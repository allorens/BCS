BZh91AY&SY��;��߀@q���"� ����bE�|    ���
)&�XKV��LlԪ��mj٥k* T�m�U���Ie�����I��MV����M���MZ�J�X5j�i���M+hK�Щ�mZƵ�ڍ[*�M�mVԵ��Z��2�4�KVYm�f��va��F�Z�,E�d�Y��e��K!Y$��B�V
��l��р��&�ɪ�+Vi[1Z��XUZ-�jmT+ -�R��B���,�ƚV���m��m��m���YB�l��2SR��mlM��ƹnS(��J�L�  �>�b���ecvc�۶��[v��명��]-i-�tdW]iۻ�v���RUֻ�}��� ��]���G�P64�i���*�    �﮵�� �W�vP��A�^�zP�h/{�x =���������� ��ڋt �����=P9�� ��� ���OM-�f��65�Ym���   	π }}7�y�� ���W� �=���w=�  w}�+�@h������|� 
7���� ��}�x �|���m��-����Elڠ�E�   n��  �_7���� h s�  =7�� ��y�޴  o'{��� |�xz��|^p@�9ޞ�  ���  zK� l�J[H�S,ȡ�_   ��4 ��i��Z :�n@ {�z�
�
�{gh�zz��j3�=(�L� �ܮ �z�F (s��]����D��B%�  u|A�p`�}C�wh�� `!@=:wk=��t n5� ,�1��ݚ������Jn� ѝ��-�h�Y6�����ط�  =�  h}��� ��� =h=�^7� �n�t  ��Gk@�� �K����⇣A�ޛ���E���Y�[iW�  �_P���  �;��
j��� �ܶ��C�q��Ǯ���{U�At�������y�${V�3�&j��k[m|  ��}��]�p g����mqF��N�\  ܫ  ��\ 9s�
l�@Y���/yO+S�iM�jdfc-���  ]π(;�΀���Qc��F@ΜN�3�UP���@
�W(��� ��   �	* �=���JUC �    �{M�(� �44��L��TA�@M �2 �~%*J �    1 MTQ�E6��=Q�4��	���#PI꒤h�SJb�қ5A�i�� �G���/�����>����~�^�c^��͜W�O�U�NB,l�h��   ��� �$�UU����Z�m����u�m���J�V�����������{m���+�~�ϭUV�|�������V��������~5��j���~3j����V��-_��\����-��k�j�2����̫|ͯ�ھe��+_3Z��k�Z�f��־ek�V�e��Z�����|�k�m_2���k�k_2��+_3o���+_3V���̭|�k�[_ym|�k�j�7̵|�k�[_3j����־ek�m��U�f�-�e��5o�k|�[�kW��|�W����_2��5^�W̵|�W�ھe��U|�W̵|�W�7�ھeW�U�*�f��m�e��U|͵�5��6�o�֫}�[�*�쪵���o��V�ʶ�̫k|͵��+Z�2�m~��[�j֙m���վem��*վf���*��2ڶ����̶�o�Z߼�V�f�kvZվf�V��Uo��V���o�m[|ʵW��־��m�-V��V�|Ͷ���շ��[o��j�f����������j����o��[|�Z��kU_3m���ڪ��j��V���W�ڭ�e�����[�j��3UU�-j�yZ��-��2�|���m_3j��W�ھek�Z�f���6�����W�ڿ�|ͫ�m_3U�+_3m�o��k�k_3j��W�ڿZ�����|ͫ�[}eW�վf��5o���f���k�-��T�|͵�-��U��>��=s{�����1T}����pOOc�HU��h*�ˬ-9I�Hk�ƅH�6��i��˧c&���.G rX����e���׏ Z�2�kzis{�HQ���1�{�+&��z��=Un���2��jbܑ^V�5҂���f+��[r�Gzj;���6vc�	&^+���5�y��6UM�F�CX4��L�Dcwb:i��tw7b���
�5�b[{����C�`-���P�AG^I�M�a��Y1�.�c����C\f��9�ܭX���tW3i�j�)�b�mǉ1P8v���	���+IyJ���2��5(Uc���%��J�B��d*�v�Ro�ĥ�t�pԵ!)��N�R�e6�84dLd��8>��ǐ��fM7op� &e]G`����i���KXtn�l-�e$]�02��h-"	�W����n���&�:3NMf�f9V����̨��$R�����D� �� ��*�1��Mhö�dzS��1;�v�I�A��j��7�^S6����f��4ӣ$�W�`هf����8&�sp��˅�^Kc��aN�,�5��&ȍa����C ���wuސ�=����m�I�%Z�g��b8Ũ�H�y[�]=�@�X�ǩ��Ғ�WG{���W��:H�R���H�#XL�x�p�q��@F��E�+���u5b �&�/A�&:vjءS`�h���e�ws���H�1�1�c-龻פj������nRPJ��4��¢�*��%d���V��W[[6�W��?ƒ9
Ii;�[6͙*d5�Um����OnG���p��$(4d��Fa�t�u,9��k��&�%��k`Uuo;�R�կ�-��*��1o�������h�k/��0��6�p���0�F��ra	��q����ynU�����cb*2��bguC�xm�fU�.�G��8��G�U[��nh�-�,�r��@�/h��4k����`�]\(����k8�;�Q��k4�J�Whư�^?�^l]��bє�-Z� C6Z�e��Z�N���ô����+�-�N-du�mG���`w��7X��T[n���7E���1�(��Vs6�)�c�X�z��8�Ӵ��Gz�<�k0"�a8��n���2S�8!3+\D�����1XYՙ��љF�*f맘�I���[l	QVl"
��G��4�MM3+t�Jv�E*�+4[���%Y+-=�*�glMg�+sI�uҤS�"�4�t���+D�SZvʹ)n�4�=��b^� �0��A&�lP��[�Hn��ӡ��2�ƙں��B��$s�4����S#ą+�r���C%�;Xw��n���Ks
8�m�%D]��aa1�f�{�x�Y��U��"tmS�V��3Xuֻ#{T�L�ɑ���ά4P*��1��}���T�fcx�Eh�
��Nnj�R��U-P��Gv�Ye	��9@� ��Aө��VJX7[jݧ�3	�9�¦f�p1{�f���PMVK@�Tw��R�TpM0�u�*0�=�ݒV��:��E���&n6.�[��p���DZ�@*��u�ōKb[�.�;��a���M�0�X�u���M�ĝ�ge��nn�h�<���d���R��u���^�_��h��ٶ�KH�w�(QYM��̍#V޶�T�7�h�⭚Ԥf���]b�6<�(�Q�N^L6�=z��`י{�&�p��Һ]��^_a �{[�Z�tKU(]Y�i��(�hm�5�cFȰ��Z������y�7�s+���.�6F,�R�Z�lV�u���=�i�z6��6�jX#,����� �����M��_<4�u�t�:B�;+ke��,����+�m�b�*̚�Ct(��F�,�sii�U��n�8ok	��'�1��!�K�m��̳��eDXl�73%���.�,;��QcRUg(LA����j��6f:(�∃�3	��X֊tR���YLޜۙ�6�E�"�=ς�a|��U�sַlnZ7�el�Gl�1�wi�X���N+R��t�C)Z�Vnfʛ���'�!� �v��n��R�J�q�Qb)=t4b��bj��4��`�Ih!�����S�[P�L�[�2��%��ږ\��2�0������nQR��{���Զͧ���K#�u4�h,ZKŠ@Bd̂V�Bm-8��#v��AcGu҂�w�	�S�ZP
K6׀!0�@�*��Y� �{�rk�Il�^P9�m�� Ӫɘ���J�w�e��w�u�}����5h��*�X����2�I.���v��P��9(d9�����P
;P��Ql���6�!!����/rkm�b�^�h[���bؗd�#c�D\e��e�Fl��(�;0�g�4h+Y�U�#!O�j;�1�[��0��Y!5mJ��A��VP*Va������rع"1$�rC���V^49R)��VQ����Z\i�R���^#z��M�*��+sP��£%���3E/Jʺ{"�"��Z�R���	��PF\��Bq"�67"��4b�+���J�5�Hn��VD�Y�eǤ�[���C�o(��b��u�&�;�t��Y>��r�f<��E��d�3n�H�D������=��\9�43����02�j��%(�B&)"T%��U��k2���d�)��z�aX�olۣ��Z�C)�����[4 �͈���J�)��gn��ha�g-�Z��z��-���]*3rc���Jb�X�C�o@uf��"�HE╕��t��df1�S�<z�8�5BV�5r���E��w35�8�
^U�ۊis*��q!&���h0e^��yDn�z-%��%֦���ViYrć,�pB+����ׂ�k��ܭ�h+kkh,Ew&CG�z7�(�����v��Q�v�"j��ԖEQ^�{��75�����*ϒ�]촕*�LB���	Y�=�e+�T|��"��mmۚ�ݬA�ѩVʰ��%�*3k�F�Pk�Y�ǖU['���c��J�Vi�r�B��Z��^��e�n�]�j��M�qZ�wJ�[�^v�U.�*N
+�^����bi��J��������[�[lY�'Q��ܥ!���A��$��2�;�w&�� Z���,�S��wu��׹6�ID��&:��f�sC�[���cx ��A�0S#���W[c,��ǿ&�����I��f�-`N�1��� 7V<-1{����"ڔ^`���sl���D��0ɳ�)�ç2������nl��^�ܔ�+4���xK�TIfK���=�a*dA\�����:Y�A�&c�N5��FVݔ V\���Yb���:fܘ�j.ia�v�#�Ö�4K*���w��;f��2Q�w^J9��k���x��oF�u��r������GjR�OM��PFV�i�����gU-�E�R���! ��Xt��%��w>ۤ�С�6Xն�Aki�DYC������.�����R�.������&�x����WY*�d�,�vws\Z�(��XG7iQLg��������tﭕ�Qˉt{@�Z��GѰ ��JːC%EA�cv��f���s�X���BR�y�6% ,)�B� ښ� ��!��hmL���G-���u�+$�2�t��Ί�Ք��XV�v���2f��-��e��+JD�%��0�\�� �Y[��l�)�e��HS�)چ��Lٸd���0g�l�y�u]"2�n@����q��	M��42d�	mk�Y�A�J�4(�Aec�T�0�8nԷb^mӅ(ٹ�Fi��e��Çk%a���v�B�FV�@y��Y�շB�PI���SU�Z8��+��vK°�X�2����hm�A��nS!��f�'[�&[_2\�z�j���e+9��n��6�U�����H�t~��]7���8�$:�����3��*`�<�:�q*��h3@#����k�NfV\Y9���
]LEY���MLo)ھ�r�l����֖:w�ݨ8�Ѵ�:��)e:GE( �j��5�����v�;r����-j������M̪�;1�-��]&6T�9�ص�]X�����|�f�О'�7HwE��$�T�f`ԭ���u;xZ#fi
`vuM������.��v���AgKe����<
��yn�ج�wKf5��@1�۠��ы#�HT�V�U
ͥV��ͼr��L�6{��^B2�F�ۃ���o���Wcz��%m�r��G/M6�9n�
���\��k��v5eef��6jӘ�7���3t�/v*�Lp����Fe��ƣ'�/0V��O'ju9��Gd��em^3�pX�I�I������5tq��a�K���bz.�ft.ۨLU�+����M�o�����=ORAݠ��f^�x��f���8��C4.���m�F�(P���(����#,���t퉍������4��؇r^5	BT�;���G�e`-�(,y� ��S;-��O �!@k�Wb��� ��D߈z��$l=5�3��R�\��b�x��G9Z�&֠���� ��f ����YWZ�h�EP��R�FSE�,i�
�Qڱ�STޘ���Sb���(S�%<���ڼ�L\l�	�)6�$�&�װ�Wx�js
�^�;��g�������f� �:�[<�s>���Ŝ|�7���R90hqM�5+��׸$"�st��S�ں
��O��q �dm$���L�aT��S%^��B�f�ݶ>wx�n�9Go)Su��f�o!�tq�-�����Q��Ի���-����p�O�$�ق��Bt�l��T'Z��V
�-�]�75�D���X)\���Ve��nS��4�r
�+�8�Al'�ii���ˆbA��2���u����bZV�)&��n����X��کu��y�s�E��0�ѕW1z6�Gi�1,,�Tua6�Ɂ]\�b)k�Lv�x>x{>�{���F��N0�&\�*[M�w@��� ��s$Z��f����E�;^l�gU-�ę�&�=Ĳu��<m3�iL�sͽi�?V����[HT��#���.R��NüڱW��6�&dׄ��j�Wv�j/����z�����tQ�4�3@���nl��.����̤y�`źˠ�*����p�ׁ��S�t�nb#�*���`��l�=Z����"��c��C8%�xcy����l��Q�w[���h�����ҩ�0e32ˌ�č�ŕ���[�j)���hA�h:�&����uʆ���4,��.���[,j��9�c	=W|�OU����j��ֶ\�ѐ����Pd�p[̆� �Ձ�-4C���Tڠ����v�\Z�V�A	m�y�;�.0֑a{�q��M"Fv��Sn���7�Ry�\�Z�{sj-�c4�4�m�$"*n�L�J���_7��
�76�yrDu�W*����y`[���5e�Pl���
��M� (�¥�$�&@@Y���̨��^jwZ�b軠���+n�6c����0�*!���q�!��֨��11̣�#NR��-�VC2m�ynB�*�V��3�t��6�v
��w@[�GQ^&$ԫ��0f�sn�(v�)���N�v�L�Yܩ�Z�oPM�h�^b�>T{�m��r���O$� l<�1w�Ѣ�ff�I�˨fл��57$ǮdC"z��U0j�&�V�1a]8�S0���$3�=�Ks��	4�:��ݖ9��R��{fV�r��\��e�1һ��T�N ���I�$IW 1U�ޣ�6��U,@~2�����n�6�^45Iu�5M���1V��$2�n�����K.�X�Yt�N��)SX���YD�/��B�Tڔ7\oJ���*�G��(,BH9����
Zz(�]�������]�6b�S~��jb�U�Ӗr��$Pڀ:�j4X@M9*_�e6��"���V�1�:�5�-9h?����Ftn�9X�{%�t�� �	�z�Z�x�:*�Ӳ��w������ZН��+�Cn�4@��a��� d�f���:#�H�k+��&�}���-^V�����-^�lihٽx��^L�n�̭X/27u�����a<(d�̄�������I( �ԴIp(�1�sdl)�d��ulh��7����ۼ��Lf�ր2P��&�\�#�!ڏ$a�5�>v�Е,m�L����� ����sPe��&�6�`���im���<'�/-�k�h�����X1=�3r��[$�	J�-�ڬ;n�S�IV��RIP[[�=��n���G���f�0�	&��Ë_���1���Z*��q��,ڕ�vKI�	�C�)���69s��ƹ릖'������؊���	+ldأ������n������=X�&��[O*Ֆ+q����+M)��Y���è�m�{�[W��b ��M6j+u\�X�`�!�yh��ݤ� 5��閐��u7��w ٫70(0�*�r��r�Y��hcN� ����tv��A�ܚ7~X��C@�ʈh������e�G.��tkZZt�(nhc�Zn'(T���{���ĕ����&�j�,}}n��������#h]:\�Խ�^fiqF�\��68��3y�,C��/%�璻h��[a�7t-�H��򆲦����[vO%�N}��Õ\�\��c�p{E��@���z/gaұ]�h�/)��ك��eu][4���+tǢ2��'	������+2hY��#�3� �����`R�l�=BW
xF��ۄ;CQ���讖�E���ԣ��d�c��.k�`YO�'��p핀�`h贛¹�/d���`��"	U�Ɓ��,Y��5�$PF���;����q�m�ٟ,��m�`��[�QV�w�������F��?�ɏ���}G�t;��s��]�j��i�tpɒ�kʁ�T��iz/������v�{��$�i��;C|r<�U�6����E H�>�D�uV���7�nY�)�-�R�E;�Q����x�v ��├׹����L�+lo�3]�/�CQ8'Q�$����l���jbn��Ϥ�`OEƐT�̜i�4�`�OT[���Y�DcC��97�7V%�J���x#�B�Z�O��v�n�D��U���zR�JS=r6]:��\���冷,��G՝L��gkXD
�Ӓ���[x����uXu�WŅ�j�y� sU��gA3e���ź��7 Q6�{��U���5!���{�@2Q�@��r7��X�;E�OAJ?-���s��84on�����<Ki��eXô/�Z)0X������F#�]6��5���g���Pp�����z�q<��L8sp��ar��r�=*�n��m�"�T1����&�8�3o;2�̋-ѰV��Q� S��B7�K`3�{6n��k:
�"�S�ء�u�Tn�#�Iζ�-8"㕋�^�u�56;��6�:��˘�oH���j�;v�pQWKl�>vt��ńMÒH5QL,<Z�ky����(SY�ak9h��w*��n��_D�pA�Xf����{�k��d,2M�1��q�����:Q�P��]�8�rk&�[�ʲ��)fn7C4��;�l�W5���Y����*�J��ގkvt���[2�������h������4'ϪPޒ,������"ݖn�Z%]��P2˽�s&i��3V����Ѳ�؋��vk%

�0T2�ݵ�#�`�4� &j��u\R*D7�T�5��S�]_Y�5��^n�	b�Ww^u�#���vK�dV���Jk{�r��(�îV��C��h&����klK+4���@e�stT��ՒS@qj�4[9lcS���=����^�#�Q�ٶ����[�f�Yc��)1f��v΋�Alun\[ՠ�n%Dwt���q�t��E[K�`��Cak*��]�S,�7O�Y`I$�[�Y��NM�G,�E�Vs�TiA�Z��zh����*D^S:o�Mکi��������Ө�7.�OAu�,u�X9 ��zR��g�������h��3�̦j�a�$wbGh�ʾ|;�%0{�0��/g;l�P�t��.f�ޢ�;lݫ��m,S�5ܖRs]��ժ�|v��0�'�P���O)R��[�us��4+��-y��j���J�r�������&&$ֻ-ؙQ��ϔ�@
Ίv��z�r�V�k)�$��Tݖ�񧪑�2��g,틔��/3Mӝ#��G^�|rP|�-婹vj��f��j�l�&b�y�����.���b�y��[��l"��N��;��oh�48��gq���2��"��I�=)L,j��Zo���:�an!F��o���\�wVż���� �߅I+vV^h�g!N�\����݂�:�\����؛k+�
��FX�V#�C����x��F���Ɏ��ȥ,�������4�t/@�xW��������Χ0�
ɖ#O�r�H�Ԟ���-?7���;B1J���t�g���+e�(D�j�^��������^ʺ���׷�Q��݈�)I�LI�V�#�`i��:I.�43�2����94VpbF���_]3 "��J�t+��VnW���]Vc��v��Y� �E*�F�,*b��d�"h�(h��=���"�:�WJB��)�w6�)�ZP��@�)���r�V��=�eaI���Kz�(v�ma�@�j���{x���)(�nQ���tej]�<a�r�fv
�e�o�6��N޼Ѝ���1�f���[j�Z���7�W2�����&^�z���P����ò���-���i%��5��a�0wnku!�h��W5��n���K6��ynYN�z��m�o2�$4�4`���&���p%k\X5��|�␴��1��k��Y��_7���m�Ũ�Wr�u��|5 ]MO��βK��
lv����#���������>^�{��2��`ꧮ��م�c�die<.�>�У4;�`'u�j��Ӧ��f��W��b����-���F�]��ۉ�:N���v�̚^o,$�#\�@5���c�h�t��08�b����-VJ�{�,^yHډV�%����bܾ[יܕI��v��}��1�"�%�Y���f��-L���p)wL�t�K��i�ɴ��ETrk�'&#�|v܉� ��#-G�2�b���8��N�g���,�RN�o��W�M�^�i���Vo �4��&]fy�����;΃`z#��A���.��ᾷ/)S{D�[R��8"zK
�?dʙB��PE���]��h(��y���ĝ-�DbZQ�7��n�S��mp� ��8-�m��Q�u���O�Aш���uJ��LQ<r�$�����Z�B���K�|%-xF]�3(�; [�v��x�8�9���>���[E�';飃��V��*e+y���9V30�]$2d`�v%���2��o{!Y�_	Qhԕt�Q���8���:L��z;0c�W���sn��Ñ-R��e_U�ܲ�J��c�m@�Y�8�,��YW)݅��J6�5���\c\�;yt�``�2�f�A�vR���T�j�d�%0q�u�
[�;ch��f}S"���",� .���z�_ko�>T�S��2sսY�Xn���ծ���� ��W��5e���=*,�6]j�݄���:�D_g#!��#�I!�����:R]ˏٲR9��* �-��`5�Br;�x�d�:�{����:�T��t�}�v�/[����.�*���k�+�% ���m)�]�h>䚽�}J�u�i�t� 	����kՠhT�t��V�i{���!�t���+tl�V2�8�8�rY�bD>f���e�L��;K��S�!��W-9���g�m��A܉Q���&gթE�Z�۹	�����	X�'vb�q�w*q�<b5 y��moV(��S��F�[V��r�R�N���T����Qre�}�.Z��Տ��1�p�-^ZXP�mq]���Ǜh!��^��X��ܛA(�{3�?C�"�z����.�m-��P_q���0S�.v`��Q��]��W[rg�[n�3��^+1Ӷs �L֖��X����"���H��ƬfvH�:�p�jt��Bk.���i�m�\������;�j���2;���N�A*g�*�X��ƺ�Gn-�ڽ�=��Z)W�`��r��B��㔈������W��%}���"&F��c��ٻ�G�IgfuC��:�4�EƬ�4��`����B{(q�=G����0�۬J�Sn�^��w�DE�բEKEZd���Y�>"�@�ZB�4�,�ʽJ��[Y�;	]%w;cq�)d���T�L����锩����Q�1��k�[���Ut�$9�J���/3�9�U>�
յrޭ�z��;��$�WuȘ����gs)��1���Unq���-R������.�SX�_a��skhdH,�3gn-�#�-��i�%�z^geQ�M�X�ƻ(&�+��:����Bp.�Z�=���;ZY4�j���O	�Ps���:�;Kد5�Hl�8+w��>}mm���q��_e�I���+V�' M�ҕb��J��f��=e�:+��2m�m[ә{�v
r�m�.S>�n�
�p����6������t�d���#F�jqH������y����,wׯ��x�z$��^���wj3���Nj{���S�U���9��sc�e�c9CVݦM��T��S�T^w�s:�J��|�H�9��ي8�����@�/��"y�������8��ˮ�����i)���%�0���s��#m�խvB�����aVw<��~͹Y���L�bx7�h�t*f�oX�0��&0p���w���E�b��qY�=H�;��{@���@ax�"��"�8��/��bT��hY�����l��f�|�p]լGM5�KYeVFc<fұ��;d�Τ).ߺ��p�1�m���Ζ]vu�e���GT��0�<�ٓ�>��:�T��c��A�R����r8q�����V>������n�b�5nΕ�G��'�u�RU��Z븃�a��X,�D�,�<�����+'0LP��bZ�fb��{J��2<�2���P�ܩp�4'����*-�Y�e��G{��j�*��O&(4hU�L�y(:��-W
�"��{�0oUٕ�t�L*ͩk%[��P�ՏHbd��S@�YPr�:uU�ù�b�WI��n�*�����N�öR��
�bi��g^��8TOrgtиgϤRrpS��# S ۻA/��ѽ}K*��<��E��Wqה5�q��`r�[��T*�Z�(�k�Z�ٺX��#AR��rF.ћ���\���յJ�� WWG��dt�W�H��T˅�)^2PapEӉ���gS8���)�0�����)M�v&�&�K݊�S�o�v�:w�����ghFZᙁF�^p���FFf%�+h�k�Jhtަ�]k�!*�C���L�9���m�bs�eb�\��1)6M�N����P9�(r{�Шt�5��l�V�u���oz�e�a�#���Q��]�_�K�UԳ�����W�̶�Z+b�N��g�jXbͥ��t�)�C]�)M貖��SYL�cqД�m�\�Р�[�[V#�܃�D�p;i�F��Cw9���&�Ϙ�W�u�ި��T컗4:�;�S�1��g~�6�!C0Ê^�=��Y2���^�i)��1hq��w7e(F5CHi:�W����\]Q�o2��Q}�v
U�K���t Z������*��-������j�k!]��3a���j/�v�q��w��U95j,��B���s_w	�]�S� ne� ,��]��zn�Ȓ��:��Qitd�ɨ�Dp+$���K ɑ����'{�xp��Uc��S\�L�l�&f򮼔�Q�\i��:p�r�T�0��LL��]f���hK��S�%nT�k*���f��6!�(��;�r"��͓�!F��豩Y8��j�����6I��
��8��q��)�Ur�3׊�l�4���\��ُ�������Q�P���l7ϫ����$�([�"�MP4~�9e���b�r�Xo3/5�6�I1;�����M#�Qr��b�VPI�q�%F�W��l 3W^���Ƈ"��۽�\I�3n�։9s��>�XGB�Ӝj�7)u
�]2����3;Tih��f4�.`؎�f��ju���푻ئ�H���eM��1b}�Xl�sרGS
�BS�<�s:�
]���u��<G83صf�*lY|���-��z�"�뭥$�瘸��x�L˰�C-�}�xj�����̵s�F�P����"l��:�`��b��x�3V���f낺S�U�ݭ��\Fn�M�0s�25��E�<�{AΈ�{��#����^��+k�:��z�ly�p�Q�8:�!��&�^��x�5��v�2���6�7`�7�a�`�k��:�,�M؇D34���M䃌���,�N�]b�β)�	��"�J�ھ�-�>���pK��i�&�U	�V)/�l����SP=�^#Ϻb&��8&" ��Bc"�l���6�7
�� �@S��ƛ5��g
�MB��Y6�~��\r1|(���ʅM����=�w4���~8����l���rF�FdA�;�mnt�����X�K(i��l��K:�bk.��:�`<EG�oR�ee)g)Q�AA�2�Bu�o���ֻ$T�d� �v�Ф�
��0��N��֕!�)�"�J=�+�s��}Q9�N���wҌK�td���y-L�`*P��6HJ�ѣ�����
Q ����L���d�M���5�5���ə�H+PZ+�Yux��8�<=��u�ܤ҆@� 7'�q�,X���o`ŗOm�9X3p-�����E���=��
�wf����C��O
B�jr]\�*R���rT�g"{+v��SV��(�-<�i�j�?�<���5Oq��6�v�i����2N2���-�.�̽�Q
�9���D��6M�y��iՉ�Lj|�>��ʳ�zߑ,��ց����9�mᨖ��o��ɲ+x1 ��!$�x��k=����4ƺǻf�u(�5�mjf3c���x�˨^P킲�b�w{ek���K��s0V&z#Z��k�wW�vGHpt��\�v�<��9�D�̡�=�L�d�)�U&��{�����7i�ǉ��*�������V��q �E��c9�rY5`n��H���W ee��4��
��]w��v��;[X�!�Qó�������a �MM/�&rG�_���ꥂ�i�tѲz�Դ��������#���`"J4�R��Ƨ��!<x��!p:����'o
���h��������r@���[�at������k2��NQ1�t�Â x����t�ʈVEsg>�6^�zкP�-�)CFv8�X9w.Sܤ��X1�%��־r���댺����W�P'3�8�ϒ����\샤뾽�Ak�P���Y��ߘ��y��5է��T����N�ȘM��[����{r����T�dy��ֱ��
��M�wp��=m�+��r��׺�fl�IGx�Rl8u%��%j�flk$�2֡{r*�)����L��.R��S�)���k���
@�\aEy��R͢�֕	Ub�9��LqH��_,%`��J"��MR�eoR�Y��'҈���Ƴ��1@�"�Ll��wMܺB�
/����
��:1��&]>[&�'fQ&�kWt������)��(艘y��靬I��q,�� H$�~�#�~� �  =~A|��P$~��H �	�������,���}�X�}1��4�c��cʺ�����l`-�월V��Mm���,ML���K�r��̬G^�������ru���5V�גܶ#�;5�*P���n�фVń�ܺ{q��1�G��3%M)akބX�����G�YY{b]9��k��C���s�Z�yp�<�J����xx�36�q�xYV���퐥v$J��UtLわj��S%u���\��.�kv
�E��� ��B��HE"�]Kz�&���,�k���zê�Y��d�-&��x9������C{�H>&��K7DM콺�8޾��*%���Jf�āL�ul�B�t�&�]��T�z�˕���
QՎ�2S�єD���"T}�f���A<<���`��r�npX��f��՗)b��N�T�@n_f��S-���B��+`�;eh��3q��K������Y3+wR�}��IROpu\�)�S9��n�É�m�uK�����T���et��6���L�q9X�*�k�N��R��T)i���x�S`�9���Ρ$%��b��8���p���Ƒ���A�GN��j](B����AL�tlR��,7nӁZ���w���YiJ��Pl���kX�s��И�t������
��^�f�-���sGJb�`��Y@ݫbT��,NXc��ۮ�mT�* ��Y0ʍ�������[L�а�ϑ9}�.Uͦ��Ε4�3q��pW�,�d�-[��rc�/h�ǔ�:q%{�U��f���{��[J�2�qc@�f��G(���w��dԕ�3qR���vR��;�P2�7m�p@C|�䶸��& ot��u�kCE�Ô��#����,9����R�j�5;2^�V��^03�/�:kB����=H�.�k9�+��]S-S�9�e��fi�#�B��9WF��|`�R�Nܴ��s�A�j���w��L�\��/��C8:�V3,�-1V����������p<{s�S/��q��R�V���9Y#�hf�yH��q�YH,HA��cH���h���*��9��3dko#9�����N2�,̻4ZI~Չq���j�O������@�p}glB�X�mn��֚��^�(G���fX���9��!������Mh���cpP���i�f��YYG$jMa���1�:��&�����A�&ڽ��M�2lN���A-��Y�.�b�n��Y���J�ӗ[ ��R��:n��V)Sh��\��LZK���b�@�c	��]g3�v`J�waF�qgAhi���Ir�J�kݵ�������P�:I=(�B7��l�zUI���Zet8�;�h����������U�uؖ{�ui}�x�jv�
A����bÙ��ϭ�Ed5ۑwV�Na����U���8ZK;Vҝ�TE�n���n;@�ff��<\�z�&���5��l�K��'ɵ O�[1CSu���MĮ�Ͱ�l�p�1�(E|��\Yu�~,���V��SY����@� �7�ו�Ev�����R���"	�9].��7�,�����q\ݩ�yI]f^��J��� �Ε�R��M��v*���:�ykg;�x�(v��";���.�� v��9vɒ*�qT�#�Υ���rI���Y�+8���j0������d׋s�1"
�ŭ3;-ҋ]�����N��	��ˈh���L����c�4�+LE�wjd�)2'��19OMӧo�TL82���sIKV,О��aR;�w&��ާYK3�p�}L�,bغ}��ͤ�M��9�Z4uK��^p��ȫ'_{�N�I,�-�Ȕ�U�!)8���
hn��yB�����Q �x��d��FJ��s��K���.$��x��]:Q���]����6������6� ��a��T���Ҭ�gM�.�-�ėS��rɓ�h���^����M��`:*�b�v�Hn��Eq�z�0�6��Ç�H���\�H<W���-fS�O������Y��Ա�N����U3n��M���:�V�����<�r#S��v-�q9A����p,��ζ��_`��rҡӴB��Q�.�JhdA��>��7�x�Mc�1��z �ϵb��ԧG�V�����uBU� ���y8���� /sm�_e1z���H�d%�U���V�@<:������P��*�&�.˭�96�4m]*|���1K;f����1�
�2�n*��,�ϸn[<-���++���	�Jt�L��v-�{Y�`$U4n�n^�z(31N�T&jx�p�tu�ԕX�X3�Ν��HH��T=�F�+���k��e����:9c�Z
n/Tu�Ҧ�Ue<�]>���m:��;�Z"��9�]
�n�#�J����")�i�@���w��e9��`j��`�(�iR.�F��x2�~S�L���nW[�dH[zz�Y�+	rfeHZFc�Z������o���g5��ۍn�yZMw�a
kd���ˉ�ɦ)��Sx�,�NՂ5�p]&�TE|.	0�=O�W������n�l��'�:TB��/��7�]��W.�=fE��-#�H��o`�t�N�ՠWE+�]�˕�MRy��p�RSc3���R�H���릯Pr���(��)V�1c������U��J�m�ZU7��R���[�k�N,�H�����w��ql��(!{�L��b�t(*Dk�)��cB��q]ND__RH�h���Nk�1Kݬ�`"kx��Bކ0�@yԻɩ=�{ �^�3nIS˧vS�[kX{2�L�}�B6�W9�>��m�密���r��g
�вvC�e��C'-�ksh'.�%�d�sU�n��}ǦB�Q��RZ���O-V����]5�t�F������%ը����k���a'&�pm���Z�'9	(sK�1�kl�����z���k�-�
;2˲��l>�}�Jri��oM�@��*[�D��9�̶݌�ʌ:#Y[����!��l���Cp�E�|�b��	,-3]�c���ݣT�W�*�퓇[�����ʜ-3̈́yd������0$/wRٓ�J�6H�Q����,T8܈��L��ۯ�D��1�z�V�*$��8/��K����������ː�|V�X�
�lSE\{����֛k���d��v�:T��/0ޱH�ߞo���S�"���w� ۡ��`-T-��`Cy�4�i#]��9�����Sq��l��ԅ����o�`�A^�0�\�l°l�;6��y��s�9�\��r�6���˻/T��g�9{[6��hPtVA%4�7���6��4'D�L�WK;�ϩI�P1���)Wj��:���;��(�ow��ܮ�����0K��1�J���|C �,2nt)�]�hcW�+�gXF��,&j�+���Α�3`�eSޤ����`����2S��PA9�w�� ��g7��Z#R	�ڷ�{�����L\�pD�f�ﷺ	�[6,te��\qWfk貘��V>즹�ɠm$���eܜ�:��Q7]�֎<knt�����Z�އN����{2����cW@������9��QwJ�'v��&���#�c�����Q]R<��pa{���k*�Z�E�O++r�l�}\�����ѝ�.���I��wJcW����h�'��%������]���Y�V��~ c�=Zk^R�9�P������ԗS1m��*&��	�8����+&�K+�6қj4���cV%<�7��NT�֗AP��r������78�un��;ir��$E�&3֩7{M��|���S�᫼�s�vk��k�2�|T�z�,�V{_.ʽK*��/�E-N�
�	3ǲ%38T��G%HQT����a�7	۾�u0pL7XW \�s4��5o�g]1�M�hY/��[�Q�xU�{Vr绬���q]�8dfX9̛��s;y�s��a�o��d3㷡Ԗ�5�;:h��?9� �M��9.�f��7-�4��@,�}F��m�q ��m�g: gP�v�
�*�y���H��Q+� `�3/'IeP�f]P��� �v�T��dE�/�G��MŎeu�%��Tz�0����ݕ��.��`�ܚ��8Lò���˨JA>Qc�9M��*]�c�ݔ�U�Y#��ԭ1�m�}́���C��O��3o���F���(�Zj�h-'-���AvA��Cd���7�ɵ��޷S�J�-b�(�z���8x'����1��d��֨�˩�m�5׋-�����9M����j��<�V�9�Jo6�v�����kK�<J�G���\W/y���;rh�՞R�5�5>#���;'!:�R8��}F�i��'xp�F�0�J��k��xߴ�vs�Xw�a�)QN�I+�����/fK�)NQڅ����Mȸͭ��Kth�x\�<*(��(\y/���}D�Ghײ���c:ˣM�X��J97�G�Z�t�K�r(�M��k�(�	��V�ȵ�
̤��sc[�0mJ��*4�4]}��}t��y�l-�[��\��4�*S��7@C�v�ND�\.m�՛tp�S����R��6�Ǵ��IfKpU�!m�^Έv�Ŷa7Nr��������0I�mj1s��w�rJ�W���Y&�ۖ�� U����~�T������B��s��b�$���1W9�-��i����)MG(,`I�����9ق��;}K��=h5VhJ�ڃk��4WX�q�Ʈ���Z��s�ucf�\y�6(�_we�c}A��U�q��y�ˈ��2���/�8�6y� ��s�.)v]d3�w�b�ʛ���rf�b���#&�f�3�w���Qa���O�*�Muojg�%l����8����iHj�O����U
)VeU��%0�d��>.f��f0��"���ҏe�(H�2��=C
����U�b��]}�\2��l�u��q��҇*�U�}r���w1�a1�G���V�c� ��o����u����Ƴ��i��L�s����G�7At��lb�.�����Hk��t���᷿c@�/L(���ZӐ��2�a�q��2Xl�@�⃼�2B��T�s���Eep7Nͦp����Nڿ�e�.%j�L�WqM5�)��&>���Vjh����m�9��y�rpn$�}ۘ�F�U5:op�:M���h�9	�����\[��D-�t"����u�ӿFp)���[��n��3A�{��M�ќ�-�,A>�1Щպ;r�oi|�Ǖ֦�GD���*�`�q�ӟm�VxcJg�X�D��i�Z����e�%�ԲAR:�%�iWf*�E�kQi_�P��<���#5#Oz1��o3�o\�{z�)g	h0�Y�l��7\lP��N����\GH�`�� quѧ]N�`r�$Tv��j/���4�O캝��H�	�kH��0h���:m�ޔ���2�F�c.V�j`e��I�*)����L�Ǯ���
��g�%;�b�b=Z�s���(;���Eove�{�/z��	��������X�s9]t��i�T�����i�����.l���zATt��XD�3pv����|uC�8�G�-��p�%�tG1�WP��Z�-�}��*?f�&�DL��?��ye����uL+��pqGK��ӊRӅ�KE֛V�f�a��4��]@�]�XLEt�(%(�)�;�	���ܾ�7h4]�7G熓�� @�T���i�sC<�gU��iܽU�{.kpf���7�*"�rM���;V�b�����!��-��4"�`�������.)�#Sա�B��8�J(�;[�3[�j�U�AuwmBr]�C�e��,8T+2�C�s"�u��"B����B�1���
��Z8�6�rr��,�e�Kj�g	������t�2l�ȸ3\��Y}���O���\�m�1:�T�v3�lY��Xp-]���L�^�3X��o=U����ln�ko���/��+U{��}Y�}q�9ى��c�g<�ږ�F��ز�B�=�XĢ�ͮ�?k=%	��5v���V���U��Ӻ2�ԅ��x�ү��Ό�yʏ<�/D�&;6�y]�!��ۧ�DL�����\^��wۍB+.Ö^�7�IT1�(։��61:�W��}S��2���6�SP��n9���2�� 9�C��~�F��+n���}Y�xV�4 +U��,d��Q���o)W[��%Na���K)��E�:,�t�c����,i+	���",)+
�|�S��vMѥ���oS�n��J������N?gQǃ�.؃VL�s��Y3q�i���U6G��8��J�E�y��8r㨁2	ܖ����k�ݓ�Pʏf����<�v�?���;���������e����o�b��,�Vb=D[��T��N2$�Z�I��8��V��)�����!4<��Ik5��Yƶ��]�#{j��%����'X/�3nZ�;Јvyƒ�}ЩN���PY��XB����#��<4.u_c�`�)2���d��8uK� � ��t�'Y�P^`�/�1]7X� F�c��h��/A�õ��^��@�lIur�
�)�l1��DڎKn֨�I��QfQ}�@f�B�����ă+�s,�8����=�ݜ��*��-��	�
uۻի7���$�bʫM��!�52eѼ��{5���;(�;:,\\�Pg�Ői�#�nm5(jmڮ�xL#�Xe%�a��Ɩ��Ѫp�-�JL��*�Ugrvy�z۔.�ŀ��+�џt#;���������qH#]����U�J��1��D�7�7{H��5�X��C�,�4�((B�T,S�瀇v�u��u�a`H~����I ��)����~�����?yy�?C�?����h�M�6lٳG�:Q��^DT�d���'��ك��{���'�{�/5�݄�U�u�`�ݤ*`�.s��XL�d(P��ڤޙ��]�G&�9&���H�v�\7{WN�O�V�̎���4���`����E�t�iJa�Cm���va�]�����1wo�rE�c{�&��T�������l6�h|$We�J�'זۭާ��v�Z�`M'|�.��,#��ujۥM������ÜHؔ��3{;i҄�S�;8̽�]��uQٺ�$>�*8zgJ����PV�I�v_Ay���eխj{�,h��*m-]R�V�.�dƓ�ay��n�^��t�X4܁b*��N�S��I7��9Wt�];ʂ���3{�"]G�wς��kn����_�S��X�s���%*�z`\�Aq�֨�a���&'��A8���>9���g+ٴ���j
�E�v���V�Mwc�9.���x��Ķ)�+zʄv��/��f�9�>dd����F=����Fik�n���z�3-��}]]���ʲ���+�]�y�s��v-��k�8����Y�l���,jrgS���'�/)Zy3�d����D���+(��W��ʾ��/�\��x�U�� �<����ή�®=�VK�I�K�r��O{�wPN/3R5cI��yt�	�oX?(�As�/W�t����b��Ӕ��x�v!���c��s����:B�R@�(�;n�X�ժ�6P�rF%՟�tꋧt%ƃ����	Κ���r��.t�gu�ܱ�\ӻ����]ww	f�(۸��v.���ru�E�Q�w:nrw]�+��������u��u�v�Ѯ��u�MC.����k�wGw]����{�Ӝ�\��N���.;�Eٹ�\�\��Rt��w�F����u͹w;���nq��r�w�n��u�7wNu�n�K����΋��7\�9�������st��;u˓�"�뮜���K��ss��w3��;�w]˘Nw��κWr����˅Ә�!��]wt�w]݊N����;��.���t#���#3�܉��nݕ�rS�˹�Ίp��c.�.JZ#s�!3��wG:vN��'ww;�͹sQ��:]1�q17wn�s�t�h�oοu��v��=%#32�CU��ԽԞ^n�Z�V�g^�]Q�^�z�罺�q�.���R^�Ψ�7�kk^3}g):�O��Ӯ�po>k�L��4�T3���#��en^������~�^�q�kfz�D�On{�T�iA{W� ,T�Vy����<t~2RW�1�����e�x���B��(e};�~��k��u�I{�}�h�;X}�,5'o������<�W��a���I�^���H�JK��ޠ� &.����ޥ/���R����IeJ��TUҳ�w�f����٣�\�w��VMf}�_���5��?N����dh[�uw��"������nhy�"o���S�vy���=�����t>����)j
��Nq.��T��B�r�c>�Y6�;v�������|��ݬͺ?�-��֖T�����yڽn?m�P�[S��؝V����W�r{?�D�e��CÜ��t=�;��t��z����y2]S�~g��m�[�;�v���%��	��c���c���7VU��)�p��*fʫ[C3
�R��wZ�s�&����A�ܭ�+;��u�����Ciա�B�����8C�:�-�d"�Ѣ�Juv3xK��=����5��q��mD�*�#\�F�6zX�tì�t���s�9}�������eJu-W�]6�_�J�Uk�wr��2q��!�V�W�P��)S�S��V���e<��WL��ٿb����mM�,V!�[���j}5����ButH�[����u뫀׫��'�m���yM���͠���R��O�gl��Z�:�ޞ��� �~�L��p[����v����q�/}u��5C��'<uf���{�g�����{�L~�ku�k��1�٦�!�E����ɾX���L�o���|�R�=�ѻ�ۖ���#����l%ٖ�Uq�h��J���z��3Tǫ�7�:��Y�t�{����Ϝ�{����d�Ƿ�}	�M�Ҽ���+(^�;��'�Ar9+�ք\�>�+�ʕ\�=[�eV�������6���/&׻��򆧵���g�{�U��}l�]���l?_Z˭?�M�bn*��w��-��K<cmw�#�K4��٦��SP�8Ep����5(�[;�fL����n����Wʄ�a�Z��&J���U�ۣ�����CU�n���Ӑ܈t��8VV��Z�Qf�����/ǹg��\��R��M�7�m]��G��̫�jpn��zf�3�H�ZkU�X!wP[�k��`��Tf��C׼u��¦�^�z�|qvű��ޞ�wxA<����<%ז{��\���gmF/���v�)����N֫�	����B����^����ɽ��-��n�R��t�N]/G������<�����F����Oe'5_-�b����u+]S��V�U��_���<�%�p�'��+U�A�|���K�#Ԓ�	L5�]�Sj�>T��^X�D���N���f������~Ӟ'�**q�E[�n�ߧ���G~ؓ�5~�W����屹���d�$���*~�*���#��;2z����=S4C�0F�C�v��U�����.�
��ⶨ��"�\�Hr�>��{�)�6;$`J~2��%�O��^��hˌ�.ث0E}�֬9vwY�HM��8����\1��bˏ|: �q�ӧ@�k�-���<����+f��R�:��3�f�Æj�Yh'-���u�á���on���;�QQ�/-'R_�����}=�IMl��x��K���WI��b���f�U&���y��t�x�y���U)u����3�Ƶ�\�����=+;}�}���o(�Z�r��/f=q.2���vQ:��fO�C}�G�؎:-I\(_/PCJJ�]$�Z�y�;��9/�6=����s�c)	�:�G	�j�L���Ü��5�<�h���u/�=JK��s啤y�
A����:�t��}}IN�\��U��W���=��ҷ�����#Q�~�o.��� �;K�z볔�U�ɬA^E���k�%"���zO4�O����}u�~����&�4Lˮ��S�RsBo�ǧ�z�73h�g�M&n��R�ʺLl�L�<C�=�0�w�׋����Vr�	^�-^��wZ��[�hu���pՏWe,�|����s�V�|+އۺ����^�W�=���Ɍ�G�� ]�;"�l�	/$�Q�VU>�7���Iկ2��N���֘Y:���듓1�>�N��1�jViˆS%[��gU��2�L<�@"{7�p�t7�{���#3k'!Ke_GWv�ӥo�s����٬5��szD�l޸N�rO�m�|_ h���E��ET����Z�fi<�WJ�hu`����Pw��v�N�\�F���=t�{/0�Ï�����I�鵨ͷ�/��U�>9t}ֵzF�V��ʲ(elJ�=�Dn�8�k�J���|�i�����K�S�F{�m�v�����[Q�Wr>�g*�N�x��z�����6UmA8�	9u��ޤ2���j�9�aEmq�5�<�/W�{������en
75��f��u����1(O]YX�I8�5T�i�z�K}JUeong�������2��=G�0�>�Lk����.`$/xu��x%|eu��Ηc�İ�g������C�.�QaUyYHa�/G	�s�{�%U��#+�3/u_�ֈ�{z��*K���l���T��y�9P�]+=�!�����U�@~nV�����[0ד�uu@�(��H:��=1��ؘ�e=w��nC]Q�- `��"Ř4L�#}�z���U��
��\x,�|�S�Hr�z�c��gZ�E�&���u�Rq��0�8/�ݡ����q'F�t�&f�.�D�Y�3�{6�7���)[8
��]��aaN�`,�0���坞a���9�'��>ˡ���8�SYGQj�������I���ڬ�I۵'��s3Ϳv��ۧ�����z�}�8�r���+�@G�yW���\�Z��w�!˺�½���h�����e����5�oWҕ�O��62�͞���k�U�C+����;~�\;29��?SF�5s�S�yJ�2�.����T���Y�
]��'�U����Ƥ̊����yb�PR��C=�!��=�t{<s"�r���(M*Ŭ.
F{�ڒ	=�����.G���a n�>����{��4���i����}I���J�ѿy|�C����g�RW��Ӊjw�yw���I�����W��d�'�VmԆ����
�Y�_%މ�N,��ڸ���������tx�c�Em9zmx�y�K�ޯG������]�	�F���5x�{��1�_h�z|#������5;P�7�Ad	K�]���"4����^���'k��k&�u����@��X}4�խ�b�]�����M���s�w�������?\�u��S�"QR�8<4k��Vd�&�(_W>�A���t�{h�b�̡ug� ���+*RoMgS���q8%xﳛ���=BZ��S+ٽK������{��˹����1�����mv��IOI�c�7=����^��j߇]�+@���^�e�ZD��V�L�x���'p�����f�T��d{�%��.Y]�w��\f��r �؞
�K����h�$X?Am}>ѹ�+��'�妾�kP]��јU��*�*�=���B�6@��D���>��mn}7��N����r�^ߛN�c"9�<@��N�Sv�]>�Rj��'�{iy��}�,hX��=M��ڻ�#~����&��_���{t򝿅LJs>�;kɅy��IM��_��g�G���8p��%YL��ݕO�T�J���Ž�=~��8�(��Etd�7k��v��K��a!�IORъ��tǾ5��f��^�;D���_@�./��x[0ۤ�ͦV�lN���6T;\U�`��d����_u$a�K4��G���N������JoY/T�A+0��}S(��:��i5z�utH]�Đ)_mI3�$�����q�uq�@��n�w�WD�}%�}9S�Q�ܡ��q*R�M[˫7�*�л)��C�V�u�����S����恮�}O�^��������$���Ye�BGz��>��:�����gq��K��ή��ay���[�@
�X��q~�D,Vy�����޵�.�j,vX����S8��4���\�ڽ��]���ؽ�U���vC^���m�=�:Ϗ��JNU����Gn\�t�o?VfDe{�ɟ�,J����o�����o�v�]AG��c͂�f�����7ݳ�Ub��P����h���4�������=>^�8�t,d�b\��~�i{�c��<d!��ߒ�t/G	�s���Id�߾`���M�aʜx��%O��N�s�UK9�L<<)�m�|Ѱ+_�׆l>�>������_����}���7ꉄj�,�PCW\+��(Jl�XϦ������VYN�����(����#�}ֶ���K%5]�`�[.�<fjRU���;v@�p�<8Y�gz�d�@��2VP��QKrh�-Y�(�g%v�v�Kt�Gɯe�D�x�"���:h᠒1hU}[�bi���B{b��wU����e�l�s�"qj�=[7�6��?z!(�?nF}��d���{=^�V;�¼����Ul�������4�?=��������X	R��7/���TҐG�����=�u��l�n-��p�K|���k2lJ}���J����}E\F��z{�|��ұ1�vzJn�hr��1tժ���\�V#��:<�V��$�7O�D�J5�V=\��{�K��d�P~��J��~�Y~�t��O/N��S��j��D�G�����E=F��^�v.&��h��^P�\�O��޾=w}/�ƛ�fG~��ߢl�)��;��S��??J���y�ś���3`6�n{q�3�.�'�w�߰����5�<�/W��������}��D|<�}���<�J�N]p���O���,J�S�o._|�W�<���Hɹ��V2���kŚr�x�c8���<|�mh�����b+�R^vd�xd%��B�Q�}������e 4In-��]c���C������k1��"]"�m�p����sGc�4�.O"z���Su�:����<���<�Y�s'u��s�%u.���xr>�V�����;bTܠ��T�&���z�����W�WJϸL7�1�������N�Urݡ��.��2;!!�$�U���?nv���X���^^82k0|w��_�S$���6�5{��ueJ�^�5�TO��a�H�#�Oc,o"O/�t�T�2��~>�ﭚ�~�a��7�Z�z�]���Ǧ,��z����H�_	ŵ�uל��_-4-Z�]ܷ��eЊ�K�=+�Q��$>����_������k�rl='n����O��>����L�U{�^�7|���:O�����U��>�/	޵���^��7�kº��'M����Tr{�i��#~ѱ !�t�G��G���j��(���1{n��]oYZ��ry)缷���[�벹���V���TVNt�{_�Ql�1�i��ҝw�x���<+��Cu��;!k���n $��:d����6lٳg�����Cj5�k�B���E�f��s� 	8Wv+=�0s&���y[���Rr�h�r���*�i�D�9j�؍)I ��':&�ی���6+����-\0�ۤ��#r�x��Z��(�y2�<�0���P�wI�Kq�γ�/�s���68��ٙ��e��&xfedV2�n-y���Ϟ�\��ys��7��cI1#�����nQ���P^�ص�̛�e�ԣ�s�3���yL�ݺ�㎮��]�6�i�'9l�otsjvL���ʵH�g]�;Qu`��g�c����g��<�z:u�S��}q����1ѝi�y/����M��ARō����[�����E����\Պ�h+����_Ϥ⮆���NC��f����8�=��!�X��N��0�L��'[\7�Y�{��.���d�=��*��'�(݋���kY#$��6�{�I��J���`���5[�S�V���(ӹ�C��Gy�6����P�[�p�Fk�&��z�u^�U�,O;�TAu-G�!8ȧ�ń����J����;>��)૦Պf;:&廎l<�x6ҹ��`���'P�k�'ʄϢ��zJ����X�H�,��<���d����Ht�r�j.�`;[��iE����7�*�L]�A�	)e�����1����A��2� ��5�ؠ7@��Eƛ&���λܑb��o4A ]Q�q^��i-���ف���kM��0
�ʄh�҃"�K6�$n� g_-BQ�=H�#݇F�Jqt���ͺY�hڲ!*�r�l�:k0�9s�՟$����a���K\�i�ne}N�c�P���C����l�����/66��8u���8xqГ�ԥe#�N�:��c����)��΋�U��KX딍{}�w9Ӻ>�2�P�o:��V\��2&Se˔�\�Qy�{l�{x��ɛ�vQ��sn5��#x���*����U���e'�S6��f
�-빐Z��Z�jPA\kV.畀v�R��Q�oW�X�O�z�si��xp���!{S+��`�%��V!#�7i7۱" $Q�Cqi�����2p��dT͂ZmN-����	ɵ7����5��	�c���k͘���3�:Q�9՜q��p+"څa�H����ˣ��:����*WU��m'�B.�R��S��՚�z9%��^�[����b�����PwA�ٹ[�#C�ibY��ө�1'��ZzU��׻sg9��Dt&�s#U����71�� �6�d��m�"�T¬U��Fu*oe-���X�M��i"��LR�pP=hg^�{G�F,���%��r�E�*n��?q7S��^ />������]IN�&w����1��V�u����SC��2;�xʾtv���Rɶ�Cf	�o{,&��Afk�,3�J�2:�h��ˍ}/���l4SlB:-��Y����^f{GZ��cW:�`q�W��^(�GLssusx7:���Oan*H���)�A.\97qK��gvM:p�;���w�� �w����;���.GH�u˸��&iwwi�s�.�فg]������wN���N�N;s�,K��у�놺I',t�8w]�gR��Q9˺��w�:�p���܎9v���i�wGgq�뻳v�Ύ���E���wq܎r�pDwu��wu�.���=��v�˻�;���r���w:~:���r��yv��:۷w!�=��������λ�������ww\r����C���I�iΙw;�wkӄ����y�E����qu��u��Ǯ�����\1{�y�ܽs�n��ry�O9;��r���w{��<���/{��z���n�x�s2B��ۂ�7/wrv�r�������������w���wk��qv���{7����w��޺���v�����w��פ���&��^r{���sy�ǽ��{{��xM9�%�r���;ݷ�{~������yח��:^x�y���x�oqs��`���%�����b%ywz��!��K��ݼݝy���<���R��
Ns������<��o:G�ּܼgu�^oE9;���o=�{߯�ǿ_/;��w��!��j+��Xȋv;9��W�49so�����Ic���<����2\����Vj��LVJ2����+d}��Zܧ�'�+�����^�2/�B������[��8�{e�6
c��d[�	���z\>�g����W�q�~��a�>����\��=�o5CFnz���~W:���1�Q ﶱ�#d���Gd�Df�WL댴&�ڝI9����^�35�ڬ��������?W�(�ff��O�ѻ ɺ�L_G/�#���:3�(���BqA�混E�*�UJ�#L>��_�o�e�/��n��7��{�B��\].����}���7��=�l}��=����A���g��T���U��%>�=[�C3�H��MCGn��@8�}�#��hY	��)��1����z&������U01
Vu$l��-�|�2�k�p��Ը��;��gӒ]�:G�P���+)$�w��6���\GC�Qb�1
ǕD_/S��ݶs�|����
����`%8������WG�}�sno�>�_p&� ���b@�����7��_��E�9�y����6L���Oز}����SxO�A�{`6�A������XT��>9�vU�`�;��
Z2��������ز�~n3�k��6"���}�.+7�j�M@t8V�sǹ����Ng�q�	����+��Ur.4�3hڕu��,�/;�3ܡ�㚀aCΉ�����z�D��n��J��W��W[/D�p������%��b�������u�?|ל���z\��@�al�l|H�
h�"w�`���
��1��Ƹ���ڱ���+�=|.Q�Vm�"L�p�sNU{�3~j�������_c��tR�Է���W���4���;^֯NER��u�n�_@���O�N�,S�֌�8�џs���>V�	^;�~t�TG:�(������]as������SOC�WIG}ʄ��m��CT�xؠ�ۛQa�����>G���{����]��׫^�c���W�R�T��6C��q��P��Z1r�]w��z��V�m~���e%y��W�=fy�_
%�+���5-�=8�=���������ʓ1VnaMxGf����M׻��Ν�QB stb��b9Ʊ���3e�8�<�p��y�%���3} 7�����2�]������j�>���~��mV���C��# �\l���a�� v�iC��R�Ú�y�F��3ޘ��s�^u�y�������7�H��"|��aOx�/�9%_�"!�FG��]�"�2�B.ߪoL�@��n���ձ�c�+�K�w��/���r(wNIu��vb��0�������!�*i#k>a+�1�y2�`�ԙB�P=%"L8�9��b�0� ^3�7�7����>���}��:�ᮡNS�]�V����t֬wV�NB�J�x����c On�NsPՙ7Xm�wR�-��w�pژgVU�c�ۻ�"
��zTB+��V��C�$�gP�]
��,�#����sl�u(P��p�D�+�v1�0-3����:�sZz�^���9��9+��=�Xn��`pkT��/��A����@�v����r�2��
so��{�^�Ї����,�������Ü�i��6ٍ���~q�}�N����:��S^�Bz���L=��e�B��Ox��mu_'��8�"C=4$����Q�nR�Y��͝��0W��<�V�¯�i�cSF�:P�5�0XI ��(`�B��U�������JAx>Z�Ǵ�]6�ϩe�X
��1'J��Ы-���r���24���:���i�a��ټ���Oёp�9q�+�tm���x�������NR9�Dp}�] g���z�C2O�>U�eM_Pf�2�Rp8s������d���Z��cɻ=Wど��?@�̟Q��>{0}����H��p����@qb�T(����A;���a��f#W��@ga�&�]�`�w_����0�TB�UF(-�������,"&��0��В*-w�����qn^�S(�ض<�5Պ%�䎇q�"E���g��1�S�R﷈x�Mx�fζmTZ��c��І�_R�^��t`G���g�]�A δ�S:�3�Ê�0���Z7^��:�];��sI��k'G�*�Lj��"��(8�J���'kީ54���PKqDjs���PH�b7溦)h��c���-?�D��N#���!F���9��\t[%���q����o�l�E��a�?W����}eǇT�T������X��{�������w_��a���ENe^��} [ϽwQ�ܨ>+W��)��1y�� ��z>�A蝺�s�\mCy���7>�.=z�=��z��u҅8�R4��dbB���Wq��q�{<����7�xf.20���Ȥ��6+:�B3��i���p��uQ�>��=�V�7�9��m�@pZt/D���cN����5�@C��;w1J�0��Zx#N�]Ք3�^��c�����9��j�y�l�ơrj�|,�/��s*Y���M1�2�> 9^�2��.��G�^�x!f�ݕ�,b�-�>�t�c�B~ژ���D@4˥I���xp�cyͩ�~��!@P��\�J���t)o��E�'}&��8�F'*�Ԥ�XdQ�՞�V��ͥ�����r����~�\tT�;�j�yJ�~!E�%�1'N>�C� Ue�����5]SpJ����b<kWj	g�E#-3&5��آ1Z��᛼��0�:�cN����C؃�t�WC�gGy�CDu�\��ĺ�Y��d������G><����6x�f-�@����؟7�!_|�\�-V�^t��xvl�'4h�{��{sބծ�B�Xӄ�D�'�?��`����m\k��Q��[�@��V��@�_Y�=Yf���Wo��l�ҟ@���t_ۓ�C�*#x��_xt�,O#@I�.����ٽY>}
�6/h�T���:{�����qt��	UtZ�TB��T�D�5��h��k����Ei�_a�E]��'yGWs2S�z�@Yԑ�?RBBGzқ����Q�	��&X*>|їJ�^)}�;]X���]K�R�n}<�+��@tls�����aG����/�^���٦����¢��z�ě��z ���P����\�/}�cb��W]�P9����H�c�p��sP�{��:��{�Ȱ�a�� T'���r⾟O������l�ǃ��#���8�kt�r�т��f���Or�y��o� _�M��?�l	fsa�'����4H����~��k牻(��ûS^�,�NQ���X~��[9�>��`.�x�U�F�	��9�	��Tys/�ŕV���}��ǻ� o�a��B>p/��6q7W5n0�Ñ�9���5^U���k^���3�<�I�C3�y�A�j�pW���S�1�'���w���7�d�Cs�.p�d�+��z-^�@������'��ӗsȺ֕��-T}!��4�Η���#k�E�Ş��̭c{�wn5���;�G�m��R\5�k2<��:U%�د�?}w��m����\���8P�C:�1�Yl��f�X5иq���8��;��gӒ\|T���"k3ެ~�.�������-�B�m!
>�1����n�>
f�O��-X��A{v%��<j#����`8�9m���xpp]��H��(.�=Ցh��t`E�I�m�G�e�k��MPydt�V�����;�>4:ګ�4�����>
�Wκ-m�"�q�a��RʸX�������V�8�/;�+�͊����jL�O�Ф�T�$u����ӱ2A��� ��L2+��|\}��_����ff���v0yW�=	�m�gt�v�j�w?x;���6p����B�H@� k�<���I��:���tuk�>��t�U�<��x] �u�ga��O��*��Kί,����v[]M{S�n�h��{�{�C�,X�G������l�;�t'���!`���8��sjp��	��^�|`�a�]��՛j��f���M�hzL��>� L!1�޸���ݐ����X��Z1|�1���ۓr,7uٝ"�l�_G��������挊����ч��l����+ú���UY��oa�QU���f\��ErD����"�"�T�B�5TKd��V'�S0�;��5��+�gL{�ӭ9hÍ��7 \x
���o�Y�.�8�El��Qo {�"Ď��j����X�������^�H�	Ի�2���I��_H�f_}��l��,|!��t��$rl^�Y�1W�����lUͩ�X�����h;S�s�pfe}|~)_ov,ϙ����Ḅ%��a�s��X��~����>��{����8�o�4Sg�}髍�v]�bg��N@O뽱݂�o#x�ϣ�[,3o�*��� 6��}뜒���^�aV�z<�Ӟ��He�>#X�� E ��_�_%�~:9Ͳ�=v-˥�^������Fj�7����y��N�N����r�#.��b�mDpΐ(�\4XS4��v1��Eo���C}�n��^{<�y�-�����h�����0�_�uk�఍�C�=��ˑ��_��Y���g{	>��k~�z�e$p�=7� ��0<0���(3�]@�<�T8��f1º�w�l�]xo��[��/�9�LU��y
C�'����W��'��!�0�wO�0�\V,����ͧ��f�3�q���gO
_��;�+�� ��6k9҅mm�
��1�;�����c�����Ɋ7g��o�g�#H�$]9�V
Yk��ϊ��1'J��S����v/�}�}f��2�'i�Y_�Y��{��̓���23�Zڽ}n�L��b��W%9{���<�GI�{zʩF�M ��6G
ymJ�ё&:*�]�bt@V�3#Xm�ϸr���p�ӻ�֝���Ƕ�9���)���̚�{b�4�.4��-�{���V���~ ~��'p������Bq�C=zGG�ܬc���������#���#��ˏkF������j�E_n��zp�ށ@���**A�*�h���P:,&�,���WU�N.�ӹ{{�e_t�8��9�G�/�G����R�F����gD�fsO��e�����*��S�>3Weyv�������#��J�똿�	�e��C�Q�4L�� h{��kDWE_�V����q�q��N�omD�hz�$��BdP�?�A���u�ק$�X�G���8�W�N4m����+�s�9�RӀU�x�f�6=��5��l'�sU�nO����9%��˽�"�㕈^�?{~ూv�/H�8U���Wo��=��|V�!��^�����MX��q]�ćs�s]�����	��몒����z+¥E}$O�����m�GE�҅8��AÏ��y��T��|�}�zsv���YS[c1un�EY��g ����@��Cbܟ��PY׍�;���ݟ���4(�n�u�3H��@p�ӱ����cN��60���C񯤶�A��>%Y��z3;*8�*?��{@{ƅ[%g��w�.��-�u�hybE����"�Ui�셨N�pQ9t�5��u5wq~����s�s�㽈?X��Y�ڻ�R��r��^�dj̭�/{�S/��e'U��k���|�:�s�:Et+�U ���N~�A���N��A�fz��L�Fj/��q�/ߣ��|i�-~/N��א>kMm�ܑ{��=a�)��.�,GX�)_����4ˁ���E�GM·�sjU�H� m�OJ^8~��x��ʿv�1#F��X�
�(V�X��V���I�m��'J5['�(���N��E_��e�y�O3�i�W �}~s ��(���F>j��<��f��69�*��I��v�:�����t]c8#���ґ���}�q�F�&��� �=;5�E�`Kw��p�����_�6u�{X�������jR9GW��j��7��=ﺄ#�H2��4$Ɨ�Lo�o����G�x)�)ӽ9���	�s�}�s���Ҫ谷��N>��DF}AH24KDQ���mFd��/���/���z���Δ�t)��);5)���p�ݔ���ɪ3��$q������}yO�0,�*i�#�
���^�+�{o�e�[ ��vLXG���1�ۈ5/�ؚ�������������^���.='!�c�s�uGo��U��(
�~�������i��qJ�܈�U�� �.�xR�.��\Ev\x�{�j z�(�Ŧ����M|�QෝY���떋}��`0���S���o+�ek;.�B
X�P�g]��O�+W�f�u��H���$� &���q��(8w�X����$��v��O"^�j�A����f��W�j��2������7�U�a�w�����f���Cӓ�[�(��"+vrC���y�j%���	fpl0������4tG�6~򣒧`�����b9G�Ot���Z�@�S���g)�lt����F�����#���������ae�z*��k �/�C�Ϻ�/�Pd_9�l�M����j�f}3�>���Af��$TMn�WӝIU����Y�b9ї�3�+:�6M2��Vk�p�&��FN�t�u�7�lL��v��^�����$���C�����#n��B��Q��L�CU�l�i�؎�h���8�����y���7;������#~=��$��%����:��VE���Ţ�Q��z���}��Λ3�E;}0̮S��]fF�� M����Ѐ碄�8��P��ʸ������4;�gޗ2W{y���3V�z:M��e����r6G}�$�<��h�����#o �}�U=#�Y�=W�Sg��MY�s�wu�6LF�F������A�F�6p�Ç8x��}����<�ǝ���'Ǿ�҄�df}��؎P���{+�]BB�N	���!Y.�ؖB2��ut�Թ����ŉ�DoWi�3dT^0+^nR;Z�Q��%�=B|{�X�^��{K7Mm4�QN:%*���;�{h+߯���.(PT��^.0�Čr����^9��;w5�ɷW8��F�:�l�(��Rv�p��f��F�#+z̑t��k&;����*´�0�y��vN\K����dx�_i �315�����}����+�A�'W�ƇN��)��
��V�P�uiC��i�R�^wĳ ���� ��(*�5�GrIkR�]ų��������[��Ki���c�-�^���k�Fv�՗rB�%�u����ҁO2�����;Rw�u��P�v�J��Đ�R���[�r�N �4�GV�в�8�i�h��`�����D��k9�����Ѝ!i�c��}Y�ԙK�u-�L��4s�V���3V+�;q^���Q#I�Sz)�o"��n��,!�����/��i�%�c�ZpɖfI9p�}���ײ���!��fp���9jt�!�u#n���̽�x���"Xѯ�Ǆ��V3e��b�O�a��P*�+`���y��9r�B��1�c�YiS�P�J��>��{��%͚������(m7ej�Y�lLk(T�u�;��Izb+vԛ��cE\��n��̝ٲ��P���	�P���@�v[3y; ��)t��h�Ruh�RC3�����������u
�YC>c*)Vs P0�$`51<a�����~������AУ:�<�zg�6;�c5MW�^��"2�N�����{M7�/)s[��ҟ	5*��w��Nr�|�K�ui%Y�*��T�M�5%�Otb���*�l�d�Aj��l+��HU�)�+��
��y�4���u�r��%@�b�Ol��L���3�0�����0ĜA*79�;n�C�1�B��d�V��f�N��#����C3C{��/e���SS�h[�;t���3�Zjgl�Ẋ��]�-��٨&=��˜���-wz����6�3�~�;ڦ��yV9��]��U�&^uZ:��;O/��2J�����?_��f4���r�4(�r�So�G3��f��VuZ���7����o��#;G���|�4.�-�w�V�g�KEX��粉]�ie�\#'${�kboc�r.N��BwM�&K͡����	�ܩ��r�Є��\��-N��\��|5MA�V`YƎ�ΝG��r�v�p� ���̺�K��{G��X�}q�=
���z9�}o:���3Z֪�Dr����.ܧy����qtTw'ϩR�+i����@O�2ە.#��^2̥�Q��꾦��R�!�\';[W�:[��>R�g��'u9��ru�d��yƧ�����$�?,��wB�^���|��7��}l��}��!Rg<�v�EY�j���D*-۸@���e���?|@j����F�����wc��������{��{�2�����ׯ�.�&��=�Ļ�q�צ�Δ�����q)��7�9t9\{�Ow\�+��]��FB����q�΃��r�qݷ&^���.��L��(�vn�ܸ���"c����%z\<���z�{�C��!{s�Ι {���޽�=����9����t�u���뛎q�wn�N�7w�������+���q�޽@�ח�qr;r�R\ws��6�1.��3����wvwu����ܒ��H!6�]ѓ���^�޹$���02ۤ���Q�]��y�.��o;�ΠN�xK�]��w8�:�bS�S��qR�+�u��a�t@�\����wnr��w$$3��i)����w+��;���:�\����P.�1Ҹ����K��..�r�"D��M
	"���9fW���y�j��M����'ICz  �WY�d�����u��e����DU�[�Y��W�gBUƑ��	�����uNYy�����>���'R�*�s'�&8�o�rY�s�n��3��s�W�خo��G|��X�����'^��[9��1@��	q�R@q�n�J;~�bz���ϛ��U�x5�[4��yG�=.���Y}�����`����9QBj_�ϫhl7��#�y{�U�FE�mW���Rs+�f^t�3�$=D��Xe��hQ2��'��l�}]^�¼;��d�z�ϔM5wjwb*��K����a�^�,�5F+���Xefвdx)���pћ��5^�}�7�ˏLy�gm/��]7��L�X�����l�ס���\�G	�H��Z��'��m5>SJ�9������w�,j�ټ�ޖ�����*�װmOx�,z�$���\7�7�l3�}�mޞ	q��=���]�˵�r�n�ޙb����/��S��7�02������읙��Q��9t�>�/X�F[1�1�o�~�S��2᳁L�(϶�v��k�uK�z��{��=lS��)���,����h؁����w��)�o���}�hO��¦��f�^�v������W������d���\qm*���FLA��.�ܭ���_n�1�F]IF]��
�"ݘ��$�����-+�;5�������uyN	s�o���t���\�v����2-Y&]B��8�u�GW�Cu���C��{�R��� �2vW�u���*7�U|g��l	撟+��t�a���%�'�RPg����ž�sU��Q�}Շsh�k�ǫ�
��+��#,�Yβ/Фt=�#t.���'��9!��0�>�eK}�z��G�b�6��Yb�}�n�ة�yM��(Vۘ	1���T^��m�nv�ٻ�=�~��bd8t����K,b©x�����4�I��[B9`���B�M���U9y�*��<�AtD<����2�xWP���+�������r�����3�����x�]���v�mxWC��|���'��C=����Vч�������]�z�T�L;���������:�Ә��	]GE��<��R�$�h:�M��3�{+����g�=7Wl5'���ێ!ge()�a)���:�Q��h��}# �@i�d0�U}�|�zpw��8�%�3vXޏy+�M�9f�F��D�zq�V�	i�bS0���Ma�W�Ȉg���G*Ǯ��S��V�rq#�;��_|�~�S���^,3����X���>��~�~?h�چV��������t}v��U�;mJI�$��
�/��ɂ�I۵jĬ<���~�>�V�^��W��ըC�p��]\n��2��f3�T˗�n��+c�w�I�}��YީFE]w�v�3���t����}�5�p:�v������leS��G�$�$� ��[���-�w�������DT�U��s��T�G�:�-�/��:��^�=����k�����=�^��`_����5�3���Z�b��}e vE��wQ��	q����{y}O�#���E��>+��L�Y�ـ��*�r��i�>�}�_p�7��mϱm�Q�1��pz���h>�h�3�ʜ%�c0O��64x|L�@���f˖�+����ǲ3v�W�
�9��P�T�~��h�ơrj�=7�Y̩f��FΜDVx�my��v��w@��bg������hP��rhb�d�}t�o�Sq�z�:ԫ*z�<]�ӱ��o<k�s&TpF#a�BTu�PP���,T�|�d���3с9P�NLO��+*�vl�D�f�����"�2�A�������O	���h��h�~��qe	:�>#T��f��v�vܼ��}������Q�iXbz~�OUx����T���}/8�B���*��o>�����8��Q��z+�*#lt��"X�����F�Ɨ�}Վ'�8M�
�q4�7�Vu"C4��ajƚO�_�����;��-�n��͔�yK[)<$�����$�w����E����ݍ-�+7d�#��E:�3���R����U�jâ�J�4+.������6۲�+݌�W+m�n�D0eU9#)�$� A)�}�{G$a�w��J?�:�Y��ns�}�u�x�U]��TB����
�R" ��~x/*T���OV2LN���t�S�v�F�Φ�`���@��	�	M�Ah����
�SCs"<:'kެ=ޅ}��#������ �N#�[>�߂V!{k��-�m�P��at�ґ�Ȋ���!w{��0��Lܞ���,J�����_i��W��~��9��i��5�;UP��wl��ӫ����S��b�|��&��w�8�(=,WK��W��:X�^����̞����������j�obs=qm�p�a���(m����6<o��O����9?W�\*��ݴ���>3ʳy���V���9S���3/g�]>�ȫ2��~�;&C#�o��޹[�&��[]3����>���p7�v��|�F�Q�#��l����ϩ�}���Oiذ<r'�n��+.������|�L�F��M3�=X���I�,�{�5�C+5иvV�"|����)�Wot]e�B淧n��,\s�J�BY FF�~S�d��ݶ}�S���΅��{?��ڱ�k<�"O*��`P�֌!0�2�R&�9R}	[�]rk�/]��.�e���\^5|�0��H�
�z�S�c����^��I�����<J�����;y>��̢�;P�7�G,�ح�C��H�PAs�&��	 �E:�P�(�?��﨟� $� $@$ � ��k���^:��=_���Б�w����� [O�P�m����VE��y:1�2�q0��b�8fO^�%���[�:	����3Wk��P�>��z(IC��0����w���R/(φ�cg�{u�'�^�g�4f���Rl'=���#��F��>��#�@=�&����[��ˡ�X��ժ$�ghR<��B�\�y�U6z<ԫ4�W���#�6p���*��p>���e{��M�ކ`O����7�t�;s�����?����]�;�~.��an��g���;�מ��y����,<$�y������X��V�5W�$/U���.��j��WoJP�F��D�t��=<Q�MK�X+hl7���q���J;�+��Ei�+�ݎ��W�]F$x��lq�2�hQ,@1CDd�HR�y�uz7
���5�Grm�+cG��LF��;�Q�=�n�E�Tc#�l�M�^�D���T��OT0�<�������1�.�+��|7f�J`�zs��Ok�-�[���w��?A�{�����0<�^�֏�h����K諡kwr��2Fu����c�(̙�6rI����=6�U�2�c�K9�񗘋Ѡ��v�'�E�j\�iuF��>�H�лX�R�.���8�OU4w��"�}�6�1�d�-c���`y�Iه�C��[��u/f}�߯~/�����᪵��mV�@"�$�� �{>7��w�Cx\��o�>��~�� ��ȿ��v�xD�6����F+�HGw�{�[�N��x��nc�H������Ʋ��\�z���,CӜ��x��b#�^�͢]��~2~�������E��Q΢�dP�Hr�#&f�>�¾�S��%�g��{=�V۟`�;םX�q�ְ�	��W��<�u�-�zOӱh�����;w*vP�c:���7##��!�o�\K[��6�+c�2&:E3�>V	U��'�fh�a��P��<9g.8.�]��G��������:EB��W1���}7��z;�H觼hj�:OA�@����8査�=��k�[�b�n1V\��ا6ʕt)b��*|f1ܰ�N�&�Я��3�n���$A��*��y[,�d�Bp�;~S��o��Yc U/�N���g��`d�����d��sk��dծז����"1��E	
K�@V/�tm�+�O�p}/�u��IVqZ��JiO����?��"/���h�%R� ��~�,l�W��W�m{��}Sޏt�`��*}{r��k ܥ��+̮�D�l�y����+{{��!ye�SR��O����)q���M��/zd"@��F�A� ZV�ζ�O����^�1��js~��Y�d�8[
t�ei��c�yW�68�����}_Z�%��jՍkh�5m~�?��G>K�����;W��"��WQ�k�y �"I��({`E8Ox��F��-	�E�G�c����w�1�0W�@�SHń�#�R�1�NB�.
>h�)��>�����v��s��� ��F�����i��Tڐ�W�*���r��XfVO 篂���sЯ��b!��HK��:�Ѽ7�+��l����A�O��j���9�W7������5{�CU9%�M��	p$`)�_NeZ8*��}����X|�>8�X�}��ZӃ�r߯��lwS~T����z�7'�T~��|pL����M��~���1�w�H����}�kX�����1zGBa�ض@�)����t�*��9$0�"�dR�R��1���!�������ޝ��O��UY\�(.Zv3���zw�Y�>&h�f���I����3aW9�6�i�p�U��USe��h��VV�x��"3&Y�\3=b�Z�o�ݚ���������ˀў(B�!B��9;�m��KE�7
�ԠeBߏ��&���L�i٣�~T@k�G[���o�u��i%�-�}E�v��#�4S��b��g`��3��e��٘o����f����Jeq��:p�e�u�:�m��3&җkF�
[��Ӹ'$ޛP�g�1�yֆ��ȶ��C��A�		H		 I$�� ;��8K�^u�BH,o���z0K���8[�-yS$WM�.~S��S�b0-��_A�og�Y�ܺ<Ӯ���I�;B�� =KD��S�<K�|�Q������7��$�U��{S�]Co��oӼ]g��w�3�����������_u�q���B��:�����yl]��:��~��{k ?�u=8��r���z7��T��N@;@uG�e	�_���Ն8�V�tukf���0��9�%;p��s�}�~�:�谷��� ^
DFe�J�q�)���=}z5�Nx��i��Y���U�;hDm}��=���K����F���9
+*=�v�Am�%�uٛa���(@b=�dӬG+g�[�V!W��G�llHc}쬹��Gޫ�3seߺ78���F>~������<%�E<�.�?~.���{>�u����0-Kh��!���[B�k]@�5z����3q�3����=2��}>��]���ZK�fwf�#E���{�z�#�m1߫�Xmm��g"����,���s��O��<=��}����~������S�n��3�M�}���z�r��ڳ[��+y�ݫ��[�uH<*ؾ�2��|�C׵���r�i�@�}Áen�4G�mc/z���C�����bi�<��%lS���P
�����V���>��ؘ�iUx�0�dM�	u�m�ɵ��֭&�m�����;��	���#@��y��ն�7��o��~Q�R�8_?:�pS���}�xo���v���Y�z˨���{�Fc,���*��hgm,	��9�Cf>���<����;��nl��r���ދ�/�^��ǎ�A���3��������I ��-�)�ek�PߡvB���P�w���P��}9%��?!�FAnb7յ��T@u��"��n�6��#:l��w{�L!����r��gP�#�z�K[��ԇ���x?-��^�Z�G�}_��졼���dH�F/�#�X���t6�`5WWN���O�*������k��~^�觬Ģ�r�7>���f�M�t6��9�6ωJh���O���6Gy!��In��(��F��Lqt❋E`�B�X��#3᪛=������}.�={8LF�@�(9�\�v�������C�n�{�O��)����N��.��X������A����A_�_��L��۪���1z`C`�b\/|n�ƣWIg��	���X!��~?{��ީ�ˇu��g��*�>F���7��i�V�8e�rmt�}[_�w�T�o)�2�y½�L4+޷<k����k��Z��q��2;Ιy1�'d-�lE+6��3�g1ِd����P]H�ܙ�j5��M�_1w�"-K���,�uo;��������Zѵ�m��E��kQj�լ[TUT[wϿ���E;�����'6����P��#8� t����K�^|E��ҡ�L{���ovV�6o���)��[1c��0�)�$Pz'�8�{"Ib�=5-��fׯ����q��]��ֺ����qcU$b�u�b9�1q�l��XeX�L��V���'�]�Յ��U������/�+�Y�7�CK`�^�!ń�HE��`��ס���^n�zTFټ��w����%��
��Г������[7�czPgaia��m�����
�5���9$�A_鳒U��CF`2���Mq��a�����e�zs��/}Y��a^�zs1���n����[��z�:�$�'�f���\��ˣ-����0��*�Q�n�C*g+V[˪���������/�3H�m�ǀS���Ӑ=�����} P�>���"�ex"ryq����抯O���ޓR���G^L���W�2�#!�G�t�f�|�,�X�`�a����"q�-�
�]�$"���c�.���~�B~*�l"(D+�y��}��\���Фj�;5�d�bu��Sk`͖0l���͝8p�Ç�
�9�*Z!��Na����,nL�fP�7�-�y�':����٣��A��]�Vm�Ź��V�<]+W�OUB�uÃO<�9WR�]�%K-�;�Q�
�+�I[MX�])فJ�3&�X�`m��+��Ԭ��Zx��Xv6^l����]���h}�*g��ݴ��H+2�Z;OIZ��E�� �3G��f� «�'�vT;]k3a�"��	�2��u5ɗ��AR��r�	��Ov�l�ˤQ����#	Ž&f������$9�ۡ\�K�8@y`�O-���g=#z�/��X˹B���m����	���ؓ1��xh�Nմ,����*���d/�W�����U)�HT���I��y����^L�y����\0޼::�������Y����'R`���d�wk�����N���%k�2��wٴFꚟ��L����w9� 8f��*i�s���.QIn�I*޵��T�d�j�)�C�ԼL��������3��K��D۴���W������
��B�[����6���`�LmH��d�Z�"d?��M�u�'A=W�r�"�כ���U$�T���ػ/K��Xmv�8�t@S����00������� �Z�h�ո�ʾ�#iÓ,�S�̽n)���-�r�仪�&u�ݗOb�þf�.\m�Qd.��';zf���i/�JΓoPĚ�Ȁ�U��hW��%aU��뙭�����\}�v�[P����q��hʜ�d~y�K:��}��#r���NT�z�MwryW*�ݦ7)=���ͭ���I��Y��GO�J��+&� ��9%c��b�1�`��p��L�����!�h#�f�R�)[�ɢ�qq��������5fV<ɰ�D���j;��_�6Mn�Ǔ�kʦ���agk�Sz���/�����������0���"�a��Cpfl4k��ЃmG�0�9,���;U(yHn�7K�׆�5�'ܸ �Oi�d�'&�ս��qsY%�r��.��O�a��P�}� �fR�����&���pz�Y�lR�㧗4��'LfN]�imaحVM�FO��sܱ$��ؤcm}�k���͚��X)�̹�%NI����N��ל��8�b��{�ֈ/�b�(�#�V�yZ�M�܎��ԙ��w��V�tfL��'����k��;���*���7#yoEqqh�$]P�h�4������/4��U죮dx�zDwX/�k�� ����{8:wۺ6���:2r����Z����Y�Rd'F�빗�%�W>�n*����t6I��\��Z�j
T[o�=��A�F��Yt�o
���
SE�u:ɓC�Г��V����W*(M/-�|��s'!��1�6���E�VS� ��Y<�q�˩F	-��I��<!1��f*E���²��>&��~&���Ir�;��e������!
9�QQ4�; l��Ý�ɗ85r�;�Ɛő���.nh��F`S�:�Q��1��n�S���y�z��J���wR볎�.N��$� ���H�ܗC;r;�LAS�S\�B%3&�;Dk�t\��R��˱n댢d���A�q�]���α�ffW:��;�i�h�wv+��]�r��u&�]��t.K�DĹ�)���F��N�v0��ౌd���Rsn����˒���WfC���'v�wu�9�4	.N�D�'wg7�9�+���
4�w(h$ɇ]�:tgwGJ�swu�&�ܒd����߾��+���IPӭ�.�6�Y�rmn�O�9�⳽�+���J� ���T£u��ۼ88It�6�y#]vk���گ�Q���j5�F֤�$� H��$� W��wy�&���4��!�WM���X��y[�w�*|f/�yM��(Vۘs�� �z[y�����b���z ��!G#`WM�yK,b©x�IҀ��t*m{�첆;���RO+�l�W�Å�(0v:���C�
\+��Ѿ�B�O�v����VU�y�m�go�w���_��G#�"/���G�%��D����A�*�h���[dLX�p2��^�ǽ��N�#5�ڨ&!�_�51�	]GE�H�6�*�
'� މp:�ͪ��I�vO�Q�8nrL-<�uDw��@�g�wLF�A*�A�^##�Mɢw�|�(�\W��q��g���xO�hI�}�r��u�	�N it���SJ� ��NC+"d�!>�Ǔ��y�c�����T�� ��Sg*�<r7KӞ-�P�^���A���#��#��/��R�}�ۏ�aO���S�]����T�9�h૟E�z��o��
�g՚�zi�k�[hD�M�.�ծD[��OӼ�Ƌ޼�u�D|�~��R>�iq�`����-�>�
�K�AX��-�e�w�Iۈ��8m����A��2v�1�Q�IA/L�C5��:�>�;P�3��c��B��HMZ���$�
z�l0�w�VK͑�S
c��'G���X{� 0�VNo�/#F[l��m�ځO�t��>A$�I�j�V��kd�m)Uo����m9�Z�(�d��ʃ�o�ż��n��ϗU��U����A�aNC�(Q.��P����Uo���r��T>���B\.Fi����8�-;�N����6���R�ه>_�M����W����p�A��k5�Ǆ
�j�l���h�x�d,7}8���3��{�ɼ�k��c�,a�H��#�&\�x�|�
v��ѿ)�\]t�~�p�=�ɡ5����Cᴽ�W{;�b��}eE�H�27s诧�����e�Y�l�v'}&׊��5[�s��9ڽ��T&����L��l��	���<'c�Vբ��U�O��\r�7�<����os	��j���-��6�g�9�M�O�N@U���C����:��ޛ�K�w��)0)[��S���u=8��(�9]�~[���#WV%L����������ڟu�9���\P�ax橸D(�s�=gps���������[�H؃
��
"���y/c;9���
�d%�s �>G�V�G�v�F�����?R Gf��������ML��D���ȟ!!+�J�U�7qՐ�����.!�݃"��L���wߚDv#W�[���/�U0�r
�G��$n�!+"&���������̭5��d�����k\qWf��ɖ���D��:Pjc�hЬ׏�E������eӤ]Xt1�\�u������/�}~��������-���m���h��6�V�UE��$�)"J@�fv��o�ЧkI�GGX&;�&~Dy�N���io�+������[��s������|�ʑW�{��n�V�~���.Ǧ��bTTW�zT�l��k�����.�����9���w�Bkw��S��t�Pcy�$ٶ}��1Zj�10��}>�Y^��`�|0�[wYc��{�����_��'q�j�`�{[Co��k���2�u&G�<����j|�n�j����pS�ϧ��b����o1.3~�L@-�ճ��V��O�la�2��w޻f�-[g���tb������f��P����w�c�XdX档�7W)�q�����e�y_�����w~,Af�4=#�摈�ї�ґ�2�E��e$�}�v�d^��ގ=��܆E?���?a�ܮ�>����!LFEKu�+k�;��2E��m&��}>ۨ�ޒī�k��nf�����c㾁�a)�lO�j�	��'�	q�[\#��bwIhM���/�:���Q~}F(b�&��3���$m�4:ګ�4�l ���9�P�h�l{��t��b�(�gC�Ӽ��:��O��c4����~�L����1^��*.����=�f�Z�5�u�޶�b��s.*�J�(�-��bZ'��os���7a|"�=mk;y��v�iB%lR�i���:�U����D�$K�mjf��m�ڍ�j���*-k�QM���zxrj�)#��rj�W�U�Tћ��%3�\a#W�h���}�
؉�n��/qڻ��,K��T�I-�b�x �Bᔪ��KgcOW�6��}.�7����M���r��벯<�1s�$0[4$Ɩ��I��V1�.��<;ϫ�����;��Zj�O�ٟ{e� �x�X���|��%H������/��k�����y����d���~�tM��u�>c��ս�qc��8	8��p�4YPd�+~�����c��Ҡ���-+q�E��ثU���\�(�^�8��2�D��1 h���Q]û'��������`�����^�C½�_Nz;��U$b�u�b9�1���5�U��d��f\4$�s��/}׃�ׂ}NNC�y_;ݚ�^-�9�X��!ڭ�~��1[f&�0g������q���AE��2���/�}'�7`~��V��_�҃;��~�P��υ�^	'���;���ݏ`�;����
���#(`�Dz�Mq��>������!鏣�<u{���Ɔ�Y� N�8���c����&4VⓀ���m9�VTg�GNy��5a���CM�l��-�!1�I���q�I��ȳ�ѱ���\��J�z��듌 ��Bt���c�6oB�6�w[攺�2��칝4����_^�~������lmE���m���E�m�E��V(��$��r��Z��ꁋޖ����"y��nŇޯGQ�/�>�}4,R��S�
���~��J�S��U<�z�=h穭f{��l1�=�|�i��6�c�v���h@�zO�NŢ��ڂ��N�$�������u�΄'�uD!;ʦ(.�n�&�uf�|�,�X���3��H�ye8���#�]��}�ޥA��uӠ�7�"����t٬�!��#�������:��n�<]C�Lb�z8��W��:�AȔ|hIB;��M���X��V�]�T��XǔѤ�B��_dQ�9Cl�=�ys+�z��q�`����w ��C�G�WM�yK.~�Y�T��ĝ��1�h��R/�k�bۛ��n���{`8@�tYt�~@�u@;!K�
�~�cW�:A��h����`�N���#��;����xWE��U"�?D6}���p~��a���܌J`b�E�&�,��~9�S^J�:4.��mU*L��H>�uȫ�p/'��Ճ�*��54��u\^wTGyz����J�;�)�Z'!_H�(���n�S���Q�K�/&�z�d��<}}[��>`g$�3�f#�f0.���oD
�V��Y	�Rj`W��n�|h`�f�Q%�[�.ވ�evE7�U��;\��ަݨg�w�N���F-XA���_8�ɦdu�[ w��#/ji�|�@?%I	��	lkh��X��f�h�~sy"��{_��`�HK�Ri�@�'r�{���]!p<�BJ�:�����u�h��{��Ma�V��D����Kfh����/���G|�,#޽wSq�n��0��w��b�����,zs
���ר�SpgD���~�"T�p���r�X'chX�����-�o��S���Eڟi��������Z�ݮ �ޯ@v�G�TW�_��׃����4��?���*��{\t�J�װ���GE��N7��?;�S�_׻���x�dz��F⺖H�Ҫ���O��hG���n�ʮbtu!p����+9WE��S���2��@qbZv3���cN��+d���(Qo�Qy���`P#�jK`�`��ᜯ��T�j�E�5�V�+�����&'�q��K�o��|}�,����#��ˀ��돷�B{�ŵ���)�\���E��v���x�Y��-�ۘ�U�$F�p�1�	�.:�8V<�Ŭ���"�����eu���=��*��I`>���r�X}JOE�Eg�A�'� �ة�;u�h���cT%�&r�_�o��l�׊tA^�HX[�Lqاfr�|��\=PٽMw��iJ{}��5�퉔̭h�A%ܩSl`O����3=8��]r�]kg�Y�m�%��61S��1��V�dV�z2�FC0���ڛ��ޕ����_����=�;����6�F�[Փ[TV�j���������O�N�l�$>���olfժ61�qU��w�3����`��@��׽.�	=���Έ�eZ���j:V�!�~�mu=9�r�@���3��蠳*#��"�_]
�<��TȦ���3����9eɆ\T�Lo���Y%;p�C�����񴪺-o�!:��ƕ��~�=y���m�c-�lГZ|�
�,�숍ѝM�
~�
@����$�Iyr��F]wt��^�Ь�4L��QDP�i׼r�}��|��T=���To�D_����+Uw���k����K��>|��˶ɷ��G�-��ڗ3u�x�_Lڻ*"�f�K=��W�z/m�U��@�O��(�tf�3c�YA�`������/��wQ�����1ۙp�}���8|����j���#�m1�r���
��6<o��NӼQrj���[�qm{ʴGi"#�\��^[~��
ٿ���)ǳ�1-�ճ�����x��*�B#�mߧ�hk<��Q~<L��{��$$�HB����li("٨h�M��?�����E�Ǳ�\X�.;�x�>y+��Ѕ��e��5�]Fp���
��g�ؔ(g1ە<�����}9v�v�+Si��֐�pL�������Q�nc*ܩV�U����;./��1���S��#�Kx2i����r�,8wy���|�  @
@�
DBڡ����S��+�T��G�r4,�2()���1�(ˀ�g
PΤ���L�O�!B�pY�Z�]f��y�a��t.��8�z{Ԣ<nN�#�bX�6����yT@k���:��q��_K�mI��h��ר�L�)�:��w�:-)�lO�h@��,1?IB\j�Py�Ex<ݙ(wl|��	�VE��ܨ�b�&�9�y����mU���H=Q9z�ƝЕ���>HE���[C�س^���o�d�7��3<��7��CaI���gĎ����X����p�����X�
��ԘG��]b���B�X��#3U6z0y�XkW�Uݪ��ן������6��G�}���~�0 ���#�<�	1��u�x�r��t�pGa�}3�3�uٗ��;k����8��4j᭖�!�lht�θN&l�}[%��*ѹ��'�S�l�k,{�����ib;j�_܄���7�h��P��# �0t�<��������S^t�Ǻ�E��GOsZ��y{�U�ʭ�TaEr�$PD�7ưʰ6�!�&7���W�\*p�����Y�RB���܋�-3�H�3G#�4U8��Y�&�j�Yղ���-.OĬ5�sƃ�v�keu5�.�yMͷ��\�s�̰���s�haR�{NR7�8F����$w]�6��J����in�3�mn��;li���� ��H55�����A���k�r}}x6��/�d�>s|�u�ס���Q�}͎5�Wc�����ݒ��e�����d��t��%���NF���+���~�e�g谽,C�Oբ/��l��J�,ȹ5n7}�vz��0����x�W�٩>�U����ϥv0-���T�8m�5����lw!�O�n���G�ܕdDy�#0D{�5�NÍ�K�Y���!�^��}�\�]/kB+�E���ط.�
�/�~�s�]��}�Q�*b.`�b~��ᇞ3�-ߜ{���A��Q�tʆ�3L�mخ�>�"��-���{��jr&D=(��f=��ur��#�3�#�X�*�����PC��ue>T�������ow2C�!�M{ݱW~�(:'c� ���T0#c�EC���cKf��d4XDtpx��z.cZv�k��q+ٶ��E���9@zpIb;��V�Yb�{�����yMa\�I�]��Q3x���Ϛ��@3$�w����h@.:�C�Fx��Rˏ� U/��~������/��5(��T�r�ۤ�N�H�I�s�_5lp�Y{��x�ݺ�[Mc�����{��sfA��o�5��g�k�r��8%����]A�&�%����\�&֠2ъsYw�Âj��`�m�I���z�kt:�EM�������9{Lʶ��ӎ�$D�BD��" ��Xu�U4����>��u�q��G���鯑 �z�E	.�޿J�S��`�����L���,SҙH�'s�)�
��Oxt����D�~��5݇ ��x`���Z���Z���t_�v}W�LEz�J�|Tg��<��pAT�Q6TF���Ց9wO��������	�2��0�X;�#��J�H���ϒ��iJdǖ��Ww�үՇ�}wh�[�Ur����ŋ4L�="��'�h	4Ϡ߲�_� H�Nh5k�$�!���WY�ν�/�����X'!�8xj;H��ȞN"(O�M���s�#=��Y�H����'����Z)�k�G�$p�����&�t��^�9�h૟E�<Ob&���B�+�Z���h.8����-`n�lh^�YSrU��b\z+¥F?BQ��g��Yu��L���;�lwg�n�:8�.=�s�8y^v-���c1un����U��
��^����R����)�u`����`���z�B=�s��,S���2����qbZv0�s '.h��g���6t�Ç<|s�6��=��Y��kWs'�m�c�Kdlܛn�Y�S1�8�s+���՜5�ތ��ݺ&��q�ژ#��TۮHֻ`<-�cT�U���ꙕ��	���jJ"R&�d=J����v����l^�3zN�b�m�HuaJ����M�, �<M�*0n�;���V�Y0�=�w�;����TD4s�/�Wy'V��k��r^�H�T��n��K�%�ކ��H��%�͏8�q�S/��zv��9�E�i�l
�����U�f�l�Kf����T��:&ֱ'���&*��v�E��%��W�����*��;����=��0>x�U-S�b�V�f�(�����*�ܖr�s��]j=Q͙b�1F�^Pp*OX9��7�`��K�ƆqQy�м�.�����;��Y[,���ͮ��΅^i�ä��!K^��J D�	/!�F�I��h9xR	7�m;�5�����ֹ5�,BW=��uX�{3\����k�C�P�*PTޜ�K����ٛ,��"�Ub�$�l&w-�.��HSnf�K�phu5r�����Y9C��V]����QU�2���E(y�4�A��m�;M�Ts9�� ����u���X�E@�U�Qbya�\��� ���ֲ�p�)!kF�7�X���S�%�5��qJwW��������E�-���.��&���w�[�ئ��)����Ml>g*0����*lV�gG9�,���g���Hl���W�`U�K}\�]2�vV;�9�P�4A-��Û9�+��d?1M��/{1_;��{��ˮƪ�-�s\�N79hmW2^���ɳ&-���A��Yk��V*\vsi
5���[��ܾ!��ٴm�}�"����s&��N�7�b��Ɖ*XI�״���1�?n�	cl��ǐ�0l��bt�Xv���H�n�9��4�]1�.�0��d��4�Nd�,�pʴ-�j�t����.͵��@�3c�p��z}0P�&��:�Xe)6���^�pӗ�*hϙ�;��w�J\g�-�I��Ӗ6��>D����]#!v�Z�������2��������[PԴ�c���R���=�n��i}�9��&{{Vʇ�Q��oj��	��O�yN�f��ř���W�֬�I[�2��_mI���1k� �XB��w���;.P���]��\�:o��F�^�����({��*���g��]qꇬ-2��p:EE�@0]_[o!��)�VCR.I�uݯ���B	�ω.��$��43j
ǗBg4u�d�7.V�R�Z^��͸��"k7W�.v��6�d�B�!_�f(����֑ڲ���F-���[��������J�¦nM����.�+��Іpp�ri��A��X�]�8V�Їer�;p��SKj*KK���QV�<)�V	 U,:
9���t����C��lͥt#��-�	�p˸`�G@�N����6��6ؾ�˿�6 ���www];�"gu��]Mwt�)�pȂC D�v���;��H��Ww)��,��Ď눙�WjG\��N�snt2`��\����9���cwW9\�AL�w\ uؚ��$�ٹ���nY&b1�Wc9�;�����n�
 �����$�wt&���Iwt�YL"s��4ads����� ە�ꄁwt���@$�ID�B�4�3sv2�4�B��; .\$�Cf�Nk�&%Θi�����9���HM%4�@Fs\�ۗH�\�s���ut��؜ݰ�u���M
��!BRLD��?[�����>����O�{������R晬�\����V���Q5�����4�o&.=9g4��̱96��������^-���u��@$� �D�v�����lg����hR�[�3y�B���S-��#5�7	��w��gX�'���<w{r��qw��0H̳�í�̉t��*0������(S^�'qM��o�xD���\x����wN*��y���+o\�Z�eD@�8�k�}<%�]z���t+�ex=c߸S�(�y�'�O�/���$z9��'��A��j�� �ة�;~�T��;�xf��w��� t_����$�Q���qU������F�3�zA��9�Xo��+ c쾣����_̹̃sP�Eu��y-ߠ5��{���r��Ϝ�E�a���Ӑ(z�s"��t�z�/g1�R���4$�=U�*c|}�7��9�~�-*��-"�RK{���W2�v��s��=]"!�A��Z4$֟#��Y��"6�u4'U�>>��Zθ&o�5��Ll�*�+�?@v�������#�����[�#���-y+�2��>
�==�Un$,�n�a�J`�F o���՟�%�I��R�a��^�G!����]��&V`��D=6kP>���]�c3�!s[Aw75%�^i�D"i�ܩ��P���-��YLQn�A��78N�@y�����S�A�v��,�(ݔ��{��V������h�B�b{NFKi����gdw����d4e;�;�>��$�7u[y�˫>�,�����o��U��Gì'�X�H�sf��Ía�����'��5�s8�^�Q:��L�C��b�h]GO��~�kй����b|�{{Ōkl��^f��2մ��_C`�ͅj���,�00�v��3S�f:m�1�&o�r�R�8@?:�r�V�v"����&߯e�i������o�����)U���h���w�İ��sP��2{ʢ�Ѽ9V޼Ժg۷ݏ���SX��&w���#�4hY�g�
G��#�.��A
Τ�+䤾ɟA�Jn����鉕���Ù�/�5N.8N�tX>����B1��#n��C�[����>~�3��o(�/i"��[g�L�)�:���Б܀�����蘏�b~�z�d���i��>�d�}���	�^�#�ʲ-��ъ�.:M�g���H��·[Up+��Dm�bn�7�7����&v��)~�U�����jc������w����4f�:
M�=����ܷ!�褳=Y{��.^��o�&$��zG�q1��|\�D�y���ўj����;D��������}�p��?K���=�{Q'ʏs���l��+�-pb���W ;X�
j,�[�VZ5�K�]%�pm��n�Q�ΚF�%z���J��X������g={6�-�]=��Q�f��˺�	1��Itȅ�u�V�K���������|>�ֽ�Y�=����Q��1�[�H`�5���Ѻ�<wܪ~�-×^�m�)���)�u��_��Q���+�7���B��~�X��^��P.d��#b�K;V:2*�צk�.W��Y�ħ������a!#��%Yp���M*�_m.,�������՝j	z�}Np���wX�5��Wʭ�TaEr�$PZ'���W�(����3����ύ]c]���C>��j|�`��F�^����+��R��ס����1��r������:�|wx���2��!"�1>�''!#�]�}}�vo�a����������}�v�*q�>��a�x��v��-uz�FAf��3�H�xKdǼjUe��\�E}o�r6�f(��JL_��No�Z�Y}�*���t)�E��$��$D��0D�=�S\a��8~w���F7��.��M��=��Sl����[�v�\[�W��ܗ�A��J��9U���ؘ���]�l�4�{���B�*P��e�g�2�6�c�N�#0ش m�'�;�(���LX�+�x�a0�W�p����]���9�i-�����0>�2�b�O4�Y˾ꍗ�u]�&��e�#�N��'S1��ٓ(V'�ƻ3�I���.���)�m��9�A*dg{7k�*�9];,��w�qf��1P��]��q�u��u'x�1�u�����6O+�;�ݠ?8���0E}*X�Θ�#G�i�-��p���	��-�	�J�G���MR�U��ό�w�80}%�z�u��"������hb�l�9�h��l`싆����N
��@�]R�~��U�,�=&����VR��Zϼ����O��k~�of�}�s�����kj`k2LGx���j`�0���3(�*UеL�w�FqXjk�7����!1�֠X��Ы-����X;8�t�Bc���!	�{*�D�Te�H�Я����;�K�;�>��2��G���#�j۬���X���ww�.[}Sq��'ʼ�`H<ϯ��0��֠ty7A !�_� ��W�%u��F��cZ����|�*�4�A!.���ez�&^wTGW��@��i��#�l%Ta�������ξҪ.�m�q�E��Ѣg����LK>��w+�ׇu���x.��).�c����$^�����:����C���r��Xf��kq����;��Kյ*�|R Ϗ���{W��r3��r߫�dmt#�XY��^r��#��9e�e�m�͙�>h�jU�0d5rA�=�{)�Ua�l,�=��/or��d��2�Ʉt��.A�`-qF���d� 7�k���,8�S�w �Ƈ9˦]z���5(��H��+����W�A�ޞ
�ԏo�`�~~���8{A�	��+C�r-�ɂ���J�|2�,AQG�-��r|̍�;��xJ�s��ޅ�U1���Ke�v����\A����+*n���!�q�.�|�]vmF��\�bK�+�Xj�9�T��
q�9�p��طM>��}��x��kwC׹�wm�Y���b��B��ʊE0}u#��޿���u�c��p��V'N����`	�'�!�~�Ǚ��{��Xþ3d&~�pQH�28#c�{���e#��f��5��}�7�=���<�mm��\B�w氭�a��J���$F?��߄
?;�{�j�<U�u��q�'�]�p[uг�٨��sEF�#L�nf#тxK��]A´jF�Cي/%<��Ʀ5�.�'}&�9�z1�P�>�'���h��G]
_r?N����g���]xz H{��YJ���^��v��縪�C��~��A �zA~sc2Uc�9.��UykC�����6zvj7�W[���נ5��w�s)NYv%��q�y��ޅ�~�qGY[����*�qX�ZkR<�)1�]؇�J�뭯á��[���d3;"}q��>�yhY�~������5c {B�^«r�'�P:
��r~	�0k�V9̫�v����0`B�e6��-f�A�r�NJLR�_mr�K�����w=g/X�$ ������Kzj�� ��GR' ȱ-����1�tެ��Jv�d9�>�ξ�[�C�9��ۻ�mٟv�%5�L؃�H�<�:&~jLV�_�v�K9�cw:�=��B����#r۽�Q�����,j��r���	��_`�
��g�
��<��4������lu��Ut�A��5��'��b����)
r�1��������A�����{��b=�Á�k؃܌�/nq�^�cb����*��_֠v'�NY ߦ��Xj��	�+h�b?���~r��C�����K�����U���l�G�\��v-�"\��������q���U�Y�΅{��ێ�����L�=�6~�6����_xo!N=���p��م�b=�V*�NS����b׻���}�xo�c���W������A��Bǩ�E��,2#�/=B-������>�q��E�m�\<���`��E�� �B�A�e��2����xPB��yь$M�9��O��+���ɭ:���2�Ȩ|ڷrz4�rK��~2�dP`T:����t]J���D��P{�>��*E�r��,BS&�
�գ1-7���ur��fOi,�	з�Yǁ��Cr{�^ut 2�z�*��XN�yӔdU��#���3{�8KW�mKz��&8:�	�;��u6���n���M���������*�����sO
�~��uDC:�/过<�l�)�e?GP�~w�:-)�o�ʃ��v}uqs��3��^	m�sYs����اcmZ�Ud^�N�P�.:O3l�B��7�����|���K3z�+�����6�&�*�PP� ���\�w{��fySFo�
�3�U�,:c� 3��.ys=}���٢bzz	cd:q�&��]b���B����Kga�y>;�b�ǳu��M*����O����`d�d���B���xR�Q���ѿ����ܬc�V���U��t#4G^֠[���u}{���/�w���";��6��K��#Fx���$�<��z��</��w#��)�;�<��}U�H٩M�X��Qh�$H�0gD�`[\x�Έ��V�G�V�MO3�*���Ƈ���X�V�_*0��)�E �N#c�a���n��o�gA'ק�m�{X�6 �����|\��m�ú���+��R��ס��j�{�&c�핗.�b�p���~�"�5�WH�px)�����l�\�KF�ߡil���8ߣ�
\�)ө�y3V�ָ�*!h�y^Bh����u�:t����4���$8�+,���Bס�kV��4	�N{-���\�q+��O	�T˰���"�
Mj��c��7K��MK���6M�ك�����V&s4d�4k*��ӄ~|6V{'u]���P��n��kЯ�2
48�20)�<%�@I�����^��R­����a��~y~�!���r��V1�����=�追s�U��Xr2�M"=&x�=Y��z�x��g�>{
�Oq��ezh�-�P���n>rr<\�y>�4%I�wx�m`G�+溪!y)*���[�+�gLG�:�(��p�D�+�n�<�23'��+�9�Oh'z0{�db�u�;�w�����;%�E;(B��QGyLǗ[�A"�i�Gp����#�m{��G�{7�h�O��
�H��E}%�z����>DL=^w1X��5��d4[~���g������o!q��G�f��z�a��Gq�ºm���X��V�X�w��s���{�*�Uz��-������a���_3$�H�I�A�m@.:�C�Fx�~;��亦����c{�=�Ǔ.��������VE�/`Z5`�tY`
^���8y���$[��S�����נ���X���_�����;!�=)���w=�ୋ〞� g��Si��^W��^�<ͷ�h|`��*��{o�b]SAa���g�W9��U���2U��^̛+�s~�/e� Yď�׻����u�Ip@A|6\��U'wbfn^�C%�s�g K8^;������f�=}�6Ѓ�:��Y�cjRۣb$�����v�-=9�8~�#���EH8ʝ����ɺ=���S^J�:5t�#�D��5���v���ׂ�D����X�L����0�y�Q^^��M#	LGa��"�Uo�����uo;�a������b}��|?(@p�Dĳ�;�����3ӈ���i���+=�Q9��`/T�"��C���|�Nǯ��0�l��<���DT���ʹ��U[<kbi������/�x���C�,���術�./�rK��n�P,|�����#��Iy�f���Ŋ�ؽ�T�G��A�ϖ����X����3y�V�G�����>{�!?�}��yVQ��T�T�'�)�z9�T�G%ǟ:��b�ϩ����un�������y�<|c�yό�vH�!����HlW�����]K�(2���8;P���[�5���w�I�\���>����f�BE��`�`��p���V���/:(qRB�v���v^�F�Z�á��m[��|E�ʖub�Ε�w�;ZDk�/M�@�r��:=��ɚ���n��5:Nz�1�U �G��~��ݴ���p7��f�� ����_�v�7�D��=�1�)�,U��9+vXiۛ]=�<�Q��F>І�q`�^�Te� �=�T�,ҙ�u��gF�Di�aP��8F*Y� 1�M�����tZJ��G|��2� 8��%����9\�q�M·�s���I�A�Xs��.;��c�c��}�"�{vfX�k	��k>�Z$]�w�q�g��r�>�'����H��Aځ?w�P�����57��Wfd_v��b���.ӫe`�Y�#�j[c0y;To�X��ǜ�Т�6���"U�������1bn���	�!�w[W�WZ���������r��.�Dh���]�?v\��1���n�G��9 ��� ���7�L��;���ћՐ�Jv�g�笮�`X�������q�blⱾT��_�R�ܘ��oʼ ¥" �6���m��o����K*Ƕ���~J�}+t���׵�:4�(��޿�SW�D�(���\�a��N��E	�X����m���n��^���/���.�=Yc�ڥ m!!r4c����l�������Bq��N#�p�{�T�~�$�/��ǽC��{|�"��J'��Α �����kİ����I�.s����f���pa��-b�}uN?�W���{{�-�dp]���d�bl����:p᳧8p���]x[�{esi�0��*!��TK]���K7a��T�]\h�.y�n�d��jBڥ�C.B%e��� �fZ�!�љ���h,�m��#��q���N=J:��G#̰6
HV�#��W.FD�)՗[��k�V��+���32O�pS3���'V���B�5��Ree���Kb��W��a��0R�#Q�ȡ���݈ued5:�)�8�3�1V�aѮ�S�
�fn�t!� �i31x�"�aX@ʝj;\W)֥0g�P���d��a�9(�Z��S��N"�S��h���ѣ���\�0���2��K�����ڪ�� ΍�rD�-��T;�a6�<Gj����.TU�!����\��x�P�q:t*�Ee5i)A>�\�`�;�h�B9̥Xg�,S�6:} d���0�	�2λi
|xT��F+�G�"
^R�Ε��ܷDT�b�H*�ma+�wyq��`91�y���I���Y���L��\����U�@Yw�)�V�'�
Ʃ�e�\��g�W��r�Sd`��I�9�*���=���U:��멉�y��~�W�>�����ǩ��%S�Pɸ�du��;�[ڎ� WB�h�Ǣ�U��� ��N�o_�41�ɽ�4��1A�휫8
�x�H�g$�vլ[n�ݮ�nA ���؃�3�Uv�C�DY�^����l#9AD��,�5���{wx���F�=�4�P���ň�vm;'G�ڲou����d�2ܙ��tFź��
%�N�t�t7��^KyK�u1U���BwmqUٹ�2B"ݛZ�i��6�:&X�6��~����O}���ބ��Ϛ�:=���0�y윏'����5xfFr_'g>�ۭg`�6����%�k�2�wsI	�{n8��Q�Y�x��GɊ�%,�W������sB���1����gX���ǿk����o,���-��mRϱre�;���6]7p�޷@�F�hq�_�}����G�r��%�rS�J�Yb��J�'&�Ik��뫆���'�
�+�z�`҆�8�"�)'�f#K���[��=�Ɖ�"s}�gKx�J�.�p7WJ�ImX˨�l��Q�d��p�b��9!u3@zkRs_NJ�mn1�065�Va�H;���>�H�p�;ydJ��r�+jJ�b��ϰ�����t�1��WS��O�]��˫�t�����.�o��9�*56���|�
�������y���c��ܶ
�`���K��S�w,A�r����B�NS���f���]F]7���uGV���ڭ{qܧxU8�����P>�xGE��r�sU�Jt��yfi���H��Y��
e[�2���9�Y��ٍtX�Z�����`�W�1M�fF(�s�Lݷ��S�z9�Ѽ�J0�%����8��_v��͓��0���dK��d��p�:�*.�g��w+����t#y��*M���2��Z������r�b���_����_�hBe��������#I��f��b	0Gu�#��Y��p�s���D�IDI�#�}��`W��vd	�".���$QD�9�s"�	 F�����,D 1�1������Gu�C������"�M&��i$�⒓2X��DGu�����BbD��n����a2`D�D��ܤfe� % 0@9�I1�,fNN���Q�)��"Y2a};E"�%��%3�\����A9vH�`h�{��(�Y"�]#˞�v��ȑ�W����M3)�� X��������x]jZ������壳�[�$�W8�r��Ó�����8|gi�۩��ݏu�.b���zL����O���Z3M��cɯ��?���{Bɟ�Ȝ#Br~�)ߠ7��_׼����lC����`DԺ��}�������l]>�ȫ2����9�3		��_z��M���{f/�ey
2��
!a��y)�N���g|}� �Vp�������b=�p�~����g�y^�3}]�A�U�x�E���y�t.���FLo����$����#�?�`�:�N<�S��ޯZ�'G?�i���T@X��<5[�ϔͲ����j��t[n��8t����CL�ȳ�hB�z�߱hu��?Ib\u���`{�"��'F+�Ƴ|����F�����t	m����s����2_�i��p��:��ˆ����Z�mD��u�R��|���Rn���%ݹ�����}��_Ï:�@���!P�WaW]b���\+�R������[�ߞ�=tw]*�U�Q�]��j���f#��b6�`B�)Ș�-�x���@��/�-�[q��sm�O⫠ ��ü�����o��G|��$�P�h=B�G���P�;�4M�97��Y�c�c}�&jȕh���lMa�2����4�`��1�#�O�&E]L-F�fL:�i��C�R��t�j�hU�Er��㏨�r��d�lց�
K��ogeJ�_>,�tS�CB���h"���FQ�6�n�I�Y����GO)�Qu�,������y[k��CUpv$ka#��E�p'zj�ޙ�����S~������;9�Կ��69f��Ƈ���X�V�_*0��)�~�P4V#[��T��N�ֺ��^�����0t�)��<?suص�޽�.j�\Ej��su�b${i[�؊���r'�ݶ�4r1���D炑L@�7����7f��[~��ǣ�*�ey�ժDTA�#/�>J���C�H�(��	Uu�X����9�
�Sv���"Ӊ�k�V�=�b(v(:�y�1�t#хi�8�
�}{�S�>���*��0�e`�Dy���k��c���3+�ч~����Oq��L�N56�Ǯż�n��*�\�G�8
�����ı:}�:s�V��T�'�Zb�mDp��Nq.<�2��c
v��OW�d�Fj����uf�؝z�>��1>��K`���!�Ψ�"�ʦ)u�p���	���l�V)��S|���ˁ�ʼ��OԿc=��3|F0��(}%z� ��H�kΦ4b�l�|~�f*��=���P��C+>ל��{�5-a�+ܽ���p�����)�y�̺5s���M̃��l��c��@\K-��c���u�*����Ը�N�S�j�(H��b��vؒ!���v��xf���S�7�v<����&��-�[cPG^G�d�����5c��r^iz��]G�V�/�Ф(��hj�:OD�L�AȖ�I�#��e!K,Z�FǤ�¾~�9�މ+��@���1��I�G6��d���>4ѵ ��9�Z3�Ӫ%�}5�+���sD;t/cg��i;P,c��U��`(�c�q����v;l��@�B7��q��ex��x9�����B#w�s��t�Gc=ON�#����B�	���=�x�A�Qum��Uֻ�Y�b���@A��H/J�[F���P:,&� �k�"��Lty����ݟ�g����`�~��/�U�������4<���j.w7U�fyz�����^�ʇ�T����%+ޝ"x��P����H�,�I6U�|���@ϧr�{��	ʞ�7W��>z"��@��yPO~�L�#�*���}t���͑t)�� �Ke����8�vǭ�%ϺN�,������������~���9��0�ˎ�r_t��Ux�{e���+�l�_<C�U~8.��k�S��>[,C�zF����q��z}��VQS���hW�$�˪�J�]��t�4��U�ܚ��$�Sr�75} ����6�Օ��]=�X4`�}��c+y�5|i��;�^��ۤ\XUђ��M�w��)M&�jÓx����^EjE�R��u'y��G$��Q���r��)�ƶ��S{FS�	J��NF���=~�ʎ;2D��o����΃�o�ų�S��ʎ��r0)����s��������񘱇�bs�!W����G�!�z7��p�e'�1�P[P}>�ifk{'�to�g����Ho�43�k�*��`��3c8HB���7����s���7fL�m%g3Q̿�W�M[�g���˙g�v'�
b=Be�|n�P�RmK���G���)��g��1��^�|k����?SE�5����{�eE�H�0"�1�V_��1�^SaoB=ZC�&+�w��}�n�"���I���3��P��I�l� �l��9˲ˇq{k ��L�&q��P<({�����p����ϩV@Qc�z�bN�縪�C��#c��D�c�3��x�+������p�·�:�.7cl�ȕ�B6}�YC]OJe#tI�W��c}���vkݼ�6��5��{�BæbO�L�5���g�X-��f�����rٳ�	{��	�gI{5)�}�{�~��xg߼��1B�aPR"���I�>G�Q�z�|�K�/�8���*	�#��S�Ú��b�J԰��m\]�l�N�9tUd�^��m�q�7��/ϮKZ���g\�`�>�B����<߽�,�A�t�Bܣ��^n�P������>#�eK���ۈ F��:�lkxqu���_Z�^<X�0�*���xO?���^S�#�B@��	M��,�}
/0I�]4L��P'A�!��A3�����R�I]E�^�3��^�X޽�1\��r�!]FxY�F�ܞ��4�|Yd�>�ܾ�+=����j6�2}'!��9��z��{|�"��JZ~��9D�~�fn�-�!�سW���x��?B��<����,Y�_.9z�	��n�;�����B���m�|��Si��Nv�=�g�,-�f�o���,���������];��V��Cy
q�Z#*e���Ϟ�/V�q��,
][q�7fQ��tS����2��C��%_�1f;tDy���U��1�<4���׾-�j�����E�@��f��3�#��1�yC��g0,GtM/r�	��PB�RF�L�-�3L�r*ո�ϧ}]}9%���I��6�����Dt5Z�!`�^�� =�L�}5c���3l����+�2#��ϼU\^ǃ�[�;��+�]��/�p%'���=V���{� G<�8\k;�q��:	����ujUk�EA�U�ͼ�X���ڸ��G�����2f	c�豏�����nJI\�Mc�Y�5iF��=�u�C�>�������V�*��Y��(�ğ���*n>���Տ�,/�U���{ ��p�ے���O�V������Y5D�.�'�]ƥR�j{��غ������נ�zC�!ϊ v�A�[��g�x[�_;����)�+��i�]���vJ���2.K�l�g�S�GW�h���_�_1�@)�y]u���-X�W����B�2�;c�
�~�}�:��j��-���#׳��n�h��r9&4�k��B$n�$O��['�:������b�U8b�?�������XY���Lv�~�z�>�*�/Fs�|���L1'���t�vǹX�����A���lH�$k�B<<TXG��3&Mp�dD
�w���x		���ڀ�����w������`���ft{�u��Mf�w�W��A(�q�{�J��f�<ĉ�,1�
��jS/uz7
{��+���Iru3j��
�Lu��xoVuo*��u1��h��a��(��R)��rr8.��5��Odi��uP�A�o��6������,|ߩ��l�ס���EcP��D�&=�P:�5�xe�8�ݼ��5�v������v;��R�}^��Ox�,\�`d�"F/����Q� �/MϪ�PQU�΃�Ui?f�+���f?M�����#.T���8D�`�L��)~5�pi&�ڃ �E��=�S��y
~��;��3|L�u�䇚�)P#-Ej脱{��FY�G���K4K�X�9[�s�����U,L�Www���2J����~P����z��X���e��b�
v�\X{��X�����I�j/�����Ϗ����^�G��/��v]De�Fw�Xͨ��u(Q��L����W"-`��;�vd�#f�W�A���/@c�s�.�U��E'�R[P��!�uD!;ʦ)u�p���	��s-)"Z�}��^�o1{%�ް��GA>�0+}"@a��P��=u�Gȉ����V;ν1݈�	w�՚^��E?�H觼hj�1O|AȖzk�T	B:M�M��l��#�sSS��Mxfხ�X��[��O��;��rt�[[s�$	_�+Z�(��΅+8�~��*�0o�c��L{K��egԲ�,R��;P,WB�u�7�r�ر�;]79뷝��V��ĸёBC�=#8���v+O�vz���9H�g��R���c،7�96j}V�.���x@~���?D�"<��m{~�P:/ɻ>�íLEzM۟r���۳���P��#��8 �"I��>�D��Wx�
�0��������>�ic��x+C�P|F������j���Ґ�O/ ������Ӵ'n`�& ������ګ��d����'���K��MUL�����m�O���2	V�i�m���fiȦ�Z��z�ps--eץ_gV����cAS�v:^e[�]��ׄM��nu��b�Z�-W���TB��2ax�ädkM!�?
��|�}&���>����c�\��
���� ?�O����$
d1ҩ��-��t���D`�R*�bq��7���T7sN�/���us��{��sҘ5;҇���5E�aq}�]z���pk=1������C�{�P�2(	̫�]Ϣߪ�.<;���b�a��17]�ޯ@��\�R��}p�5旒S��!	q诼*z�/��o>ۺ��(K�h�S�L����x�k¯�>���}�og����M���G�ǃ9ȏ��@��ࢷ�e�����Yb�]��7�nst#�4@��x�)�
�ӱ�Ә}�|e�|M�-��d#�9�!qG��i�Q�Cݧ'���w�Ҽ��4_���XM[�g���˙g�NĊ
b=_L��_���w_{�]�:a���Lg
��jN#L�9�4_�t�+{�1Ȫ*4#L�nM������mL��9��*��e\��~�GO�y[$]���I�1�3эʅ>�;��c"�5�}��ۜax��H��b=4������<|��4!��j�i�wט�n�7��Z���p= oLG(�b��淶��ٮ]&�|�	B���5�c']vr�n\}n�V����%(VJ�u�{�29-�=R�o�������%#��cFԵ֏I�z�GN����[�z綸��@��`6�!]u^��dK(ZN��縪�v;����=
�3�^nSC�nGj�0n�p���:�H �=b��5�u��y-ߠXk���&o��@�g앻��f����QnOEveDm���� A:A���4$Ɨ����f�d?U�����o}�7��.����;g����Ҫ谷��N0��" ���^J��E��"�enF�X7労m�;Ъ�#��6��X�#�)Q,�a!#�iM�_-������
��#�}�&o��a�X����S�R�i��B�נL{�R�((�Ah�DvL(ч�ڬ��c�SM��핰��~�`�L4�T��f��<qxoX���TEh�P:�~���H=�Խ=*3��n����[JF��,#Xf(	�g����
\Q^������z/���G`[LCw�D���R+G�n�ރݧ��
�����X\+ܪɕ�j	C��g�՟ّ��v�uG��7wm��^����-�ճ��V�\s��F����#��>���! s����[fB�B"�-��,�����
��$�{vw1�q��P�C��5�:�6t���	zWV�R�t�|Xux�<U��.�8�&$G�����h5U�D��~4)�����f-i��YX�����i��1kyS�ƥ���dں���!.Y�'i��v�Bf���:�����^��]��L��9��S�������SV�0L�m6��4����������yh츷����OW9�n��y
�:�7�4�e,����R���'b0ܖ`B{Y+z���;��;_�FLG����s��-��2F�t��3l��B���@�8�=om(;�י���{q���� N@����.6vxGgM�"�����g�x�sږz�2n����ż�aa��`5W�H=@@����v*JE	٨|r�*�s��?!�����ʨ�Ԩ�}C�ɰ��gĎ�4LOO������q�0�+��|^UXN�)�t����G��Br��3>��Fy�Xk��~�=cg	��ف�$ y��7=�Wj�7�N[��pU�$����,�N�<.��
v�}ϫ��\�E���X.��W}���K��ì��x<���/���X��\y�����l;�_��BM@Ԅ��F�4xx�3����}�R�[vVf���A�0�s�SR�VV@��GvBֿ^���D����yh�4\�ɳ��6t�Ç���`��1�ea���pv����{��8rt$Aڇ"J�#��� ������T�%4�e�_>j��źp�����#Ѯh��z;�ECǕ�a�e]�(̦�b�W� 
�)��(����lK@�֫)L�뾎���D����}]���W�.
��\Uڑ�t�� ˫0��ӽ�����*q85���Z�V�/6&;���^��b��S�c�Gr>Hƞ6�2�����2�^����>
�Sl��޽K���&�\<��=���/YW���+/tsti���f�IIi.':��w�6�K�וW���/TP�A%2��m��y�Ne�+n����״�F>�L�R��7S"�v��DFm\��7A�%�b��Y�Ʋ����_^죑�wzj#�p�+9�^j�45�0$ӛܲ�X�)-L�W#��;^���o����w/�ˮ;GV�7/�ПFrZ�#��Gr�cN���$�lU�7������L����H�-�����k�3����9�|z�^�/0,BvX�8kB�m	@�j�őF0T:�_F���V[��67�(
k#��Bh��}{���V�8e��j�[�KF��*���-�ov1J臃���yA�V��9�h�T�;�QEud���e+�ol�zre�����!H��N�=�S:څT�05mt�u[�Che+�(�z7K��uYc���uL|d]�66�/NC�;�_���
�q���^9�����}f��N����A,ea .���xEԞ��ۉ��$����S�6f��+�-�������.�[�X+k&�K+.b3�݋:�&������[�˴!�{r�+�K�We�C�KZ�6��m*ޝW:����
H�h��8f�w7OF/�z�Djf���h���������`ei3���ם�n�0�w��6�bo�*�Y��JN�3��Ҭ	1��0W���VF�u�����r�/	��7��K��p�E�Fi��eut�LC0�̾���3d�|�m��X��������y�f����C8�;�V����-��d&+ޭ���ώ�F<�:(��CZ��y�z�X��ǹ�Q�:�o =��8<I�s:�`��c�S�͡a��<r,<c
�ӱ%G�X�� ��YҨIv�Z�y���j9SЂ�����wE[�����f�C{/NԊ��S'��3O=��_,���d!��NPdQ�V���<Nq�w�RE�z$�'F`��K�̭�]K|NS��J�Gv��S@�":�gq���*W����fTk���V�����cz��E�tl��x�]M�7Fz_g��#
&�W��<�cWA�w`��NY������.*�M�q�j �j�}՝��k{�K�zo�ճҝ�-���Y��Y��0��oK쑂���\�
n�f�?d�΂�D�wP;��6�+�Xv�I�F�4�����JH$Ф�d#>������>��~:��3""̑��)+�ۓb���7H����t����9t#����HS78�!c�
;�� ��X�΍����܎�0	�S�幮s	ˉ��N��[��9wqr=��K��+��=�쀢��p�n�w9�w(4ɬ���.�ή��f��/.!��&�s�v�����1A	�((�Ayn�t\Ԅw��`�u�i{��{�d,��r�D����旻��AY*"Hؓ!E(�WaE���"��]ںh4bK��b1E%�c��nU�LB7'w7�A�R~�����[�<�G\�-����2jK����s�TνI;:WY|N��eN䦚��0����@ۨL��D�)���O�%	]���B�v�h�.�łsM��a��N|�0�g�R�y]^�¼;���*���3$o-���V|��ek�0ƪ�!	)��;��ưʿ���#�H����	'!���+��4=�kv�b	���b��շ�a�s���b �P���[�9G�dz(���y}�\�ɹ%/�X�p��Ħ&{]I�Mz���Y�z0-�~"a7��+�=������"%mC�b�L��{9��1�kJ���������2�=8���~�n]8���ʯXt�M'wZx��^��zv��J��s�F[1c6�8W���E��᳁L�+>mX�+;�rR�{/D�v���^ת��o�ڸ���9�}H`�l��'ey��v)�Au�p����U;����]�X��0!P�m.VSh�����7�'��EIA���� ��H�x�'s���Qꐁ"�WV�e�8�?�߫!��
GE�hm��|c�A�_r$0C�a�'�-z�mCų�N��'��{\�N�X��u�c>3�)�R�(\)� v\	�LC�t�����0x��9��PI)i;���<�+Wf�n�=n���b�3IޖnS���/���w�]��y��/�(�C�*�}�%M��6_�&u�Ŧveײ��^`ܧ���r!n�W�c���ʒ�9cޫf͐�AҜ����e�޹�K/�����o����~��>}uܽ�䎇�t��YK,b©x�ĝ��z/����9`�_�p�w]�O,1:ϟ\wW�Ńp�3$���?WP���c|]?��SӉ��w=����{}bbn�z�}�t���O��� 0~����E} ��b��=�R���y7a`��h��~x׋f���'�s/&�$�vc�s���"w�=�>n�
&G �%��3�{>�Q�����K{aM�n\lVm��"n߷��k���N�;�)�Z'!_H�(�I7�
EW�'�Ԛg�/Y�֤�/�q{��3�{��-.���8����r�(
�PZ'!�Ma�V6D�"��w�hழf�o�����s�?��KN
���i�nzZ��҇�7�sU�Y�.8uNIyQ�_�Q��Y��0[�^����	�8�P�V���_`��FB�!��X�a��-cv��~~���>�����'�Z�ށ�Sr]�n��z=�R���'�P{^���c�zP���E��Lp��ʯ�����\��wy��魱��u{�}��f,a���P���0컃�['�Eo�O��fmSs�*�2����v�xNl���g>�����-�Q��{��D�qm���Ű'+��ĵ\yr�tҡ���{�~�[�w7�c�-�O,�ݬ;� =rR޳�q)N윅m���f�'b�*���)�6�Vhx��О��9s�G�����\(����Q�fi����,KN�d��㱸e�'U�������(��6�Ց���굸���6Mέ��Z���2�j�☎����4֑��T�~}S���Y1�r�bza�P�us��8@B78H��%��m� �t�~�p��\�XR���Di�[�b1
�|(œO��K����P���Ts�����t)o��E����9�z07*��'��^5���Wf9���J�E�kAc2A����@.6(J��[V��J����z�bN�g���U%�s��9�.�Z��mI���c�wH�`#d�K�;�?Y�뭫�y]j2n�ƴ��^����N���=�uņ�#�p<��2��w��=��
��1���1�8�>�cs8g�zt�Nm�����<��`��񴪺,-�D$lA��D
A�Z-V��qU˟�\3�-E�rr��(���1�3�#�
~��$w�%7��Z'!E��$��$���J��*��{_t;�x@b�@a4�����IP����b��)i	�@�˭�%�O�����%��V�]�ؚ=VNj˭�ߎ��</��({���I�W`kx���
7Y��̦:&4�-�>6<�>���4�t�Z-���)�U�E�J^,���]AxճG�f'�V�O#Q��+㼢������ڕ��D�V�UW��Ǿ��c��`���c+�**+�=.*NCg�ߍ�����򸊾�(a?_����ժo��g�ُkr'�ݫ	��V2�l�lL���r����Ϝ>7�X������v$�A�T�^_��Q���S��E�[`�g��.��L��8F����+��w���4�R26fDxv��_;~���LC���ճ�S�������2���2Ñ�P3&���~������Oy�@�������ޙA�|桢���/�E��9�Af���f�qA�;�Ȋ�	�n����v��e��ˁ�3�+��H����e��e��иM�qq�w��u[H1�F�����:�~"C�����#lV�^S��NH��ݶ|��XJ~��jc٪�Ė{-/�W��H�~�����Ag��ہY�Ёq�R�m�Qh��N�b.:OLRn��׍<�Q���<s�B�ٿ����M@�] �� ,��q;5�We\s��V:*W�6Q����G{�xͩ�ۏ��ZG5�"����Z�!g�8�!�H�y���	�f�;S��-#}9�h�ݜ'3�_��yX�b�1ֵ��cWH�����+���5ʷ�>n��K%h[c���4l����9F�m�&6��kUiW:o���yBsx��0���Y���4��[MT貰��<�m@�k. Ra�ʛ���[ߪC?|��.:��fj��Fy�Xk��~wU���b6�ف�$d8�L��QmL>�2Xc�f��%����ǅӁ�
v�>�������?WX��!F����Rׯ�vs���%	q�aţ��J;�T'�y[d,���ZBGzқ�w��׺��>18s�V�MZ��t(�tX$1�`��ǃ*3�~++hl7�B8����X�V�S!E=�t"�NT��N�10ƹd���o�a��$�1�FMKe�߯`�^�Yf���n���d��]�ޗM�s1a:�1U1_a��o�a�m&G��T�NCG�%͚\���7y �׽�KQ��@?�����)�-zX�����U�}������}�ɜ
G�1����Һ���9�|�I�n��~���s~���;��0�7װl)�E��$�����������`I��'L��P�Z�m���?Mi�}[/�-�]Azh��y�z�[�v�\R��v��ʪ�뗛�g{�a���.�O��	Q��U��l�l�pѝNY�p�D�+��9�Y86X�g��LdvӍ��̫t��ḯ.:�l�(�u���L	}�WGS؄�n��Ƞ�hm!��4snez~���K%�,f|c���L3o�=[&]ckr�*˒��3iM�9V�n�f�un�-�ɏ��v���v#����F>�P�^�	�իo���s{�ʯi�>šm�?1��h��kT�����b��"��S�����{�n�v�Rg�+��(#a!�)�a6��O��
��O���뮠�)������0�P*#�Y&�Ё�'�W�����i��s�β,"#�{Ɔ��1~1��� =+���(����w5���.j
�9�X�VR���+p.��O����h��B�ۘ	1ޓ��#�����^�\��n�ݡ�K��uL����]���Y�*���	;P1��*V�`PG,����0�>j�}��6{3��D@���u �|TX���X�:6ǹXǀ�~#����>NR9�ņC�*.+��cn�yo%��
�q`�� o	� ���E|$2�d���Z��~M�I�G@4xMc�p�[������q�b'j�:,.��l#�
�B��
A��K�&gp�
�l�D�Z�͠T�W�"���������F��á*�PZ'!X# ��$�
Ew�µ}7��E��;�N��]���u�N@b}�q��u�	�N0it���r���-�聆�+�dDx���M�߿%ߝ�)�Wd��D+B�
�m�^;n�Z�1N6b���Q��%�&�����Sԡ�]��	%"�cC�s^8�]ٔ�iQC���QC�Ⱦ4��\�e������Lwi��_R���,,*s�e\;���)1	��ʔ�m-��L��6�>�����W=^U?������A���u�'��,��ߢ�T����_�Y>��l��q���q��˼|��}����/
�?x��Io�Sk�ؑo���߲��/lz�{�}l�Z|����?zf�nm<��z��ʌ��"x���7ꩍ��!N'�Ɋ���>�Vw�WlC��*-���K��b��7�xf(��1!��G�*Cb���"�^n5�L{�zEo=�8'��ӕIӀ��^��{�Ɲ�l>&~�~lw����YW��p���rc�HB�%P��/��CE�:n����zo���R��� 9{qU9��g׾s�6�3dC��nx�R�P�vR�C�"���zS窓4��r擸�b�ϭ��s�M��b$��������Q�����~Yb�}�l�w��I��r��6T%W�F��v�����=�#ܽ'!���d��<>�P
�����[V��J��K�3 Iڣ5��o49SQ��w�ۗ����r���ٰ�#����#��;�@��==��q�u��w��N���"�����wC/�>C��l>y���b��f�ǵ���!c�*wO�2*O��ށзΈG��Y���r�wۇ�����H,�r��/]u���nW��\��w[�ow.�د�Jg+���=�mn�G�6�΋���\;��URݞ���y<��ˤ�4=� �?��%�w��ӐWP�8�HO#_I�.��Z�	酱�܌J/�N�Jv�z�s��
J����TB����
�} ��pR���@J�lg���{���R�x�@_��*oG�U��chgRG��S� m!#�iM���r_`�	g�/��c�G\o_{5i6"�4���|+g�[�%��"����|�!?j�'�*��v��\?,�z����m������SS�X݈U�����Bxnr�[�`���X^^�+�{�zd!��E}Yq_N]Pp)a8�����W^l����G��;���*�^ޑK��ն�=��U��0,�I̮�A�p�]{f%w���'e��A��&<T��z{��U�W�@a�ɨ�H½�9]כ^َ�t�W���+��d�6������Vt��Z�(x\u�jZ0������J/�"G{ǅ�:������2��+��ڰ�v�]�Q�`��ɱ��!�U�;N��;��f�)�u~��y�U���щ�ټ�FVv��R�Hظ�lau�M�Z�����V�OZ����k�;�r���(cܺSwC5ܷ�E��w����\N�k�ޕ�h/5	\�jw�5�7�W��TQ �&��O�"�����o�8�N�[s�b���g�T��4�H��j�VO���{:�����>��P�x�Cd�W�r�1Z�������	���������֪[��a�w�}�_�G}��������vU��th^�)G�o��޼t���o�#����F���9�R|߿�m�Y��O�ԥ{���ٵ
_��%u�7�������]V��-�,�z�u�k�l�]�ӆ��;�3]�)>^o����� �z�`�s��^�&<���ڳל7y���|���+�����A�\�a!��D�i��y��=�!J��s'�κx����Y���e����w��f��m��塤m������U�����_%�!h�]7_J�L��-���Z�t܈�����V�b�z����.�"�㴠E���Lhy�W�G'ª�KK�����[��������n����[�K,*ksmΙ��*�L���z	�Sܬӏ3��4+�L��[nVf+�t�.�N�N��2�����˴�q^Q�(���";�`���٭J�qV�x�PT�)l����vҷ�>��V�=�el��H�����Ϩ=L%��
���{c���=4��5Y+T���{�b��(̗�Mg;�NR����|�׿~���s�3��[5��69�h�\���>���B~�j�O��,?Xj�����I�Y���ٸ�"�{���J�������!��7��z��Sooc�w�%T��]�N$"��׽���W�n������n�P�A�*{1%
|f�(]��w����`��c����_b����,1�(>����uh��N���xA�K5���3j���o��ߜ�j��ʺ��&��cp�-o仨3L�=�T�ʺ����|k�v��}˼^��NP�Y�bh�".�a��1*l�l�Z�s��s�+-X+r��}�n��y��5��P��F���ۄծۡ��E�~� �ƹ7���D���*|y�9��l�F�6t�Ç�8p��
!휉^�(�:���S!oJ.J �bV�-F��/s�Z9�n�1�f{��#u�(�G��	�J���i��ҀX�w!\���P���\7Rmo�`�L_-;wX��@��s�}��6x{U��\P{).�"�9Gr�
!�-C�f^b��:���1Q%��2�@�-)1��"�`܅��'3���w{�>�+y�;s��C��{VF��O�����ݭ�!{�ئ3/���9;,�g$_wIA��P=\3����V����GO�:��vMX�S�rY[�^�����L[v��+���r̼Fl��B��V�K3���3�L�ו/-��C��cN��2�����F^�:�SKɲ�A�\b�̅�oR��5���w.l�.���%3���z��|�4��r���!�e�[�6�U�:�V�ɓ.q�[��s*)��4{��uM�c���ӆ-���xn�L�)�3+v���rKT�UttJz8(�����S�R��+;tb�OX�^��e9a�]6�r���K�B}}�-2�.��bYY8J�l4.����q�X�,�]�1_W�fSaeF�ԩN3j�-��z�P�ۿ'",����QЬ]��������d;�.e��6�@��[wO!��=Ks��D�~݌;9��-[F���֣�,���Ü�5F)�r|@B������:��x\�-W�C2�bt��J�л2E�Mv
�r�������R�5]��3�����Gx�$x-���A�d=Vэ�K�9��^�~Nb�^��H��p0=fq[{��ٓV���i��Ȇ����Dl֬��.��\��GFw'n��+]<�(BC�[یk��%Gt�{��Ve���i�R\{9���p��Q�b �S3_+ʈ�̛%��t�YF�u4Y�����
S18]���nݜ[�k�o`�s�T�/��ت[��fm�,�d�9���*34�=v�0%d�YO	����Z�)���\tDdso	3hի̂ ��U�|ZA�(�u%lH��"��t6C��-l����+���+[En���P�p��W��}I���)�;4S㎶gY2��b�h��,h�J��\���K��p��:N�s@���0��O���-�.�9>ܾ��ə5��r�S���ܕ��k��RYؠ�,k�9�����0�[cbfur{	9u��6�b�kV��K\�Kp��PXe����}��t��-h@�L=bc��¶��i�5u��f��Z��By5�=Q1g�b��|�����cA��J�,)�[�t1|��&T�Օ��b&K|Ak���^�o'Dq�­|��nv_Cϵ�'�U$6��JU�I;0���r<&����1)0a��w4���A.�)81vv7�uސ��9Ƕ�o`�+v'ǁ܊=$M|Tjߏ�������Ow����@ Q���4�a\��A� ۢ~ۄT{���M�$
';�n� �ňJQ"�c	r��I!�����/5�I�\����J�s�LX(i��RQP��M,#c
C ��5�t�9���$���`X4AA�h�2�˶�ݱ�5�cQ���h5&
$���zA1�wX���IQ����I$w�k��6��\���I)-��\P���!����4iM7�s]�ڽ6,Q�Lb4L2TT�u��.h���!˜���  "�����M����G�F��d�a8��]eKr>��j�l���S�#�$2��%��3�Nuc�4����`�~�x��Tw_{|��}�7����d{N��t��G�:ްG�����Y�wP�Z�X�{vU�������{_�8�I���yX����ԃ;����W���k�;�����xt����J���ի
��!�=jK���}�һ�3���%z��?�3=�O��m����E�4V�^���41Y=3{�+�Z���(=��[5y}���]�kV��s�z�u��I�7�@����C�ʭ�#9�s)XY]ySt��k�uޟy���w!g�R������ścé�?����v_u����ID��������\!V��&����ؗ޵��4U\0��C�%�3�Ă������Cvjqn��˨qA�e��I���Ǯ�}����B�b�\�r;��Q��\pRxm^�/y��|���������Wz2�����v�.��@��EN]�-4NF��Mא��O��q�15���y�3�u\�� �xg.9�})ˊ��x�#�h56�u�Fw�Ӟx����wG�N�N��N-59��A��3t7W�WR@#r�:��[��w���&p9-�-�,)��;:m&Ӊp��_Ļ��-/�2J��� �b�,fo�'�����:�}��;�7��!VU�Ëܻ�==�nzC�b�ǡ����,�c���=4�Z����C����w�\p����I�B֝��?v�ȁ� @{'��N�w=i_��и�������;R�zJ[�Sb������@�7�޿�z���q&c���a�#En�;���_�w˞��]K����z��=�_�9x�ǫ�nף�5���ëA��a�s���_ж�Ƨ^H���|���^>W υ�����Y��Ѱ��y&Vq�n�y����.�/�x$~��b�F٥�>4����ܬͱ�/��s�t��W;�o�w}��45$) ���y���ΥB�g{66ѭ��E�M��?o�>4�b&@c�=��u�~Λ���J���(�*��\ئ3�����t�yJ#��n�l�ڂ0t��d��}�/��{F�M����m]�$��k]gWqTD��'K �[��,�=:�Y�}��2�{�;�+*�|��aJ���?j��g:��"���]b����e4y�;�7c�ت�z�;汆;9f�>� ��Hɕ�&��
l�õ��sB�+0%@-���G���yZE
���#�r�J�:�ǱJS�OW��z�kb���*˯����,���T��a�z7e��&g�.�u��b};_o ���:╲����z�ʲ�^C8���_Fέ2�w�g<�Z%�Oh��P���#�߹�W�n���v�g�\�N�/^z)V�ОY�N��&$,�,eII��H�J��mg]c�ڨ��q}�eǮ�/|ǎ����ί�e�CY��H-���8'��C���G� ���g�%(ά�����۫�8�P���b��@�br}>����R5�O�Y#��QdO�;#���__�ٱ��<��Cϣh��tt��0���g��#�s�3�G[��){L��[c7���ˍ��S�o�z�@�'�=!��='�]V�缔_�l�T@4��U*�ǝ-)e�˛���st��t=[p7f��¾��wE��\s��ʄ�=�H|�T-������_�sJ�>W<~ϩ���ql�pWoU��7'�N���lk�{�͚�=>�U��(槧�GSL�THOl�˔#�8D��oQ���TѼfug^��a�tH����#��[w�\�>R�9v8��p\em���&�00��R�x�:�#�Ov��Ϻ�v�r��e�����zk��}�>�'�5�H+�W��=�Gw]]Oz�3.���T篺{������8bՂ�0Gx%?x�O���:�#*G�U���n�7�����B��u�.�Z-W�6W�[
d.�U�2�������3��y�OuOy���{�K����ņ��{�}3������~j�x��U�MI���%��}ˮ��k>�O�v���¯��+���Y�u���-������z�6��^U���!c��n�N�>j���>A�~��+[큽##j3S�,;�jWH�����na����&xK�5~��8��m?}�<zP�c}�;S��bod�}���~[�P�?
�,.e�-����׻��@'���	2�Z�a�N�i�+���:�at;ޑA�Ala���R�#����5)��c�?�M�&ێ�A>CgpE�U����o�}&�p/��H6�YJ��d�`M�y�����v�پ<�8���b���ڠ���n�{�i�kړ�]xu���4��Z��c
O��%��L\�Ք:��wn)���*�&]k{;�9u����&Ŭ��WM��y�6�9Nk6mǕ�������j���9��
g�����3�T����,�j��������v��y��[�r�ݠ��E��y*�u��swb|jݵi�P[������e�7�W{=�MFȀ�����J��1v]�����)5'�8Wk�T���q9�ft*����1�ן���|C� i�����~�n�-���vO���w�}�E�u��ը.��m���;�h�(o@�r{֋���#ٙ#=�r��Ͷ��n�>�����ڼ��^��<��I�&�tg?OF�[WQ�S���xzE�s��R����w��j«�#���IWyٮ6�;<6ER2�؟g����Ӟ�4�!_&خj'�~���-�l��̾1��v��)�h	c-�����=�9��bf�{�N�n��/�e�c�j�}�G~��,�A͝1V;����'ޛg�U���|7Z|���.�����4H�wk�Uy'��2��ɵ)̸~�n�_l��*N���m�` �T�p�����J�l�l�:��.�G����T��W�uɒ�Sʴ�i�t���ei��KG:w@uJ�$[��;ۡmoo�7ky�|Ed���wu-�P벦jY���U�,Q��G'Z�]���{=���,�a�O
|٪�Y��پ��DXY�2�y}KG�cy�?:e�yne]YU�����p��hbs_����u}����x:��Y��?r���?7rӻٔ>��W�����B�qJ��V;���/��!7��j��dj���g>}J��vz�F25+���}]y��ى��F/� !��on����3#�I>t�b8���Z����3���^�~J-�w����b���O��땿bq"��>|�F�A��[�[��Y9ۙm�M��z�j�ln#���p�|rS���B0�{��AW�o!?`Yr'#�(�;��o����#��﷬��Ȫ���/p���;���	�Bz�7��o�+�u�t2�l���Pw����Yd��|���F�BT/Vj�`����ڝzҞ[y�#k�����o�2ס��:'.�����v��ˍ�u��a�����:�����W�+$Lz}[{�+��t���u ΀�`�hU�[��P���I�bs��9�AKv���R�y�\��:���m����ſ�!�����3g(Sє�_�9�Ozc��|U���sqM]ѝ�s���P�B�f����ҵ!ޠ��h���S$��x�Z�.���������#��^+��w�����45%Z�D�p���gߞ\�йC���ϒ����n�Ǆ��W>�{�XKa����=�Z��[�"P���dk�Z�ͷC�ˡ��A~����f�N���Lw#��{�m������P�X��?G�?�V�.�5��PS՞�^��N��w�i���n��/j>;����a�Ɇ��oމgǷ�;�7�ԟ���_D�TO����=���/wK	�R���1f_5�^�h���γr.�/}[���a��!X$��4p���-�ep�.z����<���؛�d��������e��d!�����රȕ��oY�܍�r�O^�U�Ԭi�寻���Wl�UÅ/��F���JiC{̂~�2�@ڮ��B�?��ڊr�f#kt�2�v��]~*�S׳��(�
��l��wQ��d讳@��w�E����
�e��L��E`u�ufIb��S�[�S��E,�" �K\}�X9�S��J����/e*�&���A�8��y����|ӛ��� ���.�S�U�" @a�٫�:-v\׷E�t^#��O]u�3�W���ڔ�[�F�g�ڇhH�~���n��D���.��޹�j�)e�������&�G������X��0bj��uY��d�@`p�5$6�{����I��z�Ϻ��zc��$�<�v���}���-��X���}~�Gy���z��&�A�b���Ӓ��x��ڭ�o�~�����v�C��I?
��.��6�y��[jo�w�N{EtO��Wވ�V6]j����Be.����S�
eWO�UzN�h�V��
�Uߠ���b�y�Z��'�}0uz>�{8z��Fl9���o���/|�y}cf>�U���5kaZ��x�7�E��(�WF}Q�1�>�X'�;��
~�#���{�>�=S�����	c��O���lE˺��ML���]��:�5vQw����؟g��.r>a����uKRN��峒YYS�e�o�� é����n<���3�Ϧ!�c���"�m�+�V:��lE�����x�����«.�aO DT���+�@$�hf�M�9�.7'+��������?W��{@�_����<����}U����{]c���^o��#�_�FY�;{�~�L��xal!|���W�F�](���Y��e���M�����o���z��|[FB���Y	�A^����?nt��/|�8�o#�R|�Ί�����,���-���C7;��bF�u��!��Z�W֩�r�/�Z�������Q����|f먞H�up(@�87��Au	�R���'�c�V�	�gf��(W�j�r��=ٽ���]��3��^��OD�X���ښ�n>�����f����7�e�T�!�����ףܧ�v����1�ntq�}K ����k}�7�W����no�:���DS^��9��|/������_&��A��}9]Ӵ7�mXX!HG�}��ǩ���*�9]��9^|S����]8Do����u�&' �7r���2,%k�<��7�;6GЕ��]���s��=%����Ey�(��Q�1;y�u1�"�Y"M_A��Ab�u$r��1[xh���Z�gw�� U��#�8��G$]�{i�^S:	U�ܥ��ߪ�O�k%�%IP�+)�HW��H��}_XV�s;��{�|�m{ې�W�*���<�p��b�\����5�B���{<ኻ�����p�_O1�'1�������$&��g�j�n)D�_�N����(S�=�!y'�{f�jWr�~����ms��~�\N���sޡ���8�h*�ｼ���O瘩��P�c��*���,�a��������*�U�Nk;3�����I^�ש�oΝ�}�[%�N��W��M_�R
�?~j-�&y	�s=\�m��7��_g.����\��9&�KN��y��9S��g1������R��Ǩ	<�_&��.�ڂ���rs0�kԉ��<�=���� r{پ��t�����o_bc8=ԓ���w�h��;w��/ʳz�����q�\Ã�u��mlɏV�i���:d��f͛8l���;\���Q�1դ�m�V���+����$���k�dnng#��y|Փ�5���"vaKH�$�]7�:y�mm��{W0)�$�K\����a��ͅ�H�xE�3�ҥٗp����=�8�񚢺;zv4�nD��Y�_A�&*�b��&A��:��PHO{���T�>��ok ���tQ�d�Fa�+S�N��]<ݢ�՚sf^�uy`��[�GPJ����,&b:�b ƛE��v��Y��m�tF2_n�Uw�Z�+uy7'��|g���3�6Xq��'<�o|ؒ�1;����S�&qWƏ��q�%ʚ%��B�܉e����j�R5J�����;��J+���[u5E�x1�Z���Ff��Y�n�7�_nט�E��w�]��� ��*��SksT�'�X�m�M=˺{2����b��K��CT.���w܄�U���dR���[��ka�#t#D�C�����Օ}��L�H#-���̙r@^%��#�3�=|<��Oٜ˷x4V`s~]sq� 3v�Yx�TŹкL��8f8>u���¹;k �j�����0�e]KB�s\�8�Z��K���βWho�����xn#83r������3&�3��uf*To��u6�sI�+�����xc��g;�R=��"�)G��)�1>����(�[��a���8�J�̢�_
 �V���Ã��{f��I��n����WT��g	�d��$�$��tQ̵��,RӈB��=��xQ�n� �Q�t�!�s40�g]�p��"������+2:�@��pĺ�p�u��}�5��u�Ns��c����A�8k�+)�;"_����;4v�J��Yl9�ݰ;�%��	��1:Q�:�lYe����#Э�
���V�����|7(��e)d�ͥ\�1�׋lY��Gfj�~[�5��x�,�5�n�x�Z��J۴DƔzN���E��-G�f7!�q>6�m^��;RY����"���/�����-�۸#�-<w���+<�?
�X�ۓ��X��1V�]l�oRB-�ۈ�c������j��I�u~���u�r��]1p浧,K��l�.�`�>��*�+77���ڙ���fսJu��g�kT�cVE�+��E�]�W4'�GL�Q����ҭ�&.��9�Z��%T��`u��D�W�lK{L�]ّMejSe��^�7Q��&[�q�� dr���F���*Zf��[��Uג[�� �0���� ol[����o�s}�l���-=�����&���L�	a��Yg���N���;t�:4�m��	[SY-&��(�b�A���.�C�^uM=3έ��>8�d	ʷ{[2<E=Z����I��í�ǝqWR�Λ��T]����K��4��iu�u�PU3E����Q[�J^��M��j�]@ �MGܩ�<:1�����rN.�{y�v)ҷH�I\Ҏ�uu�:R�r,�x�Wh;���;�������_ n�4A��hP��	7Ii�~m�O�z�J��0i4�#}wQc�a�p�¢��T��1c#61�@�Ri.��srou�I����hѩ5;Dm5!]� ~�?])0���?��k�v�ӻ��r@��[�����{yK������q�ޚ*%L(DQ4�����m�v�d1g:71�]�u�ѢKʹQ��uм�͌IQS��ow�wr �ݹ�g:�7.�7{��W�幡�E�^sL�\�s����I\��9s���lr�(�1�;����\5���K�:�3#r�bƴ�bז�k$9��F�	 �$JEو	1�8�KǼ�UrW�k�X|��Үᤆ�B����q��J49*@��c�0�G*p���4�M�{�����:1������a`&��jb�}�;�q��[z�ҧ���?z4oӰW�[>8��)�ژ���ݏl�t1�H{u�]�ܸ�o�k�[���7��lo}��v���&p����ëA�����twS�\��M+��ꡔ����o^���w3#����W�=���	��f�{�Oj;�/S�ZS���T���~Q����N�l��t"p�y�g����}՚���k�"Dt+!�{쯡�}W��q�ޗ�/_�X�4������[�ѳ�v)Kw�t:Į�$w��$�x���J����^h������m�ߩ(��A��nD�`CG+�u���|�1ϡ��4V���l73�g����.0g�M�u����W��1_v1�����{q�ˇ?m\�S)�qĩ~.p�R�k�~��C�?S�;};[�?X�à�z�K|�w��ϣ��9��[�5qW�Sd�On���e��E�U.�k�[����׋�Y��b��*�)o3]����qD��"���7]==L_#�H��+l���^ ��8gL�9�;�ڴgK��!�FO�1��pv�]�p�|�4�z�;W@v)���9~�P�k?g]d���/kK	�:i7,������	4�g�E���^̯����	�bKO4pќ�imE���Q�V*o�Y�q�޻A'n�iݝ��/V�C$�$)�w�pY��y�Jf����:����k7���cMur�ֻ���`��Lo�E��Y^�3���d��u]�S{��|ۛ��ϡ쁏c��N����;�.�ٓ��3u����P�G�2�w�����u|��ڔ����3�0.Nߔ_�P�[<#��w]i��_O�I\�Nֻ�V���k����� ]&oy�,�q{w������m��޸��>C��7��Ow�f�v
O�ו�	!��F�K���[=s��w���n�:�w}[�|���5�a�g-w��;�P7:rr#1����B7������d��B�b�� �89�n��gz���5oc�K=&�WA��v*�G��su�̛ȵ��O�o�ȇ4�x�Mb����[�޺��"l�1���o�mk���4r��ϻU�_�̢�	1�+��Ȃbv wej�8.��s�ݱ�Dif�[�Jă+6��}��N*�N��T�{{cED��z#{c���﹃�N,��<(oF�	tHZ-P�>�,)�#<]WC��v��^��gz�^ygۯ=�O�$�!v���㾜)c�k�oJ��hB�����b����yz���1!�Oo����bL�E�Bv��g.xZ��\��rn��|�@������^��W���[��cU�ܼ�yo����!�����(=�4](,<��T��~~Ư���Ԍs*��m�&���)h����6��%�V��v��4one�>`�\��
55��js�x*��Zo����r�|}����{�P~G��T�g��\9��8�m��Gb�=���m�J�O�}Z.��=�����/(��=S,z���s�k�ͪn���5���u�~k3у9�A޼���܁�ꯐ1`Y����j��u���b|h[�����_+G���-������:W<l�pC�[��l/@k��$���(Og{ٙ�x-�wO!�T����ecm�0C֊J�rf]�Gy��h����
���K����v��K9���x8���@Ҿ�"(�s�F�]M�46�5��z=���$|��W�~�W��m�w {�e=�P��wǫv;���>���quuU-���}���=�/hu�#����L�����{E]��'~�[�]A84��1IO��5#���Z�C�:F�GAC{}�{S�]?d��xuh9��>~M������W���K�X���Y���~����@��M��L~yZ=��������W�+=S�-��_����/�WD�w�����e���a�����&]�w<�w��Z�w��6����ה�n��ks��}�.x��p�4�)6�	�����y!71L���~+::3�����[����r�ƹC�J��W��v�)���B8F�S|
u��-y�ϖ��瘩��V{e�#ja��u�8�:'�kc/��f{�}��{�T��k�o�-�~t�K�P[�_Tp����+žc����}-��X9�f���7e"��>��@�>u��\s��2�#ɕ���D�FP��O9�_��ϯ�X(^*x�e�U��t�pgvPu�8��3ݗF���e��m�������4Z���գJ}���%��qv7[3����Ԧ����(�E+w�M�S:�Js�S���[ԟy
�}����}rMܴ��>��ɾ�7;}�w�}C=Hy!�=BJu��BA���rMe;��*��S;�FbTd`��Y����w�}����!�^l��O|+x:�X�_��I���l��
>%5�zrVv�^�[�Ĉ���0,�"8?T�_{�Pr����K�=��tQ���?���[ֵ�m'�����Gll���`Dl�xn�Y��V<ڑ��}»�g��v�X�/]�M��5�-�X���=�,i�����D�$F��z�Z����9��K���=֯�M�iT���UC+�Ϋ�D���-m�/g|�	<������޵e=��,��7䧯Ѿ�wQ��n�̬ݩ(Eθ?1��Q�����5����Ի�$t"�u�מ�]}���R�E�}�,A�$�9@��hnA�b�;��F���ݸ��r]�N���ݝ���&����o���ܹ���[�vv)��'YG�Y��h=��n[B=�0�L�ԉ>����C$l�y�}Y�1e��+/"HF��`Sn�<�#}Ј6���`WwL��<-=�ɽ\ҷ[��w��V�8���tk�\�R��n��\�L/j؞�Cf�x���!����q<��W�����{n,��[�=�ں�({y�y�9������Y�z�>�x���	���	z��^�+�j��ֳ�}A'¾�_0�?b�[��YpÌ��{ۛF�w]g�_R�������V)��ϧky��t�z�K|��m�X����5=ݙ�mY�v��_	���{_,'|��O�5⫣'3��{TϷo�6���U}�̭x]^D�_P�Zv3G|$g4Yۣs���\{�f&\�i������h�N���;��eP�d!��lI���n��NU�ɺ�ͣ2���k������|���Z�d}بG�dh�c*�g���T2x�gx�u�f��6����E�nt���HǱ���;:|����l��%"g��·���=^�sk�箺�U��V�Sa<��ψ�z՗��?�io♈bn�:ߵ�.�q[5Ir��ͳ;0WT̶�:�N>=JQ���>��{��,�j�����O��b����K����e�k{wu��:Xr�f9-j�2�l�b�M��$���bYW�d�5��X����Ro�z��{��~��߾�йh��v'�����k��{�=�[�>U˒5s^]ͮ��W ���=�ޟ�MT�{5S�R}Cj�n�J�������\�î�pm}�#�w��������;A��N�M�t��8Μ�)Vm��J��v�����X�#���S���Q/�f�Ѿ��G����}8�,��t�Y�5O
�z5W�tO�E��#�Pmf������|�������̟��Go9f��!45$)4%v��fZ�O?d��.�۳�X��xs�Uyv=��z�WK�0�?`΁�������;�'=ݸz� _uA���]͙��꜠��B+�������_�������+�s�]�K�E�����🟱���������؊�����żBK�������b�.��������_���g�J��2�S����R�f�ݼx�����i��hpy�mᱹ�!�^��>��)��
=������1�v���w:�$n-�R,���^n��7R{��R���e'����.!�Y�bEXt^�.������y(��}E:���Zo>��km���u�����/r����n؜�]�����Gu)��3�ؤ{���qm��֭?*��c��ֳ-��#�,�? ��!��.�t����C�����KO]>YӸ�W���w������]s�0(�����T�}���'��I��&f�X�F�9ۙk�%�^��{��7��^���N�^������~w{~A�~6NH�~����=�Y{���Cz`i�|�ki�;�U��=�J�W��<NՂ�>כ˺�}+lm���}���E�=3�}.�7�=�Gμ	@�6;0�5`y6��}Y`k���t�ybV!I�f6�þ�{c:�a�NA��s��^����T�%S���i����'y�3�Ƽ�7���Ǯ�?�0���*�x�ߵwp�^�L�䄏���ؼs�a6׌e=ϑ��̲��-���#87$jE�bb��|��Ŝ��]�]�r�fy����C�r�L� �d�Ԓx�/���#:Γm���_<�S8#L�\����8]35������y3�����V��3X��_-�������B#�S�T�$*%�Ź�í�����~��t\�4]�#_1�-�� ^\?&�_��'o�ק������ɞ�!_j���]6dl���?0ܜ�CO�~o+�<��4Or9�ٞ4���|��a��*���ث*�ًb�U˫�;��=uU�jz��|�j��S#�����,T�J�=��ue%X�ڎUپ����ȡچ�~�'�������ŇCz__ܓe�Z�?@��P}.�X7=�w����)��C6Ku��B���So2��w�kQ]�^�+3׽r�{]���e��\4�ռA�X�mL����ј��׵���o�ϣ�V=���}
6~,���}��}�f��N+ށw�zCfc6x�S��]��U�k�8W�^��pG��Tv�|��'s�<N��?z�w�*��;o��w��-y��ic�W ��>όb~�E1~�����yS5̮��5�jCʥ_[�Cq�D4|qv�v�vN�P����������YO�_�ۇ���B�R�܀��`��E=rJڊ�[� ��Qp����1ii�[�֎O�ڊ�`��Y;�%�]�	NWp*zzo�H}�U��[�����!���kx��|{�^���i\��Mr��tS��՛:%���忂��]})�a�#�\�o�f��=�����:�T�X�%��a�3�\�`�B6~�G`0�n,�~��v����.	&�w��3�\���/PJz�Z1u���e⿧|�q���~�
�x)[��,sK��Z�;-6z���`�3mdk��#��R���=���;Y����&���G֟�梲��ɇcs{�o�>�syz7*�0X���)��#-�=���aP�_ͭ�����<2f�M��N���\.͸�\`{�2��/7O�w�y�ra�y=���Օ�"�%����w{�c��������T����º'����tK�XN�=���������~���X��W+��^��e��$*�t$��f�"4�s&O><lٳf�6t�m�����5/6��%¾�����]����� �t�	n�*��]�m��/'=���8V8~����'%ÅF��!�O� n�+j��%Yb�[5k������hm�A���21B��y��	j���YKz	U|��zd�AR�g�qJɩ�/�Y�rz)^�sP�6�|{�/",2��V�9ͦ��r���:���Uױ#�I�U�d|��tRGM٧�e�[Xk���ړ������1)���Y�e�$[oR�di׫2�_u����P��Vr_7[,�[�X����>�v��+���27r�B��3�S������t��5�q���!~�t$�{�,�,�1O:��Uq=�Ѷ����Sfȸbx���7WH��]�c��[��Y�z2�X�Ȭ������N�[$lf���I)YM.�[�+���jnQvV���/!�]�1N�L�k͋' d�ʅ��Ϥ���Y�R�T�)�!�Nl˜]��x�;�C׌m�t=Lb��֎a��#'7�w�b��<�G,�!eك7R\x��ҡ���i떹��������=C_K�н=���o��հ7�4e�vvl���^�Wu�wQ�:� ����:2b䯴VeHn�q�a	ȊY���r-{R|��A���I	�QvF��s���A-�ܺ�K0ȝ�4T�mrI�9v)k4oT�@��@%i�\ȱ�g�s��ֻ*
̏���S�N����fi�0M/v�n-5��8\q�Z
@�ۡ�}ћk4�u!��gpn����/oc�N�pё� S˅�c��^
�ՂCy�x�~�.x��ݮ{[:�6!��V��Kkʸu�+YM�Ѯ��/��#x�����7�e]7��a.��ʵ�ʗ��_!�����]RH�O
�(c�=�l�F��1�	6�{��u�1^�c]7:[8L�a�}Z�M@������!9�+p�x�Q3dhr�����;�o�8�~���Vՠ�8>z�"A���)�v�۶N%�`#@
�#����jE��7��D�۩�<�(fqwD[�m�S�x���[��H>n�NO��\ʕ5������R�i�+6�y+-��0�vH�s7������c�g�<��ʰU�t�kL,Q����7R���T�8s�E��ܐ2
�Ni�2ģ�%��n���P��D��
>��Q��i��!M;�]�� �9V87b�{C�L��wM�����ս���K@K��M��m�n������^V�`͏q#��̝Xn���޼�k�����NC�H��ۍ���]Ñ�FʸO,�tШL�׆0L=׆I�b�,qxL޸�U��&
͙<�GD����E�*db����'���y�[1^�<��.�,�������r�Go��ұ:7.ݻ�VF��Ѻ|�:��J�����@��J!Z7�9�ԣ��1�Ļ��p�pwg�Z� �_^�w]��JRf�ƭ4���u���.��.��� ���
�>���L����b梱$�����D���L�W;�����56KW69�r�%Ú��.��6v]�u��cBMݺss�#t�ó����r�W��dѮl�(���+��gut�����77+��מ�]9�r���.�k��[�����;�r���nt��v�ݹr�ţ^r"��r�:�)6��u�\��]�p�k�r��'{�ׁb�^3p۽�r󖓖��u�Fuۗ;��S���v��d�.ݸ�.!����r�n�sn����t����n���sni*�]��י9v�E�˻t۹�\���N;�����!�˧\�#D`�W˹˜�r�%�r���G,N����t�r����:�s���ӥˑTj��� �C��d�&��Lu\��Z��cղ�m^cx��t2��j��Y�ugw�'Vͬb­��Kz4�kwWvN'1.���Uȝ�NT����{�gM.���6��ܟ�}�|�1���)���x�v�ni�"燽����:�?����M�_+�]\����~���~�x�Ǐ
�f��Zb��%���!���:�t��q��M������q�W��/D�5�E/�]1(�lp׳��箺�s��zj�jm>��s�_�%���^��2��k��t�;1�0H�\��k�+RQ
+˛���1Wu�Z�і����ɽ��_�������'���������op��H�]�����r��#}�����U�@-���#����@A��y�-W������U�h}�<�_t��C9.�w~��|�v�Jz��U�!OL�tR�s<��ueT\5{xzz�`��S�s��Ӌ:�O�թtHE�p�c�0M�]&
X��d=���̓ο%���_Fյ�.�=�M}�!@Rh.�?��Z��f�!���2�F"R���=�{j�8CjW��XRTv���_#n(�rn�lq�ۣ	�mfs���=�R^�����gxdk u�m�s��wB8%����b�Ӹq�6���s�PCr�?��.l�(���v��Ih���=xAh���FU���꒎��^)�
g�-O�1������yz���%�L(�os�����؇�{�C�	�����r+��_�/��+��E����_�^{�1K��n�U�ެAn�@,t��Bۣ%/(,<���xa�3^a���<�zgego������ڠ�R+]j�z�U�����4���M�������Uq�'�^�����Km�2ն�����u���O�?O�_�yi݋�]����c0N�U��ؤt��"8��\>?{���p�Y�����ysK=W�y�3Ao�N���^�3#qn�x>�<�Ӵ��@�RS�j�������M��p}�_T��9��r������״�׽%-�+��_-��9�~�G����k������)�g�M��Ƿy���ys�ܦ_��Y{C��o�7����,/�!J6s�9[���>]�G1��"�Q��v`T���B���؅�B�����.�ky��<�9v�{����9S��̘���m�V	�J�mw
yYVo&V��mԚg;�m��}��7kNq����A鏍d(Ԛ�7��8']]����è]^�ڿ'n�/[�{aou�w���qӿ�X�~�Zvsݚ?�{$ܜ�ʿ>~M����v5�W����[~X֍�����{��E�m��FAA8>�ϧНxzo_+�HRC�#�"m�NS�>�lmFvgq]b�:�^���.�ϱ}�7�7����Pq8�[{�X}�7�V3_9(�B�t4���ac[y;y}u�|��k}�hH̍;�r��O�}�|=ڢ���;0E�����XY���2�M�S�/�t���o��y��ȼ�xG�7U����w��f~��mf�G�)x�B�?g����2=�?jm���ܾ���-R���ń�v��/���U��b�yޗ�%�"��P�}C�����u��fa�-����b�{s�|}�C���Khz���}��
|�Kn>ϖ!t��֯Q�I	]���@������]�&��kڱ�urQ��*vt1��Գm����7is_)u =�gb�����p�ss�#�Y�Ԗ6t�+��'o5�f���a����XftV�a�G}��.�g���٣�~wW՛Í����I._���e�*~�[��؃�XF�՝��]�Ք��r:��n�B��� �m<��@ٛ���9Bxq�ׇ������(q�i��U~|�g�{]����g(�OMj��iWϑ�Q��ف�J�7��'L�oEyﳬD�}��۝��=�����{�~��wB�ԮwS�ʌ��$�Q��K/L!B�`' ���W|�U:)[֟��CJ�Չ�^��Y��-S+;v�b�n3����	!�R�T'c}C7��M��{�p[���޺�Os/&��wt���_)Ŷ3�F�E�������O���j:�Z��۩�wcth�����ƺv��${�-��A	�12���A�����nc�gy����,Z�Ч~��	����j�͞�� ��=�~����]>��v�+�r�>������Пo.�j�_��͕��5���""l����`��!����i�6_�}�F̛��q͈�7Y.��NY|��r�2̰����te.���&w�_P)�/-s�^���3�2�v��t.V��!'Z��	��6�M��L�;��p����f����������ε��J��Nję�մ�*W�O������͎��Xն�/�u+ɛ������׹���������J�?7O�ky�����ޖW��^yT�u�}�ϻc�f�C�ם��*�0=���\d=�`�K=	mtM��-i{xKa����;������^B���̡t�����,:Q1I��{�i�����
��i䯌����Ӯ=��^������	��z(/����/�W�z��x5Ay�����i��9k��v*�����!�����!_���U��BE�%��xw����f@�m����<���=���2t+���h��fߛ��<�� ����zz���T/��M�t��K/*n'Ƿ�����wf=|T@��Ƿ��`��g�-)e�ɼ]��-��]q�u�Uv�JwT��t=Cn�@���Bz>!5B{�w�͠�7�.c�7�?Gw\��p�s�������e6�t�%7��n���^D�4M�*���N�-�Yڸ�~8G�l��y:��E���W7&��#�?g<� �B<nfu�х�9��-ab�^�Ƀ�^��C����4E��n�Z��Y�v�|6�`��9��_���Z�s��Wu�6��w�o���6iCF�����
uϩ��>����k��m�Jz��U�!H�#w�fz'���4�����Ѣ!B�|q�%�p��uS�j��$-�&r)B�r���F�^�j���2ΐe�;x�}��؄�jHRhY�9����]=�վ�Q\���W�#���RcWUy~���^����i��x�!�y�,V{��}(Ӓ��[�����0*��r�u�b鋊�oT>��b8v������c������������c?gm/�ni#552MX���쾥y��]�<��|�R�Z����U�����H������N{��7����/xH�{��|��6�.UmR�z1KSPfz��Z'�l?�u�rh?IleN���^���m'�u-��m�wa�7u6]}����. �il�,�)��ɏ{��wA����Frqdd�d8�!�]��v�/{K�ٻ��4{�@�LT�%���c��^��0����5n�m�(�r��Ǵ�X��� ���M̀Wt���4��tY�>f�݌���R�� ԍO}|a��G亿W�R[�C�g*w��2-Sg��� ��Vz��{�a���2��-��]]���~�x>�<�}����9,\B2}{ꋊ���8=�G�����o�mXO��[�Ә������������m����l�]�3����7���41�)�)�����Z��?0��܇G�羨��3��B�B�S]�s���~�˺�;��=��_��������3�=�D�ު5��=�} �v<ԟ��?��f�~�~U*V=/L�u�ǧ��Nl�3��#���u�>�����_+�Ln�5/�<X�>��I�Pn%Z�k��t�a�˵b}������;�K��.�_��q^b.�ީ������h��=y�XS?1�A��{��ז�܉��Ҏ�uwT�c�d��blw��k�5w��/����Wv|>���w�v~�n��~�})�p���UO��������;P�+]</7CƁa�0����َ����3�՞�]��"�:�Ƕ�B�v8��8F��E,ƱD68�J�}3�E&�/]wb���ҧ/�I�}Hv��q<iu�� [�wV�u�:����U=~5���Ŭ:y�������+���;U��;�J�uB8��^��>���� �Si��N���X��D�ߌ�{)jPj�v����n�YoԽb[/��g>�Ň_r���AŁ��Vs'?=j{1��;��Y�M߂�f�U�;Cޒ�_&��KC�/��˿<l�n̙[��i�kiP�0,��}e��!rOo���5��>���Yw9�S3���@t��\�v���u���v����FȀ~�1w'ʤ�s�~l�Jl-�ǫ��6ֱ唯�OO��k m*��j���Ыh�ы��U�UL�|�M߻C.t�x�����ɣo�y{�c�𴇴�����
�f{��Ptb�	�z�k]�S��kS~O���牫���r�q3��t�=����o�t��H�T'c}_f��)���N	m��g��=���+��F��D�x؟>�x_
�[�HJ���C;R�֫�������	tџMݷ5j�m�w85m6������Y��'��Y����� mǻ��yZ�z�{��3��t�:��͠䗭�s�"^3��R�.�tz�\��Lm�1�)�݀��𣣭q�6My�=��r~ߍ������j�z, ԝ�S�~����DMG~�Z{�{���;G�$;��S��T:�0]I��{QW^���ާd){2J�!E��n���>�B& ��
~��=�kM�LS�ޝ���{�/i���*��Y�X;o-	��䟘���`8�<�����/�Ŏ�8����Ig��دW�d�+�9�b�R���\���}��M�ea�����0������ݷ�d��t�I���O�؟N� �z"�z��VVNv�~��Ovz���5ٞʲ���4,Oe	\%���]f.�av�[ܬ��T�nY{+�����DHN�~��Et�{3Ӻ;���5��i���IW�[W�W$�pm;�� vYt5K����XY�jW�����v���F��G!�z�#�So8�W���k��v'����P����)��kR�n
���V+�o�-���sPK�Y6�)fXb�[wE�G�c���D󔕣gc���ZY��z�Ъ�����L�����.�"�N���J�^�d�����>U�X�w�.W=�U��2%�ڇ%�qF�*�����H��YQ�3l���~�֊������:�t��|/�sc��x!�{oe(�VEb��W_�o���6���?/��>�3�Umd�7��kg����Wu�����G�r�k�K\��x�F��Ƕ`>���Bv��T��z� :󛪩���Ww���-�V�zlRr���m�"=���&��
��kld��e��'��B�_Y��^o>�]Է�X���F�̸��{.���=�r}��J��~��[Y�kቮߑ�|�[T�u��������R���7@�x�O�b�����N$��F,�=����A�{Q$�t����UE�vح]q�:a|3���k߷T��!5���̕BK���ٳ�
��x��{�����{��F�cfyz����yy| ���u�Ձ�^�Hin�Ig�>��E���#h�|�?_���y?Ř���  ����k[ko������}[Z�[?��ׯ]������~6�]e�el�lͶelͶel�ٚٛYe�elͶf�elͬʩ�S6�+e���ٕ�+f[f[fV���ڦV�5�6�5�+fm�+fUL�̪�[,��[2�f�f�2�f�e�elͬ��f�e�elʩ��*�V̭���*�[fkfm�6�*�U��]��6�-e��*��-��Y��5fV�ՙk3Vdʳ-fj�ՙ���2��Y��*�5fZ̭��3Vf�f�f�ͫ~{{�o���Z����fW�m�ݕUL֪�m���U3mU3[U2��o�_��[U3kV���vmZ�kmS+Z�m�S6�S-��Z��Z���Mꪦj���ڪ�-�ٛUS6�l�US5�ٛm�f�m�����lͶ�2�m��U3m�̭���m�-UL�m�}{���ٕUL�m�-�ٛm�f�TͶ�3m�ʩ��r��f�3[3m������̪���������f�2�el�ٕS+fV̭����ճ5�+fV̭�U2�e�elʫ����5~>������նڱ����U�[jG�p������������C���������������S�C7���|W�����I$�O�����!� �5��_���m��U���[�5��f��-~�O����?i��I$�I�?��`}���s.B 7_�������� � ?>��/�DH m���T���V�UT��m��m��U+-UK5�٥��Y��m5UJ���+6�����f�UU-KUST��f���eUR��l�m���m�m�ŭ�����������N���_�v�ݶֶ��ֶ�U�*��v�������G����@@����   K�0_��p���`E�?d� �>��e�H����I$�	>�E�:��7��_m���o��m������������V���W�g�UU�ߚ�1�Y�A?�P0p1�@��$��\J<~��}U���m���������n�m����VB@
�k~�O�} ��>�?��"?����`�   $����C���$�I���@}l� $Gԟ�q� &��}��`��I$�I �$R@ n��C� K@8����7���	 I� �|�$	,��;���?�� 1�#��(+$�k5�����Y+0
 ��d��H_{羅�Q*"
���ET
��*AT"�JIY"�"���m�e$J��cf���5�URl�V2Hlª�*�1�S&��l�j,��ݝ����V-#MRh�km��i��U�aV�i�1mj�6�V�m�E�a���ce�imj���Mom��l\D�h��b,�0͚�1 i�[Z�f�,�) mJi�f�Ʃ���5�6M�L�[-�)6�kͱ,��,ԭ��Ҷ��+m�i[RɋkP+Z�m5�5��  -z��u���ޕJ������浻:л����g�i^M^�v��2mJ��m��]�l���s�6.�]�<y��(Ouۏ=Gw�7V{�l�SU���Vأ��Z�   �=
CB�
.>��=�
�H�=|���CB��-���x}
(P��}�(]`k[k�V�k��ֻ]���zuWn�o/7�{��6���=��赝���=V���3��]�SMT�M���l�   ����v5\�u�]:��q�n�d�{k��vk���n��]��ʽ�s��4zvfj��On����{ۏ;�S*����m[jiяsRUm��"�ͪu���W�  �>ۥ;����=��wwa�c��{iJ�x{zSb��wj����ӻ�wn�g���ytq��kE��{f��(�@�F��l�
 L[��m��R�M-�2�+mJ�   vz���sM�7[wpZSuʧ }��yR�
J��zUE�˚*��u�	��U��gz�����5Fcct�f$6ʖD���  {��B���c�QT��5$ Zr�*�Z��F��v��' J�������� P��\ �Zw':� q�mb�f�f��BSed�� �X4����8�Mv5U�4S�Z�eP�U��Gh(��]UI�����ny��@�0 ��(KY�*�+m��Y_  &x  T{�}:h
�ypt(K3�C�(hC� J�{��w��  Oy�@�<���J  f;��A�W�wu&ef�e����k[Zվ  �� �k�f�@���: � 4s��@ uӀz7f���� (Oc��l=p {k�  �Ҋ�f�H�h�5 ֖π  8� �(���@ ��8= ��{ ��n= �J{�.  {��ހ ��Q�(t�'^� ���p���|���R����4"�ф���h  OɒyUP�  ���R�   M� �*   z�$��  f�矏����_�s��W����܃ٱ�+P�#�Q�춥�D��b���U�R^������S?���um�[oڵ�����Vڵ��u[j���*�V��Z��[__�������_��9��V�6�ˍ�u��!ɉ:�5��Vb�àP;m�ɑ�u�Z��M=��GZm�n��a�N���R�b���MR\9�2� X�ӗzp��(�rň��#(�h����!�:�in�RI�dKĉG�,�pT1|�D��N�9�i���dmC5�-�kM(�[N����ŲD+!T��H �h�e���R�Κ���+.MjC!7p3�-�r]���Xqe����!���"�3jS�p�օr�jrՂ�"��ʗiC�묋oFT�4����^�ºrK�7T�i����=��Cy��I��	�� ǩnb�4���+hG�wha7Tp����X%Lͥn�T�n��tw-�4�s���wT2�a�k\)�[D��w��-�`L˥dVPm�k���Pt���S�n��J���Sw������,��^t�M�hN驛S:iEZ�F=�>z.-���U��k%� ������MjjM�u�Uf���M	P�oZ���h{���K&������m8�W�A9CE%����av��}��l�Zo&1]�7Z����"T�qH��xR.$�Q��n�k�,f�3�E��X֌6��գ��ch�ćfe��Pl
Q���o.<;#�X9�,KK5���:J��%=W%j�Mƪ6pⰮ�K���u��h`*�-a��Bu��m �u�]X�Bp����)��3wu��yQ�j����̒��ՊfZ��W�������b�X�[�Uֹy�����d�+U{���P��w[͢$����oUD�wb����ej�h�!�z�|Zp�{0U��é���E�`h"�A�hR�=�n �;G~�p��R�1��e!��x����F\�^��t�hK"J����'�qc�Lw.VtJj���]���vf^4�`Z�K7�,�m��=֥���L�^���K6��'z.�D����7,���n�T�Cb��l����6p�Y�n�U���F�i�Ѝ��lY�^�J�Kne+pSm�Wa<���a�$݉����#-ֽ���ݬn�*�m�8kS��bx�JK��pG�� �֜�n��VK�x�sp!�=�
f2c�ZC���V�5u{V�ذ}y��V	t�5�jj�nК�ޜOfK������(`h��賎���w6*�C�ް�����Xznǃ��|����59jA�sL{XQ.Z쵛���{�ʂ�Y���-�l����R^�f;wY�NV"�6�ûg4�-���j�x�hæ
*B��\�k�X�u-V���N؆f|�B�G�ط拠���|e��5^n�	ym�2�z#��1�����4*f�lpF�WgnR#v�r�َm�D��om�8$��em�z�I,4t� �x����ɺ�#en�ڶ�1LO6+��	>�Jw����(l�w:�l�	�
�S�Vkh*i4)�W��CN@$!h�F�VfY2�X�е��v����]�
º[A,�� r�aO�t��7���"��V�k���GK�uܫE�t'3c�-8q9@
2�,9l�����L�N���H�MF�ۅ��2�/V�������AVe���`G�[v,�"��Ez��e]hö ����8.��-�lV}��F�tFfY����l(0pX	�orI��D���Vk.����&V����-[w�\bڛj��6\��Â�M�ZB�J]��.[�@��[�|m�����V��t�l�XX�x���Y#\FX�>�ӄ�#Y�����#R=sl�֜ĥ�y$�&�Y��m�t�f�D��tE䬍T2��t$��n�u�	%*�El ��Lw���%a��G%���^�,'�D�3��!m��/]��铅���Z�`�M�[��{��(%�5#YV���[�7�)��)BA�f�,�
�6���PaSl\K6��(�V�(n9wwVl`	xKR�a�5%�P�WP���D�D��� ���T~& N̠K&'l[	����6)
X��/oV�[���#�gK`�3oU�PX�۵�i�uc&-��a��Wq��
�b��i3%�k-jܦZ�q7!Ӷ�۳���F:��ޣl4vQ��AG3I��%��4�D�%,x��k�5б�d��];�P�����7t��lB�V;��ڹ�\��m�bhVB����:d	kn�]"�@�f��Q����\m'�l�E����T�4���͗���ؠ��)�h*�jX�H��- �4m�A���V�mܼGqlXf����+T��U�F����#�6�b��'��К�R-;+C�U�.�qc��pkIP#��W	 WU���\��X�ѫwf%x�
��o��!��)Е�v�*C�hM��,�*����Sd�A6�����N�aե��	x��a��$��=�36i���7���Ţ�f�̓i�2�j�]�I'��� W�F�������:��W�r*�9ymn�h�ȝ�{nU��/C6J1�mإ���S��X�#�����V�Q�4	��Pt��MCP2�3��d����	5� ��s���^ʺʓi&�u��d�"f췦s4���bP�ݭU.�᳉����W�R	z�ʗ2��tA���NŻj$м�*�ѵ.�֭/�+�+�Ћ(��E�ܑYU<�"�V)�y�a���̸i�bҩr��i`��e՜��$��asa	J��ɚ0��"o�en*Om���͢�q�'QSI��h�F�hջV�:p��v��"�,���v��	RY�ʡZ�b���deﰮ�%x7B��Բ�Õl^p���f�W�uRiH�=ph�Z���M`�Ɲ�h�ᙂM�c�/[˖�.�1c��H5&K/H{�o$��0�4�u��i���� ��n�ѹ�ծf��H0�'��--6�hX�B
�	l�9�b�.���LD-իf�65|N�8aH�,�K$����4A��n�CqY�R��cY��I��FW����w<6E��C�ceհ���ן=���P�m��{�6اD�n�F%u`�v6�G�&a�*�wd�R�xi��
X�ۘ���,1J�"�эϐ�]�3a�y1Lw&��J���&�^n�U���)�ʴ�[	���>H�PZ��[O��#7��+�1S�:���1�2�,�,6���� ߍ��i�F�����f)��*8(�ˏe��H�*h�V��AF��e=P%yN �ݧ��T9�KlA\�r���wq������dH'���ل4qV�&i&Ç-ơe�{�+i��#D��)k��M�%:�J���5���7u�v�n1]�I^6%���5r����,`zf��ׯj8M��݆���N��HPcӛ�08���[�֙I����*M�FV�F�ȍ]1v��w�]nK�m3S#�D��9y��2�nVP)���Z������4���oH�X���*�5��-��!�VaKm���(f�������
k�X浊�TL��S	^����Ok%����#v�u��]��ʺ(uf�gktV"Pφ�Y"Dࣷ��t���͑E��KO)��$`Ͱ��e Ql/�	A zR��D���uso
����ǩR��Ի����m�q�w�(F�5�P�l�)��	���sP��ދfL��T���h�s5^$��XĠt�B�A5b�ݴૻ��z���F圦J������͂���5����)
2��.a�G+M�B��c/u�����c�N�ۼ��
{��*7��zEjuq�ǰQɠ��#���^��{'�\_;��if�]�WA��UqV˫{��ڽ�NP��Vx��ACہ�{/4l�a�Yj	2K��%V$x��̚ɺ�*4ݤ>�H�{sT$�C�w�\��9E��H΃|RÐf�R���kHG�xt��1�7�	I�:u��!g�,���.\ˋ)���B�`Z��gsШX�^�IBW���(Ț���A�&�p�J����!��.�����̩mZ�*洮u�%�fZ���ڻF�Q>�9L��5> &�U�=��q��Q{BDљh5oR�1��avȝ��dE�"��r+Ot����	.�b���7��r:�"ͧx�A��V⩦	�-�ƕdY��(+�6䚍i��V�l����k0_$�q��t���dr!Vdu)-�ɺ��ݵl�f�Wˬ��,���Ay����T	.Q���!���930�=ͨ�G1JJ��b+��LgɷZ��r����ò�3a J?J�W�2a�K.`��˙J���m�s5�aT�H�lӅ�c1��^e7XU�%J`9a��T��'�a��`�8o-�;1��� ��j���-��F��6�X�m�F,Y�,`Pk�T��Ѕn]�Le�9�˭�"��f,,N�B/.�if��˕g��-�t	&^�#b��\&��0F�V
)6�b�{W�!�	xMbq�-P<��ŀU�n��\��*�978����ԛE=�Z'u[�)'�ن�U4D+k
fKѦ�9c\��r�^���J�f�iP��jS�wE'rYU�㳒���zA1)��vn�n���������X��ȯgZ	X�t�O���xލ-0��ވt�̔(E���l�"]��w�)I�b5ha�x�śIkGD3��8w� w�3��H�l5���JɅ� `{z��H�M�a.90�m
P�eK��<��+h9�I3�V�I{��b\ٌ��{IXR�b3�+F��{Wj1u/ ]&��>"(���9���)�oLXp��d{.*�Jl��h<�	X��!f;	,���ĵ.����,������ˍܰ��]��h��Jجմ�&i�y��Du�of��w�U��n�*��d	�)XA[n���Van����/1�jGB������8�5����,�	f��P���9��H�%�HZ�Y��Y:e<ڙ1���9��h��\�q�+RrXӦ�=�r[�v� �׻w�QP�	u����"zq�t��陔�u�hF2�M��F��Jٯǥ��" 2��MH0�ؘply� i\��[��1D��v����^��Vi;&c�A�]f������k);��p�T�ce�&��!zr�j3GE���f��B7p@��'1�6������0VXx�,թF����5;uix[��/IV�կ�Bׯ�wm��%���i�r�U�F.刔im޳��K>K8=d�qG��t��pPA����Y�cae���ݚ]=�,է�%Q+p+�ȫ.[-m�Ӊ����?+t�N┺ơK;{����!t0�	�kvQ�X������E�HtP���`���?�S
@�ҳuq7*�)�^�YF�*�ȕwv�+�v�A ��$�c44(�r�
ټ�h]乮�SS+(���3ko+!ڂ:1fX����еtk0^-h�:d�p�9B$�K���1��Q���Ե{
2��W* Tz�B���&n�X�ՁF�4�J;��d�a�<��	4(U�z���i��i�A;�!GVM���;�n��5`b4����A-�����ѭԲm�5\6ke-��1��z�(�jǄy8F1�;OA��y���3o��`�F��А���[�.cI��#FG�-NVh�2	�wa�y�[I��F̵,Պ3�E���hl��v�ܒ >-A���TVY��T�h=m!���#ӎ]XЎA�����4���K"�~=z���j�����YJ�( ��P��^��q��@���l�Ri8|�7��#{@���C6	�06�6��|�TW��u���.Q9w�&I[��`�T�&!S�e�KT�E�!����X�QRոF(QS���� ��X�X)��w�A�R�SnAn<H��Ce\Z�Xݙ�I$���]f�ŹY�idhaɩ邬̥v&�v�e�%*|���r�f��*7rd�5��c;L8E"7�f��ḾbI��sPɚB�^4�n�(�|07�W�ehy��N���`�!��0R�n�wT�Yŵ�#����	2й�ajMyZ&��")�xEu��m*I�qY�2�E���ha֍�Vv^�ڛJ��TJI^�-dm��ˬx^,ٶu]���lz$��(f �%�Ti�`]	V�X�Y	�F5�b�X9)RRa묫VNIj�c~��X��OPˬ3T4�M���Q��f2E/:RS:�FE*P��E-�y*���3���(ljJ.�?��"�;B:�lGgSwa`�_�q�H���8.��+h�BM-Tl"�0^��F��J���ܓUùe(-!�V�5�י�Yd8v^f��0F����E�Bhkx ����Cq�:�H�3 �2;�H�l���@�R�h��e]� ^��'0���H�v��핢��Q�cZ�IX��K!�0
ph,J��]m�Č�I7)����E���FP��
1e��b�We�az��µIю�'e�t&홮ȥ� �x�Z��%-�*�&� @�݈�Dk�ٲ�kRS�f�^�l����L�Q:�Y[[�dм݂����A�� �Q�V��1��!e���u�hGK����/n�w--@[
�;�r���M�פoҶ��"<J��f�CZ	�:%�Ԅ��E$V��b��x�Nm �nZ�n^Mq+��n��9���YWu� ��hv���-��[�Dӻxq�wW���oͲ��u{,S���mkŔ�V�M!J�å.�O�[�Ҙy�]�˙���F���s#�����Goe��V����WJZDl�VޢՋ̫�P��Rd
���|���b���j�Q^L�]5"������cwu��)�\�$G������������,�{���Q�U��~��t��NҜՒ��@�+��'[�}u���Ty���.-=ev%�v���Gp��v�B�S�m�R�Y��uި�5�3�'�j�ה%�6|�ߖr�ڄ�.��0i̾>[�fs��$�E���47qT�p��W����ާ�!W����+3����-=w��e$�o#x�+�[�mZ�(���K���Z�(j[��;z�T�ޞ&nT����74֣��vMC�^���Gߥ�Ev��+3�Ǯ<�¹���0�vW�y��N��E�\[-1}u���Ν�؇H��/b��E������2�A�x_A���Q��'��Nk���7��q�F��UjlΗ'>V	im���o}�c�^VP�ӉJ!��I'��fGr��֩,�!Y!�v$vDܧ������Wa�Ok26���{e�1�,TGb�˯��h������j��d���(��'����t������n��Z�IK�]�)��Uby�N�ema�\��S{����߅d14�ʊ�rOwz+S�i�/�N��F�@�Z���5��	�{8;��r�
�}���ت�۶�dR=�kQ��=w�˸!��0��F��ϱJ���Hz����jĩ�x0��
b��
��t�{���ǉ軝�GL/%K��ͨ�4����kq�:��V�S�6�wݠ���H��1R�,;��Z�.���G��yw�rl]9���-��oH
�sۣ�{ �� ��nTշ�rޫ�pٺ�7�]�<��x��Bܬ������q;�Q2�5.ݱqi�9�sq��o��v��Xi����/%<Y]:���+=��oO"���n"�Z��yةeXjf���VAvZ�y�����������:�aޠ�l�]]_�復7�q�^<]��T6�u����1`Ѯ[�RPE	�`�0�]���e��g/?�>�vl���]MՏZ8s@ʫ�U�3�z�2�"����(�6�3ՏZ�;�ݘ
J7{�	����|U�������Neg+�M,�n2�JxS��RG59���=��Gv�j榥�"�8�:��H���5Wm
����ù���5���Ҹ[��aW*ԓu�^�ۖ������/'�2��+��'(�E5F�(�	9�u�����cR9��{w([���o-KY���\��5��cj�N�V�]٫χVM��sp-u��CVDE�[��}�P��}��Y\.������G{��T�=���t��N4/A��x�7�N����Ohed��^��j	�+34�D�
z�nv��٨����맴�,���ֺ_%u4uZ<�/�;�5�¬,r�5������6�R���#r�]w��b�Z�v���XF�� O�g0,g1�R��[@�^�\֫�ˆ5�b�g]���9-Z�p(`�݂WV��,NX�[�\۴�Z��S�:���N�jyd�۫뷊���l�HF���+�h��K	��5���r���4\h}u1�ZX�ݚ�8]�]Ԅ~5�lT�[rF�dcq��u+�{7Tܧ��wS�w�i��ǩ��)R~���}�1���d��e�u. `�$>�$����o�ew���HMgjP5�-WD�U�kCG8u@�&���,��;1���}Q]pwҏ�Z��˙�Su+lY
�紫�[37i9��bې݉�k�@�mp3���)��Y3!K+�W��Y�:h���������Ci��(���@�!�������G���Wv�NR�.1��*���D��z�t��dX��V�+]�L��}��ʁ�mV�(;�0�7�χKZ6��Y�;���ԛ��<��N!��g/���M�9��X&"����ɖ�Kx�R9\�!5Ի�'os�nY�I1J��jPP �d�G��D�n�AN�v𡺘�y���;�����aU04^ѩM��
�=5^ۏ<;u�U���	��98�=L�;���;�cX�]��L�2;r"��f"�._ܭծu3���!� I��[Va��4�	��-Txc>��	�֜y��2�Sôź�gMܮ\A��yX�=�޺�gK;���x�^�lx��:Rx*�E�N��<����X��َa��Į�gdG���M�805�bƂ��1 ��e���wIL�t9_;� �Go��MT���wST�w�H�Jk�.3��J��r�6��!p�u���F�s��.ۧ�P�Y+�kN�+k:�uBr[�ݩB���t���W��:���������ށ=tr�c�8���H�y3���q�gh�X�^N�ڬo�k�*��Q����E�G�1O��o��`��oMT���{J�0�I�*�mZ�V����NdjԶ*AfR�.�F�3���Ek�yt JnRٳ�����M]�8mRset���N�Q���{��<N�0��Sz�=V����3�Ղ��Z��vu��7�&�B'8�o@Ϣ
�9#�7ϢGݝ#�1EdD1��5
�VT�(ÕiWr7V�u�����3�cXiIb�� _ ��ˡ��B��A>�]��%���x�de�W�YhgI&/u�z���(���MV�����C��8\�r���kB9X�ù(Ф9�By1�K�#%��|b�>n�a�%f��앃w1�9�_=��F��g1�`m;��|�Z��;{9�ta� y'Vr<����<�T�j�9�W8��9��Y��[z���筯��������`2��y�L�g��� ��Zwr��*�c�s;�ʘ��q��9���X���q�J���q٬��V'w%S� ��X�u�V�s�T��b՜��q�S���tV��M�i�V��f�]�;�Q������WA�#�#�~YKx6�WQ؝�6�Gs*2���*A�e�1olZݧʶّ���cH�� ��SM��s9 X���1�*��b�G����.�5S��&q�|��h�~�˥��N��'+Kԥ��(x����d5��۵-s`tڲ*�>3�V����"����j�\�itڑ�^ǳ���}PɆ�sdf�g���:�f�����tT��_�
	���mfS͏�E��FE3/����'p!�4�X����H�A�[囐}��\O��^h4��Ry�am<QMX �ԺMA�Of��~�]���7kC�ѱ4ߐ��.}xu�m�&�1����J�Wޞ�0h�8� ��[�7W+3�������^J-�/�X���CVϧ)p��g9��U/���d�h<�P۬�u��N
7��h�Y����!>[���k[ۓ@��<f�� ղ��H��[k�2�]K�Pn��(M�͙�yB�K�-}�)��0g@��$�z��@T�ۅѠ<��o�w�t̜�N/��[����m��jx�2"mQa�8w8���Ɂ^lK����7qi� �B��Ў:�{j`ډ���ݢ�
�ycw@��Re�C�}H@�)�#Q|v�O���*:���=����L��+��Q��7k)O���Ɨe'5Cn��*�n�I����'���VM�~����ɬ\��M�G���I�{VYT���.Gaԩ����q�OˏA㜳�񽹤aω�KR�d>	��Y=Ycz-=�Y�K�K����u��p�O��mv�Sl�#J��T5O�ܕ�uμ��xΈ��Çr؈��%��/��Up�\���5�\��;ej��ML�3iۋ��*�j�PE�F^=�bw׫w�������Ԩ�H��1��S��-�5�8B\���t�Z�2���B�f��D��>����(�J�Y�y�ry�v�_-+_4o�%���	<3q�4��H����̙O�x�U�)�rw�C��ۛaD��b����hm+x1<����}�`�9:CX��I���}�:]�d�]Y1g��I֨��W#j�k+V2S8���o�U��x	��	g.�v���{7ݽD
�x>��^֠S�&�x�9�}��.zK��~�]� X�A��&��f��Dc2VH����S\;��i]��9�H�w;R�<�x�b�!]�Ӯ�s������]��7Ӡou�2�((Lǁ��8V<[���ѣ6��b�ݧ+��Y.�v�����w`�<\j37��|��W\tsab�A}6�ԝYx��+�}�F���r+��Sy7�x{��=zo��,�W#��0�vոr�{Y�E��o&����VT�����pÕ��厹����5�E��0>Y���������c].EF��ص8�F/wM�dw6�{�4�頿j��rnm.$n8�$�DE����խ<5f��bH��%��W)ME�D�+]�r�s��p�	|���-U��lNO�5�G��o%tZn�8.���4�:�$���3{/8`�@D��:e�I�,�5ō&E��L�����y��ɔ�Z�)�V�K��؄ʷ��.\a�y�6Ųa\�md G㜐��:����*z��&LK�o/7�� U�4��.ԡQ��f�pܾh=�t�ڰ���B��}-�oh�Y�L�GCr��ŻB�ax�(B3qK��z�v�T5�q�4`"h�U�}ļz�����չ)��˝=�,w���k��M��=u{C)�j��4�M�;�_83�ݙʁ�k���zM^�f�����I^��t��]9��逹 ��J������z��B�x�l�����ACI�u�9\�����N|�V��V�U����/��j��WRi�ʫN�m:ۢ˴Y�Vo��]��'��ng��nu�m��B�Ռtj�3�������0k�7
�e<�nv_}W`�h��Ǔ�w�{�{A�B�6��T*��|lW^�6<���.e�g=�-CS_$��*vD<�$��I/n@C��Βd[E��i���+=NL͆�yN��z�frc�*dV;��8e��:��YCo|�T���=�L��r����#Y�M��}�Z�귤^=VmP�Fۦg��PۚӰ Y3�=���n�}�7RC4��M��c�y���~�p��=o��`ҟv�3<�պ6Unͣ�:�f �/2�V^�e�\!�wx�T1��ؒ�w+�բ�7%+u.T�fE������(�v��oVhy/�Fﲌ�C�F���k�+'K��*��⿖���[߹c��J�n��]��L$	y��d.����q��RaŢ+U��n����>@�6��Px����>k:�-���9E��/w��r^�n	���7��)WG��5��Tm�������7C^�&�N�i,M�˃ie�η�Κ�|i��s�]�D����m��an�x�@y��s�z�G8O╙;w�1(��vq�M���^�J��q[�R�܏ɍ���y��QW����3���;$��}�1�1,(��8u��y�cW�s��|���W�D��;TUdn��=��ٻo�Uj�g�`	�1ʞB57�ڈ>�e��tfb���sMN����M�s�S�(���ȳ�w��Z�j;z�������{r7-��[F��W�����OvT��xi ��E���4�C�G"�7r���,o�x�@��H+d:��mc[�õ��((���Z�Y����j��^��)J)<1eN�Gt��7����`�[�L��m�F�ym��wse'=�GʆvbKt�¯�,�.�	�}���s=9qF����FH�a3�Gs��j�T#[Ԯ�ذɷ\���ٹ-Q��0�I�0���a�P��l�B�k�F�
C�'��&��$�Gu�pr�.)��l\{��4E�ŋ����akCgd�õ㗉Z��ה��n��Q$�;fV��+�g)}�(97V�=��и�jX�8�u�Z0$��#V����7�¥���pwK�[�B+`uۋV=��*�iM�a`�K�˫�n��C5��85P��
�3� ��Q���o`e�ۂ�l�W�zy�W!�J�vj
�7��gŜҪy����fuY�yZ
��; �C�n_���bu��.�l�����M&���<��[���g����W�G$o��_+Ǥ�=�ڭ����J^��2���u̣Ϡ�f��ܛ42�z(�Y�����Vd��;�b�E(w���,�˷)�F\]E��U}b��in+���)f��@���F��7u$�tH5]�&�*C���[�2�f.��1��8�7OE�Z����l��b�fy��wF�L#^����QQ�{�h�⫆b|]��d�sE�J�P���Z�a�oB�����#uo�s/���>;���|��LF���������{;7Q�0�N.5���\���mء��s�sD�y3�Hx��h�l�Z�JX���	���w#��.0��0�3쎣2�l�ς�FG��V�r�z�≚"�Uvz��2��h�G=3�����-�L u.ZwE���dd��[_�8��D8���u�' B�N��l�%7sN]@1��y��޻�|z�I���7"��$+��OG��;��b8{7�gp�H;��)�'b!�O�F��p�7����M�oi�L޻8nJ���Cvt#��b=��w6-u�WC��̕��|-�]�z	�`��JH��wuα��=�o��',��)�Y�_��TM�J��I��\���"��r�X5B�sa`�V�&nd��dqT�K�fծ�8��V�^>��au[�?ewK���Rw�$X�[#���\t����dkL�w7�>�=�����E-��(~L�.��Ni����n�p��F�܄v,�wϴ]W��%�Z��Y��חv��ܫ8Z���Z�r�̼=��]���-�{��{�o�k�������������ws��������/���꯫���r���Q*zI�Wq���ػ��(Q��o��]��b�|c�kK.�o�J_x�SG%�Q�f�&2�AD<4��"/�t���OmӞ���̃d�������[��c�;��XL�1�w�ޗ��77a��U֪�6���{��Y����K�i|)�n�E{���p��Kϕŗ%�o���%�Ɠ)Q�3�]E1t�_og�+����t��p�1�=܀�U�m��!;s���orI&��� )�����
��w������1����-�%1�6(��gj��XH��m1�-9�I�=+���&-搙B]��c���_�ls��X)���
P�uZi�7tM�){Iӧo�`aڼ���ڋ1�1���g�o��z��׎&ˀ�C�E�o�ö�\LWיK���Z4|9u�͇�V 4���y��@�M/�c��N�H�X��ᡤ$���궫s�\���7�${fo�HԦ�7�H��_�3"%1%E}M�3/(�tC�S�&Y�+H��9�R��Y���ŋA�},%ϰ.��F])ܗB5����.Cq�,k0�:B�6��pD�5g�r�%���'I����E�`xA��Lw+��&RL=a��6��T�("31}�C��p��V�ԪQBw��x��E�ǋI8DOo��N̸k�&���b�촤S�)S!�R�.Ί���vc���vnEi����"�T�2��B�2�e[������]n&A;�Xo 
0������=7�m�[�{Ъ�AV��wR1�+�M��q紀��涅}OH�v��Z���}�N�Swt�]ܙ{L� ���D�Xhnw7o|���.�JY���C���[�a�t�)$���+��6���S�	���\�v�v���&���8���8y$���Èg.���w4����'i������r�h�Q�v�xK��17qG	;si&8�����G������;gw<�'ҴUc�DK�0�̉3}R�MhM�1��r��h��ze�s ��0�ӗw6F�k4(���{W3�@��]��Tܽ��Y-p����)�X~C��jɮ�$����s<:�v�����ƓcV�<��ע.L�T�Lצ��xgM�0�̊u#+[[���b���Fɔ�H��c�drgPϚ�;�Q��ʓ^�c9�ɜ$/j�[
��q���xaБ�����E㽺�X��H]�p��׌@�=�>�v�C�j�X��u�g^9�b�W��x�(���lW�F\�
Ÿ�g�9(�w�b��(���t{CNpu�,".��X����聦k�	!��6�8	y]c7zv��[ZڳK����.�Ds}�ɍ>����K�O�Iǃ4��]�؎ie3�dK�|}K.�
���5�)/��D
���;V4��/�y2�)!%�����觽�.ӳܷ���t��v�u�m��<�:�vmA��a�c%]�E'Ev�is�Ý5��e���-7�����ڟ.]z�kr)�\�kb�7B�b�9��ϫ�5ՠv�do�G��`cg�w�,'��
��-J]�u��	a@�w3\��i���%?�<�\ˣq�Vı�tGv��Y*	��V�V�[Qf�w�Z����U%®��>Q�<�7W}J�*u�C��7uwS�1,��__,�2��5�Ը����b�O�h���C�w��w�"�s� ��V.Q����'4�C�rg��bk ��b�=; 9��>#5b��Q]T~�Ԟ���^X=c\���>�WVWA��-��2�ax�-�!԰�{�V���K;k�oot(�t��4��Çd�9�N�[J��A�%Cvp�s�-�.�i��w*5	�����ZY���.�9�X������WPXH�M�b������k��ĩ�����b2���7,�u�<ڳw�#u�W��	h�yY��n�z���܄M1Qlom@��+ J�hen8략��E��z-��s�u�3��
^k��v��C��>�6�u�I�Đ�S��S9lY��r]]�Eŝ�I���RQ��v�d{�S��{o�v��y�W:W�a�Fh����z�}z3[��T���M�|���=x!�i%s�r�{Ìn�N���]��q��y�h����9�ʠ�fqN�"!e-'l*��1�k��צּ��aJ7�\ugF,=Z�
�]��V��D���İ�k�H0�(bG��-s�L<��,<�k�ܱ�M`���u<{�Q�
�y93Mc�6.�`;�m�Q^��g��qབ��Y�X=�4��\��چ����}�DFL��]�j^ׄ�2(Z+^b���N��[o���f�+�yδ�Z�9�;:G
�����v���l����9]��j�JT6='-{�#���&@a��x~|����1
ꂃ�`R�f�Ҫf[�<��K,��8vTX�B�;���J����釫&�=Du,��s�E�5�50ƒȬWKIr��9�蝤H7,�β����H�/�N�:�V����tܺԜ���3_3��u�N�ӹ�+]t��W[�S ���a�.兣6��ߗ��ŝ�c"���Ǌ
N�m�c�]�������V��u����jcG���-��7�P��9�S����p�
��U}���Tɺ�j2��u�W�:�m�Ju:��l�Ei)���R�ț�L�_��Bp]�����w-D�v���+P��ܧ���&mY��}�}��":�$�|un�]5��V>��q�8&�b�K����@M�f���_�Iw���#8�ڇ#���m=��ݛt���(<�[��&d�SA�.>:���l�ż0�}�xfXp�k�UZyD�=YGl͊.��b7�&S���V�Z6)�������\At�'�V삂�V�\�,��;j��H�
��7_)M7��þ�̐�qh��9��mg�zиN���MÒ�p���51�bXgj����92�j�]���u}M���Y:28�Y�ݸ���ؙ��T<��]�m���ȋ<�1`��^9�>�3}�򷽓jFZ�Hv_RP7��k��.Љ����f3��o�%���Uu�ʹ7����ĺ���w���-Pɷ�0�O ���҂U;1�oOs���ES��ޅ{K/��NJD㙗B�=��Ȼi�2��"_'V���Y9�n�e��������d�Gx�t-ŝ�}}�F�a�9Z�=W�4�|.c��C30��;�8V(F��iV� ���P bu���Y�L3V��\o'J�@j��ƞ�5� �&�0�ɱ���Z��h�h�O	{Ӧ^��WSOwӰ�âĈ��u}j��S/2}���ZY]:վe��]�V�)Ig�j�SErY���\�jҤoC��tl���w�[P�]�fU�6㾮��|O��5Z�-y���{.r�/�����tYJb_^k���܀Z��KF�ݔ�W*�Aچ�J��X�t�ov�!�v̦�z&$�j�P�C(H�:�C�x��恵�oO��:�fpI��	��ڀ;|����V�씷�1k����;j��=���,����ze{�?8��zsq$]���"=�<T��I��yX�k��+4(�.˗h~���_.��:!�3+�����N��xJdc�.�������w�P_b��z��u�=ʹ��$GD��ӊ�i�-x��d��ۙ��9fX3M>"�L��_B/��	�	��ုo��Uϩ�ȹXo;;Z��4�m�}/]�Uh�s��G4t��^��l��>�{s�m�;wz´o�EAc��>X�k�]��g;��4�ckT��N�n\��������Λx�/���0E;
� �z���/$��^
�n�������}��8d�n�6f�x�9`�͏��ུ�Ӑ�e�/�G�n��ȑ��1���9X�F��F��ھ��/��������<�/&N^��.vi��4gI�u�X��f+E*�޲�wa'&+�,%����hI�5��#�������S�^�q�ȑ�Vs�ψg_4k����9ro8m��[R����`Z��w1	�`����i�&�����/Kʛt�Gۘ:R]���� �.4�w{�����35��k�-ݻ�ô0�<���ގ���[b��Ǳ�~��U���@��d�<�oVTRtq��@��
�_>}�0�T+�:6:�N6� ���D�#Q8��(�#�s����eա�(�xo1���cL帅�AK<����E�:��f��޹�We;o�����$�s-�B�d��wT�X<�T�78����c��U5�w�k�]� ��v����_5[��`�Y����g�� V)f3�q�xb�b�lL�q��{���k�V��k.���ɩ���9i
����15�2fR{[��(�����n�ҭܢ�t
��v�0���@T���A���S}���
�0I�֎B+�E񖘬�+$�a;��Ꮦ�8��y'J���C���S�U��s� (�21],N�f�����ۘ^M>K�)h�7d���	S&��ŷ'��:���
�Ř���w���"��RV&�w�5ɖFD0*�$�觯�W��=�y�n��f��z=��u)r�xlf�*�{�	v���>��G*m�)���]�J�[�7(j��������p>:���l�[�:Γ��"iN��Bxx`LX�3���ȩ(�m̩�rr��Jr<�;����睒��������vQ�ǰ�����2��Y}h�(�f��4S�!�u鸪ާ	��b�N�P �*��ݸ�2�]k�%jZ�.���Ƀ��7���I��y��5L9F�7{�����Uu�:�ԥ[�)���ۣcL�K$t�j�ye�p���DDS��\'��=�4�=p1P��:�B���4 �z��)1ŗՙ�/3Cwإ ]��%��\U�X�[�h8+��L���X5���O�؛��A��2���C�����f��+��i��*c3?L]��6��l��}u�c͗R�Mfo.4�8CW��rxDU���XWy��u�w-��I��N�ZK|�+׋���b��ۓ-�]�a�צ�,nI�w*X����\�oi���z9 ��&��H�ոm�c
�7�B�+	b�s�N'�D�Ĉ̼���ݦ#;]�&�T&P�M�덧1��&oE�+u��儧pŬ#8�#��v�7�Vn)�h:�nb{�Ep<���Z�_T2DR��_͡�u�����nb�t�Y�G@�ɼ�⿣rm�az���y� 3��N��07s�2"��p-�}�*���WӀܖ��>m?�O�u6>V�pd|.��;;un�9ǲgR*�mw'���S�	 ���K�\��>�����M�3v�;M�xƽ]V�-��9�;K�pP��f�їڔ5���>I`�p��F(D����xJ�pU�<�4�`ܜ��b��:��%X�/fS�����d5��	�&P�K��oU��;��4��}�Kz9�C*ʗ�鈒�9�ۻ�5�a��U�ܷW@,��[})\�y�/g1��OJe����b-��}s��9�c-��8�V�m<�����Y`�m�H
�5r�cRB�4���ӧ(<�xϟm{��\K�������-����R�^����������2�Pm�,jjvd7�}��t���ޏ�=��/r����W��`k�E ��&��׽΍��B�cy�)of�k]���JV��ħu
�S�y8��yG��;��n>r�o[���/Ӈ-�����Fx�G_Rsףi��}9��o�C�*D�n��	d�(6��-��$�A�y��[|�j�иVn�_X��iУy�5�rD����e���Mw3J��/r@r�\�Y���MUq�@	�^����7u,ˮ�(�	ϰ�}�c7!��t�`�|��VB�_G-(]X�y5�r�!�U�N�*�87.�rϯ;C3�m�:819K���j�T�Բ�tp�6@�|Ӿ��m���YP�``��v'Q	��Z��ƌum�.����u�tN�u�@���]���xa}�yl�AB5��¯��s�Z�+�.��5���ͺ�˿��z�M�&��+E=���jܮ�{G��`ڋ�
!3W�P��!\t����ic�,8h�er�G��6�Y�1�q3��Yr�{)�RQ6U����:��/�X�_xW�����V7�wu�hYp.��v�ŗ��4�#I-Z�<[bq���q��N����z���"�f*��2:�����;���<����.X���zo1����!�����ٱa7����)hz�ḶQ�#7g	.�\-g��Li)��C����]��'>X������o0��<��3P[�e�tJ�����.����m��s�ذv�����֧���Dy��9�m#)�鑊�ڲ�(�k�=t���,윚3Y�5��9���o��T�@�z�ףYn��4�O�A	�X=<" �3	}4�8i���ܜp��0�n���.�8�P�����l�������=
H@s:��8����g u�
��ef=�*]�r
�]X^}�gTПQ�n �S#$���.�J��;v�[Ym��1�����}جh��%	��!''޴)���nXx�M���2p�)E�dYbV��j`]W�
}.,�jܓ��Jo��˓N�¶#�ՕwjJ�K	߃���2��x�C6�j�mӖY�U���o���d�L���elyd\���ƲLV�S�h�Մ��=m.���.�P��=gv%��b�	{���{�@�^�������6d�]��n�h�N7L�JE\�n78�)��mX���*�p��nn��2r]���Ӗ�9�H�n�0�e^��v�%s8t&ܲ�u]�*�Gn�G	'� ��-ŝ��aj�OFw��t�Q�r��p�=.(�Vq�&��㛸xg�UW�}U�}������[�m�^��N'�(tp�@F�c.ĕ\<l�����^df܊�E�z�P$s��Tt�踒/	X�Ҽ�F��Յ8�1���l *&��Ֆ������o4�ޤŦ[�B	�ne���1jC�c`����+�*�z�-�f�hũ��9���3��)׎���ѕ�]�az9����;�N�'�*Kqu^*�m�:������r�TnƷ��c��9����{Z�gM
�L�[��$c��q�X��M�5�`�Ҁ�̬;�eL�{��&5v{d�b�O/���"��=x��5��G[���.I�dCR^�삕�n�r�T$;3P��j!?�~XS���RN�tP�n���+��.�����R�RۋgbU��bt�ogθP�rHSwV:�B���(S��(
C�^�n(�	�����]�Ո������x:���Mb�|��
��2ԋ��P���n\%�K��Z�l�w@�.��b��{��\ҿ�2�?�`��y;�'�^T�䷃����VW+�N��g;�WS�:t2r`��C��%���!�<H�xΌ�{��Y�'+�Z�:����P�ZX�­iq�^��h"�A�M�����Z��+x_\�f�-o�w�]�ꀧ��D�h,���7�8��ohވ;E秦�XExc�u;���]Q��
�y#�]�j�o��P�Ȧ������������q	��)1rỮ��-�\����W9�67�&�!���9�����]v��uwu�l������%\�M�ӻ�2��ur���ۧ+��������sr� �	 �v.�J�Ît��s��k�:P&�vWw\�\��n�k��b5�sM'8��Q'�s��rHѹ�[��wr�b1�7(s��L[��H����[���X��6��]�w�ݮ\���w4r��`��+����ӑ�r\��;�Ԝ���.�v��f���s��r�I����s���)q�������c��+���$.�ww2j.�uܣ���ݠܹsS2	��E�3����~_�^���y�}??~��ls�6	�V���n�������+���Y�Piw,�4��r��]������E���6�	K;;��~�y�J����v��:6⨤�Z���F����ѩ�E�}r�U�E{&O^nv���uh�|;z�������,7��l=����u+�>��j�fM<���£��9φ��i��=iL5�Z<6ꅯ�ҏ��l}���������OՓ��8x�}�^b��l�Ks�>M�YE,I
�L���S�n:�[W6R���{ӎ��W�@oz��,�ʨbΧY���v}՜b�T�B �dNhn�8�x�m��iJ3q���gE}W5�J�с�7����;�\:����tڹ��=;R(�Hݴ�^8�k�s'K�,�<��� �K'kU �qwb#�:-�n{~yLGZ�[f���h�)��y�Z�a߲�;��Q�`��!�=��V-a�Nf���gGXrWjo�[�o��J�=��-�n!��f-Ҧ;"�G@�b�����}P�:ꑆ,����sL17�y\��%ťo�G9�9��6����4��l5�@bI@Gff��!�wq���Q��]\̲��9XW�`4�Ղ@Gh���wM�˨@Wұa:���%꒣Y�^8�bg{�X�t�K9�����'���|`b�F�ݗҏu�-�+EZ��+��|i����ޙ-U��{�|Z�Nor�m���b�)�pg]���!�S�����P{�����	jH�9z�X�)�!
�T�j#�����&ؿt�����K�ws�(d�NwQ��������P��:�&������ULa���b�	��x��P�N��i
_v2	Y.���HW���`�MZ�D��b�'�k�Id�d��U_˱�����Jx��L{�#ȷ ��Q�딏VDr���|�F%0����3qUT���
2�Mep6ä �a�V�k����&x�΍���!���0Z^��Ef�����R�nW��!��b��fΤ�s-+ :�Zc�)��x1aTEOa��T�zԌ�Fz��*���SSN����;�a���vxN4�l�� `���r�E7vE��Eb���d�D�F�f5n����a��ZT�#��ة�zo��-7���q���"�E���(�����+X�����:�!v� u�b�g��뙋�47Hw�8z���>x���k�ޮ�r�xUm��_Z��:Iw�۠�����B�*���
۟y���*���b�o�J*���7C���Xm�W�j�> ���"�+4"w!���fEN�O�	Rȼ�v���#��6��Փ�D�Y�r7e�q��N4p����:�	���i)O��!z�*�JҦj������M����|�͆.+��z���.��w6��v���-p�#� �,�K��b���N����D|ǵ^o�i*�?Uy�pײ]6}�/(�8��`���%��F��lŨ�Γ�bÏw�W���2pI��W���e���p��V;w�ي�<tA�_R���|����z��~��h��s��.������[�7Jb���;c돵ä3>,u5P�g�V�w�ǣ��[��>��,�WL��h�ۨ�t�p�Qb������w�N��:�`��7���RN��v�Yɥ�#����k:7b�S�V!?p���\Kw,���f������׫���%��`��bQ%Nq #�3�������]vhfV���n��xe+q��U�ip\��g ���mͳq,� �0��$0��2�7
j�n��k�ɢ(z�wj���p�[�i�p�4�}VJiL�B�31��Vh�4��­*�O7b�wc�QBCE��/�^���N�6xL��I٣q�W�]E+~��Ce�t�C��M�kui*���.�8]J�t�vhRĹ�U�xS@x5�Cg��zXx<e�U��קv�A6�
r�i��8W<��=C����=t�W����OF�a��Պ�ލ��CO�]��lWa�"tς:ē;�v�{��8���rt�]X�t�顡�W!q���A��{��&��7C�؊���'s��o/)$Άw,zcmZʐ��c��=�P�]z'-����|������5��S�ݚƹ���dұ�]+s.���V�wj�e4l���}��ݮ�.Kj4f�Y�7����fNϤ�x���Y�?1B��#�=6ʊ���σN��h��f ۤ��:����z��:�e�t��s�7T�����a�Ip��n0��s�=��&���Ye��S�2�Wj��R�`���3������B`!@��=E;�8�YhP���e�$��tY]XY���W֡�'-�ȧ\g�s�i����v����mn\�Y�#���d�S�U��,����-��ލpaQ��{/;Y�wj�ש�j��n�ʋ�jP��\�ia�l�&�¹��w"�u��v\L��;"��q�����VhF-�;���2ss���@jh�
�*�Xk����iD�:��E��ٔ0#<s�9���m!YE[�*ta�ϒ�z��)�%�}�?m���{;l�3����Q�r_Hs5a����d�.��m9;eR�cq<W���2w?n��gQ�F�Y=�x����A
��|��h�:5�4�/od�/s����̨�� ��;AWIg\��2�f�L��!9��z~+�����Ӯ�y�����
imR[�@�̝��˃�kN�lƳP���dJvٌ�oKG��ۨ��Ṫ�${�G��7�i�Q���ٙ�z���&�f���C������K��2v��x�l�G����.uc��d��ۍw���,��
+���	9m�D��	ﺐw�\�,>�����K�e���tnNݹR�����ώn�r���Ӥ�P(v}n�.טn�*��*�W
}��ቪ�0�P������:�k����k֘��~W��@��]Pl��=���N�%Dw�[W�^��s�M�	Ƨw��)ql���yv.8��˃^�|b�Z��(�/��i���xr=7��s��׉ G�g�#�ߥvey�3�3���2�'޸�#E,Im����Mó���{څ�]{2�^���V�΄����E�YgΩ\1�Y��:7"�������Eʎ�y_2�w6���xV��S�م���oMfF+N��;����3�^��?�vw8�S6��1�c�����䒱�od3��
��i�6�F���o�kᝫ�2���N)5ͩl9`Kl�X�n�%`9��Kr@���c����)7S��i�ah��TV�n�R9�ͽ���Ys�A�Ú+��q`˽��Č_�=�
J*����t��7�ṘI�B��|N
�>	y��>�}(crE����43b���W	�f�h��I-��O�߆��ۍ!l�&���s��U�]a�����$��t�z�mm�T�����x��3
*c�&�F�KON:K�_k���^ �tn�(���l��4\�	�����9�e��?!����i���@bI@�s7�����ϧzg����ئq��n�5�l���.+�r4��Kc0�-�RQ��|��ڱ��%�p�fGr�7DLI��El�5;�#<"��3�m_��w���;�����ӆ{Zڡ�u,�.���D�?8�̢*���=G���&3��4W&���"b�\�ż����rj/Wna4���@����3GƵ��qg	v?36.��ޟx?oW��G�B#�/f���_n�g��/ :`�&R�5(��	������m���|��n�Y��VA�\6��mL��&�m��۱|b�3��(F@b�y	�H���T3���LX�0�z�껊P�C����}�'c��В�!b�B����i���|�s�R���
�	�����o��ǎ���î)�EF�ݗښ�ݯkY�ϱ�\'���j��B��FM�\��n��[޾���N��u���ky�$�|����v���T�MF�˅���F3���P�P��N���xg�)VO*�����)*}ɬ!�+ה��T+�W7��N�<��y�C	Kێ�·Y�>���А�L��5�2�1j�Z�ј��(�ۃ?90¸��zh�0��m +��P��#,�3���
�;ZG���5�s�+a�&�H�}�ɇi���w(u�7k��KW���!h�s�jj�˷��'1ޮv�a"_�ט�����lX�h�g��YecY+'�`��:��%�ߧ�MkF.4���&��e���������ۇQ�f(����I�N�:	`�w���͠=��C/`�M̍W�ӘF�׾t��~Q`2��S<���l�i��$�;oz�㒃�K���،v��Z�����R��Jb���;c�����G:W��~O3lV��ӝ�f3��w*�b�D�ft	�{���a#ж�%�7�$^vz���
^B��ֻ�DP�n��oN��9;1��f�иB�U����ef#_p�O�&�[��P+�ޢ����*�-gj	�r��k�gu�q����"�Y�a����5����I%A�-�T�ɛ<��{�wyVr˗2[�2IF����5i��z����@�g����
\qJ���^�0�#�3.Ӹip���r�:fvf�u�v��V���oƀ�K��#�֐1!���A�����bH��u�K���gJ�t\��Y"�x�6r����)��f�yd:�p�'�>�(2L���l@��6ua��,�P��s���\)���W.�F���Ysl��W$�WQJ�ݑd[~m
F��n�%�^�և��hA�87J�^�+;�7J�Ƈ{7zH;���Ͱ���.�I��:��.�����;
�L\���+�0\e:zk>���U��܋�X
f���z�;6ؾn��s���l䏹e�;�~���vK=�㊒�_YvR���CH�����kU�=��zJ������*`���4��:4)��n��.�j�p47)]+5w����/��g`m�==��nV�&K�3���u0oc�{{?e0z���eد���m��m�]S����P�Ƚyv��d�
Φ����P!ٌ�N��C'=��:>�V u5~N���|��n����,0�lr��"�g�p��b�P��(�{RJ�	��9X�� N�^Զ�d̚y�J���#eQ��-���VJs{��]��Uk�mk��-�{S�:b��1Ȏ��ye�s;�nk;ͷ��}B�z)˸��h�Gr������w�\����$�(d����J�p���gz�|
����;h�ζۇ�����=��6ս��E��pgE�:xd
��VҠ�������t�_М�{�� �:��̰)�8�U���qC5��kL���T~�V��z���*�R�� sw�>�eu��I:��������K����_n5:�)4��a�l��-�}�r���u���GcPk5P�S�\j��m����2�������d�� ��� �*��N�uJ(N�����Õx*˅i\U�L��Y0�a����۲2��3_r@�_m�Z�#�;G�:>�jT���r��6gQ�FqY��T�m��&��p��M��ˇT̊�2R�W��2*��}Ӌ�Q_k��D�%�4.:�C�����m!�%�QpL[%Xu�c
8k�ڜ�x�q~���{J'�����i��Ⱥ�v�[��������k���?�R���_^����L��]��������2|8.<�v���>�]��]s^L�]mt�>�Zy���گ�R�&��Zu!*�$���Br���ඬXv~����=�BE<�J���R�}ô���k�{�"x�C��o����.�ʞ��B�ܕ�o%*)IV��T��+F�<�	 u-P��A��8�Ɇ=��U�~���2$��V_�R	r�����?E5z��޾�.��w�^¢ζd7�Ѓ(YO��!���s;�}t�<)W�S�w9](wB/�c��sӱ\�n����}�}���G�~�yf<�Ez�^U�p�Ϲu��q��!Θ���=��� a18{����ٕ�(���6��2�%\U���$�f��,���u����Fs���ȕX�Pdj����';e��z�C�\1�u����vDug-��R�kfs��؛���8�l��_P���������oMfF+N��;�GO
��5H�����~���w���b�r�M��)Y��I:!ibd�V�,�����!e�	|�uN"�N�沒S�R�g��7_Lv�;T�/�Y	9�Bc�p뜋��>u����i��!�u*��}�b����논-����y�l�$�`,vo�k�E��
�}5{I�S�|V�)[w0Q���5�[��2�某���\!q�*���_GA�M)�ٴ��ֶ9Vd���S�f��-��L�=M��6xX玻��#O^KeC�B+��urc������x+
-�XrEĘzH���v������!��Нw>�>ϕ�ʳw�3 ���֔G�!���d�[�"^��Y��6��>��v�(�R�L�aOV�C&�/]REJJ��a�O:׷�0���[.���'���(]	�2zN�G.�\Gd'�\ _S��D���ڣ�XV�^�՘ ��΢e��I^L�bّ��(.�]^Ǹ���E�Q�۲�<YQ�צ!�u�h��ˢh����r݊v���B�K�.�pj�(N��)�i�D	ϡ�/n%0:5f���Z�O.��v� ��YB�oSo葼��S[�_n��5l`᝔�[�d�&6�أ��Am�VooIv�W��5�����Z)���a�d]��c�u���ej�pY��*�6����TU�Q��!�)gf�;�j<%y���n��b�.�߈�ջ޵���ĝw9�.\�j�wx�_�ٍ�,DXf���'���z`���O�m
���ho3�����篴�aem�%��Na�t���z�w$�'m���]pM��D�Z�{D�Ƃ�y���ŵ��7;~��>�
�UtU���[J��m$��R�U;E:0� 8K�#��u5)�(��;�T�Їa��,�d�O��K�,�oV��Y������k���i���k5��8����
�C[�WZ�F���5窴n������ή�c���_;z�f����eKa;�nƊ`�I8����[,���U����P�V�Z�����p���V�R��ڱ}q���M�7]ڳK~Q){���V#׫�l2\7@�n����Z�_R�����v��Xʶ3�ѹ�L�ܸ������{%n�]@�s8�H+�H%K��fJ��:J|KU�����ּ�j"�A��'֫���.��n\2��9���l:j�������vP���Nu�S��w�\X�ݾ��Ǆ,��3i�,[O���ͬ�wp�ȚS5���'Ѿ�(�.��"rf8Պ��x�$Ȃ�)h�9�蹪x�є쑉�,�X��[�����;�gM!����7N��)�Au)mc��
�ƺ�Y��RP.h�q�Q��]��t�܊\ϭ�W�W?����!]'z�Na�Z{P�v��1��Lt�i�<�%�=����BdJ�Enr��Q1�0�[�z�A����w�*i�ƭ^��� b����4.�	�@w��r�e�.�ǲ*��a�ߏm�w%�f��@����Z����,AyX���p�}G6�'�v�]���B�ȗ�{=G�=ͫ��\u��p�B�5��:����\�׀�9Y{�f�����#j�NCg3w�ܐp���p�7�U��dSg����S/�����>��b���9�٠/L�$��`b�ܖya��	�+.��o%�+x�0��]
{n��r����ڱ��o!D����6��7>S��ٽ��w8�1�۶{l�W�4��(�Z�1�mtw��*2���ߋ��8��'c�U0�N�r�o��v� *ޛ2��Qť:� W�P�4\�3wtkst�8ciI,\�K��rdS9ˮ�wpuН��sN�b 4dHwv\䜺H�B!]�F��wws#2wr�%.�70E'5�7+�"U�;�J���;����� �ۚH�r�D`J�)I,����n�r����wv�t���@�6��.bJf��� n����2��f#����fhÜ;�hB!�v��vSn�R�v�]�Hr�'u�.�$��1˻�D2e9ƌƙ1M����Jn�)$P%.tE.����9;p��捄1(A!H�.뒈deݺ$����A���-�P��KD��@�FJ�
�n�ŀ�� �!��I����u�L�}��}~~��~?~�qo�z����!҇f��ʕ�-�Gy���˛ٲ��?�����ᇏ;FB�M�7�t�B�3���2>n�W������o�^��z|W�Az��x���^-������E����ţ��_�;o��ҼW����ޅ�۾u�}��-?:��������ە~�_Z�����1��>����Q�����=��8�f����o��+�y�o�s�o�>|�k�~6���_o��hޗ4�ǌo־]׃Qo~��}y��o^u�o=��ץ�o��ߗ�ߕ齯mx���ߗ��>ր ��>"�0���XY��>�Z�o�A~->��=��ǵ鷍�WϞ|_M�ۼ��o˾y���ssn��}��*��˛���������ҿ��^�<h��v�-�|^7��_�z�z�;��_D���Z@oџI���/��m6������+�_K��߿5zoj�o����[�_kA�=�^��\�����|W���o>|�o��k����y����j��ݼ>�o�x޿����x��z_[��m�P�@�+�~��4�^���]aG8�nor�O�]�~������ߟ^��߯��+��~_������x������~/��{k����W�_oj�h������W��^7���6��sz~������m��j�����o��}�"D]ļ��z�U���Fu���~��w�QzW�O}~5��7�nU�}^]6�xߍ�}_�~W�}?[x�����oj�����_^���\�w��������hߛ���[}w[���~|��}}<a�\�ڠ�q\&���s[�c�M�n��\�^��_�}/K~/�u�o�Ƽ_�����-�׫���_��i�Kŏ�����������w���~�����nm�W��ϯ�����{����1��D��F����Gye�JKx�}������~�^4o���/M�ۖ�_�����~��j7�/��^�﮷�oj�W�?|���oj�oW�|oj�Z�믵z[�\��uy��^/�g�vd�2�o!�NC� �]��$�jǬ�"��e�ke�d�K������s'e�}ŧ�|m��}���J��K����ޛ��5����^�;oM�����Ž������]��{[��}yצ�_KF�oR[N�eM�M,���ur�6�}Qs�R��o���ϧ߿Cb+�+���ך�{�\��wy�չ�����x��v�|�~����}��u�|��+���~����o������_M�<o�������zx��������2G��s5�6W*�������WXK���X�����l�:!mM��>ƕv�����<rZޛOM�:am���Ð�Ȱ!lu���]Z�P�^��e>@�T��+j��#^ .-=�Nw]g�q.����nm_lə��,٣qY�Q<ؙ�o��e�/!������S'��K(e�Ϳ]{m�ޞ1����oKE������o�������9�|k��o������{_�/{�ߗ�}���{���_�����$2�3�����{�ڡ��ϡ�����,�����ϯ��k�s~�w���o.����W�~z������Ϳ~���x�[����zkr��?���ګ��ߚ/k-��~��_Ͼ�	�C�b#Dy��v|��ur�ʤ2�������������7�Z/�u}+��W+�{�y��^>+��_5�z��/������_޼���okƾ��������������W�6�^�}��签77��տ?����{����6^_SA�W?6L���]7��u�T��{�zY|��/!�[�����齯��{}����5�ڼX��+��o�;���Z��󽽭��m��_wy广�v�{�~?=���Z>C���q�#�c�jI��������޾�m�o����>y��������k�ν-��~��y���^��s�}|�}/�}k��}{�����zU����w[���nZ+�ν���o���[�~��zf!�DxG�9��̔=3ZOҶ,�~������ţx���~��y\�KE|���վ����~W�<޿:�c�������U~/��m�u�{����k~�������r�/k��o{�+���ޕ{{x�(�����+�H�/:�^g�8�2U�U�f�7*d��-�7�����2vJ�x��ڼo�{o����U�ţ~+��������^5{��-��[�{��z��|W����w�5���s\�����ޞ��H�y7�l���]�B߾���U��]��v\^�?�)e��[%�{YKz��%;���szmϫ��5�]��~���_��m�om��o�����}z�\������5�ޗ�G�����_�^>���Ϟ[Ң ��\�b>����y������f�5fv/���2�7�읗����s�~5����hߪ7{�}+ŧ������ߍ��=v��K�oǍ���?|�-�\�m��}���֋{W>��������ֹ����}�'#�zco΍����s���|�^7�n����o�ܴ|��|���oM�ίռokƼ_�~�~/KF�����ח�U��}^�����_���5��W,|_�~�u�����m��;���|�}�U�˟o��F�#�7�<Z�X,�b68���J=�mWὛ��p9=z�I�i�ה�he�v������3�U�̞�9�`��cvL� oi�Ӈf���.Ż*��z�u#qc#̲��6�b"z�t�'���\�k�\~�"Ž��+�������5ﾽ$}}��z�,A|��[�~|��7�nU�����W��nW�����}5�����ok�����}��o�|o��_��_KF������M���w�^oC_���??�~?�����|�}�w\�#>^["�2N��_[ޖJ�����׭x�?V�����{����>v�ן�=[�_KO;���ߍ�o�޾/So��޽-�]�m��^y�Ž��;%)��%/!�����*L_�(Ϗ_���?�_�?~o��_M�x��y���׵�^?�����ʽ��_ߞ�_��Z|�/^o��|[���/?^Z����y�׿�^�������z��~��D���o���T�G�P�}�G���!�)ν;[����_�罽���~���/CQo���ޟ;���k��m�wm���+����zo�����}����n}{����ux�w�~|����5��o�>���ţ~����b4D!">�>���������'��������[�5���v�ήX�^���kүk���;~��o���}yzm���~���^�6���[�����o�ܫ���Ϟ��4nmϫ����}5������#���}Q}V�s��&&V�{����e���A!�=hD`�B$Z/�����o�����_Mp�+��~^v-=��+����oJ��o��������}-����~}�š��߿/���D}��?}�>���}тkԶbK��S�w�ﯟ��ߟ4^��ۛ�~|��w���}�����[�~�}��}+��Z��}��}�5�/}v������-�^w_�Z{�}_�~k齽�����k*0G�����xg��T0���U���߯>~�z�oJ�h.���o^��j�o�>y^�������������/m�^?>u����+���{��_CQor�鷋����_�鹷wm���/����� �$|�|@�ب��\n�U-���~Y�7����ĝ�M�}�5+�oc.o'e�����Z7�����Z����x��|���o�s���y���^���?�������j�\ߍ��uz���z_[�^��n�� �"��%���w�b���w�~|�>_���6�o]}��M7-���߫�x�Ƹ^��߫�x���ޭ��ֹ������[�_�x����j�o�{W��u^}����+���Z�|�R�7�쒆E�ru�&���e��	�׬��<h����N�.%:�4�vb��6�'%�(���0�˥N�)d
�	�X��4f �ˎ:gj��\�������̵O:�v2s�&U���Sΰp��}��M8�(���{������-�E�v�m׸�3z��2�U�n,٥�����v�^�����o�zZ���������^������/M�۟{��ͽ������=��[��m���[��ߍ����������/�Ϟ|[������<Ѿ���kǷ��wg;۰}Sx+��Hum�}">� �� |����|W���o��7�ż~��woK�ѽ��}�ׯ��Z>�y��۾u�+�������o�ߵ���}*��|m���߯��ۖ��}�����K��W���ۚnO�kg�4z�.�q�#�}"'�x��zo���o׳���ۻ��}_Lop�_ݯ��W����ݼ�ֹ��ּ�������Z7ׯ~_�}/�~�ƿ?~�ס�-�ֽ/���/����X��~������ry�:�>��D1|ӟ�����o�ߟ=W�ͻ�r���<���r�߯>w��~k�_M�ە�wW��ƍ���-�x�k�_�w�Qok�x���~-��s/���7ҿU��m�����h���K^�ٟ�x����}���>C����=Z�5��o���J���������_o��*�������5���o�O���_j�h~���|���j�����߭�/M��
�.�7/�;������~���k~�}�}�[�q7���Dh�Q���w�Z��￯[���񿗋�~�yW�����_߿~���h6���ר���^-?���k�~�-��{�=�����o_ݾ�z��:ߪ�W׾��n���s����nF��wފ�I��Fi�} �">����_;���~6�7��ޟ�����"���xDHc�D�]L�w�G�}�p�c��{��&{��+�v����Y{}��P�J�3U@�Y�v����*���ؾW��T�|%Q�W��9Ὧ�y�:�ߛ�q��kq�Dx�t���UUαx4^N`wh�c�Eu��k*��a�;H��3���o)��7��-G�܍�q'	�tW?��*f�͋��N��1嫑f iM�I��B۞�����;�<2%��)�j�󺛱EZ�{�!}��=\_7���J#��H;F�w'v	�Y���"f���{��Wc̥7nWu[N�R(:�/X��rx�+ǵ���:vw-���vrg|�[��u�1:U���&�U�4���{p���J�웭��sb&Pu��ac���yT.{��zj3jg�p�0Q�	��+|s��_��}u�7��lA~V���ȫ��QN�k�����Zf��3���e���l��|��Gy��ג��$\���ٯ���o��Wr8G8&�8 6�qai"�g��ߑ�X�p�ڿ�2�KğL��~��C��9�A��>�u�mm��=�3� �d��륤S���۶����+E���`�Ǧ7o���1p�����Z��q"1�����Vӣu�G��U�0���o��ַ���*2ӨrSs��� h�(2��GJ'�&h��ϱ��-�Eଔ���]�Mu�q�Gh�t�7���i�"�Y<ɣp۠9�{v8Es��4�vLpB�L¡�Smf;v!��a�J��e=�+#f�Uuc��F1���o�垼g�Y#���s�:�B�zp�{K!ZtP�V�
�p�Y����	�����hXbҧ����
d����R�h*�1e��$�n�h'6�^8�{�ҩ�n�b̦s�ي�����Ү����'a뤴�C,��Ib��k���ag,y��Eh
gzFfltf��[a����9"�r�T���N�U�Zzc�ܹ�;"�蜼��嵉�M��J5�̓8�H���X����#rx�s5��[���WP�O�������P�|�{,nN :�g�x+^�D��Y&\���k_[�5�ї�u��3#0�ۋ�Sѡ&�'2|Uu�G��t���]�{�onݍe-m�ȠY��C���W?����d��)��%�5O�V3��8:zC|��ʒҲ��e�n�!񸍙aX,2j#��_k����s³'�u�ah�|I4h68o�;aY�����<Z��A/���j��<�5}��h�L�eYL�<�W���i�؏�b���{�m��3�&�rQ.1���g�!��j�霈�ʔn��Z����r�������x���������lkx1�i�N���R��+�:^�޽J\�,/H�/�'�k�g�sI�Α��s�(��(��[i4���e��J���G2���A.9"�s�U:8�5���-�1e]>;��&���W|��Ư�����<-��CRF���Uk���N�1��}Q�$R9�qGTS��m�W<�4p�Q�v�:!��H-�\l�ݻ;Dq2�ܺFY�����x�g٠��[}��r��}X�v�)Ȣ��-�ݶ��r�3^$\u:�l��p`�Վ���c-�R/���#ӫ��R��o4�0��.u���;�ᔼ��wI�:�'4Ĝ����l(�������z�8�tw@N��<��-�7����u�7�'1���2_@U�R�S2(��n�pGP��4MD��	��:�T��$TYc����+N�2s¤�$����#\�N���a��.t	�+Z0A �i}��}?�k���?avppǝ'�7��D!����K� �\c���8=
�a؅o����n"�����FA���z��YaV캋!'�uI��U1\�k\��#L�����27fEe4T�*D|��+�ހ���%J��]1�{���^9����:�7�u�Y�*�u�+~�?�z9z{���I3�z�:ʭ"KD��vb'���S<�%�Κ�q��6��R�I}^�2�1�I����x����-�_y�7��/��,�ٖ��G"�`�wI��\cu��㺫�����ޚ7�W-ri,Yel�Y^�
��U��:�|����X��
�S�:�%Xz�=�1������˝�{&9�)!�r���"f�G��5pƖ�-�H~�T����י�ؚ����mz�߂��cY�J�i�=X�
���f�*
�O.|��<���9}1�`C��st�����]]���7Qıf��u�,�E�d�*����:*��z�.��XsH(�VƷ�5�z�v�+��ӡB^�1�缎e�]�{
�Iv*J����=��J�T�K����3��N�znjttQ<x"J�A�[t�D��*J��)��ܜ·�����ގ����¹��m�Uv@�5����Y:� =���'uܮח�sz�J0C��l��ucxⶮ(�;�D9�c��@��쌸sH�)�DI�j�k�uvmT��� �2���
��\i����o[�ó�N�1�ޖ�1��16b�e��v���ɧE(�Z+�I��j~T6H��O>�j���Xi����[amYdUNں�/��m\�껽�uɲ<��O8��g#$CSr;"�4�����{�2��\��;�O�K�r�'����Kσ���_X�A� ��_0hymnt��g+���Bc�p��o�����C����Urlc 1_Cr���-���Lt�z�ND����
�[s��fJ��=[wtz���_)��0�'w�:Ӝ�m���~��O�+�k´Q�3�]r��_>�$��}s>�9�W����?��*���{����e�e�e��7S�Y�:��Τ���-�����&�.e���Z��1}��N�E��VmS�e��3�]�N$Wt��/�1�3��Pաyl�J�J�- �r���7���=�
������a�6��y4����rQW�����O��ܣ�}�+����2s��������s�%*la���
����E6�=A�L�pT���*/Z�cR�b1��=�08��B�mck���R�V�ч��M� fW�a�i��N̢���V8��|P���2�)&���12Ok}��w}~�n���?�3�\J�T<O���qWa�H���ED�JG�nl���1���w>Z�e��#��'�󬹇j�@��G|]ΪZǦ�ْ}S�6���Q�uP�:zt|´��3�1�7N�
Ϡ� >�zf� <��jW��v��[&� c����۪f�s�lȜ��g������+�{Z�{%kJ�B{�}�<s��<��X2Z�	'����΂���V��M�ƾ-�9��s����kU��Sj�R�=���{��������W	��!b�#�@�����׬Z2].�Kv=�8��dg�<���v��Ƕ�Yј]ҋ'��y։�|�Qa��z�Du�p{��F�,1�Bo��״6m꬘��v�|[�LXb�%�8��.���u@��F"�~e�0t+�B��4k�J�Y|TBr�r&۩�:9��}e�ܬ��y���M\㌱��L�'���K�FM�����d���"��eu��h���`s���U����#�u��/�Ҹ(G��ug���}ʒ�0�x�\����ٚNȦ�+ ��B��_}���GN�.�lŧ+���*!Q�L9=	��^DL���*�&k��<�����k#v�f=��H>�=��m�����Ӽ��Ԑ��&�J@��=�b�2%٠l��a�X�WED��刯�:���=
��y�����R��oL�v?���T�;UeCj��g�|�f;�]9eN��.��}�f�"줙�6ǅ�Sdk�+�͔�lаťO�6q멍T�Jc~݊����=�i���0��g�y|ٮ�5^���`ܭ��
����E񽝩��
�688�,�2��0��47Y�*��BM\Nd����>���Ec�����n��!��/��a=8 �4�Z�ˮ����������/m6K���栫 ��'ib9�!�n`hc��q�_]ѿ��!�q�,+�Xd�)L�w_1������p�����7�����s���4�i�w��[eÿC��N�8�V�{oᮘ!�ʳ��ed;w����F�=���)0$��� �:�X�6g���̩FQ�#S�>��ä1�A�H��Ň�E��Z���t������n�ۥɃ����LYw#=�vU�U���F�"��m�4�
����Y	dpzںz�P�=9W�Z�]ov��~�������i��(��|u�	L.)�qW�lԦs���`��@�j�d��Xb}f�/F��G �W�z9��
�=1aww��hӍC��s�6�t�=6�2�]ʉ�e�7�ɓ��q�� �iz�9eϔլ]��K�T�'�Lغ5�z�a�6�D�:[��+�Cٺ��r�QX/ŝ��)\��s�q5��H�=�����e^\ɻ[}��45�Ot5�*ca�d�Q���n��t���C�i�r}
e!���z1EWS�Z��u��d��-ԇ�Do����l5��ҩ!X��OF=�o�v�b�K�C�����/��F�g�@c�W�L}'N�4��zN[u$绗ɮC��EV�էE�о2�3 �K0�
/I�ܔ[�+%��)ڰM�q�]���I�ܖ�7(����ѵ���no�nS�3�@��!h�d�OZ�R��{���'<�;��9���i=&Ҵ+ �&n]̳�{�����Wf��V/�]|��m�'C���ǤUĢQn��Z����丹����v����[l>+:Hv��X��)�ɗ�j-�*,!Au5n2�xs���,���3p]��-B��������@5P,K9e<ՑB�f�ĂO`�V��i�!�v��gMl�Ws���x9��w8��1naT�zm��U<��|��nv���E��]�hge�$9o5>Y�˃/��V+��]�s.��_fԓ�T/f����9:�;&�6d�7�>n,�F<�ˤ�3�ƃ����u1u�oM��Wbwm��x�d]�A�F;���cs�h��o�(`�zc���{.�VrY�m|vP6���ٞu�SA1g���{A��(S�^��M��l�Fp�afIa�����1d���5�"^e�!��KY��p�ƶ�LU����➴n(�7d�����Ȝ{u\y&�sJ:�'���z�Ɛ��a��dXd5��^Z.�H�p�c�o�.��F0�����̽]��p;�����|�z�ľC����d=�����g�]�U�kt����]��[\:�.�`��t/[�{�O&&�m�q��޸��^�>�ϻ�HRmt��S�rCZ �1�g'^��8�tf�\*I��Ax/����xq��25|�E��Wb�xc���+�w������Y -���yW�n�Aw��u����v�M�����}��H`�����s'hf�\)F-�!Os�`�b8�z�e�B���77�_b������+���ig��ny�㶐�kp�������*S�+��E"��u���f����r����+[z��J����03$�f 7�ݸ ���P=��u��ٺc�C~}r�˔浔'��O�߿_���~������t܂��Hn\�H�Q�1�$&.;��`���n�đ�H�d�P)�2E��d9�B� �!I�d��8���:\���r�	�1�c(ҹp;����a4M�HM��!w]\�tJG-��N�";�&(F)�"Tw;qJf�Gw#!4�g"��\�4�fHH�.WH�RBd�;����ݺ���Xi��(�)�[����Hd�� ��&�$���\�f���& 0PfE��ن�M�vDTd� �$P�ILL��d$4���ta�+��"S�!)��bR@�$���3I) BĂI]ܖ#"TD�HwnQ2PiN렀;�7]І;�r�&ġ�����~~���Uz5,�Z��K��WT&��|m�+���D)�n���/*�eQŻ�ݎ�����,'����::�M}U��_j���{d^���Ꞇ�C
���$�}Ps�3	��Q.�����.P�tK�������T�Gh��ڋ������isE��Hu�}��_X����.��Sݎ�6��9�Hq�%�r������S�J���P��L�5� �L>צ���
�H�,����+vH��KxW���G��^:���ot�4�ydh��.�o��n�$��1i ��xE}�+���ҙ�<LeG.�FӘ�\6�yV�^^A�}yl��On�R�Đ�Y��A��Q�`�H貇i��:��!̽�[;�F�yxկ��g�j�ɍ�2$��6:
Xpd5?��'܅MyJ���:�U_ �,����o�<W�)��P3M�KF���,�ѓ�%�a�(C��w)��ن��*�M^�q�W��=f����Z�A�Y�t�1"~�u"+
' X��Wg?F{��\�t�:��.Lp��n�3{���D������˘�TDu��ٯ���jo�c�v�#ÓT��5�@�g*����V�����b����h����D���۞�8��9���P�u[�	�H���o)�*�шG�n��uuw6i镼��;��':�<���5�+�f�u�%,9�8_��W+"�
'�&�j)�d6�?�$���w�b����Ǧ����Q�W�t�,��]Kb'��U{k�������n�,8�Ӄ��jT�.��)_���5�-m^g�i���y�A�͙`+��G"�`�t��eE�X!?����J8�$Ef��A[T���Я
�tW�a�G���=u������I��&�K�a������ZY<!�<�g���3|aụ�`ك�e|V����C�e�e�u;�#���̗�U�9���Fk��3��;�鹇���K�B�@��M�-V�oܘ��e1y���g�z#��%���?���r�� ,6�HĪ�T� ��z��ȑ��w'Rj�7w굔��
��hg�m\Q,w�3v�����b��o���z�S��x�����%}`�j�ʒ.%��Ti�����\�O�=¤giG:�S�hrθ�/C��gg�2���⃪ԏ�~����O>��Z�cr )a����]l �^�stPu�9���\r_eVr8Y1h�*��Թs���̠�o�[f�#�ȹAXd޿*�dլn;yO����Ă���^�OYMЏ���"po��YJ��M�v���3/'۴�sd�/|׀:��:���n��flm^2�5�g<ǋ39����W,���{l��.��b��zw�v[M����Z�'>�8�/�Ͼ�����-�[�y4r��響D4����偯 W���A<Q8�C�Ϗ�ӥ��h��Cv��[1d�j�F���WE.ylbj�M�1��健�[V/���'��� ���DT����0��2@��M��B 訃����4V���� 9��}}�	Xzҿ{s�E�zƝk6���;��Ũ.|-}�G֌;�9��~����fW��S��ß����+�˰��}��|oC�lB����k�!j�Jj�������q�kYc�W@��3��
���.�9ʭ��Lfb�k���p��*�}�<-���T�~"/[��vN$���p��':|�����?�����BUud�8�t+� �]+�FS߂}ڼU�{d�]��crE}jSs�򘎸m����׹"�NH��ޮ�	�Z�W&���L?znT�����q5�랧�G�+yQ��t��ț�`�1e�v���E���M�SkA%8��!9��u�3g��44&�+|r9�gE��e��/���?�fG��^�2]\�h����D2q��!U�z�A�\Tz�g�҃CZ�p
0w�k�՛�Ahm�U���&�\Y���]uXkUn�9�T>��b�]�;��/*� �[[����Ȱn
G�P���<5h+f��ċ[*�Yz���b��eO��1_{���^�mi���6,����<j!A�%�?@��f��G��V�-��6tXs�i��E��C�؋��\b�̶7�=-���[	49�&f̴t�qm�Xgk�yh�"��&y|��3c�`\ʫ���nxn7]������bY���@J��11<����{km�ܾ*D��9���8����5h�
5��'�])�G!1��n2;`��{�嬄gcy�
ۣ�w���1O���J��M��t�. !`)�&o����+�Ƅ�qk�DL�k�^]�C�}A=W���7�+��{\&�Xy�G�t<���T��ԗ�6�Nr�X������厸׏��<����Q�Us����W�>��ь}?9"�&be�:u$�S�m��?Wl�tzʇ4��E]��(��<62:�i1y���"�滫W�Ek��r�2Um�?��ac���M	�D�4.����U\]E���310*�I:5�ݻ�e�.�-�g�ތ�g�E������v�X�l-��wo�!5;���j��{)A��Ffb�1�u|�{y�"�lo.�@��kr���]�7����f�Z�l������?�3���)ec�S�t8y^iko��1+�T�&Wm�-�}Zq�1dR�2\�@&;Ý�[�f#������>|����ORv���vC�<f{��0���H�s�n~ǳ|�K��ۢ�`���z���Vb�R���s7�G����
��f`��3��Ͳ����)����5���4}��g:�l:�ۅv�)j�ݓ�ڒL �\	���L\GZ�&+�N�V5�����9L��;fU�u�S<�u�����(��$ep
�k~9�mq��0]gzxDqx�i(���Z�.�(c�M:�o�O�+F�v�+�_��ԫ����Q.��S�*����:--�� �BÆ��1��F���J�[�P>��a	��i2�����5w��+�Xo��
���n%��Ծ9��&��n���#�� q��fN�m�^���댣��z�6:���C^��1��.�q�[¾��"�	�l���yS���9z����9�F�+K59��� I�Le	d>�mv�x��S~���'�\�b๶K�Up�9�wHڻ&Co7���5 i�3!�`��W�F��P�1wJ�ju!��d���}�YCRw�cO�va���۽�� I��'^{���/��~#�g��7J�9j�=/��=e��}׌M��^G�w,�f]u�����$m�� ٸ�����v�3�)8�wY�aqR�Vrf�Un)��ωBS$k�E�5�Ά����U�U}T5�J��숬��s�y)�ſH�Tz鋳+�0\e*zk>:�e��j�v�Q}Q\2ָ]�? ���6X
f�9`I��zo_C�o����n"���=P���x�)Qw������p����c~J��N�CqK�KB\'k�we>�A�6k�7�߮��;����<~�Q�0\v�gv��_��N�h�;�9q��Tw�����&�jv��1wH{i=jw�X�r����J*"�s�4��'��y
��dċg��b�2�Y�;S�7�{Μ�:x�GY�+��p�̱�&~�ڧgFA�A�͙`+��EG)L�F��/r�XU;m&UW$yn�.6��1�:�4��ˡ^�ep��XxJ
c�Y]XM���Z��0$A�/k��}�Ч�6���>�3|b�vT�B �Ϗə�=H^�WS�]�w���"�	.��~���v!`Mތ��e���{p�������is�Ǉ�J{�����Z�^�1�:�"�]ĳ!��JT��!����Iʫ�I��}Y���̷����ׯ�=i��?x�pS�J,˦�ۨk��9z��a���?H�x��������Z���V֠�5ĭw��	�poN�2�8݋י�ϵ��|�_��Y[ˮ$A";�8��z��@��G��dt��Z�>�������X��Y�v ��R05V����V7�}I����X�6�a�Ӊ���s��A�'��N��8W2O)�DK�u*�)O��L�P�F7�-���>�c�6clU�5�zf�k�s���7�A�UHȯ��JnOʆ�'�M��P��,5�|~��-¦2����y�U֌�e��b�*�:���	�л�;��d�����L���dˎ�3���O+W�+�rw!�꟪9*d�e��@��	N����܀d-!�â5��Y�b�ԭ��-4��w0����p�R��&���2ܰ4�j�:?,��՛0�3���^e$�a���=A��l�s�wS���Xn����й����?mCyv9�鷓��{�jm���V��6P��������L	��Q�?p�)��l��~��w��m͉ng?w=�<�F�}ڸmTl�p1�qfr~�<Y9}���ֲ���Ν�p�NȖ+%��犫z�'4���pn���M;���q�.��W��n'd.@x	F��T>�t�>��I9�C/�������2�He9��9x C��èw�Q�q��t���r��|�Tٞ�Ϋ���\Q'I����N}ڄ�-e�*�'[B�?{y����p��V�� s�I<h��w�=m`�n���rU�ﾪ�""2lo&���'����w�T����Qke���&�k����i�eF'G@V̱[�-,�%���Dqwc끍��nuC�b:�W4����H\���Nq��b�Syw��[�p���V�X��!V����gGYJ�sr���
�L�cq[z�ƶ�&X�P��ʭb�݇�]�)��N�̳ud�h��n`�����9�C/����1�A��3��v�ʰ{�^���x��D�:y���)�1Uk2��x�x`�V+sT+g1�I��v���#��c�0�*�S�F!�2�3��5�v�f����ڤ��̹����e�Zw��졸�f�Wt��I��:Z&��f�E��Ή��oN��q�}�����S�Z���v��ɫC �H���5�n�x�&��f:�Fű�����J)5�=�wq�}]F��Ց��b��|�5���L��ªRg/!���E嬷'Sܒ#h��!�*~ggƃGh�t�7���i��+�̚6۠9�[��Ӯ�᫲$T��_Iɸ����,Sp��:��Q�b<6le2�r�M�H��Wq�R���`{���ƫ�Q[�jZ�������9tvؒҥO�u�,��(Y�LN5y��g�����&�҅T�.�f�Su�N챫�vN��7c�*
�LE�l7=~y$��]y��moa7!ߘ)����}osCm$��S��4P��뎷��'f݇.��$��9>�d�r��{g��6v#��.at���Ã�N��(:��2$Ta�q���P�(H��S�|�q�����U��<���B����LUfu��1ר�f~�WA^S�JsO�րz���e�c׷�8S�熻)z�����v��>�ܡ�aE'Oc�)7'VZ;]��t=���� KD�@���8�s�n~ǳq�碦Ł��hҮ�	-N����O�7z,(���,�u�|�9�U{�ļ:��G�Z�_�u���n�l��崥'�9Hz��GD��4���T����Q�֨I�N~\5��Xc�w+]/��T�W��&w�g���U�n� �<�
���dK��T���}׳�X���%�ֵPY9�|�æ3����3l�Q�p��=�e �9�j�ewҗ��o#	��mjP��b]So�o�r��<��k"�qc��J������������
�E������L���X��.�-���K4������n�>���κcY�+騣Yn"n�\9�F����]��=�f�~irݴ�n.3�:H�u�w�U������_3;TQwW-�]�h<o��e���=�]����K���Yw͘��͙��$�wK�����Ė�8R��N�q7� �uHK��<����t1�ڕ�Wm�m݀8׾��ī�ۿ8�������ѺR.pCg ���Mށ8���tM�F�����'ID>�(0�x�Q����߇Jf��1�u9=	�p�!�M��,2x�e��4�nfy⹤����HBZ&��u���>��v�&�X��/]Hd����p*/��k�Y��9T2L=[�A�%\����G�C!5?�"���/)S�X�{�s�����Sە��X�{�_`p���h��D',	5N��=��:���|a��Y���ә�/ak�ˢ��ݑ�hh��VX�J�����4���Y��dE����uU'hiE�ŝ����qս��R�7L�ݾ�3�C�3'_4o���u��T:����yV���F��l0����&t�<���D�>�x���N
�c(c�u�����l���������Շ[�lܤ�]�ϫ�8�=˫�(c�
*��+�y�6��iHN�Wq��X�ٸvoZҠg��N'E��1�W��C�s*1��ܘ��uGy�:�h��lk��oV�΁L��Ek�o8�ї��iLΘBK�![z��7�Gu�����rX�ufi�j�^1N�ە{2ڷ�[�k�L�)el�E]6g]3�7�r�Vs�`�5#��H����2�q��;#2g��Cg�j�7��N���j����=@�%��s݊�.��хl��M>��kmR� ��ͮ�*���.=uPr_'�َ �7J���9ҵu~�j�5����@ \S\�m[�Y�M\�V�Mj�v��$���y�wf�:��l\�6*��Z����km�vP���J��t8h����"P����_���n?�b鹷;p���a��
��� �ͪ���};��D3K6^��6�vL�]jv�1+D˾�D_U�~�W˱�7\U��o�` ��C�ǔ,-�%�I�II��8�\�&�����*5�w��r+�>7w�Ǚ�i_ggP�u��[g}4����TE	�h��:`x7�a�h���ӻ�W���r�K��e�;�7��3H�9G��[ӕ��I��[�ə ��P����o^l{�N��sC�������ϱ�ڇ)9�u�ֆ�W5���y��mb����G!�&�>y�`A�ڜ����Y�<��4y{��H�L��G���Q��C�+]���QCyX�C�����l2��t�t�4������MJ��R���s��&������V�|��Нٲp6���6��Mb;�:�v�ɝ������t{:\ 8�(��WX�C��$�N^�y^6�/L'f�P�[�w�^sS y*���g^Cѕ-�=u��SOe�k3/h�*g.�}Ԙ��_`��H���j*��=n�٩F\]_��Q�Qc�*Y�I�Y���2��f�]�W��l]n�J��\"���;���.R���GGٸ�T�Ǝ��z7�����@#6n�ܓ�Z��%ҝ}�x*Uɔ���e���oAr���v �}p�� n�^Ű�1U���g�"m�Ⱥ����U�y�WU�v)2�r�� �����e��AXNU-rb�Rݢ�ePK'E��2�\��y)��`๦��CIG�7jȴ�[���Ͳ���#z�k:�yx�����M�d�T��j��p�X\L�A�&滧Թ�.��A#h.���{��P�����czh���c�Bc](1;�����%,�#���uh�yH�o����%����uS��Ty�������ݧ�uM���bC5�[+fQ5����,��*��X=��W�{P�Ƞd۽� ��ck1>ۜ����"�y��v)�6óo�/ln񼓾YR���1ep%�@-յW��j=Q-m,��GJ׌�j�`P�kiu�خ�ӽP��(ݻ�'����z��>��� 
C�2CcE"�\�J���t$� ,�H�̢&C0��F"-�v���4��&���(����0B�FIF��1wt�N�@f#$��Q"�3�HI���L��&�@�0`"I!ː��Iu�d�Ja��
d�"H	(��"K1�8IM��	"$PH33%3A)�XF�ۥݺ`Y�@( �L�)#0̌F�2Y�	(LB*F��$�Hf1��Fd2!�B��#�B��B
L3$���1��D�`3M;�0� 4�u
I�&RlE�٘ƒ��EI �UP�@ (PDݡw����;��N��P���2��}d�s�lv9t�R8OdHm+�o�o�_�j�M�,���e-���@�]���W�U}�ԇM��]5��@��u�����8�FBQ�.�҅���TFҠ�=�8��j71�����+f���K����ä!q�^��1�)8([���2�=�:C&���M-��sV�����
�3�.5��]��O;�8�z5��-Dc��w���������=��5!A�n��qP���_e�E�ˮ�Y����*xs��cn1�M��#o�U�ީ�f�'1w��;�q�;	��\������*��L$V)��e>��2�q�3v�����Ǚ�َ��K�V��N#f����d'�����x�ZʰŮl�;��
Y��l��^i#����I���\�M��uLȥ2R�5?*�l�G>�Ja�P��h� T�]\�6�Vܟ�����2>�ڲ��V}
T'���p��:S>P��nr�[��Ωt�ո�î��%�T�������}S�}�S%�,y���"/�'j N��閡�u��@��=T��q�q/�i�ۘ�y�E.yld&���d)�`iymX�G�E��rʍ쫘�ю���]�.��`�0�5ٜ�n�Gp�Jv�D�]�W��ף�e��q���St�y��[���Ȧ(^����������-�r�uth�=6����`��b1��0�!m�zץ�� Į�%T�̹K��j�����w-5���^������vk_lbk��s�[5�j��A��e;�k��]��΀t�6���0(r�@�;�z��MV!�=U�1+�F�+B���e_sQ�чzs;��g��y
C�P��J5����}��1=��5��a�`�cATxZ��OM�S�pN%��Ԍ���[t^
��35BW\!�Y����Z�M;����%�U��i�t�h4�mQ��5��>�eںw.�v�2���n������7�tWٹS����j���'/e��K�r�r[6�����#\B�&�o��8����nH��Jn{bS��Ϋ��7_Lv�H�Ӎ����oދ�M�o�vI���.���ơ��v1+�X9�ӟi�����3�1�c�h'#r۝�Ƃ4P����'Z�]>��������J��!���ʉ4�o1R�:�}���ķ>�/�}q��&�P(9'�P���f�L�~��U��7_Yt�����`��n>�*l���=v�ߣ��=>����*�\�;@�>d*�k���2{��ue%Z�k١���n:�\Np��ʳ52�xN�B�Q5C7d��B C�މg+,����qf�'ьˎ����n$�+'HJ�ܝ��7�{��Zr��<uAt{wd|�o���۾=�Ƿ.�b�EA��5�Nvg�'�Z�T�3`oz#��>������M�ȏbUÁMTC��Ӯ�n#�:lK?!��	P�'甖�#��ef���r��=F8n?���.�EG&�-�&. 1aPۭۨ�0Y���瘛9x��>XY� �OQιH�dr����Te�d�ɺ�^L��EE���܉��Ƿ���@ʓ/%��5�����Q��<�&t�����|�ϯ�҅��V8z���z{����>1d���飒��PRz���e-�+L,=�����S�"�M�l�ĺ�e�Un���&:���*�c�+͎��q
�l]FƾXMK����9�>�L�o�:�[�hXa9{q˝0�W�k�ʱC��٫4.��t�P���Ͻ��s��%N�(K�%�:8���@
�qT0�g��Q��9��sv~���H��D�9r]o]��'uKA�qY��c�����y<��_�D�	� ��\�FB��ɷ?cٿ���s�����u��m��V��ɉj
i��1n��zf	Y.�iaͩ��/��_k���Ȉ�{���Y�L<�Nm�;롽�)��e�Ǯ�Urޮ� ��,k�[�kt�:#��U
a�m���싞9���nkGv�d
���U(��i�%c�������}2'�FX���8�j�@I�\�{��	��z��<�n�Yޘ���/Pb��������o���i#�a�ź���o.SF�*D�����5Z�k/���C<�
���#PR�6;���T_��Y�d4���GM��A�Ep<+����?۶���o62�J���GV�������̂�GjW��?P�'�$�+���䀪�:u���̫����܎�ǽz��1����j}����lI	dd,P>o-���b���|Q�����(����O�;�O�&廎]���uÉ��0S�Bof�;���nluU`�y���4T�@b~xH݋bl}îӌ��f��s�.�^Vwf�;��P��O����=f��Y��;s�-fo��)���w���-�� ە�X���'�ɵ�Y"����=�� ����*�U��v.U�������Zr�;f�Y��]�سs�'҅I����FӔ��&�U
ߤf���k\1�#qԵ�3!��O�� �<�cn_ZSw�~�N�E��L�',	5N�]ԃ����WE0%S�/K37���x]�[̻��D�և��%\-[82o��pɤZIEޗ|�a�����&ZMt�u���x��m���ێw��ͳ7��@�x#u��>�'}҅�]f�8^�*��j�c��7[����eZm�Q�lU�7T��b���{�<���gx�T�߫rD��8}n�!�x%2�r�A�X�,5�H�S"���Lz���(�yv$�u{e�K)��op��#v�f�o���2^�����G;�8�����]�+�6�W_�<=�遦�1B�#|Sm���$�σJ-Ҙ���>U\�%ha��J�z��-�*���ӎ5������VcDs�f�\-�K�ļ����r�|zF�}�W}�C��ӆ�R��d����2�F
�V�`�Q,Q��d!��}(\
���y��}ܷ��	���#?����4��
��:B-9l�;����數2�=�)��*��#Ϋ���wR����bC��.�v�y���R��W�������wU�9I�Y�����f�PǗ&�Ǯc8�޻�f�����Ϲ�f6��M��#tI'g�-��vЫ#>� �;P� ��D�#F�H���o����L��Y0�aq���.3������]w`R�پ�\�O�>H[@i����	w?�i���\)��d��ڢ����:fu�*�!�\�]�I��j�C�{���[�t��N<zE��'3{��XQ^��cy�ë`}�/����JI��H���]\��9�\;^����Y�x���ȤL��h@�nwnXl�-·��0w����i��]L�-2�9�z��7����NJǽ�[�lN���R.c&��fEB�)H���$L�}4:��Ml�&o��TI}�4;eeq�od�kR;�N)����u������T�Ez.�{��їG�/<z.�0ˎK�P�-\����W!�}3��T�y�r�ׂ��&�"&8�w�q^�A�+vaC�/���L�#�B-��4wna��͸B*5<�3��\��W��K���M+��m�ͭi��l�4��>lo�a�w��?3��N���uܝV��΀t��dM�s�p�kw�>���%���.A>��J��k�hUF.����.l}�麬��;������]^!=44�j�v�����S�E5U�k4��RĐ��U�*)���BL�pWBꩈ �<�%�Ŷ�i�;3nn�\1�Y���GV�Ǖ:m2��!0!�C.W�;��E9�e�"�Q�_�kh,`@M�fB����R8��ۦ�Ί�ܩ�qe�Vkn�d���t�_�ı����r��v>�ܑ_Z�����b:��pcr"n��O+o/�-Y��̳�fG3��t�]�gaV��WLN�Y�;�^A�����޺-$�*q޾٫g9Hx7W���ղ��P�6�,��1������Z�ӟ��8�`�poM�g�jλ�z�yz�ZR���Jؘ3qN�JL��Y��)v�=��{��Gn�ۚ��غ�m��� h���ژrtB��+�X9�ӑ��9^5�y�l���͋������ֲ�!�n��ɉ��'I@\�
rb4\�8]ó��v{z2,{B�X�w�ޥ�V_�~Cj-���*���] @GfwL�~��Uk1��T,���;�v���?�0[Z�#̌;�����Yjp�V!�2��[`����#U��V�u>��I�c��2]m.���;��Ʈ^ތ����Qb8�h�r���Z�v�<qw+|k\s�.;�5�5[�P��xmri_���Я�y�X=��b�>��t����4/U���V�����7��|����o���<n�gG)k��w.9�L8�d�h���X[��E�=���4Ԝ�:��ކ��a>���\�޿L�/8�O���z���;���۷���)Y��u̝���Ԟ�����zuJp�W[�^88��[��땼����k8ov�4ړPBR3m�3˷8,G�9/[��[��H�s�@9�_t��,9�N]u��/8Xŋfw��Eu�ۮ��@�S��Y�}v�o���au��u�5YV�:j���r*g`�O0��ٚ�����Y}�J��UW�}��']R����
�Kەnҗ��-q�gϨ�F\�W�`絖���xfLqN��v+������e�ڢr�;S/YO_kĽM<���;2�{N��'�Q���ݏ�g3�?�l�	lu�Q1ع��\ظu�n#���N�0��p��n&�rH��<�B����ө�P�ip�6+�oo�x�W��q��uuI�>�����Yj�?p5\mK��PUF'K��X��/o�d�O�#��򆱴�:Oo�[�G�)�|�^���ս9�;���c��3�/�M�j�8[P�z%��C���C��^3��}<!
iFO��5����\�K-�e'�����o�TB���Ag��;=�wIQ\5��e��#�E}y����#��Oq�{���lel�T��ej���8�B</�8����#�P����ɥ��`T*t��&������3I��y1��[	�d��F�qP���ʀZt�Zf¦�9څv�6����c=C;�Qzx�M�%3�{'R�2�y$���e�JE{�M�"�_e�)X��Om�;̬��xku��t l��4���ZY�y��\��}����W�_x�Gt��\8tf���<o�� ��]K�r'Q~�u;��^��6�U��i��Op[�����;a�W��n·XZ�.�l�:a��b=��-����$�T'�5�1)���dLk�'�ص�ʱUa�X�G&�im�/1��:,*/|�O΍B�
jpv�ʨ�dN��*�@]5�4��2�o5�h�[���VeGS����[�����ÕC�;N��57����U4�9��te�}�$[q��=蕃*;S��+�����'�X�n��gs5���bFbW���=�x��-9��]�����b��υ�ѢH�Hn<7<�,W�u���5�t��x|Bڞ������m�P�	Ύ]wvwv��[5�_1M����=�]�j�ol�}H>����uS�ݽU8o*�gV�m�ﲥî�����]o���<�Ntv��@m��Bz����0�{��*L�/Vs)�o��͔�S��.�)����S� ��oN���N5�qW�5��L�y�cd�����ky���Fo�Ӫ�p�ն��^�[`N,(�pe<���t,�L���Ҳ�5Oݫ�6W��W�}q�r��kr�*vU��e�o�[ˌp�c���z'xʝ%�tn��O�>\�/�'`��[R�ϕ�u-�)<���[x�j���]��707�^�!8w���]%|�RW�z�>!���2�v�� ��w��n y�<ק�M��Z�r����������)�C9n����"E��;Z��U�-7��`M��,�!u@�� h�w�[�x!��v�ao[�a_.�pu��G.j��h+�T�<Q���(��]����z����qe���Y;��}�u�T�L4�p�1: �R�D�N�e�hNĎpڀ�~/s.#)���5mF���MQ����n5��.n�L�[�^.��[d��&9��������/2����X�*��N��F�exl�����\u�͔��������i��U���<>[��y�O�*�x.YisQۛb����1�l,b�ͼ�dj���{@�\�u�!��%Ц�7�n��i 5��tfnS���u�%�nD{gyԦ�2w���������RUO��)�ef5|��r�N���Xi�,�ؘ����71s�3(=u��̥��WK��|��5�/�D�Hr��䋍^�)8�>���[����D�"��*�3*ˊ,vM�ח&�.��u���!�m�����4nƏ([E��jmotv���H��(0ⱚš��{U��w<���:7(�J��'����^�w����3[�n��#�V�f�]-�msڋgi�Ց��A�I�r��Fqa����`�=��z��-X�2P�Z9�88�F�%ϝ�aZ���a�V��rH��g��m�������q��=bcU(SW�)�fK҂�P�����}�хX�b�F��n�8XV����Wn)`��xO;����:oi�ҩ�	�E*���R�ڢ��y����5�qs|�[:)�Zzo�hٸiY�7����ja9m�g���^��~�e���JX���	ku����0;p�������J��t7Dڹ�#���<瘗H����6y��B�h�Tx
w�"Zrf�5�Νv)w!��_g_�`y��M�E,�l�(���gU��WbJ��G]1L,ٜu���� h�g6�����wYJ�
�Mx˧��{�`CS���Y�:�(TI#r����U�G��L.���BnT	�ƻ����*����>��W�u11p�{]�{>������h��e�P8Gݗ:�7��G�w����Y�5S��yl"�NZ�w%��/g�ʖwv��+���Mhy�th��i���ٷ��n�ʙ.\�KBu�� Є�yW�(e���K��U�V�(����w .�:`�cϱ	�xt�F��f2�&F��vb�@Kr��,^l�h4�T܇��|����C2����*F���+N��+��F�j����j��mf��w�_�q�U��&1��[�:�ޣ [epZ=�]P����=!Yo(�Ÿ�����7D��H����\��z˩�BK��;�}9i�\���9��+i�L���u �f���.�C�?�n�}�]j]�3y
mV�b+љ5���N����fU�\��t4ML�"�9#��v���s�C�<��2W<5��|I�Qv�_1κ1�k,�R
�5n���-���>.�q��P�;���^�H��$�Xzn��PK`��5��^X�����R�T�rymn>�V@M�J����t&7>�|���j �����(��`1kC�̔:E�K9�ٶ��]�jI�����M��yXr�S)��`;�思���oZXn�*9Q��b����8pن����n�(��o�W;POO�cm��B\�?�|��Ͽ_�]��ׯf f��A��\L̓���ƻ������B��\��Α(4'v��p����9�Li�s����@!�DD�#"0����PD���E��0�&R�B�$X�%;�LHPQD�Fs��M���)�e��%��� �h�h仹&guЧ8,F$"l�n����D�S1��2#0�4�&"�,A3K��,bDɴFLGwI�l�L��F@Ԙ��F��c$D�k��h0�Fa��Ȉ�u�&)%�2 K�ą)�A;���1DL����Δ���J�I��cI�D�BA-�sFD7u�29y޲k�'�ü͞(o�%���r�XSi��#�W	C7�L���ˮ�N*l��7Wn���]�;�ƭ�hS�E�D}�C��SǞ�}���L���sO�)�+*x���-�����B7�����:�̱]�+;S<��Z����y��~�im7Ûg����_5�nfs�����F(���̩��t��ʹ���b��l���3n>S�VZ~�p1�ҩ���%q�Ҹش���>s�0�%]-nRu��)"{(��� �ڗ;*
،J�����5��5j�`�Loq[<�jT�6���5�B�LsB����VԤ��u��G^Tރ�]�����k�rmk�p��8[Qo��Kb����W��ޔ�^��*�њ��vr�h�ip��\sֻ>��m��)T
���,��5���.�EZ6�˰8e�̆w�>�-�p���D[c+�,�ȅᔶ��S�e+*~�q/���߻��i��1r�_G&���;��
��}}:_�1�ʱs݊h�x�Y�u!��1�@,������s�r���~M����f�ާׄ�e�������ð{
ֳ����Խ�r��,bt�δb�F�'�I�'��db�L"Gwg3mҾ�12����mS�7� ���K^z>���P��in��>�ʨ��p^����7��t�����o��1��E��<�Λ(�_ǐ	�Մ��anNE�=���9�F-��申J�g+�V�4��w�YU�ȞC��v:��Ωm۷�������s�,ǉGf[�U�i:����7�Q�ޱ�Kzb�1L�f�z��g�;�=�m��ތ�ټ��ʷiK�1�}Gk��F��-��Nz۪ؗH�r�����sE����"���W��x�g�ޞ��I1y��<�.���J$Or��x�N/ Jc�(��\�®l\:Ǹa]P{nu�5Y�z�g�;=O^�d6߇[��`��u;*���Tl1��"Tu)Ɲ';��ė8�|��fk����H��ul�9����T�)O���+j����[���O��{f�c��JB�~�s�yݥyH�7à�Y���Y�|�Ng��^|מ �i���,f��������]�Cybg�y<O%��̀���t�hf�-u*��jٹ�F)��g>^�[l=�o�n��q�9� �Q����zk�y��ݵz�콻�Un�7銆uڬ�}��g)ڦ�C�}�7�vQ�'57����k��ۈ4�H���IC�nmK�����]��5��-��zv
O/�5���_)I%�@�������b��X('�S�P`7�G5}ob|z}��v�q=Я*�3�g��ٞ��vV�Е�N���|��Z/J��;Է��iV�L�LS���5�P8�f�y�7p唈]P%*�k�v�DM@��W�q��c�f��4��3M�0�t�ˉU�1|����y&&�=N?�3U�]ے�%��|�T�$Ħ�@J��Y����91�`��R
(_���n�w�̝��[�io'F�8S_&��5�_k�6�w��&e9ͺwM3�)��=�-��~����/O�wg����؞�ΪCz�&X���[��p�Z����C1TD��+�v�_nW4K�@�6Ӣ3� "�U����Y���Ӳ����tz!w�̵�]�D��e�w4��!ȭ��]��V�Z��{})׺q6��zmɛ�M[�_;�D-��n��8�.�zھXW,�kR�{�#߮�����	�I!ӏ	Mf�c5�R}G�P��}����n���v[~Os?W��%���1����*���+c'��Vda��x3�Gx���E��}����!��|Bڞ�������k��k;i;��+n�*3��T*����I�n��=��z/l�E ����:��y5{=�cY8���]��z^�CZ��b��e�m�îz's��@p��#WʞE����X�;j��U�yt�d<R��qo/5��8[_&���ճ�)�>y�#@O?���
(>[%%��ޝ)<�pֺ=2갗J�;��
�����|�et�_
�>ϊ�b���o\�Śռ����>����͵��gU�2�r�w���Rѡ5k*��[����UΣroy9�_b�)�z�|`�M�e����JUC� Ks/�.�(r�%ܲ�®]�6�����5q��n�m��N��u��^J)��fg�A�)-Bj0y��rn�J�[�t%_�I�Lg��& /v*�`�!ԧ΢=佮����߆p���<VWX}�p���6.Qi�9|��WBv�|(H�D�I4y�d����3J��o9��i+יm��QVL�G�ꪩ�zӝ�b������r�'{��֋�����a��c���씭�5S4�T�җ?t��S�����ÕC�#T�y�|�S�i�+)�;p����w�P�r��IX}W�_�Z�g�գ6��,��>s����9h�Z7g]���}66;�v��j�{gj��f���k�f*�m�Du'oj�r_>/�����3��ƻ19ԹϺhz�ϧw�֖���3����>��d3|��T�9�����s�3͇8ܯ{[?4����N��l3�{v�U�SEV�)�9� k�g0J��M��mW6.7�
�v��B��3�*�+L�n������w������uW�N�eBX��cb�or���u�]�۫Y:�y���%[.�����^�ԥTk('�`2��aN�_odwU���OnoD�����[R�ϸ��9\n��������)�.���Օֻl�r����**��n"��Ҹ,���,nE���5�:N�7�e=�'�ݛY�i�!���woWg4S����|}�_x�����R
y-ŏ�+�:J�)����Jܦ�b�ɭ����=!�L>k6��d�Շu�ܬ5ܳ�᭸�k�|�JQ#��|�xx�	G��ҷ��*��{R'�oV�����_e�ֻ>��m��r�HW�tVZ|��陫X�]Vq����Zx�u���i_�ޭ��EE�2��9حem��itbq�檆���<�b�ߪ�)l�m.{����3c�J��p��w;�p�Cs�t蹘�m�:x��CA+}5Իf����!�˙��\*w).o���0�g\q0�<��)�U�8��<2s/852��z���[��5o6�7ʍ|󘚆�k�s���C�Zګ��ȖM�]�-��c�y�����'���\G']-p�ロ��7Z�O�zx�j9���u6�~��x�.F}X�lm=��\�iK�1��8��چ��#]L�i%��18;����{_	x2�9D�w�)�����\�1݋�;��H�g"�3u_`���}��(�C���u��|unWe$LyLT��1�.�p}��;9%)^��&���^?=��x�r}2�\���nh������*ekSEڜ<�[�C�<l��L����^v��:��p^l��O��~u<�k�ZH�.�u�3(����ʁ)��Q���Sͅi@-Ղ�֫33�a�>���^Qd-�_��ո�ْ�ꆮ#K�Y1+�[��%8�5���sZ�=s����^�ʊ@l�s�:�6��V�u����)���Lz�+�ثp�&��t������ 6J�� 
츕���ο:s��1{ꛏ!���nwh�M�j��cM=��5P(t�@�mq)��l���]���_oi���Z�,��b
O.9�]��6���	���A��޷
�F�-|�Q��Zy��z�1>T=�+��J<$^�L�����:4?������D)��)�Z*#J瘎ͮr�Vf�1�+<��C���b���<��&�+�L�d	J4YO��vf���:�[�՚A]yGr��m�|�o��H&����n|:{cn�����W��]���;�N$w�Q#'=]@Ir�����P������&��y���ļ�aG�2vvڶvΖ�<��0���u`�V�]4���*�m��}+w��"�l��o.� ��n�n�쨳2F�V����[��7�-�|Q�m�*V-b���(��^�w��ڟ*kf��֦]7�5�I��qdLk�'���dL�l�j���wZެv���9ٗI��њ��UZ�N�,p��7j�̑n�n�r"Śjur	_F���-�Jmg�ڛ��|��z|k�<�sp�j����gj�-[�\����s�F���@�t3��U��Sܞt���|��)U�H2���X�����#���y1���U�n���~�j+ao�jpv�����]5���jT8�f��61־���$�ψ[=ih�V�^W��]�e��x'&������	�}aq�1�Q�6-�l���W������P��H��������J5x��'g6�%z]+��ص_D&�_ι�����W2��ނ���2�@��1 ��=/z쪉J���[��eㅷ�������y4���J���(>@v >U�),WE�Kzh��9���anϫ+"�7�},���l�̾��l��c^��n�)O��E��,�u����BZ�<wZ^$�����z��̬t��m)�Ʒw���t��R¦%��VZ�1!���J\.kx�8mB�=��x�צƤ�A�z�{���{N�{�*2��s������p����)JQ#��}%|�RW���8�w�\�2�����[r\��F�jq{�[c+�(�ȅ1�wI`��\N�;+:������K�����$#��kJ��P��)^��]�DB�J�IYQY�����K5k�j�{���G.j����
øE�MI��s��i���:����?�nWd�w'Q��L�ܓ�q���f��񌺳,cv�q��a�Q�6�����٫u;|��k�w���ͤ�����:�l���.��n�y=s,��F"�[���Xm�Z��.��U��y��7;�竮�sQ(�5���f���Fb؛y�
�����V1m6b���.��8S/o��kQ����f�5ʂ�5ѽ"��tz��OnW�sՇ��Ѩ�'�����6���1�lŻ8��rm��ق�Qg�����r�s<�١gG�]7Օ�oq�K=05�U�嘸%k��$��^}d^�0rו^\�� }k�v�iOd��rf�˙�~�*�g7:��` Ir���Q��7ʽ>���u����.�o�+Ԛ"�Oo:D5jՔ����2�}��׌����Nu��ێ�h�|%C��o�3p�����v�˭�2 )�M�����#\,�����>���x�����0�	�M�f�B��"��캕nK�*yO����m��1���Xד�}G�����E��+�{�jq��r��gc�P�\cO�!�{f��P�@n��Rm�:�P�TV-r�Fa�)Q�M�놶�-�>���{�.O� �ͬ�={1��=a�s��8\qK�k�������z�dk�ڶ�S��B˄�����-ު͢�ח���]�+O5�gZ{����z�<�O�u�g��	Y���5.َT�
�w�с�{5K����o��Ұ���z.Z��b�PZ��&t>�JєY�*���V����7��C�2_U����T�����/^��7�+��(��6q�\��=���cKȚ�,��X�a���g����c��#`��D�������ft�!A�]��
I��-�;p���U����i�&�,��S�%`�]�A�G��^)T���:���T��Ѳg�yb9ؙsv��x�Fĥ�һ����f�7��*9��(-�E�Q������^VS|[�&(wf1@��w��IL܊�������{{�ZB+=Z��U��V�{ݚ /*j���~��R�Y-s��qꦛ$]��{�*ʤ��4 i*+�s�r�U�|{t�2�panf�cM��������3]���ڽ�¢/M^̾o�x���} a��F�̜��X�����uv�YXv}��j���?��|���j�q#̷�0MYJnC����0W!�휭x6o��A�T��]��#&�a瀗63��Fz�gsXj�����[/J����wP|��u{V{6�cpո�u�B2Eۗ�"����8��V��^1.ڛӖ}y���j�sԸ��j3�3���}q��%��r��]���v�oR8��0*}����NZ��F5��q�FP�s�;��/�tݏnzt�����C��V� �iNxM��T��E�KZ��e	�,;��m��=g����A�9��ae�i��Ti��ӂ:�݆��nn��ݙ�*I���MQzb���+����t��JK�"�u_�����f=NG}�_v�h�yB*[�zu};��Չ_fv
���u��~�k������`�0�,�hM�c�UН��{G$����^ޡx߄��D��گ��wpF�mm\�3�-ce��r⛕�F��Q�o�k�os���i��stl1���\"��%�cXha�VnR׊��u3��̓ƥ]]R��cs�X� i]�y�?D(�6���E�#�*E*�=�!��h�����<�wP|���[��H��S~w+/7�Vit����p{0C<�7�QD��o[%����ܮ�T�P'UHA�uES �ڴ��Kw�7���qws�F0U���J�8��.��)�Ys�g��V���Y�N�{E71|�;�o��`dB @RWP	��{���I�ep���h� )��I�n*W3ᕹ"ܠ�{�ӽ(`���+LoPJ�DWMR:�5'Y��׉Z��Q7��'���h���꫆��>�b�Lڎ����
�"�;�t�`����b|!]f��0iˢ������B�c�7�,������h濰mj�gq�L�K0Ⱥ;Y�*���W�Ju�+��ڹu��$玦rS����{@���,�ڰ��ޱ|�4s.���K�����ge���t���͈^+s��U�I�tEIo4��*�#Fa/M���f,�GQk�z�iv�t�ov<�G9p\�4��\���4se7�6�O+�y]s.��kZ�M��� ����}����׽�ćځ�\�-���|�^}�6��{-S U�K,^2[#�6�6�|1m!�s�*��Mv�\�mq����3�//��%mË;� |U�(|�V�4�a5�3bI#$+%0#]ݓF��#L�̅����Q&���E�����h,a*77Fj*�-F�,H�S��c%D	�w�1����)6�5��5$E�4E��&���'w*"dc,lm3d1JE���[&�$�4�,E�5rۤ��DE���wA�P�QAZ4�Ƥ���B�"ę1��IɱF�!i4lk�D$jLQA<v&���$��9�  @� �}�w@��Z9 �P�+��*�y���w�8c���+t���R��a��-��S�|�.�&��4۱[cdy��i�9�0�˫'o�{���4�����k��u�����j=E{=����N,:��结:<J/>Թ9�Z��<pv�ʭvoX�&{�����sY�����Ȫ���}�/O�)z��>P���\��ݨ�kgC�̥�-]��E�-��SohJ���2�>S-�_w���m�׽�&N%^d�s
0�%��)��u�es򨛜���:�(�\,F�Ɣ��kqs�{�7Y�p�����9(;�`ꍧSQ����Qn杖�����l�s���M�;O��f�齲����P����*e�\���!�q���렪��Jƶ+�p�Zi��Oo�[�G��Kt��(����N%��C��YSү�ʯ�*5��pը�k�M<�����x��Ӕ��'z`��+w|����O���`��t]D���)<�x�T�I�]5~����Y��<���2�F�1^h=r��X�F|V���v�i̎ �����Q��42�����V�p^�}��D�J��9��r�.��%N�m���O��u��T�,2�T����ל�h�\�&�U4�mJ�֐Ά�7��=���qn��۷����C'5)n0�����u��>�:����O5�oTb|h��T(�O���}�Kp<]4����}�[U��/��|��`�-W<�w�s�35:�&��k��H�\���wcSy�@.�)P��]`�TP�5��cu�oXU˳\�>7�%̦�4��+��(O+yb{
�P�]g�<:������;^-L��g~䘚��k��"c]��H�o�Nƻ���*��'bGD�aܕٗ���歨�V�9:5)�����B��S��y������=s,��S~���ҵ�}���j��%/xK�y������[��K��{�O�:��]󡘫��V��No_s�W�M^�-oB��%`mj�T3ՙ�4o���,���v�F���Pq�yTf	�x$n1�;>�L�ck���}׳n�saQ%E\�2G�9��sb�L�����������}5܆*G�u��ށ������c@�ך��zz|�tOz����^�_o�e=[�`��(���5|��/�T]�_Yp�����̢��kB�F"z�<���e�&1s��,�Aw���qm G�&�E}s�U��z�q�m�˛�=��]��:,���9}�t.�^�]�Z~ոv��}��+�.����_Z��������=��;��C7S�I8F@���� 6KRv�ɏ0EY&�^�?/W�5��=X�y.QLps�L������}=w3��"�R]
躖���=5=95]����H���᭸�j��R�H���LW�R@�&l^f���^m�g+&�J\h���>����[c+�r��}ݐXf��\��C6�\P�U����h�T-������z�;���NY��
�t��XD�:I�����42Қ�|�>E���j9sP����w�\T�ފ#Q��똽���FEYP��?�j.�l�&� ����a��}���a�9I���۝}]�+�rE�1�9׶��l��I���^�AڽS�K��Zے����ۡ���ծ�^�kZ���ݺ7OOs�J���<�����2��)���A�U��o�Y�*d�.�R�ἦ����8nvr�_��]�->~�X�۝y�&-�;��\��*��P�n+|�i�BUaq�GMBn5¹��dO1�k`�&R�~��
_��LSؐ�L��O�r�ێN�k�.��k*�a�C��k�1�M�YPdK9p�Kne��y��'�%�N9�}Gj2�c����3*�C�5ݽ����o�=�1/[,�׎������lc�}q������\�
Ľ=�/Gih����v�T%C��˙S̈́齾Ws��vj�o��j�]�z���9Uຊ��uTFתkiBWg���FF�0k��v
}jw����\C�]n��ϻl�E 6`�@�:�k��>����o���X�+snڬ����5k�i�ä����
?rs��>�N���<��F_H�A�����8wETJtu'���<p����o�IP���LE��5�x���q��!�w�]�-�r�/����6��P�+~�.��>>Z��4��1�V\L�~tq�s�ݛ+�OZt+�H3��>�u�wt���֥�tz��y����(51}�}�_1���(Y���`�h�}��M�e_i;"f���<�7=ד��N��/k�H8��7"�^J�P����$�\�s{i*�Az���M���_#����m+��V�{�����7mNt9�Z��B\d�:C����G��n��U\s��zL�{�6���d2@qv�ghWͼ���3�,�|
Q�-�I�9�!(�%��+U��h���]�v�7��6�;��c��D�܆�N��χ5�x�
/<;'�r�k�d�y��p�����mƻ�
f5����/��\�a���<��qBl7�o���o�~z�T��N��k�5�O*�]���5J�ȫ}�V�v�)Ѯ����{2��h��N����R�k�|�Q�NJ�7}u���IgV�m�����)L�SohJ���z��o�r^�#��
����kw{�������~i��L�J�M�v�[W��끊;U4I� �%���i��хs�Wj�gt��Y~޿-���<�G�A���m���C�]Rss��t���D%+ǜ�H�.^�is�鯬Fyd�T��)kӰ���N�HIך�N-�v��p@��Y;p/o���u��b�4�2�ӶM����kB��:gG�/H�>����;r���;�*��[����me)긡P��.o���fl;��9�H��57��,�3iF<�=ԝl��*�5��]F'J��+�p�&޹�l���7w�&y\��zYkM(�� �P�rꍩr��(�'>���k��,�M=pv:h>�pg:hd���KQF��b��&���������Rޚ)<��wT�r�㑑�B���\+޴�#e��ҔH]��*�-��̀��#�~.�����} Vao�b��ǹ�J����.
I�}w#�Ĝ�,vAN^ˏk��{̴�Jýo#��&�*3(��Rφ�B=�Ř���������q����zIs5	�0�T%(O܆�])�ÐL*�$������{�()3N�<?I�kS.����I����k��+29����sy5���n���k
~�Q\�}�yI��f��Uj���MB�
Z�P��I���q��m<)�0�+���Yo���� >��n�S޷{tL=�����l�Uatm�I0���r.{�.��R�����!�oO�e):���p��k���5�'LK9b�:���2�4�qf;7+Txm��e�Z��?�����yZ��%��eb�����I��~��-~�i��<���l�~���ڽ�qS�c�����oG Ue�n����2���W�Л�.��nW�u��Z��������$�o\�y���̽�r���g�9�J9��.�{ �Yk=��SN\+�a>�O�=�clv.h�l(u��w�C�>!l����_��#x4�01���Nx�c��][p%BV1�W��N��������cf���֊U�q��r��unqX5Tp5��R�iBW��J�cb��5��i����v�8]��Z�vz���/Vd<���y��N���'��w�����-Y�fWan������jOl��|(w ;
��ڔ�|��������2�w\�ʒ�O.����m�)D����QPc��4�D�(��}��'����z��Il����:��Q�B�ﻢ�u�cw[(+w�,u��ҡqN�j�G���'38e�8L]~�&��b��{�
����]�<@�Sow��I�=r�h6h
�+�y���f�ﯞ�Shu*v)"{�鋆�t˕�}m��aπ]����3Z�]Il�j8�,��(+�7��޴�����1^��Z����&���j����Y��[w�`�C���<�"�q�yP%.��\�!��|v�sW��;A^�%�n���!��sOzV�0㥝w �m��r.�l�����7�'f��-��S��]â�t�p��·Q���l�+j�+s2y��jڎW1S�T.��S�^6m�o���4ۍvV�#�ށkc+��]�X�T�Vٞw���^=��^�ܫW��Z�i���ʭXn�P��Z�&'	O�B>3�h(}S|������=��g8������f�P�3�)>
��*��wpbqz3M�P��_�ڢk4O6:���n��'H�ӕ�����[�]i#�.����.�nr�J��LA�<l��蝣�Zs�Q���>3�si�m=�w�{g%��\����S[J��nv_>y�&�S�v$0��˻{���v��eުR���L\�l� �-�C�hX��9d�\k�Gix�+3�Q�m�<x��^]0�����^}F]�ޭ5X�(��n���9�(2`Ȇ�M�=/v��ۣ�v)E�ܕ�YR��>�E��7�����1�~��5���랉܎�9QH��A�[R�:]�����خ����u��8�R�p5����Yq�>��'�w�P���P%��[�Mu�C#�l����+��/�[�Z���\5��վ[J�ʴ����.��s�apj�V��Db�w-�-�\sƻ\^u�2�Ѻ��z���]n܎���?��	-y��Gz��-�aޭ���['3�ܥï_]7���FQ
c�J~Ǟ�m.{��[֓Y1���Gَx�NǦ*��޿���öf!zY����]���f-��$t��8�Z�\�S|�&�;��c�������*�Z�Q����J����l5oMT���Gs�N�&��г��m���'����Rņ�P�p6!�?wa��n>l����s-U������i<����a�ȴe輦���XD�ãNA�=�z��-\/!U���l� �����Seo*VIЄO^#���=�(�2�kQ��E²
��t9X�Z�9���Tq�k�o����(��s=5T|��pz��=�|����h]��Bw;�.��}ù�dOt��2o�iv�y-�o;e>�y�H�k\kF�N����+���v����6J���dRҹ�iv�a���V����|�#:`���z3tOu��S]h����?T���g��u��8�_�o�qm�c�`f��yc2e����8P�f��B�b�仺�����s �V1e���1L��M\��e=�n�_�\*د�sz�=s���}7�r����Tb�⳹V�X��6Rx�Օ;;.
�N�Ɩ�D[������I��kh@�\aq�2���)��Js��2���;w=����*�R�Z�ۈ�e�8[8���N���u-)�pu��T'q���T�wo�躖��I��5R&�:b�q�����٪/E�JR�ALwϦ
�-����ޒ#�<Xs"����\�nK-7o�"�ؽ�(�!LG|��	KC���N.n�<K�W�&�uA�WV@n���|���[��Z	���1��5����7���S�Ե��N�A�^�}}�� f7�y�T�I�!� ��x 6�6��E�f�;û��<�M.l��J��W�J���͋x^1q��Մ��K'Ej:v"z�4�J�O��������f���Z�je1j�����՝��{D�>�o_v�Ypcno}�m좓�z �n��:�c�e��X1;^rk���WC9��K�y�UpF��jYV�׶�2;��}m��IU��a��wWR�n��u!J�xaw��X�ei�LA+��[��c�&��BL)iZ�^hp@;�������+�� ����8�R�J��:�(Am(&�dz�U�n�eޛ��)��ޙ�ob���~����Y��DT�*U��=�y�/�*���J�d,���d)0{+,�Jv3�^����X�ͥ���l>�����V4o-�&��n���|d�+��;���0��*�¡g�<ݐ�l+k�bY�f�����ƒ�À���&�6���32-�0�Ύ7��-t9;�@y�6>Z1=�\��ޔ���Ù��������rǳt+�����#4���[u�����ZV��ﳒ,��ee����K������P����o7����)�|�W,���tc� S�ڼ�y奿�m�1xy;�d_f�n)h�[���G���Jf��i��\d��j�T��ǜ��J�������C�[3-�Y]z�WDК�ĳ��w�O��N-�M��E��y�$�|��K 	=�{�/���oZ�k�S!���V�x	�Z�f��X,��I�tޙu
�h��)�u��r��Q<��c�<Y�Wo?�m��������sU���*�a:�m>������R�	�m���$��F�#�xmEi�͘l�T(k�Dr?tc8��a��P,IP��y>����oA�5��J��g1����j�����O�.oq֌���aڗWf�����8�tOPV{�z��;�]6��IQ�1l���em��j5bQH���pu5|�qɑH�����jݧ�1�=}ü�����B��f�v\���4]!\6�p\05'�＠�(�����3�G�h�cdf����-�<b����-9qz���Sٝu@B�ޫ�*�bU�A9���o�,Q�V�>��
z�AcI!gl��B�*�_���b�M�P�����Rֺ��6��ԇ��I$b�NN��Y�`�K2��7~�G��dʴ���*��ˮ��.�����iL�#Rz��L�;�B�o�hˏ���x�oʝ�s0���8Sb�|��3i$���@u�}ss^-i>�pV٦��Pm]΋*��<��ј��R�s�3�&�����M�1D�y��������^J�-k�*����q*(��<U���4QE��㜷7���˜��s�nnnr�H�B(�#s����v�`,�\��������Dh�2�b�I��E@FƣwQc�͎\��i�b�#b(أA��ncIQd(�Q��lܹ�PE0V�Q�&�)�ō±Q%�h�&����Y��Ѳj5�1a"4Rl�Ţd@A��R��2[����"�Yݵ���fD�nh���9��R�SC��jE��5k�ҷ<��I�޸(��^7��M�	)�h�(5��\y���k$�f71E`ܠ{qA"~���z���;�ɕr_���Ȩt�t����+c��r���]��PQ�{�Y\�s���>9P�3P�����p�(_]�86��'�&�F�k*\�V����=�;S.��䘚��k�e��&k����\S@W��yM�ʫ<���>+{��+UZ�I��7�Nu��2��Pw]_GKƠ�;�tF1�������ʈ�Z�7���N�b�iŠ��ʝ	<�s���>�7���8���������b؉���t�"ⷩ�`�K�sZnr�K���7�<���r�ת�W�&#�7_s�ݑ�O��u;1�!��8��ʁ-��'��S<��u��]�׳���gYsG�+�C��	��U�睏b�j�c�����\طI�����_f>r�^>�$O]����UmKOWt���_�N�u�1ŗa�j��р~�y��0�D(Aga������xx*6EaWϠ�@Lzo�2i�����*��ި�2��,��Y��1�����uw���SMu�9�n{�p{/���w�ʐ
��H�i"��hm��ᳬ^WS�Ȏkv�L\M{�l�G6m���t��羌�yw��|;�s�ܘ�Y&�ǫ���)�Ͱ�moPg3��(o.1����5�P(t������*�jRW�_����)�Vg%�Na�ݥ��_�᭸�j����P(t�wϦ
�Z�'!�7فOb|u-���������}��g[b��3�l���E�x-OfEk�>����]��Қ�3�n�)�a޵��
���9v�w��h�7�Y����>�E�y��9��u.{��X��r���n3�z�+z�FUiK�ۘgF8qǍ�GhunJ�5t�f����!���<�[fq�Ų�iT�Ud�g�q��+�N����V�rV�d��ŔAL�ɠj��);YiD��������,��dO�᪄�t.o-)�{`����j�>��{u-S]ټ��7*�':��T5�_j�z�FP����bɪ��������f��XWڻ�]�"B�o)�"m� ^� 8��>�pL�%��J�.mЮ����͟"�-��/M&���w/�}�P���ۣ�_C�&��R��2���1�&��]����UweX�l#v����\d��S�3�6�s]D���Z6�S�ܮw�R��8ֲQ��� ]�W7�Y�ֽ�%6'������Ss�y��Q�V>v�y���_]�g+�l>^�L*o$�}˰�������79BT>���s<bT�ofḹ��N�}8�}������'\^|Yw������1������}}[w`��ƕ��al�8��|����>s�8��v�ʊ@l�� �wN@���4���7�a;�q�
��J��_��ƞ��I��C���l�:me-���Kײo>���-<�]R��R{z��	O��3C{�`�[(��}����i�e���~=w3Q�%x�]�|k��e���q����2	%��tna�{UB\d��

c��-9�H�Tb}����UƄ�P�OUuewr#ut����*-�����S�%*=��\��,d=�,�Cޚ�j��´Wg�@�n`�}�ڒۖз����u��FV�&��t3�R�)�wS��u�s/T���y�\ǽ-�M	����sdYn>z��,P<.4����Wؘ k�W.a�]���/q�X��5 wé�p��,�͢��Ud�q�7�p�J�faz�J��k�2�	�{����\�'W%�/{Qi��7���R��Cd�6WdV�@�\�eR�ŗ�5u����<w�j�,�&�q���DZ�kUK���=�k�R����X�;ꈞ̨�z��7V֪�q��-p�<pti���i�f��ow��Ld�;=s>��3DK̨�Z6�5:��w	KЩhn�٧!�߷eG`^��̜A�֖��|�Oe�.��kc��VRqy�^��=3<�/z{���~i�vu��\�*�nszLQ*�Q��z��V�V+8M�\�Ϗz^���}�';�0�����TuW�(���z�C�c��p�jkk���k���\��;O��n�;����̈��\��YWs�,���Osٲ����hlS���6��x�	��*lP�m��a�C1*��θ�ַg�b|	��-�Wi�ޖ/Ylb�,Cf�ȹM��V����:s�Q�1�����=,�xӥ�r	�_[�֔�y��Y��&��[�^�����.�'���m�kq.�\8.���O%W\�N*�{(�@l��!��w�eTJTkS{q���jٸCz){�F�8�&J�6{������;���������?a���E�D��=����O^{*c|��?O/tOԞ�K[]��P]��*�-y��G�̕i�ٳQw=�a�2֮���u�v�q=�m�e�|�15#%�aQ�ѱ{Z��[����ި[�k�J�;����&����LP ���v�z���݉�-�W,�5Իw ruxeD%��o��L>
�d��������w�\��ԁAŰ�Q����7ܷS/��䘛U}	�^\��%�r�{�q�Y����cb��@w0:$���R|���{'<׶9��eg���w�<����Ѳ�pv����]�1�vU�{V�����?G��&�xu9䧫z��꺎M��p�=���ghT��Ⱦ�}�h���pz���<J�'Z�W$���:�>�jS*�]دM�5������rg�{�����7�)P��fd�JF!d�SVDa�j��^��G\�<�.��{�Uz�ѕ;4ﴱ������c��c��{�s*�XV��ՈznH���*r7<��Q�'b��i}V�Ͷ��J}�g�إ�����ǳ<���vY���~�I�â�����b�/"Ҥ������{U��������63�u����k�6��MB��e���!6q�ḥDv�m:�*�p���Q˛���o+�.}�T\���O�];f7���*��OWt���cb2��߲�Eг�&�7��泺�|���dk�AλW=V�{�Ǘ;U�)
bh�[�d��΋�v�u����Ol��@����PC�/y��SG`�f�{E��{��31T�q>��Ryq��p���R��P��}�w��R��)�OcUa���bb�N�U�J|j|�>�N>�����Q�����8�x���W|��z4>���uAM(u�;���T ��"�wy^��hK�ft�<ԍ��f�is܄Tŭ9Q��}OQ���eLX��R=�]�
�&qԨ�̺4�h�kj?J�p҂��ﴽ��ur %�¥d���*��h����@�I.ytszx�h��9Jt*1��٘k�ic��03'F���j�����WH�z`��1�����3�r���&�q;�<=8?�ҕW.+Ot�ձ|��:,u'z.�Uz���<�J.�s��kT���q�¸�R��1V'��|�y�c��x�p�X��+�q����ڨ��{��mƻ�,��]�=c�>�}��Uz��B֥��q����ē�5eDb�W�u�p���j���ZT����؜��q.߾�ՖK�|�:�����r�|����'�v*���1X�V�>Kz���V��P{�d�yBy�j>�����f{����箯.s���p����Sĵ!�C��~���mašv16�<�mi�+��%NϘ�W�㐨>�ｼ������!g_�_nU�6ߚc�6�>S�*�<ѻ��^��P�
��K]'�v�:ٌ�ʤ�jo/*e@�ѩ��N�W[����+`��T���[���4��'��z��9u.ݙ��;�x~S�0,�[�Ip���6/:T��t)�s�L̗ij�iE2C�ׅ͊"��eQ�9R��ⳛ
:=f����nt[�Z��c��9��|ѝ�!\�V�7�����4,�_�s��oR���*�˦U�z7V��-�[9�oto)`o�2��{^5��J�F�{q�����O����o�tX��O��Ƥ��#(nK�;���Ғ�,7�w+q�'3�v�=<����ؖ�l�Qs����ߟ	�����Y���Db}����J���6���o��Z��[��l[#������(�H��W��Ih��y�>��wd��~�y��p�kp����}<=�e0o�����x\���"�g��j�Wt�&_K3X8�x5�/�+��ᜥ��{���m_��?O�>9����
sNfE"�O�b�i���׽Z�Hqq���r{���^�IKң��=p��������>������z��Ϳ>ɾ^P��ya�t2W�Lw\@��*'��_�j��gu1���C	��zB�����K)�]�gt�>�|׵��Œ��>؁;��W�t�:=��lx\g^_�;~��Y�;�;'/;��U�í�E{�V'M�&�B�T�O��.<�߆�u���	��l��#`?�0�Z�x3q�\bw��]JWnJkd{nB����ڋGM��{E�p �3�!�[��Ro�p'�Ո�B3�x�G�ǽft�����*��w�'V������i6��Ҏ�J�ғ���WP�H�Y�QY�V��z�$`���%�(�P��4�*��iv�(��z5��U{����P��z�3�+EGzrN"�Û2��L:>��.ù�uz�{���ˁ����3̲q��=�&��U�k���>8�>�e��"�3=�oo���=l��E��m�ó���_���x�dz���C����X�qT�ꉙ�>w�r�'%ՙ��� &���u^���3��V�O��҆z��+Ӟ��*�Tֹ�zZ��+�_]�?�4�:��#�iK&#c筬��t�X������)<"�EET�C_S�]���}@>��c�s鹅B�񯸲OW�a@��QQR�Y�q>;�}�1J�tll7]>��IJ�G�>g�7��q�TF�Ω�p�?q {������x�Ng�GT�?)�SѮ���{�U���+���z�9Ӟ+������z����2��PB9�x�W��My�p���7���p�� w�����m���2�>��m��q����׉���"�{>�S��tD�\du)��X������xB���ψ����j�zW�YU<����pTNdp�^Vtg]b��Mfm��0]kK�4����H
��Eևy�A�����IR�٘����͡��W���L�Y�/q�{J<�)�a��uyn����QRo�;�y�E�Y�;n���3q�}y�sv���u�Ы��'��7	�1Q/��r�a���A�s���y]��E�1���l�:�G�c��%�@g{���~��iK'��a����պr#nW�Vo\h�� �Y���Y3�ߵ�Ω���q��꿟��q��ʱq�ʐiO�U �|l�©�f�w�<+���]Z�2�}�{��q�؄�^E��R�쨞����7[,5��C����q;Ӿ�����mH���u1]S�'N.�x�vڸ�C��q��9�V��9�
�4���+,��h��s����N)�h��i^��AN�\T�},�[,�W
R�x��x������QO�㖗%��'���T�l�wl�\��(__���Ɲ�>���Mz�[C�{0�[9U�����>7��͘W�����JO��:�!����������P�۱������Z������Z9�z��ȏ]�����p�]�"C$�!x��}s^�T�ٜ����
��;���]#=���x��r7�<^����m�ׇdD�pV��K��X{}=�kz���B�T���C{d⽇��X�:Qf�������l�ʘ�K�l��园�����H�nudbT7� 'mk�k�'E[�<�Ҩ�o�R�L��K[k�.�^	x�L�ˮF[3UI��������V�-²j��;�������GhI|��d i>�U�����W�ٲ:�~����L/�,�(N��PVY#Gc1���v5;�i�cp�pH��鞿��1e�R��"��87W�-�j�m��������˝s���V+޻\�rd�.n��n�]!p��Z
�g(�:\�8�>���#; 璝͒��6�2��]�[�vu>��,��og^�a;Mk��}!yA�u�!29�۰-�ښ�)��[okq�;���2�B�wt7����U�M�ة�jY#o�-Ӻh},F*/��KEh�f,5�U�t�'6�=�9��0q0w��Qj�э���ZaE�:wpN�3�b=���y�][����]�m�Z�f m�(N�炗7e����6�9F|�٨E�u ܌��3��9xU�)�u]G8�ʙ�5.��.�\�}�Ŕ�`��9�4�x��[�)R�>L��tn��r��]E�����Ve^���7"T�MU}��y��RoI\��I:Ո��E�y�B���}'�V:ᓏ���U� ��_3�sv���K��:�Y5��6f
�wf���H���E�s��o<_�����!�,��>wc��}]dM�v����o�%;�X/[�|�,ُ���O����9�=jo"��$uz{�V�:���`s����}��N�3�����e��1HҲ�Mr�f�]Pe���cflմ�G)ͮ�+Ѡv���a̙�M����Zx
����5[�� �J	F:�vo����ǀ������X�pK(�E$3-��h�i08�v!��g�4͸�{�S+���gnr���$��y�� ٗ/)<�����ˮ�.�5*��w���7b�4���/p]���5X<���iΖ��m�$+�|��|����&iVuܵ.�<��l��Y��)��˥�l'y����ctɣR�҆c!�܇WV>m�W�ӹ�ݍ����+�Z~�`%����*%�[�]tW���g��6���o?Rw ��6�vø���҅H"rP��2��$���UY�v��b�-��˻t�y]ڐ9��	Oؗk�u�\�٬�3e��Fq}7���9eZ՚��cW����ӌc]jwIY�^3���˛�՝��ׁ�^��.�vQ�"�X<tF�pq�����������T�JˣM��i=��/ژ��qWc���)�}ؔ-��ܥ�������2�<ؠ�³hie���7k麂6�c�1�qwv�h�e�X���;!NT3@$'ZV���!��m����ʀS�8�Y<oN���w��Te��UYv��@��YDp���\�x%���j{�R0_�ki�ث�)��Tɽv��74 > 
� *�� 
�[���]�
+���c^7,n\��%!�ۇwX �&���"�I$nsb�͍��2bwW �wnnN\�LX�Rl�7J���i�\�/;�P���Q�*���6���r�X��ر�76-�]���5nNlm;���;�rݺv�������s�ݫ�b�ܮ�����m�k��H4d�sr�nn�����1�����s�s\3�WJƋ���r�^5r5�\1&�k�sr��^.W��˚抑wnj娣nk!����
�����]���8��\V���;j�rm�+���M����ʵ��-s�j}Vj��u��W9���Ql�V�B=�	,�''�Ng�9�����O.���ި<�{/H�|w�3�3��o�6˰l]U�uG��.�*=IF��<O�3`H��j#L����ϝ����zЋ��Z�?Hү=냵vά~����;P��������=���"d��E�L��Ftr�R�;`z��%G^s9�X����nߺ����#���T�%�Y�F�<LL�WQ�떏����\���QY��T�2b��du-��οs�}�>��>���~��Ӹ�S.g���nL��9
�������6��;7\����<>��*)���Ss�|ǫ��|`�3(� ��Ӂ��O���d���9"Tj���c��|��ϗO��?mǳ��w&�σ�~���@{v/�>ɓJ`q1�N���4�a^׷�0��X����zt\m�����zo�w�?Uq���^�q�;_y�Y�=�'�{q�3��\�]���(�K�1�2p9>����q=��L{��<9��ddB~�ޗUdy{�3u����Y<�����WX�� �g�ߨ6)a�i��*�;�.� ��+�N�7�k����"��J|oF¶�������!�&�/&8�yuq�-��馩��&��_K�a�o7���a��Nj������Վ�G�a�m��n���#C�2�BRSt%�'�њxq*C�s[W�Vp=��ܽ�aH�����FR�͋��g�uu�S]�����?D�aIe�4W�дઔ�]Dd-�U��O����	j�ЏN��Q��&�A�`F>^��^����P����+�}���x����YX��+A�����q��Lԝ��;��r�y���C2y���~+Ԫ3�=u�q�:6-�'�>U}r}��}T�������+�ʢ"�����������������[��a��n<���c������O��Y$Pg����κWᐮ�Y������xhQޏS������#UNQ[�:g�Z����z:�fю���f���2����Ft�nu�ǔ���AoՂ�=<d�S;���K��Rqo]����i��@�Ϯ�@i�2o�<���	X�w�"9�����N�����s�:c�^W���Ѥ��z���TISq %4}$LJ�pu���!~ɽ��1�X�`y�|u11���p����}<=�e0o���7�,�tt���=����6D�g�i��\wx�D���mJgG}��7�*6�~�o��O����C���́�<�d�e� ��5��R{�����E��!��+zp�t��ԟ�6�N�q�Txs��3�o��C�eX�O�T|�ɹ��i�.;�-�n#��m�f�3DM5q�	}��#��[���6����cu�'c������6�돻�_����3AM����ܿS�X�>7�����w&.>Mz�����g�P�|��G��vns�gѣ$�:4��@ɇ�'�b����yj��Y�Lu�;�d'�]��#�J&�k_�A���xuO��Kz�{4A>���uZ΄U�f��e��~܍�c�k�Y�=��Ω����qϽޡ�=�bt�̌��{,���]�=���������q�v�Va����N{t�:���3>�2���y�B��m�V��7�nr�8r|����r�z?:j���׊Ç{�^���"O�<zʁX��YD���ɺ��
��F'[��L��*�+�~4����g�J�L��&t{�]��t<�6g�+���i���ϣ�/ǳ�}q�5�u��*���漀R|hǡ�T� >�3���,_]W��9��U��i�xq�=LoJ����.+�-����w%��q?FBˑ�ŗ.�_��1��'�Һ�zr�TSyb<c5��$e{�+/:5U�wP��^��^����o�s�1�*!���C�F@�S9���7z����������V�kn��ԣ�n����_Zě���WOkFQ��ų�Xlm��	-�n�����c��]�,��.^���D����<����xȕ8wn<���4��uJηQH��&Cx��:�p����L�PmM���؟=�ٹ�/rv�'V�2�lN.9�~�#���k/�������=���ʈ�uL;�_i ~��cC��	_,^�kjj�������}����G"�ʢ��֑Ϗ�<W�����{�F�ޚfj�,�C��KM�M�B�}ّ��rH-O�e����3��C�Q�������v�t�~��׻�|�N��\���}M;|�;��>!�u��"d�����]��K�*#���?yY�.*�ff<;�s�6�ݻ���Z'V:��{caBӃ#���L�B��������R�9��xZ�}벵�J��]O4�fr��=�>�M�O��`wC�ܱ���L.����vU���FUTd�#�}��Y�'�=�ͼ�	�����P����n<�_�����_@8���MP��c�u���նw>e#Ƚ.;o.7�rz��9�vTO_��pN?�+��9�}�X�	����-��n�}ý�wYLm�+����ޗ��J���׸�'�^/{�pz��f���p~*=9=��Gv�]���(�G'=3�� l�rrN�4���.�^�dxc�^������~�ۋF�r葓"�&@>������7#���])�i=cr�n���PG�S�#�ĵ\�T�/_TȬ��q�Ѥ/LĮ�Y<��2����x^9F��Vz�7O"�]�5���+��YεR��Ib�yK�,`Li�����3$���B|��ƥ�3����
�k+�*����YS���;�ø>E��j��t�@��}k�E4a6�3��V��}Mb^`������O�ӶY>Wa��Du������r���-ueY�Go�l����^���Fx�zw�(>u\�M�
��R6�.Y'�� ʨv�Wz��dov͋J�=t}��Ư]��ޯi��H�{���9�^�u�\d�R�'�5�V`T��޽&k�B��B��z .�W�U�>��|n��7���w�x�9��C=�UT|f�s8G3�񹌉S�Z��z�z���p@�FPJ���:���z�HU��ֆ�����{�Q|ҩ�X��)��ۇ�D}��d��8� %��D�o��%y�&g�}�C��y��o���1or��W��}7}��^���_}(�~��<.����π�ϿWQ�-jf���ܞ���lV��[s�=���Ϗ�H�G��K�� �������g�*��ٿ�I/��^0p�WG�}�J.�g��]��k�w������z���R���=lꜙ�,� ���i�^�ۻ�� S��߯eAu�祈��(M1�C�	�����$�%��dP�/�nU��H�-�A�վ5fV��G4˒���e�h���)@�1o0�Qp굨����>mK,͚P6������E����g�}-�ޭ�\4:�g{Ã�i�2�Ņg�v��;� ��*�w���BS�<��~UR}��^&��{ޠ;��{v/�>ɓ/�ؽ�xF��;|�J��v|n|:��
��Ztm{�������.|߮ь}�Q�����g��b��sY��Uӂ���;�p�>%W�&<�ᵡ��>Ӣ�V��ަ=�Uc���\w��e�:U:��Rh����ҽ��X����B�ʜ7Y;����'tÜ�q�N��]l }q���!�u��z���ff�*�^�;�R�y�c��[�G��j�~�u}��R�����T���y�~w8�	^
���Bw+ޓ�z�5���,������'�Iv[��G�1��VE�;���G*ڪ>���tσ������{�e��Y�qݞ�B�Μ���Rs&��skM���W��Ck�3�_]W�c�ȗ=��U���x�P�zs��~+#��=מ�R��W�U{�
O�C=�x�E� �(ȱ}t��qfT�qMՉ�~�ޏS�\_��5}�U�� �����5��3lñrQ��|I@�.K�#�mʍwP}z�^���G)�I,ǾՔ ��3�ź�Q�u����
�W�`�TQ���Լ�qJ�%���}л�YSaN�bm���R�Y����nr��;J������y>�MW��p4e�$�����;�����C����d�v��%�ԧ����^��+c�CO^z�:OGB��K�F���!�3��007���5�Ě�{�n����MF��&��b��_?W&��z�ۏU15�.j 75�E���,�^�UA�=��Ýԏr�h>���en��G#o����?[g �s��G�p�{נ\zs�i̒Ѫ�퉍[s�#|۝Ղ���$L�*��G�l/�܄�wͫ��~�"|r�<O�̀m��ژ�Q�t&��{��9��������30��U����4.2�.5�S�|�R=?+�0��:��W��;_us�y9}�i��>P+aL_�}fI�|OPɇ��a����u�5��Lw:�Kg��t�(����^VzG�΂��z|����ʐk��L>�;�׫t�/����QV%�e�|��Twm�Q��=���=�i{��{�x'��ɡ]�q��ڀp/;�E������MK�9�k��ȓ�NwJ��^
U{�3��P��z�wۗ���9'.:X:v�#�%{���~?�x�����Bb��1��8;����[�q��Mù��d?;���U�f>�(�#Du�b����#P<��n����o�vg>6z�#M�ʉX����r�99{oo����Gzt�ޗ��ޣ�Q]���
�::�.���^����1�<��l���������L��z����}:�	��4g��}�(+]Ѿ���s���*wb����N���Y�]z�.G��ٟ ����	���9���'�9���֬�0�bJ!�H����j�Z��co�-tc ,g�u^�}n�/8��<���"�	�`dp�~�*}ݱ�/�B���L��R�o�l.ʔn����T���*��Zʂ�Lu�>x��1+�[T�B���ћ�3���=��l{�M�����À<���`��=u��l�-�c�8��%Oj'�-ߴ�н#�{} =7�1������ )�?E�^��y9�a���
I�א�Y���U��F��>��V9�LyD�֑�>��\u�F��z����3��.�3*x��^��=`��i�D�"gޮ㌿7~fy�|���m�ȃ���#� �����Nu���~U�u�����Dp�� w_j������S��,:�{�F���.�����B�Sw��M���fϾ>�d�����t�&�K'�L����0_O��\��Y	S˯mY3�\�_����ś����U#�y��>����;�����K'����n��e����?6�6��D^�ӳuFE��2r޹Z;��R�[������Ub�:�Ws���p�7ʹ��qD>'wʙ�Q�z�}B틧��z�"E�'�C�߯����U�C_4���O�Q��v�����2b���G�.V�X�tF�"��@�ݽ==iZ*��=^����m�{�j���U���>��w�d�O�TAf�j,���3���w��'��Y�m-7s�|�����y���ޠ=N}�1;�ۖ.�L�\�/ƫO]��Qx��_��?|+tù+V��㾀@���j��������}�<�����\����������������i�?��vv�|=t=���:,ү��B�`U�G�C�^�4D�;���39ί�ǽ�z�wt��eN�9�a�	�,Z��㆝�k�n�f�[f���U�v3'<���j2=�z�>�~:�xn����Y�S�����0�ў�w��#�4�ث׆x��}7[�7�X����.�C��Y������������u¡vT���I�RW���0��$��籞�{et�3ЮiQ��'�������{N�������[�5<@6Jj�^���Ռm���uO��~�I^��$'P����|5����W�V&����/K��z�<�a�w~�Y�>g�˳�%FǏ�`�x��2�c"5�w�G�ԅ\�ֆ��^�[G�-��"�����pǗ>��y]UL�{5��ju#t)��=�s�V_hˁ׶�b>�9x�K}��d2�q�X�R\���v����6�L�Oz�e�;Plv�8'˺����}�gw
ȗe�k����4(26ڣ�L�ϵ)#��ys�a�,Z�WӄS�����G?\�U��%�P@J�����I�L�9�����CVy�א34	�2w݃��W���������3޸:n=^��fK5��|'���^��qr��r�^O��'����'=�ׄp���>�"}�=87ޭ�~�����e\!�8�q0���Z��Fr<�p�]C��z�T?r�S�Hg�����ꜙ���xV���	�>@
����~V��ȑ�4��ӽZ*�����)|o�~ۏd?;�/J�4W����D�cNzo��|(��U��I���&O�ǋ���hs��JӢ��_�oKӮ��8o�h�|��^���(�ϨD�AΝս�U��p���'�z%a�����S\[t��-�m��{"7��\v���55e��ԅ����QU���?P�/cʬO^�
��T�6p]���g�J����:-��\-b@�=�v��z�}��2#�^��~������s���Y�p���fa�>U��Y�\�Q�	��S>�R�=�6��^��{�s�]F��^t�ϖW
���;w,����ċ�#�_F���o.omd͓��n��.�|��9h(�KJc���ЊWQ��,���e���֕�b���Yu���p�`��=�M9f�ֻf�$7gP	$Uս�wc�k8<#9��x�����^�z�Sj��C�#�!*�G�Z&����pα{�۵ r�3[�]_}����k3(_�8i%U�N�&W�B���oJ ']�u����\}e�8��~��%1*mTy����o^ι92"�υ��]EW�ٸynW����?</S��o.�E�[��y�n�[���s6���k��s��� ;��Q��N��FogY�,��|�0�^�������[�Unm�xx�'�2��'1e��Ѐ���1,F.V�z*�ѫC�I�Iёd��A�v�}���Uz(�:M)K�*�8�s�B�[�j�0�%G���=35^R��W����c/3��|�nh���+�c��W�J@�Ƀ��W�}}�T+%K��ɿ@�x�_�`�P@�5V(��r�����]\��V�T&y�\<��F]��Hf����VG ٵj�H�gj|� �o�zիw�����~�3jލu};Iw+t3��v5{��X���v�����
��4��)��3z�5,�F�{�ņ0����z��X��n*���zM�����cJ�>+�N�
��#��IXi��ҧ5@���ժ����[�>468ˆ��|`����Se�b8)�U31c�%��\U,�Q�ͺ4��
�xC�B�"��/�r�ՙAJ��0��⨮V���ݼ�-��Ec�%rvOI�x+�:�TC��5��)]յz�:�G��WՈ��
��Uvl��`dS}�4q�Gx]�Zk}n$�=�{�lV�<��C̐ryJ�5�N���v�o֖�
9�v�6t��Z���j�8��˙y�b7���,%�5>��-�a�����9y7�΁W�b�K���<SYfWQ�Y�v.�I2���.�^?n߅G���|�|]C�ˈ��2=;�Gr$�<79�ZD�y�_)�@jz<�rYn������L�(��w�mw�s�ښ��x��ˈȹG&� �$�1�Am��9���T��I��ڐ�݄ݎ�D��U��P����]��L�O@�
�;�I�񙏁`۴��t�NP���Y���U���йv�������w�#-q��o!8f�@J�ӫC$���q���c���'�)/��G���7u�.*��Gr�=�緬M�3�6��ǲ�:ְ��uL��̲��/~\�4$0�����1Gz�0`=3�p���|����ឨ0gD��ܾB�h�f!5=�� N5�*R#0�������'E3}�Ɔ=y��׻�;�o"BgSgUlX�P���_5C/�%n�`��!t�P�G��_xNU���\�s%��[Hʯw���&H,7v�a��3r�ty��1�Y����Y��fu�1j6�6��r�`͐��G����&�ժ���WeEt�|_����Ԉ�Pr湹���+��.sEs��c�;���W���W4�<�5�ᨹ����,G,M��G).k��+��s�(��k���us�ssnm�r�.WM�FܮE�r�b�L#r���撷"��`�-�ss���ۛ'+css�@�̜��M�\���p5;�9�w�\�k������¹P���-�w-��7*�E��5E��wv�r��6���Eq+2b����\�]ݎjws�(���n�b
�79�2Yݣsr�w5��v,�WCr�4h675_/Gݳ�+��bJ�'"�>��鷷hj�����1V�^���tS�Y�x��b��#T["����"�YJF��SJ��٧�TnҪ��\���|��W�L�o��3ވ����]!fx���G�`W�&j��z
Z�}�P�֤��>�aW�g���}SND�z�V�x��P�zq�_���%eX�J������u�-zxͳQǰύےW�X��X�U��2���n�M�ׯÆE��r:�����.��7������3~0�G>GĕFX
^�Kn^���R;.+��"}7	Q��~�C�߯FG�י[�z���� t�:u��e�b��n���
ݍ�$Gvo�����9�������n>��q'�V��/+����p�o=�#n>�SNd��@ϣ��~Y�녾��+˳���|��E�6>i���i=�вS��r�8��{'���z����U�g��=����Q�%��A��!���J!]4xt"�_�
�mW����'�>>��>�m��6u*D���o��>�<��3"���Ff�6=�Ae�\k>J�~�^����3�e-�QX�k{�%_?&ͦ�F?�8BӃ!��d�������m9��ݖ67#����*;n�Z5}]Ǒ|,uv��Z�j�QP�<�#�Wi��P�ւ7�]��{�,�x:#d����9[:e�-05C8�Xx�8D�i�z����葫�wG֐�M��R��'Y򡠍�!=��b��]r��D��7�[Uр��ъ�E]�n�}���A�y;��Pu6�>z��E��eH5��U@ɇ���b��[�[�e=��{W��wT=���!��7~/�����N��q��x��u��7��ʑ�Y9� �^3��z�ʻ���(�DI����?ի}��t�Tg���Ϸ�*���T��ܽޜ��U�k�k�.5�r�)��J'l����ʭ y��|r\�uN�x������?;����~����ڬ���5%�ԧIe2�e������g� ��}GGt<�#f|���)���5�=�7WO����;ݻ��n:���VT=���>�C�T0�p�����A��}V���m@���ڍ������ G�8�1��W�T�P��9�+��R��d��3Ơʦ/��W�c��"o޼���Eo\U��]8s�w��X�ެ}�w7���~�=�>��
��F�d�Qa�����m+����GV��o�]6Sꨟ���}-ߴ���<�}@>7�yQn��`�)v�w���պU�ФƼ� 2g�lJx�2�^Dk��C�+����#�Nx�:�#O\g�do��Y�F(�u���';��hц�+P��ܶH�Wf����~	���'�<��d����֓�]J�'��BJ_-��4�AD�r��"������z�(p.�_V�Y��O�/kص��Xm��.��n	d�@���9��1�^�b�Д��������r��H,��Q���A�^�<|\�Ku��/Ō`��R%��1����i_�T����U߸�hj��>�'ܽpv�S2)̖��L7p:�����������|={����ȱ�"�׻��^J�:��p��|G�����
TĿ��z��3�z�d��Q�˖�kؼ:�C3�i*l�d�ȹՓ޵;ۗ��w"�7^'��>}� �~��j�z����TN�vk;}v2=A{�����=Y�q�6׶�=�5E|���ޯ�� =��ʐk�S�W{%j�~���z�I��40~�P�&+�~�k`����;=m]Co�\}����{��z�~ܱ��a�uEo���^����&W��Y�9>
�l����f������~7�j�����3��KŚ�+j�en��J�]��ئ���~�g��:����χ�:���`ү��|��{��Y@��%t����{�+��0}�����U����8�g��J��a�	�,Z���A�@y��Wz��_��B:�}\̏zׯ��޺~<�P�<�xVvT鸲��3A��o}�z�{\��&��߲�`SC"W��
t[��M#[W�|�d�
��y�N�k�r� !��;�k��� S���y��^S����
w��v�U6�N�m�s0a�xY�(_"��X�mݞ��\b:Ԥ�s=vn�bAp�gn�#z���GP��[Y���������Bg�D{�z{}�Ǘ������p�]�#n.Y'��Ϊ�� �\ǖX���i�;�s]G��,��w;��+������^�u�r ��{iFEk��R��ה�$���!)��uMσ���_W�V&㛿qϣ�#�����']�f݈C׃��t������m�lj����-�3]�x�޿RO�hhG��y}V*d�p��_/I��v��}�4��{�o�U3��f������-��į9���S�zx>�A����:ޠ�ynS������Ϗ���~��V{�Mǫ�_3%�D��i.���P�;یӼ��繛^���Dx�w�+#B~T��>�"}�=8/ޜ���d�el@29�nǄ.��4{���R�����uu������ǼoɊ��m_��?z�>χ���XC�re˞��>��2,;9�HNC�P�A�����N��˯3�s�����|���+��Q���tNrol=�Q��Y��'�=�=�&��*jKcӁ�Zpo�o�·��\�.D7�ce���T�����e��B��c"��U�yo"Q͒�&�~J̓%�9z��Cځ�:9�������,Pk���=�b�R7(�o:�(.�TDh��\�]�dƭ���}�tݗh�Z2	:��T���N.k�$�����c��~�&nWwtUn����}�b{β������Į�d�V6�;���t*s��}�Lz�f{\�6qj�vW�!���#���O���}�����fV�*�����5���7��Ȅ�ˏ;�����~j����u^���^/!z�w��ʑ����;$�bz%�s���Cл3Ц�p�O�+ m0bk�#����z�5��9��W
Μ��N�r�uY�'B��+|gj=}n��ˁ�s�|�7��n����e��Y�W�hZ�|q���Y�V]\�H$:���.ܒz���t&x>��T�����_�Î���z���V=l��{�}�xns]�l�Ҩ���P�a�n-��`\�X�U�г*Y�n�K�����i	�e��eӽ�A�1��/G��s��~u�o���(�>$�X
^�2ۛ����0������tR�iٜ�Dߡ��(\�z�g��^eoz���� tۧP��f�<��7{���9�W������]�'ޙ�����o�~Ws�,C��=��\8��z�ۏU15d�%?z`S����s�@��p�+�gu	[y�%�Pm-x�F��,yWx1����m��m��O��2NQ	��@a�H6�K��J��:��x:�v6RH
�v�6ٝ��p�˱Wr@�8���P��ʃ���a/#�����s��:��x�F��V��Me��5��Ofx �G=>t��3�^�C5��&5?RG�}9��;}�����z�����2����YܕD�v��K6g�2N2$�v ��2�HU���<;`)~>�&3�W�7��������<]��������v��3!zA0�6����q��*|n#��G�jA���Ok٧֎U{hǹ�G�>��PFWO��F�ju�>g��~ۛjW=a|`�8��p���gz:��<�ގ��E��Pu6�>{��P�\�+�Ĩ���Lu�l�Gn���ߔ�7w����-�ܭ��g^_�'U�/�#ƹ������ʑ�,��^�M� ��1��k|�;���.,���}�����]3߁���U^�L��B������^�RZH��%=��ռ;W.��IZp9�a:�TE��i(��ж��_R]�{�{��v=]�h����n��G?S���²gB�8sfX�<�]z�4�yΓ��o��ԟvOs��ܳE���뤳͜���c4�];+3�tYYP�O���g�v2��,uL�����yA����7`�3�=me^Sc���}v"�YU�_^�w��X8� $N��;����[�:Y���o+]�����W"�nZ�כo3���v?IU�;�wk�\ib׃%�Q��E������Q�8�{|�Q�b��d�G#�2�쭪���������z�܈~�x���H{�!�	nT>��X� }�f���w}�;.��i���_c����*���/z�o���o�u�[�7<�.J(2J���Z��պ:�Uq�d�eKE���O���Q=��~Ӑ�#�{>�P��g����鮯?e���fk��U��2��}P���Z�V9w�qW>��r=3�+��HҔp*c=nT^���+ji�XgL� ������D�-�|e�����7� �_��5hΜ���w��][��1wM�{�����&��\N�g�F����A�����D�%yMV�x�3����޽ҽބm����r�>�⏞���B���О��2gu�Jg�1_K���
2.�#n5aW7�5�:c��w#��~Wrs�|����Q�l?]�4����2�S)tˑ�oO�U���=>T��m�#՛��ײ�?:�6����=��}��X��T�}�Am�9���cVR>�{�������*�7s�>G~�/���\<��]��>��s�_����)�ߙ�|\��+��t�J��(����Q�cj��N�����5�f�fzPEۗ%�W'T�ʪ��*�!nT!��pC��>����]�L���1�*�8����}}��v%tW��֠��+��v���v�t�%���:7s�n���-��b 0�\��`��%�@��6�]>'�F���q�u5�0�<o�0��%ޚʽ	D���|��/]�����M3�g�㳲�/������V�_?�9}��/E�b��.��nĬ��{�CЪ�������47voLw��҃'0w�	�,_�Y5�n+��0��v�6]oEk|�r��L
����#�_�Ͻt�{>wHwy<+;*t��Y>Waᵫ�N�F{��N�^���w�ڻ�<�5��b����~��P|�1�����i˙��VV��Ga;x|O��eл ����,�kwp�z��#}#��F���N}�u��.�L,��羛����4�/@6N�)`��2���P�莺���a����{�o�=��	�_��3#���I�`��A�݉n1Ƽ��dA�e�6
5
U��R�g�l���|}�R}[5F%���.�J��=�����ޑ��ި9�a?��f�P@HzH���I�+�v��ҫ��=����k&��+щ�d�;c���ߟ�������O�'~fK( ���I#k���C�>�/n-������:�6��Y�<��S����ܮ�0t������$Еش�`]�B�ڵ]��(W>b��87.�W�26uGG�1�4��K��z_n��pè��Y<�8��������M���7�khІ��eb�@2K���Wt��-�z�2�Y���Y:�3��R'�Ӂ�oޭ��_�&�ϦT��:&v�-_�^��u`�C�⤉�T�ڹcf����ͫ���R�=^ o�:���mt���|�7�k`��϶|Jf{��*pT��E^]/��K�q��q솪�^��h�C��	�ۃ%a�������2Q�"��Ӂ�EJӢ��_�f�>7�;ˇC���Y��؅�V���j%Q��X���(�i�7|J��\���tZ�\O���H�3w#O����;�/к��?W�F|��;�������B�{*pޖ7l�/A�0ז�myM2��3a��S>�]H� _^�~�{�;ԼZ���=�l��T��,��Y���]V�:)�鲾��,���B�J*"ˊ�L��k�
�M�$c�^���=u�qy�	\�q��y۫��fɽ��z�g�N��F���um��;E@c���c�M���;�L�w=��zR���~�y�����LX� y������}SND�z�V|;��f�=��&GG`}k�n�T�~������K�{N�f��败S����%�jx�ê*��s�?]ke(*h"�H�Nd���������;��2,�-RswO�.wv��Ik	\�;������./���渪��g�ɐ^��d�RԾCW���*\���g�o�̯S���7ƣ�{�E� �,ȱuҺ�ȅ�R�f�ױ��޹���N��gO���{D������}Cǭ��{���ø%�GĕFX
^�^i|�U.ΟZj=���2}	]D�^�:%�^��{k̭�P�מ���N����B"�� �ɵo�׆'Vq��4z*�n6g��u��G_�D��yb^W��~�M�DmǪ�����g9�W=��.}�3f�.H-��q���a��E����9���x��ւ�g��3�#�i���t��@~����d�#����"e����t��Ћ�~�*6����H�Q�D�f)�W>D定z���>�d��z�
��9���Ff�*�R�h_і�q�J�n�)�������o���g�s���������f�ǽ>�އ1{�O��(2{`d��>��ލ��O���]vz}z����w�,o���c�܋{���~�=q�,_{*A��|J�0�����Ȭ�>�����Z��#﫩����c��p����Ng�^�C5ވ�^	�{&�w��f�E���MX�TG��L��tWy����� M���n�X�ͪ9We�F�)g�>	<J}Z�b���n�٣i��.�v�Fa�f0����Ƈ�>N�{3t�(����\��`vsK+n���*ݧz��g3ڻV�`��XfE�	�Tj�GH�W5��u�[ۍd�|e��&0�'&��_�B���s.��L�ۻ���:Ovi�M�y�SwX��n5=��t�ٙ]�8��k ��6���}�M�ΞiK�V�/v��0k"@l[)VA�<�5t-��]+��b�q'-C2��uJ�\1l��q��h�⨐����Y�y�8+�ܗwj3ϼ�|�F������;t��H�M� �}DfrU�kq��]J�F�G9�r\OXۮ��k
���O:�-��J�;��go�L�6�.�����`��͋l�^7%�}��[ok{O\W���IL����u_RI���D"��VUo0��tLc�U��u�b�{',Y2�1�6�N�h)�TC�}t�͡ ��:���[��P#3^s�6A;(�
#�[��	��K-܌�j1b�[��mə-�����/N'|�n$odIv���O=SR� W����6:]���ޤX�K
n��(t�F�Ma�� ��A�t�-Ny�V=�XI܉�<I��
jzr7�x��gtv�"k����`���K��Gk�����%լ�Z�Rkw�c �9�1Uz���:6�' L���Nk����������R��#0]���2�\sC�J��_u�
/�ϵv�����G�:�et��s��')YJL�YpXʛ�;�R���O���S���q�E݊��جj�J.���/i�j!���o+�eb��e��6[5o�S�ͼ�2�یZ�ݶ���w�n�#�}����M�e>��Uۅ@�A]�`x^�oi\:��� �N{�n}"�LB�-��Q��x7��n���3�� �&ud=�j�>�*h��\�$��r�gL��+W��9YgS�*&=)G0�%v�r�.��Z��"���3��]�3�e�8�r��\���-��m�rG�y�5�I�6�Qf��=��<��$/x^�D������
�,�>J?.�Z����P��ym�$z����&_l`�h���!��d�U~�-U�:��Qho���ZĢ��gϨ���R��ŷ��r|����g��-vud�؞���Y�-4ֵ{q.��}n�+�����wEJ�>t/-�X3r�t+��nJ��Y˥FLdЛ"��Z[N�
�T����y�6��ߟc��뢯*V�s������7x�چ�rX��	h�.���s�W��tK�U Wº�j R��]��JP���{7���M1K��e!x�w
���z�b��G"���=�#��ԏR��J�邶���%l�0��st��l��P�7_[i��»�7KY"j=�����t���}b�Po��߯�������޼����뺹��r��&71��n5�&Ƃ�w#c��8��.n3t�]�w\�ܫ��I�ggS�75ҹ\1WCQ�]��u�!�s�p�s�q���9�ܝ��rNb��Q��.�@w�ݫ��ۮ]�n�.k��˔�wQΥ;��HN�WwI�n5�G1�r��].sE'w@E����s��7w��+������幸�1N���q�vP�@���N��m˻��v(.gb6(����9�b�]p��Ν�9�.\�擻q�̱��;�\�]wm&D+���:�s�\���$\�6J�3�.�ؤ�n���s%�h�;���s\�S��W;.`��s�9˻�)]wN���?�׏����;�o��z��O��o�<Yw��WT�i"na�=�Ē!�sxno�K�^M�s(�WXo��i`<��o�ګ�����	�����[���.����g����o�W���r�����gŃQ����.��59'�p��Xf �t9ɞ:jW�Dip:�\{R��2�.�WΏ�|e�s��q�}���Y��Q��΋^��n&Xʁ3�uO���4�y�}�>�]0���=g�3'��� }�r���Ͻt�yҨ��X�W��S��'ˠ�@�.:�D>�s��E��}[hr]c%�+Ⱥ��O���q�cC�{�O�n��r���I�d���پv�ȮO[��"fz8�h�8Z���������DZʃ�n�C��V}���;���=��Ǹ�<Q(�p��b�竧�T�ү�I��3�6NLo�R�O��}���O�W��y�do��<�����-[ӑ����~B�h�@6O2 ��~�>`7^��e��w�qW>��r=3�+�����EO<}�U�^����^��#o�5�4�Af����1-�qe����#o� ��8w9���F�ld����W��\Ϗ�t��{����Nd�7���2$�)�+t�z*r<�N����F���J�"�rj�{�D,�]/֮���k�7W�=U�N룻������k���=�-��zO-�M��Җc�k>�K���s}�����_�j����k�x$��w�e7ȃ;�m2�������*1��ur�iվ�� �h\���o�z��yW�����A������&����pe�w[�2D}��^�Pkѯ^���Tw�kЕ1���i��>�����@�~��iK'���z�G���y�է��H�#ncӽ[�6���f���5�~uro羠=^�x>��@�!�{B�k�<����*m ��m�A��x�P�gg��n���||��r������~�Gz��9���p�c�n����5ˮ��5�nX���ˈ�`�G%�p6t;����t��9�/���Ǘ{X�c�g��
+�wJ�4��s�&^Ǖ�O_��5�fp�>;;s>�N��S�t\U���~�F�������y��� �z�G������|y?U����1Y��p�'v�����=�x�꽆���߫O�W��T� �6X����z�z���|��9'�FvT���LG���[齬>�]ΩR5��>�>�ۈ�Wtn+�@7���b����~��e1垻Còn���yf}�c�2�4�>������If��hʨ�Q�Q޹bY�n�|;��9��G���C�O�����������=��N�G˹�TEd��4"�Z��[��#%=��[�g����y��v6j����,�D����N^���?u[��΍��et��Z������+�;�F���Sn�
u�+��1�.cY`oJ[F�i]�3�������z�����,w��`H�w�T��k˩�_��_��߸��q���<��ˍ�ķ��g�ސ�_��p��.��E@�`�~
W��q���w�s�8l�_K��'|�s���z|��Fyﭣ�w�i��Њ��G��۰��g���I��L��GUa�UW�p�w�rw�#<ƿZy�״���������ꉯ��� 7���g�HW��̎ŁG4Lz&�����<����oz���?;`{҉����N�z�q*5��ؼI*=���j=53�Fi��/��n!\�z���p�oɊ�������z�>�� 7�ɔ�
.7?�ڶ�v+���������<O O�§K��Wt�z�%/�?eG��1j����.�\��Mn$��r&�����|=�b��&J0ʑe����iѴ��)}��>5�v$ﮊW����\n_k��S�z�W�{��7��X����%,>����7S��Mqmҡ���� �DMw�����kʕn{I�|�xz���7^Y��;��<���͉�3g�K'v��/L����:��Ǹ%{SVt=\&X��I)�x�t$-��ɜ!PP�}��+�Ǯ�rJ�7N�ŗ1��m���dv׀��˭<�"�f�@w+��M��NĖ#�x��۽���[-����5}�k,Y�
�ACܹ�ʓR��q�ɒf譭Zʱ1Xqy�s:�B����+)�^�qu�}{�~�׾3�C�/�/U���xtg��f��	�¬��z��w,���kԧ{�N�D��E*�\EeV�����Yi�+~��W�'>��k��^t��s���v ��W��N�Ai�*���z&}���B������p<��q}^%2�}����y�9�����J�����g�1���zr�g�o�cv{&#�u+'�K����e\��ӹ�t�Pg3�RX}��/�g��{� ��{�qnH=FX�>E��U^.���>Ȩ.�U�<���8}MՉ��~2;��cw����=�׌8�QH����@�AEI�����ܣ�Z��S-�}S�W�EK~��^elw�i��RMçP�ez���أ5��nunQ|5e�'�f,L����^/v��u�TJ���!��yߟ��q���]Q��W�/��J9��'�7>� /MArD�u��q�����E>B��?[g �s��e�ty����=�v���O�%��-�3,�Z;�l��"b_�
�t�����܅F�9T�0#kBV�b�~:'r\hJ�3��Ư�l��\�d�9���.mK�8�j���y2'h�ֽ<y�j�X]��9B�f'�gr��5���eH��Ҹ˳���<W����MM�M���1�7��|�6�K
K��+�UQ�W�&�-OZ�Ԫ����w��O�Nx�C��s2,���^�
�T��n�rW��_@�9~��J'���{�![����	���6}^MЪ?�8G��N�.�t�G7!��c�����.Ǧ��=�S�Y�u1��;�g���C�Hu)�|����ʐk�Ĭ[�OްL���{p��E�Oq�\S�Ҩ���Dr��y~	��K�Hf��{��dе����F�X�T���t繕��/�;Х� ����ݨs��D���K���m���U^�L�Lw��w��^�f?�.�7���3�o�<���ק*V?�Yr�����t���%��Qò�R�+�8N��[�z}���+�"���w�g��Kg��gE�/Iӷ2�A<G]z��N���Y�P�0��=p���g���~�ާ��}R�u|�\fR]��YP�L�l��P�|9��^���NFPh��]a�����z�VGU��i�x�=,b�~�x���!��9���*IRp��]6t=���Md�V�S\���w|eR�m�u9�s�Syb/z�-�O���P��c�r&炌��������+X��3n�N���w������y�|��}��h����Ŀ_>�轋�]�*Q�i��43��݃u�3dggz^�*���-��*��� s=�"9gm�Fb˲|���痹>�T���F�&��6x�<��� �X)(��%���'R\����� {het	)Tz���UD���{�&���^��=���nj���i�U47!Z�:��x���T�X6KD ��I`Hn��k]X�qߕ�\�֑��ۿ<��ewk�L�ڿb=���4�����e��Y�PB(�H�n��/ō�g��X�U�ljν�q�K������}�~g`�wI��Q9���P�KS�n:H!yM:!�n+�y�c���Oz��\G�Yq��c����A��y��Ө��R��&���ߪ��{�t_=s=Jw���O����\��Y	W��Τx/y]п�u�}��>}�q�T?]�>����Xʳ�w��<e�4'c�J�2=���*�w������޸|m�m�c�p����޿���f(V~Q:�*󽏪���ۙ�)�*��gg�N��/O��R��m��o�\y.�ȷi���u��n:�u�w����{*'�<�,!왾>�9,+����exmº|O�ޗ�s{Q�N��{%)��r��=�eo�zM{�y�{�5�̧�Ǜ-.?8z%i�or�������%�qb��?�?<�z�]�r�����sBJ��סt�����:@q|�}ګLl�u(V"�+O���ԁyվ�<KoȺY�쀺X�L��<*vW�X�!�=��|`}n�BRw+kۙc[���|�nXZK�����t���NH'����^�`T^�dxc�^�����V;��8�E}P�Jӂ�P�u�E�GD��<��tZ��t��ɭ6k�,L
�N׌��k��s�]{ǳ�t�q�y<+����K�+��v�VT�n��U��w����?u��7�s��>��}�"�W�ｔǗ����U9���Z�ٛ�++{Ќ��ndw��d�5'�ѕP�:�F��f�[����^ӟo�x�oO��P�fߗj�^�5��n��u�C�n�+��U
|	=Q2����P�:ꛟ��S�~�U�������V_dR�,�L�ߟ/H�|s��Hg�<�L�
+�*2���x��������r�دnߝ���Y�;t�_��hh����v;�4�{�;�Lø�\�iA*��!��mx r�؍�1��Hd�Ӟ��5��C>�y����Z�0%W�J,��t��s������"�T�^��{x�xވ���.�}�>E���G;�|�����=�D��=87�z����"���#�wi�"�茙�˸G���D����o�r���P�}�Lg�W�7ޤ��F��[3�A��=��UV��wW��]��x����
��6�����܍��b�r��&Yf�=)ebF~],�6pҼ��j�*�L�߳1	:�'�]s���j�����޷V�1�3;Kb�����j�3S�ۏ�FIhoQ��)��oea��8c#WW���`�JLҖO
�2�n
����yt�z�%/��?mǲ�W��1�\���i��l�}�y�F��@w�=�=s'T�*k��\NqR�轷��V���=�^�������n|���'�0��.������^ٸ�>�8o�>%T�j�և�:�uWs��5��Q��{H���C��w����\(}��{�V'��*!{*p�id��6܃���"f5VDʓ�3�7��!\uoAy��'�����*�P�{�:�KůM���<;+���-����k���.]~��t�ۃ1�5��u�Zn�_�Yi�17됡ܯzNG��_M��z�E���y���_�������V=9p~5[�Q!l��L��reA��q���M�w�д���ܖ���t�y�׾�e�eg޵qݟ{-
Μ��}<�:O��鱿�T��ayw�5���ֱ��
T��k�+j��z��7�/NC���u���H�F� �����X�LW�Ǽ=��ͭ��^�����fT�t�V&�����ޏS����[��g�o�Q(�>$��&�<�6/~��ŗ~�k9�o�й�ؒt=��O&��/�sc�+MƘ�;X)^@��a�F�0ٽ�ކ8�ZŰxK3��9�4���Z��r�G/	y���)*���V�yn�&zxt�p*n���R�f0C7Ln>���/�Ǩ�l��U��V+�������Wt��|�/jb}�~�.[��^��<�;�4����:�f�$Q����U�[|�x���7�a���Wq�+�����q7>����:���q9��@�.Hʱvϵ�[S^"��\'�.P 7*�����Z>��r6�
�O��ٔ��H7�K�9Չ��o؏i��}���{޽�9�5�%�$�G:_�
��t��������Z����&e$GW�VmE�ܯ�}��O������
��9�3ӿ�^�62\��\��ÑY��E�nj��{ݦ��>7�R=~��o�h�{����Sic�#�%�G��v,�������2<)5���Q�Rc�>N�f�R�]�Ʈwz��w"�����~�=q�,_{*A3Z�nn}�s��u�#�'�2c�bwL;�U�nϸ�o+��yח�'U�/�#ƹ���*Ε��3j��{:�h��j�V��q�)��E�.�EG�J!����t���W���靜�{�E�̻{HJ��M~��f��&~��v�-{S�`G������TTFC���x��ؒ�p�ڗ�ѝ w$	��8,�U��Dɫ��/\����[��O8�0�p�BE��Rىv��Re�ޮ��"P�e3k�v2�E��OK�.�]vȶ�v^��䑀f��Ԭܚͫ��:��}������^pS咉�IT�/Nt�_�Dw������d������D��ϕg�>ɝ���t�,^	�
���xUW�,���J��Hr�����>S,������~=���vC�F3�gMO�c'm��Џ0�/����䎏;�to�P�y}V}���E�S����^�=����e,�QS5|�]��"�y�~Hu�B��VMW��E��.鼱 /z�g��3���=�����+�{�i��OUOvy�(���'J���8|��]0����{j$�O���s޺�MN�˾��Z�u�c[���yQj��`�*��<��K~ׁ��-��hj+�~W�y1�7&�C���.��ya�9�eq�nF�y�Yq�f��,��>�'�n��/ō�9�&��v꼣ޛI<��M�<;�K��UVO�ZG�v��J{����v�s���n�Q��8�*Q��h�66}�O��rhz!ڦ�hs��r�6�W��yY��>��/"�2�19�:b {<��Ǚs� m���?W/^B+qM���+�k�Z��bẩ��[�F�">�菣m���խ��-[j����m�[n�mZ��[j���j�V����mZ��[j���ڭj���m[j���m�[o�U��m�֭�km�km�m�[o�Vڵ��J�խ���mZ��[j���j�V��⭵km��[j���Vڵ����
�2�Ι� ���������>�����	������P
���&�T��IPA"�P�6ʆlR�"l�q]ZK[5���D%��4��lڳ6�Um��kmX��h9��e�t�ű����kZ��d�V4��d[T�M���l���URZ�M�����! ���Hfe^�H-��Zjw9+[��tF;��$��dv��j�m��o z�:�Sw8 � P�`  �   /_p}�>���� _��n�\5�x �;{�B�eP�a�7u� ٝ�Ԫ��t�u��e�QΚ�նm�F�< �!]f���[zYú�LKX�T� �wajj��́�tZ���t�� v��h
hW�F�tHw\�4�Mr5ѡ��:�� h&b�l�e�;�xz9�
�a@��
�n�R�� �`i��+�Ws(
հU
�S�I3VZ� ����a��܆�;���(f����l.`��s��th5�cee���������ݍ�]�tγ�
��t[Bn�v�s2��-GwU�jշn�J�x ��A[�B��*�` &�.��w4;1@�eu�E�m�؛-U����Vy�5�,�2�]3l���9����;@��w�PP    &*%F��d`� CA��S�)R���0&L ��&`M��LMIUT�I�      T�A��J��aM6�� �0EB2h2�CD�Q��4��mH$�H4�J�� `�wT�q�Ö_�p��Rm\f&�ب"������tAU�~p2 TU8����8>�LDU��WU����c�?ğꡒ���HbK" ��I d	��(��J$ T`!�"�x���]�Bןo>�L�Ur�.��	izP)�İ2��R4x�D��ϫ$�BBIH��׷�(l��(<�5����\��e\�-ݛ�d�]m�Ь�ݻ���	�d�:�흣淴њ�[�]��6��A%�\-;��Ĭw۫�e��v;)p�PR�m��Rt)6�7o/.�Q[ݚ�2�ܫu��&�E���*�"�ıj8;� �w�	HfEۆRFv�.�i?�]:eN�^�2���Ֆ�s,p+�`E�R"�R�]�/z�#��l{�Z���Z9 N�p�ZA�oI���f~���r�w��՝����zmiw���XRV��R��P����m!�&�X����OW@Xz�@r�쿠���e��,�<K�Q���6ݒ�V���4(L�E@����bed���0�Y����]bv����-n�}*ɣ��d͈6;�êoU��ɈK��І�w��E-L��*���!��K�m^W��x󃍗z��Yt\�9��N���v�ŴN���76- ȜH�AnT�-oo\�`v�k�i<�f�F!�;����Ȯ��(m.�:�@:�����E&%rpЗ>�V��ޢ�1�H���_�Pl����*���3�;�<XqT�(��w�5�9I"q׼&�V�=�M�,�2���sh��<��D��eG/G�Ĭ���<Kt����U�c;Tɂ�m:��qf��
��۷�~�S��pF���$�J񽷘���Pp�Ye�C�,���r�ے�7z)���[��lΜ�O*�c��2����X4�V��k"�Zc��^��0� ��fM�.��w�JHʼ'M׌�yf;��5�,�J=s�A�����h�*�=N�m��|ޥJ�U	WiA� ޝ��^�zr�R�5v }��|h`�6=pl���"�����B�ߝD-��^�H3t���V��JY��&�*�s�(ލ�Q�pl6	V�r
�Ot���XݾV�=��x��+`&�|�����{�2,#`Ç�wF����3�)�YJ�΋�5��̸^�;�vĬZ�L�Oi���fQP��h�mD+U��QK�/!��m	�	T�5:zML1;U���G�Y�� :�a���;"P�z�	캙��ZBv���,#�Z���éC���Jv�?#��H�N����Y�V7�/ꡄfA��;V�lΧ��JÎ����w��T�K��V�Q�&��^�3�/L
՘D���#`���K�f%P�.P�Xn:�-ʄ��\
\&`��C�lɬ֠�v�I!س�^B_�O@(b��n�t�j2�����%�	^�y#���5��I�:rŋD�{��Ĕwqk���I9��ٳ��;1���W	�Q���G9 ފȍm��ڵ騍�t�s�&H�/M����L�Y����ͩ�H{�*����lz��MbE��h�R��e��V�
��b����ܢҤ�y=|�u�ώ|�� c�^Ð���Š��l��̻��.��w���G!5@���͒���(�V��S��!�{�4��Y|N����F݅{ًk6�7Q��چ��ڰ6�w�D6���Вy�(���v(I���[�H�/4���j���U`�-Ț*�-^&i��A�62��y��SԮ�a����[��67;6&֛�wz]�Z�"lY�c%+�	*�G�/) w5�R!K.S�-'���/F�9UV^��&Dʸ���46�(��zR�q!��mu�Z*���Y�U�.�k�u���A�9��a�*�#V����%���-S���8*��B��h���ķ�,l�ӕ�C{��T�q�ع�%.v@���m97�,�د
b�pB?�v�]�Fl���jhZfU���u��K����H�T���UY��X;���?�W�>yw;���H�-��ޘt2n�ܗ(�� �&Pz2�6���M� .����Tm���iD�G�H�6nؤ����vs�7U�sV��	+pe2��/~(�xq�X`p1S^��R{�����6�;Uf���B¬y�P�(-�_S:b�X1�{�TU��Nmc��X4L֋��؅3UN�n�oES��������2'CE1&{���9��n�����5$Yo�&C�K���b[���n�����M��L�'#2�q3����GDhD����櫙U]��_mH�es�x�z$�,8�uע�JE��`0rJ�V�9W���6�8c�I�Ob,و���5V0�ohwl����
6؆K��s#w:�dNS�@�s��!0�oW���l��x�6�:� p��,k��&=�mؔ��UJHT'13/\u�6�7 ��slTv9A�r���QQ�S4>�]��7��x6�4[T���mf�!�b�4��ɶ8��!��^@�0ƚ2�e��N�M-��W�Gݘ�سyb����./��Ň�`���8L�?8Z�neAf�»���E^#��d�X��f'�i�8��.
��o(P%k���;�x�|,f@D�S14ux����*�n(k��Zp��G��gQ9��.���j�;bŤ�㘳�����U@�5�-m(T��GU���cvŗYr�������8�1�c�1,rȩH�]Z��ͷ-`ދ-z�bk��v�wce*yf��Q���|q��n���e:.�Q�n6V�[� ��,3���Z�#�l�UXlm�W��ua����#ė�]�*Q�g6Ѝ�m*��i�mky����,pq�Q�K�q��bIW]�e!��i���`��ҎPڱ���`Whf�c�n66m�݄Ld��%4*P\z`Ql[��e��m���?]��K��v��>�	�1��r�����|���X��؍�X��U��8sr��>!ӛ�gVi���)�\3Z�)p��baB.. �X��Y�kV���隫��0�m���v>��З'
�>:�)#��s�^h|�ж�%���-`婣Յemv��Il�J�Დc9c�{d��zV�u{�,i����:���0����a�5
�Uđm��FU�u㑌N�����IR4Y����5�ވ��R�ז�������`í�+�E~��z���`e~p:{J�[Ժ!㿻�E���΅&%�Ď|�s�m�gsof���jH�CZ�]W��������3Yçh�r���Ӷ��$O[Q���<�eM�Xh��^��wKd5iK(��F�=J��qω}���st�3����GU�R�f��d�sD�pfn�%e����V�}zf25=�wL���#`iܧ��	GwZ�J~�f���p]��*p�2W0�CPg�d�8��$m=Gc�7��5��kH�&G�N�������7%\:ԫC����yo~���`n�E�%�1n�F�J�u2�:�wj���S�"��^,�E�O0'���4����45l�ՖKxl�K�vu������Y�Ē�]�����☥#D�G;�j;fj����1��F�N�Xn�'*ѻ5cq�ҙ�:��hs��|Oho8�
�l���%���n��H��M�2�zv�C��{�1c�1[Xv�*�ӻu.<.߄����̼ ��9S2`�0���۾��TA A��l+%�wV��\Vr�	�־Xc|�P���|�
N�/��V���n�[Xr'�*E����"���B�s1��G���|b]�q�g��^��ݾ�IM 2���+бM#��(�γ׿k@�W��EuOuܞy8�i��>bJ'-ob����t�)���G�/�aH}Yp{��Lg�n\"�O��C��>_J�J,�X'uāܓ��Sw����o��M�U�5��C&\͟[t�	`�����WJ����D-ŻV����P��T�9���cU�Q&]���N' ۾N��!��g���!b�#�4�ɵXq��՗BɄK<k+)�4�����Y�!���H�3(}����A1JZ�\;��7U�p���K��Ǌ��a�e��~�����}f$��-�
�2�N���4%G�˕�og
�S�]v��I>�ՍН�2Jn;�[;�j��k��ę[����ښɇĿw�b֨6vy�B�������q0{��b�|{0����ʻ��*���%-'ٻ�r9�9��+�%}=g
���8IG����^�6)�9�Q��v�E6��=�Rv\�58�0�V:gmf�%/�3�]��gG/j��������9���V\G8���w7��ȴ�٦���*����d��W6�e��wp8ɭ_Z�3_P���mmgeJ�SI\�z�$�"�5Ѷ�m�˱w[ؔK��-W���_�(p�-�S)�Uњ���ʕw7�k�D��%�F��{�;D��74CeecP���c�h�>�E�� d�v<���3��iC��o��w<�����OD���?�C��g>b��݀��C�U�E��-2%d��������|�Ȼ�/,�ݜ�+ذ95A�J$Ŕ����@��.(6?0r�4�����}ˏ�Úw�����\S�9��f@��4��a�咒Ί���/&�s�nF��t�툚/^v�"��Q��cra�ա�y)��C:fl���A�˽#�����{‥/���ej��i��F\}6r�Ozq��D�!��n�D��]�=7�0:,�I�!�Y�4�ʖ)j�گ�jʢ���P^� ��ڽf�e80�/v5�F�����.�{%^ii�+H�^r�"��I��f��J'��6��q8��y36i5�5y7����.S�y�,r�R t3=�7K�*uW��i7�Ó��.Kz�͘�ۚ/$�>��vM��j�rac'�J��Պ���z����sp��H��t뛛��?���=�\�J.��08���;e�
�Ju镗�i��Y���j7�vv(�|����4�&�5�wY,�w�<��H��PA��CQ��vb�f$®Cm�V���=�l�OvS����w؏\D�^Ρa$��<X��{�c��Wgcf���nk�J][�uxp��SDaB�{��۟].�u6������玃z��*%����+3\���ǾZW��B��N>���/��v�R���U\t�O?�ޱ覱�y��cы���P��|�+v�݁d�ݨs�̙�����P�c{.��F������	���˪f��(n]W}�	;n�q��nW����˴�ks��e#�������k��ɩ.�+� �!����(�z����T�n��;��)L蛱����{z,85��f�̍a쎭G']�o�A�S��h�`M��g1صT��hTze!T��
�Vf�܃�d�ϴ��*���Tfq��HjY�Y�k�?-ND��_^˔��]f:�$�/X���3�w�lFuqy1�|_���7XAS6��y�W6�P,Q- j��5;kN�9 }֜t
QhB�`�e��ʔ�e�<��]��kj���U�;P�ٻn�*s�Ka����z�<�N�5��J%�LH�"u���6t�];��:F��5ُ��]A��*k�j��
�Jq��:x�f�%��T�5`���p���\]i�[�sU��[T^To缓�x��+v�M��{k]�Y2�����,��X>EY�gbӯ7�HN#5	���B�z:U���Y�"ǲ��ފ�Xq��
�͍�#aϫ7[�*p�w�+e�nA�s�� �fاoV�Ď�
[e�[��]dC�/�)P���9�-��ߵ�ݠ���̋	�\��;r<.�IY����y�E��.���rm�gt/����ۣƇ��ӻ;��nl�n��EuF���C�͙]n�ݘ����X�:L�^���?o|h�W���³�!����6.����1�[��Vhv�,�HR�]�i��\h�J�6)o5�XWm#����]�IWԕ�׍��@�6-��bWZz���]V2+���)��W�-�l>��寢���hy�����}'��C�yf�N�H�\\x������YƆc;0wa=�zr��o��Y�f�pں4��%ٝ� ������}�"�g���䓙�勵E�9�O(��t>Rbrњ-���2x��%�uβ�k,l�ʹ��N�˘�_?�(0f��`����Z֌L�ԅ��f��
q]e���۳Ky�oQѫ6��9d��L��d��Dz���0�d���E7ݨ��g.ɇ�V��7��ͧ��tdM��I�O�-����β�ܑ���J�ɮwH�4C������vr�Wш�͝dbc����Ճ��ƅ-�4�c���d[���x�\������~޲S{���l�0a~SwE�%�B�;|��_m��`�0$����h�q��Sɽ5:Ƒ�mE#͘�it� 5IY���6T���rvڱ�m:���z��_O$�r�l^[0���3���o!\�Y"�7��E��t;Dudv�b�+��j�S�z�t?+�vwNv�}	�g�wN�`�D+,��VS��Lt�g=����6����Ό����+����fK����F<�:�T�n�2{$�b��B�ѷ�IA����s-��l�$�Q�ͨ�^}h�+u��G@��;���i�,l���U:�h���u���Mg
aH�uh�JŗB� ����W}�0To��1�N�+��޹һ�κMיs��KT�픭q���nY�q�֊�-���t��z�N�hti��(��c.#['J͌!�@�f�$,�a�\/'pȣ̭m���)2��F�"L�#��2�+kjJT�r�gUq�Fk�ݼ2' 3`1+���G$�I$�I$�I$�I��#�fNs�9z��<�a� �\2"T��sy�ܭ���90^���:A��2����N��M)�u�]���e,gN}�ꡝيV#0X�Fn�*���駙a]�#B����\%��{)��P�N{\(t$��^^++��r ���t�֛���R���"�Y�X�T쉹� ��'%[��{��_"�/,�#����n���������ڎ�n�\(�2�k�M����
��N}Go��]/w�8����SJ�����1F06��/�m8�]t�9��efT�L��?h�b�N�/Q9���:am�����}�m]��
�i}t��b��5z�U0DF�H�*ݽ�fcH�)�,���7�.K�����"����g@�T�JA���_*_�m`�sn�X����eR|�`,�X�_��o�w���٦�ن���AU���֦VTP 4�TBj�8��|��
�Q�C���ۦ��֤�oL�y�"�iy�V��M��4'(�q\��^�u�3�{�4^ZAj�w��;i���|�-B�n�v���֘��o�=օ[;	]�tU�k��@�i�۸����o�`�Z����*r`t�=��oN�U��vF� r�ö��N5[?Zz��k���*�d
��ŋ�$�o�:(��F�Kud!ӱr�I�w'Y���;5��|�5���R�cu�x^�A)/��p���hA{g/Y���CȺ�n�ճ�qh����i'��L1=��
�f�Ǟ@���f����'�S���AS�cK�ӌ���[��x��
�0�l8���&L�)�Gf�����S&_s~K�c�5
�>�����B�Թac��~�z���I�@�G#=j�������_+� G�&�vv���y]r�o�D�-�X���J�&q�coo�O�w��GSg-��gL,�\:����.̊\��������d+r�m}�}�x�y$����|�2L����{7��9=�(�<V3/v6���x��TԜN>[�.,j���l�,z���5f�Y�����H���T����n!�ﻪ�T��u*L�$YF�A@0ϴ[1�:x�Mt����ZB�!h�*����`��mp����Rc,����[�h�n�űv�35�&#�1lܙ�����]�4��Y�d�u&*�6�WK�>�� �&R�_����H��옠��3u���8*�k.dS{���T	��_}�d&�yB��d�2ݬ��H:On;�:-Ўr�7�<�mH�W�Ku��.��F���U�]ʺ3p��=�Y�V�WW[��.�E
R*����}|�|�zR�gN?{��1�xh�Fgm����WM�Ŵ����vwo���|�������a[V�.�u�K�dc^tOCvf���p&�rZ�j?�^��y]�x�}�&��ek�T��2��z�쑷�CWnt6R��TƧ(�;��#�Wr��v�D#��z�q����W"z�)�3P�q3CB�Y�S���䞀�,�b3QW��f4gL���m�]]�k͠#��N��+�V�`�ݴ����!gp����3L��'	q�
����6�	qYV����6�JeL�)��#ZÞ�5��r-/�&����){�Lf�]d�{,�n=�a�_��ۣ�&jl�Y�j��Qp�e�a�{m�%u��G2��=}ZZy-u)�S��n��A�4\ݘ������b�n��GI]g�-���M>Y5L���nS���[Vۙ.P�����"���qD�bԁEi������7�uTz3�_s�T쉶3 �{���q�y�
65N���t��d���N��,�	9��dGm��B����(,�����јi�v���٥����,�������"�gWk�Jy��	��{��`!��^��
i�3�NQ�8b��Iܜ���KM[�s._J�тA��qA۔6��a��v>�C���p�AGzg婿\'�������pK~�<�WT�)�M�Z����;�kÜ��=��hS��xu���D�H6��O�f�'9f4�m5�2p��¶�L�r��-��I��ؓx���R�v�r{�NM�5��Eeh�~��]E&�*�r ��SON,��v;`���Q�����ӓ^25�
:���7x�kś��!�	�bb�,]�/oKz	êa���w=�7��
|����\��׀�|�����cp��)J��CP5��qLP�i3�.�{�����
�F��9���{���r��*�\3��j�$�<"+Vņk���I�z�I�f�W{���a-swh{�y��IdtuUR�mUoc��\J��;���X��Y�]faec,�}�C�=|��}�N<��T��2�OnLY�\��5t��ܥ�>3I|4��QS�}3�>B��Y�"W6+�+��B�ɕ�;%Y��;s�=��Ę6't[��(�Pj��i1\&�{}kJG������K(�(fq��}Oz��ۮ�C!|7wne<��m���N��Vz~��~���`5I���٠�~��kn�������l���$�t3���b��"��.h�ƞ�
�_�9Ί�2N�:*:���L멉���%����˺ѻa!3��|�*i�NoGY*H�%�}�3ɸ�;v�u�ީ[���uv��|��Pk"k5f�u�����.����/qBh�:}اG���=@�l�7t4p�¨�Z8]��ǅ�YZ��1�n'S�򄎨L�E"s��y�1��&J+k�ܶ�Y�Ƭ���3�����yf�>�kc�׽7![j��_���KjE�::e��tjdJ��.xT�Z_�X���n�h�of��h������^ ��t��Q�=)�+��{��e���nu�>]2#�k�;��<WI�y���e�H�,$#g&�y6��3���,g3V�-�?M�F��%��_j'c3�m���ݹ���!�ܗ8�e�_����4���B�m�/��E��^������Ҭ\��w��nHU��M�yV�ͽ��MQ��A���x���4N\K�����h��t��|p�I�[�K��$[P�
u24��]NP});����S���{ �]�5?�E���6��I�����l�C��q�(��Wa��]�/�Q�=\���5��%��QxG��Z5��S��{z�m������0�]�������k�
Ca��Ti5��K�K�b8F�>��Gr�VFb�=˗�W)]rf����M�	Z)<]�n��diYR�����KTI$�R��,v�i�ǍV�:1�BVr�&д�i,�^:�,֎e�l��2�j�f<8F�h��e�R&�|� WAX���*[wc]��v���4��a�a��vZ��ہq�8T�9_	�QPt��e�b�dr�)A�`1�
�5����H�AmoT?K�ҽ����ԅ�Bʬv'szN���,�j�@�CkRP2ɧ��ȫFY�xH�\�8��Q6ӹ7�5�y;�(W>��E|a����:��ʐ��AOl{+(m�����1�X��.j��*�%��V0N�lC�k�1��������զ��m�����:�*��U�����U�[�V$˺Ï$XH������E�	��;d��C2�yb�6�@#չ�c�ѳ]��JGCQ�w��ڻ��ZA�*�fLg^�;�QxN��go:�̡1+�pF���UX�[c#��9��Kn^���8�O�k3�v�%hv]�*e,�l8�j	5��5�&n��7* �u)X��e�W!�lM������
O�*��=[���b�E]�B(a�9{������!�GuL+��Vܳ[9�8�`���Op������OM����N�N�R�����Ju����l#c-x���B�h�bU���Va2+��5��ވ��_7c����te�!9\ս,�-%]��;w*�^w��UX+-gsf�v,�ٵ�\9�.�55 �Sؗ��"L{�|ڽߔӞ�"b�9D/�Q�k�^��C�	ū�|+r�ʗ��2��K�N��V�W��0�����}��D�MB�m�s�/{����1����[.���Cڹ�%k�wI����_[iV\x�4�7$Ǫ�wb�e��{j�|�H�3z��6��4�����ʥk�$~�v��i��t<��ޢ�+��_�f�0�y�6��o:~��d�$9�,L��`r�4��efk�]@TVkS�YБ �|h�J�(�/��L�{ڱ'mRk�#�c��|�	�F_g�"�Ov"���I�fձG��Vl�ސ>��zo-^+Z��訔���wC����g$�Ws{)�� �:�M�{C嗕1V��!���eì����ԗO��U� �.����Úrn' �>q"T��D��P�)wt�ff�P3w����S����+;�;e�B�V)U-�{s��1Tt��q��̅���J&���f��eD�����(���*�ʴiQ������գb[s
86��mr��E�(��V��Q��E˚�G�eeDE��0T+�D��V�wJ�+���Z%�Q-���-E��b�z�.�4��2���j�.6*���ecIm��ł�kEbF��Sb�G,����A���H}�R���8Or_���%�vQ1����������W$����F�C�"��6�ox*��G��~A�J���վ��Rc���+�3m����T;�bz��7\6nK8�$eѨC�2�K�z@�1D���J�%;�����n���a��6a,ђ��5���Dp��;
�׳���R:��h��/�{"�O���ʷ�/�n1D�Ƣ����Q��C.C�vC�PoS!ָ(�z#����W�e�'m9�Y|� .Fz:k���z���dD=��E
�u��q��|��;o죨~/�Sed��9��-uo7U��m��������&m�f+&���L�:�f[��S��zK�k���C����M�Ă+���s������UoODNA��I:�u��;6� k��S]�ie!�6[�r�����4ƹ٫ݷ%��;�p�7">��q��fӫ�kl��#�������N�W.�F�݉��U����>�q0���6↓�]��v���[o���9;0���2�7�����9J�I��<�aB��e��;���B-�e�G4�N��p�G�;��AfI�NXɚ1�d$ �5�ZPr���ꄏ����ܺ�i�T0�ŉ��䥈W�G1�E�������8�9��V! י���W�o��gB%G��gn����c��W�T;
�{'��ۮ~��+��o\�T���[}$΅�����c�V���z�nT&�t����_��eY띁�;8������!���}��Ś��ʇ�U�"/gsM���^�j�F\�5^���Ff��t6��o9�Ƌf���nw2+h4/zL�B�kM2B��Ts�B�4Z�˓
5q�G$;�tm��]u��^b�+���N��q}5�Xq�~���ۻ;eO��J�^#/���ʘ|����&��=���5�o�>���(�[r@��w��,{��n�J<㗜�RJ"T�Tq�nH��"�߯4Z��g�j\n��{M�u�.����(�7C/p@q��ۚH#�Tdt�>��x��K5������Sш9h�]z`�6yó$�;����=�e���g5S1��6w{Pn�G'���|�]������=Y��0(qA��e֋�x��0>���tTTGw0$_K��&��]��'��76�Z��ȫo�][�@���m���۠,�a~]\��&c��;�3�ۢ�+.*JQAe�%�+rX�<Ƌ�5���y�̭��^'���X+dU���)��)D�c��P;9G�ڎ>�ne�t_�L�Y��6��p����:I�h��g�P���%eT�y�mC���,Q��H�P�5ubV�8%we�lGh�=�3u/8 QA�\�{;K�b��q�|B�S.�z��^�y�NF�o������,�|�SfS�P#*ö�%�
���o �j$�zob�s�<���ɦ��E��,���j{����w����z9涔�TuH��SP��O������=б�j
�]t�Q%�,GXo�R��J�)靶)�Nb�:!���T67�Z�"u��.4sde9W�Ĩ3ώ����"�@wt�mT����@������Emq�Ί��2�b`�WA��*�ߖ���G7k���p��<@�����oM�OpG��WxI0_�w�K|���g��,�����|"�D�u6��i`����*�xF����s�i/\|e��c0d"]�.�>�O��Y>��⍝�I��p�5���8���h^�25>��NIZ�9t��n�B�6t�D;obQl������P�=�����uD�fԪ����1>�z ��vlX}%�p���$�2��c���&�φd�m��լt�5�39�Iż*9�W@LTB������L�4�6�#N�W��{�]U���O �L��Lh(�t`�O�{��gs4�m���j��CA���4D	5ߔ7)pc��ݡ̣�YF�q��N�Y�9ޫ)P�mow�c��#g�f'��*���P��d�8��eF#.m�9��\J�;��[��hpg��������!!�Z�m�>Z�tR���Vf,�u]d��,���h�ފ^�x�>f�Į�%�_7�Qz���ß]�|��_r�����	[���+XW9l�K
i3{���ݬ0��4�kvm���1H���]�s�WX�� ��4���w<�ɻ`��ʭ(/2���,�뺮��5���l߂⤹�+q�&e�.���$HX��`hI��=Z�pق�^��{s��ڭ���Ӭ��m���f�z�}�o��;Q�)8{_�������e�u�7���I3���y����5�+ΞI��ݷ��}�e�&m�w�*��2�Q�n�-x��b�3��هy� �U��c8;~�/��M���#�=��+)l{(�+��UIo��]��y�d�DU{d����VK������E����*bQ�\��$� ���4��;�u9�=�5j/�"B�����Q���W�,/Ϊб�4�_E汮\K�oy!s��:W��t�e�9���z�lrKrY�1A���fp�Y�帛d0����üҢ�6���WU���]�*����ܵ��{,U��)���jy�{�խ՜
�,�%�p�N�oDb�Q�]r9tg�1�7D̅��svb�O<U��V���mLMӍ\w�:J����g8x�I���Բ`Z'�\�z/F�o�7f�Ǔ�(�ݘ���W;�[�s�F�Y��In<M�3�j�"#(6�$�7��`�J/M1*��[��{k��Y�C���r'� �&ox]5m�cb5���~	�QB�;ܪM�]���6�����\U(�(W�����u8[i�"/k5;�J�;�U>�I�^�F���,�!b��xv$��r��ÉI�ux�z�,��W�]���t�,���y����x�#k"�F�����zǷ�s�Q��$]�v?O��d��j��WV��^���v��>n�0��3-�wJ�ȸ@S��Rڽ�c�Nȭ�1�wb�j)>�Yf�i\��o7�r�w�H�z�8Tp�v��u-�c{O\��Ț޻��ݥ9
[��-zb��N�ML�I���ޭ�n4�9Sop��:7��7R�i�0�tT�����S��-�HE�ɧF>֢k��S{33睂g]�� 9,ـ�To-����z�4��0�)#��~���)*7�������	>>�Y�LȫʽD��Y�bI�,ͩJv�/n2��z�B+��'�kRY7��xB�׀�5a<����Rh�|j>/�������
�r�U��������M݇��q}|�6�V=uA�0����WRK�c���~���&���_��ʣ,��m����,�A*C���NV���P�ѳ��9Jt�n�����3�{oa�S��06B3�6׼@Di�61��u�dfY�v �h+��d$��*
{^3}�CD���G�!�D`ָ
�&���2�{v�ɞ:yC��Xat�`��^�mn]2�1
@N�yt��
�.	�p�[���Ճ���"���B�+فh�,_*�Wۺe���;^�f+*�]�ﵚ�1-�;Uy{��] ys�D�˖B�M��Ѯ�h�"�}�	��M��+]c,�����5�H���vӖ���ؒnnS�H���ϒv�o`�I)5Ȥ�u��:	�����S���ǚc��J�i��^��3�{Y����D��~�M"B@�h)�b�Ne��4��h�uLn�r��E!�a�i�Z��X��H���UCHVi����1dUZ�X���AL�L�DE��bU`�m�
�
VQ�EDZѝZꍱb��EW�U�*ư�W�)H���AT�V1ejJ�(,,E�(���Z"*�AE �X��0�Q����H�`(��-�Y�Q�镐�Qk-�`��`(2ڋ)YP��?|N|W{B_����>�M9F��*�C\�3Jl��n�,��ek��G�օ�|�o`=�;q1�Ǯk���WI��ޘ��\��)���Z�%��K瓮$��	��7���|�Yn��A����׏����
����$�La��R6��Y��H�j.3=2�
��s��\�gMoy7�6#y;9�OE��mB6D�o�dJ%��ps,�
���3^1��*b�%g���)lM6*õ�x�8άvb���;.���e����qSX�H�A��p�)�N㈂���.�{�nt[�k���w�j'��!�[�}[�`��p�?����y`�h��NAS1�v�KIgT9	���2��)�#�*��
����|*.��9�6�u��ږM��yb�|�������f�O����k[������z��q���%�x�/�i���ӎ4$R�QfZ���镯�EtP�y��v:��Tr�j�.�H]�c�*��d$֞�B�env�zj�3�\���5Q$�[��T�re�$�5�j�V�t���n&`p�y���_�c�ezw*�	��EAilՂ��Y�g�xF!� }\�	��u5zVU_���RK��s��k_^����zI��P����S�[��%����orTi��}>� <\RwQ����^U�R�5^H;ד�'�}��d:��̗8�����$ƀb�nVG+��"��+w�+�f���d� �LW�kgLJ�K��@���c~Q�r~
xM�YÛOD���&�F<)i.w�3L�ع���/xX�����*��X����=@:T^�Vh~"����U���9r�H���U �Vb�tb�m�x����Q�p�v.W(t؊h���8���L���$^[��'ݳ��j�ܼ�z�)�^fĕ�fj|w���	s��;l���RP<����X�l:�
ʾ�6K�E�%@�$�Q�������Q�i�KM�1Y�-�:#�K	g:I��-�:�d��F�.y�]��L��i{p8��]�Gg{N(��<B���0rb�����FXmlK�0η7Gf�k�>0�bw��e�q}��P<E��Y�mR��AG}�d���H�svB'G�'���������ֽ��s�&2=$XAM'̇��=`(s�AI�z�۶I�t����Lt˭�zh��s~}�8Hz��������Hq$��zyN0��>`(t�|��I�I���s���y�{���И���l=d��\�=Bf��4�4wd>d=zI4��!�<OX
��B�tɰ^�w�Үw����z����NVW�Ǖ	���ݭg�᫐%�;jq�??z�=A1�p+��n[h�-Wh�%�fS�7��e8�AE'n.%/;���W��RO�
@�m�$<BsV�zɯ����]��x²LgI���u���Ͻ�d�'{���$�``����5Bt�04[<H
a��;��!�G1S艘Qs�D�~�޻�x"�C��l'�v�z�x�q�$:dP�!�!�i���w�l�H|�=����g��˭k�=��q&0���=a��m$������d�{d���$����Z2���-=d����{���V���߾���P逰6����C�O|�~d=��u� m�HC���'i�E��^s[��]}�<������a�7d�I�P��>Cl�d�(v������k�ߘMn��b<�=�F�/��(����(�4�d6�I8��R�v���$* m����$�$6�w���je��m��������ߝ�ω6��|�!O)�<dP}@�'�R�>L�"�z�2Bq�z�Hz�o^u^w�������L&�8}I�i��P�b2O��Hv�0����'�-����׶k �Y���߽�3�y����w��@;a�Hz&�OP=`VCl�Ch|�M���|aP�<d�'5Ld����s�y���;��}��[��ɣ�+�f���f]Ǫ�����Y��9�/>���{�5���j|���++�uJ5�qI��J�jQ��s*7+����i'hz�/����0�l�d���{`��Cl״i0eI<I��!�E�f��^����������'��j�=$yB|�a��IR��l �3iR�>I3�AI��5��\�Z�g�bI۳�	�-c���C�	�~�:f��x�l��I���������3�k}{~����I!�',�~d�a4��������$1:N0�IߖCz��C���y��������d=Cz�d���2t�z���~`)��x����V�3�N����}��}s�}�;�|�6��T��6�>�����M��@�I��5I8����$�*m����n���{���R@�����Oz���ā��ha>|I>d�$6�RM�0�a<f����e���o�z��4�sWhm t��0xuH!�R�0�2|��$��OOY!�����^s��wמs����������N�OP����������!4ud<d����OlL׹$��O����:>λ���u�����'��["�8��0:���=J�RO�i���CL��M�$���ؿ{�]uΫ�?��Z�T�ږ�87�`(uL=k-��Z�Uo�V?��M19�^��X\Z>X�B�go8���3���@C:�^{�p�$��h�m�t��Htϐ�,&��$�'��Y1 P��
��0�}���u�}�{��C�ݾ$�$�VM�7a<f�4���x��ݞ�P���X��6�r�6���=�����>��~�c�AH���`x�d�B����	�
�m$�d�L�d�l>`}�}��j�����$�N��Z@�CL���$���$;�&�r��<�=Cl���v�o�y��Ov>���<���i*��	�
�����i&��A{Bi q |�:���l6��=@6ɇ[����u�s~n�O�`,&�P5�N$�3^�B�C$�������IYP�Y!�|�m!�:�����>��~��0�d2pJ�Ih�$Y>}@є!���!�!�8�<>�4�Bt��:��s�wӳ|�~o�rOJ�N�C�l0I�2t�m��O7@<a:`,=d��=��
e;N!=H���|��sa+!��M!��� ���0C�bN$���J��=d�OOS�&��q9���Y߽��V��1 }�hm!����3�@�3�6�Y m$ē�Hx��I'���}�:��Yٻ��Ϯ��m��Md��^���}��n!�]����RU�����i��`�٩�����{ה6t��!�+jAl/l��+h�޹al��-Y��!�2�r�`��L��!�MC�hq��v���
�;fЇ��l�2|���������O����^{��Bz�v�VC���݁�I�(|��d=`)��a�ԁ��O��������f�y��s�TD@�{�yLq�'�j�d_,Y��_Psz��![z�ڴ�j�Ȯ��6�������3�/~�f-��M��/r�1��X�#C��w~��*ڪx�6ʘylXK�p�q\�]=-Cc�/N�g<9Ap�[�h�V���i�3-e�Mi��;]E���U�Ӌ��B�a���W]u�\�^'S��j�n���J����_p����������v�V��rk���̮@Q�����Kjƌ�'>���J������3�ש�ߨ�|����I�Գ�Q�����l<����z!���TVJ��29�+��3;�ڋSnJ����~~MN���4E���O`�c|G�/�oJ�B�žB7�_�"H�x�F:�/tt)�'<�%Q����T�#��u�8�v϶=Zd��i�{ɇS�I�fW0;�+�iz����3��L��U���SCz�1�v���j5�i׍�X�9��\b_j�_=y�=�,��*�T����O�wyX2y��EP�9�p9�~ܡdT��ճ�3�d��d��:�� Sr���� �ą?C�Lo<�&��P�NdWj�;���;o!
��\<L
O���N �0���g�lW�MA�ޘjo��,�#Q�1<p�"�+�Q���.�<9V.��	��;!�7� �L�k������f�1:�3P"p��A�2m��x����!lj˸��uU�vY�d��	���n$;U������WL H�[n��Vξuk8�%�������|�i')��K�����3�c��I�ۨfe[ꆢ29D��ѕ{ ��w	���Ζk(Q��%#P�C��퀇ֲ#���l{6�oX7-�hT��3��U'Y�]��H��l;��@�7���{x���nA�Z万R�ۃ\�lnt��������+��O%��&�toC�(�ewm�B1�A���P����讌cq�6�*�0E���s�T�Jr�'�>Z3��p�
�4EZ�S[Y]����@��ڂ�hWWn	,܂L:Q]qY��]y��S@�4@{���;0P�Y
��:�v���?J�y>����>D�S�s �RY�\I�y��=Y�)W��,�X�ЅUo7AN��DFB�{�f.Iu�+G,<.�nƥ%t�70?.P+='��c��)�����>��5O�����&���8(gnU�Z�ֈ���xc�6}.-j���mʻ������ݴX+:��.��t��('z�E��{$3�y'|y,&.���M�ܲ)���z��&�Kx�X=Q(�n�x�LT����G��I�q{�[�Ϟs���$ٴ��|�S�޽� A!@��Y�����/�\N6����N:3��3�d�8���7
�4c���Kg��ל�4�*�g5*���4��{x!ժ_r�A�-'���殯3�P�6gZ����@A����Dyx)�	�*r�gg��6t���r�s5�}�������F�^�o�B�������*v��A������h����;�k)N�4�Y�sN��_��������V#"�q�VE"�1G��>JȠ�Ƶ"���D�5K1R�+�
�������B�dYY
�m�R,�V
�PU��`�,����B����đT��$X��@R(�T1�ʋ��DbJ�`�(�X,"�Q@�J�dXdYAF�,P��z<����o��g]���nEIW�ց	�Y��F�U(޽Y�)X9�H���_v��b'�ߋ��ߋ�`0�_@�*���oW|�q9^f���ǯ�y}�¹�T�6[��8j�*�T��Dl.Yˡ�c��q���l���a�L쐑����k����k�H�EL`�N����r&��%~?��z��!�D+�+��O2ē��U�o�1��1�c�'ьcA���V��{��N��\~�(�ށ){9�H\X�R�Q&�n<kbn A,�Z�+��gt<�I��a��~q/�C�.Y�G�{�����֥�"��o2�nVV܂��j�	�y����
�bv�ꦑɊ%c���O�Ԥ�E�}���I�?&P��"s�����7����
6[T���O�7��.p��@ �`���ٲ"�bx��ny�}��Otsp:ό{"rb�+q��5�ʧ� �w�EuVz�ӫ�'Vc`��"��>����s��ը���Q�B�,l���Mp�:¬[q�SsA����6�IP��*k��0<�s�r��(yN��V��Jh�Mh�#H���ѡ<�0�NM/�r�2{�W����������eB�����x�Z:����sn���؅31[r������U}��y?�q���w�P�*Q�Y��\�z X��E�`�j����,s�mH�����V��%Gd�]��@�@��{��U��Ef�yy�7�[����'qW?p̕2��G�˳���Q�̗�x�����-*h֝��]Ŕ�&��x��5S���o�v།:�k��Q�}���K{���N;޹Vv3��E)�m�{�%!��˯��ݩ�`c�M��<[�Q��,��mZΊk��ڷb<����$�r�;^�Y����+[�[�L��w6��-�[3�RAp37���fC�Z��w� �����\�э~!�5�G.\U�Z��6I�tD[o����ۓf�z-���Aܥ]^�m�F@�ݾ��.���g��y&�i�*&��x�8��/g�{3��X�ۥu�K;��*&���r<�s�/׎o����k�}l_G~�mFc|�q��O6�]�Y�d�z6���U��@�مx.�N��4�o��:�PZ��e�sO��o_W�^9� �w�57ݥm��Q�:�X��C��
�<.�m:n���{�l����wV��2����t���I����z��s�G�������f>	�k��_}U_k)��]��VtM��o�{f��+_v�Y=��"l���G��!�0�攝yk�tYM��q�a�ԟ�)�^z'�o�kq���)x����m�7X֩����b�{����q��+�"�=�H�>��t1�顲.T�9��o�6̲D��{ɆiGjy�0�d�=�e�Xi����g[Z�eVF���u�'km�-}zs���Gh��v���D��Y�U�t�������Wь8ULN�VHṱ����3�؝�M�´^���F8`��M�0�q�rV��I}�G�+Q�\g������S�r�V�a�M��w+�\f�j����_:�-�I{�ֿ|?T}A�/�;2��3�<o��Fo���*ԝr���z��<]d2�g<Z�)`�uExvCdv梶^.�P�Pbq�ôn�����5���z��5\�%�tٮ;���NS꼻���u�7�e�M�� <״^�`VE�-sT:��+����p��8͈onhA�)P�S�}��L�p���,�2�=�.`4�i��n�4�r�o[��{|(�b�HX�鼍n�dɋ��e�G�r�!%����� �=�5�Q���Q�!=�xA�����Q�_0v�רaf�sE2M��}PN��@���eR�u{͝�9F�z�ioV��CM�k"�<����R]�I^|�]�s��
ؓ��U�Ϊ�&Y}�C8�ɏ%����tD�s�i�
Lz%P(�c#4��66��}��&��ᘩ�CM�W�M���I�'ۨ�1�'hA�)Lm�,NL�xqK�B/�v��C��FF55��Sp�Kat����[�~/FZ�|z�Fk�d�y#8D��������g���W�����u��y�X��'�]��#qf�҂ȬZ��g���(S�0��	�sU�{}t���DS��cQ�WeW��R�T��u�a��B�yû�M���f�X�3������=0��V�~�6%���1p*�Ƙ��.hBU���X%���GRP��J9N�-5�Lj���f��ؽ��e�}V��R�@U��������ݱp��`1�����(㙖���v6#%Eb0��S:�?|2������B��AiwG���|L|��Ԡ��g3����t�:M�r~�����o ���������}������o�/7��W�K.r8�5��uQKJ!�/����,q��� �z�6�B�+<��V&"��8���K��\�#F�N�D��^6񎞭ٓ���N��v[X��F���44�ۃ:��<w�jX]�'oz�H9f���޼�n�@���עY,��lʐ�:�է�F0Ik�4�U稣�3���$q�t��{s_j��{7����;F��zw�N��f�����&+��ө�P�R }J����Ai���=j�+��T��W���Ac�+2E���~7����e�6�?p�lp��T3m=�9��GY�B���l�^Фj�.��8/�.)�W�N��CM���=�rj�5'z����>�-��˝�z��{b@�O��ts��Fj�a+Q�t�^��F��v����r����e6pd�Pgs{xI�;���xRyBxZ�6�]�8��;!	��%
��x�\u�m�5|2�߼�������^z��2�[���hd�V��[\;��;I���\��o섬&�=[QG3q��S�luLO��(h(1^K[�k
W�#˅��7���(m���9#��<u��{�����U �9//<|r�d
}�1Hov�N�����;�J=4�,LƐݡH^^-*ٙK��TL�v�T���7��5�q�wZ뫻8J�)]Xsdξ�W��TL�*]�f�rʪ��<9*�o�<�(������"!�v'�O�ӊ�g���;&��lEL6#f
�v��>Gz�nՖQ#��;{ְ��rb�Jf��N=����g#[�Þ�kN�u���R���;��綬��ѕW�4��ϑ���E��=� T5�P^��G��n���_<2ڷKrpz&[9�Ī�`��nq�*�A4�s�������%o�D�=m-�V߶�橅ܾ��n�s�Q���d�^e�i��G_���j�-A^LMg�I��ޔ8N�cj��+�±e}��jL�\��f:A�N����.�v����
0�{�w4� ���L;�{6���v�H�`GN(18fu�^N��NE��l�`�e+)�6⻫���rs�R��Z�ԯ�j�������V�s�8�����YYŴ��Ow�)}�־ν�[�^LX���-tm崒 'z���zWd
�^�k��9=��i=�E-�%X�a���d�qov�n��[�V���y#T@��W��D�gLb�B$,H�n��?�Gx&�-_=T�k&��Tzּ����7�~k�z������
I��RfRL�
��c1�LdXE�� ���R(
@*g��P�
Aa@Y*, PPR��%b�d�@X�`��$�`�@PQVM0*��

@QH�`�QAb��(
*�
*�XAEP��X)��j�D"�*V��LϿo0t{��|����m������i�َ���r-  ��DD{Q	�w��];v�YZ�H;��U�.�rk�U�:1:�d��9�� 0���CU86Hx������J�4A:K#M,��Q��A��̷��G��{��Ǣ�L�.4HهOlh��剣5�=����Z�]�)�U�U(��NS�A����:��^�$✡�N�lZ�z*7�m�ۦ�ے̻����赲��Z���y�%%��ڿ�{m��+��$m۝MJw��.��0h���[K�%˼��(~���7@�nP���YG�m�p*��6�р��DG��  ����$͘�c�}��xR.'�R�[�U���ߴ���R}՗�|~���Tぞ-L�</"��hU�z�W�Nֈ3�3r�I�ü���)��r�9�����G;JO�5��s��c�c-.�E���s����)P����xA��N��SX�
K!*B��C��H�5"��[�)��ly��u�C��{�� ���ʆl�^�c��Y�����׼sa�ܙ�\��^4M/آz�v��{y�b!!�z���w���͜Bb��f#ܘ3& ��DP�.u"0������"y#�e������Dt%z�Dp^���A�C��S�s�zN��{n����g.��-36'��SD�`o4v���ʩ�Ki�$V�w�Իa�˽;��Cc�㎜���m9������b�aI2�NZy����GTp9Y6��
ץ��zsڹ���X�/r��J�J���D�bD�A�$���N���9X�O9׽�D�9#���A�f��f��B�{�gL*v�_MC/\�w�`��v��]����P�����=�S>��įVG�6��3�_{���b?J~�ͫ�g|�i�J��hc��S��H9�9��ꯀ�i�����ظx�,�o��`�k5��Q˃����E��a�$XӞz��������%&�4s�*�}F���j����c�"Y2Mێk?U|�9�B�+������u˭��L�LJ�q �w6��a ���U�k"NF䍩�t�1�L���J�N�Q�GF�����Zm�E�50�9�k�v�i|�J�Y�wHh{���A�[���FR<�fr���C4$gjp0��=bKΙ�ߗ,Iy	�O�����9�A�U�ޗ���|�f�Ԧ�Ha���֡s-�*9��������?3�<f{[�ڋF[m+:��Q�'!sΚ���F�X
S�b�5
�P��bp��0��k,������Rʌs̚�}�'�E���.ݳ\�%6�QMo��%ט����N�D5"�����w�tN=�#��_�=s�<�gxTX�Q��W�|�Na�cYm�#��zx���.;���r��m��U�n;*nB��u܊}�1%J�9J�]{,��k���k�ϢˋD8�e	��R�M}DkL����\G��h��ͧ�٭s�et����)/��G�kID��VJ����5Zv�7��秆�S���T�k�0"޺+@^h���~���~��1U׾�|��7(X��A��Y�="3/�9h�\.�����̈́��5m�������BDU�)�d]U�N2
Y�B�z��a�d%��6�z�P��-���O�2�k���7
��?zc8�����l������fe3������[�7,r'^���»x�W�+���V��K^���.Fcu7,�ۘz��ev=x!�M2�k\9a�@�vF��f��I΃�YI��_W�A9{6y��8=�dy�NF�^s�Cu��Oܱf�I!����W�|�1�|�q�F��>�Xy�ɷ�9=D烉�*{+��ƓWĺ羝�p�f�H5"{k[j7���#1t�~�k��$(�*Ho�:l>a�x�w+o;s��߶q�͚���D,$���I�������)���o��>Ci}��G����V�����)���zxj��H���~�,�A���ٳ/��ӡ'��Dq��h:Vl���!���⍍Br�택y[�cN�+-D�/6�J��o��z OnJ�3�՝-/��4��؈�|2ѧҠ������m�}��z�-�8�d�����W/v!�ȕ)���	��;ZϐZ�cˋ�ž�x4s�y{<�{��b�����F=Q�U!Dx�H���{�v����^0��((��^6�u]ZC����Dvt��ۍx�qqF��?(I������Y��~o�1q�^o��U��m��q|s O�-��Q��.I��:H���ר�G����dm[,y
k���g}��m�uz���Ù5�N!\\�~����ڼ�f��݀�2WX���s�����RBE��k�U�K���+���\�C��1贍0�b�?H͏�z�\o0�����{�χ���q�9}�$�i"֑{Zi��Z{��-Қ/�6g!̢�.{�+�
�j�N�d6Ͷ�J�]�ie�Ķ�L�Y�0�T�(��+�tq�q۟���@�� �e��'(L}�:WS�F���I�����fq�$BXËL6E�ʆ�|��qP#W��)\nn�׍�F��/���=�t��gM��x�.=w���g"[�������IBc�PMD�]C�2T��kd� s  ���!ׅ0��|�D&��w��ٛ4_!ǙL��(z��CJ����.�͎���O�K�y�_k�}O�Hr�G�,@���D#�*g���o9 ,'/ƺp�l@�U��dLHՑdi)a���&Rc����3DN+ME��	s70�F���@�,rҘ{+�x���Hش�L��<e[ǘ���ൻcz�C���­b����Xi��^��2�^�=�Lz,D�o�(U3�i��BKhT��E�ܤ]���J-)35�c����� ��n����zP����!�u]�㦻�߱����$H��-���-t�W�,`���]C�`A�2�/���*�.a����P-]���K[b���w\�=�R�Mw�%��s�_�?g]�'�9�#O��=M�b�����re��`-�]W�s�C	<I�l����+c\�{V]��da�-#�<���I��g�nlw���d"b���uF��HaXC�"$L��V7����v���%�(��,�憝#H�x�%ɝ]��[�3��;�3���Ϸg�?.=HC��"&����t��ʧ�ܩ̡�N�(p�%'O'R"�۶Y;]����-v��ڮ��i#Y�ײ�q'��:�V0`u��a�|�z.�J����~��9�=U1��r���ڤ�N��CA��/�Qz��R|��K�{E�ܣA�/�qj���Vf��z�+˳�!�S�����|f�Q�0//���w�нQy��ރ�C݈�xe�{v���;;�KhUuוh딝N���pp�Ty"̧{�˳f�j�N#3�kGq�:.�s�W�����UGy2l������2��Z�6Ko(�N��ޓ��~Xb�3��}3��y�/st�/�{Ƅ)U�]�2&��V݅��R�x���2����/i�gY��Zdv�G��Y3{k�k�8�T�pS��N����J?h���ܺ��ٵ�7<�ޜܹ��2WT*�ҹ�cł�m�=|��P}�9[ag.��օ+�z/�R�	Yj]��]���Z1ҚF����C�P������q%ZTx��O�8���`-N�D�O%-0���޼ut��S��X�a]�A��|er�j�H�Ggՠ�ҦU�8����[���kx��W�R��n��{h	�k�p�|"m�s��x�Q��c2���/f�GT�[���s$b�'x���Æ�@]��pO���4U��xi��:E����"|#��wj��\Q�gK��g,9�\}��
��/v�U�CX�0J�Ø����8�u��S����$o,g0'j=�1Ω��ܦ�K{�{ֺ��{����EPM�P��d�+"ł�@�A`E�,:k��Yd^���`$��1�L
��4��1����`�c[�H��J�@m3(c�H�AIR�RC��M$�M%M$�8��V�I*�T�aU�H��,\I��.j�(�-��EX�������>�g�d�ٷy����W>ˇ�k����=�4��m��#����#�E'�ml��ܨͨ�V���]7C�XF���Y���a��\���C�~b�/Q`D������~��8r>_1�O�H:��G�u�5h{�]l�U�l�0�)����4���:���;+�e�zN�oU��r'O�(ǒ��2��a!~����J�ݾ�F��YP����r��z)�.ٺ���v�Y&>8~�,"�󆽌u/������5I�Qg��p�\h��r�2�èyf�J���Aj�"��C�'V�hF�'���צ���Iү@�s�Ɓ�|�"
rĠۻ�9n�=�}���h3قmN(:Y�Ћ�wvf��E�m'��:�t۰�:͝m��k�I]Bo#�7�s�u����x���>�����tu�q��0H�IBH�*���8�?7�g+�גہt�����=�"qC�^����"���I�0�C�9"!����k��d��'#�X�J͝>>"�.>(���J��lw��!����U�Da�+l"!�G�]�<��Z��V�ޝ�4�<a�������D;P�4�
��<�*z{z^��Qq��b"x��X��HU]ZF�E;:z�4�%�b��B޷5:j�����4��{�����rG5|�8Qd=^?^"_���"��޺��6=Jr$CgKHCDe!��5�,\a�����}m.��ٸpR6l���v򵮠���̩ȅ��>��H���SN����S���T��:���(��\�J��;���I�6���'�'U�c�.T�wok�૆�wI�S\��x� �⤇E��Q��!��Y{�>�!�w����4��}vV!Fm}+������I�Ob�քq�!��u�r��H!��;ՑOz��{��TcKHj�u.�0��MLg�D������ɷ$�#A{������ʆ�|��il��I�'���A���9��8�v���I/�Z^F=xz&��$�KŔ~�y�h�}�����0Jhx�a�.�X�$�'�1zAHeOTݺՒ��;���ekz_�����oN���!dx�Dq� �!`"� ����c��X�Gsi��u��z+���6��F���J�I����0T�d������s����Yǻ~%��nCEZMd6���r�L}��e��������)��P0�x�	!���������#z�вǔ5�ʼ��'H5�B4�"��������(�C̬5���C[!�TC�>W��	�V6�+�\Sr&��*�r�b�ѮC�ZӇ�V�OX�V�Cŝ!������zؠ׎�,�nͪ��.g�~l�@.���6�/Pf����escơJ(����g3#	�������P�Q�gE@[;�k��ў�UGj�H��yP�<}�����_W�˥�}/ҋ>Z0�Q�HcZ|D!|��0�S�3RmK�����"!�O��<Iq���w��?/�fm6p,{ڐ˰ ���G��mZ�͸�۷EڸF�r�hy��r���]�	�P7��8�6���eӺ���_����ގ�O�S:�Fbf7h�E�~����⮔ǯ0��8evo�6#>���w�����6F�0�a<�"D�����{�>0��2���#
(�8F��^$W=�J��|�$i��a�F�r��}l�<{����uvz�y�G��h:B�Ӷ���U���Nɹ�=�,Q䴽B�"6�ǥ�J|F
��/����W�g�f#I���3xBsR����@����>���&Ԟ��f�����9O�(�8C嶩k��=Ϻޕ��3��<x�.2/�"`��
1����2/�y\�]��{��l
�t�8٣q#�����V�����M2�#��Гf�#c�Av,��L�g��uv����)����X�7���g5:��ordϟK:fE��n��d��1��t�vƚ�ş���󆽌s���t�Rw{~��"y�٣I~p�K�: Y�+8v_�sҙ��;ʱ���$(N�30��2��o7ׅ�gC\�6F�t�
S���	[$5���=ԏ��9=:P���e[�����(PK�t�$��3ń9��ɴ�ߦ�W�6�3��z��%���_5i���q]vOu�>#Ʊ:~/�L���1��圫�6��t׫���0�$�!�����t��kO�������bk'Iݬ�!�_q&�",����#<.]E�9Lw#�Uk�N嫸�D�/T?f��=���h`��?'�q|�#O_o������Ǻ|�lv
����mY�-~`���~s��=&��V����n֪�7�Њ�ɸ�t�;�7Wy���i�~���\\D�!���^$��S��}[�x�=����D>�58�:37^��^�͂�f�=�>KM�|�>8Q�B���D��~Ҟ��f!��e]KVOa̯^�v�6�dm[|C��{����f�v�"���^#��vUa�~c��3������<E�,�R��%DH�G��ٟc�#��$s9S"��F�0����$����D"��wF�{ӽ��d�(h�o����s���A螩���a�H������[�W!x�y0��k�{�V�k�D��,��A��O�]3����)߀�C1t�@�3z��(x,�����+�z�8��|y��g̡�����\�zչ��Kn�M�n��#����2e�'?W[O�L_��P�H���#i�Β]��B���i��,P��sR�����(v>$�'"oef���g���/|М���T"Յ�)��=�$�r�uVN�#I�Ȅa��ӧq�`!���>���g"�&��Wʐ3�a���4�!j�	����?���7������~.��?*���'H;}@i1T���]^o��ρb.��|\V<�~bjDX�D?F7 oٗ����TB��}���d�x<OP�υ?G�O���Y�^!�|ؾF�}���C��t�#����쳺��BjF��[��B"��b�Sq����#�V��v�т�ʈyMs�Уo���>5D���ߢ�8Uu��jXڸb|��^ͺ'��vn�p�� �ra2'�8��wC��Cՙ���!�Gx,<�`O7yO�����ď���a�Bk9Ys���ƈ�[��q̛�q�i#�C��"C�0f*륪���pӰ�le2.=����
�$5�6I�_{��9f�{zo}��E�{VE��B�H1�I���ޕ����#	"�)�`�/���,�A"��"Z���*w��'��-:G��G�p����4�i�:�)�Ξ���$����(�N/���g���؄==e�X}�^{>�r%<|zS�B��~.�>^���g���N�OQj��,/�V�@�--���C �㮔&D��Wk�Ro��m�c��e�o�Oq�'�;�������2�ȷ���	*>q��
���=�K� ����0��i������a��x��t�'�I[^��l����<�8�k�Uj���Uh�}�w��8�HC�����؉؀&dQ@��u��z�%xz�Sa�^N��$Y�q�#�}mz{�y�ۚj�fa'��<x��tƪ3�����-���^�ٙ�MGr�E..��q�o���u���ٳ��uƢ��~6� ƨN�3)��$�ܲU����Tn�K��ת�$H_E�RCy�PiQ���L��R���A�:hd���I��aW��[gIDʪ����)NѸY~k�*T�o�2�:#�q��W����ϻ��?\��NPG5��a,���)���nL)�Kz��X�ꄉ�8ېT&��x����U�A���-ܧ�P�9|����cY;D۴��ֻB��*мz�\�0hэ��
�ͱ/�6���/�1�̳����o�hnE�+�A��(M�{|��~�b�S�3��}���[�S���o:Z�T�ѱ2��J�GE9D�8�_Xq	����&c���&Dć_Z۲�i���;�B$�^�{(֧�o��	�W������]J�y�1n'm̾�4�8��8cJ9&YJ;V9��]AYݗ�{3u��UVy���;��K	�xLP���M�Y��u�����^�WrY�/kmd��o�	���0
7|j)5M�o�����i`��~k+8_��w�5���tzb�k�<z�[{J#�L�V�_@�l#t���J5B9e<3V�����)�B�6���I�e�t5,�t��gb�Gx�V;Z��f�ˇ�X�>�r��ؚ�m����z)�R6�T��s�g�v{�e���X�������N��	��OC(2�i��\ɚlgI���Mt��+5�'y�����J?M�Z��v�	���:�<�1mG όb�YO/8��Ú6��H8�<z@�7�!Y6e��i�W����&G]T�7�q��ꚞ[��>����w��<KG���ULKju��b�޼qE7�M�5gY$��'"R5)9k���i���.�
B�X�6d��:pҹ�����<����y�ʽ�X-w�m��
)�����AaX[��*�����bJ0*T��2Q` i�̤��"�T���+D���I%I1��jTX,����2(�R!�TF�c
�#���X(���X���"��T)h(�������Kh[(VT[����,�U�[aYP�F�8������QeAJ�b�����P���l��]�2.k:�Hz���4���᳅�mH���*�E&�X�~���!>#n��k�VRp�?x�*�˨��͝���D��}��xУf��f�r�z�2Lzt��f���V��	�����|���֯�M�Y��Hp�H�ƨ~�_P:z!�A*���{޹3��x�ҢEv�f7ˌ$����6)˙�X��<������	�Q�v���	?24�y��f]Mͮx,��Q���:�Tp"#��~����hO����*~��lC?C~[�^(]6<l��c��~j�'�z�{���p� �e.#��vUs�e1��!�.�v��3ܘ���x�����
O���z}�\����>�)�>{�4o���GC�.��ۊ\����R��ܽzmΧ��C�ɶ��me61TwS�����8-ؘ2�~��	�Ͳ�ƺr{vk��6�#D�vŢ��E�g��̽��V�����㵮r�!W�g\�]J�w=��#��X��Kp�+��ؼGP��+�ֶ�J�44��GYB�P	��
kqq��!�ʆR�^��+��}�>_i����!h/����tb�W�>�w3|���9�
L�*0��I^�ƒ�	�z?A�^��w�#L�����uy��q~b���%Y==��G���!�l�C�V�Tf�W*����gNY�W���U��^ɉn���͘�6*
�r�`S��;hYc��^a�U�W����o�ޭ��������9ּ������?����f�b�\�0|� WN��lXWZ�=z�r�L�ۇR��B�)���Lޝ��Rl�D�>?B0��9������$��t��b�V�]�o�	�v�����(��#ܴ�[����������#~�k�+��a��Oɬ�u��td��CJ�ݱ��׎e��[�瀃hC�kzm�����t^V�h�hTZM,>�?�sk�x���"����ݿ�,!�se�����r�8�ç���jn.�Y�9��4KH�!���c���!�,�vB`Iz�t�j-�J0��ᄑ�͖�A��h�ݾ�H�?���1�4�P�	-D�6��+=�~^���<9QI�=���K����P!W{�V���p�$+$AAy\�L\j3���;�#���֭��C{�V�g���E����c{&DWA�n�Ǹ�y���)�Ʉ��Ȅ[�_���w2&�)ʑ3
�h�e�5��f��r��G����i	���:F�E��}l�yq�A�g���9��O�RûN� ��c9x�|��;(����CI��I�CP�H��zi��>"��T�{�:��G���a�1�$�H�[��?[}�]�;I�C�x�.!��8�����Z�>�b���}�V��q�}n�W?��K� 	�%|M=>�׳�=C�q�H\Ǥe6D��H�Q	���+��y��������1K�KI<E=��Oz}ʺ`˴���r�ECu��9�e�G�C>���à�H;5��Þm߳��>z&�}���>��q�$ڸՋ:1:��x;=��>�i	
=܆�-���0]Z.N�؋-�� ���=4��W�Q
�C�Z�����X�u���<����M=2�W�T��dO��hk^�"���ԓ�������jG
�xj�V��5��W�qF~����]zOwQI�H�����9nFߚ늕$����\�/'Vp�Da�CK�5���_y
¡~�~�c&��{a�{懋������1�I��#'g$K����`_ �0T���L�����&�"0�@x���6o��V\^/I�A��O�8x56ZO��M]DtҪ�n⶜��JX��e~�]���mU�o�;>	U�����P?{(�!�	?���;;�c]�7yĕ��p>���*���Qg�[v�a���:$5�rޫ�5s�c��@�ɹS��N����U�7sa>�b?�KL���~p�E��C�d��{�U�w���(�;�r$xم�>�6��2B1l��s��Mgǋ#ڂ;I�<XZ�AJ���k����a8sJ�{�/4j��@?$����k�����c�,�Z�<��~�ǎ��b��8S��׽�bA��;d������V��؀��3�˓�
<�@r��8��W1ǌ��W0�.�����<вOQB,儈KX�qq�=���v��ş��\TA��֋�BA���kw���zB7ٹ��b�^=�,E�\YG��I������zyfk�줆����V���L$b�[v���g�N�:b��(��\�B�o��0c"���(8c��8@E/�\p_D�Ơ�}<�>h\BrDf�D"��^�S^ev�V�ʅsp�Y�N��lG�3P�a�1��R���۬!��|���zn/� |ǫ�x������R�vz�x$B��T�s����Q�ʼ���X��Yuz7���}� �yC��d@t�\B�����U�OvY�lCK�q�B4��=���땛��S�z>��)	~�=�x�����ղ��S�ha'�(��ի쾣��nغ���&�D)�5Y��z�gF�yF@{��4&r�J�W
rC����?Q�����	�#H��?���Uhqc��7�b����e���9`^0�4�hs�v��@���߽�?�v�'=&�ڥH���D�@��V�
���^g?
��yNL�T��u�ƴ"m�y���:���y^*����Z'Xa$o�7^4��z�3���۬Hm���A$Y�:�ҩ��C�_5�i$y�p�W����w7���͛Iq ��qQ�Z�����t�|D�LY������J����ܘ�㕓�|| ΅���-W���g��Ńp�^U͞��!��/������l��c*? �E�w��3��wѱ��iI����H��io�Cfߪ�m���"<%�x�hi��MF&A��cŤMݕbz�VI����R��=���x����4�-�pW#� ��b��ԇ�T��Q?�O!���������w4Ay�L�mi���K�up2���|��Uꓲ�j:U�)I	n�В�=�]���T�{�Q*6T����ߪ��>�MI�o|+�9z��/���6���͚7��{׋y�͖Ȟ_P��b�t��k�T��r����&�pbWK�냕橋$�*,�CϜ.����w����,r���^=0�j�Hi�8��^��4�Ә�TI��������C�Zׄ�C��	�_o��䅿�g��_/�l ׎����4��=2M�g���,�I�H����LQ�P������&Qu)�-����s�|uC�����I���q�gM����Ԏ5�phrDCǎ��I�>�7ō��.����	���z{�	�5���mP�r�����S��ܝ���o)b�	����F^�̄����QOZ�;FGٔ�n�11Q��Gm^�E}�DNXKw=?8yq�ɝ"r�!%^4FBHc�ڭ���s�Y�Fbx��$*"D/T?f��'}��OnM���XM:@q���a���~��0�ma]�}79�����z��)|���Q���p����L���x��M{K��u�uNN;�E�(� 6���:�I����|hs��5P����e�[�����q��
k�C����i0"'U�|��(��e�J��F8�XwJj���/˶r63�ߺ��c�v]G�ĵ�r����ӧJ��G�=,�nֆ�N	���T�=b�s�Z��N�ȳ��lO��<Õ{�bS짐���Ą3;���m��y��+:}x��\�ty���f[f�"���U����ki֙j�Z:�\9��/�l��L^!��kq*!�kw�s�oH$���ժ�*;0r�)�ww���m����a��$]�*��1��BX���B�Y�n�1��NCUf!�_h��� &�wÛmx�:�zbSv��цL�hN�>���w��תڼ�4�R�e�$/�A�����n�ދS�V����+�q5�>q��%�,^X��)�˙������mn旙]�;Ua�L7b������8[�j�Q�:�M�L]�2���UN����R�P���Qw|DQ֎���ýJܮEDi��U{�1�J�f@�V����ۉc�Tw�:ȸ*��]�Eg���<: ;��F�?��x'�O���>>����K��� 15�5>��Ў�OlA��@�D*����]ͥ�Ҋy<���[���W�R5A�^�n��u
8�����V[��_U���n�EkddyC]��Ā앑��R����Y4;��My�G���l>Mnf�\��s�9|�{	�e����dgZ�8x�r �w6�h�|v��3�����
�#0����sXA#�6�����I�TYՐ�s{
b�vA���`�7͵E�F�WV`�>L=k)���Io�X��y)5�
���U�`�=GJ%���U�^����JVy ����(b�dG��n�W��]齔ԘX�.��8V��xM�י���i�u���]��P��,Z�e-�P��Ղ��Ej)lh�[kl��m+
�$�ި�M	1�Z�@�̥a�V0*��PP�ՅC��TTX��,EA2�[��B#[�E�,1�E�hbQK��1V(Y�ˢ��X���E���cG2�+��m�p��Ƶ�1+���b`�*�e�������.\K��Ǧ���H��� ��`#1ræ�J�m*V�j+i*Q���.&V�,T���kG:���yN�����K��o=�;�R�;����BBA�͒w���jd�C��H#����R��J���o���6N�K�.6Xh!h�J(Y��"Zǎ��.�Y����6c�������7�#I���*�靪�gp�"�7�{��qe�B�$��8+�U*�!h�,��*h/�����cT!�_U��������m��\CTG�m��~Pŝ�Y/�Ɨ�<c�3�p������R�b/�����x������ےf`C�	����릅���ʼ�_0N1�_�{d�{���'��F��<��|�~b��=2wy�<"��3�q~CO�t�����s�^��#���*�*O��疃B[=S�-D�Լus�X�;m\i�o����k̂�J�U��W�K����_V�Oٗ�H�ЈC([����@^'�"�d��x\�4�͗�q>9~Yt$�.�5�MH�Ի��w)���6G5^T��
��:NS�9}����n�i������C�}C��-!�>��!喇)�ɯ�;���<}��1}Z��MG�M�������drI�	b��j�R 0Qh�6��[b�]��y 6�H�����YD	bC��.w����kH�I����1(��^�=��3�B<,!�y_�!�̘]/3x�`�f�f�RHm����D>#��^^-!���f"�w��<�ߘ9'�J߾��\�6�I;}�[c٪k8�d��v�7���v�d$�P���Z��n�Z!ޱYX!�)�V�l���(�Ne�?��g*M���C������lΧt�Z�ʃ���yk�s64���u,:EZ$ig�b���
�W��*�v�C̘A�cK��=F&A��<~]��]ۈpo�~��*pm���%FzTúQ*%����{���"ˋ�1�b����xs7�s����Ɖ$�-��đ}�Hi �d\����x��L�Na��yx�Pg��O�89q�ҍ�Zܼ��E܂��И�R��1d��vh�=|ႏ��˜�އXx���+���<V~j�W������d��ަ\I��6{;�b�C��z��3�؅��~ңY KB��N	�w��$Waq Go��|K�Z_�N�4�K����[u�W�x#Y �ʭ
�(�4�t��i�ٚ�8��s�}�cnO;��b����Κq�Ԃ>8w'Pb�v5k$��Lϔ��3.fc{��љ5+���y���9r�l��OK����g>#O�ܬ�>!���I�}�9�!�ÖySC�0�3'�}�X�
� |���wy��M��0yq�G5	ʈ1x�a
�����o�x�sQ�.׏���ݧwt�[��ϭ�����IZ8/���:@x�H��
�:kˋ�����滜�3�j-��V;>�V�'�}�o����y՝�v�̓���/hP兄���?��åC�kO���xu2m�#��3�b��;�(]6<���ǵk���uUqha��"����S��<N��x�Vu/ؑF_6k�!��ŗ��@�Kv35���2�)�.�����q�����6��g�"�kX�Q�Eb�#H����x�VSC�WW]]��c�Q�B�ְ�q΢3�����	Ș�-��i��52+�|kWF��<��}ы��Ο5k�ӋCZ=�hʘ����z�L��f1�0��C�ovL��qxu-<t��q���R���Z���z�=)�5��MhY'( "�A������8�r�+�?i۫jG��P_z?yO"�u�l̡z2YyBb�/o/��D���/�W��왱�>H_ J#�㼣A_1<���#bk3s�ny�ե<u-0�:#i�c�〢��:ϟC�z�3�J򢇳��=9�.,�M���ގ�$0�i�Z�Ӗyl�7����}�D�k�]|MU���  Y�l���t�`C�)����~���>���_QY��w��}���a#���fF���N�z�r�.��tJ�y�wM@� ��x�����:�z`4&_�'�[�����ZV�A|��0�*�H����G��:�>�����Gbf�>�v}�*Ƹ����=�9�--�I��x�9�u��:z��&�]�/����
�Z]vk�x��b��:� �L�oOV������z0��=Ai������T��:!`�	��|���=���㖇����-[E���
8z�1�=d����gOH|D!5ګ}�歸�dR��H�/�b�޿���2��J�k���6�xwrBr"�C�L!D�v�L���K.U�HV�#*8WH�TƳ+�r`�Z��}_UU�OƗ��ԀȻ����!���+T��+¡�߳�e���(H:}q��8Ҍz��|�	`G��]�>{{�YE�<r/ ���n�0�w.���N�Y�C���f�6����Hڸ�d�z�^n�?Q��_BJ8?`�-э�.��=q���A<0Ҝ��6���t�(�4�#���}~�ޱ���B+�K��aN�F�Cp���ݒ{���cK:|z�9hy�b�<�8��
���W�%y^!Z�����w-����b&�s �T�&z����lL
VUeT&,�w��#L����٭bcG���'(h_j4.F���&�8{�	W���?����o��vM�^ؑgd�Ig�]	�����bQ���$�_P�}��wg�:	�=_��dW./��Kť���!�M��2���ڈk�a�n��+�)OLȺɹ��+�й;��`c��9��dN/R�㏊��D�،f���.)؞ܸ��3$W��]-��1]ER���P��g&ff�
1�m�4�~^#��/�^0������*�S7�"��6ƂP�/.S"M�7k���N�؈lm�yNFyX��S�RG�;��.x�S~�%ٜ��Q��h�W���՜���"�'��,�w�=y7��ӧ�Z��$F\g�:D圇X�h� ��~�l!s|Y|��B�<x�HBH�5C�AÈ]��_w�~����=����K�f�z�z����` �C9V[ۖ���೬�1�o{��3�\d��G'��|;j�{�(�7��T���
��µ���ۣ���<�~k밳�!�J�Q��?!�P��8������J�'H�4�ΡX���������n&kE$��Z�����p:D�Lk����wJة���z���<���:��lq|�5	8x�t��PGimF<zM�=ۅ9���!d�T;�'���6&3��/r�)[��v
�s+g{�Q�G>��p�0���v��8yrvݧ�dg=��i\l�#euq7Z���+wL�:��܎�InjTv�u�!��B�i��2�m��u
�S�emG76g��C�^�R1��
"�:��@i��+�*�~��?xx�d>�%��>����Lt��sw+��Q����+�v�l������Ev�=���L+&
�GV��R�ޏDA��$�c�5�V���T,�z��Z�8sR7���H{g�¡G���d�4a��#[ˍ�g�Ċ�ۣ4VHL��̾�S�P�D˿��x�H��bW���#89U3/��OZ��K,���ޗ�qLTc�q�Q�3.����Ň��� � �l?'�~E���xٛ'��}~�]�����֑��>�ZXť��P��o���%��K���'H=~�?BN�~�B�=��jӶ�ƶ�{�Lo*hQɆ�;�6�f�2dM�4�$[�u5�_��i�#��G�B���x�>�ތ�^W�n�Ջ#�)��Κ��b�f��v�/t��_��w��٤i�����Uw%[��}Ľ#��)b����lP}���R��cAT��
+%�!�C�Qs����Ǧ��1M��s��L��(Ӱ�w#V��wh.�k�Tj=�"�]WxN
O�h�&N�VYwcpC�3�jBˤ��)������)�?��NM�l�g)�JlZ���� L;e*��O��*ތn
�s��OZ�t�pe����x��u2+.nWp-'�'b�]�S��*���?P�����+����,�1�c���f�:�`�Wy�1��el]�&����heݺR�W.}Q�4�ʺ�Cr�/b�y����ק�>��Iy`��q�
��5�w/�RMλ-�y�Z���IzR�����Uϒʧ�ȉK��C�p���R¾o�λA�Ӎ�7�����F����WwR�W	Җ��m9��I,:�oya�T��p�B�S��{հm.�]SM+C���)+�͐��<N����;��7�ۇ�N{Zsr����}�pᴴ�//���H�pt���6�Gf�f+�@i-IYiB�C���rd�r۳5Z���7y���Yv>�<R�W���N[h�x;��50�J�[���d��ʉ!���U&�z�M{ڍ-��u-�e蜰����X��C�>ǝ�5=�3��ٹڷ�'�)�]E��y���hJ�N��U�sC[WQ�Ü�n^p�rqI8�
�ⷩo#J\��.�Q�lp{:�W{T��1j�����IJ�uLE�����1�e�R�\��&e�C-�ˈ(�j�p�GaQ_(c��E�h�#�b,���*���Q�׶W�U:-UX[gIULe�2�U��V���Jb1C���ʊ�":��4�F�T��c�
�7M2��Lq�1��["�,��2�eTbc��D��u�4�VWH�c]dZ�LC]ZZ٘X�Vf�SHV2���t�6֤�
�5p��e�V�q�p�Z�VZ�Qbɖ�S-S":����I�7�a7s�˙����j�� �}����[���3�}z��N����9�b�򠵂@j�C|�.ޞ\_��������O�!���%�־�F�*�L#^S^���jH#R:��	iY:x�;(<#N
�0�Q���t�Y���������8a�!Y�劙�f8��Q�a"qsE�a~��g�Y����l�6���01[X�!��^�I/ou��KO���Xz��mF=_[��b�r��AS6l�1p"���9f�Ab2at�_��T>Wg5P���I�,��Q�0��f���'V�73��R�TXi%[�+��Y�Q�!辄�p��a��t����k�s޾�g�������'�dc�:hD,�!���ܮ�Y5ق�.���Ұs�az�k�t�\tkzp���F�No�@���-'����m~Hᎎ��L�Vɟ[�j.)?W�Q�E���^�*��\ED���VƟǈ�F&
��`�U�����1H:C����]n����
��X�>����W~�G�f�_��#ƅ����o�'G�9XsS'�Y���ȴ�׵ݕT��k�4�|�ѱ/,�zy�,�ƘG�#./��Kĝ6����{��W�������5<l1q�C�����\k����&yQ�ޖ��2���<x���د+����M�Jg�vsii���X����%���,=^��"޹�_'�5��O }�KH����.bd]܉ȵp��.�3���J��im��G�0�o�x�$�I��2P��OhLw���$�(W�V&Ņ��[���U�<�g̸�W��f��i�l3'I�g_mG�)po$3��q���,�e^����"���"J�⎛�g�LW��K��da��C�%a���;��mݾ��~'#�3a�gԉ�����z��K���:�oq�8*>�úu��Xz�|��-�cw[�U	mA��IiXax�m	���3O<���"Q�:�B���|��G,	;ݍ��N��Ƿd[S�Q��|��,ޕ��[A �[q-�}��9����)'[��+܍��E�����6f��6��E`~�#ٷ�9�5�D������P|:��H1�kW]��jƛ��Wd-dY���-1�)\�*.IÄ��mJ|2p���(���0�^���L�B�C� ����JK�1�]y��<����y��UzM�w�ʤ/�����r�UK�z���ve1�l
i�0Q�ł_�׻�����? cޚ�ti�%E���V��>v�ń�l��u���xd�5We�L��NSRZ��Ʌ���D��ϼ����a��L��fXv�X��s�F���<\	1;�"ne�~��H�"��N�s)�@�U��Gz�4�kmZ�Ϭ�8/�����57�J��x�7J�{o���h!�I,�|:��w��][����;�&��%ݨo�XM�W���]��#���H� ���#Jv��;&��	aW �Y[��+��# �&TwJ����q^u��Ú*"�=X6j���V+�x����1W�:2֓��JUN\��YtH)N���u�e�d�r�9�{�-���&���k��&��y|�*��,�.Ũ��SV7���bd~��-���x��ET,���Z8���]�5�/w�Aq�[��羊.S�0�~��yM#���0xpV�����qf�R&�7��d`�w��>u�}�����1B0�2�pv�Y�Q�����(d�z��X'�S"�����~�4`Zcjz��D�R��L.$���Y#C�Ԉ�t��O9�H�V��0�'���Z�є=�`��H�Gӽwy�J�&R.4N�j��2"�2�A��� jU�nj�ض�c�9�͉��h�i���o�jk�j5�p+�6O	Bח^J�;M���(֎7L)��"T���$�������9����,��w�Z��DY��\1��Ά=ٷ���4g9����7�
Uve��P��Wrv�Jж3��cf��^�����x�s���:9�gn���2���/�3(�RHrL|�jE[�׻��
.����δ1՞D����"�.[���9݊�4z��H��0{�-�"��D$֙�P���ȅ��iT��='yND��e�;]ahx��Q��j�m��W���j.��p���_}z.iZ���M���/,��D����"!�p6z�i}��c`\<3A�5�ߌmc�ko�T �k�t�^9�bDd&iI�{BP�a���􏠐Jqн��������߯|�&�=
�n=���^��aV"�z�R��h��=]�e��j��wLU|��@��6:☝,�W@�r�'/!AD[~��yh~�P�I?t�U=]Z�F+H"K]m��lɾ�<9����d�x)eo2r��mOx��W�j�V����f�1�.'SN*��B��E^�|FG)�ѻ\��)ݞ�P%f+�B[籖-=;���� �znj+�g�,@T������Z�ө3��(�e��;��(ߞT��7�Y�lLOI���-���a�mN��wۆz�%1�ڈ�>�*�@=B��~ŶU����ې�Lu-|)��"�Ӄ�%�:��}%�����/�Rr[�Cw���
I܏������.N<GELj)�ʓ��q&�_3;��j���������b%G0�*�=����-���֯xb�Q:)u0k��\�5T+�gc�y�^C�wqU�&��"���Y����-i��ڊ
�ԅeb��p�P��q���:u�y���!b���v��ː��e�$*��B��Nu�&��ò4qax��>�^>v^�,��*c�zk$,���c����N���*��M-�堎b���Q�Kv��t���5�u�RrÆ�	���SC@�U(�㥎;��N�S���:�{�G�/X�¼�H�劉�>=���}��{;A[(�K�-�����`�����=/�Y&^��w���ʺ]���~�������Kn����KEĝ0,�Fy�������<m�u%�j�Ba3��oF�I*V��_IO@jx_P�nɷsx��AKdA<O1i�1n�c�"�@WZm���n��@�#���3}�~�z�nj���W�C�����v'���ߡ������D��V��R����t"�4�\"�j�a9��\�h�z�4f��ؒ9::n�qR���G��2�W,S�q&[��QGm���L]W�@����Gwn��S2�9�Q��[�[T�-\�)��>Dp_���ֽ^�=p���,<�8|��[q���_�L4�����:�s�m�y7�ǳ�9�"���p����%]jx��f�ֿb�Ws#�Pi�ժ���+��-�т�$�*��=�(���Nk+6a�Uo�	�*��һhf���@:������A-'q]>"�5T������Ar���'�h%��j+�qԂ1�][��[-;�9��{VĠ\���f�h,��ɞUx�;�J]�߸b�):�F7�S�w �`'�
մL�&ea�UiHW����@9�\p=�}�)m���D��x�X_ckF��}�вl�t���\2��/g��WA26t��r)s3إz�H��i,[�t���\�I�g�e�cRb;�ӚA��_[�9��Y֮��n�8��dV��������$Q��{|��[���=��:��&\�g�l�8؜X�}��Q�vsg'w����GN"�!�d��vLCYo�e^P�ӣ�S�g����@m�(��Emi����A2�9��˵�v��-;=;ܮ=�UƱ�B "�]��afcyu�Z�:A%�+�]�I���}(��e', 6'&��t)�)��0P�窮%����ť��f�<�RXΌ����ˬAI���gV�E35�ʚ@\E��F�,kI[K�(��!��j��S3�eB��q�J�J�ȱ�mf4EƖ�\�3-dR��ҦeȘ�SNkqDƸ�)6�֎�H�R��*6ت:�֩S�̲k.j�֌Ш:����hfS�(��.�C%�\̙i��s� �X�+�LW`k-��E�ܗ�̦eYmu���1lDՂ��Qd2(�~E�dH'�՚%ߥuE� [�����熯&�i6}1x�~�ѓ3a19ڀEG�j�VxI�J)y��P::n��gPJ�"�Qȳ\k�,x����2��M�7hC$5�&N��p�Qv�[d��t	+���Uj7�����㍑i�%�>�<��Fp�/sQw���s@.T|�l�9$����r��W9�KQI%J;S�=Q��"�NCMI�[��)Cmw5���{m�=�x4�s�њ��f�e��p+|1j��;@t��
�O���e����︌�ov�Ḥ��������*�^iUQ"k�>�Gw�����セz.�'��WM���y�E
fb��Yqζ�mϿ)�R����<��Gp=a쉼�vƂ��96ɪ����:kn&����2�u�b�'�3 R�*lbu�3/�],��bYMfx�ul�@;���v*
��l�Rx�g���m�rq����ډ��<Ͷ��߁y1}�w��.��>�������:1�n�y��\O@�~�,�AZ��'�-C�G��n���s�F_���[y�jG[E+gP?�Ԧ;d9���-}�ϡ�uW]7�:�zNΰ�V� o��3b�R�v�{d�����Y7���M|p�m��f���J�1���a�����nU�T�Ф���
샵74�\��V�}�_6���)��;;3�S+%�m��h�[1Y�=f�4�o&�q|���%<��V���;�t��C����H���<7ǔ T��Z�Iw���``�J��w@�vD�*�]]�D�H�qnU�"�W�&'c{]��UL^E��2�8-�:��tu,��e�d����v/�߰���m��j�QH܆�aY����=�:�#0�<�ڀ��ͬn
�!W���v��3��Ewq� Ҵx��뺽aFI�|0X�i�ZB�Y��n0M�;�Ƣ��K�IJ�'��+Cg!F�oX����Vɩ�Óf2-:��'��VxELi�%��*��v�����T �T8��Zz�U>��Ys;x�e,�.ٮqة!qʣ�v�3�EX`��^��//�BU�͡�`�xspϜʺ貛�Z�f]+]Y���C]��";�9Ϩ���X"YB�;@p��j���}[�����#���#�E��h�C�zy�^g���Yh�����eG�hd�{ǽO�"d�+��3������ջt/5A[Ыԛ���|���#��
�^V蓽W�ɴ��E�e����x0C�md�#�D���eN4a�k���Ol̈� ��zje5IC�����-��˸����Z����P��[��'4YͿHw�1X�t�]V�&q�γ�,Z��k/g[�1�e�qr%�#]:�{�,�J�MН��ե.�y�SfmLV��Fq��E�/�Җ��%�^���\֙�R�y�Z�v���yf�s��_,�i�������{[�y��Q��V�^C�^&�UӚ�#�(;F1K}[�8��9��6uP����KQW�.��y[�Q9y�%$�%N	�O���"���6�%}��=x}L�C�9����Y�t�*��p�������y����[�N�K�[�j����.��u�~M�^��Eh��],�r�)����"!��F[�/�}����SԞ�Yq���d��&���# Y
�M��rqA͵LC�Ð]�R��U:D�Ey��>Y�h4�u�9Ξ�`28�ѱ�뻯���8K�V�p��p�1sQ������<�9�32ģ<���bp�ht�e��No�S����э��XVӆ��1멐�6:��2Fp��r�ⓓ�{j���HL��\c�
��b���JB�]c^��gy(�F(���ݾ�������p)�<�0B�-�� TN�Ӈ܎���+��<��5��Ph�uWaډ�\�s�ue�i�bk�1�2��س��y0J�~�`=RQ�o8E��v�b@�閜�v�q�{J={^=tx��j�������K���5�U�0=/��.��fL�Lq���6�Fq�W���5��Lۊ?>��{>���S�S��[�jq�Op�W�ɵ6��ם%i�N��fe��=���m�2ܮ���p��5M�Pbv'{]�ݬ1*��&�Mk���I@5=P���;O4�Q��3�f������0 �w
�j�!�p�?R΂��h��s�3+FJ�������!�5{w�Z��q��
a�����Ҫq�h��*�2m�ӄ�j�SX�˒[��yW�����$��^������͎�yZ���'u�=�1�Ö��^�	{1���!@J��%Q}����Q9U�
-2�]
u~�Y�=�X��*}��J���C��=�on��z:���!¥]e���,zF�8y�e� �"�k�e]{,�.�����{�Բ����O��8�-k���DvLhYZ}Eb�E���v�(�&��Y|'���(u�I���v���]���h���Qo��(�:@���p�Eŉ05�˟^rC["	��}o�7jE{�2�$�N�����6���!��&�
a]��.�X��8=4zDX���!\�n�U��`F���5�u�>q;�w���ھ�&��-���9�v������@��m����<������=����._�)���@��=���Y ��&!n`)�
��u؞5�I6��������>�s���L�/N�x��H��B}��
�yq؅E��u�n��w&���	��n:`�O)� �E|�.uΊ�PO�������r
ڮ<�e�6��=Ne>̾Vvޫ���z6��]	�9�A=w:A�W�i���na�ZЉ��i�50���-i]�x��� �Asyd1���*�h����b~����m
�p]{��G���ꪪ�Vkd��k��W�a� lt��څ���}���I�
&� V�������.�����D�a.a�Gn�*�xV-���fvީ�hE(�ru�gI۫���{�K2���l�_#����1:�Q��V�
�*B���h9�Q���G1a��tw�R�O�\�Ʒ��ݵ:b��TDM��V�z��3%{Syq:��%T�!�����`»�%#��������{V%�wY~�J��q)juHT�ܧ��ν���@���D��jڗY`�*J�y5PY����d;|5����x��9���	͝Mc���rd��.viӑ(q5���f�s,D�7y�s�s��������ݯ����	��b��c�ׇ];:n��_QdȂk��R9 ��NE�2D}�����y^�R��;/&����Hg[S�3����
�X���[�%�����(�
�C)�Pۺ�Dp�MZVp��f�-Ρg���/��l���G'����*U��������6J�v���I�[:�R8�V�`��%�%Eה8b�R~�+S�TA�ȐO\)��mg�.��Vp�{�U�/��%ƾ�q�&q*f���x�7�F3�����H�F��eõh��*�r�F]r�v�G�4�/\���ȑ4��Ox��J���5�C��+����΢z٥�Nc��$��#}m�ݶ����[S,U���	�U52����%�8Tk���v=*���xkNMI���S�I�n��Q���h@����F쓁�;}�mf�U�
��-%"~��!�c4�sPF��r�Q6��
e�"Mh�V+�V�1��+k�Ȧ]aQnQ��U5k�!]&5��e0[*�t�k1T,�YPR�Tm�J)�K2�4�H�G)����&X��5�
j���It��\(�[�,]:nJ�\�Җ�kl�$Z�+1��\�Z���N�N�)&�m�h�*��L�F���5���1�Kf\r�#w��}�8S�~�`����Ed+�		N*�ÙW��&pi ��15�ƃ�.�UX{�*9�ͷI�Ա�&�P�A���tU�� ����W�ھ����\=M�n
�ë�aO�z��nkC�Wn��թ�bU'�������h�^]�C5S��f���e�F��;�`l��!kU�xMEM�cae�Z�ع�^굓�Eqg3ٖ�a��z���Q̝*�A�y���3�EZ8��p<+��b左*{�`|��qJ�&vv��~�\��߳��~E9 u�� ���X�_Y����8����zL���^�s�ָ�،b��!��}M�Sl`�&q�"Q@\��h��J���f�Z<�M�BL��7��[d�A_SYtdb�{�V3�|7pB���\����ʅ7�Wڛ�9��Y����Y����0n����G�o�:y����4������:�kgZ��ǜ�D%�L.���'o���[Ncuv]��"c	�g��u��\b����c�6��=T����)X��r��V4yNG���C&���N�y���q.��Ӟ��<͌��� ������E����W�����V�dk�S�����;�s��`�F+%�)��\ʌXi`p᡼�*)�#y�C$2-�c����9���(��˵$_;��,�-��ȸ��r�k/�^*hr�ù2��a]�����?1,�I/��T%W�p���rc��:<�=ls�d�������YM�`���"3l�1��DvLht\�ݤ�&�K*9t�r��%�VK���\O>�6�c�?]��M���/5ȵ0é{|f�,7��t�W{08(���C�R�F�h�Q�����	܅���d���4.�U]����3�������\y�|3�o뻥��(�mu-NG(�����b�v����-�������EkN��d#�����]�{fd^b��-xC��f���-�N��Q�u��ӈ:T�F0Ȝ�g6�:������T�;�ϯ��,ݞ61ټ/g4��8ث�X·5��K:�Tb��Riog�mǂ)41lG��O��U����%	��u�*P��k��l�"zO���=O2�Y<�˚�7G9��U��`�LJ
������eM��6���U��f�/]:���(��%�m��%�����c��ͤ�=��ߺ�n���0nS�X|1�X����6�,���f���2F8��^�t��ˤ�UFi7���y�����E�3Xʛۊ��#�n�6v34sD;�\���Sx��c�5r|_z}���6W�/�-�.��[=�y�.trU�p�UwR����bg�!��d�F)��D���2;!�S9��X��l��pZ�Q\gS0�D��m�q���q֠'������Ё]u���_~knV����N�Y�C M�PO]�7�o�l�l�1�~�a��~$��������b�=��ި�	,I�IgO.�=��[z0{q�-�� ��Zi6�m�PL��v 
	��[�K�/l�}���7�|F�{��*�t�﬛�̈́�i�E��I^8f;�,�L5UΛ���5ث�R��y�dԄ���^���EAf��8��/���,%*�:�
7�TI�y����Z~��`��O�g�5M!Sm�M�N�af[�;ŗP�k�I���/��o�q+�l�����?����I���9��YhFU�o�j�W �2��p[:���f,���}�C��fW�r�n��^��ʽ�YCx�U>N����Ω�9]��-�U��eVpzgT�I�4�����m��f�;�N�����u�S�ij)&�ⓝX�5u�®ڷ��(F)h�;�P!���ԛ�T�]]�9'N�	zyqi�2�CF��5f�9(�˜P3�
3��"̧5M���nËE���xz�t�١��$�5�k��(8���5�b1Yϵ$|��[9\�l�!�$8�S���G��*�E�2�5����R�wHe_^G���9Z�$�DYc�\���ڽ�����2d�>3p������3Xk��|����;TE�^\��Ow' �`���DwS{�rѼ�7b����C5��{�XVl<d�Fd��]��tq�\���+�tu�mD��4��к�Q�r61�?G��u�����2�uz�#	0��&��)ŵ�ص�b������f�t����c���>��SQ��˟^�!<�]�riW���qA\Wyi��U�dE�����)���&�L��ڨ��뫔��jr��k���y5��\ަ:H��l=h�(3Xu;�K8@��x�ثt� �-aQ��V� ��5W$�;z�*��ԘM��Q�;
��j���V���D����7˾={��)�9�~j�
hV���#R~��,h��&�	�V���_)-ηSM�7�	S ��6QiI���Rn�(��)=����v�y�Z��-a��������0�����"㈖��iމ�AWP)��»���o����>��X�nZ�y:�ԇb�$�cѶI���{���.�taI^p���oZ�M�ЯiۛV�,۩|��r�7�CƄ�e���v��<bczk���Q���x��Q{�w��0�M����L�5c�L�A�Uq,�b�Lq%�=�/r���0(�G ��$+k�K"�) �:]��w�g.Vv����o]��u�K55r�ȭ[r�)��A*4:�g}f�[�gf(�LQb����[�=gkj�K�pz22���]j�B[r�U�=CU�	�<�iu	0�~�B�g�R\�
����ξ[�l^귓ё}����W�8���(��5������TӲt�O9̴*�_=�P�9��D��7hVNE��,�S>�U�=����[��<L��S0W��`�̷��C�G}|�g��.s�Z��k�"�j�������?K�O˥j,X*��B�B�L�9�EU|�D��WXVSф���IP�HR���	̪��ϸ6?oD�_	�m(0�	! Y	�TP"a�Җ!�K`a[�`�#)��3X0�'9���l5�1��Y,���S�톐����@�i@9FϬ���/�>kCxP0a�zA��
�xJ�� ��p<�2g=
Rw7žI���@p���`��55���A5|y���\����"���\U48"D$����"�̐�������bO�t��r?g�`�0X���QW��ퟭ�v0A k���B�,u��T�0h��chj�����K�I�kT��)u`-�y��� 0����;�]��2�(�*�bl�.��RhZ
G�� ���*�O�u�Ur�D@�WhHX3$���Lp*&��i�b�g�QWE��!��Y7�hn�ͅsa�|,�H!���\���=Л�����,��Yc���߼�a���Ӱa�[sXuCxy��s�O�NΈl�йP��`_t�HJ�{�	�r�_�hu��` ������ѿ�vz�p`m9� �������z��8����$]��$�eJ訢��QW�x�A �"Ǿ��H��\�h�gQq�1,�
hX�K�QEV�p6������E����F**���%l8��u����XԄ%�102�����Q[ݗ�@̉���S��ơ�TAU��;�'3��)�N(�*�P�3�_�+�����>����[����7����J�;�z�VF>GT#q�V��ut��'�F�)�J��春~４D^'Gu���p�$�"?�LR=H�*����B1h~�臠��`t�j�f�����j���4H=}$���!�Ѐ-����#8�E5'��#?�����i^���*���N]+ؘp��@�z�b�H6A��vk�N0�@fI�+��K	T	`�S�Zm�`EW��h��@<w���c���79u��PU{��;��P�.�}r7Y����[
w�U)b�h�	ؐ|���G^����"�(H�[ 