BZh91AY&SYha)5 ��_�ryg����߰����  `_�G�  ���g׫4"�	*�Z[3�  O�^]�C���>���ݺ1P7nl �-@�ȤT�� t%�UMeTR�����B������.�Ҁ��d4x�xl�0Q��0&�=ۡT��K��'B�	�	3��i�={�u�pe�z[�� !           ������ �F�      ��=B��� �& ` j~�D�� �4 ��   ��2f����CL4��!�@4 �4)�BA4hd�Od�MS4LM=�6�<(��J�2a  0�dɈ  7�!�p�"����X����~Pl*�T�Q
Q���П!u=g��Z�����6_�!������b��;�����`��H���	Cg�ĮBFہ'�0*��":"/a��Ȱ�N��)MB�I$����B�h��E;��w�����r��>	�_���ֽI����]vo��c^><|���X� c HT6[sz�ޏ4�@��M$$&x|��Qh�br��*�+�.��M"p��'G�s�Ԣ��Y�p�4��<Up~]mzp�h/r��"�E,�a�+ӯ�W���-�?)PmM��-��d�' �"�/XL"��!��д�Er�`-�-Vh��c�`J"ك�t�E�Qp���mK5:8�Q�2)F���*^�1E0�dR,���=�yu�ˍ��Z�A�+�Tk�
�{�{���´sG�SH�h�v=^�]��^�A�]�q\�����)�)�,�pB���,��Z۶��������SIõ�T;�8�M�m�Hd2��=+q���lolo�7sG0Ƀ�Ŋ]��d�WP�sN�=�i�`)��m��wq�1�x۲( B��x0(�Hz�y����c�&��� @�B���c��E��zR-����� ��,�s�#�	��(����(�W|���%�,k;�F/` BȢ�]˱q��"WS�5�6ƨJ�*Ԣ_G���A�S�u8��]��d�(�"�2,^�����f8�q�L��X0���EA<�NFv�lc�c�Ǒ8��������p�F�˅C=�z�5��:�i�|�$�򗺎��(�AD�.��ei!�Y��¹��3)����/�w��	b�h�tL��ٽ"�"q���)dY��,��Ű�~���"����8��N�9��,�"�j�ż�Nh⭃���ʃkg�r��=�A�Y�5f+Y�V+}o��,V-�J�7X�0k�[�js��"���a�4��3�h��c��6�Hd=C�u�qxT��PA������޷��/��+�m�6�lm��6��<u_Q8NE"'��s�@�''G�Q�SÊ��Z�Y�(��j�Zjr(�;n
��i�zy���{�����-K�q� hg=��K� �ᑜ�^��{�f�k7�x�Z�-��ħ�%�,|p��Pgk>�Ӊ��b[��<c��G_�~A!���>��ßͳu�7��5\����ɧ.K��l��D�U�I�+�s�/׬��ښ�&��oKYn����e�b�tfߥ�g�[�}VJ�~�Y�,qn*�Q36�:zo[u�9�g\�2�:T�{����m]���ݪ��2�W�C�)���.�����p�E��u�&]���D�����P�}t�Q�`�(�͇vL[���＃�?�`���g�n����V+3핦fe��U��C׹\]�|���,�x8�0�����Pooa�C�A�W��ه��������b����n�ݡ�Q�	;W�� ����푝�?����S�\�ɰz}�L��>����s��Ng�N�͹�V� Q5SNݸֳ���{v9m��e�fBs���2��S�o�%뫒�Ӎ��j:�fF�Q78G��s�������[���{�~��_������'�dC�qB�"���3�5��������Af˟f�Kߧ1?z��OK�w��Ǿ>�n��C٭kɳr�u��q;�y7��:��)M�V����o]��e �� ]���k�����}&���d����<'��[�}���ʯ�,���Szk�4��0�u����[��^습�D�MU�X��J	ʅ��d�jL2lY�%�ӍʯWD���;�ƏsV!���<y�<,�̏*U�=���`��ܳ�=w�v\gx/v,'6i��J�UoɌ���
#\EVIqrvI�+̏�/�k�޵�>i��eʰ���}�E�}�Rv�7��p�|P��f�˜�����͐W�F���iϾՍܔ��tl��Y�RN]ۣ"ڋw���fMNa+m�K�vْ\W�lϏ��"e۱�����y��.��yɟ������T��c���+�\6�5���N�｡����deY{_��I:��Z`窝�gqg�ώ�W�w����o����ͺd�ʻ�]l���M�5�{P�v�;L��<�|;H��6d����nVM�)�wf�^m
�g{R��&���5+T+<w[�����k�}3{sv-}�p�T�U;	���M�O�wf�����\&`�o�3v�uZ��e���d	��ls�f�f�x�u�{� ����s���Ϣ3�Z���*��f&�������]�;��ry����,��4O7q����N9I:9��0OU�b��}�:���Í#�H��a%h-��Й�qX����׳�'�f0/�%�	;n�����D�F�,����J��ɯ"�5�/��=m��UEX�H��iH*V�i���Z�hVU#��sf쒃)�je���nō@[�Γ��'���13$!a�ym&�H�� �,�LLj������|ﲬ�і����w���bJ-��h��hM����3��e��]*�%��v�&Y�f��d;Z�Ŗ-�V��n4(�r�8���!N�Q6@��V\��w����xa�py����f���Wז�-N�:�R�9��,	�
�GG]{031�{Wb��cو ��*��H�����-Ep�o�*�b�d�	���+#�ʿ�+l1��^x����=�����ΏH_��5�@�Vب���wt��iXЊ)��=�֒�>d}��ck��#O�y�jwS��%�T�+����벻3Y��]u����  �� �M�u�0t�=Tt�
d�	�ə�w�� v(h #RI.I�s�L8	q9��&��Ӝ�BZs�йhH�>$�s���L�d� �������QA �jBШ��h2 �$�q#�9�\p��$�f�rG"E�@�2!�}I�(�6�6���*�m��b������dJ�r�h�gY��1R�ԗ���ĕRJ�]bb�LL���ِhe����4���I	
����*؊��6��+��;�E��h3��@�`�*�X�MT���TƪLLԸz�j��g9� 6�� g��ƪb��Q#!$�e�s��;��%󀀡0!ȲD�������O�C��>�y�=G���=G�Q��G%�8x��bꊗTQRQuEi�Wh��Qbk���������qQuIq.%ψ3����bJ��v�~�"$r+���R��y�M����/S얝��[Y븰��0���z�;��mΨ�r��_f�`��kZr��Ur咑�ZNB8�"��󛛣�A�w*��4jE�(�a�R_|�<�s<�����0�H�]xK{�)�C ����Y�F��6iD��E$C�Uo1ϱ�1囙�\��6ߔ�ĝ�8k���f/<�����ļu�kZցPֵ�kZkZֵ�Pֵ�kZZֵ�iQ5�kZր ���C)�L���$�� �$������Fc�$���QeH����)(ϓ?7��n6�و�G�ZdZ4��*�r_3�Ú4Ơ#�Ƅ����6�w�Qȵ�Z���:Q���Lm�Q���W�w���)���΄"c����I ����oX!~+��� #ܫ%�r��������Cz1k�f���|���+��X*T��C��V��|��1-#J�L���}�9� ��H��a�u%8�i����Fub1�pj,�'�b|7Q�b�_qb8�B���Ф����7�o
�dQ�R9jl�P������u@a�%��EbI�� ��cm՝��iZ>FuZ�ʨ6�j/�u�m261�������//ŕ>e���io�$h#��C�h�����GO�>gO���*��E,���z��2�-:������F6�3Xѽ�>���g�gX�(����[86��)�����RQ(���|lQ�qV��˭���4ut`a��}��T�P�_��CSlb`'��>g6���C%ؚi n��s$kf��1����kB�J(ٰ��8�67[�b��˯^�8]��g35���14ڏEV��eq��HqȄ�j �@��h��f���N�F�%�]�!�3���)��N!�>E�xٰ�BÇ�HS�������D���o��]iiC|W犩(�J�ƹc��k�q�B����5ı���@�>�'�'����0�,x6Y�3�&a^4t�G���x������q�6M�ߛ�1S�0x|L�`�?'���t�ҡ�h~���DYM�
&H<�f��݈3���%~So��S�dܜ��yj��5v��� �ӭ�ES����u��������-a��s����x�s�fl��Y��x�^  �� ����
^ �
I R �hR�X3AGNԍ�\[ �W�rA���/h�M�K�;,$c��s��&&>�̕e�ώ�)�4-[)��%�Bѻ�4�Yd9�Hd�2u��Y���F/	�E,\�C!r�Ap���`j@��$�u~lHH�)�"K��5s4��&��%��ō$K�.E�9btB[qd�t��Y�p����\^DF��j!3D~=���U��#�l�S�V��p�c��szk��C9���a)���%��aIP� m� �v)���F�xb��[����BK,"�"e���(���!��(H�M��-X�}�v�Z�myv ��l�Z�t��
j�%*��@�F0���������̑�e�& ƚgB(�d�4����p�Xк�u��ܧEH67b�5Ӫ	e#��8Hp��
���9r�2�.l�cɀ�\��`��"� a"�0.�F�Î�䉴�g�����R9E_
D\L�
q�!�VDx[$�ؖ����������`�7d�l�d46��m�z���CC^PH��dQ���c���S�R��h����GM+A�� ��4O�qcAR�1h��!��(�����&�Al���4�Q�9>�?VF��5n�͜��袙��mK(�IK�����:�w$��4�Jv��L����-%��2GL���qr��z�	�[IW�@���u�OU�r�"�R6�F^_,4Q�>8����U���kZ�{l�7�,�Ū��8�� ��&�E+
4��}讣�N�%Tt�V a\P-.�6�Y��@��������^���[R������6������LrBƛ����ȏH.���Ұ�,�>���(����1��'!)9+�[f�yh|�O���>���%U:�U�9]��ʬ���<��((.D��P���������(j,�٭v-���x>L,�?�~v�t�0�x6a¡���*͐�	�ل0zL͓�	Ä��/<S:O�������	����l�htatك��To��d�D����1�7�ӛvm�E�(��nF�VdnD�гI��]�%f8'HG�{Y�r��V��ʍ��^��'f��x��f?G��e.�&�b=�uխL���a1ܒM��׻�q[��5�nݎtQ��1\h����{�3���U{�L�xl���)XG�M4�(%�ax�)�zJ���o�1���l��!�k9c��)B��Zf̕=�ֱ9#w��l5EUJ�H�D �&5��+j:I[r��X����쨹�v~���B@����) J@H�@� �%)R�J�Jծ�o�G��P�+b��NDݵ�Ei"RR���N����u/J��fփ���8��D�@�I�N�GO)��x��aϑ�[�M�>R�agA����l�7x�GӡԏT�yA�:Q���7&�HӃ��p��F���y���h�Ǝ#������FJ�5,�@�=d)�N��q���cV������3ƍ�����Ǧ��_�:+K�
�GU�&�[��$nk� lg����ͮ�[��\m�ˎI.��]6Svlɒ�`�A������/3��p��y�2v�U-V�&02i�Z^��;�s5���F���t����80�[^��gN�a���G{�.���e�p$NV�Vm�X�hd�['( �hj.�Ԭ5�F�����0���-j�"�45�I�=d�p��ݢf������ÍbM��(d�����I����(���h�
80�K�haO6\�8,�	sM�bP�P|sE�o�h�yF��X��K3F�$Ƀ��pE�e����<|B��Fm��W�ȏ-]�9&�h��͢�Ph�m��4��t�-@����f�p6t����F�mG��0�&�h2�ʆ���E2pQFCD2Sn�YLO��XZ�Exq�g��F����:�Lk�űh6n���L4��M���B�u{���Q��_ivL�*�Ά7R�1��9#�@v�l���`�M4�e*������#�����ƍ��ҡ�R8sp�8ⳛr6[���n�8�x��:�ӑ��n�=}r7�q R���/�M�����-D�R��}y�.��d��dP�#�p�G�kl�K�A�qu����QK��XV��T!�G%ka�Eў_saXo�[��R����|�A[�0tpr�D�Z�9˃YL�q�ݮ��ig�1�����OVǏ���:K1G�ff+�fU�!c�D�	���#7ɱ��¸x����<a<|L�C���t�6��0v<*6aD�f���k]��<�������/\��3��󰮞���1��C6v2��3Ѹ��n�
�n��mLѹ~���X�}teXՊ�A��o{�={�O����(#�
 ��
    �
�J�*M�CA��ܐJ��4�"E@�ʏ~3��0���tq�H7	T��Ț��p����k�e��!�U����i�YD8%�ی�Ti4v'Aƨ�V�,)|�-a"9��MZT:K�g��aKo��A��":l�9���h<|t��V��H�tx���!���w���ȡ֛��,b�*��<����ֶ���&����6�8p�����!������Zm����gGLyn�Ccr���P�Pw̓���k�I%U:��R8����h�ќ[<l���p4wG8ǲp�QA��RS���g��fځ����.����Z<��ߡ�Lp�N�ș
���:�0��:E�h��l4?��6��%M9�/l.��4�4a&L���P�3 UUFSkP�����⇖���rPSA˓&K)��8�gP0�م���|�2FM�4mbg��ϊZ���������up��it�]������4���c���lj�]�>���Ӈ�!���>�d�mdR���emd�Q���7f�6� �MT�����ˈv&�rwv�msH�1�*��/Ȉ��h��[�<%%��s.Z8)�t�/Э�ś��-3�4i��8QӇ������NlG�8����n�ΰ��q���	�j��SF��B�//[N4pV�M�	��X��U�<�L4_�FK`0C����Ln�.`��r��&��d�sA�!��')�X����E�wБH�'���:�]4S�AÄ�W9ne)9��d���8h����3Å��$��]M�z�ԨC�:CԼ�y[GQ��5��S�,l�-#�ZV�yx7�|cn\0}L��V�Z!����Z�8Y�֩���8>�Qҍ���	���)�`L��t�Y�!�e��%�'�c�׊&�ǲlz6M�&7�
X|x����~������i���xY(��<
��Q�(�x6di�8{�>��d��R�2�O��������r��ǿf����GT�����1�N��ɔ�u���6n\��,;M� +>;2m��_�ׄ����=~�k���B���,R_�������,<�C/e�X�~��cF�)�s��\�H���33�ܨ`=�|��n��z�Yc̵��8�t �1�������g#Jb�`����N�W&6R+'��w$� �h��U�"�_~��^}�,        �b���b�$%�tG�n7l�D9�!�ETM�p��L���V
�rYt:z�cf����5eR\�i!���s�7���BC+��ΉbȻ��f�ѿ�6������|b����GJ6ѿ?��5���|(wEp�Y\���nV��-y��	�Ť��n�g:ލ"Ț�3�w8�gAl�����1��\���4Qa�ц�����u#�][F�K�G��Q��ֆV�E�>�c�^XYh��Q�V��E�-ZQ{�y��4���͜0������L���؍|�Qu��V��-i]D,�A���9��j���]�T�N����l��Ӑ�Li�I��3�AsE�d47y8����VM5=��⌨C�v��:)�f�nM��y*m�E������D(�jJ�*EՋ`}�q�tMC�Dϖ^�'F, ���#�ih�*Z��'Ц�A�|�GZkܳ|h������h�6��8�G*�X׌U!E-����>]k�MH��H�!@ͭx��h���:xG����p|�]-Y�D��Y\¡�*�TW��&QHydg9�R#�#GV僧�#����l�Ӆ�F�dnX�<m5h�<�N6�eݧRHU7��Qi�˔�h���X4�ar���\ٗ���[Y	�F�	�N�]T1�Q�g�(��h��(�u�!$P�(��x(��3qݵՉ�&�SZE��,�/.,�@���ŲY}�=�ʗt��T&U#fъ�p����(�h���6IR��U�%P�*T���D0�J4&3�7EQ$ܹ)�b8u?/�:&7fp\��r����p��	���8��>8�*]"4=Dqj4��a���l]:�9�c����CE����~:L0�>0���	��`���0�:&�%�L���x{9	���<>���<|C����?���`�p�8M�����0p�`�>Sk�1B>8�<�t"ʪ����	�cw���ڈD���rE=��W��*se]���w�           �B�A���P�l�D�\���!w�%�VN [�����V�1F[#N�dc�8O�ӆ����⣿65K��ݟDI�F�9�Θh����Z�>�rʮ��$���\1CI@���R��b�[=��ڤ�f�w�gt�L,l��)�\ᣒĐ��ÃmȖx�Uժ,KR�rީ!�p+$�u�Yv7$��X�evTE"o������n���
��0�ޟ{юB)q�R�zG)޴b�a�.%�k%��UbX�ݾP~�P��	̈́�içl!��K4tQ��`��7D��rGE���d�s�$&xzt;�ѵ��D�#�!Άꤢ��C��5�i�H8�vXR���Y��2l8inP�zh�|xvP���u�:Q�k;�[�e��܄O�/�+��	�v�"���%KE"���֌��\45��M�Be˃�K_l��'ȱ�.b��i7��,����Ga�F���Z�wʰ���g��+�]�*�G%��.��]��^Wޣ����&�Vr�����#��E�] �R�,c1}Ѵ�pՎ[�t�h�����kxj:�3�A��Քg�%SF��,&���6;�|?3b>�Z:�G�.å����QϨ�Ful⣅3�4��g�|3���6����ш��G�f����6�"�m���vE��g��N/yg��B�G��ll���Z��GnJ���t��G����RRth��aб�3�m��b����&����֏�o�2�UQ�C��-���1�1W)h�ߓe��l�:�4�\D/x�i��X���lf�ǡ���|aF=O	�+c��&�Q0��1F��!��	����M�#�8=�'�����`�x�����`�p���x����ta,xQ ��������UN<>�l׷�aSnȤ4j;Ƨgq�X��&R,yj�s_��ټ�=���UѴ�Jd�Y/�B���b�,�2,-��{�'��'��Z���O��������+W�eA�.%1�BrajxuG��^����qͩ��[qlJ�
%�x�vr��.��x�rN9U���ܲ2L'5-��	�#B�QG��UU,�!br�e�!�4Tʮ�P���Uy5>6�&�"����[a          �BV�.���dI��mW�)�q��iIN�5-j5SLE�BRU�8�ݟ"-8�[�?0:N�4W��%\�&syK�<0	�\GD�+�S��m�n���\<�|]��p�A��~=O�B>�q�+�-�^x��..�����I'�"qԔ��T��6���!��cm��K83�Q��G�k���:��\�]#���Y7ԒP`�2��E1�7pj�-��J�Θ��h��X�szj��y��#�'N��C�]Jv��m3<��P����R������)�pg��q5v��a��T���6UP��6��)3�}俓������Ҏ�Q�b=�1�~$�E�TeEwt��g��Z<R��Dh�a�k	˒Ʃ�S&�N]e�7�h��]�0��a�������ҿ�����ч��v�7=�!�]TZ-W�mYz2Ϩ�c��r]Si�]������b�����/$�8t�У��&����m��e��d��s!�$��k�;�b�Fm�k���!���_"�pC�+v������)���2�Co��q1���G��o%UUT�Z>D�X����rH�1š`�QO7�rdˇ:K�z�2�9L0Q�a��r��g�;��R�[�m�Y�! t�`��{.��%W61��O��/Ŝ:i/bI�w'3\�m5�"�"�0�iL��V����.��+>8t�aࣇ4ם���)˔Ài���dfZ3k�Ȭ���΢����6������[F�]ʄp8T����+O���ʼQɕ��l�{��W��	��,���¶8a�fL0�a,x�f�fc�d0v>���t{8O'�������fǉ��xx�>�&���7�"�	e$$&ٞu�1�W�u����z����=�w(����哝���؋�c��9JÍ�u��f�H����� ��         �P�iZR�𛤐�v��;��|�]�m���L����z��������M�FCn8$f�Je�P[��8
3񷓔VSO�GT�ѳ+���0��iDZ-����,���r�ٖ�n&y�86l4]t��IW�~<���zJ�k���vYY�u�Ti�l�D&I2	���흾-��k���y�NNg7�l��Z���z��_66um_k����܏u!$���|���=W��4YÁ�Q��Uۭd��_Q�//X|b1��X ���Z�'�٦��6�rIQV�cc!^7��Ӌ刋�Ț��Y�aТ�GJ��*G~�<7�J.-����z�}�lԚ�}jy���a�:�HF�'���:�[�F�2����g�w�I�&�3�㽔�N�JU�(�<��+"�y|�.-#[[��y<�R����a���+[�|��
��h���&�d��^�ȃ(�Ƥ�ژQ�&�N\x�*[�ZX�ɓ��gP���|��K���:�Q3Z�t�L���Ziqۉ#w�`2q�fKةR�ᤸi��[m�t��ìl��<Z�x�~�7��Uq�rS�����X}�yb:ZgC���El�H굲>>
9���ٹ!
�h��>�m��� �M�n�&����	�����/�K�E�.�/��*����ޞ4G%QQm)f��///����:�Z=g9����L�c��aEt�}'�W��#�!�<#0�Ba��	y$��0�,�2�&�P�=�!���x}<N�'���3!���x~�'N�g��~���Q0t<(�T<0��t<m::W2띭k���+_�w�`����wf(�.鞽77�/P����{��ܳ�'��J��<��3�ls��Uf���\�ءI/��\�k	l�<����vD�5�;�,M��}�8ѽ���%g�V(��O����զ��r&-�g�H纍w$ȣ�T��N�s2i������X���-�|h��w�r7b�$�n'Y��bW��ƥ佫-I�W�\�T�M�"vRZ������K�V�=�           	M
P�+JW�ޥDd�[+��5#%�T�(�7d���pd���$|P���_�^^w��o��������	�C�rD�����T�g��5��,S�x�ui|�a���Q���	����Sn�$��){�|�k��Va����G�1ȭz����e�`sR2WZ4\��rlv���ӆ�������[�e�]:v:q��/C��6tà86MKb9v������������&;�n�zC�oj�_��¤��]]��sͿ��<�m�m��$�%���nJ6��4�%!�4t�h(���sһ���Tt2�s��q�N 9V�)!&"��.�F�rHH��갭6��guE��."�0�w~�n�QT�Qnk.ޒ���&!FL�$,��t[#O�6�3���%�O��;�F����h�E��q:<sz6lɀ�Pqn[�h��k;�F&�f��3�#M��:kʍ#�,�r�G�����\T5eBhᣅ���_�w�X�|Ŝ^#9\U���T�|<��٥-��+F��q^�u,3W��HP��Q>��օKxXZC�����
,��ۍξk���"��dx� t�{��������8v���]C9��8���ZO~c��IG�y��q/6uix�Ä޷�D�&�gŒ���4uE�U"��FŧCV#ॳGFrE,��g��,k�mѣ��t��<a��>>��|���⏋(���|h��4a��8a�>0�����|p��C�(Mr�֨\�T�"��ڭ\"����e��tn�w��F�z�RU[���=e��(�:��ڸ�{�-O��2�����	�i��0����;=�5s3����OL�GZ�+�Y{x�� U�fԩ+�9 �q�Q6�A���EL+T�_����d�^�D���e������̙{|�.�e���+o�-�70��f��׀           ��IR�4�6�h�G�iFlg�M��R�۲l��-dois��#g��>Y�YKFq5��a�|��]]6h���0���Z>Z���Jp�r63W�����:��έ��#�G��b&������E�_��U4s�?! �GKb
���uW�Th��6퍩�\�T�Gd*"�(k��V��#�]�|Ǘ�ӄ�i�)t�P������0oKƊ�Mg�m�A�B�ůs��Mm���s�9�t4͞��7!"�(�҃h�V���E#�eo���7*��f�n&q��7�)TT�P�cp�����v"ZgqZ�ս��Yf�3G�J�n�����}ods��,�/,ψ=��H��X��<�1qq�b���Z��Rfdptn�N�Y�Q4#���%�U�WQڧt�;���9���B5�fbx�ku����tv������2/��9?>KEƏ��(��$�|���zn�MF��-���b��K�818c���d�����Ϫ��:W~G�'��ʎ%��_4��2�(���������E�f�0s����>XX����M��c���Q�t�*��uPl�4�ME�T�C���vqhM��(�a}m:jHЙg
G'���q�y�m��������IGN\7s��x��l�,�pش�!���;�����@��C ��kd�$d$�A�B�P�X����|�ҧ�Kߖ'�b�:{}�QD2l�)��EAp@��1o��5t�2S+h�"��2+ �!"6f�҄&�`�������@� 0"� �
 6� DX� `@HXRT�h�`A@� `D�� Za� AHBVE� X��FU������� A`ZzT�@HFR��@l�0 �!)
`���!��L(	�(�0M0��c���Fs`�U)�B@$	@�$dx� F��HHH H� 6 64�,  � 1�* R1�6`40��`�C�������	0
�S"Dm,�c0!0!�T�`�$I$��ݒ��@"@!0! ��* S ����R��� � ,��,$�� ��! �!$@"A���"@"@�$0c#0##�@�$�X�!"d��1 Ą�ăH1 �H1�!�`� f Y� �2D�!����H!1�`D� �@��`FFa�`$1 ��`Ā�`D�`�`�`B�	��a `g5RH! `0 1V`1`0X��R�hH!�����B/`��@��"0 !*@�x	`��
��@� 0 �#��h���
�>������l�[+e2C����+�l � ��B	t�G����6��K~<��q��Ϸgrx��Y�?��Y��xN��.~��^�~��a�?�9�a���9���@�O?��;�ߧ��|b��v��
;���	<I["|C?��~t�[!��J.swG��X�@AC����v�����h��z�� ��0��=���a$ P�����c����a�\=`���'�H�T�)~�'��_��*�������<���?������a�Q>-����!���������A����!���-aSӲ \w�ŉ�A.�@H����}���dK%���b��c����mH��`����BjV(%�Tc�����n
��;�Rɇ�˵�(�B�ai�\Qi@�E �P	`-�@�$!x*h`�QB���� �� Z*"c��rB �C`���,s����6��/��쿙��n=��#��! P�! @�P�AE@�EG����Q�/�������F�A��<O�)���nC��C�O���$\vA�� �(~���;0�R������/m��=�1�
�հ3E	�P�9�֦��{?Y�CʶP~���0��N|t�O�Wd������͡�'�����p��|�:zQ�C�-^*{�����='���>�P;��O<�D��{�����k?8x��4�:x����Җ-�>o!�ͅP�0�@P�C�?x�W��r}�S�,ʥ=E���4�xÑ��<��R��} �QQp8GơD��(�Y����a�\鵋EU,	 "PO�������'�r%�/n��KC���XOP[��sH�)�7v�P�Q���W'{�Q�8	��Á? �A P�A�B��{K�㲁>H���EC���U�ث��~.}G��P����	����t�4�xz����G�������.��OGpz��^�?g�>G�腒����y��>�{�=�]>��X�����������(y����D��X�*Xb��ϼN� {0Ok8�����������;��>?�d�)��'!���6�� ��|��1B@�I$$�0Qu�x���X�x�ʆ	�{}�D��<2H�p|~N���L�='	��07��0>������ m����X�K;����O�Z �t%��e�$ ��o�y�ݞC	��f'#�|6W�#E�|��Ɂ.�c��>a�O�lr+�����}dP�
-��������8:�S֓���;N���AE�O��q2�S�����3M��<��Cߔ??9�S�I}	`���A_wy�)���o���"�(H40���