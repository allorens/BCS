BZh91AY&SY�d���u_�`qc����� ?���bC>�  	�U��@�1Za���B�6�%MSJ��&�HUD�AB�"���"��M@
R�Sl���M!@�R
��D�f��+&�5l՛[lU�IVlU�m�h
��cCR�Si�٤Q��մ�M
MZ�!�*ض�k"��Q�T��-���m���@7�q�]KI"ͫ�d���4�\r��E�CL���T��5�����R�Q��[Z�ZQ�%�M`���5�I��5�mm�mkl&���ղ�&x   >��kZ5�"�UC��UZ6�v�uZ'Lg:���h�y�[�ۮ-u�q�H
k���R)ҍ;a�lm a5�[��lbͶ�&�l���4|   s{��4���V��P��m�<��v��:��A▆��ٽ�B�+{ռ�W��G��OX�^y{ǅ������ă[���uJR�z}���*�M�,j��ZLV�)�  ��ҶҾ�E�W��zj�e����vڶ(y���^�KC��ބ��r��s��>=T(�S��%B�S�}[�uF����t�$�����_c&���Ͷm�*E�m�kZf����  ��}4�q'��}�ʔ�
W��o��%JkT[��|��l�֋�7���kKa����W�JQG���;�X�������mI�mx�|�D�M{��������!��ŵ��kmm#kf���,��  77z���5�=���{�*Ѷ���[�>�*�D��>����m�/�{���z핕���<}�J��������vv�O<�����M)��x��N��Y���@H��w�նZ��6�ʹi�[lR�   ww��:��+�A^�e�=4��M�j�Wt]v�J���8s�^�^�ܼ�#�Q"�{�g����=������YR�;����]���[H�UJ�iYZ�ZhL��  m���WJe������^]�Х�,{�;�J��ju���j���6�)�x�{�������jU����eYX���y���m�5�S:z�w��B��ֵ��h��l�  g��T� *�};�@sŀ��GKw�x���ǹ�@�����+�\��@��׺��G�{�Ӈ�)A�Ȁ�MZmKL�5
ղ�|   >�}�S�'}⻡�
;��z��@w�z�6�s�^  v�z�Q�U^z��:�={���u� ���*��&�ҭ�Sdڄ�UEh��   ��P}Gg�����YހR�u�J(S���CU�y�@�����
�V�=� 6{���A������W� @  5OlU%R�@  hh )�4b���0�4щ�CMF!�E?%%U6��     ��	*��       �=��=UT@�h     %!R4�)�T�5=O�4i��F�~O����p��ro�ʍ?�N��Kx̵�6hwzp�O.�v��e����{��}��f}����|�h��EAS�
�����a��*
������OJ������������!�%PTV㪯�qA����QQ^�������/G B8�q*�U�+�W��%1 ��@�%��W��Dġ� ��W��@�(b1
�D"\H�!S!�PĊbA1D
D��J&$	�DĊb1
��bG	�ĢbE1 ��J!1"D����PĂb1 8�J&!��
�1
����%B�8�1�$q ��ETĊ��US�%LJ ��1( �PĀ	��&$LB*�� q 
bF!T1��Ċ�� S��%DJ��T1 �b1H%\@%B$\B��q(�J��� ĠbP1(��@%\H��H$BbP������:��s�����d�ԞK��v����Z���j�{z��8pu���z��৳[��X/ �c�j-�׬�q�\ 3����}����<.�3}P�F��#,kHG�uCF���G�f�xt&I˗��!.D��k�Q�}y����3���᳒�eФ�\*�
����n�5�$��N@&�F��*�oE�����ʨ0�UJ���h8G��b�ݵr�f�Ɠ�^AT�ܩX1f�{}Ӊ9�.)|t�*v�cr}�#�)]�F�Ţ��b��W�k��˿"��!júU��˸Tg��
]٣Q�0��>rIa�]܋4��51��%��m��!���`�����㯨���%V�u��8Ca���tT�!�q��b�IP�� Y�x�\ť=������U@�Y��O�We�a��n�.\O\#��)�A*=tޡ���=H��¦�������y�Y�on�-|1�6<�,[�:�E�װ�Qoq���;���F�m<�ჺh�unkacV�Uw�7(`��l_V	�B�sP���b;���V,�
�U��5_<rB��}�H:tŜ�nkŝGr]�Vn*�oݺ�|h�"�#r��q��q�foh�����gpʕ�E�ƣx��hru"-w5��2l9�DN��.0H�����J;E�*�S�'�s��"Y�q��K��\:�,� xv5Ӳ裡����l��M�u��Ө�f1�h�E�"�c����j�B�n��6K��(N�z6=g5^f�#��3f���9�e��>��#�v���eG��Z��<+1i�O
�Ej)�����Ǩ�z�0��>2��bĩt1cǈ�d���9�nj�2�)X�?�ю(��B�x��+z5ՆR�M��]����i��+��Ó�ٝ�ƫ�h+{�m޻@ȍ����횡�K��!�or��\
�9�i�xF:�w�Mm��cz�MɆ��d�P���9PVs�(ʑ���X#l֦���JԂ��ʽ��j��نf��Z����S��P���Q��A{��7��n9(����a�E[i��E�\_V`H�hs��o4H㳚A[Jڠ�F������L�ͅ�71��H�m�^S�վ2�G�R�{��4ju�KY8����.����K�ǡ���1Χ8�v;ˁ�u�t�g[Pd���	nnPt�f�ٱ\�ʥ��4�]A��$���ț�Ա�����!�r�Ls묅�4���t�λ[�^��r�"��H��n����/���c2��2���qa�����b-���ǆ�Ȥ<)���.N�rc�Ʉ��Nu��A�f�{��wNN5�0+2��u_��w�0X��Y�L#x��.�r֎*�S%���NU�w����r��w�BgT���o��:��[�ba�wU5�^;�\�-կM��wq�eH]�C�/H*KmϮm�n�cZ�HɜST&6t�v�<iZT[D��k+�郅B���F��%	U�Ie`n��׬Q�vB��>P�Ƅ�ڐ����;o9؈9a��9_
�t-�W{{�	&V��(��Jl�%Y^�Nh�z����DP�oWiQop>�1�$;e�kDd�l!:
v��t$/h�ם�]��,kFE��+ �F�:����wE*�/kr� j��gf�Xȕ���Ge�0���P*)��{���Bh�ΘcI����X$ږ��pX�Z�,���^bƬ�t�u���q~\� ����B4�6Q���kA̢m�H�K�[6�u#o&��f]*ԃ�J�&i7Nn�t�)��k<��<m� ꫼In .���	�Dތ��:�A���|��V*#4���c�qڴ�*���%D�J��
E&�R���w��8gj9��u�������x1���U=ǙK
�yxeXx%�R �����̖d�Y��JZ�ue��
�
y��J����a�{[M���Q`�� ��	xV�j�fWX�R,���K��v�p=����8"x�������0l}��_hy��R�"E���e���;I͋i;Fx4�D\pr��3��"����DẉS�G�H����V�[n�+��ŋ���xbu�k�QA�=��s`���kN�L���DH��z�䙹uD���J���ja�M��y��5�c�<��5�x��C_m�}���8�	�׾�K�a��}p2�om���Kr�Tz���\�kG�*ɗ� ͺ��4b��;�^��;f�HYxBm��m.�WS|�^�� ǃ:o
��ɣ�Az�m�֑ٹ�죊�u��^���`���,A�R��RV�'P%��,h&�o�D�\+w�.��跹n�̽&��{���������U1�)6e��e�ٌ�M4-6�U����yC3Z��e�_3�l�7\�3�IE+8��'���a�)��6̄���9�l".]�G��u��׌�U�mʥ%@��u�=�r͵hk�.^Kʆ�B���,o2ޣ�b���;,�δ�pU;kF��xwkHף(�L����ۃ��z��	ZaWp;��c�K�1��B�ͨ����t!i�N��`��\8&�"���a+���j�<�e���W-��8I�uڒ��3͘�xzdZ8��7�£S�{a���9��^D�m��eR�7"�wEaǫ]UK(�{���%����PDP;�+�RT���{�d��M��0=](�λق9�b9צm B�9�G4E��l���r�����&X�1�ʎ�q����2(������4��W�m�7��MB��Ćb
ӱe��Ūd�;��ηa�)�i5Sg[�Wx3lT�V��U-�;���P
&��l�p]np�8��N:�Үͬ�������-?4o$��J��y�.��$H{��^�(׍s�Mp���¶U
��M{a��;G����$�n����R�������0u0ǚ�/rnN�A���w�ؗi�wj+����#�6�/�tɥm2d5T���M���zc��V�b`��MÌ<i;v�V�ӆK�����3^��.d����h+u2�e�u*�U�P1�S�.s-���'��-�����C;Y܃u`V%6����1��; �[L�������K�q��j90ɭvI����輫x���K�z�%��}%����^m�{�j3��x�� ��n鎾:.����a2�N� �;t��Tqp�O)G��m;tl�ٶn+�b[�cߛ�h�{��4p���!n+�:��M���y3�NC���k���f\�����tq���\��|���Zc=�L�������o�g�ɛ��rTވ���ɔEl��3�k*�ɷv ��: �<nu��Y#= b�Lod#4������Az�:[�d��q���e���{��P{�,3L���РP��-����h��.�nHN!���o��Af�he MYڃ7k3J�yz��ndt�ތ���w)��,�2�rs�����Ѩ�b�]��	��� �&2v�ݽ�؇ʞ\6os�ͥ��xm�t&�G���ww��%I��p3F�q�7�UB���ϛO�D�&�^닡梽��*ݒ��s���H�{�z��tF�26��n�T���,�Qf���݄8�t��\W�ڳ���#9ݴ�93+8!���=�x�d<O�'���]ݎvv<q0�&ӗ�NCrɐ78={+�lpp���RA�!�MV1Gʳcو0N��3R=�L��m�Vv��`-֮쬳u�eGǿ:�V>�Ԑ�굋.��]��wr���{�h,/�m�Y�� ��m]��ZOe��'-:m�N:�[vot�[脢���<	�Y�aVKt3���VV�Ks/�όM�n��
�{�4�1�:9R����ӶVL�:��wKs kCFŦf��k��������pl"�gp��z�y� �=�a^���>�y�^Xi�O+*�К3+L�0�(�άTYy���طa�A���VMfd�F����^�3XQW̞n���d�&^	x��h'3V滥��ڝklW���r�=.'R�E�4���2+P��`8��Q�+U3��I�վܹ~�nE�9�3T�i���y27N��xr�3hXG5�:tƬ�m�L�sH��G����9��K�W8�mL*�h�g`˲��׮d�gZ��T7y��/�vr�O�oey֭�2rwvmU�y�!x�#F�����oR�{��̊dS��)�zi��z�V�al��3\fhp4"�'Sd.=� m��S>�:fHD�-�D�d�Js$���B��>�cs��	|�'L-�R���1��;��w�H��˦��N�x�n��[5�;.�����m�[M\Qk�o�I�pt�1�B�B��e�X �b/O5vt�|�$ՎoJ�؞�|�:B�[�y���u¬Of9�Y�c��3N�׃tB�w�,�V�5�s�.�7-��Jo`�nr�@��j�ڄ���Tԛ�J�����k�b�i˸b����K����w�L���)�H���1�dG&��:��V��5 �P����,D,ʼ�N��M��b�/F��Yo�ՓDh���'p�QǮ�6!
Fz�׍jbfMo\ي�I����&Y�D�����{ݒ?^>��;�}M�v
6[X!x����90�doY2I�8r=0�"�q� �;�#�;]���t��pE�
�L�=�EL�^v7��I_%�ً�Е,fh�V����R�:6L�Hy4�ٷ4���Z��C��t	nX(u�{�a�+1��XH͈�}y��a�s,���(x[���`�st�oMw=����f�ms���1h<ɷ��wH��J�dW�pIdz^�;���bv֏w$�wB+{������j#H�!#�r���WZqm�Qe9.Ƿ�X�oCo���e��`��C��Mbے�L�c��n��m�n'����QGm����=%6ً&]�x�6�M���<Dy9"��CC��v{A	�.w[*g���w�f���<;gsjY�4#6���3ZTiS5A/]��Kk���c�P��A��F<�o�����˝ �_l#b��P6�Ɩ[�v�<��*��b���]1˧FMwrR$�y>$Օ\�"�Y�!"]��5|���`�h�V���{'f��b�۱����V6j���µa�5���
3��JoE�n��1�6�'�V�nM�ѡ�mj���BV�f��TM�g�PA�sq��W���w��>�9D0^�xݧod�_`5���OX6�qè����ⵚƬ��+ZԀ�TڱL\��kV5v"ѱZ�]�]'N�o=OL�������X�Z5���2D�Y�o\��v=�b��͐���i�����u��U�m��fn��<�Gwۊ�[b�^����-�g&����X�yV�M���4zHoXΖu��G��VA Ֆj;�R��ǝ~��5R:���x�u�Mz�/T�c����WC�Įg�e�>l��!��sH��y�VF�oC��ݱ��r�����&��}��hY^�w^�; .��r��v��W�괾���Z�`���{�ݗ�m�[=�}]�����Lh���>8�F���խ�ၛh�D��N'p��9N'�
\�3�&�����d޼��4��2p��%�5<�8MB�E�Rim~��m0��ӕ��W;��I���$�n���gf��r��ћ�j��d^��4.�G�[$��{N�C7.���YYl[8L�+0��$��ۖ���ձw�A���
�O�����9#5�aZ݌�ZѭGrV[Є��sp^����xm��^dZ5�N��nը�g�6w�źF�M��N;hH���UCR�2Ijn�*��(�3f�N��F�š���!p�&V�����9t�twP�m��3���r����q�~X����\��|0�$���Mޏd���bXW]@��^��=}Zj[�Ν)��[��i�����S�N�#�d͐�{V#�a@�#ʄ-�i�B1�a=389�5!�j�:��{^�`�	� V�o;�g';�|�N�p��6Lij;HQ�M�!��FN,ꄭx$Jn��V�B�k�B����Y�	Vs�]۝K�����5�;R����������'����{��,H�A�$��Wb�n���������ʥ��G;i���v�:�ƙ�X�x��l牷���a�U���D�/rb�4��H2��v��z���Hs�\	4j�#�A�������ՓQ�)[fd�wQ�S�B�U+rf<!�����v��&[�<p��ia�>����n<������wv9>��1�h���XL�NМ�w���kO�J���Z0�AX�\e��ۡ���L��|����&��k��U�,�rf=�-��!�Vf���'*;�:�=���b��Q���E[/�l9b�"�Z+q&�n�	~�T��u���նܜp�V�hxv(<�"��^S�J�|S��x���[��F*̮f�<�Y�ͽ�;�*��|������pł�d=���(�oh���7�� ��VM��4ʫǁ��o�І2�F���L�zc"�x'i{gkw�᧪|V�=E��W���z%�0sn\�6�[uQ5N��^�{2����g�%�T
�31&��Z)����5�Y՘���o�dS^��D��5�Ss���*�
v� WýT�V���v�$09�g-����pN�K��e�:���|i-�r�G[QwV��K��3$���g��ٚ�g������{�O�������{s�yz�!﯀��*���컈N���yH�3�7�'O@M>[�����3�mN���]�@fV9�v��w-KН(���O�g��# ]Aۏ�*�0t�<����G8��z���;�aݘtao��rɥCn�: N�J���.�ڥ�K7A�&;�nG��3L���ex�$�I�-%�vF��}ꇮ<������Y;羘�HSv�;���zs��9R8I�n�J"�k�<�=�as����c(+�'�O~>JY���Cw��~i	���i�خ�-�3wc���K,ْY$�ڐ��&�>:�mэC�#"aL��yl��.�q\x�h����b�K��_ݻr��'5#f�-���w��>��Z�ׇ�Z��w �v��+�_D������e<��)���H�*cXCJ:mZ�<U����w�"\���b&7q:P����|�;�W�rjw�s��/u��WЙ
�;���z���,�Ԓ%��ʕX#L��p����<F�5fń����{�f�l�P5���g��Uyq> |��T8�i���G	B�*�Im�iF��Vk�/^~�d )}�����g�-�ݨ��WgB�/�/������-�Z�5����L>��\x�M����ֺɔm�#d��
��ѣN�ꆰ�gnd�|=c�8���^<��,|L{��[ۂ�^[xz��O@w��w�t�����=���!+�Nк<H�9{A�T����1k/��jx��%�N8�6�4;d��\D�q�PˮK�\:���uq(�;#-�ie v��9��<3"�""g��=���Vk#��o�rή��ӵ����{Úk&
���\n����6���0*ȝ(eӻ˴�zhg�V���59�z`"��@��l��ک��[0ƛX1���"�z�
�[�P���<�=:5$4��|��N�8���d��㇃"���C��j�P;�hc`����@1�9�_����}�&(��֝��.Ouk���Q�֖]Т�)�׾����yw����^G��!�m����`y��II�v4�T���d�_���5Nv4�EwE�0姙�/M�����3q� 2���FtJ1]�y�Ss��t,��)N�&��뙘��rJ�8�vr�l��B�TC#f����5}�3���� ��xG�Y�#��8�N��/3����o:W
�\����sh3r��x�N��k��M��M` 8񷼬#r���
����8���xi�
�G��Stۥ�+�&�S����Z�2�ph����/���4+q>ʅ�V���%�M�����7k�a[�y����:ݑ��`̓�����cO=y��u��H�\��0G��M�t�$�yur��#���o��[>��o�L���������L�hYZ��X��Bn���v=���7��܅1������[����n��:h�{����+�-^�����������h�;�o�Vu��t9JD9`U�.�Sy�YCxS�G�9%����7�[Mgi�d��,z��pE띷-���7I�s۾^r�ܳ
�<W��A>>�>���bl�qJ�&�h�-�C;0�!$>\�lӭ?JH�IhA�8B}�<�:���Z�!;�����6PG.r�l��W��}����`T��/�'=P=�Ɖ�<�It�+8�NPõR�q��K�gOF ��^�i�b��Jb܎طoFU�Wo���\M=;�88�J�����֡�S,^A�%ت�
�Ӯ�LX���,2�[�b�TV��sz������b{�yݝ}������֒��%�c�X�5Y�Oφ����g������^{���t /t�͜�]n�����1\ vއL�٨��E�45v������Ɂ������q��-� �ɳ|sݢh�q0�RE����CI�Ye�ZTݫ[ʧN�2wM�ޠ^;�smHͱ]�3su=[X�Pg;cx�m�$��'	�}5���e(�
6�lN�j)nɤ㒴ЭqoH���r�|3Q�9\���3RrE�2wtΓWf[��yV�A�@��R���D��5�L�p�vN��Fw�ox)C�;���1o�%W1��Ur���ʷMs.����Ggc�=~R'uQK�U1^�&X��u:����C���v>,1m̪b�N�˷��v��j�%�b0ܲ�����7���8�g$�90b���Z�Qn�a&�4��|�R���RP��+�=��+w
 ��i3���wM��J�X��/����j����65c�"��[��q���$�#�>}2��R9`>�|��R��GU�e{�5u�����LP:�r�ΝÎ��ƟF�����|�뢯g�sӲ��pb��tU�eX�i�^���`N���v��X
|'Үo8θ,��X������ꆺf���2�٧߯�"�p��uh�S\u�0"�V�<v��kG尕��ٲ�b�X`��sD�I�Ӟ�z����9�͂�X�[jm@�u��V����&��A��P�9��S���H쏍��[�k��pb��x��q]���Cs��o���w��¸���6��q��">��0��A���>w;޹�ԯq��şKTL������k9��#����.�v�w@�M��n�<\t��t��Wc�U���Y�8Z{o��m.e�@m�F a�E�j��.3�v)��h���R�mK���J��B[��v+��R�u���7f�Z/.�s�oJYcl��^hә�]AeBi�Y��kZI�����zИ&�릆S�CF��k������,qL����[��p���~F���9���Tu}�D�ݡ�������<���7i[|�mI�2K��ʸѵc&f%p�����U1�yώi��3��6'G�% ��Z�3 !�ڄn���"�6\@e�WVrìG)S�ƕ���d��vt�gw��b��J�;�u���'Y}���n�Y0p`�gv\����T�ހ��F�7y`��/��ٯ*������3�05qk��Xw�	����v��uٜ���[��Ɠm�g����/&*��K���9�'F�(�u ��m8V|��)��A~���|N�6#�\�L��o�;t�}\��tU����h9��B�K1��[iv��e	ө>���z�\nT���Ι��-���C��i�9=.�K�pS�L�E�^���;��^3�K�����VDmX+����}����Q���~��}Q���c��0y�6�TTfg�lO�������4Q�֙yMn�o\]pHGv�,[)U�|��@�wK�i���!!�;�x�b&-�I��v��I����۵�z01*v��R��_�,�l�$���b��5T�Nh�T�/Q\�غ^^ݪ"4�"��و�	ծ4��-�j�w<�61�k�@�[�2F����@V��b-.���Z|[<��w�+�k^�u���p�w�-[7 �p�)]��-���v��O#��*T]}���\���'SzE�E�^�r��E�i.����&{Gj�5�a���� IvQeP�D;-#s51ah�	��Ĺ����K�훇�<Ǿ<��n��ˡr��(��X�Q�TAN��C{k�y����m��m���6�� Z쭭':���6p�.����K�/Ǝ{�m�m轡�^E�it�����VS�m��8{��}<pe�u�:�eb�ވi�Q{;�׽��d��M���I�s�&�Q��͋�j�z-<�tL�H,ȕvh㹈Â�18�����Z=��x�y�sG��z�>Q�g��h��oc��%���K�9���엁+e���b��g/��������
�ZG7�K"�yru�=��Y��÷g�i����[h��K&�GY��޽��a�I*+ѩ[�FS�q\�s&��<{�ܦ������(6(�H�87k�@&@��>�o�+�ٕ� T����|��"2�C��^��u�d���
���q;wם�,�wr�I�
N�Qֶ��6]a�3i��S��7�b,�2���m�}b�p,��7Z9�9����cy�+��$^ѷ8S���ܓç@��v.$���+e�z��/�4˜%P�Ϋ�q��9�\�PZ�mv��eh��OU���Fq�WS�&@޽�=���F]樍�l�v���{��`ͭ��qL&9�Y":O6n�ϧ��s�kE��o����1�[Mf��L:_j��w��GH]/zr�B�{+�9�E�W��=�c�K���Y�њ�4N�p-L|�:X���w��0�~�}=7�� ��_,���Je����,���mN5�U�2'\9���vk�I�H&I0� �s��KMB�����Gv�2@f&��Ǳ�>t����I��ѹ��l@n���	�X�6��P�KR��t�U�iR�0�tϱԴ�V�q�����	�:����i�6�L�� ��\�mO���n��@�p]�"������j�I�&;;��z�s	|�S,���:|X6��ą����W%��!��.��X�MX�iZ۫�ΦomNu��5@n�Pۣ�U�6�h�trC�[��y�B�:��$y�X�Ö��v�G��ι����o����d����\&^ۉ^f����:*{^�g�X*ٻ�	U�d�y��}�X"]��@���m��0q��Xa�ޕ2(h�y�$0[1�\�����G�c��SRp��y�\�r)*��C75[�Re͋ޥ�^45�ģ\3&h#�DM}8�����mɫt����z�B<�W���n�ج37�hY�&��s��罍��;�����Z�}�9�Q��-�޺s�<�eS��H#�|�w�=��v���פ�ʣΞe�=,G}In��l��tI�B���L��|��<�Ns�T!S͡���)�<���d+_�vr��FL�Pw;�;�kvv�۹t�^��h����DѬ���h>N�J��/dk��}�|{�ʂ���9u�Y��n����_9E�ua3���V�hZ���#w{N��cy���]� ����E�=6?�O��߹��W@5g�Oydq>��뇖��0�^��9�R3xW�?H,ތ�pc��({�Pp-r,�qu��#����ג-�l��:OVW���2/�U����r�k�`�O�>�}���|Cf#�Q|�GKB�īw3E�ٝs�Y��)�T3�a�n�z7���8���||�)�S�&���7e����-�y��.�Tf5�Eil�<c|:���Ҩ"_)'���}G����.�ԛ�B���&k��zp�����'r���/v���1��>�������\F¯��`�j��ptҴt�4�@��Ȭ�Mö�̕'E1v?���
3o��͠5xt�SLg\��I�ŀ}�2z��V�][�NWWv��$�ލ�ǏnWE)"$m<�G
cgT�Ԯ��⓵g8>�o]M�V��t��ո�E�J�7seZ����ϟ|'uT5�>����J�g����_H�D�s~��M��5*p.�7��I��X=O���v���J&�^���n()����2�Nޮe��V;&��:��#8�:m��ۤ���C���G�����t�3>�]��m:T(#��wp.��VQ!� �;�ƙ��uAƜ�ڸ��h�?w;�	�~�v�����j{����N[��Zs������JP�פ��w.��,ܵ�d�Kejܮ��\�<	>�����.��A:�, ��������o=u���-��{���x�G� y�^����b��fE��?�;;}�tz�柵%�h`��ݥ�-�qW&��B�B0�ʻ�-ֈ�q��-,L���b>Z��)j�ù�7�=��t��6���n�Ÿ�qԂ�C+S˫�J�9}s�����@<
�ƽOgS��^�!�g��jm���K���Bn<��Г!��"[�[cmG��k��;��m�|,��Ak����gj�;&M��H��oi��3�e��QmU�k�I��~�+I龶��&�0�9�/e�7�������f���Ev�{ƫ��|��Al���cj� b+:n�Ci�E�}Q��(9 ]��9Yu��7���u��K�v%n�Β,Ρpk j����Iw�9�P������2����
���f�R�X{r��/mtRý7��d�i�i\޺ʛVW�d��dA�wԳ��7E %;zr�����.ӱ�r�K/+� +��E�g�r�nIݷ��`���4;/�Y٧����!�E�[A�vn�_2QGGX���G�:p�Y��7�M ��
�X�z�
��>x��د�s+��]��ͧ]��}tQ`����i�Iku��x��gAG�@�V��M�O��!� ������9��b��nEޯ��,�uv���3NY�����^~�v��o6eU�v_sl��U9�T�a'#����g�t���yy�����G�$��o0�F{"H�o7��"w`�s�w!ҳ��Vx��~en{�})1����9ړ�S����FA��CO'��o��,��t�ܳ6�]zt��ʲ��V�Q�<^�ݕJ2ǅ��N�b�t5�o\ݼz]J���u1�6!PN�Of������H�;�(^���!�>�x0Tz;�]n�_�uN��G�t�]6��x������e��p�ǂY�v��%�Yx����#F�U%��3eGBk��C��\���65^2&4����p
Q}���Q�.l��oSNE#�P�N�J�9rd�eDT�9ǳ.��I{2L�Dٛ,�)Z�d̒9c�E$�'\�L�I:I*G$�I�I$�I$�H$�I$�9'%$r��=��rp�;��H��K�'$�$;$���QĢ��V����ω=c+7�����:8G.�D<r��!�o�����t��FfV2�u�CU8�� �(#?�D���1s�yw�(�wy�;�>u�O|�k�Wx<��}g���]V�WQ��Q\��]m.O\�w�����p�m�I�B��L�0�R���! 7Du������AQa����  ������_�����QD���/��C���&�?��?����?�v����o	��x�:|�����ӓ�+L@o���k���Z����&���|N_J�����%��4�gm5Ӧ{�� �*Zr�ު��{2Qq����x��7�钎Po���ʅ�6�m��c�0��&b"�y�ɜ�(�{9f��~�
i;��o�\���:oLb���� ��띌z'f�p���=�s|�R�Lݱ�k��/^n0Bߚy�õ.p�˪�������6�o��1�2񌦓w,9y�z�k�z'F�B1R��^3�����[����qd`X%�l@�>��	�@L]^�kwm�<-/̏Ş�XZ[;:�Tܸ���mX��+s�1�QY�ӹ�܎���fP�o;'am��%����֝�;ն��wzF��H¾^��e�w�M�vi`������J�W7.V��m4�Sx=h�V��)�b׭��G��@�Q���n�`�ި�\��<�x�k��n�^ޔ��hi�rN�L=O�i!���V�T w��n�
�;������ZqX6�=f��ؾ-|��x�S��Hr����m�S���/:U�t���
��U3DT��k(�6E���	p>�!�F��~��+僸%�`���v;��(b�c#b:VX��d@V��Zϋ�0Oog{���{���1�����3%�\:�5iJ�pX�c��D� �"�� �#Ah �(A$H ��AAxD � �D�}H5w֑�>&�{��I�e��X���5��*i��/���xl.u�\���j���N���{�[���v���j��>2n6�^t�{w��*Pݚs�Y�{�WƆVJ����Ϝ��S�˻|󌹳�py�w����Ը�һ�݌�W��"�<xn8z�������g��?z����wa�j�^�2ȲE/o��b��Ny_w#�G6�\x�R��%:t�{z��K�k�Q�>���*;ǈC�<�������l�����&��'���_���:;����s�Ǹj��a��kC�.��_����gj��s�ʨN�n˼͝�pז²�Go�]hwC���njܶ��m���f`�X@������}��ӓ`���q�x��m��Ib,�ya��hu�eम5�wV�*c\���Thu��d�)˵>�Fc��*!�N;L��������x7�u|���g�yӭ[w��4?�Z3x�&.9}��8q�I��i���k�á^ǫ�*�5�%�y�� �/i�^�>X9;s�%7Ì�=�>ӚKG��8n�?{7�� ڞ��d�R��m]���Ռ:�zU����!;G��=��z�ۼ�l{�����*h��g?����3��_2z��[T��m3d�pK�·���KN�׊�j���Q�L1��4ÁA �A �#A@ �$ � �<"AAc�p���!����Z������>�v�b�S�=��,�;l&X˜��]%�]�'l���_LZ!1�=�WX���׎���O�.��Gq�����zj|�O@{֛և)��'i���D�]f��_n�zS�v���K|���]%"��`Inf�ޣ7	��q[=ݛ�I�{���AT�k��"���e��{��g�#����J��:���C2UM���J�������H�hr[ۭa䶹�]׊n9�c	�4�����S�f՞��U���7�*��zv��{�^\�wW��;���NC�����n�NΩ��*�.����B	����E^3h�+;��W��gw��^��.�`�"�[➍�׽��0�i� ��̔����:����og���5��IW�{E��=��kc諬Y��Xs�$����I�K�:�V��$f�YÂ6�9�vOS'Vkoc�r�Yf�c�:�ݡc���}��f�aHт�i�����s)9��cq����;[��˴!��͋�ɪ�*�=:f"w��z��8dJ,}W³5��@0K٪��*0�I6���� ��u�����9�l���z
��<�R�
�; �ot���r�n�z8:s_��`5|L:9!x����z=%�\�Z��u���#�VG�3n�xC�w"�t�#ʝ)jL�]�n���*���c�����UW�4�Y��w�'X�1�Xdi��WUYg;��Y�(�1vFƇ���$�1��f��F��O���)���'C��y�l���o���vp�0��Y#_���(�aޘO�|��|����V����\6�]u
X��n���|�|�W��l��d�[q��%�'��������D�gSʋfz��l,�*�?v�sX�g��O�)ɼ��o��R�%�5Q�@K����Ϩ�y�]�u�=���R���r�d��e]�4����h��(
���o)-K� $��v����r=y	�>�[�|LxH�^�8�4H�뢪Hoc�1�^�A��,X$U�����wqP2y��U�RL�Ʋ<9��մ�kU�]��g�n�bч�7]�[r�)I�j�ۭm����H�漱ƴۮ��;��3jHrM�˝
� �T�)�0u��w�����Fs$Kj��,˔�q$���4�){��g;h�E���^	-���`����P+{,Όk�r��}���QE�ڢ���zlFv@U�S����W�����g��g�p�;�|��iǮ"�˻K]R��gP�s�n�a�p��:�s,��53�b;�I9�N��]������Z�i���Ps�����bg�6��t� ���yvk�]�Z�u�:�<,U!d��2������Ի�Kl8
��:��i�{��<���"�:P=:ŮȻ����y\�y��w޷�S
�r���W/���<��1ƽ� }Ϗ��|�F+�.���/��z���P��+�b^�~'��<]�'���+;�p�ǟ:j�(ݮ��3j�����Q:���������2�ЭmM���վndg˺�=����yhȼv�4�G�����l��8a5$��k�"��q�G�۶!�6 ��>ڳ��OA��_M���-m��$������2R���qIJ4h��YCd}�cy�4p���Y\X�Tٓ˼6��y�IFU�s�ޫ tpLg���L�Dd���lmk-Vޗƨpńr�(���ۤ�������jM������s�Y����=�z?5}%e>:6|{�FKަ�Ô@i�o_0�*4b�oA��Ӓ��W���ԥ�[DU"�X]˶ :ޘ^����i�Ք���}�K��}����	!�}�fb�a���@�����s��}ج�o�<���q��D��s���OY���c��qsR��-�Y;�B� ��0s�s<D
�v��I�9q��f�}�h� l�ߧU�Pr��0&K�Ĝ��㼵&���2Qי,5��"m�]À�w-ə�M��X��r�@	�,{%1��3fc�\��nu&4����3��Zřz3���%C�k$�j�M����)S����m��d�]y�It*�{h9�Au2�o9�υ�dF��L��9^�uKl]�������	��m����xdN�B����̙c#��ܲ��ߌ�����Y]Y�U���rbY!�����g��=�d�{���f��.���Ӝ��:4S���{��r�r�v�9�Oe�q�h�u�=��7:d��џ
Hl�$�Vu�BLQ�V	����X˻�X�}�.��n��An�������wܴ&R����&���yp!g�W������{=�w1-Zt�-��'�-�9����k[���\ [s�_yp��Gt�;l�ty2�v���))����;�$A�	���Q*·�
�*#4�@��E��]����ʃ�i[�Fn���-&ݟ4��3A"F��h���C<S������e��fỼ]�z�W�0��]gv���Nvc�DÝ��gF���%�3�20��q�b3<���%�]�sl�;'��Cz������[���f1<����S�!�@�7�'��+E>kRHs���=���ǯ����V�������|i[�C8�ݷ���!y�;�f"A�1e���K�%(��5�.���u���"�P��3c�Y� F{��g�q*u�-�N�p̮!�Tö���fW1\-E՛:�/A�ܘ�Vx �,�;�4vA��a5�Y/5����%�:�S�oM����-��`��!+qiv)-��g����>��~�PN����㻱ݽ�4ŗ��}R&ޕ��=z5ɖ�ފm��R�z�R��Ï^��t]�8�n��-g��dҧ�EW��+���3|'�}�f�a$!��:����J*�R�,�ڣۄN����qK�N<�X����$u�۷|$��Al�b7-�y���o*H�qn5K�юo�*��eF@A���c�c�.W%���q+�}�'j�n�~��:�3�����N�U����jr���c�#Co���JmPyiج$�oc�d�f�,6�|[Y��L�fj��z�*)+�����t��OW^������*�`ɛFPkZ�o�gr���lHuv^㩤N�n�������^⨰���ͼT�Kf�
���>2����p]fD���urJ�Ej*ܼ�}��g�����΂�g��/vN�-]V^y9w��ze���������tc><;����L���Hm�=�����ZEɑ�Iq˺zg�}��w��l��Wv��O�$�x�^]T��B�T㽨xSx�`�}�7�|WH:%U!~�S}��ޯ�$8�"3��F�����=��;���y�)�͈�jQ�*�r��n�&c�p������/��x��RY���s]��::��{.��N�8wV�)!6��wm�e���y�_x�x���N�6�\;�/�G��a4��OTl��W��@8��Gf,�{9TYmLav�z��}'��n�������v�E�ҝ�:�_���Ś�vm�x�bE���ѫi��+������bt�v�)��u0�(2�]���sgc��w!S�>���u��̑?)*�b��jNՒ\�{g*/����x��B����H^Rů�(w'JT��4�G1������r7Է.��C+3q��hM�h�FYrl�W��G�1�}�h��}1����E��Gb�{;=��-���xM�Rn��4����L�^A�bt�G?�O`�u�}�YT=��p��=�ڰj�v�B�H�ݪs��bʶGG�<3�����P��v^3�f4�6�x<����#����r���/��{�U��:44NeR�حD-<�a�7�*| �)��^`I�.�w��MԘ0<�Kr�GBM���2��ՋG�C���G���8x��IoM6�I��K묉U��h.��N�zu�u�ȵ���^�n=1`����oC׼Ms|�+/����+����T���*�Ȯ���g��A�x^>;��ղUl �\���C��t�Ky�)�σ^�k�W�����ҦL� ����>�(}^�cؽ���[&�Yr<��'��v�=��}��6h�(>��1g�� x��8Oo8A����dH�W0u�H5b�ſ��E^�x��h^c1�͍�B��ZzFD�4f��s�m�eզ��wA!e�`��Zhr��w���ݢ��R���R�6�:���^r�<�F/D�X[g5L���n�����:��#l�6��ݘ�	��@�մ�َ�zR6����;�l�/6t�g)ln�%ڷ��ѡ��K�hfN��8m�`�J�q�WQ7y8��nӒ�ɻ�3f �\�dG5�s����ʙ=OM��t�.c���慶`8-���!ȭWմ����0qd5�)*Ż��smbxR3W����!�[Z]�s2��Iw��vaCl^���8���@Uv���g<:쯬�gk����-]�����fy.JC�M���I�� 9�7p�lP��j�^��qej֚X0N��26I\NXIV�N|��᝖���1���׳�k�o-���8N���
O����!@V�w_Ts�.���#���*�N�Q�W|�A��Z8��v���J��ʩ�,�l뾶�Ӡ*��bL���j��~�řƞoCy�����t:
t&C�ҁx���p}�]�o�w�()��/#�jH;��ȹQ�0��:켣����ܫo6���a�$��йww� ������U��)���9��R��n���q�lp1�`����q`�m�<��^� �;��vx�	�7��X�X}H���X=}X��/f���w��i<j��6��]���c`��KC!G�j]�_�
���~��<���>y��x�˜i���[Ưj	�Y��ތ9��]��)h��83�u�m7^-���j3$�n3�΅c�U�X�m^�q�y�����fX�L[N��=+Уf=�H��iH�pLwd}xp9���vz��Lu��MZ:����M[�7=�U,�wq��D����c0��{�*�Ww�nn�Q���q�{�����	�$�Ez��Z��
������?>�v��a����0zF���������	��n]r}������α{�$��&l��.�/!=�6^J�����Y��]]��)���:n/}��<�ֿW7��I�q)�4���J�ci�~�QFY�/9��r�B��p�VЊV��`�K�A��-V�1G�{�7ۆ���Pn��P�:�>�#�FM*uH�sL�ᕀ�)���[���٪S�G�h��R{���%ꙨL�R�5�Dhb@���J�wmv[�Ux�Hi����HLWV>�pD���+��PV���^,s`�*�ez���++���Ϩ:Z'v�yZ���<�X�h��K:�jk��F������OQ�3�ۢ����{H$�l�n%*,���b��\�%���Z���)�����%�'Nm��{��[Y�{���]�&>/g��{�2�H��E�3M{�z����EQ�&�;���2x��\���ӎ3�������I繺����_�U��s�BP�}�����x��ea��zw`�X=�����w���_�?p�*+����������?�?D������t�ߋ����w����ZW塈�B�n3���3���5��J�.UMڙ٫0����}�W�g4�ݜS���#S�K1\:�a^D,��_�E��룩��Gx"�˒�g˄�;;�s#W�ij�(�1�p<h��#�{*���VJ���۽'CU7r'כ��*a��$��6�Ok�X�5�� !Xw9j�th�jH��3
Rad��l�7 ̢� 7=���w׼߸��w�`2�t+:��	I�-����D�9Rn_k��oi��#�j�9�,\#�_l���]���1\v�^��e�[�#<���{����岸T���]���5�OJ�]�<�%��w�S����SsOA�P'��^ިt�TU`��fd�ʕ&\��1B9��_	Y75��s��XclӔ�uh����-�M�/z��;#׽<㇆s���ζ�?�!��&J��V�p�Po��F�Lr��4��՜{õ��K��^̅J���:�u���������^Xl�{FnDޫf��J��%\��{��.M�J���c��y���G  �z@p�JＰEt<���\dg�@���g=G/V1&n��C�o>�T��̎����Б���*|��s��#B�(]�X�̏����>աch���S�f�_vh�.Y�	�}�^쁉5P}��RY�«�a�#6�JR�$�I�	��5�a� /8�P8⁨�J9"��P܇�P���- ɒ ��4`DA�4A|�OV�UT�b�h�b"���������[Q1mZ���kY����::=��	���\q��AMAu��TQI4h��U��G:��m�����*�cph���j��5�,V��(�*�b*�h.��L5�D��E$QA��<�;b+m4��T\�`�4Ӷ""H���w�MNjb�m�5UE4F��jH����QE4U1]lTUՊb(�14ES�L�$RD�T��DG
��SMQ�ub�*�ֈ�����\���	�Q��!���`�j���Ur�<ŃTY�$�l⪍bѪ*
��5���/6��F����Ѵ��" ��L%6�c�A5=����$A��N�b�"����RG,�m�Jj���F*#F�����j�7{�7 �M[f֊N�TrtTFؠh���-8h�Qj�l�j����j�Z��d����u�TLM���%���z,y�����WϞ��d���}��)��uJͦ�#�
�d5oz�5��X0�#.�YJ��Z��VʹlΨ �G/(m�(�H4@�R��) �]Y�]��y�I���kg��v����74��<UG��/r�	ۙ�]�傽]b9��+���n�F��:5A�ם��>[�}��4�I�+��#ؽ^�	��E$��V{�x�]�Y��Ufe�/��+66��Pۊ!_����5�4�gE��ތ���^��n�#�</����T�~��1������P�������䣓}l~ţ��ľ�7�vz{5os�bD��ۯ>g�E�E�@v��k`}'�0D�x���ՁZ�	~F9L�o��� %���F�e�q_�쮛����t='n��pW�y�!��zV�"��N��Svz\�a��Uy��U׼�%{~�7����/`(���M��:;����W#�̶c�3|3�WS��������S>�����)�k.���u�/"0Vӭ�܍�eǫm�ox���W��s��=��J��t#E��}ӄt�6�ٓ�૦*U��M�%}�վ����W����Ѻ�����&xxmu�]�⯂�DYZʘXg2s��r\�a'�_vm%LdL��RZy���/�2�y�8��_P�=��Vi���yŝt��~�w���=�Q��|��i�\bϪ�t��X��K�!jYp=62}�>J'��9Ww���P����@�e}��ډ@�!�e���}_�«��x�n�99L}�u��̦�Xg{������վ?<Ѕ�׹8�v�Д�L���s>�}��ϳL��->A}c�	��j������y^̒{��y���G�S�����E�n,ϩ?W�i�W����W�e�G3�b"g���$�٫Nb����(����Hoo�"�W\r
�w�~�}�4�=��e)�?p	oo�O�=yò}y� W�	�6⒱��,��rU�w����F�����s���WS����V:$���5���~Ɠ�t�/��z�k�\���3��H�"��֬j�N��T�
�)���h7�<�Nb��;6����^�מr��s���i������Y��:��}�b~�V%Βr�h��u�s5��O����
����(��45l�F�{Q�"_-��{v'?N�Ox8��ԝ�跚ܘ�tE�����ͩk��@4cݵ*$��hW꾩ơt�v��E���b�'��XF���jfmn�����{��<L�aѵ���v�`�^��jԁ�H%���7c*�L�M)����"�z����?m�y�8Y/�a�ƎfrD\`fG��+������ŏ�F�r��t�Ҝ�^�T�4i��CmV�ќ$ef9\�lw����[�}�9�j�?��;�3�ׂ���{b���-*�(���|��ԑ�	Lm�w�Oh�A�
������o�+Ɍ����h	�+>��]û�y^�*]����7hء���&�$
z,`�'D%�H����}ӛ�U��	o�?K��o:xޫ��<]�{�8�=+�!_�y��i��u�%M��s���S�xyo>X��M�ܼ|/[5����.�.���=�Y���{�:�o*W�f�7V�m�&�	��.3%�8L:^�{�cu�]N�A�L�t��@�3mf-���Ё^�B�L�Wݖ��PK�՞���>K����I�D�>����R���9��3��4��賳�e�7���B{�շ�j�Z���0�uW:��
�d_%�r�յ���
�*6
���m���/[z(���c��?����^��M���j��r$-�IJң^�vm��ؐw���M�#v~�����1���c���'~��JK�8RşR+2}�ے����I�.�����qv��5���X����R���=�ZH�)GY��^Y���ҩ:��˿b���H���C:��64ҰuM�J��"�e,��ٖ�c�7�;h���>�����J�߄��'�~�o�ޞ&v�Κ4�ۣ��Ż�y���#݉��B�6������ɬyڥ��
Z�+Rc���~y;w���7��Y7i�A})3t�2M�_���9(#�����Ԡb��gg�.�
'0R&��`��@�Kԯ���-\yt"	�4$.V=c�cyu��#�B�ӿ��{t_�
�J�g8�� :�J�x���U��l�b[r��c�;�����\N��D�{�z��^�y<2��=@�;{8?A��P�=P���=�� �c���k��:�4ã�<��h�y ;y^�Bqv���� ���egL��'E���WU����-^M�8y�=9�u�wYn�)��h�������.��f�b��~;˄x�Ê�V������y��/W
�2�<eo�^���ۺM]pj���uke�CY����Z�z���T���!�W]S3ճ(�w���֗���7%��+�
��*$�j�`�
�Z��DP�b���WT`�gD_�YYѥH��]�$��Iae�qS�[Qz�k}�mT�V���!F�
n����`�,'H*��W�`�C��,�S���,C�W�#k)v��^��ZK���zK/u%b�S����RB󈯻WX�@%��%�$n$��!��乾�TS���^��*�u��E�g3��R1�W�co��%~�;��yLP;���Y������Fd��F���A�"ŮځZ�D�}yb���^�=̷����l�ד�a��|r�^��t{ �4����J����̑ڻ*27
�����Q�� y�?�]R-��I����᱌��w�{��b�����Wg5]�Z�	�Y�s���mN�k��}:��p��u�wO�W��`�r�75Bn�����]'�hYz��vTᚧF9S����R�M�(�7�N�g����{��e�6o��d�}v̋<���V��H��1�@��z�GO�F��m�u:���+�О
���}6�t5�v잘w���>l׻Y�tM���l��s{���?dͿ~��y���\qBY��QD�`�M���`�f�9�ݫ�*��죬g�<4�7��Ale���Y���]X*���Ϡ�`����w����W2U��X�W�P��ey�J�}<�k�V0��^�u頶U!+������Ta{W�^�>U�ǶS���\EZ�G��=�N2B�����$,P�Ƅ��kh[+ß���VVܮ;+���ط�^^�מŠ���!V��!�F"��b���yy��љ�,�!��@X��{�������) �ش�G`���b�
�h�DلQ#r��7�s#[|0R�S���An({7�	������%��,'�w���IoW��]:C�	rZ�H�3�T"j�L��;W��^���!��	���-�|�X�J�������P�s!=
�r������t����S�V�mo��GzM�d����'��dw�Ie>}&,8j��Î��<��Y��x�۹W+sbP[Z)h�������+v/��^���2�G��������rH�?++#�4vB�y(�#n)/B��?p�֡�+���V��`�����O���	�>޿�rU�	e
�F�bŚ,��8m=Υ��S>���������l��y�&��L>���ۛlH:N�wG�� �o�ï{mf�WW�b�D��F;q@[K�g*�՚�wv��������Uם�h7�Զu)�b��[� ��2��ݿw�N����v������9�t�
���Y52n�pAejctj�2W�z�i����sk�*�Mr7K����)˥����j����^�8��ޕ���P���{���P����>f��?�S�^���B����'�g��%�S�4�r���>��������ǯb����|�g�q��4�ج���M�b�y/|�<�l]��3����կ�{j�<�<�]���&p�����n;�;ήm�M�jXN�ǥ�����*����8��=U�QV-�FJ�E���p��)���lz��rNI��p�����=��ѓ�}�����X��l����^��ռ��?�Ꞹ���]�qm,�{�w�ۨ�����!�TxE|�+�),|�uRc{ea�#���ު��w8�w�W��n$�!��Y+�8*�=Q��|N��g���o��ں�������7,T���wY���.���c�c-�a^��{�^X�>�⊏��F&[k����"Ѳ��g�v�M�����S΄�ιңՈ,[���}3k�5%�i�s�����F��7��^G�T�7~HyE_J�\Q������|���Ғ1>���>��;��s]n՟k#���02��$2�]�ҳ�Y+�]	WO�ϓ>��Om�*�X��ۣ���ʎm��^�۟�#hI����Q�$�J�`w~�M��4��n�4���>�a���v��^z%6~d�uw�-�*r�2��ץ�,;�t^������<]&d�zg�	���e�}дJ����,2�x���a�¦z��u��oN�֫�3_�tX������;Eo�|�/}AW%B'��m�ʺ��I���Q^��l&��p�:Bť����� ����¹4.ҥ/rw(ʈ^{ޥ��"o�}5�퍡}PW��ShY�r��^���\�l��V.�Ҿ����oٿ{VN��Z��S��(z���:��9��u���w�a/ ��A�r�-�ˠNH�]��Oh���9��E?J�7�w�[Q`�&~F��y�T��W�zuOYF{#�D��Z��;�1l~���ym\b�z�aW���x׽�N�N���Y~闈���qy��6�{�W�Wl>�1��&�����u~������;�EG\�f�]Vw/�q!��N�WՒlxF�T�s���Jv��
Լ/�ݱ���ޮ_>��B��
���A���ezk��6,v��5zv�x��xrK��U��d���Duﶱg�O.л�Ŕ}�G�{�&���V.ޱW���]���ܙ!.�Y^������W�#k>�۝�څ;axwmn�%�G������1��c�ڍ���i3\���tը7�Ƚ�+Խ�+�-�x	����v6Vz���;֛=�n@uS٧U�]̛H�Wt���k��\N��{�g)[֑6�Ω.��� �q�]��`�B�iV������̂���Mr:;���G�ܥ����Ư=�:�e>�4ǫޖ=�bn#�N�?U�M��.�w�*u�ժ�%x�Y�J��Qݾ��>t�G�ޗ{�{��'���i`Gg\fJ���@���GY���s�2�	S�>����V��Z#�_ں8�>��.Bn����'O"9�t7��v��ﴨ�WU��ؑ7���}�B��V������o�a��}u��^}H���'N�J���þnf�7�.�&/��.F����w,nQ���`�~��5H���7�C��N?-�zM�g:&n
����+��>��c��Vk!Q�8tJ�2�/ge.?j{��5�F��s�b�94�{����j�s>�n���ڡ����k�Dm��&�{{��H,sY�44bTg�⪗����A�@��{�,}���U-�v֊ʭC۵;q�յ�fkֆ���E�2�V\{6��_kS�8թY��b��܅����I�Z�6��d�p���6��vɖi��uz�5}s�oS�EWv�bV ]Ӕ���k�$���÷�(���*x?o��,���nצ�J�A��Au�Zd�g��h�/Za��@�M�7:�_]@��޹�&^G*��/�ۍ�v�z˙-��H�붊�r��޼��K�<�q`-m��g)����zY�,�J��txf��< �øk5nU�3������	�b�0�˳Շ2�oqos�k]���y�VF_Q����
r^=<��#4Bgk`i~�Y����ys,	\�I�!����E���<��J�[��(��~�c��<��5����7Lb��-Ӌu�| �*JQ�y��x<9�f<]Q��cF	�+���ڙR8��n�����
ʆ^J\"/�2Q����(����6^�Lx�1v��zQ���.z�ٷ|"8.�����-U�!릤��&h8Uő:P��)�,B����廐j}�ҹ���+i���=C�z���^6���VΗ�%��������3&�SmZ@}��f�@��N���@4��R5��(3��:�g_F|�=�D��_H��@�v	D��Ɓ�0���<w�=9�.z{�0�8����8�����kb��6�>�Hؚ%��e++�[��u"�t�C@�NE�x�����i��.�Ͻ�w*��n�o���\{���͛S�g$�����)=�}I�$ʹש<�����0fv��o7�X��v[�"�Z���:3+C$KoL�w�2wIE���v6��X��n��m���_��C�Kۖ�^Ki��V9/rbtb-R�޻�ڹ��5J��dӱ�t:uv������5S]�;Wg����
�����(ў�iI@�۵��^����<\��M�X]��ٗ��8;I�.���;4LW���F7�k�b3.�]����V�������Y@�V3��OJ˙��79�Ї��V����OC��}f�2��u(��xj�v�1F����<ӒG���v���B��ë�ٲ�n��Q5G�Gsx�o����KA�%���C{�c������pV�r�L�l��$��8zf�7�[�v��^Iga��<�	n#���_QF�b���Xolp���n1�q�Cg!�y�}�H�>͸���T��!�����uZ�m��
�]$#?";�'�ι'd���]�-���mSi2���k�h�O]y\V����L�4;��o`k���� �*����6�@P+��$��z	�s}mn��/&d4��J� ������m�jd��o2��F�$%�&��)�������1���`��9�.m�O9%Hn�r����{̀\3Njf����\j�]m@�6�WJ��L�I,gvrpX?Px>�`�*&�֐���v�:�AIL�I%M5m��
���:���D�������^�j*��(�
�F��V��,K�A�*�Gpb)&'�52PTKA����g����1^g�9���EAz�sg��1������&�&���ժ��&�b�i��&e�(*"��(�8�Ep؉*�����5U%��ͻ��DSQb(�y�$�ű1DQ�[b(����s&���ALE1Q+LSScj5����j��ш*��3Nڦ-�h"c�55M�P��F����cCq�*�*���QGP�)�\[i��uR�DSl���b��
%���:ƫ���h����Z�F�MEL\ڂ�����h*����-�V�"���������T4S1��*���*&� ��J|�\m�m����X9�$Aη!v�p�(*�	k�[G w��1���Q�Q.�E��B�gbmEͬUh�7}
�n�,*��\��Th��bǢ� ;*����_�-�җR��k�%{�B�R����-�c�A��}Ϭ�}��6f�N}긓�� $�/W�k��gRF	��6�^�u�\��+zuypc8�ȋ��n x�0�S"l��/�	��;2]��������p�P���|9��ν~�Wu��뽌j�s�[���Q�*N�bȜ�D������=y�_���o���d�dN�iR�����oկ����2���IP�U���ڋ��~��~I�7V�}^�P/�t�o�7�|o
%�@X���EPl�<6n!{�"ǓѣE�Z����<�*�2
����W>w�q��aQc�GŚp�������N,2�н�m;"��_ۚ}$iw��p�E��ќ�V��UV�o;�~�'Ut}ܖ�O���}�o�X���T���G�K��tU�YhB��/[��K^�3nSplc����%Z���W�����E�TY�?�X�]���}(Q���"�lZ�N�-z�� �/�S�a)�o�]J��M�w�Z��c�j�TdO};|��ԠdXښ��>�Uq�;���>�	��Z˕����>;+��G5��Tm�X"�wź8N��ب�;}����H6l���:݅�Wn7�[뇆o,��+�g�C�Efxx�״�N���/��m��}�"S��q�֍`�x�Ʀ�5�;�Ρ�����T��Զ
;d����'lM^D7��������$Y��"䱮{��D����d�	�`Hc�z�I3u0�9��T.�M�==��ܪ�(z]����f�&L#&��[PYA�5j�`?{��?����U9GB�ܸ���8����j�.�����R5��ڬ0������=0 �K5���ޚQ��v*v��;ف�L9;e\�������&�W�qAx��b�����~�H6,����1Sᔳ�8u�Л���A��G�V��ou�⼺�_^w,ǜ�q���!'YCwIғ&s6�ѻ!�,q�2�m
&X!�x8���?ۏ�G���r�����%�.�D*���E�b1b��bŬ7ˋ���X�X����[���ʻ��՝�}s��.�Fi��q�K]SZ�0�xC��|!���崡��FAg�Jǐ��5�������o��1�6E�Z�J��y�f���Ps�!u0�>jEG�������$��� a���g=T��ؗB��#Ҋ�kL>U��`J���e�h�zm������ãq�z����!kþ�*&�U�5ǫ�WS���򶣉�b��������3��G�p瑎�����y-����nf>�C�ۡ�:�]L���[�ria=s�^�Y�ӧZl��IF�j9B��l��-���	�������Y�_rwa��J�;��d��g������{<G�?7��h;���ܿ0(��k������j`5N�
�ܭM��Nӑ��������|�f����g"]��8<}�B�������o����O>p�Hp�����se�S�{-V�0f9���M��>��߾%a�4)�����䛠���pם�Z�2��	��ʿT5������<��lo`�~����3yTbL��C��B	���c�ؠ�΢6د+4�ן�Ojb���~�v�ƣ����=`?m����%���k� ��ܺꝫs0|�rg{�Z��*<e�ea��߰jЪפjN��هz��x��q�� �xq�)���=��1FA�AӃ��c��`סտH;�3�<��>���)֋0|};jm�}��:����Z&m�<+���R�v_���P`�o���w1z*6S9>~2�9�_q���C9��}^�D���K���u�y�_��^�h!b6WG���D�'퓸��6�azp���\+ag��ؕ=$V�T.��
�4�e@������N���u:���AN�9�m��,e��kxO�7"/����/�tc*��F��b�Z��cթ3��p������gm�m��Xh"{3m����/�'D{�o1�3�ӞNv䄜q����l�����޷\��~����6�=�i��1*�&��}�v�^�{�"��~��p3����b,���Z𭇆�f�gP%bA�w�K���e����׵�v#�9l���ZgcB�]9���/O�9!�XcY�X���Գ7��=��^l{�Ga� <T���f�=�f5��\z9:�WS�k�[�x�D���0�⬍��&;�I����)�Y@p�
(!R₩�/�[�m�t_K�g:�nų�c'S=,��uU]X�^����1�}g ď9�U���Wo�B�J�N���
=�h�������qt����;I��,����[@�jG�63��}�i#5}�2b�7Ъ;���d��j_��Bm[��>w�PWq��B��@��N@����1�.)�h�D4���(��U6��ymK��y�r`�W*"z`EǇ�I���}�ï^�.��%�(us�
/`��,s#�����ɍn}����["�19][�}�����,�r�@����*�t>��/��~��>�^��;W?/��2�݂gkޑ����|�r��ӏ���F�`4�n�D��\����b�
����dXV��2����� �y�VT�w�f7giI5%X���W7}¬�W/��U�=~�z(�Ņ�y���J�_a��'�y���9y��iA�\�j�)����v���	=�H����]�X[ �����!C����\k�Gl=���@����˕F�(q�F���\� i��\�*�c��A��`J�bO�:@2������>U1��ެ�N�E�YQ!�~c���w4�`w��F�ꮌ��Z"a_ʄD��M}� �a��I�*m`�竫�^�:�hDug�)?l*�Ԉ�E�*����EL+�����EzW�NPY5�W��s�#�ސgf�X�J��z�z�ڀ��-���A���{�< l}�7Rm�?��{(�[Hq���=���_�u�\����~G�ǞD^|�nol1�ڛ�]�Lu��N�Տ/SU�-��eK�)���鸝��������,>_]����UdX~����]lC���3��O�r"�[Bw�k���`\4ڰl���7�]�&BdH�_�|�W��)��o>����x"�	�)qѽQ>�g�bȽ���j�Bf�x�E����JF���(�a�T�p�U���޳ƅO*�S�_̖81;آ��p*����z�c�ڣ��1��e?a3C��f�b�	o��Q�c�����ue���d�øY��*����(^�p��ٍĴ1A`��]�p�i97������h�i�L�-� zC���kaj���9%ܻ,�P�SV-�t������}�-��\Y��YX3`>bu41�Cg�b�fPݩSL}��}���˖�8�&#]zg�E�/�٘3N[�3NO���X�b{h�l�K�ӵzs,m/73u��mDl_�U�,�!��W��n�����Uc���p��'����9�̊'����3���_Q�vW�%
q�;,�8<oъw�'s���.��~��5x�Z7�f��ۓ��Q�\����Ư U�bM��@V :1R|8��0�t!\��.w����Lk�^ތ�P���)ՙ��X~��2�Ps�&b����A�A\	&lTÒ��?KUٹ�(V���w�.`�6g67K��F�5kf���qέ����ISѐuNNe�J~��N���;*�|�k�.��t?N�o��S~?L�:'�8*`٨d��b#�w61��<{�݁�|]�Q诤�^7['���s�<�M�A��	�g��(���m8��zD�ux��F�R�y��"�C�Q�2����t��p��ҽ���pA�^9���X�X�:��D��N��Ĵ���I���x��)I���$�� ��o�sM��f�eq���VDZ�J�x3�3MdP:-��˗^�s�wݨba��۽Cw*�b�+''WѤ���q��˿j�FL�À��C/���V���`����M�����7轝��Z�����f�;wo%�n�Y�;�$��0=�c�6�i�m_i��Ԋ-v�R6��%��ʺ�_U%����c&��Nc�ԣ�-��c!E��k��вd �]��z]m�55y_Y��-��HS��)D���ҤD���8�߭���'�C��dk��?��%���˻Yf�p׹�N��XZ�g�8�z4.��~�p�3����m�T��hDy��Yۘ��(�{^��#Xע�J����c����o�������Ҫ�9hSv.�u��)Dyqm^S�>��s׋�u�:�&Ę��q�E�s���zm��2�S�V䱍�֙�p��%Ͻ����H_��0��쿫��@�z,
�ā}t�=5�pҮb��4����7[J��������u��i�t/���zǳ��/���`P�B�?0Ĩ�>�����"����e����h�ܔ+�%�}�u���G��T[�6;7�oQ�8*Dz���!Ίl�(}��UwQ�H�����`ţ�ĩ��Qc��X�G�?m�
�$�j'Ӳ'��;r��F�:`��*`u	���ܻ�r�Z�ZZ�Iڀ��f��/`W�`;� ��[��(;���A�Q>��tk�ov����^vS�3�Y��%�"E���_-w��ؾmT��x �f�A�z������P�O�D�
�%NR`j�gW��Y�{��I���ܽ�}�U�ͻkq�b�o,Zv�Ans��C�O+�X��&/	�������,���u'��𞏽p%��
L3tx���uo��>��%;n��vϷ/.Ozp�}
�OYygC�ȰN� 6'�4�X�S>��Qo����݁����'u�O
ƸaMWO�b�ʦ0�Fx�,A��D��= ��.�3�{�Ce�I��1�~�����g�'&�,��5ncw0}8
��=���!Eyf�B+��%<�S����&Mf�A�ݎf'}� �u�7լM��Bs��71axV��j�j�OP��\�{�l�6��յʻ`r�c)m�*�sNGi�<�[����m�A�~��ʲ�`L\���,_�LK�۫�h��~u��􂒫��`���N�FG���>���<{b���\���vc�'��O�3*�(�7YRpudM}�Q���t��t,�g�}�]A�4Ÿ��]�{���Axf2'q�$E���.������F��W�rO����^X���e~�0v}8��X�]ȶ_����U{�xUXj3P:��p_�*s
��Y�(��CF���W�T�~��k���#�6�Wj�$V�V�A�ku�'��=?X����E���;�c(nv���M�Daή�_` D.����J��Kq��Q������[��#�̄ђ�5v�wv`�O`�2�+;��a�e�ʟ,ӷŗnK���`7o��,K$B|}�|;�Y�̝=���]��n�8?x����9~SWK��5����	5��+��U�ipy���qw�L¥z߹�c�NS��GH^+�<�ɮSl��<���
������K%X��;ٵ���h���G�_D,���=Q,R��,(X<���cb�n��79��ɍ�P�ω�y�3���*�Ӊ��cji� ސq�����_�Ԡ@6��#t$�\�&UǷ��Q���%��X��xu1y,yP�&2lEh=BE1F�
���K�8;/#��gl=v��/hL�b��8��	�쵦_��Jv�@ƭG��Q���*±$lM�EL�q�;���]�Oý.)W���_Y��G'�Ԉ��_�a��ʴD�R",p�gD�I�o���_���0�,���!��-��Q�k�R��N���S�����˅d(â��W3����9���4D=��$�B���>����`$�B^��s��lN�,raG_rW�}.!y���Z�T伒�MA�4WEņ=N,e��s��oN�q����"*Ǖ8�V��:c!Xg�D81�3Z�:����R7)T���C�z��9�w�7��3m��ZR��s��� yQW;/$�t�W�٪ŬE�t�n�jx��j��usS<;��9ي���v^��2���.=���M�D��<���=u�m���5O;��]������+Ԯ;�%q%lȗ���)�����ř�S�����6�a��x��U�o��Gi^J�B�6�E���H��?��P=��`��L�7�]��d�"���z�E;����u��	�4�QW��5:=��gf=��b`���xo�=���񱄩�9
�P���b��8��c�K#K�X�V���$�F���~m^C��c�ڣ�����k�8N>�Q}���M1��t��6f���] �-�Xb��mN}&�Ksભ����CϛX�cEw��VO���wD����;Z�N1���#"��D+�D?*�����M���?*�r����y�?b����޾�r,�Y��S�}_I��(0�}R�8���ȃ�7��+�T�S�S.ߪ�Vw�d�ѳw+���s�C�T�55y��lI��
�F,	>Fɘ|Ur��A=�ۉ��f&S{��]��>�wL�n���{��m�V�ZQ���z~!w(?.�D�����\^a�Q��&�w�+
�"�_�ב��M�B~�Y�|��]�B�6~D�m�"�ѾD�F�χ��^�c��~�<���\m;��t�3��VL�X�4�����N�b��9��=�}�flR�{-'�(��nd���,X�Cm��Fnxl��n� �`OcYF�󗦄s��ԍ�me[<,�wM��]��;�qs�U�^�E���%с}���u�ki{��!�K����뇦
�<vs�ܪ�����#N�%��}�����yX �lA��j�L����8���v���ŵ=d�� %Y>���9\��Ұ}!���E���t)b����u�8�T�;�E��{tnxzO����0 #w��
����:d{^��o/hú<�M�7����ˏW}����7Ts;^���1g�N�О{y���˂�]�<3�]��ȆY���Us(���wI�Y"e�8}:^�W�i	�/�ń�6����nLl�ᙆ+����z��ױp��S��^��侷U�i?��r0!��w��{�2'U0�`�Ar�2mγ	�g$mA����*�C������w��g9�[׋q	K{z��y��i�K�B-�h��:���h���
���<��z��gcZ�F-]v>��h�[��Pa"��d3�f��8I��+��NS�'��N�V�J��!l��r��M��*^ou���6!���50��X76��,^>v�.w}TV<W����g����*���K�������{ុ9xb]���O$�:���o/�%�vqWn�p�k��iRU�ck,l�/W^n��t��s��Ͻǅ�O���m1�G��C�����||z��y~��r�(ho���7��S��=�&_giV�l�`θ����6U|���pls�������)M����C5���9�qH>�6�����t6���+
�5�Y�d�0�}�!����5�o\�$Ia���.⸫���1=iu]q��͙u-
��~}�R1(�MG/u^ �F���6��_M윎S��B*��e��v40�ݬR1[g%��nʄF�<�xoI"����g�٥�<8�r������<u-�:���AP�N��˼T���p)CkS�ߦ��V�P�8�R�U��մQ�:q̑�+e��]m�c��׮�x�U�I�l ����uR�@�W^엔':���b��C����w��J`j�:�mM�R�`�����y\���v;= pf�CC7�,�_d��Ugg�b���9T)�n>|z�5c^�'Y0�g�X{�{|\�U����r�IZrp����g�dP���үsZ��{79�;���r0 *G�*�iB�m�aM�ۛ1=�9�6�� p
^y9��(�����m�/Z6k�����5��gu�%o]���ħ^v+1%	�٫yKd�kA�7sz벂Oh�W���ٻ�J
U�m�]e޳.�X��җV�nظq���9����٧u� Iw<�ڙ�ڵ�t�έ��mT���I$��ɐ���;v|+c�71��΢�o����!�Ո���TSh�
("
��h�"���A�#�������<�*�F��=lUP\�EQD]m�f"�/X�D�UQG1=�	<���TEͩ"g�s:6��� ���:�
�h�b���(��EA͊��N����b(��:���**(��)	�EUUU4y�w�Rw��4��W|�
"*�
4h ����Rne�;�]r��4��5Lw�4��ד�+n�]j1[-��)���梨��93��ة��UL5��W{�0r��5��k��9G#A���u<ƪ���P�
9�4G�M�M/#i�r�[�j��B�
�\5:���4D�4�9��&xF*�:(4��q���h���\���ʎ���4�E�؉h)��/	٬����Pj�9�l<*9U=u�����+�$�?cS�޷z�l�y���7�w�wBJ(�9�;� ��<=<���}y���;��������8��]�G�	�C-���I�����z��nK^Ρ�������?�*�X5�p}
��@H��Ԧ�w�N���	1�ɂ�i9�s����tp�p!����N:,T�񜾩S����G�ې��� 4��sf-9ك�	�l�޷�r�1���Ӏ����`�b}%O��h�vG���8 ͏/q��9��Nͪ����{���}ב����!>��ʹKM�Тd1bEE=���e��Q�|���њU�;ެܥ��|�z��8���S<�Cc���aQ�܎��}chY(x��Ĩ*r���F�c�ǥ!����)C7�ǚU�z�0/S����~�l�<"��l���
y���s��ݓ�EM��^�?}�u{S�Qy��0�t��?P�X�Ήϕ�G�=��|��w�ˉ��E�Vӈ��P�CD�>�ȹ�b�*���ʗ��e�h���/�ض�b��;V�z����r%�>�2����!��9%��*�����u�Kfͨ��N:/�\6s�4ϰB���E}��5�����4�c�3'i@�n)xߣ�O�EKbE�:�x4�BiV�X���㯤�z��i�Cn��(<u�������}�����ʏ^�8fMS����X�i	ٚa��O�z�:�GpTh�Q��5�=�Ζ`��C8��`�U��=�q�����R����nt���f	ƊZ(W�I����_1�ʟ]��&d�����W�w�W�6�1#�!�,���hJ��f}�P/��SW��JN�R�%|�s�^<�������LLk-옱�L�|9�C�k����c�WƉ�<W������l�Af�$�����od���,p1z���������P�5�ȃ��'q,G+���ם�~��#>!lu�T38r�˥�1wҭzF�O�l½{��S�'�֨4�.��e�-��wf�_���@.='Dz�^�18���e��B6�S��!�m���Wl�]U�ed4#�]���x)��XK��_�?į��(�{c'콞#J�o���{��]�Vu�;3쵾�6�c;˅��qN��j�̐�N}
��ߤתa�ze4���5Hj�\ǹ�	8�`N�L`*��
����V�ϺFA�4K"l}�W������fgH��y��sTv�ʍ�ڏ�1�q���+bp:E�Y��^������@��R��%�����o�+�_���! �J�ʻ�ӑ�����l��o$1���E���.8��S�4J�T硎1��N��>�돽_�1z����!��w�i��F���~{&���d� _	�|��ț9��|,��Y��~��N���@�0&���9@8��n�zf����"�o�7;�5���θsvc��U�?Dk m� ,yl��}|4w��|��k*���}R��Ț�]�$�+��j��nٍ[�ˍ��rvN���<֬_�8�k�gy��mwzc�� ��뎚�P�����֊~3c��}6<��:8�.3��Θ榠Aބ��&"��~�ߞ?�}�ݳ/��r�b&~�;0y	�`hz�m�������"b�v��UE��C����3V�hJ�ӡ{𝤍��Q�r(P!�a�S�F{I^�^d�����p�𯎶3C����7m��SWK��Y	�n�Zd`�ږo�aN�l��4�Z���^�.#ɀ���)^B�>^�R}6��.�C������u�O���or_\�XW�+�Z����4�Aab�̝0>�WT>�1{/+s"���s��\���(O�֍�y���(��y��g��T�`�6(�?=��t]];/������^��;W6%�	���U�k���O����7��
�)�@�	I��A��C�;�y�\>]D�I̧g��Vg0��o5���:�%;s����T�	^
���4%�*v�:Z�_�ry�аwV�ޝ}�F�����isX3Z��э��P�m�J����ϭ<<��̳��/~�Ei�y�����K���W�iP='h�2E��J������$m�������:nԏ�W&63z�f�Ĵ:V\r�E+���l}�r�9k���  DG� |��d�1��8���*�?��p�tr|]}[((��_.ۈY�0�j�_�O7�]eT6=�'4��{��q��]M��*��u���MI"}hN����.�����+gtTi=��ة�-�${�Z N��Ӭ�9���ث :/�r�6ؐ�s�0��^ڳ�<MHdl�5~�9nG�ٛ���b\TPaO���!��s�s��pcyy����4S�j5/g�닗��Te�A�L�k6���ư�lL���?��e�eT�9P�Ϯc?%~W���U������7���3hC�t�z-�+ԍ�̀��c�Y3�dH�_�J��n��=��gf8ޞ��;��1�q���bf�w����B��o�a��WF�m��acrԇ0���①�a���0����7j�a�;>��ؗ3�|�Q�[�p�!�+gfg#�~ľ9���"r����L���6���jܷ>
�ܭ������q�G�HT���{���_��յ/��������w]�� ;��E�N<n|���u��g�8������_L�Ge;5n���=}�W�~��9D�x^�wZ�{/���|���vz[�X���,�r����y����6�W�h�i�'�ɪ�@N����}���F���5���k�����7áY�:�Q�t�ݩ��!��\�� �>����V��T��n�׎�~���w�pO�<���\#�NEx��u�X��Z�����eq���1��6��礦!�Jy��O�^@�hI��^�����AH񚆤���
��Dp��T#4�O�TI�;�������CЪXn��e�>Ϝ�1>��#� �5����2% k�e�j�c�+��ǰS�B�j�����ƳG&����e�{�[3�6`P)�`������x|5�������cҌ�9Pg�+̻pU��:�����l��C��s�S���&��qRZn�}�UH�K���|g��\����`������j�МX\=GD���&���/x�ڟzȱ�b��$O�f��a}5-`����wX�4���a�J�_�&��{�ǲ{�ra�s
���'<o�a�l�' �$ThG�}ut��]J;�i��(Ӵ�tw�8��D�D^������`-\���5�R��~�),A�������>�\/幙u����,���6���՝�� �K��U�ߩA���;�H�,�%ߊ��9�̩ÐfnYނ-vUm�U�}�{xX�'���p�2���0j�q����ΣܳJ�ֳ�$��(Tg{��T*�|pu�q^����ou�W->Y�ڳ�W�>y�8~~�%�M�U���ք�s�����և��v��~�!(�����辽�_1�����*m]wN�>���՞���0�WSs��g:>�
�ϣՉ�Q�]4����A-�z�{'�DC��Y�h�^1�r��*_%�xtw��i��,{0�M%EyFԜ�/7�Tz���i�h�z*��t���/���g����/ =���8迺e�g7t�zb�ި~C7�6W8����=��<�̌��P+�S�/�G�P�l2|!�uDxFV&��ɸ#�\V��:���ǰ��U���S���{'Լl��`W��a�QR|������\��,�5��;����X["���먰}����]�5/�B�b��6;�3x&z ����'�5�7���q��!-L���r���k�1y[�ezٛ�yMM��Bƻ*���'!ʞ������1G!NK�F=�@�ꂄ���+E�`�
����$�@��مz�:sF�BUy��ru�Wdw��ӝ��8A��"K����(:p��1�<Vz%�􃰍�����=e��"|n4�e��C�H�ϙ�f1N��j�	"��c��}B|�`Ό���g�d�~����p����s�ܝ�:��}F5�{�ќ
�%��y�-ƤZo�j]Y�s,<�~ּ���g���Ip(�����қ,�2/��
�%CV/�J���մ�����0��
<�TE����2yH[����w������^�{�{����׿���
�}��w��2ɾ�c�A7����pLrwP����p:"U�b�h�Bhp��gp��B^�eD{�DzVa{�q��ۘ6<��|
�S
����U�B�9ȸ><4�2ǤU[P�v:�0��V��-�����&��Ք�Z8�<^������b,�s𭇆�f�{q�B,ێ���[����b!�B��e%{⾻�ӑ�|���5�,3m�`-gѵ��gc���B��ڿQD�m���c�9'�:n�.����R���ws�~�S��#��G��w-��O����<�^��zA��� W�+���d�����T��5��y�m�tq��ٵp("�w��/l/G0���v-�S�c3�[��F��W�r1��O��$60�����ގ:Ԕ#u�Dg��9(
q�3L�n��~t/D�$oN�,�L�D4{{���=Y���k�r=���8��xt�@�*���娚���5��o��G�9�,��i}�N�g�[ׄ�-��<��XJrnP��y�/c�����^[R��x�ɂ��6}�S�6I�φn[K���u�Xkn�6�9A�%��wކW{I>�������x�����*U�;�a����/h���<V�Z�^ܼ�����V\�ih�Ҡ�2z���z�f�,����ڻX��<B9��T�۫[���γ�\��}���?�%H��W����6v���� !�9�QTE88�/`žX�Fb��s��\�J�;�g���Fm�'΢�����1L.���0B����\��'��@Q�y/`�2w=K.kyyO�{�vM��ַWI�7W�cʇ���k+�(�W ��"_I����7��𛷖������6g= �O��IN��5j1�n ⭁)P�A�4��;!���Pn]ҡqњab��ݎ$�j�#t�?^��I����]�~�������0���j���<��S���%��7Sn|�@��j{�DvFyB��	�TP>«>�²^)��Nl����l�Ufc��&@�z�S"���՞3�4��B
�ݞ��K�[ؐ��
7�U>ܯ7Z��T�����2~`�eJ�=Wĸ�cң�]l7:>9[ӫ�pc�;���[�O�eV﵅U���V</��� �����)i���>0χ��OR��S��V��qK8�Y�.`�C	%����v1ҁ��mm&o�o�BɔȜ����/)��?,��m%O��I����ʺ�s;>6c�n�H1q�7���r����~�p�-WayS.�a��R1ά��P�3��s���J9OI��9ۚ����|+ou���%79Qf��[4�����vβ�\����ø�49�yR�	+���ʯ��A�H$B*��{�������ߛ����������V��ϯ���S�}��9��ߠ.Uj����Zď�+ҁ�������5��
FF��&�b.�"pu�0W�Ϥ�F��߃j���n�Tv}6����d�f0Zž���g#	
?8�5�!	.C8P𯳫�l��-������BẺ��s�Q�Ud<��������(���t�f"��._�5��U�Su�7\#���*rE�v���AW5�yd�	^���;=8m1������)�>�������+�B\v��ȃ���1K��IM}>�B�a��]Gzz=S�qO �>F(sj�Z6$؁^��@tb�P2,����n�1��u���yO�����t:I�2��;�U�1_�49OnT.T�Ǹs���T�Kx`�+mX�YIf����'��Ǖ�wQ
���2����1�F��ޓ��C� v�_����>Ç*��c]�*�~��$o��Xc�ؒ�ʌ��>�Mq5���	��`��}P!�Q6�
.���r���`++nBP����ķ*�:�f���*�f�Û��;6h��L�u��^�{^~a�|F;�]O�`�T��r�!�j�\�j���#���g�m������=�;f�ǳ�$W�����fN�K�
a��'G$���[�+2W��q!�n2Pq�x^�7�n�F�.u#�&�s��|����	A�AW�￿�����{��r��f���6T(�24�D��p���E�WOҴvX�oI�ob�|�ϱ�O�jw�ÎM�oc;��N�Xj�H��V��7�KX��bEEF//-�iH�Sl�q��!;�cﺾo��E�fw�bU1���z+&�c&|��9�����f����oyWb��\�l/M^W�Y�Όu6�P�Ղ`oքc~�l�=
FAgKI۹뽯2=1=�v����D�#�D�46�t����x+f�oQ��,35"����^����c��LOZ�s#r���}�VԜ����>�5��s蹿�ʶ_ҥ��c�X�� *����(�ƴ7�bw��"+��;�'�����v׭aX���~��~5-���j#�r�9n�����MLٶ���K�H�����~�~da����K�����	�0�#��CU���������h�\G��#��nb��?C��61KeXJ��O�&}�P,p�
1*"k�]��^����{}{n�:�WCG^�Q����r�l�s�>-|#�(Aƿ}���s�SC|W- +�O=JVW�Y���-�'��JVj�e� q|���t��'xV4O��ɛ�a1K	�r�-�OjF��?���e��\H��w\�:�=��j;̓X��oۂ>V*Y�2)��:��i�MEqM�8�t��Z���	��t�΢n��&_:���`B�XH>���w�+�%����d�R�[�C/&ܻ9�l�N�L0��`��`���5ُ�9;������#�PA!��;z-Q�Pn &��������F�̙n����m\�!ղ�9�����NfG�� Í)��(��y]rͧB���M��V3�I�÷#��D�F�t[`֊<�'��nS���x���/_mx���`ɝÑ3y�o1��]ՎE�A8�d���+�.L����A)uyL�j���pɀӲk����� �5y��+cV�.���v�j�������G�3u�v���`��[��;�[�ӃD�3��Y�QpD�zK��0�LN1�g���n���칧�Z.�{wY@}� �WTy�����8�]%�c_�ǜ(-�[���.�x�c��%Q�Zf��J�z���"*��ڽ=��!��������6��A����Ą���������«�+�[7e�:���Kn2^[��w(��$�̨�����{�%��J�� �˝�������<r<��/-ݾ5�c�/��{ T�gT�!=oޤojhz^O�:k�(�*���ϐ�}�7��R\�/6��sP�={�U�+�6{�9>��fzE5<=(���K|8멐�5]�x�;O:��Ca������G��	7Cț9�����s�l�qX�^�p�x���0dX�%�J�`��*D�߮Q���'%�Xd�vA�wk"�bJm�8��8��f�&Wk��]+�W���T1vh��q�o��s�W��{�f�*
���/�i��<R�([[2-�9MNH��R`����n�rg���N�w�c^�ŭ���r���	R�x8n��p���Q��L��F\(u����P�nRD�Û�z�7��k,��p:5�Q8���.�Z���B�vv*3�6N턳��t����C�O�<���{	"�=��h^���ۉxޔek�o��tdkVs��]�\�seq��*���osZ������:�\r�x%�oj����g&�/�l��ƑHe)�F7��tmg��s[�]��qL�G=t�ٻD ��Y6�����-}�ţ����g��{7${|��7+޾ܺ;�A��Xe����é0�C��Nf�*m�yu�ǔp������]��:�dGf��{y���HM\)dRFl�(}ԇ%�Å��V��}��� 0e�Ov,�z���2���Oi��Lӊ����p@ۇ�a�����p�5�[yp��8��}r�p���??i�x����g��/PFl�}�7��AΕ�����|v�!�5[��R۾�z����V�_s��������%�s��I*�ϝw��_>}�肝:�)&
�����C�.z�W*��'|1\�w��˚�kG���䞠�^�6}CԇT@UA������͵��4��G]��[z�zẎ�8z;<;<<!�)
#͊�� *��#�w��<�<�2�S�cn����OXE�3�W:�(��"��P\Ω.d����*{ƪ"���p��0�Pփ�l^d���WVឱ��T�؉��Np��s�J<�C� 4h�-��,m�|�v,X�m�f� Ӽﮀ� �i�3-�+Q3%11-Q01�1s�bH�cTy����|9�R�嵊{����i�	wb뛕�i�P��E�����IS\�'�%<��xSxt�����S�ː�w������z�25E4�ˠ����|���\��ܚ��ש�SՈ#�f��:��ݣ�*$�b�|�V���I���(��ג����x64v2�����N�(�<����{�l���n#z�~��:=x#��l�U'6�����]��u����� ���
�}�����C�z�P���ڕ�Z�[�g����f����7j�*��ӡ�(�p���M{I�`gIF��Ё.�I��/�����*פn��(5�8af=n�R2�+�.�b9T����}]�x��Y��.|��H�/����}�X1�<V{.ߤ(/G�#"���������k5���{�a�*v4[��c:/�yXK�0B�����s��ڄ���|v"b"W{ov���9��tB8��@_����'s��B��1�
tD�V.f�
��_p��WQ���\�{6�Y<�.�sn�;��������P0��0U#ַ�#0{C��B���Q$�;}�^�b9�{��'��a�$_,"�˘~���ըM�		nC_T��9�EQC;���_���1���j<��D��a��E�����4�gݲ���e�j/�)a��)y��yZ�[�3�<w*F�TO_��2^꜓�j
�7��
�����շ�w;>��>�6�I�Wv��b/H��?�����Ȝ�{�Tܟ^���%$��<cu��vTc\��b��o�D���+hEd�;�:_{������\-�;G���r�$^��AC����k(�ɶ�������rM뎝�&����lkX��R�h������ٜr��v��:?A/_~��^�&˻f�d�e�|�q��|뾻������e�|��x�G� A���>|;�{ؒu3��d ��1�Xp�cv-��X�t�r*����1,zr)�^dewK!�h-��x��c9�A����^Tc��n������@q����𝤍�:��c
'[�{�캘�tZpxx�4��RP��.�sH�ƕ{��r�MCR؃Y	�n�Zd`^�Oݒ�e;��oz���H��D�b6���FM���X����E`5X��.�o�5��A��k��+wj�_u�r��?�K���H7��1
�]���Z<�̌^vnL�o2&�����;Ǎ��8n����u�z-�D��	��q�`Q�p��/m_�(��~��x�M{�����k�+�rL�Cg�3�NȚ �	I��3�~���O��L�j�|�jCK��w��ak����ft'IN���6��+�&�l	V�@��y���vVãq|�yY�f2\�G�f�#�9�oa襡��t�y:��x���b��*�	�t�J��'r|E���b!� ��/MI�Wۘ��n�[Rw�U��%D��U�a��j��x!�q���$p��#)^�:�����_�ö/]J�g�e9Ւ�@U�i�=�0U�r/�<����3!�׾�(e���>��r�A�1�R�9��~���a��|uz>ѫ�Y쒸h���k/5_�ɋ���^g>�VQ[_���J����w�׿������`VX��<�=�����?��1�g�bӬ���Z[^����P��
0�w15��A�G���0<k&p��z�*^z�&�����(��[Μ�����+M�u/dv�zo�s��qٳ7�߹׉6m�8���i�20OEE��R��[�0ł�ǷŌ���`�����K��.�!��~����'���6��c�Y2##;��%�R���<i��X����Q��Z����,S�!� 5��:�g6}��4��}1�sK�M�v�#ۍ���:��*�J �>>�ey��M0�aUp��j��n1[�qo����$���Xga��ؗ0
V��w?7>D��#��	}=ʄ��-ϾUV�Z��]�:��N酶y�c"�ɻq��N�貧$����������\�vQ�T@h�u#�]/ՑH���74�g=�*�4���-�����:0%^S�}_OX�[�b��%�oe���l�QSk#*���Y�⮢ƺpjp�\��v�k�l�fL
�lI��� 9��vg�ci8P�"�2f��]<���r�{�����3�zp�����k5N�շ	�~4�pw����[� �7~>��{;�(с�)��:�i�{9��|���ϐD�cL�A�r��-�UnVp{3H�z��(k3�[�ι��16�~����/|��;���?�(� }��1ը6�v=#��uq�4v�	N�_)|i㡰���q�Q*:�6Lq�0:W8Ү&EǞL�G�8�	�-�s0a��Z����͍߸�rc|խ������.#�~���v���&�������K
`A��?cK��8���t�
��Z7�h{�b]ȤFFӱ_�,O�>��/��/��
д�J_¤i������v}�HV�/w�#f���V��mmOY�,vw��a�\_�8	8������E	�h�����>��y���s�����bL�Ixc5;�1�u0�j�H��V��f�kհD��^�|U1��`�n޼���^7���Ǟ���ж_����q�r����#y��d(�W�>��dǳSb�G읡�T�_<���x]�5N�yIO���Y>���!�y>��R�.�����y`ɘ���5;kW)��=��6L��HT��5���^�olڋ��;��>jEG�/@�|H''������v���ڂԼ*!TܝC$Dx234U�q�X�4�C�+���Ʃ�~��������*D��� .�K�|+@�o
4=��!'NuKY}�m��� �^[hI�	G#�ڵ��y�9�v`����N-�0�����{�ݷ�^:��f��lǎ��Y��5�vˬ� ��=�������]^\}��g�FdW�?� ES׳���~�����{z������'�#[�P.[~�s�/�^��*>��?Bn��}�/Y=�ڽ��N��&zW˦P�3U*t*�r�v1���r7k�@��ND���G�C�TT���o7*�h���7;��	�<Ǻ���R���<p�P��7�)������NL�f�_V� �E<ƥq[�F�Q�
��$)*� ���pם�p>�ns~.���P1>3c��3a�=�v��-�+}�_`�2�|Z_�}� ׁ�Xr�J߭{-�����:�ڛߛ�
���c��7O�VLv���@�L�C[%��z:���w����/+��(T�FrO
��N���xG��R�<�;�76���T�+A=@��t�~"z]N�vx��ǰ��Up(:��n3ȩ�	Z�NR��rL�X�|h%�`�8?��5q@��ޚ�dQul��"wu+��H��ת�E�۱�o=+���v|�\(σ45ʌ+�+2B�%��[��������[���r��e�/x������@�s�w0�p'wQ>���ϑ~�����6-cv�N�����	W]�`�s�j���v��v���D͔{����mu�M��HT�:@��˴�̻�.�׌Ժ:[l�k$�LX��tW�YL�W�͑�-���Y�O�^�׭o(���N�~Cgw>�8�e6�����뿟=������Ĩ����_9��n�~'�r)�Ri�f�C��7ըM��a!8��X,���5���@֝8�N�a3W�Q��<��爡t��U�朎���[���͊`��o�4ۉ��z��4�(`����+E�NI����X�["����}k�Y\�X�|W,�=K���G~�4絏t��o�b�vzD�����YR�f��T�(*�\bq�ŽW���ľ1Hn��=��̸Q�IB�{J��浃�}�w�o�s�Nl�X;)��ߏ��\3�ء�V�z{i�@ۊ��g���~":P~��Tչzݨ0SO�V��{f���~�9���\Y援ǖ4M��'�
���3��
�>�8ݷ/�M\5,�M�P#�U��7��LS��oo2�l����9�'����#�*�gR��!b�/c�>�r�w�忼^�ħ�d�T
��9~]s��z#^E��&K%FL�鯄��vDz.���}���b�,s#+��΢Iˆc4�5-q��׷/�kzTkt�`����5�ڂ�!��_3�����^_,�s��j�X?4�ˈ�=�V����Ǖ*�Ec:̧Y�͔1VK��s(�W��o['̥�u��~Ĺ��%��4l�2���J�̾�e5�Wl&��Mk�Ï��{{�>�亂�3b�,.;�`J�M"���
��[o�|��~�� � Ă��Ͻ�v�n�~<���3�o�k�e^��L�~��Td��P�LQ����8��N�
^�f��:zK��e���8�z)��(��ߓ��nw��QN@�j���r� ����z�W���;��/�<�$�=���lf��O���C������8Uٌ���HD�J+(�o<��w����`�>�%`�������i�'>�X���M�'D*�МE�b����
�zѕ��z��S���|�����&X>�����U㵲�����4!3cn�Fs20L����9G�S��:�X+�A���S�g�ꬩ9��6�(����迲�a��r��Q��2��2wFꨧތ\bO��CI���z���``�S"sՎI�٨��n��xZ���`t�8(i�r��^-�_wu�i���VB�7q���C���E�ߕ�am&m�.�P�`g��[
0���q:(|�C�%M�����)_@m�Ϭqb�{AV�8�n�˳[}ӈ�p�%t�2S���'m�3���3�HT���b*�`�����)��I������cW�ǔl/{�`�u��t������p�H����<}�1�PT_F���dʻ�/�v�A��u}<w_���=�ى?U�ųN�*+��6�4q�lM�5�`��j�Kx��_D��,�fig޽}l���J���dD��&w%ԭ����A<��|��
��Ģ�����|�z���﮷����?7��5�����PP����"r�����E�/M�8$չnp�
�=��0�{�Gj�N��p_ͬq��޳>�����Ly�����;[S�_<�$}wg���F	
�í�QG���3���8T�*�g�GP�`=���~��G�@��,0�5��:��i~U��w�[���͙>5P�S�S���%��v���j���z�T�s��Y�D�0��䮃�%�b���i��5>�yB����[���_��q�Q*:ǦɊ����˲n ��vUW��O[0`<#*zlT��2�Z����K67�7=��oo��o���wb{��Q߷�9,��(���9�D���p\x�^�����u3�|U�d:� �*�}5����`v��<��B	x�7��88'�0L���&&��
,T�yMt˞�V
;:I�f����>�^M�9#�y��u�09"�Ƽ�$8��.(����?�{��,�T�����(���b�m����_/^��'�;�0�L8���@\+T��of��rd0DƉ�i�nzOe�#�VL�˼H��w�4mc���ցb��N�%ɍ&�z^�%>ʙ���tN�6U�3�7��K�G�7S�����?[R���d�&�0�W���E(ǡ	>p��vg�����QxXkκ0��K���8��^���x_�>��;��*��@'�߿|�����{����~�¤\s�h�~��|k���VD_*F`�~�#W1cgѮLVM.��J��z�_.U��5�kM"Z�MNVF�Wy__`�Q=���,C��^ߧ ���Ea{�K����,Ս�Sfrg�(O����t�5��lڍ��*;�,3²�/��oǪ��ٳ�#q��o}{�x+�����Iw�"�9�!WE�leb��4�C��fd:�U���	&���lq�z{�4f��FAM���b��(��`9[R�k�5b�|�TF���	;3&Byj�wN��w����!� �7�5J�UV��o���x���6�W)ȗu(���Q�"�c[�(�^�+�W�gI:�D�6��;��"4���x���4'��S���-�~S�L�f��s�b:�8���N�|c�0�!*(I�r����T.��M�Y�`$X� �yA��3z;�~w�s77�R{�m�"�d��Ć��X�gV)T�Ů�����#^�Szw�~�.�g�������b�Ƿ0+�d���%�p@>�2>��a����V�V�#s�Λ�n�P*��:gB? ﳍ���y�ق����`���08	�*__���bo�v�I�����FMc���ٮ��\��6�J��K6QM�����yGr���Ksr�b����i�n�q,/uù��GYՂ���[N�;y�|�|���ؠ~ D
�yף�<������"����ɳ
���/�tOF gdM}� D�'��	�1b����s�IY�&�-r��]W�]0A�cTz�ds�m��N���r���f1N��*$_D6z=�|��7��`���}��i�u��j���x�7����c9;�Q��������}�]�s��l���N�bX�^�+eo��9�&������sӟwQ��¶�cי�U;x:�*y�쉛c �Y�gGH����)�{~��ND
�V�7ƂBKt�ڼ�Kc'\k���1=�a�B�Ma�w�Ȉ(9LK	ȱ��i����l�v�� �[�'ԸQ�޸��v�s
�SA���o޿����./��.�M������EJcw7w=鮟EK�*��!癜=�c��:J��к�����+��{P\7�� ��V��S��0JQ��MU�Txz?*��^+'Ć3�p�u�(�H[�A�_kx1��>̷?y��i�����?w_�⿿�/�o�]l���=��-	B�"��L뮈�)�U�/~n�ӱ��u����@yEן��Z�n}�g�r�5��p�;$��*�z3ږ��׷�導G/��P��2x��Hė���-3˶w����fL�S�����_>��%�����㆘��Hu����U�w�x|}��k{ �}�G�ky��A�ɛ�����D$���{�
o��n��֗{�+E�v���wL�;$�.�>L�C�xMM�1{��K�F��{�>�2u�I��ή���w=�=������j�{Gk�M� �I����=���
`�"����V���xl=U�^Y_��4eؔ���n
�=J)z�F'����/��v�y̙[��Z��8S����N�����p���X}�U{x��^�U S�]ـ����۳1�m��"c5�y-v�v����r�U�a42'�u�d*����{���Q�b�#��޼U]���6n�&��|=�hï���TXlO]��McB�^sd-����6��8y/Dx\��Ŵp&=����6�]����K�W�Υ|�;Sz�m�wZ馟R�ŭ2����٭Y��=;��N�=����m��Ⱦ��E�+M�u��7�彃��0�}�]*�^LQ�M�������{D״wSz�'���x����V-�D�t�EȾ�Y� �q\��������.3БT���l0�N(Z�H��[\&�!�I��}�3rQ�X1���A��e���&u<�Ѿ8k�ǑbwQ���Mz(�O�e�芘G7�Ĭ�:V��`*�Oq;}G1��<�ǂ+Hqeaŭb%�5{d&�]}wc��zɏ#���gD���9 N�Pu�����X�b	_��śڪp�p1��f�{�]�`=�a��K���7��}s˄������> �U"��ܾ֬7���$���^�4EKv��jfV̏m"U%A1��a�Kȫ�36��,$`���c��:��D[�-u&c�{��wu�D��=sE�����!z�VV��������Fһ�骪
��t�gj�

�3fA�^Zv+�3t��-o	t��/V��g�	��C7���n[N����;tvl�1�'�'�/��4�.vŝ�#�������-_R�sx�����w�� W��xw��֯��|y+9�[�qT��Y�\��z�$�;n�L��nk��֬��V��+J�U�7����[��b�Տ���%b�5]�Z�r0��w�g*D&<�J��.ΐ^�%s��� Xo��ܐR
�<�n������d՝�⽿x�=�e����V
g�W=������d2�<FVn2�N�67�d�z��^OhefQ�����a��,jܖ�*���<����6-���-#/D;k�A�*uI,ռ�+zF2[�I��:�P�Q����]��;EotkI.��x��=Fc�<#����9�ܞ�Ǟ�d���g_^onᛅ�`�vž$}��̾��T��qЗ�"�aP����n�x�eIw�)$�J��s���OAU�H�!QE��� ����]&�ׯ��/�y�%LLX�i��)������c�����yy�u�Æ�:ئ���N��u/\0ΨJh"�����vF:<<<��
)�Oq�X�6i��*�
���w��QUuj!���ͤ���I�ƥ�FJ�(�u�rq-�#�P[5ALr��CI姛P�D]�QM!O
�tV�d��m͚�����z�u�u��8����-Lu���Ϯ�UJu6s1u*
6,h������{�4�N���H�F�n�E�qК}IÖ9�r�5�M��F#N��\�Q���"���Mbq��h�lm�\��qSz�r�SK�9��+I�9Um���֟#�RS\�F�#�b�*��]��\vɶ��r�r�EѧNب��Mm�AQG�w￿G׿^�y�9�<�N��n
S�-+��@!'Ҵ[���j�C����tM,,{���y��Gwፊ��^��G`�"�@��r�9~�!�B���믫��������?�}ܞ�:�z����`hx|��0��4���Ss�������%z�ㄹ&}L[���#��7M��B�f#�T�39��.,BE�t���VS��*�fE�b�.I����{�;˟8u�����d��Ӯ�l]�Q������՞��K����������u������ �Z��r�yљ��	 � ���������㾭������Sp�Mp��}V!��](�^�����s��W��8�CL❑4{�=�\z�1/_m�����
�X^A4mFC.�zm�NR��C��� �`J�1�9F�jŽ�S�?�c�$Oˍ����U{�ϗ��	C������®�l��ͿaC=P�d]���]qk��=@t����~5&��ۘg�m�/Ǉ��������O
a׳}��Ҕu �1��5�=����h�#�Dx��u�8+eimz�yp9��f9q�3s�C���2��`�͉W>�<ta��f��3�aB����ԧ/�F�ב���+��B�_1�X
����a�y�Y��F8�͆���%4o��h����k-P,v#���va��{�ư�`ޜ�v"����M��x_:]�1�P�d�*l��.���s�����P����Z���Q��b�Ft�a�}W����!_g��~��__z��}�w������ǞDZ�8�߰1��S"o��֫����N��vb�W����D��&wo��~���p�o�VE����Ͻ��;�@�Xo�����6�2����c�[3JU�����(�4��T��c~���鿸�N5�U�0n�΀�߲CA��Bueh���cr霗��3��L�:B@��U��[C�����|$�F U\7=ޓ�	�f���W'�7���"wE��÷j0������Bդ����"r��~�xA}=�ݜ�3�{���7���Np�X��qy��ö�n2��h*rK�8B��QR�6��3�IZ;xxmU�1���8�ٵ�!��,nT͹M���a�cU�*X�-�;!��|�tH�s��k/2�k�/;U!��ֈ�Ԣ�p{]Lg�����\���K+��p� U�lIl��3���9��=�0sC��H�1�(9��Jw�>��yߣ�������&O�}3�8���O�I�Gz�K�u�3*&��~��	�f�0��0a�J���,���mɍ�Z��ɣ��Ճ�e��f��AO�w�F����Vh�^����u����h�8W.�OUvD����=�}~y���)��?�y���&K
�U�H_Ct#U\3�2�f��]�g�LȞ�][��]�d�-��&�Rf ��Z;�������G�G�s�����'��}u������~�V\BS�1ë�,I�HISb�:Z�*��ksN�x|�Cѓ���'L·q����}{_S���~��$��̂�.?��֜�5����p��D:d��_t���&X��=��Z5y�N,.��b�d�Q�d5�qF����4%ݏ>�����W�Lک��O����X0V��&o��f��\�'sϼ���
��~�,��[I}U�uS Ԥ+��d�<,H��CЫbjJ��7�햆�}#z�*����,7J�~��F2�Uv��.G�=���L)N���#FȪJ�59Y�_]�}}��mG �Z_�R�8��xD��Z�oUn֣l��}�Pzڃ���5# ��ɑ��|��vg�r�����g�>�L9�.^�T���_8R�.���e��p��ߢx*;>��ڕ�"40�m�R�2�Lf��p���u��r#j����I��=3�9��6��݋xߠ\[�:�$��%A��R��Ҹ��A{�{�^���μc������q/R�S��UU�z���E;�#3�=J���*&�T}%��ҏ]/�V��0#K��v��[�Tz������t+$���rfc�\��]�sf�%ַ}׼l4�nˬ���cR���kc��"N�r���:�e<�g4�k��(�C���v�P�b7Xv����r\���e�n�w.h��y��=y���_=����P�$�P>�iD��^�!8�RP�a]��b/J���qǎ��p����s����R�)��iǖ�{qs��B�JJ���5��Т�E���9a9�B��^yQg�m�o:�~-�Ѧ����Z�㔶_z�e���>ڿ'��@��X!�'�;���9[��`��n��fd\샏�#V����4�n�=���==���L��iƩ(�v��L��m��s�~ǝ�Q���TǪ���/��rX�g���O�i�v��h'�|��B�1t8U���3�ŏ:���rX��yX���o���ө�S���hT7�|/aF	��B�E}~�He�Q^=��;�UC�>R�,���<q@1�ɼa���+N�3������r�JӴ�nWO���ϼ<:��pQ�%��^U1��7o�/b��_Z��U�IUU	z
�^q���E�OpO.�X��$3��F��D��T4J�&�P/���7ըM񠐞��i��O�^G���bD0-��SBr;�٘k�P�`�B�+l���
�9�/N}���F����װ-F��:�������j����/G�f�,>�O2�x]yOz�65�xSw���"�o*C�L��%���:��U^�ÜYN�M �ڵ�4�����鮹0l[,�6�9�j�4�v;4S�Ȝ�u�A��|��]`�n�9�����|������P=�����������W��q��B������l��n���PP>�b#Ғ��o �GV;a]���-�ju�Q���l��V1hO�9��{/ai������w�NZεo��w��yb_Ct,�`�}��\�$�n<U�jX�{�Ⱦ�E�������o8��;Q�<����t�|�X>vc$�n�5n^�j���|3m��^b;N��T��z��i�(<����Wկ~÷�B��d!Y�>��JW���0�]k��^�����)o���ӈ:�P5M��p���_�N3��!��o ^�S=�=9�la>F��V��DV:��?u�G�F�}@_����y�����A���N����cbive��o�MI�b���)�������\���B�v�Lc�r&�X[���:jw�t���n<�>(���	�/,ѯ�ߠ(�%�{�Jx�lc������qh���=����=�'K٬��m`S���gv��_8�a�n��F�Ir���ƭF�|�%f2���Ψ!F��ةO��*��;e�W�AZN����h�O:+���#UI<�~��wg g��3�x�gCS���b-�٩�N��et�ÃK�^��������$�������������O�臟���ۓK(o�ޒz=s��G������D�/ߞ}|���}�}��i�H�DC�,℘��I��PKz�5)ۏz�h�_R7�x�]fw��5Q�MC��n#��
¡$*_p�����<�@9Q�p{�Lu��ړuӳz��/�N��=�z�������QA{u�_�C���>��߂�B�!
��+�5��w,=~���C*�I��ҟ���s'��U6'��91aO��f�{ SPe��T0���R�`��~q>u�+����s��3�gyx��V�μH43k�5�b���D)~�Oh���^�t�q��t�(�KB9����"�Dr�b�]���؞�_������aw�d�ܷ����L��&���CD�6=~���W�B���X�*��kw�nm��kl�&Q�5Y:yuUu�P3���ΛQ>��M@j����7�hxX���K�溹gQj����'�%'�����y�~��g������JV����R~D� c���_<��[��f G��j�{������h�S�UnV��D6����z�`�ږg��������t�IV=��=�g}5V��Y
d�p��W�ݚ�"�Z m�[��0�ӗ��1�>�Z��x��C��H�-6c��T�b��B�E�n��Ω����2��0%��#YK�'P����j`�u��Vsc;g�!^&�l��gEB�j>ݺ�(�'�{���#�>��>�6���8�ǋ��T@��z�H�N<n|���~�A��a�b��^6T�v�N@�Br��Z����g>��$?��{ YdA��c�Ϊک����\��v�]��5y�m��WZ̈��z�u�����%@����xq�W����<�uu�7���u'���uE(k�N���yx}�S��KL�����AA�Ί�rV�0˥B�:���k����XݑF�_b�_/`�<�xusH�쯥��B��&#kf`PBJ���������Vh���[�&�EE�n}����0zt$o��Sf4.��N���̂�h\S��|cZs��q�;1J}�ٲ"���Gz3gXZ�R�<nB�j�МX]��(�䍗� ���
10{wR�y����{v��0S�b��KՖ:����/,q�����B\`�F�Z�Z��٤���4�\����Ǡ��*��"��:q`U�2���d�����Ց���ߡ��Z����;�=�i��{��[;n��謙��вPdM�ĨS���U����v��=-�8)b;�Nb}��#�Z�u��툴��K���A����pز�V�JJ����עtV�.����cf���/�]����ǭ_o��ޣI=��ß��}��9�}�*R�)�E��ݧ����&����͡��Ι&���.#o�*#\ۏ��hL�Ͼ	X�T����ݽ{���_z�߿��ϯ�yo�[J:�Y�o�*Kf�ڝӐ��l7��j*�A�5���c�S���=�
X~�p�7�ꏕ�G�r�xm���j\v�#+�婚q}1����}��"��tw�3��6�MЦ��!�}�0�T���)��]�4��*��c����vٿD[���,gTG
�NgƩ�s�*�r�v1�o��k`��o0�w�ϔu/f�^ױ�<+�T�$_�tD<n!Ҫc�q��4'�lb����,�&tNv�^�T�3}yv�N��aH�<%A�y}�C��פT;N�+�^�ro��p�[�ex�1����׃�b���ƃ���|h���dy	��L���U-�k�����r�����>ȯb+�vnGo�ކ�B/b#�H��q�S���sl|{ʀ9Xe��6Ey`�%�g7�\�:ǋ�k�7Co�l½s�_�N螌3�&�Ax-= !i�k����٫�Q��>[�藰_�����{��} �i�S�g!�n����c�*�T {�˻~���n�M��8�D�[��a�P3p�^�g`�̽�Ӈ�E�O)��CP^Xl���y��Xsѓ�K���?�O�KF���d����5��<d���;{��8], �1�X:۫���Y�S����)+��r�[4I�S�|��x����w�Ϝ���ȶ��$H�~��?Aa89�0Mx?�?`4���/��e�.χ���4r~���f�ҽ�w1������R�ܵxN߉٪բ&�Ax5�.�� �V�#'���0������~���{��nr�~3")ك)#��N�zb��D\/�4K"t�O�Ce�?{�:�߂�.��}�E)�;i��������@�5�Ma��숂�U�bs�W�I[e]�n��)��d=�/��L�[���:�=Ǵ����͆�/��謝���T�t�B}pȼ��|;�֎��ON�,��}����Q�E�\lgÓ��t.�!�~�I��x��ڛ�]7ՙѐ����+D/ɐ�6��
�WLh�}���pc>�Ÿ��a����c��{��V�2��:�|���y�a�;'GNE|ȯ���_r��"�']�)��5n^��@qh�������jsn{W:�8E��1ˤ����2͌(�<�IlO���9��(!{�_�nۗ�piUI����w�{Y��p���9��~��?��PWq��K��'h7�˧� �s�	����MB���VY�6�vT�ď�p+��Q�{c�}�	m�A���ߵɰ`���t�GXJ�r��t>�j��Ԙ�o� ��ή3����&>�� р�<"�<U-���A|v��j��L6��8r��R��[2�s���;�tE¹?�}_ʿ������pf��$FsU?�k��5-��'�c���>�$F� �KbW��\r�ZdΗA}w��1z��kU����"�y��8��҅������'�Oh�_�S�s�'�υ>����B�+�8x����j�Fy/`�I�����z�&p?P�Nȓֳ{\z��UA�bC�]� :�.��v^G=qF�ߩ����o�S��nw�j�B[�9 �r�ՙ;�w1[d���\�N@���c�OxԘ��I��P�Րϝ8���YT��*=�����Vw�'Ë#4�fn���B��DL%"#
��jo��w����P��dZ����NV�b4��#[%�=*������Y��7
<tTǧ�q/��4,�>���b�z���PZ�����[�,�ݞ�������X,�ů
����eI�U����4�ܦ9e�voR�������T�=8\��^pc8�ȋ^�����Av�D��׮p���"�rێ̕[}��<��`=����T��u�q�3p�|��o�X��t�z-�+�����.*�~��wL�GP�y�l�.(q1�{j*�;F�j�����6]��=��Eda��}aK'�9Rc��-?z��_���mc��<����s2M�,q���xV����ʷ�[�=�'��gR��c���4�szcxJݼ��P����'K�1l.���}���M�nJ�o��7�e�l�q���Z�v��X9�`����vٮ/�Q ��^�]�	�������U٥U��ʜ�l�ۚQ-���%;��K	_b���s v�m��u���^Q#Hve��a�0u����;�T�x���FP������	P����z[�����pY���4%Z���;L����]bδ����%�so½��e��T&nL�'\��;�Hvhq�_�vp	��>������1��~�<�^jq����� ���k4�tt��ӷT���%�.�Ӽ�7W]̩�����v��!\��.�cR+b��<l#���Z��Xj]*u&���1��4�2����8<��v'g=���^Yu�=/P�n��,�n�*����
����7�z	ⅽ�5��@�[�6�1 昛�AHNhч�A�]<�rj(�8.�E\�z�������z�pD|#��Ɇ��̅.zMh�s�M����mG�eC8�'gGFf���5Թ�A��G2�_H4_;�'��s��[�;\;�=�a��gM��)�"j��Ð���Q��M�b��\D���uf׽=u�2�	�O��N��}��Z競ST�	O8�'p�(�g*���M`��*�]r�^[�+��5:cj�\p`�ޣӷi�s{�lŔB�'�gr�xT^�4)�@���y��m��������k ڸ��+�Sý�I�÷d��rN��H���Hzt�N��:E�z�=�#���g��z���ޗ��bk{�6��<�ے7���y�g����|��cug��S�f3�8�7����R-ј#�����4#͢^W<u�f�8��ʷ��n¦-e@���O��Q䎃�ǌ�g��/g�w3^.{�
�C����$ޕ������z\��6K�݊�6h����d�m��]�6��V�v^���:��TU�B�E�J�L��r����]����+)	���9ƣ� �{51�~��mV�����U~�ٞc��ʜ��(�gu�'�)�J����0��O�"|F�G)���8�nC������{�haZg,����G�n'�1/a(7�v0�
��\��u����[D�r�{,�ŭ\�ᑂk1}ft��f��q5��9o�z��65Yf�o�����vV��̳5鏣�2�L�q��ʚ�	8��۬CζP��N�8�	Z�b�3i�ל�c=��\5h��>(��{�za>�A�ެ,����<*tU��U�]��A�y(��%�rI$�T��7n~�W��qu�3V��lQAlQDMQV3Fڹ<���U��.Z���\�#R���i�G������Fؤ�w[w��s��T�MFآ��A型U��65:�^cy���W"� w�G����z<<��Zt���Xں��N&��9�5��N#T�thuA����θ\�[-�y�<��+CAIl�͞^��:5�bQ�G�sW��9�ѭ�<܆���-Hj��S��h+E����]�����D��\tZ�����.�հ���E�$E:�(7{ED�ا�r�n�s��V���jJZ�m����snh�`+y�5�<�8���nl��D[4�5nG��q&�`��A�[f%�M[45�h��E�o8s��5��1��kIU���[Qm���#A\�ES�a�yrZ9'#�9�i4�l4��[p�E�!�v��r
J��L:u�F�A�;�ϯ~��<�,e���L��G�n��8�Ƙ��T���HI����w��vf�$v
���8�����[cx���� | @���M�˦�(͚[�P�g�ȟ��R�����nt��y�p��1����E3=#��6w�^׳�J�X�|�e�Q2Ð�!5����`��%;�ō�F��R���f=�zj9K��z�c��0(��E|���?��sȜ��?��}*3t/��������F`cCJ�������}��\;��d��ߊ����ATFǽ��Y�`�~��Τdmc�/r�A��q_���E���*�r���ǟ7��^�ؼ7���0^U����-Cˇ��tC��?�xW�1u;,�8<oюus��.9� ]k���;	NT�2�3xݳ�^���y���f1�bz��^��@tb�P2:������:�����t:M�<�%�]�����ٷ��G7߭bXw�$o�=(�>ǡ�@�����^�V2
K67��]WRq���:b��}mDn<��a�kf���<ˉ��i�k �<��x.�D���:��yQ�;Tܼs�꺾e
@����� ��]��__�M�/���?`L%0 �E|���w??z�z�D���I�����k;��{�a���?0��۔���bM��]ܷ����zg�����pW��i�о ��hl�ΕY�G
?���d3&q6lױ��y�Q�{I��S�#�kV�X������O����nt��}�@�}�Qfz�ɝu��~���o+nB@C�Y�����V(�����f�j�кW�����&�Șlh��MJ�^9c��lA����8�	޹�;�qa�5"�
�/��R��m�\�Z�V�V|�f���.f�	�Ӌ�����v�����VD^r�L_�҆ �UM�~�}�q��}���a�c6<k��L��U%@�S���U�W�ݦ�5�4ߧg��n�t�;y��Z������NAж�;
FAf��3�HH��jwN@k꽰���^�����=쑾Y��*��>�d�>���fڑQ�}{��¢��I����:#���b����"��9C2��k�^���#K��ޣ�R3��1Ӡ��/�Ч�ߠ\X|�E��Iw�J��X���z�avN�w�2G�)\B�]�7�!�>�3.���/[x5��9�o�+�+���*���8o�����1Z��>�W��KBGT��i��"�ҮpNq׎�M	�BԝZG��\ۊ��F�ބ�D����R�V�CB�,xJ����Y�)�P�/<�>�np��]��$�#Wkj:�;���0�{Zg���,��Ւ���,���yYNmS��d�H:Gy���.�0ڭ�h>���]����y���k4:�.=��/��C�M&S|�	���&;�s����\��m����7��g����iv��aӕP2����������k�G%�`z�f�g�~c�}����\�7�r ��Ćf�P�g>9X�h���Bq�);�����j1�r��f����7^�_���
fI��RQ�AQ� HpT��<����zF�0���{la�GdcI⁃Y�
�_@�;�z0��g����'s�v��c��ʚ=��Cԡ`Y`�g�+��o��F�Jr��+t���
0L��<�FE����d���@`xW��WEЗ�pv\B�8�H1�݄�5y�^�;��ϓ˅
��rR�v'����^\�z_}:"Q�S8t&��N	�퓾ˈnY5O��@�
�S�%J`��"�D�� 㘾�����9��FAf��%�7�W�}&�P/ko�׉Ȁtj���$RҨ��0�5�e�D��D����X,�Ņ�[>5xf=�D`C�*���)Sf����lW�ыHk�p��y9it纓q�/S�mPb����;e��YE�7~B}�s��j{�^g��Ovf�m��9��U��2�1୺�*0u:Nl��J���Oj5�q�^�z�9�}m飶��{a���Jf�X�o������(|���O�.��~~193��}���3������'C1���%�f��;�nͶ�<�j��ɬ��ڣ�ɑ����"kUc�V]�qv��k6���˲�U�{�p-��X�#3�6�	��z�=�#���Կ,MD3��`�/��E��������7�_e����b�,�Pp�5�̾T-m<�w����ŝ�*����ᘫ9ӑ��S	!��_�\�tX<�8�x�2�Һ;Wr��/p�b��p�c2v�;�x�Q3@�#BK`�R< 8��$xVw�쾦v�^�Xs��{�*K�S3Q̴ �BM[�d��T�Ä�P��#�.3㔄.����C�l5�S��_�UM��R�yv[R� �Cϼ�LU�^4S����2p���m���}�b}{R�j�lr�P�j��E��xns�u�LjqJv�Lc�r$���F�\ٳW�+r��u��K�@9����J��佣7�+��]*��fڐ�Ժ򚠾8|/�Y�YO}G'��Ac�	����]'>���l�;[�@╾��)˕:��fg�^0�kG��:Z�WQ	����bO��Bi
*lT�K���Gzp�)ۅjנջS�*7{��n���}H��߽�Q	N�^T"$�Mp���o��w��ɷ��5�D��i'UJ̓�n��&���p��Љ-�3���>��#�� ���s7����}���CԘ���s7�{�m�aӰ��w���^LN]����b����>��Y|���[����.�I4Ů�n�Ԯ�\�o��:�췮�>o�k��7�� ~0_�#�]~	�����{�����9�*(`p����;6hu���8��/ƅ�C��@�}j�#�z��;�r��XҴ���,�{���|]6'��90��O����]X�U��zF6�=^�`�B�fF��y�1�[΃��:�9`襫�Wʽ���1|�ăY���ك�+���]���������,�
����J,e������2v� �[Ȏ���<���]Rc�j� Ao��t��MD��zs�F��_P�e20C�S��pߩ�@o~�����n<�y�r���˭���:��d4�[8��@�t�7��ύ�(�~�m�P1\U��[Cï,�N62ҁ"Uon�I���8��zj-��nͨ�Q��`v%�F���
����[���Y}?Nu�ˮ W:r�t����X"ƫFpI�r���UnV�v26����ю�VԼ�����뉁؃�Bw�R���W�ƲЅ�y\@v�n�Y8��UX�?A��a�c�)���<~���aHN���]i�q��%'��=��ȃ�xߣ�˝�^ˎs��/�U�����}���e�tx�<���duV��A�|����I���Jޯ>�~�{-��d���ul�w�SΤi7������=�b����*��\-���uI�XCf����Ȼ�`�?>��a�ʊ������C���[v�����e%�2t���N��[�)�Ν�����﹬y��R�i��_��&�W�;���ԡ�&�Y�� �΍����'KM�~Ȭ��'_)c�������e:yċ��X�]�4~]��\�~�p���
�7���6O��7D{�dk�)Q�j���{<����l�Gt��I�A	*n�:Z��A�|�Ͻq�pf�*5�q��{�Ni�%LWC�����by���g���9�V��W����BC��/.�^��y�~�֟|�O5�s���,nB�^@z�X]�S���$l��: O�	��8+�U��v1
Åcό?b�i���}�<��爝�G��ፏ�-�=j�������m��N�ٜr'L��ч�>����]J9�N]�/��,�yr})XX�.�o;�xVm���<n�V���Xe�вd �]�+�*�oa��f��t�g���l���+�c��l�kH�tG������[J�# �C��8=!PB[5���NgF���\���5:����>�Skh8I��J���#�[R�hD0й�[���{p��1rj^\��+�,=Zj�"��f����H;/���s�/I���E\{���ǢN.�~�#�\����wD��˵�G�F��Q�׈��{h��0�;D�Λ�N�׹�0D �`�+��w�������y��z�ț�0knw�l�߄��d���B�+�}5�-ult\�|o�b89Ͳ�7b�S�@�}���\�OM̉I�g�A�^�``�WR��Ⱥ�1�o\A}j`��s��ܽ�6�{o��ɇE�1�W_	'|L�����"����A���׾`��x���`��Fo[�}�!ǜ_)�����.U=y����l�v�1�e�����I�ㄤf}�H��EԠ䛠���p��F����Gm�ik�	���m�dw�_G�tP|f�#Vg�LI�'b���o� �Õ�QrUF���;.��3�TT��,�ؠc�37^�SzݨX_d����uQ;d�A���q�xƸ��&e�2������B�+���)��������Cف�k6a[��
3�	��5�H���W�NmZ��ζc��b��������x��K��D#o�S��cm׼E��]��P���gZ�����<��$
�"~Aы��J먇���M�Z!��Is1[mк�s]�+�\u�>7�+߿r�W��'��'�C���7�{�Ce�����sfd�N=���W�'7o�<x̜�򾎷��������rp'�����|}9-�z.�du鹈]������y��Z��S�S�(�e�w8��9��Uc��wi�8�ky)>��k����'!�(wIz�{J��� ���*H�l�B�����D�}�~.o�'�=�ra�;?�wQ.����鹚*p�#Rk����?B��&����J|	U~%��8��WxM��a�9�t�I�Lg�D�+5�c�6DB"X9�!���Fu���x��Y�k��[=,fV��к��e�j/�Xf�j����VN�qc�ڗ��$��ݷk�}n`M����M�	*E���\��E�ۨ�);�B�b|ҿÃ�������k3f��D��'׏�SȚ�J=�t��hX�1���뮠��)ưU��ط+���yc�	���1{�U]X�^��F��U���:�p)	��t��|�X��Ab\x��k����ꌻX����#���=�~v0���Q�l(��CD�`�"� �4�uy��Wa�:�أ�����c��J&��nd<�9X�P�Xdd�wS�cV� �' o�>�hd���x��վF�wGp\�Bah�^"���hr�r�h/-�`��#�����d�ɑ5"r(c���7�a�>ǭ_m�K�P��v|����1h��23��s�]k��34�L���9���r�U8�,��֎��^�^J��~��E�6�,3 Ow��'�Gw�������}�6���E�a7�����ue�λl�R&��nQV�V_'�k�`:�cӒ[��$$+kZ��D���,O an������2�P�g�o	���?~ @	��6ӊ9N}?_Уc�] �r��W�
0y/`�	<W85�2�^�&^t����T�s�~뛢��i���A<'�:�O��/��켎{�6�M�aF�O_O���Q���͛[���W�4�O�_�\����'k�;!t��P��'���4u|`���T7:Y��ʌ�v�l�>����s��9���� ���8Uٌ]��y�(��C��OC���<��:�ߜ��XqP�`�u�C�w0���S���#�m)!OԄ�Q@�����VB�:*aY�&C�:�T��+6ߖ�tkг�����sJ�8+Ҵ���G��Pe�x�71৆��UeI�c���Ps!��䆱���	設\U��s9�]oN�V=�Wk��PO��]�ȟ�>���4����`םy��,�aM��V����ɋ��K��*Ϫ���ܪ�7q+��f�!�q��;�ң=Co�g�z��k�`��iq�o�B�BE���
�}|%��o�V��U��Ive��DeF���Y����!C���wԠ_�q�xg���r
@������^���T&Mk�&��u��fӎ-��2�z�4OrW$rѷ*����^�.�����CN�h��܇rVD�:w�)ngfgo,;Iյz���ɬ�@�i���.�5�ZM�[O�jZ�I\V3��k�=/���r�h�;���1'U��:�l}�@���h�G4��#v�#�q��H9B0ze�%��z�;��c�XT_��Y�g������(�,t���<���nl�X���g`�-u4l��-�,��]�E���`�U�9%�ъn����+|��0w_�Xڈغ*��"}�q����d���L۔؃c>� ����5^��;������}�v�˞���@��A�+��P��vYs���~\����o��<�t�Mq��(�n�,���Q�\�jl<j�#BO��^���?�����5�\������j�{}�U�'�Ɉ�[�m�
��&O�}2�V�z��k�?.�uP�_e^Ĩ D��[7��e���ԯc5�Mx�Ͻ=j_�?z�'/��H��A���~�n�s�O�����[ݎ$��1���o���9
�N�Y���Z�1���O�pT��P#��\r�{�%�z2�ޏ�AbĨ�T�	��x���؞^��%^@z��:�䍗�3S���U��}�-߬$>�)�J/����^��C��	�|��_ U�®aA�MAY>'��0~��*:6r�<�9uZD6�l@���ʕ�~��8MNyG�ܮzS��
ē��yDM6���o�],�J�<�0�5��Y3k^�F��f�[Dw���Ӌg�z\mL�����H����G���7��!�������y�M(/\�m{�G�y*x���f����n�^�޴p��k���_Vs2��r�%��R6w1��Q��,��V�8�#�t�z��[�v��"���y}�-W���X�OtYx̃~t�A7��ۺ;OM�S���ُ��5y?%�D�L�M�������{.����t�]���`����Ѹ`�q>��٨�]��嘂����)m���k�ْ�J�L,w�������y�P��J�)�{���yJ��)51�J��}ރ sϞ�S����2�.[�-������o�^|��:�mGy_5��C��vޙ��ZA���MI������l������Ո�d��o��1�y���r>�Q�����ќƢLb︭�k,�d��wt���w�M��u��k�b�e�|{����;����i��A�&���Ƭ�smA�^��0=}��V:��[�͖q��{�P�W��F%�/v�m�n�s=bv�wKF�˖��Ct�r�������|t�R줍���qͨ>~ͅ�p���{���׽=\�M��AkO7��Z6���R-�jXo�s����/��8���	�y��>oм��@><MKZ�]���)�XƬC���gn�H��%=A���i���r	�����������z�o��|��][��C����ڏCim��݇��F�h���9��Y��t �т�.d�*ݐ2D�Q]�f���o�v�V���O�-z���뾓��]�_9;���l��"[��lK�$C�3˵ғ�jn��r��#�C{��l^���z^����i��[��0x��JϷ��{X���w&)3��ϡ�|嚡��V�s^���`��(�5�M�O��&��n���ldK�l�K���YUo]�����뻡�M�JR���:P%0UÎ�x��\��WQ�� ��C������2
'�Hf�`�tJ|w*���7��ak�"s��u�e_��1PWG6�U/JX����j		*���lf*4P�)���r �)��KJ���Z�v8��M�f#\2<�R�9(��)�Tfl������ܫ����������T_�֕�8=Ȗ`BGp�����s�咊�PVi���s1SXuO�ڛ�-��	����j��t�RWc.;\O$��6\�w�{gm��<Gf�Uc�s�`�Đ���}k-6տ�V�j�F�;�#\X�^%� ��p7�[���W5K�M��+;h�S�-]8�]d���"n�[�E+Q�v���C��%>��'�Y�|�3������3eН�q�o&nd6�T�z�I�Y��1H瞢.ns��9�y5IAl�
tit4yr(��β��Ί<�I�X+�~�Ώ*��X��-�}N��Q�y��:�J(yD\�w>Z�:شh�g�����5�1�΋՞�m��t�F�F�s/:�Puy�9��c�u��8ml�Q\ö)���y��:�i�4v쇓�-��PRۛ��6�®lc#8�[�7}��lk����slX��\�F�F�:�I��\�	��ɪ��9ry�j�N�i�P���%�RsRr8�{\ڍi����y�@w&��[S]N��M3i)������ձN��A�Tr�u�\�]Z���h.��l:ӥ����4S��;`ѫMccO'�P��N��5ktku�<��"�v�V��k�Jr5�|��[gE�Pj���k�	+�%������I@]��RQ�����w��(�A�r�rՊ��i9&�1��zf��|q����ne�}O;gb���̺��[ׂ-g3B� �����=�O5Km<;Ս~���n�ϝTvX�|6�OF?O�"�Ϟ�>�_I�����y
ޓ�K�T�$TW�*ꛧF����7��U�_�529k/rG��s}y�I���?l���"J�'�Xo�C����D������;�~�������\L���{�slJ»�O�'?��R"B��>!�Zڭ���:g=C ��D�=!W�Kgr"E�(����<w�}��<��X�}Y��8�z4.�h��y�(>���rO�$Do٧{i�~AY^ծ�or�t�7��k�4�i�|lt���i��݋x)ߠ\[�Jw�NU��F���׽��od�gJ`@��c��M�S�	�d���.8=3L�m�ƺo\4x��˭�-�TW:�1�t�W�r��wԣ��**KbE��Bi��"����8��絴ڨ�R�릷�ǌ��63�C��s��������`PФKJ�|�t<<mzE���x�Ob����WK�~9d�h.���
�����F��}2bLؑ;��n�&U�~�_W�Q���0��w��}��yb�����{mM�J?\�3$�N�(�F�oҲ�LM:u�&н��τ�����Ź7��;���r�xq���<��f�г�ك<�^�U�J z�/�;�IM�c�e~��>k�3������t&�5��:�\H2�=w~�0��;[�yg�np�7~���hf��H����J�gsc`i��[K�#��� @��Ic���P���Cs��c��װj�%Z�Ԟ(>�l½�=΁jwD�`3�'�g����}�:\z�5'�#Ѭ@�,PTa��;<Vz%�􃰍���:Jv6�%#��I��!�>���=s�vt:��G=�@���X�诤�u�C�8��&�-�禆r��Y3�o:z�#���4A�1|�e�C21O)��
�!H�E8MQ��츎r��n#��OO�ȡ�m!�Y��pt�1ֻͣͳ��(�^�L|<Ěy+��]y�������ы�������ns�����bo8�HN|�"�71axV��W�P�DF�BϮ�~2�j�TN�]n�9D1�����朌��}b��l��a���Xck>�]���ԿC��2�v����;Z4>�T`4�
J��fWF��dy�a���!��`ſ'�Ȟ���?��<2�b���LfU~P:��Uwﺶ&�
1��Q�Fc߫����.b�f��8zƭ����uT��Νb7)��>�B����v+³�c�xJ�ȻX��������f4rJ���?\��o+�.�~���͌Q��f��kS�N�����x�t��Â����8X�X�!��ADr�sg�Nn{i{�G�u�]��+�[���I�]��3Q7�����i���6�s��F�N9{Dm����ǵ������^��wZ%Q>���"��}���QU�~���_����н���:��xQ3�&��9������=m�F�n���Z7i��j_�Ѳ�V�)U^B�+�����,A�N*���i
��=�J�·9����c�KW:#�xP�XV�O�ܸ^[R� �C�3�>T�TD�N���y���<[�}��������������
y{-��23-y���Z�F��(X9ڙ1�7��1�"�"��C�펑,i�>� W��qѕ`��;�x������^̍��+�rL�܆���{$Uc�q;������]�)�a&ԇ_@U�]'Ge�s�j2���#�9�m��6N]���Ge�2�T��͹1��N�;!t�~��h���Q�n�Sᕾ`Ŵ4R9�k����P��s�U�~�*��쨅�*�
�T"$�Mp���Rdڡ��������G�\�KvT8=�&:��iI�
�������˅d(â��j�t׸�O���n ��TF9�D�h<���=�/�z��w���
ǻ=ܗ-�?6(1c�Y��ч���w�u��&��Q��F&��KS=y���L�47�1��U�'��%�-��kqCś�+�uy�iؿy��f����=Vo^Yn�շyz�[�_>/K�A��3�}�і�*����X�j�Wq�_��fjy����uL���A��}k��}���j��KV���@����yO�6�Tܼ���d�'b��\/���6s��9徱�Aj��U�U�c�Xbmɏb�����h&7]A焂��*�<��t��W�a�����*d�^���<��1��#���ud�9X'�V�{3�8Mp��BJT��������o��D�d`��*U��ϝ��nㅘ��ٙ�R5���A������Y�iV�8�1���ul��ȫ3Ⱒg��A	4CW�jw��VZ�˔���V�<�!��0}&�r0Wζ�!��8̙�*,q�,՜%}�s�9�eA�}0�C�nM�,Eрpi�6���V��+~�c!��q��޳�~�ϸK���N�X���o�N1���C�������dF��� ;z�H&ݷ*fܔ:��n�p�ὮIoG����#O��T��l;!������k���{:¿,��������ة�ojY�����7wx��[9�;N2������|�z>|`kÐ�?r��(�}A
���\�A�D���Z�c��7�k�Ъ[���,Htq"��D1��:r��zY����Y�����8t|�}�k�ou��kX��yQ�/��b8�jʒ�|Oxg-��W�t�6a#{2�2:�~|��A����=s���	����S<��uc����^�Y���%k����wOh���"i���0��ZB�/����dA��1��q;�c��  ���cS�,oI�j�C�o67A6ܨ�3�OZ������T��~�i�d<�d
��TV��Y�,d���>�{<Vz@� ��]Ӡ�gR�1�)��3����mW��{����LX05��_�k^[��p�nB�j�������/3�X�ȟf�wGU^c����	7�e0>�0y��]?J���'�/,���0r�����L2�`���g�l�����!�7��w�(�`��2z��@WR������̿On�u���U��o�l��t������P£�3�,�C�*�xC��?y!3�E�����ர�q�]���J�ч�1#�10|߭�ڿD��P�)����8=!kr��z.|�����s���7]^�炶mE�K�`��_�T.L�D⣳��쭩Z��{#��Z�g�9�ّ�m&�C�h�b*i������\�|o�X��s�e�nż�S�@�]v��HU�`��>�w&���M{�xS����y�	���#[�$Q�pcS��LӖ���Wн��o���D�$'޾�-k|\��[��N`�N^�X�:�9�Uj�|F��߰,��IC�����1,�Q�wa��:�u����C<K��ѐV�Cܭ�
y�ؑA�]{��qn�w�-�%��+�띍�����a*fO���� @,j�+i6"z�����nF��o�;f��s��A��ƾ�!6?�_B|��G�.�|/��"ŗ��~�Ody��a�lb����-��rg�5�!�
����_]Q}�řlwB[�k1���b똡�u�o��?8���ޱ67����J��d[=:�71��D��BՃ'��gc��{&�M-�kU�����`׶���ݨX�&f�i�7>�)e�}�
F~���Yb�u�*��g 9Xe���U�Hԝ��������߿���?��</�-~I���n�Z�*f���@�:�,�&G��Öv}�k�%���������)\�o�j嬵�~�H�1��j���>��.���~����E	3�۸��<q@1�݄k��������g�Q���%�ϲ��Q�s~.�j45N)����p�
���7���T'�׻�����-�ey��5Dg��1��wZ��ui�ވ�*�;�3�;>��YO�Q'���W��ppo����#��kr�=�.}s�������~�V�7�����t�,�ů
�xj�j���#���7���j����̏YΙ����F���� ���6����]�\��.<8���/:�ʬ�K�e��=Y�p7օf20ӹ���G�����篈N�n��#E%�sr�Z�-��
�p(㿮h)�� PťK����Q@7�ם��D�G���a�⬸f�1��RDW�I_�B�sNGih��l����9�����.4�Iy-N;������G^�R|�n蝁?`=�(JJ��}w;Ҫb��A���!���j��;Z|�]�'�鎧���N���;cf���
(*}�Eq��]l7�V�GE�b\*�ThO}��~�N�o�(���
�c�t���t��e(AA��������l_+��="b8NEl�W!��}��Dk�r��zjܽ��Pe4�n�_�9�O#,���ѩ-��9��4���uI�'���cG�|$pcR��g�e�����R�� ����#'v��GD|���?4�'�@�ҶD8�����=D��$"�U6:mJ���ѕ��B�P�������"!O�Ǆ�����YTH��#�H�� �i�tзR1���u�Lkt�_�������Fީ�{݆��\�G@��M	��%GD�=ò�K�[F��1�+��^��dƧ~�7�*w���izv�;����3�Nȟ@#�_�}I�d�gl<'�0���~ñK����ˋ��G��'�Ņcԗ�V�u�)�������s����;����,����x� ��^���8Ө~����$v�;��&͂���Q��8����\�mYH!.���V�b�ȵ�u��ԖMx����U�]|�?E~D��3�sP?�Jє�)˕��_�r�;!t��W�����}�?4u|}j+k�y��`��[Q{�ӈ�,n���p�J�ү���*��|�n!gʴD±�	C��V~0��Q�"�{�2J.�l�����力�NueA���zm�;
��'
��M��´l�ߏ�L&\N��y�׵a;k��q�/������i�x୕����b<��GG��m�!����#��"�6���ؖN�H����ǳPd1;E}u9��Ӟ_o�tX�ydE�֠��<�Oa�MW7~}�g�䂽u�9KL���>0�|�8*d�^�U?NU�%����3�ɕ��U�]�H�M����)ul�װNk��õ�'U�RO�,�������8E���*��z�%���N�o��xS���qx�[.�r�t�60��0�d0�,��r�}t�4��C�
��Z%�}�ϫ�`�L9MCrCj������jJ< ?�* �����@w����D�c�*�pU��M�O@w�\,x+�g��V��+G;X�b�F(�,�zQ��c�k`�d�z����*]�iʱ9��|sOf��(�������=����yy�Ƚ�f��ҍc�7/v��� ���z��9H�J2Ȅi��sf6�
̹�����vc�$����/�Řzm�����r����'�L��6LD	c��`�"I-s�*��-��a��m}Z� Ǚ6`~��6�;�yS�+��n�+�6ϚKԳc�ꮕ��5��Q���y��>i�~X�-����?�x?����|b��s��B؏z���	4�z��6�FԴkzS��a)eMZ��HГ��������fk����lB�AU/��%�Oju��E���~5�FǤ���q��H��$Xׅ��k��#+��e)��9��qS���0��v2k67A6ܨ�T�n�|�]�{�&b;�u���{�{�>�]<
���'Tة�,�����>t��Dt&���to��:��C˱To�罏l��U�"�����/����iSښ!u4Ӆ���h����k�k��#7=t~Z�z�`�F�x����?,��s{�}�U:�#i��.���=s���`�,�.��J��aUp�_M6�Z�Rbň���nl�oA��,��/��F<1�Y��
�1��9[y���������'A%���@�A��?�/e��{�8[��\�S�x=ux���-�u��-TY���˂*��}�r?7R�LrB��w��2�-vִ���x4�â�a:��Eb7u��Z�8)��oi_6xγj��߀��뛌^o|r�߮���H]^�ͅ����[gb���^˳q��Tod�X��7�E���J�*�n�g(.a��=���E��jMú�M
]�[����'�=%s���On*�]�y�2��飩Z��/�[��tϫ��I��6�����͊`)�ر���_X�M���CA�j2�^����{�7q����=���˳�W��	lm���xxJb�ڗy��sz�]D����}'�����Ն�#2t�nJ����=R���I���~B1`p@��ܭ����M���4�Ӽ��2�Af��7�tu}�tm9����D�\;ʖ����s�Ay�v�R�9�����v�pl�^�ΠG?X���-�U\U�����Z;*�KE��x)n,�w0����X����YԜ��Tl򚳳���υ/��$p$1��9!�ԏiV����?W�\�9H�4S�bt#�o)��b�����-^l�I�8����pMwe��nG��.�Ӟ�3�B��:�X�E��I�/>�ajݵke��/%��z�/I|VA*�$�eG&��X�U&"Lݓ�u����Y+�n�N���3e�*䵢q�鱾��%�qT�ssFC����+i���@*VSZmf)���f���&�i�yN����� ��/�N��%��۸�j���Q�f�0'q�mϢ4�BĎ���CzzH���A�-�(�M�a^\;����Y��i]˳���z�u峳���:oI�n�:�P�C�d�S6� �\todN$j��A��2��9��H3*��υ��c�m��V������,���.��c6 Ì�fލ�eGġ�]�k*�p�#��|=o����~hMQ���y=�C=��Z�!�d�)^�7jtu�^������K��d^ܳd����0)��j�帹*L�;'nD��7Ӵ�}m�+�p�X�fͻ�[���]��#�9o-�I����E_��ɗ���+\z�,�0�,B����Tx���n��\a9�r����K�K�1>R�����h����bk��h�-�r�a��8�}�Z-��r��d�܆�,����ERr�UV��r�mb�!O�ݨ���1.�t�7��_:3²�������ĥ���sO'�<���:Z��][T��E]�Q��(�k��V��}sr�����8�����i���,T����+���'�d���Y�z��F�!��v�u՗�.�'��4�`�ΊE�t��rڠN�bqtH�x�G;�*2�E���ڪ�1�/Z��S0|��`k(��W0�W;s���f&<}�1{��6��W^R@�����fevۉ��S;������y��T�/{�oo�5�eu��Λ7��)�3��N�Fۨ�;��Og{�_t�9���$9���4��&�����4�[�>E�1���;u���v�x�td�����T�h��!�tS�YnE�|�s��ʵIe�Q\
�%�;ɥ�؛5��9�V�y�v�%�X��Y�w��Y$ej.�s;�4�f򺷉1���]A)x�x�pxj�΋��W4�sV���TZ�5O�91�XMe�)��k���Z��M���&Mɚ�o�����:{m�T'pO{�o�������2�n���\��K��Oy��J蜃����Ձ�W�WM�U�8|�tMԹ	�e�U�-�g)V����Z��UcɦNӯk�P��<r�o
g��x��M���n�c����3�d�����ir2�������}O��NbȖUjZnM�Z��Ic��C�ǦM[������S��_R{�5���g83v��z�SЫ��K�e4l:�B�v�d�&�ɒ�v�V-�Qj*ú��yZN�#�Żp�ՁS�ťD��c.`�v4*'WU7�G�ox�wwwo�t��é$@�g�x�I �Zi5����AISI���?'�I��
���x}�^�'�5Ms�(J�wwu�A\�c�JU��s[G�CA�1��������9�QMZ�M��t�9j���y7{���^�η-p��7eժ4Q�<��<��
���u�c���U�l�J�n��5F�Û��]9�A��rɤ�U���4�RuFz�E-:��Uru�k������7|�F�ƫW\����4�N���:*"�lr�.M<f�����LDA�0u�����Qm��g��sd�킚S��f�m�x\���E����h��G|4����h�K�9���mj�6a�m�&���\�q<��661��0lힷ8Ѻ�"
��d�EQ�X����V�UmN#V�΋f��w��1s��A�VګFجQY�&��:�T+`���E�m�F�ti����QKlPkl�Pu!���w�n{k8��<�⾆n�Cd9OFuqns�6fH\�CP+��)8��y�����͘��}w�d���g�� 7�P��50g��?�M_�U��8(c�5�z������E��o�ڮ�˿T�52�U�{i��4�9�/�1d(��Mv����wW�ٛ�����s��h{ëN�U!�lS@<�WLpaV�Wyr�a��*;��:+|���^�$�wڅX���Y��oMd�3�pw����;W���=�K��]n���=�A��=͊��+KP�ȸ�Y1v��Euh��kλ��m��4u�� `��AI_��W_ӓo�~+�a�E�]Yꝍ�	{��Dgv�����u�e�ڂz+����z�ʞ�w%��5��?,P���²�-��m6./�|���VU�P��=��x [j!iZ��2;a�{��F�!��$��ĵ�%�ܿ;�w2�Յж��Y�=A�������zYɱj+G�8p���m�i�֬��>�/�H:b��߷n��˕�U"���*w8V�&�B7m��A#���,wvM���Kw��2FQ��l�0�\�vHa����|.f����Co���X�t�ӽǧg\��V[��5��dֆ�\;�o��3����ɉ������={c��1��6���,h�7��P���m'��ODv5�vL��aT��>�TQԊ�̻�P������$>��Z��]�����x�s>��;�÷�6���<"sPӒ���W��uh@}RG���:��ۻ�N^T�/��t�9�1���]�k���k�YO@��_rˠ��]�جVz �u��w��&`��S�ׅ���ieS�
Y�����} b~@����:wk��9�;ȝ�h{�?,Y)��^�u��Tl.���1*�N(�<^���"�n��2�@��,i���������_%0m*����M�:�+�x^M����.���p��]1�Bij���}ï/Ο��R�q6��{5�pr���������aЪg���zob���B�P����f�yY�o1"U}�cZ𯟽j��>������Xn���Š]�>G��[^T�	�\:�ܘ��o!/O�|{j������ƽ2U;���p��#j}�(V��]�X�MW��3W�g����	����S�6�a�s��z�{����F'�f��Ţw3��zCUt�B/����{s�����։��.�K' -����ׄ�W�o&�����+k�{�'V���;��?b��k�{���K�B�������x����}�jv����J�������Z��'7�y*�lUN�ż�ؽ����p��`�NE�,�1`N����xV�ݼ��٢��
���T�-\U�[���@�7b�y�!CJ=��4�����f|g�Q��gV_ZtUŘ�����F�{A�lu��C�!5�>�m����O�tn���C�r�99z��f�^�p%�`G�=����6p�}s,7t��,����]���0����2���ɷ�zћw_#�yP��	C�O&�m�a9�Н�E�0�j���0�}�����Sd����;��c�_wY��ɂ+���A��*G�UH��#V�-�[㬜���,���8dq��eׇ]/E��Rs�4y׃4$"��>�����\��d�R��]h����L���Oef�^������A��T7��q7�S�#���A�I�P_���`B8��{�v)�x���˗底�m���s<�}�vK�a>�i�P~|/�q�4�G�z��N.	}C��R{$�J=��BL`��u'�/�"�)��>����N�ܕe��߀�]"�a����>�O_ښ8!o�N��{C��˄g��9���z����4j'��T�՟z�7�
��B �����������u�|��H������TK
��k�����w~$%=�B����C�﵊�kc����>�U���ڬۚ��+U��ә�����-��O��=�A���l,^a��[}��Ɔ���j�>D���d����+�e��j���?���}][x����%���FKY/�����vw�齞�Kl_�ñ�� ��z�UO�����Jk4�}U��CA�GD�/QB+�1|)�>�{�"�4B�m�6/8]���7�C���QK��¥�O�y�m�>�V��r9av�aCc;�^q˻o_߼1�7z(yYkA��=�j�e�N��*�Јa�~�ۺ�/'��^���V�0Y��.�Z�n�U!|�M�f��M,�v��5GW`]�Zdf�T�܌�ޮ�aD�|}����YK�}ޡ�se��*ɾeNa�����>w �"DVڻ����|�fǔA��cr��\A*w�q��[n"��gԧ�o��r��R����߇_�Zϗ��;۬�$>3��::����f��q���r�/�?��v�
[g>���>���l7�[���%F��hO���]_�/��k�������/-Œ������U[���u�����hU���o��\�<O�8Ԇ�����䷽sy� �Ǽ{/f��r#�sPD�t�?3���
����CjG��X~�/��c�`���w�� L���\3{�'=ƺ�<�`Z!PU�
<��7paPOes�x׭��}����/V�x�`�4�`���^�Y|x*�����d3B�`��՞k�q��&�l��uŨ�x1�7'���]���������+%{p��5S��
�W��k��kb��b�"א����,�/l��9wc����1bj�M��	`��{޵U�g&�����ͮ®��xUwc���cY#6�G��S-�>!���x���[>E��ZF�{6��g�s0��j����!��_���.Wf��[㚵�zY���n�һ�� ����U��I�mM7;"��WÄ�}�5�/;�b���}����\�����|7֕{<��W�я�ϑ>���{y*��~a�F�W�l���:2s.0�LJ˘Gv���&�ka~ͷ�L�L�n���U�ؖ����_5��g^�RWkB������Y�k-ܿ;���j�м�#�v��⁍���$�u�J
�8C�
_m����{�u�(��NN�a��OMA�����N =�ܔ��qz��x��;k�v�A�YO���}W��x���6lC���d�����Yk<�k58�Z�7~���1@q�
c��������Po�E�� i��}$q��O(�F�6��툝Ȫ����:{�$�����,�Z��[~=X+�Y!�>��m���-�i#�ʵ�yaϥ-x
/�4��[�Yc�;�?A=S7_O/�c���J;��W�H�����ǟ})�������U�v,n\��|�������ںz>>Փ7k��u3�&�{C-�5��{���BC�j�S�F�pQ~E�u��ܞ�}��p�r9>Z*%�HBU+�.ت��a��{Ľ���CX/�Ëp�?\���}n	>�0�����&�:�L_:6�	��z�=��#���{�5D���~��ā�z%�߽au��:��r�0�I�}�7Bb�Փ�8V��v�w�V#4�.>н ��\�&�w�Y�V�l]��L�z򣙬�������xc�Ւ�1� ���_]-oM�b��ꆷ��fO\j�T��	�0LP��}c]/@6��}�*\�W��Q��mo�(磼d���_$�c�-kk�{��\��&�нљ4!P�/s��{���e��Z��|\�����[�ƭ`
�^#����0�lz����T�qQ�!X��E�,�!N����eSg�ݼvV�E��b�	����e�-{.�͍;�1�/���+�(�M6��#�__Dd���Z;o�툋����m�	:�F��PChKc���zBk�#�ETa�5���:��}�5J]�y���l��3�%�`G�=@�1�%��A_
�~�W���&�==~~��6;��Xh��nާZ��5���K+��1F�=ݛ"i]^���f��<�fk�;��JXЊ�b�t9i�v�Ur�N�۴:��}Ћu�-�Jnfֽ��(�����fS<�o���v�G��>��޿�p{-�����3X�Y�q�W�0~��;;�Vɵ�v�"�ʬ	뽹��U�}�Q��_��5���d�>�j�H�G�U�,��w���_���L����{`�7�(�X�n`%��k'*�����8�C�D��w^ex����+~����Ճ`���{��g!s������ͼ��S5�sG��A}Pо�������+��WC��*z�4w�~�:�{כ�;3�z�%����A+�`��1<��i���g�i�w]�
�������Y��|/�	�	��+ �JF,=24g?��/�;��*���3�ż7�׽�������_z�Ӓ���EJ-n,�ul���Lc��YP,�֡�ᆏA43�ή�S߮������̈́W�vޡa��{�l��x��W�O�b7]{*��G��в��)_4*�����{��-v���B#�_{Ӄ!�ѝ;��L�Z 	��_����~�hcӰ��>���ъ���h��r;�WQ��Ԏ��܃��U�
f�������WI���TuXD.� wF6���,�4+[����p��I|�`v�n����{�ʛF����?�/�jgn8�֊[b*����ey� �H]�Ƹ�H�YՅdO����k>�^c>��o%���F�!�ؼ� ��q5wۮ}1���2E��,��i�m�υ"������W��-���q�\j�.�6|b674x_t/u��6������I�F�����r��}q�=�/]���9q(j�T����'i����Y?��D.�.��zY߹�Y�v}u����	���R�����b�5�ڮl�5�!*�'�\]U���@���u �Q�-
[���,�Q���,�Y�JMO�Weʥ�`��~� ����5���H�X�H�:Dֺ�.�"8�g��I� Q8��i[8��B���8z޲�oq�]ت�R����tg���k�k>�ops���]`Z�`���#8x��2���5ܖQ�7*��ّ�Y��<�9NV�(��i'�o��lp����k���6%��y���kPQ*���K)�V����a��G_�� ��(���{ ���Z�Jo�AYE��`��@��]v�%eh�.���{�>̺�/�쏵I���N���'��/�:��X
�,l���g@岨mۥ
�*#}��<b�z���t!�aT4%Bik��`k�q�B��)m�`�^!�	J�rn�q�x�z�\���(��'|��c="�pk~��ýϬ{�-aogFT���"|�u!��A}�8������j3BU��䤯�T��(�c:^)��p;�T`�˦o��ˈV��l�/ݮ��U�����J����;nk�p~�Z�Cv�����!e�6�4��H{R����� ��FvFV�*�z�U�'�g������w�Y�6 �����yM<�'�lw�^ԏvT��~�Ǣv�5�<�"C�g�<p��≦��M=	�*Ղ�ef�t31�4��cj*��/�6�ޑ@��-�W�S��k��e�m4&(�h3��}�����F�m�TGe�0PF��;��	!�Qk���f�_�P��u��{ѕ7�p$v�U�,�p��`���-��;F2e�n��6�Z�(���wk4G�#u��nb�,��|R�Ὠ���7�:UR��u7�]��	��H�k{���)T��ӊ#,�K��>�[ʏ��wk��m�ek�*��x�;ǖ�.��m���&���jy6"��t{���q���s'��Eպ���Z��V403.�H֝�=Jc�c��7xZU����+�{!��GHi�F��\֊{�^���ˡ��S-��[it͆�>���Sqy�1��%[�5�۾�LT2=����w���o>o(x��<��4t.�=� ��J������V��=�h��p� ��t��
^�dCu�iŊ_n�
n��*�3э�Ŵ�A�Nu�W8�U�8�����̹z��n{ћ���8���Of-��G#���_^�`�%�l��xG�X��|ϨU��r5�ވ$���O1`���7ö)��r!ڳ�y�Ҝ7j��S
���E�Yzh�j9��Df�&�������h�IV�(�`f)�N��	��Jy��N��kI%[��e���*��AZ�I8��R'u|\	z��u2�:R��j^�۩2g�~��H�$�}M�q�L���(S���c��O9��[�(,Uh�j�f�r�Ncv%�����ʈ$�ou1+�F�OYf���q���-)"��ܒY�?a������M�8W��vk�[?h�'�r-JC�>;V�a,_}3�/��U��c�ی[��Z��}�}D������{��p`E��9�j�N�KQ7W-j�s՟�JW�+�u8�ɜ;n��r6�p�V9�t��Q��h��Zs�4��Xx�,�Xn�-;�ՠ}�AH�i�^4��|=3 �ٽe%��Z	Џ��\����3A7H������Wԑ�ǁW��ج�]:	�wM}(�WQM�ً���M�ݐ�{���^j�v��+��������wB�5�D�>��s#6�*iۧ'��y�|������W���Y$�{��D�Q�%�Ә��҅ͅ��q�5Yn_/1vgo,�~�K���y(Fva2j륝%����V��֞��:����]W���*�����r	�Q�v2C}:Wf9��7d|a�'%zGZ�������}@�&`_{�]����r�l�����=�q�#L)�Y���u�U��}�������cA�V���*�ve��_2���䃝0b�(��N%�W����X��f�[�C�O7m���GL'�	?�k�˿�s˳@9)��No�nmdQr�K§X�k$��y|��u�v���H�'VEm-û�{�!�⯳~^x<x����T�D��3�uS��|$�9Hѕs�l���a���P�vu�$+6�_n��_RV�xE�ζ�B+7���x��!u�=����Q�����m�����.XYt���w]|&��7η�]q�L�:��0��I$��C��"�p��DG������{�-n��/�q�Ѩ��f�Q4Ѣ�c��v�k[[�E�ˑ�AQh(֍Pc���<<|:�M0MQT���]p�X�i<٠�Q����b��6�l��c8vxxxx5y�Xӈ�Mhŵ�I�Ah-�V3��sDX�j�:��(�g�&ӊu��F�U�U�q4RyQ$wu�1��(6�ڵ�����<㵗M���r9��SDZ)������j�b1\�+ Ѯ�Tr�AD��đ���G6u<j��cj���;�ruE6�w�kV�F����؊�j�5����Q�AU4Mu�r���؈�64ƛh"")6Ԕ�����lS�j��ճ�X�E��.l[:u�-��nd��r���D�=\��2p�n��p�kV�45kh�#SUT�cs�=u���ʹ:��X֜V�u��*���U�3E3��ͷ,�V�M��E�l�s�9�9U"��P�Bo)�Z,'�j�ܜ�ӷ�򸚆o^��VV�N�M���agqK(�$w���%�T���vi�y$�FH��lU�h}��}��g��W�Aj�i�ꁦ�>�7��^z��M��6�Q�Kw��ڟ|��m�?c�5�;���d�H@@�c��Os"iT��{��tN�۾��,���(�ϓK+-�,���ro��3�iD�Y���<9�xD!c^��z��Jh�.���J�@.��o��m��U=����39`D���<�;��A�$���H�m��Sc��1+3���u=v�`j���a.�^�kNJ�˽��"i/X���W3G~�=硭4��"��|1�VI��aU1�������+�X��5�Ή@�r��1:q���L�~b�j#=oGVJ����0َ�S~�Lq�3�E����]j�S���9�qͅ|���ߴ7�m��e���T9�ݝ�=�{�v����v�J��௛B�]|X~�\���Z����G|L�<����-�<k���K�uyx�����6BK�N����˕P/��7V�Ɲ�Z���h��ܖ��]#|��X7���-�n��׸�}��:��6霔�z�jv.��ʋ1��h=s����s���~tM8Ppn�}�N� �WC�)}o"��r���=MاS�����m���!��,'�[xv車/�=�]gʝ���H���깿Z� �m|����iPҍ��mp�m.>��)R�gu{�Gm�;,6�g��o�ܗc��C|.��7�����{d퉺X]{=��+x��Q�ew����R���̕����0��G��3�zc�"�ǎ;�9ZʈHa��}�p�-���ɷ�yu����YQRnTe{���7kԔ�&4��?�����|�X��V�g�T����0��t�];xO�c3]*������z(�X�ngĶ~�d�e��b��R*v%��^���	��%d��
ہ���;�h������ǵ�т,�TO�[�
�X�q�t��t�p0�Y����\D��'׊{2[������}��#��ߓ�֝+�;8!�b�
'��TKՆ�hh���8o043N��D�qs]#ku�c�>�|}ժ�����[w��h<��;��Ê��.{�9{Ǌ r3�?s�k{n��pz ƚ��`!����&I�.��i�F��F�!;#<p܆4̥��G��6kl"�J˂�"����0������]�R\睏��ժ�r�8�]�Fh.��J��e�K�ubOa��E��%�i���-��Z���B�rHXoP������t���22-K
���cz;Lz���Bt.�����=^��6/ha���V�ǟ��w�(Ez{��s�~�?`y#���|�^�s��0Վ^�z+TL��H�S�z���(�����)�y�?0�pK�3�^ߓ��)��v����W�VE�Nđ{�|���*V֋�%�E�#��H|2�[��ȕ%�8���f����t�������ǔ���grY ��aOE6��gr|�_��vp<�cH"�¢���FM��a��I�b7%Og�b���d���㌙��O��A� ���x���7~�2�6��8���Wn�od�����f]�(��@�7�%o�v�R�9����T�ߔ�?i�%�6C����'��ǳ�Tƽ�1��u����i(���#��I��%O!��:�z�g��o��e��⎗lL���Uj[�]f�ZJ+-un�(])��a�#�.C���D�Ӆ����u�r��:6��햞�yY��<8���:�8k�LȞ=��LGM�o�P;�����������v^KqB9}��>�C�+
���l2J���n�r��Jk�&>����v���~�4
W�'=�SO��B	ѐc���X')�J��l,���C����d�[`��կ����{��<�X!����g�-X�B�Q�HZ���7^�
7����Bƺ�i��X�{��iҳ�U�eA���.����&��w�8w�����U�e?��~$�5ĭ[׾kA ��P��q!@���m��	(;�,?TK�74G�"�'��1X�U�8�Tƪ[��_��=��W�خ�&K<q�"#�n��RR%�K���j����]��˯�T��Ne{ER��Qb|�,�P��_������;}��%���:�W�7�۹��P���>����:�L�A�H�������O��a�}ŷxދyOȋ[�����!�o�]g�ݼȫ>̮w�d֪���!K�y�,�ͭZȆ�a(�%�g�"xG��z^B�q"�Wy�7^�y� <��^tqC瞹w�	�f��:uN��Z2�uc�k��v�毭lN';HZe�1� ��}�/<1燠�l}�-�f=�*�W&�0�x�b����B�.�D�;���X�Z��*x�|ş3pXk�kE���Gfw�+܅4o��1c�"�z���A�_������P�*�6��4���QVk"d��]ue�H��n^��wޑ@�-3�AX�)�Z�m'oU%��~�zlV���0vr�B�z�:�&͈q�%�=>�-/���A����A}~�
%{��:b���qs�ұ�Ej�Q�ꁧ�����],�����3��Y���,y/f����k��Z�s�$�	0P�9ޝ���3G��vb�^�-�#�X
���ǟJZ��K+-�|X�[����E�9�W��|��9���4.�!s�X�_x�ϥ4r^�u�
�N�D_D��R���
����İ�x5F��uw\yiH�i��ꓚ�Eq�z:�9亝��b�tC	p�駫v��$wN���"���,D��&eu�_��g$��*�p��.�ǳ>�=�_���ȡ�Q~���IQ���ߩ>Jʲ���R��^����%y���5j��İE���x]���1�z]U"�q#�`�����j�d�;�|���+9�5�����6ױ��������aU ƪ�Z��r�fh�n� ���6v��?b�	��ϯ�1_s�/�e};��P
<ړg�~b��1$�k{;~��s��}T���9^��WɏU�������u�U���qG����P��k7��MBx.�W��;��z���l;g���lm�m��U�b@��RPܪ�[y=`�;+7�h_�y�ӯ�����U��jQ�b�(�}�U�x'����W^�Vn���粬f��AHr�\SO��+��&��������3K?�7�qČ����ş6�d��r]�(!�-�S��;���gGy�o��=b1uL�ZoA�P�>�%��K��{�\6@a�����6A�#�H�<��~�r1xe!��6����u�����~���[�&
�}�U}57F�7��u�cX��O�T:윣�piVu�v&�cd�������W��û��#1�,"w��FA~�zNZ|�چ�����'�]}n�Q1�����r�i5n��7�ںpD��z��ٗ|���cWc0s�]�����{.M��6G0���k�rg��E��|R�M�ۙ� ����eЍ�M܏Ĕ�W��Q�����㒊��|�\-�[?c�T{��TMU�'�\_p@��lj�l,�?{�c�Dq����^�ǒ�;��[���f��tJ�4�Ge�y�
d��`��F G} �}'�g���쨽s޺�[�P�3�w���[Z�.��+����D�<���|n�"]�^_w#���^����*"��{�����>x�Y�[�N���n�4��5����k{��څ_ܒ�9tW��Z7����ٯfg�=^��CU!��u.y���^|�G����Z^=�vg]z�]>����Ĝb�^I3����Ne�_U���x9i.������#�G	ZE�{Fatyv��MJϼ���4R������i]rܥ5�:\F��w��u�x{�R��Z�\����M|/"CӤ4Um�]�e��^w�"�U)��yF)�(|��	��+.�~���Mg�I��gj���~�L�݁2c�z���t]�t�;|�1��bB�[H��0���Xt��{��&��чV2�x�����,�w8KZP�t�n���Cz���1�}�/��������fv��x�i��=}-��)b��-��X�VC���$lݽq��Z����	��d�Hb���SK~2�z ڿ�*�vq�`yR��(R<y\����!�P����liVל�;~�.�{����x}�~으T�̛ꟼ�ٱ����^�!�6���l�n��59�=f�[�Z��f;{z���x/o/t6`,��D��{f������&j�~�*�{=�Y�v/�Iy��X-�X[��`H=P*�wş[�y�����=�i{���`������
'�i[8���0�/ܠp�ک��I��I;�fs���=���mk<9���]`�jŢ�~�x��%`�����(��&^m���{��g2��;���UGm`��q<7�l+��=�k7$w������^)�k]Î�U_ܒ��ک��j��w���f~��w��ȋ�qW*~��ٮKj�c��#�S7�t.���C'3��A�<E��qŐ��������k;��pe`;C.*n-&P���y}�����t�zl#tۧٺ*<�	hIǘ�vm�z_D�1&�v��]�&J�D@��Ѻ�x]Q�E�v�KB�M�ULj������=�O>��Q}&ؾ�^��l��3�}�(�܂Z�"����k��s@P&�n��{ؠ��`�
�9]n",O�=(n�ug�o�.a���������V:�Xȩ�W���<^�H�=�j��\x��Ux����ĭe#�n�^O�˷ҧ2c�ʋ�y��D݅����{"�w�Y�7�T�$[�i���sz`��v�f�2��*���^�,z⛱�!�Q4�1(ߦ}+D����������Bg��^E�p�nJ�BE	R���;��5kUmnz��^R���{��Jy7���O������'�Q�(W�1"y��O�F���!�U�n�ǲ�
.w�����^􆗥�{�Ӭ��F|ߴ,��Rr*����W[��Bγ�{d�]��l%ܵ�Y ��>Ч{/#Mf;�����zO��W߸P�I�>�On�fN��Y�ƾ/V�/���sB��w#��Y���y�S�_\�b���u��y�3:+���+���s��J�<sl-��*����3\3�MF��p���VsSfaކ���R�L��s���Ӝ9V�W��o�������N.-�����n@WCc�уE��^�H���5�?,5BG���b;�;8O���u��F�wf���5�@���:p3b��Ha���Tգǻ�o�5��6��[��T�ߴ�O��4�zAtW��;O�0�9��	���:�Ǳ��oR��Ɨ�{��5$�1�lPl9ױ#��[6z��?0KӐ�5��yyr��]����.ϙ�8�y���*��	���{=���W���őY3��X�\`�1�59�m۷�նlX:°�����8�����R�>{�6�����v�vLx �Fr��Vsy^��ŀ����ܕ���=H���WU�a<TU��b>�y�"����K	�S*�Tv�b���.�{V��>�n!�b�w����]��b�9(e����_1� �f�ʚ�fD�/Ic퀪Z�Sjaos^�O�����ᓂ��{�U^%�p�_O�y6n�;i���vGXȾ���x��*�ܲvUkQ��}�������)�,Ħ���Suv�zw�s'��__������@�,�y��q�'2��|Syp��\U���xƳG��^�<��=�;�ԗ:t�����ι%=r:/{�:�^��;1��ջZ���� ˒5_h��!��Ch�����X/<�a���0�|8xj��%����kz�{NL��������"���)���*sǽ-��Z~�w�</��w�aB-Qڇ�!���\ P�i���o�� 6
Y�v��/�5kx�	�!�<�Pf8̾ͨ0�y%�t6�J͘������o����ݺS�e�e��X2��w��G�k��o2;���nT �%�kq�~��R��8j��ρ�yK��^� �7*��1��v�<��҇wH�Y	�+�{}����&���9����xe�Y�j�{)��b	�+��x:Q����S*3�uܩf�����'uwZ8,B�]�' X�J�s���.���Cp.�{�m�ik'�J�����Գ^we��n��Ý��4GoMɻ	t��5�m��W���.n?�����)�V�T�;��L������ �YV���̢�:�ٝ$]��qr�r9v�d��D�pp���Br pݧ�\H�Y6[2	yA�u9O��,:���!%�wFo.:Ƈ�w7(z�B�sHJ�����?m9���j�{n������R���D]#%���]n��[�I˸�sG�$����pe>�.�X��6���pƂh6�n��*�V�VE݊b=��)�%�n�7\O��[�RӶ�Vc�Je�gx�j��'�/�a�D����{׶�F�49�z����.b�wlݳm�������ذ\�!�0zfhr����憫[��_+~E7�ª�7�[Ėf�D,ת�뽼��s&�퉪3��%�,���×VD�sY�ַ�T�A���.wX5gj��f��zm�S�]g�f��A�k�U��9QNT��[��&FC��ۼJ��q
쏵�u�P�o73�=O�ɷ���]���f��y뭣!��	�\΀|��v�9fqws���'���/9�q=��-�n�m�;Ʈ���z�GV
�I��w��TF� o0���d�R0��iٖ�L1h] 34/k5G	���_�}`�;�@�x�w�gU9��toi.u��Nd�/1_m� �Nq4\:�C�߮��]Ւv,�x_4���\��s��0�`d�6d��#��W0�]BƗ�9�Čf��M��Ч����434ԬǼՔ˸��`��>x_sH��y�sZ�z�%��͹^{�䊁�r�����Խ�v�hKq�4�ڜ(nv���Y�2h�j�m@D��(!�g��>h�PN�n���(��j���56ѹQܠ�I$���}'K��;M��D,�B ��b(���-�u�9EE�Pƌ\���ڢh�"'����QQ-�S墣N
��4�Z��cF�肋��6j��g<<<<</h�z�
��jj�i�b(�&�ZŪ�=cO-Uu��UmU�ZLS��v�Cִ�1E��-4�csr*�EPr4QAyn�j�4i(�v5�s���X���p�y����[\���Z*ڱZqDͬn�
����+�TUr�U=�����ԇ#rrݙ�U�d�)��8�����خ���6����.N�]Z
�����EPu�U��D��l��Uݺ�ܚy�E%��4Ms��G#I�����<�6b(�mD�UTLDQsi��� �DEDQ51DI�TrL�#�"��UCh��j��놊
����b��u�6��10$�	 H�p���w��[a�g�b�ﱅ��c�A?�I���L��M�߽�L�v�J�r��\c�{+��i��η˹��'��sO4�����@�ڃ=0�؛N����|��mKc<�/d�J��b8���o��m�2���6��6��������6�/�ٖ�Ј�>0|ć���zi��5�۬ �e�>��~���z�P|c��P���7(Rk�������{g��}r-g���9�ݭ}V16�>l�#���"�V���+7a���Wѱ61�������~��`T�/���B|��_ui>����>���uv]/�����}�=ԇVl���5����b��׷�8�{y�	=�NJ'�]����G������~ǳW���<�
�l_�O!�"SG��u�J�c�@��s+G�~���7���~��6�{�j�r�8�.a��\?1�.�V�
�{I�;L`rǃt&��=���-��\��w������گT��/�6����k�*C�@K�dr�d�ѓ ke4�Y���Q���:-g�:���s�+ݣ������8��Tcr���p��G˳��6�r��LX��$,���6�����NІ�n��H�whk;ho7���n��¥Ƿ�J巽g-�y��U� ��G�b�u����>�^|�Z�÷D���<�^�����AHP�gX粯�q#B�07[[�_���WVװN��(�v��GD��2yG�=�������ϡ��^�a��d�H{|��Z��)T�^lWb
pՌF�}K�#��y5y�)�Ï-��ܖL���n+x^w
�]��j%�n��V`�k�=�ǝ�q���η{���n�RX�
�����ଯt��6S�j�d�;x;�/eW�eOf�7י~��v8zCz��o�zU��=�߭��l��["��B�wn����m_��vƵ->=?@�'��m�նpio/#D�U|z�xK�µ�[�H�"ǽ�@_�0/T)��I�{յi�R��Ɉ��5Q���e��C��`I�Y*��I�md	���j�ĨF���q^�~;�ɾ���S�ԯC�r�OYg$D�n�;�wI֎�xɯ_�Z�^�g���Xd���$��QǑ�!iG�����]��Sz�]�gJN� �@�|�CF��j�Qc���&����c�Lܜ{=e1���} �X��f�퓶����{}�|f'pD�m=�<�8o9y���E�T{}	C);�nG!�9�z���3ȼ�X!��9�5���ل:^�.'s�+o�vj�R�ƏA	�^ӟz�{���s+>*аTWbVxF窴JYSG:}��z�}�^��|j$0����x�W��h$�T���:��]EϮ�Vi�뽖����������¦5T�|:��|�x�n�X�XĔI��I����.�/�E��k3s�tT��7�϶�a�2]��7r�z�Uɺ%7���<^���{�w����c��9p<�������@X�@Ӿ˛τW�B�o6�{�r�P��h1��͚Ԥ�o�L_f��o�'�h?\�l�_!�|���"�^~_O{Ӿ�O��w'*��+6� м��׮Z����!
�8���mɸj�V�"���5+��Z�-yQ=ef7�+NJ�L�oL�;�M�[/�?�L_޳��ӽth�ҕ��N��}9�
.�2����������7*v�kvd�Æ�����{d�¶��d���󠫍8I���:ͽ�c�EH�3H�K�ჇN�����W����5̢�d�6#r_@B��a��"v&�J��%��]��
�8�޾�cO`۽}�	�p���1@�R�~+0�
d���/]������-}^勞�Ҿj�rz;~��WGYW55�+�ֺ`�UG�
�g���MU��~��h{��	{&�\2(�f!T���9�=�:B�}~�~��I8��}�4���t4a=:3o�&"�aQ$99s]�V�`�G�����q�#��$͍9��aN}}��HV{�����F�g���p0�^��~��}�bs|��|�b�6��o��<�0\YTo����'	�<�!�^ٛo^ElA��Gq�=��}���߯�l_�ß��H�-�͞�R(��-�drwѪ��3�w�O�ζG����U��-��j+��v:�W÷=5������U�_��(�7�|pm���	��c<���|s�ɜF�f�d�V�f��?
Bz{�8L�pl��ۻ��׾��`I�]u���g{e"nE���fY������y��S����Y�7��H��7]J�������ni�ow޳�<�R5k���/�y����#��}d�s��ŝa_�kX^��ї;q/�2^�\�@��0=�z}�^���k���l8�#-���@�Ν��촼u�g}{y/ F0�������_{���$��"��֫F�
����/>m��f�.;{.�bh)P�-7�f���d��xK����Df�w���R�f�&ӳ=�n^�A~�k���ݝ�U|��Q��s�P����M6ۗ�{�l��?�}��i��9��tH-���G�����>�M;:泛u��/��Ͽ&��#��^�=oM�_�%���t�c���jP�c���;gK�:����~��rݵ3Jtެ�yZDi�[FB�=��ꀌ2���ࢱ`T���.������|�/o���K,z��?{��rtHMY�����E:��˳:D�g�ֱ{���c��݂DMpѵ�s�'��o+����t��%�8�R�*;DJ��nEN3���U�#�+S8����%՗w����x�c���Kiq��5�K�1��:�Y��R��:kO��vȉ ��{]����������w�4;��~���36���=܎�cW���lW��[��SG!u��/��߁���������P���j�wX$Q������%q��
�DX���4�h��1��)�/6��*�#��<���E�VV�ܴ?w������ZR��9� �]ڟQ��\�'�-�O̻����1����Z.�ٝ��̈́弩uT(�)Wun?#��hūH���E��.y/�Q��_d�_9�~y7,3�`��Ez�B5�����+��`	�E�r��W*��~a�T��X�^	麔s��'M`�w7^F���,�1X�9�#�`�l�͎^��څ��kӵ�w$"��P퀺�So~SMgͷ	Ef}>�\.�uU7�*�����p�.��z����?l�6��v��|0��SK~2�`���z����l���9������d;�]�k����8��[m>5|ũk:B}{҄a�]�xN�=���{�yw����i�]j�&Z�벑L6���t��+�r!��A|�y�,zSE��F�Ѻ
b��n�t|�.q�[Wo�˵s�Yz�3�3[�wz���O�7����C*�3#�zU��h��`�p�̣s��P|x���BV��#G�="�	����m��V�m�*�Lp��+p�A�^?j�cX4`yv@��z�����@����g�φ�k5
���w	E�d����s��?w�!�Ж^
��ݱ��ng�?h� i6�s�cϥ��\����DpY�u��)LyI[��۽�������=�2B����͠�o�����"����1Z�o���0g{˺n���{�,{����ΰ�7��}���kh�����sDws�r+�/U/69�5S�U	��+��A��))�Ƿ^���rA�}��A.�tV�Y�X)�e����s՝�L�3����:ͦi�Riy_3y{��ޮo�W_�1V�ij9�������������7I�[����ڼDn�7�j��Szy�|s���ˢ��gC?c�gy�xz�˳��G����i	aA�5��*�)<�ɮw����V�7�O�՚���VC�>���ow+<������%�^z�����9�����=ҋVŞ�_�>W�gx���a�Wӛ���wJ��S|�����ō����N���6�onJx��N�z�85ar�z݉Sas7�o�~�����?+����3�%T�=��7�͉c����Sb��!g���ʚ!a�$�^�*ĥ�D����i�u��A�y
��-X�n��+8�p��	q<#T�=�LD���3\�R�pl�F��!��g݄=͸G������9)����@����i�o_q���Z��e���p6�D#�i+=u��6���ֵ8寪�勛i!�A��H�pn=*�z��Xj���oC���ïUsϫ�<N�/g�hj���lr�D-|:Ez4�~��ӕyo�tr�<�ri�8�ql�M,�f�z�FNu�o�(Y�l��]��U	j���j�q�|����-_U��
���0f݊�n�S!YB���s�$��0VسE��l�9�q�g�p)���Lg�3[�#<�{2hF����m]����m���F /v�ǐ�K����s�L
�(�l�ؕ�u�]���ܺH5O�d��|��"^��Z.{7�rg�x F�u��+�h6#�q:8����Hm�����;���#�%ö�~`�п����maP}`�6�b�����wRqG����3�{r���������;�Pӭ��3���9�G�M���������W/�B�1� ��=�_�ܡt��9֏�S��U���_1 ��l�}Vv�5�`��]���*WӅ��,��%�f�|�l2ؿ���%�w�jG��eOR�����jӷ�u��{_h~��+�;��J����N��Hw�L��y�B뽣�69v�G}{y*��ú(�e�4/���=ܕ[�3�=���53~�@�xU�ۦ�ٷ�e���R���Y�.��[�Mj�L��qSi�����o�� f�)�-��'���~��~�!���me~����q��T�O��n��m���+ ��a.f����-�C6X�շ��:�1
ͽ��OJ����`'�&h��ot�/.\��B�ָ�3��4^�Y���ٝ0+�x�욫+G^^쭊$��ʑ5��E�ݩ�ŧ5e�^��+��g{�/I�{\p�ݚ�Oj�vAo,=���FB�w�C��~��G�~��+IEE�����C?	@�Q�4ʿ�������5;-<��!^�*�K�>ΧL%�zXf�W�l���K�:��!K����gWgD����܇�ls*�FY�VFKf�/�{����oّ��	��;��n3�6��N.�T�Yc�p0z�)�,yh���N2�9rd���܆�<��I����d�
D���?G}}b��o�Ǽ�Ӿ/�ϕ�A�ҫ�MLu�����y�hx�˦��[�ab��s�={��`\P��c#Ao���0hj�)�_{�����:!x�<5ݷꜲ5* ߂�#��h��uf�����qHLΧk;f{w!Y��\���
ъO�s�[.�:�yr�yUj�ji�2F丝}r+����=�������"��X����g�t}}p��׿���������z�Oܪ
���Q�������� ������>Gt@ � �@"�QN�0B�( DD���Q A�n���F �8J�D ��@"�z�U�  A*�����^@���  �U�e"F!F	EX%U`�U�UVUX%`�U�EV	X!Uz����@��  A"�����@ @��
�
�؂:��U�EVX$U`�U�VUX!U`�U�W��U�UVX$U`�U�UVUX U`��Q���@�J��yLu�E�$)@Q����w��5�_�??��?��#�r�ȏ�����O����￼x�X������������T�a�������UE~��"����?�?�=�a�$���~��?�
�����������o��@��#�� po��/�?���J� �P(Ƞ
0�� �,"*@�2�!(�@�  Bª�@��"���*�@�Ҋ�
��*�� ~��S
"��?���������(����"7��~}���?�����?����Q_���o�~���x���~��O����UE��j� �����{�Q_�PTW���A��� "�������*+�ß���?��v<c>�?�����������z�AQ_�#����������Oa��������O��C�����P��[�/��AQ_�?��*+�����x�~����1��������z�D��������a�=��${�����~�ϰ��EPTW�O�3���PTW_��������������d�MgC���!�f�A@��̟\� �Ͻ�"R�5E�
�B$�R%)"��R�٨��-Q!UB���6�&�6��P�RV����TP@U$��I
��UU��m�*d���Qe��6�h�[i������nP�lʥk5ZM�c)QKY��Y���JUN�XS5����-K&ѥk)���G���m�Y��kkl����ҭ���m��ki`%U)3e)���٦�-�Y�Y��-M�b�T��+6kY�%ZZ֙��������3n��m�6Z�Y��  ��c�Ui��]A��WZ��k�W���N�n�g�S��S^�z6�Ju�nn{���M�SZn�;Ei��ݷ����T���r�em�wJ�{���i��/V����u5�SX��ش|   ����CB�
lP�}����:a���C�СMhhhP���"G�
)�V����6�c����u�k]7�*����m(w�w{A^�5[:��uX톇<��eTW�򪽪#m6օ����=z��   >w�l:��Ì�X����on�{m�5J�u�koN�cJS���ޞ�V��G��[G�J������k��&�:���i��ۭ���ކK��Mm������m+a�E[h־   ��o�]7v�7^��K��:Y�r�^z�l#I�֕Ow'��-�v���Ք�����+҆ڽ۳�[�/jݨ=X �{�� GA�3
�)�����V��   �x���c@(f�Q��8�n�Ǘ�PX�� ��۔�]Ή3�T��4U:�4���`�3m��RZ/�  �x(�Z� -�;v�  l��4j�8[	F�[aCu�q�����h�5��;�����V� ����X�2�Z��F���W�  �=�j��Է  ��qVƍ3lAEP7/n ��wZ��4��硥���K��.U�U@ �=���l6�S=�z��)F�����a��   x`���z������Κj�:Ah:\ 
1��=z Qht r�3����
z� ��������l�6�cfյ���,l�o�  7u�@P �u�@ �}û t.9�M t=Wp��3�m�@t�m`  kzuƀ �pc�;{�{�(��Z����M������^�.mo�  ]��nàܼ�4�@z��pJP�{^���({�OxN�L����z^�� =�w �pz�N��/{@҇�Oh�*��h�B)�IIU ��F�OɒyUR4b  ���R����z@)*P&R�0��@ j~���/����������'�׬]#�?9CP�!���y�q�3�=6x���}�}��m�{�����x������`�cc���������c �m����Lc`�������y������R��&R���\c�e0�Ҕ+�Ы\��f�.ŝjR9w���X64R{&i[�B�9Q+6͗iv�]AvP���ҍҙ�6c�Kp'�dhBI�K�[�]���0o��L=Y!&��R��w�5�2�wVol8��� �.=ݽx�@[n���.���c����d-�H4�m<F]ثZz��T��5�Dq���n1z��X�� uRU,Pѐ�D[up��1��Jt3r*I�qYI�H`�Ԃ�#����6�ʷw��-�����1���Ϋl@�%D��y���y�Yx36�hb��8�5[-�@&DQq
��*�S�Ìbܠte3&�F�2�ɯFb2=V���� -⵹��$���Xu��myln����NS$O�''�ٙĥA�Z��%�l��e���*��ɸ��a��Ģ�c-(N������E�&��CD��i�	ˬ�N�M�3m\d �Nfkڔ%���)P4�2��n�C�.�C�=ݓA�,U�r���p��6���/B�kku�0X�J�;�W�{r,�ͬ l�t��t]
�Z&���t̺3p-#s�{:�gx^$����x�l$�BQ�X�3�0�GZ��0!V�;ؤ5fT��	L�/4ҬZ!�fx��T�� .��f���n�mQN�djI`�j�Gkrk/ gp���@yH*CwrҌ�X)���]4Q�ov]�u��l��ŋt൪��F���� {IIn�X�ު�طCE��
�.�2՗�A��Y�Y���� 8����NtM2���,�hLe5Zbt��Ʀ顖�
Fݖ�e�{�U��FAȩm�5�)D��JOl+��{r���67�m��
{�ա������2��Z�e�ē/.��D�/M;�kF0����!�~Ų���VWL��'f`=H�j;M
{�yj�V�)8RM�kyPe�˳zjLy�mV���.���gU�-¬D]���`�QT'G�X#2��n
�F��}��ȩ]ݳ)
kb��Zfd�v0u��'��q�4)BƨS�N�n�WR��`	����^Z�A��m�Y�f%�R�y1%u$��l�c�ܙ�(/�K[օa$]���n�G��gK��­����b,����v��i�n
z��6#`MI�)�on�!�_&����2� jR�.7����+V vw)�(j���0ވ���v�mbXQ��ZƘ��ݩX0���+�I=�m�+Z^��h�i�%\4v�9�l��b�U�+)`�2ŋظs��oa͡�oX;$�R�8leQ��Rv25�kɧG�r�f����s%H椷��#یa ��b'���.�A�S�7ywX.�32:����Hm<�J�Ѫ����vj0	���e��) ��3�v(.�E:�`��K�Y���ֽ�]��E/ ��GP�NiWV����o6P�A�fB��
yG^m-UȃNcn�(G76�k!$ˇ2��,���OX
D�%A�3%G&�A@F�c�#[Bm�T`��ә�\��Ҳ"�p��1G@`�y;{r­!4�����)��VV`.�4Z�� <�J'���:iM<ǂZSE�խwk�kf	;L�ܵ�{��Z�z̭gl��MXٲ]�=S�lɺSR"kF;X�;���sU���j
hj�oPT�f2�T����� Q�ͭKXX��X���P�W�.!�F���.n�Ҷ%ir�Y�k+&��:%K0k��U���B��en1�°�-����$���Q�0��I����H�T��-b����[5V@�VE�IA�m�ug)f����|g�r���ϐ�op�2)�-X��Ii���Mnn�f:�`3,̆�����j��(ګ`'����1�xHB��͔.�zFV���rmՀ�[R}�5r�ֵ�j�7CN�-Y�ղV�Ђ�ϱ�W�Il��D\V%p�CF��ՓJ�x)��Q� ����۫Z��-�4Iؐ�;��!бJ)��+2��V+���h\cY�nҺMң��UeV�G�x��K2]E`oV]��6��՘��5ܸ����r�nj2'���0�ƣ9"�N�V�2�qI�k����\@n�_x	b+	�6oc�V�j��V���a�Ԭ��^��l1&lF�br�h�xH������P:[Kf�
EOj�(	q6�F��P�Wz�Q���"�h�8�F��x�N�c@��5B��a��Qn=��B��f�ne��]���ڒ���!v力K���k2�������;L�ѰL�,U��{|�¸Y#'�������fJ�i�b�ӱx4�L��n-��R�q�B�t�,Clt�XnҳD!$��� b2�õqS�fZ��R?RH:߱:sS/jIZ��V@/&��YyV�ީ��
�`ɲD.l����XŜ��d�@m�k�P�29�����ڈ�u��%�x��q"�ni���(.��%�f �D
�M*WW�i���V͚�#�J-�*��-K��I�x�������(���d�F���4�ЍZB�\��U�jgVN����fq�rZ� �*��BE���w$�m�t��`�p5"�hgF+���'�5�_�7�@آRd�ǳɸs��n>�jI(^�6�)�cW47�ǭJ�m�	Y��f�V�l��Ub7�W@�Km3�i�Wy}5�;��e5Q�J�B{*�f����c�U�7^S��l�Ŏ�.Y ����Ji����t+M�7S�)2��r��4l�L���ֈ$졓l˺�mS1�qS�b���or7jn�����W�G&�7���욟1)�Y�"��F�4�ۖ����m�Z�%�P#$�б`X�pR�V[,Ve���hԺ[�Z����KP�x�'��ٕ��Yh����^YQ�{u4��,m D�8�0$����VY�Ms��@4+Ej�m�kPXʤ��*��nc�"�B�[��v6�
uk㢍:�-�û�6�Mm�o0L%�E�>�ckMl�R�.f6S2 �yB����oV�˽�y-&Y�(/�-6pa�D(�F�	ɓs5;JC�Zy**�ʤ�~Z՗H]�l�^�%ǀ+(�7[N�CKUVby5�I�P�r�JOM�d��E�Ǘt��X�n����u�KX�3��:�q����;�J�v�ҕ����'R���X����YwN�pP.j���{9��SHݔv�4s#p=8h��y2�l�e��-��!�jE�h�s]�S��P�ZI�\�azi�#�	�%�S1Q-k��Ͷ��6"�;��h�K>ȡ&��U���.-��2��6jcBe�*=�}��Y(����i"�G�ͼ�)@���D0y �x1���$�Cɂ�8{�I(D��Y�C"c7 �7M8KڏiZ�s� VU��Q[b��� �a�l��31-�2�_M��sY� kz�cjՆ6Pu��"2V:�+]D�V�BʕU�#)��]C�U�e�d�ň����k���L�gg6�{�'#�ptiaR��9���X���;h�oAJ���^�7�-̦���ժIGE�r��;�ɭ��+/%�,,t �C��L@t��PV�ٕn�+��=�r��AU5��8Pn��c��K�N�{�&aSI��+6ܳ�-�+yY �tfۚ�"��I��N�L-��7f�5�[;`m�N4ͬx�*G6��w�k�ث�+mQGi���I_�	�٤�/%��)]Tnb�2 �}�N��!`T�3�7��G`yp�ǡbKwY,ͩ��o�kp�56����[��U�Y�^�V�AX+*T�X���b=B��
�\������^c�+Az�������U���9V�iCQ�\�Z�f+8��H��V��9�p��8�2�6J<פ*'�JaM��ER�Y:a����[6|�n�(��MCh��̧f%&e�6���J��Y@��+@��������(�j�>r��BͅV����o+*[WR�5�8�h@a^�Y�t$ٍ��mսZ27��lX��Ec"����R�Q��-}C$$L7�Ws-\4蛸�ɨ�
;[��D굵y�n�*�g��;���l�I��Ì�B�����h�,��ֲrGIV����=̊c�{sJ�"���b��t��u��;��)K-u5$�C78����g�5�Wld�өoP#��ޭ��w��n֩�X]�4��v�<G����#M��E�'x��(�56�)e�.�p��{��ֹV��)��-7Iϓ/r���[ˡZ��	[w�f`L�	7l���WH<�0� �$�H�1mXe;i���+�snh_,�m=�`��ˣ���ۥ�K6�*ha�ߋֆ���,��ciR�.E�R2����O(S�itwQ?���ՠ�e��s�+c�[�`���jb2��v���_)f]i+]�(�1`*��J��!9Q�kF����җ��yG#k�w��^n���oQ�qv�NB�s�"��si��"�7fա76��aT��2GF[�h͊Ōin<M�ܶ��f�QT<YA�2CZtL*z q���� 9����n�;X�XkJ�;Z���I�SFD��e����;��˿��d�B*�ݪV�dV��2�1ކc�o��2!PI��m���!��d���X��r�bF�ƄE%���y�vd&��|3^LB�r��R,�t7N�
�Ǵ	kA�YB�̵wt�:�
�R�S$[�=N]U����ʔ��UhCt�I��{J��J��\+O�In��VRܿ��67l�z���Jfa׵V��}ksoH��Am�㥖�ʔɼ������T���[En�d`�3/qX���(|*���P�,�P�ҙ�6�2��0�Z)�.�QoL�zqKwt	�༚�z���	D��S�a*����0����G`��%o�N��r�6 �]ݚ�q7R�a��q<2S�i:֢�-�t��P�H3�YOx΍*�
5��h�YM��y��4m�pC�6�	n ջ���m�j������Q�B !O�n�ݘm�qV;�uj��`ʓ 7R��k�t��2�
l�b������0�(b(;h�v�T�T�&[��f�%���`
9��+�yBࣩ�zr�P�l��!Z3Q��[��6&�f%G30=E)�[�֫�b�~�M�0c�e��.onh�����jZ�%�I���X
�=�m6��ȫo
���X��"�^�2ԣv�k��ʵ@R�v�%��<���9z�$��
�����8w~����M ������y��;Qܫ�w
K�Oi�`�
YO̛�J�%����4�v�2�-�4�ˈ5Ge�	�V���ܹ��f�<��2f���i�y�@�U�&��h]шV�*��wA��l��7PJ���Rx¶F�ڦ�Ey��k��p�ST��06i���2F�:������.����2��w�ʲ�˙�$S��B=*g*ٽb��D��eM��tokw0ŐI�r�dCB̈������e�c)�e.��Fv�SǪ㠦�gؑo/4-6%�NTH�x�+'y��݇�|}WBr�1�ZH�dg���]n��&%���n��6�P��w.#0��0RH]K��$��]�b��llb�-��,V�rm����hz�^���e�ŎԵJ�$�ɸ(�u.'��V��T��/fVj�lJ�H�b:s&�F�!�q�wu�PIHkE��U�� d	��*@�Pϖ;��GXn����7��7.��g�� ���x�˥��>!�z���,���[K"�8�}y
Rح���ohi� �!��3��j+ 3h�_P4�L�o��L1^���1������]�%���H]*kw6b��)�*��[�(�lx�L�if����V1��B�f��,U����EY�q��\�6JAz,��rG*���ub^Tٸ ���TtX)r��`Ӑ��@�Yy�PwC>{�t,bڎ���AZ7\�Yf:,�gJ�'v�ҴX%��ę	̣�h������,�K5��T�I[�����lf��i;�*���4Z7�l�Ֆ�Kw*v�v��}Z��c����Lӥ�id��cLd5�a�S(�6.�	�b�6ȭ��t���&��X ̐j�O�3jx�G,��R�Fh5��V;�c+sZwtU	hh7Z����l�KM[ۈ��$�����R�K/7���x�d#1ݪtm�j�7� « ʱiE���C-"+["Ȍ�-`���f�
܆!�Gx�G�e���ڼ�O���[�"�U�x]���ĥ\%��1�������2�J��z*(��Qů,��`S�-�5�X �Qf­uA�,�$���0j�+[� WtO�KW]J��Ai[ʎ-��S�u�cN{���>�c�=�I{��"聧ʗ��J6򮮵��7)�7& @kp�v����k(�����2�ۭ5wikE�2@M�����m�*�`�����ԡbK5T��P�7%�U��A)�W��F�Pj�.�r��ܷI`d�f�3R%2�Kv���9l~jc�!�q�	��)8^��s��J�lۤ��5��S,���e:d�^��FCD���m�����D޷o=L�*�۸R�j]�C�v��`�$Gm��������e�cvj��VQ�ZT[>TUeM���[�Եn�n���.�
܅�K2�J$�.�{�;ui"�y�H�
:6R�V���|ei����X�mH�5�V�D��є2��Gt��)@��W@U�8����}*`�U�$�K2Ոť�����nÛ����F'�FT�{����WAP9P�Nz����a5���[<��t6i	��%f>�`�r���9U4���n��	'��'���9�ҁ�ɣ<Y�.�&����~6��is�v��o�)Y���y�_����ô~�`~����W�Vpog%�A������*���?�G��p��X�5�S�t���҄�i��R�r��>�9���*�׋��8�"� <R�ŭ���ѿ�!�Y-f�J�7}s2�j�5|�]����YI������ќ�i[J۾$�JEI�6����9�͊eŕ�D�!����p�i�7��S�=������>F�eߛ�>������ԟ��n\O���5a� ���x�'NR.�v��ӡvM����e`Du\2+�����wFK����>�ٯwPM�w�_)��o���=��4!��,#�־ch۴�k�D���^���Mx{-���V��1�v:��<y�,N5�$�.Y��«�xbŤ�p�y�g-��5!�Q�O�]�5��
]���aѢ>[��N3�_�lW2*毁u$��K���#�Ѧh�P$�zT85.�����'��M=6bY�,�[#/�Y
}�VU�7e7�7m�]�*-�5��֗]򡎗o�ǚʨі��ʳ7;}��qDv]�D�^[�[�_�$�s+em��;�6��T�Z���Y���K9µ��9���ܷ+���m�[�.�v^���)�ړx�L6��cJe]�t�M�m�e���j=����Z�G�X��G�\�lt�c�<�W����_���	�=Ė{�#��*�r�LWv�њ�i�fez�D���͛m��깠�SDL����RԹ^\�����..
6�5���z�Ĺw"�G[�(�W>Re��ڱ��a֒��ǋ���{v'�,�ܮ&΢x��7�1�B����n���w+W�_1��\7q��J���d��=)�n)��&��%�����Lu.�!����qyQ�� �����Oɑ�nefl�쇦�M<��p����u���7����(�c��z]@�:��=��qU�Wr�oR��,�a�.[��ٍѢvڶ���v�R�������,�1��3�u7K�\�ʕG0s,���9%���X܊7j��K����9pZ �)�U��bY�fE��i�Ou)X(=���;^�����V��u��u;�������#+u��t�@��RT��m���GSi����4:���.w��q���ӽ�$b��i�����v�'e,H�wH�`�[���cꀳIHgx��N��_�]��iJ���4^Cb�&i�x���:w�r�)�nQ���9$Փ|�hn�`m��BчJj�G=�3����8�a���F�[)�j��ى^�ǚȡ�:Y��i��f^�3VoS���u��;b��o5��u:�7r�T�ఇPY�2�w+֝ZѴwL�*b}Z�����n��x.6ήT���F�6$�#�w'o������޵���S'y�!����!�
ŗh����p�+�����U*�3�uE*�Yu�R4�^=�m�p:j«p��nk����ΈG����H��u�v^4�d�l�/ ����W2�=��ڃ�����(_��:P��%��#��9
m��ʍ�]�w�P�/�N��9\-EӶ����,J�|�b6���KY�s3A�5���#��v:�kX���2���[�}���iu�b��"��r�q��d�j�Z��h:�+�|�:�o���4�5��(�F>��.���lXN��������_uK�h���o\�Ǧ�\�y(�Vv'��i2�s	_�9��ԙ#eZ����ܸz���nw9��Rޞ�=\h^֩�y޶�vL���ה��!'����*���o���fk`|�;��J,�8��ب�g��lp�M;ˣh�B+n0�W�)^��& �?�ak����mr�����|�	�;x�{��/�pQ���[�����/��DZ��7��'��ܞ�j���t鉛�m�Z<�PW\y%�y}��1�\�+2�/��r�ex�.�Nn:�i�ժ"��0
���5�(��Ū��f�ͷjU[��A�e{<��� ���z0k�@3u[�����N�op����1��_žL��
w���k�sl�b�"Z���yNu�n�R4`���������n�+�ۆ��9�Z��0�l�Ӟz�i��q�4�Ԙ�RTw�_g����+���| �M����F����cx�9&HQ�3�N�.�m��]���3i%�+\��{�1���e^c�Qd���Wm�ܨ�⑞��ϼ2�;��� k}�G�tqK��YC�ov�������y9����ޭ��ϣ���ڰەX�U�&�|�x��r�of�4�޵g�V6�*�9�"a��LM�Q���O��<.��6�u�(��F�<�a\;�l[{�w��������NӍA�rod6���^��ؼRv�"�@���&[����xHBK�Z�o�F�r3���~h�yBv�TQL�	��wa$�8�r�љh�i�������b]�ůa���7rz���w��r���a��Z� P� \,�fGF
V�9���c ������$A�9��Uu�+Z�ϜǏB�ٕ(���"e#ݾ��l^�,�
%��^����r����Ǜ���zxe��� ��]��3@���v�
�V�RF��p���4�,[��.��Y��ԗ�&az�F���Rm���X9mr�#�7ټ�zm	G#�g��(1t��E�=�lt�g)\���\��bx��N��޴sg3�������T�n�==��~��弴D�}�X9k�Vs��O��1X��ދ���������c����h�����ҕsq���q�����1�b�v7��g2.wP����oS�+���ND)av�yH��ԪI!m=�ǀ�� ��6͗{�;�Q��-b^l�A74JDm17nق�8���S����=��}�_��|���gǂ�t��Çϯ���ӌ]�Dj��/cKf)�U�-�zɭ\��hB���&��,+ӳd�Nj}��/��.�P�?0��.�ޭ���T�Z��˿����\j�}o��F�؈y�(Pnu�Y�k7i�u5A�

[@nu���}��G$�r�>����4���+�e��$3���� M0���U�e�=<�$K�4��8�A�k>&����S��zuc�!"���.B"V���U�;uu��KTk�7�T���kuG��vv��Dԥ.c���f^U���3����v&�a���֍��.����g�I�g`�����:�� Y�&����d�g������ `Y:�V�yMnj�:8]B*�ц��Q0���H!2r��w��.�:Q��웝ʮM���'X�/0Tj�gK���hz(̵S�GK��� J�D��ԝ�����@Z����-E|h�^u�w���2dw�f��w+ޭX���wq|�M��,c47í�./n�sr��+��J8��z4pq���]���M�g��'�+��6^&zj�ºR;A5B�[��oi�	�P�9w["�U�堑̗h$���R@]�����f�}`���1y�q T�Z�1��^�>u�u��X�̡I���<�έ ��s�>p��S늬�y���.��q�8�������N��F�
-��h����$vf�Y����>ȷ�,���"rށD!��g�З4:��Qw���0��ڣ�C	����7�a���d���xd�\x���Q��x!�>nCט�Y"ǯ�$�sa9ٝ$m>̽v��hX�.�Y]+�`LJk�f=ξ�O��yI�������9Zul̍�f���Ek���ʁ.�7��ni�M<�[��E6��ptOZ�K}��dMq���c5��,Af=A����x"�44�7F�f)kZ��*,���WiY+�zLk�M�3=���!��ꕭ{�Y�ѺF����VDk0�d0�n�;6��|��d}u���&�ީ�Bg,X���<��:}�サr_:g�|l��s����1�!\���jjpa�I�`tG��n1�����j��%\�����
-'h)����A�����Ӂ�\+�qt�v1,|Ͳ�C�mb�-=&Э;�yz����fG:�d���#�{
�Ӈ����q �U��D�G5�`��x�ޑME�1+]BÏ�O}3x���01�2,���`ͣQ�����#�w۹���ov�Cc���b�	���m˭;��\��T�@���wV��w�k<�֗`w�E�M����wH��¯��������>\*&�>Ē1��g�l�g����-�Ŗ�C��﮹����5�gK�LE���yEX;)�#Ѭk���o��b�(�j~����%�;�?g ��n>>� 䎝0L�kB��R�Rs1�V�<�HA�a��Hܠ��4x"����[Y�D#=ނ�w=n���qw�ݾ�Q3.ӣя�R{÷U��vvd���ff<��>Y�+"�Mm���p�C����.�w�o��(�
�ƣ����!vn�;1-.ɩ�(%`;Ժ0�
z�)`˵[`��bT�RvЋ9WN��za��;�B��T����f-�r� �2����7�I���d��w0_P�E��c�=��U���/-�����˚L��՛h?Iw��hV4^T��^�hk��f�o��tc�%`5��
�I��x'_v��P��_9�I㾈d�����Od�X����;ש���]�X�Ŭf���/�:�-�/�e�JܥI���q���^�W�z���ު��@�����y�Ν����-4��o!�W���5��|we�x�لK�7q^��}�s�a�C"�)0ړ-h��Y$�PWE�Ԇ��,ٷ��N����/�T���~�f�ۇ8�����"�6 ��/C�k�e���R�����~(+�H�z�#{o�z�e;�JO�D��Ú�˺³��ZJ|q3c�>ј(T�M�T�!�|_7}��&^'A����Օ��a�*��}݊;�:H7�1m��T��zz��<���yp{-�ٕq'O�\��VK.���.�t�+�Y9<�:��|�x_T�Df��x�]�;���Ǥ��+���j�)x�˛�R�]\�gp� �v���\�\�֥�w�	w�m�&{˳�ͫ�Xu�)0Q��Uݙ�XV��w�L0uۍ5Թ��_t]�YZ9s��Xåx���i��ֱeu�oY�)v��،\#�u#�r�[b��(��������e
�s<��i�]�K��^��)F1�=*v���'MMh�].�R�8{g(D[=�6�9V1����۸�!�ѧ��#uy�k�>�Q@^�m����\�^�A
�J��DJv:u|��6=�<�{�i)�r�LV�W[�Y�N�d�a㙼�a�.e�|e5x/��f�V�z�YpT�Vu3���x
f�vG�mKӫy�J���4z�݌�k3V=��/l�g��}�s^���U��;���W�E�E[4#�g9��vw��e9s����ä'3_	\��J�,-*����^���P�ݶ00:��M[z�0�.�HҊ�"r\�ю�&�[�
��+2��J��R� ��!c��y ^fzU�:�\O�&�~샅-qvq4&�L�{t��Z'��{�YW���՞�[E����e�d�W��r7��]oʺ��e�W7�R�g�Q��^u����>/�WQ\���j+/ YÏm�c:�eR��E�̀�mZ䌱b�*�&��:�6��_LԬ1���;e�s	m�ޔon.?@)���4
�sWg[�w��7̥��[<�	�@g�e�7`��c�[�(q��4�#.����A�y@9s�V��7���P��{i�Wڦx�S������;sd]>�o{=�F�f�k���S���w֋G�u��y�%K��jj�.��-�p���;R5���o|�pڙB���pd66h�^�`����.�+wؠ�w/���[��>�I�AZ���O�7;���yc�h�Ry�G�� Y�2p���ҹV4�9/m��k� Ox��#�ZR�Y]W���z є0T�� �L)%Q�K<����Q� �]>![i5[�T��M���8C��EG�[���=�8��,8h��N�e�9�_='%]�	r�4l�s�#6T�*�uu���8Xy�eg�;�f��<����tZi�cAإ���k�������	��a�]&"�T��f�R�,lHsma��X�.
|RED�9ҹ����ص��_��KZ���ǈ]ݛ�f�VKe�G��a�YJl%�^Ȋ�rX�	�ax-kfRd��(�H��n]	ǲ��W��pP���k�<)1|��q)8P�VY��2Ā�}���/j�������,t����
p �Iwޙ�#�0�N�9+��n�����&=�)�slv�ʹ��l�3i �;k�J�mi�q�jsCҶzf�v9(�Oe�SU�
���	-U����J�wEe�kWX�;"��۬��:�K�����L�\h���<����d}�;���Gu��|;�@�y}��2y-�n��s��.�\��D��u�����������EI�tv�bo.�'0��p\ɦ2�ٻH�s�h�������/��R��v=d�o������Ε��n
�53$f��-�3�����Zu��l3�U����4\7xk�2M6�r��tR����YQ���u��N�tJ��`A�,i�EHcn��U-B�I +���^�:u�۝�!�w�OW�G���ޏ����+��Fu�Z�+n��Ed�zL�KG��]����/v�;�־=�����矟�>��`�cc��o^�y��(���o3?n3�!���jq�w���b�
���D��[����aX��_u�IV/X*�)Fղ]��vu�1���-��q��nA��v�h��:���t��6�����n�(����e FY@0�%���d����I��.��D�k�G�ڙ�3X�����!{A�ˁ.�v�/jB�'0S���Y���#�1_A��w]ns�A��N������Ӽ��s��n�d�%,�ӎ��v�|n6�t����qv��Ա���$�������;�����w�5�z���S*��N-n��G�6y�*��YL�&T�`9�K@������r�&ң�ʿ�2��3mqg�oiF�4�g؀A���F��,^�mҕ�
���w���&P,������"Q�z,1��C�����;�)tD`\ }ݽ�W�&�u5o#�]n�ÕW�m�<�ǹ$O]RS|���^��;P�B�Բ�Ō'y��ϭr������J���@G��-�ٽ=xn��˞�$�#w���6u�/���@��È��/�.r���A��H���B�nb{�#���U.��h���)�ލ׍�3G.o'u��ZwJ�F��X�3z㙰SH(��+?]�Z[���s�04�:�h���,�����ӵ���8v����pޮh��/��| #�6\��,��Ge.�ORg:�3Թ<L��p摮ͭ�	J:��x㿆Q��^�7D[Ok��Od�Xo,�I���8�/�١���4�I^���N�ע�V�N2f�扖 Gi(�ة4�jE��՗�E�)e�Vo��2��A����۹�
����뷈.��2����YA�q��45h๗c( @}K/ON�b� �;4��U	�d.ݧi�m��hd��������q���㮚�w�y�ާ����^�g��f�0'��oh֫�C��n[P�Ñ�V��6v��r��kI�->�Hr�ʰ���no�SZ����9��4+D����a��V�۝w��Y ��F9v��;���Fd�2�JF�e��������e�R԰}��uu�_6���[�m��*ʧAn��b���� �v�=v���d�[/F"ʳ����򎨇�bv �s�m������p:C��ǭ�gܠ�U� �~��¦Jz�s�J�����p�ϫ�be;�˫�`�1�q��l1������)&�Z(޷�
В���v亰��2-q�9�N�ιՋ���1��Y��g6�й*���ɖq�Wץګ�0+â� ��.YOy_q��J�C�B����fi��B��û�hI�
�S��t+ֻ��ص�BYF�ߦ��{z�J�び5�s��o�v�^��-�<	�:���C�u�+�9��p���{���n�5��ۻ���׳F=)̔+�.��՗�u�# ���5��.���� �%-bX�Xp,��e!e�7q�h~���ʎ9Ծ�5�Bsb��obMZ��F��f���DN��o�uÓQf���n�k�;�µAJ��G��ڡ�6kX�an�7M��c�w��ZB�Ec���h�R����*��Ż{���K��^�+�b��Y��n�I�c�Ok��U7v�`N$�2����ٯf��.~ǀ{s��=U��dR|�i�IP+�
�\u9���Bغ��M\Q�lKﲯ8���`�[=A������#G��[�M�*��IFyr���6���{��X�ni����m#�dY\�O�b����r��v�[��)�L��փSI޾˽�WCn��}�|�"��~��E)�H{�%�O�Mn�T�y��t����(
T�ح�"#�nZ�0���3�3z�3�nu���Y�\��p�J�K�����k����Z.\�##��G¡�I\�u�]<� Z7�{SK�q�6��rx.�#�N��uĭ���Ց����W�����uv�(�[�"�9t)�7�ޖ�g��/an#.MkzV��^�n\��)x�:ל�
鳋��+��0�<+tǄ�-�/ү{�L܁p��ݹ�D�Z����wd�/"=G1!�7�Z)2X��)c� ]�<g�egsz���n�-���(���>��2, uj`Үo���ۓ1f�"�b�fm�ԓ.]��{����x�jX�-��M�wc6+�k-
�� �N	7�?�d��	�+S�O��0i-m�#��6��L�2�pYp5�a05���WO(��[�%-wW�+�N+ݗ�5E;)S�ڗGF��\���h�B�������f��Т�ˌFHǴ���[ݲ��t�7$oo�cJ�pv�V����(�szSD�{��%�	ќ{E��ԅ퇘���ڡI>�=��Rɮ���ݎ;����Bw{ڎ�m�B��Іg)�#�+3G=ܼx_�KQ"�ů��d�U�欬w������w��9���{�/i>���i {��kf�ӵ�ڸsRq��Ӕ���4Y��0�C�ra�嶓�qW]9��l,}U1n`�Il�$lLSӇ]V$	혼|�u�G��8�S�tOm��{A�<�yͺw�N�y�1vV�T�)��Sϴ�k�M4�f��w��5d>mX;+��p��;Fr�.�B�pǋ�>����ݮe�6�:	V�Lݸ%��!�R݊`�'ۓ*ڻr�Q�X���xhK���4'5�N��s��n��:��-c��e�k�-8��%�p�d��0θ��ąo^�쨞�!���	����F4�XZEj�X&ּ���MAAVi�l^��=NIܴƒ�&���1���r��j��4�k���9�_&E����j�۔�<,}��<����������e�~<_/3��ݗb���[i�hL�z�z�4$������pZq�s@��lL5r���Î>ZM��k��ɤ.2��Qc���W"а��w�J�Ŋ�Y��ƫ��u�y�y$�=������D�Ȱ;�	�7D�cSl$U�]VE��9�7.�U�:�3�9�Y����M�G�:�n��{��t�ACx��>1��`ʜu��r�1�w;x��K��=�
vG�Q!?M'+m�T��r����	내�h��3���P<l����X�ڑ��N��z;ob	u�������K%�?d��]h>�Wn|��^��G�A�r����a}�����]�6�����'��Sv�H�L�Z%<p=��9��i�leXG��V�4�����Ft};��Y�#��v��'m� ����N���ty	�ݛn��wR;ǓCc�m_*�b��BY��N��s���[8?(C�x>ypS��5�/�}����U�{��9
ۜ(�%s�*M���6�����яrei:�����MY�"BΉw��
榐���T�����ۗ�(dQ��U�׷Mu?bMy5��ͫ��o%<u���7��*�l��4��3j�Á�f�R41�S��e�H��G+w8H�>&���!���5�y��a�Y��J�cm�\�'r]i�7K��E�]K[�UŪ�V��D�1¯:1��]:zA�w{'Ν6�Y�']n�c�n�q��ea�zqqm��!�u��.ֵ����-S���Zï���崹&�e�#H٤�Oxo�z�nEr���xI>��R}��qRy���}' 1��'@ky�5�USJ��R�0v�c�@(]��wW:��R-�x�-$��"ػA[ �vԦw,�+3���h�u�.6�;Z���/�Y*�7���ύ�I��:f�@ζѺ�s���%�*ݨ�X!+u��tIKB����b�cwgs�ڭ!�x����&�������<�Gq�[�5VtPVoi�ƙz霬Y,3�i���`O7��E�V-㳅[{͒T<M?��	bWp��j�����7>#�jeB� �~��t�v�
�2
��5���T�G�f���l͋��q(K��Q+��?X����
#�^C4J����r���a���ԅ>˶��v�<q���;�>��6�V.�4�D�Q���	�)�Ւ�n��/]��D�`��5z�۰c�[#.��Ն���RB�C�η�^Rʓ�
*m7���j���\���D�h�9��ӱC{���g2����1����#�/�яF���s�Ő����Z��3x��֛�݆�x1�P��ۑ���{B�Yꗛ��z}ա�����ӂ�������4.����v��'](J��YΡSyU�4t�=4.���4MCE�|ϡ�G0�v����`嗶��+ئ��x�ƃ�q&�/�'��J��@ɏ�ݓ�[ 7z>�UQl�X�t,=f�ͻ����}o��t�#����K�*�Z:2��ntli�#.�vj�R�*h�"��t�G�aJH@�9CuH^և&��3�k݂��{�������m���.Po2)m�o[��ͨs��Q��pC��uj�	�<�p�,�j��o��B�%%���{��^'����Q���un6�-Ɣ�1b��]��qT�Ή�r�4���Z.��[���=�m� �E�Dn��
I4�Q��'dNַ0e��pn�7�ܨ#��={�<&L��XNQ�Z����^��v���o��5S;Ɇ�U�jr��I�~��vk� @���:(��l\��z�w�]|m6�J�2q�����T[JKOr�e��Ҥ�ul��g��Z-ê��s��솰Z�Θ�)`�t�oFT���e��v%O8SмT�PH�������{�1�R�djl��F���*-�,��L"p˒�4����-�P�łNVIC�cJ�6����C�݅V鷜���6���(��B�q�[�K(�;X^[NۮZ_��ç���a+�-�>b��j��Bw|b�Q��L�ͺ4\���xA>��W�t�ԅ�M���K��&���������dWz���	G<�*Ҍ�r�&論n95��1^P9�E���&A���J	C ��*����TUKB��U���X7j���tf7�<����5%�<�q#���6�(�8:�j�]�	������:|�{�<�TG�aR#IK����뱫\��J��9��	҆���WJ��ǔ]L��vQ]�bR����7��tk��4P��r���7��<�=�(��9g�@�Lbn�;7��I�Cx�S��wV��Pj(�3����*��2V�]d@dG w��<�k^@��T���;]�vYv�9I������9
QؼnܽYW���b����ܵ�\u8'1S��3k���f�ZU���U��H˗Y�C��E��n@�Qb���m���H9�� �[��˧��{�8�o	^�3Sjp��^,�S(*�4�zM��1�+��u�o%8:`tT;	�d+�i��ߗ4�xJDq�b�Xe��c�o){��>�e\����Zk�҉��+�u\�ܓͮ+e���[���R�G#x�r��Şӆ1C�V�=>��{9�~ ����P^<�[v,<����ݻ�^�ٸ��S@�����/c6�/t�ݎ��"f}!Z�&v��ZF���T��(+x�ݝg�&[���Dk��=۽FA1�w?UѾ@�p�-D�{e�oX.��S]�un�3����k�D\��b[Qm�"�Ĕ������6�vݠ�Q,���wr�&7�|�>p���i�+��mqG��Λ��>v�@u�ve�YU
��(aS��|U�N��B�8�x+�1S{�����ܧ8�D�}6Km`��o���6QU���
��I���K{�7k�؆�ǳ�`��.��<Yօn��3��8�z�m��"*yW��ܼsr`�m��)�\�8��6ަ+�Y`�\3|ީ��OJ�}t���Ca[7�9��i�}[R����V]0l]<p�U��3-
I�F�%Y�a��yR�5�ºӵ�i�Q� ]��8�U�Y��3�mt'���9�m����34���K�� w6�]����6^ݶ��ut��{D��5Ͷ��=/l���>��֥;ͮ���@��J�e�j�*�Yө��;���e܆���l>v;�=(J��w3F�Q*�ݙ��RJ���eȮ� �;���:`�����V��ۘ𛮂&tކg ���H.�����<����3��I���v���
�	'{N�3���ً(��[,�&9������0ҹ��:w�27�fE�9�/	�l(M�l`�zھ��]oV��b�f��5%�akvpF�k"�rH��5�&����d��^���>LB�Xӹ),}�{ք�ؠn��Ea�{��3or-��]~�*�Emk��qHV��oj�,|oT�{HpƋ��tw���ye�ʯψ�ϕ�:���ڐk't�k��݈�G$v��h:��D��YSf@�XE�l1XJ�)��;�$��,�&�)�n��c�`�CF��N���۽ʕ�e]����n�ӱ�V�KÃ�H��M�H�>����B��ps׈Rs�x�~�fX���s��3t䚵�d�0l|8sm����nk���}Bh�T�Ȥ��;ܞ(.��f���v^��o{$��a�H����g=�^���cNH��V�W�`P��]ܛ\z�mw¬u�Z!����[5��Ţ�2ه�]5Ҭ9��&�GJ���<��(�j��BP�����,�V�l��_ ;.�&qj36���v�2"qw��qpS��4/B�OAh��Դjӿ]�W��r�F�%b��I���\�2���;�]u�ɊYX��șAB���a�h���SC뇫�C�u�1�U�ݻ��l�����e�GܕAc����������>/�U��~;˕%aM(gte�6[-�������s;tR�{B2�4�՜����u �E�}S�������1kJo�|�oy���z=���ұ�̭��t�=���"��5d��GI��w��f=�=��ˋN�4\���mNN1�E�z�3��U�ޝ�9%y�j�PFv�N�Vr�^���� +���nRh�W4���
N�*̦��Gᇎ����G��1�㮯$�{gG}��q�z���H,�-|���ܹ��A\U���@�����6��Owv�y4+缧�|�u��;�Oex��tn�~�揭�r���I^�B���G���2�7��׭k�S�޴S�Au=��Cר�7�Kh&�y*̈`5k���n��9ZR+��w�Wĕ��Fl�D&�,C�	��+�y8֮�{�ѱ��
��
1:�Q̞�=��<�Ӈ����� �}�����.��=��M)�yVà\ܯ����|��38"�NϢ���ںM=s;fpfq�z��ͺðvC�ʞҴ�����Xޔ�ɓ<��ǥ]���`�:��$\-�ۏY���a�z��ld��E���^8��	�l�n[zV�� =
�U�˅�#e���-�&��lЌ�4a������TF���#����	�g�U��J�	[����4˻��nt��^mh# u�d�I\�gU�a�.�6�>u#F�E9ڇwnQ�ˍ���?�ud+�.�J�#~3s��L�ջ�����,�;�<��q+��7�Ë��}���ˈ��,�+��@Q���"������/wrXUW-\�i�k*T�/wr��7R���\��;�;5Î���(*�.���8��.��y�����u��w.N�Zh8���u�/n◬�<���+%�Ownܤ�s�p�=��ܜ��2O2N�H�������ܜΞy&y����!��k������^�N��x����t(�rG������,����u�p��<�/���]�G7'5�"'u/G<�<7r�C�W'"��Iʷp�MBw]�\�+2�ʭwiX{��T{��I�&Z*n{wu���=ܗwc���.{=k�,���su���*����蜝GQw�rMW=����<֡��:3 Y9��3t=t���̊�NR'3�5�.b���U�U�Kqu,L̯R���#�Ү�wwu]C��(�4N���-1BF���I ��{�z�����Pn��Yҷr��:ã����9a��6L�UY��w:Hh%��Ri����o�Nd
�]�I��ř��M�hC���g�b�&cn*�C�c�b�����hA�B��`��x�+�}j�d5���Gד8	�>�6��p�>2P�p�U�R8n�=.R�Q]�i�^-0�﻽�y����F��ZW(�
�F.V~�����@#���.1�u��i�A'�ևq��z�U�Ǖ�s�:���#�@F؅.�keR��}��+�फ��u���������V�o���;ߝxT�W�/��ݺ�zi߭�<(	f�fJ�rej��=P%��#�^���n�T�h�3X^*uby��lv������TKPf��d��M�
U{�����+�8+�/����l}�H�EI�=m�wN�U�#�yd�o��z���G��й�p�G|]��X��j*D�a+!i����bҧ��g�L���ڐWdε�;�a�
@uJf����-L9���LT7�xz�7{���iVv�SN0�"4��=������+��_���u�@�D������t��C��x'�,�u�p�]��vV��S��sPc��֜�+n�ӿO{��O��A��jK/զ�ݦO����qO3�Kb��Lu8BS3��>�d�m���*��t!'�h��f�}}q{SXx�� N���fڨѾ��*b�u�gB	�}};�f�����5c��[r{��C���s�?k�:�P���p͵��*���{X���"aX�Q.�H���2W�N{a;$����c�j���7w�)���o���6&f�5�ʃ/�!�Y� OIMZ��n���%JA�J+����c����F���yp!��ﴏ�6�AY+tȯnϹ��Hk�Mȭ��VͤpK�qE�q�;v�����7ȧZ���#�]_#��8X,u��&��;3bܬNb�sƨ�9ٜO��F��,7s%��s$�X+Uq����N���#�?���_A�0P1�]�:�ΘjW,�=�nC�q楶���:5{�{������J+�m
��2��ʄnl"�p\�ʚZPXKSPBka��t��jVb���ŏ	�o?m��.���o��W58^�h/���p=>�5=|��ѽ �C>�ZB����OH�6�d���9S�l'e�ƪ�jhnt�2��."׼��&���;�Oڰ.�M�?j�dT5��o���Nvu��׼Mﭦ���Wϓ�&�-'%`U��{��xZ,��C�*�d�<�f�����JX���'�pYNC�y%�z�ʚPkiS�%a���=y����3]~�_�N��ܽ<&,㖛��$��� /�@��O4�JQ���Mfk�Xu��rM�l}�;�1Rw'ԧ<1>�ع+�M��;��_�b�i���\��ˢ������W�gS����G%���u;��5�U��e�p���޸k�.�>ڗ�^
���T e�D�t���uMn�7��Egv���I��GnD��	�akǟvGƞ�-� �<!������~݃�ۀ����<7�mxʮ��N�9㟹å8��C�5�̋c�9d�['	˳�*�v��H��u�+q'�cU�]����59�*s��^�B7�J���CC�I�rKm/L��5�hs�s��f�%|L�)��V�r+")��8[#����	�<��Zu�V�lO��~K�_ܑ��������y�N]��<U���YDٞ]�1����[�uG���v��ؐg�-�A��x�i�B�-��Ҫ��ͻ�F�"���Z�c�0)���.�bÔc�+ٚUj��LO	?v<�0��[���ǵ��}�m�MK��=�3�>�Լ�Fn�Yi్�G<W�5Od ��ն9�<Y���[q#�˫� �<GC�XA���䭽�t�^�T	{�r�r�ނz���U�k([��M���V��](�T~MV�f{�弎d��{����z�Ԝ�O,��#v[y����n��]7��́]�Ԯ�qY�� �L��N�a�DR�'	�����=c���p�X������t�p�����9-���y{P�ޅ��<���y�*>����k*J���=�P�]z/�C�vj'oi�UN`�w,Y�v����/Zg��vc5f
#-�+�Vt�`��3㙵ƳQ�Cr�ҳJgx�0����kt�=p�et�N���d�8J�HdCYp�W߮`{�Q��6i�B?iܘn���I�4��}6��\s6N�En+3*���ss�vBk>8k8|�FΗCFĸ[�%���!R���#+$�}�9��T��/�J���r�D9��aHp��`Yݑ
�ђ4_�
a��b(L"Hy��&}�tJ^Ո� �v\�{M�������Bt�:�̳�+�g��Q��u[��w!V�;�3�j���0�8J�޿*l��Ϥ�Z}��=J�.}~`vŲn.~f���;�=����F�S;�h�ov�-s��3nL��u}�+z��e�%ݤ�G�OWM�N#�����3���N�@juH�k²�tY��uYI�y�1J���Z���j� 8�H��Z̀���\��?�(=V��u����i�?c[E�b��$�圕�����ͬv8U��|
!�Qԙ����@m�.HŮ�o�.`� �Gl����̩r����\z�o�ܾ����;A9������m��ݭ�qU�X�!��a:����xZ-�jN;c;�ˠt�cϺOb��F��e6i-A��#��h���7� ��f-7p7>wlT�Ud/h���f-�q%���{�!�����sڅ9y�d}�r�Z6pbdC��*WS<���1��=5�gQ�iW	��zPYf�8<��E�iL����u.a�W�V�{�����*NXB��M��K��S��g,��"���P�7��'�䶯,0�
a�e^���{�Yn�
��~���tظ2��)K��FY��[�im��´�J��x���+Z��;6=�[��4߷�>V2��6���^D}�a�۴X����6���p�`0r��şdB���N�vX]�Y�G�8)��`��R�,깺p٭'pƥe)̛qWo�L74ڙ��Z�s���9�C�N�I�7�Eƽ���,j����ݓڢgK�Tl�Ơ��9��4Z��;0�z#��N�O>���c�G����	�z�MǬ�%���Ԫ�cy���+ut��t�Q�e��n�iWM�2�s��߷n^��ld�h"b��$�� �<��>���gL�8M�E��y�ռ}��§�vd�C�����V�����W�����m�$�j�7�\to_;�T���?�=�^�^v�9�)�v�k�S��4�&����w��3K^�iգ�bݷ��_�?�ۑ�r��'	���S���T�/�K2����@m���p�WS�z�s�Mt�p�{�)�|�$%H�"�L�5`婇3G~+��b]��CTVh���Op��-�#`����=�� ����� x"xY����m7��me�Z+r��RU�Ư'�8 ;{���0�^[�ʸW?�G�T�[\�V����e�����aX����U���1.vd��6���^u9�N�#[�V�Ed��v�.k�Y�ކ��t�,&�-��f�Z=�_j������2� "�k��b�����N��*��ٹ 8�[3oE_�èg=�Ahsmt�q���{�T5��tSU��$nr;�����{�H{�0J� �5q5@w����|{�,m�!��v �;9|��K���(H���������*V���a7s%���"0��b���C�����X��Ϸ�U��*Z�:6LØo[si�f����&ӢQ�FL�/R��:k��f��C���8����0e?z�srt[�"�w<�,�H\���l���QuqR���6d���ݞ�w��ԝ30Rս��ͬ�%cC��9pǲ���W9��v
ͤ1΄V�G�%N�O�,��V�9���Y�Ry�F�3_:6J�^��ʬ4���s}S(j�Ok�#��<�v.��5
]�Bѳ��##�������8U�����0���u�m�ܼ�y�c��hUX��a��*A�<Nd����ٯ_ɺ�8`3>�� y~p�"�9
��	��6*���'�VC��W�Y�w,��uC+��_���"R`!2�g���ڑ���+nnTO^g3�Ϗ\�_ ��ՙ�[	�#W�<O��K��+l�����Q	�~��8�-l��-Zw*gX�&臹���vC�3Q�YCg# "�2�j�V���m�S���E�q��}��b�5;�g���XX	�<��E�:`v�H�h��h++�woa��H��<*��~7[v�f�W�9�#�;S��&��X��c�2�>��C�}����uAD1Ĝ�XK��$�E7���js�Nvr�hF�����-��mL�������>���ĬM��#���L-wu�v,'�>q�Z_�oS9�3�ޭ7�º�'��0*4Ɲ;���-ލ|��dq.U��87�r�7W?bN⮻�7I��T�ּ|F�녌Q ��-s�B�qڎZ�����{&��1L��:�yc_v�L;�Ț�����ٷ;i �fՉ��ς��#�<������ķ4��	�Vd��k��ۈwjj�$j�w�j~�[��-î��xnD9����*���-�f�oF|�;���r�n��r[�)�T��|B�L����fTf��7|{�M\�]�Wj)�p�&3�⍻	��/��U����r��B��om���n��J���#\��:������4��rwR�!ћ��b���#�+ɚ��x(���~���="`���h
���bV�]Xʬ~~����t�p�����QN�����<��+U��W��я��H�ڼN�j�e�~eyݛظW���zrv���Wna�-]5�k�֫7�bX����4���hS�<M�`,OuB1W��߅�t����s}�ȗ�����Z=Zj��K����kw�C˅r�\��*":��l��z+);�;���_�s��o��M�I�ܦ��DTbg�»L0"�ބ�|s�Y���F��	&���D^���m�����e���ݼ
tY�j�)p�s�T�r6[`�#��q�$h�")N�r̀p��0�s�0�=�3�h��=c=V��JYi����]�7�l��"���<���e��]zL�5J�y�-|�������To�.V���õ���_]�"7l�ȩk�k����j��%��n����SW�b��mKln�9�0�xu.cr�yݝ�tM�]ꡐF
ゑ>c�8�&;���:�^�1��6��,ˎ�Xd�3*P��ն=��F#^����h
���µ�do_��N`�\+Y�Ho:y��9ȴ1I�v�n��O���g��>M`�B#���'�������_t&������I,���S��-Kv�N�6��&�2�S+�a��dd����"vj {SG���*�+�r�4X�K�rB����׫���%�VES�F@UO��i��:�!]\�"��ӷ��#v<s:�˩�[���\t��Z�Ø�1ut��pHo��l��n�n|�ة�UA*�׶�w	�-��[JEwb�_��MPh�ɷP�T�)�u�Q�*e�a������]cR�V� =��Mt�.����	W�|٢0y�E�iJ�|=3�����Z���6v�6UK�K����tz\�L;&Â���)��cq]r���k�������q{Z{�%��;V�#>��yx>��y����u��1�a���z:@J�r�7&�)�����e�e�ˬ:�5oIA��"+Tz.�:����0zy�:<[y�$��&}z����A�5�pI�g89_Vss1��ѝ���(�g$�g��l���S��i�ؔ�F���T�:�/�/F�\�%��}{@���\�Qv-�IB'�d��َ��a���j�r����u��+��W���?qr�yE>�#y�כ�s���z@S��88&��g�
�:��a5w�:����0_mٍ��˜��٦��Z��.wQ��fU^�����y�k�F���5��r*��
̫msg�n�sZ$Ӆڐ]u��;�*�L"�ڼ8_0<%��
��o�ӽ>�߼q�^5c.���$��Ǒ�;Wя��j�[�C��zݶ�t���wݦæ_��;��-9ڷ�.�=COC�gH�D�����ʍv�K��Lye�'�����3�)_��P�" HBnJ=�N�h-0�5��T����p���w�Nչ��ɭ	7�p�U�*�F���,V�2Fh�|�Ɏ��u@"�1sW�c#`��;
��׸��Kk�i�乆3�󋊙�"':9ŚN*<�ML����YSC��Z�x���3�V�D"�x��?m�{+���#�ιh�t��ۍׁ�L�3)I�"ah���]�!Fb�s�&w�mg���jvH���zq�klf�nt�xk���ܳ�2j�w;JH陯E�qS�&K���y�;�m����%X���)ص>��v�2�E+:ӻ΃=� 6��6���znxeIb��+_h%� 3�C삑�=G{z��y|��%|��es��`�!(3��菳Q�"�AwY�:r�9�z��ZUq>rR�����z�4��w�W-Ts���ԵM�0��;
�O֏7��]�ۯ�&�J��Q�����V۾��a����Њ�n]<{"��١���O3�8yg)]��=*7�t�en��%�����&26�}>܆|�P�Y0����Sp,B+��]<���Y��L��]ԁ䪱����bK�@����=��Wtl9X3�����9s���df9y�!hU��Gks��9n�K��n\��i]ז�z/�ĥ��e�w>%çg{O#�}�S�Ձ*�L�Vi87=�T�c*LՊ�]�8,ܔ_.a��"5y�+�CMkj�꾛uP�"#�����*}���sZޭ�2����w�~��
����/{���� >v�W>�7$J_#����N+w�t�P5�cTjF\t��.��ciMC�Ɠ(�˼hs9ʺ.���O���fyY�NK�4��L�#��>˭U8�H�U��-�{<���I�TS���a���ik����t�+�)�*[O[�k����Gi>��ݜu(AC�Q҇/q��`��|��������0I�Vt�t��H�Q	���N��6KN���#U+��yL]�N�v�:E��������f�r�䁥����PA�y}����Ih�ʵ�b�l�=�{1������
$ۭ��������n8�
�O��0�=�`2�i�^�K�����Im}6����%6����yn����ә�\ɚ�Q���s��qi�ܕ����n�싢P#��$��s7�;Z��z�'�e�6��`VYǋ��,Π�©�phޤn��o��rA;�{�ݫ.�b:�)d]�/���:��s(Z�,)C8`Ҏ�W��o��n��Z��v5� ثF+�n�gV��\Z[���#l��Jˁ3��>z��fC�����0�؞�r�4N��_=���L��fw&���I�u����k�{V���0U0��<�t��9���Շ�j�t���A�`6z���<l��Ѥ3DJn��@�����#�iN�	�{_g�J��� g�m+� Ѷm�[µ��Gݤ����Q��z�*�l�l�;`�F���97���AhX��=u��x-�ʋ�I�]�tn�h/R(0}�t�7|��|gB{�=�e��8r�5�=�ܺMWfr^�Mݿ/�M���1�P�ۣB<u$��F!�і��k1$��_V�����,�!]:������Ѧ�*򉲒��"q@�ò�\
�2_r��e&\99��7��s3]h�g[�����%�.ؔTAEF��<(ԧ����Ww<$���\�9��ҏ3EE�ZЈ�����D�VS��[�Y�8�J�g��ݻ��7q"r�U�՞�A]7p��S@r���4�w
=K��;��IT��w=�O2:�R���.�HW=��m��p�s2��7q=�u��B�*��5ig�	�S�:i��$G=s=G$�P�H��-�Qd�9Z&�Af�;��U�Ԏ�D���p�����$��Yx$��ȝsw%�Zq]�FN�#P�$�(�U����T�u�Ч[�������w
��p��X��t�wE�Au�+���S)!Tt��E����p�<T=�Ҥ"/���KQ:�\�p���d�s��aI�uqs��T(�%36j��{��E�"hh�X��0��f�9j�䃨^��VI�e����˟]�����v�7���] ]�d#Md��g�X���k�<$��dZ]!����%^d9��r���,�/g_[8�uY�������/�?S�R�S���|C��<�u�����<>ݹ90��|�m��o(r��\o
��ѽ�o����>�z��ׅ��&"��Ȅ�|�g�?|&#8������_���={���y};rr��_;I�!?�;�߾xw�[��O���]�<��)���~q�W���9�����F'w����~M�97���þ�������ُ�fg�L|&���w1Bbk=�y;��_�I���*���a���|
c���߯�������o��7�'N׺}}��ސ�w��y|���w�<�-���8\>��&����'���uH�V���|a����<��Ck�L������??�!�܇�S��>v���s�>���0��_�}�SxBpy>�w���!�ϗn}}��~O.'|?�z|�������������~���.`OO�T�C�?E��pߐ�Ѥ�j����;봛����>[{w+��{��������cߎ�w���q�{����OI��\}���.<������<l�����?��o#�?���o	���w����b>鈩�#��3֧]�\�4��G{��9Rv���G��������������o���'�0}C��ۓ����<&���v��8�F'~v��>����&}����S}g.���~���g艘���g�5�:��9�{�l駵��{w��1?���8�'!��nw������<&w�?�?����?�y��e��ݹGwԝ���!���oI��:v�����|�ߐ����}�#�1?\�Y���924�=��T�|����@��y�������M�=�{���+�w�V����^�z��}C��{C߮��aw�?�Ϟ�����®�y��)��&�w�c~C���y ����a�öN�SM��ϳh������5�T}�l���b�z�}s,}�����)�����<{��o��P>$'��N��nӏ>�hx����Wo>c�}w<�����`�奔�w��ý���?)�V�zcg��Ɉ��"OoY������=��Ϟ=��We=��9�{���4bwֿq�������}���[w���?w�©����x����}Ƿz��w�i���9<�xy������;rr�y�v��0�;1�7���>�F�*T�i[�5f�&�0�Wȗ+�g�%��h�� I�X�4���-c�g`�S�J�:f���u�����ǯb�ެ�:�7��*��?
yk�Ǟ%0����/	3��j�-C�2��#�T6�}-ABy�4��=uN{������}��_Qx}[6~���|/�1���o�߿������~v�����:O�9>��N}v���r}O�޸����z�e�����|��e�����n�����w�|W������^�~7���I���e7V�!�?�q����7�o~|�۟��x�����Ͼ6��y���S|M�ޏ���S��1i�)�����|Uׅ�[�ܼ~���������]��P��(I��!�5�7!���?����8�x����ߟ	�!'������s�G�}�)����ן߼��� xK���x��>���m�zݚ~=�'oY��g�%㾏����{U?3'o�t��v���0o0�N޷�?����0�����s�M�@QC�|w��?\�~�Sx}�rr�q�|�m�c?�{����מ~��LF�}b�����{o�=���{�;�w��yWyv�~'�����{q���<����v����c�HO��~��<��N��w[s�< #�;I������t}��{v�7�w��詏L}�ǟ��D��x_����}?dǧ��������~�����\}C���~���	2�O���߼��]��t~~�xM�	�}q�cnO�#�xv�F��2xv��ם����i7療z����]�~{vߪ
C������@������k��}����P��C׾��990��>���ߝ�p}�rohI��'�p=F��'?��>�����>����7��o_c;{Nw�_�w�l:ˋ�7b�׈�1�w{�11�J1�o��������<�;ô��ݏ�_-��������o���o[���ψ��ɿwΜxw����>~�����>P�=�q� (��?>����pU��������N��⒮��+*����������vN�y�@s�u�~�濐�]�5��oHra�y�����]��w�=��}O)������{�I�!>ݽ��ǔ��}��{��R7�W/����hv�܉gزҚ���?o��q?�L}��"�aC�i0��?z�˼;]�nw���\/��������Ǵ=�Ʌ<�x��o/��9��6;�e���}�>q��N��z�����~Bw����pG����h�
�r�y���m�۴�26l�;�{�F�ٽX1�eK\T�C��ɾ\ap�Q'�Qz��s
��ZT���;����4�v�۝W�\��!���̚��z�n����Z[�z���{��Q�E\}�2��pt�Ow1�hkj�����ޏ���k�;g��r�����>}�Rv�����~���N�>�!8]���q�='�J�����rr�<��Q����I=��<&}~o{;ӿ;�����o
��t�}�#|�kz�G2g��0OQ�}��������� ~I���ǌr~}���M�>��	�[|N���	���?='�;I����۝;ˏ[�xM������&��O!��������U�o�)A�-~A��=�E����!����¹��;�xw�S�s�O����]�P�����=?�m���o.��M��nN�Ϟ1;��{�_p}C�aT��w����z��zv�w����<';����99��8x�����O���>(O�
rr����|��۷��q��G�o���xC�o��&��=��w�iP<���}�;���~��yw���㿻�o�Ʌ���z>��!�
��$==�]���2��(Y�ײ~鏄���r���L�S�~���N�����ݹ7�'����������������7���yv�>�}��\.N�����ˏ�%w���7�ߓ��LB���NV��Yq�܎{����k=�p1;���������S�>��w�xw�9ǯV9\HI�����7��Lp��*��a�>�+������աɅ~�y>������a�|�vߓ˺~�O��>�%���S����'��{���ۧzw������oi���\
o��y�x����+�/8�|Nv��-��㓜s��w^
�(�~O�s��V<�~�]��������������?|��T��ߖ���Yw=_1UɅR���x�����:��ܮ�q���P$�뷷�_߸���7!>��	�\
o��>]�;�����ڭ�?�y� 9�]�<_]��V>G�	����^�װ^9k����L��DE;ӷ��ߟ^LN��r~��o��0��z����r|C���w�<+�&��=���x1�L��ϯ߼m��w�c�<��&�O�������aC���SHD���(��o�it�߷��3ߎC���nO/�Å��7����s��%}�M�>'!�?���o?#�!�v��?'&�]�!�����'�w�¸�Bq�������ѿ���PT��!ULQܾꟶu����@&2����Z�9�� I�aի�qT��*۶�V|%�s��u�g䨸nC]�c�{�Ѽ;On%!Y�N�9۸����^(�-ut�
9�&՛Հ�f;[C�f6�PO���J���KS,ٹ��잓�hX��'W�	s���L�s�祐�
C�}���|��U1_P�ǜQ�<&�$�w�����.��ͷ��;~t�����o	�!~��߾xܮ7�y>}���o�_c_�ɾ�\s�'8���]�����{��=�����w�_�ٕ{sOs��ο�X�� >�
�U1_�W�Â��|����&��kxO	�߾��G��������;�n����z�m�c�+�;����ԓ�������ޘ�;���&.f~���G�Gz���J���죧�}b��꘮}����N�m���o2�]��N��×s��x�,ro�;���N���w�q�7�yL.�x���S�����v<+�1�?E�q�D�&>�W���d.�v��©�9�}�S��b!�	�����4}���ދ����N��@���ߐ�v�{����<�Ӵ��A�����-�7����W+�M�=�'���=7�k�6Ro��������>�˘���[�e�~��̽?����#��O�~��w����
����ݿ��~��|���zOO�n@�����ˉğ�)������&�o'�='��P�y�}���'�&�t�}Hv��<u���o�_ �%�g���]{�+�zQ�����3�Dɼ���8��o�/�ǣ�>7��q�������ÿ8�����߯P��U���<
���p_����&<���7?S���c�zL.������7�9�J�]��옊��c4:��W�<s����}�]��єI'�<V�|;��M�޼y�/��p)�^8?!��nN�������]��Ͽ��>��aw�k�����>\�󴯠?y�<&��;�}�cǘ��f��:��YW��˒�+�M�.`�o�����oi���xC��_m�]&����~�!�(_��ې>����kzh�?���Ԧ�f�`��o��N��§V/g�F	�Ev��=\�:չ7�g�#�0΋���ʨx�t+��\�)�о�s)i2~����|�����ɮĭ�=1wr���
�^oG���i	�q!�c��܍l&_(�zV�K�������Y��:�\��N�ܡ't3�6Qi]��R��������L�j솭Fy�Lf�5ˏu��w���+<S�Ly�s�N;���%1�>�/�f�F�S��G���{��}p��C���;0W۷�\�r��g�f�L�x�$���.��=FBk��0�����y��v��o՗�bl�!H��]�5�S��J�]5�G�рk��w�y��l\��X�ߋ�a���8�B��-r�s�N�ɵ�Y�%�\�T�� ��¶8Rc�]w�;u��;9sćS��ӟ�t3�dژ�$�����F˯Q8r"|�vؖ�����j��e�Y�q������)k�NVmN:�J���ń���8dM!�;|΂�iR�=fV�Z=�_nt�n䭩���K�x=��h�}�g���2%�Jڭ���,���O�	�'iu�r�̼�-Tƺ�Q�����5(����.#O��n�дݙb%�w{y�]�-B�C����/]9�mݍ���c&�3#y���ީ��<6���dg�>ϛUR�sÈM��{s&Ȍ Q�@�RG�* �)�<Y9U?tܥtt}������W��'��o��΁�}w8�{V��Rf=���<�L������#�U����`Uc�U�6'�9�53y���~����t���SԺ�����D�[��>e<=�qŲ��|kN	i;(�'�u��96Ů������S~Ust��Z��̬��c��Gk3�a�3MG�X;ך�-Fe"�=�3�f���m�2�~��l=�j�uv%��S����w�f<�=]�yA��_.ysz�|���Ʒ5���}�ٮ���a���nU���/μ<�F�����F
x��S�*n�"�VQ��Lf����� �'0�l���]�y��A�қ4�5���ï��r	�ٙ_k[S��2}��"Vf2WNp��w"�h����\u����}�l������D8:�F a�PL>y)���wc�3�.���b�F +p�N%9Ǫzw���;�r��u1���eӐ�e����׏>��E�saWcL./n�YWnEC����s ���1-o�$K�tT�gzx}3���w�e�h<׽<����{��ť�=��� Z��g$�͉6�+��[zf�"�9����[֊Ǌ�����:i�o!g!��l�|��C�f�R�����"Ku��U����75:�����"Kg�#5�5C�l����>�Q3��M ��&T����%}!U������u��IH�Z����1�k"�❤4:نƇ��1�ٛ�TV�N���qw�??m�$�O^�U�c�*Ps�o��z��_h]+��H�K��%[N��ɶ��X��4�>��eAta�lP��Ud�h���%Y[�Q�+�b�Z\%e�W�_y��]�˧��}�} �;�;:J���U%����
���m�$o��#J�U�Δ����ɋ��4:{��lgu�G��s,Z8�{3J�Ve�R��׫���<�mYgz֫C�������4�ruRӣ7B,��X?{�T��;�q#�L���
r;�ۦ���"��3��Ý#G�7%���c��b��_,ϔ���h�7
1ф�|[�]�,@1)���0}|���j�e�>�N�F��0�6�d��i��2K���kNQ5��Tf>w,Y؇q�8[C<�>��۠`����;���o�Ȼ���4���Xr:L��i��݇�3�u�T���Ӷ)��u|�y�Z���lN�˞	�{�y�p����n��@!��QY�2a]�s�v&���ꮼE+�V_�/��l��F�N&	���x�À.Cܺ�/�V^eRa��ym�4Dn�'���\L�۫kW���^���h��W�`�<'���X�=�V8:���?�W�
g�Τ��6��*�h\Fmѕ�a�%�>���T~�Ek�27�ʛ?vs�rü}c� H;�����m�)�Y��#M�u��"3_�|Os��sϖ���<�^�C|�S�~�7�J��zx�����OmY�
W�\.����}|���ˇP9{c[p����>�y|)�ڲ�pT�=Q�]L�p\2��:&�1O'�+�u�y��?bX���ԫ����w���X6|":]a�lx^c��k�5�n�gS��y	�t�,�	RY�b�?�qXnނı��;��k#'����d�� ��8-4r�="�-kR7
`�����7�MdT�	*�'��S1�݉·V�\B��1V������V��h�I#�3b�R�5����&���\j6d�'���3�C`:���@�{��0�������~�n!&�z�_k�H�16s��B����࣎T�m`c.�r������p��p����5g��ɹw�8�U�����B�)Ɣ��eK�gD�&��l��^ᬝ����Z�����Tz\�L;c�]8�l~���1�Ss�L��y{�ow�Y�I�Gor��ۆSUvӬL�����{��ɸ���!�v$}�o�a�`VS�����ӕ���������hrU7�p� ��F��eڥV���x����,�Eu׬��?_t�����<�NͿ�����Λ�@�~&�����Rn�_y+�7ݳ,���= �q�W��hZ���N�R<�P���8i�j�5QLD�����N�.A�oZP|r����u�B��J1��m.�m����������4`SR�Z�$��Z6���;E`�9P[0�P7r����������\d��ÖAZ�v��� ��4>�Bks���<7>��O�U�ΰ�ų'���;�Ø�u�p�8�b��O*�����9\~���+ir�`𫴴ep_
���<9E��U��龛ⅼ�.q-y�7��[{���=ށ��ߞ�`w���W�/��x�8�.����k=��	J�+s�ΓEK��rn1�n�C�s�s�����u;���.�b�+��Gr���wK�mI�Eq�9�TT�/S̄e�о�9[��!��j�S�>rA��\%��:�߷����5�w�{Hýu�5�(xm�.j�,d%����O^3�� AX��=�M���	�7dP}e��L�����]��}F 6��\�!�]Os�A;R�������Ӗ����.�����,�!������w�;o:3�i��*os�5q!���.��<;+e2��25���>�c�1(�2���Eٱ��2�P��n�V����v�5ٛr_��q��n��.rPV�uӥ!\+�T����	v?2�]D����nk:i��B{j7z�⽗N�%Y���ൿ���l��V���Rag2�u8G�x�����֤(�]�b��7��6y�n-g��rO.�g1'���P_l讄��G���uC�`�[#|�wǲ���(��&��E�C��":Ո_Wm��"�=}	���-9K�R#o���n>��bW����!�K�20N0�7ȧ��'��#�zCK���k��n�s��#K��n�o"��3�&�>ϛUR�s�M��{s&��� �g�P�ceĠ�rP�hY��������v1񧾇׬W�]�juwx������kvPz)�mM���ԩkA��w(��B����{`[�/":�v\�l�fđL��Ǟ�:���=Y���=��fV'2��P7f�&��e��W�����Uޚ� �+��꣑��E�V�e�hT��_)�ГW�(��,��ε��d����v��S�J.��[�p��q�&]�tU�<���+}�EM���Ѧ��r*���kHY�sgQʶ�>����8�ǙaX�h�s+ a�pU&���N|��wd;�5Ք6\�
&p�k2�s����&�D�����U�9�N������?2�щ�akǟssD��p�.�[{3,kGQ�Ƒ�9nc����z�ݱ�v���5rx��p�N���;8+�_!ľ6u[^!�^;a-�KY�*��f���,,�Ys	�E�'LoE�#CQ�CGQή�{o\�;Ok}u_y�g��s��O&q�f�+Grz&-���l�Qb}'��z��fϟE�;Yo��I��Y�-��[2�/�����&�3�s^Y��#wHﯗ��F�&@��OqIY�V����m��Tƒ�T�(�pp�{��j�HR���zץS�]{u����lT˰81
��)f��H��4-P�� �N�!z�3��6�U�3��A�u�Y&Β�RZwyy��3�	���Ɋ�.E�{#��ٴ��W�\[ܖ��!Y�O@�Gt��4U�����w�Fs�?m�:�Fe�V�bASξ��]9���E�P�ͥm,wV"~��k�f��c�T�+* �u��Eks,�I�Nvq4�R�6�jH��eG	��݈\!�M�wt
:�m�p�f�{Ç��6��ʉ�D\�i��>�]������V��VQ��\��l,o2����(l�� ����j�AW$c��L���B3�f����z�MVV�hv>�������Y{+�.�n�~�c�ใ��C��q�b��|��a�(>VJi^�A�2frκ����X�E}V;M-��
l��ʌ�<A��x^9��CU���݃�9я;���Yg��V����"���w�;��7�|9�T�#�5�-�Q��˲�<��';έ8����Ɣ]9�U+Uo�� 5���H市�\���S��^V���]9�t͐_P|�j�k���wi������Uj�ݏ���;�K<0J��g�A.��Ƶ��;gb���󩋐HG�Ū�͂њr����xxWX<\�F��:ߝ�`ޥ��X#�	�ON��*�{*���[�fn��|���kѣ1��q���콤�MTz\�����L�7^k�K�G.�ޝ�6�ڝ
]��͐f�A����Ҟ��.�ٯ�i�����L�^CF՝[����\�?^�n�+����ņrq�ҟn;%�g�V�Z�$�W���-=��ܱ�CDn��ok���פ��`v���۝kn_w<��R��M�L�IYw)s�+�����D�ʶ�gy�}(�]#���μ�XO`Y�Sld�ۊ�@���4�����!�uU���F9 ���������T<����82k��6����Ԉ`nN�a��v���z�sH{sӵ�� �]��j''N�.��nQ��n��2k"�n;�֩芢2��{���4�ǀB;�� �m�'A����{�^D-�`M��D�.ݷbGMr��[\z��*/.S�iV�h�`l�gd��"�]����N�X|Z�y׫&քE�b��;��p%%�<0�[v��xVWL��� �ʻ�񶕈o�N��ê���N��0�:AoT�m�&襁�<�53>92��8��m(�S5>@��$�T�i���C�=�M,�\��N��H:P�G�k�y�.y�tw'v�NS���uCI+9j�98+�t��k�DҜv�-�rs�貜�WJ��\�w�(ԒL�Q!	0�U(S���I�FJ��S=JQ�Ҝ��<�/\¨���KS,T��*Eff*��䞮��
*���-#�3�:F�[��$��!�)=wP-�j)�i�8��N�*O7U5�N�)ȫS�%���qL��8t����^ `n�G���ws�ʓ�O]U�4�R2<�B�	���\�\�:"
�G���p�B�0������N�!�VI��RQ�r]sܳ�bQd�d*�N�n�z��jVl֨�ZQ�{�xa��R��$�n�D�K�mb$Z#�K�0���30��Y&eKS�&Eae���V�<D�D���D�B,*�$�;���VX�ht�fk��j;�bJ�"FQȶ��&ȋVV��Zf�tP������[�?����q�����{�}r�(^���l�A��w��Fx��{��sz2�T(i��bac�7i%p�;ӟ�>����y;wV���
�����DT��, O�p�w|���w�/G�^�9=�uq�'�=�>����t�Y�^�e��](Dx����EpQ�xM�<o��nnjG��^;�h��ݫV�o՝�"�wHYl����X���v��V�2��?0�n�;�Ǽ�o/>�6T�W����j"��)�CC��lW���;T���{�^cG�"z�4C:��ͩ�x
� �[Ss�v��� F�G�N��9σ�`5Y3�[:��(��d,ʪ��%��7�t���`RxFG\29;�x��Ћ-<�uU�����l��K�{��q��{x�W�D����b����4����x�����P�]�����[����"�U�w�طlX�1/W��z`������-WCx��Ǳ��:��ŷ�}u��0��ws"BP�k���~*�<ǋ��Π6G�z�a;E�/�Yw�|�̘�K�[r�ιN����C�ucg!u&2;�㘙z�Bw�C>���>���T	��x4-���M����V�rd[3��:��r�>�i%��4���Ѥ*��Kn������Jgaԍ�����S�^^�n�"��[�Mj�	t�\�ct�ε��2�"_^�?kK�W��fu&�'�4P�w�8B��w��HβS1f.�E}_}�|�����k�,z�'"*�3��,4�Y�3��0�؛�C���|rg+:�m�֟�F=^k�W1N� ���Ϧ��Ӣ��U�9J8T9�*�F��l�ꮕ:iվ���b]�M�ꂷ�@�CExWh<�a�G���=a󃮘��w�;�Ҟ ��zDzn�w^�~yfY�XD\#�Hg�"f:�|��iNGeٷ[9���;PԚ@-RɄɬ��3��<�B�Z�ev|�|�dE]t�� _A���
�A�r��w�ݷ�����%��Gz	̊C,{��+z6 ��#�]̮�؞�w�A��f�:`L����}�]]ʥ�ڌ�S�W^O��Ȭ�L%rt&&cm+�ZYYFÛ�1���݃�}�P"��G�:6&�����&��#��F̐��!�c�/����U�&g���N3/p��:u�Ql_z�8O��|�/ly���j� �s�S����mʘc��,NҞ
��o��l�p��� <�w��+@=\N0�o�[f�#�ȹi���z}�3^�m���*n����Q�uw���	�ޜ�W�3��XI��5_y3�*����l�h����i��QK����Mx$�]
g������j�Fx�Q�V�}|,��/�܎E�f�(O�3�S]I���X��Հ��{��#��5�>�����h��iF��Ϊ����u�z�;_�;�W�����͆�É���L�:j�Ԣoɰ]�g�g{��_.<`��u�L8�����/�X�Siә��({g�<�C��3�kI�rٔ>���>ve�ٱ��9\�*�koh�u7�ސO�9��U���rAU��,>�w�e�"]=��{B�_��~?ZϞ�0�Z0� ��c �,�T>
S��7q]f��������e�����#�e��ʅ�*�w�����^��_��λwb�����U��#���ٲL�Lfz�ޚw�x%q�$\
��{Wþ�e�Dh�2>�rq��k����M�Mn��.;ϧ�c��ۣ�������!�}Ҋ� 0WL^��
u�Eu�|�S�]�3����4&��^��9�%�#��^ʄ�m�h�4U�	�l�9N�uٱ�a��5��a��Գ!o�C�ç�+1�$!Q�:�/���O�/��͐�"�@��k�;��0�T/辰sW�c#K�c�g�e�f��wT�����&��/x�G0
(����'�p�ݎ��ݍh�}�#�2�,y��o�*<���E�l�(]K�FV�)C�V���.��v��9�5]O��1t��)�sbSqUX�z�2/ �7�LR3�+�l1��P�qø+0�����{��DI��*���:��^��""#裼�p����7����A���g
Zźzv�/��K����;8W<Hp�"��&!wv2����<5����P�P��Hv&�B�C�K}�2���N���F��.�J��7o79o(�뿜�Tg��$n�h���Ƈt�చT��Y�kG�e��{�U�4�2u�gP�>��w�{�J�ݠ>sr��fU����H�!�//�\I�Zt�d%,>;w����q�,���4.;>���ݙeۙ����r*j�~����^������wt��ӛY6��c�dA4�gͪ����Bn�K�{�3����Pu�>�=�/o8�d�U5^>N���h��ٖx}�u��oc���f�-I�!����\7QV�WQ{h�s��g���c��e�YVf���eV9�U�6%l� FwR��W;.KX���;�udH�������9�jao���;j椼���q�w,/rr�m��d�k۔�y�L̮�f��κq3��㋦eƞ�s�1Lr3oFp�ڡ�ʺ^^��O3�B�D�E���%�\q4u�277D��u�$�j.%Z�*-6�wwiT��LE�V��{�'��sSw+�,z�c�E"�v|���HG;�o�7���f�>���ǒ�]��8�O�Pq���r�Xȹ�w���"�k3�m�J
��D���e�i�W�}_}��T_y!}޴���$�%��^T���ں������`LV�6x�+�-[�(��"x�JV�p]��*!!�u;�S,0;�0�=Ϝ��Fc���sq��O�vu��7����<�e���~�I�A8��5:��܌�9��N�	krZ�s#����%Wݨ�+�\�p���"�O��������2�(������Y�T�ge��NB,���V��=��q��p��fE��}70f�!�u�\w�&���]�����kr��S���4a�k�v�j]u�Ȇ���<��s�j��o(ѽ�滽��ۗ�̱|Sł��������g!J��}��V��W&w��Dk�Ux��1��q��/�O=Im��3�~c�!�E	�"�Q�N���f�쌆�fnd��/`eY��M�Ƹ+ť2�!W��/�c�d-���[ž7����bÕ�0��H����8�߳�lU��uƆM{�P�a��jrT�x-�N�^}��s�6�;��t�{3�o���z��g[�J���a�̹��񈠵���uX�~`:����]��OsR��֍�Ý��$�yM {�oz�7�+�;��$��J��7��v��w�*��y�MMW�r�rlo͢�To/~^��:z�ң���}�ڝ�)[���{lX���O8�^��O�Z�>��[�4��g�ާ��~�����(S��/7�q�=����w��L*���p�Y]�c��Hy:[N
�/}5�\+�qٍ,�sӟN�Ӓ���\�X��:��u�H*�F�?��6��������N�0����uo9�u1����wa�12��N�hdCYq[��:o��8�Z�� v�w����R��$��Ue�t4�f����zm��8��7�Y��O9r�ű�>­
�3w�P���w��t�^7�pY|Ǻ�:���bʤÐ�T�=��t�a�y���S�xk3��P0a�½���
����b�8��a��u�{<��J���d�ڭ��^t+3��/�Y�o�*i�ؗ���w�+_	U��~M�j�t�t�=��$�T�p`ݻ�.o:v>�
w#]̮Ȅ���P�=�	��k�lW�g�]l��)e�j��]��sG2)���ҕ<�b5ƻ�\5�#�T���Q1��D�P�/���V^G[
:��.����k/��r#1u.�)e�`S��ο����^�{���K8{�(w�޾/�!�Z��NW7�u�B(8tqc2s:�`S�m
�|��N�(yos��i����6&�L��wjJ�VI}���U}}�)L�k�����E5�:b�B���6-5�Y�	�UO�:�����N�h-�j�jqv2�>��E��'�0�l-����7�v�ѯ�nA���6"f�$9U����F_d�ZZ�q��T6;t�C�h�@�N�cP>�5s�Þ�B���2>��8sv�Z��'�흖	X�#!��!R����n�2��^D([�`�d%�U�z֜jQ��Fy�#�*r%����l�-s��G�����и���:��S_HX�p���N ����=������]>�'��匉�&T�'Ng�շ�q/�Pi�@-����΄�\��$�w�A���x�a#`�4	�]��"
y�l"�eڭ�{��vf��#��XӋ���%+v�l~%s�/t3
Nz�[�eټşb���Ju\���I��f�lOu�1R~���\j��Պ��j�ȫ���M���jg���58�v&�7���B�����ݧu��a���܊��)����>�@]�\%P�i��[�n���
U���]dͳ�ٜ2�:t������ҼҬ�S`�8q��˫ wK4��<���^dnj�k�3Z!e�ۧ;i0�w��Vt��E�|k.7ǻ�7����,[BC����[K�_.�EG��nC��p[ף*�/���¬f� qLv{�/�.�m�s��_W�}[�v���I\v2g�ۍ
�i�ҝ�c��ۣ�et����C���_@��\k`;��q�}��$�ps�d�!�O������I�/)�g}^oG�](�U�"�No|�d򎙼 �=M��g$�p+��7Ph<��T�/R̅�;|7��V�lBv��lV_I�����6������`r W]3RM�Ö��.�Cb����AbX|���쪪� ��}���4�/R��<K���h�(j�+
�?dB�c~x������ɝu�Ɓ}-�i=v�����<����x�s��C�S�1�|���:Cm�ť����,v�wnM��U��F�!;��v]���^u)�����LJdL�q\W�]��LU�Է�����͒٤�(3�f�y���pSX�bv���s�Ŀr�t�HW
���q(�]ރ:qsQ�[�M���.����)�oRϜ���u���y]�=�������Ʋ�WMl����J1��>H�������ٹ�hm��i�AO��m\T��h�Y���}7V_�E���Z���4˨��T(�y�K]���j�A��4r��`�)>��������6�T:a�fj�`�4u%:����\��g��_I���9��0uF�:��'iِ��qGϭ*�`��x-�X�p�%��S�'��������諸z�Jz�J���4��i��������sg��h��F�˂�y�F�ˍ��.�޾��~������a�*���"��X��U�65��kk1){5NM�V���]��Q�������z5�kݑ��C��ΨTM�r�/rg*�!U��P�GA�4S��0�@�9= ��fn;]Ü�
c�����\�����ГW�
��Ф+�3�O��Mti6R���۸3�
��[B\���Y{S������|Z�0lt�gVЇ�{YV�f�vOu 6y�n��Y�0�D42:�̬��I�{����w<[�K�f�駊��}_ъ���1i�΂X:do�T��Ы�/�k�"\� ��v�NS�lm��|�����y�}U?3B��n�@�}�ñ�g�|+��oc�۶�Ί�C�4\�a��Z�NwUj���j�jwC�C�5��
x�7�����k�g39'�lI�J�A1f��=zuU2��(J��+]��!���U���5�"=ϝt�����:�����G޺(_�3~�d��,L�6{{19�PCM�`�<{��<)אA�"�s�����WOCϖ<�χwd[L�B�r�qa�T��TK��ni���ќ��қy�pn��Q��l����A]˄�J�ɋ�&Ѹ�܌��DG�ν����q�@z$J!k����S9�E7�fU�#O�ْF�����ښ�T�֤P�3����si��0��?����
d.1��E��!,d�a��3�fNKw�mTV��q1[�ȫ�2�Bh_����1�!n�m��,�`5�nc��	��$N����Y����Ժs&�=��\�$��40���o�v.����Tc�Sٗ�^k���[���Aa�^�΅��*��� U�Т_�x�t-}�CO�}��]V>~��͵���&�=ۇ������$��}��|$���}/�@�����U��?Q�Onڙ��-����*�XE�e9�t�sӟN�Ӓ����R��w#����Чg���h�;��7o+�w���d^��U's��kA���efM��*����CYq[�/���qn��@v�q��m��)��:H�g�*f�Fp ��#6�LB�L06&�P����x�A����M�9[�v�!�0pF͗CF�R�a/��~���{��݅W�����^�w��ńW?���*��|a̘�i�wZ�.S^�z��w�z$i�=�%^�:�ݓ�vT�l��]3!�=3pŗ�5rͫY��B/=�����^Nź%��2�.ͺN9`�7z��k�J�EC�-�]V	�����S݀�P��=�Z����d]�]�R�Dw��R�u�h?�e�2��x�-�4��t&n'v��u�ldIR���X���Cf���r�бW5F��ʇ�{7������D&��:�묺|�,<�Э�uą���3+#ⴹ�*��y�\e�y��g1؏���o��!��=\�����nT	ִ�:��[&���y�[�z��`7e�eo-�N�q�*WV9݋���dj̾��*ڐ�
�f���j��y�g+T���N+�C�\:��*Q���巖O1w�Eb�Hmyt�$7R�:@7��u��)ޤ�J��gqȠ�ZRܱ�Yڜ�ol�zjv���C(�!���ݾvw˨�m.�%�vܫ��A�|)
��Y��E�����X%e�U�wt{�S �4�Yh�5�9%06��qou-;ԵVJ�}o���N�+n>�Qv���8��qLiG�|��6�fJ��@b-֛;���$�KT����B�������l�v7״��ڑ��H���)�4{y��ܶ�r	m~,`M�w��3�T3��s_3�9����Z���t=�s篓�t�؇��62� ����������6�����～��H���|��*NTA�*ЎV��5�
��)�
����˒}�{�Վ?!��`R��3Uʚ��S�'��T5d{������s�{��cT�	����U2L�6�F����J��K����Ldzz�!��5�b�S}F���D��9���~uծD�+�X�i���grl����AS��XelB�i˭M��YA�y �Y�p���FQ�i���$:+�|�rs2�Vs��
��]��P(�Ϡ��P8t�5�p�-j��OzD`�\���$z$�b�녇�Tj/,����9��z�j����fh'G�l8nwYrn]�p�w�<͋��_:a��;���A-s�����HRg-u�`��y�<ߧo>����8XG�,k'tJ�8��i����ť�S�ip�J53s�,�[�X���]]�é��殹���t��Q.����{<"�y>5�];�|5�mH��jm���n0-��g��P�U:�}׸�82�<x{MQG�JW�7��ƐYǗdguD�*C��
m���ZQ��˽��M7��_�1q'���O��Bu�c҇Q޻�(��oSZ�|�y] �@	u{u�&�/���b9\}�y�-��Q<�Wv�TH�d��\t�T�S�M����1������]ݚT7�=tj�l��ت�3l���F\��� f���\�">���P���;c�״�5>�Õ�PB�}�J�HȢ�(gy�U�=�<*�3Ԏ�玈�Ri�:�'<�Q!�',4�L�M�i�R,)U@�8]���h#��G�Y�������V�:Y A&�'ni�m1P3EV�j�.EJR����y�e�Q����+"�k�d�ZVKU�"􋕫ww˕�ܽ5RI*䊂��q�<��*�{�TQ;ur�7t=/6W�CqWJ����C�QU���u#EiHg���G(M�E0�ͫ4W	�wh�$u]ES8�����f{��Ĭ�-	��D��s�/O$���*�QSB��TB��*QMAT��縔bn{r��-+L"��DVUXr���Ft������bYbRU!EP�4V�R��)-Q%J����X���tֳ�#��#wv:*�Y	35����HA��P�3R�D���ef�i�R)Yf���̍�]�j%AT�&���
*���HBdht��"N���:HX���%Q����U� χĒ����E���o�q<����t��6�ӷV��}7o�}��/:&�dtgVM(�maT��<�LS�%.�+Q����G��/R�����Yc����2���T��D�G�۱�xg(R�n������	�D]"O2�#%7�8�GL�c�jc!:lyfY�dkfܨZL��ּ{xB�׺6�حJ��k��&m��__T]���y�`����:���ޟ{M`���#�֞ s�:�w���V��c����W�����z�dSa���%oF�R�v��Zk6'�]��l.k�^�D�bg��Оg�+�Z {SG@�^0�q����6�ݑY�	T9<6���rK`u�:���J;coZ���F��i�:��%OHL)��!E��ٓ�Rx؉X�ɱ��sg��g]��t8�f�2�ߊ�=�|Z���A�L^�u�j��z�f�ע�q�>]�k%����~zc�d�t6[��6����B���o���h�DJ�W�IQ��m�ƥ.�h���̬沥�D�u������������q����혻-�㴁p_��W���qfUC��oeA���0c��s�6�,F�2��t�x=�m����~��\�F*��h%��m1�V�W�4[��R��l���Ƃ���2=\�3ۊq[�I.�]t.ut���y)t웎.�'���F��肤:��+�͕�Tʹ�9Ɔ|C�{>��u���b\�WS]��"��ؓ�{�wЏ}}}�����~s�����#,̕�v����=t�aaO0�]L�5c�7�6��M-Uv��Q5ڦ���]%R�s�;�ϔ�K���n���I��س�=
g� �X�rV�R���=T�n�$����^�B%�#�h5@������J�f0����w��p-3ם��x�̫�|�O5|s�����zi�~��ʮ4ۢ���^��~�ic�'��;�=�}kщ��bW}/�fq;,T���Ӑ���,���,��-�2'�
��pJ�Ӽ���X�;M�g�5����Z�s-l�'����7G�{n`�2�謿��]N��m��ݍ�v��)oh�6����]C���T�/�K2�OB�󕹯!��_���~r�Xy�s�:��8�Uzy� fr%��n�Ò��1���䱐X� $��T��ސ��m�_-Ϻo.���#M�9.a������g
�b�>]U�;u�t�w9/kg�TGNGwrֳ�F�V�/W<HtS��s�wΡL+���la�2��l=igj� ��IG1}�>�}cc�b��O�����p��m�T��sH�^_{�����n�0����s�eG���[8v(��E�2��c3�3�b���N/
�֙�����Qt�o�N� a�)���^�Px띯)�7����_o��ﾈ��<��NR̘ܽ�ou�3��ϲ^u)��3[�2&����L��7��b���<��X)�$�A���<�V��;(��L�HR�%qV��őV!L= -��7=���4Wv��0�MW60�$�9Q��ϒ�t-7fCؗnfzs�2g���^��Z�'�*�YU��(]K����KqO.Kc �Dd�>�m\T�-���܀�{�pR��|�fg�f�=Yrơ%V���ꍮ�v5�~�}���*���wɔ�U��ԝ���5Zf
�r���^����l���U�Xh*Wl���qUF�|qY�O��򲧩��$�f��ڹ�S��;��0���u����{u���#�dn�X磈FJ�
wjI��y�DL��j�37���!L>��<(��m��k>��f$�p,�G����{���M�Q�>v�����%��ae�N��lu���-Y�ώWOk�޺�V[��8gR�B*p8ꎋ�ۻ��r���ed �ʤ�<�>rv")�s��CB����rK|#�C6�.��V�;�,��,�Eu=k]n�
yC��#���
n֛j��r�����]vP���P�t���+��o�;�cY����v:( ��@8��0���b�=:��)�c�C	cN���a��;�����W����R���݊%��t��챸�� �=X:do�V�HV}}��`��'у�ݠ�+Բ�µn�x?��Al<y�a��}�/�ȃ���(xW	�7����v�0�����B��:���&Jнb���p�N�2�Zk!��}q70f�`@�3R	uS1ޢ!�q���y8z	�v�#s���l�4��l93�@�h�,͛���n����*x���]�S2ƻ���kP���jg)E�J�(�~ә]�I�~T��|��"�eh7f8��.��aS�&vb����j�Fp�C�1�Z&���v��2a�/+$t��é��-�6��>йh[2�j]� �)�����y���!n�x$�GqF݅w����^��s)[�=�2��<uM'�U�`.O�A�UQJ���of�C�����2	��3���SY8�N�.�j����5B*ņ�Dw�0.�zi�u�_c�����l���X�ӧn�Q��e)\���C����}�wzF'�:�/�>WѠ]Z�}Vk�
M��c�sE���s`je`��VY�b�Z��a�~�RX��9���Bz��!�)ҟ��_%L���^��6��[�\��v	i��ս�oa�`�D��X��yx=�Y�nx%e�ک�����ĕ}w���k�Z����ܐ��9��UQ�}ܗ���Z���@�{�^Q�g`�cZ��y/
�ݞc����P/ƐY�Р�Z^yY�{ڧ���Mб8�����h�7i1��q���ʫS��]Ebۭ@����;�
�/
?���>�P���?�>ڊ�������iDaf�Ʌv�`tSt��<��F�a[ڗ����]�4ǿ?L,o�u�)^�=�i.�	}��8,�cܯ�Kû+��~������Wu��S&�*�.b��t��|^�̜�MX`ٺ½�����<%��s>������^[�19cc��/�P�Ld|�6��,�"-�C#]���xmls>	T>���F&���4����滤קޘ.�ԫ�������
<g(<�h�Q��c7�k��x^c�:[�5�g�ˍ�����/���)�e�!>^�-�y�|P7�	���9��f�}nE�nL�:�P�1��>]y<FŦ�+0H�!��G`��#�j�em�[��1�#
�;����UR&(���;���&#��h���+U�H����R=�/::7���eB&�[��~��G�$(���.�&P��^W�⟯��F�3i��M`P�z`ZA�n�VfpK�1��3�xp�s�kK���jP(�I���]/9t�Ho:욱�.�q!�u��ert�T7ܮ���9DOU}_}_B,�X������1ƇQ�	�b��#���!{c�ht������׎_f�\�D����:�ڶ�˹�\�x��8���n�6���bиt�:|���<��m�d�]�-<���������"�Q���J�����`=�Ng������1d 9����x���@-��R[��w�=�嵵X�3��xi3]uq��9ߛW�2"u��7�9�V�M�|gR3B8��y��4�0,}4,�|�а�{�J�;��:��mu�w����f�N�esN,K'F��c�덇Z}i\�5¸/�\6_p0�K���i4�ȃس�!luā��5OcJ/�f�	rf8'���G���5��W]V:&����۫
n��c4��1ξ](�9{3��!K�۸s���nEST��q���%����A��)\��s����'���/]�7]r�,T�N��T������+=��\20 O��(pV�9�x�R�1�t��w2��2~��7�7E�9�N�˞������6,��ӣ���kw',�ٹ�!^E�k�2_m��E���^f�l곔�SsNhA-�m��8���76�2��eF�MY>�CH&v�f56O�i�򦮞o@>�����C��Q��}��ͻSP���ݚb�8k��UU}_4���<�j������������5!�K2���󕹯!��MɍQ=�
�ͣ��+��f��q�G�2ji�I�Ip
���J��W���Q�����c#%��"R�Ie��=[6^����'�[^X#M�%�#�ÿ:`ך�4X�������T�*&i�UF�%JF�7k�c��ϛ��.������]��c��t��`��c���r��͞H�Z�;k\Fb���ɝ��D;�S�;$n�h3L|�%�H�H�E墁��(�;wڶ��hu��±^�.9gܲ��թP�g��%q�V��)(}^�uv��^���u�{�s��1Ht�.:�t��m��<7��\vBW����{.��������d\Ku_GTu�<���#����}�^F���@�,u�B�~)�}�����ƜZn\�d���E�h	��}��ț�L�����s��p����>�{Z�o�ch��xy[;/��q�f!�>n��W>n��=fШ�X���6�V9�^�a=��M�ӌˣ�����x��*�(��ݤ�[Du�ћ8����	����Ӏ��{^�#�lS���ߔ1���0g.�a�n��R��VJuҞ���+��*n*L�-'ϕV�v��wXǻr���� w��8�q�C{�r��0:����﫹�9&C�vq=��Ϋ��%S�Ό��so/�O-�1�7c�7	��u����й�I��3��H܈ӊfo��p��9
ߓ��d5W=ð}���qR��n������t]��8	ޡ�л��R��Ļ�k�~wy�Δ��)��[��]Y�3��Jy7%�Fإǯ���U!�z�%�@�'�=3�%3v�N�V ��*�� 0��x��UM�N��{�X�5�R�Á^� (�lwdo�T��Ч}��\��.�����{J&�Um\�:e����=>�F��/�ȃ����p����M��	��{k:�p��.�m���S�?g���ݧ�!4��q7&��5&9���seܖ��sK�PC����N)�{��G�f��gPK��,D���m�����<�k����ޜ��kT���?�d�J�{Snw��/GN.�Mq��k�Q��=Pᚕ#�	t�^�!�Q�SK"^sk1�j1�Q�<�.��\e��#CEJ!ʆ�w%�Vv�x]:[5ǲ���LL����gY���w��P -��vh���:_��;��tY�&�%��q��ے��5���m�9u�Y��A�H܆��K�007���;0/���W}���>��\�w7O�-��>�/bݡHJ74��=" &j��ݤ'q����7��˰��^鬝�q��^K�/!d�R����ޅί-��Q:�ÒNb�4ܣ�{��Om���
Ni����M=�b^�J�۸M�f52�o3aH�=����bN�ָUp�pr�X�R�#�[,d	��NWG2Y:*4�𥻑�Y�_\v޼*�ϗ8tr!�v�`n�v&X+5-�R�ޕ��N8�f7_@�g)t��iO��?*��l&Z\��^�F���9]��^�[�0_�^e>��*}�FV����Т���pf�a[Wz����gl�F��7}/�{ݍ�M��'=��Q�ey����E���v��E�F��y8i�\{6�:J)J���n��:��Z�n ,����o��z�F��E�K��f�������↰�&�ϡ�l�5�dM�޻~[L���3����
y[����AQH��-X;`P���5D[��W+;#���y��{F�Ũ��s{WOWj����%,7mwhM��2a��x��h�7VnveoV��M����ͺ��D]�V^`:�3��=r;���}����N�Mե��H�7F�����a�k��u��d��sv�m�!Y�n�I��M�S<�wĸϺ�K�0ކ{��]���7�ّ	dy�Qܷ�-N�����u��W)9�I���")2.2V���6�b�������]�z��8��z���HR��˙K��&�N��*'B��_s�������^rP�'�7:�J74��H��[�_J�����٤u#��J�YZ�̵K�+!�T�QS�%���ܱ/1j�)�ݫ����#i�ڿ�-�����4�6n�N^Kq�^�'bu,ە��w{���˜�*6�]��m�Ց���׍���Z�U��A��낲��ǣ^!��%䈼��y�F<�M�OE'��Z���l�Q<"�J	�ߟ��.f�<�}J���S�
��o:'��#�ޖ�}J����u��пeo
\4��%_��˵Di��5b�Sbj}�J�z��"�r\��%Ӑf�+���EcͷPM
��Qt��:�D8�|Լ��tNd=]��a7E-U�d3�v��ز��ǳ��:}�y	�/��p2+N��9�>ry���u��%�ǁХ��j��9р�ǂ=�t��̚�'u��r��`۔w�ӑ���0��2.�˂;�j;	|1rVz��A�Iv+�F{����~�8U�'v���ykӅJ��U���P��`h�k8��Vm�2�[�5��t��웖�R�k�u$��XM�-ok�ˊ�:�&��x��O�ŏ��ב�x!ˏ4z�Ϥ(2v�ۍx�a�]��.�ݳS^�"�<|0�06B>p-� �m�`��9�݄�lçL�ڲ�?,g�X\��Q�q�|4g��W����T��hm�H�Vci�X���f�C�^A�gv-.�o�^��	2m�P8f�(�߶"�
����b�ҘjWv��՝�u{�^f�̝�ٽ�[s�YU2��\o���s�;�����.xt��g��jpm�R��|��n��[��Ulz�����Pn[
H�q)S�c
E�Oޣ@T�}[�J,�����R�Ҷ��l��Sk�MK�Q:�j��s/� ����d�X��Z}���Q�A��V6�Sr��,qCh݄x�
��1��&��%$��nŹ�
��o��1>�<��=��:���6;Gp�q.-��o:���Ou����ՎF�_T�1�2ND8�D�y0�����X��R��ۚ��c�&ԴMN�L9�"����,]$�ַZ�L�#;q+Z%;]9~Sj�>��\�.��pgHu|�Fb�N���۽��%�i�yv�0a�)Wm��\���:e��i�[�L�v���m����v6qR&�6�Z�|��qK�u5����B�G�WF�}W�
�L�p�u|�d}���'&A��Ғ看�
DZ0�w�>X��\����nਜ਼����p�ץ�/F�4?����l�K{��d�ɀ
K�mۤ7����g�L
Oh^ц�tK��`�h�ɀcNXmȘ��[Sf�&F\��m�g]�,r	�waX�I������|�a���bgJ�x5y��t�S� �*Ծ�a\�@���[1�i;��v��Nz�dǜÝ�r��l^'�W)�k�	v�B�prQe�I��q(Mw-��׽��)���闥E��v�}޸_2�/h�$�y�I�<��-�\�管��|0]�bB��n�c�B�
22��otzFD-Vu稔�ĺǞ(��WO>��]쮍O��_up����߮�Ղ�,-I������*b����A�Ë�o�����)�+�޷��vn9G��͠�LC/�;�K��@	v4�uS�7L��R�j�yқ�O�$�k>j����\��e�aU���o+N^��4SD��n���Yf�wU"6�J�H�B!
�hs$���4M�E	�eȬ�w;�i��s���Vb�OAq)�
�$��;�qs0�]ەE�X�9���Ъ ��r��������Т���YXNy�U�s��!��,1J�Z�%U.�^�bDY*��wqZ$밣�5L)P��C��aiwt=m�AO;���rF�ȃ�i�*��Z&J�RE�P0҈HP�Α'�NF'J�J�,�*�D��Y!i��Qf��	BQ�hJ%*U	�Y�P�j!�f��`�#��!4CKa*%��2H����L��$�C#4�I"��9sLC�FKV���ZKCD4,�dv���3�-C*�6Z��@�H��MD,�f��Z���4T��Q

C$N��dIiS5Ȋ%T"�16F�g(��5E:Qs$��������������z*]�������$�7q�&;�ɼ,:�-u���g������ufѝJt��9��@��3�-�깿���W�WEΑ)��5Gs�mR��kY�׹�^�9�:��#+n��ojl"�(n9�ӝ'I���/>�I��z�"���x|Bڝih�;�2�[�Z1R�g��=�g&�5�Tae�I�t���g�<�,��P�Wօ��9͓�}ix���7Wj���dhnn>ě�x�t}n�dka�{���;1b��u��1r�AWt�d��*G�{��4�g;`ge�ٶ.��޷�_>�����3�	e_ZOXw��7��%v�D�]��e�q��7�Uv�F�k�#\.��Wg�Ҋ���j��3�Kq�f�.)���)a0�#�+��Ư�����h�8޿����G�v 9ȑ��r���wi�!r�j\B��8�g�m,���a>�nu�6!	D]-��RǋUtsI��"\���������DqM%ٗ��Y2�Z{0E���ldÝ�:��S;�=c/*�a1�W�({����iǒ��D�:1ս�Rt���J�qp�Z�xeXI��e�VRf_X|����e���3]�f�
ޖh[,u
A>E
M�F��j~J�Qg�pӽ�����n�����D}�|;Qm8��d]�c�R���Y�z�	O�Бui�/��ج�q�{��bOj]<c-�n@�4@�*z��ީ��5�vy䜧ϼ��dO�NDY}�]鬝�q��j�q�]ls�%I����oY��EԲR��[+Q�P����#:���ݜ\���}C�U}�f�}����t'U=�շQ��p���A���=����z��.e�hi�r��y�wl���*��;�ۄ��:����4zw4���^B�|��e����;;M�o"�U�+�ާu��v�ʉEY��ȉ��l�����7.�o=��:��7�Ӧ��C��S=�������j�=n���5����n^���{��Ʒz4oq?T=�׶6~��Kz���Ϭ>׹��{Ûa_tT|;��]�ьڒ�5��e�{5�`7�Z���Q��K�W�~�ytkhQ8}t��^�yx����y�;Y��IA���l��ƴۈs{���u0�G�RV�n6�v3���.��qϻ��J丠�������xi	�{�v�j��b��γ�0-��y.m۪�5���jg���"ś}M�eq]���o�n����g���p��O��q7$���c"U�V�gj�_h���Y��÷������o_�����+��53�p��,�0�n��.#�j���s�ku7�&��>��S m�^�b�z`oL�9HZ�9� ����ף�M�E��n5�4��[��6�z��=ӹ�����ob�v�D!(�M%&�zf������������|��WMg4c��V�2�^9j�U (��]Ĝ���SGE���/����Z���'�90�tRsM���ds�%Ot����ktr�\�t��s�����-q����iY�N��k�V���V	�� �6F�X���ɜs��Gw �,�����ׅS9�.p辱�"����hP��+���j���w��=΅�2���.)��kg�ݙ����o���N�R���'E=�"Y��7	�`�e�K��Ef1�t>��Yq.���s���	泷-��vz��vJp���SãC������i��� �1��B���gR���Z��2�u�E���=�[]�����u�W۪���r}K�}�}|�vk]-[�M�U����P|�Ys�.�}��e��'B�F���5th-)�5�Ts!����w��D��ǃK�̀�'�S��K�o�c�o�+J��v������v�g��r���6���GFQ�ԨC�#TNe����m��]T�������↰�m��e���
]4��;������_cޠw5��J���ks\.���잹��5E!R7
Pu�ec��P�eW�@��Tu$���)�{�t�Wd��h]e�n��Gc�=;n����~f�����]ZM&CZ�E�S�R�k��o˸�=���ns��
edA��G�.���-NT��]�j��rZ���/o3ut�K����ݛM�ۦ�;I\��7{o�k}����֩!���un��a��GYE��l��x�;��HE|T��ݔ�*�{��[![Z;9����kB�z	B�Ƨw�;)���r8�� n��݁-�{���̨��_3uw�������5�oj�RXrD�(�D���̴�������f>vi>'xepD����#|���H����>�.r�in�����1�j�T�����y����s����/'���v����f���ӗ��kŋF��EeM*�W^�zu�:���ܺ�z�NTۻE�f�\��m]%�� �կ,��g��^�ߞG|��O}�Y�hͧ�l�ޞ�ysZ�^߾y����ԓYش����Q��:�U}�u|<��§�V�ю�;�o��ŷݖ_��$�X7�+{�T�}MQS�i�֖�& ���x.�kә�J�7��E�4L�q���79��{l�>!N�s	8���]]����j��q=ܫk�&�%���XTZ���g�>Y�H�r'�;��J{�C��*��e����r��wW�u�K#���ܜI��x�+��78b�i�ì�m�Ǭnٙ�ĕ�t�g�(+J��knfq���ɾ��i@�~��r��7xY�������}s�$d������M�����A��j���)r���l0VQ�6�)c�Z2��LRO�=�3}��@!\f|���Į�!�����s����ٷ9������5:��mŚ0+��g%�AM�wF�w�ۤ�a�Mӿ�:��T�v�2w��U i�Fm{���!gL&�fv�]�s��>��1��Ҹ��~g~
��,�`˙�c��,���Gu�ȅlՆ��Z������I\Mʣ�.�@uP]�>��h3ϸK�m^��q��2ridK�]��N79Θ�.���D'�\x��I���:��꿣����Qe4��-K�:�r����W֮+H�c󵴹h��e�\����s�>�_���%5��H�B����������f8ٶ�}rR���vpS����\7�b6_V�0j�������s���8���=.h�㚺�x&��Q8�����)�f���r�.W,8v���.vr8tq������u8�Z2�ԺK��U=�����8wq�3��sw�m�(>0�������b�ȥ�ݕM��C����z0���;F�N�G�ǳ<�.��{�)t�[���������d3]}Z/���qq�Π"�b�qfv4�ȭ�﹛���0��,���eQ���}�HݪꔯS�jF�:o�p^�Y��ޘo6�e&J��Zwg��1�<��r�V�;�PG`K��v�V"�ۏh�҇r�ӞU�/�����q4�1m}�����f��,�[]�M'+e�ae��V��G�j^����M�|n{W%rim�T,�	o_��C�U�5�.:�5�)3|�K�t�֖Q5�U�7��V�7g�!��v�z�u#�Pu�ה7� Q�Y�9�6�[���M��;O�_T�iL��W;t�w����w�d�G�YC�\,������g���L&�`��&��-��w4Ow+}akT�#s6��8�\pMb�ݾ�	=?O/tT�I�KLxƷs-zy���5��M����@P"R���C��jdXl�V��"�2.��')"�۲�2�\aS���	Ta*�2�N}���oQViv=�Wܷ�g���Ob/~��7�&�.!�
e���zD�\G��'��ƬV�֚N�]��=���O��ˤٖ�㗋 B�=_H.�1��&�V ����_�ͫ�WR�.�����G���;%d����gk6޲5���SoSf�g{1��+Κ*���&�gQ������2�	t7�1u;���[�.�AMǗ&��}­��:=���uC����v]�Py�`է҇��j�"2or3���D}|����d�ڮ��K��#��ue'5m�琲;T�>%�m��\�0�:43��(&��V_VF��W�wW\*�M����Od]��Z���f�DN	qy*�;���7)��Y�%�mc⩜���y0sɸǫ*K+R}�w7���Ԏdd,��KK����s�iN�Y=c�Q��Թ���ӕ7d��K!��O����v�<���[�MI�t�F��y���8�l��w��0���Wbh�9Տ�$�jܸ�p=��G}P�k�S��&8����Y?F��ܧm��g`ۋR��zk!YU׍�(�!e���_[�����F���5��g��]M�=����/��EkF�ER�.5 ��O �qIZ2���[�k�Ǯ�Em��2��z��_"-^�jDܺ��L���eE�ZIu~�o����������6V��9�r`�w�Y�����3��Dt�]�
��F�[��6��Frm����%�_]�ϳ�Sk_*a�VR�ÖvT��zwJ8��S�<��躒�m_I��q����.��z�/�7R�U]� ��k/MH�7����։�3ۧ�+��;ﱙ��5�eBN{�	,]|E�q���':�k�h���V������z��a2����9.��PU�ھ��<٤�#�gy�$��4�%�%�/vns���0��)s�Z�ͳ�p�0�\+E�����(��j%��7�HA�O��e,]����^�'�~t.*;�N����=d&ٺ�-9y-ƺ��n�6��G�	";��|N�����{U~7�e�o-��?�WO�B�G�:�n���Q�4��:~5���=qU�t�'�m�/��8�fV�E+W���q�/�j6r8tq��yU�\j����n&�E���5IH���rn��ϕS��kY�׹��x2�N��l]N�;]�)�s��kvZ��)�dD�3�T�Z	�N�v|��dvuc��tHCg�P��	!j`*�lc��_�O�k�%�t��[�f��1C'��l_t#�d[/&a��=��(W���mN�}�%�깖;��N�P)}]����+�4��������r�hsš�A����;w�n�7R& 궍�!� UՓ!����]uQ����+K]�ا���N�A��ɥdhq��+M�C����7����S�'�O_n��jQ��ȞYn��:�%����M����&��R�iգz��.�����3���}t�tjV��}����S��ɣ�]i醷>���v�`�7rj
��QK*�&��޻���;Vo�����1�_]Ym�s��>�]�����0ƭ�ڏPñߝ��\���Zz�<r_<v�_����Z��q�x��J�&�I���U��Ji�ܙ�ݗ���t��2ridK�]��w�޵2���'|�/��mt��E����/�>�E���5�4��e�������7F�8�&�r];f_��:@�g�	GN@\��;]�)�4;j�L�]m�\���q=�Y;��{��n1�Y * ��	����,���+b6�������mgJn�%K�������bԶ�Z񱡽�w.l���:W��}�t�b#w�e�{�0l4�5���M\�e3�BH+��_7��,�����c�e=���;/��2�R*���ܬ�X�(��O>5{گ��7ݓ�B46)�(�<I�-�D�4\����+8�	vs7X�E�D����Q�=P������\��7����S�}�G[�٬�]0�Ӻ��}p]�:Y��ѝ�g�u�;|g"S��=c��x���D���t}^�W�ް�p��ty����Nvz���^V��Bhf,]�G%*�X�4Lyb}���5KZWǦ��^x�IT9d<�~�^�#E�7�k�b[w���R�F#L<�8h�I���۝qwK�[kIp��w5�N��U�ET�tn���JN.�f<��u\�!� i�΃���V��c5:w��n�G�����RrD�@�M���2n���G,Tw����F�AwD�X`���q۾CZS*������V�f�n`k��'��k��f�K���h���X���u�Yb��Cj�R��Sna�k���Z~��;��_J��튭U�Ԯ+�����Eq\�
;� n����v�6�;�cs����^Q�$��eMv�7G/6�v�Ǚj�fH�3������y�ʆ�[w���+���A��l��{k��yѺ��.�»��ΏzZTgh0:�AJ��-�ӕ�4�ZVh�$�W�^�X2�,{\Z���K��ˈ�ӳ�l;z����-@ys��N�\���_n���\n�1�c`Mo3�v�3il�G �umvt��H+G8J.�&�)�G���ƪenM �vKq\�sc��ھ�n�h(^us�T(.5����B͹W�[V�79L�v׸L����py�"Jd���A��}�L���<�TMp/m�B�)F�ec�7�WWA�#�4�vɀ�N�+��!�[w;dyy��dF��3����o9B�r�ebg�#�}\�����iE�܌+Yّ�Nq�Tن�̜�[��LV5x�����+6�;�t�XlcJL�Z��2��A�N�sG.;�3��DF1��e��_T�S\џ���FyP*I�X�\|OZ����zj��/�G,c��c;���-�ľ�J��,�;f��c��p&���U6�J�B��1���f�G`x��Fu0>�ڥh����gON�v��J���#���KH���t��u�<[fU�3�WR*	6��u��B͋�_N`�e�#{��|�S��5ݮG|����4e� ��j��]��sY��֓[M�q��BX�Ɂ)��n��3�s�Fcȸ88Ա��]p�Q�~�N��%������ۯ��lt�-_f�'�UR��x�^�b*f�ufi�j�[L��]"^��ͬ�=B�6�nbݐG ��kL��=�$F�Dӡ��&D+*䘨�(�dI��,�KBȌe��e��NUJ����U�T�,��TL��-�%	����)E�r
���DUf(��F�"*2�l�Q�Aeba�&��$����.uj!e\����U',Y��i�+N�E�0�mM�"�4�˕Y����G�A��a)d��k
�̥eZ���U�4X�����G!"ʢ#2�Pβ�S�v�YE��T�:�Tr(L��uPȹr�RB�3et:\ ��I�P]&���(Q�b�NRBEP��SK��HL�"��\�$V�Ц\�C�ZZ-BV�ӢiY	�Z�H���
�* �8D����I�,#6�TT�Z���Ĝг�+�Ҥ����I�/����>��
ʗ����4�28�9v)v��q���P���@:�f���;�}�'F���������WtZ��Q�a5up�����s�Yu�M|T�����ivzvH;K!n��*�y�����>�}q��d$��B��C�<��V��K��K"�J˲��&Q�$�tS���-�K�LGrw�z�
�r2��6:�ܪ=-�����f ��{/��9��--��};�F>��s9B�e�|�|�!{���ݬ�-㈵�E����;�As�aeK*������,\�=�[^�X�Ƿ���Sf����u���,q�����u�kt�["�Ν -.qoJd֝���3i��a�g�����v�z��H�tM�h�Tl�E�L��qN:�7�jv�877�c��!6�;O�_Wё6���S}t6�k��>x�2+�_3�n�<9�\+W\���܈��O��<�b�i
�`���s��N�pO��$�.8$�u�n�T��h�s��>�w���n5Y��B���c����Yo�U��۞&�����C��n1׺�d���5kBv����aKv����r�PY�ʵ���N9܏TM_��:�Z�]�>S8�a��� $o5�:�}�-n��]yx����7Ss�\emr6���=�����e*ǖ�E��EI�x(J]7[�q��Ȱ�-pU9F���밽�<:�8��鿱����
ea��%��%�|{�!���]�X�����q�nh��^}/9��^��obݱP��(��	���sTlf�cf,�=���R9�*���Quq	�/"^9y *@QS� �s�ss4���]I�֑��{W�ǫ	]|�w�f������m�<Y��"~���z�lb[�*q�:��'(#��m�՛˯��ĝ��-p�67�u=-Z������\�72Ŀ��Q8����!�i�Y�%���z������4�<Fzyv��Y���!�2���|-	��eOm�2����Y����T3v��� ��k��������|.��T?_2���Ⱚ=��s�g�A�D�KN��+.1Rn]bO��^�z���r�è�V7[t`)��
'Q�]u�y�u<I���F��Z�s��z��n����'=�3�..�Zv5�T������L�}���Yc3��,��ĳtW��9v8�܋�Y���-�pݖ����x��s�Aئu��o�S�X���Ȍ�ۜ�r��}}��+,�W��v��l��ܲ�s�;o����a���i#p���>�u���!�S��fTH]}t���%��d�/�P��Bm���|Di��W����R���6:�gXj�AW�F�A�
�+F[îي�0���d�X�ϕ��]�Yڵ��$��`(,�����B����8�����#�xv�җ"oz��a��q��J�nI����JNzRXog\>��jhV�h`Z��a�g4^:�B��'%k=��o^7;:B�BU��5��ݮ�Ӭ�l�M�p��݆8ޢN��y�l��M�t:b��k�ԕ���u�:1ͥ݋\K��W�_l ����(���̼��S����(��v�(��d]�q�\J9��P|�)�%;�惸l�_�'-�r�ɍ�oxԝֺx�^[��M|\�D��/+��sl��庞T"e=gm�,�Ý|J�0xY���}�/����U��4��.��A�xy����R5:�T��7�fb'�p0h�ۗ�<&���]�n�"9�y�ԗr���^qv+usV�!��̮�؊`k��ͮ�IpYέbU�+f_m�$G�U}_t�\��w��v�4�W���e�s�5�rj"qtm���~�E�i^b���R�2�Y��:*=�2��_Ż9�:9��p��R���cuZ�)R8��rD:�XB�
Ҟϻ����S尝��{�]�3���nk��v��\ˏ_WzN�kӫ�V^�Ms�ϴ���e����v'}���BXz$��>
��(]�Ù�ݸ��U���P�}��ae�I�P�.2��Y�_�n2�Oz;}�6�ҍ��9u:��P�K�����XP Y/i ��9G�F��C��y�56���;���������@���D����G-ϵ�[�kl��Qy����S���2e�ዣ���+����`�u[�>Ϲ�]��u������ܚ?3,I��ؽS��sԖ�<�D?��(�����٫��+Z;�z��nv��H�&�z��jT��q]}�_dʽ���=��6��7'\.���`6�f�Yk\��{g6�l��(u����7��+�-,�SaX�-�#U�l�D�^Ñ��,�X<oi��6�5���3�����𴫏��9���rFv��͔�a[W���|��~������C1�G|�2�NG��!���S' 6�;�>�Ǽ"{boMf�����'_�L�va*�� ���E���Q�Ҿ�,�4��s����M�=Cf��)W>+�<|��C=�O�}Iޟ^�F����2�z�k%��-ʶٗ�Kq�>Y�H
*z�'���֣�ҙ�Ջ���ܞ2ںZ\��7�����&��qR\Th֯�2�h���%�s���d$��˜{!�����\As��b�f�E���6<}�f��U�,DUM�l�}���:���[�6;������u�\�3�L+�Qk�ih�e��C���v�R�YH�x�g�<R�B�9cI��9rW&��ko[> βU5��j�o;��U�����Gۆvo�ڥ��U�����sr������jԔ�ۃ�[~�oJb�ь#ѽ?9����+1��{^��=QBsx>� d�mm�����ۡ�E�ZOր�z�[}F�T�B����-�-�X���j�3�o�C��rƭk��b�;O�.�z�qh���u�x����κ��S�N�u����Z]|z뀰ud���V�����¸���I��x��g������jg�[�=�Nou,fy[Djuѫ�j���g��p���8�>�}G��Hu�)�5�D��;��Bv<k˧�!�_s�g{�+�5��jen�Cnoj�Fo��uB�O�_�r�L���I,\pId.���갓܈/Z*4̡��ų5{ј븳���Gc�=;n����Q���s�kv+��� ��f�����|�<��NR{�*#��{����˰����n
<7�$�������s��ZJAwq0�R��-7�;b�	F撸�霽��he�nrJ��m%(2v�S�:����������M�y��W�PT�dc{���R��m���ۓ�G�������O�-9����C�W�9�Q9x�
QZw�%ۗS���9P��OV�v:�s�wy�]~�Wy�*�y�",�M��.��6ݽ�ԗE��}���=йO.�5k��F�����n��ycԺ'y�e�9�3V��k���z^i�W��u�rz]-����c�W����w�]�jm���1����&�bb��kK�1 �Fp�V��:�����|�e�ϻ�^|��>��j�)�C<����T�z֯v�:[���E:�zv�,�T*/�oC��b�Nt�w��V3t������V�\�OX��I���'̦�o�v�˂�v�ʟ.X[WW��4E�z���J��!����&�C�\��1:�ǃl��{�d��P�|R�=n$�}}�N��s���v�g��v|��b:7R"O�aF�F��j�*"G;��W֡,����ܜP��&�]�=��m']�����R�����?����;��kW��{s�x�������Va:	~틔m���ڑZ���nM2k�D����I��?m{��d�bW{�4�}C��D7vk�׌Π�Dܓ�:�9����"�j�%��������w_�L�'�Z�'�1��t�B�Ď�5�֑�8�+]�@k��Uݛ��H��~?^oy�h[���T�y]�@y	y�Z�t�7�Dl�viII����#g�����2�-���k��u��.�fK&f]��H+q�غ:�8�I}�v��\4�
t��hfk8��ZhȎ�o������Gы��{���8ޢN|K>����ݛ������]{�ʭ	G�~���=Hm�)�C��h�/J޲8��5Ҝ�R�fnh���algir܇LE|\�D���W:1��V��A�f��-��I���[�ѵEF��>��x׍���mX�^��摥��
|�kY����;�OCݞ���ĽF��Fq�!e�s�5ɩ���z�k�V\����\��
�/O-^�/��X�
vs������UG,j�S��=����6.�ޒt�9n-�LΟ�����/S尝��F��x2���������/nd0>�8����*7hԷ|�Bw�22�+��i)��<�֑��}C�zr���ίq�ⰲ�+M��@�#CQs;�����rV^��Z�<^B߷��~r��ܾ�	gh�9���h)������G�>�P��1T{�ɋ8�����s��A�-�U�L~b+v�G��"Y��;(��� ��Ǌo�e����/z�D�w�)���q^��u�\9�jFA�����ޏ4�@x�g�\�k�ܮv���ķx-:.g6L-��F����%]�[r��Iv�l��k.�!�O����@�b>]E�dw�甥Igp���ϸ7����[e�z~��������
R�Z��~�%=��w����_ܓ���5ٮ\c+��{���-{Y�����(�o������q8�_�B��٫��ұ�����5�\�;��wn�V�*q}��R %�}������L���P��݁�'8*�i*�+o/���Nۤ)	G䣧�}]H�S�j#����-�̥��XΣìuۉ�R�%▮6�_��	C���7���$'���:�qn)�gu�G�������W�2�[�j��n��n���e�)�M<��qm��=�����mUZ\�n5���M$Eu�N�^a��/�>(��%c�k�:�u�Ϯ9^��r�
���o*.���>��4�C)�_2^x�L}�|2�����U�t�Ǔ�Y$��
ӕea��#,�6:�g�{��e�/7�v.���{��g��ж��w��qQZf�L&�=�Ɩ�	]&���E�d��E���֚h�3��AX�t��H¥���!�ΝEG�Y�U��iv��F���[�m5�Ƨg���.��G����˱�wX�yc�Ÿ�KKD�%�a�?^s�iN�G��h��7�E�7v����ʛ�CH��_vDvb�z��n�D=���o(��XPW[�.���#d����Z�r��{��b�����E@��⇯���7/��C��
�+�+>��l�%���;=��}��iL��ӯ��Z޻�Κ�6hum(�������8ks��9�� _dm�K�a�Y�(�h�h����=$���4��p�]_&�>�p����s� �J�y%5��r�j�����2h($�q�%��;v��'�UZ@m#e|Q8��n��N �޼fv�RWMʨ?3A|�Np-n�c���眎��L�P�4wv����K�{S�ns� �V���r %�����݃1AW,�c���1�X��ui�(�l�|�,��h��O.^�N�w���{6�G��fP��O�7/'nK%�� �8L�һ���7گY�(�R�Tg����;�Hp��٥�vi����LP�׺RVE�T�pU�J5*]6
}+WjGfԤ0�	�j�]�uĖ��Zi�D��)b}�K9J.�ۢ3��Fky5�k����#�r"ͼ*9�;p>��}�� vb�.�j~�w*��b�/��,EJ�ok�7��ց��j�ɯD�M-�0+'.Q�,D�E�L-T�_Q9fdf�£�RLФ
t;ܸo3��A՜��2���]���pMU��~yHޥ�~[	漣A�v�B���F�~4��pj݀���m�:�#R�U7x ��ӝ��}�	�C�[��x*�8�gU�T���7Ж¬U�r7O������9�|N�i��GL�/aї��e�M�:I� �. '�e�i�W0-1E�or�"�'44��b�M�u'�)��GU���msCUYb�8*Y��:�s��^�[S�ݺ4j��	���}�G2��+��c�<��#����7��m�2=��O5�<��UHrݖ�[��SA\�o.�Ƴ��
���*V.��[B�.fS���`S��&�}˻�o��m���OsT5sc������na��i��㌣4t��uozf���u���Y���L��f�ظnp�:gS�(<Q�m/�*�t�n�)��m���Ԉ�;��b8�����T%�/$uB)m��V]��v�>Ѵ-}�G��n�nY�Y��*n���衴%m��RX�O�fa=Է��X��Ӏ�9��P-�-6��Io1�#�mA{��]+�.�)^
Y[[;��U$�)�X������fK�F�-9Le,�lf��V�'km�dʝ��}�ݖ���6�Js�V��OT��j,J�>�׎�ԓKg$U�}�������7>h.�[��n�W�\�M���K��Io� 4���FDw��,��>�(T�.�`_uVw's�=��t��M�.��n�;ud�\�
H��tI1fj옅E�I7���ai;K���ȩվ��a|Z�r&�C��S79d9�o\������bݬ�op���ᓅ[���R�'�����vm=v`��\�u�ݞ�ݟ��B����x�܃U�v��@�C>��v�Y��z��������v�)�=��9�{�iX�^-��w��<�TX��5z��Ɯ��V�o{5D�K��v1����=�ƧG���.�Ț��
�"������'y�3��5|�E�uu��N����4����TOh ��:nS�����3���ξ���,-.h�{��^'�u���n ��6O,V�R�`�<Y�[	�<'�3�q%��=U��O�4�Dkj�ZŖ� k\��}��kUs���
�-P�>�wY���T�.�}�,�TY&�{�ko��Ρ�0�3 K�`��#� �h
$�
gI*hu1	JJ(�I�$R+-%,�	W+D9�ND:����bQ�\J��*�.��.\+P�ifDQ���(4�Bh��rER�&F�&RI�Εs�b��f���F�a�Da���TQ�DP�%���a�j�Q(���(�  �V
E�Ԃ�vd$�X��2�',&�:��TDZ�PE%,��IP*#$��("�*���6��(�A0�$��B��6T�t�5Q""�ɕ�.A���9Z��`UI��˚�Q�9rԈ̂�V&�갳�TD��(9QTPE&\��օAEʢ��"�&FdvUd�	TE��
*"�m4YU5�QU!,�(Q%����J���S��QEU�RA$�,L�5 �DUH���K:��:E	&\�WV��*TTWY�*�aU�B�(�Pb�E�A����ó��01�v��M�wmf⼹g�4p�g��K�=��9^*.ˉƸ�ܬ}ݬ�ڮFu�j�bN���*�_�����,r�[��ͷ�����k#���D���%��o#����M$۹f��B�^��ܭ�<�	�n�;g��x�oT�f^D�r�@�R����p+v��-�����H�y �v����ö�Ֆ��n5�"�ɘ�ʞ�>l�NG|�Mx����}xz��wr6�������bN�[1.�${������j5f�{��s)q��]DN.�����|mw�%�E
�.��\��٬��X�a�'�i��G`��~ �.��U��K��菞&��g�ym[�Z`�
Ý%�ɾ�,���!��k��ͣ�2�ݗs����J�Q٤\kvZ��)�g�L��
+.2&����8s����P��C�%P6U6��{T�c2%<���@Pэ�nJMˤ��
�u��\�L�ڣ��r����`7d��"yg�t�BG��}���P֣}кܪ���(ɇC�G�D�I�*���Q����p�Mo���I]�@���`8Nj�ShLh�������}*�݋��
�)���o]:��u���
��;E�m��&z�\ee�9����f�z{�IO+���h\;WN�p�W�y�w-�t�:bJgu��A=����5�FD�]�;��;α�^�!滟bx �n�'z����]i醷#\.M=?�'"
�4�Tu$��U�9�d�.��@��E�m�|\5ٮ^3:�]rk��5ٷ�[u\�4��2�6���+>}|r�!�I�������äʙUfgz�ܢ�-#�]ɖt�}�5���I�	���ؗ�7	����wB:e�Sg[mݬ����:��nzd�Ym�7q����-d�e�B���I�T�-�.+��͸�
��*z�Aqׁs��G�	N���J<#5���}���{��w)���^}-Ƽ�d�IS�\���sl����Sh���	��z{N&���Up��x��	.N�.��;Z��չf�uޛ��V�5m3�K��E:��.p���p���>��^0��5�0��dWuiT�\0R�[�o��Ӕ;�d�}��l&O"Y����׹��3���{rɧ�E�M��]]图݄�G��B�Ľ�GE�4�-��Igz���7Z��$�����[�qM��=N�l�a�xVwQE��J"�	�����;�+�A�g���N�l��T�jtZf��ͷ��w�dA�m�/��p��L������b��&���*+q��*�ܺ���[�y�w��+'Me�|�a�-����q����P�ˋ/�;}3P'n���%�������W��~ȓ���_��Ϩ�U��:��ݞn9Wm{=֎�::Ӗɭ;��F�Sq�7����}P{�Z��\I];P*[���H�eq\㲁�����kr5�s�i�@�6�neN�tW!����<Q%>��J츃t�ߖXn�V�$�9�]�k����-*w0�gb�v�
�2E�����:RK���>�lԶs�+Z;��S��8s�ws��gT"���5}�i���o�kv!:�����g;\Et(�\ټn�O�L�鿱��S+���V�|'�mSޞk��0�=���o4�4�z*�`|��w*�����y-F�����l>1�˧.������MM;1݁tFvؚ\��Pލܝ��d��cwҬԱò�ر.J���M�E)k�uG8������vٷ�t���ejg^
p�t�
6y��U��;��l�ȗ�nȥhQ8��'�|:�w���SW�Y`�ԎS\W45.t�6e���!R �툐��/D����6��f�4�)K*�{i���9=xں����&�Y�e�<n�=���X�=�p>��>�ީ�=���]gs��z�vs����8qT. v4�� [ы�f��eɯ�q��R�F{#�;����L����:v��Ӥ^ع+5!S�#�U<A�]ih.�wU���K�r4�TI�g2{�K���B}�����;ݭ�e��u��p�(7��D��lB�Sohݔ�(�+N��12��i��z�>-�s�3�mũ{�K�5�n�&�8D�fz�u��Va���Ɔ��M��l�ݟ<5�6)ӭc��f&��L�;�s8�[���uԠ.�N�Dpnq�XSl���{<;��WY�p�vwlf(��D�Fs����/3G��(;B�Y�j��yUs=��o�
��Ԩy��,��5���ϰ�Ml�%Kg3s^��:Ԉ��,�I�+�ƭ$��&�ޠ�#�-rVΆN�s�����U�(�éƬ��鞨K+�|s�V���}�˻KX�V� ��m�Z����լZW7&���Q@�Ib�K>]a۷��mJˍ0�u��O#;�Wiƭl�s��fv�%sr��ʄ�W��h��4�L�]���)_^�^�6ND�g�ݓ��B��G�\���z�n���Ը��q���SK>����/vo�M�\;b�BQI���;>����l)@�j�6�v���#�⋤ٖ���^,�p{B�ؼ��m�����9u!7�:�������0��nmOw�"h��M�s4g�<��s�(��ؚ��'\K����}[�uU��q�;�Z�u�r/�������yA�m�돎Uj�5�����6)��Y�5��2ix�7���V'L���>��+����;S���K��p<M��}�4H�/a�E�e`��r�E��f�o�$�L[Q��X���?J�n�,ö�&�)�L�El\�<��۶��Z�B^��*8��O�ゑ�'Qjʔ퓃���x�>�o�V���ʋ�y�c+ەY/��.v�Tޣkh�D���򃧪�KG�����S�52�T3��G�e���=���ҳ�v�Y��c^������Yṡ�Dae�ʓs��v&�ȃ�=�o'������ٽ�%s]Ø~��-�[��ȉ�l�&47%&�|�֯�D���:=\���y�lK�jo���%[�F�ʑ�㮝_�j�t�hnv��
��T;zX�8��;�����pJG�м�gm������Ƶzl��8{�s9��ap�5��y�幮��5������srh��A|ʂ�t֨��2�vX��O5��}��{�,$���\-��wܻ�PcUo���X
s���-�gD��2�+��L�铑+Y��8޼nv�t��|���h.X�:�f�����M���!���IȀ�Y/9(y�����O���~��R�s�*��6&����4�҃z������g*�bf�����%�W�&�3@�[S`-P|-'�M4in�{=�Xdo�5��t��,Xg픫x*V�-oAK�[�O"o+	i�.`W�|��7WVI�2�C*@��%���RԦ�t�z%�^ƶ�A�[]�l ����.|�R=�m�5:���9=��f��p����hWg
�����Tί��G�	O(B�$��O�a��7�½�ѯ;��NZ��^|���f��9��+�m�]����_gf��G̷+V,;N	=q��$n��\&�B˨�x$�;8�"��1GGNwQ �|Q���{:�gI}q��
vqs�G`뇕Q�c�W��S�&]c���Gԓc����o��OJ��3S̵�͎Ȗ�:�C����Vk��nNs6 %S���Y{�E��Pwy
�7+�bW�������n�p仢�m�!����o�w#��ʲ.^cnF.~�P{�[�g����ɭڣ��Js�m�s��]1L��>�z*9�?4/�y(3����헧;J��s�ml�6�Z�6s�e��jg��u�wV��5<m.e����R<�p�(���}�hk�{rz���ǯ3�7m��a����t��M����Xа+���y��jcM�ڳ�jv|O�Qf��f�ݲ�o^�Z���)��#P��xĢ7���I�����:�J��t:��VWL�ל�&�tn��#�T��X-��Y��cFޕ�nQ�w>Ϧݟ}C�U�{N�7���t�9'���p��2���l�n���y#8��P��_�,dpIb��٩l��N^#NB�K�+�[��#
��M\ܪ?_2�N}����L�V���7�w'S��Gy�u�]�8�k}�q�ΰ����	TD��7�<óyo<�����z�3�O�c���6e�x�ᬊV�A;���M����w)i@�A�۵[Y�NN��\$]&̵-Ƽ��!R���5UTE�J@��N�sͱ����(&�~;<�N��'��TaisW	�琲Ѵ0��P�LQN�Q>E����1��{i�l���|��+Ր����ã����U׽5\_�f�w����UĻ��|9P��]�4�r�=���m�\�l@�Jg�&��jӗ9e������ʨ/^�ݰ]|.����ֺڝ�LXW�����yp�b�7��ZN��8 �v����"N�xO�ݧS�^�x(������A)��W�,�<����!�6
z��%�^�{/�b	�%�[��o���{F���nbR�\�v���L] e���-��wȚnj�7"�m����/q'�|��	��!�������-r�8e�ݯ']Da]������_�Tae�V��X��ܾ9��u��U�e�6�C��Q�F��{���+뫎�	dG�477&�^6s�5�-V���yt)�W�5�w=A*��:����
�5;Y�p��7-��_k�<�����z��|��S=P̬���<���UlG&��y�;=U�5�gOwy���O���3�S��P�jW�j�a�ȯ�=޸Թ����s�G�5ٹ^��Q�\7�{��.���3|�Od;�/"FJfgʺ���ݙ�
�E��E�5x<2��8^xn���s�Ȭ�{��":���X�?z���U!��	n��{�X�ܫ���<<$c���b���b��������s���C���s��g�H�����ՙ�%!�ņ��ux]F�	�tйȅ����>��,�8��X�~���|��� �˛tTm��2���k�������� ��oH�,ӫ)p��up��Ŭ.bb+�q�'nֹ[�⾌ף��\�ۦr�l����>�ȳS�lG=-5�'	]�Ig�%z���A�p���U�w&��&��������̮HD0.�l\�쫷yY��	;_y��֠����}��{�<�#�b&���f�c7�/b
�' �eO�>��eˊ��
סcg�tt��{�ע9Q�>�cS��a9����݄�T1ڮ���.68�)N\���@n�����at���>��=�3+�~`y�����WZa筠_ظ>�)�	.�T}7fS��K$����T�Y�P�<�x�=���N��3���G��QϽ�sgմ7>�r8X�S�ȏ@�@���
&v}��,�J}����r��ʽᇱd{]���C�����<Ȭ��;����Y��P~q��F�%?��ݕ�w;����5��_�EIoLG�ƪkT�oW�ǥ���C�e���r7�ޚ�q/WP�bJإ�ߏ�{n��a�ݐ+��H!N�sׄh�s>{��2���H��7��/���UR����U�v^����̒6��9Uã�D<90r��2;�o`�fL;霭�_y��^�:�4v�m�����o���|�ي}'k,ͣ�H\�[2;��M��*6���u�.�J'~�Q�*K8z+G���{ǯ�7��O���L��zyEe�Y# V��
�(9��#���41�ֈ��]LkfR� �BR���e��2b݊���hMh���/"���)�h[w�g�ԼD�w֤�Ы�;Q�ش;�1*��h˸LQ���x��>��^=�<�tH�]�\A���e�X%�k���^�V%��z��t1�of']/>�R�ɟz㉦F�l�Y��0khmlCiH֫UwmycK2�i�`�j|�v-�()�{��L�Xs�G�VE���,g�<7��d��1��Ví��oT�Kz�͝+�j��'iX���Q��^ h���N�bsPZ�430�Ҷ��pշ�e���/�(Q�U �#$�6�����͌�2s�MACZ�2U&BW�1��R��畡�|�+� ��Ö1S�Q�N�Z>�"���Q�gvJ
�
�P 5����\���������Y�/l-��Py��z%��1��6�|�]]��0Q�r2#������s�4�joX��0��abڕ���K��ᓹA�r��	�p�Xy�;ғ��ƹ�J�(MU���[�0�Ud��EF.I���t,fCِv�(0ۙhBaYn�U��쭅h��؝��p$z�e:��q�D�:�����3u�{'�	��9 �U���u��ҳ)V�u!�IJ��Ob�!G&1�c�V��YQ��Et#U�F�%Jv��s;UL�÷o����L�>�z���9��ܨ~gR
�b�+"Py|h�
+�؝�3�/�m��H��؄�c%_u��y��p���$睫ݷ9s��=�K�|���x��V��l�f��׽�����;ᖉ��5A9{�� ]�5]4��)�j��v�#��fΰ��@o��VS��lӛ��7�M��Ֆ(��s�Aw�%6��J�x�7�cMQv��&r�R���E�D�|�Cm|���XNZv�ã&��ޭ�K�8�.Hs\������ �X�C���f�D?Kш9����f�����"��������c�{�[^�@�=������`����.gi�}R�b���c���]5���j�j�+��2����j�f��K6Ot���"�ʵ��")�,6My��U5�2�־��/��ei�k����]kn�\x��ع�m�j���Z�l����Pbu#�M�����W�ͫ��]+uȜ�ŒAJ؊=Xl���;5=3m��U������w�f_!��� 7�9�\��!��i�Yp�]�����Gѭ~ɈZY�,*	!�*y��m��j��Z����w˲Q�or�Kj�V�V.ͻڱ�[�Y��K�
��晌�"�����b�+X�"�������@<�Y�%p�������\��`�9g9&f
=�g��\���Y�5P���q;9۱P�-uY�*iki��ڨ�Yn�h��	[l������!�{Z���҆��r �&�ַ�m���C����;<2�B|�흱�Z��JvN�������?�w��*�,ʚf�:dv����ʎTTUE�%E��(�eXR�)2*���$ʒ����R��AT*d$d�R*��BD��2�\9U�(�5�:jU�@�ڤVbeD��JH�b҂�P�гT��QM�rP�9��3�G*��]2IXpH*"
�:���"�P�s0�SVi�F�EDR�ȕ��S�AY�U$Er#�\"����3����)�Hk(��KB*��Z�$#���he\�p�%[.Z�.M2��D�#R��*�D�*�J��DEtVP��\��QL�eQDQӘ�$�
�r�3$B�UȨ�F�*����H�C���D*Ԉ���4S"�Z",�9*�h*m(9$br*e)HEP��eK8AgZ&]$��EN�%U��RH�
*ԨK@�.TUrN�>0�  L��9�セ3}�[��v�8���5��ўx�mbQ�3���w;V�pl�mQ��v��{݆г��#�p|���Ծ�ʞ�?�- �Y˯���EdSy��S���	c�o�	�ul<�!
��jy��ns����K��L�H3>���d�ʆr�o֦��_�!����<}��@�{��'�;>���k����Q�c>ڡ��d�t$Kf��u�5H�/�k�؊~x�b��ar��)v�9�h��V���^�2=n���ɺ��#izՌYM�/���,�2xu���z����l�u �ղí���o"�W3��eCB쏠���d �3�PE���v{ҏm��O
3�y^X���G���� 3�ם���D�^'C���2��bK ��/�Ѳ�{r7������y^`�؎5�2�d{~��e�}�v2�s'�s&����W�!휓�����&�{�Z�K'=S~�Ul�=��3���!�%^# �vC����k>�����r={b�.�sn�n���4����D{G �v�+"z�}�W{�Ӱ�� �n|z�G�;��^��՞���T�D�[��wX��g�:���v�*'͇ۍ�[3���YED�LF��r�:x �����%%%��O�@e/��,�Q��yo�2�S�L&�xvҫ�B𛿳�vtD23�]+Y�9�^��֞y��b�	����u���'�wI������W�T�7��X=A�5��޶�|���A��:&����]�U� ����8~:s���;��y�_l����$�X��	���7 UK_�c��E��y���n�|�10��{t{r���0Q5�^�ϰ�������?e�|F��fN��7���a�������>�z��˨�e+F���ՏB�1)��5��{=~>�O���q��س�v�<{qR-������m�ƃ�M��N�<����3~�&���,�WQ�=t�sw�������|�W��G����v�s�g��'���#~�=��!�@�3Q!!�Ö��z�׆{=y7���g`�=l��T�_��D��]Z/�z���1i���c�<5@�jC��K�S�6���g���)�ȯygH���ዅj&��ݸz������x���S�fr�
f%.� 7D�R�}�\/na��iQ�����fK6wv��凞���,�}���z��>�Q���w�!�C���6	�4y>�xh��eKW��b࡝�.B~���Ԥx1�##��f�u�'\���!K�=n� z����_�K����JDxO�����e��ca*���a��������z�{��fj[����C�-�U���l�<U���L�R��:�a	N˧P+�� E6S�r�L�]�ĕ�ɫ�aH�6�\,��X6�窟r@^�|�LU�YC���:��fB�ŵ2'ư�LVR���s5ˆVk(eԺ��\�����:)1����p7s�4H�Q1i�`��
�>ȓ[7N�����-*|~�l{�2�>^�a|�^�>��k��H֎�K��;z����}�ǧjɯhs�q2m��ߤ����a�bخ���^��tQ:N:�]��M�Ӂg�;<��fa�?�U�f�O�w�c� �n}>��9䧷sn�g_��9ʴ��G����O�?��&��ڹ���6�.��m��.�TT��h�v�e��R����+O����w3��~���]U���߹}Э��[�ĢwW9e�]F6�/��7f��glo>Sދ�ݞ�CEטoUz&�W�z�Ņ��Ǖ��<��^���,���Xx�~���3?l�w������5N|n��Gw>u������H�N߇�ｵ��ŐN�qK�v�����f���j�%���A�W��@�>c����Ӭ�9��^���ȍ�z���kc�n��tw�k�r��^��3�v�dY���> fgƜ��j�Z�n)�<{�s���Pƙs���NwUm�Ϣ9�y�߻�2�?c��Vz��D�/�< R!��v~����MHm���4��v�4޹'�x�,3I�aݎ+sN�1��y���(�}ehs��9��~n{L5�����R5�xv?_[�e<��J\ʙە��k��2�_t���;)ovO����s�i��rB亮�3�vb!�ĸ^��Xʚ��fP�Ÿ� 6s)C%r��G��{�d^E{���~aw��3�O��22y�J. ܲ��X~�+�?ea��<r�ܤ.<o�G���.
��)DW����|�l����Odz�����Hc;x����w�%�2RG����=Bj)�22� 眎CYW�!Ӟ��C���h�n=u>�7��Eon��"��/���M�>|�ח/�����D�)ϲ;�*N&��#!����Y}Xx������q�4�]P����,�X�tx[��rK���d���۫*gm֓ݸ�ᬝ�s�ԅ׾���'��-N�>�Ni��#u���v���W|�M��d�U^4�:�M{Б��T���9�gW�yc!��e�?g�h�-���{u#���D�T/2����}|�O��no,#̏C��C�*�{;=;	���}s>�[;qG=�sqմ7>�r8y]�����{�<wUly�����I�>ȫ�Ho��8j4�2b���;�����K��G�dWg��?D���`��܌�~!G��G���ݨ�ȗ�ly`�M�8,��+����c����!�/�=��g��#b�dG7 W�[����qM��g.ɺ�۩�Z,��NVN�����E\�&$tC���D�����X��g{����p'B«�A���II�=T�K��0�݁�R��X멹[���⾩��Y3s;<�����yw�9��tθԦ蔕N���H�9�q�p{����[u�O���Nv�E�z���g�x_�Vp�zD��ϣ�'7]�u�w&��#����e�$k�qq�n�f�@�z,Q�&�c�;�m�o����w|vs4�D֝Ʀ��x'}�j�~�O��1O��B�ǆܨZL��wÚ��w�>�~㨓h�!��w"��~̇�!����O���d�!�ק�e�Q6�N@T��ｏ�G��g�����lzv˯���EdSy��S����K7��C�a���������%�H�ȡ�ϔ�3���A��r�������������G?T�-{�d�.1֠o�߹F@>۶*nPAD̥��&��f��~c�����R�i���va��շ��M�w�xv{�x*�=�d���\CY7P�}4@���V���1~�\�<�}��Ԫ���o�7�;>�Vzv�hS����^��t�,�WC8�~'�T5�L߬?u����gg}C���R���W�~�r|��s�W�3���G�"}~����ٚ��ʑ*`� ��,�Oz�k���]N��	���;�`�J��O7��8� ]]���A�Y@,���ǩ3}E�v�*�]��f�ۇ�HE�U�hM8��J쏈`X%�A�U���j�4�� �~vs�e���Y)u�"VO���nB�� {ڏJ��HOuݔ`uF��֫8�4����<6;(�lq������݅��\˱�޹��rg�T#>�˞���ب�&\�y,�t�F�Х�'�d��A���yJ�F��{	�1ߙ�_�-�ȣ�n�"�`=�+FjT��N�X�D�zVOWK[Ჭ��n}�{ǥ�{�;}(J��{ۆ�Z��ݜ�C}�M���({O�̅W�:0�JN��/���ts2R�T�)Q#C�3��9�u�z�����%�
�X���B�}�ܰ����p����cy�{��^s��Zw�$�љ�L����~��e�|F��fK�2~�[C�2�C(=���2�P�w��GZ���Q��o[���S����xz�k����{r=�=�='b���5�:j�<�����R��� h/�M+��.�u��7y/`�_�oz���߻���Ǒ�u�����;�I�$�lo���d	�)��G�rn��J��u���\�Ao=&v������Y{�n�n�o�W�q���r<tV1'( �f|�9�!/UI�K�r��}��7>�
pK�>�f+nc!��z��]*']��]ᇣH�4ӣAKr�/-i���_o���<]���J�r�F��Ys}����R�E����s9�EΌā�g��$zI�A�z�3f,[������w@{Ԅ,��2�+U��^���w5�.w%w�����(����s���>��w޶(ϣ��|�5ݟv��2f]с-�o���ĺ�)���Z��+��Fh��K�;^��:=�X<�fH�X�Ͻ~ȫuAա2ذhI�׽>ݪ��{�҂�۱��#��pXȎh\�?cb}�R<[�3�����x��y/�~��������t仵���}IZ�ϖ[@��J��A�>mg�d?W����k�����ͪ��<����fUT�G���T�5�<9����~"�
�A~����Y�!yzŏd<�y/a4�ޞU>����Q;��ٯ6�H�=�������]}CE�\��j��~���t���u��u^�����{�Uʺ����VMN�۩�`{�*ɮ�>��w�e񚳨�4�}��$���NϾ�9��_������W5��*R��N�S�D/��p՘�-��+�ԅ�JN�5�����$�u��,�뻿U��ζ<��;/�ϫhn*r8v��(ݶ��G�����]�Qζ�D���=cW�zw������ߟ�B[�"���0�s��:�6���9K�oVm�B����CG����םooeE�5�G��iV.�X�X�"C��m�=G*V�hMq��F���e��|��۠��*j�Q6���{�q'�,����������؟+��C�bc7��G	x�T�K-��ڐ����<;*�� ei��ύ��:؎��������z\{+��(��f"�D�^�?M\+T[�"�����2&�c�;�29��^�_�O;޸�ù]�՛��'�$���|"�=�Dd`S&�Tzhy[�9v�իv��}��TѷKrw��Y��S�E�N������|��ψج�W��/� ȅ>U��;�����g��ݫ�fJ+������|��"�w�z����\�#|�N��v��D������߂��x���g��G�w�}}{#>b��n
�q���!���";���9��	�U�^��-�Euܻ��]b�^�tL��hH󮑱��(��sW�6#~Ӎ���鞏�̝���Y~Y?�O�2F��>a&�e��MP􉨎�|Ɛ�޳�=�,si���lzcQ�J��{�{<0z�@{}q�.�T�`5P��GDk�;r�
��j}�Qu��Vp�y�Mz5gfs�3�'2�#�w�2=���{~y/�U!1"=���
�����,����X�ě8(�v.
#,�B�~�/,)^֋f�f�`]{�l��nui����X��{@���*�,���l�³��zR��?$�mu�av��gM4d��Z�d���D��#���k~=zn�d��O�;��5FV��v��p�;�I�h\�j��l����%J�ڇY7>�~�s����C�\˼~�L��*���R,��;,�����c����F\g�������{; �W�PϮg֫�*+��.l� �Z��Wx�o����ŠoԂ��/sҨ2���{�ز=���G���w��i1�~���uڪ���f~D~��TO��~�g���|�*KwZ������c����"�>�(e�Q�KV촆.�o���j������?A�a����g�b8_�L�#�ۊ����&�*��D��-㑾���ז���j+;.�f�
����F����~Z�ۀQ��{7g�8��VU���>�d����J�u�;b����>�U�f�۩���/��>�y3U�����]�_��~�V�ہ����1z��{�>���C!�ק�e�Y0w�S�7=^̴FjK��H�@f1�v�Z�s��ׅ{��-�l/T�27�R��+����	�oފ(,�*w{|o��zFHB�d��zf�W�\p������o֦���S�}�D^zEǦ�?���TJ��F��P��|��q��tt����v�g���+�U٤�Mo�EsN�`Tx�1�囙�(�g�z�GD+�`�Jju�*�k��w	�q�:��Q�u�_}�A^Á���ML����R�d���)�q]ܷg"\����G�GJ8�a�v�t���>�N6��ߏ_^��7�����K�FC��S{����׊v=����8g���DH��#)z͌��4<eZ�Ͻ[���x�f��y��=�����{*zs���������~V<L�� ����q?��~2��œ�o+���܇�aqۿ;9\A�+���B�.�c�	��l��3=�Y3��H�4�v}|���V��N���b���m���ϫ����/���#�d{}�cW���~�̟<��^���ɢ����f��=YT,D��g����r�A���Y��k�29�d4�vD/��_�.�1��ݷ���D��h�g��򮇢��ќ
�j���ʻ~;��h�۟��Nw +��7پ#ܻNT��I�a��W�G=qNɷ�%�U��~b�g!}E����٥�>Ȟ������J�Y<s�39��Ϣ=w�r��)��Iv���n��A��"7
���bbϳ/�@�s���懠]Ox_�f�W���a�?z��{.^Vd�=�7����LMG���R��M�Ȣ�&��x��"Pő��<��}�Zi>��j�U�7iɏ��n�8�RN���Kr����t&�-I��d��]w'�e�xYT�t�/���Q�uc�u�ж9݆I�ɝ7�|Ӳ��[]�`�ɆvH�!��q*�ܬ�� ���/���5�w���\�j ���Ddn&2���H:w&���M��� ���ޫu��[<v�N� ����:���S��4�`��X����x�5�>�h\j��R����0�`r��'T��5�,!l��/��ʔ�ͫkp�t0tvi`ޤ&,<��\�]�8Q�X�=���i���N�L���g<����[ëY.�J�%@�o[��R����'��eX5�,�巗E�1'��5��2�)�h*0䊳Q�t
���׽?sKc.�y6���{���QY<]���J�9�Ί��z*�͗f���n���_l05��i��_o��2:u�HQ�K�Y>�Cw��ɐN�9�>��Fy�_ꔨI'�e���e���q9�^��Y7F��)�u�<G��:��b��m���W�Kڢ����~Qpj=��wy[%�;��Z\eya�4y�ޏ��|j�!-U�l�s7�r��B�p��Rl���ط+6��=3�u�_n))�*$�'��`�x>�{�@M���;P�:�_+49���;���KcTL��񽌣nњ�;�u�O.�C�M$\�\���l+X�o4�IC�a�M� )���^Fµt�jV�h�%�������Sw�����v &Kܹ.	��0/g#P#/5և�Pw��+fm:��w1��R[�+�I3��,ah���v [�j�S�_t�M���-��N��fRk@ꎑ��_��v�܃�r7�JՒ)�
�!�^%�y;Y�;/l�����o'W;�1���z�없=f�'/L=��r���)1b�lU'�*׼�qͶ7�� �;��͹�Y��ް�+,�J^t��9�S��cyW���C4���-);�a{�(g��M���K�_)������
+a6Z�7E�YJ?B2�r܉��>������g*9�@i�W����)[��Lq�_N�b��=V�s��`�{��\��	���5�ȏ��G,�{ޞ��������_MY]�*c��w�����=Vd��1.��g]B�K;�jv8�!q
Pn�a�"����>�4���3�� ���A�
7��d����>�QO������M ��m�f�<)f,�/^֞���n$; ��]�Y��Z�c8�G2�f�����`�+��_4&ǮPj��ɀ7�0: �_��t[���Z��ko{��=�ނ,V�"ι�.mgݗ�վ��4W>J�n�bTx��6��!*ࢫـoVe�4��uN˵u1���t͖�a9(ǥ$��B���ڻ/Y�Pe��9���g]r�ǒ���e,)�K�r����[h	��
�l���n�yr*��S�͖�e�,�(�.'J�Pì���,Rwnn[	΅PJ&G@ڨk4+%�*��L�B�w\�P$���+T��Q�pҕ��'.V"fHTi���kR�R�%K�p�'M0��N���P�z�TjAU�5#�]�t����2�2Qb���F\�D��U$�EVQp�2��]��PJV:8�E��EJ��E����Z,���f*�$ή�q�ꔨ�҂);��Z���.�r/2�Խ)Gq7r/aJ��%QfXj9���Jċ��2:���Vhn����`�,<��(,���V�p��e��yȮY' �)M�̐��j^��ZY�:98J\��¤%=��L�Us�sfe"�̩��ՑAYej'U��(T|
P� jqI�d��
�5;]�jt�]�``�����#^`�ᴣ���+�u^o�v�aD,�
Q�%3��DR��>�Q>V?|)\��2�|r��؃^�y���3���x��#�b=�#��fn��u��&5����^��;S����U?"O�^t*���]߮��U ~���{z�9��_����u{N�ڜz��%Wgk5kѝ"�{�$xZt$�b|�����ӫ2�n�o��g���#މ`EN����Q����>�R�g���X�<��)����jB^��5M��r�ʥ���q�6������]�����Yӱ�u����<F��l���]*�G��C�e�R>��E/5�tN{f���`���Ih�{��~W�3������2@��z��}����"e �ϫH5{~�V}�x�<<'�[���t��9��5�Q�?cc`z���}��;ٛ��1Z�;�@y��^-4��|*��P��J�7���v���.Bk=c>~� <'�ӾR$��&�)����v��-���j�USp����U
��M�*�.r7��ҭ�_�<���e�n���u���:{g����������K ���g"k�"��=�;د��ߤ���9�5���bPJѾ�7ڪ]�|'D0�� �n�#7]�;U5�j���!O�wQ��Y�r�&�ܦ�@c�wM��s	����o�l���5�
��$��2��Y:�լm���r)����k��K������ްgh!���u\�.1��:��ֺn��w�]�}��}��f���OK����p�+����%�X�F2f�-�c�Y�S˕�s�{nJ�dz�ς߼o&�J�i�����Tw�tf������ܥ�͖�=��rC�9S����Nû�U��ζ<��맠����d'��|2�sS�g��B�Wh�����p��ȍ�q:����/��\��~y	f���OpPн�k7	�)q����`�7A�ӛTea��ύ��:ߺ�Һ}^�a;~�|B�©�{��ţ�Fz;A;�B/N�p����)�Ȣ�������~������8T�}�G���"}���z��\{.=������ ���np�ڿU���UZ��V@��zLyQY��o�8w&��ew�����g>��s�6+*�7@�� بQ#nQT���^��^d�j<��R!3w���\_���p�^�0w�s,��+��r�F���{Uǳ���s��\��g2��Ps'��2�l�3��Ee{ؐ������r#}��fs�Jc���7�k��bW][b�`�%�wܰ]/E�T�����S�X)V9�\D���}�z��KE���&�0���-uf^d�]W�;�"I���̖ɦ_�	���Ѿ6ڬ���y�����]��[7;sE�H^I#���;w�3wV�]n����',�7�>	�C�[�n[��ӮG㚸8����q�];ўt31��c�����q��c7�5SB�ؚ����6��r����,�5�s>dz�<�,Xs�t�O{f=ļ��k�~ut��������4׵�f\[�m{���w1�)}�z�I/z�4��=���ϣ�Y�9��{����#f��.� �=!�eĎ&+ơu�:��� o3c�<�0ox�t�'��[��ީ�k����
�N�۩0=���q�~�y���V���%<!�W�=���C�����3�~Ca�\ϭW�TWn\�!=�㷻�\�I�>[�� ���b�mzVD�t�Vߧ�]2�i��q���G��Q�����v�0+�>V5-��S�O��xTN�EC%���+~�Q%�W��T�o�^[���+=2����Zr���G�_}��o8F�*�`n��FW�<B����#`[��20�ߪl���Mq�>�ؤK���G��疤��h�JK���q�JC<�s���1M={;�B*�	J������#��ެQ8��9[��8e0��E���+a�`������UV�%�L���։~mv6Q�����p�IY���c�R���ա=r�x��Y@���zS �k2��V���q�a�X��`=D�Ev�����+�*vhY;�������\�{�̘{���9���lC��|�=���a�{�n^��< a��'��>�T�δ��V<(�n,�V<��1���!���;�>�;��~w�;YfP�bV"��5��n����%~��@�P�u�VF�s�3�^~���-�l/T�27�R��}�yz+>���t�-r�N;�Ռ{$d�P&Z�Nf��I(�w���SY�b�O�lǾ�ZU	�5�����շ�c�'S��o��;=v�;�2��5A�BrW��#d�_���}}��h�k�������~���p4��⭊,����*)z̓m>�p7|3Gn�H�Z�Cw�\+�|r�� �{�z�؟�?�K���e����'ߊ��j�x�叫�Ϲ#n<���c��������l߬bn�#�>�L�y�L���$nE�y���a�i�`2c�l�3};C�m��22�d{}�c>}^�a��3ޮ��;nQej�V.U���;j���"�e)��l�����;�N�^���~'�L����g���.���ݎ�L����sF��q��k�`�/-�Qї��'���nTw���Z:��NtW��2�}���"b�ދ���Y����?��>]�榺��H�64�����o�Xk�3B+y�׺|�ޞv���O�}'-k��_����m	�{L�:�D��C�l��O�_|S�r��&���xǮ,�ߍ3����V������gc}�Z�~Us\��b���}��ݐ*�&��X��p�+�S�@�#�0�@�8̅������,��;�c��\�~����:}�۩R��߅CѬ��~�I]ѾvR��^ۻ#��O��p�L�Ư/mN�<��P��\>ʺx��3q���SQ�J��EWvW�6R�{���f�S��v�)D�4׮p���N���{r=�ߟ:��b�~��^;��b�nO׋>O�r�k� `|���t3\D}	�5-1�z�Y�W�o�|�e⬉�[���le���𛋆���S�i.i���as�iA�A�Y�WuLx�&��|!h�:rǆ�Ox�&�����s�[��T���!��C�Bg��9���U;��E�~�H�3t��w��G4z7�N)���d��_�G�:9Do�'E��\,��������zc�]61m�c�[��l�!r�m��D-sQ�{��F|=�t=�0y��i2�~dd��\���h?�yL�Ld�o�"��J5�
�Nsܮ�g���n�#���W+j�t����U���؅���L�qW{L���z��u8�{4�~_25V9�uI�k˚�<��_�"�m�1|�&�*�M&ҵ\�a�nR��T�e��ԣw�;�,�����;������_S6g �y�j9�������Q�xlm��{3wr��=_M��{���p�dR���,Z2��j��R���.}	������U�)��������ֺ{�w6�d�5U>A�R{$�MҮ���~"��dg���i��;��w�Md��{�%౑�W�O������jϦ��:�9����.D�
���=H	�u;��t��^�e�>�˺�~�MW�sq�n�\u0=�k+��6+��G�V�Xx�~��<?�G�y_����I�=����N��k>��9�Dg��n �n�r:���*E�D�j�t>*�9n�����q���q�4A�O� �,����:��ζ<��#�:}Vv=�"�k}��^���^4#E|��C��YEL�A��ԗ3�V������߇�߽��#"����s��s����#���|oX�j�r�p슧;q5FV�`3�w>u�uW�dp��FoN�.o=V�Nd�_+'�ܟe���H���ŐN��"�ӷ\200<�9͑D9ώ]��l�>��?�S�;�|�s���7��y�d5��-�9��Δ>C�m"E9-^�$q���r
X<��]�\�������U5)iX��ER3f�����:qN������4=��|3��m�wX�7�d��:��Mն1*���O��Z�.�g2s��]Ѝ��)>�܉ȍ�z���_�����_Q������~)[��˘���]�����6��<l�fTQ��nL=C�Ν�E{ö;�2�C�9���br�� ,+o��7_��{�����ED�>�̫�ǟ]�x{�g�E�7�᰽S�G�S/��+��ܽ�m�x��^Nz��W�H��^ꙟ*��f[�H߈���o$����++�Ć�u�����������f�^ʘ����v�G	�m[p��!j���bj)�20�~{�b��5jP~��Q}�>ӝг<j��u��{��织�*�=�d�]�T�Ψ5X.���bD�*�ߖ;^��O��E}˦��v�\��fo�w�N)�����`=���ӷu3p��nj�{"h��z�/���O�t�r�jmu^�2��*}>�^U�0�u��l�?eԋ�T�7*YS��V���M���+������좁�7�/ݞ�������e�?g�H���ɸ>۩���N�55��YG�< �D��ძeań�c�x��x����S�bϮg֫|v��z�������bŹ��;���Iq3m�&fRB�c��91]+��Uٵ�hZ���o3����oF�l��Ie�+^���n��������J��{��n�4�u�:}|�ڒ�f�^0W
�u���-k��X�]��c�����3�x�{]]��ڎuΟldǽ�I�}����Sf,U�X�������{��Ֆ�o~�d{]���J�'��d���l
�\������$7��Wz?^�?1Z1�Ȫ��Vϓw���	��~����?@���{�[�Gl���r6=�����$�7�u�!v
��5���+;�/�
uy�[]�v����>�"����/
�o���~�;-I#a�ӕ\;�,BQ\�\	Q���z�V|g����{�x�g�Ϯ���	��Oޣ��O����yVY��۩�C���b���^�������p)\9W�eT���&G��6;�>����*�����WS|���c���P��g�w�0���3Q>W �=;�9u�^�\���lT�2Et=9�N�	z���uط=$o���<���P&|�9��K°�l9f�=~�7ݾ��-�u����F���K�G3�h	��7���!��(0�fR���݈yķ�W+*��ڦ�C�?=9�}�.Rܽ�N�8������9��8��?Y!5��ş/�+�l����`57��1�c��&��5
у�BE�T�c�F�#�Hk��z��E�ʴD�%� ��G�|9G"5�6�<����P�u�A1�D1,���˘�����[���{G4��ƹ�.}G��s�j��ds��`�4��w�f�Pbʱ�VV��+�Z܌���I�7�����$#��p^}�mI������޴��%�|Հ�=)>^'��K��Զ��k��a>��J���5�j�,�=Y�?�y�����Xȇ�Z���}~����ٓ��;�Sv��k؉1[��/�B�0��@U�u�}7��k���J�_�#�]�c�^ǽ�N�[0���ݯj8�Q��ޙ���2n��U
�ӓ���xr�t�Y�&�FAy�i��i۾�Տ���$�݅�U5ެ����Z2#��;P�ut�W~�ӿ,v�6n��	Ι�:/���A=��wѧ3�ο_��>��ߵ0����0���f}��2|Uw��t1�y���P��p�C�թ���3q�垝�߰�\�k��y�I#Nћ�m��*`w)�۴�g�
��mM/j9��ފ�=��n�z��c��fn5y{ju�?z�ǲ㙥�FJ�[f\}�z|6K�����õ�t�֍���IhTqV��y�3��K��S*��큟I�ח���uz.%߯If�����}w��{�@`k�N�?d%�&�d�.%���]i���G��@<�'���ј��t�ꙧ�0�E��Uov��j��b�K�K�7�C�}SR.���&�1�d\{B�.'��ӡ=sхh�--�yw4�{���+��MU
=]\~(+Q��X��������FNE���+��\�o(�WD[9�i����{⩰���<��\BE�p9�s�3�i�,�1��P�"ZnN�5Z���q���fvyM��G��>�[�����G��������C�!�ĥ꩟\�&OC5N6�q���O�->õ�r�}o�f�)�gN��_�\}s��H�a۸y�S1>Y~�h�e܊�۞�����Lφ��uMwC��Y�{�T����~�$��N��ۚte�ڛ)ѷ��x�׬*�;�$	��# �h{��r
9�pS���դ{þ��1Y�"&9;�)�����?S��S� $8]~c�5O������2T����\Mg�\V���N۳ݾ�J�\{�|x1��>����{�rI�N1C	6�,��N���F�E�l��P�ڴE�Ƽ���4avvgz����y�����'��fH��!�چr&��.:�:g�sN�{+ו=^��Z��yp�4�}���a�f\��\��~�MW�s|��E������3>�ށ!�[�.j}��{	K�Do��w�RC˒�I�׷�?'w�5�\�Z_�W�~#-T��-:�j�Q���/�٦^{[��Ar�c��'-u�%�IJYy�0�QJz*�H��?d)�[	���\f�Sq�2�����dc��!�;��ꎀ�z�#��j�~�w.�kx��Y���ia�&��kS�n%�t`�|1�齓�n5�MG�����{z�݋8�^�F��	�6��sw�<� ��<B$;}��N�I��햪����}{��/�:]2��e���r�NZ�sw�U�eVuغȕ���.(���nIχ ���z*�	>�|f��Z:q8/���i��3_n\�'X���mؼv/��ܚ�)*�����5}�[��l�(L{j%�¯e�f���g�ð�j	_�~[��C̙to`�<����Y��z_+츽�;^��˦n�qYhm��ː���������n�AS �[�9
t�^Dy5�W^�y8�p�܆��T��"���b���d?A���3��qpd�mǲZ��--����٬�C;�soe���xTA��d���.�{Ks���
���2@��Z���s2Q�5
�W�.�[P1���G �a�-v�'2���������b�y�DJ����Ҡ7;:\͙�( Ҽ�i�*>�uq�ޣ��򡳛۲�����O&� "�%�5ۙ,�2���v������"�Yi�٩��j�D켈i�m��M��(���q�������
Km����>�r�zT}��iG�F�r`���S=�^ÁV�Z�*�#��j#�ur@L�[4Lݬ���Z����)ꜱ�/�<��a�W*�r݀�@�Б˝q�G.*�.h\��z�h{��z�xt�OB�n�����}�ǁ�"�9�
u���� _@'�fs���u��A�;ܐ��W.C<�Fc�率�z;ۄ� 3̛`��h���ە��`�]�Gu���OQ�U�bS�C��j��x��^^���������KLa9�K����I�C3+�׭�e�Rwm�;��-���W��s�ٶ�R�,Uo,�qY��æ�.�mt�^����Gk��
�k����r��}r��<��A-�v�U��V�[J��x�!��G	�`��y�Xd�S�8D����I2~�ѝ*BĖ�X�X\{���5�ʕ����Wk:]Z���}Y-�{�،�_�bͺ����9��O�&\����Z�<]P��6�'Bh2���M~}�C��6�=��YD��ϓ���_ʒYڳ7�(��+zǼ������kL��еӋ��'n=fX�y���O�~�T�ղ:�*�17P��חNn�jׯ���$zz	�,�'zU5b��i�k��.N�A��v���M�J�Oޯ���wu�x��K�5�!h�k���m���`��v�U��wj:�4�����.T�g;��w�n8��J
��s5`޴�uȅ�lV�V�1��<���a�L8�Y��N��<XG�I
�3T�.P���]3uۉ;�d�uNDG�z稳S����(�#%��r�	dE�t�YU
�]�]�r���rOpŕ��5��IDRdI�]n�Gu���LD�P��$Em0�*H�̢���L�u#+=�%�\�(����	��{��!E�S����A��kT0����pДI�u�ʪ/C���0���ajs���FNNQ�[�yD�wS�^e+]��$�O5�u""�Z9��2�w���2�tI�wBs1'/J���d�W�'H�����I�$��NC�������H�/U/w'R=w-iN̈�D�1�=GU
��&��+D��(+]���·�˹"�y�E^VQ��yh%M:�J5"�:�����x{���֏{�x�ſm�,�- c��gZC�)u��P�8����dE��՘�MR��ڼѵ*t	�!#ۂ�M�S�W�_�-����f2����b`Y����~�����s����ˊ�NkK�x���G���}>�5�7!ґå`����{�F�����j��L�;���.�'��*�t{�����z�g�RmI0���1���g��Z�̗��w�:.�����;C�g�w�Jo'Hk��͢kr���=m��o���]����B/�;u�00<�9ۑD9�9w�	z}Q�kxU���e�X����TVwzH=&�W�z�"uǩΧ�����Z��V��&N!�M���U�'r��~�ˣcr��}�eڳ[v⽐��L=C�Ν��E{÷�s,�[�p:J��p���.���z�^*��}��Q3����-�=��ȯ���a�����O���̲3|�Os ��3�^)'��M�;���y�zF �=S2}WC�A��)����(S��{ؐ߃��DmW�d�rs�}l��ĕ�enc�7ѩ���U�Uê��(+�X����#"��繊(dsV�]n����>n��n�x�8��f�@Z�xw���C��z�¥��.���6&�/*�Ŏׁ>�i���k���:A؉c���bH�zS==~F��(v^Dn胒`4�H�}��T咘�3(�����,uL��|(mfj��[q�/��Vd
���˽Bf�Ԙ5�1Ewk�g�v���+���-�'N��wz�0a��]�s�7�ڧk����`��N��Q=݄�G���{܎T���Y�s��X<'�z�bk�n�f�0�4tG@1{<@���t{13�N���6;������|���+�������;�q��uR=
���!���A3���<Q�����q����K����dd��N��;��S.߭��~�����T#�7�5T�U�\��To��,~��mXW ?����6SC�rU�0�vCO�d&}s>�]��ê��K�q�-`�.���e��ZW�����ׇJ�zRw?����i��q�ر=�Ɏq��t�N{R�QAz<�"�}������
|6��~�CO�w���	���Ű37�x;��,�9���ǧc�����c��䓿�"��m��A�݂���y9w��+���;�i���C��̧�^�?j�/
�x�������ז���h��ۮ��回�,@��յ;�~W��+�N��<9�0�e���fL=��`��Oޣ����l{1O��e�w=�������/|��r{��+�8�Gq�}9*>����q�sy������ީ�}��yR�Bw�ȷ�V,3��\�Fy�[H\*�M�z�귱���Q[�j���{��f�ڡ��{W��1��J�Ua7B�D�T1L^ED�dtv��w�����K�̍�Ψ�y�|�{�����hf[N:��&x�}S��oJ��ˠ��yBXy��u9�y��yI�N�Y��3ެ�>ȑ�z�T� @s1�P�A�lzv˯���&���#x��(�^g���w��=�z�6��X9�Y�
�D���3�!��^d6�g,�2}�M���K�gƻ7}s~��b��{�l����{ vG�؇�9A�2�X��١,W�BJ�E�{�7���>,�Z��k|�Y�?b�;�<s�=����F���/�+��e�w��sR/�D>]��ߏ%�� c�����sQ�G5�&s���Ώz�؟V�#ζe۸��>��������M������O?Z2܏��YMz�C�>b��6��2�jG�'���r%Q��:��/ù���ٟF�|����p�(�Nv+x�T��d�X��~��e��^r7�����;�X{���=���X�܍̟o�2o�=�B�U*�����O�e��A���g����}�����_S��`����^�k1�E�º�����pz���U�JW~��cCq�w\ܫ{�<�+y �S��ٝ>����cY���W�G#�f��{n�gv
��q/ޫ�n&���T����I�(���q��F��KJ�m��]��1�dĐ��ۼಫr�[��sx�q�����ʎ� �Tr�X�e�U�3;��;���D�`�ȭ�cZ�xj��[��¥�-��}���|�q9t�h�pܶ�3�s��k��������g�/�dv�,s3q�Y�u^�b�?Z�~us��v���n�W��(�K�V2ZZ��g�H������;0�^�c��foW����~�]F��B�+�|.�&���D�w��d���y����s�U�(�#~���)���5�}>� �^�:zս�b ���/�F��x�3�z�W���'�I��%��	h���]GwLds��~�g&/ɒ֯G���#:����>�<�G tR�:��3Q#�9Ö���{G�O}�y�
�ۻeJ���}W7����'��s�����w�-�W�?��#ͧ�l0��#������}�+�ڽ4����T�U"����(�{LԆ�{&���x�)�p���q�N��Fs�~H�LNd�3>�R�|棐\��++�Z�C�����}��+�f^	�{Pd��ޅ]u�/��ޤ�P��w�H��t˺1�o`��b࡟sB��l1��=ᮃ�㎈���.��vڑfoՌU���LM�Bk�~�7�,����?�y�g��ښ��5��g����f�v�\��,��	�Qk�x��xQ�2�h����Ƌ�𜯱`����"=�ٻ(P9�ӵ��E:&�P�a�2��	R�fh���:����k:�)|3+�lE���ެ3���h���Y�2��<��rQ���#܌�k������??b�>�n�wM�9$��q��~�ا�\��s���k=�zkM�#Kҗn�=U'��2�g���,{��=�Y2�װP0��C9�״G���T�e��ǻ�������>���{�7�9�t����s���.��zk����yU#~�`{v3޸+j�y�ݎd�w�W��xS���+�y%~��{;=;	���}s�k~�͚#�*{���я;.F{������u+�
�q#g�`��DU�y�]2�O�b�K��s�O�ε0����5�sx�f�[rO̧溞~�Q8|��:�|��TT��]/ ��S���~��&%�z6��(���h���n^` zW}�pI��{j�J�����^�Z:V���~c��>��~����f�h�����Dh�R1�߇�o�����x�	�z�^���Y�;H��Y�yD�W�t�3X��I�+��lԐ�z�^�_�N}�=ny���_�z�D0�[�np4G��ƚ���+*�߯���ZWg�X�
7��.���n�Sȇ�ra��t�z+��޹�r!������q�å��m��xOǱ�\�o!U�s� 1C*���+��iCmcJ��g���/y-3����bZ��]9RC�~�n��b��ά
^*�T��O�o�ڔ3h��б΂OXOVo�i�*��҆��W|�i��r$�(�oe"�k�%6-<Ivm�h7����ٵՈ��
, |*M|�L��l6n�����o=�xO�s�\�"��7�+���ojU�/ܢׄ�u۟D�BfZ����2��f�yo�"��i����F�[=y繧��cНO��`��U�CrNq�M�_@�wF98.��r�-���j���4�������\靖^>�m�=]�d?{ vz�¦�uA��u�T�\�Zn�9���'K1͚]�yh�!J�w�T�Mg����ǃ�z���U(ey��/�%]��:x~S?d����s��:�.؀�m�DnW��*�>g�*}9�,˜^w�=�O��=�y5�u ^z��/!�:�"0�Ӟ�7�*_���3}�~�0o~���/ݞ���w�z�]�~�L��e���K��J9٣��c�[�wmԋ�W�W#e���ed����%^#gd=Oوu}Ύ]�q���Im�]��d�V�����r��!�V�r<�+"z�^DU�z{~Ym F�O�ElҥxeH��������}ul�=�]���b^��9�p��>-X|���j߄���g��?��P8��陵���Љw>�'��̡>��ȵ��~#�ﶡ�R��酃�kjat��;������E���ŧ��"�x�^��4�B�=��6u��oR����Z-r9��;���׉��}��	}nx�������zG�E�ɼ�I8w(�@��s=�Y�߳�7�e�_�$�7�h�}P��શuA'���>�=���޲ׁ>��������/�7��§a��zF�{/��)�������89�+e��GZs&��g����2�1�{ �̱�̷�{2a�{�~�ez|\{1O��9�0��%j�������ϵ�Ԭ��  O��J��������i��o2��p�	�{^=�oWk�*�uk�=r�pߤ�e�Q6�U� �s5>W[cӿ3�^�^Mlس6!�*>�ޤ�D��U�c�s���ީ`�F�d3"�g�!�g���jU/
2_ZJ��F�Tf����iY��8mM���b��O����7����!��/�e+��ݐ�V*��.�~|@\��	�Ω�]�ec>�*v��g�o����7��2=~���(0�KõM��#.����9y#�e寮W��f�A����5�&q?<s�޴�}[,�/�-0�yYY^4���7z������P��R�ρ�5�~��)�oa,��|��ϛY����H�w�n��기�N���f��pns9f���\���cgxeԯ"{}pg���~��\����*Sg��t}�`5y�=���L����`�}�,>���+;��=�v���6{�V�����ë'md�����{���������s�;Us|�|�N�TR��8�t����/�R�A~ۏnt�²�E�^N�gu{ܖ��鼝�X�G,�z�O��d�ڡ*�N�'�ղ���|q����4�ݬ,{���Wth��?(Y����f!�>����U5�׶.8=�>����N�5�=}.���_Zw�\�o<>��T��A6����ΟN�~[���~W�G#�f��^ۭ����Y����e��	nyw�/�Ms���q�ՙ��3+��=:����~���y�I#~;FU�����SC}��Q�ڐ]��D���j���~����j�����~��e�3Su���'�(�$i��b��U��'��M魡�? �@x�p��,'�(5�y=~U�w�TU��sNq����yc��nCaz��w�̨�[C�� ��~�tz�c��[<׋0��c_�1s�!��D���)>�܌�\�>����y2,������BA��Nf'�9F|_�M�v��F�\G;#�v�y�ɼ/��3���s�޹`�?<���r�� '\[�J謱c�&yuGFp&��U�G��55.#��f��Nv�{��5
͠�]b�
�#t�����O��^1R�
��kX����]�Swu�e��"CI���j!3{�:���1����Ѽ�r�yLw[4t2����iׯ*եE���8�+$7�LS���G�o�f%�UO�U5�f�+��gMO�)�gJ�ט=���Z��Өk��C�ڜ���,^�/�������Jfgޢ�����G ��dVDW��N�����fH�Ƿ�+��ݔ6Ύ7���4xO{��Q���;���u�]юK`�O����_sB��~�����	���Ϻ��O�E�����'�)��� ߉!w�А�Jo~Ym'�B��n�|�ws�5.�a�4a������N+�W�տ������6�b�&ߥ�)�̹g��dl��哓��{ޕ�Vx�h�/�S�y]؅��=�{���{3_�
����gن�S�	$7���g�������8��{�7�9�y�.v�e�>�˺�{����a��������閧{7O��� 7�D�C��լ�+�y%~������;�!��������ff\�u���f�[�3�����[��W��j�l���"�s�l�@�ʟ�A�Y�uU�uN9��-��ծv|wj���պ�6쯽}0���So�T�b�,�c��~�3�1~*��|fc�ψ�w���^G�sYʯ�ְ����lu�S�d���%,㜬��E#���E�:�3oN�X����ήQV���:�-7/��v%���UPT���PX����s��v�pv�,Y��z���<��7����<��m�x��x��Ϊ8�g�v�1��~y	]W;�c�KUw�p��/a-+c���.�jn���}>]���g}$׍R��p��Bt�=!�/�ڸ�u�FvUhQ���9^��T�ʼ�y�hyu��#����.Շn�����S��H��q�s��~�[����Ȳ#�ۤ/"Q��c�ʮ�ty�-]� o�F1p)Y���~�[v�Cǹ0�!{:w����\�/���\�t�z���0���g�wӔr@��P�j���9nVB�^�{<r/"��pߡz�Ύ�V��j�]]V����[��N�}�؞�]�y�Z����w�E6�3y%�~Y6}�!Ư9��}�oZ�����\f���ɯ����p�ܓ�L���bCtdo�S�s����)^�s��;R���{��︛���{>�m�<��[��X�o�>��������8E�U�~��g^:�;厮|��@��z}��'!5��;����`?TdO;wS7�ɨ��)TT ^\�Wn�0w��ۚx"덛a.�%\>j�\�n��W�������/�c6��l���6m��l�A��o�l��1�cm��������6m���l��1�cm�lc`���q��o���h1�cm��6m���1�������c6��l��c`����o�c`����(+$�k&�{�r�0
 ��d��I/o��@Zҁ��J6����Ym�AUZ�*U-a�	K`b
*�4-[Z@��T6ԭ��!B���"�"P�(B�h��m������і��;+늎m�m��/v�\�Xcu��م��f��ر��R��QV��,d���^��;qŵ5��IL�l]�䵶Fͣ0z�_g����KKeZV̶���՘�ͥi	JF��'��5�R(�U���k���Y��Z��J�������U���۹Z����F�5�l������Kfٚ��=�  ���򜭶cw�=��e����cw����.�g���m���m�yw�Cі�p���Of(�<s{z:�T����[6���ާ=UB��j�vն�Ƕ�m�6��m6���Z�)�|  �{�٩ֻ��ï]�5���ᣯF�rz�=����\Q���m����@Q��E�a� �  P�N��@  ���
���F� �w��Y�lVP�2��b�j�p  wq�Q@z5>���}�U�i%�']1Z�g88ֹu��\=V��3��z:���3��P�b���۴iU�6�q��H��y{կU]��f2٭��d�3j�� 7��L@���tu�CZ���0R�v����RP��e �-�L��L+���ޫM��F��.޶����ۏv�j�a�=�^����-M���Q%�k2kU� ���}�7I�;����n����l�w�{�T�m��S��{
s��4����r�u]��H�tz��t���=��w��{vk��v�p��mr�OzkҗiQ{ޞ���4l����v��m��Y   �<��N�t�o���*V�im���מ���f�;��Wm���K]O]w���Ѧq��ۺZ����2��T��F�;��+5���e,����'yu�͜�go-6Tm��SH�E'�r�K>   ��Ф��k����֣զ��oxw�V��iW{f�׶©۷mz^h������o{a�N�S���]A�x{gYk�Nk׻=�A��uz��=�wnס�mh���[X�6&�M�B��    n>���}��5z���owrvʭs�]�ۺ�ܭ������(��N��s��GmZ*��חu���c��k�(%����^�b������nݮ�:Vu�;�����i�kf�m��d�n��U���    �>���r��{�t�ons��9��z�mJ���I��e�/{�׶��89�;��Csv�V�<�kO��U޺����]�Q�ox]���\��6z�zK�l�z�ը��Z��h�����j��π  w>�e�yء��ǽ=2:��gNݻn�%um��+ڳ;�nZ�oV�-z7,��z��S��q[�.��^��Kܧ{���[EmN��JP�l������f6v��{M&eR�  �)�IIJ�� ��fL����H  "��	R�`  "��1�U5 � i"Lʤ�0���~�������������q����x�����O�a=4�����W�}_U}��?���ﾨL��BC�@�$��$ I?�	!H��BC����O��u�_��ݫ'����ݽk Y�+�VR�4�x\��"�,��miѝ�Ʋ���4���o"m -Z�(;�]�H�z`ƅ"w��i7�Ũ۫�p^4��#tI�B��B9fԼ%Vb�s .�7�[���z�+�%Y�P��B�8#Z�L��,M�jy������1VMU�J9%��ߞ�l䛎�7)�V�׫6�RfʷFi!����x>�u)(�7Pk���Vf�����ͤ�:��l�Z��p�	ތML�㎅nT�����%��ʶ���*��k]�2�و����ܧ��vE���i9V�^壠��2%�"6\e:��,cB۲`ϳfH����JJ��nM�v��!�l�Mm��[��  �gFSi�X��6�ը�'n\3e�2\V@�/!8y{��Qpv'���@��K��\� ��r���ma-j�aC�`r��m��)��:�`B��/fbʚ�wjlm�m͠������a���l%ǨL��(n�f�����G+Uȣߌ����`Ǒ�/�����]B(˧���.�Y��E�%�([Ul,wly5ŗ����0c4A��@�����S0�U��&e�M[Wl]Ų��5���S+ "��I�����%Jq�l��5�@b�/F�e���.	G �&���0����=#�7S�A��Ĭ��O'�Tz������v.�醚�ڔ��ݍB�$�7�xɬ���3������=���'C�MъA��ţHu�2���%�hH�F��˷A4'z��Ű�:l�\`K�'��*��V��#K�cd�T�ĵ��?��{5�-M`CSwtIJ�T%e��>���2J<�X�Y��X��J4�ڒ$��o)�x�c+v�H3&��M�����|��e��t�� �����wEc����,���-q��ń�ua64�I`@�:I�CQ�HֲM�o0rXa��f����F�����Uyb���V�Q		��8,�n��e�l�����#N�UKr0`+r*�cy�^f��m�r�6r1��*�k	�EP��ڒ�D%�a��WBb����A��YN���掘4Z{��d�ڵ��U��f�x7bC$0@R�n;���z�����wt�n�����"�gM<Ż
&����Z��������ݔV�>��G�h�IJȅ�2f����BmMX��u�0�G%�g[��N��U*V�,�X*`�7�^5�AfZ�^\H_[!���ʶ��z�U(�h�4�
"�l��K���I9-�D�&�;��ܨ�[P�Zo&�){��#aas5x�EO}�P��c��29�Ű36B~h�!8Q��S.X��|Z�{�N`��M�����$��񍑺�r��k���ӎ��o+�4<��p��]���2� �����j�ݰ�Ժsfܤ�㾘yYoe�"�e=� Zpq��_l4�fe�SSd�յd�&柋�t&2��F�:�l&TCU�Bn�6�̉��cW)ѭg^��m"�d;�$Ac9�H�=m�F:˩���-�HrH��Qc�C"�
�"�=i7���T���e��d�h��]Y�f^�nT��=u@Ճ�veT\x�J�wR�(���VMb�LK��B�mD�ֵ��
;��fPZ�iѩ�lʶ#��[�<��7>���N����tʥ���P��e�/r�!tM�Uy�J����j�-:UNQ�wD���
���/o�	{�ҔI�n�T�Y�IU��-+�V���rg�0\ܱ��*�[�����!�#�3c]���3���N�,Xl6��t3N\Z�U ��	$�����Crd���]��u4`ƨRw����ث�ُsN d��m��d�6��,��*�p�HZ��:�1���ռ�a�㓢�^˹�]��ۊ��{��w/l20DV�
�7�i�J�vj۷V�c� ��6ehW>B#AU��h:5'j�L�n��@eb��ۢܔe��P��U���9�.m: �-@��=���k#�ne�uƴ�]d�G ���u���ij����6��{��ޓF�n
R�񹔨ѷy���bD��VX��ñ�ũdѦ�)yq U�pm�E1^����W�@���G.��^����[4�٥��GXKZ1m(^��!ѶudiZ���,"ma
蓸n(dj�b�;��Y�
m�Ӂ����X,eKz�&�d�8�H�x
�b�J�j������uً�:Jv�:�"!zF�u�N��e�2�3]���;`J&��#J��-Շ��B�<���L�c��s; qL�= gE䭈��u��uf��!X�,`��2
�4(�p,a]1�t+�#F�v*T�v7�ⶣYB�]�u��2���
� 9<ôi��5�5�4"E�/����<t�d!�-� [ش��B�-#U-��w&1oқv����7Q�r�5T�OmG����ҟM�\KS�B�I�L�%N����(�yr�h�
�"�Ϝ��@���հ!�Z0f˫��WN1-`n</.��gct�ZѺ�?(�w��,�0�,lQE �R��ݔ��K�tS�T�N,�-�4a�4�b�m*�1њ�6�z�1k+.�f����h���C�mM��"F���"f+D-�@U0a��kۺh�-Rt.�L��Xӎ�'�'�UG�n�-��+d£0@�`�a�N��L��;x�Ե�1H��s*$�Y �)89(;�%�V��Q8w[?;�t�F�e������:m���?9���WB��=�6GlK:f,:49��L*/hd����SM[.��q�T��Z�(a�8��h�D(B��ՒY�9�JQI�^�GE����՘iy�YQ��E�2�u��⣁1Vv��Z�Yu�jm�@���S7i�w��6�<R����dݘ�jm�Lѥl;[f�������ڛ�72L�WZ� �u�G�]�{7^�H�t�цejy�Q��e�$�T��nDƵer�-�h�q���k��O	�A��	װ�X�ڦ��CY3T:*ŹZ�ӡ�67JC�����G���Z�Al%�ՇL3/$ԁ� [{ohX�Zb^��N��t�,�ll-f-Q��*b�f]c�u���¯V8 �"���	�Z��E5��h����E���Yǘ]����l55d  uH[�yImB�����Ka�W�Ǌ���v�YaR��^Q5uaS��f�t�k�I�,͚��Cj�M��lX�hZe���$�s��96PҠj�̝��HEZ#Cz-�W��i[�aݚ���&\�]=h�kn��Nc��T�F
e�32V�a}�Lo�7�[t�Ķ��h $m�##��ETtiޱ�iU�#�J�{m��Eyl���F�O�Nfc>ZqØɞO�ccg�6$�D�B�4��x�@H���B�ݳ�BJ��S\���qЖ��¡��y��0�I�Ze�ѐ\'͛0�W�x��yj�l�����`
��܃��0$���u#�7VM�#�8���٢X��X[��N�]F��kg<��'r��p1d�f��⌒c��N[-QY�>��IGX�nn�D3N�wq�ne�K0��0�I�?BBY�d^���8��\�Fx4�^�j�!
` �D= 9YE�q��u,����f��Q)�f�5��<ab�-��ݬ��u�/�d",Y(ز�͋(ڒeYnD#,%�Z{`��9{�X�!]�$���q#+]��Ae@>�9jӗm��-x,�0�!�Y�H�;�iMf��S^+Cs�t����y�F)U���1M+�YN}q���c��X�T��6��n�t5GZ�1��(`g��6 y+4��LἼ:k�*f���c�$�� 0},����b��XZ%L`[QѬ�Q*����#Ndi졙��[�e�Y	�ӊ�X�"6�:�2^���L �/^��r��YxY�٭-��,Ņ���8;{�O�������[u����ш�eލ�T��ES"�G1(&RR�z�4�J$���a�xp�p���e蠪�V���N��38����g6f�g�ChG�]��2�^�Vf�jb[�ęzE�����b ��"� �v�2�˻��:�x�+Q�	={`���^�m�FUH�^����6e��S"��q�t(�m�o+4|�ۏr���bAl$�͕�@(^�)��ql�[p5&�u���$+UU��ITiIWR��魺MH�#j��Gt�6\�b�`V��`fD�Ʉ��X!;��a�1g،�n�����^�olēb���[�����W+`6bY�Q��re���]�IJ�jU��.;XA]�r�0uVr{��"�D¬"�[Q��Gdq��2�f�w�+RJ.k�"�F9�:t���j@�o�i�7Y&�b"��nXl��â�RM�{GTfl{1J�V,6�K��2����&:��<�[�):��0#���Ab,��t�;v��٬�x>_Ou�yn���o��0���VlM���]�P�)�B-a�Z��,�LQɃ�.äM��^"�1b˶Q h��yy����
�0��hgL�t�h"Ҭl�'�Cʏ6(�M^ؚ50��M�XY�Z��{���˰�.�dx��*�ɛ�dj��W��2i��.��y���Y�q�����6����YycD��)�̧�#�)[y����h1fB�m�y�D���[
��m/6���k�ʶ��z��`c�ncۦ�V5���f�!^�D���/�
�%;�B�d��1[��FռݷJn���Y��˶BI`m�OѪ'j�0�U�N�~��)��H��#Yj�ܒƦ*ܪ�L�OtX�`2)�����!����^��u�a
����h���ڀ�o�QA�Z�KTYu4�%�3^�<U���hͦve�z.���k@�	᳴Ԋ���F�����C2� �*��౰eY�j���7r<�e���^�Z,�6��Y�D"mfn3��
P�1:��1��of�[YSm�����b��F�c��3z����t�Tmu���r�M���q,�U�u �q	l:����4�Y�N!�u��C�]@�/�NZfֵ���a���-�/dL]��R�e-Ob1�񁈹=�Jz���-��EM{f�!;��J=/mK�0� �Y�Ral�j�_d;�T:���t�T��wM��4L�Ee�-�i�OTp0M݇{%_�b�ڢ�1U�*�v��bn�y�v㖔��Un��L�:�������A@l'�`p�3�,�x�M��h�F�A�h�0�4�d��o~��Z��k,}6�֤�a�d�n�"��j%]O��MnR�Cm\�v�"-kEJ�ꦮ���5j(�e�Rfō���KR�D�� �+Ǔ~���=$����th�)���L���z ˟7,�6/,ʙ?<�̻J�T�V�u�+��SH��h�޺���K)�O2X�Sv���Yоa�G,�Н��	�82�X���$�ǂf7��nC(�b�2�
�Ց���%�f^K5�	�[��Y�]��4�;�
�V��e���(#Q�X�N���Z�6[$��m��Z�q2��ZY���4`(��!��,պj�#�`�ˎ��m�yC+#�q��ff(@���@����A@]]�hң,���\Ia(	:ז�U�!�MR����H�,���uQ)�g5n����cFH�"7>��Y.�#	a�ы4�j�� ����UZ�q���[vK��Y)8q=�ɻocO3T�д��+��0�i��`WZ�?,�s��Y��L�3f!�S,+yW���X�(VH�C
�Ç(�Bl�&���Jw�%X�x.3IF�nXÔ�zp"����vnU����b1�Ksr[Cu,m��c]Z�IR�맚xnH�Z��Pn9���(��eZ�"�Z�U� V���m�F�8X�3abaIt��ܖ�� 1W�vB�J��1�/*���W-J��b�N�Ve�n�ʥ���<�xvMХO���Иf#x�W��c5�B��[����-��h]ee�wg�c[9�դi�(By2ኯ`��ek�n��6�V�5���z;.���E�"��:`|�^踄G.8�)��Lѱ�e\0^�ڂd�)�tP�4欵CHӠ,�>M�Xn��"�ƠP+��g+r^aM�n�B���#Q' ū]�i��wh��81cB��Ӓ�ī2�A��i�p2�r��HyF?��*��QIL��[��K�V��-dXP7#��ςr5kp؂�LR���T�T)�Ґ�ܭ�x�Z@�����y1_�b�4>Z%�!n���%��n� ��:�Yu5h��^K��Z�1�,l���f`ʺc-�Ѣ��!w1��)��	c^��{��$Kn�Z;�6�,҆࿭O�\G@՗hWQ�K.�c���Qӭ6-�m,z�6�S0��oeBEEG�U.enI�c��,(5K�"���CTh�n;�I+(�|��P���pm�x.R�,�� kM��B�Śa�i�5,�yO@�qV�2��t�e?����!�K�j����{�<������n���6���@���yt/C���Wlk����ف����[PYE�* ��FF���Gu|���9[p����@��je�?�^�9g�xU�r%(R�@�w.l�����<W���b:^�ӓ�GMh�Ɗ�]�����n�/P�VZ,��"T4Nft���u����7�e1��k��)�!T�4�����(L�y�v�s����K<�+`�\��{�#���u�%�0�������$���=�מ�| xۖ��Fo�5�u�s�.TN���yX/���kr�}0���I9���J0d�v��`O��w�	Ko������2���sn��o-���:�ɒ������mz�ףq�o�`�:�χ^/�Nɇ��ք���}kZ�ycy�Q��+3�da�ڴ�N�$%Lv��
i-�g�	Z��ҭ�^�=oT41�hmp?7����%Tf��-����;�_fp�2���.|TOn,�E���;	αGik���rBn�Ѻ50Z��	��%[/�\�gL�T�J�*ۛ
{c�+��L'Ȅ�Ϋ)�]���f�uoX׶R���ݬ�}B1��7�S��E����y���9Ve.�5\=��[��]��8�d[}�1�yN���C�r�i��r9��jw3��AD�Gi�����m	�IɻlS�^*��grgP�����E�yB1\1�+{(���0yz��ʣn{%�^��ہo�<7�B�vVNT�c�[n��9���ُ­�<���=�А7Yt��a�)$�-ĖD�muz�c��9�8QY:���[k�[���to�y��J��^�
�J��ȹ�R#.���w����Kw�;���:���ԏh��}\ĳw��<��l�?HS�+�y�"�AR�3'T�R����lWq�s
���y����t�+���E��]ю��]��OBcʺ�OG�jˊm��%v��B��+{R��%=۽����3����;EA����\mw��e��o����ƬtiQ%�*
��]9وe[����q�)P��6\�yx x^y-�s�9�G{�V�#���q<�:m�X0�#ckʘ�eZ<Y�������4h����5��/��m��c�L��Ov��]�62�};��5Z�̾�S��@oF�p��J�+�a�:����z��
����6�����<�S�^�V.`����tR�ʛ�V>��%�S����<=~�=�y+D������1���>��ӹtN����ѫY��,��3Fu��p=1be�1�b{�Ο.�rÛZ]��b�E���,�l�̬�ѭlĥ�{�Z���u�I�@7+8�J��h���50��ޢ3$m� ��f�QE�_�Y�t3h��ِu�5<᳝�����4rQ�M�wXaZ��j��Ǡ��SA����I�j�[�x�H���
���Fӭ� z݈o��2#�����斂��"�oP.Jl���ō��!6^T	���	��H�'wY�5��S����V�{��t��f��3�*����:/�M���Ĉj��+`��On�.�=��g'���zb�p�]-�;{]�wi�av�CQ���J��q�Z$>v-��؂�2u��ݱb���J���u�����p.sfNO1M����ͧ�����-��ിstN��sۨ��	�����^�aV]8����Za�ΰ�df��ٰ7D���V3����ZY�<, ��I����{<˜��X�j,�cn�>#�R:x\���rPƈ�"���C��3���4�mЧ����֚-A��s�<�J�-��ݼ]"�֮�b+(9Y7!���%ݵ���ޥ��*C=��ڠ�}b�q^A7j���=��xC/��]ö�ޜA��u�u�^ֈut�����z��N���v����ai�Ɉ����P�I]�N_A�k�[�14W�����$�{�
?�>	���0h+!�3wZ+������s����O,ؔ�ݼ�+\=���:�,��e8{�l�8�Z�B��Y�����gX�q��9v5�-mP
��P̈��^z�<5!/���j� t���6]�-�v��
����Z`�w�4{����j���H�<'=ŷf��rp7�fp�uҺGՖ  2�OR���qVD!<�Ʒ���z;�.�f��(�̥�L�)��ɖ�{�'�ں�U١���ǌ!����f���eĆ;i�a���p��|�p�/��ۗ�{�1
�gUПlnޤ�2�����cj�sf�pW�1CA�W��f`�ƹڎ��u4�<4�nr�N��%T�I5�>�b���N���֗��4�񽻂�NY��fnn;�6�[y�_��8�	�K��|:�k���{۴��+��<�:B����K�/o����u��#p{sp]��}��!1������yNiO�:�^�b��o�m/wx9'��T�à٣I�ݫ^�	9p�;v�����DYjo.�+���i��n���i����=d��͇�����ٟ"��k8��Y���A����"�m	�V����^�������W[�빞5�Y�����2N�`s��IV��_�W����������k󱣐��nX���Ǯf=6�93ut����v�+��h�w��5<I��qzAw}v�T�o:������ª�}*nM�J䅅����l탋k�\YI��*�x�$N.�Y2�1��۪3XN�$m}�߲��n���S�-M�x���}o�%p�`���s���]X�ziq@؆�(]�yV��a4p����ZF1k*�
�ki%i��I
S7���#�(]��Հ���*x�:�=&���jp��ΩhM�M��^�9m����R-"�w�rKyX�4b&R�-�j�Z
޸o��<J��A�c�	�izz�@���W0x���b���ڱ�oQ;��=�ѽ�"!�B���i<~~7�oَ�eV-	�H�4���pk��P��v�+<�+ldw���
htj
��:k�1�H��1󫭥q��ڦ�2�40�D�������v4sg7i��1� �	���R�X�z��Σ���x���%��E���cE�h��N�$>���l��Z�DQ��Κ	�FF����ϻ��d��yn�Wmw����m]n�C(�o,Z{�R\Ʉ�f_�,�t�ܺ��w+E���� N�I[�7�j�h� 	���]��K��i���wG8!8��n��C]����3>�.-����R�Cf�%�n�;-s]5���[�b�h1<�M�{�����;~U2w0��y�6kHu�J�9vf:���c�F��`�z����u*�(2��XAlpO��+և����Du�g
�W��sY���'P���s4�S[��̨̛�.�!~�+�t�ܽ�w15�U	�g�*V�/3<x����%N�%<Ŷfb����5Ŭ��gm�0a�ԾW�*��.;�S-#�H����IWB��z���k����X� |���-��Z˲Eg{Uʕ3!�MM}��M��-�s#ȟ��k�!W��l�7#��=��Y�~d�0��ڻ,6�T �;L�;o@FgSˑs΁���,�JK�_V� f�H�f�D�o��V����5�D�8q�߄�o�a�,�]\�u�\�w"|��ާU���u�4^��FR8�,���#vx�x��\�+����ݬ����*�wA���O6l�g]x��cţ5�<*&f���С��3��3]�s+)����f�s��ѕ�� K^|K>�k(Td�V�������{w��-ƴ������,�a�3$J�P����FK�9X]`�� u����G���	|���"�99��{�p�U�Y�b\QPiN�k�,�r��9
 ���k��&/2z��|��59+�3��Y:6�d�l"�K%��ޮ�OB�g��&��8��`���tsm���j1�"��O8F��X��<OF�M�ts��yrz��}ٛ��t�H����28m�*Y�v׈������']N4��h'���s5:�q^�ڤH�<n��:����]�c�xu�^��/[>4]d��_1tV�f�Ipx&o��K�%����wB�}�������Y��Qf����.�u+�B�W2]ɯ[��]�y�4��{ƈ�;Y�#l�e�c��X��C���S�Ľ���=���h�����E&�h�W���b�S�:;	��R�]*��l=�ZW%6��9�o�zz������Y�Q��Y��s�qŭ�Ǻ���+��ɩ�Mwo� ����
�ہ�QS��i�������ݶz����8ϥ���^r��[F��!�>��j&���>�*��Y)�eu�����Kٚe�����m�oxY���	2�.*.ၓPNg*ηÔ��`��;ͽ�L���î���<�9od� �r������a��@���,\9����\z�lu�#U��f2�Yrj�S'Gǥ���E�H��S��]�ƺ�[e�B��`�v��-r|�d*�!�C�zk��� �:��z�83�v�i��:��Ի1�x*9��.�O����v�U���㎬����)��K������\�I�fWPerά�[���ِaܹ�`�7m>}��V�+T7MG.��M\:�+����q�D��p��u��6� +�|O�������08��e�ZK�9��}�	�$Q���0F�R�Onδ�t�,8e�p�/-͏|�0��}�����H�9.۵��@���QE-��B��d���������o]�A��ˮ�7V5��#S��$��z���]K���>\�iL姘2�� 3sL�7���h�|���]�.n}�|�����(Y� �,�6��	`���N�{�o��r�oWRH�fuʏ��Jdc�{�N�sS3;�>�\E��%��.��U��h�b�ؾ�Ӱ�Z[AU�=�I��)`�JL9
��B�e'��]�����2�p�sӖ���+{K�KO�|�x�K���`*��v�"��zs�6�eh�{�k�U8�ӵ�o��e�.���(2=E�e�5+���I�Ol��q�����N��������� G���L��>��k"������dl2hl���>t��Z���p9[��l�}	��|.���Y����t���ЍȜ��n(OyY�YV�n��/��I�k��G��㊯,}U�/0TsP3��}�B�1�/o]�ѓ����A=���ݯ�ޛ�2�o�9o��D����1��왊��⎷��n�a�ggR�Yqҙ@�h�}���poU�7d�C�;�+���#����3���e�{��-�9�iߖ�7\[Qo-Ŝ���`ʰ�TM���)c]�|%(�k�,�p�]���9e���+6�����,����6�N��Jf�FϞM����es��`�4b7�`M���"���ۍ^p�`y.�Y"���,�-��dY&R�}xp�`�+8�4�Jfm��U�]`s����f����;��]�6���J��%׫�*bK.1�C{p�u��E��%Cjel��Es&r�/1uX��u�=��Oyvf�9�$b�0�[�Yn�,�|�K�]�+�D�ݻ�/6��v�VQ�ѽE��{�-�����O��e�$�.4���M�-4�;���v^u�q�bՃ�[~j�[�!,\w� =1����\Y��-F['�V����Ͳ��%�-�ي+��	�=qxҳ�޾����-9f�9l��<;��! �#��g��ȩ� ¶^��v�����Ai�N4�쑗���v�ؔ�r�ܦp�7S�{��
�O�U���[wF��@���L�@T�s1vxbo�e_ui-<��ڋH�p4s���:�PI�,"-���� +6棙3����M��I��栀�M��n_+��=��^v�b�_e+h{s���Gs���L�֕ul�*XF�<窎ce�wW�K�u��}V��p�d'u=�Vz39YT+`rn	�����q�\��go�/O2�| �AAm��s{�c�Y�:��5�E�����']���ɤ{��h���	��)0����M���v4[XP|Vύ��,�CG�ّ�78,.�]��גuӐ���}Vx/-5�{��������y�R�H��͐e���i��ES�aL��4�����ٮ���Ж�M��UБۻ��FwR��,G�����03��g�)8�-�dY�Qo��r���-��5qN�M�gK)��V�Փ�s`���mwvrJ��}!��DU��m�֨�C��*�������N��s�Ĥh��3W=�ns{Pp�&���wo��˼��o�x]��`}�v���-G�m܍)�N[����n^�[r�WZ"D�� jn��@�u0�e$�|	�vjNq�S��^l�~G�2�Yqz���L��'���*�k��xQ)�R5���4DŸ�}6`ھ�*���w6���㘼��o��s�X�ů[�0ݡ�l$	�u���;;7Ll�2^ks�՝�n�y��}�7��'̶d໅l�}�Z�y t>���5V��+��v���r�����M��twz#ƴˈPWn�����e'\�r�)�}�ҷ���yg�������P��%r_wf2�V|�Jg]1u!h]4N9S}E�|wbc˻�$ʑl;�PO����Y������+-����#�K���{f�1�OS�J�x�6ܸ���J:�V^�]wn��=C�%��c�Zj}���Y(��=D��i��j��%�.���]��z^����SU��E{Yx�1�����%���3|>��M(�;˯2Wu���ުx���
��+�^�1t�� ��ϛ�J�m�ܶ�m��m��e��m��m��m��m��m��m��m��neJ�Z8i�l����\�E�;3F�Y��`Mnײ���,3e���ޔ�B�Q�;���P�7ݫU�Ѯ���/u�=>�{���߽���B		���$�ߥJ���/7�R҄���{���6 ���6\����.����(rѲ��M�;���2JeVcJ�z��n�л?m�L,&�:���Rm�2n���xz�O�z�ѐ<��\X��N۱�M��P���'Srg7��ٰK5K5�`��b�Q*/�{��N��3߰	X%�.���\��GNc0�kzv"�OG���D���!2�_PGHw�	q�_\a������+���`�tk�}ո,�`��h�E��14���W#����'�c�%�{�M��v|����m��^�(꤂�٤K�P�nlq�i�P��ZqU�|�ۈ�ߕ߈���V��7_@����;����5:�ӵ˕-E�v)b\�m����4s#��f��4	��|�is8���ߓ�e,BX�f�9xSvG���G�!M� mC�v�p`����yث���|>��� ��#��]����偼�ԥ��[�\�dX-��)W��C��.\�Wn�����vI�an���j�3i;��L����>�O�(vg��n{&��]`ͦv�V�]9o��ɀ A�ٰ���NiR�4n�SLU�9��p[�WU�}݈7�K�o�fA�ੰO��>ي
��}�*�$��R�Z����H~#H~ҏk�_a6=�b�$y��Y]�7)k��:�k�iou�݂a�����؅�e�N�M�]��^��a�xR2N�1��G�R~���lha}��l�"ٲ�]��%��=���$�����8ɸ/���<b�:5���ecY)B7��Y�\��_r��v-�`�i���V�MfOz���3�*і��v���{��Z���3V^v��3}�&$�N��w����'c�B{�aG�%&ϸjRc�qdV1�r�Yc�7�I��ө��t�UҠU��.�6���VB�r{I��/q��o�;�qK���*V��� 2�3�oz:�繷���*=���{��R��ǻ!�0|��u�2�g��m��t1��MΝ�=����cC���]2��	�n��Uw'���u�a��K`�/���|��6�q�!��:� ��<޳Ơ$s�%ۺe�o5(��|8�|+h˼���lI�SU����;�$����0�*H,��q�k=Ֆ�v�����j��lVދ�/ �C�E̡.��U��
<�M;�D�$���c�h�j��mL���ӏ�f�N��A�ˇn����҂2�l|�fSc)8�8ԧ{�͹�͌������t9�RNP2�4��
�5y�	��nrc^&N>��5�Zi�f���4���8���	�px]}G={�pk����{>�>�*�^#/[א��*�A���Kc9l����۴-MA�0K.�]���u��B#���zB����w׈�0nc��뺖���|N`Z��*��r;܄��o����db�.��n�8�}��S3�d�4Rp����b�5ͺ��K{1mm&�9f/GP��ṒN�[T5��Q���I*U-�1_Z�"��_n�i����V+m�u�T��ö���zKֺA!��4�S��We�0��˩���D�.)w[��Qx�%�}4�|�ds�ϝ$ax0��	�X�w��a\����s�&��2�����4"�T݀2�d�W�Cw���=d]�2�=�9Wo��a����lʱ��Ku����m��js�q��U�޴�,��%6&��r��*왂��p����e
3.,NXه�[�(� �fo[�Uq��dܳ�xL��u0�2�'c}7d5e��h��P���U��lax3)��:���e�n��Z�9�ز�I�����嵖"voQ���Ұп�cS��Ev&V�7�uo�;�ji֭n��fm'ݻ�y:��k.snL�U��T�0N�Րh�)�E�r^���m������(\rj��'Z��o����If�Mw��z��'��RόW'*�fT�/�)@�u�_jR��+a.��R�q���워�ݽَ�E/{����y����³To�9$���Ě;$��<H;w5m'��QV@[ږ��i�����S[�_M�f4cJ�H ����8��e�+q����w���>�]*82�%&�Q��7���I��1J�G����NJ{���;r���hS��|���c鲙�J����P|j:�'6l�4u���潱��������F��1�m]Zgp�;
]+$oH�H.�9���3����om��]��'Ǡ�}��R�Oh��m��|1F�_!Xof��h]��D���>�.k�t���(�;������;���"�/h��&��B٫z��{���ǽ�iխ�l[���ݶn�<۫���2b\F2K:e��#�u���u����̋��Fv{h�K&���bh[��� ��r������H9.fּ��q���)�� �[������e�)=u�ۘ)�_��!�3�Vi�qy� ��������)H.���t#d#|�e0��>��Gϱ�옯.���>%�iK�+���軹�Y+���J�x��-Q<tحΦ���om��q��AU*%�nM��2_+�M���5�݂W4��k/$�6m7����_B=&���=S�������o����3Ֆ��� v0���A3��W�F�w.��y��\@u�i���]�L��6�T蘥�o��N��N�X�a�묟,w]��=�GJ�ȖJ�*-|i\dЍ�v��R�2���k�qK��s�/��1dFWԇ!j�I����	o����[�
��.����y��xKv������V"ݽ��b��c�·7{r��7^�Z<'^Z1���]��e)KM���8�P��]=�]��k@�侭�Ū���ڰ;x����6ܖ�o�o�=&�x�a���G�Rd�v�Ea+'z+s�a�[�}����!uc�v~n�b�9t�,u<�����2�_s�#�d���&���L]���p1@n�K�0���p�'��*��A�/UqO�Y�$5��x#�b�67����QN��)��C��$wqz�!��[��g_a�q��.F�f`��-N���D��W�ݽ��1�z*[���\)���:b�SE��]"E@�y�3d��\#�c�`t�bs7��O݀�Gkw�QTB2Mt���e�%E�n�*V��2;\��*r5�0ǻă�d��3�Rh�������9�w����	�D �n���0%M��ۑ�P��C���}���.{�F`|��L���1C( -��g%�{G���BT��Y���鹽l��e'�I�3ϛ#HքaqD}�P����ՙX�aK8��8.��^*�$W�F'-VVx����U��#\vv���_+1��aG2	:|�Vi^�L}�Wu�Uz�p�#�)�h<]6+�ATBE��kC�J�����V��h��+i��m�zwe*�%�3)���w��m�
��v�m�M�
j黗��j;�NQcp�Z��ŶFң�[�1Pk�xc��JŰZ�!�A����Z��s(���q�rW�f<��1�	�׳�����n����]���iή�o'پ�od6�N��z���]]���i �u�r#COTp�Ӗ���~�Ǘ��v�e�h�{+�g׻a��r+����!�4A���d��Vѽ��{ژ��(Z� �S�n�T÷�I�?9�����N�#�g�����Ai��9X�v�w�m���F�e���^�1���_\��ϸ�vV��� �m��%a�Lj�ޙy�� ��VB���=��g?}�[a׷$92�uZv�#Hȓ��]��mK��z*3�����v��Ȼ�3))D^+��a���Iؼ �L�w\%'�w�[�	1����x�:��V�{E��2��@Vu��s��]��o���o�5Ա�*a����Or2x��uo���������bO3mZ��q
��ң�%Ԕ4�}پE�[���2�dP�R*�JvU�Y���-���߯��.�X��Q��Uf�',��;դ�vvU�m�b�<̺j�-q䫒�3 )�����V�S��H�����d.�u�l��8��|�7�� ��q�{Owu7]n��cAt�@Z����b���a�w���,��NDm��[d�&���rU��®�����ۥf�����]��oU�A�S�V�C~���}H[W�m�@�`*�Ptt�����������ѓ;����:���6�<�n
��i�f��)ڸC�|��F��e:�)ө֝����&���2���Ýѯ�uwq���R)>alG:�Nۙu��7M�N��]�Kj�����T�)��	�S=�;�gT僫@&�`Ŭ�;���:��؉&�81�ӹí�'�%�ۺ�5iw|5��d�&�4U�ҷ�8�rz��Ҥ�E˾=����3W��3#��EΝRy���oK|�4�򭓈	�K��ju�C;{�ǻ)q�l�@�DS�R��yC�a�i���)��S���
^Z�*<ܤ�O �n��>3�9n���`�1?�yOZ��vl�D>�7yMX�G�w'���sޛ(�ET���̮z{V��^�x\���m4�F���M�2l\�̮�5c8���nEF�
��6slФj��D/K�	3ğ\$��g��۱�u�n�ũ����s�;d%vw-��h�dj�gS�����)�i�櫓��g6�,une>���_|t�\�j��M(_ÅnP��3a^{��#^I�Л�.Y��AFzQ=*��Js�;xe(;i�Jk�7MO�)�Zxo��B�B��
��P��Tڬ���\̢�Ŷ5aiU�8�ç3�|�JT�i� r�G��Z�Kr�(�������@��[�i���D��P�e��K�[�x�����
�&*^i�9�eXƧ\<^�c㝙ufD�slL�2�3�xCW9j�t��4d5�õ��z��d����3b;�9]���R߉��*�H��Ô;���']�G��$�)�J�랹���]�A)�LC�霺�l�c�;3k�*ȼtK�y��9�_h����us7�Wn�I��	ۘ�!g+͖���cmh�o;����aY�:�����W����ʲp�OI\z�=�ԫB��<�9d�bL��c�r}��GF��zb2a�o�t7%�r�-8��lK���8b�MC�w.�I��,WM�n��I_1[���$�Ǳ�x[��R뙨�k����iN��z�V��w�B���a���u��styu�ѣo'�>|����o%��HЏh$R��2+�gq��/	����q�}=s=�௕�A��6��4d�<��h�u,]��T�7b��N��`v�S�/xq��h=(���:h�Q^�^M���6�k"R�>�W�y:�w5_C����Ng".�i��,��#7y4FvT-fm���J��lSgk��Yo��9q��p�L5y�jzqw=W39�ie錁G��=���D��[���o��R������u_#݉X�p���wa�P^�wh�|��9b�`j��rm"����a-�e`>�7�Y�vD~�Wz7ŉs\8���!^V������	b��ugtWN����i<�+S��ُC{$�x�ʲy�����2�t�W,,���"-R^�%,ǰ>>{cq���#�Џ5�]��V)�<�WZ�ֶ͠A�
���"��ɼ��®�v��jg1�Չ��ja'+)���`����?gK�@c��I��B�8B��s5<�G��`v)�����)�9k,��
���+r�bɥ��c�Zr���6&P;@�Ù�Lol����塧Y���qib�����-L���4[�%٩)́.y��M��:���'�$�u<�����١ƱD�\�kOR�OyL�=Wii�7j��)���b�Gb:�,W@q=k(�-%�Ai'!�ov����X�����k�pY�Е�;m�K�t��Uà�}��վ"�Я�/]1��c������N�캶
�AvJK�ɺ��[݂�X�v�q%��oK��2��|��i)eoj�S\�7q��`���,���J��E�t�h3c���})���9�X7q]��]}���.�We�/�D�� #F>�p�$��N�n����i�t>��{<O��T�Q#6�5���e�o�ǜ�=�i֟]��.ǔ�;p�3�n�����5J�̚�-������)i�����J�9ҡ���j�+�9*rP�fc#Ft�$��(d���r�fܢy��<�[5��>uȘ�nY���d��;������|&�Z�N�zFX��6���kGSϜ���P�F��Iu�jҪD:L��GHއ4�syo�:�����̦^h�g���vs0U�0s�.�S-�B[2�(!;�hwR֪T։4��t�Nv�칽��p/=�sΒ��kY�T�ް�Cqj`W9��f��B��l򡒛�"��y�w�;�����&�kV���:=YX��S��V��p���;J�i��1ꮫ'(ݵ@<� \%Ay�k�Ȯ
��Y��.`�'
-YU��S�6�[+�;���K�vRNs5���4}$���9�*�ޯ^�� ��Ⱦ���Ǯ�����F�/�'��:��ԅ�er���v����X���ܟQ1@���n��zf�����	��4Z �^;]��ڋ��[��N��>�f�{��Z�⍘��ij�X�A'�w����Ө�$G�}��×6,�3�o��v���5��ƣ��'cu[�GzNI���/ԣNb�����e��J���#1�"���ۘݗ+CO������^m��Q��Z����5�������������꯾�}�^�î.:ie��N�_7�[����⥵��{� �r�hK+*k]/��F�����V�v�4���u�g$�# �Զ���}b��Jv�m]]��ը@Ex(��󝸜�0�[����l����M��z�y��7���o��ܙ��:��������W�er�FV�kVHr�P�[7���C�9���WD')��|�B���^�G)9�%�[��ԇ���y����J#D菏;�xa9kCق��7���=�ӨY�	q#>�y| �Y4Y_\k"��u��扫.|x
ߔꛔ,)>��a�*����S�X���v���U9�Aa�΃ON�T|O$�J	,9	�U�]:���d:9wXw|��i�v�+t��E��Iwh���o1KW����g����@���[����gC�x�I�#'[���ƚ���'�-�=��g<���ͬPW[�:��Y��{['٭A!�U.~vѷ_?B��c��O�m��9ͰVr̮svR�|��	�
���Y��zs-�Rȶ��b�k���j���F�p3����%����U�����u8q[w�t���;V�2��X]�l!R�r���s��t��^��m���h��銈�FsӔ�k�z�u"+����7�r�8�v�f�+Z�@���{���ɶ���e�ל���g��m/�w6��_��2�԰ء@ > * �JԶ��X*��Qb��-�Z�ձh�m�m+c���a�����U���Z%�y���Jԭ��ڥ��Z4F��J4U�m�T���]Ҏ	YUPQmF�j�*F�J��Z�Uiw�LEV�j�[jҖ�ێ"�4Z\k�iZ���cj	R��c�e�5�j2����.�� �łV���l�V�ҢڴEU@�e�h5�Y�\km�*��iF�Z]Z�Ƣ�X��SnDF(��)*1DQT���F��#���b��
�
���e+(���j���V��Z�+U�Z�-�m��������E-Uh�(�Ԕm,b#Z��SZ¢�Q�*V��ѵmT�����q*���m��F�UA�ӓ���c".!Q"5%2�Es-�E*o(&%E�&�V.!ED[�cQe�k*�F�m��F�F�
ªT1%E1SlӧQnd���V�}�ו��_�kV|�K�ݛ�t��
�֎řG3�1�NO�a���IW���68�R����읪�]A��MS����jň5��Jǆ���P�y�cz&JU�ѡ*�Q h��\3ٚ*�
��䏗a���������t��#4��=�~�	v���T��=P�J�ҩ?Y&�aq8�0�>A���nvf�ҍ�b�]�7�g����ք��x��"�@�=#�i�_4�1���ve쎕罭�K*��0�.�k�#�9d=��Ϸ�(y�f�*��෤�COvt7����u1����V�t�{�\�i�:߂̙�ts��oKK�,\�����<���I�x�I�P�4a�k�/�L<K�|%���y'������dK���
�ނL+]	ς����q�&a�1��x�8Mp��+\�z[���!�g��{��:ݏ-�/�^az�6Fw�D�!Y�j:#����z�{�p�%C��PKV��!Gw���bHR=V��}I������S�����N����R��)��Ê�k�ݏx��ǳGQa�{LP����*�DҜe{�qi�涸u�f���8m�AZ�8`��h;j,S�r��e�ͼ���T�s�h����uz���v��&�Mb������]�bY�Zz��7��n4�Ot�
��Q�$=���b�p���v��g�[f���JD��>S�ۧ�vw�&�o<r�T�I�T^��^Y��~������9����h0Bq�"��Z�WF���&�>�� ���\(��G.n'�:�F/����^�'u*��|4mR�htq!���2�Z=>z�Q�]m��z�|�[fKҷ�߱�ɴ�W��`�Q�ϧR���ji,�#��:;�����kt���c{1g�er���>�;u�hu�ؠp�Ny�^�\ϰ�
��B�.$E_�O z�9/������B�<�`��b��T4)�z�=PV2�������BF�4zy�~���|%
�\�P���Y�VNg���z�G���K���3�/O`�r�g'g��K!�7Q,��w0�x}����[����[իh��;�Mw�/�<��m_����r�g0��r��Q'�XĪ����ͅ�w��u�Z1�����c�l.��^|��/�sNS>递�OR�]+���7�bL7Z��K�F쳣 w+C�ѿ	֍�O�S��s��Ի�a�^F��d^�>�py�`��;�Y)�Z �)/�z��ĥ`�|vx���;(�&�m�nR���`��	n�L"ا�L�X��ޫ�Ƚ��q^�ЩX8��źn3ݧ���b�9��y[{��o',�Z]�{'<�0[K{�ٵ�9��!fS��]î�ݭX�kq�y��H\C|��N���f�޼�!�{|T�ь��Mnc�S3*s�������s�8/��{b�E4�\�ӧ��m&�U�����:���6����%잫ޛ�K\Ž�MB���C�=2������~��z p���u��ɗ[�Z�H�+�y�(��uoL��Tw�~7~�0�iYh:8$�`����N� Ҙv����wu9�̰m;���{�o�1�Wy۱c <2�&:|�3�Ixi(b��,1Hg]3}r��]��2�&��C�<(Wu{գ��涡|����k��t5Z�)}�e�]�&r���}}<�Ҁ[��+jv��-�ٚ�y�- �2����s�O��S�u�i�CO�'	���+Ȯ��o�����\3�9�Z��)e�${e*�}Y���xK�T�=��ʱ��� �%��׾0g5|�oU��S�7�آ�P.)��˂�6Ou���ʘ߰{"�ѿx� �ypUCycԉfO&��WR��
���̱c��9E��-���X�N�U ����;�d�1!�/�ozWN��6We��X z�� T+��4��f�A��o�-�1g�nox-����O��֎S��ST��=�O�n�I�����:�r��l�	$�9ݏLG>��O�lCr�x�Fm�q73�w�����`L�/ac�'}:����A��̇�w�u�kjS��okwǸ�j�M�2�ҡ64/ڹ�6�����{�*Sʊ��Yd��u�|(:���S�e�V&HJ�ԯ�{f��m�^� �ǁ�SHz�K6r�MS�oԘvI>����
GS��i����X|{��,��yT9X;�$��)�D��	���L/�?E���<�X�)uI镈��t�����T_�d�Pڰ��޷C��Xފ����d(��.������CV�噜��oM�*{���{i3���ZSь�n^�.���]yƍw��=$��j� K�Y��ϓc�z�um;-Z[]�w�9�]���<�Џo$%=�x`�c��H���
K;n�h�y��*kc�5d���woʰhZp�.��y-��X�wR�y�d�n�};R���_��yd�.j�j��w��n}ɆO�Pn��Ua���Ce����Bx�9@�g}�8�l����Ԝ#�ף��k��ܢ�<)����D���&��aT:���6ϫ�F��֋���-i(����R���Ґ�d�*�ި����斋��^#�J��zo��1�v&�z�:���/��qg$��0K[h�5�>�9��5kP<8-���m�D�,Aw�؄ŕ�Ҭ�0K�D�ǥ�uo���c#����UcQ2�OtDl�}.B�h��{3j�s^A�;�\N��,*���S��o]�]��6�/k�*}BY���g�nAF�L�1҂nl��.��2��|r0�>����]�����&2�H�YvF��N�)���ߢB���XӔ�n�	
o!ucpP��
�˜<�gN��)\�Ʝ8]K�E��4k���j�r��Z�"*_S�#l������}�A���>�(bɘ;�I�"�s�	Wn�8,B��A��/e<��G;�g�����o�����yZp�	�B�e�8���EX��%[�M�c�O��T�۽B�Q㞫@g�l��J~u��g¥J�|�B��L�8-/��oy�1�x�{~�X����:�wO/ ���e<���@���Q�2�T��h_f�7q���=�+D� ��iv�`�}r�ǝ�~�n�oD,��Fn��
�*���<dR�hk=~�7٘���`�E�8:�ȯ1~8�nu���^��W����E>�4��������J�y8%u�0\�{�P��8a�k����*a��P_�^�}qpr�Op�W�{(�l_d�v�д|����]%��N�l��-���9=�P��4)4�B��0x����7X��;�܌qN�"���-���+�Ͼ\��r[��{�]������e�FICu)H��4���J2v��CY��p�]��"]P�������n�{v��m;�X�:���Cs�c �b� U�����i�v�>Ks~��R���\�m��.n~�����4�P���#�`�%حƣ�G<���k�B�Y*�#�gj���7+���P�f��n���S��ۉ�w�lhsi{�u���zx���##հ����,�!�8���1B����*���S�� �!�>޻�ܸ!^{�Y�Nf�ce���R����:Ԗٙ��A^��@u������0�UJ�7b��V^���Tv_�i�-�'U����p�)@�'��t{�|�����E��l
�޽^����F��cYxc�}���b3��S5��vt��C�pp��onA�1�S��#�i�:�z��f'6��=Y9��2��au)��5B\H��<L���w7<9L�t/3s����ษp�;��Tۂ���6�v|���#���	�՞y<9X(1xvk���|3-��^
&�^��3�u�g)g��,�H�~33��������\�b�Z�oz��K���n9v��o"\��)�H��}-T�x����ǚ�z���v�Y��[LrE^����O�*�*-�.cn%�v������vG�b�l1k�I�T�2b.Z$�{s�N��ނ����\�aw�Ͷ������a)]��e~5�ÿ��\��P\<�ïf�R2�4.�r���ץkޠ޶ܓ4��� �V�T��ѱ��,p����<�x�:���<�ꖠ�C�#����c�"�0k]U7��v��O�t��m}�X։�����t*���m!;ݓ�~�8jr<�����q�$ǵ�4y\C����@.�;wV� ��M�ؑ�Pyz�zd�냆��>���:��c���_��f�H���J��}�����c�u鸤��^�8� �L�����j�29�<�����H�X����y�����wH3�N3/2\�7=G��<��.�$�ۗ���Ͻ�;��]�˯U�,��J�9��K��ފ<�ޟ'���}�����^{tlE]�;8�2��.6{7��snw��GK�'N�=�jr6���^����i�[���u�d��6�˧������*�Ms}R��	%1UcQ��ps�/�ϧx���:fj�{�X�n��vw��Ǣٺ�n;o����Y���n6fh0u��]X�"�J����s�i�S�ᵹ�oW9D�L0�T�ŝ�>ܺk���;R-�����mO�ڊ�K�1'��Niή��T�[�'-0�VPe?>>�yw�B��s�=A��͐+��K���:w�4�=�k��:�WA�C%h�NDG;[��-�?�uI��yuxy�����O���n9�v5�Gt7��g�/�r��-�rp���cRs�L�ʫ�mT�8��U����C��Y}R%��i���w�L�	�_`չ�/=�S2��n)��1G�/��J�����Tu� /e�m�F���,$��y�d�fy�a߽*�t��D�Aޭs/�4&�{�{e{Ş�<N�����f��''�s��AWa8���������y;Xx�v�E��&:˜�Ku'/ӱ���w�:}(�9�z��~Ȥǻ�J�Ś��e�V���0�O=�g��^�6ѕ�h�	���ާ�Ǟv^ޤǨ�v
o�N���]Di4`����3�'�7"�����/�����n�[ß6���r��F񶪞�Lz�F+�Jy����W�K�B(\Y���kn�;<�����w	����u��y�)�3d��ӕ�G��Q��u+v��h�Z�H�>�E���q��L^7�^�Yy���7^��>����2���=$��̾�k��9.�^�@@���y�I.�7�X_d�+���|:vz�����F����{�\Y�1G�/�\;갤�9Xĕ�#����f<ܩ�5��|�KD��S��G��� �Y���֯`��������%��\�9�]~��r�$�ލ��lE�j%*�<�l�g�X���� ���!Ʋ��Ή������K�kx:C\�\�U�[�&�vf/-~�??N���/{ ެq���,��7�]�N_���hT�z�GH����Y�*t�v4v>sg���>1b�����O7�\����4u���V���3{ �J�_m��x��o��΀T��9�=�!�w�5�gf�n��C��Y=Y�Ka��M{v�&�/�63N�E%=/���V-�ạ$o�������з����ezw}Ԍ���g,f3�:�Kc���hVU�_4/,��a���J���={�F����)Xn��
nv��w�l���q�nl~����1 �G�T�$��/�<y��oo�|+�x�(=0�|����gT7�~�<�rx�</)w�M�F{"��#���@�3�;���E��NӺ�kD�-{؝��1�{���ɘ�,β����҆Uҷ�yٞx�{a��zT^���J�$E�8���z�S\Y)���Q|��t�=]���qYKP�HF3��7���\̘�y,��b�u髆yt��E[�q�����^��,�N��ｰ3�>�}]iZY|oչ"����+�w�t{�'z�:�|$��w��oc��k��U�����R�	�bJC����7��tdE�+��pf.��7���Fơ�;8����Z�.��ԀR��|VVC�K'��bf�����P��Ӈu�-�ѱ�`t�Ǡ>�~���O"�ZK�Z��kˋ��!pd[[�T�Oa��}0Q<���C�m�0y��7R��^J�h��y��E�՜�LN�����t�X9�N=U�*�I���w|;
Ds(�}�C8��+@яu`�S�f���xzm�z�Lf��80�T�.	�`��Yq��Qُ�]�Z�?]��Ó��4[:�t6\���u���M�mbg-��o�C+NY��b���0p���4Mv1����(d.�0zhIRg�\�~�wb�8�^�k�0�l7��b�t*��aM�b 9洌��9\��qw���{%�\��b�֋����#��^��OHӧd� �Nh9�f�{�Ӫ��<׾�p�m@��+/6ΰt��J�oz���Yj�M���j� %�,�N����*�b�V3�����(,�N1O��:�/��R��f�wq����{n��]���i�1�1�H�dd����DI]�k���/纕��YGi�ܬ�N�[�4�,vY�9]��璍諂��D���Q���+�?�@���j�xIc,Ӎj(f�zB����<ο-�d��ʍwx���&��C[B���8���Lr7{�����nS�R����.�����R�Ȳ]��V�œ�Y��ftEq<	�d�U*gt�:J7ۙ�ÍL���y2�W���rc��rgL���JӅd� �#a���Պ�|o�pf�v�ZUV��>�3G7�dob43���8�_P64�:�\;z�6b�aPv��ܽ�n����S�N����dfQf�
��B1M�G&��(��uv�Z᭍��R�F�/��}�j��l[���fV%�H��VN1�Χ����f3�)�p�On�	։��Z�Ĵ���Q)�<Y���'SΉN�p���;9W�S��Kq�4��VQ=3������y�V�x��1�\QW�)�7��ϔ�o���>g��3��̪��Ĵ�Rx��6QP5+
��j.��303�!�%Q�Oxڽ����� �馰�w�X�FL�G��KH��.2�CsMH��;�޶����m���7��
-ɞ�8��>�.�~���,�K���c�9����(��X�%v�+كX(���V3�4-Y�m�.��'u�oK�ז�y{nJ�x��N(8MS��)Ĥ�\�9�|�<�_�=�Թ�_,0�6�ȳ�W|E�i~��e�%GX6e�󝡂����P��"S
L�[��{�qβ����>���u���������$U�gdL����R��s��(�*��:�۷���`j�[G&ؼC�#W�Jw9���������#�̑SuÛ�M�%9��(rȔve��3�훃�opާ�U��줶�l^@�+z�F����� ���lm���3%���c
�I���;K��sT�4�a�9�^��6��i��k��~
]F���4~�J����Q��Ĵ�l����4�J��bZ�n+C�EAO�.�b��̗��asI\h�-�-ũb6�"%�J���c������\L� "řimQAEr����X��2�%
�E���b�k+hR�r�b��%Q۬�"��F�m��MfU��J(�U�m����YUFUZ��J���Tf\I��b�K-��,F���U�]��6��[ڋ��(���Rւ�D�
���D�
Xܸ1��A�D-3!f	E���X��fJ	.a�)ua�H��m��U�U���ӌ�iX�j-l��r��U�T�S�3(c0[E-lLfe2�
5�"������c�1��QQX�-8�QA�j�j,Qa�\��A��h��D�e�*��0����T�m%I���r�°m"� �"�1�ckE�e��7��u��G�O;�5��0�1nw����֗����L�ޥM��5��:�;��ZJ!a�٤u�\g}ƺ�F�5����������}Yۜ��������5SCk��\K��ܳB]g��~Wcn��P.?e<s�d��𙽋i	�!��ܡ�=६��۪B}]�@��[Š��7݀���6)~Qm��D��܋�hɊ��u_ǟ C��l:��:���Y��ھ��S7b�2��5������z�V����68*.r/�^a��r�����rz���[��=�]�l,	�;/;*���b�z����vT�A6��^m�y�p�[~�ҷ��N.�RS�_t��vV5�f���V�B^':�ߟ=�=�_�yzl�7��`6#�!&<�m{Xw޾�\u��fy_s�˅�N�{�j����>���R��z=]�~N����^��X��I��j��Tٹi���I�7�5z(��qԯ��3�����d��e;��
���'��cW@L.w��w�����t�3v��� ��
^`c&��A�j�3|�m�YX��e �C���b�Ehg}�f��c�A�����w�y�Sنg)2#�� ɋQཁC����c��K��1[�[��rI.99��a��?nߋ̣4�K��V�5�-��z�`��5ֽQ#~���<��f�c^r������	����r�=�|����wL�'7w�n6]��F���(:v{���{��/��ms���'=NS������@�5����K���=��N����	<�fP��x'o%�v�'܀����������x���~���dKsrm[�*RC'�y��WR��v������P~s3�+��{��{�tfa��dV�=��m4�L߯���
��s���t��S3a��6��c�w����8t�<�7��I�vT7�Us���-o��К�j,�_a����u���k:�;+����0D� �8���=�X�;��c_�y�Q_&��wSZ�Fb� �}�U�/����`{����yҝ᝔��J�R�*s�z$P;ڍ8��K/��k�m�$7�֙��\�v��.����o�7��d��n�xN���V���b�ꦹh��5m����[o3���7m���f�N(g�,0�hǸ�9GmJ�4��WzS�u���6���Z���;m�M+���f��l4�eWIT�Wx/���պy�	�o��)rq�^K*�}�3���tՙ�~�3z��X�0�p=�T��Ӛ��>�᫧H�_��>���pNys���Q�r�:�c��;�v�o�\~����I�@���w�I���s��/Def�^�jw���{T�����WM�y��f�s���c=9����u���ǚ���]˲�+Q����k��uE�/��"��ی��;�g��R�%6�QW�k�p����ݴ*(�[�WwPz�-p�3�Jz�N�+�yɹם*�����X�����3<z�����Z�-pr��ĕ��w:g�Ǜ�8f����w�ݗ�Z�6=[M����;���st����=�&��iWx8z�����?��޸�����_v۰���S�o���En�x���B�;ҁ�X,}�$��WC&o,�KT`n���V�B-���*x��*5X��z-xT;0�a��j�k�o��\�b&Z�r���Î.c��Nj���ˬ�+�r���.[�c:;��3{*��w��G�A�Kۖ�סWF3f��˞�tZ�w�����yݘ�>QV�w@�S�k��v�t����^�%�����w=��Vozq��]��I�;�oT��ծ�J�Ԑ7k�������}�����d��!��إ�p�����v����մ���о~}�j�'YP�������t��</���M���d��5��H����@O1��Zƾ�o�<n��o�s#���pE����g��n�{۹W�o�V�쪐r�^�c����{bczҶ��Om]�je7�џo&���]=m[C���5}o<�;Y�̠�ó���<��1������:g�����ߝ���y�?��d��d��'�xfBx�d�ne�RO�׹�e�y�|�i��{��}�>������c��yO��N0�'���L�A{�0��:��}�PXOP���u��P�<�O|��T<��'�Oڿ�b?�?5���O���wo�~�����~�sx����W�*�����|����XI�ϩ�4��(j��d����'�:��y���I�<��:�ĨO;x��OR|�<I/���n��7�?�����Xm)�F�n��ѷGj^���d���Lv?���P���F�B���%B%��xYVW;5�M���y<���l���]Q��Ix�m�Or�b�����=�W]d{�x9+Wg�P�A��OC#��Ѕ_
�zT���v�+]'�֝������޺�4��{I��4�Ԭ���&��q�~J�oXI�&�b��8����O��'R�����I�6sY:�d����e~�����������+=7�Cs�Z�F��d�����x��䕓�R~jM$�7�'��'SygO�T�߸Ad���Y:�ɳ�a�I�T��J~��˯ؕ{1iE1��zL����a�'�=d�s�8�z���י'O[�%a�!�?2�u��YɦN&�)���:�� ��?O���'R�>���9yOO=׾�����;��H��N2�}�H,�0�)��@��_�=d筒z����$�	�l��'�Z�Y8�&�lP�'yLd��	C=��j�»�xa����V�����?`z�Ԭ����;�{d'ƹ���2i'9`u�M�rw�!8ϙ6wy
�=MsY%I�CP�|�d��������)�y�����nv�zɤ�I�O�S|�u6�1�P�'�6��N�C�)�ORM���ɶM2w�`�$�&�9�$�m�g|�V�>Ͻ}߶y_���_��ܼ�>4Pm}����Xv�:��:��I>I����}�I�o��8��Ԝa�;��	��3�:����;�x��X�'Y�O�6�9���a�۽��V�&�~.��N~��wN���YUl��h�xJ����J�Ԭ�@�'|��a8��k~�:�OP8�?sW�N���ì������'�'�oY����۪}|����^���8q�i? t��'�OX��r���wTI�<9���a3��
��VMRq��j�Մ���~q'Y8���d���l}O/����؜��o�M�;���������}��8�8r��Ğ {;܅CL��Y��C�~d���Iě�̒�I:�d���Y8��'uMꇬ�Bo��E���>J��$��;�OJ�-�Z[�9�Ӳќ��]�9�d�ϯ����NRm&���p�Z�iڅJ�h����^����Is2�̜�/[X�Djwn��2�}��vcQ���� ���.��]��X���������W<�盛��>A�������*���d��&�{��$�X{�p���M�6��)��
�? ��Rx����i$�Mϼ�/�I�a�"��ĞН_����~B�	��w�D���_�e���=d7�2m�R~����d����$Ĭ9�:��1��d�N �;�6�������C�?$����	�K�?J�}�o��z����Y�OϾ"
�Up�D'��O�s,>d�?�g�d�!�)�:ɴ�a��́�6��/��a'�u��>è,�A�0�'�Y�0�'�|/G�{�(� k�~�O��Ϧ����m����ԓ�'�E�O�>J�~|I�{�:�zΦ��Cl8�oϰ�6�ԝI��2N!�N��{�~C�7�a��$����]��Z���߽���N2m+!��6��O�������&���8�����Y4�Ĭ'�Ri������T����0�|XbN �{<�$����*��������1���s��P��9�>f�O�}�8�������N�|����d�'�g<�+'P<I���ÈVC�c'Sٖq�~J��!��� �Jy�ylU���
�Yz�s��]������~�)8�Ĭ�?sq'P�S��	�߰�'�䞲s��'��Nk̓���p�䕓���+&$�?e���_}(]��V7�*�[��w����_����5���[�:�Ĭ9H��'R��;���l��I�^d�~d筒u�'5d����������J�����ƞ~���q���@��m�ve!�4��o)�'�3�M2Lg�2q+��Xu���<���'P�����q�L��猛d�~rH���������pA��7]q�����_}��5�V2��aRq��Hz�Y:�+	�N'�p>f�Lvg��s���^`x��N������8�z�������~���QO߽*�&���4�g����,�����O��r]{����w���[�߹m�Wa�EX�y!���PQ��X1����dc��2b��e���"�cW�v��ߗ�9k�#���.��t�)����gF2E��b��ҧwX�O�9��y��α�\���V-�q�٫���U,��+��ԃ����2y������d�	��>B��
E��d�~��>I�ѿp>f�N3��:�I�?��'��ߝ��v�������������|~��'䓾�8��M$�d�N2x�o��!>f�7�2,��sVJ����ϐ��Jɣ(0�'ɹ���S~�}�I�o?h��\�.��k������9!��O����Iרy��l�0�>K�:ɶ�<��I��'�6���i�Gw���C��T�&×�+'�Y4e�d����^6{k�3�A�}�|�����8IY1<݇�I�N0���
�ɴ6{̜d�=Cɝ�i:�9��4�����a�<Ag�C�N,
��҇��>5���8�[���s����oy�$����:e'���>t�5C�X��Y:��?s�Axɶ=���VT5�ru�Y'<�N �7��*$��͇)���ύw�5�u������]׿~����O�y�J��{�ܑd��'���'XO�ߔ:��CF������'�{�@�:��~Τ�ʆ�s'X�J��0�'R����n�����~��߿~�_�2x������'�y�_,��=�Oω:�Ì�o����q��ߘ~gY<ağ��2��N���gXO��w�o�-Ǟ�c������y�p���� ��������J��,�N2~J���C�?2k���$�&ϼ�/���q�	��&��d�=M�>��'O?S��'Xu&y�y�w��7�ߞ�����aĜAzwxI��ns�u����gRq����<I�'��?r����MOw��c���I���d�T'��"��Y�W�}�񡟮=�f��mXR�Ķ~��ֵ���N�}É�N��xO��>C�:��=��N��5�Sl��;�:����;�Y:���My@�����%d�P��Y4���y�?k�<=���;�?��}�7��Ao{�V�ǋ��j^$:�j��5Y����.nw/[7ڝf�\N��5Ӿ˿�[tj�{ud�i�닌_ew"��S��N"���H�ԩ��H{���w�ż�g��N�F�S�6��`m��X���CE1���f�?��&���$��?�z�u�$��08��M��`!�N�Ow��a�9�:�a:������~��s�_�����}�}�_�}�ג��x�`���{�y񮒲c��u��L>B��:��Y��*k~�:��o�:�!��):�ԩ�l'u�2�}d�`�.����}���)���W��Z���_��z����'̟�w�~d��3xJ�Ԇ��䬜a�72����q�2�$��o^�:��WSd8���ܰRu��P�Ad��{���ך;�]w�����L������ӏ�0=`�@��ORs�RO_Y;��+$��9����!�l?%d�KHz�Rq�2�	�N&{a��$��}��N2�/����yy��s[ٞg|��{��}�o�Y8���>�@�N���'4��|�>~d�'�;���|ɳ��T��k��+�|�d�ZC�8�����>a�s�߾�W2�Y��>��}��|�z���!�'?Y�ē��<���=a7<�x��M2y�0�g<a���	�m�s�a+	�4�IPP��>B�u+#��{�.��Ns����T�2i;��z��k|�댓���d8��i8��w�O�xgp�'�&ϻ���'�ݓ��O�6�ݐ�|�~��U��J2���jh,�޳4n�߽�����d�(O��T�eI��R|��SsV���^{��|��~启̝C���ԓ�xgp��Nx�&�>a���u4�����~�/�?:;�sϷ�<�7�B~Cĝ��������y%J�a�ԕ'̬��I�OY:���8�߶m���N0��0��ho��>a1:�|�$�I��{�3�����{����w��:q�lR?}��|����P�C�&�o2N0�}�IR��u�"������'�>��'�Co�d��UZ>�}U��C�V����b�<�ݯ1={�[M���[&ݫ�w$[܀���ƴ�e�ݵ�fP\xq|��bJ㵘Az���ӵ�6v��G1�̋�{�S[mӓK�����M����9��E>]���i���N��*Q��v���ۆ���u�Q%�V����Gs����_w�I�X'�a�N0�����8����r
d�+�RI��G7��'l>�$������'|����+�ﾱ��}L}���W^)MU;Z�ߍ�{~�c���z��9�>M�q~�a=aP��$���u��Ý��'zʇ�ԇRzɯ���'Y>ݒ�C�w��յ�ߨkӒņ5Ф������j�$�;gI���	�~a��d��R{��i��/�RO�u�}�PXOP��a�N%By�6�䟙P�����5�y�& q5�}�Y�s�{����μ��8�O̟��a>~d�V������XI�&�>��m��P<?o$��u��xI�������$����Y8�	��s�d��Mz#��|�}��o_{��
�wZͤ�O��R|Ԛd�72�zϙ6��8�?%f����sϱCL�Ad��'�q��Y���N$��+�����k�Ukw�[��Ґ��E��|��&�0��=d���ԝ��8�?;�䕓�O�?5&�q�	�1���,�	�
�߸Ad�����'PY7�0�N��*k|�����i�Fw^o}7��k����k�d�0�Y8�I�'�w�8�z���י'O]��J��CE�����8�d?&2q?S'�~��.�%U���h-ů��7�}�R��o�~Ͻ���m��VC���I�T��2Ad�s�$�X~���>d���I>~da>Osy%I�CR�����)5-��d�=������ƺ��w�}�y����~C��d=M�Lo(u��X����Y;���� �3\���O�4�Ü�x��N��N3�O���d�����*OR�����<���w��o����VM���8��OSfI�N���C��$�y�Y8�d</0<d�'P�{�:��I�;�<d�L�w���$��;��M�h���<�z�oD��ɬ�W�)Κ9�gsgW7Pn��:`�������	�1N��O?G.?E¯p_�S7�`�_cgc�I+4�{e̥�7�gTѢUۓ�w��،u���p��{#�ae����Ӊ<{M�I.�T勖�O�}������9�?��'�?�k	PP�Y�+'�,5h$�O��
I�N����,�����2u�'~��z�~~B�βx�>���u��_����8�!ox8��Oo~;u�~f�<a���a'l�>�d�C\���2{x��u+%@�'|�������C�$�g��+�'X}�0J��T�?oS��L����vN5�a~���d��}���6�����u�d��<��:���;��q�IR���q�d�+&���d�T����~r����޺�?���`�ߜ��\ϩt矾����=�a1�a��u�sǸi��? y��*d��͜�C�&��4�8���*T�������̳�_}��ߑy.�����M�����]}���=����O8��߲Ax�l7=�:�*V��Xu��ns�6��)��
�? �gԇR~I��ɤ��>���ﾕ�;��?x��l�L��6M\�o3�Y<$�vj�����6Xu�����o�M��OO~�3l�C�~βLJ�\���Ltw�:��)��Oq�Ԭ<���O�3f�s���=u�w~_�����:��	�'y�Wē�s���'fXq�x�M�Xm�����0��d�'~�́�6��/������}�PY&&�9�Y>J�?}ze|���=?~���o�y�����d�+��x���G��ԓ�M��E�O�8�2�z�I�l�a=gSs�d6Ì&�>���'Ru'�|�8��:��=މ?!�q����u�OMk�?s�o�?~�8�d�C��2u+!���xì�����O̞�w�D�N07���Y4���XO��72�2O�S[�C� ���G�B���
�D
����3�{,o�~��}����~�ݓ�8���ޡ=I�6sXu�I?!�i�N~��v�d�'��������2J��yI���a�7�C�4����8�?%N��99���o4����l�:")�Vvda�T)�����XZ~�+'9�9U�n�F쪜j�/+~<�"n�|�}{FK�ZO�U�E���Jn�ڗ���M��Ȅmq��-��Ӿ�sh�g*K�L,�-�������Z�ge��,ܸ3y���l�fl��G�D�$3����^-����P�}4�9�O\�>{��,-g����V��Jv�mN�]"�bڻ�/ 3p��Z�/λ�����H�	��
�*��:Y�9��~O�)�FȂWԜX��?+y�5ܱuu�R{87���Sq�5(���cd�f��*�(��R�%GSCBL�pWk�V�8V��+Hj9��e�e����=�1�0�T�ԑf}z=R�E�["�;+#	]^�����E������)����ԯ����%=�S ���T���U*T|V�K�/I�)�f+�
7��\f��=\Q�ުC�΋�+5rmq�\�:�j���wL+����hkLf�_`|v���d+�U�ܱ�u�ۀ�E�\���1;��P��Yշ{%l��s����|�5u��{R��#�d_-��g�{݊��m֜�ش;������E{�0cϳ�r�����d}sq�.V,�YJ'>b�kvb����ݒ��I
���P\w@����b]v�e�	������Z����@��-H+ni:qv����w�X��C���l�_Q��mv�;%���z�U�D�y�q�{���esʾ�RǩВ�r�LX��;�.;�:������'R��B}�I�����J,o��̶��\��\��Q�o�L䥰v�4��F1��A���.���ؙ>���!Hy9f��q��2���
FN��9�����m�S7Rޗ�/9lC���_��
+��=��=j?l��9��3�q��@���3�_�X�H�Z�<��^�{����ٶ�>�1<����ߥ�����s;��^U徊���`s�UN]������J;�n�����+I����T��]7����Q�qcM;�\xk��b ��"l�/8��Ҿ����{�u�5�n&_܆��>*�j���\�@����h\nnF4��҇k��A������$�=�@]��5��5_���ٔꜺg�ȁ������"vpG6�ts�ݬnzE��:��O-oM8�g &���W}�b�$ڸw��@Xm��(�]��y���N��y�V"�k�[ڰ��)��i^�9L��dܵ�n�#�q�\��V��x����yĜ�	���7�^�0�V���D_Rk�Y�Y�	Zy»��Q�"�[6k�h-�?ovz����Lp�����fl���-:d�(v�=	춎	�#���Ӵ�c#6�c�7tx���ɲ�J��8=�t���aw��wp�R�9�4��}t]����KI���hs�{��[;9��c�ܴ�m���`�r�䜂���n_kO7-F��y닮�m�o,���U��{}�@��+m��*(.5iP]!E[j���h�L(�1���+\�����,�&*�i�����.*�F"(*�"�b���)�*�U�*��`��VGWL1*oZ�AQu��9eQ��`���V*1�5�DKh�Smh��j(+��9��Z�KJ�IQs3
�qkUb��X��M!SJ"��[Z�[30��,U��0qƵ�y�U�`"+��N	s1Uˈ���(�k
�vX��`�KZK�]jWYr�V�Q(ڲ�5������"��R-����)nb���(���wnB�Y���1�F���b:�:,��̥R�F�*((��V��V6�a�r�1�%�"�$FB�9f-���TF9f�SV4�7j�M��,�(4���ʕ�6b*��q)���8�R,Rb�(e�@���`� r����:�iGx��J�6v�kh���rpP@vB�.(	xtf�
Y���mƗiYT���\r������%��ݟ���	G��CԜA@�
N2u+>���8��o�ì�	��:������s�'��O5�I�$빛�+'X>��V|�}+��Ϯ�����Oߜ^7���I�.2O����PRM��2u+p�E�Y:���A@�>�N�d�a��@��'�O'=rI��/�|>��(ϭ{�u����ޓ}�_����P�VM����Hz��:�*I�g�k���&;��C��J���ad��ݲ'P�o�;�'4������}��� �e��1~ɇ�x~Խ�O������'��=��N���IXz�j��'PXj���N��SO�q6k�������s�����N2u���{�X	���{�?w[�\�tΝ�ܿfw��O4��� ��Om<��Bq�d�|�VI�s,�	�l�
��)5l�$�'SfI�N&����6�r�Y�����w_R�ܧQ����Yk$~_������C����0�'�s�μd�I;�'S��I��d'��'7b�8����J����>B�u+&�P>a�|�_� ?P͏�������m��ik�}�o,��w�d�_�8�g9�n^�l~^��E��b �5T�uY��V�v�yf�g�R���wc�]���Nι/���(��`��x��=�P�ݓ��e��E�eW�%]����ݕ]$}�l/���s�;HB^�랚�=4�|��w��ӯݟi(�'�}X������a��yc;���i���{ ��s&G���c��6�^D:�Q�-C�b�{m��(��6C�7��Anf"� ��f��}6��p�>}jf���)��J�n!�P/�/x/��᷍��ߘɝ�(dȻ�X΂������s�˚��hv>3Tb=����� �{��<�v����s��s�'��_Kq�/Ӯ�c��C���\!����;���]{�s�?WL�� ����=<�λc��7}�9����y�y��&rc ��A�y�K�۾~�����s-�v�?{�k���$��-�6�p] �s�w�Gd�}�2�S��r�>J�{d��fC�wE�V�XZ#gs��S��S+�{>rw�%|�����h�'(yv����N� ��N��{���C�bJYN�G������FV7j�nv������m����Tu����*�7Hy�=�2���	�`�.L�J�k�N{#�N}�uw/��do�`t�lwD�;[`�J�gim����3�Ry��ηl�X�M
?oSZ��+��9�������ۛ�]�'�T���z�ǗiE��S��uF�aA&A�y+��-�3��|��lĲ��MnԱ�{�q\�kr�b�4>�&_����Z����Y!���)��Z�=u���y�;S�e��t�����i��I��^<�z�9��n?��%o%5b�`w)q��8�&J�WTѶ���꯾���8�Q-��_�=�@�� [ſ9�̞xb���R�}�O���R竍h)���Ng�����|�ϑy�퇟��rw�������B/���-�.��]�lTߦ݊����ժr���1��0{g�f�#Ε:�T�ָx������mʧb�xv>����q�%�i��'��}R����;����N&��C����ν���Vl��y1^��M)�y��>�f��휦�Ծ}�8hs�t՗�����L1�D'�)%�D�O��_b�Y��51�^��^q�3���)��y�-p�>��Z�2��uo6�u�]<pe�����1���qny�]�0����^9�m��=�,��/=�b@�U��E���;��������+od�(3O_��SB�q�M�&�������^�W�%����c�s(^�aL�/9���	�Ԗr��7.��/�B���,:yqV�֕�����+��[� �&%�VV��k��[Ô+6f��s��G��y��úw����&�2��W�F!���ݧif�Һ7�p�hvI���:��9��Υ��ѩ߫諭No�]��bc���N�Lf?l��b��]n
�F�>�U�r��{rl�>��iZv*}�]!���K�s�0S�׵7���*��z��Y5g�1t��wE ���O@�=K�����I�`�����y��򊷋��h`Vx�O���O6�;5�;~����=��9�X9���f�.�=�.�n7]{*�H����7��{���WE�[�s^|fgx��to):\�w�f��3����Տ9 mP?k�Vy����a{��/���B9K�����׺��ϫ��|�Z$���h�c�.r��|�h���E|���mr�َ\|"y�ʿ�Ƌ�>��{ڟp���gN>y��1�&�ڋqW�n?}�"ݕ]#��%?�OX[�,�W�'�nf{��ﶮk].w������S ކ��}a	1�zU��Y^��P�\�Ͷ���}�ۍ�a���B�λ"2S���"�e5�Q�_)#�'.�]F]:�gֻN�q̛U�gʍ���b�$Ls�ݕ,��D��e7`��e7b^y�z%�KmkU�;:��/HeF�uq:�t�U_W��ru��k?����l���@�����ǫ��kؾ}<����r����j�����/E�G|�{Zk��Rxn5�OU�t*��5:���n�GQ�X�@�-��n�L��ٵ��y�;>���f��0WR�r�3K�w	�����^ϺG��'n}y�t�"����(��<�w�k�o������m�X\'�$�����Sw�=�(6z���u�����.��9 ���ڮgX�)cRd����<�M�<ini=2�3��w�=Z�!ph�=n�_�b+���bO`��K�I�Ǉ,����}֣���Z}R_�e�]������w�����\�%���W�O1a}L����>�y�y݋j*�hhާ�9��ky3]3ݷ//~y%ƭރѳ��Ka���<�#�^��vv�/ׂt����q�]����ے�`E�Y��
���/ �jl��J���s�� �Wf&�1�����	C,Y��q�ݓv���������㏞Wj�Pt�+�����ť|�3��N�V�=��-x/3��p�/�+�V#�##����M��������������أ����{})�̓vS����{~�D��_;�b՘Dڬo�W�{s��N��{֮m��y��Z�Fb�*_{$��A�o�1�N��;�O>�ѳQ�v �k��yٲy����:I҇�T���KS}�{��@�z�mc\�*���e����Y���7�f�jU�;�YW�4��rV������ygm�T�����������z�S�\gg���e���Jt��&=�=aj�����8�Wzw�-m$�&�Nyy^�A��~�j�W� ��d]�k����ʓrq��f���1]���T
�!���_Hڜ_;��#���'m��Z=]�Z0�dz�����^�0-��w9X���
���{���eu�����.c��/Qc��\ͯ3��k����)ds=��w�5{�nŝ�A�V�WD������3yXKD����oUd��X�U��{���4_C� 2Ժ��f�����8�ӡ1��i��gi�'�X���w����Џ�O��ݹZsU���O\�
�r�N��BkAQT]L�MP�-N������߹�.�{�+��'&��i�st6�}V�1��;�|�#*�]������ۍqt߷��[��	Ͻ���u,jhm`clu\�s�[��~z}��nG��I�3�9�d�3%4�y;�|�}�hV�u7��P�|��ɕ{�Cv'����V��X��ϦG�.����2ǃ��c�o�c���w/({iU>p���k��5��d��b����L�P����>���a�9ݹ7��أ�pUG�+OW�~�c�H�(���y��7x{�tr܏4�^��*������`���V���������55Y8)��jr���;D����v�J���|;*��;/�������m��O���uW�os�����Pq0�ԇO_�[C���7�tG���X��'���|�ei>>q�`oN�@o��ǵ����m$t0�7[�M�E���u�����C��Y��Y�o���:��R�p�f�{q�C�+����`����ϫ2���,ݘ�鲄sk�wTO(u!�-��G8��Л��A�a!i��%�O*9�s%��`�]�.��z����n�0�t��}��}�Jϱ��Y�7�~���g�ݬ����L`ױ>�W�u�w�Z��o�[ߝr�md���=lɠ�_=�i��Lg�H6�G/˼j�V�2|��Kpiƫ�۾���:��v$_���r��S�e�P��*�0W9�ɨԝ̯{ѭ\�����"��-c��z�uǒ�%�JL�k��qaxM��y���L�������e�W�go,�ҧ>v�Ǚ�O�`Ix_�U�G^bJ�_9�=�p{S��>E[��'ʮϲvױE�}��ٯ_��\B���7K�$�|6o}��i�����<�/*w�o,;������xm!� G;o"�����9�l��s�u���zȝk8-�y��n��)�sMT����uϑ/෋����{�9�%��;���+���d[y�y��� �;P#]J�>_��_\��,k=�������P��^
����e��z#�=�o�P�'ƕI�XձJu�R�+nbZ��}ٵz��KP|&�;2�˷�Q�пq;M�pJ��(�rd�4bvu�&p໇t���;��2/g��e��#zM���E���}��|>�ǽ�6=9^��$�b�^hr-$ۈ7uH7]V\�>�B(l��6���{<c�u��و9��K~�����{X�
�7u�ar^N�ȸ^��KZ����ϻ�^��j|庐?V���f�~'2��^}��d�#g��,{R�$X����Sz~�ϣ�dS�������K��oy��a�&��[�a��e{hqZw���L��|�1�}���k/}L��<V�`��K�=����<��.=|���Yi�mɗ��Z:�}���S�Qͮ����ü��~��:_dɻ臨Ư����l���wբ���u�����O}�-���58�����I�y��N�N�no��{���s��佊b̯}{N�pr��3.mt�c�ݗ�&��^�ps��n�ܛ3���}�.��)d�[�V1%p��N�������+\<��G����_:J�<�MwRy��!ZT�}�:m�mB6����C;�bV��'��t�ٷ��7W ��H�ø�^!�t��
���Xd��>��}�mx��c�*���MP}âVby���ɦ���]�(d���꯾��u��zm���w�z��Q��`��&�[,����:�2Tg�,�.���c�2�߲��Ruw "����T8:T6@9��z͞�ځ�|�W_�K�d�{��^���`)��&wb���m��t>r����S�{�h�623�����$�}�>�y���ſs�\S��f�ҹW1G4xy"ߟ@.�	����T�˟�a8Z~�Jn6Y���%�I/ʻ��7�,q��n���z��
���^�f��>�K[�(���IW�w���L_�TJ�L�ڦ��[�V�5�{,��vl��ovUX�#��<�48^�G;+�r{JwSxvU�<NӾ�mO*<��rr\���
;2�1h�1�򅹸u>5>}¯���p=�O[W��kG�Y�m��`���w��V,�m�Aħ5d�>�����=�{^��g��yCe�o��E�aG2<�&z��3�t7����}e�CrZ��[�)���`^��ڎ�7ʛ����n}���!�qqZ�@�%^��&��<0Udu�.�x[Ә�E��ʥ��2q6��l ��[˼Q��]W���FҺ�Vipu�}&��=���wZ�g�!��֥��d<��c�˄��\��<t��%U����y���z�pn�9������+&g
�-YTe�	b�Ïz�S��ʋ���t�x�F�kn$�+١�A��ǽ�8��"c^�$�OE��3�v�a�r|�9���.�f�ɨVk�$�V�%��9��5���X�*ë��^p�(�r��G;]�u�a,��6]�q���zZ���MfZ��L���=�x�Z�J�'T��z;�V��9�u*���^j�;Hw٣�^7ؗ�SIý�<si}T��h�y-�����2�����y(��4���L�W���f�=r������+]� Wz�*�8����x:�y�`ϓ�o1s|�{����e�:\�z�W���Wup���)�t��B��4�ng,FC�Z]K_R��K8Nvf�����q�O��熚��nG�|�e�ݛ�2�Ǟ�y�}�s�weA*�w眸���%^XB
l�7��Տ�D���ј�3z�m�*7��n-F�*��sU�F�T����ƯOn��~c4��h�7}2�36�@��}�No���gܳu$�|5����ucP-�)fE��J#{����Jx�Ԛ�w2����/�%6��c���5|�\qD���y�:n!���3Bs[���y]�.+�s4>Rԧ����Pk3Y��{����f<昴��pX�b�^o$�Q
�v-*��t�<�d��9�&�'o�_���ƶƽ�=,�;����t=*��.�l���L�	8�ڮ�C.��g������ɽKOj�(uv�f��M�즚2;���K���(Knٴ%Nq&���&s�uA�D�΁k��D)
C;j�M޴��&s�R��͞꠽}�7�����(z���/m�v�d_{7Ǐ:��e4�u���c�07��ԌP˖����1JC�}� �e`ul�I��6R�Y�N{��rα �J������aV4�r������Ӭ��3/ՑJXr��=R�#��<�Ж��.��O+;N5�%ؒ��j�Ы@�#�ӡ�ޡ䷗��ܮqk�ڂ�!r���jR��b���p��ԧc�W/�9l�Y9�;�V����\�yA�)��.ŧpE���FGo>Z�yҦ��}X�<�U�8�ܫU�lr�q���@��q��%v$9U�Ʌ��ЗX͏dx7ۖ�?*��;�H��:�M'lh�"��+��'b�F�c����J�w����gM�����ف	Ϟ�mH���pV���v���s�ݻQ��(�^w-�6���m�٪�rW����A ��G��Qd��O̢"
�i�XfQ2��Ub��f+��t���E��8�J�a*;�Ņ�M5�YU
��`���XLa�kb�IPmTDaU)F%���ȷZ����l��+*[h����(���.%J��Z�R��"
QXV
����)�[�ZiZ��(���
EPX��`TYR��1�(�Y(��l���(�J�VEF*Ĵ�T�EE�JԨJ1�aUj��E1-
����F��*�lӴ�²�H�Y��hU@�c�RV��-�UU
Qb��*:��FҪ4��̓�L�j�إT;�>���5dV�u�o�{lH��s�c#1e���{��,zb��J;�Yr�z���^il��K<xv�e�nR�ǭ�1w}�}�}T���7�Ц�}M��m�cq�3W����pɝ���ެ/{�;E�s���8^�c2�3�����L`] φ����㬒o���v-�$<.wn������ט\1��3�`+ah�.�*jqqJ�^GY���:�E�b{�
o{�"5�v���Iyք�3���-pr��(g�e�Jff��m�~�:���z	��A���o�^��=m�졧|w�u,s�e�����]��l��Վ��5ʜ���RƦ����{�Ցc���]�۔�l����������Ǔ���E[`;�Xg	��z��W�K���۪B
~��-��|\�ʙ��y�Cyy2<Y3��Wp�i�;H��陸�#���h@2V�s����i��~O<,\�ͬf�f�"��K�Ҽ�O�g$;��5�Ut��l<��t��J7,��=��xn̿k���9�7YW|��{"@����Oy������/rd���nvI�RM6o��LP�k4�9?��=�{7޲Y狮C�5�>����Ruu���/q�L�d���ar����h*,�du4���q�'�	���/��> �&v�5��z���[}��ђm�"\�=�B=�N�v��z%l�(�}-����N{c��Z�#υKaI]��{��pr��Eq4qo��yF޷��.o�q�N白_��B�L �~�:,���l�ϻԽ��%TOJ���E\���;�f<��q��ԟ@lc�s�}]5z�pC���⇢�ݖ-��gg�=�g���g�~�sS�b��8��|�f`�gz{Oy5�a���T�J�/�y/��_e����yt��@B����������xM����S#���g/ Ϋu���hW"���{9.>BӞ��z���[�����/f�����^~@������_�u}ϴ�F?p���iu�`�2)z8�Θ���=�񽡶�_�����R<����f��P9�A^�r�ĕ�d���S��{S���x:����Ҧ�N��e�����	��L�%#���ŔGh���R����:˚�'�A뙠��W(�`h�N�V9���=�����Qi;����.tjǎ���sx���A�;7\�]�p��O��^>"]��v/v*/���o > }��M��7=j�:ϳ_�N�1�E��k�����+9����\#ȷ�+/w#�&�����U�j!�
�^����yN��l��}bz�s�w���Y��O���&T����>@���h}��~�*��j�����+_{����n<إ�t�M�����g�"�v��]ثo��%ɣݴ�n<�ŝ���9��lD���n���-�M+��G�3y�JV���3s�}�r�����/6J���[�g}�{ r���bYU7+2���N�;7��K���"�-�ԁ�w�����M������al��7�l�������g�J<��Lކ�=���'����y���j���+hMy�\�G��ec[�����o�=1�sS=[���J&<��u�y�Z��zs�lg>�ǵ����懂��H�Vm�m�z%߇7��|[���v�WRn�e�1�%F��~T�+�U����Lr$K��>V�+*K���3�5�@خ9���\�����V���B\㶋��s��7H��pM�z�e���(L�ʋf]p��	�;OxxU�o��{���  �}���z#����&rc5zG/��/�dݙyX����zn���S�*8��{Ӯ��4��>��jq�y��=��|׳.��u�U䨢Y珬�eËC��_�1�89K���)�ӽ�Ov�*�|�D���5/��g]�x��������>��'l�����X\��0�s�5෹xqݵ�M' ;�a���e;n���C�G�Y؈�����%��f���s�n��=�=������l��/����#����'V/e��^���m����̭p+��K�s��L�f��1��}Z�ɵ=ü���v6��j�.Og�36���yy2<X&rh6�76����Vʜ���z��*�f�����`-ǆ,�������Y�/�:�������Ʋ�P5TF:꿏>�-���<u�k}0�T��v�Sx=�����:�z�S�����]\S��e8�
�ȉ����h�	+zyv#+8,��3�dƁ5��V��&�����ϲ����M+�mIwHJ/��W��tt���3<c�-�=Fo��q_rV��9����j�a�e�RHVt�0���r>�ŭN�����u�M�V{�6o~Q<�?M���������TIĆm�jܭ�\�k���w��Xj��w��2�-b���ZY�g���~�Q��ݼ:{�8���W�q��{]3������-cۚ�����krnɛ�\�N��ۚ�k�O�;�u)1�`=~^�vVkѢw����s+׮�s�ˮ^�gg!���p=^��j�ɝ��ힶZ�D�[)���nt��	����y _��W�;S<�A��f^xG+I���o�we����c�3n�긁�H�U�lZ�{����s@�;Y�0B|%fԚ~��Oc���� ���V���굮�����Q���p�/��n4����c{:5:y��rpͺv�!��><��N�WK�(+�.�k�bNڡ>��/��{%K�I�	�\��B*��lW���O�u�)���mߺ��>}�<�,o<��o<��'Q��"�X�L!�l4�6SɴÞf	ބ$o��_�л�2&G�\9h.�Kh��l��R����ؗ	9�5�%�]q�j��-������7k�pv���]��6��s9�,1�eFpaG;�}_}��W�]���b��n���\���7K��}���z�>��޾���&b�u䉣���y�&�xX�sDs���'�T��7��+�#��";�.,SU�ۛr�p���[�֡G�����F�^�{��5�1����J�]��ikCi$�Bg�3x�T=�Ol�yN����,OW�x�LY��{��å{������:���r,��T�,����{,��(	��,��q���ݖ����o���ǍB��]�������T��k/�]3�J�=�:N��7�֧���`ކ��;�Ծ��r��X��'�]���fw�t��𾃇���{.yfL~��7������ǣr� �I��{�M嶲5/�Ά_?��,N�yGṩ�~��l�/x�`e1�Sd�U��������}�Th��/�e����ǯ�;�1惬u��p~��b�:�؜�ǾWYKt�"�f����!߳�gqqIT�t�Yi�)^�K�q�����xC����2h���="�ܱ؇�r����N�ϫ~	�K�y()��f	.��t�S�V,���A��c�v!:���?\ꋞ߾���}��������{�o���7K�v������pN��U�&Gu�����d\_���I��`����������/Y�v���ʛ���`��z��WyS}����$�=N�Lf?o���5�����όo��4]�y�_p;�/�v����'��U��+�I]�Ns�}O{p�9m�Xr�kqt��F���|P�`��lx�Y��6.��M��E=�S��OJ�ԄQ���3��_M��y]��+���r�?����~�x籆�*���:��U��7D*`}�����y.q�&T�tި.������b�W��O�I��m�:Rz��R�%ƇO/��7�"�^��T�R����6)R�7-�E��n�X�"�=o���坔��9�=� �5T�y�6��*`����X�e@}�.��c�و9��-�>p_��X:+i⮧(���0B�U�^��h»2'Z��SE��~��v��`/������~���6��l���N�r��Ȅ�#%&N�_I����-H�����S#�]�72.�n�S��%q�����!���E�/�μt�t���_}��2������#v\;C�ٵ��׼��쪱�KA���Ö�+k�/�{ҳ��o׆�(���{a����n���>��I�����ޜ7���/J�݌�u���o�t��\C����Jk������'�o��kK�ٓ�K�������K�1�gó����q�;��j�x��S}D_{��Ķ�֣��^I[��8��7}=�~/��[��+x7:|����Wg.�j+��p�wH6��q#=�e{ޏ	%F7��YW�[H��[fg����c���߀�Q��4 JȘ����zl޿o�v��R\��e1�|�ȣ<]
�K�F����MSap�	��!9誆a�-�y���xu8�~u�E0�ϟ�O(!�x�
�µ �u��z%#É�1u�3�^���웍=ȸ��s��Y���նs�k�H�R���)|OP��Es5�#^*œ`�C��GV��P0�1݃OOv���߮���z����U�Zlą�L������[W�QA�p;�ު[�Yv�Szs��J��J
�+e�7u�:E��
⨩pѕ���vR���$���kc
�N=�,���=�U�M������W�4�㓻�n��}�0�}~I���u=�)	��ݵ/��ODF���Z��E˃�A�6���&UѯT��6����M>���{���s��=r�,fÏ��t�����lk��Ob��痬Пo#��P8M)oO�g�<�>3�=x���)�V9r	n�Wh�~��k�w-�+r�>�I�Hd�j�)\��/�5�pSg��.b��]�m�\��i{�o�{J{᳕r���v"H��a�}Q`K�_y߸�J������aE��1���;˂�A���{��Pj���Q�1|����Ua�<P��=��!;6��(љ6"�Zqf�p�m1^�oOR8�P":��)='�r�BA�Y���0ˮ��j��W8h%�����J�B��W�!�rƓ��8�"#���)[H�R�E�e�Z5�YKWv���A{0�$fי��K���J��т�e�:@�矏 W�p�k���NCA��3S��'Xc�r��+Z��m?�+���x�&k �.�{���g�%C��bCo��*�p�<FmJ�F��M��D�|���k��7xЊ5�̣�U��y2G���{�a�5��]zz��Ɍ�<����d�M�^�G"�Z�!)�f#��e��h��fǝ�m�
���2�[|[����:���Տ�{6��r��U�ko��������+�9����?����#
,�;AS���i�C4\�+<z�&�@���9!��e���Ә���u���j�{�%�����2���uj������1Bzf�]9����yK�K�,+�3x\�pyQ�S��e����~�σ����gB�y'fW�q٩s���E׭���]`��F&���� ��ß���N
��=�4[��F5��]d�|Q�v��x��G��Z<�!F�Z���N����l����G��8�9H:��e�O;7�.����K��٠���߆�	�?��eO\Bx����M��q��鎯^��걛D��A�pa6B#�o���;�Ai�a7T�0�J�ܚ3��pV�d^������fvm�w0>���W��՞�S
�A۱B�]_�`�s:�S}��,+����+nw�dl��5+d����u
g,!�2}1UJB�U>n�Q4��=;�#b�Z�:x)��I3��/'ųL�o!u̦GJ�1X$�u�%��&%R���S�����{b'�N��DhL����2휥���1]WE:�I���p�	T���i�k�t��ѵf����v����%�E�w|��/�$��_w����&�\z�X����b�slcm�2��M��0@�v�� � ����AR����Z�(.�|��YV#:i�q���6H��;��o% ��+;�ژv�)]�GR��872���U��)+�*B:�_!� ��zb��:����Ճu_*"A[���`��a^�6�:�����y�ם��i��1X��� �����\	�7k��P�П���ǱX]}JfQ�Ap�F��R�X�:���B����8\��}��r�|��!��{����5��:y S>-V{���Gٚ��i�#*d�Ϭ]_k�z���$92^���pk3��z��I$˰����臽�]�h�$�Kj���;c9iL��s?3.w'���[�"�Jw�&�B -��u�D�f�+/�z�TT������3+���|��{O��|@�	��o|.U�M٦��򺱼h?Ax�kb	���;��9c�n9A��_Qn0�|������������zlx��)�>Psc���W֏`��{�;I5��:�7ou��s��=��Uͅi�����+�-e)�Wۘ ��Dc���x�*�ow�'o���q��8�9�N_j�4�m��ȣ�1�줾��,ch8ja����P�9o��������}DM�Ӹ;[zk'.���e
�34;=ݖ�Fe�G��s�v>��t�����!I�uT������sx��/l�,���B�1��S�f�'�}��+��&܁Zs���~��3m���r��ff��=�9$fM�D�J�]d�=�-�ag��s�;�2b�zJ7����2Gw�z��q}nX	���T�)�6��� �7��p��+�ٱ\������4c��>���Cg���<zp�DG��ҧ��W���5���-���Rv�RՕ.�fm�@8U]&��|i�S����k6�O�4u�]�l��S��9�T ���3m�һ[r�PԶnu�g�i(�����[��TQ�8̇�M`Ƭ�E��ܬ&��d�)P��.Z�09�e4d���qY�ϥ\q|�༽�w��r�,Gu¯4[��j�&��ֲ�P�|}J�����B�}�UX��v�%��yua��G��uß)kx�ae�4����x�9sY�ɷ�
����8b�۫M��fg�y�m�r���CV��&\ \�s8���*���_/��$T�����1��c8������H���l"�������9���	�g�;���csݒa>�t"S�ډ�Z��Y��27\_#�^T%���I�f���o��X)<Lw]7g3��9�8y���������V��D�铫�{iYM��>�][ݦt��9vmݾ7o��vu�TU�Km���U^�Z��	���x�H?6���qi��u���E�6�h*�\q���"��ڮ&8Q�k,chT+(�bcb�TAX1O���2Q�B�J��(�E�L����(�UJ�Z���LB��UH�e�QQE5l��f��B�@�W)��Ԡ��V�1F�eTY�1̹��j�.Z�$��**�%P�TQ���%���sx�W�(�E���:q���m���1V,r�UQ�C,��QEAƙh�(��c�6ԥ���qF�mxY�U�m[k
Tm�F:��\��E�n	��9��iK(��
Q��)F(�km
	�b$B��T��(��Lj�Z%�ʙcb�DM\E\mZ(ZZĵaP(�6��H��UQ�$�ho]�譣jKl�0�b�%JVe�[����m(Z�w۫9�S���k��2���
�z������1tq�\[�T:7��(�n45�?�������E�&�yϊ��K�ԼsNS�r�}	+�:�q&+C���,J��u��'��Y���}��S���ƨ-!ҬJ�1���S�X�ef�\KpX��p��=k�(��y���g�|ā�η\�!=b��{*\LpT���+�s���X<��ζ{8��l���Q�uk�>muU�<]�o�7���]+��a�y��I�U���v�����"n����9��ڬg�=��	W��D���[�ف}��'ס1���O��a�s,T�̶y�v����P�n����\�871�Ɣõ�2���AX�-�^
��
��t���Y�O�k�w�*��'$4b���0��s���{A�F�$��~o��~���0�^�p��-	'������ ^4���Ct$�S���ΤX�)r2v����s���j!�P�m%CJ�p�B�ꁐx5��&��H��Sl@#%�+�x�a�쥕#���(�Hr�u[�L���ڰO�/��fX���rxn��<gj�=Ւ�^�}����}H	u�5����p������/�9��B��f�i"}�	ux�[.U�8c���2�Ȉ�$�u�z�������6�:o
��q����@����!��Ư��]��.
��4Kz�t������N��~�����5��}��A�uҝ���/M�6ה⬨�ٹ�D�p�CI�xѮ�8w'j�>2��?+�a�����spk�c(k��hڙ/�}�-�ze��<� 
�}L����^jX~MN=G*��Ц��=
=b��mً<C�î\ã�\��K�٭3)P!yl�ٝ��+u&�K�4lS����g��LPs���c�H���.��(�1̗�Jhz�ݖ~k U��|��d�gm��|��r�r���)�R�w"}��t�+�ƴ�� ޳C��W���#��>����^J�^
�R�p��n7H��h͸��75ޗ2�G�5��C�d���`q�o�����~�Y��۹~�����wwX���9����i�/p���|�����=a3U�_[�\.���C�'��F����){<�F��{�f�|�	�^�vee��eC,��%�L�;�x`��:�>�Y�{[0-��н]�eK�ZJ���.�v�A��p����K��=lY=�}Ԭ٠]V��s
*�ge�܅�+Y�̜����ʸN��c&��n�T;j���#Y�#�\^�Iwќ��%� �=�4����Jm�i]���0��V��	�;WdR󯡮ũ�<\;F���;&A��`���Η�ݸܩ�\��k/��~}��|�g�������|r��l���\O����ͥ�*����g_�ݾ�^q�z�b�vi���]�fGW��9��¾��-�gȼ��L�Xb��5�y���-�þ��Ǆî��I�ũ����v��{��^�3��^+Q抬��z��G�'`��}�Ӧ��]�&V�P=�yU�n�NO��:��2�t�5�
P�'�K��z�y]nwL��Vًۘ/��MR�S8�	d���݋���T�#���]ڬ4�-�s5͙۬8jQ��@�6�o]�[S�/��&��r�d���f�2�Чjl�w��c�]�}�F����$�ߕ)^�~�,n���)���/]��oz�|�lo�_t�CL[8��b/�"M�vi��ܦ�)\��/1�����}�=��sw��f�j�Jތ��#t8p��J����iU{��2��E�.�;�*�
�W�:�]��=�7�g���6��S�-3T��oH��\��� ��VR���	g�A�U�{���
���r�pn�t��2^�ٹ+(L~�I�����]��U��Y��+��)JN�]�6o=4�W�yt�/��SOou	��t�D@�)y��P�:����eQ*<�S�i�Vh�s��������Ϸo��|�����������}�X�H����t37�>j
5�LR��oI��+P*��.5�2sQ��0R4#�%�ɫ'�Unz��s���|E)�}YY��*au�)[Swg�II��>�Y�OY�S�I�D���{&�X0z���{R�y<0W#��7��K9"u'��k;_/i�mcY�p�y/a{��+����k���?N�8.=����P�}\��7�)c{e����(��D`�c�+7��d�s�;A"�x�V����)��҆�X{v�go�����Ɂ��x��=N�x�r.������'�>�q�gʴ��v�l{�A�G�}K#m+]V(A�����A�ws��w��|'U����ϯ,�PE�L�m����=/���+ۦ�"�)Q�%�4!��<�4���½,Tsċw��e ���{d��<���ڬn	F#�]P:$�&�]�.���e������=�h2��/l��
��o*sk}���'ڪ�CR"�oY������C9�T��'��f-A_pv~��좬�Y�*㶇��{G*�7�+k��Y�Z�x�}�qU��=�,nQ2p e%t����:f*��=emvf��=1�*K~��;�/��כ���TMM�Yh��O���ڹ `o��B�;w�;�j ����jA�n��压��C��g�~�����S�u~�oye/�ɳ�!WY��Pn���a;���yb�E����j�5��'X#%�n��%��S;t��d%Y���w�䶳��r�Pw�P�G�5��u����#b}�>o���ˮ�r�q��Y�]%�xg��[: �a����) )�ܵj�΋����_j��-�1��&nt:��0o<K�/!¢LV%[���Z�ĪW��zi�vا���kם��!��?*�\���x�Rq��L�d�{���ra�v����7��.����f���@T��xAo�R���eV��|'՛�ķ��x�2
z���^^�c�a
�+O������<'J#<D�{(��֫J����)����<5Nd�5�M�&�t��eV��uTɋ�|ϴ�����&C�Yzs�6��v����ڱs�8f��j��]f
����7��
���`���ʾ^Hp��1�-��j��#mw��U�ٙ}3��3ք����P��a�]R|S�<.�K��/-����v.��|�a���~R�b���WO�Օ��oEɞΡ�ŕm��B�*�p���}gw/֥��Ϥ�g�}�U���7c>�X�nC%养��lsX/�	�k�#R�>����}f{��qz+��4.���JPnh���r��tG��L0�t��U}UD�br?�v�Vc�0�P���V���p\��_5;�cR�����s��;�75�����ުL8Q�x��K�)%����� ]c@H�"�	9T�9PCe���Ǿ�_�Ҵ��9�>�?2-���ح6	�,Ui�OE��xLʼԄ�}��M-������܄c�C�%ol��Fl:���૬�Zĺ k0���W#u{�X�.]����<��Խ�]��g���{}�T�{�z��Xh��j!"��Vy���ý�j��k[~WbƩ�i=X��-���X��~���=q�	��0O*�Je]S�$�F�"n�n�ĵ<5U�W�|E��f�Bx��;�o*1���^8���E6�dX:-ٹ9ߴ^VX�\���<K��+Qb�< {��>�ܩ�ә=O>�
�d��K�������O_^�^y\��;��W���1yh��>l9_۬x���E�y�KIۙZ��Ԡn�ҫ���BWr"���CuѺ���6xO�h�ί*�x&\��*�T�Λ[�X���մ@�-*�4]�EmL���=�+*��s��h���3x��o���f�A*��˾���6[�z�,���T
g|�uh󂔟-�a9-��,㮭��9�֫#�����g&,R�/0m(��.^4k=n��~��̌μbK��E�������G��7����w+��O ��5̶ �q�o��쳆���c����rc�\�]���Ŝ��^o�F�|��V4K���c�����>��
U��Lz���k�����vP�����Ko�Aw)�L����+�r�=��ÂgG��d��w�`��X�RŚc���I姞N��	�u�&�'8��ۭ%QJϼ�PV}�n�5 �������:��ut�s��׹�x{��� �0���i��C���|��}FBc� �Ș���(�>"�����6��[���O��8��Siz�7��#yf��+U��[��.��úw�,�=�v9�?z..��es�)Ss�S(5�tc��FT��x�ՉJ�YhY��|�CAj9n�9ےzջ�(O��ɼ����l����YC�'[Ñ����Ȏ����^�eƩ��gM[����ӠW��&�qJL�g�~<	�u=�6d$,��!��݋��9l{�2��S�:�1����r"R���3ڼ8	\��(A5�]�a����e������s�<�����g��׊�L���r�0F�;1(Ÿ��XN��uv��IuA�?U�X�x�x���F�J�|�3�
��K]3GUu���"�O�\Vu-)M���ufz�J��^"��P:��}�ޮ�c&{���]T�_e�6�v[܅�X����}_UU:J���۝M����H���P�u�P��Px��ۨ�1z�����L㦃�ٻ��S���/;��
���9<,5��I�vG�/r���z����F��W|/�7�9���;9�.���;�7�uL���E�������^�m]q��8]0Wv_l��7�2�p�~��d08S mH�A즐�:�4��0��s�[Y'�B����ξ�/�y5>!��=�v�foLW�yB�)='�r�l�BZ��{��	��w�c03[�C���^W��y��;޾�5�K�,\��^#��QF�y��5�p�-���,��y�k0�'឵�i}{E2}~u��]��H�(J���yỂuW���O�Lmc=�������5ىbk���1�:-���HFA�ҹ�=]	�S.4�ך���T=�m��I1�U���U�%��G6xU�M>�B�<@�s�kA0���R6����ܗ���7�W�;�c�v�/_T��jRn�C�uz;���l�� � ei�fly/Z��s�5OB����4Z�8�m6]-���UGY�"+�"���
(j]�T�i��W*�6�L=��t�غ�u���fM. ��3��d?	,N�;m�
�5˄�c#�3?�g��VJos�~A��9E���}�}T���9޾W~?��h�k�L�b�C�A�@4�������}�?[��#�=QRN>����Kxv�k�]�^6%�̲|Ȇd�� ��\"f��[�c�s�2��rY�wx��C�����f���!�.����P'��:)�34�}���M�t��#s{r�:te�J�LS@ִ��C��<>TX��*�X�D �[�r�<�4��6:��|pMm��ː����٠�O	��&�Rb_��0��u�|�񮽖5�V�z�c%�������&�~��eP�+�r�B�pZK�g��kj�
�Է=���%yI�w ����c9�j뤺o*���x"�tg��zD0f�X] WS����L՗����3�Q�Y�X��c77$:��0o<N}Q&+�n�d�Z{u��>��H��{��~J�\�B3���X�6��}�.�2r���n��ǘ�v�;Y�S��&��Ї��w�P��И}��
�]\k���ڭU��L�=%ؠk̟P�2��L�U5z ��ɬ���y�mg�Rl�+�6m��ظR#���j�X��O��Y2���m�݃)՛���
�����|�E^���Q�n<��0�ż��A��f�0��D\�ڦ��������,y����C�l�Ar*w�UUUuOgs�������y)s�gI�|�@�#��Y��5xPa_��«%_2I�M֏D���#X�e6i����[�Z�Tɋ����߷5�m�2[綝��e�#�w�.��B���u�C�
�h�Y�����bژ�Vלh���!�n��k��	��Lt�D�ά
��s"ݏ��*�!Yh:��
���a�71�Ɣõ��S��.P�^N�A�#U��/z{�/S��P�W�c>�p�W�� ��,AX�Cr��5;%xqM<�o�K-���{�FM>��;�!�XPX!�x���>2�%�Ҟ� _ӟ�� >Ȅ*��K+�Գ�gx��ڃ�%卂��{��!ϩ29�Z@�]Q��+�����-HH���ۿT�<�g����{����hFr�N�|reX��VO� N�2�psLϞ0��3w�L�o-�jxC�t2�:��NO�W��瞬�;=��5�_u*�+��;�f�Svc|t�b�r�!.�6�g����'#�����>s-�O  �}QZF���)��]�������]�Ӯ�`�=��X<j���Q�.�>�Z��n�<ԖR�p%�c�5»�LxI��9��&����	A�/0�e5�f��N���Q ʭڻBh%8ٵ%�JR���g8�TG9̪��_n{FԘ쨟W���)���nEqx�pMDe��_L�踑ŤHc�;4�6`A���2� Wt�̀���ue ���I��Z����3��]]���͔�4gmꔥp�Ns����}��惃�u�v+��Q��5b��2)}3^�n�V�p�M����������.��k�.`�F��eb�þ�r��.GUҢn�	%m���T��Џë�Lh���_ֻ�=����:��XPX��;ܿ�X����N��h�3���`��hQ՜a׼�
��3�Ӽ�&L^=��%.W_\ϣQ�/]�j�;�Q�L�ļ���g�M'�N�Z��w���= ��zE���a�1�ՃtW;�f���cxE�M.�r=�*$G_�4��N�^�(�V)��W�p̧lݣM^;��Z:�a���k�5��M'�"��7:�uìt��$l|0ힲ8�[C�׳7/j�����I��8��T�[w�
@��鞼�(:|�dRR�QY�_ �}��$��fb��F��ή�}��Hax�<�G����\�5��j��kv�tz�bS�"M�2YC���zm'5�A�'ź983֊�Sv5u;�J+�KlwQ����Pz�8a{���[�:fl}ڠ��)�jO��L>�^�-���������o�q4�+��l����fRtUl1�ck���ܹcu�w�G�G,��jj�7gBC,�v������S�}-u[�깈S��")1�B��p1��^�]���C�%�,�'^S΁�ױǵ�"%r�_ơq���n��6�;{�|�� �+y���J^ʋ���#��
�&��;[��cjnn�>�s�.�A��z���>9�,(V��>�RLkxw׳91���(��gx�����w{�d����|7�����Y}IV7��j�C���4�WSPf˽=w�n�Q��mcVi�{�{z��a�Fl�z�P_q�7�9	��E�J/uE�o�q�mrV�w�i"n�w[�+�_D�E�Ǜ�Ȩ�^/��V�G7x�0;�x5�@⾰��p]��N�kg����'��B�*����p!��T7���	��qLg:a�~�4��*d^�%z��&�W������Vh�������
���n�Xgή���S8��`R�Ѻ��Y�f�5�$�&n�^L�ۏ�I��ӌ�Ԟ()������9���)�<�c��w"d��p����ڹ��Ԙn��{}&�Gt��tz���W/lM��%��݋)�Nܣ���-��nKm��2�z�W�<���T�˙YRձ�m�q�6ҫEU��eDj��l����jV*�LJ��q�F6�J��ł0KR��mdm&�V�l�*֨�1�F#D�}pq+�ә�T1��j[d�*R�B�8�F"E��Y1Wn
�6�)4
���&\���e�����("+&�f��Y3*��ӊ���K(�mm���Kta�RȲ�R����Ŭ+EI��8eM;L]� �������Q�U��JF�ȭi�b咢�FښqUĬ*V*T�6�*�Smp�*�n)IF�����*5�m�R"	�r�FѲ�QaR�L�[mcj�h�5�(ɻES�n��.�P��[k-����ikV�PmV�IQH�-���i1��֌A�*�,�6��F�V��p�)D(��Tl��#R�R��R�TƢ?P&�C�I�ܽ��F�z�����%�,M�6��>R�w� 5��wț\82[ܖrt�[}Wum�;dl-��\ڶ���W��|ʣ�rw���<�UWBWDE��f��1kx#�1g�~�ax�\ÿi��,9ы^�ns���X���KF0H�]�x��^����x�O��3��S��u{,����3�C;��hz��G�X�W��N��I^�#��^Z)5��Cۨx�3m�_	�_^Ǜ3���}��8)M�1Y%���� �,�u¦j!��]A�����¬疮�b./��p��w�@�>�# o�e�3k<���B�bc�щ~v[���[t��>1�<��H�m���0S�T��AWK~#�x�'ܰV,T�n`�	,���3n9x����w�K�L*����A�]��Ca�b;Y��L�L�[��W/\嚲k��<�]y:���E�������֓�.V����v�A�Rjf�dzuh�VSY(3�8Ε�S0Ok��]ګ�0W����])+���Z��Ԥ#�� �	�w.��k'�&��lz|��r&�w��z}��8���Y��6�����^7�0a��r��_������uI��5=P�e[�LZ;�U3�U���^m�`~�+�J�]5���)f��㷥�8��R�v5ڥ��c4�9%���}���H� ��ضo�N�<w1<<�^gןs�Z����bW��:�uNmN�U���^�{���X��k����NET/��T��aѕO���yA=K�x��jȳ�[��Jh���m���[�/l�CLb�Mت��n��xX����L�:��/���ۃ�_�r�����P	
��j��
�-��g�~<NS��}�!#'4.�e�z����"���ߢ���{�m�6=�#����Y�, �F��o]�[Sƙ��&����#�iY^*�HU^��x0�]�К�U���({��$�#:��W�U0�xƝ���ݡ�A�~�y_D����U;&�˘p	�a��o��d�w)�	J�=�/�׻%��s�of�Ǜg,��(8d>S����0r�V���$GG���w�o:���c8�{c�V���_��^��n�h�!��El��'�{�Pb���:�4�J�XD�^�-s��TLW�gp��^�v�foL|�kD2����땭�~�'���Y�r^xL#ƶ�fks�0�u��~+�Ő�4��P]=[J��<�S��Lu��Y������}�7B��`'#ג��G���а��:orۼ:61�$�9d�{#�<X|5cqu�VUZ �W3t��~R���v��ky	��.�9{��;����a��ja'�-B�ob|��󚜑������}_|�̷으��J-���c�(ASD��(��,�ߊd����#�jw[�U�}�N�&�ekXaA�}����{����5\9�I|~���}E\N�x�&ha�F�9�\k���ze�>O06C���K���GD`��YY��x�T&�����x���q9j���m����6�\Щ�/�
����87��53*z����]�ݭ��#���N]�s�`��}�\^7Y� ;c���P�0eB��t��1�u�rpX7��lp�����VI]�^�;��vG�0,O#5A^��]n�(;�f�fUJC��C�8S^�U��
����m�;i�T^f������|CG�e$�z=lQuK_p2�	��n��က�i�߳�Ș��w��FVTg1�A�_EV5 �"�z�0����ϬQ��*x\Bx���Q/_�-�����8�򃚈T�_�����\�<pxu���)�wf��&���]J��k8��a����x�cx�kLV3*����wᡸ�4eL��eL��WB�5B�aq0�$ط0h��*��M޹y�ܾ}ڹcq�2�>J0IN����]^2z������D"�i���*��L���{rf�Ѩ��j�����-�;I�b��v�x��|��;y0ӴU��|}���"d���ы�C�/�i��S_g7�������of@��
_ĺ�y�e��6Yd!�]7�{�<�El��`�#�E���v�k���2������Z��o��(=Ŭ� ��srB�T�x.�����]���&6�Z��^��ۺ3-!��$h��<".�˃�0��[�|nۘ	(N�B����x`o{E�/M���A�-A�g����p�W +�n�[��K�K����=�^���Sk�-��=�5�ډ��_���^3���f��m����QU�hCW�J�Ą�Wȏ�r���==���'���Q|�eV��Ԫ��1v�u�:75�oI�嗧+Gp�瓜�;�¬&ٕ+Q�Y��*v-��«k>q��d�]�>���o�ā�=�w�{7��W��{�2�VZ��8$��f����õ�2����)Cn�Y<sѲBo=����[c��P.��j�;e�ܦJ΁1�R�0�(8W�5;%�.�y/yQ�Q|�޾��<{�f��aA`�F����U$�OU_O o�� �h	����]v�g���p�]��Q>t�ڔ������,���]͞­�*C@�/&0{6��b�:S�T`����[�d�k���>ǽm�.B�sn�Ք�J��aܗ����&�wD�FE��s�`L���
nm;�L���(��)߾����6ed��;��_?eC}�	��N.��]%CHK��:�~�W�]�K�2�K��f�zgtŁo�TAim����ic����tP��'Ib���1���1���=��y]�m)�j�7Yn)���)C�"�cӓ�U�=�,K�*�]z"=�
�^�h^4�O�N�m�*�;�ō�c�u�ڜ^�spk�!�9���z,㞞N�����鮸Y�y�w	������U��|��3aA�>��5�#`�
�~��-m�X�n�%��2�zL<v�&8]?R����",�`�G(S�Tk��}Ƙ0��'2��4�}&��=�kÆ݌��Vpq�ĝg��IU�":̥墓������=��b+Gey�ټ%�o3� ��Iu*U뙌V	,����ă��G��
�z���>HS��.w��X�������o�8�}�-u�xtX��|�[ z����HL�|CFs�B����q���]��������,x�ډ򂮼�24z�gڬS���Vu���/->�h6!�^����:+�TR[|���X8���(�����ak��U���m�9�����2�=*hr�{�^'���ʘv�f3��+UL����]��?a���5�I�<W����s[��1v�+]'�?W��)/gd\�՜��TX:%�d�/���K풼1�f��ßC��8�+����c����fb�؝�X������,�|���I:�Wآ��b�<�ЃA&'��޴pE���W��ҍ�9/{}}�۬�
�P�k�%a��8\�ٴ��4��|�M���sqv�i�Z�łz�OO�"W��9	��¨me9e���c�[����Y��]�t�w��'�)8O�X����S(5�t>qs.T̵�/�ՉY�����j�J������^�X�\�":4�{K�Ϫ���4:� ޮ������h#_���6{ݗ��,z�����\ ��=�)E���Ƀ�������{zR��nڈ1Уy�����bN��7|�bWX@*�"� �����Z��ߦ��Ń8�/c��+2�.��}ĝ�Ε�2̧��ŀ<��^�C�"���J��g,B��(< ��M�F���Fױ9��>�L���׃��b���<jĳ,���&�٦J�SWr���5�C�+�Q
���GxL�|4ebq�	ž�5~����c�KҸ�I�@�]r{�������=ꌻi�)����v�S�0ur����S�لG��q�Gu��fF6����F��&���z�Ǜ�ev��%ӷ���9E;�}U�Q��'�۳;h [�sG�g��P�ln9B�e�UN�SC�E����go�R�˯*/Nvۢ�T��-�K�+�2�^�G���x*+dT�=#Ơ��������쾤�v�,�qy,�C��/�*ˬ��!��=����7�>j
5��b�����@�7�T���QzaX��m�Wz+�<Hq��Z`�9׵E?���E}�N>�������G`����I�	�g�V�L~�0����>+�Þ9N��nd����(�ԁ�/�ۀ��aX��O��C}�2_����m�rԡ�ӤԳ�e�M`>Rآ�=�&�-ݩ���e�K��"T��l��ĉ!^�F��=$]��0���#
,�Y�
��OJ�l�t֐�}i�SixmVx�HN|7��Lʁ��G"�>���FG�!������s8�Y�.Ϭ�!|]�W״��P��*�:�4�^���:�պg�w�k1v�����9K�F��	h�H��V�UѺ��&�Ƅ3vXX�y��Y�`����)N�lR�ڼ�:̣��C�}���+Llwvc���{�9�F�����06���C1�j���)p�AEb�`Z�����t����o:�3��RW�l<��jsCy�,�:�n��9cs;�T����d�Ջ"�����U��׿���p-dW��/+�5���C8��G猤�G��/孰|�3M�u6��e�-,�����s�
��R�U�_4��z�?��â�us̨JaS���М�kl餅{��b
�pv{ݦ�yo�
��`W]}͚��Z�øo�ul*r��r�[�J��+r��=�+Y�R^��� ������%��~�	B��
�r��M���o���N�,�<�%+���p��f��鼣=���@�����%�*:�f{۾]���D�X vz���-H:��srC�9uf��t�qzyB]��nLU��{��͍��fd�՜ꭍ���#����G�����>����n]z#]�o�P7�'{����R�w{·���j�O7�*�ѳ� SÃ��G��.�,s�����	��"u���Į�'�7�c�l���>f�75JxN���!c={悞�蘒q�Mo7,Ҩ���ћz爿�V>�@2g? )����;�njN�!�r����޺��X;��+uo��']`���PA�ed��B�5b\(2����h��eX*W`��-��V���ۛ�kZz��sw e�S�ڻ��Վ��ѝf���[B|w�;���L�mb�x�7�}w��&���JA�2����w[�����������Wj���He��\5Cת	S����q���V��f�1ڧx*�3�{0��j{p'S�C��4��%�pI����a��u1�0�{�2���hZ6t��e*ot�e�r
�S���`����Ic>�z�(�_c ���r�E��w<^�$�=���o�vdo]�+2�0�'Ǳ,����O�� \��N���]#��Wg����+��s�O��g��]Fi3]�%CJ'	t�nS�7��.	L����65#x��X�����ʦ��V�}���3�8��x*�Eh�t+���ٖ0q��35l�*�t�,_W,ja��n)��\��ɝY��'�g5��K2�K��}�OX�>�:?o�<E}��	���Ŏ��]cw4�spk��!����'o��`&y�{��-��u#M�S�����1���" B�v�4������� �/�o���i�PƢL��Q������M��`G�w+�L)OB�M�PW#b�7�n�o-|"��ݵ*�o���҉���ڂ�S�h�;{��M��,�4�εY�7������[����^IXa�p�*���GWN��ͤ鹦�����#f�r�HWc�	�{�s��������||���b��]�y^=D�c��>{|��7�r�aQ��wy�~�SHz��,3u+�vѾ�W���2���N�>ҏ�����c�f{P��Ļ3�Vkr��"K�R�ĸTd��S��O-u�C�K���Sl��D�s�A~�Cj�^{�+~���變\ʣe���[ {��UN��ß�ζ�_w�㗭Vi�:;�������!�����>E���}pU��ǆ�E���$�[�	��C�S�#B}��g��pƼ�\�|(��Mz�9�z��/	���,��b6L��z����O�PkVL���ګ�Zp�.����Y�u��(�g�J
�;t ��&�����m�<��������y���\���1�Cx/���D�?��� ������+j���٧�8G��`p��������X�J�]bf6�����Ԯ��b�Y���c]k#YB}}J2G��JB}Y,
U]'z�2��|���^�(Κ�I�2Ҳ0���`��>�,�l9�ra��.�(y��7�2�,�k7Y��������|,����ݫ��C<��&g�S��CyO}��Of�M�(��YD��V��՗z��j�0���{�R��X]�솏u�-O0]��#A`Y�e���������%���%�Ўf��j�����cL��&.�^�Y��JT��L�5��R]%��>/1_0�a��:��7���XG5��$�X$���cc��BVR�{`�xzo_hj�����1�SÙ�M�2������"q�Ã�.<ohlo�3-=G����d<D�w��;��kw;Oy�z8��������Υ[Ѵ�|�'_oѷ��J���O;3*�.sNw'�z��F��I��wN~9l
 �y�����kJ���7�������V-I�T�`��c��Xޖ��q�j;|V���A��Vv�1wac�/݃�Y���i��1R�S�ʶ��Iխ�QѢ ����D]�k$���G���o�����)���ԨE�MvvѼ-��H��� م-�س4b���=�0f#�W`�ޯ�wz��<�׃V&u
y��Ս���5�W
w�3��ʹ���
n{�}����j�1ԋ�c*��ż�!+7�|��;��Z�;Ȥp���X<$3ڄ�����V�*J]@�&��y��ż%��H��8�r�5�B%j���<�zί�w]�]p�	Ӝ5����d=��]v]ڐ�خ�j�Rn�tDt�O�$���ה�ʰ7L���a��ڼΰR��n�U�7en�3�O,��TN�ROk���b�ifm�lbQ�u�3�5܎sV^p�c�:.3���]\�Tl�����]���;�U����rɑ���f��O�kܲ�f�����]{h~N$��=۾0��[�����Zg����\��� t^IM;�I���;c]6�:e�D�#��l��-bT�1�ӧ!PBةx.�d\캉�q�Q�����b�JopZ�Ev�В�}��շA�u7b�Wf�[�0;@ST�I�2���[�V'lY����u<"\�z2�Sy�Cm�j@��ɖ'��7�=y{Ce��S��.�8f��۵ۛl**�`Ǭ:Σ�0E���qȹ��$��՗Yr�S5�1�;�O�k���Mv%��wVG�wi����:��8�h�9�n��a �4�.�o=z&od����qy;v��\6��Y�G\	�<͙V�ớ��|#ӗz��.�|��QڍrT]ƻP���AGۉa��Ek���m��z�s�՛��{r3�� �kY���iNL�x}ՠ�|>�[wp<��u0�m^k剪G|'��<�x.1�uV��Ž_�q���%�Wt�0NL�0��T����s@��k�A���c+t�x/��
R;/��[�*��wǗ[%c\F�=j�g���˾�|�po����b=Nk�m�V:#�ol�ocP{�t%��$�OGo��=��Wr�/_Ko�^ݖ�e�z��*�Y�?�T�8¦8̖Ř�RT�9H�j��G,��ڔ��W�h�*Y=nJ4���B�����fLZT�4F,q*"�*X�h(����n�T�RV	h����(���e�Ym@Ql�s0�E�c����Z�B���(��!fR����e����1m�0v�f�fSW2�PD���)[�jE��R�V�m+nkX	�բԨe�Z�ź��٦���n��f2䩑1�Tk�3
ڥ"��5��T��\�kT��i&��[X��W2�]V�G)kJ�"&e���e3
��(�p̸�$Qm�*V��+�V6ʴs
�D�eeLLJ9pµ�f�t3n�L�J�����m����S\�F��*Yn��Ĩ7I���J"¢��l�aP��LIc,T�����a���6+LHX�@X��.Z�QG3܎mTL���b����A�A���*��6�;h��+R��E�V��1Q�n-2㔴�Qm(i����WY��� T��MQU~!q�Փ�ڕ<�Ĳ&k�ޭ�2P�N����6�i�)��%��0s�����N���a�	�Q�&���؏a����Uk^nog����]�f���W OP�hs7����?	�u=�BB��]vL�%]���G6C�^�'5+2y�@EWUc�0��X��Ѯo%O~M�i�{�*�$�ݮ��|Gi�:wo)�����#��1d��>~�<�*�;0�.�FH�C�o���ջ�[���ϙ��=>��H}s���x\1�}2��xXn�'�!�ɨ��O�=uΞ�����h��� a�=�Â�=�r�TI�{�*��Reб�B�]��0����X*Z5��{2g��;x�:z��Ƴ�@�ӭ�d!��+��zG���ՒȀ��2c�s=�ܨmOeU��u���(��xV��&W��vu�.x�<�
5*S��Ez0x>�y2s)��yEB}k:���D5��+��xL.�ν����E��/�� k��$�4%��:�.��Hh����V����0�J���*�%�~���^�5ѳ���k����e��间nU���'�3�fx�/N�R�ٖ��`�W��^(����ƅͫcƕ��x�yt�5\�L���^WqP8��|/&�ct_1v9��F#�|N�|�cJT��\�.;�X��ģ!'��I ��ƶ�.�Hb��\��Gc�Unc��1��Z3��䠭��\r��Ɏ�zK���٨�_��S_�bu0���GDg�����}^A�0��Y7�C٭��@��s��^�J��7`��
�u8K��Ϛ��</��k��-Y/˩�!�����}"�Y����]A��2kl� ]�*���}MBw�t��՗LF��1W��X����n�hJ׷���;�+ŵ�/�����jN� �
Ų���a�u�4!����ARer�^��$m���!i<>�8�jN
��=�44:�"��!�I�筊.���|�R�G�v`�jy����3�a��
������8�����m�6h/�QO�tw�Txyz'���;�������l�?��[��l�,q��o�71��+�6h*ä��"ߦ��#5��/�:�a�RѮs�>��k9T����z�qxhɓ���s�	B����l��s�vkfW�^f�ƥ
��^��8ŉ:�u�.6Yd.�Sb]����@�����z]Ћ{�p���č^��k����>s��Ռ�R2���]/���9ު9�=WrKˋlC��4}�9�>~x���Z�t��G�J����}�T������b�q�g^�.g��9��Sw��F���Ue'>=V��w�"��R�w��)�o:&�������dp��C�vϮ�tэ�׫��4���;�b0�|����R�\�1x����םn�du=v ��!�ʤxDv7��<�R���V�5�R�Mo2s����ם��7�д�c�9t��w+i}1)Y�~��q�N���rؙ�|lo=Z�����V��r.��誓���p�����9���|�vM��Uf�j�*�˜���$�M֑���T-e�2���,��9V�o���j *K]��|����Mv�̮L�Q�g��M�.���~�{N��|8m�2�A)�]����?�ȫp炳����+��=z�2%߭<��w]�J�+-A��X+���7��4����z�n(�����Li��qh|}^������^��	��c3>��U`-�3��+8�0��9]�N��xI4�[ǖ��;xtFk5�����e����\r�%������51ⶼd���S���l@F��Г�Jg�<
��B��]%CHL�8�:��s~�����ܭ���ˮBG�*�ryz-�U��ӂ�r¬e
���,˻�䗶\V��X���d�9@9y�1܍�d���p�����,�n��v"�}6,�N�/��8e�ڷ��!Q&�b�v���k+�Z-�M�Ib��:�ǵ��`��m]���ܲkg<Lb���X�ū*�8�k�c��{0���*?p򺘉l��;m�k�~��SW��>�x��� �fK��������g���M\ʯ|'���yW2`�v��\~]���%�&�J�<*��^}b�L���F6���\���u����(�;�mqQ�p��g��}��I]l^� �� �`�tiV���Py��mD5��X<�f�'*L�-[S��Uxy�g:(8\�(.x"�"ɴ��P��T�� {8���u���پu��,{M1�T���Q*�p�}N��z]�3��IR"(�R�=�7�*�v1�o����9������z��t6DEefa��~��i��s���d{�t̻�U��l�*���b��C��h�s���dq0��3�4�y��2=�fӬ���~��۞�(�KO�iOh���G��\��AWHyǆ����滗������'^E��L?z���L�oG]%xd�.���O�К��g8�Rgi�Kuf�INI�N���*n����ϱ�ݪ�h�dԑ�_��p�\~~���L���f�bg��&wQ�����Mw�E��{��wnMP��X��ʩϞ`Of.�I8,���;�)[��N?�R>��o+���6�G�c�}������8^mު�4c/
��P�)���'��ٗ4�B��"�׵^s��ϻ�� <w��ijc�o�wc�53��]d�+|xf��(:�>-�qr�a�6��p�ޞCo8�]{U;E�5�z!*�z[����@�!����L��W�6��=���[.�]ѵ�o�Q9[X���5�yҐ�d��Iީ�ʏW�-��PV|�'y�OI�s}�D�*�R6�B͍x�K�.�+�\��Tc"���@��*�7���j1��j$k��&��Al�z'\4�bfl�&�ѝC�9tjR���Z[ޤ:��)N&�#���E�P*4k���U�從����Q!�7\�����g��muF_�n5���z�Y3a��t�ydU�	%�gE��*�PdVy,d��w���t���P�2�S׃��K��
�L����x�s&�(�W
^�ڱ�<J���o�u&:�ӮC���5���C-[��u� ʺ�t��Y��Rg �rלqbsI5�°�����k��r��������@�����{3�e�v���W|�^?õ66��:W)C��r�����㠍S����d6���web�+Ǎd��+��M�qna�p��Wϑ$�;�jr�仒T>̭ۜ=�^ytjN5%�RXW*�8��閻��U-}l��]���|}�o��B�?�W:�]e�</��o����ts�C3z`����F����1�_U�_ s�:�C���3�R�!��V��zS\/���9~s��ξ�5��
J�u�ޫ�>aF���� ��֜�m!��V
���&u�px�:b�'�bQޜw͢���]'��+6^�] Cp9��C����|���v����,���v�K��I���b�og����J��G�E�b'����IiU��j�?EC���};1�3d�0RW��W���JC	�\''v$j�z��*���O�ҡw�2y㵞������,�9f��CJ���P��)^`ʅ�A�M)�V^g{����R����cc1;��F�k�c�z��gB�y$!�W�c����'q�}�
����_,���y����v����ӂ��wZ5�.GQd]�C�v"�^�@������{&�}Ӯ6w��`cн9� ���������LWK
���ćY�<7�՛9��-q�j��p!�=�������݋���+kND%f��i�9��^�z��[�6���a}���swΓx�PK���#��,ꜫ�m�v<մ�{�k�xU�[��M$�N��@���o��p��<|�Z��i�zu�[E���'Oi�����������}K�ofUB#K��ފ��d�U{1ub8)�Ej����}�}Y�o���Z�m�'*{]�/�!����j�5�}eV�����w�۵^^&Y^[��a�m_��:��2�
��8,�<K���,�>,�H�~����)�gjv�Sݷ��*��M�}:��dz�hǱ�H �Q�mf_��n�8�>�l~�0�X���ؽ���ul���~4�R�*@�چ���EV�G���c���K����ǯ�Z��0�7�$�`����+�gY��ىJ��g�g]P�*�ٟ}J�ݶ'�A���D���WSE���y�`}t���ۃ��n)����c.�r�^eځ�to��9�~j+4v3pZ�k/Y�ý��u����^fUP�1v��;��
��9�+p�����{�ˮ�ը�#l�^u�Ğ�CF3��=��A�ŵ0
���d�Y)��ܡ�g����<���[T�9}f�Ϳ�H�Q��o١.:��ۉ�����>B�漦餐<skN����%�S�$�g&_C�P��p4[���Z�غ��J<��|�,�L�U��~�.4���tbO�Uo�ܷ6q�ڕuf+j|c�s��ё�A(m�4�a�^��<��X�l�bΫ���p�2^C1����~��o���m�y���+�g�i�����y��R���S'lͻ�Ual/���+X;�h7��<sY����%і��,��c�p{���Df�_�t�m��t���-ϾIp�7�z|�o3�]�k@��p��Ȅ6$�R����u8��\M:N{}��8H�v�f�@�`~�E`���ʼ��&�e��z]T@d��K�K�	���aV�|;�4;+�W{��=�V+ O�J'8�x=�u�=�r朣3}t���4|�p�Ｇf��@'�}*�̗*N�Y�o�4)� �/*�!��|1�4�7��S7��x6�/�:o1ȧ��u�>�T ���� h��4����l7O����;���~�k�����t��v�+��^.g$Pp��P_���E�i}���h�(�>�����KV�+����s*�O��sXu)9���c�H�2��0�}"!�畍�����\�6�P�z��h�KS��"JfT��LVIf��&g�\��˲�VK>w8jI�X����w6��%���;�e���o#*U�*�B>��{y�^�!'wO��B��S,S�Z��$�ɸ�\Fz䮾��WQ߳q��󩍉e�4�$�����6p�o���޻�_V��_E-��v�x�}����[��(�?+h�;:��n��f*��d>ޖ���� l�����˗R��]���MD;>�si�kBƦ;��mV�
ߊ{FL�#ʇ[��|���͊�MP̼�>��c�oH��p���u�E�ڕ��zu�F�>��7-�!�Y��ڽto=�c�&���\e3�FsL���lwj��/��0��]��v�ICR�XiyΕ����g�L����T;�`ԃ�>L��2Hd�Wiћ�m*��k�r�7Ӽ臝�:cL�N���ʌչT���k<ЕT��������z| �\��+�pxo�ǾP�+D�Fz./�#h{qϮ��a���[�ט2�����eG���[�|}��n}1t��[�&�J:p��V��ֶ�#�Xd�:PM͞_ޗZ�g�����`{���
g�����9��=��2y���W�0U�N�h���0Y�v��&r�s+�Ṏ'1vz��������ߩ?.�X�a��Y.��2a@ׂ�Ѭ/�.��]E,wE{R(�q�N��W�e/=���<�"�u��w=Ԯ����{-�[�im=�����͕[�*fԀ�PT0�J��-��9�M`�8�s�q�in�EՋت:Y��f�AY�]ٲw@�c3h�:�馾ɫ��E���|��ROZ�pg�v+�~c����+B��=C}3a��n�ydW2a$���	�}~�.�޺�e��ן����g�R�?_�qJ�LW���^.�U�L��'���x���de����M���{�XL�k�ܮ�r�γZ�Sg��"�)��lvQ��l�\E,(�jѾ�����|7j�fz�4�\.�l;�r�4�U6���n�%ѐ��B+d��W��5H́T��k��w���O���E1�����C�r�����y�+ުޞ�{�9){;���`��C�΋�r�xc,!K�!��hzף\/����%mL��~�c�~���7�����L���seL.��)[Hnj��VP�@m�ּ'�5*<�x�F��n-W묩��%=�
͗���%��c<'��e�}Zt�j�y�n�������K�"ŵ���|D��jC^�E�P��tG����>����k�W[�e���[��l�hz����#+��)��̥��%��fG�ӷ�ٯvTB�}�{�#f�2�5O_}��M�=�D�kdwM�8���ƫ'h<��Vm��.��Y����6$��SɎb��WC��F��D�ә(mGO���r���������� t�?slu��s�7J��քLԓ-2�v�.��M�G�w�r�N��޽]�*P��)������M��� �F�����T(�\5 �06�W��V�����˝���^���R84�jUT�a<�w����������h�*���a��셏����7�pP,mR�(��lM�[$����=d\{�#�/U
�{��Ym��(ˠ�{9��8��t�~X:��>��D ������I�;c_iEu��3Q�)@i1]c�i�6�l�V5�8e��Tm�o(Ą�X�t�n�]��ȴ���K�Sƅ�������g�����[˱g}lQ�j�����ё�tǶ�mYM!|+
�I�y�ׂn�r�q���j����>*�ܛM��u��U�������!i�Ue � ���L�OH�@�����ë5��:�)�(v��1�o:��MM����-�X��t]�)��n�E؁p���F��y��/n�ٯ�<�:9>1�>�٥w� D0�����=��GZ� ��j�s�r����<����O�(oo1���j�8=�6u9�V�t�Z-T9���bJ�	�*oTi��8HB�1�ާ�e���8�=�Zd��e��)������v�s�<�6�>|}�sU����ֵ����W;u�D_vҢ�-��0�xq���K웾���N������n����Z/hPS�U 11S!!�S�q���IC{�a�V0�v�N�E�(a�s���H���F7)7I�`�R�̩"9��j��X���"���1kR�e���3p��L��4�Ǻ��E=+^�f�e�!��lr�Tp����tst�:ds]4�]��iM��7+���ӓ���a��i����Oz��!t�-�z7��ɜ�K�p��F���oI��: q�<�,�ُhs�r�\���"��5��3WG� Q�/��"��w�����U7T=�,�_�im� ��6�=��x]O4z�59��
.���&bZ��醮��`�[�"�oF�Tz��G��ӳ��쁭���B��Z[��퇏�+��!r}�����Ҷ�g����7]��f7�`�q�odz��N��C���=��崙�O��r�Yεϴ�[�^q3)����
��7
�iһ�κ �:�Y�,h��y�qc{{�j@��LR�v��q�8].9-�F�wep��6�>�WKaa1.�uf.�,��S7���'���VQ�+',_�sN�����u+i�Z�T�ȑ�JP�T�=��M�:��ɯ����	SY.Gorhy�)}S9]��/�Y,2��f�k|�O=��x��D�(
�A�j����"�unbL�l��]k0��ɂ��Fچ�1��aJ"&%>�f*[��3�˴���#q�P���TI\K��hfWX.#[[�ܨ��Z̉��(�G2�\�+�1�4��Y*V��j.�\st12��S-TVaTR\)V��r��V�*���7w&�0���ۍph��
�8nfq�Ӊ�a�1)�+c�`�8�s�֖�+SVɖ�ieժ8�6��4���.�����X�LAr�+j�Qՙ��(�e-mR��jl�"e�T��j�k�uk�D�SWFZY+T�+���-�3)X�*"Ya`��%�3.j㢖Dj��TE*
2�E�Ji������j6�T�J:�S�UR�(5�-�CuK��&V��1�i�Tk-V�j�YF�c���kJV�V�2���)p�FbM�G,v��ܵd�U�V��հZ�R�Z�Z�(�KZ�Vm+"ȹM�X(�*Tm�d\-0]�2�ʶ���E��TR���KMd���Y���)F�UH�[mES2�(T4��F�C1���m��fۦ��[,��0][�v�.ڮ�W+�˓02�U+��R���������o�5�n?Q7���l���}�xY����S��t���餔wL[`#/�9���2��I�p7��9}N��'��Z���E�k���P�k�����B���b�C�Pu:h��h��VB����<�Q~����2W[ᲔdhuG���I4U`���h1/�e��r~���(�=dk�����S�����_22uX�Ϧ`�_<C8��񔒯^�m����bg3�<)3�	�� �X����'�����A�QU�M#W�f��k-h��b�9���#��]N�T����Nm�Hz���=Je�H�J�S4+�Z��vޠ�Hi:�o۾��#B����*LK�[FMPV2a��9��ܼ��	�ՙ�E���ndq�r�(t��(P#Ү��<K���r�z؋5�*lK��|�^�Z�+�<�T~��>�Ǵ�xD��h
��ۨ�,�1bA��ꐸi�7��/�(���y��jwԄ��y�t�c�@�چ����<�C�G��,^��׽�Q��(��o'Y��%�([�p��L�r��ĥ`~��0���{YO���l|6�ɣ�A���(���X�$)�r�>PK�u�_%y��q�묺�^��]��d�g<�������=DAf�ޛ%l�N���x6�<��]85��(��6��H�N}��V7�*58��^������0v��2�)_C��l]߾��NN���
w��5z���L�N#l�`oET�@��$C�]H�Γ�q�v�
O�ٗK��y�,�$���Rb�L��]�;�n)����Z%���
�=}��;��H3�^��y\y�ػ��D	��ӽ��_����%gz�O�
�O�T�
18i��kw�;J��˧X3c�^�U��'\*e%�3�||:���>�|wb�����v�!ܾ�E�IpV�*���]�Xd�3R��,<zvp'����%ͷ�XC½����8Pj)\e�>�����U��F�[&��݋�<z��9#]kK��� 怐VD!�'*��->���Pzk]%C���U�1<����t��e�v6�g˦e^mHH�jx�%���l��'��/��k�Otw˞2�*�P� !.���a<����g��|�=�`ɷ̪�-@;V������N��i�F?"H�[A��	�3��:�cw<[��5�G�/�̆��[e����GVX[]��
t��hgG�s
���v�����f߫�j��= <�����g������(so�g�K��mI�ⷖ.����KR�Y���CZ{�r�mӬs�z^*����N1g{��mr�w��?��s��R��O����g3;��I^���@�UZ@ Ь�ҭ�/�+�0�EW��[��.����ݵ�(��yB*�>qOϢ���0e}<�y%�_a<+�Ѻ�lz�I�/}�G齺�Xu)�|*$=N����ck�u�q��
|�L��Jg��]�>Z�RuK!����c�	��I�`�ĝ��-����`�rC��y�5|���^7�Ӯ��
!���*�/f*��d;� {�s���dz��2�R��}�6y������A��sjC������->�=�g��R�Rq=�#]�|�]�|0�O������{	��1G\&X��֕���Nr�}�%o�F��+x�L�{Q�>Mc,A1g>fV���&N���E�V��i}">=�).I�k���+r9-%�ySu&+=-Ѓ>ԃ���|d,]zK���b���L*��i>�N�-���0[>���q� ���|��VC� E�xS��%m��d�y�jM�yw���e��$�0�<7^���~30;Zg%�KJ��&Ŧ�v��ݮ�*��x��*�6��'LHw<�:���m��2�kT���	��/�#��B���v��7����{4+�AQ�uߴ������__Ft���-�[��˃�+]'��}�(ߟ��oI����|P��a;Or�k��Mg��	�K�WIީ�ʏW��N�܄Us���fh��>�-F��C�0V��H�فnJ4��钼�ʛ�*�Uy���,�-8��o�wl{��}�um��f����A�����M�٘/>���}�̹�ͥ�r}������{�|i�~�=<��c��꩖G��Ʉe%X ���&���u�?�7�͎r�ȝ��/�M>߫�>��B��y�}=r�(��w��t�"��	�}�;�I�E3�����o7��������S����R��}s�ԫá˘B�.a�~#�;��o�h��=�{暟vٯau��r� x��f���=})O�TI�W���N��;)?���=õMv+Ԩ���I�_R�TX���9�:������	�fI��o��m��Qv@�h[�J?CZ��� �]WR���u�B���C���=�T2�>�|5��c�;�S�,ϻ���]1H8-�8/Of���^Ƹ^W��r�K��uHQ��i����K�����ǯ���p�K9��6�;�F��L^��Y�^��u7��ms�-�C0g7{è�W7Y�/-��tܸ�lu�Do�L�{��/�.�.�=��s����m�Vw��# �a�T���Y��nm��_9��2sU/�K�{��?q'@���1�W��k���&?	B
�Y,O+;��|�n{{3͕�a���h�}���	��墯��Kȱ�S��J���[k�7�9�K�c$z���9Qb��ڶk�Hjv!q*��tG���ڬ�R�.�E�I�<�� E��wXx�������J�S�=N���=��
��]1o��`����p��dA'&��6�nx�JL�Y�!cI��C˄R�1r���[��u����Zwvx.ooS��.���c<xN��nҌ��^�!�`����}�ʜ������j}�X�f�!~�`@�ip�/�'U���j����!G��G����Mwp ͼ��Yˤm!F's��ud3O�]U����N��)A}U��"V�YI��O7�a�@��&�T\Ҧ]��g��sojCԲs�R�N�+�>I�7�;Z���ڡ�bDVT'k���x�u�N̛r��wzX��&,1=��M��:��6�o{��q�<�q�W"��0^�����Żg��:l� 5�Ob��:Wu>8=;lΚ���,yz��z�"n��w��x2j�zM*�ꇷ��F]G������hlrS�]$L�s�1�?�}t{���lS��Wʽɠ{��j�6YH~Ш��
�'ԏCı�^��9[f���+e�7n-��^�V�ッ�A��� ���o���ݮ��{��<-��p\6D�R��RzoOR"�4�K�=R�׾�~����t>�W��4��u]��˱X�:k~�"��xls���wOQ&�PR_9��g�]3��V���02||��m��259�]�P���[aD�=�`�kQ��K�J�R*���q�C��*�^a�8߶�;Z��C)1Z;*\LQN?x�ͽs���X<������ګ�N���M=ɧ��XV��2=H��F�䯍p�`��\�v-���c��~�h[�;p�&�e��̉ƮO}�"&`Lt����V_�:�N�S{B���;�G��s���-�rc̷kO���ь���$�+-ۨt�p;*��|O��U˧cE]�Id��k�`�����0���V���� �j�Ho���`��W^�vo�f+y��D#'�p�	�+3V��oM���M-Hq���3�"K��yu+�q��{~FT�Ǝ*�z�7��홝ԳT��f�|4NQ�J�w�z��S�urj�jѠ�m�^*}oc�B�雙��s��7�9ds�����A�}����۲I�����.�� ]y�$ՑjNU+����k��`���J��ثQNg�L������Ҟ�@�˟�H��S�"_��b�諙�fpM��ӽr����U��Ίa�� 5��𤋮���e����({��SX#��ʰ��j��8�inv�I�ȩٖH���4)P�N��e*U���]`����7���l��1E������{��C�n?yW��O�<'��ʙ`AuS�̐��\
4ዐ�{+6�񺗱ƒ���к�/-����?
���#���J`�HL�5rYd�`��eꊓ�s��ZF�ٔ:�+�p|���t,�0?THz�ˤ|�^tr���ᒪ�A:�sqbX�3��Fa�i�GS;�a��͇�,�l��n����F]n�o ��7������ăܲL��g��Qo�:Ў�����{r����s̭WRk���Β� �*�R��Ō���u=�a
������ZS�<8���,�����S�{�īc�]�٭����R�L^�h��d�nky�ׄ�!{%�?{��=�C�C�r�w�.���;{j�x��gq�K�U�;��$��iݺZ���5�R�b�v�N3gW!) �����55�m��׷_�Q#��������C.f>7G���
�C��>񃰙Z�*ժ��"���W��{�Ep���-�@|����Z��<6��˼]m��`�0Lr�>ɖ�v���h@u��`���lNub�	,���(����R'/m����+�r�3R���7�B��.V��uÔ��rQۆb�����֓�l�8�[��!�� �����;�r���囓.����;�wz�3h�+E&n��^\]Ee�*�p��;��K����qSz5�Xi��L����*@��}2�v�x�ՇHP�-66^�(֌.�+�\�������z}�L���VM����sBB�[��um�e��5ԁڸ)����[3��N�s��Ԕ;f8ċ�S��T��+K��k0��FϺ20r	��� pp����L������������r�K����#��1d���ZՑU�J�$��=ݭ���3����&��Y�WJ,9��)pk&Z�a�xg�zb}�
 ���ͺ���o��0}钂��fO?"3���h�9V�б�b��Q:�ޣ�Y�^��/1L4��٘��Q^�mI"�8��nJ�y�V��]�%ֽ�V��]�`k�U���]4'�{yr�7�
���[�§��(�2�꜖����^nx�ru{C��DU�K4�_[�M`JW!�@�y�t"B�b,R��D�qb&����i����#A��Z6�P�xR�Ti�vI�M���k�����i���~^��d{o��N]�0dh%�����8���j�@�6�=�1�)��=����+���5u�;�	i��ヮb���K��wC�w`���3u��b�zO/>,!���<Cֲ5��v�d�Y�k���}�Y����@糈�=����!hy�b�
�]i��V���eeiw�I��#�~�I=ibr�c8���ڢ�=~E��U��[�մ�.�d��"�x���Ge��uy�(q�L�)�X}�	�:?]��yX��ܜ%���#���k�u߻ٗI���X�2$VsOh���׎w6�����>��8C��pY�	�x��ԇ=��1Y���:��پZ�R���*Vov��:�W��A�	�`�>����Y�L=�P೨�dq���R��(A��
x�O������Ι�46���8�fX����/'\U�ꭣ*�2}f�P��'���pd����M�����Ws����m�kF���o�z�Ԅ�h�Ѱ����	���[Y-u`9y&t���g��±���S��BK�[\BE��5�O�d��\�	�Vu�ݢ��N���n��U���GM���ҥ�{��)���˙9�v���?�Z7�a�d�]38�l�o�{B��^����hg�9,��`�\z�<p�$�>�v(��lW��C4�����f��ۜ.�����G��8U���&�gL-��u3�U{m�3��9���=Y9���^[8"�'�I��FNo}S��-#����CO�#��]M�N�ɪ
�L���I�h>˃z1y������~|=2���m�Y�ԡO���[�A5��U�g�X�\������Y���p@}���z�g[Lk���S�}\!��}u=`1b�~m�E��� ����}���3w��ţ�� �ugI��/!�zd�u���j�=���T��]�t�˺N�y�F��3n��'۾�I�
Z�c�˦tc�[JbR���b��GRe��_�����@���1=9�9w��{�X�eoK�y�Z �HS>'�t�%X�����ݑjhy�e�>C*�����K�I��-����8��U`�����z��o�{<� d��� �!4��Y�f�wK)�U"�b�s8�e	u�1PR��Ӗ��N���]�&{����niCs,a��վ;z��|��/>/�G��D�ml��If/���+�|��y����n�KC(�h�勜pbl���o+Y{��]��w�� `�cnpW�s�hh�E7Y�2Ŕe^�x�3�]�t��p{<�U_OW��3��Z/ą���i��6��:�9�\�0˭��8NkH��)�=1B�bF{��$��[��l��u�ʔ+�^���z������eE�g (p+,ldP����o*0k[qb� _[��,����q��v8:��1�=I����냈F��_;W��w�7�Gs�3KY��'���\؇:`:g[Ш��:�=��_�f�G�xS�����۔��J}e���G1��;\��ؗk�I�:�l�rE7��\��p@�W9�ۆ�EK�֕m[p��ҭ!�t%���\r8����8�o>�X��
(�Or<��p�Ӥ�kV�1nؑv��`�Z Ravc���%�R�[=L*���2��j�7�`A}6��˰���8�n��۾������'��-��׌��������x��n@�L�K'�ݛ�켽��Rn���Χ{�`�2s�H�5�+4dҧ�P����S�6/�u0+����|�zӻ7�ݰB��>�W=�ԍ�ݸ����oQ�\���G���b�ijz������Jg��i�q���ԧ�y�Ew��m�XwT��%��+y�\W̈́����xr�ț����1h�:��Zu��6g".*�dV23�MЖ�dV��kw+Rz�*�r�p�ڢ�<D�F�Y���L�R'Bz�D��GQs_%�G�	t�᫵��WZ����h�9G.��>��(dr���yy�L�2� �J���x��_��l�z7�]��k+O<���Sכ�e��XG�µ�-{��5���H1�;�����K,G������8�oljFȂ}vw��A0�&vnS�-�5�˴���c��,*�A�g��yQ��O�]I��F։���S�ڭ�x��>��v-�s}x����)�:�WZsU5KG��D]M�ǾE�[=���S�e�!��"��"��ks8����t�ӱ��cD���m^�K��6��R�R�� ��
�[�xA�T��l�N)��^�+6G}X��ƭ���kn�1݅��᧮�:�M�Cѷ٥�����z����%nZy�xL��*�݈��E.X|���u�����9�������8�o	:a�:+ʷ���Kk�Ub�X��z%g��0<�`U�VS�g1�[7��yrW]eδ4���w��g��V��'x]��<.n׶pۭ�5ʁ��{a�PT39��Ꙓ��eJk$r}�3�3j<so��D�g�ډ�^]���w�Vs|�:K�1�^#��<��A�F���Ȉ�C�զ��z��ٴ�uMZQZ�Q�G-Cj?�S-�֢�wK����)Z���5L�әh�eX�"&0��5�i�.	U-�َb`�Snf��+1�f��ij�YQE
���ֵ���,t�]fkT�镊�*�6�9��Kb���fe�����XQ��-�Z�M���̨��䬭m-��1�*3\�-��l�K2��M77��iQ�ݔ\P�s3-+#[�Ţŋ*WY���QW
�mk�LsT5�4 �5kJ��,-�,�z�TDR��ʪQ�3)P���-��E�mZ�j6�D�UDM꘶ҕj��L+4�j���
-�[P�eu��L�%<j��U�X�Uʱ��mq�����V�8�p��Q���0�mV�uB�����e3)��Wl�n9��k\���e�VV%��q��(�mԫ[�m�J����%B����u�k-K�+bV�En\D�RڱmU�Źqb"m��&�F�e7�
�U�P�ҋj�1�ffL����Pr���ՊZZ�WT�L���Z�X�4r���YXbV�Xb��(�Ɏ7-L�r�V�E�ps�1��0KQ��re���q��!s��^C�^��(�H7�{�VNV�ܽ����T/����"�i��z7��i���\5v_�K��51WM1K�=W29ƜJ����7s��Wӎ�a}cYhL۬2��s.!Ծ˴���27�`�ڧ�xמ%�L���d�����:�m٪S��+�i�����Y��5M�h��ȼ���p��[Y9��\%�L\fia?
�WV��n'S iL;^fS�~���nŉ�������Xϥ;̷D�ez��(�E�ڤL�!��.Pp������`�F���n�T��$�ǰx�=Ӻ�}p�7�=$�&�W��_�( �4��"�U9�k��S�u�'xn`�"v�9�׷�l,F�����w�Z���Ҟ�@�.~��l�S�"]zN�.�e��+(M�-li��>���}O�WYB�ĺ'a�rvPRr�<��X)vo��2^���\S�|�@�N^�o=Y�a���5��]A��O30X��,v�y_R�&�J3'2T�Ի�2�^]c�e�
�r<�2[���e��L�%!2���٪����tŽpl
`Rv���V80��:�[���G�x�!��,礸,\�(%�G<�^��`|���q�v}�Nx&jam_n�\�0�kj?*�
c.��s���{\]��w�Pb�a^1�n�d���a����~�b�}FQ����"Uw�Z��3L疮8�
�R=��]����\im���3��e)�����s�bh�?����%nk+������2`b]��r����j9�M�:4���=s���<�+!���.�k���]�a�mS9Y�%3*S�Q&+����xK�_��zz]~���f�
���W�Z �{U(~A���g�פj)���q�;� y��wR�
�~܆塚/ #Fqs���2ߕ��e�5Ʀ4<w�I��´��x-��]X��t�{���?[.�Nѓ�t���Y�0v�²ݺ�m�x8���%��<'����<��/w���+�'���L�++}u��CF8�=�-��X4*�8K�b0��Zk%O7��~��a�Ihd��'Y�}�j.��[Hz!d�+t���7s�h�I��f9vz�<�ȽLQ2�����ʥ���h��{� �i��r�S>[�yW��
�I�k��e�^�
���!�x�*�P�H�f)|ו:
��8H�FB_�.
>]{�YÎ����	��6K�:}��ձ��.Wg׈��a�:�4FŬ��^��|����n'<b�p\����U�^�!V�hS��XBW�8 �t��	Jy� 7�B�3�K�I.�M��{ل��Z~}
gݰ3:{ת���5٨t����|�JƦ�6:��1��hiTzW6{p���MrU��k�}}��
����^�u���5��eTY�ex9>>�:��	�k�H�R����'�4M	��<k[���r�b��rs�w����7��NS��ِ��Nx.�����n��z��r�sFA��]���m坳U��������M>2�]����X�}=r�,�����n�kϋ�㵈{C�[�e�"��|Jr�8,B��(:t筰.)ZɊ�\9���0�Y��]�/�>�<�S��׾0o���},�%w)�	J�=�/ �F�!l��b�ڼӻ� �cs5��t�/Ummu���;>VIw��\�y���ޫ�\/���)x儃�雉�:���g�@ղ�	�4�&��.��*w���o�X��CV�����Wf6��|�\Y��1��{z!g�����B��A�oIιZ�Ut�3]�z+Z͗p*L����Oa��&�ܽ�3ޙ�y�D=���y��zek���c�<�V��3�j��+]PS��������Ϭ��^7����0WC�9�n9������h�E�'���p`�7�p:�o{��kk�,�hM^6E��}��L{1�|%�>�Oy�S=�ױ��	0�\�>o�f�o���m�n�1l5[5p̢�UƷu9ggj��:v�p��/�͐}��:<����di�}��y�6����8�tU��o"g��W�En0X`�_���F����de��z$�
�����*�Õ�\}���{˴���`5�p�%C�z�@C���Vu+�n�i�c��1�GGo����W��5�"���p�D ]�'i��a�i��ݜ���,+�7��g5Q Ҝe3,g�Nkk����J243�xz%���h�Y�5�j�Y�5ֲ�E�WF���hCK�g���v��=�8yx.���2�h)߳ӛń�=@�f����OZ�U�n�
u��>�uV�ƈuSj�Pxv�/!��T��g�v�GY�C��G�,���!�`��g<ʼ���`w��߼%�N*�v��*�N��x�}�������� T_K�CG(eL3E���M�+Y�6�v+W��4͙�����0J��O{�����`��;(���P����r�zT8f!�te�W޼H/zp�l�"V�u&}F{�;S�FT0^��۞�a�+�����1�7�����������p��e���6i���!�*�/��rL86_�n��f����~|�-n��Cdb�Ӛ��왶�gXP�.��_n7�cv�]1u�8�u���o;���̈́#dM�Qޏz�t:�vѵ�龴���}��<�~��6��k����t�r�Ļ~= V6�QA��O]�<�"*�F�U�J��J�9κLz�;Sp��:�����r�st�IA˔-Ę��˦tg�ܷw�t�3c�sپ��,�Ӥᖈo�S�xAny�9w��ej�g�Vo�%�!k�b�R���wE���/�^�Ѐ���wz�r���I���|�����<2���"�V{�^O�`��>����o��9���ӎ�Ʋ����Xd9��әq�2�3�����'�t�I�tI�>��çk�edY���^
�׹}iX�阼	���*uLm_mƹ���vȒ]c(A�b�
����q:��#��̧��R��;v,t�*�c�h�YP?y�m���wy���%P ���)g]3}r���JUt����x�t72]��tb���vxv��&�񰐕�=�\$�t�yҀ�@H�"ؓ�OU��Z��f�n�n��3E�a��Դ�iUD�2.V�\����E�	(��d@N�mJ�[YSp�z�qS�+����E�ɘ2��Q�j�3
G+����,
pܧ+_mM��۹�y�;��⥵Q��E������6?��I�;^�1k�(3fmu����p�z.�(�ux�v/Z��a4�f�_d�n�U��{l>�8�t*����u��y�.SU!��ӂ�>�x!�hm`�,R'a��Sй<7Yn)��v�8F)7��s��;�_�>{U�<�z��Xh��kPiB�u*����*�:uL�<%���c[:���|��6����b��y��z'㞞LIU�`x?@�_o" �[]�2����.�ِe�����V8Py��o��m����!�K���s�)J��r��ʭS���kWp�Oӧ�^V�vωWr�����o��s���ʙ���:�LQ�7i_x^Mw�9�\W@��u��%4r�蕾D�	�\)LWY�grl:�Ibـ'4{�]%_��CnL�o0T޳C��Px�}�Iu�mY����}n�/�R�p���U[k��0��S/�|{���H�� o�uT�^O-	��|C�:��b�{r���{�{/����~�8�L{�2_�����(*�8��|!�zOC@�[^�QZ�|��LCRyu�Pü���t׫�w=�of	^r�5X�=���d��e�ݵ�i�X���`a�t.�|�yH��i�p��ۙ*��a�ճ��涤r�7�A�M�4N>sݸ���}�ؼ���P����hVox��۵ͣ�݊�PL������h��+�����.��%vTĽn��*j9I_X�1�1՛��i���v{6�n����)�wMչɧׯ�� �Y��0]��P�Ԭ�ϳ �n[�݇�`�}.S%�J�#;�\qW�Y~yے{��Uޣp_Ce�����/,���8w�iԪ�U���p~D��dT��W���a�G��¥�i�}x�(P���Y�3>����U���&��\��Z��Sq`�9�h\�S����x�:�-���z�z�1��h�����@qb�S������/E�z�qv0�[)@�>��'��f5v���<��vG�� p����ۚLCv�����b��|�$�{ɓ�NS���fBFNh]Dwr�Q����F���@t��<�2�{_�n��g7�C�����,�Z��Nzi�1`�:Nr�^A&��d��������l{G`�Yh��O���*,R���t�Nm��V��s�p��//A95*�����g<Җ�
��Ã�,F���vi�����ܮ��@�x�5���H['{}��3��A����A��Z��U�V�v"0V�q�$���6��/�]�7���0~!%)O����4m���nW�zKÖ}r�yS@򹔖�8öJ��'� �2��'X�W��w	�V؝�IY�Y�N��O�)�{�0�����5���lXk�HDh<��2��3!{0�o�vns�Bg�x�q��צ�N�tQ/W*�j|��1�價JnY�x��"�@�H�%�k��pu[ Uޣ����=�hg��x+Pԑ&���½M&W=�C0oLPy��t�k�ޓ�u���,!�@f�;*۔o��;�ϻ�H�i��4�=��g����;xF����}��
�X���%edG�`*{��7kw3�>�=B
�v|��W��`��پ���̠�.�R�߱�2|е5����=>��5�����/rLa5�봭r��nN��K�G�E�x"2{B��/OfI��M��U��5�c�}V�sŒ��=A ]nC�EA׫2b��-V����6L�����eo���g�Q��ٶ�J�R���C�u�v8��*�O7���>�Z�Bo��+��P�ڃ��S��|�!�3��g|�����^�[�`\�=���<}��,���(u���<>�ʩI����e�#>��v	�몴�}ktxL/�:ٓ��xC�(h�w�	��F�u���i϶ [ܜ�p��R�91��W7+B��wX0�r���e=�g<�̍���v7��A�mξc�܏�;������{m�9���Kŋp��fv�y���R;���Z�1���M���UL�j�n�Wd��Gwڣ�䘸��H�t����<t����-��ުK`b�ğKΟ����nh�`�@�Ď���h�b�Y�2����^'6��=@��>o���͌�����<��x��ـ
�"�O#���n�9;3&�CY�.�O�{ݼu�r{x:7z.�8׆����%��}Wq�B�p^$�㸩uͯ���W5^��F���ݛٸĳZڮ���6��8aa��e��`
4�<ɷj��r�5/�8>��.��xq@�&�иi���u���%���%Z��Z�%R�Nң�<cX�o��n"��ϑѼԧ����9OùT9�wL��([�1N���kZg��^�˽\�0��Z��~����AwZ���ͭ����I�|�eM��VJ}�_��Y�E��р��9[T��
cY��� ��P�;(��ח칅���l�������w��gtwe}NCw���eT�ج*a1�2������������0uE�s�ޓ�rj���,{�4Ϧu�:���9�Cɗ[�*�������|(Ɇ�!৚�7��KZ }H�:�ǵ:(�&�yO]s�W�6]�J��;�N:.�ZhL�R�(�&+vv��:q�znWlV��_[^3D��]�QO&nD/���P����6�֥��w,�xF+]���V]�Ift6��}��]>=lq���ҋ�q��kG�mz���Y]]��LiL;^�zpIpV�/�`��{)�L{%��O'�R��Ok�]�=�r�������t�9r���d��==�B5ڧ�i�z����s�o1��!L��J�F�'Bg~Ip�����@��$��}Ru�4��ѯxc�?[�����8��N?��*��'��W�SZ9o�E�!5��������Z���.����:}ϦAyQW3�8��<p"�xıH��g�o��\��ⲱ�{��\��[gR��/�P�����M\ʯO7�����Be���"��V����:�e-��-rb�5A�j=X>��������]`�r<�2[���e��T�0@�X��<M���w���� ����ϳx�3������b��R����)㾊:�Ll��U�����y����mn	U��X�d�$�r6)���}O��L�u�]\Ɂ�THz���k&w�w�ޏ�\���t��a��� ��2�(�R:���w��3��3�ﻦ�.��+iГ���Q2��u�793汞pI��i��t�z-�f>J�`ͩ��4f]�8��Hbi�K$��yw����y��Ɛ�>�ַ͡'�d��H��<#)\3��M��H�}Z�խ5�nf�Dg^���/�����=�z5K�n����[�x+\kh�T�*����O,�4���T�З,7ś
�4~���M3�CQB0{��N�@�cxB]�5���=�7���-�Ԏ�o:��N:�����Y�;ycӘ�kJ�jӷա0�[�HZ�i;���AMSTe3�÷����C���kzf����N[qJ/o6S�x�n��������C7�8CƻlVQ^��j<��k�Y���j_��3�����f�����v�S��y�iP�>eƂY�o+��J�+��m[�ŇV/-��;�8�x)]{۵n��7^_74w�Vxrܬ�w��ʏ��Mw;�����x�@FM"\�fσ:R��6��7.տx���#�)u��&���"��2��t:���a0H7Sq�eŁ��{���K�cBiS���|�Z_^W��]岃,&2���<;V�s�� �I�]Z�Yr��5����Փ/kY��\�i�H��t��יw��]�|P̅x�֎�bj�fÎ*T%\V+^���,ܫ�=w��1�����F�9�f�I3c��VFTT�m����|(]�l�b�T�*#Ϯ{[e� ��i[癔�t��@b��Ŋ�w�M�[�#5&-�=�1�w�[����4���W�.�8�]�=���ᝯ(E�:)iʍe�1�1ɇ/���h�I���eh*�'����Y~����[��Ե�c�^��
{����8�j-Gu�o���u���x����=2��Wx��Qݼ���Y:n
Tt-y&�ǋ�����C;H
3�$f���N�y����E�zB[E���%[R9���[0����z��R��9��0�_I�;�T��82���Ԯx��:���1�.�dpGM���ïC9���������mge"�]�j�Gar?���t�S،�ٰJH��4u�P]���6�ר3�����T�ʋ�kTva��<TM�O����í�Z|z��״#l�qZ�3a���*t�Z�%��F�9��ס�o.{�@�ag+BK-�K�ԓ�`�}�讑n��8U������#�@���q{Pf^@WC���Y��*{ԝ�oVں�}=�L{��9�b�����R ��u�Wa�$�ֺ���#�!�)�FW$,���,�u�h[=�\��I�EYV���V�f�����l�����j��a��%z��C�_\�C�A����!7T�dS�~�i�&�-9z�V��z��o��ΚU�^=q���n)v,5\�u���%~6�9ݾٗ�NN��˝;:[-��*��q�1	��@$�A��V(�b֨�Z�֘����Ea�
���5K�����(�U�J��XU�i�ikS�5q�F#U�EJأ�a���mq�cjZ-��(ѶV�U�Q�Ʋ�R�#Z*�TҶ��L�8	Z��l�+�e�X�ԥl�ZUkm�Q�ӌ-�[k`���c5t�FԴ�5�T�b�m-���cUAQ�[���QF[s*�aYZ,j4r�h��Z�s���X��h�V��%S-1��j�m���£j�,H��QAAJʉU�9��R[��%]T�Kk�1Tf[Wƪ"�+iw�-ލ)��qƴ����%X��R�r�ih�V�aR�R�[V��ե��[�\��₸��
�Ѷ��Z-���ʋk
����F٪\�(3ƘR�Q�f%�T�%bV�m`�Z�j�V5Z�Uh�4���PZ*�k[-�խ���n8������+r�*��DR�"[X��¢��b����)U�Q�*"�� +�(C���ӯ�s:��u]̀k��؉�U�����,�u�1N`���F}�r��s��lgW���ئ,��U�\��MOM�-=N��3v����
L�� ���$��Sܱ���8Rμ3z��d�{�t�ػ���=;�u�x���R`��쪙�g�>;�pQmfb�4=�4�1�hÁ9�7�nZ�D݈gn^�.��|���q�P�='ܠ�X�����뗦cږ7��;���ٝj��p��'	�Z�r�<7�pCm <�d���uݶ�>���u��
X�6dO=[�;�G��N�[�ۭ'.\����+Qt z�p�o�V]yxq<����)~��wfbƘ�]ګ�+�R��V=\�@�R�v� j,M���#�K[�~��89�[Ѳ�SO��]�g!
����-�^�<..��Xb��5��r�uǸ�����K�<z�M�5�w;�f���0sK��z��񫣡S+�v�)�d�Xm�5��+M!F�^�&zu7�lʨ�D5�^3�����8&Y�B$k��pV����׷{&U�h\&��JL�g�d���S|6d$!����}֯����7�������u-,����%׹'/ +����ǐł����k�l��_kR�N�`��Ͷ*ڈ�
=��+�^�2��cR��|��Q69�9����/��z������t-���o���?p5�4��;5����7�][��l���2z�,շ��'�s�Xn]�v/l;뺺��9�\s�|��{��+���/��P�}�Є��	1n�}[����/�hs&�1�ʋ{�S9���^��^���zŬU�-��s�6��޷�*�����_<DU����].^�7ᷪ����۴��ٕ���횟g[G�`�����u��K�B�B�O$7G����[�����|�=��T3v!/���^y	��޲'���El��'�x���)��V�A}�_��� k�غ].t�/|D��ݞ�~���腜jq��B��p�x��*��GLjÕOs9��百�^�=2�ɂY`����u;8���'���1��*au�U��\��*^l����vo�J�f��c�fN��ӣ�n�{s%M�����}���a�n�k��*��u��&|���r�{�/s��������z�:-���_	��V���|�u�oU�;�!Y*���k���8���>���P��z�E��jB�oϥL	��{1���AD�A��?S�����#C�-�����vR�@O��K��9�v�E�]��j��ޛ}ק�M�C�շ��hΓ���4LMfjX�B�|7�����ö6�ݬ�4�\��,s�n��X�ŚՌ �%g��:�uNmNE0�/xr��U~��l��q:��̭���H��ћn�U(��u��#�2s���P�~��~���K+��hR��n��҂}�:���+��C�|'5�ז����ۊ�������!�v�Y�D5�SuңňO��Y��L�.1s#��z���p���a���1�����P+�#�:G�e$�z|��F�[`��ձ ����"�	�M$�3}-�t��>��銷aV���<�aQ�p�N��[�~# /�z���}~��e�S���Ԟ_3�]Jh�P�H�������t�X�Q����#��"L�)w\�j�y�<���
�K��ғ��R5cT��p�L��WB�ST(Q�aBmg��쏔����sٛ:y+j���c;	d?�D�33ò�S�FUC������`
�����T<�G�֓�+�}U�^�-���� ϽU�z�p�4�%�c��>RA��=7{��w���m��%x(:��[��m�^9�)�w*�3�`$��ₕ��:��)g��z׷qd3���:xeP�:�)F�)zL��X)���W�,`8�@_b�K����Y���ga�6Rѣ�T�Uؙ�� ѵQt
��[P�L��6������9=�h���GSt2c/��B�驇|��$u�Z�櫵j�[�3`f�ش`u���l�j�8@����L��)�����51Ӯ�e��.טB��8Wq\|Lf�������YUxi��R�-�~�����ڻt4þ��GE��Sf��6�|�eU���z>�oM�u�t���1�%R�l7�2^����N�;�j�`�?S]��R���~5C�6ݚ]�"���i��j�ܺu�v�Sx~W]�k$I=˶LWn�T�P-��pJ
�]]����ws�FS0=9"���^�
.)<�=��f{"�c��
�K��.�%b��,1K:�s�.�R���y����f�u�v-c��/EE�PU�0�:�E����$�zU=�u -�$}�w�����Ru^��FK򭁧�s�]6}B٧t�(�&C�Ɏ��)�
R���e�ג���◄k���!�w<{�u��T�lץ���n+ OP�珢+G
x��^5�7 ���o
O���^�|�=�,���^�o=Y�a���5��E�X��ݍ����n`�b�+��;�0�5#�'j��b=��=է�=���:E����]	�K���|��
v��G|�����"{w�s��p�>����䥽ƫv����z�+~Gg�������e�K�i�p�Ą���g���ȳ:���vIjs�Ɍo�X�X�E�n�b���R�Prvb�=-��L�=�`A��<���6�}\��ɹk��>�D �T_ƕ8o���V�m���Ş!�T��s�.a�<��a�����{����
�~�k%��)�Y<.���:�6�~֋9�a�x�^����T.������0�uc0�`�biO�h�d&���B�:��9�L�V$p���'����}��Z�$ϸ�:yM&+�hxR�$�׿JA���I�[]b����d3�B��n�\_/j�(w���h�<��dr� _�`�~WS��g?r�0H��Gε���zv�=P��+�=��ۗ�g�����
���!�zNu���%*Ձw�;E\�ߓ�le'����K^?.+Rp�����#��)x��
�C�&Nzy:��$�n�������(d�!8p����\0��QJ�䠧�n���`ӣ^�M�1n�R��wz�=z���-�d0W,����r�r�]G�6��E�����WZ���9���syf�>�ϐ�g���4���&�k��#ʱb=1K:�f�`IeiNmj�ޛ��q���]�y���z.F�r�������Z��c��]�uv��;W��uti7�X���'_�X*���o9��ی���o��X89o��%w� �����0�B�Bϑ�_Qܰ�m�!�ʤ��)�;���74���g��w;tc��1^���ʥ�O�W+Q�W��N~��-��ދ-gV��P"��N:0L�ٕQ�k2����}[g�5�D�p�2�t9�ܑ�'�E����+�Эi:��U�=�"��]`�e�z��L6����v=/���>W͏f�VX@,��/�F�;�;֩�9�X"�9����*N��#�kַ)�R�x�/o6�T~�+���������B��g��Z�(<ӛo�╬�;�����������ꃋg4�?\�`�s	�a�dV}��2U���%*o�m8{%�bF�f���w�Pz�����)O��:�	b#��B�Bķ�$�`�%��W������{Y��Ώ޴�3qf�c#A�z�zȞ3��[ H�1�M!Lu�i��%d.��{�'<��+�0Y��CT�/����w�i���ޞ�q�e�l:QxO3�w�^��5��2���g��K��j�BA�V�嵵�<Ӣﴢ-C�rX7�g�9���mf��m��|2�d����1cY��V����΁3��wA��x�3%��=�v��\�ar�}�}	�`�tm��_��b��닡�Xo<�[��}��=���Bȩ�<���δ���ߊ^+��;�oD8�}���}OVp<������2��-v���n��<k2�>U��Լ���3�[墥��]*��dQ�:*0>�a�>o��g'j�kɍx�8Ms���Mr��nGX<v�5��z��F�w:߃��z�ɘ�?z�5&-��Ĩny��Gic����įGE6xU���}єR�o4��gøZ�+<z�'U�����S�N�K���c:�zȂ��W����#O>e$�8�wY�'�lx�PP�\���\�sPuJq���!�>s[Qj޹�Xk���y�y������y-�5³岮��bxІd�]38�D<�^+�R��yz��z34*��h��<����Ԓ�=}v(�.�����C4�����y;8Ϳ�ϝ����)ԇ3�:�tU�M#��i���X.�9�U��m]���}/�oٜ^�z�	����S/���� 2�٠�����O �n���U`����YI�R�
0��$�{w}S����L��Do'I���I�7͎�K�U���*nտJ�ތ��_iJ�j��uwu����Cd�b.g��w`�>��G:��#��i����e����_	�.5R�{\#��c3�O���r�r)�����o����c2����I�h��F�4eL��%��C(J��T(Q�Ħ'�V��Jsޛ� W�Ab��}�K=�Y�A�3=\���C)i��+T�T�W���wc�E���z�P^�-�wKX�u���<�g0t�.�����EoNH���CSz\]�Y�f1D��ю�70_�64O��!
�Z<3�Jx�_�}���!�Mӊ
K/4����a0�\��-6�
��3���C�F�'Z6}+P0�.�y�9w��i��*i^5���=���l�̈́-sA�_IxΓ�3J�JV?Y����i�G�K���$֬�2� ��=g9oK��/a�&u����D��O ��� R��Oh�����5�m�Y�8�8�{7ʆv��ݞ���LJ��6�C�jĭ��e~#�2�t�C�n����5�[�	'����g%0pdK���!�e�(/��LVWWC��cJa��0=9"��S�[f�ԡ����~x�[C������&:RX�JK�	�Ԫ��V��t�9r��53%X�:�nU/pͧ�i��O_!�uN⋾:�T����R���$��y��M.�Q�W��Wd�w2=���쵕yw���E��<~x4�[��֚�{ha�+MDJ�� %\{x�l��'OZ੔;���c�:�B ���]q1{���*{Pf�2:�B����=bN����øS���Pn�ih�}T��=}<� ��B���R� ̭~��|�����=�;���>Q�f��CJ�p��+���U���=n`
3{�٬ܝ���q}�MA�X~9�󺨲N��c��ϧ�}S�W+@K��N�
��w�,K�_��&ZY�=*����D�*�L4�ɫ�U���Ր�f"k�4��Ч�,g�lu�ɜ���Pt ���l�]u�jafe�pj�*|�y�2d���ɋ#tE%��^��e�ތ{|	Y���H���*p�x�}Gឤߪ<,�¥����C�_y�=~���Nwa�O�:T�x.TTM`��%�C�ئ5W�pz�f�r�:���f�rG�e��	�3kZ��c*7e��zU?Rbߑ%}"!��+[lX��9�}�+�U�೚o���B.	~�&�5�R�}Q&+>��
u0��A�y].x�|��H���T>���u>�_�'���<��d(����yhL����~ .�%v/`E��|W6�-�43�(0z0����߯%J��c/�;�^P���>Բ�R�0�p��L#��%8���om�ʙ�V�]SZ�3������7E�\�^��IN2�mt��f+��p��(��˽�W½�٬�_��pa��p9����5�������҇姅iN���o�����z�\����Aa�;�
��M �g!L����jt�։�2�?�i���������+ۖ����6�+i�%%�/�칕\no;�7}zRs�X4-8K��0��d���}���fA^��A�a���f��Ý�ץ���|2|����㹺��9AՌ>-tJǡ�����鴽���*�CY������O�0v�?;����Љ]�,�&�aT:�����\]F�c^~�S��3;R+iP�^�D���'�AI����qM��Q��`���vx��p*cF�׆��]������U�nY���di}��%1r��fUE�D5�^r||#�l��5��x��}t���~ssmxת*�R'hE�49��٘��8�X`����5=���[�� =��I7�An��olI��;O��D_Kd�(p������~�禜�ŗLs��L����m���A��2�Um��k�e�C֍!:;L0��������g��$ I?�H@��H@�?��$ IB����$����$��	!I�`IO�@�$��!$ I?���$�$�	'IJBH@�x@�$����$�0$�	'��$ I?�	!I�`IO�H@�~�$ I?�b��L����|P � � ����{ϻ!����/�9\0�oUr�$ U ��(�jU%Bwz �
H �  �? 5�L��      jcM�*4 ɓ&@4�12M56��= �i�0� &�$d��zF h��jh��0 hsbh0�2d��`�i���!�*H�h�И�4�L�bb4��3I�~RHIG��,wĒ&��Z$a"	�$��a��V��P$�>_WO�~����������u~ynG�Q�T�R��&pH��P�E�[^X�pRFP�ҤJ�1T�!��e��իюI���2p	�{=�^�U�UUQUUUQUX���������I��Z����������������ϳ�$�M8u߭�0�J0gEm�^u[:�ʩS�ڻ�7��.xG��U��{{6%��jt�)�&�"֚;vo�1��[��n��������)�UZ���2�!_����-
��\�+��l���ST�&ި�R�&"wF�L����#E�aU�JAl�*��R�p)�Tf�R{T�n�S3JR�SRps����4ֳ5Zs�29B�&�F�d���n�f�f�M�C{�]�ޱhˎ۪m�5tc�C����Z�R}�]?y���֥9��������g�o5J�4/��߇������ν�9�Qv�[��M6��ܼ�M��qgrK̍�{>hڈ������׋�����)��7�U�(�Y��j �%tʋoj�n1�א����{u�xt�r�#)evc�4�o&���w��2.%�VfM=��z??������;��1��/��W���H�[���mZ��ת$�F�xuh�"I9#^ݶ��OL������'�SaכmK�D"DQ�sׯ��Zm��c�m�ni&�M����m�޶�`|%�����@���-�۶�6�6�v�na��oM�۶�6�f�D��PK��˔�4��Vک��IUUi�kV1�U��U�h5X*�˂"�YaR�q*Ԡ�X���e�"{��<�$##$_�	܆���y^��)�#�����E@�%��U��+U�`���>�� |��
�{z�׏�6v�ݲ�;e��݇�UjW�$������X1�Q*ڋ�������]��d+�g8��V��=�9^�*(,(%-�Gu��ձ�Bs#�pA���||��2��SA5��E�̓�H���f'��0竳�B�=?��XN�g�B�	� �t0����p�1$�0�P̒,���X��D��i���l�����E�G]L����)O:�$�4��0:��OWw�;|A�N�D���Qw{����cgNwtu��M1yl�����mR���
�� iG��<�y#�h�G����:�XI�:��l��U{�%Lhr�"�0��q������dfDo`k]���I0&���+�\\Ќ�+`�8:f�z>8Q�m�1$<@_�Tޛ��pX^�fy�e^�ˎ�B<���)Mt�����[��Ń�h��Z&u1\s������n7�W��mZ����y�!�}O'��O�}`3�����v��@�Fc���8{]c��Z[��^�x�������I$�o�@��|�򓓍�?H�'�{�����
���wc�F=�
���g��+��^�BOpb+D�]�˚r�sL��e<�֒�1���"b��&�k�>&ػ����\ݻp�Axs��{�x��n-3�t�n��8��u�ќ�Uq�U��Y�^����ݺ��ؔ�fN��~z��KZF�Ti�!�/a�SՂh*�:���\�̗�}�A9UՉ$��D4#��~7�'�p��[��qŦ-�ΌೡE�P���E��T�s�i0�2L��lns���-��q��c2ݭ/�o3#'��l�V�� Od��c"ǐ���\��g	�G�l3%���cC5E������4SƋ�Sy[jҊ�.�:���{gi{�ni�� �oH�~�Z.&��"�1Ɉ��X=���I+�w�hp�9�@�o��o6�=Mw+4g��.��Ӵ��-��8i�f�~���ؖ���������v�;�������9�1ʽd��D2���Ì�o�c1��OZ�GyhI��8�o��b]T����.tr'i���0#�y����eC��D*�2#�(����k;�D�=�Vu�u
���k�|z������s��;c#i�31$�_��(J=?|L���l��ةAH�/c3`����z)1[�w��V��s�pk�SKZTs�]6DEJ�lJ�@�&l)�j��ܠg0-kFV��ޚ�FȮ��_(����=�]z��p��-[0�EN;��
o�1݅FW/��c<��V��2�+N�!��-(�`�\��:�\9i�&�Nq�Z��Y�E���!鲬�g^p�q���J�ʵ�p�W:(t�/�L\R�� �$�'
��#Zg�12�ȓ��E�<�yȷю�ԯ��Z�����#�"�S�£�"��&(�2e��D-C� ���pH#�I��Q�-TI�<�`�;��e���N�HA �3X6|=H��ou�A5hH"���CA�/���H�@�(���B!�|Ã��tt�vQ]�N�,Ifb(���|
sS!��UB��f`  ��B�� U�R=J�Db�i��E�`TS>��^I��Zc�|'����,�7���=�۳6c0�r!�z�%�0d�r��ם>l���rc��	#���ٲ.�v��^I3pR�=��J�((�n���|Ph���2�|j��n]�gX �=I��"
����.޾���O��Iބ��p���|�Mo��-�پ|�Ѻ�o�|�W� ���0j�'�b�br����i�a�l��� UUUC���"���7�ߠ�.��9^�ٔ}�we�<���kj�6{&�F���Z�%�͸UqZ�X�Cߚ��dw�<�b�l�#�خ�.ql�=a�e��d�aF�*]�R#�X�c�.�]Q(��;��;HM��m��sT�rن�����"�FE��^��:�e�*6��\���{���;Ml�O�AV�k��UUUP���.gܾQ���Ҏ�
�.Ҧ/�x*�5ꪸ)�u�t����� �g���ެ�Co#9�����
�&��Q�a�Ay��ݾ��(���vUG;\�7�<�O�tٶ�_�M˅7��T#�7����� g��<��c���>�0�P@p�(YB��
�UQb� %�$&%?�!���ɮ!f����L�rY�qfpd0�O!�/�=&�|9I��t�',��R�JXba@��!�E�ҁiIJS�0��Ђm3����h�AEDT"��

*��"(�QE��QEQH���(���+&���1
�8H_*�`�&��[�oʒRq%Ű�y罄�H"V�=ډZ���ne�+�ֿҋC��������-2�'��J1�cSa��٦�y3�d�9����a|UK����E��.mk�L��Y��"D���{v�Xru�v��Id����&hq�$J~P�
�Z%Ӵt?�a�M���'�_<dۄ|&���}�����eLγ��J������'�#�z���#Ш�JX�R04=�H�	$f�gQ���0%<��]��li�����C��֙�F	f,XIkd�8(ǝ��9�
�����</�E2����x�?�KD!M�-6J��0��ҿ��A!PHB�����b�(��IC/!�-.���f��k�����Պ��e������n�b���e$Z�-j�"���]�����季���y5<_Q�ץK��ڴ�d��Q�o���s����9�=���73`w��-<���׶n�/�ͮĤ�D���%�M���M̝�����ߵ�0,��ze�eƸl����=�Ş���ӮUl�8�N�#�;M��ssA�3z�G��j���D�/M9�tJ�v�O�$��#�͈ѡ������a��ujE�����|j"$��9A"}�z{Ȩ�+��tRҪ������71I�%5ŉ��挛�$�I�9��QQRtK�O:H��;��'�!%����b�z����jI�����R�!Q��)kY)��yMRI�[j%#3�Y��2bJ4'S���N��;�h2��(��������tD˦	إy�R�J6sN�|���_��1s��s���:N��;9G�s�H����:���¿e(���΄�t���Q�Y�Q&��{�>y>�N�0}o�h$NO�\k��R����xy{ѤT�D�N�FOAMR������i�{27N�oG��g��5T��Щx��s�RU�]]m��7�g��1�����R�H�5;�i��s��z*����lb�%��p�U��ߔ%ܩ��eXU6��\[�,`o���Ĩh��2�W���s1�Nm����d����2Yţ`�۩�U��^3a�8TJ��	P{��\z��]�J{g�������"d�����)3LM�q��d��Y����U�WG�{��G<UJyشG(�����ޒm���.�p� Kq�~