BZh91AY&SY4����_�`p���"� ����bF�      ��(R	T>��(��T�m( HP&�i,��A����[U[4Z�L��klDJ�@jkhV��kVmR��Ѳ��k%|�,eUU
��4jٚ�ƑKc6�V3Rͩ&��#*�m�Zm�U���Z��ZU�mZ��kT�f��JY�LƊ��Z >�z��l�Fƚ�jR���U(�wV�[l��V̪&��S���Y�T��Q*�hIjZ$���ERVV�d�dR�m)��ƛ�<��jm�-[�   Y:Ϯ��kw�
���tt�;�샵����ҍֻ�&�uRM����j��V�\j8�0-v@�f���P��T5�5j�e�W�  ���*z���I�/zN��m��(8z�mj����zs�C݃�gyھ��Ok,56���}��5*C�z��o�k���>�'�J���{ު��IU_|�a5�m�4�V٫i��5�>  s����R�E}���J����k�>����J�V|=�/mR��u���JC��m>k�<��*O]���޻�]٢H��O��}��>�m�ۗ��|��Zbm�{�}��%/c��[km�T�fM�4ք��ԟ  �Ϩ饴����!>�ί�w�}z׷w݂)����v�f����*��4�;��}��ڦ��}����fU�׼�JLڶi�����U#����cE�G�.ٶ�&�a�5j�imel|  .��$��^����*T��s�EzV�Oz��U=m����Ѽ����ҕ�g���f���O�z�-0��#{xޚN����y�4�5�;������'����ZЊ�I���6��  ���J;5��^{����Z��{{M)[fl�{;ԠQW�p{�J{w�U���z�f����/w�TG�V=Fnf�om]��z��U��m[cúI�m��s��5Y�����͵5[f6��π  �|�����7Nz��U6Kuz��&�W\���ǵ�����K��iD��m� >��E=r:{���W�O�45�3�Q��9C�kS6�[6��j�   ��tu�a{�y�mU
�ޓ�Uֶǭo)�z�ݏ���z%A^�������7�����U�z�C��=�7xq�*���k6Y�35�5��5��`��   1��(R����������WT�p��=��z׺�o=����뱎��y-���w�g�U��B�fޯo<Am�n��V&���
ZdU|   ۽�]���zVw��u��%�t2�k���^�m��<�͠ep�:�����{��� ���z*�u�����^]붪j��        j`�*T��4 �@ "�Ѧ)J��  �   ���)*I@     j��@��( d    '�����hh!�0 @�	I�(���G���4i��=�����~����i�b�|������������ݿ
|�s����ߝ{������u����
��PT�� �� �����O�����>*�QU���TG�qU��a*� ����������,'�d�3	�L�f2�̦d3	�s2���&`s	�L��S0fas)��f09�̳e3	�L�fS0���&a3&d�L�f2��&a3	�L�.e3	�L�fS0���&a�3!��f0��̆e3��L�fG2��̦a3	�	��fS2��̦`s!�L�f32�09�̆a3	��fc0���&a3	�L�fG09�32���&d3)�L�fG0��`3!��fC0�̆`3!��!��fC0���&a3	��f�L�fC0��̆a3!��f�2��`3!�˘L�f0�C29�0��Qȃ�3 `�(9�0 �\� f	�3 �dA�9�G0�� \�#�s�`S2�L�9�G0 �D�� s�dQ�	�D&@�)�@s .`�9�G2�A�L�9�G0�P\�#�Ps(dA�(9�0.e@�@s"aT� 9�S0��L��3 �e�"9�0 �P���	�0��Q0��G0"�\����0f\�s(.a 3*.aQ̩�&P\£�s(.d 3.a@3(�d�#2��\�+�P�(f \ȋ�`@3 ��s"�eĘ��0���0��̆a3	�L�6a3	��fC0�̆d3	�&L�fC2�̆`3!��fC4�fC2��̆`3!��fS09��̦as�L�f2��2L�e3)�L�fC2�̆a&��L�fS09��e0�fS29�3�L�f0�I��&`s)��f1�?��$�����@f��}�}��?dsF88�$�.�5���<�L��b�1f�ɉ�a٢Լ������n�,Q��+:���-o���V�kˡ��l''�
^�D�F���v	��܃Z��lֆDZ���d�GP�\%+��Ѣ�mO9�bzV��ޫC�b�O.&̼4�/N,�FD2"J��S���v�` vX�,A��p7�f����l�HS����He�kpkzR!��Y�k��A�x���Cw�$!˭ȡ��X4	13b��*[S�A�@g��ɭ`hk���x�Tw%�;2��[�aƙ��n��%]�b�m�M�6j2 S����`8v��e�n�4�ݢ�6k0�nL:�I;ank$n�B�W����[�e�Qc�x�0����kyf�Z��n�h��Y:�(F�cVE/;uIL��ki<��l�7QSeX�p��JT���*-j���,�ң�6!�%���xȊ���dRQb�2˦i=�P�QYZf�bt.POqIP�l֛7'�B�wsod2<Fh�`�Dٸ�v#���Ղ�6L���E�n��Dby0�/!�7l튔I�{���바�(l�N��[lmִpX�.��ie�I4̙�n��va�J�"�#Z��cY�&�7QHE
��P�[iٮݷN�-�y����s����M�	��5�f�7,U�J�X���цK�ܫ�^PGZ�R��uh�h� ���G
W4�"
iܤʽ��Z��HTh<��7u�ɂ�^�jB��l£y[eP�A�n<�k
�^li&�-�
��4��d&�^&��,@Ŷ��]�!�H/Q�d�;``xȬj^��ڡ�%1�Պ�w��)�&��p#�=}�+4�Ig��(I��awo]hܩo.����nJ�t$70�י#r�{w4&�=/v��̴w`�
��:C�#Z����G���,��L�+�R^�j��vV�QB�A(����+���8X5�l-��v\�L<1(��S6n�B��j���Yf�	��q}�q-%�km邙+M$ot$M�.3J����n͑�Zn��Ӡ�f�U#�P?�%�%s'*�-S�/�@�XӺ/�Ŏ�r��پ��h���ִ͊�
�'v�,@�4̱N��n�GIK d�TYY���YU�ai�;��K�Lu4�������-��Vm��ͷ�2�V^g�$R�X�Rea��Ы�[v���{��5VEf�8%�;0��q�ot�I�9fMs4�������W��īb��} �wh�1�POsd�'�`ɋke������*U�6��n��i�3r�B��z��Ԡ�km{em�Ou=�-�P:�M)��\c(�lŚ�h�h��v�^�5��lXSs0E�1X܏�x���a$�n�9��)H�E
��K+n4�(�m҃A��:��P֩���M�@(��F��%K[�mjl�Ǒ�,�Q̵l�`ڂ���'p��ԍ��I����{0Zy�v�oś�Z�w�ѥ'"�)�
<�Y7'�o��n4J	�J<�E8�0VTz��o���B�báA�g���u��k��+S�і�2�j�BkI��v��L�i�b-UL��!3�#���`�H�4�8*'6�� ��6a��С�1xġX�N��N=�m�Xw�E8�\�[q�h7�Ú�4�x�.]�釷�P���E܃.'F�ܖ6=�1R��E���0����ޔ"D��rP�e��An�\.ռ��-'x��.�*�4�wxSfZjU�H�tG ��ֵ��G`h���b��$����;�%L$�L��r�2�L�{e^#/7օ@^Br���P�/^��Y��Py�Y�L��ԁ��ez��ĕ��IV�󗗹.�Aԗ�9Xl�X�b��橗�h709��df�7~^�eڸj-�Đ�ֲ�x�m�5�5z�:�m8.�:Cl%S4;�z0n`7mfL�6�1ɳ2
i�-Ĕ�,!��NܶF��t�*�ۣ�6��Cjn��IDh�٘����6�a���;�"�*�*n�#d�R��owJ�;������l���$�V�:��{75b�j���b������rڲ)6��J�,e�������Z-�+qU�����"��2nHF���'fѱ kh½��:Bq"pӽ��3F�&
Ҏr-�%�v���Y���0Պ�R��iԳ=�
*��iq�j6I�E�.�k���6�<�Fsb���)��lu�+f�Y�;4!'EBf�R�l�!��Li6��R�+���2�q�^����=�Cn�ž��u�e<��\��I4s\��d��x�4�(�e��x��A��x���U������W�{Λ�6�mpN����w5�I�֒U���tmn, �-E�������&���*�n0n�&��e8�՗�՗­�- �O���@ޢYŖí�%�������sM�͊��M���ʅ4�K��1M��~u�^;щ�g0�;�!���� �Vii��µn�tŠ�kasb)�lJ8vV)��N��R�N�N�ݍ�QI3clɧ �.%���.Թa�J��*��j ���T�;��us�ZQ��L�tm�D-M�K��Z/��^��f�2^���;� ���6Y��B�?��/[�N�J*o�ݍѴ�V�JY�潷Cy{��J͌�(��r3�ӵ�<�d�z\�ueyn�)��9P�^��X����؁�w�С�/#�x���m����*�>�ů�w��:�Z�Y��P����VFE�KH-f啑����q�8���W�h���c����M�65�uznf���OM���kr=��^m�J�в�檻	�H�4t�\w��2ȫj��(F�o��"b��T���V�Ɖ���a�R��J�����\���Ӏ�5�z�f�wBv&�^�w0H�ݽ��mA�"�`9unm<�`��{D�-P�kw-V5�se�ch���U����H)�	�4Ue�Tl+c�Q{/e��J﷦T���k�Tl�"p�X,%-jG7�f=��F�+�hR �[�5��[E�J[�#(㳸��ڔּ�y.
/-�q���^�P�XN��TՌFEɛ�=U����alu6�]����+�&ȯ$D'����¼2cf�R�4�V����YO.2K�L��V�Ev�֭��VC;z��W��:lYPb���B9��	{���u˕�y,��v��En�Ql�#��Zh7�-�͘R�4�2-��cX��3�}�ű�{��e�X(<mٗ��R�����"qb��ii�IW&0�e�7Rމ�x_W]`�U�1b4���t�亊IMژ��ח�DqQ�$�wB`nZH9��/z-Aa�u��m�Q�V���4��0�F�٫Ȍ�c1���ݼkiব�$�rՙV#7�$[2*�ЩY(��:��kq�X.�n��"H��Tr:U�Ш5l{�V��Kˤ�7x� ���u,������Lɲ\����W�3q=tp�Hq61+�Zc�I=��Q8��pұ��>�G@��B�v^�O6�pȒ�-�R��*4���Ц���g��V��-V�I�J�2��6���v�XyU�|C�oVn��ju�<
���X�Jcfĺ2�F6�e2N5��{����]��(��BEұ�����蛂��BkN���V�l����UQ�^.S���ьYn��G	CEk��lf�r�V�7ieǍ���J�&�#��.�1a�*2]���8r�U����k2���R�m�b�wS,���r���YFZ��v?�ky[����?�l�J����E,�۪H�#	/B|���e��t��8���6�z�5���r��j5�Q�y-�clS����ZsF-��CZ�kE��kZ�A$E�2Inm����AǥY+)e��f�j�\5��\�*n���ͬ�m��¦� �jfa�^ޟZǉ���"Cwԭ��'ph�qJYɻL
��e������.X��BM��O�[oI�Mk��nͭH��e�̧�C:�m�KU#��]n]eY�@�V��D4#�����ep�f�'v��v��Z5�J[��Z�e�y�����^�
�Jᗩc�i�aQ�FS��#E�E�#�J��N"�n�9B�kUGvP41�Q��d[xT��Z���t0N���p�3�IݪZ�MKr�l{�"^�ܴ����6���[�(�HP{n�Wr"�u��x :(nf�FjQ��-G`P�٦����H��t�9V�4.��� �~�m=���F���(S��	��ݸdkݼa�ɸ��J�x��'���5oV�d5D�Ybb�ڱSsU��E�2�1CukyGUd���	P�܌ȩe	N��:e�F[.���ƱǯP��D7�I4n�]�v��]���:e��]x�Ҫ�"Y�*c԰̮����:�^�;��4�V�ic�c�h@4�r�Zr�[���1�<q�m�{��եI�W(ɹ�s�/��^��2S�7oi���N�!�M]C��}ܰE��0��n�[��xv���via��/��H�t�:�km�.f�BJʈc�4�W�y���X�#fn��D��Y�M%.��拍U�.����8+�_4��qcHo��oE2��e��k�(��n�M���^@��f�&��k�%�-��'/^e�������(��Jp��� Hf���S��s/1�&3��՘v�աn' �]����N+ʴAz`�t���EQ:�b#h6K*�U�Df��9���6��xNP�-��ź�pk�z��ˣ�D��V�2,Gl't)kӁ��p����;t���Ɏ�Ҕm�r�1wZ���ǹVq�T7.�B�X����P�Ǯ����B�Q�Z1{f]q݆u��M;:��gUn@=��f��4��Ia�3D��XCs3;�[��_��tL[��Lb*t�m��7#�xz1��aʛk�	x�� �ܭP��~Z�
ڵq ����t�f8v��D%�F�A�U�V��hF1����#�Rv�'X�n�f�T�������|k���z묕cCł�n�Y�"q���'&�j�$d�Э��ݜ��yym`�R\~��f�
	�XHa�ؑ8��Cs��Ѽ!�`Rܐ	/P��-�ҙB�"@զ^m�:8uR��匌�e��M�d�5C(�a�P9.����(����ʫ5�a��F�C0E�M���,���oM�si��Q�-e�d�� V��=�Z��I�G�vPSIna[��NT�-�-�����:ƍ1+qd7y����уv(���p��Q̓q�WY5JȲdf�#�w����X|-p��zZ�i�7I�f��X˄�D^9q=݅�in��+��x�i̢76�o[����7O�f�\��)k��ǥ�9�j�Iӷ6:%��,X��f�$<��eV��@zH"S�"m^��!��Z|�钯!����.h�̰Id,)��UC\���iɔ>�@�a%��U����d���˭8����OL(�!�Дj�(c�A��]k{Xk�Eu(R�/9��e��Oa%u�R���ڸl;�R��"�3�P8���
=���WW��fv!TO���'�ya�\P��V[ͻ�WmV�+K��V5�Ӊ��k<U�`�6���- ��h�%�jz�x�Zz���M��L�7�o�tn6cI˘�A��p���t�r:�7[gZbCM6ս��0�ʈL6���`Q�iU�'Z���T�]!V�a	Հ��1q�;��e����̢�'��e-'�}oF�8�2�h�h�r�nT8iK�Z�;�c���Z�l'�.^��*!��R���[��&&��Y��)�\5��=Yf݈&�Cu&U�u軶��553o36�f3T��ta�j��c���޼t����gm]��D^�[KЧ���/��8���T�V�3��%�F=ץ�O/%�IU欘[�������xu3���2ՊJT��Y���Y��Z&i�W��d��m���=�Y$�5��!1�t3	g��fYH��͔�;�Sc�,f��֚�d�nܻ���r���y&���F���t΅J�7XeiKho2�e7�jzVM�Z�Rb��������$7qe��J1XN�m�9D��� �[̀��efk�b�Ja�U�s�co4쳴cM��bۗ��M�2�j�Rx�v�z��YU�2V�c&BV<�ݭ��4:F��;.�9hH��t<�ʏV�
�`�a�9��[KJ��k�.5�1���H�k�!v�sЭ�gn����m�I���5�B�$$u�K+�gq�45�NՇb���
Žډ~p���1�۴��:18U�U��v���);M�Yy$T�>�� T%���$�����k�����j�!�7��vPF>)p;�V��<=���������k$�}�=��y�Pw,s5���ewY.�Qn����z��4)eӭ��;n�D�YYcE]C�C�-�YN��ܓs3X�oAmI�H�����؁�ݮ&]߱cj_sh���4"��h�\q�0��j�N�v5 )��#&��.��%]l�m�<���ڬ���E�m#^���[N-#0�Y���\YF��.���m�T�rU�"c��e<C�-s�Auy��t�+n�"�]��D8�y�]g�Y���PvGX�ŔmѷN��~��f��M�\�v���:��fx4e!��3<�Cq���&KGzu��BƖ�����($u����=���
̧�.�`��z;C!1� 0� � �O'J�m����iS`�p.O	F��9��m�R�ͽuGY��:��E=mo�52���=<+kA�2���_� ��9J+Z��=�O�,�6��W�T��JQ��O���1�� M'E����m�@r�IU��U�����[Qo���s����?g������;�|"X=|&;���gwwwwwwstq�&��2o)@e���N�g��b�J��D�g>P,�J1����(�[�*v�ݏ� �GPl3�U�`fZ�_Y�e�6�u�H`)��iլ��*m�C
t�º���v
]t�[�����WN��e2�t�*�!xj3��lu���uM�+xeC�1
����P��*�gGg0S���ENt�[u�.)2�1p3��k��s#8.n�Rk7��CE@t��>5;fcTiҲ:��l2r{�c��!��*
�xU�FΩ#��
��Ȍ��];���OP)�.� a����-�h\4`^�\�e�h�&ul�}���;�	�}AHy�p����h_,�X��$(p�ʅ���˭��4���Z�3���cV�KCx�MCv�jW���b� ��Y��t�\=�$��;;t0�Ge�Gy� "J�Y�M�AG��݆;�A��9�r��U�����Z�vsr'�bj�n��+7`>�ʹ*��f[��՚��J�H�)���%s7���(�ⷪ94����H����n�HK����4�-�a��`Y��5W:陨��(�"z�~�:uN�(ytW�Ln����J�W`�j��ͫ؆b,7ֵ�7�u��㷛Z�8iе���b����q��������*ub�ލ*�w�p؆8�֑ܴ�Y[�pC���B�8U.�	�Z�u���7�h�B$ֱ�����w��)�0r�1gLua���#ғ^��;�*L���i�z:z�X�B9[�y��M_L��5��z�AR��lא[�BVt�`�驍���Vq�i�|ġ)��fW{�fN�('�W�P���h2k7w"G&2x^f�dmL�jML47t�QX��)��U�-�.7�9d��E��lCw��tuK�ӆK��$��%9.�v�Y�`K���r��Q�t�}�z�<t�n�NG��R�є�t���ye	X�nݨ9��P:��iZ�IIH�9��=tzlsGVVѦ��Ѳ�D��h�ˣ]�����*mE(���U�*��*2�/)TlNSvWf^VI�>��\}1-��o5�;q>��m>D�	���C(�O/�)�E�]
�#sDsk]�n[�|X]x�s3Vnѧ�@�u���2tZ3���Ljԟf��ȵ?�;���/ob{(�r騾�#��ѡ�"��3uS��kT�=]�1%�v'�px{a�X�3t��nk��i����9�A&#z��9C������N�;W/Ol�ח�wN�gA[G��sM�[9����AG��QZ�I����hTd�ÎT��a2����H�nR��M�L�JH����ׂM�L�>�q���{����C�
b�Æ�9I�0��"�����5�{b	��jz�EK)�M;�S�pe�96k����Iز�@U�Nb��o5U�}č��ܱT1��jܬ�	�]�f<`cs�p�D���H���d5�,���t�me�V�t�b���h�M��X��m�]��n9�ID9Du�vɛ[���2��u�gKU`�5��j���S���M�_vj��&�a *ŝ{ܻ�='"�
1 �3�M<A����a�:;�7���+�&��'3d	���1��K|�,�s�z;�T�b��J��Zv+ȕ��$�Z�r[E��Pg1u�s@p�:'y5���<5>.�
��^P�HR�{S͌�H�f�յ�����%���b�\u�l���m��D.�������=W���aP��=���漝��)+�F`e�5n�����.�8(�K�å�}P��ڝ�B�Tv�]�3<5n��ay���ef��06��8�#Y3)]iv*۱�����1}ڊ�)r;1��t��o;o
��s_`mu��3aeO�d��itk�B�`u��G.�Y�7�<g���[Ƞ{%��.���-a��z��]�0���,5��V5�r�9���o�<��Ϩ�r�@�Z//k��h�g-�:�,u��F�^��8xSx����U��+��T�=�mj���µ-�����7P��K̝C3�E�0�Mj9td�7,�N���1���Rc�����4��x$�ʤ&���o�$�~(̫G�>�b�a�Vp�3�Ժ�u���*�۶u�1�Ss�W8m.�]Ώ8Z=�u%��GI��U�e�Z{q�Ca�#x�U-��K��Z:(�b��R�{��@�
�=���p���$��k�[��n��ŀCНɹ�\ wD�[�XK5s��������z	e�����J�Q5��BY�˔�Ɔ���)u�p`٤ӁV[�{w��.�V��zZ��Y���
����������c��#���J�m��Yr�]8����F�`t�|C�;dMG��wk;Va�*�	�[7��g�)gK�
i�:�cHz�v���ER�:풐�;7iY�����d��9:���يK�5a��O4�:Y��&�}�A�����wQdD�}��v�8�d�Ӗ0����7J�x�[�[|�%��^T�����@�G�).Z�s1���ѣ���Q�u�i�lX�1���Y�rw�`cIKb.�G��ֺɄB�x��E�$X=�v�.h8b��սk��^5v�9����i	1�ͼ�Ce�u3Md�ȡPs��uygR|CÍJ�v	�>{�7�,��:������%���rM��+x�Q�+o��N�:�K;M�J��kU���6��t\3g�hj�z�=��h�+�Y��Tdc�\�V*�a�S�9wC� `Ր����ծu}�].����?�H�lI�,����v�c�$�ل�˵{��L�jM)�~���b�dr��w'u}՟Aԩs)z�³茵��̓T�PΛ�3������c2bJ-u����1Gq\oy堂jtfE�0��jø�<ph�U��N,B���z��o�Mpô�i�x15���|�E#�B��ue�]�#�`���]Lr�Ka��^���	n������8�i�{�ik[(�wt��jm�]�ޜU�B2��f§F��̛a�ͧ_��B���:��ӚSn��d���l"��6��u�;�ҥ3;Gк����丯�Jy�w0+����1�!h���)����z��:P|���h�Tfn���Ym>7�Dl�u�3Z:����V����
=}��.���ʕN���-8h��9��\��ե�J�%��j�h��p�cXVElgxۮ8���B��+y�( p����Mj|��)n����3n��	�kt������ޫ}T&	�bҝ���ِ�vr�x��!��G#�f7+k5N�,P�6��t6�!���k֑Rg&�uP�ѓ/Z�{X29Ç�".iuaI��˳M�갣m8�r`��r<?2h9��9��4>��錔_���"�[�;�P݊Μ+q>[2&�m�զ��mw]/`7��XR�
s�kzi]m���,l�%Ћ��D�P�ۄr��"p��ᧇ�\�.`_W_N�ܣi�D����j�vs�L��jkCT�Ɋ��j�v��B��p�t��)���S����z�J&f�=I�%�J���fRTڛ؉8�]�`gH8����:�TO*qv9cT�৹P��s��-�=�쌹:�D8��pT�WC�(�Z��T�K$��3�\8��|,����zU(+�^�f�}]�n'���W���B���Ƚ���O��ed�=-k]	�x�=k	,�4	p!N�"�X����ɼt�o�u���UH�z�a�W'��u.�*hL�ua֒6-11�јޚy�a��i�{0ɏ��7��of�`��,+&����lLcX�c�N��=�Z5�Q�u1�s;�h�b�����CksضX�d�����b���+};�4�v��R�X/N��f!Fq�wo�`�N���yL��Q˽�S�� �K�	L��t^+��:�q���I|B'�
�-Zٌp/�¤4�b~Ͼ"z���&�i�c�HN�@��ެ�J��h��o>���L��[�uzd=]��ic_;�ûxA��(u�g�<���X8��������b���cs�_Nv�.�s@*��E�������h5��x�9{�R�z�.^Ζ;Z�4���~�g�I��{��3-3K�>�-+]���g�f�;б*�܋����K-D,Vh{��������p�}q\�S~��۶\��YH�
�dd]��d�W��;O�_��'¦��@ڗ|п6���Y��1�Xq�-�E�����ۇ�Kۑ\�����]��v��8m60_�=����}��;+%�t�Tq/�k.up "�ue���X'G=�ďs��4	,uѷ�����L������a�>DF6�Kݐ�3;�Y�]܍�Y�S�N�9����4�cΥo���%P�	2 ���OU����nw^+�fmή[�oQ���MJMXq#�&]�%c=����u���+�s����|x��$̃��v�.%�t+�]h�P�x9�Y�'O\�[6>F;��[����.�wt�ሶP��E��k���nĚ{�pK�����#���%�<���Z�5�r룸+����E��?܋��6��y�r9�wX���*ž��K�y�J��I�z�����&����eK�K7Jc}u׆* z;5v̾��Y����D)�7{����y�Y]�I�ި��,0v!nB�l��5 �VXO$_P�4Րp1�1ZѦt6�fS�(=�/�>V�	��Dr!�[�c�;�r��r.̜ ��y�\:�s@��&�d'/WTl�8�EA��I��-��7���ԉ3����.J�ŋPt駵K��`��uǫl>��@���2K��(nu4]�a�b�3�����������4�:{:�ʉ�i
���Ʊ���w�#{Ɍ��x�J���KX���A�H8gvd@����E�%u��24�['�f�
ڻ�}z���-�x��M�ut��j��Kq�Vf�7	yut���G.�%��7wF�$���DT$�+�����)�Yb��Tl�6���qco:�:��n��3+�U����,Ż�JB�u�Q�ܔ^�����Z�ҝ�^��S�.m_r�]�����ӷyoF�W- z7�VT� v�:�f}��/-=n����-u��mDrpeG7.�[hӬE-Tx(��ʘ;5*,,tݴ{,�P�:�������̙]�K�vBL�'9��f���Kz�ˮ찓*�3⢧�1B�A�-��a���XG��r���#1��g7Kr��짅��/{$�����0��]:��k� ���*#9���S����5���:%m����|���u�+([ppX�V�޳ڋp��JuM�G9]o]t��Z���д(+�s[HyU���)�l��t�.����7�V����/W�Ck�r��-��:24�9�\�5+W�Ԋ�T�k�w����RS��U�=�j<�\�<�o==:e�9O��Z�wY�v�wvc�B�9w��4G,nm�Kj�mgB�n��8]W)W57DR���zs����"ܓl,F�Y��[��M�cE��q��*��6*=o5i�MKx6�c���L����3Ŝ)YZ�h{�p�R�+�Κ�����k/;6*��Ij"��O_S{�����8��)h���Bڗ����1f�ysBIf�Æդ����^�,4�L�9�M�B�h�xt�o������tm� [S�d7GnJ����F��ݜn^I%aѕ1Q̂�"�!�Z�N��S��8�ܫF��t��e\�ART3��Ra�yŚ;�gEƳ��y��㐣j��ww��s�XY�Fp�:u3(लrSn�ܢ
�sP	���[K�JY��c%Ѽo�h��m�)���=s82S�Mޚ=�.�j&v�	�@�y��V�����w��pv]L�7|�Pcٜ2IF�Őh��b��)�-�%���z�2�,� ����f�.���m :L����d��<����ɥ�|���8 :�f�Jg�F)��
���{AU�օ܁��X�w�8�� Wh����O;'�V���c#pf3!�9zM���p�����`��kZ&�*v\7ڴ4�u$�-e���B7Ri��~[Z^i7]!v��N�!�����w�(�1�4͠�F��q��'���7w����Mۧe�EtW���n��4TJs��Z�ŭY�采@l�	��uP�����.;�/��]̐.ݲ������QprW��T���n�Ph�2M�{�3�D�'1��^e �<ǅeq�n�ktB@�H�YY)���jvj�8�����������qx�Vn,�+����3GI"p����r`��<R8�����ǵ��sq�m�o��7r�M��:3O9$�]r��C{���;9��ypE�2e�G[�>);�Q��nT�3��G�]���dwtqǫ�T\�.�Jr�3���4�2�#�7sTwAͬ3h�lO��D�rI9ȓ�M��N*H�U�V���u�,�+b│��Ř�*$B�ҡl!AI!��ή#?:L�D�VU�,Sb`�u�(\B����F�a[FH��1�PI�K�$� 2��"0�)����e$�����ɉ(Ų�6�1��U�N�	�`�ITE�aH� ��� �%~eR0��G�H,����G��?�i����� 1�$�H�*��Q6�z6�$���F�k-��y7~�aɏ�bZ����XI�6J�T�c\�#m&�8XL��2`!�
!LP��!��5��J�B�a�k�̧&4H,v;1T��?�����_�����H������w���b�" !�����������C��fi���ELxɏ��
ׂ�g�sV�2���Ly3C�ި��
<S�Q-��4�����6n�:=a1I�W���}E���Zˁ>�����M635fv<��k��y��c�E�R�յ��p�:��\{�z�r��ħ*ٕ
�{�&A�A���^�fLn��!vUZ���=�x2��5wݨ7�dR6hC�{	rya��*�;}lԙ87R��9Ƭf����ʹ�WU�b"�v�0�(�e��`�5dLY�z�P���/*V����F��X�u��Sc�	�X��􏆾5%�Jʩy���ܚM�y<��0ͨv1C��	�.5]�jRK����ٝ�L�EcND���aü��L�ך��:ovQ=�;Z뺊�OgQ-��2�K��޽w�\#Bٞ=ڲ�u%�[XM㎞=q�Z�t��5�Vc+΢\s�ݪnȭ��p���֫���7h �$(RF{8eӻ�)���G���Z��y��[X�;��}�juн=NU�XB=����Re����V��J+��c�d����{u/l+"�������}��y�EǓ)6/E)��D_[��R4���P�Z����EZ�o���>1�xxp�77V�'����)�uI��T�5nơ���T��Ry}�"k�+��V�[}�ҫ�,��#�@;����j����}��o�������o����������||s��������������������������������������>>>>>>>>=�>3���������~?������������||||||}>>>>=>>>><||||||}������������>>>>>>>>�>>>>>>>���O����������`]��T�t���LF�"�5a�Cǚ�XQ꛻�F��(�Vͷ�k��o`3{�e0�ff�Q �U}RV;NK�ٌd�U�TΝP�"`���uQt����+ߟH	кh%J	�yΣ:��*n�6�&0�f�T:����ԫ�'���}��A�ڭ��E�Ɖ]j���1��u�ά�V�iȭ�ԫ"����t���P��N ���-w�GtFq>q��2_a��<A��p�G��2b<�!����W+$"�%�*v�6��R2/�h��UƲ�	aê��`<6����*�Dv���&}��ڲn��ɸ�W����b�	�u��uF�a]P��V��D�q��V����3���;���V(�(x��M4$��C4L��Z���f�Vb��i�oXڳ�z������h`۷)�f_N����.��W�|��[S�+�Cn֪*��ĤYހ���.����v�F��Z��x�wu6�D��,1����Mq���J-��ښ��י��hS�I7VKe㳴�W�z���{ו��aS�h��1�]������#��fC�P���!Äc�]*�mM�l��f�+�u��
[�.�j�5�An�+|�
a�M:���"h��r��"�x���8�)J�K��P�������a`۱�J��q�6��+k	P��	��ؚ[T��f��ΟO��Ƿ��������������Ϗ���������||||||||{|�������������������������������������������~>>>>���������||g�������Ƿ��������������������������������������|||||||||{|g�����ǯ�����U\��Y��{��y��v��C.�K�>��;��.]��f�� ��BT6�c�F�s�ӸU��0�Iގ}B�.���BT|��-o��6�j�,޻|!�չ�p.��W��]D�*3X�Vp�ebmV�'f�-øUA��ٵ/e42�%�.UaSN�i},P�²�.#�

s����RS[Ǯ�&r*��MK�;
��ܰ_.�%J�K|ے="�m���s%0%*��dz
�X�����[�ue�Dg�
�J�h>��IĖ��<���Ʀ�����4塻�M���D�7�f�yԖ�+5Gu�bZ���Y�l�f��Ć�w�u%iu�K!�c�ʱ�N{�-%UZ�G;�6�8�h�i���k�`=K�������ɓ��3;�j�)kn�!`��g@�e��٦�R�#��*F�6sI<����٘��������O��)���5口j�������$ŹN���%�7��fh���ڑ��oV7��]8ɔ��G;��s���@B��n�סe����-])Fo*s��-Y�t%�B��I:��>ֺu�Z����b�0�r���e�b��<%���ն�;�Q�X|����n�1�^S����W_h�wp�D��Iq5Ǝ���\������mЧB�5E��͐i�:w�OT��3�����~M��gE7��r�i�Ǐh-F���ۺ��n`�"�w ڌ�ªs�6�en\	��+]��z�T愳oVܺ��P�NR�yBY��\�I5�B��&l�{Xk|WUޚZ3Ҍ�뷮���`��3s�q���:ىe�|:[��H3G�ѝA閺�j��wWDv��Ȃ�U��+6�t��=�Fk:�!�;�2���qޫ���;�gX�@��xe�{l�9v��D����hi��Ҷ_��L�}W�+3q����Ԯ�p��u�E�d3���۬����T!��/{N�����ؖ�:^B�⽾t�Lpk�S�ˋ���w!�e^��4�+9JW�](N[kgg6���K�õVȩ�2M�Z�RcW�
��/D�j�X�h�mU���ű�K\�t\���hF���ǹL�� ��²�f	]�/��U�I�7��YW������;u�2��bw�u�%��묋	���,��')X2������J�pn�^�.��4:v3:�3���-t���uطkV�6����q6�[�o/�O��M&e� p�#�uǵ�8���c	���BA=2�e��gRvq��sn�V������8۾ٖ�U._h9Sfb�rAD���V�l	��O��[.���0��3R�R�_m�ΗP��ˍ�e:o��S��A2�ƅeκhhO$�_�C��׉_b�������=�PHs�U�sV����bU�馞�X�3��)���,���V��آ'
��ns�͉G�Wv �e����*��Ǡ�]o��L��^��]l���in�!�L�.[$�[[�t�=����]h��]�u5#s:l�&����Tٹ�E�}�Xn;���f�� �t6i�\4�%D�>
�{���u�Bz�ՉE��%�vW`&�D��	;�c�S�m��uRQ0([���;8��֍ ����t�9\\���lr=_��-]
�H�͊�ؔW*]X�Ɠw��em�ˉ�ZgK���ώ&b�K���n��ʵ�Gf)����xw��e��=b��ݭ�t*�+�냐x���320T8/H0J�ԫ���v�ccFe*�֧�3e�Ya�̛y9�{�"W��.4ζ��
GT]2]ǹÞ)�X��V�7Ҩ��`�b������GP��&p�O���ݴ\h's|��p��r`���oD�;]\U
k&�'3�mp�R�PP���eKln���8�4�
�M�A�ʝ��m\�Wg��0�z�
Ӈ^�RA�(uJ��I�pn�^hv�N��s ���i^���VwL��zl[Z���Vь��I��.�s��9�e�+���T�K$�p�P���3B��;���s7����,,��X,�D��s0���^\�PH*�f�V5܅�H�q��;��� T�����և�N�2b�������G�����"�M�@�2c���r$�0`�y���o�[�.�PzӨ����F��b���o�V�����ױ�C3�������G��}�7_N��pl��ID71	�ؤZcW8.�L����	��O��n���цn
�k�[aU�2T|�R-�عu:w�:
��b�M�ŝ����N9�VjOX|�M˜f�<� ���hgR���`�p��;/��4�.���B��e�6�w6�ڏ�X5A%a@-�;{�zoֵj�ީ�s���H����M���zU��Q��߫�"=�f��L��+���z�I(Vf-���84�>�6ʭ/A��g1��ҽ���D,ʅ8*��፠q�p.�rp����pUG�ʃ����2K��_j�e:Q�WX=*��Ҳ�Z���FB�oT4t*�P��æf�^��M�JElu��ų{&�Ƶ����jn-�����^�277*ڛ�sm���]E�H���uC{���e���Pǝf�v:�"��Q�,�=W3��	�WN�b�ܭ:�<�GI��[��K�S$�ܙ`�;7�IM�{�S�ŋQq���M@9L��.�z�*���r=����^�u.�);�Eb惥7wJ EуU9r�S�ӹs��N�u�<d�Po����+N�ɉ���F��7`�[���̽�e'2��z���	yrl�wӖ��;2�_|.P�x�г|C�+ǽc(���!���ݢդދ5�Ε�YSi��i��K	`�^Ӽ����lU҉�3~�Uu��T��X�S/{z~��2g%�H]>kf�hͺ.#:���W��Sޕ����B-���0[3�'�Ōu�������:�K�M�a�EE��.�
�.���L[�NW��g 6\�̼ˣ��Wq4T��5�7h@K�kF�o�X�-hWi�02[��C���b�YYZ�Th�\޲�+��L�ZJ#j��_C!�s�<Z�Z�,�B�q��ѵ1,K�v�A�2��m��{y�%��uۛ��*O�S��1<@k��6��.P�Y�I����h��)&tok�5����k��^�V��_L#����pr"^˻ ��Y���T�ΰ�N�캸L����#�Q�����z+=9܆�e����{�6�R�,���BP���z��h���ɽ{g�B��')j؋�
�U�V^VR@�zQ����\�q�1�n���4���Q5ϸk�g������/4Nxlr�mv�R��e�o���趎A���RG;�.
�E�%����0��m�9ϯ�p��6��g5��:⧘����{v��@�S�J���iy7��s��a��1��I��׮��:�
�8x����+�st���A	(�Srk�]H}y[�"r��FPXj��ꥱU\�.�F$]�}t�x@faW�YCz[��7ۖ"ݰ���y�2���o�����0uz�Bi�F�<m�����w	�V�uc�����b���L�07�8�P�-�0�"2:�ۆi�q����ݏ&�W�d�ك�vr�=7��!��mt��7+}l����:�j���].QŅ[�|ldR�O��JcÅS��]zAv`�E�:�]�Y��xi���Φ/���B�I����f^�]�+���Ҕ:ʷ����AA�sM"[!,�^o-���¢�F#�V���$9L�h�Ӗ��-[�`9��^��*x�t�=x��87�d�\s�ބiC�`%�φ�ҧԫ���yM�W�#�9]4�'1:�/:4U�������}�8?�]������ć��82��ÑJ敼X�w��݂*���S��B<JYek��PTl�̬F��nT�b���b���H�*ޜ��8cݖ��v<֩�@��V!��D�bXy�����Ui����-im�Α!ۗ��U2��d��mnG�Hթ:�eM�lX�d���l
ox n߽��bF����.<�(S�ԧ���(����;�h;��ޅS;�����hXZ�۔�*]�_	��p��trt��kF��]�l�\n��ت�KV���=�5�G
���j)TD%����J�7�e����R����E,?�)vU�3j��7��V{䚮I�ܨ��\@�!C�m�K�#�`��v��f���F⸠T�.uJ����qF����s��;��2U!=uws��de��0�G��j��o떚���5�ms�޷�y��y�:��)t[�b�,M�7c+��h1��jR]@17�cH.��|8��.�k���G�wo6z��W{|Fu��$>���sl�ܩqd�G��S4�K�[��6��9����i�|��]5vl�(,[�{.�Ⱦ`�.i�ջ�wdRe,2��gts9z&ۤ�p��R�s�%p��ڲkY��� ��u=�ނP�^c��%UN�G* Ӝ��H�-�\8N�q����hee^�$�6e�]Y���(��rn�^����[E���IY;-��Ӷh;G����gm����um8��ۛ)a~h.��+_.���5���j��	c��R��ND��\��n����������}�f�).���n��H ��.����0N�6`]�/��1>�]��{�s�4]<����[Ȇh����
��;O-[��P�u�o3���F.�°2j�/�L�ϒvl���a��*҅�S�b�QC�Q���\�"�(ue�QM;�#q�)m�Ƶ��6e��t`ܫ��>b���~Qu�Q}�U<��H���SoV�����3�V�Tޕ�-������#cѧ:��Q�Y���RVRܜ���υ�B����n�z��b:��0��[�_z�;p�xm��#�N\�U�8Ӯ�( �Ic�����|i.n��\s���A]�^��c��mM��w`�����+ݫ@qG$��˛̥�1�,q%�(:��}4^�:_>�B�RI�%�W0o��1����^�>��L�9�]��un�f<�ol��hg*�;ErYtGrxk����@��2��[7q�+��:g3t�C 6@�j^�:�nIK�#���F*V�aɺ1N�)}V�i٦�=\����<���,<�Rj����6�;0�U#40�7��Y�M�p���7yfq���Rv��Z5�&.e�[��e�uo'�QǮ��+w!ij�
&񩵺E�3u�c��tU�l��Sz�P����;��
4�h��ȼ��'I��n��4Ԕ��[��h�'���A@��D֣����w�Igq��E�u����Q�i#�q���"t󣑓��ڲ�����u�7]�����p&��۶���|����0H���$��g�E�	j����I�FÃGZ64���L���������y��{̯���?o_�������������z:�r��C�֠�&�N��UD��4#dDHJ$!�	�
A����t�*�PL���%Q���MJ�~�X0�n��5�C��@qXzX��͊N�a��թ��eu���]����l�ej�8Q��wn�Fp��M���P��î7Hua��$��f���FWX/T$qʨ�]0��f�]O�@�p%�2��;7{WrVict���R��RC���7.�gP7��L+$�B�	��s����Vy��04Y�ɽ�ǋE;kl�q/,6H�~�ƍ�z(P�� �D	7)��Y_�ΥcX��t�:.��U��N���LU����2��C��tpL�����2f:裩�\�E���jA���K��U	�!HU87H���[XVlP})\um��{7/H	��Y� ��NWo)}��m�*d®+|�M��6TM:��Sn�O���f�ˈ:�2�%�L�����4**5p��i)�y�����M�yncN���D����/_�	w�R䤵�+��mǘ(��̨16{��g�e�2��ʘep�1��W�@�9��Ο ��lh����H_{H��������fQ�^�U���f$�z���.��@T�2���Y%��ee����<S#���]�MgQ�5,�N��7_-�u��ݹ�T�Mƃe�̒��i9'K*����\0B�,�ZL��.F��B	���B'���H�	$�?CJrUH�-3$D� ����(�ĆDJH2B�(� FTr$�7)�9Ü�[ssu�8}������Zb���b����ؒ��������TUTRy�,�}?oo�����~?������PD�EPz�M5E�8�Jy)��k������$�:�-PϏ�O������~?������0P�Uz�i(}�j�
�j�i��&(������"�V����N1�"j�����QLM%Г1TET�D4EU--%QCIE<�LUA0PĔP�#�9P�خ�U�L�U4�!AABQHEISE%1z�DD�E��-R�lH�ET4Q5P�QS�P���`.�)i����5A�-RSLE_s��j�[K1� �A�֦�m�m�����˕��b���5<2[4�̓0|���j1,��TP1��u����4�KZ�c[mZ��)uE�1��6�Ƣ��psV��E�1���6��l�Y�b4F����X��b#YŰm��<�G\2lj`�[mx>��V�d
��~�eg�O�V#?�{ݏS�CMz��鈭�Gk�����2�M+z&5��mv<������8.��-��`(�L�d�}���ꙋ�ȯ�������^�����.�m��u���r���}[�z��;�l��g#��%��άfxy���mz:�=fK����y�TF�sd6Ի۞W=V�ќ_�쉏��#=Ի��3�vz3��4�w<��v|�p�Q�%�O��k�{6	�`�����p�_���#|�9A3�^=���s���Q��.��ݬֶ�J�{��=��{�M�}<Q�-��ɸ��?����z���?| �.T��W˶�u�V1vv(��E綼�\nW��-�?�L�<��.]��Wِ]z�2|���L���c�z+O;���E��Ý��� 5Bo�N�
�9׌�'�I����Q��9f��`���^��5��k��/�����X`&��K=Y����S���v��b2�gׄ��u��SFX��V\Re��́S߳����v����`ܹ�P��.l��v����}� ��������]��si�Sw&��`�)5�qޕƒ��3>�d��#A�r��A���P�B�v���ݼ]%_@������.��v��5ٳ��M_|�n��IZG��:ێ�֚���t�3o�v�����uK�^��}�Ҧ�\��월��{O�.���`]$@7�b�� �e�����]FkO��e~9�8���t�z����P?_i�����-Do8�įn�����j�m���~���`���U|r�ޢ�5\��{0,��R1���?=�qL���u�=y�O���ꜳ��w&�w����S�w����ef36�E������׺�ڃ�sW�>]ҽ��JO�۾<^#�Lk��=m�m�Z^�k� �]�Ǻ�������q�y�X��G���T�nӇIޞZ�ޜ����՟����+��(��7�oð�ިهԳ�~Yپ�aw�7]��U0|�U���}�z��q����{�S>�~���������Oy���m)G�D]Q�-���l�+�{��\�!��o�'�s�-z�GW�N%���T����R����4��_
��r�P]�����
�>H��l��δbB�B�@ζ��Օ��k'+�t�sZ�����S2���d�A�3ebWSN�:�ř[2N������OS�g�X�ih����sƼ^z��Ğ���Z��/���OG��3�����};W�7�۬��d��{5��)���O��D]z��%l)�N�g-�dޒ�<�����xg0�a{z~0������Y��t��<�x���^�^zƽ��}:���k(*q_��v��;���	�3�%�����<��s���(i�
���������c����ab:X�����5�K{޳��1���7��<U��;O�_׊�y����P�����ie,Ss�Y�%�ﲙ�y&�Y��h�F|&�sNZ�n�߻�U)3���V{���X�Ub�4W�]%
6��7k��3w} ~��kI��^���_?Y}ណ�����my��x�-b2��fc���d�۴���h�4�k�;�o��s:����W�N1\��ٯ:�%��:�:E�m�QF��bwɎ�����);�v3�u��t���5iB��8Y{R-�w6�!��U<_�{%z)f�s��Qa�.J-��u�蹺�������-���<��M���"\}E���]L���������Jy�W��m9��E�ADf���ڠE�n�c�j�8�U������A����^$��5�n$�x�c��av��)�_��0��~�ם+���O߷|�Np����d�{�����̋6�=V���v�՝���wK�uz\w$^��YFP�뚃{L_��.�􆼏mw�kUEu������}�ߢ���vt�U�y�Je^�؞�����ukb�yy�9S�;/h=�pېl�l������h5=��T�v�,ӆ����?A}S��#=�9��g��Pd�a�d*ؿ>��\>�]ϭ��ᶕ��%��6%��4��g��益<�[��*��ɺ�9��䝟�"�H.�MЏ,{�R�ócOfU���(��<@Ɔ��{6����ۏ�|#�r��S�y�V�
nyW}�������:�Q��:D��O��?�)��U�a�/o�%��)!�O{���X�o��l=H�F_g0.�����8؍>��r}ԔV;-�QR��=(-bf]��;��-y;�����a�K2u�ރ���S>�Z�oG)�Φ��T�O�"��9����Sɺ:8�u�ˤ���L�]q��e�X?n�)��������7�ə�cS�~�-q���E-����/$Z�3�e^y-�u�D�_F=�*�W�uZ�Y��A�C�~1>��i�z��6m_���&һ�2���<��-�m�uN��*/=$v�x$���[?:���e{Ư~G�[c>F�3;�fǤ;�iw�ųe�8�{2򢅞�$W�挓�휃؉��11?�}+-�r]�5+f��RK�A"�5{t��s�x�R��Oﳻ榧{�BQT'�������Zq�W[9�j����\�w�|�_�7������KL�Ȩ�G���Dd�m�Ο)�aH<=}[DS����gݮk̓�3ڞ�ea�=*��k�޻̈́ʲ�3���}%��G��W�ڽ:��`ó�ZU�j7'�S������<�O~�W�Z�\M	��_|�v��>��P�t�v�ٕ�|�NB�]��Psl�C]�ϻ�X�E�wL�v�kD���̵� �W��l�5eFe)u�F,A�k&�.VwGyZ��Y�2�]�-j��C�G[A����i�ѷc�L��Ʋ�DX�\��V�涺,�jΎ��)�ԺU���#���g��T��z�[���O4z��W<�6�e��M��ty�p4^T�C�4I��o#M���E�mG�J�^�x� 	�?U	7�|<�������˾�W{��C�3��9�g����G�8�@b�:xe[~�=3�V=�s��<��V��~��8��ڙ��:�M�ڬ���Y��;\oϗ��Զ�-�:�dr}��w�Y��o��p�ӿf�ȿ� ;�o�lW��\���1�=8�<�͋�>�7�;+&�A���2�-��=A�L��V���ED��~����X@�F_��\�F��t;�C?.���oo���(��l�j
�k᛻��Q��+J/`^�F��Gu��B��`�<�K|�z�~������l��r/Z��^쭧��[��T��u����qF��������H^�imv]w�Ô9�ͭ�}q�?|��L�Bz���@'.�萗���:�5��.�y�^��*�5���/�n����MG��WXnt�\4 ��+mYSz����o]�vLc�d��a�o�i+X�P�������39dװW�e�b���G�I����spp��g7�A���L���r)5���Л�BEFK��8��h�f{��'x��0��+HK{���%҄t��Z�g���_fmux�Y9p���lz��`�uvk�)�\��P�}^{=<���gw�ǉ�圯ھ�SH]]�S�Oy��"o�Q�x���<����;̽>+d�͋{6�osד�����G��~[���;�W~�)�����U᳗}=�{����W�;6�گ��tz���7c������f�e��}�!�����m�7yf������O{T��OVS�V�U�6�6�9���n�lr���,���K�=�Zur�V�������k�f�s(�k�mf/C��I811�����1��>��]���3?o��X�׍X@��X����YW<����[�n#�Òb.yw����/_������@��bn�'��IvB��[v�LN��t�w¶���� �l����d��0���w0pU��S:�Vn���~��^x�R�m��`�[b�uܮ���ۥ��gW�m���mj�_B�a�l|��s2�u��kQ8��gF&�R�ټd ��������C�0]�E�É��o\}�	�`�:vy�����/�=���.���8R���w����Hsc�8���
�	����)py���<�����1Oȗ�B�X뿠o~��Ӑ���M�|#���$�����8���=,Қ,���K��ф�w����L}�x���4�]�<����I\�Kc�T�f�9)o�=ކ�=��Y�_|僒ߦ����JpڷW ��vi��lXQ����+M��g���e���Hs3�ط��d���1z|�&v�F}�u�Nг'T�yXi�o�LU1�k����t��K1ߌ���;�?|�	��w��]̎��;4rl����"y,��{�EO���������P2���і2{�N[�Ǐ0�m9=��i�%�
���}ٿG�w�{�UCm��2[;�#%D-�槨������ܥ�5W'm.���fN�����햛�lBͽH�F�G_@/9l˂�\K׷��W�����Jgg3+ �1@ �n�V�Gcc�^.�WIl�3�L�3[��c�"_b.��eո���IZ�ēcm�r��a��B��ˍ��/�P�M���j�+^�6��
C�d��觽����p.�`,� *���~g��:��������U1������N�&�E�a�3�?t*��P+�/��[�˝[S;r�}��]O#һ��qY��������~����7���W��|����X�yЙ�z�Pb�|��~���]�iD皯E�|��{up�[�m!��:r�?x~�hb>�3�dܩ�^˯o
-��ݞ�G;J��Q϶���SPϪ%4���g0� �,��ǲ�m��d�f�Q��x*�쑦r��k%�Mw�A��&�Y�'
�Bt��/�����k��M�Vw�O=��1�U�g��If��3�{�����7ٖ�oc5I�{8O���5�5Ǽ�R�Y�}��Kן"��X�o�:�k�x�����-\���z�w�<ί�S��}�x���X��G�K�w7I�R�v�)��X�y;�H�jR�ET[�ϺJ��eA]m᤺Ce�J���F�"!k���L.�j+��G�Z�K���L�����Nt�t)�a��޵�%NXU$��2Q�����[O#�X
�G���a�y�1q�l哕W!��;'�	��u?W��=��'�+Vk�m�]B;���lǙ	LnS{A1��VS(~kiL�<�6����-~'Yo�U����+T���\~�:��C��W�ڪu]�͇���/E]���<
�5���j�}<Y�-��ͨv��OZOc�����>j]���%���CUy��Y0|כ��yi����P�Q�K=\o������&�;�t��y�W�q�}�﻾y}����~J���2?`��a����������f�z�{d�ܢ�9�3��������4gfc�*���ȵ1����h�;��b2<�f��i�P�����v�Q�`������>�N��X��`�6�\�l��+웵��760ƿp��4����1����n9!�}��d�/�c�xx�֥�U-�����oP��+�f�ĹX8y��SY�O�����0��Ʌk|��	�7w[S[�Fθ6c[H|2����ú��a����\̈́��yz����W|�I�R̡�C�oe�{�%�{cV������խ�w w:sø�5�����,\�G}�M�%�<�4�˸w��e��9m�2�-�����r=�HǶ�'2ںÔ����Z��ۖ��<�[�6���t�Ogb�cb���/mK�ø30hqø陷���Z�rQ�z7S��K�;�8�͕�jeMZk�WN��)[�!8*7��K�j��{���Oh���N��*����QV������BYLR5Վ󴨥hfE&,1�k����A�a�d*��u a�
<�������a3�&��yIu	�eۧsL��Fc�E;��Pwe����掲�m�)l�7��N�ă<����*���֙�Ev�x�%�N�s��{�v�aŖ���om�zd�tsGi�\\�M���,�3��B9�ᨡf��z'�O�N�C$=N�Q�xn��Qr�w䐀I�hasee,$����3�s��*]�M��+WI�ݧ{�'0���f������kݫЋĥ�:�j«�?���j]�cݦNin�'��k��/l��K��d;IY�;].w��\���h�
�X�Tv7ԥ��Q�:_<|Ժ�5����&��ĩL�:�(�,rӱ��5��Cf���V⭷c
a붺����W�	6���2�$��FR�P(��y�vKm��1r��U�}C+�U�7�kU_����i@�oiG}G�*ĕ�W ���*ܧ}�L4� �fE��xx�ت;�m���|���Y�Տ���Y�Ӄ�SL�������5�1�u�ʄs�E��FJ�V짤���U��`R6G]�RA��k���Ws-�n���	������oO{��xR��+k��}9>��/��nQ'w:�̅��;BX9���C�cĭ�_�:y��2�ou�cs�\�kjÐŶd�r�U�u2r�y_�8
�]�}MӤ�Oy�p![�+/��7�խ����]��uT��Ma1L��[�O�"���W���S�늻��y����(J�n�M6ʏ.wA�q�U�q=++ m�� �}�Eq�_^#+���%�����R$�r�WAm��\6��A7�b�	�:f�/�i\�fQ��c
�ݞ.+b��Ν yJ�Tс�םxc�f*<��,: KGcd�5wn�*ҵN��%�j��<�}�������*Aۮ�ot
宷f'���GB(��b�6�&o1f���ӵ/
���^}�A�m�;>]Y��U��3Xo��qUӲ߸{��0k�H!��CxkMCY|ZO�,��jf�ϕ���F�@k����/�:�p�l���P��̲r��flA��ra���Ѕ֍��G�*���m�ll�bђ�j3���y�1o��p1�[Fϭ��c�ڈ��M�GW.\��������~=��������?Gϧ�-�F6rA��iرlDjf
B�QZ-�DV�QmmZu�Z55V��������~>=�������_��϶h���EBceל5Rq�b|٣���.�+���"�֘�lQEDLz�"����N���� ����cQ4�����͚�'�I������y���>\���䮚���)���(h�G�<�$���
"�JR���
�����>�*�`�
""n����#3AL�{�)<�DHU4�LEUD���2I��G6H�������h��+�iJ��Dh"
~Y��(��:f�d�E�h�UPE5TQKT1T�G���E%U5KE4T�h�UR{�AS <���L�i]�c3�����ln�µdN.A3�"	ΚY6+�U�� �r��EA�bE`�J����������/i�D�e�u�����ckX~�N���~���/:�s�ѐ�'3C�lmሌo�oa�jd=�P�hJ1����f�#;o�Gq�v�^|ųIi'�6��^3U	�^_MtQ�L�Uc'i!��ܳ3�����>O�y��ey�dϹ�י CH�i�h�$6�2�1�^�ͱ0A��U6y��d����+�/\�謁�'\	����Ŀ���6�?j��{o�#tj�k"ho)��/{7;���U3:��f���U M�q�v1E�D���e����z�e٦�^E�H�Qz�.s2����G��6�}��`>m�bY�q��
�Q�\3
X�{&����в�>�s�0�C[����={7���!��غă#^���u�ˠ
O��i�7)�4��͊�B��'��s�F�D9C��Σ�Ɯ����K����E�XH�I�:$��Ģ��]>��Ul5�rr]��pY;\ua��<��{������`'����Do�h\s5�s;og���ĸM➼1L�~�-|]��V�VLܭ��-��{���O��a ����P����nl�4�t�H��+��� 4�����ٵZ�_��l�엶�f�)�\ǈ0*A�c���l[ۣ/o��,淘�u�9�����O�BV���G��Y��ܺ��U��''k��6r������o�e�CFN[w�n
��R��?"Cʜ����kS�T���O����rc�y��%xV�yy'�7��g�����U�<�;�3�����U/�	y��0#��M���[7T��bg9�!�p��,��cGe���Px=8@kvcl	籢c�x��a�Ob�J�uΩ�/��y����̇���I�}R+OҘga�g��Z���r�9��=W�=C��?L@�1��.;aLmO���e[���}����|%�/��Ǥ�@���~q��υ����;0�p���9�-��3ٔ'����&��X���� �$�mB�bͶV?�,��k���;�n�3�2����{N��K����t��|<�(LS�>yo��#���F�W�p@��	�dfO��b�+Ͱt��6.�X,:Ɉ����:�7ú�Z��S9p+�]��15��O��g�W�]�&
����m����[�M{5�v�с6���ɟ��}�?3k��ӌ�>YP�'&��z���j���v�� ���s���.��f�ZԿ]���~�7�jFڈ����ɽ-��0���h>[����Cl�����vb�S��3��n�j�ީ�#���6�A��f��V��^����˞��}��'5E��v���.Sg{�E�m]TQ��R��y�y�I�F��7dNM����|�Ǚ}f�.��Z��k�=��-��fSX<�ñN�z�=����}SsU��i�"�"���h���g3-��x�V�����[P]O�Q4�K����
��Y�i�Ď��C-�E3}0�3M/.!�jD8���y��z|�b��y}�����IP�w���K��W-�#��#�h��{�˜
��l��M��VӬ�C�^J�n�M���r��f!��r7d=fӳX! [h�
h4X�=|�`x�Q�����3����/[j���IY�;�oF�+ښ�\��뇣�bsf�݂��@A���d��	`f�<���0ΌoWK!��z����y�$��]Q�̎��yӢ��w�r��,�Y�����A�5�h��5\�eF�=u�z��o
Ԧ)�EIe�� p�d�Wy��П��������th����*o��3C��[(&fqVP~=[�*��W�0,a�@k�\�������	� 5�|:)�
����eԛ��Ŧ�}(LC��
����A�u4Vʞ�~�����j=��`�,$-j�����+w�.HZ8@��'�7��͋����`��s��t�^B���>�ԩ�R^�
��渹E�U�h=�UF_��Cy7��!��|�C6�-�0��wa���1l(53��Z}-FB>����}��ƇeЋp2���oj7�-7���`�f��=�q�w��q=�t�x��﯈ߠ�8��]pe�g?D	�3m�\�^�y�k	�ј��d��s�$�Ư^����ԤѬ.�lĤ'�R��9ս(単�~�ϴ�ANCq�պ�Ӭ��&6�W\�%��
ǹ�(8a<�K8sfP���`�t;e���Q����C������&*�x<�k%cs|. w8;���A�- ?���>���<���W��o�hR���z�M;5�S'86���*3J��-�"��H�c��2}�!��}�����F�}M���y(�z�����NE�:�:��xC�qG�zk�8����ɐ��[�����&��4\�k
�p�Ի#'r{�,��Ed����O�g��x����������g�i���"�D۳�A����*8�����}�e6��Ia%f�_zY��R�P
�q#ŧzUc^�Nc����Ě�C�_��v�����P�ʈx�'!���"��Jv��H;t�s��2z� �c�d��M�כW��6[U>.w}Ʃ�x��y��[в�P��p�5nG��c:���C�L�W;�1��[���� �ZvCϣ~w��y-��n� �۪��-s�T�>� �[L��;6�.e:[#%m�wUQ/��̄��ʲk&<��R���%=�E��j�9��T�~k�|F�0w^>�ܬ,�O!�n*}��G�G�fS�Xp��@dK)� ��/"8���D���_���$������|����*�y�����V��,$�}�Ka�B�4����Y��J7[�K.��ײ��+'�3�r�[��q{&�vhu/�� 2�h�j�`�.�ƻMӬ�\iݤzq޸l�37��fM���x�]��� �� �������ɺa!���o;Ctx`�Λ�G�D����{*C����ͼ#�V��1��u*���8���{Jr��[G@�u�]��`3oK���%��e=y������w�����]�3����?�i�5Y�֣hz�E���Y�U�j�R1�0���[��XH�謁"���O0��\�D��Za�q�i���=���B�icq�F�0�~vGD�ޘtN�z<�?�~��R�k/G7=|Kߞ�������_�A.�:-=nܾ��2��������0WI��-!���������k�ݚM�������/� N)M^����/@c�e�v�����)ۯ�cÛh��bJ�N3E�n��W��j({nb1�&.Y�K�!��\?���:Ϭ{F]�ˉ��"�?0��<U�����W��Fo	%7�	����b�mK�ǧ.��S ������h���
��_��~�4�� ��b�qgdn_^����#׻o(�CHmz�sC4��ƴ���ѦI�2�1O��Aj~��Qv#�Tk[�꠾�\ɮ�#k:�T@[��`�M^Yɲ�[T�eO���Ʃ�xi�DO�� ƅU�ՠſF5�߮��1��������J[<�t�	�P����P�44G�K�0~Ӵ��Đ��P'�B���9\����g5�+�Kc{�_�|�|4�s��0��h��"���*�:oD<x4q��o�K*v�^b���x����p��g����wηk뭮~_�����f$�߷��t_E7�u��M�T��Qc �cF��&ꘛ	�Jl�w������u9�O��ԟA���A�?y(�䮑G�q^0���酛�B��!;����ap.j��e ly����G���F�_\�Ց���}����vEE��/��wf��m=SJ6�c��,����-׹vP6$�C	 ���@�	w�*����h��]�/{�e�Ő�λ�c=\*ɫ{�\ޝ=FS��2��W�������i�4���=Fܩ�?*��y��x*T]T][�7c)lr�q���=W�%�=����9e�1�X]�x�;`h-|�ϼ�9��\6L_Cқ� �oH�+��<�D��i��S����G�Uy��dx�{T��2�O�r�
m��>�;����?Ѣ��{I�W��(L2��#��t6HݎE�<T��Ƶ��L����ve��L),8����{0a�7����$C����:�5��27U�纜5����}=%��.�\\̮���{�
m�yE=��2�#?�������:���[��`�}���E�7�3��T����9Qf]e9��Z�mv\���!��R_h������!:�$��t�a�h��Yu�O��{LeN��ZW��.6�z����%c;���)Y��Ž��Y��wV2w�X8�m���FC$�6q��e;��ܵs<$��{o��=�v
�Q�ׄ|7Ú�9k���s���?�۔9q�{�o{�Ҳ�IW
a�<u��n�荂��@/:(���io�'�MG<����&����?�ܵ敄�1b��u
l��m7� �Tf���Y�
0���d�\��Kk�brz��Z��9��_|_r��f��������@��3.�!���K>���p�!�xiꇿd�@�p�m�=����Te��.d<w�j��c���:ـ-�uʮ��s��+�����|VP��ʱ�5}�@t�����'��3OY���9��=��r���׶$Us�1P�8�t(3_�5�Zj��9K.Z�cS��v�\��E2������š�*>��n�h��i��.y�G�M)#�}]B��dP�3Y����/��x��F�՛�~'ke�-al(>@��e��eےg�v|�R٠ö �[d`���깎�AD�.s����%>�F�n�3�1^��r��3���t�s��.���n�U]�O[�1��6֕ka�v���b��QRK��m����@�J����y�6�L
-9�ݥ�!�,)�l���%��(о0a�Q�Z��+�,�<3!��i�vsi! �ʧG�n�?���V�b
_�C��3�=<��vvK����2l5��P��1�b��������mm�nҤ��T���a������7�L[W�+=� ��6f�&J�;0�Q�q�yE�t@1(�lJ��H�WY7�n�H�+{l�F�o_=��w�ʈt�&s�
(P ۅv��d�;�_LAr���j=�w���/��:|�➧eI`�2_��4�����1�޹�����;2dA� S �弬H����.mx���Һ{�����[Y�O�D�~w�b��-���ʊ߶��r��[��AN�$��8�L*�_W��2cBTߵ�m�؞��f�q�h�S �vDW?��Q�t9O3����j痚:�_z&��d����ں-<���V$��M�aA�={է�k@Ϲ;P���0�mȚ�=M��q��-5�v9�Z�X�򵠺o h�F\Z5�#U۸�:��6�����t�jh�QA�6����l9�J��i؜sh�Û�������Py'i�Kڧ�6'�ٓ �������b���l�m�?@��jN�x`j��0gy^�;U�����������k��/5c����cn�	���,����th�|�_�|=<�����M�v=�V��t"`���p���{��]q>-:eV1�^W7��2��l�C�z�f���7��3[7��Y�*��K��Q�V�bn�3p(CN^�n��9	�v� 37���Վ�la ���j����̋r�'�KSL�r�'6������|��Z����tw�V�v�}9�'�1�K,����d�GKy՛�/*#y��2���;��3�?N慜$�be�{�Y����޼� �J3�r
g9 t�� <�=�xy�Y�K�]�C�Q ���aK�K.*e����n���
��WnU8+:�����Н:����9��F��0��u�t��{���s���L3�C{D���g)�b���n-l��!��F�ŧ�Q����$`t��v-5��bh=q�E�yS*
ɜ/��O��+8&j�J�����zwt�d��,�S:v��_�w|8%�8ý�Ȑ�ח<=B��*�=��_W^N�sY]J\c,�U��ܖ���C�v�㢣
�)r,���P�� m�w�gr��4k���1�˳���v��55��.(��r��!
Jֹv�0��<xhh��,d'�34�0``�x����k�+6�i���=oq��j���Anʵ^f7EW1���PP���D@ր��_��l.&�8�t�\¡Le����QM�Sږp�D6�A��8ϳ���b}c�K9�>^�q�K�1�DP. [ʤK�E"��qy`����}�;c���/Xs#[����u�3E��Pga"��a�3<�P�����oY$l#>��r>�d���=�N{�h#���'������ 6*�ڷ�%rש�7���[O|�{LU���ù��VfL�j���릓��c����+��Ի5�$�7��]T�n����q5�Wz���|����p�O`�n��G�k�x7����c�(�[r1l��W�5�ϙ����W��_*����
"��0��B�C��5�� �+},�ߛ��C=���3藱�Ss����D��i9�ګ�ae�3Y[�;�1CPj[�Cp��kz����̓�K�aZ��蚏uP����5=W�*uApxه���{q���HF'TpWK��lW$�3�m�ʒ�*f(����mD%.����t$�����:
�-3m�s��T����#+�ȵ��Q�\E�O�x&��8�Os[�M�v�z	>3F|0&j��eL���漢��j�{8��Ʃ���;J�:(Tj�e�r�1}�op������@�r.�����{�A.��/�E�'P�.aބ���}��s���97�̆��+��-���ca�иG���ɧ��gAZ��WbYr��|��SZ;/�5YQ�9��z��>b�As��P���O�-[�$C�����Z0�\!;�o�O,�Q�J�>�]�ݖ9�b���MC%PK���4�w��5��˲����K���C��>���b����B�f7Z�Y�}Þh�E@������(:;�cl��s�X0,��[$�3a!��#����6�d�3�Q:�������+��h��������؛S%�&�R[4��772[�͎N쩅$��C�v�+����Qu��,����.qb���%��֭���]N�R��Onm�*h�`xEp��u&Mю�HpA��K��dt��\��J�]��;7�	C52�ٰ����
Us��]g�o�#.>2Q�kV���p�汜����%8CCat�Q�ec6�=rs_Y���<�RT��*ݥy{�cޥJ���$2'�6ü����
&B�oU��E��\�k�U`�=
��uBݲfk�g^����y�.���b�)Ǫo[�X ��N�8����p��2�'����!���+qWK����+e��^��J�or(����9�>x�	f���������	�"��J;p6u��$�<�� :��FΉ�]	����n;�̳j�[z.`Ţ�I�K�`3kB��y��(��:����u��ӝ�X�Ǯ�(�ӫ�6�id$�[��4)��,�V�V;��.��i���PSEaF�"R��H�X������Tq�Y��B/���l>M�ŘK
�4�XpA߷�T���"|r*R]\�DW*�ң2������-%��.�SYj����f�:��b�u䲅d�����\x8�QUs�eJ�'�v6�0�ꙹ�N���;%�{����f����M(ZE�7�ԎV=��Rj)}�
��vn\�r����i�]�l�*,��Z7�vL�[ a���lzXt�h0��Z�H��z�T��2�D91T7�RB������ÀT3J�&WK���e�>qB6����N�Ӛ�Quڽ�x���h;X�m�][H�*�E���n���Y���'��s����bMը�Bki�VN͜I-��/7�c# �it�Yu�٠Ý�.�Yױ��M��&h.��M����[V�ނ��M�}1�;|���s��e�7Ի��^e�.g]�o&�oד�,e��2șS���9�u�8�]�S�N���x,����e�-���E�UĻ�ʜ+Mڕ��նE���oJ���s�S���H�h8����u+�(f�T��o��:ŭ�a�sp��d�1N�i` 3�».����^��qVذ��ؼ��[l�^*��ᝨ���A_,ň��S#Ļ�eҧ����[9�یvs��x�aɀ�T�Xk��)s�M*�wY�O3q�;��"�a��v>�[u�Lݷ��+MFX%ZFb$��c)n�ZvP���%���=Vr\��!��,�Btv����[Y�$bB�̚�'����P�p��rIġ3����fǎ��e,0mvZ+�Fsn�;R���@ 4��,̥���B���:�N�^c$�vä:|5���t�z	,vМ�Z4 �����xG��2w�7��[i����	����̆�s��"񽗼�2�=]f���d���&/����_8�,�1d�`���+�X��f>��<�jj=����[��2Is]���d��e�Ra�� 0L�UK�U*T�-�Nb0��g�	�Z1�Hh��ߏ�$JSH��IP1k@L������۟�����������������~��3��h�
bhi��"�T���hy�)���Ϗ���Ƿ�����������~��(�d�h�������������	TE�4R�u�u�321Q@]4TKT�MTCDCE%kIB�E�4�5�T�T��ǽ��(fbNK���(
/���4�1AM5TT�P�TD�D7,PSQHQKd�CAUUAAK5HQASEp���MRTMH�G�IUE�+CAAE7{DEQO{D���S)��#M:w3��ZF�F�Jyh�ƙ�����(K�5ICL�R/V��z���s�:�/\��V���n[�AKz;�vI�Z,
�[
n���J�� m sy7\}]i�>n��M�4="=�	�\Tnv�֏n���}��"�(q2d��P:���Px�"��DP}�}�w��D(���y���S��*��K���[)��4ic��j�ݎdC6�>�<��꘥7;@L5��-.;V='��#h�J<6
41��H|�S8Ckq�O��"/�Na�Qs���C�܂�N4�`���!��=>���Z����hw1��A'[�ʴ6e=��9;}K~�;��V�_���#�P��R`�a'bϏZ<f�ʜT��oN\��D9�g�Z1�k/�r��ϒ�)�%Q�Yy�_*����r�}4�<=�>��0�;����M��35��'���#����}LZ|��g�= �ÃZ����m���SQ�1^��m�m���5��v��/�R��-��.�*Ή���1����6��vqQ�L�J�\WK�=�*�8׳o}��z��Q�^(12)ߤ���B��s�F%+^�l �^��O��r'hj�"b�|���v��x٥�3j�,[���St��l]��|q�'� ���P�(,4�#v�����U;nD�C�#Y�/M�0�we���<}z�Ĺ�P�+Ң��	|��h���k��:iPI�.��ڠ��ݥ]K8�M�ȗR�4�|�z[HǸ�c�dտ���OP�t��y�[�S�$���ѼZ�G����ûe�q��#�ih���v5V�j*�SsPExj"�6t=R[ŸT ǗһPۘ�m��u���:lͷ�������/?����?�����QDڈ�������-��FT�hë' ��{�C6y��d�||�!?V@!�+��s�h���%��f[V���)��_��1���+��&.���t].�Aiv��ª1�)f}0�2�9��u���Q@g8v�
ޘC�F���S�k�Ֆ�O��y��M��.ۜUR�2mT���N1A|-� �Ǝ|��4.����6��n��Q���'�O�����J�0���L����q��c�ه|:%�Cg������B�iTa�n�������	|o�i�ӝO�/&��w����&�&
:�.�ᡀ��O�]�#���>GFno+mu�I�%65Ƴ��Q;�ofl����ٕk�5@z����</ʇ��`�k������@}k깦I�Ч�U�nT�+o��<�����
���D?�覗9��#�U�FRk�o��ϕeޛ��h+��6�l60��]�g$k�p3��޲'�&xg��!ʟ7<�	�*�����i�����&@X℁Y+��uw�ۯ����r������\ )�<����J�Q�g;S<�B����~��*�h�c�ZE�3���6+���O7w/��Tzh4�e�<N����������|��ʢ�+Z8�[w�e�X���{�����9+Yѩ��2����7�	\f���_k��V�k�۴�:\ʵ9��ņ��=�����\���A��|��κߏ_�_.\�9��� k>�+����n��{7d���~���%��ۇ�}H�Z��x�\f:�t�'��v͠�-��R�=��~��EJ�
k:da��t5�:���j�6f�]d�Mkz�V>��4M�ބ���.�_�|�viq���p�ol(��
�G::�|/�y[�_���M�({%*�j�Y.慒��T@� ��eC����YY1���t�����{U�(tBe�L�k�F���yu��΢�݅�P����5��*�0o��&��c�h�!�4�羈�酋d��PؾJ��z��ο<��Q�W%�Z_r��w-f�x᭩�j��PF��gM�@ML��2��򧋗y/����ݥ���`Ӟ`�U�}�C{Lk�,��Bv֖w�As��~Zx�]�����p@��2�;�u�(��F��(���۩-����{Z�=��~wx�l��+�SK�h&Fm��D^�� O:|`��2�+���t����@%ܶ0B�g�n#�����@��>��s�?����j����C6Em�^R�`��G%��ꎽ���_;[��]\D��|�\\x1/7�Q�Zb�v�g)�єˮ�Gb�x�4M�TU��m�l�5�s�7:8q�XtB��:-d{N�����{.����![�2@Z�1�"���=��C���a�> {�=�� =���� ��9�Bj)�isc91-�zKoڣ���>�a�S���i�:y�K�`��cS�>a-�F�K^F��OE3Ay����j~�)�<�O���pb}Zj�����y%j>+޼{=�����!���)�>���+_�1�|e���c�^�X�����:��� �\y��1�wt�?>(`C$�Fh ]tDu�	hq�F�;���Gu�<�՞�m���z'MV'���5Fs����׏4X��>�M��iq��x6:�����V�~涜,��ok/S����+��20��XY�]?�r���15E�Q���^�r��� ����<CRfڞ�i��p��r�2˟�$]6+�їw��$����L(jŃZ����S}��v�Ԧ��sR:��U���2c�o�Y23UF	�Z�r��N5�:li¨�h[ѭXk��(b� �h��v>�nh;+m/�e�^QZV�G�@��QVjm{6^f����;v�L��m1�i�"��A-o��1?amc�ұ��ӓ����^�^��뛗��8n?�����_�_�I)K�r�goS�_�1�J�I��s���������᱋���9S�1K�Ba�*t�锹���Ôg�I\�t����6D����,�;:�eap�|Y��&]u��������p���dRL���~EG?�
�s�QO���������߮bj��p���!��*��NLc׎ǲ���S4r���r��:���<�J\h�c;�Zk���;*1]o\�K(u��ǜW``7�:��:5��O�����A��� ��
�6Q����~6�����2�]�=ˣ���R9`�L]߃9`ZC�=���K�^\�O�Dk*Y�5�2���;�a���Q�:յ�.�-�G�Xy��#	�m�-(�V�\��ֽ��ڠ2x}FZ#�Կ�t��h�Q����AF}K#Ɯj.�x���vN�k�Z��nZ��K~���N��tx'Є�Ak���Xi�����ԓ�F���~n�t��Xy�M)�o��^�����;�x�x�	��������?�ժ�;�����,�ƞ��Y
�ؙ���ΰʎ5p�^S�s���0�?��a�U����NS�=@����]��*jq�����ג�ƶ�<M�tL!�*��y�gL�,\MG<ñ>�Co�l�"X�o_q��,F���=]]@�;��$���@BC�$��n;o��}m2MR���;()bh}�
�j�Cm����,ޫ`KD����[@�K�s9��6R����YJ���ы�>?�߭W�%E�*�
����6/����j���vse�L�t���Pe��.ӛg��A[Y\�>��N�K�S������� 7�y� �?��<�5����qz�K�8��w��U����d�0���&��90�(��Y�
7P���"6[i�����Q�K�ܨ���k߬v���V��YB�f�� mU�Mk�~'�[	���fܨq�O`�L"}���G#W�����!c8���<(�z�1�|<�7۽3�}$��be7����8����nF)b�<�Ψ�BLZ٨�Ң��r��ND�WQ��__��b��߸�J<��e5Y�H�]6_�l��08KH�nԐsf0Y���q�ҩOu�U����{�"�.0�L}�I� �)��`J=����#���[N��>.�:C٪}w�]k������;��j�Z\[�A���B��aC�Jb�<�e�L�n��V8K�^��E��ݨ���9��%V��P��������y�FEP�hÊ��U�,�%���5U�Z��R��U�V^��F��H 5��ه|:'�3
��Ш���4w�zy�e��Ga� ������ܡ� ��6q���A��������=��3�p�<��B�ǚ�t�9�?kT��׵β�-�q�'�J͉R?����w4ۈ젨��=��������u��<��,0E �H�A��3�j܄a�;��}�ۧ��]�F���x��=/MS�Ү�������֥I,�
�K�N����u������*����p)���������!M�W!��S�P��t����q�h/�(���&���(��O��X<rxo�ˋ6,�/�{��ѽ�Qι��(β�)�����_�"��K��딬p��~0�av+��VU��R���*�73�ը��G��X6v���l{��3�P�1�؍����P��s�j��}��乍
﵍ހ�{�0Ɇw�H��&���4,�ܞ.���m�ZG	�Sl��=��D�r� ��+�{���W��ا����c�`�+���3���|ZZ$�1/jެ���ɐ�Y��Y'L3�κͫ�d�V��p��E#Ր��o];	=�b��1�"�"��Q�-�a��lz�P�;��a˨�y���m�lV2���������5��4ڨw7�2M���4"�y�N5���I�\��EJ}�'�mc���d�V5�>��s`-�e�Ng)�i�l[N�����;�&������k�7&��=J��n`���C���
�e��b���y��Q�0(f�R|��;]c��Ĵ���c�c0��L˟��Y�"5Q��]7��0�m�>jQ�t͗��0jHuS��ڕǀ�@il�W}n�#��B4�څɧ��' �$�ȼ��y۽�>*�K����-<kz�Øиܗ��Z!���W�x��rru����/Ӈ�!�O��{X#]�mr��[�V���X܄�n�Yj�쬚�k}��z�^���T���9�UT>�=x7J�R&�qj����1��l��E�!�wi�,Ғ�ъb��t@Qj	�=a��c�bV��<)���;����b!>�=�Ց,d\�,_�_����<�����Ϊ��"��P���f��j6S-��E@-�U�f3I$�;Xe}�z�|Dm�w�gzF�j|������9Ug�ܺCO;YN�\_F�{gNK����}I��n4�(3���4��;A
�k�<����!�qLz�x�G#������8��Ft4�����Ɨ`5�#U��-�����*0��V\{����q�+���J{~hw�P������D��\�AO�Sl�����it����|E~k���9V#���ǝ������=6�,�~N����(��������\Q�4m�8un��3���fB1~��3�h�A�e#�_|���p�2s�{�~B���,I���T�|�� :kM$��Vrf>�xД���d���^AiD�e�({�I�����*ޒ"}�<h.����j]<�zw�C�EB�D5k�Y�-��Vk|o�Ze��O���+Uy`�ڷ8:���i\cN�GD`���|��zYK�ؤ��=����u����b�����TݚE����z���0-	N_[�yD_[Y�!�*���C���V�vlV�?�,�Z;+s�.Ӈ�ć<���V4��7-�� 8�\*�8D ��-����؈���Ægv�a��a�ڦ�^j1-�8<��U�+�їw�2Mq�sq�uHXS>��<��v'-᷉�4t�g��x�"����V�k�ɕ�1��N���,�M���c;�f+������s_�Y�kAu$ny����C�$�߷����S�����[s�鍃l��k^i�OEe>�^�r6�?�����ɷ���8������n3y��s>��N���m\*��@ȭ�F��5ݓ"�=��e���=��?-��ྞgi0SRXv��t�G�cWz���=��l���^i��nD6.�|�[��ʠ��A�&�iw*1�6b��tVU��
�d₮�"�^��mB⮓��iO^�|�[�]��L`?�8�G�����BE�ݕR�EN���9Լ�u"S͘ս��)�9F,^s>����X�5۰��<������兟	�y����y���A��:s4��CL��VXvlsbz���=��qe�1-�LC��ط��a\# �y������`8O��g.�Aj��3X='�du13���F�9���l�]˩m����X�0�G|�ҫ���-��z��IeM'�f��]*�����i�^�\M�yo	�ҳWw��ӌa�̞X�(W3�6$�6�\G�>`�A�g�����+�:\j����Bp�y�^�i�b�����:�߯ʀg��W9� ?9���ã�k�Ls��pOk�G�a�ؐ-��$CQ�a����_G�7{��˲ ���9�Wv�si�\O!�6·z�<�(?J�<�G�\�[⁭h����W�:b�t��++���]m��1��!r�f҆��W�w掂)�z��@q�S�/.���u��u��"�8<��"n(���X��1���V�.�Y�K8���w�!*�TS�,���2��ꥁ~�Bh�9V79_v������4<���Y�0�����^�*m�dKe-�rwB���b��F8�*st������i&�]��_h�0+­J���aϩE''�U���9�K�.�_&�>}C�?S��~g�i�]�*�y�t��?Q�x)�j��AB��kY�T��N��Wz_6g*�h�*�Eq��T4ܥ7Ū��]8k�zΧ�l�-lY����z)��T���+�ľ~�XFܹ���&���%9*<���ؼ{Ur7G-����q-�p aR�������ં�a3JXV�`��<L�4l- �N��Sv�J=�H卽�[�!���@,�~�v�q&~ӹ�.B�6��Ռ5 �s��*}D�+���K0�M�s^����N4�;R�>3:m��.��[#?	�\.���YF-�8E6�S�7��:�������Ǌl),�����9���S���En�V"'Ni*f�v�� Hδ.u.��ry�p��G+�۹-��%��ykop�#/� %
���z�q��սl�E35K�g[�5f\�����j�4'ܔ�a�1�Lr"������L��)/	�6J*֕��s��j����}�u�yDBvؘ05��s/���M�ÑX����c},������ʘ�a�
��R�Ҷ���cH�Ur��N8[o�t����F��d�v�e�u��K���mݩ��6���� w:�bn�{�.[�u��Nwq��ļx��-r��w��������a�$X}s�N�!��:��ign��> 8���K���p*TM	����/%tZ1fސ� ����m3Zud�V!�R���[��1_dt�p�r�ys�HtB��T���}w�W7�K�q.�v�lE�\�[#-��I��[}וwEp�`t����'�������x&!���U�Ajwf.T�+-m��)�l<9���.�M�u�݅�ugR��t���nV�2Ա���������Vذ��J��0��19%�����#���k����t��Y�q{)C���޽'Z����Y\�s4�8UKRu<�dW�J���Vz���ԛ�a:���s�=�5���@3���q��'���f��?��ܮǆ�:�[��`7{6�%���wJ�v�ʘ���i���/��v�A\�E�}*K<�솱�2�u�D>�*Ԭ،��[�*Nֆl!����Vc�ܠ�o{�ɱ��X� ��E��Լŝ��fD;mŨYkujs�.�:|�m�Oz�Mz1�.��#N^��4��W�ގ�[P�8�B�z7nN��wc�o3��f+i��Z[&X9j{oq>85���MnS��O���$���HfZ�t����4�#h@\�n�^M[�Ph�ʀ�gqy�m�sA�x�Ӱ^X,��#�B�4hkI�>! Mˬe��+pu$�]z�qqT�J
����_4$��7doa�핓x��T��D���8��\.Z���A�a�p^;����C���8E�]�z�e#/�,���;>�c��|[���t�2Lq�{x��]�jZ�r�n[6��N=s��ެ��y��D1���F��dT��P_-�&�E��J
�r� 6��l��޷}%*��U�6M�3!�SY]1A�ʸμ��E^4�s�����P�ϛ�z�Z8�ƣzLNn�r	��#;���V	I�^.��u��x�o_j�|�����N���f�Pk9ɶ[*��Ϳ��]��_��U��Đy�<���M|�!AO�<}=���ߏ�oooooo����P7̘�Z���奪��}��	��SIǏ����������{{{{{~�_����'dz�����AJP�A�M4)@��EDQE�As&#��*R��:���")� Ѥ�"��.��'[u���4�)��w��}N�z�Hr �2�kԼ�T&�o\��^�z/Q�9��:�^\��Bi��U�M��r4s[��4�%']`9uU�C�$
9&&����kE���E~���4ޱl�|^c��G��� �i��#O*(��O�O#c%�k�1)�a�d�V��9QEU�HQOW�QW̔�)ʊ=AG#���:)��+'+[w�Kno��y��5�}r��]�S�S6�����nH�إ�E�����d`?xҫҗuu�w�-��������*WP�Q7�U���&s�7�ߣ��w�z�q����?��>4�Y2E_L/�a1Oj*y�`ͩB�[:�B�-�I�)��"��� �
٠���vCx�Y�1K��Eq���K+���H�g˥q9f��s�k|�k��S�(N'��� #o��$=�Dz!��mX��sT��;�>�w�ۨ\�X�C��{����ŋ,#��a�g�� #�u�+��L�ۜ�Kr^�6�\O̳�`�݃˱R���.�fZ��4� `�o=��-�O�ޜx`N�2�·xR��ܝ�Z��dnVb��^�H�-���d�kg�:N�q�F��:*ה�@x��;��	�-h��S�M#y��}�N`E]��z�8Ǝ�3'���i�����ag�0-�|��	�V;U�I��m���-	��҈���~�w�n�O�����D7�E۞Ø!��i;[2N���k4���p�{�$=�rp�\^~��>���T�y��a�ݐ��q��,��(�//���˭:y���-�ԉ�3p����;i�&8�@��Vi�O2~�G��w���YSN)����ɓ�RIǕ�R��'~뫡R��z���O�f,]4���ٛ�֩l
G�����G\�l��$ś�Y�t�����W/-��7��]1�����*D�󾶔��ꄼvf'׸�c�>^�
_�λ~y݋��v����8����߿57�,"KM��nS)�N5�\������pY0A~P?Y�fDz����Y��/�xC��MX����B}��#��qcתjZW�d���d�2�ݚ��W��̬���G���}�,
�zN�Y ���	��Ϝw��t��<UV��=kb�J��-�����[
��9��P�6�9��ʠ��C���Z�0��c^�W9�1��A�*��ܦ��/X�*$ʵbOK�ۘ1mr���ڧ����F]��	�	��h��4�q�\Y�TS�C�Q��u���ۦ�3#�k�ol�!0���r�y��w�t��N��-��q��jxz
�-Q<��6p�A�L镩�(�ⳓ�nZ�4O ��`�}�y2�,6�;�j#~���K�K��:r�̜RnP���jR�Y���O\���{d��	�2|��'�6K������t�*dd��p%�>�>9�3��-R�kH�3M@��V��9m�j��\�[�L;a�kqŷ�EL<D$9���q�-��q�ʀ���*���1������q�}�����K�u��5�1Z��w>�μ/f�%nwT���w���BH�H�,$r���%�XlV��z���ۛ�i���5���%�r4>��+�w�3T4�ź�4a¤T%�oT�*Gu��A�8'C4�\͜y���Xգ-�Ǐ�t7��g�A*��ܵa����uْ��K�JW�� �c�_���¹�A �^����z�o�~.�KE�gz�	��&"�C�����`P�|�S޻k��oP��1�����݅��	 �m��Ov�ވ�і���Ua�΁DA��sԙ8ϟ�3�G�(T�n�-r�_M��POѡ�@T�5~��w�C��v�'��^�݁A7b�%���ƺ&]���'������N����Zp_�_Z����?;����;Wޱ�颻 i�jJ,6H˰-����ʒߩ15E�Q[Wc'S�ɐ�ϳ����J���Jۛïa���N��j�^��P���'�[��(b�����`��.C��hF�0>��	<�ԷO�dOi� ��B��d�Ī,M�3��8~ئX�>�b'���q��\Xv�16.]C\�`4*$\Ag�!�+f'�ޘEi�B��\w��5.��2�hY[;��m6�L�*�
n���o��m�I�M>���hdph�X6�<��N�e+�J����gx��3�S�ۮ 5r2��NN.V0�6�X���8���ь IM>� �#������n@!����-׈L�gm��������(�nx���,��%ei;�2+���`����ʃ|�%������W(�%��sp�
��*�9N��2��e-�d������7�K���\{A�>�g��a��I^���V�)��r"l87rf�Ef�N*g:���p���tE3�5:�9\���^|������p�s�P�����tmcl����v-=��3�nQt�c����d���`i%���l�*�H��/�xS?H=]��sc�����ف�j��ޞ���M	���[�s?�¡;�N{�9-]I��Vh�C~��$�L����s���3�3��Ȫ�TXm��:{[z NAN��3Ia&�S��q��e�G���|M����tO��i����c��-�aUJc�+��C�q��e��d�c�z��o��r�@ d�;D� ������������^����tWt�9��K�,};�>#��P7�G�K}_�`���"��|��~�[�qW�J}�����g�%�Dds����y�3b�i�'z�	K�`w�`��Y������͵ںGtv��L�����z��=\����\Z44˃��K���W�ͼ�}T��1/�NcL�j�CXhZg�f�P�U?�b�z��6a�rt�HFD�dR�ꪭ��R�OOO�K��8���j~��o���AT���˧֠�艉B�[��(/s3���W!�ᩌ��HQ5�bB��ǖ`<훮J^P��؈��dؓp��=���kt�*�c��!������/kp��I�rr�%�*�R����O�[WI��U�CŁ�UCzE�,�,�.�xX�X#�sP��-���i�BV.�ӋwE-����}��?�� ����V;�%3�WB<��r��s��,4WP\��[�ϳϔa�2��4r3y0GLSy���A\m��biu�Y,�Ǟ��)>�ܡ{iVk��YP�}y-��<�Qb\��e�5��w���C䜽�9K f��c�>FΊmx��\�Z����^�{yClrڍp+���%��e��K�ɒ4$����8���m��v�l��^�2�:`�V�1��O�}Hɾ���]�f��O՟�ܚ�;�̐�}f�|��O�3�{��(/ށA[҃N����y�t����#{eT����|z}���?�c�X��oP�����M��c�<�#B�a�:���ù�iFR�͙mݦ/��Z�F%0��N	�bZ�dlk��FD?#��h�a�=�]9Tk����x��Yw��8�媜�k==�7
��F�o���]��L1����_���T�~^���$d�~�J���ސ���v�(;qV���L�k`��\��!��s�P���ɖB�jC:�b�� =2TV��S������Wy��8�U=S���ft�.S���E���]�F1�j�c|7�7,ե؉t!��b�|{e�� �8D$f;��-m�eI���Oc�t�ɹ����>�o2�s����)ݘ�Si�%�}2����7%���7g}z����]��������r�U]����u>��^�۟XXko���f�k�o���= Lf��QgÑ�v�S�D�ZӇIܗAͦd���G�o�9=7��?|��Co/*=�r��9��w�9Gh��N�4�����G?��_uF���)����,J}圂��ݼ�>�3��C�?y���s�;��L�����-�nX�.�!��9�N�*6�������l��R^!n��Qz����;�"�W�sZP���d2YuKM�lV!��C��2��I�C�Cy8��g`�3�S�t�%�c׆)�)a^-^MV6����٤��1��Uׅ1mD<���90q2�F�{/-�,"+���S�@;��u��@�!�Z��XV��e�
�e�p.�mYSl$Z���-�����+�G���󯪣{s�}��.�'A"�Ÿ,1G�?�v�>)�5�w��S	�Wl�6B�}�g:8E�jC���8��6'�Z�N�g�<��ގgLq�lL��P�6��H��,m���U��=(�)���=���FKr�gE4'ns}v�����8�HñO�rQ�|��⾨��ڮ����ЏnjD�i�3���Nf�=�b�]�ki�s&s��8u�a�gL�>�<���J��A%���xμH�>u�N�T��,�r�\��S)�����`=�t�L�O�ajUҙ������aVWӎ�&-8�](�GtSj&�+�;�+pѿL����:��ދ�_�+�'��`�"/�7��y�Η��%��'�m���\u��Kimi�7��n�����5=��PͲ-�����t��B�B�Q�kƎ��\�ᮞ�>�X��H,#��\�;����Jѥ�֧ �K�a�U�1k=�z#�`��o^�~G�GsJ}~&�Th��0E���fk\<v]��U��F'v��T1�*:�p�4��g��F�>�.�u?=1���gj�<�ѵ9:pE"�r��Z�0�ws�b2���㾲,����a�As#[��u�af�Чk!up܎;��q�(?J��F��qD��x��}��Z_'�k \�u��T�f��Zj� �R޷m��i- �	M�@�T'��.�ş�����̟?|��4���ø�,6�R-%�wC4&��"��a���!�b��i�T�� �X��0�xlZD ��81u��dk>>SQ�6ä-�W�L2x*1}�*�/VS��Zzwq���j[��)�մ)�PNqL���}2-z�;B�!��˚������\�z��!tܲdb�.덼8w��h}���jY��ǀݛ:��![��n⽉�Qjm�qul,�T�N��>�>���Bo��hy���,<�nk���R�T���r_n���3����Kw�%�[�-N�CE9����&ކ��hn�[Z��-�~������Ȼ+b\�]T���L�<4ۆ�w���;�3'; �hCt�K���yEi�`�^����Ϋ�SU��I|^*E6W)�{k�Wo.��O)Ҁ0zl�m���m�ʱ��&�W���E��T�NQ=K\����.�}V��kP''%ο��3�g�nB=~p�M������S�1B�s:-S1�<��wx�5���E�s�P<��K(ts0�|���"�b]��S4�ګ�SZ{7�/L�.4Dũ"}���6�Bү�G�kߜ�d����$��4{ީ�n��i��(�7�_�������a��z2���v>h	]s�����[���9��MM�Vf��6Z"�݀�����I%C4?0�F��PSЗ��^ǩ�+�'@4.�r����F���8<c+��`���{�׫+O�(W����c$�|S ��^5�!�b��<��#I{7��"����Y�k���͗��C���(J�ס�,4�!��$v4�mG	�*�tj6Ú�e%9}%�׮8��t:@�C�1��z�,2�h�/" �����ci���� c��~����	�|�g��:
�i���c+�iPV]-7�v�Nb�w�7�E��g��Z����ө��lT�;̃-I}:��ն�?A�|�I3:̞iz����+�4w]�cåwְ��q��^�z	����PoJ֞�v�ܘ�����}��������h�V��1��	ƻ�fk������L!���,y�gL���K�>�L `/2xX6�_��ѐ�C���4�l���M�׏�O�}̲��3$��F��0�C�A|اEA8���o-K1s�L�!F������QV��}y:a�������.*�Us�i��'�;$���	�Ȝ?�>��_zJK����T<��J׽Mbٕv��XM9�C�\"��ۊ/��(V��X�ܗ���!l��r9��i�l��ˏW
Ƞzp>̵n�Qi�s��Av�ƚ��8�eg�7���S��\��eC�ށ����7^W1�}��w0���Yi@<�`��
y��M&��@�"�u
�dU�2�����&CF��a�:�Mp��Q�L�)r�.�.��k.�5Ss�~%:\�Lu��S�R7c.�<�o<��]�52��t�aכ�F|]�C��`��l�1W�,e�����@�B�s�-*���DX˛u�w{)��1�bV��,t�C��I�=B'��Ǽ�b�����U�FV�f�m��9�`_ёu��H��َ=���q;�3���eCtS��z,��Z2����0�;��6{�:�oW-U���9���twa�	;���k�ӱ�P��
���c݈n�4ږ��2���v;�M�I��O�����x�c��I=�k�7�q��s�'�J֩i�娦K�~xz�����R��/]G�y뻐82�bh$y����sU�q��ޭO^� w8�Ia#�Z�����6�8�ǈ&���*c�w�mG��+��ǖ�l�A��ڭ8��#�
�{7G�Se�(�o4���S3^8+y�?�oG���W����}�g���6���I���𭖨��5�:�����c��3���&���F{3�a�a�b%�_�pߝ��|���}�}3ʢ?-"XVz_�5�~[`��w��Y�u�W{2!�1��S�l�����Kf�y�S������r߾\+Y�'�Ƌ���K�}`����=��7��/�5���7��3�(����G�$���� k>��
�~ǹ6'_��g����l�)��Z�BT��{��A�7K�!��F��H�l4���hO�ߨ١Z��;5�s8&=�)�s���5M=JBbUH�|�*�}�ڃ�%� ��,ͫ�W����"��߆�m�6��=��s&�Z���c_�N�r�>�G}ӭ퐺͋�YS���o��5��7\��g7w[�VWc�����m��$�\��ُ��#K*r2����C����ǭk0Ί"�*�+��c��l��}/E��_u���[�M�W�u�	����)���&pW���R���t�w�Jr[z�� ��gfu>ͺ"��4��k]��sM���-���˝��l�Z�ŀ��(~���)�d��zF����@ aJ��r]:�QX���{�E�vsٖ;9��˶�*a­�C�HT0-���%�ǡ��q��-��+$��ز�r�V�2�\N�X���<r��S�eEW����D& ���ZT�����f�H���X��%gV����]����	6n��T��Ú�kU.�&����p�u�=6��q�D�ԦoG�� �&�ͼ�T�Q���ukl��o0]s�jW]4[�\�G09�LȊR���O}K����S	u-!���q%�ի�1ַ:��'/�v��e[םBm*ZG;����8�b�\h�5x��1�k�w��՜=��]���"o���>Ӧ����o��ȫBy������
1���{}��ɤv���tR��b�j�e;��Whuc�� �LX����&�H�w9v�=zn�:� �B�g&�U��j�yk0=�:��*M�8m��{���۶���K
��N�5�൙R�B�e
Se�g)�NY�Lǹ��T���������ێ�/I2�ʂ)
�Þ�-v\V��"�ٹ��d]%W�6Z�ֿ2�k,G�m/��9V�m����������ˎr�Gj���h1�K9]'VL���7p+�T�ok�9s\��صK��Mɕ�O].vݮD��8/�i9yIS�E��Yl^+@�3���{�+(X��L{�; WRLn�[V�1��NR�y���%�Q�ƹs�=�k�e-���Ž��n�ii�Q>
c���n˻dv_ˍ��H�-�;e:i9[�h�ݩ����I�r;��;�ZK�E)Z������ڜ��� �v�=6a�}�j�Sțz:�fјGql��]R���чi䥂�-F�e�~��^�I�1J^�o	]R�3Z�}�&y���(��fٵ�W}�P2�p�>j������ Aˇ�aR�r��\��H[.7K�k�:�f�z1�25/��ފɽ�K����'X(�gy��"��5��ϗt�����]p:UյnF�cfS��oKU[��9�J ��L��l*�X�;��J��R�tZ��"{+�۳SU����� �op�8y�zO4[�eY��6�:aӚTk��.We�
�M�9O�R��&�n��n��®�:ɶ�V�v��vB�n��|��XnΌ�������!s~��c	�˽���*��߂���m�3�$V�23�:��c�Rh�wC)�'����d��o��Q�X��иk1�{z�}�,c:�Y��\�,ܝ[�b%7�����(n0�0�")D�A�J$�d�j�M�[[hdm�c����NIl������A?��堤��:��</^��]{�S�h�J9�˒�a45��x��}>ߏ�oo��������~�ZZZ��p��������Զ�G�9ʂ����z�u����z|}>ߏ�ooo׷�������}�TW�Ѷ�d�)�'���h:���z�i�z��G^��Z)�����Ͷ�(޸k��4�u�GSAT��#OQ�3l��s-���P�=$��S�OS��WRm��s��w��?->����tr�#��
8s{�GD�F�Z֋�t��55\�|�\���i�m'�9-z�8Z"����\��Iͨ�[u�WV�uuS�KHr�As<�%�S�X��M	�Ԛk�]A�kr.��S��I���#M��F��#��'�0ST{m'w�cݨ���h)֞��H�$Q?�6 �d4�a%�f��#��3���k�7Dѡi�㝰ZNa�k���A��`�&���\#{�f��1�6_"�V��Y�M8�0�!p"�	�*$������~?��xs�RP %{��{���4���x,$��犪e�qt�h�MG�B�s-C�!��U0�z���!�F���H��;X\e�� ��Sm���f%���t領���h%�\�g)7{�V-顲���{�~���k�{�с@��"������w?����(���[��d�-'��p�c��Q��/`i�m��c�X� ��t
��<xȈ����a�]Էb��Q�77]�1bq}�oE�Mgq�t�j2��Nu��2�^���pHz����3���%P7UXFo[�`�"Y����--�0`���՘�(��a��C���`���f�̍Ɯ`����9�ڛ/�c5����1�bD�(�vٱB�,ϕu>u>
�@./6���Gi5�tD&N\�����ػ6��0�4�k2���(�F�{�뢧#�TC,������o��L�x-�l�������Ƹ#���~~"�<�A��)��g�;a�[���3p7}#]�nמJ�{x�/���T�Q�9�V�?��D�O��짱")�+��d7��Y��w�_ɏy��8_�L$Ե���0�{Lڊa��]��0�l�ow���O�4�Me����}�ȷ����s[쵺����NY:���i�Z���ݒ��{Y�����2-��ύ�9m9�/7� �/{g<,�@������s�پ%�XJ)8|3U	�r�i��g%��3s��	�D}���%TTZ�*%�e�v�Sy�r1��Iأ�g"ԇb�UK�:d�[�^���i��bجu
.���Dq��zQ�3QA�O���/�#�JO[����[r�$��r���Z�v�S���$哞9�t5�v�.[���m@�;E0C�e��c]:�/��+�w��=z��O���a���Zf�>�+����RF�A6z��=�%O���a%��7���ޚ�r��Gk��)?Z��@�Y������U��^��bߔ�y����z�����_.()�+`�rė� +�*�80ac��_�.�}ji������q�u!�4r��rT���'j9�眳+2Y�w����Qj"�攧�:�FR���8r�ݧ	��F����{�봷89eA��N\p����j�q��"觏r��A#�	�ٻ}1�>Ί�*�@�É(�[�ݖU���G�L4i��h�����F�FN:�E
"7m���>ll���a*�Λ�6�G
~ʍE��ߩ-�������&� �Z��Vxv�i���t����@�+f k/��w�C�(�R:(p��Ξc�H��E
����r/-��'��J���8q�h޹Gx� ���:E:��8˜�+�V>�Z�p�ڭw��	�c�����]w���s���."�M��u�43��3�1��O\�5L���گ�v	(��g�U=���u�q�<g�uƹ��=3�G,�3���1��
��|��a�FDQ��A�#\�y��j)^kRK�������ugw��?�h ��H�jK,�n9[r�W�qd��¼{��#�hbr{�Ţ�׸�0�1%יE���~Tk�#z:}(�;Ǟ�"�:K�ڙ���W�����2E�6�-��B�gK�zj�%rZ�����E�rb��3�)yl$��K��11E�?�*��!7���'xϳ&�E��!��9f���Y�����g�̷��m�w����碡oß�p55O�_��d�ʄU�YWLv�5����=��PN)�j/Y�������Ω�f�8��Qv x�d��n`vKm}����A`P�y��O�[P��Wv��)�<��fa��۞�+�S�i<���W-9Z��H���4X��!D�{�����k��|���4"�>�]�w�5�c�UY+��(踞4 ��,����m{��_�����4�u�(�ȱ�c D%>)�M���(�$��q���4�Խ�����&��u�%NY2���k���W�ܒ׶�|��S*��BC%wp�8���EԨ��8�YofGEӧ7b8l=2*��AVvN�fX�q�k%N��7byİf�ݨ9=^��G��潿�	��Z=G@v��5��њ��_(�ަKn����j~G��\�&������q3�\e-�;���R�l���;E�7z�l��{�3T���Lu���B�h���'��XO��;1o=@]^��@�|�xP�9̻?��2 --�7�F=\d<�4�W��<��dܻ��j²��`�M�ޔ3�m*V����-�f|��6��&���M�񣞑�7�n+z��T�.	`�}9(�Z�a~H�x�8N"}�:zX��S���_ȼ<	��y|K�c�h�iV퓖p�>a� R�T3P\�_ly�>���mX&�f��� �;�%ح�Gm��f^w_�++��=s�QL�6Kz|7��YA{��*�I�=ʼ�=�����Sy~����aZٷ�4�9p�<-��8���BG�:2�.i������U/��~�!W��D�u�ot�ur�B�'bM�#\����PB:�P�jQb�Y�6��υ��U�;s5�c��1�nf�k�kܙZ��7�Y�@����!R�{�i�%�5��"��ߪv�>[¡]�vNr��ŵIw-�¹Q�œ`km@@�%n29�L�|�w2":����\��͎��gn�Z�R(�o�
v���[6:2����R��8l�����Ku8���Ь��<,�S��X��8%�O��;�9w-���:e\İgg��{�|}'D�I��&�͌9.X �q��M�6�wid�C��֯��v~"5������?*̲VXI=N�m˗�M�
�N�U�t'^p�`��p����nX�.-t��z�2�h���/:�|�c�i�coe����K��5�q*�Ʊ������	��Yb���M/�������wt��y��Zʵ�F�b�C�EF4�'^�t9�>-��N5{yK'�f�m��a�n��lZݡ�,<���H+�s�N��{N���&�����U���fxv�����din�\�=�mf�Nj��h.��==�KU�R��l?�����-69���d<��.�YU.��WvT�t��ɞ|`�������~�*q�o�i�5�>h�h}b��[�[M�xe:�l��[mk�b�������)>��g�׊�o�`J� 1���a���D'օS�-"{�m��V=��T�0�I�sz�����W'�K��(��랛��@1>�GP���f��|N�vQ�c���U���&j�|� [V����ƺ�*5��`3��ö�V�KsdC���hˢ�!�r�З��~�f��/�iﻋ�BҾ�ڽ��PGqL�RS����M�D�,�R���M�5l����JQ�i��:����m��f�������1��K0�׸�vH�j�I�����Q.�z�?����x���֋�0s�Ym����}��0C�ĉk�J������>�k8�mg��-���uq&7��8��j�4�liaw�P��y�#�|��>T��t�)�:=��6���kNtlo!���{���ܴ(�Cj�t^��x��	�	p��!F����fVe�4�ժ�i�{;Vj�^�#����;��)�S��|�F��t���q�~~,����7���8=���m�+GO
�|J<�����f���$d2��64b�H*��,�d,��{n�{/��f~��#+GoK�)1��j1�^O�@��v��RC�Q�3��x���b��`��������k�H"�ۺ���3�ڜP|������LĿ����l,Q>����(�qi�dHʤ�H�`*I`��@<j�D�w���ܩ��۶���K�|X����s����u{�*ֱ�2k�+L��u�),�3�F�U�fFW��pU{c��XbxsB��T5˼i����,��:�u���|Ǚ�#nWS��I�:�x�b�i��U��Qc �㐪pǞ9ȡȑm<�Ũ��lKM��lu�f�VT�5qq��Mt6rGE��R���L�>t;m��lVj����F����J�]��j}�*�aK�qi��q�^[f,Κ��eu�ŉ�-}Y���ߤΊ�j8/�����g�h���+z��&������7='�	|�Cj�F0��d�ΚV��j�O�<������91�^c�T1�,�v�f\]�B�r�s[zr�\k/?{!��E����gluQk "�;�|�6�@�д��XY"��4Y�̀��N�V�݉]hV�������ŊL�ewDt~�_Fq��h��k�>�є(��sz���z��Q�d�o�C� x�4���r�0��4�F���'65�l���awK] ՝3iA�˚�)�g�
�%��s�$a8�|S�h~y����d{B�Rg��v��g-v����W�eT�.)d xϩdx֨��L�`(����q����á�9�����U/��5N���S�T���
��k�dA���1a��`�ZD�;�ޯ�2Ǳ���n�����(H|.�d{;�l��8�w�8�0ʃ4\�_9��M�M�b6&k�(͎��J8�C�=�Fa����'���9y�cl�RE��`�_���Ш.���Y�M������'�Y����SӁ��cQ�cqW��K$����p����)Q����J�.�:���Zh[�N����ܜ�.���@��4����N�˽{!Ё�W�X�jJO����s~5�^ֶ¿�u$�L�����6�Cz7F��n
��Χ'Z�s�T`6Hq�x��C.>ۗm>�wZ�ˠV�9�';{�u��~?���,����i8}D�;n�]�
kܿ��jj�_�GKߋ�^��K~q|�<m_R��~����v�]�a՘!�q�-��n�}�i3�,^��[�AT�[t�֌��󶋛P%g3��5�	PV�nn��
�yG)�\��6���'�.�m�#0~Q��[��͆Y���:��>'���|̶5�	�>���}t1�(��~G.�o�I�ë�F<�t�:�O7���y�\H} i�:��=B���O�T�q�����ѱ�"�7��^�(r�s�q�ZDz��h<��h��2�Q���=ǟ��X�	�]SmK/��/<�r����o
�6�&����L�C�A��;�}��p�.��f��;3�p�=/1�>9��b���0j�P��h[�C4��N��s���Wq�kq��b
�t8�mV��`��`	��)��k�vaL��Q��n� ��"6v�lu�A�C lgV��UKi��j�r��5>ak��O��֫�%wlL��i}���^����G�M��	�ˮ�[3:�R��T5v�~��/�bL�`*�i��|gײO�o�(���i9}-dU?�_ Y�.�jS�ۘe{�\A�=s^�XOR[�v�����W1_v]��6s�9'F�(<7.�w�2�˼�1��%�H^â�5����E \�W����������w����D:�-}�f��n%�(Z��>F�����aU��j�/s=�����n��y�Hy��Hai���~`|���~��Xf��j���gU�Zɽ�y���T��L1�����Lxy�5g������e�0-S�d!z[%�vj*�d���L�ˬ�k�KL���e΂�;��gF0B��qS�S�6<�u��픮UI�TFNW�D*O�N:�2}�!���)��}����Ù1�w���i��tyrv���.Ȫf19��9
]V�A8��ʦ����C��S\�c˖+̺���$__����S+�l+qV��mV07�4�3QMؔ��JiJl�VP�{Ս"qT;���x�ٸ�g%R�p"�/!�/�v�������NT\m/r�#��"u��ȥ�}�t�Q���B�κ�]� ;c�~sP@�B��&�߂mH4f'XW��S.���'���Z+
��b+-�c��yk�W\*/&^4Rz��R�u0-z����fd���?A���Vń�w�y2�~g��w2��'i����R���Ÿ����ˌ0?v
�6�C8{j`U���ߠ���Md�̩Rq�O|�5�w���M렰��l&&�=׃��Y�9m^R��Ugv����6J}]��|��o|�WU��xR��OS�x/�>���M�D��[6�]Ӎ�}ŵ��%A�ΆH��Lq���`Wن��PC�eph����aO'�I�~l*f	�;�Z1��e�F�����2/v�y�d
�#@���=Y��<��*�r{'��k��ȴ�Æ�qV>d3�=��^n�=�1͈��>h.����f�����'ˊ�>���n�;<?f�j*$t��Z#jC�-s������z��ʄS�Ŗt�:Q���r�����o���7*�*G�=�σ�����Qȃ�Rio@�??��.9�C�*�̓N,:x[>|P�]�ۥ���e`$ q FD���߅z~�+6u=+��e�88#��l��/>"5�y�|���pu���]��'L�OZƄT�[�kk��%_��C����@�5$s�&N0~y������5<C�R�p�5Y��7���衎�y��&<�oV��9���H-�|�~4꾶��~�э���?d�eZ�u�@sZ�k��ъ��.��F��p37��I��J�!�%%ؖfQ�& X��"7]�r19
�O8�=�����0��`PI�wa�ұ�n����#�3��/�\�R��G.:�_L���v���ლ�-�C��f@\��[&B5e3�y�gG�I%�-�%�'�p��9I8:��8��4��.V�h�D31,�s4�+��㬫��������9uN�'6v6'j�nحQ>4S��t{׶�����F۶�QL�~/f�j(��@^���[���V}'	�8]�/:N���e_s�p+(�X�;�2�Y+�79�J��O3e�׷��q�"�i��q�駕�f��Ї�q���uub��%�l�i��l�qt*k� �� �Z-+:�O�nE1'�0�%ʹ-����So�4i��ϳ:�:Ej��q���ۚ3�m�H]�9�J���9W&�]�d���7�8���"�	r�v�����h����k��Vb[w���5Nʋ>*G�W���bݓP���<4�_\���U�9���V����M�נ����7HQlo�o^��S/s����a,Ѵl�d���]ZX�!4r�d��̫�3hՋ7�K;rZ��2V�9]#H��s�]��Y�/u�h�Ƃ�}�뽂�����I=wq]\W����n��j�,�=�"o7c�&Z�c/J�]4we�yHs���;H��ܣ��9�٪Ib�Fǰ-�=:� ^p�V��%�.W�(8[�ЧW6���mӬrڶ%��۝a�z��l���g���;��i�
Gm��FMT$��8�4�
%+ⲥ��ܘ9d",T�Ќ&M����\n��T�$�&��\��ʋ��sc՝r㬐�|���H�1�T�3�u�1��]Gn-�����`Ɏ��a�H�i����쨪j�,(��T�0��3P����n��SB*�H��r8E\���ٺ���{4����^�x�6�T޷�V>��G���c�+P�(��r:PqXR��s)���!ԩ���$	C�����]Gw�G�B�5Ϙ������.�!BrK�C,���������5�UҦ��v���n���xi��tJ���P�nt:᧯`��U���*E�}��Q}r_c��jj��era^]����Hs�+,�f�v�����^��������탰�V������Y��;h��)ܝM�˘o'i{ҵv^�Jdѻ�KP��S�Jɹ;�Q۠�p-��Y������M.�w^4�g�\�u��Oɔ�Ф�Gc�F��_D+uf����6��t�6�ń�y'S���+�݆s�:�al^�')�N]-ZP�[5L>�]���"���˜�䙝�/�Q�H�7��)�ï�����!�C�4@D�bm��������p�֒!��ncOOߏ�������������_�߾���R"����×�=mu��5��EF��ӠnZ��ӟ�O��������������~��"�X��b�������3�i�5AS���n�~mƬF��u\�\ئ��墔��F-]�j�:��V�tT�
������Z�'[IO*t���91�Ӷ�k� �5N�TCOQ��MSՋ�j�(�"���(���u�K�I�{����RĵTsj+l�m�X޷��Ju���Z!�-b������ъ��vĔU��\i�#���)�(���&�y�*����ӽF����)���QQMMMCm���&8Ƙ"��i""��F�Q�/{{Ƌׯ��kgz���ջ4"4fL%����Q�Ӽ0Y�O�]oY���c�X�3�:d������G�2���^���t�,˦?�8����l���s�z��ג��D��lM��cXW@����n�wz��&��9��4Ϟ��S��2��b�B��逡��9eCm�\�<�d��w�q�\��(�.1�JׂhSu;S�H�N���oU��i`؟i��m[��Ax�u�Y'+b��7��I)�6��I5���<����8��f��R3����k�H��)��f��M>�.��R{�(-����j���{yml�>;O��@���c�s���T2�#��N4���h���e�3�h�%�,�dj�P�6WT�K�в��2�/m�s�������B?>�Q|�Zg�wK���+fui�ݦ�!i�?,�ܣ8!���Iƥ�Nؖـ}1.�Q�������1����Rv�9��S��SD�e����f�
�<.��ke�)L�x����@��.d(ւ�������/���)�����o51Ԅ�ҟi�GT�l���Q�����Q�����b,廐%����8G@ư�Ꟑ�Jjf༰k�f�r���x��fҽ�����n�R,�j�A+��׸3�v��+�8c�����sL'}�3��8s�mZ���+���rl���Kb�	�Y���:�%x�׋�^�t�z��� �;&��&V;j#���tb���o0t��]�b �!�Eׄ#=��S��r�kKa��B��-����4 Ʊ8_v�J�WP�+�b�$#{�Q���kH��8�S�����Pf�� �	���=H�M�m����m����+� _@-�g��?07o�m����q�a�-��+�[�j��=_����z��K~ ���z�a8�j5l|Zj������m7_
��J�j�,��z=�S�w���nׇ1�t43��F}h��z�ۧ����RuѷӃ5]<����\&R�J�R�v�[J}�i	�Ѡ1z�����*��[d}�T[������ϨB�'��2mO�e��0 e�:<�Zn�M��+.��/��3 +_����ח���._��js���1�(�T̟8�C�f�B�iA���_ܡ�)�qyp�/&�p���3����>;t�;AjK΀���(d�u��I� *|R;R<�n�0�9H���e������-��SO��F�Tk�:dhd�ӆj�2y���S�^��̆�ݿY/i�OyՎQ�\���l"~��;,M���3ZX�s�vǞ�ك��gi���awJV}��L����m�v-��Tg�74�.�j���.
�y��֛�@�̼q�Õϖ�"+�q��>:��{ ������9�l�l*$�;��xxU��;/z_*�@ ���C(����Mo]����t��'(xc_�Qp?r�1|�/	��Y5�;���{w{�f�X�+�Ct�:�I��_'�,x�p��<�fK���hL��uo"LF���eCoQ�~�Q���+ޓ+������/%����4>@	���L>zh(���}�������].DRu�=��Dﻶ�qc61=������\����{NŬ��P���,-��>a��I�f7��唁<ޑ����{s�P�r�md#4:݋�b�Hބr3��.}��ȃ�P�@/}�����0��;�d��Z�c��c�ŕ��U��$4���uP�?:c�ɖ�-�����:���}PG�<�D~XO����|���՛ �{qj���1�i��W��♠TZ�T�z|^���=�"T�q,�o����@�5�j���!���OX��iE�wnhJ(0�j��ѭP���#r��?xO��ުw�����v�^T#/*��ƹc���؋@��n<�t�7&!�����T*�^���5��P[5�i4��Ry��W�^��ι]��C�*j-*ր�p*y���NAoGE�����4���>8��!��hW�.χW�V��n��%��n�23���CI��*�����+Y�j��K#��6ZP�:ƛ��t�����N.���	c��|��0W���琦�VԆ��t2R�ʹ�P�{Ս ����"9�}!�5nYó���n2M�1�BOtX!�D��xgh[P���S�aS�汳�66^e&��3�oZo,^F�L>�{c$�-"����i?��,��m��3�7bv�(�9�J�y����uh�R��QZm�lP�S�ZS�l;M[�O,KgK�U�vAa���&�D`�ƌ�KM
нs��f]	�}S�Q.}��o��B�ْ�Kb��=�s��	4% �2��[�X�K�d�\� �B�����H����i;�6+����(VtT'b��+t�����F��y�P���lڛܝ��h�h�ңG��Q�ym�:�3'})��n=�وYcY�q�a�r08�Nv��\AE;Vt�Xc����}��jDם�t�h���Eݙ�1b��5���\��ʍ�̉��[���� M�C�.� ����/�,�3��o��v�^I�kL�3o��E[֮-����Ao
�86߽�o;θ��㞣?,�M�<F�X&<���[�:!�����a+�\�L7��?��R�9�B�] ΐ+S���*G�h���D_�ܾ��Vm
II}����SF��
�a�m����a���'q�PВ�4�XJ�fv�oV� ����b�G0k�I+�1{��vt�7����½7�^I�4G2yRy�<����5���2f�<j�ׂ'���8�G�� k>��YW�N�G�_$!>�~b��R6y�F6���J���5x���/;��u�������ޒg�2]pߋ�+���D>=�͇2}�n]������bBSi�Q�������2��v0zuy���L�+�3?O>1ǟ�w��Qљ�L��z���Ot�&��M$m�1m�����\�U����מ����S
������y������9�U���}���]w/w�˃����9�_���>�[�S�=�
�P�/ތ�a��v�0�sRӜA�Ò۳�����$l��t�$�,Y�5h+*��x��T1NC�O\
C�<N�"_��(�!ա{{�3�dkoTQ�,(���&E�)>��"�(�5M�-�CU�d?�!�������h�X�a�c
ѡy�AG�;N���j6Kf�"�o,���U���gT����j��+�YT�p��^��x3�L!��Z5�;-o`=l0�ħEk�rN�H��o}C� s�w{2[��m������װԉ��߷�q�]ՕwY�dkVxM�w���3ۀ��������u�S� ����w0Ή����Y}�i�B�se�ŵ4����Q�����P�S�vc˴���@��N���ޑ��$�����z9OYS�F�>�����[� ~r�����u}Ԏr���R��ɭ�u���B��w�2��{s3�s�]��0���ŬaY2�=��l/��%�xq|�b���ʮ:I�Ul2ǌQ .��n,h�%��u�<y��Ô9�H�����#��&_��V悮�r֜�O裱��Z��*�����\p�i�zV3G�uF��[�ѬE��w�xe���������44�:��@��^�8ºE���D��~/P��a� v�{÷Pf*���46���
�H��F'���}���ރ2�/ݦF�Ի�t��3l
�+�S�,�g,�]��H�{]�E�5�� ��
T��ќ�2Xk�,5;;�hP63��kMw�Sn�`�w��O�� ��������Y�g�V>���#<���eBF�b�����g�mzZ-�R���q}c���h�T����̴$[�ץ�b�Z&B�o�)�-�IU�I��T=��^�Ji�,.��|�3n�}�S�G��i�����[*�Us(:�W�FZ���R74���S��b����ӡ�.��֫�Z�ci�p�H�bå9㛼�0��!:r~�'�'KՏ{����&�J�ޭ�--�xn�Rb�sC{쟱!��YWgKW�L�M͖�b�#ř���⼠�$k����½R �}�3������XB^���1L(�1�ݰ�)z�{R�lR�u�Sa��VC�;ن< =���d1��l�N�6����UЋ�Ɂӽ���k���0��,�)EYjS*�ri��y��i�?8m�Fb�=,2̈́�g:fˍnl�l�
�%>�[�-�7w&z*F�c\�%%W-=��1���-@p#OK�Ժe�H!�Y���Ry���z��Ȯ�����z�a�0:�.Q�]T�Q�^�}:�Pa��t�,7᭥Aֲ�;�����z�m6�Tͦ)��s
Ԧ)��*Km�T[�B�!G44�Es����<&�7P;����w�����cHSf�/)��8<mW02��\�8�>�G/"�L�d��^����N���]q��#�LDsu�݊dM��<妻 �-��K]%
��ޑ��c�����S�����p��!�z p�ǳň�5�`�p�S�ΏKbJZ�s�Zq^�����j��;wVD��j�[������A�j��z��1�^��G����w����!D�텤��\�gkQ|���ڣ���,�,��Up̥����\�&}ǔdZ��ܓ-�¯�gcԏ���Y9k}�,�sZ�a�]���텍�yj�q�w���V��0�W�9��*[2���y���>-�Yy2a�zm>4鉑q�.��n^��e����y�o7���:�n��HnWl�L�>=I�dD7`��^CGS_z��Dg�_�V~���/��!4�Bӓ�[4��k��v�}��C.��>�c�\;,����Ч���֗�$����}GZ�$�MҮt9ظ��j��<�����%�X��ڿ�:/�{�o���g��+��,oK�:Q��\��v^�����ʪ�d@�(s�nN�%�ږ��c��Hn����j�U=�f�6�g��|�=^ Q�����/��W�+US
�"SM��+(U�\���cj�O��m]P�b̏B<L*��(Ѥ�����������*Y?N̨�˗���U���5��I{^�=�̹z���͕��b��F�L����ґ�	�b�	'Y�[X�NL˭h�Z,�AjQaV`RnU6���/��"���7B1��UǇ<���#9س�1Xn]� �4�b��:aET!�m�s�v�E��gE��-ŨDx��@~�T.k�ޮ�ܹ���>�`�X�ƅ[	�ٝ��E�.(S���Ugp�O�l&R��wûH��ܦ`=���[&��S�Ξ5n��|�e\��|=?�V,���K�:�GF�[d=��P^c�s�����V�]վ��T�
�@�SSЎ�y ��泟hn��s��/;����͸-��V�{;�鏫l��u9U�<�of}��Fȭ^g�^m�.����b��*tzY�Q�xm�9ƹ�B�=�_�"�Y��7u�i�2d�8~�y��6�!�+<B�GǮ�C��KH��e��F�Hص��_����(s�z��ч��dG(�	[�AM���x�����$e��6��syViI����n��k[	�ϩW��tΙ��Dx�p���
~>yP���&қ�|/��/sqP��3�� �1�ޞ�3�?Q���[��_��ꅮ9��)���.gI|]=|"��A��,8ws����A�M��>J�����`��'���'�m�]w��9w��r4d�3rm�� F)MR�I��f�5����v��a-��%��ǎ+�F����蝳��F	�[J2��~P���ݻ>��������j�w3T�>I��;�89�Lo���F�h�G�;�@�j?,�N�bj6�4��P��TS�;���M���������V�a2�@a���)lÆ�ON�	�,j�_|`������g;|�q[���c�����hYz_�J��c}U�����nւ|��'�������?�U`�뇖Yx��u��e��GFP:y��SWH��N��VO�m=�L��*V�NE E7X��KVgV�=���M�C��ǘ�K��մ_��=N�� �oxte��u�PB�3�ރ��!ԞQܝ��ny\�QN\pa�0;���{��Ys��4��ap��融�ڐ01��vA�蕏�閹�)��h���F���,Np��R}P沁���Gh0yy�:%�: �nCE(��g��<)��ڔ�]�l����c��3���1L���:��R��z��3x����m|K�?��3~�q�D�����<+^ڌ���]�l�����}�C�\dw![żB??�P���xd���i��Q3Ɇ����9e�aL�]f��ݸ�ϯ�%.�i0���k'�c��ܨE��P�''��[n%�'�% k�B��*�{ʂɨ�̐����\9�G�L��_�ιV������'i]ҚJKa�sT�l���Q����|�;�nhF�p��#(e9���[�kd�_�����^*m�6��e����k�>T��z���~0�p�83��zW�>5h`͡;|H����Ǩ���tZ��3�}"��2���ayႉ�]L�7E���wgTJ>ޡn5�Z��3��L=�V��t3kOmDTa����B�H���o�t� Jlm���ҷE�&�ڲ�ͧG�}BQE�Սam��#�;�e٬Ӣ����-�0N`/�n$���r�^���`�!��`ːf�8�|lTْ��D��-���5lʶ`�W#`�=�Ռ\��X�V�^>�Beب�bҏU�����^ݟc�*��b��ѷ]�������
��\�6��{�\���9�'���ko�R�/�M��]
���E�;�������]M:{i�i;��|@c����8�+-��z1N����K�D81��ܮT��݋Ŵ�vo,�b�W&5��wg���f��7U�@Ԓ�66�h�h�X��W�TB��v곇Xu��EMn�B�w:���;tv���T�rI��7�a�;Z���֑\]��Ŗz�t#*h��6-
���Mj�ufI�+^p�#A1H��S2Z�����b�tZ,H��vk��j�%��M���݂���ή�D�M�g/wL����;��ջ�oD֫6^�k橣$ ���#Tw*���'t�\��� S9���y��]�jn�m�m�RgGz���^}cB�c]�ձcYk�P���E���X����-�L������rf��W%H�Y���gY���I������R�8�7���`�{�jI,�ϛ��ͼ9;f<m��y��oP�(�(㒜��z�`A�״���b�R��#֋4�ur�,����R�&D.���/?ld�Y��n�S-٫d�<gf��y�3wX��o$����	�9��kX�=q�-�	���f���W�N�!�kBƉ�3P�Y�8H^�N~=Iq	����x�s�`�����KN����$�j���{�#~�v7*��"��ݝ�\�gtS"P�{��5��\4.egt���M�v�h�D��������ݤ��]��S)��-8�x7�\b�"�"�d2�U����zz�V���o���>����ud*���������%��»;��4�-戏#��ے�K�''#��*�;$u�Բ�e��
R��f�{;�g�S5:��)�7�6�f�,�r��|r���bYT�Cc�v���d��ۆ��U���7�
xj�ܓ�q�3u������v��\Ջ&j7b������-����%ɥƯ��9��`�yiq��%l���wU�fm{��(4��2R�6��[cV,��]����3EK�]�Vs��R��v)�`	�'bغ��N����}���s9��§-|�U:�*i�s+
�M�F�^�U�A��;@�b^�*�r�z+SV��!�9���X���,&kEҗ:<���eQ���r-�u ��5�L�unWNͧ�:G�tǛq	Sn@�K�7��5�ǋ�Յwc#����/���)�0�-K�o���iį%�yW�,��1��6�jPf���CD�lTB�4�&((�)�z��)��SES���#���|�PD�3IQ$TD}>ޞ�oǷ������{{{~�_�DMPULT}�{b*��N9;�1��-QUD�MQss����}�>=�����ooo��y�1ƪ&m��������E�]ڽZ("�rT�U5Ds*��)�[>�f�bfgF���ՠ�=lU��LII]^�a��*	��b�h�("��*������1������QAE�x�R{�Hŵ��$�%:5��ۛPm�=�X�E�\9T�LLE�n����Sͪ"���Qb���PPRD�CT�b"b���-UURQ��oe���m������Z4󘪈=�^��<4i*"�J�7��
��`�l4�QutG*9Y�]E�shѢj"J(�(���*�*��)�"���;Zj�X � ��*J&���IELAM�U4Ss�������D�8��c��krwo��=ǈ��gC-�EЊؚ�:�qFX���-],�Vn�N���+��"k��w���\nu�U�Û+t�I�ԇ^����{��7�Y$�B5{�C��Џ�D����av)؃f�ך���
�|����P��L�լ����6J͆L#:��7E��r�o�&4�������V9a�>�z����P�fIټl��5W�*O�K6k�{��/�T��Q.T���'�1�t43��5�[
D��=���1�!�n	S���3��y�.vp}g˪�z"��q>��5�MX�>�ޏay�%�F9��ˍ�����;(ֆF�UM��P��e/^���aT��}N+[X�S��
簗McZs�w��{iՌ@��`Y�O����xF��4�(oBd����mnPк��ؖ�����c:�߅���Gt�=9|���
s��G��QcF\F�K{_��,yTvTT�-sX,Z�զަ�2ͷW@��\Y���Ȃ����L�~��<=�Ll�p��'5�K�Y%�<~������ưbl���.댲O#��(�z��K�����w�<&H#��4���ˋ�eKUM	����m��:��e��0���=�cLsm ��
eKËר{���|u�����J;~K��&S��LFZi,w��ĝ��ЭDS�WY6c�gcyV̩��!ܰ��}��D��tǢ�9�Z3�5�nu���Λ3��|�6	�^*aVЛ��nlbj,�BS4�$�


Õ^0uޢ~W��6	&��<Hu�*0/{f�^�o����&p��,�o����ǞyT��2a�6��X(�dd��	�G �!��{]<��LI�M�&�-)w2�0DG'7�tz���]��Q�,�y�թG�Ӻd��;!�����}��W*=���`���0x0{�,�Sȗ�S�������`�犒�2{�_�;V�U����S^��3���y{�&4�ށ@u�BM�\���_'&0s^��7X/��׼6��R���K�Nw����?	��E����ʿC�<�2'C�q	���f�ֲ�ݽ�n���X��=?.b�P:�qT�L5E��K>�Ϗ�"=��Ȋ/'u�FX��u��;>�gH0���|��*� ��Ff��%��^��ތPϾ�E�T9MFܝ���Hcy�r��!�m+�e���^��71���T���6z)A���!tհ�ۊމ�su�a=Ɲ��C.�"���Y�(O��x��156R���D�(d2��e��6�n����_q^���4��1�)Y���0.�f�B��c�-��~���3ĪxqV{󻴯}����p���[�(gV�]��ɗ���bʪ�;�0�>�1C�5o��[�Uc�h��K:��3�gטu�zb�>�톨��+~��i%�q��T��%U�g�<���4��vn�4���j��7(v�W·j��j���s���o7�xӻ�R1����7?�-�n��Z���K7f�9�;2.¨�2(���d/ѳO]�=z���j��ܩLN�D�W��G#L��\�+�;��^5 �儆��9��-�U�};vq�1���ץ֔��v�-:LL� 6j�J��gN7Q�n���uȣˍGK�"�1��2�]��#���k@���9J.+�eT��I�(���R���o#`&�-���N¥�Ę��x�wÂc�a4\*�=���Ϸ��4��3ZM�����rO���N��S��=Ƈ#ȿ�X�W�P>"6�;�*C�������9��I���<rok"s�^1�;(OAd�8Ս2��͛#���~_zw�B|�ʄSˍE�WM:���zؗS5�-q��m�����T����Qȃ�`lo�Es��L-�_7]�Z�iTn���s�Рe�Q7�֍۾�cT��F5��y��b��.ā{EJ|r�Ff�۲0&�����
���|c�ǹ�E��:t��="�3E�����n��*�q�&IrX�a� S����fwglӮ�:��Cv�PZ�)�R-U���9���޳�r�F�*eg'�*� "�X���;&�+��U	���P�q[��lˮ���4�I��ݟ˦d[����<�P�QS�6̍�F�q~@7�x�u�f�3L]�~���7<���T;a�����6͸�o�}caXy�I�_h{ӽ\�߾u�--8L�*�3'�������e��[ވ�����jGW�f���Ƈ$�^�g��6��2���AV�ѥ�ӵ	.zQ隊a��E��e^������L|W8�s���0�$�)lÆ���I_�����N��Fױ�ߖ�ƣ���F�Sk4��#5�P#;{!)�!tڮde%r�-x� ��akQ�|h�cI�/C��Oq��7C��9�׻!P��X��&\��I��
�j�L߹E���݅[�YT��;�Qs��?�'�pfAf�u�����8��*���7�+5��e��qV�a�5wzB�R��W}������ڀ>���������?��)Ѥ�$�x����	1ݝ�+3'�k�.45����p3����R�1����-3�EP�!�呓G�VV0��S%s�["��^}|�\�w�`i%�?�n�6��^c惮**�����k����O_s�*D��PWSK4_Zs`�ܘ^"��f�WDl����w�W;׷��ZJ�	���[@���)�̀��<0��l|���Nx@o�5�}_%���o_#[r{&^�����B���v+���/cg�j���=�ϛ����\9�������2��:�_djegΆ3y�}^"��ZEY�s5�!\�;Jn>T
�(�0�h���.fkU��h�ډ*Q�4�u�L	�RXa��<Ξ�q8���m �=��"�M%�����|֟.����.'�u��5��@��9aW���{��C8-�����O�UI�eß��T*���Y��ܨ3";���PKq�#�1k}R$@~����3�T5���ر�6��v�7#\?'�OV���!�3�M����ta��v!�޴�����������I����99�{��A�1;�)ja	Lp�w��ϴ�9��
c}�
,1sCQ{��N�\�қw$��<t@^���G�(@#M�x=تXF��*}���Cμ���vʴ���XW��/��v���1t%踶��S���#p���m��k��.�\���B��~h����y��_'f7��Uy9u�Ģy��4W�c�a�W��gt�e��a�jY�l�G�UG�R��WI[WVl*��R8�#��4�}��wfԻ	����%j�~{�]�Ć���rF��RV%�c5�����f�նˮ��V0�''[��
��UK�|�6�����k�	��-�ӹy�)	��'ܶ�0�v�ĻKȗ��Յ�DVxNMW2�0nw{|�aC&C����oy��.�Lhj�A���;x���p6��k�C�W�����z}?gȹ6E�Ӻ>�2w>��F�[Y!]\��\O��к�rl�Khz�|�.W�{1RGo4ni�2��[����y�V�#{B�H��ܖ�"�87U��<�sSw\�\܊��q��֜�q������'܍������I�kk�<��O��y{���z<w �#Ǟ|7�j�Q(َ�k_M�;iHV��Qzfs1e�f��}�r���=h̍�E�)h�j��e�m�*�&!�"��-Lg�t>��޿Dj�����QXj	]tsAcO����\�7sY�`�͜�T�F�1�`�XbN2��)1��+{fe�k_��3�V��A�Te�<�"�����xm��'j������L��\M�8i�o�n���/�n��"������ĵm�����2Aܲ����z�ޒh���������,�?���s��s�C����ҙ]��-�����q]��D̾M
�򫺞�ӝ�F��x�I�7y&5�ej̥��Y�.������V�[��"�76�q��ޡ��S	��-���x�-���
n��8��,��^Ɓ{��[��W���3�0��ԕ��&�e+��d�V�捝�3���^��^,��]�=�'�!��Z�c�T]ΐ�a����k� 3i��S���"�¹_�Ou���9S e��3F�i��=�;���W7���h?���q=^5M�%�D�\i���p����w:뛻2o�c�y�^��t㯍��U�b�|,�E=���N2�����n��2�o�-V7��H�[K&��,*�'׌�k�?��ۛ�he���6u�W�?w�R�C��DP��{y�W�Y�+i��8%<�?<�74y�#(��^��:\m�N���4w$hs�4^M�	t�fn�lh���slW\�c7����y?��rl��5+z=w��9����k��t=c�،Ή��]��9�<�h�g�nG��>���	�oR�FC�F�	Q1B�闁1y�FOM���p!0׭p�fSY]��͚U��Ӌ�߂��>z m�e�:Y�����*onI��	�S�w;#�Oz�C�+�ycG���z�S��� ���97!�
�v��;2�2��&���U�b�a^�-Fd��c�~���߇�w��Kc���^6����J��[����쾇;��}Jt�[�\1�71�/uG]�6��j��z뱌�/�����^������ٷ�F�������� �C�$	���z\�,�t��=s�:�"��P~�w����8�`Z���#s�>��z��]�F`v��<1�[������LN�g��Ľ���Ŷ��i�}���gK�	����Ȭfn�Eh��5G4ƫ/��""�H����<���b�0_F{*T<_*��v2Km1��j�=^���&��er�h�Ԏ�<d�S _)7B��b���uu6�r�KQ��[�%��QS�T6�f'\WW���"�8�<�D��,sR�QY5$��{^V(��U�P*����,�$�h�_pvO�+����4��|:��n�����r[G$�T��T?r3�̾����:���O��Gj\H�]K��K���䤅C�ٛ^/u��^ʜ��+t�Ԅ���ڝ+��'l=VyPY[k�����wz3o��]���r9�g�fX�Zֆ����!�̵,�8�_>�ve���}�=�yo^�~�u��\�?���ԯ�d˓O�B��_[C |\1��xC�u������C��+���|]<:��G�h_]�Ŵ��
��*�z�����[��n�aMr� �7��@ĵ�'.&�{+b��6F�|ؘ��j��>��*�wcm<����>C��ޑp������Tِ�MK�#�Mn/:�"�J��oѹ@����ezB��/Q-T����J�2۸Uf��"�UPm\��T�[���j֬� W��@EuD	6�n��)Ѝw'u����2٫���P��˓�$�u�E�um�F�������ݝU,�ce7mgjYc� .����\��V0}���\\�%��U�"�_��T�X_�fz��3���X�pkVj��꞉��;\77i�ۣ;�|cVP�J@/!��|`g�1�'����H�)��v2^2*���޼�_>ZT���m���f;�:ý������tВ���)�Kփt�&���(��{[��1۹��=Uc�6��N�5|;ݬe�pE��1�J�ʙ��B'����6EiF'��[ĝ6']K�s�,��s�H�U�q�V&-j��f�CyW����Enb�jS��w�]�����o >`�$
R�y��*�ȿ>jm��x��Z�!*�]O�6��D�찲	�p'-��ھ���g�Uu٘e�э�"2A�9K���n�T�m�k�l����#g��敩3r�}�x�Ė�i���qy\NV��1=�+{3�3y�U!���d�
�]�G���i=��W{7�ws���Wې�*v{��WI���mS�}U���:��r�R�f�\۞kq����fc��c��%"�l�yUt������0�Ǽ�o����н�j�����ʮ�����C��x[����V���z��zb��+P��ݷC�7�jszN��-�@E�fӊ%�f�T8�*����9!t�<��회C�74�����ڭ,��v�.ޠ2
F*����Z����H�{�q=/�����P�z���l��,�mfKxOlF�U��^E^2 �Dy���/�Q�\��_�)V��c͂��ceI0�3A�m� egP��R\U(�	<h��.��J!�Tz��]�
0���oqN���{4�mgR�\FW(���Y�@۽z�Gv��uN7�S�v+cI�K��tY3jd��$���u[�M]��9,^�J����o���D��Ջ[��1�G��1��=&t�i��Sc�7��iL������m�Y�H�ދv�tN�}��V�U̜��⊥��cc��y����zSɣ8(�p����,[;��٪+,<��)�<��L�0N�C��o+o��T�gkZ��b���"4ȡū�G+���L��c�RT�쁴�Cn�s ]Ѯ��{�74�[C>����vP �V�f�5�v�%��%�����'[r��[\WG���Y̙��xG�'��o�r�q+7��)[�
$����I���Vm�����-Ir�,�o^$��K*�]���1{p3|\Sr��|�!5_L�7�G]�L���w9�@Y��rx]X@�e.�LS
�{�-49���)Ul���o�m��R�_���]����:\Us)��>]H����,�t��x �Vx,&�2����<)M�0$Ҋ����fCsb�vݢF.�۪�j��YXf���\5s�>�0�RXg=�m�2�g#����N:�޼�f�L��^5��ri�ww�H㭻���`�,2��8U� �/�u�£CVs��7��oh1�Խut��%=�q�}���}�j��pS�e䎮��pN�Ļ�]`n��_�"U��LZZ��9��3�OK۵�&o�M��1{�o�-�geq�A6�K�5Q��IV�	�4�,���w�ܳ���z,����V�r��2v��qM��7p�v{�z�P�8r��;8Q�6�ɉE��n�\u�:>������*��R�����E�:0C �A�x��*�ǃ8�=-⮄&R�HW�5��
7��,Ӱ���Խ)�S��*�RV��u�k�p���S�w8���Q�K��	��7/�+-G�՚Y��D�Ң h���55g�@�������ΥNv�<�lfA�Ö@��\�C��k�a�SW�n�ո�e�LA�[��+�mev��X�ڷ\X��|�WTg��7�b}HP�%[|��B,i�x��W���0�y�Yg���ΏKyh[�A�}���+�ֈ��-l
�ãS�\XG���(�թ�2�ݬ�`��Գq���T`L}*���O0���6oqX��U�-B��/]��[��^u���u�T=5��®���;��VS�&v��m�^��[�Î+���t��ڙy�!ĺ�m&�GL�gU�dW��/5E#9�8{#�Qq�QIu/�2����B�\�p�KNu$��}Z�u������p���t�lkK)�R#�"O#�8���t���p3����9�Y�^��J��ݕ�{zo�7��y����(xB�DPTUU�,�QI1]�T����'�Ś���
0`����
�Ϸ����~=������������ة���rK�3U2u�EUQ�u(���TAբH�����.ppu��D]Ƣ�����}>������ߏ׷����EWݪ�)���P[r��S��IEE��ST�AU�ESUr�AUT�Z�T�EUI���&�H
�i��-z�Q��*�(�x{�xQD�P�T�j�&�$�ֳ����N"���f��ՠ�"������"�OV�jK&�V��3TT�A5E4EMW\�&
��[����5UT���q� ��"�*��U0�QEU0T�KS�AT�ERPUMEzq���"*��H��ub����њ(�b�y8�$��(�b�����"����lDA5�h�H�&H�j(���
*�"�剚���(��	�&�@"H"��R�U�K�g���d�/�-���NGu��!
r���t1��(G`Ռ�A�}B�$8���m�ۖ魒3�y��?m%���.����/��6�����i�-쩝R"=a3�b�i�Lҝ^�k;��W]T�vs\��1�9=������y� &a$L<SiY�[y���ۿ c�r�;S��Q��[�9�0}��U�����Z�M#�1ב�+R�{٭��+���h��%�<k����xCOf�c���T-m�ѩLZSb�u���q{Ÿ��#��g�M�C�鶊�ǵ(H�N�89�^�=�Qo '��<Y��.�*+4���v;��]�ӌ��a[�fxnض`h�2�/n?��;�J��؜"���^�٘��F���3z��=imyS�{�TK�F���nU!�iq�#���t���}��ӥ��9����
NG^�W�*�O�c�z ��,U�u���v�k`��bIن%�n�s�Wg[�[Б����|��s��%%�VSէ��C[��N��K����
�a3}�L�]�����3��M�����Y�o�X�uC�Y�B�lW�~7�rF�v*���L]'�^'-��6���k�2��fV�yCqc���b3eq��;���.�]��c�N��Cw���4����=>o7�����qO٭�Y�����Ժ��yPJ���9*n)���Xr+.��C����!�UL
{�'�\ⷭ��Ե��oCq���Q5~�N�����ѹ��<�&�g~�(�{?P��U��VJxG������9z ?kD��u��������粼���{���9͇u�0����<VR�z��de���u�
�]PS��
[8��/!�x�қx�L �U�� Qq�xd;��K�)�E%e_k)���n{�K>��ڟKD_��S�V��>�^��XW�V�I���-��,qou�lscz���S��yH��Clv{Han1ةCLB�vpZ����݅��z�NF�-|�wsV��dQ2��uǞC��\E��X��}\�|-g������q��C޵<Xo��ܞ�̋嚁��4KC�"�1{vaZ]��G�+T��nk�1� ���/vИ�M-q4w^��M#��.���2[�������q�L�������z���ڟ^wG��M9Ykty-�� ���O��Eԗoj�M
1M��]3_f�TS5Ñ��;�oTX�9���82s{�|0���د��Lo�Ʉ,�͒s�d�vr�C;;w����}�7��� K�֍w�oo�v�g��޻���oݝ�hu+�����+Z՗�a=&�9���i�:&�! ��F��/{Tl�l��P��QS�R�\Oc�t=c�p��ťT�������>����TLbK7(ڕ�
��)gޛg_|�x���������k��L�0Y���u�1q�핖5-�nI8��^sV��0�XQy�&n"�����͐����C��¥_K���	`/]�/��h|0dk8YJ�9��>����u��u��!G�e���ֵ��d��w���+lFD?Tl�wX�f�Y��YqآGm�|��oz������SF���N�G�l5v=�h�ӽ'��GU�nJG$�ё��9�ú},�	�8!�����(�_$H���|�Q9}����R
�&�򀱫;���٪ �[��Ux >��|H�]��qXfE�L���)�|���-+m@å�c5�%�5+x�ȾP���琚˞uekQn�敷�7�;ru�r��n ��;\�j��ݏ�/���!�\�<Qo���e\�����Y���}�*�=�e��%\���:)��Hq�Q������'c;�R��~&I��D�$���������X�_�1P�<���Wy�S�Z��� n��TZS](h���޳1�(����/Z1����ژbņm
�k�����V��ֿL���p�
ޜɮ'wn�ڲD%�>�Xd��x,+��@@J�dp�Z��3�x���m�Jq�ִQn:93�x�VCi��e�Z2YE<@�F�U��SS��x�/b�j���	#'��F��j���w�SpAU�5�y�vDM*�w�#w%�ѹ�d��qu;v�Hg�������SC}��CΗ��`)�8Pfr.r]d2U!�S�T�ͤ�t��"��O�0����cҏv�|�~'��iė�H:�؟lJ���z��q�7�����l��ݧc�%��<��Eu>�e��q�q���(��0)���yamӪ��b6|v8�)q���|)U��wQnbs|~~�'~;�n��ڀC�����
�ū�5��`���S\&� ȳeL&i �j�m�3���`�>d��S��-w�n�V/�,4v7͘U'Իfҥ����4��E��zX���R�n�-�ɫ%�d����AJf.�]sy�����������s�!	A�޿Fiw�K���0����=�W<C��m�+i�h..�E�I��ި��l��B77'�mr;�#�.(��^s���W���Yq�]K/'*۹�S���:S��#��˙�f4½�-���E#�瑽KU��y�"���CEŪ̺��B.�����7�b|ݝ"Y��ٳ�̎)<�h�*h=I�&�v�c�W{sy]%��FO~�q��Ȍ�l�'�HD?�uXf�;�i� q���Aq���T��w�\�o�$'N�
!s�w<�$E����h?n�F��j~�4�}�-�\n��s���6��on�m�"�o��7����̀om�F�h��'*�$�W��N��k�� 6k��K�\�zv}�*��0��[���桍3���k���ʺ�)�͈H�F8�`i������o0��-�������?h�+���S�@� V��*	�tT�f�c���R��������σ5G׹5�8e}��_ܘ��M�N�^�fU�-������;$å�Ԣ��Kc�y�%,Kv����Q�v�2
�5�������?_�=��g8�i*{�{�����B���v�oS�#hz�x<TK����5�&k+
��U!ުn�g�5�Z6uE\��m�N�6Z����R�4����̲�Z)�)F�t����A�7[���k�d��ӋyU�X�6�UPZ겋���gc���]���k�g=v-Ȏ::�*J� ,��ƭQW��[*�Ќ��c��s7H���,�q�e�tgx=-����rVT���ڛu�{�ouy�*�����=W.�ߗR��Ӿ��*�u��/sϖ�y�ٻ}qq�������H��Y���j8!�Ȏ�\3�{�����s	�����8����w&�ux����⳨gq��ސ#?9^�<�Z M����l\Jߪ{4�ϠZX���Ab���jl��Z��튘��vO�xN���ȕ����g��UWr���<�[j�m��;�d�=s��u[��`��]���0'	Χ�u��9j�([y�Q�ǘ�Z��ʇ�g�KB�R��ՖL��"��:�/>�[tؒ '#F`��{�ì���U6�-5}�/��lH'�}s0�^0j|�<�:`.�.���ۣ9:sX�S.�X�o*\������������@B�)�ώT���D#�_47nO��ȹY"�n�omǪ}GZ�A��j�2콚z�՗�芐�O��=��:�0�����ݦ�7Nm
~r��q�Pv��)�z��]�ۻW5��{���UV@;dO;��+�V�����.�vh)��c=��7��[����)6˭v�l^ڴ�����ta�܈P�98ۗ'�VF�y���-k��
�*#T[`'k�ZA��Ka�:q�L&�kѦj3��*�Vt��H�DaO7��B6���\H���7p�l�S0��A��tN�^(15>}��\�/m00���U�Y@��*���@{k\Ϸ<]����{�|{%+O�,�&
�e{���U��q�8bߣ�gl޽qƷ3�Cpl�p��^J	[�[{�A�i���4
��J��tR�G+*�tT�Rު��� �ޣ�s�4��������ڤ��+� +L����l�f8_e�=���e�׳�{А��0uo�����/�%��rr�]��$̍:�Dc*�|���S�@a��9@���4��򁴫���^���gu�^��	��z�j�j�u�s^U��V��,�8����a��������]�{jBt$��}�s��H��sm�NվЯG��@V5�ڙ�|���um>⑹���4
ҤoJ�ZQZ�g��-F��bca�I��Mv	�4EW>�ǩ�yE�����ԑS�t�Ҷ�����T$3SǮ��µ�X�Β!q�D#1�W��j�u�
[�-�6�Fқ��bw�F:���f�	�+��F���MgiT3��Uqe�ȸ�1���SD]7��-k荱�ߧ��0�6�Cb`���ܒ��:�O�~��c3����|?�Ȋ{X��.�=��ЃFK�~�aϛa���� ��]�W��x�E,v�c�ѽ�ͼ�����/�j�~�g:���oK=#�l5^�7w;�$"mu�y�9��A$�	P�j�OU�w��2{����M܃�Cֺ�Mu���a��&9p�)��H�z0S�Ʊ�DL����,�;1��t�zmI6�9cC]�#�tH�����?v`�>���&����Z�O�a۪�}���'۵dgN�%i�޺�'!�eǋ�H2�Zcs��n�5��e❃n�m����:3'葷��^�����]"����sn����d6t�����٧�MV�Id��
{�Y��lW5�u�>���|[�������C�������$7v��-|:�f�4Op�����#kem�M��zj�I�W��Un��0׺{�)���=��|,���/&v�5�����md�Ur9[�[�|պ~�d�����	M[�^z�Q �.���-�$�އ\�u�x+�aix��|�"W^PNd3�Р�T��Ή�!��!q��p=f�Q-#����ȴ�Kݱx�߆���˧۪|�W�~~��@2�ts�#V�� T##��{��Rճ��،LK�H��ŝy5�r*Υ���s�l�,1�}fG��m�CX:�+m���=�ח���R�S+3p��Z�c��[G�h� ��Iu&j ���K��fOs_^�J�N�+���4@��� w*sC���S�;]t�U4XCgq��ɉݝ��i���mq6z7�{|{���p�9���7f���A��,���9���~ca��l��n��k�����g*<.�q���aI��*�x����h��i!m�Z`W�$a"���8Z;��1����}�y��� �<4�e���*�e�	*E�C��>"o��j�3L��-�������f�"��|����Pɟ@�V-�M��MM�N���l]N�dU��U���pe����`�c�ð#��E�S��d���p��*}b��<�-�Ǳ�������Ug`l�˅8���m^�F�&���A^1NÃ� T��5W�����]�8�m�]	���}��un�ұ!�Ů�v΂�͐#����DC�u;?t�HC�.њ �����Ḟz��3"N8঒K�W�:Ԥ�l�=j��A�=�eKWF��`�";��1��S(w(�zCy8�{,XR��[�c�[C/u��[L���~���v�
�A0,3�kzR��Baג޸��P��j��S���������5"�Y�"�{�_����^=��.io4H�wܔbzz���3kzsv���\Ϛয?�Z���r�h D۪�S�.�bǄ?l�;�(�g;����E^#t ���h;�I����93>^l�T�]��`��q��o�7���hO�0)j��:�t}]���DTr�L����O�޶3��;o:�>�49v2^^�d/J��ZhTb�E�ݥ�� '��*ġܶ���M�-t� ��fQ�)���S�(]�w�w�f�{.Y�_Q�C=����B�}����>���⮓�k'�!wT��>�ۡd�Cۧ\״ G��]���6V���*�D� ����;	�sh���Wm>t���QB�P�<��7h9����ݑbwr*E�F��ڹ�˪������2�ˠkA�����z�)�!J��)��L}oA͹.�؁ U8ˣ8n��5��0>Z��y����ͫ{|��")IFM3�M���vE��c��#�5�k#�b�����s;E�M�7�z��RY& �#z]H3�sʼ���e>ۛw����P�|�����]q�.	s��z�� ��H:s;e:{ߴ]��x�Y����M�T$Ӻ"�֬ :M�07U�<��]r�8v��0[��r��ֹr�Xid]me��r���s-GßCs�6�AC�-����ܥ|�;�:����A�Z���8�\�.�s�!^�=�Fc��E1�Q�Qxh˵:��fFIܜz�H�Eo���N�jZ�n���|U�s0Ĭ���n`!q��R�ˏ=[J�y H̼ЁsJIdT�0[M��]�[P:S�!5J��miJ�O�"�C#��Ֆ�b�]��P	�̺�9O0�n����'8���3)��2�/��s���Z�;�-��ni��J=ݴ1>�/MEA��n�gT�@��gub�2�p�I��������\�6����S�����g��7�����_T�FCy��iҦt�#��t��9Ü[A�o5B�3N@�k.�N�Z���e�b�tV�xU������=���4�S�x� ��V����N���,ڳԵjM#(��\�J圢s��2$�`��[m�<�o��Č��p�������{z5P�R��V�m>��$�ǳ��]�c*��)�{��M�7�h�ހ�c��oE8儢Ó��4��z.mN�t�_=��l���z���t1o�]���۫WhY�˦�Q9]܊-*آ�,ؕo�G� q�e�
oОW{-j=�[֯J��]4X֘�vnT�KwS��Û͍���ljy�$a�����e̹s0T�������Oa#o���*	 ]��ʀ7[�b�Z��!�ի9�+{�©�O���6�/1X��*�)�+rO�3�ә�s^J�4�8�Lc�� FZ���D��8=ǜ7���rPn�Wb��1LX!5Ѳ�;��E��%(	���3������1�ڗ��L�����FV���d��T��$��q(��lI#��Q�XL
�U(�L��$I�U�HQIED��UTF؊j������d�����"h"g��������~?����~?���߱ESDQQ1QE1%Q�1�������EԸ��%?#M�������~?������~�_��f>Ǝ�QD��DSQILE!S�QET�UEL4���f"�"!��������1Su��TTEUL�Q�
������ryRU��h("�`���"�b��������
���&&�*��bj��&�A�!�����(�>ښg���1�������^�uu�D�U=g�Q��d52TUTQ�������
���&	b���OQ��f�&*��h���UL��TE\�m�d�ZJ")����11{�TML�B\���5�OF2MDT�MU)�1E�#KLTTS%%PRUUDSEQ{�UET�DM��QI���\��cpVU�:KЮ�T� ��S��=��\�P���O��ŷګv=Ulơ7{�1̃�rz3��Sk��l�Z��s;���5��@��a�[	�Ců�������&����� ���;D\��.��OiJ�}��k˽/�l�w�T�I�8ӌ���wX4r:�x���)	���W���xlm���>�7�6Z���B�7N�j� T��'W<��.�ܲëcNX���C)�H.s���v"mTt^mޑY������R��ʊi��c�Kc,�;&�0`�՞�!�@nM�)��7*Hm�r��;N�(��[�3#��DtQ�)ʃ�!�]������\,:.�Z��Ӽ8��Fe��>i�Uh��l���������T�9�W�g�!_=��`�<M�<e���b�$�Ѿ|�$�� ؎�%�@J�8�P���6դ�ŏ^�ڻFl`�ث4|AF"�v4���:Gs+J��I[�iؽ��fW\� �h�km,@�r��7vdb����āx��a=�{.�m��n�30-���ٯ�p�0u3nf�W(=85T���G�X�ۊ���Rّ��7�qeN)2�=A��nԻ�bb������<��1��K�$d�������z�� �AL�i�����Ys�b�L�!o3��lIMi�4s���D�ᬍ|�".���4�xx{�Oo7*W���_KW�W����K5���{���O� ]�iY��%A���Y>ݢ_ֆ�0�p��_�&T��3M,�ca�>��&7Et�ܥ��R�6}N~(��򋪋�u�L�y�+�ʾ$��,ʙ��k;Ts���ڮ�������j�����v��+��P�g�Y����"м]�g�[��Y����n�R�F��Yf��l��m�j�E�º.CI�z�.U5�9M��W&��27�q,���m#����ʊ�AL�=��l�wJ�|�<8��O(}2��+��jk{�@�����[�kp���t�����H��f�7M{Y������o_�#"w��xguv��hSo��ZZ�F�Y9Z��i��#��[;ٸ<��S��#�nB��y��E��a��K/37}F����Ҳ��l�3���v=�s���a��b�f�u0�7w�';Yۇ9��w0�Bm�\�M��(��hP�+!Tt̆p'i�ʚ{Yj���ؗ��T�V�N�_�~���mE��b�m>��R�����%�n e�F�:ÃACt�5��-кJ�Up�]��vFy�L��<=f�Z�3���y���Mr$ʴ��T|F=�l֜��7��y�0�T��}	9�����ܔ�ᮆݹ���0���d
�M�q{�6�L�_��o��\+v�Ev�jElvQ{�.�[%z&qT���0dնf�gyq#�Ɵ���*��ז��~w���볍���uQ��?Y�~Ui�~�lᇁ�Lr"��n�7]V����s���l=RK*���~��)G�[�S�c�� L�,K6�U@릥t�������N�fΘ���)�Z�_`c�!���F�ؔS�n̸#!�v�u�X:��g�5s�|�4�R�� �J��Y�R�.�5�{j�g�Y�%A�v-YUxS�l�I�1���wʷ��+��;X����[*�L����kE�j�1�H��"	پWɧQ��<Z�f���[H��N�SG>{��e�X����T�T��v���`�,����h�K�c'��]{b28�|c�i��F,�.���ә>�Ե-����Oj���ٮ�0y�%�*���fNʻ�+9������FQ�]��n=�I�JI�ܹo�;t!���L�C�"xA�X�4��bh�M�+�p抜2��6���^���{ƱotԤ���v��GO��E��J���g����k{I�u]�q�+�b�v��-�t���`(�-������ �a����7-���j�UaE,1��3M-s��A�1!��;�׵V��)h�庮���Wg�m3C�,�����v`����������#o]���������G��9�}��a�sc�YS���^�1j�>�o�:ë��4ɱ�{4���᪃�F	�W���5���m7J��:��Yz�5���1Ϫ�iş�'��L&�w�VS�^+���>�lR���Z^�c�a};����Ü�y��[�*̮3[V!�si	�	�`�'_C���+������忒�zs{���>�8�R��6��w
YNt��/��
�{����z�k��d#��g/*�Z�}c[E ������$�Ğ��LxЁ�n��t?�gCֶ��w!��5}�W2#���>�9Ӵ����<l%�4~oy�\l�g�٘	��׾��J �5�S��';3+ϧ]	���G��.����;S]�&5s�zP�ΌL�E��%7�b����R��\t{�-C������G�Ѕգv�!�����p�8�d7u�/�q6�h�wg���>���!t,���\u�[�VL�V�f��m���p��b�V2�n֫)�a������<'�#a[K+����)P�'�x��7n��=�5�kDH���Aj�psl��;^׎Jp�{Q���r��9ZOS�f�e���l��ove�EC,���eq���[��[*�k�8�{���a��6Iu�JhWz��uzx���;��`����71����ٮ�s:��޵>�%�Gʂs�Ǧ�⳨8?�����J"�t󝨞��-�Gu<�L�1hИ�׌Z�[��ڮ�,�EF!x`(����=z����s�#��j�Dc��x�\���{՞���k��Au�ϳ���"�D��Q3���o@tZd�7
�|87y^������~����'q�y�v�aq:�t�;A�w�[��-�ԜN�ـ/쿻�g׾p7�iG�J�SFH��TZ��t�� �uü�C�����ưm�E��ԲW^�
V��������}B�;�0C���q��s��6Q�4G�CCX	�*�[Zx��V���0bHvu�嚲�h�(p���ԇ�������֛mB.����}�����y]���1�əWP�E�ʡ[F4�Z��.����mG��XJU��Z�}8/��Qѻ��Iژjl�"�,�Sx�<eX��t���;W�c��u|1s����bp誮��=����(����*�Q}����+<�����bg�n.�l��T��nñ�R��M��ĕ׷*��Y��&Rjm4��������Y���J��>�$��x�_<¤���7U��X�;���/�obK� ��]�m�t�,�\�r���Ad-�5y��lu��Yث6���v3}�f:�Ҹ+���,�Qޣ�ten�Y�>v����>dk��c)�R�ph="�	W�i��E+�y@f�+"WT�y;�l�.��vo�����h32b��s�=,*�Q-��ޕĲ+c�;rk߿}�~k=n�=�3��=�Se6���A�_e���
��0w+�Z}ze����c3`}�s"��^��3}d�K=d�|H���s��;G^r�Y-f>ι�CK���l�W'm����ye�����<ຓ�V�o�j7J�+稩Z�1��/�{`���_����ӏ弝���b����u�� \lRS"�;���J|V��'g�x?�w.�v�Py���5) ���������O8��T5j�:�#/�����Y��f�Evg*��v�h[�M5���+G���S�pT���V�MNa�Z�����h�ue<�!L��ߧ�����c��h�Y�޾{�ȇʘ��5�^ /,�U��/u^x�8��g���hM�>��2�~��͍�&�Vh6"���-��D��ͧ}-\'z�ڗKƩ(��=h��ML���l���#�H���T0c���3;��$u-B���X���\�_�F��T�=�Q�9�������,y
���u�n,�2��yD��Zz!0�z�ˇ6�o��zi�S�0�Z��er9��)��`����"�Z[oc־������vP;}5}���'�{'�jn��oUX�-��ztO��v��w����Y}B�<�D6�Çg[����$Z�c5�Vf<�jWf�x�3b�f3p[�v�n_F��O�ᗆ�S�c�lo|޳���L(D˴#5�m..U�t\�:QrVd�S��V�[Ŏ�Ѧ�R�4yF�ӣ�4�⻯r#*)���x�����Js�x�z�n���ߒ+ag �2BUuBͼ ���
���N�rf���8:t����;�/5�]�]�|3a-�8���ko$R����&��|�E��m�^Y��K.���^'l�	آ�ţ���x*�)���]{D�D���p}ĭ�&w�1��B����(K@���*�7��m����nlul)h��=u��n<I��>>�K�+�|Y�{��K׭o�����C��{x�ww��X�E��ed�~.��_�:}�8-�d&��d��DE�ɥ[Zr�#iV�z(�)��V1�M�g;����.`QpaJv�x��*������X�Y�E�E!0���Nh��nx�śQ���\]�3e��
�fnR�E�k改m@K[�A�p͏�X-j��#%�u���@x �ΐ�\5y�����}b��Yzo)��� xP6!����Ѻ�GO�c���۹Oy��G�B��S[J���RI�o���F�4s\���f��
tmb7���2�t5I#
Ƨ!Z��C3)�q#�-ۜ�e�K9z)�;�.��٫\�Oz^�oj�#�Y��<�rlbW���JV2���7;%���ء������W�����=���̺��M  0 yc|nֶ��;_7e�\�t��`�[#�z�v-=�hյ�>t�LN��o���_��#�҆�*�\c����[�r/*^,W=�"6��jȩ襳�1r�(��� -���Td�/g�C�U2dA
������}Q��D.�j��ŞS/m4��
���zˁQ���jTF04[$6`B{��f�(�5����e{����x�w`ں�Y�*6��SR��ze�'�$�@SPR�_Sc�oV�[,�%C[y?Q��5wo�T[�F�;V�ǭ�oL��^jC�[Y��RЎ�'�ǃtN��
��ei����ݺ�M�i{���za�$� �u�ǽ8U�1��,�� �����.X�3E�I*�g�#ٌ~���5�i@'r}��P�^Vϙ���W-��&�a�\���m70�,�9���W���Er����{>� V	�
z")��~{"���]eJ}�~�:��������O�]-!�c-�H�h*�ab�ۻV��M�6�X+�����Q)��a����xu�3kt?�Zsw��ܙwH:�%7l�����(�S"����6*�}�e�Ѩt<�+�����4��)���C������CNzy:�V��� a�4clv���V����#1�n�����p@������w���c{��+�nO���%������2rl�I�L�W��	��R�7E�m�*Hm�X�]Ѩ���**�{���b�ߣ,oP~�����|�`, ]�X�/����6Hyޛ:i�Ӏ7bn=Y����A��:L�d~�W@yy5o��os%���F�
�P!�{����a�ټ%���0Vh���*�C��O$I����u�W��1X��\/;�\����Õ:�E�p�ӗ=w��@jl�b��YLR�U�3�ڰ�.�8H��P"�[Z �؁�׼���ƨ�R���p�@����yx{I\��@��-݆��~�9��Kko5$����k)�`{�h7_�����x>��`��-,����B����F���G� �.i�d���I��ظ\}D������jY�J�D�-j`�G.p�d�����y��9�%�[v�_]���s�5��r������:&BS�H�=��gt���%����9�h�p�h���Y�7d��S�m��k���J��43���9@#���;�G���Z;�K3����ӡ�K��qHi�M��pg"����u��q<�p��SAٵ�vQt�r�f]�ЅӬ���x�}ٽ}�s�2M�P~u6���ѥ�l�c7�]�u����;ѽV��������(W�M� ��|wy���>�@��Gu59��!=Q;GGL#��M��Wn:��̢�= 9lZŻLgg:=7;�����U��y���d���$!^f���zI��c����v�2���F�1�F:�6��6fףu�I�̈́���L��l\�7����j��$sk�za����J$^#:���7��x[Hk�M�X��J���:�����wv+�����r������O�C�1�Z�[j4�D�Ez�fM�Ԝ�K�l�̀f>*��.�"u�.�7R����kM�U���BQ��N-�0�I+�=�,�J��K�
JX���z/9X��J]pCՐf���i�λdb:��\s���T��B���,ᚷ� �<���e�L���	\����՜�f�]4#=z���*^6CBLK��WHw��#�S�e&�åe
E�fGiԆ��֖����V��'"�ʊ�y̥�91ʦl���#L;ZMw[\�r_+�u���6P��5��4{`�R���^K}S��]�
+^b��3RA@:S	������]h�ᕓU����+�A���ê�镘�Y*3zev�Ɉ�':�0-7YǢT��s/(QۮV��@#]�Gz�p��
h�\ y{��_=���\�`�(R���V����r� +�SCI2.�f���k����.�KG|]�*�z%,�dV��&
*9�k�0lGחUd�˴��{�V�(�n�;�rK�i�t��if��J*rk&Ն� n�s0��2Q��;k�F�^��iV�+Qs4�1��a��b�!�������<�zz��l2�k5���;V���>mZŶ.���eY�7n�BS���|�9�S�s]�V���i��E�1�ld���.Ir�]s6�ѯJӬ)h�R4D���6-®�?b2�vѦ�D��+L�qʼo3Qeq�8%n�ۈm�)3{�9o.�-IͲ���W�>�;dYr�f����r����@ƻ��1�.�!���X�(`��J[��;0i����uO���c�uI@��W�(5��h���ήEN�2���J�Y;����ӛ��'$�f���{/p`�������)��k��1MU��F�����F��8qi��W3A���o������~?����~�_�f�"(����U1EL6����$i*�����4UQ5Su�g����}�_������~?������ox<�L�1MGPj �Q�����}�AUSE5D2TLQAUzڦ64�5QS5BUG1�I+�f
I��$������j��h��"*#N������fJ���=g�A��4梚���a�*�ՌQT�m��D0ngu[��32ET$AM%USTiq%%��-QZ�E�/V���4z�*"��R�)�&j���*����5UE�ٝ.�4ii(99�(h)���nm4�T[&�X��&��TSU=FX����"�G\5PQE�1D17�
��("�!���Nv]�8a��L����c�
0޳��P�F����O+Pd�,�p<s3]����_�c�������d�y��qft;Ƌ���=���i�;�<璮�nT]�h,�0��:��M�H�T��>l�V��}�|60�<��ZQ�a�8��6��,|��2��3y0�D�6����J+���=X���Z�BA�^J�ж�Y���ͅ���ݍ�OQt�OϵK���]���������q�E"���t�8�P3OI���̇�����s2|v.<�)����y�����os﫩*"�e�qf7"t�����+��mEv>��W��D�`ȗxGd�^n���&�w3�ܺ��d��z��(5�곷t�"[;ٸ�6�WLv���d��&m�v��u'�m����<r���B���~�w��v� zVM�6r����
�״ו�v���z�wlq�/�w��2y�>�zx�&�o����<�lh��ĜoX�NM����n��Ȱ�ǻ���y٢塤E���j�u�G�K�E�gQ�������`Ӛ'�a��`�����y%�@�W��*i��B�y�L�Xι�vʷ{G5�������je�M_�*���)�d_n�T����6@�B�lf���i�30���;����]Y��������o7�y.��)�e)�.�ߟ]�<z��XV{Fy��"���ǉ ��2�X�/�Wz�s����?��*@�T�C9&��x<_Gu��/`�0+�w�2��ú������͛�E_p�Ox[�.��lO��(}��>j�})���^��)���Fp�c���f�H2�\r��mUz�?���j��jyU������Z��j��鋹��x7CRId%�Y��jP{9�uQ�Vq��d@����V��:�.���h��G�Gh�K+�<��ʚT��m�wz��G�N��?m�0�4Y���"u��z/m�z5>_l���w�"t�荀��j���Fٶq,`�'k��b�ųy%Vb� ����Ufs�����Z��{ے�Ԣ�v�P	��U���5K=<|w�(��!��QO?^�|Þ:��:�u���g��p����>�5(��n]#x�
1�B�fhYӓ:]no\�!^^�̻���^6�%���E%��eE�%�i�P�x�J1c�v�mI�z����=�*"6���L))C)��{{������A��Dr��z��Gf�FcDs��Ё�K��uR髃&��j]˹\�G\	n�%v\��	v ;���Ǐ��H�e$���v`�lߧ��̍H��GHwVZF<���|͉�2h�3�r_n�����&.0�YɓiS��":<��#5�B`^��~YR~�u��,��.�	-�v�k�v-#TF�\U�c�&��O��b��|h��`rjcwz��FI�!�E��m1-�Yp��/�׆@���ո����mUV�V��e9T'�h�����ݸ\]�_�t�� ̫MK.��+u��DH�-��F��ؖv�^3�TTT3�{��&�)V
6���h�ɰS7/���}V�D�✻<['�S3Ґ4˫�l2�kI�D�P�#w����!�:}j���j��(�(��sU6n*'(�V9��x�f�hA��"�9Czh=�H\��]���<J\^+�Ն*�/�J��s4Kc�'O��.��#v j��*���a'��؎47�.���ݕ����\�ڷN��m����=Ӭ.N�z�o�]���g-idg�BY�G��n�(,�^�B��tA�s�к_gwK��p;8��M��ֱ�a�ƶ_MG.�,�UEo(�@eZ�NaT�n���iw3�i�==���{�b����6޻��ެ�f��e�ׂx��"`�,�ki�/��Nɛ���������ls?b\ioYU�)VwUE���'����g��B P��S��v�ݖV��<�huƁwm��ҕ�z��z��xVFb��ה*�Dwdk�r��kP����l'_��(W��s�29��j��dC�ً�ۑ�r��ީ��Q�Z�[��x�����(�F!���y>�/���_����|�O�0U�V%S�s�޸ l��y/3��9�pW����^���P�hp����/��M\\�#�u�Ξsk�����ε������a������t�̷e|�@{�غ}��;Rso/"֠�[�8�L��C���gHq�<��Eд�����H����J͍B>��{��>�ո�W>l㕥�~We�{r]�)�����Nw��B�n��n8K�u[��[S7�������w)��T��?�䶮+���w�[3�@co%�M����l�p6	�oI϶��8q���Ǽ�	.Ci� %4��9�׊����ٗs��+���0��7=��o~������!W~l���~x������7�G�Ʈ��)#clb�==���|ͯ�̐����_����Yf���v�����ӕO��{	կ�
S��*ހ�Ԓ��H`yg���b�>޳5��� 7n�����1O�r����b^�r�+��=p���]0tE�7��7D�F5�E�K]���>ܭ��І�#�>T��ϫ�_gئҫ�U�Vc�K��[�5py�oDp�{����&X�	ҭ�WW<�
;����ʳK��dH;����@b3��ʴ!��l�p��@�������JW��sm,=+�`̉vFT{�x}�v��CgIw˕k���i�Y[�����_z���E#7�6��y���*;���ݨb�5����r���9	<^a�1�`�HF��{|�$���� ����cM�m�E1
��<�#Zfyd��mӘ��wp��Ԩ�n�cL��Ȏ�Nv����]���':;ٳ	�{��+�� X6�kN0ؕu�c��+iq+Ǽ'J{Wjt5;��fJ_)g4'f2����*�
]��bt�s�x�"�����별�Ӟ�}��{�V�iE԰y����ۇ�)n�{�Y~{��=�g���,�L=U��ܫ��!N��'&���ϭsd�3�����~�Tq57U'��{�a��%�i	�T�����Ű?��*}��I-!�)#���1f�v��6qc����Tz�tU�`k�gk��y=�,ǭ,m��	�{�8�Ό�С��ӥ:���\�f
�x�}��3"�Rf�wR�ͷ���uޗ:�S>h�Y���+��ug� XGK��7�&����E��&�[�d?��t���U&:]����)�;Bk$`h��xA���{u������V,w}��8E�����K�У2�,���Sp�B�ܕ�R�咕yf?�*��6��E�K���꩹�f]�aϚ�ڟ*��S��FZ���l%�R�+k#�Թ����;���^���p�m!�����v�=;�R�����Kl`W�(�s+��6�ϵ����GI��r�jo�~i��<}�_���ٺ$m����is�O2Vj�foL�n�/:���'Xv�7�+���eܯ�Bc��5ThZ�ߙ�ĉ��� @k�Ǉ���i�'S�rDl��������H�o�]��&
ٲ�|Zu�A��;�~���<��ؒ�vE��Wrc����{���I���Xz��on�m�ڥ';$cS��t�0�W|��D��9��ŷ��R+M�ȸ`trϋ5uZ��ϻe
ós�o������a�� ��2F�l>�-0�6t�,e+�к޻!;����U|j��I�ZwU�N8�Kb�^�X��cɐ*7kE��g���؈͘�����ekR�Ƭ5���^��}�w��� ��=��6�����P�@��hq�m`�i.�]��*���i�6m�i��ɀ3$9��@<�g�Yp�`�}�3���異[�-�np���+5�V�P7Ọ�,O�����Ck5���6�u�Z��}��c��idMK#���Ѡv��5M\�T-���3���n�"ݶ����|������7^1Ba|`��o��|g�n�����:�)�L��e�[�6��c��B()@���:��fVl]6uɣS�]%�ټ�Z�<�tB�s�;b�X�w��pІ͝�\nT��ʑ�.�1�x�>ǘ�fc32��y����BΒʣ;ގܺ��v��ϋx�x�6|K\{3F�u#�-�n���)��nf�fM��[\2�a�Δg���7�2�Q#���W��hx���������iu{�mA�ik9��3�Q5��
��r�t7�R��������끷/a=׈�A~B~j��S��>��Wo��+��@؎;8�t�k��J�mE���e�y;G&��j� U�M�*��G
�J�,��i-+�y"�c�{�����S�Kz�)_P��ձ��q˟6<Zf��mjkk��	&��RG%���eǁأ� ]�J����]�����
sN;L���5qI����#�q�_��0\�'�=o�U�9����ɘ��n��נw�K��=qC;�����{��h���G�˺��ޥvj�L��w������-o��W����቏:�"����W3{����%���s%��j}iL�qݑCo�@+כ��Zj`��^�2�q��y��a��z�]��쨎F�0�2��Q�l��C�i��Zɡ��ovueʌ!,ؾ��ޓl�v��1�e��b}�ja�Ӝ�7f�8���Թv�I�����,���&�2+�,Q�����5on--޼n����,:�d��L,�Ւ`d�N��~�\����$�k����w��an˺c���<6")��w��y�"�{��Y���m��-ǯC��hll6t��E��ɡ1wc{��bMNJ).���^�k�S�.�ŬG�TKEG*�n iJ���<���nǂ~�L�aa/�<t �[�~0�r�g��4��. w5x�=F-������f���}�O�0ag�J��<T�U��V����`QÍW����;�Za�o׊�[��)����g���e��2���}��+�ʝ̹�ї��m��k�mf�8A]�Ĭ�*���!]�-�N:o��bIG2��7�\3�k3^LR�]f웱�i�'|qVRUs3����ׁT0R���mS봼�-�����!��\gmW���s�F��78��Oigr̅���۫څ���/�j�%�����0����"_=8��Rv��-f!O��M����p�b�g�f8k��]aPN� �
� ݌���sc¾;:�m�����E�QcWt��:&]�q̵��Ƭj�lh���}��X�8���k�����������W����v:��W�{J��%o�t��9�A7�@�ӷ7;�~�b����m�'��"�@��i��#�i}���U���1X�H�ލ�m�����T5��rUθ�=��GCS��P�,�;K|��[ث��eJsk��� �'t�6�ub.l+ʲY�fÿ.��x#ĵ�U%��s���!��]�̥fVi������2U��k1��.ToS����ܖ�D�k�3��ߤ���lP�ퟪO|rX�r� 8�餒�ب'��#�1����	7*��~�F���:�1�շ��Q��*�){����_��ھ��y�<4i%�K
�أ�uPht6���Љ�"&�VqWo�;_�驕u/��3f�p�G�Y۶Y��_��ym��fy���_�����O��TUEw�A_�~?�H��QO�Q����D'��=��3"z��@�P!�a�eXaV@���aV@�U�@!�eV@��`@�U�!�eOl� �P!�`eV@�!�a�e � !�@�!�a�dBV �@!�d!�a@�P!�a�eXa@��d@�!�d3a�a�a�a�1��0�0�0Ȱ�0�0�0���0�<��2,220,2,00�0�2���ad`Xd`e`Y�s��<�� 6�D\2 2�2 2�0�2�0 28@ @@  � �T � � �A �P � � �T �� � �D � �A �`Pa	� ��i�@$"aed	�@��QeA�&Qa���Xbi�Xa`�P���!�I�`�!���ʰ�0� C �2�0�*�(�2�2�0 C ʰ����0{�=����EF`)T�?ð��������~��~o�������C�����_��/��__�ǿ�~/�DUE�?��?�j��+�����+�?�>�0���i�S����������~o�z8�������������?�~����@`AA@Y%!�� � � % a � &P �@ �@ � �� $! 	IF �� %$ P� ! �� �aX@� Q�	B!a $dB%$P!�	��	�
T1������������-"� ��*~�7��?��~B���pt��#��oʢ�+������}z�'���=Ï���c��:���QU��?�?�/���N�TW��Q_�C�a��?w�Ey���=�����?��L����������=Oנ�Т�+܇�~����ETW� �(����A��?n���Г������ETW��O��P��+����!�����$ ,��`�g������^�<�;2_�Т�+�=���̘���?���|_��<���P�#�Ϯ�E]���~}?����$���d�Me�xǼ�Uf�A@��̟\���yT�M%*� (U��J�$$P�QQB(�HR"�b*�"�ATB(������ٛei�
�I����MI�a��q��M U�f�X��A��5����m�cC33,��a6�,���:�f�(���U'l&fR�[fj��f�l;k�Z�SZ[i�&�l�R���k-����fl(�kQ�T
2�%%M��D��AM[,��[V���VY,��M��f��h׀  ��l&��r��-�u�)@U6���dh57l�
��en�v����媍U��*J��Vev�mJM�p(�����d	L�J���5m��n��m�  �xP�B�	$HL�����$(Q�d,�w�
(P�B��yxy
{�m2z�D]�n�vmi���nt)��ݭԥe�3�]:a�-��v�B��F�۵�,aE�Ubi�5��o  �{@*���j�����h��+L��a�6�ڪ�� 
�zʹC+��1ѝ-e[]�nu��)�� �J�*��5Ji������E-i!�[m6�� <)Mj�[�V�K����K��M`�ER���5RGF� WQ�4���@R-��QE*a\ԶEI�6U��j8W� ��(IN�v� ��;�GF�nn��P��
J�f�j8 �����lw:�4]pu4
���P;;%�6��-V�Z6��U��U� ��5׻�r��P��r��ۻ�������V��0jF�H
��J�ݠUQ��M���N�&������l�jL4�m�x  �CT!�L (��q�P�n�n ����(�m:�  & PsR�  �,�  ��  uRt[Zhڢ��*d��   ǀ  ���  ��� (ml  ���  �� �����5�ۀ ڻ�7f������ .����lm��%UP���   ��P ��:�
 Vf @��(  Uݜ 
k  .��  �w� wm� I°  -t3M
+YK6��Z�kY'x   ;ˇ� 5� su��  �u�Ҁ�� ��p  -%�   �X0@�9�� �O��)Q��S�0���C� T�5<�P  E?�
�  S�OFUJH� �OT�I�U)�@b3T�i���wq�QBFPX���LN@3�@x}�\0S���'ؾ��着����ľw��+U�m�5j�mm�j�km�}j����6�ֶͭ[m��������g�	H�%,$�Ԥ~��m���;����տ��h�{��}�Vv��b�jt���e���V�X.����V�K��n-X2��E[0&U��کD
.\�ã{��ZGn�7hU�N�����\�`ݖڸ�f��֮z+�_Q/��E��3n`���f�H��n�^Sٷ�q2��[I t��\�K6k0�wA�3JLYu�M�?m���lȑٲ��y���ƀ ̙�u\j�[<�ܢ�r^�E6)�m ̅BQQ���;�7�����x�4�ل��/V�oD?I�.�Q�t)��*��a�nR�a�1L��en9�d@�`*��h�Ie��V8%ܲ1��J2�
�F��,Y[�4�%+E,�V�5�桮�����!JVO�k-��� ���J��&��+�D����aHb��)RV���hn,�~ݒ��6��L}%�B���lf`+��Չ�-[��Y�����nC���3X0#4ExJ�~E�<�Y��9�����OQ�����;B�����*E�(ֻ&n6�bv훺����E�ߐ6j'����J)��r�ޅf��c]+ ��ʉ�j(b���h��%R���A���b�8����e��X*޹b1C��MYJ�����D�)ʽ�T6nT��!���~�Ŭ�nj@ɺ�Ǡ��c7�7i%%�����C�&��3�*��H-m$h�5�e�,��r�+�TI��[;���%f,R��Y�d��P֠ ���'�v�L[�,��ov԰$��E���[���)-U�%]����� MdҘ�p%u��/qZ�lPd���Y��;Y�/V9����֭ne��H8��`�.?�QCvբ��Tю��^�4����J��t���
]vE��]�x�b�1+��M��e��)�NEa�Y�,���܏c�߻w/�Yv�X	ax!9�)e[�v��*�����/N',;�H���Vj�R2F��P�hPc, �꽨L�ư�n=7������o>�J��5A(S6oL�7(�鲘�{���kheA��ͫy0T�N�Bf6uP*�)�� �)�� ����Vbв����x�c ]�+4��pXGT���o2K��u��L�{V��Uv�1�լu�k*�e��Znئe1!�X�5g�:���� ����n2�2��P���$c������L��|�33n ��Z���[�t�C[��JF쌠�q`���
�VpG�C@C���op�6�]�ug�����6��wn&g۫T��� FV�X1n���-H�bu��&I��k8�l�ܑ�v�T	訮��e���5Z�+vd�T����n۽�9V�`��5���I���ML��m���7N
6�k`�e9���9��i\��#&��n���B��J���ŋ[�D�n
&�I�bac��1���VS��6l�V2�9����K%�ܻ��!6ޝ���2م�KSV-��˺y.M��j"��(Z,7/El�7)�U��:̱1mZ�3NK���F5�dRM�����ie	�C��͹V���DFŚݍ*ѭx�@�@��˃�VJ������z���Z3�r+�:]��Cb/z(&�tQ��r�3�]Kj��7�P2�Mɥ��L��]��Ť��Ci�J�߯Nd�a����'�!�wn��ځЍ�Yl����W0�Jm�N���8�>�N/���ޱ���2���==��^�ú�F�:)	��]�^��-�J3öLn��mCX�5��ڛnf/��IwF]�׮�g���)�]��Vi���32�[+K�afe��l�w��ne^�u����sϺ�]�i�S]p(w+Ts/�m���坠�W2���M: T���2����n`j�Ȳ�i�fe�@4�Rm��{��F�ENS�X��0���hD�D��������[�7a
'��`�c�)�cv��y�$!9j�d�zbI,���� �]ꙭ��ygo�"�Q�Y���d�R�t�	�A7�����Bi#`OWǻ�3猘��xe���Sb�52���l��oL��*�mVX*�aP��d�k���^�	޺P�c2E��'a�{���b4����#kX�C���4�]6N�0�C������IJʬ���6ü���%ɿF+��2�P�c�:B�{.��`ުpЭ�hYw�:�F���^�%ɨ�U��5;��YH��ݨ�[g[/�"�R��q�j�Xc��A5{oFM�C�p2�*T�+re�sE\e'��NG�6��x+Q���i����PŴT�ԍi��]m���B˧Y���n��s��2�j��a
�6�T4�A�w4�-�mH(iM��/"ˎ�9B*��1Mɗ@\p	�����kWA!i��[��HCIP��^�#.k��.���%R;A��^����^C@�p�q�7R��%S�r�Ď �ˤ��Y��m,�)R&C�B�.mC�B��B]��5�[�-BD�e���� �<���P��B��^����X�w1` �B,Ӗ���:u��%��v9yu�����Ū��an;��ϐ���.'/u�~ �*����c̈Ӽ�@hl��iO/P��N�%�f�����+�*lwZr�%:����96��w	M����oS4�õr�S,�ڶU��z�Jn�U뒴^5���DC��$kk^��,y��de`��)WLԽ��,���9Z�Z���²�.䂎`�0]���o)�X/p$�4l�ZuXm�˗,eC�m��ua�:�ފ�U������CSh2�T��c��� _��R��1��(%S&�3v�ƴ]1K��R�H��wz�n��veLN�6��c(�C��-~؅�)@�ʄ$�Kv���J�;���v��Ŧ����qfXP:��J�7i&&�Ы��5,Ӳj�8������֐�$'4(��Y�Y�R�Egv&n,���Ɉ*���WF�)�e�͚Ȧ�� �n�Aˬ�����PǛ���r�d�lQ@`Xj�m�U�ZK(�F���j	���n7[k^Z�r�WC$���wX��!�f��H�S��4�30�AxYp��W�EYaf�����{���Q[4�Y���A��+uJ���`��ͷ�61ޣX��֪��ii����s2�$�:���V�n���"Ԋ�ʹ"Қ���S�7�4(h���흊�X�0�N3����d7�DB�t���KpФ@[���?m�2��-�K~�d�s*���2��r�nZ�A�&��TD?��3f`Qٌ�`��tL�)P!��
N÷������ݚ0�W�f�7��Ub�eFH�M�����
SS[��Y�d����,%�ݪ�+3�Dl�g~1�����$�R� Hr�]7���R��u��##Oun��)���䘵A����^\v�g$��W��MJD�f�=�VPX�(���n֌�4��\m��`R	��u�y��Igl��ˍGY� ��TX�7f��kd�%2,��
�ͳ�Q�3n�c`h�m��D�x�DͲ���ó ��VM�B��CE�wB�M`Md՛[D;1V"of7h����5�E]b8冝�H6±�e��#H��k*;������U�m�GCQU�%
x�ܘ�`�ۂQ�{�e8�n5a���L;��q��އV�`[YZ��)E�a���е'N��8r��L���;�fnE��&	�flw,&h�(�r�a��j��K	ڈiJ��6�+j�R��#@VҧjB����IK���ϐ����-f^�b���){n`��'ț�V�f��RÉS�N�����*LM�6���$�Kmc�P��&R��V�gu`v`���A�I��0I��k+BU�tP`U�ƍ�>'N�3�Ѥ�Wy��L�e<�&=J�kN�·c�v�Į���n�a�KV,�Mb����n�-�O��-�+i�3�h��O&��&��=����%5�a��I�	H��*(���֕E�rI��v�=w,d9j���ubhp��od��=%�QUZ���o�ɦKcm�x�t�{R7 I,�L�������U;��v&�4�l�X(*5�SU�	 ���fڭ�	��ɒ�Ǻ�����/IÃPiRlZ˘X��bZF�cʽ� *� �7]�,*�Y�nD�cY��y�^�
�]�a��j�ʽ�I7L����wH}��{�m8n\� 6eL&�1t����଑Z�o&��7n�M���w[M�	"lC>ܩh$�l�i�б/h�V̙%LdhJ5.��jx���S
���WH큆�5���i3n�+f���]`��P�6O�؀�)aA�s ��%��t��-"���Զo�F�U:��$��v^ ��wM}&%l�0Xۃ�-�B�@꼧	4V+LB�,�(�(�W�/p���٦�y�1)��J���+��B���X�N�ZV�5x���b�[��c͙5b�ȕ�[I�Ӭ����1�@�Mn��5C)��@���̦�B�{!5L��&���F��_אǯh��k ׿7�&�
�C�T��"�a��K6��&�� +� kk"2h#�o���ŋ5��jbb���5�fo�q��=�5�䭘�[�>ٗ���~��BH�M��A�.Z�����f���3e��7Uf�;D��������E�΄���Ks+U�IQ\˼�A�����]@&SU��W��)c��cS*^�6I��{���ҙI�P<dۄ;F�H��/]�qm�2�J/�N�*(�Y7w*��N��0�ʳ�l�Q���L�%����Ԍ9%(Q	kH�	�J����"��!�M�����j9r2D���J��k]�ӹP��2��Sqfn��/hZ�ځکX ����-���Ca,G���,*�A(�X���p;bdҢ?1*]�iYuk ���؎���h�v�mc���"Ean��:Y�FЙ�\׈A5�w� i���÷�8��`���c ���1�\�M53aD�ܢ6�HXbZ�i�R���4�/d��1��f̧SRt�y��61����HꛓV�uqK�ܧ�63���K-<�fee���m#�ɮ�i	�!8�@V� f��6�	\Ȳ�SOH�p���gUXd6:�$�Xzv���8,��M�Ӈ�A��n����	��J%Gג�h7W�y�e�Ԧ�X�t���{%�Oӿ�{��[-T��X84 ��X2���\����P(ŉ�ܻ�F$���v)�+���W�*��wr� ������3e�c^bD����Շ#�N�㫤���rPڸ��Dj�"�;�����Om�[���Tq�0�ͦ]F�L?�23.�+\q�{/Eh؎�H�v�j�CR ���É�)�{���Y���̭+E��TfX�XU��K���7JS�{gc�E
V�7�#�u��eԨ�6�Su�<kQ�Y�٥(Ӷ�g�ҰV�	��/�q]I�E����̓,�$÷���$	����j�u���)d����Cj��%7C��LSc�c�i{S7��p=M䳨�D�����`	˙�6�j���7��{���++%lA�Re���]G M����B��R̽�q���bU�/�T��T��z���Ւ}��MΗX]!|��/^0�7��+H���$7S��B�=Sw$fm'�l������X4��25�膝N�lu���e���<�n��bgs�{i����T-��]����d���^PBj�$����v �,�ǫ���^��m�C���ܨ@ r�d@M��7�]Ixi��YY1�q��$	��7E(�q���
�t�ܩ5�u6��)�+���^��.��b�-���=U�[�k��b���R�5�����U�dE�Y5�P�;N��DAa��M��z�:eh5NR�uj�Ba�\�����v�`�#p�h�v�U���T�6�c�5 v�07�Ǻ�<Ğ�����yI�/V���!
d�n���Yo`x�_۸�3�C5SY�f��Ҙ���w	+x���q�����:��mb�
�P�G�M&^칫3Ö�V6^HSq�镅�zb�ЙV	��Z��6ٵD8^��aK(n�/>�J[��<&,�-�&����hMD�۬5i[
wQ]�\،é��n��4�6f6������Kw/�n�
�ot� ��#��c{�Df��٥XP7-���	[�jiU7@�BQ�j��XMm���*9�NjZf��RD�qM-<�v�ę�r�h�����#P�f#W�@�*N�9�M�N@�|��O��0�������,VbV���d��+���6�b;�sr�< I���6thJ�0��5��_�I��F�8a���z�N]A�h��:�Xn�Z�틵�=*:�x���t�C�����Fy�"�;m֜�tG��F���F�T�W&&Ų�3ªP�	��i)]�Ӵ��)a�E���)��{Q
gj5��S.f�̻�7)�Q�`�"�< �Y���ˋ6�����R�N���BoJs��U��n��X蹗�
NX�ѷwA�Z��̩E���Y��&�p�P���L؀O0J�k-�V����-��4��[T�-����1^��V����+wMG\���sM�v�6�]��+hĖ��B�4��v���TɻD<����NTj��zE��2��)�]��V�zv3X�Ă�Z��X���sZ@);�;��4�3oPT�P	T@�۴��t˽ՅY�>�ttLQ��x�`"*�;(fdG# ����� [�ڪ���j1B����}{��?Q��[
ȷ���c��]��7wP�A;pҝz�Kʉ."򳺬�X�B�'7B��ܣ�1�Ҿ�+���(�jW<:7�g*sno�L��We2�.�w%O���~�.f)�T ��=�)�9�5js��� m��@�ø:��b2B]���޷��ԡ��V�`�n�lk->k�-G+���4�5�fT�˃Ӱ�*����L���&�J�:=�`9���wU�u��&a��]Wm9A2"W��F� K��
�k[�}/3
J�fڵx����訲D̙,����S@�w:\������vM���Y`��Ǯշd]R�i�����t6�����c;�m��i��n�����_um�U�4ڝK+Z�O��"؃1B+tSvp4O5��������MK[[3��Ь}ޛ��j��Or��pB�������Q�s���$�b��V�����<����wR��/�a�[�)Gju:R(��]*��(���sE�yz�Y���KW@��-P�i-�AҘ3�7��X�=���؞����W�e=��o�O��F�]u�z0NS^���ݤ*+3�M�2�¥19c�'�%$S� �]���J,v $[2�ܣ.P(1f��`ڮϞ�(N�)�U�+_ 2h���㒱,.��6��
�J�i^��c��� �ټ��ԝ�i�|����'LS��K��G�m\5/;�}1�	�j!d�i?6��wB*�c�+�T��i&��]�n�υ*����s1Fgz^q�G�^0�i�{�W!��z�u
F�!�Ot���}�1��#���*7g���gX����]O�anfJOq43�N�T���ܿ$iH�	C�Xk�.l�f01剴�/4W�s��p'�Q�]zR3�l��������]����ކ�9��׏��9����`Evw(��v輆�K�A�t�o.
p��F{J4M�vx�._e<����ۛ�$oY�AvD�F^�����i��ll%o*��	�(�0�S�ȲE�w�.#�pS���r���0�L�Y�Z������m�z3�z7�¸�:�c�U��w@m�Ou �SRӵ"�l@�P@e��u��d!5��Z�[4ۻ����e���}|��pN}噺v��7�U�{�^}��YϬ�Zo���e����rB&:��M����E�!��G׮&TӲ\��e+ѹ�������*ek�Cm@���dS���mX�¹ڗ���cc��@c��/C��Ir�Nӱ!�0��J��h��Gg �R�}�u�nB��3��;��=�rIa�L��Q��i�Gs6�!��_#�$���E	Nf��8�|
�#���m�׊^����I�bre�d���/8�,�Fv��&3z�_^Y�[}�m�k<�˺��ǯ�|��	���֎3�v��	�^1$�a�v���wy�7i�k;�j�(pyt� ���hǲScw��=V�Èh�TP�{�CR��4u��: ecg3_|D�c�;���$h ��˷K�h���n���ltu�wiH׼��t��&��\�^��@���\��\���6�}�n��v+��"�E!\^α�U��Фf뛽Eo>8�<�hmf@��N����nh���+�FC��:[�yܘ�	�+��	�$�M�����>��R|�r�pO����8�O7u{�����@������q�����go��j�uuedyAa{��Q���KL�Iݷr��ˋ=��(���h'���e�1k��Z�T�F݅I�dƲҔ)$Ď�[��e�I���as�%Pxw�Jmdo4:��1{'oHc�F��rݽ*���O�G(V��'�bܷ�ow�)�v:ʫ^��9
�Y4K���RX�+otl�18����G6�m2X��k���- 	�Z۵�u�����<�c8.TK��]t��HXr��ܘdܛ4>���f�$c��rm+@���(K����Hq�
b�6#��SA3�.���5�R�Z��f�i\�7'`0	�q�[�	���/�r|��<�~�s��:�ڜ>f�Zg���2�n!�w,zeR���~�ق�oǑN�\�pF¼�*dr�\+���S*Z��X�uU�H�����I�zu�:}|���ԩ3#y{��{6�",ئH���$0�|���9��i��ب�gА���-U�ٔ�/��=-�|m�v��mu���]^�{.촄r��|�cb��=6�Pyݕ���ũ�GW�OQOCC]N�J2�%����J��"�,Y>j��1��N�̩r:�]RH�geǅ¡�A�������r1Ұ^�"�ZB�u>��>Q�5��oinLB�+��i��t�ނ����͌K�()��
�un�;Ƭ�<������kgJ�:���* �'h�+'�����żw�[|����g���ǂC}�օpA�3ś�H����UofS@�M�	Fsv�7Qgl����1�ų�{�D̹˅��gS!�+�c��9�t�0y�[X�8�#���4[�QS]��}��|m�D�?o�!ٛ�iJ-Y��&9\GSYuj���馦��XsLR��n�r�wO�Cޜ[���ք��9�VRopv�8����*��d�Qά�����ቻhs�I�t�X2s�Jtooo��N�j����e����p��U��o��2���C�e�[Q*��Lwc��G�"����+�s��[�S��<'JV�Yt��˕lWyL®���/�
;y�,��Ti�k�9VeYw��3-]�T��fv�o`�U���uJ�Fd�X�y�P<���!�6�����fg%*�!�����w�Cu�˰�l
�e�9��9X��yV˭��Ł��IZ͠�ZA�E9P�|Z��{���Z�i˱�1Xl�c�O����-Űt��Y�y�g�{�d
ΡL�G�<&�Z7v�Z�k@t:���Ȏ�����_�LmZs[�n�ޒ)�w�:�q#�d��S[��&zﾹ�(&ō�)�k�f��kL�x�:?[dt�4��
��B2����X���^�ر��˹��2�ks�+X])5[�4k�}�V9g_`�^񝂠�f�'i�
�f��R۰��$9Kn���j -�Β�u6's� j�4��%���ˊ�YS3�kM�޸6�mr*���U;^��P�{HK켼�r=L`�o�yu�V�z�C�P������A�F�阃)WW^�����&h�K���+�������/��;���1� �v�b�(�Yo���C{�Q���UX�B�Tk^-�M��q�v�_[W/%[R�'�>��=�SO:�,M'}x�/o�����Y�=�7/�2�vfN#�۞���.xi&��Q�7M���)�_�︄�vI�8/R�4Bb�˪�w�3�m�Y��&5�mgm)� '��v�.��BĒ�k ���R�6Â�r�찲��֓F�#J!�eJ��'U%Z�c��U1"�Nr��֬��\�����[���5Ή��Nʾǩ��/�D��[O6 ���}�(��y��y�醦�\����c�E���qL�
bVc=����wZ#|�|vTF�o��� )gr}lc3s�)��>��Jb��^d���f�������Nƣ5���u�����F�Y��رC�'����&�`_w�A~cv[�x���KQ7Gb��A���C2Yukr�;��´��N4�������v�/�rQ�E;ás-�>]W�ր�3�.�ŮlI�/�b�����t��V��A�R*��s��a���Tr[h��o�x�k��7)=��3B�t��VMW*�	�F�\�X���Y���O5"S��X���0^Cm:;Sr��f��0wo�����ٵZ�:���Jd�5��wc�n�����x=R���>�nq�g�f�(E5���Z�5���ޛ�׳�}���bb�p��L���f
NX���_.���;�xӚ�Am���¾��̴���l��+���V��X4e��=|�铖�7*�s'uc�l)i=l͋O]�#f.�(M@���=���r�)�1�1s2�恓d�}y�:*�aM6�rbQ6ݝ��e�}���U�K��ƳLu���q�qW�}y6:�m����E��W��0�����VI�,6��j��:�K�]�:�����}����ͷյ�1��q�rXx���S^��A��� Q"@b>��y�*���s�r�Y�	�'����Y̓&�
	]�{.mՆh�h��juu��W��P�oe_i��t�*��o2A�<b�R��bՓ�؅���u�W�V�3M:Z�)�5�g��i��{�p��Gc�ä/:�u]i*����������7)pMM%���w����ȇ;�����o�id�{Lw�6���.��n�p������R.��Yv�����Ɏ��Rܳ��R�G�������ld�͖L��˒�Y/vI�}:J#��;8ظIn�l�:�wM�ﳯ�LVnlo���v��in=�&;�nT����"6��=�.Q�|ub:A]ۍ�رs	��£�..���s"�,#v�������XO� �K�;�f��(�N��KWf�F��o��u��U37�͡��,[�%:n�F�B��7l|��ΔUY����K��s7l��Y2�~�Aҥv;�f_?T��s�P�غ��3��!xЅ� l����^Ei��g�o��0]�L椒�]^7���z&�tCYW��ٔ�i˾@4r�wpқM�t�e���TV&˽@���ʷCi7}�Yy]s��|�ދ��h�Y�7J�2�x�"U�V$����]�E����Z-S�6ٹtZ4�LTfX�������9q'�e�|i����a�'��?X�4����s%X��|2ڽ�1cQq��n���*�)��%��HZ�TM?v�s8�+:�%�[u��!�9�k/h��E�Ts�'wO�.U/�3��&�y���=I��G/}2��%�Dr�u�Vx@-T����[���8����t��[Se��]3yHʐ#���s��f��ʛ���Zʠj�i���R���i��J���>�>��;�"'��եٯ�U�\ff���W���J�=�W�����ƛ�]�e�I����wk��b<D����!�KNG�í*���Z�gN���3��
�(R��r�s��nf��7G��/�� ��Xr��jU�Q�["�,�ε�8�ri|n��e��5.V������c_h��K�������:l���W2rV1!�;�T���>V��8�I�7�+1�>�ߍ��ؔY��ͷ�J�F�ؾ��_�ּ��΍L�tn�(����N�.�=��V>�-.�*�{��px��w��Ʋ���E�[��Gs���r�)��$��`��n�@+�|s��x��ܼ��^�Um@��Ɏ��W�.|�B�b�鸇V���������h��h���V����P�q�K{A�������{z�!�sC����dqÝv���tū/�n�־�&�Tq0�ָP<'e����ל$n�R)b 7(�.�Up!�.�r�҅��|�m3`r3K�� /+j��)pF+�[�I�ոz{Ժ=y+�:���TG�7����G��B��:�hFT��V��|�c]G�J���IqB?�$;���EI4z�n�{Ǻr�(J/3M���$��m.w^���}���қ����o+|�ܹ6�d5�¾*�����a���N���\�t��]6�����ݏm�7�s�$BbsF	r��ܡOp�.���S[��N�B��y@�X!a�YVۋ���C7ݮ�Y�����Z�ʍ:TOO$�	�f�z� �0U�u���/�N{��L�`�C7�Ǵ�=��T7]��fܾE�l:;y��7�K�W/�#qt*U�U���<�ge7������R>��`��m���^^'z�-�����y|������W�`�u�O]��]F�okC�n��i�b���zs�b�B+9��p�1x�;"�Z�Ύ�.��yt�;yvf<�bsK�j�S�gJ����žҲ�����9̥��]C�(�ݗ���A9���e7	H�͉A���I��F��O���g���坍=-Nޭ��ph���Y��2k�[������G^�gu7���V�#rN�1���D��g�/b�����)v �:$PZ(��Eu���E8�E���q`Il�Х��	�Օx)�d�$�a���E�@L�į-��4�A*���#��Lwnr���2!#�O�F��ozj�8����zmZ汢��t9	u)ܸ��̫����s��{�|'dXމh��n�uxM��|>G.��*;4Zsvؤ5*6��۳6��J�W?tP\�M�n
9nt���ǙZvKˇ������>*aY���{�bJ����rF|We�R��V{ݣLi9�0t���uLV��+/y���d7�I3���̬P�g�����*� ��vh�Bî�m��<�+EwatZ�f��e�/$�V���5��9��q8Vk�x �(d��{DS�k�s��Ux�k�W��v�t��qHiI��&R�.%K�Gx����E��3v\ڽp޾<��8D;F3˶m=_L2�nM���E��Z�ȎůT��g=�X+_]m�����p��ȥ�r0ީ����rM^���au�M���	ǼF�ɝ��i/��\{~!�y,I���]��h�|7��t>77W�g�ENo*[�pvɵ�̦���Gv��7Њ�`ɫ)���kU�sY\3t�xX��Cq��A^�mNs�M���&#��	2t�q�RxI���a/�HZ�]i�mV$��z�`m����l����=�8Y5�<;݄��b/�����8���΅[���o�.{w��PnR�p�S����}U��}�}���UU}_G�}��9��v���.�	Rb�Fw%��]�����/U�����.�8:�'1��XO2�5؊ɫe?��u�xu�3N>�жX�ڹ\r�e�(ϱ��k1�W*WF�R�U�i��iX,עv���&��M+���u�x�m�lG������7��VPX.�u�=��q�q�{��[�E����nL��l��[�;�O�p��Y�U���´����}��	Ó鷴Ĕ ���hZ����MN�d�y;��H:]�X����>o�;�)��M�.����l;��\p�2ʅR�X��:��C{�h����hR�z��Y����������%��l(�JԺD�e*VR��o����w��m���p���ɱ!s���-��śU7H�+�h]�oj��X��V;ku��ۖx�����Ő�`�(<�9wJz�M׌�4 9W�7����1*��E,姙��́,B��R�Ψ5�锋���-�k�O�ڴ�䈣�$!.�j/�r�}`�0�`l}��X�7kP����` �����9q�Z�����x���O5�o�7ș�s���eS���ٸ8��6��A��X�>��ou�q$;U3������ź+2:�)�1�1��ƨ9��!2����>�.�7y�4�������)��T-+�ɗK^��dP��J��A�ˌ�������as7&P���$F@���1D�m�4�ӫhe�6'Ī�YC����5qy2wUq���dtC.�?2)ԮԢ/P��RcV��*�F����K�������y�ʃ�`�� ��!�\���-�B���U0��]��:���@��z��E|5T�+�[��,�ٟ2�f��z|��N�2C<챎8�S�qo0f�����������6�䔆#�z�%O�rة4�;g8�跆�U�){�1J��W�T��N��'�ǭ"{OV.�΢��a�l	�b��ͣ��ӕ���6.�`�3L3g������Kӭx�\�9	�S�ⵌ��v]I.�n�J�AԶc�[5Ru����eB�؜�����m3:��q�4J��h�-��h�	�d�|҉��//+n�vW!��F%H�KVw�6�a��\�zA\;Z�.�\1t-)�|p2��G'<|�{b�ѣ7f��p��i� �=]�c+�����ɕ̶ĆM�Zӥ�թ����ۄ� �-c�듸�rv��w�%��+N�w�֎���<��ޤ����d���^�5\*���=.SK_PUc�81�5�7�f�f����F�s����<u�´��d|�,g^��By�ֺx���΁�g���J�P��7�y����U�'��Q���Ğʲ��܀�ye���tZ���S�&D��TPj��r����T��� �#���yc�w+�f��͌{w`�e»_m\hf
Ui�Za��l5uV������!;7��ۋ,�y�S4u��v��<��K^�Y�:�^������(`\�ou���Ô5�k/�2#Th$͸pV�1N�w��� �`���T�9����r�0j��e�I1�z���2��gN�Sq�T�vӴ��[z&�t6�Z9R�H��)-�?H�\Ǚ��2��c-��)��A�k.��b�Iڏ�Z+tٜ��kf�6)�Κ��%�(mvŷ\D��(k+�	��:�q����7"3:mc�s.�f4�,ݢ��x� b`dJ�+y-�T����0�1޳D�����Mk[;b��l�"�"��мxڋj�`��n�CN�#b�R��E��x9��Ariv�M��l���7Z�dnwj��>F�d
V�Mj)t:1t� WT��[tui��]��r�3h���tf5�F[�����gv�{�y��%ҥ�[
�W�R�D�i_R��YV�Vc���q��]0{B��+!"vb<X�Ǣ딗G6���1��hA%	���aÊE����`]Ӛu7)��'�R��M���.<��r�i*��w�[��$�����䎜��I������b��͘	��a�rR���ޜ�r�Z����U���7ז�Z���z���҅
0!(CV.���
d㿤�r�.ȴj�=������R>&%:��|�\)�kyA�Yt+r3��Ҫ{Փ�,t�y��� kM���@��×��]�����M�[���9�+���i���*7Kj��n��-�]�̇��8U�u���D�3�Hl=�0���ǃ�X�7���?�ǰ��.>��O��î�BY7,�X�w6�����έ����cYX;v�!F��up+��n�^�{{1_+؆L���bo�Ė���+}]K���뽝ئ�mu��	�f������k!��ۗ:,`��ZX�ڰ4��׋M>�+tv��9��Ӫ��4+����aTj��aڣ��i�4��
�vR��{�
�3�BT��66�;ڼ�v8�G����w8)x1�nS�Vk]
1h��>�����[,L���Z��@>]Y��.ȶ��B��V�ZȲ����v*��9q뺴���,���V�	����+�Zv�*T��J����\݅��<�bݔ����ބ���cަ]�9�z�:�؁V#�
�2n�*c�h,q$��zþ8��]�2�V���s[�C���R��,��^�.�}ԉ6��l�}ԅ����S�9V�߳bE��Jc*�Kj��t���� ;�C)`�b�����+A�����j�1��+V�u`�Q����k�t�;w��=5�9#}�6{7Va�U��[!�xt�G��� ���X�x#���I�>W�u[�ʰ�r����I�J�V�z��Pm�٠s�������Һ�(C��rK%2�=2���`���V_I]��ʜ�."��Ss"2�v���s@S``,�E��x	���s+5
ƞ<�ڮ�&���ڛ��É/S3��y(4452B���%�w���.�1g�-1W>W`�ާn������O���S��b���VS�Hg��\A+}Kgl&�}���Z��W��)a�[�Ӄ-qܗ�7���g�!��g<˺Su:U��@�6�7�gTj��an*k9^Q�C�V;S}֌�u�\���|��ԥFc����
�֤��y/O4Ŷ���ղ�K��ZN,�QNcޭ���㼰f�9�s�Of��aIp�
'��`y+Q�\�I���E%���ec����e��[�����䘝.'�&6�m�{�������ȶ���
�rJwY�;'� _e*�j��32����!b<"{;�w��霠��ږ v{*dhSڴ��86O�@H�}^lT�/�T��pn���-.�	ۦ{�U����s�y�,]��7�6@lfjm�b������:��W�o❅���=�f��@)e�Lc6�B>���UC��q��xX��V�N����,.�w��&�UjV�w�F�u:�ra��^���:g��E���m�
]���[Z���m��eև.C�=ړ��]���V���S�viZY�W�qe������k���|�7C�ء�=���յ��!?������WLA&v��i��&^���CZJ�Y�W�/(}m �}��Ψ��������]�U�%`vC�³5�\e;L%�4�֝�����`����O��
ATT�؟
�.�p�;������V�������4R;k\�jQ�W��Q�B�s�{x��F�s���uB5����i�|����΄���X����dV%��k�ᶢ�5�ώ&wΉ�0B��r����)�q%ݻ�9^Y���	�2�������v����Vև��sR���ŝ�� h(�
��Nb���SxvT��1���>}X��W��4��̱�;㒬`�pK��NE��z�+�[ڊ�DqR�y	�.'qtN�EDǎ�v�=v"�g�otř�_
��E��Uh����ؒ�l���6���a�;�Lָ��Xܺ(:][��>��haw5��Fo	����N;�&��4:�m�I���\����wf��^�IR9��� D�w^j�]K:��g!�6sV��yT�e%@*��]gb[�a�AY,��o�\2J"q^Sx`2�*zu�����
8�^ k�&�Zi����'��G�vM:;O�x*�n���7�����X٭�Ķ���!�{ƐL-�����7�11��G��K�9z�3�1�L��ԇi�+���hb�|f��.�;A� lA�Mo+3�r���kI2��%M��D��  ��lO��u9���6�&�5�V1�l8�?g"����M��,�<�/h�:kh�m6{q�Qԁ��d����f�ɠҭ�N�7p�&ob��t�	��܅[M�e뾔w
v_VR�Zt !xf�Rm9y�۠��,7� �b�}�Wi�v��܅�z�.B+�بtˮ���	�+��0a]|��g��	Q6��L�}�(�w�9ݥԾ%Q�RYE���Y�ҰgJ�v�-�H���z�^^�Ms���C]�%nn�}!��8�L0Q�*���-N�|/r�j��3Q7� �tY 1h@l��z3Ӱ�۫��[=u-���w��ED�������,sg�awq[�z�	��Eu����C )/4k��Ș&<�ދZY�q*i�]v/��mkb� w:E`�\T��C�nMJwf�����u�c0gu@6|^�7\�S�4��~���4h��������[(H��`f��ث[���'�������nb��]��I����dΰ$ی�TjP���nM!�b��9���.�%���+7����V}bor�I�Mg����@�A4V+\ �L��6�ڧ�UK|#�@껭m��lr�a�ӷ0�'�m��}�҅�Z�@�4]X��X���8�N���DT�󶇷س<�JD���{���u�dnԚ�w�F<B����h����.q�� :7q=��k,�a��`�d��k1MV���i��c\�Y�Ը�&�y*�0c'�(<b��y�շI�q]rkT[\�7ih`�摃�Y�k�L=��L�f�:[��I򮙎�D5׮5 �Y�n�(��\��;�+7�S��5�$��ܱ(1{��!t�H�/�g�e�ЈWU|���D[΍�r�FS�m9�*��֎������e=�����(_b7t�]���v��m��r��`�m<Y���7DZ��Y"�8^�SZ����5�,>�����9�c�E� 
]�u�l^I������e#tC���m�I:������=���[p�5��:z�$�GM�6�^q,�T�;��훼��Qz���T���w:U杻�7�_1��Gl�hYƂ���unaRa�v�gVb3�b�[ҨG�1]�ßubN�,�쨷��>�OP��;e�z�������4n�Q{
�B\\B����M��K�f�sͤ���>T�ϡN[k�R��VR���']S�vx�mQz��)կ"j[�g͝C2�۴i��;U�f�qub�ڕ�c%�:�v�h
�9���:a�(��k:�M=/sx�|�yI�N��ܣ��B�B�WHQ�ze�$)�A����b�[q�u7E*h�u���b���&��j�֝��T.3�IÒ��n�w�bX�9Gen�7B�F�n�'�e�Vn�����s��=W�ڵV�����Q��ņ�#q�:u;9�֒��̯<��N�������1����H��!�b�;q�^�t{�gwo��528-�	�E��0@&gZך�4D��;T\���Z��Y4��	����t/J5�pw����u�3�����p����<f|��[�춵We蜫E���ܮU��#��c/�k��ߊ)��{&���0[���oH��g9Bh�����!��v��ݩ:�Y����bx�M�=��)^��,����xo��]ʴ��e\v�3��t}��@h���5�f� ��@��^Kڱe�,�ؐfѨ3o3d���q�����dǍV<5�,f.��|���?��[c{��bV#M��Э�n��WJ���MV�!��)��r���*��r�di��뫵��9Mvh�J����2�t1c�\�� ��r���N�دm=5�ˮ�n�0U+���4�*��`�sC�J�ƫB��V��!�u	�����q�����,�c�2��Ʒ��u,�s����k|���or�gL��������i|��̩wA����Ɋ���tϛ�֌y��o@���-�&��lC�Jz��G)}��I޺���ܷ�<���R	�Zӽfu�K�nL��:�$7��]-�]-�<��>l�{	(�Vc�z�I�����Ime�4�7.� ^���,�z�d�g�ur٣�����E�.;v���F��[���WA^��V<�ڳ5�/�3��Z%u	̓yE��W��!�Vº��绐��Z�Z�7W��{��5�N$ܠO��Fh%�p�Y����q�[�Ww�ᩬ4B���-�Tgƴ]�Z�u1�ﯚ�G#��Z�@ӭ���XK2V*ٱk����[�se�3rb5
�8�+��Qb�SO%�ռ:�����Bz�^��D\��<���v�3��][E&jVH	h(˹���[# Ћu�6���5��]��YΉw6f��MGķ���9����;a�{��8�X��˦�ȕT�u�m��F8�����tt�/pT�b�����mB��V>�s\���%i2�[�O��m�b�|�k=�m
�႕� 	U���/��n�V�Ӧ�ta���2,����4Sَ�9W0,V���rv�ξǪ5̃Y����@��g��p�P}ki�/���o���X���)� �V�ݓ&4lS���iDڈ$��,��۵���WtU��q��u:��M5�mv���A0��S!�N�Z��ʳ�_UW��}��UOگ+Я'�X�E���L��\��Y�.�u̧���֙������z�SF��3i��u�g2�$�ẛ�Th�X���i��!9;}�Y6%�F����E��V��4M��Z��HK]�T72Z4x���Ӹ����c�+`I����۝1������H0��.F��L}�w۔�b��sl�"��k�J�8�`����Wgs�,�`����h�9lT��r�i�̔��9�d�;%*8�b��lP�c���3�S�o円8ݛ�i�F0qwgOc���੆fvM���FY�]Y6��*l���ˆ��lXo��c=���Hԣ�Ovƴ���q�SOpDHӦ��Vu��6.��u���{�+��gwP��4�m��ǣ��r�A������5�ʟ:F�J�W����\�<�x�;�A�u���Ş����2rr�<��_tU�a�xT����ޯ)�rnJ�"no;�
ǁ�1*�t�h��B��.��\/�x���yD�ǯz2\�R���Q�:8ɸ�ѻ�%c�t��`wr��Ս,Z����Y�z�6*P�b������l.�y�����OZ�&x_  �)ф+�L��ц�L`du��|nVw��I>z,?s��l��]�Hz���[����gj�'�����v�ĦVq��{S��xs	���QP��Z�]�ѢE;� am[�R`�����_߿���4I_˳I%2]�14F���@I��(H���((�Ҋ����Dd����guʂ((�!Q�(��d� ��ء�D̦
JJ#cF!6�F1���XB�wH�d�Pb��(��Ř$��IH�Dh�E�FP�`����Ed1�c�b
6*mt6�E��(%6�ƒ�5F��$���6��IDA"`�4��1�,�A&&�N�0�h)�,	I�%!2*
˖��R`�jFQ�,���(�@�JCIQ�E�1F�(�T���3�Jŋ(lF���h�r�0I*64l%�cl���{���^�������_�޿�?��Ú*���Т;1���4�gv显/H����p�~=A�W�r�ϑb-����Ǔ%�+���݊�������1�VG�B�+���R��B��Y(Q�@̤^]�u�MB�}�����ӔD-U"c�����l�s�x{��ܫ� TGsy����I�3St�ۯw`(h���@;1]?��I�jY+r�*:��Us��FJfb�F1}�"�tJ�e���p�jp��{��Bs���6��K�6x|��+�Q�A��*�R�TF�M��8Yj���糠�}P���G:ۊ4����-7��3�T�N��dV.�QSU[�s��q���2Ō����%���|�=� ku�^��7�X�ћ�ʮ�Sil(��p����y�W�&�U�l� Z�]t��tɆ-����.��nMz �L��}:�<�"���ynpj�����_�q?�����5o���f֠�O.)߷|���7w���x�*	��ٔ-Q~5�2)�[�@�{�S���0�<xv�C`h�-�L�w��1y·��C�)j��}Mf����}��(7��+��KS+�n�<B#�{��%L�;��ͽ��u�ܵ$ג���l�;r�}@�K�tl�m���8i�*�s��ܲ��7���)`���"ɓ�*+�zx�̑�`�m���3�"��G|^�tv���ΔnO5�1�JL���^@�:�"\S�l��l�
�'�����6ܾ7չ���u���лL�䞷���!�����|�A���w�/�\)WO<M�W���w bt����5t!��?y/��_>>'heϛ�h{ˡ�kG����.8H�V�#��P"�܀������Z�n%6L��p�w �bDBG�ȿ��xr	H������Q*f6'xlH^�E{#�\%���@��7��W�!I��`��<>2�p�@)����ă�[I�riV�.%��ڄ.=��#���@�:CL����Q��!��?�"�ܓ�:2��ǟ���h�U	S70����S���K�|��a�F�cM�l/���Oê��
ر(�R_��&&;e�|��b
ca�BLT=U�3@�z�țzd]��U�\ٜ�S�_u\�w�Mk�j�� *;��.͢. ���n����<�c�LC�����u4?�Q<_�$�c��zo�Ee+�;��{�w*�)'0��3�LV:���6>Q�3�F�]<;fX;W�Q9�F��k8{��C����k�%��q�'��}9+�S;r^V���s7���	#���=�+�ˆ��!��՞�VC0�C>�rvI}�+[�'�3`BV�ۻ���;'M�n-]d�Uk�r`�X���+4<z�5�����\������fYA�j"�޶��'�Y���{R,�?1T�7�z����<Xnx}an�*	U���=��B_^�UÜ�׺��ի?����N�KK<��z1��hZ��!��m8P��t��I�`�*H�����W���(�H�X97�gl�.hW'mY�S�d�h��g����(�ą۳M�����s��=����������&��B��=~�h�q���5� :���^UG;٥��0^8��ܽ7
��!��*�XvBwo�0���Ɉ�?8)WFenB�����ecw2V�<��X���G5\ʘA�vO`�]5�����A�+�܍�H��?tV�����&[�S��T�U��Dr8��طj�[uPB�2D@�7�� �/i�B�m�-�R�����#�hZ��1];J�f4G
����c� *��:�p��o����rѪ[��qSt�4p43Ұ���.{��y�V�0�	��D������,�tx��)�^J{��*��-YA��"N�˩�P�i3�Јv&�WY\!�rf���汻����3Egq���䷥"����u�ON,uYf���Gb���I|PUc��]��Ðm<}x�����t��ؔ�m�sdVa	ïu����1Nл�@-�D
8LV���X�τ��xP�*#w��ź�� �����E�J����k��n �qV]�7*?U���g�y>��Uo@�%W+�|��rUz�l�K��/;NJSRv�`AJ��h�0�x���O}1�d�f�f[	ij�C���D�8}��9��d8R������&�Q��A�/�:̪F�#��8��x~ԍ>�,�Gekc���<��z�ܭ��t��䣢����T�r	��S��\dЎu5@5o���g���qXFl�Φd*�2���8�oT�d^��G��Cpz�K�˥-o�7n�%5���k��E�ɘc8�kHz�[}m����u�_e0��yb�w���;YHn�.wxN�rb�:���|:�s8��2�+��(F�F����ncF:�Q]����������HEr����ġ�9��|��'��u��F����[�.��4����W&��g��vu�֋�=��l���d>�V���<|��;�iÜ*Pyޞ{Aik��)JF-�s��v��r�� q;�3qg��EB� {��;m�^�^����p��n���23��>����I�_�o���(K���K��]h:����e�ī5���/<���ېW�ټs��wh7:�Q�����8���zTP�(�8_j�ϫ���x/��S�4�睱�t�V@�"��H�U!ԪB�yfg>��rDePyѸб�%��\9�k䝤c!��3�~��	��'�ىHق�fK;.U�騌�xпh�����	��A���Y,uZ����ok���0��.�&ʓt!`��T�3�J��֫J�I��Q��:LH��@�1oL��oY>2#Q���� S��r��6稌�r��z�����.&@Zjؘ�][F����B&7��/������6�YGjؤ�e��4s�1`���P��Ёf�7Q_p�R��y�/�=����U�-VGCΪ�T��Ӈ�ʔ_vѢڐ7.�_�lg�咷 ��$1�s�g�f�ҥ�&#y�d熖o���L��t��O3>���b�����۸p�M���d��2 ��1l,�$td���1vu��B+�3YP���ytR�j���4��F���*uX�k�;�!H�zLޮsTD`ELhq^�,`�5�@�[������'���Z:�m�!:���$/Z��{oׅ����
=�D$�rNg�m���u(ʡ]�Ox_p��U�kvGª[�;s�6\X���Cis�<�vǆ<����~2�С�9c�.�@�6��]�����x���Ԭ{<��Of�Û;au/h��5;H�z��ӱ�#�̹6��c:Nĭ���sc} �!t�ߍ�W\��ٽ(��CQ�铡gvش�窗>
�ӯOK�S�e�N^}��:Ӥ�Y�)�uW�}_���x.j��6����a�!U����Y)���S-�_n��(h��G�dF�"�8�@l^������AY��}��		�Ū���zn!��������Ƌ�s���qkP�. ��V���ggnx�������K��ѱ��n_�V���a��h�f�G1��5âV��y�S�Z�}�зIV�&�׸�T·Z(\o6��:;N�9e<ǐ�e��6g&0A��Ȝsݯ"����3D�&zLdt��1���T.YQ�F§]��@�/:-��|�u*o{Cۭ��8�\dW:f�`!��#k��A[O�s/��[۲�,tr����ycN|�:���eh)��p*I��$Tt�P��_�;�3�S;�m�PhS�Q��;��J����E|�L1��q$��;�o,O*�Faq��&��>�~���(��O����Z�ui�E7-o֬�����Vvo\�rW��9����̣�*��U%Yb.�H���!Ԯ
���
؅�;X�6Ԇ�'~�S9�ݏ>�9Ujj�3:�r�܏���ռ���6ݙ\qEM��tSH�s�
1�e����T�.�Å�\b����;@ܜp��;9Ǖ�>|�pT�6�P��J��������WV�y�a6�%a"8s�H�5��8��Ev�$�6���P�0�;
r�%�d)�mP�OξF�AB��gK��Ɩ�"Fq�;_*���
�&��:�]B Loe0�9����O1k~�~[箎$�ߧ�����M�ީ+���E�(ڤ;��L����D�!�<uh!�>г]�R۩����iu�0��ȋ}ma�D�K2�Z�v�jE���*���;��AcA�}Y�Ui@K��:0_���/�\UÜ���n[ab�b���t���ϊ�no[ݹ�X��mLv��=���;]�qJF1�E&6����^�D�n��ÆÔ��cW��V9�ܽk�
�@8�1a'8�L�(�ąѦ[?Zj��x�q��2��,�r)\��.�)[���;4:,1O�'M�泈�*��rJ^��G	�X���ܱ��R�4�s�33m�-����|q�{�=����T���s�da�V���%[ۆ��A��ـ"UfХ��T9�n��;a��uw�F���d��I��TbGB���mݴγo9�SS"�S���R�o�H���w�2�[���"���@V��j�*C9K���K����wd�\+TL�q�vP��Y��|NA/&>��W@)G3���.;&�X�ȓ�t�+�ݘH�Q,�t��hej�uB=���;I�@���62-_D%w��:��飼rST�<����h�{k�T�q�7g�qb:y�Ӽk�Jr����h�W���ˈ:�o�Uuю�*�M�I;�1���7�;����%#Xv�B���>,*s�)�ͳ��wpjM:(��UN-�grȆ��|�p�|{ԣ��E��{��w�ᛐ%��~B�ul��>�b�n\�w�[��I��u���C:ǫ3�g�;]ʷO�nvMF�o�0r�,r2!�o.*jXa���^�,Z�lb3ႀ=ׂ
�:�?7�7��=����k��1m��� i�����Բ�[�5TQ�#CwUB�8o�z&��&|�]zl:��ٛZ|Z�}{��
������92�z�"�{j��3��r�<j�?y�aW+�\��Žjs����U܀}&�ۼއ%P�npV͑�n3��:U/�'����y�w_Js�����uWw�����s���� �q$�I#Ιt�)D�F\s`¹2y=���nvL��N��v�Ze)/nۍ�H��u)I�]xu����Β��\���/tv�OM�|��w���G蛝ģt�9�iz����e��s��vEs��'g�Ү�};e٪m���hĊ���H���27�����V��4�A^�p8(�=�Ɇ�t�2.g�ɖ!^�*1��=+�n���^;
@�*W	����ڣL�PO\�X�[����o��`�Q?���D\��n��9:��;�w�	�Zĥ�K|��.t�ϟS\�R	�Q� �|V�����
�:��iݷ��a��ަz�̹����c���޸y�l��D!�o�˦+z�"��D!_�;.*�=��Sj�0�s�{���� 8���/��A\6�'i�h*L�k��S�b�e�B�ɉ\i�n���\udQ�r�Zj*N"f聈�:\�q��U���)�g��{\T�k�����R�"c�O���t˴k=B���J�k��LM���\@(:IZE��SB+�t x�F�0�4w6w,l>S\���m�P���oi ;�
�j�lW�މ�#y�ap54�ӓ�`���;=�e�}@G[��T7��uB�c����mKds�x���|�T�Rh2Q�q�D���AiTG0d���7+n��p�w;}ˡS�n�F�=��?X�=s�O��m����۞vh��G��V���)>7�SF$|��ZZ��Z�5��̮\����Q�� ���W� f�*��F�n3$D6��J�*{�����:ϟ����g�������Mv���B�1��� FW؛Å��\���H���J܃,F��A���+��uDE��ͣ�kY<��&Q��e�.��'��_9��W��Q��UC�����|~����y�5�I�l��u��5������Δ��;��1��n�}Y���L'[��Ɨ��\3!8^C��Y�R����Y��,��,`�4qP�#e 8J _s�bs���Qح�O*3�88��_Hͳ6Zk��#�9���Ab�꧞C(p��lc§k�J���sNH��EϷ�C%�{��?s�F��c��:��IX������)x�\�Q�v��]V���ϩ�O敾9�yn�zk�����Ὢ��D��v�1z����|C�=}�����a�ƾ��� �xS)��LƇ�5r�9���B�Posۏ�8���V����aS,GDd��}�>x��pC�;��zk�V���َ��S��lgл~<�Z��/��vӈ����NE�enF�*�h�sj�����4=wj����������5qq �_v���	{�sS��D�W���=�9m�
�^lS���պ�pGZ7�*�VF�m�ZQ�[���g�6t��M�NkwKF�����I���؇Wxz�j��n�u�ŝ���-z��pw40�����C�&	��x�N�L;����X�Wcy��VC�n^$ѩ�2�D���P�5�<;q�X�[���Kt��7VtC���AU�D�]S^�z¡z%a�|;��oE�cv�R��j��k�X]AWN�N=Y�3s���0��
L<��[}��Z�����C2mb��r.Y�c�L�r,�}�ܮ��Vǣ�v��s�����;S��Y�M$����g��+��*t��ۮ	�j�Pt0�4.4��P��ףv���a�#��>+C�E����[}Bbv@�l=�Z��N���KɷP�4�[�ơ��ݚU�Ά��R�S#���A���}�*�豯��M�.)��S!4�Ҭ�f�L��Tʆ!|�5˼w25�ùI�v^���Li57��XqT2ED����&ڇm>7��㹽X���8�Ȕ=s6;�v��ŉT���)���� �m2� p���ݵ/�A�r�3����]3C�e�O)'U(V���c�q�gϼ��dte�76p-Da"��xa�5�M�t��n���5_[�QlB�#�.��d[z�&+�K_F�}[��:c���犈�g�t���^����� �Z�2�tf�m��erR�:�<�0�°��]v���+�f���F��o�K@�������{E�_UҊo��k7a��FR�C��������2������#�U��p̣C��N�F^67�*�2�3F�ztc��0�y[��ԀW���W֖����}��[����	��h���+Sp=0�<h��ǲ�#�r=}�3R\�-&mP,Zq^� �O$�5���b�=ו��"hœo�4��y�J�W5+���r��;K��'S	��m[�s��������nUc<D��,��i8�җ�)�G�����D�n91�>7��C�v^!H�M>+����ͺۮ�v�O�pGТ�e�/��iJ!8�z�αvJ337�g��9����\��_DƋ��r�Q���&�ȩ���Ὑ���Z�n`Ks��2���w��'�5���s��Z����[���Vkn����a��э��u ��G{G�����碔�v�.��t���B; ˕����P���]���XY�\\��[G�0�)�黼�[�u�*���2�ؒ����a���6����3�S,�r4��8KH�rJ�f��5�gd��ʽ���S�MJ�j{�
�O#���ʨ�R�&�k�;5gO!�¸u�v�U*�Q��i�v��xg]j�U���8d�9R=�"�/e�%;�gzh�eU��s[���U�0=�#�M]G����{	N�U��m_֖]tkQ0��>�(ɚ��1�>�	ɘ/:yxd�����W"[��(|+�C�,d����b�p��(��4F��DhLDTQIEE)���4d4lF�bɎb.r��6]ܢ��fb1�0�F�A�ء3N��d)�$�t����F4F+79��*K�,#�쌕N���1QL#cD��b��
 ؤě�$)E)F�X��LE�F��(�6�5DQb2I�h�ذ�R!D%�� 	4�1h����2��Ɖ2c���a6��`ؤ����sr�K	�,m����BA��3bM`���h*(���\"��@��"��3(s=�iS���K�.Z6\WV�;��k�����ҋ��٘b����:l��,tu������B�\Ѵ��"am�������r:��} |��^�yo�7�����y��o�����ί��W��_��׶�k��h���U�|W�W-¿���^���kO���{����nU�r������o���H�����Tw��ɱ���!���
�W�^}��<ſ��m��{����zm����~����h���^.W��U��Qo�����W�^�ڹ���������Ź\��W���@ G���9	��(�lm�������~+���W﮽(߯�x����-�W/�}�~���򹹷Ͼ����+���y�|�ڼW7���ҹ_��ܞ��x��w���ο��כ�b"�����h��tvt�*�:�}ʇ�Ezk�ſW����z�W�����������^փ^����-�\����~������{zk��������nno������{[�ͽ￾oCx�|�x����h���y����߃�DCD�����C"�T�����m�k��m�{s��O��-��O�_U�����oJ��?U��z�{���k�Ϟ^���~7�����^�%������m��Q���~y�꽷��^5}���!��#3T+�v�LzË����j���/�﮽��������{��*����+���^�x��W�r��w���~��K|W>���|�y��5x��w�Ͼ������o���ͽ.W��@��ި� }}"0��g��M�v47����S}���"G�g��"$k�~/������W���~�^ւ�W������+ţ����(�{o�����-��^=+��1o�湮�S#�"��"�������D��6��6��hz;ʏ5>���"$!�ލۨ�-�]������7������1^���[��_���+�_��_���/kF�����������h7�ί����\��\c������GF���� ��#�#�t�&���l�{��_�!P���"#��W�>��n��x��}�~-/��{�<�ռU�\����߽�9�[s_�;��K�߯���ž����������J��?����/�`����#LEx��`�����վ�ڍ�rM��!�'Єz�D�}#���5z~�9_����W�~7ּ^6���y���_��o����Š��{�~~z��~-�����z���6��ߋҽ-���m��-�W���;���o�s�?D|^�z*=&���x�՚���K��#x�W�Cz�dfe������2\���]ٮ�㵀h��BI� ֌��PU`�;wxލ���)>���nt��m��p�Z�P�m�N�Gg�ӝ�p��G��s��[�rmgo��+���������{{˳?�����_����z��}|zZ?������zo���Z-�꿿}_�_犿�;ҿ��x���^=�y����+��������x��j�����(��D|���}�W�JE?p�G�DFs���Q_/}��o�{k���տ��Z����W���zk/�<�6���|�_��������?<����n����ڷ�{ԕ�{R̿1�DH��G�?n^��W+�u�m�����/~�{U�sno^�y�_�x�+��������w������������~���~|�����.�W������͹���b�/���������ꙫ���az9q#�"CﶖTb1�z[���m��^֍����o�M��|��i-��^��-��u�|W��k���s7�y��|���h�Ay1��"�} xO�FV��]��S�8���E�>��z#�~"(D!��k�����nW+�n����^���o�����o~|�׊��ۼ��||zU�μo�ܹ_��W-�����D�����1�!>��M����}���Y����;x�<�} }b!��F��-��~{����/�������\�>-����~+�������ߋzW7/Ͽ|׵ʹo������\�>|�^?<�[�~�����/}�Hޛr����43�Q�'�8�z��rO�-����_n���w����??ݫ�}k��|�y|_�ѽ���^_����Ư����J�W-��_~�^9��x������ֿz\�����[�|{[Ź]�|�cx�����r��t��lM���C���#��1�������*����zF�\������^��o�����-�\�k������������~{|m���KG��?�_������ޕ��|�U@W�����_PURx�]�\���Y����.�����U���C�R�}�u^7�}W���=w⽭�^�;z���^-={�⿚�7����|^+���/�����o�����w���|W?�71��ׇ��l�X��|G����ۏNHK�Cî3w���1^��|D��A�~�E�����|^/m5��^�ޕ�_�ƿW�k�Ѿ+��o��+�~�Ţ����ޕ��+ƽ��׏�r���^�y~*��o�w忾z����Uϼ��F���Wz�hݼ�3��y�E�q�[+���H%ƽ�lQ��eo�e�,�ׁ��3A�V���z̀W��^>�b^����v���*r�L�5�w����c�F�]��"�f>}C:�3������Y\��K�d��A P��#����}�^�����w�|�^����x�}���ە���+ם��x5�y���߽��sǶ�Wƾ�_�����W��|~_�������m�v�m��o�U�3�秦���Vp�U�N>�,}DH���|���_��.k�}��zo���-��΍���[�~��{������?޵�ڿ�rߛ�E�6�s~5��ץ����o�ǝڋ|W=��������\�"�M�vL���2��|8z#�}H�_~���ۿ���M�~o���z���������o�z��_��o�^}����W����^-{��޵�zW�^*���|�wk�x+��{�W�����^�}C�]�wh�I�^���KzW+�}����sQo����M��{��W���_z����_��.W����W�|���/�5��Ϋҿ��^5������_�F����_�[���#�wȿ\������>B>��~��x�}v��ܣ�^4U�r�׵���m��U��x׃�o��o���5�������+�^��}W�������܍͹�����{o��o����z[���嗀O�(Y,�oFN������ ��5������/���}��y�[ǋ|���_��k����^�v����}^{u=�⯋���^����żk��ҽ6��7�~~��|�{W�G����������o��o��r�ٮ��~�㸆��$@C�����y^���_Ϳ=y�j-��{�}�zۗ��W+���~z�������o��n�����o]�h5%箯����|W��W�W����_��~^֍��U��ς�~΅�7z����¬QE�D!A}�������ߗ��+��_�o���y{U�r������������������[��|�꽷���|U��zW�������~{�o��r�{��{@ G���*��4�|�Pp��E����y��_���[�{Z7���ޕ�|W��.����[�r�W��|��ק�r�����[{U�r߷��W�����}_�����6��W=����O������9���۸��݄e��X���+�����nF�ߝ�o����ּ���[�����כ����������/�ž/�ŧ�����=���W���|��������^�����痥xP�$DBr8w)=���#q�ul�̎�K��:^f�c���ڕ�v�w�IB�薫�V1����Uh�r�ջ6S$S؅�_d�qo_�!�^'��9ѡ�/53�|��b�i{:Hmq�'�Z�Z�!��G��f���U�����:�
�2ܛ�O����=���������<�������71\���o�����[ڼU�μ}_[y���[��y�|^���7����}W/濿>|����ޛ����W��\�/�|[������"7�_E��}��0Z�;�ȩ�'S~ӷ��\w�">� �� z7�>`��G�}_��Ǌ����~���b��o�����^+ţ�u~����^v�>+���"�W�����|���6�o���}������梽=���={�U�mzr:���9���#�|d����)�~���?/�����Ѽm��~z�_[д�v�[��^5��/]�9���_��w��ܽ-�ί�����^5����[�r�W���-�~~�|���Ԏ��7G������}�O������ſw�}�\�5���ǋ|W.U�������~+��~|��}^ޛr7+ߝ�}Wv����E�+�z���h��Ez~x�y���s�yB���\>���}�*����;6o�� ��uZ"����d�ό�"C�j`{ni޳�/�����Y}���HN��q�︰���3��T�f*1�8�]��5GDq��:Bs�\m<�3��B��?��f3
���B+�f��?w[�b����U+<��L��McM/{��374W����0pT�W��:�X!|� �Q8iy\ T#
c,�g_^��\���ϋ_m�KU�w����w&��KU��� ��hxP{���[<U���T_+%��i���5S���薛�JŜR���}'Ρ���[����B�a�͍EF�W,1��-N8/�O�P��",Yv�Oiv��IgU��:�/K�:��E��+8j���W}�=�K+�UɅ��*�����g�awN���!Vjt�f9�J�gY
�/x�-�Z��"��_U�㇌�;����j����L[7���j�i���R���fX��Gc�������� !��\���r�6� :������gTSٖ~�1��ӝV; �)��Ź����0�rD��8�v�@Y���a�=@Bq3`Q|FE���^L������)�8��P�;�T�+]�z'���M�����e@n$G��8��<�ݔ#���B��_τ���mNaS6�BQ���\ �S���~H���Uu�Y8:QP�eG	A��6�a�<$L��:����ᮤ���lTCt��ρ���]4��6Oq��:~�B�v7���kG�_hs�Q��g����ր#��t@�J���P㢅�����|�c\�ʭL,&U`�;�gRb��o���3��9������T��;0����JF���9��$!Y#���䱛�p�ˢU����U*�~����P���&;gk�o�
�ɞ��V�i�5�7^�����U�"�,��\=7�%�d)��mP��X.��쩍��*p�56��Q�r_����z�Ud�{��4d�9���yHn�H�j���"G{��u��k�%����=��sդ�4z����dA���[�1���|�;���̮b�ĆnȏM�Xhcpn����9��]��Pf��ܶ��i�Ο}�}V�e�ks~�a��Ef�;fR>ӓ��uQ]��j��<p�pk{��:��r7�m���V�ŽXn�q�NO_�bF
���\��zs�'j�?�KV���Ѿ9N�1ӛ�z��>�uGM� ��si��5��A����kB|%�g��y+|/R��[ٙx�Q�I�Gs�;*��굫��m�v���Sy��a�S�FD�� �U�5uB�G�_cz*	��>��yT�C�?�/����ʫ��{NCVǼ{~~�D���+�p�V�˽dں�>�қ�!�L�i{OZޕ�ͦ���R�̇8��q)���=�q����럫vo����
�:�7�*��H��p���[���U�xXbo�M�1�D+#��OM�[�W�ζk���6��7A܁ד�bR�'2�F��.&�le���w6��M�wdl�1����*�\0,�/��x4���Ӏ���{��kJo�e��Ϸ9��JY0��=���K�㐜���c��_[�r.���"#�#�(��3���Z��s]��[,aS�q]rc��e��:}���t�a�k�%��J�Ш�n���Ni�wı�ymַͽA� ry�Y���N���K�t������]=�liWMe�a}"[5]������rΊ��>���	�\{n�����DD}�*a��͚�9�!�^���Ī+��l�9Ud��HJ��Z���9j�W���Y�Pw�R������C g����fc���ꕹ��'s7.b;��c�jH��%�8J�K&�KGMOۗ,���3�R��Di�6�H�%'V�J���}oC���Bwsg��8&�#�`t���_w��]%�9u�k0���d�aB��cB�U.��z�Nulor��( D`p��21���?5x �����}�i7�Ɠ�A[V�0|��C���;K�bAq�Q�[��a|�K#p��7�p�,����u2�a��\��uli��=�B&�8{U�Cf{�鈘�p���Q;�F6�~���L`�]��T;�=��:��9�ӣ@`N]1��M���
Ì�s�Ҁ�Ut���=
sJ�*���HC�e��
v���L5�C�qxFu�p�'g��J�U��Wlc�}�sʞ�^3�Xb�/r*�Q��V�O��-�ZV��3����g�>y�����6aQ���2������;[t���#U�T
D���?xk3-��Yʲ��&�I�4��Ȫ~���8�Au����[��>�|�����K� �F�²-��sc��:U #C��L���y͙S�F�[:p �.Q���j��*��%`[�(j��D}������r5������~`f�G���{���Er�`�E}Qc�@E(]��X%�`�$��lJ-oW�Yxn�3���p��Ь�Tc��2J+ �Hpe;�]]�ݫ�1}���M�FGD����\<�]6ph�7M�"��o$gݳH�$BY<�+x�(���3���0����ж���Qr�F/
�G�r�i�-��?`�w�r��T�k[�5.q�z������Ȁ�^D�P�'��9T�d�4�?��~��vnIo���Q���;��:yd5J�/[(Q�9*�*�:��1CC���1�
�Ko�b��ҸQ�wO;��8�K�eqlh.� }n�b/*���i��$au<*}��k��G��K�jD�y#�6]���W^��+���l��]e u7�X�D0�e���(���H�3�.y�԰%2\k����X�Q0��<8r*��&F�$�NYS�����e�G.��֪V"���9����q����ɨ��A�y��3ﱨ���on��3�8cc�$�8h��	¡�Ǎ�8�L� �k/����GΜ�k� �Vc��
7��#�m�H���-�M��Эj+I\���U�'�띥SX0E�`�!��{F`�[0RT��Cm� '�t�u��犧82�s����d�C��	;+��?���ꯪ�t��g�U� ���f*N�pp`vpH���f�n:�jE�^�]�j�����f*�v2߻U�w}ǰ��e7���a��-n-��a�>�|��:���3�qr�)WJ��,O��f�|�����F~�ڥ�5Y�cd
�yʷ~7�eq�=�bк���m'�٬��6��&�\�=��DOК����`��"��GI�ggh�u�+��RhU�/��e�����\"�4`����s��L0�}�j9�.��Ν���f�ƃ�݈::�[Xywe��0-���e��F���V8*�ju,�u��* wʍN����fvVMy�"c7|uv��� +�`
��"�W"�e���q�����m��Tj�]����pX��PT���F���G��CΒ�K�wǲ�g
�9j�O{��1�����+Vl�Qy�q�&xۂ�VS�c��5�Y�#D�.)�4�;��l���-�o���+����`��R�T+�$8u��r�@�dJ2�j9� �bDBEq�˳[s�9�{Eг��#|��2J�O*�þ�����[aN�0��q��M�`��:'�nj��p�����U�5:�,
��{A��=�҆��#ʽ� �w�r�v�r5�t�[��M48K��\����O-����q�m~3:wv*����i��ۂ+`�/�}�����2w?D	�D��D�L�f����� G[���D=C��th����UΉ�fRI�������9������o��M���Ҷ���חQ#��s�(��ԩm�I(�u�+�RB���g����7�4Lf%L��<'�@JZ�e�/�W��$�}~����O�uj>�h֍30�2����І;JyU���r��ʮ�Q4f�BY֪f$�-��׋h� Yf#�p����k��W���΃5u	�Ne:�fm�R�/xPq��pZ*O_�bAύ}Z�N�9�����5�o�b���2<��������*[� H�Rs�cOG;��׌�",=������K3�k���mK��*]�%
L��p����1�B�p6�7��c#����5�+a�F�W27F����lH��sǳ�](�:!tsPf�c�O��Vԛ�&�z�������m��b4@��3�����Ӧ�����Eĸ��Ã�%|eZ��d�Eq�[?&��Έ�S�6{(b�X�2t6�~�Ӂ�5�5��S�[ |��|庒ji�N/���M�-�{u�����F�t�T��0����r�Av������rOXф�v���n�I�u�Uq�7������o�:^�7�G1m��+������]�hͧ��Q�*vm]��s��|������m۴�ov�46�q�ǰ7��i�
f��U�r{/Q�e���Yxd���k`�T��Ӷ���N'���eY��L���05����1_/�qm�̾��R����ʽ<u1G��n�OZ��^c��X�a���&�!��R}f��4֪����6<�|H��z�*p���9�1��ϵ�y_.�QV����;s<3o�ټ/��I�����h���EN�}sx��s�ȦC����}7^U�T�QѮ�����ݧd�P6�ױa��J����|����N�"oٚ��ͳ�-S��|�f�Z�������d�:���pD���{����C����h��|�aj��kS���P� 圹��2�ppn]�I'j�lw�n����N�ݳ���j�c��A�ն��:ƎL��T�e.��|Moԝ_X���ٽ�[�4�T��vn�{�AД*	[�(>�:9��k}�+7��˹��Ax�r���#�3v�/i=��嘸�"	ib[׎��΅���ҥ�q.�hё�}l�MJ�'a���b_GL]���ɯ�=2��/��L�"�ȥ�"�)i�s)�W�&�O�M�h\8�H�`��;Y�k��[y�-!�Ǯ���n�1,ҫ��s-�*h*�^zV<}����E0����rR�F�]Wg$���PA�M}Զg)(�	�ݘ�Z��2th�ѳ��px>����t�r�X\Բ5��8i�p ��m
Z�ga�m�-��/u5��'�+ͼ�s��	��fn�qk@�|K�`[�o�7>��o#��k���^��+�H�J�I�x���;�uy���H�d�����[]ା�|������^ޞ�3$gD
���ݖ�)�E_4�rs{��ԗx��zPƴs�1���2\�4?H����Hv�5pn�Pj�������:W�a�t���� ʝ.q��	>�]�fr��|��e���5n���
�	(G}����y�fL���s���t����s[�ڳ���ʽs��P)Z�[���&�T�5��bŐ����,����Kt�:5�{�P���t�w,;x+�G4r���5�X�8�I"�)���;=!�v�k(d�.�'����ţrKO!O�̅6Mz�|p�Q������2[��a*Ky�w`���*�๢5�^��6z�#�iU��D=�(��4��R?4�_U۠�p^�0��L�g�]Næ�v��3(�]�tU�ic��^lЂ�!]�5�Ԙ[zƮwoy�m�}oz�&+��R��tU�+����V��u�v5n� aA��/h��,w�J��H;;��$�w(�����$�h��F6��wn�ˑ�����E!;�T��F�"�wWJ���I!b�m���q�EF�6�\�� �\4T���d���4j'v�P�	��A�L�*�\-��4I�QF�ܹ�b���u�(��J�h��x�,iO;W6�ŮF�,A�\�H�<��̨4m�EIFƄ�U��\��mDI�A��%���z��u�������n�3�o��m���ڱ�}ӱ�d�ζ�1��1־b��	�7�->��}�4?il���{v_?ﾯ����^5���M�T���Q��*W��|9��]�#Y�+p�c���o���AG%�B�0�X��紸�_B��`6:cm�����~Pҕq7�el�f܇��;f�\‡���p��]B�K����P��1WTV������e�xɞ��o6D� ���{sj6;��	S��d��l��p��E'U,Go~3Wj��6��	��S�����_��7q���X��Y�-��%X+D�y==�B���) qc>�+x��`��6!�鉎w�FE)�0C�ja��=���_�0y%��fi7���<���+((�i���f\�L�{�E���4���A�/a����� ��s*sn�a��-�7�)U��#�{�F�t<������3佧'�:�~�s�k
�S#f0L��
�%t��i̩4�a�!���w�N�l��X�&$���7. ̈́���B�ؠD�������,��
�K�c����o�e���d##���¹6u�eįì�|��/��í5u+���^�T[(��:'p���0,l��5(C	��*�KC�������U˄nJ�G�B�ef4���Uh���2���/\~4U�{H��	�ݗ��doi��x��qpf<��ϯx�+DV:�v�����Q@���������*���{��p�Ɠ��~�'	�AT�-�*�{L��x@�}��5�XfC�-ɚ�er�׺���M!�xY��][s���+��3�^�������\��+S+c=��V��qӀ銄���C|a
���1[����C΅��jq�X.��2.V�[Ԍ5n�vB{h,�TQ��'��LVZU�.����J��K¸�����G>���V��(&�OZ��`��G᳜�X����n�9��#r+踝u	N�U�w֩Ҳ�d-X�C$��j�#byu}z��{<�v;�8Z��$b{V#��(z\�����ۦPw�j_�f�ʈ�����H�4׺��"鳃D!�n1�P東�}ӔQY��ݵ�:ޡ9z{7��¡�ǐr�Ck�t�
��1aC��wRxٍ\�3���,ptv����ƢFȎ��\K1-��a=$g��S]�KQ��(Ƴ���ZG�9k��CiT�;/����,�R(��q�9ԢbFg���W>�xyUV�A��:x�����>���5e�1i�Wz�P���̪�n��(��y:�u��KR�qՇR ��Fi�\�`�A<��GB���oEཷ�()��=Nn��}]�٬oO�5D��W*�Dw�!:��>�+p�@Y�լ�)K�������難=������a��u�b�(��<��]�E�U���R@v<'�R!���'���j��9<S��L`�M
b��qˠ#� ��������v�� ��4�[�������N�vGWEȻ5�믷]0�Pn�9�����msx>@�����k ӄ=�w�3Ep���忺��g27�����
0V�z�0~��5�H´�w%f�F�T�i�d��2K�1�U\��X3_eB���ζ�}ʨ|u
���Pă�a�,��ڳ[��Mh���P�	B²��@�_nR�/x]+����JX���@p��Ё�8|�/��<5��3�H�7�M��lW9琖nq��r���-�t��p� +Fm����&��j��]o��k�������1Z�l���&@�q���kD���#x���9D��.�1�n���e�ܣ��"��(�7�;j��e���+���|݀�{ҽ-.??�����z��'OY���������l�TY���VhD��1B��s[��μn�k���u�]q��+�f.[X���I����5>��U������2(������U������Lq��_���	�@un�@r���+;q��O.�k�r��]�;q<Ck;L�4VjW��A��u\��[R
�������/���y�yK��g�L�j��� �k4�_#�j�y�[���/���	=Ɣ	��ɮ��e���֥�Y�����>��y�C�*ᤸwܲ�
]h�f���m,�ِ�Nvn%2�>q�'��A`�N�CӬ�ׇ�|O@Y3�c:Xr	��vM�D��%V��:��B/�:H�P!E��0R��66�X�
˪�Rf�q^O�^e)�:
U�G1���]���7�h=�ހ"����REt�xC`��rU7�f7�pl|~��xsh�%a�����P����5&��:�y`u�e�4��Y�a�u�ifb�뉺b-���F)�w8�����3s�s��K�jh�Sԓ��)(��u$��K���#Z0�]�V��:��uXxa4�?�i��u���ڏc�\1^e.���s�A@;g"Oq۝����~ɇ��y`(�?ce�H2{1�]h����:�������H������N��'�=�@�M��ۇ�c�	��b���9�X.�ң�1�?+�PسI�sW�jf+��P[\/l�7���knM���ta�2Wu�ch�5v����-�=���nt��j��t�_����e��;�d��wn�U�sw���͸��ʉw��+pj���_oT}���|%5:�s�����ٿ�j��2�N�s�w�C+:h_�΍�N���N�&��=Yq�fF;]���25J��+�^��f�t�q��p0Z;�������8#A۴��h�w`�\���6ϩZ�AD�����*�#�oا��V�E#�U��*S�Sì�}7�����彿{z��(p�]�R���}0�����2���z����-���\��]$�g�|��'n�O�������?(�ba��NER��"��&c�X�W���-���C�X�U�<t�/��2��*���|�1��u<LGeD��J�����-y��1'w\�40vI\�:�A�ڇЋ�Bމcw]��;�b�:r�+>SPO �ݮ�u��v��#��*����ߘ�89\^��E@�����.��|����'��)Vn�Q��U6Xn:�ok\a���0W��bD�zW�v��L�r46y���m�҄.e}��U�g3/l�Q#n@q��z�h��*U���S�^!��5 B1���T��\Ӫ[Zj ��U���
�������0����E���1!�5f��p"�D��2'g
=ku}�V)h7�m*4��=Μ���y�ǏR`�l��/+1N��.�:� �.c��F]�\���TN�ǀ�5l̫�8]��8����������=���*\K�R�U������O��6�qأ�!�5o���xfX\,�IX/C�ΚkYޕ=m�W���i�k�yO����ꕾ�zK�rR��g���}�jtK^o�p��;֝����".\Gu��iئ"O��
��
0@�1�J�l&cpܓ.��E:�U�����0S�U�k�w6�d�!9�#Cs0�,����0�fo���K����/R���b$F
v�ó����7�gLD��;�ٜG�h�.��˸��!n��v�؝����Nsr��bՆ4h���i����(�1�WU����Uu�\〵�$�{�:�����'\Ͼ�bk6����$f�>{p�'g��ү���ǧiM��z�`�)�˰���� ��4+�x�~�yq{�(�����F�jf4:�3���{�5G��|���	�|lGw:z\k�c1�1�������v=z��������6�&m��{U���!ɞ����\eTr7˯끨�7g���wLp�Wֆ|�(��N��1�n��%�˞Z/{"�]���!���W/U�=qI6]� �T��XuX��Q[�˶�ˡIV���U���3tdN���q
�3�c#l��e��<ڶt&ޢ4v�y���bT�e�2M������J!�G��7d��jì� �2]?ꪯ����G�������Q�&��&���1#��$��\�\�Ct�(D��x�i�h;��Y��7�{�SK7XH�H=�hy���.�(u)�k䝤c
�9�vogiN=��LO�s���䡑����[�KYd�ٳʼ$�^����v�'�\+L�Q�G�s��]�ߩ·��I��Ɋ��q5��G���R�󏉤���	\c6����=������U�%d�tk��ϝ*�X@�u�s�d�U��ˤ��/��j��ꊜ�ș���WT_�aی5G0X�oj�ϔ�:�t ���)k�(��K��;eu�����!TZ��Q^�E#9"�ڝ�6��9�E�`��_>�.2��mh%�b�IH�$h�y_*�����4��'ۻ�3������T.�۫���K��7Z���_��fi���i�
��0!]�X3_eBb;��0�F�&�K���S�]35^��ck��zg3�Q��y(֋j�pp�
�a����W�<���ᓥm�
{k����Dk�Z�gT����_%�p����'��̸.�g=Ʊ0 ��k����+�r�:�+]�����`O+�����Zt����ù:�Ϟ����'Sv��;��J	���ǹ����鑐8��w`���WD�S��䱧��jZqAW�I�;���yJ:��DG�G��K�����=1z@��7���s�^��F��`�{O}%�|����Q
���+������Bߵ(B��p4���!�Y,1���'|)��F������_&qT�2x���G�-��~�B~�)p�#��}�/;|s��-������"����=��Wq�#:����jY��8?������@�u�G�ܘ(�Ft��8�)�g��1�Ud����!�6�OJWq��㞾d>'H.�.SY�8���Y<>w��-{w�+
N�C�e��}�ҕ���v�\���Y�}as#jHnf�j�2�em���NuMN����q����yW'�_��|XyҨc�3_(!"@W�]F9V[jD-��'1I�%.8&�q�	Sˎ��=	� F2f��M�7A��e.v�^Lu���*�m ଧ�>%#��~b~�.&�]P��A\� "a�2W5�+��ν��kd���s#��!�(eA��Ù �wNA+$�|�L1��q$��;/L`�;�iU�Kk�B��Օ)���T���l���;܀G�����R�r�li�zX�:����	3�l]�����=�4��iGUW�7�e�����ݗ��>M���_m]>�ӂ��EKh�z��D}�}\ž�V�H���/�*��⏅?��f��ʥ���x[�ɮu����	~r<�՝�kl��s�v~�'M�/�I��.Jӑ&8mMT.�ʌ
�.X�4�D���w���M��J"h1�6b�5BLT5?:F�A�	�$w9?>��0�&�+��|b�6�q�����ƀ)���&���צ�ۿy-�Á�~��<�"�'6���X.˧��+�2���唯~C�vn3m #%H	9��u�-��"��0:�[Xi+V�v|F�k��D/����V�;�%��������钙�g�>u������NEw�)%+��������`"�q;=-,򩜇b_]Gj����+��N���d��$܈�>�O�m��� ��(%�\U���8����z���v�Q��Q��ab�s�E^���qK��9�Ƨ��[r���Q�
�f�M�|�i����0[Q��]sp��^�'
v�c>�0^8���*���	�cj!���&�l��;���z�th��=jъ��lK�<�W=���RF��i]w5�.3B�D�P6�ˆz��Zb�Q�Z�赻F��^.��7��r�W"6���
�;:)$��d;a��{�]�ͦ�u��P���\��؊�O't������ #��R��p�Xpχ��������N����&��?��enB��
�{P��]G��^���v��04�Wt���d������QJ��""��_�/��ڄ�K��"5�8���W"�ļpM�=<T_ZS2�t��&�挀�9�؊��|b�5e3�{�S��l�9��"è�{Z�;�W�лQ�4B4�7r�SʧD�8m}
�o�G��ʼ,O��٩B�E�憐m�uZ����j�:��*ɇ�ޙ(�o���O��7H��?��^&�ϵ���j�/�Õ4q�5u�%۳�Pt�F��z��*17x�D=�#�p��|ٮ%�9>Q�m���V�f���lPJWys�s�T�l�5���1p��A5 =⪆���c愞1D��L=��{r���@���t6��ojO}�#D��L��f[�QdY��hnf3g�_ׯx���m[��Pa����$Wu<�~�V��Q�������J���ֲ���մ5��u+��s������fw MXmp�i��Qx;7�c���@uƫ���qY��Wu:P�pk��U��_rX�f��j�{2�l���D���Ȯ*�eŎP�qqo�����F��+偂`�|�K�@�Z�T���w���Q<G�Qrf^L��=HW[���E����%�GҎ���+�;	e�#���s�t�B�;�f�S�Fֿmmm�SBu�i��y�k]�A��Ж6�
���K��h���dҵ��]��S'clc��j'f�)���񒥛qB��5�-�jJխnq{ˆn]�fv�`5\�are�8v�����^t��i
䚢'���[�^+r[s����p��O��\D��Y�J�p��"�T��QKB��C����p��ݥ���/!Z����-cݤ���3]��C��7�xdy}��3%�t�<�_$��x�u�mY
���of�\�K�WI({��ݕ���s�#9��e%�_C��{x�9���h�Yχ�zVA��ey47o�s��9{L��`��:Q�,�W�a�ձ���+x��b�p$ʆe�+Y����צ*#�;D�[z�"�m�77�OP�k�wjR_�+9��f����:�Y�+�z�b�'���^v�0� ���ܧr��m�F5�"�����W�-�#om*�*W>K._[�U=�.�ͯZwJ��O�y�|�6�ڻ}D�=ٿ^8�9��.'���w�uXa�1n��<W2u�m����@�\2�� ����Ċ� Й0%�Gbl��%�j��Ե^���e�E;���59�����%k�����[��:�a*g�×K`���9N�i�3��tz0�{��z��+X�3o�<�$��4�/<j��+�TՃ]CA�Y�+2�G�� *m[�9�g�� u�V�@m�d:�����wWMSk�Ζ�G�z��Zꇪ�u�ESbZ r�/D볬���5�]��r��IP1�H,��؞5�fne:#�QK�1��VV:1��f����p����.S�q	�xNcݡ��}sx��G���� D\N��)i���n�.%���_$)~ۧB��zJ��7����U�tyɂow\�E�jVV�L���-�v-}r��&.���B��{!����}�PӡW������ôc����&���I�.��2����f�0����Ϋw�mҳ��o�f��rf	�cY�Gs䋬�X��Xގ����'�R�!㩸�q6���2_?�^e�����F�|Q�t�[��ŷ�p�F�_]�,�Ag`�� :�3u-�.ۆ����;Y}��]��Ob�@�.�5y�<����Ν������X	:��ۥ�^�����s{�i��ju��%z
�熆�9�j����QC9z��k����xX��fi�)k�XFIZo�U�u3N�;�=�2��}�%�H^&=��5�uv�p	V��y���I�ؙ�I��#�����k��(��~*�ۻ�0�
�ІŘTPTE�F��ݭ �ƭ�r�LF-�EF5�®]*,(���� (�+��K&��eͫ���IE����6�Q���sE�F� E���wm��X��ѱ���4r�X6ME����,s��[��#b���1���r��]���'�}Ol�eGV�rA�*�N��e�r�/��|1�$oB���P=��6�2����5ک��sz��aC�Z�g�W�}UT���'Vy?nb��?����q\��
���-�pz�C��r�n/&a��R.�pDM	}
��νcPo2�東 TZ��:<1���kl��	H�#r&a3_����)�r��l�nL<ݍhR�Ԭ�tBlãq���F�Q�r!�1֪��؞�g���r�N|r�����۹���lj$.*�2�9��yu��/NF�L�dT��B��C#�(���[uΚ����<��YvFߊ�7����Ω3�z�H�5>�y�l��n�e���rӹ��6�L������"���8�ۍ���q��<5�с:�3�[q0�ў[f7�Jhh������,B���rPȍ��F��B2���6��;+�P�����tzv���1�(�'/��/N��qS��ic(�e)D�|؉��uH�����@���3J�U�*��&�gg�\=�%���Њ�S�����̸����V�$��'*I�V�v�� �;=Wt�Y.J<�F���0�do1L[}V�.@��(`���)e����,��1�]I� mZf}��Lxw�L.hw�n�N���eG�\��4'��\���1�N1�V�<9��V���!�/�a�~C����!�y95�W̞��MAb7�Kk��s#1��av��Z�SP�SYP_e�SEjT���eZP���2�t쥸�W6a\����)B6}��i�ۜ��F�^3�
�[#�爺��>fw*��o��{��>j@l�dX�0��T�e�L�{��dp�.'��p���ܷ�?�����)n�D'��_9��s[ـ��V+����&��[�>��n���ο�$�"�`�eB��8�\�i���8�+qQ�o�j�U{��3m��
U��"�K�[���xJ�^����T���:�s���T9�D
���29֎�}��xk��Mw���Ȫ��1&�GB��2z*�t)2�s����i������L�c��Oo�_��z�c�[ݹ����1�n[�!s���o��φ:�I�j�\>��b<�]��o�|�a�����̡��a	�e�;鹆���ݎX�؈C�ƃ��o�M�W2��f5��޼�')���Po#����aZ�2��<̮��l����k+6@�O#����e�B����O�K�|�U+_l+pk,S�+�
���i�-9|mU���f�Z'�[mf�-���"��:^l�:�݌-4�Ph`�����W0�F��t;�ࢎ�[!X��{.�*^{ư���ѹr2�婜�,�}����]Eʄ�+F��^��e�S�
ף8+�%Wv4��BA��7���U�sO؎K�	���/q��T%{��u�6*=�}�}�j�s��m�Bܭ.5�����;� Ʉ��;9�S�@:�Gvh�&�3ٷ�W%�����E��.	�:�*,��#aS���&9EC4���雅�d3خD\멺��̹�[�5�b%�t��Ĵwr O�O�˺�nT6l�����ր"�IG���T��jc�\����rC�X��|x|eN�̈3�p��&'��a���\�̚=uO"���]��lkHl$kt}�`R˨�����6�S��G����W�ZW��5z�z�=ʵ|�r)C��P�Ѿ50�\��n)v���e�u�^G��#Z1�n�g���Ycd�77�0�2�{x��덾�j��4��`�LW7@����̂-��4	>���B����]v�#{��B�=/���Px�]<�]C o�2x�X�v���#���5ĝ7s/����ɳ���r���B��C�f� Pε@_'P�9��3zd&H�@k����R���Sn�{׹ېUٽ#Ջ:�Z�B���b�xmWL�[s��*�q�_7p���\]C�݃�!(G�V��vR��=����{ ءD���6oq13�uLJU����v6��cT�I��|*m�gGE���k�]�>6C
|˭���8qs�BG|;]v�ފKٓ�n�z��|#�z;/�z�+M��䲤n���4ty�����*��q�U�}�u�$=���KJ�Ż�&�k���#�iV\#]�׻���lჅ��2�P�7�*��8Bo�}i{O�/e�3CP�[��n��yZ���0�q��T����|nz����C����puB��M�5�@U�fB��
�}{�n�o��:�����t��/ ��r/0�=�m��U�|Ҡx ^�e�R�7�����R0*,�-f��%[ۆ��A�(f8�`h�������*r�%�	�uBÊ��\v���%�*$�CgA���/r6�#Q�U��r�`H�q6#2�v]�{W�Ӻ�[�����ۀ "���T�<���
�d��.���S�a���'GX�����}�=#�7�a��ۑ]m� u
�yJ�o�����n�(�ב�Ü:���ۣ\G��a{NfX��e���e��H�S���&�L�]�P��wj��������ۘn����;�5��p�;�l�/��,��iIS|�~�u�vh���cB��Qjߺ�n���/vodBL� �ar]��9n#�O�}G�˦ ��]{v���ֽ+�<�ՙF�[�Q�<s�.�t�S��9��R��N��2Vv�VӼ�)-����睵���q��Tޗ�oK��K\��ë,�\�i��}��W�|��l�"�W�9���>nk��ʃ�Cߓ�as���a�:ŽݭYꝲ�\��W����L�Ψ�{�O!+����ڈo)�9K�W��P��68���G{.
YG=u�w�����-�o���r���g�/;�7���'�sl������j8��)(�Qz�hZ��NK�7�H�k����CgZ�]����\Cu<�f�����Q��N6f�\.q=0rtSY}U������zS��Φ��`굅+7cjS��H�|�|*��c{��j�!;j���<U���in7o��e����1	F1h�,�m�3��i����V]���pbZUy���_Z�jyq��.������(��T{���8W4�SZ)8|'�G^J�����=���|ZOB�]����U��l�v��f{l�M	\	W�:;*$���M]�P��np�'�b���+'wh�5�zgX#"-냗��z��P�LV�A�@��J�V%�l����b�V��]�eLz���Z̎��!*󠱧i�!>�|Bx�R�ӌ�ʼ<��⋦>�ڳe�U��{!Ɂ��땃Ǻ��YT�{�ԑ��V�}}c���V73Ӟ�ù^'e-�u�q������}ws�Ș�$��껋����Z!�Z���z��O0t��Yνp�}�]
�F���A��U&�Gu�͌����S�yv�6�s��;�qo!t[�?+�1_r�2��Ժ�3�f�f��98�`ķ�Q�n�����U5CtU�TCw6�f�/�[�5n� }x��w'�Ō�ڼb)�Ŏw���r������5�Uz�8�I-z+�Ӳ��oE��_+�Lo�����X��_rY�r����"aR���оr�x���U��g��~^��We|q:��Uy9��U��ַPkp�W�d�T�C]�]E�����'�l��\t��� �,�q+��f���=R[��f�j��qv�憪Φ�4VC|wC��P����/��-�!���=�y��)K�'Q�״|���9��1��W/2�ݩ�_s�ކ	�mQ��(�a�Ϋ;Z�ߩ��4��(ئX2�a4����r�z��O��S��gv�r�Ϥ��@�B�N�)!d�w>�U��W�h����ϴjҚYR�������{9�]����wt�]����#k��8��^��T��s>3x��ꝵ2qk�=�x�R��k��
r��X|�Ru���to������:�k�i�����M��'%Zd@B�^EQw��,�$~�1|��^������TN�K��w�"&]8<�-��Y[������7|��;jP��$�)pXo%��Ƹ��w�V��jb���ҷ÷od�M�q�U�	P�X�sY�&��[��es�e���s��ү�iK�M�>�7�Q��2�����2��6 Ӯ\�Q�1��ܘ[3��Wpf\��]Ɣ�p�Gsy
Y1s�;�0w&�x���tC�b1?8}���2�	�^���6�Y8\�%X7����fө
l�����n%c<*
�Kj-߲�b�y���ݓ�(�b���X�BQ��E&��U�4D�6{.�/�\��<�-�_9��V2R��(�-�;	W�x�U���$�����,��EЬ��u�YC |�����(�.{��"'����x23oOP�s��ε�KtcD#V�u	|��%0%�7�]�:�M��}�}�s��T���wv�t2�B}T5.��&��P{r�ss�9��*���cۨl>���d�Sx��^�5�7��dt,|6�����+\��=r㈩����kStE��N-������^���QE'��Í/ͬ��v��j7��WC�(�{���pi�0���+h.;Gߏ��.�g�~�#͑��)7XQz�թ�^�gaڎXwo�7a�O�l����k�4��9��(��'��c�+[��޷�j��VR�7cj"T�j�,�ò2�ǡ�SW[��[�?����i�㷵
k�n���e.t^ik��؂Vܤ���x���ܦe~�Q�]�Xy���q�{/v�o�⣮V��ìQ��2g3�ζ��S����2"�,�\�>=�Ҹp�*�d��6i�J���\f�=xE	��	���L�s��1t���K�Lw ��u����U�m ��=�,C6��=N\{h�syz�a\�t��\��),�6U�Q��Ԧ����Ӏ!����^�4ֲ7}oq��8@Ż�P7|��K�v�W��y�F]��sF��wl:Z�U�W]�x��GU]�u�9u;�n�n+���}Hb�;�3Q����YWc��޷�ԇ{d�'�}�]3B��x����Y;�V�����ݙ�ɕ����P�쭗��U_�Z�&q�/ꎔY����s���g��������u᥵li��To��[Z�%�w=��;�ޠ�'U��CWr�`���P_`�}�U܂ap���(�h �[v��3����:�r6���6�!!�琵�V#�j�N��BՉ���^=�Z���B�_66��#�o����kS��KI�އ���b;����/'1{�ꉋ�mc������j->I��Z0��jÕ��Aqh\v�(|
]K���'�t�����yq{��S�p�����g�Ϲ�Z����*�G�E]��.ۭ�c�竅�{��V����p�m7}��U�=I�ʇPfv��f��d|�ۥ,����Es���3 ���Z�̾�0EM��gYUԝm�����n���2��.���v[��<�j���Cf��b��J<��y�.h�:^R�B�����Ģ�<ۅK޷:�ou�Vw69u(!Yމ�<��XU�~�")�/7��ps�U�}k�Dl�����a�c���O;��O��F��r��ꃗSl�����y<��U�o��oku�s��D���e?���p���*��e}�C%
�ޥ�������E�Y�ƻN2Su�ת��{ю!e�°�|v�\:"�]E��1�����uQ��}Jq�r�_Ϲ+�ú��Zr���2�%Qs���s��[�f��ڥY ��'�d��v_wHOSk���.��5(����F9�hƸd�s���Rby�ݻ��2��ݰ��p�!��.�-�VLOkЙ�9T��8�Ĝ��#K�%�Z���F���Ok�rbn����t(��M�N@qt�_��=�����ir��'-������^���xN��Zۓ�Vf�b���׮�%&;/��h��]��K�����*�vr�$���*R� t\x���{V&��QH{�{��+
;�TQa�n�'{`9ۗ�i�69NQ(9.��	��̾�s
W�����st��A��7���*�������э�Y�>U"wق���f�$�>����lp��{>��O.֛����L{�<�������)�,]h��GC�\垊�!X`�!yy�c�yf�{.��"K��攷��F�æ(1�Uu�"��x�����J�;���͜�WsV��\��v��X�MΒ��X2L��TŃ�����%YX�GM��juEv�(�����͢��T:��[�9-�;a�F�3i��7čLm�*�Q���H_Jo��*�W�KՐ�Y3�(�+z���[)��E���e]�\�ú�6��~I�eNoB��1�Q�}I���9ή^�]q���/�"[J��	�����K��d��R���+r����g��>f��ӂ��S�]�v��Јc�K&)l�;����
Bq�^�!}���hk�W�̺=V&La��d���=N�d���*���l�6E�S�'p]�=��L�S�l��#<���譐�yb�=��1�]O��CH�'#Xo)�;L5zE�Tc�ܫj�V���.�ѬZN�렺����n��G�Sjdhf�C��l�2��6fgM:��<�]qH���u��ݵ�&��6X��C&la�8_ev�z���b�=���o��X�<¹R��&��F�}\�z�G�r��3��̹Q̪W˔Π�o�w�h\e�¸���(+�S$���9K6A�u��p��PfbQ�>�/z�q@q�F�{��CL���̭�� X���ū�����s:P7V�J]�������>��W�9R�N�;��!�F��ΖS�u�7yԊ�V���X�ڧ�f��x$��VD��[Ҏ�(�6��k:e�h�\��>S����'؃M��UY{�8����헕5]YV��䃰�5M���6�f�R�,�Yc�=���8�3���w:)�a�ziA��EjeioԔ΍�5�J�S�"�Vb}�5�B�����t�У63Qf�$4���3j�V���Ô�=e�_؍:�G��*��6�}�B�s���w�8N�AJ�{.u<خ�K)���vԗi�=�1܎G�͂0�4�g^hŜ��T�V��7�E��W+�����A��Τ�u������Ie[��+����>di��bm^=�iK���ck&!�H�!s/3���hS7�yB��i6���K���HpG��]f<i�,�ޕ%�&�&�����
�k2F�y�*�����A�/�����{��lW��X��6��3j��-���V�$��d����r<q�wn���f���0�����
�yu ����`A�w)�W�����--�E�LKE<�NL©	k,�z�3&fjf*��*�dՆ�(�Mv�9�o�uLi���!}}O335�Y��;Ğ��Y1P]wV>��Ε$X�ܭ��B�Shv��������~��n�sc[��.P��E��M4!�:t��ݹ�*9gu�M�ܹr܄�E\�%\���u�F�\ە�E\�ڂ��Tnk��B�.��s��u�F5w]tۗKE����b�W6Ms��.���ws�s�ۃ�\��\��+���r�u�I���\ܸnn�m�u�1W9c������рJɹWLXƅݨ��Y�r�p�ɣA&()�[�9�� �
Fn:E]8���[����w�N�~�s��G������R���1T&,̨��;|Niʐ��ޔl����c���ﾇ�uw.���&y��o������N�G9��M[̕�)d)t�-]�ᵜ���_dN���.+�q�T��,9Q����d�)���o�p�vu,�(�,[I�k]S�jx�w>��:��esú�0��Ye3�Yܘ��)u7����c�U�\���lTE�,��W�_5%��g�;\��!�9\^p��T7"Z��SF�E�ި:�57�9��F�8��Ȅ���w�]�P���+�}}ג�ΡZ��������M�.��],uK�)-�xq�����&�oc��m��1�U�*T��|��=�X���^��=�=t窽�L{ȧvᷴ�������Uc��]NL�x�VENF<�Hڠ���/J���K!���~�|��L��Y�(������"TWE�����u�����_t����^������졔��O��z)l��L��f;��hyv�G`�p�b�.}]�r�:�j�mѮ�gyJ�_���]��ໞ��l!E��<x��X4(w���M�օ%��r��C��01�6v��Zz�S�����`Y�ڙ|���Xݙ������9��=�þ�a�U1�1��@]����P����hI��wP.���3�tLr�UT�0�-�0�N�=�,'�q\�6;o�����z�kTT�g7�W�7r����M-���;fo��X+�r��5MNtM�'��d��s���5�O Wʀ0�=P`��w�4�f��8F#w�Ou΄K����t�̅�&�Z/a!�C�ݪ�)���}+��V�3=
�oloh5�7���t_ͣ�L����!�价 F�py���HI�y_�h������`�N�-��y��S�5��NE���d���µ�L�%���B�qM�>ĺ��Q�gz�~��k�E�;~����Vw�ql�)������{_O9��_Y�Q�t�3ᇛ]������1��ѹ{G��_qOj�����1	/v��
���"��������h8*�.�\�넥X.�$����d]^]l��@�y������x�x7}�r6c)���]�y�lT�Qs�hȵ<���q���5��t���A�,7��3f�Z��6���TY��n��l�/�*�� l糹�S��aM_�y^�I�X�cJ�j�rp��aT=�I���h����([N+�w�Σej�Ҟ^>ݸ��Қ�|l-�Nff��	��@�ɨ�e�NA�ث�v���|����v��I��r�ɫ�JgsY��GOU����b��Vڽ�����8���Q�Xl���T��R�3�Rx�z2UӨoWa*���zf =���1:b���f���L���U�s�M���yG"ʚ���_�/�����%aZ
�re�;�ڽPȫ�ڙ}N�Шn㛡���+���بnw�����F���@����ݿ�f���;�5�
Y�:�lKâE�Q���>�=/�nw�les��m㝋�]iQ�w����*q�ɘ��4d:��=����:�����x�̯db�f;J��9v�R"s'�4TV�Ie	mf�]X�N��|%[ͨ��
>����^������
hF
��ƺ��Ԓ��2u���,4fV��F�>OiPv����龹����[��<���I�����pd�ѕ�wCU���FT�G^:���(jvZV��5���f��p���6�Q~�Qy8꯿}Ra�@k{�-�{�������9�C���u!غ٘N��k��X�ϩ�TE�Ǎ[��wR��s(%�1\5�1�JU�/�k���_b�<��\S?d){�]L�J��Wc�z�y.������㷛��_���k���ڵ�F��q�w����Ղ��QKt���uo�}��.57����{�z���g��4 ���+�c�Ī��	���N>�;�㶋�J~�����Jdeqp����8���,�w������VJ�Oj�UCO��F�*rM�FU8|72�-���wl%�.���Q%��d[��[�׮gw)�@֨z:����	w7�8�yʗL/�h��҉܌��pn�§gwى�^�^�}
o#cf{���9|i8�wF~������Bi1WY�W�i�r����3<�76�c��zi�Ը�+͆�bzD�w�z5[�
[)�C���)nP0�0�[�V��{E��/=V)�+)Zܸ��-�4�i��5¢��Cy���9@Jx�v���&2�Ӱ��[y.�Gn��I��2�ǵ����.�WLĦ��7w�e��仪#T�l[	7
b�9B�殄�d�s���|a9��?D�ʌO2�
�>�a���;�Sܽ�r{xq�4��B�4k>㽒�k2,���Uo��+����Y�oN��v䍄���;]�󄰽@?sg���5�u�m��1`=�q��83k]�r�U{�녦�8-�Vd9:2�U;e3I{����i^�Co�><�t��q]M�9QQ�2atGOsl�����s���}��ݞ�j����X��v�7LGe����Ϧ��|�T���;U}\����b��r�)��o�l�E���iltCŹm��5�g��Btt{���{k�Wr�o�(�|�����^w;ީ�л�WE��bT�m��I��v�����Q�U�mJ�ZՅ�G8���aC}K�0c��B�r�Øm�|�S���N���;Ɂ�K�+�[��]�(�y7�Ц�=�rl�
����qX|*�a#vE����ì��+��j�5�;���ͼ�3�ґZt)p����i
�l}qk�dπ�w|�Y����*��������Ҥg+T=1�K���	����>�ʘ�5�WЯ^u�UgP��+Ѫ�<3�3���J�,͝Qw�\Y=�ɕϟa<�p�o��ҚZ$u�
Wã�aù��F�襄�6�R�	�^
���_ы�[��ҿ���g8���u�Gf:W0'��חkq����Bʈ��o��;��R����}Ԟ��%*�7�\>�ѓ�5�[���3�Q�:`GT��3�����Ի���}'J���yUF�7�	n�zFz7��/��1�t.���{Bwz����B�3'�w���A!�x�.����f�����~WNx٦��[v��#�"���˧Ж?��|w)�9P��mC�*��t�g�>�4���Js�Q���H�ʴ_�l�ku�J����m��G"W��[��*��Nm��gΰd�Q�NNK�y�
w��m7̅�����Z�.U�¤��u��	'ݾ!j�)D�����yl�#h@h���۲��C\�6�Py���Dtq��e	���U����[`���r�5]9�����^61�����K/V證� dd��I����sZt��$qO����]G�������}a)iI�໬�'l�z����-�/��qJ��7�������}�EN�R`�~F.\��ޤ�ͯK9=ih�-�
;s?Z�u�j��f�!��^f�z�>v\�K���мߗ �j�S�죋��^�(湇5k�\3��2μ������GϽfN3�]W�N�$�W%Ͷ<">� �Ǘ^��l�ge��V{��ʪ�M��n;z���c9dO.��d����Ƞ��}�*�d�8�_OԹ���[+U�����b�m�+��5��|�3UXº�S�S��#�l������j�t���-+�����m���!��-s��g�nJ7%:� >���ޞ�4�eq�bģ�hUjL��B�ng��>e'�sY�n�Y��S5*��j�v��!-�MJ�mu����:����c��:���G_��b��Y�V�B��1�b�PZ0���@��;�f��[bPP}kp�^��e�snF�y���&la��[��*̹�R������b����;BLo��^jT���R�8&j�L�B�yE+t@7�1�c8B�	!H�)g����D;y� ��*�C�	���b��Z�ʚ�ٖWd��]�������V�Gͬ��V|�<(��7U{���Ͷ�9̀�-$rT��Ƴ4Q�aRN�����W�E_LY;���H%踏M�P����/�����X�c�mD_+�;�}�[�� �	Ş��\o9�=�M��{��Ɵm�J����T}�O�l�q�;^���]cٜ�8���F��G�	e�k?Ί^(K�X4�H�I�f��\&�u�'�ro\D�X�l8׊f�Õ��]y��u�D����;���3��N��^t����e���1���35rj������=��_�K[�u�i�NT�qR�}kj�b����[�[Ǻ�����ѣ�k����R�����Wo7AT8����c��
��NWڛیi����l�N�RT�.���t�\�����BUA�_J��X��'�A�J�by⪗����Q�X�s��"�ӥ�Lgf힫z�`A=Ѿ��W�+1��㈮|iN��S<1eb�W����� �ف�#����h���W�M�2m)��Rﳫ�z.�s_ceѵ���T��[ȫ��bՂ�.��y�p��z�3j.���|�>��N�]�ם�T[Y�+��rm��#Y�����8���7�s����e�8������I�~Zo�*-���t��Qb��[Z�f'���"�cmK��_4ҷûod�t�eta�� t,r���sq��q���˜�p/6��w�b��:�J�	��T����̛_'~�e��]��ec�xTz���W��'0�t�B�n���B��QS�׳&k����0�#�enb��[�p̰�c��ɪ���}��s\�H��bq՝q-���=���B�s���c����UU��'է�H�����������B�s�Tڇ�VC���'�l�ٿ]Qy���f��97��-sp�k��;ݺڢ��o�5��VS�V2#h+o"s����������<[Z���u7s���d�WSZ��F�k��%��A����sX�ުp��ʱ�]E;A�=�3[<�S�춑����ߜs���\7#�;�옮o�%Q����Â�כ:�3G8�K�կ8\J���ʁ�֭ �OC�.�	��*s]�����a��]�j���eF�X��@u�t9W�S�Ÿ{��RxA��z���k�:���V-��`��QC�~��y�M�l��M�ƅ�	���;P���P�o�q!M�Ⱥ���z���^�.or�3��9��nV��־�8^lj��t	�'�Q��D/jꝯ=�Բ+DI���V�@Mh������>�ie5�:�0$:��J��T}gND��q�����O�)�ao-6�r��k�q�}Q�J�[ƾ��+-�}�˛7;/*�{��ga���\v�Z�tiO.1�ݸm����ja���6�~���ܻ��3��+{�k�_Q�Ȯ����"ҿ��ݼq�	�s}w�$vp� ��u=�xE	���6:ܹ��
�\��L%�U�_uD&5���D�7�&9�����ΙX!)�����]�e�bs�+�tt����d��}(�w*m�Y��'��TT�t.�1�k���!�ۈ�f,ԱAa{������}8��h��^�����Nd6�������t��f�)m:N����c[�3�b��8$%��x�ҭf~���@*.A�Y�o�����mdwmt��i'r$F0�]�j�p���)Ҕ�ǂ�M��;D��׫y�j��׮+.���^d�ɝ�~]͕����Tơ��Y{���xAŪ��������v�
��M��1��$F��X��q����m=l��ݷ9���u��Ňu��\� ��<����ӧ�6y�Le:�.��/f#���ƒ�L�.��@_#����۵:׽SB�"M]z�t���vƺ��{{����ԳZ]s}��Vl�
l��A��`
�[;�6�E|���t�}1��ݽ<���i
�Xɣ8��W���'�o�U��p�1��by',ܜ0f���dծ(R�AVa#���fQ��/	�q�w,��¯Oax�  ���_fT|��n��;tqz[Յ<lm��λ��{�Mqu�Ļ�n�i�{��H��}���� qڧ��G<iھ��I�v�x��.0V��������U�
��vjs�Q��̼>w�=���[�\�PǏ�����2��M��&I�^��X������d����;��j�\Μd�Ǝuj�Gib�%�,��q����	���׼�rǭ�Sn\�]zd��sv�l����Bb�괥���E�I\Qb{�-�O9U�%�8:��V�=7�t��(��� cj�ʤ�Y	�p��{dt�#�gbf�����0J�V�����%�ڃ�6����)�.6P�!��[�zĞ����$y\�E���錹����>�_�{�2vѧV��/�|���f���h6�+�WYZF��|��g�C����E̩7�Е�ە1C���}�I�!w�S���P1m'��Wep�d�P����#z����q�w%����2���kHj�|r�.{$e�u����ɈމW�ۖ�l����j��]��Z;a^+�d%O�gz�GK^ް�-����AYl��Z��p������eV���PeZM�N���G�R,��r��	��M��B��g�����oY׊C�*+xD�����5+�r�V�	��Zq2�3�H�N٤�3�on��l�}�jٗ���;/R��UEM��ee�H)E7���wC�k��a��_@s{4^�!uiֆwL��A�>���(P�f�6TMp�����"�]]AܖJX�.-�%7y���괎�����7����:�}�=�?��]�(�÷��[ړ�J++���L�\b��S�������)���8���כ}YfR�=\.9ͽh_;:WwDŸ��K��C���4�6���@9�H�[ʆ��L�M���2裛�m�X��ﺻ0�Y��oF�p�9�ˑ��qʷ�k*��ӛ�|;Yl:�9c��Y,���&�'�ގq�������+���vԵ���Hpe��Yni5�����E �A �5DP��"��-CS��+�k��]ݛ���S��\\�9� �:Yp족i2�$@;�63'q�JS��%9��2��;��7wG8w]�Q	���wwS��d�ۮ넖.[��wvИ�� $� ��Ȼ�
�+�����,\�v�:�]�K�tNrqur�s����.��e��W+�Hw%��:���\B��s�EM$��Gw+����Rn���ƔB�w)3�9w]n��L� ��9��!Ε��!��wsdw�P�;vH��;�9�8�a1B��'���"���P[��]�f8)�8[�k-g-Y����y�gkV���'�]s]J���XDu�����5��ulg�L��C
��Gv5G:V��h���V� ��-��*��y���2��^��2�����J�RN����UC�'�<�x����^ �U�ݺ닾*ZO��ukL�c�4��R_29'��%�#�E��Y���Ёs5�bL��5����_^=�����Wn�T���Բ��/�r������jSE��0Aڒ���O�o�V-]�4ꉎ�m�6�B�7��'Ւ����阏_��s+ϔ�g�ѕC�h\t���]Kۑ8,ݶz���W���N���פν���ކb���?��(��N��0Q�M&�{��I�ғ��Zא��%���b�ۇ�:���ݍ�,bqk�����%�<�_YΨ��iS��7���Ȧ����x;��ֶ���cG���MQ���N�}K)guý��F�ա;�iwc���5�t˝��(���Fѓ�`�����:�{�J�bj����ME�Hp6e-|^W@�&��N9|��X����9��s�����)��U���x�p8wx�4=��]{{��7fߎ����9:��遷$��g&M7���N�ʒ����n�=���R���wg�W=���u
��1��u�ꄟ;�����b_Ly]��`]O�%xEv8��y�ߠ`�*-�*�G{��#�.�.6�u�WZ��N�t�kR�|;���2]�L[+��	P��@~��e��5{J8��8�{�`���5ʢ������б���]_+D-��	U73sr|��h�`�pݼ���2Ի���� ;C���[��q�d��'���Y��2���"/{�u���b'�'�Юcw�v��j�B�
r����(.���b붪r70�#7�x��[�1r�l����ki��@|NT�u{Xjݞq ��*s��3�YG�7�h��W�R�c#�����s2v���΋�vw������K�^N_޾x�8�Q��/'_�p�pq=)fI��l��pӤ���4:~{u5���r�+�b�-�L<�bB���F�{�c�/�H��wsL�����4�s>̻n
�Qšє}�Éj�1��۬2�ц���)�]���z�^��[����͙�O�Y��f��8���"����zxE�_V��p1�����Ù<�g7Ok�ME˓=si;�м��O�!*�|�z�e}7�߲JQ��:�k�劓���+f�I���)��]�ު�z�ḡ�f���dn*qc9w1s���j�b�]/o��Ży��j�u:��΍�R��M��$軞��y����a��B��T�y8��j�op�㍭��ˀ:^��X�u[�Ou-���Ң�Z�<����p�sU���W���o�m���~�=�͈��_B�y�T%E�ՎQ�\���92����65C<�׼���#w�n!�����酵�Ъ6:�Ku[�ED�CV@���$Z��>������6���۷�2b��2�%�5��jʘa]tWS��h���:�]4��)}���F�O��K�.v�@���]T��ɫ;��f9�t��Xf\�S��9�L�N�F*d����Æ�zvoQ�dg�2�*9v�Nb��nd'w�}�>���Ղ�o��׽��N@��s��Z��"4��N�O����4�;���r�w�; �wyi?v�A�9�!��S�l��*t6.��⶟;v�{p��gi.@d>	���K1�h�Fj�}�3�}�S���o	����������
�s��+��-�a�Ev�X����"8��&Y��c���V\6�Tީ6�ʯ��}ed:�h�l���Czm�&�����׆+i>��/���jq�:�!T6��CYN�F�|VDh%0�eR�f�����ܔߊ�ڧ��j�ϤG���^���Wb��V�:u;���lL
�m�뵯�'*1=5�'��ROW��u����Nٝ����c��S�-�A���[Aqӊi��]K�=I�=�9���cs^���ͤ�k��eD=���,;��m}<� ��!{iuN.�f�=Գ��cs���Jp� �Έ�{�ݭ��:���!T4�حi�dO[�].T�ޭ%.!재��)e��&�b�l�����D[�iq*�i�`偡�f򯖸0����k�w��j�ѥ<�p�n{P��p��Hor��|\]�͎}�}1���&P�("��*��n*�t�B>�8h�X��j��*8��(��:�n���b燦d۹�2�s����vL�S��jL4zi��D�5;�E��(��8q��Fd�Nw��ޞ}���S%���P��](�=өk{�g����ï�ˌ]*��pSJ����9C�ۣ�T�hOOK��N�%02T���
�\��L+/�	}{'v+C��yԀ{oFLR�i�e\a��B��t��>���/�V�ʝ����n���[U��;�[��S�Ìg��A�s��ivz����2�R�ȸǛ�@�c��-�wz���&o��9��s���4�\T�J���j�W��9���V�;��;����'N��d9�3@<��F5'��y��C��0�oB67���y��֙ǎW<�J��BO�낗��<ڤ�å�^]����=0F}�Q���Ux��V�5���+�̅���ν�Y���ߏ��__$�Cp��Z��v�X��y����{ʻ�R^+���Ԝ>������2����T�[Z=�ą�!T�[�+�z�˛՛�Jx}h>�^J���\-o�͏SHRc/�}jen�z�:��>Ru
o3�b��oo*�N%g\;�=:�Z?\�ʞ�J�^�#�x2�.ʡj\ C�.4/�q������#��]�4��Xr&�H��n�º���ۢ��%�J����Z��uu��b�xN��<�k��k�Lߗ ���l�q��s�����4���)6����ꜯ����y�����V��L\�܋�������QK�8�ɷJ�:V��k��>of!OvZ����ۏ��t�jq�%Q��R�ε_Y��핪������aX��qV)�mk����fw�#am�q*�=�*JLW��Y\��b0����E��U��5��\mN�>��a\��7L��[j��r�7M{�Ә�=cU�[�u�����M*�z7z��O��*e�ц����zm��9@4���B5!���"����׏�_t��u��{�\c�T�ʲ�����Ƭ)#��-�zщN	���ˀ��I&ʙ�z�TCy
���܀4kҮ���T�QB�7��ޝ=�)+rj#ݰ�y��˅дQ}�V�@���2�fhs?l��k�#�u�XpR�b�^�.�A�P�v���u=�1��R�[��{�*\h��J^���W��]rq�CҬ\]��ȂϛN��z�(�Ζ��*�
,7�uq�H\,�ٷ}��s3�0t0���/���h��4]�ٵ�w"�����G�*����m�s*��b���9�Ӹ�l��C�����t&�e����s��ٮ0��dL4��/�K��_^38��#uɣ�S$��5ѻ�'RS]w֜�_cP6������u��YG��G��8d�\���Vlc��|8#��x��SwܫZ
�����z.u�̯�X.1�U�d���;O�q�n�/'*1F:��ԡ*�|ʝ�\���)�~�����{�jJR�⧎[9x˪6���F(ĺe��sb���mBQ��2���<��������;cj'���*���r¦�josZ뛪�#9j��Qp�_�'e'
�k��k���J�\4���Z��<���͓�͎������wՊ(���Ɩ���g����ۋ��&����:�9B�I]FE�'jV�]�,Y���m�-e��۷��SM�V�<:;,%4bc�(o��ֈ1�Ʒ�I<޻R��)�[�e�+�����s�m���Ѷ��W�uİQ�Ӽ��m��=�T��ӵ���;����%�d��ۈN�OVv��N��]vE�cc�*m]h��ý ]��t�];>��A�Q2�Q��F�J띗k�PE��d�+�W�Qͥo�]��i��Ti}��xS4��w��,Q�}}Rmc����M��+���5��p��W�8��u���"�V�w�3-pu�K*%1]2����2�ҝB�څ:���Tj�ۖ��wc;�'R:F8�]
�]�"�Oܷ�'5��sH�}�_7���k_�p;��q���^Ҷm2�lCw����b-��a4*�@�eu��E�Oc�=����LL�j���t�1�츂�h�ꁁGI6-F�Y�pLb�n�z<v���xGo�)b9�U�;Me;F��̋�{4��ePÃ"m9�k�e�U�:�ǵ�A������!G|���׷�r�ȄnE~��84��9�ȴ/���V-]�4���z��ϥ���f�����?WJ2W�Wz�B�~�ڜ�f��и�Sh�j�>��^L���S��ј���a�&`T�N���JM)�f�l�2����S��T]����単�`��+v<䝥iYg'Z��N����ͱ.�ތB�w{tƠ���N���U��Nz����!�TA�C�®���PV.NY��I5й�_s�ٷ��M��y8j�`��v���7(�1����~�߬<���~�'�˅f`���r�6���9^�|ݭ��:�!�{��gT�p]f�6��b�÷�R�]6;�Y�Q���Zˈm��oM�:����ct\\�C/R�R�jJq?R�#'�A�\n �x�u�kx�>l9v6E���P��٫Ʈ�
O���::��pe.|�b�o]�-+�p�b��P[�R��͂���1��t����R�W!�o�Y��N.^:уiy$\��mn�ʫ��y*q��Ց,�K�k�+��uǠ5}�M�D�=�Mj�G��X���u;�4sqk�݈���R�-�S�,����y�4-�7͝��_Öd:��|�:WW�S7�*|<2
Z*DYV���j:x
���3�&�ݸ�+)*9P��a�}e\:���x黺c�k{�z�I����,�>� W��Ac���~-�Ǻ�hO���;�<Յ����\��k�eӥ�b���;�f��Um���^��]���J� ��#;}�l"%��
�wcB��"���{�^���X3�y��a�����gmV��V��ٝ�Y~�b����p���H�B~���o=)v��3�\�����݃�z�Oz�a��Q��gnT�<f�(���1c���w�_��V�1X�G+�����`J�:��ճ6*B�6��v��������8�ݭ�������+e9ّ�rݼ��(Y}9^�Ny���^�꿞�p3*YG��9�\
��n�cS�0�ȼ�)�~����w��E3irg�l��R�����QZ�;�6:bNs��PN�<���5NV�B��[���]�vs_:ak�ڔ�.V�����A9}}.����_Ѳ�n57����q��1Q�1��VѾy.y�].5�ꅱ*���1�����j=|�U1�Iuaq�ʥ�/�Hr(��C�+{��5n��Y/�e���w����Uks/��§�(.m�Z�����WCݼkk�����v�6��"~����f��:�g�W	��>;��W��D"�;�&|��v� �w{�e��>�Z_+z�Ks�C�Y6[A�6�1��\*��g���0�/�����&!QR�b�=�`0p�J�hw�Z�oscަ���T��Z��'5;���sp��C��Y{hҊs����鮕�hK�CI��ޡS��pW�6[��y��Ζ�Oul�̻�}$�tL+�Vr\5�vM�t�"W��7q#�����w��;�{�c�l���Y!X�"8�� ���w�EX.P�z�=� �����5����]��8���v����1�]*�b�Ò�l�$S�&�LF�R�u�/ZMe��蜚�ܖ�{L�H��K)�%������X�D����)�h��vk�sZ���V��3�7,����nn(�[I-�R�i��RU��e�#��63���o�e��O8^���Z5�gj�>t[��W�+�J�Ԓ���Es7(˃6b���zq�o�RԽ%�ߵX���׍�&NG�:Ⱥ�b���Ë@kWk�M�kK�Cn����,�bn��.#�9S�oY��9�5��D�Т;v:������؅�h�ox pv� ��u�Q^d�9��5vot%[������QA�����ߧ�&U�%պ�\������B���V��Y���2jZ�e9�U�+Im�Êu�8(I����)����}={�t�lV�_lM߻A��7)����f�[n�E�N��9
�;�;���E��1)�ϫe�\�m>1�%M�t�'sÎ�����ء�w�,3A����@4[����*#V�t�J�˼�T�A���v��:ѝ�d�O'M��]��{x��)��e�[Ὢ��k_���V:���Z�7���aN�3ǼvW!�l���P�#��Z��*��컲,�������l�3U�k"����3����:��OG:�����?�8��D�h���Hⶲ��� ��h�{jX�(��1�{*�pyY���i�&�S�CǹVn�5G�����p��8����-u�}3{q�E#���4˄m��8�˱�kz�]!��Fq�����9z�ݩ�4l�/�Z�ѫ����2���lK�y�j�B����/��e�7��Bܗ���Ҷ1��Dq�A^W':��v�]5�}��)�5xjh�Ӷ��+T��쑳۔�l��T�$�f����LzN���&�.ok1�N�/+�Kq�{2��9.,-9��c�R�S��D+]V>m��r���i`��+�0aǒ���as�r�3�@��xq�צ!S�ԆL������nC���;{�k��f')�|�!P��s��ψɕ�Ƅ�]j�3���֖h���{wyXop��۟v���s�9��ȹ���-W3Ս���y����l��r7�\��
��N�@��t�\����V��}W�f}���>�ky(똺F���\�v �ua�\Q���ڰ9��;*�^�}��C�+�۴Qr�9�7s���rܝw���u���Wd�.�"��XD]�q!�n��]��l��su����I&����,Y�RT$���9�)K���D��21"�0gw����s�� �\��ʺhh�.u�	3H	3��L��9����LJcBF]u��$)�
5�]4̹�a������d4��7:�s�Ӓ�JK&ws��wC(h2���C�M�\�2JI�� ��R�s��]�A��Iwr	]�c	�v�1I1)!�sp�b����]�!
K���@�8�K& �R��2D�q`dcr����z�����~ߞ��7|�'w���)J�j��6��0��mm�J)��*�\5Ӛ/8�E�L�'j�k����'���v$,�ы��]W	��jV�ۺJ��W�tԤF��S��k����FW1����L+�S����ŧtTB�S�RGq�$lt4kq��ϯ�%����Z�ڲ�.̸	�%��:Z��sn�쇧�"����Z،�ab�/���٦ҷ&�ݸ
���}/^T��TO,��1F+����y
��C�^sE\ʭ����Iα=��ԭ�7v)�f�7�ѽ�O
o�U|��k	�H1y���D��o�.Ҽ�2grOwnsD�vl�і�w�C�j�yN�7_~�%�Zʃ��Y�e��Hו�4dVc����X�#�����.��.��eF��`���H�{_s����~>}��~^���mT{տqr���{���T<�<3���o��tMLG��X�$r�P�C�q�8����=�k���$�p�'`�4Vk&=�~9f��,�֨����]3Q�k,�6(wy`��ë����ѐѢhж=��۟k�k
�3�1n
本k��Au�գ����'f�)4\�\�C����Fh�뱟���eg:�'Otgx�[C��}�h^LN���bZ�[j���9Bf�ī'	�'~�-��W4�w�md�Q��D/mT���j�*A�ɇZ�O��w�o��'�^��r��;���o}�J�rT֪"�'q��&��9��HW'Ӕ�5��m��oj�dꅽĪ��vT��3�l�G3��B��n�ɞ����-����KY���`���+��Pzj��{e�h�I��t'���rq!__%��.�of��ҷ÷obr�iloa\��yݮȫ<�N�Cʞ���s�����P�sf�.T��څ=�Ж\'{]���>U��鐵݅ٗ�NR�=��Տ��h��:�ʛq�i�*yfUʘ���Pa9��[�p�s��db#1{ŧU|�d�tev�W=�T�>L�O!\;�U3 ��im[�p�P�.6gkczk�B҉7��VWܨe$�Rj\���'�l�\���m��c��R��Hp�HĖ<|���M���D����S(7�mn�����l/vVV�l���C�x'D�#*g0�q
�f7���O�s��v��N��n&r�r�v���3Q���N�do|���sÔ#���<���m�����-iŀ�&�9Pu��+�7�>J]"�Gܫ-NU���.�bBC�9��1U��נ�V(��o�
;e�U��O{a�9]�;(��Qh-�����.'ϥ��y����+��O7N��0�j�/�:�s=����u7�5��sσdx��.:qM����^���t樻�]��U����B���o7�����6� ��ܞ!t�;�����F{��]!�=���R���ô�w��i���n������f���'6�\�T(o-U�����}=]q���m�܊oj!M�[xl����7w�7���ħ���42٤�tS�zw�����s;�5͟{ψ}sPF����fs_f��Zw��R�R�\լ]?+z�i3�P��q��\)f��=�����Ʉ���(����.f\*�<�]�9ȫ���!S��Y����+]�\u�})˻����F'hI�v��w3��W��	�SM���ն}��0�vE�$:�#�`�1�P�d��L��D�Q�M&h1��x���9����/(Q5Lu:��V�r��Ǯ���$	]8C}�OJ���q��}\s�{�b���)=�ߢ�#Pܲ�%�]3�O�V,:�2�X�E�	5��ޗ}�P�[�����ƪ�݉�r�+�v��N`�����t����%��X�̰�c��s�ش������W.xMQ�wn.1��|��Nv�E�=�6�e�X�u�N]�����B��L��fa:x��iԍ��+�+�����툷�9؅�i*.�9�]��N�����lJ1)w�vO^5�흡ѳ�TR����f�90)�Ǜk0�+{<�#��RTf�SyN�7Q�]A}�S��^NFù�eMn��|��.5lO�);nup�[��X�UO[W�P\Y�D���:���p��γw�|��Q�ܘ]��\6��ȶ� �y��-</={^��<9��J(b����mY�_b�U�*7��Uy�7}�j0����%�A�����=�������{[�G17"����M��.T�8z��ؠ?�qw�����?5�;K��/*qޞ�sC[.��C�-��}�.��}��vՑ�u2�l�^C���Y�)L��<��V�u">�֜ڒ��0�8��yf��v6���YgnK������{���3Ֆu�pɖ���O��|�vO*�y�,����;�,��yϊY�@t��7�$�:��B���k����Mr�6��Ī��vWҠ�JL_$(��:B�t��
5�<��o��<ҿ�.ʋMu�t���%�-���Q'f�[vUF�w�Wz�"ԇ��/J�٤�W�r��?;���W}�tO:�Yљ�Ċ7�`�QQҜ��@��:�O����W5��pᩆn�p�WuqP8��k���+m�ÿR�c�����]�a9����z���u��%D�����cas�Qn3 ^���F����.~
��c9X}����a���^7s�I��1�:����ug�}�`6=8 j<�	w�M��=���c���!U��N���n6a�]��"�g���p�}(��Tk�����@y�p{��4E}�>%�>OD��,���lgC������m&���sɮ|%ӣ�	�ʂw�h�n��N���)R؂���{;�A��^���pL���Tw 61>�;�2�Pv�ة�kwV7k�v�����~y,�;����Pn��,��ϥ-qa�;-�����&�������K�93�:4�վ�=�C�����QS��Q�q��fG���N~8�ӑ'��*1��_D�?�����'���c|�t��'Ei��Koi��%~��ϗ�^ v�#Y�s��<r~zD��wӾ;v���}'<v�j\FS���l֛� o���������СGtg�[����1C��Mh���q#�qtET<5�����u�1����d�Z�Z~�����psw`��5�+���y�!��<�R���ɜzn��U��M�@�O��~5�ח���Wu�8%O���Zq�����y���Z)��vf����7޸mC^H��c�o�\��ݝ��q��jtz:��GS�#K�i���{��d��ëW�}�l��}DS7*@[y�Y�ɉ�V�W��{e��EJ�,���A��z��|���૸��n���T�yE���Wk��oL�cK�ǭAR��T�_L���x�K��y޴�y��=ǳ���U�U��w2��t�F��(t�2Ͼ�B�צCsd��*La^��	h�6a�n�2/�^������+�6+̞�W��2�8zPT���7�{I^�.�Ne��
m�Ł>;}�,1$r�%���z糔����wi�����$2�����7x^K����Ł������zE-�/��'�ժy����nn�]q��h!��ݺ]K�3J�/���%N�߶��U������O�CP��d�Z�_W���݃ƣ�cz�S�ݛ*Ҿ�ޕ=���z��3���{נG�.CɗD"�iS�Z�2)�iӽ�oY>Or�����5�����S7g��ND���t���s�0�뉺c��=�L��������W�GYͳ#�F��=�#>&��vDs�vLdG����c�T�6�>���_��Uxj<�#a�/�u	^V�w�K&�΃5��c��'VO���q{΄�ߞՏ^P�+�g�3���Rs9�6;��Fp�${�l�G�q��a�m{���p3�����1'v|A���?z��ϴ}�����z��^�۱CEPpF�� izmqOu�~��/z��E!��n�����(���oW"�����(vϿ1���́���i��=h�w
�'��&�rv/'�{���b�HO��������xq�~��.Z�܏>�G"������R��+˝�^@����f���=��	��z�ns��l��t���}�u�[e�1��l�|�������ty䧥�=O�\����X��)o+�$�~;B2�u�Od�<33��v�iF��{C���{y���Y.�k�K����o+��W�ʖm���7�5n'��vX��I:u��D����o��Ka�!�Y�%l5�mX��]eg�/tNaw�?7�MϼX����'��UC�i�l��/W�툹��G�x�^t	H� M�i�oמ2a��p��q&�S2�ȩ�@��ҙy�P�g��c:_�Fo�_)np�pND�̗�az9��m]��C���W��Ġ��8�7H���چ�<�\y_!�d��Ǐ�zx�6g�z}��؎������wҫ,���BsQ���zhWź@�KGە�h��{cw���WG�]�9�$W��QL�o�tT_�܁{��^�g�0XĦEG���"fxs���<�}��>ts��i��3�Lo:���G�w�G���>����˒}
ⓡn}F�HGklN�z�x��S�ΰ���x��>��s�X�Kև�2��9+�%��ޏ{.Ȯ
��j/��
�;����缨�H�w�7QLLSU�o�s�܄��ۼ��"��G��zjE>�s������o�^�1~@o�e�SL����:ja��n�Y��8Sj�8_�ٯ16t����\f:��B��N�G�������nl�����.e�3ax�n�;ͯq�/�����N��ą�������AfI�醥==�W�]f��B�
�����-�R�9F�.��쌎����~,����/V�Veb�ٸ%2�����a�÷�:�w�}�,Y��j�s+��P1<B��nE�b��:��<F�DrE�[�=Q'.��u���yApP�}���he?]�F}�����{�X/��IG."gð�X�._��Vwd���ꂿT��eoW��q�>e�9��,�q�{�\�'̞+}�q7����|zt2.�<�����W��N[Ǩ���C��L�>�c\�������N��m��^��������<bݑ���
MW����>�>�;�}3�vg�FL��s�9�Q�M�/�ǵ�h��g��d�gΧ'k���Ĥ�����?vc}�}���U�j1]1q�:��L�'�]ގ~�qsM�}����l�4w|�Nz��{+�\G��1�~�� �H�*M���j]�xe2�6��oa��/C��+���	��D�y�ӑ��}��c��*�~�(���P��(�tX�x_��{&.LIB�B���L{��l��7��q�G���t�{�F�_�}~��N�eƒ(�l���z�O�H�g@��;�pproI����w6XT�!y	�������|��=v�x�9>q�sހ�<��Y�x��7�c�Ͼ0X[u]F��x�9\����[V��:��C>���s� c��eQ�+�x+o��N�^g,.��a�w���<�7\N�|���1Os\na�� �:ո������]m��O�|��.��V^�Զ����ZH�%%ww�E�4�9��pN�Xrn�yh#2�Mwv���:�qd�B�f'[%sԆ���8p�:}7 ى�H�ɒ8w^Β����QC}����X��ۉ����O��s�Z;��<ܤ|�U�n�sΕ��n�<�i��^�{���w>�@�D�g�&@|j/�b�N����{���W���ֲ��l�W]yG+({��r��k 
��)�Q7>o�6�͢�vN�K_���,W{L�-zd�>��4|��b���ް)�ty|=���>%��H���/u����8�68 .6�';��ע��	��34�|=p�fG����/��<o�{n��Q�q���2���7�[���
��{n�$�(�i~�}Hu���]�����F��3_^����ǃ���O3^�m�Z�P�މxuϪM�������$$sbv��e{��5��\���ζ}���.�\K�݂��Fs�����]h��V��p���$z�)�vVV�;�WY�r��j�xtv#��n���g��/�d���{���|�t��s�hn�tL���QC����;�N��4<���'�Z�1����[w��~������\w��w³�*��DS��T�_}�޶,;�ǯeX�o��_�s�o����0V:g�1��U���lN/����s27��:��4,��n*���"jgX}C�\ťլq�`
"=�9��bij���Մ�wn�S��%�RC�� �8u��[�]�|�-g��l�_ Gm.ܽ��f0��*Go{�����E}'m,��L	u���\�!��2��V�X���Y��;X�TQ��
G�L҃i� {qo}�qc���}lK2g`�����q�T��S��ԍ�7�����s�wK
N<�WF9��b��wv�2'�v���W�;�sU�c*���1]�B�]L��-��W]i`��ܺB�]�[�D����}���R�#}a����8=���7�{�U�,�D1�>����xc��kCΐ����Yh���2�����^=�jF�: ���؍fQ*K�Ǽ��ݾ�$�)��>4�۵�V�Ն�����@V�<g=���e�gt*ה�Q�A�-����yȫ��ؼ���{�٣cb�d�5�1u��f�j�À[�t0oi��gGC	�6^�,wv���B�k]�(��O�3:봋-��;ն�y�3��\_[��f,���c�t��K�i+�V�������d�g+��3S��Օ�-i6�mm*5�x,�-��Ś��^Lڊ�$�{�ds���97Mh�*�6��V��c�B(9X��tmt�j^N�n���ʐ���,���of�X��d^]&�^8��������=��lж��'�V{������9�S�J��ž����/	@<�n��n�2�K���G� ª�|�=��^�
H�w�TO*��{1������,t����o)��gW	�B��6۵���c��a/��>���4s�d��:��5I��Y[��tn�\�����d���H-5�G�}}mݨ��u�!�J��^Ix���9�=/NGY��#�=
��K�T#�9�tY(�:���g����-���+�:��'�-��k�,�k��i� �7݌����]U��V�s����F7ϻ��Qa�ۍ���ܶ�f��\�^�����{ەi�F��+�v�`�Hd��]3%�)[���:��Ջ{�3��\��C��ejʠ ��n��̴����}�,M�����ӋQ��2���#l���*n=�7e�TE<�7�����9�6������K�d�qv���D�o:�l1���iff�6/���2屮3vᩙk"|v"�Z�p�YY�;���G:�t�Mh��v�iT�D��=�U$i5ƺg m{%�>aF�uM$;����x�Gݕ����ϧ�A��y��]�¾��v��j�lny�7�c|���7X̰���L��۵�7�\�;��7�eCFAV|�T�n�[Yr�Qt�+o��97o��ԌLMQ��J�bg]F�8z�=���,�T����)����h��%[���������oy �}ȈL��G9iL�	�Y��L��"5�f�@�ҁ�(���s��0	���]�'w!]�&w\ɔ�']ƙ1(\������)&#2,��@�R"$�&S��IDQ����04AR$����룻�Ρ�B���wp��L�c��r܄FY�&Bd�˕�0��눀4�JEK$6$��;��wn�C6�\Rf2��S���ȥ�!4d�LP����;�!H��w\�"A;����&D����ȉ��)�Qr� l��P�!$�L��Q��u�d�P�sN�ˤBG;E0̑#����1��$1���3	NniK�@��s�C	K���(�s�&Q�ۀ���	��%=t��7s�js0-p�.>NV����k.��-���� څ��`��h�Y��z�ab��.��3yz�L��+��L�J��Y����ϰ�{��R;���x�c�q�IgVz��n^�U���e���i�u�����X��Qs��eJ��Z@���Ӻ_����ë�ǽ1���7��DǳѢ�V��צ�?G��fʐ̑��e����^-�<~�,?9c����w��]f��^��i������ϥ���=��D��Q���K��dmCV�# ���)sH0Lg^C�^�^�>�9u ^}�EG��пz�n|󞸙�QjhT��9�w}���4��Z�{v���%�B�ݎ��޵��x����q�ː+��XXv&��Dr��hF��y��3Ǭ�ϳ[�;�U�G|Gt��5�~U^*=3��N}/h~�X��Ԥ��4yk��eE��������C�����ׇ X�N�Ʒ>51�{��y��' z���&��+a{/��tNln�_�S�$�}'�z�n���ͽ���Qθ��c����G�<ԉ٤�Z�	��m�nHm�_:�9R�@J�I|t����a��6������^� WЕ��5g�4�|�6
E ������zQ��
Utq��X�1����/C�*˰z��*�CoGQ��>��J}	���\�j�-o�n'YO��������e"F�[o��w9ժo{���=��.k9Ԇqo^a0bczݨy�؃�&�J�;]Y� ���+S4͑���O�+6���SՂs=��ǵ�
�6�~N�M�i~=.�������i�-*�!��]����Y����^��q�i���<x�ñ;,e�m�@_8���@�_�MǮ����7R�u����o=8̏��S�����2 ?w���,V'�hw�c
���(ʏH�ed���	��W���s�_��u{�q�:�{خG��F��ng#ܝa���غ��Z}98���,������d�����2�ё�z��m���:�O>��۵Z/��*R��8U��X�z�S7���⩁5<�~��٘^�/J螧����\����꽦�uQ���*c�U ��)��?Q�͒�[sP�LSt��¼^�mCG<{�)��4�I���j��\Y[�|:R>�}�ݑ��4S����,���-���^�[�7�U��H@���
�=2Z�����g!Q��Is�<��{�tW����Ϝ˓��A��p���F�FW���1�>�g2�Zs6}��*��]~�����(���.�ۗ"�U: n�f�sP/p�z?,�o,8F��Jj����;6�<8_�������<��g�S=lW����u7ʞ8^Vu�)⮸OK����Wd9ISA�N\F�雏��R���pR��=��oE��d��M�v���UJ�+=+�əGVf��q~^����N�7����Ҵ�@/
��c�=T�.<��f�ޭ�S��nq�9���y]��9�1�ul�G�͛�}q��bb)��7�|;��3�n�N�o�~3����jGC̫�+��x�
S�s�+� ��?@��3�v��^V酞���^�U���pw�[^+�.y(����Ec�/��>����G"�@JrG��y6E���.e�h&v3v��f׸������7};{X�����3�;��w^�TY���{n���N���ς�t�gjsk}[�h���<�V��>Ѿ�mV����.�ϸ�%e�#���x�w�s�n#��qWTp��wN�_�ߘ��v���s�C���W�^Miw��i���7�q�,�����V3���ռ~�ƴ�{���R�Z���q���o��-�/O�Jë*�2�kK3�7��]�yݏv¯x�Q~t�yV�
F9^���{�-�1~����8v�}|�f��ĕ���T?U,nL�73��GM;1��oW��|��{M�������f�{�M�χ'Whh��J���)����{�W�Y]���Ll��n����ԭYN�B��C��um]H`i��5��Xs�����&��S�]�R�UK�õ��z�!�Y{k��4s�dg:,�w�;!B���Q�&�J�0-��Tt�HT�`|�Ct�[w	�	�-vf�-#R�v���3�1]�R�0Jq!n;Y��(B�	�*޸yW��v#�evG��<.Z�+Pg�ޠ)����E�"E=����o��>9�I����Ч�U�M"��G�zR/IGt�7�����~�Z���Su�r&�vM5�|��o�R2�v�&����;�,'��WC~��g����wMG�����o�"=9�^땻�[����9�~"��)]
�%x�9\����UmZn��P����s����Zwg��=�7w`f��}ݙ+�^���G�^ۤLO����"	kgrc��7I�}z�NH��s~�;�Tӭ!��/����=�QcbW��$�t���0�)�m��{�g��6f��}w�-�pz5y�.=�^!�@����~� �<��$��l1��CY�㱄yG��$�>e��j_��To?Q���q�K���.d���|\�L�.-��X)K�5֝�P�����=�
�'|f�^�&�K�O�v=��T}1q�'Q����=����dv�O�n@�78�g��$���I��Nׇ�3kG��'Ei����f����#��^ v!z�-Ӄ�#�����Ya֖bGq��W�b��A�|*����<{���57�͎�P�K��em~�N���)]�
^2�a���}��	��V�}c���y��pu؋�!pt�cy�_JX���v��y&X� .�UՏj#-ȧ���g��܋Ou�b?��X���e{��5��\����`Tb��@��Ș�:Vļ�V�z�-�����1��w�6@��-����x�����r�*.<����:=X�M�C�ղn3Ӿ=���\G�Z2<�R�jY쉜zd!�UP��pzá�Z/��z�x!�U>��9p%��9�F���~��R�W{�e�F���~����\f��{f����g�9=��әevn5£��Q�ɟ9�ͩ^7��4�������w�>��Fo=���X��uS�P���F����"\��u\��"����ږ=}��br%W�ў�+M��M�{޾�c0"�g����U蚜�F7�z%Ѩ�쀔�șl�o�+��m0�z�P�^�������Mw����~�@m7~���;�p�L������R�z�����6���Y-
�{��m�2=����v=;H���c���XϽ,�z��.�@lթ�O���u�ګu�У㩕=R{|&7�?%qV��9���VG�| w�ˑP���2��z�ԓ�O_�9��1|��,�1H؝��T��iX�s���3�\����4��g�\�D��2j�����I��=5�9��&╻���xe�S`wC�v���k똛��6�N%6I�.ԼT����	*�'�S%�Ä�e;;��J�����+w��bMީ:�=�=������wN}�%�Q��w��ӌ�I���yP���Q�o���U��Ot��:�>�e���tC��ZdTo�|{!zn!;����G��yN}.r��mx=pk������z��(���vK�老z�n������'ä�k�j�c�4O�/PW1|y��r�^n��#�=>��`<�_�Ĭ7_;0�ѕ�a�f׸�w����`�Xpbk��cn����o;fO��S'�=����D�9q3�v���xn3�P�#6�Mj�̝O�I�mw��pǶ��G;�}�X�~�e���f�=��Bߴ֋^ڞ=�>��e��7^�1ELL:9w�+77�3���f��7�mO�v�W�^��{��z�#q��ݶx���H�*=:���*@��[��ߠ��.�`�����ò2gT�ƹ	���걹�?_���o�x��g����7q�[��L1V�ٯYw������}98\EW���,o�3��L���\g�:�>�C�ƫ��K�7^�5�y6�\���[>��q���fo�S$R*v*�<��M�F����t���\�Y��z��<>
�5Y:'9�m���^��m��������ά�C�Vv�s��y�����lbJ�U�%ںק�We�k��bg9�럹�&':�dމ\��qq�(�sJǹ��K̓�8=�/(Վb�1�x^��*�:�dcT��t:��
���<��}�#�,���5!5^c�Q+�c����t��u��G�6Jm��8M�&�¼^�v�^�����9�n7���u�T?JF�O�vo��z�/�U]����<���ǫy�Е�3<�7���V�=�PѨx��[�ZG>~��g}z�Hq�UzK�2e�\����n�sٝ���0�謪O�oA�Zs6_�<m�^C�~�q⸔oޑ���ܹ�����ʹw�N{��{(��PwǮbaz�YN{�FG�Ҵ�@,eB^�=��W錏N��ήo��6ȱ;���=��׸�nd��N�'"KG�麇ו�b�����}ǲ�6�W�x{:�ۧ��.��v��yZ�a��@��2��]�B���z&|��V�CK[�~كX��'�/*��|�#O�Ç3�{��A�d���pS#�4G�%ؙc���6��n�7��Ura9�q�i�q�<}}=���C�N�5'v|FG:a#�mTO}Q�_w�J9q3���+��|4�b�j�	���mhw;[7S=&�3��P��������N��k}�q7�s�}��K��/=jcn�F��t�y^���/R�
��W.Oyd�xzn��*��:'{j:���i�Gl(6�ݴT��4�	��͹�1��۳�f|�UG�Up��<%_݇�R�."��]�3�LL�e�+���I��Xv�eyT�Z��5\�ͳm	>��9���{�\�r�V��_̎#�6�|T���''�N��5�abp�k����Φg�<�7�N"�~�{������QV}T����ޯE�eo�=�H���*�ʌ����8��T�o�_�H�q��Qu�fV���:�|g]2������hv}�Q��zi�E�۵Ʊ]1��=�>	�|f]G����'����F�KV��z}�}>���;�%{"T��M�Ck�p�ƭ�j��(��_'�V��G�����qu�;���~����1Ч(���D�Pgݑ�����b�J�������2��h���~���l�{�S��߻��7+��r�,��?E��;��^2�����>�r��H���'c%�3�XN��So�ٌ�
�9��7��9)ө��Ö;��l���M"X����4O3b�*y���*�g���# �ٹ�tv}߿Q��wfap��������O��p���@�<��B򍥵�1~��8*�g��z���{%��{נ;�fA+�h�h����D_�����8��d�tϥOQ�9?٫�FݪӵwֻM5��<ޮ4�
��vo��$*��置C�gC��R�rC�����Yŏ[��;r;W�hp���^>��v�C\��]�x
c��W}㦌����m���&�md�%$J�GO��L��1�q4)�yMx�*��sX W�m��T�'õA�s�\�ƫ�Q]oq��G���D��et���}F�J_��To?Q���q*g�3�$���1��u?a�{a(c�1�G�3kCì�0̥��m<ˏgԽv\�G�I��:���+��������S˲�Z�4}�B?���|���~�'t�����Y��S%~���^�x�u���s�6R=6�R���,_�~?�2�W߹�b���^F���c��+A�)�[�7��u��^�~9Y�+&=@��m[�H���w�<�=������k�^�#�7��z˫x���=�u�<��%��r��I)����G�o���9����y�!���R�jY������(xڙu�'�)�X������5�/�}T�����r9���=���ˎ�k׏8o��Edk�)��{���fdg-�BՉl0nf����;�ɕ��϶�x�B���~���^��q�Uj�b�tJ�f�����'�y9ܞ~0�ڈZN�6�S~5�C��ȶsjX��{և��3�=�Wq�� ���٘V/J\٣J�cy��/8�85y�c-=|D>�	r������4��ӹmd[ug�����]|�O���-�-�6M��qC2�\���ZrӇuq���w.|tM���=�]�FG8����S�,�0ud�ӈ/��׽�������kz-��C����7��W�`yR�v|�S�pT���G�e�����9�,%���!`U{��{���1�ȣ5�xV$�K��S��{} d�_�<8�5Q�Cr��eI���K_�����SѪ6�8����$9��_�x���½����<�I�����J�߿h�7c�ю�;�����t#�=�qMҿQ^}H�5�~TD����^���:cJ�a����.�#�?C�"��Nh>gt��K�IxTz��]���g�TK�{�@3����Y:S�'8r�u�MTﶊ>�1�=su���T\�2+\�f��9�5���s�����D�_p$e��jl���@�&�J�q'ȫ��k'p����Z�A��Ǻ�'�����?�v�C�1�.=��	���r�Q��$>9���;�f׸��4Wن�˛z����eaG��>@G'��l?Uq����{ݘ,c�8+�t�>g7�ڇ���P���ɂ,c�����>q�zt����y������7��Qߗ�5�κ�kE�mOɟ�}T�?V���g�"�J���K&v��sk��r�q�3V5�zcN��}�5������G>�P�����W/����n*}X�����w�I0�*t}��7�Wzإ �ȴ�,1�'hxu�ٳ$H�����	�9���`œ���p���j.ue��:j��Wzh���ۮ�ȃ%w:W)�6�}cKErDf��T[���	z'�9���k�怜�ن�:ͅU�2���&>����L�Eۼ����V�*��fd*���0r��9�S�j�`ͻ{jGخ/��=�E�^U�1��Β��m�C2��΅d�jjx� ���M�S�����Z7f^=�35�Ck�<�5e�g�J*Ri����|\�3lۆ�tSۜ����X���Bڰm�6�ұ��S�R���������M�y�k/�>�$�F��|fP���p� ;�ͦv�F6�Sߞ�W]��`D嫲8�j@��掭{\������{ .�cѺ�#����u�n3�_p��yvf� j�C��q�LfB��<����p�q��+rt�%��\)�y�;��B�[�Y&JX2�I1�����"7I��-[i�Bڌ'�B��٫N
ǱX�Vl��wME���_��H��Ms�o��7a�@�3f4�p�훆Z����b���u�/[G�Z�lm�˄�ؖ�m
���[<��,��E�2���M=7M-;�ev���
C�1����mL����1Z��{u��D����LZj��7��񬈟�q����v�S��	
�D�`!.�]Ĝ TX>;�ZS_�h�n�p��|F4�u���MN���k����)V�(`tif�
x3|�Vr`�����-����pkhRZ"���f�Oy}�.e�.ż��!+�����+ܑ>%/5��^��byL	�5�ܳgRb�R�\�
I��9�ɬ���!������<{ɠ�6�a��Su��լOM�>�5ܬ�#3��b�0�,4sXp�u>t%�k�b
�R����	�I9�tW�Nű6�Y9)��z��b���6������0 �o!=#{V���aw|睂�λ_N�G��Z%f�ʚk@R6bB�b��Ѷ���Ƀp�ct�
��z����{���:��
p�"�7�=�{���o6�(]懕��`bY�T��F ��l�0N�ۢ8ۧt6������T��d�C��)��:$p�֠�0�����àJ\�Uv��%��m���3�V�/)^��yP!'����N����릗j'������Z�J�q�ڢ����+����9���^�Fcw�k�ݗ�kseJ4R�ۜ��5r3��%�sZ7(�����-�k������ߟ߿������)�a<v!!]ݔi��A%�+��$&)&E�ė�)��`$�H"dQ"s����#f]�1@s�ME(F$̢&`)�H��3&	����7
1�Re ��!!���)�$�Ma14�!%F,�A),�JIr4A���ww!�$�LLD�dddbS�g;`"��$h���`�SDI,З7H�fH�9��1�M�����h��,��h�A3Jb�D$9�h���)H�H�Q�2`%)��R�	��*4D�
ad,hCL��b�4Q�D�M$h	��dŊ�D�
K
A��S#d ��Ĕ06J(�FĒB�ˁ �Qe˘DLc&��0j$6B,67+�bF$D���ok�p.���n�m�U��˾�CU���=y����,hq���.5.:���wn)��jv�܌���Fo���p*�B��Ԅ��#\��e�Oﴸ�5>���~'�ӌ�(��7�j�n<�`�]I���r�-�\�����.6������29�Ϧ�{�~��x�G� ��~�K�����ѷ����S������l���=uL	��0�grg�^���3��F���C�fD�՗=o����e�-��~�q�T|c���F�M��e�'��ҙyU��F�>"sǶ���X�[|P�t�z27�+�g��{�ë��8�g�C�  lMC�1M�&�G,�{�</R��w��$0<���Q�j=��"q��;�>To����ϥV�e��'�n}�k�0��Y�P0��̒�J��Aܮ��h�sj5���^��?IE3����_E��ȿz��[��VZ�i�7;6���O�3��h��uP�*Z9�����ﺢ�s���߉�%��x�^1�mӿF��{{����9 Tz��غD���tdA��;�Խh{�*�0��+�&�|3'��2�ZU�Y3�8\/fA��Mz�'"KG�麇�>&%��*5χvB4�«�B��^�o�V�rE����8��[Ȍ�{Jw��n�e��˨�v:zd�q��Wu���շ��oRT9J��������r�W���x)�zd��Cz�i�y|�MeY؆M��5}i��A���I��nt��k��k����\V�]���8��=0���6��o�9c�!ú�&��2�������4�/���~s�pP�YTB�� n&|��M�>��lW�f���:���l!��#���$��4{�g�c�Q�~t�AuC|r�+�IG	c�`͇����}0:۟y1��{k�o����������~�TY���@~���U�լH��pOR�@��ݕ�]b��G�����t_��V�q���zX�L�eK�Qڽq���W�Rx��:�v�Au���h,�3�)��
�	x}*P۝�2�kJ��
Ӭ�������N�
�=X�խJR*���5�dZ�Es>�p֚|�AG�� ��ҷ}ic��L>�t=ȥL%�i̸���#k�(��=��SG�����#�l���e}'0���㸮��ɝe�$�k��ǫ���^tt!>�����v}�������;�9MW����)�9N��0J��X��I=3>��j+����~/6���>�y�����9��7����^ܖ_D?Q�*|۳�6cgb��+��rK@[�E�SrS.�h4o���=�����{���s}/�ϯ��V'�T������� �hA:��Pӆ~Л�з0P������N�k�Z.gv3�qu���c�7o�g/��}y��~�����i�"��Aݴ�si7��6A�c{�e���Z�1�WT�"^m�)�����\��ۓb�0�u��Ξ��]��+ä��eHfH�D�h�,y�P��yʐ��ُ=Z�oݕ���c#ގj��u��GI�Y1-�0X{qT���V��x�l�+j��>�LO��$q}{��O���R>������"�S���-���^��D��S�������(*3��o��K�]�}�}�O���~�:�7��X*�}z���&�����^9Ot����/r�L��Q+�G��3ݐ&��^����@yc�����W��=3��x2Ƿ��b|�vx��XP=a��������>�Д�7	ب���6_��:|�X��>ۢY��{�8�������߾3����r���6�<;�=��fW=О]�������GuB�(v�Z��Ħ/��� vQ����>go蝯�;��:+M��_�����~��,�[��uu�����ٗ����(��4+}�p�z�;%��f�W��q�5��� o��J^�oq�GH������ _���h�����
�5�{����:�*��mb�5�G��R��t�v���=������`�Ob�!��t�]����������~�c��e��7I,����$�c���rv̥k'7����vR���κ�<��O�g�-s=6�xu�s��+K=W�(D)�4���_���t��zU�c�������v�_y�b7Ϻ���,m�3�NƧ�X;�2�Q�<9��zp�^���Q ����	������^�q�x�{.;���;��QH]D�~�ȷw{���ot�x�^3a���'��\z�e9��ڕ�y��i�~���W�O�t�{�dz{h��Ϲ(��B�|�c�^�"���l�"*y_\��}�,z��C��3�tW�8U�	��7f/��f��.�Y�@O��Gt�7���s,��υ;6T���G�e���+���
����rg��}�^���Z��
	r�=^4�[�N���ǆB��yd76J��eI��*ϕXW�0�b��v�>r!̜�B�j��i})�{}`p�S��x�<��=q2fȠ0DAk�s����aωh��	�x�i\S��x�N���� �r�SʧDL��77�]�WR���L6��H����;�#�^�^^�s9��9��W���ت=V�UEy�֪x��V��3GMK���=ei���|{�6ӱq�׍���l9>�h�@y�R�qc3뫫;ů�i��[#G� \�ٙ�qNĘ�㌨�!�1������Qx�9��ǖb���b�ʹx(��5����_6�X�r��o88�[E�w^��:��w,1�o���7��쇝��ue�X��b��xF�BIYOF�7Q{,�[� �Fr0+��9R4�JK�����&�N}%i�>G�"n����.�'ä�k�k��ǌi��P��t5�/�,�ɰ�GTz<�k��ڱ�.d�@J�r_���^��0�3k�R��F�M�F�����G+��N�9z��/}H�����P���Z.;�'�\L���ڇ��<������
�l�Lr�~����`����J]����K�sRv=��WN�{Mh����9j䝩+,'��5����ۇFKW7��o��j}�W��߶q��z���_TU�ڏ*�G8�oQx=����{�NN��W�����&w�΄����~=��{�d�N}T��<��mxU�Y�%��Y�*(��\��D��=U0&"�X���n2gȼ�wa���"�ԭ���B'c/�	ڊ�a�����������b��{(��(�
�nM��⩁G�/ҙr:���.�n{���І8o�
_c{Ձz
Go��aU14{��p�#�=SD�	_�U��ttEA�p�~��QN_ {���3ٓ����3�l�o�}ǲ7����x#�YN�nzk��%�aNߌF>�(��Y�w�J�KF>P5�����l�9�D��r�����vp#���;�^���(��';Pl�Z0�^����&��8��:���qe��r,KyҰ���W��۵$W��p*�z�=@��P��WH�v���뭽���x\��p�ՓB�;�`�O���mCF�x��_;�6w���S;�z
���A4tL�B����=��~�=�d� ?�U@3�o~��3e��J���u�����(�f�O�}fJ���(��2�7��ˑQ�t@���10�Qt��s�:2�i�^���t�K�F<8ף|�/:ɏ{�9��N����˹�QD��ޛ�}y^&&"���k����t���"�;H�L�G{U\���>t<�"\����^��ϑ�S�+t��|/�0@�=���|�\�^�>�q�ƭ�A��2x�!{��wc�G�(��rQ˙c�oH�t��#�m{*�������ۻP�3k��/���ۇ�i�_���d-� x߽�q�����=w�L�\W�݈��l�x<'�:���'kgCٞ����9{c�Y�}Ģ�!g��wB}s�$���g5C7�;�S���'��3gi���Ү2|+Mƹ�Ζ^��
>26v�����Gr*/��X�Y`�5��]k�܂�W~cd��|�wֶ�k��3��/�}��g�+���Ni+�Np�6>�׉˚^s�a���Υͮ4-f�~��a��ݭ���|@B�mr@"�	�sj=IN��%7��Wv��f��7;��$���m���e���1�JI���ܭ���k3R,��۪�����뽧�D�m
�E����֙"�1�W������=�hvG��F.1��D��z���خ���/]TdUȭ�S������2ǽ�]�����}��=�P����AgϢ���a)�Ω�9Hκۋ}bVV�zn���|ϳ��sϮqu�;��q�n�Җ:�{�I�Ԭ�z��5q�Xk�,�l��2���7�Je�ڰ�u�Q�=)������7W�'��@vI�T��锾�>B���}p6Hl��̑��l��s
�+�M��1M�Ő�V1=����*���}�iy^�~>�����͘(=��Th������̍�yB�^����l�C9��+ު�X��\�º!�\H�K���G�"baz�����Wl��aҗ9D����,z�����~����Mx��yǽ|��=�T<�M�Ih�D���מڏS��N�:�kYs����<�Q�ґ�τ��Q���3��W�}� � \��<�]2J���3*��뎯X�w�_16=�?A�u������))|S�1��F���@y�pyˈ��v�S����������e��)���wDoP~�Ḟ9T&��w�9H�YuNeF�df7�lL3�����]{S�vw+�h�:�OgHo3]zvga}L��NP���Y|'l=:�K����9��lݙe�b4�f��ѵ�l%3��f�%����7>6p>�����c���=P�fG�wg�
��9Y��0��^�[6�=H�#{��oʎ���9'���ׇ���>��p<3<��S�d�VJj�>اI��;vd%M�`��`�{�V uz�5����S���#�{�+����z�y�n��e�.��c�z�pX��k�u�~�@�������57H`�{��<���aK"���qBN~�^ة��L�B�GѪ@��H���w���g�}����_�Z<�J�eW�o�d���^}�ӊ�n}|6�=w�g}7��7���r^�q��x���7Ƣ���za�f�
�R7r��vz�>��"�4<mW���\;��N|6J�Sά=}��)����'l�1��'���g)m��}�j�s���+#}DS7���S�"2�ȶvK^^�=x�`VxeE3�}��_���x;H�yO�ܯTx�u,��q.��-��G�&[(�¼^��۸���vO���(c�;϶�P�{���!+�f��ڇ��G��
�zd77�=�ʓ�E������3�R/��4��ь��/�'̯ =Ϩ'כ�h.̣z���f �{�f������z���g�K��וԝ���(��1J!�7�����ƾ�}�Ws����zO�q� R�4a^6�ufL�qα�mǳ��<��z���c���%hP���Ħ>Ĥ�_�O�y���q���p�ԑ������_�Fz|j�<��Ū=��7cs�QY5>��π�}�\�Γ�	��P�z�u��>��p+#޾ ;��Y_�'�fi��ghY~�P���F���U�"~�=�p�p���/�g�U^7�����dV� K�_jHV�3ݹ`T<�tQ�3���c��G�.V����#,m��ٸ��~�R��.c�R1�ۙG�ja���%���n����+D�#�u\FV�w>&��:ߣj�=y8}ێ�깾C�̹�h�]q�9���t3� � 
�Cݵ��en�p�e��>����p����pNx�槁��/o�
����ȅ�Ƚ�"z��<�N�D�9s>Go�b]�1B+}��%��V9��ͪ�q����g[ W�m�߫�Ga{2
7Ω��hDm�ƀ��꟧�5-��?%R˥k�6�p�T�n����g9d�,�g[��"tc��K����9���^��[g���#���Ճ�p���O�,��g��)�1r��<	���+���P_�F�x@��E�5Pvf!�ubn/��0��Ƹ5��vOj�9�U�T�IK6�3�cvL�|���=5󷽏��+�����;��<h~����Ό&i���T+Z�V2\���t�����m_n%��Q�.1t��	+7���B0SG����N��Y����z����}nw��^���N"���l���=2�Ϯ{Ō'Y�}�ˠ{<�K�F�ϩegOu��N)H��{��w"/��*mTc�Q�{�T�ɴT�S~��@��R�į{/7�;<�G{h�GUC|e�cK�`������5H1Ч���ފ���PEs�I�c1H���pL�p��6;��DmCF�w�G��W�t��n����~���(��z��`���ƙ;��o�oL����2& ����9h�sj5�Į)ϩ"��J)���N��J�H�+����\w;�Vː=��>�� y����v�U
�.|�@aa��e��J���Y�,�j�'ޞ5>[�arЩQ�+'��L�����uN�
gzba~��LӞ�чҴ�|�8���v�BT���{F���1�>�~�>7{�P\<��ND��_�u�2�LSS�O�=�,Q�,�Q�ű��Go��6��r|-�k�7�g���U y�K������]�2��p�<^WB/��<�'�V�U�5~.�^�E�� {�uC|Y�$ly�(���-P+��X>��lܫ�g�a�Ṋےe)h�GdOg�eC ��:�$�@��MW*}�+J�'�Kp��4��b��涞�	Y�g���[8_ұSH��6�Y�zw�v�� ��ט�e8h���v sdR[��VG��]Ŭn�A��� X�&�WN�C����L��[&�$�(�_E�"[���A�]�z����y���v���۷x���̒� �d3���c*ЁB{o��>���������'�8N.E��d��1�vk%���H��NmkGl��5�y�u����0��Z��u���w=`m>��8�����,B��2�|��	��m�w�Cq�ʒ:�]�%*T]L"��K��q�@�{��c�j�cқ[�[��-WN���e.���nŗѽh)�ƹV0�4@޳���<��F`헰b-S�:a�u4�1���&i#��Q��Y�ѹ�mmF���f��]�p�Ƕ:�M��$��Ƴ^Z��7�ɖml2���`N�0cxn����S�[����1�P�7Y�ٓ(�>m�>�Ipv�n�}�o:��;�[�2n6c�s�N%�Y"@L��(�z oXy�2�_+�ge<YΞ�*ДT��>̩4-Rj��ƍ�h(�2��7:�(W"�����ڕn�u�����6�l5�)�3���(�݄a��.���P֑�E��88�ɡ�Wf����^�}O�)n�Y/��*���rh�`�o �lS�/���R����%��.�$��݆�}��-p�ȫ���$��`�.�ug1%�S�wE�jٗ&���%^�W������i���D�w��m'�}�f�a�e�YH9�����j#`�Y-���s|0]�Ӧm��)�E�n�"�S�{�^�pfj�m$��6�6�ݖ���]�Hގw�QIR�3,��	P�=���^V<m[o��gE�1wV*�E�R�����W��P�!��70[�C�����l����\�=��S��y&��x"�Ss���/:�ʺ��uZ&{�Z����`��;�u$w�8l����'{���gE����XB�V`�J`N��c�IF&�m^ɽ]x��)ُ4^$���O���>���$�PnK�U�DԳ\Oq�嶷n��OBn���<fD�E�긱�w@��٠�*��B)aᙃ��Y}��"�PQyF�%W5��kx9��Sz�T��)���Ui���|�*����3NeHq&�[��C�<���y�>�g��,��=%�M�AE�]=���_*�q��PpF����dec���c��t�e$a��=����w|�]uJFU�۱�l����4f^���\�U%X�wy6)�C�lQ�Zh�e���M��QpX�)E�u74�n�Z��v��Vo+1G����1�䀊jэ��v��t��fd�QpY��ħ���.-�]]Z�Fr:��F��3#ض��i�t���{q��@%���u|71p�]Eκ�P=�l+
�T��y�4���q,���m+����>�@�Q�L���i�(h��
�@i1%AQɐRIL��c&��&f�2&)�e���FBH�c(�\�%��i��HA9����b�����2C,0�(�5ɖ%�K	C"�	���ɴeˬ�i��`bD"��GwF)�G.("����d�,a,�"b�7DFC���	������(ѓi,�0�Q�JC 2np�2���%b�dd��$��4�̰ED�4F4I&�ɣILb��bQ���H�&�F#\�,h(��r�42!Jc	�f�hLS#F1DB�ȈѨ1HdɬEK���h�ߟ�������V7�֖���M iI��t����L��18���+�Fg����DV^%[��f�����MsE�������W������n�W�'����f�w��������/eF��vdOLCv2�g�b\���T�C�-�>8J	��~6�����Ǻf󥀶�q�zk�D�~�.�9J}�6��#v=��Ͼ{�)Oݑa�uXڥ�pË�g֞����\���gK���L���O}Ր���p=�x��Ni\�F���#
��7'�RȪc+�������<����7�p}Q|�����7�����oċ�z�Ƿ�Z;޺C{�l��=4�ȓ�O]T?P��Ь��R�S�U�≝�'��mR�ю�����>�:�=��X
������%�tiN�j��˷S�=~��U�V���'�MF5�p���f;��څ�O��<�w��_�uj�s��r�W�5#�z�wE^�7���Q�@,���i��g�Vd-*<ߞD�/Sf��Ieq��ޙ�~go{����=KH�yV��@l�ǤS${>�My,y���O����~��1ݙ7
����a�D4&r7�4ײ����IcLʃ�T��į�"���N;��!�����ѩ���Iz�8+��	p�-yu�,q����'��DbT�u���z��\I�����/�z��$��E�{��0}h�S�7����$���-v���ׄ쨮���rI��LR�Pᣔ���@�o�\{X�&���joc3'��|��5m�M�]�X��J.o���q�̉�_<f�X��ۉ��ꋤLe^�=P�nׅ��Z@�s<'���$|2=J��=;L��_ �=�S���R��NZ�Jb{�z���&}�1[��8<���L<5�¼/�U~9��0l ��V������x[���S��D���͏�͢=W��5����"��v*���6��"27���!�����1g�o��I5�Y/r�.&������6�&��cL�.�=p�fG�al�ܗ�(]Lz��Q�f#>�S�Iҟm�8�v}��^����5�_񥍏Ɩ;��X��?E��ڣޢ�^W��_d1��W�}CKۚ����pa老v���yy^����Q��r���-�4(Azx��l��}���7�������m
��Z-{Mw�O��Ւ���:t���.fc�p�鎷;GڤmT�����9������/�墐��!m�G�r;}w�<���O&ŗ>���<'}=}3��5�_��}��c�q�zb�b���#<F�˅l����P���[����}�{��󹛗����������ޭw£{��[�����OΣs��l�x�Q���J�Kuo�Rӹ�������ѓ\�Žݶ������H<ݗޭ�n{cǞ�(�r�F��ޝ���y]\�W/1���ek�����Լ��J��K��Z[�)g8}|��Ln@�W�$���2r�z�F!�^��%*���Yy�"��R����1Sȋ>E����n�1��z�0�_�yZ�c�+����tdo��q����\ת=�eK1��S� -�#�2�D���HE�p���ŏd���gz���L{��i�~�6������{��\X��~7�\�c���F\���l�JZF���$s��ȍ��¢=����x�:V�H�籲�˹u�ƹ ���B����>%���@�~5�6�Ed:W�7���+�5��;���t ��9's�=7�'|@������<V�`�z�Q�i���@vR�����ߌͥ=d\{�P����;���<��K������^�'"f=q7Lu�g��YZdn��Ȅe��ǁ�q��u��=\}�~v�Lc��OM��z��}�D��]��>E_�u\fއq���l�������v����3������^��/�t'��懘��F}�{�\v�j�>0�4���f]m�b�)`/�lgraV;��#Y�<�e+��M̯؆ů<l2�o��3�i��6���K�Àl�]@:5t����J�=fv\��|�ʇ�H���nK��N�z̖���q�4:�ͦJ3-^,�a�5���ZThC�8�_�g[�qnQ��}�V"��>�1~���p{����������d���'���b��Мމ:s�:���׹qU4M.�N����ꅆ�T;ͪ�z_�M�u�B�v�~�e�뀍{���&Gó�8^F㦽�H��[�>;uIp�3�X�.U�����a��J^���>'�o�� V9�zp�b��c����}�W��i�j*���{b�Td�J����g��)�1j���}���Y��*ށ��Y��my���7�k��-���9�-����z��`L\���:ϴkT���5C2��ާ<��f��*���5�{��;�_��7�\md{�<a\o�S$W3,�Y󬉧l�j2=H����+#j�>2���_�Fo�WϽ���Wh0��Q��P��z��q���5���O�~���[�d�F��چ�|��q�g����3^	luh�P�~���N+���S��љz�a�Ext��% �n��)W~���>چ�}m+��u�H�?IE2���zt�Cvǔr�F�������3�/���L��J�Qs�sai̍��Q����vq��׀ږ���Gw6��/Y\�}ܣ��UwR7?MT=qW{|������ѥx��]M�%,�Xy���m�t3�5r��T�@�T(����N],b���&���t�[���E�VG��ݓB�E�L�=�a�,�(��ҟeOZ=˔Lm֔u+����S;���zO8۬*�.�\���]"f��������4�,�E^闑�0�k���}R����ŗ��L�O� W�dy>�����S���{<n�#��`�|��W��G��/Е\�-�U����%��=w T/x��g��r��y�U\�ϔz��	�պc�����W5~.1<��G�ȁ�2/��)�D���b��뎜��'�P��/�3��pf�x�n�<���I����O2�1z��.7ԁ�<��;.݋c���9���o��Ve}�H񸗇a��x\��ǝKoL�,{�s��[��OXb���|.�!{�>��vO��������������Js��^MiW>����L�D�^��#��]� ����tn�������r
?w�6@�~A��wֶ�f��l�un�߽��������u?*��tb�x�q������G\G����IF[F�9'0�������W�2�{{���A��{u�y3��,&�iَϹ���>�z��o���Nj����h�,X��U��)9���%�p֍���7%.ו˳s���܆�1��ϋ�h�f�r�N�Pi������t�7ٮ�z�y�tP��ԯM�Q�F��,����L��eu;�]BJ�7�-&���=�<��2[�vЕ��F�ed-f�>Ć*]�o8�]��8{���]��ȏ+,�ol)�5^+'�&�鸚�k�ø�)���P�mRk"�:��Nx�_f�s�؞���u~<xnﯶ�(���V��<��wO������\�*�ɠ���Ty�>�Ϧ����j&�o�ym��Z�:���z}���dB����$6l�m�T�-e�3�6XFC�Vē[�7Hu���8[��+���{�6
�i���a�{3�F˓�y1-�ʩ�+�a۱��Q�Dꊊ���J,(�|���*By�w��R.w�j#ۙ)�9�_�������>����m�h���wf��BZ&�x|K[;����#��U~>+i�ߍp��"bצ�e�L���\��Ş{;t=�_�@zk�bbb�V���ށ0��ܼ+���W�:ə�z߶ z���m��|�ږO�X[fl1��D:�Vɯ��>�x�4s�Bc+��ٚXa;u	���m�^ �G�/�|��i,x����H���+�ͭ�'|f�^�&�K�N�yc+{N�����[���I���۸�;�g~��ӟI�;q��z��z��X�X�5f����%��+�Ԕ�e�����o��$�i��X\1gJވ03������^h��oKr]x�M�b���?>	�a]ke�;��o�/	
��o��N�09��Se����M
xn�ɼ�g��{�����(n�A9�ւ�Y&L�hQN��t������V���lxo�]����q��w�,57����JX������fc+G�����,z=�Zn#z@�_ݶ���V2~�|J^�
�<�Сo�֋^�]�SQ���^}���:]��=��+j���β7�#�\.����o��R������8k�3���*�(JQ��^!涧ǲg�c�;ɝ��@L�u;��k��9����ޣ�^���}�Dz�^�gѫ=|2�(��Q��f����}ꇱ�)�a<�}:���/�:����!�Q[���)�)�z�6�Tm�5e���"��� -����"ϑl�71�#]~�;��
7��ް�
����p\c�Wq����u~��%�ע]��U#�j����%��ܨ�7�#���3�ﶼ<��k�v�Dy	\{"7��W�<:���2�5��E��d���}@Z�t+���ɏ�{�}��mCT��f�C�Sg̠[�����Z�Y�:��/�,'�o���d�Gx�� ^9M
���� ���D	��U���>9<
혟zh�"��3��{�=��\���IL��=	�6�M]K4���=�h_3v�l]´�D�ve�M/U�R2ٱ���M���qR/�P�t)n�o��;\���1Rܭ�W����h���5hH��Y��}�8�[J���Xt5tZ7)�f��ݟ�WvYɟQ
C+���c���"b������%ᯖ��WBY
� ��Or�^�>�L�5&��Q�e���Y�3����I땦F��;��]];"9]��H�2�r�Q���s·��K����;�M/O��9'���M�5en��$�?i>]ڧ㡱2|�����!�N����{##��r�x�<��"}�Oa����u��B/ޛ�����7�ڧ0�z3k�n9�5��r�_�B�Qdo���U
<�V�Zr��Y&�������ǋ+�3�:vaY،}Q�ٜ;����ѝV����q�W{��/O�X��cz�$�gr5[�ǡ.��d�ۈ���o��c2v�vz�����KG�7�z�O����Y�����?.��z���Y�'U ���\kO�ȃ��.1>Ŋ�;���n���;\��q��0ጫ~������v�C�l�;��F�^���l,��}nZ>�j��߀U�>���D���њ����BΏ�e����vG����O����^���Fo��|ado�S7�I�Re���P2����X������hd��@iu�?-|�}2�]�`y����xujep�nW?�jޛ���W|���ھm�:{Vt�6țLsYVVrY|MX�N�N�Τ^���ə6Ba����╍xT��e�|/-m�3yd�]YYWݪy���� Z>~�S��O��K�����[�^q*�b�δ{!�����ᐅ��N�j�;��t�	`j3"��D�a^/sj5��uǱ�Sg#�'û"7����(TU�3v��כ�:}��d"�	J@�O�ȟ�U�ߥ��ȅ���Ī:�׭#�k�]�xG���ϔ�+O����Ճ��>��<`�v�U
.|�@aa�/Ʊn#�|=y�R�������E9��}��%��qw�ˑO*�/��!����x��	�+���A6#'wv��M�m���*y�%O��ʟ�r}8�{2�>��老z��W��Y����j�g̘n�Q�F�\{��J�K���y��J�8���
�^�L�#K�ǻ{�׹蛨J�2�L;��u�kO����	ПB�]�s�@���]~�\�zs57���VwN��Vx�=���3��fl{�7&��J������n���~�TY
�ޯ>�v��^�j��y�h�������ʜ7�J9s>M���a�\�t�i~='8�_U�ި�5���6�3�Qf��r�Ѳ��S�CV���Iʢ�V��X��nYˡ���f̡̭ 	�gvFh,�R���AL:�OR'��J�]u:�:{�Zך/x�YJ���Bu7�PC�-���GI��g��/	r��g���y�F=�{,�������g�Mp��ʔo��P��t�Oa></�c�����Z�+k����vp���rg���3�mg�@�4����?W�q�4��A]��L�|�}k��9�z��c'=�;f�v[�O��Kg��w��{�U�ċ�����ǲ�u�{ט�o���b��l���$(�E{�v=7ޅ������UG��z鋌��ɟ��o-��~�������yU���Tͧ�F�V���;�wx=��ʍ9��M���x��\;�2��u��\<�.��#})��Y�T�U���~�B�έ��\�pc�mZ�2�{!���fPf��,	�n�U�"�#&���~W�W
S�뻼0�<����Z>�sN�ϼV��[���(�4��EHo誑��w�<�Ǿ5ϴO�9��C��϶�S�������}#M{-�;��׉b�b[7����*&�٣�oѓ���؊'��i���9��+jЛ��׋���ϧ>ٜ��1�7 Ac\}c�k?J�Zg�C��D��	����ӐKGv=�*�,d:�e��7Z|��{�s�6�ֶ��V�Z��ګZ��Z�kmժֶ��ګZ��j�km��j������ֶ��mU�m���V�����Z����Uk[o��ֶ�Z�km�mU�m��V�����Z����Uk[o��U�m��V�����Z����V�����d�Mf
�|?a~HAd����v@������xʠJ% ��T��D��B�
�)��QB�8t�!(*�PAB-�J�U"�J��*��J�d	��!RJ���J�TIJ�%J�TEP�T*(J	$J���(�ۡQ�����B�`��if���TJ֠����R� 5p ��) )�
�n�� n�  �  f   n���k[���Ɗ�
�Y�8� ��mHm[Y�7v��@kk,ԩ��V�l����Q j�c�0����-�����[�@袕�9�d�wE���l0�4j�E+fIk�pPQ�� mY�V��۠�ћY�j���]��k,�lKj(h[P֥Y(٤�	T#���94��T�"��
kF�Mj+FF��tΫA*MB**R����Ҩ
�k4 �Kl�1�*4V�H�k��4�m;]��ҊҒU � [�LSB����i��f����6���B[h���#K6ҩSlkA�V��kcMj�-aTڱKA���!h�Hn 3Ut`X��ek��cJ����Uf�J�e
�=  ( �T��41A�@�A�1��a%)Ud�ш�F#�49�L�����a0CLM0��R��10&��# L��Q#@M22�dȓ�<�����0�ڐI��Ti� F#� h�>�'��7����|c�2Ɩ�Rm�UW�	C�"*����������UZ)�!AV����>������*���A�(*��?9EU�� 
�#%aV�z_t鵊���˝v`

���9P�@F�a��L>�;"�ye�H"��M{+mx֓J�zZ��5�p( �Rf[D��3X.�57]�&Zv�6Ѻ�**��۰��"���gIQ�Fh�5��NBn)S-k��a�����E+
�X�4	Wf+6���2�CF�p�i ZSkLl�5AE��L�1��l�)ֺ��S]F�cm�ܻ�25,�ťK�]�$��f�n�bfm2��Y�J`�"�i��Xj*.Cv�e�_ky6�5��U�7T���n2�`䵵z'�=�,�Ә��ª+$�l]M��5�c��G풙���y��i�c~�IE�9(��,�IC4��[YM9wZ3B-䭊I�1f�f�Jw�UZ4�X�@*e����e�c�¢�N�CV�U��Z�&�Ph̬���Q�	r�v��"1Y,]:���RS�FVGSY)��e,�{�o-�-�7��0�̳J�#ejj2^U��kZX���Cd���v$�@���.�rk��.f<�֞��&���v��P`K��{1[��-d0�+FnGTc[	������n�ۊ���RZ70@l�:>RR��,�U�W�w)m�kE�5�r�Zϖ�f���=-�	�4�K{e��3��&�i6�\Ũ#�xE쬻-ۑ��b-p��EG�A�n�dP�Q��Yw�E�-���h�������j���H)F&i'�n��T2;�23�[ʘp@��m�z)�PI�^�U0��g+vS�ݨB�e�;LA5�ĴUG�7�Y֠{��O��wB�PN*ܶ���(Su�(u7�a`�+N���	��@�,�1�B�Z�`�)V�������`F��R�T5V��!���ͫ�{M|���&�$��p�6�IRa˺�L���vT�����P;���N(�<M�s\�.����'Ch�0l�`�&Tt��1j�.��ޛrj�rJJ�VoC�I�kl���"ڕ/䕚ǥj�G�L�O���i�؊�nP��R3B�[�-誆����,�S\�Ҽn��7K>!�RTN^�H��q8�����v[F�	)1#��m�e)��Py
Y"[����B�.����7JGF-fE���";kDrn��a�J)��Y6��"�w�����+.��Y ek��)R�k`ܒ��2m�ޥ���O�J��gi`��#o�/P�KY9���Ӛ-�Ǳ���o6}f;b�cô�ں�#Ix�f�Vk�v0�N�휬�b�=���v9b
�é�K* �٩��քJ��VbuWi=�Tͣf�:��E�]mȮ�RC*
�in��(��XTgB�i�����`0Ǩ]�MV���g7�6��[�A��1c2�8+K��jm�A���1f�/%"j+l�n���(j��mm�ӳP�Pa�%(d�#śz�w��Y�T��ckc5BM5���h�3��9��0)ejגn̒�f��d���T�$̧+F@f3��O[X�xM��0�5��>Br�������uP�ӆ���t��q��Q���E�����%\�[Y(�%�L]�uw+pSso�S�I5���-┭���k"�
f���Z��Ӥ*	�F#"&��M,*&�(���J'c�W[���na�˼�l��P�R�AM�%��1T�q$ͺU�n����l����z&A��ȷJ=r�$Z	;	�fT,ة��6ɼ����*�1,�o�:��Qm��ܷh�������
�8�����E&��s�
��(*Y��A�33�`�j��VFVM���>w���m���%�;T�fK-{04��U0u�ͽtRQ�OUm�O������c]��@	���t�t�Xy��ZٲlEc�3\�u�PVTRA,�sl��j�SV77?�^
0!(0Ve�c)�$T�i�a}�杆d�ϥ5���p�&�/�%V��Q")�����i������I�ն�w"!�Jv�	g3v���n�-f6�mU��x�|�[���~Gl���i͸q�~R���V�{(�Ǭ@��f�ѐ����cȂ���
���r�SrU#jG�����3^k��F�i8�	7kC�Z઒ò�h�Rct��[���y���X�.�M�r,R�p�u� ��
����f��K6�lY���H;Pl�V�,kӷ�*xK�W��1���{���p۪-ʣ��4�b�c�sB������#�Ol��G�SV�^����p����S�S�.�x�bɕ��-�w�6�)���U�ې`;E�0S��[��eYD����ȭ^!Vklm�5�-�i�feL*�VY�g\*��ƒ��Pm\�Sl��'�nR��<߲ޒ-�V����=�Gn&Y�FIz˹!��A��7�%�U�h�����IڻpT�u��iOЪX%�	���X���C2��c&C���TCe踖�u��ɓ3cbܫ��e�i�d�_����Ӑ�Wq���X��m�(̦�D5�x��UUX�wdܵ:����0a�9����Y�}�uк�VPM:t�EVu��e��x�%5�lml�M�Y*Pup�<Æ=;�eQr*,�@Z��[hݣ��{���l�asa"�<�V�!�ՒS���'Hwj������a(޸t ܷ�V�l�!j0���(�c+e�Ȃ��u���s*�S�I�ųN\"�B�����a��nRQ���wYW���F��v�bݕO%Ȳ�Owd`�#)QRcr�Ӈ�
�tu�hiV��Ţ�)V�aD�l�м��R^2�ք�-�V��f�+0�整��(N�mղ2��j�4��^:�:���YP]�??�J3Sڊ�C�Z��䒙����k,����nJxZL��kHׇ/$m��J��V)l��Im���VV�w���T4]�n��%kt�X�;���0'��S�2	,w����DQ"��ƪ܇A��9���0qě�:أ�VqP�J�Lނ�#�*�t,�	̔SV����񱌍wi[ ��3�nV�v�����laTZf�MFk�8Tz�neQ[�7�
��Ðgي�
�دv��+2��8�@+;�z��]�s.�H�XL6V�����Վ$�[���W0⡡�^h��e`c,�X�h+�$�2�|��-�]Q��݊Ip]
�9[{v͆L�N��y�\;w�*���8�SdFؘ��8�T�r�UUՙ��,p�rVi,--�T�,�3%-��e�n�d�h�C`,1PM��6N�6F�R�N�c�%e��q�61#{ʸzܤP�Эͼ
����Qm&嬦�X����֖�V������j��ɣ�Hֲ$�v�b��kΆuAvY�B5Tm�c�33f���r�P��lKi4�t�kn��&[�	�˗[�����Q��/vml���S'��X�:ի���3@��J�i7R�X�Fe�i�Nر&�� �K����E��-��r�	vEm���ɗUob�t�aܬ�i���N%J��irf�)��);��:�n1�JQnc�cF�f��%�Z���`�⻭*V/7�^�zN��b]4*+�
z��8�T1��k����ɮCYb�6l׳�� bI4���đI$�I$�I$�I$�I$�P�4A�Zh�ٔN#�&�Owoe*4r���I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I%�	$�I��I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�E�q�t `,��ڻ���8Nv�bUUUw���;���g�:�[��F���3��r���O9j�a<6%?�x�:CS���	]��Yh�X�bX�o4�m˲z��T���I�**�(����{O��z�����o�f��MX���A�}��|�DSE#���wQ���)3��ٛ�#���&��rOz�SwFA�#9쾛����el��w�)Q�P�j�ҹ_����g9�{����ޕe�e�)�c&�E��Ftux��'1IA�Kg�6BY5�)漩X�*�UDf]��3�KR�P�rS�s��W��R�ne;T�e��3nڬE7�Խk*��ˊT�N���F��Sn�$�D��p�ɋ�&�u��D����"� j:����ڝբ�4�/��(6�:���=Kx�n��w�]�j'-s�!n�]n���c�2�oX���yf|B�PK �Y]�6.��ZW���r�uFt(�����	VeXGrr��us4�e�-��Wf�tZ��	��c��I���8z1�N�l�{��
��C+�D�d�wtкwkxN����q[��ɽ7ak1k��ʨU���v'�tUgCi��fI݁շr�A:v�+s3�=���Z)\�����5���\�y����W���,�(�[�Ḥ�q����W[[)^N�Ov�²N�g�LX�����V�]ǜ����op4W��<�ަYv��n���И��P���R\��ŨK����v4�u����޻>�"��T�$�}u�Á@ٺu�ɻ:/w*ub���z���[��*u�	�췍�tH��ڂ�d�*�j�8%�7)8�\V�+�+m\,�qRʱ|�-�x��uB��<��{8�0��S�p��]K]U�����:����ՃQ2��;�ˁ��O $Zߺ��ɽ]%��T���k��8��>1�fԦ]4�X�I�uX�8[.�f�d��z�V���Nu^�obY2�'t�T���wX������0�]ǨF���-c�ǫ[y"�w]<�.�tլޡY&мp�XJU^������c��̨�ç�KzK�-1���Yk+6�xE���p�}�����+�5-�<S�ح���.�&�C�K<��ԇ�M��%v��}�cgX����KW9�q�o ,)�X����<�~))��]�����|(�t8�ƫQ�5�Y�flT�_o7��iE���Iz\2��WL;�.����+O��]�b5�-r�ov�_>�|�efJp�q�f����J	���Fjg�';S���un���=ktrǹ uF5B��I��h���W_4�%�@��ѵu�n9�X�Ԭ �WF�mXc
Ҷ�m[�����wn�x�')����-Q������̽G����7��W.
Q�cNk�6Λ��*�e�E�w�����1����QGV��s	[�^���8iֽ<�PUG4Ҭ����`�>�.�����&T46ͫ��BPŇ^�&��j�?��ck�������y�"�<w�y�>]]���A]N]�s�Y<t��Ȼ�9"�U�ƥh�U]�@�E��������JqE�K��K�Z5�{>5�b�bN^�@ԣ]]��;
�g��k��g�Ӹ��f��A,�^���;:+Ȕ��sl�^_;�M&�J'%�*�Rٍ�i�2r�LBf��y�WAW2�\o��e#y�ҽ��j��&��vwo>��צ�����u�uT#o���1V3̺H纵����H��s��u����K}\�L�lL�a�Փ�u�v4%\DD�U��Y�0��A�C�#Է�9HJ0;:�=�ͮ�1���H��}�W\�+3��ݘh��&���F��g"�f[J�#�ut��Ct��Vg!�,˪F�տ�T�O��-"�&��dwy��ٍwZ�ǖ& �_.�p�M,����Ir->wjK���jֵeb4��	X=]���o�@"�/��f���t25);�}��њLe�F9ܜ`��Z��<P�+x쫬7}1=�ͺO>��sDH4��lm2���������6ã�{C�8#f�$F+ȧM�s�;[�CV�e�v���ö)�[�u$�N�Y��+r���]N��λeY٣m���]�mә�_su���˽#Jz�/B��"VvY�r���;�޽���%M뽙��|���a��t�h�R�)jʵ�R�R�� i��̏�f�[�H�GT4x�fY-�ڥ՛PT�����-f])ح��l�(&��t�Ձ���)�Z㩔��k6w!�4�5qG��S{QWًrv�V��*h�,l�WK��jF�#�-�0�nf�	eF�fS��M��X:ܹN��gT�'`��؎R(�J��/X�Ǘ
���j�h�W7��N���A]������ni������Z��nɘs��$��גE.�^�-p�-cX9[D�>�T-1Q����:��zG��V�;ǏV�;��Y���o}6�R��H����{���0�!j(��7|�^���`�#{������W�=[ֵ�v@>GK+Va��,0�<��Ud&�jW�6�3K�PT�:��P�;n�.��2���&]�|5�zE=�]�+.�����@���]$�/.R}�KNg��*7t2�ڥ�ݑ�w^U��F��X��2��'+�Q�|m�S���%S廔�ɔY�j�X��7t��fM�;��Z|�u�V�l��r�b�V�.��l��F֤�����T֥��Cr��``VRj�)�sYv����xo�\�m`-J��Q՛��c�#�f	�\��q�*��b��W@>_wji�L:i�[��[R�@�,��*�n�p,ܻ0�8i"�%��G֙�nm\���٘��]Ѝ1edb_2���vzT�&��Z��s� S�Pp��N�a��.Q�Ԡu��.4���B�/�����E���w�%hX��᫻|�J�;1���B��*Rx���s�����/�Q;rS�M_;��4��yK�SCe_X'{.�or�*�%�]b�S�A��#4b�i_�b!/C.��r���:�]\7�{cW���t�J�/Z�d�oBn�`��ݝ��sa>���=�zM03R���z1���9��.��\��ߋ����qү�D�ۦyʺ�[:��c�5�?U�P,֣�]e�5���{��9���}ڐ�C+`{u����mm�@�g�%�W+%�o��U}�@�=���v�o�<�pv�W�m)�`jh�G\JJ	$� "I)($�  � �$���L �D�X+��M�&��
u.Z��m�o��wuI$�����ɞ���| ��v>ѭ��\�]�q�&����wv�!0O���A�Cux�=��S�9��q��WA�H�N�5�;ˬ�Ϝ}YmM�V����#��u!8�Q�Q�R)" )m�� iEb$�I$�I$�I$��'�~��c��-�~�=�*��$Z�X@ ��� u&C*����M�Lf3ٟT�}�P���q����KV`���ճ���`W��%�����i�4]����	z±5y�zU�f�5�U�z%zdi�Yy��߲��r�P��w�z�Gh!��V(���yXZyn�Ĕ���csC�'��2,mcaR<�&��e1�*-s�{s8��d����Gy�&͠��]�Sv�Ah�kQN��9 9]�#�7�jV�e��.�]���1=W�)�e�_>� �r^h�ԥfNtz��й�
�
�}��N��F!h���+����v���l���pT9�L��}<��ӗ2c��\�&�����a�٩�U�0�7��z���o���L�b�h���8��ƍ1.(���#�L���Y�	��Ȋǥ݇}XQau��KUD�ej}����
���W{9�����+�;�9#���B��v�,y[b��>TfMB�FyR0��̤K�s1�Њ�t��r�%�Ȳ��6Gk��|k/3�Ncp�i��׏�"��}����]g��:Z�6�2��Y��y���-���K$U�ơ��Tx�DoF��f��&�V=�(ӛܖk�H+3#�D�5
�u�\f��3d���fv�(2L����MV�Y.�P*&��Zg�ܖ����%�ͪ@
��:�K�4��S�[8A�rtm�y۹F�Uɮ�&�ڛ��*"�L�c�+;1����L�7l�P�	eWKk!��7,�am�k���R���Z����]{��Ⱥ�w�L�ev��(��P��(ʢ�:����J�Ӽ�x�JVV��w{K�k��E����ͫY�3�=��)�^�7��\uۉ���7̗�x�ᕳHG���ړ����h�k#/c�u��mC]��=2��Lv�'%޴u����
ǚ�'�m��YX���V�����D��w��X�t�$5}z7	�����K+��٤�}m��鳚���s�N��+�ثpj��3[��1mU�yN��\lLk�w�D�]8�����nG\5`ɛ�#����7��[�aH.��n����Tn��\K�0Չ�>0�w+lPH�5�N��-I
��p罏B�Gqۛ����r�4Բ
R��3��m�8���8�X��d-6\*U�b���[.��{��)𖛃
VjRU�Z�\i��0�L��4i�7��U�c��^N/�e�PuqB��UP	u3�F�û�4�V��ˍ8��O�W��6��i��#�S����S����u6�UP�W2�I��[�ͭ�Quo������G�T�o����7r�28QO*�*zt�)��3�.#2�mL�a��]����3~MV�+yn%c�rŹ�I���:�}%��PA�z��A9ղj�ZZ0T�q�*���z ��g��)El��hmc/��^��,�o���Lcj��sm+5�W����6�3*�]��
��	5�X�9����.��ѽ���I)�2�B�+�a֜�Ҫ�;X!t�A��˻�I��biLs��f�P
�olٱ�SL���1%\�-�*���V�d��FP�}�X�V���$�� �w�Vm�G���q���u���]X�*�I�+��'˵N������[���6lbT3#�L"QO�����ț�-&V�TH�,�s�b�qo�Ѹ���it����,y�E*ǂ�����]�Q-���Kz�����X�Վ�aKN�ƍoi���iKȳ$�2�飮�.9�"���2��oy��M��WU��y٧ ��"�27y��.�g��FS�u��W�;]����+���*�v���3{���T[���5�-��ˏV11{_e4�)��p�G�;«W����"� �@���)���F�����ob5;d��t�5o;�.����=S��5֫T�ֽ�J���f��m�7*�m����ީ�)F��f�����X>�F��e^[R�L=���g$��w\�Tu���i:�6�lu�
TulIw�ؔ�S��Z�D��V[�k����m��!�u�{Y�_m;����6��"�Dv����l�� � s+�lr�N��n!''Z����N-&0j���(m�'o<��;:�λ������r�,-j�;��ʓ�r����S�U!iY�����1i��u��d���nV)���afdN�gW*���b=H��\;%b3t[��F U��K2�X�J�Э�<h�.eǹ�
��)
�"���(�
h���ռ�N�cV(#�'4�c�ج����*�_4�4�胅���!"��hmi�)�˷Qg��T'K.����PV���P�伥ӵbn9R�-�N���q��d꩷�6�NBknH��7)^ҙz��.
�Sq�@�+��X�����!֭���zj���e>��W��W�(ۨj��R��N2�<�LJז-�GJl�?gL.��N���=u�	T����'\{l��sws��)}U����N�Ӕv)��i��ԩ�ΝT�L�JW����U����Yʺ�Ǥ��lE���|����9;[����vucT��h��0�3s�n4�|Y��y�n���9�D�9�'_�ַ�Nԕ����b��T���82�@C:G�Y�3�l�ޜՅ6]�Iaj�����dq��A���	vޱd���Xɷ}k���p\�I�8�b�r��X��l��"��7%Iu�����8GZ�;p�O�9ub�$��S��Wn�ښ�V"�S���+r��2�����:���x=v_*`�wuّ4�a����cܫ{�i(���K%���^�[��D�Z��)�}�'�R�)^fk�%�����ֵZYf���y4Wwf�Mi]�\),�1*}%��J�rl|`�}�u�����!<��w#�
�3��oV�Zw1�e�W*}ʃ�x�>��gq�fP��S;0uz`�]��Gb�Κ(G8mX6��=�ݮjM�3�=�\z��vЪ��-e]v��%]q���/��!�P)r�=9�V��p:f=��y�%��%J*w�����˽ə]r���jipnF�O�K��w��uZ��In��c���3�.��W���{��:f��k3Cn�̚���W+��fgŝwɒ����c�N�[��'C�T؞��]�J�|Gl�%�u��p��Zͥcw���A3cy]���,�8���b[j�p��)��n���d�o6ގ�uW���X���cX�V3�]Їm�ƪ�\h��=jZ�;n��箮�m�ؗ̖/����JҔt��$+{U�}o:TP��=9�J2�l�T��k�Ґ��N1�l�H:�����;]��xfb�"Z�U�d>\xK.�]����I<<������kU�0i�G ,�p;b�V��ԩI�m>7{�/�,���ۚ��U�ҸÆ��-t�EMqw�gP��qd8lH��7��Fo`���ofe��vEN<���X	�l��7`��8l��ɌЍn�O-�{��뛫���#x����+J^�z��u����A��3��n!�I�FDLy�y���˼?:�I$�I$�Wyu�cvn�'&�uQ�(i׎JI+����<7v�Q�ʤJ���5D�X��T]q�6�l-��e����]�9$�X��q�b�+���sWy�FĒ����J��S��{o�k3A�.�ߎBe8�pUmqĴ�p�4v�i'i]�+cu��#;6���۶q�������Ӥ��DCcX��2��G��Oj �Z9䁲�S�LM�z7$��Lv)���bSZ��B��&!w"�6�'8*��Ѷ9������9,S;��W�=�l�;cۻ!(m����b��w2��:�5�y4�SI1;wֽ�V�>��HX�u	d6�͖f-
�����&�ۅ��J��F�DkU����]�&+�	�5�u�5�q3����S�e������7�G�ݙ�A
I!K�'5���% Q�s>&� �� ,[O��d�$R(��f
E`(Abőa���AdH
aFV�YY��Ȥ8�I�%T����PP�+ ��((�§V�������bL"�eDjOY*DpZ[��"��1H��B,*Ko����Y�H)R^G���q��/��>j���/!�L��)�x!�$;|7�E��Fp G�ou+���A��N�����$�<"��`����̮c__�<�s��u`y��ѧ͋۠{+�idB4���T	\Ϫ��ꋝ ���cA�2E⌒���P�Th�X����6�$-"���Z}��P0�$䃚r�]�~�LWT�I"��
�\��Ǉw��P�9��h�a�*Αɮ�3�πqI�r���r�"�h��k�r��c��~3t8V��r��Ҏ�Fkw˰���rݷ:�o0>��	ȰrAL�\Z�d�$��(F�ݡfN��;�B X�:��Q|���B� _g���ɧ���#m�a!�T���t�X"�N���jh^�n�6���,L���ܴ�s���zV�{����Dgz��V��ND�o�mi����y�s���ݾ�,�[^S*|o�ʡ��:_J�<��f2'eu[�|S�F��Qx�cj�J*�GU��z�9r��8$�;�ب}Pf��;j��}4[���Y92@p
&gw�1�z�uצ�s^b��CZt�uꦯ����>+/z]��F��7I��/e�\��Hbf^f���{gW7��j���[y(���N6���t��=�j���7A}OP���)��s�+-�R��Vg��u��!b0�3$��/�׃��~Dgp�~ *�Ε7�б�ϊk�]^��av1i� �sg�|��A����P�9��1�ّM�:�r��-�7ņl�C'�b�]>�� ����R��/FTC�#w�;�]��MH�e%�V{�n�Fb�HŇ��c�)�V����| o{�S��_�@�U�c`ir�zt��~OT�x��bd�V.,�t�Eb���^���tϞP�d��'>�Rn�-80I:hZ�ӓG^dƠ�5+��y�azy��2�:ޛ�kB���Ǔq/Y3W�y\�����1{�E��F
���y���V ;́oa�����>�`����!P6��7{@�h����:���^�uQ:ON�z;wUO�Bm�#:��������M���Yx��G���t^���X��
q�d^]�mmuӼ\�Z;�!Ƞq�#�&���`(n�����^�H/2t�=�)x���|����Q +r눬�Y��׸C��a'+����{SF��+��?ģ��|��Z;�k�Nu5��oh�sk�O#�]�3ݨ�aY��+_P�0���]����E`�-�*^	 �,��£.��ϝ��@ưy��@b�7�QF����SQ�s7�Z�[�5���Z�#3��� �XTIa��ڳ��^��<������t�)�l�X_�4ϕ�u���1R	>~��e�<׍vO\E������]�T��׬tE¬t��Wo����%Ϋ�Y�T���&�>1i>qGBJ�2f_[�|�F�Ͻ깰��5㺞����M��5yyIB&���ܛۤ�jմ�R3]>O76�F��ڭ�Ƒd�i�0�~��1P��5}��^.RX���pW�Nl����g��G��Ȼ��tۿ��WO#��8�&>^+���`��U�i���܍3Z���l��n�sz�b�[9�68��\e$:K*��:ؽc@�5�],��J)�X��y���kH�����q���P^Cd�4����ʘ�[J��/�ƕ�K�g<�ߵ.)V�DIǎ�j����]��>W��"�	��ԗ�7[/2:w�`
���+����)����R�M�I��b��[2ɤ�[�J�:����L��9��M��+���S%Z{}v�`��vĪ3$ޕp��������#��`z))�{q��ܫ�vJ)��t��8���oPZ�Q�d^zf
Ku��}�Tұ&�sA!�	�6���<8�z�@�|�g�3���ǳ�����|�;UQ���7u��#�h�m��nU@0�A&��F��Y�əJ�|��[~>t0N>���}�����U�	;T� �!��D��[���*���z誤�!�W�س�O��/'��1y�Y�E��yvX����F|"�.���TCưV��r>��6��2�]�^�2�.���(y`�훻�c"(�Y[������κ\���E�4x�c��C��π[٠N(wf��o&�}u���[�^�_;��fk9�Zp������X��H$�Юd9���E�ۊ#2��'�cYV��5�L��"�����و:����Ժ�(7�s��%��&%�+�\a��^z���1F�3j�����TX��ub�Ů��`,v�ժl\eP�1eП75�h��+�<Y�f��4�}W�L���xB�|��ߛ��X�hi�ίhܾ�f�8��q�x���Ӝ��{�8lOP{Ӭ�QF4�m]m>�Yj\+�������Qp�O��"8u_3ِ�1�f�!!'���Id�/�7��vU��UG0�4oǍ��n ���ƹ��s8-=������gz�-�'��˪ׄH-�[�C�w̦��Z0-������XUл6o��'��S+��<v�j+��-�L��-��2�@�&��,V�����s�״o�Q��5�%�#83E<���>.?����ΩyP�j����X�i�M�Lc�o^@7�+���@dC4�j�ι	l��6=�}�����
��)^{@�;�5�|��p{��7�-�'&躽�n�븢��#v �Y�:�wg�k%�n��^�.�Mq�º
��@ǻ�*�.�7]6m�Q���:�4� �0Nv��FLM����'o��wX�F81�q=]���ώ�^�fO2��AJM�����������,#R���UQ�2�{�J�#)�B9����9���B՜���"�e��+k�����W9�?Μ���!����܃I�ޝ�`�6Cu�����G���;&��H6A�z���Oy��������gU!:�f�yDm����S��;g��T��뭺���:�G��n�N�Te�M��S�Z���._B�'���	.h<�\��vM��N��enK����bǗK��r��R%J��[n�n�c*��rx�{��N�%5Gxf�,�Q;��06tF�.rI�{�]2�����-�rs��W���]��s�΄���nे[.,5skQ/���l����8:�� ����̦���b�F-��g4�>�(=���[�5н�X��|���\��gy�F���єo��Y�{��ޕ���f��]$fgs?�U�WR���C�{����=�a�_-I$�I$�J�NB��̺[���
Ô�w\B�o(�B��M���5)��#
��,[�Kb�˗M��H�����Q�"�VCW�5YI]`$匸GX$�̉c@Z��Ya����H^^;�h��yf���]���ₔ���j<t��-��P��pT�|[e+�l�L%�4m�ʠ�I��m4�?���A��5��(��2��"�ԔNV(�TJV��p�̯�'�"�j�/�h�N�Tn��7�T��q���v�2�Y����ݡR�P �Bۻm���%F��i���7c��8Ѷ�X�	����60��1���Tv1��h�r�$�z�z���vF�w�#�G=������|��T���T��T��SS���\YUq�L2�jV�T��TQ@Y+EF[*C�+��͔Q�~k2��)2�&�0���_1�a��0e�J�\1zؠ(j��L\`��	�¸Jf�*�
8�UU1E�Y"(�)*At�Re1�,�K0�qE�V(`j"�uk�C��P�
a�²6 ��1�g60Ԉ�s��d�=��r�<�}�5��v�Œ`ܚ��#^�)���x�ft�4j�u���EVx�]����[̛�3lV����(�ι�d�-�z��kq����vk�|8_��]��?Q�de�2��v����~f)H����a�w���g�-��_��9���� ���t2~?ǥ��?T�Z�:���ֽ��v�K&wY|~�Y?��~�B/o��-\����2]�_lTm�ɬ|a_�^���b���P�a)�ߤ�b0�
:���w��i��8�#���ݥ�;çu*�aeL�m��������[�,q�Y�s�U��ᓱ��o�&��w)t��g3u��ߦӞ'�����k���v.�+ٚ�x��;���Y'h^q��ddv�w�t�g�&}W�Ʋ1���g�Y������{/.�~�>��O`�����|3�9��w�u"�?z�*<��<�hl��Fn�
�����������ŭ��؃�G,�+��9��ǟ%����A�+��.K�V�*�ut沢�>}��@=Lcc��^o�:�3��B�Z���H��{�1)?|�����l}U��؜�7�:�M;Ԓ�=\��q��v�A��$	���Nκ��tR��{h� �ms�}���!��T�H�ȱ"���_CavT_V���bW�*p(մ�t�H�E��:*�����������^�nD?�φEmS���1����ֵ��Su�W�u떗�ܿn@5|9\�\�v�v3X���g� ���h��N�U�V�1�)��C��o��xJ�s��y�y}�h�q~���jX�qR��D�V-��P��-�:ISs�n��y3r�{C����7ԤH��=�UxM�>��j?Hg��G����b����~���Q�E�U=�;BXS+rVl#��h�-���C�ϴm�X.d^���^Sj�.�;3�D���6� ��z���%���BpHĻ= �.�㗻����䇃  o<׾�?��)}I����Q`Uc�[���[�+\ߙխj~^�����G{�����R�z� �x:��m�����gO7�����@��o�����9
�8�:��E$<d���m���u �!�i�Yā�i�j��8�~����ߵ���:�&0Ρ8��8��dXOXBd�o��	&Y0������L>L{���}�<d p�'�>d3�@�{L2M��6�(��&�'�2{�q���ϐ�����uu��y��ϡ>`}�=d0j�E:�u��'Y���u�q`M0�$���2c �=�N�{�mxHv��>Hi'��0���z��'X��� hfP:ȡ��N�`i���]�}߳�s�L�`zn�i>�C�l���z��<��OSl���dYr�u��l������;��:�/LT��'cl��n�f\�����[�-�]sHkW/������v�I���g>y�k^���Aw>���Ad'<����2I�&��񒚤bg��&�0�3�@�N�4�8�aY%f=��@��{�c��_3�5���=��N���8��=BVe�a'��<��@��bH}�'�2x��!��	�OY��8{��q���$:�l8�|n�08��v��ؚB`x��d2�1|Đ�����i:�c	���}�s���e�E5��>HB�l���NY&Y���i�g�HQ���$�$���IĚ��s|~����^�2|�`{�I�'�CLY�|����!�L�5��q�He�������=�޷��2C�Y�2,�o�'�3a:��϶�gt=Bq�b��!��Xc�OX�Ѭoߵ���&Xa��%1d�d���$19C��!�>O!�/�!�!Ć�py׷]��o^�m0�$<N04�2�|���cx�!����?gm����c�C�&���������[�\�a�����C���2�'�x�I'��Hu�?XM�3�N0$���w�y�wϵ���2�<gۤ��qR@�!P�Y�q���I�0��6�[$?O����w�����/�@��~ݬ���R�ڝU����|�v���\QjT+��GS=]�����9��N=�2�U�o�> }� 1���w���4�m�f�����I��a���I�Y�y�P�@�'C0�o�<紾}���{�d�,2C���,�(OY��'�VT����X`q���P:�eB{�y��{�{�k�νǶY<I�P�ˌ�&��d��c�AC�=��ɍs��T�z�8��"�p��7߸@�=Ւq�Ԝd� d�9�ْ��$8���6��&�d���>��\�X�y�=
Ȳ����!�l�z�4��'&��$.>ć�d���e'�}�}�y�y�9����q<dyC��'u&����8�L��|ɭY�I�b�������c����>�'X�HL���@�d9L�6��>I:�4����2y����$5�O_m ٫!Ă�BM$0��Ru���i6ɔ��a}Ϸ�{������}�:�I2���I3�Hy>�q�`c>��@������ |�`z�ެ�,����n���Ϸ���w�d�$�&�OXC����u �I�C��Cl3�x�����]����s?W�s7]N�Y�U&�˂��7ltql"^�~���d���f:�K|�C3)�lZ�|�y��]��3��n����v�|���E��|���8o�k��fY��@��;�m�m<L0�@�&O��$�&��~����i��N��}Ϲ}ƹ$6��Bz��N��$�a�i!~��d�I��Hm� ��6��������{���<@�C���S)��j�B2m�Rw� a�<�Y���	<dY2������i���+�]��k�y���3�T	��`|yg'��y�~`=d:�!����d�hq�:�7s��y��{��Y8�z a�Ű�`gVN ��e�`T!��T2O�C��!�?Rv����fgY�5��m����2�VM�<d��Ha�I�>�u�<CԬ���P:����[�^���{
�l����t�a4�:��&�<Œ�Bm!�'�X
|��}}d9x�]�\_~�[���C�a�@�j�m�a����C8�B��qe'���q�a���=����n��L}�{����Ğ�>ϸ$Rz�� ��=B���L�P�}d��8ɤ��a&�!�����_5�w���a>�!�>RM�>�z�����YC��P�v�'���T����P��p,���M�?nQ|F��_~oƥ��37:2&�;bY���Ө/�w9���Rg�v��-��y�g��;��^y�����$ C�!>���@�ϗ�aC���'|�� �u�{p%�4�n���Ίvoe#G]W�Ƶ�S8-��Ӯ�ٓ�����Zqh���z�_���]+�Uw������K��r�y����
�"S�]���ԣ�t+V����\^ބF9i-�+z�)1s֌>�	�Wu��E�aJ4�t�b�]��S�鹖�zz�+�%2���̊�n���)��.9'�8�W�('^��#�[�c�7�ʧc���JD��[��/zZ�f�w�5�OzI'x�c��^(S����nJ���;Ph/�m���� _���&""#�`  �s�5��q����1�cw��ͬL[�c��m�sc��G!#��C&o�F3l����Ĥ���ʋ�;��*���P=�p�=78R��8Q��Z-oq�m_�����!���Nxb�W+z���Z���9 ���Ы+��h�j�s�7ܽU�j{]��`��ov�:��煥�`��ύ��xF{v���.�����.�v��E���U��>���ݷ]~n�c�v�'���ҿ~�0����f7�/�p��l��2�z�����*�E���ʴDe�[�R�뙍qL��wj>6]����9���7��� !$� �@���@����E� , �@YQQAd��y�ϯ3�9����ɽ����	]�->M��Te��뎪���m�h��2���K�þ���WR,����K���Mcy�˪|tv��8�=g���߽��`�Px$��>�v��8��Тu_�*,��� @Y��3��^��ЮoQ��Su�Y�$x����}E˶#z]q�����To�f!Q
�E���Hy�M�y��ܙ$�-mP�J�W
5o:��!Ok�����������*�^xR�����UP�-�'sm+�>a��r�9�|�3�٭}(u�U|U:l�V�+p]Ϸ��CG[qX�u�fh���^�/t��t��
��MN
�w�2���қy��R��t8r��un����T���iu��:e�܏lZ��{R�����4��,�tH�C���0���ޥ�F� rk�kbU*aQ���7��*��&T6�Ix!}�0M�h��Ql�[��_��L4��������0a<&���: �Mt��k�܌��;���	�l��h��(�v�G���)�9���;v�(��t۬.��k2����W{UUN�ǧ�p"^鏳i�gp��I{C�7@����ܞΜ��܀�s�t��?|���+9��I$�I$�I\R�Ɍ���F���+V]����ϭ�-�n�hQ��
��:��+2\�f"��x�Vl��Ȭ�qE/#���.�|��i�YQ*�re�1�J�-�)b��l��	NJ�|�x�8/fe	yT*���daU�4OΓ%@H�j�)Ad�T�[-ǙX��YW��p�� �1�#�����4�pK�T�B05b[r�f�ϝ�U0@Q��O0��૤k6I��[ͬ�D՜O&�	���P���c�o~W��][��=�v����������wY���D֑�i���$:ʹ�7��XM<SWu�<-*�ui��I�CUt���A$�wHE[eݶ��;��ut��
��������)���?-��j���d��8��w^c�d���J3���9� ��)
�I�R��SVf.1O(eRdA�cp�L3���^���E�q��V\�Ԟ	�f0+S�ŷ4˃4�.�fq���i��c6Q��p&&�&<˜�Uϗn�<���Y��,'��Շ7�`��Ln�dȒ����W�|�sB�m�5� Ç$��'jX&2*���SQt����h�r=�Dz!vi����8yP�x��X��Fro��KVi�]	[�V�����s9B�v!��ۮ7%����Ax^"XQ�!���V-A5
�h[D�/�鑋9XzWZm�w6��؋ئ;4"��/���;��`)o�*XFQUշ@�qN��f�+޾�x�u�<�AQzʪ�C|��j�x�M�mY��Ƕ��kP�k�;����=n@��0�i�v[Tb�au���O\�V��?{{ﲬ��>����1[l�3Q�-�a���tĦ�īX�9^�[]K'(A�	���[*w `q��p�P�����{��!�N_~V�?��gd�(Q 5O-��[��SN��F��"i�f�!^�����Ђ��uE\V��u��;Y�*�oyɋƁ9�h�� �9�A����c�@=D����( �KSK���WP�t-9&/<-�ݾ-��u�td�S�f��ڵ��8����"��N�zΡ�}Z*���K7{���K��i��F��C�L�q�9�d�V��X���ϭ��]���{IƳ�����Ol[�Z�����U�.*��z[����
xi����8�hUq��t�����
������ �o5|�3��l?�f���ZS�|WR�%����=1��zO���f�Mxh���9�Q���]�S�Ag=��g���Jo�*������~0�����}x�`B�Kt�[)���b�ʼ1Q1�	�h��"l�( �]�o)�R��D���MT1LAMf���T"�gcP�n���n������(ޕq�j���Zv�\ޔk�e1���E�z[it�S����#�B[�yw}�9k�������>m�Ӓ�C�/��?���E��	8�j��-ٙ�8.��f�Q��r�ΥZ��Z\�U}��Tu�!;f��,�.�`��YeNR�+j�oF����	^V���*����C��cYǫ��q��; ���G����m�y���̢�/�7���B�ްrzLK����rYP��M=>+շr{)��p���įS]ז�IÝ��p�; �>��u��L�W<�l����d��,U�7��/9��/��I��#5�2�zD*����A�uYd�';���j��0k���|�0�-m8Bf��]���K���<I�֠ݫ>o�\�q/w��ґ$9��t����\��:y����I {�y��{n��yhˏi�u��ʰxk������	��5(�׫��r�d��ީOk�8)9m0곔uf�y�uކ�5���Dׯ=��X��w�T�����~mt�E 1�xRǢ7�ݴFuaa���鳛�qp$���U��ѩ��g��.���q�tE��d�������^�H��=��~���(���i^����mB����}�+��ݬ
���U�(,�u����j��o�OuW���:��Nnsn����-�Joj]a�f�_L�9��50��zE�rʹ~�DDz(b<��ӆⷞl�`ϐ&(�p�48l+�\�N�¶ѳL�U�]��y=LWl��^�^�w��`K���V:,������<W�SdbAӠO'U������-�f:չ��"a�|"�����v�K:kt$��2KT;5gb*�P�@���즰��&�׌y���*>������Ɲ�#&�
쵲E�����o;&^�(�_J�/Nrƭ��o>j{�S�"-:˛}\�R��^���\�<Yt���م
�_>��X�5e@�JB՘lO=Ԯ��������َ �ڸ�M�z><"��K�͎d���g��b��`D��^��j���8^�X���S����Ǜ.L��IR
}�³c䨡�c�e��gwY��c$��s���3~�w��K@�lSt��(o��(ŅvR��^#}Y�T���)�]�
�`v@}X���]��$�W���%��O���c�Hzax��[N�W�^M�|\�� lcn4A$L�9��n�u�;ѩ��`�Yl��٧H�+��t�)$�p��G�}� �K�mJ[]Ǧ�bw���٧�$��ҌA������x7�i������_V�������k����7j'�v� >�]~���E���U�!�c*;\�( 0�=V�TU�ST����Y�RC�\�Kc������e[��n9�v��]SH��cλ��F�,p9��^��7��[�����x�����\o:����w_T�a�h���Z��`��OW�8u�s��a��'&�J�L�V�F�m$'�^ۥ���VZܸr��3[�E����	���,�۶���ޯuT��Br&�6I��ܾ�Dz��{RB��A���-t7{����s��������s�1Gk��#�;��Ȓ1M([s+1��{TNp�7a5^R�o���j�ڈXޞ�ǂ��$=Q�2��:��Ci*���2�L� ڋ�;wٛҷ�ĺ�9 Bu�c��N�oz�p�q�7]^��Ғ��Pe�������<��iS���y���i7�\˹���-T���b����X:�SҮ\rw��`��+y�Vb]��D��f���Nƫ�ƶ��X�E�����c�>�T��_�ʩ�B�E��m��
~ߔ��ZxU���].�U�*v�C��7��b�}&�]?}���v-l1?;��1ѽW�6Rw	��&4��p���і��\U3n�H�`�a�f����*�V2��}����oS�����t��Ω�G7A��?�t�?{�����h����XQ��rD�.�ⴸ�.'3�Ptg���9�6r٘ !���&��yC�o�v�獈�gط*ۿ^v<�s+�҉u|���M]u�+N�j���{���ޮ>q:��tT[q�������.�1�:`�����h`�{9U�WrR�J��ԯ�u<;��R.�|�8���M6���%WY���&��FwE�!�i�<zge�Y|-	�=�q{]J%W���s���UJ�;���r�i�UIC��F-�+������;� �^ST6��V7KD�����\�a
��a�v�f�͍"�`�%�L�RM�UG�*��YT�F]�{J�g"ͤ�`!
�viik��j˳�΄sp92��˕Z��[��ț�HWYX]��K���$g�Œ��N��W��������,N�8�Vea�Q�q���Cd���[
����ԉ��og<�Ms�T�����R�p5ydJ[���٫
ݝ�o�᦭j�%��R�ԥ��땺���ue��_)�wd[p��>YU�F�Ռj9%��1T�I$�I%���0�b�t�v�J��uT���Q�a]��1�f]G	&g��ʣK&�U��f't��^[�Xxꋻ������%�iY��WN�Y.
�3F�̊�c��(�2f'�꬚k7qմ�8!�We��%YM}n��3%T�db���iPJ�fʲ�8qg�%�U�l�p���r�9PaD�HYǔ�,�_O�"/rhY4ـ�.�צۺ��m�*�6S�8��޼�"�,�3ټD�˗d��e�S�г���GS���j�s�8�y���F�bd�
:�(SSQS3�ELE
���s=��6��h,��i����ͳ�`���e6��0\%\R����%E+����n
��QE�mۅqj��t�0�UF#�8�2���VeK�`�Rx�
b����f�-��D�)F\�[�a��B�|Ur�iP+*�m����rs=���B�B��ΔrZ�:n�I˝|Ndu��=���#�����S�
�{���kT�) �|u0�g�MkwVG5Q��X7�Xy`�85E8^-��z��v�ĥ�w�霮�VW�
�ߥS[9�dr΄QZ�2�F�6���l#&��Cl�Y�۸�,a��7,V�U�]Z��rC%k���i�i��O�f{k_���#�
����a�5u43�Se��hF���-�$�_�=�2�ZQ���H�{F����3�q�l�u:,V�{s3Z�N�7�d�ϡ���%k�,��1���x��Y"��z�f��ƃ�:)<]-�p�� jV�ep����6im2���V:����N(�5(����DlQ�F�l���_����܁k��gp"��r^mC��IH�)UǦ�.��	��Oyc\�=vwT�ʮ��I�-�\,*�p�&��r�_����������f��qf�� ���2\����ۻUl�Y��j�\���YBR�����(q3S��%��5�7�k��(����9�TM[=]��S���b�_ly�y�ԥ���Њ70J��i��J��<9���.��J�<������R��'�˲���X��1�=G��z"��<�Q��Sxֺ���<kv�"�s�Y�����]p��NZ5%7���m�5hZC$zJ���\���`�^���}}o}�42�H;��Ȏ��2�r�m�Q���pq*�ac"�q,�/q���9�Q�dd+Bk�k�|-K�x)"��%�x�Yr����]aK|��>�Q�&_���t�no���]�����2M:.���ۛ�%Tƻ[��5}ݞ}�����yZ��wYc\wJ���#�p�2ޅ�p��as|�9���8�9�t��u���R��ͼٱus�yP��b�O�D{���g�W����㧴d[ͽ�p=�
�1���W|Z���V�T.�y��e&-:��@�41%��"��n��j�5у+:l�m�O-��!�V�5o�p �����2��.��%�du�Et�zI�.�Ewi���[�`���㨮�{ԍ
(bO}kOc5x���;�3-)M2�33�m����H;�F�.��qwe#���%Zl��ҳ�V�>��k��N�/�=����&�U��by�OeM��d�i�֪�e�&��.�ioY��4�ܗw�t�̱s�lթ<y�M<�ވ�%0���Ҙ
�dLPۋ��E�X���0���a���mۍ��rVo��ւ�5�T���+�0�78�����Hٜ�*j`��wEe$~WY���z��1�1?y�l��k���v�+�Ô���9
�`k�>���מR�C�O9O^�^S�o{�|��vW��|p��L�W;=3�q3�%C�yK觷�2Ns�,,�j�����Q��UOL�6�����N=����qh�� ��l�^�c^��ָ��?{���9a��\��u��5Y�����f�d{Er�8ߔ9��񃐗����(ǲq���u��#Sێ�ڪ�^�\�z^L���]܍���7�sx�cBV��/f^Z<&.6�_R�R�]5
�[�Tc��2Y{Ok;��/�]VIZs�w'-R1��;�űW�c]߀��e{�F��N��堨��i��>5�PhU~�������+�m��٣Ǣ	�'H
��ϼ�4E�xE�7C��v�37q%�1�b���� �­�+���Ǎ>�J�ĳc�"�n|�UO
w�٫Pb2d�a���Y��zN<{�Qx�{ e��"����0�̭��//On�8av����G��F\�}��b�U�������x}�k���Xo�_%�y!��",������>M:v:O^8_<�\{���N:������YOw6g�DY��G���)�~�鸚�0���1*��"�L(qJ$H�0�������4�!əe���<��m`A^4��#U����ƈRr�U-��V^����U'%����u.������M�l��7hS��=��u���D�7�a�ӳ�i�H�TY�$�Nv���G[a�1�}K���O -Q��ĕ^�[�mnK�����77����)Y�p�X�5gN�n�M{��U�쫱�|�����1GI5�4z����Dɒ�y�,�B�C�~�)*g����(T��k�+�������!�Y��#g�HJgƶQ�~��]y���i}r������_Q�dC�g��3��J?$��
�1HJ�0���z�F�kN�eʐS��^'�l��)!vp���Ŕk�v��9m�R�������a�QH�T�>�:�^v<�̦f����6� 	yrr�/k���7�u�[+�_+�u��m��&�PK�D�x L˛�l����=u"~�U�f�\���f�S>+��3��0�4��Ŝ4Rnr�������#�Vx�k�z�f��^TaEs
}����r�L�f!�NyK�;��˲��g�R�)��Z���$�R�/.�s�s�Mu�=�՛WC�����0mӾͪ�y�ު�M��A�(���d���*��L)Sp��S2q�� ���=��7ʌhi�<<��(V.=��>�F{|�̾�"�?;��_(B�f߮i�I��3܆U�ٺ���g���LGu���2�񃁝�F��j��S����G�X�A�QG_V?��2j�>"��e���]o����Hcy��q����v�e[�����lXo�-�������b����Z��>�w�8���սh����ZS��Ю>�V�H� ��Z�?1�a����6fjY5I=�^�caz�|)�z�m]z�ծ+]��t�b�Ӌ���Z~�6_[���@ڼΑ0��MsR����R��
�$���q�M��r���ŝ���(� ��x����2!GN2��o��v�Y[m����W��u(K�S71r$[��O��8k��M?�k��M��D�_o-8t�mz��iJMz��X�о�ǆ�(�/yr��y�1%�8Qׁ�J�ڭ��{���1���el��B��r1D��u�~�",Æ�CH��NHx�{;��.x5���4�4�=� A%2�V�]n�vƙ�b��v\�:��dU\��B/�L�v��O�(���1����*���A㸘��s¨�U��R�������UȜݳ*i�G����4o��F1L9��^Aj��O��A��{U��3=%->դ��b���:����f���GqB��[U왛�<%�����C�=�,�㜄�.Q�IlUǥ�&��߮��f��{K%Y����k�[�x�۬UH}���m���J0cVp��B����n�b]V����|Lc��օ������Ǜ�����v�m{z,>Մqqӣ'��!��Y�D��fL� ;x���r6��3��J���ְ�cÀψ�:�^Iۏ:7o�)�ij����_M,��\{�I���6��~�P��P;A|�S��큊�V�h��u��ZʩcjWZ���ѵ/UrT�5��:�5U�1X����9r��ͫN3��Ǚ�{����h���|�]����=���v
w&S�Z�U��iki]��`��y���p-E^��v�T��c"���z���{0����K���9�ho+K
IV��W�nήs�PպJ�n�d��]k��$m�A&�L�)�o�a��be� mΙC�ej�vxV��@��g*���iq��!�٧�(��Y�זj+�p��y����ػ����n�x�g�����S���;�-&�V���w]ٷ��،�ݭ���?�W�^�ԏn&�uJV+J��tgJچ��u��E|��*���p�;��E��4ؔ�V�����s�Rm�ѽ���+�Ћ���@2f�$�I$�I%�\���X������Q^�͑{�!�k
ܻI^��ՙ'ڮ�]�:N����픫U9\����ޮxOE�+Ə �ӆ��ޭ���=N�\kb� ��.�1��0��"�V��4��xow`�@�s�k;k���i�r��2��v�
�M���qiy�];��.��(�[�Z��L����Ѯ�r���������I���w�Kr݌��0�e�[q��s``U!/��^Y���c�{�f�t�b��ǵ��Ī�7^we��]���ڕ�mh��;T�x���ޚ{�!�8���i[�m&K�nfv6��Gۉ��tQ7��ʔ�:w�]xB��*����-�"��鳥��]
�]�>���e�Zۚ-�*<�L=L.EJ����4RƳ�%TM�0Ԍ\[EA���y��LZ(��DUEU���DM�#��I��1�8�[���T6�Z��(��(i1�b)mT|�V�ZUm�����Q*&��1up�QDE@�����0�m��)Q-
#KU���X�i�aU���e�
(��Q�!c�U��)�U�,
�J�����k��zɨ�RڱY�Fu�(ިU�� ���	w7Cߎ�o�v��h_%��$a�Z�Þ�@������fm��4p�@���!ŏk��cYCN|�ެ��=9]��ύrI
8t��)�(�6},y1��k����S�����q����7��4�L�2����ɳy���_N�K�I�� ��<����^�o�t��7�"C�	�ԇ!��}�^.=�Q��sF.̅	�Y�:��ϹxٟTc�0���'(Q
��ذ�y�8�k6l颌����^9k����*@_d�[p�>�N�)�����!�^/��V{�<W���7.��!Ś=�B��H�w��15�r�5��n}�dKa�&����v�Vf�!MVUwv?s�Qy&RL��H _��	��)d�x�Yذ�2�p-��=D���Z\_�FQP�|4b���{�3��ڹ�sC�[a�#Sb�b}�{ۤ�
�	~#���g��w���n��6�!����,_�vW0�خ�E��(���>�13�,�%s�a�y��>��B}Q�&��6$Xs���}8��͈׼w$��p�v��ȝ4~����2׎�B-��oN�����_mYfǦ��՗�x|E4b�)x�+r�����v�D3�O}�|cZz4ş��U~s�N����&Og���M.�`�8��BZK��CK�a�&n��?]z�&�Ӷ���t��G��D�:|F�ǈ�yG��OV߰:<Yη�x�`�p�TFy}׌v]�]u���t�2]1��*b�j_+��UN;qs(l�x����`����4d�2�x]��{�w-Q|�]3]�9LTq��&����/�mA�uJ5A���9�Qʌ;o��Tx�,=�so��:�<Y����d_��Íٛn]j��W��'>�]t�s���K�?U��	��~zGUK�������UQ;��=�����tt��颈Ɇ�2곐X��79s�d��9.��UŊޢ*�=&\*�q�r�v_��7�㠊#�5F���Xw�L�Wʔh��P�Iݢ����	�*ٹ�5�NV���+�8�skԺ�1�Ɨ���٦�����dQ'�x�A��X|Z�6��윾,+v�[�����3�yr�H���s���q��y��
������8Y����g1�����;�	�/2z<�S�u�0�J͢�S��wQ��vh���a��O�}Ƣ=[�ʎO���U��)݈�6���hK.��9m#���pN�!S��u��1���åǉ:p�C[8a�'��ox��u����4�r�^��}��N�x�Sn�z�b�0�䰣�L>�H�^�E��/.7��Lhl�V��D�Ǐ8k��P�A���L�<w5��zY|����@�X"���N?wP��qb�,Zg
#p��u����2u/�������DHxTB��9��)�A�n^�G�{T��L�/��������fΞ5{�ۺ�ݍw!�ń1��ըձ��C~֥zb��	��5��^U�ܫ��|�;��a?q�D7[�_�℡Vx�����H��%�:xD"o�Kux���V:��n"��J��9~x�ngE��n�]�N���ym�GƳ���
��m��\�c�׶h-m�(���ƥ��ޤA����?{y��.s�w�*�,#{�M��W�?�����w�4U����}4��b����5ꎟdƠ�fW�3��>^�j���j�헟���e��hw-�*a_2����X����&���yjR���~_U���;G���,1��^�g�sZ*�>�k�u��
\�]+�?l���Nf�S6�Ĵ����g�>:Xp:0�j�������a]���ܲ���]n� %ͪ|[@���8]�ݣ|�ٵ���J�q\GƼ��c�v!fR�B����u�zT�G�#�a��������6�l��G�*��S{���0�����_n$Q�!��r'�<�4,x��MDš�q�Z�t1_^�Z����E�Y0eUTs�'f�ܸ�h�E{xtItq=&��<�c�au��Iө���(�{ֱ.oY��`�Н������5�]ԥ�.hw����I�}�m��X	f�^Xz��H��%�ty��q�_��J�����.�x�"Ӆņ�l�I4���������o�G��-R�6����dn�i[y�bۛ$uV0��V{9JϹa5i��3Dw۹��6lA�]c�2�߫��M�Rg����� g��o�8�#9�F���?C(y���)�K�7�/�2�.�w���Z���}�4�s�����,R�>�\u�����SfD\�����KA����w����nXF�3"Ⳇ�yLZJv0��������G��5n������x�Wrë"�jr����ѽ�^�R\+��N�S�:Y��4Y����b4������-s�QU������rz�Y�3>ӆ�i���0͑�U��^m̜H��a�Wێs���^So���i��!��2ɩb�k�a��;�rf%W*�HK�/|)��ag����_��w6�4���妲UP�Dg��V���C뱷q�4��=/�(HU��}P���ܸ��;:<g��R�\�]߽״<p��=�țm~�b+7��cCN�3����W]�eТ(��
^|hC�xaD�7���%Q�d���\-��3nQ��U������gv��DI��9�x�gd��]�L�@��"��d��ݯ����_̽
��jpq5v�b�Q=�`��U��io�[�]�1�-��e�& �x9r[j�[w����zH��(Υ�-�D�*X7�¾����U��O|�=�d��~�9�s�4�~���:l�V7�?��=��&��yY���'����V(�7����%b�Vp�;��dċ�pb�=���u��Μ�&c@�^S0dtM	���4��}dy�X�!珋6Y<x��C9p!y��������_1����螑与<q����Y�f�W�p��n�Ε�8y�H�z��6F�\`�ğ>��5mo��@�~��Y䴢�
���e2Yz��*Ow�������w��"XՄq�V~Q"��i�L����S���&��/+!��o{�җ�C�t��WS�c����C��ה̱V�̐W�CU�v���";��$��Ɇ38樂�c���4���=N�n$]@��=�I~d�e������|��K�L�p;�T!�5G��Z?y-��͡I}�)鯏�W���^t�Ξ�<�w��7�F�].��t��\	��0���Hq��F{_!٥ח�H�P�G��r��K�"���	�Ի���.�c��y,ύB�M�0&-4	ڌW{L��Dl�P�h�n,���R��Ҳ���=^k_zv����>ǧՙ8�/���c8!�#
7��&�ѣ���d;�M4x��L��P��#l��t�Ƿ^�l"�1e��_5|i���Z�sï��󔋽�J�����D���2�jDW%�y r����	�w�n�hi�o�jѳ��:`4a��vS8rM���5n�8=�w�FC�͗ёٲ�f��.���/~�1�w��q��9��@k��.dV�g^]7���f�b�i�����\/�5
{P�g���֝�ϊ ���8w�pi0w��Dڟ�%�)�b\���gc�L^����~}U~���+����z�����~�q��X�𵒷����hw�?��b)�־�H���V.=>�N��>)����i�E�<�>4eGYS�u<+8U��/�&��I���t��4x�F
AOM6x�z��8p\���<s<�J"�V&3�eC���e�;Z���Vp��^w�n�}��v�:nvI��Q��LL��Iu|�5G�V�5.g�Zy�+���*Jd�*��)20�E.zհ�'����*y�*���2���{�$P�U��h�!�`�iuk��9Vv|�s���i;3E*�R��G���!v'm\u�vY]�j�y�!m����f���l�X�%L>*���1+KwIW������߲���mRM��f(�O���s��h΋kEɆ����[9�tu����\b���c5���Zo5��g�f�.�(�u1Ɲf�]�mH�V-�um���Y��vtw|-B}HT�OX}�.�
�t%�5P�����Y6*m�,�̱��y�{�B9�8I�)L��2�:@��m��7����N�;LI��ӝ%�G8�ʼrV�[���Ί��Y�wr�F�T�Z��v$nX������>��7ed�@�x@S&�.f�w2���gjƮ��	�&ap����^�s5\�5O���[��(B�y�RI$�I$�Y�7s#/8�9P0����y�+����z*�Y������kU25)#%����ŷ8��r��9�nށW�;ީ]ܮ:�n׷}�Ƥ��j.��,�z�17j
���2����O4����o����3�y�P�P'[ea�Õ�����q޺��L�:��m�Z���n�s��㈖��!G�ޅ˓ŋ��*C����{K\�-٧{�r�:F���Uۚ�Ա�2��uֹJ�v��P��1T�܋e�[�+]��V���|�r��͋�%�*d���M2�%.�z��1�]��ν�kVq�`��d|�f��ִ�p�շ�3�mKP�yhLUЂɒ�����j �c�;�j5��ü��s�w� ���^��x�ځy��u�A�o��n}}����H_p�s�NaM��֒���6vCJ.mDb0X�k�	���#Z*���9�0�@U�����h��`�����DLU��	Ĩ1g|œ	�`ÛTe�b�"b�DV(0DD^%UQQ�
ǩU|hx���U���Q{B���_�Q����2[H�QUQ���SL�f����PQ6�p�P�D�QX)V+�����OQ\�Db��n�(0wJ�(��c�מ����˳Zﯻ����|������UV1R�u�l#��I�~�&���Qdi���eu��VS�^�Zh�g�p��*TÑ3U��p�ځ"5�9g�.p�`�z����9�YG�[�a'#ǎ���k�Hf�/@�-�.��Y��G�҈�B�WH��N�J�K�d�rɞ�.	�l��yq㜸�ǑC��1�W��8��S��2ݐ� ���|�.�A����CI��Tŭ���j����?=4Q�@�;��I+�%nz�=�K5X�~Zr&g����`�Re�f��ȴ�Ν,������������d��U�m�p*㥟s���m�~���"Vq�329ְ��/W��UfGo;�zũ�T�zWyg$�n�H.�kr��;�hѥ�ՙ����#���ǔj�WQ;�?Wm�f���uJK#�-%��DB'�چ�V�a�5�v��vh����vc&�q�:�{�nr����)Ɏ���=!��f:c]y��[�	b����L��!�L�7/x�;>�O���hxц�4,�X�Q���(��ѝgw9�S�=qn�I���2*���l+J�b5��לH�q�<~��q~ɤY&�qx�|�������#���u��Ԫ����FcMQ�t)��˖纝!O���r��]h��3���鹋�2Y�*a(��]�3<��f�t�
\j��u0yi<��OE��E � Wl���U>�[bpG0�L{��|M�����C�72Y�U�OB���ZYS(�)�B�fND�(f�s5Zw]�����](�6٫�.I��Y����	$��m.x:=;;*]/K�[C2�vw,���wC 8�l���O��3 �?Ud��g����Q��
���6����q����n�JY-�+�93B��ͪ3
L讟VT	�t$-��Xz4���I�#�d��{А�q�NV�W�k�C��yY��N��:z���!ؑU�KuA��(��	�+��}���A�����)	�W+E���8�̧[9%n9ļH`��>,����1�a�kQ�qW���$物��?A�B</^(�oV��fu���1=4��h����$�n��E��U^J ��-F0�u�aOun��
��6��R���2��h6~�x�*��<�f�,n.8`�|}k�Ҳ�tf��B��FG���*���W�Z�<�.�32�[sl�u�*,��/���y�������8��=7���L��;:J�z���aM,`�T��4ؗ����o_�~���hDά�=4������p����t/�����!���f$S��k�B�t��UFD�$I�ώ� T_ԇ�f�o�*w]��h���#Myn���Zt��DratMn�y�Kj��
4{e�1qi�<D��tqζ(�UY�,f}o�����2���L��	��yŉ�q�R��ܳ�)�Ⱥd�ka��.?ny����F�It��u2Q��h�F��Oƌ�,�6"�>@��A�������S�����hѣ��4B�Þ����'+��S�6��N�*�#��ٝ���H�zuI��v�t쎑���Y��R�2� ó�Yf WfZ�6ۚ���j�Щ�Zx�{ѽ`�a�<�z�w:"Z��P��5KL(�,3U�	Q�]�|������J�܁0-��0���WMĎ�=�z͊��2��K�ya����maϏ,٧n=HM��o��:����d��ze=�x�y*a�.��,N����C��J���[7&M����2y����+ ��Q��v����wכ}1o��,
��}� h�����ځ,�Xs�f?C9���秴p�xYFC�OsQ+U�<u��Z��۪���3�^n>>hk��������x�Ee��S��y����y�ӧ�=�$8�bF��b�o{*�l���G��܁�8�as���c"%;ut�jc86{Z�=n*sb_ml��0���+{�!1�[y0�����זx�W����L���[��E�F�Y@���J�� �i�B����⠞�1��M�!�;���k����A�\L)��/"�tW�-ّ�*�#<���#fVn�fܫ��HFO�t�8}������YDP�㧧�ơ����QC���T7��"���yI�c�R��o�wa2���;�\N&E�s�*]%^;�/䃷TgGM�B>Ԑ�[��4���Dn��G�tl��B���+��a����p8B�3�d�L:w>�æo1��Vh����澅��肼t)|Kʴ��kv�>��S�d�y�+�/��U���o
?g�r�ՂnH�zD�c�no���tU)�W;0���D����̮Q�W�F9~}c#�39+6���ۓ�~�������F�9��X�ӣ[�w�㪯�a��v�̋w��7�#X����;����B��S��WR�Π���-w~�l׷Qzx/5Zb^8h�����e��H�(�f2h��6�T�1q.�ָ��GN��㳘�>�cj��U� {10f�K/ۑ�'6��5���"\G.�9����k�w6x����H��a��#�� M����m;�L����HӅ��Q�oJ2��^;)�υ���wn�:�������ZY����q"���}����uT�?Y��O��|��$�ouZ��22��K�צ�4v�:j.7�5�e=`T1��w��ԁ�-���
@�^]��<����`P�/���w.�3+�@��g�����Y�P�CE�?/Ej,[oT>OΣ>Vp3*�u��W�v�K��K�nՊ���r�$��zO������7���p�j�.��=Mry���+(��ޞn^����@P�*�ִ��]嫖�PǗi�,�"������>�.S��5f�j��R�0ޢM)[�r�������>��m+?q��]�kwa^��y��L�w-ɝ��9	pzit���L�?m�ʦ�^�4lᄫ�|3�����WS�g�>�a����nu^m�0��}k�l�!o�yJ�K����F�=tse5�+Ԅ����7�H�h�g�5���S�
=�Ȋ�E17�ZBΝ6|QU�K���p�G�6X���:�Ҹ�����q��&�}�l�K���3L6��,�s1��pq�P}����`��LΟ<`��^����M�.(��2hЫ������3/QU"��T��{�M~�a�?���|B;����>z�Z������_ �u���=�Y�}�X��zikb˭}�cer�:��>>��O�rF����K1�c���GJ��2-{��zC�=>�N���\E�G�����u���)U��F�=�Ր�b�8���P�S��*- ��xE`��<�|�}r�%��>���k"��G5Q���	��}��k�-D����r]	 ە'�J�S8b�^��NUH�BG�'�#<��k�����gǎWx��l��V_/��/񳌢~�3�Ob��q�J=�B�ٟw����j��z~��?x����:_
�>�M��c�S�c*�ei��<�:���9�!��)Rݵv�e4w�:qX�$�ܣ��M�[`�l�1�4��}G��k�js�Vʭ�y\2��������!ڻ��N�~��!:��^I�yTo�(�Kz_�����c��ˋ�od~��|Ϸ������Ǐi\p<�`����weU�����t��_NKʇ H��k	�M��N���H���"*xS��?OM4-2Ơ|��j�v\�y�O��-8||5a�-K�7��R�3��m+�����9	\Ʉa��\���.�m�VpP^�+L�����|�iB�q��w0m�_����˨]R]+|e�ʓ����n�y������:~+�}y��x�K�sH��MZ�C�q��������z)���r�x�	���eF�lߞ^�m�9q�Q���L0���_W[r�ܕ�yY�ɀm:��;��sgD$z7r��N�7��z�����b�q ��,U����G�%�8 �C�qZ�N��γ�T��.�Q%b����L*�)��8U���ngAv��鐌�l���=v�I�K�]ݔs��|j��ۦ��DQ&�3wY��phM�����R��e}2��ށ��6a�*]I�T9V�
�ʪU+�Oa dwN���.�&0,���Ms�!vh��kZ�Z�r��Z2�[I늫i���jݞN����_KZݼ6�P�ך�V����ኁ{rR��A�y\����<�\��ƒ�/!�/��λ.��5��k�.�\6���&pD̕��J�L vj"8ʻI$�wwwwwwu��'/�ā�l�V�B~�rȡ����E����1	��"�6�&���.����qr,9%P���`)�廳f�P�i�J�U�N�K�N�(IJ�����,�FEX���B�.]��)�8���,J̬�U*/;�����u3.�[�LYv�yi�B|*ͦ#!5�Bˊ!��m|���ŗh8~�2��3?�Rcm�sarݧ�2+�&�4~v��i���i�
�&EW��p]UWʞUKC��u�5֕f���Sũ�e?�KQ8��D�Ĝ!B�r�9h��IUԡT0Yt��Uw&Jp՛X��H݌N���̷����'Pe[e�/PIZۯ1��[߾��w���AQwIcڊ1��1*`��"Z�EkQX�Q�Wi.l�V��V�,�!iQDQ�bPXa�Tz�Tr���!��PUFұV
��-Y�c�b0�
��(�A`�C�(,(�"#"���TQC)U#�$�1��!�J#�+Y�EQU։DX�r�"EEE6�H*�)�+p�Z�@�Z1+V1b�ŘdyJ�$U"� �O��)�+h�A�o4wd�6�ܜywY1Λ��mů����M�M�ٮk����r�V㗙��j�]����7������H����s�l_������Bh���Ι��5
��j]��n,#uY�m}��/N5f����U��e�5T��A�ۖhb�HV)�c��Z��i,(�����~�fg1�r�\^&l���#	8x�D#퇦����G�ӣ�ޝ2����<wUtyi����r�t��w��ia��x������M�����'!ړ�����Su��"�p��Y����iK��;;(¼�kg���bm|��!dd��&r��a��:��]�cI�<t�������(�B�x��f���w6Q�&faƻ�J�L��rf��G�q!ٶ��꺊�P���Ԧ5��C��"�yr�Ԉ��ӽ��%#�]�}�eJ�z�W�ߏ�rt��@�h#ٯ�x�{��ծ(�
	�q|x�&tʧǈ���z�V���7�{{��G��`ו�#0f�2��zQ��r��WV�vJ�6�0�,?QSsP*���O����*n-�%�~At��~~3P��_�Ѳ��7z���2ԫ�,��p:���m�>�i��Q`U���gK����f�\N<�Z�*cg��aT��Peml�?J����U(��Ө��N�2����&*aK���eCȁ*X�G�t��\p;v�)ً�xgeI�j�ow��ݍ��h��1X,�rd��]��������-��^�(��-i�����owc���v�4�N�J��WXN�*��lwobB�9sU*Ɋ�T�TSH���'5��,�W%�w6��G?���t^~]�^X9�-?�@��J��Z�5�g���g�k7�@mi��ڷю/�oN���x�n\�x���26��GM�˸w5�k�u$���M����UsoAի"Ξ��~C׏�������o!ϴ��x���]��bw�C�����N�'�}�D�?u�B�T�s�+����dS��<�A���H�v!�\������}��/���<h�����c�2�$��jv���v¥��k��a���>��4t�F}H?,9��<��Z����a��o��P�?X2֘Q6�]/;��7Hp���%?�l��ly"��T�,�M�+��ʛ��ݢo��+��{A��Wq�Zj��5F�p�b� .Э�L,�D��o{�4�G,�\6yTu�u�Y�+:�(��	n�qS�H�b�6_������:x�ب�!��i��u���`<���o��Q�#b��E7ftіz�C{��{n����N�ĉW�����ڄ)��(�;����*��3vL#Ey�ϵg�FZӚ��6}p�M�5Gb�ͧˁ"��RU	��f\e\ۨF��32g'�C�aOUX��g���G�_�4	���i��p͍�(j��{۪�8ن�\h���M�����9q��oλ��m�9B���V��+�S������	��yb�4̥c�p�LA����3f��+���ݦt�嵾�*��h��M��j_���j�Ś���=9>���u��2��ȶe�^!��%����ۺ�ixwe���6�4^lX�N��(��R�k��u��%�ԩn���?z/x�	��ߕ��J�|�J��&�)m�<sU�o�5����V�ͮ|u�g�}�G�Sj㥜�x�m�ê�K�ݾ�ig ңt��8O��t��>�#C�+4����,�rg�e�����k�#s=Ԧ�B��;,ғ��7�@L+ �0<����gW��|E�d�-;<�#�ˉi�$z��L���ȑ��\a�,����tT�=��s�3=���d��ؾ�+Um��7�M�#J��a��ڭ�G���_	��׵�弸�&Y�W�v��]�b�|u���N]�]j�|kT7��GN�va��,V�\��V�V�=�Hі�:d��8�V��A��8Y�Ӕ{U����etjQ��s�YU�+A�yku� � Ĵe�}R�Y��vT��O	X��Y�i8{�p�{ �1"�o#0OJ��}�x���o����~z���O3����}̸�_�%2�6�]	]Jj`d+�':��^{BD:��t�9t�Ԋ�Sٽi��Q2�G\��<��4�DC�1Q�ZQt�N�T|��ވ��^�9�gH���!Ż��g�8j��_q�2�N#�pk'؁�|�Ƈ"s{����Fj����֐=k����G��ߘ�K�[{��P^��g:���]��X�a����8��9i���&z�?�^Y�\�h�vv���,"͝j4�=KH�������\�Bc�byӮ���޼�J�OUϜ�#U��!q�Z��L���d���y�
&��B� �l�E���{U^��b�]�0�ZY����Y��[85����.���[�v�Wh�*=%d{�a5�yi�ggP�0��9��wh<���,;���\�g�dGHU��8n�5�hy��1�z�oƲ��*#�K��8���קԳ�"�u]oF�L�BW��'��J��J=��`�i�<|o�LZY�ţC�k|�Ȭ_�ݻW^a��p��,)�xC�~�n��ƹ�ƞ�;��yW#�S���N�tpR�80Vl�;��&�=���?t��/r��1���_j���6s���V뼩!游��e$,���<�HY:����\��Ϛ��<t�*T��' U��������m�A5�G��.{����z��o�k��R�/.����.�Wu��G����qO.?lƋ5��g� �2䨴4���k��yvh��)Z�~��V�3H< ���v�	��7Nofv]B�w7&�ˉ�A��׎̽��dS�}D7�����0������G�������0�ꠦ��7"!b�D!��r,;�N���mQe��!q����.Ό���H��#^�Z�S@����\`��US#lI��S3b���Q�r!�l_L���~�\꾆��Z��z��5��xwW��xl�Uz���x⟪:GU�`���x2f�8h�~�'�@1x�\�=]7���᭘�U>�Q�!��iq4�(�qY��~�W�<�7X��_Q&��8g%�Q�966��A��N4=N�WrI�Ɋ�@�E�$N4��8�sx�Iڌ��^BY�ͱr�Z�N
pz��W�$}�\4}�woD�:jwK������6���_s�(~�Ԟ�u����y�cg��&��S7Y|���ߪ�Z�{�ڟb����G)�����-jg�39����V��o��`����*<#���?s�8鷶7b�Ѧ�|A#L�CG
������Q���ט��`�������
�LI�un
|t��P�/���{}v;5s�W��f^h\KW3�*TOH&��6�Û]ǲ�X���eqX��Q����������)j㠳���Ѥ�銦j�y1V�KMu�"Z�q2(��چ�B���{��Mr��oH&�?="����|p���M��+��$��Σ{*aå&vj`Lw�S���7FMeT�rzH=*�&�u�����.���F,����5Ī�}`k!�3�o�0u6�f�Ӑ��O!8����`���k�yT�����NϞ�;K,u�v�M{o]�G]�W�Oވ�Zy=ف;<��Q��^�?U!X��� K��4�>���)������+y��x]f��yq��҅p�	�w��t̩�]Qb����*{�9�|n>;J�/�H�V�����г��O��5�Տ�Yv���\p,�b����/=r�߹��x�?3�Y��
�9^s͑�IrMdê2�jdφCl��m|�O<�u"��.������k��O���-%�4�m
:p��oJ5~�yѧ�&���r�,�D�Z����:�g�O�WPG*��g5�ղ���Jً�k�i�b�<����Q�rz+��דxإ��\[��ǀ�[\)��Xr-�hq�}fV�f�\㼳��0h}�ά%}fV2	°k���S�z��5�:56���F�����Wt�޾�ݐD�/ۮ΂H۽ư��}������{���z�a��)��U�i�}��ut��ͭB��(+I��uS��+�5m:�;_k���������׷l��]�Φh�CvՃ3[î�����R�p2Zv!�����Bhl�*�v�嵽%T��-�ܕu뵝�������Ww#H�ko�d�|�e>d;�_�Î8�4�o53�hYʴ��!�G����@y��t�<��er�����2��&h���qف-'���cJ0�P#mot�`�^�/����,u�l�-���n���P���$�I$�wws	�/�d��U�bW�Of6D����p���,�pv��dq�9�b�X���VJOأP�3��Kr��v�P�����F�)����VU���n��Cw����[������Qp� �����VԺ��mT.ۧw�
À�v _c*ѱtJ��E���ff*�ƁW�X�cAa��WmTb�-��[B:V*YFear�a��a�iS��j\.D�e�t��	ѨRVc�
�;�&U�J6f[���X����&J�)�c�qf�"K�Eg�Q���e���3*��BR��)�;����4�4�Ů��ąS�*ĎfYy��cƮ����g*u���\��y��}�{�����F"�D8�aR"
)�����"�R(/
�K��a��AA,�"�1��
�,PYa��+���"�"����a�EQbɫN�*(
���� ��M�EDB,�R!D�L��"��TճL���,Xe�dX���TA��SvJ��T�j�D`J��EPX�iY`
	��d��B�a�� $~��K1�T3���a��G��IY�a�&k}(���6���}_{�&�94soU�w���V����ů��`��w-�h���cRpLvY=^n�ml�>���S�
��U+ŷ[
��)䧾+w�j<��
۹���fi��r�%޽$��0�+hH,���9�a��̑����p�\d;��|-�\8wT'�V>rʠ��݃X��fe���*�.���Pq Uy��7tm�ο�<�	�S���\\߼�7P7�U��y���Ir;Ay��N֞U�l.�]�I�h�8k(;���^�G�՝��,�")�j������D]kPv97i0ř���UP�GW'�/��WՑ�;�6��,��.\�LM��E�U7Z�ʡ)��
v34�Oe�+��St�mk�J"kn��;�V�W`8��[�WL�ְ�&\b���^9�ˌ������f�/��7ۮ��zS�!���ҧ��K�ʥ���}V��|�#rr��IY��1��n���s+pa:o��[esP�\�\k���d��"m�U�`����ˇ[q}���;�)
cS��+0o�����mA�n���>l^��e�gf�~q`|rZM�{�����b��N��λh��Z�q?�}_R��o%�����=�E&���u��1�&a��p���Q�pk��j�9���s>^}����Ns��p�#��{vx�t�+M��=�P=����?��fI굡���q�������i>l�Κ{����3/Njۇz6ö��y]�-m����ͥ35ج����?9��\c�E��IE,��Y��:���fe2َ��bҨP��0�P����U��5���,َ�|��r�'\�p)�Tˏs���T����=9 �$-u`�m_�*�\y�u�ZAD�;S���_>���y���BI�V�����T��G�<���6���5f��Q�ݯWt^3Ff�8o����QR���=+O.�x�!���=Lԙ���c�煄��A�����kO|��)A����Dغ��~�)	q�q��C\V�P�u�_�}z���I��&�ݺ���]qI�zo���=S�HC'�`]"��Ȥ*z�T���°![x�rܣ͚F�M�t=����@M�e�5|�l�M]#�oM<����*���i���U�]ף�F���>�hV��)��5�`�Wm���1�:�:/�Z�įz��7���6ZBg8�����=�"{��ߢ:;s��	��(�/[y�� k���D�C��1L�{7Uͣ�A��xj��˼DB�n�9�]��*m_l�k���+cΎ�h�����$=L����к��~��2Klc-uh��ꈶ*�]�*wjH���}�U-���[
����Z�����vx�1ͣi������� WF{��v�Z��#�6f�I�"��x	��Y�o�f��1���櫥*���:q
�B�v��6�)�gV8/j'C!�8u���n���M�w)�r�> k��ֺ_Go8Du)��SIO�z"�)��>[H���$��\��'z-L��m�� :�#�������$����J�m��rw�<qt8'�.�V���P%�������^*S���͛�P{h�����#���w�S�cه�@b������Q�Jo�$ь�m��雂�V�Y��Ӧ�OUzw(5�T����`KvS��R׭\�A 9y�y�7;��L\���ó���s��z���a��R�w,��Ǝ�h�����V��9IX�>�b�)��ww:��+T�ot�ޒ`f��c�8�YKJ�z�/��+d�'�O��g�u�#��ˎ*�k�6�v��lEYz�/xË�6�`*�[d+���ӄ��\lu��m�ש�xff��3[}����h�\��[#���w��ql������5k���<������uz��9��L]24�2h�t�Qe{�k�Qz��|Ў�$�wqY�|�-���ѹ�.�[gdԫ4k:M����=2D���uY��C��n7=��ֺ���7�u5�ж���G=̷.�q	t$�.$��j�$�V��B�/���d�Ç�Ec��­Z���ѥ���o��n��el�`��b��N���f�K�m�����R1�$��"���S����F�6:�y��MA��#ö��S�q�w7<׼��I�bn�KȞJ!���p�˭b�볢� ��A��t��,�B^_c��:u�������)�1��Uc��<(E�Fr���o�.V��o�I7yUυ.�d��1f����&e(���4���S�r�xR"㦻�t3x���uk\d��9=����&�v��Aa�jM�L^��z0�S��	G��7t\��dL�9j[�|���k�{��.���{+�&���(�T�n�K���؊�"�;"����N�C�p-VR�ܵ��f�`,�
Į��
�S�~�mLw�>�%"�W\�:�ޚ�m!�u��#�a�qZ@�Z}���<�"�K�ʨ�jV��2�̣��W�-�u�����l�50�C�wU���:�[(�n�f+��`i�|�5�;'3�E�A�NRʨ��RV�PƋ6�Zt\�t�f���}O�Z���ң�*�^wq>����΅�9'K�^��AL���y��6yJq�@����2�vA�����Q�\-����5oZ?B[����Q�{�lvE�v5�BD�#��>���)��V��������/��&�D޼��񒼁@ɉB�5�ޱ�T�u*f��i��12�,�Z�U��v�dg����)��V����b��
��T�hK���3m��k ��'���G.�G���z[�哋�N����78�Q�tD���csy"�dD�L���ّq$���h�p�S:�����hlN7��;K�������vp�2�]i�\��.�-�Kk̶��ae��	]�O	�C��U2Bo�7	�qp��Rո�RB�r����t���%��f��������2�ᯫo���ɂ�MdH)ۓyP�ܧn��EMF��÷�d�ܧ����ub�n�B�3�`�In��Ht˾z��E*�S�-��'k�yI�%ύK��+_�ˋ]Q#�VFӾ��ۢ��NT�a���e��%=Ҍ���by�i���G1�Ԫ�B82��p�c}��@S��f��ۛҶ��a�2ԠZ/���#��95͏-Rh&gb��w��a��2�)]�bv�@�w�F*����e����9��t55ظ��AHhCn��X�X�Ε3��U8�����k,���.h�����=�)$�I"I$���Vݬ����[�pmbj���`��n����.N^S$�D='�:SMW�"��7��)�MЫ�B�*��y-�YG3�hG@�eI��L@�_^2��!�mJʤaUXs�LP�Be4)ؒ7�Q*�^Ig����唐�ܩ�ϰ�+�$�9Ae��Has�n:�*�xo�*�B誥�U�	x#�K���WF,�X��Vv�t��Ҹ�c�]'�.Ҭ���Fr�Z����xM�,�c0��l�ʰ�`ˏ4��[m�0�V��}��@ꪱ&�,H��OX�d4���+$PI�i1�TQAb �Ԩ$R���UJ�Qd"�"��Y�<L �b+VAJ�mc�Q���Ŋ(A@� E%`,r���m�>!*Ad�
0#����EP�Q`��0¢�UdR
��aY!m��8�p�VIƠ�I�N2AOb���s�2��n,�Y뵓�a�G-�����r��Ei6%���F�y����A��7}B��wh�I��k�������phZ�j9�Wv��z�ڥ�'X*=NG�wp����Q�Z��I������ �7�!�^���ϱOw��A>/4G�P�ؽ��`e�@o 3�j�'a؇���.���:��v�bޅpv��\�zj,G\a�D�0+.��mo2|���*j
�on�}���J�G�N!��-d��di�|�R�.3�}{0�aë1z�5�<��'�5FzgXc��������L����o�Q�̉�uϮ�R���X�=����nUK�i:��p��w�|��w��`����D�ښ�Ν��9/V|��PF�6V�9Yz�/��ʱ��1�[Q:l�^��� �TC jy��;�(����w��}b�aa�͎]j�1���j*,6rwq[��cM�Vyt�z`�@������E�����l�p�k[*��d��W8%L��0W&�˻{���t�0�!�.�cKZ��-e�����V�f��Y�;6�^��M��]z�A��DL�s�
K�R�4gVvڥ��]���\�����6m��z*�F*PP��v��=ys�(�^��*�˩���m�-���˗>����&gw����TZu\�����1K[��Z�Y(�૳G���v�w���}��=�ZPM�+�o��_2u=}=,mf�v�#�7eE����Ŕir�=�f�����ݜ!k�q�A�B��u���t��z�3[�PWtM��񉱝���a���-cJf�T�WHYxv>�[Moe�3y���B�⽢(��a�8N�e_]�Dm��X�!斄�w9%:�w:e\�l�Ȇ�\�Z��hu~��&�c�v�{��ikPt�v���[�5J�l��l)9�y)S1� ��gW��}�[ �WgǦ�o��t�1��
�&Iop��5&��6!��u������XĜ�
ױ�7T�Ǜ��+d�uu�Țl��5�I�#��[��#�F�"2�˯N�|��Q��3ϠشG���q���{/w(09��;db�Y�5�_�Wu�
��Qsѡnq/�^��2��2�sHsr�v�'l�ܲ�X4H��e�����x���C6�Y �F��6
ӗy���c�1P��w�y|G�)uE,�}��7wnb��A����:�`�wY���d�����eNU=(��Wܫw��}��t�_g,�G諲w@��-b]��ep�����X2y��o��*�o\�i�_^�"F��xfD|X�n��y�)��՛]I�{��%�mDύ#6�Bu�lt8"���3x)�TQ��'i�+���F�&8�dkA8���毞�&Z	 ��Ψ��|���d��YڞiT�������2Y�z^̻C@���:r�D����o�W��8L������:��g�=���W�n�׶*s ����+��r���i�G'evR3
q�fC����g:�dl��E}*ݵu��K�@�v���w.�-ꂶ+�Sef
��{_s%ᬊ�|K��,�ӿ|WB����X�4���V�a��G^R�B��H�~�o��z�Y@�.Y�O=Y6�`��=9��%�������8����N����6� �Bh�7f����|�e�q9V�;�jyc�i��!�g���3],F�%S��ygTw�gt`���n�����ܽ��PFw�ę@���j��9�8�s��d���ҹ��&O�]:n\�^kP��;\�D<,G@^`��8�f&�����@�����S��ܚQ#J�_r8L��5u+Ϣ���2��~��oinnF��g���tQ+���}�d�Ό�B�$U䥔�~�ݢ	<�S67=�j�>�Rʚ�-��#K)ڴk�\Ί�p�N���3�	[���{�.VFv	�7�����G�/q��Y�x�ƛ+S�(k�����?`$>�t+��5륥'���O�X	��=],6���N�dE��|������Cs�9�I#+^����vSm0����oH��FOU�D�8��d>����������8��4I¹�RgVv|i���l��)���˺e>8�!#n�-�!����U���K\���&9�Ms\*I�h�5&�u�ܭ.��`t����' ��<x	�u��{CE����p� �1Z*6��ɎQV^w,0,�F:�5y��i��#�>�����(�jBb65{9�z']�+����I%p�|�X]�lt��ⴋûsfzyЈ�Cy7|Tn�r�s�N(����ƨ�o�9��K������@�'�	�b�U���޾|�-��U�q���b�!5z���V�K��W�LX�����hd��:��cg�{�C�|�>�&�vL�ۺT��,Q�nS�r�ԴU8����u�>�SH���K�b��E_*���q��_����:o�۾p�8[4*��\t�l��J���J^(K�v�
dnp��	���M�+ֽ��L�C�~��K5�����f_#�E���8+F�uξ��������W[๨�H�4\��G�m�=�{T)=G��]�=[���<�{0�Bߺ�r���:u��N�Y��b�u�7�7Z��bח�*n�q<9/xUէ�M�+�v�ÞS.���Dm�s�m{��+f��|�	�t{~0�/����Դ�MG��7|U&�U�|����[�?�8�]�h��S|zf�Z���'���z� Nrq�=^��.�W�[3c�^r�:�Yt�>Ӆ���=�&"�j��I6.�}��� �u�/)�7�����n]�:]�<Fd�d�^�W���$�^�j�E��~��Q�����i�ZV�x�O3{-�K�}�#+�!M� ��8��4�ÑsLڞ�\�x�kV��GD��.�Xw���"�1�רsΗo�3\GLV��]�N�%V,�����%VQ�V᚞q�Y�M�\t2�2^>J.�J���[����gFV�v)wV�bΓ��wU.
�V���X�W�v�G�55�u��&�A(��hpz!���f+5�S�|hm��ݨ��5�U<�P�;W5.���		u4^m<xF��6ɫ�ӕ�$�ov����ٕ����f��F�p��63��W�C��o
��{
���y�u)E=�&c�˃rw/_cr�b���J>X��|4.(�jďm��i&�nU����(�F���{��b�SS�KrrYʺ��K�����	�3�.��N@��ʋ�np��=l�#�]Z7�2�F�u��1uHm��Dj�n�c�}X2��o��f�ιYඑ�܇	ڍ(�ʪ�^P��U%'�3��~��w7M$�I$�I$��M\M�ʺۊ��y�C�Gn7�;�]HN[,����5R�\j�����4�p�^��S�Y��=�'��$����U�NOR��WVWR��}�_E�}/��Z`��r���g�*���Pn9����F]�'���ʧ���Q���Q�������C�N���d�L��|o9M�w+�;����{H@K�]@�WH�G7P�Ɍ�̂�Ӯ�Z���߹�8M⥔��j�|f},��N*�������-����{t{[�2�^��̓�	�G���q�Bk`��WfY˓g"�v=�XLPr��a��wg3�W;<���a�F��A�-=��7sZ4��Hr�$Y�����*�T�" (�Oa��,�R��(��P��	0�"�5
�lYR�"
VJ���(a�TQB���(��`a!X#*�,**�T2�)AH�J�P:�͡D��`T�*TE(�M���0�ű`-Ak!P���{d�Ab��ReE�]50�
��d�U%k8ԆDg�C�Y�|�RR=�-j�gM%'�U�����΁'��3���� �@�ۉ��	���x��	pMl�"y�foz�f���gCsVpq��c�s�o�0h靧�Xͪ���o��/�L+���9��X�mnǭP��N��2�L9[��w-�fv��n���]DU�G�����
fk-�T��h�7X(�J7�ٲz�oB����YlIϽv���˅i��O:đw�"� v�l��o�a:�\٬�"��1�T�r���}Nv�S�Ŗz�j���Ϊ|o�}ghP����U4��H->W�Ż�%e�u<�_!�ae��v��VN�����ڇ���0Y�����~�Y���\"�����V����׃5�@����(t�F&;#x�'S�]m��'���]]���d"�A<�[f�ќaU8�_]|i��%���o/���13����:��R��6��QN���v��u�ٍI�`�fk�g��O�L�E�6/�ۭ$���P\y&ʋ�%��Ŭ��3ѧ9���43x���EDに˲�x�uNP��Ulݩ���0�̧�9�p�t��Bu���ª��̞r�2e,�ڣT�Y�(f�Υ�*\�fs�d���9��=�k+�@�u�����Ǉ��X�,9�s9�s\:y�ț���麌��X�s+y��b�Sp*7�	z�ùB8g�P�}�#'�0]�Ν�1��B���j�MR�b�6�Z�e�� &���~���+��(瓙U�R+>�d�'�?�����@��2u��;F�1�dy�H�^4�cHT�n+U�e�0_"b貱�3���R�&�9ٜF(Ӯ��}��طv�v;�f8v=:�Dk���j����{��7�nO슢ƙT���8S���A%�ֆ�桝eJ�c�_XI��u�j���]��:F�z��M�r�GY�3ԟz ��
���|�����_
u(W��X��o#��D�3Oa/u��Tc��ZG�qEi���
v~�x
��詋��;��c��{}��az2ɏG��#ʏǠ�x�  ��<V�6���o˶iU�a�t�$�PX�T1�6ftsb�l�-�@շ�܎�;da�_�@y�F�5Xt�
�5�Q���p��ݷ��E=�*O$-1ٛ�/v[�ꩾ�
Yp�z�nM壩5�*�%�6�۬�Z��n�V�e[���|�S�-Fd<��IR���������f���ɫf�7�����pGcO'���`_�(�8u�<�k�'iz=�N7'{9
_��A��uX���_:����ײ,�R*ϖ�H��{U9�|�D�Z�i��d�0D��jsy[��ƀ�ἻT���$��f�Sk�6��c$����q��J�a��_3����ыW�f�S=�F2�<���H�6[g���{�+̪��b�����T�A&��>ᷗZ�Y�«��g�3r��X�W[w��q�|kX88��5+<ԩ%ֲm���
�y��.1G�}a�=@��[��^������?���_�S67=�����s:5bU���Y���t�=VW���>�����<�aa����LՊN�y�����v�)��R}����@�ftD�z�⮋|�M�/S<A��km_�=Pr�t��	,��B�>QbI5㻞�'W!O���扥2��or�X2æ�Dޑc"��B;�[�ݻ�l��yMb-w]Rw78��e�݆f��+��\�jz&����ܘ�*�bp$��CU=�pR���%�D�|�����d�΍o=R�]�$Wbʍ�"��R����xoR�q۵��6���W��btA$NЈ춣yV���D�g��#s�'i�LΞq� ����W[A��@��葚�������f�ҳ<nD<�Sssp��\����$�Q^ox@ٶ9x���1>�T��>8��U�e[����Qiߋ�1�q����m���Ry��uky�C�/���G�$��ڮo�����*n�׮}]p��eK��ʢ�dp� ��+�Kdv�pXW+��g��R'Ï`�{�}���:�V�[F���A���{��hgp�x�ԟ\ەn�^������(�F%m��;�����ҝN�����#6�"{��xk���v��|���kA"ٰv���IJ�|/F�k'���Ԙ��3D�E�����.79߯|�7~�8��q.E��=� x��!��F��Ǣ2��"��%�W�%���	�c>�BC=#�'.���P`��5qY���Ǫ`���묌�X�zPN�Z��6��t�X�C��ö�-r%�f���D�W�����\��ŕ�)�ؖ3t*�̮/N�O�x�>��Y=d����G^߹V)�^0o�"��̥]��ڗg#���.�9��%bW"��5	�~�8
+�<�n-��z>���2��g<d�a̴�V����Jʲ���rR��g���r����Vd<�̪�<�ɝ���"�>���F�Y����k�!����}-��@��1өH�r�C��~X=����tE�D�J�O-ڳմk�iX�Uo=����U@"�/T�K�R^��W����~�|�(6�p�{�c�f���0��W��������n[�vV�D:��tlxJ�tŉ8m�:.Z�SpL��ؒ��i>�ڶ{�g"�s��L�w!��vd�y�;z��%v�y?T�-���oG��}�Y�uSQNj�&2pBӍfv��K�1EFW�&Z�;C��3��[�r4��ME<�#S���)췬3��3��c[ie6�J;�JѳW1o6�:�Z�3+�Q(D$o�7XM{����i0M�P�\���+b���ҁW5���E����4�|NW�*-�]0���4.y�l�ߡ���M�[x1O	ܜ��Xa�w΁��DA�I�������I�PUZD�������.@���Z��E�e�jK8Nx�V�宧�K\��4eZAAUl�f��(����"��XK�5��#`�+:d=��i��U_#V2�#ln����sL>sK����P�#1�9�o���7��&w��o���`4�,�l�(*��4{Nyg^X�  0(��0���*��шIZ�?�+�7�o�����O;|�?���t,��y�D�|AUq���?z=\����a�����Z{Y/���d�2Oa6�?*�&{)t!���H��q�U�G���s }�+�U�� +�'eO\�,

�W�(�!���S+��&��Y�=v0œV��T�w��������km�⹽��RC��.)P��@i������z�����a����>��QAUm�ˢX��Zj���=���B�d�`�}�GB�������_���DY6���<�x�~�f�B�<�[���

��� !�w�p���3�c�g�I4];�z�u
��ي=������b��N�&%v�k�(N&�A4�����*���DD��ƍ�!C�(
��bF���}y��b�,���Oa��?p�ø�\h򢠪�4��iݐ��x(*�W��ف#[۬�g�1�i4m3�h7��;R���n�,|N@P��᧓ۦ!=I����٘}��AAUz���l6����%^~�hb��U��_��Zǚy�m�G���֙�A��;�:�Ln-OWI*A��yꁷ���ӐZ��ȇ����������@m-���`PU^]f��� �~�j�5.��w`A�'V�4=Pl!�L:�;�,C�,/f��B*����C����<�n�� "����lH�s�p�#v�b�$!l)ҏ:R��Q@<�"���;\�.�p� �ؾ�