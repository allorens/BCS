BZh91AY&SYZ@+�v߀@q���'� ����bK?h| @    
D ��(�ҙD�Y-�AT ͔�5U!fTQJ�m&��	H�U��Ԓ�lh��+Zj�dT�E#}��$�Ҥ�$� �T�"�*��u��$�4�B�T(;2��H�@T�4)$J�J�*�i���� �yRI�� Ȥ�+j� `�U!u����R�J�ZQ(�0H�i�	[0���l�JSCJP�QIT��4�ld��u��īL1�R

�$� �9}T�4�phh���]ݪ��n@7I\4mF5�(� ֕N�G
Qvs��4����-D�RD)Tu�DUZ�x|��  ρ� (���(;Ch)@
U��@�)�.v�Z4)L�pR�[Nr��P�w]�x@�w�� z�֪���}��O}�k[P�a���J��I   ��w�ҀQ��p����{s����r��N�R��W{{����=��C�
���:*�)�/S�z��K�<��@[!�ޞ��v�$�v�F�����W��  9�}� �K���
t�ǷOR�U�<��B�����)^�v�=ʥP(^x�opƽ�� J���=U {��AB����J��R�	��(  y�gO;| R�˼��M ��x�$�u��<�(R�������S����B�����|�=��G��]������[�w���e�6�"��T��mb�I�>� �|}(
kXq��U�h����J�r{�҇����� *�z�Au�K:u�(
Λ�R�X1��
QnS���{b�N�@�P՚k
TH c���� �í �� 	�g�@��v� �� w� ;�p �.��  6��ERRٶҒ+&��y�� 9� 4���@��� �� i J Cj 4`��� 
�T�i@�U%��i� ���Ww� 	�P �0 tw Զ@ Ѵ0 ���h�� 	�n  A����DM�4�fB��T;ϔ� q� �  �& wt���.�8
�( v� � tq�   �    >��    �JR�� b Љ�0�**2b`& F�2a20jy2
J�~�      ��JR�M ���M`�I���T�� �  D��(�"��e=L)�i�z�b<��=5>ϰ�g٬�����>�v�!�:�$֮Ms�}��tN�9�d�w���E8K���^�� �� �
�Q@EO�AW�@~��ȏ�??�}��!�?���<T�dV��$�_��DW������CQ9"��������81��fpv�CY6�md5�k&�M����س�d5��!��Y ��g�Ő�v�d��k!����dŜk&,����Y3�v,�b�ŝ�!��Y1dœv,� 9Ʋ�bɵ��M���ɵ�;v�M����d5��CY6���@r�œv,���gb�ŜLYزg:ɋ8,�Yس��8,����&,ೂ�&s�೵��;k8�v,���ɋ;LYƌ�Y1gb�k;pY1d������9���Ŝk!��YƲmd5���s�ɵ�k&�q��Y6��LP����L`�0.1[&��k8�M��s���Y�Y6��d���ɵ�k;k8,���ɵ�8�M��,�Yd�a�5��M��YƳ�d5�k8�q���5���k&�CYƳ�gɵ�k8�@s�;k!��Y6��gɵ��CYŐ�YƲ�Ő�v,�Ygb�kZ�s�gb�Ő�CYd��k Y�CYز�Ő�v,�Yس�e�ŝ�;v,�,�Ygb�ő�LYس�gb�œq���b�Ő��mg�k;CYƲmd�ɇ!gbɇ6CYd�5��!��Y1g�4gb�5��;LY1dŝ�8�v,�g9Ʋ�k;q��YƳ�d5�δ�5�k;CYd��k;Bɵ�k&�@,�,�Y��k8�q��YƳ���d�ɵ�&�M���,�Y6���pYƳ�g�k8�q��YŐ���gbɋ;CY6���Ŝk;CYgmgb�k8s���;CYزb�LYس�gk#��&,���gb�œLYس�d�a�5��Y6��5�k%�CYd��k&,�Ye�ŝ�&�M����ŝ�;Y;v,�Y1dœv,�dœpY�LY1dœLY�dŜpY�d.pY�d;v�q����g�Bɜ�YƳ�g��8�LY1g��k Lv�@,�Y�9س��mg�5��k.CY�YƲmgmd��g9Y6,�k8œk.v��+��0\b��q����k&�@,��,�Y�Z�����5� @,�,�Y�YY�Y��M��Y ��mgmg���q��1b��q��� fM��ɇ&�M���L���,b�q��1��k&�CYŜM��Y6��gɵ�k&�qdÜb��gd�gmg`��Y88b1W"c� �T#C�8�E�".0q��c� .1Tq�#� \b �`�8�Q�
�1q���Tb ��8���1 q���b*cS*����11�)�Lb
c"8�1��c�8��$b�*8�U��6�5�`,��bɋ;q��v�CY6��d5��q��Y6��Y�rmd�b8�q���+���B.1ddزgmd��5�k!dÜk;k;k M��YƲmd��ɵ�9�gmgmg���� CM��Yf�3�8�v�@,���+�@��H��~����=~�d��7�?sBuW,�"�L��۫{�u�B�M�ƀF`����B�������"�ݲ�ey�EN���谲�A̹65OM��â�&����8��ʰ��W���ӣ"N#��ޚ�a�S`д�et]���x(RvJ|w(�ު=Wca�Ne��8qd��Ѝ$��+���R�޶��gH4n�oH�w�9^�s1]e91���l�ߠ�p���Y�c&�z�f�=}��\ZYq��$l|<i�S&,+2�"�c$�v��&�*�h��;C)
�*-��nL���t��zj���Inmј�^�b��Ly�s ��[jv3�R��)�E5q��v[=΢��U����
&�RKk$�o�_n^0�sox�̧V�ZU�Ή�+z���j��F�j�	�1���¥CMkZT���*������TG��s5w!YU��f�Q�ˣ
�s�\P2���t�:�
���٬�"Hi���P����V��L
DK��D���4�MMt��Y���]�#����g2�ܠ��8}K��ȗc�Wb�]��j�� �ZB;���&*v2d��͎���í���0����GP3�	Ҳ�*��q����2��Ң�n�n/y�r�g�B��)�km	xV�S�[�ʮ��ɘq��B�d<�UyF��4+��e���Cͩ��O��u�����a#^1@p�J�pk,^�Vn˛qZZ��r���X�e	��o�Fskx�*�$b�I�Y]n\1G����j�����/8-x��uo2��i�8�Ԣ#K�>Yb��]c���<�6
�Z��Ѫ�U���ťWV6�����lX��̭��?5޺�s�#��Ѷ:�b��O.�A��cx���T�fR�wj¶�;�t�x���r��q��n+3cy����� �R�p����r���ZO,�#��8@�iۖѷ��׎�l:�C*�<�VmYYo8�ɅrҲnGp�\�ˠ�de;TjwdӇ-S
��/;&�mm��̊�F�>���&�^�}m�h�xk"/on֗�b�G���h˘s�<�p��9�]R�M� ��ŕf�4,�C��o(�`���rJ�,���_V�%s��u�{�r��˲�,'jz��s�[ȮY ����$����fw0�=#*��6�Xt�ep�O)I�F;���a����%ev�ׄX����دq���+��&����.�+�{v4��$��M���%@��ܥ�Y<�a5�f�E-�z�{r-U��mm��T9��5f�|�>|h�W:�A�D�R�Ŭh�4�R*�g ��6����%����]nvY�v�!���m�������$���h�T+F��P�+D�"sJ�F=�HqQu���n򝢳�@�"ܮ�-IyY���[:�mV1m�kdD�xk��n��$�����U����e�m[�L�wa��U���N�.���2M�ifYz �y��OK���0N��.�.n�Df�2���7j$p�1��kjn���#f����v9(�WY�tG���5���z�Ժ��Y�!y� ��zB�`�^eD�N�\�o\o�WF�N�.󼮇�����x�WF� ��c]�C<N��^]��u^G|�2F�"���1#b�}|%���{BdY��V�͘��:HM$#M�#�|�m�ȭF�o^/2*��\F%�-�#3�.��n��Fne��=���vkr�[�t̙�Iˤ���.�\W��ˎf���X��Til�5Z�Bi�����T4D��7uy���,�mn+�J��J�]�O]��W�uZX�Ɓ6��'u��ז�*��Q���[�`�̀jFA[���4U0%W��{L{R�LRl39�wk*Q0�ƃuk���D�a���+J+P�ƅ^0�O�^P�ˡu|{t�o�-�Jb�REvmPHr���HwL�)�B�{��8"��i�U�nau+$9�t�n螕'*���u��^{�	u��Yǅ��n�Mm��Z���72mhn�=�.�D3��j�5�Z�uhO�Ҵ��{/y朴s2EZe6CX��V�f��սٜ���#�)0Vpr��o+�����Ӷ��D��J��N�2lڳ)X���������g�f����;#g:�3ύ�4���4�#[��i���:.�R�	!��t���j;O&h�n�b�A�P��u�Z*�J��a�5[���d���R.�_SJ��˙
y�%%��c.��e�JѴ^�S�]ԁVݞ���ىV݅�3AAd�󭻬Ɲ�ym�ݼ�TJYdU3i=�yU�;O���iv���,AJj�b.�w=y�Y`��ݗ�K��q�YubF�6�Zţz��lb�Lt��^&D:��(�ѷ]l"��"[y��yP�$.�e���NºIS��:�zNm��V���|�3 Wy�.��#�4E�6R��LD���Hl��'2���ӥ�J}۲mF�7]j�3y,S�v<0jճN�:*����(�*n<׉�T�jC�KP9Ĭ�<�3{Y�0��K�N�ݷT�f��կ5�WV�-&-G F��N��T���UK1��&�ln�����7}��yq�o�4�(mW��BTS^�]����[���zom�j�Th�xB�H�Y������QXh���'�J�B-|+R�z$n�����Y��g`dg�0ݼt��yr��'&L�a͉ӪzXѴT�����8J�W��3J㎓i7�[eS�U&�r��@�sm��.�fz�f�m� ���se}[g�d��8�k��}ya^�y�t�c��!+SI�YJ���"s1r������Q�6r�nb�ߕM{B��{��k^.�]����YL��Z۶:�����5��,�Aս+��1�(+-�"��ͷF��Dz��0�5��.O�T��.��2���x��QX7��H�z,U�;��6f��Ru�6��͙�IN�а�ݔ�r�	�yv,氾u}�ʆ�I����Z-nU\��f��qW&a�0�b�V;��ܤ�`;�2�45�4i
�I`!4meRЖRh�i�ԩIk�@�+x��&��XCr�Ŭ���{��.��,->4�p�yH9�$y�B�1U�z��W )Ⳇ�l����D��^�;���vr�^j�8�7a}te��W��7�A�	�.4n�_��QU�^H*,"��N#Nh�2�{u��%���[�P=y�a���ݼ�Ye��2��DD����pIT�fP���c��uyzL�P���q��V��4���p;L����F���[���0����S�y�D;�u�"��D��]��\��0�-p�W��k~�W���1����9�9�k� h��t��`��H1��Ɔ�
�iM�Dy��YHJ0���Xh�%��%�0N�0��Z���=�ƵZ�j��*��̈����]i5�d;'ud��[Kx�C�*����RԪ�R�ÁP�f�e,AQ��-�ۄURR�ʇ��Y�B@g#:;ı�h��U:�٫�>Y�bC-��xkr�bj���WpP�]ʯ��0�n�4�Q���cۧd�t��Wg^���	ݴL�Q/r�Z�8��Jc�Y�~���맩	�V�k��Y�.�$��$�[��ުf�G���Me<H%��r�d����օ{�����H7�҄r�9UThX�Ȋ8v���ADf�"�8��0���CX�p<�܍�Mژ�#�fa�FVЬݑ�H;'p���{�S�ݭ֥z�(4�k�u^��F��Z�$��uz��y���-�Z:밲_��u�Tbtfw^���U��*���w2�PZQii:L*�i��Z1�|��W=ח�f�pWK�wN��&��Jwv�'��~w,��JLENY�X��U�F`��;T�8f�pS�^'���r
�$U�Mf�٪{)f6�j�a CO�i@�*.��e����KUw�BWI�L���u]aբ�N�kUndR��fK�rE1�{w�Zދe�ٯ�+�pm.���ݵʩ�1�[L�N�2ü�n�hZX�����,4���u�G�WŊڡ���*h�J�X�̤�.g����7j��b�U��p�[f�-�V�0�E!�傦��.WZ=�G_q~f�Pyp���;�io+I����l�(���woi*������.�7Xf+u4�Z�iX���r�Ι7V!���;z&;ʣ���{,�'�M���R�cs^!��=`_z�m�K��j��ͼ%o1ܨ7ԥ*�u���ћ7��)��WTc����PNc��M.���T��,-�5��<�FD��6�ewD4݄�|އu2��n-=Ĳ�v�/���v�R�P9�۶p�����G%*j��ne�ݢ0:��I��^����-d�y��]�L���d��\+�����9�#j��\{J��`ʵ�-��>XH<.�=�7�Q"ˉ�c��A��kW&�vh��UL���+��է�*�kUf�`��f�$;f� �ehz�Xz�p1j�����]�nn�<ۆ�k��.;�v��yba�ę�Ӄ����wh��i�}�uٕ��|4S�p��hb;3��h]��LmJ�q,���wt;���
��E'o��JM3�h��3&JJ�PrS�n�2���K�5\�m��\hvڵ)�YVes�D��S5%��4�n��7������zXP/2<�/z"{���pl�Ha���k������ߕ���-Dr�i�-EL��$h�'syn�T%p�Pr� ի�\�]��'��p r���+�j�ad�Qו�4��d�S,��_��u*7`­]�Up��<�f*���^&Z�Q1��-U�M��6�oV�mv\+���t2�Չ^���V;ӌ[�Y���b!��D���TLҵR^�
q��5J��D�g���LRU(�KU������M��H�Ԙ�6�J��J5�K���X� =��A�*���ۍ�Z:$ff'�E>>k2��7X2��qۧ�F%S��[7�v�YmL�x݉����7u�*���Ø���*��[�s&�wt��9,Y�_tcR=�v٧Sv�Q�ѮT6�A�\M�"��1��7��\��[G����e�m�wm4i�x��V�U֓�n��Z���)Vc̓j���=j��c�҆�r\��S[�1�"+��J](�A RhY>�n"�en'�:�؎!���Ӱ,�U�!�����TdGS�y֜=�3�r��i�]�f���ʥ�[��i#�gog,���@ؒ���M���,v�ґ1�c�kt�ZB+vZnK{5Ds&(޽��������NfEY�n��(�Z�+MS���1XlW��Tݒ;:-X�5"T�sGb|G��{-0M�t�˕Y�,��kf��e�BЯV݊��c݌������S4�Rq��U���c9�s;am9y�*�H�u�q���#�i�s�\/Q��,ݕ�q�n�6Η�%y�'���!T��kn�3��4v�u!A���Q9m)Y���AREVN�c5�����T�����Bݜt��y��/��}8mltHPaX���*���j�	G��Z�d^��c�+Nbeb*���Lo��y�n����*���ÃJ@$r�דE�L���fL�l�8��v�
����7d��&ƻ5�����-�Y�v�;9P3*�ڵ۽��T}K��Vb�A���=��RW&�������K!b��W��+;�%����w)뜀�S8��1_hZm)ɃG���#�R���ZD��j�L��k�l��cQl��x�tV�����Y��`�V!�N4��ː�2��V񵽪�.n'�J��$�y=k3[��U�J7S7s}T%c�Vt&*�����E�b�a{�\�y�YEs���[ud�S`��#�ܨ%�\u@ƖMH��ǒ8p:B��kƍfk�=�i밎s|�����n9ϲ¼m���q#y���!7B��kջ����[�Z��ӹWOR[a�Xy>]ɵ��T�6',8��o��Je����e꼬�x��-aD���ݭ椴V��:�Q�9� ;(��wfelL���&->�Фf��J�A\9�=ljT���Q����iZ�s�jrt�b�GR�XKbX��#��O���,�\F�j�YKR���ִ�kYv�տ,�mn�k-^'�t8���[iA��-j4�ȍ+4m[[�y;J*��}]�R��%iWf��bv�W���e�+��n����UiN�؛]�ֳ���+E�kȲ+�v�Ҋ�RZ�ښ�#kim��U�8��l_jMrY򘾤mO��10�hꜗ.k�i�%qV�����b)f$���� ֳ��Wi�@�>�:��s��^iy:U�b){Ҷ�]j51,N��v�*�'i�\b��I#I)Q�E6��R�Ig)��x�%�5X��~W������D�'�	4^Z��,�\駊ȪM�����J۳�}qۡ�n;Yb��k~�ɖ�άiZ�;�mׂ�\�ԛ�0���Vnv�K����K-@]��|���I�O�r�rz�gs�%�ȭ�R&��Z�+y}*Չ*T�E��VWn��_fъ�l[����$��q`�u��J.�ib[�ֵ�倽J"WSIZ��n�m������4v�f�7�WZ�x����X5�4�ԭ��b�0{V%��)��)v�t[�)qki;X��gM*1X5[8�ɳZĺ��� �}˝�*�B��+�y[O��TՃ�lD��,GVR���Ex���֒\$�.WIZ��)k5`/Qjؕ���Y����e��5�J�Z����aXJZ�J�ƕ#i51$�%�E�6�'ԚQRF+"�@���Q-[k5Mz�A�O�d]'�کjĘ=���iR�����<j)tf�b1{�,��u�W�\AK��y�r@�Z]�^^ԁ�^K���i&��v���X��Mu�J5`�[�ܞ�*X�-ߤ�z�J+�ԢGĒ䩮��_#b�s%M(��v4�TR��ݫ�A�S����ӴA��'J�DMZ��ژ2��ԭ�E��W$Z�5STjbX��%�v�ĹRՏ��E���]"ѥnru�i"7WZz���I+I���bE����7�ӟ��zy���_z~�O��5��E_�g��I$�I$�I$�$�9�8M�$�H$�I�$�I%I$�G�I"��Hd�$�t�l�M�I�I�I!�\�I�I$�ʒH��J�I$�	$�E%�$m�R�������:�6��㑌	��Dg��D��F���cd�}l[���h�:���1#�U���u�[
T�Nq;��&
	^p� ��(�IC�ŀ;�ͪ�6��W)f/�	v:�`<V�x7a�W�3tS͏��pG��P�3M�K���)>���h�ڸǌ��3{ݰ�;[gmJ]�)�wb;�e��'�;�e���]�Ȅ��bS/7=�i�!޲mo1�u�Y	��I�n�X�-e�
�J���E�����i�/��1��@Z�-e�JZ��q����f��X����J|�����_.8�\�X��B[�E�^��h��6�2�,s-�5��Vb���-j��<-A�x�dl���w�#wה�8��v:a�3U��5^!دE�ڻ�47�MR[��.� D9v���=9��6�Чʈ޸3C���6e]խ}7t�{�T�b�Șa��&Ǹ�-�c0[SՂ�a�V)��"�.��n� ��9wv�M��ګp~��!��s���-bKZ�e��G*�m��Y��p�<j�i�Ӳ��Lͳ�»���w�ڄ@�H���0��2����8&�N�zɲ�guM�žǎ�q������2N��1�'z�EuL��g�b���"-}Q��VB�,��Z���ࣃ$���[嗇|�	��g)�P�f��m"�T �}�ۼU{��B�Ş�2�U)ܝ̄�0�6=ٷ��ve� �o%L�7�'^�7fq<4+4'm�d�`�;Z�^I�r�����fc ��6^A��F3�%e��鵼7�t���1�ԉ�J�]u���
nc�L��mV�)n=b�ʪW����ؽ�h��j��Ue@VԲ�]�y$4��%��st�)����oA�ok�Y���2�nf��E=��'3���1�뉴DP����c{�%��0*[��A�M)I�}���^rj��nQw���]�r��W5ۮ���VY�N'�����|�|��x�E���ԝ�u���?S��Y_v] GZt�x��q��y�P��XiQ����)�`KmM���K��].�"7k��\��dl;H0.85:���o{;/�Ð�y�i���Sk	�nd�")��K�q���oI �y��@'��x'��qgi��<��姩�Gs�J��kB��oW싣(�۸��V�"�����4)s�o����y,�� �m�&���G��3o��*�*ᅾ����]�R�!CIB�6���
�8X�WI������md�|�����Wv������o_^��a!�z�HX�|k;)vLNq�$�&Xw�����oFP�J��>�S.o�2�.�A�Iޗ0]f#�D�t��xuP�1��;�ø7��o[��vU������v�˶zz�C��ʔ�!7ӃW�+K�)ڹ���U��5�	����Kyj����xh��>�;Q͞E��1�*v�����T��ۖVa5�<��j�j��H�D��E�}�\����/�k��7S����jD�OEhWTf�N7�70�᪦m�t�J�z��u�w`޽{j���Z%g]���le�|�H��1U�YԳ���]���G#f�������*��*dSqD�p��ֱ��.j�K�Bx��Z1�+2��0gD�S�β�;6�
�����ǧ�����M&�\�z�\2H^\,]�3����8us�zf�+8 ��U{N'Z�U����;U�,�Id�C6�y#��83:$�cc���<0�1a	�� �ɟO���$V.6y��w,�05g������){Rb�W���R�y�U���y��O3ܠ�s�{wq��XdMvz���b�Ђa����[�r��[o�bԟ,�o�d����PovG#�Ԛ����ݎ��Y%źbS\U�l�X�j�<`ݰ� ���r���r�ywb���0��Q�����{[�Md�x�ge����j�l����] �6�I�n�z�V]*�h>��fUaR���qڻZ)�z��s# �']�� w���u�i�O�7�zI�I+�w�Q͝}Ei]N���y-AU�E`Xjj�p칲��Cy.�N�Nu��:�ft�$g�&V�Ҳ��0V%\d�Fp�t�0gc�4&Țl�<5p�R���Y�- ��Ψ���L�x���FX��a�ח3+p�֩p���s'S��O�<�Gwp��#�u�u]�4���-�RN�5�Q �єxaY�N�z�X��Us\��mT�/�5iW�*s6`��7���W��D�=�x5^#�|�"�V"t	�����(q�Q`�{ �#�c����U��Z������r�ؖ�L�[��o�%��#(<��A̕r�Ȳ��on��Ui�Y�w�S�y�5�E[�T=�]��ww�҃\��P�%���m+��Mgne���T	���)P居�5ל��s���ei�"��;d��.�	]\�S{���K̮7mG�ܩx�n+Z*��a���z^\`�{��vY.e�d��!sy]���`�I�&������i�#���a}��.�F���׃Y]�YEd�*_�[⭡R��R������N�-^�
��,t$�0�8�炤έJ0:lr.�(iȜ���Z�	��Z/u���m�\J���O��q_������O6�:�^;��"Ɲ��õ¹��������xi�ډk�y��R(9�&�&{��ɮ���F���,rj�aV&���{�uj7x�u�n���%�:V:�U�W1,d���#7p`Ԓ�s�f�4%���,�cncx�*1����y�UP�&�nb��e#�$ᵙ���jYN��+���9��>�`�IR�b]��0����9Q��go'E�j�"a�LG
�V+O%�ͺ@xݾC�j��"A�du���[GY$׳��eI��t����o)��@q["�Ǖ��0_��x�le�\�����s�!�{0�mm=ݹ�j�]c�LHi��ÀY����T�Y�����K�i��g6&ᬺ9��uܳ���n>
�.I�Nm�Fq�R&��3�jL=ܶٲ�C]�ںAW��d�V;b�Ԯv�R�����_+�$[���r8�5��U+�+rG���EuʝR^�;�;(wegrM�SR�@����i#����F���g�A���ț�[7Fp��]��C.m�E+Dv��*�ok�w|��뻜7Ċ&CO�Ed���Iwn>,=���CD3Cb�t�gNn[vs���3
n�w�	2��,���Gv8��Y�Wn�_�qס|$^͠F.��0z�B��2��`Ȼ-�i`��;��*����Z�VU����ܤI�J)l���k+��x�<��Te�)�V5��;I1.�9L��]N�o$J����pj4.#�:^�v�7n�z�u�iUT�;�b>�j�io[����G�`<�##��Ⱥ�R������k�x�B�n��:�z��\*��)�/yV󎡊���ª�j�p͛P+02$m�R�W�c�N��`6�H��ڴ�C��6n�&$`�b>��TZa��; ����RY.�.���`��x�
�v#j��pbοmijܜ��!�k�<�W=��սW�1�r�*}���ۡ"�k�]�[Y��������̭��&�7�n�/t��9Rᷔ�Ë����Xagr��H���G��������Y�A�y��{Z*f��.1rw��!ƕ�w�7ը��3�ػ'S
��6;�Gj��Xd�|Vs�%D5���gUqw�7�,����/R�t�e�,��[���c�#]0!�Y��\���
�5�T�K�r�ҚP���\���kT��&�vF��34�Q!A8����<���3������9�E<&���Xo�)�\�*��Kۉr��	s'�\f��m�ދ��]�}���;m�.��!,�r��x�,���/kddA36�F4o���]�b"�̋�.5h����V�ۢ),�D�f1�h�c�Z��Ad����Z�¢r
K:��E�e[u%��>�۴Y����*^��#]��^k�@$����%�[u�sU�;sv����}-KN�tN���"q��ʾ/,���rRc����̭�1�F��:�H�r0�WPn�h��X3N%9��8p��l����בPwL��;t�5��4d䱗uJ���QFɴHO4sZ�J!�P�0N*ޏ���&:�e�<U����*�'i��g��L9��c�Gb�ӹ㹇�R.�d����CuvX�n��׉]$�{�|��G��Ҹ�A!mG�����k��6�4޻���Dof�k�*���p��2��֨Z���u�Q�h�r��z��SZ�W��Ve�V�{4^uK����,9��J:�۷!Y�e��K�ki?_ӊ��Y+��GH���'x%{�6�+8�hˋ4�(!��6���z+/�>{�Y���u��tx��QU}�D��Ol�5%d�����\� �w5���w�ݒ�<�z2��ʪ�b�~�]��MV����^`�"��fs�؆��Ē�uuʼ5��C�ك{��`a[��MɎ����t�`nP��a����ܪǝ7��S�Sq�fCO�Gw.��yo�:�"�ιh��$�!IIҎ+������!�,�F�{�Q�2%^9�O����]N�j�L����1Ʈ��AX��P^������Iu����N�WR���j�m(��ɺ���3���[+�L��ap:l��ww�=9X�/Gf���U�^��t7j�.�AK�,�wB�X�QČ�HmZ�D	��銌�[�*}Z�Z 70�;@����	6�p�(Z~n�UB��������P��Cz,��.L� �O1��v�y�mU�f��B��)=��U'f&�g;r�q��.��e�ѓks�;�}*Qە�T
�xv�#]9�N�r�AhLb�n��ˤ��JYrZ�4�'�{�es��3��pտ�a�[���س�W��{Qk8�ۻÊ�rH���9Eᣜ��mk[�ֺΛ�\�P�������,��Y����(�nh$���[��5�Y),�ʱ�����[эݡ6�Sە#�{�rо��zn WWF�^�ӗ�fAr�0k�X,샳L[�AH���ztk��]q�ܡ�[G4���-UC6�S%��wz��9Xm��4V_Q��Ž�P��H]ty�)Jx�[O+��&m!y�����v��}��ɸ�!�{���ؓ/��"�I�.������x�;;SyR׫1��,������u{е<�U�u�7�j��c��Tp���B���̮��G�A�5�:�	���f��F��)ok;���,��f�I�����	)�u7�"N��s�.���v�r�j���>�^�v�ͫT���St�8{o5�I��F	����#j���px"�,S�JT�7�7е3;;ێM��Hl�n�ݨ��R�p��_I�X�m�xݧl�9[�Aތ]��Yz����x�t�ꮙ)�&��F�c�u�Ty\7l:�,h]6��5�]���ΧZri�NZ8��0ٳ]Q�y�UV�\9�bl�Ι���V:�X�Qs��Q��� �&��`�%�]�gq88��]۱��GU��H���J�j�BgR���:���.��򋫁93z�K�:��K��v��]�J6ڣ���5�=�1��4��E�yՐ�xݛU'���\`<�����0�;ojŎW)͢��.ĒC�{��w��O),s�aY܂�w�������r��G��&�K�m�K�E��ڙ��r�B��8�N�c9&Ov��BT��d0Co_<��杜����)��<�Uw+QM=e�f���,֘�ǈ�9�뢳�!'ڕ܋���ͦ"	�y3���S��8���ٕ�OD�Hdj�n�Iq����ޘSt�wK���l�Gh߆���Q����=�Uɣr�J�����ג8=��jb2��J��6��یI!	��Ox��'[8�'oq�ɷ��I$��{�`���A�!�w����>V�7#�	��5�:CȼA'���Nu��'8���q��i�)���d@C���!�S�d�D�e����N����`o�-��PȧQ^"�	��s8�dK�qL�1�x�|���L��:���#��ٜb��������	�q,FE@:����s��� �+����f�'Sȧ1�1�p�9�\_#��7n��אּS����`'=`�z�M�N"�]Ay��A�W��N��.Dy���NgP<�����D~_Q�f�AC���ϫ߮A?�rzUDD��/�?h���?g�~�������UFm���G�]�kޣ؉�@�4���)P�E�Nwm��].yK���~n:�i�ܸ�7B�/��sC�����Pݔ=�������ԋo�Pm���t�b|�pN�M���*Rvn�ܼ�V��R
���R����5RC�C}+�Xժ�+�v*��BE�X6�gmi�
�w�hc�s`F�;�<�^��o�^Z���v�L�&���l; �y��UhO�؈�M�'`�V
%�5eΙ��������yY�G,�c����F�W��<�JuL͑�&USg(̡����{�H����Q�����5�^�����o#���Z!��סu��Ҫ��G��$�X�,��g`�l�]����]�7����VҙV��zY��p`�9n�e�qc��Җ�:��n��o`YC��f<&�(�{z��Vmo�4�0��O@�-�ww8����D�9���5!��j
�{r�l��f)#]�G�Ԅ4���*�7R�moa;n���j�T��X���盚(w����v�5oS
��-UX6(%�ERLNN��f�X��m�6h��m������#�. I�ln����9bo�i!}ҳ��;M�gCtq$�4��5��y'���jZ��W�6(ݖ���;�L�{������1S�vP5҉�p[\ft�d��W&xlz�����x���zzzkZֵ�kZƵ�kZ׶�kZֵ�kZֺkZֵ�k]5�kZ�ֱ�kZѭkXֵ�k�ZֻkZֵ�-k]5�kZ�ֵ��ֵ��ֵ�kZ�kZז��tֵ�k�Z�ֵ�k�F��kZ�ֵ�ZֺkZֵ�cZֵ�q�mֵ�ykZ�kZּ��tֵ�k^ZֺkZ�Zֵ�{tֵ�vֵ�xkZ�MkZּ��kZֵ�kXֵ��=;vֻkZֵ�zk\kZֵ�kZ5�kZֵ�ֵ�kZ֍kZַ���ƨ����V�f!�r���-�+p�����TN/
m��[iut�>�^�̊��	e�e�vF*��ͯ-�5㳫��ڣ\{;{"ܱR�d��}^ހH�mt���ay��K5���ONu]NKM1�Q�Ժ�ŐI4�&�x����7Ԭ;c�og;I y:d����*��P��}g���,e<x�ԋ��h�dn �9���=fQ�J�5[�ecα�n�$-U#YV��x�RG�A��T�&��f�j��y��7riw��@�YpBN�,��x0�X#��.����T�y�JF�pJk[m��$]*@� ��r�([��܆��}"')���t��|H�ћhU�O���OG	 �P��.����6+�T��r]�ݹ��5y�Z��a��f�U%8���[ǩ��m��bBx�#���c{ٻ�������F9"��fi��|�r�:�y����7�n񩌅��@	}ٲ�Ac|M*��ך7%�+a�Cx�p�'<�u��Y�֍	�Uut$�ew)��z���Q�{���u����,"�9eCZy�ŋ'ӎo2���s6�vL��`����dT",ۄ���"�;�0��Q�$zsp����}���A��-K�O��D��s�oo.ޞ��׆��k^ֵ�Zֵ�ykZ�kZּ��tֵ�kZִkZֵ�k�Xֵ�vֵ�xkXֵ�kZ�ѭkZֵ�hֵ�kZִkZֵ�k�Xֵ�kZ�׶��Zֵ�zk\kZֵ�-k]5�q�kZֽ4kZֵ�zk\kZֵ�-k]5�k���k^Z�5�kZֽ��kZֵ�kXֵ�vֵ�xhֵ�k�Z�Mֵ�k^��ֵ��ֵ�kֻt��ZѭkZֵ�kZֻkZּ5�kZ�ֵ��ֵ�Zֵ�-kZ�mkZ���=����<s*me��P����S�Ql�M�5jo13Vh�+e������ZK���<��Q�S6;'u�HN��V��r���ؾJ��Ps�/,uO^�͵rf��n�YO�R�hfShsw��;&Fܙ{��ئ���2M{� rI+/�h�.��l-�6��)HN�H��T��{ˣ��(������[�B��c�н�r[9A�0� �){����l�t�HX���źWb��vVfgjO^.Z��%�3�t�R�0P��� �=�u<�l�YTJ7H��EQ�/`���VZ�BwmRG^�0��
<�Z6-"M�pC����Y�<�ǥR��b>qUX��I�]P���D@V���\�z�*��]Ӵ�v���7�u[�{�m<(��$��������n����HzcG6M^�{�j&妪��X��o(i��rW�]��*\�o�K��WQ��o�!�:śD]��)��=דIё��(ӎ���M��/�݈�5[@�����wԎ��m�5�*�^/�]�\p+�[]Ϝ�e�v��VB�w?U3�͉���9�����c�f�\�s���9�&�أ��n�ǳ�,H ���}7B���\���#��d5;*=��żB�z�$u�R��T!��'4e^ի���ֳ��RN�5�/��/�]����r���2��hu1���vk�"a���e�G�&�<�����UMlɞ��̜��2:yt&Tt������	(�ד�A���w��8�@Tx���+z���6��wV�+��B�����LF0w�]�����$n�>���؋7P�G*w�tC�V����T|��\��7���V֭mH�Q�*���g��u75��#^��+���N�ҝ��^�2� �>=�%!׈͇mpTr:����{\�[�<%��y���R�/�kU�O�����<�|'b>�o��v'��e��l�S����J��+����C+zH��N�kM�	 ��a��Lq��>2
��fywl{�H�p�E��;b����V���ļ,�g �j��k�퐆p��m�o���0�z��熚"�ݍ��p8i婷B���&�UJ�F<єF�f��&�b5W�Lu�D�(���܋x\�Z�ӡsj�Ur���y6̳�X�ν��˞��ƕ�FFժ]OiN�]WmJ���#ǉ�ud�C�䖂:k�m��;�����#���zu�"sr���\*�<q����qx6�N�c���� ���Ҽu-'T�����������0#VOFOn��B����F��!s���z�z�.�U.�"q��bCkl*�]d��b��w��K�Ǒ�-�[���1�-�m���/*OR�E�3f;�v��L�i���JZ����3
�(t��[j����wR�WZzX�r��X1�1��ΡQ��r�<45��P�o�k���#���c�*�p��l�H��Wo8 ���v�ȷ_n���޽J�,𙧢���q{��j����Q�w���X5��������u�uU�̱*�vmZ������T�d��F˧
3+6�v�9�e�iWtw�*��fʑ2@w�v����K
���,��Ǥ�ؤ�/��֡=C��]��l�`�|0�7
��#|]e�0`�y���L�R!�q\�QZ)�K�s<]�9š��7�g:4{s��&�4�M=x��!n��C9"+tnM}֫"�;"�����5@�W��j�zS׵]ѵ�1��N$�����m�[]��Ԥ�D�c��k})"��\Zя�9EY�2ƛU8N]'fdB&Ԯ��>2����Se	�zm����+��)�Fd2����%����$�}[{4�c�7 ��l�ay�%�ԕ�Mm��յ��S�k���Q�tڼ�v�j�;�@�ot�$jN�y.'��+X�4~�3#`h`��	�P���"���{���KovK۷�N�t7q>�S�S�|N�2���U�g�E�%Y>㺣6����XO7�L����V!]�b��N�ݢ���o7c�<���U7���T�m���|uԱWe�G�k�q;�k�Qʹy��u@l8%m��ぇ� Q��;�;x��qr=;{�tT�K�u��)p�'��n�4u�o���I���ޛ�����/%at�z�ѦQ�'�j����J1vj�%&�EFu��;���g����2�0n�0e�i��h�Y��{��-]>pS�ك��r�n�1u1�M���[Km�k�k�ȑP�@��J��㡘<w`<�g6�p��0�ͥ��iU�uZ����ں֏G�C����)�K�qV������6�į64�Y�2�K��pۨ,�v�׊VVe*�S�8����/19Kfz�d���+�)�}|_*6�`��My�;s�A=�2Nw�
��d�X����c�/<�+��u1��2���|%���%|Wsf�{�B· ���i�i��K�"�m�Q��b�LG�$o�+�����%w0������n$�`�t���u�v���b@sdn5\l�cn��&l�r���hwM�;*11���U��r
8�G�B7���;X�����1݀���BL�'f�5w�^K�j�_InS0�[0:я�.�-V���w�`�[*�
��DX�+�{,5n�A[�J{�J�uGV�E�8�/���;B�^z��������|�p�[�o-�\�̪�rc�؊��eh��KF�kpMѻ�&�UI]m_)
-mޠf�y�\ɡ)Dㄞ٢�.���*oM\���P$c���7���_����n�IK�uM�7��2M��*<��;4̮�/A���JSF�YôH�tJB�8m:ֳ�kn��r0�-��ea�]o�!��u�i1��Y��$,�x���d��J|7Ҏ_fy��S*-�y�.��z��l"�lwv[bu�[��G@ج��W���ë��vWC,+�̭�ݛ��B%���2�.Wr�7%�Y�۹L_v����GU�\�H�6�[۪��!�ZN�F��pW���=7[�u�+��/�9����r�{�.�mV-I�]\�9c�s(;ٕ�-�]�>`:
� ��&�It���Rc�U�>���u��b^�%�����7ݵfV�V\]����K·qȓ��^���E�y���:�v�-=�����Oݏe1��W�<�¶�V��%��4�t���E�#�w�fT˪���&4Ek��pɑK\(Va�΍�_J�Ϣ���0������,pdZ,5�k7|¼=��Xئʶ�TU���]��ZS݊�7mh��l�ed'����.ܱv�:�8.;��ww°�m�U ��ǻ��&��uܱp;\�"`���6���)gUB�N�n^��(�U}��5M#�e�5Ʋ��G�wb'�1 �\�o����,z��c��H-��Th�<�GQ��W�ʹ��j��~�3��QTI���WR�Q���8Soc>�����j)6�F��0bf�k���q�4�4�@��K٪dY�8�GY��r.+���j���
�"7-\���t��)�i�rP��ų.��}��	����OC�h��8s\�r�z`�%p�t'm�w�j�M�͌��J�TPI��3��)n�r�Y�(0��%�"�D>�V-��k�s���E�s���њ����|��̵�2{l�=W\��t�S�8��e��c�yQ����2����o�E����[kK�䷖jC4u���|��q)����}KV7��'f?+q)e�5�U%:I�T��)R�#*:��\���F��.ʖ#�	�$�$��'�(�u��{%5��R�-7v��(�ă�����7)��u��Ħ�-��s@�Gz�p��r�<�.�����!׽|*�v>!��;��.S|鎸dZc�k'��u[����hZG2��3���B^�ct���/7*��j�V�Cё�򦦆*�%K���]K�6�.���a��U��x�Ю԰�똫!��/�3�rm8k�S�t�쇮��\S^�AVU�K`E�cS����5�;��)�`��2R�2��N���tH�����hn�L�Q����0nk��N���qH�3]��!����j7̼��K�����^��(������j�+}ݶ��A`�@l�o�dgY)P�9
d���n5Zœ�e(�N!��.��K�j�R����:Ln���PUK�=�2=F0zs�z)��N�d���3H�l���v��#��.��3�d4RR�d�8���Y峸{ӮT��3�eD2�l�2t�uE�]Fe[�h�>g�
��J���f��J�lmgM��X�i�0̱��056��(K%49�7�iչ�s�6�P��WK,ܴRʽA��ҝk�JH��{q�e�6N��˜��7w86�z�����:�KII�ȬV���W9�o�����z6-�.����^]�����@���N��Q�uVfp�Ʋ��r���r�H���==�@S��J$3Nh��5��J.w� ���w�<�UtL�hae�h;�~oW5o
���#��1�>u	�viZPu���Ŷ5o��YvM��������tڹ :w]�ழ��x[�:ۼ�r�ݝ,�aN�ge� i�5S38��q�97 ��.�'��^u�s#�-�$��O������0�53M�C� ���e��� �ٛ��bO`J��<�LS =��I�e����1!՛ES�j!��;���Tr��<�Y�N�$P�B���e���۳32�^=@���Ѹ]:/�Q��]�Y� 춨���4{~�!]l{p*�i9ӀSa��X�ј�ϣ�Ъ����0u�[�u�.*]f�����^�k��G7,(ug*�*���Q]��И�8����z���f�X�U�!��'�K�+�d
k��v;+��N�u��KQe��U�`گ#�����׽R��2K#(Y%S�;JQ���<�_%�Ȧ����vrѩ���0�	O:=9�la!��G\ֽ�x��{��󀽍��!�,�ݭ��EE��ރ&�}ö�L��4ָ�s��1S�|5ێ��B�ch�	x.������� �ɐ������?���5� ~�zH ����$�_���JF���T�7H�"1(ܣ�w����^=]d��;�|xH�h0�A�[-����N�B
a�4�?�e"�	r�)�$I��O� �L��q��
�FB�qlYH8�(�a2Q-�5E$��S�"$E�m�r��F�R �
F%S.��dMm�7��W93�SE�چ.!��)&ؑCf���cA�-���JM"Ӧ
��T�Tila�X	2�e"$!!Q�I�4�J ������ ���-�B�ɎDK�^���w���u$�!�@�$���Z޼�p�����M9!�c$�����c�\��Ւ��y�ʹxV�+B�UZZ�F#s�V���w�qoY� �f3�.��F<�6��F��=K�2\���(���S/e��}���'�Mo=m湗31<�|4���͉ܳj:�c���6$N���-ˮY�UrT�B�_u�o-u ����΢��*�Z ��1re���E�����%��n��}#�VA�a�����ݜE�J��7D��	mm���HJW��fC�7�
�;���Ã��5�	�qn�.D(�����-�����R������rZɻ�r.��n�)�5��yRX6IB��AAݹ&+�A
����x$��tfӃU9�Iޕ"�.9e�őS��/qw]Laxr�nըqުK&���M�i���>��'Q��%O��vbom����������ɗ��m��@�q	)+��ӷ���v��:<�W-Qi.,��-Μ�7��OJHm�0��}��X���$�h�������#�Y������Fm틵�,��Vpn`�e�&_G��w�߱�E�Ñ�KM[�]��r�/]\�t�F)�m< ۤ�P �ᐖ�l�&R�M�r@@@�YR5d���e�&��H��&����b81��LJ�]��>���)���z^͢�9إ
-����-�%r����S4�< �T&DYP�
l��T��"�0��!@S|e��j�%D¾9����כ��*^oDE�{w���"����FQ0�-�X��$����㸡ox���ڸໟu��sGY���wD��y�w{��������%.�N6c�0�< �L�a�8O���fGI�Z(%q���&	q��F�ff �R@����0��4a�R%
���z;��x-�>ϻ�޹�",r�8��H�a�2��6L	��
Ai�Ȍ��M���T����B�l9$(B\�&KFq�[eHZ	��@K(F�-�
e(��&1����$*�q>F�K�z���w�ǹ��t��wQ�QqDZ(��L��*F�-`O�w�s�=���H�1��a�Q��i���L�G
.G�J���s�$预Oq�N��ֽ5�kZֵ�{hֵ�v�۷mx���I&!��*�)0����[0�VAɚR��n�8��8�tk�8�oooomzkXֵ�kZ�ѭkZ�۷n���$��2p�a1T�X�����k�=�r��
*�^�y�ܱ9j�Ҫ%�Q�3��E^{'3-��<��]A=��fr�-S��n��aT�"ZVau,�����"��ZJ2B1=Т�3s�r��9K[��L��Z�!	����A
�CH�i�kYaQdT�Y�9]$"�����
��|�k��+,�֜QKi�B�$�U�Ε���t�Nn���{��"';���Z�i���܊( R��O>n����i���µ��>p�߅ܕe��g�K�t7\�+��B>���YUHV�h��::�"��O;�^w�g��={�׹%n9;�Q;��Ͻ@Zw^�^�UM]w��^�=�Ww��"�GN��\4B�f�z��u�L��O�s4���hx�BB��wq�I1�NI���U�+�v��yy9{�em���+�0B�h`��4�) P$�B�Ơ�q��Q�d��!@�#lƚ���י���w/��K����=�Xd͏���+������k�����z��wXs��j$�˩4�[	Ba�@��Â(�!m�`�ۀ�! 2c@�S�HI(Ƹ�nNE�P�DD#0TR&x�i�[��p�b���Ja�ʎ�8xx��f�KV*�Z�Q�T��O�|RY@�v�kMZ��w�<�
���Z�I��zTޅ{����^\�B��Ej�O�6�<�#:�ޜ�B��`
�����Tu*F���F�Ϳ�Z�~?E�}�5�R_G}���ݦ�J� ����Ne�N|7�Zb\˓�&nqVW_���_@���������0���}��Z6p�ն4pҽ�cKd6N�T�7ۂA������ ����EC2V/�.�\����o�0�M�`6B�E��@��e�A\еֽ�����Y{d	یB�y�m���[I8�o��)g�l>`�t���,��9u���g��>e��T�L�W���U�>W�
gM�S�a�Q!l��X;��L)�Sjb��2s^أ$��H��
��˷|u��Q�g�̼:]��kQ�@o�0.����q� Nʜ����z��1�3�cwECB֛S��Be�"ɼ�2�sqs��m~g��O�J��6�.eg�[2�m�6ކB:/���S�rH���Y��6��:s�ɷG]�����B�������c�l��k`���Tл��]�.n�5ٺ:E�ML+3�v��I77���y�(2��f�����Y� P�)�k�i���e�%�Iݤ0��K�d���^�@С��#���J�U�`역*�}�5�b*4���`� 6i�+�8$Ic�q���� b�L��N�y���=y�/�f\���bT�D�BuW���Z��o������I�T侒�i#J�v�pn`L�����HT�g�7~z|{S/H�SL,�^��²ul[���@��d�Sl7UGPS]�ߏ����������}��ni�/�3�E�X���"ޖHl �u��,�J�XV�O�Nٴ4�N��V�72v�@�g��
���YrDk�(ց��pξj'I�ѮsF�)l�g��,9�!��Io�U�	�ݜ�a�`��MUy�;��7d�~c(����yH�vA5��!�v�߶[��܂��kj)f��ܗu��<����Њ�1�v֮�e��N�T:x�3�ij�dƯ�a��6��`���&�.���ը���������zH8\ܗ�����8�s���Ð}�j][yͩ-Iײ�����ɇw7����I:������z>��Pg½l��6v	���&F$�!k��o�ma(�t�ey+���w8������ąx�R�%fKj�|Q�w"���=�W;epxf�;����o<u]�o��	�ʎv/�S��8R߽K��ycl�o�m�z�Ϲ�1S�}�hɥo2�6�$e�n����<V��*�[�[AG��t���e�.s�T��8H�r�Va�LW�׊��uP�?�(�R�rUuV/ʘ��.o7����"�y≡�طv�ƍ���#su�U�j�G�UёYһ��D>�,{�@)指�&ײ���NB=��c�mZ$e2�Y�)��fP�l�g�w��E���k�t�.Of�΍��q����sVN%�xgB�VN�~��A*���@)��9Җ��}��ڇ�_.iWf��9[��*��2z�px[�rP�f9dv1	1�r���{�v��U��EL���zn��H�VǠ�/&�s:�����ayW�V�#���kd���&��n�Po�,���9s�d�q��I$��M{��۬H��xs�����-{�YAT6��c�{�}��V�{��VJGԌ��s�F.�%�M2(��[��Kl�X\J�QZ����<ڒ�P���IU:���{m�S�
]���h7�qZ�8�(�2�u�Z�&��
AD���pcuLR��9:����3K� ���$pB=O{�ۇ��:��T\��N��N�!^R՛�M!�2�{kW��)ڜHW}]m�Q��m�a	���z�#������ϳiY��D�$جOF�U}�y�^�d�Y�>w��H����s�����׺��Q���F�_�����Kkooe*��(�戕cՒu�a:��� �!;k'i� �:�#$k×�y��E>V#c�u�X�]�J^�-�{��vs�{z�+�@�9��\Z�dإ����6�Y�s>�p����iNo[��|��O.8YVK�P�Q.����.fA���i@w��6Z��tʑ���SJ�Vᾩ��Y�{|�rTݽ̊��L^qwO�2���8#��3�D�K�h��x{1�j�­�Ige��OR����P'{�+i�uV5*EQ.�lף���з�0F�<42�����I�`��`H%�~���n�q�ک�Ճ�S;I�4�q:�:���0_R��^�s��dj�S�
��ϲe�e]��:�$�@jB%�_dX^У�ȴ�D��#�R���I�3��.��F=����*�)	�Z6)�!�
����ۜ��26�99�r`�Ub�=~�5=��ׯHM�JBF�VnH�k��5�l+取�����u����>��ϣ$�2��4*�u)��P��n�>�R۱�qS�����XY�5��J"����]-ĝ+X�T�M�̨�%a�զp�Wr2�4���#s䶌�fw�7�|{Tܛ��N�Ź���K��qx��Z����j�S���ΖH�
i�(-ob�V�Gb��KwNӢem(����ĊR��;K�CB�|�x�'�uX+�t$��+%�ܫ-F1�r�>�&n�����)�S�����	��H�9=���>��h�zg$/ �;��N��s^䃤:F���gP��`�|��LC�;8�l��Ʊ�n�V,���������/)�������jt�Toҫ�i���2�$_�F$��'�/̜�e��V6�Ͳ��Q=�j��6[x���H
�Ą�eG�d����Dˬ��>�����I$���$2=��� �u�!c�Զ�&�L�-_=P���k��
��W�d,��
#D� �L|�X(ʐ��;E���̱�p��o��}�|��sMo=��*c<�0�f}�W2)l��F�ը�'L�QE��۝��vv�ǭ���מ�̛I s!_l���w�a=����d�b��׳+���|�}��釘u9���t�A詇�Ӛު�y��(f��+)k��ȥPq�h�iZi��Q���}�2��R�ZB�
�!#y�P^�S�C��۽Ŕ��F�`�8�
z@z�TL�lW����L��(�{�����6X*�-it����pM���sfM�Շ4�̵m��UqҊg�Ԕ�U�E�t�Ř�������y�f`F��V����p��Z������Z�\������.��"q������&[�[�QeuZ��\.������
����wn�j��Q����1���T�c�Q�n�ǌ/4�0m]��<�f��Ƣo$f�L�M 3���7�iQ��ޙn��m2�!�d`�.�T�����+Vݣ[���gׁz5�-a*	J��8J��ۗV4��lgt&w�r�jmn�b:e�t/�K��$Υa�*�eIGdFC[T���̩2U�d��*��b���+�?k��K߫;��{v�l��v�x��w6խӒV���A�����e�`|�'������[��?(E�ӡ)M����J�鳥��1������Zj#xDT�ځ���a�w�r>i�6o�t�R��>��s>�2�L.��^u^����L-���	x�,k�m��|�4S1^�3jߪ�����ZKW���V���|�J���K`-z.|vb�;\�Mͻk�vW�TΗS�m�nt�r�U��}W�CwYҰ^N�Ⱥ�%�,\��Gm�۠��"��[G}�ړw�Q�v���m^���;����&��uE)�ټ�w�^l����.F;0Z���(op��w����gCP��P���e^CݎM=�i��ɲR��L�"�~���}W�o-�z]�~�z,�(���y�h\���^Fa%!�ی谗���Ż�Ag/��|��*)�
�b�j�^^"�(�������X�\�H��BA$G�)N� �l��4��R:<A켐��rn��%����R�҅>H�H;p�^��#E�aTP��Xm��t�i�Zt�M��0�XJR)����&�<���n�}o0_�E��/E���
Z�s��(e���Ey$e��+m���Ylݑ{8����Z޷w�L���Ð�k����݄���J�}`���f�_kM�������u����퇣�R���c.w¦�^��nV�Ԓ;Vt��m��>ěQ���?�\
��-�!l
5��U�b����w���\����ɪ
=�ͪ4۽���-��Aen��!&�����T65��:k�p^��V��z��7�e�"���[���lͤξ��e�UR�N:���Ύ�ۍ4oJ�5�Ƙ,�7���"5������*�	gL��V�Z9�&��q�#O^���/8u�Gde�7I[�⼔;�oEǁ�Gc��Q)�z��HWHג&F$�=!CW�m�ͬ�l�ӈ���FRX��Z^5z
��Vz����T������%U6z��<���������U�i��6 �ȊP���Ӟ'V�Dҍõ�-����l1}���s4�� ��k�6�N�r��/����'Ű��+S��Ui�mp^ї��`ʑ2�߀�xqCȫ�(}�A2#{�Z�f�0hXeKN�[��aU����X�؁p0Yg��y�j��Vt�~�y����$�G��5Iu��V���Xd@Y���S�I��h��[VQ�6���U^<�i��7�8!������Cr��RJ�ڪ����S�K�g�
�*� �k� ^ߒ�$%[JR6וu�m�>S!uuNN���'��A&d�����^WgR�0���2�UlV:�Ѓ ��
�0�\Z�7f�����հ��Y+�	Ns�.^�Vq���ٶI�7J�`�Nz��;9oj�B�CϽlqu:��z�qy�"�r��S�^M�\���aʝ��s]�V&q���o�H��I�ov�@;����&^u�L}�?�8�ãg��_u}��Kex���0�L���MNqdm(H�*]�V�ﬓ�������o�9Y�f�a-#�oI5�I9U�)�c��Ғ��;!��fz� �%� �t�$EV�U来����H�)6ʴo�^w� �^қ�/�d��R�:u���\
�26��gb|Nz��	#mOUM����O'/��g��_/�`P�@9~�3�h� Ky�+���D�XKًрeCY[��:��!@�o�nz"��ʑ�� n���	Q���ټ���X�t�^�e V0`�k�A�q�<��k�-�ed�8��j'v�JLsI�Ҋ�'g�ہ�3�s�bl���7y�7
����j:cyP#8a����ڿn�����٣��GG�����#�
l�5�&����3��W������KX+:=p��v*X���˛�Ӄ=�� �����*iF�� �t��$��)����tH�].�S�L�Wƞ�P����佥f#��Rʱ���mr��1:yʗ�3�Z#��(���Y�F���2����
��%�ũj�� {O.��R/!�+yq�φ�hf�Ѳ�7��Gi��h��`�K1����T11�³�#�YmJ�Y4�$�>9 r�EUm�Q]L/��0�wwtlTl+�^x�r\:�֖�V_G٧�
�^�{<��ٴ�Mк�%:���K���U,�N��7Xۉ�\�1N�(cWE����X����OI��0��v�8;2]*�r�vJmi���4�W(�]Իc�K���"5n^�;�+6�D�w�@*�L����j��8�7D��c��ٽ\�֣�3/��!"���bܠ��PP�6�٠U�]�t'Vo	ZMk�^R��V�c�͗�:�`뚓�%%;��f�j��ugr���>y4��N����#/�X2�	)kP�=p����R{��������������ś����}v�82޼�cC�,�yn�e��h )�kp,�E�c5ӫ�<���`�+w������QL�u��c��=��3�r^��ݔګ��5�W7��ۣwܲ��O��h��m�UE���Z髃s�4d��"�=�A1u��MؤB˰�K!�$=���Q�I~�^��k�~����HD;�*��]NG-�j��ЛZ�+���V���7ʸc�$8��T㧻m憑�x�b�;Z�����Z���.�1����U�����G���^�y��8�k��u2�J㧔-�|\��T��W�	��$b�&���K�ԁ�JS�.���^ӮVc��VA��;�-�uo���MU�Yj@�^u�K���oe^��m��p���������֙=��Y̧��߂Ƃ{G_��AÎ�-�J��ev���r"��v��;*P-꼜2O�<J:�Rn�%�fP7�D\��򥐛�&A3&6����c��{�g �t�r��0��VgFkZ�qA܄�*�>JY���T7�.�&���
Ԗ��Pؾ�<��AD���T�iY�e\6�E�t:٫�d��f��P�u9�~]��R.XgYe�k��u��7d91n����J4�j�;�����SSlǮ���щ�n��%���Zt�%˶�V]��0�3|�ۺb��W�+-{w�r�B�(�3Ĉm7
���}�c��,��.�ѯf�=]��E�3I:�
�om���H�u�-.��y&g7�3�zR��h9�����z�v���N�h"n��a�GS�\\�&лL�A*������J�G�+X��P@���{��x9C��o"�̻χ�W/����]���1�I^�{�x������]��������'�f����sd�r�ۧOO�Ƿ����������Ƶ�MֵӧN��ǮgFd����2LAؕ��zS".�t�u�D<݃�����uő���������\�M�Ir��0��i�Hwrp�dNB݇fa!��lt���������Z������������kZ�N�:k��âMkS����������s+ݷr�L���t,TK)��h��2����w=F��+�+�)]N
{�n�;�)�#�$�o������b����n�y�=�p�{�q��G�qݲ[��I�}�����IQX�9��xw^��(���D��7!p��	ރ����]h�N��[��K��uGZ���*�e<�{{�5a�$��sįuبEb�y���2�\�:TU���w\�-r}��S�A����;��	����u"�W(�TY��u,(�y� �IU!�r���A����A��{�$�P�;�p�r�eUG,ʪ���"�zޛ�iH[�\��\���Mk*�K̵�(�W�ݡʧ�
��n�ȋ�\�����*|��i��W�qұ��	y�A��;�W�#ԮTW�,,ԡgI�1�72q��%_w!3�Kκ�wH�I.���&�C��Z|�m�,�{��p�ݧ�,�E\�-a���G;��2�g3�=�a=��"Αq�	E�m��q���=^q���x;�էv�!�}*bdC�j��t�Ւ;&�;_�a'��x"����[��W�"���g���ƞnS�g�a% �7`��}����Տ=�>]�Њ��
�]w���N�/b��5t=��`�nyx������U�҇�g(�����/�����ac���|z���Fg�}B��������w�[7d��u�=��s(/�}1��Y��E�y����̓��o�k�	UϜo!<�ޅ#c!���=�Q����E� ���y��-��1���O	��n��:;͔�����܁�kC����W/<����9n�=���[�G⻢[���zi�	�U�q�-L���{w��P��1�C�{2/��gb�'���`�8�~��7�lu>�1�w=�[�~��7�]��V��Iȸ~��c�h0��Ir�jܣ�xy
>�m=r�ן?Tk nI�	�]�:�K2�c"�t����N�����"���^og5g=S;;3�X��y�.R�z{Q�=���W��3�r�/�E��4���O,��!����,��\=�v��*%�þ��=��|�k;!�8vv�u&%��:���G���K�5x+�98��#d��{�Q���4���،'D/o;r.5{�J�ة �f��S�z�*���'3�@��v�^�т=��b|�v�噹',r�v�v-��Y�ޕ���\��T9�Z7,Y��N�Ty//8�����{Y�E$�/�.z�v3���l�/�@����1Q>�:�!�x h�A���Yټ=���n����v8�UG��A��4����N<����}���t�9�mi�;hzS�K�
���3<����zG/��^��>O7���-N�h�u�z6�K�J;8�ɍ����|��Ź����O��?���q��Kx/$�hk�QiNm�POa�b��h.�<L�'(!��?� gh��z��u~��v@lst������;?�6�� �'N��6Y�e|i��fD�����p-�ʑ.�������_�p/���ί#�wF�n�O�uI�ٲ��0O��-�8����o��Dg���\�KO��r�c�1'>�|Wܞ)�������Ζ�7�{�դ�|�kQ���A���x0;���ٶ�,o1?�*H�v�(�ڢ�����Q����Nm����)��(������t8�%���U���2/����lx38��/���z���'erYg���8������ֻc�n�IG�����}��0�����T\>��y׈�=���y\�.{���I�Ǉ$�`/��ͦ����bϲ���u��[<�b?'�����wZIv�\�4;�v�+���VWY_!		i��+�WG�5Bot����2l��L����t�j��0%zu��J�	��×�+������?���F*��j�zۼ�ר��/D�� "�7W�?�de�|��d]L.{P�r@�-@>ƲO~u��ܨO4t�?�鸷�Z"o��d�ܣZP����8�7�50����gd���6�H&z@�\����/�dxL� yۗ]���Ӽ<S���Ч���br�#<����2�}1�>���7�m�7H6o�-K�Ԙ)Ɍۮ�$���okjye������#94�F'\� z�H
,|�kA�U����jdԾU�����G�<db�kXR�%�˞��2��v<;�������I�5�&J�\�����)�^S�zvF�����ؗ\���%���[�B{mi�zw�wgNY	��T-�w8�A��`���8��_�[���Ek�� x�$g�߻�'����i����i1�M:�S4R���<P�b�`0!Ǚ�� >'���PXsg�;���Nf��(�ܲ���{]Z���v��[q��>����B���o-m�O�+<�7}���%�g@�zՑ�'V�oJI;�fX��zD��@ʌ;[By/.�8t���S�g��;?{�,#�k����v���2v�x��r�Cf��$�2���wL�"\m���-{$�DjWW�yq�7e<��u�ڢKfCC.����T4�ڨ��m�BP��[��;�z㡂ʝ5V�(gY;{��[��jn�_���������5/��� ����2A�z%G�;J���x����3��ϴ� ���gQ�ڞ��$;l�qL�2w
N������^�����/`���G�y�\n?5���y/,�r�DC�K�#n*�A�����p�
��hyh@��y3��_ ���>��n�����X��ٳ���1��z�4��E3�3�aA`&At���:6���O5����
紫�75bv�Y�ʷN����n�W��[1�cռ55���Sjq-s耔�ç�6�F��Bm��sKz���n�q���Ⱦ'�Ja�B9��W����uY__M7_���
�;�}fl/u�����:xz�T�Hj��f������d�� ���-��8�7R�a^s��ϸ�qn�Û��0���Z��"�����p�k�y#�nI�%�?0��������r�S�t����S]v�ښw��P1��O!��B*���龑<rzQ��%��-~�{�%C�O���_!G+��z�:�ۺ���xyC�9��a�s��ȍ�8Ѧ��,NwP����T�v�7I��K�uyY�r����	�%��-��*0�q��T�w2��;2Q�x�$�o�c��"�&IHu�bŜf�K���<���g��W�O����΅5K�v�scW�}���������o0�7��+�vRѼ&���zڎw,���x�x���{{������r �n�9φ����&4=,��� �է�"�: Cu��OOVf��7�]���.W����jؿe����e��!n�A�9���P�W��FOqK�Gꮺ̿V�f*<t����=����mJ=�䠲�icHw�`�Ѭ'�Hz�$p� ���O|�x��ï�w=DqeL��YY�<����7A���m���i ��;��ܽ��ǠH�I?�+���?��[�)1���!�L���"nR{��7*��l�r����\G' Jx�ɰS�F�P�9��j��tj�Cɀ�_x0���Lt��
U����B��n�	����p�ҝ��ٔ�*�w���S�������n4��x���gtq|��Ǡ��p)�gwP����4m�q4�Wp��Niݾ����Y���ef�����N�lo� �q�����-�#��5��O11%ݭ��I���Y�W�Ql��Mez%�ѣ�N�����^0/�b%|>b��H�x2����V��.b%�'
X�kъ����ps�J ��~�[�����U�q���"����	_��߉���e�"���dy��d��8�A?q�9����՘�7z��*����d�o^tR����=��*�[��ظ���UAUg��T�s8ӢP����\����̶�le�:�f�{�"�۾�8M�i�kN�Y�Եe��ѫ����?�y2q,���M������@�_\�7s�x���ɽ�wO5���ȸ~��jA�P�m�z��������E���,�B�T�l�¡� pqz����aG5u�/�.�`�
*����>Lu�^��'��a��>=0�\{��#�j`��̑)�U��N�������=�������ۼ;��<S�n�\�:�2�g��|�g�sXd~՞��m�ή�_]\����׹ǭ,U���V'�̓O�W��U���I�VQ������(ɟ	��V�6��F�7��<�&<=�t����������r<�1�λHa ���\]�x�7�9>�Gl֒��'vvg^���~����N�l�Hj���� ��<v/k	ݠn'�v^�m�[9����`�b%�L:lנ%�8"Ԍ���pm9�`�p�)�-���H^��r;����w��x$�p�_�e>a���Z؇��f@q07/�3�	�Oiٓ/�]җB�b����8o��T9�VV��"O��P-�?�T�/X��.�h:��/�Wʜ{���<5�����L������J�cz�ޡ���³�)Z+츟
���|>;�%��[��C����.$O�/x�\W؋�.:����e>Νҵi�P;=���!0��u����ZC�t�(�dc]���
p��{r|8x�����>�����p��6�ߣ��I3G!�WuUU��*X�~l�@�hb�툁<��Y�)��s�N&�>	����[rx���2�4*A�
��xy��xy47i�/�W�CsP]s���!��m��`����N'���o{Ilrg�!�NF(y4C�7	�� �)�:�a8sy��7Wr�gNm�*a��g�ҁ��ט �ȹ�Q�t����p"'�"��ؾ2|�'�"ƃ������+�	G7g*�Ӕ���Ƃk;;��+ t���e����-����稧��4Boq�t��&:�m�qͬ ��=�Q<�}ʇYO�Gzvb*�dGj����̟�^�;2|6ab�����#^�Q�CN�Lt����+K��Ea��g�����g��p���Es�IW�y�Qzw�vD�>d,8��.�<5��ʒ�БB�엘��Y�3xy�n�U<^��K���b ��ɤw��Ui�p��;�F��>�^^��dY�1��3)m�Oo|9=��(QM��N	u��|EP�1���=�c�*��v�p!�n>z��Ƒ��˷\�q��f�A���-�^��_����NIN.��L;#�Ku���|����=��zOÿmb���̚���Y����.Q��%��ݳV���z����kxV�2��(d��x��꿖١��3�/��4��I���i�ݜ�z�"�i�3����r�
��q�sfG[kEu�w����fo��9��'|�N�k�v���t���Ւgwo&�w�����ǆ2�x����{Г�XP[��g.fg��u��'p����[p/n��0��w���%��9טvn�)���wP)�N<��<����Uqk//-t�mp����[#�0/����:���<%��)�-�
]���y������7ؗ����^O�B������C2נ�Z"�i�l����T?�����1���M�3��=J�W�s�ǆ5�e�?��<�C|��7�<����D�C��d׶<���='��ަ׻�x��͝(y����ʢ�R��.��/jg�����'��#��>`)�f.+�!1��ݝ�*�����"1�����ND���غ[�t����wR�Yc��g��*��>Ô�P��}1P�F)���څ�4È.��}0��6|�%	������isB�["j�����������+�ڮ��B�P��|xY�|���8�JzB�0h��ֻ&��U�]x����Q��ݡ�\.��I`���^�.���'��-RN,���䲄h��Ȍ����$2�/�ӆ��Ƙ��Z���S���3#��w�v�����r'��v���,ע+����ǻC5��n�Z"��U���d۽g��(��67o�y�6��͡�	�;�%��'U�,.�x��ǂ�U��JW���*m���q��:f�	I<���^�t��Iøw3�p.����~�S��~��幽��y�1޵�����wf:ے\F<9[j��ML����ާ�����:���ʧ��y����6�J�j��!s��ȗ���f��������ˀ��a��ŕznG1�b�<�zhY�e�(�r���L���a��k�{��QÐN�<��vܴ{�ű��B!�C�?C�����:]63w�)p(vF���<ft0�Ʃ�?���M������*fC=���5���`;z �-#`#_�?j����~�J�
8y]�%�浭�O��^�v�C��O����]+[z�<��!v�A��'��(ݵ��l�x�LFuof����Ѹxx˖=����t���k�(4�
�Q�ΰOh���%�?���6�ϻ�R��|�s������.�
�ԩy�@�t1��9���顶/�<D��O|9����F�F����t�3�M���C�9�z�|��
��W2pk�B3�~��-@���NҟE��t�ƎBQNo0�YϽ���kU���Ha����|~� �o[J��绥B7a0K�B+^NSV�eY������c�{�!��Ⳋ��]�������pB+FQٻ���;��[���46(�B,���GRdgv
��[��5gF��\]u^���H�bu��ua+{_It�6�fQ�5�ݪ�d�Y�K���=�1U�������vwnq���]��츑$	FFFF�I"7�����]y���n�1>1�=nyP�����-������s�9|�������������]����9��Jr�����o�zo�:>$>�Ч�Z�b�9i��׋ǩɼ������0g�%B@ֻ��sU�O=w_�8)�z��7��ʝ�_>1P�c0��5=-�)k{������y0�~����kZ�aqA(��~�܄�P��{�߲�{x�{w�c�ѽB�a��ۗ��:P��<s�0��8I��]��w:}����LR��lgV�T{Y��Lmn�V��N�e��@��"�a�e#n]�O�#�e�]]����]����=�/|��7̋��wV����L���[w�F�K��
>5��/��A�c˶hx�����/H����<BW[��6xx����sb�'��R�o\:��l p1��p����$���۔3s:l�S�eb'O%�']k�r)z	A/E�Y�$M'�VQ�1�B�Tk㧞̚�w���J�+��L&\�q�6KW+�W�͛��W���;�k���] �ppp Vn��-�16�����fv4vލo��c���oP��;���6-�}�i�齂��Ϫ���6%ȱ}~����n�;��Nt�=�J����
�/fk���+\vIV��v|���k��O������9�3;/@�nYSH��ڂ�0����{�Jr���.�C�d����k-y&oE���"q�\��/ABf-\��St7:�{�.�s��s;�'/�4������V�M�i��btM̰/��[(0dL��� g��)k����68O��o4�̥BoE�E�VJ�W�
-�	��{8ո�;Y��T���K�pP�����9X]��Ă�G՘��
�/���]�7'^Q�pɗw/��ʟY��� �ͥշ:U���L��3R�	`�Cs�٧\;����]�q%�
7E\02ܮ���୙�M�.�[׼;��1[��)`�+��-��|0u�^C�ޗC��o;�V)0�j�ٙ�搞҉�'�B�nM(R�nb��nhKeQ���Va��]+��O�����8�kѩi�s�	����|�B��&��'c�}��m�h��dge�y�ͷ:��Я4Z���Wǎk:�nE�d�ӇJ�]E��+��;��/5��b�iYe�2��P��Vm���*��w<����hu�2�	5Z�&+(�[:�,1,Vh�9mfg����\��18��Y�WS3kO�q�u�Ӄs`���UWi�{Jȥ�j�>���df�n^I�c��%�Џt��RPD�����},LW:�6m��ڻ@׹QǓ'}ﳦIrIP]�U3�`2�Y\��G�R����;e����
r�N�gow��3�z%�όnӲy-7�[�t�n��	ܗ���q��9ƛ�iBq���Q)d5��e*�]�mK1�����㣎�4��6m�Q&�Wr�&�S�Y��R�W3r\�h�u���vq������ZW�E̽���q��r�As�][�liY]{����uρŧ,������h�p�x�X��+��bmZ�k�+�^��R�Y��"�-qsT�N��%^X�/�k}�)�M<�n�e9�γ�:�{�v����U� R�3Ҕ�3���Z�67��@Q�ʮ'7�z��;�N�tѶ���@���nLy(Zh��U:㭎ͅ�)���[6�,7[D����E��o�b��х��p��8Ϫ�˫w���S�����Y;s_e\*2�[^f�%�^�J�O�l i��=L�_>�uq	x�sܳj<0iw��GՆj�Y��z�&�Y�U�����=ު]�5�wJ���ѡҥ��ͭ{�=����%��Mt��3�jG�����ܛ7-�]K�,�o2��Ԉ�<�e�����r�*s����Եv,X����f��qϧ�9̌��L$a�"��2��G��Q%�t�(��
��\@��̙�I�t�����kZ�k_�����N�:|k��X`ɓY\.��|z�u�W+;y�^v��\��$��\���#���<;{{{||xkZ�MkZּ��||||xt�����R	��2a���HёY�h	|a�$G-C0��N�t*���ٓK�?v!U�E9���t2Q)@�9�h�����K�`r�"IQUO]��49.�T\t��)V$ir����E�ܜ�
	@����me��7\t�<� 倴�Us�9NSQ.�uVf'B*Ғ�
�QW"8QTW9|�^eETd��iX�s�
�ZUE&\"�O����;�HY��,��9�QDL���VW!1P�}'��!"�8�Es��*<�Eu�IR|�i��wVP���e�\�R(��}m�H�L�����A71�,.�"���/G �'5-�HK�UEȤÃ���(�DR�.Z$Qdd����gP�#���U*U�E4�˾R���b~�$��n�t��4XmBX���0Ӆ�q�[�&6Zd�ሂ�a�2@�Ջ���ׯ��N�J��k�� 3�� '�rT���u�&�3�L&�Ar�$���hl�溗Gr���}A�7)L4`Q�,�-���H�q��W������M�/�����ϫ���P���Q��H�#�E"a�D��1��(ٌ�X�_ ��5�����/{ׯY;ךՅ�P�E+�R�^�I�c*��z�ĥ;��P�q�}�.�a*s��?��ujxbٞ�)P1%��xo���(��F2;�kH�(L0W7�`��t�Q'�a;�ɛ�� �D�Y���d�^ڑ��=��9�aI��L�^C�����܋��xϝ�鵨;�+�-Y�?����8��nNZ�D���0�;	�ｻ{<N�jvmn�9�H:"�P�e}gI�e������MQ�u����t|�÷�����^��������0]|�t'���)����KO��
X<�$d0����;�+7�F���yW��!��{b�}>��6�U�ɨ.���ܤ4�Ͱ@��~r��a8n���8.-5lN���!�ϸ	�okl*2*���1���_�{���]ʱ�9�똨u4��wB�L�|���H������� �la.�[�T<'Mlg��s� ̆��p�su|�WGH	��(���hk�ۻ5�eJ,�=mKpU#B����?� <������;s�Z��s ��u������V�=WI���Q ���)�-�2ޚ7�g�!�?t�ht}�rX
�`�`���{*y���ڕ��2�W�tQYB�1JB�M�4^e��sO�rS��\��0�
0�����Е��'��^�>��Z�jk�m��E�٥i�R��0�P���O�J��x��-��ӻӈ����v�"�*�O�p >�y8� �G���   v�z��7i.�x{nnq���n��5�l�]Q�`����v�����
 Ƒ��0/w��e;��û׺P�`�1uCN�Ios]�6ܟ�[�4�~�q�b�R��E���ؾ�%C�]6Tw+�'P�d��gy��_���jv,�aTrQyj�˞��2^�z)�s;��w����C��&d]�v�<������L��O��T� ��Z@t�v-�c���z|����փ�d�Mu�a}��ť5VL�xx���0n��}� ��
 �'V*n���I���������@\i�!e^�|ss�x{|����tշ��4.CïL8Z�Hvn����}�4�ܓ�����[Ԫ�	|��е�IO�t	5�wP,�5�����6V�0�C�M���FO�+,g�٬���6�f���
��OBN����B�ʼ`[:y���tځCVR�ݼ�La�EF�V2�tQ��yú���;�h�{���M�hc~�ܯ���H �0����!�#��I�şHle�k�mC��s'��Y��c0j��^}�#E.��H�}���z�w�D���O����v��CvwS�XىⲞSBlإm�,�i�UX��O����O�}�ڦޤe�ֵ�WU����X\$b��AIs���MF�t��f���'nӲ��v	����S'Y�GN�]�=�k{�T�V\x�̳�;��u�9=�'��:t�8鎝
��G��nw�w��Ô�"O2t��(]�����fM'�%�"�T�h���co�~�졙���<V�[4	0����?W��<E[�E~�>�;p�������!9k�^G=�vG�_�7 � P�qV�P��9zn���'f�Ԟ蝡C\�*(⢏��7�!�^|�m��	m�j�Ʈ�>�����ns�p��REكMs�
�L�njyu�d�n�c�e|��{��0�~�fi���������u�������+_����k��.p8�Q-�~����=�q��n� �������|�UUp�do�֜�ë����"�-z���XH
|LR~a|�y?c��9P)�z�4G�}�w��s�l��+�/�������F����U�c�̮�qI���Ӎ�hkЙE�n�5��g�57�r$�C�=��p.!co�@��@%�2�J�]6�������ʅ�K�K��Y�*;���-4xz���g�n8�t=v@-#��������������V؏ܥ߯�pCB��d[���Xf�2�{4���QÁ](����~O�W�3����[�0�P��[� h��ҽ�X�/����2(�;d/�aӎU-^P�mv����jp���L�Y���R���a���7'�B/Z�Ԧd͓f����`����B�}ʖ�,�]�I��}��W[�LX2U�V:ne3�)�w����h� >���H����Ң�׫��J�s���}�_)��d����ƞx������[�m�5P(��s��c+��&��$T[K����)i���t�7sץ�_7#��3rW9��=->$EDd�?IY��<�j�o62���;;����ogX5C�vv�O!�����%M�qa ���7)�q�޿y{�I��|����i
z�9d���5���S]���.pxzXL�����]����8��B���L50ݍƉ�u�o4����Ý�1����!8/��V�%�f(S����|V��닌pꜥF]�pƻ)���zN���#��A�tSmޜ����3�����z��0���}���;��q6�f�ai��sxz-3�F��'��,� �fUA���}5�}�N�������]�K����.��	.�a-��Kp��+�G�c�̀�E���;:	ƥ Kw=���U�`���m�����T��/Z�7ٸ�yG�!�/ώ.� L��"|rx�1���'�������c���ڭ�ͩ��������c�^���S�8.)�G)�r���cnHW�����l(殞�3rU��[�y,�N��5��;�q�r���V��d�|k&�l�j���t�d5*�w��46ƻ�H.��3ԅx+��32�ʏtr�*��%��J�zk�iy�.���ѽB�e� �ԱoCo^�(`�r�+ׁm�:���� =;c�Њc�:t �rrk���%��[��U��Q�[S�s�wjy�ʑw��1�oi�xy�����S���I��('�Ms��ʸ��p�4�|-p� >=茆���� <��0�y4�n��z�g����PI��oM��^�ő����@��L2 �9��C�\Hgn���x%�M^.;�dp�Ǧq)�'����.}�����ݬ�	��Z��X�6X9/�8�K�Ue����CE��U
O���A���~&{�Wcx��}��u܍�b��k�k�0͆��+�ŧ�-#Aj�H�����C��i�ߘ����������Gr�WGzKm`o{���zYRbw"�r$8�f��3��k|gX��"'��:���g�!�p��Fk6����e�գ�����=�Wְ��a/pǤW".@��f>��sb`swd�7JD�黍�g7m��#�$���*��(N�B����^���%�!0[�����"��/����$�ŜUn�'8z�h0�&D8gv��X�޲��wB�pe�a����}h����f|
ϸE���3[���d�a�}�g.P�CZ~��L�SV:�/`��avV��;��u�5��u�����,�z�nF���g^j����.��m����g4��6t�)���Z���KB�!�;������6O�ꂜ01M#\8f���h���4�
���TkX�L�����m�W22�l�N�7 �K�:T�#˶t����nR�ӎ7{�&�'� |=1��+���Ҋ�h�����@���n���zaQp��m.��t�xKwr�gР�(�z`Tb�7�O}�]���Q�v`$�a׍���/.��^���y_k���Z$�㫹��[�n��꺢bj�'}#��zx��;j
VS�$O�'��c]�[�#n�\���	�y��12�U���Ŧ7
I�>i2������E��0�8�>_|�kǄ�>��z}��ȹYt���Y��'�����/'|e���Ȧ�2�s�1Eם�n8О�����K�7|�qo&5郲�ن�R���8܀~�09��ȱ�}�r���@�k���#۱��3�wÎ�P:ȁ�G��-?AA7sܮaHd��v\�~�L���y�{�]�Oh����_=��4p�dp�7��;� ����s���|�@9�UG��K�0��d�U�:�Xo����1��Ț�Ñ[�xsM>(p�\��u̅Ӱ��C_1�Ln�S�\^
p��kۤ���	���S��~�?�;c�R�b��E�:����i0B��J�F�P9��?]=<�g�i���R8����A$��߫a�˖`��B�I��pΙL�*d�6���f�[w	�Dܴt�V�{�o)���V[Ѥ2`�Or��->���|�r����W>�v��������u�/7����7Y)�Q���ӤS-��;�=[�{U.:xy�(�,���5D���P'i*�#��Kс����y�о"�7��ڑϕ��~�U��3,��<����c���l�a@��zJ��% Z"�7���t�.�8(8�uL�qf{u�㚸x��~1X酈���c!"�S��5��W���؈��ׯ�'�{���b�6��9�	�
��ot���Q�j˻oG��^�	=.�)�0y4�ј���9���t���{	���l�n�>0����}����`��,��H�{�=4�	��a�a���(�۱�ڮ���p�>>5���7��e̽Q�g���?g�%�$�ln�'�T�$ڝ|QG5T�Zd��׸#Z�����8'�@�{(W<��1P�V����@|�z-�s�kw	l�N�ȷ4�M���X���A(�~�Ù���x]μ��+�qZTY�F���|?N��͛<=6��F[�<����� �X���fy��}�%�a��8��n+���QI�g��N�,ۊ3qn��Pq�����ɇ �@�~`�ۃ��GO�J��b���O'�b�������gS9�X��^O6�lN��)!@����9[�ݕ�G���.L"c�����l)Ӵi�� �r��!Z��#f�'t\���^�y�. EX�{�97�2](���-�k��G)o7 ӣ9�y����kv�̞�O�=�@t�N�ȉ�7���^�vJ�xy �_[��ݚ�	C�	��6ȳ"U���8���Q|���z=�ە��w;��zk�	�7�0�������!|zc�zQ|��a�;��Y�[]h�b�w�i�k�h�SO��	�_�� ��v@,�]�7�=�u��1�p��jo�M� �����;�.�&�'7J,nB�ÀҤ/~��t���$x�CÓ�vx;:�xkx9O�lU�Nh==j�#vi#�ɚ٘��]��tS*d���w���z1�I�s�pi���7H�����v�[w<�Ƶ��!�� V��>��^��>ۆk���p6�ǥ�� �C|��D[S �.�a��$�y��x��2����?H}<��\�W�|a���@srY�}�I����.;�"b8�f�Cڮ�Q���rn�ަW��a��c�n�^�Qx�vH�4\Q��1�g��kTgV�bu�xy'0��#�%�H��碥��c�XZY�<���l�|����svjb���v�f�%&��Y1��� ���]6Ú�,���|��S=���n�����Ρ>���՛�+̓�Ш>�Nnm�74�`��	c��:��(�¤��Y�˖GCǝg5�÷-x����r�;��o/��F��PsiݮA����S�7��и$�����u��4N��j�����w�ޏj/�Lt�A�Lt�@2 �H��s��O;ўq�X�����&�ev�f�dY9��H�	�iF.K���9}��4G�4��j����z��w�g�sM�<�ݳ�(:3��-��ո�v�m�g{&o�r��yqVo���� sy�[ }���<�s�r�n���վ�:��{�V�=�ذ��ߴ�_s��������O�/�h�k�f��?Bn�:����t�neڣe����G� �&�XΪ<�E�ο�@���^���t�2L8�k����}|���M+�Kf����rlogx2�]CU&�(�����l[ç��B9�M�Pc�����y�����ZNf���(���U~��=�n�Zs�H��#�n���D�-χ���\��tc_����^�}�����^*�G�����(����K��<`v3���oӍ*�<��w���&�z��ڙgL���[dl� Z������'���s�Tc,u�2��h��S׵�ߺ�r¼�����������;�|Oh1:�K>�c�F}T�@֎N'Pꁥz0����Xw�_ݴ"}t
��h\i�|0��ʄG��3 �r}���\p� �>�#��0���%��jd=�r���e������֡����w�6v�j�f���FI/0�
�rK	L�+X÷H��C���'W��������֠w/�4���3�����#sO�7�wo(�5}����nr�F��-�r���ڥ�n���?9\<Ӥ1Ӥ �  ]�ί�=o�]��\?����[k������qN���+!�7��6�|���4T��k��w�Q:gj�bx/�C7���BP����el�$�kM��^���=��5��W����7kQz�{��@��pc�}0�'��{,b���}n�����̎p[`B�ح�S�Gc��J�G�#�B��Z�{2j��^�q�|E��u����۬-t�F��vUjZz��FNN	a}��T�VE�f�.Yc� �|kc�=_G��w)�>�sd�&:��o�Z�4OC{q��|���(a���<�{niq�!�42��`�}���+�)f��ixo4�1��l)��j4����e?����Q���1�;�3��E�ߕ
�Z?��"?�5b^K����P������ѳ�'r-��1��􇶎~�!�Q�~���%y]��W[ە{ߗ�O��7ھ� #*�no2q���dW=yrT(9�/N�]�0�ȯ4�
%�6�a�.��Y9u���tޙq�E��[fa�r���o��nosX��ݼ�A�3E�H@g��Fo�us�%�赣Vz��҇Z��G���"OU��Ɋ=ۍ�V��9K�]_Ht����c5)Ȱnܸ��b��bX}�3{� Qe[[��R��b��^<�9`fy�g+Og:�R�V蹚I���V����r��[f�V&�`����A�7Cz�pd�U��� ���]I����+ks��bnar)؍wum.Q�Bpv�uM�o��;]tk,�Ѵ�T�EҾ4j�éz1��e�HẆqq�oq�8Z�q���r.�hJJ,����𸦞��#w�YW��l®5]bs��woZ�Oy����m�	P	fN��JxBXӬ��]��}d<�ƪc̨�p�=�.7��bW�d͸w&�or+��� �!
޴,��{5�x��6�1Ĩ��w6em��Zٜ��Z�����P�`⍃�Me��/j��i�M`0�:�܃���d�Z6�����R�pv��aUmR���M��U�j�q��}��֟B���[������,�o�׏}�O��Ӎ\��.|;p���Kbⴠ� 7��-����*���۝�����_Av�Z	V��H~D�m"(�!��/X��G�odtv�A{������۳�#pQ�����D;�T7��#�vv
P\������>阊c)+��ho��`l�h�U勢��2��1C*��`�t&�N1���+R��S�H�� X�J�	���B���We�w������ѥJx��{*�ɝ�T�;$��W!؊��V>��ӽ%��K(�j�{[,��v��Jm�K�۶\�̦����s
[[�ET沞���sj�.����`�����:�[(�5���5�2*�ɛb�o�dm���O1����t�X��utwhޓw�YY�sq�o�(�����Y:e����^]eD'Z�š@��r�͹�3��9F
����܎�X;j���ocHqHc[�p�]��3���Ղ����J1���}b�[�gHUPZ0�Y�6U��@��޸���@���c�3+={���\�]t�x��~��5)�>K.��Y*(s+�)�a�}�X�^h�g�d�vk�!r�39d��j�G���WHP����t�tn n�[4�i�e�M����~�
³#(nQ�)���a��S|GM|xM}��F�a�ݰ��58��;�s*��5.n�.��ab&h�,�e�4�����hHb��;N�r�ܶ\Ε;�����5�T%�g�����"`��HXl��[{z�r����̍�v��ҋ�Y�zPRn�:C�pҁȚy���,N���u�3���9�9�n�3��ݻ��>I������ڊ��&��ΈU�?=�H���>ִ�dUPPZC����
���9��`U')eDD��0�
�:����a�#�:ݽ�����7���ZֺkZֵ�cZ�Ǉn�������g�%�����*�ԟ����U:��̟�rt��1mP��\�����������Zֵ�Zֵ�cZ�o�ݻ|v��	��$�@��$�t9�C*�����~�G�
�d�HsȪ�Ȋ"�+dr��*��C�����r*~P
*�2�
�ds��;��j\.Z!+TB��D�y�QUTT�"Nu5�J%�Ȋ���q�bp����V�	4՚��9vr��" �D��Ȉ� �v�r��ETr�D�h#�#��TW8U\��U�I�m�z�j�J"��g*���B��(((/ZuY3�r�Q�!s�UwD��r��J�F&%G"�K�\�*��֪_�
tB��EL���D�Vek�¿!�z{�QQ�QUʨ�>�DAAQV|�I�*�E�r"���Bt\�J�jc�ʉ���#Ϸ-N1_f��}kQ�9��rJo�3�����8.WB^<�Y6�93)	���C�1W}�	�jj��uX������>�"�:c�H��>yg����׫���@�I �O��,����x����W0�%���=��D�:�ou;��b�(�+#���F8O�㡃�l��^���~�R��S��%ԘWdx��?<�\?R��=w��j�J�_�[Z$A�����.1��U���Ԋ��)�����3����';��? �=��Ag�#Q��s�� y��{X����.��}f􎷮vSU��cl�`����B��ֽ�歰��Lc!2j�2C0�@}�"Ţt�gFk{�;�/��d�	��j�^�P̵�%�ȿ�3�ևr�R�mos�?���,�\�f�C�#�'�0��گ.�A�Q���v詙��.��e:"�:�w����/�E�ӽ�ᫌ�ń�|�"�s�Ox�Q�2q�\����u{�~�<�}�æ����=��;�=�T�ێg�~���?�w��R`yB�0,!����P�R��KǙ�G��gt�lt��mN�ۈ��:�k��Ԕ�p��8��¦����g������CA��g���W�Z���\�㢔�������P�N���"�3-l�*nԻ��׻.����ml�����k{c|NB)i��nZ-�@E>�eӻ�q<�eS;*4�	���}���#;��s�g����=g��9��|�8�W�&������ӎ�$A�VDD�{�oI����{u�� _�ʅs�+�����Ui�6Q��ZHS?�^�]d�0UƗݳ��{ǅ[�[�7m�֠���RQ<�ް;�0���q����l�ȧ�rn��O�G?a��5ykN���Sv�s�Lx�o�Ä��� ���������� s����qkC�>���7�;�7��������1$~#���>�r>��X�S����IGVk]0���ȝ�&О�`)�6��|=L�����4&1���t8�qI���3�+�ֵˬ<�l��/�ڡ7V��K���(���.�_4x��=+�i�i��ʘ,5��M�c�����'Maq����ut�;#[��u�-C�e�z�����+O�0$s�/ڹ]�7�\��{��t�sE^����"[��\���s��O�p!w��m�c���;|�����k��f��W�������o"�)�l�Y��|ԧӯA(-!G��-^�M2옩�ˮ�����v"=p#���uN5�<�"�};|�	�۟y��~�$87�&���*�?K�z��͘p��NŇh+��W�d��*�1��މҍ\�8��U���MH^�&:HG�ߴ��5 �˲�����9V�Md�gQ���bw�y�(�^�9���Xbe����N�e���L���k|^�������ӎ�H�ӎ��p 	 p ���6w�L���\��7)��:�릮�Y�˔�)�Q`9H!Ug�^u����=����x��_�H^H[�K�����ɴ�V��݄�Fes��v�0*��(��7��Ԍ���k���P�
�A����^��dxG�*kf:b)�󵙾'�I���zS��K���ǔ ���F_L> @��_/_�{��7d�^]Yպc�x��{�o�Ы0�wz���sW�r�Y���1��~�"��Ëk�s�Z�SZ���5Q��g����{a�}s�< j���j�8O=w)��Y��yi�����h�549��E��8�f�\"X\� w?c�z��_a	P(oK�=�)����5�]��O4Mu$�%��Kp��zn�[:y��x��?.� �xEX���gX�.��P_?�����O?T�E���=w����-�,��ٷ��v׫_y� G�����Tk��0���֥3Y\��b��Ȑ�/z���cwx��<�K`1i�>g��>��9���t{� ��뵚7J{y���xM�;½;�]0�7 �K���y��g&���^X��8th5�O��i}�4팍A;S�w�����-��ZP�d�W$et뵗^�n���$��
_V��� G��B���������֦�)�`����]x\��,��7R%ܘ4�uؑ���t�޹��;猶s{5m�w4{On<��	�ӎ�c!FAI=&�u��z8vvT�F<6������H��z����<ݬ���l�{9}3WAöN xv�!�oTτ��L	m���ZɎ�v<�}r=
�FU]<��Z���߳��Zm4	l|bj!�dÃr|�d�rz��"Ԋ�1%��}n�Ԍ��=3L>S��꼻�@ck\�h4X`|a>���j�\�U�.�d���͋7� 쬾%�I���Hp/̟��i�S���e�{��<!3��p��NpLxswS�^�T1kw���[��l����*4���P�|��C0��Z������$��^zf�k<��78�����Ŗ]�oU����;#�=�k���]�H<��S���z/6�6%�kY81OD��gn�t�ќ�	�-�����|�)颔rqB��(75�\�n��z�l��T��U�r�n��7t�t�/�RO���-��TEq���j���ϗ�l1Û�W�)��-6fY��"o3�ھ�r�e}�~x��B5�:�x�c��gܮ�]B ��՟�b�l�	��}�|Y���=V7�f���a�V��@�/ONY�v�X������'�T�5f.�,^��%c^F��������+��K�V�v)�ڪ"zNȳ݁Ms5�{{�k�r�YNA�������!7�o=��縬�j�J���N���{Do�t(�N�t**+��7r�O���	p:Z����]~�I�ܘhm;<fR�c��x��OP˗���1�y	Z��8�s�'t��b�>gwM���O?w)�S����Ű�p>�b��zC[W?s�����ENCٵ�g�����H�2$��&���sw_��K��A�Qz�w�xa��a[F�:Z:jZ����'����cxT_��=c�e"��4�T�{�P7'���[��5���&���ϲo~�v�lU)$����K��+��N9��'�ʆt�Uವ�W�J/-K.{���0N��uI|���ǥ��Nõ4���"G����cǺ�~_?>ѹ%_�5�.��b���YT�
�Nv6�ӆv�������>Vt��$b�a�B����cӠQ#����N}�8|��{�ԯ-i�0z���Q{�{n�-m�����v&}Ƃ#�Ά�i�=�?kU�tg��.�V������ә�{	@�JA�>�`&��`��͡8w�Ьy��=�{4����蹇f��n�q��ad����}.Ƚ��DS"������[]s8�켫w��D���+3L�q�Q��W��Ls��4wt�Q`��nay�ݽy$[m�ڷȪpXu8Yq�;*�g�ԭ��hѠ��c_		9r�ss��R�^Z��*����8��oW���8�󎩾ro���K�>n�\t��N�t  � 
}�m�y��Ϗ�Ņ�������z��HWn�<�3 ��1J��SL��i���3�M�ht���ż6��f�
�i����n�ի8-a���S5����_q��!���x�ӻqRg]��"%��k�p��^9���S��=!��!ܯ'�?� j6D�t�t��b*�'L�gm	n�c��^��%(��8���_W>Y|������|�3}ߎq���{Z�iX�q�?��<�a�V9P�ύ����{^b�j�39�!�b��vǱ�,�M0���wZ�a��5�����l��� lε �����y���қÚ��B�+%�^���'�Vp�[�d3g:e(��DAg�/Ã�h�Z�^����,�BN*��3����Kw=��)���9�8��#�F����9G7�v��s������1�-/�k������<Su�.a|�y?=�u�	�y�UV��(l�u�
�5x��wv���G�;��ژ�>�"Q��p՚�OvM1��l.�[zVӷ]��^���{� L�f��t��{XZ7���BgzJ+��̥�.�|��x3�i��­w�����bTP�����WBʧ�șBp� ����0���mm���l.H�W��o{sY�n[��3:N�^�Ip=j�H	�ީ��Z>�`˝o��]+S���vkvr��V�D�z��@���t�2(��8�G�3������V���+���8�L�X(���HAt˺&U,����k�渵�i����p��l����^�#[��A.{"�ũ=�Ƿc��3L0�)���ͨ���ݷy<O�臞��[ @�6��o
'���:OT�L<�L�����`lx0lì�-�y���	iX]��8p���^D;' ��6[ʯ_���t�m��> �Ϙ6�%��A���g0v�v�9�;C;^?�1��3\�=��� �sɓ��pXo�.|y�����6����;�c��+���=r�{��ƣb����9o����O�_���Ó��떲��n�qJ�g s	<��	��IK��L#F?�LE@q2�|g�kH�~�h��W���b�IO������<�E�-�>*�!Z���|���E�eO?X`q�����e��6zp�d��}��y�q�"�p��z6'��@���~��Cu.��8f�ܲ��l�={��L�S�ſ?l0㓋x�*�E���
	ƾ*���<쏶�~�@0��]�g�sWcD��r�aA��6��6:1h�f�靝�z������ �ez�K��K���`��֠�o����oc�M7O��	NOی3$7,U�&����%���#x���RmU��瘧"����3w�JƨD��T�a�lw���`(k���;fu�:2ь"���pv��D�"̉�}H���2B���l`:J70i}��5�5ŗ8�Z��n>8�P��8�EC�f�fi�k�gy��z�/���ƭ{+�Fұ�<��?.�G�V1�n{������gw/gf���J6�=�'�O�7Rë���߲��d�H��
��'��7M܁�8V���������kJ'hp;%�U�S�G2ou�0+�Ԙ/'�Y�����`��9�B9�5��ĵ�t���8t���.Ds��Uꖭ�L��b���Z��^ �zi�f1��=�S}q�(l��E�2�1��L<6�Е�^��u�[�-'�$st�wA/A����Ur�H�\k�'OC;o�\��EK���2'_�`Kl��� ��q�`�]P'�r5�?~�f�r(�4k�f��N�]�pma  �^D;'�Ծ�Z�<^�|n�TC����*����xk��s8��O���G����и
�~:cX~�D~Y9jFyC�N�ڕ�L�p��M0�		�[�L=����� �S+�iF�|�
_[���������̨�g
�W��Ϩ���D��fM!(f<��^��^��&>3�D�~���=y�������-��&/ꌶ��B	�jwҸ��c9IuE1�t�>t��,D�]&���������sӔ��:$}֩�
�z�d�Q����Oy�ͦ��":P����q�pf��n)bל����&�]S�53�Z]_��������naq�۵�S (l)�����׵��odV�@g��o�LU�zk��e�[���q���i=��s�<�¦X�9Sl���:x3.#��f�"���K|�
t]k��P��ƽ����!��-q�*�o(��pP-�T�j<5a{�]�"���F������0�w}��u��ӻxP�=k�«�q	q�_P��>B�yV����o��H-zںG��owf;����Ӗ]|�W\�&�'���y��!7��Ҩ��Gs���B��ٸ-�}�*��ɾ8O8��-O�[��u����TW�'��ߣgH�o环��zD���4��fm�k��[}d�����j �7z�x����9���dW=.J�y�Qzw�xl�S�Ӟ�������n#<;H��v~`��T�[�n�l�4�T�t�[��
zc�dsP�֯Vy�O	�c�A�\�̒�f.ᛎ�;���z` pqls΁�}��S}"U��U����,��}q��;Qb��]�������">�M ��5�$:�^=H|{��^S�J�d���_���].+�4��_��p�������UI�z 򼷘x�Y�n�݀�]c��^k��8�U�n��\��Q��-�9ڶ�c.�b以
u����Bgfc��l�:EY��1s�OBmOL�5��z�\k�i����{~oo�:E��8�$$	$!玻�|��u�{߫�M��:���Qm�$ ����\0j�����
9�8��y�=��ϫsOf���N<"�N����I�K��֯�[5�	@xu�0��g�q��[ܮ�:���|�����S�'Ǡ��)�ֻy(�H�:�OB��������L�<�!������䴇��,E0g�{#r����W ?���&������%��<�Hl��N���^�U�e�[��Z)}�$ǇXc��
|���t����X]�3�ez��K�����ћ��}9Ts��a�\���,��ێ�!�&xE�"���ZŽ����KgI���5ۼ�p� ����P�{$p��y��m���\<�B���?����2_����z���R�On�ך��!���`ۅ���%�IQz�]�O�͏��[�/^hMJ&G��A�Nx]�z�ێA�%	��������\� �YB��ǡu�kTX��-=��i�}�������6D6��9�����Ӭڄ�S%>�Ms����0�s��u�3�� 4�ȶ[j���̛� ji�ŗ-Y����R���бT�ވGgS�����������ti��'�N�K�X�d'z8��$y;8Fq<{����ִ"K
��U����.,].��QZ�?H���𵌫�U��5e2m�:����*���⡩,E���ʍJ�&������t��.���]����s׎Rw;V��:]gqRr<i˔�,�����6b31��nuP��斚S�f�ڞc��vWC�!��,�2��.
U��ü�˘5���	����iv�E���m� ����p6F�E6�����t�o`��w3���@��1�W��L�|M-��$���դ/}���k�H�ʴã\5��(��;gr�w�!GS�]
�jr�����"�'���(qD�~�+9*}D.嫤μ�3�0KҴ�sp���qTΖ$;Z�5t�fBh�)0�ͽ�kI�ŵ���҅�Y-|�Y�7dn����>�Eb��v%67}�w)���#YS��Օ�2�a�t�k�x�L�y�C�IRna��f�oy��HnT*Us��;���������.�<D�b�Ym�yo��	�`BP�6�J)�rd���!n��SYFn�]$E^>�`ڶ��c���c�����a���E�X��w��Њ$�6�6�0L���1�*gfಇp�^Wk_]��֌@6h��f�����a�`���J�!zc��K*P��H;J�vK�܁�6 ��o,Jtq>�L�*S9�D:�a��n��d@����]U{x5>���a4*w�U�(�H�7�ʞJw.|F��ˌ�iTba�j��3/B�Z	�L�2 :nowm���NT��miu�fu� ��{��k:l<�nMY����Y|7��и>˄,��{O��p��c�3����lo7Ѫ�#ۄͮ�����v�ƸA��<*�L�]�m*�|9�r`�W��t�p^nVVO8�OugN�j�mK��P�Zu(3�ʒ�;2n;����k̵�)Ji��Νp<N���OBlC b�p�n�9B���оu�T�����}��E��y���}M�vH	BL��:� �����b&Б���x��9��y�`iZٝ�~�ck�!3Wh�c���jy�"QU&ȫ��3���+oI�`o�{�MN�9v�t�+t�A��Jު���;��x7��hcW�����maY)\z�WNw69�2wl��
��T�����KGj���B̒�0a�3�&7���D�yC#����6_.�*�-��6Ջȸպ�Ȼ�'k$n͠V�u,�b��[c3������ἜN�p�_
��:j�N�ƓGs���cn��Fj�����|��.#�HT��|�~7Op"�T�*��yU^AF$E��s�"�"C+6i�B\�EQV3���ӧ;xk���]5�k]��k^ָֻ}�;v����=B\�E���}�e�%�(hAM'$�o�,̈�i*��Na���:ݾo��}=�>:kZֻkZּ5�q�v��{{~�o���G~�z��(��%3�E�c�:W"ڤ%&X�,�p��T�q��DQ"����C�K��""t��8x�!#["�
f��8TT��"�T��E^4ܽ(�q29Y�D~b����T���D#�ߗ��
��vikI!��r"����Q+%Jԙs6~�UO��E\$��\��9�_�Nʯ2��R.��:BMY]D��.��(�
*��5��AIs�C��*�HBlΊ�DW.jQA˹�,:�D�eDG�'��
T+�B
.sSD�ʮ!\�u�QfΔs��돯���=��#�$%9$�q�.#'�bA��iJA���qĈpx�M:S�j�9ꣻ%A�n���P1X�q�՛�r-��b�M�!\��/E�]t3��pV��M��x�p-'{J
�ш"4C�F�FI���*O"%RpĊL�ʉ��\��59'������z*��x��ޠ�	�c1
(�Ө�1�$�)�[P��&e7�"�!��Ba��ɹ�[9�>Myq�t��J$�B
�"H����7�y�/2oy�z���*>iGu��#�^t:���]]��Y�ٍm�4��_��k�@E����P�.y`! U�b;��(���?�Sv��x��>7i��Z���E'��ʔ�w� <�#(D�~rg��%�0�LR~a�/�~����w���Ӿ���'��Ĩ�6�����ޚ8tz��S�l���+�M�7a�,���y��C�K�K�Q|寺*ޞw-^�榐�������#Z�&�W]&*c����5��3����DOe�zf)�5{3���.�/]���C���K߻`&��N����5����n�f���H��s��sBb[:���������s��O��L��za^�u�
���uE�un���.P~/0�Z}�v�z��m� ��/϶�N�y(-��2Vļ�_�o�2s:2m-���@�{�E�X<�H��'�}�	��<�l�zZ�Ff�����5��'6Ȭ�Z���.M�|$�~����}�|l�üpr�=��:�T�Ns�R��']�C-.O]2yMՁ���I$��l�?un��b?��k���[X�O��&O�����f[���3ն�;���.Y��:w�3V#X�%vpy�U���޺p*�pd���W�&�{H�T��ٔ	EH rD��U���UZl�^�m�]zM㸍���I�]@q=j�2=к�y��st)��y�T;�i�2��}\�{�"Ŏ>8�:t�	�	d/=��]�Ϟz�A�7�1�q�#vz�!Z�ע���+�13T)�����>މ�����n�/�=��?`��s�=6�q�Ȅ�Eo�s Gwm�i�/C��'jw"�c�]Z�]ٸ\���2\!����l9T{w��k>Jx4��<���8�)���>D�)ߥ�����7���`�.�x�K������9E���/�Ü��ú)��j\�z��W��m�B�<%u
�+�)ZO�y��~B�G����F�E�F���q^_U��D����x.��,�R����皤���~�����DwH�rt������/sI�ӃK?��� �����WԹ�Ts�L�R+�u&�(���y�b�p���k��͎��un��է(t���q�iw�ja�rt�%�{��0��X	�I1^h=�՛WJ[�ݽVn�*�w�gd5�ü:י1-�7:�Q��񊰶G7K��㱜Dp���U���ȿώ�]��ga���}�%�z�* F���-���Z����f��?v�����pz��^��"^h+V.cuqu7&��\ư�#]��R�H:-�X�4{��J��rW��e�آH5����\|f?EӚ�
��}QS�هcwx�oPi����6`�խ��>�Ui����}1T�ӻ�hdT��듮uu�u�z��g���N:F:t㥁$DB0AHM�z��ŝ�ӥ᛽��d�W�5�4�C ���}/0����K�e���1%�� �I�f\m(����4��b���>�
gZK��+�=��:+C��a�ʀ|�D�F*$t^"t���O���8I�K�B��TZBsn���ø���4Agh@��]����s|d��v�藽�{��	�\�d� �����3#9�2F�SU�Y[9�"]W�z*/�x�ُ��߯��ej@�G����zS_y#s��G��ȃ��I�t'��J}k�����A����jl���/�c��q���[��']���n���P�/�A��<m����j�v.�;7ck0k��J>�y�+�N�1���a��DPv�5sm����y7���<e�v���'y~ށ-Ԓ�gNm�0��u[��;�n�j�f��ܼ��#��vPC��9���:����A��%��B��=I�ܙ)� .5+)��rx�|�}��eL\�:�����sn���^E0C���������P�����C�GJ�q��'ۑm^3�����"5"���TD���Z��GՆŞ���x�y�a֫d���P�=}S��ۨ�QzB]Զ��or�(
�K��9��H'ʡ�Wu�/zt�����$��&���I��<��{c�t�Ot��c��ڕ5��w�����qy�M��=���t,t��L"H@�<�ד�]��^�܇���Oiö��A�0�U���7u�2+���S0fV,:�O9��6.Pٞ�'�I�ǆ�l��g�sN����0�7*J{K�6Μ��͵�_u��>dT��G"{KY�\p�*gԡ�0��s�'�y��T_�����w�v�ygH8�zqU����$�.�>'�w�>M ��b�!��ǰ6>=�Q�?T�Im��Z:-��<m]��l���q��S�2[��]k		�K�c����`����7�¸r�׺�Z�`%�������|��/}Г�_T�ε�s&"<�tG���*Gl��ot֔
�=�����K�N�IoH��*1��I�b�UY��C�	��:[wɞE.i3���;���f�!�(G0���u�S�3V��Radħ���kג��S�L5߳�7{}�Nmr�y���֮/8p��-/��o�>_p5_,"��g=y,���-��ݑe�6NuP����V�����[��@��ׯ�ʆ@ft	�~G�Z�僑U�4-Y� �߽Y�h��v��m[��!+������9vj��I���r�w4�!s���X<�9S%^:R�Bgp��`X�ʣ���\�g0�R���X���@�jb<
�]�>ꒇq�1789LB�'�pvV���q�;ٸ�彌���p�@:�Z݀wn�����.��3�o�Q�w)yGm�\�z�����eBwGQ/"(A����Q@?1znCxf�M�2���
J���O̓cڜ�1a�=�DS�}쮮�rd[�f�]IeӚ{�+�E4�"�ob5��tJ��{�8�E�SmlK?�r�Nl�fS����,�|���S���hd��s�*|�1)ƀ��3'�O,�H�c�M<5�	{�H�^n�os�syߛ�-��Z}��2:�O�h�u�P������Ú�wu� ik������.�gk����c;E=���z���\������Co���o�!�2�`GT��s�JH��Ό:v�iVǖ�&�(����OC\<溘�����%C��ͪmb2��-Cɽ�ޒr������b1�W�c��{m	�M>>4��r|{t�Ǿܻ�e�SyY�N�	�t8��L����_��2���r����>h!������77Nd�{�˺�~��Z[@�C�?��Z�	�Zc�.�C�}Ob�5�hwP%�i��$��#����m�LɁ�\ "��i�*��'�`x0��:�C��	�����Z��vK?���Ok�����8S0.q���o�����	��K�z�=�S�
�9S����l^o�P����f�^ͩ�c�){S_Y"��a2�������yk=eU���ܖ[E��;3;�k�p��v��5 ���}�ݧj�o&S4L	~ ��<�{��ݻ[��@S&M�a0�
 ��ua*�.�,7��8�`G\�q�����W�c<��Y��ǉ��vL;Ks��s��G��`8�f,~�y0��|��G咸זV0[#.y>�=�u�<S��V��� ���n(@�A�-LX�wkǇt����8��iᱻ��l(��ւݼ9�cNos>�`�cv \��^]��<�[���z�<e�.�7�G%�l>�;���L�����߉|��)��z�-��T����»�/������`�
Y߯�"����C�iY���IY7� 5��L'�^��u5�B�M��;�Pz͜��]R%��fj��a�и)�[@��]���Q�a>=9�#<���y�����z�ӹJ�v��*���g]Ex��A���1!�{�:b���]�M6ЄY	�o��/��{c�)M7_���P�8���>�h���PP���-�!U��!�1�>ӫ�;��#�;lSI����Ď����:�b��u���%���涸7"NE�� c����m���᝵�p���`��Ⳉ��m,.�
7���S#��Z_�/�^˞h���N��W��l�ީǍ0`X��)g+����/u��t���2�����r_����V �N�	�6��Y���v��S/wdo{�:dY(�ź�{�F��5��JH�4��A�"D"Bq����<����������/�$���g>:�e���E˥0,��v\z1邝�մS�昽դ��sЄʦ�����m7���In�Ӈ�mJ`j�J�+ys5u�(�_���ìtsL9���-x/�}"H9<^V?�su?s�>���l���ԯ1���1V��=�0���SK��"�0B��/�}����tׯg �`��q=[Qn�C�jj��w�h�o�<3���]�͑��I��A^�|uXi��z��qH��vRL�ύK7g��0z�Λq�#>�S:��>j�;7�p�C�q"9�O�<{��n�a83��\������v��䎓�S��İԄ�����ۦ�'��#^�9gn8IQ��##���a�$_s0hK�ꑭ�[!��Y���f-�قQz��������Qn��U���pR�!�4z�ƴ�Ƨ��C5�X�˺5M;����O)v�G^tŷ3O����ّ[���~��)i���%`�$� @�dE���+���__&��c �F���~��{r�S�5��͵�e�+n��J��d\�Jf�,��vl�$MWq�Zý�F��[��THm�t�H%ϋ��x�I g\������,���u`a��Y�L�K9Y�ozD��,��=�P/x]�-�Y��!��to=�{OR8��PX�M:qҒ	{�fo �{n���ݻxg�o��Hi���b����X��'�$]�E������f�s��&(����[�I3�����Ї=�n��X�AA�.b��lg9����Ej�)e/�#|2^]}�����̵�w��i���od�eWʅtq�&��kا:�P�W�¾>�n~{q3��v��_��c���nKkW�a2On�y��H�����~gO-�h�P�Z鋼ű35�x��P��ɸ[�q>��ʟX��� ����@��3m|�,��M'g��o,�van�uo'�2�F6��9�Ъ�X/l���CnLt�[����l�t�w_n(�1��!�˩�\-��.�SY�~⯂./�����R$�[|��6��0x˫YyGw:�����v���}��L�T���>m�||}���f sjz^S�6�v�Fa�ZI=���� w8� ��»���a� �?"�V�AC�$V�-"�ݎ#����cr���C�4��M�-{�_Z�X�3��{lι,10W0�ۺ�`0�n|�:nvV}i�?�%QC䤵����}��'�yc��4&o�8�`�r���"���d��cܬ�Ki.��]�� �8���T��>�yt�Ky�\΢���݅��Z̺�|�"���ܼ��$�C{h����<���N�t0���9�}�9�=o���"�r�Y;���gB�ʖ���� ��������T��|TGOl6�)��N�k�,�D���
�G��ui�ֽ�v��w�ADد��"_�gݳ|�tI ���C3�f"/�M�:�w>�A�D��o����<�%)fk�{gwٹ�����҄iM>�WT�>{��г�5>VEN��*�@��s���F4�o��[��lD�<��84���J�ӯ}�Y���^��>?s��oM���KK��5;��^�f����""=��]'��{�yu��G�y���m��=C�C>]�	,87s�K��uG1�Y˓���#�_���;l(X��S]�ʽj�*�GԵ�ߵ�="�JY�W�P����]����I[`���q�c�r���ۤO5����T+��P�c1�K��u�ٗ�8�r��^[ӯ�靠 ��}�%�bS�+̃N�M�y�	MA(�~�Û+fzr�4�>���S:�og��.�t�=���4��!��{���	�{��('�:�(̮����4]��k5'I1�IX�K�.��|�����sָ��w����s��k��#�t��3B՛׼���7Ѷ��NJ�ު'��dT����k'&<��CSl��)3��43�Ӛ�ge-ݚ�|@ȃ��x(���b���g�u����������Px,�O����k�a�f�vDs�J�~}�rX��,`�lbj]�_�W�~���biӎ�$H2�9�7�ף�w�䢹�	T�yGhi�n�g*�z׍��iQc���@h��s��6C����Tt�� Z�=Cr�I�&]'�r�wBeCz�][�C`&�h�;�՛~�Ó3��wTM��A�i��f5�Bc�knr�[五�vF�MwP%�ݐJzw��}�"/h�N������N0���o��V��<�_O6�ƽ�D�~�]sy�����k�v�l��k��������>׆p��-�
��_�a<�Ph��>�f�y�ڬ�X4�>��.T[^��j��o	���~����?/C��,аg:�=���I���&O��n�QW/��'�������^<��ݷK���I59����hڊ��;�|��i���������OM�g\��|D� ���W�k��m���o�nU�v�u�||�
J�|z)s�F���O��1��/�;7~W�aY�ƌ�n��\�%�޺�}wJDV��:��P]��ŧ�^m�s}YL���Ԫ���=��=�5�����?��
zh;��fn��l9��eq�a��ڠ������N�7�v����76�p��5ej޻���3'�FphՊ�3���c�5wn�b��I^i�I��ϙ֤��2�.�z^v�����L��DW*�T&:/	!F(CMŚ��	,f�5�a�ne��"�wrUe�^�idn]��\5f�WJ�<�ǮvvWuݶ�:v��8�Y[Z�Pik�\ +Z�����N�2���6�v�5�$u�ʏvX:Q�CF����S�� �M9zF�X��u���Jn���6��ۣ)a:�,������J:%*���N�7�%����,д:��.�dXsN=��ܸ��!θq��R�A�d�8o*�U��z/6Ez1]�ST� ��M.�ʗ\1�,�bh�ά�',��:{�B9gk�����$�Żn��|b��y��H�ҩ稁����1���wi�2=u��)CTD�\_n7KE ��*	 �.Jً2�n�얺�M
sܙ�\u�+N[ȴ.�1�i�|��Y���e{����j�oPf��z�n`��*1T���!���wA䂦�tgL�b�0�;
D��.��p�1B��(�u�O�ur+��8< "6�r�����uastt=�Xi�����:�S{��A��A}M�gXY�p�T5�έ�UP�!�����%D2���aov��N��o����� v|�t�dF��Jp>Wc-����K[|��R�~J��y�͞JO,�p��{묾�`�k�\N��`(�?yv����Od�l��(u�����sF7I_�Rĭ�R�EJ��<}��l9�u��#����khl�~���sZ]s�H7�*q'JW^>�7j��bj��^�E�u�:�d�2뮐��b�xt�Ƿ;�X�
���*=@�t��o0V����]t�I���K�e^M�c�h�LԄQ�}�[m�1���.M�L��՜Ɖ)�t.d以�������n^� $�[Z2.��t�	�.^�k$T�VWurؤ7�t!����]����y��p5��Z�-(B̾����tu����;�I�7�DZ�b¶���)����n�%&���:�;����2�5ʋ|��9i!TyӺb��i�Ǹ7��{�*A'M�_j��yT��'h<{T���.��>rw�˔2�i�m2NVwgC���I-,�ߩg�Y�$���W��Y��)c`��m��ޫx�W�����T2A�]�Wp9��j�U ��mC���L�|{,��H�Z�d4�i>�33���<���յ/�J��v�;�^����\�7�6�.q�Fs7�T�퐪CC��Z&a͹@�\#�ڧy.ɇ���]�n�Lnr�Z�-{Y��Y	=z&�����*=�g�u:��ӷ�&�r�{`�J��s��
$ I�T\�Z��'�@�1�D�3��)ƈU���n�{��<��>:kZֵ�k]��k��w��{��������U>�!�C�]l��VIEUA���$I$�&�t�ӷ������ֵ�xkZ�mkZ�ݻ|v���D ��˜�eE�4Į[LK`'�"e(��1��8r
*��Ј��?wukD�B�����B$�(���k��sV�LU�%Z��UW
*�%Ti�E%a�]�QRt/�TG+�w|�U��L�ʷw#�P�fTb�!ʧ-$�*-YX�	$(��>�

$�]���Vd��w)�-"�'
���,�Dr��a¢�,Z�i�r�9��Xe��A�N�LQQ����o���W��i�o�6��]V�J�*y��y+y�̭���Z #j�5V3ue'�q�of� w|qSR�߽ޯ/W����37�{������2r�l���^����>3��.�,8��a�;��+��%q��#����͸^wO'�&4����/EE�y�*䙋��]�-�1pq���:l�Fu�,��A��a�!3=���D���`��K.{��u��7�t�~����|�ZĠ�(|~B����ǝ��ۼ�ä�;L�zs	���u���%�r��ϵ�9���@�N,V��7��u��\���� T&r8�Muw>:�e���к���N��ya$>n���Q��*�����!:��k�>Qcs�r}�����]�e#Fri�T��zv�d�In,;� >KE�ȏ�_Lk��H��~������*�'�Y^��su��hh�Ɇ=9w>����+v֘�U��˙ų��=���q�d_a���l=_�tׯg��^Q#uU��~�:K����z���U#+�}9$k�+���wV4|��3�(v�Ic��e�9�v'���Y��-�JS:���H�� ���¿3*n�p�3)�	���)ɿ�>��I��]G��.��Zv�(4�"'bv�#/,�u��m(�TZ�ԨI��F:�uG�2��2��A6��1>^�#�J�X��!ͻ��bY�N�nN���Q��xX��9m�Ao>�j��\�۝z�1��d���Dt��I����a��r�x�[�%�9��p�1����S��s4�=i	еE�9�L��B��y>x�=�%Q�bV�1��N�����L4��ˌt��2��_�n���"t���%��Ѝ��!F�dŬ�8]�}�/�A������S_|��7���⻣B+۲��]�:S�Պj��=���������m�Tm�"�p�`��n�ɸ�Ȩ��F	�nG���/ۄ�� ��d�mJh��n�����xķ0Ņ���T���������U�9^���	�׿c�l!�W�%��K+���B\t׺�7������������ؿ(�s��˱��W�[���6�c��ܓ	������L)����Q�K��[:��}��3��r���!H=��n0Fܦ֠��8�'���P���~�YgXb��X8���q��XuX��w.�P������_z0���>�w6D�eW7�����dW;m��-�W)z��go,y:�����^�ǖ��0(Ƒ��z` ^}n|��qL1����Q]�E�uȩ]k-^'���ژ�
�.�,��!E��r��p[�ܙ���&]�EL��B�w8BL��e�F�:G�ٛ��+x;*V�Ke��|6N��ԋ���I}�J�W��[���ͽ�<%>l��Jh�Z�$���̖u�O~��u	:q��D$��z���xwǐ�|Vn~-8��;j�C���b��F�p4N^!{��ܪ�;k?��}�k�+U$S	Qc���>G�?�~cj�ݽ[v�.�:���%c	䧓�K.{��� &U���'��nC��snz siv�#�a�&��siiQ/�%H�ܕ�-.��v-����Z�5��x�;�w�8n�s+��tI}W��f��;X0�M�00�"���RFx�s���/�;�NQijw���������u�3�>�|%X��an�Ɖۚ��4�wo�	��|@8�Ԩ#��Wsv�jxδ�&���-l�z�l�g���~ ����T'�*�N1���En��3�\�*e1���n�f���8�)���+�߸�Ly<��+"��K?{6Y��@����J.v#d���|P4�/1�g7ވ��g9]r�;C��bO�Zq".;�"R��:n6r�7�&+M4�UPw���tܜ�]�׆�{��avH໧͢�m���y��o�-$A`uOt>��)����Gjq�3f������a��{2�G�a\�X��b�e�T:��.]J�u���u&k����bp�O[�_����������U��g�xo�yX�f���ieYD1I�����̹�!x/�H�"��>h�A^\��u��G�lf5�3���7v�rT��fؕ���N��7U��K�X餻Ys�nN������'�oO.8�,�H ���[�J�v�+�8���:9�G<�s�wVO�!��3y@�l�Ru|�W=��$���<Ǧ�Z�TK�[�z���{gn	��")��}:�P���y��~��G^6:��+��]�'�\BsW��B�K�<���AJҁ��~O���Y��a'{+k1�T��T��-�d������Ys��`���]|E-u���X:���<�F�#�q��{�Q�۶+)Oa�o4�p��P}�1I������b��g*�+t��^�s���7��i��[\n�i����l�2%R�0�@8��ג��-~���X<�.?��O+��Í ��'��8�[��B��J
�r|B�e|畆��>�?�;�P�K�K�dkt��X%�v��)��|]�7s2+��]��>��)�O��H%�	�l�"[�gh�����{���t�%�B��ɛ���5��8�����u����|�'G��'-�S-��P�<|�
W	!�s]�gu�i9�]�~J#O��`��Y�6
���S�x檈��v`���$C��.��	3�K�=�Eh�|2�9ϓ�8/�My�g\$�'�;��ЅZ� *ၕ0�5�������.�6�z$�`��ݓw��
���oZ�HД��m�̡�8�v�*��k���[��+zX�nJ��z��ӧLY7�|���ֻ��5f����R���i���"�&�t<�;A#����:Es�~bU�KW;���:�6�.Y*��&�;X��I�҄o�T%N��􍈨s^Ȗ}���J���"�6m�G�0TkH����%�޺��绣B+vS	=R���q"�-��g$bƹ�}dw'r�7{{�kC?x!�O�ӫ�a>��g���=�A��WE0�b5b�	�#
|��7�qU����*��y�������|o'��y��ϴ����0{p�fr�Ͱw�ln �*��Ӭ+�f=[ռs׽n��p��6`ya����ې;G �t��f�N�.G4ٮ-��pN)(��{�>M-�=�*�>5�~y��y	�xN/!b&��1ux{ޣ��%��']���s�Q<��[��kg5E��-����zwnyMݔ�K��1��-���	�; �~��w���2���?1\Ȯ��}I�k	F's�7f��K����+wt�ū��ύhzz���.��?�o���'%�PP5�xwgg��A�D�B�����nM	��9�5�6�A?]�[�7�O�&�$=���n �5¬��/Uk�e�Z
�� �K��a��C-&�7=n�_m���]��kV�$�Xa���1.*H��9ݛ3h������G�/z-9ܥV)c�������?����g����?��H[]��$|�m�pƴ���g�;�P�����w6���~h`n�C�`��h�6�i;D��p`�3���s�n�qO�l�+�c����~;��u}B1~�f!�+�^Y���[���5qS���d��T{9�2��i2F"
��'�H{�M��[��9T:G��6*�bI�pT1���,6�Ʒkߒ3ꠦu��k�>j6!ؗ`�p֔g�X�<�,J��;Y ����N��o$f�.pSlKB�*-(6�=�<.�$	ɘ����o��
.��i����>���|i�u33z�L�~؛>ÙUu�%������>�+�0��c��,`��D��C�X����thE{vR{�	�O�jQ;xP��[��%����oX&�y�>�6���[䂝u�|�շyۛդά.8� �����e{6~�b��i�P��������~VEϖk6��҃��j��)�a�"�	�?_r�gN����ܺ��9�C0���ۇ���2�ٚY,�f1���q��E�ᕟ\�.�+a��8��pte���T�nĒL��/3����+!G��y�	�ʫ{pD�F��y�qp�ܬi��0'S��t�eж��M�a��;z�Tw��,�X��W�R����?����7K.�Ct4	���ع��h͂ ����]�r�-����Zd��q�4���g�a���~�`n�eWʅu��L)� rq������OQ�<<��,�'�����ށq�.�1��[�6�[c�'�Q<�ܧÔt�8�����G#�Ǯv�0��a��в-�ސ�ɻ�X�7MF�#p��I5���@��*�$�'a��6�ve�;����+�
W͗���L��cy<� k<5e���0�jN3�y�f٬ޒn_m�C�t��P���s�\��Ο�L�W�a�6�zh^y���%���+���"f7�#�N_	��*�5��^X���������R"s����(�Y���-��*��S쓷tt킄���A|�2���]�ԘP�2_��c�����֐^��0m|�P�9�чt�X���u�`>?E���S�H���	=���,%�g���^��������n�k���D;7\��m����k]'�4:c']�CӪ�9��p�m���k�e�#���t?�?q��:�?b�D�7��j��U�Qw�f"��z���D����ݣ\�\ft:-U�._2�0q�-�%qfe��Y,(W,�3u����#[�Ϣ�_f#�,J�#�>T﹛�����ȃ��͊m�t{(���䬃Y����J�M��j�k�7�wh /��?�x��^]�қ�I�m��b�\�C�<B����c����Er�k��m�[�j��s�Kp�Ӗ7��b�g��!���Mx�0�vt�|p�!�X�y��ߐ��{�ڏ�uAQ�Y��n�x��=�����omq�����<�<��7o�a��垵lK>����3S��[��,,5S�����q5"�0����!�Z�
��Rw<�q��.�Sv�zkX��1���c�����x�ax-遠�A�e���+���͖��eWʅs�������͵�W�{U��|�_�w�N*൅χ��f�ܣ�5���P}BSNPu��59f�}vOFa6���>���7z9u�F�c���|��Hv���}�*{�|������]�kE[px�'o��)�.�xn�C�Q�����+���֡J�?�H�<����#Q��W:r�r�ç}��@M�9
|�W?0�ʧ��1�n�R	
�j�@r��l�@dW�L�E�;�O{�zĻ*��	�6�o@�����/IE��L�-�
)i��W|t���k�E�V��~�.*���58fG�O�u���u�&c��cXA,�3xk�c����y[B㷂v�S�=�����c����̘�j��9��Hm,[-Bԏ{u���[w�d,�\�N���`ٯ�S��_�� 7�uy�Iw�Є/���m�4�����D��ޘ�ۜ�V�ԥ�5�hwV���+��y޳*��dR���-���|�����k�/v����ϪA��0��.V��wq����{U�=������f�W��� �Y���H�_�!ٶ� ���eE�;
b�ʲ��N����Nl#"�կa(��nD�����$�5���P5ӞT�����R�U�>u��ZYٺ%�� +�_l�KI"+�p����Ũ���{��
�79#�}�����۹���q�7)<67#��*�>�>�'H8Z
T�!>�N��n].��)L��νm�؞ʮ'��������=(���*�^�9U6�w��H=��XJT89�)���g��2x�TF{S��ͼ4��S�؍iiA@���sq�ꜥE��}G��_��z,)����>���[��=���b��F���k�?HS�k��1��'����E��q�nӺj�I&v�kW҃sP����Ql5�{2���}�E�>c ���9�UW��ߠ����[��>'���G«m<�|w�8�ƣaf��,_:����ǫ�����6Y�J�=�J����2�|��O�{������7���S��V^pI��hc�,ܸ�\u7(=�zܔ��F�uT���R���W��=:q��:qI�	ם��~���|7�ޢ��>�9ť��c�yU�G}ߟ�a�++�Er۸<�jm-1��������.+��0��Hە������P���H��]��l����ᄜ�����%|���q��D�?������Z*��T��C K=����O�{rL8&z{��Q̺؞�=�R`Z{\��lͫ��)fN�h�/Σ���xLy�?6Ðۢ��'��D6rܞ�Q|}�`�*�ǘ��Ź���m�H\�i���Ь��˹�ؼ"��@OS=��	C�ڞ���{3V*�w�^{T��/C�	T~M'��!��1��Q�����:��w(��l���D��5O�����=V�`�\��箨�|6-�@�ǐ}g� �_t��yQ��E�S3�jR'�%���}}"�x,4ό��	s����[k�`�wQ�u~o9~;��m"��<	������~� ����s4�dT�d�N��ι9
�<�^�������v���N<C���d�ǃ��Q1)�%ɗ�a���o�E&����|v��p.��3Q���(#\�}A)I�9�
Uw�z��S���T�M���n���,�\�%���(�M�wy:m�������U��u�d��)�C�v8/���XXۚ��ݳ��/+7~��P�$>�/St{(,ؼ�y:��"x��Y�y����agR�������0!�3��9T3 ;]�3w�֋��\�.���rK���$��W˚�Ì�jtb�Lk5͎f_	┐рa�L�V���yU�j���a�T��43ǝyK�9��r{��W]Ճ6y�ܭ���ӗ��.������y.	5���u�\�\���t��l�X��u��s�Τ�Еx���YyVW\�Sx�g��wk��K��l}�]Ai|[:����	��
ez���س̌8���*��^�H
�el�:c�e&j̥����-Թ6��͌��s���3RC0�uv1�c7�r�be�ݍÒV7������}1s��5\����%���D�]�'o=M�afQ�!������v�L��8
\#�~���I]}��&3�Vk�s��tG��(�f�a�Ƅi�)��V������������U;����P3�r��u�C�\�?mi|�ٖ���͊]R=ę��P��KR��b7�؆v�\����<Eu�
�x� 3�:�	v��*��J%[۫mS�p��23;ۧ*�%դ/5DkG,@��!W�[}s
V��r�<f�n����i\��S�5�O$�N�bU�Hvt�MZ�.��؟Bƈ�΂�W:V.��rel�;9I�a�a�فZ�e�'0���}�qǕ7t";��R��̾������d����|v��/�m��C��!J�^�Kz�
bM�-�ݣ8��[�XV���F��4�V�['���;�w����UC�(ms��X����S���}�/hٍV#i1��Vꔅ\�����s��Z�Xz�_�Y��t�m`xW+��}�Un���	C5��nn9�*�yE��#��9���Ed�+8���[�:7wA��]��&��)�Vf5뽜L�/J��]u��I�D�Щb0j��4��RԒ9w)}e�{��Ke���DFC���:��8�>5�JW�v�2�ޓM�W�@��}�[W�������Ձ_S�:�1fV�hI�ѐ�uܨQ���պƝ�����VMe	}�w�f[�����]���d��믤lW_|f��?|6�'11����ɝIY�N�{Q��\k"��ofp��μ��z(��&N�3���a-gp�X�.U�-�}:���m�[&dj�R+�WD�K2��|�*:9�sm��VFv\��1,�&�;�7v�N�_Bnh���A BH��Y\���{��1D+�RH�����k29�=��N�����ֵ�k�Z�MkZ�ݻ}�|q��]����32�&a�RZ�AJ4EB�k�v�on����ֵ�k^ZֺkZֻ}����{���}�}�K��uM�[.J���BvV����Px�-�����"�QZ�&$�Yѕ�*��B�	�'!l���f��D�'S�@�kCBȕ���XW���
�|��	aTTUN����z�8w�E]�|�
���zY\�_I��˺�*�Tr���/��r����':xC�y�8$�uJ+u�Jww"�O'*��P8>mwm	G�,���������Ü�<��GB�DW����� 蛺����L����8P(���,s/��%�q.!!q�*0Y)r̉FBe�L�/�� ,���D�-�
q	�b���8�]��j0������u�Oe�\֮uqs�r�	�z%*���utZB��mb��5V7P3s���&цF�4Pd�n8�e��p�LS�l@��4�%�DqFˁ�$i���r�]�n�z���xde��/0ʐS
J�M�a$�#qBE���6̆0��>��x��ds�w:/Xu��ʧ�~����S�N�]\v̔*��$83���~�<|�U������Hbю�q��9�F�^ξ .�hC�Έ�V�u9�$�o���IK�����R���J��$�; ڳ��	o�Z���Y1iU=Mn�a:T6k�qX�1U2D�3�n.)����	��{�l��N-�è��tg{�#J�y�O�t�r��nD�����>t;���ޅ&�����������1�/h�Q��*�#�AǬc�(�Sn��[xulc���f�P����Q�C�W���ҹ$���W<���j���˭̍�Zg
���ߧ� �]�sui�w_�Vd��we	��w���'��0���6�{i��N���]���<�ڻ��=�I��u�j�h3�쥓KT�ot�&�FL��iq��r�g���A�}�a���μ�K|g��-GN�i���1!]wW����7s��Þ�������6�o~�i}���Ɋ�����W�����b=v�v�1����ۣ35@7_c�镧Q�wR��7���_=`��ڥ�}���B��~���1��I�����P#.a%�N7)کw5�ѽGm�UV�n�e��}�����8ћı��q����F��&�N O��wǫ��ת^W=Y����l���<¼E�ᆯey�N)�)�

�w��&���r����Rx��|w+��˞�6�`q3�v�����zC��pj=$���eA�l|�?)[JU������(g�s_���^�ChL�����w�fȗ��նNѽ��H��fw�'�$�cxppI�V�}���tZg�Y۴x��E0�Y�o�6�K�9�wM�I�I�B��.l��QQ0]Ɯn�W�u4�g`��(=�"&��U��f^*����y��{}&)ϻc��okSm�nU-Zi���,r�=����	�\��HS�T��j0�m!��\�_�������M��-_
�/�����6ۓ�:���C HG�1��Ӱt�܌1��j��㹓�~�V�ێɶJ���3��>�Z��7�u�?q�ˢ�x"h�f��)d)�e	�w6׻jXU�h��{�n}B���2-�z�+�Y��D�T�sI�42(o�q�c��ʵ���k���$
0J�_v�ne)Pi�:�� �	�י�ً.q̛n� �|������~Q��F�1�5�;��� TfQY��\uu6�l�h�gǇW�<��hS�b$7���g��r��o�\�]~������J亃�2��u��C���"��D_ZWI3Ǆp�;�i����=Ǻ��@��;�FY6�y�����.��U����L��;�œ�i��ml=�GrS��y���F���$�ui�Eݼ��7��]�7���F��<���UA.&�u��I�c�Ywa�������͍1hR�'=o���i��3i�C�3���,��ڧ� B]�k��v���2��f�x�o�(^q�\e����*a����3�v7{!m�2�'�+��4w��+���;C@7{���v�ye-2X<:7k��}�QE�ɤ$H'N�'}A�{��v5�b/L-��W��Bo�����`̩/��JA@�Z<pR�`���_��ݟS�B�P�����Fd&`�u��#P����/өm��xw#�5�V�ԶU�Τ��cxeu1�t�G;��XY;:�9=�wo��o�
�`�0/�;Kr^5�ξ9�T}����7�����ׁ��^��X��p�DP�
�^� �����3w5��w�if`��f����WC��VªK�d���C8C�\�:[י��si�gW�S�{Gv��>�I�sB���'X�
zQ=x�n�^o��6���n����S�HO�s6	X����uL��� N�n��7���n���W0�5�W�@[����y�s�sw\�%]�����]�ݭ�@ӯM����.A)��=Q�emށ~뎫>0n���.LgI��f/�����Hn�T��%�����At�xD':����)�s?^��5 iUop���bf��p�x���[�U �+DuW��^r+V���M��V�6a� �V�vϠ��Y<�e��j����u��F5�kN��l�}�ku��ı�cہê9�=2 ��=_*l�ltrQ��;�M�i�F��{�ň�ƀ����7�wx��3��gשu�@pT��ݣm��A�ֺІe�F�˶�q3�cG������2�����X��۠���cd��Ҧ=�<��8�m��-Η��97-�x%�����f�@�,�'UG�r�|ȉڬɒ��v������d������������3|�U��5�������{�db;<�~�R�L;p�x��}]ES�;�}�׺�O`UY;L��;��t�!r�Yv��WČ��FDW���d��il�@$M(�k6Cop�xSA��/�'��� w���{
�
�R�����I����x��h�m]���ro��A��w��3���F���u��+���N��N>Z�>���kQ�wn�@gn�z7D7��P2�1�{�0`�\��rC.E���l�;z�QS䐁��v�g�c�,'�p���F�L��5zNa�=��y�W�)]\'������>��3�4�𛫹ޝ��j*�3��-w�>�U�~�=�Xt*O�n�ܧٞ�Gb�]+ï��a�^�L-��v컆��(#�;�W'���P%�D#�Y��jqq���%�٧�4�A�
�wG�yn;F���(��.�-v�byUΓAd���F�V����ѯGwIޣb��ԯL~�ݸ������/�/i�nҐ�%�H�g:n����D͖�"���%"�:y��^^���w��2��wv�B�T�XyB�n�h�,�a��s[}R��+�^�8����|���(��\v���eW�/�rܜ̑nuȄ:���ɳ����&_��YZh�$�E]�<��+��	hm���j�S����0��S�suro7���Z ;���V���;�z<s�l������d�hrY+�o{+:�]u�a>���/8����q�u��^$�Rn��N� �h�� �n�~Cm6�ެGW�L�~9����M��7�r����'���^ݠ���#)@��la�u����wYg0�����!s�G`0T����5�f�{���{�w7�^Ɨ�����z�������i��:uI ���������M���4��(��'`�)
�a���y�[��4rg7�9uGR1M�-q�;�z6ΌVQ�1�h%�:$�*�5ڇ~���W�������#��E��#��3	�����H�����-� ���)�릾Uh-ޢ�-̖]e�csKj^t�5�Y�������¶؅7,��M���.<*��҆l�<��ck��B6��ޮ���q֘����1Ǒܙ��b����)-�2�p��ԥ��Q���<�OQ��>���9�6�c���yyy VgZ�o}�7�<.��jz�ww�}p��Ԅ�G�oo��&��9L���f��޿l3�0��|���������0��WRw�����p�W����(
e��G�i�쳡N(%`�_t��=�^����P�0f!9N�^%�w���]	\���EM:��஻&�:P:ױsZ���5ƌn?�I���hCda*H�?wKeVKtK8��6P�;��!��D]���TI�RB�^\�uqe���RUy.���Z��w<{���ۺ�O��\���2^�&08Zc�E�djU�ia�����>`6�d*]M7��1Ws�'���X�b7&4�َ�o����5~���wt	fn
Z���z0�m��o[J]1|�)S�F�.�'gs}��W(�m ��,�.���W�D��^�R�:3���,/ݧ"6��&{�����m�FΗ��V�Y�R�b�3������kmsD�}Ҩ�l؃u���erY;��&�w}��c,3.���(ZE���[�k�*���9�{��F�^K��:
���a�4��i��zV���L+�-¹]���������8�����}�dկ�
�k� �hu9��]���*���3;��^tO-�Uܩ�ܑ��+���z�(4d6a����=�'b�vDN�F����,)�a�q��G��e�e�dM�d�u&�V��.˥� ��d�͢p�/7����k���o�W�W)���P�y��Γ�7�����&�;�(Ù��V�RY�y�K9*;|.h�����2��L2��ط��g��8Ur���EP��0��>���'w�i9���f�9N�Jϻ�AX�����6Y�A]�MUf�z@�ͫ��sNi[�8:G]#æ��o����R7�V�{7�WK��,�E�tu�u�~@��S�]�z������oի"�����v��l��Y���N���]f�o�C.�c	]]AwuB��cˡ`m�����]V�P>�QJg�����F�ХT�}x�����vcFmc����㼬O�j�.P0�u���b/�޽�(Z�
kж�z�w�����2H9�h܁��w�o�����m�����l;սY{z������y��p=��Q�îռ!�K�/����t� b�훷I.Mg�P�W��Bh��	��wBx�ލ�3�<o[��\�tV�޹&{���P3j��	xe{����-/hi]ԕ�ln�î;v��6=�u\�"�!������M"��$�u���K���-��F�A,a��õ��q��FPlvO7�Oniی�am��Պ�����g�>����`��=�������B�� ��hunAoK���&��`��{�iWO�'��m3�!����ź�<p����������}�H�Q��;Y6t9W{5�ln�� ����nĜu�k$���Rdp~!�l]W9�Ֆqn��5������XM:�u*{�`7IXݼ\E���8H7�\�pƖ��@�5��2�zXY���b_��}���;��S�͌'v./>�= .B5A힠b�O����K�3L^e�@v�}4t.]hao���h�.���v��W�}���ƑdL�Wq�=�u�I闉Z�Kv��j�5�z��|	HnR�< �������~Mx�*N�ʷeLZ,�4�\��P�9	2�F�n=���a*:`IL�sF]��Yp���w���?��DN]�8qz=�SU�����Һ�h���ӵ�g�X��5G�'�.*�]n�5𪇪�{[���.��K��w,i��g��w2�um�r�p���0��*����aTw�sx�y�����5�{{�w�v�p����y�����#*�����Q�x��(�}����)�J2�۶�i)�S����~�s$]wuz�˲"�Z���>l^db'I�@M��wu���)m��5S����<�i�0�̵�8v�d�̆x�����Ú��9�\V1��M�cKv��K	���a��(�[�����JDf��]t�
�U@�1*뺻���7O��[V;�[Y�nF��(�A��C�ip�(�a�z�o���J��U����ؼ�U������v`܌��7D�EnNCp�`����>a�=T �M��u*BG�|�<;Ew�='Sz�l1�K�L���r�U+^h��έ���GW�ܥZ}��u��*i�� �BVIsf�\Yne$V�9�YK]L�Uj�	��Y��:[�fw;�f����f�٩�r��bŧ�M��)�[T�6��p
a���7����Nfv�wZ��h��u�8���1�p�jDv�p�7ۼ�̈e*-���{V��x/˭�������t��P�b��o"{X�x7q��=�GtЖ^���8��ΝجYIe֊��Wcۉθ,h����O�໤�q�ukR�o��w�L�q8���kv����}�WE!gT*�L,keq�Վh�V�v��s8ӎ�-
�*�A�7u�/ec��p>a칱p��;E��ڦ੃�o�����Y+l�kc�j��v������X�<�P�b4��G`Ē��R��}J��ݬ����ۄ��/U�̨i)�M)u���j�ƭ%��@��/N1hu:z`����ޮ�VLL�۽.���B��+�ғ;O2ܔI�lr�n��>d�w[�r��8�Ւ��d��mGqGA����N��e]���/wru=�5x`�2�J�1��O�!�x��xX6�˚=��-�Y�X���W� �{%n�0�u2f��r0�7�&ЕE[g���vM�Z�(e��J���`tk4���M�iG��F#�OVVk�ŤM�������m�X-5ߴ��/�Ӛw$�p�%)�`�ź�P��s���A�R["��q��x��,>��.��B��h[�����h�b�u�:e��g/���u<Y�e�:V���*=5%Z�嘵�k�ț���/�TʬN�e�G�	'�,��%�N����7��<�|'mwGM��vL'Gm�v./3ʬ.!B���;z�����̬���Ϛ�ă��v��Y9��f��F��껢*mԴG�F	}�P���I+�r8��n�����Mʵ�	wDk�m���}}�u��+׻����\�ͷ��J��=80��mK�t��;���Nt�}J+�����3h�wJ�`�͛Ǌ�FΧ����6�����D3���R��z�t�.��i]�n�Mw�� �9����S�  *X_| �C�d�x�1���p0�:�4h�ȵ,��95�:I��&���u����b��7�����_k�#U����w�e�wJ�;�P�gf�B�.R����[f�.qe.]���v�Ƚ��j�b�(�5b�{8k����،Xj��؀���rer�NͰQ�/&�h���k��J����ї}q<Oz�Y��J�\�+[�]�Tsm;$�r�ń/���x��2�á��j~E�%Q�Q#��v���7�~�����kZּ��tֵ�v�۷o���_o�#����x���B^b����L�Z�Β�:��#	�÷�{y{{||hֵ�kZ�ֵָ�v�۷m|xy�c$�y�g �t~w��b�U���!��ȩ0�9@TIl�L��PC�T�i�'R���^W���'�L~��\��z�9(Ԋ�EL���*���C�@�4(N�	�&�.W֑NO���9TPQN�,�@D��Y�h�*�Ų�A��r��.�B��&��U�C:UM!
L�Ud�y�'��w��\�(�.�.�l�����Գ��!�I��W��Ϣ��|��4�����{ݚ\F���(s��ܾd�k7eӭ 9�3o�nc�aA �آ�7����^^^�����.�7�Ŝ0�_�kc�kgƘ��AhCL8·Q$��psHܞ�^�c��i��t�oUj�n��'s�yJ��D�K��ɟq6�dJ��ڧ�{م�ϊ�q������e���	;�q�ڂ|Kz���cmb�:-�����C?��3|�A��@�ڈ��yt�c��f&�5cYgѾ���@Xz�Wn.��jZz��y��C��ƶ�ti��S��b��K�٤C�ʨs^�w��V���S<�ƞ?�m^����eMw���^�Xi޵#pz���ɓ�}�ǔ�Ɍ{[���Q&��J��˪�O?*YU�4�i{�Ȼ�&�E!��:/�mL���8o�na��(�*J�{�;����F�t	��n坱b'm�e��eٵd�R�t���zI���= wq��R]NhϚ���4ȝ�<�ii�j7U0Ħ�ڠ�)�gkKJr;�PWls"��� ����j'�u�&�Y"b��=/�lUcKr,{��Eu�	X�uݭ˺��S.>#f4-ѕy�j�rN��U�Y�]k%����6X����܊��D8�kh��'�W��� Lvjw=���}��yLp�ϺA��'��7��[�۶�nf�q��n�3[�%[psS���q�����6aI�x6�$���z�>�u�;{��w���l��+�kP���r5�uz0��s�d�N�Gy�wLL�i�ZN��	Q>H�fbV�!��1va��q�Yw�T��R�$0�of>�����w�=ZW�j@w:���d��Wl���,���RMs�P��OA�J��$;�A�%C:h�����z3|��h�m����P��.��[�?o��*%s"%�&���t�
�k���[`�L��9@��Ei��zZ�ƨԵ��/�z�d2��=<��ǅ��l^�'�n�L����J8��1�*�71nl�=�)��2Q�=�����W~qwF�O�Fv]Z�s�I=�W�{Iz��b��K8�a�������=+��$���'���n��H#�wX߷i!n�bĮd�Đ������f�Ŝbb�!�WO��;ĊH�=�����IeA��m�K�����,v:"��Tc%v�|1w	9��}!����7���Z��sf>����(Z��yyǟ�����̹����z��F$֝_goC���m3����	��*~��Fm������`�����"C���3�ۑ���_
�5��p����]
|����d��u"��PW����ۉ�nr�I*�qoLa�t=vKb	%ǹg��y?�N��M9!�}�\��I�Ť��󼹜@�eN�Vh������CI.��O*���qz��;�";Ny��@o^��ºu �a�o��u	���C0g��D�8�W�jٲ�6�2�i�6Y���x�~á���e��w&�S�E[�3N�\$�̥<xvu�l��W��8qmp"��y�QQ=�*x��-��6�ě���g{vq���ޤ�k��a��NX6KA���7_L�Lyu��R��Ud��7��ݖ���=;��� E�C�8Ҧ6�����_{i"iF���u�K��Sv�a����G:]dU��O�V<�2��+s��*WF^��H��ݵא���U�nt��P�4�s�;�#�Z�8�ȬY+�u��!�ۼ̦S�:)�T)и�m�a�{�c�|f��z�nv,UD�>�!����V��knIųk�6�\x��y��0�98��e+��w/���l3o<��n����,�nF�)����X!������Q�4��Y��Q�;T�ArA��� ��f�xd3�1,�����bpM]{F�*��ͷ�Y�.�^}�T��!!�h=���u>��py�n�U�U��1�V΢/�ϙ�QW55Z[zB .��P>�0�`=o�s_�^,̉��n��8��R�c0F|�s����O��iwSW��1���i��v�j��^Ҽ���E��3o�����X�w=\���`W��1��E��:7-\9���P���ʸ0e��
{�n�·�3�]�(.S0ԝe��;$���^�P��.��*��q���Y�+r��1�Ɍ7c�q�����%hᇠ�W����7���M:��"�����o��JW�-�Eƪ�ޠ�ߵj��jB����v�8;;��h�L�5�=�ء���f�U�����PgFӘ�@zӾ�f^c55� z�$��5�IS¯2�.����o��x[��f�i�t�3���>�)�[n�km���F:�?{�?]z��p�*��XToC��O�e>6��%R3�Xm��M��ω���P�nbG:eo&P#����J6v�P���}�;��d�B�}�q�����f,��F����jA���d妢;�G{�����D�7d���m��f���;�o:��⏷e��u��l��2 �H��W'@O�C���G0�:Yn�s���(��4`kg�}nd���i��ê:淚e��v�uF����b�U���[aU�p���J����4@�^�+g�\SK���q^�br���P�(��H��p�W�o�Έ�=N������Y6�]��s$:�6ϠWX���`���4xf%$
L�N���-���$�����]P�1x�G��Т�"/�DMI����/5�H=HR���v���&�
���F��p]}=��8�Lú�UC����F:��������j�W;�e)X{n���T��
�,li%�HJ��bg+ug�]k��@�}4��5Mz���Z�8p�z��;��=ߧP��e���=���U��W:�.�f{��.�r�}���V�+5��ĩS��NW�����ׯ����+�SL�F�:EY���6ו�sN�e��*�&.z��i���^6A,�$��zHn���˫�'F�-����*����6Xt3Fs���SmNqՊ�O���5�� m���:QoGg���]���T6@�?����e۹���ci^�#���Fcz{�%=`u���{��V$���h�2�x/��	��v���u��X8U�w�������Ϲ�{�r�c<�&iN�C����0`U(Wk"N�n���f�nc�=h#���E�Ro�<mlX�c|1�uFkEiGV͝/�>���.�k�)����5~Yr�~���r)2�%�k���ߧ4�^W�$�U��M�p��;���S#��7�|\֫��D+}M��P{��=U�S��;>�8�!����6��Oh��Fk<��d���l��	�*�����J�=W�7��!�T�{V��nr2p;��R�������l�񁻘W
�I�Ӯ�췗tt������W�9�Њ�+��;s2,V�-H����3݌�@��&��I���M��G.E�w5x����N��f�\li�D��/O]z�~�Q]%���b:Ԍ�M�ҝ# ����kV��'*������*�2#�]&���_-��I�5�L7T�"!b�5������� ��P�֪/�l[�n��n��n��	�����v��W�SA�]���������4���vE\�z��&�t�_ZL������ɨ^�I�u>�ga<ß�U�FED��;Du�yU�{�wh������ҤV��T����ܧ��5eO���@,����Y�w,����קg�0�>�ɾ���c�:��JF��̛�u|��3f*y���l��������x=vKbW����z��S�F�e_�%�»6�n�9��[�x��=Ԉ���h�Z;��0�ʛ�:3r���q����bC?A�Uq�hܺ�P��@r#�/�ۅ�K�	TM칬�;�NTU�dR��(�Ą�Kf<{m�uá�"� ���g{{w��ōFH��ܥ]M�j��\����,dc8Vl����s����)�u��r�;ӽ�T3)�]��D)/�͵ϛ)�J�M#��hN4�x�v�	�Λ{0_Rj:�Y�%����q����P��1У_�������~|�5�'^��S�_�Sڂoe,k��=$���v����P�5���^�R۬9��!\�F������6����{X�{[� t3�lk�,�H���	[h�f�0��[��Oѷ����>��R��ͧ�ӏqmw)VgQS��Y_����8�R"}�j:�V�ԉ�c%�:cq����޴5O��>c氌 �9TȪ!��Iν�͆�fY�K��'/{�C�R0ҟA�Y�7���h ƍ�CF�_�Ow���S��ń\_��f�<��9�7��]� �������P_h��ڰ�A�ӷ�nG��f�����~'JB5�9K^����Y��Qk���y�w�ҽ��ݯz*榩rڽ!J����2/r¼{c��f�_kuj��\e�pנL �RhE���Y��볁]=}��Fh�N�=k.{��F�83)%���3#N�N�ݖ0�<���J���Ԛ������M�d=�E����ni��hx����(�nc�1��Յp�r&E�� �5$㫸+�����}�����.>!����-�w���ϡ�l�_1F��� �9
�:���Sx�6hUq���Ǩ���34��
��H�H3OL���J��@�a�c�=v��'+Fr��e wWr�󤪟/�rߎfzE�u~��=��Q�ݒsA^�xn���N��{��1���H���N�3�0�^\��r�é��<x�%�qF�\���~1ܓ�c�M����ڌ�4�n��H��q�7�ruH�$r� �F�J6@��T#�u�\�{�P�֣��[��n�a�6S'C��Q��z����Q��U�i�)a�M�M�{{�b��l!��ƀ��6��D�;Rf��|��:��7��\Dq��Q�	wIՒ��Ѷ1�a��g�=�es���b6f�p�={�6���'3���v<�!Pe�F���VXȪ��.�M�WےsXm�C,����裂��^��|�uxث���n�Eϲ�<�)활~w��@^�Q-kygA���R��ۙ8iY�!*Ω-�(WM�R��Ù��M��횥���ӛ;xq���j�����?��&���z�������?��e.T	�! �R�	3�V�2�0�l^O�=����`���>���U�tc���yt���@��|�vݛ.L�=�9|}{W��T�3���J	������!j�"�bjMz����y)�8��t��L�h��>l�������P�׏T>�;��2r��L�U�E��ڛ³s4�'i����JV$my�ٹW��Y��)�P�X���X���vwI�9����{B�5��/��z��[w T���f��q`QO�s�Ѳ��� C^��nU�nv����o�6�hkAJ1ʼ=����u��0mz�e�w���Q��+4��]��t��rc�,m�Lwq����*|R]fp�BcF�g�W��oM9�:���85�$F��O{�{�r�\�lUX�Y�.՝å� �TyQ6G1���
�!�>���}B�{�X�eW[9O�H%z�F�EUd��ͻ(��<:��Zk�g��io�¦�wB;�=vV�Q���b�u��Vq���+�����ڧۨ^D�6|�-"h�gM��^L#�jD�
�aR���m�\K�w��dT\OX�7��J�oKd`}���7V5��j��ػZ�2��nZ��־=ssar�`��wY�mL*�pD�a_RSR	��h᫾���kp�a�-vSC2�6S��W�0�a��b�FE�E��|6�+9M�⭇�9�:���h�a���FdR��Ut���s��5��oM�.�Y��`�.���i����лj���kh%����\�/+�Z2��r��m�xnoS�*,�\��ރ_$��2nV�[�o����^�OM������Fص��:{��Za��M2�d�[x�O�{�w3>�`���G��ta����yB.��Z�J[��n"��;��k8��Wod���}i��K���&<�%:U�mm�L�N�^d���#��*8(�P5p��=]pw;3y��[��t]�%fR�s;��L!Y5ki��
�x� ��i�7�gfاnʏ/.o����J�Pv*	.m*�G��r��e����-�|�LU#�������r��;r���7+A�Э�wU�^��;֏��*��������W�/EU���U��+��W��r��2��sx��o�0}o묕���QnqlI$�,h��h#`7�ޫ|$�RwCz�7A�X�y���HJ���<�y��ߺ�C�S�ږ��wӘ�m�W�E�s7)�G�9�W�����GŲn�����Wa�̃�]>���ov�����T�r�Ea��K�|�Ӧ���$5ׇ;6h�u�{'Só;+/]Zꆭ�*]����L�Vi��f�NU�r��DR�7S�h�ȟ�{�Lv%��8{��; ��kFd.Y���˼!xu�c���Y��c�9bq��fXc�^GxB�%\��	*�d���LN�&#�"PKUZY��j4��k?�{�YM�Y���:3��6��h�������]��샑�7jZ���W6L	حԕ����4T��s
�ª�q�d}�k��5AR�b���z���19��aҲ.�T;�)����b����s�:�����5�eo35ޘ:�э��f�mp�zʃ�s.L`=i�8�C�k���[�������ff*N��sT��`��&;ĥ�u�����m'}�S�@!U��V	���u�;?'��쫺M�����Vm������c%>�y嘳EoRX N8��:�r�//@�]�݌�%<�rI��f!9�**��&��A��8lI�H��J��%�6S�%s�<_��>9D�$�Y&�L��|ݺv����|}4kZֵ�zk\kZֻv�۷������5��g�9!L� �T�u)���?f�ooo����5�kZֵ�kZֻv����o���Z��Ȫ�/8��T�r�Gt��H���Ⱑ8w��H�5�iQc7F]���d�3C�N�w�xEv}J��;�/��}L��B�#+YA!c�Nr�sNr*��9t�77CL@U+�k����>p|U�:,�wp�D���+-q����x�k��<
�%�����9�̜�L���紻>�V�t��0�P/���'����R��3:r}$(��г���_Iz-�H�Z;��a�S(Nk#���KH��wE�1�� Ƌ�N'#0�

$�A�T����c�d�$!p���@m�Kp�
�xsNk�H�k"���%��P�WQd��gU��2n���{Csj_N-=�m.4��kq��yS��v{ �=	�F���[p4�p�J&PJh��d����D�=��"���Wp��tzS���s�����;����=֓���R�#�@���d!D�Afq��zx;��>8�yOs�߽��Z��L����]��Z㔞L���v��c^-ԙ��mf>5��^<Qݠ�*��OV��$�@�1�u�Q�q�/#`>zo`����w�[�RԷ4�����r�y���g�J���q�@>��N�pur��`ຬ�:I�4D���"df�=�GrU=7�3^������"�"���$ya�1L�@@��}+���}ܢT�El�Y�i1}�w��Z�quH�#K��@��r����\�������337���e&���8`����I��VJ{ͼ������B�����<g�x-�������E�m�I۴/{O�$�h(>/ ӑNdd3���N{���x�D�0��'N�{�p����f�	�Z=YJ@ا9B��8[̊�3sN�T���a|������F�Vj�C������j����e��S����r��f�e$uX�h�T�[�q� �;(#äR���Ўe��T��u�"3*rb32���Le�ùi�[ ��.��?q_	'��~H�3�M���}���g�0��zZ�I�b�B�Q�;�ƃy���W	��4s�;�<s92��(��Fv�윎t�� ��x�pb'���h�o�������Mʒ���9�CE�"|L�	����|ڂ�	Ouw)���
%sg��%��|�%{�?+���WΪDff
+4@�[-���]�Pڌ��I�H���`������]�i��o\�X���~��D������dϵ�N�I�s�J�M�E��)R��n���M��c��;u���n�21S��ׁ�˦�UǇmv����Kv�M�Y³�C
��F��Z��i�"3�B���;}���˺+���Ƅ�1������{��Y<M�wf���0��a,�o>zAWLw�����A�:�T��͕UIQesչ�[�g%xm6��`���@�S�ۥ{���l����]_�^��=K�ʆ���ݘ���ߘW���+�9��;"��=�f��v��`nF���:gj��S��0���A�����&yF��������x�tW@.��a�FX�՘��į�^E/Iy~do79u�s�F�2>;��O��&|>0�Q�R^Y �;�ۖ���^�������٭��/j-��I�6�.��y�cp+�[��
c�[�^^���g%'D��u���¼<<b�1��{���jO��	H �8$϶�㴊�f�K�Oh��Tr�����<SxϢi�.���t�E�mqz�Gr�^l�sqIUn�! D�H@s]�O�pM�ȪQ�/HR��H�!�K������;{�K(��ӽo��-�&��U%��m�q��u��l,- 2Kӻ@�{�����F��{W&�늉u8����	�4A�ur�y��beZ��9����YC%j*iU�G��9�f�o���挸��7j��;�,��[H�pp!��[8��_�Oww%U���ܷ㙞�z�M��s8�=\�^�4��WRB6�n�r�1��3ҹ|�u�E���3��?���o�����N �L�X�6��h��nO?�����lt�96�FЫy��U�e���'��6=)��!�PW�h�O���N�V���bU�/|�}d|k�[0��W�����d���5���7�M�|9�������=}���Zݱ����N��5��7(���v	yљc����g��Dx���Pƫ$��0:چm�6v����Ju�M�c�Z4��U0���C���7��VoU�ݵ�k�K��S���~c��}�5�J�F�N�Ӟb�3Lܪ�8�N���ڵt�V�{ g�`�f��@p�fr.�n��#^�_���gfoI+�d�5���Ѝl�i×�6��ӐCE�Od���D3���zH��ur�s��/xNǎ�!Pe�`�ĭ��|�3^VQ'Hv��j�f��|����W�'�5��6��F�\B�9����y�ڑf x�U�V4k��y��R.��w��&U��ihW�س��4����7�G>׸b����77��\R�˾OK/�N�|�ț��;��KU!$�i}���Lu�Cu�����kd�T��*Y�G#���=UzWR����,�N�pT��v1ٮ�U"�٭����z=wלl
8�U w���OTr�n��V*���r��VӬ���ё<��e��C�E&7��7K�L׈��S���{%�Z72c��D�O�߲�*x�-��T,o[����n��sD)�.��ݎ�.�N'��!�\��I� CýQ>�*U��ӷ�]�Q�؊����o7���ՐΈ�kz��L���v6�	�c�+�ع�Y�@�7�a�Wi��ݕ�B�uGWg��0S��/���/���cù>��H�P�����Dl�[kSK=�od�v-[mHig:�w,D.�QB6ʐL�pO��#��,���r�9���& �#��0��f���u#Y¨t�DhQ�=�m<{nOu��:E��ݾ�ٲK���U���Mg�>�j~����,|i"�����iȢk^mUK����}��Q#��K{���0u��C�C����ܥ�ݢ���9F�/��.���\�z�D���:���i��4�k�����w�ՙvQ��3�za��D(�F#D��T��$�w��s��]jװd񷍙��Ĵ�|��l�kο@ˣ
�;'_;(�k��&~nj��{��giy�"M�UI�ֹ�Y�r�<�m8�Օ�u�\��|�@�龬5��{6��(V��}A��c�0�<ͪ2�;�Ռ&�vM5���>�S���s	ͷ��!����lī��������*�BVބ�չ�j�`)@��%|)�]��vq�Sh^�^��:��_G׭���
�Yx�BĬR�fn[{w6��� &�E�覫@�UM��ҋۧK/F�q��A�f��7���;�IGL� �����o@�Z
S�s��~`����J����,�n#WW��m�ͯUN<�c��=hb-����.lgz�2'jF��Zvt��,�jŕ Ua�Z�IU�^�Xӛ}7]�jݞ�ba��pN�4n�:i�q��=�ʴ�U�F�fC����]
�A#���[�YW�r�Y�/w�/hPdE��ݝa�b2O>�_���7m���rwr3Vm�{�L���o[��g�~V+4F�ފ~�f7��)�*���I|���^c����^s[�9o����������;0&k H��<o4����K�L�߄�]���l�4��<��}>�;0o ���Oіn�{N��;�R��+^_)O^n�m�m;u�tb�J!�F�s�̩��ӷƀHUG��� �H����6���q Nw�=�e�|P8�b�|գ���JiE���	B�1Q�V�.̫��?v�@�/����U}���@c��6Jg������h i@�!(��D��`�D0ٟ>���(�s7���^�B��+u�rv3����g,�f�V#�p�nݣ�nv'���ts��~��z����F��[y���ǟ�##��gcMQ=�׺����;�x��xw�=ǫv��g��iXvr��Qٱ�w61U`R���wX擕�N)�N�XA�6�����-y�D��vBM{�V�cl���e#E��<�U�#i�G ��`��)�h�s���7ov���=����zy �{�-O�������7Q��sx�9v��kB���K����}��Z�8Z����/�O�GI����w5�9�&Et=�Us>�W%��"�����d���d���m�vn,���~�0�,s��joT�F�;��Te���_n��fn{^f���'n ������GQ>ɹ�S��~vS���\�����a��[�x擜چU¦��Bꠎd��^ɏW��sŅ�+�dH���,_xZ�j�"�8zO)v�E��[q|�w�Nݚ��7��2�(���T��M���1܌u����i6׹�l�&S�7/���f[�B�J�����A�y�ƋN�q���[�̮yJ��xd/+��¼<=x�O�	M�����m�������-���{$�ώ��7/m�y�6��2��Z��tzc}��YB�`�1���zW%-���QU���'V�,#�}�pp)� ��I���}�=��7�s:_^)�l�j�$�&��2`� �������(ݾS���鉌�S��F�����Fp�}���ě������L;a�{t�B�6^ڵ����Al���:wN�ZR��a=5շ�}Ri�ی1���ڬ�xf�tw��W���7S�Ep�<��hH���0�l�c�6��.���"2�ƫ�����3W��P��'8�.%9�xV]x#;^ ��IHd�a��%�ќ�p�[H]A�-W�|�H�n2�*�2���	�0�R�ʺW��5�dd�]�w�`f`��9����j���p1��	�H���e��z��?�������`\�R�¥��Y�u)w[�,����B*!���`!�2�����ou�5�����`O���^C~��YK,��oj'Բ�r_vd�,�훹�"�K�؏u
���ec�����h���/��`~���+f[?.F�k���H������)��8���O(�L����m$QhsB� ��Q��Wu�&��E)y���Y��^��kI��u����4���)�s�łhp�绔���������r�t���.��w{0��z������Z�\ө�g�>����˝����P~��w�E�fxvP\zE#*�#}�W�t�^�SøI*���p���1��T���X,�uku�@`�c/��b
Q�O$�ǹ�)�]l�����٣��7���L��L�:��c��XPL�u�����bZ&H�S�A�t��@�ޠ挀�N�n]y�6�5o��zL���kcoV�1�[Z���}�U.�g�_�h��m\8�����wgS�r�y�决w7�8t���ؒk9%a�$�i2��k���Y��g�=5�n��.uO��z�UD�Fz���{���M~�l
3��[]Oc��5<g�e��0_g{��@H`��$��\�9ܓ����C�1q#�k}}����;�����3�x<}Mp�L���(@
�$`��W{�5*x��$ �-���#k���"2�Z"��JHM�'CUTA�w����<�ol較�{����y�ޘ��PF@��]�T���fXͥQ&n��b;���o�t3ˤ���j���&�$�^Ya�۽�w�_�^�m�1h�gm1�C\�n㻆�;�^ߠm�G���r�,�X\h�1Yts�	�[�ǆ��"�{g�E�l4v~``��W����6i������Y��i�����n��h(�X���.td3��a>�,�̓r.���խ��y��VɯYG���d�t���� �>{QsΫFS75���5Jo�Nn�!��iX1�UfЎ�"� ]�Z�=�;�G�6:�y�/�S�S�;�vح�t:�-�\\L��"���C����\��)ʼ��b��3of�3;+	�W�r���>��3A@H ^��c��=vKg׆�m{U��%�4�CI����β�u{�"��~uS������.᧫�c�g�
�}A��8#�Jw<���`p+���y�:�ݹX��o{�d@�o.ꆶ�<�.�.��V[l��6'�n���1;�����m�h_.�L/V-�*��WA����A��GpՓ�Z��(�nգ��xV���&���2���j�q�v��-���5�[ɜ��(�zu�=��[OhG�A�\8UL�	�dax����-�>z���ʎ���qW�	�NM��*�{����L��-�vfћ݋ه�����H�v�7-�UyS����	~��d�:����9��L潜9l*k/5��\�Y8�řC10jq�ٹ�p��1�V!LP�R<\��5z!�ag"�[�NP��Vz-�K7C�����ڡ�2�ϥP쾊+V;T���F�8[\���'�;��Z�`��4N���U�f[4u��Q7];zL�]m��3u�;�V�J��r���{�*�p�U^��ژJJ�B�t�e���8�ds��VA,JAZ\���c��K��k9�C��X��y}��k:��v�W�[ٓvfHm�w�C�³�[���^T�6�S�O�"�+%[-��z�z�v�T�wgv=�S�-�^m�/R�Ng^���ɉl�ڒTR�:�J8$��{�9{P�qU�5��j����gJ��^�1gv|<�Ψ�n՞ZU^�l�պ$�E=�V��6�AoG�K�Gn��:w&��$�Ȗ7T���nfli��g)�eI�j]k��ge�L�� �h��O�Il�C����U�����j�x�p*�����-�U]�J�4I4\5����/�t�y�۷2u��&N#��)��_�u1��l����Y�gZ4c$�+w�;��ڼ���2ڣ�E�m7:�a�+�fz�ov�o�2(1N��^+��Q�Mk'^p�b���rS�j�]��O��s��/LΩg�C=�P��B&��;���b�%��������Od�yՉ���b�\�wE�VK���s�:�ړAu��Jʇ)"�.��M=���s�d�9Q�iD(��gx���!f�a�ގU�E�ě�|���rfĀ[]̌λ�a{Ou��x#�;�̊�+}�vR^��p�NMQ��9X�}��5|��ͺ*�Q�.�]�%�\���X«Ǟ5hv��a�W7���Yt�.�F�c�,v�i�ꪩ���ʙdv�T��r�
�Rz����j�y�.Wp�ـ�q� ��m���cw�,\6�F�Vwt{&;�2njG8����/u)w�d�K����L��R�q��z�@�T
�����Ҧ�3��F�y�9�Q�q���BR�Z�36�VM�l_>Ͷ��YGy�vA}ۺƄh�.��U���Ȭ�ӊ�XԇMLޘ+�n[U���o&��
�fbtr�E2(��+��(�
����w��_q'�Gդ���*�����ݝm;|||k_��kZֽ��kZ�nݻv׮��B<�H���MN�O,,�\�w/9Z���*��Z��v��������kZֵ�kZ5�k]�v��^���HBf=d��ޖK;��� .����[.����99G"֝Ԫ(v��Ny�|ɸ�K�m8QB�6C���rr=�v�E�®Gr�J�i��T*��_I�
�VL�U7��be��]��*Wih�$tu*!ʕ�u����WT���yRg���;��~w��E�y;��݁E=@z��~|��w�x��;{d��9QfWrO3.mʢ�/]�9�y!�;.萗�����E+KD�2H�s��SW\<���ʇG�^�-D��^KT"��Y]%��f�
�^�e?K��E;8ᵭ�{�GC�.��ޡ����w"+�仚���YL�oW���ؾZpj��t+���xy��3��R�,q�h*�.�������z�uϪ�~�
V+���Y�Q����W�;�&v��6ʟx�V��6�(S��o���=�	va<�	�:)���OM%Y�<9�Nag�O��E�5F�̰�]���%�Se�>��u�_wo�y���$,�3��H�jqysp�~Z��|Ժ���ۡvj���p���������9�n�G����N#��ܵ>��Vm7�++����zg�#6�a���w��D�2Fy�76�Vi�\xy?G�ԉ�S�v�|6�l�m�e�r����m���|;ۘCb�[zw|_g����k�ʼ����Z���Ƣ&�ViY�=�Ě�n�S��m�����
��ppI��Ƿ��ynh�;"����\�K2t��7�y����udt^wyH\�{QkNe�ngc �-f���^���ª��њk��8e�O���iZ7~��$�㡋@�n�w8��T�w���؁w��T2�z�#z1L<�ɣ�QM�蜤��h�P�j�n�
A)��}�D��^�4s���r���"N#�XWюdpoXQ��*�U��8�o%���nMN�e��Dxf�5њ�o<gD��~��m�]��K8��C�<�Rj �nOGc#�>#�����go%D)�.�W_����`�n)�q��:��(���zLN_)(����lѾV���2�B=U�̐f��8��Ůd������{��{"\�� 3��l�O�@�\�)����~ɇޡ�ڡ��l��[���O�=_�8#l�r�=���yrYb2w"��j̏{'bz�(�"�gvg�~� ��g'��~�"�O׶]��n5Юy&�LS��Mj���=�sr0q�8ipWG�1J6v�V�a�\l����yx��N�dv*�r_h>-;�Cd0���hD.�U�#�/�����h�w4�a��$������OM��
��Yq^i����%Eδ�TŬթ�X�4�킃"�g6���ޥ`<r����HrB�5NbeJ�vP�{d���v���R^�Ux2�G��.�����Y躥>��}{[}r1+q��t�>�L��}B'WRM�G���'�	o�)�4?zxxy��f{V_,\3Rk׹>�=WG`�*عKRR����32U����TGy9�����v}�&L�w��D�X�(Ιc�o�oPm{��r{
�9����>�Rr�VwNg)�����6�V<�3ۯuI-���CC@�t�K�ǆ(�(S��J�;�N�+l��^�U�p�ҽ�MgS�jE�J�|�f��=�j��Oݳ���a�L�0gs��]ø�{�Sz6%��g�-Xy!����^J�8*7%U�¹�z��t��E�������M������	x�8g%�*�bNR���%�J�3�=�3R:���7rƽ��\���e�.�z�����g3��>#}K�?A��R,n�uw/_)��Y�Yų�����^}��횜qlVe]��ܱ��cd]�O��B7;%�"e���+����7����Z�ٝ:d,j�gL&��pܳ#��4P�+ F{�������];$Nc��:[��m�C+��7)���΅�#�.��6�ZIl8�#x;͗�O�y3�V��U+���t>��h껛qYo/�a|۩����S-��%�"�7W���������O����n�U��K78L�t ?�O;Z�]�6�6o6���і��GW��'����и�L=ӎ+bA'coV�ӭ�d	��a-���e77�I�����k_
\5�,�0K��>s�۪��foc�*?c��GH
�����o�����g����Q71Ѳ�C��QWۤ��@�Zsۖ���(��Q!-�W�|��_f��[5h��'`���h�A��pLl7�DtdY4OG��UX:��d0��*��u�-��1���$���pN$�;��#sڝ�J���m^;bKQ_��˷3(v��w��u�;@������ӎ���|f�̘��3���u"u�QE�0L��8tQ�q��8��?R�$:�ƾ5[?���N߲l.����ut�a@��b�<S�q��nH�]�ｖw4�Oֹ�T�uR^�b'�5kYJw}6},�ek2f�̩��^�Z���l�۾}��g�3�����i�ۗ�4��գ/mQC|owH�RM�]�T�fؾ����Fx&H�6��e����w�w#oc�6I�t�R�.l���Z�y���2V0vҩ ���j����߮�������\Qٮ]�h,�>+��N9��*�O�M]���"�*==������s�i9$ڳ�K�E����C�,.�Lfo��"�����op�G�SM���G���ٌӻxsW���n�_z�"^�7�i���r{�l1���Sܚl�VwLM��=+�.S��|��w�o�*ڽ�~ߕ�Yߪ��R��o%���̻��@]��RSbR����WwwIsf�����
ƻ���kaS3��oE��o�w��|I��\�k� Q줭Kf<������Q�Z�j��1������>�6o�m����ʸ���|Z<A��i�m��nJD��㍐[�:�i���o�FǶ�e���z�t��n�s-yW{}������=���Y�ڬ�W��0F{��#j}
vFƚB��!uM�S�]�B�'kPp��Wl��e�Kg��Y��n
}ߎ��?��[��0Fr��u,�c��׼�&@��n�f86,��8�j�,�!��}�����>���6t��h��2�9{i|uj�]_�՗gqu���3��v4 ��Xp�h���]N���Y�����t���?�!�����������;��o����L� Ӱv�v�l�o�ǡ�c6���y<�Q�}�ދ��u�eim���0�Rh2�����ݱP�C�K��e-�F�%��K����>7J�tRH*B�������?#����6Qkp��c��f�U<,�ھX���җ/�h�H�s1A����;��ǩ��X��-ԍ9�R���ā6q�a��MB65(�w�]�N��$�Kڟޤ�#Ք����&Z��ME��^f��
�=����	�K�C;���CufU�
�o��wg���H����nv"p�b�VX��jǌ��':w�Sk���꣩Mq�^�/]�̐f�%�N���Ծ<�ә9kI�섟����=^w=)?�Gu��%M��t�
$�N<h F��V,:u����{�/��oGQ�C�PѶ`n��a�{���Ͻ4�i}K�$��9hY�]w���޳�����SˬL���}i�-��F�K�຾I��!̎��u�����fS6 W�
���o��2�ky�\c���ݔ��YD��]��e壽d3P�w)v[*����CgGoA.�:������W�L�<��}�ߪ����x�8(�����b�XAKN8�b�s�T��u�6�6�KU?n_�,n��n�Qӷ�1~�/'��,��#N����+fΗ7i�t�M���z�ٜ�T��J7b�{\��܇;{g{wI��Q�
빽^�r\b�'�+��u�k�!���leQ[�mt�֢ъ
��R=L	G���׺�뭟+��|��nĴbC2�9��÷zo�3�ah�n�R`�G{i"k�N��f��j�Y���M�um,+O���y`8�D��s��s8x#Nޘ��Mt79��7�g��5v��́v��0P��9"	����Px��ٻ=�dVͬ�&w�ֻP��i�7�Hx�O7۸3��$�4Î���X��(�_��K8vq����BAI�Ӊ�zE�K����
}3�aj|��k�5�򣙆�]YK0��pۻ5�
Ҥ�'Q��}�-�`�"�ZK�l�O��W��n��E�]5X��i�g�]�0��R���n�f��8�y3��twn�q�)	��έ����2h�Gw9�������ȸ���Do�����k���\���2ս�s;�o���"��37ޏ7�
&2�aj"�=䧧O3>�z�3D
T�$m�)g�i�V*jjƶd�JmQ�u�D�4�h/�	C��z�\xw8�nw�j�uw_(��Y��l5�N�h�}3�yY�Eӗq�2b�p�g6�d�r�Cv�F�Z �)�n')�<�V"�r3V��8��ʩ���m2�j�q��Y^���@g�+]{}�3.��s�s�Ғr��ƾ��T��PsFZ��i¨�'ѡ:�:b�kH�˭�7�v��S�����x��B��4d2m���ǘ��+2/����XH�B;�E�Rm<x��&{x������{|�c[e�Z���W�Y���]�C`;�"	��R� c�^(��e_ٷ2(�4�Z9���m��Po0���������9�{�.�T��e���J%�Ië7n�0޻oO.�7CWs�8堉��c��l�W��7��:��*}-�nZOy��d�p<��9�j�EVy�f{<l�9�^���o�u_v�����Q;�@G�ﱭ�=3�\�G�E�B�G���*��͐��@̛����3\"A\3��ei�*��/����Ƃh�9M�4Ɣ@f g�u�N�f~�����S�_|>N*�b���WNW�(�|dn�^ t91�Ő;��[[����:�~G�߆/��.f|H9>'`����1��p&0|�[6���mdg�m�:�O��){n��t�4���E��b���^}�us��lS4��7��k7��
�Zݚ�j;m�����gǩE�VR���S�2[ulU��#]�G�k��ȁß�`*��;�5�k^pz6��G���j*��r&^1SW]��Y�7ʦZl���D�8���P��ʮĪ���:՗��wK�P^��ҲTf�R�
A&��̛�u>��:�� r!���4%q��F���f��0RS�ܣ����[w��q����Q�uC7\[T_MY���λ�ZY�_u�����KR����g7������ꔱ�f1����:��OE�(�[�^	��lxǕ6Ғ���p�sێǛ6�o`����yG
X��,�j�<<f��y���4����؀8b�V�)4]r���m���^�F�Ŏ���m�|��v:B��d-hY�k���Kb���,Y�ctnkR����`��v�l���s
�v�*C����7�׺R��4�O�[����#g��+�,����w��ۻsY-"�N8�곙�mi����5��s�
w�6f}���3��gz�Ӷ�Ft��x�n����4'g�k��>�aɳܻ"	�E���'b!nr'�6��R)HW��Ob������Ba�.GM�l�̾��DVc��zO�տ�m�}[A)�6��; �����3��,��4���݋xG��l���]�_ePJ��������]�9w���7�f��N��o\m��K�����W�5H$,,^bm���"�z/�ǚD��^�l��t:#�,�����E��ɲ�z�n*����GvR;xpE�[�d�:���O��Q�q��g�U��z�V�BMVxLU_n�����5��R���8�����H������'�H��A U�؀(����?� ��@G�DETS���DUS��s� � ! �� b�*���`�(b���)�0b�*���b� `!*� A��"`�+*���b�*� A��`*���(`� A����`�b�`�
�� A��Bb�*���``*���`,�+ b�� b,
����`b�*�� A� b� A��
�� A��B*���*���`�A��b���g�`ǜ�@ �X0 �`�X0@�0V  2 �X1V  �BU�`�X1 ��`�X0@�0V �X1V  �X0@�@� 0V  �X0@�`�U�`�P �U�`�@ �X1VU�!`�X1P �X1VE�`�  2Q�`�U�`�X0@� 0@�`0�0 �`�X1@�0VU�0V1@�P��N1��H2@��2EP��P��EP�1������k@:@@��@@��D��T0� �1E2��"gc`+�C&@�1E� 0� � �T@��D2@ִ�� �F 0�0�H 1T��H�
Ɓ�62���"�b�  @b���n U��XU��X  1V��]`*���b��*���(���b�'0��8�ϯ�� �*�#  ������������A����Î!����?��z��?�S��>�����o㟼�?H �����~*"
/��DW�~c���8?$��_��և� @���ϴ��ä����؝��@�A;��~��0���FU �"��  $������������� �H�	�B
�@ ��"��`"����
" E� X � �`/ڐ\U��@��@� " E AX( b T��( E`�T �A�  DX  �AH D� ��� *����A��X*��*�(�"����"��}�	�����G؟� Q�$ �ADI�4�_����	����@���b����x7�O��k�?�i��Ї��i����V���>�N���" 
��_҇̃��!��AE��}���
 
�� ��?4���^A��y�l���@�H���>�����_�}
�#XwG'~�?O�������a��������DV����$W�|ξ�Hr&.����	��~x����}��w�D��� U�9	 ��}?Hl�����}8���Q~c�����(�?����}��}��(+$�k6�_���K0
 ��d��H�>w�IT��j�EU*R��J�Q!*�U��*)EJ��$TQ�d�J��T��!!2P���ET�R�D�j�RM�afj�T�e��K0��[fƠZ�,lڙ�ٴ����Rm��٢2ڶ���֬Qfa5m�*�l��l���զF���K%����cU����[KMeI��i�Y�&�E`M�jL�6e�4��bmV���ai��ژ��5jMf��4��a�٦��[lլ-�-��l��kh�  ���t�]����Ͷ��=�^������.��<����]�;Ƿ�^�*�]Ǔ^�kӦӬ+ѻ�'m�����l��q���uz�7�j��v�'��m7��P���֍���%d-��k,���  7q�(t4vȅ
$9��E�БD��ރ��B�
){��OWi������7r�Wc����km�s�i6�{�����0�w[m5��^�����m����cX�ǧ��6�M�Mm)Z�[m[M6i���   ��W�v��.:sOw��ڭ�mv�ʫ��J�Gc��nڕ�4��tԫ�ƶ�%u��wMn�T��v��eK�;�w)յv����w��m����mu)w�\	魌���m6ٚ����Z͛�   wO (>��� �ȵ�դ[M���ڽ��^��t�U��z�[�WJ��˵h<��J+:5گn��]��ׇ�{�Z�S��X�-�&M����)��   n���-+H�6Z���׵��GW�EE���N�,�ti���z�Tt�eZ�Π�tE"���=
��j��"٭0�l�66ͦ�E�j|   �<A������TE���P�3�{s�ԕW��uR��v�MHT�Z�����ܫ+e�V��n�y�\ ��Ww��{5�m6�&�]��1V�j��  W�@[��� �Ǔ:P � ��� �,���o6@�۶�{�� ��w��^�f� 
=<���dj�j�-2�Qf�Y�>  ;�JUA�����U@oS��C=� zt^�V�  ۰���B�]����A��]� �����{�����w��d,Ͷͨڕ���cZ5��   ;�} ��������L @{�gB�P=�i��J;��AѺu�
�秃���箃JS�Ƙ z\Ն��fZ;��ki�V��  ���V������:�g@ pf �dw�N�wyx )T�ާzU(Oz�7 =u��S����� �"�����)   E=�	)*P&�#*�z�  S�A)*P)�PJ� 0 �)IUQ� 3S������_`�sj�Oۺ;k��h���h+�t�es���4��ϯ���z�^��~�{���1���m����1�m�ߌc��1�cl�m����~��/����y�1-���B���MћAջ�R�'�k5����]"Ό�՜���:q�̊��]<��N=�S,�r`nȉ� � �SL��Z�+j����4Y[�dY�ܢ��1�5���V��wK�V�^���X�"mٶ�!�V��Ф7m�� l3M�X͛aa�J�:���t�h=t�t�悭��8����W���P�"�&�"����F�3m�3HXRgh'X�Y�m������3��6:�Q��DSw�/%Ӱ�����fY�߮ڣH�,6`1��7fn|�[Gmh��)@wf&o!T���[�-݉j�j�"4Dt*M�Q��$���ȊG�/"�xN�Ѹ[v�1�6��7��Y+9�S�����̎��m�F^�ݢ���|�bu�$��c���%��ZŪ�m����H0Dj�Ѣ�KU5��C�(2�����Q��)YhجU&�ah�P�ݗjn1��Բ��[ze�$*��dظULH�=�%�2�ε�ѧM����R�}[���j�*R�o����n��t^����ݤ�)+�dA��&���{�ˁ�e��2�kn���c�y��of���Gv��48���ٶ�E�yb��t������ ��,Ct2i[�
���T+,� ��Jm ��-�cv�Q��)�[d�d(2�S��^��'Hc�T��L ){��X)�0i���jL!f�.���ԧA=M 	¨nűِmMrX���Op�r���Il^QhU��I�Ena��v]��q� ��D�aV��2n�Wc9�-�N��E�]�H&�d�d��beYa���f]d�N�։j�9�C�iG"ub��� ���� �:FͰ�<hXO�er2R�WBK֖�J�Z��/)�R�c�o#��y��wYB��U�r�97C��R}a��v��m �-�ܧ�t��U�TŬ��ux4����״�T.����4���lt��Z���Sw0�)����JV(+5qIxZ�����IhT8�ٙ'K,ꕧ��
�Ǯ1�r�i�˽*�����R�1̲գv��z�JC�)�W�
�{�^Z�Y�i�g$��@Hf��M��,8\4������^�u�3�,�z��mשT�͡���)�l+Uyx�aE>�|�]�`��Y�Ô֭t�4�.+�{�M<uBK������ʆ^M5�7#��7���.H�l����H���Kq��Ө[`�&hOM5
���;Z����G1��ɍf�p=s�̭8��$���W,8³�1j�R�w)йN��X�ͺ�a�J�p'#�
�����{&��,m�Vkb�~�])�
�CY��ʍ���Q��J�x�m�����a��{�V
ʺ?8��M�*dՀ�b�`�fVv�{�%m�<bܨ�{��/�J%I'��l}�=&Щ��k��{D��*@��gBu�����M-��0уσ�n�wtw��e��meL)cd�Ӗ�{Y�[$U��6�e�T�P�.��7j�0�M�"ƛ5���ů�:�h� G7Pt.!��l��ygG؄�NNz0J�ٔ�<�
\�-Yh���Wi%��@͠�d����#
ϴ�X&�X���w"lC���ꖬX�U���ѧ�寙�s2<�y۶ʭ9si��-R����E(�.�I,�" �W**ͬQ�`պ�t��uɗ7tR�����WY���}�[CiaK���n����mw��޴��kʕ����	���V�0��͏"ZN��q�5{�)Gx���ż$f�*R%�&hZ�S��$� c�gh�l,ѡ����V��U�JJd���P�`���)�1�oQ�Õ�Q�jj!$f"n�)��fH�i嬪ؕ�Y� Y�j܂�e�TYR�Te7��l�j�CncK�9�A��;�� YrTZ�B��NV�E��@!z���on�4�!nIu����3�tT�����K���ƳD!ɫ,}3T���Z���^oj�/�ڱ�f�G�&�RNfV֟��/`U����C`;1�]J*���a��T��������mar��GhB�G�n�w����Uݲ���6�6"�{�
�����L� �-�7q��thY��Sn��yR�Z���m�FAv����@ (l(�w�*l��\r+8�Z
.�b;Tn%N�5��o3�̃p��Od�Z��`a�0:���z��8\������a���P*�f� ѣj�X��$ r;VE�;� ՛�U�*�b�Gtc�11n7#��T��
`���e�ǻyE����)ՒhV����h�aFʥ��"�Kr��sV��wZ�xW���O[�#����Z��ɹt��7[T�q`�Ѕb�x�嗹�gה�1+U���h"�E�XsB�M���.Q�q�p
֩�O���/1�B��G�A!��IRy{7& ��A�1c��{f� Vܙ>h�-��41:"l�<�-
ECTj�'��̶�)�K�?,��+חy[Pۻ���b	HS�댕)h.���%nSPՌ
��әgEY�CNQ��{CZ�B��x�m�x.����DG%�AeZd��ow)���Sq�����i� kZ��A�W��ݺ+K��H"��h�u�
z���Q�Vh�1�=������� m��b�
w��V�\��W1}6�f�(Q��8�

�;b�����B]�|����edn�E���F��{���b��U#fTo:F����^`��|ܵI�wX�7��q�C8L-��iV���72(A)��Ɲ�k-h�m��������_.�.6	v����u�O���]��p�1�-���f��xԉ����YH�CK#N�:ڷv�H����Xu�ԡo0Z�T���I7YqÔ��P�R�JHF���%� "i��YHA��'3t��	s ͎�&���y���I���Ix�ͣ���:ۭ{���lT�Q��6�k̛hC^f ��E�Ȁ�t0��(B��A0Y�X�JS,n>-l��1��4�A�N];�SE�0�E[Y�⿥'R�*@ܣ@+Ca66��UZ4��3����,kt��ʚk�T�buR����:qi���̻�]f����Ū˅�K�M�PY�jaF�U�Z��*l �*�;{e�r��m�oY�*��pֽ�eK���K9@*=�J�v�z�M��V���Iaa�� od�QK�H��7��s3kL/k	IcYv31P��WK
��6�H���6d-��7Cte(�2�f�`i��2�".��b�=.�����a�o�f�T<2�֮L#��M�wb�+, ��,X�h)NÔ�e�vuV(4h�]û ��D�0�6���eh`ͼ�ͅ��T@����i�
�oQZ�Pڦ,�[w��yg)�,���&���y�&㽺�e��%˘n�'2K"� �9�2� 7)^� ���*�Lj�gRu�E>��ٳ�iyםQ�ۨ��p�u����%�]-�Cfa�����a�/h�0]�8��楅�d]���e��1l��Y{�V�zv�[R)��D��*)]�ĕ[��O�1�*Z�4eۺP�D�PPW!���0IW6��v�wt�`'�2�݃me(\e̺�s]b�z�B��'� ���C�Z���5�u�M���fj�m!t�I�B��AA�(}����V*�3��]"yM��˿���[�-ٴV4��n�kh�6��)]��i)^IM',�˛B��V6E�D�z�	.��3�7/p���Q�a��5�7�+Q�An���ݣ��	 I(�k�
��f�V�ۘ�!ᥠ�Z� Kٕ�"��1(�#y2�j����Y���3kJ��[��]a�� ���{wWM�(�Q��HsA�i��L���h�A��+Ǌ�J  ֜�9� ��*V��!����*�Y�&ve�bBXl��o2�U!�8�A ���*ɏj��n5�W<�ί����C�YGf����0�*�.�m�^�R�X�F�M���;0���WOv�+G��H�����ر�P if��2�f�nk5���7XZb����َ���MYd�,��lt��6sG��F�4�2hr�?YV�e=���h=����૖���
'�SWm��:j�%�����%j�e�ɰɬ��b�iE;����F�`*l�l�&ň&�m�~�2[�`�$Ԯ
��5�klb�R�c�.M&=�`�w^աO뭐
���g7�q3�i��F!/,��L@+��]�B�)�V*e�#
P72-l5�fPm
[�t�e�"�(�f|�i��qK�g�E	2fV�x\d������&-٬^M�00�+J��I+�[����Lt�e���E�ǄV�AU���jZ�Sڴ�5�i��	P��F@6��U�%���PM�f�� ���A�g0��Y`�rb	,�T1*�z���1���MX��l�2V�+P:B�{�V�Н�� ]�Y������e�YE(X� ��lX�3�k�
�`��0���meo�"��e��=����h��Fw�X%#B��	Je�yV�%Ь��e�݊�f|��mn�6Pkv�k�I���pe6>�e����!�7����Ѐ�{Xl�+Y�h�ID6iX����+VFQۭ���Ҫc��T��ܬ��v�cIآ\�mͱ�*���b�ݸr�*��v�t
F&P"O� �u*�4���
]�5��w��is!S�M��t��M"�Xᕮ���sѕm��Mb��S6[ i��1c)�4��O�r�#Vb^�nTOf i�B�w��T�j��E岶�;�k)�6�;�ħVM�[�[�(m#f6M��	Gl�ti�,͑km�:�R�yt��5�投�a`��.M+��H��X%kWkp�Z�NV!Bʆ���1��n-��!U3Q.Ibm� 2��m���*���%�����P��nh��m�V(����w��̡c\˱�;պ�F�#�����7nv�Ȁ�y�Q#1���aj��<�I6�Z<�AP��m	�2:$y{���B�2�����Uzf#��޿�۳i�����7l<�M�f���fK����"�U�j=v��ܴ�4B;�H�*��v&۔�]8�:۠Ƞ�ǆ�!V��E�n�ph��tYP+M�NaW+Fƚ�7.74�{6ĭQ���J�rX��&Le(�ݎ[�,�8�����P�����f�Ml��aȃ]�X�i:�Rӑl���w+!i��ŋ ��S�Je
�lh���w�)�v��5-ܸ"C%ͫ[��-.�DI6�j�,��-�M[L�Б�X��D/.8�m�h��2wouaS�S�.�dOQ�U��V�_<#@�d�oT뀔*ŶE�C����v&��6ڥa5l�y[N��V���Wk��E�(bN���f�IaE�7V��,WQY#+-�f��+6����mQ�,�m`e�ۺ�&��a�SxU��݊Ǩ/��%��I����q��d���)�
�*�D���k��/f��Q)�Զu�G��M�#C�.�Va�.}j�ay�:-���r4BBi�*� 7J�OI�P����kO=�<.�՘�ҏex�R�hXOfmF�	n%�&�9QU���W�cہP'-M���de�ȰT�+#�2=�u6��YQf�	�cij�Z�`D��v[�-��l&���S-'��hpe�V�I��`�J�qn뱆��&�Ӓ�4��ܷ�A1�f�2�;&��Ս��H�h���Gp70�qj;NY�ɮ�mfjn:l^`��J�	����6M֚ےl�F��̸���{5�t��Ñ�,��Km�V�!o�Ԭ�y�[�*�ymZ>���aPNu��&�<�B�Rd��GQ�Hl5!�/��"�rbbف]]�Vf���̉�6��f4���1V 
k%�;�,��.f딄ܵQٻσ�s��N�J��1h�IN��e�i�]L84-�wT34,���������)�eH�r����[��&�m���wfk��̵r�Tĭ9>�3r�*�OwK917o6m]��!Q�[�[�����8s�Q�$�'Bn�0e�3)2�Q��fK�ͬi\ө�"V�Mә[)`Zر��2�+�V4���f�ͼ�������P�nA`�n,r��Q	4C��h�,�)C�]�,9����x�f�Ж�	Kwc幣i����ĝ����$�ӊhu�c�+n���kl��,�ȭ�#S�U��]D��v�M���!�֙���-�,Z��ԣ����.��㎶+��4�fԣ%� n)��4yM1Z0-7����W>+5?�#"�W�Ct4	���ܵn���t5]��6��2�Q�[N��ɱ�l�ˆ����A8�jZd�f<5�2�Ʌ֚��&�		Hmc1�W��m`9A��P87m3��J� L�c(栌1aI��wa���K�t����J̨���,x��ZZW#܅6��*��B��V"��anf����/K��e%�K^]�;�S�Cl�Jl²����Xm9,VV�o(��ɷ.�h-$Ȱ�2W6�K��@
dj�wXF���S%�/��� إt����X���N��!�^9�hl%Ħme� �NQL�=�7.����SZKZl5g'ی�BQ�gs�Z�fAX#w�^��5n����ta�2��8��������Ps"�ZVj.�ҟ"��E�'-��&�{bJل۹[����'M�,3)�����,��yvP1&�)�ĸ�`�-J��"�%��؇2|4����L�mJwJ�4�,q�B���Y�l�1���Zԩ���1!r{��҉,'x�=d��GB�!����wnE�;egMh[�w�6=��guc����i��S�;�h���]X��mqI-
�w���2�^s�n�d��qZL����o�S��m�6N�ɦ�vLjN�ιJG�b����z��[+o�6�5)v����Ma�2���u����Ψ,$�ܥg^���pGV)��\6�Iqs�KGhYY����Z�1������C�XPt�<�3s���+�u�l�����x��Ϟ�����ii{H�ȣ�>� ����� ��0��thLz�3�YG�䳼�TN����n�It��
U�S��vլκ�)�z�
����M��T�,ǰQ��]�ے0�Ya��YB��2�᪯j�V��4��d#@�.˩�/6�sv��m���X2�MaV�]�sؤX�0��ҞT!<��(i-c|�: �S��n��'m�kz&�e�o��;�פ�[�=��3�r5��ҵəen��u�t���`�ӫ�����e��z��^�}W���"��=*�\�u�I�ﳠ��5��Sq0؄���Y�Ԉ����E�v[��c�wJ�zl�J%�Q��;��f�K�=�"#��D��)c��s<���:4��îi��|k/��b�q�X���Y����}r����3�#��8���4�*��̻�e8��;7�[�ߡ�靓��&�V�	�Ӫ��������x����N�4�p�����Q���<(��X�*�e�FSR���>�,L�o���w\٬5-K�b��v���PЮ��ү
��Oa����S�5�;�a{5�V�uiR���8��P���T��[~&��P���Ǟ��̥Ne��W:i�ܹ���,�L���遘\2���WG����,�k��_]�'c�[ܷ�@v�6N��b�sۮVgZ6'.���� �0���ͽ⫡7F���,�e������Ni��v��ED�;�|i� mѢܾYYqU�M��������j�ȶ�^�CPK��ĚwY-�:��g5��h�WH.�{��o�ʂ��l��n�ӳ��x,#����[|�ù]�7pU�v����#�#
3� W�[��D��u9�v�@��8^�[���/O<��[+1��i�N�aC�M��I��Q�h�07�^:�mh���ob���b���qV0�f3�IP��$I�3�c��v�[�t�u[Ts_5�s� S���v��|�L�[��`Wʲ�h��Y�M��nv	m��*3&
�j�*Ě�=��r���*u`���24YӴE#�Xx���\�J�U�}������n�e딜o�����
����4��N�3Jit.\�*s�̔V(�2�ؚ�:��q�.i�!	Z]�඘�c�$t�����j�Vfu�Wc�OTM�7)Rt�dGV��V�Jk�6vz�m��P��@T/�ՙs� ��,	�l���-3[��ձ܍�sy,�O����faf��)b���;���J(>�sgT���N��-w)vQ�ǇtihҊ��j�Qw�yۂgS�1)�,G(n"Fmч7�D<���6��Uܵ8W)۶�A��|ʶi�.�u��VZ�W�!��E�{{�|;��Ո��Z�logh�oV���K��`G���T9�q]��%&�c�y<����ܥ%LƂ��K!�w���K���:�K�:�i�Y��	B��t��m^}���fmu@D���BW`��A���ֹ����r�BF��z�鵜�Bo .��o�OX�X|r*�����;9�����tu܊҆�Pn�8�EL�w^��Y��pX�9@_܆wzN�غv�+�����ʝ�z�|/qA��h�r�|�A��U1Rb5��zc�������srѵO��MZ왆ĝ�[�w��,v�Tl]���ښoL��+2��sr��jvT��K�+I�����ٜ�i��vj�{;#I,�y�q��/*.�\-�9�8T��Dwq˱�Q��-�)t鬵%��p˔f
y\'9�t��I�I�� Q�\i7G�\т��'%ܟ���5\���)^P��<r�i�]��oA�HE����6��]�\��}�V�oS]F���\��{0�y��xJW�Vxzj3f�i��%�^WV3V����`>�hT0V�Bi�Bvl�{
\ B��Ol��*a�"��Ie��.:�SJo�3n�w:��B�e��qٻ����K4�#O;f*_v@�y-��mr\y��L��t�Ȫ9x�X�������j��m���I=h!Bί���˽�{G7f� �;��,�
�JP\+i�D���C*�]u��#�������k�	�E
��v��8��4������-��:��Va���F��ҕ�{']LyY��z�dg��{M�k��}�)����//M;vsJ��;hD%���JE[j���.�M���횕m�������*jݯ�f�A[C;$a�������Ҟ�Vn�7��~I.N�R;B�Kji�G$���%���d5��J��Ȗ*t��p�\��2. �S��s,[���F&/��3����=I�fg
�o*yB����b̫W��;�<^�D3Y����BT�Q������0�2�U����('(@Jv��]1�ӛ�%!;�I�	�6�5��P:jZ�KOZl��WMo7[����E�	,��x2����4gSV�g�E)��@�֝�v� ��,;��*�ET��S&��0�R�L��ņQ��������D�B8����u��R2�֙͛	���p�쨲W�&��^ϑ��/���w;�	\ �����y�(�e�=v���x�3��\y�8x[`f+��+��U��"�$����ݩ�Y������(:U��A�J�)���J��/w';���X����d��+�f�0,6j�<�GD�F;A\� w�]�a\��3�
�m��h�lf�=SyJâ�]�s��vV�R���6�(�w{Q�M ��G�m��Kuݸ]��au�j�n[캙3/�ͷ	o�WzK�J��LB7ל���#����f[t�#ĝ����\V�3i���y�0��U�����~f�r[E�l�L�Ā��B&o�wV�E��K,�1�P��ز%�s����+ci��"̀�K7u�:�;�2鉜)�m
���z��9aE:'�1i�f[�5�Q���X]n�u�Ȱ��σy�8 |���p��V�=�2vEi��L�p����!��e��jϱ�5��:ڹJ?W6\�+N���΋oaC���W�'�(�Y���u{�@k�툪x���Es�3	J�ag�m��2#e��$@9�;��CZ5hY�3[���s�z��U<5Ħ���[%i�4j�2hu�>Q�VѺ�昺��pw
�V^*²G�r����N�Wa��ˤ5�e�\A]3t�lv��<ov����/�)��J8��g����"��5)��.�g������N����$���;�u`�7���2%$�^���4R��vF�y�j�8�����������������u���)��`��`���z��CΎV�h���ʙe%����RZ�7 �vc���r�s4+I�A���+��c��{KnF�c�Λ���b�1�QUҠ��b]|;��9�y��֮;D����(�TuB/"Wc	V����+/�(7�[A��.@*��T|U�ú��`/cQ�����\	���-�O-)v��V<�u�f�p岐�>S��NS!Faĕ�'�;ؔ��|�X�Օ;�3m0��TG�����7�[���4�)���m���J���k���n�o
Y�FE���u9��NG^�aJ�j��U�j�M�ٹv]ζU���u�+f��MX�fw,sR'*�9�
���)#x��f�j#q�|� �좭��#���$�e��9F�4ga��n<C�)Ze
�q���Nk�`���衍��{�,w���r�����\Y-U�Mͤ�JL���|����o	;��t��ۻy���O\J��7��;��r�ĭc"�]�'�����m�=�ﻍ $1�q��$z@����ڒ�-%��]��I�-k7F�U��-Ѱom���2�%��Z�]^��=f��V�iX)hUo��E�w{�O=:�a9�x���Nb��;��Y���˷�����.�æ�<	ڒ����i�IG|��]���Y��!�B���/�>˙�.\��2�A�Lz���M}����ٲˀK��V�ޛS�Rk0��[˖�N��n��&%�d�a0�8��oP�g;�Z����	����4�b=�(�lU��Ε�R^mr�5m�'Q��[�h�㨫_,���fqV/i��]O�2�u���[qZC}���1j2���{\ջ�����\�� WK�^�+��my]e:ٝ϶J�^�lp�Wt9I����h��I��w
뾱�0l�{(�H�n9�ٹY��,Ĺ򳗽%=S@da�_78��o[Z�LfN- r�d*3f�9Y���ؕ������%nD�l��C�5��4����FI.U��V�V�Vd�v��K��g����X���(�"���yc�+������*�R��p�ඵ����m��۩�]�z��X��!�LJ�ē"�
�u���HӾT��%���ƻ�m��Q�q�^f�96��"�W�*��꾓fS�=C����2�p���_�y��^w�=��e<��x�f=�c]r�գkm�0԰�]��G��31�*�1�`��uƶ��ies%��T���q����U�2��f�2���Ya<*v-J.f�E�q4�>�M�$�����x�w%�T� 3.շ��%��-���T{���*b��
�k/w�'l,�%vGS�r���P�	J�R��k��R��a�������x&N�\����2�KO#�%{�C�i���]G���d��{3! nkS%9{��T�����"3�{.�[qU�[]"�F��������	�n��zb�V/o�_*���K����7R�n�]|l�����@��8f&��z�:	�Y���(Pm*v�ƕ]�\'��p���[Yay�5�����Il�R๱���'tx��Denݚ.g,Y[Z]5�7:�;z����X�ɐ9����=��J@����]<�rv���(��TK�.l^�l�Ve�!��Kb�d*F:\�}J�ݫr+KAPk�S�it��1񵑩�&غWRTO{��bU*�\�����tƈu��a#	�]�� �m��ȫ,�4D�u�J�8&��'�r��U�ٜsj"S�5�h���e����Yۺ��M���
��]�\�0"��CA��V�	��e���<W�`
��u�z�/uJ��E���2�
%��FN6X��HenH�X���mTR���	Ucc�H�Y��Gx_�E$��Q��)���y.D38�f���Q8j�$��W��B����ƻ�,��]r�m_G&�U#T�,�x��O��e��1���X��g!9���Sxր����!��	(��w�lv�ZG{^*@�S���u\rGx12�E�H�@�n�Y��Q��2��\�t@Z�c#kG�`2��̗4i�:�(u9�����Q S�y�vjT���(+|gvc�mv�������	�d�\��꛵�.�+�`\�=��8�뾴��0(�9oX�%����m�΍g��%�����Nٰ�B���j��]�Ã�7��k�1��nv��V���U��q�<��9/D�-����/m�OsO_c��c�v��h�B�9@;F�Ფ9�<����O���:ne7��>����itȟ`����@A�u���m�$��t�����E���Q�Щ>v�[�ӷ0[�׹�n��T�6�\�	���Ik�w��r:�%f*I\n�PM��4�m�O7X��`ӱ����S���UE�������B�Ct����i'{{��<
h�ѧR�+o(��ބQ}Y�l\�g �Ņ�8�Z��3p8*�(���I❫aV�$io����c2iƪ��e��HW��i�`��D��q�w����I�V�����+76t� ���,�r�+�Ɉ������9�W!tO��;a�Pw�[��f֚��`��� XQF�p@Y����w!/n�:��R���MQ��1Vo�
U�KT{�)��7È>ɋtLy���ޛ�wR��F�]�.(��{}��xn5+|Fnr�2c��.���iV^6@����g�婻e��6����[���9�⑫K�1���2^6����eP�w�Ydڐ�=�0:g:˭�)��`������.�^���Ra��9���^�1��8���s��X��(';3F\�6ҳ[;71�:N�a]1`Y|^I��riѠ�j��ەٷ ��k��VǏbP�^�ն��o� ;�u_U�D���
����86�jLq虋s�u&rA-�;���#1U�u��pZ3��
¹�3�D��5�RuwKC����ܻv|1�[[L�K"��VȤ�'����~�i���k�&��{��b ����Y���t�(TS�
 <�f��&�����Js�r�qY=��;F�Es�7�I���Wk�4�]V$��ۊ��.��ѕs�ʈ�Ef��.۹Qk��YD�9w�&���O=�.�����-������ME�rs�Y6QIp���SWD����.NG����/;�,P����ZB��%ݲ`N�z{ICB#�	X�Xj$}������[\��M�ޗ4����N��4P:�;�U��Ó9�|�!�*��Xd;�yO7m9w)v�:��2F�)1�c�dNL�jwl������kFAf��	�c���D�ﹹ(�q`��ƴ^����J��N���ͫPue��y7�'W����ׯ^~{?}��������m���c�}����.���-�MrlKb��jE�v3�0�W!��,*�5|&H���[���+�[x	�hfGJZ{)R�K{R<P$
*���w(2gq�������kR�@�к�m��X^�g�n�Ns�u���4�޽�\�0�����&f�.A�2��A-t���rn��'24�u� pXg�ij�b�{��<[2���d��x�vma�4��λ<�i����
�HZ����Û�E%Uڎ��Q"��12�]2����{I˼� _C|U�Y�#�fsv�;GkOb���V7It�~r�秖��ٜ��A2n-Z9qs�7�j�0Z�3:\�j
�i

_BU0�w9���e!���D�����-V��7/7(0 6.�bÖ�|w
��{��N�|L�FzsM͹�l�1Y���1��nX1��M�9MR�}�N�w�@hz�ާ�v�ˣHʴiS���4�Bo"�骯9�:T>�780�^&F]�`��(�6S��ی�|$�f�.���,��4˜�B]�bT�=��u�����b�Wc5b7ܲ�`�fj�����n�n���%����̻ P�{;�\�\���(v������k�^e�k��V	B�ֻ1� Y-���b%u!gz�FL�`*�c��Ĩ�7jJ�L�3
�c��\ݩ�X��f������y:�<.Yڿ�cobl��f�L��Ö��Kz��ݶ6N�;WT���ɸr�7j�w�1���1ܺ�t��OVpSB6`K��@���y��ٴF���w%�Fo��J�KI�@w��y�<�段r�uz�3ZF^<�����Z�n`�8�W8�]J��J���LW&/%C�w����``S���5s�4\�Y�p	�f"����(��e[Yܲ
�.��\{f�}z������!���D��}����(�i;Z!��t��m�n�:���㵝9c�*
��#��6̾���K�K;�,N����7�o�j�C�g�x���Jk�r��gM�C�J	F^M�Ù�ȏ,n�^L�=�'�g]<�G�@5�]%��9a���F#���4��&`�X�:���Cg+pѴ,ZZ`�V/�`{��i�c�WsܗnB�v���[y��v��k�I�М�][z�V���e,|�52��Љ��+OV���`¡,���*�fE3��Z�9��rP��N��{a7�]KnK��-��؈k������-4r���B!k8b&�ݜ3��/�4��Y�����l9���YKn��}Y+(RJ,v3)���A�񹛈;D�C)�{b�*��-VHd!ωXY�q�����:�gA*i�Ԫ�S��pv��,;eeuE4r!�7�����[��kI����t�2&5��;X��5����;�=�&X��B�R���h���[�q���P���^^�8���r�W^����QD���*ћB�-�St�?n�z2�'v�&��z��="<(fIq����'mWt͗v�EbE�=���ŧ��j�x�H�LY��]�6����Rf�C�EtTMZI8���8]�,�r���=a�1�Nf�"
wW`�P�`��]
��0*[�7-���b��Uj7{S1<H>V�to:�8"u�w	x�m۽��+,z�܃k�V6r��,J��v7�;>�����6������e�rm>EԻQ�7(J��p�Lb�LHIZ����8nee݂(�Ն�x�s�VU#V��.
�WB�'K3����]�|in�Fes�R�J�̶�э4t{��0��-/���Z)_Nz�{�#F�k��Ń�y�"����X���>�!�m�����a^�j��G�U-�	XRb����L
����Z�b�9�N�Dww��.�˕P�*�;��MeWNW�.炊x�̗ج���Yu��<��(��+rm�k�7��J̜�*��=��V�y^9m3�i�v-h��X��^1�u���'��zO]=��B1��I��z[�e�F��|�(���k�^ wX�v�G��P�(�WO/����E (�tV���b�n�^����Ɇ���+��JMaz�fe&*�¬=�m�[wX�K2!MV98,��]�˺�;��P��*���V;�)rKD�o���뜳:�Y1.�DN�T��Vh*�Y�Y��PTN�f<_\y�)��(+��٭]}ʅ����s��T⭏7u����zdٺ!�u[X3GA����==[���ha�e�a�{��p��(u�H��l;%;$�x#���RrB�+�]��d>�pSArJ�Y.��W)Le�mZ}���ڷ����o���2�5�Z�)�NhƄ�&沧p�6�Fc�qv+��u��R��+�Ʊ��Q�̐���Ji荔2��aL�|�L�̛\2�K�2����O�I{�������YL��L��.��֎�:��h���l�T��,�TeYm�{���7�lk�ս�v�*
u���R��LrK����`�۴
	�Ёk4eڷ��8⦎�.E�lUۊ�GwG�\xiX�pu��w��l�V6a���_"����q��1k{�T�gg<�l��T�he��}B�4oa��Q5>��H619V�f|m����;M��oE��;8O�]��.V�C6������R�����]�ة��)@�2N�N�˹
ܗ�������hU�a�}�u���K��m��/-��m��Q�|/+��_w���G,<j�̜ �) ��)e�-ս�Y��h���Z�s�#�i�m6[e���nԥ��Y{��r1չ�0�"sS��X�TӼ026���n�����e��	�:��c��ܾJ��ݗ���ɰ0����R8�H��Jt?pU��6�)�b��m�.
��Mv�;�_e ��܎�c�}ܕ�4�<f����KF��^Z���\����E7���wV:杔��G�-a2Y儬œ9�7�f�c~�f�k���Ո<����5g!�����\�5�OD��;X�`G�����tf�3w-�yM�ٙ}��j���ݱ��WAy��[���Bto��}�2uC�mQ�5����=��R�[kfR��ZS,$T��U�Xy]'ol�b��ތ��X�q l�+5�����P���F-h.�G6�]�9zy��er0�]�HY��U�l�u�I�G5��I�9����p�˲�
�2��²]'/Z}]1�c@�kY6`KogeԮL��"�%�kr��	j��=8��W\4R,��ʸVH&�[yĔ~�ts��B�B�M�!d@zGOv���"Jy�jKmV�����B0pV�2�e�|E;>��v s�	��5gKb���5�TNq�R��#Oj�Ù0�5d�������b\�~��\�e����/JUEu���+���e
Վj�����c++hN��h���Ve�6h�Ż5Q	#-�[�d��aŷ\��,<�Hgm�'ג����t�mn �`�y�54I�Tot��Tg��E2EO;�s��k��������Y�B��(Vָ���A��w�� ��J�d�t�t�lQzsn��76A�8��oX�絣J�/r麊POUٌ�.4.�{R�dhܹ6j�g�hd@�]z;'5�$+�֛;]|k�`���6�ͤyJ]}g"�-�ٵ[2���X�&mu5��Oi`{��(ovT����{Y7*��i`�}�j�Ss@���"GCM33EY�u�6��g42r�ň�a{ٵsm���N���V�u2�U�oEٱ�v�$�X]�M�}�B'�,��i`���y�����惽�(G��Q�ގu�h��۴B��|�ee�H�t���Q�#[��J�An�w?&Fl9�I��]Gs���ٔi�>��/���0��Qˣ��@K����t���U���Jޥ�`�ُk�vҒ2��/�%tV(�t�M����zT�'\NWt��5�|H=v��H�;�c�oo"%>+r�%Ʌ�+G�xҘZ4��v��8�b�ڝ�������Wp̛��R�f��oK�A!�ձ�7#�ه94"J��u;eoU������n���P��7uz��.�0ѕ�8�wWu�v��ٹ.�"�rw2ɨ��v=��%AN�윳7~6����6S�$�'�y9j];7�¹�$T�W+r�M��U�%��ܘ[g(J#�̏u����iΦ�����%u��b�n�fZۮe%�a�\�`��T�8T.;o��[�L8	h�_���G�V"v��77ELY��*2^#w:��\�w��vZm���hP�"����}��s�Vf�I���-�S�@���4�_9���+��R7!)���er��kZr���Pd1�vhU����0k4�P��\{���QܹE����X
��R�=;[�ͻ4�:7�(�IrJI�m��q&�h)�NU;��ֽ���{�[W��"/k5�� eVue�T����f<\Ȭy��R��E����aզe�_!:�7]�9B���6�ur�5�L1srFz^�m��7c�����w��ѯE��Joa�M�[�<^Q-���u�_B�eMk/�Y�4ѽv��p�w&8���R@*����Uq������V�s��:�l��[�A�(67\Tm	��sz�=Y�z����WK;w���NyFLU��<�u-��Z-�6�J��|u�yt+��,I��vk+6敚���2��Չ)b���+��C/z�Iq8 ����\r��u�u�V%cF�ի�i�����c������3�Y����Kvq��c��c"�Y%��n�E8<�0�	�z����a��dqn�T�u�,)��>nM���Aor�nsx�{��-:�"�c%L�\�ᆶȴ�B��d�t��S��m�Y5j�[jH*7�{@�Acp���T�:��l���Ճ+B8k|i�G�	v�����R�{����e,N�OeB��L^�2��GU:c�ܲ�)\W-a��4�RZQ�T�F�,G�a��n�N�r��
�R�����@&u[h�3�q���ц�ĸ��̩��Ͷ�\)Lu����:{�6X
�@řs��5"kI�c�:4��Fn���wHTF��ng�z��4��,p� 2��Ud�ޣ��(KZ�F�i����R�4u@8����M"]�rm؊��*�ۢm��Ak`��-i�ou�K@9{Y�
V�f���'��C�Y���Қ9.Ƕ0v�w<��we\��U��Q���4j��[reYC)�b���k���e){@��V �#9K����tnquq��t���9��'b�͕:��˼��N��M󾁇Ѥ�V��*m�z5҆�3�c�����KL����f)����p��hµ��;�n���B򔛉��ep6R����V�0J�R�_3ַr����aލ;�"�լ-]�u7���Ip]_�%<�e-�pI����w��Eie�CI�+O\���Rg.��ø�={xjd�A�m�&@e 
���&a��c��ʹ�J3Z�!��ݪK���R� ����yt�� ��؀{�A�7QX{�5���/]Kz�C��U�Ba��f��6��$��ڢ�鷸�����Yj���&�*o�(�P�d^f��n�J���Ð�t�\�����̀^�X�.oCU/OSB��ȯn�.�psKU�su����^Θ�t�d��:��G�$�%{[3��h�m��4%�ѕc��k�k.�M�5ƻ��+T�הL�[���R��*��3��n�R���m^	�'Y��i)B����Ƀ \�a�qQ^�Fާ�����'/[����)����Q%������	x�~�D�h�#
WD��Ǚ;)Iڔ���������N�0��d���ki�d�z����R��Q�@#�C�J�2Yt�rf<xmHU��K�x8�G�=����>!���e�#��x���N��R�c���Q�
�n�(�g8a�n�V�䶬Ezch���6�&��X�t�V�`%VfIźŻ�.q}gmV�F�.�`vֈȝ�����2��v1^o3]�p)ҵ���z�"���f3���T4��v�\否h9�����O�zn���K&�y��͑��)���� {j�4IO5���+���4�	A��L��WAe#������+��T���E�Oa����j����8�Et*,WGձw�*.��AQ����]����>��YY=U`u�x�#s����t�5z��VWX����[δڲ܃2@����;��C�`���>S����Ef��V*ŋ�E;�������7��m�{��^ud���yz�B�|�1g���}&H]j�����~�ݵx]��k��0�.�&pP�M��
i¬]�&֨S��������kOd�-��ha��Q(����]�ub&]Bv�@}t�`hԱ��	B�떝r��m��n����L�g�h\ʶ���&ܮ/.H#�p��k���֗,o&��\�]���Wol��	�����ҶZ �*٫�x��� �[	���}i�7Zw���$}���R�.Z3.�Ċ��G0��½��8��������-}z��Jq	r��R�sǍ���3v��p�wr�׵E�@��fӏ#��9^���Ƴ���_;n�+�rP�� �h1�i�J�����o�+S��ұ:�H�b��V������ۛd�5Ƹ�}���.� �gWU8r��6+-㥙�V��bmhGr��+�K�&��h�f�C}�w%����F�n��b�J7��K����o�r-ޡ���#�pcqF4�V�jͫ�q�]h�D�'�%�R�kk^¤U�f���e,]�Sn�9�}�g9��A�V9�C�rL��Z�W-��@I���GG�Ra��:F	�^-���ؕmu1z�p��E���A �{|_E�s�q�PX��B� ��ǐ�ӭ�"�V�����{�@v1L���+�?W��}_W�|���S��{WLǄ�,"qz�[o@�<��L�oy����wo�TEʇ]*���j��V�R�y5�G+|z"�]��^���"�4T3:.�i먊���w���Ԙ@�X�컋�vu+ıY�]I3z�U���D��B���ʹ�2���:�U�|���9����OS�Ғ�Ε�s�ld�8tꧫ

�+l��Y���8��{�
Rҿ.7��q#���v�Z�q�CV+Fl91��w�u^�B)z��E�v`I��Q���w5�Մ�	�2�4���΅Z��5���1�,�t|����p՗�6^܄V�;O�u��r:U�)L�lu�d�:�Wwjn#���E�q(#z(�.r{����,{�ީy�(��#{�\�j2�Tǖ+j
�;{ٹ��	�\�J�_^�auVK`R�Y6Sew64��Y��D5@fъ���*�7p��_��IAR�.�Q���ՙ�6k�si���5:&��N��F�X6�U�p-��=�,��4���T�wƉ�/�J��E�{=��О-,l�+,vEƻY�v��x���ҏiҹ���'4���-P�R�ج ��˕�2����6"F�+fQ�"��qܫ����������y-��56ܵ�9�S�{%s��D>��z+(7�^7)�}4���q6a�=[)n�uc��Յ-��9u:���#��zZ��!F�#s�ZŽ�0P?h�P ���K�E�r(��܏��C�U�Yz���5us;����r���PDE���,ʢ���C���FVBVa+H��Q�DRd��D�(��Ay��{�p�Ν!P�HE����3(p��%Zy��$��h�<��<�!C�e�R*4Ъ#��s��V�Fy�C4VI��/8 ^��%uR9�%�)�(�z�%qw�"B���9�,��s��R֕*���(���y�Uw�(nQ���U��r�Dt�nzqq
u�!8��2׏"�<�@�$�G�"�˘��t��0�d�wOR
N%��R�̅K'=tr���O$,��r�掮��^�UC��ʍP�"4��B���fqK*���h\�
�E^�5��߭�r��qۣL���v��Ne�ܮ�rP��N��T�ݫj�|F͞rñ]:�J;g"i�N�5��I_#�,y�9۪���v��FaT��;���R�ιS7Y�� ���:���Ͱ�{3��v��&2Uyh.�@k��6�������႘�X�����t�S
W��p��eޞ��0<��^�����Q����X�_i��*�9�ł�3ؽ�+�룇:��Vc���I,�����񋄜VX�^���WyT
U��ճ^����6f�wbl��9e^�PW_N��_+���Ɲy'43}���b�{�"��	�2��Cǧ������y��P���s^7p!C��;�z:Ӹ�!�:��o��Z.u�7v��O�-�⮧K�d����Ώ��Ꞡ=���+*��V�=��ʩ��\L��UM5]j7�t�k����ݧ�ͺ�w��>�3ThO�quE/��װ��0d��7��]�t����5��7��y;�lŵ�W�������4>���?l��������1tL��X�=ӣu�<d2U����xC�'�_�Ͳ��pm�pCV����Kw��ʐ��+�ၚ\}g��{���w&�>��|��`�p����gD�� �ٲ1���)䋩��;�\�_W�j�3W,ڒ�i�M#������Z�$e-\Y�]u`����r���8M����ʝ�C-�h�\R�!���8���ς�	�`����u�mR&��y��:գ�����>�l�TZsB�}E��AV9��1V~ƽp�����ا � L�{5�X��:��·����j��K�4 7�>�*�Z�k���R�E��ײ�w���/�A�`�c�+r�j�QgY�]��-��)�j9�g��ۻ�n��z�ϩ*B�P�����2��91}�ʉ���P���zw��<-��1J��m�Q�E�<�v�*m��@"0#kᶼ��8���V+�]w�<��Y�?<ͨ!��2v!�@k�u_@/��-WTb�����c��9�v߷��79������uB��ɨn\���j� �¦/���~md�_5V�D6���u���W?X����0p���uy�`S�yW��ޔê�]��^��%!�V�2)�� �{>�I��MVa�_ײ�?����W×�+���WU�LV��ߘ�Yln��;[��-��˸��r�s!U�]/�j�t����AV�M���^zr��^\ǈ��$7�vƂ�uq�OD�W%Ffv2�P�Ƙf�^ɻ�nԅnt��3e�!7�M�x�4��w�R���P��f��\�ŠbH��Ғ�@����T��3�1>)��,ʏN��@2r�/q����	`�1�c܎�D��1Y�'<��]�-�k�<@S��'E�K����[�U{���d���.�HÅd���軆g1ޭ�����{-;�)�I�@i��'�(���W�/nx�]_�Dy�ut}"����P+��m�L�;���f+D5: p5[0X�)�F���	s��k	+ΠW���#���'��zhE,t��~u�C�{�{o���ά�Z*����+K'3���T<F;�9hi��Zftk�//`�j�������,�cA��%{�����w���rY���=�C��EU�UGu�8�o�}�V߲S�ε�Q�\7&�ig���Ge-�ғ\�j(u�ǂ{͟)� �T>�N����*���~�!�ҍ9v�R�n��EcU�Wd��wFM�M���1.�	��l��)�݆}�]��=��>J4�v�(�Жk�4c<'��E�!���%x:��f�s0F�̐��U��ӱ��q&ۃ�5���j�a	�Ǭif���͑�0��R]G�͝N�]>����o��ZsM���	˷N��JxR�0Cr��[(�_ʬ�t���l�� �~˦(R�V��X��w9j���1�Ꙫ���e&M�e������ŶV[�wKxL�3��_]>5m����d�ۜ���(�O��3U������l�}-$v�c:��+���{���!�6<:�o������/R��@L�3M� ;�g�wV��P�e,x+m8k�z/ #���*ݕAe��Թ]�L�f.d.�|��!�߱�j�������&����
u���i�1�+^���X��s'��v*�WC4?*�pҼ#ȯd�ʦ+|�}��eD�Z�9g��ˋu�>�,ZL&̮�Ǭ�R��[F#ۊ�\J��@!�G���Ǽ)!N�, :ʫ�}ޠ��s}�C��i�[�Ӂפ'#
zp}�]k1j��p��)����zb��7R7�v�X��m�S&���Ώ<LS�jv�}1\Q���X�S����צE��M���.�#�X�kRW����X�ۤ^���1���68u��zxy�c�%���Fa����42qfw:ǯ�J��u�Aģ@�b>a��d�ewM/�bs_:���0+uySkEޝ��1�߆cg$�k(�����CK���a��HT��t	G��a#Qd&s�3{���zf�2�� 5�ud���Ɓ��)��a�k���;���E-[��
dyճ�m��h5`ਟfP��ke�3�h�T(]��+e�W�kk�z��Y�Ȁ(ˢ�����\��ra�&;��TIҼ�.�ζ�\X%'��&k�R�֡c+����3�d���i�,�+�7:Ӵ�Z��{���+��b��y�n����aI��un�Q4hC���N���c�엇��`��n�廻f�S%�P@�W��� dH_��4e��%�)�h])�����*������e�"�9	��*Ӹ��s}j=F�:=���ƌ����x�hf�A�h�?knm��g�m֒�̰5��/me{�}�ADu�����3�({L;n�.׌��Y�-��ϛ�=jwi�^z��P�W/�1����C�Y8�sC.�0'涼U������Ǵ��z���p��ޝ��"���]lsu;.��`�����{G&lC�QC"��K�r�g�����sc��k}��/N���<1qN+��j�����i9�	񿰰)m
���-�
�z���J����5.�i螦���T������?���^K���W.���b_6��p��dYnـCĭ���.�=�ˇP�M8*S��"��oU� �N�/��y���٦�����{3�D��k�{�o��!=��
��k��멩RнkX4��O<�>w�u��+���ێ5�Y�+7$��J��bٳ�;Ocy��̏v��r\-����t�]����qT�!���;�����%]G�֑�)|#�yfk�:��?y��@��g����?	�(��=,���[��9�p=ݽ�KȖ�LY.��uڶ��������r���,F���v��ɟQ,�g�K���Y^�<�ީ������z��;^�n�3T���z1)�1#'	��T��˗O),/}�����s�¸ ��ϡ�,�1��{P����~�1�"��Ǐ��m����)�T����R�������f*��8�<.�i�#��Z����
����P\�J�0ݧ&$m��G�@M3:� ul��LF��

���[:=�7[���n�A����'s�o�3[�y���Խ�l  5�$R�$��"�ʍˀ����<�+Y��D�,^�z���+5�uqtE��U��;�>J�ᢀ� �g{f���n�޷Q;�뇅��f����'^�]��vj�w����|8X
��x�ߒ�
�"��T{��M{N2f�^q��\�i����E�<}ܶXt����}t<�GE0������L`��ۡ �}���ね�4�5Y6r�)A-�����Y�4�n��N~$�n���Hض[�.�L�j˨'��VV�Q����_�FG�+�=�ȃ�0rٴF���s�&^p+������]���ʻj
ч{���W9]�[ƃgy5�*{�`ՆQ�)���ub�;Mȏ8=�oU�A�Q�US�N
+������ܵ�����AWr�]uc�JO..풔�ו�6�D���Z��o�L�J��0O*�9>�JcU)~���k��ݗ��I[^���k>��˱��8�>�� �Fz��*||�=s�UP�Vo�ݾ�JSOH�1��Ͻ�H�1�١��_�|��+<�]wp�C��mW7�A/{��ܘ���A\�&*�=�Gܶ_�ł��� ��*���]V�1I�v�({34�+�Tb�|�$��``@oUk,�S��V�D{�C}��R��N��K6R��P�����ީ�x��������eK��m\l�v!�L�;W�ژ�5�r�o�� ��%/m��g,
��v��(T/>�T�VdBю���rų?�W};W��{�+�치��#PN�����|�P=��|Ү�Z7��ׁ�U,x_�	h���K8!��hTe�+�d�3��p���yyp�zK;��d܀�>]Ǯ7���d�˝h]/i-ԟ���G�B�λɒ�L�����зݑ�9�*.�AX���}bt�k5B]稂��3�� ��v�$֎�Oi�D�]Y`���ej�dzs(���±<jb�Z\�g�m�J\՛��v!o��LZb�̧٪�G^�9�#��&����ݢ�� ^9�����6� !��)T	�Z&�4��&��P�����{����'^��X+�o��+��Cg���<<�0�wB焺��I+���I<����#�f�pi��a�%��dƈaC��%C��ճB�]T���ӂ=�jK�l���go�WX��V�_�gq,ۛ#��ZL��8]͝L�Z�{�d]Ԣ����+o��c�w����`���Qvk~0��q��^�w"!��7, ��Q:v�/ W�������r|�����z�N�������?5�vc<+�1��p���b�fU���z��;�l�ex�c)��1O��F�?���V�o+�������=�����&b��7�I���[@׻�w^���C��ޘ�x��������]z����F<���MS9����Ӿކ��p���_���n���c�xRB��
*��<�x�N�T�r��B��I��^����v����X>�;�4/��Q^��#�'y�/��t�RR�����ijs>���F��Z�ւ�z,m����{.��s::!������٭����Zx)Ȫ�@*�3�\�4kk;@����WXJ�]�Vs�֬��˓���I�W
�Z��u�D��݇�	�r�u�i�!f*SM��^u$74\�Tv�b���Z)���:�V��
��!�`�A�� �Y:��r�^wZ�Y0�}�m�u�KJ>��X�k�ݑi��h
�G�Ҿ+_����\��lp��K�k�o�,���6�Nvĺ��Κ��V�����]XP"Q�l���2�!"�3�8/������ϓK}����M�W(�Lݒ:�e>���_ua
�C��&�����Ɣ�/J�U�f<W^]y{����fq�?�5ݕ��= �p�Ћ�����X��F�i��"QVl��=�qΕ~��r���c"�w���m��7�����m�d;�f�S%p}8%#V���~���q�"�����/�h]9�=p
_l��T$�=Z�ψ��7����ۓ^}��)b���s�i�~�����#��i#�Ⱥg�ҳ�ٹ�B�?T6�Ix<���n����}y��� ���s����~FV�=��N�k�e3^���K��\��܃�[=�ˈ�m�k��
��Y!>������9`L5P�V�MAɰ�[G1��b��υ���%�ȫj^`ι��Pvylq,��f%D����y��Y���be�i�D��#�X��VZ���� YB���Z����0�:�w�⬭���a괮p٣�ctVb��N)z�X*J}��l�µN�.��x�Z�����x�UPC��b6ޫ�>��&��`�n�_�I�
Ќ\6U_t���AX3`����sK��[����=��;�+�Q�qXϞ�1KӃ(�Bsこ�M��e�k2Ͷ�s�`�t����Ư��L@%3�r��*���뿏���zfۋ�ٞ5lyN����r�߷5���}�@]�\%
�<�ٔ�xV8��A��� ��G
����
��aD�\_���ϟ)7*�m�i��c�K�;k�B <߆S EG� nm��.��k.��=ɍ�f���]q��m}<��^|�\F4%��#g�h��vL��M�}��S��
ŭfR�nT����~�n�3T���z1)�1�Q�Iډ�~jHS�"o[�mX̙�>����h��l,7�1 ��Ze�Y~.c)5pŊ+��#E2P8���iީ�Dm?m��`F��L:��f�Z����c��5'
��N������0�|}/�ng3Rh�p@n�΁ � I�׳^�9�AJ��|��э�a"#�'0�;����˜�Ru� �+�����H��UV���"�����M�P��<��ua�]��WYI%u��]ג�s����e-3z�ъ��ӎ͕N6p����a�]�����k�Eԯ�j3��0�\l��	�Q�C	�-E�l�X�s)��z�mdg���Yݭe˜�/n�O��� hۈY��ƴ�]���nv!��(��.j�iv�֘yۉ�=x��{2��N e� ��IN�u1��ګteѭ� i����<|�d������śO1\��o5Ȼ淚�����g����|�ɭl��G�>i�{]�ڛN���APd�=�r�D��'��${TB��B�ۘaY�DM����O��*�[������g%8b�֓�*\�0��;�,Yn�8x��'WgiA��ar�g��+�Zeޛ��H�ۜsN<��1���ЬO��ֺ�f��|])Q� ��J:��*d�ŻI���O�̢��j�2�5�3�م�50tOb�٣W"�JQ{"�(l���w��h�ҙ���ۘ��jgCS[x��o�}Ηn0�����1�v��W����5�A��>!p�Ĺ@����K���mX��ʽsщ�*
�hzg�7:�Ol鼮2��}e4jPtiR�]�A�>�1�Z MBx����4kwC�}�L.<5�9f�r� $qf-���%�F`}o/��)�N�J]�%�jۙr�iR<�,;���s�Xor6�Qn����7#�8]�]֞+�!:sZ4]��Y�f ��J�c/8���񽋮^�G�SM��V�S<3�b��24Kɥ��JA��eȏCEi�G����"ڧ��U�X��i鸌����-��8s�D�Z�ΐ-v/�v�y}�1oj⺻���x�Ԍ�YLVWPۥ�-ͥP�{��Œ�S���:���QQ'��C�)uwۆ�Dp� �P�6w�c����{��Z�-:7td�vn�ON<��iYA�p3�I#>�S;�o:"Y��49��W�e�}�SPg5����|�ISKffԇD��9Ҭd��6��*[ys"tc5����Hc�p!A� �����ƕeD����&�owW�����B���3.�Zh v��a�Fd�'c�D������#Qw	j�]��ԫ2p�b�^�ұ%5:M��N5Y�o �`��y��tq����=��|�]�O��v����V[�IT�1�Y,�vn4n���B�p
����㱖�8**Gy���Zv�й8��T��	J���e�]�ǝ9f�S�H�]Z�ea�̜���)&�\�u������ -���ĦdY�����%�Ҹ��f:���=%ꅢ��
��Z����u*�=��uk.8�*���h����/v���p��w�Ҿ%�$��M �W�#S��6��f���C���A�W�5��2wֺ����}�~���EM�x�
�(���̈$�sPI�k7]0��v^M8x�p��*�Rh��]iAmkX��%��I%F��q�,�)	d\�aW�ܱ�w
0�.�r�$!DC���D��V��qe$�8Z�H{���U+1·�fsO6T�I\�#%8�]%��VEq[����DiȜ�P�j�����9ĝZE�8�uS�����Y��Hz$N��2.�ҭ�{��5m2��V+�^�F��Ȭۛ�ؑqU.�f���(��dj�f�d�8�7#.YBpNJY&�T*��ݖ�����jf�Z���y'*��î�S=U�Df*�n	�H�:��̌��q#���U��UI%0ļ�ez���WR15hHTQ�+N\�6����#�H�ե	2���\�}{(�t�E��X�ݥ��s;AQ�	ܭp���t�)�{SI��mP)��:Z+��;W-G�	��r�'wK��n����
�����/�}Qߩ�aT�}���$��&��Aղ��_�z
<@�v�t���巯p���F�O�k�o��`�0���oB�P��DCD[}_|Ǉ�}��!�^]~�E��ff{\������|�)�P��nN����F=;�ڭ�����~��aw��<�>[OĐ=��&��gF'�8���{M�97�N���r~���x�U�SO�������<���B��g<���b;]�|�ӝ�����x�n�[�o��w�������I�P�w������bw!�-�~&�����s���=�;�����p.<��'�>��@~y�����&�\�������_����T���e��0s����w�;x�Uǿ��&�'���y�7�99�۟���m�=8�I��������$'z�﴾�i�}�ސ�M}�v��'��㷈Rz�ב��MW	B�fo�g�%�C�>���}�Q�O>�~����o8������տ�o�7��=����=&|q�{������NL/���P���;��n�l�w?���UU1D}�
������L�R�l�F�B�d<��n�r."��#�� �0�G��x��v�?������~�I��o�����9P���97�'�����O�}|��%w�����}��ײַ�"D{�D�"#����nT�'r���S[���k��">��A�c`�<"�'!��7;�s�O�=��aW{p����L?#��&_��ېP���]����� |I�]�A����ӁM�	?5��6�����}�=�~{'UwO���5l�}#�>cDv���}���{�����?�zW�_>��O��C�k�7�<w��C����<L.��빓���0��|��<M�����A��}C��i���8�I����^�o��z<g�-Y�W�^����b"�"'jc���&���v�����;{O?~}�;z@����~v?]��ݧ��'��o����G&�w<�������&�y޺<w����z,���X�DH�!Z�휘�v�(��?%��� D`�;螟��v˧};��n@�v�{�������w��}��©�����8=�&��w�ϼ��ӷ����='뷏;۵��9�oiʟ�[ro�O�m�����Λ��IR�!�b1Ӕ3��=��y>���Ȗ0����������ãZװ��u���R��*���.碚��W{[�΍dj��lŜe���J����������%�:�4Bj�ޱ2����3�Lէs��Ǹ;�$�'=��$7*XğI�_w_���W�/�}G�[~�S���z�n�V��'z;�����{����0�^���}q��7������x���'��>�p|O��~�;/�hs��߽��$���ۘ|Ut�+�����H���>B�lzq�7�n@>!�������睃�o��o����ߧ��|@>~ؓ�o��;��P�����G�m����D����=�W�:��Z�|��G�H��荙��	7�$=o���nC���N��N?���v��'��<M���8���!�5����|������i�_�.k�|G�>����9�����}">˿>���G������WKחy��?U1_!�W�C��F'roן[���}O����{�����97�������7^&�e�xu��������x�-�����=&;^��ῐ��}G��d�s�ʩәѼɧ�x��`�|G��|��zO�o�;������9'���w����&������Ǥ�F'x�`��n~���#�;U��I�.�C��� ��hނ���>���M��~}�=���]�'c�1=�#��#����|�xG�G���>����D��Ȏ�����~��n���x��k������~ x��������1&�>'';s�#�{�N�'&��|w��nt�+���}��~��Q��od_�ͭJ�%��1��GQ�oi����k��+;���z��	90����=��������;��Г}BO�ߑ������}�z@�I�������DE�;]Q#�>�#��oٶ}
(#~�jgz��D���ӂ#��oi�ߎ��?��v���;O���%�����G�&��&���߁��&���ߜ�ӼNL/���>8���9�S��ѹE���-�a��S�������ߴD��6}]I7�|E��DDGgOуzw������NL.���[��~!ɇ����oJ��iߞX��'�oם�?��|I�v�����������z򏠏�}_}$��
B>�u��p�s57��y�����L}��?|E�Չ1_PU`"~��=&i���r{p��Ʌ��ǻ�?�~�&�ySx���C�~�w�$��?�'�w���c���!U^G��a�K=0�+,!�}�ҕ���i��n(K�Y�o��%����A��fz���]sQ" �G�KD�Eq���������f�r�Br��� ��j�s@խ}l��w���k�*e5Z �*�b�X��EnX�V�L�:�#n���p�ˊVx��۴zoh�V̵)N�Ǿ��p)�����v������ޝ�������>}�;Ӵ��{���G�8�ǣ�M�99n=j����{w$��'���~���N���9���n@�0D`�?=�着��>�޾J\}�7�r}�ߞ}v�@������}]���Ͼ��K��}��x��}Mz����c�?��&��?���N�q��<@��[~���݃�}w������|��`n�F5&f��~�VQ8����n�Npx��q������O���E�ϼ{C�a�m���oN��M�_��m�ӿ~[w���>��0�{OϾ��c{C�?>��~�r������~��$}�	e�H򨽃��Y���y_}�������S{w������;�1?��������<C��;�[z�?�y�$¨���=&��L4w��>8����$����O���o��M�9>�;����;<^(���q���}�#���9v}A&_���wX��N�q����܁�'��}v��8z���'o�{��_�;Ӵ�S{_��0�v�g��<����\J������o��9_؛�]N~���4&l�/����|���w�?��!�����{���w�=�8��Woo��S������۷��;��x����v���|O�K�����=&����������<>���}޶��nwMN���{;�"6߮��x��/v�����~+�M���>z�~!��bw��wv?q��������rs�w��׉�]�S�>��90����s�w��n@���;}t���Oo&�cAW�Q]�������aT����y��q���ߧ�|t}v�w�Ͽ�z@��������nސ>$�w����~+�M��?��nN�`��x�ڭ�������{v�<չ���� #�F�;�u#w�����_BG��L}=w�����9>�������'����9=��N@�>|��w���Ǵ;����te����߾m���;�߇��_����?wۏ��u8��0G�!,�^e���z��z���cm4�>.����|~���ފ�v��9Ƿ���S}O��=���y���q]����£�cDw�D廻f���.ޤǗ*"����B�I��e���,dw�93��3oN@[6���b��1[��R�ۼ� ��W[8��].Kgva���f�A�)���$Z4�O��-��:�n��}t���E{t"�]k	�x����k�!K��{����C9�L�+����m>���H��.�� dY4%b�!�g�'H ��(�k�{�]�6^�x��L���̢z�N#`��<h0��4���Oۛ#��3��PwQ��[�[��^#S���KI�����t��]9:zFZ��v�fU3^�W���	�C�&Tݐks�^e���U\���A�)�`au����U�u�z����O���W�:^��~VJ+���Q�/���yU�u�5]��b�ɸ�`������C3׮��:�Ǽ�;=~�8�I(�zu��}Y�V�������L�1Ew��׵��T�c=�P(TgN�iD�߁��7o�82MX��j�ϩ����y �7����*���뿏��k��i�4�j��\���^��f{��0W��!��@]��B�^��Ӊٔ�xŎM�,Y���wb-6�J�m�]�j<��� �����r�gә��3C>7lV�ഷ�l���
0z�;Oʷ��+�� 8^T��g��W�G�k�}�خ���4H����`n�\�����7�ޘ�i��s݂��VU��8��[7�9��k�;:��Ng���
�o`?Z�6��wQu*������&=�}������֭�z���A{�D1��v�9�j)�j ���囂�jÎ�u	�L�n.�C�(�j��3�H��-uM�o�l{ĕ"�p�uH?@�L��;ߛ�L�åLm���Y����$�K �Er���@�s�d`����p�H3�i�5%���1���`#L��3��i=�)��F��lU���� q���v�8Β��l�*S�J������h��A��_�	���6��31�yv��!�s6&�����5�qo�;�xR����.��Y�v�!��䥖�yzh�d��f /UA��S��0�D���JU��1���&nT �zSf/E�7q*��*yOqA#p,pW��6��k����dHB�L ��ā����QZs2֕8(C���a�׃�ۂ��5Pɨmւ��``�B��'v�*m��@"���ش�P�\��U?Y��v�={��l=�cwX��#V�%)�&�t�}�_@54�j�1:��(a-f8�������C���z�s!F�T����̝�� 溑饗H�۝7�xfZZ�ՔQ�3�C=Cf0���+-��Q|Q�:����Y�M�T����_���y�c�����up��e��aV2:���4�[W���;��5�݆�#an#����D�f+�yz7���(RMe-4,vó�"yV����P�M���u¶�W�uLձT=�P�Z̸�U�bdufq���i�>zz���/0��ǳ�2唣��"�c}M���y#��82Y�>�g.�P7h���۔���u�օ�H�?^/v��pl�;�:Ǿ��;��۬����{���c�T2��ϕVW��xo��r��$<p��lŮ��D��`\AA�-��8#Z�h�X�S��Z��򥕲�-�Ƃ�ƒ屢��g-�l��f��3���Yg)��&tE�!;�)�I���tԾ���)u���~M���ꠖ�.�S���j�6���CǼg��\.�?f���MSlQ=�]�n�8Q��~Deh�Wuhʦ׷�����鏮Ly��e�P�@����y�F��t��Y_|�M���ߞQ�)���>��SJ�:Ih�]u��c���g� O͘ʱ���-秃}��dW���c�\�Yuu7_�d���T|Cc;���G˸��o��='�-�9��\���I�iˊz��C7/O��=�р-ÚM7T\�" H���@�o'1��9��,�{�|#{ו�7�C���$Y>�Nr���Fۺ�$�ﶤ��t��{�Id�/Rnb����{z�f]+un�&���ݥG�d��Ŗ\�h�W.���wL�n��V��5��ƛ��t�ڈ�[ǫ���nU�ɳ�
�r��pR�L�b����+�J�}���Ǯ�|�-����ǌ�^��:��W�݈
��)�=�E���{���ED9�����|�^�� ��٠�=~�Fж�7�j~��2F����Kʸ �p�4����sYih���ཙT�3�&���_�3y�Ǹ��U��!�{����_k!��X��z˟�j�=>�[�"
"p���)�o�2!{�����?xg�������%!\��C��$2������]���E;~���9/|�{-�4!�:��b��)�y1N�����u����]�;~a�w*�?st�y���w/���V�����'@C��|������`��'�|}��	)建���xK��������S-�k��n�Q;ý��h�e�_OL0z�J�eG��?_{��`ei�^�z�v�9�K����iFlJ|��C��u��|7�|hm.{Ǯ��
��m3���]�x�x�pW��X��Ѻ�~�;aa�P�\��-1�t�݋||)���X�\�-�LN}L�r��,��T� f���3�����R�!Rʠ����P�R��@�3Zo6�v�S���J��
����ojF�/��Sj^a�#���V���@
n�77+(�����~i�9JI�WM��u�h�J�s=�L�9eSk��q�>��U$�2�s�f�Ħ����TWö��[����&����d�L�7����/�R}�;����WZJ(a'7�1���Jew�w���N��.�ؕ�53/y(�X4�G���{�ᯮ�)dk�^����U�ҹ 7�G@������k�z���]c�|<:���;�ٽ)¸����O�{$F�tE�;�Ey��D���r���&�Mx^'�e�H�	4�@ـ�T����`~�n�1�o%��s+��Q9%�׋����剟7�{w�=K͝3�@��?����|����>$���9j�;1�Y��kpm���SPuf��?tJ����Q=��k<�0F&B���nm��(r����/�-Sn�k��}��� �ុ�Z.��]���=��G���t�k�c5�kP];dKȞ�=��.��k��d�x����42�ȳa��J���.�(<lWR��Ke_mw6���z���6;A�)^}���a>����2�����C&n�0�h�WM�o��ػ�*��>��MV�ns�s�Q�ɕ�(��կ�zn������q���x����|���f��;s���㷴�&]�*��]��]����\wU^� ���u�7�7?}�ժ�k��$��6�_4%�Bqf�2�J��h�*}o��s[`;hf�foev̍��Mݘ��'Ԭ��S�Θllhv?�W�U���r_OR�����KEu�BՏF����ɗW��u��𿗛����Xʀ�we
�k��ݫǾՆ�/=ٞ50ݕf}ƀ�tUpB����q;1�`�	�W���[u0��uvuŬ=�ܘ�����("����s�f�9���'���qV�ഷ�n���^ץ/�/z�}-$�ސ=: �z�_�ϧ��t�7��o���������N��qtV����;������ݙ[g�B��P���c0�7p��t�����_v�j�K M^Oh�5IX�X[�n�Tz�*d!h�P�|Ԗ^@�e&��*m�khFaXE;��x��w�,>��*�pC�A�ZSS1����}4�<-�v�Ƥ�T&������3��������}m��^����:�̭\ G�S��{]���~��O^<4y=}�7�B��&���7�O��j!�D�s�a5��|vs��"k|��z���~����������^�_6� sn≂�0�_';F���mő��R���ܠ���X��Eh�ec�U�s��� ��E�һ��ڜw��.vʎ�)��)L��j�`��!u�21���Ϧ�oJU��jy7�����u���Cc~fա�u8�7qn��w�rZ���{�V�7�u��µ�~�����m�=|W�fY��~���a�U���Z�5��.��'����/����z7��ֱ�@�ROt������[����l���~��H��2d�&�~�:���(:ۊ�����5���C�����u�n��{"�;گM,�7�
5���pQ^ϼ�=@����S�e��f���2��u���g��@m�"�d
�s5�6>W�X8L�l��V���a[��Q��������?�L`9k��Z��}�����ꁻ5Қ�i�|<^�}��|{�7�t�Eӿ}s;ݾ��^�۬����~�$vҘ�l��B����<"����'�u�kܸ�
Ww��
�U(1���E���p�+$��(h vqx����8���������5iY�5^����/w�||r���+�Έ�\'p�C�^��[w��	�][�U����j6`
�L�rJىD}0��*�_l�e3pܦW�ڿ���������]P�*��%�"0�5��"���%�^��������#,F!-q���r~�WE@����ґ�h�p��TI�f��tQn���i�!Jָەۭ!�����M',c�c���;3�+��2�y�����9����WB���oY��u���;)wub��t{ħ3�>�1�n���Úx�U��۴�&���n�i���~HV��mb�i�ח�1!9�H33Q���CwW-�m0w=�2��
``�#����z�+<���Q����ke�wW��K�Vxڣ�;����j9� �릚m)��%+�<���6���YY��%�3/�����k��v�����d���:����3���^�\ ��c`m��q�CSKF��WtK�WU����E�g�YӨ���}PC��8�`�wٓ�B���(�k��������T7,
Q���F���|#�T�ܓ)hwQܮ4�L����㊮}��M�j����t�B"�h�A�pɢ	ln���!譃kq���_:+SH{����nZd�V(��Y���aV ������ϛ��DB�x��
y�pBv|�D���]5��.*v���QST�w�
tg3VwX��E������'�o�w9<xj5�{	�݉L��"MKzV��ʈ�}���o�CŮX�n0i,<��x�dԵ��	�7��� ݭ��p��F�ˏ���uK;m�Z1T[S�ZZ����� ({chX�2��l���sY�>���굎��]1t�:[JS����5��/E�pvS�ڀ����wB�5V�:�s��kt'�&՚��ҕ�l��<|D�Đ��Υ�뉗F[B+���:i�RشJ�Vc�I�h��Gv�
?.CE>��꘲S�˦fXm>�t􎫖s���_e���T��*T�]1��Mvn�]3;ە�J,��Ǹ�d�+v��Π̥�ʆ��bYw��d��:N.�Fu젞.m����^f��h/�f�"@�I��\�۲k��r���P��y�,�f/#��Φ�_��X�]Vƻ��k5���,��Y���0뢠1�E�	�f�L
�!q�mo@%���OF�M�}B^Y��`qf�Mi�A��qͧ��c��0�撢Bsu�@ϟYVx(�:�{t�@�ę����1m� ���8u����Tw�@����f9�mg�b�n\�ior�z��U=�L�+�FՃ�w*Mv�3(&鱭͙}KN_9���8� t Nk�I���կ
�����*��`���>*��ĭ�����q��b�%���P��ݪ�5`=�+{��C7�ľ���7����q�3j7��(��Ml�>Z=o�;�>Ү�*���u�@B�4��*��aZ�6��UN�Lx{Vͣ�f�Q�����#o2��B���
�WBgP���lYq��3�賀����f�9+����q�]G�3���Ƿ��[p���S�O%$�Վ�L9���9&:�u���kf�ܠQ���	lξ�_|�������׿}{��z��S#V�ME��4�(�L8�b(�E9fp҈�����&G5	Ui���;���ET�RYi[ ��[M�g#���e��)b	�S�����Wi ��P쵛**�\���DdEd�Ea)Uhg,�V��%n�����:&�*
Qm9rR�
.��
�����a"�Ib��U!3�a�$��Ҩ�V��KC.���(�,Ui���'BL!-I8PQR�N�2���(T#�y.mX�"��F:Vr�B���3U����*
0�BRɔhQH*��mZI�9�����K$6rT�+L��YlB�B-(,�Tje�	al9Ҕ̳��j	��:�)*�E:Ut����N�Ў�"�L9'�p�iА�9D�5����EB�P�%�U���y�[snix�������|�Pt  ��6B�\��P¥B�.�S��ҵ����Qη}n�D���6'��^����j��y'ޚj�g�Q�k�Uj�����d�K���v���d�k�b�N��y�%�Wx���i=��{���c4nf샌�9��OKv��")�mP�F@�� H���z����JƖ_�z�l�+�J�9[���y��oƀ�(p]^�gˀ p�`n�ў������P���*�V"�����~5���|�pCG��+���Fl;�4P�P�vr7F��q���g�z]{˹��� 0�^=�^���B[m9���^�^��]ܤ�qb��}��{�S����=��H��1�וx �6�;͹�:����Ғ�8��	=��x�N�
���鹙���RuJ���@w[�=t�]���U���.�ks���+�����5�Ǝ��a{�=��"Z� v���X��K's�o�9��g�d!�#o�M���m*�#Vt[�V#��fC�ZsB*5�Ԉ���`ߠ��}�K���3��ˑOs�$dE�����VR �ⓐ!��+��o�\>ʉ���>1���#Q��k۸��iY�,_!yԥw-�'g��*ڏ]hӽj2���!l����u.��P���Z��=�nB�3|��H����h�X1�ƾiw(m��)���k�o�t�6�=C�(1��仸�s���v�Ҡ%��fvkF��%N~�菢#��<��բ�As��W��ԉ��f�����;���ѫ�~��WF�!��.��O&y
�T�W�7>��[�j�Β�؟>Cچ+��}G]k0=���V�5B�bS/Vf��fu&Or�N���_�t�m�s�G�+�Z�8����s��>땉,�˝��Ɉĺ���^;/ܩ!4����M�@V����UQZ�Ji{A�컮�VU����R�H�ܞ���V�0ǭ� �����Uu�D���|�����Ou7@ܧ�s��{���w��g���u?W�����K1�(���e_K���0ωW��K�f�O��2s��K|����!3�t��6��(nu�����wP���m{U"C�с��y�pX��غ��~��& k�k:"�B�?o�`~�n�0��y�=�J���^ـT2�ή+L��(����,O�y��:���(o�1t���(mDl��T$�(�gD�W�de
1fe�
7J;�k��~螦�\�����GI�G�l�N�p���u�8P�
��^����,ELn3�I0|�X���M� �j�,�}I2l-u2�m�|�M4��k��WY����O¤�߲���=�9�ź���^�p�^s�!謄7��N���]5�e��F���i2%7��ngn&1d��"��
����U��WڟW���י~#G�+O���_�fX��Q�y�|��~FV�=�lUt�Z���.��k��N��N�5�:�J�6����#q�T7,/�M�r,����d��Aꪶ�W���TKW���o�g+��']Z�0![/:A*�����
���w�ZK���h�����_�8P�Wlm��g�~ɪ�0lO��?2��]������Bd�ȷ&�Hy���X0����+3O��f�j�j�F���K��r������^�X�A����<4[�L�r�Z~�/���U�6k��<8�����C�c�
�-�S��z!/=��B\�aN�����*����=�}9���@s#>7����"��'P�G�y�V�~�-�H�	��U��e�bê�ឍy<WR$9 n��c�Y8���(<q�u�?{�1z~�	���L/tɌýn�3�1�]h�JrL[����� m[�~�O%�R	)�L�Ρ�#DzJ���6�R�qN�{vOz�Y;l\���ÕO<��v�5{��Ws�
��W=ܻ����B���c�	]���7׮�}x̔2e&F1z�} @q�P��6���q5�fWk��f�1���sɅP�ϲ��ouƯ�R�%��+��_8 ~�2�g>beu:��������n�W�}U�}�S:d��{'�GOiX��"_Q8�@��T��Z��+U��)A����E6=�/|=�y!��Ʋo�q�z�N��w��Y�P@�tV��� *8�ڝ�<)}�灍�����7M@7����{�	���c`�*��Q�P�	�)V�N�dk����3s�pՉO����K��h3��a��RS��?E\LĎ�4i*�$��L�S�3��1����.��*�s%-�-�Ӯu���.S�`ܪ󙍀)����I�ً�g�|u|�c��5�8̬=��u���mA	ɒ��18��n+��l�챲v��u�P	ɋ\�F-�`�/-���]�a�]��n˕�U��1�~d����6��.�M0����T�g{�̠_���d��8Q:(�k�(*��B����{�:��Z��M'ə�T��,xqd7��"�-�0r�;����|o�>'�����5Ѫ���`�{�d�p�'�u�Yӻ�@���֊�����>�U{�n���߶����J�0#+��>���v�Ф�����R�60ef�W.���ۦ�"�����u��aJ�������w��%�u�)Ív(74��Wz���J�qR�*^�@yb��)L�R�Z�ۃ
����eϔQ��[g�m

+wښM^ds�Ho{��J�1'�![F�i]�]������:%%�e�xw�'|K�1�	�׶ǢUT0/�(1���E������1���V��dtv�̯yj����ǵ�^�DB�_K���(�;���r)��&tE�>N��&�yn��~�	ԩ�:*�F�D莂X=^�K�2���ھT3��o��2��.��S�Z|�k�Ǯ:����X�i{��z�:���
��Z�$}������~j�:u!�e�3�{Mk�l�>��8��y�U��a�\8i'��P>��SJ�?�Z5��e{]�B+�Z��o���m<r�8����,�]]M��d����mPUe{�s)��g1�[�=�Yٽ6�3�F����%9ϥh�r��9��#8ʿ*�y1�{�,� ��f�fx�Qtl�ìԗ�N�W���|&����IO�4S��p۹p�D�FSQ6�N��c����	V��Č�&C��9�_0;�Ϩ�i�a�v�v�x�,�-�G��cD1ng̔�&�«�e���ܶ�i�<X�K��R#�P��^[��l\Knl��ZL�h�MU�&$�x{�8M3n����_O�QC6�9zVݒ
�����30��
���pT^>~2}�����=�ۡPMyg�-��
}Ӯv��70]{h]&t	2Jԇ�Eoc�J���G{XYf�խ�����v�M<Bt���Hd�ꡉ=3{�W�����]C�6��&�@*��Cή�y�@~�~G��_mf��u`���WZ�-�J���q����)<��8Z��XL�3M� ;F~�qꁥ��o+��h|<{1/{��2���p,��� �����a�.��pT��*<�J�&)���B�a�:���|}��i9+Ӂ�ӯd���k`���ҵ}��(�� ��N��L�X�e�7�Q#�{=$�}�[��˯'�,^���X��[8T��
e��]��p�w�{h9�l����'&dn�t�&���vc���7).�~_sJ3aqէ ����'�xU�9���S�1��ME��a�`��]�jW�X:eP�+u��?����B��!�eL{b�~��nz�dk���&�� �^�#�NS+��5�4׽�֝���v�Ek����^p{��^�O�E.���v����x�^�������U}�(��Z�F��G��' >)	ī��'�r��Fr��w�-�L}6����ݒ:¯�S��]}Ƙ���	���W�^�A9�c���D�԰Q�xsޏ=x7Ն���L��ѣ׎���r����eH�[�@3���
^��m���ܻ�"�w:M��9�V�k&J�f�2#G����C$�C�P��r���m3�%���Q;9�>�����e&5�� g�� ��5FBgk]Ei�w��Ja���u���s���t<'�y��+m����u�F�t��s����EJ��"�;��x�}`��i���X���:��R$jv�Դe7UR%�# V�@�@�1*�*�Ӄ�g{/
Ua���[�k|����a�j�>�c̗�������'�ejDw@��H��*��;���j#�rސ=�s���FHA�g���ZK�3,~�#�Jt��Q�`0e�"�Ȇ��ބ��xO��v>g��5bӷZ)}��/��qVxx�X.��E��J�s׮�S=�z���>(z��s4�1��*<�
�]�F'@97����P��IȨ���Ǣ�kv��.g`��mg���j�~���'��YG�&W���կ�����%�83���J��}'<f[�b��{ʬ+3��f�5V:U5~?6L��_�����<���-i��/j{ܘ=z��k��7�s���1G�g�%�U�P�i��q;2�/1�7��>@�U�z��	�"��"�]�Y[c�T�if��bb�<�zI��F���u��RL�wz�V��x*�KBP�o��=�����WS���X���Z*tD���]�	L��w1w��m���-�=!���+���ҭ�����>���(Ǉ%+imF-���R~��Q�w��}�n��oV\�D 9��n��Mmsu`:�J��z�?v��}�8��J�O���w�������{2Y���j����@���]�u��Zؾ%WR��V���8����e��Q�YT���L��;��1p�S�]sB�I�kG�-�f`�f{F���!��~����uѤ4S�|7��K�}����5%���@�f�qӸ��Y�ufƮ�%p�S��~�D��Pՠ�}ܩ[�ϗ˹p��T�쭈Y����vrx��5�OR�-�mz�ư�>2��̭�p�qo�;��i�pJ@װ����zH��R�޳�/��a.<���*~�70�D������좱�U��<�~��y�S�AV�<�������0��%�>y��J�����`�?ݦ����n���ym<�_M�_H�̿�>獼yd�7�8
C5��!�ݰS��V�<y�.wVX���*�"�Ŝ_*��|i��8�F��jڂ))L�6��5�=�h��(�ef��K��]ֺ�B�wJx�zr��7�\-ʅ��g[���� 춶��ċv"������*����G*���ut@u>�z��]G��6mLx���g��}Y�$���O�1�w5
����G���:�q�4n�n�8	�諭���>o'.>�wr���L���ժ�1x}���m��y@���cd(�/�x������L�4�uv$��2�s�V��}��6
��qWd�*�΍z͇��~50�c>� �$���?=~�(`ݜˇ��TE��.��7��hZpd���.]����l�����ԣ���-�b{�j�z�ږng��5ݾ����6� >o~��$v��c��
膊k#�gOt+��WN���B�IzN��a�/^�*�-d�'�.�W�l���ঽ�[�.��Տ��>���<��ek��>o�j��ѵ�6�D	��Z�9��Ý��΅��w=8ŇY~��F��ڰKUE`���:���ȟj���گ�/�����7�4ݬp�*�o'�>�x�<+`~��G�S�A�Exk�+��-z>�[�6�C�u�Js�z��ݺ���]��%=�t3�˕7m����3an���	�>�xJ��p�*��d�+(��+��i�3��.Kх$���A��=+�-:>��Ue���jF�p�r=���8m�y�Avh��..1:`!N�7I���A�B@=��9�4��3+�|po4��s��Vgvd�Ukq���w����u*!tn���%���Wħt��	򶕕6�y[�2�m��@\�ltuڐ
=g[ӹܹ΁������UUSo��ɽ�X�þ���W�K.*�+�ܽ>ߛ�3��*ߓ�����K0
o�����$H Hp>�`�TE���v��R�#�3�>��xm܍��6	b%��V��E^��l���>��������,zӱ�*��h��3!�
��Ş���B�R^��|V�&V+�>,yy�!�Dv�&-r�^^�\B������~]�.�NWN�z�+��krM3Z�R�Һ^�yf�s�z�_k�r=�����_�9�
�Xs2n%�Y�`Ng�4�է�n1�oю��k��]�.wA�@�epw.�Xǭ�r}����,�ZxԞ�~�ޯ���f���F/��A�+�e>�
��qb{꾏k-�V�Of�|`���S���=����K���m/c�r�P�kJ�iG����2��B_d���������Gyt�����k�+��u���Y��׶�ݜ�b��臷��+k���Զ�B����%�����|��m�ܶ7��R]WXmq�_Ѯ����{�].�Z �
��u,ޮF���T��@�g�]u/A[�//$[t�5��M�Pvh��͈KJ����wv�Y�(S�=�@����u쭇;әs�v�)��'Xr��=ȝ���Y�� \)^�4q�V)-��+�(������_7WA[{,1Vi9,{6�MZ�̊�f�^5Q���h۵7�����|�ڤ^0&��/#�!�a�8�`:�8��Q�����tR���i7����8���4}:ڕe;n;����h4��.3{E�;od�T�g��v�����Ue7�"���6�G�]+�T�V��h��C0mv����D�� u�g�mصr���Q�1L�����eӀ>���8j�Jnk<� ��^�D�v�):�Ʌ������F� ��Ά\����^��u��i��Zy/�_c��� ˤ;�^���E�u(2n�Il�ӲE�3��(y�Bӥ�ڴ�`��M�ͬ)̰�T.��0�h#�;��R ����RCZ���N�0U=�2��	�1J}��-m�
O��C��,�ۦ"���Q@�|Ԝ������8qJ����놭�LE�$�*�!X��h���iŬ|�j8�d��y�Қ���NXH��͞�o���D3o�N��j�p'b�0�[�g��.�,%Jy/LN�a�
��j@ՇB˺�t�R6^�+{>�OA����<HE��]B]���qIO�h]
�#�	�u�y[z��;��R-�%�A7i�X��e��/�b�fc�138�B>�of֌Dm�5o��rX'vT��s��L�q2�����0�͑��;c�<u�r���:�I�B��{��Pa��y���e.@�T�ۅ�CE�k�j��XCNef�4�s��,T&7�,�Pk�iӭ�m4W'r.�M���E�����xF�*s����<�������{�mFH����s����e�e>|hm�ݨF�k�2�epq�겤|k�qm�!�_)�o�I���ԛ�kU-�X���V5��E꩗I�\�1@��Ճ�W=�W�B�y6m�Q�����o
<�
G(���j�������o����%GB�7�e�N�_wףx^/(5��`]Ӥ��X���א���b��$\�����>�}x����C�P���׺��F\%R�ۖ�loMp����X��]��U�6�%k��o�n��x�٬hY`s�k{+i���n¾\����*��Z�]�9.�Jv�^a�yow��=F�7sMJ��d+p�suW-۫�[�d���FR8���S�Ҋ�Ei��9W�8�ey�J��XL̤E��kgZr��M�H����N�z���U5�g�yE{R���zS����"�.w�(���o�'���3��f\������
�ޮ7b�5�T�lR3�.����C�����AD��2��*Ŕ$P� ��"�D�s�Z�cݧ�fY)ڢ�����I*�E(�E�R���	r��̺af�dDY�"f����3�U��̩I3�U�'JM��T$DT�@�-�Ows�	�DEP��22�L�D��eЍ.uB���)�m
D5�X"E�$A���gJ����T)%$�& ��gJȲ�Ԃ�U�7wshT����4�e�J�2銤jJi&���9(F��А�d�%�&ʚ��TJ��)f�ҍY*���U	D�����N��Q��0����,�,.R�R�H��S"�k$��r�H��]"�\��"���%�T+�\�ft�\�T�����$���\�4�"**j%a�zp�BGE"�E�E34�sY�5=q�5�YFeE�I9G4֊VE$�M�T�"2�V�I���U(�͹Ĩ%iEejQXRs���y���IXU�t,c�dO`43%r���u$+{{�<+�0�A͕�"�B}�ؽ�P�@�G)c-�2�<jݩ.9�+���n�/{���꯾��Ψ�q����U��"����m<^;qV7j
��%ΕM5��Y�{�(t�-&�d͸�??-n}�V�^ڛ�՝حf
ـu&�l�$2b��q+o�-�󛅵%+���߮'�Sͅ7���K@�r4Y��AeY{�e��?Y�'uڵR�?<|�x[���X��Z]��F��wP���ܜ�蟃J�N�jצ����Xֽ�naKW�k/�[+��bW2)��4,%�$c!(���l,����҃�5��������l������#�����{u�ARF��~��&�V?\���`}uC�r)��[��P���L=��~�sNh�f�H[Q�+����|��(��wX��R.e��OгCլ�6�6y�p�;b�*٨�!�w��eת�󔷒��/�'�ݸ���Υ�ڔ�֓�m�;
}OE�:��s���W�D?���H��U�R�7��P��rMT�Ɯ��4�VE+pj����x�P'��N�+*�^�B��&��z��N%W�����W�����l!�0w ,��h��2	����p�tk������wmp�(����V�vR����@�W���U��K�r�	��z��Y��^�\�����z��V�Hg�Maa��T��{���Q��g�m.EVr����V�2g��W��I����!Q�ݐ�/?d�k�ݮ�X�����-.�����ҝ\Ml��mI�}8)=o�cv}�~5^���Z��.6J�ƽ9VIb��_^ݛ�g�W�l�򜌵\��}%�	��hw�E^�sܤ���d:F��V����=Bz�_�	~�שb�S���y�׊�խʊm�;~���_<^:���w>Vu�{9/ @LҘ]I[R�R�֌lW�~��O\��]E^�N�C9<��R�1��`t�X$߳=8����;�!�)��N1�uD��T��x7�|B�����?��>V�8ݝ�獏\��/a���կE���z���Xy��2*Q15���Ԓ,Z�����*vvۺ�mHqYܬ���q�jv]��6.�W%��T�,�aNK���u	�
4�oF�i
m�XM�5Q���+#eA�_Z��qu-.�Q�F zgw!p��>v<m�ܵ\��OR�a��v][�o$�^�"�]Jq���}��U}_{�ϸZ����{�4�n�#���[c+�uJi�>�܅d��;}��6��������S��1���!&���o��Co"��f����K-E���_��@��|��{$����%��oCb�z��*02��~���y��{Vw��[�2��5�qUM��jt��ޱ�%�>���'h�7=�Ua�k�={Y]���}6�������rϣ��)�X%,'�+f,��K�|\/d#M����dy�P-ey5����y`�j��i�w,>[��Ͼ祚��2���}�	�w���XMS����Z]�9bϢ�ϭgSZ����ՑZ�]��L�g��ރ���mmw��j+J۳V�-�'G������v��$�Gկ����ü�.�p׹F��WM�p�aӴu��uX���K�W�*���6�TOۯ[��ߣ}�U������yNbYɯ�[:�����V]i�X�����n�$K��WMjʁR��C^�<�@�i�Nǁ}1~2��Ѝ�0�k��Y�g&�M�P�/�l�T���W��R3�ȹ&Ԕ�A���*��vX�Ŧo���4ʧ�7S���V!F�����.&t0ڛ�g�|�:nMj��zmR��^�/�z���^7���ez���j�ed��k[n��mY{�l�^�3�ȫ3Ӓ�X}��	�VV��bN���Ӂ��<��~�M<
�la�T�0]
�NW��z,��׫�t*8�����,��5��;�3�9�?W�jy���:�u�V�J�q"��Լ����JV��>{���l^C�SoЖlo�I���6'>I��\O�ٿ�Ɉ�򯔽�/c�1^!T��
S���_�xʛ�JeK��
�dv��5�Ԭ~����:�d��_���ⷤ����Jk΋�����&�4T��-�Sc�����w�_K��6������z�W�O6o=�r�I����/D�'�V��{�2� �]��@8"_n��#����{���s|�5*5�2ۏ4��q��ghR�=������[ף����LG7���gYW&�d�q��j�_m�5��$*\�Gĕ�:��.��y����&f�X��¶�[VF�edu7��ҟ 5�N	Y9�Mu>˖0 ΀��F�o=��7ҕkuwF�AM����3W�Q�������j�.�)w�sw�g�܋���+V�2{Y�ޯ��O���{�.O[��Imއ߯�8=Cs�Z��-�<�m)�կ�	�]ޥ�!���ḩ�Sp�?F�'�/�<���߭+�V�:Q[[�[�Υs��yo���N׈5��}k<���2%v'̿W�A�V����N�Ë~ίM�]Dʃh�N��C���!��f���ކ|���M4]_�<׊����a��ugnK.�bH1�Ȝ+˻v=L9�x�Lo��>��j�k�S{M�!�w0t�+5{nޥ���%�㏻���oj'!:�d��?���=r�lB��xl'��̧���#��U�
�%�@N��In��V�T�,O.!�k-�y_Q��ߜ�frW�$�nw�W�����ϷE��+^�V�^{��t"��j�MV�H�~{���zǪ!�5pσ_j�L_w�zc���T^~ޫ�=^	N��'[K�ש�Y�;�ֲ�:���[K����@�!���&�u.g5B�Ye��%oT�vW]�&�ܨ�M�yn�ĪW*�b�f��L�Ð:�WG��-�V��X-W�-���mBL췴�g�>jY`����=�_UW�_-�ڰ'mr�.|ȬYmݸ���Kt�D��s�~�B���&�=|�G�[�9]�=^՚�)�t:����/C�ldBo�Qi�yx�#���VpK�]7ռ����#�s{�74:լ��4ˌv��S�*
�H8�e�q���7t��s�8�h�Z<�-�\fu�J	[�$��|�.F����@�G��:�ܲ�z�x��U{&�[<"*���irʏOs��.�xX���n��}�
Y���g��r�p��{8j���x���U)�Y��q�����Ė�C�����y�||��<�?��b4�imJK�|����o��i��÷--��冽�=Ƈg������qz5�/%��qϨ=WQZkR���Jw~�D�M�[{�;��Ԭ�=/D����{��r�����q^<�8^C*߽�x�W/qo�n,�WG<�k�D������V�}��D)yj�7y�­2��9��I8]uf<s�l��ea���=�egɠu��[}������e%�F��z���j<zSk�2t\�֨ns�0��W��웽4g ��:X�9��k�Ac
P�U�uDQɜ��-��Γ��̻b����=��	�?}UUU�����Y��U��`d���KңV,��cb��oͧ�n=,��[�����v����������Q����K�Һ.N���c�M��#�5r]���G��:r��[x,,�Z�9n�*���NԺB�k��=�;��y�#�~�-M�z=P�7x|B�T��?�1`q�M��'�{۞{��6�����O�]�>G�s��{������7!�/����aR,m�Y�;�fr6�Kb�@N�@�۸7�|�J��7�s¾m�S�r/}(��M1��3�3b\l�u��?�J˿�}�%��oC�g�8��f�K$_,2���UHܮy���[GZ��Ήh�kW��[V�k�݆�Ӊ~�pwf'�������<�TL5l�{P2ۇ����k�7y�M��k}}��Z��Q�Nm��Dk�S��&1��k*�.��]�%�w�(���y��ΛN�l����k��B���*��3���$j�V��fP��N�H9ٻ�%����H�E���(�&�꜡�W]8Y�A>������@�y�!F��U���§Z�դ�[�x��$$�N���j���*v20_��������.���x�3��Z��&y�ޯ��N����IY�j���R�೤N]{pĺu������kW{)|hL�g��ރ��[�K���|7=�Vm�����p�3�b�w�Em{��}J��}-�C�]�����{(��ߢ�Y�q�=��A�+KG�U��U�^������VI��]��k0*�I<�9��=1��-i��J��u1���9��t��X��@��n<%��7:b�)2���{��}��?{g���mY{�l���7F�ƭ�����ٗ��.K7:2�;���ߞ���j�-����G�1���wUk�JG�[�ǫ�W�dyk�Z�Ҕ��k���[��黌>
XY�l�+�L�a�����~�?��T���y4�n�G���.z�Wo�؇�h�y��K&_�r2�ڤ��LOfm��)i[7�簻s�J��n�cU�/�]���M�0��?c��ߵ0nJ�����ݻ���<�[�k�.T��$��]�x����^�^H�FBa�C� �a��hF�`�"v����B\-�K53(l�qnEt��f�9ܫ2ef,��8�����ꪪ\�!Z��Z4le���F��[B0�{%g���3��P��صHd�'@�;�
�n3��~��:sQK5�-�RS�o��c�sq���W�y3E'��w6��5�I�pˌv�S�����^�ˌ]�=9�l{q�X4�{���Uck6�r���Iش�m�;�g����L��F����.�z�Gqwl+�|^�Ks˛���Zx��f�z�4�|x!�o3y�t&�49���{�+�;�}g��Z^߰�o���Ҟ�Z��&y�S�"����+W�4�-�R9�������/b=����R\�ÈO�UG՟#��[��	J�&JHo��+�ܘ��Rw�9觙!��i_i���Ëj��Ӥ�f��^���o;m%�a��(���M5�~˄�i��Ӧ��ƭ��W��t�I�[X��>���\c����q��Z���m�u�n��k�m�}^���Oq���wC�/�ʲ{z�<�J��W���2�mÒz�lʫh`ɵkҡ䧛�>�UCz��NfEԑޝ}�`}4Cw,�*��l0k��0B1N�Cz�NF�4�y��!���h`��ykʔzj�X������n�lJ�I�=D�ɝ�UW�y���vRkv��]Ԗ�v5��J�cwo~����Tާ�C�����/{��F�l[��2NA���$�_D��R�^O��k-�y���pO�M���3�%,��mv��Ռgۯ/�O�j�T�%BۥY���X������_����޵��������*��*���W��q���<�bSt�v��f�{��Ⳳ��z��^o��y{�o��o�?D.�ͭ�~{���{�،ԧva�I��z�~a7q�i�D,�j�Ҩ��榼�+l�il�J��_���
�5k5��e�;�}	�b�z��ag 1[x���P(;�Գ�5��w�m.Y�~];�O���mǝb�`zC��k'�k3)�ZR8�|%*�N=����n].�'}{������2���q�~��{;qE��^�[T�Hn��̫=).y���kiOz�����B~��l's���^��Ʒ�����i�#��7\O7�w���Wl޾��4��ٺ�����M��Xw�Cr'�+�4�lb��9�:t���wx� ���wr����xo�tA��J�B�!E
�)�×� �848�[x��];��꼤�� �%������|�.����Q^h��gm;nsY]�u+��ɢ�lE\!:0-=9��>�A��f�Za^�t#��Y�(����n�y���6�������V�Xu�TFE�7��aT�L;C�J	�nfJ57��ʌ�x�J/�z,����"�ϖ��T�YhBxc��.Gנ*���٘���u��d�ps��E�}��^I�]����9١�Ku��L��ʫ�D�#�S�K�@i�Fɺ��<�y��dXE�����j�:�c�:0v�"�|3a�7ʎ�X;:�5le�Ǖx�β�P���l��c��`�|z6�W��P�xL�;Q�;��ec���j�V_i�ve:V�a�r��͛*>��Z8�'�1����4e�wV	�V�)�hK>�����1�^Z�\4�/t�R�J_ �'6.�=��+�䊱��%w�����!8+H`Nm]�(��F�J������/X׆�)�m�h2>�;�ʨ�ήu;�3�+���*y|�!SgDZ��;-5�؈
�j�YD*��j�p�O6��s�zqV�e�N N���8`�H's.t�V�b��=k�e�V>UWs�gw�O,ƆfdLi�e<bAST�g��s���R�P�s
���3�h�]���w�M���,e���u}����qL�X����%�6�5��`|��i�y]�<�7���Ǹr�l�T�{bG�=�I��7x��!n�{Du�B�3u���#rd���\��6f����	4U�$�=1d���m\�ȃ���ɹ}���lIx7:@b9�ev�H��"���݄ӎ_�t�.���VT���F�V��&#�4��Ir�j� �ܫg]��4.x�	+2�4�]�i�X�����Wy1�w��Xm\odHh&�%ͣ՚��pd�Ą��"3��YʦQr�[��Zo���r�˽S��p�JC�a]�3tv���zd�gFQΥA(�+��k@!�fR�r5�mձt4ɹd�;��e(�R�	A=�w��1c������52�Qa�әx3k�J8��k3�$�ȥ�ݐ����M�>��h�Z3k�r�J�:�D�'2`)�ag�0�����Lw8��[L+�7ub������"�e��ib�^���n���3pmb�NE��
}n�s��LޒS�s9�F��u`(L�ն۳�$\&ԇr�Z��丕L��*��
<�lSWS�2���`��k5�+��G՚���+|�[�9�;峹�E>�ٻk1^��^\��ȎXHk&[g �a\�ʾ���֮Eg0;]'2�Ӭ�+�i�Ѫ��sE�yKkC˝z,�:v_O#<s@�8�A�
�`YUEd�D�0�+J*9U�kC��U�*��K����a�ʹR�:�!���HŕR�VJHEpNma4U$#�euN\)B��+
:Y.�瓔������*��%��.TQTr&\"*��u6�����`dFM
�Xr��΅"�VE�"�NUU��DU!Ŝ(�:TI[U�(TW8F:DI���Z�\��-�!"�*2��p� ,���Y:�EtȠ�#��d���)$g+M3�5�er�*�JĽv9�)ȷ6D: ��##��g���-�wC.T:�' �UT��
��]-:y�vS9�m�V�t8&d�YNp��΂�4�SX���z$U�t9�㜢�^A�l"��HT] �"��Z�4�Ş���L�J'D�+V��ˉ
bQiHZҤ�239UT����$���������YĽխƦh����?s�r��x*�v�c�ۋ)`�{W�S�wV>L�u%�����9s%���Cs��� �}_}_}��/�{�/O&y�wdg�ާ���{!������_�-���-�w���bY4��z�kkbc�^��i�z_�Uz5�/%����r����nd��G���k��t�K՝.m}k�Ζ����ytU�'��^��?l�p���s{-�B��ڕ;R��y��Q����V�����&yrj��g��y�)]�����6b
�}*5R�j1��߼�K=j���������_�����ܪ��v��M����;zE�E��!�"xŵ9�����v�����i�m��|��tO��on}uD�e���qk~���s���5^���ԫz=I�x,<�}�~9Ӑɶ#}��K��^��OǑs����5�z5�Gv��:�5�b��{��τ��Fm<�>�b0�~B��vLo�*��Vϱ�3���s`��V@�S��q;�[�̬�a"�٢���BV�Y��=I�B�ց^rsjE�����"��������(������^vT�����10�vI�Zكza����[g:�*�q۩%�!mv1j�Eb��pw��rK��0mL���꯾����h��y�9��췾���FC{7�޸	�,�������qz�+�z� 7^QI'�`w���>�o^�>P_M��C��z<_����j�ϟ%^���;�������� /D��V�ا�2�
�z�?K�8���W.\;�k�[�X��Qi�-���>���N;�Ug�%�T��L漧���;���{��w�ģ4���Z|~�<�˽^�o�=�{��XO�։�U�:[��s�Ov�=W������؎�4&s�]�~>���6�哸`�d��E"��W�oZ���Ҿڇ�aŹ=r�R��O�=Dw�Io|A~r��7�)M�=<�[��s^߹���i_m[��ط:�6�uM�Ի�f1C�Ҝ��{�K��{bg��|�Ln�{�9�{muv�G.	�X�	2�*�\5���%�3lnĿ"��6�ۭ{joi���+@ق���Q/-���V���<��C#h[�*���`����/
䤝��vQx�Z��[��1�+=�,��Ѭ`��xl�[L��Z;��1�}Ue;��+"Z�+ZΡ��[���L��{ҕvz�3����o��iTL�ĸ���^U�H.��9ɂ3E6���)	�����}DM-c"woͭ��L��w)_����_<)4��Ղ�ϖ��V��u/��u�4%����uu?4��y
צ��놃X�?o��z���{�Mo�sQ����� �q0[qK�ֿbr���{���(��=�T<�=�4�y�̊j��MHU�B2�DNa����J��s#��;��/����M�ys�4\�o����s�;]
�7ڞs�Ii�Y/�keTuz�>�{s�.�����l-���t抖kH[6V9mD�y0y�� ��n�#;,�{��9}Z��BI�l��p�8����v�̀b~��L��{�݆�ꬑb�Q�x�RR��5��r��m�S_=1As�ǐ\&��R�+��O���g%�g/e��1^�[�}i�.-�9�DJgM���wy,�D闣[��zmZ\���kT��}px�~詑;����;����I݃������ Ɏ`�����z��w*�vO\C����3��L�S�W2�H��S{�x�QCS�B$��OFaGմ�+z� ��B�$��K��+a���*n��2�d<�������r��\e��bY����}�}	nzQ����v�_��΅��T>�Z����3�K�	d�kc��3��*����{vc92'ވ�hs��c�{\�2y��ih�_�ma���Uu�w=�G��^�����L?n�:��M=_K�e�'�|�tܚ8��_�9e��U�LW�qQD����nz�gmc�M�Y�i�����}�q���C]�o��r���{����ս�x�pk`'rV�J�K
[�x��On'�iJ��P�>'<�SnV���xl:z�A�!j�)T��R�ϖw���s�,\!o��V�:�"O�*�K��Ǘ�w|G��S�ϷE�I��Z����,�C7;��&���f���G������%C>�ڧ�~	DŹ��xjE����ևI7�G���{��f�硽�Q��:�5HU����$?lJ��I�g�oR�J\N�=p7w�Ou�/C���Bo�Ni�E���xnٜ��bx��ٻ�PE�y�U���-칌�H}2�[�� �Ӈ+[�IJ9��������Ѯt �8ز�o�oFĮ�ή�r�HNR9�ͽY�:'��9�7��J��"2nV>F=�S+DYݱJ�'_n]�z�Z�r�"�:c������'���{��6��X���R��^Nw4*�V�P����\c�}�/^9c�����5VU��w��ݏN��Ĺe7�ӻ��z�OV+���v�1U発�=qf�b�Kk"=�n�n���_Z��;y-'�V3�.ͧh�ֽ�y��E�+�n}Q�<j�1��҉�K~�V��������/$I�v���J��lU� jwQ ���4!3�Ye����9��j?UdV�zVR>�#�����?L�ϗ��k��l{w3z����a�^�3��ΔV�h�/Ծ�Z�q�S���ٰ�mn@�hl%$��ej���٠���g}*������[{��E���7�V�UF�N��k��"�?l��T:U�8=7�ꝼ=�V��u�/mͨ��8�����t��[�[�+@ك�C�F�e�
#�Jt8V�g��=X8]�biN�X�'Y��yץf�-o(Ǌ�n8�-v�ʍ����"�e�səq<�tեV���\ؖ����b'�/��}wki��N��6 h���*���� ��&_o0�hP'O,|�s�I3�+��r��������_W�wQ��O^�T�^��ކ�C��O,�o��Wh�Q�vp�Q���B7�7���n/l��M����MB��p�5�E�<�:n��:�}�rr�m�p�^���a?$�^����b7�%����Y�IZ��{v7L��^0�W�0�j߸b�����5`���,Ϸ�$Ҷ}�����#^EX�t������SuP�)���l��2��]Ӯ���R�o4�("^.�p�����\�?W��z뼼.�	w��or�s�nz,��EK�ӕ�B+|�0+W�����F�L�y��z'碫ݾ�W��V��6�4+�՞ۓ�㛋ۊkn_�ޟ�U��&��\6�ek�W�E���jv��T%�%<��/����^Ks����j���3�����G���{F�zo��)i��V1/jN�ڴ�22�{*����3�����L�iu����\A��З]Nl=��)Y��r_˹�+���zLh�K�Y���o���mu,̮�&�E��a�O5Ȫjڒ4�v���/q�2��J��#;[��&T�v��q:��Oqz��2����ޥ��V�[���oh7���ꪪ�fΓ����q�������T!���8�잹K���;'|u��A�9�Oj�%�t��:�j��my��ih�߳ط:�6�uEi�(a���1�<{���چs�:{�5�]���C����,>߰z37�-ґ��6�:��IH����Ju{=���V���7���wZ��7}���DսW����R*���{Q3�ڹJ�cw<����i��W�����P^ze����� K��E�Q%*�;��V�4Rh׺����J>����q�D�#Уy��K��S��������BQ0[EJʍ�ȕv��}�LCl����Tp�v�ib����uNj��ڄd%�'�a<����y�$��a�ޱ�w� ��=�z�
m���S���
�B߲5��JƟ��+�/>�@�~s�羣�~�Ou��;�|°��9��������(�R6��.���7��K�M4 #�T������\�@:hM�&#ۼ�ڮ>��^��AOh�pTcֈf��~�{o��E�Hc9{�ه���sfm�[�YI.�����]Թ��Z(`+�51Z��C�.��A=�z�ak:����Ȯ��}��&���.�&��ODK����csB��V�I0�C���]����۳��x�vL�_e�Q�!�{_��p��9�Y�.Y��v���ɣ>V�or�х
j�A�j6�*�v!ޫ�����%��̾Y��<d����g*��w#�)���Ɣ�᧙9I�-�xj����5=n�X�{���hz��f��i����;	����lb���m��{��\����ڨ]�Q[�����e&Ѡ�;n��L�����o*����d���~�E6���qϯөx.v��WV�G�/V��)T^��zz��^�~����gX�SJ��V�c��/�}ܛ��n,���oֳ��YS�[�Sm[�{p��`X'w6��pW�[�T���`d�݁�佨��JW������<��g.f0Ud;)�PR�ؐX/iǦ�����>z��)TD��ժ����PG��v�n%����gWȍ��X]�����Y{���R �4�Le�t��6�;�&a d��л8�{�/)�����nWH�	�9ۻ��bR�{B���͋Et[H<,>�J�q����A�=x��Τʱ�C9�n���w@�E�)�^�a�J�G�}QKG�W��9����z��߼~a_wӭS���r��Dt�*t׼ jOE�M�?t_zZ�}�[^��5����)�u1�`6rc���߶qnڭ�*j���~X축�x���
��r�S��^ߖ�Ơ(_�2�պ�D��w5;��w�Ou����?1P�U���ge\·mW��חSV�(;���7����sB��k4���q����7(�j}�v�͘p�lZt��ҳٿgyf�.YTߗ�ݢ�����L����&�*O��[�zY���|8��o�Ϸ"[����o�����c�e�6�W��8Z�.<�3Qm�����c��cf�JK�y-E����Þ�Z��2{Ԏ{����)���Rg��w���g�>ov��E�s���"��`��[yt]����h�{Y�kT�b>��V��~>��=���&Et�1���k՞F�d����J��7�Y�Nw�F�{�'�h����$zԩW�� -˧������u��0{Qk����I�nQ����w����\�W;,���C)A�ۦ��I���Z��j�<6b��qF�a{G\h9z3�KaK{�Τ� ژ�}_URZ7c�V9A����M�{�lm@�շs��ytU�'����6��%a\�z���7��pxGY�鶽Si�:{��mR�%���ܞ[Gȟ9�n����w�o�!�.�P�a��MΩ�VK8O��5��%zpo���6�ۤ����ke���U_�o�$�J���ϔY���V�����r���~z��<�M<�������)9/,��*�V��;�(�,MJ��Rq��k�JS�^k��{k�z=Q	�x,8r�nU7�������ᄖ��Lo�J+wb�ֽ��O�o��gʶG]yɞ��~��faDy����%���wd����&���|�ƷM2k"�eJ��[{��-��ĩ�Rl��#Of�V{�9��i��Y!=`���P1{ܐC�\�_zϯү�',z
�j4��2��sR���A�!�����+ލ�y�LQ���P��u��zfSC���]�����:��O%�OGb7�#y����h��/��qg�d��5,M\;�u)\�G���z���D;5e�	|Hձ�����]�W�ml������	wjB�1�[ύ��h3&�c��+mK���!8�9�.�vT�gufȷkOE�
�6Y��\e��ͺUj�K<��.8��p���B�����5�Ǝv��B�ܩa�\.�G��c&�uӂG����J�(����4��n����{@���qv�J�7��#/On� /m�� 4��hR��R�w5�Ѹ�<���!��4�����B��b��XÝ�w�ͧ�a�N�5������5f��-[̻�Wl��=6;qrm�(lo3�)��kI��Z�:j�U�E>߲��h�ef]��3KT�l*&�4���/�s<P!wg�訞�5�B6G��~�Й�X
�I׫���}v@t4���$�
o�I =IZlV�CF�;�D�#\u��V�X��'��)_!�v:Q:�IL�]Qu��l;��aF�Ԏ��h��ا3�|�m���|.(����Ԭ�}�D���2��s�b��G#2�E���9�{��PJ3��Sk_dι�R�����*��)��z�(eʙIN��oP�s���a!���Irړ#��t����.�|d{��.�e��V+�ŭ��4��O��D��*,�Tuv��(��16��lըJ��Z�j��9|�����)���,����� nQ�&�c�> ��xSۼY��kHn�A4c�� Nn�5�,�x֮�(����Q��$/�Z�jȎ���"���VY��+G41���Cܢ�y+��b�M(���R{*���u=�ښ��u��1�Nm�Еr����է�#4������.������٦u��b�F�.ƻ�H����J��j*]ѣ(���Ea�=��ۭ3#J�����z�+�ke�r;���k��0�wt�K]ia@���i2�1ӻ80��V�芼��9X��t!�50�����s�ܢ,�k��]ݸ�+���p.~�z3vK�P;H�ǝ�3Mp�*@��˱vN�̈�LX�	�b�F]
=��ȩGo#̰�n����BH�4^>�[U���o�޽�j��-��}��^�\� '�D�n��7�{Ձu4��v�R�xk]�uֶ�mv�#�Զ�5����.�MW��@�Bj�W���-�=ˋT��t�m㼨�C����@w���ٰ���fl��k/9�}�]���^��8��4������y����������+�E)J�$�+�P����央ܡ,6�ծ�]�X���W":̈́�ԦIE�d�Ԧ\qj�N�M�u�;�:YWo���hĲ��c]�X@ʵY�-
�T���kk�PJ�\R'N�'�Onm\��������߉����t�Hed��I2��%%%�',�-J�HZ�Y�d)B�%b��@��E����
%BD���iE�$]�SZJ��R�a�x�d���D$�w;���Qt�	"�$���@UC�n%�Ii�*)D��+KC��KȵB�e�tr�ۙ�"I!D����fUPU�ܓ�r�E5���()��r"�(.*�e�D����+������J9DI2�!
f��s�L� �T��V��Ш�"��d% ��J����B���{��"-,vY� ��2�R���!Q�9C����W�Z A(K,��Ⱥ��e�R����I!)\��A9�z$UP��U������DDF���!��m$��PY^xU�]*U�p,���DtU��U@�>�}�4�֭�o��NsAo>�H�5u�:�[r����ӳc	n�����D���Tμ��Wu%�3&����~�����;"����P�Ѥ��q���=�V�Ľ�x�TS����ʕ^��j�j�Rq9���?LnU��tm8g[p2�Ϫ�?g�_�e�y�R�^^�����VD�����嚴�3���W��}��=�c��^�R�ź�ʔX�^���JK�|�g+Z�؎�"g;5���\.lr�{�nir9������%��ih�^\�-��B���|'q��J��-�cb/�{�xvW��E]����g����Xssط:�כ�E����4�ٌcv%��j��S�Z~U��Ъ��S0K~��O�[��7�zwc�6�j[i�x�c[e?�@۝��nmD��~Ռmn��Ih�׊�+���~���Bi��U��ҍ�Bu�kY��4k��`1�AoO�%0n�*W%���_[���ɚ,Mz��0Ni\q8賠�k�WV�nn�AU�3�
�Nt�\�Z�'�7���Z�h�|x&����[�=ۻ�|G�����m�����).\�5f�ļL��Ŷ�0]�b��L�"Λ�����鳩ɗ�Rf�].�՛�~�b>W�;���ۜ���������,�<�w��՟�(�ҩ+Ք���V�'1���KwXm�Z����������SP܇K�S0������Yf�A*�T�Kq�m�){7����/P�x6ϳ�T�"��hF���w��v��L^�ew�޴��'~���e�w�>aX~��:sEK5�-Ǻ�g8ŇY�~��}Ayf��,�]���}�h�I�l��az&���iY&�6E���gu���o��8x���vK�N��cfD��ȡ�������������Y�T�	Y�Gxx��r�4�ej��Ok�����g�6� K��G���z�3��ף��>���|G&yߒ���-춶jUo����gg=m8�������˅������ҍOe�˖�ʕI����^��!��U�)���5ǽ��>��g��������#���
 6v��=�]9t~���W\�&����%�y���r�J�d��^��t�PQ�H,�a��b�,x�
�rmVنtQ�Ӝ���Y��J|4ԧR��t�ǯ��N�S����\j� z��0�x;z8�-�.0�V��M��L���X������j{9b�u���Ǐq�J]J.��zz��w�Vx�{�o�|���;Y����>�I쵾AN��;��k�c��Dx������Sm9מ����R��Ж}����K}K܄;.��5b*���ԼV�����7�M�*]�&�R�Ym:�w����t����������UD��z�\��z}��]�n)KU^i^��V\<*-�����XX��2*膕+5Y�`֦��O�[��f{՗.���Xֽ�ض꒶|/��23�J��y*���^Cnf�Σ�&+���_?3���D!;����z���[Nq���0��K��[��
�&�����?1I�F��͆3ՎL�hkͫ��s�L��#9�Y鯼�慚��m����Ag8}�����'L�Y��g���>�S�C���;�6�,o˞\3=����
G"ur�	��'�L��|C����⡓Q�C�Κ�~�}S�:{=ռ����u]���Q���u3���}d�!Es�^9x�l�[��S�S� �]GQ�C�8lr�,��d�A@�����]����좮N<�zpBkiq�;��VM��չ{�~���6��>����j�Q/c����z�y���dK��,�ڗ)ꪖ��^��\Ȕ�.s���}�z[,�iX�d���d��=;���dV�zf�>�y�.��xC�����i{#���MJ�Κ����s�W�n��"��z���*^��7��5�{ʲY3�����3[|&��q{���Ƥ��C�r�T�:
��\\AO�u�¯��n���˱G�W,ƱY١��U��R�J���6���̕�x*R�Sy|��rb)�����d*xί>B�]��l>���sa�[�6C���$�&i�ؗ�Ӷ��t��)���!�e������3��z?Odm-�󙵎��X߯硯\<)4�ʶ�0����48��u�Y�2xd6�w3N���F�_+^��)��kע�~����޶�;t��)-�kǰ_P�˛��}���9��=��δ�m�taK��6�	��W���|Ǫ�tKzI�Z�KlV� ����l�;F��'zb�IݵʻZV�ټC�����]�NW�lĩ����d���K��ɘ2ٜ�DA�X�|2�_�UQ愛ng3B�?��9j����l,��|�j;:C�z?y�N�g1Qc	秜�~~>��1����zi�
�|�������VN���iI��T�y�1^����GӋٞ�*���9�M���͹��-!n|#�9��Ү�:?�QԻ������fP�ե�����0��',z �f�����~��A-�I��b�����=^�LnhU��$�)��؀��TL5l���� �wO#Ә��׻�7�P^H�H�j�,�O���=���{�nx�J���m��G[�����H��m���D����i��Zxԙ�Wz�6��|\����=^�~��rY<y������=k,�ڴ�G��o˽���&s�;&fcTn�#�9/>��\?W�[_w��b����y�[Y=r�U�7y~�>���w6�����K~=(�C��w�sܦךA�V�����!U�޹��xu{+�C�%�7�սf�ٜ$�s�ȯ��Q�v�Tފn�I��ڳ�#�������}��Y�ݑ�Y��}�j{�;M6�h1����&��A�����w
���K�����m2�ܠ�S/��J���R_e�0VwFI�R����*<ˢ#�Y�⮼���=]ҽJR�N��:t��]�<�զ��Ɖ����'͙���wp�=�3�������<�|�s�����5���s�1�YO�w�T�m�7��7��{�;�佽)\�p1����[��4��n����=/_��xXN�� ��W�R���J�����_�n2��ǽup�U�D�y�/���n��ab�T�r@J$4�^�o����A_eXs)�k��"@�@�k���ʮݙ�;'�e
B䬫s�?��-�n�ٿz	�'���8��l��>ƽ�9�P�8�\��
�B߱�94�ڿ{o۶2l�6��.w��g}��Z�CL���N\��f�{�[q�*SNfw��V�<����g���0:���ˌwzP����-�^�CUz*/7�M�o��勊���wh�ޯ�z}ƞyJ�Kn#�`���dqT]������Y�zxh;��W�;�Ի�;:�Fs�[[U%٭�Yp�d�1v�)�fK�&�����L_Uʀ4Kp��K%�(�w|�e:��w[�.���4tU�{�����e��w���َ��^=���|�T���ߧ�*���-�������׮�.�dε_;s�78Պb�Q���^��=�{&�a��L��,{�-�xj��]�S��u���]�B|��NR�Nm4���S���$��}%����y�����ޣ�1�QwQ�c��ǘ���[������bc���R�\��bg�����i����~d�kZ^K;��;��_N%��mZ�eT].�:�Ŕ�^�u~�O��e�ܧ�GƷHj7\�l�o�t;��Gb�s��ֺ�k��{~*&7�[�m�j=4$���N�7��p�i��=�C[.��V'm`��ңU}%(����]W�ו�S�a����c[n��kV�
���"�=U"Sj�y�T��>نwJj�����=e�<*ެ�.ۼ>
�_j�9������7���-�W�#�_u+�R��y�_=����uI\C>�}�&�S�xy5���*��T�wӽ�)��{��i�ܿ���O����]�� U�bx;;�˶%_u���6+�>^~���������3�>^��ԫW���;;���W#Y�>�zj�A]L���^,��Xv79g	P�%��8�1f�c?}�D{)�3�m��O�q"��������-�q�<o<5��s.Mlm�}�}�v�uH���=S��b�<���Ks}�RM+����@~cu��^�'-�>|�q_�����{��t|��#������k6�{#��_N�	3��K���0ZQ�gl���9�4���״8�mA~��PƏe�K�i���qLq��k��j�יj�n�5���mǞ�Sꇢ�a�e\
{C-�N��W��W�.�{q�W=���U��U����D[p1�~�q�U��[s�B�q5���n��^�%�ƍmv��z��'1^�W�/.<�c�9g[�Ns�v�<��ܜ�_]ޯ�Jzor��{ڣ#���_�4���y���NX�c$���'q&{�,\l�!Ϫ�;p�=�/�T��7��U��>R#JOf����}��p��s~��!�q_i��.v�Cځ��柷e����,̈́�ʷ8�I[�`t4��2��1G�5�am`���Q`DX�i"R��
�/�2ƺ�(�ND��(��C������Q�u�Y3)��ά��,��Ń �XsJ=�혠����l+NJg��zJq���j����Ne\���胮ƻ���or��y=s�ڸu��v���v=Q�@�:G��%�Pk���ۻ��<{���u1�&�N���t�ڛ�K�j�]�t;�$�h���W5��9k�7�3�ڹR��؇��\<*O��,!zj���u�G_�xR$	q ��$$�$��Z�Ҕ�p�5����_[���ҬF�no-�Wn�w���}��/�{c~u��}����"�s����`�~����Ӫ�ui�a�z�S�sP܆�k FBQ_�,��`X��*@smEf�[䗼}Z/ۭ��m�1͹��,��ޘk9�=�}���V���U�o�y�?�p:kY�m�vϘwz��v4����ո��h{>c�=�����W�MG��3U�h�I�I��
��֭��Q-Ŋ�3��M���d�d��w�������Z��]���g���糹�||3��\��4�W�c�s�ȍ��"P�ń�aqy~����cв���?�t͝.�:Bn_m�x2\��+Ѷ���U{���jv�5�.�eٕ�XU�*�ޢ)����4�99��n@;m T�2�¹�X�1m�O�_V�V�r��֨��;�U���/Dq�V�<d�3K�^;}�߮��'��,��sݑA���{U�%����>���>�U��.��\{W�;��Rҽ9���qau��>>����kk��#���yp�D���jb��������颽����}�⟫ܦ��iyZ[C�[���faAC��a��~�b�Ն��J�n38�mS�\'�O���5��Xy���5��{ܡ�XD_EU��R��T�o�n[Oε�5���Gc�W���^-+/���>cv�0n�4Gj�P�>7w�<���[Oo��ڲ��k��Z�}z�������`=U%*�;��T�%��ݯ+�t\P�=r�VY�������R�o�黌>
�ڦA	|�!^�Ҹ�v+��]69w�m���M����l^|����u�S2���g���_(� ٗ{z� ���i�{��0G�`��P��#������:���hmu^Z�H�XX��v,k�l�8�-��#��3�J8��$�a�ܾ>#�ؙ����DbZ㫍p�3xiǙ�v�@�u3��r��s�b�Zų{`BT�� x���:�K&$�b��̫���XR`L�v^p�X�ɍX-^����UCg�׶ſ��O8>���g=�{BT��-�\��ԜU��^�}�1�k���)'NKF(v�-mqnaxl*�t�0���ٮ� M�������7�����؋�C�]3�;r5�A ��.൚A����28I���>��PM��+��n�)�۽KH�&�gy<no,�WK������T�j�c���ŉ=r7���#!�r��b���!AQ�n����;/e�s��Z�8�dh|,#'\���1�*��Ri���f�6p9`o+dy��C�9��aٔ��%;�fV+�-+�%�m��F�-�۳���-����׋{Z��J�Y�^潥��֋+VM:|u��,���w�*�]E=R�uև�A�sCɧ�vc���kF��������5�bkz��ލt�jZ�7��e=�`��$b"DU��|r�����3\�P�TU�'�:��3�6�Ҳlco8r�m�@~R��.�&3t۷t��\����ٝέ�*�	�kj;������ޡ������k��ݻ��=���M�w5%�1I��_LY�Zk�qɵ ��YHd��V��Yl	Q�ٛ'��dޭ�U�F�wb�{��ٴ��kJ��c8/�L�*.�nԣ`�[ �Ӥ�A��"2��
I����`��f�N�\}s�θ�Ǿ�Ft���{X�g������.��fGh�!����b�ܥ{
ɶ�C�kv�ǅ 8��y/I�:9����Ś�d����ىu;�i%��i�\sCiVS�ʺ�]�����3+����ro���;��tG�ޤ B�iҡ|�9�#A�C�.��9)W˶k��qp�TԨym٦�����a�<����đ��M���U����r�L�_�Y4��a�1�:��W�`�^�餜Y]e��	��\�Mr��e��q��F�U|�QZh��ӕ�dx-뇖'�B㡃W4D�0<���%p���0�tTT��r��F����o1gb$��i�ƣm3rZ�7�7�ր�i�J��rU`)*�;r#�I�f������c��sN���^<$+s�:�U��h3�1����.�S��G��;qU��$��ܹ�Hm�o3�4�/M Vnܕ):Ԃ�����4��w�T)`w��r�n�w�3S
���2.Z�h+�Ό�ői�ɽV��έ�2�	x���!�|q64��)�&��-u4;���
X�[��d�̓]���Ҧ,;��]���JYy�o5t�o��^`��c�YX���@�p�~�> ,W�B�y��WRR(�.^�P�J�qBP�y�򊂒)��W%9�VeEL��\*�;DQYJ�Ҍ骵2���P���eTp,2�R�.QE�dh�G����d��͠�)՜�,���L��6�$Lä� )�Rr��L-Y�e]�u�䜪�˝!:��qv�)d�H˲��ts+"�F�g*�6�!8�-�Y�B�\�.�ʓE�b�\*�%�DW
%��sp�E)�J�bF)���.��Q&��B�(�["wk�$�&\�2MD�T�Ke%Q�*1��˗-�D%H�Ȣ�ª���#�A�J����'")�T&\��O�I��� �Em�#��{���fuH=��H�gF���*e�����k���8c�v��>Amu�P�dwtQ�x���x\��v]�>����������v~~�h���-p�x6ϲS���*�d-/|}~����&��idK	ܕ�y���KZ�^��[�O�Ӛw���`
H���Aݾ�U[ܠ�I[s��{����܆��<��<������d#f�Ӌ�i\ۉz.�twzԛFG"6�=/k0��㕓�>����Л���{���?jԩbQ��"�����t+��he��e�F�e`6����;�����?@���)�qlfv^���~L��?�wz}���7��;�}t6�������A��Q���p�]�Jℓ~�b�nw���{�#_E��������Nq}�\){��^��9ư���'/��d42�b�s������_!R\�҉�S�lF{�����O����>�������s.t�y��~�f����o�̟h1��	�P�ßE9���`R�hq�w�{�uϥ��u�y�^��O]_�ȼ�ީ�O����E�T�7��6[�}2��� 5p2�p^�.����t��yΪ��^��Ȅ�p�܎�.B�cNP�kN�q`}���ͭs�st�ެ�w(>�-A�����r�����W�ݪ�e���L�=G0�#�Ɲ=
 ��o<ts��{_d��K�.:��v�뤵���VW,��4(�p�b�i��k����Kg܅�Deގ���B���!z�Q��-2���d8	��,/�c���Y��"��J�ɫ�ۇ����v�>S�\����>%��P$���&*�����{ȇ����`Pb��c_���i��M	���o�"x�=����p���q�F��Yp O~3�F����O�2�\�^�՘�J�^�����?:�W:v�7�m���*��u�ˎ��a�8�2m��u9��L��n��^�p@���\��� ��:�p=Θ}>��ӸJ��Ӭ({��I�y��`�=�+}7�]�GO��@Nv�����߾Y�!���O>Ȳ򫮸��^��ԍ9'��hV�r�f�FIh��������d��P�{�#��B1ǯ���m�Z��d��:
bXC5�S�_r��3��t�ة{X*�_��/����:,��R͟D�o5o=�r�{���q�/��q�����e�*>"�ׇK�*<鴧�����n��"L�Y4��M�j�2�Ve!W=��߮�W]�}���MǺzێ롗�Cٸ�Į�����gl��ra��+�[j�`:��U����Pp�\Ż�}qڰ�y�)%}1���3>7���/��7o0Կ>u����O4��gFx[�ᶱ�S�L�!v�U�Y/{�+^'V�t5��a�A�OX�).W�HZ�3ۥu��e�w��v��7��;c��X����ݳ�.�W��W+�8N\d�וV�J�}�Ft�Κ�+ݷ�X[��*���w��V׷����e|�7)g���Ss�*z1̼V��W��.��}λzy�6�\��H�w��g����[����.�{�8�Cu���-�73�I�O���6�P�i d�����k3�/a�t�!�NGvV��{h\Gk���s�P��e�ѝ�W]T��p9���>����Z�Im�����:\z������G�Wg���u�P��$��e�BgC�q�o'VOr�nKU�v���Hjo�i����Qe��/���q��漍㕆Y�֤��נZ�fV�
κ'6�jY���]OSU)t����{����u1���<v�;��D^��G(����y�)�@���%�A�`���l��2��??`���xls��Vr��L�%�g�b����Xr��=^=���m��h��u�:�1�&t Ҹ��M,��tאP����U����c�lc�V$v�|w��CI��wQ�T�guQ�@�d�P+�^~�L=>|i�w-���9�qxdB^[N��28+#�;�`�f3�#��$=����Oޢ�X�[�:BR�{�j�@g������__\-����E��1�Y�6��L�4�w)դ/��7�.�l-��oH0ѩ0m�J�KSc����e)���WSs�6]������L��sOqΝ������5��b�Ij@}�!V�z*0�W����)m���A�9��h��m_I���OGL����c�$s�r�R׵�	��� oCv��޶�{ç'�ДW�dd����!�Bj�L_;�&����Q�Q�B����Q�d��z��a�)A��;��3�������s�j�X����1�]w"��>��7�<�����yʱ箒^�tz�=����T2c��Na�q]Y��(�=��i�y~�<�Wi�T�.iB̬�W�~��Jv�x�Cڱ����/��ٗ/w���g-��3%��n|���8n0�3u���u��E���Unj]?={���Ҫ�I�:�}ʫ�/}۾�>��9�8��_�A���+�Xp�n`gGU/<��Y�^��p�A�����. z_V2���q�ʽ��OdΏ<��.e�zT�5��2w��Hyஊ����G)XF;�P�Z��.�+�;��>�f/���=���[lS���k|�"m�b�,w�2ѺrW&�/w TB�z�W�;��^�9w�{nM��za�9��@f�PΨ�,���{(Ǻn�;�ږQ�V�ّ�j!�}ٯ� {X�˔W�t�	W��>���`O#�3l	~.���E����$ڕu��{�w$ze�0�l9�����]�Ky���a�Hp	\%c�W+����5�R�k��3��O0��~z+���s�UDp%Q��hʦ$��ET�O��t~�ou�{�Oq��T�&����m��������X��� ��(�p�$�3O*�Q���S(..ߪ*j<_Y��:<��,�{��jJs��C£ܨ���|;Ѧp�9 '5'@��@�-��xs]q��㓑��N�k�g�}���Ӵ��s9�i��8Uǻ����f�;���nE�L���^U��f<=�U�y��֮W@�Z��^���Y���뭳�;g#�w	���ێ��4.]QgJ�:���{)�%)�7�{�@���4/���9����d;���c�t��q��.�ܮu���g�ѫ�W�]�Y'�!�9F6'����E�����:�j���܋��q=Q��{�B�'����k3U]�U��n0
���t��dr6v�:^טm�~8����_ݿ�~��h��z/�*s����I�@9��O0P��-���?%��`��G�J�a�2�����NwVl�y�G#g�u*ZJ����o���±��}�<'6]�&�k#g�Dx�Q���9�^��TJϬ{�4�W�W{���SS�#��?m WW/�C��7�e�W}Y�����FmdPN���W�=A3 ��d�kP>wPC%��7�8ViVD�_j�Vp����1��÷v�]��+�sEZ�F[T��]��p1C��ueo3�����!�T�|�/k��Ȯ<�.H��������;����׫*8��'y2�ow��7�~��XX�}>[��xLp^u�u5�7W�.p;��JQ9q��
��/G}.�z���>������o8��=qZ��.d�f�{*ͯB=���b�Y�#���Ma��r(�`g��E��ށ�uϥ�
|4p�o�R�޻�k�h��s��{*tX$�u�l�G���Q�#����d��z��^�13�<�:^��T�E��߾�8/:��q�*_�KAȟ�R�M$y�s:�wi��uytu�� ��K2����x�#�O�v�>S�\�z�~�3�[(V���a�%�g�����=���򽘓r�������,V��9I���;d���+��=^���87	�Y�D�1����-���:@>ޘ����}�?:�W�����[G9I¯��.#��qp�ԍӷ��yn��q�5Ɗ�|d�q�;+�ׁcig^���l{�m����/lTk����[x������w�K�,�" r� h�h�����W�7�1m�}��[�I9�e�X:�<s�Q�3�2I!��;��~�;��cml�~�܏v[kR�"��Թ:�-{G�aõ�8R�Xtm�ɸޅ����`�XJ�G_**�����Bh^���\���\6*j����x��v["V��+.f�Г;)N�����g�J�D��	��Z�_z*��t�����׵�n�ӕyP���TU�w�v�5��יc�v'jM�wR�Ƹ�����.o�c>S'�����R��]z��sT�/_���]�G�'>Y�ۖ��R����Gx ���@oz��M��s��>�s�[Յ{�~�t�i�f�{R���T�K)���^[~�z��(�}�}ǁ����0͟|��gs���{���Nt@S����W�����'0���(J�}�Ft���2��gU2Kqf���U�_G�����G�2�nS��`��Zz1̼V��{������L}�a��w�~���Rq���g�ˎb��{T���5�w>*�˪>�]>v�<7(Z��s����������{۽�:qW"=.�cQ��N��ov�zo��9��,�u�k���|}V�G�q�ip�M�w�#�׽��ǥ��I��՗����\f���|���'��� ���l3��s�a�yqw8��=�S>S[!���f��|7�<���ﻥ�^��q��k��+�Y�� �Jt?Y��{� ��jm�(�R��m��"�jX� �1笆�=��
5tD�9ly\{���d�1�&���'�8sL��C�x]gwe��N^��N]��5�m}�J�c��}�j�eP��m���B�7E'Ӂ��qv^�f�lqBV��[�[���3�@x���:�R�	�ӝ��h:�{����u1��;h�ۈ|�;}J��֍�y95z�{�T���f����� �H���ْP]�??`���xs��v�=�
W^���Hמ�k&�ٮ���_i�<o�D� �l ܁geqU�0���ۊ��5ѝ�"�<�I����>v;�9Z��Gu!��{��ێ��*㺨��2 � !����<�S�6��pOFfg-��7�&wu�}�9���N�q�נ_��^�W�b�T�� 5��p�uў�t�W�}�T�1]+���jh��m_I��D��t�q=||���/��}�C�Ӟ5Sz9�EO9�}�npU`��het�5d�5��Q5U&5��d�ϧ�ox:������*��]�c]�Z��<@��VI��J��Y^�x׋kn�����~}C�fx������I�4�{@5��Ea��ʁQ��T2a��'0ÿ��0����m1��/���Ce�e�z}Q�wÚ�=��ݪ�3{��Nϡ����vg�{ѳ��D{�k��2��A���is�4=��; T4��0��F䨟8OdF����}0�eP�@��[!$���)�]
Ĥ;��.o��E��9�)<�rQH�4�n�<����!o\�4����e&�����ٟow0U�_eE�׫w�8[W�/"wjD;>�Zlc��)��P
�(y{�wm%.��;�@���w����3�:��x�닒�c�`u�z1�Gs^��5�/bY~XC�c!3ͯ*o_����:�����i��L���8s�xOR<x�uee�gz�)���L��(��M��X�p*!.����ey�\f��}x��x��߸R��_�*�WҏE��
<$�G>�!�c&�/w TB�z�Wt�;^�~�h�i�
�<�O\/���ב��s˞>��*��#PeS2�����~���0�{���$�_I|n�ש{N�������>�;O�:�?^�'� :~!��)n�;��ŗ��t�מ�CEf�j�[xg�J���ry����zo�r�2�]��F��[ �bN�!���@ŵ�Y��}�=�U�L����n�Ӵ�������_G����f��A�+^�A�m�����*;/�\Bs��i��Z�u�c�ӛ|�t��7�q;q�wƀ:�y\U���D�xw�r3|h�*�7���54."���<|�l�m��Ǻ<���/��٘�D���.���œbcMCdiu彶�;���0^���z���5:�A�٘m����S��%فe*y�V�u�H#vIr�K��lژ�vM�5���/p)q���2�Ai�&�@��X
��@��l,�ވ#y�G۲>���&ZWT�`s�늸��Rn!L����^�Q����W,r�D0��H�r��Q4���]��d�zO��W��`��������7�29�1藵�}_��~9+=A"�����]���7�ՙk�t$���}��M�u�{���=P29צe\a�l<��íF�٣xc�TĹ�\on�qW^�"�x��y~�i:�>} 9=��}t6�L�����_A��J}>���u�^���Z�j�\���}S�N��^�?}*k�Ǿo�������/w���~��XGFwW��fF+��x��!���L���d��>��x�}���/G���Q/��C顛�C�+;�
ܽ�~����k�:��c��̹��8N`0��XU�7�W2���\�]�
��ܽ������+Q���?˖/�T:���ߞ�ח(вR�3ƾ3�zed�eP��Pq��D�+�	ڏA�v-�ʯj[����뚧,5�u��u�C���%P�D�Ȗ!Ku4��\f��yuA�K�*���od��z���u�=���?����u���h?F��-�	(�Dc�f���� ��{��؝M!���j1}�"]D_;�z�p��6�p(1��c��Z����W�@���㰳��J�]K�z�Ө0p����M�_]1ZE*��*�A�\H�C�&��j96��I�sUY+ib6�v���K��9N�98݇Sr��*�V��%�(�ĢeG�Fl���٣��r#sq	��l0�u�t�K9�V)Un�0���\�3�ئm˘���'� Ss�a��|VŒ$M��d*��&Z))I�$�V�VfZ�{���2a��Z���>��Xѣ�����j�n�Hf�c�Z��%ҵ�9']��"�ء�S���o+x��<��c@ɬ�Z��Q��c�X�M��&fwai̥}]|e��K��Ǡ�;W<�g���uɴ���Ԗ\w��.�Xz���Xmi�7h&Z\�<�7I�wYef��Z��ɽw�\�ǹ<8�ɱk~]m�.�}���4�����y���w1���䖲���m߸��j�D�+F�	E��YAe�x��dr�NM
�u�zư��R}DN���mj4jLqT�u y�[z�쮷u�uf�Dϰ��YDe�zgV���;PIۥ��ҿ���,Զ6�ٌ�����%��<���fahh̓h��Y|zU���5E�Yt��x^Ym�Z2��L1��mpD���,�3�t�JE�i�Խ�BG���!V*�[}B���h����mZ�^`�HtY�-�|���{H��Sz��`�H�R�q�r��t�a�p�zI�Tv�6;��T�ЅV(}�����h	o�1Ak�[�<"v����Zき�Q[��ْ�s?o����}+����Ml��������]U��Be��e�>��;�V�a�s�K�IW�;5&ʝR�ciJ��"ǮҬ���w��]wWSư��#&�|)�qA�	q���B�i=%�Y���m^�-�C��S{ij^�P�򞖰��&�=���:U�x.�;�xp]�X�r�[ʐ�0�sz��Y�p.�g勮iL,٠��=�1 R��2A��r0P���y�Ģ��ou�ɺ��������t.1v�E��"��-�,�'��_�Tڄ=o�p�w�::
$��X���o��We]�U�il�����W���JS���u5�a�7h4!�r�E� ���;g�T�e&�M��V=�TZ�����Q�c35��5l���S�d�^Q�z�%X���U(�V+�̡\{��a8��Xһ���e�c�ݢ���NL�|G�cBv�]���/#�awQ��Jl������&��X!Clgp9��Xx�:^Tû�ӡX�oh.`F��r���6�㧴��%���fq\���f�0�+��2�i\*�3;k��˫��2�is�Ef<��|-�V(t �]{A���N��l��H��)aᔃ�e��2�X!`���5����be�l^�Ը�N�I����c�)Q��M
���N�T��I�˕��$r��V�B-:�E,�R��C�J��UP�A��q 5*���t�\SlĪ�YS1**�H�J�Y�+:qKIG.�N�{����w7[B���tH���Gtg��gb����(��u����.�yQd��D�,�99�NI��p
��v8u����`Y�X]�/<㓛���rJ�o"UEUQR���"��[�H*�QAS��.�_U�s�����:OTzS���G � BBt3�rT��(�®wA9^�¨
bBL�x�B�(O�������	y|(�<���N:�=�9B�8+�H���/����ޟ?�w�]�W}/f���u}N�X��Ւ��Ȇ�D�ͮ��0I�EƇn�\�PV����Y]S�aE4��c<�z�u"���T�ɋ������5�_q���i~�<m}~TݶǦ�z��1�%z;������=޾#w
F8	�������h���L���υk�h`�{����~��sYm/���M��N-��~�0�zNp@N���d�r�߁cVuhྞ�l{�m�Ӱy�t��EQ�)��w׺�>�2�SF���i�h蓊dD�H$���qE���if�/�����^�ɫ���'ּ���?���y�%�N�Wފ.g�P$�*	 �������)��@dU{��	��ՎŢ���j�M�u {�k�ކk ��޾���%S�?�,n�Í��jr�n�B�*��+��0�°�n�\?&��ߜ�&M�����:�������xt���v�7�5�ܬ�QOoX�
|�N��q]��\d�5o�WUa����M�����롙�����.m��z�pv��Y�=����d��'�{x�����Z����BU��������I��2_[�ї�w�{�-�뺞/Oe1��`�7=�b��9x��+=��oU��O)�~7��&�\I�Q�q<���l,�A�]���ߴ��΃��e#M���{�$^���:v��|(����ՆiiQl<��#s�w����i+����|�,�W��/m֜=d��bv��I��-N�R'[c��ྩ׹�m�-
G
�� z�Z��#nMln��7����K�Tyd[��eK�x�7Y?S�U���V4����Fv����r Ů���q�u���NQ�m�u�U%d��3��~��_��(ܺMm��-�VC�:��d&uM��
I��՗���*�f��1}��J�Ԁ�|��h���w�n�L���Ol��jb�HNn�q~��_�/��_�~�U�����5?u'�Ě��ex�<��d���
E���H]T�s������`�!��z#���o���c�"K�"�<ږ=y�<�M��׸<k7��΁"E����L�����(_Ο^;̅��=E�[�/^Fy>�7ܤ�S_������{�Ӕx� '�c`L��xS�<7h�VBY���^p����3�>�V��t�r;�Ԇ�~�7������p���A#L���ɮ�~�����m���]٧7O}٢����ϣ�sOq��v;������uD�j��2�5�C�}qԇ�S�r��{�®*V��q��h�w��7�<���g8��u�S�$zF��D5�X�&���z�لǙ����Ԉv�Z<˥�6�7m+�*���1�%�G4kc�G/�g8�̩y]=Ս�U~�R��#S�Y��U�J�F֥��,_^3ջ�$i�dV�{���-G��M��+��B�F���dJ	,�t��m�.(N���U���[Ẅ�d�$�|6�TON�B���Xj�^��!�ɫ�16�̗Ǡgt;5^�"Qי���y[Wu�1�(Y���)*(�(9f�W��=��#%���~z#W]Ȭ���P'�;z���[;|.g�΀v�9�+��e@��%F{�'0ø���qE���c�Fxvy�g.uH�����Z��->�}C�ߺ�t����ۅٞ�zx/~r�Ȧ3%��n|��D����A7�4�ڽפ�ǰ����U�Ks�8��U��}���VQ�D)�p�����+:�n>�S�iK�y��+��V��<�Da����;��N�����W���7��3�N�Q<f=��/�L��G�>�2��EK�����#h�p).���]&W���m�%�����V�����U>�͞�E�	9�V�F����yNC*�d���;�*3��bF�td���e�Vb�򢽕:�^"���eUD�D,z�R7S�7u!�ۙ���?X}��ʯ>W�;|Д�{�����i���H=��In���ʡ�l꺲#��̧#���wTܫu^dR���T���E	>�G;��1v�]H+�/���1�Ι�,�%�,r��Iy�/līA�� 9�EӽS�]N��S��sc��wq龐VF{xmQ�)9Fb9w����������nzG[��]w���1<���C�ѾyqW����ry����zoܨ���]��i�%�9 '$h�Q��y.s=x���T��������m����;H������^�3�i���x�fV�:��5}�2^�p�] l�ʁ�J��_,���뭳����s�w	���޸&r�3SV���/I�zƼ޿=Tt�uI�H ���ӝ���Y�C�m_=�O+<s��Z>������aT�~�n�SӤ�|6��+������t��L���������tZɫ�c��!����u�c�=�����>��t��g���7躁�~��p��F�����fQ|r�EJ!bG�tR\�r%m�jރG�nZ�n�MǟP=��a�����2�s���������=��<旻5�]�����W��=&`����OՕtܗUa_F>�:M���N���ێt}3zxR���'��'!��Go�#rƯ:B�kV���s��ma�/��1J�Ϣ�����K����
IC�&Uݽ��PʿF�W妴�99q28}S�8."��9x��Y�^��t����=7�������ܑb_d�lܭ�}ֶ�cp��	
鷈����6�Vy���M]�"�`��($��Ȥ��V�ٽCk(�ڏ�#��]%f�2�h&��]�ڶt�Z�-Yu�#ƹ�Ӂ��r�%�vqk7Ұ�l�٤k.�^e������-=�Nc���WB�
?{s"�u��J*�l/�|#���~@~�2���]v6G���~��>�җ��NR�/�l{�N����JZf�A��s�(��N@j$wOD��ꎏ,�M�����u
�UQ��wMe�p���8/:��w<��(��G�Z ��=�����HEe�vD��j[���E@h�mS�z����'�g��|�����:���gĻ���s�}���y��*kC������@�������T�\|�4%b���O����}ʡ�=^��o�<+��wɱw�mj���u|g@�(���S�v�����޶�G)8U@�S����kt��cW3�o���w�g(�n	ѐ6Al�Ger����Bν=����J�>�"�{+5�Y���-&㳮'M��\U˚,�"U@�%um���z�S�`N:Z5�p+|�<���i[���Op>N���:k�+"]WL�#$�l�5��J���Z�s޿y��{ܧ�ƫ��3K�&9=����ԁ�q� o{�k �}��n%׺f'���.�2���{5����Z��v�1P樛�[�d��+�@��.���J�3Fc9پ�M�#������lK�Bt������6↽d���_J����vǗ�w:�5���L�S�(�hY}������4���f�p�P�f�6�F�i]�6��)����'%=��9Ղ��}G>��w{�c��ܛ��_'�����&��X"c��������e�=�'g������>�U�K�Qo�ں�Lc螒�=��ȍ��|�}��r�{��t��{�+���(�G�5�����1�1�z02��k.�J{.'�� �'�0�����,�S����r�FSډ��}��̸3�F`��g��S��w�u9���R�2Vg�{r�tJ���G:���G)�ڧ9m`��̺��9�a��S"�U����@c�/E�������j�Z':V�*#ܕ�S��(�\1����н�m�oN@���>P�vF2o_�n{j�i�EtV�3Q��������N�����/�T{z��S�:ۜ�k6VV��$�����&P멖�%���3�8��_��J��<�]v�cԮ�j=�=�Tv��I��v�ڔ)#@�Z,_�*������C��uC���C�������	�>��v��ٽ�|l�y��o��{�w�ӔYaX8��z[2�\;�ׯׁ�tܹ��O�C5"le�u���+*��@����ں�~=^�~kk']��	A�0�F�z���%*�AX��zs��|_^4��o^mX޽Q1�M�k�����D�c���yFց΋�T�0UCy�df%���Z����끖7E©�0�A��&s'�/a�����edr��_��@�}}q�Ӕx� &d-�vWAw�ט9I�Y�Y�Ξ�G�Ӎi���]j��y��CI��u�ULVwU���9��}N��(�k}w�}w�+��;�w�;�ai��*:��l�>��\t�`7�zDW�: 9�oq=��a����Jq�==��n�u/N���,�P������Ȟ<O�/�:�+a�>�8�9G{�;�)�^N5^����=��7�$5cj�D���t�5y/F�Q�Wrb�}fO��s�����d�{���o�_�Ȩ�B���J��.c��	�-exe9�5y,bګ
��)E!Oc�F���t���A��wO uu���G���%W�2a��0�+�0����j	�y���\�J�Ď�{~��^��q�t����}5p�~mm�3�l+������G*{^��[�7#{�,�-=Gp�7��^^��T��q|��R�n���+(�S��̊/3�m��7�-aj���]�7�QH�o��+˕�zL�.%:�S�Tf�w��B��md�u_�3{"�rH�ѷ���ƶ�XE�;��le!KuQ��;�%�3��.B�Ooj��0%\�Mp�:�;��Y���&d�yq�,��:F&O��)�5�F�9�IScN���λ��-g碥 �0g�Ԥ1��H;uǩ6��kfP�쓇/��::OI��NG)Xb;�_%ָ�.S:��{�B���e\[��K��:�w���ח(��>%+�,z��,\EL�7NC*�49z c� K�2�}v��F99����G�E-���]!��漌\Gs˞>��@�#b�e#UO�q��/�����{�fu��W���=�;d��ԃ��:� �\�u�Iu��UeF7��sҡ��z�z��6��e�\Kw�}���v�O�I��|;A�-���E�������l+I'�#T����7FGa��w��}g8�9�t�*���F_�ul�΄�yx�T���}9��x=
�ā��]P(}(W���mh~�]m��t��3����l._R���u���^{N�W�p�,O�6C�H�����A��g�xnF�,�i+a���e<j^�Z۳�ř��*w���.sIQ�!���\K��6�Hj��b��u�-d�;��S���1�P�
��י|E��w"㛮'�9�� ��z�T}���P#�ߠ�*^�a�3B=�.f�U�=v�I��zX�y�bSU0�q�4jK��8Xv�tkp��0�BwK9�nx(�v����#�r07�ʽ[NU����p�.蔡Z��\,�-q�8�q�O�-v)ů3~��T]3z��t���|���$8K+(�_�z-�����n����Nc<z��	��6�@s��|��3C9T��zfU�6�7}��^���Tz���թ��������Z#�}�ߋ(��]w�H%Ǻ��ꑜ���U,�	�"�F0��^\�*tu��
��R'���+�E�������o���l��5R�`I)Vw����n{ܗ��p����ắ����I~�,�M[8%>_��ΦDg�z8z"]>�O�zǌ_weܪbbG��2�C���n*���-�=h��0��c+�Xo�r+������]G���Ԩ��eW�:�������})�]xf�|�)�yr�%-3Ơ��;��G0F\^�]�MS�\߻�f�}���*��X�wMd_W~��C��Z�sʇR �r���b�^z=f��W8�oL����L?��Gl�=���\u���h=ļ�����opd����I}(	�ꎒ{�2*z�>�~�K�r����v���WC�b���p���W��E�i���Ap:�(�y�����]��N���s����x��*�:�Ƴ��=�۹�X%h��چU�u�n� 	�k\+$�mY2�%�1���z�[�Ѻ[����2�K�]�V���fʶ�Tx�c2ۨ(��Y�F�X p�6�@�R�b�%��Se
r��}jH��]�	*f@[g/1��O�|���m�5�yu�����r����0d
;+�׾���z8^ҵi�ט��;�&��,��X�9����Դ�wT;�}qW.h�h�P�4I][F�������vz�v��7��PF/n���tb^#��w;c�=H��q�M���@鮸�h�DS"�@���2f�Kh=umGl��ک�tz(�9WP�Z��oɫ�7�ԁ���'�?�z���f&���s�������7��b�wk]O3�o�/�z�����9|L���7����z{�?p���m/K>#�ί������wR�ว�¯%�[~�z��,}�ub� R\=v�u�6o�]ى)����t2㺆����za�X�S�pG��\?:��X�V�*D����#���9�><�����ڨk��<gWm��uL�F�'2��*�a�W���8���m��Q�
��ɝV��r �k��D���}뷧��hv��ೳ.�{�8Ne1�KR�+֓����^4�j�%�Y|��QXO\� ��DӼGD��Ow��綇k�IJ�ġ�G��q3�(yؔ�֟�;���SU�)9)��Fw7�*^̫�,#�X�H>͂Ҧj
# 4��6�;�Ǭun��ʮ"Ҥ��̾��L��5k6.	�������V��*l��{i�L[��o��3%��R7���R�I��ym���H鮊�[��y�7��*\�i1��|c7v��xi��l��1�Re��J�o*�j�S��<�+6!���б9����lǕ�$˲-�4v��A`Y���p�[����e7Ҋ�옕`{�Cwf�&J+.�%4�C����U�wv��t��|���÷��["�����U�&2ᗁ���>[V�ljd,z��[\�݄�N�z@���d��r��oP���U�=�]Z��ܣ]��Te�5o%��T��WW.��a���j��g��[�q�& v�0�W� �#���ry=zf�*���4�լt�����<��m���~��?eЀ���ϝK��B��;�~�n{S��9
�SEu��(f��fs+R+���1�Guഐ�������ob�7���n�zx1)�۵��,�il.��ݼ@��Z���:�]�*$�.�]�N{�y���Z�����.��R�B�m�͆%f���]�.��{*z�h�l��r�:#�κ҂��cC�# Sc:"-�{�k���'t$����d�O��E�zE�1^�y1]y����Oz���#��_:��������^P�F���'�J���������JE�+d���S���OF]�G&]��'fQ�+�g�Tx�9r�y�z8�b���B���/7O-�s�%ҙ��l-|���V��}����Yڎ����`	);(�7mu�K�T-"�2lV^�2�����%��0��dS�R�`*��4㓍gu:p�c�⍊l�X0����xWd�WLnws(-�h)+}yv��=㓲��������aK�w7;;ȉ��h��^SݑÆ�pӠd�̔x��]�]XP���I����eŐ��E���&u��m��m�:�Z:�B��W\Ŏ&*%��L��S�X�2%]B�pSY9��)r�������-Yo;E���N� E�^v��[5a�eJ�"�ָ(C�˽�ը��`.�F|)�.��]y˖�A�+,Q������k�C��\���f��K���Hd`�C��$C�sQ]]5�4�EY:�&v�8��շ�X�iqU0�����Vͽ�b�Țz]�{1��jv=��8���L��;��L>iQU�q-fʌ}� h��1�>�����oUC!ƵZ�\���SZ��)E���PN����P�m*�;8�5��u�� h�u�s7)<�7ygv-y�^�:,���3��"�z�7wA4��zwM>�k)�Y�]s���լ�-�q|�c�/2��mk���������^�7��_��gա-p:��A��w�I���V�u��u"I�\V���G����\;!�U��ή����WĐ(|\���Ȩ�^�"���#��s���7�;�N�ys��Q��/�9�*�79W*�֣���1㞅I��*���z���s�i�����1�"��r��s���K�E\��E\�"�2�U_�y�G�r�1���V��rI����[���*�.z�b�EQ�x�#$dq��C�&��N@�U\��i|�e�5<�\�wr&\�r�C�r�� �B�"�����Nq"����/�!]� ��r���DTEE(��T�@���|e�ET]�GX�E<�*y6,*.Q
�VQW5
�U2��K�\��dAY���"��\�9�$PC�TJ-%!x�Ç(�""�UQsVDTDG=i#�9���$�W��=�Ȣ��<��(2���ul*._<;Ώ�x��Wu�v%UQ�]�'! �ź�Az��(�^�/$�(��J'5nw3�)\+�-ω��B����&U䲞$(�:&�.z�#���<�+�'��4	� �F�[.֌O�Ϣ�zdŉ��x��p�'E��(x$P<-n�$�[W�C�Bw��P�v'�k�F;�D���c<�o�������C&ø�ʤn(�9=_х�	:\z��㸿}֮3}��sqR�/z�<�J�U)�J}$���	�qS<�.�������~yE������:Hb�f2M��~��ޅ�=
�f��t�3��jH(��X��H_�S�ϡ�h:���<������4����X3�{���>t��:o�z��8���F�É�ǣ��P] D��6;۠��׾��P��j���̬�G
��R��Zr���l	��@Of�t|o�[�짺�]Y��1�j#���\:k�z�r;�wRMǻ����b����� �/'˵�Ǐ���g#��K����W��R��54T;�o����=ǎO�߻����4YyNS�S�G�p��g�MU'zn �6`wRT�83��P�EC�m_I�<���g8���T�WO�Nd�=���4�=�RmL�Ս���Bx�_d�5��CMUI�V���ձ��Z�*�31����%a���ꌊޡd
���+��9A�1塞��x׋���?\��v��Q&ޥܓ��M�����@�v)x�����1��F�~O�2י�Cf9���frv���N�{�;�Z�5'ph<�)��+�x2�z}C.LNfp#
]4T���,�9{�(Q�2Ven�uу��v����f�S��`�w<�f_1aj���}C�{� s~]�7�j��~��W����{?cB,ܔ)㟢y��}���O�����	Uv�F>��o�V:v_��3�=�'+�|9\�dW��>�{گan^Z�gE˟a��O�FƢ�����������ʫ�/v�>����ܔ���XU%��/�_b�P�9f�!Y,dc�\F���\s<��SqfW��������.��������T��zq�.�,�������y��I��NG)�9,c�K�q��13��8Gc�o�׸��r�}{q��^3�k˔}�Y�)���,\T�#qNC*�d��4vh���I�yFu�U�״���b��O����Hr��1q��現��)�U����~��u�K��/oן��%����h[��^�w�k���Gh���;m���}�R�}E��e]���3�xv�[�G�V�W�}F^��Ϣ�\Uķ}���O9�v�M�����{L�,����y��(Ճ�����t	��l�!��F�u�[�iC��+NDwI®=�dg�;�j��}����>�ЄƎ�ԁr�|���˲Lm����d��VF��&� ��^܍�SZv->[[�]�2�=ҀkY�M�]ױ��]���H:�BOu�ܶ�k�
� Ks��au���ԧ*�c<4bp��:�Gv��(��|����]p�sc^ť{�Tk�d<��]L���n�T��
�/M|�kC�:�lǺso�S�\w�e�v�p���֍t���Ps��١q.��j���Hr��s�s��U�Ͳd��qV��]�g��ͯx�Z�Ϡ����=�}}qE��(��;f+�{]F��-d�O�"�[N��RZ1�>�/�^q�b�!��6�������*G�G?_I�FG#g}Q����/�I�^	��J�y�#0��0�yoe��ɺ�>} t���4����_!��nfWo�F�8����W!�=�Sஶ�����K�_}y~�~K���1��o�u�w���mS���E��8�[m�V�x��wBsıqΩ�#�q�:��u�+i��T�a�7�[��^���<g�Wcמ��Y8Яv���q��8�|�㓄� d�wS�8/�S����S�=��²s�;O��S�ּ���tNm�>}43^׸��;s.t��'2��?P�E����dP�51�<�^�Rc;
�v����W���%5ށ��>���^���)�yr��ωJ�ò�+]{���4<�����vX�}��P��T�+�q�Q��9��W���\�9�u��7e��a��զ��K��.9ɛ��0t�:�K����*�;ݲ�4��4b�y��ϯ*ٺ����8�u�J���u�4Y����h�
�
�^S��7s�s���H��A�=@R�K�k"��s�8ju�B���^�D�}�v"�GSek�Z�/���'$���1���=�H�.7������>��<{;jl���\wH<�}ڮ�W��a^�7������'k�`%P�[����ϟ����}Ǒ<^�'��(5����K6�V��,{�v{�&����c�+�w],F��n��.�S�v������}���n�';��w��Rp���u���f��xۂ`��d
���5��x���Xo@q���^�Їe%l{�6�nwR�n=�pt�u�\UĹ���" 5B@�0WVѹ��b�u$6��yR^�x���Y��&��#�����GOR'�g�� ޫ�E3�9�-{��K������yo��W�*N�'!���B��j�M�u {�k��f�
�޾[��D�����x���!��`��f:�Λ��ب���WR���/F�e�M�I_y��d�wu��"V�z�,M�=w>����Wu������.|nx+����+��®2^�[~�~�]w�C:W�]��,#�@�x�Գ+��S��`AT0����N��=��?��7z��*`��ʼ����b�6ᵒ1�5�h���a�٥�
��p�Y�M�m���G�A���/U�Wy͌W�p�������蓶}����vݩ��V1,�o�TƔ}�!���L�b\G;���Cٽ<J��j�X�Oa�,�>̔:��_��{$T�<����h�n��=��oO�:k��}�qB���t����2�!���3�i���8�3w��UŖ�����j�v��� z�i�%�^���]�>�4;T����{�C��s��\�d,��v/6�D���ﷅ�����U2�*�S Ty5d\J�\G�"]pƧ#�+B�=�;\�J1c��q�:[�ݾC�>M��*�]:�n������
��r��8�����G��2�w��������~���Y%Z�J%��3��<�2�����q~��P)�_���NGJ�V6����l_�쭦�h��µ$Ft	�y/�H\UO'.̇^�F]��w�ڡ䭪�j����AS{d���om�7�zd�Sp��#]����[/kL�q5��56���g4�B̽�
���{��2�9Q¯�u p���������3��їT������W)���õ�M,{qV�!�s���wRM���#z����==�Ď]0-|��F�ڠFF&x�8S�NL;Vݽ���A}i�g
Ux�唗1�
@���]�< :��k9փݱj��x�rc}��r�V]��uK�]��t~brF�܊T�܌�V��ƞ�{;V�G�6ĸeqC@ɘ�!�˺v$V��&2V.��w�c�=�#L�ʁ@��M,�P�Ϻg4���k���!�� w��v=q��ݓ:���޿��t_�RyH o�u!WR���@/�D,�P�W�o���O���*�A|��n���S=:M���*9ղE�K�t���\���C+�a���bO�/Ô��ȟ{
�dP�_�����'����u�� Ts�t��s��;������S��Sb^�W���VϢ^�����]�!��H_y������˽��ތ��Ī�L=��a���o���ŗ�*�6�Y��裘V�k�
��_|�Wi������U����e�]����L�Z��z��o�>������{��F�W��!�>>����=*��>����*��۾�3!p>���Q�������t�8r��~5Nq^��p�A��\�;��=����G�l{*��uGrn�}w�|׆t?s��3ڳ��&��^�Z:|��pJ��?r�9,w �+B�����T^H�]-{,0:r�=�����1v��G�Y�)\c� Ζ$�G)�e)��a_��<+o1��Z��L�e�����1�Ad3P�z///[��� �̓D����#��X��/(6'sm���KWr=��*�U�aQe�g:ŕt�)j�%����9��*=���E��KW��q�v�u�=Kv�E̶k�΄�&���wu%��+�+�;��J;��^��C�3h��w<��貉*��#_T��"<w����^߹��Xz*���Gz�0�7��;A�>q�Gm����>u�A�O��l�Kt�����v:6'g�ug7Ώ@�=���3�d�~yqW-�a������TF\>���M�UW�M+���T�^�=�|�����]P(t�o�2�.�*�qZ{��ݮ٪;$tk��b�V�bW3�_u����P,ۂu2�n�T��
�>�y͗���}�_��E�{I_3��C�M�t����9��m�\���4.%�nI\	d�hK;���<��[��׺�U尮o�fW���!�t��q����
}}qW.k�ڙ!���b��h� u�E�kI�����no���o�U�Ŧ��[n����7��� �.�s��:�7��%H	��7�қ�>s��)�ʎ·�\SR_�}@t�W���|����cS�~��-an�I�dDo�r��W�E��������Ӱ������%�z}���q��;9ٞ��\�	ǌ���n���#)ߌJ�s��_�_���԰�^�[��-���X�{n�KZJ
��j��#9�E�-�$&;�f:͢V�N�[r�Gυk�٣�6�t3:JB�-��m�s��vz�j�W�u�u�eQj+��v��^Wg7�Q��x�i��N����1��ͣ��,��d�w��/	Áq߯/n�Mv��PTsۊ���~��n9���[�����9ư��rr�g�T2p;����}�����PdL\��˞�վ�q��W/@/�̨}43^��e��2�K�2�n�g�#�,�;ɫ��M���o�w^�r�p�� ��hr��@���K���ӡ�k˔}�����~ �لu������%�/�!��]�L�El���U�]P���Ⱦ���]��zzо�!/,�K��b��C�W�X��K$V��.���E2�e����>�ǳ��p�OS�Q��6m���޲+�o]ש�ͤ`z�М�j��-�g�=I�C�К�+�>�'�ӑn��/|�=yѕ��c[W��^�C΃��=��u�:�3�L(�nb�S�v�¹A˞��]O*𾜉�&�`��u[G�>:��u�ˎ��a��Q�p���fl�PvW)��g���*[{s�ٝ��.�+C����Nm��߻��뾸���4Y��D�� h�}�r����7}(���9"4%F��V.�
|��n;EJЎ@m#e�f��Xԝه��=���:��c� ����:˰�t������0h��м�H��eb�6��gT+?�=PL��-l�~];9�YF�C6��q�޽�ŠT���f���������ù��T�|G������O{���m�V�q�}諗U�3�Z��,�]�n����<�ݕ$?=E��>:Иz����ҁ�����t�q�W<�=���~�8���aY���`Jl�د���UԾ9F��[��)�Ty��d�~@�5&t�#�
��w���c��\.��*��"��6|:�ꕇ���/B���=\�¬}�FT'%1�װ��6%��t���C/z����&��c���}1�1�z00��}U�D���
��9K���~夫�O=����Wo�я�oO�����m�
��z�=ޱ�,��p��Vo�q��7�yg�i�>�ր�{�����A�:���ܦ�j��[X.#;2�g�s��nuozeu�SVn�ه{U��a��ng~@��Q�Ցr���u������m���ن�����ލ�i��7�N���K��7���g�x:�����[��3�P�Q�}���	�T*�i)^��W�z�$�H�V��
�·qS<�/�r��x��ިl�^.\P�q�j�ط��=�+,��j��d%�ovi}`]u"3�¯�Qt��R�L~^���_���:�J��}�7��.n���#�O�y-!OU٤��0?8ed/L4���U�ov<bA� Ɔ�t���=Y{u�+��k6/R��.�ssi{?;��=�ez:��&f���+��RAU�~�bJ�2*���x�פw8�; �n��u��ݽ�u1���<v�����]{�v�IgYD���#�Z��w4���Ǹ��Vz*g���B�>��9�s+>�G
�J�a���{�9G��"r�{�f9�(�����K��8��+��\UA�ӿ,�tאg�������n=�Dm�]�=��5߮���W����j3�5=�7����'0 <<��þ�0�}m�t�i�9ӵ���h���X��=��_<eM���U{�\OU)�$����������*j�K���鱲�]�+s3�Jt���9��W�u`�>��Aw<�rD{�p?���,J�as��!�Q3��w?M�p�����+�Uܘ�����>�����2*7�Y����+�.c������S�s�r���뭷��5�ƺ:pe|��Ç�S��~}C�{� saw���G�Dl�*0���o�.�ngE���u#�՘n���荮*��l{䪻O��3{��NϾ}46�fz���k@˒kG�
�[��
{�We�*b	Ӑ���6e1ں}&ؙ�72J���d�gt��r".҃��^�iǟK�L��u�����\; �i���T<���50���h�,�}Xz����e�k�\��66^�S6��b��)��GJ��� �夫�L�r��Jq#Bϔ(�`'c����V^VR�ord��c�r���':��|-�f�̻����,YV`r����W[�e�Y� �c��r)\��Lo��L}�`�+��>O���DC�=B�Z�,�������Yo_�Z���b�MD�X�p��wJ��̆����j�3ƫ����(�����D�+Og*v*�w�,�tT3��OO_�q�i�Z�����7�ֹ$O�-j�nw��K�_%4��P�b+j�Q=;(Wt�;�ɑZ|��8�R��Wy/R7%[YJ���yR�s�(��c�ߗɚz����~�W�Dtk-�Z]P��i8����6�
]�}|Zn
����	�:���/�y7�� z�쀟b�+��aކ�������@�� �vG��K���N��c���-<��ݺ;׀J���X��� ��7�pB-����ys���8�D��j� 	ݔB���#xh���A��6�{��]{wB���*s�apv�S!H�TҨ���Cd��	ujK�viIe�B�Fr�����.���J�S�X�tjY]�S�4nulG����4��i��Z��5��w-��k���.����w�SV�>�n���)&����эYjQ��͵z�9͎N�%%ˬTż��/���N⛉b{�u��s&����r�<��	�+q�{r�2�AL��nkr�=�����G�I��Ǝ�wWA˧5��n��������kr�VT�S뜴��,��BD��Mg��sz�<��"���Ѵ2�9J�c^�Zg!U+���.����;�GMY�2H ���W���I��}��˾�cLW�),�,g��Y���2M�hܕ`V7�H6��}��	�n��e
t��K#�[�c ��l`j@	Y]O-5kD��κ��P޸?�ˡ2=���v���>Ô2X�Z�T��0�x �h��\��P��QK��3�)��:O�u�b[r�a:,�y��޿�E�yq7W1��j7�%��(u�d�e��s�o(��B2=u)1�C�������6���,i���IA�4R�C�]qHy�V�s�l�i���-]�%�\Z���QŲ����kA����Y�i�f�v�P�Ij���۸�P|�U�ԫj�K-JU���Gn����tj�)$ܭ1.)���l��_n����'<�V)�a�|��{�2�$�4�f�˝G�����P�2�������Ƕ��ٝw�A��ͤ!���[����:jD�@A��'�M��MI9��FL$�*�$�5q��nY���a�ٍ݋Z.�i��H]��	���}!�wnf�.�^�u�N�r�s���=iS�D�K��$
�*�wO�t��B��n�S�@�\��W
2-ֲ��Y��	ZG�Ngd�E"e(��"�!��"=�B�U:��^�<���T�e\�T��nǻ@�ra����A&���p�䐝yk(�zӟ.^�s2����)ՑEqD��U(-P�q^t��E�]�����.�Ĳ"**�+�Ȣ"��i���s�*/���E>"�z�-��E�Y�<�yۑQK(#�|d��Y�|aN���$Qz#r
=�wJNr���r���띸Q�
<��L�U���TW"��x�9VBV�d8RH<e�dp�Y%���(��$PT�!�Ȃ�ȬZ�9ܣ��B�>G�-���A����:��y�t��:�Q��v�Z�uJ�1B���� G������P:2��5i�;&�˱��);=��� �o��7�Ƶo#t{	�q����`���u��}��R���8��tO���K�-/z�h�ܬ�8�,�Ti��ꛙ�x�G3�Z��D�����]�Ol�/�z���o�ݽ��ב]��3���N��=�^����Y�`� {U�~��^��׳���x\�v_T{�F/T�d��A�=@Ζ/��y�NJ�͌��s�wu��{�0��M�W R�z�W���W��V��6����</�@)bȽ�����_���rAy��g��T�}��{����{�{��#��1�\��N#O���ᐢp��c�{:6�%#�I���l	��Pd�����\D�}��<�v�MǹQIRr���?g�	�c�~���g	뎐験�Cs�-�<9}�n��Y>Ⱙ�6��۾���||k���#.:����uP<\ �$��@�_J�^���Z�������k�	�Ie��2/%#ވ�������wƁs%�U$5b@��Ў7��z(|����Ge���z��p��T[���.�i�W�׭��+=@p��|��Y�m�' 2}���Uc�ȧq�f�J��8g��j3(,~���S���l�V�͙��v��N���jݵ\l�e�[�܆��u��IrK�J-�;�O�ѻ.G:~��t u�W��t��q��ê=�}}qE��8�Hj�NىnJ����y��݌B�޵U���̚��l-VC���۞'��g���7C����~���y���;���
�,�	N#��g��ihݜ���4ѕB�����\��>�:{����̏G�_�+ ���u��/�vuzfz�7 5A����:<��A�7��5���X|�@rn���dwM����`��<\�o�M�T��}G�7l�(�Op2p9���EK�p�FƢ������n��S�U�익CyV�c�TV��ڮ�߯p�G�埋�u^?�JK�s���5l����9u�3���,r�r���z@�k�z%��@/�̾2=����1��T��g	̸3�'�adc^\��I�J�tNF5�m���^�\�,�@��\���})�ן4��Jz��T"ڋ��FfD����{3�;��Ѻz �T;�������d��0�c��4難?u��z�)B���V���\��:j$�j���3��p/&XN�w��;d���}0����/,��O�Y��5����.2��@�{�u"�
磾`�ݷ]��(�v+⅕�a��a��/�kX&�]@h+M19��E+�D�X�v�$���((q��iיّ>u.��s���wntE"�Cթ���6��m�B.�x���ɠ3���h{ՙ��𦅟]hx�h�$�}3�H�P��nbOJg_���,W�{���׊7ۮ5T{,�۱oNx�����8ڿ*n��|{�,���3�L(������ue㯈�j�/�2<�:�=��]��0z9�[G9I®=�ps���{�(��nl�$!au��*�k׏ifw�n�ޫ��F�c�=�����9��r#���q�냦���늸�4Y����(l{rǇGB��pn�L�*M-�,q}^�qEiY�1ʡf��.�lz:z�=��q;��@�����5�ޘ�>=�7��OZ������g��W�@1����Qzr�2��Z�C������@�	�w�7���r�������}=^S0�<�b͂�pVEK�n0�5��ɻ�=��2f��� l��y��cY;ׄ��{��@ꡗʏ��6:\�<5�������/꽎�5� tWw"��v�e���wzcD��w��{zG��_i�UL5c+���86�[�j^�^&�s_輳����Y*��v��=��oO�����ݷ*;��}��̿���Ƽ�������]G]G6Ix\��@���S�>���i� �{"�m=��s���T++:;�E�������H;��P6��]mN�j�6�'y�ql]<�+t��Ճ�3sv�����?���q_̣)��t+x�Xm��S�b]:�8(������yW ��W��.��s���d<��[X.3�.�+���x�]q�9���0�h�W^��qG��,��Ցq+�q�]pƥ�����Zh�޽���k��C�;�$�\��2�{ƌ�B���n"�������0��t��bbHup��{޻y�g�
�����ϳ�_k�����$�S,*�3��L�r��x���ז�L{����j��yG
g����Du��^��y�1��,�ԐU|g@�ȱ芕H_Uy>aP��Vl��y�]�g��A��k��:��v����v����m2N+�$k�I�����gzm�jG�;����L��������̮R|u{���uG(Ӕx���O�W�F�&�����@T-�^�0���;n)�V�s���}�Hi>�2�zv�W��V���npN�t����g�ί 9�F���P <<��¢h�w�[g�3�{��W
���׻~�}����D,w�tͳY�b�Ijn	a��^�zpg�|Vh�oM�SڍL},M��.��J��%�� |HX�%[�9V-#��vҁW�M%��Z�J���c#C��Չ����Q�h�[����lT�1ž�����qW+:띫�vi�*�IP����dڳ��»��#)l�4��y;S���[d�b���kmk��]���A�������Mq#%��M��Hj6hw�ҰӞ|����N<��˕���b�!_5w&}FJ}={�Q�Q�,�\�>�[3�7�CtOG��]TG��u�4�WZ��l���ض���Dj���P�� ��V��ʁQ�ĥ�w3o��lt��5[���مR��q{o��c}y~���*1�3q�;/����UGL��]�Q�z=���t�r��h��ދ�#ZN�°��ems�B�������M
���������nj��W�6U���C]����?c��n�t�%���W����p+\�����OrkP�^����'b)��3Ts�F�s�~�p�>�Z:5���ܳiͭ�U%�3h)���H�%p*9;\`z%�ez�\f�!��1v��G�gĥpe��r4��ד�	��)����q-�V{�z�4��63�»���t�/9�#���IBz��t�����.[мAsc���fd��a��0�{��=�=�Dv��c��שV�u�	�w��-j�ׇ�+���法��4�p���_���tx5T�@5p�r��Mi2����ǽ9:L�ޭ*_s�g8��/�*�V�����%�Z֖Kdy3e�t�����͖��;�8$��Ά��:j�GC���S01���rKU��f쬨�[Vf�j}NW�<�<�mg����(�fIAqv�'�Wx�9<�}�m��5	�f=Y�b�r2��X=����ף��p��r NH�. )�0:R7d.7}�p������.�y�W@ߗ�sx�^�i�\{��ˎ��{���E���x���8��#"&;��'������J�1��;�;�p���\���4.]Qf����f�y�ח;���Wb�!=t_@1��{,���w��<��|����_>����s]&��%�ϩ�y\FZioP���Q���ɫ��c��"3V�ȸm������f� �޸�i�Z�{ׄ���"�b��y��+�nZc�8�x����ަ5)�6�=�u�y{�J�\ǹ߷�Y��+��\
�u�U�C��6���ZN��M�X�j[���ao]�E�zs�<_������\����;|�\r�"*�<�$�m���T�����e��j�e�5��Fs<���ќ���}�_mW
^��z+�O�׊���?�����M��ݵ���nb��z�Q������M��KX�-�c:^~2Ee������{�8�
��z�F�8{�;�}�s��F�;-��������sٯ*�6��%>�Ӽ��9uҔi�XP�#/PA��S
W����AL� �-=�w+XwJS5׾��RR=��~�jt��^�=���s��_Ǖ�0���T=qav�uqC�+���;'�G�-j�hul֛�������X�.W.�K��M�a؇�H\v��GM[?db�45�eg�<���������m���T8�1�n@$�wM?���s��v�k�xs��?�,˺���غ��o|�a��P�ED���ug��Q���p~����ǽ~��.�};��1-�t/\��{\��O�Xv��	�A���������j>�zhJ�t(A��I�<�T���YU������ԔX���.+��=^�ލ3��p�	ѝB����mu��a�T���V楝�=�^ׅ_�J���oz�9�)8UǺ�z�]�������nc���ttq�U9;�>�Y�=w���d��y�^��;�Z�=s���N�*=�pt�T���sE��oӐ^d`��n�#���{)��=���a�,���|�}�;ǽ�pq7��wjk���*gȋ�;�>�lך}�	oM��u�o����L>54T;�m_I��Dܲ�uמ�����;��c�򺾔��Pvs�wYC�U����\�.�q�e����ȫ�~^����O8��G+�s���W��i:%H�i#��R�I�ޕ8�e�ww��i�@��+��^�N������I��r���t����>�y�5�����7�0��N���^�x��~�>�)y��W$t�(E����ʬ>��z��jS"�Cu��^ȩ�w+�y'�y-&�;��އ1���"�9ׇJ�G�ѳ�_I�	]<+FC��Ϫ$�=ң)b^��5~�\�P���]'����#ϕ24q+�=���f7������5�'X����Y��/O�2x*�˿J�}�G��:��F���\�����v��	O�X�U�W|%ጿ�Դ��Jp�W*3ܯ���^���oO����}ە�Y�׫�k7{���^�ŴǷ:���Ӂ�_�c���h��+��[!;�/l��N��5:����Y�w��_��[m��xg1���ω�s�P˙~4gj�uP!��9��n b�޴�r}��}#3�<���յ���{q����.;]d�=B(���T�)����n���thy��h���K3�%��3��'��m��z:�;o�5zo��2ϭI`�,*��DųB+޿W�S��-�z:*��g�w��_�z�x{�up��<q|��v� ��c�O�(+Y�U{6�h��^M&�(k`o7%c���s���jj���d�3j�j��)�Z�-:������V������{<�my�9����/t ��w3r]Ma� �b����;��!VY5��5��t��t�0],��w(�H,R��{��c`�e�3�ԙ|�%��+`����`~�i�[��jP]�~~�A����s��h�W�@�}}q�2*=�o�7�����5�w�D�3`�P\�+�0��,��My}<�.�Ev����u���^��W2Ⱦ���_:���d �J`z\y���K6��7�ٛ�}�ٛ
򍔽��Һ�v#"��{ަ�oL߉�h��S( �:'b�a��������cށ]ٚ�(t.���D��t�q/�@��)�_���t�S$54=.w�qѧD�ic�U{}z��Fz#�4��D;��ܘm�����s��(�����������ʝ�D]�Y�/M�_\��T,'_�q߃�]w"�Ϩt��t�k�+�z`?)ݛ�!����$�|Ǻ��;R�y��T޷zYF��~��?~��/�uX�����#QU0������W�{ӽk����Ew�x�P�F�eC���¾��,�������#�Y�ZMu�ݸ�����;�ǣz�
^{��o���z>S˟��F?SM��R/�,�g�����',W�	V'�?����X��A���k�1���㏮RV����z8�}D�����jߔ�,,xĬ{;2�ێ����H����	�
�.d�Zn��@v(e�Y���B�Bc�.ӗ�%3�y���*Uv��LT�\�S�>��%�����vk��}X�}1��K�?j�KE�#�'�TC��ѯ��:�_t�>yQ|��Uׯ�1�<zt
�W�'K�=�t��z�6��V�K7�]F��Xnٔ=�x��ٿx��n��$�Vc�'��V���[�_	�u>/�P�P漌_sˑG����>�N�qZI/�Ţ���Z7E���A�����q�d�����ȝ�q�~��L����ˎ�7^��|�\�)� !���w�W$�Q*x..���7}���O9��z���Nn�&���VU�G���.;�|;�g	w@	�I�$)�0:R7FB�{}��Fa�>����F�y���;����9�®=�de�ճwN��pB.���6Cu��:&}��)��Wvw�7ۍ�m��-�;���ُGNm��t���o]�.��h��5�i�7�*}'<����\�����JsN@���e��upa���ǧ8�}Q���늹s\'�~��H��>��e�:"`�VѺ+rj�ɇ��D{5�	*d�7�Q�?}G��}o�c�6��1�co���6�1�cm�1�co��1�m��c��c�����1���1�co�c�6��c�|�1�m�c����1�m���1���1���c�6��c��c�����co�����6���
�2��_>S�� ���9�>�J��x�UR���HH��RUTQ"B���H�HU)I(E)J*���T$��@�(	(�U)TQ���E��R(M4���P�5v%DI*$��EP�(�(��B*��WZ*U:����(�����-eH��Mm�ʒTT���������PUR�D�$QR@�*)$�"JU!U��PID�
J(T�%**QUB�E%* M���T/l   Zxzj�d�;���59V;1�St�lWs��UZɱuL�uEnU;�.���F;m��V�V�UXݝU[8R��D�*��  v'��[k�d�����㵪�O7���EQEQ`X ��(��,�(�� ��;���(��(����(�� (�� I 9;�(���RV��J[e\   -{�TwJ3F�]��s0.��kHì
��M�uEi�N� )ҷ#[[IN:��Ym��rhݱ[�ET�RED�"�R�   k��Ԣ���wrԪ;:�a5u�ZVW�����[�ͮiن�&�[�U[]ݫ��ݗf�J��Ԯ�e��sE��N�Y��l��R���R�UR��)U�   6;ջuví.�s����)[��:�k�R��Ỷ;�:k1ʮkmg[����N��8�«k2�t[�Mi��wl�swl��w]gm�b��һ]U�R
�U$��Cx   c��Yf�m���ڧ[mv��w��v;t�U���a&�[��Bڥvk���[Swuv�朻��b�v�rUj���&�Z���⻻,v��ݔ*
lev�UBT�T)�  z�hۺ듎�uKd����Ҵg�%E+��T�i�j�'t\�Mݦ՝n�Lݻj�����n�B�8��UݥK�5�n�[mmt�9$��QQ%f��K`��  y�lDU�,Қ�T��m7(�:���k��E�R�RZ�T�n�r��]�ε��i���s�]����F�WgN���ܨ����N�3��J�]�EU$D(�TJU^  wlS�64ٳ�wK:��ws�StJ��[�]�wm�b�:s�v���һ����j�\h�V��wwu�����R��%܅u��kkwR�֋n�iHH
���	lʒ*^  j�yѷv�f��:�u�[k�5�u�Qwvh��wp9���:d�]��k�U*[3�]ۦ��m������m�Wt[�U
�v���T)���*��db41��$���F�=2b@�@ �J�   S�i1����   $�E1�Q! bN�`�ȆF$3��M^�V3�F/Cr
��8,X��冭b�<�E�D{ޏD{���{�	%$�BC��$��BH@�XB�$�BC���?g;���2�҆}���e�&&QY�YN�2�c��(���X�H�#C�]�f�)F�2UHT�r´���qԶ��kf�OB�󩲢���52^����[��ŵl�"h7F��Z�q���Ù�ESN���b܋0�,[`h0�t0�F�fQ�B�y[�-�w�Xō<�nG�t�^ܼ2CH���"F;r�4֜��QFM5�:*0n�D1�f*h5�<3,�Pm�)���6�\����>�:*��D�˷�gR<�(U)��yB���VEMD-j�R������!�5v�̈Q�\�ş�JM�:(�2��b��.���,X�!���y;x�� ����.������&`�H]k�f�R��.3�3)��V^V�Y�d�����(J$��4�*�6a�1�4 �yV akI*����v�ݬ:);�ha�$�З�q��nJX�v/F�͓C��^����IM2�V�x m��)������k�����.�mG���iU����D,|umb�VҲ��!�f�
x�&�n�4Vk���hʷ������2�����r�e��X]�)��Z{��l@�J��$�h�x�%���!�@�4��3�Q���5��n�[x����=#�yp��ZeFY�j��p��[y�H�n�p1.Ƅ�Į������ڐ��[K`6���w/7)8� @*��Af	�^ǋ���
�m��dw�]�bk0$����]��c�)��lC�fA��%Ѥ���u��E�2�-+���$�����lä
F��/K�Xb������ei��}1ص�p��c �M���mF7�6�2Kffle�*LݬՔ�k]dya ��h�4���3-��:Qi�����u�GE���G�L��B�Y�+8�1�tP�� ۷�����6:z[[�6�aD��Vꖨ����ף
�k@Y�cM]ߕ詆��WQ\|9�M!�r��/Y�J����*`xU'��e�x76dA�Wx`�gi)����n�6VG�Fa�E�d	��v�$�̫��G��X+̫5�f�ȭV֜n�CKo ��܉ïD��9):F��?�`��l�YE�n
�wS����ò#ʓk�q�4���&�bj�UR�6X���[��ҷ���ѮAh����m��jn��Um�2Æ���E�Q[�ua
��T^B�V4�F#����YYbe���ڈ��r�͕+*mH��ڷ���P��,���ÄޓM¾�M����r�:��\�q<��K �c��Q3.�mky1��ӛ�ǐ[ڋw�-�ɖM�
$̰�?����ۦ��252�m忊ͺJ��D�$32}�n�f2���÷k�&LӒ$Y�D��Y��C�7����!�Q��W�H�U�R��d�PI��UvU�ct��)�2���͂m����m8�d�g4B��P����Vɨ�G���k7Q+�+0d�S(Vl)Ӊ^Z�% *&`T2�U��X���4?�lgS�ȱ�yR��7� 7�LS�ʕi��z&]�k�N�ŕ�PM��w]���]0���L���}6���m�h �2�=��YJ��Źɢ[���:�Mݲ^�
'#�1�Q����8C��q��v�7x��U;ǈ"��gS��2%��mI�Yd��ߒJm�L�k���]��l��Q膅�,^:�V�#]�����O�=��q��5��Ʊ�5�*�F��4�k,*��b�Y� �ͭ����ua�Hn�J*C�y���U��^6��B�i�B�U1�һX����)d���֫&S�C/l�dM��W{�	Ge*G^[�!	�[����Y���ޭ+!���ʍ�2��>�J�^!=тf0;���j�Nӽ�j�b"ţ��V່5��MƎ\���t4	0 (,Љ�0i�n�J�tIs4���z4j�:1�u����\���b�q�<'r���%��u�B����*tXǆ��c�I'JD�K��1`�2%Ҳ�f��Lf�LVQ��bce*�`�X�o&[%�T#�6/,�2��X�U�F��cl�UfY`����ڰ6��G(HMB�@�-V](�hx�T�[�n��Q[�;���c�.��v�S�(<�� �����V��U4갭����J��B��Q�M*�[�lշL��U齦 �ݥ�����%(i�]�^
Y�#�7btj�j!�Ub��Ђh*߮]�F��w@.`P�/nԐC.V�Kr�ý�H=T����N3��q]˦u��m�
tU��
�EXZct.=m�&��m*� -�1���bôw!C-���/��:�cuS��2�V�6�M,����0L(	B� pլחi��[l�J���حܔu4���Cᒵ�4���WX�k$�ot~T� 16l�)����EoWP�>��/wb�F+0� *�"��GD��֧�;
�A���\3\�R��,��˼oc�cgh�v��JB�:�v3hBPJVAK���h2�� R��ڵ����T^$�6HZ���"�WQ��Ef�K�^Lo4{��ků+r�����4�R�2b��Y:]�["zN���W#I���N̈́m���<p<v��z�d{�d� H�cc(�7w��"����fd0V7@��u%�� "��&Qv^��i���.����m�$p����e�"�ll{����m�w��lM�Gv�v#�$k�l���Y��ƼC.��Xڬ�,�e���w�'Yn�[-�t3#$#���Ⱥ���KtE�x"ɍ�^G�m6 ��,i�s���I�[%\OP���P����3UE ۸CD����-�@2CrwH�(],��r��]"��K�)G�n��	�ַ\k��Kc�Kr�b���!�`x���D�[�f	�L1�`T�]C��&�v�e7!jcO.�0ݢ�,XG�xPve���E5oVER�-���Z��8�[@��@V��u�c ����<�����M�P-�񳵤V��Cn�{�a)9���-*5�r,f�d��k.�nP7,m  
u�E��.���Y�Lt����1QШ���@/�^`@a�Ŝ�i�x�V�<�֦�����zԫf
��������U�*ҥF����V)R��)-Ux�Su�6�wQ�Si[�LLlH���e�J�`gH�"]��v-D�����!J�U�J���@�DZ�I/N'B���iU��p�w!N�h�xHT�2����J2��V���aI\@;��$�<kP�A[Z�f&JY������V���@0�V����=��z�lJ�m��3(�UӔܵB*�m�ӈ#z�Sr��r��ƭP���:cb�� 3f抎��HI�F�ࢦ*�'�y VnC�\��0�R��:҈��A: v1A4������Wn&.P���WWgP��Ĉl�ȕ���9�wD1Z.�
�85[�B]9��p��<[��R��X
J�,ɍ̄�i���*��q�����j�Ei��X���٭�+��u����;�Q�ଷ�m�:h8�i�z�p�yj�iF��%(k4��q,z�VFkz�5�j"��j�at���QbQ�+�M v���nf:��U�%Dn��%�`tP�ڍYf��������QX�����D���nR��Y[�6��KР1�,�����`�M՛x�*�5������Qm?�^Vކ�P��2��&-Ԓˣ��̥P	�qN=��a����ɱ��;��p3�
gor���I[#[�2���p弬�II��K@�F��YV�-V3��x������J�aWN��1��a�u��ʔ��[�°V='U�X� p��9��P�}3	u`'Au"��J{[�]l��5{d
�L÷6
Ei�wW��IQ��)�٘�h�g	2}f��!�뫿����f0CA�;t҃p]J�u��.S�w��:�Ж���<�����N��AJ�틕���hM�6^<�0f��8�k���rV�z4L�fVk�U���7L���r�DJ�#�}��)`������ocʽ(w�^1P�yXiX���l2J�Xдk����["����R���45�S��l�#��+/K�s"yQn:��t]� ���x�RY��d���o_�EZ��ۓX�� 8�T�� �+bF��{���F���ZۧB�rh�^�Z�ؠL�	Y�i'H,,�J�y�]�e�@�KU]L��#�NLЅ�z��J ��͋�i-(��d���͆�����A�"#3�kj*8h���8ᤝ��e�v+~ݲ#��n͐�@^cU+&\͠�X�5V�xU�5MKmawk�U-1�a.�Ƅ���ԪG[k�KZ����2�x.���*�Ll5cU�"R��ӓ�Z�0F�f�l�.%�Tۑ3ou��Ѫ��[�,j9)]ӶaY.�eՂq��-B)���M��º�G�.Q�A0��kU6��Ī�P�WL��;Q�,�.�ݪ-��:%d��F���Ā�m�ݙ����
{E�q���ٵ2��u5^�r�����S��D�t��jr���!ڲ�u�Xj=}2J�-�����hq��(M����G�6Rn�n�n�{�AcL�̌Z�,�������ے�l���B�k���u
�V��G���
Xi���T�o.�15(��yW�7d�Tk]�[b��3`������Y;�Ar�݇��nooBc��F��c�ַs^<�̶���Z�
�oNAi�RV����ͷg
����pF1��7m���m�apc$^k���H����L�y�j����A��2�RM!����nЬ{���T(���,�QH
50�3s�H� �U7&�3����zM���I|XW��c����75��JWq�����$M≼ɇ��֠�X̺m�r�6q:��f�%�Z��	�.�û7b{�!v��WP�����!U�]��,�7s�`eҸ7W������ĂLe%��+Ƭe� ���֦�r�Cy��aI�y�V�z��u�V���6`2fQ��p�4����	-��Ch̭�.bʼ��5��l$�;��ٔ�ww�֟������YQ`�Pe��]'x��7��4�WF҈eH �S���j4���
�x�؄���nŪ٤��)%)0�m�Wx������[����ѭ�em;5��t��&0ݍ�X�q�6J�����tK6P,̥�� ��Jl`˒;.�9���mb&8�����ȯLx
���ݼ�m�z���i��x����65x7M��ʱL?�X-�Jsv��VT��f��bJTqGJ�H�5�	ѭ5l9��&d�cwP�WH4��I�o@�1ˉ�Wy@<YLe�ӛYm�3%�Z������������/k�F��W b�f��[ð!Z!��D��K�0'��J��R�.	�n�������-�խюZ4UE1�H�׹��z6�b#lGZ4�`,f��V�����N�,+�X���pf}'�)���b�GJ|�Z�^�wG.'$���gOҚd�cz,jl&�NT�h�n,&�d�v��L�wf��
)��0��\Z�zL��fJ5f��حzJ�����y�a�7RZl��H�=\�܈R��a�ǘ��T�l߱� [vm�$;�
h�hYz����D�k{�U�ۤ1��uL%��D�F��3nkgp�ݥ��nIZ^ee�qElSV�2���a�I�~ڻ9V� M؝�dm,Ri`D��۪iS3P#$wOLwzHs5L�RZ2����[we��Л
�&��SU��S_�Uv�)ͧ�uM�GD8�i�FA��If����[k���r�j4�v��$�D1z�9Cp�-k��Q�[[b��Je\L'/C�(N� ��n�^U�ԡ���f��$Z�a�h�X�uzhPBR���Y4�T�-�c�m6�ٗ�Ӕ�>TI�R)�V���$fb�yyAeа�T�mD��+�u�I��ZY {
�[eطB|����V�/2\�i�E����zą)�ћ���U�fݨK �ua�foՔ�U���k�����[�m�E��C�D�W��c�%lܧ����m�%�3Mͭx�s0�!+!3.�Q�˫��WR�4d&XBӣ���mP�c^4��-۶�zE�t\d����3-��F�<V�Ǖ%(�Q��ի28Σw��t7wj���GF��[p<j�#���]į5Km[��,,bQh�hbԬ��I�i@c���n�mZ�0[oEEYY1�T�uڤ3r�r�W7P�pn�;F�Zٙ��IH� ���xnK�[�m�4�t��"F��V�
♆ᴌ�<���0�V���6�Q�x&�2̍(�I�a�YR[�u'��Vn�U�B�QĬ!��Ks2٦�"M�\Z�d���W��s�:,�骬S����xM	#�.��b�ݧ���U0^�$�*4��{,M��>� �od4����� ڭ�
F�Ȯ�'�e�`��-]
5n5�b�)�(��ڶr�ww�P���2]�-�,��Y�%2V��U��O�ܽ�D%K2�j[Ha�����F1#�9b�X�a��ⲩ��Bw]����$�^7j�d��me�Nز.h[HlT�����R�P\gnG�U��*ł��v�X )�]�IV�yڪ��T�)�!�N�Y�	F�|�`7�FY�@�Um�	I���ݧ�sz�.ݛ4S2g\�¢m���#������F檎ᳩ�J�ax��8F�E��R�S��2�V�
LZ��Y&i"j[��a'a���=���;��~��hn+W��z�ݨn�G%�B��f�i$�]�[֞!}W��wѐ1�ݼ����u9H�zup���͏_m�F�DS�E��!W�o�E+	L����M�e�J�P�3T���m^V�R��὜�Ē�'y%])���9��Z��2 s\�,B� ɺ�(6����,��v���}m�>�ļ:�*j��;�<�)y��Q&�ʲ!F��N��B���Z ���m5�U�̂���sv�X��b#w��h7�.��5VE����ʌ3nȩT��ޡ�е2�g|�mj�]J�����V-xX�M�����E�»b�B_m�w��b�9��W�����Ԇ�̢�w�(�i�y�(�+e��_%����	��d2��#y�GU�h7F�B�Я�����yM$�3q]Ï��p���ܡr�B;X��i�k�Z�*n��fc�os�ٗ>n�°�:;���U�Xf�D}6<A7!���\��.�J66#g�^�Ǜ�C*�y�����'[�RX��[X(J�J�7�Ùl�Η��qK�3����dY�� �Ai�Sz�v��tkBf�Ν@#v���=��X�*� ��/r�[aʼ�w�P=j�����;�@��%�*V���r+F;=�+gw꽵N����3]d9n�h�VT8%78vV�C�](5R�D�K:`������a㢶2�J�K-�덖+
��R�;r+��Υ|X2j'[[pP]C+Pղ�!b����ӝ��(q��q�l4��]�ȥ>QhR��E��
7���k@M����t���=��f�.�վPF��]yP%�g7�Đfw-��5��+��}�-����)����F���$x;j��5��6������uî�>��"����閞�
���m�X��v�l�44���ZЭ�9w"�+	55�]��Rc�p��;[ಢ�/M	 I�ۡۼ�����loh��@�w���ĬY�L<qu�Ҹw:���i�:/vq�ݧ��m�����MFM_ga�u��ˊ����b��n-.齥,��- �v��X�A!uܛon��[���Y7t"a�;J���+�n�5��w[������RFh���]�ZM+Μ]��Cvڬ���G�)�)4�]c��3k��.p�������rŌ!��z�!�RoRC	�d��7[���M�;"[ˢh�!�K�r��^&/�[}����:�2/�Xϛ��� �?^��8���=@�������S����f���d��T �+inv]on3��l�[��CL�6���m��t��_P�C\
� :�M�����)NY.��y��\j�%����+)�t���<��rmV��9M@�&+y{����o1/�4Z�CD�-��>�u-v�d�.�yK����rYw��Ƚ�o���HX��h��x��-�ս3MpȦ�
Y�^�3���A3��g��!ɝ��)�yv\�wX���nX��%,P̰�5i੥�B�4�����9��
�!e���k7����Ν7�VkU̅�`t���7��xD�QЬnn쵱���b��m�RM�J���v����}��!�	���b�͝(�G{�e<yMbL+y�%�;k����wb��]�j6����
�`���+ѥ�c�
�l��ѽ� ����A�Zw�)�q�������������;9]p�
�ta@c��F�IcH�sGo�}�������s����n�v�IԢ�b�.[<1�(N�� w��';%�k��*c��B����yW���]�B�3O��B[�1��W�8L�2`�u��U*����PU��oM\�fA�]�;.92�2wa��9�tV�G�rf��I�;�	d��V[����i����d��j�إ�V�g�׎pp�J�����0����w����9ͰGZ�vL8���JK�᧶�Ϋ�B+P�[�_K2Z[�ZQD]5��ʙ����,�O�t�JE:��c@��K�2*-�(n&���O^no	@�N�DoN�K�������ACi'؍e��Rnڊ���QSN�b��]ov�L�o�򱱖���e��2����,Q��&�(]˫�],++�� ��y]f����z5���8�X��O;/NV�Q�m���b!J��.�q��+-iK������_k�"��9�偱(� �i����nJ�FmZ�ZfV�)�Y�P\e&r^I���G2�#�]'u1��݇�vfJ:��	��ڳ�l��l�+�"��\^���ѪW|��[�S}��hC���V�����8�VY���t��֪�3K�B}��g]�.	��s_(b�v�_S��r�����M��;��x�u�%s�%VvgV*�9�{�Q�E�K��	����u�YZ�!I��/�z�(�1�ݦ-�@S4��&{?$��#+yVO�%���k�Bbo��0�rh<\�F��׻e=+�Q�e%�-�y�7�r{��)��9��;��f�W�7��rFX2h1u�n���f4���K6���]
ŋ��Tm�2��/����d�T�c�y�V�3e����{[k�W�V�ӱ������)���WFhĸU�����O�<���'lʚ)�aejn�a��\�}ܺ֙Ҋ�	�[�v1m'�٭�՚��5]�ІT�̻}ţ�9M[9y�ح��z���֋Xe��g�]gj|:���n�tسnR%m[�ծ�#���^��o���˛)=�YE��A�a��y.n�v�گ2�ٝ�����ޝl�k%��:-�����%��]	�(��):��V��y3*WR2`C�ËK�����9P,���j D�F��yM��4�	������������1_J�7�����3���V�P�D��B�r�WsG�o�0M��av��P;1px]C ���v}�|T�c:�Ū�&F�C%kQ���>�N���ֺ���/D���/4D2������R����iL�B%�q�Hn;��v�g���(���_�I�b3�ߘ��q�y���e�45jj��_[8�TEj����)V�6�������,@\�)C�Q��Ln���tes�`�]��Z�9EY@��enp�C��»ov��$<(<V�Kl��(_ӈ<6���ć�
�HUɦ��D	Y��1��eK<{�T���N�p�r޲%N�.ݝ��1Τ,N���`q�yi�~Zl���Y��V	XhR�,<L�Q��*;��Rk���Je[j�C˭��)t��r�S-B�C#~N��]IP��1��$0t��p�0�TP6�[�Ú�G6����lp�ˑk֞����h�v�U+p�\����4f��)�q֐ܚ�l��v��ϻ��9X۝uiDFA�@��b���ڻ�V��2�F�,j
�}
�fə�����X7��}�Ǧ�fj��fk��q��c��ksxM��*
��AC!��V��8��Nm|�kl��[M�K�(�:NN�>�S�l�$�e����W/{@�;r�W-t�"��Z�D%������]'��1���]0�S���%�Z�"������Z�왯ti�έ'N�Y[����TrZI�N]�&�M5@��&noTjn�CY]���p�C~��]�g�0��=�$���6s���n]�\yލwx�������c7�d7�p7�jo:��D�`dS��k��Bn�e�6��^��IsF3ϱ<#X�{��J��p>���O��Ɯ�f��+���p��u�]O��/�
������b&�_K�Ε��2u�en���������u���W��3`\0Hv�U����?n<��;w�'`��y;�5��wt��քK�X#��e��lOV')�pj[��ɊL�Ji�y/�Z��w}|.!2�.9v��$2�m�A���5�_p�`��;q���1����S��i2����klޚ�����{܏Kq{l3^@^
��a����!�[{綇>Й���VL��3�:��nrN��<���Ck*�D�6g7oOV3 7ɪԇ7Ѯv�S-���4��h^�_�D���J�u�٨�+������]�/u�ލ$����Fq=��F�Y����R]M�N�o��Xt>uo*�}�TV5Y�̸�12m%J�K���|z�i��o�P0ܛN*b�^JAg+����7Y&Ѧr���+�u���d��+���s���a�0A���Wx��[e�W��g�U{Z��}Y�$vK������f^�o+DWnN�:�o2�r(����=ٴUI�άElk#��'��7�����cz��Lx4!��kZٹ�k�)�#����7��9k\�v�N�p���ޠ@�i1�)bD��c���FX=(�����U%	s��Gxpͳ��V+��-��R��_8;�Q��B��3�^]d [Z�rwr��7:f
�D�,Q�9Y]��d�k��˝w��WK�&��p�˚�ʙ�NU�9�$��������N�^`bn� ]�s�gfI���V��˅qt�.}�;ч9}i�j�J�J�TT"]wu�)%by�;*>Nuj� EY�\�7�'{"(:�3�������Z��{��l�v�k*�H:ܥ��=A,�$B��x,�\6+�N��Gk	@���/����{8F�Nl�9�ǹ�T/K��m�[W&�=���(�G�JW)ul.��(+��\��w2�N��Z
#;��;(W'cGi�ifV3�e��h�ec���w����t�pS:뒼V�f�n�^�Y�S<@�y;���4�8�J�;��/���zF�{����围L�������N��C��@#����p����@�c�^=��8UC0�h���,W�'�*��56ھ�Nk�.��*����%L��F�Q`�1=T�:����^�X�P�����%����s9�8��,jOaJgx�s���7tf�b���_-��j0q���
blQ� �Y���#9[��9tѦ��B�aЌ� �^��S��� �Oxk�����k+pO�V�
:"��-Rv6�1�'��)�H����f�19�y4����qyHm��8����KMz�9P�vv�D��s��Kmwh)�@^P�­2�da�z��<�b򡫹x 8K`Ǜ�9t$h��{H����w+:��3�%��wvʓ>4�7�Q��#��g�]�V�t|�+�m,��}�Y�wWp�����2�Sˎ��ވ^1�#f��)�t��Z6��c=]+2�	/z�4���bPR.��x�V���/���Y{5)�Ú�^�m�kv�-�a�J)i1�H��A�����-N�1��iÁ:W�`"���	)S��8p��:oM������&��S> �;�g'g_h�}}Wz�8(��L%�t
�J�԰V.�a8���EJ2/���b��/���]�7�ʉ���!�	n��=�|*��UƲU�p��vg�)������cV��kEm�7� ��c[Y,Y�@3�^��[�L.yd���"���P�6���4s4ӺW�R%ҹ�|�6
o{&*�3�ɮsw�`:0Ak�J�%S	 [U��,}�MCL�cX�;�|�k��K��O��u��]��mܠ���2\�y0gG�@���i�*�0;���g�C�!V�ˤ59��V��y��P��K�u���M��>A�EOr��F����'Gs�v�.�w;����s0Y�Zke,v�\�=;t�v�8a���{��]ShI3��1�6��ijh���@��q�A�wy]�N�����:�w�o���T�D�5:�;s)�|2��B�^�u)a���3�8��J�=lKT�[(�c�n���6r
:9o^V�U.����7���4�KN�ou�J�F���p��GԠr��]�q�ĩ�u����+%a��+��� �L���^ڴ��Z=���?X��cl���
]�����u|��5��� ��>3h�(nWpK,bk.��>�Q�Q(� �Ө��kou8�6)%�*j�c�Y"�I���:�G��.����ᕘ�ZW�GW�"I��1�Ү8�i��؇`�����S�J����;iɡ�yq��ۇ����w2=Ζce��;����)em���]q�c�gD%��,s|��s��Yl��v�VR+�sP ���4���gp"+�T VoV�^I�@1�n%U��N�:-I]eOWuM����\�s�EE�R�v�y}��jsQԮt�Sx��r�	�rQ��}+�ER��[�Xu-Yokn�ma�ZKF)�H���(Z�9��>��(E y��ܧֆ�`�1X���-�rT-5��[b�jc;��Ԫ
x[�stҘ�'��a�y��si;Sc��2'˻$��7����6;������v�Z�9Af�	ĠQ��H���<�|7f	�T�zrZw�r*۫ʸ�x�fu��
�NJ�SoI������DY�{�b*�H��l��]Z�p�s�����;�"��ٽ1%�6n�S2N���*�.�1��̸n�M�1 ��6��(]�z7��];�yD��мw����;y���֕�@ j���W��497�[��S�2V�NW�+�Kd��͢� �*�Y��돺�t���d�
ɰͥNl�n�tk��K�s[�h�d�� 2sۥ��2��n	�.�I��Z��&��Χc�sFU�|��%Vm�<C�Vi�sw�Ԡ�8-����9��Y[E�;�^���uӍ��uK�,��s5�VӐ�4�/6��9�/�˿��M����e����
-Ipb�>*Y�e�2��ά<��e�ޞ�ǎ�ck�ot[�~��vw��].m�� ��O��n=(ۗϻ�\�X���m����v�Hq\��n��%�]�/� R��_L��#Ӹ�=Q\~9��nʝ༜ҽյ��5F�\��2�;�\�!4��)^j_�����HH$$�	&�����_{�fǵ�~6t<1G�b�[[q8�WwD`�.U�W\�*����yWZ�f6��1��{X���W�>*&�f�۴�f�Q�j���k��� �/N��ӆu�۹�y�č�O,o^0��A|@�&���Ů魶��op����|5��8�rE˳�5�u�f�j1C���qD��"�՗�y�۲��T�j��|�MرM�d\�v��TuՅ��t|h�Ғ����&�q��}��o3y�c.�r�2�8d���U��0g<@�Yk�M����+r�'��C�Tt����:g�wS���J�� �a��.�(e�ҰS�c+����(��t�<� �U�x4����tmi�i�ܧzX�4���f��8o=�:��hE7UI,.h�Κ��5��!�(��;�{���F%�,
ܙ�W$���wV*,jq��2����`Ն��x&��eH��d\P�;�{�ޡV�*#{W���������s�M���C�ne��B�<J�j�D՗�k�*4L�}��i��2$��3����d
���ĺ�(J~�>X�]('������`�+5\=�Y�j9��/vlM�-�B���.λx8�!!W��S�%�S��pV��K�}���S��2���J�1d�G�+�g&���ܰ�x�㧝��z*$���s5�S�9��\�-���B��|�
�|�uF�5��$�\�S���	���Wb.t�[�:%�w �9\{� a����ru����S�x�v��f,����pc��t�d����.:Y�>��#�ү�t��}��#OI���w���)�G2�I��ށt���>�)�����<���ϥ5սݍ흎&�,�ܓ#��#��a�Z\*gY���t�X�Ӝ�Ю0+�tn��ҘNPczՐ��1>S�魛�-7�ec���Ƥ��k;�|��XVj�[u�H{R��fZ7j��Jl`*�;k��&��/M e�=K�4�L�����i�:����.��	Px�o=9�Uc=t���,�,e�5ro�/�p9�u���)���5Y��� ����:�aN���*�a�}V~!�k�5�r�,��9��6��!V�G�#�[I���I��]��U>N��6�
Z6��-�M�+�W��wqp|�q�;�e��E��&��
n���vi=�R���[�v8h���
�)Yˣ�ظkY��V^�����oh9�P��ֲ��;�1�9�u�F��ɮ:���"꺾=�j��}ң44�P��>	��X�/,�&�hnØ벇�7�:�Z�Q8/�S��l3���J���|F^^��q�L���$-PR;��S��^�yQ'N���:[�-[�kN�8n�9ŀ���ݜ�fka�):f��vVI\���oq>�)پ)u�jE�ÜhK��,�����M>��N
��w��ڹ5�"�W���	Pb�M��8V]pʽ6�J2�\�_m�ʚ��i^�0<d�|���������]GjpL�˺tY\���D`ړ��E��b���6���!��mrݗ��Q���xJ��8K��C;b�׬��²uA��3�vV�é5�7,�᧓-�&�1����y�Ggd��b�uut�y���glm��=,�o7�Qi��WP8��E�wr,��`n�֚�g�R�nP��e��ˁMfZ����N�U�V8�Ma�јe.h��h���1
��$�ѩW��v�y�Z�����F�p���4��;����}�4�g����*ι��+��2�5S�B�_],2v��D��(�Z �o�+���D����J3!�y�H���:�.��2�4T˲��T����U{I�װ�Gz´���st\c��*�z�.`|QG{o;ȪF3XO3��2��$;F��F�<
!e�j�u���=}�	w��\0@4����#
�p���;cOG6Q��#y�� ��me������WIQ�y^�w��pq�`S��k"W�[OEY�2��O;,V�0�m���X6h���e�㖰���X��^䫥�P�X;��{B�Iq%�fJ���W�F<���o��t�*���k7ى� �b���E��C��S"'M ��
���y��q�$U��F����}�t��u��$�Nժ�5��;q�i�$��b8����v\�ǿE{��"b� }/q���p,1�8"������Z� �.@�)+�]�����V�'B���Ws.�UJ�ʉ��1�!H��z�e۵���p%y�H,�4��*�b��2���p�9'���ç)PT�mڮ�[p;��Y���T4��x.�"���M�C��w=�j̬Ј3�q�J)�-�t�d;��*������wx�$}1W	 ��,����}hX���p���/C��M�R�kN����=�G��iVme�%	�T=��kj|��'P�L�X�Rau^V=�����`��G��)umnAW}Ղ`�)oepU���F×$ٕ�+դ��B՞��[W>/�����=cee_O��t�o-ugX7n�k���������[�(Xh���](*f�z
�Vf�c����i�d�
-��P#):כY#�G��\���[X��p��C; �B�^`�ɵٙ��mc!E�l}��{��1�L�Y��yb[���B�v6U\��k�Mi��ƾ/.�gp)��9���}�,����NVt�I��3��.99��nE�t�Fq������"�k%vl�4��&��ܥ���i�AѰ�@�D��	���.��7���˙�^=c��Uw���V����x�ֹ�Ƶ�m����A��\/����.�5`����n��;��|ƶK#s�
掫�A5��Jp�aTm��-�{��ȑ��V�k�4vWl���-u����N�M�P)[a����3`�ǯ���n>RKS�Y�J��:����)n�e�+1��-��Z%.|�ha��x՚}���<�IgZ��-�g1����Պt���j�-��Ҏ:�HJ���V;�=��7�>޳.�%��C����,]{��p�6G(�:�ZR��;��cU�h�+|�ty�@����E�1A��m�RaѬ'{5Нse7 ��u>�*��6	�Մu!�
��l�(K���T�:���#� �oU�Êd�)�l����G:g\�~��}���zz�.�����6���.ۆ�u�;�G�ub$��+{'>u0;
/Ƶ��:w��ih��oo�&,_�0b.S���l��0�� �i�YY����64�ŝ �Y�ľ6�a�xpgυ���u�`Dj\9�:+t�:���7r����N�6VoZЮ����]�3�}���o�wT�Ļ�f^d��RK��i�*�m��Y�a�o�܃\\�J�ʕ���}Wό��*zЩ�d+v-c��5��i)Q�ذ�qua��.�hIGV�	/k�6�} Wq�`�u���:��*�Աݍڷ�p隨�j�c�/8���*h"��� ;6\ne�ɯC��V��=y��2�E�r��[�Wj
�+��5�X7L��%�J3V<6�����%J���2�c(q(jn��H�m�&�<r_^lq�C��Պ���	�`�ǀ�n�=j�;9%R��,�)�f����'
 }��̕�G	v�a��K�Q�M� ֪�m����o7Z|�N��gI8Wn&���!����Zԥ�����h}�U�7�P�:%sv����R���v�ƚ&�[�n�KӉ|��f����<��Q��2��Sd��d��ߙ����*-�;p��!�S�o����[g��e�-C�Xx�h&���ZO���M���2���GGQ�#pN��AI2�����iJ��˚鎭!��2���++]w��]mAR���:�v�$������n�� ���Cp�4֧]c�hCeh98���W}�&fX�r�������q��|��w;�(^��WGYK���T�޽ ^"�G6Y3{�7n񯁽�'o^e7��$3B��B�`�k��s5V�B��Vs�V��f�)��Ns��VxΕ��(��Sk��pf0(�,M�Ӽ{��=X��BS7���B�/7Es����L:�Ku/k4.}\��Ҽ̍q2�ֵ飣�}t(b�E������L	Օ�a�5��;-Xs�:Μ�Ƙr��\�YH+Y6�P�0ڒ������O�D�f�Za^l�V�"ن�1r��`�CK�t����j.Y/p�<M�vdJݝ#��h�B��B��u�_p�7fN��͏�f"w8�/hk����d>��2�҈�bAJ��f�!�p�rD���:�&��\v�8���de�&�dw��q6�j��>���gm�6mjk/��>V�t,;���q�C;o6�l��,��X%��P�k/���^ZzC㱽��V���"(]�}����������� @���K����[�c�N�o*dέt�S�)�ֈ��ٜ�J�Qƍ�FU� �uf_��顜du��ҥ_�ʹ���V��=����S�ڠ�;{�`B��#Yl\r��,Uܺ펆_P�[��I>����6G.�qf�k��Ӕ��>�{V}Õ����yT[H��j旎Lו��<޳���K�A�46;p>R��(E�2�v@e�^�sO}�r��#�V(B��ٴm�*+�� ��3)T����� �ir��%[Sv��(5S�h4m���&�ַbQpЭgh�8t�v[T�����]av�Io-��8i�X0pt�Y����bbWv�}�`�SF��&g&ƨ21�pי�p��W]�h,q$mo�i@s]�`��i��yK,7&��t�c��|!9Hb6�D�L4��4 ��o�jA2��J
�6�����:�B�롼/�\�u��,�5u�i��3NnvK۳��7On|�$�۫
zU3"��s��x��o6R��8j�na���Ћd�V
��\x�l]�ivҏ��2�V�9�}#=:^A���,�*���;�����Ye �u�euej��u�w5v���ri�lm��fY�F�c�$y����2Nw]�<
��]�Ҍc^R��S:�0���Y�"[#�2�>¦v/�O_�+�#S-���f#N��)���]��Wܹ��M��=û*!N����m��lVDe1�s��19���mn[-�-C����f[��m�V�t�g��Z4ޚ˲��@7Hg#'b�ϱ9H�]���3|�h�o�s�j�J��X��r����٢m+Z�T��zGgx֡�e�"wq�\:����d�y�8_�h�6��.VR��h��K0�V7o��f���3P�]r����X�O(�am�|�䭢��c���j���5�JL�Ԭ��l�i))�zL�sQPJ����5�3�d��|@?mrU����O*�¸h���x8KR���T�����y@��ӻ.���`ks�
����-�ǘ|�U'8�����W%�"�Os4�%hݖHjub}���@fK쬩�23{�E
[� S��+�]�̍s�A{-갗V�՝�[̵��<���W��9�U��=]�8�ib��T�85n����݌�@�A�2�^^�-���Z4n��;ee��]�q�K������Z-Vm�8p�C�n���L�;�8#6�kӗ��Ǎ��s:0PtQ�śC�M�6�r	Ѩ'�I]�q-�ӝu�o�Qk�"��̴�P=���b�	�+P�8�O!)/+w�ktr7���զ��la�юu�zq�V#B*��������\�ꊞ���qy�qwJ!�p�P3w0ͱ(Yb�N��z/�j��Nr��K��Ẃ���8ss�[�}���n��9���u��e��7gV�o$l�shX̳ ��;�݅�WV�cXk/�]iJY�,4���Y�OT���sJ�b0꾉���[Ζt˝�Q���q���ۆ�4`�Q^j�SD0�f��@���W�3��ȧ��K��\��ᚹ�}�%�e��r�~]�l�Zl6�]���ˍg/O�"����Q�s�Z�5�DF�2�ԣ��H+)��Ӂ-�@j{1��ٔ6�Mɑw'-V֔�����GQ��͘o�Μ���]��y$+/"���Q)���G,;�J����Z7Յ� r���R�O9t������u�NL����p����P��y9�iU� �1�ts�~xrn	�*��6�fp5����R���F�{�{i�����#9	���С�
N5���=R�M�1����1�YZ��l�utK��3ou�(3G\s}uv;����~3)��Ε�=m�}wpMn��j7�Υ�O6n��焝�arY��G2TN�Wf��k�q�m-�=4��Ci���
�����+�pF���{:��n���V1�s���i���]nVQ�K�q��&cw5��w���"�6� �h_��Pڃ͟ s��¯���xљ���mn>]*Y��;X������G�����
Ѱ*S�6���a*
�\R��W�6%�=�ُ>
{E�2i5JEa�O�5ϖ�&D0����q�[s� �v�w��H��N�-Gٶ9�|ζ*�e3m��Eg�@��
�6����6�_5le꠆2�:+{ȏrr�9���?,�t"����h��u�zr�4��t3(�s0�����]�s�}1ـf>H�I*L�CL���f��{�8�5�+t���bd���Y�G������yK���-�;o1�	����N��G���Ká鹃g7+,:i�g�%Ϋ�}KnŢ:"*�9��*E����]e�E*�_]���y�:"�j*�a�|�\�WNR���俱�w�?T�6���9�ˊ�u8;]������J�?�=�����zÎ�+��V߶"`�H�ϰ��}��4�����M�v-Fb4�$�������Y\OQ�N�z{�XLw��-t���X���id{�^e�8T�o���O#(�K����-w���
�֔�a�zyN�۫i�s���N��6���˱���-�㖖��6�X9g�ugWr�GK�)�);t��c�y�¯�Uq��9��I�[��F�L�ʺ3e����2���=[�,�Vr�
�z9ۇv�sY�P �I�v�)�s��8��0\�Y@_u�C��82�V��9գ����S���v��81�1V�!�(���$�+5ܼ�S��!l�N\g+r�ݫ	�oq��:��mL���퓖�}��`��n
~�U�S&��.����d��=�4r���_%r�k+Y��Q�e͎:�
!� >��8�&�=[��qv�;:뵛��*%as9��-��w5�-�b��������^	���Gs�^�!f|�C��bA�&5�
���a������¾�j,h�e
֡	P��5��+�����S=�}���la��ʱg�/�L��oN�ӌN����gx��ۂpb�Tԅ��
�g��d�7R���9kTH�����2�]�E��X0+�S�&���iw`K�> |�M��D���kC�Y4afމ�Hމ7��v搌��0(>��\*�3?o�3�=�}����b>4R$H�#��UUԱEDKV����#b�]�PX��Z+�+`-KF ��EUX�m��6�1�6��E+h6�*R��j�(�1Q�Z,K)m�1�1�*L¢"��E�1AX�%b��)mrܭ�Ī�Jƥ"���8���m�s�Vչ��
f�TPP�Q��nfe�J�UKj̶,D���QE#[J�W@����UK �e�U��@c��R�Vc�*�YDmUjU�
"��1�DAQTX�V�F ōj��LB���*QQEZ6*�`�mT�����UDX��TQԂ[*)-��n��UQEX�8�Qj�*�F�j*
EmF�E��iZ�Rءe�-��E`�F����Pdr�c*
�B��h��i�QU������1�����u�Z;���q���O]���w�@��̴g)b��ʙ�om�!|F&PH��[�
L�����k���< �?��9�ݯ%t�S�bu>����b����uT[�2�k��Ğ�y��	�&�#�[�.�)�)�B1���:
�3���K�ً���2�٨�T�@r��؜�$��nJ|+Z����Xiz�=U�w��;�~x��騕�8����Z#y���&��V:�1��nF�����<)��~�l�T��P�(w�ۨ�K=������ޫb:*���r�P�'�����1���l6{]Sږogڽ�Rέ�uI)���F�K�rY�}ݥ�x�p^.�`{w���N����j[Q���]�F,P�Ḽ�{]-	�%^��RⲭV�[kZ��Gn�j}����t��5L�M8��L��)v{b��f��ҽ�Y9��S�˼��׋l�&9�	G������Y�%�'OT�}N'Z�����DbN���������1�͊��n�7n�ʹ4@;E<�.������z��ee�%z�e`�2\F�",l�!�b�(>��θ��;��;����"�4�:t�d�;mh��w �q���u�c��)�v�-e��Rֹ*�x�R�ړ�9�[eYW"��LѴ���]��.��z@�np�c�f��0�Q�����gCz;��o��5�� p��,����*K^%2k��A��X�f;~[\�YΥk]���e��ʪ��f�4��Tb&1��E9����gƹ��;���b����:��Sŀ���m)R��n���i��������v:��:2��ѯ`cQ.�d%�W�o��;�W=&=�O�rY�V4�\�6�n)�7P������Mі���̚��~��A�=x5<�*�9�M���u���
Wf��ݜ��Mn^�"�\F�!p��MJ�aep��X�}p�V��\4Wb*��8��Z��0��Ц)���j%t�b��cj��l�z^�ŐosX�f{����a\6-7t����ama��Yk�c+����iӏڵ��������t&��^hd�wS]b�F�\��N��Vf�+˕
���n#��r���������`�rY�(.ו���2�P,j�s��=��>ت�)ҽ�8Zx�a�e]������®��tz���a�q��%>�]�v�l�pW)(ͱ�khJ��g=�k<e�k�[n�ٴ���{4��q�7�)dS����c�ݬOog�R.%vwH���nc]�&��Y�GFU���j�)�v�G��3[�3i�.U���3/�mA�p_��>u|����ս�mMS����5�{�i�=���D���m����7Ƃ{�9^oV?u*1����LɎ����Ww��Śz�A	5�]�	�ێ���*��b�GE(3��Xj��ʻ6�C���ؤ�Xq�ʢ�v�Y�m�N��S<0�]�dR�/Gm�WV6�k7-��!7��\b�1I�E�c��d��$f3�E��z#^�x�[�{�֝��q=<���F�t���{ٍ���c������Υ����C�g� fsoS��5���{;#7�Vj��I��8q�7�7U��T�ՅKh��1�b
��x)�hsY�Y�y��@ޜ�	^]gr�"{2��=)<��.���Ա$�\�h��N��APr�3.T�z0Х�t.�cwXR*�כ�x/-��w�v1��ݮ�I�
p}����I�̊7]V�ډ�����V��ݸ�EX��u�V+C[�ҁ&]Ԇ����/gSk��[�KŞ��ؔ�1'����ٴ���=>����a]+�.��tc'/S.��+-7Z,T�aF#<ɡ�p��^٨��J��c�&z�USI4���er������I��zɏ�l�K��gP5_v�ߨ8W1�ٲg��>:�Fa^>��������^��KwNt�g��(�ʞ��w�>�����J���feҽ�u�EGr���kx�eU%�ܻ2�n�z�[�Ŀqy��oҊ��k7�sK:�>rz��K]��X٫��<wS���Y�%{ٞת8{v��z����uK�Q����r�g�zd���ε
�A$ys;��f{�1���/=���,��]�@9<���Сt�:�.��˧%T=I����M�}��ې��-�n[�����+ ��z�ڐ�����`HV$��v�Y�,����*��*�WX���]byA������4������G�Wj5:�Q�;i����>��[�����*�h����r�嵥R8�c��>����ÝO�vu���@�T��*�ԭ#K��'�dIE�y}]�Z�ټ̬)	���g4�q%\���h�.\�zr�J�GRc#�$-B�����[��7������:vQYٮ��M��ggǎ�;�����Z�i�/zL��%E>ҥ9����Nl��{�L�[}X�g\ƴq�����kZ�l�t���=#-�Q�*A�Y����Z�y�:޼�f	�
�x�{5������`�zcx��OY�Y�)T�Ջ"�^O{���yV�#y���ٻ�/��5��Z���ˮ�z��̪޵���T8�����t����(�1��
����/6�A]�����sS�7�ϩ��_G+jW�lNCo;s0���lJ�Y�
{���_v��d�+�����T�9�.��3��u�lfU��jٛ�x�'���<���oҡ�УY���x�Y��-�k��r����.�<P���دrŢ���o��-Tl^Lw�T۔�N�5��GuV$�ms3�Î�zɓX<�Ӗ�uY*����љ���^�FWfԙϝ�7I���%�/�a>�A�G(p��Z�]�5�F��js��������޼2�6���(عc��7i5؝�˕;���V�s\X#�'s ��˩�ڵ׫����\�.��Z.ݯ>���K#���k�9�zT�\���^���yd�y��Te[���m�?u�y.mUOI��2�^�Ƕz�U9�u[���sI3�O�����x�VW*��YɬQ���C��P"�nF�|��59˹�f?*f��K��iD�Q�И�I��︾�ڡ�J����RhY��[����T.�㒀ג���b��!j����Y;uK������We��n��*�gN������+X������z/.e)�텮LRO�C����s|��^��cc\��E���8���<g��Ck�uJR�y\rn�Õ�\K{�Xڪ�c�Ȍ�C��D
O�:��wwз�I����K�:�9+�+|�{�ڹ�|�bv)��:��S�����I�ds8\�Cy��+s(jy�U�\�.u��3��.��k���<�I�T�r�b���K,�y��ܽ�#�c~���(��M�Q��F�#H>z��2u�\	1��I����w'^�=�'��F���UiS�ku^�_+���ݫ�f�S��dVvӮ���g>�\�g�A���Rᛇ�ż����O��oq���ֽ���4Y���v*����Uyޗ��5̆9Xi��}\8�n	��:<�.�/چ�AZ䮩���ck@�j6��x%��n��6%��$�9p�!�	�InY�&=g��¶}h[�hl����k���'��j878*Ӄ����q�In�پc��y���-���);��3���UFs�]��|*<�-�ɇ�����ѕi\�WM�w���}����}A��{�8�1����Q��\G���j�-��|����?_�z/ͩ�Nu|�\�p~{�j<X&�<G���]cgJ��!x8������=�ޱ�a=���c�Q��u�Ϩ]!��O�g��#�}\��%G]}�ێ��«ā�E��iD�+vo���fZ�-L�۰��i�)|����fߛyQ
h(ѷ�*R��m�T7�=�X��F�����7��d���V2�3���L^m��fS�8���+��K���\�#��W��"��?o\GJ]�h��3��Tm�+�^�·N�.�<u��m�C]!�7��������v�[ںa��6.n�KzIO�$*k��%�t��K;�+�{ן]������"�^8Y��uD7A�fGN�ò�l���Jrj�K@P�+��J��+��O;\9��K{��n��rz�{r�n�xU�>�tQ܍�{\��;W;�O���pϰ�~|IM�_�a��]s6���щ�!�Jޣ�)��������Z�suR�OE���y���fS�sP���p�+zjV�[��Y2�JT�ڪ����n=Y�V��M���yE�:
��CD��q�.��v�"���}�OMܾ>u�چTkc�)���;
�g:����ئ�9����)pW9�N���wNr/���'J
ƴ3h\�ܑ��R��]鼪�������b�UG�3����d��Ҟw�p����m�ŞX�{�{��U�1:�'=�j�z\�O�<��=�*+;���/��&��o��j_n��'L�q�t�V����̃p�+$p�&��0�'!�cmLP9S/�!�������P�^&�u;I�Ǵh��)r��覞$�P�8����F%����f
����,��a��o^�:���cYVb��ky�[;��ɍ~Mp�Y���ݧ��^�º+'
�:����W�Pa����Ƥ���Q�8�V�ͪ��օ<ow�ד�ݽ.�g���&ӭ�d'm��ۭ�s���]**����ҫ/S[o[��;{����57�F����s�3+����i89�i��֣�$-sp��ZˌiodC��Q���i�_F5s}̵�{�v�z��mp�"Tt�Rb{B�B�r|����1���F׶=�&�)���2���p�v��uW��Q\/�y��H��;��}8�B�RW��;Kh�C���Fާ���6���9�~'�A���K�5�Q&�>z�-�5/:��ꡝfL�=�tQ�ֆϣU%	LG<�=���x��,���П,܊n�n)�rX��t�wM���ޮ����܍��|�����V��f��_Bsm6�]I��vcѸHH"J����������X�љ�L�ɪ4:��ݫ���{�R�V<o�nKC_u���qj��;��Hu��3ϛB����<��P�3�G�s�����Wi ��|�����S�0�ዤ��]_v9[{W�V�ڑ��4^U��5 ���V��w�"V���2c5Q��\@R�������-�g0�wf�ZS��y�J _f���<�.د�W�s�͑W��
��1�x����	䕎��9�n��+룮J��e��d����[� d�3[��0t�ۃ0�QP��g�k<���6y֥��3�,ˠ#��ulN�N+T�|��\Tc�Q����¡�s�r^z�R6{e���fV4'�S���tq8T��_\fʊ�U���n���\��r��n��w٭�]J}��m�m��\��O��T�}��t���n*3gmL�Fw��?z5}�Z�J��8�7=�7�J�pM�01�~��)��X��*���R�c7���;�[�����$�?6��Ъ�R�9Q%Q:�TN�*/�!�v��Ӱ�`ʼ�:��m��̵��I����F�*���u��4rR��J9Yf��ܬW�e���j:w-�YX
;)�;1�I�X���p�2	)�,ƷF�Y΀��Jt:��,���{�x.���L[n�Q�
-Gf���;�]��R��ݺ[k��	�r�wlBcp]��R���t�-��4ď:e#`ؘ��ِI�E̲���PV5JWoj�z�ޱ+6���["�����
�-�����˘� ��Uc�� 7d�SwM��C`�	1�V#��p�pǽ\E,�3u���22�#�_����{�8l��h�179��â{	�ht6��\l�9Z{��Q���7�Ý�F��Ne	9�ǆ�n1�����彛�NuLQ�F*��(�������s�����J�Yy�WYS4���a���]��O�Fd��f�-C��<|�k�Hr�(�(r8�Hn�3�kU�*X��p�B��ox��s!�[��4_J�P�w���w.�v���*v��T_fb���˂�q%�xء�8*��Eլj�mF'@����Y��w&�
�ep ��y9�Yt���qV0�2�pWB� *��)g7���O\�����Zxn�,u�9���]�q��ܥ���S��D�Az�
me�vMvm�5g�IR!d��%rㆎ�l�}�)�80䶈�36�'��8�����س�����2pH�s��'Ce�s��L���*�2慄>����Ȏ�Չ�gt��Ө�\�F���\�#����$����� ��-b.��wJ"��*�霕�n�vS�r���.�����nܬR�3��.���Ӭ���\��eئ�ʌ��+�6��+2���u;�n�gT�§cU ����Lޗ�2�1 �v����e�h�v�X`."�&Wەػ�r����3y�`*ԥ��*�q��D;��YY��ط6]�v��1Pt����n8�p  HJZeœ3\��p[��R���ܚ]���Y2�rz/f�W�5-��Af��:�sXP��^���w(��얨�X�S���s�Q��5}����Z���ñ�h�҇/x,�ƢI����᳋3h���D�ovV�� �r�Er�]�6��wөAǶfu�ޭ����J���GS��o��Đ���ano �U��xf�i��K <�f'�2�vDqe�׏	}��-�i08P���YӚIg����b�D&�=9i,/�:��V�7�;�ٛ�$��:��f�H�./!��&��Ws4e�5�p�ƻ�K
��Շ��ҴR2�($so��H�k2s�S���N��3RJ�z�S���Hӥ6��͹ۨ�ܬ�+������|s!�N�Ė݊ؗ-�-��s&g#yf:�����J�n`�(��u����9S�P��9�%�&A�$u+K�'qh����.��z�sj�ͷ̌�z�[cZIlqj��Ɋ0B�:�7��0]ܕ�%`���d�w�>>q����Ъ��TKUH��b���PX�����EU���)Z)t���V�Z�F�*"�(T�V#l�n7%EQ�[mB��R�֥b�fQ��R�hZ�D4�i��j1EV�Da�CM5E�&3Q\V���-�TS-�������խE�G(T�3&El��1��j�j��Z�aZ2.Z�"�Z"PQ�*ڥAj�iTP�)aR%���!Q�������3%V4�e�f\T�h�Vڲ��,�ж�KmKm�*����ҩl��u�*�*���+��%�
6Ȳ�e��KE���UE�r���ʔ�Ҭm��)eAJ��j����6�Ub��mFZԲ�cK��̶b,hR�
1���Z��Mfb5UR���5�km�l�`� I {�R��f�ބo'���r=�O:A�k��{�i�4,�޳��>nT�#9ۇ@l�ɢ.��$a�:*��Ssrw=��)uN����9f8]I�s|�\^V;�J��D��}��+T'�:��b�-vN�:����*[;�=�Jf�Rf��No%�z22�*�SE�CVPN�����]�oP��Pu�@䳂���ɖ�Oz�T�)ؓqλ�xo�Jd���O�^��+��ҙ�:==�����B�h�N�Rw���m]ٽ�{����P��M �6���=>���5�����5$6주֎��~w/���6�9� -Cn��5+���O��c)c��yѽ�����`zu�ep���C�A̙��eej������՜��=g�U5R�Tf�&;\�ME6
�C�������z4�V9�4uEr��b��϶���z+���|)�Z-���:���f��wɹ��y8׾�'��֮��>�^.��սN3|��ހA�Nv�u�H��w2����4����X:�2�<C�K����+��A�a�<龍\�,�U�RueB6C��1����'�UͲ�v�3MmC�Wǲ�k�Zu�-=�.젷;*�F)��f�9��;A�`b#_t�d:�.�N�i�+\�Ol�{���
�����P�Ԣ�G+��f��ҽիg/�cdT�y����YMz;���	x6w>�=�8[g�į;h�"��C�}�hJ�yp{�2�}�~�=�*9z����M�.f_;�Ƽ�WN��,CǼF)Cn:���O2��o!W�ЫI����߱�f�6��UF�ۖqY��]s����k{܇w����Z��>��k/ءLRz����ͽx;*��=�Y���ɭW��HL`�4�	�R��p�E�Os����;�o{+�\3X:{�T[A4<sJs�T�{��t��VU���+�T�C���j�׷nC��:a+�^W��ɫ�����r�Ø��ƅ�/>����e�V�#SQ��G֕�-'uF2n�2�S�y-NOE'Uj7�'����J�/{�n�k&�y�<���{�SK���M���yP]C�@Lj ��C;�^���ՙ��\&r}��u�w:�nq-@��\���d&J�Q�t�����,����4:�%Yg%���X��*����g��
�aL�2��)[8ڈ�j�A�u���X/p�����I��]�k|kO�d|�[0Mbf�ޛW2��:��}����ʷ�b�����cz�Y����1$�nu����T�#n�W�w��p%���:�o�nW��r47$�:>6 Mm<�װ�d��=X���N]q�ϥMT:k8f{x�Y���jN�uX�z/�t��X����@���h��P�yLm���:?*��:ǽ\���8U3"�;��o�q�� ��I�5�`�.��G�m���ܺ�E��d�_N�RU�ԜVU�Nqc��_W��c-1��?B��=��^��M��ZJ�����O.*mF����}����*����Ϋ��e�����й����LS��n*#�$*1'J_;�"�^>�2���+i����I�X���s`p죒�u*:b��!������(`�S}=��{9L�ۈj;6��W�o4��c�����+Y'�q<ՇSL��yağ2�?}C��d��=���_tw�Q�����^б��	*(4/ûH�k>9�"v7�+s���u���u>��x"c��t����u��=}:���і1.z�׊ѭۑs�˄[r��;R}]K�p����ɝs�F�2,n�=Y�2Q.��(��w�M�˩�v�)(��]�M�hړ���{ �m{N?0���)Ğ�0�=�,'�M���%I=f�{�I�>d7i�+'�,5i�����,��f����_]}��FXN�au}��~�1&�d;/��|���<�� z����>x�c&v���&�i;�	�i�����XN��w��LAB|�B�|���b=��B;��:���v'���nc�{�C��Z�<N�����Y��8���́��l�p��Oz���:�d���'��N�x$���ڒD@=O3�V������F�}o5j�D�8ʒ�i'�N'p���z���Y'S[��%|d5�8�Ԟ�0��a�����2u�l<@���M�z����b=���5�8"��~O**�緭���Y'�v{�ړ��_�T�2�k)8��'Ν���@�?!�XO�y�I_���	��=��u$�yL����:dA�]s��sw�G>��&�Y��'�x�~�d�a�����RM{x��}���Rq��N�vj����?P��	�?R�M!������Y�_��>�?nՑS�����#�0����m����d*d��;�!Rxɠ�h�$����W�$�ϲE����Rq�䟟��N0:�CCDz�y���gb�_m;����-��}��6����8�1�w�8��15�0�'X�p<IĞ�����'��￴m��'۲Wl����0=-���`��I�U�r�m����JD!��!��z�Y6é?y`x�d��<�	<C�}�:��1=�u��M��'�8��T?N� z��'~�|�i���#��E[C�U�R�����1���I���a�	�������Bm<f2q�R{��4��s��'�8��y���I�?C���N%Bw�?$�'�Rr�}����i}!�C����Fn�t]���٘����K� YnU�-5��y`��tA~꺴��m<{6�c"]�R��;c�[O�d�_e*48��h�Z��&��4��2���_-�1�u�m)�wN�Ti�x�Pm�"�-�&:�.���\�/<F���v��0�n:�[=�ef�J�끙�K�^}c�����f'\a:�?XO�̛M�gY'�Y�:��Ow�4��M��x�Y:��y�	�N!�Y��$��>�d��	ξ���f���Ӿ�.��p��>dߴ����'�=w�h���w��ěI�*��N�g'�T�n�Y&���Ad�ﰊN$�*ny�	ĝa���~���z�8}~�ﳼ~s�&�OXt�a�O�O����N������uĞ?No����06r�̬�a��d<M2q7��I�M�P�$�{��N�`y�_�;�?8ܿ���x�.�mU��O��#�#�=S��d�����~I:���d�N>0��:d�x�����:�u7�oRT�H(z����y2��d�o)���!���g����T�ӛ�'+g�C̓ơ�'�X��I�NyC��2Ad��}a1&���ԟ<a?Ozd���&�;�P�����ޤĜHl�u
=�" �'8��U��|N�Ҍ�ڿ�P�'�SOx�5a�i�|�(u��� �C��d��v�,�a��s��7��Ԟ�$�&��	8�d��k�G��=fMⲰa�����O���Z�ϢT'�+'�,:Zz�����M�>M0�f򇬝2�`q��<~C����6s���O4ɗ�Ǿc����E)A��^�2�l�V.��|$�m��od�!��~�*
G�u
��VML�q'�>f�,':�݇�I8���'������I�Af==Q�%��\�j�+���B�c'䟐;�p�f�=a���p'P�'sX$���'XVO��xe�=d�Tެ'=M�:��kvB�4{Ј|4�7\�}�GU/��?F�'�t���N�y��>I���!P�'�,�{�C�M���	ԛ/7�*T�G��+'��
��OY;�{4}c�Cع�q�ԡ���D��]n�Y]ہjMm!��� 㾻9}˽��9���T�Y��8����[s�/%�I���5�Sk{q+�t���y����l�j�=��ƚQ��Y�%N�ӹ��W�=����)Y�����F�SGt��ݹG��u�ܤ�\��K�O�Xb=�"?y�CI^����g̓���q�Y'>�4��)��
�<Af�{�*Ok������?^~ԕ+	��'��>��k�@��M��������y��Bq�vn;2~d�0?3��C�=βLJ�_{�Y&:��:��)��B��O���a
�Ě�jm���<;dNY��m�w�.��#�{�>����N��+08�o��N��'Y6��?O��N��>ΰ��Xl��:��14��|���h~a�O�v�����l�J�]\��q�"=c������4ɿ�d���q6}dR~|`j��$�����l8�h�<M2u'~���d��މ?!���è,'�w׾]��9��~����ጟ%d9��<d��'{́�'̛�w�ےc&矰�8�u7��I��&ٳ,�$�*jnì8�jn�3I8������:��w����y���s�{�־��]���|��;�a�m$�ӝÌ�J�w�u���>$����'�=y��I����O\d�'S�e��m7�q�x�4nÈ)'=��=���������y����$�
�Y>C�N%g}��N���a�m����ì�>0���:�ԟ>���`x���o��<`l�%d�O�,��i�����w�N+���g݀\�Z���c��{�F�RL5}C�N�`n~���'�a���:������:���ì�|a?CΙ�>��w�'Y'��kz���$���P*��G��/�}D�1��ǎ!�Os)�'P�1 ��>��'�X��a�N>!�� �q���d�a��aԟ<I?CΙ�<}I������{�Y��{�&�x�{�#���IXq�ݡ�T� �դ>C�N�̦0�$�bf$�5�>J�ߴ8��'_����4o���I�>n`W�^��_�1g���@\+��R��p���u9[v�o�@��낦�QNU��l��nBke���^��q��F�F9�ʾ۱:��ޫ�}�oLZ��'�*�3�w�V�����<�N�	(�'jj�[;���(����D������ɜy�Nu��i<|d�����N��M��څd�&���%AB|�!R|���l�����ad�$�kt>f�N2��O��<��b"�!� �t|#3s�~�2&�f��������z�$ě��I��'�o�	�6��o!XN���Ԙ�����!Y>Jɬ�q���&�O�u5gЉ��ǥ���덜s[��}N~�c��će�'�����������O�<@��rN&�=I���0'P�&�����w��J����J��VO�)ǣ���	��H�ĵ�S��x��'��N�X}l��kt8��2<�'XI��L��u�s��4��09�N�I<Ag���2^�a:���z��=��3'(g3��}v��s�#ӉY:I�'��t��|��y?P��I�?!ĕ��L=?y�LgP��2~a�Iô�N �=��B��OY��1�Dp���6����|r����&���8����J��sgrE���������lՐ�����Co�'���u�L<��q$�T5��:ì&�|�db �Sߥ'��P���=8qk�s�EC�M%C�|�
��M}��6�:��9�$����>�O���$��xj�q��T4��l8�����4�����z=� ��r���̕���߈�g�i$���p�'�)ϻ�Ĝd�+�y�+4w����i���.쓏�ԊOόKa�R~|O�T6��&�1�({�C�#���#-���j�O������{I?!���8��z��ܝI�VCg|��O�=J�����zɾ��_2M2l���N&��"���&�r}z=��=�E'פ��9�w�ah�G�?0��<M2q�g��u'�.��~C�7=�M�OY�sܝI�VCp�u��������z��M�w��a=��1�#��D��i�!}��F���x�n�0�R����0���Y���u1c+DW۸�)uE8�B��˾}f���<�DN3X��I�)p�!	kr�[4"�yA��c�Do�̑{�IP�1�A]�gcL�&a�>��)����ޫ���؉g�I�S�3Q�7�o#|���~��'8��P�$��5�0�	���d�'��'R��XOXq��O�L��9=�N�s�	�i�N�z�#�>������$,���r�	�_{�~����NRu��a������Vu��
�nÈ)&���N��x}�B��'���Bq�Xo�ï̓�1����z}讇�P�#)��U��m�$I�O;;�$���O_���h�'��|��d<f�q��q�z�Sz��	��q'YX�̅I�N%b�Ͻ {�z�0�⤂�@�}y9�׵���p��I�Z|����w$������jN0�g�����:�X|���
C�<I�V�O�pՇSL��q'��y臙LA�T�,�}4���C�[��M�q�>�P8�M��XLd���u'�O����&������g=ޤ�2-:�d���!����.`��C�ǖ���"��=��Zg~�k��q8�<kY9�!��:���<���P���|��M����'�O��B|�d���V�zw��LABh>��� ����ݽ��Neӭw~����o�z���N�Y'�=f��|�I���=d�Cw�2q'��<3��P����Ğ$���$�m��O��B|ͤ�w��N������;���u����=��7�1	��J��T��Rz������F�u����v������':���C9��OO�<��M��{�=� x�l��DV}��Zv��{��Bq��Ϸ�Y'�l>��I�RM}x�������'��:|Մ�����|�A�I_=��&'Xts���G��*�x�إ�Ơ�Z�����}oLd��h;�B��OY�wuY6gw�l��o$�RO=�IY>�`ne'=d�f�N0>M��0�a��H/Y4���ڷ�y�����跨۝���R�t�k���ϥ�%�c�i��rrft}p�8,��H,ݠ=�ˡ{:����Ex��-��g�7�����̂���COEt�{	�E�uk	tBW��@k�O���%}mn��MV��/�e��;��Ux#����?����I�X=�I�	����l�A`o��T8��7;�!Rxɣ���l��?��W�$���d������'�?>&!8��{���}�7y�O��|w�|7}����:x�Ğ��,L�Cg��̓P���q�bj}�:��{C�N$�{�!Rxɣ��ѶL���I_̓�=����y���;�s��퟿w�:�?{��}�� z�ǌ�m����O�M��'����'_>����{N��LNs�:��T'{g�I�*��@���M����I4����7[��o���?~�{��%0�N�Y���0������[���'Xu'�,���N ��xI�!�,�i�x�C���N%Bo�d�'=��3�~}��ߝ�q��;{y-X_�,{�=��=�茎ُz�	����~~d�Vu�x���ԜBkw�4��M��O�'P]�7�y�
��E�{�=s��B ����U�}�FT��)�H��C���!�!�v�����=d�'�����OX��i'�xe	�i�������TѺAd��p:��O�R)8����N~�Ů8{�_o]��_��Ϟ�zԞ���a��	���q�������N�������:��O_ӛ��+'��̬�a��!�i����2OP�l� �K��~���{J{�}�n��o�{��q�iX=���N���w$N���p��I��u'�'�t�$����{�u��o�ޤ�:�ݡ�+'�<Cs,��N'>~��wm��ȝؽ�c���D1EBC��ve2u+GﰊN2s��9�'h�0��	�>�I�����'��O;��d���wz�q!vw�~�~�5�����͡Y8�ö��=M�1��'|��>|�C��?���8��(y=�H,�a�}�_�Ldٮ�Ԟ�$�&�;�$�m�9���w^��w7���� ��&��AOK�f�f���)��1��Ҡ�6�� ז����}(e�BZ[�����#3O��v���,�M�	�0��b}�Օg*��ܒ��Z���.<�� Pu`oq�4:[�Nc��;˷�5�M&�n�^�ZD-�7����cV���_�Y&��w��	��>B�|��@�ORu�RO�q5��L'P����%���I��g0��a���{�=��g�kD��_�R:3'r.�|���>d��Ow�u6��7��N��<����5��B�|��A�$�'����Mn�検f��z���Cpza�D|#��;�c%�w�;���No-(�zCNu�d�O�v���'�4��`N��M���$�9�5&%a4S�+'�Y4@�OY>�1��'�la�|�y��Y�2�W�]4���Fv��É+�C��'��?�6Ì���0�'�<@�l*�����$:�����@��I��z��I5��
����q��N���ǿj����ӿkO���������N3��|I<C�8������8�1+O�ì:�9��M$�
Cg{��q��o��'�5����Iԟ�����XN��|>��<�{�����o�sޑd�
��ORm�b�Y�ٷ�O̝C����d��{�d����� �L~�I��{aP���z>F=G�G�xW�*�����K߮���	�N��I_�'��dRx�@�X|��Oω�N2����I��?3:�ϳ�'�V��:��15�2>�G�*��4Lqc뺽�������s��a�'�:w�!Rxɮ{���4ɳ��%0�M�dR~|`j�&ަ�,6Ì&�OL�Iğ�,���N ��$�a�w��^W5�z��}����h��" ���!O1n�}�uG��j2��°M51Y*6��y�׭⽾�Sw��F�!�*�QUe�h<o1Vf(O7kL�y;`~�3��݉>�q[̋Y����٥��vv�ܬQ�Ȓ�K:�K�la�DGÂ
T�N@����wm�\�Ӄ��}�_T���Sê�Pe���ѱ�MH�ZU��y0&΋���b��ꍮ'-�Mgˤk���ms�5�Xx��O�/cfs8GF铊We�u2���Ǩ����wD��]۵LY�ك��UY����d�.�Ν @h�e.�%�oa��U*Ob/-{��L�E	������7��t}��//�J2ҙ�q�M�B�����bvng^/c���Υo/S��AV秨 Ÿ��r�����!qĤ�}V�ҳ�Jy����b����w���ҖU�R:���ջ�[}�`�ڴ�=�K����U=��O2U�}��.9c�
�;(.��q��-0��L۶Qj�mX���W�9Lt&`͝��n��2M�2��a\o~�ͧ�#���wZ�<e��8����t"a�#\����W,��u�V�'|m_YZӭ���2�R�/_4�)q�nn�}>6�e^ݙӒ�GR31� U�5��^�[�'s���Mg,t"��Q3�{kqg��敃)��M���w���׉&�O7+�V�p}���kU�S��:�別[���v,[%����]v�;뱭^�V_o>f��eZ7���l
�
nBGN�n�̭B�ٛa��O^�� Ul�0���5RJoI�"s�'�v�u���	�e�6�J����2�|��r��>݂!Ǔ�����!�wX�un�Y��ާ.l�$�Q�u�L]�o'ܩa�aZT6E�1d7jȽ�݂�OWXUڪW�N
2�O�����H{�vf��g�:���A���F�u�Į��z27V�d&�Ռ\#��uB��!3�<���Z~ʗ�jښ���닇P����2�-=AA�:�foR�V�GR�Ѳ�T���efZwg��C,С�jU�]j	�����z��D�C�Ʋ�(	skS��3��CX����_]�g�}��ەև��+�t.�M%�i�|)W"��R���jV��q�����<̟`!K�]a'Y���˒̡�2����F�W|�b�U�5�:lX�s��FQ�b��յ�w[ ���pY}2[����7���mZ au{�a�6C����d�)�X>����m��uͰ��u(M���^��4ZGՍ$�(�7}zW�x��y�Gn�}����k�9Jg)������o6f�R�l��-�v�B�j��ƓM�{3�DP��yy��i�XJ�5��,�� !T�9v�bW%���̸��%�%���:�
4c(��B�����x]-9�=���5�m�̴�R����#xT��eN�ۤhL�B�k���YՊ�x�m�����C��K��@���j&!6�_>y-+�v��.���pAQ�ݛJ�SW(�Φ
@dT������y�-���� �Ǧ�#��p�d��Y�jq����;��y�@�}�h��-'����?{��+�T�-�j5R�J5j�E�m������Q*"#VZТUKE
V(Ҋ���֣lKjZ��Z�*�Z���ص�"�B�EEJ5W�W+E(�#KZ���jYc-j���m��m��)QB�)m���Ts�ciUՊ,kTPh�e�,X�X�(�jVШ�lB���)TX�k�[Bԥ������ЩZ[VҔj6�´V[A-���kkj´�6(�A���-K(�-iQ�QRֲ��*�m�mF�l��Um�j!KZ�Z��\�ij(5�lQ�E�[im��+j*,��m�m
�1jS)GZ�QQ�Q��J�Z�U��)EF�V��B�R�TcR����Z�5���[���[km��AE�#�*�����Jب����[J9���b(ԩicmmZ��KA�U�KF��h��#S0���TE��[X��ԭeUH�m��
V��D%h��w��O%�3��	�:/�,73�Û���*N{ƸHl�܈-�8<�६��f�E��Y�A��^f��  �2�-�۩����{���}�.���~m��v�oʯ)!8���t^3�f�:�қI��N�B�/�!Qi:�R����8��m�S��\э-�v���r�������
T%��Pm>�W��b��I�_*��}�����بܦ���:�ýڳ��K��rOk���hR%�3+�T�a
R\��̄�uFK:ǣ#x���oP{\f��'�V=�3gh;�\5mc窽o����̽�J�bcB��:h.�#a�i����>��(�n'��Vr�W�MV��u^�5
��#a�soӑ��Hߝn	��{�Mc���+�Nk{�⭫�r�79�~.���b�Ez�j��,�&�/g���R�}u�Qlm^"�S�T6:�Lާ�tx����C�������V�;6�#��o�w�O7R���缡�b�8E,\�_3+��1K'���T�'SG�s�U)���9Sʼ��k_{#p�.'�(����ꎓ�Nnӊ���{�3ݶwWKF\G!]YRu��
�K�g/j-\���!8B2�t�գ�	�M,h)(4�s�!!V��*���OU���_��D{�(���r?CCps���T)�tu�]yq(�^}+-z�H:>mN��b��n���a���h��=�������ȚM��&��O.��mRqZ��Ǳ��q���O3�[{���+
�Ν��P�0�	!2{B�ڳտ:2ijs��Z��+�N�9�Kxt���^G+;��K�-R��nb+�Ez/�d�S;Q}�~~�V@^zI�s��'K��p���7,>�P}:�Tv�{h�v��G_a��ܕs�:Wg%jI�m5����ߡU�:�䪂u�J���G`H=��}<x�cv�m�:ɋ~|Ӹe�p�n#^$���{���\�]���V3xϪ�nQ�3{=�Jsq=�z�A������Ƶ��;��ՠ��'�5��^�[�Տy��f�5��;�=��z�#Q/:����A��0���3h�MЬ�^�'�>�5,����b�,B�/��p�/��\��L�S�{�ulM1��Rge^>vKU2Vo+�6��r�)_Lme�Z���T�\Y�7���j�b̒�M�/6�j��e{]a�b�hR��xɔ���-�j9�9d�Ir3�`�/��DDU�N��O���Vux�9�b��xrY�V:�'�7=�l�>���՜ݜy�(�s2�:
����v�4�����>��n^m��X��Z�����&��gg�]Jb���y�g�juK�T���CR��U^V����7~�q�݀��X�k��1�ܳ�Mg�d�]�-���p-W�s^����s[�LBi�N�W�"�����:���؂�j��뗙mZ�n��ǚ���pf95�����{u=B�;�edt���v�[���;ۉ���N��*+;Gs�����h�5�v��;�t�8L�\�e$���K���/'õVҚ�n�6TVU���n�=vz�2�Q�cN�OK݅so�ZZ�?���Õ���m�{+��XEIȧn,յҊk�mk��;�ێy�:fŖ��u�ؑ��XOxg�W�;������'�u:�nU��*F��a�+]�ǅ^�Q���k���� cn'B�#{��<��`�8��5� �Ġ��!qK�W�C�mV�ƍF�f>C2�K��]Hj��v��Z:R���^v�O%�z=���sj9�c���^s�5M��$���e��;My�W4�z}���'3z�[�ˆ�4��8�P����A����m�Nh:�Ѹ9E^0��^f���]����$ە=P_�j�1B��'�����F;�gr�Za���ۋ5��)���`=tO*�����w���=�[޺��z-�p��.����:�1�dP�tQ��k�Y,rW�V0t�rq�̻�}ς��o��9��%�ǥ�[�M.�a�Ox|��X�}k�P���Ou�)x����_����o�bS�O#_l:hٴ���g����u4ްy����o����_��`	&0�ug��������g��w��R�*߱�8��l��*)����KwO,����/��6�[���;���ܝ�ˉJ�)fc��dLv�3�ME6
9��j��Pq��sF��4��n��1�'�g�vإ�=�9�X�n��<�^Cr��]���" ��D47J�á�V=�p�ujt�3B��nܝZ�ڕ���%D�n��&e�T/���0���1띆գLM�*%�EgN\�s��UU}_CY/wkj�O�]NЧ�sy��8�\vK�x6#��ѕ82tf�Fac�.I��+�	YY.:Ů��R�R�d�y���y�j�d�]E�螙T�xX7��OR�۸�sU�ue�E�T�b� t�d\��˽�by�Wѩ8�er��H�;�{��7ڒ}���7�'���^0?�T��"7#�����'���L-���^���$�s�K�������M�zִV�^&�\��<���N�2��E�h���Tָf��e�:�s�>�Qs(��F�x�tN�㲗	����B���Վ���3;��{9��ۆ��n5��n�����O*�s��L_$��RX���4enk�D�v�%vm�nS񸽗J�\�?*;6g/�)�N�ث-*�{K�I�����[�j[W2�>�~�=�:��q�f�	�ȴ���3��_޷�CΞ�E��[�g�^A6cU�-+��1Y�G��T:��F�#��wJ*y�����!Gx��;-�+M�=�A���h*����.v��9f>����S���9iZk�;{��\\/���wȅ;Tڼ�EM�/�=�Dz6s�O?˦���_�����|��.��Gx�<��r��$�:��oo�ƫE)���]���7�e�>�k)>�U�a�˄�l�mE�]+ci�9��N��5��w95أ�s��>ΧЏGrp�F�d���*x������k<ߥP����G��[诛�s��c ��YY��Bg��]lTrCC&<�ӿ+�:��u��T�*ob_oUF �V�*������β��r�O�X�*!�X'�Z�LZ��ږ�w���#5���|�G�j���:rΧ��^��Q��ikB�Q�������Z����++�ԁ�V� �sؤ�}QNk%E^54�ڝjւx��B��m�m6v�2�.yyX��E/6�)�A�A�pb�п=�6����$�CgJ�|�HM}�/{J��s�n]�b��⣰$+ؓ.\,��^]ME_�1]06�pިo%93Z�Ѝ+q�����L��.��nЉ�}ݸ����!Y����\o�j���S���d�p鵽7j���]�*���9/UN�d�yk��P���p����v�Pnn���Ah�ɋ:W��}_@Ya}ҘBM�̮�if�;{�h-�ò�J�uץGLRa,0�m;��Uo��$U�Л|�{�#,���J��è:&j�u)�%n�X�+=.�d�9K�!>�M�{\9��k��v;Kh�D:&;�;	�i����R��J�B.��/��$�5�|�Kι�7�Z�5��*�!�ӂ�\�n�yOa�AC�U�\z��K8+|�,ܦ�g`[���f�p�x��y�j�W
�ى�C����5�}}�ˤ��*Tj��t)(k������!f�U�~��T��<� ��"%l���1 ���&�Q̜[:^K��r�bI�(ܰzɬ��+\���;��gj��2w���M$���^��֙NTo���)���ӵb�pۮ�5�Esv�oޘ��y킧S~���Y���=ɨ�y�Z-��jf��CK��.�z)D}=��+��W��C�J�6 Y�Y��oF���|'pı�uj6;����1R�:ed�Mdwق�ٳ;��9Lr�v��ݹ��q�fo^k�]ݥNff�F�nS'����nP ��BMq�=�x��iY�K(,v��Y�+w
�遼���ޏD]����n}-��.i�9[���;w83參v�&�Z�|g���I�wvھ�����|������6TW��V�[�U��E�+��C�+9C�	��f��.��{���޳�>s�����*h�d�쉉��$�4ѴN�*m�im�o�!޶j��׬j4{G+�ާ��� �n�݋o��.�\���MQ�3o@�y����6ʮ��~8���\er^���ٳ�-�z�^Jq=w������{�����_��e�$��3|����7f��(ݾk�V��(�A\/���	E'��9�W��N���F��ނ���k:w��䷟յ�M����d�Ձu.�H7e_�k��M�[�lu�v9��D�-b9O1��v.U�l�5�tjn�c<RpN��']Xs[X����:|f��G��Pۊ�̳��^�Aͷ]���QN�T�H��s0e>��.��y(����	�i����rMp���	�t��$�{5�w��l���P鶣2�Kj�c���k��A�- c�V˦�t�T����V�y؀m�1���������k)��;�}��{��yT�<
���n<Y�PN������jBxD�$��3��g�P�����Wv1��\��׌)}�Oe�'�أ�̐�`�V�Ѽ^�9��KϮzvM��l�+���FÍ��#_fȬ9QP��ld��'qZĻ��WZ&�{�!���O86�2�b�Po�޹X=���Pf95M�f^��������g��\��yZʜw6<�j�U��Ƣ�)�gw�ִ)f���z�N��Mh�sš�z��z�,����T�VVKAA��&u�{M��	���8c���%U^���35=��ݪ��y���Gݦ1��p�T^>��W*��Y~�Я/y�Ŷk���3�]ʇL���b�[̶̤��	�'Z����/i:�.��}����f^L!���ʞ�R�>U���nP\3ԠΦ*;B�|��"�K�]�6�x_=�����5r�ևJ��)o&p�9�ߗ�N��u���ʛ3��YN�-�ʽ�X�7����Y�kd��p)�-�w��)wZr�v��"�P7��ilp�8��9k0ڊ4�+E���gtT�X��-Э�-#�q7y��FLȎYF�.�#ޏz#
���i.f�s>�݌�X4nQR��u�4�LE�5��)F��	��8E��u5��) ����J�,�v9�
4l?�PO*�u�.�ޱ^��T~��}��s�O����3S�3}�k,����E��1��ٴ�kU���7�o�j~��t7�f�j-�5-�����IXu�by�kͯIFO�Kk�gw�S{/��ƾ�PVLr�y��l�r�½K*r2r�]� �oZ��}�����Pu3��ɀ'G�����J�aC�c:ã�9JVG�?E�ܝ9]qkK���'Iϗ��8߆��L<%�ӗ�O�B(0l]��d��"zp����.%q�l�l�KB�X)v�u\a�����Nۿ�$��i��ѱ,�:\�͘�!]�sG�,�Ĵ&��5P��Ȣ�c��׻��'�i-FE���Xķ`�Zd��3ˎ+����� �9֡Ϫ�z��U���o�����bv�јi�&���v�Ŋ}�1|�	}�1��f��fj�]���mX��xJ3�R �Wf�)�����O�����9͘�wi=u�H��=]H]�s�gz���f��6�c��Xo1��Kt��i�\ސ:*�������x/�p�Z�/1�5�'hE�/4�t�Lᶷ%gR�\���s�:Q��؄5z+�<��;���AL�*[7Ps8�7���.n��V�p�L��q\C>ԁ�<��`���h v��9:��h�3�y�����Nn��ǚL��&�Wk.�����g�N��r%CQ:7����f��niv�t����uJ����i���,�Ha��n�s-P�[p�$��a�^"��\;�=	!ڐ}Y�f�H����.ER�9u�ח��uC���]�<��6�UҰ��`��h�x�6����ٻN�*�.����5��oq�-�	K �fG�¤c,Wq�����[O)m�n�vv��gu*�I�蔳�g����'�(�q����5���\l�
�rm[�U9@S����C�-m9;�nΣ�r��!�)�U%s6.3�WG.ƎWR��R��U�ar�ĭe��d��Y>�f�4�H��ռ`�eVX�GY�Wc*���6�u�h�Ŷ������}GrN���>g��F�_,]tlC�����We�|k���/�GE�*��s��3zj%���v�a���Ի���Ӆgͫ�)�Pq��X���+��#prh
b�瓫e��7����5�3�luf���S���ڰ�Ȏ��������b{,(/4����zJ�}�/�����S�Xk��WdT�>m#]�K�Hp��ݪ��7_v�ԁ���]ֺ���*�nA�Ʉ����b����N�=R�4r�{�D7��ەɺ��6�;)\z�I��i7X�nwZ����shj���G�v|���PeA[L�I%��e�����Zev��I�͈��d{f&�0p��1�{S�s�\��t�nmp��wo1�l9�ԓ�]�36�!� v��U�)>�X�l�ֵ����=RZ�'�� W�%N7ݫdL� ̔r෹���o�*�*Ҽ�;�*�pG��ڙ\�$�*�Z�A�ʳX�f<1��xi��u�2��;{n�N{¬ �F�7Nu"��d�w\�pt����.I��b����'�E.�lx��0�V.7"]/��UY *��Z0�G�`o{���s3F�Zu�P��E[|�B�ŏ^n������T	�A N�#S�c%��֝Xh��;��ٽ���48[-M����S���=KI5�����v2��DeXͺ��N��`��4�	���щ)���X;7��:T���v�)�VJ������B����p�}���$���,;�7��7���t�x��uŷx�Ո@�n��&�8*t\����7��u��oM���0<��>��+���*ëЧT�p�s<ߞ.}�����}����Q�"1���mm�V�
��B�lb�-�*1b"(�VX#��խ�m�ҍ�J����F�UTѣU���V�" ���F1EkV��(�F()����QT�iU�ȋm�����U���L���--D�U��"�#Q�[[kZ�X�J�)JU�"�)l��j6�`����#F��Q��E�A*��bEF��є�cQ\J)j�eF%�%b"1UQ���h1�T�X,�Q*ՍeQDF9h1QTX��
$DZ�"�*Ԫ �R�eJV�%j�P��EbRʢ�V҈�Ԩ��[k
ؤUX2ڨ�+UTUb2���V"�VT�EDJ�1�(*�V
 ��6�Ԫ���U��DQUF"[X�Ŵ�D-Z��kF��[U--J��Z�U-�j[h������b���[-*
�(�Z�UP�V�jU�����,Z�Eb,���PX�-+h
����V-lX�o�����l����7�6��r
�u&oKtk戳[��owX��W��q�J�I,�:�����4d�D	���)�w��  :���ɕ]+�s:��?����+��ά#v
��/�����Z����T>κ���v	̤�w�5a�m��&������c���*�s�V���e�66F_ݎqB��/us�.��#Cj��o�;�!ŏ@`vZǃ֮]c��2������o�]�2�c��8���MG.��%�����c��J{v_�K�_�0��M<WK��j���Y�h����z�u��QZ�v�ƍ~uM1˨�q�R����uvC��U�DP�=�6�猣C&0�ڒ�uQ��f�:BIy�Qf��W�|X�.����wh �`�/�IDP(s3�	9�/ >���Fk�w�����]
dS����ۣc�;���(q��Tm�۹����I�R��J�]��Q�^>�PZy�|��Cm�镅���ț�Z�Q�3G_&�N!�nWZ�@G?s����(��bPvQ.��Ǖ,=��C��ph���Om��{;�go�\�Z����� E������+:�����9��Jg�Q��7<s9�uL��V��5�ӊ�ZY���QV�=)��7��ļ���gf����:�4^���s��u����m������VOY���=6v��r�W�ok��.�t�-n����g0R�O��c���.Y���K�{��D��%c�*T����k�2'��qÖ*]��̴*��:G�uϛ����.�q���O(����~}fϻVr�kk��;BCL�0���ݘOY�s��m�K�G=P
�BU���/2�����+ۍ�Q����I1�P��]�7%.X.F��Y'|p��W<5T9�z� "C+*�tuE���$���IP��D�ю�^�NKʞ�"
{���U{��q�ܶ���T�8U�4׊�^\�B��Z��O��,�ݖM>�	 �ʩ��T��]��_X-���TW{r�ӥ�p�(��-�͚
.6�Ǚ5S���@�ŪBFH���mYv����\3˕KU^4�p'=��������(t�����/ws�]�wlb�xk�;�Z׎�;����ob�D����q�d����萢�G���- ���{F.W�q����:]-,0�jyl{mU��p�M,��فO;g��^�wOk
JE������t�t�z�@H�!��o���i�k��p*��׋�'MQ{ԅ��̴��"�]�#l��.i�D���E�F� �<�Ɇ�EMɆ#�Zs��K�@e���h����ݞ<��g��CZ�3ڮ�ڇ7;�u$�Ǥv�ca�8�N�Qg;��"z����e뫙b^L���
ɜD�Z�����]���{x�����=��.h;�3�˙fZ$V(�Xn1H
���=��e�+�n"�c�/��t�=p*����zx���L�WR��r�a��1Wy��):��5D��y�����0�;��o<�K�w2]�C��i.�"�[�=g���iH��C,c�<�άd���)��[�t�Ke�B� 1^ǂ��H�g0�,��f��2t���d\hT����v(���(;[5���LT0�H��)jMyj�'=�1������GR�Yʽ,k��VS���W\����c����^$bj�RÄ�!˔�]R�ڒ��c��.!��ūE'IxhB�_�x�U�4K����:�ے# ^���E�K�W��Hr�[S��~k.���K

�R�nER¶�X��o<�9���ғ}�xe,�܀D��lN�*!9#+��\U�;(���N���UB0<��X��Ă�W��踲5+{&�⼼T��h��Y�ZM��"%����P�:Fl��̧������󽆯�����ԗܥ��V���5yE�Qͽ�m���H��\I�*U;:�Q���ܢ�Z�|�΅l��eZ���#�an��ɠԦ�$���(c��j����y ;;7�Z�U�l�B�����Gd�n	�m�7j�v\�Ѓ>k&N�������Ny�뒮8}�Qqq�Q��@�s�>J�c㻑�:X�Zh�=~ta�i��=x��t=�{:4m�i��8��.���67��c<�.I����]yXs@S�V`�y|/�4�K��]��wV�S�h�1y`.��	��!l�`�(;�N�B.���6{H����b篏�m�Y�⋳WR�#�L��x��q3����:�+2���@K��e)�ib�Sy0��f1�wk�����du.
T2U@t�D�;˺�wu��w��Yz��O�Nc�7�6�� �ͯ���Q�akMh--#�Do&lno>7��]����J��tp[��a{��\��1���ġ��yd!q�P	�������kz%{/��<��[Hc�yZ��]�F�W"�NX���q�o�`�/]сY�)2���J�Ϳ{;^'Ԕ�R��S�B42z�ڇؼ+k�����'4(�(С޿,��ўw��J,1�&EA�"8���sK�r��洛�q��䬦@uLj6��[(ґ�ޛ��g�� Ί$I����͊����Cz!��i��?������(a���Z]E����@�x����{�BL��L�hʕ�N��/J�IK�Y�gpa�+\8�!Q���3����/l�.�NA�:�wB��=r��Ͼ�G����ֳ����Y(@鉇
��Y�pZK��G���5ژxO��Ɯ�ta���A��3�pKٻ�T5K��U�Nq[�`�!�%Q���b_�Eo�+��� �{/i����[I�v{���3�x���b�/�f��p.C]�_Ӛ94a�Zv���㷔{w`�����ճ�[0����H��7�O��V�j��{�LOB�j��7欍�:�X��,]��8O�����SL�׃�������jgV�`��+�Y�R�b�M�kf��U1ӎI��ߙ�o�R���:u��/���/)�7��"8��϶6FvT�Q�ϻmх�Y�l�բ2�ؗ�+�X�z�˪���'R/�g��쮉c�3��%A���U�_�\\iz���B�G7k ��w}/�ni���y��P��p!
�N�TOfo"�;�p�1C,a}QÜnj�ê1�~�����	~�0�\k�X�ƥ�J���~�tKy7v7�%�H��x"f;$���A�a;���n��sbPpT�E���Q���s��S��'&c�VS�G�:l�ӧZ˔����!��u~�M	��� ܽ�<�uܩO� &>87'ox��Ԫ+�<ȕ���pX��sb��4<�2�ov>���p�� d�qb��ə���7P)5�u���G�ެ��(v�a	�e����/J`=ő�\�7��y!��})bN�yE0�>�������}���X>���/�<�և��}2�Æ?�oxU���^j��FM�����r��M�lk]����v�z�Z]Zy�`���H�;�ַEs�0\�ߎ�g�z�������:�O����ˏ�B��"��Z��ء\u�u����o�0%�U�p,
6��vW�8.������"x��9u.��#D�l��0)M=S0��K��q��U<�I�(;�F}�1E�U�7��}��g�a�R��`�*�b��b�W;oJ�7gu�C��^X��M���Io(BΗj�rQؿ7Dh�u,H�Y�wJ[�y����H ~�]Ѽ�p�ks��%�|�ecP�lt�큊tc��_/%@��s��4��?{�����D����><��;^���������	�ĄU�䍜9��H5��7=���u�y漡��{R��5���R)x���"w���Mi�����j�r��O�~2C�_�[N�y<��y�5�]ƽ��2�<]��|ço{ R�o���(1
�7o��:�DM�&:y���Pvc�͙q=QF���0kJ�i��S�l޴6�$�9pmvq��J7˵���.�1���y6w������rS䰰{�X����VE�ڦ©�O.U-G׏�=���u�J���i��/��Y��$\V]pW�Vtd"��q]1�pf�tl��,gŢj�ZS�:��{5�>:��)��yEb����p��KN2���yl{mU��f+��u�#p�ࢺ�SC�<�P�$��:k�X�OqW� ɴ%�Q�,�q�Z�f��ގ��Չ�1�V���{v�'��7�SA�x-�uA�#b1D�È����]�Ւz�g�yOu��ڤ���'
�+<X�Q�Ę��N�M�B��E�+���$U*RΜ.:�X����7��-��[.)�Y��ŅK%�;�d�@�x���R�
��z�0r��9Ҧ�Rg��`R�DfO�����3�.G�M���h�g��%� ���
�gK]y
��=��i�5���S�wǝ1�|]h�p�Y��ֱ�p��;�E��c��*�/�Bi�z�v�D����F�P�.x��n,����<��)5�r15D��pײ���tw2��g^8q} �P\:�#F�b�@��.�r���O���5�����j���@+[���^M�}k�u��M����3�5��&o���j.�n������.Z��S����
b�c�q	P3hn�nj
��_/���G��C�mަ&�P��]{I	ゖ��uE�����9�k�Xa_��P�(�1c��=u��?ow��0>��NK.���YD�.��^Z/.��J�w
���^y�n]�*t) 	|Ju�Ǌ(	q�H�BQ%�ԏ��y�v7�y��K�7�P����O
Μx�A��Z퓍��W:��#���B��B�8�p�緦��Ekk�L��~��ر��k�~/����t�T�}fv�C6OGe�b78:�D�ݤ;��p���#}��!�m�t榅�U<�v�{��E�NgC&҇/�ߖ��67��l{E�OJ���ۆR��H%=����X̍����h�5.�3�l�K��j��WKdZ����(;�Wt���Ce�r��o�J��J|�N��yM��(�����)��Ҙ��k��#}��Kҡ	�y�e�k�m�*�O�pFJ�}⻱U�\Jޜ�����D�
�
J Ƽ�p.��.����&2D�"�w{zI�CSJ�v�41Х����V��s�!Z�#Mh,%�s�"7�ɿrx���}��	.�ԩ{»�Vk��m5֘�o"G�c�go:K��Y�;�x�uoD�B���Dr�d.��-*a��h��L�N�ݯj�tsm�v��Vԙ�p��Jv6_A�݋3��[����(o@�X)�h9W��~%����{��NEv+��t�F}ԉ�se�7��D3n�H+���Z<ld��c�.F��a\�\[�љr^�� cQ�0����zR+N�T[�r.��7N�l�%����ZV��MQ�{y�k�@ϧ�D�㼰P\C҇y������<e�����R�L��Я��[rN�y֠�a��:e�/$��W�:�� )��pP�^��J�ajã�Q﹃bi�{qo���Y����`5#a�r�Iq�I�]Zc��:�ac��os�u}����z�w��N�Gg�Z�,�ț�F��!��"��bh[k �ڱ�|aW�t�m�'��ɥ�p�������n^JEײtLٍp.C]�X�8�Yf�m���VK����J�pF�L\����C_7��xjƃ��%{����3ˆ�j��O����l�
 �|�ݻ�I�FA(ڏ�����/�{�jz�DWs��Z���u&p`KMьD�������tl��1���X��ƪ[Mr��q�s�%Z��>��zV��Y~�V-�^uG=՗ea�l{���L�s����]�,Un��fr/u_��u
pU��Lz��=NY�.,����v�[B���97�K�(T��;���up�*J��w�3���T$,;:��PY �D��l�7�g2��Yѣr��T���#�_z=��B��6܄�y������7���~���,\a�E�>���_M��)�;\��W��=w(��۔�������lc��d~�yg�E�;>�������7+��s��i��^r5n�d�[p����� ��҃�R�0^5KOo�S��0�ٝ���C��|�;z���a=d���`!P���\��>��y� �ı�5��^f�O��p��~�IamL��W��e��r���� �#�p��$������#2�1�l�{��Pԏ
�]�1|��Cm�镟p�.oxS�G/H��ӧַ}'/+�mA�dD���h<����OX�\c\�wZG�U,=:��ڑ�+�݇FN7��@���^8}r]�~Z���#aZ���ص�p]D���P�1+����w��)H�p�kڲ����:!�8GE:g,T�'��-+e-)Ҙ����/T��C��W�yo���G�=jN��1#uM�
ea�6&����ƗUA��I_z����e�W��K����N|EՒK
B����ٚ)�/~|J��i�d�i֎�)���n�������u��t'��u�|�� q�P�;jY���#C�-^������� �LŅ�v˱�ǳ��m<��V�rPL&�>��J�]Zֶ����1�j����Q��ϒN:�������oc�z���Z��d��1%��Tw�K�[��졝M�&f[��cSr�YF�'h�d����u6ۙr�oԤ�*�OJ��t}�tU��S��16�ھlm��n���VQ�ϵ,��uWFc�C7�Zko��"�]�ɴuD�e�7��!�t��ݢ�H�K�\7K��
��-�s5]�1rݖ»B39���Chv�u�Qxn����cG �ӽ-��G��&͌����W٫ �k8%l`���aCڸ7L�	���۳-�۱�.��� w�3�ʚo���M�ݻ+�^Q�s�|�"3��5�	(����#���-%�2�y�ӭ�D��V��h�����r�C���ǔX1m1�,`�P�I_+�[eqz�]�6��pfg77�-7MwZ���6�LhI֕K�4����9�L&�����8��/��j�G��%W,-:�ݬG�c���aB`�(���,�P�o@��V��/�`��ˀ댺����V�1	l�
�Y�w��7��8p�ճ��E�k��p���_n�X�������z�$lu�y��z��9�k	f֜�Åmuw;:��U�x���|�yö��*+&�#V��b�wW���j���4]w{�n�PЭ�7:�-pB�?��51L��ˋ%�����%\�f���g�x,��u�w�(|���JXx^#��v������u�w�JV͜���-c�fU�<�r�|�)h�`��h�o�d�kWw[��ۼ�v4<*-=��� Z�u���	ec��}E��q�8!�ڬ$�B�&�7n��}�vM;WWOh��e<�9ٴ�f��'\�����Ӳr��N�V��h���|�f;f�-��λX��F��`q��s�:����rfU7i��xݼ�q�a�[)��{��{#$Z�e.1���`z��[*���J�T�\0Q��ۣf�2H k2�[�eЊ�w���2N	��67�ݤ�|�լ�=��2���k�:V��d{|��`k���`�:V��A�Cy:��@	��_;�0]�=6L�{�HL��f��'P��q�ä=̩Xz���4f���4Y����VN|.�pA�<�IM� 	Ǩ��[ú��u�L]{ �PjՔ��raK�N�u9��[���U+t�:�]�Y��*��b�t��]pX_>������'2�5j�����t1�Њ��R��`��G���O����em��o�Z�y3f�[^�:q�'X�QgU�:c���N�@�w)�ܮj�x^N���d���z�u�I�:i�m�bT���I���n����*"��QD����E�Z�k*���[J�kEb,jUE*P��ҢXQH�PDTE����
����D����Qm�"��Pb* �2ڊ%� �
��B�TX��SKab"��(#YE�[X�[QkQ�l��S�[JUj���V�`Ķ�Qb[EKhĭ�QTP�Ub�ѥ.6ET�bTm�Q�X�Z�E�b�6�Bڊ����Ub1�(�DVj#l�j�`��AҨ��-b�VZV*�+l��Qk*��%��� �K[����+��X��屋�""��E�jb`��aPDV!Z*ZPU��UD����*"#"[D�Q �Q�U�UTb(�b�b��ܡA�X�TA�Qi[�aYB�bJ��m��Q�+E�m�S�(��,X"8�EU�TPU����Q��Q��(��
���1����K�*(�H���ب*��V
T���#mE�T`Q$�C���f��8�^�]�kg&ή<>��w�l���5�Z"�-�s�f���;F:WSzSS8Ҿ˭w�Ȍ���#��n�]���_UUi�/%�o�B��J�n����w���wMxoT!1�)r�H�Ï��^e��L�	�}��M����*��bbk��2�;=��P�lt�l+F8P�Բ�l�F��P =遍���Ba�V�/��v������x���\��cG�)��� [*�����+�R�r!��7b���6X��k�P��>L�R�g[h�N�o��ު��~r���"��F���9���R�pmy�^{i��%��z�y�5�]��)�E�;[�o�=�:�0k}gFB,-6����aֶ�\vq��K�ba���r�u']���E��v�b���f�(Bf�;�3��ӌ���c�Edwk�,�ku�jV��Y#�7ȳ�,�$�z|��z| ���o���a8E��.�~��m��5�j'Fab-#�l�Ĳׇ�)���V���l�����Q0��F)Y�Kk��ec���BN��BJb��'4޼�C|K'�a-�,R�=a�5�E֡t����.���+0B;�raGz�i>��v����\l]������͠5�F+���̯{s�d��P��:)ק 3ީQ*�{�"�~���{�2���[p�+b|�Q���\R�[�����5�w�Y�rU�\�^|��(��(p!�Ƥl	���K�{��vM�/��d�b7��@*���E���/`��ּ�:�ݐC �%إ�7�x�2VT�nt�F���XG)c�u���޶�a���B���H�H֖TE���h���緘���~N�Џ�ט��Ý�<#�B���]k��7���w{H˺���.�3�w��B�t�2�*L�r��X��֬�1>�s�n�lx�Crh�\e���:�~�Ɠsw
�ډ@kD���Dm���R'��,s���٪���PY\5�uw©��n$�L�G�{)y9=v'�y���z�T�7�M���ŏ2�؄�ו(a�ƫV��w$۰&��D�@�������|א��Eg����^Z�Oiٖm�K��VJ\=�r�R�����vN�n/ĮsDT����1��3e<F�H�<"��՛2��Mդ�cO�R��Ǣ����%s1��ϣt�Zh��;��Ws52l4<�x.����-�܌sw2Ɠ^�,U�T���͍�`k�cE�p��Օ�#|Y���e�~V7r��U���@S{U>�b ה��P��j�s��rkk����� �:���H��{7�'ZՏ�`SS%��ru��2�!5�$ ^X���VR��:ϫ0',�m9��͸��R���ٿ�=��E�KR淬�బ��Ն��蕌�/,rޯx�]�G��Aߕ:�W�3\�ט)r�N�%$Xa��q����\B'D���"]p5*��S$\-�5�f�7�+�3zt�	��D�p嫇�̵�����<oi��,��\�P�7�ս�V��^���F�#�9R�%�lJ22g�a���||A]�^1��P�t%��%��eg)�́�Ƽ���d.P=lu�8����L/��F�r�o��
㷳֏�e�hP�j�%Y9\\Vݥ|��� `������Z���b�����r�Uƃ�*�÷r�A;&�������ѡﻑ�])c�0���0�k��=,-��J�k5diZK���'�e��m��$:��65�c�tˠX)I��������� ����P5�!�ݩ��v�m�ҡ�^��ޜ�P�`6�CF�]RC8�Kk�Lv�;��q��{���6�mGm�P-Jܙ�,&e5�+I�C�*���]d�4-���V6<���"��4��t+�-T�1G��e\B��ԡVi�n��]����w�;��m�)��֒
���m\�95uv�|"*���jøxƷ;�9N�z֢p�Y���$d۔_�`��4�]v�l͟H���mG�h�����jfX�j�rw諭��&q{9-����h�8"�D�����Q�ZM�Dk4$1��0�r3,O1���)A����RE�{/�xMS�g�I��1��r������𡥪#M�̳���M������=B
��������p�ecPά!�����+>�Z��F<�oN��x =�[a��t[�k���T��˕�K��¸�l{���~3.����O��>s{j.4�:9�	�<��OV긯V��P��x�Z܉��<��{Ec�=W�M�w�vsɬ%��n����:��-��;��s�i_��B}�h���[�ܛ}Ζ��\q㮈p"ۯ���P򿱎1�s���`��j��ה�vC�������!U����mgNN�&�NL�.,�a�7�F�XT"��~R��p����UF����"���t�.	��c�����*dG��/Nk�͵�#�����l`��2�os^w��HCH�3Cs��(�#��W��
�������������ܱZ�������j�:��)P"^�nH�^��>��H�_*��!��ה��AWfB{3��.��X�LRcS����1K�qOy��/����j�:d]�WM�	_]L�}�^�Grb��+�0��o˨�����m��1�Zw��`݇�1fgњ�`7���_}�,!:�YC���k��F:�j�!�03�'�W��
�%W(�g�X�v&� �2tw
o5ƲM֔T���2-��/���W�#�� #aZ�=�
���k�v؃����m��ya�J'Rf�:��w��)vt`l֑t鍸�vZ$V��R��*��{�{B���E1Nb=S1z\{4O
�rt�9��3�&��4�C:�va��:���|�+��kssF`�:��aP�xHэ�[�hqn���K�_�����t��l�)�WkFݑ���Sȋ�2�쓅ߺ@����p�%��Ō�J��4K��(�K����SZ+33�<��I^㤦N�UAB�8]�H�#�̚MZ�<.�1>!�gѸ�t�{/�X[��K,c�m��P5��G��~k�`g���/bjP��>Y�&���>*M>���k:��z�*0?[���Y�k���5���
��\�<i�Le{�X�V��9~�>����}c�8�[�X�E�T�]2��P�M��#r֍�ũDPz"��WF.@yֺU907
�p�Oev���xCwc�R:��b;�r���|��)ܙʋ�a�)��D�F��Oa厞&�-��d��}C>��:v޾s�_.�0�eMA9S^��b���(į�p<���Ē�>�Ky{&��K�%��)ue�ܾ�{ޫ�Ю^cM.2��eQ�cI�2+�
���b����r�R�ˢ��53�v(��TnNY۹���ϩ�f�Me��.O��@Mt�_H	x�3^������+���_S�kT�ץ���7���l�X�y(��+Os���U8��WY99S�qi9�f���@z	��*�P��A^�c'�j48�������H�)�g�� b�����Z�*[H��B3=��u��H�o��o��y<���v���h4�b�r��`�،z/�\2��Y[��s�\�xn
tƠ��>Y�)�Vi[�,6���%źi[����|�~�vM|�?Q��PȘ�4#�y��[��+�w_��������m*g�"οk�JE���vD��Ē�t���6ؘYs�f���ʷqЦb�.j�r��M�<��-����1�;U�]a�c���FC�/-�\4!c�����$N����v�k]Y����Tt�1���Dx%/)-�0�ICc��&*V�g��¶�{�Ln߰�p�N��p��ٽ�g�D�ԧ��o�s��3�s���������L�y�kiP�fk��I+����bG�)Y��.uֳk�y��1��7J��o�C��h�]��Y������k{j�}J['�{tȲ�_J���_Z�75�������2�x�V��Z~��Ry�&�� T6% $[w5�죆��wJ�3x'L�Gk��J۔
�=A���yaLn�;'Z6"��J�4EL��͍��r*�'{�q�i7� K��A������B���,/����{��v��p��G[z+n\��\�W��3n:2�e]��q'r�w��|tB��UG#q���p�Q3Ů<;��ӛW<�d=7���;�<��1N��c!��`3��{�Nǣ�	U�p��%ښ��y���y$�ƶU-8l�O,�.`��mϧ��AE���#�C{^����a���ߒݭ#�c*��=�A]�^|�;��XXh`�
J��1���-hݻ!�Ü�ٹhʁa��D����v�1��^�P{2�ٍ�F�փ��9�ٳp�+��a_:DB E�~���.x� ���[�r.���Ny��:�Y!d�YW�g��\�5,�y%Q � ��q0��밎)�F)oT�E��Z�g��ϦV�]P[.���n�`g���`l���))w���4���^�3���G3��ٓk�(�vF�Y���u�F"K�$��}�w�kڝjK.�r���Y�x
H��1����{���ۻE);`N��0Ag�[G8.��D�}7U��,¢��i���,t��1U������ǒ8����N�Y�Z!22�!v��9hC:������(ە-X��}2��JG�k�G4�7-P��l{�~��fDu���^O:�O=3�7{�(F�r�(��+t��+Rϫ�Lv�:ncׯL�qm>"yT�w:<��#Ի�tz��P��)�%�v#bP��@zm-�M
�W��L�������k�ç�+M�"��)n�ș�c\��bW��1*�0��/G�6�ՙ!*OIlR�|p\�V{G�7}��U@�R~�@9:��k��U׈�@zo8z4��ܞ�ξ��9�E�;�l�C3�Fי\g���8/�{+��uav2Ƕ��w`<-�:qoC�	�%#�t���{�Yk�Tj��x��U\|&�C��7v����Cr%��VX;�R���K˻[Cc��`vZǃ�P�[�8�*����r	��yo�q��|li�NT�Oʝ��s(z��K���x�ߥ�A���#Ny%�ѐ/=;�ݞ�B�'�et�s��+��u��S�K|�q����rR����~ S���7�VP���N�b���Y+��:��(�6����g�:�Q�:/�_V侑m�lr-ij9
vtrqA��F�OEX����g�����k�<%pܗ/�5�CAVk���<����}��xߧ>Ÿ�w�K����*g�;�o�&�ܗ��-M�~EG�D����3}!o�����ટ�>L,�+C6�Fvo�{�'=Yi���J<���2�Z=)�+I��Ӭ�i�Ԅ���8����}/s�uj&FY[���F�۹�!F�<v+��l��T6�-��(�#��4.�ԊjC��偂���L��m��kO:�Ѵ�rZ	姳��0.Q,�L�����ǁәBgv��aM����oۏ�_�+F&0��*z��9�^;���Ч��azW� hN�<*ԝ5����UX�E���f��r�o�݀��d�8�`˲�e������-���j{B��X�͌Qc:�!���RG�~P×-�-	����켐ӽ<`]��#m?�p�5)�����}hx�R�)����x���U���&����d��m{�6FC�^�ѳ�Z����k���m�ZrK��I܃j{A&'��]=�v�6�E��A�1]����(�m&/(>��ӹ��f�]��}�P
�Du������F|�Ƶ��c���*�W�V�̒H��t�V�Y�=�M=UWaJu�m�9����rsY���<�E�ef,fH&�������=��8�3�]F���8���I�^��wB�I���zB>�2^��e�f�f��5y*������<y��d��p�y�9f-��]+P��L)CL�~겕[��PL��!���?U��<
y���3��jg��vy���^oi��{%�<�T�Q���9t:���8�iD��Ӛ+���t�D�E��6�P?�oOX�gF"��o]1�wZ7M�2	�xW�M�_�����XԺ�q&.
��_״yEu�tO����Q�*�vaQ�'6��oHa3�_m��x'ݨ���\r�Z<�����5���H��'y)ֹ��xҺ�.{��q�P�'F����g�Ԧy���*�%�A�s�B�]{74��(x��BJ�&\�b�C7�X{K47Thqa(����Q�����
{�^�nI	zV��LFk��[��"��l�Ըd�Gld�@�x�����wY���u�O���K�ެ��4�h�����S�5lZ=I�̡�m��T�
�*��4xGR�Kl�y|E�B��dI�D�x�s=>��i�t���u�u4sa�]��{u��)v��K	ê��mG+'�t��]D+M�V¿����,.d�+��H�B���QInR]�A��ۂv�:��d>t/Q�7s���.X�w�/.�$
���)��"}�&!q�A�p/@&�����9���f�>�\�1gD�Q��s6�{��������������;a��������ԭ�`A�dnGi�0T{�-�}����bn'�iCٺ,R���o,V����[%^.H�\�β5�˫ �t�.b�h��q���Ն�=v�Q��Sih�HGo:�VAט)r��oU�"�1�Y�6;A>%=�Uӫ'�܆}w�x�V���-��e&��p��LїRKS-��rm�ٍ��VIk�܇
zL�e[��<����	�A_��U��y�qmO���(18<�V\�6�9�J�5����9��pw$�x�^q���p��\Bk;A�]*F]#2jD�����#ƹ�1F��� �nT�J�uՏnu*�/���I�.���lwV�G W˹�/Z���GI�\~�=���3Wi8�V��Ô��ޝ�����m�Kd���r��I����'i]�9Cȋ�bJ�X�V�+j����%��4w�9Q:K����-�\�ht�/9�Ղ��CM�8
h�����=d��m��c���]'.^��6R|��mټ�`^���GJb�]:�sn��,p�vGv
�+��������vZ�����K	�� �y�w$���[���z4ϣ�����#u�$ޥh���CV1ͺ����i��L����]"u,K���X�`U3�7�J��ym]:��d�57�.·�EV[�s����F,���-�^'ݹ�n�+h���,C}���qB�1��淹WQ37��k�*e�;r���RW�Z�o�J0`)�)����zMG���kui^����i�];�.��Q�5��ٜ�zAG`�����;Z����� ]q�5��k����*��b��KaK[��;^I�;b�5�p�p��wJ˱:�uvn���;J
QJk�X暵,�7ul@,[]��(!�t^��X�8mj�4��;{F��`�N�J�[{PM��f�/���ԁL��}(Ayv�\�Bv�8�O�v�$��Q��ݷo.��%H��4�6�C�m�;�{�-�l����KWV�X��\�f^���|�5w����SƝ��t�w*7�A�w�� �W*�������)Y��E���ݐ4����})nn8i���n�H����،�Ew7���}CV��y�a|v���!:aR1�/Rpu�+,2�����+E�.E��m����e����1RI�Y��H�8��(�#��>c^��*���,�����#�_S�Lp}��<��:�}}��C�z(na����uX�P�@����  ��DD�PF5�A��H��"�Ke��(��PF+�b#�V,KB�DX�����T\�m,AV
����J�l�Q����E��Q�YiQ��"#)lF*����UUE�1jc�AQ�QEĠŀ��,EEX"���"ֱ�*EV,DEF+naF(��2* �Q�,�*"�1T�AQF( ŭEeeB�YX�P�3
(�F*##�9jŶTb1F*�e�DX�UV*�b�Ŋ�	�QAEE�e����*�UE�QEkQ�֥B�,�(�����q**��(���b�E�"��PY��,F�#%��D"1X"��T��
�AbG��b��DATEjV�"�����0EV(ŌU���*�*�R�����������(�""1rƕb���B�؂�1QUĪ���E��������/�'��h��]:v�h�۔��V�[<��&k90.�3�1�;R7��(^U�q����J_nsi�[��U�����I�g	�H���С"w��?�^b���������]kcX�^k��^F>�=uY��|���␰�o#��K�j,WS��8���\'�R��Z��%�	��}�k��2��{kå	�jXpږ�Ll�w�E�V}U�B:������zPn����[�s����UJ�$F@l�9���@YD�/Р�5�s�6e�Z�%���Wq��z���ظz��2�5�_۽ O���Hk�3�7%�~�5�:Ɗ�'���}�M��ofb���l�(<�����Ǚ�j;���KZ�-�IjH��Y���z���WP^��a)����Q��x���x��㔸h����Ez�D��Cwo�Z�Vj�6��0��ڴ �[Cҵ�'�xa.����cp��8?���V5˱����O*p�FO{�B�%�]\;��gW�/��Z�J�Bx�99���x�]�G��L>���3<�G_�ǯ�<9q؞(�N=�:���yz.!��&軗Z��?eޯ��ʃP[v�S����ڣմx����1#�.o=}p��E\:�������WV��E>92q���cMڵ؃�V�sh�a�C��r���R��P:��4���%+�%\��x����}RM�K�;�4�ݞ�K��G\�J��Nd�$}�%2o1��|����%oNx0�ꫳư�UaЭG�<Q�I�H
Zo�t���u�y��7��Q,����2Y1ܨ�ũ}hdF���9��V]�[=��Y��W~ݘMp$� H�����ҫ��( �] ���W"���N7�F1�*PC�{==�e�r���w�قm�K�ȿ�㥠��-�9�{�hL�è��������'���#o:r�qP?X��g����m�R䘙c��L"k���� ������vK��B����J�,��c�L*����\�j��X2��K>�Zy�nd���:��S=T����&Á�fu)uq�Þ�k���C�F�ZD�����-c;Ғ��lP��"ٗ�ؽ	��:=�3��u!�E���"�!��l	Bu"�.�X��~��.m��\�l�\�R�Q���ǯ7������r�L�5��!�ħR�\H����y�k���͎ (�7����ִ���z+~O�L')�K�O���I A�ޢ�G���k�ҌeuO�h�ͣ%.� [��a�t�lS�{|{��^�efq���ݪԃ'�w�Wf-�+;`�!��8���䚲�q�S7��G��/�[�͐q�N�ewr*_.�\4�]�H�8�4�Tr����YA��������u,�ש��xY�푢��:�E���\g���9x�3�X��ua�jS0���rŎM
uRI|���S� U~a�ע�l���Q[����iG��1>!��W�P�>���V�a�3����#de��8�bd���OV긮f�ǃ�~B]n��Bo�ׯ�m�Yܖ��=�G@q��7�H;T���XG	���ϧ���ǎ	z����#�5�?mo-�!>^����#�op�W�1�1��P�,�>Ÿ'�;�n�gG��W������hȖ3�\"�D�QA�7�F�XR/���wۼr3e	����i����־���.
���P�o�3�ߪdGT��j�Ӭ�U�Fv��8w�T���r�6��+!��e���wZ�)H�`�;�\e�Q�Cm`i:B�6%V-�m��Q'1l�hU�dM�:�S�v�(�ލ�t�X����Ю2�npP'��s�T��E�8��xE�z��\���M�����Kr�����1�O1<N�B���ks G �k�s�J����e���&{��Z�n4j��ΐ)��<&b�w��ƌX{�p�lCۛ�:�opܘ���sgT�"ϸc�+kO*��3s��:WQp�bb8y���C3^+C�p�MCw�e�n:�tƵ!PC��|�W���������eb�� �3���8�rtppl֑.X�uv<ԕ�Ⱬ�jJ��ٯ#�,*K1k����a�7Ń61E�U�7�o�HUN��ءN,�p����}ܬpg[c��+a#�<�S<5�̕��)/=)�X��Q��/�E�+B��2�_&�"NdԞ;��Աp�Nq�X�:�IA�eX]흢�z����
1�y�e�[�;2Km�D�u
Cs��9��~ۑ������_K���Daӊv��W�������"�Ώv'�&*�Ϲ�^[L����<�+�ۓe���>&�Q��X��R�6e9*4p�0�R��{)�2ߏXڅ�7�d�F�c�©���R�~x�=<�#�>�v���Wb����W�[�o�=�[���ְ����bdp�w�I��^g[��s������Pi���Y��N�Ohp.��(��h��:����9�R�n�'7��XC{[g&ڋ8Nē��T��_=^ 92���K��7�c�<C�}sU�[��� ���- tOe�^�����7�9��33(eD:��]*�C��K���b���%�������c^�Zԩ&pI���@T�5�8Ŝ�;aͺ����'�G�u�d���&�g�/�"-I�Z�u���4��Eb�b���#`��X�y(��+��28��z3��Y��Q��TH�
͢8�O�$0�L-q=�<�L%>f�>'h:�w���\/�rX��Ԓ�:��̄⧨�~�/�����ս�%�W��%��#��A�f�V��r9Z�iuP5g�bc��Icg���Z]h�|��Ss�iźB�2c�1�`���矽�n{��u(@��L��H�DC�С�;�C��y���cV�Z!Xsdp��e#�7�-�h�{����6z��D��Ѳ���W���ٶ*\���n9���Cν��w���:|cc�bT�`15]K
[I1���++H��Wa3��Zy�6o5���<u�ܠ�L����:|�`䔼���b�IC�y(��=��Emk6r�O�r[�˕׾�5���2k�'�> 6Ġ5$e7�qW�p�
w���Z�F*.'+����!��MҚ�,+v�4s�u����5DEG������aЩ�ͅ��J�+Ԯ`3n�����|��m��oVun9w�d�I,]_v�o9v�	x�M=ڤH�H-f�����OɼG!]ݹ�(�z�S���+M��+�����C����Ķ&^<���C65{�z�Нߕ��K�ߺo��]tP�`ʇnFl��[3L�d� ��S�'Z�(����}�!�3<�v��M�Ɲ.ui�ǯΌ��}�"\0����T���
�z�o(��܍�Vm����k9t���P�G�V��a�^�=��XZ�J�C,�` ��F��{���]������L�]iN\�.�]-8l����\9U��N&)[R�=+�}�-ُ9�Gor�Fe@kg�!h-���J_\4Y0�ĭ��WW��1���y��!��H[ʆ��"�4��	�I���\��`t��9k�V�Χ�E�7H��3�V�WOi0,���"?�#bu�RaA���b�*�,�m�bʱ~T�3��w��Xz_e�t��,�җ"�㥠c���
�.������Te䣽��1�����D8)�έ�wX~�ѐz%�`��y_�@=49��OR抾�U)��E�^s�d��.\���g1z�KB��*Z��1�:e�/�#�:���o�}Ů�t�r��]j^�b�Y�缻2�����ڠ��ނ>�ꂔ�����[��/�xhİp^�ò�h���u��<5�Ɠ[��hQ�o,�����wu��N�J�O��bZ�O^�{s��s��kZ������z�o�}��_eT�62����(BE�OzVS<S�a��NX�|�ק�cDӪ�Iwc�L��K�kXw��k��:��������*��,(fQ�{P���D1�=�2H��ǵW�~��NAO'Kuc���p�����X��ܹ6k����]U[��{[Q�]P�Y���m͊\GE{~�q`��^e���>+�0�V���w�ҮX���"m\�~;;�p'�g��V$�p���f��,�m^d��fh����a��.3*�0֪�ɷ"���a@�m���z�p�u'<<ý�E�k4*�������G�����G����'T�VF�{u��#�;ⅉ�^ꖳ�z�嬥�"���UfwxA;��Q���|F)Ϲ;�fetJ���>�61؅�t��^K��#EƜ-��<y��^�{ӧn�ܠ���N�*��7�eojje�a1a�5KOTΜ�u:zE�z��?R[l��.]�׫1��#"%D�9�F�XW�|X��V�01&�f^er��~����9n���d���k[V��(���}c�x��Da\ps�7|�NHv��}�)�ާ�G��l�JK�qП�������n����3�RX�љ���8hf`sn��T���纎��"#&��[ڱ��7g�j'ٷ�y�!��1eID@C�$�j�DuL�)�=��?+e�㼔�s �%��	�]C����ǥ�3��ժR*(9�����T��Y]�tܣuk��D��r��Ƈ^��"e�r���!�?�Q#���O%������{�/����-�Nc�MJ'��0򥇰W<0���\�z[��h���a驊�tӭ8�ɪy��v�D�XS��^�D�W�t�o:��Dw��)vtCfp��:cT.�ʉ���_v^�"��D��1K�k���qb�,M�me��>��1&�^�h>�#q��!P�6�]�c �D!D�1��h��,��{	Oư F����죇h�\�*L��ӻ��J;���F�:�Pp�mn�
xo���y����y���C��`�����@m�#��N�}�t.I��:@�4v|S�8��x�1�٥�������e=F�P��7e�]�	#$��*r�;U�e�g�n��Y6S�t�K���7bKU��6Gr��k+A�3�A=�qU��u`D��˙����6�T�PZ��uшUET��N&*�%�;Fu�\�Vc�%.�gz�w{&��k�y���ʤgs֍N8���s�Ғ��٨��߾���M����K�(R?x��K92Jf�f�������,P�~ZՑ~{���ѱ��ƈ��@�o�I_g���uc/����|���X]Tu�Pz��[��5���ܡ�]��o.���˺˭��-V���ob�1���g=U�D�Ĝh{C��G�Z+��˪�_P��qN<i^钣�^�,1��-�m�U��k��ۙ�H���v��UOW�)L��f;�nw��"����\�a��a��iL�����	�my1��V������ȏ+R���e$5��d�PaY�F)Z}q!��B}�V����4!a(��"�OS���K�i;e���ΰ���΍�T�(X�]�k��{�1�s/M�ɽ�7�@�׵����;�bOgl�{y���24�]����-�\n����������������t�C#���;Oy!|�����yn����Cz�����C��y���yÝ�G�u�/g��f��.�hZ�<�1vV��J���;3�#[)jN���L�9@\,s�֜]u�}��<����]�u��[5m���B��ěu�VN�nos���
Kǭ��Z��L�-�)�ۻK9n�e�W��ma�zk��}��p��.������Ϩ�"��*��/ �Yv�+�sk5b��#�!���U�bNwOJ_{��d:���1��O�� �B�D�X������m$��H墓�.Č`b���J?{Y�&8&�6/ٽRO]��nH���6r˸yಉ,(
�;u�P9�����;97����R�]��Ŏf���̚�&�d�����G�]0������5n�j����n��zO']\}�nO(>W��5,-�
cu�h�Nh�Ǳ%��[�KV��&gN�Ӣ��{�5�e�uҵ����9��	g�q�3	���\v�c٩�.l�ޅ\K�cѻ�u�C�-?�[C�D��.K�^����Ԇ�:(9�]��!H�f��1��r�g���'��p�9��p<5��c�\�S�
gu���%Ny׳)L�3e �<�W!KL0��.���
��y6r$���Q7��;�9P�[���b�S$Z�-�~�LE)}p�kf3��V��a�g�C�=�9���
zo)ޗ}J�Ԯ}J���:o�%�*�2Y1��`�r���=x��J�����-�j«�ԺR�S���Ժ�U��[�=���roU��̈:}�s�|(*�"���k\�:�vn���@�T������T��<�_#�Ѱ�I4��l���'�ݹ
�˕�KW��,����f,�+���Q�b�&9J��R�S��vM�uȥ��\-�D��Wwi�u�[YΥ��w����iV��bH�\H�X�*���V����h����{x79�]�R�f֚��b�}X�^�i�u`��%ց�J�����H�n���/m�����g>��t�.�a��H��!U��X;M�3���T��sjfi�Y�7�
meq�a<:��l�Y�'bT�1&��Zl��۫�W@�� {&��k������<Lnf�.�S#����@��E�k���H+��v±��}��GE�و�D୧�!9�;��n��Jǐ���3AtۭW�2ʵ˵'=�������Cm���}�(�ܭ�C�T�oz'f\/;�m(�Z�ڤml��XU��J����G��e�N�RgK÷�f� e�q�t&s�9�/%�Q�V"7��C��оb*���1�5�����j��c�h��Ve��c7Y'h�x3Q"Ȭ>+���0��O�����j^����U��DW���#��'Os�4�m����>�D:7�k�pfJ\�J_^E2��f�@.�7oI�2;K��cܕ��X��Qu�#����ܠG,���E#B��M�\��#����2N�+�縲�2�M�
ƶ�P��"�b��L=M�KaF�;�}3d�W�����������z-�t�Ƕ5;�Ws���|�yV,*Ħ�v����ހQ͔'�� @d�s���7u�]$�ŝjݤ��Y�/xU�9�2h���[����y�_Y��c��HG�P�<�5�����]/�h���]7�,��� �Y���F��x����y��F��k��1W�;.���f,(L.�y�:�,�ךoiq����$�!-uf�3��)����e�%Y���e֦�&p��Zv�/�B7���[��:�q�q�/z�jq��z�ەݚ�E���UQGg��a�������w�-�b粺'!�a�l���?��Ms;�s@�ׂ��U�$�e�T_Z�m�z[�іy5eٙ{]}��kw\r����%��t��|EѤV��qݹGk�ۓ�m��B��Ֆ�Q��47�}�叄óz��{�J��#᧶s�;��~�Rہ�������k�*O[*�˛��.Y���ל���7�}��]�8���R����i�'R��+S�j�YC6��7$_]���[�d7���;E�,��m�&^{�މ�ć!7^m����`������sqN����M���Ĭ�3κ�9J�zK9��IP�X��N�D��f���ܘ:/t�1�*�9v���9Kt�|�C�N�Uj����Wn�Fq��V���][ݙw����#�Yk>J��EX��5jX��JPR���c1X��(�E��(#�"���(�TF1-�R������TQEUVZ�X"#�*�Eb"��j(V#Z������Z�b�Ҋ�ڱ�,�TA`��EQU2�"�F��Z�UDAcG-Qj�U�V,L����5J��T�D\���X�Z���KAQ�ƥEQmm���Z�U�DG-��EDDETc��5�bDb�dk��UX�*8�b*���A5
b�V!iUe-�F �Q,[T*��T�cb
�(��X�SDb(*��(�(��*�Z*�m�,ĵ�5��T#+�5� �*�6�qQ� �db��1�V�qU�1�Ŭ��ڌ[eJ6��*�T����Q\�`�"�2��Q�(�ƌ`�"�U��)/�o���[���g���տ۶%ȏ+�*���&�'c4X��L��4E��ofwl��6i�Х)�� �.��.���$=�S��F�G�P��`�e�ƨ�\MF{��-�s�C;�cQqVzm��ަ&c2��D���yd!z�P	���\t�CO0���Q�ܻfWRޱݻl�3���	Z�EӖ"���ٴ�S�wFd�IcQ08B�p�YW+[�z]$r�7�0�K����Igr�g4�vbE�9vK��[	�Tw�I��͛���xVX)��Z��+j`����͕�YL(s,gD��l9P�a�|��Bm��V[�Y��:�]�z�AD����p�ɽ,`��5jd5Ya_��D�lJ�-�1�Y5A�NB]4�����&�B�X+Զ�G�q�o�����U���v�f�)=wwm�spt]s�=<V��pgQ.�^Sb��0��#�k�P�ِ����9�Ӵb�]F��Fy�h�m��7�;V�j� ����=���:���������������I�S������g�VS�TȖdZ|�����4�DW�(�ۅ��7gQ�s���^|��?5��TV���Amr��k�叱ȅ��J�0{�F���a�A?����3x2 Piɂ����1;�%����w�X6�T)v��]��ޮ�Y�mr�WKMe�| �����̧�X����Nv�k��r�c���VG�n�s`��I�[;�wx��M����4<ɵ�[=�>�٤E��h�����P��-������P�{��|t_�'d��!�S|���GE�Z���ʡX�.�3^���蕌��_�����v!L�nԱ�o.���Νm��q����v����T���!�5:U��op�V1�-L�,tB�Q����U�����h��ӮR����@��;Eܙ�R�V�<<J��2��,��Р[r�&w��Sa	8p#��\k��m�^b5�����xo��Ih�i
֗h(�c
}����r��xb$=ť!�k�GB,r7�q0�W�ب�[w<n�0xo��G��c�z�+�r�U�I�*���]�9*���yɕ�Æ\ޱ[�uN�b��r*�wfO@��B\e<�f'n�=įJ	�N���%׮xF
<��� �xe���x�r7���Z��%�þsȷj�����ebPR�U�bX�d�Q�t�9�wAWx:tp�yR��I>W�TWm�����]�:o�<��-)�S�lv�a\p\������W���h������ںt@�%2i��2�pe;]��z�qG_e���j�7�f$��J��;��cBjC�U;X�W$s�.U�k=�N�oT��o���#&�;�8�P��n؏D�h(+jA|�B�)nZ����H�&`@m��r�1R*'rˇ�hl\��0�#
�Z<3�!�r�J���>R�ݜ.��mf��R��j�>�D�Ē���P��"\�6F�T>�R�6�Gk���M���09�P�s4k�}~9�$���I5�TJs
�8���I�Q��L>��B��-�;����{L�'}���bb�U��4��ٌ�����)����wOy�W)�K�rF��6��U��J�A�j
��^�H�@����2v�`W�(h�-jȿ=ڍ����"��LK��֤�a4-�^vG��ĿQ�U�F1;c�����#�@�oB�G�v^�`���4kfz_>tP$wڤ#]Nímp��g��3�]̳�\x=����<������S|7�J���[�#t�N팅*��c5D<�>��	bv��O����Ih����:y�i���%9�@� \F9�o��KN�(f���`"��'pߥ�d�q#\�n^���q}��a������WD��C��{��_M�C7�d}��0��R�����*�H�PU�iL����\��L.n�S��3���%��w�}�H��H��:D־�#��y-y{�[;���{}�M�yP��˲�C��]�Z�p��s��V�I,�%��G2��5�Fn���AN��-d�@b�T��MY�PU�ٸq<�������u��TP�r��N��ȍt�{|$K|��:MIξčkP���v���m��3�h5�]�_�(o]m.8+jy_ˣ�V�����fP5���q�Ot]5�W�i��yf@�R@!�9|&_V�TƧ�5f�a��v�R�0Ҟ�Ţ�GO���^J���p���p�e#Ზ�긍���p�ʫoe�0qۺ��Q�N���c�9��/6:Rk�J��6���e!�n\��Q��P:�h��4�-�C8'�����2Oqa�a�(����g˸p�I,UE�F�1؊�w�s�h|Ԯ�>���"�~����Ɵ�����`M)����.�eڊ�ʚ-���&󹙾���YGr��v%K��(<��^�5-lXS�u�h�Nh�f�Fj0��2����&���%����S�l[�MB�:'�߮��51*�gh����gt�^J�Vu�d9O����X`��c��|wr1�K�M��Ό�&'��%�<�Lo�eX�e��XxL��y�Z���ߝ��*���?Y���Mh+9�m?*s#�����&�����_K#�lvbk�Ϸ��{Ї���iN���yut��K�S�jLo��&Ϋ�m�<����b閞=[�"�wQ]Ӄ��`Wm�DG���8rw2s��=�'f�^�ݩ�׷����Q51�vup�����j]�g�,$YC�\���M��'����<�yy:�����Up�KN=�����(�5W]u�a�y���ۇ|�Mj���m�v���k��E��7�t�T)}p�kf5�Y��n��\��+�>��`̜�[w��ݞ5�U�+�F)P�7�㮝c��3=�Ɏ�a������$j��;w����&7r�	�ї�#Mh--#������]Z�.<f{%�"��^B�p��++�q��)��c�'�C�#�Yo%�K)r,�KA<���=��S��<�:����´�#�|�GC���匵wx�l��,t��:�w���EϬP#e�룹����𨣖M���N��S�朷.�H��.�Ļ��i��
NHD��Me�)�s**//��㾴8���`�<N
�ޒ���1�r!)xT �&X~��k6�νJ��M��HA0�$�i�_�õ�҅ၵ5��;*�
�� _��+H]�F'���Aꉶ5V۷XO[���پ�&�e䫉8&��eP$�C��pIͫ�τ��,3�\��Ӣ��K-em�Sf�&�Q���v��M�R�go��٩*ͥ/2�MC�v�u徫c��W��"���K�q
�E�#c������N�W �l�mm��h[k)���|�����I�\��)Ķ�)T_����D��BwI�tF�y͊Z"�:�H�Mx���n���Ì�jƷ��[��SwsFj�-,��RQ1-�<,��׶�1:�!�^+qp����Og��,�K�������cP+{�1�;%�V&VrԼf,.�;l����Nc�.V��:.j,�A�T�F�.���f���2.#n�;�:�2�c�P�#�R�b�+Ն�î�xv���s16���̡�9Tٯ_M�e2n6�j���s<R�g��=A�y�߶OKٷ�R�g�0ia`z*��(p!}Y����1�1�sT:����dw8F��=�WӲ ��w�_��6�e(�F�\(k(2g��G���)�:�U棬����#��'ٺ��A͉A��<C���Ih����_{$��KbԸz�T��x�9�C5muȿ"�#q�P����X컭V�#�;��ҕgj���\R4qU�M�}�u�yЬ-��]�t:��c��n��Ucd����9ǃ�C1a�xYJ����������j&���<ۍ+ݠf��1e�E�՚+�.yE���/k�]t��s�J�EX;-��yږ�7˝�u����<��H��N@�x��{ݡ�����X��ky����Ͱ���6��)p�D�z]�a����qą�����2z��V6R���\O�TZ# G���A��ph��Wz�+"�WfqkFk�m�w
�FA����Z������i��ߨ�m9���C�W�;:=9Yw:�EC�S��/�s8�QՕ�/]�<l<�����)�]��j~�(['Ns��]��l,���%,q�U�Ca��/���aC?�]ل��G����ua�:�����lxsnf���}�;ўN��X���P��]�6$�����#����^R��"��{� �ysWf�n�9���{�ʋ��X�;)�D�ΥKyV��3M��C֒U��T�W5��h��E�OtDa�k���O�֡�e>F�݌����$1'�`7^�y�s��.�|����ӥ�Ƽ��ؚ�X�/���>�S<,��qbF��Y�I+��x�WX��YK�Kz/�}6����wsX�E�<����[U����zxB&��:�����b$<i�=�\ُ��k�S�֒5�Q��I�6˒������]����8߮+(�έ��,')�S��	��OqY��bؙ�Z��[֮k�s,����s��=��dc(�M7QY��Ļ�yQ����g���M�ӧ�V�n1R�V	ޕ0����׏������^�[Ø�z���S���ƢP�X.
�������o�j�pgdk�%�f�r�mGؼ"��n�������ۙ�H�x?I�v�N1ap�黩�V���P���=�C5��L4�:2
㚼"�F#`��ĳ�wܑ�L��\�A�c;܃��Eh����O��$V(�Xqz�쉿)���Ӟ�;��yYn�Xb�_6�#�Q��$�K��L�W*�.V��1��@:����E�7�4Yd(��xr�(����4v�ͻ@�#A'�O}B�����x�#�������t���8�v����[��mm����KD���&Kԉ4sXP����ט���X�'��Q�݃ܕ�9ǫ�l2���s^{}pٱ��g�F��Z���6��lb�#;;/k[�uU\��B�?9E��9�^������Ǎ����ŵ,8l)m$�R;�u�@�ӹ�=]~��9<�K�A��cE�	W�h�Z|<:�"DX9%/'���{�n�xO�א����-��1X��fmx�t��'������g6T��z����tu>+��/h�~J�غ��vЏ�4a5����'���X��NASZpr���g'��yv[l䮙j��
�O���@�>'C��޲;@��vHjNO-�����:������@�^��Եh�K�c.��bǙw�h�`.5� /6% -S�R��fK��ښ��)��)϶ٳ^�[K,������O>2��g��{���5����>!�w(%��x�%bF��2��7�������%Ǟ��b�f�ôT<�S�6��d*�O��Tf��:)�M�����h���B����P�RR\0�<�jDl)�id���g#�t=��z��[�WS��	�K�(n��\;"â�ƚ�����-
\|=yZF�f-���@8��L��d�`��t����Zp0،x��Ӫ�M
'�m�R�Ց'���
X׬
�
b끠��$lp��t�W���y�[1��%oM�NI�n6�S��)7v8�yj�,���R��ۀ�\�}�j�,���00�C�GTd"9ٷy����`p�Jݯ}�=j4�-i���sH��Í���\MFz���;��c��d⥝ь��]ȸ�s�8�J|��B���%��Ȳ�� ��am!��H��ݣ���|0"���k�%·)�7`cX���`��S�!׎��̋F:'B+����ev�5�Wh�pw
b��l[{oyuꬹIt��mdrjbG���I�]z�3�nO.�ӧ��'Y��kL�٥v�fb6)��I�t���j��nl�Z.��ZX:T��F�ⰸ㡊�|��Eu�X�V;�\7�Kh�rIC���N��뮫���K�D}�LmD�jO�oIGt)�sNE�vbE�9vn�ƶ���G*��,�ψ�)F@�}J,q���@ySZM�C8�5Z�p���Þ�P�`6�C��z�#݉�ף��e��Lh�5[����&-3�,v�ޔ0@ٚ�2���� 9�@����%W��jٝ�xִd���l�%�:��[e��qϩ��xA,�b��Չ��&���������<\��4`5���]�\�9VY���m���h��ć	�'���ڋ����žW;M�hA��bW��S��3�7Y)�uЊAgH���Py�ħ\1���䀬���؜���61���<��*�]�*6���&�Σ��z]�z(v�X�sܮ���s���sK�*�)s��\e��H�����X9��_�[��y=�:�͑�=�H�kf��_��ꔡ��6#ʛ�1{L�6=��+�|gTl�e��4%���-�׌�eA�@�%K��n�.��ڑSYhA�b���6G�뽇��G+T͔��9���;�.%dі��
E�v�f�8��[4�c3�M��bhf�}c�3�W�T�׉�Z �/dԧ�,_.��n9J����p��g(0�Gw�ۜ�C��tI]���W^���:�݆�\9�p%����ťZ۩X�aea繴����)x�R��~q�к�f�Q5)��y6Z�D���w�`��_7��O�`��Q8K���:`�<��]���w|o�Z���}-�ۋJ�m���]�Q3���Y�o${�d�b���%n�;g*u�d�r�+`��fwC�l�����C�6,z�Լ\{�m`C4Ca�r������n���R��VE5��5>�����j'G�����])�J��CBҝÓ8,*�{��R�Mt�L�tw�Y����w�%bήm���iG�U�p�}zD�����L����x�ا�rS+I�y�7�Q��aeIPt��E�8�V�]Ś�h�;k�謁�]�����t�[9[�-���8���q��$�}֑D�jG�D�Um�}Y�6��6�Q�.Xt2�Rp@�>��v�l��u�JDc�5u�S�:�kf���S�Y�Go5J���j�o���Z������%�-��C��8t�}���F�\�P�ӐZb�J�Q�̭�&h�7(���陬^�����*#��O��W�Y�F�A�}�����LO�L��2Էt�]!W�t���*�И��i�u�y�p�%�56���4
�}˧��wUۄ���u��4\��`����U״����#��H\�,S��Ty��_r� �ual�t��Rj�v ��k�n�nfuk�V$�핸"�Vfe\# j��)-�zaF���]Dn��f��דUNC�В�q����ue8E_n�tS.���Ss&�PU������1�Vpq8y��Of��wV2� O����;E:��uǞ;Oc�^�����v��[�x	��v|F�ء̾���Ҥ��j˼& kkYC*�9����ۅ��4�Z�Jm�ȡYF�n���J�M�{�r�Z�� �@�V�j��>�3Zv�6`�iҸ���S�O����&gjݦ7��k}W��lAta����kݥ�Ma�6r��8W`-9o;��N�tпʼ�W4_�Tmy��h�J�ϐ.�8+,�fb,t�{���#�wB�k�@�
���#��mnmҔH�0�VHGGD��;AX`-�ͭ�'�w�u�[�(f�K��J��mM�E�:��v���F���F�A�]�BM�E[����^�Z��޸5$u�ܺ(�w
y�s�%e�|� զ���q:Y�ߢ^u3�éE�\��8���!�Yv�EhYA�:e�͛�ױbܭ���o%�G�e�+�29�ǚ໎��.���\��Ņ���F��s�6>�`!-�H�u������eUUX+�P`��"�QITE��e0UV(���#Z��CRV��K+c#l�(�QF+[��ڂF8�V���Q-B���µ.RTEm�q����*�E�b�1L���UH��X���m,R�ATUDD��
�X���!���+B�@X����R���6ьc
���X��Z�2�PX*��IA0�E*UT���TdTE��6�k*
���E��.2��**�
D���a��e��H����4R��V1DkPD*U����b��*�DX�*֫iV"�YZ(8�.Z2���-,E����ATEQ*��lEF8خ���h0��(�"�����E�KeF,U���0�V[b���dZ�c�qUr�F#Պ���Q"���Q#Eg�w�|n�=���=߸���������+zeJ��YV�4d�AB�w*��'`4�dָfto���Ⱕz�h�' �m��0Ws�@����q���xa�U?,���]CS���+#����\yX�8����M��`�.ukL͝ʨ�q�-=����w�C��dK�EV�.�Z���*Dv��*n���|��3�J�V�ݲx�����u���;�:�L_����P�nfx<� �}��w��uK�	�͜����y^/NDk��[]r.c��k��!��e��˺�bG�p/I�޳t��pf^��{�b����P�A���+8c���V����X"��D����qI�������՚`!d����bPur�vxE��ʖ�����S�Fz-�����/�7��V�h^+-��
�c_�Z��ض�W��/ibc9׷���-��D���!�p�g9<F�qÖ#�'���H�����ź�k�N�[��)!n�,�O�v)�b^�Gy?!�j��Hi��
� �=a��
�]#�<���E;h�h��<�#7yj�|�ˏ���)뺡	��.^$h�f[�l�/(f]ѹGGw�3A~O	��d�u4$a�@|0/�j�L�~�g!*Vn��.w��χ�l�RV-s��&݆�Xo0;K�KnYݮs����;٭՛$�����S�nQɂ�Jw9�z�A�a�i�Kzދ��K��f��6�ݩ�r�΅��ƶ�fYi�6�d=��{�s�m�'�=}���*x�u�=����)�c�bJ�,Jr^S-�rSyڢ(�z�Q+�t����˵�|>ԳL4�K\|3)�7�P�vY4�c����Z�c5�POG riZU�+��.!�W{�p�p���p��H�	l�f��X$`3��y͉���퍑���Coj7N5<:�,��ơ���F1?��"�����}(�+�0g_wf�+f�7�\C�vt0�¢�b7�[Ø�;��TϰUcQ(q,���B~�3�9��Up`��GTJ���;�3��ӌ���c�ʬ^��̤�>>�Se���� �����z�-@:�@�@�)�}0�s�^��7�0�Ѱb�,s�2�N��r���o�]�ĩ����PD�H�Q0��)W�8�_�e���z`be��~�.p�X��CK	jZ	;�e*���k�eYҝ1��Qoo��[9��&%t�W����bn�n�4�y��2]�~�4 �b�B���[ָ�R�|�8s��|�l�^(��j���`5;W��C���9��Y�w�!t���
��g^�Wj�
��^�K��H��ŉ�Ð�h������i��gl��el�.ڔ��=���&\�:�����w��{;/R
9ft�Io
ݝ��ΉW�%
E�-}�jAo]���>Պ�ö�a�r�td)�� �k�
��⮵��{��Rcaw���g�9]O�Y��G�u�(;V6WZ���̦*�R9�bPUqK}H�V�0��Y+g/]+�s��G��b�̕��K�ccǢT�d�MVK��3R^
��r2�魅{��v�+���Wi�j,�p{9�Lj���lIH�"V�sU��g',��X��Y����P�I<���x^敖��2�.��]���@�U� QpSx���{u4YoRG��䑕�nS��͚鴲�\�/-�
_<T��>jX[�8���b�j=��жUc�%�C�8�ԑ���X����3e����I���p���{���QOy�;c뵣��ఱ�%3��3~�h���-;����P�RR\0�ʿ^�]j6I/�{��~���Z�u*-ڜ�w�S(�x��gF�g�2��f�p��w��|�PH�D��6���ȼ�Q�<�R���E��6w
x�\}�V�;�R�_o+��y+��X'e��,�R��-ivJl�J��\er�Y�4u��j$�Y�+�r�1ً�4v����t�c�M=�.a�����Nw�m]�H
�m��Z�%/�52�\\��]�h�oVk���+$u�2�t�ʵݺv`�彼�vU
�J���J\�UP_S�L�~��7���R���2��vNtW1z�[�����ʀ�ә��1i���GIDמ�p8Z(��-�܍v"���Ӹ�z��sI������ͯlƏXQ�akMh,%�s	��n�8��o+�X��E����{Ѭ�($Ӱ�[�r%�޹�Cq(u�<��B�Δ�W, ��{sKH�ܪ,}�7���Z�Z1?D�<7g�Zv8�e���FܨEչc-_w���[@��R�Lv���#����7��"�`艊�0�jɯ���pb:��U��˴�;�zӯN�|���U鹳=u@ǒGR炩�;r`G����ޜ��{��"��ۿ\.}����o;�+�"*#�Β��Z�+Lv���7��jo�}Yai.k�p����2��u8(�� -p�a��u@Ck��%��L
]���|��/�wcֻ����ڀ���[���=ϰц5��Wy,���*�0�-	��֊q<U�� �|j
�dG3e^L~��3 18����� �Q�"�J�A=X�0wQ�Q��m����M�,��s�9�F��<������m�R=NV-:CH� �V�8�d4V�ڰ�8���Z��m��\Ec����V+|���:M:�@R����l��ѫ��'f�8=^E'2���%�6���Z8\�m���F�6�_F`vv
�KfS����h����}��@s�������+�Y�@� ��ފ�����̖LX�{��#S�T�X�����'�KX=�%dv��e�a�U�c��V��\�X��Յ^���ܝ��!���TٯMLu	Ux��̏��}���oŹc��ʕڥ Lwm�]�챺��dh�w��/
X�k�jc�U��}�q�5.ߥ���|�a딆���	Q�Ʃi�yLwc���%����L��ά��,��#g��e������޼��Y�@!Ⱦ,Z�\�{\O�uݠ�����(��d[л�6��J��q٪�^PN*dB����/NF�1s���yz4��hz˺՛���V���6T]v�vkH���>�t�b�PW�L�Y��S��ƇV�dL��S�S0���B6�����ֹD��Ӯ�/�����i��P�1�rR֑g�r���Uhv_)��@�L
����)V�R���rV:ޣ:#���hA��2��Yib�p���I��
��C�Y�y��gJ��xM�Fٌ��Wk܇��.]����2�rPQ�|��diől�eE܂\��3�M�+��X�Ȭk%��j��tT���t�]�or���o��i`��@��kRt��
�]D�b��&lf�p�-!yA蓩==�	��gFx6kI�9)�x�D�)iH�Z�6;S�;δ��'0.�2�yK���������7O7ؼ$4�PÌT���]�DB�rJ�^�W7Y�R
^ek�sǵ��@=X�]�d�I1�P���w���R�č":�}��R��!��x�gc2��|��1�]��GW���,��,_��I5��*%9�[�GIh�5����.��9̀��T��ݱ;�fOQ�Ҽ��,��YC��������X�ǟs�&�m0ͩ�Ȝ���d�\���� �[�����漡��{R��1>Nd��i����뎽���2{�ђ,h~M�"��F��sî9�����ץ�|��y�p����I\�s|�ݶS���������~�u�\C�Vtb,-7箘��;��<���3C	�/��,�C9y��y��}n>�شX�v��]�Q(Bg�S�c#��ӌ���<�=�9ٿ���k�I�#�R���m)ۃ���y�{�38�=�)
���4o˴�s���
�i5O��m��N�a���u��Xln;���-����U��؄N���t��:r��^����Jd��vS��+��q�ґ�o)~������P�K��R�;}�Y�U��E���3�n)�ŀ2/���b��7��t��ġ�q�!��Q�m�I��gs�"|�Z��3.�i��g�&Z$W�D��q�@U�O�$0�O�Ħǡ�x��w�����ԛ����B�'��^ę�*U.\�7�1���uu���oc���oJ�P��$:Ԗa�P�O�h�F�#><F�_%آog��<'�W�����Q���P����d��������]��[t��[�.˲,L�d��D�q�a
��Z)�i�}#.������{<��Z]h�a�U��*��zձb�\S��9����Y]�'[��u)�����ﮍ�0Tu\�ٯi�7\�w<T`���ȶ����bH�lm��m̻r����o-�I@&R3��mi���3��]E�fǳ�$�C_�7�ȑ����&����׻ܴ�{cu�l��:�Yk�E��|)2�.BǙuy�u��]d�C�	[�oEww 0p�� ?l�|Ğv��cEg�����y�C��q�,��QKE��Fs�AG`7�:�-�<�#6TˮÌmb]{����cw{݌LX�i���ڥ'��]s��9O�ȷ��49	�=��s:����x���/q�>�xto��:�itmN��p�D��.
����LG�]��6_ikf++����ɗ�̂v���i-�`��@�P�+"����j��^ɒ��b�v�1�O�k�����+���dM�5�J�ᣤ�~˨�l(;#�L��vPÆj�G�~te�ٽ�m�6�λzd��_*i-eq������ ~lo+�k�cE�p���>Se��
���hSe85p��IT�:�����l������L�lqu����R��v�L�:�Ow-L��s�(�t�gҗ���.�����[&�1��ù�κ�Z�IT��V&�I���~j%oNx0�ꫲ�j�Cő��ҡ��n��}\�aP�z(�Q���k��|���mu�ϳС�����I	x�$08����D��]S�u��'n�=J�V�����h���c��t�����W�wRђ�:�%VtH�t`�,H���
��;MT\�n"v�7�"���|�EӖ"��)�m��%���R`r���g]Z��I�^.JUY�WAq�Єd�����;�Fڞg4�vbD���13Cv�;Ȏ߫{x�љ�|;���+���kr��١��+�Li��j����pM��C�O�iy]���:����9TĐwU�̽�h�N�i��������0��ky�lt�3�"�%������ch� ��7�)�M�pN{�&wR��=Y늃��Gז�ixnZ�95��c8�5].����/��S���)���l3{s��i`���ʅ��Β8֤�i�p�0�Cʩ|��f)��$�ߧ"�n�RӰ�x����b6%q�Q�!��Y,Mm#ؼ�7�=x��5�=�=-]f8��S�9��q&��3"��p/�v%Nh�Lч�r6�{G}5�(vlѶN�F����^e���/ђb�La;�&'��@�g��F����azj9l���[��;z�X:t�+&Pk�;E��j�]�*5d|�L��	�����R��.m�}���vǾ�^GҍT��ˏ���2t6E���dFj�h��<��DӼ�z�,1o��z$,z��@~�`v~klyi��y:�z���l{+�W���3	eU�^�Q����P��9����-�sv�離��ǎ	z������8c���.�ا�g�5]\��Y�q�:�Ō�.��5KO;�7W��Ŕ%'d����^�!,�e+�����P��t�h)�)=.qhd�coB�Vƅ�Ԍ�	�������21un���6�DI�y7����6D|8�RN��Zc+8�x/vW
�\n�������1�G�(��&��]�q</�p0q�6Y��-���n�"�����G}��B�|X�)u����w|8'X)�*J# O+�u�{��˒?#ܒZ}�#]TҘ:S/N{\�m����뉄"�ب�;(9 p9�\����u�̹E��!E@,lV(.1���]P�A���+8c7�Xk}�v27��M�N���*d�㚺N����ԁ
�]�œ�(��bPur�vxE��U�R�C���5�l�[�=s���ϯ:�Kr���+G1��V������J^�d�W�t���@;3��	����1��N����G�iQ×�<D�H��e-)Ҙ�����8Q�؋���i�y
Д�k[�����7ؼ$4�
q��va����5�J"�s�J`��n.�U��u>e�^�ۅ�J��f��&�)by;��(�_��4C��3N�0�,c�&��N�wn�[���[�"����rK}w���V5��I1��F8��[k����o,�
�tWkJ��]и�FϦ�/��LpNס�y��X���w������֚�a�>�=��ױ��l�WYx.Xq+;��/�#��!��]ya���5��ɹ��@p ��{*u���bE����tZ뒞 kE�giV���n۹��LS���J�y�ȸ��޺
�k��4�Ŕ>�Mj�ۛ�%�k��k��Q�P�j�X݈��ծ�ۢ��]��	��I�E���ٱ>.%�;���$�-<3Tr��ad�s뭵�V,H����Y�u���`�b<�@�2Q}JK�_C��V�[�IC3�2��[8��d�+n�Ҫ���U�B�!iH�$����u�l����МQf�}K(����m'Iu�g�wa8��mG�h�!M���M����y����a����c�˙����:9�2��n���19��㣘1��a��m*A�cy�hr#W��w]���옧�c���{��#1ȸ�y�{P�r��<�ǻN�8�z#r�u�Vq�YU� 묶f��KUt��e����Ea��9�*tɷ�n�\CW/�7�VN��-w��{� jc��xz�^��OӍ9m�ub��M�s��Y׳b]������U�����[a��]ύР����[ʺ㍞�9�3kq;�s+�x���ݼ �\�]�V�"����2�ut�-�O�G��篞Gd���8��X�y��dX��I��覝;��8�({iN��3 �;r>������.*wp�܊�s8�I\�n����)��":��(֔SY����w׻O�t�:��s�6�Ӹ7�f?Z��س����2�IH���;)�]nK���<�Q�Z��(�y���p|�,����r�'�S(]nv���`5���'�];˭�Ks���V�M����������#���;K�=���jޞ�CD�eN�+���/.�ҫ�l�m�b���XU���Z Z*@�a�u������Z�wTN�ĖE{M�u�J�#� �pz:-�U���tgv�U��臗WK����R��99�תRk;C�qL�k
o��1�F;C3&`Ln@��w�'C���Y�lk���yР~�b�@�� ��}���H��-�/�Z��}r�N9�7[�[c�l�.f`XܚQ�M÷ܞd���� М�F-k4�����,(c2��C�]d�����1�QgN+ꂵ��P'^�
�F�P�v��y�R��Ɉ��iv�d�+C{<ѬI��f�5��Mj0u�Mo	ԥ���R��YnQ8=;���&���.�jSS�(�w7��e]���[G<�y��M�;���6�����N�����%�n���N�3viY��mǩ�e�j�,{6�c#�]�����%n�Ϻ'�(�c�G:y�8.(!��h�8���y�c�d��3����.W7��^e5I)�|B��:u�u�����J۴�P�v�D� > "�����R�,X��V�cZ(��2ĭ2�X�Q`���qE8QQ�Rƶ"���*�(����0b��T���h�����B�TE�AULj""�kG3jTDF"�B�
�TQ�fe��Qb1"(��E�%Qq(�-J��QkPQV��Z�UkI���1�%d�V���ETQ�1TDUc�q���Ҏf�����TAb�(�)m�,%�(�,`��,b
��+Z֊���*�U�TE��҂��"�b(cAAF	�k%q
�(�UC)Z�DDEʫQQ"�� �ib���A���eR�YEEA[h�TFe��b
#�4��(֬\nZ�Ҧ���l*�V".[5��Q���۫��(���V��  �A)�G:��޴�>���*�o4@T�%9���v7'�m4K]M'\S��8�L���Dn��wGK�hj�ޡ�� W���{�盞�~k�mɲƨ9����^�Hׄd���6h(ו���t̨�jB�z�`�P��gu��j7O3�{�,��]z}h_)�aq�
wف����uJUf���'��̀�$\Te�}T��A��=t�k���u���Ƭnzgh�^nL�NjxX]�29o�����@o�E���	�T��ΗKNG�a����cڦ�X�S�{`�9B����y̡ZRP���M=�I�D���F&�B_(��
㚪��z�k��d���苑�u0���V+��t�O[��JrG=�WY��uS��J-�"���3�o��Wj�&�a(;�/��T ��HI�*�L��tP�z\�X�1��++��}�ɮ�ƣ6��lH��^c�{��ɒ�<F�Ix�B�k�;O�u��G��"1�W��(�#2ts�Z=M�̱��,5�����{��{Ȁ¸f��W�.R�������#��42���|�v�
k�+�c�l؎Æ��(j�뺦�V�" �L˶-��^-��7��1i]Js9�N]	�m�o��&fK໒�6�Nu�Q���u�|���=w���oRY^��S�д�6�h�P���ޛ�.����x���0�&ޞ�s4�v&��2������^ݾ��Kc���7VK�ϣ��~��u�WN�}WŊk���4�J]q��7ҙ�=!1�A�s��F�Z����j�U�%�ڈ��-�%�ŋ�&2��ņ�T�7.����3Y������}����DL��N
���>�(�Ũ+D���Reȸ]f�Ws�鄇���į��q��S�1��$��R>ry�֓C�Eo���T#Zʺ��ƊZ�5��s�Ӷ2'�N���h��b��Ǳ+��0Ϸ��:�,�߀�����c晾��P��ۍ�oʎ�zǹY��\����}���E>�+/*Bᮨ��:�>�1j���l���U	��T,^7�<��y�B�;�܂�D�<t�q�Y�f]I��������lh�)w�+����:OW�E� m[Z:k�*oy����g����q�+=^Se�U⋿�j��ږ+��ւ�H�{�H��pÉ�;yp&��9nm1�^���wٔ�c5�ޘa�΅y���cxA
}&b����N�^Z�g�,�F�-��.�lw͚ۅ
�#p�҂����g���&\	�݆��,dy�e��H��Jv)�r��D�ݏv�+���K���-�K}��Ɔ�Vț�Y}�G;���ޡT�ҙ��[���l\�$}�X��4��b�,�s��h���<��ͅW}�bݐ;��40����-�Tٌq�# �ւ�ZG4�!w��ww�+^� ��)))J���"�܍vmQ���Ny��:�吅��P�(�M<UaO^�*7J�7o��<bx������e�+uLY�77�W�9,e��.�JX����qO���O�(�o$�^%F�
\,#'���7�KU��ul^��-
:�1�"�sJg�YH��'����V�\�L���s�\�f Rt�5�9蕔7|���<2��ۧ'�q)���h5#a���!ﳍjN���mïՇ���_a!v܉f2��lK�Gb���ʹ��b7(C�Tl�o��K5�=���n�2�0�n�6��4�Ϧ�j$��fD9*�bV��RFӛ!�Z6����߭�89����R��X}~��cA�#�781[Δ��7Y)�T�w�kp�wc��n��iю�.�
6r*����2���V��G�X��������!exE^촲�=|+�?x�`맵�i�ݎ�M&Ref�z�9ܷ��j�$����f��>=����|"+���J:��X�ĳ.dʝ]k�<�����dVf�՞]2��c���;����/5����_#��pJ�L`�i=��N�~�E� _�«N���cҮ=b~2������M�b��l��Ei���O�d vx~o�t���U��V�=YJ�꠸�U�nrsB}x���jg?.Y+��XSR&����'F�:wcs�B������JߌXU�譡�W�
���3m$��)��s)wUvX3�+�W�q�e�8��t�p���;�"*!�(i�ǣ�Z�(|����hߜ<WV�{4P��%_�uj�m���o�>7�'ז�b9�,ݸM��*S����Z���ꤗ�F��t�h5�á�G'���y ����O�w���/c�og��֣����PR��l�����y�������~l"W|�]�h�^��w�ŧ1\<+��՞@R��������֙b�q��wZE���KNՉ�K���{��H�����[
d�Rs��\}j����� EhX�Ğ÷1<\�X=K��/4���;T��.��a��b�.�`R�����t卿:�̞"N�Z�:y�ú
��I�bJ�Bܸ�Gs!����KnĄ�ݒ���>�p����1�~��i&��T\��������J.��>BžC���^Q�$$����j+���� e_gV.��S����ضɟG[1h�=���x!�T���ͳ$�E�0�_.��i�.��&3c���q�������`(a�R�Ck��k�c}i��78��}��B��ΦDnE�\<(����q$�X����G#��4k��+��;I����JI	�"E�6�\T������Cc6:I���0:1��]�;�� a�;�r��#�����`G�@��y|�LpT�z�b~2�Տs$p>�t'M[���-�UD����$06e-!������ɲ�PsHg�et� mU��|����v�����:ߊ�r�h��Yrc0�Csî9��_�4�x�Z�'=���Z[~��1���ȝU��EŁ�[�׭�Xx�ǧ����<�뽏D��� �f��i'՝+w�%���q3�netW҃%L�uH8�t�����1���t*A�eξ���t���Gp�6�Y
�.�<[�+� g����R�@o���iW�\��:�	�n�e^�\��tf֑�������S:��08�?��$+L,8�F"i�\�B�1dP\-�}1�E���
�r�̔�WJ�{�]�D �����&�̦_�ip�&�.=��� /[�w�Y}�L����)�|���}9	er�9\,�u83�WG(�:�����ZTB��E6�'��1\S�R��w�HB��r���º����ܮA	:��	)��q+v�6ac��!ϒ''<�ԫ�u�r�u�,��[����}�Y%X�� s�����&��ᇵ1�����#Լbf��F���)����f�S�L�*�ޔ9�:��o�e�nU�V��C�<�/��D��hu �u���K�9��4�D(x�(O^=��Üex���*��gk-[�K�"0�պA���[����<I,B��ٶ*(i��5���t��+�y��;ɋ�!ŎX�jE��7U��V~��b�U�&�IZE%�ƍ�ۨ��߲�OT0����*�����9��"L�d����r]؞���Jy:��,
�"�i����CTk[x�j���D��)*�F;��(MI��Fuɳ
��=����܊� G�'�jħ��'T��S��,)�
ݨ�b���J�戯d�LM�n�k0�=�f��z�-�o�S� �li�����E`�������
V�צ;ˢ�t��"��&�nn�b��E��y� ���Xx�F���R��N�J5a`���H�P~=��Z���B+ck�L���~��ց�t�"<#˜�ٝ���,=�fk�f0�r�}���TF�jo�%��r�gOQmK�j�Jq퓻[C��5t;V��-��Z�s1��[�+�x���͎/:]��]$��p�n1��ޕ�eµڹ-�5xgz,Ֆ���ϗ����|�{�J���V֎���'|��Y��A���
ՙܩRE�a��s�p�W���A�EIr�<Ŵ���Խ�M�S�
����ݣHMgj:��ܵp�kf3��n׾0Ù��r���`�y=-��H���1p�t�u�P�*�^h����:���w��f1֥�a:V�T��k�N4D�#�s֜<M�_����+�I����K&s�=ͺ�)pپ�G	��}��zb�<���gI�7���z��Z9�F�ǖC-�1`Նsz��W�H�4�NQh�Owb��u�(��uI�Ғ�A,r7�u��r��~*'�~���0�/f:��)o��%��]����ݔ���=:��Ϫ��.�=N�/s�ͭyk��(�iڞ-	6�ip���>�:�~r�F`l�I�%�|߆��`�}���̻��*�����j\���%ﱎ�wJP���yc��'c�b[�繫裩���{���Gj/����aiֻԳ��'n�R�]]1�q;��1������xD��9l��!���3>��+^���)e�YPa��j>ѪgY	Ҭ�k{�5���@�-�ԅe�a\4�[bV�q(C�Tl�O2hx`Yi�s����}ir%�ǯ����/]�>��ư9�����d+��u#��VY��#hK���R�H����gv�漍t����~��bƃ��/s��ޗ�ٞ\q\�G�҈�cЇ�Y}{��؝�!�{FיXg����p�ecPՄ?�`a��z������VE���6pU/��k�V����롶Hb"jd�8zޗ��8����0���b�w�t���$Ѝ�+���V��'=����rvK�>��Y�U4oL����e\���<ڷpI����5�`�]��C����O�vLnߓ̍�^�6Lo�P,k�:ɜ_�=�z����4 �֠\gD���jje�7�.��jVw(n�y�E4%����:��47���Rm�&c��"v�G7�`1^E�`�g���V|Q����Y�O�]�T�N�l����P�V*�L��ԻJ�������"���D@\���Ŷ�5u��&��`�ظbt����#\�zp#�J�A�&k7U5<�&?읶������we��X�z�Yb�����C��,�o��V7�u�g����4�EKY.����P��|v]����6�N�IA9�f�d�fil��,w��wy�6�K��aJG�+�3rPv�B&:�q�I��!�,�i�,	�2C㮙��P�*%���S�v!��"G������Xg
�?���u�Y�w�or�D1Y�.gg䓼]>���Sz�E��z_�>�b+"11��q$v�gi�h��wk�~�����8�:�����:�pUV;��gF�b���rSd��g�#bZV��lN�{5a�TO(#�]s=��X�ϰ1���:�C|y���3��0�.�>��kRS�huЧΩ����pDE�T\I����������>R�Α=�·�����.�֚��g�9��=��<��[�l�#D�k�Z���yx.0�,_��I4��Lf��h��Q��TJ���D���Ό%2l�uTB�8^�0gǗ�O���t^b~;UJ�
�4�X�ܛ�����M>�w[���Xv͔�[6i�me�y|�4�b̜2acgc%�q�7��/n�+P�=��;��c1zJӶ�w����ĸ�#�H�.�`���U�Ag(��j�ul"ښ�;7��empn[�o�"��\#`��q���.�+�B���1����g���Ԝk,� �N�\��u�͜a�x¬3N�U2�t<r��V�*�Mɳ:�wN�B��4W@e�a=7Q�|�+9})<�}�qT�E���ڨ׎XB�:b3<��n�Ok��V�ۛR�]���;�Uq�-�lUC�;���8}(2P��*wlg�]-8�u�3[݄�\��<��������&NlΊj���;��{P����U��d��u��L�{r���x���-��7�"�UɄ����WS;R�2Ìs�h�X�aa��q-jg
�]2z��ሙ��>SJޜ碡\9�TPUD垔����3�o��C� K4e^1�:[A��B35����	�+��jd�Go%�3�h$��`�x��Y)_N�*���ʕ*^��0�9֏W��c"ۥ��-�eنِ4u��w��f���3V��@Ek�
^'��}���p�b�}(;S|�wU:x@��}p��y����r�������<ML�'�nzب�����
���U��k��v���'a�phQ�P�e��z�^��j����`y�M����-�\0!cn/PO��}�m�%Y;}��+}Wj��&�D��Zp�������H�zݛX�so�E9w�;��{d�)�f���7hJ<'2F��s7f�U��[\2i�Oo(���2�8{U�]!6�1u�����qOo�~���5=i>���rV�x�G�]]1B#=�S��[�أ�	�+�_T�vkm� Ȳ�SA/�C�	*"��n���d��N�[᫻w���yy�ZY�<R�����U�AH jvb�7,���yY���~D>��.1֝�Ǫ�u	L��á����we�}�b�vU��G%B��N6��9�����#�׼�iF���T*G�X��\.���M�&EY��[�1�� ZwҮʸ��՞9��KiU�\�kMQ�%���̾�o7�����`�j)f45];Qlŝ��+S�Jޛ$wm6��#��Tr���O�6�\�>ķ���bt׌D�<�"��0�t�㎥���Ϭۋ��t�gJ�IS�����:���D��P�5��7���:�UL�k�N��6#x*m����vL�g����έ�(�>?8^��!o[rwh���śPp����8fyYyH\��P�Z1{�f+H�ȓC�����;5n��;|l	�Wq�=:�s��&�yY�pk������X�S���aY��A�y q7�]�y�{̎;�)�d��(⾮���E��ñˏ2Q��#��h]��X����{v�e�SK�uh�E)�/*���
�e�I*D�IRaV�6��$f�M׽��O0E$�fԮ����P�h�Ǩ��;�Ǫ�=0W^�n�Oy�a��)ҙV˝�:J�3u6o0�̔�3yv�&N��bt��Ad�fŹ����fi�\�롨p⩻@Gz��dpב�eZ���������ob�IP���;�����登���"Z�r궫�<��VN�)��q���&�/oyWp�P�� _Rub�X+1�KM�4��������d�M�;E_ܚ�����k�>�\�J�n���tGv��	r���Y�������g7�=NFh�b=dm�t����Еm4�Itu�<��J���ω�l���6���s�n�Gi���;��e�������h���J{��k����%P�Lзo9cpG�;}��+.�P��tD.��`V���{�'o�w���=G2�7�p�b��|�1d�y���ԙͦ�ۭ���a�V,��K�n�)�ޥl�����JC�d��L���R�]���]K؆���yr�}�K�^]g��'�@؛�*��n�Ed����8�(�܌ ���f���#1HG1���Z�����Ѱ���|"��@gQ(��U�(�a��p��� �ew)sz��T&EF��
-�.R�h�w���U��of��'}P@kW<�H�é�0IΛ�{�K]\F�K��g.��u((ڴ��5���ۃ�4���"����8
��*��Ab(�QUUET�
cQH��hQuj�(�����eJ�R�Ub��UQrرQ�,uJ��UA��T�+h�e��b"�"���,"� �
��"���:eq�J�����TR����V(�̪�*�(�+-������&!���"*����("�U�1(�+V���Je�UGVQLJ+4iV�QD����PETc����TEb����(�5AX(�X���R�
( ����EDb*,F
*1UV
���i(�"0�
[`�*����KB�������*(("��\�5eQ���b���+V*,E��5h*�b��Kj�R�:h���U�QU�]2�"cq+lTA+𪻻��K���qrpJݵ�%��W	ә��no6	l�N�t����ĝ�\���l�[�d�4<���<��j%�u�ꈃ��F�	\�����$F@��y����Q%��ץ�%�5w(^Ma͡t���m�{�ګik�H4�\M)���lJ SRFW��4~��VDY~�ڮIi9�+�x��Ema�^+ �p,��/�{��4E	���7C8�	h���ٻǗ��N@X�e=5��p�P�b��Eg�X{%r[3�҆"P���_X�^�˻��ө���f�qі%e]�T=*/����8z�q��Кhw� tK�__�?-�}Z6YC�,�Vj�^�X�N�'�'��"VN� �ʞ	���\���b�se0�'b	����������v�p��PE���瀸������_��N.7O]v�d;�Z1#�	~J��r��ZɅ��6�a�3���0���!�J������yN�nJ�o=�� �j�_`L;�c�s�/�pVl�sڄ�<'�buyXd��W��̻�
�� t	f�scn�ę��3<2Y0�.s"����n
�吁��t}d���ٴ�/�7w���b
x���B��y�I@�i���S��5�]%wS����[���k,"�3�h�Zi��p��݇%�yW7�ݜ��#դZ�Zf.)0ҭQt��A_[xs�+���FMT�ͦ*�v���ٚ���$�* 8T1�&,��6v{�Ӽt1Qo�Ⱥs�##�!�X�F�[6U�n����/�`�.]L�G~J��<�����am�W�k� �{��d`p�n��-j��]�1"Ô˒�}=t��#�:���
�u�z��K�����9��U��|a^O:�O1���B5�ەa��� ��5�1]Zc���6��}6�e�(��tڣ�m8@S.۩
�,+��!!]�tJ����%���?\SC���_N�>��ӯ��hus�����)f�Դ$5ا$}�J�A��: �)��w��p���<��Co�a�c��_���C>�F	{����
P���Dn�M+�zҫ�(8����1Ly����WN*N��=x���N���qPԺӏg��01ӧS��R�J�Z����ͽl���G��N�r��W����e��v�����2�OU��(�����R=U�sɭ����̵��J��G�B��ef�zPU�2�:��5��N���\��	��u��9�W ΋�"�`7ț�+|����ܲ��R���mY��f�����/As��}�w�7{���;�;��i����c��Y��P�k�=F�]�v���� ����{��v��<Md��Ow=�.o`γW����ܠԺ��	�-0��ݕ�����K
�=rb��0߸z�<�7�ǰU��7����c��a��XmJêS�����f]�|�Q)^s|!�&z��I�B
��;[#����E�bԺCUÿr�܎�2��Ư��V�`�.
���3q3<<���]�֏�/���{b	U����cq>#��y<�=��&E�[!�[�Ƕ7Z�JG�+��t���g�U�(��Menck���ȵOF"DS}�"�oVZ���D���h1jXmi�(W�����D~�'�j�X:\��;����u�ߋ�8"�|��֮+G1��4,J�-���Kn{Z����U�{ml�f�ԢxU��[ν�U��.Ό���,���W`!��������v֭}�P.N�-����5)by����!�����9��_��=m��O�i޸k��e�^i�����X�/��f�Gr�U�)3]ēIKI�(��d�2 *�DdѫWy�fb{$�����Rn�/�͎�e���c�A9*��N�� �F�m	��ץm;7�G���Q��SS���Sy��};y�V�һ�N͖�!������}o��[�oM��Qi䚺X�[�Z�/qj4�V�CP٥�P�f��K�W�����xN�G�j�C�Ch��I�ī7��3|�!�r��Ex-���=�q�*}���JKD�����d�.������h!>��g����]!�G�7ٱ��eީ�x�oY4��p��}�N^;6�øYG
����,3-�\v�r��v���Yb2O3q�4>���`w?е�#��F���\sŞ��5��urS��+����WBԣ���b(��"�QYu�o[����3ҡ����U�5s�괶�5�*���̼K�^V�f��sL�*�ĝ�A��k�W�q��*�{y�<�v�ަei����h>rz��'��}��+urRX_#����� �_H	~�)bE@�%�7sfm��BM�k�Uv����7�2�J���A8Na�SC��g��E:�W-2�jF��k�M�l,Rb��~J@v�\pa�q+zr9�LȆ4�6��QGX���,D������҅g*b3#]2�Ѱ�����y��@����l/)ݡ��.�0c���;��.�M8;l_+��	:(���������F���Soǆ�ѡ`�48?-5��l��}�;�Uf6*�]�Ek/)J��S�U�G�m���y�nq��K�QK��'�[7�t3���Y��8�8�z��!�;Jq���'�����E�QB�.^���:���fX�n���ݩhB*�L���+�'Fϲ��%��wV��z�$�G��ƞ�㘬-�v(��JՍ�ֱ�sWX�LŖ�ww�6g;���(Pޥ�1U�m'�r���|�/S�fJ�ޖ::?Zݽ��gb�p�Ջ2e3�c�԰ᰥ���H�aJ�)�U�����+J,�a7M�����O��U�䔈�.J�r]؃��P��ɁR��\F����޵y⥲p�'-l���Rw+��B�h�^lJ 4H��j;�rl¿GD�|�:�{�"ߪ��srf*�I���q4+VK��,)����\^=�\战�|�	�$=X��ڻ�m!�̋sQ��z���lq��G��z!�/��Wv��gm��q�u�&�+��a��:�mMB�H�_��yx:�ߨJ��d�!����DX�#���|��	<��e�r�,�_�V�����1[ ��*�=����	'D=#��V�=�8��4pLX�D��őa�����k���ù�d����K��;�*�{v�������i(K���1Ñm&󱮮���M����|RnQ|e^�dm�����Ωy,g;��b�Ƹ+���Y�j<׼���{F�Rzr}v,t��xd;��~z7�v2�V
VH���=�P��ä��4c�{/2�J��=��%�X��/���Z�>S����0��|�.t�sD"�Z�1[��%���']E���@'��81p�����V���a�3d��U��uf��7{�i/��qi90���+����&��T[]r-9�Y:ࡱ�Ύ���3�/�g;��F��i񰺗"�C�x��q1�밎)�{��*�u��z��SlC�Wֺ䜽�E�y�j�x�nm���Ȳ��H"��چOH�ΐ�s}�B�w�d�����-/r�'��c���	<�7�@�ґ�k�点�c�� Y�W��z��WUrY��΢l1�^��K�������aʄB�{H1��$��Zy��t�ݹ�\��z�a84-�W�h;�VXV�:1�5�[�cK��`Tf�ʲ�3�r�X�`�d�ҩ�#��*D���Rf܊����5؍����;�0M�'�S�"}��h��a������.ӑ�ľ}��zdM]gV�W�W)r��Y�����c�iZ��z[����Zͳ��3�x���]@NY�!��'�.��;��^#��ȥ���r���^����(�����:s1��Ѣl;�
݋�j�vz�zr�����dY�NGdԖ;6r���o�:�c���8P�oK��I�w
���b��rs�"%���"���;f�Ѿ��G�����g��XϨL傭4�O	k���嵐ݘ)V>���{�U���;f���TV����s��yN)��U�r;y�f�,�Aº�����ZgV�i�F����yk�Y�M��V`��{���d�H�ڃ���o�eNF��|e��]�����z���y<;�܎\f�ےԣ��k�����S����z�&>�
�>����ccܵ��c�IS�$\3&!v�K�Nk-K��v�;B���D�A�"�W�F���"��c�>�p`�}���ݻ�&�1�{�{n�p�;�|y9��bKG�HV�R��Vw�\��v5����m�ܮA	9r�A#q�&0F:Ϊx��
��fPr�B٘�0�>�r��gFZo��NZ�a��=쉺t�N�؈sY#s�����h/�զ_�+�Ã�R�!k[�ڝ��6�h�.t�V�Ж�G�9GI)�m��杬�3*[']���9r��>��N�(Q�3@B��u���$�"��]}{Xk�L����@�t�'���<]d�8u�ѱ�oz� ��udL[���ǖ�5�S�1��4'r]�v"�ĳ' k^pS,�b�NUqXY�ynW<2��͋����\}j�D~�Eoԫ�<��p��ӯS�%��ܜ;Օ�����h��7�{;<U��
]��٭5v鋷W`!7	���3�˸�7���a�-)��P���CP�}K͌a�S�o�7��!�pr�y냍���6�dꃃ�� ���Ɗ�Z>��ۥђ�M�k��k�K�c6sEeR�w�C죻�=���K,'RՂ�F��xJ�D�?�P*��!��Z<�L�:�gY��ÁN���y��SMƲvd�ۊ�Na@l�6J�Rtס���k$�w�Yt�}.&8,��zn����gR}�vS���ɦc��Ğ}��5'My�u�Z�8X�PsJ<�	���y���K��=�qz]
�}�U�c��[�	8_ݓ�f1��%i�=�HP���������w���2���_��Q�N��+���#�pzޞ���XPa�:b5�kc�EmlW<}�oI��Lzl��fxUf���q'��A�/�QdȄ�yS�b;E����(ĸ#��.~Az6`�
�V��VW��J֓�h@�5m7���K��u�@�V����(�n�4jԼx�^�wI���ۧ���:���%�V.n�h.E۳XzSl��+gm�w��׷,��GUmn(� �Fv7(a�hhc:����*D��(!�q��=���ത�İ�YS�\
٦�w߲���x�2m�����Ob+��Z�q׍��#����]\�YA��DߢY�Ηm'�}t�8[	�8]I븄_,p�;^nC�:'õ!=I�V�j�Nga�n������ogOh�%9���3}�$��u�1:�!6���Id�b��|���36�����c{��gd�޷��']XsY�Ý}���ZAǩ����Q69ƺ1)���LV���gg��Z��3�mI�+,_kH��Y�Q�P�!��p�+zjVͰ�+�O�S��u�J�9GT�g�0�
����>�%�A�M��J�5�n���+��'y&�2����f���n.{.p��}!���Q�9���Y�mt	z�:�n�-����MG.3f�7����Ey��SC'��5B�}�n��,́�f�k^6o2�˧��lk��8�e^�f�����ge��9��9��#zǧa��ܚ��MTR��{}��n��b�8ޣ�7+�%'W�xY'�V��u�:�Uw�W7$�U�s]���E=�����̊�I��	��sU\�o�Wg���^�T�ے�^�r���kx�\42ѩ�F��4�n�\��;����Ee\�G��ʬ��ʋ�k���-hO+�9U��(D��x9Y����z^�7��ok���"���/ͮ�b�P~�_�<�3��D���z������+���{����74�k5���r=\=�ަN�d��V��u���W*r�/S[~����;{���hW�ui�@����w��|�NZ ܊+�4*s��pJ�[���ګ
8u�=�]8�v(o��Y6{��L�ډp����!^���ȾW�m�ĥe {�Q[ח;&��|��'4w��']z\����t��Psq=��D�;[B�x�g��f򋎕�;rN��D�v�1�k������<�z��SU�4���C^q�}��6p���C}�/�:�O��w3���݁$ I?����$�iH@��	!IHIO�BH@�hB���IO�BH@��	!I�D$�	'�@�$����$�	!IHIO���$��$�	'��$ I?�	!I��IO�H@�BB��B��LPVI��m=��@��v` �����������( �(�P P � EPU( *TR��P�*��J(�
 J� ��E%P $)@����
B*R� �PH!(H�M"%i�HQ*�UQ%Q$�R�%T��RD�R� P�*%B�@�i*��Q*���(�UT�EJ���DRPJ�	DB�R�*QUPU"�%"�U	JQ*U%I'ZD�QBG��T@J_   ��ֱ�����C%U$X�Y�-[�m�Ye�1@6�VԬҩ���ȶ�Pi�ڔ�������U���P��C�U PJ��JK�  b�Z�eZ�4����JѶ�Xh��XA��Pj�m�J6իV�SZL��Ѣ�`��5+dΜf�V��C�*vjW���R�)*�/�   	� }
B�(]����
(P�ΝP� �0v�(���
nۀ �B�(P�î�@ �
(\sp�h  n���
.��Q�&�iV���6�ҦD!*��"�֔)|   ^ն�� ��l��V�b���kP��Rځdm(j�ml6iT�ڃm���J����- ���`�jD�HD�QE
���R�}�  u�^�P3m���	jL� ҈�b$ʲ���U���)@���X�hѭX,�
5lZ+-��[MT�k
[f�!)J*UAUIT�  #�.km�5T��Y��A@ڕ�45���-m@leX�m��)0Z�5�l1�4���,�-�cLR����XR��T�EPH(�[x>� oK��iD`�)��B�`6��m��J�K6ժ��X���km4�b�i�L2b��� (U�k)@_pҨ�Im�UH����� 	�H�C0`*T�ǹ��m�F��j�� )iZ�P0��E�� JԡCHʊD%
�"��E٠�  #�ѥ�5P
j�6 *�� j��� ��/]TPPq��UT*Ķ�TR�hb�E�*�R�QJ�JB/   p*@v h�dV  �M��J��� �!�EA�j���5 -�ţ@��ʦ��π��eIT� ��F�OaJR�  )��2�D�� 4ba�J�4� ���R�x� 2 MD&(�0<S���_=k���(�h���ܽ���i��1E��U�ֱ\f���vc��R��9���$���BH@�`�		�!$ I?܄��$��$�	" ��ΖE~x�k����^PaEY��ƶ�[��J�<G�&�y�Ρ+�sQks���pT֪�l�]���W2ڄRz#�Գ��j�~I��	W�fD�ͱkTCN��$Y��3��B��YY�.TW5�*�2�?f�wz�;�kA����t��t!zqՑv�*��w��V�.��uu2��&�Z�Զ�'�ֳS&'Y��Jv�)���ָֈr7���*������EiYg_k�E�ZZ5ҨYˑ�7J�PD�xo-R��Z56��1�4JD�f���$ʫ�3\���n��,L�9IoڎJ5��j�5q�,´�.��mۖl��r��F4�F��^��IQL�٩�t!B�;
�ڂ�W�&`�J�������Uk��,*Z���J�ڬ�F��Mfaͧ��\V4�Ln<�W1I��,ǫYY�(n�nΝ�y��'Dʇ�r�˱BuAC,�v��fA�1(SR�e�������:
��L#���6�*�h�,m�|C��4�<D^��8U�mɞ�H�cY���Gѥ�����Z8��y�MVs1]\[t5��]���Lp�7�re�jo-����Ô!�����y{V`�PEn�̽%)���)�̰E2��A�����g0]-m�g��{\m;x��,��RyV)n"����
h5h���>�(�)��A��X�=���pպ�����*��woi�-sc���)4�� vR�CWO�i��~g����AGxa������*�HA.b�Nd̢���t�;"Ks`�v�nz�u�*�MS��i��V9�U`fV%yWM�fcH�0JbZ��K?pq�F@����w��J��}Y��m��!Z�&5�t�U�"P͙�eO*�8��,=+�e��v(��,�I�q�n m�o*f<ݩ��k�D�z鄶�֔#�"�\Mؔ�Z]��")�@���1�;�$��k7)
kFX(޽�$�ˣZ%
n�JϮ9f<4�]l=ݒLU����ݡ|�z��̢/O;��2��;ҪcJ�hXoFY�b¼�B�;�I��İ��8 �&ݚ��)�r�ekp,�9�v7UJ7�e%��T�F��Y-�f���,��E�
�ϭ��r^��
�3	���B���N�/��O]�7��[��eVC[h�V6���N�n�l�xB��C:� ��̢�7v���b_Т����3q��SU�Y/2�2w�("��GV����M9
���P�fγSV8�%���(��e٬�
ԥ[ �Պu����僶����8A8�CRCY��2��l��!��[��N�A��sxV�R��jf,�R,�e�hљ�f^2EW��e�ݔޫؐ�����U�^�ij�E"�<Oț+s
�N��z�^`��[ٴ��X�ֲ�%�L͢	wM�^�^Z��O���隌*ɧ���a�� ��;RV-��&��[����ʫїZ$�gD
�I 4nl���f
���;����+n��Q�P�M&i��)0�`�:�JF,��̕�T�T��l�!�J�*k-Q�����Bc��Iᛑʳ7p������c.�n���r����A�h�խ}��8Z���0�g�����v�k�����DU�] "Զn�͡���s n�On���!{`�Sw��jf�a:/h��-��nYp�w�E�ds��s���eg���ϰ�|E�Y�z��(|����4�ڀ�Yב���ߝidS;�c,f�2Q�̖6��(�.�����)ˤ��jw�㙰+c
f�CrMu�]�[cn���Y�FE�SX�LfM��N�!=�d� :8���ۢ�"2n��
�R4�0K�܅���V��f��;��Cl�+w3(��.����Υf��O.�{�*;t��K���n�U�[��0��ӻ�nȤ*���i��"Gh鶥<{�J���A�-aٔ����5c�2�l��-�M�N�$ �-�[��ѡ�YddM��]�.`��$+��e��Uạ���,f�S0�@�tq-�Kt&^��I��Ԇ�e��ĕU1�Hݸ��"E��y�2<@�t�O.��/ls5]h���jc f���SW5�
�m�̰2�ݧy�^�����:��,`X ���V�U��x���xl[P�2�
��)YB�vf&��~�Y,��A�ˤ��+^�e��nV< ��@�6P5���{��Qx	ŚJ\��.���á���'r���)f��Ԛ�'0�㨲ʂ�+4wNd�8����|�ըF]��:4&��p�E�v���IH8���BfTl�V��*�1�	�cIvtV�cj,�nZǆ��Ժ��SY�zU�@ǣJm��*��kF��EڴK��ɓu@f��{�lIS�MU��[eV.X)`��H�{�Z�� fν�2�jO,��m�/�H*���lht/6�P�P�6�f��ec��\H���TNށX퉎�N��k@y�^����a��l@�i4�^��$U��|lP�J'����.R�ڠ�Y�^��X��2�inn�k���g��9��FV@-m��(TpJb��(��5i�uI2(�2���]7�*ce1W���)�4��[�7�۽ʶ���жvk·L͢f�%��	ܴ&c�/12M�Yu�Y��l�,�<F�/�V��6��fe����x�e�&
D�ҋ1�r�LIkh	�fl7[xwt�-�o�ZN�3�M�&���/ɤ�;�=�j��6Q8�V�� ��j�,���/]��]���An�z���9tA�"�[�EZ�1��ˮ@4�(7�a��s�3s�`Z����
: Ѯƴn��͢?��l�J��b��ߡ���2�wX����l]^=��K���wCJ�C,U&ڸl^�쏶��R�"M��QC/v�Շl��f�AW�k��\�Xn8��{��Bme���+(s*��8��ֳ�c.��ě2�X����:�JM�v��h`$SY�2�Z[����_�M�Sh�k�齖^+����Z�VunG�4QN�̶^m����FN�d�Z��:M&Q�S.�9N�.�7A�t�#N�Ѷ��d�_.�t�a�F��n�72�:��jh���Jm�ݣE8��Z������N���[ķk�l��M����m���$�.�HEz4c��!I1�HJt�uMt�ˡCq8u|�ͲQ���u�dä|��2�4h%W&���mǰF�R�^)Z��rɳ��#^�.��B^��lR`&����tt-1�EN�����b�j,��tʳ\��l�%Θ�m��4�k�h�s=?e�°E�u;+7osEGN�X��
4@�&���ٷ�QX��(Rd��^e�r�рݪ�5];�e�P�5�Î�&�b������Ѹ���;X��:ͥ��8+�⮋�9L0�YY,i��52U��[C�XB�wu��q�+f�ɻPjy6T��؅1��n�Z�.�&nԧ�j����B�^B�=Lf,�O,�2a���w�m�<x�o� hb۹7Jù#T�B@��`��VeIx���a�٭�<ܤ��ـ�����m#��M-r}����ŭ��[^;�a�Ŵ��5qE>ېK:(e�I��4�Z�+9ؙ*���WOci�+�!�fL�@\�H-���\Ȫ�Ԗi's^*;X,4[ʳ%e/��Y��R؝JQSq��]
T��N�e��τͽh�3�R���M�֗��/su����2����2K�F�e�����HC�(�WB���ۮd��� �+I�͒Ѽߞ�n:F���"A�I]`V�$6ʛji���n����fP6��3-ض�w��dHSu�u:�R����wX��YKQ�Mٕ����+l�:�f@0	lŎ�M�R����Z��l��,��kI)ꡃp�,+�6jkGnzC�ma6^L���tE�V-��ژ�Tn���5R*��9��2M��-�&,�6�j� ��3c���GC��oNT5���9m�F�;�ر�$(Y���lZR[D��yZ1���P�s!{Z���y�-�Yf��B�aU�(�e�J\{ �K6�ԭ�Pڬ�-��V;[Lᱨ�J��\��f���v�1%�Įͭ&,�6�M��47Eާ����b[�Q�&�Fw�u#�n���C�KP.�Mgn�t節�«XI�mT�]D
�2��,������p�$�:�S�2�L/T��0퍧A۔N�]Jj�����1�Se�\Ӧ�n�aL��E�A|�+B%�T�8���t�P� ���А�Wi�OM.�u�"�����:��H�H:ɖ�u��dZ1��D[.�T�� ���Y��@�	��t�DS��uz���8ՆmRĪؠ)�:Ƃ�gRz�^��=�SU�Id7��cfkj�;yf"�U�WN�ζ	B8���*����3/̤��pj�i$��T�p�h�h�e���Y[��p^�҂��0SU��`ۙ*qe��E]��x�2���I���xY$Բм�,��yCD����,戎��W��������/XX��o	�X� µ"���E�4���i 		��T��ڥ�+��-T�4_"���c�:��.�LRr�+c���n�iU�6�����"��ŧ�me�\���8a5�Zqn�1���vV0b��U�Sd��v�&�Z�b�F������4�NY˰���u��D��-X#���yx�蘷(��l�� �֜��T�Œ�����&D0��u��Uӷ�)�()�����ka:%]��0=��ca�a,��9Rç�VBa�ff�)Z%h�f6�J��;������4�<�M���1��8l�.�a�v�:�}��5��!�p���ܰļ7F��������q]�c��$���l�t :;r�����&���u��i��/R���[�m!CyV�X��e����v2h�z*��Ѻ��M��ѽ�
�f�f�=��Z��nd �K�F��G��g*����a��*�v�F�72(4`���L��d5�Nd��XM0�Y���w[��Wcr�\��x����h��Ĳ�[MA�^^
\]���mu�4�PW^f,ǫ6�< � �X��x-��Z��n������[��'t�̑�h��~��-/T�w�* ��:�H���n������ӧ�P&�;�xd7�nc���on�z	
���.j���Z�+nY�$:$i;�D�΍V+ʻ%lW���Ot���j�B��bN�7G1l��z>F�]^ũ?��q)��[��ݣb�EMe�h5�0n��8�����y[�	�h`]�iY���Z�S>�n�ݒ�PXr�V+�k
-K"�XR�4�V�ɋ����m3��`w6�%̊�9g�*�κ�}���[u6����``�o�g��*Ɛ��Ш��Ja���ձ�X�f�C�����-E7"����yf� ������*ܘt%`�.Q��+�����y2	xbJ�$%���C�{��tr�KbT��k�R��L��1�ʕ�J�:=�K�h��z��W�ng0#�/)V�v�_�ܨsb[�~׈XwVn���EɻtT�t�fL+'
�Qԗ�Z�v�W�UԥI G�,ں��F����aj���N�W��di�l&Q����4��u*�-[�ǎj(��Z���>Wv[U�,K
h"���e]ن%BJ��-���o~,����S컌Fcۺs�M��w[P��uy�4�ٵn�+-��g���Z����ky ���"���a�x���N�{|�*���؉�]����We�Maf�h	^��YfS���ռ��ݥŲ逭�ڻ6.�n�B�aV�d`�X��'ox���GU��OR5���3��d�����eڧ� �/)����skbt�Sϖ-�y���kZY��Z4S�r�O+�u�Ř�-�)�[[�lh�A0U��*�;o��V���(*��iJݟh��=	��Ei�V�]Y����n�m��}ս���|P����i!X��F�d�Km��EКj:�b\C>M��V��Z��u��D�Ѷ^Չ�YU,�
��v�9g .�Wbc����ʽ��V�*�+�����N��S��h�q��Ϥ�kXׯ ��Ի�ԙ	aucdR�"����v#u���=�e���&��1k�Xut��4k9w�5j���?C�n2X���̑ĝ��٧V��DV�cD�v7�n��@:Z�%Ƕu�����ӭJT�6��(�雍�%C��.��ͬ�[/LN^������F�-�f��"��n9YY �v�-'��z�_�[2��F9q�l@�`���!�`�x��Hqd���{$�u[3���:Ôq���ۍeչaQ��f5��L63j,���@�扷�A�����r�MtN����Ar����dֻ2��v�āT����N�\�t�|��+O8���~x�4�rm�[��N�^�2�[q5mL����� ����fr����hU.���#��W�3N��-g��_��+��![c@�4�QK_ ˷�aWi$��z{�=��n��y��hat\(����)���7"���+�Cen�9U����-y��:�[wY]�Sy��bGs,�ֳt6��T����"򒗛7�
�)�۬��*gNJE7s%f���V)��*�iP���*�l���"��Tw ̣Y�N ��ՓnK����ch���ߴa��$96��m�ET�Yf�7�V,(j���h�� P�-d�ަ�mktq�`cI�#���1�`�Z�	L��.�}�PY�[�09e�iڳwm�כ!�C� �#�K|wV��H�Af��'��F��rACs�s	O�#�m�Eӓ	ub,v�E暽,��U�X (�c̢�6D��h��ȕ���ݽ\-rY���d,��VV(��K0N�weC%���F<i)���J��o�_�ho8��dK�ʛ�R�2j.�*6'1[��z��q�vQ+)M�u�p.���������ܡ�*ӽ����5[A����W\`�XV��s��Y�W*�g��H�nJ�O�44L�N]��k��o��;����� �k������iK����/V����k���׽T�oU��!O��:�op�8З�gʆ*�E�ؚ`R���8�Q�l�1|w
��FS�va��r��qI۴Hl�a�*��d�Ң�u��1i�&�ۜbr��2`S���UugZgtwgҫ�M�T��7��ݒ��8e�=��W��ţ�->;�+}I�9û�K�p��/H�;��������0N�D�bfF'[jJ�U�J��50=GM�1#�j��Y�n��_:ʢ/��BhFœ�7�Gc��6��i��jV�pJ��o�v�=k��~�q����0�J��ɫ;�����e����f��vq��_:�y�T��i���;�u#��򷭃��I��6�>N�����ǎ�B�f���&,a�՗;�՚�&�ֵ��Bں�1�w���IK���Ԯ�U� �:"��km��g\�q�0���yu���)��1�A#�[9�[�k,�,>�h�Шf�Y|�h��5aSTq�Cl',�3��;(�Jw�kc�p�5,�Pn+@��ц�<33Bk�m���սO>�0�u+n�bT���ݤq2s+�� n�ކ^�j\�8m�:��[1�V�>����q���x�m�k8ڰhZ[�tZ��-��OAw���wӷ�j"O,�L�(�#���N\<r�Q�Gz��9���͑���<���/�NHs>��TŻ�O�+ӹ`:Wۙ]`��.����h�Z�ڒ]
����h[u˺!�SO"�#�@e[C;fIf��v5�K�)������0pʝ%��j>ɺ�u�e�7��@Bʔ/r�Uљ����
c�C#���C�֋s2�XS8
��tA��l�,F���ǂ�:?4�HT�5��%��=���������R܅�b@� pw�M=n�3X)�r�n�X��w����Ggk�:d��8H�Y�i$����hlѵ�yWP�w�zu]�m�3������fQ���ˡ��üj.�/��4�[�eNe�B܎�9 쭂mcj$�}��pnfp[P"	e�`L���K.qU{�z�Ы���d�VRR�4��im�V���f��pQ�s�8T�5�Q��!H�̭77p@��`j���}g{0g��3�iӒV�(�_	Јz���˚5�T���������<I��z8�X+�y� ��z���:��9��%�x����2V"ߝ�x�N�9��,@u���O.u����f�\o:���D��%��S�K��0�����*h�]K�5,'�+h��I�Mנ;J��7����%۱�'���K�R���:���r�Q3��%��{x���ɄL8�������T�	Mf,#����
\��ޗ�hƞ�9mr�T;Q���͙�(�7��7�:J���#gh��"��kk�����P�*�K�����T�룱v�����rp�^�5�%�hj%}��P���3QɘzT�����At��I7ʀluj@��8�m��6��w:�R�k�d�4Ru̼˵��+ot�u��4��d�kYd��9:8�Wz^����Uw���
zQ�/st���㻴eޫx��,��M_b�H�f�<�m�w����sie��U�4�p���oϥ���)� jJ�&Tc�C�pe`���U�i���(:���yq��c���:��]ƙ��8`�ǂ���<1w$���%u5X��Kw��1������c] ��Άg�EM�.��7�.%,��@���Ŷ6���\��^o^V��.G@{��r,�v�ǵ�"5Z�=�}z��[6�N���&Y�邫�+�֔�����-c[T���Y��VWA1�K�GfK�+1V��{!Th���]�s0E���B� 3z+��[A�X�m��1X.
7���X��*K$^_v�h2�n�v�ͩ��Zbv򔩹���%Хt(�:zĐ\����[gIح�F.K�T��P�k[����#�C|���rبR�1:�AOU�H�y�W�g�Z��E��՗� ��r�����<맧xv�+
i�%�L��7X\[�@^��xI�J�u�,y|��Gc���--�� Jĝ�$�;e�ϙҀ���9��Tg.[�kG1b����8�4���l�*�7��㌔�	��i� �G��ki����s���r���{�`w����Ok;��:Ŏ�8��m�E6�eN�F���xg-A�̵�%G��/krn�&�5�[]]�,�5���ʪ��(��&��5�Ƃ0��[S���M�ϯt�,�k%l�ÝH�gq>֭N^B�*Z����-5�jX�ڎT���b���!vÆ���dw*�Lu:�^�4�Y�4\�hPzo-�U�mԠS]Lr�Vv��)X�|\��{��(�7G��<���*�
�E'��q;��%��nӃ�����_":ƴ���L� ��;)ʯ��К����e+)��q�L��0PλL�����y��o��V����b��8�Q��D�C���35@4<���U�ܮ��&��*�S�f�K���	�4�
Ή��q�q�7�և��p[b�mG2Ô_%�9��]���R�[�a�ٙ�0�&a꼭���9B����GJ�9f������h+���t�oVo:�J�XC*�D}�[�U�������%M�=�7V��WrE[|����r�G2��׌TM���3o*t�I�y_�=)xa.l.����R�(�6����;v��,'Z�4�Pi�:NV*Ⱦs;�� 1k�29m���Q�]��<B�,��qW�X0$J�ʘj�ћF�m�7�֡*%���W���b���!��p�3:�`��F��yH�Ǒ�	�"Ɖ�%gLᔤ�]�<�h9R�g7K�WR�Q,���)�ֵ �[��XTF�[}h0p�IT �K�\٨hS�\V͹|�U���[�R4Dz>��P$}��Ceb����'2x��:�t�ޭ|xhZ��4����mIV'C��LU�+�^]�X�n�8B���N��_h�n�6��ԧ�t�#{O�����q��O�S�2��,����;Z�76�����;��-$R�D)-���v�����.���F8,�ymqMQ�I��w�){4�B4s+����ci�Cp��l��;x���o�^���;Xj���ԝ3�䃹�V2�ߴ��i��ό͹O>Ug�X��+l�6�ZA�5݉g����+�eI��������B��af4	����&���9�+�:�vz�Q�L��8��4�#7(ؕ�����9W@m��SI���F�5��/6+�,S��6-�QY��ܼ'�4j�r�5�Ӟ��Vna�)"_*j���jm��Յ�.�s�d���;�A4���uά��g����YXb�ĵ�l�����]X�튓�Ң����ʘ/���*�L�W��~c��bګzLR��`��T�H��[�W	���u}4М��8�It��F�IR��VEze*-i������3&sJmgk{]6����vB���b��*u�g%���2WAn�%�t ��� ���l@���Cp�J^�NE,z*KYܴ�C;w������
<� �b���x��"[܅�]��WmX����ݛy)`��\b]�l[��2�us(ŏvը�^٥�)�=��q��9����B�7N�z	�=Iu2�I��_96��A��A��u'�V�4���`.�`���	�1��%��ڱ��!�v����\Z^�����<HHܡ��N��sUX+�#\sG`�m�:w�����ɝ}��\uR36��vu�q:w\v
L᮴++/r�μx��2J-��Ҍ����>ͲH��(8����7ե��Fm..���E��f,J;��9|�Yٵ�r��o�� ����]&W �������2ŧ.X�j��7�Y��i�#s�97*K�~=��V��ww����-�ee�i�2�[B�#&�.�gŸ\�:�cV� ��w�k��	N"v�ڌ%����l�)�mfj��ƃ���C�vIH��t��e6�i�E��ԡ��0���`�nX�
��bN�P���光�s]���'y���Y:u�j�R*�
�1�i���ф��WB���6һĺ��v��WX�=�ʵҡ�z���)���9)��]�A<�{���HR2n�DfEÌh���VI�W�9�'�SI<g�9�D3%)��Yڍ�
��i��G}d��/M���*�SS��G8v�v[oˡ�i����­��n� �kf�Xn�v�-�-�8��\�C{Y�6k��|F �kh���Y�we�E!Q!Tw;Gu��"U+�T+�c�|�U���r�l�@1�O2�Hy���ډ���e:S�T�R"��+���b���YaWe�͵G59`XC,ş6�h�F7�e�'�C3v���̋6�Kvjk�4 ����t��w.Ƌcpܽ.�vW+�NP�����d�x�6D�2�Iݙ��1o[U��B�R����p�`�oH��lɠ�m��]J�����U�t�V�ˁ�؛:-{��7|:`81KGj�vNFX����6��ɆZb���4���\��'^PÐL��;���ֻ�(]�սf����銘�+�X�nD��vM��7g�iU�+�Z/Z)ƹ�2����ơ5��]�*<� ��w[�6Vq���"=P1�x҃��wR�Ʃ�v$�V�Y 5
Y��j>w��8V�*J07kG;�G��hh�0m��;,���"/N5��N�ظ��������0Eю�XF��}m���D�*v%M�	���5���A}�^�Q�K�J�xXTL�V{@��S{5�WM\!Ȍ=�L����k�oq��(�)Y]�=���<t�j�wY����>8�<@U+{�p����ތ�I�bI��X�tIU���z�5���K���ڰ���q����uD~eR�Cl�a�t�ݰ5�xOt��iHp�����}D���yMZ2�Z,N�aM��u-J�g�:ӧ���P�h�7�ӣo*<=�1|���܈����F
�e�F6��� �r`�M=���9R�g-��@�����E�[�3?;w�]�j�j�E����T�ٝ�jV�.��,jN5�6,�փt��# ��Z�G�;��m<�U��/HM�C��E��!)���L��)[�m���o��w��.�o#�'�m'��`u�*�����<���g(¦u�n�͕l�[�6�<WC���@2��u��(��A��F���3y�:����y��"��`Y*��Ymc Wt�%�N@4+n�KC��Z̛��4C G�Sq�����f�P'h�mIW��n�關�Z)�b�2��������V�;�Ƹ;�����^T����Dx���v�7�+]6j�r��U�r��q=��֧��[���ޤ�޵�]+c�t�<zѳ޾����gI��'r���!��ܣB�Kri�\� �/1'Z��ji�9Pf��R������\	M��l��\���:�a�²n�/��b9�m�����]n��Y�:��Ӡm����h����3K�2y@ᩳ�ↁ�U-�1��f�ݫ�N���rj��#��GyMWK���;�2�Y�r��WC6�Vs�C���z���;@yȃ���|�9N�u�r�+0�V\��MY:.���=���r�.��i ��5cR+:�oi�n�����W\l�;E�j1z��ؑV8�f��6������''����=�Fr�g����j>����{��ڡ�hϰ-�� �׻�5wk�7��P�����qa�lt8�d>���!qt���)a���ayXs`���[��76CsK2��v�--ХY*�G�5aY[b��v�l��!8��*֣JN�z^hF��X���{uu�`���T�#��hћ��w��SB���)C[�������%��]^��9'�Vh|������T꛶��J�nb���<ͺz�!�h�&�{6�d���&�9���a���Mt3��>p�����2�2��)�舢��z$s���h��"��3�`j0VF����u]]q��,6;#I8�B8_���qS���M&���w���<p���)C�sw~P�L�J�"��i/9�d)�S9�e�-j���˺`J[����A*�^Wn�02u���k�z�8����T���s����Kx��[�o�g��6\�~�f�I��,=)E�fa�����e��Y�����|�N�d�7�����}�K���g]��M�NN�&��Ax�,P[F�#x(=P�%wr�kkF��Bھ�r!fU�ss��q4��>5�/��O%WY��~�]���ح�U��f���}f:oJ�)�X(h]=�vݑٲ�i؂�
Ĭ��v90Q��ρ;ӯTWa�v�f�:�I+7��u��#�Ϲ��#g٪��T����:4$&gv4o_�z�P�A��+KyI91b������,�{���6+�;7�m)Yi�g�WJ0+"8#g2R�S�'U�%�:R�����O��d{
ؤ2J������ ���	$ I=���W�����g��}���~�;x�M��ϚhPq��ε�"6�Rp.�.t4�;Goxv���m*S��'�f��98��9x���5]ZT����\T�r�[�3^94�bjkOT�2�[u�O.���R�к����n]��zq��nR�U��J��>����s1��T�������@X(�X�&�(^��e[{t��ڹ.M&cNc�T2���9�ڕfk����B�*S5��v��ㅔ9�if�S�B1(�D^)����D��6vn��{t\ڔ������Lg䔅�k9+�"X�J)��iL�94S����Cٵ�oK�2���R��'>��*}e2�Y�n'KS�Ǩ����M���jJ�[T�#2,��p:ᖣ�6�	�X�^�꼹J[�t6E��#-��	A��c�e'�|������
X���̺Og  ��+C�*�j/����v�Nm]p�D$�qN���*%�%�J��ҹ�
�nƮ���n���)�Pm,�靗�qD���z����	DT�����박*���` _e��j�ŗ뼸�M�环���[+�
�7A2��+E�����/�,���]b��]S�o�^ܫ.^��/��Z��4�Z�p�Ok7�jN���1�[�GR�ܘ��@i�â��3v��|Ⱦ �¦!N떹����ֽh%`*�+,oR�B��c�]�wdn�#fj	R�X��z�|,$��D��/�1͐���io;*"��h^N]Jj1ބ�����#hC��nZ:Okev>�FÎ���k �j� w>[�Ù�n>8L���n�y�K�sX��c���<t�n�|�T2�tjq��J��MD�f�x�#u
v)n�V;S�MU�����giT^v
Ss����F-�ˣ��u���� }b�U�f�tq���,ܴT�����52p)͸�r+n��k�n�Ke����f�ش��������`�+��E-G�Ǔv V�ҕ�m<U��V�L
��K٬�05�0�/A#���m��&��y}׬A�m.Q����ʛ��r%+D'��[�H�L�j�0��Ĳ:=�́ު���67ih�\d�(OE�'� ���dPg�ݝ��+x�zuC�ˤ�������d�C4U�Zw��\��A���z��%�)v�����Hu�����R��u�v�;��q�_$X.�������;����\b����ݦƜԎ!:�v8�E�H-�5��>7��`��P�	�r�ʵ觬�ĭ��y�wס�p��Gt-��.8�w��i�Ϋ�Kå�B�|�e�R�c �6wJs�\5:�d՚=�En�T�;o]7�4r�5��Ѵ�2�XM�� ʼ�w
S��Y�aR��Pڗw`��ƃ'!ٔ�gk�f��2S��Jkmp�*����t@�8�wnv��V��GwB�'�x�u	�U�S�ܕfg^�6��%%�Ȯ�Ԭ��M���n<��ͩ�VuY��P8U;7zN,|��������P���ӡ��ݱB�w�3QN��V�N�,���sVS��N�kM�H���[��+E�˃mf �I55�I�1�6���Ċ��IQ>��6�8�jnr�ٷ-%�N�R�R���ջ�R����\�kY2!��/� a��!ًMΫ�C�6�@/�Ԗs��>�YGBb��Ω���f�U�h��[�]�v�ªA��* �,��<V�k����ll��	V��n�̳:�����L���/#�����KV�"�g|��A�vWgu���3��Fk���G`5���V�l�%*���g\-�A�����X1��}0ܮ�3n��	�=�� {jqi*c�F�yjwvf��p�o-�)������m�At;Y�m�"@�g�.l/���\�Y�E
��g۔fe�����0VڻtvӤ�=j�c���7���d)��L�V��6b0t��sIҁ�����t��F�91���h�g��(�ݝ��V}���w��N��u+{Ka�C	�Ӛ"�t��o��)}�j����*r�d���x�=�k����w(h8)#�n�F����F.Q�Y�&������Ւ��eȠU(qV� ����z�ݜ3��X��ʌn���h�cu�<I������sCK6Sqټ���.�4��Ng�v	�o��Bf���҆�N���`���PX���a?jU�"��c�����AR���샊�r�uq��ח�|�n�YҴ ����;��rmek�f��[�2l��0z+|�1��b�ँ<&���e�;ބ9J8b9��E��<�#`t�x��f�n+B��o��7��qh��d�'n=��*�J���io-gV[w!�D��Aj_v�8�U�.:���:n+���S�ܫ^Z-��n�T�̦l �*�,���[�t(Ws�ЏF��'nh��eO�*n+$�����ϕn��;+���}�h����4���j����h/"��}V"4m���L��ɆN֯aκ���"�%ѹX3뵦�EI���ae���3H�y��g��g2����p��t��v;c�;k$Ł��'m�jq��Z2�V�l!f�wӄ�g/��4s��5�E�dW���I唚���/*`��V+�K��/bT(�md=����CvV���FM�v��G���9�T��P���f����s4b�ky$ �����7(��nQ�`�т���� �y�N��}�X�Q�r��cl ��f05g%��Zޅ�,\㘈���+�U��<�[�s���N��(<�N�+�u��r]n�k!�5گ�J�)�X�,��ʗ �\,�0�>5;�n�;�[�
�hǒ���ጓCI�{)3����f�j�^Ͷ�S#A�e�\��@��#o;77D���4�M�Z�gOCX3J�+}��Pn>��i�ӯ����[	�oQ��	G����uqY�ն�Q��<�D�0P�r���ӣ4r��C�����UՏ�u>U�<3��J�Lu$�]>oB}up
¹v6�w0�\�1V�nnQ�;���C�����;��[�SK-�+���,ry���˧KӑQ���ަ�|ɩu�U�\�j |L�R���5[�o1f��urv��Y�����|�,=[f��ƨ��1�����4�	V.h�&���x�o�>gh��2���gsE\O/�e�q\7MM�).�SX�Ծ�JY��n�V�JyCA�4](.כ8٭���ti{Y9�Ò�^nu���$z�0�V��OnQs>ި ��,�֬�0�mt{���LxM�{l�D9uj�uM̕՛�8E�N���;RM�\ք#�k"g�w�����D��K�]Y���EP=����Ƽ,�s�h�|#c��L���P��k��iջ�؀}���mn��ʆ���Yf�4�8=�y�Vx�?��>�����T�aΛ��uim���j�t횇a��ea����Z�Y]�\�;�FȬ�D�'$������X$���3+��9#���xU�0��{���z�*�R�AV�zu���4��+9gb�cCP�f+[�V�F�Sj����hm]n=9Uy���a\d2�(��[�)�JH�Q*<6�.'���Z���ܣ�z4�a��lW��:�H�Lm�ؠ3�l�V��j%�E'�v�{�/N��7����{WI��w3L�����~1i�[K7��S�a��s��Vd武]�6-i��Vo�I���nuN
c�B�#@Q�8��Y�/G:�KO����h�;���B�9�ZS;m#���*ͤ�� ]���Y2�:�dÀL|��R&�Vцsos���4mU��Fk�X���g���2ilnn���
�/�RL�Ӡ�R�^m��<[��R�c�%�W�M����9`qֈ��Mw�;��>��Sgj��
��k��M��Ci�_Gy;qc�
�<.R�-����jm�9�3�Z(:�}����\ٵl�M�MD�s��hǄ����!����ӕ�X/�ǘ�n�K�OK;j�]�w�ޖ1q��GG,����lb��͊}���Fzi�C���k0�5R�2��u[��Q5+f�g{�58�{o:^e���L��$�b]�S�ڗJ���ћS8emiԹ��]�.�o.f5[��5]�F�}�˴��@f�T�5�-�ĝmZ�6v㏝�׵�ܢ�<m�[UY�l��P�oP���蝶D�[�f<��<pM8�����v��핻%�f�9�g+hi��^І�F%x/6�p��O�*�a�[���N��avܜ5���k'�Q�c�AǸ��f"��=��ˁ����Y�0�}�U��IZoT{��w\�Wk1wk0��rL���G�[�Gc�yܱ��{(��g!�y�]\{t�������|:����f
MI�9�d���]���)CYB�U�թ��m�L��
���<* 3��5�"l{�*��%�e]��v��}+*5u�O���,�D����$xc��v�����)�8���ӛF�ŧ�deD%�Ϫ�O[q�Vv��[wR�4��vs���z��LT��&�7�}�r�ŧ�PvQ�a<Y�2��\Ǵ\�j��e�Ωw�ĎU6h��bmf�GJ�6J+h� �)w!��1�I�T��0�к@%f�l�9Y�ͣ�J�W--I�Z�8���\9�&R�G32�\W���nIg����&���.�V�ʊ\v�ۓ�&��m1q%+Q��YQl͝mj .)r��Wt�b��Yη8�YR3�0�엩>������Un;��g]�*:2N���<�[�FQ��U%�H#����\��YB���h�ol�}O�2��,Ivۺ6S�B�GC��Yц���6�r��I]�:V#+T�.\s*ţy5�i�jGM�����)��(g`���P�N�(ȝHvZ9J۾����T�#+8O^,]�������i�I}a@��'yZgQ�b���-����am.����q���BA�a��{*�~X�B�������#*��B�v�T
���xb�:�w
�Vu-7gi<�{�W*k����S�j���jQ�06d��*Zm宱�<Z�˫����W�[��q�Jr�e6rf*��PP=q�؂G{��3cXkm��Xr��t�z��j�yc�Ⱕ��X1��(����J��֨%��xKt���A����(>h�����R�#K�IV]��s jL@C��ǯt۔�Vm�mk}R���+2��%\�t���@�����e�*Л�
Dm2 2�#AԍiQV��oᙈΫ�r�|�Θ��hp
v����jt#��L:�y�s��v`�wcڎhl\����� \�&��+\��cj��Mt��s�	���6�;p��Zck2�#J�n���/.�QM��/N��E%�@Gv���X0mE��f<FLyP��:��!b�[�0�/l���t:�3�fq�5��`A����߹��$5{ٰ�z��H��;�ZBr�c@���X�=\�ut"�l��Qe���89@	빷�V!;�����q�i��<�F8�<K/�0R���%ݸ����7�ˑU�;�Ck\.r�î�N����**nt�f��� ��6�K����-u��v����ɣk��W,��2H�_ �t���r��B�^W%��x+	��]2>��*+G��gPk�F��w[m(��pm�ycv�.���A�Z�9���[�,�<�qٰ�J�8Sy.a߂Ў�r�mw+ʵ�����\���K'+a�2�]e=ˑn䜆��+Jovw_>� 7�L��C]�Oeb׆e-3�M��W�?43���
���������3&�F�ݠ*�Zj=\l#ީ�^��pK�*�X���UyK7woFi��q���6���$��,JD���x��ӄ�6�h;�$v_�:g�f��p���t0v��q	�Y��۫��R����|aYY,��Kz�;1����u�ĺ�E�ɒ�vi�%tPa�v�r8���[�O���(��fż�8K�Y��%�3f�Mb௚��J�ۥ���^�ld�2���+
�U�/���(�un���͏�Ѱ��]�Uɕ��S�M2�S;F��$�1dt5qQ��|[�(&�;ܲ���Ѭj˺Ё�z���\i>�%�r}p�ܛ�ܸ���w�N�J�^�';H.:8a]9����jv'��E��Т^Y�[T��[O��D�X@ou�v��0Q�-i��Δ{p0CSe�XoRծ*�Yjڭͥi��Iʊs���SW���T5ظ���]2�ƨ-훪t��c��gQ��0W"2�\:Pp�V���J�g!�go4+�ڏ��LЎ)���;œ��%OGldK��g��toi��[E���o�@T���;`�����ci���U��>��b|]+YN|�*q��^�����R)���[?_j�U�p� d���R����b�����[�Ԓ�u�r�����<"j���G���
9�lT<7k5)�K�n'�I�4զ���Y��ƈ��&P��@��U�*��z75h�oL�7)wH_vU��
�#��]�Y�����\T���Jo�ޣ8v�'yk�<fM};d��E������*|}B��J�ݢ��`��y�4 㕨>%��W6e���GvU�6_utä��cm�`6tV`���Wmv�U�;Vا����;�B珮�K�\&S�e_4�U��p�a�1�Z֪��.T�:����ړӝ�W��Jɖz��d-Э�VKnsy;3��=��uٮR�S�����X�i�ܫ�y�]'E�ϩ�ZB�Q�MX�yK��X��Z,�pd[��ѡ�m����\�q�yX�;�����iu��BH�T��/F���#������{�e�Ǖ`������3�����Q:4ԍfQ��q���yQf1��x��غ�V��کP��m-ʶ��t���W�
$��!6��l��6A�G����D�. ,Yw��c�_k��F^}��2��[%'ܲ7Y��Ղ��ݾ:�%Ӗ���_]��ABk���T���C���C�R����a�ĵpT�P���!�/;-i���$�)YT%91�X�*.�;*J=K��VIeC�ū�\nFn����@���
��4���{��k0
 ��e�m��#���6�U��}�o
Qq�v�����V��ۣy�gLj,���2���E���O`�37tjM�
L;��h�#9��WM���ִ͂���k�%�0�Y���Bj�鹛DO#�I������G�6z���e������4��su��S(n�W�"(2�y%���RweC%e�(��N��_r<�J;�]dd��GW<Ҥ���,�#�㣿�dW��7gQ�5�9���j�^HQ�0ř�6)|�;��Xpq��gr���)�z��#p�}L��S	�WE��}��8�-�b�޴�ȍ���+��Vѫ�&d��6�L[7�t3\'Q����CcYD"kfs�0�F2�4lfFD;{p��X�7Ň.��	ْ̩F��S�{z�Vs�lE�ʘ��,������{�"(�4 O�e�T ,#Y�^��gOP�U�]�)�I����J��ٍ�43Z�9i�����5u������&,����V��w���u�խJ��ŀ,����.�e�jիhh�NYT5�w�5�d�R�53[)W^���kg\*fu���-VZv�$Voz�״�2�m���k�;X���k:�Y�ֻ�ޓ��g�3WM,ӕt�M5���Zfb�ٙX����I�v�`�+��e�U�Tjюe�iKN\��Ũ���Z�;[�kR�� �t0�VM�l��f��kYb�eKS)���t�]u�jժ��Ԋj��M�{�gl�,5�VV���j�YW]INj��ԧ3WY�
�-�t[9���Q��T����e���5Vu)�E�,b�uɪAg9��kM*:��▭X֥[-X՘ԗ"��Z�r��k����f�egS@i��J*�U8L:��p��T}�5�+�Ԅ�c�z�P���wDT
���9Ӎ�&:u��Wm��W�e�� ��g=�}P��,}���G:��3.B��T�B�&�q��D}��֎9�¤Χ����e�����H��>mr¯�`!V�~?}��;�7OG�.����{^y�Y-����v��]��3r{�k������e8 �N��S*H��+~�AA�[��f�/f)�#�/WG pt]:p�K/#���kh_�����R���x�G1|���\���|����iT]�홁J^����%¹qr������&�]1��4�*ƹ��8���H��6�������1LԽ~N�
t�{a�5�i�*b��u�U��s�.�qp�H�;f�0�����݃cQ�"��S��Lg��8fԜ�wzR؉e�Sm�6�Q[��>�װ�O(�,w�XU';���v�ܫaǬ6�C�o/{&���u����ۋc��M	�ɒ#�z�c���K��>7T��my:.������^�s<HIʲU�6��=�pw��(9^�d�3YyI�x�"5��~��ޖNe�{���_���/f���F:��[׆������:���\����3�{��9z@i�ث�|����'�PKJ�5sn./�P�F�Nna�X4u�*����2:� �ɽ�;�WcA�M^�P��4�+]F'�xu(�$Vz��e!��+���lXo���}#&k�-��(oZlM�Z�{++S���݊CR%%S�3�F?Hb;��Qr�͟`2�@u�cch�R�>�EPg"c/sj�ǣ��ܽ�Iq����ة�P}rte��R��P/��q�6���裻KA��Kau���4���s�=YV�F���P�Z砉�\3�k�z}�N;~����i�3�X��j�ݴ�H�0�C�
����:��L�!����N��u�O�?����b��6;�~<қQ�{fab���n�]H��t
�\�]�x�._�8��Ftd٣��v�"���uȨ~ip�g�ɝ�V%����tg����|j�r�!g�"���>���^�՗8��$�BC�:pΫ�Nv�(T�B�gr}a�r�C��]�x�\-�����{��wT�n}l�G}-p�r���\*����[d+��e��K'XN�!��7Q�v�;�V����V�"_�aȚ���	��xˎ���\5T�si�P!�A�]/�v��-����l�\�02�D΂�a��];=�J'P��i��#��L.�Fs,�|5�ً��XTy����.{��]a�ó�p�Ƒ����Q`���+�*������M\�;��;����B��PA�Ff
����O8��9��$n<ڼ�T(n
R���K<Z.�t���Ǽ~xWw��}uʀ^���s��h��͙ݙ{��[�
�̆���
��X)����3b�T��_�8*E�
�&�j�%�Lv��Aˉ�{g�l�fZ�59�*`�r�q,뮪��a�UoE��1E/N����LV~�2U��ߥY�S(3��,"b�h�4K��mFˋvk��幇u0�j|�$�UF��[AFa�bsM>�t�>��9g<ja��o͋G^�g��bZ�3׾}�~�ee�^����+"�Fۯ(��m��˂��:���g<��Y�&�����3i�K��d\�	��*­��p9���zľ�o��>D/<I�6�).�0�9���w���h�J��즘������+��9]2�q�*��ZH��Ɋ�#Z����^zf:2�Z���+�S�6����"S��鲢)m�ؕ�.�iT�G���u�E���
��2�]�ˬ�k�f:%zB�*��>��,Jz��u��6Է[�Ճ���u��7�v��1Ԅ���K(ջW�c�U�������O#3������$�c�SNd�v�0:3�D�yr-Ɣ���N8��3q�r\6�Z.=c��Aq��a �q<s���u[\/]�y(��]��K38�ԺCɵ=���{��Py�̨���#�i�<������{��P��]r]ʺM�&�3�U�p�����Qc{�;r���.����dc]�T�Wv2c����}���o9j��!���[��$TźV��rTz�=�gEk��2���
+��f�����73�5�^i �� �A�%
����!�C���{ƴV��_������^�Z��b�c�	�~�Bv=1��3�%İ�s����*c&�-�QH�71"[�X�r�7w:����e��xR���%2��&�+�^���B�<u�Wy�ꬹxq��r=�.Ve���׊#�Qλnpr�p�8��eh�3u]�bS�R��Α���q>���z7��+��1��Ъ&u+;��Q"�Zy�)T�<������B��,�h���|:94M��n���B����]�r����
m�t��ӱnq6Tl�*���NN]���(���B�҇��'���G��+^�����}mJ�˃��KoQ>���M�ً�n���v�o],���,�ޘ�m�^n�E�t���n��ey��u,;b��4�b�G�@�>`��\5q�i��72w ���F��I���뱷x3���/F8֜9)�ڹ)y��;	O{��Dܭ��Y7ʓ]��g��[̛
<ܬo���ؾ\��kG:iNl��"=w���-�t�+���3#�h1��{�݈�`d�Z��\��./ΨvN�rG�Vļ�1���p�J���ƏxSr��T6-�5�v)ʁ�"���@�	�p�����q9��J����b�tbj�Tg̊�ϸ�N�G���aB���fs�c��T�1�L�n�s�t�E<�qu��&rn��x�Ȗ���1�=#Oi���2��X�A�g>�q�a�Q��;BZ3������A�	�h���0��[s]�J&+�z}��%���O� ��i�a\xh��,�HV��7hho�I;��y6�x��r�;.��Tt�O9����['Ո�������^-�)*O�L�B����E��|�ׯ�=]��M��>�7�b�J��c%�FaMn��ʟ;�lλ���a{\*]9�0)O{TS��N�L�W.,K'M�l��u�v�\389,�`!�Px�����5hZDU���d(�5T�}�N�
k�*�~�IVl��L���c���jk�*��| Lj��e��v����.�:��ʗ[0�ө\�cj��S�z��j.u�o������-�7-�=�.�;3F�Sy^�Q��, �#L����%�1�v_m]��e�{�v��:ċ/n>d�kb��V��n�U#r]���1_Z�o�Q�"�T�`�D�|�0�T��wmR/;���C��zi���^X��Jo�
Nv%�˃ct��rz�,=�.�'�\$�Wr�]P����ZTvh�v2d��P�Y���U*���󨗼s����/�9�HبХ,���PY&����;%��fQB����>F�8�u�nv�Qv��W)�[95��8C���_fņ�����l�gb��޴��m4s���x�z�w7���}sCH��;���*Vϋt��u�ca�[����ًu��5[�7�^`���@�)Z�є��+���eB�	��.ưE�	ۏ�N)��}6��>��Kn�I~����W�A�;c��砇Sʸ8k�z}�N;g�Ar�ɗϸ>�ϳ�^�5k�]y��vHV��L�:��L�"�i.�o�	W��B��{�̜DQvz�j��B��e��8v�3}��U7.H�#�R�J�BVH.M*�_t�u��~B�#��[��-�
wr������2���%9�fL�˒J{��a�wxg�E +`\;�r�����}�Ӣ�4��Q��$M�of�^�b���\�]dv7nJ�o�ôĉ�#-��)X<L�4�c��y���H��3�@���d�<����m���zi	Eq�g���̫\u�A�%9qWT�Jݳ��%��yh��xRI�5�YS9t��Γ�ܫt�]_���t����d�M����\F/*g��n7�uB�K���#��������뜋�������XY
��>�q�Y8!M�=��q����\���s+��2�IҢ��Ӎ���KUL6tR��4�It3Z��D_���=mW�� Ԕ��k���*�2s�h�7���\�P�K;�كɍ�y����"_�u0σg���F正0jH�@�+`DM�s�r]���o���	�O�K"3�f�B�|��1�Ӊ�l�o��%��������K<H�,U����.�5����#Zk��L�����};e nW�<�ٵ �Q�[�LSU��.2����|���ޱ�cld���Po�ׂ�1�v�,�R���x�2����9Z��3�4k>��ѩ;]���4M9>��r�ƶ
��:���E�[����ʕ,������I�.!�{v�x���K��X���t��{�.�Y��jZ#b�p�?{�(2��g��[{��[�P���ڗ*.3�����1�</bչ��ǜj"�%�e��n�����v�d�lW]xP�UwKN�q]N���e�e���9��x�l�Yף���� .��{�5����
Fĭ�����=�Tކ:U�z-
��y0��N����R��cPg�nQ��b�6yn�+�u��|�_�Ϛc�?���+t�k��xk�������u�|�"L�|��֡`��^zf:2�)��Ѕ{c� m�(G:;��1�h��B�jU�_q�_Qs�sUc�`s�^��A�]�3�.":'B� �B�n&�K)�Y��F��.��I�r,dڞ���>}�Z3�����v�a�;�eJ��
���BmjX���T�#`<^�
	�ul(޶S��Jn,��9�
)F�(�Qƺ>���؏���u+��*�qh��Ѡ(�\>c�x^��>�R�j���l-��:F��[ιQ�v_�*#B�y$E�B�*f2qX$C�*&+�)�Η-p��=Sj���m'�Q�1׺f�i�uH@dC��L�y�eW@�Q�E��D;j���Ϋ�w�S}��Eh�:�����a�fb�e��"��b�<�VÊݞ���y��בoN�K��ODse �gAp�a ��l۴-�*���kǝx�V��������l+�Djo�;��',"\���;��t��؃3�)`fʻs��]�]�R��]WN�:�ԫ���D>�zUE��m\���V�����75��W��(��λns�=C�쮵�#=��Y�+؃�t��h�ơ��:f�}�78a�"�j��Ys���}Y���,%K�8��+gq��N�)	z�JHf��v=��ߕb�7(؜�G�Y�[E$=N�����=�*ky�Bg�FYR���ٚph�Pu֪���t~\R��:�>��[=0�
{B��a]]n�ʥ�ԍ����U�Z|��kG:iM�XkIt>�F�e
�}�)�c�kҬ��''���F��[Y糢�2H<�l�edu�F�G�V ���,"8�Fϙɭ��FM_U=c4��
���sM͌��@��JzƠE�;����uC"v���J#ﺣ�1�"�<NcRĬ���(qN=R�aB���V��:�/ x㾙���r'k&6��&%rd��z��}s-��mf=SP�B�W:�C���s�G��rFYld�v}>���-_�+/���^E8���>��!+���A���Ps�>+�#<����s+f�
Ii�7+!w��>S�@��u��V<sx�T���.��Dk{C���l��&�R4�9�K/GVm!r�n�%��;b9�3(�%�1Ɲ�@a�[���ݵ?�zy_��Ϋ�P�+t�uΒ_N=, F"N�VXź���Z�����W'�l�V�n��$,��'.�_�����Q0'��b"��R��8,�]K��q9	K�R�˳q�6oD��c��b�IB�Q�ܽ7����W]l,oO$�"e���Du79�0)OQN/�;�2�\��dੱ͛�bL���<�6�;�O�����6\n���dQ��ٰ�(�j�2�31\�b<@�Dʫ�.�������K�Ѕ[t�1�`Щ�<�w����ΞVq�"�ʦ6D�]L��j�O-YϷ�ecg۪aP���	4�Ү
���o�
�Nv/�x=�1Σ��L�;�XI*Fʵ�2�������l�=����6o�sޕd��>J�_�)u���'/��^�������id]���P0ܣ:�I��6jUs:8]#E�(Mh=wKm���<!���Vq��;��1 ��B���
�+�ؿ7�lt`z�	O��>�!MV�'�a���e�)i�u�^Н�R����D�b�ڢ��3�퐜�gX���=�7o�Nq�T&d�tTKX�	���>ތ�.eHr��
x�^Yd�PV�'`�r��,^��36�Bb�:t%6kQ��H�bR�2�n�b�*�Bv�%#i����Q.�0k���fu�#�g��a�U�X/zɓnj�nP{h���W^Q�r:U�(����aC�]l�^�vr��%��-J������ẃn��:�y����
�wq����(�ԈATEui���p�Fk^
�]����s���؇R�"�]��+���%іx\�n�#�ٻ4 �����4w�jP�2����aQjak�ǗX1�����Ǜv����W��W�z��=��ŹY�jS�rn�nӝHswZz�J)/�]@�ַ���� ���C��h�}R�֠��b�d�|li��E�svo�hF�5)�oG��9��TtZ����6�=�����f�Sp�Bd�Tj� n������
��;������Z��tE����@@�桃�I��+���\�i�ug,U�=˚�|	�����VM2�&R�]���!�嬕e}�u��VHwҞ��k~��&�H�gZCdB���(�Х΁����(��-^�:��יAKO85���M��uhY�R!�nFk��j)����낳��ɵ�34*�V��8�]N]l�,AOkX��xsX+�GPgib��5���y�j�m����m�[u���e!�pq)е�)K��ĴneU�n�
|�|�<}ȶ�/��꼧Wwj�GЬ��9+�ҙ�Իt�.ۮ�Bf�$�9�=��sKr�B���=�|�VwR��f"#߰+4������ �sN5j�mcl��>O)����KId�xN������MlE"p�z�ǆ�ټ!� �f��;����S
:��i}�i���޻��wZ/��A[�N�B������lk�y�
�|����C�/W!��<o���!�5t���%Y�b皀)m<��O�Mވ!J�sxq"�Gr��mXz�}O��t��|y۽��3,���Tk��!���S!�T ؂�z�yf��,��j^$42��H��lV��S�����X�2�,��3Vs���h��3$7Wk��]1��:�fR�5�@�hT�Ƶ�\sY��>d줠��)��u�$�t�l\�?7Q�09�{���!� vy���c���f`���0M�"�ąJWt���Q��7R�z��f�f���9���}������<s��@(��J��f_8���6{�˷�[J���m<�%�����L�efv�y�2�fhg �FzY9+4.7���� ���,w�f�L��a-Dj�AY#c`�Xˡu���ƌ-��n���u�ɵ�6�+r��(�A֍��8�X�A����;)�i���YF��]]����F��z��Ϫ���fn��jZa��p��lC{@�� �oY���j�.�����%f��8��z�JZ��YSj�։%��sZ�j��r�N3��m&��E%n����kY��l�f��ZT3�²�;T�Բ�Y�W4�r��ʓVG]l�L[��cV����FZ͍�q��iؚΫ�3Mu]&V����X�Z��O"�M�2Xd�%cb�֖��V�ζ�Z֭%��3��]�k�������VU�ʷa�H�;]V5��YkV���n45�JcJˬ�r���ֵ�CjIZ�Zf����s4�;��8i�d�j&��:h�Q������Z�C)��q,t�Ֆ�ir]k9�͝5�e��*Z,׽��d�d�X�l�u�2ɜ��%f*�M���bb��YW]:����ʵ��ɔ�fkY]dT�U�W[1�t�-�ܚsl%��6��R"���I��;�G�ݦ�c����Lf����6jESq�)���:zt���H��4��**��j�3Z�E�����5b3�u��Z�N����e5��O�b:<C\48��u�!q��[����Dd�#kk���:o���p��K�������ThߎƘ�R砇Sʸ8k�{|t	�,�l��D�2�<�J.":嶠�i���vHJ$t�*�N�2�i&�ڈ�8���"�n�^�gW,�c��<|��b�+Z���]uZ�R,#�R������>�9�!>�:v�n,t�U�`wSc:�Ȩ���2Y�w�;2���j
�l���8� t)�u�VڇjʹEnne���꥜�W�^���9<�T�g�u3�>��9S~R����5�������"�o��k�9z�<v��_�����T�:�#Tu�\��C��}���Py�w��\bK>�IJu_�߲�P�FWU���j��pBT�? j�nX�F�f��Q槖��(�{��:�v�V9I�q^�V�����U\dϨ�$P2yקK�Y:�kq��"r�R�:%�:�E3�њƌ�� s��J�(L��s��@@%@���R��:
�åb�H:�
��v��H2�鮾�Ky�u��m�[�8|�C8M����َK��=��d!b~%Snx����o��y1Q-[�4+0�����I]����.��_���)�Ў��J� �ֶ�u�(G�f��&�ZuyG~��.ep �=pE{��ؙ@�0�����t�b����>ٖ�MN�̽n�{:��`��I9�K�<L��螭�w��.o��(X�
��i��5�u���Yzj1������G�K|��Qo�2z'gK����h�.B/c�!F�ӻQ��ʼ�v��uh����μf�|˵� ��]]�|�M)��e�5�U��:-ϔf*.[�E�����Us6�g�os[;����1�����}��x؛E�h��Z�����*�p�Z���+�j��|�r�>Y��_K�qb':�N*���uO�țs���X��J��7ˠK���'��f��l�t����B��>�+e�����W�U�$!^��T�Ym*Z�3�4���rW��`{.��D�0���V9�P�ҙ1�*m�9R�!Ę�̸�u-s�1�o*�	~ʈ�=7J�I��"�M������P}ζeE��'v�2�>�n�A��"Gt�O��V�j������K�T|87�Ճ�ͿN�0��gOa��h�n��r!t��١��ܙ���$��d���ʂ:WN��.y����}]�*�a��vF��Z**m���HV%�Nn6���/�\�0��Q�u��\&�s:V�)Ɍ�VD;���&Ĭ�Z�����<8*�A%VrS��/ouh�Ƈ*�\�*�lf��K�F�+ R�Ꙉ�J� Uʏt=��:+\����7�Msl�Fq��y�u1r�]~��X�r�H�PdIW@�38��nL5bC��	�4N��ԕ�cmK6Az��3�҃3�p�c��:�)Ĕ+������e�U���v�&�Kw�������w2(��5�]�(o���)�6^�Qp1^��8.,W6��jԡs���[�f��y������������C��!ǵeh�3iU�WMS�K;���~�o0W�B"�8-Z�>�k#Nb��xY�f��X���>l���R��W��IJ�0ݣ�F۱�C>�دh�rjFAVNC9��Ō(�7G��L���Tb�����zm�k�zOLӃD�������3�k�r_���n#P��b���-�����6u�Q�p/ݨ�ߙW�a>Wд4s�����'�\((�L�4��UaU�7�kw�#9��u���ר��y$u���-�\XuC�v3�=R�ϊ�6�6���d������yt��,��2���b'��RU��ۙE�J�� �RL�J�m����{�'�;�<[�aK��Ow�W�v���3��'�Nqڎ�Df�%Z[���]�U��i��qݴa6�N�zm$��vN�r�Y	[p��£�BWw��8`M��)�%�b�Ѳ� gJ���✨dR���m2$�Q�q��ә6��ٕ��q���K�ı��H�#��G�ODܸP�����:�/ x㾙�[���q�\]�$�V�z��oY���ٶ�\����ч2z�2��X�A�l�҉Ι�������;��QI*���U��0Z�sME8���>�8!+ �z(1�,݊7��}��}zdԯ�~F8R�򘞍���]�>�P9 ����ԗ��$T�ʂ*Et��/�n���R\�b:+a9�΂���^�^��Y]V}��^����W�A��Η�X!�oS����;/�a�Z���w:�Sz��_g���W.,K'M��7abS}�
pqS^?(�Һ����9��t)�q���d(�3R��w0Je���:75�6�.�滒�,f���./�Ê�Hܕ`������uPw���ܺ�ɡ�ev���ގ���O��aR��U���n��pBŏz|����K�~�>�e/�v�`ɸ]൅
����w�z���u�m�@�sW��*sсa�4u��40��3�}����ؼ�&�����a�"�u{�^_���\C���d��X3��nuΙ0sEI0�d#����ud���>�k�n�Mw΋��{����ӭаxtr��H{5�~�{U����C��"ۣ�E7c&Lp�U{c�*rWC!�P]�Vtru��\<�W^�V���s��sc�M����/�,���&��h��.��`V���[Os�z��S�x�i.��R�砋4���B���U�}�����2f��t#u��&9ۃ'���bڃ�>�u9\H�p�.���)����d' �Y�6(n`i��#3o���|��늷�~	�͇���>�F���/.�LR�cX"�у��씒ss����������0�8(��Ї�V��7㲚0��z&�AE�NT9��]�pu�����<��ARqt����r;$+SC�P�Q��: T�B)�D�f�s=%��<\���SEC��U����i�P����q�{*��qu!@��B�BF��Ś��v�ޣ$����bϯ� jlgV)
���g�ɝ�W�q�5�X�{}z��{ǫ�h���8�]`���Ea���H9h���}��xS\�4t�^yg�y(��� �%A���o��N�4�����@�sP7+���K�0]�e��&�Հv�n
�z_���E���=�KK�ﳞf�='j��[K�H���`�m�<i*�rL�aoN�j�̺���3p�Jĝ1�6��W�Iq�]��Qm�Eh�O�y`&�����c
�X��C���M*��p뜋�n�U�B��W9���cʹ�g�t�X��r�2��0�zEB��-�(Ս�U���AԿ?	�|�N9X��NV�t�Ɨkw��ٍ2Ӡ�BB���wAJ�S����]K<Z.�t�������Z\Û���y���R{i\�
�E1%��D&}��C�sV3���
���X)���y����Ǜ2��{Z]&�g"���F�[Fr�a��z�϶e��S�\T���9��1؝drV��z�♃r`L�.z,��ci� �W�<�ٵ �Q�n1N�5OtqT9��'��}~5�ا��A����u��t��1��N��wj<�f"f.�l�o!+Go���(��|�?]���>ְ>�eևS��)A��~��klzdԞ��.V�p�jzU�{u{5��@�dT��P��;8��[��,��y
^�Ko�;�9�ן_�ڌs��p#:�OU�5W���B�V%J�vSLuCŵ��S�d�f]�Rپ�Ӵ�v�e��8�Q1,� *��A�s=��+�%oޝ+�l���_7���gg�o�U���������Q��i٘��v�.�3��75kU�5H�^X��,Txt������I�����ۧZ�'&!�Yϫ3S�F#�ؠ� ����]��O��ԫ})�Scd�K�L�B|߱��Y�J�x&c�)U�U�%
��K4��r��M�]qb�dM�P4_QS�sګ��)B�����z
��v���C���Ģy��(1/=C��Q��"�ХJ$��d=�U{,�vs��Q���"a^�OQhv4��Vh��Ȩ�~�\Q�**8+��G��V6�;�*�0�����Lj��I�J�\��Y��Z=�L:檺��Z"yth
vx}>Y.
���n����M�zi0����W�}�ЭS��PH����!d��#|z���d�7Ѻ#���v��`��H�-Ou�5|�(�~�)������w=�&\]�!��=0}͛3j�I�o���
 �K��>t<�g9ٹ&�)g��>���\b�������$&P�b����+�7z�f!3rU�����b�_+^u��)�����6��P(�]�9ˍ���V��)����)�Uni��7�\Kդ+x*V����V9xdi�b��~�ϫ2��ՎXp�F=�{n2c%���j�_��^�H�teЙ뢷�] C����ާ�v޴���Q�����F�4�ͨpQV�"
C���cj���}qeel�=�Q��șݾ�S�Qfd{}����7�Dlu��(�[��R�Q�X��`8{]2Z�c�Mgﾪ��	%�������V������]Ҭ�|�9�ѣbu o��G�_|D�HS.�y]־D����I�L6v/��]	�w�#���s�2|���>�5YN-`'�J��A�<�6 �(N�%�+a�5��s��G��W�a>WК�ٮ���(���{8(��Ľ�λ��S\�^��`FD�<g�wX$U���-�\XuC�v3�=R��Q.[���Ua��VG(z��'�U>���=�Q�]+$�P/dR���n�v+d��<LVvRjT��z2�o�z����@d���Rѡ��U�������%�g��9y�@��d��W���
W&�/e/z
���{�$�(*��#��h�5AG��*/��j}���.�;g��Gw1s�t����d{v�ؘ!*W4�S��~�O�����t5��1�^���{TȤ>�W;�w��P �ܡ�j�GG97�g��>�:��e( �N��9Ί��Qw��e��|79�U�Pږ+���B��s����(��cG�/\��^�G����0HQ�:���u���f��Cd�h{p]t���ښ.ɬ����6���M]�]��M�\wH�w2�n�-?V�k��pG뙫vå}#é�u�֧n�
z�p:�cEgp]cG5Пt��.	����l����e�U���Js�xa�x�Jָ��٘�]5�r}_z2�������ɟT8�.��S�%vBc"%�'�N�)]��L�ce��!灨sB��W�cװ�(Z�L������OS4k�Q���jQZ#�6�J���< �
��#Yg�P[���� ��Pw��_�AQ�������քl�!�ȗ%����^�_�G�hk��oiW,X��X_I���mbH��ДWv�I�rK#/��obo�l8���A�&���sJ~�N}Ch|�]+�h�C��H��4K|��%˵,
*�x��_No����n�����_PY&ޜY�:��t2���3����2{ɲ�s%H�
�2DoOAi�����R�t'}9�}^��٪��Y����Pe�K�>|Z��cU�oYl=�Z��m�"\!	M�Qr��v	�iXh���rx��d���0 �~��]u�B6%m5��'�b:<C\41e�&b����M������·}֔F�n�x�9ӊqUt	��v����W�H7㨡�.zu<���ڵu����/�wW"'�4t̮�d�ڽ+	GGx>�=C\��{}	�-㕙A�<'�ZM�B[Y�=:��Ӊff�9ώ�v�U�1ˍ����n6����c9p�K��<�k�\9�f�6�r�s1�w2�Q�ek��X)��]�S� |���7��*X��ӿ�V������GXm�@�#�BQ#�w�u(� X�Ge��h�[~��x�\%�Ԫ%	k��b�J��X	�P�����3�Ua�qu"�R:/HXUB.�7��[|=4�Z��Uk߯D
gQ�~4��Z<ߟټ����]|�cг;ϲ7����4V!	=ib=��UQ���4zH�Ȱ��_I�n]�P.����uo�9�6�5�/^	Z�OI!J#�>*}�/�@W
���hiU-p�yo�L�
�;�[B���F��3y�s;�r��.���B��	Ϥ%B�C+�UcEW�.9���e�݅�Dv�s�[��rTb'�4�`��� �@�p��7���è�
�J�}��ՙ�=��׺����x;��9�4DS[��S>�a���b�xs��J��}������hs���F�]V���@��Jb�kVm�P>JI��3=�-r}��XR{��s�!�a^�O�b��[
d��ޓ/)e&�޼�(�d���Z�e]A���'��F��~W�Z������x7Q���ZC!����m&��f�RZi���ή��$�b�0����S��re-�T����H)�S';a��6��4Nݹ��O�P�����j��^0ʂ�T4׌._��w�J����1�F�WM��#7׬�y&fK��.FfUm�E�خ�&�(鑾�^.�:�,phh�u|U��5��ͧ{]a�{���ur]���٪�{͒Q�C�r�H9�hKMw6Y�C\���_q`X91V�Y��d�ch!�&n��]VG:'�G�����c�v��`��;V=�-��`����I��e��u�e�bcX�p�]ewYh���**�JR.��]���7�����+OM�������+zc���t�H���#WPp�R�2z�uiGDeP�9�����N�)m[�+ ��J
ul��X�l>S�`d=3Gm���ٰJ�	�����*"=ݹ�Qwں��=z���r�@���6�V&vV��i��w��[t�O@�SV����:�yes��Cv�MџlN)��9�/H���L��u�;xqw���Zk���;ڮ��v�G	p�;�ھV��lK�u��b��Ι5K��㣘a�o"���ЭhE�,뽌j���p㖴#�b��.��PݍQ��L��\��z��V�6dU��:����+9լ��"��w
��.i�E��׷6�9m� 2��<��.���@�W�����^�ʕ3�^h����9b�+SW����2r%:���ٛF�>YܐU��n��;ޱ��u�i��^��w=7Ԟe�%���[˘��R�{����"�Kj*�)"c���W����\׷]���6kt��n�q��w3d��[��[�����zf�h�wL�koh�=3�oZ�Cup�{��H:�E��Uh�Hұ���;��Jap-�e��߲�'�w�kWQ����5�P��ڝ쫚�ó*Zp�o0bT�չ��֥l��|�
�vL���۠�6S�TC4E�A���
��+ז�;��la9 ����q�;7���f�2��1k{n{v<{C��t�\����l�"�1i�-t�Z��ui��hO���J�vVm�88�H���-���\�	���<��)�)}+�g!� L'��knMSK�P.�n�()�j�[&�,�YY�u��TN��ֶ �lԩ��W�J˩��
�5��W|&l����	B�|轀�\�x �ӺT�P�3s�cY��K�th^��P̵��2���o�maF�;�V�:�7��h�c��ѓ��B�/$Y؃o+E��8�뵶�P��`YC0���N�$ҭ�'��E�;�W0���Wa�v"FoJ�u����s�^0h-�(h%%�r>��0���]��u�,v!/޴F�C�Z阯���ibq�pڙ{��Y�ݵ�Ug<6�J��@U�)���kp�L��ְ����^k�P��y�f���:K9�\۠���`�R(�۠�1��hq��/:�Z������{]��=*�!/"�Z�_�^d۫�U��Ї2u��`���Q��w��wnVjR�Y�������w��Q\]J�\u�fN�h4�(��)����(Ҵ�mvJ�KB��:��.��V����MuQU]R����DX�)ڌ��o�<�S,�v�2658d �.Nt�aVe�A��Ѫu�Z͢њ�ua�*&�L�������c���W$Z��`�ө[,�Z�eV��HʣV]sK��-lhUF�Z�+U��)q��:�ԭ*��V�v��WA�Z���geb-V��UbK�e�E,�����e�͍�����b�7��%������S0�lTØ͙�8�(�Փ��#i4�6�Ӎvl�����j�[3:��ΫM��[]��f��,�Ē�2n���N)��J[0ĘpO{Gc��q�Θju����ך���3f�z�oc�]p��,��U�q�h6���%q��!yӽ�L&��)5RȮ�8�u\َlf��k"�:��Õf;6+�e�6��c���f��a�]\E-c36u�d��I�N��y��Hq&vg&�1����Tw��©jy�?9�������Y��E�Q<l���Tnv�H��p����*��w?BB Vs�s��1���o������L?��d��S�p�@��C&�e2m��
L�T�;d�h��P�m���d׳�H)�f�Y:����O��=��U
gY_QĴ��3ɯ�V=tv��O����9����}�}^0̰�R�޼�l4�!�-��#���Z,Ù߬2���-�{Xi4�h
)�))����(�3̚�\���aL�������2Rfk�L*���g���)�Zfe}y�)f�v�2�<��G���Ϩ�0�<�����y0�Y�c�C��6�"�ޠ���ha6��͊A�IL\LЦXa�39B��=�-&LQh��
Oz��k)8�0��G�>K+���M�[_{�xtxLӔL<d�Y�57w0����ɣ~��RO�����p�3�!L4b���Zn�gm��JG���'-�d��RA��L0��@
0u�|b�&��>�o�J�� t	����%"�S����0���M�y��Ob��>]�IIU��@QO33�Xq�u�u��ne:ɶ�D*��S�Lv�3��Ɇq��A�}�g?W+��˾�g�<ߵ�g��
AN$�D�VRA�{٨uP�g�y2�YlɯXe�aH�35��e�ai�2������0�S����u)���̽Kd���hq%9z�p3���>�����o$��: ��G�kw]�)��S-�Q�d�qe$�T�B��2)-�m���c�B�[3�Y�g����L:���Y��nL&�m���?�I�=0.�Z=ҪV�{�;v�|��p*<* �)��\8�Y�*KC]݆a���C�S	<�0�7��P�q�aI�Q�l��:�1P���L�):�I2�J�1&�]���0���O%��[��7uv�<{W�ou�9�,�N6�IX햐S��m��Xa�
H=��߬4�a�*���Ʉ�3*ù� (��҅%�a�-�uSL��C����@������d���-�֙�'>��Fm��_*���L S�T��̝o���2��)�'ޣ�Y�d�)��sT)8���a�'��@�~��]C*�:3�L�[��(a�aH��]�c�`�^sǵ�T�����mKc:��:YڎKJ�/:m.�f�1uG�m�ۻ�HR;j3˰7s��Vp���:��;���-!�{ܳk�����h�*>qL��X�vʒ��,�F�^V���|��9���_cJZ�S�d��)W*k�u�t�wn�g� c;�s���y��|�j��������iH`3�&'�-�UˤP�Jr�[�KB��M_,���2��)�Mc:�Q�a�W��m%*��+3�����2�;�)���S�-��qjH���,��%��c�c��x�̰�-!H����2��=��e �αqfS�-۬$��v���v�H��
On��zᤖ�0�d�g�,�m��}*�	N�)}��j��.s���x���òiE�=�.Re:�I4��*M��D)Ɋ��h�O%��Ԗϒm��>��"�R�0gז�) ��I��z�ho�L e)�VWjR�u��/���ngǷ �i)�@P"�.<-Osv5Sl��C]��HJd��ܬT�J@S.�d���3&*|��O7��ja�
vɓﻃI�d�Gٹ=���~������I��g=h����d�#������}ﾼ��:��]W,�:��
En�i�|��e����A��hd�mE�6����In�̖�&*Z(|���a���O��y����0�n��]��������sK#��G�D�=��e<��Ru59�2�@��g�~�<�=���v��&�m�KI��3L6���>��SL-��E2���>.�ŘN��Lb�L$�ǱϽM!��=�3m��^�J��@�aI�o�)8�0��'[a�o�a)O�)�s��@Qz��nM&�)'}���+�}�2���&�o���,�Kmf�-���>�~͚��|!T鯩_T'����F0]�LO(%��*�I��%3���d��&Դ�))�!�����'qGǽs�2��Sb��T�% s��8��i�
��pN��
=����C%�3��_C�\��}�k0��{t;�)�a�a�M�
Aqu��VR�#�!�u���a�aԶ��ٖygXR)�݀���f�JH9�y9�\�,��0 p>��w�_̾�ڜ����}�,s����>d�{��a>IM�f�높u
e�ɪr�S0�8�a�qDs3&�)U&���ْ�tì+�B��gSL<̥���Y0Ϙy-2�'��^�yy�g�mHقcGrS��z���"ŵv'[ҕ~ �K���k}~�mn�1Ulh7�wɊrP�o��wU�Mk���ݗm�A|���v2���n
�6�p��{����9Ǩ�s��CYג{��Y�3�?{� �O$�֣_�H)�'yYCihZA��CY��a��\�e'�S1��L$�gqer���B��P���Y:�b�hJ|�wBβRAvg�'�)� Ly��Se���:�63qq}������N2�D��0�L;tN�_wפ��$�n���hRAN&~�Î�-�L��}s�4��>��v�(J@��ϩT��X_j�"���멚�H9��K$��mW�ϻ��>��{���	�UI�q	�[�u�l���M�uÜ��6�l���o�u��C�d0��$��0�ԅ��Ҭ�a� �d?�jX�[��ӝ�_�=1�*=�'��
a�ai�nèe ꡩ]�au� f}��!���<�N{0�RS��=rRN!L�/�gVB�q����4�h�W�<�i�JT;��+x���:>իS d 	���uz0�
�@Ɋ�
f��q�KMf��S����- �j���<�B�r��,�u��7�%&y
f�G���I�Y�~����-'��������ε�v��{��>�6�Z�d�l�Y�@�S�/6R,�% `��&�Ө��C(}���Wh0��S]a�Y��Afd��)4�$�mI��R7�&.��[r��/w��y���Ù����ǧP-)I�gj��2W.JL���C�jH9���厪aHJV�Y)���-6��i�4��M!I�&O�y��aN�Rg�e �+�3�c<�1^�Z�n�����9�g>'2u-����%�P���;��A�!ۣ'}s��Y�Ka��\0�3h[0����AL2�bo��hZ�sS'(Xau�0�U>JC��<�Y�)�S���u~�*r�cG��V�� � ���U{�}��.���L:��v��2Ry�����C)�
C>ݚg0�
�I��s,4�%��2���I�0���W,RRAL3�Yh|�B�>���}~�t���s�������ILY����PJI�)�ֽ�2�Xd�.N����O��ņXWhY:۩��m�P4��>��Y�JI�P[�M%�Y7��R|���+4j{�X|�������[[D����'n�l�N�-Y�*�L9>�B�x�5O��v4V����u��y�V�7z8�2]9�
�W\�ܫ����#V̧�E]�U���V�ž)�Xf�Z��,P��Ω��������-��(\�>��n�Fot����1��<��לǅ-2�Y�?7B�&R�H`.��'�`�B�X�/�)lz�hJ@�(�uRR�>�0AN�������B�ju��9�Cl)^�0e!���Jo�Z�1b��kh����$�� \{� �������C=����Cm�ɏQ���+l�r��B�R|�BN�5w0�wD2���B��KM�l�<����z�QH)�y�_�|/�+%c��}�}�W����ׅ6������a�E�aL�jL!���8���@QB���0ӔI��,�Ǭ�!��fXu�jb���JO$�UJN�I�
M���<�XWh;���a���rV�ܭr�c�p*<>O�����0�{ٰ��ANz��8�C���㸸c�%1e����HJI�)ΨyRaE�.���ޠ-'53a�a]�dɎ�Xq� ZS�w�s�i=�g�o�������:�Hx����i����(v�N%v���0�]�ғ	�O{�t��Y5븧>m��N�0A�il��*@�S�TRٵI0 �:f/�iS`7y�wWʻ�1P<"E%>9��P�A������T:j}�>L�9U0�Y��E<���w֠a'P��h/��tB�q3>�̼d�a��z��2S�L]
k�`)�(�������+�ly��o�n�� |�|8�4��T)�a���l�̳�[/�E �3�a6�P�O�f>�y���0��8�C�)�g���4���=��]��i:�_���M^,���_MCϯ`���G��v��}�W�(��8�(����a�d���*�8�'P11�%3��u�v�f����l3�\�e �L5]�q
E!�����e�����z��jJb�&g�@@�p3��M�TW�{���{�%guRZ���0�	�P��]�B�e�b��W)���s;Xi��gY)1
�(�2y-:�3D�JC�Rk��!L2�⽌�䴂���L(��#���tK�4G�����=M�q���Ϭ�A���;�sꆐ<�ϋ��)�|�)'}E��R�C}ŋL<���v����8��S	���t
�y���u�a
M�ƷX�5��������,ג��"<����x0ֹ����w���ef"oƃ���E"A���Ofi_nj�;.�;R4n5�،l�m!���#C=�:��î-�ۀ��V�Sr\ƞ	S:���1�U�)�Uy�Q;��v6(L-ӽ듵BVq芉��+�� < ����o{��$˞�
C�v�S�L�2k}��[%9d�ѣ��)�
%�ê̤T5+���L�sřH,�0���)���R��а�m!i3��C��:������#u�v��3����w�s��R��J}[�̖����ɇ/�-&]}˙gY>�\�,)�2�y�����[%'Y��\ʪO���J��$�4�0���B�e�KfNz�e&2����U��.�ʭc�U�d���ע�CHR(���,�:�B�L����,�kVu�P>JI��aLϪK@\Ͼ�0�
Oz���v��2�L+�)��.i���L��2�fRh��(
.�--5�8�\�؍U�}x�x�\�> 8P�����f.�S�aʎ(�O%�2b�m&�I��Y�%��:�����$��͙a�T-iO�[�2�ΪJfM�p�):�d�l2��з���'��R�϶=�3�q�1����e!uS�D��S��y�|�7�)�w됤Ɋ�a�l��a񚅳l��&��
AO�35���e$�d��ڨuP�u��}3úǽ��<ߎ��f��'�T�(�@w"��<R)�=ygXi>ChZ�#���-a��2���-�{Xi4�h
)��R[�����[<ɛ�ɹ��a�̰�h��8�I�m���񪷗�~�;�ϼ��>�9��ʪM�I�k�$�:�3����g��sp�<�H,ϱ�!��B�I�PZe�̴0�NOf� �.3B�a�����
��������a���O|�b����̍�^�� ��1�9G*�ۆaH{��2R,���������~��RO�����p�3�!L���Q4�K@�wa�I��a){�!��%����) ��f��cG׿���]˸�"ǅ��T 8�f����yRS�T��AN�j�oqd�+:��T8��)I�7�Y0���gޠ��$��f�S��o�C�v�8�1�0��پ}u��[ݑ��˒��\{� |ϠФ�L]��e$�1P9���
ff;p�e �ٯPa�aH�7�^,�N!�-��n>�y����a��!�k~���l������7�9�W�wNVB!���vp�9�8J�:^f��#c�hJ*t�9��̋�`P�m�E]kC�}����8�j�)�m	ֿ�b����1��GzQT�o���za�1tRްEgu�|8V�O�E6d�a�ʮv�z]VE[�W>
���'c23�H�?����΅M��>�IN_�-?���f�1}�}wp�aL�0v�qDu�qe$�T�B��2)-�m���}��ٹ�Y�g�����0�ZB�f���02<:=P�/��ywm�k��p��3���9�σI%'���6���<����8�Y�*KCGwa�Xe�&;P����O!L-��U'a��Q�l��:�T0����):�I2�k�ěev�S/�����]h�:����}������k�'ii<j�q'�I��g�0�Sl�m�-��{A�~��i�بZMwvy2���eXjwW����B�ݰ��LQ.�i�بu5��@������c�u�'��^�Y�?n����vu��S�v��i�
a��t�l�o����a����Q�ꬂβS�ɏ\9���Cޠ��J�@�~��]C*�8�&-�([6I{׳�[�V1�f���0����_o�R��L��<f��j������aH��3��̖ɢ�t�IN^�h�u�Z�2j�g�}`e��S4�1��F���0}E��R�KB��<���f[g�~�9q.�S�d�T~}]��j�Lx5#�c£�t)�g��3�-�a��6�"�Ҙ|�C<��e �ɬ\Y��@Ó��Ry
gݩ-�)�T���IhS�g}s=�d�o����v܈C�N��}T�.H| ��H���raE�1�ܤ�u�i:�ԛez�S�Pe�3D�y-�f��|�m����a��ɉ�^X/P�����.M&�{�C㝰�eIO���t�ŵ7Q�������ǫ�Y�� 
,Nz�E%:a�-59���Lb����))L�7땊��H
c�e2|�u�l�O�<ߪ�C>aN�3�����ͲS�*Ob� �"�|��(^N,��ڄ�%w��D(����=�}D=u+>���aԴ��fY�0ϘR(h��L�l-0�_v�R���j,������R[��%��R(|��=a�je'�S>�z_ӟ��ԍ��[�il]|<&<:<%�7���Y�h��2�IJ�<�'7fSh�L�o}A���=��:�a�6����
f�m-!N}�� ��[-3;B�C	���X�xT{˾0�#a�a5�2�2灣B+�"hּ�!G�ך�Q�M�T5d���gݧv��jOQ��@�-G�/de��U�o�p]|g��xZ\"R9d�S��k����t���U�*�U�{J5Ֆ-�1J��gL=7�L�M�5�VWD�C����oA�S\��I��B��T��̀��)1�{ e'�b�}�d�l6��� e)�%#���&P_&�f���m�j�0�I�Wh��a�]	Է5/����|�Qv���������x7���9�
Z)2���./��!T��[v�i��'Jg]]�
,�e'QIOq�y�58��Q��s�2��S�ù��J@�>$����ب 	���r����	���_�|�9ϼKCi�L7����ɖaM�ɪє��0���7t)Ժ�N�)����:�Wa�u�R����g��u�"���
a�ai�h�mC)U&{���3��y��5}^U��>������>�E�aHOOg8����%���\0�$�ݳG;p�N�L�P�B�q�9��� ��1ra<��RWh-8�I-��a]���Y��3�hs�������tw���r��q�aԴ6�Ũ���~��%�i�h��b�'�[{<�I��z���̠(���+���Ϧ(X_�,�m�5��2���&1bβR�~w�~޼�YϜw��o|���O���n���jO2�DϨ0�L=tN&^N���Y�m�T6��AN'>�Î�-�L���=@i-�}A���P<��iI��U%�(��
O�IOXu���v���϶}�;�n���m �+x�q� e)�.��*u��}ʖ�u���r_l��B���o5�z�e�S�k��]:>�B�AyN ?���QfV����]ۘՋ�ΗS.&��c"���(#:+a��s���\t9vn56oD������W6���t�y��VD蝇�!��2�T��t-{�}z���}Y�xFj{��w�
�6�I9�����.�)H���p8X�
_qx:����hx��t�Lp|��y�E�ݛ�C�).ܖe���jj�S0^�'WL7@J[�3�2�S���"��Nms���"͟ll����y1�j��Z���3��*����Iͽ9����;����Q`⧝Xp�̽�v.�@����=䒤��i�M�ܳ�᧕Z{�Q��% ˷�-�T��;�-��D����j..6UHܕRc0g׷����Z����ސ�B����E���*Jh2ܜ����k��𠢄dd6�.�m�Q�T�ݮ�iq�C��^u��cۦ؞S���f���ױxf�h��ɓ#�k`���ሹRMB��3=��]մm��s
����@�
o�M��#����M�9�Pm#]�F^���睴���~�t8���(ʜ2D7=Y� gHBmt����hnw�=�.Ӥ| �~���f�����Pc�*uK�Hخu
�u��W&u-������'�����q�(�خ�[��AU�ca�[�ϯ�@�8�^b}F#���\4`�ٺ�</Gsy�p�w�t���3�j[��ǘ�3��rZ(��NJ��<w~i��Xt�s�u�\	�ľ�x�*��~�("�5*�j��zTD$}sl�Gd�N*��ի�s/'���+^��쬂@B�D�[V��EqGϥ1*��$k��=��W��"4yb�sdv�sr2�Ȁ&�����{w7켹�G�k��D����J��PWM��
�xk�'5�D���Q"��T��;�ȶ�8F�������>���� ��.lB�����U9N�*��VwjN_n�(�j}b�)q���E���z��cg�\�ទՂ�G;� �4��G�����"�����[�q�gfVP�e�w��2m��W�݂2��q�Fo����!g�O�z]/yԃ��w�a��}<�T[�+i.P�٫�'��wEg�9�S��~���]�_�r�!���hiU-p��[�K6V�LD�Ͱ������@c���T�#<)�[���pBs�r%��k#�HP����wk9���v�W��TT>H����.�j���9
	h��W�jHN+�HV��ղo�_�ۨb����vF�Up�wO����S�hB"���L">�a���R�G$u=1������(�ۥ�Z��3{#��7[֎E�pT�3(�s�h�	Ӊ�l�S��[����i�T����e��*�^�D=��H�,V#<]C®%�CBܯ!3�� ���OFk�����V�� �Q�p�Q�G�^�_F��.b��'��⮡W�
c���r��9g$n��&%�[�Q�W�:���`9\�?*�+��k�����>������5������x�Ui�k6�JӜY�H�M�7{�;��H�C�j��E�֖�أ��h���/uj�U�m�n}��=��ǅr��k����2�
�Ľ#���+���j��L���e�`[��0��2"�no^�+�ީ&U����9�Bud�#*&Tr���  �{���z�����EKC���9:�u�n�f� g��5�xIS������]��̕��z/(
��^OYQnPv���άS�UwM@��s+��C��1ֻI�;<�q��)�Ѧ:�G�`���_yu�Ph�gR�������sه�T�`߶G~�FHo.�i��q'�{k��6�"�I'�ʀo���85V99�P�W';��-!ݝ��gL�����v�������
� >ᮍ/�p.k��K3���c����Q��ӧ��ە�f!������fH�c�7�R��|@�P}Bv>��P�
S�v�XeњA���\�w ���JX�	M�9���d����-f��V@��:�b-��"T£�𻰵=h�舼�~�s�FtV�x�p��܅��_��#��H�ḌN���N����u�+�!���i_C��Ssq�:
�W0�{e��Rs��P��r:�e��˴���R����uԷ�
�DYO�t���]��6
��w0w��4����nD����;v��?8(IE줂�32�ut]Ѻ�7��h���N�ܷ�l�x/J -�ҸXA��o9��߭��|�G�,�1B�v�VW�ʺ��Qgw���=`<!Èk7fx*���	\��k��=>�`%KeL���u�cළ�:��6�d�7�hy.�;{7�[�巗Zp1Y6�|rnL�VP<�}|�<�1B�n=+��c�S�:�*��U��s^f��7:�M��TY\7�M�R�3s�"��oC�s�_=��A�7gh˰�p��Bka{&�I�f�e0��*q<J�@�3eA۸�yr�Eh5 �i��S�[�Zc.�ʾb=:j�v&�Q�wW΀��1K�k�x�Z»�WnfẲ�`�O6`�ٖ]����LXm�O�[a$����j<���^���iF�#z�R]wA�Vb�P-R��X΄��n��f�.l�%�x��Y.��gp��j�2b`�xz�����A�q��uZ�[q�{B�<�H.F��4�B���v����_K��GB�D�y�;U��Or�\�n,�z�!��h�A��	ѣؕaÝ3;���U��� ��|�v�m��G����+�n��)�G5'e0և{�f������s��,c�\����J��V��:����+]s	'[��-�%f��"�5�w[�o���@wD��,od:WL�p�y�}©�!��8�N��s3Nj�dpT��c�n��'گ�e�-�o2A�%;�^f͉X�8Y-� ŕq.C]�`�����Wʦ���]un ���-�N�;��k��I	1L5%���A-�7U�
�r���V��v�ϝ�/#aE�
B��ժ�#1U��v����c�Y	��e���*�^U��@^~�Fn��!�F��G�9N�5ݝ1�t�U떞kP�M�>�f�Ԍ�cQ��niJ �M&�{k����o�u\l�ӱ0�v�t\�H��l&�q,��dTK+��C`�W{F�P=\L�.��}�0隵��;/�8�h�K=�ڤ.�f�Jj�޵F����挫�f/MZ�r6�G�B ��&�Y:����b���F��ۦ�q*�����2n��k˹-
ERwF�U�����Ԋ����ưwǈL�m�t8���R�Lx$������g^�:��5/���W�(���m6��At��5+�`�Ԛ5�[�]e��&b�Wl{��rξ �CVD8�c�̫��۠&bzj!��iU��:���b����l��NޫKuX���\9� Jx��#w����=v����0<9V:$p:V��gc��
P�Ћ���L�1(�R��SX���U۰��j=�v��$��xs��tܓ,I��T/�n�`�hS\���9QB�7K���txR��j���N�-f�[�U�W�uB{�
��Xw��AK�r3��	unu�Y�:v�P *P��j��l��I�٭i��Y�c5\T��f�s��Qs�\[VZK���K6��*�Y���2�b`f	a��;�&�[9.�&Z��a������H��.�Y�p���3Ӵ�*�Մ�kf&�8a�4f�ƥ���c�dZ�t�c+(�\�X�`��Z41:��]wK�Шұ���c�f��3��˓2i�	�l1ٝ��
�p�U��Mvq��MZ�;ڨ�*fl�����rF����h�j�6�i�����ncK*�ui�YY7eh�N�iŰ̓3�hi�ʳ�4�fWiن�2�n�Uu[3�뙌¶��M89�յٍ�;Tf�l�4ū��Y]�fմ����&��D�0գ6%��1���*IY�i9�]���39������>~W^��+­�E��<扬�����s�鋢�Gb�rFf�*F��t��m`X5`���:��wG&�n��|<��kUŭz�^�6 L���?	:����Baʻ_���ײy�٭}qHD[|s�,���I]!G�Ŕ#=��Y�)VpDV�g��+W��m
��ԯw~Z����[{��-~x�Y�O4� �R�t�B�*��������g��0e��F�>�>���n'��ԯT��FŁ��7v�y!�v-�&ʋj��N�轚��̐�����F�˼�������uԢ��<�E�4�r7�ڏ���{�+�Z9�Jq���S��0�稡�6#���P2����a^Mz�e*m��A�\gv�莭b"�3�%�Ҹ�L�0;�ꕏ��6}U>�9A"�W��Ir�l	S��ćYmlď7�j��("��Dt'�J�s�uC"v�Z� X��VR�ix|��-xp��WPܿ'X-�{���Țܗ���-Hݎ�du�E��霊x��*���'��5ഩ�y����=CԪǘ����}jg>�p?�7*6=�􉄝;��).&~�<�7z8��5���b���M�G(�K`�,S*���f�Ҙ�K�l�o{tV��HM��R�S}�T�0�+VI�S�Yb��L��闵�9ޢ�t�T͐*wp[�w)U�7�:�V���3WDh�W<�c�d�kHt�1I1L���P��V�<@��� <�q������Y��Aq���FΠ�jĨ��&힎O��C��VT�ڱIv�^y��._%�V�QC$�?Y��F�ii7ʝ������o�p���C"�^G�f�{S4��I��m$�^ؐ�s���S�(V�"�6[��SB��Le79�0)OQN/���a!�af9��\����*2�b��S�у�I��\��t��S|�LL})�L9HE\U��N��T�%F'���I����`�LG�C�"hk/����
*�nJ�W��z)�f�G�V���9[�lj6�X�S�����L����(��k����(�q���:V��irJd����ųJ{t�~�[=a�j�9���a�26dF9j���u$���=��_I��l

.�{.���@�
o�M��&GC�
����	<����.���Fjh��#s�(����h�,{�DG�Uު�>Ţ�^�P�w9A�RN8CR,��{�5紉N�����^ �S�b~4E��Uc.������w�I�N�Jf��8�{����K�_-J�Ӱ�U+t�^��A}y��U��Y���)���@k�ça�K�qV����Hj]�=pݡ�R�`s��.ԧV���L��� ���à�&�����|i�^���Ζ0�L#��V�]MdݶowZ���< ��w98g���:�z��2�Z�����z_�|�l=���o�v�`Q4ʧh�g����Z��)�ٿ!�B�3�ްE�	ۏ8ΛS�U]z�v���^�"q�[�����%��ͤ�ؠ�2�bԅ된�5j{%DArF>�:�w�����TNf��go��&�Tƥ��^b�؁4Ai$_;Qx������JbT%�jf8�쪧�v"�(]+2ت[��Y���ѵ!���P^��!X!*�NpR�A��7�nEB�\]��|��.[�a��:�_7�|��82:�������ƫG$����k��W5���{ٹ�ٚU'@��:x|��(��Ln��ܟX�d�J���h���ȍ2Z��Onj��*�k���OZ���F�^��!S����.!UX����+�P�"i=R2;�:��P�'+$��K��zn*-:q�1]j��s�N��@�����|����R����tL���s���׉h[gȻ5��Jo��
��_���P�$7S�}���~�n34-��}�u�I��p�l.��gMi��
���va���Z���}/�"
�޾<�;B�J0��\�v��{���k#+[���ve��E \+����8�y��=�M���]�Då,BS|�>϶fU�*=�I�p��sf؛����s�諭��^%.���fb�~�tEF��隹Np9��ȿC��fMCs�r�p�ΜLV��
w ��ߺh��Av�JUt���;�Ds����/�s>Fx�T>�[���2�`,����0��1v7����Xa"�T
��|��PK�b|œ��8�Z��H���=p�'�6�Ы�_rbU���`����u[��7ƬQU��.�~WEi6y��7+�"GL�]�}�&�az`�b�},����.-�)�.��`cu{5��E'MX��Oi��b��vr����Wx|�(}~'`¼G�*\�5��k�� v��|o��(R��L�br�}�y~���Iw,�����+��ц ����qI�/t��豨W���*�Xxٌ[���(uM��"��ٜs0�)U�U�(O� �`����I&�P�����r8���cZP^�ܖim��fW���8ߗ�#�$h+�Uʹ�|e.\	��nG@�r.��޵}�s.zl�<��h�6N�U�]�;0�x��4��X�����դz\�]�;e�n����p��X���d=����wr��TM���v{�R̹�|��}9W�.�p��E뺐�`�=�{u�j��O�#7��,C'Ν}���6]��8���g�Ӧ?�O1�0>qP��ޝb�l����WE�q9�	Y�"��<<<<w3g�M%Q�ut(޶S�.BSqe��)��]��*l��j��:���G<�ܛ:�X��F�D	iG������rӧ�����6FY.����Y�xg�Q�Ǽ�m	cd ��T<r*�k�0h���g7�\]�!�.b��.��mw-��L?o#d΁p.������7O�t���_׍�)
���UpSFbp�%��]|��|��灤 ��K���I]K�O^9���2�4!@�;S�3C����b����ml���3���'D6�^�X@b���Z��~>����{���c�>��4�Zt��1���*�����.�㊬�a��-s�g����xu5��g�����S�}T�*�.6,a@������NŹM�Bj��H�95������U��xR��I��ZNR"p'ՓB��Z�� �z/ ����p/�;e^ń�_B�����!�f*�����bD��\�k%�3@����A�@ʖ��Q�y5�P��� ��l�y)��У�j��QW��I���X*ݸ!k-l����ޝ��Mɯ�7BT�Dw	����^���)�V�.a��9o��ܬhv�[i�c]�f�9�28ݨs���1ML�tB��nr+
r�b�
YZsd\���s�;�����RI�0����ޏ�Pܝ��j;�{_+�n$0����Vx���g�%ʁo���o�u��u՞�����8�0E�d8I����q9�r�|,W��m�����TV'er��-I}p��r5
㥩�α��@#����<3�O<��)Tt�4'��^���Lݛ��:7%]��KAG���?}���}(���s`)��c�	�<�^Yk����T�^~no��^դ��ʋ�;
3�>��*:9ɿ[.��=^�h�n�U�c<������w[Cռ���h�<��|��ICʸ?�����AEԸ�lve���R���r\�kԘ�Y]Vf�A{/J�q�C�c#���ug�9z���h�9�fԘ�����L���;�"T+����y0���\��m�T�c'=�����zU�i�d:���[Ѫf��y;�$&X�P��`�E��
+¤nJ�X��v\K��Iu�K�ౚ\Tv��mȰ9T�`��%IM�l7W�P��9��dJ��q����q���o*8��"�X�\�r�X0o��$wM��d�ԕ kO�fU�.hs:�ᾮ:�
?�Gb)ev�R�	�r��X�W�-�Qv��vp�[�x�.ȋ}�L�,�m�qS�F� L�"]ǥ	]�;�F��2T��#W0h��V&~ {�����X�i��0\}�1p���E�r/ج�7�m	�U����5�o�b�6o�����%�NvdO�U�f\h�V��9�T��P�Q^�G�ꛝ͠a7��7:���r���5*��W))@�/��6j�ݒ���e&(	�\�׼plk�S�ABЕǎ��d.�wms�:ߝ���j�7�j�%z��J�*�X��X����Qf;�����[ܶ`�ޗ�E�s�SL���:��6�E,��@�� p4���(M6w��&"�Oѯ^�a�#���҅�L�)w�n�v���t�
��OZv������035���y�Rk����`ц�=�(ې��٫S�*"�};�w�-�쐌��'u�ώY˫~	�fc�9&����W���C^I'���b����Ҙ�r}�������v���c��<$�p�}��u"Ԏ�AzB��`���9�J��T�M��=�ml��{#5T��4���H����;2�J���!b6D�t�V��HY�Қz]R��IC�������ۜ�n��!���噶c&�����=͑����nY����T�ـ�\O��
���s2�gh�B�+8�;�C[x�umu�{�1��Q��z�LoU�h����\]�q��)rl�N�a�ч5�,@����C}]�jy7u�17t�l2�����[13u����������iޤmnJ���(V]�+�w'��v����§�>���}~<�{6鞪=sͬ+���׮l�\���\5W9!\�>�q����zB�Dڢ��+��9����Y�l)�4,�(9<TT^*qæ#���`�NB���=8"�� Խ�~2��]����z��|=t��EٯD�����|�>.^�Y� �DSCu0��\9*����Z���v�v�[�������
 �� ��Ny�)�F��.7�D��e��\ʙ��_����6����t9���^���D7����a��3��­�����sٛ�V�{�<I�������d�q���������|2�>b���Ծ!z�,Hl�ٺ��Vwv	�� [�b��T�h;�!2�6uȘi?[�x�~�����ŢM������:g�r+X�#��u�~�m��;��r):�:�7W�]�3�j�3���e#����T&�	.f�<�Y�D|+{�+���N����4��9P�N�.p|�ʕ2���1�1�wz ���V���'49qи��U��^΍��uH@V�!K7�z�]۾q�*5km�`�v=�
*u��*�:/S{lª�X��	+�+�b��&"{'@<4�ۚ��ʊ��Wjc^_�x��J8��-�3Q_�x��B�V/�+㲚c�4~��+t�rS����E�滨Ou�z��g��sM�[�k�x��vvo}7]����^�P�J��T}EONܖg}�挤���Ω&)ÿk*dc���ˬG��#A_wʻ�p�4�W˗[�m/\jRXS>١���o"�5��0������(#�lʋ��*mm�S��P:T�kԏqY!B�=�\��c�=/ӱ�B�
7�ح90�CT�7v���Z���7d�����VV<]0ެG�{.�-S�Q|r� �T_D�ʔ+T�B�}O��a�0EE`����ޮ�]�^r��I��(W@�38�k�*&(�77���s瓧�[�Z��n�h8�Q�?F�G�TL�W�HW9"���1�@�E�T�(z�ɋXRBl����7���뻥u�'s��,@�03��zhs����R�^k��_+�f��Uk��Vy�G�fn+id`��u���s�p�	q哢	3�LJW����,�+W���w�MhWu6#pi�@O�opvp{g��C�u�X�͹Z8.��ťjoPyg"�V�e��%����b��}(y�Ƕ�,�1��ْ<��jsK웛IPM�< wM��E;��)`d;��峄��ȝ�Z���Pѵ�U^���o�Y�-���^m���^��aA��c����*�٬�:Ռ�Ϣ61ݹ�r�r6b*���ޡL�ȫd�q�a�ر�7v�y/{��[��l����ӟ
	=Ƽ!��c��;�ڕ�ٗ�CO���rTU�-���AN��#p�_j>n���6F�$7
��)�ö7�o���\pV����Ү
�Z>�=Lt��c�n��o"db3:tS��Z�l<���a]Mz��7i�Vi���R�V|*�g�9A"�D\�S�:�o�Y"�t��K�L��)˽@�w���
�%F9��D��E��葢Gg��y�u����_U9�w�,z�F�K��t(6YNs�c��T�1�L��6�x���u��!���6;��6P�D������Q:�Ъ=^-����l�Ҏ����S�� c�:w#�/ɺ��APCK�r4�-}z���%Kl������i[��|\�z7��W�z�>K���`�z������f��?�|����|Z#(��Ԕ<���8=�5����H<��]���m�{4�V��s7�J���w�$�%:Gn���si:�IY���ɑ΅=�F��]�M1��:��u�F�z�d�y��%���n�f��f����p��PB|��sL�3kn_ɋ�8=%f֍"����GVЀ�+������}�I�u��AeNTa[[Τ�Z������}X',�\z�dYMՖ���\X�t!ӷ)^
��w��T�e�4����(+�%Z/����!D���^0Vviєkv7���mGm�'��^q��xS�r�oh�&�uAQ�jD�Zs��'�%;u�p�7;9cՙh�]#���4㗪�YVR!!ump@�Vdb����zVt_L��v��ӯ�gY�a:�YuÕ��ܭ�ٮi&�ȫ�Z��g=���q5�*��oM	;��B,�RHj�����%(��z���.��1O��9젶Z��,J	亇熧���Dǻ%���2��W6euX�z��3!�`_+v[�GR�)s��R��3�jmx#���:�� <Y��ϋ�;¸�Y���N,��f z����\Qf���Γ+:J��n��w9j�J}���P&�V��������|5��fۦے�W��7��w[�v�q����NdMncWP3�z�Nl�4��]��������ֽ�f��F!�R�Ft�2v��9�J3�k��=�>��&<�ά� �9G���o���*��C��
g㷼h
�l�hV�]�wu�IE}�:>jMٔy��xe��z��g>�dAn�Jٻ�#�e��fs,��M�L����·ofd�:����xp�l�X5���_i ��{Pr.ى�k�s�Y�_vj0�ղ�C�^����`��u���\��Β�W7��JsI�C�y�*SZ�Ƿ����W�X%�<��B8H�B�ᦟ2�����=�ʇ�^ �Kz�b���r6�(k��޲��<l�\bg;j��CFӲU���F�@������f����z&�j�(�G9y[����}�/����h$!�s
�V �9k�o�T]�*�ͮ��'\���x(�us��V-rz�J��}��ky�y�_tQ������b͔�ֲ3y���K3�_T{V���� h�o��D�;��SL��	$GG+CޤO�á34
�h����sO�w�������=@���d`�|��Ks:��!VpT	Z���|U(v��U��a�[$g��c��ϥo3%��,CDmfڧ.�cF����OGn�4�S�(w�N� s:�]F�s1u>��ı1�+Yخ�[t��W���T�-����I	�;��N�(�-���@�ގ�;���E�{0�I'�e���: (��>��
�f���[�v}�Հ㓮�:�g���	�.�jw���]%N���u �%�/�
:̾�$EZ�Ԯ�]�03D����o1��xڂ8��SB*�UQiY&�,Uز`�es-v���� :�0lj�����a�U9�.�Q����3���[*哪LkC\ l�k,�ꍌv�f���s��;6T+��s���̝l$s6��V��l� I�i�if��S@`�3�8fNd�T�eQ��Û0�9)fc�Z6vi�ʸ�9S�c�4֚��J\�ƭ2�3��*�&v14�fw1�ggl�ں�f�1�qZu�-t���1[b����Չʒ�gg;3i�9��l�`��1�6fܭYKa�ô�Tfg��c�M�a,;��lcq&��EM&c6a��L1������uksf9�un��c:X���3�1�	�9]���fd���$�8�qS���	���cf&���9�f`�~ � Q�����Q��V�s�!�z�57s�<�&����㇫r���Fl��nK�L�O���زP��ݳ��=�wG�~� .�\�����d_�켇����sq��(�'amTl�c#���-{��,�_N���_k��P�[�B�u]��gá�JR7����xR�0�*ՎϚ$w:�3n��L�}��ا�n<s���������w0HL�f���1x����>x�q㻧gp���Wt*v���3��g8�T}j��j6�_*�7BT�h3a����Q�����]����^��573(��w�#!u�}�^�G"��pot��r{�l��ױp�T.�i���{L��K��+2D!��
�'�9 �2P�G�O�o1S\f�8=�T�z��#R��VnkY$a:�l-9�Pm#�'�.�?����5�U#l���tDz�ef�}U%���z�jG0h��(��fņ����}Cfh��bHB�4��P5�\���
�}��N57��rԶ�c����ڢ���|]��]gX���襞}~���G
���.BelV��Ww�K.rt(�X&b��b�|�.q�rk��<%��:�R{����Ys���k�r�f'�Ju-k�����v�y��[�5)
K$6aK$9o��cN%��~�=���`�4����� ��$�Rǈ]=nH&뿏���T� �B�U���!4�o5�SXKV�U������u��F~ ��o\�7��_{�6�Y�K����(7!9W�8� ?~��g����#�z��F$���7X&�k4����Н"CH��eGXGER�>��b�$�-[�kR��>wI�[̵� ���R,)��*B�BUB��^���qz}��y��*�<)݌	��6���0�}�6veX�sPB�l�N\W	G/�xt����ʛɚ:B㉭���4��O���7*�[��@���]3�>��ʛ
\�@WD��
 �*\���P���е�Z�\be��E؎��^��p,j�rB��}���pE�^�AP�"g�V�!��r�$FVãA�ؐ:N�׌��:b8��5T�s~	�P��C�N�b��*�m���0z�{�=��Օ�ރ���K4�]���PXc�?*���w���M }G���1ƕ��2J/ ����>B{�¥o2.�xM�R�K�T>�lR����\k*�8nP&���:z�1�e.bo�00����z���̐�UԝqS�p�rjwf
�#<]C¬i6ȠN��;�h�Kҩ*��E
���6�V�ΌCh���k-�Y`�C�W6�C���ݠ� �f�wMX��N����2����-����Đ�{K�)�z�yS7w��f����Q�v��;�F;�x�޻�/cn�^��;7�FQ
�{�������R�Y��~��2��^c�,����yn1MW�4S�#j6}x�	��nC6���iJ�)�t����}t��fu�'T��ݨ�L�͗ �wY��.@���E������KK{��R�J���lc$��n��oQ�/qQns�S�]g^����k�:���v��=�W-����$�"�T7d�Y
�8a�_�k�޻Q�q�.7�٫����FD�jx�)�>+�4nXT�j����l��=�ф ��Q���%�'&��u��M��o��#|XmZ��2V�ɘ��T�z'|�mO�@��2�H�6ʁP#�d)�;y���K�e�\�ʱȾb�+ʙtZ����| �s��W.@}�Y�����E���c,rq��*���;N��s�,W��'aA�[2��>9R�EE.r\Iu��Q�5�ͯj�vmԂ��/�0x(9l(�oc���JL"�j���,d�J��nǻ��^��xM��=ڵr@<��L�_S�QA�Q��{*�Z��L�w���^���O*�U��9]|:}���p�C۴c�a�o4T}�
�g�N+:]�5��^޲��:/.���sZJ�P���7ԁ�;EL;�*ݥnT}.]/j��Eq*~�W���j����}�t�oзVB3ƯP펋�������B�m$�A�z�I`�����UB�Q!S��4V��:�u������:M���;����%t+Ճ�o��<��9ԷŢ���~��*|V�Y�Qgkz��y�M���G)~���ӹ�|�Ce�� ����BvMmc��ɊUbC��Ǳn�h��̬���o�Q���o{\�>��P�ʮ�1)\@b�gE*�,�ƴ�lRi+��o�ܱ\�M�1��le*�o�aAz��-H�Ud{Gf���3�V+�Z^W(�mK}a��>�l���.6,a@����˶��6T4Y͜��ś��=Qr�`|U�[�]���] ̾C�WMVS�Y�}P[���H)��:�u�A�����C�h��=55&�]��m_B��ΚS�#�H�]��*[��=F�ר���i3�J9�rǋ�\���M��S�uC�v0rG�V>*&¡�*�g���G����A]-fu[MjYZT��z\���j[���
�%F9�T2'oܭD؞���8
Z�'����;~'O���B�;��Ͷ����	�����P#�}�ԩ�͌_6w�̸_@f�0��"7W�/��9����N=Z'k�������]B�v�k��e�d3��͒qY��P�-Ix��aN���`T7bC��{�r���'܌l{�U�&z(�T��:�/ {���ȷ.]\S�}]�]�9ӄ�o�9����u{'P�s0(�s��c���������q��&5��l�P5T�֮�É�Y�'X�=���
pBW�H<e�靅��MX��]'Omp�F��
\�mX��9 ���'.��5ʩ���"�Mb"�C��:'a��y��p�U�'{7X60<8q�pfWs�G�f��h�+iX�D%9r�gKw��ĤV��Nu���˔�*w�`R���؝��.ˋ�N
�n���yLl�4p�"]K����J�s�Iv�K̊�F={A��L�L�W���pDMk�A��#����Eņxƫ��չ]�[��,z��������`1͑*Jh3m��Ҟ��/a:��������\��s2�U�P�c���.�('��y��Q���8�n�&�<=]I�8����r篚R�,On��9�zU��C䮕��b�Z��h���nw�0������d7�J�iСLg�O"q�5v��4o�%��5헊�p����Oo9v04*ӂb�C�;0O]���$[E#W��e��q�1L�U�2�_]�J �I6_(��Zq3�7�� ֌#N�@�J+�K�ü���hK���z���'xƊ�#��=�U�n^a�LFf��dt�I����A�93���(�TL�Z5����I����a��-���Pb:��@*¾͋�|F�F{Ua+ְ��A�|���?n���1��H���5>_&�v}�46:��&i�`s>-�NGy�u��m�Y���4�m�h&��V�{a���v�s���7ꝅ�(�"�*zf)K��n�v���s��W@�S����U��n��n�dz��|�Ө��\�<k���D��R� �8��5ջŧE̛�q��RDف���6g��C�: D ��E���Ew�>}/8��o7j�[�g�����1��n\��H���+%T)�
U�=Z����TTAj��䯹n�\��ip�w�)�'����:2���5Z8�g�]*ZW��Y׹{e�m�S�~� �U�%ʀi}
]mϛ�������/e�˺�B��4��*i1��f��P��(�������p/�Us������<,���+��4<`��H�c]7Wg�m+���}��J���|�u�:��z�?u���5"o+�͊�j��W��׽�����p�q���oR�9%�b�Vm�7ph.�����~�M�R��Κ��)&����bt�u��rF�	�
�]��(tp���2fab-�����t�wYS�V�"x`ÐE�v�TX����U�f)�N��D�s�7�0�Oq�F��6��m�����?�~;�.�tJ{��qsW��� ���u�Ǝ����n�HHW��3�58Wr!#��7�R�J���P��Uq��O�Qɝ\`�+��e�K,���p���zn��;梮�늘'�+\�nɁ�6�Ounu�v��p-,%�^����@)�͡��#�J���F�	�j�E8ݘ�p� w-�x�����\��L�$Z>�.�0�;B	� ��Q�*�g\��^�;K�&(��,n߼���좬������+"�Fۯ(���m���S��8�6�,����c���%k&�k��k ��Ԋ��*��z2��Y��}0�=�Uĺ�T�X�!�b�n.�J,��`*���L���6�V9���c�4~�L��<_yst��~��#T�꽶7i#k�l0��#��B��[.�$h��UrZ�_b��t+��w:0;]�CQۏjx���G6������
u�\y�������D�0��m�ݫQ�j�o!�w���<�U��|i19�73�zͽk.�|.�73*.{����U��¾�ֶd��*�1-Co,�����7���x�>z*�"rP>���̉��F�@���zY����#��	k*du�j\�ʖ�c�W�+
����>���]�TqΕ��G�u,�j�E�ԋ�M��
��gvs��Qc��-�b��.'��O��b:�c��%ܩ@ɸ~�7����GV��9ې��X.���� +��4�çJ�)*��7y˵j��#M �zu�1n���%G�ʃ��^y2�㭹
L[�9t�Uؔo���/(X��I~(2$�+�T�d�D9�r�b��nC�w�qW�=�xkT�s^{+w-^�.�R�:����6lͫ�q%
�$T���18dS�|�sZ6��<J�4�i�Μ�T=��`��Ce�EE�#�/���'R���=y������f��Ir�7�鮡�)���.7d���u����bS�Vp$V��=W�y]ѵNx�޻X��oi�Mδ�&u+�<=Df���,ce��R���{Gf���_r��\�U�Ϣt��Q/Ï�:+�'T���]���aq�c
m�����i��a��>徾�#��K�)b���XBuh��GjI�yY棩�azʤ�����ga�`z>��@�sZ�-��6,�
�4LXQx��ss)C}�]���#�2ܓe�޹��F�R����Z�qk�u񫙴�o:0-}dB�Ows�'��9�����K�M�Q���^�AyB�JC�SU��� O�(��0�
{=��8+����Z|���y����x>V�[�zҸ��S���5�P�G�2��:U�����e�a�Lh׋{�݈�y$�7WQqa����H�J����a�1��õ*��ӗ�YJ�67[k�M��l)�S~�.T�*{��E��v'T�x7����N�ɪ����KR� ��G�gbc����E��α��������nm�9�F\�LK�tO4�*�`eE�A�8:z�������T_���s�G��
v=��E��5s��h���0��[r{��`�|~5��wF��>| ����U�*�.�{=��U�N�N7:I�6�ɴC�u�YJN]K�k����U"�O�`C��8f��b֗\�a|�y�1�/������yy��z$X�s���0�]K:Ha������{���6�]/�&W#��R�gT�*oڢ�_bw�}.ˈuV*psf�ܘ��Q
��Xi�"��z�R�)�� k�����(1�t ���8ڤ��3rӥuf��$8��q��j�<-m�J�CE��R�;���u�ZSgL;0�s��a��o�cKs�F_)2����	۳��o$��n��W���+.�&�]��A}��MW]��W�|v$�ַ֗.g�V�C��U�T�37<�w0H	�#�C�"u�O��莸����;RQM�آ���]+����{����\T/�X7�ۑ|�`0["T��(g�殿J87�ܽ�-ȑ͵ff�M,�\=Bŏz7��';���f9+9�W몱�1�hbR��Q�F��w��iQ٢�2�#�X+�T���C��^˪nv�$���j�)Oh��F�F�)e���>��Kڼ�=���f���LR&x�	�6�����XZ�&r� �P����XWٱa�#c��3G�Ĕ*�N�^[yBq�:���]�r��_��2�JlmQr�s>.�	�!�u��m�X_��W�ƍ�J��1�&�DL��m5��Z�џ#���p�����H].ưE�	ۏ8ΛS�˓����]���k5r�u���W�D➳F4��O*�w�n8� ?��=19םH`0'�q�ߥ�����u�L�r����%�P�"ҡ:/���XkB5U�*X�D�o��*uGV��]�Y�CnlF��У�%���z�+��]�y��\mҙ�RW1�� n>��r��	�o��q�\�Moq�[�n�
����W�z�	ujj��1/m)���rK5ĹK	��;�2Sdn�b��*efGU��]Â\�p������G�S��n�\D��2�ܕ2ҫc�>x4�͵��%}rq�ʥ�lnR}k�1��H�����M��D_<(N����BT�D��ns$%�y&e��m�K�˽ᖝL5�I��36�(oJ8�'��%��L��}��b��U���Zj&�k�f�p�թ��]���\�p`��vk��K�/�܅T���r�|����<Q�w;�N�]	cICn�0�5<�j���wBnޓ4���-R�f����n,9��t��k�8�_V����ѥ�WliQHY�_fTԩ�ѝw��v�־L���I��N��Xa����گ���Ie�X��KT�ݞ��i��,�v��	�C��:S�J��oOc�/�Gxj�v(�b�].����3��Bu��y�6���A�$�E�}V�Pe]
'~�O��ʹW\aW�m�"�]՗1d�Ei�5�ZX�M�w����M�p
�,�_VE��K�N3��Vm��1�s1�Xz~�zkFNu�{em��6BJܴ��j�+��Ņ3 HҀR�;l+��>B�#B���;@^��%��c-�փ�V��J��);*����U-�54c�.nmDW�2���5u��G|q֞��:�N�[+vv��*�IaH�sf�|6C�u���:^m�&�9�.��ߟV�n�ܴ�J�/M*{�3-�ZV�E�]�EN���1���.s:��9ڔc�e^=:l,ڝ��*"��L|����P1����;Z��\^�+���2��HB��wh �Z��rv���=G:���'�vsDa�h�-,�@�v��uuX�en�.�H�{����ut㇬#�s'i���s@j�]٘JE���M�X��ٙ#��D�uv���m
Bn䳳��;�5m�M�K�t�u��'����ڱi*��-�{����s�;J��Sw9e�4މ{$ 뮳���S�Bū*\�}AtM1����j[�e��b�w��cr�:�j�&E������=XE7�N�W9���m�3�}�E�ә,QȖ�un8��Ӏ�����b�j�wc�rmg@3+������/k���vNvϟ0)��z��1]��Z�Y�����vz�ww���[H��{B��{�y1h�j��lG�0�h��V��t����+Z�m�)���yv.�|�uq��IW*�훺�cd�b�	y��䋍?3ܫ�
�y*7��U��ސe�X�+a
�ܧ/��������d����KN�D��r�*�����kg%�Ej�8��SF�9Q�r�5bh�%d)̆����ϲ�*gV���(똫V��q��4��a���s�XM�8c��i�ͥ����k�f-kc0cU�WD�ci�9�+����f�j*`�[���ѵj�����[��́]�`�1�cV��4�cMff���s��뽛���r��	�sp���<��U����gin������ff9���1ʁ��7Y�������z�9���v�g7���N�K��+�µ��s`f�8�yn;��g3fll�v�i��{֛��&�5wwf���61�yvvfن��Sz���ͼ�ٜ�9��fq���c��lz�����z��`���;U�nKuu���7g8���7q�o�^��t��'�h�f��Uzs���(s�k�)=�hI�Fn�)出��:���Wi������U���Q��oL����o��j����-�BT/�Z��>�{*��qu"�+��+%d��үD{�H���D����Uvc���TR��ew�N�eC�3P��l�N\WH
��%B�݃�I�\ⶩ�i�S�+*g.�*�{-���(W��K�����ʛR���
��iL�bv{��:�Ղ����]�����x�d���pC�r����5W9<Y
��O��g<��z6��C(�4���Ώ�`i�u�A��}���/��V�5��U0\�t��b]�I/s���U�5%8�Ey
�$T����W������/%�Q��eDd	��LZ��N Di�u0ۯ\=�F正0h�4��`��*x�]I���Y���%�U���]�-����}89�aˉ���= �^ɝ���:�	�
�#q,�LTsڎu�q����$Zx�#���t�%[G~�>pE��_h�QaZ>��N4_kqi+�*I�CJO{��,�ą���qWP�w~�C��n�ڏʼ��"�EM�{1�.'F����]BCF:�,��W��5�Ao>ȸ��ƭ�ڹ^��E��$m
S�ͣ1XT�$�I&�s2yt59�
�������*��m�݅���fҬYX4ѳH��󦼫X�t��d.�ӱevq�u�%9�K�őb��hv�Jgq`χ���->Ԯ�'��h�r}YJ�`񭂬d��E��j6��R���@��}� Wf�kZ����q�]{���k�{�p�#��'�"���W���Գ~���pj\��x�FZ�=rݢ�FuZ�3�5�}�7(i�>.U���m��kȸޮ*��ćgm,�IU�f��B|����'T�\Dl]u ��%	���6]!�p�\]�j����k�R����@>����V99�P��ʙ砩�L�Kɘ�^���9=��6�aE>�1���sB��I�S�c&��*�e�Ns�*-�]J����Tuu�K��b9r����p��A�b�ԗڏ��j��f۴�nBSq`��Ӭ��{ac&��:�ڌT��[�u,rf��v@^�S��-Ұj � =�3���N�;T�=�U�5�'i\n�G��s�|��FY.�҃"HB�L�N+�s^�Q1@�72��6{:�Wû)%Wc��\ù�L���B"lz`�sf�ڸ�@B�̅�]R"�y��iz��Y : *�+n|}Ǯ�:�(��
�����c�8�
G�&�R��F�f�\�c�Z����#��r�HT��8+s{$�*�#wJGf(����H���t�)Z��9{��s��-o:�Ea�5nW%�6�g���%u�#T[D��)w|�sw(�}��Eh����3��r	������ L�b�<�B�Eq��g�8�ǔ��D�-�}��D(Fu�s���1=�YZ"��Ux�� 1H�<�U�˿Or�盜,��,��b���6��|G��	*���,7O�(� f�<K��y��q{�#�4X����fE,'!��\+�"P��_Ӛ
���3� m��\���7e���8_���x��,��d�df	�)��qk '����4��0��g.6��O5#|a@m��a�{�+�MU��J#�h��׸PQ�np�Ok`��ڌyW�u3\�-����	^I�`��/̢��P읎J���Ӽ��PS̵�Y��:g���녔䓯�����K�`J��n���
�*1�T2'lr��[�jrY����Ƶ�X7P�C��q�]eB��Qns�c���<Fr:�"ܙ�v�""��3w��7Y�b�b�Q����OX4a�Tx�?,v�峟J8���Ȳ�O�NJ,fؗJʱ��G���񙽍p=�Ό�� #y�Mo$��������{��Xq�׌S�~��z�v3U��>'��e��'�
6yK�B�YH�p[C"��s��Vᘪ�h���X�d+��oJ���74
�q�z�q�-�����?bG�KW���ؘ!*���a�=�b;��jʋ�;
u�L&�]+u$�������W%�eB��p<�$��
S�R_���Da��Z]+�Shr���,��p�;˩r�"�.'!)|�(��N:�7��s��Q*%	�]U-ͭj�n-�����n �����[�o}�.f)�)���ĉp�\\�pT�6nɀ�.�9H�j)��O��\FN�l����|Ȣ/Mǈ͆B��Re�'s���=���+T�W8�/������V�W�p�P�#Yg�5����"�ՃcQ�"�*���pVc�l���r&�ƽ-R=M�,��i_gBM7���X��%�';����J����.�3�l6d���u9W����f�����^��Ѷ�d����X��� b�C��^���4�g��yRIdY���0��(��#���I��6j�rg���4Q�Bf܅����,�ə=�1-\�gq�=�i�:���] �z�47�lt`}Cfh��bP�f���,F[p�-��Tu��NcQz��ϴ%'+}���ܻ\��mB�&d�쳶6p>|��qTYO�<���7�f֖�L�NoV�S�0�ҩF�4���ww�����|a���K��H'96�-zy�=c���d]u	Hsh�Ĺw���)}��kl��������J�!)�6��x3���9�#!Ǫ���v_��w���g���}~;c=b����b~�>GG���hq���$.>��nӷK�ݾ����Y��IS\W6ˇ�W�-�ޜr�|�4o�cLu5Ǣ`�t\�dIS�ٷNġ���=�}��E�Fܰڂ����B�4:e�	��Bҡ9|�@���i,�y��W,�c��<|��	�P�����eU�N.�Z��(/HT��	�H�j$�̃Z�ݒ�%Q>���lgV9W�p[�qL�ʱ.:�C
��{}{uN��X��W�NA*)o�6ȅ��i����A�E:�S�ryp����җ�Y�}�7h�>*��%點�cs���h>�@U�>�<�UK\.����FU�B�Y
��>�q��w�^�N1Sir�V!�H�Q
D��:MU��j�i����_����S��`�yYZ���=<F[|�y]��������J�=�ຖx���ZPXt=��B�0}T��h�����'��{��ý����*�'n�q�YM�0I��or̙�Q:2�=��L<7��fb�d;��<�j��v!�{rB���H�3��o��a�!��� �F;l���C;㨤qnqz������Xi��2k�W28�q�Z��8�u��9j$�9])�B"�I:�E3�p��Շ̆��J��
_����6*瑫Yo(֩�)xE{�~�v&P'E�aq��3ΜLP{g�l�fKQWRF���xR�86�h�����x����&ɝu�Ι��<�+?Z*�ϥ'Y�(3����kGП5�r���X{20��VQ{1s��km��$Z>ː����Y:��Q�L�͓��S�D�ˢ��es�{;�q�MWC*����JH��r����V2H�>Q��ۗ��E���(;�ynB�k��VB�T{�7�o��w:����4�tn����
�=��S��{�lΎC��fg��\�/L�Q-҅{�I���|�_�Ƙ������H�6`������eM){']<5q�1
�>����R�hL�FR�
��J��Ϟ�A�{\�7�q]��Ї��D�|\}EO�5V99�P�k*dc���k����4�K�϶<�A�N�<��@�2�<�OL�Q:/�r2
���U쳉�Py�̨���T��똡�6:afU�i�y2f��٠/{%iU+6|xY�?+0L7Mv�,�D���Y:�eg���k�ԝ�����"xP�YF 4P�hzyg9�rҽ����q�0��s��͇�]e���|�D�:�q�2��.�?���Pa����v��;�\A�F��w�x���J�
�ڏ��j��}�~��w!t5J=MDcu�d�v���c棪��%��ɇ[]R��9��"yth
.��=���Z卂��ݖ;*��9��u1r�]~�l�B�y$E��D�+�DFN,�s@\��g��W*����$��i�R����]빇s�ӂ����5��o��2��_R�݀`}t���J���.�:�S@����=�P*�n�
t�K&�+�@s���y��4-�
_��c4͛��=0�°����D8s�۞[F^��V��3�LJf�w��c�G�4���˵u��r�ie�V4��CM�L�QxY�fPB7z���jDk��`�f�W�\��<�R���Gf��c%ע63�'\�R2
�r����@���\y)1�:���t��았wSY��eE�n�N
�L�����&σ�#_���h�Pa۷�x���-�ৈ� 1ڏ���{	�;�G:iNl���'״k�h��}��[�U�d:fZh�Қצ*����G�A&��%G��&l����,Zx"���B2��$� �E=�][X5�
�}[y��՘p��EC��T�`�6�ca[�{��;4]d�6���>մ�E£ֻ����2�WQ#���������ς��#��s��9�Eź��;��5�%�T�uv}}����~[3g���1=A�>��(�撛�.T���j[L�	2Tc�uC"uB�a�ˢ��b����K�ı��P�C��Q���H�
(�9�u�Z�+����L�G�\h}�\s��H�W/�����\��Q�㨡�J�|���c�=�g>�o.^FO�#6��mRJ�d�;Gغ���N��x������t�=gτ�=2��O#��Ip����7A��Q�Ԓ룓ܰ�P9 ���
S�R_���S*&�ҍ�3�Б'vwm*I*��_�Pq����΂����yy���"�c���R�!
�]\��J�/M��uo{v6N��r�������K��p^{��|:	������"�M��N��4�Ǳ�E.�T
��C�}7Γ������I�؝����Yfgnr��uNF㽫�B��/����ַ)�������7֬�mȰ9T�~��4���$
��o�����D�P90>�BY{���wG��*#^;��K=�립�Z���Ң���q��C��Ir�(���p !fhϢ�}�3g%��	�Zآ�ʈ�.�}�F&�+���1�<1	���z�!dJ�{HV�bQb�V���龑F�X3�ʂ�&�����BM7U���,{�}a�Pe_��w���"�<:��1�W�,ɮۭ��٨zx�^�͛�a�2c�z�N9���A���WD�xuڑ�L�t�>�ZY�pm9�ۦ�Cc��$�zsf��h���t4�cڵ3:jͅ=���{�t:�29�F٤ �B���
���b���я�l��bt8rT�����j��8Tj�I"6��b��TT�����}.���ڢ��SA����Y�62��_J���s�O\U�C�3�@���>�F�����ì���g����}g6\S�&1m����������8��X���=�� @�z&��PnBr��ꡊm`/�����Q]7�5�� Xr;$+
ht�u(� _�Bҡ>�x2g���{�������!�X,���b�+��c�3�U`7N.�(W�*B�BY���6�_E'��mur�R��E����+�C8-߸�veX�jX��6�˥�j6z����Wڹ.�W1f|RLd��{kt���w�9�R׉&֦��L�<t�X.��n�43+v�*Z���*պ%+�9$v�sp� W�;:�֩�FG�-m�V�(�+���.����G��f���[ xU!k7�Cu8� ��T�b��w�G�[�rtu^�r\��wЬS;����*����pb�սxR�Z�6(>�9���}~<��%�-�Y�\3���_�!\���wZ�yǜj��4��`N��,5^�@J�r%�������<|r��&�5�qJ��n�p�;�ʽ�h��ƙa:R;�=8"��S�N+�A
�3�z�� 7>��碴mõ��1ؤ���T")�!��D&}�Ú3X3��O���^����pF,�>������kK��w��\(= �Q��.79q1�힀m�������r÷�'������b����#,�R��`�R�}��3�e����q}2�:/������EOL��ڼe���E�����Q;:UTdV�g�n�0��hB�� ��G�'�u�)]��os�O���I���~UtWT�zS�K��GA�yF�娓L��ud4� �/|Q�9Y%Þ���������L��Q�8E)�R*�z+(�O��'��r�s�F��s�A��뭫KVWM��;���^CFƱ3A}�T"D�a�BJ'%r���T��IK���;Մ��k��j��Љ-�j��z��d !�b1m��$�Y��s�5�i��
 �ߺ�n��][W7i���GȈ�8kR�2b�39
] \��c��%�Y&e[]��yr��_IZ��Q��2��(,�Or�u��c��۠��M�N"����J��鎯tK�NU�::�	"{教M�3}7���u�a��*�Hv�)��m�1�˂�;��w]���D̵Z�^f�nQ���n�+�)�r�9dp�g�F��+�T8�Ը1An�c�y�p��'|ѹ:�i3v�>ٓ�U��8�*T��LN>Tj-g7ё�R�<��73���*��[�E��YE%Ew�*�}wY�QKnv�����<�ku���@7�X��:�;�I�ջ�iM��_i��5�Ã2�Ĩm�//(��d<�k����@����S;[�
��[�Yx��u�'t��@�$'�.�K�0S���{�͕`�	�V�.䑫�L-��F�Q��팎o �GZ�]fP}O��J�i�z�ncnp���H�^Q{c�=f�\���/K�H��]�nƬ�j�ʽ�V`��m,�7�3��-�_[<��n�l���8�Xܔ��V���^�/3�[z)�>GUx�[�\��k�t{��ZW�S;�nS/�h	�����=�M����6�'��J�K%VT��G�&M��<�<8�o��A��[Q�����G��ӝ�'��.�I�f���-8$��V��ڲDt�'U��ޖ�<��NΦ���i5C٢�\c����bLˠ��X7���M�ۨGnCm`�t�K�w|��3v�\So�`Lz,�iuw\_r���Z �k�hJuW�rX�Q���6��ܰl�_U�fmK�=t/I4,���v�:-Ŧ��+k����>'K��|��CfQk��j�ر���;���YXY ����z�9�@Z)��gjUm]e�R������}A."ɩp�궍�%^��8�#Q�˫�,p��|���!(�7�3�j7��-�#P:���5f��y���u��ăkb���֞�
g#�Ea��X�����ݱ[�$�.*��KMm�n�Gy4"��iGn�:�V�ɈHRo�0�Gօ#]��ʬuK��ц�k�j]��� ���3�B���'�X�:�K&�ˣ�f�d�2��ͱj�6Vpƣ��{s]ŝ�ut#��^��v�!8d��r1D�{t+2���p�<��k.���za;���� ѓ1�S�֔�\����{$�&���vB��.첵���v%X�RFd�k`���]+3*&Sy��j���(�;�2:"ŭ�x�Ef�9�o"�4.�ǩsx@����ΈU�es�J�I�6�I�c����\�����k�si�Nr�c�Ѐ�TK�
��P��NQnb�υ�W3��]3;�d��'����v�n;�;t��y�v�s;+^��1���C��n7�;�7�86I��[��7N�[�7g0w��6�P�`U�B�]Ԋe���f�k��M��z�uʍ��wV�Mٛf�����cva��7��{kz�����]�fs1ٛca�P�����;޼����M�;�Yó֜o'N�=k��WT&;�[����M�޷�i��a����gV��ɺ�^����q�G3��1��y�t�*�1�40q�-6�u��[�6�67��Ú��7�9�ޮ㽓1�ٛ`<���Ιu��q�mz�fw9�m��&��)9�j�j둵����j޶U�U4r4ġ����ǝ�w]�摅��)�u��RP�_�ƞPN����1h���뺎��u*L��X�����~��}����oU�Kt�^��tV��J���i��zF��˼�3�B�Ķ����jU����66KT��5p:/P�3�}j�Y>�F�\�rZ���Lel8���9�,��>"1\X�\Ȓ-� �QS�pj�r/��])��c��S��ږ�����2vJ�W�%&�%%�=C�*#�}"���D��܌���w���g<��s��Whg/���)���H ��m���z�y
����\O�<8.��	�~��w��88��y��5��<�t��k{=K� ;����Z���(/N�>��t�b��(��=��Ee_	�M+����W����M�WB�O�!A4���� ���M	�y��:*�o�t<|)	^e[��%l�|��FL>T�؎��U����`L���Bv=1�ٳ6�)Đ�s����2f2��}�כ�ق��"<US�uF�4Fiq�sРT=l�V�&P�y*.�zz�������m-Z��5�Р��p�l����d(@λns�\���|z�P��븮�d^
T̻��C��K	�R�,����H���lE]e��pc�^N96�9'T�W��r�x�dM��;ܷ�k�w��r�,��C,�%��oJ��#�>ܴ� d
=�L%\�9�oT�k�������UXH=n�M8@�^1�Tڳu0)�3Ua|^�̽�$��۪����>�U�Y�6o��Ռ]������]��i�{=�^���J�{y�m2��A��<V*v'�9�t�>_�(_��5a�g!���b�F������Ȝ�a���$oLy0�ؾ�m��{Ӣ:/f��U	u�[?.+�k�u���+lյ7�`����1ܵ�lJ�|k���f����|�̫�O����{5Ӑ6f�x�(��X�3�`t��w�G:�`y�E�9�1�;�$�ʳͳ�,2��uC�v3ܑꕁ�Q#	S�p����/6�I*�b�2}Bz�"�W��Ir�^ȥ=cP"�d8I��Ô^MF���{7�����f�3�{<�KF�YF����<�I�
e�9�9y�@sT{b��2p�q�{ܔOL�~h��*g"�'�J��A'��F�
=@eE���j¬�����yߗ��V�+�LA���c�@��&	ӹ/��}*pBV	��T\mWe(iȒ!3��[ϊ���~ܡ�j�GG97l�u��p>�W#@YJ)ө/��H���	�+�u�W��]2a�]_Yy�A��I�=�s�%ux�ڔ�e� ����܁D�VP��y�z��*���b�q�|0;��*�����xmF; l�ӽ2��OR�c�B�Tr>=n^mk�^�Xu���i�p��j���ec��Ih�uhC���c�+�rN9�Ksh.�������t3�yy���>�7ЌR�ƴ�d�j���n��m9�K���`
��jj!N��"2���0
�Q.�N�O�¹q~�N
�I�7J#��s��+wi<�K�`�&��.2������E^�����j^�f)�y�\p���pV�j+Dy��"&��4Ӭ�< �*����-�_���Δ9A�ʱO�P���z���G��*��!�D�>m�o���Ձ*=SC]��'Å#!�'��r'����ظ�J�u��4�0���lM��6�A{}{�l�M�ɓ#Ղq�
��V�t�"������jCR��I1���Ńhb�dt���6�٨-U��.��غǷ���Am�q
�?L���)e�Ӣ#�uz��tŢ�J鷁����������9��{N�d��R���������DA]���|:�q�j���ϋt��%�#�qj�nvW8�=瑀+*j�~��e�u��Z��$h��k���~|8 x�l(wj���`��&�Or���ii3-��(�U쮑Do�����
CAcO��t�Ժ�+�[��S�w�2��J�����y�hr�V9�-�=>bːKd^����ّ�¸�7{�>M���k��dM4CV��z7N�#�����݉Ae��G�S�8���ޜ����ѿ�M1�N<���cMmm���f0^3q�g5�+�_�jܼ���.q�P��n���!(��)�#D�B��⻢*I�6��֥Q(K����Ep(��߂b�+��c��{*��Ӌ�
@��(��<���̎,��c��5B��]^�Sc:�Ȩ�O��������zQ��P}|㢪�L!� U��o%�b���s�����)2.�W@>�{-�ۥ�˾�t����Lku��\9m.K7n���(e�� (��(�����(�眎��n���R���b̾�-
�������x�?J'_��H��M����42:��<������!�G����4�[#�E��阮���(Р�ʱ��5%8_UԳąf��JW���gs"{G;�]���1�G���+%���n�L�!�4f��0jO8��[L֛%���N��{7z��(A^�1؃��DfQ��=ˍ��DH��>ْ�Wny�YÝ9����&p�����]=����Sek�l@eQ�ו-�F�r�2��s��\tl.� Ѹ}*����.ҏ=�)O�����v��8	�(2���듗���[�s�_n4��6�̶y:�\��n򌍣QCi����9����kʴ��K	��@�p0�-��z4��>C�vJ
A�h�I����7���yr"b����u23��>X�r�p7<��Uu
�TO�UÊeE0xU�׻�ؙeH�E����͕ ��bJ����7��w/(j�8�}��Y���j=�۞��p�:���qnE'C�����^�v}�+��h�-Cލ�c��Ӿ���|�[Ι�z��l>��b|�k��N�oU�-҅{�I�Z+*W�<S��G5�+o1�4���u>��p%:WZT�gR�����_�o���-r���m���\�<Ʉ�r�~��*�C�}l����3�m��'����A�ԗ;��+�TgS�y��Kt�N��q4�:�(��T���܇�jz�V���uK��Ӿ7F�G��o��.<����"�W9.$��
���
�uK�`}oU��L����#�괥��}.��7�)E��`�	M�� +�w�6���-Yz5N
��J� Y�Q��F ��z�W<=O)k����	B��h�<|k�
�(oQ�k=�]�w�iY��.�bٹ
�7X�J�O�Jmc\���đ� S���j��/,<��t��X�ʘ��/f�a�h�A�n
�B%vr��r�Iܥ�4�3ln�9���4XT{{�2J�w���,�p����p��܅���Xl�@YO$��������Y�	K��C��M���9��wm�G��`!�����΄z���亅y�<�|C�y�g@���m��1 ���۝���t�"��T�E��"��*h�������fb�ɔ!��b����E._��jAǴ���/;�}|	+i`�V���o�_�\)g��۞[FB\y��ݤ��»"��Z�9��^��8")ix7���0Q�G��(�R�׺�2�����2����8l�"�qU�/�h��h�9���G<H�����Wo�I	 �|]�]�v�>id�05]��\�l��5n��t����2BC�R��v'��Ѯ��.�Β�ʬ�/95���{Ǣ���ԡ�]���G#S�}CG:iNl���>��b3h���;U�{�X�`@ꖦ�х�>�,GvE
�]����8s#nr$z�'�e�G����|��gD�B5Q�꜠��sINE9P8l�Sڅ�;�_��c[�u9l�u]m,����
������K4�_*k	�Y���i!��غ>
��eLy��ݹݡ��lRP�=�_�>�#��z��JEk�8:F�b��ێbڄ�>�Of�5��f���<�N��qVm3���.y�l�,<�!��$b0Ń���F�w����h���U8�zUtL8P�}e�ۖ�b����wT.��ĭy�E�ظ��\�,:g"�'�J��D���J��h~����<ܭ�V�݆��n~˽P~���O������&
t�K�$DR��GM��Al���'8!�p�Y��U`>�����GG9*���	��{C�A��P(A:u%�z)��[KVn�M��׽�7�S��@��AAհ���AEԸ�\)��v6odX�xo�cz?L��3��(��5�ϫv�;uH�.��P����DS�3�����g�>i[8/J�'O[��L�W⠭f�;tY�%��
�ռ��������ױS�y�\��ir���Ɱ8��%P��k9s�����x�Wc��~h쩜5���m�p!8TCur|�T��[W��y�px�M7S;�[�٩��V�qTFaG{ۚOan�u�����P�훌��2�}��^Imk�uH{Gw�Ə��t���te���>�£t��ܺ7��˰v���-�]��7T�����u����Ec�r�+4�9|G=+s�>:���yV*�\#h�*��@�� e�\
��(��!�yW(�%+ؙ�H�c��]�˩ �"`�r!�DQr��t�'���W�G"+[l��G������Z=���Ng�㵝F�q)jI���)���-�b����-F*n���	y}s~'i�E�ˇ�����~sD���3�ֈ+��J�%$-�����4�{í+\���g�m2�;ۋew�U�*{.���}yC��1�8��>�)��ob�b���[X�9�~S�A��m�F]�m��k��Yw������:���0��q�>�y.��L�y)��r\�[ʽ/�q�<u�����r�wy=�����;�BZ�4��Z�����r�$bDUu	u@F�{m�-+��h�vh���lA���c\�*��ӒC�h��5T�h�(+���1j�΍�[���x1�#q�3Ctt������-#��B���ᑓ9���wtl�6��#qy:�_=�m�6�����;Dl<En�竳��_b�ڄY�L��Wfa%��71j��4e�ӥ[�Q���(�@Y�PԖ���p��>��H���ڹ���3n�n�N���J�>n�nEJ)�� Pr)L������<�qkj�0Wdm<P�XMh=�=�<�s�8�5��%ћ2gY�w{��]5�iR�o[�QL��T��C���g8��Y��Օ��;O`�~���꼠.�N��n��K�H6�rj�'�9�}e���s�1��Έ�FL]�%�n� fR�@�[p.���5����f����i)ZK�ؖ�[��\]�zm�o�C3	]����wI/8��y�$(�X���O�8���h��]�Q��VUx���c!mMQ���k��׈�ک�Uy<����_�ފ �	U�nrA"|rgf����o��`)�/����m�v�d9,���X���z)����I��3��ތ��17��;���{+�
i�r�;¬��K���Yu�=Yj���ܓ�z+BPo&�J!���
�&��rfۤ�=�({/$Ȍ��M��"r&���/tS�97�pk�A(����`M��P� ������`��2�ǵ}ԯ����g��g�죗n�F]�K���T*��X?X�Q�͜dd�K���ޑ�k��P�&�q��X�m_���}3P��5=�wch�����q��{*eJ5�w�Y%�~Z��ANݱ˩Y����{���IU���;�2CHʰ���,����O��R�Ua�پ�85e?"����k�xyI�Ӏ�rJʑC���U�ѭLM:..b�V};��Mr�Z�$�΍O�ES�D���8X��0$��G��̘l҄����X�9��{��ҵC��&����=�'�4��n��m-E���-Z�a�ɉ�rsC�
9��TS�8�M6��N��.﷪�-��h��É�'rě-NU�[�T�C݌yrD���<Z���c���;�I\�<ڝtn����H���CZX@�Ҧ�\�7�+���x�6�=��m��h�x>#:�����.��p`�]������*/rS�YET��
K�0�`e�Ѽt.�����9)�e��]�(�@ŵ��C��Jw�B��o����p�v76��pR�Wsn����,�W˗ۓUJ�ٻ�n��ey�F����0�RL/p[��iH��ڸ0� *Ι���tv�;�hH\]ZͽK�tV\@��p�3v��a��MS�P����CY�����sV2��7���MC�f�l2�fպr19�m�Pm�IfC|�]z����ρ�P�Ҥ����+݋svc�5���5eA���M�ۻRY�0��`m[�M�_!����]��p������g	�>�n����|g>ODNKe�ŏ��<�=�@�+���r��6�6E��a;��
͕P���r��
T�o+�b#o+0�fMHԎ���>�@ݤQs�s�Et�5U���{��D	�^�Պ_k&�v��L�=��U�KwGy�2f���츦:�.��ڊ�=S�p��OX��e��cHS�L�-3\�J;Ǆ�}���ٶ�Vv�GJ�%j/v���~|�����P޳E.n�Ȓٲ���:�Ok�kG;�f�[g�5*�X̾�p��6�tNi�nl΁
�J_Lq��[��eX�L�@s�Հ��p��z f�R�u���+�6�e��	�Bق�]`�;�Ԯ��%v{#3���R��V����;��v�v3���،��my%f���8XB����G�|�+Q薬:����:n�%M�DWm�;,�ɧ��[�qؖ�n�c��+���`�H�Pۂ��-ʱ���=;�I��߯��M����ż;Z�뤿�5�׭/Z[��]]�����z���=t���3 '��K��#������3�}4@F�����8���򧒢}X7;5:
���dtޓ�\��#CWu�(Fi�ź�q��g,�zN%2����SKzeή�;�B,�t�:�:�[Yc����
�3��О����]��S�-bA}&Vjַe�sR�Ӄ\K��\��ٝ��V��<^�Ս�KXR��)ų/ӫ����8DS����]ݩ��j��B�!˨v�KE's��Dg�۝/�fn�K����^X@ESx�E�S;%;�����C��N$-�%M��h����Kua;u���̬���:�'f$��Vо��\�Y�cͥ����⥎8�ݶ�F�N�K�J�MXw/���jU˺ܙ��V��1����T0�n��H��ǎmA{�8��P�@L��-�_e�׵�Ɖ�םٚDl�MQ�qwL��bъ�l�4$��޿��\�ܣ�a����;�f˨,���ut��XH%%G���+lU�W+�oPU�����̣W) ��%�q�s9����"L�7��DF�x�Y�.r�B��(�84���ԕ�U�XX[7���M�S��*9�zC*�j:�pOr��8��z�cprL����j�m�k���9�v4�Ct�s���W{�o{Z+�;0�{�V�z׫N��d�8���Z��7�o04�V�;��Y��d�i����<����yc�U�i�35N9<�ٞ��c��Zݛ6�X`vt��6�׭=\oZ6��m�3NW9͜��lc��v3��-��V��4��w�8�9*��em+Y���Wc31�Ս3��ɱ�76nsev�ޞ�k�ZN���30I�����gy$���kf	;oj�Z6c,˵��Nj���, o��<j;��+�YI�]��_v.�o\*�M���b��sI�;���B"M��=�h�� Ѱ��e A�gG'Ez�d�+�����|V[ӓE��@�{-��Tp��.k�H�Z����}��/�"ĚʯyDϟ,�7�st(
�$��H+�Nz�L,r��@ɤ�ͦ]&\����5Ԛ9�4�$�L�3TP#'�*�� }:�(��ܚ�S��9�L�q2������{'k���^Ц����hP�(��S��Y4�0a��4�j�7�`�����V�9�G�b�8oP��jT��lG��o�^��	r���u���XM#�(�|gSf��"B�u��c������!R^~���7�=�Ղ��X/�=]�}�V#@���T:{�Uob��=�}n&}U��l�C՝���+�|���8�Ma�9�U������+[�6���F����l��!��:5���=���Q�M Z����0 2�\*�{C��]���]��>�u^q�{L�Y��9��=s������Ž��k���
጗sqܼ��Q�[����a#4i�_V"��� �8�.1}7LrVv^�W'����9������Lt��ro5{d��H��$4�וC�3��Y�~�5m�e�)V��k9{�)��a:i�^�*u��p�Bk-XyV��ͻ+���/6�m�Ʊ,��79��`��Rha��j*hs���	�몢k��P�\f=�ݩ.4������}�Y�ضܽ�����Z1O�T;�/�n+C���=�=X=Z�c��]�A�D��Ai�6��UY�n�/�$�a��1�t��2Wrt�"�ꁦ3s�'�z��D/�O�����O�l*�:h��"�w��F�KAn*m�;��[evRkYE�����x8>�YG�V�x�߅��J�9L�u�.WUNDt�7�Hn;;{�I�y4�ƲϓL�9زmu��M���,�HǍ�$����3���N���)wj����o��R��p�����u�:n���Z����lQ}Z�[H	N���`�Q"	9 ������W6��V�����D����2��Ij�+9��dpS	`�,Ǽ!��<���tb�������_c�^\eX=�n��XY1'8�5���#XĮqE�E�� j����Dj;m亁�CaD�����b���ԽY�q���s��`�rS�Oa���{��P�u��Y���4G'5��P1)��.��78��m�����֬ư��E`ݜqON��D�G$�c4,CTk(l�D��u�f�r4��ȮW��������D�/��V��P��C:��ΐݩ��5�v2����999�s=�9 ��EߟX	�D���$�u49ÊC^��.���8捽�:q����Mx�u���QL�
���C��9���V��*��W��+GV�����X����x�U}M��ibǛ�Y�D:؈u�vcT�����T��"�".Ұ*�]�>�l�RgbT5sk����;>od���p�{�5�(}�6��]zs	�ۢ�]!�ٵ��#ӷwN[���&9QP �� Z�}�m݈-]̲l�l�F�Y�#* �V	ָv�6�]D���Ά�ċnE�V��=%#��2��^	!�ѝ�''��O;��^iem���}Bw�&N��M�\i�c�}�pw	��6Q�9#u�|�>mi	�����tz�_J\�ߟEic��l�̾��᫖�-�{z��v;QvT�vn�g�Mx�<%uVys==n�j�٧d�>k�ޞb�+����&�_�V�2�s��˶z�o�g��0��L��N;Z�3��n���S�FwK���eq�e>Iʷ�'*�U��-�O7Y7.��p큃nR(H��oO:�j����ͺ��c�*:��-���k�}3�=/�PR��U:����^Om3�nx����)�ws�i��=���T�?)"���Ѿ��kQ[L��g�Z⪮��'K�՗�����䐲�sK�Wzz�����b-�I:fyI�+�\��3�[�sJ�3/��6p�(�
��*���fceOj\Fk�o��q�X��ҵC���&Zg����f��s��e{5`��]Hc��}�E�aT����x=�5cY�i�)n�(mi����摡��	����w���^�U2�u^T»7K0��w�ESu�OV���3^���`��P�]�1pڹt��9B�c�bV-�6�ptnu��{�m+\�-������tnl(�5�z���N)�R:�Ta��-jw�jQ��a!3k�$p�S[�	7E��ʢ3�nV�$7lcyyK��!�8KA�	�Dj��=��	�nN`��|*��@�s[a�n�IdgS�,k�����p6vh����,`�SvQ�LR�݄ݢ�ۓ�Hf��Go�%��SH{��������F0 s'X�Q�nٗ�6(Od�+{Biv����E�p5�(S�e<�ѷ3U����Lkij+e��`�����*���q)/6��fpE����n>._.�ē��ϥX{�^gw��@δnU/��k���m��vLMY}7ֻ�4��!OZ��rv�Q^vԌ�ЯJ�-)3#d���xm�����<�|[��F>�-�n-���~�4��;�'�����+�2�;TBi_c��S]��9�]u��lX�te��/^���ǔ&r6~�vx��+L�ҩ�;�Eoj��7���
R����}~�0^�F�W��B�	,=�XKZ�������4J���]�ȾFљS.:�V�����t#*���j�R(Veആ%�TL}ۼ~W�������[���}rBlӵ"W��b�F�LRw;��#7
}�C)�:�����o���u`���v>�!b4�Om�����޴�t����5[SȘz������>\���r��:����:�If���
0�X$c�W�bg:4�������e�ڽF;5�UylJ���`�nh*��3�s:Cӱ5mP���\Ҟ��������.J�O.����4�"9���
�T&�Պ�o����&��T{Wk��R����N��)��*	��7W$5�T�w�N��������q��?9�EW�����s;�ذۚz{���-�3��\�6F�
��ԴF�чVE����$���D ���ApnKaNgsL�[ˑ�m\P2F�e]eW�te"��nqB%O7}N�v{��*�Ւ7%�H���ۿg�ۗD����`���� C�=*e�V�{M]���Ԙ(̍�Ӻs}��ەv^��4��mH�&�9�5ͦ͵$�8��KC���2��!�V�HR p��t��k0�rc�=Kf��m���D,خ+L[nrVܭ�:�Vv��|���/B�w��IݫXma�˜���7�lW�9�U�NS>�{Nb�"�\�;�v�kRڬckR��NƲ�M3�9ذB��hnT�{�;j��+m�q�$����+_I�%u�����;s�)GE*�W1�������}##iEѾ]'ڭ���H��G}s.���i\g����
󵥻���.)y�C��S�Z��}U��6h����H`�VJ�?Kwޤ���v3E7/ܲF%3�%����ۛ��f�y��6x�ܧ�Ҕ^��/�����!c4�Hj�ѡ�q=��c9OQ��r�U%�r5�|� Z$K� 7V܊����ͪ���\6[t���K��{sE6w��Ά�5\%�ȇ�G|N�x/��=:��Sf��c)shY�o:6�ڛ���Q7vko��aY�[B�*O̖�𠽛�C{V��@%�dr���c4%�gQ˼�1�Í�r�w�,��WV�y:�1���QC����.^��vm��N���+���]����3�3�fІEJ�ս�Y%9��Q��(���I�oa�(��2ʔ�{s%���=��U�K*�MbwW�v�J��o�Sč��{�k>���)گ��ryEN���#�vՊ�v��|3)Un�.���̜քe������l-ؖ�[��\]�	�E�&��8J���w��%�F����SZBef�^�<I"Wzq���e�eEc��ۜ�*�}�@�uSk�`2�<���N�>� �y)m�:R�tr��{+X��EΗݹ5��V�̦\�e���
AlCd�m���{�{�Hǹ����$`�I��r�7��u���V"�䉫�W-��;rF�hBS�>�<��[^켡F�b)k����}�y��^KQѠ ��S�)Ex�]�{�����U���̹���7MҨ�.�]�۔��U��VTt���]��0��x�R
�-��i[&�];� ua�2Y��
HJ޳���c��X�t��)rj�0�c��8i�٩rz��G�u��{n�6��"I����ᬘ���#�6���{��>�4�=�{Rҩ�
���H�q��3{ykq�>x�$�+_��g[��s��z��]�g%d��i{R"�U��F�1��{F]:r�aj9ѭ���>f__[g�ǔ+�c�"�Md^�w=Z�?X��z�=l��үڡ���$KNo�Zݭi��]y=\�r�"_����(���M�_�9�9K3YW�)�g]�:.0��.u�R�Ǖ����T�|<5T��u�ԗJ����31׼�j9���W?7\
q<�]�I��������s�W��	$�&�&��h��c;UfR����n���6�٦�c���^P��"r�)�=I.8�Z���X@�h.ܧ�7ϩ^��ɦ��؝��6�/�˅z�$D�	�.�ty�u�rDnqV�!�[ڻo����s�X�ո�D3��:D�1�����^Cn�eeV�3/�o8��3��w4xᾳ�����OPM{��7��c@����m���iS��1g���!��Rgd�*S;Hp�����x:nEh�gp��mAS���:�`��p�\I$�?/L��η��nag���t��J�O=�W�+u���tC<���~�y~�H�w��G��t'):�*�����n���Vws����vV1�m>s֬)ܝ���~�+sҷ������};�RF�ܙ8����gGշ�ӱ@pޯH���k)�ō�ڮ��j�4G�ګ��`&����SuI�H�p{�*��9��^��6j�����}WB7��6�|�C��q3yO�%}��V��[4�`_q��j�C�Fv�|Һ�_*}���ܸC��oX+1�j�ʶ�e�(�5@�pU��΍)V����:�봻��ռ�1+��:�͞#ë��QW{>�^5Oc�oHF�`.�������H�Mlq���Zt�:Ø��U5���E�F
�q�vOV���iܙ�\V��b�3�;W���Pl��R��*,���ʋTF^@P���j�Y�.̩��"�HMѪ�8�'}Å��T���!�r�W(�wdk��3�k4&F�n�f�+jJv�[�8Zo��S���3� t��:l��c(��� �!l͂�>�yJi��Z�I�/{m\$`�p��c��*C�o�<��T�r�#��J�P��}u}�e��U���5�J�᫥65�aq�Ȗ�	fΔ�|�ܡ��E>voms�O������"<�+l^ހE��z��"��ޘ����#-X+2�[O3�)�Y�7-DV����X�\F*�7�V���V5ۯ m�1�.�G��:�f�۳����m�ѡ�l:]��Ȭo7/��_���<�!Vt0*`�:h�ҷ�v�JAp����Ʀ�@m\�k���=����;�<ͽDP�ܢ�X���[�ƶ�a�������7u���i�G�!w��%�J�un�ݔ�+�t��
V�=�v��-̽.ZG&˽;ܹ�R�V^"��w��yʕn ������ľh;cw�ٷ����H5��ƥ'A)��lѕ�7�\x�Fvч�ό{׀�n-{O�Z�.��],���L�c�bŎ.��2D����x:�-!�v7�J����}�*�cV1\��'4wRW�+r$w��Hr�+�*��ޓn��уUw�f�ɡ����܆̜�k��!:6��CW�,7���:�����u�@9TbCy�;�7w:�tBkV��+[�d�24�gS�8>�4n�ܣB�sh��y˦�'2���eoJ.���]]���'j�V�<��Nsr9d��(ax%�]f�ѝK�I���1E&�gΡ��r���VCeuu����� 켊�*�sKn�n���X�tt��]ԩ�n6ý��_�|c
��u�����DR�D2�uj����@��/�K�䩽�Ԋuf!���p��v9�k|/�{��C�О�ժ���F��e�e��E�KI��0�J���[0�:�u��c�÷��l�@����������O[b!=�Tə�Wje:Iׇo��4�n]M���(nͽ7�u�k�F%78D�#�D{Q2�T��Jt����[ۃ�$�����
�`��ё�z+/H�r�!rv^0���lS�]���)��{�A�Enn�X��s��2T�r�n%�r���m�%ok��{�Jc����������k��;V�<��K�E��4�Cf��klg���qQ���$r��w;	��fbts6�j�W�`���#C�Ҩ�WQ|eu[�3/6>�B��%8���K�q.V3E�I�Mf�GB���WZ���S����gnM������%)r���f�2hȥ����$S�55n�_V���e�Kr�2gXӐ��l̮�	��RBGn_���������a��8K��ӹSY������޼���hBi��s�M�ӱE����k���Zfv7և&�oS̢���8z���-<�ްv�����������7�s{���ɦt�#\�Z��z󽥤��^��85�k%��ѓ��iǸG��晧��=iZ�ehv9���򬓛�کӵ�V��Y�1�Fp��3j�Q��/5��7�M7����w����lkE�S��u���p�z�����v�X��7��^�o8l��{�ѭ"��.����oK���g;�]z��vh�V7��z���K�=�o��ow�ՙ�%)�h��Z�Vu�t��V�][Ɍ���0Uu��k��fN41��)�fT��Rg2���!g&���v��!	n۹���sw�Tᒮ����*�i��1q�F��p�������4qO��7�ި��a40��娙�q\��E胆�-�x�ۛ|E����u�OF�6/͹���m����M�x���Y��Q�iN��m^�2��ʶe8v�˩ ����0_S�EW��8Ni�iJ$��٣��+FH���6ʿVU� e"��eN�D�J���s�O7ms�l3�G5�oo&�͊P�R"�v+)��;u{��flho^�[i�Z���'�s�q��y������NS�s�y������E�oV�j{��i^�'zշI��Y��>�v��"��E���ku����T�b�=�Rj��WX�#%a��a�d�Jg�Ӌ��x�L�%�#{�0mKPZZ�]V5[V9������N�k����T�(�t�)"j�����|��U:���͑}k��W��tIR����(��u6��'+����|'9s���ٷKv�����ʃ5�I^atY�8L'Eګ�{�-�Xbuzop�q�I�L̖�c�F�v�sP�	��I��<}%]$����١��!=��L��n�2Q���V�.��=+�#ݡ��C[sX�M��Sj�>3�J�iX���*F$|*����5�}�EN��v��R7����wT�pOqX�rJ�h"�/j��7�.�f�;�����S\��I�����敬�-|{[89�A�!�9k�6�s�Y��J^l[J�oh�� �9��oGcT3�D�h3lO7T����N�g��M�[��-_�ћ�O���߁*�k�|���qU��ǐD˰�o�n�N'wU7��ۗ�*yB�C]zkq�^)8���'W�ޟoc�K!�]2�),�΍X��+0�;G��.�5�"��1P�݊��v����mtZ�J�%w\^����kN�����	�*�c����C�w��+���D�+Ѥ=Ѿ!�Y��׳G�.��*��6��u\�]��S\����G�t���}���
�Q3^|���|�'(��ۿNǚ��r,��kw�B҆��2<�7|��-WMkU٦��[6kb��l����o6��:���*a<�;��wA�I��ҧ��V[�|ۦn���=�Z�e����JDL$�-�g�X+��[0�;��<�| L܅�V|�}���W]H���qɮVV���˜��}��U�����w�r9��覶��T� D�Q��������ua�Ch���#M�m�{Q}1�NKt)���J��^��E�@�)й����Q
vXT��ެ~L}���j݇/%ߔ�R�H���:��yj�P�FI/��7�\�Jc��՗o�4��m�2�l˿)qA�HX�S
��fw�WS��ς���'Q0�>ε�`���}�����B�h&�DԞC�8�w_Tok�}{�:��up���4� _3//�6�vgK�k �ɏ:5��,ڥ�X1�X�[k:4�����9n8�\f�^!Y׍(�\mX�䑥P��������*���x<�\��NzW�*))rA��)DFV�K�
�?k4N�r+/����Z��q*'+�=�FCpۣ��M_M�2�ns�rr��K厧 ���NY�ٽ"B�}��5��er�Н�Q�*[O�y��]�n�N����Ù�(9y2cNod����CuY]�I���J���C���7Z#�/LG�z��Q9o|�Y;�ZK#6�q}�%�Ď|.��9%tTꈛ1P���Pně���dx�ڒ�N��Ǩ���9�4���&�0��LM̩�]�Ǜ�-9:r�:�w�E�{ct��ݺ]�7�ϊ����j��譸���
Z��^���N���Zt{�d�uEʁ'@���s'���O&�Nފ��(�WE���Ȱ��i�;�M���!&�ǝ�qQ���r��Q]���ENvn ��V�Yc�8�B5�S}�������{һ����y4Ս@���n3�r���mE�@H��U ����2�a7���R��ky]4��%u�@�����V�9씣�B��5���w��������ĮpZ[�˿���H��8�}r��b��Hẗ��gG#�r1~?<�i�US�)Ex�}}o��Ws�}��UZf��u �Uf����:�F��y��&N`^Y�m�m�Ư��fe�\�q b"�@�j�N�g��&�ЧA���ZDbd�<D?u���5Rm�;+���l�P<$Qvf�*a���W%����F� ��s����L������n6�i��N��ӇD�r9��+�Kl�nU��?r�#5]��j�:�>�S�W@}��j6Ѫ)Km_+����`r9%c4B���F4hq�A�`,=��7����/��������Z&_[�C�sr(*�gg��:��禨;�s��,ї׭��p��I7���QO�ɢD��2"��*u�ST C��t�tm;{�t�u��3���S�К�C���������4�lݜ��[�E.Ϫ�����o���U�M�奋m�==���3��VN��y'!�U�S�6��;{���]7��@�bq!��;���ry��d��3�l-��>J�=��s
�+*�[�t�BR���tem[���9�0�=l���Y��Ms̈́+,`�S���E�6�I^á���L�z��1��m�QN�QvM�u������9_V���1�6��|v/L�x͉k*+1�����o����\�柶��)��.s]}wsP��)ms7Z{H0<'����ٌ9���C���i��e��4���f�;�.gT0,�i�YY�n�\pތW�9��Z��P�㉵��L-���*���ڼ����w���m��w¾�E��}뤕��OZ-�&�b�!v�Z}9e:Lh�(��q[���q�
�T�	ޣ=�SY�8Sx�+t����)����-��y��ɹ�2\p��6�𐒊-#|WU궯�J�F�g-\��w|���䣣Va�����OE/)`\ES�JQG�"��W!����_nK�;��YM6�簎>�!b4��~�^��U��h��M݊1�[��"�Z�U7Ln^����������б�����M��M,�L륛�6%�H���\!��#�ntkv9�kD�/��6p�E(8�^���=�K6ܻi��"�'׎6}�U�P�XM%�ȿ.��rò��L�����yն�Vk��V-͜*�k�|����s��8�{1�uŽZ�h�2L�$*k�2B���=�7�5�c�J˞�k4Ω����E��y�F��Efki+�{�ك�p#ՅE�����S��D͑	���J��6�� �׋6�We��1Ze��+�w\a��0������8�	�"�����a���w7�@P)P�WΠ2welܻ	PN�t���7ÄUq�	few!7����$sGc5K��Fma>�k�ogG�۫�u�u&��Y������`��mu�Y��N��έj��$M-_	k��0�q��H�}���#3�Wۥ�o�R�zrk�\P��L�ԧ���l\�x��7����*rk��c�:�~�E߄C���Ϧ�>k�zP�k.6����0�=-p��nv��d�&�k̦T��Ǖ=�Ǧj��:�R�I�;�J����	�B7��s���]}�&2��6���Ϯ���W݉AXm'~�;s�;�E�3��!tX-(��*(v�k��٣�z�p��O�����}@m[�/%ڞ�9g�`\@�vf���tãt𷶴���sԪ&n��}\
��`&���}rCl˿)p���ոp�w��s�p����P�b�קYV��o��s�{������UB8�\�:$G��tu�b-L	��k��:�X4p	��������!���3M\�n@	nH|����un��vN�_K};0����0E�tq�.��`ӫ:M�������x쩈�i\�|FfZ]���iÅSra��,]dם�EY�����(����n�����1�_F6�4���f^_A��9D.�7
o7csI-��y@�qAP1��
>�.Њ_�L+�hj�������g��6h�+�j���~�ι�D~��3}���U�-�rh�sޗ��OERh0�E�X����kqI��B����f�#~��Z��X��r��)��υ��G$�tT׆����e�tv�]�0�j���oM��Ew�Ӕ��cb�r���y��G�\P���x�%ɤ�j��"�^u�~�B�3j��@�ooۥ~����>�f����"��K��kyr3O�\p���6ʺʢ��39ۜT��d��(rU�U��l�a����׳V�t r�R���VR7+C��%�����6?$�����U������g�lP�c�8�B��P<7�o�o���S;�+N�d�f���fu�>>w&����C���pJ"N�cM�7պ��]�Z�1o���
�`E֣��x8�8��R�~vy�LR�����ݤ_k�1�h�*w#��}#
���n�Z�U�τ5�7���X��0@�;�U˒rX�jYU�mjV6i;��YM2�;)�n[��>aǝښ��u��)S�9���R��m�j▟b�]�/��ɝ1�|x%k��1d����LWl��TJ7��D|�����L$�����F�Fcٙ$j��Ҵ�4�wVd(k�`KW�$���ϼ�c~��S�Xr���0v��s�����c7nO�3@�柹@Ď���xSQ}E���\��M[c#}O'��on��Jn�R�haEyT$cR:�"�.E�Fʼnf�3;;�RS��������Z&_[�u`�nEP�J/sIo��������:�P]�SdoGz��Zh�h0�E�b�������j],�!U^���vbz�7 ꓚ�т�eIf��]*`�Z��G&GI����'���!��U�*w�R�'K�⨌�����r�ӬЫIRh�{/oS̼���bqS;���s8s3�.�8��(�^(���S<�Ӄ��W�8����Ǭi�����J��
.�i馍���z5�bX�DܽŒ����Z;���w�p��Ă訧�������FN�L�Wi�)��|"��:�¯�n�v�����J��L�;Bd�Q�2�[�kOi�6<��h��4=��s
����Q�4_N�W��yN���"�G���bMeW�Vk�\�b�9C*���^���㤋�����mg�N����j-���Q���X��ފ֯k�j��\����]`����m#r�����f��j����afTgW�͔�_%�W���g=����j�b�T�j�g��MX��]cP/%����pv�]O�qL�Dվ����z��6�'�����⺯U�*�3a�����Y��F��};��]�蠼��S���7R��\&�Ft<�;�{�wUiJ�i{���HX�+�74�W��H�td0��N���Ӻ󩤪+F�?g[�M#H�5��{%C� ��2�ѱ�P���(�SU�!"�ם[4�ie=#U3̌�B�]�3[5��۫=N��:GZ�o�>��3lYz�π�t>'y��FWjO��j�Kz�)B�Q���!�kn�5gd�t���sc��īiʄX���i��U#���I���i��p��136�р��	U�G�{O����,���if3Q�3��5-VT��R��KZ5�tI[�<e>f*�E���ΑaC�8���y.��R�w(��@>��T��m:O0a;ۡG"7�v��~�Y��!x�Z������H�����e���cCa�6����[Q�+s�<�mp"�T�}vY�I���V���y���"{���l.i/��D0u���q컟m��|�������x��j0���u&�2dZ�uk�֘�
��������"�ZkX��>Վ���ݖ�.�ΡI*�0%���|�p"��P���B]1uJ�9�4����縉%a����аN	f�x4+NY
ۮ��/�+�ɹ@c,s���%��r�N��{\a�rF����R���p�w�]�LX�(��2�N�`��]���Yt�����#l	�Nd<c�mQ��q����Z2��2�LЮ�E>yvH��U��Khnپ{���\飮���kļ��t��e���V�vb�1�����������6��+*�*���9d��;�֌tأ�֗�mto�mӺ�H�7l��A���K�L]��H�AL˾M�d*�ծ��th�a��%K��K�@@�夷�� �`����d�����S�G%��dVxs�=�&��s�5���6A�O/��S�tSj�mfvn����a��^���j��Sݚ%ݶv�9�l�ʉR���m�Ù�ebs�,gAG��i���84_dje�,�%=�jo��jb��5mج��p9�$���V��i7�onqN8�_T�c+%'�_a��2���6mֹuU�2�W�E�h3Y��9��!�V<���-U����w���k�FnJ���Zٙfqߴ��vWhXr�� Jt9�8k���Ñ�:x��$˷�q�,�2H��8��`d��e��4�W��$b�/�f������b�ys rUњ�k"Ɇ����̫�⌃m��pgL�I��Yؕ�9�r�\r�i[��x�$��]׎X�I��z��9F�׏B�W7{��9�Vƣ����X̗AX{)��ʹv1�5�r�ﮑ(��MI�a;'3�ԅ��سC��)֫{���I�^PSE-<�+�͡������=:�h���[���[�p����Z&_<��M��V<�g��ù)�zaHen=�Tɯ�����GE[��峼���@\�S���Oݚ���R��ս� B�wm��`�{�,N3�=�+f�M�/k$�5��ܾI��{���۔�6�T˚ƩRcWz@�uc��d����#��Y3)����Z�N)}f�"m5�Y-$�75�NoM�Y���T(�>%1�TZ:�1U���޽y�s=���EC׵{���
�T�ܳ]����r��`�Yr���l0e�Λ�WoR�Vs���W�z�k#+L�څ�jrj֜�1ZRA�-�)k�%XZ�O{�3WZ���4��喫;�3�a���Zi���31{�z�;�OofyγQ�ڹe�V��V5-)\fժ�%��YYfMedխK�z��]kRN��-��S�kM9�4WU��*ˬ����X��tK�����fw�oie��.�vZQa��ee�RMj�L�x�4h�y�٫j�V���UKMd"���uf�GYt����-Y�Zt�b��B�:Fdʪ��U�ox�I�+�KKW���ae��Y�-%\����^t�V�[�=��޽�Y�+ɍ�\�f���*��s<��\F�J,E����b��|�!����	.�6�>LU�Y�����k��n�4�s��ˏ�}t�Ӝ�}�T��ƒSLMQ��[^
o\P�n�4�ah�/�����r6Ƨ��u��7��o����a�̡#1�v�'ѽU�P�Zh�KA�0Ȃ�L��J�Us]˴�{�ҨQ�k���t0�7�Q�Ձ�)��5�)��3�/����Ƽä�r<��5К�v*��h��|�b��~c�u��9ݍ%����|�E���9+�����p�S��ռD�^ҿNex9�I�Z>�j�	�fP�(��_Dh�N��[T�y�;��N�"wV��q���Wo�CcA_n�����q���.)�8˴�6vgN�
�r�OEeN��&��(v/j-�j-���J�g����Y����I��4A��N2[�
�W����a�n�.r�7{�ԧn1L���w����])�EΑ��9HF�GwM!����`��h�´0�98Ķ�{\Z'�=gG��eb��m���$VTB{w�0&eZr�yG���-u�n�zY��]�t rǦE-���j�U>B�opn7����dr.A�k/S[�ƞ�ʒ�.��5����a��H�W��A���ҋ�$��p��O�����X��d��PGnH��-
���cl��G��͉�	�#R���:�v����8���w/��R�H�������=�Z�u4E�IOr��'TW�M}k��V��ɤy�q����e؇���{QS�&!rk�04��z����WT�O���o��
�ue�����ϰe@�M^�x�j��A�[A{�H��v�>���F�~�Ղ���\�2f��²��5��8x��CU	١�\cyы����{��C=m�9�=&�uz�՜�?JV�X��l��0⼆���WA�\�F��by�Ì�"�5�)������֜U�g�Ȋ��SA�D��5F�g<�C9{�jߣ�$c}�ٿ:�qn�E0Cqρ�H�.��Q�[`�	C�ٳ�����e�&�XyB�a�]���nx==��;5ݽ8�g3�cˇW�=��a<�%a��\þ��V�BT�#&�r徘/E��S\P�k��ҽ�5gǔ2�jp!�6B���ݜ�?H}Zb���#��KkJ��s�(P�O7*�lݴ�[�m��hɆ΋dZ� D����S�ɷ(�;���ѻ��3�3���DWB� �ɪ��^�7	���Wo��t��v�v}������D���g9���$m�V��%_��S����B���){��'��ܥ��·r�1=���<�og�^�{(V^
U��n�e".t�7�&$k�5�or�7��>橦Sq�y��Ҭ��p�(o7Ԧ(��I��;�ֽJ�m�=��M-�O���	�C��X��&���C�7�dD�WM5�Uܻ�9�U1�I.�5cd��@�����V��d���{�5ntζ�$a��#��J,�D|���]�Ʉ�ߔs~â:}6�htU�̆ZE$MK�����!`H��BR�=��[���:�ҽi�S�B�Wb�j�Wso�a��*�PA74�ʄ�H���-��*�M�ć'#yb�r��o/���u`�F^_7W*�P^FR�F4hw�"��^yL��uz2EQ�݈����5[`�Lzܑk�l4:�j��.�o�p����3j����IJ��O]�f�1ē6�ɝ���BC�tˇ��f�zɶ�0�Z6�d�A����)�X8��3����$�x���] �R��ҹvb��\�-`B\FtiV5s����H�sr(*�ε����;��{��e���~��)�Oz:��)���2�fC���w	�gf[��y�����*��c�W�|��t�9���`��Thc�)��f�s⒤Vw%�/�*yDM��m�yB�a�T}�[�ZX���Q	�!=�2%�ny�:�
R���Up�Bs
��@]��o8�D�\�n �U�*���" sPj�C��	�*�+6��9ӢG\[.��>�yȯ��#�Uy��ЯxB��,��V��[:��g��j,qN	�嗧���7;@��ׇj-�|��G�叾�w�Ov(	���W]۞N��	�
t'����G�+�Z\6i;֭�)�9آ��͕R�D;�J��b�E���;hH��U!��r�풺��{B݀��w	�L51YFs1�]˻���`��7Y���(�²�md��O�9�]��Ȕ"�&Jl�VH�/�x�
�3�lrE�y˧e�%z��z���9͍�R���Wsky3����u��;-��/X{I��sQ=�C��i�[�[2Te7%������~S�A�6焆�P�}K�QCL��z�yv0�WJ/V0�l��G��8w/�Sм��S�JP6`���Zpa�7�:[����U]e��e^�M-ykL��W8n_�`1(օr�9�8���'��O��̗;��h��\�ťue�!=�cY�+��F�ō4��0��Gװ+��8�=\3�[�iZ�Z&__Xl���QcH=͝�ַ��V�D`�`h�BFb4�SG>��X�����RZ{c��\l]nB��,��(�LF�>I(ÊC]	��`P�-� p�9��uk�L�϶^`[w���DmkN*�C�ury��ᒆ��ǕyWj]F�;��o��@]�^���Y������a���Gh�@r;�?)w��5���|r9�mY��Z�n�Ԗ�~��7O���P#�؁��#�4zu��uh�qжב�\2�%;U���y�h�YK9e��'�f�ĭ�:����D��c�o0l���sA8>����IA�as�t�f�$!����޽�����\�;n�	M��64Nީ׵�S��$Ճ{m� Nx{����0�=��9<r�:�w�r�ݴ�S~M�|Vn׳]�{\�as�����o����k�E:�E_�*�|n�[z�v;QvZ�ټ�S�j�4�>��I׽{=cM�)W�)���}s�P�ȞT"��Ӏ��R�Jl<���k��酔\�'W����o�vP�OF7�^\��Pmm�[���خדM��!4պX�9읰9(#�$`��2�q���M���Uo#h�W���+�c��ڶ��y�w)��tz�9��M�H�P��U:�(�����o���G��}r[f_@Q�\g]F��$�)|�-�~�t�a9��-#��}VWs�/��=3���6%y��t	�Ϸ�ND�z�Ch}��~�@H��v1V�z�tk|�5ʏ&A}�&�!v�<����[�a�yAT(�5P���C�*���DJ6��&j�Gu- �>˺}��{ U/�Gr��q7�k#W��Y�5��mj�ݙ8�ii�W�&���ŻHJ���R&Q�J$�*"�[>�a4fI�)���������IrD�,�]
��'�svyl�';���(\�m�I]��\RJ�'���g�4O��w�I٢�8�5D�,��O��{Qk��:��Z�2��x�C.�E>�'^MD2"�5���G���/z;!N0Xy�ՙ��u����t/�NҬ8�|��-Ŀ:��;��=���C���	�v}�U9���(]�6ˢa@�cb�r���7��ɝ�� ��"RB3}M��IQU��s
�+]�"齱�PWۥ�Ƚ��c���#�f�f�e��pT�Dw�of�W4�*��VeQo��{8w&�f�;^��8]-¤�{�z�e ޭ��f���@�`�Br���GbWC��&����4����n��Ms�6�t� �;7k�[ފ �{�;RLcyw��#�=T�TbM%w��W�]$�%>X,��s�b���MM8�wս�۽w�	<J����!R�
H�|�J����7���v��e�1UI���/(��3O����x��ǢO�����I[/8*ૂ&����h+����Y�R����6������(s��T699qYn���TQ�����m����GhHTԺR��9��[��6/���M�PnY�ǵ��e&Mα��s�6�(KJ(�_"�p.���yE���7䏟�n��%���Qѡy,	eS�JP{V��}Pj�u�-}�V�vu��]��^����!��}��J�hܿr�$bS=r���Ϧ��Z�ӻ��)����?��>P������j0���HƸ��ɕ�V3ֳ�c6��sg:4����5\%��X<܊�q�p��SVuf�֕<J�k���;�5㍟oG~���D�Z�dD�v���Ək�C%�b�7�Mf)9���:Ug2��S�Jl���`���ӟ��zZ�>�����r�:�_=�JZ�N����v������Gj��m�S�'6��{]g;$5hk-��7o��Ru�f��t���8o�����!�oԘ�O�S�
�2:.Y�ӭW�T����84�?]{؜nïY��V*=l����6I��!Q�)f��G[k��j7ZӉK7��-��@��(l�XX����T���ܜ:��d��4���9���&ڙpD���mj̊j悳����bWt�q�Y�7 {�dv�a�c��a��ʼ��9�(��bJ���\�r���yS��qjg�L��w�GA�^Q��ۗ��*-Ȥ�9�9u+��Y��l��x�J���/-��&���`4�蒤��Pݓ�a^J=��{5����;E�=Ga���Me>���[i���X��Z���R�~;)�:�G�T��2�_yu�PV��������S�����+>���w%�{�H�k��WD��{h	�B��Pi$[*cԺaY���ǅx��8�y�>���(W����z
�t�Լf:%zBS��E9Ս�9���EͥF��ޥQU�Y�.
���U{,瓰����W�v��T��<��!Zx.Q�r؞e]w �����S^t'a�
vh��i΁r����7�� +��k�E�r��Y����\��E���sڵr@?g�2H���V�� �(��TgD떼�p�р��S��l(��;�i�����=�N(A�|�l
1��`C�C��g�84V����G��_�v�s9�u�n�e��[����9�J��M�n������!Qq=�Iow5nK�E��w���=(]�g!fQ΀�t�\�ر�#�p�+���2�  �"�.�lPs�yӎ.Ƃ�l��E�m2�Gz1��[GeNvup&�ˇ��櫌g�E*ps)���o��:�,:];x��<�ЭcV���l�@���o��^@���Kj*|R.���s��ؚѽ�M���G)b
��	��'Hd�`���W��8..����G���9�E�����㱸F�O���g��X_�:?g]�89q�c%Ǥ��,ͥW�\ B���"�V�g��~��Xy>��m�K�T�s�c��c
>��F���B�Et��� _��٣mX���a�녚OY�%��b�J���(�]��G�E�@�������eCE�ك�u_>��ZԔ#5��8]3���qj���lw�PS��F�������TE�����oj[9w6��-h�M)͑�4D�/��pB�x�(vU������/|}�c������X�rːVSM�~edu�F�G�V�D��5Q���� m�ý�N�1{؋z��!�&y�y뮥"���[��8V�Q�pT2'y�KF�J��m��C��ۜP�t��ٚ�4:�L�9��V;MV>VM^�syY+��������$��BH@�rBH@�BB��$�	'�!$ I?y	!I�$$�	'�!$ I?�BH@�䄐�$��B����$���$�!$ I4HIO�BH@�B����$�����$�$$�	'�!$ I>��$��b��L��Z�|6l�� � ���fO� ĚwǽE�j�%%B�)D�)!()$T$��TI"�P�J�QEBD�B*��)BU	"	R�E*��*PP)J�
%%)"�D
��k*��E-��"H�JH��(*)����)R�T(�RE$*��+ё*(�JTE*%R�UUU%"�!)BE!%*P�*����I@UUIH!J�(*AH� U$T����퍙 �  ���Kh˳n��vZ�m�;�:�hl����۹;��:�*�G+�k������[c��m��j�S�mV�Ke��q���t9��wd�R��	)%U��  7z� -�Wm����fͫ�5�j�qd2k��Q���viSl⳥*���w@jv��t�7f���cq2�sN�m�]��5r�"���"�����   �ʏ&�E�5΋erW[�ô�[�ӭmôke�˸1�.�uW:��.튮��u0�']xw)�z
 
CB�y]

(P��ph��B�t�D��A**
�e.   ;� �����h9�� ��t44(�СB�
:��(P�Ax���C�������7mû��]�c����vwn�7Ak(ps��m݈n%R(���.�]�U	�   ,��kZ�ݝ)V���1��]�l��B�F��H��v��Wv(CuZ(�upM���r��i��:���J�ڤI M�QT�U�  �iU�n�;ueKX����j���.�j֙Σ����Æ�nT�p�-Xwwm�Wwmt�j��g@�Us(δ�k��J�+l�I@��5��  n�����3�rdڶ�9�ʭJ����ۣH���Swgj�q��e��Z���u��)�k�������]�c�P�EPR�J���  �w�� �P릚��]wt��N��:�c+n5�Wl�il軴Ӯ��m2���)[�a�v�;�ƺS���7e�+���Wf�*B�@!*�TP�[�  2��l-��]�iZ�X�Υl5�wrR릶��;���ݗ:78ٮ�h:��]�;v�m��l���l��.�:�-!�t�ق�U�vj��m��  7TM;\���][b]�v�9F�݆�N�V��dk�k�A8q"�k�U��j�N�є56�UE�]�wu�t�-n殭x �? �*�� �)�IJJ� A�OE<���  "��	J�� E?"l���   i"LʥL�h'�Z���@:
��� A#L��I��MXO���������^�g�����$�	'�5�_��$ I7!����$ I?�� �$����$HB!!�����o�1���cרZl��sM4J�Kӻv��H�1ڷ�k�6�ɅV�Z4��71 c�9yX�*�ݩt3b6�h�͈�r�>w�<�{2�^�N���ԡǬ�i������J<�r�B����Uo*%�j�9M�J��D�nCZ�1�w&|��+sR��5x�l�����Ak�v٤X~�;�+��Y����x^��T)R ���bRDU�V<�I��2�ը6���N/fi-�� �6�[��4���Vp�0�:{�R�[BSl
�Bh�Ue��n	CkK�D]���<3�	)z[Êf�9�����~��EՈ�3m f'Ө����v&�Kqk�����Y@�Y�������it{H!�G/k#U/`L<��Y����ˎ��	�Jڻ���_f��6�㬗�e���[R-N����"�(Z�XDv�J���u�;M=�R�E�w��N�X�c�Aܬ6�m�H�)�ųee�����WhBհ���I�M0�^bj+�VF�n�;�!5������ķ&MJ��	pf0ೂU�,�`9(�Y���4l%�8ݜB�jmf����v��JƊئ�q����G�܃7v�Mn��V��J�u�v�q(C��_סI���Ô\�Q�Cn�0[x�o�@P�ɍ�}lX�li��DaMסXخg�b֑��[[��ȳ#�X�5ɗ�$���o�I�R���ܔ��QN��uU���@������9���Q5mf)�ƣ��Iuk�`��ӔḮAhb��7i����B��
�#Ѻf
D��+bn쑊HiC�)nn�6�H�e¢z���"Bh�Zu$� (]�:[Z�[���Gzp��e��Y���E+F7R7V�+2ʅ<k@$8�	�!�u��� ͭ�OV)�V M�5�ū.�b�^�=Ph��,p^^XB��՛�T�	\������Z�b���/6b:��,�T�2ZM�a�clq5���%L�slK�k	ܩ�֍b�AK(8�lf�Dd�[I��I<T�۸�쇣K5 +5�ucB��I㫐
V��oP�%��)�����(�t6�JM;&ӔS�
�
#
��q^��Ȕ�Z�	������*�[%���	qj�F����UqG*m���; ���-���C[V�U%�3!�7��)�ٸ*�oh��YE���Z���}F�ݻqi���,F�:q3`��4[mPQ*D���ĵ��e�YeXX���t�H�B.�Y�a��5tqf�t��^��Sy`Y�$.�G����%�Q}�����@����]9���f�ˡFfx*�(7�Iܣ�U �ff��M-�ܼ��Yęݎ��\�_����X�Uت��7����U��F���k�Yn��u!�fo�e��Q�εa)�k+h2���$3,n��2���߭ѡv���Z�� ͌�ˠi��6/M�m�eH��I�4�V��:�dǷ��w��m�d���H�P,�y������i��oR�`츖+.��>�L��U��V 2m��ԣYd1�Z�/h�h�Z��H��j̄�sq�Q*���z��
��U��M��[b3�n�i���b����v��X���"ʃ\���w�{�Ln'�1H*U�f�J�l�X�jlK�h�K�.A�(�ks)d���j�}YE|jg"b�����;�sJjA��%�ݚuMَ;˄Ӧ������C�v����V����m���nGn�jD�x�h�85�4m��Vb6���,�����+hȦ�w!��w��IEi���V�f�%�Lfʐ��n�+K+
+@�Y��]�[{uY`fج�mݕ�ܤ�3���(���Z��*ͣj�ț��<�^)ui��"0�.9HS:�6�A��b{F�i��n uƍ.%� ���.�
�ڥ���#�2A%Vb=T�ҹv(�V�z�7ua��"5�U�єTh�Cc�`0p���T�/nKֲ;7�"Z6]B��^Ե71�������K������w����+%�+aɀ�+�3��etI�cU]H�� �p� �ٺރ$3%��f=a�q�����ؑ��_c*j�yA��G3Ei���#+m�xy2���<p�:�Ʃ�A]���s���řzĲp�UJm�Ǘ�Z���e<K~V��w4�3�*lr��"Tѹ"�(n���H��C&^!��G�ż����6�i0��͂�˫C2:'j9z����&��I�CT9�e�,�U2$r� қ�O2W�aNV=�4�Q,\�U�%��q���ch�WU�*l����l�0a�f��HV�zkDѫ3�3F�Z\
�]<ͧ�CYm�6�!1$�,���*g$*�,(�L�N� sA����AE�c5�Ov2��A  +دK[W��2�����lU�iܠ��,c����#7"!��:J�l��+7f͸+B�H�
N�m�*�Y�[gI#U
��3v��Ъ�@LN°.�췆�{�*��DS�yXEH�>%^S^���Y�ܙ��h�#�,c��X�V�JF�7E�QЬ� #�a�Zf�F��7)��-��#a7�SwXcU�{mպsw-�e;��Z�	͖���Q�
�@)�<�U�E9fαY5��r�)6�,]Dq�L`��=��,nb�(5k����2��r#��.�ɚ/m9IQ���)��e���X�% --���:A�vU51�4!L������^$�q��*�]Ŷ�;Y��4�tl�g�×�D�N;Yt�:i�5�u&@���Jl'[�n�Z����ő�ʬS�l�`����#��X9�E�[h�yk4S�3)5��5�{�vdH7vh�ƒ�r��Ǎ�3��m^��9�E5t�Q�m��X���-y�(v��`EP�3@Aj{Am,��Ǹ�R�q�i��]��(A�$���S~����uj�
E�nĦ�M͵�^���Y��d��D�BH�,HI��q
8���\�qV�k^�T���ll��2��wJ����)��6�P�uƕ��>��û���|��T{��ZeA��w-�����G�mf3�E}VTy���
���i֍H�a�]�:��_k"�V��Q�nV�z�5�X���ò2����U#u1H��J���
��e	KoU�X�,O+C��m��3 w��=�m v2����Kj�tY��՝��-��.7bV�֚AVܳu2*:ލ6���E��`,�'Z�h_,�W4KHV5�r�l�~�Cn{2����M[J��� ;f�-��$���uE�WX�n�^�ܥ�r�ZѦ�%�J�m|�dk�0��FD�#u���������Te\����GLs.����"#%n6h�%�ndUi��#���ʮ�Xۭ�%��L�[y�e5�]�-��a�������㡠K��Q�D-d�-��툖�W��Y4vd5[H��jۖ��0�F�֒��YQC��*����)M�3N�`2���f��F��4�ה��P�P��)�kjT&U�f�tͰ���!X�ݚ+{�*bjÛn���0
��)���룀&f�V�.S�Z"̴9z� �z�[d��9{-Ƴ~Y	Ien<{��X�Z���TёH��SD���[��R�[a",���Q�xZ��62���J��)��Ycj�>xv���b�|A��^PN4�ثp1��mD��xn�i ���P��K@�(���&�"�kNl��#{I�&x��ו)��]G6T��[Wb�u+�w�����Ek��)V5ۑ�bL83j��J���T��"ô�^�Z�u�+7M	�9I�y�%a�Y��Rp(X���1�MԈ%*9�#�%��V���N��!Z�߁eƀ[�i÷[���ǀ�Ze]^h��P(Me�Tjږ����{{�YXx��Э�b*��y�j����jӷMXE����C#[A�"���U�j�Ч��CZ5�ki�z��5i��%r���:pm�iA��H�)�i�V>�(rI�ܲiS[��kX���R5���1E=0�A�VZ� jܻ� ��Hi٢��]��5K�(��+
�ƚlx�6�<{	�T*��A�{y��VodʷI�Ԭҥ��8f҂�ͺ��(2�l;�*�QV�nK� ܓ-�*�M)rP�3)2�`�$؆�Ű���d�KvXR��GE̢��*nԑ�������Ƕ����0t�@&�YM���3�sE�yVq��U�!ˏwu�щb�]c���V�U�`��c���m3chHG��Qůf�-�ږ���$Vs��u��D�dq|�H��7��{[F�J��j]�[�ִ�h*�I��e�F,�'[�ou`r��ʲ�J�R7�+"��H��G]��E(f������Y�MMhj-��&*���W��Az��}lS�=��)��wt�XC�*�m�R�YMe�5��kZhu�;ǋVn!Op�T�����ԑi��죫-=#���77E��M�Q0oeJ�R�^Hpf�(�{�c�b���+']#1���e"��Y�i�zV ����6c4�Ovc��d��u�+pb$5�.�n�����L���b�jq'WZ��T	];��"��f	P8���UM��)=+���ٖ�k��q��;�d���$���j�Y��)GO\ ��n���jX�U��ƥ[w�ȱ�k
�N��D)^��ά9�%`��3f�� �t�κC��oqȁ�+~�r�b\S.KD�B�RZ�wmfș"���MRT��Z���P (��4�;1���E-Fe[fb���c)�1%jT[�+�aC�[�،'
�����K1�J��*-(.� %���LY���6��4�%�'Fj�{4�۬[�m�����*�y
2�j�3EJ�/.䒞�����)^hғ*ãe�Ϊ��И��N�b�[ͤ�m��H���^8�tM��m�nl�.��`db���ȴ�wiF��2B�lٺ�f`���2��U�m�&�)�efY[�ٓU��j�����G.m6�@���Z25V�Du���owa�J�R0���knT�2�f�U��S�c����+LAM��̢H4S
�J5v��ti�c�a�m�,��vBƭGM] COO��kJ���[��eͲ�:������y(jV�w2�[G(�-B�[d����:̷e2(I�:����\��r���<�Fj�Kp�m���+`Ъ�2�;��$rCYI�njx���2�f�U��i^�Zqʸ�%%�a'���Ѱ��ҥM��f����*R��g���0]=[p�A�i�
zskf����b�B�n��``��y��n1�y�hl��a��Su�Fj�N�ЅiJ��V`zi������	æ���AbηX\gC�*�hǆL,���r�l�fT���!��&�n�SB��a�1���N��+ :��#�A����B�h��Z��t۲�i�(qd�1�hm����хPp).�{��5w��OFf�n�yV*Ö����!����˽ƪ�\su6�V��sT���*�Յ��]>�F�X�WL��$Rgc�V�RS�Cf)+�{j�,2����Ҝ�X�4ҭr�B��a�R%E�ri'e�<t&4��b�uKL3�L��ڂ�l)��f���7	�˗s0$��+���X��4���Nna��)z�!A�o�N�P��-�XWlE�fœ%YbY1麇)r�f1C�)$L���k[u�gwQ'P*�ZeR���H�;�m�e��zU�Os!���eL2���U��[ŉ���f��ĥ
�%ZN��U��m[�7`z����4ހ�-;sc��[�*�9�"�6iڒ�3Cٯ+q�F{Y�@a��kt()�֤�@T&� � ĉ�%]إzm�c>���8�)�`p��4��4�ڸԪ���Q��l&cu��n0n�Gf���E��Yfn��#�B���F&�ۭ�"�	#��..��+JZ�З�%��[yU�[�%%�l3w1	[�] ���)`��Y���Lcc�o̛i(�q��~�a�e�̊���s]
�ؽ�ʫ.��v+Mݘ�@GJ	�ځ�3�9��~e��Q�Օ��=E]��-0,�O(@V��m"�Wwm*
%CVI�J��U�3-�6�b��1ӧH���W��z�ʽ���G��C�U}�{�s5=4$���ЫMԥJP�XhQ��id�b�٬��+ZVٙx4�ʲ�P7x�r��.T��IV�e��f�Ur˼��_�&htO�c��w�)�pb��6$�t��t2l��t�.�$q���n��@�P���yxNrEI�8���@�n��qGJ0(rclYQ����Cdջ�K*�#��<t(��r;D�f&VS��38�F�`�;�xi���Գk&
#	�T��!m�6wr��� CM�Z1[�����p�6�&��M7Mܹ�f��C\׍ �^���eI�V�J�6��t[�����M��b���qj��X�^�{
M�N�����J�r�佬��[;e*J�T"��㸉D®�ی�U2ɽ��Qy��CL��IU�69@�4��h]'J��eE�of���zd��m��P��Uum�k2ؗ�!,���2�"N�cX���,V�h&�U�З���ỽ- �۠�6�`ƒ��	)���Rj�5ɛ�A��co�X��EKm�����C-a��A�K@͓2I��H�2��=����D��Df��	qB�ʗj�Ѩ�����)2w�$��L��*�롭�O*�]]ϸw%I�hB}�2�\��\�Sw��C�
�hf}݌fa�q`=��u�l)Eǀ��]$����f������RZn�i��]g+�Q�I�O���ޖo�Gl���,�3nPWj8�r�uM�HV��t��Wcm��H�t��;�a]jV� ����7ju����i	�A��;�۝���J_,g;�-Z��\-p�􉆌����)�p��ΝV|j�㦷`���:�9��L�3�vh�ݽ�J��<�q�e�3�_oG*��P�;������8�֊6-��Ml�)]]�7�>��d3��{�$૘�GQ7����{�s�v#ͷU�t%��tjQL�P���P��;l�o�s�r�����R��(*����Բ���s�q�t7iՌ;��n���2q�y�u��*�η�.f|�&�݄��cJI7�n�*�ڴ�ϔ�osaHl�ۿm�w_��7 �]���lk��C�08��E3��uZ����ӧ����f���#8
�[('In���KՆ�h�N��5M��1�
j���^׻w�/��tL��;�c;*�t-�Ӌ��igJ|#Ǻ�3yš4>��aT#Q9��e���k���v�c�:��-a�e�M�������w4���E�< w���Q�oR�b�]]K�x��amS�7�����6ɰ[Ɋ�&�7���9ŵ���+�0���Yc��(ev��r�NU�޶��e*3q_IFX���g��4+̽�q��#d¯f�͖En��ZF@��V���F�
R޲�C�ǫ�RXwNȒ<G]�%ok'�n|�N� ����n	 '8м�n�<z2]�bէ�Xn��m��v����bY�u�*8㬩��عi�@�\Oh�M��#�8JJn4_EVw.Nz<wI>����2�{�í�w�pX_Y�����ӆrL
�(�5�[`�q�t	��Wi��+��{x�4n�_����Ǖ� 	\�׬��	�?'c���"�
 �0�R?y{����=����)�f����X��F�C��I�v�ɳQ����<��顧Jhy���*)hr��C��'j�~(��fwT��ۼ�������trz�.f�v�z틠�O�i�A��v8���p�رM�r��;n5�nR�/>��(֣��u��PN���o��Zق��;�v��t#S�b���B����>���J�����,��{�X��u>?Xx�&�	M�&��J⩂��;@[��6-4�7�{������@��Z�7L�tY?k;�,��&`�z��Т޺t�ͮ�r�;lޕ�p���pc��r�fू�4p:���"�Sy�{�u�����t)��(�Wd��W��[��.��C�]�3��{C�ܛ[��n�F�\ȷ�oI��%��ֹ�͖vc�*|��i�[��H��xM�]%�p��i*���:�Hgw	M��v�esO�^
�8�U��+ʛ!��N�em
�	�(��8f��e5UڨoT��	WaՖ�2�ۗ"�em6�ivSC������;�8��ql��$ytVC�sR����;o�=9)[q�e�+ ՝ҹ��5����rY�CE��ǼV�<Ѽ4�{M�5]Ӯ]Z #K�Ⴓה��T��a�w��VdEm���R�NJg{�.�i�3Q.���7����ԃ�Q���< N��z��"� ��_D���˞�Ee�a��|��=�.�'%v%��Cˏf�*n�.X�h�lR�/6�7h_�o��K��[��2��1�n���h��P�F�:J�Ã��]��!�K����}�t3�n�`�=��6�NEF�Lw˳�3�Ax���PVԦ變�(�}�y2U��Z��#}6�4�}L0��v�GCT��콬EN�����.�)|n����q.�7��E�����g`K�jWu��wu���|����J�g�Γ׻*������N��\�_����p�/\��u�?^�{0��q��"ȹ�c�v�
�[���z�ǡ#a>�KL!w[�l���e� �Zy����qoX!ad��(��ݜ����;
���Ef�OC���=*�鶙���FĜ8�9��]׽.ܷ���6��U���>q�}�'DJ�)�/�"�[�㩝Cht�I�#�8td�y�'����� t(��� �"_��dM�ܬ\&֋�� ������]�U�:��"��&�$�Vs:��叇۪��;}AAc��.h�k�r)�"�.��B��`��t,-�.����]�}��Y	���ao:�3������9ua����{�R���?��S��%���)�h���)MT�"��jZ7sZ�I雙 hmuE�f��իfq{ތ�È���~�m�۟ �)�b3$C�,��8�|�G/���sJ��CU�M��9yq�����z��'z�$�X� ��$�Uot���h����u�iev�.�����Z� \2�SIG��-u��@�S�Ü�݁�f�U�B9c��O�&��ۮ�	��t�m���U�� �X��C4*V��pZ���47w�����-uJ3V���˺��Rf�ɺ�Tn��J�*�"m���s9�uh�FP[�����꿌���*��xJ�/�k���]��!���$�v��7.Ɖ�_� qj�it����)��XU���vfȮ�_�\�>�#�.Ky]*|.AD:�|��XiU��`f�U��O��˙N{���'�Njz�~�D>�����!Z��u��6�g_'�n}+M��X*";�u>�w�Y�R�	�S���Sr�Y;D���\�N�>#>�o�\�Yf�M]h�N�7b^�=���:�*����F9��߼�{�u�<��\9���|��ʵ���g2%�Y�lp�]|�T��s�'^7�f��j�J�T�3rګ�%fwc
�'P�k��I��ݞj>x�s�;o�B]�ÜB(c&ǋe�����Mg��3���M��"�7GwQ��wjY�+�����q�]у,��J�*V^r`wY����|��j�s�G�t��cS��<q�#�����[����.�\+�*�W�b���-�W�TyS��ٴ�r-��T���]���GX��$�;9ڮ]���ts��7����/���;�*]IԈ��B�s�������u=���jR�Q]s�Uc�kCX�s<�K��T�(��'i�a[��z�s櫢2�vT�oou�Fu�6��&�w��M��L+������4�/M�V��彪�����R"�Z�p��V�x湔��pH�un�:0�Ҧ���F%������]��jul�1;T>rl�ڧ:Q����k&)�{���������5�9�a[Z��8MsV�@�E���K8R�F�E�vS����ժ��aP���������5X�^:ӱDv�OV.˙�����v5�r��Y-�#�N�ޠ(vѼ�ι�3��� �-T D�V+��!��	]\�A8�XX��+�6�M���ݷ�q1!�1�ʰU���>�1:Ҫu���v)\{�e���5�-���J$pw7���,�K�o�Fk93��K��h��b77�&�d�9�38�t)��w,Y��Ž4�KV���k���NJ)ر����U�_(I�Xuݢ1�[ɮ���2��ӭ�֛@�9����t&��qs��9\�P�YT++-{Hr�Je�y�����ѧ\�|��9vx6z%z���o��e�ػpt�<�5W���*d�V�:��޽��
�r�]Ɖ�ٴhj	m,۝��e�����I�=qĜ;�r���|�n����]P��Y�/���Ιo.�u�D�������!�������(�N�q��ݷ�r��h�g����nu�|gRʄ��f�T��cq��:뮅����'se�%���ّ!ܤ����i�K6����Y�M����Q������g~�]H.�k�5����
{lp�Y=�$eY�I�חpS�7����U�������|ž��f�ow���5gr�thQW��6f�b�Jު�:�Wk���y�ȧP:%��\>�6�w>��Ub�0�Mmoj���e��� {����E���a�O*q&��r�
��b�ڬ��]�&��r���~̮{�{:�|�AN	F�oEL��d\��Fi;v��\׆-w�E���;f�][��9��(��Ր�c'Q��H���"CI�1yrʼ@]ڡJufW>.��J�L���Ueݦ��]�ϛ����2��\��-��l����
�k�Y]��Q�9��w�������t:�{�4;��t���j���UJ ��J9�`�;{Gc�c�x���WV��'t�pRu�о��.6eoV[��q��C���+R��ve	%�+�r��5צ��#oWj{B�c3q���u�U�}�p�*�W9`˾(&�����u�jۇ��̅0w�z>���>[	��'G���M�X�o�,�����l��an��o9n�V�ek��G(�&��5ؑ�f�,���<�B�d��ޡse��u�s��{�g`w���  �/�7����1N�e]<I�f͛�2�\��;]�^EW���`��8	N�Ȓ�`�D��:cA�m�H�ƹLZ��!A��J���*�N�!�3$�6���k�x�uͬ{�g_+n�@����i���]�Vj[��V�u���i]�N5�k1��������R6�Ƚ,��c�U0j�c�"ܾMi `���C��̵��8��q�;
 /#y����9ˮ�*�Hp���Z�K� \ц�ׄ�^cN� �;y�U�����F����֚�m'APߢ��^���<ē��0�+,4�ӡ�n�
QSm��L�́���U�s}��˚C��6tY��u����Rd�O9R]6q�찝m�f4�<��쾽��w������,���!�z�v["0�omQ�wa=3Q8'v@.@m�T���5���\e���L��KkVRQ�Kh
ҷe���A�U�Ngh,�6,��Z.��P��6�U�pR�7S.̵$���]���n���%�Z��[HwLx�N��1Ͷ%���0�S�A��n 6���J�) ���u�9�7���U�v��ɚ�S�����=�C��ˬ��4��qg�*Ւz�nl/C���q��:�ʙ�vH��*��k���_P(J<i3Ժb�p9{������CM�M�=x�����Zy3I-��FGt���u���L8+5Z�RWY��D�yے�BP���f"�-������[t��u2yf�@��32a����9CC��"s^Wn�LVo7��5҅d����s %���I��	��(��]m)Q�i�}��5���J4��j�� �^Qsv�e��.���ٷuܩS�Z�` ��5��BV���5 ���t��a� ܑ�P
}d.�����n�,��6���5�.:\�����ǯ������)���CzsW:�&�{B�$��΍T�dԁ���5xyS��+j�b7���̥֪�^@1hU�t���Z�~�f�m�In=]L�z�p��Ŏ�\J�{uB_gtv`�;v�]\�OuQ���ӏt<a��`VRWSH�V��Z%�љodX��t�β�˅'��e��f�!qXY�ӸJ=c+���(=����ڙ��̬ݎ�g�u��ŷL��KF��"[qe��AM�G>֕N�zH�e�T�Om��{�6��E�/:»lN`�Y��'Ք�J+C�Y��ۛ��Ϟ�r��d�t�X�I��0fDxA��vnۭO��5ˮ �V��ݶ�6��� Ր�sO��n�����\7V[���|D.�G�;����o��\�E��E1<���B�.Gf�狱Rewwj�l1u`��;��Ԗ��(\+��m�^��-��|�=j�@���U�xM�Qn���i�R�:���{N6j��kuP2nE����&�c���.�����$��A;�ͮ�	��'Y.E�1Nznȸ4s�$�[W�v�B�"���6;j=]b�E��y_C���E�S8��F�B�ɻ��w�������W�Y����c�=FD�[,���SA
���j-,k��pi8j�y���,������+��j�6��A�C��׻ ��2����妈v�#g�\�3U��8=�^��sLV9��	{��6�W�R�?��p6��P�ϻ�F�'u�LY'���u,Y��Д��q�9����{�"��]�����WL�[X.!��pbqB�����[�,8G��q��d5}(n���.��X.f��Z�c��~肭}��+XC.j�t��v�5��F�]m�H�t����y,_M������']f���J�>�F�F7�lv���gd޴���\�gK�l\��y_�W���dY�9Z�s����w��1b�ҹ��P]]�oRuo���:�k��+�c�5)���V۰��,8�"�h]tY�\����[�;Ed|�T���O*U��Ƌ�N��sUʾX�:z �s�W�go+��"��u�9�c�����/�]B�x76��`+�dwwAY]5uI���\���*p���+��iv����V�q�y�v�u4')|��ڎ+�u8gn��o&2�S��o5ˉw6ӀKRv8�,�|�NZ��oj)��֥ �QȨ]�/��fȮ:3Dz~��9���N�;s2_4ш�5��m6�ٷ�2k�co<���Ub�/����[t�[I�����/���ΧG���5w�tgoR��Z�Z��u'YƟ(t�:tÃ\���� =Ge��N��r)5�%w)�5;����׋4�-��#i�*�VT=ص}$d���h{~/�|ן_�o�>���e��R�HHH}�}U��q߽������Y��c�֣OpC�&�	0����Fp���R�[K6�$G��	Du�F��8�[�h�[�ʇ��nh´�9^W 9f��N�}��dW����>�¯��*Ұ�|�d�:`�aSk���L��� ;[5��ee�"�rc�ٸ�廛b��o6Ti-Y���w��dky��+I��m�|9���އ��OU�C�	�3��A\��x(�W\X����,�|�2���P�>��hui�f��ռ�m�s��ql�"(�^��:��m jE]GK����­4c/E;R����R91����|Coq�MnZAb�%{��z1�qа�����Bgk�2w<[R�B&�Σ�w#a��6�7Z7P[9���+d����B�ZY�����է�P�8e�)d��e���'2ya���ϱ�ĞS;����ג!��SF"�8^�E|u�M���0�٥3�8�yc{��Y(U���� ����.VU5��]h�FK��f� #�����na�㆕�W�0-�H���̩֑�2.h��N
�����:�+9�w����1Wj��meУ�<�J��mDқW�o%{[G��?rZA�3�eF$�PQFp
8h:t(^6�6Ʈuםii�%(/�F��Y���$���f���*��o.*ŉ:��-
�F5.ٗ,�ݦ�#�ȻΩe�շ��б�Ǖor(�!,���۲�;W�D��������4�T�]���t1e<��ֳv�K8eE�<�d�h$� Y:����.w�y<8�O���]�]�"Ŝ����TA��5�D���7L��;Z�U�+�+)Ј"�Բmj��Ʈ�,؊�dn)��N�Rs/��pZ��f�
iV;�VWN������pn���r�c���E7��!����͓	9WK*�f���!C��dH�[U�+���j��������-7�X���v�W'h���-6��'ժ���F��YIdAo�lT�AZ��zT�і�f�3�gU�-�IyL�7�u��]�eۼ,��ŋ+qZ�ն)��)��X#<���I5���F6[bX���m���̥ȶ'72�Y�����,t4B�'to&�͛��y����EJ�0t5�����/F�>֜�s2.�ա�Sަ��a��PoL{����h����ȫjWA������肛����J�.07��`őt����2lت8��A���p��9�����F0v�߻ �Kϙ��%m�3��01��q����C����oxɅ�C��hd����7�.`۩u�9k�h�N�h^�T�@��0�f���Qn����ُ;��Y�S}�+�`�-umHd�(�u3��V��1neNCV}��}�Nb�;bZ��c��;�S���%���,ւ����(ό��++�"2����N��e����%�0�3-r����Z5�l�-��ۖ�"bӆ@S�F6��X�mc��a��Z�P���]�c�2b�!����A�;��i�t�s�їe;���Aު�M�u:�V��P��\M뙻zg�ZA���b�\͂��68g�qk���曛�&�}΂�Y:�ݳ�t'�r��ۡ"W,�h�Uj��C�Ov1GWe����cb�����N��ڏ�as�;�����4�Cfd-���@p��Hp��!
�$ŜTI͚2��`ͮ X���eE\�0��r%���Y��K9�cW3T��1��2vk�y�_�;�����$���C�Y\�;�Ϻ���yzj�����WU��3#��&��c��.ʬ�'C�.�z�ՑJ;�ݨ����Tm�퇵mu���t3�����.�R�Ɇ<�r����Wf�3���7�9;˶��c�J�k�s.��Zcw��Ź�����7� �9�8g.�o	�Z4pR��MB䷺.������/xDð�kBNV ����,�8�C���� wP[M�t�2�wKF��OE�"�n&��g]�K�[`
/7W9��9�0.��v�bv*돺h�z��;���ؖ��p�Gh[]y�Ni�F�6�qk{��
W���;��� ���E�XS.¸��N�_�.��^�Sg^wu��)����1CR���5[oa�ڻc5.��3.L�Ka�Gnd���K�:�H�]�}�)�9Iwq�����h��5ή�`1�+[�RRԳ���fJ1[ی��]���n.����Ij��	����3���y���*����Y`Vcu�`����������Eu�������B��Y�BA�|�<*��U
6{T���i8�t3dL+���w��5��B�zI7=\���p(2��Ϗ}�� "�#�Y���#��v��������7{	�X�b���NG|̮j�|9��5�+��kT����7"�������R�$�1.�`��>�ܱγ����u�#J�q�)RƜda�4)Sn��b�le�y���W�q���1���������n������h�0���\�8�����J���(�Ϭ3h�w&\C�j�(X7r��,f�=]�(e%Hb0�[�z�[�����⥩*�-3x9CR�����0Wnp�A%"��᣶ї�`=%
�.7��y�����ѐ�����-ǋVNkj���e�ŗv�t�йQX<Z@���9JD��#��7�9KpMU|�����xzֲ���5]���(�h.K޳�uM�V�,L�&�S��Κ&W)K(��p�(h;J�6�}}O�V���w���[�Oj�RܖHr�& �s���_���iZ�GV�=OZEP�8�;{3��ĻQ���jm�#�%�0�ސ;<�aU܊6-��'��ʻ"B��[��'e���L�G�;��#K���{Γ����{��Su]¨��.�uھ�@�L���T���Nj\��܊�[��]uiīo��w}�-a�Πs�IB�wO@D���� �
�	^u�\ۻ�M�NP]�`����^)��V���|;�˸�e='9Vh�FQ�j��KuҎ��=�o����]|;Q��l�����]b���a��'[���������N�����9���.{�i�{/I�g�qИY�6s(�F���C+2�J#<��d�[�t�`�Z�T⚇r<���ʹ���9�����v]��C��;z� 	�s ��𦫺�1��`�K���	���训N��(�����U�VZ��}٠n��K]	{�d�>ZVu��PC� �w%EG�1udl'q�$P�H�s���լހڤ�i�`�"ˡn^n�gr��4��)h�O�	GON�lU�In�t�x���p'���n\q+"��v;9�Ft��g]}A�!I���!,�K��]/���O�VN��b��+�H+B����@����«0P��z� ��8Z��3+�	�9Ŕk�Y�r������w$���q���W7���R	g1ˮД1	z��_Kx�a��^f�����T��眸�y_AC�ܭe�[oI.c�.�[�%��R�����Yj����_NO��Lٖ��,�B���r�vl�v���v2`$+�:��K �Uw&P��f'u����uioM�;�r�����[���)84]fJx�ꨖ��Qg�i��Ź���H�����X"�f��E4���B�i�d��V�Ʈ�KEҸ�.�H�D��z� {gN�j�X���r��=��5��$�v�:MPh�xMJ�˲��`�tk�Nl�hv 9���4��ܯ�Q"lWiLk�Wp�u�1b����f��wOr��f�S��K�Ę)A����d7�.澇��B3JQ9t��b���cd��a��á�s����y�-ι��jt�vL���k*��K�yg
YE��r�_s�q�VdH�fWs@���8Aó^.}��#��[�f�V�8Ί�wzuB��&�.���{[�/F��ld����hö7�d"��5;�/^�(�A-[.��Sw-�G� ��e	�B�R;i����Y����r^��8�5���o�tY�fm�|$̚E�a��̩�Ͳ�P�/^��N�ic�Em� �K]%����R��p#m��"*N4�,�4�0�B�)e.����LjʭV��ܼɣ)�����\\%��w��ķ7�C��}��⺄�U�׫�%�ޒ�@��l��!���ZT^�"����F�gc+e�Z*�DK�5[9u�ؤxnU����	��C��f����FӘS��+e�<Y�-��ow��
qY�.�*_g'�ʧI�.��®��Rm�}�����Ziak5W_�f·3���]�ѽ�g��U�ll�o�:T4�p*PۙTx4�����u��#�*�����*V�d��J�kT/�*�	Ek$��sr�X����j�����.���!A0�m1} zv�uذ��+�[@N6��k���`�^����R�="�����y7�%s�ʘ�Dmka�r�{K%;��:��}V33�ۖ�t���闹7Mw79'�U��#�eZвwR��xkE򌖭TM�Y�H��I'm־ʂ��G���n�����,pCy��6��̾P��ה|�nv���%��Es�o�cf%M�P��oKK��+�9�3�2]�Y}��wI��;�O�Q��sg�T2����]��0�tS�+#z�'ڻtt.�Q,dT��.G�B��	C��᫩Y��.D�}�c���aٗQ8h8dx$�Mc7��;��L᱆�i]FN�xҳ]�	�机���%�0c2�e���ʺӭf���+.�ɤ`s�T��MZA�亁��"QR
��{ʤ˫�L��Z���)�X��C4ieۡ]֑���"�� ���j�`ыLrA��5gJ3�e&,�ʾ�Wh+Vz5�C�X�Wv��2Va�Kg�h��S/+kdâ�R�Ȗwe:�������-6�z�ݹC,T ���U9@bwө��++ �L��u	���ތKq�oi����eqd�-���kcmdu��:9P���g�͔8�rۨz��8��zf+e))�����Ҁ�p$����ͮ8�R�]��k���Ve�T�P|�iS���R����){.
�t�9܍Ѡ���zZ�}n�I|��=�\�5_[�]"c5op�'"�V��&W$���|L�G(���뭾w�x����yEkh��Yי�����ć1<���jJ��� �U`e�T�	3:���HHcwxu��FoD-��)Ƣ����ghF;���W�n]ɼ;s���VY��V94;��_XL���]K	�K�B٥�K��Z,Ω����ҝ��Z�mdڼO�v���H)7u�I��@�V�ַ��!�ʀ<��l�]WY��G;���潺��I����9��B;X��� u}r��ܤ��M/5A�̩F�;4�
���LNdu��L�ũ�ѧ�g�,=aJ����{\�7zl8���{�U���0��s�ԠY*���ַY�J�!��/ 	���=�rֺ�YpV���T����Ȧ���]���n:	p�
W�h��o��]]� �y��/���i�0 ��o�4/tQ
�q쭳]Ok)s\g:���v]e@�O�7"�.�����ٗ+'ݼQ]���.����^���;�Z���\��mE�r���
�V���ǋ���:i��Θ�;|����c�uqٍe��a�Ö��u7���Uw�&��Q����օ({����p/���8�$2�*�$����
Е	�����O� =,�A��g'8�����Y��xR�	�.�H<]�%���v,c;��<*�`Kz1��͇��mww��i�l���6�r���y�|�A$�V�{�[���֖��όĖ�Xx"ͷ��N��`��9�˩G-Nǯ�]��+X�f�fу�����|��P>vz��f6M�컟*�uir,��ɛ}WWz7�G7�#�|@d�P�Xg;�+.��*ΧN���r�H�v=*���1[x�y]|7jt�9ܻ�?
F����Y������*���ڲZ�\��N��W���w��>F��p{���:
�V��6b�!7 u�)�e?�\�[/��\f�8V*蔬��I��}EL���
f���M�u�&�ZoZ�1pL�V�TE�*aW9d� Z �q�r���J���6���vY�&d�Ž.�>Ѹ�8�P�;����@i��={��K�&ᭋf�+;�S��X��o��3�TXW���s���y�@��6�_)���ZTa�·���J�3�J*�QX$Dn���Ou�um�$3F���T6��eC:�-J�H��B����Tx�̇��Vصj��!lջ��q�� ��l��Vr _ ���c���4Q�i�N��1���xXS:i�[Z\g1�`�A2U��P�b&DŽ�Y�<2�T�v�f��MQ����0����j���\���S��"�U*�&ը��SR]u��B�\���&(�-�ZCl	�<H���Efc�j>�.�Ǽ�X���r����$|���k��ɢ���X��|d5Ϫ�R�֬�k��T�;�۽Q�t�l%��>o��[���u��1�X �2�s��v)�	ʎt�Ck�XÔ�+p�"`�Z;��֬ׄh�/�%rr�S���1��i�Wr�;)p촦��8j���4��4��Qε}�(K�o��6��7.�8�Ai��y��G,�W����f�qj�fj��@!r)�и-���3W��u�=͝���$���uډ9�,l�R� ��ͺWv�xt�r��J���+���?z��evF�'��uM��JΩE@;���zP��6����5j��wmɫY��f�l�-#�)� �"�õˣw\�V�'X��������縷�u�˴��S泗��̫*w۲�m��|S�Z�ދY�K��[�b�j�6:�m<�W:���"XAp�"�#~nmJ���J�f���׸�����(;	����=����or�<�C����u�z�f5Ǳ`n���/"�ݞ��v��u���W��*&�bR<����yx��Kܫ@m�ƾd3 Lr�A��&k�΍�v{�B�v��R�Y�� �!�{B�'Z�n�R����[�� ¯o�p��M�$r��ч8`֑�j�ef�q����u�{+��[��}@gQ�foS�#�Sa�hm�|ݧV��v�b�R�@!�=t����xJ뗇[�u���A��N#�*�ѭ�j�`;��Q]u/�6:R��.EkK{X��2��m�:�{��\MK͙6�c�w�ܛ��4Hu�x�]�˸fjV�w2�/yP�]���w/��6�
6>�{�ʽJ�i@����m>�4[���U���%��㋊���8s�.��]Gt^�ꔗ0x'�!�,�ǭ�'�f�9�s2�3;��L&p��Eq�U+�R��;0��J/-�q��)F����NK%�'�m4� O�;K&��G�P�b�ՈW�{v�y\F�r�}Df���F\y�M��X�m��d��/�n��=��*1������m۾�)����\�k�g�4%������d��| E��F��6�B��cF-��bԭb%h���X5���ki+m6 �TR��,P�E*�����i��b*1uZYDj�kVV�V�5�*m�TkP�V��ڭj#��0�eB��,T��b-�ʵ�-�h�[-���U�Q-Z����KkeZ�X����P[ZJ2�b*,(�6��f	Z���)l��J
U����j�SMW
V��bcZ�Tm+�+�6�ZԢ�� �kT���lR�����Q���-�pS"�6�,-ZƉZ�mj�\�c-L�2���Yj��)kj%�EEkKE��KJJ��e�J���Ɋ8�ml�Qef8ɂR�*���h��5�+r�S
��l��Uq(�,+ZVUX
�k�1)[J�
�Km-2�c�c��iF��/�/�����c�|�m��H  ˫Μ#ܐo�M�}�:���#�9<�SǠ��y"���/���>gS��. ��}���8�tU+'3�����I�B�V ڡ2�[��a�ԫlm!����絑�ދ��[�U�2��*�a�꬇�Ցs�9Y��Ex�gƫ��uDqH��\C)z�	�&�j���B;Y&���7��<�x&�Cy`~��r�%D��%��0Vn�v��/5'���,LJ�ʦ���M������\�gVs.���g�#ʂ��,���ӗ�{�KgA-&H�'���U�^����2�#��u[Y���`c������E3��Qe���p���xD���Њ��E�YC(��\]��d5�~k�u��R��r�����ν�^?����tBR��J*"C�/�%bD�|_�U�s��Q#�iA�<�;fM�����B�0лL-�rSL��g��C�w�5�L�Ʃ|� k�c�C���PZ�����]ޝ�1���񔝑W�K*�|��L;Te�'�)Hi6K�-uUQ��x����k{F>�'�k�3��䳭�}��~���p{��,�2��n�k/M	ע�ւ�����v��
�R嵱u�-WA6����]-�AB��U{�n���^g�V���1����d���
�Wkz�2�U�e��5�mB�����F@൧�s�]��	��Sm�:�n��;5v�T�2,����=wE�w�ίU}���5c!�ۏh�@8��ս�;�2�����WQV_j����)a�1���	�i��{�g��*��:q�'�ك���x��ɮc��ǖ�s=�ꪙ�C�+u�	�>!�[cltW�����[����vd�ԇ�����ۙ���5���fϲ�r��ͩ�IX%�x�P�W�2�������6���>���&�?K�ol�F%�|��p��,��[�C$��'֎�./���e��q���L}B��[�{��o��4	s=�M\VY�&9����o�k�0E�«��^z{�u�3��	M�����j$86�y��и��)�I*S�"��'"�;\�y�}����;�/<z�d���HVIW��n�oԈ߱t_^s6�C"�-�	�Ǳn���KB��+D�\��]�ޱ2�RP��G��t�F�Yz��)���sw'n{�+�93�S�3�N5���v�p4��+1w��^�ևK��S�{��X�j�6�΀���?u��dv�<��
�c�f vQ�dv�
	�UX@|����xIl�����`	ҷ25��돻�֯y�4by�>�y.�c�BiGB}���
�{�;���)t�T���Pz�_!/{��S%��[��(U�ԫ���n~Qj�W4�<��{��^!ÖGcUfD��e5w٭�6_%#q�5���y�3qm��7���aW9]�2`�;0�a%5n&J W�v�e+���)� ���w�zf�W����9�e�2�	��r卂�^�6V�lI�X�]{3ݼ���'�d#���}�w��]��=r�(̠*>V2E[Z4MƔ���ˌ�]�7ݖ�޺�B���ޱF�)�!���g���xLĪ×	�<�	���F�'\������pI~�X����2�e��㮳((k�ٞ�S+2��1�y(��V����J�;�eGt|j3�6Й�qڢ팫�[���{HO(�׆�(u�95�^��,=��TU��FP�:,�2 �߅'XK*ԠOY��`S���E�r䮣��9�ԧ�r�%�uF�W;7�i��;�5��HՏT��^��,����j��^Q�����3���m_���|U��[O39KT ��
ׂ�A��NQ齙GvI%p:NS�P��5Q	��Ⱥ�L��d��4M�·D2�H��-�g��8t{f��f���ه�C�,6,�i�����ծ�(�P��t���+C�����֎a����ĕ6��m�s���NR��u��n�v����քU�p�A��e>�����U��z��IO�=�g���}�3zV4���9Ҹj�Mq�v�o��4�����e�ٶ	"�XU����Z`�{Ta��d���_%�PM6��3^�����^�����>��m�i���]t��1���n�\L�G�C�_;�n~Ɵ����,��֚�e���	�"iXW��YI;��AE������.#(f�gWo����L1~�s�n�Ne@��R����Z���vRDd��*�W���6f�䏹��Z���W�����{a����Nŧ`rǍ��W/ٍ<*�0�VW=���3(�Z�l(�@��������+���.=�{}�CNۙ��r��G!x1`cv��-w�V*��V�p�K�WS�a,�H;]��r��1�F�Pu�5�ǈ����W���U�Y�O5�����,k�����E��a�{��ڡ#�^������t���Uv���H��'�6�NEEj7��y=O�㲆(b�h���%d�w���^�k�u���J��N)��5}Ba� "�vM��u��0�7�X�=_&]
�����Z8�D���صÄ���U��Ś��;J���+ojwD��]��֩u��e�QV�lr�;;h�Xt 3+{��omr�Sk�:���%*�u�Z���N.�Hmn��.�9w*�x��EIك�i�����n[������|۝׭na�/վ�ô�}c�xE�u	�;�T���
4F�iG�7�)S�=�-�J��;��n��B|�)����)���|Y���i�!=)Ϋ2�y��;\�C}�����m'÷��j�k���n�����)��!՞}��J�m��}~��3f�Sf��:;q��N���O����};���]"VP(W�|J���#�����i���dPQ�����}en�W�e���f�#��5�]��5�]��b�Aq)	��`�)�c�@�$����o��S{�ڄB��2&%�05׼�S�˙P��Vx%��x�C��~�����C!HSm~����*O������|˝�3�|�KR�TI��e���2m���w�4r����D�i}�|��uv0��`�+ņ+$yPR��)o��~"�nk�u�/��� ��Pb�(i&�R�X.��8-Y���mPzy�`
��"�^yk�][����3�u�8�|�Ȉ-�yPO���WE�^ܯ
��6v��S�am�(���c7�B��oL��%<F_J��fz�k�Q��1ExN������om�@	��wu����HPCdHdO/C�;��|���b)���ȗfMu�Z�}Vj ���6����$&���{�o;�ui��˹����SNwj�i���osOJ�\`<t鿤ɔpT��t���/�%bD��b��}Sr�����ZɆ.>|�[�E�'��S����ha�.�- :�&ZύQ����hu�sxS L�v��F���Jn�g��l���)�ucj��	�L��#V7�4���閰u�ц�|wf�췭�1�0�04�쮧�7jzV����g�})Xr�7V��^@���_N���8�Fܺ.i�g�帴Z���&wUZg~�L�:K$T��֣)-K_��JL��;0'���+���t�US�
�B�К��-����������ӯ;[|��X�����[`�}�s�?U���8�����%������`�J*�[�e���a9���+���5�K6�1�}��2�>�ʨy�:����r�C��UG���+c����p��;}��B�mx
�j�"y����h��hCu�c�l��~Z������)�������u����v	~��$u�����q}(V<�%o����Ϻ\h�%ֽ�kǯ����G�O͙[,ݐ���xh��}\�w�yQ�r��.<#X�u��u����ElD�V�ʏ��nz�Fz׆K��V�z�30�.���
N's�r�*oTy�2�j����e.�Mߌ�dP���^�G(-r��ȑ����g�����!�$�ESe�`$��>D��DY���m�z2+[�d�n/%yݚz��zWk�� cE1�\$��s�>�A���oF]65гgX{tO�.�2g��#��p��^�Z���w��y'�_�*,�D��Ms����h\6� �����*��^��nf�g�������F��V�8k�L�e�Hv�/l+�)�:zj�e�����e�� �>�z+>2ck~uZD�q{VK�*
��F|�SV(z|����Z�h���/w�y"��Bc)�̽VDϩ��߾銀Em9r��R�b`�FE�����Vh���}����kR=�h�_�#@��V"��E�P�Tls��A򱁞�����3�t tX"�Pxw�{ښ5�03���x���]v�+�V�̭<<JIhc%.�������#lg���a�I�}��.�;�5�6|�vc<+�㮳���r�P9v$���s�+�aO�o���%�ITxM��!bum*�^�օ���u��E��V
���7<=&�畊��Ù�7Z
-�C���G�:D��z�j27�iul6�r��2�������*Q�F�vt�חO�Jě]=(ۛm�������8�yV7l�vL��`�ܴ2]���"���f�t�����=IX�~o��ɋ��]�2>������_���ϔ�<��L�T7�,H�HY:�YW�	�;ZR�pm3���G����{��h^Uy\�no1J��$;�5��HՏT��CSkN1Sw�L���� j�a�*���G}�HPF.�O39KB	ގkK���uZks�Ny�=�۳V�Z�P�:�*���[��ئ��o�_Z� o؇S��UC�~{�Y�vz��	������o�l(E��}j�,�Z`�{Ta�tN��u�v�j_7t��B��ނWg����nq֙�'�[�%�©|&���+t��{�62d������:�w���LZl�Ij!Y��+q�~�߈�+
��e$��s�`�VW��!c�G��=|�����[���~Ņب��By?J$P�݂�	;2-�K��"[�y������N���3�#�r�~q{%a߇Sx�>	z/hrǍ��W/ٍU��:{����m�llbW��MA��Q=_5k�Ⱥvج?uN�ˎ���)�
/�έ#�x"����=Q|j��w�]������-{��B�Gۤ7�v7���نY �ᠡ;����#ݡ�KVZ��F�c�5.��zY�ͪ�+����:��c�
u�4�T���V��.N��h�8:�kz~��|���؞��t�pĲ\�}��=3#;�{W{O߾]Y�X.��ZR?��%�}�L�(��+�q\�F=u�kg�\�Y;��x�iZ=Xz*�8o�.�#>iO5+Zaw+��5����5Z-��\)U`S+v'�I����|:}��-`%�N�=�C`��}-����W�yZ�c�.�]�mG%88��8g���6G����X;���0�ݓb�yzG�ւ*�s�Q��M�{�-X;�7����<y	����,Y����v�R��|��@��(�x�[�ٞ#��z$~���PWd���YK��)f1î�6���^�w�g�' �տ.~m�w��r�Dy+����QUٮ8��;�E��/a�Z��7-�U/�y��w�e>>�ꔷ>qM�##��(�`O��+B�0�)�
;Xz�j�/��W���+m\��� 	���kj]�J�����kw�^���S�b�~��t.���ҬzE�M�Wn�!k6��A���J�j
�w�R�'|�^�qO+,	�
*�u����T^�X)bi�¾�v���c}�� �غY�)�n�kz�R6�5E3.@����יM_9�4alK�#3;4�+R��q�p�K%q3z�v�at��A��}��x�C��]�w.Lm#9����4Gb��n-��Q��c���DZ=�O�YƏ9��t�9޻h��neԽ��W����0�i�7��<�x&��o؍���i��%��_o�v˄���4����i}������3���`�<Xb�=뭍�_E����bX�����\�e[�A�$��Z--%2����P�=�l�#}���vS����pad�{��2��3�W�+�%[�@��`�ǨCt�d<�7x3]�6�<�9��M�V"o8����tçK�.��ṄJ�Hv����H����K�T�����Z�]z�K�~<�Q��Ċ0f�rX����rSL��g�ZnK��]m�-�ͅ�׹PޖN��9�I�_����wN���p�H�M,�	����\�'�Mx�h�U<�;��s�>�Q��Z�U�X�5�,��������g�})_�T�j������P�+��C�U��x��ѡ��>����>v�<%'=�7��*�^�������}�v�/�{�t�q�JW��K�5k�n�4�M_;K7ltW���˰��w��qTo"�C����$�^:�?�����;%��U�!�%&@j�	ƐF��1賹l�/jr`�nG����-ŧ��4���;^�c}��]p�3��;�;�<��(�3yf�O:V�V5Ґ�[F�Oq�e������8��u�ٔ��V�^���򹚏h�Rj�6a��t�Ѻ�Âg�v���
ΰW,�C���	NVWQ��O���z�n�Sk9`���$������f�N|���1�'K9/�ڵG�:{�/���Q4n�wQw�y��Ƽ��%�M�� ���p�����[m�Ae;�*ub6�$�4�U�w5��F,�W�u��NP�Qb�D<PU��o��=Ո����*ꃎvH��7e�"�w�	#�v�*f6���d�^�h�����o$0vۮ�X��̎�ρDFW���Lsn��c����Eӣ��f�����{���*:��֫%� 5w��@�u%Ƶ�[�D�������\)�8�*�2��A,�Q���Za/��զn8�`潁	P�����r�i���\p��k����Wl�G^L�|U��;�u��JK���ҧ*�g�L��k�yb�J�q�����Wr��]g��-Wl&8�f�uMř�p����e�+�-m#�u��=��'��fPJ�`.�<�P5t�|;��6uM���ʘ�ˠ����rf��G�}v>��:��7�8���ҳ��Vh��<�$:+�s�J��[���d�Y�K|;�̳`�i�,;�B��������4�e[ʴ���wJ��RWsQ61tͫ�����̕1V:YCP�+��=6����(��=r�vbE����9γ+�%�*�i�E˻S)�o(��L���7�g=Q��L$7�y�W�|���M��:���v�at���G�gQTyK��1*��д3X�=D�89���������6=A�;}��]fĠ�8��B����O�S��lhS:ˆ���.���' �IK��=&��<EՋ�3��`v�N�C����A���+ڗC�����w'[��t̢Es��O��D&9��U��R��֭�9���\n;إ�R�����T��I�Lh�7!�X�J�U��ǽp��m�MK"��Af
{W,OXJLB㵨�w]���8����M��D)U��+o�/&NWT���{`t�6=��� B��Ks&�u[.��`����n+���y�5��ȮeM����PP���q�`���������X8d�������d�o��͛����|7۷NWzLt�/P]v�M���g�Žx�8�yю�K���Om<H&,,�p��2
�:ڭ��ҋ��T��W,][V�c|*ˮ혦X�C �����wnt:��=�e�жG�s
�����-_v���ߒ��C	�*�_Nw�>���Ku��_�m��f-�@��8=�y�Iگ�e;�L��Y��}���OKV-�����K�ʖUmAj6իE���J�)r�V�E�[l�ik�e��R�EJ���J�R�e����6�R����Xڪ�UTnfWQS��c`�PQ�B�QpqJf\A�hRգ��dQ�*��jUV��IZ5ڕ+hV%kkB֌k��lF��4S)[L�aiDQV+ih�Ɩ��V�P��%J�)\k1E�b��ؕ��j�m�ʶьG).%Q�TZ���F"���-5\�Qr����Q
�,q���[�-�J��[(-�Zш�Օ����cm-�Z����j�����#U[Z�ĭ+E�҂F-��kF�QkD�mDA��QLq2��\�PeZQ��aA���-�8+�*1�mQQ��V����iA�������b�
e�)j�UAm�1Q��������[[-*�Uk,j[h;������wx��,��򋻻[m�{3�ʹU\`*ӭ7,u�Y,�u�Fy���I����:ev�Ν\�C�y�gq�s�{r���;�Y.~��p�����𒲥�x��Z��2��N览ǵ��s%K��S��h}ҏu������ub�3�.�{:��%n���W���� �����
7�Ә|�wx����EcT�3�*���[]VЇ~Yg�K{e?+������FB7�u7��R���:
����Z� �D����������\�䕢\�!�9�s�}Z/��E䧞����>a���Ť�9T���UNYn�o=tE]ל͸�T2+���Sy��v�x�']c��t�f!�zJ� ��uoXyj�7UP��tx޺s5����7�=�O7�&��)ˋ9���C8�I���n¡��Y��e6�Z��5�'[Ӧ����d��u��+6�r�]�0+��#fy[N�N�d��9��o�����`��%y�{��z��O�Ճ]i��宫H�Z�w�lɂ�T��3氒��4L�
3%�ymzwF]�$
h@���[�9X�R/��[P�!1[^�̘<����WµF��/����>�����=MS�x�.�8M�ip�f^O�5Z{�ՊC�� ��I��ù84;�%h�r���MiY�� ]LLWIV
�9we�o��HTQ�2�c̀&u�95yG��-<�I�[O����S�{���F���Z7�2�K��ܭ\��{�	�@�E�V�O�2�֋����9|��(����f���^�3B=�y��Uڏh82�h5a|v� F�`��Uo����hwOV�d��L^�ۏ�G/9��Y7+�#�>Y�(O�|��Nj��@��veV����;\�}��oi��r8���~�Q����0�zY2��a�U8��N�����[��q����^׃=:Zca��O8�����<��q�L����T7Ҹ�BGzB�:�YF O�y���KSr�^pw�}{q��pi+�ꏢ��f�M �[�j;�k�L���F�:�5�ֈfx���kw�{I��F���ҁᏗ��U��V��)�C���8c�������N��stA﫵`Xg�5b���RQ8kq��/�tL�O��4M��
]��"'|-���?[��u����O�kK,���k���|�W�:*r���13
��j����	�4�����J�t��Xo>u��8�o�,�&�ۅ+��+�h��Z�3������&L�'3��KKnsWsE�cb�E�R�o[�1��v���W�U�J�;�rĘǱ�VN���y�G�f���^y��{�����
��y����4.��F���GG9z�eZ�u�Iꃗ��X��y�q����5�7��>�����go.�z\>�V�Y���o3Ɣ��W����N�F<kJ�YI;��BX{M���ɛ�[8n��P���Ӫ��M�;���{��J$U���#��ڎ�$T5�����A�|��m,"�́T&�^�6W�+���{%aަ�Iش�|��P�u���Jw�T�_$f�c�Ƶ*�fl�B�P ;��|E�C���?u	�9qО�E,{��ž�.{�Q�]r�m����c?b��u���JĤ�h�/j���Ϭ ����k�9�\��9�8*W�c�K�0J��*�#�:��X:��7D����pv{��Wfd���;��D|h;��e���T$��a�TV�c��*�U����f���S\r�c��I5�ݘrڏF���i�2�X��{/ͳ�z���`"�nɿ�u֣�P҈���骳����n�Fm�*�g�e�:/��N��Ǎ�Y��f�s����)��>�@�R�q:��e��˩�촩�'��]��;FBGC�Z�@n[���cz8J��X��'JY6�ca�틮�W2)���ヱ���E�Aϱ�*�΅N��2�ߙ�w�oW�n��n��Ʃc�QGc�T��i�G��:#o\,΋Nۻk%�Y]]���M�zh2�Ӽ�T]Ia��y8l*�P�f���I�2M��e��g��v�虙�d�7��]�sy��ݫ7u�gXF��A�U�a�C�<�F��	L|�Wog'�n��Z��=�O}�Tqy�	��%`(W�|J��h�a���X����̮�t��f
�`r_D�T0���H��5��šJ�Z�p?�h�d�M�%�^�O���d�ǂ�]:��[[΁�L�U�dZ%�05׼�S��*U���H�&�>�r?��%L���i�$D:)�`!��7��Pޯ���x&���޷����[��u�E��Y<N�Z��F���`߲��?9w�tx8|WZ	��;��y���������̞�3��x�&�a��x�X� ���P�M)M�UŜ����f���;u���@q��Y>��!���3�+���Al�yj~��Ux:�GGc���w"�8���z��ۡDd���m��"8c�2�
������9)+'��X�m۱m�d�[�U��}��^��A�%<^9wRʱ\����u9(%k����K��]m�,���v�8TT��y���<�Y��c;���SgE���s,��ĮT�N� �[�ʇ���7���QM5����mA໣ý����>j�J�}�Gp}���k��E"fN���*����@�Iy���9=N�(��oR��E}j�ľڱn�9�:��G*\�i�ܝZ��χ\G=����[r|��V�ʱ���&-�J��5cp)Hi<�/�U�޻����Ϡ{�3i$8{�H�寢������z_�n��<��J�r�:��`�h��i���W^�yx,��J��uFw�"�3�u`��C�ɝ����t�.>���4�>�!�TV%�g�2�꿤z	�#kpVG~�����p;�o��MXx���m��j�uW�J�Ww�ﻹ)�ʃ����߿0;���|�޾�:����6�a%d�*Ь�]!��bީu�4���9�0���W���}�W�=a�]XdrP�NU3���0�Jݺ%x�)G��{���S
�4�{�f���v9 �t��'+�4_�T=s<��U�!ج��r`ӛ)�_���N<�cw{��7��7����^>�5�菐�~��x�҅c˒V�r��d+-��s;=�䤆���:)Y�z.$��l�$+�I{L���DS�����Ŭ�-��v��{����<��Z}b)�D�C��0-��誨[їG��݄��>7�Z�[R��3���z�0]���\��˫�b� ��d�iP�](���-��7:v�@�
u����c�9c���Z܂Q-�5��r���IZwW�?��%q:����.�X�J����+��ݮ���թ���o�9լ����S/�Q����p	]�qZ����aP�igXW��Sj̅��2����nNQ�[���a�t�U����w!m9��u�4��-0l�I��u�ݭ����k/؟�^�KD��ذ���-uZD�q{W�&U��p��|�A��&��m��4H_��|�5�ˀ�R.��e�8�s�+�2`������]{jV{u�?	�Z��Buh�F���o�|!��ܨC36�}�P�To��_%7��9�=��u�g��{��qV�{���5ҁC����x���]o��\*���Wx
���X�yq�Y��ӕ	�v�����9�K�����zo��8.�+��u~�C���7����E 5�u��F}�vL��%Pq�6']P��k�3D�c_=J�ΰ�0�#��������j��7�*�u��>�B���r����ETyD�������xr��'/)ֵԙ�u|���,��<��k~%�v����QL� x��mL�g2�{֖E╡Oe�ՠqLPn�rO�vT>�ϟj�t2�:c/jm�6�p�eM�b��ڴE`��p�]t�w6	q�gX@�@��͸n�fBJ�ߚ�GXN��M�Q�4=ȴ���=�,NzNT��bѶ���i9Y9�N�Z1��X���UGt|��S.�1g\%��W�]m�e\]u�39K[����=�vۗͱ�N���o=�㾕�^XCHwCI>	a���ئ��o�UV��
����Á�VU�Nvʵ�he��{�A-�֖_�'e����"�,��^��Z��-0C��w6�3w��v�ۼl��ll��W��xv|�]�ǃL���P� w�9ڍ^�O7����'֧֯�rъ��P��t��k�b��x&��<V�L��}�V�/�L�dK&�$�e��P�(Rn�2�^<��r�!�[�D�;�V'fET��*l��u��*j�?Q��Dg����>+��5�w�p_�At�W���g-����`r�E�߿]�`Ct?}�39���"�
'���o��f�
zp|⸊��_{�9��i_9C����CNܙ���JȆ:�t�	+�M�%�WS������l>噗2s���Ha�\Dr_4��2U�pܗb��%�R�M�%g��� ?Vh���[�\�^�����7��ІBãХ�ݮ�L���@�ƶ��r���F�O.�.�Ǚ���eu�U��˰��Z�c���!������Mޗ�v��Cz���7^n����(�����Y2O��S藜�tG��i�ۖ<E�4:�{ٖ��#"��ڽ0�����*�E��E�D�.��N�4����v�nN�YJ�t�ޙ����0e�0�Dn���G�N��!�Ut�0��=;��;�b�'۹a�>�ִ�ܗ��w�b��N�#^������)Ž���g��;��p�wΠF9�T���.uoԞ�FS�+p�e�]�g wv4��;�f
{&3�1�.�;��g���J�d�5|#�"�#u^]�Q����S!����=���nN����զ}뻍h�w���3��qy�	�u�%e�xa(Sp*�E��������l��^�o��p5��I����-��~�VF�{�c��[�ZT��V�L��<q�a�Ν��C]��R�dx�ƫky�>�dB��2'.���Vr��NV|u�4e^y�s�j�!�|"��K�Ɛ����o���z�u�|�|�x$�Q��钧��>��u	mx�~2����露IK��x"{�4��J���xha�ּ�]���S��J*�o�)b�W�+�^Ë.V������tE�zh�G��!9fK�ʪ�^u�q�}<�g�e���lt�I���C'vV��Su��&��ژn�:;;:���3�*�f� j,�(�yj��u1�U��3��n<���rv�.p�a���}��ru�FO��� ���P�M)��]-%2�KK6��Ĺ.��W�����.�'�gp缀�����G�>�/�W��-�"���������첷+8/JY^����f�A�M��L��;2�����IY�D�� �!��ίc_s�M���fz<��8�٦����',N�%��p2��rfl;]{�L.^ �{��8�JV�i�)B���d�|6m�>NȦ�ՍN��P���W�z�y��{!�S�&=��0%�9�W�hxJ�R�=���.^�.��Y��˙c{�E�b��<�N�z�Tt�ٮ}��°� s��HF�L�3��BȠ��X-=P��glm^&`q�;�W����n�
�f}�H��:���M����;�U0E��V�	�1o�<Ka����≗-�o����ᖠ۠�������%������s^}n?g�mN�NehV����|<j��a?Ow.�]gKy-_@m��uՆs�z�>�@r���a���t0I^+��_?F_W�3pE�Pі���VU�o�vB�݉��Y��\22���yzk�W�l�������4�����u���6ޮ�{Ǜ}n�ok�|���u��a5ݽ�p��w��m�}���	�%!t*=����p��[�
�to�׳{�o8ww�| �Q��"�4Αuǆ�����MUv�����a�^��kk���E��&=�u*͚5c
�}����'����?�Xz5-q�tH���P�x�/�
�RJJ�Z<�����֊�X�}].
�{r�*�>	
��^�)��V4*������Α�g-[�`�&���`K���4�ŝ>:G��J�.�w�?T�UP������η���s���0M۬�c��Y��X��mz��z�w�����tts������q�0����O�Z���	Y��ww΅��A�V�8k�L,�C�5�q|com��<��ttn������X-�Vl� �]˃��'��ڲ\�I���b���.�Q3�}Y�ؕ�7ĔԤ���*��oĮ({(�}����=÷�(q��JƠ���_nM篘�[U��஫؆��b��]$[�h��E�ۉ��;�G=U�(u��w"�s��:o~�`�x��[P���f	*���s��)��:A��7>0W/���W��\�N��<T�2��'�E�;&�d�����b��ֵX"\��@.��s*�[{�\"A�n�_(��P��:�9tGh=�H:�k��޼�ӱ��x���=|S:3�q\#�[���ʩ<�o1��gM�j��JࣟI����n�2{�$�\���yWX���ݼЕ$$yO�Hr\�gdV�n�ߞb�{�����>z6���e�p9�M�-�j�V3/I��x,�\�i5Fҁ�W+0��ɚ>zێ����)J�t#�{u�E@$3�I�'����uc+�X��\:�j�+i"�eRO��҈��	��Z�,F6�9�W�vDB{����n|��ó:|��o�}��֥�}�s$�cX*U�\����H��W�L��ӧU�Y4b�T6�o),R֜��EG��uWR��I��QG(���4V������n.�2w�+�uv��9q�*�{�rmGh�%��b��B}�kC��gb����մ\��a >�׀�uWR8g@4�r���d���>d�.6V�=��nge��y�@�f��8�9�D����X�z8��ӥ1�V����
�X�u�����>K�_>�_v��.�ݶV ,K����WFUw2lޚTYҍcf饖r����8�ZƈA�f��U�i��ҤhpZ�����7e�#�.��8ث;�=�����#�c�T�S)���q3���v�#�+l�K/p@-�'�C��"S`������U��aq��fVF+�i �:�Ro�OGJ:3o:�[���Qsldh�I��r�.���va����"p�+z����!}��њ�Ĳ^LG-�_=f�_9V�d����Գo��mn^��V���"���X���eMJ
$l Ti�S��N�rgJ5r�����׹;�_S��w�f�P�ұM޾�m�]3����!bm\���஝ں7���)�QV�r��������9X���<賻��ͮR����Κ�#y��:Ӌ��F�Vt'�$]Mm�/kk8}x�S�@��������n��.�*V���}�]�J��[Ʊ��Ć�w��WK���nU�x\��F�e���Q��t�ƴJ�gbY�7i��S��z���RsڴOp2���|��M�&K�:M\q]V�l%��w�N.�����R�62�;y��cx��qfu��:���p��o�e���+;q��u�S��l+I��f#�m��oT�VTS)��k1	}�B�r�Y��V�fR[�K`,v*�U��>�21�V���;�Vn�<��pe3π�ګ���`&t�z�gq��y�	x�J�x�;"�r�����#��8!��g�t0:�����)��(�.�t�X�W�K?��\@���e�9:���o��K�,>U���9�73H�R�TV0����"�1��E�ZZ~������,��ʊ�Z"җ2�ZK�k
Z�*�[� ��DlKK��b�[m��*%aR�UEQeh��)j�Q��U�DT[h��EX�Bڈ�F�d֩`�KJV��jU ��Ub��6�k
*�5*[(���l��������ڢ*�ڋ���h�S2�q�EBڨ���%��3-km6�Lj�UT������֪V����*�T\�(��K@FZQE`�+n!�TL@mR1n\ƉmZ�+-�Tj����
��j�*+*��#Z�J��
���h�L���TYmc�JE�Q�̐X�ڱX��Z�EQZ*QmAX%)PR��R��kaQD���#�VڙjµE�*�(�ED�Vڶ�b���
�"�Q�U�Ib�*�iFV�PcU1-���
�b�Db �T"(,V҂��V��"���`��TFT��*Vڪ����Xe(��bTPT��TF[U`��#
P�(�G]������s/w�7�-�	F�J�&��--������f�c�mC:�.|�.�V�8oE�۾}��Y�/�����|>�GIn�7�������3�*~`zx����]J�^�Z�G�kl�r���=��^�����Y�5�3d>���T��*�q�3�V��Jԫ�a�P|�2b܁2�/7����y��j���sV�Xg���TC��7�J�M	�
M>u�߲M�n�}(�]�	J8�<1a����ۦu/y�=a��~CAy-õQ�CA�\�Wi��'�wx����XHՏWKD���Z��Z7���2k����M62�kxo���y��~����f��ߺo��^XC�1T������b�.@{e[�9؆)���R'�w���\'5�x�3h6�}R�S~�xt�Xx���,����"�"�XU�����K�,�މ�9ƚ��� ʣ��K&���B���m����]��~i�Rs*�2�˞*5R�~�4b9��6-����|r�L2��B�]���7����x֕�ܫ��+����q�B�v�ĸ�P�(���������zP��LzQ"�w`�����#9+9�e^M��/*߭��Y�I����/7�niv��s��2ӘxV/��E�ӣ��������%>S�n����Ky���Yoh����C*tctZ����ﻤJl�s(U��+e\���l�x9=;]V۵b�띀榡���着�����DĬ�.?��Q"�Ҭ�X�<�������He�t�����\�	*�]37�sl��z�
��1���Qf� �OQOQ6�L���m����M� �rի���׾����-�S�;a��~�+"��R+JFh�/hWS�:�=�o�S��ӣ�Xc�m�!�
yB,s��M���2U�p����§ܔ�R��rܨº���LK�>��x�.��}�J֣�.�����̵�.$o�%BM������JC��$|r	*dpF1r��b�
����'��Me+ߐ7]�߉��h�`"�nɃ�m����ڡ�w�z��I�%+�U���Qҿ����߳�a{N�,���Y�wQ�5+&�. �;[�>��j��^Vw�>q�ҎN۪B�3][�������2���n_N����}���bV������̼�z4����f�;���u�o�7Pm���wā�����$�����u��R��]cLʪ��wzk���t�ؗ�-��D�
�
n�����iȥ��BRz��)H��>�UA��4^ƔS��`�b����k��X5�t���R�[e����71_[�bSCm�k�&�E�wh��;#5��3v��U�>]�;f:Ż���VZ2�.Sŗ���UЬm�e��}(97�55��_U}��2�����ܻ�e�:�z��$��~�k�هeU���ݯ�3�]o�<��U �;՜��|��+gB^"
C�� =�ME����ȅ{��"���ϫ<�쎲6nǖ�݅�׬9V����*�H�Wn��ڧ���Zupv~�Y�Ȧ�0��]�R�,y �S�R7ZϢ���Ip�0�a�>iw��}�U�~�~E�{a� =�V�����VH�T��\�][�A������Jm`��,�S&�f-J��qs���5�׃/�ʮj�^�%����8/Ze��Q�
��_'��웅�C=;7�<��/��x�p�ͱ�;���rߓ���t�r��S�p�p��򒱍yห�9���]���8�i�ꤳ5z��*�(?u	˓��o�Pք�,�U�o֧�VTpr	���a9h$�ކ����Y�[GG��B�"�K*�RwИw�.P���U���q�>����9��CI��閳�m��(R�=�����˵�%g�N�ج�dVun^�l�F�$���O�Wj�/�ֆ��]f�}ŋ��.��
[5�11Aon�	�<So{s�6�e1}4�⻘f��Ql^����LM��y�ξ/&ͫ�΍�E_p��Z䁎�P��Ú�qO�]�ocڻ��I�O��I������{�N�����d��#V}u���}.��@hY�yn-�τ�����:ԃ��ז�﻽���L�5�g��*��ά8�q��+ ��ULdv��P�t&��{�C�w��w�A�:�Խ����g�ʩ����K��~��X���n3[��E�?n��b^>��wCJ���A�_%����OXsZu�|5��%��u��3f�?	�r�3�ָ!��� t�VG�pO]m��t�`j`�~AW�g��궄;�88.�~��b����q�y��j���ְ��@��+O��:%>@V�_J�9�'��B�o#w99ek���Κ<7�z��ޑ�D���*^XSIYt&ςB�4�����XЭ�*�ҝq�F�h��u�G��+�y}rWl�|�u����H�rTIYt8�A�T�7���;��a�4��W��A�G�y�a�׵�s,pKk�mF-��o���t�be.#y6����O��Xw6��]{�Z�B��,ﺜ]�,Ld�D:��ϻ�a>�?O������o����2�k]7���V���k�V�m�f!�*w(~�Ks�-&~���Afe�B��'�^��9F�kV5�q��:��dOpBX�;��Y�.M��lӺ뷻�`���L��j���(���;�qc�,&i��~����� ����U޵��3���ݰl�+-ϫ>�ZE��wܵ�i�\���6d�Aq���q�.�`I�7�=q��+�a���Æ��P��׎��6���e�8�|\t�vǇ8�|�0��4�z��8׼�� �"GtU@����>�3/}h��r����ȑ��=+�7Y�+T`���O~2���X��J�CF���2���u0�H�2Q̖Bۇ_����1O%n!\3��{Bk�r�6#���=<w���.��a���r����ֳD4u�g�BIz~��7 �_���r�j�bǽ3��vL�� ��@�Q��yY+hLf�0�����YWL樥3b�_��#�]�q�J:������=��9�yh ��E���ou�{�^�!Ou���J���?�r�G�&��d�:�>�V5�8Q�Tqb�u�I��Z��:xe��ד��a#V=U%�W���+����Jy�y��wX�b�і�=$�qV�S�ν���fg.� ��氆ҕ�^L�!���`K�w�]��&v�*��� y5gFm�e/v"�G�����1y��q��gM�W�L���1�h���
4��\�s�I�2T¤�f��q��o+-�M�^.������;�tT��d�qp�@��R).�dxt�vr���2�V�'F�d���������~��n���������D�H���=D����6��`�R)*��S����c}n���-2��]5��%;�{��W[�e�3�K6�p��k�$+�a���g����3�O>n�?-ML^�
��3�fR� @^!�+�Q��O5cT6o9�hV}����q�bx�o��V�<�_5�.pǂ��;-).��&�E Dn��Wt�Ň�w���T��,�g���T��y.�o��To1��y"2K}�UĂ��>�NNbM�-Ё�����'u�w�����;7��
��1��p��b ��OW�=D�^�E�Aѧ�1�GP�~��'���7/�����_-��;a��~ϔ��5b��IX��h�%⌴���f��L�����[�P#޺ćE�L����*h2���J����B0:��X:��7R<��/(�z,Vy���-e��й|o.�;{�!��v;�̵��č�$�I��j���QZ���Bݥt�OD����;�[y��<
�7���Ue����s��H���Lk�5;�3yoqP�첉R�R��gt@�I^�A!EJ�&@mnP�r�� �u���@vD�}��b�'A��Y}�lu:_'4w�w5���Mc����7�2��Zdl&���{k���ҭ�]!�j�.�*wZ�9��C�/C�i�;��L�3�}�� 1���m{���.���Et��_���Zi���L���=�MC��3Z�VI��Pv���cW�F����;n�}-�f-��B2�	g_�s�O���"��{�
��YT0��	ҶuY�<�a�������>�������]�^��u�x���w�#U����$O��<b<������O}�_���{޺D��-����x�e���׏�YW��.5bׁ������9��m;�aߥU��:?o٭ߙ\s�����D�"%½H���`�+�qX�v��ȅ_;�E���{Օ�^4�S3���1B=���Yɕ
*�u��\_���7K�`?�0�ȳ+�yO�O���ͼa���I]�ߏ}����ߗ��@PY�*�{���� ��v�E�0�1��s�ӌ?!��|�'�{�i�C�2�>J¦�f'�̘�ľoI4�3L�1"���|0�H����c�/O~�/¶��=�5�z��_ԅg+��d�svOY_S���6���$�y�h+����~�0Yԩ�w�+ɶϓ��Lk"�'Y���"�q�%@�SFXu�g9d�|g�7�Ͻ�q޽�����|�;4�I�����m
�tguǬ���R,�~�~LN2z�=O��Ch+�&��4x��Ri
���Rm1�����#&=LI�;��VF�!�E+#�J h�w��Zh�^Z�f,_�y*������蒀�S�lӧ�j��i�j9ot[lˬ��Q�������"#O8t�i�J��{7�~���my�Lnr~�ٖ�(��:c]��.���K)�����أ��f�#��TVj��}��Dq�*+�o��Y�/��<}�� �
�=�+;w�{C�Ak?����
ɳUL@�+8����)6� �s�u&�Xz�0�Xc�=I�YP�{�@����.��7:����;�I�ް*F�����x���Ӟss��iA�m���R)�=}t��Y+�j���m �a�P��O�Hu����X�2���?!SI�w��6ŝa�c'�9�OX|�3�?^�D�!��/�b�����ö9�[�$Nwٯ��ϻ[�w��a�|�Ɉ�_�m
��݁�GXM!�)���ɤ�=f�8������@�=�'�Wÿ��q�qS�1�AOO���4���߳L��0�u1<��|�yLٕA��gN�_��� 8��Ą@�:KA���I{�1�J�S��w�?2���b}�M&�i
�*{l�B�z���'�H)��8�N�~q���&�8����ө��I�y��럍=����<ֿmﮙ?&;`W��bDd��b�p�gYd�9��H. {�}�k��Z��I��)�Vvͦ�4��O��l�)6� �g�1����2W��&=e|�G���������������<JͰ��Mn�1ԯ��d�����Y�4����;�h)�M<�3Ă��_N�?SĂ�w�M���i4�乑|`T|�J� x�#�H�j�S��V'�g�������]�����>La�`�0�f3���H/�:�z{��I%fϿ���Y1����M�RW��'��}��6�AH��2�R,�9ߵ��)
�3�y��L�'��O~��s��o�dt����I���������}\*���Pr�n0Y�+&2��&0�x��R�E*g��z���<�xi�A�%@�kF2u���ɟ����N�^'�߷��!Rw�{�����O����ߥ�ù����|a��6@$�{�Z�S=q�gp��h���%��i��Rs��i�ɴ��wH)��ɉ��gAgS�<�xu�'����3Hq:�O�ϼ�c�f���׿�} ʧG��DG�G�}�C�R~J���ǌ�����s�!��bL~N�EĬ�3VzɈ�xi�d�_��nÈi+%W�l�I��u��*K����G����R�>��l�k.|)�3zG϶=�Ю=�Ю����]*s�Jf�F�K=��>��,�q���ïnEy�:�d�v���Z2i�-S���H]��˘-A��D��K���ʽ�Q��¨B�ѵ;��q9Lɝ8Duw���|>^J��*�a�����B��]?���6���?w}�6�`Tx�jT?!�bCÝ֧P�Y��'�<�4�!��ݼCI����i*E�w���i:�Ɍ�nÉ�#�d_���Ɋ�u���e����;Y��bO��(t��큈)g�ì*o��f��J���Y>9��6���8���涓�+�G�V5�ϒ��l1�a��1�Ă�ȥ�`<C aa���Ǹk��?\���}_����Jú�I�OYYϬ?yM�i*N!]���L�M�Y��Lk�'��SϨbJ�d�3�k�%@�Wú�Rz�=`T?w�*}d�ǉ<��� ��m�?��S���/� ��#iٖ|M��h|�'9C<�� u��ɼi���f���6�O��߲xΤ��'���Ă�z���jm"��Y��_�(~���+���lo�����f��>=g3/?{t��R�U}�AH�Ʌ���ʆ����i����~a��4��Ԛ0*�9��>C��O��M3��:��W��c�e��(���,_��זݾ����|����g�q �a�s�ĩ��XV1�&>��ISHT��l�IP�)��^~�1���=a��i
��& |��������~�?#�@F��}��]�_�{��~`�k�Aa�X,�*vg����xw�ju<H/���wZ6����ֿ$Y�RVn�!��Leg9g���*T���1�VE&!]�_�̞:@���|H��@���,{����7Ϳf��1��d����������9�CO̘�����i"2w�f&�6���'穉ǜ�I��'wCxsy;@ӈ)�R�bTR�̜#��$}d#�wM?����������4ퟒc��y�R�?!����T��]��2o�6Ɉy>��gY3.�s�i'P�Y=������)׽�D��Ăʞw!��N�d�ɧO�#g���FzWOe��n�o{��-^�$��
�k8ʇ�<La��c>B�gXl��H/~C-4�Ă�7=�'P�<J�I�����
§]�ĨT��y�n�*���|��R@|�&�����6��*�Ӻx-c��ϣ�S��ڔ��]EV}����z�v�a�y����!�Fb�)is{���{S��{��)|k� vй�z���xvd����Z�%���D]p��p�G;f!�s`��6�o,����We����^1�����| z7��/5�n������~��g�J���R������>��>v��+�O����g���1�0�c7?Sl�6�^!�}�I�u=C<>�=H�����N��m6��Vo�{�����y���u֓�����`/B����]��R���ۺ"������2x��w&�(*|���3�%d٫�������q'�����}=�i"0��:��G������}�>"��h���c�������ǻ@Ӥ��C��2M;@�)�{���@�����S��M%|;܁��bL}c�|����=�4�ʑ@�]3�K�=d���'L�&e���ĜB�a�}�a����{�{���}���3�+����kG�x� �utɧ���M0{a]�+�'{�t~C�����i����=Lg�̑g�+q�-=M$�'��f���_�7��M�H��z�9��Ƴ�_�����l��PG���#�@a�V���v�ĕ
��s$_�`b�扦u�S;d��6�P<OL��R~e~`T��g��m
��<��
�9y�H,��<�~���7�u��w�}�˯�a�1=H/���bi��bO&�c�E��?& bVN����ܲm�C�ÈmĬ�L��H/2|s_k������R~|g̕�㙓�_Y4��'=�]�S{�o���<�����{=I�
�&'K��PR#5hx���Y�nn�5d��b��;@�9�����Hq���B�i*M�N&����M<���Ak:��w��� �g����Z�����J������{~Cȏ����}̩�~d�g�<�r�q+1�2���I>B�f�W�Ab�:��$�ɦM?2}�i���c��!�W������O�M ���z����:��Y��?o�ڽ&��p��?"?:y��C�� �a�{���xΡ��q���ĩ�;�)��N<|2�H%B�V�y큉+7n �_�`b(�Y�&{a�g���3?t~��~����M��pf���"�����|~t˄��8��+�w�M ����֧R�c�~���bA�ڑM��������R,�=��@�Y>M�9�Ɉ*l����Y��U����˥�i/�P�N�p�:�ӥR�1����9JP�]M����BN�
"�Wi�Z��g8�O.�˦2xRgs�ėS;suVp�,��|e)j�X.��]m�o�gƧ�/�w[b�㱡(���uAڎgK�'.�vg]k|6����L���*�a�D�x�"�wܔi�
�]smh�Co�Tm)�*��V3�t
K;��6�]�ٯ�c݌����U�M�]�)�q�L�������H�g>O�N������˙�>.`�tS9'2��,-Y��WXֳ
�V�
k�d���s62�&��%��̵Y���,^T-I2�RԼj�K�P;�Q0��u�5���<u��n��|D+�`�����fffD��a���:�q�� �+q&C	��nU�c��v��I֕�f�$g��Fj�Ư����Un!ћ@;�%p��ή�S4���>7�8�+0v��}B�Ł��ܺ�R�641u�`SC+U)�Ϸ)Q�öBǳ9���5Zi��n��p*���2<�vF�ɹ��ur��7�b����jNO���/7��J��}��e���YDVCVb{Cw��凲����r<�V�R�a�7f��`��Y��M�C(:���i�?n��a a����\�Z2���Yd���L�ۺu�V�+��s�	�K,w8�|lp֭��
#�l�K�.|�l}�'ҝM��zdgi����L���9<߭�ɣ;���h���k��*��ow*E)�X�d\ ������붂��ٽ��7Q*�Q$7g%ki�v�K-f�zm�0� ���{X;���^'�H�>����� ���	ï�C(IW�r��SyEc�pB�5��"��K�a�*�N�H%K+\�m�r�y�j�ܷ%��e�a��!6��L�x��&���s�^�I�8�ږ�.֩�y#3;Aٴ�l:��]c2�'2�ꙌT����K�@��Ĺ+1"����y�3̅�i�Y�ǉ9�7]�]� _%��靳����R�)����Ok����%�cz�����s��a��;�O��O5�`��u�YT��MY��+��Q���VL��im���C=\���̫U3���|���=,�vӂ�<m�J�'hk��9V�bⶐ��&��`�����·O	�_V%�wnvCo1ܥ�:�ob�{�I�o�ճ�l��Ho&kcjZYˊȤ�Su<���]30v�%��/��EیO	Q:ܨz�J�e���Ŷ�L�
�C�ꣳ:u:+w6!9XG^ut���h��+y�jkR�M�nL�֯o����*%l��՞HH2Vp��+st���[ub��G�V�k{��
��IV�q�GDB�_�u*��&Z������ֱR`�m*h��r��y�N�� �W.�QuL��;��cY\2��L嘷��Z���y��+�9r�B�w�n���;Wҝap��)�+.���ik���s�u�Ζ�.��9�'�wf�u�������;�~�O��1eJ�RR�
���Ar�m���TZт�F1E+D
Ũ�AJ�KV�V���V��R���E�,QUj�9B�h��(��@E���Q�
��D-��QAEQDc�IPb* �(�b�ȤX�5�TX�,�(���Ad��iX�T��U`�QEDUPY�V(kYV�F *�,�����+\KDPb��l�TQ�VՊ,R,R
 4��QX,bV�9Je�J�V¢�R
�)��kZ�+��V
(,+*�����1`�[)
E1D�,X��D���� *V��D\�Q��RX��(*"
-C2�Hřm�,[E
6�F(�E`�Q1*,U1A���(1ŌQ��E--���9j"�3�[-(-����X���"�iAb�[J�Vc�8ʨ"�aET��T���6��@\j�Fk�����7���ǹ7{�������iV_;�il��;�Qr��@�7��j" � ��5�Ls�v�zw��9�}� �����k���,��>8~��PR(�S�ގ�|�>d���a?&ߙ:��ê���ɹ���Ǭ
���gsRx�1 �Ú�R;�i�bO�O��N���4�Z���w��vC��{7��޼S�#�@B Q&3��$�7E1 ���7����!���Rc�T�>�Sl���C��M�~Jβw4�0*M�S�{�I�z��/�5��x��� k�O]���u��߻�O�3ۮ��̕�'��V����v��|�C�+���|ʇ�?n�H,����:¦��l��=C�x͡�</�����Xo�� u+
¦���M�~J�7�����߽�m��̾��ϬI_?Y���X���
E�é�Y�Lf�+{g��=e}d�n�I�uĞ�_=��4���Y��1�%H,�7=���<f�}�i�"����=�����w3/���c��Dp��������l�@�Y6�ڛf�Y1�C��'�+�Y��6����{hz�"ɣ/SI�'������&�̝L~O��M$��Y�ӶA@�c� �ݳ���}��]���0�"���dwd��y�rM> qě�;͆$�k��AO�TJ�w��m�M0�7/p<LH.3�,���c��&=eH����i�2\;�ۜ��Jb�G!/�U��oz�����a�Ĭ�?Y��0*N!|��m�j�`Vx{�i"�I��L?w솙�J��~N�͟���_�5S��I]���I�VT=M��&�1
F�����(��0����������������g�bI_�>C�����aXjk��bR���ᴛ~偌?Ms6��R/��s��
E�a�g�ݐ�?2Vx~�C���&�_G՟y��+� �}��-�a�����~�޳\8�PX~k�(c8� ��yC�Vg��6n�=dR�����H/,��^RT
��߲u�gݲc'�s6�I�+Ԭ���i
�_�����|@$|O�/�A�ʷId�	��}�]�O���q�0���@�+��L�3�$��'�l4�~`Tި`������8��'�ɏ�t���>�$��,�PS�T{>�m�Y��Nk\��O3g�k7�[��%�|{��SMu�WS���}��6�^<І�f�[��Cs��wJ C(�Td��X;�Y�'��R���;r��%��Y/��	;AՕ�d=r���sy���r#��O����<35�=n;�0�;/�����>����1���,����d|	���ާc�>?@�Nv�z�Rc�T��`J�d�N��d��Y�x[j���8�LLd����2�S�8��E�������4��:@�+^���2��ѽߎv{�_}�M�o<|a��iRW}=֠(,����M�u�f�~a�cÞ�a�f3�1<�p=a�bbWfXb�XTճ��L@�_�i&�r��y7f��
E��7�}�.au}�����s{�|��R,���R�d���H�7d���?��m%gI���0*����J�^���a�6��b���Y�q8�bAx�O���J�R��߼ם����:�g?�~�����(>�/��D}�ZI��*�m
�tg���'���?����'�3��w��T���<�4x��Ri
��$�c�g��i"2c�ě�wL���q�{��u��S?��Y���R���W�U����hm ��-��H)��f���Ĭ�z�������_aԞ?0�a�9����$Ǭ�~� ~J�̗|d�IY���<���Ro߽�Y�Hĩ���u�o�B?|�0���݆�R)�>z��,ed��P��At��P��'ɤ:���M`T|ʚ򟐩���;=�&س�>Ld����f3�r�z ��qO}��5t䙷��ԹD�ԅ|UxQVk�i<xɈ�0�%y���1"��:[&�R,����M{HVi�& |���W�d$�:���c�
���{��li+3�yn_7���v�����8���?3��(�(��Q��ȥC��CI�'s���ԕ���I�+;�&'ڤ�i&��R�-��HT���������8�N�~q�~��i�_X}���f���>;���ݺ�܂���">���t�0���N��wܚH��t���;��:��&��ki��y��I�hbAk�5�~j
b���OhJΧ��٤�H#�z��<C��{�Y}�9��u��>��?]{����=I���}���g��5f�1��~Ì�y~`V~��'P�VJ��w� �S�4���_�+%w;�jL�O�y�a6��I��g�̋������w�������޽͖�+�Z��*�15s��GAլ�}��+��TŰ��Cd�W�ļ���*ߛP#|gm���̷�t���S�;;U	e6k��سhZ��muA
�sSnn7׽��6AYW�nJ<2�`�곝�z�6=>]{ʏ9���?~�>��k�ߐ��$��Ş��1���!��~v~�i��͞��E�Y��4�I��&0���M�RW��?w�<I�*
E�����x��g;̇���B�L��{æ��{��y���s�^ow��&e��t��i��Rc8���P����Y0Y�VM�Y���c?>MU �dR�S��H/���m�������V{�&~w@m6��W�������=��W��r��m{��>�"v{�O��&� ���p��S=q�3�|ɴJ�b����
���4�d�c���R#'_�g�3�������Ă�M{�:���P�|6ر�ҿ!޻��J?�٤���!S��iP>J�S��Ch%@���4��l=C?s��i���'��(%g�P�g������4βo/�
��!���_��ԚAH�����O5~�?{�T�Ϳ�6G���N��W�'9M$O���zé�����0*<�sR���NwZ�B�f�z��s�Ob�M��$�"���"�Ŀ�d4���Y��?S�G/�à��}��?O�5{_�8�!RW[�����i
���^�����ϰ�
��!Y����q9�M�jm��Rq��g5���^0*~��X~k�%a���i�a��17l"�����k�Q�.��q�����'�i �O��c4��%a��4�d����X~<��4�'�W�)��M!Y�ϲM5����~�H*q�yϵ����q+��k�I�x��P�w�*x��F�������z��P;^�}�HV~�W�AH��>=ˤ��26�2����Aq����N��2i��8��B��i���z�0��X{��<gRc�S����Ak=I��?K�����W��f�WZ�;_������=������
�g�����t��R�Uy�̀��S��hq�� ���f>�}�i��n�X����y��I�����a�m��1��5���U�~V�X�H����=�������c��析����c?{��!���Mw���T���4V�Lxɏ;d��T��l��i%B��Z�� ��2�=a��i
��& |���,��8��>i	�o�~o�{�����#�2�<ϲ��k�1���t�bx12�;@\�9���a��a��]}|]��1��֯j!��ؖ����;;7kiV�C�X���Wv�k��ҍQ*��)�kÆ��v**w�o4�ue��bt���h�rw�}F������k�}��������CW����x�|`/����g��;�i�0�c!����� ��~5�h���bA�wZ��f��J��̆�1���Z@�Rz����+"���_ K>?}�����������_���O�>J�C����1��z�wX��u1����P��&&=c�LH#'�y��6�Y�'����'�S��o$������9�t��q=��" !_��nt��~��mO��� !3+�x�t�0*A~g�6~�ߘ�]Ͼ��M�f�1�%gY3.�}���N�R�o�ޗ ���%>$T�����wt�"Bk�������sp6�oWTX_��!�X��̚BT<d�d�Ԟ�7��0��3l�����8�i&�a�"��I6r��"�s�}�"���뫝�_�ԛ�l���u>�g}_ ��T��~�_6~a���6�m��*S�O�a�4���75zϝ��
��L���g�O�C��3�i�M$�~ϲi1��b�{���YP�Jߵ���}�^뿼�9�9���N�z�����ܕ�!��邌�Ή���t-Xt���ۯ�᤯|��貸��=����K^��.ك��J%�;Q�C��XH����U��hq>��u�_p�QL�`�)�IwYK�`O]p�2�[_<��-<'G<���-}ƴWR5��h�Gڥ�V��ŽOg!�t��V��k�&���R(��ϔ姎o��h�`Wy)Mfiñ��{y"�ϊ�[���j��0�����t�^�a�kep�\��:ͧ�(�G|�q�kwT'K�����Vh�p��)��ï�/�9;;˥�p� �~��+��4q�����ݾ�l���8��pݗ�tV#ʆ�gl�J���&�g��wJ���ͥq�]{�Q��I�(�ʬZ����W5�hY�&ѹHr���->������u실V�՗K����f���BX��e����b��Pٰ3�7���#|\}�7Ͻ"����դI�ZWe2�I�W�n�$Ծ��y}ރR@����G!��-o������O:$P�݂�븜�^H� �[����S� ��h?s^�GY����OE��α�z�Al�H^J�)^�hx9��,�D'�➢j�݊��֭���At��bB�ѯ,�����.:�觊v�̇�JȆ|`�k r���3�u����F��,�+ռ����ԃ=���/���3%YG�%؄:�5au������\��}�4��VK�v�>j�[�ܰȿ��{ٖ�=��	>�Ҡ�_y��>�gxDl#:g���y�ρc;�k�pJ�Ua�f
���LG��Tz�v:h���z��(H���Qϥ(��'o���+ڴ��{���-��\Llt9���s�v�z��7�'��=�Y��cW�F���(�Ӷꕃ1�n���B'�_������qε�;L�ގ�D�忓�7v�:�)1瞼�[J��\�٘����ל�����9��^j'�[դi�(�5���u�0������Đ���
�c3��zhrP�#8[%w%�:e�K,97{�=�X��G<ܔ�y�~�������Kҽ�`X�����������Ɯ�P�*r�.o`�>���f�G`�_�u�lJɲr��2<�󆕲;P�.]ŀZ�#z�42��8:��������'L��v��*�כYV���}Ҹ- ��V�G����=^�pY�W�t��I�U���R��Z���xvf�^��3⯫�O�m`���ig��:�ο�9�v��w��.�)����/S�W== ���>�-�f{�։��EZ6w�s�x�����m�l���{9������`.�9��w���	�Sw��Ì��4��s^����R��l�$C��|�B�ς�kn<�N����U�B��6�?M�+�#�Y�=Fy/;�Wx]���x~�!�wEs��c-�����'�n�r����[쓯38���,y��0hM��d�hr7E�ʏ�;SQ�tbc�e�ߞ�9d����X�)���As>��m�4�S<���)�>��#���KzJA�"�X���H�
`pf�=�� Jm2h.T�����ms����Re��\ŋ�mhV��եn�.{S����p�V�"-���l� ��|�o������	{��?}��UUzd�k0�v�w�޵��lfįuRo 5�/ʂ�{+�t�tNV7K�j�s�/|\����|�d���M�uR������
sr���|�Vo.ۇd����o����%[�P��;��Ҩt�8$5*��M��=�2�py�sܽ�{u��9z��.m��uӸ��zKԕ8r�,�=ǝ��i��g`:S&�L;�<6�c3r�����s{<�JKw݄��}v����S��f&�hZ7f_�e�77��.d�E�Q_��n�<Y1w��%�o9����[�x��/�X;�b��bu�a};�eX�Lg����7����bܩyˤ���{<�w���0����h��׏{xv��^�;�J��H����>��cOyɵ��v|W9��j�����똯R�O���ƧY��g2�6��}�/_�*H�i����|^��ה®��)����Qw��f62���˦�Vn�D�OE��eo�Q+�y:�c[6�JÚ�b��g3�Nr�ޭ�������߮vŎ�RA8�V4�jK������o��lΣ*v��I%�[3PW��1�,v*���b���cMf���O�{������~� ��/~���Z!�*�Ϸ�y�]���I�1�軙��E��o���.���X��>�1�y��%��N�����<��G�E�}�2���v�o��O�&H{��i�����J�����Rc79�{`�qZ���`M�$�8=9Er4��yN��0�L��V�?X��7�N3��9sqJɀ5�Qh����5��䚢��K�ӨG�g��S����_9�`2
�G�$Y�u����J<Db�Kf:͍�����qP\��M��]�u����r
��_zx�Wt���|�ךO�@��}i���e˥��W:��o؟�W�|��O�fLӚ]����:�~m{��Oq����摬�k~R_�y��wnߨ�YuĲ�2R�u}OA�<�Չ�(H�VN'(�=`�O'`�6�Sw���Ǣ�z�n������ʄfξ�hW�J^�oN�Pu��ǯ��_�gʶN�wM	���]{�ڷ|>������:b��)k�p�|z�;S�{è\ǳ������U�e`�s�����g�%�_m_aɖ"P�dQ�9;��,|�d�f7������y읲GU�k3���Κ'Tx'�_�{���CpD=�5��B̬�gk����M�̵�K�٢d��烪��.s��6?W��`f.ZH9'f�1j���J�	�5��=��:rL�,zv�o��g��d�<nFe�V����t�&�ڥ�+��Z�m����7��]=]��{�ѾW� ��\BD���{�g_
�'1�Ož�*�O]�t�7$/dC��0}EѪb�N��1ݏ3�b��ՒS���1����{��o��m}s�\�s>�:e������|߽�s�ݬ�y�4<�;�Ra;�Md܃�J�\��{�*(��x)c'�Y��73\���3_�̿e?|��;'׆P};�����r��6�&�6�k�ޫ�O;}�oWz D�\��*�}�V9�3>3$h�����L�����֮ʋچ
�Ĳ��]8 ��f�=r�4�'�΃3���x�fq���K�z<	��^�5� �)�h�t's3��qe���Ֆ�Ef��ұ��_�D�X2e�->���d���&��mg������yItK)\6�� ����֔3��}�}U]��s�1n�iο����Q[C����7ܷ��쯣{�Nw�-�NgL�""�y�4��ԭl�:Y�s�Ӽ1����t��y!��绅�~�g�^����R�hrB6+�ܰNķ�Nρ��)���.Y����ag�qE��N`o�r�x�J���y�W6�_�1Q�Ղv�_l��ww&77�C�"���v���[g�{)b�w}���9�Gr������9�OJ�����vmo��2'��_�,;�r�����y�Odd��\~�,���9��7�y)$VP�w��*��U�G��~��N8�\�,ڔ��b>ݹ��>�]��X���g+^�h������}M���b��;v��|ߥ7�U���)���W,r�{�ڌL��w�
�b�rQ��	��/J�Xoo/���u�Ω�{ג)��Ӎ�k��?=rBe���V�)��I�`ڄ�Y��%����5(d,'���L��y[ǃn��4#�w����;J{ZN�i��|�����/�E�D[ՋFcaQۧ��U]#(�n��\֝�D�]�j<:���:�Co��;�-vp|*!Y�xi�4��[n9͝E�E.X�D�+u
�ŝ�Y�Y�"!���ͳ�9-8->�k:	�Ll��^n�}�ևǢ�Q\^�5uøЃ�'28J-�c�3���:@�w���Ԏ�4c(<�A�X;fZ�ӌ�՛�a�1�2��B!�=/W�f`Gu�mwQ�I�C]wVQë��h�G8'��a��cdK��\�ӳ&tDT�w.���W�Ʉ��@[����������u�y��)u^C+c)КN��=�mV��T��5z�S�t��6�sC�*W�敍 U4:�՚N�Y�`�D���	�72eiK��V�n�v|�ܭ5����KE�}\Ԝ�����]7Z�i���M�>�V���w�΂���S-�Jʋ�4)*�0U���X�
0�Y���X�\��Y�2aV��Wge�����W\�_:wL
k�n+�&��ά��$06�l�n�ͮ���=k�x:��Q��	���\y]�m�ۅlc���o���#V����8���NY6jF�P���K�PS��U=)�s���� �]#W7k,���`�(�4]�[���������Ӱ�tJѲe�@�`�xo�*���h�����)]u46JG��[��^e`��)X¢��l�Ž,L�î�+.,Qp�;�IWSGOu=A^<�A�+a�η�zP�5
c�V�Ym>Feg?�W] ���^Ix�����Z��1a��*,�&�cZن���W]����7խ	V;������-t��q-ݒ�8T�p�B\Q��n�3O�h<� Տ=��+ ��À7�,�.��S[�!ݮAd��:��J�h�q��e��6 ���β�u,�{�C��82�It�4Q�hu
��Aґ����_
��،S4^^K�c���Mr��t�6Jj�q�JJ���H4��*3��f����f����i�=�o>�WL��H���P�� %_������S�V�t�r[�J��qk��<�&��b�	�'iT�e_��;���j���};\W����WuͶب<���3b짥&aBn�8Ք�͙͡�Q���4�y�����p���A�|�9���-
Ȉb���K�������wgb�<
6z�����мE�����1�p������l8.�q�o ���d9;��Dr��&VI���/p�n�
�p�#�C,fr�
}�w���V������į��(S�XL��ֆ5u�8�˫�pM������weÚ���BoMtЗ�	O���C�4 ���Z��W����X0��t�k���'և`������~uu���j�QPe�TelEAUb���Q�e1��j(���UAA`��m�0X�+R(��m%ciX��DF
"ԪĹL,��p�J�U�)R�j[E���%�m
*�R(,X�H�V+0�V#b5��UA`,1U���Q��
(�QX�%�����jʈ���"�*[h,�A��
��P�Em*""UFe�������LlA-Qb�YdUPTV*�V��b�6��Ic"*cE�
4H�Z�FEb�EL�����R�X�[T���,b���(���TD�
Z("ZX�
ъ��̸(�q��X�B��Tb�
��Q%�9Ȏ\�R���-EamW3�1Ee��UQER�A\�&�VDTX,X�",e`�1ATD1��"&Z�0�L��m*�ؘ��PX��V��I���d�b�Db�YUX��H��@QD�H�***�mUc��TQ��b��{����k~�̓�}շr��s����y���Uƃ�c&K�7�S}쬦��0��^'XX`���S�Ӫ�ކ�9�UU}_WL�Fw$a�#Z���y����]u�sg$y";��<�5��0ھn�S�|2����	�:%Y��I|�[���s��=l4�ng�$}ێH��o��Y��}��C�3~�(s���ӻ�G�n����'w��ݯ[�ΐi�e��)�Ȱ'a�Rg�r/ʾ\�0X�Y���zCЫW�q���\�:�b�l���_�Z˒�g�`�}T��_����c��(emGy=��qN��Ǆ9��t>2�\�`�:l�IN�<���Fni��讈�=S���|�Z��ԓsGk��m�w��tҫ�)�:��5��7u�!��O)�V7�G��{[V�{��;�J�N���mb�X�[�_�Ʒvv>���bid;�X;��&�vR�A����~������LW�;V804<��$�W6���C�1��t��T���5�>�v�^\�;�����#�=r���Y��#L�"ٰ���B�݇����;����P��4���_
�Pc\��!���[���?Z�~���%�!+]\���u�T|��He3Ee�΢(�9���`ˀ��2Z���qo�F���{��xk3z��� ~�:p��T����}�y���X�����)�=ίE��=^yGcݍ	]�e`ۃ+c�*9����ݏkx<�û¼���t��wۭ�K��_��ǽXztX9&	O#/;�rz���&�.�|�Ɩ{2��eشx�v�)Rh�9e��_ں�Ηy̵cv��5������^�OL�i�.�{�>uc��~��-uc��ۻ����Kez��¦>�@S��w9����>o�ﳍ���K�̋�ђ�zA�l�sڼ�^��U�t�ٽ����L��6G`/Et��d�s!�wY�k��r�w��M>ml�z\^W�`kBv�X#��`/?Z%_�g{/;$曻^���i�N����`3�0�q��J�跟ᗃ�}�
j��$ԯ��}�d���.�R��bz�����_�J�p:�C�:m�ZsCN��Bݮ����c�Ov�U:���Ѱ7K�0$�4���ɽ��f�:8�e_j�ϡ{���<�V��Y:*$�by�h�m�7u�K.�9���"�����Eׯm�����;�P֒�u�+Gx�=�j�C%����嶘t)�������|>��m�SW�7�5(���������k���Vk����6��8 �m��M�*=é�����m��u�<��X{[��Q�{&�7����X�D��ڼ[��{r��9Yހ��a}<}�����g��7��-1�~����Ϸ�s��sxT�ud�pM=�v�y;>��d�U��v��M�ϥ��{�*]����9���E=5�ݩYT'��]��Q9-��)�}۬Θ]�)z�l��Bʋ�=��zts|����8:&E�x��{�H�i>���"�#��l��T�k�`�>�9&	W���˸j��J$�n�:�;g^M��v;��K�]0���Vs�s-_��أ�;+՝17�:���>r���}+�C��	���i{�S:�y��������E<6o��u#q���O=cd��>9ƌn�.�"�D�W��4Fw�m�]���A�)�7Ҏ>.�tj�y��hD�+
w��XGl��cuP�����Y&(���A\6j�z���HXN��&��Y��/.uԂ�bj��cCF���-L�Y<Ɩ�w,����SXhb�r���rs;
�RT;oW�| >y����U�+ǘ�wz��ĝs �:e��7k�z9���y�EN�ɥOqs��/�e4���ڪ����=�.+S����ϣ�\��'n:o"��y�����ﮃ����Ӹv):���sʌ�E�/ f��s���M�t������G/���ۖ��_�ҹ��*�Mv�\�u]���W���[	Y+�M��k��~��f�7���w�u Ӌ|r{:��ZVu<_ct1�~+[��N>���eS�-�1����#�w��<���|��/m�oN�=��Mϵ���%pr'r�bv�]2p�Tb�2��՟I�穽�)���x�OM�O������m�q����ږ�g���Mu�~N��؂����l襜�1kc�����')Nk��TƩ?!v�{��{8j$;^�R�%�=��s~��=/���u?M̝��[��uJ?#�n��w0PI����5,�z��;�(�~,Wk��ӴC��;��^r����]1yYJ�ݜxS�yb��ٝa�K1�И��;�Rt�8j�����ͅG�Um���u<"�=�c7�˻v�I�a-����﫽�y�fj!��i,F����-¹�յ�'^���c�:5����gy�2K���)n'皷��
�x�M��v�>���GK=�=��|!�r�^��ҳl��W��H�����Ϝ���!4����Ի��s}qo/b��G���ڧW-nI[�t.V�����{���@ u�S�~])l�KKN^#����1^>�Y�N;���THҔ+#c{��CC%�X��WKl�}	����R��]!�̤�J��JJ���AyS5]��d��]�=��s�L���t4�^�A�N��e84���E���������jz��'nZ���.s�W����\W75p�Re�+���5w���f;r�_�V�k���u��N�w9N�7g�r>�Z�<��uĲ�9�	*�3���S�/)�}�/M�o����[�I�V�������,��̈́8v�M�7H1����d�F�*wv.�y�&�� ���i4�����7m>�N�o�0E
�5�<��]��[�p뛲�;��*��s�D/RW;�eа8V�nr0孏��.+諭�E='y���=�ۏo^��uc��NA�Fw�4,CEԬ�̉d�$�+ק8�`�n.���w���w��6�{����=V�]��̩��Y��I���ݴ�jvsw�}��}�_����ߵi���)~��G��}\���w�0Ͻ�D=cZ\j�'�j�Gϊ��Z7��y���{ee�O}>r�d��ɻ[�I��/���Y^LNn��<�Vwz:Uo�	x�)=&�U�c�ۛ��ivy���&�,L��W��sr�G���3��}NI�SɁ���OW��&y`]��=�l����u�a��WW����Z�����sƻz�5@�Tu������S�E���&�/��z)F�Z���c8v�o`ޮz��VnOO8Mo���'�>�:z�?���g���3v`��ɾ�C6��AE�ye�o���7��졿o0�82�nlF8�S�KZCV��èL�B����KF�[��}���p�L�s���)�ǝ��Iu��_esO������V!��6��댷��Y�r2�SW;1N}��x�=;����{��ﾯ��z;�V;mߛs��S��8t���v�"�Q�D9�dO����yt��s�.���P�E��K��z��'a�$��^�S ��і1f�S�r�y��ו�xu�|߇F&1��\���J��U��|^ߓ2�s���n�N�aߙ���7꿹�3���,��<�[����[}���ٷu6�9�ׇ{kjM�ǻ1�wu���j�r
�/�b��������Yu���E�6U��;��n's-���cޗ뾴�5�UD=�C��,v�:���N����4sө%�t�o�ᥞu:�̳/|���mvdO^��'�U��#�[8��f��wh'���@���7���pȔ�G�E�T��}I�r3}S�,M�z�$���8���a�2fF�%~<�T�u8��a~'�ϒy#�N����^��2�t��OB����x��>�2`+&uèT�P�̏�w��RR�37K8���hے�K����m�IS�V�b����o6��"�#8'.v�Aኺ�Z$̷���v�Z��RW.��d��i�֞���S@��k��&���][�(ыq������ow��Yy�㿁��H���0�s�}}NI�U��0�[^��nf�c}8ʫ�[��vֻ�`.�=�90ߵJ�g2ՎrIc��R�ck�B{Nzmw<�.����x&Bh�s�=�Fݮz.�/Vz?mlb�_r�y�[������X6�s������/�s�|cu�Ij/0���u��������LͲ���Hڕ�Y2;�膉��wat�8<<6�Lݜ�>Ň���*�rʯa��K~b["Y�_�z�9�A�Lۙ�}�¶��Q��� D�ϟ��߯P�v|^zA3{|��Y�}:��a�$�|,s:#^�}E�L2|��F���������1;_�(Yn��24��D���+^t>�:�W�I� ר�Jvh�ll/|���X�z��1�w�U����r
�6��R�c�ʱ�jvC�۸)�D{H�jn���M�a4�7���z��.+Y$���*X�w,9c<�'����im�oS�� �GyU��Vg�d�1M��Z��9�{:XU��y1��3��Ŕ�h�c1-ʻ��"$��S�i0��"��rP�OyDsd��=8�yw~�}��>��d�����mgOJ�v�*Ð(��ܰNķ�N��,ŶU��'�};�2����Ǜ����y��������P���-�wP�	[��N�����7Ul���fN�0�r��󿺩望���r���'��}�mEܛ.���i;�Z6��PݙW�YV�{Փd�������r�2V\�xϒz��ޣ��{'��%��v���H؜c��|��y��i�`��[�`ǀ�%�ݲ�o���o���`��+��)��l�%v��JNH���SS=E��>��s�E��k����2E�Y\�k�������Խ_������u�̹[q�����!��I ��xr��-L��Σ����X:q�ٔ:nҕ?oo�xI�<�:%t�U�X~��Y��ϵ|�QtGmX�����ل&����ߤa��yo�X�HP�
ʇ�������i�{��w�񬧝]0��ʺ��c��V(U�z�2Ǳw"�7˩�=�����mLPq�Ů;]�r74J��]�=��>r#� n`ū��r��y�+��W!vXg���:m]gc�{~�j�hse���������w����G�~��Х��6Gg���(s�m��+���Y*��%�f"h7�Y��gd�lIqZ���5�7)I���*\�*��sدu�.rk��Ǆzy.�	��nZ�O�J��M�ƽE�[�ך�<V���^�O�\�#&�'r7��}!�d,�%-2W�U)ԧb�ţN�~�jwQm{��	����I�	\��gj�җ��ꇞ�_�e;���";��{|�Y��~|��sإG��o�[و鴚��m���������u������z�ݤ�n
xv���磿����ǼFk�o�7���Eb����;7���f^�"�z�?��5?��[���w����7�zI�}�}�s�e�7��o�)�{�1�C�F/y���E��<R��yۛ�B�mxW�������.��*�9=�6?W�<�û����C�Ap�c�r�<��#y�����b�SG�?h���3p��M�]�ͳ|-�R�2���p�@=�N�68�Z�F˦2��� �f�e�/�j����s�I:�e���\�u}.�Bn�������×,.��V�@{F��
��M�Z.�Mon1��Й��Վ���d<T�n�$�rSLH~#J�1�������,=��Q������H���U�4w��V���Z��B�L5�%�|Z�m�=��S���[�/���OygF�9��އ���2��F�yy����$�mP�I��fT�;/(N,�l˫T��\K�p���r��ld%'9��0a��3qQXXcl\�(��}�k�*m仾���M4�vim�i��f�����y�V�;��<���
3%b��Q7 LK��D;r���4��9!zs�=�þp���u�H G 6p��k�W��a��Rs�n��٨{l���V��s��Fp�2�N{oyu�� Nh�U,X���g���y�\�D,[��l�=���\��j��]���_1��JA�:���u��E�>���'��]�!��e�T�cSu�ݰ-(Gz<��ׄD�ˤ,�F��Ȩd�\m�sRS����aٺ�%��Y�s
��E���n��n�X&�@;�^�N.|7�_������|VfY=B����쳷��� 6'2���b�����*뾠Ў�c]��-x��9
�� ���N�Ç���t��J����6��RÐK�e*��.p=M�8��G�� d�f�y�Y�ڏ��%EL���|zWuuR*�\���:Ye�U�蘎V�A�{ģ�t�k���MK@gf۔��{���1d�m!S����Z�t�^�uf�V�*HE�\�+�P�ԫ��Wv�X:�|��,o-�E�U3L>�`DA�1R�{�[���"1[�no^Uհ4�5G^c�N�W��N�
miI_%%������*'��Eޮ�o�d��0c-���55e�v;�Ps�n�5�-[ޘљ+����������]��E}�����7>���2�j��Q�p��oPÉ�t���Z$���;��]�ݙI�������U����b��Q�y��,�r�Y��\��}N�9��݇rix�n�o��.[��I&�zfjj�8z�GS�-�\�8�Z��Y�u�J��]{��hA]����tRk�I������G���N���tǵӻf�:�?�Ӂ"�uJ��YC��=��)��u̮�aԻ��	S^S������]���j�(I��r��w`��Pc2�]��'�tqt�SabM3��B�:л��$��{�����N����[ӈ�飭֪\;f�u��v~b������_n�mX�Zm^��׹t1!������n��G�uv�\5��͂u5|����o{�����߱��P�V�UU��QV���kA����(�VQ�X�P��
��
��TETb�E
����-
���+�r�A#�V
�qV"*��֘��(��K2�.dRb�*(�k1��DE+DX5��m�QQ�m(�[e+�̲���d�n\�m-3��F`�*�hU-(*�U�J"���Uc`�"�+*Uh�R� �U�QE��1�E˙X����%P��KD� �UH��kKEX֊(�FZZ"��l*VQ��IY*,cZ؋-�cT�(����V8�UUdV+X"���Q[J,QQ����X(�Ȳ"��)b�iX"(ĭE��
#YT�J��DAT*X�E�b��e��PUZ¹B�ʈ�-�%EQPF1DE*4(Vm+X��-
� �ff#��a�DD-(��*��ffRҋUR�-� �T(���7��W��o�V����޲�}�vQ.��M��Ks�t�|�"e%D�u�����Y��c]���i��ָ��?����o��ޭ��R���u������K�rSɃ��9<��w"�],fx���msRC �o;��X�w������s-_�ۿ�w3˹�VW]:f]V��E]����8}����GwR>�ί�ku6�좳)�{�\/��d���7���v�㇭���������{��FjV�X��צ�K���s��A�.tV���L��|ݡ�����rdmC7~�7�<��V�5��W�Q��W(��Y��KY8z�.���ʴ��fNSbsڽ�h�1���y�.��v��1�r�║�������n��;m�ϫ���C_t7&tz�_�)x�1*JS���/r�`�g2�?=q�mwi���Q��/�WNm�Ƕ7˶I�z�}�d؄ZF����'�]��nS�l���Ck*��y׆:W�+��y��:�K���$N<��݋/ӱ4�䖶nVΣ]c�D��L<��J���`#�t��Q�X��&��˴U�\�l�ﳲwu�)� �§d|�3��+�P�8���T��)�L"���J�iun��yC�z+���ϵ
�[����C���ﾮ����lW~­��\��ܱ_���}=��=�/��_��V�.r�/2��-�/�����r#-�MuIۧ�@��zƿ��N�{b�3O�������k�se{�k���yߣ�ފ{*kJ��>�5筵��r�6D���d���t=�h��Azy�꧱˜�Ok{�����.?mGvμ�x)A{�0�LN��/����Ϣ�rOo*9/հAm����`�>�z�v޾�uC��]�Y�/��Dگ>�HDw�*k��W�^�t�O�S7��w<v���nd$>����>���X�O<�����W��ۿ�C=Z�s���l�<t��d��u�ԖZ�]ˎ��+/�Y\��h�=�ܗ��^F�H�z!�;��R��L��_����e����o/��e&�_��ԛB�EaO[4�&כ�_]�]��/D�k��;��lm�=���5�}|��ڻ��68;+���J�ӱ�zi�rʹf�M�0g���5N�.�˸Q�p���ת�1+yD"��oHd��7��R��Z.��L��nd�#��嫉�μU׷ۡ4����Iɾ1+�m���҈�3>ވvx^u:7��;hMܹ����[�Q-^]��~���ɂ,	��Z�>#��^�a��ښ�Wj|@���19C����RL3�3��yi'�>óɬ�o��Q��1��{W}h���Շ7$#�%���͗��G�]��/x��k���|��W�{p̡�=�uW�X�`9}���h7Nz4��i�L�7�@�ř^���m�{�7ý�mՀ�#xs�7�~t*����{��Y�wh�X�W�қ&y��s�Q\��E�V�{+-�zy��U�3�ު������wΔX��/�Q~�x�nؕr݇��.pۯt�}bze����#��z�5Y�躳%d�Su����%wp+ ��c1G�����{V��z���)��8��
x��#C�1+��*��ѩ���<�A��4uL��Y���*��o�^��6L���M��m��+�M�����Ԇ��8��w�#���:i�<r5��<ѱ�Yx/�Q�nCe�C�\|Py�pA�4;�Ŏ�}��6����@���9���~��HZͦ+m{$��9&	O& �ogH�+����m#u�F+��J�!�,r�w_��_ں�Η�˔��A��|�oc����n(�l»��{��ow��R�4D�Vc����3�t�}����o��\wJ���ak�.W���E��$�U����nFi��וxWf��{] ��&ݙ#p�L�5jzۘ�}���!�����N-����+��y����ح�5w�v}&�.+
z�6�L��\�u=Ȇ<��nh}}a,�vm���f1��^H�y��I�r��%Wv;)�g���M�Ok�VǷ]{�0Fy\�J�}2W�s̃�O�Ib����6X�j�f�i�m��2�n���[�-�IW;�ҍz�5D�^N����e�է����-�����o���<�[�^\�p�T��g�X&r���T����&_S7
��H��.��I�<�>KN��vvR�;x�\���*L\�E����m����#��lT���zyח�Un����g���v����fN�빭�\�T������a��v����������F{�«��~�����u�fu���f�]��+]��<��ܙ��a�����æޯ�sz��u`�N	��wh+����Ӛ�l�]鈅"���[]���n}.�g�>�����ݼ�F�!���GZ��|_s�M�;0r�mL�F�� ���]Nc�=�9=�����<��͓t(U���+�Oa]뮧u�س���}
rLSΏ:$��rH8��޹�=�f������.�ʄ�ep�R��}��V9��B��Ҳ��{�J��y����U��$�����]���/~�&f�Xۯ{�����^�<:����v̞:z�0݅��Do~��r>/8��R��5�&�g��s��}]:7��nN;'���2���v�� ��M+K>���n�ﲚfj�?@{�w�>�R�9�<��*I_k�n>���-�
�}jc�O4����Rez˯�.��-{|P\�zg-����|�86�X5���A�u\���^I�V��JB&�f�uɓ��ׂG��lT'K��啜`�R��T瓸.N"cZU��-TW־��ok+ �����ꃙ�9WG������7˴;�7|���ӧw|_��f;˚b����eb.�*�5�)پ
�G�@��|�r�r�i~�J�<Xo}��5����{�8)�Uy8=հ�r���@ڡ���z�\�w�[��pM=q`\��hO�+��.W�������OH�S>�1��R�y��aj��m���f�75���`�a��;�X��n��G���|��SB�"��H��1uR͎�Ww,�:S���wz�����+;��[��]Y�q{�<s�֨}g���'���齙UѥwYG�ObK�}�W4���C��R��k���ܝm:��T����f��ӨI^�Z��[�C�y��SZw$�����a�Q�3��p�N��lԫ�5�&މ��h�վ�m^\����o<�.�=�91�`�������<��z������.=�|*@w��0���mwzh�ϱ�=/k�s;���^G9z=:��S��R����Ϲ�<Go�}�"�+#\6�Ur����3R���*u�q����K��w�����Yݺ��+�-<b�u�Ƚ���>�7މ�ҷl�W���uϏ�>{o���X�^}�[�獳�2f�j�������uB��:�bPq��5�����d��Wfi�g��v�d�5�4ߎ�=�et�َ�9�R�K�oT�����͑3hw����%�wxoG��{�~�&U�Y^�A6���Ry�p����r]<�`�ɸ �tGާ�>��銸E|w���/:�N�/=+�8�ɐ�]��o#j�6oSL-��>޷f{&|���-I�p�Kݳ,9C4�9-�UPl�r�=�*�]���c����%l��JjG�}Aevym�}+�l�wV=�5����]D�Ӑ9%\�}�Igk�yS/�~�%�^����9�t��kp�������;%����ݬJ��lP��XsA�Mxs��S�7Ҧ������M$�<��,������G��ygc��QT��L,�\���ni\��ܪxςT�k�>Lv����}�a��M�1/�:�H� ��K�Z��2�xWw�_r����іocQW�3�%�إ�	ƪme����вd�Yʑ����(ovՇ݄㽸�Śhp��7bN{�}�����D�ǖ�����I٘z�ݤ����[i㻛�N8՚d��#ow����5�-^�f��vbS�V�{�|ԯX���0���U���:>��=�ݛ�'��Od�"�ʯM��}9�?`��JLO���\�L��&f�}*�؄�� 矈����տOr߹D�U���;��k����"��[�p�����J��ci���Vs���"w9��rmpv���]�!S+%�d\�O��O_�c�sΗ��WgJ�eʟlt�q��>��Q �d���gA��*�0,/�BUVy�VATzn��D�R��O�5����H߽W��y�o\���1�݅�܏�z�ګ�v}���d%�2#����躶�tV��㚦O�#��@�R�|�jƣ��JM[�yw�E.꘣���.���X�2_�rꌻJ��z/��w�M�Ph�l�]Kk��{L���e��Y��,8�Z��%V�]>yj��6�OaPk�P͟
7iS����,|�&#�}ċΥk�OyU��tb��Ք�]������_�|�V�R�ƹ�n���쓪�=��s��U}O�>��=A���R�Zo���.q�[�r�䬙�X%XuI�W�N�H�����9�Yg�|��Ǳ���켤�	�U�g�����2�Q�>�Kvo��ڤ�X=��Rf[�f����U���9^����͸��˯#3�h����`>�=���Mw�*���;<e��2m�1�;JS;�H�;�+��u��gv�٩��ѧ���Z���[#���Z���7��t�_�y8����hYT7FD�;0�����s]:�{l��j�^����'qM����E=�|�m{��s�l��p�7R��]��*��r�;�N��c����y9�\�|�F���_���x{������7�^;>7t
�r��a�����+��,����^�;ዟ]�=)6�~�$��Nu�ɯ����%=b�wX�3��2�~7�d��t]r��%�}�7��z����;�Hq��7��N��.�WD(�
�/��&��u�n�7��eL�j��ي�edJ�s�+5��^tκ@�#s)%L�G����}���\�TV3o���˚-T�"��KsY�9�[
�զ92s�	���U_w�w�;�mY�I�������w](ٝ�&��Du��e����sm�~l^�m87�� u�>�E�2x������F6�y+�5OsN�H\wn�K�����NF�������n3���v_f^v�`����.~��G?��VS秎\���>�UޏFK�����1uf�N��<#{��b����D���C�����0���c��hjJ��ز�+y�黣h��w.ã�Cr�#��l����:�R�F$K�}��S�Chd�회�+p?$rt�����.��[@��Nf[�}����FS݉�kΦf�^{P��IWU;�҈mg��ٿL��~��;Y=���!�8����������~���v�*�q�N1S�e��c'��7{�c�u��r��I�V鏳澿��3SR�M��������Ԓn�ܭ�Z�=��pUwd�O. +j��./4�;+:ȸ�Ws��9��tmm=\�yX��;K��G]ӣM22��43�,r�%⵶I��ă;6���F>s����5uO�h��	gj[&���ŕ�+�����L�3>--�(��v�:���Qk��ul���y��p�u��'67krF���oQ��Z�L����ӕ�}1��2&�
�ea�u]e=}��j���Ň{8އ��/�tWu���b�{
h�7wj��]X������ݮ|/9>�#C�ß"nY�v��uof	(ʳ�D��v֩q���{��Λז�t�Dow*��Q���s�w.T�
���ko�@.��@^�#��Ěu)�+ǋcT�.�h�� �u1m�����O�s\F��t���lі���K!�[n�YyS5��R	A:Xh�E8inN͂���QޭaV(��rg�1�v���I8��IN��n���;�{�d�m��!�7�*���6<c�s��tv-���[3o+^,�B�<]ewqcmQ4���W�6��.Hu�ebR�,�쮌�7K@����7V�p9��f�ԇJݿ�;fbJ���z�����ݬʕ���r\�u�2=�Dn���8� &�ۀ�D��+�5�*��KqS�!�9�8�sϵ�x��Γ��˘�N̙�7�]�W��IE'\�nC:^ԁ!�X5�i�2Ȁ��$��x�DX�hst ���gd��ma��+�{�G]
��7����u�,ƒܻ�����R"ns���Ok>����}̃{]Lc�`RnU��u��\
=��:%R��>y��ζ�:�u��k�ה����F��S	lj�7]�Ʒ�ea��1�ysdfGsE��H�B�=y�,Y4��(�*;j	�\�͹6�5�LɎc���S����F�D��/��cY��j�d�1�us$<9�g����FiKm��Ò�= ��o�)s %S�v�����,e@���Y36SȒG��R��Xt�9�x�����'�}Il����PK�7�����sb�[�o��5���w��]B�d�<��;���c�e�ޜ5�����'��C��c&�bqb���,j�ix�����~����Ԑ�Wl!_\K.b�;/h�2Rr<\D�ˍ0�r��E
���1��PM���l��tt�ީV{����"\�grh�Ts����\zS�:	[��Ԇ�̎���8�ƕ�u�H��B0w's$̭�뽠��:�<��Ε����_3e�7��ۣw8Wr�t��:�Nc�u=�.���B�EvZ���(6'#}�k���H��Vdޘ����}��o�l#�(�g[�*K�7G(v9�ф��B�,���u��S�Ί2�3��&;�:�v�'`]�-*H�K��H��Q6�(k�U���:XW��Q��=vMp���"�5�m�#�]J�v�R!�E��J�[�L�z�N�|�V�'�v	���xq��}A@X��+�YP�J(�lTUA�\JcEc�VPĮ7.`�T.\DLs
�
�*���e�����Lj��n8
̲���R�DFڳ((Qr�$Q�eldm�ˉ�Z���3�Y\�����1k�
*��UKK3&[U(�J���9-�Kl��b�b���TİU)U�8
&Qh&\ʨ��F�Q�m�ʃ��Z�%��U,m.\e�UUb��E��IV�J.%-��h��*�$�*Q[b6ؘ�ت�����)�b&��QŴ*"�"#-AD2�"�V�d`���r�*�bQEaj5��Ƣ�\J5
L�*,DAd�QQW,(� �,[e�V�#-)�(�? �}�7s�N�S���!}�)�z��L��,�Uו\����g6swu��B?n�
���@.Ka��/X�f�z�p���5�w0�U��}_'��>��lkY<�'�=�:NQ����g�?R|�����ܻI�ʤ�X#��Cqmd��+|�yw	��q��;	F���{-�]:6����1g<<��e�W���T���3��^Я>H��b�k�}ee����*��v�k~�`x ]�>z)�)�ڊ�KrC�b�o�Ik=�Pg�(d�+��ms㷽���	���ھxm?�����f��#�������e��J�b8��]��>��/Sw�}@@�p�G}�;�ׯ��~�ӏێ�<���Kz�ďT�'!,%+���J�*[������|U�WB9�o�{�6���R{�w�;k��^�π��W��jt�3+���걮{x�G��奜�Ҕ�-�ӹ�nؒ�����Ra�Ҿ^�a£����bd�V�b�BB�3V٣3.��[}Cۋ�hҬv4�C����"�{V%A�떴�;�)��Vm"f�QcNP����5S�&i��������ZZ�dDȴC�]�����!�.�����wg%�@T.�_r�o�����g>}��G/w�rq�[�ĕ��W�G���\��Wr�Q�J�1o�}��)�C�F{���w�' �%\�}�%��seX�3���[�4ǽ�lb�;�ܮ{cs+;�����*܂64N��i�ċ&�S}�7��l��}I�/�&�<|�8�f��(�^�}^[�2����9�7*��ׅ���Y�z�ݯ��]ϳ�}���SK�,��ܗ�l�i^z˹5�>������[���k>����*�.s�&�ר��=�v��۹�2��<����v�v�T]'�-��Μ;�_z����^>����u76U펏m�j��z�f*�[S�WV��ӫ�Dv�j�����C9�c��%<��]��'��>->��ٺ��Ǿ��1a3�n���])�M���t��9�+c�%Y��r�z�f�X��*g��ܚo)��}�k���.;���8f�7�zv�ڎ�:^�����S��F�-K�d�|���Dev����:u��x�˳6���:D�79t.M_��/�/Mm�!Ŭcm�eu#��!�u��z��$�������^����t/\�nOdG��_M���q�V:훧���{��j��{��j�ސ���˻L����I�:��{3���;Y>��{D�k���x�c'���r�ʷ�3��?�4��v�kk������^����aO\���A'��y]�I��y'�#���yM}�����|\���[��`k�̮���[\"�q.�ϪU�3JS���fo�{�}�/nʿ����(G�5ձ�8?�U�~�	<��u5z^K�;�ՎZ:fgyl���^=��K6kܳ7C���s����or.y`ޚ�R�����S�`k��*�j����c��&P��:k�1x��ں�����;�)ؗ	~���nSç���+�f�I�g�Y�˨2��ꛃ��L������ud�r��}gw�QW�w�*�3x�Y��8/��:�)���	� ��jM"�YsZ�7�y�哸K�g��e���V6�7T:��y�gis���9�)��p�<���q˖������ٵ+���o5u�G����zdX�����<��G����;��V<8�ci�bp7-�{�ƻ\K{�pN6�;�V���`���=� Tx'�d��U"�Y�ٝ��/s{��_���J����ư�?����Ng�\�r{h�i�ҩ҂�u��|�|���t_P6�+~�Q��^}I����3>�c ��0�k��v����3�{��c�M|]ʾ y�J�i���	u�=����%��٥3__һ�=���WI	Á�v)q3���SX����ղ�;:����Js�C�&�>x�g��[������0�������)e,�wF.��=���ۜd�l8t̟70�دp�s=j��Yo�P]��n
>�A�d�����E�ѯK��s�Yp����1���
s��n��i����8ߨr��	����{v~���:����E�P��xG�/���;�����O�o��k`2��k��J���f����7�µ�OXK��k#)�+���>�s��y-5w�o�>REW�l�6mo`�=�3��xyέ��+b��\vs��l�o��u�*�`�&�nK�M��s�_`�λ9�U��6侜oOdX����{�g�ne{���C��J��K������n=[iJ�]� �o,��Nn�V{+�w��p� �l�(��S�/*����}��7�V�N����W�~�7&�Y������%_�u��Fϳ�420����N�D��cd���q� ��{ζ���T���ӧ8x}#�^��b6�{#��14�^ʲpC�~�6����*��������y���:��%N���'l���71)���F=�7��^�Z��+
.~��3j_�r*�=�׫��N�<}~�ix��+�N�px^zg��+�lj�y�y�(:��f�B�o�d�����5�W�<��y�+��yQL���8-m⃤}��s�� ����rG)�vyǴ�a|V�ެ��u���O��9���}�]����ǥ`�%8�ƻo���O�q�=p'b�R������]}I��.&���(��(�������Pz�Iv�3�����o�	�o����&t�s9�T���+[��t�'Va�R�{R�)�:������%��N�\��8��F&nɿX��]���8�5}�Vv�����܌��ow�����<Ð��}��9����}�R�#e�)`�#��=�.�%���./'��G�����|����m-_������#x�[QH���sV���hS'��g���5�y{;��*/#w�f������_���n��\��L`M�Rq�����{k7�y<��=.S��X�^�I��q��1ۖ��V�d���|z�-���@�~�M�~���f^��:�ie��9%\�}�RZ��%	��`Ozs��MY���۹�W��ۙY1���Ձ�īr
�6v�����J/��.}�S��a���L��|�f�~�1����ټ}���1��j��z��p��v%��z�ݠ�K]��^sJew�Wo�gӷ�#��sT}�����rW~�[t"�e��Ut:>\)s�bמ�X{�kz�VBp�"w�%����*RQ"H�����׸�/)�0����֭���*�wu�Ѭ��J�N�:�k�����tea�Q����ZT�\����E;d�4;�Euk8��P�B�1���N�
sË��G��:�;.B+�{��W����s�/웵��Ѵ/{wB^����n��p���}n�͔~��Qr����%^����{ڷ>���y�=
 �nwY�a=��]�[�r��7Ϫ�ϜX�I��L���ʫ��eLP0UWwCë��uss��]��
�b���5vt�9�+d����\�!g���L��	��<�O{'���!4_
��;�F7�]C[5w��k�k��Q�)��<:���E�0O=x�n���q��\������\���o��{z�fes�f������|��.��$���=��gx��9[�Cy:҇<~�r�����H���-N���W���0R�vG��Jj@��[�woC���9�yg�.!_%���
r�$_��1�"D-JƳ�2`��R�bR�eY����1)پ(ϵQG��}Eq�!�
�ڰ�f�6錙�]U��߯ީN��Rۨ�|���=q'��<�q��c3�Ͳ|�tq�����(9{:EV��-�CA ^m8�R�HZvML���o�p��|:�vv�ρ�m'��n�3݀}�y�,^��r5�N%ȗ9���X��׆�k$췜g��oD���wX��Ԧk�~w<�"�������x�0W[�߅p����r0�!���ɾd��L��o�,#�	�[���~�X��z/e���u׶����
�"6�nr�}y�t�p}�F	�d˔%{��Ui�U��P��6uht��N6�.��{��T`�t�_0sr���O.���mW�mx��8�HS�%u� ��y/5z�j�s��Ǒ�����=a��uo�h=r�-��=,٫���^�
����3�z_�"C���,Ua�,�[��y2q������fr��xN��'j0�M�u+�c�'�y����G�h���J'nS�b�.@{e[�ַ���tB�kp�Gw��r�<5חmu���x��d���$Wő|�*����r���j�1����y)�z�?p���x���D+�K�u��-v_i�Rx&���U*Ms�V�Od����������x��Pjf����4+>�`�n7�h�߈��ZW&YI>���Ӓ��+r�{Vέ�n�y(�ԘS
�	��k���٘G75�u������ˣR��n,�e{5׷����F��5ش���/����p)�ٵ�����Q亠�Mt�:ۍ�vv����&�Z��ŷW�C�$#��o3''X�w-�{�����f���d~<�U�+@Ň���wzX��o�+�s�`��"�Լ�m*�p���xgU���5��z�X)��!��ⲽ3@}�ŖV����c��T!p���F����K��{���О�Mg�ԁ{
z���dX�X~�s�Oo���n	l������}���[da齘��+�x:�tԊґ�@�Ix�_WS���]��vMs�.^߯T�d�-wx E�3}|S�e�%YG�v!VK��Aw-��5��~�.1~�Y��o"����\ë�銚��eD��>�Ą���&�m^�X�����꿔]�ՅY,�VK�ێ?�?F�;.z�?@���V�6D߽�k;������nɹ�u�O������^e�|Ϩ��}}��O�j�&}fZӣ~ν��;�fxV'u;�\��Ս^|�@����ܙ!D��Gs�por��Q�eU/���b����u�n�e�]�e�Pþ��VKeʮ���u�L�̹9�v]�po=s�c������>�gXG���.��]��
/a��z?D�����˽��i�f:�}z���b]�+�2;��;).抉o!^-${ڋ#s/�tо�"d�1c�x+f�	�"���7�r-�w՜�kD�;ڎ�u�gsE���y��^ǃ(�*�]��l"������w�Ѳ���'S�᝔����9�����q�޺��ǻ����?W��cTo��x"V�x �=0Z6:�nN�Q�T�r�N�L�ʿ��;��uP��U����~��mo����N��]�@f���ji~����f���Gb�5[W��o�D*��2-�XDϙy���.3��O\������IJ��_�%c#HW�F�ܠ�5T�J���u��i��FP�V�g�똥l���Ewx,�'L�l�2�`]�`��w�l��Y�;���������]��i�t��Oݯу���dA��dd��\�k�e44�AJmR\Y�Dx��h{��t��X(�����I�՜�vO�;��R��p9_(��Al�y��U���G��Jޗ3ח��̴��Dd�{Z�o(tt�r���;2��D��|���"z�~�Cr��zZ�v��t�y���2�k4�v=�,:���5�ha�.�&�����/���3�{Ν�7u.rV`ߔq�VZ⇖܋=Ԉ����6��J-R�7#V7�4���QtV�^�E�ǳ�-�Y����h��z��T�N���Cgq��U�q��wI4r��<5d$� J)G=ˊ�%Y��KFI���)��0�
������]+��@0w>�t�[v�EԚ�8q�P���wp�6W!���I���VUu�){S7c�B̈́c�x[� ������v��ݝ9�o�`��9��w\����5�)����gk��R��#ǉ"��у��(�uu��0��	`�ǝS7-I*���&�yG엽YL�[oM4���ظ<pc�;KH�]Y�e�X���hz�k�(]��06�XQ��L�CW=�eot]��C��Mx�`n�/w$�	��D�@��Vf�6�è5�����Y��b�,�g��������VC�VV��7Υp�����S+9i#��z�u�\:j�R�������[z��.Ys����5��*�&�njK������-�uԡ]�P^#[\�3��0�����X��qƓ�7���M�lO��n�.��5և�vë���\d�Uh-�6�>�Eh��D�n��n�Yl����+�vR�1w+Cj$��a���[OV�x)�3w��}-T��Y��|�0LM#+Dy���y��Mj�g3�d�ڃ����7|��i�&]��* �vπ"1�<�7�����5W؏m�¶�T��:�7��[}`��;XrV�t@=h��:��8�w���r��$�8�G�fX���v��	�A�]�qYՇ3�܊H!�hJ��2Ϫ̽��!|��`�G�e������͵������~zʜKt�ou*
�cj����f�l���E��Z���wC�>���#��/��]�!��&Vq���\�H��.���^�T��Y�����o|����´6�ۈuih ��c�7U�1]����!�x�6x�58P�j$VJE��Y��./�\:F�+F:�>:�7h�bi��tE���+*:1$6@����=ɝ|�$F�ݒb7�h���z*��=St�whv�ַMlB�]Y�f�����Ɔ��	���^�2a~3�5���Ns��]˺K�╹4v8t��˫ew.�:�=g��S㘲�*ƧO�  ����+��l���ͮ�����u�Ób��=g��b4�M.��s��b�b�c��zm�{#.mq}��ۮs�(�u.bmL�3��K�W�]�[0գu)�I��F�_G�k��� �����g��]Vn��y��m>S��_rډ�dZw
";3�jB��klD9o�RE���g@���,��֠���NV�[�6,�c�x'�P��eGs�+�h9A��iZ@d�bf
|l��ef?�V�ȳ�!:�S���G��m+�c�kw�s��i�#����#���P4�<�>zD:y���ݫv���wР�0��1z��ʙdS���o�[̀>�a�^�5���F�X�#��wg]Mw;�%�_I7�A��rb�1PE�(�ZX.Z�+�p,QYZ�8�V,\n%�UDPb��#mbĹ�*�cb-h0EX�h�2"����%�E����b"&Z"[PPT�U���U"&fL�lLJ6�Qưna��Dm�PD��kT-��T�U?e��:l����Q5Kt�V*�iX,TED(�*1��[.��Y1+V�*�%��®R�[qA�8Z"(*(%ekF5*�E
�
��ժ�*�(�m�J�F9ekUAPF*9n%�UQ.ar�V��kZe�`"��� �i���5h� ��2�5h���!������e
0J��ۂQTY*ḭ��V�Q�ˊ�iuk4ш���ZTjUFQJSN9��2�\LK�q���Qf4D���k�wV��yj�nv��v�A3Zq2�(,�jVu�El��CXѐ�Y\�l��y�"<+�p��Xǝ����9}���X�C��0m�}�5n&wޗ�07o�~��+r� �*ڗ�4n�ړ뷛���5�Z4=R��k�tg(�5f/Zz��g1U�u�u� �=\����>�<Q��e���,����T�1���US�P�:�[�&�Š��m펋^/uT�{��Vz�8Q�\����\�Ϥ{{j�v�X%�x���+*�t��Eˮ�US͆'ڪ�] ��
��]Xg�P�'*����Y��]��W�'֎��$�
���9x]Q�.����	�Ʀ�\�4�SB�}�ɃN	�~U��K�t���n{���8�b�����L]k�tH�_M�x����X�䕠K��P���^��V�-Vf-=�wS"��L�����oꪜ�[�[�"7�]�s6��	1Ӗ��z�^��k�2}������u����bJ�+��N��-Pf��.��z�Q��c73h37����(�i���}+����q�$�|�p4��+2�U��S��*�l�uf|�ד���n�{=��nVc㲙�U� ��~T�E s��?��	�E���yW�CC;�}
4�gBn�vt��������51tU�2�H��/e]b[�SW#ޫ��/�35��w9wX���-1΂>,f���'BTc��K�F��n㽬�x�;νw�L��;�3����%0l�I���<y�W���㍬�b~�A{�>�ON��l�"�w܋XD�����^>5��=	�5����{��B�{ࣜ��h2{��D��B�����>[��/�C(q�R��.Xڬ�ѽ~Kz�~�e�;-s�!:�X�b*(���>���#�*�A�c}h�C�Q���2d[�6X7�7S}���T��T��V8�b���k>wWH<*����b��p�0W[��\*���݃z��=c���:|�G.~ߧynҶ]pwXj1\l��K�u`�ȏ���-���=���'�S�����~4♂�5��u��Ǆ�AZ'VҮ�e�h]\Bg�L�����/��:>n�u�c=��4��r�uҏ�a���
��o�s�- .�;!d�	e)x�<�g��L�$ÕV��Z�|v��d����]���X5�p�w��R�%um���^^8sy�t�ۆ�\jƣ���G�v�]�b7�%SλB���<�����~�Xr�<��3�s�F��ܻW֕./�J^L��~������}U�����<�4%B������V�>�+4,8�bnN�,2��t<��C��DXTu+b�s�ǧ�i��t��z���}��򠧙. cy��t���m��\�~��U:&���o=���֮hiϨg��i�ɘ(�5��]m� D�|{Q�7�����'g���BV�i�w�yF�Y϶N�=��EE��9{�N�w���}l��^�&c}�v-�,���N�H��v�]�3��nq֙�'�M�R	����āՐӗ�il����R��N[���Pٱ��4+]8�	�;�'�i]�S,����۩z=U�嫝���˥�L(YG��]�>u�M�9�X��h��E��+>��"5��<z@f߄�u���"o�;�&�*y~���z��zmsx�>���������3�Nٯ����F7C�6�hs��Y�� D��l�d]�����2�.o����Թ%��נ;bL�~���U5"����qUD�!-]���]����&7ɷ#����.�����*h2���U�p�T!+�Lu՚n�+=e��m���r�r���|wi^{�v������~̵��#rT$�m^�2��o��*����y?�m��Nx\�ӮcǝK�<ǔ�u�J��Y��{ ��^��f�KIh�O��lFd1�X)�b��Z��T�6�-n�y��Gh��wS�k��s�he�޺����
x�8G:,���ݰ��l�6���κ5b`λ8'/�gT�^��q<�IգM��N�k�_��W��ڦ�M��`�Xa���&���Z���Wڞ�y���K�b�'۹a�>��'^գk%�-��x)���F�MJɇ�_��;'����v7%R�Z�=0iG֑�C���7f��>(ϭ����qϝݍ#X��UdE���{:���{�:��y���?z���}fu�l��\�og|Hug��#���9��Ǐ����k2qۙ�l���>�/ �Y�3��!X<J��h˕cr��u��ڞ�>�N�8���L '-�z�d��7G��[������Mg�֝��~�a��rt:��ΈDo���U�cy�66����.���5׼�S��MO'�8��-8�w�6UnZzQB՞��3ԑw�A�Y���7��P柘�;�R����d����m%'P�kǇb�%�yA%D�'��Vrg>���u_t�w�Rg�Þa���c���;���ɩ�<�������<�*!�,����A�F�l)��긳F�����C��������bѲ�\�Q7�v�ڵ����9�A���J�� �9gX����/�]����	7wЂF�]^�n*�P�,1�l���&��w��Jw:&�E1@Ton��u7��2s��4�)E��a
��f��[}էY�a>��>�դ�xOު��a�{n����4s�^��9_(�"|ʂ~�i��u��i(����첷+8/m�
�W&w-'[�0��nd�*u�<V"Cr�2[$��Z�V\�}5t�g�^��UN�v��H�Y���u��>N�%7�,o<�@�����[̴�3�q}�+�=�����l柒���A��c:R�q`�R"��z��q(�*#T3��o�R5|r��1�K��f���X�hx|D�=�����˵�&y�����,z�_��t�r���w�-W�����ܬ+s���kGGL�3�г���V�Y�a�n�Ӈ��,���;=o��߰��g�Y"��μ��M���ߪ��(a���t&�<K}bz��\.�
@ܞ���7&�g�mW^(zϓ������}'nn_N�J�-�����;�k/<{]0��(��_@V?X}J�>=JE�˸^����M�$����PH^�ǻ��%eeծG`2�x.��R��ژ4~AW�g�\��Yg����N;��V6u��3"�Wm}e%�:33���0�-�s��ov�n�Y�a��%����Ntdu_N���<�	��.�o��s�2t�&�}z��wgUGf����N�s�R:��H��A �	8�fB�ۛ V=uÆn4����uӯ{o�{쵄�����^gB�l?{j����.����%��v������/k�Xv}g��O�q�Y��,)��B�MP��^Ҹ�ݸХP��z�ڰ2�	.S��uD۲�5~W�m\�l�iߋ;���8ܕV]���EtU\��rZ� b\}��6�^��?bg۴,�J/ho"_�qg>���w�Ƽ�ͯ�v�Y��SOg��F^��}���h�)٭ܗ�=ƕ����G���"yS^��^Jf�$��˸\n!=��w!5W���0suO���l�"�wܴ'ZD�ߜ�yl�b�T��7���u3�SRf�w^�,a� �D�8�MB�^k�n�X�R.�9���!1_ fv���p��I�[U��וcB	Z,Q����D��)���mJ��Dvj��@��g^�j ߱L}��}�۩h�I��H�b�w�-`wWH0Q�ߓ��6)8������uo#M|��f��k��Y1*�.~�'yn���t�Y��「
cyį�����_]q��z�#�����ܯ9m3]t�&Y:+�[�#����Uڶ���x�6����|󊽕7h��r}�OtK�T�Pz�N}���֓��eR<�坬�Kh,�U%����xz��2�5.���>rgv��}oT��']��f3u��v���"��	�5�zY2�I^<&�PX�έ�]���8���ѐ��n�� �Ж�pVE��F�kj�=_�~��/��f�~7��\I��!}��OjAѷ�t�Q^�-	m@��.���b����.�Խ�z�Y=a��~CO\��r��P����,Ӛ��]�,+pA��jǾ���^�Q�PX+�%�/�� ��V
G��.u�KUu��$c��i��uO�8[�&�y`XeW�\�b�(�5��اK��o�)`s�멚�^X�².�}[�f�*D��A�3�"�>��O���g6N�<�#�E��j�,w*���c�h|�v���j��T�*�����E�eg�w�o|�g�n@M&@�h�kn�gh�\��������A����MOˆ*jƨl��v��]����u��B�󩞠D7X�����m��%�U2AE�:Ju]ҷ�X�����=�}(�W;�V����E�
����V�ݏ������>����D��WE?#����^K�y�e��o�W՞�a��?l96�%�IA����*��f�웹���tݠ���2�<b�i����G䞶��B��e��Zttn�i"�eG�����:��3�IQ�ђ��ޗ ͎�
�.#��F���s۱��f�[��B�7k���z��&Hge���;�����Y���d+�_�xUD���D�
'�z�ϗ��PC�a��8�Tȼ�W�7q������S�:��?x)Y�X.��%bRo��-W�x�B������v�<1�7]B���u+��4��#>��G�d�(�.�!�r�î��u�N������qgE$�W�w�d˭;{�8��4���-.${�*n6�ġ�M����%�+b^Β*+n�z�Q"�v��O[��CԶ�Fi�JfaM_P�j)N� �ԿD���{sy�����dJWZ���ʏBϬ�Ztmg^���|��I��i�R�aմ�����ԓ���<5Nʯ+�܁����v�R�_ƷU�OT# �XV��y�z8?��S��[�G��׬<`��5����.���H?�Un�c�
�5���º����\����w  ˬi��w�h�w��s>��t�x�vYc���4VJ��_��c�\�r�X�AORʂ���'1�z�:�ٛt��5��P>8�p#�W�<�t�Y��M
ˎ�\5n�R�-�V����d����b%R=|\����U+��2}x�N�5%��!�v��ju�y��.���q�gq���	vv��v>��@vh!wSCO)�Z,�⁪a�{S��׺��Ow6�;}΍�l�K���E`�r��⿷��m2!W��o�]a k�yY���uf�^�=/�xs��X�E���r���q��w�B7XG�gL�M:�����O�W�bo�f���Ԃϐ�8��<�%�D�F%ă����\.��.��L�Xp��G�ݐ���[�R2S�+�\vb�ǈ��u�F	㶹f� �PcACI4�6�긳�������G�$���3^]z�/�W��
W��oLy��L���Q�
��A?X)}��J��e?8u_M�N�Y���;�;���o(tçK�.��vd:
�Hv����Yk�*+������t������aW:�u�0������a��]�U,�{��̛o՛����#>���:�/���q�҂��]'dU���e'}	�C()\;��na����I97k.��3�>r���������8{-}/Y�v�d�<�Âen�&O����]K�����Y��ؑ�
������ZB5�.����fC���	���Fy���M�
�BjsFfݥw�s�	й,��k.��޷W�gH}璎��'X�T���n�yM���\����)�*]��{sm�ۓ�27�)�q�R�o��du�ᣯV)�m�>��g���o5��9�r���8m�&�Z���/��o�~o���YM3>ݙ�t�EL����dmn
����0�u�MH�����Y^��6$��Z��ޱ9X��A��lv�倧G�\ןH�7Gd��%�x�H=]֓��4ޮ��p~�R�]Cb�in_@rz���V�;9w�u��:����^M�IYe�ǋ;S��D�>��k"�����V�ʦ���՞�����~���\küX��&9]t�e���fi!�����1�*���F�P6�Y�XU�`S����A�c����W�i�K�R�+�C��]ŝ�+��*^Y��i+.�pH�RS�[�[��F�I��;3=It�V��D����m^�dV%�fo�;�dx�zJ�+.�w�?T��|	�;rY޽����<]���ѡ���Hتa�qx�r���5�m|(p;heM�μt���g���6�JMxckC\�=
]Nz�>�tB��>���L5gi��0���M^��]ְ�FDGv���%`�O>��eiwܵ�i�~�-�~~t��F3-�ÞmX�<n�e���O��NCU�L�.L��g�ZA�r!�j��a�tD��`��1�N�5M�#o�,Gr��{V*�j��G��*Z���F�k56�O��Ef�����չ��t��Ok�D
��,�)�"�܆ޮC-
�N��!����e�$�%�z�5x�e[�ͤ�$�8��_<�]�͏/�d�Af�mj��FGJ��8y�F�p�07J&3iዻ%۸]"n���j���V�s8�ύhVi�Fu�]�z��9R�8���T^�y�)E�+�.���z�bή� �$�,�B"���\	�E%��fr��$@��N�:�rF����j��E�t�TU�������c�s�:� ����/��d_KVD�/^[�m5{���~=�J��2�n�� Y�pt���/Y�b�\+������
�=AG����b;�R޳׺�
x��'A�o2����%�IH��F�]��9C[��o� C�1��gxj��;8�9��hm���or�R�Am�:���Y}`F�>l峮�j�J]��Q��V�@U�Qt��T��<j���K����~Y���e��X����lK��fm���n�x1ᇻ�\F��*f�ku�
ƫ�K�<̣�S �[m��$2��F����5���\�8,IP�X���,^<YA}N+U|�B�wW.��u�lxF��u*��D|�i�NY�
���\�=�g4"�w����ҫ���wt�0zs[|h�ݮ�ڶi�`��>B�q�&Y��:�k�3�t��ɒ�;�R@Gm	8vГ��k�����x�4d�	K�r�1V��
4)ћ�s%�0�g�\�t+��*�d,��[#BHt-gN�1��Q��v�-W'ښ��Y���A
�9��r�h�b��*$�����g��T�m�Qq
9vJ�P^٧q�wVN�e����y,}�$3��ioyֲ֮i����ϰ��byö���{�y���t�؜�������`��̖sD-ʅg�5
C�=]��Ă|�J֮ofk���'o3�k�\+E,�Qcg8���{Q�"rY��K"�X!ku���M�]K���8�c�p�bN�7L4�{�Uh��d�+���i��sy7�il*�s�����uwh�Aj,��ʘ6eg�fSx#�t����RV�6oU��ң�Eʗi�s�Hab�}�a_ǖf}}���G�L��=V+���qJ��7�fsf%i���2G{���<V%}L�o+�Z�����
q_ϖ줜�w�|ˮ:�&�i�z����ڮ5��7$�7Khn�̜oG1}�X<�࿹|�u�������Y��
ԯz�[<�^�߀������fUҭ�Z�v�&����x˕ۺ���E�I�u��Ŋ�r��:�=ܑÏr�u*�yh�Ʊ�Nx�<�v���]5���R+y������<~��%"	 �"�L�\q(��b�\��԰F�b��(�5j�S9jR�c\³�k)��j�"jʡ���CE�4ᅩZ��c��:��e�+%���Yu�Z�[�ZU��,1U��.J\h̆��EZ��u�\)�-Qj��d��r��-Vڬ۬0ĭ���UT+4�ŋ��WZ��2�Ń+A�s+1-�b"*��
��֫b,�����Z���.8Eab(����PQTQ����6�2�U�����"V�c`5�6�0��īm����PADE����kjV�嫪��#��QUUL����,Q��,����Ucie�DDQ-����)m��U���5�d�*��4U�Es3�jE�Q����luJ�2�Z�q�C�L[h1�#mU�k&�T\jcX�ɤ(�,�tj������U1(�Y�"]dr�Mƈ"����k[����?���|�i��ִmV�T}X�-,_[Imm.�c�HGCV��Ą��RL�39�;�V^+ˇ��,榡�N��;�k��~��J� D���!�
	y�E�`O��"��c,D8�e/���Vڞ)��P[`��j�٫{mQe[�|!�n�����|[������j������0f��&"�򱒽��ƍ�;�fW4Ѯ����{ ��w	�ª�T���Cdë�S�[��o��yk(bUa˄�A�O�q�S/ݗ�s�cZ��c7\��Oy��v����V����
����0=y,2J���lN���iW�W�ٓo#~���WWL��*u��E��4��6������,���'���+�:'���3ɒ�F�{ϔ�]{����Q3�@k�j�\��Q�	��UG��uڍ��UA�:9�/E>�mj�X�V_u_!�8g/y
8$�%�:����«�g��%�=L��"qU�3F���.\��.�n��}ufr�0G��sXB�<�,<*
�M��,5���O��m�wI�����{g�T��^V�֑)��)Ԋh��O��g �;,���	Y��z�V�.�m�4�5w�k9�uLS��m��N��=[��q�5��&�N0�Z��Cd�F�=��� R1+Ɨϼ�ޓX,�{�]b�ir��/���Uk�s��w;�%�Ү�աܧ�h��*�;(KU��}���5Mi4��<�](lY��N��W$���e�3�K6�pʛ�{̊/��]ӖϸO�m�ǆ#�mT��mv����x�e,���C�-W��j�mn*j�Cf��v��������!�p��UCdZ��ީ��Y�L���x���WE"��л�n^��<��A��T��K�*�*]�fߺy�79v+{��A:��"�
%���^�����z�^�M�,��d�!/A�r!��g���c��=ULY�s��Y=H,��)�&ש��c��� sɬ����y�ym�C����:�觊v�s2�)Y���Y%bRi�Z'���4��U�����w���XC���ԃ��L���SL�3%YG�%؄c��u����tB��r��t���-e��Ýx���3�7,B6�{ٖ���č�*cj��)-F�x��'��]fb���.}[y��)m뷃�
�5��iu�߉�j�Ϋ����	B��}���z<�;c�wmaL	Z�֣ޙbv�_�/jâ�l]����3±;��/L��d�~�pQs3U>��+.����݅X#�z.W�����+t���6���ɮu��sma�׆�S�Pʎ�#ܗ��ls��x����oy-u�{#� ���=<��!���u��9p���Q�W[uh4���q�Ԟȳ�&egTV+�B�|�(�5�o�rv�R�_ƷR/T#�S�+pm�(��7�xm\پ���9�js���^�feh�j)}Q�	���ӑ?z��G`�Y�an��˿-@W����j���m�G��*�qݾ'����]=�g�G������x�!�t�F�;��&�,����>¨F�������8v�� �e�]#S���wk������
4p����N�UiZ�,8� �'/�=�E�o;��dB�s�d[.���ɛ��n������a��ŵاu>VpL�QW�u���/����`#՝0f�m:���������=�W�mB���&{�بo,Ե.X�F�K��Vi���8��}�}gjfJV��'S�ʍ��f�i�LϽ���K1^.<E��!�)r���
��CI4��OtW=���Z�|�-ڪ���"�s���{S���d����9K֙��|���AoȺ��8��C�-��3/����8ؠ�_��K�;���yC�çM��L��T��t���z�w�����5h�au��:�Q�WJ��+���y��7(+�ms��w����ׅ4��h���:-�O"i$�]� ��DKm��`�{��W7kcw�	��!ie.X{Bu��U��ұ�cM�vnF|��!�U�8]6�]�g��:������&�%�&:����j�	(z�X�s�nQ#�f�Ǻ��Z��fXְhaSۻ����w����ѕN� �h��r�֡�<΍��y;"���c>N��k��^y�\��Q�vϸ��V7���}/L�����U�9m�x�[��z��'���ܵ���'�5i͇1x+���?+/�P�6�+�W�8�HG����в(�-��>�[���-�+��3y�� ~��^9$����so�N<�F��س3��7S~�	��,J�7_/o7<�c��ܧ�v%�C����f��FjϽ���vY��齟H����Gi/s�;Y��{�[�bM�a�-�QV7�����
T��C"���/~�c
=+Aù�X�c���_nW��c��&|1h��V�ƪ��՞�]��/=k����`����=��o��U:6x��x4��~W��jLf�Z�)K�}n����ih�]��;��Odui�5�B���D�zC<s�*^N�H�U6PHW����ݳs�F�o^f���N5v��2�w�u��� �[�{:9��b����ڷ
��o����_C�^U��s��]i�E�s��v ��]��_V���$�|+7��Ǝl����(�Wn���͘���c^-�#c�o(���̕ǁ}l��7i��j��|�X�^)��H2C�	��˭,�|t�7�Jˡ��zÖ�|E;�s�j2}k�U��r�p��u�<�=��@�y�8B� �%���n`���g��^�g���RcA�e�`�6��D!�w\o�}c�8��KT��0Ds���o���f�O5)�]k���� )��Dܡ���W�@|�b�<wܴ:�"yk��Oُ��\m^��rOԻ�+�aSV$L�!��^�F�o�/�s���W�����K��b�F�߃��x��UY*�!
YE�'�S!v�\A���d%��T����j;�o*1�|�ߌ�(G��H�b��KY�A��Q��b��6��?Psd����^��a�ۄq�����}��X\&�v��C}C��)����Ο��DK��e��`�#�g��;��̠��u�� ϻ�ɗ(2Js�����n��n�y;�2����Yޗ����>�RDg|]�����;��
���7�;�N�Y�W��4]F�s�j�x'���j���]5���cM��+͋�6��Y�f�>!
���i�9���{��:�T<^γj�M��7���Zp)xN Z9s3��G;5��U
��Hk���;ۂ.Ȱ��+��4$�ZY��_^μ�I<f���v(��:&'�	�N�N�.��%����� �~B{)xv��M�b<�X�7U�Sέ��S<=���jǤ�J��(\O����p��W�/����&z�[
���ٯ
�׳��fdR��sXAC���5����RJ	a���ا�ʬ�#bv��al��OI�mx�\�0s���R)�[�>�kŜ'e�׶	Y��f��6�x�utш"��-�X]
�_m؇9�>y�!X�a�u��8v�Y�\֔s�õcKt�AƟ�c�Ձ�P�k+�P\{��B����Û�4+5�1[���]{���#��{@S�b�ȟy�һ>�YI;\M8����U�+F,=
o!�,Cܗ�[>���Z���m�׊��{�wþ�L",dKx������W���5앇�����͞�yq����t�
�W��	,x�J�+��Ɔ�8]E�(�%�OP=D��2+}���un�n�{lP۟V��J������S�:��?yJȆ:�t�IX���Z쪙s�6���h�c���d�Շ�K��'�
�p��t�	��I��=�~󝑐�Tٳup����nN7�u4��e�5ӂF7:��gmJ3\�p����Z�3�ŅwB6��5k�������Dq::ݥibS��.�U�5q����vN;Ƹ�٩���x@V/��HQ�hS��I{��W�pzf	VQ�r]�FX}��Q���f.��G��]K8hW��	Y�{���8�]FB�w��k��F���&�m^�3s~����y���;��l�Y�g��^|a~���/� �]8�s�CM���zfZ�ަ�&��ۥ��5�u��ЩZ�����.�W�ʏ~>����F�g^���|��5�뙢�u��L�w���([Bo��k�cW�4}���UHx�.�[�,��(��|=8b�V�^�iKi�\�Q�^ṷl��]�Ӄ�A���Ve�<xD��q�'D�~�AЮ���1ށ��6���x���Č� ��q=����o�>Sk�������mR��ߏJU����F�]N�F��^_����	�=aq�+�/��452Mt��~�yU.�V���e�G��`	|{ZK��s��f{췀�Q�p%���״���^�+y�66�����"���/=p�7��r'W0+�K�gz\e�3�A�����搭�k��P�5T�J��waW	��4���^��vr����q�] 9kF�H�O8q�w���=|7,;����+k���_n'+J�vi|��-�$��d���,Of������$VXM��a�Z�[����_<�it�q�#o��V�\�ޙ�1]K��.��'��l�����nW�k��45Cy`~��r�D��t
OOqD���6�<:9�o/<�fy��Ōg�S{���x��H�'���k�x>T���|�8o:U�~I')��~F}�h!�8((׾_�y{D�O�#�h�/Zg��V2Q��z9ŀ��y\���1�(i�~t�X3ٶ0�WL�Z�o(t�6�OX�\~� �jZ�}��[Υ��Ғ�H���ioj��@V�R®u���'S����_���7�lr
u�^A��شJ�&Z�j���5�����^|�i�2�x��DR��t���k)���K�PƁ~'�"�w3u��k@�s4L3[hxAH`�����3����r�/{��tm�v��r�� ����R��@n6�+�>���!�Tgxв(�-ԫ�	�nE7�m^�H-gV�,�j�q�;��>�H��:���Lme����UO>(a,܃.�L}~���_�? �b�<Klm�jǮ�7�*3V{���D��\�Ϭ8���`	|��'o"Z)�����9���)�]�E%=�M:�rıH�a�"6������y���͔�T�`�h'R��E�Ê���{�*�;�e��­u�w��U��պf'4��4��-��0_	^Mp/iY[���V��[:�d�[AuՂz�q�sOt�� �k%�<d_Ք<n�4�+�
��>�A�ԡ�_y�uڋ�Z�&rr{��N��C�e���W��ᇵ�r�-)�gg�U{M�z���g���V=�Ƽ�XỖ��Vx�$�4��~W�=�$���J���k�菐���]�A)���*�����γl�,:�
�2䕢\�#㼳�*^XS&�.�vTC6*�r��!�u���U��M^��j���:qY�D�fkN�Y��q��Jt�e0�כ��ٞ�v�Ae���U`$��eF���H_�P�U*�Γ�Ŝ���5�X��oyʿI9�r%^���d
��u�g�E����̶;���-�s����}�\X�����J'��eq���{��� <�v�D������7}�k��^¾��a-m~��~�7�a��{)E� ��� !Wu ;�@Q�i��φ�R�����dWݐO-��rpOP���cXɃ�*U�CD�(�� Gt@�>�k���j�]�����	�8��AFu%�N=�ot��!�L��t�I�q�2.сr��h�0���)At�B�0��ز���e�z1n�B�mgt/�r�o�N�Ll����5�H�[�ԙ�=�l��b����nZ�mB�I˦�zw��'ܳ�W[��錕�P҆��h��eQ���~�-�%�����>��"���'Ք��$�[�V_���[�a�\C>��-g&bU9p��#����}+e�>xyr{y<�Z^�W��0E���\�:�2�(k�g���d��a�S���=\6vmw��c�m���{��f�j��}�4N;E�q��1P]���u����;��
��g���:䀽����5�)�À�{��Q��D���Pū���v�k���Q�{wz���w>����fu�-�}C��ߣ������;��w�%�W�yG}B�C�U����u�aG����K}���z��b�qK���������G5�5KB��^ʂ���B�x�B�($���	q��+���D�͸M��`s���R)�[�>1�,�~�>��CM{�z���w���ZD=QS��j�,��ڣ��d������vC�_vYi�?X�:��% s���it�}�)X4��9	��w*5k�*j����I�\5�1o�S��Q�y+~�u���G�n�7�ғ{�Z���XܔU�8���moZ�f;��9���[�YoU�6��ʱ���K��3�Jr�ڎC3���Ӻ��YX#.){�s�/s��4;/�J�����>����w+�����4��؄ԭ�ヷn�*M��2�J��7�/�q�۠uJk�+�ac{*I��^���h�ޗ��L�=0=S5X�;Z���>[y,�U�n��Xyቛ�Dj;���{C
��$�<��pV���� r�R�v#�O{���h�Mh��]E�o*�	��C�C���ܬ��f¤�rx�X:NF��ʓ�t껫��cAG���+���m�0��ryj�:9�:כ�\*�b�e����CP��r���K;��I��v�r��v���Y]�T$��% R^;��ZJP=4�YW�(8~ЫB����f�Q�f��q
ʾ1�*�>�b���no+���s�rp��J8\�3���n��١o�F4�PM,�T�ss��|��nZ�T��O���4������ai��uO�� n�j��V*���:�ÀR��6�w���������=�ފYs-�NfMY��'6�qSh���㼠�����700�g�[�_��s��Z [�l��ntӖG�]��	�2X�ʊT��W/�w;�vK�V�T*�sú
\�{����)]<���dP��C��rmv�+/���A^R�Mkaj�rprs��[]ȣA^[�ms�0�ݴ��ڧUr�@�ه36]#O�PZ�e�ٯ���k��cEh]c�e[��_v�ե�3��pM(ue)���<�dl�z]C���l�����5+��d��+	{�и��E�.��x�3�nfvgG��>W� ���z��/��#�����ug.r�2�`±N�l��[ZS�M^@z�ن�r�M�YZ^41����{�W�^W:�Lj��5��,#�F�c�o�����&����&3e�/�Sl������?�e��M}�IY0D��sˈ���Z޸�\� ��r�E��O���5%���n�<��bu���S�X�a�K��X�����XY;ۨ%.�9�sn���B;ZhVR���i1F����(|^兒�T�\qp�`�n�s<a��jwY!5:�ݭ�&�ūS
�.��@���o)L��C\}f���ҫ�(wP�7�ǝN���Ѭ��Kx��+�t��{}y��9����ZPͽO�&n��я����۽�S�]�Bq��:ؔ*�L���A�4��o�I.A]܇(#�J���J�qp���O5��ƭ��!����c<{�H+�����o]� ]�iU�]L�-6,^���8x��uVE���kA0���+on	���o�j�>N�RLVc�"pʄG��ö�n^1�;�6�*��h�A�t��w)m̆�u����j�rV
&Q�r�->`5ٚ8�/���u^��<����`bc�S�����uMat�UPE����QGE�
"EMUQEAt�EMc��b�.�8�fH�(�����*�W��(�6�AF:������WWN�\k�QRҺ� �Z�:h��P�`�]Z��bi�Df:q�QunR�9j5�QRڶ�r�YPQDm�WF��e�*"�EQ�b��K���6k+-ƈ�EF&5���jS-b�EFi+m�-u���V ���R�UC)b ����F�Q[l��Xꍥ���"V[aX�T���q(Ōպ�-���F[V"�kn�&6��[iJ��ʅ��Tq�aP��"�+s3.�r���-Tֳ4Ҫ�Ղ��V�WK�f���������keeT��(�"�U)Zc�e+KKQDDTk
V㉊V�Fږ���A��2��ZP�*Uj����Z�*c����.V-[,U��,ˍqLjZJ ���J*(��PO�k��_�f7�a�jΖ��LǮ�<M���dx��=��u��t�+m�psQ�ԶN��tirnsgu��d���*�=�7�s��x�z;ǫHzV��S,��\N8�������Z1a���*�Iz�����ٕ�т��y��*�v
Ϥ�ȷ��EzQ��`X<����9p�\N���I�<���np�*�R���,x��P�r���sª&6QK(�ti�H8��H'(7���WDg�����ˏ��)�
v�̇�
VD�TԊҎ�'�+�p�̓���yg��>Jj�[�P!��H>�.�s��F��EE:$��˜���%7�fJ{�[2ݛחS�]Y������������F�{ٖ��q#rT$�}E%�w�[�i�Yu�YҊ�`~y:�O�㲆(.ǃ-���2�X��~�wiKU�G�f?^��*#�j��P��D���'u֣ޙbv����2֝�ЧT� o
~��q_5����Z�D�P�C'��k>��j�h��g�����^1#ؙm8����̌�c��s`X�[��e��fQ�_9����Ȼ������:�_��L1T�«w|۬���^쳯t���K��֐P�Ɲm
L����#����kR�@��6vp�[T�㎟Q�g�����C{\Q���ω��`L�l�I�B��9d#S.��꼳,<�K�qɍ�=�;�{���EV�S����uA��]�7��h7˭r��r\�sy�V٨�.(v� �=��O���O]����џG�Q,���S%N��y���ݳц��(�-�Y�B%�k�Ũ�����9��h�w;���5.�_ sqL�v���f)ó4�����V��+�� 5\B"r���\5\V7�г¼:��#Me�-;�6šxmGH����yY��E@�=��/.��Vjw_��D=;Y�9v�X�Iʽ�+����T7�z�e��Nj��~K��I 0(c<e�q>���ȗi�(�w�io�������`ήX3~�c��:x�u�F	㶹`�D�WM�i�ޝ�a�@	F^�d��Ve6����V�& �ӽ�}ea���S�v��=��p�â��7B�)e
d2������grНo(tçM��(���u#�ד�)�-w�Lb$u�/�%bD�~�X*��M�$q��A���jrSwMJ�Oe�֚h��|z������ܭ��`H���P�.5�P��o��vEt(�f���`�W�Du�k�oG��_T�����TEw)ˑ�_5|;�{�j����K�/ǁ+N琙=F��Q�4`�5wY{⏱��c�>�ꚍ%uΰΉ�6U�Cr
�qY�]�,����
Y�{l}���`Wa�]�%����&���F��^��%�|��Ս��!���ze�v����5���җ/Yy78�{ }-�=��\���\no�����+8�_JN(��aX�W�-a�L�3�в�';<a�t�;�Kl��y�ĵ�J�9t>�H�o�Vz	����ߪ��"�ՎU;7����i����F���&�"b[{c�� ��5`�L�����}������SZ���S��O�#�$����|U�Y~�C(8N��9��<ua��C�/>��a�u��peӣ[ǧ��7�Jݺ��⼋�G<}\^}u��>�r���_�Y��i����~~�k���R�V�gDVY�=*����gz���0V�y���q�Y��&P������7��&��ۣ�t�X��*Vώy0�B+�SI����N�Db�Ey��={�?W�+Էֿ_Q/��Da澾f�W�E)�	�ކ+G�!�\$ˈ�o�<[Je%�A�'�:�RL��]:У���ۯk�;(�,p���W��K�wqEm�Z��,�6��|��P��k���´���+x��]������d��J��K�	�G�'�[ǨQC1ξݷ9�U�P��z����_f(��<���V���J���nSδg�R=d	�l�t�7��˞�5�ocn+��p��ӌ���t�ٷ��C��<	�PPM��Mp]���A��mZ�� ��7`�TjWS0_`F|r�N�N,�C�����^�Yh�}Y���M�rla��>������S�
�6�ky{V;v*
��F5��Չ D�=B�^k�h�r����V��̞�.�6�f�,��g��¸�_�V5�̘=��^�7�Z,Q��[ύ�Y���-�%uOv��c��޺N�R4�ϵa���c&h�Uu;K��~4v���3�h�W�61"�����Ov9�Z�+O�(�Թ�ńM��f����Lĩʄ�A����;���h�����\�K�ǗPz�9��#��ϙ�[U��P�?�= ���r�$��d���7^�=~r��֗>�t|k���j����le\x��LTg|]�����<_��.���H�es�5�v�P#�wl�}+�5��N�&!�@m�V�~;mp�rV/���߱ng�����󭔲�%�w��!�TS<=B2���-�B<��P�W~��3^�\ W�7WB7��*��Ppy�� .l;V����d�\ZL�r7���:]�:-�H�*j��t=��$au��s��t�C=����xp��F��7�>���d&u�yV+�*�ŽR�b�_�iƻ�^`�e�k�Πc���ԒHo��`�-�d�S����̗��V���B�<��<��-<'���?c�c���;yD�Vb`��ߔ}=�zsԆϮ]�W���6�5��|�tC:�M�i��׋9�vY㮒Bm��,��g/v{��I�+��x]v=ENTX!��0��ɱ�����ǲ��t�w�άk's�pȈQ+�A�ԞM�R�L�_��j��Wk~���0`��<j�7"ox�a�x��AHO��|�ٽ�.��ƴ�ϩ�RN�W_8�F�]�wJ�Xy�̈́�����m<�f�mV=��[�D�;�V	;2-�K�y�\N��~F�_tW@�N�W��ǂ�Z�N�|��U�4C�e�
��k�<l�W��f4�����[�v��,���y�̤���Wt{u��@>�ˎ���O���̇�R�!��]5�-��]���8A]֫R�@>(������ԃE�e>����z^<73�f��:}�M5<�u��+�L�L��zN]���U��\u�*�[�#5��Hk �h������S+n|��-n�̋O�xL�cv�z��{F#O�9��zo4��yG���ƙ���};�}	�iY�_���gwZ<�3�l�Ft,�ۙa�����.�j�6i�_��]Z����[��6>]&��v{L�3'M}Ϧ_k<��� �Ҡ���{����O�㲆(.ǃ-�������+�7�V�C��+�]�-�c2��֡�*7d�Ӻ�Q�(iDP2����|�͋|��\Z6�җ�Zuts�3y�ِ?U�:��{O�:����8��@��aGgm�!fb��[��}�\�oS�����w���Z���o���,����Ӟ��l�/>�F����f�s�2��[��l�Ν��bL�#��=�ߖ\�7��C*yC�U�'U���O}�qy th�S��l/BO�^��0���pa8�@���Ῑ���5��k�/��wp�R��'���K�LVL˟z����xG���-.�����Jvէ��Ms�ǥZxh�*f�-�JȜ�^�ߜ���L�QV]a���#���~��8�����<��Z�d�/�����b�������X����H��.&�+93TW2�:sʎ-޹��#s�i}ڗ���Y`y�|{|��c"����+Dv]_r{��4.�u�#S������o2��Z��{��g��/���0���a���n��R��&ݢ�ti��7�j쥵�k/\R�q2U�_w3���dG��:wA���jzG&��Ռ�o�t'nq�ga�ӆ��G*�AZ�t"�B�fu�&ΒҜ���5�ʾ�ފ��;�H���k�5�^��]S0��ՑK���;ս%��{��g�w%݈�=�ݭ�W�0���j ��S��z�7���>�Ge�����fh�Mw��^x�,k�t:��]�F}\�!ұ�����I��v:M-�^���
��]���h�1�J���U�������-���`2��r]�Zm�-a�_7��� ]z+��i��gxW�ׂ�WU���������ֵB�r�J-
T�jƘ��zVi�ʹ< �a�TИ~�҄����{�z�d>���&y����'b�Ⱥ�/Q�V}u�:���.����N~ԧu��;�[�hYc�m,��t��>�H��m���z	��kpR�OU�B�'�����T� (a�[�X��5a����3��}��鳲��U�6�Y��y$�_{/�d.�̓����8�SQV
�-}���������v��͡��ؠ��ڣ�S��9S�F��������F�ܦ�����e���v�`�N��F;�J��iܶ2ҽ`T�S*�D�U����^Ak� ���r�u�[m3����֒��i:��[wZ�H
���V�y�U��j^˜[��{����\�ic;��ʎpNkg]��8��"SI����f����g��⹎��`��܍(�!��>Ϝ�4��O���u�'�PG@�<����ڧ�,����䌃�����+o��2��X�]_e�)˗�g�q�X�B+�SIX.�tw��ΑTYo�J��)�JF}��謁g���s6���v�ߚw�΃�0��4{l���>�p�$�t Z�u!�*��.��B��Q�k�;><�$��/����ww bX[lΆ����o��ΰ��me�hCT������S����(�;�V�M�F8��yM��g���8k�M�I!�5L���
r� ���z+6\U3�-*_oB���R(�d�<�u_{�4�f
ʝ�F����&|h��iy���᧸��)u�����f�!d�{�2�|�cXɃ��J��oҶ�!��;��:�sr�I�32�,�����Ջh�a�V���ї�P�To��Jo�P�z�~�-w�-l&��q��ff/k��M]�!��,�]�lR������yk>��J��.u^�D}��Ԥ�c�����'�'	�2��Sfr�U�j�ĤY3)ȡ����Ϲ�E%�0:�mVj{[h������4�{:�sꗁ�����[�e�t5a�������d�-:Ԗ�&\���U��Ѹ�H�Fp��7bQI15� ���\ڿ�I��S�@�Դ0E�
+���]fsJ{½Mv2'ƼW��Vk/3Z��x�u�ĕ3݄۔!9e*�+��W��ܣt�\�t��r��ߴo�=�8]����~�������\I�$w�,�k�b*]V�~;5���Vw�VN�����|���/��]\���ס���S<=B2���-���(�u�K�sN�9e�WNWٛ|� ��W ��B������g)j�A�;��P�.�֊�ʾ�f�C/rY�a
�@SC���&{��'W4N�t:!��E6[�>��g|**�t�r����\ݛ��9=�	YȯP�T�֘!�Ta����v�W�;��t��.,�׼�OaV|�����<���rp[ W�9v��`�q6�5�+�ml��ܯe�(����
�}`�����Ⱞ節RN���h���
K�Rvz�7������]�^Q�f�;�9b徔H�s�I�q1:��"�AD���� ��@��)��]�]YS�N����}�^?�;�]̼g�mh�q�R�XkN�}�;dX��8�0��(��(����7����&XFu�bT�ڴ��iU��!���\J��^�C�b����W��cT\�t!l���wt�;.,������Wc{���8��y��PMߋ���L�p{������rǍ��W/ٍp��>�D)�{ݘ��\�G�ҽ�l(B|U�!����\��S�觊v�̇�R�!��[��i_��F%;7©���.�h�%�
�d_�r�w�.�_9|T���bݵp9��[���,p�٭ׅx��j�X�;_��V�wp�~
�ݷ��᳾�SC��uGC��H�( �7����#����y����Ὤ�ڭ��vi��`ϊ�(=�c������f�2w��O��-`0�E}�lN�G%(��Bw���b��_��u3��<�)�T�ϝ痊�������P~Cz��OV5xh�7���G�c�f������r��ޝ]W�.�E��^�y@n}o��7����X����.3bgT]����W�-S�ie8�l�/r�/�/]�]���xe3�Hv�5�<��擪�ds>��g��3L;=~Sf�`��ƆNT���X�W�<�5}���n�����~��$ I?���$��H@����$�$�	'��$ I?�	!I��$�	'��$ I?�H@��	!I��B����$��$ I,	!I�H@�hB��@�$����$��$�	'��$ I?�	!I���$���
�2��ƺA�	��������>������{�� T�(��D��Q5�[`�R)@�UJ�AIEZʩi�"*%J����}Ǖ{6�VZ�6�MNV�ѻv��m�bѩMZK2��V��e�Y�l�͙*��Y�Zͦ�$�B��n���+MTemh�&�V����e��icM�cb��F��T���*-)[jEl��ڵ�[`�}��Lf۰�  =� ��mF������N�j���0Z�e
���v��9���t���KVY�������զ  ��mÊ�C�@�8�hwj\�P����6����ln�
�:+j-�'MT��� vx����iL��vP:�ݜ�uȳ[
��v��`Pt����hwkQX��j�5�i�� ��yf�&u�'C�0��Pݮ: � P;޽� �P s��    (w�{�� �  z�^�7w:,n���JA��K[f�x 7{z��v�v�]�9i��Ƶ�m+\�֮�ݝ[��ܮwc���������N�WVܝ�N�ݸ����ݸs];��R����Kf�m� ��k�]j���jewm�pڤPv�wv�CRmշ]k����v��nˬwd��ۗ�UB���j�wg]�˩۩]N���m�f�MKR��W� �W^��Q[�sP�+p�3�:e���T�N���sn���Zi-UZ���'m�jv\�v����`��t���ё[Im[f�� ��[h��ݝ�7kmki��Z��m�˧kT�wk����Z�u����j�������u��Յ�.�]\��6�k6T�6Z�x 7�G�'n��k�M�]���U
['wTF��t���s���1�4�;�(攣��ҵSQ`��� g��.��ڰ6����P����sv�ۀ
�6�A�#�:��	��    "`aR�I �h �  ��0�IR4 �M2bh )��US�  L  L	�)�CIR����� �44aA	�&Mɪ~�FQ�4�'����I&b�U ��  ��8����T��[�ê����oz�|-1�bqƘua�'+lAA1�4G���� �
t���� ���  �������44�g�"�h	�D`E����B1
�A/Ý���k5c��0A!ol	����T��ꉃ����w2�$WO)��
�K�M/�0+�/I'dq;��Rfm1[�SsU�y*V�Q"���&�C*S�u���k.�^:Յd��ZN�e�֬��ܠe��=(:P5Iwv
�I���*��X+*��c�C�5
`Ы9{iD��j'��`��mf,�;D���;��>ͮ����s�����X�5:��ٖ��ٗ�V���B!�lK*n����K
�@˷����wx՛Lu4D�����$��Az�h�:�^ə7-f�H�[+J"��X��Q�{%jOP`k�cq���%7/)�9p��Z�`r����k*`�w+6�g��W1J�c�N�ơֵ�L���TY�0ejKM}m肆*Djn=�Vl�Y"�z\JܚfPH(�[?B+�ᴎb#V�dE)�i�Ҷ�P�QJZ��XEͷH��q���i�r��7����b�ڽ�C�Y�6�*|ebx�ИS�ԣ�UЄ���v�il�e�y�5j쥐�Im⚶ �gfHöeA1д�"Y���Ci���**�,�kw��M��E5Y �)챣4V���]�W!:���X(6K�3͆]�Vi+�%���/H$ѫE �lփ��yW��v�����`�V&��V�˽�G�ȡ���f]f37�e��Z�&�tA9��Y��Ř/Mif�`����p�ώ�I%+U��U:��o%�`�gu�N��2�� �kR�t�����5�
Z��&�Zk%Y�i�wN�9���؞�l���ef��V����ګ�^�y4}a�eV*,Pbr(�V�5-!'JֽK1V�^�PR˶r�c�Z#�6�?��l��5�H��N=l%]ԕ�V�H{�7M�J/p��R�'QwWZ����$���sBͧ�����������5L�2V12���vDD��72�U#z~-X��ߵ��tb*�1�Gc,n���7\���:l��:�8B�7	�w�!��:3t�wyPk�%�-e6��'yK`�r��X�^˫OX
V'#�����7A�N+�i��m��Ѷ�4�JT��$m�P���`��L\E/U�7�4P�0d���JҚ�5}3&�u7GB���cm`cQV�x�U 0@+$�i?���(,�1�[u���J�n+��pڳ2�[ʟ:v%ɒ�z%n2�YˢM�1k$kO*A*���V�4,[K/�v�"��QZ62�f0�5m틥�Tb�`꺖��ƅ�M9n��p1/�:X��t"P=�B��^S�������
�7B��S�d6N�z�m��G��l��02A�j�q^SG.n�-֍r
 ����-B��}��q�P�٥%�n�c�#W���9�JT-pܒ�D��^ӭ6����:��6���ѨV�X�3�e�U�3E�V�wl�	��eE`f\�����Ԏ������W����V�䂍 !����A}i���WsT�e��=�-2ҷ�����I�ڍ�� ii@�>�k]��u�X/LQs0*��������V���I�3%Et>���a�pU�Ԋ��^���ީ�g��Ī�w���2lnA�[�zt�%+W����1�jْ*�4�j�M�����4�.SYz�����.�T�G���*Ƥ��,��e|�p����j���+E!��Y.:������H�YClTۥY�-
=[�h7i����ժM;c6�F@�b�,� 
h��4�t����㱴+&}���a�b�i;�%��F��K1�J�S�FQ�4m[��D�-8����-�
�R��N�̣af �b�Fڕ6���l<�m�j����.���)�9��43Kp�f�L��`y��f��x�N�"mez�������7�j��vf�\�M�a��,��f巻�蔎ô�tpX���ݗ[���2�ٍ���za�r����(,��)���t�5����ot��B�S8X�M �T�+��i�rnE����N�/%"a,+U��ڙ-�;T�\o�[�XZ�jkŭX?� �ZJ,�%aT�
�`������/��MˏhФF�E���Ǉ6���G�I��Pq���j�kn]����Z�n�hI���,T4�rj|���j������i�wFl�TrhU����-\v&�u�8����+y�Qv��'$�m⧠�H� �7.�Y.�*�Ê`�b*��r� �-a�{��@0
�41�6]bO%�!��g)�a],4˚ɺ6��G�]^���r6�X�r�#Y$�@�#F�C^V�n��FM����h��֦(YH�֪y�	��̽�0�kj;JQw��XKv�- ٬u6�GM�ܒ`v���YPJ�����J��Ռr�iU{*��f-&�oa2��7bkLV<{�孬�ε*�[-�5�6���KY�Zۑ�[�2�5浚S_N�ok��&�Գu��a�WrZa���0i��jΝv6-�yLU엘�w�D�n�&/UZ��֧ڤ��ģ�!�+q�fS�P�U�i򖉒;��jWx�<�eӶ���1�!��L�A�2���h����cv�9���Y�iU���2���N�A��'�Ä&�6�n���ͧ5��AJ��/i<��ô-G(�K�i� L��N�h�:2����u�&��et�Y�� s0f��Ÿ���,�$���e�sw�q���(�a��Y8��a���\�B���"�C��<�"�)+KB��XO �T�m��"�S'�Z�sV�BۍV�rk"��͎�!��#�@�;p:�G!8�4�8��kw	
��� �����I��j�n1���)l��W"6�L�$�,ie��דͶ��ckF�lJR(�=��k�Q�toV�,V��.��"2������Ja2R�^nɚ��U�H|�l�RB���U'�V���m�.ST#�`2�+n{�u�ݭA��+m=�Mn��
�O
��([yG�)���DwE�\��
��R�wi��My&�ڴ31�j�U���q�dA'�m���^<mb:e��r�u�nR�Jm�pl$A�(e�JŤHV��U�cӻZ��,S��y��y��V���L˺�%-{SS���d��Ve���+1n�p�Gl�@��E,anYmc#�:wP�,eX�$݁P���106ʴ��<s�{F�KcL�^��*�s�-n���v��*����0&D�[���StԔ��� H����F��NV����X7m�#zkr,��A;T�Yy<��]�5zb��&�&u�.me��l��EZ�y���l�7x���ޜOn+c	Ǒ汚ۣtr,�-��]2[���X&��U�`�X%��^^��fLxov�0F��3��ʐH�k�.\��6�a-�u �&`�t���圐��++!�൉a���9$6�Ř���O�s6`q9u(	*�è^f׎^�Y��	֜"4e]!qe+X�%���*<7x�Ifn�QT��M8��yR�MU�1�;�i^�ET0V1tlS���f*W
i�0RhSYyL�y�w�*��oi��䕂\f��Od�4�4P݌֨�	�]H�b�1�T����������ے�H��Uhmk��6��AؓVɐMЮ��5,�W�Ap]7*��`mևT�n��ur�3$j����Y�<��
�AV�n��@m�s��)�� I	�<l/��μ���(�X��Ŗ���KAU��Z�$Ҹ��e�pInh3@�F�#�0�
�i�BJw��%�8����(Ų�V�(v�Hݖf�5-�6�V�:B����HV�v��z�ZԴg��5r۵�.\S�1�YL��X+�q�;�����i�d.�����;�[�R��g	;��)̤�۹�J�E&;��hAX]C�ohM{0'��Mꨲi��묖wdj�5Ni��C=�-������"���`�Fs �� e�
�^�SB�- ݇��c+Q��邓�`�MW�r���y�e��gv��{�DJe25�xX	$��3D�u+m�u��΀aw�(�ڷY�^�#;���
�D�V��6��K�.��HX���f\�Ɉ��Gn�FVVLw�<X���-ࡡn��B
[[*Exv�]�������N�U����ej(0�	'�d��l����C̋`z-��V�չ�-\E�ĥj�]Y1���ڹ��;�ݙG��*(c��57�&�J����Q0װҡ>)\�-�r
��<�2�L5�e��L�4�OPLZz3%�S���oɊ��5���K,ڔ�,h-}n`�g9�f�%vV��D��\�Z�����7XY��K	��)n�T (�1�� ��VG	Î�V�`��G,;��X��M�:Ylս	9{)��D��)&i��*h�������TJ3(J����[�37T+Y�n�lʱ��q�.�
s6���E��-*�)Tiy�Q��$���Al��d���w
No,d� n�ה����iBU��k�9t� B1c5`��,��XqV;�H�����'��zq�bE[v�P���G9�%b;�kŀߺ��t�����YRc�"FK%v��3�kd��t�ԺM��[������F��Bѱf�X������-҉�ր��by�c���q�Iܬ*�$�;��H��D��^L�[�:T�ҥ�k*1���BTI
W���p
�&�Zf����܊, e��z`�%����:xRyc*[;���Em�`���Q���ܤ�b��$�ܬ*h�LlZ�q��Y�x.��Ia7�U<&*f�eCu$i��k
�UԬ�Y�4������6XA4m'i�'����[!CcN��ͨ'I��H@��Z��:�n`���2m-��̪"X�����+�L��4��Ui&�f�Qc�^�*�8(����H�n�7ۊ쥗��3u1M�FGAY�2j*�ҕ�<�� �4����������r�ʏwF*�BMBnj'I�UFB�[F�4�J�b����aL��P��L_��G����FF�E^f���~��֊It����܊J��Lr�Ĭ��S��SyU�)`Ȏk�7zWl�,�A�rS���g�p²mL�	�dM$�+�3V:8\�'8-�]h9�S�#�����F��-]wGS�i����c��N"�c�d\F�^��I��lP@e竐w2[J����e����ukk�����J(����ukf�'*䥤sD@ޞ��ڭ8�O&�<�XY����.�%C�v�ox�ʘ�����e
���f�0�]`���쮝p�LoT�.fCX��a��sG:�҆�V&E]�yj�5�9b�*��d�`.��{z�L���b���9x�V��|���E>�S{��an�d7,���u���<����{��2f�w6)9�f�4���ւ;���s����so�j��T�`>��YnK3��d���X����gz=��A)���Z�q2x:�٪���ֈ�n�AÁ�;�!�в������\*�'ݩ�r�/&ܕ�I�-��5�����ȰTƈ}�R�EJ�١�L�a
�LXӡ����K#���T�윛v�:����ڻL�ҡ�v%�P�oGqxi������D)w�0��)jOki��L�b]Zڈs�ۘ4�a4O�n�!�M�v-j� ��*�Q�4f�f�C7o���:�7Vu��
�q�]��,��+FV�N����ؠ-7����y��1X�*��|r�ib��w)�[n���P���*8��k+x�X.�Pf�� �C��Q��sT�T�Sa�"�Y�{q+W�Xa�)W,��ľ#v�@9���z��F��_�98����Y��^��{(ĥF����G]����-���O�՜�����$�gw����49+��W�һ���/�-�o�BD{ M]��V��f�ꃁ	5���/�s�!Yz�QK~��z0����L�H
�ُ�Pw$wqskM�c�aܵ���dݤ���R�^̛�UU��q' >z���nmf�IJܣû�>�٠`4e�Ti+���m���*+tի��됤)�ci,(F,fq����0�,��l5m�8�B�c2�q]�34��J�E��<>���%gVqܚ���@�j�]*MD҉��[��w���J��hk1���$m-�*� ��t�H+ln#���
�xATeB����K��C�9\�[���C�҄lIyEp�������i�B�݃6�E���5OCJf�]�)Ǆ�w2����ia�1Z�T:Yx!�]��w�`����I��;�2IW\�Ԫ,O:�3M�R�y�(;�";�6��wi`����s9�vBV������)��6�եb�neE�6����6�R�kS�ʖq�9����Ze�n��#�qJ�׍ۭ���lY������e_n+��1<(�n�:HvJ�jKgqb��A�)/�b�ƵTH�,�gz�ItH��27��Ն^gegX����1M���yR��j;��=Y�r�:�C8��xS�1�aW���p<�n��$����c��#@���Bkݠ�L���3Q�*�S�]��5J�����rh��k{Gץ�B�Z�=e&��,p����_eB��w�Ue�6��]��K��X��e����Ԍ��P�t�p����:�>Tz�.���� �C�h]�by����;y��:š]���RG)�
����I�ס����urN��˷����wn�(Y�w}p���b�U*.ԫf���lm�㣕�t�J�h��Tn��nl}�F���d���x�74�����+ɝڋ8�Żݝ�7k
�YׯjR�|���6k�P�@/jaWY��.�86�`z�/8�OD����m�.�٘��"�*���<��ø��u25�.*��;<��3�RB�]s�c�2�z���P�o����:m�ä��է>9�E|��:�V6f���bk�w$�v�CIv�Jؒ���U��Q:^T���o�m�Փ��e��,y��Mb3-(�d���>���5�S�����gLcp�`KF\w:/][|Z�lښ�����궁e�D�F�
�71I"weYٰ�v�p��ͱ1�p����%ӚlN���JYE�.�c�wm�b�rV%w$N��M��S�u��sqrS� �b�XL���.�5��ܱ�G�y������35b��"���3�Kĵ����8���U����Q���7"��o��aQ���Ȅ���{�� 5�HdA�{�������V���y�Z���f�"�	��
*
�Mz��W0����(����^ߌ�������r�zcN� J�%���D�E��D&���5ܹ����ӶF���i�a�(	�:Ρ��#�Q��W|�[%�3��OV�8Ā�X�g���=ͻי�t����Rw&)(ٻU� ��{R��kɫ��r�Gi_[��۠����5���;� vF3/L��7�����{{�m�fgEz�u�	QMV�����M&��R�.o*X՟A��;;�QC5���u�j%0�`
�%�+A��Qْ�}���6B�O�k�iG9�����z����n�R=MK]��D�@^�²Z@N�����PjfЧY�*�o&K�,̠����i(�I/�ϐw)	I]���Y�W[�e������1 ,�+�+Q�K[\O���3Lv�
�)��e�
����|gڷ�R|������ǝCKt'"+
�9���"3F�(��}���Y��&:�kSRl����z̴�ҍ�ֶI��<�"�I�v{[�a�5o����2s�|`�!�-���_]ڝO�5Q�١yȍ��f�1|#۩��խ�W[3x���{��B���6]y0vfQwe�V�kW�L�
]f�iDd�ꝢGX0�4֔(�������\�h �i}�2��h]�̥��{�/�ʣ9�2BD�nN���
!��n�L,�jZ9osiY������jв!v�-��r"�ma�(�Sjذe�|)ܲ��Kyc�V��&I�����i�����<b�W{Q�=�S� Y0��Bl�����m��]M��,��7�B�9� �sU���ꗄÛmT[�u\h@��������� �~b��<Ҳ�:�3���'wF�fs|y�R'�T�"z@3:TN��#bG\��ps���}-��7����K�����`�
��T͚я(��Xv�%������r�c2=�LP�+�J��4���D�bxH�1GR։+2�qPѽ:[��9�R�&��n��w_<�vL*���
d���@R�(���.	���� 7@�=ք8���ϰ)S�GL˨m^s�Vȭ��\�zxRk�IK�#ǆ��J�n�4ҵH�5�Zw��{ID��%(ڿe��e��$
4��rűu�)gA��}�)�䔷!���|S[v��8婚�yza��_4�<י�n�	�fB%�;�2�N}����1�B�F�+*qK.A�q�C+_o'Vn�����p ��Å��J�Rq=سF�F��3�9F�lWZgN��a˧�1V�K��	����AZ���i�x֔EnY13ή��vѲ��v5[�%:��y��<X�G1�\�m��ֲG�ݡ�/ �1=b��˨�7��";;�5w�Kn�v��xGevb�h�N����5&��)�DM��$g���=���ͤ:����tŶ�$�a�;1���(�S(t�0�ɼۜ�e�D�@E&�]I��NM��e}�n96��vwh�X�m��R���N�����]�����j��^^�v@��^͊�9y�ɰ�L�+ �v�y��:T2V�ڑ� 5 KT�N̊�˽�p�PX}u*��4D-ˢ�쭫!�ǋ0j�1q��`:���+�I"Mث�����@�UoC��w��r�E�&�=���Kxw#� I;�	|l	�V��t�7h쨺��u;��>:�`:ST);}�y��c��=���KYg�sdsS�E�ޫ�=DW<�7��E;N�g�c]s<�l���5�ؼ�+0�s^(N1��/��m��xS��tH���Ϋ�����&*�W��|���G_��������}�T��@�����޻GO �Q�j�Ym��ר;�m�ܯ{����Txu+��-���V�`�$��˖����>f·v��|�8��2)s9�V����O9�Xʺ�gO[
��jV�x:�Ku�ס���	{�Z��γ(�F��	-�T�[��y]�G��+I
̔\W�@.�ԼE3$Ы���t����1����bEKy��N.�\X���T8�+fi���1���X��r9��{Y�858F�27Hl⦝�n�5��H:}2�.�ӌ	µY2��.�8���:m �z6�ΗՍQA��4�q#"�[��]��8�z.�5g�C�-��ѝ�y'�Rd`�d^��w�8�r�5ϑ��:��c��,k���fbQC��̬²�PɄ:�&n�͛�ű��}n:M�(��C&1w)5$w�U*͇&:�X�6[��G^���β����V�9��J!ظ�Φ����;�Q���F��o����� au��_
rxm�pN�9�:l�"&�˶X�nhyU3��Hl9�"���BBv�t� Y�^��	�1�9�$]����kyP�W8G-&�1��j.�<R�fw��hZ[H�T��ڎSxL��N��p��Tũ�3K��nT�&N�S��B�@�f�u���ޮ�����ƧJ$�S�9�P�X�Ώ��2�p�"���cS[��ս׎N���r k9��*$�؝۾�(Vw^�rY����-Ӝ�:L3uB�	]0Nl�կ#׎�:�4�b��t��Qt3sfwr��[MWs�!�l��ӷhe�.w9:�_f�1�GC8
خ��@��#uۃ��"̫��+��]:�� ������p�n�If*H�EJ�����|�j�����nK���ޥM�k3�!��)������[9�ڪA�합�Z�T;�9���fN��s�.ۭ����:�z��62��#+�9F6/Z����6��h/�NySE����ךA�靔AMW�D@�8���ES�0r��I��l�۪��Z^-}37��n�+���/d�K2�G��Em��[��eT�]nS��X���W��y ��J�/@��Vn9w;)c]
ju�1%�9Vɣa���k���`iCK�ڶo�ױz�e�WY�+��+��8Gpد��mq�3���˫�ց��N|���Fv<�/l*�{ܩu�҉����!MJ�PI�P�t�<�#XR¹�sN5O�^c���nQ'9q�©ml�"5��	��c���rw�ၛ{�&�I�b��7 �*��u<`��Y.�R���%�}�mu�:���W&lʽ�2(.%�J^�\�x�E��U��k3��=D�'iX�Yoث)�@9A�k���IE�H�(Υ���lS
����K�sdV5]N�Vθo���N�]�C{1䎵5E���J���Y7S��1����9+���.�K/Z֘ٶ��e�@1�rk�@��*�S=[����:ᴒ��#m nTtw7��\RΗ��'_8���RX��Ϋ�����һU��ī�*�n�]F\W0�6�����r�p��Ai��U�uJ��<B����d�ieD������)V�`�&ueI�'�k4��Ёd��:����M=�딕�#����]�9��0�c��o�y�5�>3�u@,���ӣ��u����rN�K��7�*�8���zt [�)uC�-�ͷӕXW{i졁
�@ћ�P�Q��w�����̺�m�0�|&heQ]���S*ɘk��~��f����}���q���+��ߥg'F�� �D�C�oNu:&�V6�x����hw�8Ս�|EՊr�AQ�$�ޚ9=Ϸ�H�h%22�Q��ݵ�Z`<�э7�k6黒�Jee�)⸲��n.�Q�vց�����1��#��\u�ʔ��YާQ�:T����J�N*'+�ޤ�T�F`�9�~��_v
�3�5z+"��wNu���i�{Z��9�V�Z������ލ{���[z2�dG?��ټ�Ar�l��Wr���gI��1�}Z�����u���p�j�񥒦�ǘy}���U�Ok�BL���S�R�	�]fo�+7+V�BȧF�n��)�
����ܬ6��@����`���l�W�V��U��h��/c˲L:�X"�a\��Z)2���Kg�b��gN��3� Xa̫�vK�t�["&���nR�E����d�������Ev@fd��(1��7E�eN	M<�h�J\d�]f�%�2�	8:ӭ�^��CR����v�(��b���e�Ñ%Z��mS�L�N��X)�
�aW��`�X*lR)_c`1�C�����

��Z��f��}r�����j��I�{��h��4٬�� �y���E�Zx�k��B��g��r�o�b
r�ފ��f�d���pQ�*��R�tӰV��2�Av��'��'qhk��+E�M=����Q)G�,���tX/&�n�����˲.v�x	�v�NX��lX�-�*h�˓�â�l����,����]��d6���#�X����^�G�֥��c]wO[�g������fqQ!t� 4�i�W�m��N�m�5u�u)B^K��`�T�ٜ��U�P�"�G+ڊcݙ5'�����xK{��v���c��	���L�Cl�N٫��t=p�@-MC���>���L����V[���{H�n�Az�,�b�J�CR�Mi�L�-�sUq�u�c�"�R�U+�6s���r�2�^Jl��f�oU�.�Z��T����2V�,�Q�;wg4�4��!��!&�����&I) �����հ�����u��6
����[ysab��=�RVpŚZ���hpQ�ʮN�Ͱx��T�s�T��\�Ү�S��e�*�3Sh4���;9��=F�yz�v�wfri��f]@Z��'q3z����e l�����Y�X�.���ե�qm���}���kB�b���i�n@��(�\ �TR.�ˬ��N��͏wwK�6�%�ge1�p6_��[��X;�D��s� ��9��͞����m�j�1@|8���E�z�ۗZ��ӎh�J���oIk�wb+V�bES^NU�!$�Uܬ\���J�-�s]FVJ/\�rWS���un+ �u8lW;���xu�T��k�4s�N/���j櫣��]-p��n��$����ZA)R�}V���O ��Z�Wh���Z�2�y]AV�.N����9t��mU�n��a�xm���K�l*!Z�Y=�ٔ�:Vn�;�"Z|�-��L��Nva���f.@�B�y�=;�WhV�&���4դ&,{��3^㲢�,<A�������ֽ�X(r�V�|O<��q��
a�ާD��R�c:���΅0�+]��J7&��66h��05�m8�,��R:�z�����D��B���z)�uKF���a�h��Y�n����.j��<ɒ�"5-��Z�ww+J�-8���B��7��*#k:���������F\�X��*��X�sT*�`���|�z��}��볓j��f��c����S�\ �کv@�[���VV�ُw�l)��\��e-	�G�rΔ:�˹�Q�ź�y8@�)�c�u��
y�����_�"�h�ۗ*Ѯ�9�3�2{u���O���nՉ3���G7���������H���L�A��湧�]�.��4-V�k���aʏ��O7�A���7I_L��)�H��b��i���"t�E�ՃB����}�C��P9 ���<D��.ۭ91��).�ќ�rN��Z�Qo+2�pP.u;�c5�8&�]X�&P��Q-�=�;�b���㢐"ާ�A,V�K�V�쾏`��FU��y�f\ 0@��Z�����X�i5���j�D�^P�v�Z|ngƠ�S�b�i�۫jqRTru��ܘ/ ]H�raj�h%��>7s����c�Z%k�F��[�&�*v�l'j�%O	�B�6U��-�V�5j26����8��lתV9�`��+"��%���;��u�]Nfí�C�G�a8�@U�:�u�o��j�E�ؓ��T3N�����If��Y.�]CG;�5%�Q�M%�d�o�@�q��b��v��K�V�C1lk��A"j�.*���;
h�ݮ���'7s2�����hV1�O�H-h����f��C �Դ8,\�Ħ�lnJKC��� Xd�8qF�N*u�JN�u�k�|��ds^��6T}tnE�hۥ���on&�.|Tp#����s3mvli9s�W��=ä23�9O-JΨ�vV���4�-u�jН�Z���|+ְ��]�H�J�k�^psyv��\i�N�r�,�Ã7�ItT�k�#����ze"	��B��Ǎf��:���G��8SJ��� ��>;ԃ��������FN؎�,˗.�[�iV��*' �ӗx�m��C���%�����oj��m��
�7L��S�:�h�T����U�B �s���H��._�ᦸ �|�7u��+k��|���`r[�nŐ���t+vd��尶y3���x�;�@�p�L�Y�Mt�b`�%� ؾ�.y5�t��쫒},oF+6�)_e;f��Z��P�]ܵy�^�/���;��i�NY�9j�O+c��N/��%��1�HiN��R��\�k�LI�r�.倖I��Vw3i���&�uv�(�l���������3�����V���/�f-�[+E��֪kr��]����K�@NgX��bn�\9�RS-�ިvQ�`<����u���1�F�F�[cx�'ge�AjrNb"��:����6&����s&i��
Ty´��/2���������TPȫ4��3��̾v4�5�K7t���nE��*�����*�SM��w\����}ZX��-��}�S �B�q��kY9x��G��pu�V!'��ͣ�Wsn���u�(XC�
#��Y���4 M�ɀQR�,OK�Qn)-���v`}Ww ��ER�,�Z�����;w�&�gb��\�h�Wid �
��U�:xnc=�
�v�ۉ�B���E�P�n����س8Gƥ��s���\:�]��v4��j��'|�K׮f��YP.�W�]3�7���/(�o$5C�j�U���Y���I<�H�m�ZW�t2dr��IT�s�x�gZX�z�t�PlB��C�͗��,�J�3_H��LTT�
���eKr+_5b�7Y�h�4�g+xu15�g6�IMӝ��AW.�+&gu-[@�m��M�v#�VZtA;��/�NڇFC2i�`��D������:���8��_ܩ_B� f[]�����Ы襮��o*������	�,5�;l_"T!�	��˻҂�ZKA*`��Ip��By���|
sX��h�M��e:�Ȗ#ˑ����2����OZf��]L�ҙ�n�@�I@�F�q������ܼ��5I'8W#5����>kM䔺-V��gεd5�]L��]\�FP�7�kz�2���������`����YF;�dg0���v7�v7(�l�����S�,}Z�+⛒�ß.�Wc.]Ja;��i|�X:�zU������ԥ�\53c�n�Gj�Z��N3�5i��x�_�6OU�i�vj�;+�(W=<�X7L��v����|�}�&E
�����o
 7��M)��c@�U��5׹H�]|�����͊�K�K�XpY��#["QR�۹�`lL�t�6�v�AS�CWz(CSfCBZ����s�~�XU�&���(
1hꬰ&���n}��E%���-�}��X%�a[��JЧ�O���ִ��i�t��D�Y|���ֱ��f>�X"�#r�|���4x#����O���pـu�-���15�s���a�;K,��1f�WC���%�<ʎ���m��ؠ��g>���m��p�3���	��չ�='��
���&����\�揱~M����]VL���N��2����f�a��<F�:+?@벺��.���0�M|
�.i-��e̭K��+T^B��
�p��0�I��v�t�ǚ�2���ۡ]��{osH "aX���iCXV�M'\ܥz4[2�z7x1�bvE�}%sE&� ��-r�9�37�N
w��^f�j�m+䯶���|��;��]�9Cm
��5�'gݡƟq��`�KИ�S��:���r-����s5�f� a��Q�'D���[2\�. v�����K����6b�:obD��폻Y��Cl[2���� �u&�D�MD�9���'�Dn�D� �!|�Z�k9�9�X�V^-�7:ޭ�&
v�WO��Ъ�9xT�I�涬2����B��:��ri-����ɓ�C|��f�l��z��]�ӈ:F�k�Q�iS�q�^�V�mo)�vwfk��q��d�.����p=����H�[�u톕t����ZR�����+I�:h�Z���h5��QTb����
EV(*��T��h���PUAVb�FF
�6+"��UJՌD�**Ƞe�E��#n���Z"-��TU�H��%�UYD*���Ĵ*�TU��cL�*�Q�*�KZ�*�G�*ŭX,Eb0Q���b��V�QeJ*�P�����+mb�Q��U�*�uKQ��"(�"�QX��E�EKj� �E1��[Z�*�	������V�Q`�QAUH�PDTH���*(�(��QAG,*���1F"�

VQ" �Ȣ�J���X��q-�J��1�)��U`(B�o��G��xv#��s�R����(�Lgb��m�^�GB]E!ͧ���f�c���=[��3辤��[��W�j�����y:"r��!��pqyRE+'�{"�k��kn���y�^��Ig���psT8�Ĺ���ޥXv��ݬ�a��D�j#5H\�)2u�����p̈́���3&������l2���f�pΌe��PT5Uz{�����Y]�F���޴�E��n5=��k$��eLN��ņ�	M��E���y�^4_��p��FB7�>�r��)�����"H{�^�ȶ��ca���"r�pI���	,�L���"FvQv9�V�=��� �tൠ��V\&f��T.O7J��yʳ�o�ɓKy󭿜I�V�L��(��j����ьp�ʺ��h��zɐ��I�V�N�c����VL6r8-���7Zw�9Ԟ�t�G9fG���])wx\F�c���e���`i��wI]02�	�k��=s.�[���z�J�j��M�
� ���#���3.��`�4��W�s5�U�ah�P�\�&E��f8���)��&���҅s�'W��ǫа~N�ٙ��}�x�q��Fm�a���aҊ�ܼ/�^s@�����u���2/��W|���]G�}y�P��@�v��L.b��*'6�l�Pz�"���{Ⱥ\sme�X+O�$�b�*pʹ��i
���SۉL���G96���<��0�l�N⑓S�"�jc���=M�G~��k=i�=����ۛ��vF1%f:{��z�o�V
Zuz�j_1ͪR�#"���)�9-cކ�5���n�u�N�e�Q�Y��E��-@��<�2�8�56S���ϰ��fE��	J�!s�7F��l,�/\�4��n�c���7�!�k�}b���4^.�`��#^V�����jK9�e$L��p�e7�(��5��d���&�R�S�Մ�`�p]X�53�+�E���[ױOnw���Ln>��5|��a.(ώȟ��v]\Z��؀�J�u+�U��m*�*��;�T��잽=�^��*�6!+���vT;ηoC+J�(t�c�1e�Vc�f�$��t�ew7��úg����U��F�7ʍ�R��yZZRw��ɬz��������I)ކ�FO��ڐ��Lr��Y<t0��]�J8ju��
��o���iy)A���miI3^ ��Yڌ_uy��E:�+=2�����k���K	�k0�޸&���fqà8�6���U�][���M����r�H��z��] �|���0Q{Z���X��Y�E�MQ�Ii�dM�@L���U��P�;�c��a���ŷ�$�.8�J��ǧq%��y�f�S�7C��p/1�C��\hd=��)[�q}�,��B����XS�����Fw �D�u��#����m�8%���y�k��YF�@�#��X��-I��_l�kx"�x����U��d�ELw^�u��6��a:^E9)�sg��i����7n{!�p�,���ǩfr�w�Y�R��O�LR8�� ���MBf5���v#J�7��ՊN��3��ݐ�l�(/��J�v�-�K>Y�H�΍��۵i��&Bs�c��p�-5���,�K�N��q�Y�2�Z�����/on�.2��w��r�q�����@J6rm� 5\Y�����=n{v^��&���ȭg�6k�Z�ár\r��A����zuV�Q�+�xU�|���~�p海NZ2���h[���̲��5-4����qP�Fٷ��3^$��1�v8�XP��d2��뮩��Uo7@�@�-l����gM{{6VHk.zOP�eٹa���1�9��WY$�e;N�eI�Z���a)|f�UW�c�z�1ѓ�G���=TS#o���[<1'=��)xQ�{��ԣO Z�w1ƃ|��Zg�(*
z'�⚍���<�\c��=P���B
:�紟���)���;.����G�|�v�*�
N��B��7N�Ukc^�%s;d"@�|^�����(ܺwᶩ)[G#ntK�;�Z��IVp�],T�]��4GzZ���F�ے큁��> �9���FC-�x�|$sf�2�#k��,�<$9B�/�D��}΢��[v���]�{h��p>Eȧt.5)�ߦEPxdgep9�	+>[���h��#�n�)�%��l�N�{\rz|�b`�i���4�'[\�(�cYSFQ��ilc��[Ě�=���2��Ul%`��R_9�Ȣ"��9nn_<W��:۝��
�3��h�[�f�x�=�˒s�ߨ�To�T-�>����YEA�&8�ދ��iQ�E�b"�m���ވ��n>�.��F�պc���^e��Jn�އ�<gk#u^WZiݕ��BK<%X�C�����a�x��Z�v�U�x�eJ��Pq&R�VI�j#�o�Tl�N��XP��ä�$؋�b�ǚz��%^%�����ݧ�ް�4�r�Y�'=�my8a���(DԡgwZ�%s�J݅�y�2�����.4�
ē�	3Y�Bڽ�)�S��j��96d�WA��O�aX�G�r�sZ���	e��˜�:.)E_���"#��OC:CO�;�QZ�e8�2��s�^H1m���/��>s����X�"竹�z��.h��,��ZjG�e��w$�*��ZC��r�B22G��2������!qY��rs�\ߊ#��m�5��R���	����
*������J��&�ˑ71�b���(j��:+���ޖ�+�p*�5f8Ÿn�(�65��?��� >Y�X�'��W��v�̝���{���	Yfg�B�*�3����4���	� C,\����0�b�Tq�b¶SԎ�.f��Υϯ�qr�&�C)��q��x[�=�/�I!-�WӄL���E��q�k5t!���=�-/e- �>O{�nl��[��TT8T�)X�ɄokT�=yo�fZ-��X-R�w��n4*%RJu��2�r�0v79�2����I��oa�p�Nu��+��`<vǞ�����we2t��5y�Й$衝�W)\w<��eѫT��)E���O3��eq��I0Y��WS���ے1��}�5����L���]kX�l�"���8�W�&sMT鸧!�G�rv�.;l�����g��c:;}٦�В©CX4:�]�zz�Jp�,�|������)�u}p�H�Ⴌ*ޓ݊-���J���Adj�^��M;5n�e�5��/':�+�oJ��<�cz�bE���gY�Gpn;wJJz�$��δ�9��p_��傰�#"G�/��m"��1N��/"HY�N����16�]�>��::$.s����y�Xo���Pwb�/<��h�"߰u�5���WA��N�Zǫ:Ɍ���^�k�9��c믙�4|��7=�,q�=ѻ/��S�qÝ��@5���UB�-�T/�s��xO���H��C�<��+�i�@4�;W�k��p��	l�ƃ~���pE��]���c�j�ወh��m�o�u2~nNB�z���[�eTY��@1P-X��4>Ȯ�3���s1j��8�
��M��7+�D�v\��%|�^�YFf��:�pR��v����a�f����\��c��A:�a�]t,Z[`�*�-�X��S=�n!`�7Кٲ�Yz���
�`	U��5z�L0�;��ռҏ�;����qk;�8L�wXj��K og�i/׋�+���q'#5��g��F>7ѳ�!���+�6o�V�5�vC�����'��hb�w���N*/�pm�O {H����c&�cSň�!.��=Rb�A����"�/����`)n�c�P*k��rI�D�|���s����=�d��<�pN��޸�w9���VX{�KO8ꛐ�$�7�vu/Bx�r���Me[3��|�Z��o��4�j����+���@S�*v���%�kkM��6�.v��h��	_�WB��s�wq�{*��9�W�ʾ���~~���.n�!�e۹Y+ �^Z3k�p8���ip�gF��j��k9��;�)�}��b
`Ҹ!�w�k+x
.���d�2R����4�����t�3j���f���+����o	Z;�6~��j�쵊�<nb�3s���7�b5�@2�|f�e��P�C밖��T��T��%]}�֋jQ��יW��S晏O.d��R-ɩj��M\���<�E��M-�%%fX+���^*�z8�x������Ǝ%�0m<,t��Mj��iV��5\�j���7{���D�Cx'Ŭ��N���Oi��D"�e.���t�,�Mui�ƶ����;�{���[�(��Qm��s���GS�)>�ą��;�m�@�j��k2M���`E`{��*��u�Ҏ��L��v�ŉ�uh��������t�.Gi�ݗ�U��k���/�@N"f���У/O)c"'�Dֹ�B���xo��rx'
�����J���S.�s[�!&ﳏt2U�øAm��yĪ�:���<��D()�*�7���g{�M�s5�?	oP��#e�Y�;C{o.������5��2z�+��Ͽ'�Ã[��E��%	�W'%ea]}V8EQ �W�������٫�<I̝���lƖ������KA�P��n���]��d��\�������빻�rE[\���u�S�v[ٮƩ�ʷt�SƄ�bK9��;�y�ؐN�/D	���ԭf�B�"�t�����Z�	��4�2i`��ϳM��A���!/�*H<S
[�eK��h9�?�
���k���㪌�OI�Z$.�&]�J���b߂[��0T��Վ��S8�c۔��Ⱥ�$�#�v�M�Ū'��o0�]IȎ��sz�kOtj��йQ�}f��փ+�+hfnU��ƅdʳ� ���1��^��/�P\e�&c��
�:��]�/.�}��F��I����n��E ��X�1シ��qWK�6�Ȟ}�h�yZ�e%�v�]vgX��z�"1�&�I��"�ʄ�K�ݵ4�-Zh�{���p����H���!����;�z�P˚�:<�z������h�2+�*��PA�QE��A���FVQE�(�ER$c�(��V""C�EUU�DF1F,E���AT*,V,Ekb���,�U��AQ`��(,V
(�0���Qb�B��EQT`�UEA��P��`��1"���Eb��b,DZʈ�E��$U�DEEX���E�"1�*�e-Fҥ�P��Re�TAPQR�j�DUB�1Kj�Z҈E*���b2(�m�U�j�֊*%eX�mF
����T�J�R(ŕ�km�kR���֋D��-k"��P`��R
DAER�T��²��������`�3]�.z_��l�.�͟���jun�]2�N���d�������I��w��z���	Ơ�M5�5�N���ec�8�h�Z ם	2�Q��6�iI���Vev]k��X��^�ϑ�o>q :�ݬf�K���|4H�fE��-خ����m�b���b:$�9Ka�0��n�%-d�t��O���IX�lZ<K��c��y8������\��b�{l��x�^w�C�|+4��
Ԟ�"�=Rw`��7�o�B{�i�er��It0�$���
�X��:z��o�ccL�_�K53ɶs���+�vU���=\ۓ��4�s��J� Ŷi��SS��On��XiX���6hUq(Gp��d$^�C{0�����:��=z�ċ򼙢G.e_kCQ�.�G}9j*�
�Py�f���-��T�X�s4��#�3]�������H�,�n4��j6�lo�"���D�JV1ӡ���o:�S�ܜh�֜�`��(�V2�����T�����>�Lu��C�)��kp�Ӝ��ٰ.3��z絆���C��#
��
[~߉��IXZ,�]�u��j��@����U����o�*�NoQ8��^���W%D¨����ѱ�^��r��f�f�s	kZ��>=Sʫ�e�A��G3�h�$��>>]�1��%��˛Qݼ��G+�dK��`���w��y����<QaQ*�%=�F��c-ĉ}����t��3������8ӧ��u�zGZ����]ܛ��>��d��>6���4b���36/����;���ew}�e���&k�M�wS�g���� <4����:�k�jnB���#��rߛ&m�h�1>��moo�������G.�{�Im�a�5���3��U��øX�G�,�xMS��<��wsK#K�����	��d�2�=��.3����$��NaJZ�vj�͖���T0[�M���h�
������J޴�o���06�k@��#J٬{��> �P�m��<��e��.��$�כz&���y�W^9�\����$<�N�\�16���s~�U-�J�\�	�,���3�C���n�M鋕��ҍ�Bq��Zd��(���/�oJ�7�/��fIY�aF�[m��J����b�Ɯ��O���4�M�t���iй9��=U=+�Y��[
�j<����8#U��Xz�,6g�V��d����ȇR,;�;t�f��nv6��o���2=�w\4�M5�U��y��\U�L�'e2��sk�9n_pZ��%��w8��h����G��������b3'u�ѰΠ��X�[ҁ�˼Q�is����|X�|��9�D�H,�s��s�����y}�f�� �|1������U��f��<G5Q���ʜ����9���0�l�-wc�q	���+4��ݬ��8��M������2��
�穕�Rz��E��rb�Z�bC�Y+���C����>Z1~!�AP�T���E�uo2��Kt7��:�t"���6�Q��OC�Y�1[���-R�,�q=R"�xCmi�j��o��&��D�4���%#$�� �D�PC�u�6mCι�&Djœ�e0��١��0i�i�VU��i�Yȩs���؟
�<|:z.�5��ը����N�Y��e�L��-��U��Q��I�"D*v@?J�ݜ��=	Y@pK
G/��~n�(�n=Q���ڵ��+pP|tr�>��KX�Գ��%I;1@�9���U�W��#t��!2�-��VTt$mq�Q ��*`�u}8��Xu��s֧����B*��]V�����Mܙ��ݬCS�ޗ�ƪ�R���޺�����kQ�*GL����:X�q⁦�����1q�<O��{b��8��Vz�(��^1yWdKY�C^2��z��EC��%&���{q<gh�κ�UqO��O&�Z|t��r��E,-��Q[HNr�v�y7PqO'�߀�S�P��-��'���_��Ul��Q��ӽ����9P�c��/+,!����;g��&E4n�*W�e�R���ͪ�*�׷��|w!�%�
���L]v���!r�P�E�]���5kmҵ�M�cL2,p�d����}z(������OH��ra�Tiֳ����P//��e��H:�)E�ܥm��\���1bJWb��E�W!�Q"D��q�u6�S2a�,B
\�<���c�3eLt.d|Wɪ&W��gf��{��*�3���o�B��w�)\"dd�6���R�$�`��l��Jc9��p3�l���ƺ�n������4K��&'�R��\�	XCd��)I�e��B$'&��i�BŮ,�xZ���[���}��
�:k��N6rK�"/�����e�vh�R�e�,�̗��pbKAn�p�:ۡ:��KeŖ����޵��Lx�� ��:�
��R�$!�Y^f�c����VBnbx���l(�e{��V���zϹI��vWu�K+Y��g;��}��k���c9:�s���vX�"��v�.�d�q����V] ���J��)sc�up�Ӱ��z�������6��x�-%U�����tt�����^.������;C���Ǐj#�P�r���6�A�ժ����:��Ů��جս�)Ț���@�'�wy�����QVz_�����~�*eA�@�6�Ɣ�g���25��M�x��4��>'�d�sz=�FB,�ƌ�A���u\��J����V����/YH�fD����	s��Ke�$����_ �<�X/��L��fa{�G���0xFKk"Hyɞ_;LNu�;mř܎�y��P;t�M:�{J�L����C-�+x�v���*�)f�[k&S�h<l]��N�h�� ��t�����f���=�;:<���wX�ur�$�C���i��NN�{�i���՚s��Ϯ9
9��=/:K��TXY.�gV�����Y,��(����p�}:v�f㪷/Q7�i��B�WJ���,�Ŗ8�;�/���!���ʕ�c����\����nQ;���Y�ά%7���Akxf��[u�=��T�������ٽ�z@w�Q���M>�ɴ���}�-݀ZTn]�;�F��w=]Q9��eY���1��NL��Z��4��6]>S�^����\W�۷�	����g7�oI��O���s=���Nm�ơ��3C�S��x��0_l&xf�'#T��EY�z�P�ͤ�p�t�g0ە��QR'Vh��,������*�h6:a�i}�XؠUy�4J��Z���(��k��u�5r������̊��8��*�Bu@�lVێ��,��[2NU��p5f{S��y�%kXh�pPTGK#�a4�1���b�|�9[maF����z"�@&��NR==R}�2kH�Y|�W����Ws�E�Ws�o3Xё���@1��A��F�ɚ'�%�;����Y�2��d�+,=�M��hm{=��+*eShJ�nY��]��s[<�Ѣ�jҠ���lVt4�7+�EC�x��_4�����~�,�t>ߔUyU�&'0,�6��kx���W�\���7�o��t t���H��FT~�\-z����a�v�[�/u樭/eqoa�6��؍GP���K���]�t�6��K0+�F���n��oK# 
�kj�erV��R
p�bg�ېe��֮��"��5�T�v8z��i�;/�/��������nJ�A�e�H(-�z��'9J�Fd\J9������%���8p.��~**�AUi)��w�^��ˌ�}]r�,헥��6��y�b߾�1�#�|��(��j��t��*�O.�W��?�j�i[���>����5j�d���%�C\ƃ4��O(��̛�/Imo�rA�L�:�)E_��m�zT�eY���(&���Z6��j� t� ��a_b��R�T�e'�e� ����3�<�āq=\!�ݵ"����r\��E����f�k���*�R�L��H�a�wC(!�1���J#93�p3K��a3�P��옋�߹�+�Q�PwΎ�Af��;�k�6�w�Q�/�i�-��7�}�1Y��N�s6�L#"�����z-��t���O2e��TY��E�2F<3�hU��f��˸�1����F���(+���Q��ѻ���6��+;�Mb�c�/�͎�q���W�(ԺvS�ŕ�[���F$C�7�Y�N�;�ј�h�<�})rhQss��4ᛣ�s�����c�T������'Zv�b��I�Q�T$b�w%��곙�Ҷ�WX�'�uַX�;�_;b�m��?N���;l�t�N�T�r��"A�ޭ��lǆ�9���U[��/9bj�"`q���L����rb�Շ5��_{�L�'6VNU{�9U�'R9؞v���}��⤧MAV�wSSªod����[�-D��pM���,ëer�'TS��-�_�� �9N������Y�P�+�i�4X@��)R��'�ECݍ1��}A5{��9gzȆ:�O��g%�1B+�:�ڑ�ɺD�
����v��єF�8�v<�X�uiWwn,@̭����nE���jޑ\��#oX-ۥQ����T5*2u`�9��,��7
�� ���L�ՒY��j��b�)Ѯ��Rnu�R�ҝ�)��*[V{���f����V`"�X����XvKkVJ�%ӗZ4��+��[t�)�͟c�sR�2P68��U�N�i�.:
�X��qv�cA����:�c��u��;��3*��1`��h�R���x"��KT���KͲ�3U�ݖ�yRP�St7zo��t�ƅ����F�,�m�f��J
�V3f�C�T�{������1?��j�t݀XdȺ�

�D� IY��Q��uYw_a��JU6s��v(YU�1��M�����.d�<��xFw#�ӥҗ�A[rӷ�#Dѵ������EG	���M�7.�f�FS��0#h��\��J�D��2��n��Ix�6���03]��N�]Nʚ+�J���6�˜��2 7)��m�vEn�w�����(�v,���C$��ࡥ3��>��i��|3d�s��}�}߾����sdX��I��QEE�ȥj5�R
��U��*H(�E��b��T(�
����bȱ`��(,"����X(���F
�X)�DR"���VE,Q@b1H�R(��,�0"�����*6�H����Dq,���X�h�PTTX�`��Z�d�X�PP��Z�1R"(�,J�T�Q�F"¥
9J�Ȣ�@�
����F��z��a[�9sD}ԅ8S���J��"1�ӫ���\ۤ�9� 6H�	���^9W���=O8������]�7{w�h��g��5����5���Ҟ�)<��<p˞�e��!�Ǳ��(29*(��]vh�b�{��N⩠�^�,����?(%��F�B�BdnQ�U���y�-z$��TY359@�#��R�L�j�B�����ah	N����f�]j� Ta%<�V���m�-�|/����Z���Y��:�u/L�<=�s��3�NP/ y��FPކ��g�y��r�Q���g�}��P��v�g0l��t��Q��Q��c *Z����`���ñ�#5�Ȟ���m�̸���滉�=�b��WrK��|�-��厫NV�^-��e�MΥ���pU��x���Z��Ӯ[`Y�oa<��U��dZE���ӑL�*��6gp����RN
ZrM�W<�g8��ze�:+T���v,L
��Nu�U6��#�E������==�V�Ȱ����)�zwb˫�} �-��G/yo7�WÜ�c��������"�1��*ZYC����Y�'�k�U�]M<���S��/F�O@&�9�;ϲ^vEdt8]6�ހ�N~��]<[���6f�o���b�#6ݶR |5^�VTf�S��ԉQ�����b��̻�8]�ɼ+�J̕�>��OֶӬ>��R� t�XG'�S�s�&�ޡ�s5���x¨kΪ&l(�nW�H-I��q�enP�״�j����k���U���֒K��^�ُ)p//1t�R[@��ԴdN�|�߰)��_gC��]��\��
1���th�
m��丩Y��L�
5C8�r�ڕe�!�/q��9bK�V�#Ǝ -?�����ϯf�	�&4dK;=�9�����mj�	���6[EQo�7V�M�{[���ᾭ���ѱ�pL[�ܘ6t�͸1;Ȍ	bݛ�Q9��]�TQΉ�|��5����w���I��9�F��l\v�Ro�~�ͳ�敶a��;j�9B�ܷsy�5�d%&�ָ5S�t��WɶYF�S�U[Brza�悜��T�vD�p��1�\cKf�*������ՙ�jB��Q��PT�Y$=��Q����^r���d�'²!,�����'� "������%��	����S��C�PWi*n�W�1��j���`J<�AiV,��ķ�s�bk�ܒ:�f]���ҹelz㣌���҃�!�D\�}��\f�yo�8�H�b���v���A���<:�V�C��d貸�AfJ� ÒI������I;m����7��j����tk�*���%H�P]��me�Y�W{i@�
�8���>�<�6�;��ܓѶ�f���uV-�e�S�6oN`#�ڋp��9�&FdWe։6�1��6(�x{����4b�5��FdB79���.�9�
���>)l��i��j, UjJm���y�\���6��wE�Vݝ�z^o���m��R�J>Z���zzƢ�A�tV�'���p,<X+u.V�1.aܾ�y��#33Q�t�+��G\�h3~$t�k����a����s�.h*	�2(��4B�^V���N	�/MAu����&N����Wܳ�L�:�7���W��"
�/��ۢro���lP�S��r�����R�+
�2�}�gu+�b6�C�������O���{�����W}��,����3d��A��E�2n��K�A?o+��9����nnW�BK�:��'h�f*i��z�@�q/x�ַ����23_�<�i�׎"a�{I���3�<;ա���=����v]�;Q��x�E�����1��إ���6�Nc��L;�U���N����E/�*�E��g���j�<��]� �r��fQAF�����!ѐ*��gp��2z�
#����f^dv�)��-H�֐�Y`�����<�N޼�����'!���r��̘�t,�^��m�I,�z�N�חq���Z�<P�*����bT�]�fdiczy*˹�|���E,K�I�S��|�w)a��ӛvӕ(��JFi�������=\��{���]�Z��n�˟,��
**'xrW�sV����"<[�3��/�j�!�������6��,����ɞ�����Z�V�{��7����쓷��ܒ$P=��g5s�A>��ߍ�#�s���6��qU�@�Z-��ŉꁧ�o[���m�E�h��r[���%��1��v9ܳ�+J{�3���*����i|�t"�^w)����ܛ���%����TO;�[{��e����W9�*��%&�儤	��-,��rg���P��OC˽�p����>��(�=�K��K���2�� yܸq+����(�-��6븊��]VL�U~A�Rm�m��M�W��̦H`��|�/%:���'���3 3;,[P��վ ���t�Xw&����9m\)I�iI7y I�μVn@��R�"=�^�E��|[絕	X�pB�����Yd�Z۾rz��N�q֧�7e_0ho�-:�{��@��&Z����yﮞy_ Xg��]�v�*��a�BXK���d#2w(e֙Mt^�f���( �f�\|V�2�z��W����J{���S�L��Qu�x��P�wǚx��\8v]��U�Sp^���s���m���RS�Qm��㉷Y~��I-���+4���/��U<�.W����BtxjNzY�Yk�{BN���9ò��2o��kF"멧s�s�Ip/aN����b�_!��u˻&kdT_3p�9���rg(T1%�/`��μ�̰&L4r�R�,�W�� =�H�]�m�v�];�s�qJv.�X�����!˽�Z!���%֭=��Q�k�V⟕U���� p�=\���$d�A&;=&*'�$��"���Vi!5�u�#�l>|��$dB=��;rgLe�=�����*��<��>�e+�L�|`d�q�9��W\�L��"��/;"��wZE(+�R|vb��kj]�6���(J�q���4�Ĳ����o��g���
�p��\B��/��sڹ�Dߣa+����\y��x6��I1~�=�L\Oe��;�N�uV�Q7r��uy����]�ÃN�q�"dfEvN�6�1�9`��p��.�w���5B��d(��kw�o?:�y�<��y�T۶��;QaP*�R�Nhœ�z/a.ɟ�)��5�<���ݻ�;7+��?,��6��yh4�����;�{E�ۣ��H�l%#.�0-��	;�I���[��ld�vn�死�q���e��K�4U�H/Ȉ���9�M<���ݝ���q�^=�G�Zo͉����8��]�l�ժ��.s7*���4Y~�"�+XX��O�����ܓa��+5�g�^_Fxɭ���M�Wɑ��ښϓ��ᠨl&s$W����V�V��
9�
o�x�n�5=���ћ Gd����)o(pZy�^.��=�g
�a�/tTR�w�(�]�E��i��>]IND�����y�u������6������R��ʛ-��n�ؽ^�.&'K�|�9=�7����Y��m�[;̗puTY蝳\���M{zܑ~=��ގu�H�]��w����(���ɑ��Χ�4嘭���Fn���p����=Y���/x���;�=���Y�o��rT�;����di�k�����"=��)���q[��[
��P�F��Ca�I�0�-)@�������'$+BdnQ��g��fuU[⛭��]���d}(��<np�țYo��
��9��Z�+K���Wǩc��nvw��� 񲜫ھS�Ft��nʨ�����W2��\�s&I/���3Q���/��_uq�/{Q4���U�$<�|S�\�ͅ�Vi�r'6��#W@>ZOp*�T�~uXK`����ё�X��nfd=�q��Q��/�9��"�Ft��M�ê�����20�~�b�g4�o�����U�H}�����\����T��F��+N�p:�N�����A�tM����Fe�F7u��{NG��!Oe*&�ͮ�ee坳���{b�'S�C\��_�S�1��[��1�}yEĎq]Y� nI��ۏ6�����:��7qb�IryX����Lt�a����]���1u�B�TB]l�Ռ�jT��+�`c�sA��{���W�y�K����q�q��i�`�ZWq�8�� �%��:��ӱ���Z�WQu�)��w���]P�b�W��6�g�:����=�ft��r�\�Mjjw�Q��l̗([3L;��.���i�nH�a��Ws}S��2�}Y#IZ깗l�B���;�{��Sv�΃�C�x��^6r�>���n�R�JW/�S��x֥l��f/S��Gqs>8�9-�Q)�
7�j�Wl�L�"���f��"�ʆ�М�%m5�ڔ�P�ڎޥ��p��V�A{(�,���9�e\d#p��w�����A��+�Ws/^Ro���i���n��,�V�tJ�/�����j�˺|�Y���|�� �T�:�o�ԍ޿�m�
�2�r�#¸�{y����G6��^^㢹���Hv�C��b3y�+�F`[�f�U���9��sooLB�E*g|V��`T�e�ĄdC)�k�M��3��b�lm�{�[7�Z6�3êa��&U��\6�CS���Z� �	��֮�W�p �kFc�˂%:�X��}z��*��q�)�Y�qA`w&�i'�f��,.�!N�Н�.�0w-�	v@�r� Q���I�d��]�����b��l�2�=�;�G��!eZ ��b�����������R%b��ĕ}�9l�(J�Am�om��l��|���XAm�^����F(��v��42`�o	pP��3�mW;U��p�]�\�>��Ţ�T���R���M��-��oY�A;H���4v�����^j��L�D�jE/"�㫽�S;OI4�V�ź�Ļ�%d�5����>�qIcu�H3��e���;�z�9h�G!߫r㤹X�mF�dӿff�_G.=jG��	��9X�O�w�X4p�Ca�
V��ߢbf'�3>�h�mm(��c*J�b*�Y��H�Z£,����26�j(�D(,� ���8�VCX����R��b��QUPDR(��Y
�eA`�(�TR
�QH���
DE�cY���eQ�TR)@m(�("E2�V�\�X1JA��"(�*-��"��T���jiDTb�Ī�Dkb��J,\kWVz��U�����Mbc�
�h�Q8��O �w���s�+F��=NKb��vsR6����^�-8��j��"�)���e��c7��E�r4TFd�=�#d��CȎNqt����@/��z���W��j���ш=�>9(1���r
e�zd�?&��W_�VuT{��Me�M��-�NҪR���Y]	D#H�����ع�̄�&�0��Ou� �yI�w|ݡ��v�EH��岷")�wO5ns�3���p¢���4��ʃR�8�̷�֍����}N97D0��~��ݽy�����z	 w�W�t�G�ߢ��^a �v�,zi8��+�UZ�6}Ï^�0*���탲���<!�;���U�A[��&�f��T7GwNmf��<�]T>G�����Ve���-W�N5����l;¤��'�9�ε�W����6�pjp�I�ۺ�_{��Dz&�=i�������8[����=F*����VT�l�:[Y�\m�r���:�,Ƀ�sL������W:��'"��r��~��ɸ⵬��g�	)�ܳ��CaUOu�WF+��9smsz�{څ"��~�Z5�-q�$�ޓ�.!&����m�ż-��xg�9�7i�H�c*�c�\� L��[�E���>��J�D��IVo%� ��,�[����:�A���%
p�-O+�gf06�?%�5�)�<W��G
z6����<o��'�C�xu�p���"6�r4�qkaT��]�d���hK�Q�-�R��������(5k39�Yyu&"_.�c��y���Υ�!��qe8��ܢ��; ,ѧ�.ڷ[*�#ʲ��ٝj����nVҝ��,�X�qE�{���ލ�Ĵ��#E���R_)��"�{%^���5uP���ku��ʐ�p�ШG�&FO^�h�8�[��\r��41�#l���¥��Fd\J9����
"�Կ%'x/�X�.*���?z��*����zZh{�gI�P؋��z0�n����X�r�I��Ћr�_%N�Qw�Vn�[�~�oH�����Ov��+����Ԭw鵦��K��f�^):��t�mX��8i�CS9N��(��;�ݳ�y�^PM�U�zК�4d�]wxo�%�E͸����/X|4��3�LT]-�y��Z��i�V�Δۮ��.��#lv�����MV\^��	P_D��ݙ�ej�$[c��Mu������K�5j.��7$]RA�_M���}����M�,imE������Do��ą�ߗ�r�<\rRR���AI�8!'"G��7��Dr`�od'c{�A�x�=�^,}���ktw9�y�KTEB�)��Ao@}���;�n�[p��fb�)S�{��<}�
�5f,1A��B�`�T2"Q�OgQѮ�nB/1rO.x�~��I�
�f�i�=aY�x}@Y�C��HC�+$�</�q�4s�+%O�g�о�oO�f�/(�(����*}�{��z��o	�� �j��ɶ�8�VT��3l��:��O�E�)�/�"�=5���A�߆�G�I��������VJ��E�hd����N�/�'P�C�YLX�q5클�u�āԚI������^��}�Oz@�&��LC�l�%0�9̀���Ȳu����r�g���h~<����S�I�N���������������;���
$ěd��N�̛a�:�d7�&�z�	�/�I��"�i���rie����C���W�}C�X?�]�W��ʽ���׿�Y>5��9]�U�؈K��v���h�^��U��WT�=�-j�+������*�[;V����ƪo������b}F&ތywe�FZ��o�� 9�}���.��8�M2VI��7C�������N�g�����5�m$�ɣ��ԟ8�y�y��6Ȥ�I��Bˏz4�>G~����}�z�!Ͻ}B�N�<�I���l��a��q�!�>d�'P�r��Xh�=��z��y��*��i'ɦN�����&}�{�~���HC�{�d4e�!����6���`C��=d�O���N�������`u�N��@�ӕ����}��y�w�z�������c"����/Ԑ�i��
N |���O�XM�|�hu��j}a���2�������9tЫY�6���و�:�h̀�1B|ϙ<d�쀤����m���z���q�o�j �{�b&������@4;@ϾG�F�N>2���Xq8�����}�HCS{�m
�|�@>I�Œz�߬$��6��<�ɶO�:��;�>߼矿{�u�|	����n�|�����l��O���~~<�������&��6�i5lP���'�2M���{��|��߾v��}�ݓ�8���-$�O'�Bq����:�u&��z�i�!^0���''��ӈC����H(m�C��y^��2�������_��>�����2Mj�ĕ���èI��}��0��u��O�
�s��I�8�FRq�ot�d;w�:���sZ���y��c
�t݁�OYn�N2~��'�'�Y:���5?XO�*u=d6��{E��0�ȡ�Cz�$����<��j��ǆ�����Ǵ��߇G��ݍSCD*^��Bx�8*-t��;Z��84��~c���l��yd�M�\���\��M�:�Sy���c�f�m�徤&���R�ߑ�z=�v�e=?��>�����`,����>$��|��}�M�^�5��q=<�z����8�*T�.!�Cl���ӷ�.��?oy���������l1 f�ì��	���&��<2�|�����`^Ru��?j�����Ę͞��4�YY����G������w7��!�J����~d��v��4�@�S�1%B�P��|H(c�x�]$�]��??&��)18�wI���dR
C/�����SY�~���?gy��w�T�!Xw�m�H)��g��'P�va�T��I�R)=�P�OP�SN� bM!_9�d�)
���'��O_�I�PĂ��|��O�9��O������������MP��>$<����1���i�u�i� ��l6�$�V0��eb��5'�W��Y4���3Q��2aeDE�zR���M����{"���
��:[�~IX5��2�
�=f���Xxn�$��̪AC��j}dӤ��_�q�O�3:ʛd�:��p��r�_�y����ןw��o����a�߲u<CVM���2c*m?$��X~CI�7��Hq%I���:�X���*m�8��=B�fXm��S��>�9>�� vb�7N��w�1�ԟ?&���N ]�y۷�)�F���(q4�0>o�0�$���3I>fv�I8�@�T�aP�+���H)x�Y=eC���|��y����k���|�B�� bOYܫ>d��+���I�q'�ڡԕ ���$�.a8�q �ܠbC��<2�Β
�s2VT��0����J�f����s��}�w��I�'X�N����I���4βVN��n�Xi>��i�+�T�{CHu%`ww0*AN[��OQIRq��v�H(|�ۯ�o�o�gޞk���D3w�НS���ɍէ�]�:�%�ΑY��~�5�����Mہ��P��8��6�1�����h��o5XY�O+n���+'Q¾�35u&��U�q=#OpK�#���ŝ�7��?��N�IǬ���l�q�_S��<H(
8k��k?Xu4�RT�z�d��6�Cz���T���Ɉq%g^�Ï��J��=����|�6{��}��΂��*~d��T�B����|��P���	�l�}t��e��]����T��@��ۡ����FX~���b�^:H)*Sy'���=�x��]ѳ�w��o�y�L1&!Rkt1�aP�;��Z��V��T=�&=t��8���g̗���JΤ��Tި�S�>E:� �Xzn�$�<q �<�N��u��=׺߼�Mt��?&3���� ��;�i�%e@��`�c1%B���1��Vk34��6Ԟ_p+:�Y6�ytì*g�}a�1��*u7�M!ĕ��w���������w�v����q���O����B���Xi ��4_�o�� �́\I���ϵd��&�a~�!����Y������_��Ĩu%g��w�6~���w��~�c>d�*i4��CĝB�4v�4�P�J���8�P��&2VT��*M���4�d�
y9�*M8ɷ�¤�7�4�Sh���:�����s�w{��&�1H,�Փ���:�$�l�R
J���d�*Au���0�'�u%a�
�r���,3�%eO��iǈ���3.����W����������J�z�u�����S��AM���I�<q��Ă��8�08Ԃ�Xm1����4Ìĕ9�4�Y8��tǉ+�?w�~���u��7�_�M!���Rt��z�c
��ȸ�hV�T��1$�lՇ����VOYU��O�*O���@�AC�FXn���1�Ƨ����������|�}�1��t��f9�H):o�4�8�<7���IP�J��O��'�T�3T�I�+'���i����`z�u����1��T�<7a��I���>��]�]���ܥyؑ`=�e٘s��SZ�!5/)�'�Y�	q��:�멘���5+_e���j�pኵz�0F$�H�Y#I�$*����.���v�έ�#A)�[x{$�;g��W�G�=�Ea�e���&�H"$��=|t��LH/�i���SԜ�=�یR�,�=M���R~t�Rkz��'XM\O����W�a��s��7�=9�3�������I��Ag������8��x����6���K�
�C�+:��t��� ����c�AO��%I�4�
¤=C���mH/u�-����y�}�<�Ld����S�f$��XH,�N���J��_�6�3����i�XT�vf�q
��7�N�T8�����o�>���j�Eϼg�31�i�>����G�g�v)�I�/u�i �S/}�Z�ô1�Ƥ����<H)�M��C��i ���b(z��y�ͺ@�T:����'YY=eO;�?$�'�w�y����^{�7ۿ:J��P���c�g���M����R�V��4�d���C�+�N��s�!��h��� ���v���y�bC�C��ۜ��ܟ�޵��{}�� ���1��T��&ٌ1'�Z�X|§r�L`m�}i�ɿّC�+רRq
Ͳ_��!Ė}��ueuG�f" �ޜ\�?����O$����c��l��P�5��Oj����*VJ���������(bAd�y�L\IX�Ğ�Y�J��2��
����g��_k}������i>B��;��&�*I�5�:��g�VLd��P�*q��~���H.���3Vk>9d�ړY�x�
q���g�:���L�jt���U%�p�����&b*\�.C�vt�Ԩu���d�+'��>�J�$ĜB��P1�d�q�v`m���I�l�����P+>�CI�M��ya�u%x����}�����w��wN�
Azk�'�� ��Y5�Lq�M�bC����y=�08Ԃ�*�l�y�&%gbN;f$C��!���Ƨ��4�H,6WѢ�����.�P�V�к��pOA�mi<N����0���n�{0]jqX�tA����2�՝aK�Ʋ�#�z�5쳹03�&�� 蝢>{r�����}(@��aXأ3�U$�3|������o�V|�$���+1'�V|�o�C�J���0��R
O�P�����H�i��
��:��Ă�����Ƥ�h(J�S>�H)Xm��_l��w������~�m�;<̝eb���st�$�+6��'X|§���@x��V�'P*C��4�������O̪��ɉ�
��P�R�<����zw��>����t�m'�`V�`x�8�<f�
in;0��1���b�������� m*�&2q��<��x�m���4�S^Si4���q;��ﺾ~�y�w��vH,�=�O�*�p�!��&�g��&!�J�N>��P={��$��i �����R|�?�Hyhz������Ƥ�+&�S����y���{{�{�tM3�1�}�!���i��4��V��u��R3��Hq%x�a���Y��5�B��J�}é>sT��?o$�c�n�T*x�Rz��5��uο������ ��g�u<`q�q%@�VO2�H)����ĚH���w~4��F~���-���(�}���w�d����P]8]a�r��t�yB�(O��\�VKr,�(6_�������UEH#�A���:5��v`�^��:��,�#/%ԙ����-��1�(=�H������TuUq�-��RX���c�k�������n�^;<���*��>���d���[	u,�QRR����Ȟ���if��rd�{�cso&�e�o]����"e�M\��G�-H�ׯ0Y�5�Rد�-�igf
\��܍�{�w�miNl���[�U��f��;�B_�����w���%O}�eLp�"3��tf�+�g�.��!鐊�z��w{瓼{y�����>Y�p�Z�<�t�P���ĺ��r�L{��O��#�Y�DR�dck-��%���5�,ع�ɕ�H�6G�ܭ)ɻ�p��ˌ?�[�=Z%���>N��U��T��=�c�&3-�RZI,1�0#�̸�u4�x@�/֙��<1��o�t*���g�/z)���ܻb^� �0 |?1b�r���2�y���������¨y��u�\ vUw:=ˍ���ER��^��F:�y�J��Լ7��S��ic��(oo2w�����+�yԼ��t�YJx�cuW
�*���u����vEb�,}�<9T �tjʺp ˗�ӷQ���W����*�[��_�0�4:<��b�QݣtT�f�_mi�v���H�M���EZ������7Η]��b{�8��G��V.�f���L�4`�Y�& �f��2���}^�����-���_u��RY��xN���B����b��3�Ek���[h���rV��2(�y��P�eW9-.Ǌ%�n����<�R�%+�(�\Oݾƶ��Wڰ76�,Ţø�2 ,^Ћi�d�aM6�cٲ��ʻ�w1� ��s�Qp%J
�� �JP�t�g[��t��5b����h����܁e�J�\��!��f��wƛ�]�/��o���.��3g��:�9����G;5T�T;2�z�S�@v����UݙhT�ƫt�S�L�1����H3+=#eL�#0��,>�J����x���ç�t"�]@I�N���<��2�Z�3���)ؒyB��Ue�J��N�� ���qΝЫ�3o�H<V�l���QfC�w8E M���M��V�l�~*��M�:� �Y.�ʳ�>B����1����c�(v��!Oa��2���f�&N��8<	�%&��,�@l�e���X��l��/2)I_Py����Ԋ8�s�o���f3kfH7�-t������o%\���ݵ|��r���Wo�P��L�3(�[,��B`��!��+vԩ:�h���<:(���2�S\�iu�\�׋#��m��b��B�L�Wvn^<zF3�Z��pwc��U�����QMd#��f�/�������[}��Ȭ(�Y�.�1��2�����ԞX�ƹN�/	�\#3-.�Swww����M��j";�i�cgt���`��<�Vj�n�n����1[h,t���:[�7�S�j��W5��V�q�/�)�1�6���\;���RgTu���W)\�xoJ<�ML�t6B\�F���YE��[9��1w.����v�>�PY37UF�W��o:����H�lHN��e�>йV�P�B�_��oL�՚^���T�S�:W�16V���KǓ�WU��˴��o�4ú��/�t�j[��_j�ݴ88���N�΁{��~Ϸ����ߦ:��%H(�+E#" ��
�E��V$P1��AH-IP)���[�	X(J5�
ł�`� �0Led�Z�EF,�Q`�)P
�FE$R6�d�3,U��(ԕ$DD
5m�E�Kl*)�&GADAF�VDAJ"�E1!Xc%b�FEP+*%f!����\�*E%�T��)�
�V��2b
�hQr�E ���(�(�Jy�{٬gV�Lwmܺ���GKtdj�mD��|RI��巹6�UZ�G8���{��	�%9���u��9��(��x?���W��7����G��b{�#�=DT3<8zUtN������Z|�j< OWתv/1��#t��XV��W*3
D��o��{��@+j	�YX&]��O����ZKyt�4�m���It�4y�/B�_>�T(NK����|Vw~�dE�왋�o�F��"*����)Гf.�F]�գ8kf�A���ֈj�S�=2e�r��3 �d)y���6���\�
�ye^��s�$��4�"G�����Zϯ�{K�����8]7DWH�]EJ�v.,�ā���HxN���|���I*q}wힻ��S���ګ��BnY</Y#��V}f��^o;��ꈩu�����pK��8J2�����5��#-]#[c�c��%�j�� ���ax�]�K��<�%��%;*�u2��V˶c��;1$nT�5�UDF�����0��0.=� ɍFu�[h܊�ѷ�(}c]gR�Y�bE,��8�H~z=�z<rC��z�8�ߊ�񱢅�
�ˇ��h�}��y����ַ���B8��Ph;�e�^���f���²��4�co�)ˆ�u4�_MK�����jzr(Z��0��΋~U�� *�j�Y�cɿ&����G�(o���,��w._PV�Uy�2���<cB�QY�9��6�-)I��P�J{{�P�9���j�
����)غ����0]e�CT�E^r��}1�����LR���K�抬�.EҪ��]�Q�w������TxL;vgauiTu�^d>��2g�f�8(� �岽!�eɪ�ޛݭ�P�
o֮.(���T䮸F���f8Vrؿ0^�t������
 	B�i�􉙪�j�%���c8l+�*2�aim��<��c:�Δ+EC��R�*�bM@�сi�*5��ap�t���M�kJ̼�x.���#��wP���-1<�S��[�fQo!tm;/o�%���G�T$�8�ñY�	u�"2H)�N8�,�d+��e;��N^S*^�"{z���r��'���=�9̨I�U��{ʭE��5���@4�Y�G��TDG��us<S{=�lpW�+Fq��\h�O�p���X��uu�ބ��D���
˫������ׅ�A�J����@' .��j����@scnsevuM�On{,�l<<Mm�α��4=wW��/U�zg{��Cz����|o�W��/���<	+Y���@/�xU��ztꊅ�Mz����	A�����^;C"�[:���Ϻv���>�Ԋ�p��ժ��aU�T�����p��#n.E�)TD��H�r�:�:�[�k�n�����iv.Ԫ絭5
c�3*�eJe��T�ph*�W�NuDnҔ��	Y�jzr'����7@�]��zڛ���Bx����>8mZU�Q��
q�2��s��=m����;r���wWlz�e̅�ˬ�cFyީ��S2=P؋�4�w�R�����Ck�$�ۥwl���k
��0�8$�PE��AE�M6���}���{6d��B��`_�`Zj
����Yw
Yw������>�ع/�X9�=�u�=�wÌ�Ys��`U~�蝈��l��D�����k��I�sU�;{M��O>0jB�*Tb 
��mK{XK���3Ik9FM��=�,����g���W�]ˉ��
ױ��*f���{��r�_�d��G%�蠤Fu�N�Ҩ��7�*D�CM1l��_2�.wP64��^�ȫ2�[�9e��PQp��<�'#w���B���5�U�g��gN'����Lex���@g��k���������Ƭ ��xh��p�`�>.Ф}~��Ԥ�@�f��vOK��g�V@��7�����g���>�D~�{���Z�Y��q\ɗ2�|���/�$�$|���.^;��u�b�e�tI}93�I����kDRn^����Ƴ.���w��
��4R۫�85�mF�<�]�(�o`F��n4�ȶF��]�Oe��ͧL�jj�b����h!/�=舕�E�r�|Ī������@wr�}ώ*��tiI�י"��W�N�~I}g�D��Fwj�>����]8.��RqZ�h�g7
�瓵8���%��~�iA.�:��T��jJ�B�"G
A�3�2I�p�<���=���ƨa�|l{h���Ԫ�u�'��]��f�ޭO��#l�"�T~���ML{��Jqt���s�/O^��h��te�y낆+�=��E@�x�.���t� 8wF�^Z�^_A�-�t���(��(2R��>z���ߗ���ӎ�+�{ ��^fFӕ"�keH��發��F|-^%�-�H��];��Ě�S$R޸���v1ۜNěۅ1ͬy{%X��PU���d:�諶���d���P��y뭰谄X�W�����wy�Z��:��4��v֜��F��_K��J�����nP�[]�+@b�GuQX����!��[������:�����8����{JFi�)����� 8�V��3��`I@�{�^,�=�&o*�L�M� _��}b�?Y�09/��۳K�:�B�Q�t�	 �r���뤫-�Y+ uq /�Ш� c�tׁ��K�쭤����g�~�l[ }�ts5��VT�e}g���,�EP�����7Ӝ��p�񰕨0�ҏ�D���:�����m�b����B��X5��W��)}o���8�\(
V����{�C|Y��d{��;�b�V귅
�,p����#�����.�-�P�V_�n��qп����êÂ���g�U�oՍ���N�l�]�}㐺�GOګI�i�/Sp4P�8<����}��Әl��-�_��5{
�[c����j�
����n��$�p�rzz-��˅Nn6�LduG^ٔ�Y�+j�<7�Y ӝ��3�k�6�e53���`�z��7��5t6	��wQrj��bޫn���=5���֍�w��)9G����j_bΤ��[@ɴ"=��N�_th�)L��6��""a^Y��U�঵ ���.�*��xA���^�.���T9R*&��Q�Y���SjV����xV����~>�WC/���Y����fUـ���"���;.7�����L! �/�<xOz�C[�ev���z<�z�c`�Up� ����s� 54`Z~��{�xA�ۧz*���į{��{�m{�L���U,�� �2F�g"xjYr���ޝ�T��.u�[��V�'=t&.�J�s�:�ŀ��]����n�����������i
n��=f�Z������ڕ@�����U`�0�	\�7/ʌ�~رyu�V�M+6�c�H�8�5��n�������||��	����������=|V==��M^�H}j�*��A�\2�D�����8|;Z�ņ*��.�9�Y��7K�q�L�	N�������KTV>�A�Ȭ�
���9��Ǻ�d��F�F@8bN�@Z���$ط"ؑ)�]M��pRNՔ`��`�f�_{ވ��QMc�r~���ȇZjg�w����Λ�,�@�.�3�S�Y\HN�)p�Q�-L���S�5��8+!ȳ+��n!]u�`�ԁ-�F{�Z<���s������.���_)���{�A�šG�}�W,���6>4^���Wu5T�����Z}VPI�wz�=���2&д�����靅ե\��u�[͊�|���;�Ư���wx��=(ї�s:��DC.�]Y��
���0;]���O>E���[6�w���GNI�^)ؐ�5!T�@#���ɷN�OxR��:S��/�n5P.�S����\x�!0*4k^'�Ov��2�=�.� �\�;Ջ���i��/U�P5�k�5L�æ�=�!Ȉ��,=�|���`�j��Ɔ�\4wѻ��c����\t��T��P�o�.�|�EqQ�ΧȬ�/3��$	���{��eO6�8�E�#�>���6Ӓ-kڏ(u-��d�/P�Lf��cu"�}�}�����|��̪re^��bhp�:M`u���c�Ŕ�W��S/d�S�3��.�`:���| g-�ZtIT׎����M���d�oU�z�qוpT�T60�ȊC�:��y���u��\�ss�Ox�0��ľ��7�}�O�3�?4lA�m�g>Λ�qp���,���A}��c\)��Ɔ�#��X�)~�_���r̝��w/|n�f���;�n����f�_�ܡEU̖!���^g��8v���5z�:�X�1W�8�:�B��`h�]`W�PiT�{����p�ŏ^,v8��v�:����T���������%8�����PL2%��[�'�Zfh�èvV|�%�==BL��MbJ�%��;�vN�NO��E^����R���zࡊ�J��B�d[�'��^׊�"5m�"�:*��j�fL/��́;�߻k�˦0R�e�����-�W�{�p�d�η/���S\NJԄ�t;{�\Y��`���8@��=�f[���s�~W�PP�Ҧg���P��:F�I��o��넞��V��%]&���(f��q�B�bP���Ja�ّ���Nx��H��効��m�Wz8�GD�9�"&��R��l��٪��PJ~^��E��*^�C�}���"���﹑��� �=��pڗ������t����&|�P�V�<HN ��S���J����۲\��]����se_�ֺ�\��4w���JN`8k� UU-���j�&��8>���닂�PU��L+k"���G�*#�y_�k~if�wW^�iâ�_,	b�P�ԣ�B/$#���]�q9�L���2ݑO<^W�ܿ�Z��\(e�)[��À�@U�a������o{�2P]�tߠDJ9���y�ͪ�ڍU��*#�̭��γ�-z���mo�R��n��;1X���"oC��̾��S���@�V&�)\t�b�����U*dZ��g��v�b�G`N�eU�j�mva���\d\����CE� ɶ�Z.�����δ�$�+�����nl����J�{��d�ĉ^î��[�5tك%J0X5�"�!���n�V�|��q�� 0p�����B4�Z!:� ����u���P]B��2�c����\}ܹ��5����3׫@EY�@��!X`��v��O�%�k{�s�WVό@Em�g`z�̪�|m얺�o��TA�|�ڽF�Ʊ�Uو�,F^�ȅGF��lȘ�;u�uo([� �L������i���*YR�h�xGr�Z�� ����+�sr9L�ք&CL]@x�d�+����m^_7i�r,գ��KUn�j��Zb�oR��Wj��An֪��[�:nJHc#0Y3~��L��c�vTu֠�f�+����5�rw�'�si�V���&^��]5V�'op�r���l��a�Λ��	wf��+ffI'V(���E52jt�}9���ͣ�;����z�l�V���
��׳h��w���gg�*�3�E�����H����@fa�}�n�����r)+Ҫڌ��IOgK�7T���f�����*���ɸ{�f>��'ֵ��<�Y+F���D���a�])}(��3t�C0K�fM�(cOp�a<��r:]����$y�e�ҋ
�ԝ� @PB.V�҂5u��:pWn�rV��+:���#�y��H �.��2�}$o4�@Uތ����.�*OzR��Coi��A�IpG��x�.趡O��)��l�,��a��ȔqF�j��hc��Y|���-���oT�g]3�[���AШD&�U�d>���؝-�km�c�r�umW"	���d��yՁJ�
�cw�)ԙ�d�]i��i��7>�����}��9��*A�}v�{�D�]4�����=��;	�AHؤs�݋�[�簝Ѳ������d�N'��U^�>��d�H��
˔���J+�dIm
°RTT1��Vc$���b�`
B�Aa"�.R1��b�R3,�b-`J�`Q)"� �1"ŭa1� �Ak �Q@��J�VLa*b�f"�
�I%k+	Y
˗b(,P��R�əq���TR70PR����)dP�J����FLj���jLb$Q`�*J�PE��
�s0"�WLI\d�j��_sC���>ϰ�԰��˻
F�����|�\��[��j̔%���Y��d3{a���֪��n��Z����n:mӚ��K*r���~g�_ͅL�W�;��f��'$^�)�� xA8�C�E[�U����FՌ��$�;�[��xvxv�y;�S����ε>�	X�*����P�x�x�k�]	\�K����8�<,A�1]ixK�*��r�_�+��pm+'	ۚ�9�瑒{��"��7A��V�5��p��93Ɯ�:�"���ق���l�m��y���V�L�bqӒ��1�d�F�ۖ�;sհO;���,�,%
a ��7jAN'5��(��j�i��3��kx׆�+9R�K��\L�jF�
�W���<���V��x�q�<�Ԧ#�G'�_��IuƵ_> h�a�^:��x͖s�T�T�nT�H�:&��j��\t���\��9�X
$��P�Fmf�������tN4Cf{e��k2�l}N�.����2��d58���HL?w�x��f��G�	��-{���ȶ�0��pU�m�����P��G���Ʒ9Oʯ��'��{]��8�j�Q���U\^��Khe�x�N�C4�Bl�� C:���<;(E�e��kW�i��@�
��a�v�/m"J���3Gۙn����D�|�=�*�^�4}L՜8����=�9;c¸^�|MA¸o@��]����^tՆ�����˛ݲx�+�΅����@t+���^wr0��^�.�*�u~��u�<��mq�Z��Ǽj�@G��64EQ�]h]�}w�%��W0yqR]���`˗,�����NK���s}�0,��?���ӌ+���d@1`��U��R6��s���.du-)��;��������"#L_���+EA�2��ۿ)e�.J�%��@e���H�z}X~������떾Gs� ���A��Ψ�֎w\��xM�Cp)�qP�Q�a\`�`�5έF� �������Ry}��#���� ��C^[k5\�ۀct�4-�7s�ԛ���;�xw2��Ru�£�"���j�'F�~���o9�g��L����kC<��(T�(�b @���#3�������)�������W
����U����d��e�y�;�l�1�g�e�P�s&���R�G
S�η)њU�;~3(΍m�rM�<8�C�]?�#\�{���`�V���cd񠏀�"w�^�;�R�X��p}��\;�<_͝8�p�&�_ez���SZF~��f.D�mW�;����1T�����|/�D�k�S�?a�S�1�"*�f��]���t�pw<��������"�T��W+�΃J�~<�����wq�� ��|m/���B��|�g��DI�m�5� z����pCG����\4#�y|>�+�4�\�$�4�7kzϏ7i,��S6�V��~�\<�/�_yxV�@/�UKK�"�z,���6�����]��OeÐ�6i���{ǡ��n�@'t�����	�7Xj;A,7�3%����B�TX�rtLqSO�&��jD%����%W�Jxf�����D4s-����2�k5e�룮�k�B��r��+��r�����d��Q�^V��o�FVv�:�3�Q���,�W��'/��w`��<QT�����o�8<���L���B�3E�C���zczg�-�n��{v$χ{lz�ˍ�-�]j�*����z�2E�GD��37��ʎ��F�I��o��rO!�V��g8��X�7�GT�{�G�����]f߭xW<�4<�s�HRbT��Ũ<:}���挜���VO������TU���W���4D��L��9�/*�E���Pl�@�B�ڊ�Y
X*P`,���3I���:�n���e:�ԥN��Fc�M��4+X�7��~��䠅o\ӂ�~��uQFi��O���ā�� ��,o"�K::~��)�������O2����������+/��&Oo�KMP���e$S��f��f�i��wH	.v��|��z�[{�jpK
���=��)��!��Z_=�y��@tv��W����[�h��T�}��p�,��P�J���-PsJ�|60)���tβ�2������}��.�f�4WW�'�>J9G�(@�^HCk��{�mɮɌ3Tv߮�6z��z��׷���U�)}o���>Z�O��t�L��E0·E��<;��E?*֭��F�(φ���Wh�OXپ������.��+=�r����Y�X,Sl�$�ޜ�3��*�G�����=���j�&z��Ic��GܓY�C��l�|7��� �Z�Ht��Uy\3�������6dW.���\ԛ���ʻ$K5�]u��.A��P�����gJ-A���u�2���w���xf��w]�^�
著�<�í����zȯUi�Ф K�#��u�\%��v��u�T倧Vm]#�iU�j���[�c���C8p��-m�[�e?r��,:�lnP�,��wtk�Ce�1m�g���)�=�۱��d*���� ��6v&�1�,��G��� �M��r�Ҙ���/��tk�� ����Eys��ۛ'�s�,Uxwp��}Yʗ�P�R(L@��T�W�b�̷k���������_gM_�k�Y;\j.�m���p�'�6�̑Ԯ��Dy�
�0�=���x!�#Tt��#�^�B>1v緼T<�`Y�8��4,���+�G�r�%�<wUi}�ױ/UXk�b�m#T赕_H y�ύ��;]���Wi�u�g��F�w.s�n!�oDe������ʤxM� ���D4ݭF�b���˘�J���%t�5��n�xw�>><:���#��p�v��1�EET��LF
��*�t��66������fQ�
�����ƫL -k��c��~�w�ִErD��g�R�#䠕u���'+
Ճ��9�1L���,�<u�<��N�����
2ӭ�n�)ihֹd�n��J�G������[�sS7b��u��f�n\�W��ȱ���f��(}��0�)��s�_a����c�߹�=�e�W.N���W4��Ss��� �_B��ʌ,�-�>���f�j"���p�{�qH����ӱ��`��Ǿ��"_ثC`��PXc����ϕ��9a2�-�{�Y�i��Vdk��վu��ȃNbࡊ�t%H*:�5����[.��hs���)�fƿ{��vx{x1�<�_�*A�&�����r;Ti����\V_��)N��nQ��U�K�n�j��=Nf׵4���ز�z��o ,� �G���gD���뼠<~>���*T��ș��^�x�T�f�'��L%�V�W����.�*�!<r<i3�S�^�z�:���xxA�KD�`�}��l�=gj�2]ҧo#�n�ʾ� �R����{�^U���
�+E�nx�%����y/���c>Eg]Id��^[Bc^,��WlK%	P��]X��=�w���@��+n�U;j�njw5�C�t��8���	���zk���]w�K�G�h`��v�e}��E�!�?p��F���"�T3�8��i��%�<��緹ĸ�ׇY�AUk�V~����H����BD�I�u��4�^y9ܬ��(1u}usK��B�vf�-O���72�D�9���^������!D�.词/���4�f0�<S ���ˈ�jz��2�NB�q��Pu'2;֕��C@շLU�z|�{6�����:O8�HɗJc�������-Fv$'|������,Uc͵�'��G�uu^q�Ĺ��U皘��%_"7��T�%��+&�����&�yL3P�*�_W���W���)R�_�41]	�Qrs5칫�������O�b��33���^wۣ0eȍV�_:�\'��NvR7oY�:[���3YZ�F/���u��\��g���,�b �s`9�<�͒��N�������gZʹA/{��k���6�j ��3�w�׺{��Sy����Z!I�w5Shg��	cޮ��΃�$t�V�c�@=�
[��{ѯ��Ӓn~��x>�5N��P���*���<{O���J���BN��d}�}g�q�
ϩ���uC� ��Vr�O{�I�i�M���yƽA��r��/ӔM;w�+, ��h�
�qy�I�O��AޞKhQ�)�r��]{C�|l�EHU��|��N��$4#6��w�\�-��qhh�W��l������)��Z���U�l`T������!	<N�g-����¼�l<|� J<)x�.dT��'}�RZyM�J�0���>͡��/[��~9���g��ph>���L���}w����P�}��;�{�Ò����Z�-aʤiq~.�� \�����QW�^�����x���^���upt�1XIQeb꿻^�����{dM�n㮌�Ш2g ֊h\.��=�
�����w����
��|t��n�ܱwns��Qm	D�)�r%YG#�1\������V�j+lr��\��e7g�,ݾ�w���A݈H2_Q<�	��v�6Y�ń�`Һ�E�P�h�q<���� w�RtR���[��#�����Ҙ螔��&n3a\1^�� � ˏ�����j>*���Q/O��
��X>�g�q��=ƸzB�R �w���}�U�<2���a�W���
�gav�s�*���^1���7]�����;�&����ÆE����^T
˾�
���)���_�{t���8gGX+��z�+�]!��� K�`�� ��3O�L�����M�P�U���ס�ŉ���������b�j4`����ܢ	.�C��)�Dٗ,S�|��e�:�N�VyTՊsM��o��"������v>4h��#��
���:��Ss�QT����dؼ�ғk&{8�x��^F��U�½g�qK�8*�r��kbU�;=��U8��+����xv��TwD|MJ�`�コ�R��?y�zH�`ߩ���j�������̵y|��X%�S�D�:�M�5�R���=����4�´���Wi]�z�֦���\��*�{Y��GR�$���ܴ�.��aUk�1�tT_I+�,=��v:��	����4�;	���Q��D�%L樓B����3u�k����^u+}��u1ɆHx���S�]�5C�ح����5P�y���y�Q��;z�(qf�I�f.��ɔl�5�V�wm�ɆVܫ�DY:��-����2�a�������et���C/���X�-R��c^�%��
쬳���>aˡLG��uA2�e�c���ȓ8vZ�H���ܺv7��I���t��O$^�E������p큡�\8��]����[3䨁-%���S8$�����X�:�e���;`�#ݛ�  7al��]lT/WD�j�^���\e�;��+�8�q��Iam̂��9�K�`���"u+�O`@���m�{s2l&d��.h]�&5,���Js;��1��r��� ��2+�_-��:����gd?=��>��v�U:A�{Ϻ�\��)Y	�fh �WԨJ�A�:�-�]��K�l60Q
�n�a���m���ް�ZTq��ۧ\�Z��-��{ۈ�7�T�y@��#/�q�9AP���*��2��Vr��m�KE ���F�$�G�Օ�;-�Ou����)�+�Z)�;	��7���)Zu̗�*I��sy::8��>�z���d�6���B#;�U��ҡ��d�srY҂ƚ=�=��8:�V�dCY��+wf�a�e���շ5ڻM>�|��Tn[��Ԑ�u�J4�7&�m�����I-�w}>{/r*֧|31�{�*��N���]��]�u�i�6H򼬰��=	��.�aA��{ye�t�t�6��aθw1r�us}�b#i\�4�\3�3�I���+�E�E���j8���L��qݧ6?�u-�������W	�p-w�I�������Z{��/�r�H�����g\�A�1g+�,��:��F�7��<LdP*ۊ�VcY�d��傅d̪`ɈTE�*L#�
�HV,�	SV.e�1����B�%�R��Ab2��Ć0�
��
�¤��a�#0Jȡ\`b,,��e�*@̱Lb�-�e���ʔ�0S2Ɏ0Ć\��X��+P��Eb��c& �e�m*&R�bbV��V�ff��B�����[K�q����E�e�%2�eb�1Lj-�#1*c�a*��m��-f%q
���S����
`mX�k&�M3�γ���r�vn�)�7�s�,s��ȯ?y���9��I:8�5�~�ꦉ�\�R������Z������v�6���4������øv=r��Ӗ@�J^�̰]z�y誃4ЅrT�O
��D V�t���k̹���rw��'�Z1��������>�Ԋ��Y�~5W��XW��yv����=��1;Q7Y��QSVJC��A���/���A��}ru?^�ȶxì����ת�1�F���7�᭞�	��3ø���a��=��/R�0?�n�N��X�P�_-^5���2�-'Q=֫��6�ێ�d�uL�c;�ȘkB�U���C��sL��tcmfqM�;��{� �{�{FB�.pӘ(Z��QS=]&-ߓ�޷�ω)Q��$Ji瑤k=���F�ٴ^)��A��I�Z�]���骼q ��ߡɖ���ynV`�o�@u�Nn̠<_�O_�VY�EL� JF�e�]��{�����T%:賩�u�n�x�Zn����0웣��v���]w�%�6�fqW[���p�A�WfCFw=72M��d�oF�bcY�C�/`ët֤�/��[a�i��j��z��T nd
�-���^��}��g�ʇ�e��t�7R�S5���Vf:�z��蟞?���UxP5�ө;�b�2K�t`�l�������Y ]V�5�P-��gp����k�Y~>zݼw�y��C�:�C�B�8��*[���«*�q��o�ɱv$ٺ9�t��AR��_{������~��Ҧ�Ċ�Z
s>K���\�U��_������7I|j��8^�
�%򡐑�|'_Vg�t�nϑ���Tի��47
��?UD�x��\Gec'�{�e(�uU�4�&	vUS�CBeژP́���G��i臕������C�cY��Y�5[t�_�}�	ڝ�Ǘe��3��;`xA]�V mߗ;C��[5�ӑ�~��4�E\����)t=��kAf��[7��p��K8��R��Y�i��l�@f<��fnͼz��̝��-�������GN4�"�y�QV���NF"B��j�t=�6��jI�+�9�ys�����<W�b`��fܞ���ԭ����롶�TI�f���)���+�Q����u�k)d_��W]:N�ؘ���$�l��W`��S3q/�>Z�j|������i�����k�<��F��uQ��H�K�H72���df߇�=nF�3�
9�57�������*��ρ��J��}Ǵ���T5U���kj{ӂ�=��F}���u%��c� ��Vr���ym��R�;vmF�I����_��A�����k��AFݻU�.�uTD)�;��O���0���2��E״;��l�F]T���Uq onqk-D.z�t�6���4T+˫���(�KW-Pq5���afJ۝�����������|�;:.��x*�`��᠈%���N��
[o\�k˞��l��<�k�՟��\B�攝�v���ݽ�ե���}J"��,=�̱�=���S���`��M�w��P��Vc���{j��o�.�RQ����-R�V(N�V�2�Q�NQ�-��K�;������>�Y�G<]P��G���}��M����wNM1�x��Gƪ>���h�6�\��`�m>��
����`Ox���*#�*�_�z����dS� 4lۓ9Bԇ����j Y%L3^�:0{Ɠ����h�ҡ�t��j7͡\ �i���N��ǀ�=�c�p�jA�\)|0wr���/GWG��_f�K�$�.?]�!��"s�wbc�۔�*�,����s�͌���s+C�캧U�[g���&�qAX��1���wL���쩉%�A�w�a�<��p��"�O�R�,�]$�%���^cr������i�0��/���P 	`�(}P}��zJ�k��>�R'enx���بS�j�ɩ�M�����.U��e��t{�F���b{��Z:韊E�V�8�����W����B�Ш'f�Ȳd�*���`�o�F��o��X��NN5��h�ץ��n��U%er�[ZJ絖Էa��t�]�0t����c��/ԅP�V��x�\B_�D���|+g�.���˃��lS}����I�2���C�"�:��DDpxVP���<�xy���F���)_�p���{��t��~�,��|qW5���f��W
��^!��u8;�5��RGrC�ۑU������4�@ˈ��v�G�X�KZL�Qt�i��Y��
"�q���c@�T�,����ӿYJ
��
�}l��c�X8P��|*�h��U��p�	%Z��
Ν���xY��K	tՆ,U^V�^7PHh�I,ዞ&L��[��N���!��8��f�P�Ҽ�0�Y�;o�0(���z~���i�cXj�1�c��F������7<��r:�w3i�����GH{<��b��������_��xׅ�Rp�����y�
%�e�/q��N�ᘷP�%����෗��b�k6�G=3
���D� -;���Ǧ�/����	��{gNL���fb��p����(s������B��$�y�5��)3V;� ��L׃�ȍ�X���h�ǆ�����Z�~���y����N7pr8���u�
̹2��7\���]pj/�Q�=����w��,�&pk��8z=f���O.�.��~^Oӹڦ�f�Gl���>�u�ar�>TY���8�4lU��BIF��ꥷ	Љ� T�`�\,xs5�ޣ9����jZ/�����5����N�C�r�����Y3́��tz��K�S�K�1�픪�D�+r'p�KD�u@�{���ì=�~��|S-1ⳮh��Vۯe
˪,w��n�q�Uh��m��K��Z��{۱�<����GW��
sb.��U#^S���DU�s����V����~���U�8g�����}�
�_o�$���p���B�/McP�V	]W]�㮒}��I
؋��ɻ��^Q��ǀ�����V�g����ozi<;6͑6�OQ0Ëy�6�j/����1��5'f־�{��܅'-�H�6OY#���\���|hmb�)�3*nf-O,V5���	�qq4q�X���O����4�ViL�.�ƕZ��_&�&����n�ڷ�w";֕��~�1T�S�q�Ffn��L�%o�r^��m�<��f+ف׼�]�z��Ht��}�iw����`"�x3b^E{�
�f����ԧ��޹=�/`X�`,}�}�1W �n�����[�m��aב�T���o�w��{�w=$����ZiDѬ�F ��g.�֎sš�Z���������t�B���Q��20<<+�vtz�f�5m{u��)#�4z��ޜ���/��:"��"tAô�!��7^��MD+�;��ʞ���˵8�d}[`��Vr�+��e[�A����<�r=Y�^���6j*V��J苸�j�/����v����n��	���
j���f-��:7ol��`Ӄl��� n�a�:vi���S�b���1ƛ�}�1�=���Ie��\�H���)��[�k|mr�+.�/���Z>ݝ���1�5�EdC�w[�fV@�/����b��+��-_���̍ۓݭ�vb���l"P�X8Ve�qxz����E
�U�`�sO|�eDg��;��^��"�{NQk(��`c¼@���b�L��
\֤ t�ʍ�w+$[��	����UP�P5��j������Y�͹:�����8	���Q�෶%��j��{i�^�ݠ�~rK�O���ǅ�0W��/UpUwv^�IB�41���]=�d��H�1.��Q��PAӕ��N�]Bq�&�����B\�Hx�-挳c�]lx1��E�W¬1�ָ��E�8>��ԋ�ǷW�5M�S��U:���
�-��p�'���qY��2��Xj�ՀV���e����-�4"n�0��V36ط{TN���"�.�<��3��q#G�K�s����A@ ����y�$%j數�9��g`6n�?y�U��Q	�*��q�ʳ�X&��먫}O���x�u=˕pc�^����f�8C����f�5ف�j�R�{�
C���M���Q²4��.���gX0L�j�I;x_�5jf]]���);�pd,6�B����r�S�Bv�aѥq~�}ض�
. TELG&̉z-K@��:��UU�M.�D+6�Vl�j����L�EEQ�*"#�°W��Tz�=ǂ�|qg�}����"ǝw��q`>5������쨝��6�ײ���cmYim���W���UFN`=��xv��Tc��>&�m��<9Nn{�o��,�E�4�MO �*��#^�TuA�n�po�g��&�;�h��� ��p�CL�T�O
��D=9-�@��"�w�"�ց��
�TH�Y�6�P�M����z'��=�����:W��dT怾�T�vQwm��\wT�2XE��*d��=���Q�N]�nԱ�B��ޝ�l�ֶ��k�DE�=f��U���� 1�>[���㼵t��V>�U���?�*E���2�V;��� �k�	�b��g�{��B����&�ӱ�5uB�ËAExb�5 ���ws���h�=&w[Γ�x`���N:@A��h��]�軇"��t�Fc�˘��WX�.L*�35X��2%�*��5F��1�)���Fp�	�ʗZ�6��s���8��� �����Eų���y¶�zt���W�WȝQ�*g�����B����c:y�A"������@z��GH����NZۃ"�ܣL���ʰ;s��w{�h&�d0� V�Z�0 �y�0p|b��{;#���=W����>��M�!鐊:�PW[���������c�x�ܨ'U�2o$7�s�Ml�R��c`�#Cv���ʀ�b�YTu*�lö-n�݊�֢�W�M�u��o���jF,S��QlsSx���-8�����jN=e4���j�s���wP�ם�,����<��D�i�5%���[}˴s�a���������X��g��p���셖��ʲ��W���t��D��P4��@锳j����͸�Dgf֫Ҷ�`И���-b���`o&���2R�-�4��Vވ��m^�2�x5=�������]s��X�
��hQ���/C��,j�����.��*�~J��4��3�[�u(��_$����na"�8�5ͬ�;].�~Y�4n�q��-g==}��8�}���,o+��"���5:�p!�qn4����譝�;�������2���)c��T����NRXȮ�ì��*\�]�¹����� h����l��ә3w`ܝt&N@�kTߕ��/�fP�VN��@�5{R�m�,�c�36S�ɜ�7z��"l��h��;Kr�D]��2�@��r���HN��Ҵ_*����%^~TU+TaS ��@e�t̺�&�v�4��6��wv+hfr�U���?i�Ъ�@��z�jM�����Ƞ
�w����y��6tci�:�x[�k����}��Ĕ�9��Ce^���LM��x��������_6T�1���_x�_X2��BT�d�%�[��t��4�
�6�@�z§n��q��R�6�q�e�H"\�k+\@Ҝ�WG
��z�f^�����I$z���%���V�ӏ��q�����[Y���#9����ȣje�gw"�9i&�BB�$J�u%W]r��mD��T���U�GV���)X����[n�k�5��>�$�*�B�`�ܥ\���j��f������L��L!��x0H�����1����(�������V���/� L2���l�.�r��)d�"yDN�n�3Í��GH���n���tv��4sv*��#S%J�o��_��w3�2(͸�%߾���AC���Vb婌ș���+�6�s���V.%F�+s�`�X������*UZ�9E+(�c��10ADa�T�Z�X��r&!�f\r.5�%A.f*T*�b�YPX��f+P�����[U%+�1"�2TmQ-1��2��T��ʬ1�1�Ҕ��b(�r�*�WYPUqTa��b(��6�����5R��԰�V(���R���,\JŶ��G�2�Um�*���TX�Q�� ��h�)Z����Z���Ɩ�Y\�Z ��)Ad��DLJʊVEXe�dQJȖ�c�Be�-��7��ҍT��aTZ�|*B&�
�s��Y�B�a�aKC\S܍�Su��m�d0��q��b���-"�<��rnLq�����|�q>44�bwڬ�r�JgBu�7��}̺��8�	R��b�`�(������xU/��*�p�\�U���a�+r���:)M�E�_Ǵ�����7 5ʙ�S����DU�|4hG�J�3�^9U��Y�*�2�L��R��|@!�לD�U7Y'l�#�45�E��|hub�c\>��wy��ɲ�1X����@�~<��ACH#����QR��}���M"����y�2�3ΡX���"YS�O�@|�b��蝮�{!ǁ!��w�-S�~.���d@�0���n��غ=�	��z�Q@r�M{2{�g�}!`?W�U�]�M	�:�W*�>��I�T�3���.w�����Ap��D~Œ�k�;����I2x}�/���Wn��w�Cd76�ID�;h�+��וa�f����`�����F���� �+��
�VK��=��m�ЍWN�/KT�I�����WW[vEޯ�k��ݽ��sR7˂����~ұ�	S"�8;�G -��Շ�������� +-��u�d%z��zmM��`S�ő�ϲ(��Nam��7 �����"�.�8ζ�}.\��<���Du�&����u�L����W�K�d�y58��ʣk���}uJ�Qipu�2)�>�{�Ukwn�,�wl�ت��Y��g|eR��
��T`�|� 8_��Uu�F �zN�x��C���lt<<��׶�C4n��te���YI��/B*�%PV��`�C
H�.���I�����^T������9U �Ʝ �Bˢ*��*�
�E�|.�/HD���zJaV��إ0��݈�j�]2֣����<�֭_�C:�0���{x�#�Oީ{�*��4�Y\j��g������1UEL�Vepձ�����9���ݕ��_%����S��uiV��#%�����8�[����Ĳ�s8Ҹ V��ش�t�Ve��֙�m^n�;���=��hl�I�*���Ѽ+�+�]D;�����WP�!Ww2)׹z�brz��k�o���(z��>_Y���L�����Z+!���Z�5�*�n�v`D�F���|���|N]�F�C��$^0��%e�T�F)�Ҋ�~�ˌ}p{`;g��J��0]x�V����j���g��|��j�+�.���h�@���Y5��
�|)��6޷&�������w�2�I����K�
ĵ�*l�dS��B�@��m�b��fM�^sD).6�
�ld�=���(�33.��}ko�,8����n�x0;leS�%��pd#LT*��T���;^~ǳx�0�B� b�¼=�/D^��s��FBv*�l����2�`��+G��4h�r�#��xS��=���Z���̽.Bͣ�3sz�1о��ǧ8\��O�@,�Z��Vu�Xʃ27u�,n�vu0�YhTT��{C���*4K��N�X᜚�f��hz��:d%���ұ���Eی�M�69���
�Y��z�ŀ��
�*��t�7
��w���f��^i�8��]*jC�)]�Q+&p6�u�V�UkqԘ��k汔w*zw�q5��yゕ
"�e꨼�������7���Z�}����+ �\Z�_a|q�F��Ї�CCO����pQۭqw_��b�=�D !~�o���Ն�j�Ah���@c���=�=��bT|���T��
gmQʊ���S�p�31AE.r�y�>cw��(1�?y&���5°;��DVS�U�ní����i�!�ߡɔ����0:�*��Y,[(|M���yuf�w��S�5yP��TiǗ1|n�
�5�3U���̉��-�>C���jA�F��.rA��ۿf��8��!״+2�˘EWA�V8����f*.�ߗ�{A�(_� ��كu��/p�0���(�тS]Lh(]N�	�-W=�}oq��e1���)bF��ڂ^3�pE��L�!�Ҵ���/;'lw�:w[�gG�Q|����J��� �5���@u�M�}U�n��>�IIdw�Uߠ���V�yAgՕ���E�Y�7�hu�.z�������\LM@��[��ыG�
�u=yL�z�I�(Y��x�~���,��Df����b���1?d���Վ��b�s퐪�D�jD�>��S"����4JI���vܷ̻�3�a��3��*u��T��5�nL�:S)57�N8���y��qr�[�E��z�����G�J�ay��
�� ����1f�w�7 �H� ��_*��ٙV�<r ���?EQ�C��ѷpt�Xe�����<j��������.�U�N����Ab��[Ү�������z���{���u��V ������Q	
���A��ܘ5��;����r��*��`�\X7��[�ŎyY��\Hu�������.{�3������Dvqj�� �8�E�-�3e���jGa�r�ci��P��B��fL�ṁi�UҜ��5OMr�S���dw�+մOֆ\���犦jq䮇1��0ߞC�m�ɛ���-׊��Jr�z�,R��M�F�R��蟺����˿^��[Fz��͝��;xYO��WQ��GCtmR���xS�P^]���e$�C�#LL�V�6I��_?��y�@
Ǿ|< z~C��mю��bC�&�lܼ�\-ϴBy	P��B0�<~�v0��ri��@��K�+[9�'�V�@�)���o'�
�:�4�D�p������қ,r�-W:d���]��P^ﲥց.7��_��X�w�os(L����Ȼ��W����2�x�����M++�'D%\��mGnfX�>���޵tr�X��YH�k|���4��<V�U�<���;kA���Vl'��㨕��z��j��ReM=!�0*[��G�����)Zl͝Z7�51i���J۷�jMƍm�mM*�poE:J�Y���{;���{�;�����O�B@T0��b>˪��z��QB�	]�Y�XP	Hl@qn{.�\��1�
�D�R5�����X�p�>�'�-ZN���޻��h�4W��/�����t���\�Z��ܾ�,d����G�ӡ��ɭpp�o�Gƨ����(p�~^�l��|2zw�^��uh�Y���p�^/�z���x�Ȋ�wf���9"�{�:�P� �v���iu�V*: ?i� u�2�Tv���u49���aC�p갾˘S�K�c��%זM$&xQ���w�+E�'A��k]�;�o�^�F�+�+��&Ϙv`v�%�
�^x�/���|�u����)T)vxlF4g K�t(�Ÿ�H�Pu�̔��̬�{�6��Ҩ�����X�y�G�TkÂ��"�?V �����!�ê�ug�coy.Q�љ�U����4����'�z�Һr��Y,)ܨmK�X.�+�����ϱ��n����F�~f�+wS1�a���K���x�J͂���Ғ��GT 8V��U��_���5�n
�`��bfd(4/8�ZYI��N��933T,�A�-��^9P�=�5ҝo+���!�G&r)I=L��0@^��x�EDÔ�lȗ�Դx]s�U���D+������%���h
�aF��ѓ�}.b�Mv�k4m����6NW=H�p����S��X*f�j��#[�����S��$��<��}�\0_�P�0q5Syվ�A��խU���k������XL&��`����(�4�K��#B;uV�dE*����J���[�!�j�����`c�&�8t?��`���%H9C�i<���p�
c�#��kCt��5�í�:�Tp�h��@�wf���Ͻ�տ1�V��k6s�j�H��E���N+~_\���:��^�����&�w��S�Nu�)TB�aW���a\v9�IW�Ox$K��۾:�͎�����Z�;���bJ9����K$7ӐF����`�M��f>��i�gv��o*MH�+��6�?=��Y�k}iY�B�c��F���Z���[S:l�.Кj�J1����F�I^^+=�V�TatK�(}�r�\�	�\�	d�&��\��C�`�k�T�x/�̉��*9��7P�N?t�֕S��3N}i}��U��S�`�˓.`Oe��oF�I����ա��� �3�ps����C����v]�^)�7��������4!N��Ç�UA��;+˨��yn��(�Iŷ0�>�7�Fy+UFv��Dԛ`¸C��W�K�-�.0��)�u+�0ٜ�vf���Q��$,���>�;��F�r8� |���z���㋕Up�*Z ]K�QG@V���柽��o�a�^a���.M ��	��b��סn�	<�Q�"=����J���*P��v�>�}��TV=*����7���-S����ue2�ӝ�r^T-,Or�+ђZk2ƶc6ξ��́X�#0I�5&<T���C�e�<:ϋ�>^,h�J����ǳo�S�(�3/==s�R /	Ǿ4/�/����W����Z��?m]K���y�}˺0�"���|��x���N�#�fƅJ*�e���ʇ��}W�"�`��=_k	>�q�x��43u��WB
@��T���# 0_/%�=�b�{=u\�)V���UKMr�8����뽍f�'�Wx�iy�'���u��V
P���'� �0�d�j��<J���rblv�4�ubA���}ފǙ�4�K�qh~;ut*�&���h����/�ȩ�U#�f��KW�;5i`��e��A5�Hl�L=n���Y*y���hb��EɂkT���< OWɟ�h/3u{�\�l����~��
���ϧ����
ߘlh����؀_Q�k��5�����qB�7�gSޙ�)]���=.�m��k3XR�]s�M`V�$�1�;�	��.���ҽ�o��{��2aq��YW��J���"�� �^C�v�p2:8,+;�c��5�w$�ܢ_fG��>�PeڭR���J���$Sn9��vu&�S�Z#;�C,��0�WN�<G��V�P�e�	d�K)�`K �1�W:gE�=H�Ǟ�5�C�,��9\u�f��uq��\�9 mZ�+v��z���w�����R�_59QE�ĻyՂɺυp�K�VI.K�o�2���r�4���nkW�6RZ�_Jɏa����2o�9ؖ�0 ��^Nv��b�~�h��Vv��N0��\���ա�z���q�*[`<�ݣ.���b�otJL�H.5��G�q��l;��>Z���nFoY�E�GB�[�]�D�_r�sM�h��yʒZ�/VL�q�R��J
eK,#��������*6��z���08�z ca�p4�n�u�6���� �+5f�j��Z��E���&��n�y��[�8(���mc���ݴ#	�պ���$��.6o�]Ӓ�l��p�W�E�b�������kw�uB��z�ʊ U�X�SXj2�KXpo-�5ز�N�n(,�'���Z�'f�#��^�Q������@�Z��A��5X$�ND�^oC|U�{B��4c�z^�;܀y�[�Hp/t]�p3ëq�D���V�܂I]ȱH�mr� r\�X�-��T�Mk��.�N 6��ܫ|�����jNtx+��wV���cii[��8kp'�E1Uw_T$�[�l�:�,�i��C<U��g:9GHв��"�E��յ�b3�I�3���XP�R�L��Z�]�N|sZk�eb���#w�əZ�X!=+�&iWM}g�Z%l���ҥx��Gvo.�OWb8�"*�S;G���2x�CX�L������r�� ���ײ�]�RZST�pG]|��;�8�dT�oc�͒���)��W��99���L��sD��(R�]�4���������cZɉ��&[Q�Q)h*�",�����eml
e̶�T���,����[�KhF �[&$Eˈ�,q̢%�m��Ɍ��ZTe�JV[Uq.\eʰ�Ld�,n7ĨcZµ*��U�2���Z���mL��p�kZʙh�q\-S���R�c(�Tk��ֈ�e��I��°�r�Eq�l""�#r�[2�LK����T��V�aUD�rᕑ�P�HXT�fH�RȪEdX*�ZR[��!D[�����fe�+���hҹj6Ŷ�Az����z��_ּc���Wtz��*)O{rQ[��e�R��Nْ�l�����{�ԑ�'GwOʵ�:��弳MЃ��|1���D*��R2j8lַkL̇� eک�~�r�O�dEE�a��p�<��=U4�>��[�x4��yzw�b����W.�W3�d)xFzv���~��Q��I��)�l��
NN��s3pmϽ~�n���^R��E׶��xl�E���v7l�������k��U���@@�
T���p��;9����Rh�v�L�S�yxs�*�60)�"4Ћj�Y�F
�^�Ǒ�§=^�q�8���	C�d5��Ʈ��������spn7w��� +�8�z�eϧk�b�8��^K��g��@��z'w|<�[�Ou���b�o��e٫��AF��������'_����}��0�"�W���P@4��X����H���z�ـh���'����$]O�9���)׮�R�[O���ڏ���D&6
َ���=�+�b1o,��E5c=6)7C��>j�[�h�t\���L������5�q�J(�JRv��)�Gxo<�E<����c�O>�RCҴKڣ4�im"|$�Z��r7!\1^�3{g먕"s���px��䜺ZɌ�?e)��2��K<2!�7.z�US��P�xv|�#�U��y�W�&�<���xS��{�J5������V�][��z)L�}&kj��ɗ0��A�>lda��Zi�>��0��-��L�C56�l��I�s^�����8��n����WHt9Z��ʑ7&�eX�����@(A�Q�ݔ/DR�<@�5�lu�9�H�ʇ,�c��U~|.�L��5�h�t�
���`�+�77:�'-��u���*�p髅uL��uƠGs�������;*�S2�U2��=��gT�R&�fQ5Rr=�C�ވ�v�A*���K-ݎX��U���n���)�;�θ/v��9��a4�]����ѭd]������hC�ٺ�jN���;���]���:HV�J�pi|�#�w&�*���K����`�V8)P�(��S>�BV��Țd��vt�1�Fg�ލF_�}|��a~(p$�F�+�Ї����"A~�zr�W��"�������/E�.��0*��g��4�]�望/���S�TzFl�q��,��J��~3*� ��c��1ֺ��C�Ŧ��.�fm��['(���\M9�kX�0��EX�h�+���_N�WVEQ�!n�}F����G�၎b�3M�ʬ�yB���l���>u�8_��lzХYʸ{L�x*��N�@���U屠 �Ѕ:��L`�>g4����ע��u���yA� <K|ǟ��,ۯk��	���{��]Q���S���X��F�hNU�n�i���2��5a��A��+t�㊑������*�A�V+����V���4�WHg�]��:4�<��:�+��6�-|:`t	T�Uꡧζ����03y��6��a]�����*F�V/�-x/N�R�J��5}]�͜O�7ž��EԐ�l�-�{�����n���jD֪���p�r���fh,�����f�m)x��'fiW���Sy��L��?dx|*ƍ���{�ₘ/>��_w�ԡP�:vC��WiHp�Y o)�yջg���d����jS�6w���@�/+˃�HUd6�����;[G��w5��
�2���)�2��	mx�u���u���J��G9��tך�ɲ�-���.'ƢIɜ�t*á�_#��̵�����6~K���l1�'+���ϯ�������BD�I�H�a��(��/�3���^~�~���=�PFǫZ����(���*��/��T��ף7#-�=e2�f����f���+a��`�ڧw2{�K���;���5�/Ua�n��4U���C�m�ɑ*a*�2[�1<�/��7�,y��oy�{[U�r���'�������J�	�Eu�7V�5���n�7�tԔ3��_>��"45hI{Je�&tY�����ud�rԔ�ͺ�.]<��d���s�-��9��L��V~�>�C���w��ۃ+�]P�f�;l$�_��͝ �T�j����T�%��^b�D��?c�k��4�[�D�`��N)xFzᡊ�JuBke�pa�@+���]&�o�w`[��E�9s������.�5Q�����~7�!��a�io.�pi�<��#6��:�Pe��R�\�¨��RCɮO|",�s1�P�9�#_p��ͳ&1�9�U�B��S��$ޔ�j%��W��h U��4�� >����zj�3�1r�%~���+B���㢐B�>�LDƛwG+��)z-]{C�m[T�jh�]C���^�%�a�US7�_�`�<�����I�S�8v�������E
UƫW�Mm��
u�Dhd�#�)3�����r��b�6gpR]�G�ƾ,���[�F
�V,rA�i�.�i�L���gi5����5@��U4a�څI�f��� ��Q"�PY�n��[ȹLtZ�K��xx��G�Q�K�k�H���3tz��âA��΃N�GeS:Bu�|���Z�64|,��Pp�O���V�#ŤV����~�����*z�ʫ���[V˳Wň(�ซ�\-�����ޞ���dWB�<4<;削�~6`���];0�b��_o/ɯy�-�4y�{�W��L�<�\�E�m븍G5�-��92�� ��C�|S�9�����/Mt�&s��ie�x�]i�U�%�YI��ё��dOK�.�'2��]��n2����� �,ѝ�/;��VƔWf9�tjA���7�/_d�&f7n�^��Ӏ,d��юG��"��N_;�9U���Q�Xi�g��v;�6���Е�B�9yygx8����,[�Wccm7N�+�[q<���۶FTu���=jq�x(IG�dx�z��Ӭ#[���V��C5�֕�ݙ̮NY1{�C�y��+�\"��=M��nt�V:�G�6���L�[h_)@����(�Fs�5��e�d�s*��X녦���P���UE�c�٪Û�	�Ƙ@�J�[�����4�+���TXn�������M��<�dʽ~ϯ�����D�ݛ��p��W�5�ߐ��Ӯu�jϰ{za�˷��7R��U݂Gm��p�S&ND#2vE���]db��h;��c8
m��[�^fI3�ƌ�w"�3Y��흵����ծK���k`V�M�����3f���Z�y)�X^x���?gw9s�}~��+1�Ĉ�l ����
����v�>��쌯Kr8�R3{��<��/x*h�Tf9�3z���^�z�R�>�P�t��;����Hf��3/3��"�Q�k�%\�R�+�-�YrU��E��97C�[��W����N�������@	��5��Fs�S�T�G^�VN�^�S�r��ݽ$ \�ǋ��C|�;�)�1��W��j��J{�v�>J�H�ޜ��#��a�l��U�RzuO:�k�h�bE,��p<A�:f�22Q� �g4���Δ�:�S�J)�ַc�E������Y'R	3�:�y��|��}�V@���s��J(�����u��֝��Ua�e�ĺ��f�OF�Tt4lW��2&�j�o�zqő��Y;f�n{W1��JS9,&�:i��ޒt��d�-z���ʳ�3�F'z�s�Y\k�r)�7`L	�tq���eX���]b�±�0G��-�@i�[�,��]ۙ۰�Ti����ދO�����9�x,��2��*��N:^�g��i�o��y�&�x�j�dd�"dfz�.�I���E�a��>?E>���MA�TR���(�R;w1WdR������.��_��ǻ�|�If����)$�!,�K)OQW~�W��q�K�Se����Xx����ݣ�A���&��3��Z�{�p��/{�
\7!&k5HY��++��5���f���֎ҁ��\^�	�i�Mi(fH��Tg�țʵ���8���(��k=~MY�6@�����"Oa������5�l*q�'A-b8��!d�f@��o��
*$���*��[���9j�V�ٶ���y�楚����M�b�T��@1��\W�ÏEε}+(�O<Q9�v��i"�{ �~�u���ڱ�p�LsO�ڻMF�)���g!׎謈A.TWL�����sQ��1�z�[�����Sn#�<'���M'=�\b��z��\��ts9�x%gel=b�#��I��;�E%qM����6v�_:�s�B����ŵ@j�NQ�{ �� �5\%�싄Ɨ���u�E����n��uF�BVS�r#X�F��h������M�ӑ�grIf�^u��X�e�G�	��y<�̫�s+]�+Y�˸�W�5֭�r��g�'���c��I\��ٗ��>ųkܽ��V�;���@�~�]�J}ː���	Ξ3'���Yp&lm���U��/�4<�3���� ���ȏ�|M�ф�K��^aA*�k�`()}3:��d��|�]��R�8Ϗv�=�V]���{Z�z��)󽫱�)Ɯ{i�.�4�;MF��0VM��K��S�	tЄ�كh �	h�_L9�������U���+��zL޾��M'�bR�X�-�մ�RչJ�FM���[��u[ͧ؆t4m��w:����I�t�'g�z��T�^5�,��3��b^���L^o�γV:O.;ᇫdX�Vm�[��]�v�K,I'i{tK��j�(_Pj"�yM�3�BA����m;Z@s$�A<�v�0E.���ɬ޽ϯK�������ҭe�c�%em�ے����V��З#���-�b�a��ss#�C��:9iq��G�p!*�"G~J��
&j#s�;�٩�Z#wڭ��p�Co�V-^�g):{@؜�oj��	
h��I���)��󝛇`��BJ�&���Pt0�H����7:�̋V�&�̺R��������Bb�0z�]�i��$�~�x[��U�C�r��e8bު�~�!��}�Y��v<���������=�NC�a�[ڹ��܏�Il&N�a��)z��miW�>(������������fR��V��3Jƣ�>�˺TlX��_Ύ��@[�O{kԻ��e�#1}�0V��^|32t�W�{OF��(�'	��컗�*9j��зt��up*��S�T���E�y��K�/(R�6n>�ڻ1P����ln�C.��q*@�D&�s�-%����L!�n*X,����}�͇�.b�����|�T|�nlZ�b�Q����XX��v4pW�u�9�}�)F���N������G�fqZ�����íӴ;�([ʱ�%c�Ae�`�j)�DV�]=�;��D���4t�K�}z���7t���QMwZ��nm7�j��x�xoۖ���&���	ʙ�3������Y@Z�65w&�!K-eK%�Ba(���J)���	��(:.o>j�c�s$ѡ�<�̲����lG��J��
�Q��s�.�3�v�X얻*r����L��LD��jGK�p��5.5ӐҿU~�����-Ylm|cq�*e�Ll@V�U0��L�����EDI��$�LZPQI\JLES�����Y+*�QD`��kbŕ
�Tb�EA�*EZڅPF*1V#a�DPb�*�j"*
��((�F"�QE�*�"�QA(,�+!UJ�B����*����"�TX��K"%qX1X��X��R# �H���j*cQ�DBڢ��W,�+c"EEb�DEE���b�j("1U"�"(��EUA"�EU�j�
�EU����DUV�UX�#"�,�1TUT2+�+��U��۩��Ƹ{��f�,��@�������:Yg�&�Lġ�2݅d�8��nm��~��z����;<9�<5�y��a���S[��R�7��g=��sш��+޸ٛ
��ܭ3�\葑�.GH�<i|�m���0ӓ��Nx��#`F��e6c��
�.����F�,�K�X,� H�LuDp���������"�+yq���6��]Q�� ���(�f�ۓ��p(��YI߃vM�(��+����L�ׂ�����'z$*v�o[嵕�ՊD.�U��v�fy�;�i1�W���_��Hy�t]n��g��wN���ZU9n/���b猻�ٞW�)��Q��^��|�a�q=߂w�VԷ�ܦ�y�t�Y[��XʼL/]��������	�125����uJ�9��k:��2�\�=w�ɻ�3/���5k�3�n�E74i*7�tk���ty��Fd시=I��˸�eۖ�m��oY6�]U��n2I�b3���WW�5�x��_[�︤�谓��R�Tt�/k{g:{��=p�p�ȥD:ۿ�:���8[¹��cu�V�=���%��^VB��~S\+���Ų�>4�Q�P/1�o9�f�����+l�U������o�d�yt������|�K6NL�����<
JT�t�/[�7��m0�7=Rb��6����A=���X�A|3�͚>H�ȉF�Cɬ�ް{�}Xn�?KO$����x�i���2��=�|���}��,t��<�Ҿ�|�]���HC��`t��]C�u����{���������-�]D����/
��ҷ+��תYK�Nn�7�n��E�e�'�Q�l���U)�$�{�K���A�a���>�"�W���x@�90���'&��q*����;��"���ӑ�AՊX|I�Z��u�eL1;f���5s
۹W�z��o6��2
5��kk�B��S۞�.{."�i�bmaF3s�e�--�����>��Zx�E�`v����z���Tq8��6��j*%��̋%���I��[��+�sxnm�f+J���Nq�^ �Ȼ�x1���9���}tU�%�Yg�Ok'o\ȷI97[�x�U��(���D��4XW����٠�o
����5��(NG=ήT��fY��%Vc^�v�#|�ٔk�2he^��.�.U�Ջ�P�8PF�u�wc���up�Ma����j��Pa]b���؛���*x7ax��Y�M���	;Z��#ē����j+<�9	3Ú
��s$G�E��ӵ�/#����;]�)[,�cSѬ��5~�FH*(�nRγ�ݡWT���B�#�cKyΙ���țKt��ls��r8ED�2/w�E�|ֿ ;.y\+�����e��(C�i��Sn�<;�^%x�`�i�u�_[#������G#9߹=X�� �<۰z�`	��;�J�VuTY;g/�B�s��x4T�����E+�V
��\sT2Qޘr0ܣk�Iv�4�m�aZ�g��0�C�Rc���֠X����w�s	੝��q<�(��^���3��Ny�TתyRK:{��Ye��Vح�@\�%pl�V�^|�Ӻ�כI9�wj��h#oy�g��v���D*$A8����T%w��%����w�臗ob��i�l���o'&B���8Y�Gv�=ڡ�*+Yȼ���|j:�=]�jJ������<W��?��z�z!��ڏ	�k�Y��S�&��E�T;%�KJ�+ ��[9��b���p����U�5y���:��ܒ������ ���3�2��&�΀���K'��UbK/w�cFB�)n��7�oo�?D��B�7)G�g8���,�h�	P,<�;ӱ:�zxE�sHo�ި�����F�����q�������v\�E7���2[��A�a�u�"�-WԣwD��\�7�)y��wZ79j���J�K�ǯ��bmuDb7�H'��C"�@�/^�	�"ār�6��{nk�n� ��vvK�>M�G=}\��{�5��>�k��!L#u��+yT�c�YX�p��Hߠ#KǗN��H�S*ͮ�c�D]�8$��v��tI������_ACp�>��ki1��x\Qwӷ��ކ����+��iCIiP��妯ț�őc�[����禝�w��1vQc����h���U�6�j;맞U|z�%�*S/u�"����N���R3'P˭2�����4���.�TV�o�_�g<I�F0	Gs��ښDU�3X+6�yUgCt
X1��)������2O.��ݺۿ7�۬�i��A�m��fF.-"�ժ��ӛ~۩�2;�lU{PY.�o�9�:��.E�����C2&Ĝ�w��+�2c {�~����I�Pc�E#P�rCH���(�0Q��i&|�+�t��Ǻ��w��%�;Ln��Y�֮bf.&�X��v.�S]e��RW\{��ݡ�.�S����k���5ٌ�m͠�PG#��NC*��eALn�F�_-ȵy+c�\����ż.���OF��E��FI1�aE��	����o(�S�.1+�|�f�3�QaN����/5�Q���<\�s���ݦ%-���+��3����e��!s�T	Ya�D��/�s���n��������~��kf(19:Y��<���S2T�<9��f�c�|��ʘ$T휾���\�t���p<��-n�~��P���D��{r(���W��]��T�H�3Q�py**{���.񫵺��0�b7�6�K��U��@�uicQF��WmK#֩��wC#Q�,aU~;�T�t���c�p{~�T���W.�.�۾n:0�xNEWى�{HnV8h\�3���X �rޜ��ne��f��i��-$�!w�����S4nakb8�;Qa`�Fsq�˕b�`sp����"6�]�{|�����D��?h/�n�{�l���VԲsn6��P������fWj�=$<��x��Rf��
/=��5N�M婫��J�8���4���8��<.
�ḟ�H藐�l�Gs%�!��T_�P�m���<��OLa��N����%p��U��J���Bai#\�Kg�>� Xz*f�M�?mA�I��*$1���|��8ީ �Ѩ��A�FKd�G{�s7��DdG'�Dd��&C�xggR���������cJ���$�E������lJ\�]8� 3Hj���3y1 ��,��l�=5�YV3�E��V�� ���sM�����Z87�ն�)�r.���hVJ��z�h0�{�����Z�\�M�
����ze7�@ˑ��AYMWO,?��`��^%Nܻ����J��+�T��p(����ɧ�ܸ�����}�U�lBWW�_y<&.M]���y���J��U- ��n�W����`ڹN��uJ�6�o����~�4��YԹ���vXT��1E�ʭIOcQ��B��LL����BD���fc�p)coQ�CA?gU������~w�kd+�LM�WrKW+�us#M���G�����߫A{�d��I��â�^L��Y[�I.d��6�\�Z�h�^^e���z���4>��uI,�V��R�!jbQ��ErOS�}�T7�ڌ��%w�^l��
��I]�a�^�v+�Z N�0��x�%�M�!Xe�u�����1���OW^,�\�0�����GLN[��J����zxE��i�AN��4�4�GV=��F�"ј��j${�D"��q�P�ZI<Z�Yw���|{�
�$��H�_v9`����L&R=:�c5�n+�v>�/g�x�Ҏ={��<I^�W��8��m�{�	T%&U7iU���{�'Vj�����:���/��et4%l�+� M��)�hŠh��ز��s׻.�tSU�L*�D�b4^�tez���ʲ�M�է�.�f�r3�uNrd�v��W���#�{g�t�1hC��w.�k�oa[u
�Ys	���r�����=�;��f`�bb""" �$�)H���
{|F\�@AL�=`���Ne�	f4��KG��Sxg���Y�K�{�b�@ H!�	M�yˢs�leg)��@AN�ĤF�$r�Y�������i��y>���kn�7�5�����<Z�8��Ё��z8[�d�
~��㖞_@	�PS�9"����t#��:��8�btHt�[/hЃ��K����"��ޱ	8w�����@�ی19�i��DN�`,u�[�סb?����5�3�K�7ٸ}�m����*6mȁ�\�#�PƓ����݀)5	PɊ�D��Jm3�,Ҝ�\;ʦ�����3n��'i~I��m)���D��C�Q������An��_����{)͠πC(  �S2Fc��M7���8rRX��ƫD���-�����qw�!�\���^!��f��_�����l9 ���ޘa�{�C��3���Ƅz$� �Ң�
Q���)�|�D`������#�N�����`�ME�Ⱦ�* ��nl�DAh4"g��uF  �0����
�:����d�kLL�����oy;B@L��KW	���)�@��9wd���+�u!�aH���=���J|3ۤ���?���4�յβ���6W~}O,��<T;͉O��&!��ˀ����eu����蝀  ���[�?T�2י�qM#��3���ab�ǌ� ��H�=<�{׏,���P�|���Iw�am=-@@AM�Ҏfݩ�<*]1����'b'��Dۅ�n��Qd<���HE>�#�Oh���<O-E�oҊ
o��@\+����n��]�ā���kd�A�hA��Z�Ys���"�(H�p;�