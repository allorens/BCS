BZh91AY&SYC�	�� ߔrqg����� ����  b%�     `                                    Q@� i�Ww�   �    �Qe�  �           h        ��PA"����"$��%$T(�Q"�R�� �Q)D��!$���E ���"$��Ҕ� Y�*QJR�%*EPT����8��;tD����Ң�uB���L���UX��T�:J��,�8����
  �O��E+6�(O;Mg֥�ԔHRs�y�J�*�;��ʥJ���R�Ҥy @ 1(�������rv�C��� Jm���Ֆ�\`D�"���JU)B�W�� ;���� u��t �r�R\ =������ ���J�� ����@`  )7���;�%Nx@�c� 8�ބEx 6������r�z�c� 8��(Ix b^@�w0<@\�{ �@  wϫ�Ѡ)JR%!U*�
�'6�E C�� �`<��� :��� ��x�Qp����`zz��<y�  ���%C��y��`z�(���P  .�� �z�/ `t����w�W�� �Ǣ(���@y�@d �� 0P ,���  �T�$�QU"��)x �� wgB��A݀[�� ��݀ �� 1��C���2    _|�  ��$}� p�U gR ����u���8 D: ��� r  � kǧҔ Ä�E�*%*�UJ��_ c���ݝP�� ��. 6��� d�� 1ܢ�\ m���8�� W�J)@ 8}�|C� j�U0l9 s�9�Tq �ʪ��C�@���� �       S�J��a2`����L LOɉ�IUa2`02d� =�#�!�h442M	�6J�dԔ  h   4 h�S�)H��z��� F�����P���#&������jhh��6I�yOQ���i����ޝw��a�����7���� (�'`:փ��U_��8��A?8(
+��S�@�����g����O�g�����C����C��(�EQ��Q��W@ (�ѓ���I����<�"��#�������~�/�/�i��@M2��
��CL���PM0�`E4ʨ�S2 :a:�L���U0�:a4� i�@�GL��� M0(dtʊi�WL(�A2�`�3��+�WL��2�et���#�GL��f]2�dt����L��L���+�03 i�4��4��4�atȚ`0c�@� t�ef@�+��+� �+� � i��� i��
i�4�at���#�GL��]���+� � i�� i�4�e0��L��CL���i�tʚa0��CL!��(i��i�4�d2��L���+�I��#�L�GL��]0�2:et���L.�L��@�� �+� � i�4�c	�P� t�`0��CL i�4��� �+�
i��i�t�`0�æ �+�
i�dt��at����C�2���4ʚa0�� �(i��]0�2�`2�at����L��VgL��� i�4�d2��]0��L���t�:d]0��L3)�4£� �0 �e4i��#����2 �0 :`A4ʢi��"	� U4ʪc)�  �*t�(�� �UL���QM0���T]2(�0(`4��i��
��UL��A�L�&2���F������'�g�I�?\֬z��f���QM�U3Bq�/q��<��`��1�^�&S�!����m�MN������V�QҬ�{/ܳ]�b�0h���hLJ:9���9$g���]h��fͅ/�p��MQ��Ȇ�p��7�B�z{���n�,e��ө>9��%�֕���F��"|:y)��^��S�w*��8:��S����B\Q
C��Ǯj�sݿ!�ΏF��x�S�{c�����Ƕt[6��i�䇡����]�ЁN��h�Nɣ��w@��ǀ�~�����v�X�|�k�ZVF=���d�0m�5� n��8�I�˔����V��d�>�-�S����zT�b\3w9C����{�JX�����oӀ�_��10�:�qe�%e��_p�{��>�=�bPD�C�X����+��{���4�Ý���[��[J�c��Y�9;
8�&�ݍ����[��1����:��r��p�rc�u�m(��n=��p����M	&sz�|�G���Ҍ�n�3%:�8�t��k�����6L�Q�+�Ԝ�Q�k8M�1��*�Vf�mk����[s^bʠ�a3�<��n���M�k�jow�ǵ�sX!Zr�t�_>נ`8�����^�.��XNS)l��A��'�����̵^�����s�vN��~yy��� �Κ92)ހ˱����-��1��#��#mm�ȳu#�y�n)��T���rظ��Ä��7���+	+�7M۽���l��h_n\Bb�q��B��YR�wv~Q��Z�Q��X�(�T9�=���,&�_BrN:���"C"���;�l�3�P3�瓷N�3s�Ŗ�`a^��p5m�����[�`�4	�tB9�S�x�񂲫�����[�w�w9q���b	r]6�˒�N�Ec��ҫ�՗_	�w�f#;���#w��C���^�D0e���7,�g5�)�>_v�S�a&9ӟn��H��X�lsaGOvkn�Q灒��,�=�a=�d�7Z�h����kֳL��[�x-�B�����c�j�+gU�SV��T��+��(�x�s�1ì't���цћ�I���@Xӫzf�]�gq���}�u��v0#1��m�7���V�cDp�f�!��R�
�l���`�^�6���ie3� ��Q�ɢ#-�`�h�|���3ٴ�Gt��*�;ܛXr��^w)hI�9]캟)��8^�k�e]�,������w0Ka>�Ec.�^l#��Tn� �#4q��#��	�=��۲���:懛��yvcЌ��~�,�xؤ^F4���0s�nW�����iޠr9��u����v��i���v�d�ǝ�^���Ep���3�#{�N=����%����ޓ�ރ����[U�v��`G7`�CcQ��9o�s ���d߷�d;w{#'�?	ݎ��-٣9p�v�U�v�5l���󵓼��e�vb&n�ñ���IX�u'��K�h��έ*%�1J;&�L�)^{-��?h��k��8�Y�6pI!8@:>s��5�����)g ��fJ|�����I��K"|8V��5�)}�/n��f�ۊ��if�\�:5���BJ�nM�ɛ��)��{��"�̊7W)%�tlf���c;]���Ցˠǹ�m��x���$��<���ؤz4<�Dz�������(7Ջ+���m�:QgrD--�Θ��a�k����Ğ��}���TYǘ��4Z]���db���.�{�nl�6w��yI͜�WB��]��z�/� 6\u]�������V��%`S�k�L��׎�nU�nC�nt��Z�iX"��'dB�T�ɞ�v&���HQi�h��=2�q}���0L�J�|�㮽��8c�d�{P�+��6���Zp�o�t(�3��f���^�T�q��])��C����[X/H{Mr�nt�<|�$�`�M�ѧT������o�D܉��tó:#��&�qNPh���L��qr�P[B=��w%������5�������q�\��f�)��N�v�ɺ����!�#��;��9���kq�/t�7�d�0G3r<v�Π�:�g)�Y�1ځ�CG&W�}"
\6�'����Rڒ��ҵ�2wi�Sǌ��Dɴ�2l�7O`�nއ
� �݈�+�v��-��X#���V��m��v�wJ���U�7&�GguEg41���boVy>y����{�
��'i���z="�2��ih��/���@߄լM<�.=O;�˶ë�)�:7��WM�E5���\��f]�p�,ͣ���(�ӳ:�����lâg���D ��z�ɴ0�[nK�}sC��a���*���n�j�NJ4�O[`n^�Zմ��1�l8�Y��F&�z����lF������{x��t���y����[C�A�P��s��<M{�!�Y��7����w�S�n�B=~�8B3� �M��NO��2��OnR_��	�Y3� <��"�� pA�w�j�F�:K�mٹ�AOp;�a9j��������]�i$7c�9p���9���$�ġ�6^|Ύ�M�8� �ǺE{X�O�o}&�X��MY)��v�r}E���-����J��;\�CT�*����i�ɣ��E�ݸ�LW�Z�ݣek��'�v�7��T7��3~���j��#;6��	ս�7�J�mW�l��a�oM��Ǽ&c���c�`ۍ7�4,?vV&��X/��_�A���ǧ�wh[ts6�2��'���F�"[6ю!ѽ�"����l����ϥ�Oh+����j��ȧr,�3��p%�����)���uvMH&�Kt�4�8ͬ��D��	V�z6�]�*[Ȱ����wS��*.�6M������n]D������`<�7�ʷ����^�2v��y6��9��䒼�����	��<P�4d&q�Y ܻtT^7��9L(��"VS�w�׳{xv[�0�:��oK ��^��Y���*9LZLvY���v-�f!���Y����]n�)7w.�Tdё԰�7�'��r=�`�yq���&�0��n ��P[z=5斷�\�U�d��8a��7�<P!̎=E�A�o$7��ly����sq����96�͏��ɍ9ϑ�V
�,�k���m��w���h ݰ��xК�Q�X5,� ����f��8���\ч��OP�����ߑ�E9p��Sz^��hxH��_^X�X�։��=QwW!��VU�J�,Q/v!^[��}t�(������z.*]���hv�jx2�So"R��!p����;�xW��	H7V����7i錁(8�|m��d��>���9:$�ۜ8=�7�E>�r%�ڻz��GP��kN�sٽ�q���9b�v��A2��>�{eV@�X�pE���d�.C����Ve�=�`/������-�|��Ǜ��iW��8�.˧K͚��Fs��˰h�� �p�ۻ���Ys��
K!��q+2�s�����������8A5��̣H�R��|�;+��!���OG0�m�E�
b�F��w����,�PR���sx�J\���(So�h�j�:3ϖ�G��>��N����u�o)���A�PFv�q� 7�U���.���>����Wv�p9h��Ӈ ��3�fv��>���
��<+�2>�8��Ұ	H]������ӑ�^Y�u�;9�9�����Z�Ӵ��@Cޛ�TyJ9sqiK���t.gnv��]3F�-ۮga���<	ݭF�����p�U�t���"�'i͝�T�&��X�Uv�T�5��l+T��7,&�vQ�w��A����ytZ�jf����Ί���r���g4��(����P���#�9�ԙ�v��4� �I(�=�Y����&A� #�G$ǎ���<�[AD�7:o�˓���Tݸ�JG�]��1��o\
Ⱦă�ŗr4����0���fUO\�R�u4��W6�'u�u��6X�ˇ'��5�Ҏ��疎[��ns\=M}��~l`ʤ�U���g�g��$���pԔ���P�ph��f��g'�h���U��}���oh�(������ǲ���+V=,Ӂe��@C"�;	�ڧE���0Gx�:NH����`ՠ�{�ju��tk{ ��t,��¢��v^��!;�j�>�i��I�/+
:��ٳ���h�TB���i�uó6��+�=ߖE��g���R^}�Pr�@�
`8gt'��gt}^��v��q��Daӭ�m�[ۥUi!�.�I�&1���ge��r�/XOQ��Y�N2���"��B��w��n54M[׸���c�yt�8�e���;I�N>�c�Q�t�� M������wLk|qh%���TEX�4Y@<a�V�P��A�(s�g�1���ɐj����U�P��=��цb�s�պv�������3{�ŰC�����\����Z^L�.��ަ�/9G��f��˫�x\�i�f��'Sy\�R� hw�Aw��F�6gm;Jv�^M�Ȟ�y^�.w,[�O�6��-��;5��"�<�2�(���6jZ�`͢��\9�bl���N]�]��Gڻ��U,�^I��>�[srosSvkt�R��r�Á�^|h���Û��ww�����њ��T������*G-�6�o��[��{f���j�]�	�f|4�V����A�=�3�oNoA/;�M�����Cӳn�g}{�]M�>������p�`�Ɓ���*A��"�a�{��U���Ƈ�(�˵u��t�dY���p����%k��43ר�Y��@\%��C0vv4����,�e�J�v���B��٧"5����CC�)��5Y�r�۲�p��B-R��ŕ^&lV�������\�>ג[�ǍV&�t͚]&�h&����E��:#�$e�w&���:����O�;�NQ�ϫ��`9*!c:���&�ݫ�5�|�����sF��Ծ�N����x��^�s�P�Y��3C����7��]]�9uKS[p>О-S��&��앥O��w2����8���j<p���:�] �W����ܣ ݛ�w��0��`�����r�m:G`��U�A�>�n.	�RT��T��t�:���j�w�}ve�U�����:dh��S(O��{
�\K@U@�r�X1�}�<<ua�Q�(��^r�Iϓ��7�y�5��i������v>Ҳ����$y�_0:˙��Jh廈��' :���>[�8�y	})�M�C��Yн�.f�S��mqC���h��w\(�tNGX�Xٳ6���3� s{gaLLҐ2n�����i�r
p�7�)�*om����G��J�\{4���,�����&�x����Tzw���v���@p-3��4�:�n�s��#�1�pd�%~��urH��^���#n�BWs�E��~kxsj 7� �r�&S.-�Ȯ�D�WEر�7p%!�;���������[cu��R�`Wõ>-\�Y�q	��b�����.�{�SszZ�6��_R���n�ݎK�i'�B�3������b�����g�ʯ2�w;g	3f�ۑ�ym�Ta�Ý��KpS��n��V�C�fu��~;�ɺ�m=�(>б�[�|s�=˫UaR>�7gZz-sfn.X��B�vs��P�̊>�%�6�����V��'��������)��q��)He�!]�c�q��!a������9���=���t˓�i�sF1�؛:F����{X��[p���N�w�9���6JBr�;��w���V����N&�ֵU�N���^�#Q���d;����iMe���p�ݼ4���Uo=��s�O��[��Z8▱hӄ}Ñ誚A��]uB�%�0���� R:��ԝ��'�˘�򘂨�&��:�w��]76�[�8df��zѨ�)�����H�tQ�Pb�`��pGm®�péZ]Q��EƗ�����6�N��k�_F�.����6�y%�Wk|��;m�o�X��o��)���0�Z�B����n���2Bw��ɵ���Bܼ(��SX����ԎM��eX�ec�a �<׋��$�C�P	�|�l���;�vѺ;Aڨ�Dc��B䬳��!<���_<�Sl�>�o&�L݌
�Xf�.�q�lz���㭀�����ӌ۸�
"�g]t��m2�b��s��3�K� ]�Ǽ�S�8-�L�i���Br�9@�"7k�[�)Ċ<� :<Ӝ�9̥;*4>��T���EC/� оj��m�](݃
xswQ�*�?a\��BX�x�|QƖ�z�� ���i�r��FI�1��_Œ4�n�N�kQD�d���5���2q�#�4O�`�m��7���R�Ag��yt����b���w�glP�ܴ�EK+X��4�(I�-@�P��4���Tz?4��>�Yh8rti��'�=�G=�N�l��m���+C�4�wf��]�hΕHF>���!�1��3�!��b�c����o���y�f�R��H�����8�>��O�.;�7]�P��軺���6Ť�;S'c	<D��}I��}��L�4�4؊��O"}ҁ5��vy���^;9`S*f�3i7��ȟ���\�ht�5�x�Q�҆=/�Y�蟭���=�\�	� nO`U����������s_~{{�(���H�����=_YYA�e
ER� i�hD�d2Q\�% 2S B�������T�P�UhA"�V�D�R�iUB��hUJ22�h�� �C%hJ�C!A2U�!�@)�QJ\�F��Q(C!T��r�@i
@�) � ZAiE(�S ���T&�JU�Qh
 P�D)rr%U�@)PJ���hUJ 
Ei(V� ȠD�) �@2P@�2)
@���
AP����ZS�d�����̴e�}�vk��\�jO�M�%��#�yv�͖��Xr�M��eo�x��Y��V-�f.�~aK�,�;�L�d�S2`����J�.�Kk�+!���H�x�=���=�����>�!�#z���F��k��	���5m�K�r'��4f��aXc���$�H-�[�jl�C��cV�o>�7���źi��p~kqtĴ�"߀�0�����dd��]}�v��@L��!�R�Q���x����ӺIӻ_�����}�����=u����� ���}����_�<~��l?��������~���>��w�k}�}Yߓκ3�����`�hkV�`]�u"���go;�9��%�NoG��{�	 c��`��[׼������2���t�{�kۢ[�x��=�)���q�8Zy7��^�٪�G�k��CA`ZU,/OP�G"�˳��ֈ{�Bgȼ��<۪�!˃��4sK��[�3�~!�t��n��Y���|�S�<��=�D��(s���`ߥ��>���X`�*n{p�d�"�l� �H�J�YO��	:���s��vn�' V���M�y�=�|e�a�U��������üVM8m�v'rM�%z��\wV]͞ƎJ�vɂr�^�f�C\��tkY�'O�{پ���f;u�K��MH�?��^��Y�QM��U+�=�cۃ�������>V�L;��� ==���6ƽ�"V���ȍ)v��`��/}��g�����V@�nM[��4V�+�f9~֤�L��7���^�xǆ����������&7����R#F�!:��%���6�NzW�;���>�{y��ͅ���T�>��&�l�����s�wP;���$5��
]�=>Ք�͗/{r��z�ޚq�N�7Vw��]#%i�X��i]���N�3u��F,�S��)4ٖh��ql��̓#�'Q�"{�Y��f�t�		��w��^�oG#�u?��cێ��������_,��Ǐ<x�q�ǎ<x������Ǐ=<x��ǎ�<x�Ǐ<x����<x��<g�=�/=ߎ����7���^M4}�9�}�������`�y}�Ɩ���O&L���^*�g��&_��@����f��hv���}��Oz��[Ž��`^��������x{����{�y)��Z�2�m{Q3�dX��.r{r�K�K�4�;�y�}F�Լ9�FS�yo��kn�*��z��������b>���
�|��Wft�2�J���������0�WQ��B��� Q���xA��产{�,��%�m=�ڄ���Y7W�iy�z*�L��i�]��/tͻ��n�8������;�M���1��|��+���_��ڹw�b	ѷs��g��]!ze�e��{y��=�>Q�#μ�l��}w�χB~�;_�%��a�U�2aw��L[��5��r�Ʌ_z\Q{�^~�~��=���FО��{&s�zwar��q՚���5���V��l)e�{�h$y�_��=w���LQ:���t���9�W���n�a����\k����g?J{�+���ϑ�ԧ㌖��A���ӼF�ϳ�ۋ���s�l�u� >����y�5ۑ��M	�����1���}ؽ�"bNָX����Wo����=��{�5%g�/l�~�{�䦍>m�^�|��V������}��f�o�h��#5���X��c���u�����oo��Ǐ<x��Ƿ�<x��Ǐ=�x��Ǐo<x��Ǐ/�x��Ƿ�<zzzzx��ǏO:��ߟ����_J���^�� �ϵ����B~u{H����]��ˍ��G�2�ew&M�̲<�qӈn����8i]�:�F�2�<�꼪��H����f��t�Ə'�p/?��l�=������ٵ�<��P:s������w�}xMˏ\p�wP��ܱ�G�od��E��S��Ϊ��MдvN�j�˘����zdұj��m��wG �/���=ѯ��+Gr��<5�8��o�BD�Ἢ���'xv���9�q�Gn���Ú������/8��ǅ���.>�����ӻ�_j���x�ڱ¦�^����W,s����>+�G�=~�$<����&�7�'���B���U��E�aKw�;�"ئY=��|���#uj�e=�V6��w���y�o�c"��=���}�6������1�m⽳q��3���'��{�D��lCa����Xj~�Y��.(r�);ǡ�B�1I�[;^�p
ͬ����}p�p `����\�-v�Y��{��`�o�Q�5���i��� xa�{�|�u�s�)�.
mOӁa��.��SH]�KCz��]1�w6!��3^]��"Bj���HiY䮎�n��ʧ�{9l:�u{x���{�X (f�Ni_%�,i�<{�A���X�Ԣ��+wx��<'����,+��9�U��(&��^?���<x�㷏=<x��Ǐ><q�Ǐ<x����<x��Ǐ�x����g���������g�͒-]ZNβa�<����C��Stuƶ�����A���r���:�y��c`�r/n��E��{��h���� q�d��݋صE�O���>�㋭��~�o�1�e�'�L��Ȣ�G��i���Zy���A6w�z�́T�aX@۽�m�9}�P��/,�^\d��R�O�����{�YR��힙�o�(v�z�U��'޻����+��{�8sx!NotL�B�j�j7=g������N.	o�i�>�����x�^9�\�9��9y��*��d^mZ�iU{o���U�C(���Ə�,��dΙ���;�y*��v+�����Ԫ��9}V�V?��f��edYop��jίC��|��o��g�|�yp�:vr��:����'}��rs�{zo����h���3�U�"���}Nݙ�{���Z���&O�oE{� �����K_G������:9&�x�˒$�WD\ee094LFB�����S��h�����==��lvy(����ޭ��cܱ�C�l��PِpoY��u��xxC,�����F��۱��,�ێu`�#��Z�R͡�} �M�5��wï<͘��	�}� ���r���Gݶ�ҋ�3�r�$�Άz\�t�u���L���m�`�{{�S��p�\*��|�[Lg_QV:�[�sϞ�뾧�OO����Ǐ<x��ǃǏ<x��Ǐ�<x��Ǐ<x��Ǐ<<x��������Ǐ~;ͼ�]~��3�|Z�sh��Q�l�E.��
��{��3XCJ�:x�~���	5$g����J��{�8�Nv-����V�4Q��x?Q�j��+6p��u�~�5¾�sc�xnE�<�D. <$7ssh�i��4��>�K��/{��;���`zZ��,����� :=��dاd���j����"ӿx�-���������n��s	}�"����`X�����|'�q+Ӵ��������'(2�˺U�[�����ܮ9����
�u�yT�{%����7}���+����q�WNOCa���PY殍���C	MqQmY6w�o�{�s��ҽ�P4J�=�K�+�^�$��Y�fZ���&�q寮&����a�v˧�
<|�����xS�f�� g�2ĥx�D��P�#s�����!��j�>���FK˳}zM�^{�M|t�c{�����}����>E4#�kh����^�r�K�n�)s��۴=�{��gc�(��/R^Df羚����?�~�.�����vyo��9R��7 뗎��}��޽�O�H��\��NI�giܹ���>��:��n��.Z��������lyP��C�G�z綘i��@�\�G���w���<t������{{��h��Tf�(L���<N��Pw;�λǻ���Ӯ7�<��@�=d����3L�iľN���E���޶���q�;��������Ƿ̨!6f���bHQ�O(�=�E�����3�� i
<2��/;�?��=9��ܝ��.2����!��l
y��c"��N��у;��ܤ�C�0�$�����D�c��G2�3�"�ۧ�l��I;�,�c���g�l�B�Mu=ݙ7'�K���I{����>�-�Q���m7���b_x�Ð�U�n�=��i�L��l��wUYA�X�=:^y��Af�'n����q�"3�i�Y������e~]�zu�X@i��]�OO)V�{�|��	���[1�ק�ɋۦ'��<��^�u��<'s߲��[ov���,�<�D���^�M��������{y��ޥ�`���;�}�{��Dv���m�<n�������b�W���0��^�9�Ë@�;�
 wl���@�e�K��x,6����3�5�����Wz�[���=�9�g�nZ�¢�o�`r�4�Y�A��>���bW�S��j۩��I�]y�H��&���>�Ќ~�Ha�%o���=�;�ŏ{��s�l���h�:	�Ƣ��7�-�'4ݬoE=utū�D״?B�Eg�N(���fv/MN.�O�\m��L٫˦]1'�v��[�,����^iǰ���_����ϖj�o��oC��닂�s�4כw���:�!���˳}[x��M�լ�;q6:��^|��GOLn��U�����	�}7M�T�y<��^lc9�:7Nx�s0v���A�m�S8�c�Z���|U���~�w�.����G�L�܂��g��Ƽ8EG_w��;�s��l�K��<���W]�q��9eA��m����9g�4����;�Z���0f��6��ڲ-Ĳ�nuo���xèO���A�{S̝�p2��e���o�0a�Gq�gi��ܳz�%�q���gY��ga}<���|��z�z�vz�<��de���_��;V[��q��֍;5���u�]��|������#�׫��hYe��O�������՝����_z)����徻��W+��h��'��띷������:����^+�q��ɮ��9	�:�%Y�V�PGy_{v���ɛq,9מ� s/u�l��6:w�������I۾�������[x���� /ys�oD��,�F����j�˳�^�ݾږ�]��>��[�պy�g ���m���^�܃�nJj��OI-zr�xǂ�q#��{e��g��R4��ۧ��[��N�x�"�����=&���Z�����S����$��>�w�D5q�u�;�vڇ������p�	x��jq��!��L��
�DT6w����}������}4y�Yp�;���jլn�.yg���5�W����y�^7�G���x��ڟ��'ⵅ�v����%�9�ݳ�3ۊ�<��wG<��ULxwY..��k����6��i��s�.�NGK�#�}+���<볰����y�L���GS�딯������D|�|0���p옽^����K��Ǘ9��`� �`R5���_�w~�2�����k^�g�f�z���{oU�t+����g����cs7J��x\��Xes��]���5x_�����w-�F���,/r�y�ҧ��6`(�~K=��A,�퉯���N��z;<l����6z笋zo��~���(��zܵOj������g%�����H;�fQ�v6�,��'BƼ2�̑���踪�F6|y���ĥ;��$W��p�;��,-���
�en�?`��Fw���{��X��j+�*A���	xL${υ�^wS~��|�����L����|.т�*�t� ��;%��<A1���sq�{'�s%�y�p|Y�,�i9sd|a/����s�BJU�$}��oP3�繼z=�����7;�ř{��?o,��}GY�p�^#Wi��}9l�+/����<7�hk>��϶5���ah� ��}��n�o����x��Gt�n���Y��%����	��Wwf��b�xp5�;=��L}���<��v�>{����'\�O�ji�͛w�}|M=�4���l���f�i���hxs9��L���҃�nh�H��Ic�����f���x����wQ���V�����L\}T��#�gaG�O��y���ﳬ$��Iv������_\�ț����w���7�{�8����ǏG2s�<~ݞ��7�k�o8������<���V}�Uyx@�c��&���G�X�hH0��)Vu���=s�zo�uՊ}ux-q�*^��1i���֌L2ċ��K��9�g������#ZT�)���L�$
"xߏ��-;�fx�ݟc�/�͎��`��w��d�nfM�Q�wN���y��{��g�Ǫ>�{�{b����|�`Hpx��^�gx\�C�=۸ހ1���
��z�;�<��~-`�N�x����-�q�%|��c6vr���3�����~yE=��Y���s{n��y5���3�>I{�ˎ��~�{)8��j�����⢔���
���
C/*���Z���mT�������{~�%��8G����>�u� ���}�;���u=�E9ٵ����]�׍�ͻ7�̳0�D����sW��}�}���r�yy��?M�b8�� �S����̏��z� :5vk�]TݞI��Y��p��0!��޼8��"+��/�6o��ٚ�h��`;	~�v��i7q ]����{<���%�{Qܝ�V{�r;����{d]�S��=��뗇&)��:��J�G�������!�b����ۏ���{/�;K�䛌h�ۛoZ�4}Lxf�o��AN]�����ED�K)f`{kk1�l�
(4�ö����\�_��w<\Lդϳ�n��2�x�M��얭���i���K�/t=VE���m�E��W���~D�E��+�û���@Y<;vr����[���A94����n��y�W�n�@v!�vu����A���S��{����Ӎd�0���mp�ý��W�Jb����'έ�x��O�v��u����l�{������c�w;���%];�J�����m)ҋS=����Y�7��a�Ի��$���S�?f�����=�����^��w^��J�j���[�JO�f�O�*YyJ'��ac���ˎ��ۍ�j�����dָx�^~<���˧�5R-O�-�皳�6����9��v�va��r� ��OO�Dڧ �0ϝI.�'Dl�m͘�U=�m��v��ww}q��Ɨ�"wOs��J��;�On+M�
0_y�;>9[�-sŞ�N�s�r7�)��5���˥>۾�����`v��]}�(np�����Q�4�-g\�k:'��}?�~ϹQQ�*�������>�����v��!g�馿�"������N�l���_Ε���UUUUUU�=e+3El��Q�j�۶MSA�ٴ���Y�*V��ֻ\����l(XKHl�e�6�X
\�/X��p]�uL,��,*��.�J�9#��B�b�U�+	k)��X0%@�Z�1[hԔB����mX�m��Hެ�Zb���aer�7(V�+.�-�k�(2d����Ł�Q�2n��4���(�E�(��.� �a-fk(�*�t"3M��ʹ%.��z兆�Kıe5.�[3��[�����mL���r�,�4Y��t�e��J���31\�Q�.��J]7mHF��c{f
�[�%�d�b�6��C
A�X����Kz�:0�k���lK[q����F�եXhfif*�L����7�k��"@-�;	��vnj��X5��Hd`�v�8�"�u: D+����m������ �IjۄE�4LC!Z���\�v���j�X�����R�HM�. �u�1�!Y{,ue�Չ)t#n1	A�٦��!N��B�e#Z���ke�-�Q�Zhۥ�0҃�)��j�Mh��K�-Y*����͊۝�i-ը�Z�a	mvH�(�1��dT��k�
��E��`�*�c����nv�,�[�K�)i�+��b$i��jZ�&�����G.6��U����C8Hk���1��b&�I�3��1Cִ�f����)p]����\7kZ4�hc1����f�A�ŸUGa��J*gLBmKRZ:�P,�]�Ŵ�m�4�IRb���4���R9������F�3PX�R�!FQL�Q��E��"�M
:��Wf�9�
��C@�`�T� WLGZi��k[-�e�tH$X�Ԗk�Һ��%a�E���4�I�1G0���Xj�*b�72�<���af�``1f;Yh6[�] ��470�[j9Xש,r�(���1�T��)�B%�m�5{(1�2�Ylt���[�0Y�� 2�A˥l^�(���)�.�8�ne��tc�,(�љ��b��R��V^�ـ4˩y��:P&�f��ٌ7hfme��c		מڔàk�� ln�SYn��p]D"CJ�SF��B��j�,,����59�����K]��a���uj0�%W\�n�v՚Wu�F� {WX5ZFh�����M`C:e���h����[�)�Ynm���c���mf�kŖ!*��4�cb��)Z:�.��$е�^G��-�v�U��P�a0�;;B��������v��
�&����ׂ��,sb�0B�˗#F��!���� -�e��n�h,�f<9;B���ͽV�����[{A��Z��F%�c�rfn����jp�[fs5��le���@f��H�
��Ԃˈ�d��e.�س;Gv�ii�(����4�TG:hb(kXf����-2FԍttZ�)��uK �f�a�s�,��e���na��v�^��5�IBI�����+6f[��L�])P��*LrL��]CZl��0�lܶ�In&j��@��=5LkJٌa�Ѫ�#�^�+���Z:��4)���!.L-�9�`s[�)+���HF&̩�� ��YM�� R�s�p�U�����[�u
ΌHKM�:��l!QK-%#*�:V�����Q�e,m� 8�64"GGE,��F����Gii�ܻ^�q�	�V��k�IS��#X���Ĵu�jF�m������TZ��jh���.nb�ۑ��m%��dU��[QMYYL�����7���
�`�r�Ys2�\�+�u2�&�Pn2jqkH��dٚ�^+3�����n�1r2�eJ��L�1* ����-і�M����Rh�]����2�F:��umw\ ���\�L��f��`��YaB:!�4�VM�]�&�)�h�06��Z��Kv�6���m�i�m\�h��XU���*��Y���ۑH���1vRܻ`���-�	ԅ^����]
���t]�բnЊ[niZ`�[�rA��e�i���D-�89�FW���f)Ζ�X�Z�㉌�l���*j�t�kr`e������
=^���4�Цҋ�K��h����m�P�����B0̬�b�7:����� [��4u��&T�!�#��af3u�
��Mmb��.�Qc�����j
��ɬJ�L��]u؄��ܦ�]��tI���`�M�лF��l�u����ۮj�qf&�mCZ��0��ZIZX�p1��ݑ*��Ԭ�+qe�5�0(��2�b���k�"�V7`!h�u]q�.�et��ƘF�dLʻ0�W$�ؕ�:S7h�r�fgA�tt�tŬm� bk��B��-u�V����K%cJh�v�i�v�.fKq[���YA�:�j��2��S-3�0trY�Pc0شllo6����.&��݋�VW@�Eʡ��l��e���؅��GZ\��d�!�T����f�#�<�m*:;bh��!Vf\HK�j�[��:[��:椆P��Yp��@�C��`*m�
�����ۜ�6톡�A^�"4p6��י�ۨ\٥g��e�.&�6dB!36�r6l��.e6��	���m��˴	f� l3v��JL
�Ytf�;J��=PI)p��e��tƙ�;dL��eƎ��kr�@Äs�J޴��E�l`��K�8-�8���B�j���ĹW ��k^����Ƕ�Mj&�l@���j��F��2h Z&�	�i���TB���i�k5��Ҭ�����9�]�[2nɆ�c���Ӆȳ^s���Jꂹ�h�gLƭ)eꉇvt�4�#)F�YM��.D,��0,#��j2d6R�x�0���MI���[e�9��4\���,�SQ��n���1�Á��6D�J��3kah�$9�SG�0V���ө�c@�D��G@,R�5d�R�-�k�f��*iGG1r��-,$1��44�ڎ�l��S:�VRa,���Њ���2T�Ɂ������
lv3HL�iXLck,�5���ƱW��,*�ns& �Yi���@�i+E֐�3n�B#�.�k.+�F�4��5�.Ҏ��i�Y[X��� �hح���%������ҝ�Q��f�f��m�b�失&�Y�2�3ںl���]�X$�ř�Sݑ3��Y�� %+4d������	�:02�Q�f�t�e�k�0���L�0�Єe�؛L٩�	��2ʸ�a�d��%SLJ�F�0-ķ5��n]^��Q�1+M��b�l`�ȅ�����K;;Va�,�B����LG9{d�,k�ю��.E���!���l�Fչ��z�*���C���60LP��8���,[��]�)n�.���%A�6e$�FXݥ�*Bѥ�Ĺƙ�#�9G'5�*n,�M���b�GB6�kvt�X��LӈV�zX��Gm%��Y��if�И(�ַZƗX�z�	
��6�;f�P�#�D�6�٭��YU�i.���-�3nTҤ66l�V��7R��U��dҵ�f�Mb8Ó.t��,�u����4�h�j�-"��]c%u�t����X/d��-��)5zZ8չ��e�C3B,2ZM��,�Җ���V"ҼR�r�@�q�	�Gn�n��j�U�Rn,���X�V�u�e���,���J0)�d֩mҺ2����*����36�t�q��ظ=T���.s�l�[#061�A�0�ZgjD���^�&��c��l	���U�d�t����v;f.����ثU��8��p�T���.�9��R��ֲ�
hM��ku6]��&������Ͷ]���2�F��m)e�T�K��ֶ��6�P)�B* ���f����
��[�-q�ɩ]x�u�bf�H�s�cVV��l�pR�V�4˶K��^��p�P��Έ6͉P�U��
��K	���bhgb\�\�af�gM�iY�FE�����2"�����Z�W.ۣ�!.�Y��7�&���i�����D��51kU��4�Z�mb�,��m0�5B*�0�t�fń#�:�fױ`���4l Qd���5�3�h-�5�a,�������9nj�Sk4͂��,GFؠ��#�J�M&��nzܐ���'Sb�Mrd��SQ�ulы�$n�:�۳�����H]K�4a �$�h�81J։uZB�l�.�p�Z����õ@��񍳵u��=�B��c`$�d��d�n���U�-�[��
���#4�s4�f&��ȑY��u;-� �6F�m��.RV2�Z�rRQt֗��GT�2��u�c�L�k{i�R��f��8��`��ѡc@ʐWFݝ��h<W4P��r3%��GJ��A"��v��9�`-JM5��܌)f��iIx14�\�Įf���n.�j�vMJ)�M1[2�Z7C�0ہ�IHٌ�q]�XV0�0��b`օĸ�,&c
�M��hZ�;3ۈ�7V&4�גj��f��v��-�CQ�3$�@���LG���H��řMMf炐��2V�&��*��	�L�gsЄ�QԦ.���rԷB���j�\��'hjm���v�6�jBTtU���bhG�d5���ȭ�0���.��-%��u�SS��%k�:�Ͷb��e8<$ҚX��ٰ�`l!��٘����f*D�!�����\Ř�ux�V�& ���E��3a��k��l�4�GQ�l��15Y��P��t�ˌeu�L��d�Lk�V�,ݕ��B�+2��]�C�6�x_��FKqԩ+YSHm)qphf
u��88#�?:�\8	˒C�]a�ZSm,��Xq�a'UDN�q����gl��5�3 �"�����k3���	�i��9���v�LIFmǧ�nݺ�$������v�B'L՗b�!N[n\���%��2�8��۷��qLG�1�9�I:m�qZm���hrt���%�X���C���N8��|;u�'y�DfYP�v�r&wf��.;3�H�3�9͛�:�$f8����Dp�˙�:t�ąm�G3m�N��;��޶i$�����e�X��;	��ݶsZ�Rm�ε�pə-;.��6�Al���T�Q��+-s����GA��e�$GftQ�n�3s�Da%#2Q�bK#���vqI��q6�Y3��֙���C��faCT�fzE_����v��2i�9�kq�#Ya�[,���s�Q��16B�
�]]��kM�]6�pu�a�t�	X�l���/Fn�%����8N��ټ֝|,��,ۃg)�+�F���`�\�����V�(.��@Z����ƥ�5"T�j�Ѷޥhne�D#`�Mջ��&rj9�)Av�Ժ0�Ҧs�k����R,�-;�l�&�j�0��
U�S� nB�Hmf�kԫ��ъ�Σ���
�����L:�E[�ݬ�3�!��g�,Z�%��BX��,t,Ќ&,[�Q\�k�ԍ.�n�h�42"5�h�oQ.Z���	D�j��pH٭��y�<�a���v;Q����[U�-��6m���jv�nqύ�`���hb���hktB��e+1:�靁k��r7%��@s� ƒ��tj�w2Z҃�ņХ��i[.NA.P��L�2ʱ���������%Mj۱�fj���9�iI�
(K�� �l!tN1��WL]�w0V�]i2ȓWk`�-������e��FJ�	�<&�7���Б�M�-p�J���$LC�䚂S1���,bZ�cwh�hj��Z��&e��Z��\k�	f��똌ݶ2�,I6�	k��2�R4`�e������m�*�p��Q�E�GV�]�ڒ�����ٛR�At&��u��2�M�����rٹ!P)X�\���t�D���j����Fؘ���Z�E��JV�'�����v�`�:TMMf��4M�s�%��CeF��F�	�]hHKf��nj$.�))��n�t��5	�J�P��qq5HR�9��nд+���WB7
���R�\�XKT�.%�b�S��c�fd�ef�E#.Q��&L�4R�ɪ����ڍ0;mDW��q�6z�6�6�Ff�l.q�HX֛fgb��R��k B��W ��ni�]�8Y�P"(1���l��D���)�=;�����W�e��B�S�`F��6���R��ŉF�V %����R�i,����,���ʖZC�V6�X�5$)-��UhP��`B���(�m�e�ʰi #���Im4=�1'���b�9ox�Z�@ C������e�$Dki(�,cD�!QZ޳z��ֶ{gz�<w�����ԂRX4 ��}�~�&�7-����K�H�H'�/-�[-Ý�:u�E��S�`�m��7�z$c�E�`��uT�4�D�݋�Ǆ�t��5�8�I����I!�_H��r5��jD�.�#ļ����2�8a�B �m���"�i�2���c��6�p �����Lˆ6�h�ik�"*2=ĂCU>��"9U�69ֽ�XH�/^M�E^ ��V�KN ��<�3 3s� ��h^�D۠f.>�����Mf<I#jv��-��<&91�y������� �X5���]���Bf�8`��c+L�d.bK�΄��k;&اp�٦j6=�66#ju���Zѯ�1������UR����Đ+� ���o�`p�w����GS��?^��_j��'�W��{;��;�2gT�'{��*2Fb��*�e1"�F4�i��������@�$	y����;xǉ�lwyY�ȂU ��Dtȸf)ػ)�jq�'�rq�	��SIh�q4����:�}ʝ� �f���2�8h���Lr�S�7����c������ �sn�����}YN�7D�Q�q �V d�%� 	��<{sWeʅH��c���� �N��刵�=S2?c���W�Kjf֒�Y.�"�v��F
Bb��bRR�ߞ�}�Ʈs����
�l1�A��B�ۻP.��ȸ�3tF�ǀ~�^1�~k���wH+���4�ˉ-���e�6�X_ag'A$�sv�A���հ�:1����L�.�S���р��{"I���	>+�<tՇz�������iD���
k��v��B{�O����������ي�!�_����nd��G���Σ�t�B⎐|6�#��ڈ���3:.�F����٘ �����@�Ǩ�I!�_NY����ֽ� �F�����&N؜x�Z�f2��v����@$��G�O�q��!0�w"o�o�����F*��@�c[� �-�#Ŵ��Jn�9�ƫ���>�ˣf������$̨�i��,��a��W�����D�Ϗ�������1���?{o�S���w*U'W[5.'��r�<@>$U[g���K�72i�)�Y!�m��3"�;8`�2��A5�d A6�z��1�vv�	#2��Zq�|��d��wr�̈.Ί���Fjǂ�W�j"`@%��	�ڏ9y���;��.la�I��S��e;���� �M�C2~|�9�	r���߷�h�w�^�=!�X��zQ�Ӕ����X1��=r�+ɳD���\0d�(��j�����qX�T�)���CY�b	�݈��|0H�m@�>:�q1������j�[��mlK�Z��T�besJA���ܛ5*]t���
9��z��=~J�QNK��z-v�D r��@�=�8�oqA���8՗ @$����I%� 3I0p�Y�*k^bx�U��m�Yy(gz$շ�5��A � bo'`��Oo�Ɨ��q��n�N�Z�!�����oi���,�)UŖ3f���|ӹ ��u�����2wt�g�Tv���U�I[��
����N�ӈ��&vH/���e3�~3���+�F$��_Ϲ��{s%�+�����dS�N�ӈ��C7i���fDP3��qYX��ʝa,���(�������Z���3H-撖)u�QşEewcU�felSV��m6���>N�Ės��)q�"[��g���)adك��iN���O<꧊ &آ�˝WdKE�@��J啚�@����K���&+@P�ccB�C2�+���(iL^���)�&-im[f걸C^9����YX��P���s�p7f�]лV-%�q�
�@��:�sqR�Ț6��TD���j��p�Z�fh��f�5��T�k�GpVSY�\KTv�΍se�]���Z�¡�n����Sc��iks�|��Cjf.2t]�w�NSƠ�o&���o���b%��f�`@$����c}���$�Hӥf����������W�ި���	�e����I��ٟL�M�q_ˬ/��Z�p{�	�N��!� '&|�fdO�#kf ���x�nR�vx	 ���O���
���wd�p��<l�6�5Q�[�9�Uz`a��q�|O�rb-9��$l�֙�[Q6`�[�7������B+JH�j���1����{S�'���j7�c1���\�x����1:b]��Ac��#�X0`\��rE�����Sf�
im�Ů��I�B�6Ʋ���%�N]?�!�;WN4�H9�1������Ҧ��F�z '�/f�`�-�8p���Lj���񝚸8�#m�ww�͜�le?1��p=9���&#�1Y��55*̄�zrV݇���;�b��\�g|�X�)�8Ή�J2uR����� O�&�� �w���Lڥ��C���c!z7*�Yt���b���1~-5���f���Tfԭ3�]S�$w.`@ �4���%/f��.�"�ó�Y�vMm��|���ʼG$@`���;�+n�5`��ْ\M�bA{��|�Ԗ�HՋQ�D��3��,w�umѕ��c��	%��= �3n�@.B��\�A ���y���t̃Xg2�]#]�1д�45��sXG�f&/�D�~��~}�\���r�<w��L ��Ǐ	��7�ZY�0w¿zyL{9A�?7����}���+�F#�C�?W�g���r����Sv��K��$��{ $�26�@1��]�=���C���c��.�+n��9�{$j7@$�J�& ޚ
��^f�?�ߞ���VJ�'娩�{ws�=pӔh�X��dЫ"�
׻��Ui���
�QW
-5�H�K^���d8����b��8`��p��5���j"w5��p�`1�q��ˀ��"I��ۛ��44� X�My��x�qhM�EÇg�τ6D$;��Ak��=�oKN ��f��O����s�+49X���"٘J�b��ʦØʑY���)3	��f�!�Mr$m�_���U��c�����PĐMk�/��و���U6���J������������B8�-:��'kf �b1袖=^������띸H7�u�}��e2*	�z�pptQE�ƽ3�I˻�����V���܈�H�>��whx� ���H$���բ�3�v,S��5DEN��\>L�Ee@<Y��@$M]�{����w���dR�7e����Cz@�DŲ ��y�	�d�ir�5�Lgg��
���(��~�^��4��4&�1�Q��OCN�{6&D��`�ى-Y�tiX�b���^��>	��[+���!>L�v�"$)�\,0�㫼�����OWC�oR��ͪ�x�RR���ցv�{V�XŌ5e���Bo=O���j1�B-[�i�W��ǈ$��}ׂ1�rcc+��*��� &���D1q��"��8AO�~*��mOY1���I5�/�-�^ 1��gv^��w��-��B9���@�>�G��*�����@/�Q�Vѻ-����̦Ǭ�#W��|׀	��f⎤坐H�L�k��r<������B&g|�)�b	 �OV�H'�;pbT�+��n	:� �G�ذ˩�iEw����}>?��d��&Y���<L4�D� �r[e$�_ܸ�-��RkW+;�٫a�{B�7�C��pV�sv�v�\:l�5�A�x�����(���ǦW�"x谽��tڑ��C���}첎ހ�?��%%|�m0A��Ѣb��hڶ�1���,]�ds�Ѝ�R���\�����95�nƛ1F:G��fԦIn���n����ݛ��U͊�ͦHc ء�,eGUu8�Aiu�
�`d+�h��pK&��-�b����J)�m32���T֠�����jf�f��	������-�HE���J(�K�WK���*,Һ����5�5I�a�;$�MJ�a1,�r����m���X�i�@P�%�j+��g�с�;�8`��p�Z�#�A']^G���K�;p#�}�eY|O�nL���)�u@7�q��EÄΐi�i�H��-1�7~�A"]��PI#gn���4���ϝ&��_7{f��pjđ�'�̲`1"gu� �f3a�$�5T	Ӷ�``���ƽ�Ԃ�j|?w���$�2圈,�6�}s[<I ��׃�V�1��5R���d@8���\�w2�������&��C��z@o�,��� @�ϟ=y<O�~W�:���L����@����+�Bk�s��p��%��,�$�f�}�5��1�:sb��&��o2��A�%�f 8қ�bm��m!@�ָ���Xp��bY��uے�J�7s�o4��:O��Ocݵ�r��p	r�-�]Gh�H��@*�4f��(����n�dK��'}��LIi�hdr�\���U:�����	#7f= ���U>2��6��mī8R.&.�I�w�A�ـ �O�I�������k@ �&�x�|wv^.gQt�Ag�C��ZS������&#a� ��bI
��$��M^��{i���P�߿>yΛ��X�e�d��|������Nn��Y�����	 ��p}$^��&����ߞ����6�n�Yv��nX�M`�Z6��4K�ePt��rhT\�?_~��j'@������5⁽x��o��)��E���Un�z�2x�A��x�«Ԇ��)iB@�o�@���~�r�55��ϊW�	$|}"�%X��h����T(��H78�
ɜ0f%�0ƌ�>7㑭�I�������s�٘5��e����8�.�(��(�+n�չ���O�}�#�n{��~�<�l��`�U<<��&�,u�?pޝ���**��`/�� ��}wZ��cK����X�t���7�z��Y>��3�6"�x��������v���#;N�rїؙ6�㔗�<�>���-/Iӝ�~���wǢ|F�%�w�NӇE�)3|��Y�:��tep�����&�Eu�kM���D����sI닞o_JGX�W�Q�\���'�N�z�"�bc���a�z^��>>����W�����;�E�5D}�����d�G;ŉ���ӣ���9��V�h�Q���3�v�o\CƜ��^�9�F�=4}|}������(]lOv��U����e�vt��ŝ������C���/�_B�l���iM�xt�� ķH��X��=��|]7V'}���f軯�~����G�O�-�pVNI�mWǲ�S�ev��<�[��bj�~�zp*����[��S~������x�k�~���
.���m�0�d��7K���d�ӳ���L	\q����l;�or�e
���K����ޞ=^ױ/{#Ŧ����{����S�X��i��ov����7'�3��;{���W^�r/n���j��~�z�]� ��F�\~gX���xw�i�9��L�A��>���n���B�}����H��3we��xȸ���}��.��I�s��ŊM�/�l��m���s�����ٔr���u�Ň�oLЛ0���Ν:v���5ٕ�ʊ"oZ�I�i��
r�7Iy�M�zVoǯ_�/��X�^����<��]뷒[��%N
h�J[b��JV�k!�e�����u���[C=���{ץ���}�ӷ�n�n؎��|Ý`�Έ�///Ku�����0�:l`C��+�)��Kq%��y���;:��+׷��9�w��Vיx)id�F�%�Ele�N��8�imi�mX�Y��G���v[�<��S=��L3-n�&�W���VH�N[�qe�уŖ��<��o6�{�s���xk�ҽ�{Ԭ��=�Q�n�,@/Ow�Nz�ޖ��
���^ⴶ�����w�}�K�yڈ�������cLRJqI�s�]��-����d	 6��^��l��8�/v��� �t6�zc�m�l�2M�^؜筝�n�4�[s� �r��>5���>4�ϏS�/����C��7�����3���e����W�6\Ie�ޙf6R��0��LbP��I�e՗S�;�Z���ԡ>���y�η�┥'O;�߽�S	B����
EÄ9h�E @�3���Ef�r����}��y1m��w�'���}�C�2C$�W���ɂ}懥7X]�8fm�h�,�$� �D?cY�}�5�3kh�v ��w!�x�OQ�e��x�3/x ���'��c��K���W �#�|/��"����Cq��u=$N{߮�v9)JPl�~=�}�m�$�wW����޷���>�~�(捆L�&ԡ4�dƏV�-5ı]���K�@����r�>|�,�&�1�f|�g�d����^ ܛ�2\`�w�z��OR�JP��{�}Л,��xپs���攣=��=�)JO}�\��"|�D '�S#�Ĺ(�35x"����}ӲS' 2�z<�����=��\���%�2�w�{�rd8ɒ�	��߭�GL� �R�׽�s1��`~�D}��|v�����f^lֺ�[�	�N��׾�eԦ9�������b	��GôP���"6�(u����Hy��N@d�x��7��n\�	r����7�&��1���s-�\��3=NI޸�I����I��7�=<�R����]����#%(O=�$xIG���y!��'�@g~��8fe���f�
���h�����%=�Jw��Oz�OL�h��M�S=�����p�Q�cf=6*�EB�Ma�{���a�;�ƍ��O��� �p�Z}>ȿ �*�O�@d���y���w�{��^�f�����}��L1<ߏz������h>���a;[�����V������ʐ	�0Ǭ�M
V"+n�!5�6Z�ʔK-RR�޾|�?�Y�8Q�S���N���}��%31Jǎz�v�L���D-�y>H�|>��:�{̘�׮�{�={߮�-�4.A�>������o� ��8vr�<I�|_5$�I�� #�s���v��t>���}�I����u!��>��޻��d&JQ�߾�!�x�c	��GY�y��q�����$q��>��(�b\�s]u�C�N�����JPd�~z�rn]���I������f�t|.���C�L�2f_;��]˲���G}�'ސ�<��L�3��9�>��@�𹮈𭚧iQ���}��1L�篜�v�r�#�=�1������5����4�9{�}���_.�(;�~�s[�p���3�[5�]k�Ϋ�C�25�<sl��  #�">�lG��|�VA�x�3�=�!�2{���n�L�S��3�C{�+L��^}��cJQ�}=\_PLH+ѻx���b�47gsDPM��체�e["�C��s�7��n�]��A��j�}�H�=�|���k���Aѡ/`PWD�x��H|�g?,�;x��}���ܨ�Qkr���a��l�تi��t�B\ˌd����[�+�+BV2��.V$�(eٲ׆TB��%t�6�T���]��QF��b��iQ�MA�\�g�\ ���R[3s��kEt˔"�Wdm�����H�Imsq[.�V� ғ��"����7'��u��ˮ�4�fS!�����xū��kV���D	u��"���bkl�ZB��4�T�9޾}=߇�[�Y]��Q���{9��{�b��l�"g5�׽�hv���{,*s�Ͻϕ���@G���������<&�S�(�pĳ�w!��E޸��}�){­�L��P��B����L���>G��V�K�L�;��s߽�4e���D�����~�Q��O��<��؍X����g(3���#���n'���2�	�&��}��rN�:#�H��mi�㸆�1�H��@���ǜ�Cn�JR� �=��cJQ�x��L��ve>��t�>*�M�H�V������ ">�"�]!'ޘZL!�3^��{��)K�����׻��%�*T]�Hϑ���Sk��	I]�
��|����h�)<��}���S3��G�~�w�m��ɲ����Č=~C�D �^ּ�p۩����\���� ��m��>�<��~U�efQ�lă=Z��j�:͢��Ke��Yp	�˶�b0r9��Y�G5#����{.���'k�|���g�X$ܥ.0d����}�	��"��"<���$xIDxtp�ꮂ���n\;�!!سW��({Ġ|<���l@�"O�D/o�q��IEâ[���,�� 5��� |�.��?w?��s�����;j�w7|7ï.5��y����-/�����̟�1�o����7�� �`n�[N7�QA=]o�g;3dzԴg3|��.��!�uI�;��zd�v�d�I��={��`�zH��>�m�������#�g�ue��	ػ��𢏃W\G��%0�R���=��l��ZR�^:���wY}ˬ�<���k��=$x}�O�����ƃd�2�~��}�m�ł~Eb6g	� �#�G��":�Rh�y�X�Y�#nK�D�G|,��2�����n��V�(�J�z��H�⏼	��	�Լ��ν�<��J��e�o�=ﱣryy��dgE�0�u�vxq��}o}Ӳ%(���[K�A�jz�2�{�|(�d�}���cC�2R�	��=�j ��|!ܺ��$I�hwom2�5o�~7��|�p46��� �5�Mv�j[SFhbd�v���;:��?e�����Y��:{l���{�6Y)��b�	߿^��G�>�'����K�I|>�g����v��n�� �� �����@�y�������	�Ւ�:L�ĳ�yJN�����r���9���;����Ɣ�7	�~����M�Be��Gr�^����/�P]�m�QTS��Ҕx-z�磕��et�����{8K���{��]� }�}�H6�j9/�hN����'�=xN'���]����:�RU�x8��Sy�͓{	�{�$�;/�#r�ض�t�m7�>{q:����}�K���׽�K�2rC##׼��O��<T��%���w!�S�@�����ibU6<��>�'����LA�	�1FHdc��\�n6A�>b G�ٽ0<H9<S��jv�/pt���~��&�rLּe��ɗV�k�:��ć�2=y�^��I�B}���O���D��l*��%5="d$��3�2�ə/��� 4�7���x��`ȠI	k)>��z�h��U�����@`.&�+2&���&0SB�R��ňLtBve�ʫvDd%{;�)$M�� 4���n��[kS�9m�i����H�O�$��k�H�p���l�)���UW����Uo��m*7�3nc�
��I+��^3>I$|�0�wS�I-k�r��m{X,J^����L�賉y�O�q&]����2�]�o2��ULv��wc@'�J�D�QA$[7�'�!�g�X�IEâȇh�����l�ב�V�$�nn��H�[;&%$�Q]��\Iؤ �5�(��G1�g�V�/>�1�ǵOxM�*��[��t��c�(�k~�E���S�p�i�>�T�u�N4de��xx�	 �&�L�|] ���Y��$ �] H��&2����lCm�$�;$M��̂H}ɉ@"PQ[�$Jj�k��VMO1�������b�-ܫb���n��BZ6���`��5���t� 1Ou�,'�!�;��<띉2�H$7be �I��! *�*�q�k��W�R&Q%��0L�S�b�\��79�2RHL�Q]�^�ʉ2|�y���0S]�&QA+�ۉ�k�EV��������vgawix�fD�)$L�l$��D�_Eds����,�32@���HH�L�t	�����L� 賉yH����ʧ����%�]�L�I)��2=��9;�z�-�hΖ	#y1)!^g�kHЋ���vGL��Ny�k���n�6)��A%��1) �
{�D�(�]���2�t_[hT���k��w4M?�̚�yRF`��
�ƅ�]�C��`���QMsB}1U��bpE�2�`��	�8�&Ԋ�E����
!��(3�w������RF�2*y�:�\��3	�a�Be���.
l�u�siL�(��aY��d
���T���l��MãW"���KF�&[D�@�\XD�\����*˘�pR�K���k����]F�6�-+Eo9��f-+
��aK����Kh�L-5�m�@������U8��J�ˬͦ�۪)�Y�J��뫚Hh�3��s�1�"f*�b��f�GMM,p�f�!]�B��1��~��AH�N���B޶dJ7�������`%{z�D�H��/2�ی��6��Ą�K�k6D�P瑲l"�;��3IWOD�)-a�6�滢�!$�H7�"g�$^[��$J$�vQ@�=��^�ؖ��9H9J"B���"R�/%�[$$��]s� ���Β�U<��+�N_H�(��^]��'җ{xPX�Y׋2ҷ-?=l�݃o� ����t��y=)�Yհ �I�vޖ�4G	j��H�W@�K����vu$pC�g�O�q&W�'�gD��0�b�?���u��QYR&BI#�[D��X�zR�Y>����}߿�y��o~�zN9�A�(����+v��%��
l<���s
&ڡ�cT!c�����O����h�|�%/$�Yu� �H�:�%�k���qP��L����)^VH����S�9����] �;u:f���L�o�F�D༊��{aB.c�o���F*m��l՗i�
��8.n��T�߼�F2%;�̒x��{�b�n丈�8��F:�y�C�<%e�H�o0Kvޖ��/t��u�|������Ѥ�D3�w!�d����e(�0d��d:I �;r:[�L:�����X�`$��d�&|���K�I�~%�`��A�Y�
��D���(�(����I&���hQg��$�AK����X�l��N��7�
zD�+,HU��ř�;	�W*�e�H�����k��PC?�i!U="g�$��[�CO�o7��Q]�'ҞRx�����Z-�]-�aKA�,"�ۜhQ�2&z�]�˖�`���st]�9�����H#��}~�_ߟ�&PH�� K�I%�"e)~��w�"^E��ɾ�>�RH7k��	.�G
X�B,����&���D�m��L�.�����	W��}H�� ��A2�-��s��zԦj�o�/L���@�b�x�4�6L�H$��n�	Q)*ի�ٵ�L5�h�8b���&���)����:@�@���GT�nI�[�6n�+ ���{ٻ�M�%ĐYS��FT��x
>##"�$ׯҤ$�D���)rxa6��g���\�7U�3=�S�ny"k��$2I���I2���|!�m�:����X�^s̩Ix[Ӎ���1*��D����L�ױM�*�rM4\�/�$﷡�T���S�i��I2��$H�fn�#�E�C��ӟX�y�04��B�b��@\�Cb���)	t:�;H�$�
�af�ggd�+��[��.I%[e �I���	N���d.r��$ϒI%=�"���q\���8y�	Gdęo36�ʪ�,��:_��6��BH$	/M�șI��}��(��ڙ�ߤ�>�q3N&ft�H��Z�,���h3�� JH�랉2JK'�սq$AM�H�(��ޞ�#!3�/G��+B�D����~B����	Fo@� �	+��)$���`z�,һ��EU,���멂6Ežc�wF��e���_?�f���.�V�s>�F���S�9t��;YG1�	���6^Z��=���|}��(�~ǁ2� qC9gr��m�D�H�X����e7�O3ٜ�O���<�&|�2c�)$ٽ}K~>{�<>�3������,��ea���F]X�Q�i�҃)5��k��,L��$���S�H��E�Kc�W� ϒ^K9�g�)"Pl�2�z�tm�j�#��d��W�Av<�@,�#�&r;��*�����BH(�ʼő��_� L��I�RL�����e$�O/OU�������P#�
ONx�w%�&qO>���s�Ik��HH�a�%򓾬��7`�x)f���	QIS�<�f
6���&I8`��*���dW��O��v��-I$����JK�k�<&B���8:��t��M�'�fI^�ڃ"j�pA$���O{_�$�	9��X�X]��K��T�fb[��$ϒI �o�O�ߚ=��<�� ���s:Y�-��T�1`������K�v��2�.(c�������2_�^� �>�>/�g�ݞ��˵���J����F+�;}���sv75�F�-yM��h9s��"l�����x&�>p�c�iS����w&����4�{z��ǷG��
��cX;��yv�>Bv[��Zx�wxkw)z!����J�t�z_�ˣi8I���Q {q�Ivb:GQ��K��{=���w��s<�(?�{u���*�����I��XO l�v�k�}snF������=x�>�{���v�v�-��Ձ�;�����}��M�S��ɉ�ܫ��o�j���K�;�ֻ�-�R�o�ꦛ�z���ǋ�������-V���e�(,�R�m��V{��ޏ���-S��ez*�(�L�yy�;=���OV��t���F�s��	���g>�oarA
���գ<@�"輏o�w��m���}���������#i�Mal����}�\L��@4�`��?��%� f%4+���^�#��n�yc������b՝����t��|�p��/�<�)��2��͐`7�Χ)�d]ѷ���$+R�����x�gvx?_˳�-���	;ہ�F���s��4������OO����n9���h��[�	L��X���ec��1�6������[��
�{<���}3��%�l�d����O�XV�ْ������:{��=�I��5��҂��LB\��_ws�qs��W�׋S�@�~_A����IɧF�.�����Ps.
&ff�r�2pt�毗�1	�4K��"F��-�BG�����z������~_b��-�^^^X�{�H�mĀ�:��NLN�7Bh6�X�γ�x�sm�$GG_9���v���1����xdFFE�4Ix�I�,֓6b�@���w����⬠9#��;�:t�۷{Z�I]A���!!;�y�����0��{�EfaM��-`fXU�ۏN��k��8��zҒ����':�n�B Kq����@J::Έ�:�4��ӧn��w��:�%�սk�O6�a���
��s����r<�)�d��֝-�2��<�	�y���<�K;2mۧIݶ����v\Q����"���vR�n=�fq|���{<Y��Y�q��jK��;8#,�,�.���Q㎊��u�e���/J��S��B,��hA8smK���W��&Ԗ��(��ޖ[J0`JՊ-�� �/^��N�Ŷ'6,W�����fBh��%'��B�K6��������nWE3i�Ăp]S7K�1\1l�˚͵��� ĕڬ�+Q�݉k��2閑�G��Z�;.v�)��YoۓN56΍����f�,
�N+�k��6��p6\B�V[�䕘L�5t�x�˦�L3*R� 
v�cI��o-Җ���9��u�t!
e�m����43�rLkV��:�X适9�%��3��uv��a�G#-`H�M�!a��k�Z�՚�,��@s6.�
���yz�R8f�f�ˠ�Ďy�Ppv�jU%����:��΢�:��κm)3� ��T�+#�[�2٪��	�5-�u� ��
�S �+��kH�[SV,5�ݒC�Ikm	�ʋK,ҹ�+�h�RU�ԳMv'`:��7bͶ1��lPLYr�6�3X�M0F�:E�,l�An��*j����`�Ε��6�5�K��02��Z`6�ɮV!F���m	ut�ظM�6�ZB�KN��Q��lrPNՆ�ic�s2�v�o�+���[Q%h,˫�����к��K��u
�k��@4����i��X�¦�ћJ�H��Ўu)c�Pɬ��h�����`].t�b�������� �VFQ�Vb�l���dTS�5sf�3c(@t[�����U�ʐ;�Qk��YeҺ�f��tV[��"AA��[���*Z!��1�T��0�s�0. G$2���RC]e� R�j�ʖkMm5��%�ґ��;Y����T� L,!iλ-z��R�0ƌ��%ƕָr��F�a\4��$W&R�LFu�n@Fm��fH!�]���ܰ��&-�$iq(��	3G:ʚl��,Vv���D���uD���Ԣ\�3�T�֐�5����莩��6SX�G�n&��&�-�iy6R�샥RZ1�6#(��n�:6)HFU
�ie���֌�ٮ�Jff�b�d��]e ���V�[y`�����,��+�@ֳ�wx�'�1��Q��Tcvr\��@�k6n%��H�9�f&s(9 ��k�����gX14!��1��B�E�c�p�tm�%��ib�m\�@#V�`��01�]����J�)Ic.n01��k��T�v��	��n�,*�5�l�����MV�ZHf+q����1�,B��RM3�PVP�l���y疵u6m֨	%����1�3�p�Ό�Du���CGKH틱� �����<�!����;~I������>s� >IO_H�	W	9q(uM�k{�>��K�v$�X�Ã �Ht\��
@WY�$J$���?[�R�Ͷ��IS�D�Iy#;}D��`U�W?P����3�on�8��o;t]�݀���%o���قU��'җ�A&�w����k]�+	����2��IO_H�IK�듞,���:w2�6S=*��8��3p$�K�j$�H�����$�H�4�R�Ɲ���	,��H�+���$�h�M�2&R�I.����&�Wκ�])l�J�5�|�2 �#$G�� W�;�<�Sh��'Z@>��;�H�X��I�=f�SsH�X^y����C2���A
��a�~~���m(Ǳ�����"f�`O�$Io4����Rg���`��_5(�x4$��`fR��b)��܇z��U�=-(%���LU�m�����K?��H7vh\�h[g,�ʞo�B���i���Ӛ�F8ud��~<=)�s/L^:�̫qޫ���=���t��� ��I)߶HI$��yA$������m���;�y��f$8N�v� +�� $Iv��I�^�;����Y}�5䗒�3VfБ(��]o<�Rΐq���w.��
�	��,ڑܺ3�%��Ɂ7�fI��<�R%c���mB�FO��$�t��� �7��;;�wuqit�\���
��7Bމu��ܞ���3�6�<�t���I*ǎS(��;oKHJn6b��� l����J,+��5Ű��H)ڠ��1�E�!n�c+��;;n^�7�3� �� �	�&D�%%�Ѳ;�L^I���Ғ�̻^|���gW�r$IH�
��T�*x�rN1����$-u]2$��T̶w@�H$�`���1$�(�v�$�i�ύ7�������O�'ҙ��JD0vw!�f�Ym;>iI�|̖B��IW�Ưm6�"���,��i.��C�|�S���	�O�6lj���a�$�j�;��Ɋ�'�q�T��Ἡ�L��C��L�$�L R��Ϟ�o�X+珔�E���不��{'�Bd�.�)�זWt�P	@��l�Y	$��^�iA$�:Ά�� �;� ���<���#o�<>O�F �~$�҈��fLq��m̺I�8s��mEQ:cͩ��%�ْҒ	%=�"��w���D(�\�%NY:N�Y�cc(F6٢ۈY�(#�E��W7[5�Ƴd8_�읝ܻ��#��[-D�$�����]$�S��&R��E����&�S(�%n�!�����x���';E�O ��%��)v���Ҽ�(S�t���fe��Ֆ.QIkN�;������܅BR��fX��%�4O��z0:I/%7�D�I]�Ő:9�����I?��a�%�$�@)��$��^.K"�܇{�+�����
�6P�I-��/$�S]�&RI%�Ʒd�
�Q�
y۷�K2�D�]f�c�$tU�1V蚸/��Sۃr�s������������}�̩i���Bf��n�����&Fe��319���[^���,C0%�1<�W]�3�K>����(�Izm����$^SY�$J+� ��$L�����z�$�t��Ej9��f��t���cp�dѨ����i�1W����3�re�LG'�vrP����%���yWnȩI"C�:D�J��2i2����->H^S]� �	��|]�wN�G	ֹ�Pw�z�=�m�E��� �&o��h2I ��H�RV�U��"�Zĕ5Lް�p���IZ�|%$Iu�D�($<�4bc���.���iI{�%5�"e��:D��W0�-�(�1�T�@��h�\��I%�uD�I.���J�m�f��.�SKJg����wLȃ,�V�%���w���\� �I%��bC���Vy��-��nW@�H��#�L���[��d*���zˁ2�lצMc.��r�o(�$�z/A�;'��W����^l�Q��`��C4����|���̙�N�趒��,F�ne�$�I!�I;�8��I��R�b%Ҧ��v0RX�`u�!-2jے��a�v�&i��h:5��\�`fڬ,iI��4ڲ��M\�49v`&\�;[02:����Eef,�˝���:����U)� �a�CCAf6�t78����b�Q� �F�i�M��&�`9��A#G��;b%�f�S�b�2ԛF�ee�c6�4`�kB��ܔ3Z@�~�����=��1��D�]e#��fZɵ2Bm��m���ϟ>�ci���?�@UfșI$��lKyKy��Kd6������1T���>]W2$J�&d����2�C6p�"��˻9(UPO|�2$��W�Gt��[3�3ҐH�dt���(6k��d$}U&���2Te�t��H	?�O�L��p�ꢒ�ˁ�-��^Iy#�g6��:h\��H�5�^�ɼ�FwD��>j�����)��vtL��Q���]�Nሆ�$�I�z$�H���N.vc�b����y#]�%)�a@K|J.�f|f��2&/�����T�檉C{fD�I%��ؒL��Q��&U�S�4QX�4���`b�
N�;0F�@����K��n�ڼ��39WQ���;V������8�D0vw!��>���z$%$ٜ�>H����27��4dL�F���
�rD�)$ٹR<�z��=$�Y���Я6_u� R	V��a��G�۩��A�U��y�%>���7p���|�-��E�׵=�{�i�{�/���<&?��S�wlE���h}4�=�����g��h3
L+2���@�O��__n>�[�3^�I��H�}�$	E%�u�Un$f�)��J�yC���w.�wadW<�) �n�	 JI$�������d���ǃ�$�fh��%.��o�33�	�LHJ:��B�ޭb���3]y/�LRA$%�dI$�]��;Փ���S�BK��1&RY���Kڝ�0`�U<@�J@$�뎉 �;�TT�n�Ĕv�I�%^fe�=�"	RK�:D�G8V����T��.C$�32k�kf6�9�jSW	�hml����R��A�6��=��[�Qg1�	�m��H%�D��ގ��������v�jܩx'�R	��&��������;�W�랁X��Y��g�0%
�����L�򮞑"P�OakC�_�D��é*��Ά�1D�$3ѯ(�Wu
�+�dnD��($E�����b&���jy�o��{��=A�ub+}�����Z,�źy4�y�6�9��hӴ$G�����E3S�V�0m���x� ��> ��<=� �Yr~H�f� �I/��2���11�p�W�q\�f��5�}R��,��(��F䉟$Kf��>��c"Ys��V�$��ʑG{p�=�����wU�e���@$���)n��jrIȲ`5�H�H��g$L�x��lމ$����2-gzܥL���h0uUpQ�-S#��RH:[U���Օ��hX�0,Y���x�S��J؈(�v�A�H$�f�I��뭷�[���"}(�Iv�ȟJO�e)�ȦNh
�'�Ǚ�f	g�g/'_ A'|UӒ�|� FoU�l%7�x(U=;v$�܈g횽�{d\�qbIJ��U��*W�^I�9�|�H�m�7va,[q.�+��u�%.��R$�J��&A�+֪80D�x��~�*��^̊�q�KT#�^Iy.����(���� I$c��i��N�sQ��r�%��Io��8d�1�'�>5Ş���$�,1_i�<�߻G*�*��:��G�מ�y�3\�^N����fff�d(U��P,�f ��>S(��H<�c1�8wE�Ҹ��e$��Q�l	���CU�)ݲ�M��2��I��$�I���� J��
��o�Ϟy�
!�����	�Yu��\�l#sE�ls
ݪ���J��Z�2*Os���_�m�8N룒�;r�J	7n�O�I �
6�Dϒ�1�44�]|�)���}��2��uN�%� ��&�n��2�h��co�h�nB�����3y�~�'�Q((��(�Ҩu��s���)M�J�m�,���%��P��2�S�`�sz�H$�Jh)�)�_j��V$�G�5�L�I��Α"R��#����wtꉖnꋛ��כ	ٲ�I2^�Α$�I.��N���Rr	/>vD��G�[hp�A�.	�%J�ޑRA.�|�"k��c�Z�c$k�L�"PQ��'҉ �~0|�8E�ftS�sYO��B�� ����,��/=b�er��'[��~�[�ϗ�����;�׿F������YYQ-�9F�d���F��V�e�KbeB�F�;3g,N�x����� @�&UI�Q)qգ`�iR�)nXA���]h+����TK�m��[,l�V]a.���ё�8з#���Xd���k��h�@]R�va��b�fDi�*��.�˄���k��X���-*��٢�-J��:MRG	fRm���9͕ݭ�[�R�,�6��Ԗ!�۴�78U+M��R�B�K��eJ��������u +�lY��Ch[�Ҍ�e��&8��,Kd&��C)Ե�sP&kA�[bW����qp}��C����9(_y��>	 �J76��$��y���d$�p�������J�ܑ"R��Y�����wS짹J�f�y�]�j�%�^U���t�tt��~dXs�Ҍ���s�n�'D4s�I-�:	��p�h�M�2$H	$����R�^	5L{1n"Lf�鐒I(��(�����2�[�q�fL�c3�����g7�D5d�rD��@�	H�B�c��D�;�M����[o��:�$�kdH���`n� ���z�e�c���|~x��Q���6<�$�c�L��)l_H�O��d��tI����OM���=E\��;K	vw+HVU��h�Ĵe��B=Ǭ4s�P!͆�����Ϲ���$;�95� ג>�WLlH2�%��!,;�۬)��~���H,��g:��C�����UW�^�����&[;l��)A5I�1\�Ա���*���ԺA�3CՕ���oU�����?\^c|��ѫݢM�x4_�*�ϡ�N6oƖ�*�I4{��� �(�
Щ0�*�$ 5M@��1-���Ft�&Q	��y2 ��M��%�r�"*��;Sbe/�	�,���&uQA.ʸ�)-� ���) �	4L�l�ª&zF�~I$|��l�$���&|�
�N�Ch%� ��*�t̊��%lF�I �Z�1#@T,�?k�&RJ{:C��c�Wg'͢��y2�!PѣQ�`���:I	 ��t	��y���1N�섖�t����Bݯd>��$nt�����u�y� y1u�n�p��ѻ8^WY�+�fٶ�3�5�;v�)mD����?~���*ٟ�>�O��N:��&{:>I�kf����뮁2��K��{-;�f-3l�E�.	�e]gH�JI	���;��=��Ixk�l��$3��&Q%�����e���)
�r��'�T��T��>H�́BD������D�U,v���Ԯ�v*f�&�A�@x�Uy=�ݬn���E����h��3�q.]��+Cݰ]�}���1_Gr*���������iX�L���,��o�仰��O ����Y�îq�h`���➓r��_��g,x����hE�ѻ���0�7�D�}��6%�}ޔ�~��N���s�&��P�3�8�σX�g>��J��f�:�?j��xX����G��A�n�����@8��[x��7��=�e�����yF�=�&�x��xo���=���L��m�u�8u��"{���o�xד�4�U2�٣��S�2���N���x�>��5_?`e�c.pt�]��fm�u`�y5_*��{�t���$8e�No����#���0��c<4���S];���~c������uOKoz�ר�u�}��oJ���1���g�g��!]-�cȱy�f�n�,3�w�������K����t������#��7�����꧜�b9��O=|A��w���L�?��{/����=�j-k��6(�[<�?-��$��<��G�o��5�=t�r K��z3yA���O�WBf3#3�84Z�X�{^Ɏו1nw� ��2��^�<	8lݲ7�9�fCu����7Q�x7zhۗť|RrI�r|9?�Ү�'}�Y���J`��c�<9�������G�Mɷe�Jj�US#��ny�ܞ����8��@;��xg��i!D�+4�$���j�x��\ d���=%#d=ý4�'){����2zu8ނ��VU��(� ÏE�����������@����,oF�y`� ���me������Х�$��=y�w�3הq���vڏl��gy����H6��`��R�J���n���\o�<��eoZ�aA�;<�[^�y����<���;Q���"Z���v���۷Aֳy�D�XB�"XF´� A�߭��R�Ju��֥�d�v�w��3���Rl-�hk������̽�ׇa{k&�Ѕ��e��QP�D�B�őI�TR���	-��5�:�6{�FM�[���<,�N^�'q�V��yh�[w�㷸�y[�3��{v�e�f�F��JI����Z�PZ[�e�S��"�ķ���mY�[o+�e�/{�{��J^bK+m�Ӕ� �
N,��Α�Ӣ�:s���k����cvYVU�B��?S�"��	2��D��
P"y߯��Y��s�}o1����@�BZ'��3��gS�e\6�M�-��Y$�]� �ב	/$�����$v;`3�d�Mvo�f[wKJ\�"ǂ,��&���!$����3��]�D	�o��Ɂ��2�^	/.݁�'��<&VM�Lբ�H�H��.��t�&���B������+)�Y�+�,���"�#��,Y�"���\�t�I+�q�I$=��"I�X{iܐ�F��p[�X�JI%����di���;��UA*~����f���u���"� ���k���HGl���L)���w*g�M��S\���gtIpHw�>�5oH�D��3`D��J+1s�x���X�|RIy�"^H�v��K��
9�1�'�E�GD�j]��;�i$��a$�HLVN���]-�?������h݋�6T��]�ն��k �� ����Q�X��W�o5����q�h�k�z�ER[�Lޝ�F}AC���!0"L#H�L�%�@�x���y���=�yL`3��gQ��\O��%�`�ξؗW�j�����mq�����I+����@s�����[-���=�'�e�B��6�S"�n�	� �C2�]b�Q.�f��R��6�,t"�`��M�8�	?����LH2��;oKHH\���Mn�]��3��"�It_H�+b.N9fA��&1>Z�e��Ica���`m⢩� ��f��2�Es��iI%�'����
v�! �M�2.]3��T�>�I��3 �[f%��D�M�,���oñ"PU�$J),u�!$z&�Ä�\"�O��@���в*���	 ���HI%}|�L�$�@M:��r�$�_\�������,|���U'�ji] '�\D)��a������+�) ��_�O�I g@�*���'���a���3*!��4DAt���{zN��Q6�����_x�l3�vO�R:��»�W��6xՄ�ǰOy�:|DkA���_|(ť\X�x�Ѐ�̭i���@�@�&QI��"U�{36]k��u�0[0���uv�!a[�C]j۫��Q�`�;� 2�kSe�uf�bK7��|��Q`�mlH.���Y�G)]n�0�kj�h���eE���B�B\!��4�Z
��[����*鶐��V��n�l�
��&6�4Ļ(�ˤ��nіZ-��h�Bm�e84uoV���!f��\̪5U5�ux%1fB��G�k)aU1l6.u���fM�:fɩc�\1�յ1jڣ�k�����?_?PRT�BE����Y�p �A@ ��6ĆI$[�!,��{;���gdH�IBߟ�HH�Z�c�p�iK�`D%䮋�]�[�# M�`�ߛaHI$��������|�l�v�U�: �N��\� Yس6��$I^s���H%��7sq�;��o�A��eJW��2���!'my�t��w����?s�A��,E��ld�	�[bY �%��"I$Gt���V��e�7��Y��
BH�U��	: �D3ʐ�z@	x$�]�"�
�$�firUu��&@I.쀽��C_�`�L�Hi���u�!�+�i����]B�*��u�,��ڴ��p���&�rKq���~��:�����pY1O2A%�5Ø$���t���Ff4R��TUTI��	$_@sѭE6 S9	v�'�jZL<;g� �C�3r�,�������YJ�۽$��DGY�#��)����ԧ� ���[���x�>��9|��)��}<�(x�͎vיּ�[����&��j}WÞu�Zh�|��c�]u�k��U�!2� 31,¤Ȍ@ D��(,�<��I"U��"H$���H�E$̺���Cc���$�f�x"�`�>K�`G���މ �Kd6�����s�I$W�"��K�zD�+�1�2%�&cEt��
���_a��5���>��/\����I���I�x.*��{�3���N AY]?nQԎ%'�ߝ��@~���U�	��.�n�!$�"�D $��tI���ԕs��,��,LP(�C_���n�Ъ1�6ZZ�^�Õ�).0a�A&��1&� �L�os�p��]3�1���<�	lfD�)"S��I'�7�3��jI�_�@\�!P[�'Җ�Ѝ�C�t�
#��R&6EƱ"A���! �K�6JI���d$�[�[�Ӕ���?�����9�L��b|���I��I�9�BK�.�0M;��J6�B��&V�5�B�uc�������@����r��J�Q?5�X͡B]��)������laV�ɥS�n�*~ ��>��&P	�B` �@H� �bJP9�vw�����{�(�I��L��v�w�ݑ`�"k�ꑽ,�&2̤T!x�^f`�f�im�<�����Qy�Bo����9{�[7��Iyk>sH��H;T�9�2%�&cV���g�$���z�h�ه�$����RC|���$ϒA%坐 B���^:���������?��i�.�J����ih��{^N,�f��4%�ѻ���|�|>�Һt��;�_%I��+�$�l�x��H+�0]� ��ۻ��i�jZ�j�i�RMW���V�\$�A��= �O8�BB�ͦ�j���F�l:ɺyI$�mΉ2A$!��u�x��S�k�2�����O/bR����d���*�w�z�$�9z�!$���ԍ���z���^I ��I }��g#tÖ�9)���;TW�=�|��'z c�:D�]�>I$�^��	 ��	l�?'����J������qw��nj!�_a��f?.;��:wY���	���K�^�1g<��^��˜��a{|�F{Q3�Gw˪<C�=���2 L �� P�� �*������a׻ߌǮ�wdX;P�Q�!$�F��H37��G���U�K3*$�I �����Ex$N�s̫n���9�O��?��ffL�ܳ8��
�\8�ܰ��g	k��f䥅�0�M����}ρ>Ox�"��f<S8��|��D�s��J	 �{�I����I3��I$�7���ozNZo0gN��z��F�z}��9�s�yNd�c��$J��@��IA�==o2�	A~�(;��pg����8w?�t|�*@U]�QK��HyA$�95���k{4� �I ����4�4#|�c3�b��Q��x�ά�"n45�^�;�����$�6���BD�w<ڦL�K�H�#З��ie�rY���;L�*��<���cs�	��nv�8�VU3c��.^I�;��I�z$ϒ��A�j�4�[��LD]��l���L����Pt��E���Hzh������s4+�v����N��A��n���ʬ��-�>���Z�߷@"P�AB�E�I;�R��{�Ii�BI�BdV�I���&M죳gZ���Q�k�\�%fl�E"�.�SD��x�Ya.��eڴ��GZ온��pm�M6�[W]��Ri�0�^�`�K���Ή�����ً-��k�-�����<h6���`�E�VS@��B�Cfjl�r��f��z��nWd�k�4`��MlĲ)�E�ɗd�f��v�� f�ff��i[0P�ǐP�mJ���R5/h���xq�U��50�U	a��v`�k�b����
�<TP���|����Q�g��\��Hy%�N�D��>b[ѱ�9�@2�L)
y��0�R����p0�b̋�I�̄ms�zY�U8q��:�����v��I (�h��I�y��I�,��{�67V̜�����b3�LU%I�g�($�|�x�?���/$f�:�����$�4�1�J+�&��)/j�p�
 �����׳';4��Fe�;v�J�fK�E$���e$Kq��ڳ�K(�m��l��k3�d��U+���I��ci�
lJ�&���	q͙�2�	/7^D�IK��ǡd�9����?>���#5�k��B�7M�U����V���w2�!.���J�ۯ߻��|�j�
b���̝eܼ��Mׯ�]�E�^@K��i�T��4�E ��*P	y��$1d�ƨ.w��n��p1��i����2V���/.���~�5$gJ�n�����݀G��g�"�͘o/BƘ���A�,�Bcc���dS����̚�B��=T��#� L�(�J3�%L���A
� �]�|������ν󯐥"R���E��E�z��sͷJ^�F�d��,Ȼ�,ƫɲ�fY �o3V����&ݼ|��-�ډ� n��D�Int��tV3�r��;�)��p�	�wKy%䳥�']�$��=���Ikt�dt����%���dE�IVk���H����r���HS�"R\�rC��F��6�/+�*�{�)/$�]}!K[��e4Ȗ���x�i���U�%�!!M\� K�qR����,��b�R�UU�HX� ��w��֩D		$�5�g��`��ꖙ3t�[f�o�!jH$���O��J�Y�%��Ƀ��K�eϞRP�XcN�4�%�)�I$��BI#���	�I�8�*=}ٚ�$�RA�y;�OLj��fI%�wT���>��1�qW(��yG�L1��x�������ga
�j�1�6�7a��ʻ�?	K��wT̵M'�*��	��o7�ם��� � ��P�T�A��i
Fd$>�� ���X�I��@�D�����Ґ��H�:�0N�cTj�麮o(��9��K���B@$J۴�>I$��?JjrL�9,�XAs���dZ�A.��w�*���-�/����b��%�.<�	U��(��5����ف���~���cЇ�K�6Y���[)�����ZӮv�V*��;m�>�}��y������y"u^SD�^fe�Ч�m�:۝�T^u���o�X��K�om�R�HV� ��w��*��E��n�ѡ���n� �*�6�e$�� j~�>Iy,��a�(;0-߰G���je�rY�̘:���Ud���I��Y ��O�-���`��%�fjn�h&R~��O�C����{�Ӳep��+���W��a�>J��>��%�>�D��H=k��e%���4�[O�6̵KJ`�<�)˲ac4f�Λ6ݩ�-L�U�������p���iVx�puL�͠j�����a||�����=����Ą���	0��,ȪD�� ��+j��g}{箶o0E�C�`��c2m7҉1�՟8�]�ś�q��IkT�I2����G�Q(-�����zro1`�2S;�N]ޒ�9��-��1 ͘a�90�X�-�@ꕵ~O�߷� �r��;��T����	Fsl#)$����Y��F�NIw��$'g�i�PIo҉�z����\�+��)΀�����ʄ��us��I(�}�} �Au�& H�˃����o%����B��r̓����u�e�I �f��l�$L��ѣ^��Mv�[i=�e�J�$|�G��D%>�/l��;��U��)��u��͑8���y"^�$1�!$��xK��-�m�܉ׅ/%���N*�JI���o������T��s$�-���X�.�G���~�}>�^��Y��`s<�O�p���xy��˸��t��ōyTŒ��C���٫@����d�s�ĝ�x��>�ק{��f����P�o��M¡��]LgD~����f�����wu�;��{u�����=��������>B{��>��7���t�^w���ݙ<�nUPZ-n�}֜��0�b��ijg$����A{�^z7���f8[T�h�.��
���������ۻ!�y�����gͮ�4g���I�\_�yy��N�&�>����}��?<㧼���燙,�N�a^��3v��#}g��]�����{�x	�7��.���xX���p�>wu��y�@�{�7��1��&�C����RW��[�"g<�նi~���Ӌ�՞�x��v��<�r������LK� bW9�=�{VL��G��A�a���� ���{�����V�7�\Q�>�<Z9!\�\έ�ꘘ�N�{/�N���q�R�
��n��>m�NJ����ޣ���=���z���s��$7��@�/�-`ќ,X��8��n!��pBb���5.�nz�qЌ�Z#�ã�׾�����A��u�x��}��x��C���q���7&�X٣Ҽ��pmRG=�v�2/.e|��۷X�X93���W=���;�=o(���
�(��V�۞���Ȏo�.R�k��M����9��;��oIv�;��m�E��=e�k<Q�G`�7��&û��o?s��k�?/oy��{ta�|=�8&��!�ЍF#�xI!㣎Lx(f�z)>�,����XЖoea�eˠU������.�[e�V�bSay�Ab�/�@�����/nŶ{v�;���M������o,�;ݷ�!UF3��O��{��9�UQ]uz�������^ׇRVM9VD�ޝ;v����0���D;��B��YP%����#JhoB<w�=�뾻��^�ٝAƒ֭��Y�6��ƍ�����O������z�\�^���5	�&�����,����/;Ӹ���u��g�u��{�u�[޴Q{^�g��zڈ��Gm�
�YŴ�!d*@�����f{�^� 0����d�o����w�ݺȲ�������;���7V,�K�J�9�7����Ez۳�iY�Ee��=i��h����S{��g�V^�5�w��������v�c��M��ܝ�X{M妿�5�+����Q1(�`��!��X��ƈi����je[VYa\Rr���nH\�c3��x�u͖+Y���6=��(�M�,�Kh����2j��ih��U�Z �k[0q-�YR*S=U��ud�8���Y�31F���<���&����,�6(�j3:�rB��Dgh:;�d��ܹ�%�lat]��1e�Ռ��)��0YR��jE�pZʔ���c0:�l��5b�ѻ����e�f�fkX���s��S&�)�6I���A�v��ص��T�Z���T��M�䵫0m{P�kf�/!iBZ�	2E2�qz�SSL�vڹ�1V+�V��ɵd��.�Dtay�rQ�y�pQl͉KL�Ō����,	jc���,�a`5��6rkW;a.��A��3H��%�s.6J�.�M�{E�&9���F$mԋH1�$`-��l�A�[Mu5�9ͤti���v]��+�݁��Ɣ�5��y��Nls@tt�&{FDՔ%�ŘT�0�f���u-^��-fv�1� 9�0�6�,+�c9���n4uXƸ�vŗ; �l�� Me5��uJKa+�i���Dr��H�&�2�5�fz�E�v��`�	.�����Q���o"�"���ڶye�j\X<�W�b�]d��"9aQ治�0��e��bG]1D]xe��p��,��0����T"	j�Mq�,�9"��Ǳ���N�ܶ���5���]�#L��]f�	aiPl��b�S�\4k,�Ǩڍ�5��4�Y��p�]�����v�3�b؀�ć\j��c1R�y-�E"3KUv�Z7Pv`6�j�j�"�ٶ�<f�trLVkj�Wm)F�����KЪV(�h���������r�3[�i2�V=���`����+�%�Lh�e�$�Q�[Z܏[�g�ape�{7������(�tlL�Lf˝�]&���l�MkIFihK30��[M�F�εe�@}�#!,�,�ȱ R� �J4*�珜��u�*c\���N�0(�͚�!�A�[�f�k3�6.c�8n#�у��il�[�Uщr��2�F�h�Z���Y�1Ԛ��\��5�]Xf�1���P	�퉋,Z�y�5sr.f����cb\AlЬLJ�a7F�t�:�[�\Q`�n&ڥ�dF�)��V�5�e
FkͰ�ڳfԪA�V�ӝE�Ɩ�3*46pj�-"���@kSY���+W?�	�߂Y���Y�~D�M�!�	[�#АI���kO &R�ŸJ�$B�v��슥)/$�^@s�� �r��;�PJu��4��?V�}��Ym�2�_8r@�"����QA&�P��]���|�o.�k.��:��zU��"(�qD��KZ�vN����]Q�I#�o6z'<�6��)����$�K w)�wTO5K��1X��D�k)�3*~q�I%4Ӫ$$J�v�J~ݾ�[�Mh��)ܐ]���� ���.Ig;1uP�a�j�ېҒIGclO�=1�zqRC� DQ�H,ǝR$��K���*Rg�����/���lsx�w@���������9-��2A]u�0�"�n�\�W%�9��??~	���NТyd�
��/$��cOO�O�)�9����կ1\��~���`9(�]��4�[��H�83�rŘ��M�>d�y��h��ʗ��B��~�N���b��ΒB
qa�r�9�����������i���j�w�Ӭ�n�:�x�f��������k^z� �f
Q&U"dJRIR`
T"Q$@�P(`��={ޏ��x$�K��8��)d����	�o�}���a/T���<Y�ܰgN�`Jq�� %ͱ!�($�mY�k�pD���d��	%<�= �J��*<����)�;�����R��+��y��+o30J��d2BD��}�>	/$��:D��]Ι�H'��R�#�tJVVyˤȳ����樐�"I��!L��q���q�e��O�A(�m�>�f	%�� B�$) ����w%�
�'g��hL�CSfc4%��7D��M��#���D����vNIg;1u�}���ۖ�PJ7b|��Ks�D$��4�|��y�z���-��Bc�)�%HIO�nYLF�� f�k�`@��gڗb� ��U(�h��**ߥJH����}��E�嶟F>>tԼ�V?\�Й��t��Ku7E{�	 ��ێ B@$N6�ؼ���M��ʴٜN,�B�?��NSFB���<��L˰�gN~N�yY'��qm����l����U��0����|}�(`Z
"I�	��@���*�(h(A����~	/F���D�ϜD$�罌Bd�X3�z�	���Ƶ��VZ�r�Ct��7sT"sʙ.ށI%仦�$�m�|2�4� ����Dώ԰��wA��<�
3`@�H${'3�N�>��
�N�$��=�$�;�@�>H��\�*�i�gA�R
�D�$��L�Ij�]�˓W�L$5Sam�U�n]��v�۪�~}�(�6�ˤ�3��sm0�y"{5�BA H��<HI��I�q�HM��R�	�p�3���w$��������e\�2R�N��n5���%$�n��I%�IF�ȔI��zVA<�ga�)1%ȏ�N�8�K��f�F�zbRD�=���=t4��\i�^I}��	$�7���K�X3���&�	��䋈�"5����s3 �)�q�Iy�:�	��z7�'<�q���퇄��gt�3mFY���M5&�ce<�`�v��9���#<��N
|̘�S�'v��˘��ENT;Zk˅m�>������	�2�(�	B
R(<	�Y�=g�y2w,�˼O���yy+�6$��	ܹ}�O4�A�Ec� ���- ��3m�Sֳ���$��⌳MQ�=o2�K,�Lh\Sus)q[Q�.�U��sjgE;��y�{�;��̏A7odI�6n���'G01}�#�<_;\E�v�6ɴ1��g5C'��A�='gx�ّ޿S?�'��ļI�wvH��&1뻠L�&[q맶�{/S�rK;�ً��lNA� �_lI>'ǚ�)Zs�E��b{�6�$�������0ͤ���@%D(��TiV�Xב���	�!��&I#��u[k�52����#j��ī$Q��'t;�2����Q �Έ�u�@��&
e�,��8�H$5_dω���c37O�<�p��ECD�7��=�Apg]p�����&���Yiu����ls�kt�˖�ua�-UI�R����ڜ�ap�|�>f��|dY�hJ&D��f N���#�UeL�����K3o͂�\��mA]�&�S9��l��лl,E�Z��m�qWM	jU���[)��4,���g��<�Sdes���ƹJ�4�#FcV[�b6�%��Q˭���T�E��Ԇ͠�6�M����ة�Ilү����WqJ�MQ���d��	����)
0�&�)VJ���6�%���@cBb�A���f�3K�����A����S����-��b��-��?S��ۏۄڮ&߮Ǯ�A'ůsbI �tD�f�*{{h����ޙ$-�`���wA��<�1�0 ��~�}}�+���	 ��뾙$�{z"�D�BYi�ͫhy=tE$��L3��u��$_��b ��S�5�̽H+�x$�gDC�3ӗrK3��ΔѭQN(���Oo��E�}�kh�� �|O��"����pdq���8w*[�q{I4!ރ ��'f2 �I{[��T��Wc}���R'�/��� �����>�n�"y
bȉ��-�Q�4Pf���E���ʆ�]3�e�	�8����b�3��$YŁ't;��U\�ʻ^ �A/ͼ�z��K*壢I �z��jWyg���vt�Uҷ���vV��U �&ݭ�C������c9�\H\x��X-w�p�9�-�3y�(i�a�F �ר������G#%�	pŅ��4�NcW�;ԧ`ep�	ǽ��P�&D&P�&F��::��'�f�p}�	~��ǉ:�b���xb:���r]���&���x$�m��y*�_&-Q��;V� �o���k�#�$��`b�3'HM�OC&Y`��}͒ ��C��$�{ޝj�˾[U�=u���C��S9��ě�j��;`<���W�/�b����l0 ���铲љ׺%�}�w��ߩIIh�S��R騃���5�ծ"-��C�b*ma�m�K�;<T���υ����<�N�"x�NǠ�_)��9�>5\�r����^8� �_���!��Mr�N�;�T#��dv+
a��算�@�%�]����;�|I�R���r��A��"s��C2w.΃��QMp��s'�$�����su���`�{��\�m��TF�ޜm�>���ը�/��߷&_*h��� ��CE`�G�c�S��̷vk"�!��Ѫu���� ����aB���
�ַ��!��LL�}2H^���.��z���v�6�O.$��[T ��H;Q{I��q��g�D��o$G���L����d�22��C�ߏ-���0���,:)��-��ZLx���>����}���Ͽ>�@?C�5���;XMaٍ1T��\˒�Y���MW-�����f��ϗ縭�9tz=��Z��fĂ	;���T�ճ���-��~0H$��!�*���RN�鍍�LA�ɾ��36�cD	"�;&I�$�G;"�굋����F���C{vz��F��M�Q.�\;��z/�C�"Fn���iߘfGZ}���`���I����n��d�ܻ��F[[�մ1�-��sC���$�|N^dA>'ݒ�U�q��xc���Uf��߉��[D��e\���/r}W���<P^*�f߆>��챛���R�Mu��6.��\�����u�e�� "dY� �	VdJF�")R�׮{�7�ۘ�D�wA��<�1�K��?d6B���5O䛮&d	5ۙ��|@#�_�7`��`��<C�I�wHNɘN�sKl�4
��ܚ�3�72����t.%S���>#��J�Rvowz�v�_����ĉ�~0fڵ�5;y���-�2��GH^���́vZ�r�Ħr�ɿU z1��SHR���=�(H�̈�%�}�/ƈ}�G7;ь6Z'+d�!yP���
IݠsF�>H�Kt �$ʹ�v����~g�����@�|H���i�H9d�9p�O�z:ruFS���@"�r�`�+��cuR2��m� �Ƽ/0{�pfL]˻��Tz��� �m�H=wq0��t\��&x� ��{"	��_L���Z&���UKw���g�7]�L�uD%DT�-r�;�=�+2l�c��[�[��d'8�kb%�z�C��ӑ�&����B��(|d�`I�e�w�����ᯈ���vf��F�l٨í3*n0�W)�mWdVe���\�M(�kL;V,�0l�aa�ͺU,ʣ\B���-�b]�hlB5����:�il��6Фz��͗���Q��36��4:Ř��i��W�q�X��)���r�[� ���&���Yy�5��hstz����	�nJֲŰ��fS6��Q+��)ph�53�4�ʰ
-#���[��ߓK���i{??�<�����a�o �"s��A5�A��p�����x���aJM��@�I�k+:�H�=��l�'2r�H��� �wL�@5/J�r�E[�c�Ҩr�Ħr�ɍ-���M]stO� �|���t�dO\`��C�cL�H��ޗ��0�zL�h�$��9�l��g�Ռ�$�CL#�|vw�$�A�ܽ��e���h�Z�A�h�r�vr��(/��>�Iv�F�9�������	�V���&3�b|I>=�p#��%�� ��Y1����c�.�s�5#�[e`�-Ҕ���Д�N����d�ܻ����CkzvvĒ>��8�Y��:�kǖi4H$F�d�$F�
��;�p��2v�A-��o�K���޺4S�5<㖽f.iG`�7�x�BĨ�Y��'���u� }���{`�z�=�7/�߳|�ߞ��7��x�#�`jd��P�F�׾�|rh(;��׽�)��ͷ��W6iC?U_�
�1���N�{[1��{v�kB�ˋ�c[y��%�o�A ��b ��!ӂ�9gw&d��HGOZ��M�H7�u�"�m�;a��Wc؂h&�����$HB��3��3���D���@��G�:#ɶӘ��6�����	��2���'۰�`������L�M�rC��p�`�Wj�c�b`݂�wY��tn2��C13�����i&�wt���Qu� �H5�p ���>Z���hZ����2n�cҁ�1�����gr��3̓8���'b���SF6/�ݷ �O�ls@���U�]�d������2(0V��Å�y���	vF@�'<�@k�V���F���u׫:���o���x5��a�@��d�Uy���>C��WᱰS�3c_���q�.��	�9�����{t�����f�z/���5w�{��=Vy��3Ö�0�pf��q^�e���<@s8t�
�&����z���������n�3E9=�o��z���x�fߐ�g�oa�}�y�Dv�b�7��ZU�>�R�ڨ�#}�ō(�ؽ;g�]���@x��mvob�lvƬY��P��z���3l��G�}�*��|����'�]�v�>���:q��n��S����-Y��{��|�pO@\�*�;��@�~���)��,F9���vbU�r���x��ɷ��kz���<Kٺ$�{�D������>�xo_K���+�菳}�� ��z1��xo��G������y�R�U�xʤ��`��}��7y�v��V Z�z�sӽ��D���g��+�E�.64��\~H{���Gp^#W;�y`��2�E������9P�'�����z��x]+�i�m���1��^��9���"���ٔ%�}��������	�q���޽]��7A�^���2Ӧ�b/��V�M4xcᅁ�m���ښ��WOh�
�m�z���G�pկ�=��3{�'ԯr����E�}�>�?O}.�MŁ��
�緼�z?���~�Nw��yv�^/6��r���pɓs}��Q.�]�o��="��	e����roe�Ys���D��5��f����s�w�4�l��@Km��}�9�Of�f��Yͭ��<�?���38���k����ۮʦ(��e5�mԷb'ׯ^-��i$�D&�n+4������Ye��Nݽ����a���6���vfu�VC��m^��&�-m�Z�q�n�ݺ7��022"�+����؊γ��JB�g3HaQ�a�e��XbL�ӷn��ۈ��:3C�Ͽi�ZGY�6緁O7hm����jf�8��f2��2K$���5�ɻv�{޶n%.�Ķ�I
r�-pI=�nۧ�cy�Y��f1,��K36����Q�;iM6i���,5���f۝�3�s[vͅ�[�,�4���+;mf�6Փi؍փa��H]��rvaNf]��n�[QX����n[m�,k-c�l�gY�m���ZZg-i,�:sL�Y��:�l~Gw��I��e&"T3}���U�ۈ�{c�8h�L�c��'i���{YB|�����. ���x$�w�g����KVa]1�R�!ӂ�9gw%��N 쾉y������A�-��B��J��vy� ���wZ�2��5��k�5���"L����(JJ���u�%r[2wf+��:9I;�HǞ� �{ A>Wtɏf��TsM�툈����x����wgL�KzW4�X$]��,�/���f���o��	3Q����kzd�w���>��i�̂��m�2�]�z�s�߉�{��H7�h4�i��~je�@���	}��W���l��8^gUx�mmBNo[�x��� �ۘ|	%��fI� �ǳ�Qɒ���|`
	�w��ջ�������M���	ܶ˹dLs"��"��2�|�o-[[0��-���}�{����L���*���5�ۘ��1�p��UW}S �>ݨ�Ӄ����NF��$��x�Hי2 �m@��O�g��_ao�ǖʲ��dUEe��ip��kŕ˖�6g]R��l���$m�~��N
`�ܝ�1�`A'���bH ����ͽ�Wl�lc��0�O���j̙'|�:-3��3�������pi���n$�哰A>%�o&|O��;�P"<P'\�paq�(M����z�5��	��wgfw�lWL��ځ ��v�i�S��I1o�2	$�9��dçr�A�˨�s,t��@�r ��'��& �^ ��cE�)�H&����(�M�`���Å�{������x�ηv0�D\��z�f#���w�׮���P%�݁�ȳfs�K�����D~���;�s��HT>�A:�NN;��c�T7]�b�u%���֪-)%��� u�Z7�u��efh��|G�L��L���O��fg62�aI�iv���1f2�e���h�.W%/%@�F[�1�4�2��+�й��](ZJԸ�M�Y��L ��n
�P�dжѦ��C�)�6�Z�a^%`"b�*����ѕ��l�N]vX����q-`�u�B�.I80sv�Yvل�c�(�#	Fh˹��#Ś$T����v<�%������B�(�T-�
�&V�e5Kn���Fil,#S4K6XB��`K��w����p���O���ӑ̽�+6��s����$���w-����݉�Ů�e�+N[p�M{�!���'ښ9���k����٨����u��t0���H;��gc��$��������$�k�b�4r�H9"p�읙Ɂ\�5
�fD[FuGso��:���C1��OF�N�>��z�qU� �ՙ#�h��3�N�;�x�(� q{� �t�cj3ĐsA>��H�h��ޙ)����fv[�/=��Ő]��!�d��BPa�H���y���[e7`V�놠�(�z�F�b�K
��Y�;�p�Ͻ���b���	��"۔}�g�V�M�@ ��P	�{`�	�#��'i���S� ��7z���,��yC��xz��k*\���#.-&�Ƥ�M�[��^�y�L&���(b+^t�ݨ���2��,\K�����ѓ�Z�Z;�Y}B|afdI�[ߝ��$֨�$��_}2H3}"�f��{Q�;8��t�30NY��ήp ����^5�X�+I.��s�A$�4j��oHB�����:,�ч�2f�8%��	`C��I%�GD ������I�vW:�@z6�dؑ�\�Z�Eۄ�h8vt�����2|&�i�n��Tµ�K��X�x;:D��� FI`l͗���^��b����h���4�$��t�-�o1�˚��q����χ��?��f
��>�;��7�'�7��w�n������6�_6�D������3����`�t���
-�����,�o=�dI�{j#�Pg]M��[zа�A��"	pS�\�L$ݨ�	7�����L��D��=X�7Y�|��L4������`~�
+�7��c���$o��M�$[�F[J��;�h�
��=�>>�$�)�u��{j�=����(���>x��vvL����3 ׺���Q�"�߉髉Gn�@ �֎�7Gu)V��s	+2�d���d�@`賻E�	 ި���z="�*c<w�ʹ�	�h��vM[�h��� �tU�&�Ƭi1Ǝf�.�fau�[�6�me��6V�w�Ђ����ω��Q�NsG!�&�_��{�܈ٌ$�ި�<��z���8.�C�Qچ���[����ĒI=�Q$x��OL��|s[%�2;�i鶞 �����6��ww%yޫ��l��O����@�k+��CTc���'ă[�':���ؕ�c����u�Rw"�:Y�a陁>��� 灟��O����A��zW5�ܔl���ؕ�ᚱq�؂�s��͝�-��L!'�_ǘ�T9�x�T�V�{�ε�~;߯=�g��M4�U�>�A��(b�30k.쌅��Z$�����K^V�����%�|��#��`	�u�L�W��[-Ӥ�0�!&`��(��R�6g\3U���p�0WF�e�iX�4֓m/��Zy��/0t]ݣ����$��n���DFWtύ�;�d�7~=sq���>3���0ܧF�T�5�>$��֙�z��Pڇ��ޙ#�ww	�_3m��[�C8.��4
R�h��n��@-��[�$�/���-�[�@���û������{iDᵽ<���z��xj1�O�n�ĂI�n�M�h��~0k�R�Ȝ�);L��ڙ�$�͸"�#;!�_�oؼHh��>���w�'�X$B�r��~QZ�q�iC��܍���[������(x=��@��|����~>��+ʞ� �=<�{����zb��=ɻ��U�{}�"b�3I�33��#�	��	ir�+���MIA�6h�'k��5�톖���A��h(�b4)	�!���۬�HQ��6�kK&�sM�,��9�V�Rl�Wm�5��Il��a).m13��F[b���G@ �5���)�rd� @������� �hT*UWr��Ў�%]�۫��6&1ڄ�9�V��fz�6 �%#.b)���i���X(��$i�m� Z8T���Yb�b��fl� ar`٪ϟ>C����Fr�����ZLx��͉$�7-w��.�ː�[v��Є�b�D��U2�k���E��h���as��k�,�����$�݉���,�l~a�J#O�F�9%Çw)љ	�vg�����wS�l����tp�H���N��Ǚ�z��!�p��F˷5=hUY�{.(G�$�W�I>���V�qD��2n؟E�d�$<ucl���^w�7e�x�Cd�����~��y�$I�ڟO��Nt��,ئ�5�c��*B4�u��=��j����	�6�f+j⤌;W�֡@�^�_r�`t� ����{�R$W�sn= �v���/���9�(M
����KzP&�b=��')˺f`�]��ݍ&�Q�l�P�ci���DNO3���3���f<)�m����n1��LT�K�f{��~ķ�?z]�+��<�~�l¥���A���*L<Դ�����Zbbs�x��ʪ}�����λ���6�0��~�鶍�H�0��4�Dy����a�=���!�"c�s�v���%D�giި�s�.h� uܗw)ђ���l!q�
i��$ʹ�3�oz":�J����Ag3�c��p]×i�t�t$��݁;�ZuPoE<��@�緀DuoD��>�2������Q�G0�:Sh�;��)H�7J��%6��k���G��߳c�f\����y�ܼ���u]�ޠ�^�\4l"�tG�����#}�+�0���'i�ۘ��g�L2��Ҟ{ ��ȂH'�ս2 ����!쭷��&ڃ�f`���Cm�@�{�$jEfr���v�SO�ͷ���|�U��_(#����w���k�[�ѵ�X�ӷۏ�]�:�NC+5�j��d�y�I��D�7o����� �WtH%a͓,�ǘB.��'��m���[5��ܮ�A��މ���;[za�)�����1o��"`{E�����݅=2 �F�f7N���ٙ֬�$��k�	��$tl���b!�&V����+�4�f� ��f).�60�eZ6�KqZS�\�r*��,���r�|� ���8��ѱ���F�3T�v��<I1ٙ2#����3�gg��TTl�=6�ejG�z[�WC�>&2�fA�$l;oT;x���ll�qۣi��"�^ڥ�c��Iګ*��A&|{'fo%��]�e�s�!����3�~HoLG���n�a�30w�Q�*Zy��+���F�I;�90 ���#CR0���v������0�a�%�3"1q��i���d����\�[N��O R����Հ�U8ǒs��c�}D�������xo�L��W��{�a�� ����Q��� �r>��,7�_�����lΟI��͎x)��~��,;JfA$ҝ��(��JK���4�me�g��qr:,l�4�12MR,,�]ܦ��gfA$�Y�|H�����Ρ�^�g0�g@�	;�1� 0xc%`�b]×ie��Ń[��(����H��$���9���r��ٓw���FN� G�2�1�p��ෝ�c:b	 = 9$�1����"��I'�%��	ų�$o�I�>!avo$�����jq�^�n*7;��kt7�'�G4G���a�F�hx��7�0
���ni���3p��̖;r�k�)쎉0����x�N�">$R趀H1�}0J�)ۇ�&%ߤ%�?)/u"]��� D0k)cM)ϕy-�g
����Ӟ�'�*���Λ�w#{��3 ���J�Ӽ�;����]�vG8p�}U��1��=�y�叽��{�U�x&�B��a�3�*�i������9/=@P8���	�VQ��|.�ǻ��&u�����������wOǸ�����s�}>{J��o>0�|�,b�gl�Bl�i5t�eճBp3_���O۞�-����sZ�^Me����y����w7ot�HHAb@����rT7ٷQ��=#:�ڳ��m��y��6s]��L-l`�n�=��2B����=��.)p.�ش�S�װ�;j[�ͬ|�)e���<_h��<��Q���n�����m=AZ�x%�<��6���~���qE������@��Wؙk�ݪ�l���-�I�x�{�_y��:���^ݫC��EÞz���dBn���OgQ���<����^�:��@�L;}%]r�ػ�j��<p<Y���k�*��-�'�/.Jv2' �UC����0V��cp\R��=�d��c<W�N�|��ч�����ڐ�ko����މvl'�ˈ,��;;�9y�fN5�{b������| �<6摓�PI4iʵ��_i���{	C76��I�O[�ֵ����cɋ�Z/�[ì��{bw�ѺOS623���+�Ý�mY���;=��-��1��N�9�2W|�^m$��&�
� 
\�p�;��gH�Y�@]����q󿂽n��Ja���	a%��cʧkea Pr!e҉��U��R��îj��ö�����'�Xq�"���S�������iy�0�e��l�Ή��'Ɔg>�.��q��l�m���[[Y�q�l���5�e����u�^]���۷oc�fM��QAe�d�dldtS6��CJ>��t��ێ3#I/,;����;zt���tU�I���e$��ibڄfŹ�N�,�q�6�S��v�w�}��|��ֵ�Z۳�jYpΰQ�vA��f	ɶ��ko�ּe��%��ѭ�I�e�,�9��#>�h��ܗ3�l�m7ie�Rq��n�ىfM�[5���h��Ά�8r�d��8��5�dvv��'rm�FZf1,%�u�cl��'��l���͆`�[k!�w���,�1�ݵ�#�!k6Nku�e��Y������L�kCm0FN�ge;9�r[�Yݷ�d�g�rH�ȶYm��[Z��b�D �Y׃��)�	��k��F�	Y�Ԁ
�h\��3��L�'��y/[<�G1Q�,��0.�%ln1�8�Y��5��X�7 �F�mE���[��E�:5��[����WX���-�̠Ye1��n	f͆.9XlZl�˛6 u�V�ũ��5����t��:T����6�u��F�Kj�,5��c���<�m���j��J#�݇�+/����d.6�!�P��Lf�eQ�9e����at��R�����*�F-��&5��@A�h	�qq{E��K�--��W�(���XsA�m&#R������U͈�W%hB�Ԥ*ݳ��k�Y��-6��g��m���)H	D0n�&K���M��4�f��EU��^/��-�C`�G�����1p��F���4��]ɊF�Qa���lM�]@X��h�)K��eu�%��3%�J��i��H�nuIr�Eva�3k4�ͮ���[ Zj���XY�$�	��eIj���,���ݳ��h��ٙ\�n0kɪ��@t:�f+�R7���Y�u���
VWm��`Wv6Ό[���7\b�U�̳F��1�4�UΖ�$�l�m*P�Kf��
�#�K��$��L6'1��X��[�.N�� 5�f�2�Qu8!qB676ݫ��W���ql����ֱ[W�S�X��#�e����&��àX�-Sc�D�@�9��e��m��v�2�Ck2,
蝳��d
�]`�s����R1�Q�GJ���l�0�lɋv]�����B�U̱�o<4_3�g�6Q�Z��s�6�1`�	��J�4i�uŁ�"3��8h�u6��X9��Qp�Q��AQ����9冖j�ݣ �̓e-��i4&ζ:�j���ISQq�$��H�;8%5%7WK��J. :<��X�V��Y�n�v��������o.|_dn�]���GT���Ǌ7ܜh�.cu6Ƭ�1�l#��^��ݢX�cZ��n
�L��넀�����l��s� ƕ���KMCl���"W6���u/.,����f���t]pӜB�P���:9�]�4���2��³��j��PI��2�N��-������Ie��;�WB46���aL̀��^���mˋ-���؆�V�1�n������ښ�˜LdYpK��ImId�6�iZ��G[`�nxt�Ρ�����>uCvN�>�: ��Xrz� Fvt�3WA�y?\ǠM.�h9A�C+E��`�@n��IתR��޷V�$�7�o_D���v�׏]]�A�x6#��b]���.�:nz<�"��$/$ISE@�w���'��Թ��'�zw��|Hg���رw	��2c�x�pI�]��#��7xb���Ovϰ���9x$�
3�<Lz�ڤ	8���;T�=�	vl�����_� ���f�L��^D���L��L�9c�:b�$1�S��v�����m�2��J�l3ê�sj<f�X�2,Z�&�왘;�vG��͘ry%��s�w���{�;����j��)��>���u���`���D���Ќ6��X]��-sZ��V(ڷ����w�s�p�^����c��#J�3[J�62dQt����,�ު�e�5��y���*��w���?>$��� �mG�ѯ�����k����H�
Z.�X2�n��&�=�	&��3Ag,�;�=�x�c.�d�H�n=<�y�Ļ�ݪ�F�v[^눫��1!���y��9��t�bjƖ�&#�d�!�{�͉�.�7��c�c�I"�2"D�U{��b�� Ke_H�O�f\���Uϭf����-�6x,s���0��m���]�d%L�&)� J�٘���Ҵ-�y�vۺَ�㹷>� �sz��t�4^�I*����Ќ�3�o����N�ZwwĴ�0踂z�l��n���S�Y����I���>'�;�����Zd��=sNI"�Nz�Lz�9vQ>=Q� ��ΐ A$���nJRn�	����-F�D�J�$����S�O�y�kG�D�n���v1�m�]S6��%�܉tK��p�{��I/1�A��xh`H�wr��Hg��07b���:ڤ�������|O�'���	9�.�'4���c���[�y��:�w�P�=���ē�:�Y�LN5�����>I.�h$�D�t�,��-�_,'�V��T���ֵ]BᴌJr�!7l,�*�ɉR�J��q�&�|���f.�wp��}���"�e0􈭾�6=�����3��q���� 'U���63�o:N�"���O��؋�L�շ�P$R����D�uQ�s�r6.�b��q�k����t�@��L@ro�M�tH'���Fk��׾�V��i�	�$)nSA �[� �e��Qg�!�C�e����L���p�l��$��Fft�$�e�p����5x�'��d��0����o��	���F�M3�8e�cι�U;VE���"sA�F�1Sh;+,�2�B��n�4��!�{�	G[A��V�VӤ�'��;2O��ۊ���.��U�ށ{� �Ov\D�QJ��1��F4�bP.Yܰwr��iH�㔌h�u,�؋���4b����z����5R��Y�ga�����A ��. �uOR���gN0�c.�d�Dm[�`�w�w�1�/9���wFu��6�u���� �	 ��rak�o1=W���:$���]��;o���*g�ٵ @&Z��5�U�87���]�Ē	{)�ٺU��N��X;:U����~��پq�?�-�Ȓ@$��㜣�
%��b(�uݵ2H�ސ}l�DC�r좼z�#�A �(��<�����1Wd�\t���ޘ�g�f��9���oO/�j�5S�������*nB����s|���w�ٝ�� ���Gw��~�P3f�\�)Yx"�T��i���nE^��xC�!}���]K�l��6�$�Y�źM�7(�2���',.�kc���X!�5�ڐ�$X�+,Jd�DJ�e�F�i R]�[[ˣKu��%��%([��)�6�]6��2�Ybi��v�Zu"�B �a0�b�Z�7I^����Z@f\h�iKX�Rd �jL�Hʘn��;M@�	+R-μ0���&��=�mҕ�nШ�]�f;V��ݵ�b$ԥ�ԣ�Du�֕c�p�]nk3��fm�%�(�)��{�F#����:L���#��k:`A�y H�i�������w��	;�13�V������d�(�`��[W;�u�"|MwT@�>'5���n��]�H��ײZv�ܳ���t�;D�Θ|O�� �+g,�H�j����0	5�. ��q�F��qܳ���ًhԦ��榚K+�OwT��:�4��yd��e�4���4�%�b=�#=w�cPt��僱uT_q� �sٰ?Ei�mEW�u���'2Zx�O�v�D����}�����w�)����0��h�al�d�ncsIr�m*�AaLʱ�v������;�����<r죎�lA��Cl"	 �;j�[ұ�ʫˬ��~�T?(�\a)XwN�&�N��O�n9�e�;���8"9�&X�w�BUd�B9L*�-SVUȰ��!ח�Yv�]�ט���eh�Z)���Sq/m+�Ƈ���y\,.��{�}�߄Ft�� $x�o�L�A�x�/#���������s|�.r�`��Y�t�q�A���>=�^9={��\��!͗��#����O��WgL�g��r�
N��b����Mu0���g���<�2����>/��'��N�t��ת��ec�# ���S��o6�A�f��E]���k���]0�==�"@$��uY��}%�g�$��3'v)��"�,\:Cg����JлhR���1���z��3]�gϯA������غ�!��H=9�}���:��*�EUs�$.krv�%q9vQ��.=��޶��X�h�A &{vg�����)ۦr9ܠn&!�׷"��t�MtL�� �k6`A�2q`,Gks���c����zoaY��i�z@e�]w�eD^����6FB��U̻1��O��*
e��n7���w���w�����H;�/g=������c҆���n�t�	1�=I ����H'�߹��!�����"Y�qܳ���t�L����I[�@��3u^8�*o	Q]2H$�丂|m��<S����1ɗL��Qo"	��i��b�B[5���6RP\�sۑf���ƥNn�x�mft�yˮ�ڙ$��z�m��	n��wn�?w���d�A��x|�v.��ȻS$=t�ۃ�!�7wYUu�	'y�#�>W~x��aj�� �p�a�d;5;��W��GL<��OT\A�$�~� {�N�ɰ��Li�WN��n�\A>6��$m\�%��t]3L�L��^��b1���f��G�L�/�FF[�$�Μ��3�%�<��u���j�Ż���=#����Y�N�"(Zf�jޫh�
WwB�w��NyEr���?���7�6��jj���瞫w�@#Z�]��'f��, }���*q�=~ݺt���nOx{� ��G����Ac�Kvp�>֞��n{v'���·���� ��<|O�v�d�����>���A����ո���Wڶ�-�jkp23qy���ģ5v[�@��gf;�p�t.��;�H��>'������(�k���j1�@�]Dx����	�9����o9e3�ڑ%3GSn����f'��� �H�'��A �NܤC�gm=f�b�$�F�k'vgd\3�����	�3b@'|�l�okb��7�Z�G I��x����#��҉Z�� �(�j��Ր��xN�:���f�		�ܙ$A�鬌MI�Ё=/ �P�\�%��t]3L�L��>"��!�VQ�ڶ\lV�� ��q$L�d�$ot�0��/\%�&z�<X7v�YNɳt4V�4w�����~�pQj���K�/w����G�h��\Rw��X��,b3�a@�:4�F����'U����Ju�F�A���\�����X���B�a�D�&�)nص�l)������t�WZ�U��:�	�EL���I�t�;X��51+L]��)�fY�l�*�fb��o�v�@�9W8�vk��$%.�f9,�3`0	+cR
�&�R�e��C!�Z��Ś���a,Ű��s�[@+]��.ͮ�kr������Z���[\�녹ķS"�`�`c`8[nu��[@�u�g�T�g���2Xi��m���1��{���D�����V��L8��Pu'��s��+�d��l�8I:�ioO��ڏA���іz�;��́��$����<���m��w���-��]��[�t�r�P�I&�e�O4n3�*�#���;�dp=�1�,���ݝؗ�g����,נ�O�V�#�2$|A�1�Ft�l2����Xܶ�����O���i�?���h���H#2:!��1��F��+��>����17�Q���S�Ry�t�1��E$�@r�,�w.+a�k��A�+4Uå6]��ePj.�Ǔ�~����hތ�ِ}{�������d���/=]�$��LA�ֆ6�P,��3�}����Ì2��$*��| �\3����C�Nއ@Q�<��Lft���u/���Rw���Գ!��牄	p�M<ߺk$q� )�9%ޜ�@�j܈�	"�%��I͎*<�Z#^ ��*�����S���v]��f�Dx�/� ��9�r��Ca�����H7䷶�$�G<���bؑ%��R�U슗�Vs!F-�b�M�s�J'���׀I1�}1/�N���`����['vt�g3�!��L_gD��˚y�R���c�\A �F;��!v�L�ҡ&6�p����Qvw4��u��X��c�n��k����
�gW��XAb?4н�U?8�q���zv�GN�n;�7	�΁ �M�s�>�p�`�%�p��Uz#��I7ս:4lԾs�>�׀O����L˴�gxz����%�.��'�ᚴ.���A ���I �#��V3.D��耙�ˏ�)ލc��W���x������U���|��<m� �E&x?5����_F'�5���7��!�r�Z`x��V]���PN���&y�<z�/�;�o���SˍJ�N�T�SK��ύX's�.�g����y��/���A�|N/y,�Ӌ���ӝF�����HO�[!l\�Z;щ������7�[�֩r�O��;�ȝٷf^E7}����,5<D�a:wtq���Ė��Ik�;�e������S��������՞�{ϰ��������Kҷ��2����{�~�tc�9�2�u>;��N�\{;rx��9L>��-`m��9b[�wW�g�'���=BMn�K�����Y�[�s�{.��<���=�n�_�`���^\Z����yo���x�_1@0�
���We���3Zݞ�ī���Æǡ�����s:׷�1E���w�>�4h3!��ŋ)Ay���~�i��������6����ss[<d-C����{���I��=�Gvo_y/l��ݙ�}�z�ݲiۗ����!#ǚ�\���cyLB�vf�7=�vo����ۢ)V�5��w��7��؋�w����:�
#�+�9�������S�>��F�8�);��6��~v\L��G]i{�t���w���ino��F��yխ�FO�#�=�*@g�ȷ��3\K+�r�֝�+U`6%�Ʀ߫�pk��r���w��	���/�ۼ���<fC�셓<���=2i�aߙ������qSTM���~�^?���������ACZB#�Da�b�E�u�|A�S�u#\��Uw�mF�9u���g�;,�f(�8Y�Ye�kM4�2��ZIJJYe���x��s�=���ۯ�Q�mtݶ�^5�E��cZ3lc4[j�l0�[v��MkIĶ(��n�|�����l��@I���>������u�e�kV��%VeDXe�zt�ۧQ_Bɴe�Ӷ�S�ol�{u��6�n�N��"�#h37e�75��-���n�|���@��Lۈ�i��vne��'8{u��[���+�&Y&��ӹ�3E��f�sl�kr4��=��Ĳ�m�+,���6������kn�R�$�٩�#KE�tbalۦm�ܚ֒[dN6Kk&ͧe����m�ֲn.Ӆ�nq�S�ZH����3:�'m�:ٵ���I��r۳m[nr�sg,��[i#��ԧm���3��H��[]�f��8f�&����;%����7�xۤ���ȒG���q}�:��/����o����	$}=�L�e�휧	; ��L�c�w66����)c��ȂEMwD��|{�gՁ�g�%T�p��6�� :��6�8 ���S#���I>=�0!�S�ok��He��C���I$혍i�V��	 ��I��L���ay�XP�R�T���i�5i��6h�J�n��
ֱ������ݝ8.����������H�혏�u���=�ON�A���0�߿B�|�^<ouߩ�����]%(k�H�I t�d�$����^� ���R��D6]�<�@�d�6�k�"�2�zd�AWmG��o�W3b��u�^Z_�웾���Y��gt�gg� ��h(u�2��"o4vk�'ĂI�� �E��m���a���f�6�������X�!�����ߓ�{Or�{�u �ϭ�BY�������0�rh�b*����#s;�e�m��E���v�/�/$?F3;)�|�[#��b;�jd>9�. �]�L�O���������l��q��TÃf4w]c���c�V�X`�����"b�jn%�5�ݏ�~��{� ���]ݕ�2I�0 �9�x�k��)���1�6c|}�� A��nŝ���g��\�q+#q��n0�q��p��E��h�47ln���q/�ܔJ�b� ��h/V ϐÓ���M5SL�;2�~wM$��w��8�a�җ�1."Z�9(3J莍��e&m�Q��P!u���B�g	'�W}9���qEN^O��)|�����p�:p]�3�xGM�G���ͽ�62^��c>��W�I�-�h�~���TdXK���+���n�z/>?��u�����ʕ�������y��57�|��	�U�X3��!"
�Q��'F�\�N�/)��d�?�Q�-K���K�:܍pe:�����:�)�1�Pu�1�/Z0��Jg9�aJ�vv�k�Mq�f�sZG���,���[F�H�'0���&�.5��+�Y�8ٗ\�MfB��.��.h����:�(٫�f�m26����C�ڑ�t�E��U�5ill-qF[l��+`$��b�����J洊72���Fb���kLWm�#�yI��*4q�b0��:�f���&�m8L#�Sp�L�&�s�h�~����]-�o3����A;�����F��L��.�۵�t惛�[��sd��.\���z����H-0�B
�헑��H�Q��A�3�#�K��=���v,���"��]��	'wo"A ���w����Aۋ@��Nn�'؇�x&!�$��u,#���9�5�	���I#s3f|A5�K������"UT0��Iqi"��A�	���$]��&l��WsTn�c-���L$��w�Տ��D���ȵ�Rݭt%@�0+y��h�hƛib�������0ﻼ�rfw	��8g�����A׽�'Ă~���w Suv��v�/޾����5����[&|���݂s��4��";]�%G�MN4��(wnQ����԰z���B�U^us�0�t�&wo� ND�IOxz#͌���cb�&7<��J��"{�dI�%��=����"+-`��J�3�Y?����ݩ@'�j N�5sf���^�׵� ���Fz�葉�g.�Y0|���O-YQ���J�[��.j�&�ݘ�A�-�f���m��O�*:C��Q6��=3�1�'<��A$1�����yK����<T�$gm��t��G��lK�W3��@�A�1��r	Kc+n���*�Ë�K[�v�)ql �h-m6��Os𾐯�t�M��=���k��	"Wn�<��9!z���Z�;�`y͙�A ���;�2VY��N�3ǔoXi.[�n��6O^�@�����3�v%����Y�KMM��t\�����>/�1~́A��!m|���z���zɑ�]*/��P͙���N۰)��}^?{ߞK���3�~|���aþ�TEҹ�Ek��<u"rcڲmٕ�Nѝ���w��<	/�� �~Υ�哰L��˪�l�T��s�� 3�|V���I/5���Gt=�rN*C%��� �VG���:$ZpY˧�<
�L@�|k�:$�Ѩ�Dh��˘�!����>���]��PCza[K���b�����6���1�#.�1Y�ia�F��Ft�$Ǧ����D�� @$5�Ǡ�^Fr{�A�N���zb����w" K]k��p�)h �PA�T"�zd�Ƽ��8�	�ݽ�[k�	%���ޱ^���9;���'&es؀�c���L�3�����>�A̎��Af�N�f]�*���>���1�n윗-��3�I~��λ�	��8��w[5�9Iݕ��i�ۈs��(��h�gȊ�r�4ȥ��l;L�����8mYxl�����ߟq��,�����їx��R-�pʦ�	��S�:�?���Dݘ�|H=��cJ����+#	�˞�>�>=ݑ�Տ{�.�OV>���=��'�~:��kh� �d�V�΂�46�`Y��1��T��:�\k'�w��=�WN0~�ElÈ��ؐH$}���oj��
�-��u�`�θ�7�rd֒t�E�ك�<�n��h��M��|I;Y92I>;ݐ#ǳP}}��e��Vy��C�\Ă���(3����}�&���Ji��KEA�����I��&@ ��vD/3�]�l���y�w��}aJZ��);��SQ!y/ٸ�Ae��
3x�:�H�t�eTN��}�弜�v�U�s�� \�ck�u�x����6wO��號G���D��	�����Ǣ}�Һ�D5&��M̜,�Φ�N(�̶,�2]6�����سw/��｟�n�Ə��X��d>ǽ�3TWe0��
���:�u������F`ѩ�M��% Hӧ	҉U�Yk��gI�S��L�,\Č!�f����#�]h�+]13���]�]T�[��u�D1�xf��&�¥�X��
Z�+j�B�in����@˺��(�z�t��ՠr���K6hJn��҂�邑�c{f�X�8RY��h�,Ζʑ���RiWQe���T�0�ʺ��D���.c,m���*cS�ٮEf�-�{M��в�p�AM���)����`y9I:�պ���S�ˮ�[R&���ȀA 2��w�L뛓��~������p]�f2������(�19F�:(�D����Az������W�
pe���Ԛ��9�x	�$�F��	��7��{��g��jʻZ['wĒ^d@>,z��G
s�Ȃ��%231<���ƍ���+h|
ژ�^D�Z�����9U ��T@C=�8΁L�8g�,gz<�s�v$���n��i}ٻ#p��؀!�u�A N��ɸm�*:/n(� ��~|�.�"�na,�Z����\n��X��:��3�]�]���~��#������=y<<H,w2ߗ�$
��법a�-O�3K�dĆYZ�25V0N�)���ϲ{jd_���7EL��3]��z
��o*JӺ�!S��7xfhe�33\S�g��O`����'��ΛD�t�3m�3F5�Qw.��~>M{����;Z }]?L�NP� ���/��=�����vd�������{2z��6�Z�w�w	,r��������cRf���;�(�z�e�t���U��-��A6mT�'Ğ�;;M/V�NU�x��J ˸D�Fg�g�A>'ƻ�=����ʃ��K�$�l�J>'ǻ�}2�*V����9A�r�,��3"Ȧ�T6�a�\k��c�f�\W�m�h�:VL����p������'��,f��	7�;	$���o���4�͖ح���/#U�KĆo&p�]��얕��a���/�������uǣ�x���~�k�T��H�7V�wLO�.��vc	$�m��	2�o�4jt��Z�H�YO���c��xz�<e�X���ޢvyu��c�N�Q�����ٛ�H��M�aQa�䧖0�le�֗n �랟I��5gE�N�.�Ƀȣ��v�y�J��� ���O�>#{m��|�o�ķF��6A!��|H�}I�3�����N�k�Zο4O}x��X=�wA�.!x�����S�Y��;�&�����M�t3e\���\�p\�m�^ٖ�M��Xp����t�"�3{S;S#�6fvdߍ����Hnl� �w×{۞\�� �Gn�zd��B���fp\3̂Ҷ�x�1��>us�Q �Ew\@ �}{�$���Оi��}�d���w)�.�!�;L��t��	��?&��@�)��0��|����W��I�s_!�b�"Θ1O�.��{j^f��h�$���Oy��P�HF���4�Y�y��y�(�=����v�^Α �v��г����u�=��;��6�S���]�2�G�?sUU
9���8���zh�	�N
vf`�'=�ܞ�-�&��[ �{N��l�A+�G�>��������ly�l~���%ܢ�������I�n0bV�9��H�f�1̶��x�!k��Y����v����O�����ֻ�1$�Ξ��8�+����x�L��I�u�8=�c3
,��f3Q�72Il��TL��v9�H�5sُD�OL��K�/7w)��z"@�ρX'��.��y��M����̱,6�<.d�X��m�	�ON�骋�w)�.�!�;L��f�e����$�KtA �Y7� �'����,�F	'7�H�1�gL���X�Ω�A��"�^�<�r��� �u� �{�/�&�:�����y!>:��t��٣��)�Y�U�����.M^y7���h�;�F��Q;�î�u�P��v�9[��w�����j�\����E�잦ɹ�;���v�WR㜠�:S<�'ٹ���}�:'��^��ڻΌP�{N���y�6圦� �^�!��.T�޴��=�uG������q�{��ğW��P���)e[�,�(�>�X^��^�������x�m���~�4�m���l���Ƥ\�{�{`��]}t�/���� �Eo�3Q��8��G����!��>��l��]���8��)��q^y��f*��4�� �s�����>�����Z2���kr�e����n\M�P��yfΞ�[�S��f�<���_jx2J���g�<ʓnL����h4,�	bדQWtXIW8���j���W��M(zv�K��&	�Q^�C���AC{��le���!��s�s���7�iKܻ�О�w����Z=V�gPH���j�.׼��^^���7��ֻ �I]�7j>�a��y�cO��/cV��J�Du��]/�`��M쀗
����}���/T��G��=�t0S�2Ҭ��ž���4{-H�9@>`�������������:��t}ޝ%Q��l+%�ùK�����*���52����{$~&]����<k.�ٽ�0lWD���1�٣Y���n�+��z�hg�����0��Od�^���w)ʎ)w�&g��,�����2ˆ�c��&k��"H�9�P@f���1���]㴢_+�h���gH	�(|�T8��a����������M�U���Q�jٍ6V�Z ��-l-�v��9-Ͳ��8�Oμ�޻�~�O:x	d��(JNC�e���f�kki6�s�4�q�n�E�ufffmǧ�nݺ�y5�f4�EEf�&X��im��6"s��hwkdMd�bĊ(����Nݻ{Mw�YA��%坧w"�ݚC3���9:3>�y�������nݽ���PVffdVYPva���n�6ݛ�۳�.ֵ��7I-h����6���f'$�;m��rE������8��&�������m ���ll��DK������[�H�,���R��gm��mo���N��j�m!L�j3vn�pS�rv��Yb��8r��8I3$�ۭs�� �hV۶��DE��ն�N��rs�mg��t��lɴm[l�N�Vm��oky�&ə�9 �Kl)e��=b_j���ۡB�X�#5;0,n�+�[.�Y6�K4�D+�4ѵ���@�i�[v.L�
��L��6X�f�33V�x�Elr��]�����dIF�0�vu�+H.{&C�+�	H�\s��ե�9��HV`���I�0,��v֑�K/�imY�4�-i6Ș�s��n��Q�^�GT���Tr�붕�X�(�2�&�^c����c]�Y(��*��3J��d-fX5c��e&�:�1�e�A�ɠgn�Si\����RX�eV�����ً�E�k�R5��j�K��ZՙV��9ͅ,z��v�K�Dk��hʘr�y�L�Ĺi\#LԒ�DَK�����mu�4JX�%�lM�2X�����s4�.�0H��3�Ɣ�ittA����8A�@�]���	ah�*,ep�mؒ���m,Q��Zd@&Hp�[�K,��pdݩ [l˝2i�ڛl0IV�<հ��*�K\¼�,��]�k��ŴlZ*,���9 �4���d]e4�jl�ll�E�Zӳt��
��������n�MeR#�]�2Wq�h2���6l]�$��s,ѹX�YiH3rPv�$+Í��F������ԗvBpAhi+�KB1�*v���\��H���l���E�^ewTɥTC2�`.��C7^]GA�e���9��BiW(&ĭ���Yf�g.B2�a6�0ّ���z�)��]�6l6�l ���r�Ӷ�h�4��1�-D�۪&e�aln+�͒�"&F\d۪��h�k5)��Vś��m�A�%����b��Ś�4Jm�ə��taԔ2����YBXa�����b�5�\�p�ST"���Z���#�×11����4q��]P�۝���M6u��ΌѽTC���B�����
)��M�k-�hY�*:Ĺ�J�$�e�e��8��܋�6��]��BZEXd�Y�]fb��f(\j���e��J��$�[+X��Z�t����q�f+��b)@eV���8��a\2�P�;P������t�f^�aUMv)�h��f�ia���H�1%*G2�j�&���h&�(�MC�v��SW:ư
eU��MtP��l�ש4���CQ3�*3)p=uR.�� �U����Q��,�X���Ŗ��D�:V��x3�4������nYe�6��\�nݬ��&�e ��YT�5�sm�5�F�`�@�&n�����}>A���?~<wm� oc6$�}��Q�7��s�����$��jI��N��!�/O�S�z
��(�aҸ�k0	5q�H$����Y/xn��3��H������grK��FD�� �v@�	9�y��ݢ��C�!5=�&��'{�}
�6ΉvpX3����s��m���i��y+���O��� �w�:��Ӹi�P;�rnfL�u���o,]�LoKǉ-��c����D�G�y��j홐H'���Hm��<�c�q����p������nc͙�Ɩ�JC%��R�Xi��X!�a-2�p������챹l��.��]uL���ǀ	�m��1�̫��C���+j�$A�܈=���h�vf`�F�� !>>|�x�=��6.�C� �����H�-O|c�L���sS�6�U^U�zm	�^�ڜ�X�ӓ,��2m�Zш�²*���S��V��H$^�D�� ��G��p�-q1v	�}I3QIԼ�ez�`A!�[��>'ċ<A�����D�f@�|[���#F=�f�A��.�fa�zo�-��A��f-�*z��eQ����M3N([�t;8��ݣ�;�#��B���3�V	�tK����d���A^K2;b|H��f��a`�q}�H$�v�|H��铓�f��ϓ>C���}���;V�ƴ�yt�@��h:��5��0H�u�QneJ/��߿���D�o͗�Cfdz�k!M;�>�%N戚��#�ŧ9�{ ��!���C�S#':�I��6��ó��2�A&_u�NTwO�������������"`�j��\��3�n�@��ؓ#3m4鈈ȜV�'�݉���
�n�:}4GO�_�'sV�t�CÀ��gk�Wdy��繸��}�,������v�0��M��	��x$��ޙ�=��f�S�h�(�E�+l���=_�H���A� �Lwt�A�ڶi�<k�LV�H")��060352��1�Z�=+�_�<��s#٥�	T1�'�!�����$�I�ڀ ���u�P�;��W����_x���M	������R�X�Ix4�K��D������ZÒgr����]GD
�Y݈�A$�j f
c�gq�����} �7U��ڷ��ų�?�2{hp`���"g�bI$H[�S��%t<����E/Y��	��^� ���b	U�ʙ�/v��pD�ϙ\_W�g\��$�����Ov�Ǯ�h�\��3��� �ލ�R�'`>;2�	���I':9݇F���w;5s,�eڭ���z��3�o�����>ɚ��5��݈�vs�]V<>��Zb�]�l�$�F��&XP;�O���d�7��)&l1�r���TdA$����DE�e�X$�ޙ���ts�y-��8�,�I>%��l�3/bR���J�m�3��͘�1N�)�xN�2N�p��ɹ�;�vǹ�gdH$����	�':9�	���x��3b��d�w�b��.��;�N��2F��A=�,�5���}�W⹥��I͎x�%�2�"�a��	���y��.��@1�1 �����	*&:���l�	$ ��<�O{��`.�� �C�KՕ�Q-������D���|}]�I1ս'��S�u�'f�AvR�@�,d��Ԅ�L�]wD�4��ص���KV�6� ��&�^ $���%�Y7�[3�̫�t��z��A�b�Ο�;��������{=�L+w�ƒ�z��[��d�=���2��Շ�@'����)��4���YA���]n���]C.ea����$��ѫ�mQ3����]�M)�+t٤ə�r.�SP���6�8�`��P���R��کD1K5Z���Z����-dk�D�-K̀�����b�k+����"XYM�w�)���f�����!4�P�6�u(�V�3�
�Li�؛R��Ʌ50 5�	K���Fx�B� �M���e*ih�%٬���X&����hư�\�f�h�Ё�m�Lܓ*h�|��h��)���C(���H#25�G��OoL��OnV�	s�Y�[ǉяa�[0wp���g��yV>]z��� ��Aގx��� ��LGU��1��;����wt���Du?<���>$���Ԛ�o+ĂN�s��>���Cz"���o3�!�����-N�m� ��Ǐf�L��A��|�j/�n��@�p��	��H:!�*�+z�d�~3x��ǢbnxF��KL�5��t����Y�> �츈j�Z�#���"x�
ܛ�aq�Jh��3�u��U���X�^��NΟ�֌�`Ȼ&`�����|E�fĂ	��p�F
�6�M����~h����|N�t���,¡�D2� ����黹1.<n� �
+Q�Y�������8�ry��$Ɯ��Ou-���U5��q/u�o�ܵ�J+۝�^]��11�A>/��I'��= �{��)d��iXO�[�,Ԙ;;���|�@�!]�1�/.#h6���������$��� A|�v[�)ܻ����Q\��dL��c�W�\wdM� �n8�CkW'�f�C�3]]�37�%݈gbX�S>3�/��솾/��v���B�h�˹�A ��Ǡ���<"�`ᥫy>�e0,9b��)�!m��[�ZR	����B-@]��m-��z���X�X0tC�S����/+�I>lm� �nꗡ�u{yì3fd�'ă���ۖ�P.YE�3�7J�i%sv�W�\^�P$�O���{���}~���7wR��~���9�ޒS	�L1h�P:__<Ey��d1�%�rv�5[C�<U�\�U�:o�gV	MMV���8<:�?nt�;�R�Xl��}�ӥN[��AK]�te~��5��ݳ�sݻ�-ݳ����	l�� �ǲY�8vwL�(�1x�ؐ�)㽗%���x�C�oN��|~�;:5�>8�q�!�t�S�ww%y|V���H$���7��tg*m�H���$�Z�$tm��-zb�g���Hkp>���D�wE,+ã5%�i^5�n��îÖ`Hs�uv�w��~��q�K`�헀CZ�B	}!ޮ��k��� Ckn(߰Eg��wJ�;���t(��f�E���v�I���C�_L���L�%�ytDl���y�D76[؂ޫ�c@�dYd���׶ v/:$�#4{)��us�z�� =[�O��2{;����fSY�Q������u��7�E�@D�Q��$wKW%�Ǯ6L)��*�|G�uYG,��W�˼j�)Ճ��߄�����i�W��}����=x��v8K����U����}�����u�M��bS5��x�$,� ��Jj.��1Jd���;��M����,���{lƾ�!����O��{�"��ƽνo��|��q},�G\6�Cc8�Υtѡ.�0]Xf`@d��sj9����op*���~��\���{=�$�	�0{x�#5��7�F	�5�y2"�}�k,�C;��:�TwT@�ǫ�\��#�z�M���A �t��A���~ƏK=��9�X3���Q>�͹	�fK��dܒ"�E��M[Y�`��V�v'đ���������d]�0{�n���z�9�6�Ӟ:���@$�l����m��}�Δ��J�F�Da o�zI��2��b�Tcǉ�g@k�
�I�֍y��݄�l��$e�@�I-M������Ry��SSąB�������S,��1f�����V�?/���
$�����Hz����I���X�9��zfɯ�0�^<7=�Q��=Vdf�(du�E��)#R�]\�)I��1XX��Um�&������J�m� �ڧ.tH��fG)�Y��je��8�Z[(�J��"d�$�S:��A��$9F殅Ґ���ԗ��k�Ƃm4�,�
Jɍ�Zq��Iq���ePI��=�:R�����Vp�60���ef���ph�T�u�fleѣ����X���qLw�U&���.7[EF���S���]�c�u-���<��Ʒ� �Z�r���P���&�".+Ǽ�&Ψ��z�:�L���� ⎰�ߞ�lh��{���A �����Ko(�K�Cots�E�+�.��ݙ�v%��ub6��������]���8'�$�'�� �k2�����H�S���t�A�)�����j�7��^Ǡ�CsU�ۮ��ֽ��b�ax��@��ZB	�d]�0y+�g��'o#�|Y�о�-����j<P}s2�?Z���3������H()���f��m�.���ر"����p�V��9d�;�Y8ģ�;�e�ÒAmW���u��'1��q������O�K]��<�jN��`����H��<ÁzQ���w:����{S=7�r�^0�2��whecA�UD�ɴ�j�^7)�d�6�d)�����Ø�EXr�R���A$�ժ	�=[]3^H�7:ŵ,���|�� ��y��8ww'z��uCM�V�Ԣ�0h��8��sXA#kk�LvSS�3�K`�d�t��	����W����Ƞ!	���I��H��FѼ�z7ĆQ6�	��k�g)t�c7.d�H=�q�i����f���'ܚm�f�z$���u���;Wqg�������&qH�U�@��V$ ��qYp�]SD�����XeZW�Ͽq�iR��>{��ﷇ$��d�O� �{� ����K&�h$�U]]"}{�N0tY��2xs��띁kNj�]���`��y��;>'��u��"��0�ya�#�jN��`��șِH$�I�؊�I;�A���1���"H�Ï���`�z��Fؽ�x �O/bD?(x]�[%�ƁO0'R��9��t>�ͺ���,���M���n��D3���7� ]�Z�ק���k�=�;=���z糃����2x)f	�H�Zm8������<R��vr:a�n'G�6�|:'�=eJgy�ӆP��b\:��'�;�{�`m���81yl�s����{�qLn0�9�e^���^��<r�U�[$8��e����;z�����:��g��g_'��6���}�y��F��{-�/��I� �'R標Y���js	�'ѻۦ���7R�`BVmܨJ��cT���Z�b	I��ʌ3�x��a����i<����Kz.i�~��="St�؂�ɜ&�����5I;px�g��������7i��-��zd-�Kχ����H^�=vg�g�i�F{�=l����pà9�P7�{+�Y|dS�N�/��=��vf�{豌;�q��v�c��l�,�푴�Ŋ$����gq�}�G��v3ӯOk^�L�}�B�<���8=��wwm���؛�ץ�DB�}��~��u�.�:����4㿼�i�����-7|����Ʈ�/rM����]���)'ˇ��_#�y��93�=ǧ��+9��8��}��ww�ԒKǗC�{��gp��:U�j����Y��eٽ}K雴��j|�r��x�r��[��;�+��� Ph����A]	�K=�N��ܸ��}&�`k��73en�x��/��_?�7�o�]��ڳ;N�!5�Rt���\]���+3��=<{}��e]�Y���rۛ"A�$V����e��Xo��}�$�M5�!��qǧNݽ��wl[d��s��%����2�P8��E����J۴��\�F,���ӷn��"���;��$����:+��[���Yĳp��!�w'mjL���zv����MQ]�$5��Vݹ��%)$@��S0�z�yi�v�k�;79���Bt�DQ�6���9 ��(�f��/79Ü��םسR�"�,�Ge�q�fm����wi퓑t��"R��3VZ#��ii;��y�Y9G8Am5��w'Zo//-�9m�e���I:Vns���!�s���f���=��Q^ٶW����ȒP^w��ם�9�����.yz^���m�<^n	ӊ388IN�E���zo�>&���$��q;�X5�û�)�Й,{j�����a����}�>$���ˈ �˫��:vl�NM3��Z]��'b�;P#:7�I�cW��L޴\�rxj�˪� �̷	�-�h ��cl[6T1��	� �j:KXSB���趄�٦9/�3E.ʲY�E;����r�J!��EvTρ �͸�O�e�� ��s���N,�(�ɒ	��}e�$]$;2���x���φ�r(�wr� ������7��{;�tN��R�<9��6 ��ǷO�A�v����y�E�7��ˈ�����r�#NwE��]5=6���TP�^r��YnsA$����S���_����]�/�}'�	ݐn!�㾸(zۋ�,r����>^'Q����n��Q�/Vy�D�K#�{�xH=A"�f7Ȭi ��5m7�� o F��Ag��Q	�;����A=�nNx�����������$5��x���	������F��������$R+�7���npjۆ].Рt�Pt��X��vvUa&�K�] �;��6�30Ny�:�sf �	,j� s�_�����]��f"X���I�m���^�â\���g3"3����)`��h� �eW� �FWWL�V�m�sS[�K�{75E�bC�b�F̽�r	=�]s��`]ɓ5z�3�^��,����mN�	�'E��Ob|z�n㙽.&�x=�|H7s�>;�v�u�L#ɧd�u�I�)�h� K�zp��H�3�� �Mw\�}Ϙ����c��-����'ă���\C�ͨg}�.�bpßf<N�N��9�ʗ�-ާ2V�`�)/��5�ܚ�vY��Հ�Q����oU��0]Bk�����zǨR�b��*0�2ջ�����.ĸbLm?����V��6��B�����̼��Z��^�(�F2�/:)&լ�X�F+L� �0�-�FSltT�e�7x�`���F�#��Rf��-n���QhZ��6l#ae��E�]��d�����צ8؅!��L�M$���y�����77T�ehR��qD!�tkHl�YD�ZMWT\[jc�!l��0�n�P�i��1�Ո�	���y_�=ߟe�U�s�}���Ó^6�"A$�~츀tWJ�<�y�@u9���8ӹ2LnKS�3ᘇ`�dc���Yb�ظJ�6o�@$��E�Ե^��Uӣ{���F�p�,�)3���ڙ �ͷ�H0ʹ��a�5<�̥��o'��Aޮ{���Q.ŋ���љ����D�ߝdLq��< O��67r�����~��1�[3�}��0�tYK@d����	>+Vty���~��"2��H"���B��PmOr��]�����S�`��HMW�k&Řo4�z�rj�L�&��ɰ��}���K�D��D��h�� Y]I=��nAW5��˯y���ۻ� ���[��IE3�wpS��x�S���L�ѷ�<�S1�n���ֵ5˲
��,+��cC��f��w]�	�:E�&�����=3�ޙݹ���Д�w���rOS��dE{�Fl%�w�`G�� ���	v�K��Q5Z�����czZ���'�;S>3����]�@�T��=^Ai��$��ȀA^]�܄F�p�9���ϣ3�T<{�镶r\�CP% Y�� �}���(�O�5G�&j{�g���c���wA�%�p��NX��ŋȨX��A�蓯��\�݄E�驨��M�\�Āz��A�U.�ߝ%1��Z�E���s-6sZ�Ռ�!Cf���k�@K@e���|���}����jx�+nH+l������sR�Bh���6Z�F�41��E3��S=2	 �s�vh���'Įk� �F��H��7,�͖EZ��z�=+�RL�Y�d�Er��$�ά� �k+��9�h��ZhH`�X�K��VDB{�3�Lt�=����|+gx��ﱁ�4�������L�C�r�κ��Gr{.DUf'z�F&�(�s\8�+l����� ������;2A�u2g��X\"1��Z �WJ<I vmt�'ă�][C5	���tt_��qt�1b78v�&s�S ���[��bV6U�D3t(>ˮ��]�A�H��24w���O�<mv��D�t�Tpk��qB⠖�8-�P�b��7O�_s߽Z���>|����c�;'6$g�ǒ���A��W��e�Yx _K� ���LZ���X���ۈ��Z���VbM���>Uu�B|LyW7g�A7�g_6ф�D6d-&��$�0tAS���~$�]\�H+/i��mKe\�v�3��FL��A	�g�wvgtɋĂ�GvI|��G(|�w��$G�$U���@V�˯%������˧mǝ�&F?���B5y�.]Ñ�vt'.���7��r�e�6o��g��+�-q�-��ײvh��J��U+��7�M��L�"�Z���'fH:�L�s�o$Z�d[�`�)ja<�s�����I'��V��B��A�{y|��~�	������v�CAtu��X.2����-."��:�f�8�+��}����INι�c������[o(���-ݰʞ�ۙ �k+c�w�m�d\"�س��R�T�p��>e5��I=���A ����A�l���c|fol���!��e0���J�}x�q�BǳnY��!�Gz��v�G�e?�k���ND5���ϓ��/�J�R��$��	i����=�"�5k��V
N�]�ӳ�u۴"	�5���R�|$7>�A!�����S�2Dw7�+�9K���̋j	�8>�&��vUo����ݾO^T��4�8Z���b�eS�OI[I�����o|�X�Y���^�Z�[�s{S�iI��u��"� L�At,f���T30�&�3��)j�рJ�e
��4�1Fi�68�β�K�e�]�����Z�B�9�\��n�)h�U�������ʯQ��g������P4t�%B�:�K�L����ɉ,��b�ܓg\ks�XP��4�n԰�b����ltP��L�\;\��mY.�6�
V6�b�ӕ���M�/(I�b�i�X��o.����]=���~9Xe	��?P�=�I-z�|��w�A=�9Kk���MlG��m��1�3\3�K���K�t�xr ����Ǚ���	��L�JkOt�$�͍/�c=[�l�d\&	اUF��ߐC�sb@&��=WkvOy
sf��Cgt$��=��27�{�û�`�C��@�V��Նf���f� �v<x�H��ܑ$��u�`P��:١w�c���@;�Zfp�: �����$_\YmK��V dg@Q{O���".b�`��=h�f�'(;��&N�l:�ͥTvb�	��W6
��3P Y��6�Ο?~��RN��˻ ��;�� ����$�F�\@6��^~B�2c4�W9^�����7�>&����fL��u2z�b�����:���P臸�1��a�
���bH92 H����~ߥ��bt����Ұ�ܱBv+U�m���1�V�l��>]{��A�Nlɿ ��d ��[�]K���k��[т+�3�%ٝ���R$>Wۓ �ch�6#�tW���Ȓ|I�눻�\�.�S�A���;24\��ʝm>�"{6�%��MgL@$���I���>F��u��vfD��$3�s(3:�mlz����=OW�5$y��A�$;2 ������
�8�����, �M�Ѻ03�wVf6��Z�̶�b5f�Ќ�m(�xf��L΋�b
�}zْ9w�#��[w(:Ǯ��b2G>�ӛ� ��
�� �'4S�;9wdFykGc�qs�K2J�{���޽�D��	۟��nny�Q�H���$Kյ3�b]�0v�Aꎁ��x����x��O�-w� �i.�A۳�{��gޣ�^	�'�@`I��"ד39�t��޺�+y��!So����S�4��vk�����J�n0	����ù&%�;]�\oT������j�� A+�"�~"��D�f��-��׻�LM\z��4\�.�S��S�$A���{%�z=�Q ��� �gg�d薚�d�A��
[��)vIHV��a�Ɠb&�R�u�nAJ�,Ke��vNY����gv,�gu8��H]m���"r{�OOsl_=6��jh���V�D7�-X�`��4���3�箙�y+�a�t] �suA$[������������Ȝ-���'oo�!��Rwwg.�ĕ��D���O��8O$�KuX¦��H���;��l�b�;UF�;f����c�W�a�ē�wg2dy.���<^�EY�2g
�6�͙	2'vf��j�T5ݶx��_�\��g��W����w�������;��{�v���x�������+�'�˹t�LK�v��"H��{Mj,��j��VsџH�2'�o�2I>��!\�۪h�<���/N1��!��4��MBjis.�T�p�`qiP3:�S~}���:d\&	ا]���L"I��ؐ|Gu�_�'�ɬk�0g+�4D�тIQ�"}^��4�����@��� ��1�3���f�<���<ۨ��	�y3���z��8+b���4x�f.'�SA��d��'�ryQ���ѱK&��FT_L�;ݑ�(������vA�U���.c�<2��#�}�S<�I ���Ȃ|	��e<OV�6]�@�&m�dL�sS;&اp�� �lϢA �cd �ͳ6*�;��P��C3���ϒ} ��\ӧ��������o�^ ������� �*�+��Q����b��_�UP^���a�0���f;7�`f� �H a��PBEA BiTT��c��i��B&EE�tH�f#��u�@��fHS��]=HJ�f90c�So�P aP&��@�b	�i��`�B	��P�Ha4�����b��LL3*��&4���0�&�`�0�CL��2*��
��3�Qpi�EXBa�bBEX`eE��VDXQ`n�E�`E���TXQ`dE��AX`e��XY�QAD<k�\�$��0#�u����0A � P(TUR%�����׽��>y�����CY��������C��������s�����������٢u�_����s���������_���ϳ������r��+��o����y?��O�((
�?x�(�"�@���_�?G�6a�HC����������~������Zy?�EQ�������_�v`u������;Ci��z�g����A�M��5�g�����>��������"�2　����"��� #@( �*$�B�A
��@�		HD	He!PP�@�!%		FD�BY	Qd%E��FYeE�Y%�S�@abTX�E�QT�E�}�],~Ώ����=���L�Ph���^X�G���������W�\��b��?���v?���~�ٰ�U^����o�;������>����s�>�?lg�z���������8��o�w����QTEi�;=� :h}e����}O�L~?�>� 
+�(�"�zX~,x;~��x��+�0>�����td���@���W����}{���:� ?�~~�����S��}O�i���QTEb>�~�0�D�?w�5����"����ڟc���������o_��w?h~���� �}g��χ�����@�A� ��w����`{_�����+{��ߢULX~��QTEp�?������~����L>����`u���.���'��s��"�`;������[�=��>�|�>**��� ���>������6h����A��Ǌ~�����/��2}������}k�E\�c����g��<���PP������^���_����O�!��C���������d�Me��	8?=f�A@��̟\��>X   t�� �� �     @  � �      (*T@ �  ��T�T�J�i�BE)KM/�]��fF��

�[PPB�IADUkDRV���P;:u��T�U��%(PZ��                @                            ��}9j }9�;`{�w��7 �� :'r��0r ��� C'@�EM�ډ+f�|   �<��18�� !����j�误���(���rx��!N� �)T>���J��R��JrR�{�Ҫ�J��U[l�m�p   <         G�)T����R�W�5'�H'0Х]`��((��UJ����T���YT��Δ��sjP�
�;� �
U)VƗ��C���IT	*�   ���tvn`��x ��� ��G&��C�]n :����9K�A��iȕT%"��  �        ���{�)�}t�t����m4/�� ��uho!�oS���.��i�S��W�/ZU�� ;���wh\�u��m��gZ�   ��TO�r١�� ��Vcrc�O6�S�C��ؽ���5J]8 ��}�s��[n3*���][���n�%�EUREC���         ��j�3N�}5�Ϊ�g*�)���y��� �]yJ�=���x��mS�iQLl��� �R�su==�v:{��jIE*U����������ˡc׀�U��6���v�^�yeByg����� .(:s��٭��{K�T�������V�EHT�� ҂         y�P�����폾n'ͩW6R�c�iGF�x y
�=XҶ�л��<�"�l��i5� � ����H�m��"B�)��  �)�k�K���// ��=����b�X73T��� �  "2 d5T�;���>��O!���54� ��b��@  S����R�4���ʪF�R�  T�����T�@h2d0�*ALR���`�����_��}U���= \���X|�`b�?��������{׿���6��c���Lc��c���6����x��#���_��Ǔ �r2�ӛ�39gkG{
|�k��繿�E�)�!�&����l�;��:��:!��7��LM��,��Q� 硣�Nǣ�]Ǫ�z�Z��4�欤k]��j׽���4�p���|`��;�#��q���- oFn�r����±{�H�W �qR�;2�����W��^���gON�����EN��S�l7&!F.�Bߌ��N���X �7�[���ok,�G�jP1�Q۽�QmR��L�d��^7M�ۇ~�\�Fjˮ��u�u����Md7tӏ���[ ��ճ��b��r��O%w�M٫�oh���[�6�b;C����3�JPv�ǝĕ��\�t���I�QIT��|d�0e޻z �L��ÆQ�o#ǥ�d�PAjۮWG������U���Y�ʯH��+�t��IpxU{<�o
�Yn�3���\�.���0>xV����ͻr�Y�a�^���of��l�zu$k�T�Ր��Ch#�H�"�a���	4��`�q�d:A0l,�6�φ�q�֦3Ni�@с��{��E���X'v�4S�2�Gu�"��#ʓ�^�&i�WQt�-�B���-[�v��u�ʝebb�r.����
qcoz���7�!��Gc�,�W����..�Ͷi��́�n-kc���|-����j�-l"攆���ke;�N�ɝ�P5��Mx��>�����x��A\:$��n��VҶj���Kxu%��Ez�<�OI�L��ك���a�y/�M���2�V��5`Xh�o��Ջt.J5r=��Y�,/t�jZ�r���T	�MC��$�1���U���Πk����PlNH{�}݅w�f�$ 'H�ugp:*����f��6i����Yn�T�&�1%��xS�(�ovGp�]㊳��-	���Y������c�6�^ �����Kn�Xϳp��ȋ�Y�m�����e�)Ժ[N�7n�3��������u�����i,��م�/���"�f�%�/Ĭ�.���7�Κ2��;�.�D3x����j�LIcS0�&`�^K��ƓB�x���o �0�OsQ��͏��w7f=v���N�m� ��C�
c����.�����BӺ�:���u�{����N���OM��.iE.nU,�4���Z�A6Hi���p��h��ۼ6��0lҩjNǉ�Fj���M㗈��&[���2����{#���[y͜�M� ����׸{��옸��FO`��kK������xܝ0���t*��YL|w\N��[�˾� M��٤.ڡ���	��sy��sժY�l�(�cR��i=�6��.(��bq*w�*�{I��%UkV�J�Hot)؃����`���[�x L�&]�A�t̙�Er��G&q�1�r���f���q��=�76�8憆�{�qp<�<�U�_j!����>-�lM�4�)�qB0�@��)z�" a��g�TJ{��j=r��+�]�6��sB�-���Ʃ��9
��7T�o̠8�óe��ʖ��e����J$)s�lXǵ^�<�]#NKr̈́@/��>pv�^��nÏ�Pݚ��݇x��ُ:5�q�t���6�,4-�UۧZ�^�ݛ�gV�Y,�0v��c��3�=�m^
�;���r�n�WG�{G��J8����	=.�-��!Sw\@�\o����ѻD׼քWnF�lV���5K��-|8���D�*Ű)����.I�K�gNV�On�E�	�/2Y�z���t~�ͽ��]���(�'�M6m1�C5�vvz&+.�ܴ]�.wW
K.wq�R�K��S��n��+	�z�:k���R���H���� }��8�p0��uo�c�ؕ�=4���;���uI]�����.8���侈�F3e�������8с�C�@��涮����
�e�Mݮ<�g-�ƒ���lZ[S����x���z���`asw��&��7�[�;gp��s�v�Ydlv�a<�A�Z�.��<fCD�-HoC�wG���d̜�u�/SY�b}�4-�J���\k^��P��!L��
��9��bZP!H��ٵ�����;��ua����u�oc;۪� �輋P��F�7�79	�$��r��U��r��pm}�vd���$0���j��Y_o;wjӃ:�f<a�(�z#Z�	��_p��n����u�sbG뮽��{�ob'��j;�Ս��DnP�z-/{qJ�5�����%C<"�BhY��yb���ם��8F�sF���.^/p8m���y�n��O^�����M���rI�>D�f�m�]�a	�f�{y��U�{3���^�s����3To\o�d鹻3���kT�]�[�*�`��� r��\׺0�Y��0FQ{��y��,=�ӟo���Ő���B;0Ϗ���Y�bdD�xL��!3�����ϧvZ�m�Ь��׃%0�VIc�l锵�n���<�צ��K���+�m�����׼�l�{�wtML����J�8wi��`Q�����,�p�O'��&��1�;s ż��S�/�r�����2��Gh׳nLY�1iz���9mZؘob᢮��[�ow^��aC[��N��l�!�9� ,��7;R���{�m���z��4��#�T�n�߻t=C.os�gi+4��t��]7�o<���ҷX����H1��<�YتV��R24��Jx��熝5�p�i�H��Ў���E�g�H�t+
�hV�.s��\Ū"�tv�
�=D�g=�a��Uչ�7�{+���CBo�p��e�Wa��){�v�y����a@i=�u�G��~}���]F�֩Uw�sWxv��]�s�ٻv�%�B=Θ���i齑���F�G�L��� �d�Z��7�7(��Y�"�B���#|��&��\�unō�s����tN Qf�tg<� /�!���]��K;O-YȰ�ࡼ�u�ݝ�)3i��nn��ΌzG=͋+wV�5@N�#tǑ�y�h�k�T3�b��[ �N�w�J*'�V�����kQ^�ow�-y^��n��\UA��{�\7iľ\i����j��v���E�֡�J�X$��m&�����0�Ȣ���Y^� e:$k�INe��vc�K��P�
wuڜ�{K�������w��q{C�BFܨf��
�B����qd�v��> �,'�n�VU{.4Cb�Y�Y������L/g�X-=��m��(a�{�$�(˻ܫ1wM�ĭ�Bˡk�RBg��޻����� {��s'\�'	�9�:�=�E]F
oC�!��~Q��v��2 P>�{��Q�'��,#�j'���k�v��$�s����ǚۆE֬F��������P֒4٫�g.����L�X�&���aI�r־�7@z����ϙ�$��m4b]^��p�;���1�x�����G:hX�t+l�튍ٺg]gB
�&d���7n,P���p��u��u�2���q�N��RY�ہ�qJ.kJq���l��(��|zl�N�zY^IV�wgt]wɰq�1���!wg7�L$�ռ2`	efa�@�`0�gr#M��ۈ���)�#l���n�͋Y�L4�i�{��� �K<)�Y��2����E*O����k�\#���;�I�'o�`�#�H5v�_;]}Ѐi# ���#���Ha$$���Z��w
]Ɂ	$hq����4@���X�xѿnmOx޹��>ƗF��w������{rF�gy����'v�_7N�5o7�,0v�B(:�g��1�5ڈ��Xba7�z#ma�1�<�i�$�����]Z���bn�cP�ad�Lb���I�����+4r��M������϶t�2ݬnM�'��R<N7�Z�7/e���{���:�&�w�A����l(�D��Ç���f��gs|r��$FHYŮ�(���!������
�Y�vY�Y�rn:�r	���,P�:�r�'82j�n�kd5�`װs��Ն�AZ=_�x��"sY�r���5v�,����n>��1�u�z�eΩ<���}-��ӂ��(N`xV7�ә�gZ����020�/+���N(^�{��rMٌ��m�fť���Fq|�N'.-�O8�u559�{��(o��[�����{/���W�S�bt7��ı��w��wH]/ig�ά�MsZ�<u���gEg�\�.���Wpg{��_ =Z�S�Q�<��CN�s�g>a�]��R��;r7�qt:8�3{y����wY�9���X�U�z��kt��p�W1��h�+ʭ�FT��N�!�Ni��r�YBa`�N����XŐ�kܧWwP�z�$��ŴwM�Id�;��6�(�s��tG���pJt�L,$,C7��,�`�k��J��#�R��d��KN�B�u��u͚���Mn��p�]y�5|�7���f�ʟL�#��{P��7p�'HF��9�aQ�&B�h�.!��x��c�	�y�7�A�Niº�Ü�I6�뗍��0��� � S�x=r�:�՜�Ę����Ӟh�R[�ϩ%H>P��;	"���B�uJg)J�a@�����gr5&���o'Dq���"~-TR�y=��Ԍׄ�6�6>��7�Bl��6-{�ux��!cG��\-�p6��q:6���߂K��n��Ԓ ��9q�� 2�2�l���f�M��ۙ�5v]w*�y�aq�����tI��M�W�j�A�Hp���ך9�j��.ǰ� a�b�뻋��)ބ�����d�����N�C��ӻ�).����k.�W-�j8sHƦ����¦��Y�Q���F�Ӕ�ۋ�!�����h3�\ظp:�&�C$��au��!���a�(nD�o:H�yLӿSC3;{8n����_2�z��{:���ܼb`����v
��LAKy��� �C����t6��D4�7:A���S�M�Hy�4]�-��N�=���ӻ��GgY�7V��ǓT)NT�N[�4��ިe[��	c*e���d��cA��K/9���l� �Nu��T�Ov;����&�\��|�`�י�5��nV�<z��U�όK�l��M�^����Z�n�8��6�	PW�3)E�˂�guѱ�Aqy�p�����d]�C�n��'�u���m�T�L]a��N��܁�ރ�GÑ�d��cV9�x]|���{Q�$���콻�$2���+��Vܫ8�[K.e�o���l\���-�t�6��w!tvoL��Ʊ^������((�;�Yd�!�E]:X�ˉ2�D�ʎ1���y��7�g-yٮv�R�zh�&z���S*�#����7{x<����כ�՘����-���Ԋ�uxս��c+7ثv�^�m+Z=�h3 ����Tx/�u��Lg&$��	����F%��1��[IRc�KQ�/��o��U�l���7�K<�
4@��bEs%�ظN�;:5���ʴ�~���;����Lwr��-�9ЯU��9WeM�կ^�c���0�0�O�����.�3�i�aƼ�6���z��r�Mw^Y-7]��5��s�J�{⽧�Y�k���{��='5"9�0�1�|ى��p��;i���N<i�0�NJ�����Y�ї�8��Xt��A�.㾃�T|���Ȯ5�JܢW&�;<�W 2�=y��K'f�xv���ư����{�����oCg1�3�N�l���0m�7��mv��w�F��ODr	��
�E�[�B�A���Rxq[ُ�^ً�صj�K�sY�%c;���0���ζ-�'�c�N��@��Wط�2F2B)�e�;^HD�{���gsW��gtcNoN��v�S��Q�5��W{dԹ��/��`����������r��R�>�\#b�����O����U��E�ۍ�u��*曻2���9���Q���g���WV3�^�Sn#�ݯ�g�ܼmX�9Jx��,̓���o
��v�I��ºë��%��L��1ER��ЁB�t3q�Rf[^��;������0���t����F����i�5��γ^�ӷ�3�h��OO8�wd�i�9���ͽ���P��o�2�>|v<���N�����As\3EǷQF�WU8���G�'��?N	��ΐzFִf�{��7�E%�(V���.+���f��.��8�q\�n���
�us86�\έt��.�ͪ=���N�i���+���H��"3�#�%��9
{qK���ζ�L⇾Ӭ82�7�y�v�ƒy��x��]�C9��Z+���qq'��y�y��@�-�maŔL{��s���� �Ԑ�m���l�K��:���Dh�'r9��;P��n6$�����G���V5N �^��PdkK����6���J��:u��(�է;�OF�a�,y2���������wl	=a)�VftYs�&@v;)��bTiƺ��N�[�q��cY^�oR%�M׽\����;��y���m��c)��`ˁp�.bM���a@6c� �ěe�l)�m���6\m��\l�N)�\m���v v6'��1��CE6ċ���������v�\�( *�i�*�`Ă퍅 .6�����6@0�S&0N�2�c��e���2��'˰m&�v0�`� �6� � (m;`˱��ll�0bq�
p�Hm��e4�����p�  �`�ˍ�.�@�(.��m�!�&bp e�4�6S (H�2�6]��(c.6?������l`�����s�}�����}����>,��l��tl�c���݇�qȹ�D��Pqz��]��X'�#�p�3�I���<l;�I�:n�ت�s{�>�̗7&�xPC�s
��F(��~�°x[aV{��r�}�_{/�F~���bzn����λt�ì��)���A���=��[I
xH� �f�r���]��.ݫ=������O�Qx�
�O�w��M�!y-��7�{}�=��y*�iO!�Mq���F�/Rax����HW�y���$���Zpol��/7��;���/�������jxǷϪ�����(J�q�}@��>�^}]jg<���[����L,�j�ORݨťWv�����}���	}��K_x�㖼�V���7�V��{tF���z3����g8��>���ԣ�n��|+O/˥�T]�f�>����b�52�P1x��M��F��l�y>)������@���1�x��O��9p׾N#��r������3�խ1���:�)΋G�z���ΟM	*��N �C�:e^,!�z9��{D�eacu����/�f�;|���>��X;���V��ƨb�
�ڙz�>
�y�uaJ��=����pL�p�纤c@�JΔ\���@���_m�a6�ƨɆ((��:�n!����X���>귫3�;[���1s�`��[pi�9��6��ޞ��P�{^w�>�}�V�h�~�����-�rw�s�W�p�8k��<<����O��� �#��Z�0�뾞�J��h��u�1�=�U_=/�ê�[^��bU���,\+=��y�'�y�j_Oq��<���<��L ���c}nBG���.^�vt<�����B�}"�m���un����'�� ��^q�=�qf�ST�y������~���V����Y@�}7k�g{&���oe~,PL�V�eA	Z�Ĳ��ђ�Z���W*ԑ.��G���[~�c³@�6z���v��S��{��pV^�U㯞��.�n��3D�32�#ەTQ�a�̰���\�_�C>�g��<���,p�oe݃:xPF������r�+�zZW���=�9�JO�0�yv��߀͔.�Vs9�u@�xvR�Fᓚ�7���:��r)w���.� %�s��M�^�?C��ܝ�hqow�d3��EDܨ��W��mm9��y^�Ӿ��`�9V_v����8)~��&An�'���M|'�{I�������Z,d+��Byw��8m�ga��b'�b��k�3M���H󃏣���XG���2�63�l�@=�W�Zmܺ{.�~��z������������A
�o��ڵY�9���i��:�f����*��]9C@�=��ȋÉ���\�~|�V]�Qy�ټ�=����I:��$�[�c���Ϋ����aٞ]�.���D"x~}+g/�\�Q���j]�:���b�]����}#�<<�pF~;�/�[����e����BH �R8�P�-<ﭚg�'yM��w|���W�ypJ����x�6;�ø�+"A�W�:��Dd���O��S+��|�qc��D�^
7��7��K��.��^���r��d��0
_Nܡ���ˡ�G��O	W�7޽��':�$y<V��&`D�>�w�䯯�'Ao$���7�����@�Zz�е�k��m��ӰI��~������� {5����7��vZf]��Ϊ����C�x��� ��{���b���".�������h�~/���=U��P�!�ud˷Ǚ�c�n��cm������	�ϴ!���x�z�zx�@}�kc9F\��w�v?3�{�Q���y�FX6D�uL�y�	&F#�i�[`���`�fe�Mg�Iw��isw���� �{[v�p3Ξ᳭��~��4�����Zt �L��O���j�Եw6[f�w����6�;%ٞ�R�������G�?G>a�Ӿʼxh�n�_��p��4v��n ���d"O΃q|��}�Π��Ө��#*�"k5��=�H�����J"6�f�`���ې�\t����"���t�8q��� ��ܜ����8�'��k�N�'*�OZژ'voT]?Y�=�7�q΁:O��+9�]�q��.��p1Ös ����g�V2w���j'r��{a��v`��z�X���;6;���7'm<<��3�����a0x�y�p������w���6�v��/-�৞���_�O����L�d�2���֌*RN�h7�]����4p�u�=����	�(��<���z�9�О�ʇ�\��w�����5�0�h@�t��h/��n��h�a�^L�i�\モ�:�m/xz�BR�����
C��@)�������W�>�H�Z���>�8�o�ֵ�0#��:[�}��R�����%o%5�	��CP3��� �����t�3�(��,�;{M�f��NQ�U��=��)�v��A��%|5��>�<X��R�.y7e�o˔�^�6�^��k;�8��v{^���a�JB��g�4	~�c��<��ؗHI�����{��"��c�cY��dG���4Q7w��{.]�٩�?w�^��'&�&����.�F�<���²������\+�/kŤ8��G� �TZ0��m��\g=��v���fu���;��upm�r�9W5F�>�-�<|T�	�^�;�#�^��A�/~�/n�X��&�u������.5�4�&T��������Q���-�}8fD�L���G.���e��@y�׊�Z,3��o-ݘ�ߝ���a�3����Ӯ���{	]�.���z�6��{6��y��wۯI�)���Z�3�m{�>�"�r�]���X���h��z�Bo�{,0$��vF�j;p�}kR�x���u���
�
L<����[9�V��V/��>�tu[/���e.����{�v�un�Cp�9`�6t�FL��={��<�V��Ƙ�9�Q�{p'�Z��s~5uw5l�q[�{iX�;�kb��s ҔO�{6�J`��n��o�j�}�iWVY^�(Y������MT������5{9��U�b΃��~cz���}f9D�wcan�^b0K�ט�V}h_����hG����]��,,��21-������\X��X�x#�o����t�ܳM����@�\;�r�&��td��*T�xW;z 2��_�>��[����^[e���Yx��Kjb~'�'�tW"���b�鸐j	���� (�hj�1,j���Z�AVn,/A����2��#ϓY>N�^��p�*�s�2�-;�s�S������f�~�c�H;b�y�Yh�Y׆͋Y�V����4kbi�2����o*��KD�{�6�FMO=�3g��y�S��h�/De ����X���jp;�T�;���08�Ջ{|�ݳ؎Cza�Ǥ�?e���&i�¼x4�v���_n�F��_a���BW�� V�ˣ7����ɭ�+�#�+M�n��8KYq��h]p�#1����������9��v��W�$�K�4�P��tt���Q1u���W�A���ޫ�)�Nx�m-|����:����1�H�;�懆��r�tvl-�-z���+����3Y��5�
��R"V]ҢQ.ɹ�x��fvq�i;�U�����Sݶ��>vf���$�����}���W}=��Pt:'�i �x�m�����NZ�0��=ě�U6�v (��=���c�8N�6ջ���oy}�=��];P�]�G���/��:�?"7ӻs[&��.[}�x�=ŪfL���zz@�B��!]���>�p��I�����o�q�#���w��3i�x�@�:�%��B�ȃ��Q؏?Z�.��:��C\���w)[7Onù-�m'dkw�_)��P�h>�`�]'�����3��p�kqGi�'i�;nk�/��wѫ'O�V���ZA{�Q/�+��k;Ҫ}�AͰ���:�o{]��-�1 o;�=�s�aws�uO�l��u�V ��뤯,/,�5	a�u3���{�7qw��ME椤w=��˂�r&bw��Ξ�ޑ����:H��I�q�@cEB*��t� ���z��%����\�R[�2�"���Α�bڄ�R0N�=<&�Z��6�����(����Љ}�웕����q��,Jo�vN��9�ñ�'��RK�?7��U�c���]Y��m�|���[�����
�6�T�7�x�����a����,����{�>˛Ӗ5�ni�I�õ����Z��{ɾ��`:���;�{,����G�y	A���湤�Ӟ2{&�9�ң+Yb���µ��K/E�4{���"3U�'}��&�d���;]R��u"c%{~-�Uؕ���q0rk�Y��{:rc�j�i.�>�*��`��9���A��?S�+�>��s��/!��D���xv��3M�{��w�C:9��j<�ˢ���X�ko{�����V�-��i�MZ=M^X�H��?c�����T,��q,�Q�fL����r��\�����/מ_u.�6��Қ&�X��#ӳm��9v�����+�_"i���ڏ^
�&^}�h��);!h�aS����f���Pݳ3T	
$W2��8dP=�y)X�5*�>ξ�v����Yb��������u��^��\�U�m�Rp�6!�Cx{���TmLT���99M�-�������C@�&4���1��7����!n�.qy�������В�}�S���?v�!$Yj�;8.O�=��n�ec�JuOvsSm��*]����b���T�C>>k���������SFq���K�q�.����������h|bѱ�2�ǎ,�p����O�q[ӻ�P�ɾ������Y6܃3gj �Ԫƞ�3�:�������w���/|����L��ہ�>�x�I	Ć���sk�O:�
S�$���m�����Y�ӕ�y���GqM�k��:;	*# ��������g{����xO>��5��N��i�I^�=�����z��M�Q8��Zf+��kM]�=�-��-șb@�|���y��ͪ�e�ԭ�r8��)U_^߼�R����nt�f�M٧�6{CR2�;�3ޤ��>=���G�ؑ�*к:�*�A��h&��rS5��A�3���w�<�XeGh�&e�<Lrb@�۠[�FDA;M������t�� ]�p����7_�d~��Q/h�̑KD�Y��-�r#I�
}Ϟ�ݸ�XZ~���g��<��O�]�/RV�^|yװ1��1��]���w��Ri'>iâ��J���3�=����h]:.��ѝ���Bƥ��#�9=~��|=���|��$�|d�h<���b�ۓ�?��@p�Ԏ��icz#���;e3�zn_Ck��*�]>]�`�6�=�
�l.�c����0�(�d�ԣ��H�{^��F���K���>��㮝�����eQf �ua�l�||���}f��6�'�l}���L/N����u���u�jݽ��f;�����CC:'���ᴾ�|��,�v��y�q�cL�����e�e�B����o�S�����>WR��F&�knh���}�5{gU�ޓV�#���]�H<⧖���w��4)3*(w�]�4�v#�s����qg����
i�� Y�G��b����N��kٲ�pm�xtZ��\����u�
�{ψ*+ovL��|�\{m�+�O��M�+o�����
����=)̮�ⅿ_C��@?����9�8���x
}�M�R	vn%޷:��g_x����(Hw��R���,�2�6\�P�������\yp'*�����	;u�A��ĆU��c��|r[����ǨVގv�\�toZd�����'��L�[�o����F*�����'�6k�:�Z�t��(��~ӿ>���_J=��#��j�q��3�'����k�:�Ǘ�b�j�p������q����^m�|���Q�8���wի�.-N�*m�� ������y����j�,�q����V���1	�{���KPU�oK#/F��r�As6��Y���R��68u���FRn���1<�Õ��`�gy��J_=2�Q��ܗ=��/�a��x���=p�=)�@,i�{$��11�^!�g�`�%�;f#���`M�_w��k���3M��^�z��B����ʍ�s#������ۼ��K۪>�9펆7<�#��>A�E9�Y�2F�d�u��]�C;�v__up��=��q#�A4u@C��Zգ���w1��&��ynr>�a��m׫73��c��M�	���ku��ž�pn�=��p�IQ8����#���ɔ�����|�j�4�|����I��魜���x�9Kj�42!�*�e���* ku�.9II��o|W}�Aq��ط�n.�?zTo^wX�y��>��z�1���Y�l˃�Y �P$��}q��
Bx���a����;��5c��k�}��.�Y��d� �ti+__G��75���	�`۾7�l@U,��؛={7 ��m��#xyT����2���M���Q1N^ܝ�|U�͘�2c#mc�'o�P�^��Wny*�W�~>�ګl�w����=��_�y��O=��Nn������$��<��{�mk�N�ZR��*�*�hg����r�����#�o=X^�[j��������cT��KkUU�T,�L҉y�-�ww�%N��½ȷ���t{�#�U傄�Qt�3�
�y����l`�}6�_?����.���f�κݫOO��Z3�܏8�{wa���봎�U���mg\�Tn����g<�c���o\�m2���j�pܸ�2;v�pG�e5���{
v�녜�[��c&;;[��J���m������1�3@��s>��s/$��۞B��6�m�^[r��>g�]ظ�0OV67]�-���[�M��c\�K�]ט�8���6�(��h���ӗ��+����tq��kv{7Y�.��66�q�N����T��;�`w�K7 �y�v�mڪHz�{;������������<�n���ɬ����rn����+��E]e�7�#�;1[�%��v�ޣ�J�j^�[��=��s��f&�*u���S�v����Z��rA�>���98���@n�m���`ݝI�@ƛ�x��Y�쉛�<�s��IxY
���r#�mvb�u�Zx�m=g'2������7<������8=�a���T�bq���`�nx��谩O=\��M�\���/b
;m�����u�9���q���Y��)�tzz.jƞ��	ޢx���S�SOV�l	�a86��۴ܵt7��W<�ݴ���ws9o����c�O�0�+ˆ��a�c���X�;�{o�À�[�
7N�pN޹��gm��a�']c=WU�vOGe��8�u�\�0��]tj�OmAWc���8��絯bk���g��6�ڥ�Oϝ��n�v[.h<�}lX���x���nn�q�!��-�g��}n�����۝�H�Fn��][8Z�y˼�/e�f�:'c�����ؙxDMSF�d]�L7����Z睲��=�BK���]�x8�]���lwcE�q\vA�]���!�=#<�Z;f�׬���-�xK�%�o]�m��E�.ͮF͐�r]�M��y��wD���[����8瀮ՃZ��c��X�!�u�c�Q�3���؝�s�j�6�j<��{5�x˜���-W%u�qL�;M���G�p���rps�
Ϻv��k����j�,
m�{]���[�\݆��rq[íW��w7<�7dpYM:Wz�A��ݧ���r����5(�lh#e��lmD�kGk�v���>'�᩼�\=)�5�����p�zn8���d��.�vk�g��CrK� �X�9���-۩��E���	�-��4�G�wW;ղ�i줽Tv섃x{&ې���i�� ��!���H�bb�;%K�4.�;[�Y���<׸69��	�m�wn�k����^�ܯ���B5����k�޺�`�71�k�͇�Ǌ�'p���'�u�m���h+�!�.�n���7hv�@�x�ظ�Q�<��v+��\t�ذ���*::������[!N�g��v@2��ێ�ң���q���dڗ�C��i�a����m��湣��v��:�\mvY��W�����NNs&����9�7[:BΙqqp��^{q�����W��33�wv;>.Sp>Ƥ^�mˮƍlsk��Xz��[v(J��g�;�n�<�m;�,5]�xō����\�yf�^�ݧ����iݺR뎂��tY1�,��=�-{:�����1��q�c�#h�;\D�귗�(d�x�#mAk�Â��nݹ�ň�2�zza���4�Ivk��yË�\vj��u��5��j���x�f���G]^q�:��9�F���&����wM(g�wn'nn���nG��;\����M8WqAy�cɋ�x�j�ʧץ��yYk�>Nq���`�1��`���sa�g�8�׌n,��w&[�]�㞬v��-+���m�W��-���m&;wb����bʣ��lۊ�N۲��ԅ�u��]�]�xN���o���x��`�k�u��sMVwi�v��5Sv�66������ms�m-�m���n3x�U烺�]�b`�4v W���v�+��.�9v�d���'���b�� /OL�/\/]R�"��:;� uq�u5� ���\��⇎YzE�AVN�P�q�"q�-��"��j�㴨n�q�j�'=+�v�m�G����ri�Z�\��k=���8�M�6�2��!��jܨ�Y���7O��9���qs��qm�q�n6�ϭ�C��z�ݗX^����v�m<q���t��I�7;ny�J����,o=�cz����;��móS�o;�W�ή��֐������;�;d�Wu)F獡��u��2��ۡJ�nάkǃpn:�C�7]����27RB�I"EˏO��t !���놭��8��T����m��3q�W��Etg��۷k�[�nл]��#�q�iz��y�2�����g�K��v���`[Q�5fzٹ�f�e�c���R鞹��=�:�T�h:�ӵ���G��U�n2�P�n�&;\�r\�7�y89�<r� ���Y7p��g��;��=�b������	\n݊.W��C-�
�v�籷�eveT�=��k��rf�[��>3w7�[;6�ێ�Jt����19�"��Y:.8�g^:�N<�K%&�;��7[p�;�\B4�51���7[Eٺ!.B�=mWc�����wƱ1��k�؍[l.u�!V���:�ܜ0w`һ����Nh����kn��u;��]{!�66vP�8��ƺ7������Ξ����Y:��A�[Fov
�d�y��K��ѧ��:���qj��ve�p�YnM��ʍp�3ںݰlshX�.LI۸Iۆy���k��[�:����#�c�����i�\�4sc]HÄ�Yͷp�G%�rӚ㶝�K�2玳x]���=H�R]�}ne{9��;�3����}���g����v��ԛ.�s�n�;u{=��;v^4L��]�M6����>	N�;hĊ��v86���=n�!��ǖ�8����r������s�`\��)1���r�;c�D�c.O�cx��p��1-ѡ�㔪�ks98w�.!�K��c����zE�xu�lN�9iruu����y��{Q��ێ�؎�U]=r8���EF:㴛�A��Sc��B�Vi�X�(=�٭N�-���Ū�ۢv�x�N5���Q�zy*�8��#:�n�k������+�8'�]��k��t�z�spM�|��^��v�7.���9��6:�n�s�t��c�۵<.���rEq&=n��Rŷv���u�����;i�u=�l�̀|\pݚ^��n��I���#3$7vԃi�dᮆ�V�����T���ť�=��p�v��#s{3ۭ;ͼ�h�g�M��һp���vNq�ۓ��<vΐ�zzb�����@�n��:�t�e^��l]������O�ǁ�1���<tv��97�%�,&&�Gl���6�Ɲ�m�gtAg�2q`;(8�<X���{q�c��t��`h��:���z�7eP:�':�ݱ�[%����Χ^�ݬ!��k۶,cb�t����v�<�����Ư@���.��8{6���=�D��;�L� w]�r�CO<\�/[�Y�qۃ�8����X����Ih�{e���Gc�<mm�\�sո�vݹ�u\[�Q����u��\{r��v��e��:�`|��0QwG�y�G�m�+�K���uvz����`�Hv����n����!sn �K(���э�vu�:�v}۞=%ע��i.�$t�G��:�v94خ���&��{G���(��ky���Q�z��j�����봵��u�i��Y���5�ON�����m���5�5��⍣k��r�=���V+sn�>���@����4V+h�P��$M�v�r���B��-3���1�Ý��#��{c���u���gXB�/( �;mǳ�B�m�⺍�e�a���q�({nE*�u��;��A�M���ۢ�۵m�ۧ���Y�n1��d�6��=m&��Nt���WM�[��O;V6�Q�;�-�^��Su����q���a�ؒ;q���ڱ��Gnv랊;kp�k�GW�����7n$�Cɸ��l�۞�	���(֟v4���)���`7d��R�c��������v�ޮ�\�;4G�cu�a�!h{��'�;fjg�la,�s�g�nE�	1�nknc;s�n��'���[�m��pv&*ګ���e��7;s^89��h����K�� �vG�a�ŕ\v/��u�=�8;O<s���5�ݍmwCv�׃{unE���2y���^NH���(�B�n[v�r��6k�$ꈇ&�]���c][�j�۵����<�)�N޸�뗇H��V�P3��R��q�n5��'���;m�������gx���+��s!ۖ	���%���ά�<׃wb؜nv5[\��[6�5v˷mk6�.�`nu����z�ntV;�^���'���nz��ny��:�L�c97g���!vY��m��\ώ��WT7�x��{F8�.��)y�|��mp}غ6����.�(=��s��`8v^2�Ź=v}��<�����w=�U�E�lq�PwۍvM��� v��v��l/�Wg�^�9M]'��7<i�l���y�E#<����Pt�g/<���O6�V0�����Pn�<�6�V�]���M�FvB:������綹�n�rs�7��6�^`SR�y
�i,����U�S�����z��Q�Ϋ����;@��S�� =uZ�l��ޞCu�z���-=St�ۤ��q�n֝ghs�[�L�j����
���K�Gv��f�n ������+�����i��xZ�[�6V�����u\�9��ZH�q֔wYy��*v�����'�ͭ=��u���˹���հ��Gchn���kh۴������s�)m�ё�g; n�ڋ���v���g	���W'�nu��v�؉��8�:l=���b�]G=�:QD��T(V��,���#�*�"Ҷ���,鵕���H���IE���BIZe&p�8\�[9�(�J,!V�T:�dg*��J\���T��f%a�%"�mN�M�JETJT�YIR*rJ(�H�(:�yÇ(E��2�$'%�H!�,(���3,�E4U"MMa��R�	�Ð�B�)#,.Edn3�KM!4C0�KID���O$�t$Nf�Ea-%1
KP��͙s
��\��R��H����,�J�k"3-B�"QP䨤�4D*T�-
�'���#��(��QtR���b%b�h��0S�͑��6�)��̴���JU5",HY$�W�#I˜�KZi��i����U5�P��a��ZZ�VH"au$9KNt���RB20�\W=�ox���e�c��غRvͭ�s�����h���vŹ���ۇ��7θʌ{u��!����]�}�l����8�.$R��3��iz��x�65Y��Д�WGhCv�}�s�.�]��	��|q�+a����ĩ���_X����S7m�Y�e�������pux��v��sV���W$<�{nwRV�{ZY�ͷ=��t�p��s7\�q�;vynvg<���؍��}�4�rm���::�.�u��=,�uu���G�����WWa�L��7U?������3�2M�l��AnB�cG&w7n�n�k�9���]@4������� �r�y�nκ�L<tky�\\\���;��t����WY,�s��p=����6㭲���ؙw$�	4ذC�kIjy��
�qϜG��Մ��4nS��:;�t�8�K�gxx=�����w�`��#��i� 3���,s������9t�E�-���=:�ӭ7X�f��Է��� h��I���ɦ��\���롍tm��o���/&�ۍֺy^����.��Z���[�]u�N5m��Q����r�Y	M���6���\�_/V�r�Ҽ��v��M�ַT�c9���{lv@2Dܽf�;���n1iw<%�n�N�n����g��ӌ���S����{k�8[�ò�N�^��\J��7;�v�>�[�9��Z���ו{ǀ�g�4�ӷG�w���Y+�.az��u^�v�g�ͮ����|��km�{S�2��gb�y���0�d�%��v�+��,l�n�4^�m����e��hLܩ�۝9}���9�uq8y�o;��A�Υ�W�z���2�ŭ�m��νl׳P�;Q����[~~w]��	z�o ]ͬ`,�	���gǭƷL8�vۀ,���Nr�{�m��g:tӫ3�ˢ krm�x6������۳͌y��ur��[m�ק3ӧQk1�Y{���/cY��۲;{s�x��
���;��!�g�|m�<�;)���^9�;g��9���88c<m�� l"�M�9ܧ'<��w=��0���rnra�{��Cv{c7`6�dw�	��&�Wo;��0q�v6܉���a�3�G�>��q�������8�r�nx3��	��y�M�ϝ��v<�{c�^2a�&�y�a9����ۿ~���a"������A�����b�ȢvMEN���;��;lz�&�\��"'�Mx��ڐMŘ�]��վ�`�v���I�õ��[*�or�@�*2���w��U��&L�	mF�� ��ʒO���T�R��xH7}�OĂN��$խfR"A
	�"��۽̾��l笼�#n��A ��ȠA�����'�C霃����ji���R�[��c�{�I��1�a�	"�O�;y�	� ����sj���<!Ù��#	q��	H�R��s�	��j���X��U��v(������>���D���޶A��=�� �s���"5NT����#S�`�~��c�y���F`
C`�9���|m���{�eU�)�AO��G?gyLW��K_��&OImSf ��JcE,}�.4qo�w)��S��z�����a����2�M��p$�{"�I#v��� �VTڧr���d��IrH�(�H�kƌnВGu^�I��Bb��N(�̻�I ٜʟ�ẀH��;2���I�1Y]θeT��4��h&�s�I�$��o��	���>���U��jG �^�a jŇAбc�v�n^�0o+�K���L��@���l�E��7�F��Փ���wc%��6Ѹܖ4��m�;�:�;�����3��\ㄤ4����}�i+J	W�,�� ��|��E��6v,o�ir��uV�z���:���6F�H�T�(�[X��|I��x�vI$C�l�{{͂A�1��+��:jO�7X1(�0&0�159Մg_u0H"͌���Zc��XJ*=��w���ϬaQpo� `��U�Ԙޣ���7�i �؜$W]N�loVCa˹�ƍ�/Klcʎ�$����^��`��a'�!DD� �1���BɎz�dm�k[$��l�	�8gs�I��B}80�ަ	�w�f��I�1[[=m�A �ʚ��n+6����W͂I���#�DK�\]��޳���L�B�5"��#qa�(m�Gm����vC\J�k����b�[��E���߳�ȅ�aбg�e��=>� =���y��N���x�>=y�A�sp���%&H"��~^C08��?O��Eo~�0�2�I8gr�Ks�=Q;&{]@�!	J�!{u�~`3�BH!�iA7�2�:{:�$���`�ܯI�k%&�L)��:�9�V���ͰIn����A�;�+��ھt������ܞ��e�f2x��޷��ҏ`��s�#�ħ��d��o�Y�ۻ���_^z7����vh}:�)a�׶�Y��Ͻ�2^����I+�B�q࿜�fw��m��)�A��S'Ğ3�R	9�|ߍ�7b �o�a ����vM.��w�Wnd{su��8��7m؞�KP$�F3�(D�
^vꙀ�(�d�@�Vۮ ���I'�6��r<f�ƞ���['��ٞȣV��SA�ȑ@�a�k|�
�9�o�� ��{"�ھl�$���9�~'�(�3	I�I���e�C ���wj�� v�j5�	 �p�d
':��p:dlABQI��47[槯S����|H6w���x�z���M��9�7o.��p��$\vX�$�0&0�1U9�0��u3f�q�xP��ay$%�qD����E�o118����yg���f�pg+6i�0���W�/����3'v��q=i�]����3mB��gbʎ���#�͏���I�����,L��Eن��F�<�7)�Y�#�kn$���)����v�Gn���t���	�l��6hpN�.�ɹ�a�u/6:�۷c�8���,�v�gb\��хL���lv���Cl��;���4���x}��I�u��"=�'Z�-ƺ�J����&����;qv`c���[�n�n�v�v���c�����#n�k8ˮ��F2��/�j�r���̜<��\n��ڸ	^�WZ��I�
�ӑ�7�����ߜ|�r��������<��d�n�z�21�<�v�̜ށ^'�����m�D�#%D�&b�Q�m�zX��V�e�Vv��F�	�"��~o�0waK���hN�0u�-:��dB2$W��ݰ�$�ަ ��TLen�2U����S�$���l�sp��Ʌ$(�Q�<^�'�ei�Cp�Ҝ�A 2���Iu�r� �=�r��H��[�"L�P��BR� M�|�>$�^A�W=�*+��ݍ�O��y�I8u�I����L�'Dנ������ݎ���5c���\׌=���{IƳ����p�$����R��u���}�A�	ů"����1����l�O��y������N�WĄ�S����p�4E�0=5G&��[�"+��+4��e�a��X�\v�y��^�_I�K�:V�ذ�u�dq��4+�VY��]�%M>g�e�sAï*ApC_��h�U�������!�#�w5��$�8���7c�鉿VgWN^o7�A8u�P5tcD�2
���w��.co���˩Cn� �}�^@�Fs�x�}w}{O(���3N�ы5������yk����œyr�D����'ă�^T���|�.v�]�X�*
�����IJBTUB��]u^�=�=�����$���7/%�������Q۴݂8=��0Iï"�$�;��-B�5$:[u|�$�l����)%L����e��~d���wF��+��ǐ+�5�S�|7+��F�:;{{A>98K0��DH�
h=;BH#k�`�<m�f�ȯߞ�i�<H�d@�	�{$�:tʵ>{,�{c�w�n��R$=Jͷ�mk�j�'5ջ�v�n6#EW2�SQm=�Q}1����g@�O����@�{�3(�Q&P��--�U��1�Q 1.���^�I7y��н<wv&�nP�jpGA30� �(�v�#ow�4]v���آ|M�_7�I���1��V�8��H�1	(�)����
��^�N�:�]��km�-ˉc�\no\e����\��&f"(3WI$���I>����+����b��T�>����H�#DB2�bB$Vξa��[��.M	��oa�I mm�~ ��7�f5����	w�$\fX�$��D�H�l��S���I&5Gu�d�ʮ���Ē�/[�@���� �%Z3�2`4zv��*�&n� Ի��&�7��O� ���[^�t�w3��Z��D�K*�.��X�}Q׶toh빝��"E�Ō9�PQ� �!�9aΩ��H+M�����ީ4�8b�iR}��3+sY�8��z��>O�&e*$�%�=m�|x��	�SU8hY&L��S$�33y��=yR4�7����1�g��F�4�I-j�"�]��� ��ux������T���un�]���߼�B��"G���;��LI8z�(����N}�9-�l�osy���(\$��L�P��� ��5q0�t��/p2	�gsd�A�ו� �����y�JsP����>�<D	@�1!(t���'��P�	#&�ʈ���9N�3;�$�;yRC�����I�L��n�����N��r2l������ �qe�P�|�n�F8h#�h����nB��aDJ�"&��� ��x�yW	�+wSqn)׉#7�`���^$f���U�Nw�D)�Ը��ݼ�ŝ��qQ��;��n�@F����'��)���'��x�.��=�=(���'<��Y.FO��_����^�>�ٹ�)��ۣ�n��ߑ���7c��Y��p펤���qY��n}a�[R�>�li��ꗺ�i�ƫh+r2�]�s���p�&v��8v���t8�.fx��{<�w;�9][8��b�GFv�R�T\j{��ӻ�h�,h8S���I=na�c�`x��ݎ��b1�Jt]�1�r1r�Fݭ��ۛ`�]6���
�c���n@�ll�Şvq��5'm�wn�)���;4�^as�t۞��c�߿?�>�c�úX��d� �t��	$�s]�gWNmѻ��-%��V�$�p��	 �؅�����H����ՙ�(cKcY;t�z���N��� ��|�&�楽6�M��#$�*
������ENc�l�|bg{]#bs0�O��D��|��pqn�1�W�r�K�v��'	0r�$���)�M�oQ/v�ԕ9��z�UT%e_)RL�(I0%~-�sdss���-�^��0f���� �>w͒	����˾͙�$\�A�8�o>]s��x#Q�Vf��X��8�n�V�%��݁���h�L)�3"D���I ���$����2�A��fLĶx��H ��|�`[�ZF��#�R�~O�=�Y�\��M��	oǍ�O�����l�K|Us�p�?g���+�vo�����*�&������Y�TX������43k�^o���N�_6I gn�d�4^�Ǔ"��ߤ���G	S!)	D�;:� �'�sw��I񬳱���먰I.���O�;w�fn�J�L�QC�<�y{�����M[v�'sw���I��fFӇ��H~s]X�0#'A��(�f%F��Vx��p�\a��hM;�"��[$���oĒp�]N��(L���m���]ϥk���{��,sV���F�D�S����@�BB���SL�aL��._s� ������]Yv%S1���&�T���cdof�h�B}0�D�����A�}{�Z�^��l?��lH8z� ARqg���')�ɘF
�&L��nzz� ��+*H$n�co��?��w/U����ķ�Ճ[���}������z]k���Ǔ��S�k���3�^��p��W�����V��Z��b�=�^�.�f��]9q�z�x��4�X��4�͡w���͚O\a�6�(�S ��˜��(����Vɗ��ɹ̝���1�K�G��7r�'=*���}��^�<��)�����u���D�0~��:���^{:����V�{~��^/��{)�;�O&��f�ѹ����a�K'o�Y�M�!���"6�qm�z�����};/[]�=?2���B��9q��Y�AV"��(�������M@ZU�-M���{�F�ώ�p�ʽ�xq�z�&c�e.���N���	�mj�d��y�_p�{���}�ۓ��F\��'�lV=x�V~L ����Q�]%޼����S�(�&�c�6��,���]���d����bt��+��Ujpụd�<�U����߭���C�J�7s�l�-��ݝY�;�37��c�/w���v,�X�^��l{�uZ�~�铆^[�%�y ���s�FC�L��\��B�����#y��6����.�ͯ���p��P�$ҹS�-�Ѱv+.n/u:�\{&͸��z#*��R��#���{��9������!�a�{���@$�G��M�?Cr��/@^'�a�� q����WgG���-^�dn*<��>M�g<�'qw^��sA��;�n��ɼ�?q��:�����V!�"�*f�XA�@"O�,���MAS>���F�*r����\K���QQ��Ҭ��;�gO^*3C%�fejJr$P�j&�x¼akB�e^&k�� ��YyJ#78p95N�(����eRȬR,�Y̋
�Z�p��$�AeW*\�8Dٖ�+%21B@��H�T#T�&F���e&����QJTIQ�3KiT�j(����K�U/9p�J���"�Idl�8q��j�i&a,",,(D�$	�I�TR�0�3��CM	S��R�Z#5�Er�(����F��rښ"YU1+�$��ͬ�Q�QXWF���U�����bZQ""��ʈ�
�,B�J�,Sj��3,C��*�.�3eiYV�L�j�t��K�+P�C�)eO�)k��ē��͂A>VEx�`��3��1�y���7��m�~*�|�f�k�x2?�� 7{��r�� nuk`��n�J��fd�l�y�$r���<.�ј����Gv�l�l�d
'+��38�z\�L�R94TE(#"7Gm�G�׳��L.�!���k���.w���`��J"��S�9�z�'�a���H'�]|�4�'�f�s�.�R�{ӷ\O�6z�):�Sg��(HLR����:��eL]�Pd�}k�#Օ���;��=6l��V����c��H�Ef��lf�>#k��Fh�3}2��s�5��Wy`/~�[v3�F��:���7���׻�+h��H8gr�ܦH&�;�Ű�h���:���P8���b螞~�e�ԧ�����m�#J�R���ض��{5��
M ��\���2��(8?` �#@���b(�Df�5b��~g������Q����1�*��$ᕛ��	�ͪ6(�Y�%�����w�v;6�����c=�x�ʗ=\ \�UuuW"e��|�\?z.*5����*H$��l�����4��5�i�@�,��$�y����ɝ��"A)��>l�jOi%�U��ڒH�]x߉���lj�`�yɻ�o����IY[�fd������ߋ���>$��u	���LE�?	����E�wPV�A'�*dB��sƏN�$��P�{���A$�/��$x[3vs�mUU�t��
�b����'�<�EO���q�L�F�w6	� ��#�,�zw!\S�R��(s��kX%�;�L�2�V���nb"_�M������GN��� ?E_�~�?I3�U���W��� o�IS ̣Q ��͸�삯f�ۓ��%A�y�7��C���0sm�X�9���cKZ\��uģ]����[��-ӧ�v��8�9��u�� ��&7V��"][59��Ź�
eJ㇎u��^rk)�킻����lw/h)�V�ѭP񴽴��j�nx7d�塓���I�[60v'�1��c���}�i��`�-ۮ0��u;�7��6��ݹ�ɗ�n�>Žm�y���yه�)��w6;'\�wg��D�T��㻯)�@;{�L�|	<�+;���ٳo*k��$6���1��1�L���2%Kg�nP�cH�S�|�Z[��$�E��6}��<�G��j{����	U�PD`��}�i�d�㇞T�n�Wa�f��ݭp�+	'�{��'ĝ<�Y�f$�����L�/�9�D�Ɂ]�*[t��$��@SޫP5J���|�����4�Fv/�Ԁ+���������Y�Ȋ��WO��$qא+������.��ڵo$&� g�2��;��S�x���!�ZS��X�n��v�u��З�m�\_ϘWl�0TJ*T�/�_[~$�yR|FSަ�V��)EX2���g�P�!U��LLTAR&�ܮ���R7�w�R.������q������[�ٻ���ʞ��x��Ԝ���z����*ux����W�=@�����m|$�˞E H�?�lpr�;��Fjo�=�� ��p����ܡ$NS�a�I�%�u��s��	$��(���̀O�OJ��(�J"}�[��W6L�$'�jO� ���$���u��P��U���$�9�$.��3HD�BBl:�/{��uU����D�J�b�'κ�|n��qki~{��nu�F#�n�������{mn����lh7&�i�����ls�ϟO�G	��%H*D��� �r���I���̓sQ<����s��So��H���ɺe^�	I�e�ۍ�~�:���vLH�f��o���GU�6H7y�L��?S���-��<��1$Iѻ��]�s�0ωow��H<2�6{ob���s6�=r�X޾;���c�;<5{"���79���z�$������*����&�\!G&z������78o5���$_���`|OW^�����2r�A��-:ND.��z%�*%��a{n�A}��$A�ՙW�2�1w�,��y�d�MJ��Bh�,���O���#�ں"��<��>��~�����H��~���oP��G�^>GW=�y�(�#%8�4w	ɨ�q��I�w<y�ݏk�f*O^�ma`�-�Q�紎�*A��ϢT�%!%	���]���a��d����ݞ{���(��~Hd ��ߓ�����/�D���������<w�i0�}����g�z&�G�?>�n=u���;q��Z����QDG�������P���{?;�ht�	 _�}���ap{�pL�����1}�����/�q��C�kÎ�_]���%&Q�f�=OD�����g����u����ϝ�ݡd�ap��=��}�����~���=q8�����߻<M�Bv�Nӑ�]��$�FY\������(�!��h��A��{�Ҿ���#��<������bl����w���@D @�o�>�}�unD�#p���:���{�B��9��Տ���g[{��=�bq�Ӗ��7���嗍UM{f�� �׏��_�n�~�D�mܻ���>q���~���i	�>��z�\{��!�&T(�`��<	����� ���|7_�`�Ͻ���םw��7�����߿|=@�$���3�w��x<�0�>���x��8'��|��ߟ}������<�n5m��x��VgUQ����u�)�q�W��Gl�w�����3�FX{}��������g��:i0�.����۴$�aq?y���0������������c�߄��߾�z�]�t���~w���s�~}�W]J�:Ꞌ�����:�������1���}�>\O߹��w���?�<L?���1������@�@�	�w�]��&<���/�_6>��E��wCH�>WI����Kt7��0������v��HN>�����s�v�HI�}���������˟��~@�$���f]���;�
x#��mx3g�"�;9$(*T�ELC�@>��26��ǌ��>� i�giӴ�y����L(I������z���qgi?������n�y��?���??y��=v�:L/.����d����N��79]�x	8�������� �Dx ��{��������Wt����pM�>���'��$ N���|���i0�}���g�zdӇ����㺽�!K�b��͉�~נ��2t��ef��"��u�q��t��](k�K��_�#����޾~s�^	g?��;����a���nUm�`-�g�ڻtn]�)�G��g�E��9;`�o[��!c=��Wtś\y�ٱ;ѧ�m֐�v
㪃�l	�Ƙei'l����`z�]@y[l�8�qq�v��z��،^<e�1���[�-�=q^�[i�d�^��j���C�¢v�79�m���{]���ۚ�w0b��v�V���`q�����7_��b�nWu��{84r���Ӎ�~;�]�XW^���	pkr���usn�<ރ;�������g/=%�Ow���q?/���<v�BL.>w����s�>�ȏ@>���#���ך�(�}��˃�]���wh����}��=}pMϏ]���\���p�y�O�{��P�,�� ����Y��1����q��Ͻ��ݡ&��ӏ��~��<q�0���߾}���oD'ht����{���}W��-N�^�D �M�D��IF"Q2/P=Iǽ{��x���Ɋ�����ݞXC� ��#��ṛܞ=�����,@�@�'�����=L.�;HY��>���A4��s�������:���n<q>]~��s�;�~��_�r��_1����>|��w�Ӥ$�|����������]���9����w���7���>������pM����}�\n�������ow�����t;I�����@����*>���� YGǟ���8�8�C�4'ϟ>���7��:v�?��w���}�������s�w[�ڥAp�UP�bUU*'�Q*U#�����QK=���Wn������[��k������tݲe�?�|���a������>}���1DbL-����`�<$z�������_�;���;���x�ӡ�BC�ϟ�vz����;�����뜹:�ט�Ǡ�#�oh|(�"#�Y�W1O��r��iQ�w�O�!�}�g�C�L��O�> �'�jaѣ%Z���wp}�+��x{�P�z�`�����?:�����l�:q�^���<v�:L(?|��<@�'�g�����xwR	��"o銩�R�c|#�^x ��3]*$�FD�����$2=���"�	��N������nЄ�M8��?}��<{���>8��8�B|�����S{���Ӵ�����N�(�Ϣf$�R��eŐ������(��UTn���
#�������10�����y�� N?����x�������:���>� />�ޡhz�qs��q��q���c�g��߽��;MI����|���v�����u�^������$�{��������L/˿�;��a�1E���~��=}�����(k��	W�`�����eIK���d�'�v�bi-q��۞���nZ!�n�c���s��=q�n�~��~M����vz�S�i�w��g�ݡ	�$ӈ����c���y���?~�>���1��λ���av��0���|�o��{��'�t7+��(�#����x3�,�<7������P�c�A��l!���#����� I N�������z;I���_�u�}��.1���|Kȃ����\�q��z���������i�$�Bq󿟾v{���@����H��!�ƽR&�九��G�C���$������J-$����7oǢ�B�m��U�b��L>4xZ��_��w���P?�8&L/ۿ�;��q��U�������������O	��p���$0G��>�dj���|K�q54�i�޻O����<�ݡ	�$ӏ��}��g�ς>��v���7r�u��S�N�_��w��v�c�~��uΔns�u�ׇ��ǜ�������&$��}�G���m��s#��������c��߾y���Yq���;ǎ�;N��$?��}���aq����޽���?���v�-���9X�F��κ-�	��xt�ytA΃��t=~���q�u��Ά�o�����|���a��HI�	�������v�H�}����RpwП:<�~s���&���w��q�ъŏ՝��f���b�:PB�2���Y 8����#�#��7��I�{/�=��۴$�aqw����0�ނ3;��dz���#�*������ͪ���t��z_��Ά�s�����I�ߟ�v�����>�������>ݓl��_Vgڵ��H�$` u��~���z��߾���D�>�� �$��P�	�/�υ�ym�U�Ho΂aeF�#�@Dy>��v{��a@��#��￼=@�	&	�qW�^�ӂ�|B;l��+:��L�����r\&˟��\o�eK��RZn��YY���+��� ��#�n��7;�&F���ꞃ[[�y����n�?�?y�;ǩ���w����=s�/0)�o�|��vz���;N������!���}���|C���>{��z���q$�}����g����t�_��;�̝�>w������I���w���g�-c��j��	�,m��T�r�M� $��r<�!q뿟���ƞ�gs���� ~�8�~��=}pL������ݞ{�Ę[�������C��S��LrV�@}^"����g�}�u��,����vz��iŻ����ӭǮt7Cy���������HI�~����~�K�f���s�t0Y��� H�����S��pY����;���0+�x)�ϟמ��xY�7��B�u�OE˞`�=M�_�vz��N��#�#�^�`��@Dy�O�E��nm�����?c���0��?~��������0���>w���u��c�[���s���!��(��eD(���$xr@y�����{�13�~�}���̀��'������������Q#=�}`�HB�����=N/�{��?�����s��O^c�������|v�SB��~�`�ϼ��0�_fz�$ �O׬Y z�����{�&#c矿mxY�� �ۜ��Sm�L�$����^�N���H�~<�����Oތ+z���{|F7sW��6�@=Ov�|�Y����:�#Jl�I�B-��tՖ�L�X����E���N"n�C��7Xw�ڋ��t-*_N�1��~	�B��Ό���JJq��J~�f��h���1� ���3C�o�J7c��D�OI�oG�]yu<y����\����`��\y�ջr���9.Ơ+;(˷��������Ν�$G75g.j�8bG~�������,ч�.���2��+��O�ͧ�O5������j��ukQ���Q7m��U�[bya�Y�U����>�a������g Ɍ&���@���
���D��:��[����2����<��;������,	7z��ל�����8�����\�v)K[��70������_�'�Z��Y9x�5Ox��]c����V{�գ}zz��}�D�"���f�<�˛O<�L����u��w��Â�9�0���E�#ڻ��]=ko����aڻ&�<v�Z��:*;aӾdᓋ̜��#L�KFЅI�w��D��]=cBy�r�ߟ��bx�j=���I�k��9y
�7��f��϶K͗�*P�4Zf�b��ڜ]b UA���1'~��;�6�C��|w8zB}���J�n���}fVy��^��Fq߆�7�-�.�����y����o\�.v�wv�ZbV��Jf�e��2%Y!! ��$�̪e���5#���Q��e��a�@�Q2.��0P�J���*������FKB".�9r�T ��2NV��4�D�C�$fY%�\������%d�¯QsU#�m�29���E(�JEMUFVI(�vU�$dJ��ja��d-U�и�s+�\�f�em5(,���A�"��A���QK(39T]9JtBH�"$ԱQ9��;)@��Q"��S
�L.$RTDq4B�����A���qFp����5%,�,"�P�KJ*8�v�PjY+B��Y���5�[2��-�b�eh�QRB�Z�R��ZXZ
���*�U.6�1I2�,-j[)L��bΈ�Nu6&VX�r̶�P��*�T��d*�t�#E����V�A�b���������pZzPʹ��s�+�Z�� �h�;q��7�ۧ���k�J烜���+�G��,���9�\�燝�<7[�-����nѳ��n]�m�3ˌs���e�	Iږ�ud�3��Rv,oK�ͮa���^6k��ܦ�:��mb�x�wnu�79�g9�qɻ;l�����.1��m��F�ח��赸x��v��/�v�ܪ��z�أ׷c�v�S��γp�����Y���k�pf�BvU��яe}�������'�p�=��!�t�6+rX^Hf7��ln�s�4+e;[�6���#`FkA\<V��,��ӱ��%�B|\��E�,��7�ݼ��+���c0C�m������R�Wl����)�71�&+�����َI�m<��Wۋ�$�D͹k���n��sxypi��v�f�xS�d�v8��<g/���vap��΅6��l�ݜ�ǎ�d#��okud.���wn0Y�s>.����ݪl��u����]���/'lr�����R귰���8�U��}�����S�%��e�GO� G�S��ݳ��Ap�,��B����v��j�;�y�n˲�ݰ��n���z�D"�s���s��r�����l^�g��"�����	\�m�0&�Y�����\e��7�q%�� ��VV����>��f�I��u�]n�q;]��ǜ�y��;b��"�k�5�^�s��Ѭub��m׶�-��ORܽn�ꅭY⹑��Ҥ��s�oj�r����;]�v��[���n��
�1�p)wE���]x�5m��ո�e�D��y���܉�:�3��x싰;1�������w7p��s;X3�%���{���t�S�Z�t��Ў�:���2n�m��m�x�3֭Zt�8ݱ<v^ۮ�l�������8Pz�.N�͵�[לط'9�l�mq��b�+ё�����ڳ�nu�N��U����$ҕ�fE������5ute��{����0�ݿ6�bP��Y�u����R�:��C�dv��덶ذ'+{c�m�b���F��Υ'Y.%�CnB�u�K�bTƻumۢ-՚�G�X���,���o+���6֌03�鸠��p������ZGU�����L�r8���Gwe�i�t��]���9��Ξz�=�oW�7kv ����~~_�dp�e�9����ɭ�p׬�b��I�4��L�uWn�w�yd�MbԎ�s���������=��y��Ow({�;<O��'Fv������t�P�4��|�8�8�w���O������t�������orav�?o������虁>*
��)1dx�Q���π@�<���2�������Pv��&�	���=���
x�:矿|�#��Y�����*l3��Z�hz�\}:����Ӡ�\�n�;q��|����&�	4���߾w��t�!�N��c��L��C�A:���pL��������Qc矿|���&:?���8qz�t\��S��ﲅ��V�i��H�G���GU߽�ݡd�&�G���|����G�#Ȍ���G�#��v��K�>�$������ s��?�����+����������>�������ݞzF.~���3������ ��?$< I N���~w�]�v�gif�� X#��F�r+V�I��tnSzn;t�����2ON�q��Vً��'QD���a�����O�E=�sE������O��ߝ����N>y����Gz��
�����P=I�߽y�����n	���w���F*��>���=}��_%3	)&b`@O�#��P�<	��ymP�ϾT>ˑ.ʻ�,"M}1Wl�)��/�����;ͫU�&��6N�kR�{�]߉^r1?���N��vft��Ѯxq���+T�]A��� =�o��y{��g�v�M!&�y���x��q8�I�?�|��=M���������7�qmU{�E���&`O��κz�P=Iǝ}���<L)�h�����IQ��{0eq�qy�%>H����;Ǯ�;N��BC�ϟvz���u���㠺�Cpo<(�3��[�"���U����#����N;�߿ݞ�z�P!$��������|(�϶�٨o��yQ�~���1�<����z���������r�ys� y����x�$���围��D����s�a��|??y�\z�qaĚO�>���0�z�}�|�,�k�dQ u	��i��7_B�$�gNݺ�ʯg�.�r�����y�{i�iy��:�K�qI�G�u�������]\�r�?�~�8������������~}��縌PF&pLs���0t� I���?���>�n��߯�;q�_�~w�
aC�>|���g����w�8�:z�9��::�&��;� "=�m��썬���x>n���w�ӤI��vx��I0�Qşmx)�C�q6��k�6�~��k�&exa�P2�)R��f&�<�o����g��޻N�i�~���hY4��p�}�~�����>�s�?���e����V�s��W��g�C�/�2��L����{+RK��ڧ�X�ź�t\á�/� �}����q8�I��������oD$���s>�������&`J!D(�2�@G�����Z�>�sl�����~vy�b�8&�߾w���H�O����z��~��~��������}�����ù���G��ݘ�&���}m���������;s��<�����eĐ/�;��������;���hx��K�~�g��|'s����q`\��9�AA�A"T����s��jF��ɝ��n�ܝy�ܕ���߉��K���z��}�����$��;O��:��	�!4�������N?�����?{����Sv'?w���S{���:~|���'�<���3�G\�����aq�]�#���T8�#ۘ �����!�Q�����ΰv� I��?~��<w�Ӡv���غ�+��ן�vx��ӈ�ߟ�������8��G^c����߽�ǉ�$�!8���Ώx�: � D�geL∕�|�~@B>	�?������`����c���p�߬����W��o���������3�hO�����!�y��BM8�|��x�\x�@�����g��j�08ͱ����̅U'�S.���{p�ȅ
��7�{N'��������kD	�N<�n��	ƃ���]>���w���1�����Ν���}��������:��<�:뫪��0����ރ�|L)������g������������~|�bzpO����I������:�n�;N��!���vz��4��Z�l|�M���&&T JS�)�X�zR\�v뷓[U��tËks����}���s�87�v���|�}��q�aMd'>���;v�t�	 _?�����0�;�����8>f^~�����^����>�:PH�� ���o~�������Gi���������o��;?;v�P�N>���v�\x8�7�~�������>����u���ƾ�W��������N�-�:����tu�S�7G�h$��������&-@}����g���0���u翹�����߽��������%�'I���c�x;N��!��|�����G޻���K�W9��:%�Y���4����#�@DyN?�����x�S
��|����Ng3�~�����{�)�����X���1s���ǝ7K�:����>~��0���:�������n���������|���ަ�|��x�ǎ'8�B|�����S{���N��������	ʸv ����%�L?e*��&k*䖙�ju-����5Zq�����el�_M��F7�@Y�sf�4�L�@�p�:�c�����;�F�K/��3M	������+ep+	S)B
^��X������{8�q��۞q9:ǂ��t�:�O=��]�ӷmm<E�
��7V��>�'='8K���#w-� �Փ3��9q��웲��fm��;g=�v'ڸ۸���7�rb�n�g�l��06ֵ#voc68��]O;�����5m��eݶ�ن���w�qj[nzہ��7 ��P5�{=9�{Dv�q�m��e�r��=��mECm�pk;:��A.�z�;/;\������Wa�]ur����IǞ�}�<ώd����ݞzF*13�o�{��&翫�D� i������dx�}�@v�ݞ!�i�^|>k��:�:�y��x����$x<���<en'�>����P!$���>�z�蓂g(�����!�W��Y�\�?��?O�?3�m������qN�ˡ��0z��������S�	Ӵ�_���;<v�M!&�y����Ͽ�u�}����<���}�'8�I��ߟ{=M���i��{�����ξg��u�s�����>�d��ew�d|$��rߏ��Q	 ��{<�1Q���_���I�<@�x��|�s��A�"+��{�"<	 fK����#ནY>L�DA
$O��Ǯ'�������i�$Є����$0|ϽKJ��a�ߙ�i h!o�]=I�3���������3�|~>��E������_a�y�N�a6z���Z۱���Yx�i�[�.�tB�L��=�IR%D̒����G������'NӬ�?/�~�xݡ	�$ӈ����x�Ǚ����u����?|����S}�����7�	0������I :��bfA�D(���X� ��w�Hş �(�
�Ι�"d?��ݫs4��_ٙD|���6�ͣג��YMQhW�y�6�|.{@��H�;+��\h;3�q���r�^A�$=�=� ?�?�߾�<���L�������t� I N������<w����C��	��YT�@�O�G�> ��y`�'��y���n<q>_;��x��a|;����y" @����}?t��>u�P?���g����x<�0�1V?����<L/�g���뜺\�Ȳ=|��`���ӊU� >>�}��;Oۿvx;v��BN ���׃#��| oݿPdze���ݦ:{��v���0�^|���'hם}?]G::���ô����}�?�dvn�A�C�W/��Z!oI�G�9����0t�S�@�'���:ǎ�v�>�  @�����,�|W�J��}w��t<iNGE�mu����U�Gn�n���d�u��u�k����O���ן��������x��~_>v8�4���|���G��� I ~���g������{������:����g��>w����bq���c�������Λ���u���S��{����S�t;N��;����i�|���;v��BM8���~w�x8�
i?�v�B������'����@�V�bX�_,����{�� S?gD̃(�Q31�dԜy�߽��d�@~���g�����|;���;�k�o�ƧX���<�ޓ�ݯM�TuÓuO� ��&g�z��'����C�;{nU���uQ�ȥ�g������H�%�'I����X��;I�!�����g�{�N��5�ts��Wx�ǎ'�w��j���h���=$G� #�y����
$�������=I�f|�Gϫ�egt�Q]��C� �/�?u�n�����]q�y�y���7��{���z�:v�;O��ݡ��q��UG��=d�>~��<	�gi>}����ޡ;N��O�����u	!������NB��I�&H&jdDV{;���zDs�.�$���uq������S����~��i�뮫�.��i�ǟ|��v��Ɋ�������=���s���`�<@�U�{�ٙ�� a�3�O�>g�G��!������aq�>��<�t�s���G^c��'����a��Bo~��s�e��Mf�|7�$a�>� �!���>�z��N2a�?�w�ø�F#���Ͽ��'��]���Âb���ǝ7GW:를���o����g��:v������x:L(x�qu������\�8�8�N$�{���ݞ�o];C�q<���@�7��̃(�Q31�dd#���#��[��>,�R����2b�>�����=#�Ę[�<���	!�#��"3�|�}��|�:~q�����_�g 0����\���8Vvg�[7��p�Z�Yg&������^�o.u@��r)*52n�S���� ��3�������g�{�N ������us���^c�'˯������$Є����Ώx����燗~n u�@�?~�������2a~^|��q�ъ�?�~��<L+���~��輪s��:�8qv6hu�cv�im��.�$�$�۪��g�c�����Q

`�1����:�ӧi�y���nГHI����G�>�}r\
���c��#�G��ݞ��	�;N���߻��;@��뮸=s����G�i����{��	���e��(� V�ehx$��( �������:O$�	�O￾u����C�o��^wu���z�����4����������s��y�\z�~�>v8�5�$�Bq���Ώx��
wr���ҝ���@B>|]�~��q�ъ�~��<L+�?<1%H�2J� H��ϨY.;��Ի����y���|v�;O������HI����v���Ě��vz���y>s����|/߁v���?�w��s���뮇��s�u�Og�'���A����1���߻<�_�u����[f8x@�iS��G�'��O�|�&y��������G��׎�!	*�l9�|+!˨����G�e������7�Hkm�}Y��fw�˂6y��\�	TF�S�9m=@�����*��y���3�I/�g�}�}�ߟ68�����F�;��Wn9P�\��¯�Γ�ДGG�\G�^n����m5��b�'r�kS�ݠ��W��h��+�+�^]�{i����I��o�8����q�n�`�:��wI�n3���.m�K��H�8����[��v`�zy�ᣎ��k���n��ցDր�t������;n1�UZD��j:��dKjی-h'h�9ն�fKs�v�p\Fq>��e:8sb8̃\���t����N�S�������{��u�����n?��|����x8�4���|���X�������������||;h����������G�׀~�<1V>~��<|pM�=���s��7\zs�`�={���ݞ���i�{Ϟ={��߿��;<�����۴!4�&�G�~w�x8�
hO�?}���oA	�ϑ���y�~�[�?)u^��� �sc�O�u��]�y��}���A���Ɉ�>����g��(�L8'�����B�5����ͳ�ϼ�� ��'��~��;w���P��}����=M8��N�I3 ��5�υ��#�w(�S���\���:^�~��ɼBM!8�Ϟty��:@�H�?�~���'��EU�W�H�j��y��S�CG����X���c����t~x���뮖��	�y���S�t;N��_��~���̀�A쿚}W��@�<����^��q&�}���ݞ��	�t����׀� O����[J�($D�1U�\t�]��E�2�UKE�9Љ/3q�t�K��~����]\�<�s���@���}���v�S
�~�������6�w��;OF�lHέ��>`��v|�>�>N���?}���aq����{Ǡ��E��;q�8�ο}�i�BM���>{u��=)B_O�i�Èo*�� �֟.��3���P{��`�����p!����&�fi�-y<+�>�p_d޽��`�q��z?���HH�����P=pC8&_��w��#��<
]�V��L-���2|4�����TDA	J�aDW�dY�ﶅ�`��;N��/�>|�hx�BM8�U���1�0���O����>]��U�A$k�*��TX�3b&LA�"G��혐D
꾜b粙 �=ɠI n�R��Q��5���,�	&b"&��וD�o/����E+
��˶�$���E Om�Q�kf62����(K�����L�e�ݎ|Q��b�%��6�M��mt�V+X��?�~w��d)1 ��uo�H��B����U�����HVЭ�m��A�(
)�ꙑ1 ���	��uz��Y[K����V���H���kĀH�^3j��~;�$w� T?}Y�RN_-�03���� �v�/�V]��wl}aO_���z�t����g��j���K�7��*�w��Jv=-��/��%Qۉ��h�<þ��>��v7g�*����e��{pγrn:���vIZ�N/E�a�x��+8�z�i@Z�:������a}��xAy_K��ٹ�c�s�J�˻0��>�5�Y���t��=�tq<�u�<��Bأ�V��LN�7a=��ժ�����*���r��<i5���}��?0��z�v������d�[y�ӗ�7��6
��U/�ӧ��-#�B]��V�m� �L�{�A�C*jk~�h��K����S@�� ��������
y6��]�ZG�eo�
S��g:&��d�{���hZ�q�\�l��g)���,��il��{wr����w��<%�t֭�2�Km��i�^��}�{�[7��أ-�{�- Y��[�!|�-®<ĲC��G���'�Yp�����j֠�ӗWO�%wqɾ��ڑ��y�q�)���J�/�Z6�hpڽ�9����{p+�������{�/����nʲ��[�g���Ak����N]ñ�𸏃��3ᚺ{��3n<���Ι֍������qYֺ�so��x_Mr%�/�.��O/Foud&&hD2�{t!J�l�ry�����Ў��R=�y��v��H�J=���j��h��n׬�z3���w\\}̥����g*fl�w��+8�\x���V��{����OSzȹ{v��@E�W::o���޺��?�ʫD*u�u��D�sYD��i+#H�0��3F���8\QE�r��Ɉ�2M-Q4�L*T��$r����B9&(QIheRDPs�EF)I�*� ŗ)�W"��榬���I8�ZyH�� �L�	��
$� �fҨ
�SQdx�故�FX�R�*� ��TF�IL�EJ��'*�I&�L8f�"ӚШ�Iu4�9fb�̮a)r�hD��.!��*�J�"��&au�j�	�K�`��\ �U¤��r����HTU����
�*J�AI"��h�ˡ��Њ��*P����EhTs��\��&D�*�2�i���
F%9ETU%VHr��D$)� ��*(�f� ����l�r�M�F��rr*.sA
���E��i"L����r�&է5$���������DEAQI�1��(I8Ar
�X�]8�qQ���"�:�x�
r?�6�y�{���A�(P ;w>oŌ�Ң#Ќ�FE?��廠�1��i\��w�$�y���>&���8��ٸ��@E�u}�8<�-µ �iX�{���d���z��."M�P^"�vk�����l��?>ρ<W�5� w4 sŜ8�"}z�y���⫦��旛��a�w����0�����<$ʈP ��;�^��^m���H&��6P�{'j3�c��t�Eu:	=ۚ� �{����[�V�)��t����1j��l��ΦH'ׯ��Iɫ����\d�(���0���	��y��$�>�d�|b����<�Z]S��w�9�k�a����2��S@Q��{L	�����	3�V�3�d�c���Bo����O���׆��q������,n��{�όu���MEp�;�]Y��9���l�J��qI+n��~���x��Y��K/B�qw3ؓ�ٙ�}�}�����O�oiQ�D̓
!����$��yT�y����ۛLz��� N�ʛO,P���h�wp�stb8��.܎��^^��z�']�6�\��m��ܗv�[�[�=����{���f��t�ײ{n�A�E[������ ��;bvM��"TD�l7�BD3�J؍�S0o���n�r��$7]R	��j�}[�N�6�>1*�
D�LH(WN�lH�T��q��;�"�YO0E�v6H$ٺ�&���̥� L�@��[�;�{��M>��'�k��A�u�D�6���͑��ov��=M�I�w��J�2`�4h��	$�ۻ�=%�J�����u9pO�o~'����j}׽�5��L͋�Gm'��cw�2�Q���	�����sےذ�*\'S;S[��si��W�J�Dj�����2�Vܨ�w�T&�j[�x���=�~�����]�t�:x4򻁃ۃqu��œ&\ͳ˼u��hs'���9�ї���q�$'0[y����]���0]m�g;���,n�3�A��r 6�kk�l�b4���7c��^u��m��ה^�"ql��:냚����=�\��ٌݻu6���b�9is��z��v��	�vټrk����x���8֋���8��Fm�c4;�Oi�!^��/�,#��8�:nӨ�#�,q�WqشrW�~��*���\���^[d��6�&����`�df{��2oL��� |2�[��~Ea�SD��l2ZN�-��uor���`�}�["����'�1�7��\Q//t@��p�}*a@��d�F�]z��^ok`��y5[n��A���:��]^�A>y�߉1*�
D���V�<y��9�27
��:�l�P��|s������Z%�}�
��p�>Nr����2����l��͒M����VR�W�gN I���d�����8��.��]ȿS�����%n�4�� �=#�h�De�u�v����p���ks������z5�%)�Et�
$�wwu�N�졻��͑~��@���l/�J��B&D�Q������7�,f�m��d�ҭ�V1�b����\.���W?yfM�aS��F�oY��5^����[�/�����%i�
�j�k���������׿z�g�m0Iߟe2A�����b�Wt�T�3&�Rģ#:)��A���~$�"�.FTy��;�	�.���	{�(:��$LLTL��#om�c:8�ܷ�P���w;B� �ne	"�덍�¬q�7ُ��W6�P��R&L�B��[~$�2�I�>�u�������L���`�E���26��y���k���'a���z��k�虞�pk;S�#�ג��T�H�T�V�v&��E1AJs���a�I����n寮j��'`�ۢ�VTֶ ���lA�9dB�>R$I�f�����p"��fG<�d�w/q�|Iw�(]y��uoQ鞶KݥDG�2L(����� ��F��I�>ڡ�T�T�}�a:�5q��'��NX}^���6�w���|9qG���.Z!��W���y�� sq�VI�����<��-���}���[��Q5N�ʉ�L�1(��vx��j^��'` �o<0�˾�=۝���0���s�Q��dɉQ2[:w.���r�y��q'�|���$�.�}������B�4t�����8�풅���̇`2���PtԶ��D���{c:�
D���s��l�{BI>'�;[1���9�����~<�C�����V�ZQ���o{�><�+;��U�����EN�v�D�Jµ#7z�0nY�O��	��� 0_���������Wz
=ST�O}�H���/�J��L2L(��U��q�, ��f�H$���l�	���B�V�U�D�	"���Y}�f��G+�S�Wq�1Kn:���-����DDqYF������b�b��[�	��v�L�fa��2w���{�|F{RMV��&TL�dLD���t�#s>�f3{:Vd*�4�6c�W�%�n��Nnv6qULQL���H �D"EHnߜ���m�=��z�fI]�v.�p�[�8�������2bDTL���<�I'�/{[ �E�v1�ՙ;{���td㪐|s;v���FȘ3&D!C+:���j�*�5�$��ۭ�E�v7�|B�[uF��Q?nw������5iX�D-!d15���}���� �Utj抭�H={�L|H����9�S'�D�0�׍��2�W����O Q]��2H$n��`�I��'=�U��$fK���Ң L�
"����:^d_(�KځC�;�A�����z�l���;����wʨd���ߺ����&��x�=������k�9��y�o��_�(���l���xX�� '��N�L�Ԝ�MDV������*H�q��0\���Ny{9��7Y[���m�뫝�v�Z�"�4ڿ��v�����wo:�k�;Ů���0�9����mj�u��\d����q���`��Q�ר�t�{��xe��&�6�4��X���ȼ9t�^}�����{(C��t-���{jܹ�]3Ω�9�rfCkt��vz�gs��v�=.���Evc�u�e�+�vM�9��<��Ħ�t�s���.�&m�N����^*���2�%#"bd�� ��o�㙛�$�Z�ȢL�E��Oj��gcD��ɉQ2[:kr��(e��5��=�``��n6>6z�»����#��a!L!,XQ��+ݏm�A ��@�
�rT�.�wU�ω$u�c����$�zbaL�2�!�Ow�r���A���`I#V<�$�����V���
&�0���8H}�t,B��_W�|�N}Dw4�d��T�s�:��һ�B_�߿���9�+ivT�ug�Mu��gm�y�WN���S�Ύ:۱��ߟ��3p���9���#N<��>$f�s����%X�?V��0~�@rz?jGumUL������Ү���>���{rt��AFY�~�j��k��ͫ����Fh��ote\���'����"�R�.D���M���Z%���xxvž��'Č\�(�|2�>lb؋'������r�%�՚FR[:kr�>����2V�駉޷xA�<������b`�R$%!L�B�c�r�X]t��� � ��@$^s`"�;\N���%�)'R����ԛ��Q0�H�R�	ٮ��~$ n���;�5�[�ƍ=�H$_^s`�M�v�n:p�V�iD"Q��B�&�9{c>�-[pk�!��[n�y.grc��rm�/qfg#����Fx.z��7/u�E�v�;ЌRS�"J3{BA�ݼ�d���0���%1�����4���'1�O�/��	���� �F3/WR�8����5�H��j%g��<��߫�I5�n�)gGV-!�Y��aMt�s�"-�a���D#�Y]�����B�����9b�L�D�<�P�5+z�xu�r���/�}�����/����>�}�f ��	�d��v�(A�@�U�� �ۛ��A�8z�;hOr�x�v�	�\� ���"BRȄ:s]`$��H�}�=R�NOu��Q���w3u�I_eHB�f�P��������)�hj���m�S��'SU�m]�ר�6�@�w=\u�ϟ?~�d���]~�W}͒M�v�$}��Eó�Z湰H9ٻLA���ʙ�D��B3@ю�:k��˾�͐I���`I��(H'��w��v�2;wL(��S&J���a��BH�9+v�'z�;m�~��[� <;�����Qİ��Ll�ڌ͙ѧ.sj��	��L�I��"�9}��w�6��<7ON�5�)u[��eU��.*0E��@�	�0&�]���u9OM���.Jޡ]��yՂ��"���N�wY���x �²��QY�f ��	�d���^����|�u)��NG����`́@�]�se���S5�9���FD�L�$��Go)�J�Z��[�Eנt�1�f�yY.mc�����Qޑ!)
dB���8k��n�9�r��]7g!�][M�A'vT���Q10fTJ"�o�5���Ϗ�R���H�]���8�dQ$�w�����S1�n];���3>�>��I���Fgf�I1(V�bss�իqټO�:g������ّۺaD��2��o���W5��q>0zr��NngS�E�����.���[p����B�QGȕ3@���q���*���v+Öe�A����[���{�6Ld�)�����Ɨ��"�Q�_K�q�wMaB"t^{Ⱃ�=0z�Z�\�TҺN;;�g�P�'�#o�����Mw��%��'/Q����&�^n.އ����J{w.�79������J�=�|���y�tOyKA�tyz*N[�[^.��z�^i<�6SM���MR���8`�]��B$:�����ٯ׾!9����g���Zc�ɇ�2�[�Y�S>|��J��oyA���>����cm�3�l��f���^S�9N���^~TB~]�L�re�b>�wy]�:C�z@4TsR�?:{�S�@�1��C��]:-Y�ʇp���ɮ:��?H�[FM9Ԋ-��7�9��_v�]��:x�(<�,�\��^��z!��؇��ۣ�Gu���w�D.5��,+�9������,�p	��|;�<ְ�ZR{�����n�vB��J�;⻻�nÐ]CeM����sxa�$���qvM��$�s٦��zߙx3be�-���9#K�	c��[�{w�.sj�봐�R ���ƚ�o�(�����xyYS�wx�����+�7x}ZE�Z��\�Q^�I���p=��+�/'0�t��>��UMsz^����uA�yy�n�� ��uŏ����x�t�/��G"GɈ!@Ӫ����*�Ѳ����&L'P�Ĝ�W��z'��蘿5 h��b�@����;��=�U��Q��ر�rG�hWU����)��1��Oo�`���l��P�S3v��+��/z�^[$�CǗ��;�r5�U�*�Ȋ��"�2��DUt�գ*�$ZJ�Sk3�Z�.s��V�#\C�ar�%��hEr�\�1�9x����r�]�UA�$�UQ&L�-��� �%D�� ��U�-�N�(���R[)4J��0*��"��d��x�8.DEg%Q�⥓��*�-�i)!��˝D��]�J�QE�Q�t�Q���#[r�0��GJť��R(���[T�"9r�%�B+#@�$�V�"!P"ܸ9�dQBHBtQN���
�sB�P��Dx��Vi��D�.�%Z)��)*EL��$R��QEB�y��34�#�\��#��\�5���
��QYYʣ��vyGFd�b�)V	Np�!9��!$���VY�D4H��)0)�(�*�J(�:Z�#.xʢ�y�RkS��g�{��Ӌ�s���q��mѶ����]��w�b�2��:ɀ�'���촪�sݍ��3�[f�:�[h5��ۨc�_b���ڇtHG��E�L. ��j�n��poU��ɷ��� �͛����#	]��E�9����ܬ�]8��Jo4�!��a-�m���m*焊1I��K%Y�`�R�.6('�k�q 9ݭ��GT귏h��p�q#vB�U�v5�����m˸ׄ��w=m�{ �΍�( ؘo)vs%�GK�z�T�n�n����8ݮC�{<�E�t�
�>ٹ�v`I��l�q���Л[�؞;[n;�M����x3�nNn8���f\^�z]��ob�����͋t��׎6�:͎��3�Yt��Pر��ԕ��o@	�͖65�iہ�CC�F��{���+g�t���M~\��}��mO:�6r�:˺P9���{2����qȮ�bM���mӅBQ�t��p�n�*�>ys�p^#�l���>�w�> ]ǎc�\\۷۹�9x����tsߑۍ[L'^.-� ܛ��l�^��mǮW���uk6$G���K�x{u�<�Җ�-�sv^-$���q��N.�x�=�&q�n�U�wc�:�f��7c���py����X!�ۦ���/;�K&�Y�^���N����67n �J��@ۋ���}5�g��lf�6���۴�6��[�P75���.��;k�,\�=D��a�#�ku�4Fv�q��ꛮ��)��f�xKg�������Z�X�3��n�j&�s�9D��u�l��	���ݞGq&À�p��zr�ˣh+{7;Frv���kc0�`�ڮ[O�����:��Y%���c���r�'ʭ�{^���mr��Ⱥ�k���k���v��c\��&7o5�׬��A��tv���=^c � n���;�vg�n�ͻs�Z3���@;]�fe.�̘��Ux�8^�4��̖n�+`�{������D�9n��l�h���Ħ�����{�����m�m��Ϋ ��6�Cg-�ϣ�\i��\6֣��qε�s]n����v��H-���m�%ľ�;r�����6� +d���Xc��.�[��'V��{s,;�@D�'�.&�u�.�ɞ�=c��Åw�u�0�ڛk��N^��C�ݝ[n�]�=��1�4��[s�ɋi
�jx�:��eݵ�#�$gd:sLoWd�Zە�vJ�@dt�Ii6�z�y�����Y	��6���vm�3e���u������ꍎ�'5�BO���� ��n�yl-��������X`��=!�)�Vu=l�z�h�kyQ{�`�H����>�^�`�f�,�ȁJ��k]U�w(��1*$#"D���`����$��d��y�m����O��k��ܭ6q��
K�_)��JKK[��?�vp��`�A���tD�Fmn6H���aD�D��J[oz�$�׎T�<*��z[<���$���a��s0��J���lOe�۶]����ŷm���v��l]IrX:��.�&�wa��?�>'��3��=�����m2|H$����4�R/6�`�N�f�	򦷌�D̔�S2�#��P��W�$xJ�B��5�6'��ү�7�B���cg��;R0t���o$N[i�#� .Q�l-�u��7�*������]v|��9���$�w�РA�{V�F1�S��B��w� b	�����O����P'(E#ّ1��p�}{٭��H��#*�L�Q)HFD�oƶ����P�z�,H=����$���4	 ��{^���1E�w����X'���(�0�O?^1�`��[��8�6���:��u��$�w�^�@$}��6�s����]+Q��Jy��q��9��]�5n�Nn]2�Ϡ�v�b����FH��R�7}m�m��@��;���]�q����f��A ����W�B��̩����m�t>ۛ-�f�W^i�ڮ�۾��>$;���#�}u�J�⽼�L��UT%3)�:��P'7;X�A����2m�s�5�ᢟg�3��-��������6�kc�:�ӷ�Q�����k!���EN�P%�J��G.�����"����Aw�=@�}��*U����&dB�z���F���i$mwW��A=����;���fnQ�h�B���9�&L��Q�"[5��A��ݠ�&,jA$�Κ$�33���۴.�C��,�ϔV�s�E�s�FΎ�.��ݛvkB�tu��jѐ���`ې����~�W$Ѓ}um
>$��`3�|H���=Kz�p��x��&�w[���FH���m��l��,��Tq4;^h�I#3�['ā�۬0	V2�b��
r����$��~_�l���s �S�J�h*޻��$��7['����dĵ��/L�I#3)�k]=�#���`��]A�ٻ��	"�ui��g��T~}�-Kh��)ї���W��b�Ȗ�Y��jT�j{O[��Zc;T��;"�t��3U�Nn�!
9��&'������߾����<�o>臜^�R8h�Ͷ� @��cnG�O���c���)�^]�D�7[��ci�L��S�8�b,�$�dS��:ݎh3mnj6e�ե�h�{q��v�=v�?�>e�&*f&)R��H�^m��"3��: I��M-�LNd�Mh�On�$?x�͢i�"E$��F��<'�g���g�owԩ����<�@��%��Bﱰ$��ugQާ��%�٪IRD�R�������H�1�����}�$N�]�� w����^l�sG�R�ÉiZ���~�K�;�mO�V s3�� Gnc�Cfv���J���n�6����P}R�S�}U@EU��������ҳ!�^˸�,���� [�m2�����:��n��U���-���2w�w'^ꇧ@���>@9�-��;��-�FM��$�ܽ�{�W0��*�y_u�{>��m���[��2pc�uκ�U��g<8E����i���M%�ݰA�kre���W<ַk���n�u^},�3�=���m �G8�l�ηQ����>��ط<�[b�u����y�;��ᗕvNݭ�%�^ݬ��C���z�7GS����Q��s�R�=�dnu�=�O=�\���h�^s����:9�۷]�[t�/1��9�1�z�nɨO[�t�۪�g�G=����(�9�v�#��t�3R���õ�ߟ1���"%J��c�p��C@Ǹ�n @[�ߤ�NqhK�_�� c��$���}۠�t���,X���/�2n��8�5�P+9mU�J%����D�$�7z���ԲI�{�zKncc��SUT���0L�w��j�in��d�k۵�uê�O�y٥�W�與{��@,x}=��iŋQ)w}�w��uw}]w�߼ '�ƛ �����u��<}7�2��9���٠&�!UISM�o���X$�w��B���"�"�J;�ߚ ���� ��i�PZ���S��aP���͈7��g�;F�����<���y����0khe1��Lw�#�!#*f|Cq��k�"swyش�D���p����Q�Pn����$�go]�`̢�|��kZ�lJA(Y�1�Ti��4�u�b���r�ܛ���z��b
�:��/_y�{!����Hs̞n���YS�f@ִ7�L<�+"�E�1���S���s�	/��%:��؀�������7j	'��;����hD�(�2�%11S^��m�]�`��w�*"��~�*=d�� ^��݀��7[�NCz�I t�|��߼*��V1 �-���[Ӻ�� c�Y��gszw�a\�������31�T����?���� <��s�SQӓ���� wk����3M��$����P$8�����$��`�&�Y�ӌM���Ax���r<��l���wW2�HV����5D
�J��H�u�݀�n�a�>@��{�.���4�Ꜯחwa"Orݧ)L�9D�)J��-�!��؂<���,��[C�;ןX$�.��r� �X��� ��o�G;{Uv���fe�� @��k��pIh��s$�?���\���/"��W�.~�{{�"�����ɧ5�$�ԝCSh3�]�;x7�b֛�m:�mܗO�z���g�xͼ�I${�O҉(1����Ol��J�T�3��z7�;T[�߂#t�� $���D����wrfn�p��]Б:͍���}Ф�X���:|r���q,��w�R\FSȪ�wQ) �+4�@+/��H���;��F��̹q���|��<�+�a�ά�t�/S�^wn��gדT�<� ������r퇮������������?W��w��`E�yfe�[t@.cx�4{Q'PXqQM���ɐ�F{��������Ɓ����`|����@�_�:��2kD�ٿ��P�B;UP�����~ A���Ҳ �{ǻȝ~S>ˎ��s� �>�� ����F�|�,-km��ٛ3~`͒I5x%$�y��d�H,���leX�c7�h��-Z�Ҫ)�J����*�T���]��L��kxM�[����S5%�nq���B��������|{H����A��3���59����~[���b�ީ��$����W�����i$Nrͦ%uF*�چ� I��L��븋�8�mP���Z����_~ws�.��k���g�Š+����7]�[v�y7n�85������2����n��a��������Z��t�]F�^�ŞC��~h��7�웡z �%%)��®�maOGp}86# 3��[l@|��ݤ�3�[�w��ߑ�ħ��~�5������{�=ݙv�>����9 �⽊���s��%�wu�6�Y�؄��=��TUP�����\^��<$ 7��|s�X�DB�vy�"$��6l$�s{vM�2�#|}	�	���u��	�v6�lJ�wm�\�f"rsn��I$�fƷ�"벨��5��ȟ�.6TUc�sBbQ���>�Y3LG�
�5���D�5&����A��(��Fh5�8{�n�y��f�f�����b� �����_�gw{'�߆��É̮ۚ����\]E۱#m�3>zܧ�<uO���X�Gf�1���n�m�wnv���n�7�g۶7Z헧r[u���V���	���c��v�7Y[�9�2�nN�U��<`Gq5q��]\Vz�%6ۗ�6y]pz뇲����7��՟I�^�ʶ?����w��5�W]�KC���n7�tr��\a^9�P���M��.���	��=��Ѻ-/M�z�h����y�����k�Q�8���?���Skq��2�k��'/�i�I�n�0��v�sô��z2��H�己��=�4��ŚQ:p.`c�~���{;���=�9Y��� ,��c�B�v6�lƻ�X��K��s�^S��0)DJ�AUT�=�-��!o�l@ �N��R�7ꩬ�m� #/g|� �~�o���٠����*��ѯ�/�G������	�|�A>��4� I v�0�(z�{��WG���ŷy��ۖ܄�F\j�EEARMMC`���@�7{��gk�]�y���X�[��?�^wu݆z\��D�����n�� �~G���[ۭ��K�F�Nl�tS��ƫ���]R�gg���~���y��Hu�w� Y�����(�X׶���:�<��M�!���Ͱ��ʩ���
��������Ȏ{��>�s��aƙ��Ma�aN/_fl��R�`S[b��{oj�yP=FN�&��OQ����b,��I�1���g���J���6I z��4�@_o�vM�'V���_���6��{w/�4��ŚQ��������� ���j��c���;Ӿ� �v��@���H)����%L�3;�5���&t_Vd�wDx�m6$�fwuݠ>��Vo���o�jc�S�����u��IUUAM��2�X|�׻^���qoy�-v��7{��"�:�J4�wuU+���5%#Q �)3L/\�nSb�.J���w)#��6d�/Hܱ���~|���T*�D�Q��[�i� ���jȈ����4���ڜ��� w{���N#A$@�`Be�um�i�m���J������DA����@ >:� ;�կ������S�s��)EV��
Q^����F^uy� D?�0�����B����i
32�^k`M���m�y����;�
x\�oC�B�:q��6w_0�]��9������ٷ��j)�YQ��Η��Nlh=�M�ڕ�5C�X7�sv��z���MVny�c��t�b�vv!�s���w�v�at&h1�K�P���z��,Z�U(˧AXѪSy�D��4��5ۧ`���_�$g��� 1]M�I�G���l?G���z�g=Zq����ɝa>��%1�n�`�h��-�ݫ��{�]�˗��:!騽^�>��Իs��̇=��Z*��onUz*s�U����:���f�����^�{9�!K�釖�½�B�Xn����ǯR%�sN�}H��Դ�azu{���~|�*��T�A��������ă�(��Zz=р�VD�E�vt��<ơN�a��o�W?��D�9j�n���[TjT�((ߑ��0m��M���w%���h8½.�Z�(�o������Q��d�S��	Qm�	��<#�I���4b��Os[K�I�^{M雎y��zw����r_N�׬´K�W4l#Q����痺�&@�k�B���vvx�}vbT��`��#�{�\ބ焹�����d{�ߦox���(̻�e2H<Y����}�Fw�m�{8�K'0���`�r���Six	��X�
}W�pe�즎��/(�f��@n�h�{ӻO��װ=�q�e������6����zhv'�S�G�gz�c�L�Ʋ���l�rx�{�U0��Bww}��E~�$ њ0`f�jA�PY4*�PUM�q8Q*�UP!�r�e�j+U*����iE��
!DDE��Dː\�
�]�f�h�T�� �P�:��G5dI�l��$��"���U� �,���:l�Z2"�U�UDT e��EZ!g�"�eȒ�"�B�ȕ5(֦�,"��)�J�%��ڱ"��s�4D��)U!H�ZD�XTQ��Q��T\֕P��9YP#��Q��4�P�$EYQT�H���Q�]D����D�-$�UJQQs��s�D�ĸQ&ʩ�)�'EH�G4��YZ��""��B�x�NDP�Y�M�QNZDuX]8�Z�2N$tL�ĕ�q�K���gXx�"��(!'sr�"?%�ٹ��|߻�uݠ�Χű�Ij���&�8����@�����f ����`�A��^���W~�^ŷF
f%�����<��aH�LJ�PUT�{}�� j����^�Zܭ5 ������e�טA�E?7�ͷb����ß��	#�B���y�4&]m�`��� �O7�������0v�T.�0�(��$"����}��6�k��>@|�u|�]~.�&���&�� �ͦ�Q����U(�Rh���V�:9�$�yĨ��b�  ;3�����d_g����-GR��yi f\D`$�"L�X[����|�b������,~�켾 �:�A ��m0�Q]�UMU �PR�s�����7d�� �s�h�D��ʧ�Y��v���9
<y�ЋQVX�$�V��f�bjdQ��ݾ/��4�ˮ@7�'.M��p[O2��(�6.��~�L�׿���߼����OQ���2J�&��6�^Kw��v�M-]����{��2�%����%���v���Gd�*W�g��6�����獺��vİz٬����;]��T��gvJ�"�AUR���m ���c���,��g�Ds�=S�����l" B��m�=e�EUDHT�)��}�v�
s�97����]:�%�Jg��I%��͓a.��C���!���L��?aq��P����f�sq`�y[o�E�8ɽ�-��6@�3���Ҏ�"I��ݧ5rU	w7?a�[�z"!��u݀�Ffu7�qO�:�}��Ʉ�{%T�R�)�1�}�U���^a��Vk�w~��`(��~ �w]���̞�����'���Y��w�ٓ���˫x
s��
�ws�	T\�@Ɉ�*�fzߠ�/׮�R��qF�>W��C�w����ٙ�Æ��4�d�R��k'��|����ᓈ��Z��.si�,v�Z��lX�d�cv�m�Z�/b����lN��k]�h���U�S偹���6^�����nۢ�<t�Gd�zN�^Zx�9CFG���sqX��g	����<ݹ�R:맲�q�lq=Q��\�/�l(c�zs�)&X�������xRx\���k��ڝ��8S&�d<�����gL[�6J9��!�����-D�h�R��&��b����v  ���4���fV)̂I���d�sz�����)��+�*�[G�c��*���;���o��	����v ��� �bO�����mnk#�Y�ELR� U(�3��-ŀ�nd z�s�ǠFh����Dp��wi fd�r��WȄ*�����m�y-�r\�e���G� 7ټ�+ s'�~H�6{+���s�z�$��ٷw��iF�H�$���{j`�J	�ƛ�U�b������>72u�l�7�EuR����
)D�pq뎃wc������{�`Ng�u��=�v������%T�R
 )Md�ǯsnՂ �3��A(��~h��I�n�>��@fޘj/ڜ�SP"h�R��@��m��Cب�
�g��D���c<�@)��L3ԍ�y�{�E��C��=w%�>�:j��Lӳ���=ōH� ��hۭ�J"L���T3O&n�-ǯ=h�W�dg8~Iy$��c�ZS�jM�Vz�2��;�bE(�����qRo{��� H�qs�2s��k�| �� ��`�Yg*T�
X���}��h]���	2��@ #+���@,��*�{�9�ǒE��R'��D!2��Ri��c��$��s�k��,��S�������ȍc�N �>B��m�gw7h#l��lY��
bi
bQ2��P�
��������%�2&����	UD�F�a5�?~����Q�0"4���A'����i ���� ��Ϋ�!�v� �������Ԗ�%hL�����'�E��m�ⲳ�w�9 ���與�gw]������o��9��7����%�T�u���M� ���v Ҏ��o��f����0O���ɱf�7k���ո/�q��f��r�D�A	����:_3HI��X;���F/�8��(-�s&7���̂y%�2{h��7���v4�%>�3�U+y��݄���6�H���hv�]�K�%���u]>��X`$G=ڢ�u��)H�"RQ$�;O�g'qf�3��HU8��0Vc�K�!���w�^Y�9�*oP��Z#0`���n�����ݭ��)w]�4�#�	�v�熈�u=��O�Oa:>�"�RT	Rk���yTK	f�s�h�䗳#9�Jkc3��J����x�X���	/J�Tp�eB1&C'uS��	��_�2{�+��� �[��w`"I���@d����q�&���~�iW�aLL��))�-0�o��։'3#�����67U{v"v���?�nou����̞mH}�L������*�4	��Y��َmK����n�V |vd�M"PB籟G����\���,���xg�Z��_b�G.�5C,�>�S���H�kr�E��J�3ɤ�����t{��㬑��U��F�4���ϰ�E	 "y���%��;dRD�}SU2����C@ [Y�7z�w{�j�y��f�h�Fe�7$�=����*�cfuےJ�1*IQ�p�F��1z���ۣ+�c�^����2�����2�N՛�&�*��j"��o� ˝��H���~a����fu^�q�G]�6�(��!b�*	UR���|F.���{2U�NK|�� w;ᤂI����&=�m��#�h�^<@Q^�uJ�$��"e�]�R |
�fI�%�7���*��Б+��6 �+���	+��b��d�!S"�{�sw���M�� ����������UBE)$��up�����d���*�D/{www;V����x��o7���X�� $)���	$;7��U/��^�z�\@.��sw8���ץֻES7}{���3_��-�ΑӊrkC5魬I��#aУK�"������5#hk!��$��$�M����n�;�\r�=��q������cw�`%�y���6W^�G^p��iE���\iw+\o&M{�9�/]�����Y�q���F׳j���V(3/l����k"=��VL���t[�y�^����h۳v����ۤy�1���é��[�-h���K��^��y{*�v��d\���ӄz�u�kuӋ6O9���ιs�(���W����fK�K��3pR�S�mpu$�ݠ��t�R�+ꪩ���N���g��I%���&���1ϗ�B�Û1� >�c2\�0T�Ҋ	�"���yv�9S/��Qغ籕bI�����_ ���� �z�bח��*�K�7����UEA5)�]��� ��������W��7W��c@ >�cl����n��Ez	�(ʄba�Zӎ�Mp�f$N�D�c��b��{����|d]�w5�]\^�b�b�1�ӛ:�Z
H���V���o{��iy"p��I����G�jIGz����oou݁���6�x�F|���{s��%�c��Τ��s���t$�:2S�l=���*� ��u��p�����>�Ӷ/eY]�&�n"#{���`�h�4Y�Y��ɣ!{_{� ����_�҂���)�����%�����ʀ룘x��F6��L�V��Y��ߓ{�ot�;�2�5������#�c�=8��tv^Snm���A�de��S{F���Kt��́.��wޠ"o�vＶ��]��;��+F���"�Gu�ݫ�� ���f�l�Wz�3{��� ���ׁT���ȡ2���0	�̇8��s� ��ݑ�}�޺h"]��ٌ l�������-��cڎ�'tj�7h���[~�H$2�uՑ�gS~C{�݀�6.��x�+�sl�^�����m߯��aX���M��jR=���j��m���K툨�x��?~����l�k��޻�'�S�I(w\�.s�n���b.��]ݤ���w��Ic�@�*e
�D/c�I�-߻nń˻�u�98��� ���:h"!]���L�z�'lվ���8ɿ_���̕-��o7� @�������ȸ�y�bu.&�ʮ��Ӷx]�h���w����щ�<���1��]�{��>�|h��Rؼ��z�.}��H��}�x�]�m�N�����H�fJT�9�]��w+vG1T�H:3�� �y�0 ����7~3��̤:+[k��b1^|@��	��M���i�I���~�D��b���T���ݎXA���o�@���{���p�&��G8��߽��|�e�Ű�fqv�y*�g%��|�mWmt˸:�??�>��=M���}�p�����!e�4�@�����4�+&"kV���Ư[�	$.�]�S�J��fh�!SC�=��qh7ȇ�.�tfz�ԉI#�|餂Ks{��'�FNP�h�;�R@��	I"ba%�	��6�Iv�sd�f��4�{���<�Q���i� 77��"��o� ���5|�խ�??���v]w�D�Y�mm�πH�{z�"":9ߋY+����.	V]��u[�����|�����(iy�m�����:�%\qjr7b7�*~^�҆�
�{��<n:�v):*(f6��b�F�r��D<�H)z#`��Lf!)���.ŢR\v�lgx�U�sx��[۽w`tu�q얷�ӹ/:2A��i�Zw
Ǭs�vs��ʭ2������KB�6�v:�?C�}�D
��Jio��7��;� ��t��IU�̙Έ��g�-�c� <���$�t/C�n wA(����$��	�6ȧ<�A"W��z����	x�^ w����W�0�[��j���SMG���Շ�G^S�+�*�'�e�WUn֤�Kww���GG^y��7j%P��jD*t��l�X�u[~(ȍ��<w���.:��@ ,����3���}��w��8���ɉ�0z���$y�A�&f���m(��VK��o ���5� ����(��^w���+���iڜ��%���t�����O���"��`�w)�C�˄w�1��� ��M�N�:8���c�z�l�ԇv��}&<���..�׊7��w��t�&��*^ܱ_&���L�7�ܽ��f��vC�8�ǽ��
x�� �	_���]�o�r*�5�ü�[<S���"����{`YJ7�����gse��s�B�w�q+9|��)�z�/h�}@�䯦[���L�
y�!g���N��ܸ����Q��gy�H���s��|
n�x$uA!��y����Ȟ��꧵�}�K��U
iY|Ȣ�i����ڛܡs=~�W�#�"�Z�{�s�1�Fo�y�xH�;���a��v����[����b���v)n�f�ϭ��fh�'��(g�ϻޝbѳ��^�4���qj�Y�w_C�葚9�;��~�7�[nm�|a��2� 5�=�oc�\��0"Wg6��{��{�Y3Q}h�Y\	]PԳī��깾��t��I�gޫz�X��}z�e��;�N�r���]{�g��$t��k ���� �����Aq^��IM��ol`N����
��^)|ߦӶ�s������Ek$�Q&��1�[��Jgbуrs��q0U7���}�j����pj�E�3�w����x�t���Wz~@�����ϴ�c�}�Z��x�.��.��lo<��m��s���ܵ��- �yg����)�1WsN�@��H�@$�pq��$�Ef�:mn�rwn;(<e��s�<�1�N��&q#��<�B���p��$�r�8�D��n�QE�'�-,𵜳r�B�j�D�ۍ��%]s�*\B.r��Qr �
�L�^p��pER]āTQQDQ�P�ǜ���Mù9 �{m�p���Ý,*ܵȜ9J˙��Y��,������n(���H�9rs��(���dyJ���V^ss"��PDfUQ(9�������*�')*�s���k���
�Ⱥ�-�B��A,�8K8%�+�r8����˜�:W�J"�8Kȅr-C��9IyTШ*�f�UV�x��1p#�L�n;���*�I��Tqܹ��\��'pK<���pNr��Q����QS�j�pZ^�R(��(}��똷O8��q�I땬,0�����1��u/��)Cl��g�ە�`-�Y���6ɹ�!;g�ʸ��n�s�7*�
nr�`��k��>��u�^��ۛs�����c��.,���v�q��ڳ���c��P<�8; 6����uϔ6ۡM�m+ur���u���e�\S�SY��Gf��mq�XA��m�$xTi��z��/.��v�{\vW�q�g�:N��Y:gъ=�[&�iKu�] �nR�m�nUv7nm��>��A��r���-��Ŵ[��^<��)�r�;�e�tsm���\n���&�����n½$���բ��睺�7������=v�C�wQ�io]]i���j�KsW��E�sv8[�nԫ��+j�H��=��/^��'t�dxv�n���6����ϫ�tI�ڻ8觷�=8��ggsv��F��Qݹ�Њc�xwm�탓���*b�9�������zw<�����;����z�]ۍ��NXz��]vf�m��d��Ӻ�q���;tP�䮆��y��$�y綸��x%��nP��Ļ��ۏZ���1�.�=�f�H�.���*۝�݈v)����F+n�7����m]�9ݞ3�����9N{��c�&�N�x�����ps���?�p���֧�[�u��Z�j:��n��x릈�t�2soV�sǎv�)��ݛ�7ю�K�s��!�����͈� u���b�����,l�1���{�3�I��h�'�Op �W/[C[<h��~[�'?��(i7;��qk��[��vsN�RI͎�����f���g��y����Os�W�]�y�b�=g�a�;b7Q��͓���v���v��r�t�9ow=��۞�;)��pXܹ]Ss����֗����Lv����%��m�m��vw���qD�1�8�a���γ����e�,v���8ֹ�l	���<�ը=6��2��-�aNh�ԝfp��g��9������*1ۯ/,9�nut*ڲ[��ꬼs:Kn����y��hA�`��\��4mnN㕽�Ü �z.^*�w�2k���ѣi�FH{��<�\���Z�6��m�[�D{q/K��]#��>I��jwi�P˞��7[]��7o�F�m'��:;(e���6��nИݣn1f}��s��BM�W)*�tC�َ^n{�B��,m�G&�\h��^כ���;kY8�p��;������6dL��"_��k�d�t���D��9}������^`k�~�����@|�2:��) ��"��fB��	�ڢf��鬾Ι8�3���u�D�$���r� ����d܇wʺ��I��O���5)U�ˆ����vcl���S�h�߽����H�G^��@�ٔ�SQ�""e(��%L�d�=�w�k�W�(�lR :��n^?0K�۽w�n����g����V��G[o��N�ډT(A3B�N�'׾�wo7�V&����m̛��t��yx���w��������ι"������w߿�P�����S=/N+��1�l\�۰n���]t:���/����q�9�CC�����JHn^?6�&�w�&�]��k�i���H�$��7/��`��$���M�{��ڰ���OqW�>yX�T���Z�;C<`��B���j�	U�X�L�jFOu�����c�O�1߬ɞ��(�nD������w� "������݀���f(ۚ�Um�@)x��L�3!Hm!�q�Ā�77y�V  �=�U�]9Eo��#@u�2���븃J�*� H:�,{6�����<��%v�n��vv����w` �����8��ݨ���%ly �����)��R���j�T)�L���z�Z%%��i�r�l��ӆ�Q�[~` �;z��@}񑹭�'��=_��N!�#�����I�V9]Z�I�g\s;���c�u�:����o=������g[�M�{|����Շ� �頎�{������+x�d ��z��I*����""}2fa�z��RA$��(�/�Ͻ����6|@,�޻��)1����Kf�m_�J^)Ʌ54�*d��l��.Հ67w�$�Q|�Ms޳�USJoʫ��f��}�<BÓ���_� ��E�vS�T�?G\��g��+��[��=�D3)z4�O��3�n�䯷y�I$p��:IH;ؐ%zd)�FC$um��[�s{aҊs(�k^��� >÷]42:���p�9P���n�u��(���QX\^ے��K^0ꦕ�={;���z�.�"dn�~ @z�)p�;�}u�ԥ�6!D�b=ɱ����9(qA�7����m]O펻h�@v�����f��K)#G�����@?��ב%���׎I{٪7��b��۷v�n6�"n2�J��D�(R郎��5�{�=~�����vD f�㖀HG^S�RJjf�=';g�^�J��Q�D�5�TUO�'��� te�O�1׼���Lٽ��}{�|�^y�@$�?K�8�`�h�Z���Jй�ߥ�қ����y������j�"2��$����D�.�/ji���r]���ޯ��+�&�^���y����8�.H��w���$\�Fk|mAr�e���m�(�#��o��Qx�"���T�6��ۍ?  ���j̗�et�i-����` ���lR($�w��q�a��r��&}��v{$�`�ݒ��l��nY1�G�K�R�Z�cHD�Ks�Bh�S1��6;������2:�� >�{��%KȾ�3nge#8�mQ�y旃�>��ST�*�I��L���[6���/UP=���Z$��o?���n""�Z��6���H��R޸��%
����D?�{���a� q��_W��*�$�$�n�A%y��v��=B��O�L�2�s�a�g��6��2g1��/���n� ��5�A�:o]�=É/.3�ߩ�qȈ��10��+��˻� 7L�5Foݗ�U����
�[t� gouݠFq��.i���k�i�`#/6����m�B��C"��'?*�H�!=ū�O�����5l��(�x��h���$�?>�8>c�S�ߡ����j܆���u��;KI�+vF��XٺYl��Z��=:���	�9�a}����m���޵��\���W���m�\60g�v�;�PJV��uqг&��9]�+����z���������b�p]��^b��N��V;7=����NCa�m���wb��и�q��={�	޻9�rv��6����Y�U�ɱ�]��;
<_�X7N���8�m(qܥ�v{lۭ���ϳu�f��X_n��{���^ݼ�ut�� �Ǎ?D	��;� ���5�
e�|jr�u��Vk~ A�����s.n��a N�7_����/����mGf[��H�2;5��{'K׼?$s��*��q�U��"RX����3���� ���C@ ��+'CGn�IЖow7a$GfԖ�x*H!B��-&_j��Y�LV�m���;���\vk�� ��|�-����k����%.���$�NЀwЈ��H����n��H����GUu�Ԩ�����]�X��� Y���h�Kj���b���$�FQ�g��M�m�)�N��Y�ݺ\�P!�y0�]�Dz眷
ZJ��{|FjՋV�E?|g~�HD������|頜�l�y�mu{s3���@##�]C%i�%�����X�>���?g�{E�gl�=sh2-���?s]����In�Q*vn�����7�p,F�P����۹�n��^�SS����F������}` �i�I$�O��p�-^пr��3|��TU����`P�~Z[�$�Xn���+��]68D^e�H���ky�A�$A'�Ai�VjH��<.a�}�4j�W/b�]�E�.� �"����J�Zn򤖒��w]�*����cmrG}LR1�H� ��0��9}S�nws���cfv�5�Pmۧ� LV��I�~�$&������7�#�<t�1���lQ-r�^n��b����-���{0�n����x��ۛ���>�&u����l]�O��^ouݠ:�AVŋݮӉ��y��Ex$���n��d7FV"�(�f���L��n��~�`�ׄ�]{��@aw���}y��w�K_-�k�Le��Q�p�蒢dHl%��ߝM��;�Dǂ�.균�rܤ�K�FVoI2�ddf\�t`:J�)�C�MnC��a��O����E7����_q��x9���a��긤�cc�W�x�@~�����No��;���}7h���J(���z�QB���+Tɟ%ŷR�I ������d�yl���S���!#fyԗ�&&H�"
�L����݀�پx����Y꼬�Z�x��M ���E������2vL̼����	�ӹ��<�95��v���]R+��v�=���\_�{�ϝ�<r��?o���|����w`�Dvk��Y3��c�dk��@����AYJTj���J�|�1�m� r^"�n��f����+��;�m���6�DD�j���2�v��OE%�\.9&%D�ESd��.Հ����T?�A9��O��2���� 	^f�ݠ FGn�H��dP�)LȑM.:�\�s�>��wd@�Zv��D�}����7��gn,{u��Ys4��;x�`��vz�B/%W2�dv<.�Q�tUc�f��[8"N@e��2Q��݀�%�UT��D��Fǽ��H$���î�~\�fn�;$�On��^X{u�,������m�?�߮�n��F�^�F�s3ӛU��Z�x�V��.ɴ�&���׷ ]����}j�da4�/���� �c�=P�D�c��yir�|E����wi �û�%��QJ`1 9`$��'S�UW�^J�yy�ϭ$�@b��,�:_e?R$�e�R�5��u^��x�$�O�D�7����"R\^c�A,����Y�̙�ޮ�}n� ����#a�7���}�%���BL/���a��B��L��]I$�9<�$�����1v���p�L�st�H[�A%A�̉N���'���v�9��ξ�%�uU�\>�5�fw]�?utT����^{o\m�=��/r�s��W��9o8�Z2!���i��k�p��"ߓY �p~6�Fv�L
���-����?<�Hn�t�^8��xx�l4nnbg�<�F��ӻ^��a1&7�G��kS��eӷ	�7=���#�k��t�Ӳn<�u7.��1�;�۞�^{+qķ@\��������NZ1��i{[<�����\�DQ箝�<��/@I��\f���..�� "7[L��s����Ϝ�J�d����bv�y�K��ׇ.�n�???5��bv��s�g�'d|��,5��u��!�/Y�)��ڐ3c=R���߿~�ڴ#��hV~
�x�$�X_eI-,��l����h�ɲ��^mq������>.�x>��Y1(�Q&
�L��|��$/���.��q�~�  .�ٙ�w` �Ө�̈�O^v
K�F퐑�DTʙN����舋��w`�6
"/�+�ZD����ǩVfw]�`N� �P��ș��n�����vf\F�E�[��,�� ���b���օ�ؗW ����#�M���A4EW�;�˴� A���x���*�GZ���Ѽ�M  ��7��"#���?���Z)�������0�PCV[�=G<��Ynܴ���@ۣl���9n�M�9�t�S�Fr�?PMR��1�? �o6o�/��ٮI	���Ȼ삎�-�'��U�`�G�l=��$�h��"����<�fA��.����f�h~bCy�-�^�9���GrP��!v#Qʹ�a���ҷ��~�����y� �A���w|��]��݄�H��[�"L�u�.8���)�����"qn���,3��~� ��}�����<0�m�Wl���H���v����yp�*T)������=ڶ��S�٥�b��^7 tv褐 FC�uQZsF��9U��";/��I
�� ��>�0�=β�I%��T�5x�����m��$���~�I8_e?Ru�^B�f1,�K��ݵ��d;�C�nQz�㊞�W�I���mZ�)D�XђL��
+V�Dj!&�[d�	i��~��%b}�ZU��G�Os�z�	 �����
�H&"R�`Hm.;yR��v�
�V�{X|iێ� d>�׈̷�Mf�Z�V����h̩1�(�Mqo�Ia}�K�$���[�.�~��+9X���/�v�F���u��c��=�*(��F�����<Ϯ{XW��=�魬:�T� ����!F^��f�B����M��r�7.���}��c��
Ցʶ�'jVʹ���-H9���l+��ͨs�i�|��w|8𲆻�>��*^��C-�f���^,��װ`��v��ah�7_��d$�Y�Nv��F'�����}��fʉU��E8-���	�����}�۬mG܃�bH�J�fM��c�\>����-�~�{)���>j��C|ո�qdgx��$��&��)�73�(X�e��%���b႞ q��О-�8�.�v.���`�6t��������u�[�^��37ۓ��}���5��8��8�����ƣ�)�1I_q��yϱs#	��sN��l�?zm�+���H�L��t�D�����]�`����"�u��ϯ���]`2S����j/�@og����fwB�p��'F4�S��3��c����~8&ySq���:�{��o=�g�����e�OF0� �1���9�}5�=����{gn���\m���[��?��[�m�h�n�8=ώBuz�Y�ާC�qmLn��Ecƃ�L9����nr�"d���Ir�{ֻsg�3�i�b����{K͡o���H�D�&�]�Fv!���a���뜰G>���m�7,�k�|5ar�޻f�vL�}�9�[:ηjr�E%/. T��:H�s�+�����(ôН3��wU�+�*G Oz���wp�H��0:t�8�	�x�y�d��(����Z$�7�;v�q���aP�zEW�8�p���\"�+0��rj��*np�Ir%Fl�8�Xx˹@�x��y<�rD8�"��r;��f���
q8��s�G"�Q�	�S��')����'"GqRl����8p�Z�QF�p�$��Hd�p����UkHT9x���=�����3�1����DVdJ,�� ��wr�%jW(+ �sȉ!��haqP/�����+��q���(��9YW�8�9EVa������"�(��
��Z���M"�幜�a�&E�ǃ�4[��79�<(r�&y�l��qE^5t�\�x���5$�g��"�T�J� �AA��8˕Q�ˇw���*�Nr˹JCP疕剓�,�3���� 2;q�$FC�m/GT��Eac������a����4u���=��|�`�0�3�z�bgzx�]��~
Fu��P��&%:&���t�K�_v�kq����(�C7�}��:�`#a�7� ���A��f�ވ���mӤoI:�	qIR)����l� ��`�n�:�o���}�ң�Ҩ�UO���mx6cO�$�����%��cnzv�L�uOԊ�	���=��EMLM4ESh��$�#��-����|��I?������v�A	�J��S��u�߁\ҳU}��&�Rm��z�����XON[e��һ�gEv�w�|��<׈�����]8Ȫ*&fI�R�4i������Z��L%Gr�t�^I���0�G�^󿶉���ӷZК�G<еӯ����]�o��������[��^�+�ӝ�!��y�k��6T��
96m�{������Ѿ%-�6eH�3D�e���v- �:{r�����{O:��Pq��4 s���"X{qɈח�\W\�^�mf
�	0t'7�ƺU"�5;cu8{L/[��Z�^�^v���Ԛ��(�P�jI�W]�8��I��w;� ���0���}��WkFE��%����]ߒONЀr
(D�2&e��rZB�K�2�s;:7+�S��0n�uݠ�c���u0j ޭ�bj{�=rmպVZl�v]݂@F�y� �vfv'iՀ����@ �����}�W*�
!MJ��lnb�(hs�T�� }nՇ�/���L�Eǯ�U��^R �W���L'��(!������#ú�
I$��~u�23rp8{��U�w~Iy$��ےI`+5|�-u����n��4���Vu�@#���6�I��a�eV�jA����8Р.��W�7�Ӆ��Ɋ�F-W�
�
yĎ�F͸n���,�ZnvܖC�����g�n7.�!��d�UI��}�I>��Z���8N�uu��C��q�S�;�u��϶7��{qe�F;ZZ��;Z�&�<z�8�E�����	</v*]�=1Kۭ�ޣd�\�/2;m\st�]�Ʉ�@��^К|Z�Fy���e�^�mr���8L��:�
�[kq���3���{{tv�<��n�ټ�����ճ\�$mQ��T��x-�)TMM)��2!ռ|�	�u��  Y��Q�K���r5�z�;�Ým�J��Y@"eHF��q���}��<w{���Z�>ܞ�- qo�K��T��tl�_W�����R��Ҩ�UM��[t�l[�� >7z��r6��}�h�u��`"��7�Eb��RQS%(���m���G���u{�˧h �/���8��� ,���sۊ�#�Q˘qY��ɫ�}����M�M�7K����ūӼԬD�܂M�|��o[��	 �gw]�e�S�I9�
P �H�0JS�D�ٵ�S�ҙ<k��q��Ϭ:�mZ���4��������D3(��*v9�~ �|�O�@���v�M<�tYG��D��6��PI+6��HEA�*D���&/�__]��Kw^Œk�\�r��Yd8<6ݙpY��--�귂����s�(�W���wom�?yF����
W��c�^����b��vg���^{+�u��{� 跾��3���"/f
�ʫv�ũέ��dm�($I��u��v'� �^�s�`�A�E��Q�� �Ežo����q]B�)#$ș�Q�ulÝ�+T�8&�L�c�%�%.=��N�E��*�PB����������$�LU6�����(���I�H����6�@��~a-��ߎ� ���U��C��2�G`��>�1&h#+b1(�z�`]u�k5�M�a��nŪ�������o�xքELTR��o1�|����ŀ�䚛��D\sS,fjo�Cw���{�cA�;����u� ���P���~�|�����Z��q�5�;��֯Ld����RMH��s�˻ lv�� ,΁��lT �����[x�U�Y�������Ee6iQݗ�8�e��$l��F�^	��T����˛��]�;
ۙ�v�O)�m�^u�?p7{y��E�h6�ś�A, �@cS���<�f� ����A�۾� Z��f���_OF�+�I~I;o.�%z�� D�B�UM��߈��\�f��}5�z�O���/���u����r��zi���*�T�)�2�)�w\��l\v���7k"�<���杯���ݢ��T�(&b��~���A���j�	��|�U2{v,��s�R��ݻ��K��,\M��|T��"%Hd�ۿ{�ꭱz*��|����tK	$5�:%���o�\s�9Z��Mo ��WQ1J$�J��z��|�n AK��
ȕ&HG������j���5����)�:QJ�jjI�4k���뵻s�&i 2ߚ^$J:�4�I{3;��WS����OvŪNz�ƢoE[��m*D^���wV4��"�Ь������f{.vw�����r4��אE,��V{�y#ǵ��$=8c,�	A"LI&�A�5���7����jiM����{��@/�������݂����n��s�17[H��^[�Ium[!��OYթ�ͷ8m�-������>��h�UT��[j��י�0fgsw�n[{;[��U8d?c/ ,}���gm�][�aZ�`�?��p�^��Nau���muV)$��B�eSH���nIA������v����5@n/��>�4Rm�i��ngs���>3���X�o+G[��π@|l>�Q�N[~����%��g�_�r�T�xj鼎 25���@�vo]ؒK�a�����ou$���~�TR�*�(����{�v�����^!l=2/זo_P?k��f�u��$Aa���J�r�;��Xb����_8��\@��Z1_G����s���x`OdA���DF��{m�zYݡ��N�I3��Uا$���hDA:
J+\즱kq��ۚ7k
Cv��Ɯ=N#���ې��v4ۙ�U�@�k���Sv�ہ�:�)��80Wvx5ԝ�=�D�/��k<����l�+{���J�`�q���b�퓁-Ȧ���vT���-O^������:Ɦ���c��x���\�Y/T�3�7T�Bm��G����v/h��7u�M؍>���w����X��#�G.�k�[�s�����K�vۑ68��=�D���&$�'�f����J�7���H�n�a����S�c������ݙ�w`NF�J��	��Tӂ;��� e��;�6�������I���[�I����e�N�	�������L�"�UDD̕M����J� �cw|׃���xeQ�ۦ�����w� ##�[�+���_D�
�&�M���ɼ�[X�mS�� e���� a��� ����ޞ��yW��
���O��uM� V��@E���k~�	C�'�6�cV;��w�v B���d#a�y���L���L$O?#K�<�͙�������E�5n�:�Y�<ܼ�z���H�7�l�"LĉQ2��V����"��a�c���}>춽;K�wB��ۻ� ��[`�dN�T@@&LI&��5��t��yXU��Ԯ��. �{����<��B���j���ѳ�g#�����'��>�Xe�c"�i���Z���Gn<�8$sk����c���� �����}�~ +���ܟq]��jz7�p&d ���i�Ou�� ��y��{���괮턗�#{v�D����Y'ƭ!a) 7t���w����%ُ��U���� ���H���=3*9^����|��MXb��j
���!������D�n�-TK�3ṝ�Wh��y��x߈fv��&��w�Y#.��ߦpjX�� 8-��Tg�6{OS�t<�u�ƥή��v�?O�#[�P�RU��׍�� �����;w���W����@���r�۪�"�:y�0) "�jQ@��Ҝ�o��<�.1=V%��u%�Yx����w~I%�J��ׁ�2�=JQ�*$���k�� vv����ǝyV���S��_�blr�9��v9i�ݷ�o���1VD�p�"Fl�����T�G��M�N��e�R���5��
����[����GV��� �'^T��]��w~Iz��A¢!$�}""Y���㐢��eD{�q�� �޻� B��i���s��i ���%͉ӓȂ�"J��'yݸ�n�{��P���mt܀�{n� �7z�� ,���Tg��<�a�"�Pؘ�D��<��s)�u�%Գbƞ؎�.6��%�.k�7;u�:�}�#�}QS?�!ǲ��@��;V$��H��O�B7�o(]��7J >����ٮ��B��*��[��D����FA���g��g��J�w�� n�d��{�%��~���~%x�5TR����j�C����Š�ڢ�IA�k{:,]��q�5-! �7z��DB���a~R�T@O�D����qץ�;�����n��� �Qݺ��H#���>�ފ3}3�g��_�.u��_cɷ:���#]<���6g�%ul�nk��l،Y�aP4ߞ./�qPmM�a�q�? ��v�"׺7�̀M}Jf�B��m0H��/O�L<�D���w[v 	��L�'^S�-�N��}'!��ߜn5�G��r�8^����7����Pv�m�*d���cp��2
�$�
e�'5�ڰ@ [��0@ >Xu���/3��L���� �n��h��A���R�V%��7K��,B��m<�{]�"�v��� 2:���������y��M�-(S*
�)�!w�[L ��i�@9^��V����_{� ��� @|���oį.��L�32f"f(����ٻ���:� ��)*����C��Vu���޻Ᵹ����y`!Wv7�a�NxI���T�0������RW����3��a$ַM"W���oԊ	,���@=�a.DSo����m]�Ur��T���ůel;v�ؑ�u4�/c��ۣ�j�;m��Ղ�X2��4�=#�~;�}�����|kK�� ����w���?[�9�U�������!�1�dO�+eHh�6��C��u+ט��Èf�g�Oō~��;��5�'��1�#�~��8���)A[��Gi����c�J��>/�?o'�`'�����p,SW�;�<�{fO8����W���=�T��\3Q��G|'��R�u�{r�{�)�h�9�3H��"6�z��h�_�кC^�ЩZϝ�ɈB���3�k�
��x���8�#�<9���S�-C��l��Ȩ��{s�y]��w���O�n�5�����{��[��j�F^�ua�ɏE~��R�	�d9���ݩ�5d��D̓b�V����B�?�[}�#vA��ub�y��-�:6�b���w��s^�!��KA^�.�O1�\��f������x}��z������A�,�O{|�&`��������^ޓ�L�����y�`��n��^��˒Y�i�&�<����A�
o#!�vk1N���딉��7|`�TI).�%CS�{_k�-�:��X��I7�?.⧭��ԏ]^�_A��,���N3���{_�G$8�+��^���O{53��}�[����o�.K�Ή�K��:v�x<g=s�q��&�N�#%��C�+�%���/A�z���{���3����J���tD{0�nt��h�{RVr����mf��U�;�������	EE�9�pW�H�8�HT�Eh��&���R*,R���n6S�M�Ar���r	�㊰�ܹ��s�Iq�1��\�N^"\�9P�2L��k��Ç�%q*83�RyX�B^�3�1�ӷ���
AV`q̗.!Ã�N��yL�$�J���#�(��U'9�(Ң��I�MD��Q"��*.2��⻜�Hs��2�R�3p姊IŸ��9�<���-�����3+2��L��%�R�.8�"U�W��E��]P�Ey$��4Bۍ���Sˏ�T�L��IP:IT�(�����(�Ed�YTx��v�m�8s�N|pc'o .��H�d��H�[e��H�,�8�S�8*����S�l��n�NC�!�\���ʒs��GwE�(��'�qEFV�))n+�q�!�֝�q���PҢ�L��aK$�8s����U�Щ5�����.X],K�i��۞�n�����㸽��ڃ�'���n\r]9@��K�ˤy�Ob��&���<�z�r��;�,��=�ύ��u��/>š�3�騳Z�"��ջiE�=s�y��0�B���1��P�&��c<s����Gf����<��vy�V��8�8���V.2�0�:�bv�f���\q���x���^�X�&�n:�h�Xc�6���ښ��h���E���X {�Rp/�ǧr��W�8n�qq;���h�3�9�L�,��7l]�mƎy�f��bv�oT��]�7��q�p!�y�-\n��=�n�r��'�&���i��Q%�ɹ���gv�vۗ>�W����d+]=�dU�c��Apa�狮 N5��l�<,#���Ũ=ɍP�:�kk.uv;�z����yz�)�wR=��=ql��5�%�&��������iw�EOnώ۩��v���ۉ�\�-s�){Gs�:{=�5g^�Pn{�gv��1�nlu��8U�B���a��7f�>��[g���M�FK��Y:$��'4�Ć�
�{lU���������ez��kث�y�l���[nn-Z�x��32��[�۳k�9�yg�y�m���mq��dڼ�r���gfVl�-mF�Ι���Hҹ�ϭ�H�N-�%�;q�ї<��jΰOvi]y׮e�lYp&N��d�/[�;�I��k{s�����Jz��Ҥ���p�d�ȗgF7n �&T�AKЈj�w�0�;t'W���Y�j/n�nK�,(���.՗-����vfۆ���gl��f�xw%;��<\1�n;tU�gƠ�j���-��֢WI��n��縮�^7$vy���W,���̖�'99	���CGۮ�剧�;�:XM�{=B��ۜ�{)&��֏Z�ι�(�7�u۷7Eܼ��'71�kN�%�Kfډ;��r�Eʝ�m�qM��č�(�+�u�n�.7nR��5��
�Ȯ	9�6
$�ݺ��H87<��K8�̚�5uv5�\�ٞ�+�O.�Mbz�<	�n��)^�I�ܻX{va���䮞3��6q�V瓬n�<)&���m�n�{<�a����*v|*Pu2d�&pg��N�v�Vڷ��R�d�r�������Q��g�+�����|M�g�Z�N�'�X��rڰv������K�$�9�t��I(�H���A��%�N�̩i����w��Ov&��gl�����F�����}��>�Uѕ$P*$T�V�6� �����%%<j�����/���3���"*�ͪ�U��=}v)!�t�` �ʈ�)R:[�t| nos�""=^��4�M��Db|߈ Y��w`�͖�LJ
���3�׎H^�ꛪ�Y���|�� f�sv�@��g,��p��0E�����HP��$ȃ2&b"a��k��ZI$���:YݓV6�.���H5�ܒK����D��l
Kh@�ں��X�3�_И�.��J�h�P��vѣ=�EF�x�lDuف	O�J+�6��	0�xʑ&�&���� �s���` vc������*�8kN[lR$�wsv�;0p�RQ>�4�����"xR��TBԷy!��;��=z��^�žו��vf��\p�?nݏ� �v;:̣ʞ�/u�����Ђt�U@��db�U)JT)�1=��� 
������o� ��Gm�ʇ�)/O	ӊR�b%b�c�g���D�ʒI%T��]��w��ՠ$��� ���m/_�?�`)i?Z��Gz7��˶y�!L�ԧ�m�i����KVm��l���3|dD��w.��S:Z�10A,m�l�o���s^��㪟��@*���� _c�C��v�_�����?���y�Ҹ���^B�̱�m��[V�nD�C������z�ɹ8�s�~~�΋��TL�q�߷nՂ �g��}RMܳ��]L�Lv_]�~Iy��E�a�	��xʑ&r��9|ä:�Q���$�Go��	�|ؤRS}�*cS�潎��/��b�&`	��bk�
w�i0@ 跞�[���Bw~0L���N��9�$�N ��AOj���mw�����[?T�6�^���Z&��{!nD��a�U�������\8����_[i� ����,��1JR!D� L��k��'v�b.� k�6�o�L ��뼙v����ly +���f�I�F&TG�J������	���ŢhӇ,Ȍ�@%�_�@ >6-먆���wi�977^�j�S��()��qxF�q��g�ø5��gau���!=��װIؚ���'UH����"t�\[�P�A�o��%�޻���l��>Vg��,$��z�%�rL�fDʈ�����v	�rމ�XE=�/ E��~H���l��R�v�H��#������3	�"L"��_7D��fw;V�B7Q��G�c�veb l[��� ��wh/�jlA3 M}D��z7�퀌򞕸�u.������ �[��w` t_[��u+�1C�ΰUf��(���[Vi̧�tP����ޝg����`�=ٻ���!��se(wE�^Ű�����>|U��ł����IЬo�%_�EЖ�uh���6|��ٴ�K����B�Řq�e<	Q���X	.��&����}m�ID�:{]���[clv�QR �L��nض�lJ����Ob�:k�;b�o:@n�ιێ�����NB��$�J)z#w�ЀA�������}u$�ЫDQ<jM�F�vhׇiU������@D�f�H�����,����x>Y>���=>�+�: ��޻�$���}t�H�Q�E�1������ȭ6������&�p��}wa��}~k��Ez��kѮ��8_guݤ 辶׃�i砤)�(X���%�?t��~��IFy�^��� ��`c��\W��o��ܻ������5�T�z*7��� c�����Qw'Z��{[� 轶�P->nU�W>9bc�G\l�<d�+;�l��ϥvV,G������	�3f�z�P~�x���tqi��v� %��cw�v��,����^����{p�64F�����5q�v��\j�;�y�q�Ym�ۋ$�a�] Z"l"��N���n;�uڼֻ��Q���X�Y�N�:��4�R��uض��Æ������q>z.t��p�W�O����#��nG���+����[���ռ>i��G���Ӫȋp6�w�v�bDr���o��?+��>�r�OMݹ���g��LK�i<O&y�ˤ۬1�m�ƹ뱗���n�˺�y����ߛ}FM�8UUq�Vۈ���{~�` 2���ْ�U�=.�l��I��E�m���*��$7��crM#S�ݮ�k;u���F^��C�,|�!���:v^{��{ �fM��1JX����`|c擡 \�o�<d�l�ǡ�m�@2��a�"�&���eUL��d��s�k�j��I �ʫ�-$ ]r��|���]{|�fv�j�P/!ռ�a�!�"L"����}��Օ|>��F[�7`}�ߘI-�X��X���.l��)�n.���UB�3d��hp�R�n��+�]�B��R������������e6hė������` �=���nw7h=X
�P9�6�c�s�M���mW6% ''��J`�@�et�<�FAѻ�TV~?��޵��ɹ�v-1��}�;18�m*�g,g'vvP��g��ա�������o������dԑW�9�G����W�ra� ������;�w��f(������b"	�������u�������Շ� �ںw���e]��]NQI!���v QLٵR"b`&)K!s���ⶵ�De���G�s.�΀>vgu݈��]s4"�"M������L�m�<��*+�52U[�wX -�Ϟ2o�~���~K��'x���d�����m":���b7��b��0#߽ˊv6͹������k���cp2Z�+�8��фL�3�`��!1&%B9=��� ��n/�������W/;�N��;X䖕�o6M��;Q(�(��A�s�JDݣ�/�����$Ovo7~I$G]u0�A.*la2��3wb��9f
�$�2ߗM>��������	 �W�#��%� �?*���<E��1�6�ʅ�-β���ξ���~�*����uo�!b6�����ګ�����1	�b��f)�9�U�K.�+�����Z ]|ߡ�g��D��Q�f$2x�����8+�=�]�[�  ��o��o���q^&�"=U�� Tͺ��"*UL���LE�i����;۱�^]�Z [z�d |d[���(�eg�TΑS�{���n��'fFꭸ���9�3p��{s����Ԟ�s�H���0'�&!L�<��f�$m��Ia��-.M@�ξ�uf:m�r [|�am<��?D�M�M��n�I�TŘ"��[�{4��Z@$�Ix��tK	6���I�\�;"����m��}}��(&�)ShOy�� �	 UU�e׹�Eߵ����ɐd[�?U��%T�"b`�0&Y��6�s���(��I$9�y�H��z��� ����j���������\�L��Q1���a���6?W����Ŷ
�u��SMo=����~��=����G+:��0.�����=8A51J*i62���{y��ʨћ�F�$�r�]4�	6���V�o]�Kw����##�}��<�r5�:��BQ��^W׭�]�����k�ٮ�"L�&"��t��B�$7WTx$ ���? $oo]��;	�7����]����D�³o�;�3}J3)��u�6���2YO*��Yo�?� ��� =�)�,�'�K��햲cb�Շ7ḵn�i�Şi� ���X �i����������� ��o�n�u�C蝗(	A5@E*���6��"������߄��݀_[�
���;u���F��V{q�~���b��D�2��}wX| .��6A�궭�ܛ���'>t�������B���e/��Yܩ�n��e�9Q�ۤF�b��r�QϨD�X!�9F���	u���}[�1{�0�
�0�����=�K������s����f�j+6�BB��JS$[���Vg�����8����v���h���˜�nru��X��I�k�Y�լn/=`�[��e�h��5�A<��[�����a������UX�#n@谬򼽔�s͸Ix ���N����-�m�sS�$q��6.�㣷l[�0�\]S�n���u�(vN��`{���r�Ǜ���[���q�ګ�#I�f�秌��y�zc��F�gm��pU���kn�]����f�H�LbF�J��n�'7{��ZC� ����	�f�aʶ�"On�7i	kX��
!I�f��*�x%YAN�g�������z߀>.��_cl��}�W�}L��]��EgMT��f$����Ew���� �g�L�{o��ګ+�V {{���_ci��eIJ�SS(�0x_!�'�&� ��v�>�[{�� ���'�1�dDE�n�a{'NQJ	��"�y��6�L>���Y��u�=�SO�.ۿ��u�6�PWi�bT�2����/I��EDɘ@��=q۳nݶu�\i�Z7�]6�.w�o`�.�t ��!��,����D���x |�� 'k%v��g����eݠ��m���=�DAUPLR��M��mx�'������~���g�]P'�܀O����}���!_|���4���c�Q}_�c���a��0���?ZV����ʃ�Z]�i
.+{-��� ї��� ��󘆁{��f�"��|�,֪�Q5R�
��[�� ��|��}>N�<�٬��$�u�6�I�����1ئ`O�)&a2cgy�=g!�_zIA �� �^9h���w��]�?F��r@!:�m��eIJ��je���{��v��g�9:���uh ^�t�I#���K����[�o%�������ϿK�'�ʕ�S˱Χۭp�9�Χ��/f7X�v����������UTDR��Oq�� lzӣ�ww����zb�=��*��>C�u��	����:U
�f�T��ήwv��j"�}�3?{֓ �ܼr� �wz����^�s���o�a��{b)AUPLR��M��Ɲ ���ZA%�%�U;��
��3�"L*��.d-�R#����޵bƻWkZ��V��g��X1�e�ٯ��!po�K�v5A_�m�ؽ�a�š�z�<|���[�����ѓ�Z}�𸳹*g��ya��D���L�r���{�/.:��+犂���Ķu3G�/����B�%�<�ʱ��y/L�)�V9}����K�"�x����}�$Ja���L� �|�􃝠��:���/���Y�c��\|sW����P3E��m�ܒ��ɔ1�j� ��?��Ꟁ�e����j��x��x�!�
�r�҉�}f3�7��=hϏ���k��Ҥ�W��R���^��w�or��5Z�t�< ��vK<�+�mN�&���<t�C�Ln����`��E^��n���/g/W�������p`Ŏ�>��{M��tX�Άq��g��c>��y�Ӌ��=�b�8M�,��]�h�����x&��9�)9�R����|��\&,S҉�D���xP�;5��qKh�s��T�q=��Ô�w#��G%�f�8����o��`��x��=w{o<������wq
B�'`�w�=�ڧ��%���Y�i�SR��j�u��o��Nm�5��gw�ە�����}*[��24_Y�}��c��Լ[�ӯeTC��]��\�f���\'o�;�t��	�כ"�٨��>��=�p�j�	�_�{�)����z>�xh�i�e[��d��9�����o�2�����83�U�$�V�9��{׏�׶�hbVHQ)g"�!T��SRD.n'�����EJJ�'��G��9Ŭm��6�l�m�g 㳹�'d��|=�pv<x�ۗ ��Y�AYs�xK���%��:��k*��L.UT�E�<�5I%\�D�a�V�jZU!�]%+M$�P��(��JiY����mp�!*�t"%�b�"�9ĆZ���K���$�EV�΅�Ȓ��1��O]1A6F�"IA%J^$���X�
�P��9ÒHT��224L�"�*�%Id�Q[KML��\U��e-L�XS����p�Dy
̉"�J�����$�HeD��i�Yi��b�u�dNr,�D,U+�,�5�9E1j�[�2�R�W9r�BIUi\�EHPӥ�I��i+L�6el�q.1�d�2M:�q�<x�ժ�`��-���"Yd�Zjy�ܥ�"����� ���uy�r ��>mQ��n�,��T@S3&h�β��.ы�`Iy&�uCH�;�z��I$G_e]�@;����zE8���ǵ�A��N�U*����TId����Z%��e?4ͩN�����䐊�n	%��޻�$JC����b�Q���o����q�������曅f�[At�e���i���q����7�����~:�I�k��}�h����GE�z�*�q�Qs��{'��� ;{z��<i�`%d�"Y��U��E!+"���{�,�n��wo]� ����R�ڞ1�}
����"ql��#�L���Tٵ���	F�y� [kO���]@�޸&�Wۼݤ�^�f6��g�"�J��Q3I������u4zs�؈�~�z��ٞ���K�-_=<�10h�9��;�^m+�s/�[�Ȟ��S�={;%#��e�L`A	�s���]۶[Y3��""*�����-�S28�׷v��%�Ȣ�Q4(B�p�6=x�v_4�aI�\��o������v@#cs�	#����UF��5�I��Ag��u�m��ڥV�/Y�]����7iL7\�p����~�"�@�E������BI?���A��^ˋ���\�{e�d��q���+���iB����(�M����y׽隿ss��vynv�;�@ ����/��0�;���8�~��f� {,�(%UDE*m;�� ���n� ����Z��+���� ��u�e�P*��j��	�*��{��FD���O�#���z�� J�o�0�9���j�E��Iq��%�v���R�b�L�l9���@����{��鷁����Q#,�� �����p��C9&{&*P�jh�Ea�S�3��)0�MJ��|��㼤\��w��=���F�o��AΓ�^Lu���,�7|7z���"� �"Y�^�ټ�9ls�m٭�N��o3۶��rP���n:��0���s��]j�rP6�룮f.7��j2:W,h�!nV��ۖwr���q�ٵ��]���zal	�۴=3�3a!�����V�Cs�Ʈ�ű���饞xƇ'7h@��K8�x�ٜu�m���-�.6�k/6�l�xy�k�v�.m<[9��+��n�c����N8��dN���㣷d���3�r�e��<O7,'�J��LE�-�*`J�@�&t�e�p^ �i��	v�7ђ�g�k��2;-��@:���>��"h�I
IE��޻�K#Y���r��b��Rq}wu͂A>����I���L��W�S�%�Z�G��e�a�s�z����T]��us����%��L��ަEq�"�0�2I�4�}��g\���Ę��l	�w� �=�H}J��P����"n�L�$��()�-�.�m�q̺��m���e��wsz��"�~'ǎ�Г|̕t��GN��Lݜ?s�]���]3us�Lv��svkf݇�[�.b�ם����w��\M�u����+�����|�|��Ӧ��G�=�߉�����Q�TĘ� �"[<j�+��QӲ��.ߦc���0S��:U����h�����Aڊ�ˉ��gs!R]�A�|VY��A�6bu3AÂ��*�=q�ۼF,������>�w����t�m�v�"'Lv����ĩ�d�EV���n�I��OV��Gm�I�w�� ~B󓟉+/�@Dw���`ճǖDx�w�L	�۸�A6���Ȼ�N��� �fW^�B,�!( �@�ݪ��N��a��}3�p�L�A÷p(�}|�J�'�)ORF�+�.ɥ˸�l���I�@�l�6u�ܸ:n+ȗ![��	�O�A+qO�~��������6���cxvj�݈��ִ���	�]�jx�bB�RD�k�'�6o��9�[Y+r�	� �Yw���̀ ���oOgC�����&��QZ��B-�5yR	�w͟޽��M������
҅����PG��YqYʘ^�j�vY5�ރ���N���G�EJ��H?�i�_��NXy���0�7WO��g.�}o���E��`̂A�2
B����z�ZY��d�щ���I���l�N��;�1}�Q�Is�^ɮȈ�D�*BJ`�y|����0q�]:�sR|N���'�:�i�A�����M!3���{���B;�u ��F@aͬ��f�=u����WmU�������ls���߉�L��Q �����@9�z� �����Nޣ���0ɷu�:�����n�����ڿ6������;Q��뼦<GfoS� �*�;+yK�-;���x>�� ����"XH�s^��ssz��%7����㼍�hɧa�F�	�x�'ݙ��#�\F���@5<��/����eo�7m�A$���a��t�Z�Ս޺7�Go�4���B�d^�r�`E=�y�qϻ����T��z�.MZp�^j�v�}�wJ-��y[�w���<>T�"Q)
����A�õt'��@��3���#�7��H'�L�����x���������,��{�;�٦�n<cuƈ��sc��N]��0L��舒L�R�%0s�-��g�n�u0H �S�v�k�n-�˜ro_�����K�(�H��	�4h��zI��DK�G�R�ڬ$���lA�;u �CΝ�����*�l�$LD�AL	���� �3�	=yjaR�]�~$���a�F�۩>8��2ȔL�Q��ۀrA�b��{;r� �N��$�|���ͧ}RA5z�>ڛ��3b���l�Ǖ �v��ӷ�ӮKOu���LM�ܩ��o�65��)b���!�w�ۙ/Af=�%Hfe^���PBҹV�?:�3�_{�p�ǭvy�N�d�w�@�ڡ�t�$~|�����.��-�٤�l�iD�m�śq�T�	;sѮ+�SeaDrbN��(��W��rB��W�����fz��ٛjIyvS���C ��nݖz�r;]ûo���wN��e{v�.�������&EێN�c;U�n�gb�t\�=g2v���]q�l�km�0�hݲb����giN1t @���G��๹�O*]�s�rq���%��U�h���:en��f��]r-7f& �y ���}����DJ%!�}\�$�3�@I� �|��睅�=��]�(`#L�P�[
$�&0��`�|��&�:{v$E]��׮��	�2(�F=|�&cc��=J��]��a�$DB�Ț��$�u���� �����j!�O�۩��_0�v�%"&"T ������Q�wQ�r�09@I$�x��K��y���\N�/A �o������fA�fB��Gkwd��7���5��� �Nvy���I!��6GrS'������A���7��6��G����9�tgM�v!�ѓ�
�u;�"n������ޘ^�����g+(I �n�0�$�}����#M��;y���@H ��f7�E��T((��ۮl�\O�PM��ɰu)���?{���{{��]� �{+�r�s��:�EZ6h�?n{���k�VY!'��}^���tS�Q�Et�;gf�9��
��B2�}$��f�$�}���S���cN�,I��p`H�"RP����l�O���I>3|T蓗�wu4�I�Y��A>w����f�#"DHF�+�k����:
IU���I��l�	���3X��Qm؋����l���)1��N#��$��r�tOcTBV#���z���0���Ԫ�}�X�
#Ѕ�*��=(�;=]g�y�j󣭺x���k�m�e�tJs�n� ̓!B�
}Q��2{���$��z�r�-�^Xu,t䇷�͐|�7�'.n"4LL(�!R��� �u�S9��gl:�2	�$<���$��z�`�̎�����?Ff�A#J��$�+:�$�>#��A����CQ6�Nu��/�V/w�;NHB���-t�{�(��v��m`�1�dU4 ��ۋ%;���{[yGsoO^�yUS��}����	��ץ�k���R%(���`���nr33�0���I���`�A8�r(I�]�y�m�IɛB6v��I��L0D�P�B0&��u��{r�����]�7�	�=���[͑�/yK��+��֊F"b�\8� �Ln��m�u=s:s�=r�n^�[���O���]�(���/�n�d�A�9�$�q��g&��ꞓ��;���z�>��+(	>6ֲd)$#aH���l2su��yq��a�m���V	 �]Y>����q�.�,MGs����(�))��(B�Ι̊� �w͟�]ъ�5��֒F��o������0I��JB�ݾn��M�<�����7�BI �o1�|H���~��0��~�|�\du�S��=6�_3������ټ΂���<�ք �d���`�{4�[�qH1n~��ʼDt_\$*"
R�^�?e��?��݃%(�خM�	��a���ec����C�4�3JFjߏ�.�9�k�'7:<!�qmp`��n�Lp�_����#A
B���K��$���2���`\�E��0I�����?�Rm+tIQ$ɘ�-��͒ssj�X+Y�LvܒA>m�6	$]�s`�̝�� X�55^+U�`)'��"��Ͷ�$��u?I=���X��Ǜo�����oю�I�@R�TW�Q�Y��Ӿ��s{����`0I���i�Òy���|j�=���a�r9`�(���|߉$����סּu�;UӒ����:��r�����<QG����g_�m�o�0m�o��6����c�l`����m�lc��p6�����6��`�6���0m����0m��l`�}��0m�6�����m�\c���6���pm�o�`�6����0m��������m��
�2��h�P 6V�������?�����<�|�  @  
      @                     p 3�UT ��*TzhHT�U*B�(�PE B��J��J�H�(U�E@(����                                        ���P0�}+ˮc��r�6�&�H`��
�v�F�n��Zs�J����F ��G-v`S���p����  y��0�C�su�V�Yx &T���=4r5um6�jDNۭR��p F��.���=�6jsu�m{�ͫڊ�$�U�  � �       ^���9aU�k�����mfӡ�����S#u�E�[�i�t���׻�oT� ������ y�< z ��   B���z���� ht�� ҂����N�^Y@{� )�����'� x�v�:(6��tQy� 9��z� ��
J��  � �      ��@n��zP7�s�ް�(<�;�{�� ��%��0�s�A{t�{=�*��� .��rw2�s�(���|  ��ﻀ:��Ep v��[��2YN#N��U5u�!S����rna������na��)TR� /�  �     =  p����b�s�+[��C�u���p pl��� �;P9V�WB�� 04ZΊҮa���U6�E�  ;Uy��T��g �N�3�t�vr��E� �u[����@�1����5((P�  �    =   �i�;u��sk�#�(:M����$�`������ �֋nF*���P� _|  z�� j��ց�� ��r;��)�P����:��:7 qv��;�&ΝUͭ��
.�˥ul��  P  ��2R��b &@ 4�C �b*�	%*R� &�L L&����UJ�~��R b   4  ��E4�Q �     e) STѦ��� 4  !!��Bi�i��2A��xD���}>��}�}�o�5���$��.�������L�?�		�H�����$ K�?��� ��@$	RH��3�G� BB�x�������'�O�a��C��������.v��om��`��gc�m�����6;�*����h�HH@�����ԝ�}�4��}ߗ��_E����	r�r�"�)���G���G�/������|�"�CI�s�����j{v��j��$�6M��
�[?�xު�&�6�v,W��3���#��1a"�F^�N�n�UD�%�V�0>�fMigj	�n��G��뗢�f�˞�雌cI1Np��1f�Ŕ�ov�격9h�~������6:b3�8��t;�>��hC�[S��v�/0��5�mͯ;H	� ������{ �͆�\It>�Ӹ�<-l\y��#^�gf��ƹnٜk
@�wXZeя_�Ό=��Xɓ�9�ئބX.�zb�˯� ]Յ�M\�X�w�˒��J%J�5�:v�p�g;xK!��s��ӖY;�H�.喻�����)BɫQ!��r��O�9n���O++�%7v���ʜJ>�'nq+��^I�����bA�t� y�ѲW����F�����P(����ԁΛ����ŧ:d6R!�-"r14�8L2rG��%���NR֬�-4,&Rס�����ǶIh�q郡zݡ��I�c�����l�gz'�foN���ɬw^�
&�4[�4q�]��kv#3�"ƕ�B�pm�60ZƳlu�;�f�aȒ���ۣ݊f`��&��㑕0��yU����ȴ��3]�F�֚��a�Tmq�e��LҔ�f�
�޽��nTY�0�7�{�S�����.��X#���{�\ق��q��0��{zoZ�!;��׹�4O�Yn��N�۶����]�nǩ����7�4�!;���F��yBcW7ߣBD���:�{���f���\007ua�ٺ��/7�hLb �r�tܥ�m����xv;�	8s(��;K{��c�n�؞.�V�&�.�yo��$���`�X�sN.��8:]W��r����;ӭ[b�3�i��+�ӈ��B��;)���_�w']��N����#����PO���K�.vWF.;�k͉kԃ����97-�(kG#�wZ��];��V<z�=�~�t��ʚ[��-2I8�<�%X]�emz�]�+��FI�c��D�v�uR<�O�ڛ̂ԍO� ��>��w.�t�6pF���ib��B=��ъ�8�d�x� �.?�o1���M׋�����M���-���v��;�jF �W/<H\������0�c��ۧF�pO����;��G}.=��r,'��^ �B<6�.���m"���a�7�]��Ą��	jN3kW$*v��pdn���d�}P}A!�̣f��#�2n53�=�w��)���w�s��{�8X1l�v>Ĵ��IM��Z��
x]o:)W\���`;�{6 �HS�o,�F��t�9�Yͧ �5�t����@�G���o��ua�Ss.����@�mF������v�&��!�K�{����q#�b�Wr���;�ԤФ���[���İY֐EX�s�lŦ�Z9�XR�$v,��Y�j�%F��zk�:�Yz�gr�6,,�=������!��:qW���lWKk4n�9\����ڔ�hm��;7�(�=�zH������c�[�k�!*�^��o3�F�����	P;m�� �Y���'��4����?Jt�V�v��z�onm�r����6����m�<>�X�2����nz��{n졆9�f���U`����j�������d�໳#I���Rrc9 ��7���!�
�f�]���plo�#,�2�+
�s��8��3{qaE��h�k_�z�^���s�&8��\�p�p�X:�.��x��9)�Z�4�?n�ۚz�p��2�t��"��Cf��
:�[��s'BG �V�w�,���vl�㯌�`�igwc��,X^A��#�2e�+<�H�&j[KxsuE�)�M�v�H]�d�lW' �9��oN<gv���#9	�U�UpA?�;��r	�Z�\�������}��[2�!縳x�-/��N�n�iQ09�GM��y���G��V��gr���y���vUj��!ؕ	�N٨]];�E�b������ڲF���=��I�qk���31v��ųa�М�[����$�h]�w��EJL/&���׆�3��p=�K��{����j��\�Ç�<^cl޷�Z9�@���mw����p�l��Y<.5�dnvA7eب�h�^R�]��������P�����<7�~�����3FòjV��^��1S�7�P�E홳����id�f(/���/u8��=���'�ǗJ�=5i:��lk{y����H:S��$�P�Q5�min!q��&���.:�n_���y�j��95�y��X�N"���{b�N0��2�Y���yS�T���a�oA����e���
;J�D_�P��_�Y�t,R�nVV���٠�#�z9������wf�A��1���ݑbҚ�j\n��;o�1؍�K����Jv���	N(u��8�v��N��V��xfVx}��sǲ���Y
5	��׵���o�D�y��x��q��4�8us���6D0�I��]�u�[sp�5���Q���%n��O[�<�=vmC]���{u�8B�9aXn������#�m�>Y(��G�gd2#��t)��zq�����h��vj� ^���5٣v���v�3ED�Hr���,����5�ÕU�x�K9!�3��{��f��y��%��uɭf��w��-���&��B�U�wz,]�!#Q%e7@�4�n^Ca�z~�a��x�pݣ.4y�����j�J�b2cW�oo�V��l/�B�w�3�r�Tv�rM�NC�v%n�mKX����F����g��&�V���aܫX��,63Pw;�2�c¸^Ŵ�B�ᐎ�5�'Df�i-�0ҏ���(i�9��h�D�y�3���*���p�T�u���������V��g;ؑZ�};Jy���!-��4�[ڦm̼4�שa9�s���B�09����l�
kc��}�F]�;9�G;WqVsK;c6f�T�i�y�B��eY���}�x����o��,Xe���1�+)���<wt>
����=ʫ��sn���%�ػ�M�	좥E�^v_�Y��4� ʱC���+SGk��u�b�^�ʢ���c@tK@`����<��7q�N5���T�[�W�by�64nE�]p��w�97�Q����ʃ�˖�Q�T���F�H���u�v�� ��<��j-�r���(�<�9����`ǧGkj�n&���3��;6�J�e=&n�]˹�������֭�Ʃ��g,�»����p�E�%�)nF��gN��I\.un��C��طr�翲�{{��9hwp�ލ'����b@-��^����Xp�hR�N$��&�T�gw[�{��LA	�8��T�y���{� ���p�.�l -�vJ������`�p���������mݘw#��{^�k*�m>Ѫ�
�a��6�tNXs9L��ݤ%Jh��sm�>�̓4�ͦ��v�6j�v�3v��AdճZ�{z���e�Ä_ݍI��Z��f�ǝ�mRN�u�L��K@'���/�	^�)f��e���:��9f�jyӪ�"��l=b�ծ�c���XY��
�N.)��� U�����:?Wõ5�5˷KwyvS�4-;��ڄ�qQf�n�»:�,� �H�峃:pTs�~)�m�BX�=�����u��>�^-i�ׂ׆(�Oe�Rh�#���f�����/TU^��2�����Xbm$���_=�pdѯ ��:���}��.�Ŝ���)�<� ŀ�n�)�V��L�Ă�u�.�m{L�#��$�%�.v�a���ئo<��Tu���S
�}����SXZl�V��o5��F���gn9�z^��vq�0��]�S�HǗ'��U��۹ͼ����L.�f���s{��}��v�#&�56�hTN
�����P͓xG�I�5��t�i��\gb�ob�+�ApG֌bv+�� �@<�8��2-e�Ś�j���������bo�'���P��ׅݍptD��4�ğ��'�C��t�wzf�*��#��F:t�ɝs5%��b�{�A#�F���㬵��:.\F�ݳ��xJ�+αdp�y�ݭ����8;6f�fp��"�9#Hlr��<E�EH!���+�nl��pbT�T�Yf����+K6n�n���ͷ'jm�]y�����+&�ŗ�v��sN�"��e��1���9cٰ&��A~�:B{6�,�#�9U4�_QќZ�����s�V���:�yJ)��ԳyW����7!�x�rl��\�p�;�����N�4Qf��؀8�>ܺ�::�=��*n�#$;F�k���3��n��2`B/.Q�NAݬP��׭uSI$>G���.f��v�3�z]�{9vH�f����34��MP���鿖�7���㯅4j����X��ł�����zȲ@�Y����)���7��B�� �	�9�+c�U�5m��7�:Qq��wu���=ٮfhO�+Gj����eΛf���2?3���`��K�'[�v��>�(!�1�7���a;9��N�Cm����t��r�@���7�XPǷ�|IW�F�r�{Nsy: �@:�4X�)J�:����6'���{���m)����6���=ܸ�(���\�q���%��OqwGp�B7s�ųv�=�u����Aىt�Q���fC�r��EzJ�'s���Okq��3���@�H�(UkKV��ÍOۋ; cvod�_���,�W���G �e�tkGf<�;;t�l���f��ު́�;Zr��0:j���fH�^���m�ȳc�7���	���7����k�/M�vT�Ba������|[���@�1�}�yC}ϗX��{j +�&�6)t͏v�ȶ�;�t<�yH�ؿopͣjt*U���f=ݭlG���������8��w)�2B���kǏ9Z����=����i�VH��<����'Y��yٱ2�L�Ù��1P�����$���t���:�K�p��IL�8u�Xv��~�`����r��%���ш�y�(I�:�ӂ���`�S��pܘ����EĜP�]�k�#'r����5a�;K�����4���q��1uU/�ö �h}�tD;�d fj��	��L�xX�����` �M �>���KS;z�v�N��VLE��c�T��K���cΧ^�gb�ӵŒ\�Fp��Ve�ж!2�ӡk:��Uܝ��k;z-쳚	r�r�^����"&�e�3��
s�$iդ�-;�+��e�T?G����é|{N�{}	�i�fm�����(�ئ�d�a���=��7�s��M��<���� d�u����˵�Is�T�(R�͏�ΦnK)�&����%�����AT��3`��p��:�NvV�ܽ	!��t˻Ɯ�[� ë ��Zs]���F
���\/1�^�am]�ۚ����t�6��bװC[c��B�^t�u��ݓ�W6�pŏr��3��LWS��飌;�Z��.3H������N��#3fc|�qu?���&� �9�vo>٢��Q����0+��i��������\�oV̻�l���۷�#k�Uےs9{wV��t���цR;Q��sxk͈^bƄδ�V���!�I�]O6Q:肱�n�ܘ�:
��Xά��U~�=1�Zs��OHh�&4���"��9d�׺/Ogp�SA�}v󽫦?�?�á)�t
 �5��C^�y��l�%�dy�;h}:zg*���~"q{��.ǯ�v��6���:3׺�չ��0��o��ݺy�(s��D]|]6rT۠^ֻp��`-n�c-nv>��v�<��wR�]8䛋��,<{
���<�oLc��R�é�6f˝,��E&5ݵh�N���Z�Y�n��H�J�{�<E��n�#�k�1@� |�Q6A9�y�M�l�`�S&�����G"���h��1s%k��v͓���r��@Gt�U�UY0�լhXo�'$l]��XY�ɶ'��f:�V4U��$1�sp��n��@F��1vh���=L���I ��M�7�-��@#�#�cG� ~C+���`��0��0�����](�������sFu�"<?,��m��Cm�6�v� 1��q�P1 c;le�6\Sce��
ll�)��.�6P2�ě��e�.����$�	�\`�S��6�`�q�؜'ˌm�1�)���& 	e�@'����m��C���P ')���4�.�l�Sc)��c �]�bv�m&����(`l`˔
l
c`\�q��Cce�l
�� 'm�I���1�SHl .��`Ӎ�)�pe0aC!�	`]�\�` \li����eC`P�ebp!F�_��������}>�����}>FG?�!B��G��k�X׮�$ K�>)K�H����5�A`@$ K�?p���tO��c���<�����^�n��l�4�cw���x�0=W��ǲC��T�^X[�:��l�"R2"�M'v��:���Nc!ӎ�nM
�o���/�&�hwKbC��kT�J{��åWS �(Fh֬L��n͜R��e�IM�]*���#Ð7u;���aLk��`s��E�����1ۼڝ.�8͈����ٳ�FX^6��{��C�.0�su���O.o7!%��U	����$�^a�5̌��3�X�B%�A���u7�e�c���e	LU*�2����s��� �r�~�����,��,Ά��KZ�d�X'U�ڽ��7;�vms�
�97�=)���`f�Y��s��Vv}�����Ǜ��&eR�-��@Nx1��\J��{w�V��W)X�,M+�b��c6�\�F��@f�j�!��^�Y�4[{�:���	q��ݞDg��^�/D�|����vz 3�c)ni�5���
x][;�)����湴"fXtBx�{�P���~� 8#>�V�˹���^v�h2�)Lz���$��pn��2��{d�[��xg������i8�"B=	;��X�������Cj�T�/6��5#7�<B�{��p_<��e!��VHw϶v^�[%�P^��i��H'-�����*��T���Ķ��;ܽ/z����gt��>Q�@�Iw�v�w��yf�>��r��gm�!*_i��,���w���	/��ɹ'�I�8*-�ɝ����
]�p񫣹H7 �_i�\�6��{O����z�k���q�/N�o�٨��h���*�s@Rh��g���Q5d�u]���������z�yl�L!�x:��y�z{n3x��=�Შt�X��T��4�G']m`��	ۭM��QU�6����3t��r��nn�ᐡ�6٧��v2�W��4[�ؐf�����K�74;��b]�y�=T�iC�ɦ�
��Yami�)=6�V��^����c峷7NO;Vb>a�EQ�wWp��tٜ=�5u<�{	�������ȣ5/`v=�8���|r���x2��s�:E����yQ������꤄l�o�׹�ٚ6�٩͑��;���Ե�#�5pZ�V�ǯ���2N]�#��M�oT��:L�
��o��v�eV�:���ة
�R��)D�V��:�J>��{�����烆Sg��^��)��ܹ��/j��)2��(�(F9����ǒ��O���o%m�?���ь[��Ld�z���xe~��A�*�O�g�o'!��=ǌ\��z]E�>����.��ա�7����
��^{)�*��Q7E}�N�;<-�A�nO~��x*IR3V���}G����hG����&n��tpbm,�ub}y��iG��B^�O@3����n���+)�h�R��m���y��2p[��� �#����.s�h���]���:��\�t�|��x�&�N�[���AiۅhM�o(��Nk�fB��xa4Z�㴒�ڡw'��n*�����l��^FQ�ck�0�/���׳�Eay���ѷ��#Mx��ì���2*s�Z�Cf��&/R%��[ӷ���3ZIiRx,�#�9L�p��@"����z�z�x������Y]������<���n�ӭ�v�=��l�?@'�=�4������➏ݺ�A��<���Lр��_O��0зF�L�VXv���9ց�*�u/nj��L����ތ+h�7pnf��"�4�L?aeQ��u�j����� �G��¹KI���Zb��A���<�e�H9u����^Ş�t��Z��z�V�~�D�OS�a�0���_a;Aכ��Z���͛��nAv��&+p6iD*�cO��K��k��=��q���=��6�����CCZ4]�t���2���w=w��η���Z�N�^�tk�c}�z�����>����v^s��qoL���dN}j=&zx�Z��탐���zvC�o��5	O{�f]�{�y�9nX=g���q� X����+γ&�'��#���m��L�tYR�=E�e칟n�E�ɱ�U��叅����(�Fx���F'<VvMe���Jc>^�|��q���2ܽ�A�i�T�+οZ0��v,��Ϭ;�J0��8��7`ȡSV�(�)���o�{�U�N�y�׵�NY��4M��Zܪn ����l��5Vqɋ��f��[ƞ�>랂#<�-�/&���2������޸0y.;lW��x��d��������ijٌڨ�%�6[ߗA}������3�6�ȬLl:�	�63C����}p�q�hOh�;9Zf�DU)��d��A���$b�E�D˸�F�EAxc΍N�1;T�0�眼xV�<���P�[���s�	�'��t��;��Q��z+$ʷ��s�P�Hr������؜��iAT��`��_Q��GՆߝ�K�*�)�nrsV�EVX����2p@k�1�~�F��׽���y�Q���H���BJ���}�ú�NC���~���k��vM�~���\6����1<��;7�l�����IoqdH�C#-Y�t��	�&�\|��lɳ/���+�=O�|A�\��$���F���'�{�{MD@��m�mk;e-.i��H���y�J˪ʰ�9�v2�;ctj差a��8�ݺε7�.�X��������L�����k+�<����{�q��J�7�}�����}�z��n�	@#vѩ�T��j$���N�\���p�ki�/H��w���V�w�mwh�v ����k���|W�X.>Ľ�9KړǷ98�vL����Q��݉���i^!���{v��aLd�wW�V���{�{�{%���5T��Cu]��0��_[�%T�k�|�u�x���ݔq�s���ZCb�`V^ҋ�V��~�\����}9��'�/;��TX�!H��Q�&�\S�vY��B�ԃd�;ݥ���>�1����M��s���S�yCe��$C�y�z���s���4���U����{n�U�W�O��u _D��]�1�쿐���/N�v��=R8�Fu�x�\Sphҋǻ�H|�mN%�C�I�=ux�k2��+ ^W������ݾ�������Kb�����Z��}�r�U p�;}"�G������@ wfݘ���<T��;�Ѻ^�Rh-�kv�FN�:p]�o]�_�2NA�����m��f�ѷ��Ѹb�i��L�E����I��3�-��Yp���h��S�&�1u���ǟ��΂{�ǰ��qm{�=�{���ҧ���g�����Eex��.����y0�)V���Y+�-�~��ѳ���g�����jT슙��#;�V<T�EJ��8r�sY��}�n���x��ŋ�L�M�L��J��}e�e��c���֍W}�{���;ɯ0'ox>�t�_E5��@ݺv�+p��Qdը��U���Vw�����.�f\ܣ������_@kɯ��Rd:��j��o��'p��.���t���15���j�Rc�k=�UdK˯�ɲ���4�U�:��ff�Ǽ�7�E��u����c݈�gi������g�Hs�=作 n�b����]�l$�9ǚ4����19�§e;<���M�K�(ͅ�i�����_w��� ���8�i�C1��9�^73���K��m�:0z7g�%��MJo{���ɡ׆w���V���~+�X�I� �4��i�k�g���r�����,y�w�4o�u������b�D)r7O[�h���9�r����pޗ:�uM��6���(�t#5��F����&�t��ǁ��Gy��>�=�z
�w���-�s��'��M���`$���r<���r��jE��:��K��-a�ک-n���#�Xp�{/Q9M���1-�b*\�^'�Jd����wO'%jbZ=@��ޛ|�vU&�$�&�R�-�2�M���@������V�}���8���N�k���γl�}nJ]na�����&PI��*���3�{�Ǯf�ax��N���7[Q� #/f��y�,�[�z�N�z쌽�A��x�7�r��zVMy�l�'��zG�B��|ԯ=�s���g���s��/
��Y�d��w�D��:��O,���E�lcz��gU�u$;��;U�2Y�i"������Y�?^#����
�gX���J�..Xu�a�l;^%7�o%�S82��K>[������g�񺅹F���El��=fn,��3�|.s���(�-��;�:��o��0iscM���,�����H���HC�9ywwnQ&����=�n����v��G�o���a�8��%����M�36�Wr�{����;�������.�;P�^J��ؖ�����QL$�X1j��L把w$׳���*o{���̘��~һ4S����c�m?j�'�L�I��wa�{�t�g_gf�{��8�K(�U�I�ҾcY�@�nA�7���Rǲ�aZr{_�>}�D�c�BQ���b���{��]�z�bRdD41ǜ�b\�9"��$��A�<��{��� f�|*��Di�_��K��Vj#߀����5�y�s|r"�����׹�6�bEϚ��z����ꏣ�%d�G����N��=��"�
<�s���<8Y�q�d�`��	�����}c�>�������b u��BVY&���}�G��<�����*��g=#N
)�iK$[: '�#%D�UJ㛚3�
ҳ�2��%���QC�9d�J�{^��1VŤ�U�[5S+%���*P$\���eA�>�W�{O��=g��"j�2P��f�ja�0���0�c!K8����A��V�X~����LAY��=��i¼3p�8����}�����;g���@���)=^�>��� T��v����ȳ��k�+̴���i�[�BQt�9�-�ai��0F݂�[�P�bYՑCD�u�M�[���^V;q�Q=���t��Z�V�r�s=/��{��չgq/�uw[��}�8�d�{0#�o�F��yW.��y#'$�U��Le��˷Hכf�{�7�z�jW�*��]2���c�[���_����%�y�;߶6or����L^ڹ,���8}���8�W�����-ۨ�A��9�+!��=���<$����ī��4%�n{\d��y�u��֜���F�?�uޛ�kV�����6�nM][E�I�SL%{�[��j�����79�q(,�*:;s�wikQ�zt���n����^���G������NԞ@��q�`Lj��Ĩ�;^�^��^�;K���g��=8#�g"�
u5:˴�ȴ.IJФ�PLfM�z����J���7�U8%�����fh��U��.�R��1DM=]z�s�JJ�ޥ�o��[�ƞG�y�g:L(�h���9�]���$I�nN�杋E���E9KL�pn-���ѓk-�H���"��7}���e~Ōu�s�w
���xtW�{�����knm�ݝ��ʴӃojn\����xvMnV"�j�V�F��*^�Y.��|b6_�`/b�,��f��(�Ww)�؇�l}�b>����Ț���;V-�Q���Y��&���Uk��i���\�(g�x�6���^&d���]��Iއr�&/@���hy�6S�����+��v��g��/�w��V��*m)+	�{9�)'�R��f��V�JW;���	��71�P�cݓq���j7a �TѾ�Ʒg��ʘ�h��m^�o�{�n�:h��@��gM[�!;٨z�f"���vɣq�ۺz��;�=|z�$9$�qw�v����.g�c;Ӌ��~�f�^ӱ���goL�����mc�jH�� X�7{W7=��$�zy���[%pwi�=���S�u̞��Ln���7�jK�ab�Ҝy>�p�! ��i��{OA;}�8N�ܾ���2� ��rwt�2��+�do{_?.%-�6�Wn���ڕ�o�cy�o(9kՇ��Ȱ��������ۭ�yЈK(�R�G��0y'C��{/�۰>��r�᚞r�2;9���a�zu�6����ߎ�5M1�K0�Qn�w����uR�-Jk�Y����X���w}����� ����XNl=�n���w�����3[&�-12�W19�X�++N(Fe$՛t�M3����Փ���cm[����=2��T�7KF�B��37Bzs~}N��oö�<��V1�K�{��{
;����`3��ˎX/Y���c��W�^s��YU`z*��x�W���c��b��ǽK{�5�|䐐� �e\;�0{m��K�b<��� ��%���^��1�c�*�����������Z������������������������������Z������������������������������Z����������������y�7]p�Fڍ:���A׌���n�;^Ƽ�ʛ�9Pwm���K��痞�ؓ���n�g��2��X�zn��Ɲu�ͬ�T;un���:���:���L�˷=��ql��=���JbwmΌJ�'Y�vp�Jm��l�u8v�컘<);V�.��Ux��	�ۈ��l4t�a��&%����q��F���:`5�凵������A�m\��Şx�r�э��\�eK�뭺j�v^�m�OV���Wm����yv�z�&����i�fz�G2Y��.�]D�����u�c�n�N���9��1Ǒ��V��c�ݸ��m^���fLǣ��0�����b6۔�Қ�k�.����n����n�xN���ܘ����F�s�h3��K�CjS�7oN�GZ8�y��Vo�n}��6�Z�j��[��n#k�yRٻ����]]�'������	�"#��w!���u�7nR�t���˺7���n�&K��N��\�����X�طnNn[Ub�W]X���r���9�=��g�Fw�����sK�rۣv:=�V磍۷V;F�a����o=�Y��C ��Wқ��n�ɭg���gh��Z|g����vN�;��v����@B��>�7IY�"��N�Gj��n�q+:,r�@Qλt���{1�{��56c������m�;�G�ݘ\�;��b�N1�n�]��gY�<���Sg<�<���铓������^SKj���N�+;�;nN@��n|O���\%M%��e܏l�熊k�Yj���e,���,Yz���NҞ�x�C�����3��l�Ӝ�N��1�F�V"I�=�]�s�Y��4U��B�]�
�y��am����P�bRx�Y5�F�&��:��t�yC1na8�I�� �q�ۮ�^㞍V�]���m�ڞz�u��CE[�t���S�Z�܏3�5�x�ãcj��ӡ�g��۩��n{�d�����<��4v<o/m��ܚJW��g)`���A˹�99q����Nu�6m9�R�@n�۶�rն�d�F6
@�^����$G����9�%�`��;1���]u�+�vvz�;����q���yv���f�ٝi:�a�:6�����`d��'\g��<-/���̜����[��V1��vc�ȶV%�rGV��<ɷi�ݰ��eG��˒z�=�/T��m��s�D�XN�=��s �Ӳv�/l]�#��éka9�F�:��t����\/@qˡ\=�`y�x��v�(78{&Ǝ��rsܻq�g���O��-��GCrl�Sl����\�2"��b4�<��u�*�s��<��{v�3�b�\k��)�8��i���ez:�n'%<��e�ηt�؞}��LA�u�X���/Oe{]\�b9xAre���;3�u�s׍�=k��ƹ-vxeN�/k8���[���y����Dݺ1ι!�]��\��۱���xsv��ޣ�Mgim�.��;ZNM<����:��8�κ8�,���nل�#��^���,'���x�^�μ�s��i����<�u�ٻq���)���=�'�)� z�-%��fp�+���sbn���z�n|��Ƹ��pGfݯ&���"rY,=�/kO ���|/;�=�D��-Ōrɺy۷'��s��f��Kq�=�M�����X������������mp��,� ؽV���n��oq�g��LYb{�z��'��1׍�e�����q�z�^xۓs�uS˻c����z뛭�o=x�fE��[��ͷXޅ;	쵷6R���;^��`�g��o=K���-�9��Q;:�L3�v���ƚ��6ɷ�tM�u�`��-�x�㗓D��^�3؂�	��S� ke���q�FD��[�Ne1�l�#��7g���DdR�9�㧱���A�*F��.x|Ÿ�n 8�l\��n��a1�W��l6v��lS<�zF��qe.���nYƭ�%"�m�k���n��9��p�F�	;�v�٠���v@F�!��\c���'��=��n�kn����m2Z�u�Mk˶�8�ob�L;ڻY�X�ϭ���8{m���1��ۣ,<��ջ�;n�� g��v��N�l�װ=r�7��0�$nec&��d�;u�ax�N��Q؊x6Y�"��q��S퓷:}�����2�� {�WlƗnG���Zu�qv�/m�-���gu�KV*9v6๳@�k�7"Mi�%�pr�B>U�Q��.�#x��m]��/2��;�{����%�w8���7_n.}m�SWq�g�����Ş���<u@��;@rt��l�ػk��q�J�ۨ�(��f��u�4�&e�ȝ�ۅ7=��F�N�6�ҹi]���zs���\^�=1؆RpǤ�m�zS�n�e�,y<�V]]����-+�"�ݭ�\�u�ۇ��{um�;x�ۤ�q�r���9'V�d����[a�]s�6��+s�Xq<򻕖'\��Z�屦$�r�:�A�g l�Oge5�󶋩�wl nL����g�9��ۆ./h�3�δ�#��[C�����ή&���y�O��\�K�M���4x��D�c.�b����/f�-��,Se�z���-h����ɨ�^����Z����]]��6�TFa5ּsqW�;[���ㇵZx��8��^�W]u�]Z����O����{G��[�������ۚ���G]=6s۠-��v��#��;e������}�vg��ʹ��B'���Y��S���t����7:��rl踧�MW_)�xa�ۆ������\���ܧ����W1��;�	�i�q�p���z�&�n��O�\m]F���q3탮5��z�p�[��Mu��ncq�M=�ٹw,��-���N�>M8�=�ca�lh�gd��9��̜yY㜊]+��. �����\�ƞk�vb8�������9�7 㧠생�;p�v�����n4�n�zK������C=��sa�q�֘p�N��>��q�vgn-�m��)�@��rf���IS>kc�-�w��{Cpd#e<v�Ж(8��]C�
����w[���nv3&�v�ǛQ��!{��Ѷ�D�l[>�m��;t�<��k���0`l�[Q���z��]W�ۋX�y*��wlK4��c�FOa�	=���lg<���vvar��ݔמ�v�����۳���{�q���9�W���0���u��ݸ̆1MX7S��	nӸ�A�]��+�X�kr۱��e�VwG`��f�'����s�[J�l���0�j��c�W��f՞�C��O�s��ͬ�m{O<q=�vp�'���2u��h���5�h�Π�m�6&��mR��\�Xݔ�cg���/].�۞t��q��۱�S�]M�sM���u��)݄׏,z�x��Wb½�xz������ڀ.���M���q���+�%��=�;[=�n�Ƅy�Xnx�J���Be��
V!=�T+Z�v��uD�A��c���j���k�C�q�mu�#���N+�s�{u��ףcD`�l�-������x�r' a�ҭ�:�s�p��M{V8�;k���b��&�����:�#nv��VŬk�8W6��9��wnPWs�\�����֖��F���kv�6�N|<�&�s.s�R%G!U��l�¬��rE�m�������n֮5{O���r⧭j����k�ٺ��+̭/ra�#;wf��a�۶��{i�D-�m�v���z��<�.�ϖ9^���P�˵ʩ�0t*�p�&[\�y��>�3�XzOF�u�������;�`���8�C{x��گf=���4�Ȗ�������'�m�+��m�vE�k��9�:�	��]�*엎��\�J�=���_a�q�]�����q�S��e{m���w{��e�Zq=k�B����vIm�����v7g\vōӯh�䮑pk��6q8�;��b�\�ny'n��"۳��M�6�z�Tt�%nx�Ggu�n7Y��̗l�㵍n�p��JD��w|ƻ��Z�ӭ�lu���v��=�\<s�u��i�qc]�{up��a�|���W���W:�^zѣ��z��A@$�[u�g�Φ1�g���Js���vU{^g�.Lk��zkv��x뱹{la�s��������7&�Pu�E�I���I�ݬg�S�������B盺��:��Ocu^��6�ce�e�\���O9[z����D�Y���`�\P�<�mW;����ڙn��e�5'7�V����m�M���ɤ��Gn^:�Q�.҅�[(/OHN7's'O�1���;U�;�ۅ�;{R(/gbv��v���O��F�1�F�:ջjF6^ݢ��.,��3�6��o=VÙ���:������\v�ckkCÜu���e�6"+<���6ֶan�m�v3rv���n���]m�֍u���xb��8���F�,ԵUJ�UUUUUUUUUUUUUU���cս����S! .\��vPQ�$�t�.ܮ��g/0�wr��r8�
���D@]�Y2��N<q����d.�'qu��v��
"zu�ZW9�Ur�&�W{A,��'��#��$T!3�;���*9vkx��Ruѡ�����\���<�U®R��RAUUs1���֑Ns13�r� I�#����"^�8�BA��.�HL�wH�P�Rol�*�W�!���ϦUE�w|D��Hx���u.=<*���s�Ҹ�-D��d�
��Hֹ�U�y�L���
�4
OQ�G�~����T�Qr	�\�\�P򲩕EP]�&�p�
�e�v������[�E�C��r�)���!*�(�2���)�zga�hky�]"����.�i��}��{�Ϳ���_��UJ�UUUUJ�UUUUJ�UA��g��ˏk��V��9�պ�X��/��q���)����ٶ�۱�k�1��/�)m�Id�9����ˏpU�O-U���]�tl6�:�-Ɗs�xn#@q�gqvv�[q���v��T��a�ݬ]�sjN_9�Q�wH�x}�1oU�q�Oۗ�v���ʕ�%�=��q�O3ҩN��-	�g+g�����룞�Z%�8�ݵt�b���N�p��]��pn�g[�ۇ��k�u��t�g{�Lq��Yw^3�o<�<�:�m�/C�ͷ��q.��k�ݍwI�m���*�{"�;k����N�Q7Vہ�x㮎ۮw:���lV�u��n��ٔ�Ot�ir��6�8½�&̦Kn=��;1[7���!���3�U�гv6��lv6f����[��=˖9���a�Cs�.}��f�m��;2�t<\��7���Q�	+sqQ�z.2��s�۷��Ģv<�����prUƜ������Վ�:��g�N�\�ݩ�t����gn�Y�9���L�\烝�g=ۓ)nh\����"�R������>��XW���NӁ܊�[[H��I~�"��JB��;���l�b|��Ŗ��0o�88�q���u� �� �2ĮgX�:D�ر��/s�Q��u�od{��v����=2
-�{f�\��ەʹ�V�����m�x7]��qۃ��']��ȥ�Um�MF
K��j�y�s�|m���7)��g�R��7�M���m�ۧf�9�1z:���p�ӏF�nv��#��`��]t#�p;��Y,b�Y�+úy�Z�bݍ�L�8N{\s��͵�N5i�@91��[��M�7��8��k1=��<a�m)%�ec<��Sue�R�4]=kQ��u�Bk�Z����{���ϊ����rxw�c&��g�{gm½���aNy0���^�{�t�\�繎^N�۶v�<�M��Ϸ'�/*��駔F����wY^��k���x����/GKے��u��K]��:��.G����㹩������b㈻����������c��+�D<���e�Q��'�"H�DH�E	������O�"US��ϗ��^{��`��ޕЀH�*���m�~fnw�W=�m��ܹ�3I�"u�\��X�����9�w�_�g٣�y�) ��9��I6|�śz�x��~=�f�q��X)+O~�v��9u���}˶��K�d�ρ�wܹ�H�z�h�P������]�˧W5F5@�$�ՋXؐ7�� �o���wxί/w��@A�w.`t�'��9UvEnL��Q��y�y�dZ��δuY�K�Y������@ ;�s4�⋚|Z�tM2s��%1�D�4Zs�;��qce��v;P��7N]q��K���x�J�	m��y{�Z��|�2���_�@;����)�[��:n�`�s;n�W�',D��+(fG5��G��U�s�\L(�1T�G6��V��[&YF��klk�s[[p%)(���x�^��^܋J���hK���;�?5�{���1�o{��I$���$���� ��y��7�6ڙ	q<83w_��[i��>w.� ��zŃm�<{O��|@ؐs��@ ���<B��PM��5%i�|��j׳ӗ�5�����7 D@�����D��U5�����a�Uu״ k��@v�E�b/������{��kS;����� �/wn�	 w��f��]=��=���m�ʙYISC���[}g�y��pO/���m+�/#e����M_~���uv�^���C��2p���!#���exwU����ʢIB5���Dno��P�p�IA	}c�g����� �'���` �t� �o��s|8{��H.�I��T��ώ���<�ˬH�S|�U�!�f��<�#~��S��of�Ffc�ͫ�^	�.����b�LO�E~>��n���9��ok�K����ߤݻ@|3��i�@ �}˟`}�t�ԑ��嶙���]��=�@�;��� ��=˘�9��~�I���[g��k��#r0m�Xԕ���o�� ��]}���r����:��s36$�ys ���Au���24؅�}��	kG��3=qkH봫����0��n����=~�����M�B؋��k����=ˬ  �7k�G���>��O�o�ɐ� ��)	���]�r�݅�0��_hoZ�쑵Øg���@|}�.��>��tI'I���<�_$�9���ȬՁa:��a"/Y� I���d�{�w�u�a$�/�������o�'�������X�
&L?{����t�H�� �?{=�-`����ހ������q����j]�����ܐ�
DyoM�i��Ț�o�Ȼk_�@��	;�2�a>������|��~w�Jm�ٓs�����n�`}���nA��嶒;� �L�s`�oͱ����IF�\�� �-oH��30�w�������]ߺx��T��cN�b���̽-j�ͻ<�)P]k�$�d�n.i�o�����n��I�k����� ��]ho��nq�&b�'�/P{[˦�M�۵�e��B�@RXW�zL��6!]��d����s�X �w�� o�����W���sW��Ov�$�5biJl$I� =�sY��e\�=�_^[����7�r�b=�s4�o6��*�:�[q�FϨ#�.��I$���d�$���fg� >�ܾ��r,Z�����o���{D�J�eeÞ��0 �}�N�}�7�a�� �$ Ͻ�BI����}}s�}�۹n�Ć86ga~Ny�\��Ap��r}0�-�=�����:̂sG�h��3���~|���f.ᘻ�7<9��$з9�8㨫n�<d��h�[�o7�/̙3���hV��]�l�q�6�Y�e�_:o�݈˽*�D��@&�*jkQ�ULW�Oc[5�=m�������sW�/����q�vS��+�-��� e�����s\��Y�l���n�]DJv�s�jV���j����u[LWY{pN�����=a ��Ɔzp���ju��HQ*vU��JE�Km;������sZy� #}�.dBf��1q�m�^��UV"" �j����85�cRV�b�o�X�h���s�� �U��I�I���a$���) ߷�g~��{� ;8�AÚ|AIa_��-���$�"�� ת�s����iva'	9���! '�}�~���l�A,! �-Ԧ�$N���A��;�曼�{Z��  9��� �g�g>:�����ER����K�r+5`XN�� =�_�NO�e�>�b�e�O�{� O{�S!�$�>I����������v�Z5I#����Pq��ok%�=�sɷ��kس�4�^�5��~����(�D_Ckr�$���"	's��\�b���Ut�����b ���ȏ^U�L����L���ց+Y��Y�y錟�z����#Oi��j@oe&C�h�mKm�����^fB�C�TG�3F��%�cFr~���u��$�$�{ܤ�I'	���ه�\\�q}���y'�}�kRV�`?{}���g-zA"F`]���sH�X�\�Y$�7:��Xh��і�_�b5�w.�������6���� gm�@ ~߹�uC����M� �}so�=m*n�S��M���6Na }��3!C.ON����<@|K�\ρ�3����~��X{�3:�yZEMůB	hDn���P}����
��m���㫖���]M`�������߇�*�:��������� 7����Cq{�0���5ѓ%��Cy8�p����t�Vr�e*r����y�����Y�{�;��;��q �A��@ {~�bX3�Yy_.c<kݝXYu�qO2ϋm3>�v�- 3~���A�<���X<ߧ�����[��ă8�'!�%ǐ�| �x�4.둰!IdÖ:�O"�b/N�,ˤF��;f���ַ���~泋r!k]#N}�kRV�7���z��b���'o��	&<7��Ȉ�A�|�Jo��ߕ��H��'Ś��-�5~�2.���&F�垬�]�\6MDw:�������9�S�	=r�Wu�~QĐy|v���ŝ��:]���]t�=֎����L��=�;M��vKry y��-��s���}ɬ��O;7�-V߮[� ����گԪZd�|3ۚσ;��[������_�6}��30��ݲp�K_x��q��HѰ|���+(f�w��m���\ ���5�1�v�@ {��� r{ۙ��H����V�)$d���%eW�_p� ޹�f �wsX�H ��iBA��^��~��w�n��"�v#ʹ��)Oq��.�qZ�y4�'{�;�w�Ϋפ�x,5YP�6k-���B�]��s>�B��j!�U\���=��3	$�ד�mҳ��ɳ=����^����;ɘ0�o~�@�޻�]ZǾ���ʙ+N����$TrV�/-�;�7��#�����N��el--T���MDyRW/ڟ�k������s.6 {���w��.fg�3�|=�L�`-�{��Sv���)�	�?̜&�~���	�OE�ֻ�  }���f �~�@���Fؘ�u�}�=����Y�@:��~������]- 8��rY��z�ǳ�@�vw���> 7�[��wY����;QC1�7�m�A��g���J�� �-���0{��w9�w�m����a���8����m���� �L�s��?N?T�9D��N}���o��@|��y��?s��h���i�k�|ѫǻ�!��ڞ����n=�~oi5n�˷�w]�Mc%��y.ƌ��|v�/��ċy��'�%��_�UUbk�ծ���V/;)�J�x��<�=��o>�Ső�n΋��8��ҊvN��ԣN��nr��1��:G�qt���q�C�3�+M�q��˶�I��j�I�������5���z���<dۻC��Y���;Q�s�8A�:��.�F9�s��7g���]���ŭ`�rp�ɫ����C��l��k�׶���;q�k�i�lf'�����(/Ј��(���T)ս�Q�?*����䃦wخ6|g9c�6/o�����w�����agd9���2	'c�M��XQtN6qRW/�0ֽ�� �W3�]W9]y\ HN��b;�o3 �O����nk[�X�=�c��hݒܐ�g���$���@8Os;��v��m�>� w��O7�UΕ��,ǈ0������<���������]PD��ޭ�@?��}�П/��6���w�Q�kT첺Z�QC[G��� �=̹����ɘ��f� �=��x�H��1,,�ۯ�������#	d�F�qg��K6�M�F���(�鸝�y�X�X{fjo����E'@�N�L�x�X��w�6�Ͼ퐞g;ۋo>ٯ��|��I��~��#Q���<����{�:MQq6�k��y�vz��̘�3w����]��V-�{��a�Ü��]�r޼���(�uM>�1��.���	Qh�	lK���0>7=�LX1j����x߬�(�(6yR�/�3�Z�30w�p@޺��_g2-�o�ܱ� �sy�`���rg�ou��nڅd�S>A�;x��.�R >u�b���}ə�Ӝ�כ\�w��v�c��H��/�j'K`����@~;˪N��^a 5}���'�i� ��,l��3����vY+qV�Q&��;L��7�k���dJ��*�P	U"�eT����et���|s��g�6|��2`�A�)��z��웗��t�9���^�İ�M(��P����b˥C	���?w{o�}[ OĞ��2�?jU$��~j��x�����Ȉ�[2e��U\����w'����s�=%`_4�0?��٬�^q��Y�7�kt���?���o[���J�b�..�xd��ץ0\0�5�~��7<�/jȓb[���K-�]ՙÅ�wښ7a�ƾkB'�W��t����-����X�p�h�5A�OEs���	��~��bge2�x	���5�X��`�:��6�<��G��t�	��Y�n�"I0Æ8��9�{]��vx��3���^8�z@L��#;���;��gzUDhY���#�;���|�^��:*&����CBf�J���B�g6f�^&��|9��1n���~钌=0��	6aw����|���qM�@����7<�`�z�eow�����mH���~�Ӛ������ogh�&4����(�P�͕sٌR�RFk�>ZB�ׁe9�bM�	��R���]��b.13�8Ccr�V�&�Q8-�"ӗ��r�9FK�E(����Y���;�5��O��Ԓ�q�p^��[��_��Fk���7�
�#�D�:��xےQa�����xiDW㲩�.��{{؏��V��oO]ૹK��� �����.���w��{(�-����&I�)��ui�D3چ����B�"���x��u(����K!�3����X�eB
U��AP�7�H̴ޚa�E��^�����qJz��F���tj���"�.��7tt�ݸ�5X�1QP�c�%�6�*K�����P��6�o�+�\��.�8�t��Qwܘ��dEQ��by$'�����"re����*��k��w$� �VD���H��
$�(�I�ȫ��Br�Ν��B"
ndzNC��κ:e��s�D��.�\��996�����'s�������U�M;.S(шWiĩ"��:	V�I�t��e�EP9�9]�iӮ{��PsT��AG92�E�*�f��2��KU�:亚$��cǺa}�:bJ��wbr+�K1+*Њ�@� 8��+S������w�x"�(��ݡ\�&hzz$�ND�&�ϝ�:�W�ӥ\��&�Z;� '1���un���m��{��������b����,oK
'��+e%�&$k^�y���2�m�&�ށLGKU6?&I����S�ћ����vs������*��j��͠ў���A��oX�����ſ/b͟ 5��� 
}�Y ��ə�Z�2y5�|��;9��S�d-��<���햎��Q[�'���e�r��;�'�E�&[1��û�W��{�= w~�f ~wkW�7�'���fѓ}�1`�>=;�4^���ZXZ��wy�` n.�ϼZ��|N�|��H�r�#�����<��o}u�0̚�G�A9m���ܺ��@���d$������.)i?�� G��Y�����0]�&��u~'�m���g{���8�-0���I��I7��7?{\�r/����>��ڠw}�z��ֽ�����6=�8�:;�����'=֧�����VFL�j2o��典���I�#':��	O�b?���~ɟ��3>����̙����_5���&���@���^2	'񜾥�7Y�.����ɻ������n;]�����1O7���d8Ӟ������M[��~eW�j%���A�9uC�>w�՜�A1�\�2#m�Cήy����~�b>�ݚý��0�Y�TJ�e�|o���$�j�-q������I�LﬀL�N����$��4��5q]o����7��3G]v�IeM������ot���s�"�(U'x|�چ"""|������rg�fC_Gڜ�N[f� �VMO����'�F���A0"#��S� �$_��_�;_�P6�s�/�۠{����H6��J����ٮ�m�%K��5���?	M�/\���!$D��3�o���q<��=-��֥{J����;,����/���{�nZ@$�����vx���-�c>�}G�r��_,����ٵ����/���m��akӇT���	��nx�z�^ȹ��d�tuN�R4�uq�̓����=�A�v�y:KÝu	u�=��=��`�g�gq����"�!L��e�[�u�uaJc�sq��������u�m���u]�K�=�ڮ�Es��{W]]��]�4!��֣��d�iw�m׳�)��1Q;�4]V�ۡ��p#���۩y��#.u�s]\8�c������W��	��G�,�_�?�k��� 9�e����<E����T��F$��ݬL�~�+�ÁjQ���s	�������Ә�z�Pt�4��7��h�sk���稲>}�/��c�/彫7B ���	�zb��>zr�@|
q�wrwU;�K�@ ����M��yM|��k��)d�VL�~�Y�����!�8J)Ɋ p�}���$���8���([���	���Kܙ��)���NV'-�1Oe���߹�<��~�@v{;3> zw�h >=�s1a�m{w��k4p�Ucŝ�9��6�y1X�v��9�����6Ƌ����e�zr'[����}7ܘ|ù4NI����'���|��F+�U�oӼ�@aD`>�m���k�I���ռ^�����1�WϺu/{�Z�H&��T���g��	���/��~������C;xE^�c��-���Aϖ�N��S�~���o~�I?�8�-��o�3>���7'z��ksݻ4��\����6�5�gn���y�vI%§���)���A$�UW� ����[��g�T(�[1�������]�u ����@ w�浀 >/��'j�{�#��?ğ�� ��n l�K*t3���X  �y�{�cS޳�9΀�۠ ;��3؍�����ڞ�{]�d����c�'m#�m��㥻]7Z���^x�A�uuN��]�]���M����(���+���|�˭�~�`g���m��n#,����@$����;NȠ��$�=`w�}�0	˾wTr�J�2I���$�M�}Ł?}�蟵�-��@��^R�%�6��2I'�~��a$�n9�<�TF^�9ƴ[�X�kGC#B�NӼSe���ϸi�>���~�C5m�mT��u�h�b���MJ{��T�K�;3��� ���X0ܿ�b�[5�UmjX Z�9��9/�"��;��G�$��wZx�/v�fb@�{��ѭ�IQ� ���ff`-�Y�k��e� �K�r<"#��ڻ��y���{ވ�{�I��N�}L�Ēo�'����y�z�5���9�QI"��D�t��b�P���x�� �2׵�>����˾��λ%$��C^Gw�$'	��l �ߪO�>����j�z��s��ŀ��Rv�j�-���d�z�G{~��O{uF�$���d�I$��H�N�rw��{���Tk�4���%i��o�X��nפ�A�Ӛ��;J��K�`{s>�����u�
�]R�%�l/�路����~�!'�(��� ��T�d�ﻧ�O�<y>^ËC��wI���O���)�o�����&��b�8v�Bΐ�o"ȳ��r��U��,�[���ü�Ł�]��U�-�����9���D�����w��R.|��Nv�v�'�N�T����BZ��w���7
펐%������cΓ����ن{fS{V5j�YS��nw�vy��S���ѝ5�I w�6I$����I���+��N{:�Ox�{�߷kz���x�$��T�a���&a>~+�Gy�>�ާ��@ �n�w��f���9:��k=Әˢz�*�٘�˭ �Ϻ�	����L'��^�3�����t@#���0Q��L���V�bA�M�e&�}�À}���� >�߷�� �_l�����Mm���t�A1u��m�_�a��30lA�Oo&w�5��=�b��}n�@���d��F���ǝL�ə��y��ﾤD�F3��@�Dl�9�m����=I�s�nz����8;�5�鍇�j�I�N�5��o����mDq�dM��>E'��m0�h�;-�:�Vo]��o.Wv�׏��;Y����\�݋z��D@��q�7='<s�5g�sUn��nT��1gR���:�vܽLݹ�C"�Wu�R�7a�M���e�97f�-�^��<2�@3����6��m�w���El9wnz�ƗhBh���9G$�BhEèݚ�i��{--a1yx�(Y4Վ���M|=֎��Ӫ��s��zV�jm�fi�k����o��`| ���ςvx=�מ�rk���Y� ;��o[��ڬ�0%��2oа7�eǗ��~c��DO�Na=�V���}�ǿy��[Q浺s�^٧,��,���߷�m�wӻ5	$�0�w���D�O�;�HA�H���f}�d��S�	�l�|���fgNu��͠[�֞b�ovf�=���?�{>oQ~��'�I���~ӌ�ʒV�g��M�>� �9t�}�����{ݠ;sy�@|w��3|�7=�4��/W�l׎�v�%i�bh�Mr�t[����e����u�B�����՘������_�_������׳�� ���b��U6E�D�q8�-���c���Ł��{��&�~u�f�gn���o��L��܈�q˭��z�t�	���[�� ��9������l��+:Sɶ�z�Ed��r��[&�l�:>h]b�}�s�I#p�{�ZoD����u��{��M���>�����Y*`K1�a�̸�m�ܵ���g��a,�w��t��� ����TM��a)%,��0���絼��r�> <k��q�߹n�@��sZ��-��������LXf]5���N[f`?z&�$�3��?C(W/���(zBN=��� ��Xސ��fa�?]��\��_*g�շ����ڬaS� �^����Z^��/�5�-t�
o6�v	�uY%i��ӻ�\�Ü�� �9��o��.����FN{�>�� ���Xް�l^mvR�/����@�~��]Uf���?�(D@���I�D������H�GZԥ,����&�Zu�f�ۥA ���5�`| {��Cx��l����02/��X����=�D�;�t���$gxm�Ñ�0��{�ncXyz�=%�,��շ�U��x�{��F�ζ��rw�6�������"�VZ��<3�>��o��Gl��7u�� ��70�H��v�M]��7 ����I�ָ��W
YeTa��y� ��tQRߴT����d����&I�Gw��A�I7~��C�OI��xφ�qnCk�1bnK$���L���7^Wiط�ʹr�񙩷�#눵��l��נo7�kOD{e�$ۇ��`�Ϊ�	�z�Y�Z��b�VIZy�Oo��uf���T���s M��'�@��ka2Z���h?r@1��G�e�QI~h%���@?���tP <��U٫��i��}�ϰ`��1,�kݶ؄JӮS5�go�J��_9�k9�<@���rf��d�Ӯ[�絡����^z	��syh�1c3�[N��ʙw/aw�¾p���?ՠJ�m�t�b�:�T'���	#�����	�m��cLm���w~$}��9z^��b�VJ��O>3�e��|?rꓞ��{����0 |=�LX3�>6yT���npe�u����'ꨚ&���g�3۶��=��kW&iN���j#�l�笚�G����z����A��9�o1`�=�b��D@��U7��Lm:���O�4����0bÞ�Ł��F��Z��c|��U"9A�ܵE,ԯ=� ���d�I�I�w�Z�%���}:W[�W�b�VIZy��o�M�>��%NSs[Wb�o�ڨ |}�{�d 0��,�c�g�b�-�j�5�w�R��K߀�<f�����,m���z�t֪��o��z@#S]��ϼkݲآ5j1�&��$����z_��w�{���~9�4�@߹�u%�a�O����P	��o� ����������u�Bǉ5�6�i��a��"ͧ�
�'��;NJ�,�ٺO�6�U#۬�xv������}�2I�p7��+�ձL����^��6o�¹���(9q窍�l�}�Á{n�iU�� ;4����[��͝x�FF-[���%e�\R���Se�*af,s (��C�"����^��y:O�;��������Du�!�s���rI�\�1�����ԭ��m���mK�!�{�'7�D�5�y*L�m��h�mvo���A٬�Ql�S���v�[1ay �E5���[��Ұ��m��C�HNVV��i|��G*2i;�lLn�M���u�ٚtSe��&f](�'LA�Y�lT�3r�B�4^�1��A'�s�pC��|籿on�@6j�F���{_�:����!��V��4ؚr��VJ�� I�u=���I��}d�=�� +8wb8�Td�#;��ٷw�>�7{��fԷr+�U��s�ӹy��q���GD�8|�nt�=&|�<=BY\�I�]Z[���K�<��<��l:�sٯw���᥁y�+[y,�3R�5P�b�TA^{��O�����v�l��Vǃp�v�<�7}��;�=�8���Og_�^i^>;3�P��2lF� ��u#$N����MY�r&�]��^�Nnl".�z�{��[dqo�:z�V��q�A��������}:$U~�����D�Q$Zv�:�tR��aG��Tm�/$s�n8���'H�'79�����E�:u-�5P5���g"��s�p�f$hҕ�#���Q�_:<�:ug)��11eI�TJ�Bwn��^t�O�t�!:VE�R��^E��盂�v��!|�w��%��I��}D�NT_�;����
**�!}��8�eQO0��s1�\�#���U���HDAf�%��t�QRQ��A+hE��:�A��z[��b]ΖHE楅�	%(��NE�
�)8���LeQ�y����&F�i�J�<���Q$�s�B�w#�&��J�I$���L�Q�ߗ�/��e��m�UUUUUUUUUUUUUUu��������]U�ս�ڻ�ו���Y���6ϱtB����7V�v��b�^�[Zx*������v��@<��xcۃ -��e�γ�G846��)w^�0mn1�7x�<m�ŋI�P�J�T�THV���&�NS��n��ε�ޝ�\c�v(G���gn�^���ݩ:�u��ř^��hq�u3�sx�#6�'U�r�/Wcq��͞-�Z&���{iݫ<�6����A&��9�E���p�A�D��y�̐�g��p8����b��Ѹwl�\"��bN��h��k�:�]��Gb�+t�Y8z�	��y�;����;]Om����vl�y)�ۮ�:y�.z�a�va���F�4=�.����wKۭ7'nz�L=�6��c�3dB�g�a��+��f8:�g5nM��<7l�4�5q;nۧ&�����x�*a�]�1nn�[XG�rvh�==Gg��W�u�u�.���u��Z.^���#�M�1͞q����n��������|v�F�h�.�Am[��q6�6��*u�\���Ϟy�zv{k%3��-�D�"�K��V�i����/�=�&r�J�.{k�];�c��8y��|V�+��[.n^�7)� hvz��a�I�=���\cm����aᮺ��Z�܆-���7GY����Lϗ��V�ͳ�A����RɜO��1��-���lxsЛX�]��;]& })s�����s�ն���V�	u��ƀ�5���hc�ָι��x��DDv�6q*t�݌�Q�ǵ�v���/7]uj�n�cY�;z��=v���
�N;6�Wg�=�ڭ���"L��q���y)�=�y7Wc�5�k�p�,�X8K��c7GnC5�o=i�'�=�0{rk	d�X�z�b#^1V��K��Z�Mu�C]/���sUUU]�{�o�UU�ܵCT=H����e�;y0��kݙ�w�Hת��÷bx�U����۱��t�:'��O=����{d{[r	�+��|�v���v��N����^�E�˪سۃ�Z�װq�k�Ά6lk�<�i^aAv6^!<p�qn�����>=�RZ-۝���2���s�@O(�I/9kl�(ܵ�L���?8�k�'*�z-��<Nr�6[�v���{��=�\�t�5�Z�������b�7f���g��@�{�J��	�{���a-��c�O�>��k 	���k�N7�s,����X�b=��3����E�W����g�p@ rw�7�����(�x5ֻ��Kmr��(dEe���2KX����e��l߹���z4���f^��N8�b�DG�D{�,窅� �tjf��0��-�ܧյz߯~ �� ��33���3Y�[�ᑶ�5f�³�Q�r�YZ���u� >�2�W�jcy���r� �{��x��ɟa����5��I���9	]����$��@�۫�=t/nކ�Ct��y��T�������4�َ:g���c����>�s�	$
}�k�M���%�c�x��ݍ������o7��uR\�Z��a�ȡ'���%��4�?B6n��z"�I����w�|2L��<���ں�N�U����]���W�n�É��#v0S
D�� ���.ԟ� �}� 7��fB	+����.r�����r�[m����������&���cl���7�~߹�����s\ѡN��X����e{������ =�k0>��ww�$S�-����c�s��I��HKX���+�J����qk >Ü��7�ﻯ	�w��O�@����I��- ���٫;��}g�F��#d��\�<��#r��Q���D�V��)Gk�vΑG��%kw��{1`����k�@�{�h9m;����#��f,�۸�6g�e�DJ�VY���;uC�������ٷ���o��ws @#sܱ�o��AC~������D#���b��bZ��>�ң`bJ���*ў���Wm���Y���.m#�({�a�C��<g�5������4�N˽��[{	`�8��6���]�~�B���d`F�ʤ���o*jI)$�	0�=gѤ�����$��� z{�7�;�s�/S��~�Mi0SN� '$5�9�T �;��d?4��/�Χ�"��9��I=��4� �}��{3;w5#�p=<l�	v���@��`��{su��z��a��6۵y2��P��˙ ��534A��<�$�����`Ds��	t1�]�I̭�$��*��8�qr�IZ��k�߷����|�˹���^�[�-a� ���@#��z�.��3������9U���Z��DU�e��wS�@� �9�f���or��YyM��J�����ܤ����ġ����ou������̣�7�w��@ �n�}!�<q��lPo�����_7�m4{��0�K��\����eƺ9u�B*�!������w�§:2�B{��5�d���;�%���z� �ۿ�ޮ�;�������vR�H����>�N��)����r������������a�ﳞ��61�M�B�5]���X�I�[�x���/>+[�2S��i	-L�����e��G�;��6�  �o۹�圽���t�.��nS@��3��7���k$i��������=۬qdSӼ�כ|��`���z�)$��U2p��路�����wL@.�8ț���J�\5�o�
I�G��� ?��s��3͌�패���H�;�����w06g�e+����c���~��M$��K��I����Np����-�R}��r�Lw�����'A���K1�@��� q���pk�vY�_4���[@����)��H��Z���'��w<ha�[>���j��ҩ��9�b��:��*Դ�i�P�S�*�j���q6��ǛG;7U^�m��խ������w�����{���4CsX+�����b��)��<�7\����&�\�ǎ���f]��t�4qm׉zz�썙z�e�u��a�u\�v�����[�;i�g���0�-΍ukc��Kۈ�v�v3��d	���:����u���`�۱"��v�9�,�v�c�	ֻ��7f1u��5[rX�;P�F�[Vf���F�7�B��5ѭԛ!��	����L�;Y��Yw���ҁ-��޿^��I _�0!"��h����vW��G����퍱w�\X4jE�;(`I# ��\�%�}�}
���ߩ �O��.` ��@ ��&��͋�e3ٛ�[mh�0��V�6��w�X|��9t�� .�u�?^��z{�� �ys o~�t�!�8�%kU�����Z綉| ?w{ϖ�� �w��@ ����&߷��x? wɉL�-G����Kc '�q����w��g�)�{����˘�� ���@�y��9w�5�}���' ��$��[`Ź��ؽ�Oj���T�!�h9(�qWL���{�N�T�l������`�@�=˭ �����g���F�o���	���x���[����r�Y-�����wY��������O���ָ=*�	#����Qb��S0�mN�\����W4qMS|���a��}������55]}?/��}�Z�����}�t�ǻ�z�A&p=޴M�ϼ�+r���m5�=�Z ;�w6�6 ̓�H��x�9�韛��w�U�[�{��-Zѐv�IZx���������m���h�{|�w�����t��i�x� �ۤ\�(�P����-���" ���̺/Z�B�� o�$ �{޷� �I��S!/��Q@��4ֽ���R�XH�n�ڢvс��Ƭ]sOnUzl>7tV�S�«lW�����ϯų5�9��9��'�� �O_��T;��g:�)mR���n�+^���`U
�:�	��}f�&;�4����q��D�� ���lM�sM��Ջ��o��-�-����:��� ?O��I���&B���$wH���gpD���+�Z}7Uh<9�#R/z��A?o�z���l+��8�k���X�3X������I�_��o���o��,�h>��ߋm3�e5]=E�k4�"""j�捂IQ�f����,߷{�,���[��/Pﳻ��V�dO*9+O3���� ��<GH���8�;>����<o�d @#sܳH70O�K�^\v�uU%n�A�"�[�Љ�φ�s�ݑ=G8�r�v�-�n���"L��13D]}�^��z ��o @#sܱ�;U�^����{�ox����w1`-��t�����5��u&�F�4���C������&=�~��| ��,�0}EUo7{��y�{���j�-�}_��\>� |=˥C�n��]}�� |vo���>�ܳ@kK���	i$�o1��o����w`7�=��� �G��f�$�=�����g�|����M��v�d�&1���e�le��uo�{jLԭ�s�ܾǗ}�$(������y�
Wns�w��4��o���U���O���g�\�
���~-�����_P�ƿn�z��N�AK�� d�S�D��<�lDG�#��绰��F�#n���6�;q�d5�፴�n:�me$��ώB�z�u;Weyݴv'U���|3�����x�$�s�w޴W<�j}�w%�w�� ���yf�`���G�$�����>�ܤ�%�w�{�������I$���h;�w����\�X����^�̝�t�C�v�>�v��������s���k��wޜ3ݚ�@���Y��@��w�����О@ݪ��i�;����_j��@�r��  ߹��7�H�~��^�Q��N��h��5yk$��̮�[a%x�/��[ t߷��G�w�]
����|@|s|�w��3�#���b��WU�ߖq����j��{�k�����r\��A���}�7S5�J�}���3q��:�g�ťo�o�CK��I%��9�n�m��'�m��J>�6y/q���t��ht�s�2�wg��sڍ�V;nܤ�f:M`�li]�!Ηg�"��sj\v�x��p�
m�u^�<�At/��r�N���ތ��k�����b�$�n��V��ٍZ��E�cm�^��0X�q��k����\�t�5�<iY9@�n4j��v�\��ܽ`5��X#3dv{^���5�7I��k�x�B퓋C��˻tsٶ�\XΫm������Lo�uP��{��`��Q��x"5r�,p"f�U�_,�߷��7�Z�� ����<o��b��WN7h�fT��'���N�"!M�s>���u;�߹����y���n>�$�ew��g~�}7��� �k�����z�8����@ >F���{[ɿng�m��u�S>�v��|�Fv��g��믉��fs|��>�oۚ� F�*������5]�p��b ��ZJ[ �J�$�#�ܚ>�߽�y�j��<�z�I$�m��$��r�I�v˺ٞ�%�P-i�$v;,N8�ĉ[��+�nD[��ݨ�P9T"�����˜��r��m��.���`������ n{�i ���2&i��gw��`�߷3�Z�����H8{.� �L�I���{�ޘ�45�q�?y���7J���'ȶ����
���_L��ߋ�)Z�U��6�#�Ta�2%��ǂ4Tn�XG�� Ky������RE$�_�ֵ$R;��qڣp���	31���b�H�\n�+OX��{�p@��]}A ��*������D�>�L���(�Eĩ��b���n�̙k(�f����MԪ|*Ua�E���f{��m�{��ǧsOɛ5��������s�,�V��iF�D�w�2���iF�J��{��;ij�w���_�o�m)�4��)�ǹܣi���=1XX#�&t��Q�f�̙g^ZT�TJ��Q*g���6�1m�y�Lk�����-�Q����r�5�ph���ST���<ɖ�����iF�
�w��s���m�h������~����/��n�����y�Kv�6�z�ۨIbeVIl�����������ҍFj�w��<�m*EEM***h��9�:"�J�2�T�ҦW{��[im�tҦf��^�/&8�gK�Fz��ekw���*j�0�{<ɖ��M�2����ħ0��)�"5l��g���;kl6�5L)�a�{��OW��ߟ�j���}�me�aHj���e5M��2e�iF��5M*�w��3���Q�ҏz.�q�92v�N�}�ʿ������g�9U��q�i[Q�s��L���MQQ*j�D���w�����*j�M�2d1��}�=
��_g �ͩ��ۨ��z"}�&-�N0�ݱ�e{|&<�Iz�������p#�A���؊�g�z�o�Y`���-���O�4��|Yc�|����Ҁ�ܿ^C��k��Q=�};�W������n�3I��9$_���Y=a�=H�"A���ˇ��o�M���&1�n<��d7̆�5^qz�XC�k=�x��ڽM��{;w5��������{� A���_ꎘ��O\E��B�|2�#UF`U��m��Gi]�F#XQ�3s�N�W{"�n�uk�Y�������[��x��3�e�ˑg,����lUo��k��>	y�����L	�n�P1�F�<=�g��N]�ɓν���$���΍��;���L[��<sm\���gb@m�Ǿ�<S�>^wYK�`����k��>ҷ,��*���4l�#�z�J�֮��|�L�����^����A S���K��$US�K�2q���BW�5{n
t��)ҟCo�ݽ��׬^��(�MS�
~�j��dbǳ�|̻ɣH���|+{�W�յ�볻���q#xi/���o����.a �Pde�ϲ[f[ͳ��}��yk{���Z����YI�1�����"��7^đ���|��'��ے�}��/W({J�y��zzU�&Ad�3eVA���d쵗���:7H���f�U@�n�����ؗj�5m���["k5���3�iFQ�o��Ϛڶ�ٖ�ۦ65��w��L�*�w�9;8	��Nd����T���y��vC�3E�e��W��
5�\��i�Qj����'�	�bh�I9�����x�9
�(�NNE�$4�"�U�&B<˹��^�����B��QI����t�Ca����tԬ����TkN^�����P�
.�jDT�5�R�n�<�,1]�pTO	��m��zY����II�Rҭm20�Vki�̺�1���r�	��v�uL<���s�
��!YQ�#4u�P��+Nv��=��
����h��9r��r���K���ºE����uݑ�J��H�/"���u��S�r������_$�}P��[����UHWdfI2�BtԹp�֐�_g��]�[N���j.�b���8�|�?�߯!���!�����5MRe{��L�M(�a��j�Q���3m����g,�Tu:<Xf�ձ[�����r�^�M�/9ϳ7me�]nv�8�������[�nt�<����������Q��(���}yE4��s��;��Ķ�v���t½��&Z�hh���t���T�~*Ua�E��Zh�k��3���m�j��0���gw��Kk[�_(��Z�R�k-i�l�������Tš�T�N���T=�o��Kf⦔j4���g7�^QN�[J���rs������e��ʛ����V��mQڴH[;v��nCB�s=����B�o3�|�>�v����Z��e�T�����3����i[Q�1ST�)�e7�^�M[,h���Q���w��amq��V/:ɖ������5MS
MS/�߳���mSE.g���)a@�b��|?���{�\N��Ң����Ou�v�+���'��dͨ�ҧC)�MF�e����Jٴ�L�M*j�C�ϯ(���T�t�MS�q��ڐ�nşI|$�H����5$TRޑ�X�L�w~���a����)�j���ג��V����MSE̗ǎo�i�rs�κe�iF��j�UP�����V�iM�M*t�g7�^QN�[J�Y�Iu��a:�1�i[Q�{��L��w|�i[T���T��^�m�b�T銚�Rh����=yE5�X�MSJ5�D���Y������U_�Ĩ��qP#x��Kst��!��p��G`/��}�zsp�͞�9�u�b��|U����gX�Mfcw�t��*d�۫�<y$$��kM(�a�S/�߳���mSE�a,��0T�4F���MS>/�X<5m*U4�**h��9�:"�J�/����M�'�E�D�zH�k��}�BO�2�4��Uo>����J5�ST��[�g�F�'�A�I�ۦ#�>�-�FPC�A%+$��(!T/2si��^{���5�Q��m��(�T�T��<���xh�k��3���mST0���ST������5MSE2�����2�4�Q�\�u��X�+;�\iF{9�3m.���R���5�㷔SZiF_*���V1,�V��,t�Wx�L�O*j4�Z�o|�L{��\f��o6�Ŷ����e�2�7�^�M[-����j4Owɖ���45MS	W�K�Fsu3��{�gmL�T�Qw]^y-b�f-�����k=w�#o[J�*iF�D��̙j�Q�ҏL��3��91�&g�{i[8�4��ҍQP����)�W��J5'��d�TҍFhΎvY�f	��H�[J3ؽw6�9sت�v^0(�z�����Iu�X���5MSJ5(��<і��N��*N���g�~�m��v�F̪iF�J>��kY��v�iS*��!�:u�	��5M+e��+����4�Ҧ�J5J�T�������o�����X�e����Q�\�{zE5l��MST����9�MSST����߻�i[Q����}��=i�[�����7�Ӳ8�苋�L�����l�&<ܗ{/Y�Qvى�♓(�`�Tom�;���ޗ���;����}���Z�3-��mR!�����a��s˕/c���lq���v���D�\v:���;zݫv�r�t׵e������z�ַn#���j����Ϝ��GF"��;yᲿ��|�w���q.��.�IP���=��Է���v����@p���,�z��g�ܻ7lu�F.x��]��u��]�ŗ�=�\�\��K;�lFf��h�..�u�xCf9;ru��mIn9yK����V7j�e���a�c���|����0T�>֘�N��v���,xj�TTTҢ����-SJ=2�T�ҦP{���m-�i�J���V99�u���P�3�eի�SQ�1ST�K���Ѭ(��E����#!��L3H���h�k��3��0�T�0������g��V���K�VҍF�L������d�TҍF�j4�T=��s���Sa4��{�_l��޷�S�-���c�Kls�i�}�m8�[��X�4�Z
�SUQ*g�|�m�mS����� �I��{y�m���^J�	>�𦩪aMST���4�0����ST�{���m+j4o�癪�+1$UN>�=�2}$oRV�y<�7T�q��QSJ�*h��x3��Ҧ�J5Q����u��ٷM*e�T�g7�^QM{�z�`�r��c>~KmG����@�����T�4ST���f���`s�#Ze�S9�߳����aMS
����=y-�5d	���_�iq�Y�>D�I�t�a�1i�T�N���C��w;ioqSJ5Q��g7�^QN�[J��k������M��}
���{^8�%F�:���z�x����%�ugY�ĕ;U�����R��%����?���S-SJ5�STTJ�}�w6�1m�iF�)4ST�o����J5���vot��j���k���������)�g�|�vѶm�h�gYd��u��T�4F���5L����[�VҍF��#3�Lל�ؘ�+��ǹ��q9��]1Tq�L����o����6{!4��sa:�U����]���L,[��	���k~�ҧI�ҧI�ҦQ���ƶ��6�4���MUC���"��J5Q��g.V�y�sa�kx:�4�Q���.��M�R��4�Ѣ��������mST)�aMST�ﷂڶ��&��h�
`o�ί�z�����4q�l�s~�pC�a����=?�������P�1%��5�g�U�4��\s~��lIgXײy�cB=��24��1���9�͝�o��n��*j4��fo�����αT�8�q�Eb�$��h�!�k�x��A$��0gPD~ϋ���؆��7�l��j��XF��J1�L=�s�44F��~���;�۪��J��=m=7���4+��Y�0�{fn��ę/S���nz<,�L�F�&���7܅��(0�(5;~�i����#_;|>�����VG��n����da�=4�Y�q��
���c�l^��1�4�^���]M��Zgy�{%�+ah�Dh��XFZ4�#F(�o������CiT�u;���=�#�m���&`��#L3Dh48��{�'�!�@/~t,�G�9�� ���D��+�.��/���JI�/y^��K����µ��ќ�qv���>���g�;"t��2n\v�k4L�a^���q,=k�k� �����Cf���^�QMi�F(�>7��bE�d�IS��&h����τ��+�� ���I�d,��(����rh��20;�sX��i�"�܁�^�u��J�&�O���_��zh#95s��x��f�����40#ڀҌ�9��+`��׹��>w���������)�M��a���y�M-F�j4��g{��"�������&��k��݂����8*42��m1B{oc#pC'3v:跮��Gk-U[U�~���ֹ-Al���ɴkuw���$�{�����A;�o�؆��3�ހ���{�E1��`o���i4F����xXU��"4i4F{��,alPaX���51ù�ya��Y�M���������2i��h"q�l�}���!�"7��t��c<�j����6uk9n;��`��c�l]��3L�Q�l����`�l �"h����1�{��S�rk[E4ph�Pa�g7�`�KMF�MF�j3��{�X�i!jֲ8?�B��%���ܟ��r��Wr켱$$��Π���G�{��@�,`FA��7x�߄�h��27�JK����rg#S�.����F���z ������:�����:(��g���y�E�4jbl�4�d�u�x���HH>���F�{��ѥ�����b��Ua�E�[Df�>/�LCiX�h��/&��ҕ�;}�Z�S�X20&�zɦ�C�q�����˂�#�������Hk����v�`�/M�ޟ��� �vמ*�U�u���z�c��p�7R����}~����a���u���4��D4�Q��s��i��A�4F�����4hh�^�7�wy�+�3y��i���J&�JF{��r+e� o>�w��&14[An4\������6#7ӵ��T���=�:�#�ph#!�����L���D3u~��Ca�=�J�/��t���a�]�QpiaV�YDh�Dg��o!l-�#�9/הa�����Wp�3����L��ӌDR�܁e�Dq���yF�ɬ��;E`��c�i�����_uÖ�nXbPiFo~�r[��Q��v�פa�lA#�F�Ά{�c��j�����G���>Q��潼��m�4To���&�4h��y�a�ҐD�����("?c�̭{g�� �-dG9z���X��Cj3�}��i�F(�0�{�4|0�A�W��{�슿�@�v�����݊���K�^�`��$[�PN�bZ�Ҿ��۹'�c��=���!�=��֪��B�.*�Akb��o�xx 꿚����c�w-۲���P<vِ��xnn�)-�tn�H���sհ�u��<�����E�e�c�+����r�.;u�O/=�`�#����sƺۖ��d��ϔ�x=ۢ�=nv�6Nnu�҄�d���38"�.
��W*;��W�;��פ�D��=rg�<��v}k^��8�>Wum�Nҭ��������c%CO�[��t܃Y7	����{�� VZԒ:��%t��F�t~,�&��1��u̇�alQ�bGe��i����`FF/��M1��S/�m�ffoyb1!����\�#�=W��0��FK�F��w�LV��4ŝ{�4��Q���9�yᴩ��5̞LV�1F��&��zF4���;�s�Z�Ci_{׺�m�{�[��5��@� ��b�EI��3GE��E���1Rlw���!�b�w^�&}݁�q������0֚Q�b�"a���4Ѥ�&tq�M��Xoi�M�ƻ���kS{~�g��[�X�G��̚�JQ�#w��M4q�lCg��� <W/�p��؇�"8�5��Q�!�F��������he�{�x4�6�4�Q�}�y�4�ؿls��͊4a�4vg��0�6-�s��1�������Ȭlc���{Y|����?o�j�p���/f��c5Qe(��&��<��%9h�\���~B�9Z���_��ٮ{!��"�! �stA�n4���y�-���{���2Z���織a�4����|�0i�I�4^s!�Tx�%V�i�l�}��3�@��U<+��w�o�53T`Q�Y����X�;��b��\���b+��I�ں���*����D��Z,�}�$����UJ�_+� ��1=��ҍFd`M�{�4�iƂ!�!����2�� ����ڮ�8��yFZ��a�իE��%����?z�kH�F�b=�w�,��b�4F����N�u��h������4��5Q�ҍFw��2+L�[ϸG]�RҪJb��-���{|�]���;�ze��)�܂"�g���!�4�l�߻�l�dLѹ~��z<��=�V6��Saf�X4Ѧ��3���om��x+H�#9��yalPF������Yi{���ü��T���V���b؆���@�!��#F�yF��U{o�o��&0���U�;C�vٝ��g�\r�9����f�<�'M��q��U*�2[�%����*�_�Hj(�iF_}�d��lCh��n���0ѡ�1sW��7X�|��3�,Cihj1��{̊�[���������m��2O,D�E�5�&>��M�`��G�#���H��<l�dj3u�^Q��4��jcs��V��З�`�G�����8��<�%V�i�lϽ��:�ؠ0�(5;5�ɤ�X����
��M��٤�W�����	.۫x^��wx ���vNa�
�$L�,Q���=��"|W���	~z����2��J���s���!�{Z��!�C}���4�;�#F�/(��A֣l9?}bh��Ii�k��ޫr���٭�؆�F�g�����l � �&�\�#h�Q�b�=�s�[�s1-�X!��i�@�iA��k\����I��P��Qik%1m���c�a��!��"H!�=�stA�o^sE�:h#'��w@[-�j3��^Q��4��A�w�`�F�Dh�k����jejV�O�V�+jD�rAyrƱ�-�n���079�pб���w�� ��?�vb/8��1y�bG&�y4�ZQ������s&�4��M�#����qHf����!�"8�r���0�6�f��'�����n$������ucX�`F!������c��Zd�u���LQ�4F��v�4i4F(�0;�sZZj4�5Z�{}��r�\Xf7����-�XX�Ghp�Xf��6����<���{�0gDh#�d�����j:�x�dL��ׯ(��hb�#����!�h��8�&J�U�i�m�ﯹ
�{u|7�Y|�q�iF�G��ܚk-(�`FF/|�M4h#�D$;�w�3K��-->�[�����[������]G?G������e��v�!�f,<�G(cЕp�F��9LY��[��!$O���#��+]�Q��������+�KMbk��ޫ��F�ҌCg�9�d�+a�<�����p]h��'�Z����4F(0�Q�߹�M-&�JF�j3��y�[-��3g�؛c�1I�o����=�5��4�B��Y���h�K*��X���!�����IO�m!�bg����$	 ������6C��y�-���8���[-lg��Q��4�1F0�y�bF2m�-��0VQ6��k��X0�(�4��.e��z�9=��0��Q�߹�,Ch4����� ]��o��j�����ɠ����nV	�	�c�l\��������J2���%�[� 4F�[f��_J�{�G�#�G���t1�m-F���=�dV�`L�c]x(�c�3DbG'�̇kv�+9�#�A����2�7��8d�=�he�##5n���0�6ku�nr���A�����F�#D=��	���Ua�E���܇Sb�#�;9�ɦ�ҝ�-���r��-���~���A�Ƃ8�I��@�pC�7-�
8��8rݥ���6֫;����%�0�&�9ż��7$s�j��H���wֽ&S�6���~(/u~X`39f!��Ý�0�k��B���#j���zOr��k\���z{���A%uEy34,�p�:c8�kg�����O����{��X�������q��ޙ�,_���$�+�f��wrn�&�O��;e��-:��:onr=�NgNԛy������p��kG�I�5���B�Cżh�u�w����=��2���z�ʽ:�}]�XQ~��G����g�/�յ��b�r�I�@���TSf2K��. b����S�<��xx���zs��F������a.]T5؇~]��n�͞�������k���ѩ�)�2�3�,�T����[��У}�0mS���໒h[�f�	Ԃ6�:6쬒%�X%��X�,�;0���kH�jЭ���M
����C�RL�\�=S�徽��李�U�G��8G��>ӻ���:'NLi��[���Z9u-ncbfc��öE=�dc��d�;&̈s+��͇'��(~�-_op,`%c�{�H���[)봴Н�-jUK��ð��Wa��q�l�Wl�Nb�?9���t/ݵsG�H1s^�g��a��f/{�;Xn<�ڮ�pw�}��gO(HЕ.�B×�;�6#�o��8�����GPW��|�� ;6M�[&��" td$���1���_����>��ӟ�h]"����]��p�բ�_N֤�X����dH��:�t��"�C��r&���Xi��ܒJ�AE��NU_*���r�D*"M"��e])�;�L����JǄ�������"�D�e��L����9\�UG�h�d䁣L�ӳwtL�e!	$!�vA')J���'U��.UЎY�I��I���F*ZaIQ�d!FE�XZ�U�Q��,$Ò)�˂��e��*��-0�P���,&�[�W�J)o�E�D�r&��*D0Zp1Vjd����$fU��&!\���j���C�wCD���*Y�FM2�Q]�ZDr�dfBE�e�fbibZXY�u��S�I�x��ft��*�G�;��~������������������:�Q=��9�i�N���\M�9:��uF4�*�;i"��p�u�/kg]�k���a.�k����2S��8�յNݶ莳d�ѭ�������}�y������"��S�y�8�qˎ_j:w��`n��YY�+u��e1����d�'ml�}PzO'U.v\��8���՜�S�ۑۛ<؃Q�WOg��my��g�d����[9-�����O99;�G��óJ)`��n7�|�f��{lz��FI��dTN��������C���d!Y
�%�I�15L"��ˣ���k��:���;vz��ۚA�ۢ���|fƽ��1��)��m�0=pr�cr`��75��;���v�u�ݔPoe</c��b#�k�[�}���箃�]�^����ܱM�=��[�!)�<�Lx�Þ�5v��
]n�����ьvk��������n�;�prN�nnM�q��9ڛ]����暘;�+=��"Y$�xY��볍�X��^g8��g�[e������Ady���u����5ݸ���S:�\�ʶ�^���׷�����a��F���k ���k����@Ld�b�'��<i�ɻg��Z���[q'�����]��ϋtT��a�mnäG���t��/n��\���'�K�C�� ���\�s'cn:�l<;���9��s�/:Γ��0�hӮЅ��z���ټpe;y��E�h݃ɐ�D�-C�g��ی[3k'O�����s/�:��X�)u��n;:�L��&���ѳE1�{u�\I��tt��׶�7n����?�uϷ7��8�>�Y���Ό�l���f{���=`�g\��6܇H]�sr�`�Sg��kx8��;q-�<����v	�6��2���k�m��r�v9���c�Vuu2�l�KW8�5�UUU���w��t�>UUW#�y�z��N뗭�O�.���������ȚΈ0ˮو�ba5�2�]����.�n}r�#��v�rs�9.��s���8��v3юЎG���<ױ���c;
��-�S]sι6p���<��qx�vS2�E�x-�9��\c�%p�:�-��mQ�n��ݡ3�sz�77��luK�;J�ɛ	��:��p5�.^�a��]��n��8�܇�ѓ���;M�Y���lgQ����}C��`�40#ڍ(�s��@��,h��{w�a�CDb��{��N��Wk1tf���!��5Q?��w���km$s_��'��Id)�lCh��o!�划�}���N���`�`���F!��{��c1�����(�ZiF�0޷�W��`�^�Ǝ�F�gG���`rJ0`�"4���}yLCbG'�Y:�ZQ��6�S�潷�r�ӭ�8�@��;�d.r�&�n�=4�ֻ�3�4M
�����}ٴ0��PV �ڍ(�ǻyL-�4D�&�۽#Cb��1A�߹�M/Uc���嗍��6��Fc��2��Y��ECa�#A��G'��F�H"{�0gD�G��� ��h#!�sw�-�l���;^��kCJ0�Q�{~�4hh���f-��f6E�UC1B�bdp�F�T!J��B��2sY҆��������n�;nA��`ĩUXg���4Fg��d1�mF��n�i5���C`C��2i���A�pԣ���ۦ#��_�܁w8A���ۼ�Mj�crn�p��&+ e����2Ͱ#Q��/�����~�:��t��|Q��CZ�kԽ�q��{]�d?URǢa?9�ux��ۚ��S��jq���7x��Oަ���?�/3X��'�b�b�h�|W�ޑ���#g���ih�(5]��S���sG��{�ȶ2ؐ��uz�KHS��m1��gy��<��D$��0e�oI��#/����?�g�P�����H�@D0#Q3u˼�i4���0���h�Dhƍ��Ò:0`�Q4��_+콅Bz��@ID#�����Me��20 _�̚h48�G�!�w��}5�L���#Gf/yF��k^�:��7���c�l]ϯ��֚Q�Ҍ�{��lV���ޱ=��ek���'��F4����w�4��j4�Q��;�wyL�wL�C����GkN����}`�Gkq�"n^y�ȱ���b�4M������]��\1߾�Ch��yb! ����3�"84�l�绽lCfw����Kʼl4T޻�a�l<��sZ4�%�.A��`��UV�[E��ﯹL-�m'��3sKM����YiA����{��M1���!�{���lCz����X{���:���Ȼ46����Zk�3��ƾM��J5J3��y�ح���=�3��Td��i�Y������Z��O��rju�*�/Uষ$kC�ޱ+����h���ZOnG;�ݣ|�[��\ɭc�H Լ��h�h�Pa��0e���iA�ҍF|s��`Y�����V
�%9���35��N9��߱�_����I 滬�h#�f��� i�l����{w�a�sX�S�ǎco�{J�u�01y���Yҿi��$t`��"4i�3�׷���آa�����M5��{~礷]��XL�	{��i�m������@�pC�n���0���~n�2�6s�kJ��8�;�t�T [/��f�uu�y.�����Z��;U����J���[|��_����x4�0#Q��J2���%�V�1F��&�۽##�s�ɇ����L��3ϰi���ҍF�j3��y�[-�3�����c�3DbG#�v6G�Dָ}�˳��\ �ҡlCz��FM��怶[2����(�ZiFb�;�=j�{<g���^0u�m�!�I�UXfQ�������܅��(�4��h���Q��a� ��3'T���Tnip��xq��1C��y�.�� ��׮�=d��nM��B�@e�LZ׻�L�뗎��]痎MZiF�Ҍ����ح��D#Ggn�4h#a�=�s�]6S��n��z�{���pl�̯_{7�����6�������^�F��a\���DLr6�Ρ�J��^�x�4Uc�@ ��K�5������_m5��?k�Q�*��ʭŶ��15��lyb$�! �0gPDy�.���t��q�h#!����-�lCj����Q�!��a{~�4i�A��u|އ�G��z���ڡS5B"�-3yyh{k���C{a��wJW8ܼI�Lk����ߡ�$n�1�F!���/!��F�����0���`D�����h48�j���]�x�̱���א.��'-�1�G����:�s?�q�06f^y8��쵹z�$�vd߉��b�I����N���Ś�iİ$0?�<{�#9*�|H'=�q0s����$�2E�GrV2����513DZ���H��0��-�uĝ/�l�F4��w6��ۉٮK4�P�z7T�#����eѡ��n��ׯ&�k��x�t� ��]�w6����AflT��K�̾�!�i�����p�O�|�q]3QL.��Iʯd!MV�v���vj,����Y��&l�9�F�� {����򪪹�����[���u�I���������n�m;K�'���W�v�3÷�n*���]��::|���;�����7m<#�\���1�x678�n�m��\Jr]�v�/�ݺT��.KvX�ٶ�TݗAηn�7i�=e�gǤ�vJ��1�Ӹ늋���+�x�@���4�1а`�����Q��.L̝͑V�T��e^r�v���W��1o�5
X��	]R�e���"���b�S�4ml� �J��K��������JK��2�ra?��� n,X���^�*�z�wY�t�I	~����mfQP�隄r�K�`�%ET��wt�>$�k0�
������cn�)���D�[Kpa��E��S��E�g�:��TI�}B�A��Y� ��&�������DV�����.|�s�Bէu�?���`�H�'~M_�j�ػu�~$Ϲf�|6/�l��j���F���#R/� ���ځ�I�AR]����v*������\��߸6s��ؤ�]w��{W,�	���.n d德I�����k︈NʉDJ��N��^���w�{�]����c���6֗�|��ї�3�~�}`�@�[��lc�&��(��v����x JUĒOwr�����&�Iɜ�4tB��w��_����&E
luۃ(�e���6�!J7P��k	�x}�k�������=2�D�u$��k����3>�ăUۘ0��	w.��	$=�{5ӷ�O��}� ]�H1��jť�!���~�K�&�/�3!>��`�w3!ܫ�d�������^�XD�p�5�E��ڳ�\���4g�_;�`����N(�g\┵B��͡w��a%k_�׽����*�]�I��$v���Lղh4��0`�~e�@&��5`7PM�����F�E���6\�]��@ ���Oo+�l������D����rГ2�D�B�0Q�s�iU��I��Q��ڀ�贈��&q���z�&�d��©�T�雝y�����voKyn��VW3Ir{[��r�
T{8�D�g�~���y�ߛl�kً'���X[�bH�(Q�z�.�ݭTI;�{	$7�œ��{}S1y4&�7.]�-���Kn`�$����eW)$@�Hē�8��$��b��k��V��SZkd�UO�`\�3�lp��)���=�y��[ήu
iqLГF�Uxp�,��ʬ�I=ܞa�D���+ �{���$sj�L�`r������"׍�v�U7v�2� D
�A)%B����9F󪛆��9�e8�K��+��(Wu�׻�6	=�<I��s�&/ O�Ԫ� �_rw�<���S&h��Y�Q��a'���	+6�ĒOjO�q1���19�'���².g	�"�ض5���V�>�{��5BO���}�j���>�X�v�7��S"&����ƽ�1��$#^n���#y��:<Tq�0`��wY� �U��so^ԫ�	��v'�N��nz��'!�.w��X�"�`TT�G	���<�o��'91r���B�DJW"/�Z��]M���UbuuĒq�y��qe+���Y�g}�]vO�9����E	�hЊ���9\�6MO������I$�i�	ܞ��	9py`1�lt�J�M�ӄ�XIZ�O^����O�sF����Jn�����$nOd_���JK�+���Ggy.��]sQ��9��d `���^` O��3g�]qHʓi�}��n�ԓ�G+RUnc�7�FI\�Y�Yu�gL��D��� ��.�	�ܳj�}��*�dIO��W�}����ѳ{o0-�zq<&l�CS�@�؅���G۩V��wĬV�]��}�H�����~I$�y��m��Tq"&���V�h�=�wW9�{6�'��pO`
�e4�;ԁ��yBW;�P���v8 ���ϭ8�n�f��nv�L�x����zu쁧^��w�[U�UԢ�ў:z�k<����z�i4��}]�u��-Nu����s7�6�.{�A��\lh���C\v��^Sn,�c�V��52�sGL��tӆ;hC�Ӳ&͐}]�oƥ�s��9+�>��'`�UU�/s_ɷ�;�Q0H����K(Ԯ�{ƥ[���B�Xi��q���'�[s����=��c�L�Q�I���z��$gr�K2ݱjE��s��֑b*��2"k��\r�gw� �v�]1I���$��=�,�{�֛K-M����IZ�z������t��8HS�I��&�߉���R��/1����3� ߒ)~A5mݒ���`��G`S��d�Ji]�O��oUԮ0�y`& hS1=n�w�[���*�0%��=�6�g�6�v�g��ϼD��̙�&hU`��$�_%W��sy��!ycg�O8�	$n�vMߕ0h�8:��_'�^�1Z�.C&�����W�ӿ��'��+������ �ݎ�[�A��R}�����o��vZ��<T�YQ8�����P��{4�kp���� k�J0
|��$~�����f7�$���#��w��I��ǌ��|IsQU���r��C���>'���x&�b*��2"k�ʸ���D��-,n:��I��mOds�j�]P@����P%ȕ1U5QSD`�]��*����ޝ�2
�U��7�${k��R�g���_{�w{����-ME�gp��^|Gڧ���Yc����2�W�ϸ��j�F�w��X�A�m��v�p�"�-���WyZI��0���D̹�DLЪ�+'�1[�=w��:�A ��w�$�mua
�d]pF;�vUwX5~r�@�`СF�}����lA'�4Uz�R��#9�η���|�&J��C�;��X�YO�=� �}�g)�ދqD��K�x�gt�z��L���R=���7b/��3B��^n�|��u��	��:i=�	ws�c��%�ﷸ{On,���nD��1I�"v�$��ʏAρ@�;�5��?aZ)w�x��~��f-�g_M�w���8�t���'_��l�y��m�{�ťpL�MR@\r�`��>+�������P9��3V���b�RJ�f�E�j�8U�1!>[�!3��B�oa��:f��y��J���V�����ԾÒ�(�BqI�T�.on�b(M���,0E4�1v&L�<j)�t/2����"���Q6O�L	���2[�}؁g]�m<0l�oT� ���*Yp҅���gnj:��Y3��l��^�����G(Fq�#��~���-��u^]�H�ʝ����}�1S�a�3ü���d������x�A��͢�q9��:FM۸�鐏<�����;��}���a�'�w���zv�\��vcZBr�섦4!>����vd��M���1�o�R��/��]YLF���t�Q�V�P,ܣ9YT��g�mh>`zօ�<-�[;լlZE=W?��k���iԟk�7�#�v�ؕ)NS�����
5AF�ۅ����6��D���+��������ۇ8��9�.�"��o�,`q�<Y$��q(ĳ2|v�j	2����"��"I~y��((�A�,$��AeB����ү�:E���I!!0�9EP�E�U$�H�uJʑ	(�*� ��t�O��aU�$�QTMH��K�Y��
�����3
MZF�Ia(EVQ�\�J�Г��t:e	~����a�G/H��ZJ�&�1�,�0�
(��QPL�5+0�BJ��	Ԕ5Y� ����e!�R�I�bHjr檁I�fBI�����CY��H&E�QjZ,Ψ�i�b
O�
�Hr����zIU)%�*֬�YT�>�ʝ^7.X�"�2�����U�����%�S����%����#:�EQ;0�$JHA���'���H;ׯk�gϾY����:l�9`�"h���U_:���P֝zs��g�]u�� �����M��fni����ز[֪)~�"_����#`��Ue�)����\I;�fx���C��_�0~[�8c��ћ�(@�۟���ǋ��{{u��9��A8����T�Q�uZ�yͧ�)������#{��>��R�� �H��vT�|�htr���M�E�'fX��""��X|��O��ˢ��K�$��զ�>%�+kr�Wvv���c
�12�$M3B�0��ۂ<H<ҡ~"���غXi���$�έ"�o*^R�@�`СGA�y�^3�뜴O�5;~��W�-�P.��hi���u��;�c���j^B��n1m���C7�3�b͢q��S:�ç�����������.�+a\��[t;��WDP3��x^�}��̏���К&�3UW�u�� ��_,Ð%dC�ڛ��-�q��j��@-�Y�P�Vz*v9E��"�T�UGj��<�]���v����.*��Hx�m����ٚ&�>�}àѯT����w��A �sZ�d��r�K�;&��&)U��$�J윪"E���#:����Q휤��W�S�q:һ�Imr��GUMf��gN�B��URDEE�w��A�Y��-:��d�mU��Kk�#oW�'i�IU���sqw��~f�Si���d�@%6�`$�դ.�i�=��g �z6�w��#J!b{~�d;:v��ܤ��d���� �y6��έ6aE���z&��xIE�Բ+e�V�x����OUN]SV�u"'}@`�����'�+CH�_���voG��䧰"oBK������UUUP�>��<)����\�-�a�i9�K��n��c��9�ي�Ԯ�d���ݸ\ݸ��o�9�ذK�;��f���uh3���/m�]�)��v�n�U6;�.�ˁ�ݸp��A�\�&NT^��v	v�e�X�q�� �s����mڣ�`�7ng����'Jmq���l���/�T�]�N�A�.��~|��1�|��Ke�E8�#�]��Uz۝�R/X��bn5ݮG�Z�rT�v?.{��R�~�����k5��mk�{<w:�٬���;T3w����F�b�տPd�=>kӍNΧ��aϤ�]>��H$9&��7:��#�7��fΕ�ys�����q��&��� ��=mZ�s�� �涳�$nOl-,4&�畒4��k^�WE�=����o��H��,	�+����7�i���殽��5�m!�ErUn)�3}$�*��Վ���`�8�`$�����3��l1�E��T���+wN�:��g;������]73��(܂�J�+����[+.��9�E�GU~��w7�i>���D�]߹���x��(����f�8�=+�3UY�ח`���Ux����Uml����J��;�t�
��4�l����V�p���y�lmȪ� �K�&.���3�p�+������m�AY?lY$��Wdg!-]h�g_1�f܋�&�A������>��w���w$l��s�ϛ}��4�M��{��yo��9EJ�q��n���3����/P�Đ	'�Z���y��'����W	�9̋�!u��&*(�ݷw�H����<GD�ʡ�W�}1��d�B��[[َ�a��]y�y�G:�[��L�� ��<�vx��o-[��rIK�-�Ygy�iTU�ESw3�I�_�$��,���v�P���2�L[�9�V<H�!W
�0D�ʫ^;scO1s�9�{=3�(�H9��O�<�,	��x�I��{ĉ,��@צj�1;˿F5���=��������I�����nc�[慨2���@^��!4r��+��J~�c�oI���Hϥ֍w�l�];����{��O�$��Wg���=�&܋�*���^!�ll�sj�׏Q �u`�
K��;�%n�Y�q�<��^'v���ƵĞ�}���h������n��ڻ�I%�Ռ���fɘ������d�M1>�(�5�&�|\r����5�K2KSN|R�:���Es6|��11>���UKk����� �|��f�꛷	���+�]wd�o��Y�";<���7V% Cֿ���ϯ�y�ͿVI!��AQ��,͈w
�=��`�\G4�ՠ�A�ߝ��W�;��Gf� �����Fv͓#с�,��JO�#���^�����I�Ų,۽o�ю���ܝ��Y<���5�յ9<o����c��8�w���iW>�j�]��
̬�˛po#rdMU���ݰ�bޓ{�����,d�碊�/�u�s���o��-�VZ�yf����]v���ȰO��kN^g=���<�ާ*r�ܒ��+̇Vv+������Ꮭ�>N������*qJZ�s�d���SE��n��(��A'�z�����ѓ�fw]��lgl߉ȸ�舙��5b�u���#t�.'���C�Y6H';z��5�+�R���{Y�g"�7V$�C�h�^L�ɂo�N�� �}5��O_��1c��&MI�l�z*4'�\��$�w���v|�6��1ȧ��������$�@Ϧj�3�2��@8��ˤ�����fCj0�3�l�O��$|۫��KLG6ӯ��*�7�z��&�uL���IU�;S5�Nh��	c%`����|�$|���J��wٰ��%�O�nq���:��wi��ߟ��UUq#��<����َ�Oz#���᪣�7N��n�w/7�Yq��ػ4pI��u�<\��ټJM�4�����\ݎ��r��5����;�<�P^l��Oc�㵞N��l�A�Wi�9s���6.���96��M�۬�Ξ;�w�Ǭ��K���/9�>nA�Ԓ�ڳ�*��)v$n�Yg�j�:�l�%�<��@�b�\�.��f�z�Ѽބn�O��2ʜ�5���APd�?�6���'wz��	$s�� 5=qkOk���.�� ����<:A��9�I�}��a0�'�v�ɚ;�����]X�>o0`��H_MGS�R��z.<B^����5ui݂I<�x0�H2N���FY��,�JZ��>$�\�b��^]r�벫u���|�ͷ����5��ȃuyVI ���a>(�l�;��~̙�'�k�־mii�͢8JBU^���� �Y���*��|㟸\ڻ� y6�` ���`���,��w8�3j^�ڎiN�����
;b�Fyyy������Q�Ꮑ�"}35X�]p �s�+Q�ٰ[S=4&�҇{����N�r�T��"��~k��}�'{~��*�{w�x[=க���oL�K�]�*uh�c�k��p�߉V�a��=���{�pO�Ƶ�6�=SMm�}�I$ww,�	$(϶l�J��sw<�==b&3F�MLA���cGأ�A�}yW<�;�&*�A �6�$(�ٲFEǺ�Q1�O|��#w��Bk ~�̃�:�� [�)]��r����
�';>���G�h`Ͻy<|�r6]�HY�=��v͂���к_s;�2��jb�Pt�D��F\r��S9��t�V��5H���������dul�G�=yy�AG͂���y���v1��̚mE��p��%���^&�x=�60��7���;&�>=��d��r6D�x�n��y���:�N*/�q�s��ߓ� "��� �Z>W>_]Yۗ�n��{������ۖ���}ધ�^�H��,�{8'��>=�T�y��V�4{��;^ݾ�\�-�M��Z���6�_��E�������K���u�K��m�8�̪DEh�MW�,�+�$��v	�y�Q�����3��\<��\\`C5��F��;�A'�k Ȗ^ꣵ��3l�dU�߉�_����œ%���_&���6� ��U�*�2u�fu�u��Qm�-m2|W!mX�)b��X.y�b5UQY��{�@��U�����A�{��?8w�`���dز�xD�����l���L9E�k�Cz�l�|�z�A��`�|f��s�W"tɛ5���	�&f�1���$c�`&��3W7�-ؕH�5o]�A��`EH&Y8"�LDMx��P������(�5}VA=��������W�z	��f�C��෸Sӳ�E��p*��dh�Ay�qf�*#�+�����Q��w3���ޫ��5Q�n�.���oolXSN"A���5&=����` ��+�����ee�$���	ge�Qۤ*+��\�^�{Ԗ����G���vb�m��pm�����7��5�������o��rѣUX� ��5�,�m3����3R�u��>$\�aV����REUTVa�l>=���Tt�i�m]:�K��=�+;(_���f�TX�׾'�i�͢B���^�O�^��Mw=��L���ٷ;�\o,�$��<	 ��ji��v�U�I-�z��?/jsyQ�����V� $�w;*����}���.'9��XՉ���U@-��_sZh�����^)�B���	qe�{�4KV�7�0n	�إ\$ņѾ��m�E޼���y�!*^��%�=�/�~Ȟ�{�F]��S�޸����vM��Z�B�\�d�^��1Bz��;ok���8�#R��;�g=�rpjW�_5đ��ĉ�=�Ф�n�s�;)Ybl���\�,·/�/�qW�wظL�'m�1_\�^)x)���\eI�2Q�v�#H+s)Ou���.۝=�����f�%�g��w��]�r̡\�����$�_��Eg�^����.��_��鏔��h�zf�N�p��^�\�Q�Y&�y�ѕ,k�7rb���o�0�X��;�O�0Ogg@f�y=Bxҵ�$[w�(ElMh�6$�C`�۱��M�y�ч.�s���=��_(�|���.�L�Y{p]¬�����ʿn�
�\�y�{ݍ
�>53_�<�OU�8',\���Tjb�b�*�����p�7�Z4E��:X9e������-�
�܌�mo�Q���5Ll�U�ߏ�Y囀�3�9��������7���ZXo��Cn�Ϗw��#�u_c����jo}�s�_�����tD����8��0�7��������r���W��;�y�3Ck<)����kt��;��x��x;�]�#����R�����~xWh>�̈́���:����%�E�V�7�z�w����jz���^o#r~���C�����'Tp����O���F|�H��
I��`dQd�(���y	��Q�_�BΕI��[Վ�4�"b�\Y���h�TYU֒ʂ�bF��_��-�Nj�!��U�Is:�+DUR�3jU�
RR�Y�mXY��Qg5"Դ�eX�����R��]T�4L�TP-J�M9)e{�J��D�Ys21��Q�f@h������Hb��d�f�i*���(�K'8�w3��QӥPFX�VK*��,��V���]RKP6K"���I	=!/�*�"�O"�)
|q��Т+�j9s�UE�E�.d���	�OR���J�r�UDP$!��DUQ�)��I�:� �6\.Q�ʸJ$���/_y�yUUUUUUUUUUUUUUUT�iz�u;�r\K�on���mDv�:8�s�L�K��s�=��[�g�>ݭ��h�&��TڵwOE�t%�8��;�|���V��q��N�,q�Q���c��.�ά�셷<�:��]�ɩQ��;�`Һ�vܜ�V7Z��M;��t[&ЮB�[�Ŗn`t�m���)"����k���;�ѯMr�X�'p[��'�����o�$7��w/[\�n�*ɻs�q�uq^q�E1���m�=��z�V��ǭyv�7�˃kN+l�{n�yS��&���%�
6�TJ�����è���s����{C�wn����m�8��m�gp�acq�v�kn����5pM���(���un����J��:���	�I;+���r讍����3Y�m���AG8U��8���7�Ku�]���ݚ8U����rz��q�V�m��u��aN��R(1���ۓۤ6qs����qΤf�������-l�n��t��Ƃ�g.����\k�7�o7;_��l�6x坺6��2Ụ������(9p�+��{E�mٚ����Z���e��M�����r�uԶ�5�8��;��˫����@<	��nb�-�w;�g'\�;�۴c�ћoku�����5e��kH�r�������J�sȧ�:�$�n�/l�Fq�p�*{�qή�k�#�(��ͽl��o=<=�[LI�+���'�5�j�M���)��:ѩ�����w����Ξʈ��gO�n����A�Վ�7t-ii���C��+j37>�WM��0g;��v�ƶZ*��������緪��ͭíZŬ��=�W�%���*���lx<��ޥȯif�D�>��b�
����u�n;Vŉ��υ����ml�i���r��'/��m0v@9�Ľa�`��^ׯZ�9ŻU�u���Qk�H]�����K��UU��n�s�.�"v^��p��3���:9���z��Q�5v@-&�&7����;n�nu�^�'e�\n�!�xۃ9��u��]��n�.�H̛;����؎k�7��i��w	���:�/\��3�i��:R]��d��8PB�F�//��c�m��\��]��]�/LN��<9V󮓵�n}���e��<�Ga�v6y�8�zy����.h�Ԋ8&��U/�v9P�;��?��"jL{P6�vZʲ|s�����f�WR�f�{0|6-d�$dvO����"f�]Z�H��qâl��xI���`�	��`��\�q:틾\���v�{�K��˘�����M��mU�A �q��I�f�$X'����*�'T�����'�ū{�3ܑM��ӏj���w�Ho��0rck��	p����h�v�V�N�'|�``�����p"��"B�`���vA<���޳���G���tX8�k�Z#��%�ɺpG9ۂ�(��
:ۊ��j�Z2R�e�&���X���b�#w]Y$9�y�����Vݏo��ɦ�=��id��ƬjXϤ����d>��gڷW��M��oJ;��fe���h9�������q(���Z�`L@����PF�eֽT"�ܚ�ƛR�c��d�y�_��Y$|�o& $��K�r���!�o�>@h�Ԉ��]b��� ��	(k�p^�r�d���Ao��U� s"b�DMMMfx�{���w2b�������� �Ϟa��d���ո��#Ȏ�b:QDEW����0�K9�b��d\Q�����VH$�<�Q�ɰC������G*w��>�=��F�zf�� �����jݔ��·u�\��J��ǭ���T_�-��M��us� �B�ݛlVݙz6¥�~'ħ�w��jD�5�X�=>�k�����5��3"̗z��R �@%�o=�Gn̓��zt���ń�� ��IRcـ����
+v�-�n����Q>}y�c�[u���k��+W�oq��9�C4�"�	�Z�_L'���+�A�:�^+kJr�f6deDG��;�I_�����^�9��C]�{�R�Aԭ�"'[�a$��f�$�oX��|�W{n�M�����y�P���ˮ�8��D
�T(�����7י�O�z�ǀO�͊�.V��!�������qcgJ��$�GXK5z�ԁ(�UK ��A(Բ���\L�3F��W��Y����nآH'��/�-	�
)�26�5�<|�n͂E�g$�DE���{[֛~DǠ�5�n{�g��A�6I�ޫ"����̾��-��H�F�
��-����\�i���V�"��MV�)��V�A
���n��94z$^�"�b=b�s�`��/D�d���� �{uU��y.V�P��2����r��@��v�9��P;:�K���ai*~J�-��<�86�k�X�/�cg�*�S��Un}��K�ڿ}s� u&�U6*��`�	��&�o.WX�ة��={�`�^�Xs��Z�\m��_����ۥ>P@�Z�H���ޮ[�luj�3�_e�-��$��5�3��RWBYe[b�$��B� ����wowc,b�@�S�$�z���Q3 �S^�ӏ33n�M��+$�;�ز�bi�fp�\k�v�c5	��_��뺮��	���^x�\�Lf�Ή�D��}�6�~���d`h�P�~wמs�s5ڰ_>�>�m_�ە�r���WE}�� �|��un���?�ﯤ>�nX���T�$^�v �m`�x��r��kd�΅�c�W#�f��})$ɑ	� SW{�p��P�}9�ip���2_�p~����FD�_���m��m>��}e���Z�L��	i�em�y�ݞ�����LN��ی�'��������1�ug�7=�=�;��b�rnŬ5��#��^7=�v�ϛ!&�Yƽ�륝��.����֬�p7��p÷c��]qr���x�GN�{3�hI�6ˠ�vϭb��y�I3��5����A�Wn�z�>�9�V����z��c�P#vZ6��.�9Cq������S�È��������ۿ H���zm��	� �\�	.ܫ����LN��ۻ'ă���|�Ls4Ȫ1555�D��A;X݂�mu�fu"A$���fI+�j�I�K��=zx'"a��4jMzʛy��}{vI;�u�;��	`$RM`	 �ܫ�"���0dEzfj��]B˙�oĚ��@$[��w�;�r��C��Ǟ�ꉃ�К����wRV|I�ޠ��VVt-��P�v�/%��X'�����X���}>��� ��d��X�օ$��|:�'ʫͮ�Jȣ%�[*��g��/��W����pa$��j�I>�ޱ8o�˫W��&��)���u^Ւ2O����W��]�L����렠dt]Q�0������0��A�I�o[�2���Ե�ҩ�QhX���5Yȱ
P��%N�9K�ҩN��r�H��U}�B{�`Oۿ]�n@KF�P��]�hu�̃3&��MUf8��d�z�Y%���n�#��ᗭL >����4{�µ~x>��Ӿ�]����}7Jş�@ת�9.Qh��6g�X�K�T/�u�d�jL����1�Y��s�b!�^$�VU�A!=�Iir��UT��[�w{|���U�(R�H��G[E�X�Am��['\�x�btNZ�eNg�1��r�Bߟ�k��O ߓ w}�}�2�g���꺲A>ڬ_�MC�j��1��o9��2 Dgn�Y �H���$��g���GEͺ�'�ό�	�W�»wd��M�c�eM�d).�CT�D�^��Z�,kN�eY5�E�X�"�D��̹�/1n_�d�dB�ʅ]���uƗ'���	&������^ �ls2̚5U��z���1�$��W�H�@ֹ`�AZ�����^��~P��"5MMz�Sٙ���v�{���0�t�睋�w�,��v��19��.rs:��#�`wQvN;=G+r䌡np�#�yqo=��K�j�Yn��qE���-Ý��g��f��ڰF��@��r�Օ�~$|s��qc�cz�e���?����V�b9"w�H4�{)�I�M�H�Mx�6v:{e�')�=)O,��q�:��BMD��7�ݘ|O�KvŒA&R4;D��>���@/�<$�ݫ8z��	B���U�]Q{���J��N�-�>$���Y ����x[���4j���Un�v�>\��J��qK��zo�� G�,&p��{}���?:�`Z1���RY�b���b�����G��<��iwB�+RR�Z�03��&;��ɨ�2O���Hv-��}��`�}��6�����+m@��V(Պ�J���e�]���d�s g�cLR��Z�Muy��tr�;/�Gg�/�=�`����`��M��dU�.u���,M�����M��x⋭�1�j� U�bͱ1���ٮ�3�Z� >��2O|�\h��*]�D�|ּ�0`��Fff����j���N��Y ��U��3Kz�U6	��*���`d�~�U�&�c�)�th��ڳ{E��$����$�j�Ē|�Bpʯv_���&6n H���%����� rM��qqtC�W`���X�J�W~ ����9rݿwn�x�b��V�Ny.��(Y����V��I3��mmE��ǂ����_���Bz��&҃y��E��~�m��i��ە�hW��n����ؗ/�/������U�&7#no2�='9�ɮ���s����96�.qOQ
3��kv�m�Jr��u��=��]�b��m�'9�u'FKk�W��{�/����Z��;`�-]�9(:f�|��7;�M���\\8"���ܯXVL���{�s����{	x�Qmɢ:��ƙ���c���נ��8�׬u��W-�<�ۗ�8�h\�u�-=~~w����LɡQSUY�Y�zρ9U�H$��7�����J��A���
������S^�zm刍�pñ.��������>'ǟ7~��aʸ�^����M�a�#��115Y��X�q�y���Cގ;��j�j9v�yX/]�Io��Fl��d�ߟݞ���b��jr�JI.�(\հO�%�e-���-�1���5�z�I����}���ĀBŖ.�[��T�>x����\݌���f��ʚד߷�K\!SvW�����h���y�u��(�TQ;!�$����� �*tV�um��$�I��A�eY����8e�cu[j�U��y����3&dШ�I?��V{�."�����<�ŏn��س;ϓ�[4J�G��������^,�[UC6:F뻔�:��3~������U�%}��0|^}�,���bc�.�ǃ���sϑچ,KW�=���y�hY���iĎ�]W��� H$��ı?��{.�mj�8�Z� ��1s��95�3�=s��ǭff@$�����oT^X�ea��M�`��{��ص�Y$����}�-6���]?W�[���^���幀��wU��Fv��Ϛ����ז���#�FyUAF�ѝ�5����t�V��/#���>��bt�ۯ������^h��ox�{��$��e�$���vA8��<�	]�=���V,�'� B&W��]�$T�ŭ��y��$wU�{w��I��cn���W$3hj��G#��[u�5;��i���w˦��Y �SW��v������_{6p����s�X�ݰ����>�7��g�W��݊v�tc���&FF�;�=�*'�^c�}�g���UcoeX��=���ڮ�Pd��[����/�,מقo[0,�� 1O�h��!���`E������k<�U&�F61{�zd'� �tS�c����گ�cH�%s�mD�T9�;6���QR��f���9�Yf�y5�n:+���q�lٙ4���lBC�O5w����ɻ��N橅է�F3wI7�������g/�;_�'��I&R�>�%�&��AZ�a����U�;؈{nk[����xy�uf��{��lT3��K�m;ŏV�j~�*�&��p��g��\�'�/�o���ˤC��uǢw�y���\m:X��d�^l��s�n�5�I~�.%��t��;ن�5�aǂg\�@ɹ:��-V���w�Ȇ���.�8�Y�kw�!PI��MFET�Bu�g�2AV�����ٹLg�'��j)�Y���TdC�Y��
�Q��ā�&��=-k��sF5��S>���1�g�d�ƶ�rO^�������{O>99F�ů<�K.�ݝ���cN���in6ɝ��+Lc�&**l���Ƀ�>��gy�)8vl��,x�����S���뜉�����T+�V�w��!6{=�xG�i�����hBf����+[z��bM��m4�6 �cR�
��QEI��!a"bEJ�'C��dh��"�TTE�QkT(�@��=�.���	��UE�T�<�̠�*�ՔDDVX��ʪstVq ��.p���*>"GtJ�W�/E�kk��T4��D���-K �[�۴��\���^Uʔ<�j�y9YʷX�dw�efr%���?)�Ȕ�fr�̮]>$�rrrT���.>^p��]�������s3[/�9TETWrTJ��-��L�rr5:�*\��NDՠF�H0RB�'8섛��N��<륗
*3#D�3|3�Q��"��dQgǕr��<ZT"
rr�K �r�D��i�ꉖ��UW ��P�dU�Q���R9�"�y�5l�L�]��?�5���I�U�	n�v	���M֢�Q�~�~����'g;�U6��rŒ|H����O��3:�}@Vu��[�#�@!-��u�ZM����g4�½�\�.ʰH'�U��K|��]��}�4�������Imq�
_>ӎw&�k���t����]�Q7���7}�nʱ�x�\�$�� �|Յ�/��k���	׮�2M�SDQ>� ��y�&\,�ZEd���%�I[��	<����,�X0�x��q�jC���A���^���I$�M^|wS�m���cf���H9��� y�Y����3��ۤ>�gwrmo[^�2r�&����I (��W{f�z�"`��X��q�)�^Ww������^�?��v�.X�ǻ�9Z�ͨr
)SU����ILx�������>Gj�,D-_��o�0��Yϲ�Yq�9���<8���� ���Ĩ�ɳt��t�K�0��u�펅��ע+��:�ɵ�Ω���p�zخu�,�Tw��r(T�3T�.��$q�Y��Tglߍ�Ď�U�&�^���$�w��}�B`��"BQ=$�﹪����評R����^>Q��`��ս��l�[`��ؖh�Bjϳ���� ��f� ���:3�a�&Ay5c
9�7�"`�P�&��biu��]B�=�&泳	�{VI{�\�2[���muŵh�u��Xޘ�311B�*j���(i窬�₎�{s�2}Z�fB�ڿOn�ټ�ic�SF6���W�6`#g�;�z� n7�G��M���9�s��<Sܘ&�U����@�՜̝�9�����׭��m��P��!pI���n��G=(g���[unݹ9�v��=v[��۳�۷�g&�On�p�$2a���\I�2k��{q�qׯW�kq��=��uK=��U&3�D����r���;aĀ�M���ѕ�/]��wmq�2���1��9�����j6�����M<Fz�{�Q׿�|/��Mz��M�z�i�k/j6�����y�/]��:�w���=n��=����l+e�.����R�;*\7�}�?��޴A ��fN�޲8:�Xo��� ���Z�ԁ誱2Inb^�<��F��z� ���`�^�]�O�ڞ�s�/6��`��"9,OI5��ih㛽B�."�8s��n�HY�VH$v�X�d��hMA��a�����S��*vL��kl�[͏�{��r���������9���BL��E�4��I���Uy���r�~.����y�0�w�?B,�~����M+��� .��WY�<���A���y��;�Z��^�N�e��Pl�D���
���|E,�	窀mv���:��l��VO��앁���Ś�%j����H0k�2�����қ��{��1�k��nxDo��VX�/��գ�۷;H[�3Z�I_?y,�����Ŗ����T�_�<û�6��9߂G;x,	���]�}�_+F2^��nzR��u���u�3�P�&f�۬��	ƹg�����%��J#�]Yk{0�L1٣fjA�'��B�뭐���X>/�{<��M�&#�U���wvɡ�!&����^�}�(���TNA3sL�}7Ww��mv{�|3ۊh�'�j�1
Ϥ~mGmv!�	�6t�2���ܑ���y,v��b���=~~��<�&��5^�M]�H���	Q��`���<m:�³+v����O=�+�\ѥb%jS4yˈ J��5��)�b9״�'�<K��� �V��*���K��S�D��15�:��$�}�,��1�a}yX\�����:L$�ܸ[�G������Ԝ���g�Տ�5>C��y- �M�Y*@�ONѾ��(E�*�L!_jt��|Wܺ�������k��>�Y����Rfy}X<]�.�F��~�~ P�u��>�]���ﯔ�����o4�����
IjzI��rX'�sz�8�V6��6�E.��$\Z��}��vZ��a�7:�T<h�DqrI�<�M�u�ƫ�������L�#t\���6��[���Ď"EMA3>��[]�	>(�ٰ	 ���`�U���]v��I���ތ�0HRhI�U�K��'��Ϭo_([��id�$���ğp��1��Y�wm�g�.v��tiX�))�_�0z_�  8b�<I��~�0�� ��+Hq3�Dɪ35�=.��c��r��!xim� �N�+�@'ǚ]=
8tL�Y����Ȗ4&�-Ysڍ���ݛ�ϵ�&����e����,y얋t«��1�UmEN���U�A8Xa�����=�$8��`�t\�}"��115W��n�H$i}�0]���R0��w�~'��r��k��I��	YMxڶ���2��0�5e��e��]�6ݒ�m�*,tNJ۲�k8��qz��Z��]�_�����W�I�\�[Aq����s~$�Ud���b��3���;�a���LW���Qf5V	&���k��b��R�zt7g$L�D�zlR�b�y���	�V�������d"Fv���Jk�b����H��4"*���f�3���~�0j�L  ��t����� ��_s���{���&��UQa<�I=�.J��O�k�X!���A%omX��>�.��[5|s���51ѻN+\�)���J����Y8H�K|�G�=Y��}1��x)V�y���5�$�I#�5#���۔�^�ˋ�w��e���k�a�eP��Eo6`��9wkWo��b�8����6 k�!�ݪ�\�2����������� ��ۮKUv�`y�W�����.�3�<�Z���y؛��٠AN�4���.�T�j�б<n�x�󸌽���qqs��ls ]��[��Q�ɺ�TFݧU�KgR����7=��Z���FS�ݹm�ty��zU/���s���=R6B[���oZm��Y�����*i/^t�t�� ���1b��FG��d�=5��k�4�p�x$��ojϏ����x�����ZB͎�;'�D��*�3>��|�0Bյ`�t(�ؤmK�I<�n`>$��'���� ghY�_��\�iퟺRm$u��$�A[�VI/7����e��O�k��<��;������`��S� �{��j�a�Q�dy�㼶�Ēf��2��w�s����jQ[]D���?��u�s�]B�[qw<'��
�j>�߫��%��>8���I ��߬�O�o]�:cEI5��=���[B��W2�"bj�=���`�8�l�Xc*�LB��'��(��nkU?n�Ɓ]�Xf/.^����c�T�ĕD��8r�9:�&k�eEꊦ���rڰI>�߮�I#,����hW4�0L�"fxLEL�d7jş�ޫ$ᾍM9�.]��A涬�ٽvH���d9�b��3�����DV�[αm*��=��H'3Uߏ��j���S��	*[��!E@PHRhIU�N�ĂA�om��3�wq�]S^�ڭ$�;�v	'��.��[3��B������XϠݭ�llu�T�������|O�rA�֪X�|���8�� [3ɫ���o��W�|I:�n H�8��o�t�]��~�n)�5S;���<�ښ�6��|�#�mز7�n`&{6�ec����m]>jN[P(�Ks>�����H�]�0��u.'T�]�gEtة�rl���V"�h;9uB�b4gRyU@�N�g��z��{S��sZ�,��d�\�w�#�|r�2����_u�����vI���&d��.� ��P6x������ �n���O%ۃ '�nh�Uzr�o�19�[d�1�Y���F��U�ol�&���z�s��:��z��x�ۧ�rx�NG[�V)$vDM<͆�WZ��	�q���pH&$�LM�����9�����o���-l٠�F[�U˝߉��� ¬gPd���UGy��wN��6��J�ٔ>$w7�|=�X�/�O��=ca'��-D�U`�y���ǖߨ���ً�Sֳ�i$��������Dҩ��T*�����z����>w�y�T�p`���X g����|�S�id��dQzLY�C���a!��ږ:�d����w�ĦvjS9~S�uۈ����,{6c�����ٙ����o|�w4�l���J;%��?R�	9{�X.�G<R�o�X'�Vf	9l�>$u�]���wj�L@�4���c�`US��kF����9���܂y��7�N��
X�,�3RLO���}�I�Җ�O����R	�������:���GG-��΋�0HBjH�5���A|^vYS�T�z� �)��`�w������(��m��{�Ʋ�zD����y�e�ȳ��*�Xwi��)ʕ��g��̝M����o���UkZO���1�1�:5�]� �;ytA>$=�vI�"$	>���2�`��Q$:���^�%��I�E>�����H�޻ �	�v����0koM;��'yaY��s��/�]���>ػ;ZRĚ|l+����aT���%-�T���G(����mą���:���ֈ7fA���xv��*m�䣺	�{=����nN=���K;p� �V�"�f�:�fv	I<���u��o�l�F�t�^{�q��}���I�[���w=�ڍf	����d��������o�Y�ֵ�ֽ6<d���XÏ؎��eT�Y�WG:����Zu՚�1�>��5�1蛛�X���s4�2�RD\�J.��v����b���.��'k�!��V������'�f�"A�^��ܴ�B2)�0ё�(ٛ3P%�y��X����W�^<d��^�z��{R��=����8��+/��{���9�k�t��a�`������3c�������Vn_f�B��Ѹ}ݳb��`��]�	�_y���{Z���-������&��X�<��ȳ0��Qj��$�(M2<��r�Y��ۛ�+z���
�V���\,�nZ��L���h�@Cڏ�zD�S�GN�o��֣i����oY7��{g�=8��r:��}��l�ʎ�S�e�ٗ8r-c~"`K��<�ײe�T��jo�Y��.K+�EJ2��y��W� ���{�[ #�e{�ƺ�G�NF�`D�����V��,�ƻ�,����V'��[�l�^XݿMM�˖2*�[v�����01��:0J��G�/���=XEl���{'�o�1n��^�8���L����5��TAp�jY0���8R�V�Р��Ns9Ay�u#��E�	�QUG�ȼ�I�;�g�ք�Z��A˔P�:���J/=��k("�Q����QA���{��UPQIJfs	l�S��We2�Q�a*Uȉ���;���wI�
"��
�jr�,+��w�u!�ͪ��I"�ċ�wN8�ww
wFY��L]�=@֪$�G��V�S�	r���)$��i9�Yۢ��;�C���Q_)͔s�!�A\(�e%ETB�qV�\��Qw�É�%K��L�w�*��I��(�*DJ��N�Ӊ�Qr�*��qx��y�Aj��?��檪����������������-]O'KƦ�Z��rVwX���na���sӦ�e����h`��:,q�ϋ�`^�D=7:n�w<��ŬW:�׃�L/m�rd#Z�]��^��q�I�
�����.�h��25u��v�m��뀎�s/p�vM��ƆWv�;�ay,<�9/gy�Ŵ�͹%�;&ۥ9�6�i���շ=k�g��Z�N:��j\��[�{b78�aq���+��{��$Vo5�kk�Zyw�'��s����l�c�#�s�o�����v�k��t��6<{g<s�.Ӝ��7h��t��#ճuS�؄o%�vk���Wt�+��k'X\��u�l�$�{Ae��C���=F���������pp���Uq�m���DX�<�Jݒ���{n��G��9����{fd8.s��<����
�wa��y�S��́Ѷem�v�$B���mk�=�Z�<ti�' F�����v��m�ώ��X�v��F��ۮu�|lAGc�;c˞wV2��s�cu�v�9�5�^���Ū�WT'81ٸs�����Z�c�ԧhw�8�&�ǜn��K��lv�O'�f��ۺN��X��nv��s�]��]{�Hv�o>݃�zm�j� ���n�o\��vy�0kݽk>J=p�џ@N��
�KGU�� �R�t���t�3���[Oi�8m��1���2�}b�J۴X�>ϡhU�ۧ9������Ov�y��ۋ�\�nݧ0��Z^(ojݸ�B*nr��ܒb��.ͷ#Ӱ��3tݯtt�o;�+ra��:[/7e�I�A��3��Y�g��`��i�M��"�=��K���Jfg�Vt����OO=�*#���hv��� �N��upO���w%�.GN���'Px�]Z�"n������f�d`��f���\H5UU_���UU[��v�_n��<��y�rq�.D��tv�YKV�t�/Q����]ȵ����r�;N�xq������i����׳�駛j7l]�u����z7X�>��e�Ჴ��,��8s�ݸ�.;^�=��S]@<�+������;��ŏ�Ɏ�0�u7-��m�i�[���1`ی�;
�'c^�ѝ��N���V�ku���uC��Z7O��쉃t�mN��5v:X�V�o���o���ZIk���/Ͽ=r�аI#�v�x����Eq�S��HK��Ψ�a�&�jI���|������&4FM�OS�@!����b��r.Z5}�851��!�4(��E�ۻ>���H47R]g\� O�MݐK��x���3B*�h�ow�3��7�g	��X$#��fH�{U����H�]v	�Lc ��1UDY]Y��u���'d)��ڤV���O�WfՂ&��N3#b��A�9ir^�;��͝v�a�%:����<-�+�uٵ�Fk�.h�I115O�]{vI'5��$U����6�v��`�S���Smg�����T���jzMv��Z>���	`���:u��ҵ"0tL�����ҕn�O5t�Ƀ�\���F\�5�qݿ��;��Tl+�Z>��4����z/� ���	+�j�:��_�w\T�D�*�Ϥ��P1>��������d�kU�ݨ��6qՕQ�z��>���`�I�Y�VHΘ$��4DO��*�X9Z0MD�A�v�a��^v׬����f/.zj�&s��C�u�dL��5S4s��4Y#���FF���6�@�噀�7;j�H%��ߏ.�r�'�rf�A(X��=GC�(�뷙��n5S�1d�x7I�5m�й���;YT-�{����ƛMw=�zω'�w��J��ӱ92����I+O�{@����t�Ng�u�?	Z2�b�8ҝ�р�
�ڲA{�W�Og_D��t�ц���,�-o�uR;%��^�;�Fn�B�	��c]�+���M5���]YEv�Z0���oˏ�G�X��;ũ�1}��)w�| �a�����᪻�n�&�%� ���`��~��9�
�MD��1>�4��1w�1~<�ذH-�]P�Ih�H�J��遂A�F���L�Z�6�a��-���O���I���I�fdK{�^T]i�!#r��[J6#Ϯĺ��\���5�Y��wv�f�����}.Q�������g����^�Ck�a���"3e;��|���$�1e'�r��[Z���f,>5�cgq����AKU�$�y�X3 �q�$��}����ѹ�AӵV�e"A%��I��g�f��X��Jk�ad�3��b���P>s�kY9�dL�H�uX'Ă@�������YS:���C޳ϳ��s��X"ƶ�߄�����x�wp<�ͳ�|�X�g3y_(~n}�.fz��ݑ�o�ۄ+�`�Y�w��|�[�Ϧ�fh�f��簟-[wP�����ڀe_P�3�,	{jΎ[]����O�}������ 5jezz�+���N�<H����Gֺ�q��Ew��G�*�=�[\HosX0��J�ڳ����?]����$���aVNqf��*��^}��]���Ǥ�Zf�k��6��ɬH+{j�"�������� f���f�И����w�I!�m��%#�̕6ன�LN��!gmX3f��j�E3S|�)��=v�6'�nfH�[W�|H�޷�7��{���dX6.�?�;v���,g����	oU�9��{;{4t�B�]�H$�vՂA#�z콨�E���y`�"������#� ��o��ste���TR������_�����;��g���T�=]q��,�r�m��F��4�bjWR];�|�*l h����[�#N� Y�k��\�j��m����ѥtk7g��sٮ3���i���;`G^�Fc��}3��磒���Q؝ۇ��N���=c�1���a;]ճػ!s�Y��n�^wZ����w=��q��y痶��t��ˮݣ\Y����=����6}��d�Y���%Zu����!t;�b�Q9.�ƾ|~v��&S���L���nf��}533@�z«k�	$-[bψ#�z쮔�U��U���ֳ��{�V8��A�U��]R�Ov��nFZ��	�;��d�{w�� �a�7��t�f�N	�4&�f�g�ǻ~��U�I9�)�銖���[V	��X��*%�3BhL�T�1�3�jO]����A>'V��I+�-�X2o�"ҫl��Q��fbjo;�%��{/v�/pɌ+A.{*�$��V	� ��g�!s����U�jf��J�X@TQ��8���1#�N�GA�Mݺ�e�<�Ė�`&�|�;����.��j�h���X	�ޫ�r�e(��I�<�u�V	�z�^:�H�Q34W�:�la�4;1���f�V��p���]�A�և�e�����u��f�o�'{]�\�t<f�}��>�E�{0����o��o�?v�	+���` ���nj��fo:��O@� �
��D�&S��N�k0�A]ъ^S�n.�U0I#wz�Ir�U��r(L�Y�n� ��p߸*'� �X� 2����0�uM�~o�C\x� �cl,�&v��B&j�Y�y���-�|;� ����ݗd�|s[Y����mX$I��������5U�Ȋ��O���j��c��Ö=�=�%�cW����?J-�s��lY��a �|W-� 㘍1M5�[�`���0�"C��Bf����l��W� �@�VC3�y��s�^�H}ܳ<I><�׌����\����[Q`��*ff���aw��a��m�dL%��[����dd�=� %�L�#�:���J�[��~���6k�ۧ&�[ײ.E�ԍC�j5J���>
�ē��$��Ղs���T�xϢgz���`n0H7\� �|H:�ՂI�޽(�{�; �|ZWم���"�ɚ�U3Q��3ݒO=T,[�SF�h�|�vfx�H/���~����^燷K�����jrV!��A�ġh�m���jV�i�,hU��l�q���1BhEMU9ffHZ��$��`����9�'źX0�Ud��HO�j�ə���{v|��73%�ʻx0�	Ud��;s��O�k��2����xLQzM����%o_5;��6�o=t�m�s�Xb�^��q���|IĶ�K�볝Q`��*ff����.�خѝycUh�Ă*u��>K�$�˒��dCO.}XHn�g�뛁�����:ƍ��o���x���qwn�۽�S�.e��QW��(�fh݁R���}04H>�Rh�>���4��6�dQ�l=��H3��,�.�w�A>)�X3�dKkv���Ӛ�(�c�T��,G]t��ۄ�A����VB:��R�|���EQ��%3��v�d��T/Ē\�F^d��a� �T,�Tٓ=SPh�����v�bqg�������>$�t,��,�I�Y��L�-�u~'�B�HUDԈ33Q��iH/W,I l:���ՒwuU�J��0�Κ4MTMA�W����LneVe�Y9��`$V��ݜ��]�'�f���-E��ыwu�מ/3� �Z��c������b��u�X��m`�A{j����7Ύק�=X��*���u��lĎ�V79����n6⯞����Q|Fgc�ۺ�0J�Rb�n3fd8���Oy_{��UUUUR�O��Zq��iAS
;cNx�h����b�a��Z��f�ki�h݁�7.�9�6��r�n.�zo���FN��J`��6�w�Z+�Mb4�c|�����;�{����7�q���C��..�Q�u=��ٞ�n��)�`�۩��m��V��7]K�^��O^�=�s{�n�ό[�����x�j֠���ݞۖ0��s*�m֞��9�a�y�&�`�Il�����^Q5����go�m6��k0�{j��4�О�O۵�߈&߾�3���jãV��Q�OZ�W	�im��� �u.Y������3����}G���㝰(�VYW��f^<C�ڰI�Jf�_M�d��I��V�Ղ}t)I.���"fj39ڰ�E�i:�I������ՒOn��I����޽s���[&ʥ��J=5��y�~�������'��? >;����n���\�sQ��̈���>v/qם�/m=�.���2�-��I���}sGm2��)�`��""DO���NŒ|F��ߞ��訜x��ͼ�u�{��0�{^Ճ�0I%5 Ϣ�R�A|�˼yQdL/ٸOӯ<�산^\��{��3F3ފ������-Ξ�b���iǛ��"+����#���en���ɿ}�	$���W��߮�I76^����e��vI����%���'�x�}�Ɍ ��S�v��T�ǨC�T,��`����(��vYV��f���x�m5v�Ǭ�|{�U�I[ܞE��5�x'�*�t)I*����35�m	-.X0Jk������	���%k�d0��wf�2E-8ݴn|Z*��e���Ɲ���p�j�W%q�K.uup�*��]�?|�o�b�#7]Y$���`�7r���.t�I>��w�Q`��ELԃ5���9簜��6�V���}��${�~�J��=F{� ��v�/f	$ˈ��}+�A$�\��$���ń3C�x�}�vN�F��%I�<K���[Ͻ�`;���oy&��w�"�K��A&�B�>}�k�}���;f��i��4�f�wLl��jhYc2+t�ԞӫP���.���&���w�=�\t2�i�| �AI��n_9L��x	�����~���tYrݼ9�,��fE�X���%)�����t'R�USx��	n��\I�[����#���8ezTk&�s{������w���r˾�k띝B�|Q�ݳ�TB%D�d�j5�`��2&��R��������}!97;��ٻt�s9��ꏴ]x����Y��S).NI�Ε��,M�vQ�睂��}�o�L��B;��x�� ��o^�z��غs���$�B��O]rUֽ�m���nʊuX�d*���t5%�=�|U�G�h����E�x`�����y��/vw����'3�5���l�f�ۤ칓6�_p�}#�bGb��f��D�򕮌m��9[[,�a�9��)R�%Y�#nZ"�\���4b�����OچY��8�s�ac��s��[6w�����i�ÞsM���9J��X��"�<���^�Rr�&ų�H�bZ ��G�sh�wD}^���զ�A�d>�rM��0 Q'�� �j[�Bo�w꟬�붛N��NDj���5	'p�b�෸������X۪���H�"2Ѥ� �Q$!t#�h���C�̜��L s;��Er�5*��A$[��|�:<�B�8!½\�F����
��W+�9��x��3�IPR����;�Μp�Q�\�T;��$QAy�t�ʋ�A~����:�W1j+�=8Trtw@)���{�yi�2��L.Y˕O;�fr��*��:K�Q%15
͔�\�IGq��T���"t4+��B�[�[��ۘG��*��YJ"��s�i%z��#���"L��a˞�r�r+� ���2������iD\�\(�mX����PQ̗D��.]$��S�"�W.��vU+J�����.�9'=YNwg	��U����J"�:�8t�r�gS.����F��	 ���O�,��I�k�d����C3��SVQ��5�5�������kZ�2n�P�O��� ��Q�s��������s`gH��aD-Z��>�� �yX�����Ꜩ��]��I�+W,�I;��͌=��/V��p��ET��ڻ#z狶N��˱���m��=
G���ld��?\��(ED	��|�˰IW,��H��5W9J&)�]Y�d�w��aD��Bf��SRl��x��O��;�V �ɬ�|I���%W;ƌê� �%q`�>���U��|O�VذA[�'d����)6�'�w���8$�(�MP3躮v�w�����^	+^���Go+fEn3Ww��i��އ6�N���ٜ��j�D:i���+�����N꽌?y��h�
�qۼ�R�ee��nVK��x?�"q��0��s���ËQ�PJL��ּc �ܘ��ī�:g�ׁ$��ʬ��c9��{^[���<�S�\n�]�QYIT�뎻f��8۫nH'��
�h+e��z��򪢌�_�,��=�vA$��X�ʺs�α�=:�2`����b��
'7u3���y�ՃOn�a�A[ʬ�	���q�]bk�K�'ٹT����O5`���$����vwmTGV��H/yU��ܕ�˒L""&����`�s��3׊9��"g�� ��ڲ�J�H+{�Wb��W�{]_�H��H2�D�>��n�H:���ʮVz�{VU�����$���2A�y�C���h���M�oƩ�����[d�1�4�mE�]��^]�@�܇|�rb6��=�Q;un�5n�ú�L#�g������m��"��6�+E4Ы��q�MPm�G+�u�u:C�Gn����:e�;�'=�n{���f�n���ۮ�z�N��wF��M�˚���w^Δ�����̻��u����X���4#�爲l\�@���W8�:u��W ���1�����F���cY��\ct�E�Gn5#�nMшњ��kS�]�K%�3[i�5e�Z�����Î�뗑�#͜�	5��GMf�TQ�x�[�,�H<ҫ>>Z�f���\^h䶃%kW`��h��� ��=�� ��d�����i� }�{���H{�0`qj��ߦ�s��1 ����V,(���L��u�����s�s�\\�w�ˈ��ڻ� >3��f���&�T�7*%�Z���if���{���_����}�`ӝ�����V�������G���8��K~x�M{�W "�B�*�ǎ;�ꄷ�DG��fdDDB9;�L��'��J�	�zk�ŭyN�*�\��s��SKl3l�%̊t����;v�u�=�u�����~�ډ��5�{4����̸ �O{��n��˿q��\�-x�{��6��{�0�z��[�T��A��e�N�=��{{�1Ϡ��F�Z,�w֯�&b�dlKqc od>�N�l>�R&���<��nՈ����@M���W����SdJzb�s��2۽�Z� ��ܙ� [�ꮐ6�����������!6\C7رa�
Z��3�� .o�ih>�����×�S~�w�@ zw���`	�~ҭ�U]�<�aD��d��u��:�H�]��ހ7�� >�;�t w�ɜ����ffo�9���ߦ}��*�rʬ�bZ�����<x��I�M�V�|�W��}�;����f7� ���J� ��fa��o��[��7S��+EQ���Na�������|�ݾ|�;�-h�K�θ����~��sX)o�M��rk� �ʵ��>�����o�n�'O���2E�x�3��}:��LF��f}�|�ôs�_�6\�P�$��&I�O����!�9�N���>}�;�m�}��ۨŨ�($�b�YY ���9��I#����'�����`��r�bHl���ɛ�h��|*�%2/�V<�]7��s"j�,e��w�?_`;�1����b^7{R�OpZ�~4��ވ$=�b"A�~�̈�+^�82�q�C=�Oz��%�q S��K@��sZ� ��'�Ms3����$��oJi^ǲ��t����X�	>?{�)�&���a�I��X�����2�'#g�M���z�Vf�괮8�����]�]��G�-v�ö,��7"�ĖኧeP�:��*��m��[���hl&_����H2��v�&�2���*������30wډ�:Բ
[��L�q+�NNv��{Uk۫�Cb@f�����ɘ1SZ��.m>L��+�9���P��O�1׹��7���\l����7�I��p�I�{�#a"�}������2��]�0Z�����w=�؀Aۛ�`���y3��B��3�u.0U9��c�IF�T�	��F�c$=�����v2�`9���6��ދ��c��L�-d��~S߀=����K������ˏ��p@��ե�~k:ׯwWzD>�}�sy��@��&`�y�i] 3km�7�S2U�k�؊�S�V&�j�v�%��n�N0C�^�'Ad��l��X��પ�!(g��sy�` ��=ɬH�{���=�w�oy�v!�k�t���,����3 ���vU%j�i��ik�����S;�kxޝ�&`6��U[�;�u�kMk�Z�y��������� ��<σ�>��Iμ���r��exg���^�� ��y3���i] �6�� ��}�������w��p ���W >�W@ �o���oy�z��_L�ޞ t�zbXY9�,p*��ۓ��ү@��kO��"�r��$M��K���||�4��=�f,;ّ��W0��h���S�s����Und
�F
�SQ{j�M�K��9	��Dq/a^��u��G�3ߩ�O�;�������UUT�8�kȇg�+��Z��� ;\����T�/v�<�䡆��K�l�π�8 ���v��.�'<�fIj�޽����7u�M���Zs�`q�6�N�tgmq<�F[�	��\^f��sz�aշ[="��9G<�ճ�V�g��mo\b-�F�����\Y��f�N��n0�:�wBF�dR�mjwϏ��n�`Xػ*v�	��@�[�d9�����8��]�5?���~~��iV� 	��  �M� 3�t�	���s~X���x^��X L&�I�q��:H�m���s��f�wK��z�֑�g�� ��-��{��,�.�=�{�|���kx8O8V����|���I$�~�! �'{o����y��*�9�r ��Ub ����uψ��*AK~z�3�����u߻�@����$I$��I	$�?w�7j�v�� q2�[�M���-��j9}�u, p�=�ud��˞�I�[�?ğĎ����@����|�H�vEӍXRwo9'ť� ��V�{��=�m	p���=}���޲�ʫ�v�����| w���rw�����OkzA�r� >@��sY��7��I\���ˏCٹ������SӪ7��b����4�a����h��_d=�&�$�m�������s߾��}���g���7F���<U�k�.������� l�s1��#��?LX1��y�����j��|կ��BT۱���y�ŀ��=�� x�n#��S7{�[��s1`�ɾ�b�D�	GZ��f|�����iw߻Wo�$��հ ��� ��$��O{�M���@�Fǰ�,`������'��:�"	Z��Œ٘���{]�}�=���> ��;4�{߭oK�Y���{ä�r�JӮ�"&8����=c���7(&}c��"$�8�PUKU/�����і�_�<�}����o�ˀ6��t{���֓� �M߻ퟲ!��RC�WdV�6�ܻ� ^�魩ťw�w ����$����L�J�q��{�w�ϯ	\���ˏ���o��x�����>�u��J�� �z2��n䚁be) Ƹ�Rh�S�,&�\n����f	H�	�-Tb�"�.si�k{��/kY���k���@���g� �$�-!����Y������\N	f6 ��+����n������l�]c����H$������Ee�e�C5$����ɲI���B9LgGۿ|�.�%�L� 	7�t�@#;�f,7�,�p�@�!pN��T�;mΧhzM��j��CQO���R�M���j'Ҁ����_��@�����g�����js�G�{�&f�`�o���@}��QC�-��ds����=V�;�R]��s~�H��3M�x��3�����9�Ł���-C�WdV���<d�$�s�	$�7=�|O!]s��� w}�@ g��Ł���ĮT�	mǈ!���[S}�։�٠>��u�� �9�k  9�vߗ}��yhw�w�;�dBfl�|�pq���f����w.f�������=�]��ŚM�{M�W4�h�ʷ�A�w�F ��-4�sV�Ω!UN�P�G���x��n��<��Z=�  ��[oH�9�Ń7�{�0ܘ���n ��&ت���:40����uw��t�ۭ�j�r��ff�~�}��r�j�m�xu률����b�� ||���Op=ނzsJyUq��Y�`�Bj&�X)+O}�{�X|��Mx߹o=�c�|�-z �{����9��2D(mGfE�oc����z"E� �"��>5��4� ���k�_�IϞP��?4�I&ߺL�A�H��s�zt-C�WdV�`<��_џ��N8H���@8I�{��&DDDnuS]L�|#:�G���D���dC����J�mǀ��3X��=t�_�7}��|�����ְ {���$��]�j�g���`7��S�DɕT(	!u!�I@��~�.HB������i{�K!�Qe*���D�������tc�:�2����� }Y@�
4� 1� � !$�Đ� ��� ��p�/���gɠ���8�I�iG�C!����}*$$!_�bo���5>o�y�c�x:rCA������H1��ed>�@�5�(��"���ikdM��
�(ڄ��nҿ�@JuE����%�	���|*��O�!4��>� ��o�������?���Dĕz>��?0_
��G���H��P�O�����]>���������~(I�������&D��_���_p~	��1|��A�`�RI>�P�i~ ���XtK-&����Ȳ�����0~*��k,�~�>��h��~�Ɨ��)La�~��B$�ϙ�SyR��O��CK�?�� ��� �� HH8�[lA�
2
+iJ
�K�?��������X>GA$!_ 4���d_Z�C�K��r-���k��i��B4��?�~1u����F|���2���x��!���@C�?��~�=�
����Q$��	g���A��H��/�#��~�G��ѣ����EB�����S��ߙ���/��Dd�/�|����+�%���p}���jϨ�R�/4pК|�?���x�mmel(i��߭v�!�Ͻ��c�wo�c6�|~�g�?��}��Z�c�� ����f̄������IH@��@}T��m]*�L?��|�v� H�id��VIY���B���]2��8Ҁ0�hKHYB�E$����1SD�����ڤ����BHB�������~���$i!!x���%���I�ԿW�H�SG�?��/��ߠ|�$���1}(?�>�� ����(C���w�h����
�b>����|#a����`��� K�?%��_�}� L`��H�������?�!!�~�������������5��#�H�/�!Q���}H�@m5i&�~���@���z�&-~�܀��فq|0�k�H���_��[����n�b�鏠�X?��BB%_w���?xW����U�l�����a|ë�@_?���5�_ݩ��Ȍ$�g�F�G��C�� ��C@	��&%����
��:�#�'���?��-�����	~��GԆ-�a�����S҉-�A���H?]VM�!�����D���|$/}���ܑN$ߕI�