BZh91AY&SY�G��߀py����߰����aU^<L��  >�@�P�   ��    :��EQ$���(�V�6���TѷpkL��Z�fր������H�  � @���! ��F�� o             ���  �7^�W9����{M{�=9�n)پ����S`�9'�u��ꀠ���K�>n��B^��`�����7}��{���Wy��{�k�{w�s�!���gܹצ���$%۹���ؼ��hg�@ R��)��>�nӧ{zy�q��Y�zj��|�]���\�َ �ݪ�]+q�/

�z���5@���﮴G=�OAM���/����N�h�ö]fθ��yK���n㦌�t%ۻ.B@�G�@l  vO����\W[v�؎ܚ��oS�_}�i�l�c���V��}�{�M۹n�� ���%��Cs��˻�I5˓mۺ���o4kٞ�㻚ӛ�;h���v � N��K�놜�R�n���^�-����L�s���2�a�P y���p⛃ʝ嗷u-����
ۋ�<"����z�hw7M ����  s���^v�Gu�w>�OO8|.z���G]�s]ە��{�k˧G �#�C{ǣ��S�:�<�oE�����N���{l�-]�wnI]��|�                 	H�             ��jz�*(1�@�JTQ�4i�12 M0JmD	*�h� �      ��I2=J!�����M 4 �ѠD��SiS�I�h�Q�zL�)��<������*T~�a10�4ɓ ��o���8I��.���d0���΋ؙ6~��Xg��E /x(��a� UD�@@?Z��_ΕE@���s�_g���������ߋ��{�g�lT���4���l��#���5���r��x�0v�g���ͽ5Tت뚋.�9@Q����;?_��W���ο��:���j��j�'s.��#Tc'Vj�b�\.���O(�Z�9v�
+�J�U�!\+�0�T*D�[�k��UH��}�r�U"Wj��la�M*���2��z'ZVT��j����/���K;����)�C˅���)�h�O7��Ř�`�ħ+U�$��J��Q�8B�ƭ��K�B~/��T!bDF)W�jTG+Q�P��.D1
��8�,�:R�U8��lB����q�Ȟq��8�(�!`��u�[r�<��!X8�+O1Z&\xG1B��\�b���<xS��B1�F��qHRS�
p!8�*)�L���T�i�!�-4!�P��!Q.#X����))�����㕢qǏ�S�W��Ы1��@�X�G��B�\YÍR���h�q���ԩ<�+��p!qN9J'���RS�1%�+D�5��;.-
�p!T&��q��N�Mp!g5J�ϕ�k��[�O��mځ�'�Ф��������s�T�ՍʴU8�T��5��D��U,+nQԶ")�(�s�|Ū�*}�l��!�����-z��U�i%�jx1��S��u�1M1�q��ι��|���LP��-��n�%h\�x���w��1�koV�ڬm<D<X؈z��G=B�"!`�Ճh�Ѓ��FÍB�b<-G�g6�mg�s~�w�,�ֻ�u8Z疜�[�M�M�M�m��$�f�g8`჈Q�q�s�rS�Y�"U��Lq���8��8�q�I. �dF�9����v\FK�%��q0�x[�#����P�O���s9�'���!��Np�e<�q�~)����b.�sЈ�x�mM�$�!s�Cڞ���=Oc�F�L�&2��1򦧍�ܕ���]�RcR�\)��Sx-���jo}ڛ�p�r�O�1�ڵ5���O%JO%Y��+�!3�F'K!E%����(OE�'�����)�!W.�:���+�,�Ji�9�B��Z`��Z}�[��c]"t*B+��]4���bV�	H��b�R�e��6�^)���R�r.�}��ݭL�дm�ѷ��NF�P�F�U��j���H�4���*R��ߘ��L��xO;&��U�_�<菂��!�V�e�#�YFs�q1�0�g7�P-��1�&!p��	�&��xX!h��n�`��=B`�4-Pkg�&#ڄ(b|4���T�z�P���B9b8N��5k��,�����SG�b55��*JOح��K��-F�p�|'�b��!�p�H���&!i�¿��RF]�Te�R���W�G+J�'Ԉ���+�-h�	�N��D�.R(B9Z�,LB��b�{�lLB��#ڹ	����bb�SL\������u�Ҿ�+N�TF܁�
��!h�Z����ڕ&!F	��b�x�G����V��!["b�	��
|+�hB�b�����_	�\��J)��LX��+�Ty]R|㊎����b��S�Mci�ą�jy��z&-ūmm2����֪SP!r���\��Y�Rv�![BB.�P���|���X��\�B�F�-W�|�V��2�MZ��8T�C�Y�X�����f<F�l!�!�-��
��,,R6�E1�Ũ��U�C!�.QNVS�BG1A0�w�b���#�B��Q.QOºF1Z�B5�jhG�ڥ��ܥ��X�R�r��jz�ҫ]��Y}r��m�0B4Q��T�hX�.�-P؅2��Q����D��X������)�#�]\�Z�������v�u���k�o=Y��D;�+����0��iL3_�{7i�ڋB3a����R��d;�E��[���lC��[~ň��!�	�)�!���ԏɤ%-�$#"�Pڴ!�1�R?4!�1
�.a�@�����#.�6,D��j�c��l�*�!��(�I0�F�4S�#�b�hC�b��b8B�C��/�7�B��"��F�!��Z�ZlB56-@��j%�!0��*�T�0�i����|L8B���bIC~��bl8]�7��!m�R�~��Z*�F�1
��ԩ��	��h�j��-�&�~&�b��B�C���RC����"f�hBC�&��v�1�G���r�Z�琜1��1n;B\(��+�(��˭?g�j�[���	��5ڕ҄��ir��z�߹ө�މ�OP�Cuz��\�=��F�3�F!C.���FZ�B16-C�b=�P�>�-�-Wd:O�����NM&x�5��ܯ�gp���j�T�t��wq�w��tԍ�JG�p��b5ҕ��h�![|��Dl1����TC�-�b�b�x�
��HVt;U�V�С�̇�7�_��,���2��|�~-���_����<�8�2�*�\�.a�0Θq�.�!ݦ�S"�##6�ކ.O���-T���QHFT3.�29��qi��f3&�ߙ��۰�y>[.��0�`�V�ka��z�����`Q��tLF�����*[Т�m8��j�*��_���k�g<{N��5��Z��p�{������~S�r!�mL��eL:�#YL��,�¨p؈q,�k3��I���a�;D=����r�:S�g�⋘wsM�r�a�P�J2!���f�Q��cn��&>e�:����z��v*R����T�p��|�����|�:���e<�v�n]7l�
�Ҭ!�!�-�Л��6��|��sz�p�P���w\�GC�w��W���r�j�m�@ۤ��!3V5O?q�(FˊM�
1r�\\k�X���؄[���0�	ո�bs�R��<k�
tq�U�bϕ�Z��1
�p!�Ɵ���8��bK�V��<k�
v\Z�B�p,U#�G�p!I�,�Ʃ\y�\��<xZ�=�!Y..)�)D���C�
Jp!a�!��h�q�c!��;.-
�p!
�,S#�G�p!I��[ÎR���x��s��Q=��ި�؊mj��1	���#�pw8�w�SOG�����RSj�.ǈE�@�n�V1[t�ym�lB�S�[�T�Z�t�ږ&զА��#Zv�8�
G)�����HTk��.��)�!�9_0v9���'m���x#��j��Ş���R�Q{)Gy��.B��`�=��ն",���S�)��aV�[B؄t8��x\6�9�sk<���~{�w���:�i�������n��Gi�{��+5Ìp�\
q%���Q��2���8��[�-�+���q��pzԮF;�q."���pk�\`8�G>�-�e>���Y��z�7M�v�n�[P�U7U�U�HB�����hW�o0�*���>`ָƭ�}=^T�ݺ�wM[1�br�X� �*{�{�~a|+����8O�T���eZO��7g?VIौ�T+��q�i�A˪;��$k���|��H����o�=U��_˗�Q�(M/�y(�QQ7�6�0��ϯ�6fYW$O*o����L>|��ne��Q�IJ��6]]\B���~���M5�<� ��������N"��n����-E�c����5�5N���-�s��XE�X�v��jv�>��י�WSI�۪�K�<5E������&���l���#�����OS�Y��^�Ҝ�z���Յm�ݶB��c�r�uh����y�::�"���wl����b��YU��ղ�1����+��an��L��|@sYE��Y%��U���My��s��-k�z���۳Y-JH���:�QWޞ-e'���|��_z�v�)e�ic�ᨨ���ɾ/��U;0�!y�"�y���q����v�\�e���8��G_/����<�dW��|]���3�Gz�Fw�3����7�o�,�_\ :�eu��ŝ^��s��Wes���t{Է�c��N1��c��T^�L���q�oK�wӋ_��Qa<w�^��Uyu5����T�#�������Jt�o�#$��;�b�ٻ���w[o�F?S�~K���M�b�����^Y���WW�ݗ�Wy����^�㏩rt��9s�x.l�{"��י��9$۷���e(���2r{b����t��҆�jjz`Q�WL��1Ӝڌ�հ�~��U�u�M6M?[���ٷO�a<�Y�*�h�i޽����s��f)���}u�c�?.˚|���p�z�nI&��^��~s�Nw�'��m�~��m��f�'_V��z�v�Q}�=�=��~�{}���5D�~���\�������z�+�Zҷ������q����ϐTE��螭NvjK8� Z��UC����A�x��y|����a��
)�����o�^x=˩��_;}���/{򊮦�Mqo
�s��g�(���%���%��e+��lˋg�ʥ�9yq�G�TIT�y%�WakY��ZoԪ�[�6��S�?�0��Y������rxy�W��������\G�u�1�L˄�.�s��2z��/,��3z���\ˌ��S2R\q��w`�p�l"����]�%	�\K�!9MN����j9��C��.�].#�);��4Uє�utl%� �I���2!�`g5��8��������>W��.���5�d��.}	C�fyg�<�z���2Vn�����3���g^����	f���!��o3�N\Ƌ՜���p�ʢ3���Q圼���ŝY�9F{b����st�'G������x�꫻#F�����S��5Y+��;��He��F�m5	i%Z��4nW!��Wk�����PnSx�6^p�$�^�Ҿ�>J~i�v���>�;j����9u�l&i$�ȹ��W�嬦h��U�5���'�����<8����ɟzj�x��S(��V����jE��Z��h�׉����|�<��5D�*�n;���S�\I��5Kq�k4Gx�ҮS��ӿ"J�]��>N��7;���L�&����+��'�O�ߞM)���e���ia�4���~Gu�;şnU���q�׉eY��s�oc���&��;�5��v��%a���Ǚ}}N�՞݃��/n5�f5i�j���=.�Z��Gΐ�y,�>���rP0�u�L䮋O9d_1�T^o��`����Ś�5f��RIV�B�0S��~����/�s��֥u`ug{�Z�����wX�l���_�D�mE�����Ƣ�v̩,�</;M��l�F�+��W���0m�;g5Y���]�g��c]Y�l�]��*9������o�T�ʽ���$Ք�������İʻG��ϒX�gc�6�mz��!�u+r�å�sțj�����]��[�F�y$y��\�n��G�dCO�jD
&�Ttn(�8�h��'��Q3s���(��#8=��Ԗ��)}�SG�fE(��	��6��?��K�I��^�e�"���<�G��̚�G`��Ŝ��i�y�����Xj��##b�C�=���Jjy�d��m���8�@7�}7�X1����7�Ş��Ė|���Փ;�_��3��\�j%����k�Q�����P;x���,�ĖIQ:�����%�s�,j��s�^D�Vj�Ė*�͘eJ�e��㉨�j9�Y��n&�K�*<��r�;N�s1���Q��,hW�$��,o�"]Qb\Y�.��eG���hr2n2a��{5��ennU�ݎ�k�W���V�nRY�]�u����y�%�"�/�4m��L3��=h�u�[�u�ږ������CQ�uFF�V��³1�J�Cq�����w��5¹`�ܭ�9*J��9+���ejV�>J|�����Hs�7P��۝Xyf��Z���F�+4g�����*J��3�2����=�##��;����m�tigyeY��8���5�Y|N-g��y��N�rlw���y�1�I�qq�����f�5��0`�wI#�r��^n�À�#c.}Tb���x�����5�k�HKhen�r�\�-�Bּ�Q<�ܤY�a�uNz�$w�5���Q3�� �$s ש�/���>D�Σ��q��<:�#�����<��+C��2qa嚰9�����ۑg��=�ܹ�#�E�����%'���/ي�Ȁ��՜Dן1�G4���*�E�@F�,���5���v�f�-e���&G��oYy	QÜ��Ϋ�p�E4��ug��1�j�A%�kջ������s�}��|=@[�������8h��,�y�>q�t��~y�9�N�{�����tӧ'-Yŀ�+9}G�	�7�xNp}��P��Ͼ'sGQ=	�4���m�q���V!\���7FC{�uF	!>xD��y��h�c��`�^�7<�jf�Qk/y̧=�3Ӝ,E�|�8�8H�,h�<>Y�h�V}�o�؏{�L}A�cFUs�݇7q,K8�"ǞXye@o�:�!u�,�vf$h�՜G!�j3���[s�\d��h�x�㼙�C���G��ǕcX���Kt���,ϡv��;��5bj�+�#�g8򬈝y�5`�5�{�b�>�3ʹ�O����3_Xm�\z��������o==tB.�>�����{=;<��Ŀu9��e�_�:�&���}5Gf��w?��]��������5�9'��ߗ�qH~�	�07�{�o�B��W_6��.	C�F�o��\����_�������a+؋��b���y}�t���y��y2��}�{�BIk�W��Ʒ�7[�t���Ν�����T�����!®q�"������:�\]�r�v.��v����g'���7����ި�����#���d�=y\��]�å;���ϵoOB�y�=�f�:�W[����V󷫲��R�jݘ{����A��^�N/v���|��Q���]O{��#��_%]��uJ���u5�$}�^�]��������s�[�|�e-�z��D���إ~�W��j����L�\��o�yf���}Y��Ż�&���{��|�}��E�k��{��GIK���sv&&H�r���y9ԯN���+�)���1��Ɨ]_]_y�`el�VE(z��V�#����i..k���\�k[m������������Z�^��wϷڞ�N�$>r��U�p����{��������c��:\q�u�f��N��O��Ded*~֢*����sZ����մ�v��\�q����K�'���;�:�7j��U���O��ԯ��J�oy���o�����]�����$Nz;��#���H��1#g�p��i���ꨕ��j�bi�C�d$�t���e���5��7e��(T9��(���eZ��V���j,�5A�v�,��8��Ȝ�#�,�,i^�Չf*�Y�J���<U!�m1�7cV$(��me+u��F�A�54J�xd�5��fBʚ1F��Q���HX���
�(�"*��K2,������%�渲�4���G�w��&��K��cCXE�U�N�QZ0i�	����b
&�bU�5,&7m�`�:��d)"@�Af4�$�dQU�`�%q4�Q�J�9jX,�,x�5��ʆ�Ƈ\�V���iH8���5f�"��Ć���wid�FI^Va	5(��7P�h� ��D$4B؉m*2aFeUU5�E���I����_�TlEXM|K��^ٖ�h��՛H����V�kʎ$���H�%D�fKY�Hbi-ܰ�1�PCE�Z5
�����D�U��7ۢ�����F$$�՗��D��8$�I7�PXۈ��DQJ⊈*.��V�(���ى�QG�'.���
7�A�9X�"Q<�*�D�="$ưԖ*�0��ѥ�YQA�V9fc�8�VE+j �,t�Fjr�
�$�B0�;�%q#�!unꙬ�sdrR��Y�1VK��r�`��u�I#Goյ�A�0J�+p�d���VHl�B9+�$&F����	E�� �k2�au�y�ӭ,���I�MD`��/ј%���f*��hgQ�.<��7�*���V��v�河3��A�������
�o��
�r	��AzJ���Y�E!7�u5�^)!����i����.d�o"�T�'�'�v!!�PG��R�H�s@]Va�&bfR��%�ǰ��D��$%�n+�:�7�/4b(ȸ�����MxxG���1����"�;�Ew����0L�91*�Vbjə؏;B7.�	�\C�f(j'wD���P$Z�(T{7r����Q��U�֪��!������Y�e5�OB{��`#���ޟ�{?������}����W�(��}Q�U�Y�I���P�y5��=_��_��7�T �H�@� 0	  Ѐ �
  �   �     ��)  h@ X  h�  � �P X  X& �  Ѐ�  �4          � !�d��X�m2�c�9�.3(ʶ������95h�Vab��i�q�Y�lH�r)��nM���H     p�  @  )  X  X� H ` �  h0  � �@   � �   @    B  �	  �   @� 4 A� p���^���~M���(<qͥ��%`�(٤³(��$jfS2��m�bY���y�5��@8�`  �� p �  � �I�H` @` @  �  8`  0 �   �  @  @@   � Q� @� X X �P����o�I�52��[7�ۋb�[��j7H8���X嶢���ƽ暄��57��}�� X�  X@�H `0     က  Ѐ 0	  �	  � �H X H�  � � ` �  �a;2     p� 4  A/	��&՚��#i6��m�#��M�qJ��j��6�em�j��R���r3r�FA��PR�M�GpARᚆ�j¶՛�Wx��x��ې�Jg=p�TՙՊ�d��;�C��C�����PY[G�����_��������o������'�?�M���:�2��6��Dz+jB"0���:��#��h󍲆�BB��єeL�2��6��8�����QGQ�uDDy���G�L"4�"#���ʑ�m�F�Dq�emiu��iDDy0�DaDG�%Ty���F�i�2�)>�_B�^B���")Di�R2�:뮺�#�\R�Dm�G�G[F�0�R�!DQJ��<�0������G{*3ެ��be� �R�FZ�p���y27cq"Z�m�i�	��K-�����*u�%���RY�B���T�U]�_�hz�X��\RD% �����nbM���x��ƘH�ʄ6���bJ�����g�
�Q'6����Y�8�1Ʉ)
R j�����QQ�`��b���T�h��#P�%�$,D�mm"�1"�B��e��B<��! N�V�5����4�(�ML�F���R�/��+J'�Y�T˖�5A+�c[���eC,-��cv�t���u�J6������
�+,hX�K*���v�E#����Ia2���+���b[��KF�j&%QG�eL��Y�d�������"�#��4SG]S�͍�Bdc ��i �"�$h�4�^[Q�N����uk�Uc#�$m�X'[���#��B�����4VB"1�$"�*�%SŒA˔q(�;	c!Q&$�����K�B�#*�\���H�7(��)h���c&D*�i�SLơ�5jݘ��������$Q\b��F"�6柣�X���S�G	q��4��Rh�4
�A�E�2[-�s(�ȝk!1b��T,$�(�ai^1(��2���AlE����q��FX_�WT���v)h��b��	'q�r���nA��\R�dx�-�s)
\���H�X�3UB�,�RѰEʆ�0��J!di*J@b	G�c
���	";V)�DȊA�)��!QHIb,$"eD�$,��(&YI��� �h@������T�"E^D4C�))��\��r�m��B�)I�dlt��&�h�	H��$&4!1�(88ZDFJ"e�!�l����6���B2�Ҧ&<��PhO@��1��		X�np�]X�~&�j�ib�"ZGp��F7���d�A�	V�Y���GI��r���Q�Z�H�E��"����JJ��K��ktX�H����TQ�61���b�I����:�+�ح)Gn[$�VYZ���,�J�$�������yGP��S *�*EA���*L�&�Y���H��-�zo�pe�QC�,��R0����ŸǏqecD��7��*C��q��k
(4<AE�x�A	b	
����T��<������P�Yq�RBbg�4V&�+�2��[b�&eb��q�e,c+�2ADH���T���M��W[ň�����IK�,&Px��Q"�H<�R��*!2�$�kiR��L)Y
�(<e��v�5dĈj$hU�&<�RԒ,!)n,����C%Y
	Z�p����FF��B��CD�rQ�$>л���-) �T��ϊ�n�1��d�JQB+���¢<Cq*�H��T!4�H�(�LB�X�!hB�QY�GfQ��E�'����e �dLv2�bL����[�p�*
bj!���BA��Q��eI$,DH�i�d��
�S^\EO4�.J\�H���K,!Ue��L�ʉju�HG*���1����)dl��Ә��I��mMJ�VTB�%�uZ�IUH$�RGk������d��b�i;$N;�X�eq��)l�6G%�<��$h��7$����H�v�UF����Y'n����K���'R��Q�����d���J��9�����7^(6�T�mQ!5Tc�q'Y+�V	�RU �TJ��b�c�7QF�m)vJ�vJ����Ciښj��+`�B��E"��TF�j�<rH-�-���m�*V���`�3TN*������r����k�B�
�n��n!���c*�`�c��mQ��I�4��U� ӕ&�PV8�PT���P�GV5n8z�(����!)Ru��Y��ȫV�]�h�%��h�+�eN	�'!'Ryn��O#�����T�)m��&�q���lR�܅�����j�	F78����#ep�ΡM܌i
�ˉ7�
��+�����X62���i47v�eI��%u)e�%DV7��<v�Фr)+Tbp�mA¦�R�T�RK+��i8�J��kX��r���"I�1["&an["���\ER]�c�
�B��Ĕ�47eeQ�$��ep�v�Ԣ��Ĥ�m�����c�I�R����V�B�K[Y�crB�Tg�٩�B�ԔR)��]#�5	)Tu�C�9H�oUcpX���U&�'�X�F�����r�Ȗ�Ze]���ę�W$j�E,pD�Q��0v�m��4��:�N�76U�m�$��ƛ�7���.7(�R�H��y��z8k*���H땥�1��\r��20m�F����|}�  � UUQ��������  �UT|���^ �   UUG�^^^@� ��I$�$�Zֵ/��g�-jZ�[+ikG�i�a�y�:��w7��}�(�I�)T�hYd����#��DRb�Q�XJ+YD�Q�<��E$*5T��[��Gkō�2!U��5X�¹�DC��UZT7�4�I�Y(Ճ�)P�[��)���&��JF՘�Lt� �J(�C �팈���0��"�tCD��D�"��Q
7K	+P��JR�D!
�АL�����-�x�2�HD��p(4�F�Z(�S(���:1!G�AGb��(�)SAdCb�ŊB�R�JHB�,@�B�	 �1���2�!d�By28'B�)0J4��F���u�Ģp�	��%,B��F��P��UaX�$pBrK�I"�����)p�H[n*X�v�K%V���퐭(Ǌ*�X㵹'��X'�؋aU�c���R��	)�U+-T������ԑ*�D���(�*t�c�M*Ԏ9[ۻ^±)m�(mI$�`��v���~�{�wN����{�xds��f���j��s;�h�.�N��|r��'t�G�:�����b��q�����mu�c��͇r����l���9۷]
��gK�y��z�@����'�ޟ�7'��i�?F�Kh�O�Cn�No,36Gx8��?�B���d.��@�<�q����]4`p�rӢ��K!��C�<8}r_��:4h��� �%��@��J�E��6��O:��������!����!�4�t��S��"#���è��u�U����uTI6��ie���l��$�4�3��K�����j����PW+?{�m�=���X仢{�>�1�3��p��ҏ�l|x�8du&F�vpa�R�H�^!����o��pp\�|������*R9q�u�Bh�θ)ŧ���Y��:lɝ`�%��Ԙ�D��|7�:5�~t�*y�]e[�qF�FG�S�2�b��b�X��t� �`$�C�
�)�qTI�ի
��CA��hM��F�F�8bΜ:�
<(8g(�G:(z���^��$.BH��^�9���m![��8w��9���=5��\���vk������4^W.Ňpp/>��)���J4U0�Zv�񑳃C��j��ю��8{�|�T��u�Z[�qF��P�rkV)Y���0�9A���:�g��Hj�rJ��ݒ�:+��&������?>4�||w�u<��\0fb��/��!c!��M�YX4��pp<l�A��*����"[�I$Ιr�p�s�!N�6�=y	$���K����ww!��N��OO�c�wW
�)�8C�e��U2�Y ��jEO�Ho$���N_l�q�jFCE��Q!���2��e�\iב�Dym�<�p�qR+��+wFj��X�7���9v�%�	�8WQ�u��6��WQSN*ƥY"�%lbd�D��m��7	T��+��"���u��7˷u�B��*�3r��i���@թ����K!<T����W���ˎ����P����s5�M[�V��9=:Vڦg)�&�&n����ys��{'�5Xlw	'ȝbb��H)��DtA����fƍ6=xy-0P����d��p��9�+ʲ�ً���nΖW��a#h�m�\a3����F�mB��4@���K�5�F#ߊ6{��.�vD�K4�M�T�Ya
Y�8JIp}���ޗF�|v��I&��h+�uM�ˌ�ӯ#���<�<t�,�>������I�jR����$�H�㦔�1f~s2[�Ui8�׃Ǆ4��/7mW*���񙉒98M�v_��IC��	ō�pP�}C��IM�|9:8[b8H�M�X�8�Đ$�~�X�C^}��69zh�O�i���B����F��,t�4���֫��d8m��[O<�"#��8uyN��o��+J
��̈���I$��������4�#K�:�n�ܬ�*BBV���LzL-�b��o�=���z�֨��s�|7(��7�h��񱬸"@��'}K�X��g�_�}�}�<�N���YPEQ��\%_�ºV�x�D|p������RWR���x[0��cnMcr����7Y�9��ߝ k�rHD���0Cf�<YƑh�"<�#�Q�댵�z�}MԨ��i��c��$�Gs����e��#���xgfCgZ�T$`�fNj�:1�\:����^��wqAi-Q���=��.t;RE_.獥����!LlI�"Q�4F�zCc���F�M]Q�F>K�����+��7m���`�pan��b �|x�a�C�&ǥ���I �t�dl8:[,t0x5����s�h�G[.����<|p:|x���!�|�*��W�^q5f(U���G2�{P���H��&��C�ȥ%�B����I$��k�Ί�yY�s��6&���t����;v��l����<���p���
�)L�ն�v�-OB���q��Q*\)����Ӝ!��=~��_3�_�_��7�篾��Hq��٪�����p\��~T�ӝ���T��*��ϪJ�8pc�ȝu���֣pr@���:IF�0��%(��h��)س�S8x@q	t��N�M��M� ��n�XV�%{M���1���6I��I]<ð���:�$,�j�Z$ӭ�OfN.�86��n���X�m�U�܉>�FBU؍�[)0T:�Ci/#�BC�K2˭:�8��#���y�:�)����q������I$�f�c�Y�=Ku���+c��Y��Q��.�$����3�d�뀧��H*��f-�:ѧ�<u���;<��a$*�Ѽ2z%���;;��:��f�`���$_}��#9�s���^S�	tߍ��dl�P�ÏC��H'��h �c'�á�jk����L���#l"��Եq[uy�ڑYU��m�e���k�ulڭQlq�U�Kb�jʭx�c�b����d����Y6|?�	�|i��ʕ�����S��U�⟕N�j�-���)�mO�����~'�~�+���Z�[yV�Rх�W�XZ���*х�j�aj�b+αm��[�Zئ��Z���U��n��-Ka�S+1jҖ�����S�ū�WV�֮U[U���ڵUliL)�Z�Z�V"ص[�Z�V��q��ŕj����j����O��O�N3��>8�2k�'��/DuUl4����U�꺬}J�UU��Z�KR��b��U}l1�Z���mb�*�}m0��0�<���������W��X�[�-V��U�űj򮪭QV�F�*��8����[��x]��*ysv�읩wZ{���FRZ����韾�b@�����!�b}��=wT�;���f�b��/���"��gֽ��I�_�n��.e]��sG�k����I�WO7�yɝB��귚{|C�Uݝ��]�"�l�i`�2F�������gf���}��T���i�
�`��q	E�}+��yos��͙-]zۭR��y���ۧ��,�hPI��}�\�y��y���Dm���|�����W�%~��Yh��sk�d�������^z�x>���� fd���仟wvw}���� 8@3'��������������}� 	���y{�����������}�� &s�����yO<�̼��[���<�y���ΰ�,�)Lc5�g.b***	���c�S ��([<t�E�EŇ����q�l�� B	�"�4�i�Q��)J�{�]7��Rz�dL�Q<�l�\8Cl���x�Ѓ�1�R�&�8�Q�骢{4�&�>�|S�I��[XÊ٧#����I���`P���0t6�l;��!�B�Н��	���8`"��;Y�0r [��'4I"a���G�b�������lԍ\zi�(�t���L� G�a�t`����	�R w��� ��g�FZS��̼�ߟ�y�^u�g��Ǐ�g���**-JN48av�!���a�$�#3Dd�g��<F*S���3�Ғ�3��H��-�W*HX��QOЪ��0�#�p�4�6���{Y ��%��EL6!Ǵ��ѱ�@p���L1);eW=� Q���B	��a�&�?���gYI%����G���7����]uF��̣⃜,r�;i����qD���BU�^N�\)���d0���ְ9 e"���4o�%�D^��3���i��)��x�7�Ӈ����1�}���|ᦔ��/̼�-��DyG]"��.���Ӹ���6K&��+��$�2-��,h�Ֆ�1e�!���Mn�di��h�p|�{��MG\�YX뉌��1��QQPH��C\[$Ʀ�7���1��n��jes�P��m�Œ�t�V���9!U�g!j�cz�w���Q�T5���>��6�;`~ܻ���e�۫�w��@{�B�D5��E�"�U.���9"�5��z�\��mw�n���x�{��D1����IF�HM� �lK ����(`d��%&p4� 40��7M@�$���Z�k�a�!Q6C�hJ"'}$��<?Q����'��UuE��ò� sn%����!�4@�T�4Cے���9�X�F$StF�_JD�}���Z���|A% 5���|<��y����ϙ5�g�'�`;a�	Do��e��b�Wy��U]�Wv��	���"� �
�[}�R��V>p�=&�L��P�,����o�[���L���u�柖��"<�>:t><~>�r��v(H��	u���"����9P�� �P���?C��D� �1���&��D:@�\h}�QA�䍸S<g C3�`w�Y��80xp�U(��C>�4Dy$�N�5��$a����  �`<�%J�<����l 9 $q���- � �P��;�|��,�����l�X��^p�!���? �#1��ΜGzyM�<�ͼ#�Aԧi�޴ܞ���7Oh��)�D��Pǈ� �:0���a��zs�X���>�od���8}������FUTл ;Q��>��]e�Ê2��4ʝ[+e����Du�<��y�Ts�h��,H��̫?���gN������Պ�p�ْX ST��'�Ĝ����$BM�@� 勈_�IG��4�ɂ���@t���Y��m��)A\�TX�A4���;�P�)�	L�v�S�P�˓i�G�-���g��O$yi	�<𸋈 �9���P�D��)��t�#��Q��6�#��0�q�策F1��f�֊_���2}��L�L
l�,��aB�a��PP�\���<���i�<��G���t��c����Y�;5Kuv$�e�D�Q���܉~+��:A!D�u/��f�gA�D@S
�H'2%�h��Ռ�^������~e�_��o��8��":<���S1�KSLF
��.���@���,��QQPH'�P�	k����6I���'z[��(�ǅ�&C%�H� d!�����n��c�̌=��b� �d�r[�s�:A�%V�܅r�kp��>"�����#E��}��O��,���c#0��'�7�8i�Cv����%PYk.7��H0�W���m+ p��6h��HX��
���:SD��Z���9��h�/&��"�IJ&#{��3)� �f�?t(��0�4b!�$�l�l�� �H� ��7h@������A�����UF���C{���Z0�>(���N�6E����J�Ud��ӌ��ѷ���Du�<��y�_^��V�ě�}�j�n�9��r�h���#�iû�Դ�>�7����d]<�!���
HQȗZR;'q���6��'Lk�7i����vY��5g�t����۾\�v�C�a�g}��Z��fq��ы�k���̨�y+��]�������潿uTF��I��>6�R�f��n>#��Mw|�u��V�[Y���&�.��$��c���H A��qt@40~o{�Xv�����,j�&�%�hz�`�ޕ�M=���:E�<ZL�C$-�����u!"`�T\@L.��d1`ўx�f��%�Z�.��W�-�aD>�	$&,|04�\�̈q����2��L��<�F����Od����4�ADnF!C�%��|<�45�:�bC4�DH��aрX��Yd=�FJ40rg�������1S!8����o�K�ݦ�#^��n��3s�}q�FA-13��XB���Z, ��(����Mϔ��M4���̭m�?8��"#���yl<�&�)���kJ�r#��k!�"����	W��ܯ�64�JBhh~rダ��
%]�����M�L�'\� x>��q
?&��Ȑ�$:}�w��7���*�h����� ��$��|���v�xn�ߍ�|#�3��H��2A�#��bOh8<_��- ���f��݆68�F��O����,znV19"\/ꑒ���OF4P��#2��8w��,\?��!ܗ���N�5l84 cd|9��c�8���$2w��\�%u��
�4�j���]S�el�?6���Du��<~�6�v/ꘚ�hƤ�HBU2J�4��TTT������9FL���	����ɓ;�=���:UUZ���8<��;��f���8���[���}�EU^�^8�FG��Cp��7x�~:é��&���Ӭ"
 ��� �����6T7H�:h�4UX�xy����AM�B�� n��|=2��_B`p� �a���d�t��o�
(��v³v9���㿨�r6�Zt���4 wÂ�A����_���]�e����'>��L���2�|FlɣBl�a�e�abG4S挸���]Fߟ�DG�ӧ�<x�3�I���ڷ\�a�Ix��-��ޢ������_��UL5��À���G�8@��llr���\���a��i)t@�ߔ�$$q�|f����q�M�3]e(uA�lÃy28h}��e�� ^�(5C�ی9kܪ�G]�PYPK#��0�!�t�tM�rѲ�@ǡ�ۼ�n��~�U����ǚ���~<pphm��D�z��eYr���rM=r;2��8��`��!�O�ϫ-04@����L��	�`9aC��4ۂ-`f��0Fm<I����	��A�d�ׄ�a�rBM�\+m���4#[S*~W�SH��~a��SJ��mY������}lZ�V��b�j�o5�-T�-V��Vũűj��U�*�h��aű�ڲ��)X)UR���z��[�.ԝ�÷7K��.{'���O�}�M��M?0��?+���:�RԊyl-Z0����Z0��-_�o�~U�1jy�4��+�Vehի0�Z�V��u�*Ե0�S+b�u�V-]U����6��N-��\��5Ul6��j��jژW�b��զVͪ�j�ص�n0²��-Y[�q�-�TU�uV�ч[<U��M����Vb��p��_4�"B|N��!>$���o.Iʝ�9��;N�oeKW֭+�`��ylr��DLד5�-]T[���[�ey�b�űj��U�j�an����VT�K�w��T���z��v�ړȳD ���oy��w�����m�4��m\�no��6��g}�ʗ\!�2�F����oE�lH�+,����qs]q\�����	yî)�����:U�^Ϋ_�zרP��ÙW;�z��lÇ�N�i'��č"u��Эq��z�=�����]p�}!>�
%��5<�Yw.����%�ٗf�~�n�8�ۧ6��u�����K4�2����9`p����ݶ�����<�xǣ��s%޴6d::�����잼��x�/�[E�Fɨ��vDF�D�\Ìz!�q�刻{����de}��qL���K?�	o{o���>��9оsگKw��R�tqs'Z/���\O�����Ǜ>�x7qF��@���9�y9��O���j�D��JR�өȒB�j;#�N�u��&I(�+�M�XQy:��5�b$�c���bU[TC�[ Ԏ��$��Q²Z�*�E
�WT�N1�KT��Ј��V�k�A&Y����kշc�����I:�o�w�}����{�����{ww�>������ �������32|������ ����}����ywwOww�` ~���s�߾|���̼��6����"#���yN��8�;X±�Q��W
Ь���)������ibb!�T,�-�B��+�V�����uB�W#�X�"�S�6�V$�2�QV�Y$j�#�)d�B!"$��m5.��)`�^\FR�e��Be,��ϊeRnHQ�� ���C+
�$���F,$�$ɖ��KU�N42U�b5£M�Q,Ō�*�K��9
���%�&K)*+��P���ZUe.6�&�"�+!)h�a!J4�ɈbeTrƬ�&�M���qэ���D+D�MLQ��(��A�K�)JA[�<�+P�9�R&*�j�ԍ�[%�"V$����ih�IA�Z�U��+���1��$�rQ2�S+�-�&�j�Z�VJA)bQ���9`��H��#j©H<�5Z�c,��,n��ef��%�c
���R�Li��r�jv����bNd�-�&��1�EQ�c�e�/"&X�v1�c	��t�t������ӻ_�U�P�J���w����{��HN��^cG��;�L8�S{k50��-OT#ʔGF���f���Z�]�>�"�|Q��f�qKI�R�Þ�U}~���Y���m��˟���~9�z�%g+OͰ���J�C�-�_:�U�|iӢ� @��%1��{p&GA��	d���>c���n�&7Hl������9>��"���[Q����E>��@���P�rG/����+��*���0B�Kӫp�[d��=���������{#�%\"o5��g���a�,�N�,*��.A�|ۇ���;:��QX���0�	�3� ��}{�"�c�ɡ�1&�_�
�B�hϽkjY�m�:�_k�4��(�>N$!!4I5����eaZ� א�c�[��2�ͣ��":�)��:~:#�ߕ-�M�!�MCL����1�`$�!+*%��6��t:s�5�2@�&�'|.�ty����0@������nM��so3s��m�ӀC��M�~�����"`,r�|@��k>���8p�L>��޲�F2�O���.�_	$��B�.���#�:J��r;��D�q�kw����ԣ�2E"E�ea(�R��=�{ȩn����޽��ܒ�Bg2I���$cͽ�E��� P�v%��'A�Hpd �k�hzܴc[P4Dv;�(<�Q)�b�-�����=��,�S�2�/����Dyu��un���Z�+l�S�vl��,@ΏMf�,�gPE��ٛ�;���c�H׵O�/0L�[W3�3L��b��d�@��,�� 4|c���q.��Bތt�;��(1�6^��M�F!�F�"H?�b��W��X|% i?M���B�Ȕ^Z7!��#?�H��q���:ݯd�ևoX���\>������=��4�aCԮ�� H�gِ$�p���䧍�4�Hf�e��hx]!g��;"��l���'M�������@;�HHa��j�YIMX���7
�� $�I�^t���Oё�X6�0:4���&���[��2���?8�G��QGN�������.��]�c�1�����2�(W?*��UW���P�T$>hl��0�( ����~��)��([,y����3�1�(Ƣ�5��vID��3&�6�,�(�ތ���� �"d!��%H15�Q>0e�G�5�ǜ�Xq!:n��٭�OI��74xL�B���Ph�X&��	�vw�4�:@���`MS*��˃���Ir�1#���ሷq��Ɗ����4Q&��Z.*�E�T�">��9���$sMï
J�p�[��a��Zx7F��mC*N9��4�L?#/2��ߖ��DG]E<�Y����|������U��
�v�Nw��{j���
�SiIXΊ�겙���!x�NIc�����^X�6��}��c�0����ߏ�SY[�Y��J[ڋ�]�o`ܸȒ�WۉƾV�Q�R��%Z���Rŋf;iH�f�\�
!nf�WX�ϸ�\B����R��R��s�y�SǱ�i��z����4�S�䬈-غ̇�lI��5�O��?.�C���H�Y���>3��b#������K�D�A�b>(��4�c�r" gfC�ʈ,g����q���D��Rv4��>j��I8<�A
���バ):����7[!w��cR����x�2ӆr������e�Ns��UH$`'��� Ѳ�����FBG�,��zi�Ӡ$�v0�ka��
�0��H2�Ig�Y��Ѣ� ��h��t���a��hS,�;���b�8A����M�<�̯�����d2A(���$���\����U�������n�2�,<�H�ѷ����":��:C��oz�W�r��;�����F1�c ���}O+aʰI���0)��C�3L��)������J��� h�~�|?$ѻѢ��^rgS٣��q���{VXt ���R��4t�8ui���(  q��9* e	�{]M�u�'H@���E1�_��@ �(�e�=�,�-%G��ut����$+���Ӊ�r��B�>��h��M�24C�
>)�� ��"|I�bW��m櫬<ْ�d�(rC�~�{��Y��lyA��Q���Ъ���ɡӤ����x�,��.��O����e�q�e�m��Ţ<���<C�Hp�&���Se��-���^�.1�c	 ���d��r�-n_��ٱ�����Rx���z�Q&�; �
cL5�#iC�a�h4E:b��5���r�C�.�b�b>�0���=X5�a�}0�G�
�ɞ>�h�f���r�9U������,,���T}K�^����7ѡz��pl����`�ȵ��	�I��I��Å��0%�$0t�qFc |B0���K �Ӳ1�&�]ݚx� d�YiT\.>?��ء$q�4����R�2��ٲ�9���L����p=��$jI�W�s��<�H|yL�:��/-����yu��?�����ۉ*ՙ�RA���sw7�1��Y�h�XB�A�>��.h3!��eC(��6%d��}�;�P˄�H;�h{`����oK��S����	�!��8~li���lh"�/��CdwZra��D)Z!������(�~�E�f}Z���� ��7��4�$���D-�K����	�¸T��h�'����<��WGfD���EǛjF�!���� Y�t��u��2ꤠ�u�>�cO��x��(p�E��9'�ZTk#A/)��Z~ioͿ?8��Ȉ�G��������{�����f"�.*�!¶\ZQ!��!
F;�ey�ظ�ˮ�G�E^ꈖ�ՎE��e��4MjNjz1�c	�-ρ�3+��),d�\���J�oy��+i���q&�rt�]��+/�q_U<�'��j�y�+P��"X�c�����_T&cx��l�U��T�%Od��<6X@���p�~o{�Fhx�ǅ�>�%u��"j��.�[wn�5p`|0(�e�H8:��F�G!�n��0��@��TX��vV�U��;MT!��t�$6��l ���s%d)�Po�?D�R�~Qbi��'U>�!	0c������0/)�;�R�H0a�,���iP�V�A�)<;(�44D�:{��亽5���KQ�왖L���9H�	�iЀ|�Oۡ�� �ct�!�ŝ��_Յn�	S��}�8��u�y�����y<C�Hp�\j!�ō��K�reN� �3q��"��ĵ4�M4�$	PJi���Yd+�TŢ`�g����2~8Y!�P���ޯ�r]��Yd-2�85��F�v0��������կ�F�_�e���ɕ�M5�)��0��nJha?(5��l� �4l|X����F=h2��R	fƀ�l��cH� �����VK!%��_��KM9­��wx�Ӥ�gHH¨����󡡲V�װ<��CA��Y ���楗vXQ�7�xI&@���8��#D$h |}��v����R��ަ�T*�q���>��h�H�!� |C
px�'�m��ե~W�y�ձKcJ�qV�ձj���Z��V�8U��ů��j�qlZ�1UuUj�a}V[W�VWz��n';�[�Wu�i.Ԗ��L*���J[L}���}�Z��Z��~W�yO�E~R?0�~TWߑ���F-Q^U�a�E��b���]SKb�j����ͪ�S�R�j�O+�U�
Z���V�j�yKF-Z��lJ���-\�����bl���>ƙ�O̟�L4�-V�U��mQV�U��kbե�j�f�j��]U��0�U���ラ0k��c#d��O���G;�%ڪ��ĻRv�����U-XV�֦Uj�,Z�Z��u��F�|;��ntzN����'��I�)lZ��+f�űj��^*��V���XqlqM+*����W�U�U)j�,����F-T��ʟ��e_UVL��;ߖ%H%�,�IA�&(�#˻���U92�T���t���y�f�!�|�vX�������W�sㅏ�j�t��#w�=��系M��.#��Y�w�����Y�$���	��~V�z�v�)�r��;������^wϞ���i1]���mإ��Ia�xRo=�s�6r�C�-w�N��ܖW���kw� u	N��ݷ��� �y�w�Cx��śx�T��I���;������@ |���f~���=��}�@ ���g�����ﾰ	 }uS�������}` NIRK޵���<y�<��<��6����Ȉ먧�S�}��X�s��j�r�˗#���QiW�Ӵ�7R⁯;.��4� �a��qJ�E}�j�����O����|�t��S�Uu��8��
�F�DLن;�`�v4(���⇆��sRX��{�4�"QK��$ ��Ĺ�|3�A��|[LZ6�*�l�5�B���ծ��4�q�A�w5=v�I	�UV�8!�9w��S����0R�����D�cсCФ���p4��E bP!�G�|_ɥ�W�#�ݲ��6���!��1
S�9��,�)�07����#L����:��iƞ~mo�-h��ǎ<C�Hr���n�2r�F��,Ϸ.1�b�$��gBh�,��&�?_���~�0������������<��v}g�!8v�O�&q.�(Ԫ��x9:q>����T2&���{�%J��QP������\�oD����I<o
�r���m	u(��#�Z|cxm�����*C7���!�����Re0`!��đ�2hpP�2<b����&N�J�d��c�60˺Rș5����Vl�d0Ƈ��d=�!Ұ��ޒ���(v`�t4p��6�~�p�ћ�S�6��y�����yu��˰��D���E���q������]Օ{�8n3Єc5L'_i_7��ɏh�t���\�7"�Ưqh�Sy�,}��K(��Q5����&��������>�"���$��;�-Y��z���}�&Á!�X��Gg!�8#�iQ��򦞬M\��9z��n��Kmd���9ZY+5=Q�;j�U�Z
VfߟL�|�]c���	*T���&���DNض����k%�On�n�˹®��o�?I�:�i��I��I��x�#I��;iƝ���Ř����]ɱʚ����Œ���E�0xS�q2k h�3�2 �?fS�v�7����v֍��eU��lhp93�:<�����:�p��E_�K!�;<t����!��æI ��Y],y�7��0C��C��&[�CF�(����1L�YP��Z�1�[��Cez��XRagY
��T�UUC�i�صE4��o�I�/�e�?#.��-���V���x���:t�=kt�T�)wuN��z���А�ԯڬ*��H�L�ó�� ܁����0�<Ys ��#ڏ&q)��i�xL��K	���f6�$r;H!�Ñ��`r�tQK�hpv`pY��W~4:�����Q�O���>q(gO�2�˝|6=1AD5�N�H7K.�乛�>�-���{�x���:��x�hy��Y��i&
'�f�;�|sƃ� k&��fN7f��ʃXC�x0��Õ�q���q�8�+eż�ߝZ���u��u��n��cʒfY��󈨨�	]z}-��*�l��E��ϴ<t���t25��u�����!
# ్��x"B��&OY�&���9�o��2�t;~th2��)���<�Y��@�|p� �#HJ�?߹4"�m/̎oz�lZ�P�T��H~����	�i`h<9a����!Bn`��E�x�����0�7HC�5b0��R��S�Y�t��)Q������v�V��C��33f��w�-�z�6q�z:r[����ܑ��jOy��53����>x8("��*y��e�^qoέkyh��<C�Hp�lPeIU87,R�sh���	ғ�7�+����J�F �ј�HH��(�0c��Ya�>���:�Zd̑O��ʘ�tK�������x���!�ߜA�2t�-��q�����C�e��5E~ ��Y���3�#>2���@�}���^�=��l-�Œ�+[vv.v�g�Ǉ��pۆރ�A�/#C���M�,
!@p!�o�t�:7�3�4�f\Hnƍ�(�(�$&M��ݰ�O��2�l6�.����ߝZ��������<#��6/V.n��k�i�֕"�t�=X(�^ծm��uR)"q&�J6D%�񍱸Q�	�th>����u�V�7>-p���C�Uۍ3HU�.�y�o�H.�Nl��1����g<Q�|��^�W�
�#��='v��mo��b��WZ��͍��C����7��.eGFTDB(��e���Ãư�Kr��4A�"�޿^L�#�9��f�7� -�6G�[�s���v�h�]Gs%�)P��v��4@�d���$aCF�3���פ��		�v0!��y��=#2eð��>�;TJ���x�~��arCHQC��*2I>��)C/N�
ԡ!͒C�$�����!�F����+��G��ϼf��#�16�O9�����m�U�Th�0��/̭ǜG�V���u��u�>�9�j��n����Y�p�:Fj#��ГF�3[�y� �P?aVa_ڱ�$Ն�t9M}&Kz�;�CG;m��1�Q�l2C�3"O������@�0���#�	d
2��Lcm����Rz����v15�m�>���\48`�i��� ��/q��H�<�sKD;_O�a�����؟7Wwy��e�5��J�Õ�����x�hu�a�b��cY �9!�E&k�`��Fy�Qۭ=�A�(sR|!�#�����N���ɳ/2È��/8���ִZ#���yN���ǫyf���Z��E5��i�!�!R�6��M$xQ߾*�䙟}�2�:m��>-K���8v0�C�Fɑ�h�u�>6q�QrI{�L�G�<=�����;ʇ�0`Q6!�P���j��1R
d��V.�6h���80|P`�������c��_��p������~:C�hу�!��|3��G�Δdj�Ψ�Q͏��n�}kW)a�
��GZ�H1O����CK��$��r�iX�����ItΛ��pB1���n^:���,24YG:e���~�kE�:��T�;3����ƒEl����2�+�DE�X��jFH\�5�����А�K��6M��(�܉2�f��B�GR�o�<A�!TBWi��	c$�An0����~4?>c�i�!�����4�O��O��)5#O���}�<���)^yo�ʝ`�*�o���o�Ѱ�g���,�*˩v]:x����I	I�~��G��1���2<x�㓁��磱�Bz����c��J�d����9�����︊�ʈ���i�>ڢ�[�Oتi�-QX[U�y�[6�U�ů�4�)KU��պ͸ŪշW��T[U�U���U�U[Sjʝ��vN�t��U�iڗj[�-K��Ui��m��j��ڭ_[�4�>�uV�����EE-yl}hŪ+��E����n��b�bя+�Ҭ�U�՛V-�-�-V�ٵE:�*�j��̱��>���ڿ+����[l�0�>�9Ul4�U�jҭ��U�[fե�m1jZ��صZ��-��V-V��V-Qlu�-WU�"شc�U[[�4X�|%�����p��g�5��U|����q>T�.�sr�jR�ʭ_iV�6ū�S*�uKa��|;���:M��������	�ձm�jZ��W��T[^*�N�U[SJʬ������������y���j�2��R�W�V��{�����?Ӟ}�]������"Q;-t�cy��?*� �w#�LnVS�Ӎf�վR��:vtʎ���4ڽv�����|������ާ��Nm�7G9����T�9�1����!�*٣�?tSN��4\Wt��`Ą��T��'�;=�_�:�xJj�]��N��K�i��6=ȧO��2id|���9�K�'5w�N<[0��&�_w�����[��ڎ�{�t_+N�M|9)�Q�C�8Bm	ǺB�x]7��O.g{(���9�1���&+j�{�ev�����B}��]{J���5Q<r�>��������Ӽ��U��b|^���Љ�mu�u�FՖD�r��5Gjx�$�qj]C�=�Һ�V��I2�Kme�5�ov�Wg��c�Қ�eHn��!%eC�j!�"�v��+R4�!R�-�a�TDDFY�5^�ڍ���k����ﾰ	 躪�������@�_UW����}�}@ }u_Wwwu�}�  X��}Kܗ.R�r�K̼��-n�kE�:��T�gI!.��X���1� ��m���*�B�6Ո�Tġ]�嘓X�U�"?��&��-�B��Q�d-Pm[�Z��tnZ)d�C*�c�D�U\�����n���U[J*$���m5�4"%l�c@���ZP���Y�'��D�`�TW�:�+P��+�)h)����
�Q:�B9F71&	��F4��J+mBt�ܶTI�Che��\)Y��,�&1e)j�bYJ��T�:��G1�Җb
J)`����("&n<��a!f	D��:&' ���@�-H+R����E	%m�r�qe!d!H��1�A�+i�%�!����o#DqV��U���Z�e[q&�I	�@��̤rȭ�EUI�Q��YGcI��"<k2,�F�Bə*U��ʚR��n�W����P�C�9�	UUN%��#x�ix92�+����!�p�%kiEt�x�Uu]�����V�r �h"��˨�^�\�<�{N��_zi�����v�Y}�FmA��:]�⺥˴�K��NA[X��1$�smY
�/u�R�����k%by۝�{���$2YwwE�#�(|X��њ!Af��m2����:S�I��~B^�Dn�ʍ3N�`�C/�����3�IZ�s���\(�JD�f39�&i���~-k>����4�=3�u�!�=7�6��>�}E)����R�Ҷ`�>Մ=�q�ŵ��<��$�I.��_�2Dhx\�+��=���#��M1 ���� ӄ��Ke��[�Z�h��u�8�_.%�"�J�ˎD4=&���'�h���		VRYg9���BDt�L��g�>�[�%�CL�y�Ó�~^g��eԭ?d3�[t4�E8C��e�#��#|�&�4�*�pr>� @�����͟���~qF�>�8!�:3mͼf/π�������Ӑ�(u"^Z}�}���j�ۅS}>�x�/��Q%y�C���Xy���Z!�礔=�f��t�)�<C���ſ:���uӮ�Ʒ�R+��̼�ҙ�z���А�,��zd2��i��L�3�8t4@:pt����-ћh,�����IG�'��xgO�Q(��JS2�/��*Ɠ@ӑ!�(�#�XԬ,��2��V�Gч�6mL|�Ѹ�~4d!h�g�~|�v9�88!��+�*�pp=>�ѳ�B���U�C�gJ6Q��bv7�J)pE(�cQ�������_b�<1<o�Ϻ�l`���Ki���q�[�Z�kG]:�Mf�}R���R�d�>m�!��p�Mh�~M��26p�(��c�#�M�8����l�)H����R&�[,'���i�:B��uS����g:��V�h�������i9�S�A�9|9N�ٱ8C�10%9��|�2��*{d�a�~c��x4CuP���L*���%Mi���,���~p9w��lL�n�|`�b�&�(٧�X�4����;����8��������>4h���Z-h�]S��}��{�+5Y�s����MT8	��KjL�շ��x��
6kU��6��R�eMԥl��,�.d��I��TTV���Nr�d�2�s�v5��}��ԭ��������u-��V��>��-J�嗋im*�UU��3�gTft)79��.\��b{ER�l{�J�c�ߥPe>�W�S6���fF��%��򲜨��ON%'�{W�2r����pGs����\vB���9I@X��迿��D83�<d
"i�=�ʸRh������E���C�`���]V�'���uM��M�D~+�0���ߚ۵�S���J����+�kG2���ҊR}�����F5���C�-��Ӄ�#��F�:뿉�D;bn����zn�	Ν����4h�7��p�ç�1@���fKa�e�xO~��.ou�[�:���n� ��Z?T _)�	EZ�i֑���[�Z�kGN�N����M�܄rciXE����!�Y�G�',�W��e�pς�DA�C7�qam#��i��&p�R�C?|G�}t���3��KzI��z�?�Y�Hɷ[)�\&1��
˳Y˿�:�GJ<�N��u2�G��e���+��iq�B��%[p�-��쮇�n��h��)���f�u���m�Z6�~ �y�UT�ǃ��Ġ�5��P�!	L�z0?<r�!	��:��^1�}���[����L���u���8�-խh����uM��z�3,�rFF��ʳ�u��l8oh���LtX�tJ�9=,��8B��2}��|h!<Q�N��h�l8C�5o
X�m͂����-���Rbm�,:O	s8&s�a��)��0|!�C����Uc�R�S
�}��q��(�y�e��=>ϼ��@����B�	g�B0���͒}��.�
Hp�9ѭ����7-����.��m�x��2ʟ�F����9�_�Z֋[κu�8��J�Z��3�IL��QQZ�IS���h��I�N<1�����t!з~0:~��<la�X�L�KŰ��S$��Y��n,TQ-�S��P~�i鼦��@4P�O��{E\�yE������
k�R�W��J~}��&GC�xh�jHw�����RO��g�Y&�G�uz�����p4ﳣ���FGG�$�-�F�CO�d<���zt8;$2����)�iykq��V��֎�:#�^���V[#s�Nq�d�1�}�8�yA�9M�&-�K��/�qWQ#u�Wb��&�$�M�����Y�֊��А�������noB����ҪY]���Y�Ź����7���ɮ�g�#��9�/:x�o:?x�p�r�oC����Y�)��ㇴҌ~_z}p�O�X��j/�z6�!;���j�)�cܵջ*{�`���sE��=���ӯ�a����¢rN���k.�n���Əf��8g�l�d4㞇T�Ϊpu<W+�|CF��!ޓ"��a�b�S��p���!W�7!04���r�����T���8k;�/����|0u���$29�l��&��Asq���wR΍;}AD9U˛/��T�q-�2�ީ��_uV��^~2�.��ҙ���qē�&��US��/җh�����a���y���խh��p��fYr�IL����kY1�EI$��T�n�QQZ
k���_j�hʗ�}�������f�D<&�HHa�S��я>9��q�2<����i��i�i��~}�ܣ�o�9K�u��U�h�2aJ}LcϷ2���#��ӱ��m�9���փ\��`�i*7�8w8 ��}�[/�pڔ����*�~��)�Ĝ5=��aGz!p۳��a��N���P���`6��!���~ʿ|�i��u�摥���RȈ�e�GYB"��Dq��Gu��B��!c�Q�eDm��yu�yG��yyF�Dmu�P���#H�TG�i�"�FQDG^E$���DiF��Q�"(��"4��#�i�֥�m-kqH�#���4�#Jf+�0�*UeHB�!�T�E0�ɤZ�[�S�y�]u�V�YB"��DqG�m�ѶXB�!�R�aOߛ��^���q�z�m��}�M�%�P�&�E�~��6{'��s�)1t��s�an����:��U���Eb�-n�:�][11ӵv�^�{�{NA��'g���|t�N&�	Ч��񑎣nW���f.�������vjtڪ����.:�l�����&�QN6��Xp�ef�q�*R�w9��������k�q�ʫ��ej��Z�..�E�2���( ����˪������� �����������ﾐ��ꯧ������@
 ,
�����<��y��y��[��խh���ÇpM��쯷�TTV���z�۶�&�h�^�g�{�e"�����:8<2�4y�g!��Y�|X�=کZ��~�����7����a�"�톂�~~�l`�pKȆD�jK�#Q7!I7ә.��惤()�ۿ�(~�4p��쌇M+���;h!?=�5$3�BJ됍-1�qw�����s	7�ŭ��[lp��9���|~��.y�]��d`���t>r�842⟘q���i��u�խh��ÇpM��V�^�2Q����)d$${�EEEhH5g	�m���J��\�x�����>`���)�ّ��)�TB�1�ʚD�[PߵFИЈA��,RT�иjl��/LpF�0-orl��u������
>4�a|���Q���|K��Q:,8B��EUJ��ˠ���4;�>l2C�f4���}�(8C�'._p�+���F��HC*M�"�|eM?��L��uim<�:��Z֋Z:�u��j��w����8k<�1��,*��u��o{��!�C-lr�U�e�8ڲT��W��G�N����$���k���6L����oF�{�yKF�N�����4�t7<'�þ��{�����{�l6�h�\+��%���zrk<�9��T�8h��&s�ŝr=h����﹓r7�ʼ�m��Z����x܂���ѷ��c���q�V>�2����J`�'߾}�}���_:i>��xs�f����/��RZbzQLN~�ьt��a�x���ӗ�6&M7p#$�'��o=�����pӂ/�	bK
M}����B���[�SH{�
!��c��>6��$��GZ1�!		�j�b���W[$>��4tÄ[�-խh�����Xq����L��i�u�bXՕ���6���%���j`jbq�ّÖM��`���fUW�i�fS=���C��ۄ$��D��'�f�$�L)1Gx���AW�4P9[>:Uvᢍ���Cm<�:f��L��/�5��CJI��O�;ݺi�8V�����)��e)`k7Y��M$���O+��B��Ѓ�a�1�Eu�0h��,9ԣ��ҚS,6��o�?":��Z�:x��f͐�F�����H�J�+%E.\<����	��b�j2�yA߁���
�������I8m�>ރ��i�9�w�?��i��)�b�F׸i�q:����[�%�i�����b�|:u���?Q�Έ�l0|�lvg�\�>����{�H.}1�s�����0�~���g.%�ѥu�E����O���g1�@T����|e
:�	~1&��)�m��io#�?:���uӢ:3�w���U]sS����BY�x���ЉZ+����8�q�0H2)�#7AQ=Q�9��M�h{Uggj.��'뒤r��'H��I$�z��63��'{��a����n̧�|��TI	lp>B��M�9l����2l�^���IM�xx;�4:6�|2:i��0�Bjuӧ��u頇@ၳg�:}���2P�G��!Zц���n4�����Z�k>:t莌�Ȉ�9~|/_*9�ʄ��UC�����<��b� ��{]4�3�o]K��H�q���Ѵ$\�3�ﻴTTV��<k�Ļ|w0�>��ߩr�*���77�jF�G&���"|���S��V_��կ���˹DoH��� �NT�[3��Ɂ��JeAw�j�)f.ŕbɒ�C��!>���"s+����O;��b�S��p�ʹ�UQR�/}�^�FH�%��	\2���j���;ne?4���r<��|Q�^��$�G�A��уͥ94ڿrϽ�Z͍&�ȸ��)9�+1��]�xI	�6t�����*�w����~���fOt���-��&������>��Ap۞����iXݳUЁ*FF]���$���ki�'�H^ç�Ga��SJ[��n����[��kE�8C�l�(�I-xFy���	5	5�����М*5�kf���fp!$���!�.	�-D���duRJ�	3��d$+�ה��i�;�Q�o��ћdB��5Ŷ=�s��L�+�λ�%�ș�O�dh��3�<l`Q�aۗ��$�!ǃf�=�/3E�7��ă���Tn�f%�¸�Cȯ���V�Z'j�L��>2�8�n�'I	��r���c�e4k���m�߼S_Q�~��{�M��F��daL��l��K[�κ���u�T�7Y��+*g8��D��w���5q2�^��mGo�>��>�3�gP���7�x��AF֘��i�n��D=��j���:�81�C=�|�YvU[,�prDD��+u�I&��^*�Zhrdl!k���˷#���Y��c�
!9�c�&��cs=Q/������M�x�wV�*���5AF�8�4u�p�ƚt��ߦ<����G�R0���o4��պ�ִZ��]S�8��꯵�R�Y����(��فS���ƍ�Hy�'��TTV��%Ht�4r�����Vp2h٧v:���*��v�`��8i����E�Ebfĝo*���%�1U%r39��$$����@��>��u�_h�M��Q_�Wsʼu�F
8S�!�#�ea��H>0�4|f}����[�c��x�Hd�"�I�B��TpXq-4C��e�r3c݋�c����C�|?Q��4�c��c�ɮ�:��r�q4Q�Ř,�QZ~i��T�DDeGXB���"#�#Ȉ���Wm��!Ґ�Da��eDm�u�ym�Q�G��uDE6������"��DGQ�y�Z")�e�Du�v�DmF��]eH�U�i�y�Q�E"#H��0�"#��qn#KiKi����J��qR2DS��DaE:�n8�����+-jZѤDq��o��6�B�!��)M2������7�D�9ɫ�]�jF�(n�^�k���ʪR.kUػ����l�͊����{�s��{�y�ƞ�{����M����./��D$� �=�Mٜo$���kz�'����ת�d�~d9�����q�m=������v+�P��c�)�J.T�}�mZ�D�4H���kM��'��*�#��4!���7������߈x����_}w��;��Ӄ�X8y������Cev�(��V��Ȣ'��@�N�/6�4^��5��M��p�5�����zo�y��w�	���L�>u�C��ַ��;�~�kcݑJ}Y�H�F>N��c�'�z�Q�ىWC���>��<��|���B��j+n9D�CvF�n�ǌC����؝]�)�'"�Idc%�jY����.Z?7v#iEr*��KMƨ�+���tֈ��Ws-���mI<O�nN<��yof��˝7� � �
 ���������ﾐ �
 �����������@�(J����������  �	*���<�rk�.\�rŧ�[�qխh�����Xq�u����dcZ�EJ�(М��u"׉�$�%���p�(Ӷ<U��q�5!J$'%��2��VR��&'��B�2cc�qeɂa�a�d��,��v�b�DY-&:"�x��uR�
����($��dVb�؈"�D���E�j�-�,���I�E$Aep�ư�����Z�
S��r�0�i1��Ai�����Yq�(��б�`��T���8=�Uf\U,��!K�J�)HJr�r�K,w�1��%N�6�6�$i�E!�ĥ!!
� �X1�b��+�*"h��\�(���r�Z�ؓR�A�TQȥ�ƢDqdj[$�JBEB��Yj��.]�t�¨"6��QURj	5+"�;$��n�)bE+q��&AܭY^)���RA[^(�%$��!k�U����MZ�SR��6t�d�ܑ[ƕ�Je�d˂ɒ7=:���Н�{��繯Tp�Y+E���ݿjW�[�{
j3�uڅ9U
�2��8ɽ/{�K����E�r-�N{g�̧thZC�ҟ#���Y��v����uFf�����O{��u0=���.����>��;�7��AL�\f���9��zٳ���d��тO�\�rÅ9:`,���BH�C��bl�S�c���!C����3tH���*�COʚ:t���a�`C�6���4tz?i��'I)�2�H�xp�i�@����t�W���J[Z��M��Hr�M.�>4<r̕RV�A��ѧZ9p��u��UӍ)�y�q�矝[��U�6p�	�V{V��i�&�SzC1:G�g�w�u���_om�˞��"�i�	߽�TTV����e&W��`Rw�;wW��]l��>�t����L1�����u�W����ω1a�t��<�ۡ��À���p$2��뼘q��h,۷Fj�:<tόA����-������N�6�Jb�39ٗ#��&OM�ݏL�xzJ�����8�M�lh���vSY�<���jb�����YL)l?8��-�~qo-h����pM�oo,�V�Hý�**+Bk���gN���U#]�����x�#�75&<<|E��Iڭ����Bg�@�Km�ݚ,�Ktp8?��	�\֑֦��V2 ���e��Հ�Oξ&K2S�&�>
>�$�t~��haз�N��Xjʟ��a�v��zW���ʪ����-�^R&�?p���0tz�����˪e���#�un-�����g��.F��BS�K��wuw.�d=4���Жs��$젧�=>7���}�����|;����N3�ͺX�1�$��q��#Cק$�sWɈ�od�`���vA���G���ʑ~s��8�!Fr6�<>�}%���yd8<6~��i���L���E�U>�&0��^*^,~6����Ͳ�d&w�A�6a�:*�)N|V���U����ߘ�+��Hʑ�e�\~G�V��Z�kGuN��7�w��g�����'rn�:qigx��4P���&H!�v���%��ܾ&���JYvԖ]�f;���Y��TTV�����Y߹���9�/��rW�޲��N(K�g%�-����?s�'?|�u����D\�k�񩆍�Q�V=��U����պ�R��ȸ�i����a�\gk����x���m��Cg㚯߳��7�$�i�n��Hi���|ͧB�g�,Fs��&w��"8�����S��me�IR�2�c.���{��_��P�G�y��BC����!34x�lx�͒�*Q��+u�Oo��U�T�fdr��!*V��92������SE����9�I��|�kU�4x���d�=c�}ze�;���uM��l������Z�kG^uN��k���u��R�j3Xw����Й�In:���7�tSe��rQ��9r�4�a�4k����l�!icN�x$cD����d�bz�23��&:|90��2�7	��:J`E��l(� ��΄�[I�XHԜ�twfp���ݦ�����}w��h��
����D#�Cn��_�vk��BM|I�#�e�����/���Hs��|a�ʺ�l�*|ٗT�β�.#�:���Z�kG^uN��+�z����ˎbcl��٫��܃����N����#UTaUP��~��xI��ې�h�����㎃&Rǳ��ܓ;v0������-?~���݉�����m�/Nni���z�֩�l��	��3<���BI%�Jl~��D�(6Si�������>�q��,:{���V�w{a��F[y�읻��aӼH�]+��S�g�،aM0�2���-���֋Z:�u�x��㵶�U��������EEEhHh���I!�6SM�L���L�}�69~ CtZ���2�c�Z9Z͖K9�E�Q�JUer��Y����?jHBC��C�!���	!ghj22��]�$�!N�x�~�8�K|��z�h�	6Z����?VW���{I%D�V$T6]Vl*|;|<�,�����@���S~�ﲉ+�px�����+E����_h�*i��e�V��:���Z�kG^uN����/��g�v�˚N/S��p��!�A���8>;�5�B�V�7y$ٌm��Mܙr^q��������47����{jmB����L;E���`I���h���S�p�����:��I���5_oYN�����.ӓ�j ���ԧ�E��=��-��T�)S,�q��o/.�u�ӜM�C�p�N��!8w�j�w�^k��)��f�f�|{����&�
�!bdJY�zi�ř>,ӣa�H�4J��4r��'��p�i�)H�,y�]���W�_d:hy\`�`��~�����p���$~	��"�3�zg��x��������R�\P���?X�o�hkJ:�4�9�?���>0�qƋ!�_�=8��neM�Ӭ��έ����֋|x�ӄ8&�&�%�T�Wy�TTZJ>���q�Fm�p�,�f�Lz>t#�2�F����:tm�����Əp.0ˁ�n!�TB���B�����B�Q��Lt�A������C���f���O��p61������>�W�]6�>���Rڙ��)T�������r9����A[�F��`����.�����~")DDG����Di�u�y�ѴmL�B�#�DFi�UFQDq�^ye�yG��yG����u��#H���:�(�##(��#���#�q�mF�q�")Dq%V�a�DF��GQ�^DGQ�m֖��}����[
_�U��BDS�a���eE:�n8�#��DRֵ���ŭ师�8�h�,!B�"�Zi��a}M}��Ϧ)��V8��[��fe[[�l�K�\�]8y�N��D�L{Y%�����)��!�����$���_��Z�NkL�]YHO����p�#U��L�*���֪�Ʃ�N�Z��+��k�o�mT�
�362��Ӯ�_zD��ڡ�g5-��0�0�Jfet�]-Sd{���ͽ�U����V�� @UT������߾� 0	 ��������߾� 0	 *���wwwv�� �HUU_|��\���^e�u庵��V�Z:��pvN>bH�zEEEh�}�2�YR��[�c��O+O�BR�9��&ˆ^C��:h>z�6�N��>��A��5�u�z�$փc���ۻn�uat]��dj����2I�c����U��I�y}C����~ѫ�+��\�OSA����S�wo����(�=k�\���xsd���!���7>�7�!1D�m<��&�%U����c_Yg���U]����u�8�.2�-�G_���Z-h�ΐ��9�Ev�����r�,��$�� ��L@�^�QQZ,����i#��$8+�����M�~�������!�Hd���NY"j�EU�LV	��N�:�hzp���B`����t�^# �@�	�l&�'o	*T+FIG��4�ل!m"��M��C�ze}�R:
ig�,2h�ι�u�wU���a�΅p���ѥѣ-|BͲ����G�_���Z-h��)��U�>cm�Q��$��$��������r��iI3JR�e��srw�5eI�ZH��Ym����m���Sbi&�K�?u��6���9��������>T�$�)�N����f��ث�X��s�1���)'���\�d���R��[�Z���ͧ}��=�>:(��a���z��Qϧ�ͳb�}U�y�f.�J���7�I�\���{�MO?����H;��-,e��y�����3�?��ϑ��c��&��7�	$'�����hG�Yfj������HJ��x?��H$�4W��<q^W�����W��N[��'ѓq�h���h���3<�>3��p!���8�4!����qH#?���g8�bi����C���;2�s�$"{��у+eDy~[�qh���<�O����|����Y'49h��6�X���y�Ej��B���OW�I����>���deđ�6m��Hvg��'li�^c��,���$��Ã���;x1:o���Y���~ԑ~
��V�(��x<�U��p9�el;L�+`��Ŵ4&i,%�k��ȓ��I$ �7��*�ˈJ�����6L:zBIC��G�!�G�������=����~N8>2���2�-矝Z�[�E�<xGG�D��{5n�i5'\if]��u�TTV�wc=-�.�_����W�
��9.M�܎Ƿ���[�$��6�t*9=�I�4y�tC�����ѭ[^k.!TUYE�E�̇Q��C����q�G����IrC!0ǽ�NQ�};7�����2���CF��	������'�u}%NU���5�6q�8�.2�<����yku|x�Ӥ:;&�<;�gnM�Eu���TTV�<V���|K�%p�����փ绯�0�,�[sD����&Gz{�G<>z�>�
���C�a�$$!��::D3���NBA>x664}g�E��*��R>ǪWn�~���8ِaҮ�2�a�͒:9�8S�!2��.cW�<0�q��F�[����Z�E��N����H}�1��v���I�Y�9�PT?�8$L��b+A��RHl"�!n.\�cY�|����X�T��ꤎ��x;5�}��QQZ7��#&I�{]y�lQ�N�źK��q��S)�؅*6|}�1���;�܃��jrT��#z�=��so:C�,4�>�J/��H[]�߹��*�u1�y�	�#^��M<��u��8��w��Uk���s�5�TMPU�[B;!�5��he6�I��'x=���!ht~~xـ���C��'����`2�+���$��%�|1��m���Zrh�c枏�v3�5��=�)�F>���j������x��>�P��c�7�%A�V�ۼ�\� �I�8�_YN���s�]��A�d4t�e�0��?:����QkG^yO1�3R�H�l�>�EEEh�IR�-�l"�$����B��P�os�I8��#�b��ccCϴ?�>(���f��;��F�xC�G�
8w�y�ͷ�=8�d������=!a�k����r��(�+��)䪍BC�IB q��<x16��ɓG$���潰�CC����&\�<�i���ױ�B�tE8C�[H���張��Z:��y�+o�8�ϑ�n��*��m��<6͹��u���IAFkr�����BB�8��0ق�>ð�P�t懷��0 ���J
�e��;�\�7}��r��:�r�.3�DEJ��u�I���z�<C'��$t������C���gL��F���$�����5%�r꯯6_�>tt0u������΃�Hem�Z~y��_����-h��(��'��nH��̌��Z**+Gl����3'd�n�t揊�Z��>�0�ƘX���v޸Y�cq�Z�,*�����Kz5�%"V�FMh,��G�'����2� f�Ui�l�4:{�c�����`|��k����MrjT�E��h����U�BCC�ɡ���rSR�p#��%M�ś��ں�����h8<>�e�'NɧfM6tx�6V}�;���y,qmqY�u��y�!�R"#h��#�!H��"#��(�����l��HB�!DeL���2��#��:�<���#��:�""<�+��"8�#H����EyQ�Q�Dm�DGQ�SN#h�4��������#.0�E"#H��#���ۨ�6�L��XF�UuK���,�,�DS��l#�)�[q�GXB"��DGV�ZַV�[l���!E�>HS[y��L����7���e��=$�zt�9���wS��5G͛�"̉���ʛU����g���6�/�Z�O��_l�"�����6{ǎ؊��&殭�|���$f���x!�N	����3�����c��k��û��]��^�oq���^�-[oW=Nk��kY���=��`3˝���Kç=�d��o��5/��}��v?N����n�f�t!�ṽg�I~��I��b+V��[	Fz�4Q<�:��A3�-)�ie���%#n��Oj��㫭����F���wM������l����lۿ��f@�˸���E�z�1�N��T(��ݛ�>[�i�]E�I�&l��)��%vUϿK4��t��\�q�IaR=��9�+�H�IX��E��]���M�T�V�wSu<�sm%�:����-粭���F1\���j�H�V4eJ��q��*셣|�?��o;{�Rn��	7�_�o�~��>��  UU}�������` ` UUQ�������`  UUQ�������`  UUQ�K�*y�^e�y庵����Z:��<p��ӄ�R$��iGDL�*"cq+U1LTvQ��BGiDI2" �JG�$�G�+r
�8�QX���eI�T��i)�Y	2UX�E\%n�H)���X�Lyq
*��┢@�(��[
7D�H%ZĠ�A�2��cnː�bCp���I�̕��T�<tpDs,P�9R�)PH�7���Eb��T�Ij�\�x:���!H�P�4��X4� ��uQ��
�	֔�B�	�1��CP�K#K�LBxX"%$8*H��\*h��pN�&Kr�"Gm��pHB��(ҶWU��!�Z,mJ�Q��E����6UHm�c���K(Ԅ*u�i\v�<��P�IȈ4J��U��0n��BJ�ԮER �*H�1m��쪺� �"�t����,HLw+Q���Et���u%�N�"�D�d)MH)6�Đ�E���c�x��-R�3�����!�y��^~���ﯞ{}X���bz�U��ڣhk���Ѫ�x�K���w�7�Z=�t�G��珁+k=زq��7������/2{�t1�q��r�_Wv��:o-R��7��	y�����M�N��H%�l*�s,����~s��o?;�8d��$&��|;���)�(�h��>/�|�1����nO���t�W����l�'C����SHk�H�6�a��2Iׄl�`-�X�ޝO��>�d�V�>���A�w�[�b7�း�ė�Dt>�I�����!15�A��u����S��[.4��ukykq�u�󌷭5�^��ᦱu�8�'&$,[��&���hHK
f��A���������r|Gcmo���h���Y��#5a%IS�%tjd�M�GKR�h�²��M���GE����?B鲶]�>�|��VJ��ŶD`�x�+{�c%彉����$d	��������Ym˿�����G�z}��èi�ǡ���.�%��̖l��Ȏ�-��Z�מS�2����$�)!��HHK3a�/�J�9Vr�����K��a��WԪu��a�C��x��967����`~�4���|������:t���#�������t��g&����|u�k�6h�z��7��S�fI$!1��e.~�V���L��A^I���I�J���d�+	]��ܒS�as�V�ϳ�u�L���/2�O��q����kG^yO8ʴ�J�:\��[�̥+:�o�}�uŻ4�`d�߉��ؓ�	�K �9��ϋ[�H��F�Mkp���M�|�����J�dphHk#�6���ъ1K��fx�W����J p9ޤE2 ک�?I�BI%�l2.��h��rhl#�1��l6�D�����5��,�}��mF�SN2�.4�-�Z�Z�E�y�<�.�~�Y�3�b���zZ˛��Ry�ͻ�����Fmg�krj,NF�Z�r�M�J���?D$$%�*J[���?|���d�ww�{�)�l�9Ԓ9itҹ�g9X�֙�U��ڕ��Ε��ϭ�*z��
��z�ү8T��.�R��Z���ԸNL�0<��*m��#�UrQ��A0�O���b���ʿru������4�,�m+*�ɯj���q.a�����{�����G!%eݺ�M=t`·P7����X���O�o��%|%t���}�;�$���б�enH���c<0����T)�4p�s({�L���t���1��ILI#��k�[+��+�[=�g~�*��U�2�NaN-��[H�q����-h��)�o5U�5��T7�����Z�u			a�̱�d�c����O�����T���D�BT��O+A��1vضKn��W�d(d;�MnM�&ކ� �v����H���bTǓ<tHB��$���	`�c�N��{��g�iJ���o�	��:�p�ز��Ӣ���'�ŵ��]H�$l��[Ց@�FU�w�<�>h���Ak��U�|�~8,���/�<���[�[h���<�v<'��EHU���R��$�!gڄ���]r5iEV6V�?o��#�>��WՏ�1�d�æqB?}S���FsS���{�VJi����eZ�{�i�:axZ�?~�K�u�c�S���l��3Á��6ǣ�81��c����7�����N����]�!f����?u		/���<�5�+�����^�,���e֞yE��Z�מS��3}���Œ�,{�HHID+���j���gk�d���n��B_aL�ǚne���K�d)Shd��YN.�cr21䟁a����3����.�FHdq�����RG���?K����õ��gL���j�<lL��<�c���p0pr�g���	6}���w	6��%�6�P���`<<�)�4J���T�l��4���Z��֍�h���<p���~g7��_��Z�V�"j�I��w6�ɧ
Cb��C�Z.�!)Ǘx�MJ6���ͺ��E��!(�_���-T�yk�W��g�z�}�����)�E#��*b-��S���Ss�U�Ew-T�
7o^��Q��Bx<5�q���=�Ow�8�W\҅�(���N8�>�ӡ��#|�=~�~���{�ݢ���x��_������Vz�B�%��J�H}X}\�L�Jv?���!����/E'��a�O�J��!��>��vՄ������,0�T3�k�O�:	x<�^�%�p3�I�3�$0_�<�·�^c>a�����n�2�����"��7������FEe�٨j.3N�9xBd�s�����������oqL��2�O�~qk[�Z6���<��e�-��f������v'�<0���%������6!
�v�nuQ"�譟T:>z�	`�.6d�!��Q&C-���t'�NcF�n��0&hp�H�8gs;ڿd5�\��)$���a��N�����?d��wWn�:>=	y�U� Ԣ'ۥ���cC��8c����Ό�y�[m���Ƒ�,�)�DG����"#h��<�����6���P�!N#(e�UFQDq�]GP�<�#��<�#Ȉ�:�u�Di�F�DDyR�a�i�Dqב�mG[GnUiN�"6����B�lB-����V��j�m�g��F�J�R�,�,��E�L"2���G�]u��GB"0���:��#�[�,��e��Yd!�YB�|���S���~M^ܭn2���m�fF�[i�����ʛ��ڣ���_V=י�ETq�ۛ����;z������W+�)�|�<��Ċ�E���s��˵z�>�9���������BSc�)$&�t)�n{�r��h޵۱��/x]����;���>��$������������y�����t�>7�d��~}�����>'i�*�}��v��wz�ӑ��\�S.�����!��R��Mܨ��}Zw�}�� 4  ����������  Ѐ����������  Ѐ����wwww�  �UT|���y�^e�yn-kykFִp��6Y�}*#D~�$$$���r[WVʻ��.������'c�|[f��a���J�=�w=y�6a�ydgxI2���w�f
+r��֬�f�4�3s���L���3�J�a)ɳg��)��[���d$�����_�5�OJ�|t�͍��ڲ]5T0rx��Ӂ���mv�xɇ]6ҝF\eZ-ŭo-h����u�����U+�f�UUUG�W�}�l��S*��S��뮎��xi�5�SFe]G��l����4�[^��e�>�|����d�eザ�e�2���`c'��;8i���!���a�ْj���5"b:.�!�ς��@�����e;F�HCCXd��b�%��������Ҝ8B�)�YFQ��n-kykE��u��<t�"��_���n�`:Q���Xڔ����i\z��4t�2�7�ӺN���#��4�M�Q�$�DY�A6��%Hi��le�V�q$�@�q�g��S��<8y׽��{���CNt�g�q�!���t�>���3��w�N�|��F�x�M\8u޳gd���-�M�w�N��Mw����W�oZ����x>+]B���E.������}�܆t7�5��t@n�.��d#�(K��P�$j�=
�}�s9���yxW�IU��Y\�GW�Oק���<�J�Xa)�/F]�I-v�'���!64l5���H^�3���U#���h�ƫv���ZU�饛�m[�\�A�ٛ�\teV�������)S�XS�2����[�Z�Z�n-y�<�)�Uk�j!Q!�n+*����f�X�$p7d����nI$���rO����zHS�a犖<nBI�ēo���s�9(�t��J��IX��pzm�`t8�hxp�]$	��nC�8���z�F�5�t�ޮ�tF2G�Ι���F2�S��KX�m��64�϶��U*��e�}����{��E��O���$���sr0��s�Bd�P�grʩ5�Ď!�'��J������7����jyl�2������ykE��u���}��FkY�.�����c�rI$����{��
�5����e8:4>&G'�>��ߺ�H���u�z��p�����n,���M�{Jk�ɱ�۹�y���`z�lh�|pўɊ�4�O���5����G#���8J��h<��p�K�I��W+���\��Fܷ���+)��?83��O�2Ge�V�ߖ��o-h�֎���!����?�X�]c!�D����bI$����7|�$�M\�xYܧ�r���E$�Q�=��~�*Z�pٺw?`nb6.�̧�r�EU�F_�`q^��xa��=CM�NrM��j����/�®��L2�s����+�z@lk�+���d�2����I�nN����h�C\��#�c��3G�\*�W\?>�Ϭ����u�斈��o-|���7�SZ�J��=u��d]LL\*rhSH1iE8���J-���]n>r��Y�5yĕ�m��J�q��E�1�+To�I$Jq/铭/�ڊ�]V�b�r��z���ż��M���TtX��=[��dγ����S�����>>pӚsz/dVv��;j\gAV7J1��"s�
Oj#���)��C�����'d��G-�Tf�H��J¡_+)F���l�I�ɲ��;v�$dãC��P�UI��,�Ӈ>4�ӇJ��?N=�W5c��\�C�`}� ��G�27z��BT+#N���t>�ǧ���|d�L�Yd5�;2@�����UC:��dUP
�T�������-o�7���m���kk�pj�,���[o�w̱�E'�G�[S���+i���GQkE���uN��T�K�R�bc��TsWx�I#ً8C��Q�{4���}:t�8�6k�Y�)cp������p?SƓ#��?P��P��Ӓ�h_���zC
���W��:m��j��1֭���9��n<�'�8N��d%]����$�\w��������-��S�y������rI�>m��G$�EvӒ��q��Z~">f��E[YI��$��C ~(�<�l���~qh�"�l<��S��0�OI(�I��T�U!y�`��Ȣ0�����~�$�C���t�!���ݜÒC2N��H;�h���L�xl�=��h��Ӆϩ��#4�W���B�5'�����鴱�H������sHo��c���͔]I�G��L��iކ��Z,᳽�I���$����I��&���v�K�I<_l!��.��Ş{˄I���7���I҇�Q��[*i�_�~i��~D�TZ,��ӄ����Q�f�o��RC��I�폺H`z�o��S�h�������J��J8��i&Em�F3��������3��i+%�w��`d(�BU���1����&�Q*��d.��p�x}���?B�3|�N���I	���xv�KGB��h�������[��הҖW�U)UF�`\O���w��羟����w��]/~nn!1 ]��g��bҘce���6%�$�!�={{���E� ���DA4ZH�DŢ%��� �D֖��LDZZDւ"�De���MD�+Cp��4$M---&���D�$�I�$�M�KJZD�E��i����%��E��M�$�x��ȴ�����-&�-$�i%��Ii%��M,I��I-$�u�β&�-5ۍZbhM$��d�m��&�Y$�i�KH�%��"ZBI���I�KI$�I��I$�D��M��I!$��4�i9�H��I	%���ZIi	%�uĒi$�H�H�M�M$�I$$��M�$��I!$��$$��!$�miii	4�	���BI	$$$�I		$$�M$�m4�I���&�Bm$$HI!$��hI#H�H���BM�"id��i4�KI&�BM,�K&�I-$�&��--$ZZD��2Iii4��Y,M��E��I--"m%���$��I��id�m$�ȚY&�I�Iid�Im,�I-M�ȚH�-�-�kD��KE$�ZIi%���md�Y&�D�ȚmdM$��M�M"$��D�ZZD�&����ZZD�M"H�Y6��D���C���Z"Ih�D�KD�E��֋Bh�Bɭ4�M4�б4�D�MI�M4�4�M&���b�M&�#9�٣Y��#[�#F�4h�!�g6Ѡ�l�cF��FF�4�f�:�fF��fF�#[4k24�24dhhW��[�:M)�X�l�kl�cF��[4kl�cF��LѦhq�h�ml���F�F�#F#C#kf�����Y�kͣ[4k6F���4٣i����k1ّ���m�����5��`�5��`�cF�h�dkmM�Lѣ���1�F��[h��F�����4�F�h�#X#[ml�6ѣ#k����5�F�h�m�h��m�k1b#Bd,�b��C߆8-�6!��BfB6B�Лd#4-�Bm����!�d&�Blж� Ѝ�f��Лi��M6ɭ�4�5�4�5�&�[m4d�m��i�Y��M4&�4��d�f�Y�CM14��dѦ���&��-�km5�5��h�k	�ɬ&��-��M��&�hi��A5�5��4�5�5�44�i��LM44�a4�i���LM4d�i��XM�ɬs'M4�4�N8�I�6I�Кi�4�i��k ��4&�M4�M	�֚M��M&��i�КM�hM&�i4�D�MM6I�4�I��M	�i��4�i5�I�M&�M4F�MM4�I�4�d�I�4M4�4�D�M�4&�Bi5�i4&�M6D�M&���M	��l�КM	�КM	�i�)�&�4�i�hM&��hM��&�k&��4�I�4�-5���4�B,��#!�"h�,D�D�����Z-��-��"h�h�De�4YE�4H�Z"2�M�B�hDd���4Z$Z,����"h�4Y!d<��n�,��B�dM-dM-DБh�h�HZd��E�BУ$Z$Z$Z$-2�2,��Ț-&�!��"�h�h�Z(��B"E�Ј�"дDY	�4e��Z",��dMc�r$4�B�"дdD�B�!h�����F�kA4bѨ�ZѦ�4m4i�MMhMh�hMh�FHM	�M]uмp�4kA4&��i�M	�i�4Z-@�h&�"#&�Ѧ�4m4-hF�4ѭh֍h��Z5�kF�ZX�gpۚ2!��h�D-���E��-B���E���ɵ�E��ËH�LD֚&--5���LZ)�1i��F�=�O`}��1t��iM4�c����؊�$� 
���!�`��~W5���_�5�y�~~�2}����ق'�������������r�C�����]���8?��������������?#����,�k��͛�O������kC�o��������1����������?������?�پ̳�o�[ُ����M������?������C�E����"R�+h��������?���_���?��ab��b���֧���_� ��P�_�lK���ċa?��_*a`B�?�9�?��))?�N�"-4�~�k�t��O����aR;���l�#�[?������縟�7�* ~VX(����("XZ�
��ll��,͎C3�i�AH� aT�Gm���	M3s� �����7�_�n°�� ;�����o-���l�$62��͛�9	f�lZ��j3f(Hm��#l2�k���s��� *��1k�'���X���4��@C��[�����'��)�p?QI�_����R~�P�������bq��T ��ʅ��?��k���������vG��/�k�?�0���O����s��	��'�
`���������:���o���g�_��@T �?�|#<���G�/�����]�?��@D?!��H��3��Ҡ* �����hW���7�,O�)�?��`t�����_�9O�ώ0q�c�V#f�J�1B�(����#� a�ِ�䥿� *�R%�����b����ؘ��QY7���������νlQ�m�b����q0Zk�qr��P���A?�=A )����~����g��mt�* ~��~[S�������?;�?Y���������~������ȱ�~�K� ����S��?l?{k���|3��	?���H���������O��>���ӿnl�L}�����l�Ԭ�El��ejj�թ�+VVՊ+V�Z�jիV��(���e�QL�����V�Z�[P�J(��M�R�j(��µe+j5e���VVj��V���b���V(+ej�b�AAXPV+��b�X�V+��b�X�P��X�V+��b�X�V+��b�X�V+�V+��b�ԭJ5mY���F���J��5mJ�VQYE2�)B��)�VVQ[VQYEee)�P���El+f���VQYEmJ�)��YB�)YJ��ڕ������
P�
P����j���������eeemMJ�����+++)YYYYJ����j���cP�Z�lV�ԭYJ��Օ�+VV����+j�Օ�+VSV��[R�L�B�
+)��j+VըP��B�B�B�Z�J�jee2�e5mYB���Z���[VP��YYZ����eeej�Օ��+++VVVV�YYYZ��ej�Օ���X�MZ���j��իjՕ�)�����+(��VիjյVիj�+V+SV��e�jյe2��J�V)�QZ��jՊ�VV�V(Պ�5eb�X�V(V��b�j�[S5b�aX��l��eb�L�SSQX�X�QL�V+�(�l�V�����Eb�V�j�ژ�������V+V�Q������)�Sj�++e+m[+5
)���[SVSel�������B��j�j�M[V�QB�P��jj+V��(�Z�QEիj�V���[QB�j+V�XS+R�j)��l�J)��VjحM[Q�(�SVղ���m�+QEmYMF���Q�+�
�+���X�V�b�X����l�YX�V+��X�V+�5m[+��m[+j�b�V+jڶ���ڶVղ�V+5jQ[jڙMZ��YF�
�QL�jQYMYZ��jڕ��jڲ�Օ��+(V�����
jՊըը��V��
VQZ����QYMB���QB�Օ��V+jQYE
S(��P��+j�����+++++(����YYYB�YEeeej)��Z������ee
�յ
��emYM�+++j(����(�����f������e
j͕�e5mB�)�V�++SP������B�P�2�
55�Q�+VՕ�f��[V�ڶ��jڱX�V+j��b�AA[��b�AX�PV�V+��b�X�V+��b�X�V+��b�X�S+��[V+���R�+jemL���Q�+e+P�j)���e�S)[)B�)Je��+j�+VՔ��E2�e�jV�����+jVQL�
P�l�e+++jVR��e(R�(V�e�Օ���������j���ڲ���e
�����R���)Ej���������X��(�JjSVԭYJjԦ��SR��jjQ_�?���w�?���� � T3�?�'�?D��������:��,�"�$X�U?ן���@�3&J1�Y���?��T�m �OC�������r�p%?ה��p�A��}��*���O�5�̔U4������?���Kj���~ph�΃��_�������P����̅h��~�pv������o�LF�f��f�]~�:{��q��?���?7�p�?D0���O������I������������C��R�F?�w����)��?�