BZh91AY&SY����L_�@q���'� ����bI���      ;
��$�EJ+�ʀ��
R��Rld[ 4�B�U�IKmk$��$�JP*�$_ZB�]5ZQT٭��v4ڕӧl��굪4��TͶ�MQ@+j��6V�(CZ&�l�YT�"�&����a�V�kd�������k��%�*��m���Ui��{�ҫY$�lBB�J[hk(�ԥkJ�*TtB$Q��R��TIkE-0KX!هl-�Fڥ%D��P)�6�J
�(��{�c%�����   .$�� -��E:�9�[  Z��uPt���U����vj�v�T���[@: �-�֨[�p�Eu]���n��l�Xl�l�5mW�   s�v ��hZ�\�N�ø�t� �Y�
�h���t��L�v ���5���6S��Pv�����EV����f��k[*
b����    8�� z:z���((켼�� 4��7�=^jP�<wz�R��{���G��л�k� � s��4h��'���j���� ��]��76��&V6�)��   n���Z�"�oe�P�Ҽk��z�
m��O</l�kg�n �M(Z��L� �]��P���޼ r�l���+�Ը�ՔP��:�I@��On��5U�W�  �c|CEhN�����ӗXU�1��t͵ n�Z����q�$��whj�5ƭv��j�雕�4�Un�M��ז�X��l3[ik@kK� ���h6չ.r�$
�ud�AT*gg) U�e�P�3���cn��waUT��� 7�mSB�r��H;&��-a�*�GR괟  w�
(�XklP�� �b�v�:veM���.�[�smA)g9\�(�ܷ.���suUR�N�\ �nY�5��2���A��ڤ�� `z�of�J�,��
U-m������&M@
Kr�qE
;r������B�E�r�R qv��&�(��֘�m�  L�xUP�`n��UP��"��4�E�9Ԣ�wvguJ*U�v�)�1�((W1YEUUW:�f�Y�(h�V���  ;�R�0F�wJ����PR�g#Ja% ��.��g\�(��⨥t�*�G�     �   L�)R�A�������TU� 4 ����O&!IT�  0  	��S�$�P 4   h S��JM���CC@  4i�@T�j��M鑩�=CF��4h4ڇ�w��ޅ�����䘸v/n���8�W��Z��i���޼�[�G����� {����VAS�TPZ ���ǁ?������"?����?
��
��UU����_���'��C��!EW����O���d�(�6��A�l����n�ʟ́|d_�|a�T�<`O��P�<eO��<` �|aG��aG�T�}2/��"xȞ0��	�"x������0'�!�<eC��<a�D�<eO�2��	� �¾2��� ��>2���S�̣� 0��"�0�����x�>2��+�(��?,����9���|e_G�A�|a�������(��>0�����>2��#���� �ʞ2����*x0������32����*x�>2��)���>0��{a0����xʾ2���� ���0�L��'�G���|eO��<`O�P�g�A�9�|`�A�|`G�S�<e�}0��#�����0/� x�>0/�� ��?l�2����*x�>0���(�ʞ2}�����"sx0'�)�
xȞ2'���	�(0��#�|aS�T�0��� �0��)�}2'�!�(f|`O�P�<aC�@�}��	��|`��<eO@�|dO<a�>0����
�Ⱦ2��ό*x��+�
�ȿ,���0��+� 2����L�� 2�"��Y�|`C�E�|a��C��|`C� �|d_�|d�C�Q�|e�>X��0�� >0*�(��P� ��<`|e|a&|aD|eD|a@|d@|dD|dP|`@|eE<eU<dE<a<aQ<e|d|d~<dP|e|d|a|e~X_�  � �|e��|`_�P>D�OW�Q�=0�0/�����>2���¾0/� x�����#���Ⱦ2����  >ox������G��!:'��o�4��i�V۹�5�g7A{����ڵg
=P��Kx應#ˆY� ��I��5���c͡�֍�[cu��8Q��mp;t��L�g(�X�]�F�1>X7Fu��!�`3cb卸uŷWCj��k��{�t�i��5HI[�m��i-���9��:koddc�H,��y�8]r:�)Zw������%m2$7��g��`�6�ʘ6b.Sٮ��Nne���d��J�SǇ̲�j�ʧb�n3R"n4ꆊ��1�߁go+1�ǐ"�U� �IRz]%��-Ͷk#��X�YU�<Ndr�mM���0��n"��<��;-�tt��w��7[��N�$��VZ��קdqJ���0,�-^�яz�낄��l�F�L؆,����(���vŢ:��s&Q�e+Ǹ"q�@��w˝����s������F�lt�\P5wtD�6n�q�	���!y�RHhv��,!��2�)��<�����2�¸��s��R[�ц�V�aS9�m����Է�y�N�X˺|��Mֻ�Dn�xmJǎ#��\�pG�洭V2H���:�Q:C����#���݇,c�Y������H{n��'r�0�4���5�p�O�1����HHNY,P��j�,>2�e�+sI"f�˴sh�q ����!:{OMzA4*�=7Ca�4���uǱ�N��N�w�Wx�e��a�T9�x�b�)�U@�Ja|���e�r��[����u�� 2m��oVպOf�mFe�ՙ���5�[4-���ۺy�5�h�KnA���e��7.VہkC3��(��p�f� ���%�ۡ�`�cY�t3*`fm�Y-[���%�F�@��e�Cr�2��dv��b�6v�E9T]8����ړ6�C%OG����ػ(#�F/6�c��+�P�y.U��#�X���*�tr�G����v��٠��D�#j1��M�u��
�PطݏF��������!ř��ݑ@#z�)7ٻSfͥ��1��/bf�R�㹌U���W�shŏ*�#^ñ���6�4L�[Y���9<��b7S������o�[��U�Y�v�`䉷�TZ˺�0����o���3�o���|<�rL�D�wm��Ee�{JV�]�0++,��+jQ�(�i���n��it�R�	n�����yګ�0����yԕ��<�%hG%7k�gR�&�}��\΀rm��^�X�ͫ;*j��6v��7��6� �[��J0���z�ʔ��	c�s�^�f3f5P�!ش�Vٷpb�E{3e
�Rf��M�y6f�Jݘ.���-N8��$y8��S�XՃC��I�(b��)(H�����4d��D��{z��U�r4)��BN������db�N���~2'�\��!������#�BK��~���n��.�<'<�Dj۴-))mk���c	�62SK�́m:ʙ�oG8Ȣ��yO��!<��2��:��m�0CYX����o(`�p�UpX1��l�\K(�ܼ�y��Ƽ�'���nMuln4"�Z�� �Тΐ���B�2��'}.[7�7�V�Ɯ7v]���8�m��gK{��Z��h,��ۃc�fb�d�J,8��V���Tv2Q(2D�4�u8�w.m��s����d�VM=���bX��w^r�)d�ɛ�m�e�1�������!��Hk\R�-��M�)Z�b������-�`%�h�3�,�f32�Yy�X؉^),,6,�h�[��LV�Ttvf�T�cE$��v�?+�9��D;�e���;��Ԍ�ܵ�A�̼{�C�oټ-�}��;��J�Z��,�7���j�ݓSsA���Q74�঳oۗv�˧[ё*�꓀̗��8�X�$/Jw�X��QZ��4*��~8*�����wǷE��Y��WD�̂�k���cct7L�D���������T.��+w���\���;o��jMYڰ��S5��Ȅh�nH���Q�Pt!�����D�#Է�v(�8EX���w�h:C6��Jb��Ge=�.�����*D֪�f�cB�{׽ٜW����34L�ǔ�z�ӄN�-�Ѳ�d�(�qQ�޺:l�#�c��N���L]�7e\yx�݇��f=�\5����J����b(����{�1�]�Slq�^��!�6�<�f�v
X��w��V^����i���) #��$+�:�m�R�#�
���ql2�H% ��frj��+��SȢ��]y��wք���)��$�զ�"�"n�]�5d���ͺ��5�Z�sXÝ��:љ��((�3�P���n��Bm�ʍ5y.SiDhk�h���ܐb�pu{�b�"\ݔ]p�l"��D��Aٹu��vNB��&�RE	"	0�軅�Ղ�sN,�]m��VX�p]�d�ʐ˲5�EMО�6Ǆ
yfSbP[���+G�>r����on�y��KטKʰ棵0�իkN�FSI�V�8ʁ��͘�jaA�f�9$��&%d��	��u�^օ���"Wjk�w4��L\��{P�P��/��T#4٨/Uݜ8��$i*�	�&p��#[s$��W�k~5��:U�F�?rx�rW*xE谈F&Lln­��&TPϔ�ǋ@ܶe"�8��N��<Z�ɗ78��2�&6��q�v6�f	+2�;���/k*��Ыkl�;.��w�g�<8�+)PL��N���)� ����lW��fz݄��(�
��O]�{����k5�C�sP�(�8�r]��˭��/@�9fΖf2�a�7;�66��[�}'��[u+)nM©2�-�o)�P�s.�n�8q�N�V�u��C�ab;�V#�FU�k+;�GN^�l�r�ڔvm@$e7vik5z�+Ev��<ګ\R�Xt!l�&X�4Xl�܇	�Xr��j<���mf]��ӧ�pZ�v��ܢA���˚��y�rf�2BR ����C�wj�m$��A�+,^�Wq�w,��ʨU"����A�4�Y˖-c!�c	�M�N��ά�8wh����s�=�ٮ�ज��è1w���ϟ�Bh�nk��\ŷX7�6�b�<��+S�Ln�X`�7`K���k$���,����e�Y�����E��
|n��P|�A�	�.4n˿]�e^:��[8*��)�i�`���Z�7��,Jeͷ:9�.�wJ��A��f]e r��spF���cq�x��K�4���+s�X��4�c3�՛z��&�N�Т�4sFVM���&i�~�Hr��*%����;mz�\�2�(�
`������D^�7)��$��󫞶�� �:��B�
����!H�,;Mfj�e��4�0+(�ܩ���g����}v&	�V��X��G��1줌3P7�c"��I��^�I�4Ȗ>���J�x|{:����V��7AU��b�!VcX�f�<�d���8�n��f������L'�L���G�\��j��nMdN�L��"�D�����1����3g!,�w@�zFQr��P���܃VV�6�QR"�r&t�0�vK��M���C����sR��Ѱ=�G���y�.�P�س@�'p�4�b�Q2M�ۤ���?�p�So'�9����Yb�*n�:X�{��8u���¤kc"�O�Ū5]8�j�q���Ɩ[ݷ�M� x(�����k`�4���/���Ӿ�J���i1}��5=�#��u/T�Sn�G��LL�ML7sii��5�Q�g�T�ڝm͵���t�M�GO���a�������9����oE�� ��-��-�)�g�J'ף�J3gt�XVF�ԍ̠3��w�%)�Wy,<�l��S~��H|t�%r
�$;!Ř5�si���z� H�ֆ�w1ˏot���w�Y�����nl�����;Q��(��e�AH7%F�x���.�-�����Οf��E[����k�s�S
�	�v
��!�� v�Ҟ�w7(���-S#��_M���|�r�(�2Ƹ$�ŹKFk�)-�ʬ�`��&�R�I�H&�S�3�vC =L�~�1����Х/��	e�1��T��i�yS7v��C�X�1���d�ݼ���r����IJ���z��2<n�C�X��Y/;�ȅ�T��4�'8enn�$����F,��%�f;F��Qf(���MS�]jT����T޻ժ1����PNc��M-k��e�zr6Q̕xM��/�}�7r��l։(�%����쉝���!B_v��D�ԩL�[�mԊ��[2����)8�4��M^p��F���k�f�'ZOi��z�|��iC&��q�v1L��z�9n�VC��1,q��X�)n�w�ח ��O@C9J�Pt�x�����4<�m�+E�~7�Md��zo4�B�Y����77f!�te�x�47���H��"" DTlS��mƶ�%�v�"��dS��Xh�o7�2�@3��꯻i��R�}��wW� ��	B�۽+�JJW����y�6�]��`F�{�;��!
��1`�TT(����&��]&�MJ���J��1F��u�.�
f�L�J\�B۞�3B�7kC;���)�ˋP� `�6�o)����fRR��Y�,)ԋ�O2X$4�����P�2�4fY���Sh�$�o!r2S�e��Z��Q�g[��Ym���J��G͑���bnnc���x��\�:�i��X0˦����ky��2�Ʌe[0n�U�t�LRLc��ܛ��^W%�h,^Ly�Z��c�-�ZV���u�H���J3Be:P�i�^�
��n��T	�Dه�%�P4�2�EV���&�aIkZ+.��
��6��+����)�!�����L�OoZ���Hv��m�̈́m_�	���q��1']�%�����2*�W�X���	�R򉶥��f٠na��G�i�-{SMʂ�]�V�;vJyE�;YR�rS����ou9H''d�	�]�W���/ۗB�*-vH�ݻ����v�0�
�Da�FM�ONq
��Uk���͊�R�l`�P��K�G��x��W��Yr�E�&���`ѭ؏j<�4�y��K�-�z��h,���)k�&Y�i��H��kN�3�Ӳ�͈u8%�h�K�8hPJ��$�o;{8��j]BSr&���S��S2/c��[����9{���^�Fc��-��Z}:��+�<ƞe�d��-�i����
�1X�?�k���PmC+��@/�ȍeuG �vB�����6��Qׁ��Sv�ӲU��n�*0�5������.0��wGͻa�B�Ͱ�ʼ��l���L�һm5��f�zm��{ǔ�&7t�8��"V&�HSM߲��5��#j�	��t0���b�S�Yv��0N�8�� 5BU�C@㡸���B�g8�=���/e�����!A�`$er�Ѹ�qwyttL����^_2�FZy���n1Y�yiz�"ye���6tE�"T5 ���yY(��9���+(I�Z��!�FTih&���r��k����l����3^<ՓX�-m�k�R�+�B���M�w�e1�s(j"1�eVݘ"TL+�u�jƽ��N^% ��S9{#�.�)\�X�:�#8+B�R�صSՖ��I-��E��Z�Lр
5��#��4�Ym������j�J�T�`���\�c�c��z�e�&��k(���$���V��6px�Y��)��KRE
��˿l��l<-�S@B_�kɛ����-��Qٍ�f:�Cr��s/6�Y%޹�la	��m����S0
L֭��Wf�f�J}V��X5Q�����LCd�X������,�V���&���S&:Lzx7����3�d��jAD�#�W��f�����
f�X�""�qj�����,��u����ݓp^�;�%��[S_v�����MJR?8��a��9��u�n�ǹN�΋[ٖ޹�4�E�i�`�2�V����X�vr��&`�*������o�twL��fħ�<�L�Y ZיL嗯2�$f���Rْ�3(�M�2��ht6�Qҗ�-�Pc��n:�r0nn��)i��d���wI�+O0՛/.M����y�Tgs�}u����⃞�<�WK"N����3�L�!m�2Rxx�WbɽFg)���ؗc���onoG�
�鉚�]''e�U �I���p]�|U�Ui`� 4&�m�n���O&�Y�M&�G�\�n��FRt�nd{�.�=���n�����;�v��-:����8���[�2\��������WkC�z#cd��ı����&�,�$RK,���tU�Q6���/�w7�x5nj�1N�RxW����f,�S�7����B�]vA/,FcY6 �̼ژ��b*46�R��{�UZ+Wp�f*B��^"��e�!gv���	�����hR3Qݥq� ��:��
�#Iq\�8��M�Q{r����d�1$bqw��{T�MD�*A�]I�.[F.ż��΂h'�m&�����r��p�EVċ.ťI�!�DYT@U�3�D��E�0ݖ�ô�d-q捋x|��H �a\����I(R>��l�d�4&I�0X'����♥F3e�x�+M��\�(M:�Ά6A+��	3P�;.̢p�`XGQ��k��3h��oC�6)�m	  �H)/D��� N�H.��.ȱ���Q�C�,��1��д�KTIrz�h��X4
#��*���+���� ު�M+�Y ��u�*L
��y�/�mi<�`�,L\��p�E3��2�pN��T;GIQSY�	i�Vr��DE���*����T�ͲQ4 R }EȽCd�+��l�Xe&�h�h��r6a5�.YXF��&̠p��X�%Z8	@�`S�gt��ʫ�|�6�_1�_L>��G�?Ʌ�ߛ�~�?��X|}�F~�K~��;����m��m��m��m��iOt$�l�-��i�m��nm��r�m�[����6�x�v�n�m�m�m����m�ܶ�m��Ӗۆ�m����m��m��zL'�j1��I�iD�X�q5U�MMIQ�;-n;�e3�4��Y�����!B�!��j����-�S:�#s(Z^ε�2�vX2�7�����O�13��2u/I ���u健��)NT��=Yi,[[l��5[;K5N�\���#kU�oI�����N�ܨ��x�څ�n�Nr��,z7K�u�Td��Za�owX�t�]{������g<�E�5,NZ��ƫ[[Ԑ׋�y���v	ɇ�v�_[�lv�ܴ�ݫU}X{V��2�J,�V1�P�(k���Qd\��p:��®�\Ϋ��M��_���١���7��,��W`���V6���G(3ճfjĳzu��Y��'�Hw��-�'Vn+r(�Lʁ�]9y�>�޲�iM�}�a�k�l"4zhł˭[��@��N�A�h���i!����-ⷍV�8��R�#XM3�S3j!����N��t���1>�9>4�'tMk��ӷ�[{�	[k��6��&�V�p�^��E����1%�|��'P��Iӡvd�U��1>9Q�Jhc5g��-�aÕ(��n��z�	✒�ak����<�*�{���ђ�X�gmv����l[h��囐0A���eՄ�r�;�.�;E�p�Գ�e�~�4�0^�1a^L�Oh�!X{WV7�WD�s��Q�=9���w�W7J�L���r0�)p�5�K���!�)�����C��y�_��\�[t�Q�i9F�ҳ0�5+AɆ��wY$)���/�w>��7\����Ҝn��y�t�� �ݘ��	��^��(v.�mh)#�U& �ƶ��\���C�T�/q�D\�g����g_D��#����C�"�7��J�%�8��c��4\z�^Փ�oI�M��H�o_�ͥ��%݁Z�t�:p(����[�ެ�XU�Y��)L����I�Sr��\��k�U��.����J��drV��!J���v�I�rJٙ������;')����M雱�FBT�S�f���w���]�o �U~٧����d�ƥ����Ge��\�YS*ڔ����bp��M�n��3�����wN���g:�%,,�չ)��{�p9�[M�o��2���E��Q{���6F��s&��1X8.�o�~�S��σ��3�ZYy��������O��#D<YR�Ʒp�iB�ݒ���'�w����.�V;lWu��7�Ɏ�F):�Vر�%c���e�s��.Y��`�=�2��tV:�^�8D��󀥷�]�Q�\!V�AH܏l�À�bBj��%�]Y춧^(��z�l��V�]�AwN�BE_B���烶iƒ��B?T�-���w	�
w"MvYTO(���	��r[�R�������%�T�w�Ӯ��7-�� �Y��H@t�����00�7MbΕc;5A�S6�i�s�C���N�ͩ�dŉg�%cWgb�.������_��.7JsT�m���N���=ɝ���j�G�FP��k-�q�4�r�R+����T���a�3T������1:�]'sG��50�f��23.k�vS���+s���xM��7^�Ca�qk4��Yok->/�¥�Vӡƚ���S8��e�yu�`���W����}m+&��H�U�Aڤ�Ѷw0�7꛷Nf
�eX�9�!L��X�E���ﴦ_k/�`ryh�hw^{1wvP�� ���Сy��R�I=ôY։�z����Sd��s9�Yji3]W	�7�;�T��`�]\m��S��u����(��M$bJ�k.,la�.L��+_-���&��4�����8uY|�ˆ�fl��G*B�Uh�RK\�;�]/ll����+�y�A�p�|��=2�9Sm`���e���&2M\��{���+��<ܲ r���ѵ�Q	ֱ>(=�@L��V�2��kr��$�@�Ưf�â9S��٢o��F�wr��A=X4��	Z��C���腆��Ug
�]/��,�$�E%CC1��Gm4pfh�)��/郪�v�XB�+�B_�}��7��V�w%b�W�����4����Ԗ3�9��,9����wx�+Nq̡u.�����9��b���5�-#�U0	�Y��<JU�4�w��v�$��+Ia�af�:�X�m����J�}�iJ�[�����C}��^�O�>ʙ�JqqW�V
4�:��8:ݔwn��[QPy�9Ǎ�"!�Jt��d9��=�9��J�:o%۳��͎�%��s(ޞn�z����Qǖ��J���f��9Ӕ��yX��=^f�{����V!}G[�Oje=�n��y{V������I"-
�i۬t/&]����>APo܊����e�Wdz�vW�{��M����r�|�Y��ǌ-��ˣQ!'W��w-�-P��8[��(u��J��K��Ü�����+�13T8�&�UD�FS���,Q�ڋTR���M�鏹��|�U����3j���`���3�t6���YO���3k����	˨X�.�5T�v;��ze��x����U�z�s��T���{�4��tE�X�P�܊�"���Y{�t� ��=����c�p�����v�vU�&��3a�A������[/h�\��YQ�evb=�8R�b�����xAt6��J�18�AP���>��o��e!��,��G7�($Lcuyr��ꄛ���r�Q/:c�r���i��f�N�&Di�݅+r�818m�8��m�r ^=��d혥�(\�s�s]��:�=�u7�T��wLKH�m�<9=�݊�
�tC��f�W�e�'{P�{3WB�B)�w��u8���%׏6����4+��5���ed5��R�f?<��`����L�qB�b�RV7aµH��:���1a���u[)�j�U0�dY-L㶛9�V���.�jĩq�Y�P�K{�+]i��WdO� �棚%����p�ӷM3���ө<��-�sWT�n�.���U:-��\aBUvb��epݕݝ��<��șܜ,��jN4Zb��-@��F&�Z�8��E�]m`�.Y���(&�m�ͷ�k8S�m<�Ǜ���A��^{�yt6ȃa��hF,�7�5�w�J1vïa�ô���U��8c�/c�ݾ��9���C�|0�vU���ܨx��ԧ3k���jz[� ���t.ˏ*c��vؿ[NmM6��C�������:0<Y���bO��T��-`�N�q����&��qk;	%�87Z�W���׋�N����.�I��7��e<�;o[\�͕�8�ج���(���s��4ɚ{�iy� �3�e`fz'^U�K��Z��˓���r�Ժ�:�<b��	����>��)h���'Y!-�J�o&���1s�|�Čϣ��~�>�(��j��S��]�{˹�cHJ��Y��8DB����৹U4��4>�u�رHem��ʉ#n���E�d��η��;`=h!�l��;�|�^{$8/^�gU�z�k묏e�.����:��۽%�������'t�v;�t��1�z�I᧺T �Cv�N�λ`23r*��f�%�����W@�E����lv�����(J'L��b�|;�֨`�p��Ͱ2:��8��LX9B[��r�\jJ^��{00�F���އ7&>۫I���@���63|��"�+�p3S���T�椝�ٗ[-^㭩��0�kEgZho �0��������ݷ�Y�Vis.ҽb�}�юܳ�M��Ǎ
WLfE�:�Knq`+X2 
��;WJ�"�a@͌}�n������K�����8jn��Mr����������ֽ�S��V�2�h��1F��/ ,�ZR$(���gw����ݢ����s޽�OА�WH]���T^>��ʴH�(��~e)B�N��'�6`Ž~צcʻ�|(��,m"���`]O{tCyx�Yb�P�N<�����ɠ�^U ��I��"�R��Ú�[���,l[���ۆ�I}tF\V��ֵ�t7UL{n���þ����ݥ�_L��]2�"t'9c�}W��X��aB��f�v�WU�!�m�N	ݢ�[@mbS��w��+*�c��j,�s)�;�y�q���t+t?tvm�V�mQ,7�;�^�ͮ{5hֵ ��{
v������cBҶ"SN蹢�*z[���':�A1��SkD���e�C*5I�V�@,v�%xf��7q&�����:4/y���-�_P�Ǖ4��(@o�۩�v`���n���Ejl����gu9�v�η#O�/9ݬ�WhF��jk�]������W��Ù���lp�z��q��3YW���h��̤X��5�{t(_f��f�˶��[���4�w�N��<cq
���KQ�]8i� �t�
	�gT��*���d&�fQ�����4ta����}��n������**��$WU(n7kc(�;��^�k]^���/�&�Z.t"�B��3�rsnou3"��b����0�C;.�+ӇS���E-XX3`і�Y���w1�op�/rSue�WX��N���̑ݹO'C0�X��e�S[��%٤��u�ɝ�YA��
-S1aT%��iK��?|oU�?|FIvX�(^��(��d��h�5�(�tq����3�O��2��ڹӄ��`#l�n�T�p�h붱�WqV��ʕk�c�wr�K��,�"�+*�Y��^��[�mCY��l�C�ݹ��S�J4��ݓ��j�7ww����:4�,�-MS�wq�Z�%I�W����٭�o��7=�׭E��wr3P�X�;Az��:um��wZ�6�z�< ��\�ʬgP�j�;�1 ��s܇,��x���_	m��i�J�\;q��zX��W|�Xo���h
���f��cy����ţ��Vc=�ص��S�o�f�*ea���ܡ��Y$n�,��˸{!c�&��3$*�֎�0�4��ZB�\n�kl���+O!Z�s1Ў���N�Δ�\�%�M'3����9rC�43�m�)ssJp:��p2e�����,L*���`+oE���6�,њ�aT�ES�E��7rAZ�Ⱥ�]�5�	��n]"c�`�Ц�%�x�d��FН���V\I��v�KU�Z��X�K}Sֲ�L��3��r5�u�Xqe,ǹJg�K���
�t��׎�]�v�U�o_f��n���G�5����}��<pl��
�I��R���i��%x)^�qh;֖c�"Y��&vp�`�M�b<;{2��0��e��W=7�S��S2�.�>8 ���hܮ7�oei��WP�%sz���F�0\�P@�'�B������<zoK����`Z,���3W+��J�0ۻ��v�M֧W�d��ܹS�se���;��P�v�lw�K�X6W��U�N�9oa9iy
޶�SCq��۱�XŌ��խ��㾧�e�~+�����3�zR�(k�Ρ��Ra��9*�(���%!�fs�n��u��z��q�=�{2�:ÌW �Lgbʆƣ���.�g`��Ǳ�3��b�	�=қ�*f�=]¦c�˦�&��PW#�C8k�;�k�1�"��H͸,��Rt�Ñ�T)�"l]�ڝ��Y6"�|�\�����ˬ��\��N�Xt��m�^9�����)$z�X9:���t��]pv��3��з5��n�s�
r�Wb��S���͜�=��͐6��3MZ[�9�I�l�w��巉�f�\���f�)A���n�@�v��UXif3���gRd4�Wo�uٕ�r>�;�eJu:�#�������;`=�h�g{P�1>��5��m��;���Kp�d%��(Pq��8�Z�˚�����B�wR��{�n��h�0R�^�h��y�&�{�@�S��H��9�ܓ�d�S
��y��=Eݻ�ӱ��w�5��=�dLE�>�V�sz0�[��'4���P�w���A�9���O�)�UZy�o�L�j�����e��pU��,ٹl���,�R�C�Y�z���a��EI��a�Z�r)��!ÝY���<�aTѰ���;q�%�\�B!�I��n<�4G@�����G���H���J���9�S9����{)7f�i�c�$����3Ҹ��"��oF���i��P��E�+J;(Z��OD|�Ek:�ْY�Q�zÁ�pW(=��2a�z�;9]9Z�#v$����&u��@�p��؀j�4.y���;�ϸM��l{!ǔ;o��` <�]^S�����-3�����J�v%��&A����e%k$nT�6��#V�t��Z8��Y��뱵&���ulu�2����\��f�>�.�I/IΦ�iF�Z�`����˼sNs���i�Q�_̢��h��ܘ'5��ػ�t�&�eVWn����v[�^N�8SUg$�Ԋܬ�����0Su��0Si��a�h�:��%���PMKm�n���{-�R�5&��5�݋ƛm���~"���R�}b���S�v���u�+�p�1����~HO�M�(h�>��>��)�OS�"iԾ���R�@|��'�/���K�	�>��=|`��<����܏̦��>=g��/ԝ���5�x���z~����/����;�A侣�*���PT�~��߷Ҋ
 {��Sy��>A?���'�P�|���/�~����was����S�yU.}uPʖe�DTb�E��o�!Cf�Whn�!I��f�ު�7�ވX�g�V`ͽ�9-[��^�s	�oC����n5���3��ì��FI�LI�]M�6�itp��L���w:�ⴱc�;��8�W�l�Wپ芘b������n�e��5�N�</�;�*�4}wb\�ag7U��U�Q���ܡ�S�����d�qK�u������^AC#�ot� �jJSz�)n���R������Nc·iS&sH����ⶨ��yc%H%�j�΂�{��q%K���TM�8�2Qҝ���Ymgl�g?<��|���;�R�Ds=2m��zJ�̳v�+=�E<n���qpҹ�H鍕��S�|��pm���-V�Ord=V[˔�o��p<����(��V��w�i�Ŵ:ݺxKu۝�n5C�>�BD���ۀl�J�X�K�hu΅T9̤1��^���n&2�#��TPI2�Q�|��f�9B�[�OT{����MB�b�jn����\:�Ƕ�
ie�=ݚn6�b`��W+&�V�'O-7�3OVjn�r�i�R�9:��r,/6�Dw=c�C���y�V��0,�q9M�����m匤)���dsX��}�c`�ا��9����j�ZCR6���������ڹ?u)�5��	�o�H�z+���pI��&�av��(E4o9yYl�$�t�e<��m�nY���^xV��.##t%+�*�0��D�)�QwA
��l��޶�!���sLe���C��*����Q��T���v���貆�N�w������az;J���"�h���۹^�qJT��<�Gv�30m�F�Lנ��[{��3b�sŷC�x�u��`�W`}�O`��E�.�P�A��`c	��!%��:��L0��D�]YG�0�t��c�"0\�6�j-��A�~�mp�El8�ǋh&�+L�Ⱥܼ�F�:[@�7�b%`�Ù)Q�t�x&DQ��&)�8:�k�[w��2&����2^��g;�"��N�2�U���@�)c� �6�hR'(�+}�7ge'�;�:��urdӇpbh]�]P�S�*.��+3{��(?$]`Ƀ�W}�)�y���D���1���F$'8d[\�p��7�8�M;i��Od�ö��L��E��X��Q\�'K�[%�R��v�o�;{E���"e���&��:;4�Ug�}$��r���͍�V�4Nz3�yҗ�%���r�����28���VF�ׅ]dPv��ٌ�[�bzX�%\J�K�}^9�yՏfn���ǘv�ʚ�VHLU7,�k(0����Z%(�~��������jv��!�Gu���X@r�	�ڲh1eLvF��[1�B%n�x�!ם��w�ќA��.�?��]m��ɍ��Q�wAĝݸ�H۹ �y���ږ
�9o�B����3
��JdP�E)u8�B��q��G�q����WEE�9��h}Xw/�*�搸cx�R;�&��=�h���hrij��M��d��Qd��F%P��K����z:���t�"�M�S�8XP�&6j�����\ӈ`�X+@�2n;J���L�5�$撽l_I]OW�GsG�U36k�ɗ�G�\:&�H�h0�n��1��VH�ڙ�c�FG�Z�F'}s,��zɵ���/X���ІгHYKp� ��VMĂ�;O5KOmw B��Ð�lR&�� aOwz�-�}�\���
Z���g+�\����5(ģCv�I��@��kY���-��|&:ҡ"~��9vwY̓y��cbܵ��2��@�sz���vM�)���Q�>��4�1��J�����vn�V����R���8���Q���g�.���^�w3#����ZG�!&�:�5��Ս����(]J>W���������t��d�q�X
��]�����}Nܶ�������{Π�%�`aa z:�_�q�,J�3�{�����<&�Rr�+[+Z{¥Ÿ�#V��L��6(�EU%hݘݫӔ\[�fɪ��vh(߳bA��X�dg�!����k�ѫzĝ8����H$��˅�3�]�H2��&7��n�3.s���T(15��p��1I�`��o��Y+m��;^V���Qc��h7���d�N��� 7Q��dAR��޻�K]�m�{�-3���<����d�������k ���z'Һ݌���a)+X��t�ƵDب�qh��f����(lP��gT����cBi�b�+�A�F�c/eNT��q٠,���6��Y�A��$Z��$�\hQ��s{��S��2�c���,��d�m'l&���;���R��H1+��f��8�P�����ۖ487o��F¢�����v�uv�4e��ΛtoC��{����&�=q�Ê�7��cs]�ݩ�˂�'	��u���gg>Kl���`1��X��Д\˭���f�1_e��P){�nM�4�ܩ�j�>�Uنł77���/8��B2�����q�NaI	�r�5fvJu}M��l%��C5<D�M����L��nǣP����̀�*���8�(��]5��z�W�f�q��w���#��AT{m�����f3��ǯm=��ؽ�k&+t�wn�+=��s��L>�Ag��4�h�+z�z��X^J،�<i�޷�oS]f��u<��ġ�������fN-�����j���.��<��:y���yWS;x�8b:x0话ߚwB��̗��9y�14y�4��UcP�����1����WG��1��1 �K���nq��m�!������^�Y��qd�
���ruR.�k�]�}.�J���E'x�%���8W}�"묪�{��R֕3������Y<�j��>�|�/#���g����t�����7���"v�fP���dz\]��*D��M.C=���y�@��]Z��6\u�����+1:\o,�S	��y����tw]ٲv��k��Kz!I�R���tיe15OK�L���⮉���iy�0���{��B���yy�b�H�ug.�R�^�75�X뉋yxLP.�����.{R�V��w!�IΗ��T�Ucg^��u�j�bۆ��z*jE;�C�|D�;6�+)nWn����o���H��M���ܷ������U
S��I:k�<�t�d�:.8�b�C,)��/��Zs�=�i����=5�6��#O�*0-�y�DTm�u["ʅ�<V퇌9ȫ�/3q����8rz��:�wP�4���l˼�1��"IH�k8kq�n��E���]��̣����q�Y�0�ga�3�<2�q�����d�-9k6��t�����d��˦�\F�R�3Z�Y����4b�]��9L���{=� �\�2�^:-(�;�{��h�^�w�ct7X��&�uv��M���3c=��˕#Ҭ�,���{.��|���,�A�gEd�c�ډ�/�ܧx�ݭ�5�.�L��ow,`�O-�R��k��;މ�z���
H�nN���-F�R����UHjo1EB�2=�_^����-GR�is��-�S���6U��26'8�jϽ�B�3�6�Ia��i�����5���{q�v�<�eih�9�T¶���F�(c�fnesw�㷶0��A]ۛs���\ʋ�^��U&-���K6)e�zH�����\���ҿ,�m]f�ǢA����'n�k��q�\s�a�3OQ�-3Д4�s�L�q\ԝ0��5��x���$|6�/�X�׊�\©��z��J	<�����Up�*��������A;��5��]���Y֔��vZ��m���4�J.�o�fU����j��O��RĈ�2���!6qTyVZ�q�m���o5��b��c9z�pW.���ĩ��c�%�)WQu�#�j���J������G�]z�|Y��Re��u4n.,��Jk\�q�;�tgr�C:�U"�����t�r�K춖^�����iSj��N�&�N�!��7g{W)b:��d�7�nf��Cջu��m�'�5!����^X�c�
3��
�#�Ol��犫��k�]R����.ŰV�Y��X>1@���C1֛�"�	[.�i�j�A��B�X�Wc5uc������i��e:S�0��c����ەW_���ӳ��M��A1�Aѡ${�
�����qLn�z���W.�S],��FM�t.��e�#jh����]#��ZLp��2�_;�K)��'�S|�Ov75r�g�&ʬݽ۠�[��D(�������m޺���5�%���v�^ֶ�{:]:�4ڐ�@���˾�wڧ�h˱KE�v:��>\%>��EN��Οcd��/!��T�:��mj����Q��n�oG1�#+NP��h�6�В̐WY����YQ�D;�.
�7Π�n���̏���w�.�m�X�6\�ɩ���篰�*���r�2��J�v��e]'�4�#Lz*8�X7;Z�wo��`^���WN��g�;�nZ���Z�ɥ�>Kլ㙦.sr�=
,`�䁙(Z�����ݠ!���-à�M�e�>0�est��ೢ�w�5s0�S]vWo��[au�j��ګ���b��%��;�n&�E���;B���q>��W�����E�������֘��mb����L���I�����㺚5��ۏj�v����6� �rnVBQ�6���!��F�*\PW�;���1xT�S*h��2H�ʌ�Z� l�*�������WQ�"ټ)$:@��&�:
Sa\�f���!,�@��T�	���h�(=cz��+ӣ�+�ˡw2�D!��q�һ�R݌�^�r����@u{d��ִuMt2.i���T��ﻪc�ꗱ��j���H�JF�����۹P[۪���o2c�z�&�Ȃe��bq+*�m�#��8�����;4�ˆܻb��q��V�q"c�:�%�&ԬS�s'3�Q)q��*;�@]o'nM��EJ�$UØ6l;.�UcZZ�u灌K�]�`Eu3h6@�*J�uW��=�1�/l\���X&��q���T��1Y�U�Ϲ`�y'[�dgg<@��ٹhԦ��/Fk�[o	84�v�$�\f�c[xs0�;{p��N:�[��#�}+�[5��;�����4'p�ek(Z��6��9Ʊt5}D�OV1̻|��t�9AQ"5�ŧ�m�ǅ����Jm�P���K��w�Q���,9�E�sh<�dط��X�ܺ]��|�8L����4��VXՓ�6C��U�%��3�Hv2�P�v�2�|	�ł�-j��B{���Y����%�qL�*R���٥Y`�k3�ou�l=I�	��9�Fh�6�3,L�ۏtd�۱����q�T~Zh�N�`<�4���V���,9�ι�hm&X�`@Et�{Y�n�z樇7Zۃ8��|2����4�8��w�f��X�BFK0�����@�td��7.:ڶR�	�UNF��h[Lj����O
�x�N��w���0!�;S:�A�B���YQ�f������֌�ս����@����=ytZ�c�V�h�F�6G`n��s;��9���K�:T���-��
ƅ�eN���(�@4��4m7�f]�,2n�D��tu�͡�އoo��mh�CM-5R�u`e%�����R���(�ds6�M��#G2���de[��c2@7cݽb�n-�rPUw�d:v�����	d٫`6��1��጗9*���]���wm��I���&]T��k�!c����;�1nS,�e������ 
�VT�gv���eu'\���
U�]��\������qE��"=���S���=�:͛O�!�aZ�^`67����A�_��[�������I�f'���C^�6v�``��I�s7h��nƄ7D���:uf���Yp�wx��T��/���Im�{7_v��+" 8Wa�\}E�X�"q9�����R
�^�[��c��Q%�u��"���dn	��Ry��Z�.j�������*]�F���n��ud�b�:ܗ6�r�4���&��Ȼ�M���MF�t�jZ:���:��Bى����QD���L�^�/�&���.	K�<�U1f���{�t�X��t�����0v���q�F&L�,� ���������.�Ppy��)��`�.�(�-���c�uW#�F���ge:EsaX1\Ŝ(|=(���Uڏ�Y�K����&vқ�;un��û�6��2]��a"4:TmA��G[x �ه�^��/z��axVn�M�f��;�<&�C`�X����d�YN
#��9�MW��+y3�Dt��Uf 綱]��!t̽-�����=N�ɰ�{J�P�{�6�ʛ\���S[��{�u��b5A[ڛtz$�A� pT%�ʭk#!H[���.-WQ�5d��tΓ7�d�z,����'����Λ��ǺnnJ,h'���ע�S7�9��:>�gF�-{�U�Y�<E�"��NSq�3#�2���u^gl��MU���)!,�tf�9kX�O�a���ڥ�,eT�2�L2Js8�J�c��5Y��Őn%Z^5:�ar��vj�rΌ�OV��R�%eH9�po-��IU"u\�я{��f۱%�ObA�YWf�Jᕤ����n'�#U���6���x;�˗�Yq�4��ac��	���}|��}������G� 
����?����������@���G?��?���������g����}��o���>�o�����}>�O��~��� ������v�.y��򅖂��RJ�i"
A�R0�g̖W�M�p�Y�$ʀ�,����� RK$FF9%6���F�h�mq|�(�"P���(�1�F�b�!"
�BIp�<�i�	��eJ�ʯ4wt�u��w�e�\N�U'6��{*�4�Q�f��
j;vr����*����Q� ޣ��h�b^lC�VxS{�aMK9rmNկ�Y9)8G���+*v�L폪Qr����o�NT�Ae�|���r�Tn��Ǯ����Y!b����y����Z�"��(L�v�+�nA��L3Z��ؙM�ܶHɎ�,*6�.;����-꺾v���$��$�K����9�Sd-,�E�a���]6`��g"���S��/�Uٖh�|k���ƈ���8^e{�*^Q;{�+�I�d��#�U�wP�W��1��["�h�p�K�D3�
������$�F�HĦ��V���ȟ�,!gw�/�ջ?@��)�b�i`ڪa�mQq�}���aq���#Z&
�l�t�<�R5}�QS���3K�F�W�k"�ã��{T��<k%N�t�4��/�ow8T��<&������4o;r���B�Y����2p�m��K$������n본��&�����uJ�r���F��]D,nf9�:�n��I32q�vMnbB�7Wp��	C+�ԚϥM�:�6�-n����2�f�g%��� ��4It�U�������e����O�#R���[M]0Q	�[{B��La�xn��s�� Rj�aF
r"a	�!� �P���L6�,Ϛ!�a������J�����0�c%�1�(��6K)��!ơ
8"hB�`EҒɌ�9A Iqg�*$�)#0��Y�����ȗ�$ 0D $F5RI��L���"�a���e3��a,4Sf ba�2[0E1��D�e(ZȄE$R@���C�9
,�DÅS,6`��ē*6\�3F���a�(���#�A$�8�\�"���6+X��q�D�S���TLZƛ�h�llDm��b�ţF���&�j��6�՛[`�
c2�Q�����9ֳ�t㱩��4�mDkiM���5�l����T�آ�(����#�cMm��Z*��ڢ"ֆmh�����Z�b֩5Q�Z�7lM�AE�m6բ݃s�*�`ƭ��*�jѵ�1����DGZ���cc]آ.����:��kX�����։�F�jv[m ӫmE8���m�h�V֢��b(�M�V�&�֦)�3&؂#����ڶ�Z�kQ�Q����mYѭ�Z�4�1��h5D[h4�l���":'�٫lE��l*���Ղ	�����s����tV�����m���kU�j֍�V�QŬ5MAl[��ب���6mZ-X6�Vƍ�bӪ� �h�m���n�h#lE��1DD�ڨ�٣Q5Ej؈"�����lmV����֨�X*��������Ɯ�E2�R�%&#a��m��K
���I�_y���v���Q�Wr�׺��� <�H]x09˩M�q��� �2D�,�6��N����x�[��m��DS��`����=(��b��#�ȤDڵv��il]z�v�R1d��:fI�R�����3�D�O�U����z��<�?d6���(</�F���y�4�kӌ�'[����n�Ϣ�+�WGnC}�ιW=�h�������債�y�a�˟A��"�Ca��h�2�dN�w6�o�6_!Kt�z�Ѳ�;�"?.}
��?�l���=m�I��I��4��]ir�P�D�眮$ڿ�02v*m@�W�8TuO�}��2p�׉��������ګ���?v�I���;��o3�1c��j�C��8])5�aki7�k6�A|.�{ʯ������q�!?+�c�N�^\��ij:9�"����t���s>����j]yؕ��_+y0 ����C���[�w�_&`���0�]V����^|集�,����T<�;��*0.j�Z'Jl�J�jz�U��
H�^q�2���[���џ�������݋�B�-�h`�*!��W�Gz��r��LP�8�Ӹh��!<���=�i
#jk�ߝ�J�~S�5z�Xuն�G�Fh��U�>�*J��K�Й�̸藼�zgF.U�����Zg䐪�G fe�wof�� �靧{��b��)D��w��B��O_/�����������ض_ݽ���츮7���)���q�n���BȗK>�]FF��`ޞ��ca�c��|_1I�K�]��.pa�qP����[��C���/��4S��+>����i�4���\��0-4�gE�Ϙ�ӽf�,}��og�!�c��nmwq1�2���8��|A�' '��0ꡜ���q̄_B�׹W��U��p8U�Q��dЌ���tx�"�I�_���5���W%��2��옍!��ج��px�#y\J��n"��,�����:�mkޅ��wv}��D����j:�ѣ�?O�qH#Ԧ��䅅悗KM�P�*o�_\>?wlF�z�'puß�GFT�1w)Y��SK�"�=������	[�؉w϶U���\7�xA��{�-Z�W����Wc�W�\\�I7%���ה�H�`�:F]`��y��v{�:�>c�ء�u��{��V�Pר�1ï`��ݩ�wպA=�?9�1pe	�k�m̖��Te9z�Z@��"�}��.��ٜ�n�k��^��ٻ�n�N���؟G�gӫ�B=���z��˜�w��q��w#4�#q���Е�����B�R[�m�uq�z��(�|M��uPz�F��Q5����:���4�*�\+�j��|�s���7�)i���խ=&��8��pw�
��D8N�wPv"���3�m�h�2��ݷ�x���j��6�:L�}1
D�_OР�q΁�*��*��%���d���K�}�=���{�1�ÈȐ���)�J�z������(�q����S=�	B�d���5���8i�l�;�U����,�CX��fřQ=qƅ��ǩ�pn>΋�s�@�\���V��������H`�w;_������yW��5���}��4��@̽׏���"���=���_o$ln��u|7n�cy[[�QYB���Vk�Y.��
g`����*�ə>��>�ܔ �Y����۷�m�ѹoR�T��`s7�`���zv^������R=�̊ga��`U��5G5��:��c�.�=��cc��5%8d*��M�����T�L�-ƛ���0��������U8�=@����>�އ���i�$�'�ή�!�������k�zMA3'd�G�N���[�������Փ��R�LDs3��l�6�k��@��B	9��f�*�Z��	���Jm�Q�$G��b`у/^7d�mǛƃly��]%��ŅٷɰJ�f�gGC�A��cհdm��۞2zO�-��XF	�|�����O;��=qZ����Lh��5�p���V�����R+9`�ǛE�.7����������5�a�Hɩ��&9�I�UcaO!J�h�<�v��U�1>}�u��<�k&��W0R����X�,�wc/+��+����g0�&,���εMdY��_���!A��[7�;SO�إB�v�p�s�U������/~߶x���F�ol:A�V�W3pn�]k{�r��}Ep��eh)�D���بVF������a�]O]+xY�c]T&l��#�4N���k�c;m@�Ө�"�x�eA�!cI9�KQ85��\is{SV�4	wwm)*4y�^�X�@�
�<9l*l�;E"��z�8�٪��Zj2�*��������oތ������n;�(J�s ����!�]�aWG��^�AD��IQxnO���A�t+��f�Ԡ}��C�c�����ø�y�W�z�y����5�u¬�����(����)�w�8����O�m]�tW�bϜ7����}
�u����dw	��C;v����l�M�0�蜝{z#w�W��3F��'��6اOd6�ɫ~$��t�O+����Ȋ����7�z����6�7C���I�繑�l�\��޴�1��Q\��7"	[����9��x�8fM�������i�Ӳ�v��::�6G�)�$\��p�����&�s�:g`n3��%K��q�Q%��O^��Q*��`�%y����`|5��ޓ�N1XaW���T�gv.�I5���X���T�a��w�}db"-:>����$؇�F�?��1M��<��s���U��t��#�!ۘ����[:��n���a�B��{�^}�C\0jb��!ǝnm�U����}�5lSb��Y��v���×JlĬǕ��r��HҦ��
�vh4����C�{�ߖ��1��<��c_o�𷼫���s;��J��fN}0�*Ĳj�)fu#�+�����@���S�>�ovU�� ��kvM��	c���{�m��5���@ X���R��f�]�y�=-�Y��_Z�;Kge;�t"՘�9;P���">p���J�^vGu��y��w,R�WZ[�i��+S��v*(�qy�(s_�B�����n��T8[��Ji��|�;��n��v�%�*���kυv0Q7�Ďn݃����3�km��b���w�Owx���;<Q�^�~|�g���f ��w+MF���
U�h{	*��p.16��
�4&0�Z����df`y���1�Q��E��D��ˋ���FP� �gg\w=?�6c����'�s��>�K8�OC���3dЌ�ݯp8x�ow�3)��f��g��2_a���Sc��tVB�j�����@�S�v�-��s�`��!Ve	,�Tm��Ƥ�V��V�rSEx�bVPD�[�-S�;K#&;W�vk#xoO.�od*���.���Ѿ=�t���y��w���,�l���^3�iI��Z�}Eu>+�4�/8���[=�~Y�Vu:9�
���	������>����\�W���z�q�6#I��r6��x0l�$�WF�E.��R7�CK4�-6aG@�<5���t@��MP���͍q��GH�K/yotӱ��7�yc	+}��l���j����얻y.���,M��4����`p�7�F��Qv��x=�G�r�n�t����iW���FC�Ĭf�&�峵1�S��L��*�=���]������}ס���xƴ���s�U
���UL%P#� ����\*[�ݫ���+�I��s��}z���E�����8���1����Yu��mGj.�}�w�\�<[TS�P�E+�G�0�8�sx�.j�k]�:\��nsꞨI�I1�y�pͷJ��s�t���ܬ�BH)GrA!��J�Sx���ӛ�ʬ���7ǭ �]�g�V�y6�:<�`�͸��H��v�ٔ)ۃw-���Mg[����Wv�LcN*)",�X�U*aRҔK�c&��k�	��sp@�fQ!i�J�1���fbo2Z�1�HIzSM����~��g2�o?Jh���qmï�sL�/��ge8��{��˭%��N���r#�dgH���8���\$�>����G&!q�O��MC��UD��|z��3S���D��b��?ow@����輪Uǒ��m�Έ]����N��OW��d=��߆����˿�����KJ)��{��'��ʾ �3�z�}�w"��Ȏ��ȧ�ѵ��3J���b��lU��Bq�[���|;��݈?+��L���6C���}���j�Znh�W�3c�c0{� �}��+���Iw-^�Va�[5�wV��tbK��p1�ji�)+�툗���2��[=V���7��<w�+�8�q�b�*�Uֵ�����3���EEv���3���5�/磧��[��#�W�":8�p�z��U��o���V��x���qϗVl��[���q����r�������oh%<�tX�ĭG�E��xs-���J�AT������l��`����ˌ6��כe\����wf� �c���z����R�2R�/Z�y�
gY�L�ik~�Q�m��1��(�][��<���6Z��&u!W�{�}���>Ӎc�5y�m�^G�Y�v9�N�jq�B޽�6Vr�V��o;!���ݘK�{�V�d��_*���	X�}q�^=�Ӎ� L��!v�V�|u�a�_0�gsyԋY\J�{P�XJ�fh�SO�LEG)�Ob��A�Q�o���-����*�|;�<|M{�l� -�{`��k+��"������V�L�-Ӊ�W��<��ؑ���[�c4��F�#i�8�2GL��9��EY:�0{Z.73Oi���ϟE�tT#��$����c� "� {�_�i��21�il��|���K�5���N���FD>�XP�ڮF�F��W[}�u��m���1%�o�*��[YAW�q/���>�fJ͌�h�'��R��N�]�l_X1����g�ё�xO��q2gO�?���=�U/��vݐv�6b1�&:�<Kp0C9��)+;���*�t�-YW��V��sx��e��ђ{a����/��w8`Ǽ���e��v!Kc��3���O��7E�krda��1�� ���u��{�z������j�R�s7�<j�w�h2N0����ґ�6���7��6\=����t^�w��Ϻ�;K�ػ Μ�Y=]̽L)L��d�W�*1�F��C��kWE�׉��ockk�OWwB�L�!�vCU9̿@�p��5�g���'��)��x�m�:��*�y��:���]3>)�ȵawB�<�v���uL�G���/2Y؟��=�0��5"!=���y0���U�@J�,�[��bn� 8=uG�[l�����_ݩu�����8�5֨1�\u�siLw��8��}�9��3��htvH�^;`��}�^��?|閡<�z]��OTB��(��������#���%3����KV>���5Ϩ��~hø��m��Gu'���>�zڒ��v�{e料|){�����Cۇ��ꙇʵ��VO����C��������������'ǟ����}��y�o��1���<osV�T{噿a�iF��f��b�2�j\�������5�G�|���u��9-�a=%�)����
��,I����u>A�VB��8Z�ǀ�&�ݴ��026�9r��1�~t���������Q�O&j��bF.�h;���4��:�h���<vhv����|%c�6x"7��24i�뷲T�mZ#>�5���w;�lb��³�R՗L��\�f�i�\���Se��]s]Սa��ڄWn�+�Y�J����pKsX�����j^�0֨�M�vm)��:�P��I4���͖e�W0���/v��ʃd=��L��&�Ņ.����+�h;{�J��x{�{z�Y�QA�s=�{Z�h��j�U�+N�ס:h�:�Nf��N|��[�7��۵&�N���\�=2�F�칝ك�,s���[�#�*Yzl�U����\��0�]j=W2�>u{i���Y�++��V�vv���Y�2s�X�o�� �O^��S"���G+'(��L��ޙ��K�El7�NOkۛ�U�#;))��8ɾ�Ź���䎙-��m�!��)�v�Y{�@3�g9J��;R5Y���Q�a�
��H��0k�A�
I�t�/��b�=�����t����oݾ����,�$�
),P��#��J��ﳵXٳ:]3���Vc;�m�{��D	/�7p'X��XB��{UP)ڤ�=
���:��u�����E�:u���*CE��?�]�j#ݽ�����m��/<;Aa�aSh˸�:�=N�]9F���5I3���Z���
�W&4�"��D���\YI�����w6��y���U��*��X�k3{�_���5N�����]�[!=����ɺ���Z&oT�{��C��J�,۔�:M�]�`�ǯ���Yrn�Z �u��W+�-c�Mݩ��s����fTWL�z��&����b-uh��6H��8�-���WC�;��˺բv㳴�As��4j�u�'kMZ�`�[С�6B/��g)�VL�n�4�i̲��j�j*�v0���'j�^��*�/��u�Ѯ7�sl�|�=�����ʱ�cI���æ�er6ѷ��\ә�Z���i�g�E6K��u(����M%.���z�]��u!����E�Y�0����c4+͞��m{���w7lk�o1@ܫw3T��M�w��9��<p>��Yu,Ô�l2��,�)7�v�>V�;s5S����LC2rmBKZ��V��2\4�t��9V�a�V��Ƕ2�L���s��́
rmՅ�g�r�Yʪ�zM^����>$Ci�T�����a�#�N�H-\�GN�ɻ�ԑnX��lC;.��I���1�$�2���|��
��V9	hI�de�Y����<�&�Cg����CDʽ������[������E�*�f-b���tu�����[kQ�ص������]b��(���ڪq�o��IZ"(��)ֵ��m^����bb��uLUEq��ŵFՈ��hѨ(�&H֘�mAV��+�ִX�UkU4[EE51ME�:�F��*�������Ѥ��v9�g1�jv֌�=���P��]�:-�kTULF�m�Y����ƍE�W�bz1�b��T�L�5Q��ؚ��*(��M5�[a��:5gX�hɶ"�lkQS�:�uES���6�u�[4lcY��*���$�:6�������G��Z��C��+1UUۻ���Y���]��nڣ�MV�Um����&��5G�z��잮j�Z����"�^���t�)ъ(�k�UU��:"+գ�[:���ևWj5QQE]jۢ���T��;i��(�"�j��"-��Md�uhű���X����]Q�Pv5z��j���'�=A��繂=��(*�*�۱mQ5uc%kmA�4bകG[[�Wu��O�Ѷ~=b;>����Cwu�z���맛�M��h�lk@F�s�bǨ�<	�&=~^���?}�F��6���I�[�P`͛�x��NU�����p]�u�Sʺe�-`ġ��� ����u-$��51�w�8��MB��JwWqB�{K�]F�K	��wk;O����H�8�v��n7�^x�����k�ǨcJd4�`VzؿV�����q� C�F��{ǥ���4�w3Ez�KE]/3P]�E��CS����P}X;��OVj�k�>�
��F�������-�*zr�� �թ*f�{ԃ,���L�Q�y�=���w��n���OY�����]�hqm��"���j��W;��Jla�R62��s/���љ�����r3I�(�Fc�M<�o�������	`j�O݊lEmx��b6b�����OW�2���≉d�#��T��#�񹩝>z���`(�����c�'ՙ쮖ͬ�w���þ�����-���?D��>7��T	e��I��:皟"��t��Z�����+N���������Oy�`d�0�GuI���۹���)b�Û�LYp�q�Y�*^�t��Tr��w�r�F�Ѓ��DsmLpm��iO�T�I�M��Z~AGy�y�
Km<����kƯ��u�ea��o�q�a�_@~�l>�Ϭ�G ���c��M7_j�k.����<}���R��fU������b��Kr�I�{�,�jaa��Ci��;qШћ�ݷ�6M+׫3���ط���2��{sq:1tyH�'����٣`�]��y{�<�\����^a|����s��b"��!�Y�8����V(>o[}1Ǡ�w�|ǔ���dLB�q��6��>�ϨV��-��GQ��8�����2��|���E>��UBr��1�����_Ԙȡ(t�O|y����ն1~f�M�~-�n�o+��e0�/���Z䷪=7����[azu�Md�>߲m��FZ�z䞾���s&���xf���4{e|���i�x��@;@��j/����0�S��ʵQ5{|�{ݔ>+��B L�>oBif:�N���wHns�� ����L3�����ws�l��ck� �edM�Gڟ�\	���"]���m��x���p�m�9�绣Lѻ]��n���3-�����v��8�c C}��v�~kO^/6��i�����L�#G����ʅ��cM㘎�^�F�ﲯR^ō�F��8)�d���(5y#8�C6q�dgO*Hc�2`�(�b�क�l����>�*���x�{~By����Z��'�-@�RF���c��<�/P��fp��m�B0ܭ<�y��d���x Gܜg��ˣ[�������2�D�'W�F�+�I�5+�i�p釧�ƪu�"A�ZʣbÊ�l�BjV�[M�)��g�Ί���]F��Ln�����Us�Z��+�f4�<����ht����ѳ�+oOD;����{���jU�Zz+���*S�]87�M��i�7kW'�]/�J�}̮�r,�3{;�,p�h�x��ْt���p�\3<_0T����tl�]Lqv�>�b4�-^c�'�1)դhZ�T��[{�ͼ�h���M�6WV�A��b�t�zA|k�:Añ�ղ���:}2���Te�����N2<&C�����w{w��u�upf˳e<0��6�c2Ai���'T&�}YP�7����,4��;�K��w\+׬1LK���9���E�m�� ��
�����Q���T"��>S]]Pɹ��-��q~�3�U�)dw<��I�Ґ��$���r|��X:noWo{��~Kn���=��2�����^5�/�q�N���*�
:y�~���G��i�r�� ve����k���+v�g��Qq����q�{��B՘��:�_�sߒ�\kU>�a@�	�n�dڗ8�{4�U���s��DÁ�� ��i���2��,5��*�6���S6��=�}���5�]{���i?�\�f���@gRdK�p0C���~��fI�t{����Qo���Y�NE˩�=��{��۶�f8虗i �c]�ʚ�L~1 ���<����V˘|���0#����z8�6���~���g���W,����;�;3 *If�dK����>�u�9+
4�m�]+�N�9�����5'��k̓�m5ѭ��L�!Cv�Љ�q9�N&�I��-4�<h᪇���"�N��.�8o������l���I�]3���*���Pi�e�N��U�n%�lg�f|)����M��q��5W��z�+-�Ǉ�򵍝�JI�*Tk��޹W#^in��?��WE3��)öx5n!fM�,��ow�(����e���/sQ�]0��L��A�n,�i��lp�����&�Z��Q+N�+a�1L�:b��ЊbOQ���q�nvp>���`&Fѯ
N�Ifব.�֢́v�j��� t�c��V��������K�0�o_W�n��7!	�{��sK��J�|ݮ�����Յ�RX&�	��}���5�z,cü�Ԝ��	�By���Cz����-�)�{[;�D�W�yx�qU��CtKbu��L��0�?E�������>�����.pa	�h�3�ȣ���v�r�ڳD�T7(��dQt���.�n�e^�iۋ�r��]�Su��eiiՕ7c�mv�L��E�,jc�YM�D�q&��"��_���zo��9��"-�4k݆�-�������u�������!0	�8F������Ӵ.�Te�X�Ψ�+����y�	G��4�L|U
���9:/rڤ�hk[���ԃ^;�,�����÷Z��)�vk��I�����R}�K��,T�����S��{[�y�Ɂge�GC���&-fZ����Ң���u6�u-Y����gkz�SGK��R->�de�}3�,Ē�YǞS�S#z.}�����Xtz�:�ޯK�bْ��L��OJ� �M�DjB�v�0�7���5��췵�ʙ;��d#��5ØO߃��P�=/캙dZ&�}?n;�u����K]�;Jۗ��oSi1���3�k���K�gbLg�`<h�\	ų{����ō�Qr���:�㍜��P;!�I�)��Ǥ� H�v������5�n��Ǟ �OOѴd��>ʃ]K�-(E��qƄ{�&䗿��K	�27k_�߹��$�q2�[?�lEC�{�	��k��n�V�g5�����!�z�x�s��9�n�h�_H��U�B�Iw~�U���W��9�[�.�z*o�
v�g������/�T��Cq��u%Lۆ4 鼞:��j��F��on���}�� aVX3x+�;�(����E�zGb��ߧb�����Jm��=��wyT�u�a�sR*Hd�i/U�ؔgPs�Y���*�-I���08E�6>!�gO���S�4����#��d�'L,��Fi��)Rk���Ʈ{gO"���	0���t�)����Ue�;=޶S����<4u��m���!c3����$�7z�Kb���@ٓuN������������r+B�� �]���k�\���{A:�	�0����R-��eI����6���QR�ɷD�۝1�M:X�ڐ�*�Ԣ�9�=��#�����Ƶ�%ٯ��&А�y��%:N��:[X�R���s�^�p�s��C�%�i�U�a�>o�Ŕo�S1�0�\�KϜ*�a��/Z�O�b����)P�E�7�A
��|��N2Z�V���]���{M�"=t!6��ٽ�j/`�]M�K����~��e�>$�^[���[�qM!PFi�����"�h^���=�V*���<�;=x����o���I��{���d2�Lw=2�s���8�c^C�5��.����xMtޫ�e�h�D�f�����+���ƽ�)��tu=%s�S�~طvm��Cs��ӭ#3��#H�a�=\�<�ӯK�~8�Q�bK�^5�����WX���P_P�n��0��Yz_n�棼3�M�"�k��_'ۆ��v�N�ד�#�p�.TO�.b ��'���8"ͣ���Z���[;@C`����1�5�=��@;�B(4]��f-�S�R3��Y�a���V��"��Þm�l�w�C@.9�&uc�q����@̳LY�O_�~ǐ�~T��?f�k��+|��^h����"����u`�|Qbۂ�����p�j'_Om�9�.�=<�תc.z
U���DM���*W+N}��S�:6�҃��|o���_��[����/=PwE�ݳe;��R���(N�]����� <�6p����s믷�]��L�gW/(�S�,">Ȁ=n؆�șvm�����yǋ�l�w��B1�y�-�{j����2�8]��j�����,��/�}1j\�ԑ�g���U�-�?4��..�bp(j��6?s�­����������Ƞ1��	��a�z�S*H�3��{k��s����#� י�{�v𯷸o�Z"q����a�7���6����΃?�Ƃb���j6-_�)0���8�GubĚ�+#+�ښ�ӥ�Y�G�D�k�:���C5�	;^�7�M� �	�{bS�Hд��/�y�OS���dBӼ�\1l	�;2~0��?<3�~��|�[	�f�]Kw���=?U�'��u��S�i;d�J���׋���O\I�[��1e��-��c�!=B}�sཱྀ,�ϐ�ZHH��w\��9��vf�҆^&�s����E�1��8�H^�՗��<����� C� ��/��'Y3(��I�x�wŴk��&@�yj9r�Մ���[N�|�ٷ=������9�̻uI=�ݖ���֕�l��^u�z�ԤY�u��*��ʊ����`>�cD�?�O���4Bd���Q�(�E~�^j����s.Bvp�XoM(л����k�C1��c*�;���'�u�}���~a��Y�d��'�$���(����a�+d\\��|�޶7GWuÇ2LZL4�w�q�\���oVNfns�­��lx|?���|�+�j;
�!�}�j���ƿ1�Lxkf�H��:~��a(%�Q���1.��v3��v̓L���|��8G���0���2S�L3,�nQa�]�P>�VDEլ���f�Vlpӧz��+SL������w@����̒x3�|O~�o�p_�)u/�eB~_�wBx��7q:�EGV�l��oh��l4�s�&Y��x��i:"��g/��/�P����]�z5�$+~mъ]���W��2z̷Z�4�#ّe�!��@A�܌�HD[*ok��0�S�4�im{����A%i��B=M��b򴍔������[��r�g�>S��b��{N��!1���gw+|���|�cB��U����9R��T�e�b���O�~Jθv���7Θ(�)�8O������魮tW�_60G�cA�0{?L)X��nj���-	�{�m����&�A�{Ά�%ex]���Z���[=w�ƆA>5����!7���Ob�`.ɶ8�{�^8뼻�}ݻ!sre Jue_��M~��x[�]�s�<uxCo��!Ŵ'H>P�'����7Ym'�!�F@�/N�7T7�쇾}i)���C��Ֆg,�>1�l�$�+=�)[Hܤ.�����p��ɾй�:W�*�<��0�r�p��iv�T+�1��X���{��g�T��i|�ۘ���4�z�Z�pu�j�p��n��x�� ���"��t!Ht�}�|��������p�G��Ҍ�N��bY'C�yd�┦���{#2�=�o�A�loV�8�Q��c�Z���~���{��b%Q�P�r):ahԢ�<��C�n���p��\AN6"^*����𧻓L�#!�ki�#[�� �Hƅ����8���,�O�~J uBw����)=[�m�q�m7���5P6�+�}-���n�1)�L�C\�b]F\
#�����g�
}j���K��}��n��@B�Х�-@��x�� B9�Ha���z9\�6��U��cs{�<��ֶa<wT�^����3�ЁQi�¸��p��vB�:
��'�}�_�b"eh�����/��wx�8�"�_���I�����dϧ^�&g��d�,3���7�WV���(������y�G��M�d{�É��+k�.����$@:Kϰ�i�w�X�c>�v�&?V�����������?��Ac��7�{Q��`�c n�0v��$= <M;L�o�L�hDK���ʘ��4y��*C����bv�}����r�9�w3E_I`J�7����s�u�ժ��u�0��~�X�����0a���
+�m-�ЭN�����r���Wt�VRv)j���қ("��J��,UǏ�{F0����ES�7�Zp@J^ �Y7NE����U�[�U۽�f6��'l�e�Ҹ��~�U�~+�GH��H4C@S�@RP֍4�TUT�~>j�n�Y�x��q�/@���kC=X���t��Ⱥs�|�8ڒ�loC�u��=*��9���CZ���5NP|ش���yV�w�-�ä�o��5X�'�fy�5⢭nX�:��yş$�H��2�&�Fi=ʿpQ��z�o�Zğ��d�/Z��?wƧ��R����ww6�qq�׮�|�#sS��P&%�t�K#�J�]�#���9�<�{w�u�U���WT�OY���J�������G��<'I��Juk�S*+��63���rWg5�r��ڽۻ���̲�����!�yٶ�81��.�O�$É�I;�� ��-I�En��5 g�	��%o�"�9lG��O�}G�_m�@�#��Bm��ۗ��EΥ�X��.-׭׺~�uu�am_o(/��)>��;��o��0�`d0Q��G8vvZZw����}�R:W�I��a�<�ެj�<����^�1����:LK�F�0���B�w0B|��Bk|B���u�qO�0%��M�.�)�_��6�a\�/��r��i��5�\A�����=��w������{��w����z���7���������z�3;�}�Ym���z�.��͛��7j[�,�z�a绷Z�G��]�
�罕ij��i�YŉN6p��d�`ݻ#�-�RZ/��y�bi��js���M�Wvo��W�-{���k�g�{���uͺj�[oE[#au��;�;N�ݒB!�Y+C�l������������4�Lɴ<ç�q��i'Ҋ�l7�'m:̦S�`�f1�pP��T�r��avmHz��.��wf��ZD�4����Y�kt1:����S�cLV�-
��<4Ֆ�`���0V����M8@�H$�����b�9�v���X�x�뀠��טIt���U�+������9F���@�:Ȩ�Mf��{u�q<�ˇ������q��p��a��_����lgc���E�x���Z��m�9�P��:�0ݓ��ý۬>�����w8c�{<,3��u���zi�'6Qn�J.U��Մ�d��zwp���l��괠�*�ŏ��,JȒ��bf_E�|��g�[���M��R-���bD�j�;�]��9��!�}z7�����f
����^աf)c���'�ޘ\r�Ŷ�]�2>a��Ssf�.:�̥��m�t������1�]Z7S!e�F�`RYǫ(+�l;��k�3���pV��0�4D�:�p�ג�W<LbjЪ ��8������}�}�a��g%�h,���n	��Hb�ԁ*���C9p�C-�f��d�M޻�d{D�g5\Q����n*�g�W�����m�ۇ ]�a�mT�NaBۖ�f�m��g(�ow]zO��蔺S6��a@�-�K5��&��e�$�͞��Z�j:Y����	�]�Ǭ�M�9�c��;�Lֵ ��wad��A�����z�1vہ�e�ۮ��}�aA��bk)Y) j4%Ԕ����b�o ��/�3�Z+m���uA
�֪��)�gT���*�ȇC�-�|)q.G)�<����EZ_M�Y4��OX��Y�ī��]qӫw N��^�<wZ�I��,�z�¬(nK̭,��ɾ&M�8G��=��q��(�9���L^6j������F���@.f;ɪ�:�v�q-ͮ�0�8m���4�0_N0p՛IH6��)�8xqY7�6�<:�igC��������k[�%�
�!f��ljڂQ��n�'l�%�t˽�H�U%�R܎�F-��zA��fs�K�K
:ߞ�ɸ�f�V���p� �Ӽ8�'��(��/#>|pi<yu�m��� %l��'NΖ�޺H�N���E��8gm�
iGZ%���}�:)�9d�IPu)��t���v1n��g�C:�f���+�J��ӏw��޼Ӟ�7
���<ݥ�q�mktԡ������ֻ=4rvU��la��ݖ���f��d5z^)�����H�\�$Lmޗ��z@%Se�Q>,��P���T�U����Ds�����bޣ�N*k�U]���b�c!AX6n�`��i��۸蒸�<�X#DI��z�ui;വN	�W@qtU��>��Q�\�����QWNlLF��UbC���<��F�0t�t4A�]fX-�ي$��gm�nmsڣ�q�^�EqPX1��j�4�z�bqmzΊ,�[�����Q�r]��۠�븫��$��WI�`���#�u��V��1�z���n�cz�*)��4��M۶{c�wckE��Q&{����b���[&�%v:7d��LD�=[���SX����#��"=]3Q�fcSMU:���������DwX�cS����k���gOUڍS�:5UDfRgb**q�U1Eu��f��5���U�7M%U���Q�*�+]u$��3�������=v���+�\A�{��UDI5Z��&�����U�-��U�tA&�q���cզ*v5�멣mm��n�Elwf�������U&٩�54E�1D�A7lW"��4U1uE��I�WW��X�X&�k��zΉ��!6���t��E1GX��ﻭ�QMU�joF�4QZ[v��UD�ݤ��*��a��m��l�N���4�������<܀����h��=v��wz��ʬ�r�/���-rE�/���������|':���}��o�k�(.��]ի2�p0�_q�A�k��u��w��*��H:�q�-��mH�j�D8`�FH6Q~Q2;~j�$D� ��
EZ�oe���弞f��u�vvGd�ܜ�h��ʦ�p�����3���T,�1%���6��\��ɝb_�?��&�Ħ����<�y9�y7� C�<P�s;kaxf.��4k��po���
$@:K�0
*�tr�-�b�Ⱥ�F�2��#��t���DL,s�Y-��N�	�.��A����wջo���7�6�����"��瘸�#g�]��4\sH���_T�m�������=X�𨂴�q�Ѷ��f�d%�!��s�Sl�Q&@v�}kO\�o�ȧ|�PB1���E�͖�qXWdD�J�����g�RU�>�A�Y��x����̌*�� �l�6���{٩("l��f�k7_g����֦r�Ȭjބ�^A=P%�$k����{*.���a�r/�g�ۗ3jo�/d8:�DD?�ˎ|�ߦ������pH
ǰLRu`b4)B�	`!B÷��k��_n��+���!�h^zY�$Ao0�v�N�{,�'�SsP~��$�ħM�|U���fM7�Z�{�oyо��j��j������������_S0s�	�z�׉����}Q^�Y������^{���]S�J�e��^��m�������V����:�C�KY���=Vsɐi�r�a<&#�>�j�1��b��H��/b�E)����+��A���]�F��gnF�6e����;Q�s6�"�*�O�=�Ĉ(�4�P�HH�T�""!=�y�QIn�6��n(�g���Xn��Zr��$A�/A�-ᆷ����1�C�����b#us�9.�V�ixjMoEJCJ�i�eIOV��"��q#�����lD �,@ٯ�<�B�/�T��:k=w{m����t%�>)3�jPv�
�����.Rz��Ƈ-�`��ٷ�����(u�2�2I��z�r�遳�U+�5�{�г`ĝ�.�QaAgO2�
�XO��ǣX�;=�4��H���o���s��Pr�|���L g���g�еaD��瓙����$��Nt��Ş����طw�0\�O75u��Ã���� >'50̳rKnĤsx��/�Z�(�U��ћ�����@�f���Ks �ŗ�^�9�"]぀��hzr�}���]i��t�>]�K^/L�U&I�&�6��L˴�lk����חx@��#���F�l>ram�����B�=��癆�f*	�������C�D[.x��9��A�;+�py�����P+DQq1�ޠ8�
��p-�vƱ�nʠ��/��A{d�߾�-��G�����E�qb��
�U��f~ZD=���_���°ྚ�*��N\�rx{0�x8+3:��+9eM�n�̾]!oq6{D���ZY��j�h�ٗZ���İ�XB��H�g_(��_3���`[}�"�I�c�0<|���E���Xܴ���=�G��4 AB��� �(RL ����*:�^+yj�ag[���gA��zÒ����&����KcV�!k��2�WB���6��N��hf�`_Q�}y����Ϭ���޸鮯k����r�#��b�d�f���C ���Pp.VhW����n���9���$�z{��ߺ3��⢏Õ��	�h}u���N��ʜN��Go�+�&��χ���7o����LP��w9�Z�n<'�o��1�$��͛���a���W��vU�G0Bƺ���k��:�1�d����%�`+�0��qOq�h/B65������#Pi�֨W����jB"�z�_pvQ��vEL.ѺEֱ�n�1v��,X�-K5���5ݽ�7:p���
���Ȏn��[���:v�8�8���=7�spJ�\��CYYl�g�1tx�D���n��s�w����<a���~��1%��,����h]�Up:��֓�ok��}ܰ��۠*�q�,|�����zY�?j�ث�%��M�8���sV*���O��+�c8�<�>�/>�uN6��f�������&>�P��?7���t��E��~7��8pȨ�������p̮,+�!��Lŧ]��	�#���g���w�3�]��w��t�|�mT��N���;f�9�F��"���,e���R����,��Q�A��24��r��;�2����XN��Yq����]���?��=���� A���eP�)��B $E �B*g��_^k�K[8�??m�1�t�Ll'�oSm�>�z&g���cF,3��^�W�4�0��+X>f�"��^�����k�\s�C�t��.����3rJ~�^=%�ĈIy�x�><���}���y�H���w�uU�CK0:.'�&l��Fk���c#v����A!��pF�v;u��-w^��7����o���겂b�z��d�l�О�ǳ���4��4����t���V�����Ն��R��N�=��AO�|�����
b�� 0~�� x��*x3907+3�|I��.��Wvj������H(2��2]r����ت��C�������/�(�N^�"VӅ]E���;ҵ�f�[��|�кS~��[,%(2j��5i�R�`�ݠ(������?��}�>?o�.�F��D�9�k
B ,!n�B�a�f�A8�`	d���xղ�4�5����{gN}�;��9U�Uvw'w^#�,x�f̘03|$>��A�%:N��: .>�l�*T��
��'=�S��e*�����n{�4��9�2��mzc�)�`��L8�wQ���')�~oO�Yɩ=i�-�<kB���8+Heg�NE$����dIQ7�����-i�j�AyOa�Z�%T�؛C0�/�[�i����<Y4c^E$Qfb#�L���&�%��)�K'%�\���ʧq�e;v���8��`�{hm��Ey��1}{�{�����'�)���JU�U����� �R!�	�`P�Q)
���㟜�q�B�M��μ��Ǉ�)���$�����ߞu��9ϻ�xg�#ϲ-�?��M�&86ϯg��ߎ����7����C�𸔻^wm���%X%�X�e �Ԛ.�`A���-��}����\H�!�'ۦ�2BzOz)�)�L�3�H�����%�L��qxwm|ga������atd�@��Me,���-�2$�7��Lht�c]��Rrִɷ�
׫��w#ht[�7OC7.K�~���je�)�hz��~&/��}��B���K,}�_���Q�U�.iݕ=
=,G?�i˚Q5��� �1>p���N}7�'�X��\�Ĝ�%�ͤ��њͥ�Ɨ�w�dq�|������p�(9��
)Ș�`��&9��#Y.����ޚ>����܍�{��;�pxr�d�Lq �/\�o��%��4\sH���_�,�����\��,�v}�ݩ���f�󀇗�Ex����%6|�1��hljO��H��	�!�"�gyɈ���ԏ��5ǘ�EI��Ϳ��ܱIc�q�� ��U�@$g���U�e~S�$�>�i󧝑���/�82�:��ˋ�N�^�������C7�.�9�BڠM��x��۠Z↸���Θ���Z_���v�Yj�.�~b|&1_(���#!n�jrFD�Ē�9Z]c�ݻ:�R��]
 ��eiU#�ţa�ǌ6�Yǽ���C�����iF�JE�I!�I�h
A"U�& ���9u���H�v�~|Ǧr\�V6�!>5��@Z�,�3l�v>0X�o�j[�ML��텰�{�39<.���!㝰�2g�Z��e�K�uk�I��Ѫ-��8��խn�yIU��� ��y�*����L�SzTS	87��D�g�75��d�	���2�
��5��u�7;��Q���X%RN.�v*/�xt���~������l'��#{ڽqy�k����c������\�	�����d�s�|���A��!�O��1�ܮ��õ�X׼qv�a��)��E�c�F"�5�ܟR��(`����`�Bh=J��^-����wl<�	y�T:�
'e0�p�嗎\���'��ǜO�˿�J�.�9�2�7��m�_��1�bE��=<�7'�%�]t�w�$닿������U�+�o�2�RаND�fldV��[>�mkw�0�� �Ƙ>�i&5遭��hZ/qm���-o�0Z�U���YO�
}r���7�jr��|�0B��+������#'�M��� w��۹��
5y�+%�d��6�A6�L_��I�W�匥��5��S���4���_wg4�����6�nHS���l�'�g3$٠��Ɓ�6f��TR{�6��Ҭ"�	�ؠf�ޮ؅u��5L��ԧEU����81ֺ��""?�ĊA��0��B-4�O}U�]LWo5�8�vA�1:���h���z�O�Cz$���y�6ߛǡ��ɻ6tfy�Ҩݳderf�{@��)Z�(��LIz&��f]��-�z�ų��yw� `K{+S$\Ct�)ي<5niвy�,(l��#����fE���1!�pC/r�v|tG{_�N<5��<�r%Q�鷉�تK��f�.#��j+'p
zS�Vln�0f?��z�  �r�g�ގ�e��(��啕Ӈ(s;3|嗔�íyg����,:N&.�ؚ�i�q9Sp1�R��� ż��D��-�+w�w7��0��Z|kXR=u��`�3ǸBll��9�2\�Ksu%M��ሮ	����Mwu��K�H,����r�ߌ{�u�cռ4�{g`#����/�� ��<�sط*��gu�pm����Jea�Jt�	�����.�g-�k�<'��|C�`2XoyóC��+��k��
���(T5�Y���>�M��塞%�u��L��I��qOw0�sD��WMŻ˗<����{;�2 ��e1	��A��s_	�ݔa�(�a`#R���L�GOg�~Ϳ������K�Y�����j���F2�LPE���냆����7�'
�Ӓ�K.�3Ǐ\�$Ä'F�c�#���}Ե+��蕝�s5�p�m�Re�N��n�giꥠ����ȫ��%�:<���_���=o���S�B�!�@(� �D� %*4�a��0o���]�Wd������;���zht3�0D�	�E�F�҇O��~5�b����g�>ZG��'}�O�~4?!����^�!~:c���O�Y�,P:v���n=m�$ξ�9{��{ùţN��1:�������9�K��p�<�k���ֿTĶ'��簵�T�h��x�e'k�\�]�S!�1��^��?6�w,m{��?H�����.]�6�9���T7W]m����&��vf��26��X&������cя����?|�~�����uۍ�l�P��OoAб V��y/��.��9��w%�/��H�v�����b��̺�R�o�S��i�`�p�)g]�>���\_�L�{�ڌ�K<	��vq����� �O}�Pe����l�ùԝ��"��:"���t�چA��'>�Fs_3 ��硱��<���a���j�Z�������E��WA
&K�y����K@3=�aqg���R����Fq��j��+�8��<�6_\�����ׅ��	�����q��3�����!����
����~��������Q=wCU������u`�B4�)�&��kpq�Y�;f*���jwY����D����19��erU�*Y��T'#e��%h���蓙 ��g?KY��>�y��B�[���j�j�<쾫������׿�|~@��+�Ҕ�
J�@��HP��CH% ���g������n?�7��m�%�"������|F�>��hJl�#(2kF%?J3�(�Fh��4�LG��%Z��{볭.�Xxa� g�i�>)������I�#4����1���z��� �-�Ý�V�ۯpr��]�*`�S|$$�f�5?D�I��bS��]"�
�v��h~~+����=Ե�(W)�lz�\��@�t�m�5��ʻe�)�d�q=�[ԓ�ozїQ�"*���,vo����b�e"�4XsQ1e�>G�g��??/��v��Nr> O���&���+�:���6f�نD�n��b���S���M#��a��?H��>�t8���u>�{.���s��-�z��M��*�%�s����/4�F����t{�,gE-��f�/ѕ�p��_��};��8[.���ȝuC�E7P��ƻ�Jr��M�_�ύL��~o3�6��r�(���^�wl-��@����y�b�K�{c7�\O0�Ϭ����WY��q<�T��K:2{���[B'��C���@A�<�&�}l/B]��������1-��oG��K�`iP���#�f����te���FY�/��?V�?��kWyæ�mP���Q�K�=�ʉ�D�z�_Iu�w�iY ��=�j�Սqepr�{t&g-u�x�g}� dJh}����f�j��T��[V�9������|b6;��.��c��]��8�*�D��DPB�*�1 ��IB%?����;��Z��}�g�pG�� ؆*B��w�<`PZDL,p����K�Cs�4Yڸ�٤��v�m��Mj&Y�H�!��_,�-?�l �gE�6�/{qE��~�z��ނfЏ�-���١;��b�����6�؞��ͼ���n)��:_�d'ڤ�sl�vw�,`��ĺ��ez��摆+�a-^*ϩ�F@�z����l��ۭ�s]�j�r�>Ui;����g$�!��P����X�5@'ֱ�OV�K,���Zmet��,>|t���D���}����a�?�`��v�S������ �ɊN���x�T�e[\q9��y��4�Ul)��N5u@h\c<	[��E��N�35�N�*rSsE\�e�R��*��6�n]wv��v/�+��J��]�:q��E�.�og�Ƙt���gP�D�R��ʦu�v��^oq����W� �I�.��Rz�D�6 ͕I��q׌������#�i����\:��콎�4!�L1�Z�,��oeIo&��3l�ɬs�e�����\����������>�W�������{���O����{�^�w�������^^^����z྽]M�����<�����BZ<�R̤��3H#xZ���K�-C,��s�;6jU��io.��m���Gi�m��s%����+0\bta�/X�B�<5;8a���Q�ڮ����P=jIz��fR2�N&�M�U{DL��ꦲA	o����Z�R�ޫ'[t�EL��;��V^ԟN�e'�6_a�׶x�-���P��74kzr*f�YT�k��6��R��7���L�և��̗t�7�C�U�p�,�=k����-�C,|e���i��'��F�!u�=�%�kjP{���*��R��{�̱;�7�ն(���jp7t.��\�nmݩv��mR֛��E�*���θ��r�ȯE����
��ւe�>�ϧ5�����VJI��2��COn�y���{^�����m�Xs!��dk�	����`"����(s���8܌
:���\���a�:l&��E�꭯Zo��uǻ�vPiQ]F�r�k�����e��ɌًoW�٬eX�[ۇ��&c��������)�k'����q��n_EyK�e�Q�n���!���n�0�eX|Po���9VAR5��V�woN��mm�ՅȺ��#���p��*$�N�%A�ѻ�u͎�*n��IM#���/�2^��&��pp�?N�P.38�́=C6�"j��"����ZWd�]�-۱Y��M\���$6��a9�k�2�:��n�mm�|�jc4N^B�����9e�����O��k��C��&�>Ҭ��6�so.��e��im�҉���6d��U"ad�r�k�Ki+a*1���Y��lV1���K�כ��G��EV�j�N�A���5M@�b��A�䒘�&��������|���ث͖�N!�q��cSH�dUЪ��2��ݵ۪�д˵6�^d����IYjtZխ�]w��]J��޹����s�*�ɠ��=K9q�0d��g]8sn�.C;�g,:��+�\����]��)�5�+{Ulal5G��ct���sW��,�Ks2��s�MW�u��'�k:���ч�)+7'U�2ȵ��;Nv�q�ȃuQ_�p��T�S�%����En�1���V��e`E]�W0V!RҁW0��S	�F]�q���S�:�	ҭa��eA���N1�@=�����3�kn:Ã1�S�]B�=�������Ʀ��m��ݷ��ppK#�g��'�D^�:Öt���#��o�궈Ж>�ӗ��L�b��ʹ��^P�R���e��;�`z5��'��99����<�dz��uՆ;�
v6P���M�����յ�E6>Z'^�8᪓;�;=L��
H��h��sc2:���QY�N���}t���Y�zv^Į��@�����Ȕ�5V]�"�� F��Zĩ�-	MR��Lʗ����$W� &B�A�A=�%��u���SD��Wc!UZh���Z�RT����i�6l�32�1A�j��(���<�T��(�Q�i�F���v,kN�2b-b֢J:�"�� �Q��N �*��h��O���a��EST�MA�;�q5������:Q=�E#U]jd����f��ą�6Ƥ��F#m�(�-��MU�EU1H�cE���Z�UQk'��.�IN�c�W4:�6�h4�Th��T�1M�DD�QM4UA$�$���l����6I��j*&J���j���ՍQAGm_�l����֚�5�cI5!$�QE5A]f���4�UA4D��^�퀤-b���jh���Z�
�&���+g;h�*�����q�S��֫g5|��n�c����j"��"��$�����>c��
����"��o\b;i�8���Ag���=?���}����C��{4*K��f]�Oa*!��m�ᚻ�xhq���o�*����ԍ����zk"���S0����a�@��%
 i�hR�!JQ����������}~=�`�0Tߞ!�c�9��%��dI��«�%s�Q˔��),kܶ��a �yءel����j�q�=:p唆��qz��u]F��$닿�����n�e��v:�n�J�V����X�{B�4��9��Zz�3�~`~?W�ss�����}ak�m(����a���s���Z��1��s�w�pË0�<�Aˊ�|;"�g�X	\{�<$M�mbo��6�N�4��JT������z�Աj�:F����w8����&�q�W�k|��mz�|r�{�l7l�'r�^�0�u��̻H:"���S?4�Ö/x v������ہ��s��B�z��S�̯�f(����	S� ܷ�0�tE�ּ�Qq��Щ�[sQ}�ڷ�������q�3%o�e\f��tkNd��.U@ t�JL��nƓ�.t�MM	��}����j�o�r]X)������S���h���9�r��B��<�^V�:�^��c�ڈkZ��+&��zޜo	���5�g�!6_��l�9�j�e���������F-���ۘ/�aR{o��A�g^�ѦB��TFe��CeN�| ������q��z�Y.�gF�\���l�a�0&a�Sg*f�J+X2��8��xn�I�[lN@�2,V�띗�t�F���!��=k��r9�A�������o�_^������� P@)L+@�B�_~���e{���m��Ds���!2�F�'�G(o:$(�3ENNȝ�GVϦ+�מ8���/=-�ݮ�ڽ��^?�n<C.�<�����ħVRX&�IP���ǭ}��l�@����V�Q��'.��&��s��C��������^��2��^'I�)�J@L8�p�8u�����[U��y�E:���3d�����/��]�a��(�aa�]g���u
�Z驅ʛ��ȝ��e�P�4倧p���zhfƘ�	���M��D�iC��qWK���+������j�yA|e�*�?��_�� �X[����\���~��,%/l��C�	��}��;{:�^�K�Adw:�
�s{����y��퀃���t �~a�W.��?l��͍ʉw?W��M\�V5��:Mk
'�s����NU�4���L�~1���P#�<�s"TO�v�,��Ƕ[S1�Eg���٪�F^��~~�I�g��I�N�x��c�t�K�gbm�'b�e,�m=�w�zD����/���S#&�gm� :�Ǥ�!���1C����rԳ�C���n��4z*}��ҳ�̐q�� ��im>l8�����u;)U��Yl�W�o�n,]����yan�i��g��ŧ)���yL�kƙ�-~�M���P�z�z�M�,h�-�'Zv�{qu5��k�ݷ9]������	�B�R�	 �� `���������$��N��^謌����T�َ�uf�(4~���l4z�;�Xif���T�{Q��a5~`���7�w@�'<:JC�o_�v���ЫU;H��h��lEÚ�C���t�����ZF�w�)f�n�uXv7�mTounjf�T�	*������P��o#^Y�X�id�p.}Nl�*0Xf��:�r��ޢ=��1�>��l�2���lW�G(=f�'��V�S�`qmrC� `(�9[�b���2r�:=7�8���W��	6XFPd�U�4���Fc�M<X��f��j5�Mt�vNj"X\� "N�!�N��A8�bY'���+��5�U��y4M*9ҚY��r-����C#�N��\uA��.6W�]����G���'r{���Jt� s�T�E����c\f���"ۑ�\�m��4��_W?/>b�y�ߨ����3bc�����9Y\�v^�{���[ur������V:C�J�<�XLYz�#c���C��~����^�SL�3�w���v���^���0�Bn�E�?"H%�jM#�ȼ�<���h�C���?o�����ɣp��Ƞ��.^YR����,l��׾!,�\�l�C�}!���HK'+ks*���oy+I��%����QҢ��p�:�nA���ggV�avMz�d����A}:E*��o4J{i�#����t�TG�8K�ϿwϿ�����}�~_��1 �B�%(RH���y�ϟ�<��}|�[�8vv4��ݹӍ_�@y��5�����̱�Ëûk�;^���V������ =�ȇb��dN����C���Rr��6�j�zT���y�E�.ͼ��z�t;6�����v�E�K��H�4-Y�,8��,}'��~�Y������պ�]g�v���E	����H���Lk=:u�~K;�uسi��mųћݶ�!� LW5��?���e1��Lp~��_�\)��d��*zt�W>���J�)P����@�f��0]����5��tz&�M��.�q.9��5b�i�p�Rv�^CO3���e�^��㞨F��j*m�j��M������l�w�Q�;����^rz�N�L����ᵲ|.j��Cvq��$P�}(2kUr�$b��{6pM�1Y���[t�W���CY���I?~�L�F�^r����u��5A	�� ��V�S,�"w��Y�ff�'�榎v��θ�9�d�����5C&1��#��0�����؀>�/w��㡪��L����U�6!:���ޤ^��Q���ݛ����gcW47GI��씽��ҭ;K�6��C��FD�ڭڗn��o4hQ۩N۫���+(�A�&�78xvm�1���zerx��t�ze�⫣��������{����������f {*�y�35�k���|9e
W�T�SP]��^�oC*���H�ޅ��C.a'i��b&1�34M�$�w6�v,nd�q{s�$dU�V��s�ȶ:�q� �5äU@�h�:�^[�9�\�6��,�4��0��F�,`&(t	O�@������.5��/��B�����E6D�ZxHT��9�	��hOY�%��P��RS���E�y�i�Zas�c�}�C�����R~o-ȉ�M����_	�
�A������F� �&^9+�Z�˔��),x�Z�S��b�M�[y�c�P�g���w�Tt�xh�]&|(�bNߠ5��E��JI}cR�Rkc1�K�g_oZ-��谐^���r��(��Ѕ��a{���Q�9�P��5o�_��<wGC�0��,�>oO,��u'��J	{e/�4�:�����1������ ��˲Z�>���a.�|����7�o?�dZ�m?Mk�&�p�����=K��3�dK���H]B���m�c�9xֳO�޹��b�;�ͳ�ܤ�$�x���{72�t*?rW��y{�*�h0���Cw�0�a���Yk�y&.���2t�ױqZ ��Vh��q��O��a�L����r���e�|V�T���~�w'�s$>f_SÒ�x,w�c��$��{���͇��02�Bq�����d��za�Y��6�44]�������f������8{�&�Y�]��"�.S�NXE�0��xwQ!�;�3����^@A�v�ʦ��3���=��VD�.���:��xn.�@�",�|�I�q}e&1R�����S�k��Q��C��qN�y
^i,	��C�E�gӡ`r]�k��E<����;�_'7�H�#lm��R��C����ȝ����:�x�A�j�R��뇡�8���޿��%M�>�0ZD?�s�$�姎��jewt�q�~����zMK����`�	�Z4)=�G(]��ס�V���>ǖ�[rƨ��-0{/GEҹ��0�-�4_�B��h�U�N��������oI`��	*q������P��5����jU;����ˠC��nt>W�</"�@"{z{�Ru��K$�<��P)RaN*kx'1�9+����5t-��NnW��:s�|�Ŀ���E�=��~����)�.�Z5(�{4��\�n2�����ol^�;*0i�W��mvjiAC64�pd�S7O��
'eC�z�U�VM7k*l�����9՛ݖ�]r�OI�%���W�?�ig���ć�������>>_{q��5����o	eZ�䈷 og:ٳd�4̴�bѹ|��bX�p� �2����.S��ݹ��̳�%P�8e�� 2[���n��˥t����P!�-˴D�f_���+�O^������{0�x�M�ev�2���������G���>�� f��7����Q�A��V�����ǜ��IwO%�8�I~����ﾡvJ^�Gs�U#��dW���ۇ�7`8E�A`q��V�+ʌ�0�𝥛Q��
!�LK3)���dַ�ҹ�r^��>�7rʹ:-����3����~����~����3�EyEk'��3+D�7�;
S q�e�gӯD��z��f:��dǋ7鉿ff��+��H�"&\h��!�`�|/��|3 �͓�)�[����^�"ޮy�j���n�Ņ�������"��X�n��.�C���_F�f�Y�&��������X�m�U�5�Y�gw#a�7��2�>��4c���T ������c�v�I�OE����a��*��*3��9	d8�L�B�Kޠ
�W).���m=sͼ4��=z}by���(Lw&��T�J�����r��"ܡ5>OEx�[H8)��u��@ݔթ�	�$r��l�z�=[¡�)���:�`�'�^�n���2��yq��5X������D�������+��ds�B*����]cfd#�˶yv�ׂ�;��e�K��K��V�#Db�jЂqDĲOa#4ɼ�^O��	I��0̐˸X���ٺ�����v�C�sH�Ǹ���xEk�'Hf*�̆�1Jm��,�i"4rT����7�K���T{��v��wq"�̡%ژܒ٪e �I�7x%�z����i�n��5�2g�N�/"+G������<� ��f�������ݥ�~��:zkw�\^(���eza0R/��$vI���;�O^^�sX̓�{X��w,/�r�L���Rkk��es_�c!�{#� �L%,�^���o��!8z��H]���9��v�k���A�U��1I���"���j�'=8]����4[Pr!6ƻ�8���RaVf���a�j�Z��<��-G!7K�[��P	|E�j�0�����,2|�f���z��L|����L<6�Н3M���Z�vx��,����(�z��t��ܪ�[���>������p��`�<��۞�	�:꺞E7GOV5�ғ���@6�����Cf��A;3U^�����^�	��꤉��s ���||�jP��(G�7�+�H3�=�鑲g���M��S�|_�b�/ }�<���
������`kN|���'�>���]�;z�X�ޝ7n
.��P$@:K�6�>\1|h|�$��и�X??������f�/D��%}|2��m�z�'[>�BI��c�Y�H��H:"��W������ߠ7�����e�$l$?+r]�W��E=m��e��55]��O���c9U[eA�t�N�u�`�󶢅��y8�7�{^�J��X�e��t������f.�F��V���a��
�[�; VOh��iw^�lkx��b��7�ѽ�kx[�9
�	�<=���x{��xJr�V���1eՎ���s���4"���b���F]�^z=�lOt�o��,�d[�[Y������,Baqly�M\���ݭi�	,�Z��A�#8�86GPփK�2����GTl�:l�'��b���#&*&��m�j��X���w}E�cR���i��}��23��gV��F�L���X"K�l��v��u�Td.w�О�ok(⎮���CsO<�b4)\�L)� ;'�����-�Pd]	������O`W�Q����.����.=ݦ-O�Y'��%:��j�*�qw���c���P0��>zT}����ZC���������p!�t挳�7:a��ԩ2�b���Rz(��l�;�0���*���i�l��=(.!3��a�r�!�"�����ʒ���E��sH�ZF�C�[����!٫bQ5�<[�`DϚ�� l�Tz4�wøm<�5%P�am&@��C��)=l	u�m������Z����`���TB4� ʹ����K�bš�y��bN�����G�ן/���q_?S��=G���[��\��4�Ws�� ;�l��a ��"u��Bұ]u�.f�x�j�]��Ń�w��	��:������;k �ZZ��6rHg��[�Rw�p��CT��aR�.���^8w%#�2��V�3=�о�?ǽ�{�jWכ��w����K*U:���1v����3F@y�4���01��~hiμ���#�.E8�IڿChWʮC��w�Xs}�&��+	t�@pa�ᯉ�����ߚ�^s31'��h/�u�s�5�J�J~��oф�6��@�r^�y�ё.�m��r�$:׎����H���:��ɉ���L{!+_ -��1�+�pf�r	�v�lLg����.n�/i]Le�-�!��]��&B�� yO�+�f��u3ǲ�ӞbC�P,5=�Q��o��?)-��	�譞�X*YU�0((E�#2R{��Ƕ���3 ��ؤ��1K�C��?wf$C�Y!
$ךn6�5t�ê�x�XH��8�sI�j1���]��j���[;��52�_�ʕH�L�8u�8�n=3R���3��|��%�K�Z9�ԭ�
i��̎����c�fF21�����%6��F�~7���ܷK�.
���V|9�.�{Q�wkZn�vb�t ��tO��[f�'ҙ�yl�	�T.�g1׀g�{=>�o�������{���w����{�ޯw����{�>�O���sv׷�]�neiqBތ\N$�HE�	n�R�]�SE��Z�U9�6��U#�ˇ����d��Z�`bkk��p��Ip[���=�An!.�0�#)Mݺ���x�Ӭ��������N0r�a/+��V˸�w];��SL%s����2�`՗4?jM<�]I�Pt}2��A��)1ˮ9��ɲ���s�eF�ۅ���T���#����ūn��"C� �������j=�R��s@�ͻ�Ch[�}���t�7���cyP��ָӽm�t�4�f�nR1�|9lźq�ej�Ol=jŮ@qk��#s;��
�Pz��'��H���6�m��{�vW}4L����:,Q�]ˊ����"�j�]yA�0��+E���(<�zg9�̓��p�y �y�Yb�q���Ll����tOp��0��:`�:�b8]N��B�R���k�V�e���^A��r�>5�9=��n�L���6��.� �$#�(B^�'���0@�g9�]]>�ܩJ`��j/e����
�6�B�V��oSoz�̺WH�6#�L�7wvw@)HS^Ɂ�
>X@��9	�u���C�ღ�ý}S5�@� 
0�S/(k�z�tU�l�1s�%]ƃR�*ʕ;��eΊ�g_6Qgyi��\��ѓ���c�
�J�����
N*��EZU���')����u f��^;QѲ���������v��Xy�����9ӌ��W��ү���i��f��-����]h��1��b�6��۱Ƣ�u�/>n�V��g,i���M�r2�I��X3Y���(� d��6D�Q&C�L!l�{��ӻ�Xw�d��jG�9�N�X8;yY�c�ԣ���ڽ�z:�7g+�P�T9K���sC�!��I����E�ػ3�gV�j�#[�Kt/���"�%N!N���[Z�=�{ݫsv֥MI/�k������uV������Ť��hJ\�;-J&�,x��i�V�k*{ۃE}r�Lf9MM�����-i�g�@�V�yӠ5�����z�ש���m.��鵜���\k4p;s=�3��}��UZ�kd�=Yջ���O�{�a������s2�k]$ډ�
�PJ�]����C"���H��(^��<AI�L�ʠH�*����P��L�t�7�k���F)	�v���ރ|�9xve<���*�A��]���Ї���ngR��t8_ϻE>S
�g{�Ѝ�ՠ�6~�S��w0ˏ�^��u��{Ͱ�-�,Ԛ;��Xȯ;�u��v��y�ư��|�֟�`k�d÷F��:��N:͈���:���raW��νm�ݙ%KڔgK)٥Q4Կ��ҽfvLŎ�J΍�Q��� �c��v+)=Sn̝��P��Ǥf�4��uڟ<ƝY����U���ūF�����#s�N�d'����]+vvq�I:���h��Hil��d��;Z���w]%4EkZ�TDF�Emf؂
glDEQU��)��l�)�j���#b�E�q�ti#b��ōRP��t���v�Ej����**g���P�آ$�"�lQLUL���MF�3%�SgI��d���4�m�:�c㎺�������n��յA��Z�=j4AV1������U0USUl�����q�D�F�("���
�#�uw��&a�DZ�LUF�Mj("�+g6���UQF�����
6�kgF�&�و�P�ٵ��U�b��mE��UA�(h�H։�h"Y�q����u����S�-E�Ę�m���b�j*q��lhJh�(�cQ1�53�AEF�A�$�q�)������Y����UDTTD�fM��*X������ƫmUM�*i�cS�Eki�@A$׫���[yƘ��dH/��ߐ"F�a�l��iH�"ފ��v��h���7��coVh�=՗�a�%L��jt�9Ӷ�,R�9��qqY3{,jȚ�0��r����h��4�By����)��*�|Iq�$i�	�����S/!�dE 1���ǀ:
�"�&d�r�%�v��s�v��n�x��`��9�-˼�Ԝ��B`�E��D��k��	:�1/�I��Z����v�W�Ƀ����A�QqA����ZE�" �E�n�/����0��]0�/�~�I��V�������������ӷP0i�W��ký4 ��@���L�|dI�f2ԖV7a��GV.�<כܲJ�2�r-?5��j���^	�I���{����|��_������ASr��s���D_3�U��/YB������uV�y����i���8�!ã'u�.�5Vڬ�Q��8{O�&%�Pڢ��̚��-~J�S��i(d�ϖ��vMv���m��1���&'�.�\�����vm����cХ1)���3�ׯڏ&&۹�r���1U�FM������^�;g/@vp�>��F��؟d�L�F����+��r]�*�דxkm�G'���
���΃��BY�z���.���4O�q'��|�r����d{a,&���t��1��}ɾ���8��r�!��&����[�v"���D��ZZB����8���ʖHu�c��U��,w�$edN5�5�'_kG��G]wXj����A>WC*߶X�{�Z2k{�3�#̬�{��6��Tvl@Ι/9�V�gM�[�vJe]���[�cfwD(*΃9I�#����8S���
B�Vd*��i"�8� =�w]�}�f?�W�O������,�]����K�y�i���Ƽ����܋��m��-Y��F��q&���u~��Jz܌i�H�ݷ6�6���pIm�oNs�ǫxR;�jw!�f%9��v9���5�%CEǧ��0K�b�=�Jl�b4�SP�f�߶��a���Ȝ׼'�N��H��f�C"4= ��*�6�@D>���#nq¾k}�����co�1*���X��m�9��$�-w�����_)��= ��Q%ٲ��`��H#�9�S�G\y�f�,�����dO
��`K&KS(�j�a�r�� �!+�YN'�na{��E��ũ�қޖ�#�i'��*| T����LY��<�-��u�ΐ�zJ���/v�/��HPܦl�RW����i9	�^��O�H%�*GP�0��^h㺫6�����ܨ��������؍qp��^�zi��j�k�vQy�,����(��"ߣq���4����5���?$H�������?��uH����ƻ��2m�^?���X̦���7-���Pf�/8��]��nV���JȰ�#e���hFd\�j��Y~#��óK����a���0n���qӻp����2���ZRb�޺B� ӻ̅�aۥv�SYV`��r�����:X�1��ـ�;iчZ�*�7���j��a����{�H�طve����?0���;k��%�_7z�-1}0�=�;��v�g]ߴ�Sk�<ǣ��=]c�3��/���=2
���
O
��)����9W�<˗KzvH}^i'	1�a�$@;^&+��~���;���Ds;G��RZV"���몴�]s��ޞ���@m�-G�Cs�����j&Y�H`����sͼ�\Xo��2i��
 �p�Sv�'��	�u�L[e:ݏw�,Њ�t��ENϢq��M�S����r��V^�.ռ�k�S��&P�a ��%�j==�v��b���� Ũ��m����j�v.�%�7f��3�jq�{ [9~n�D^t:����M�&��V5j��e��?D7ML��Y�fwj"�j�,��X�WZ����'�ؒ��C����	�J};��TL�˯9��O���~����tLRuc�J�*�
j�q��d��Z69�������jcM���۰����w6�M�v��b�ܼ�R{�Jui�J��]�N0�vE�*�N0�{����m���x�Ɍ��wOyd�o��:/��|	`���u��5Ձ:�,��Ǫ	λ�Rs3HA�浐�K�So��G�<p�|z�c}���WS��X��ݜ)�U3���L��S�[���k�B�@[�s_S,..�,C�vu���k���{��z��;tϵ�|!��]l�ۜC`�I�0a�E'�
&��l��f��rZ�mE%S�7�><0G`@Єc;_���/�K.�0�;*Jz���c9t���iy@��δw���9p�D�z3Ϯ��d�+���~�<�ܪ(������]��1o�7�.BP#@������)�����at����PH�"�@2����D�^��]WQ�f��s5���6�'����#w����.�n�K:y�XWZD+��� �P ��Zz�3�|�<�j�h1^Ԃ�ګ��r���1\\��+�҂^�¨�X�j����&��e��3�����iy�X�ӗ1&#�(����;�{#ry��Ҩ��K�FR����0���{��g�I4��b�i�Ӝ����,Ba����Y�͛�%�&$��^�L˴=RT�]�+��W�ǚ'�-j]������4=��yO�(l��#���#ٝ���`#|���T(�4�+s<�sy�Z�ۀ��ݝohlg�`L�\>d$�=5�mcv5��7������{��3���t*F�� 4BWs��
�U�m
�M�I�7(�k��&�:�Lo��`�ٰm㹊˵lݓw5�7q���V%� Y�V[�5�9�����o�)WP����̓�λ�%Ԭ���� ��\s6e�6WSQƤݝ�v[��� <�V�c�ߩ�u�[u^��5�[��[�.�5ʨh�k�o��t�ê�E3���,`������ s�"��嗔�'+sy�z���$Զ5�B�l`�2�WB���뇭��.b��ĳ�鵕n
��0�ʴRs]\{c/�Z,��S�����ږ������L�F����ҎP�=;��4�֨K�9<��l��P[���=?��NRlg�}!`��� �f�!2��%:J�BJ�� �֐�N�F5+Q�����B�r9}��J�dQC��u���������O�fI�y�K Xʺ�~���.2�F���'�/����c�v�B
j�[&!0\�.Cu��<;(���f�6��*�ެK����Ӡ�t��U\�F�d\˖��]��B
��8Bn������.ڨD<�;���B���8�8����"��_��ƵJw�L!��l�?���O%3�RM�w3�h�ȹ��\�bS�(,hZr��'��=���uV��U��=��a���u�LɃh/�{Ljm^�pZÐaQ�s��T&%�V�.|e�gX��Z��������C67�����f�ת�)�Ǵh�iВ���PřZ�	��	�|�ӗ{�7��k�Νv�j���cj����`U3�\�+�|���H��2�u��3��c=IY�-���+�.�78���ܝ��u\��5�f �np#+m��xq�fS5	?� {�[6�5{�}��B�������"����;5[��S-�o*LS?K�1�Ǆ���;K'M4!�,e��wy[ �+�l��a���g��wh܉�lO��n&M�~���}�c'�X�.z3xw8�t9�F+ҴE�n���:%�,(h|.&%M��{�I��3a���ݛY��7��զ�i�!��!^)S���o�w�sy�"KJy���lF�ف�Uevk�.N�΄�^����>���(_I`h���r��F�����Sp��v�5��{�U���-�Mǜ���Ph�ѣ��^_��#Fm��/�ƅ��	��Pz͜O�UH�P�X�Yu���`�^JE;�-�Xt]��j�%���!5���ɪњO���O�_ ]�_:��ܣl���A�lT����#hh�a���{���FQ�9�=�JȮs�a�yy��׌�:��+��I��Gc�W�}О�-��$^����Uza0S|$GTVuE�n=�[7���4���>,zU�> u_�.�,��I��:皟"����ŵBH>�����l[U��.~شC�W�Qռ�5�����
�Q���MkTk2/">]�_b�ssK��o�T0�-�%���u*n�����=N�&��F�i�/.��ɖ�s��$�p�l^�ݷO(-*�ݶ�Xu_l�V���u�۬ =�uۺcp�W0��oٲ��I^�	�X��'+<�P�Ǟ���υ��D�Ɲ�/�5En���ЂƦ02�^�jNuD7����zOȲ�^��R������j���n�ws�����(M0�9���}��n�S�D�^V@�R�>���M*l��X��M���"Dg�8��C��>��ܑ?.�$W�R2^;xgv�xt��/!ye���k�N�$�0VW��X�&O�LH�c�/��	C�2,J��+��{�dW�o�6[;~3��Dz;���c��p{�B�t�\4pr��&->��^K%9�\!ھ��Ay�2_�﹜��圜�%�� �b���Z�^ø�z��9�[}Kܪ����YM����1d'�T�d���s��1�bbyۺ\���ś�����Ǧ%d9�sj�9f`�t$8��PQ�11�͎���s���4#�	v���F]���;�lY�`�é�U�[���K��o@ȧw������p�Q���*z�����PV��Xa���7Dպ˲��.�~z��è��6�3�ݎ����K2�G] ���8�)�
n�:P�ʐn�0����i��*	�Z�Ī��x�}�O�\��5O�$ܵ�� �ǃo9���-�W��s76���v�����p���%��b���l���|=�TN�<�;��+�|/T�=����\bT,|�O`�Oߒ/"ܸ>���K'�B����o5����^P�2�P�z�K*H�3�1��N�ʋ�5p	C����Xs�1��薶/̑���M��g��l�8Z���a'�9��오���Ja-��q��.[�>zD�d�)ۗ��o�We��]p�!0��mK1��-�^~�ʂ����4-7�U$�/�:q�٭����s�,����Ķm{J-�oh�,�9��}��f�ٹ��*S.`&*ۦ���(�
ڏM۳zYuf��,��;������ @�Ƙt�L9�C,�sRݓ=#˝h-L�IJ��^��p�2�iz'�C�3�ˇ��-y�!���=��Ol�&���K�����۸�7�s�/r�I�ҒǿlDh��S�q,X������l~=�"�=��<��X\�n|�v������<�n��QaK:y�*�`��(�~j����#�3��`)rnI����X.���xN�.��T�-�㊅�1'\u��\������?�R��L�y{��O6��1�^}	B�F!��nQƔuT�+I-�uy����jj� ��}�~�>�X{V��?}���}P�51�%���Y2�:��i�-�	JF����D���*�á��N����-�p^�(+x,un�d�δ'`']��_�ޯ.]x��\�Ϧ��X	��h�����N��?y���h�ϼ;+�kP�J���5�d�4�Rݾ{ aw6��D:�#e�ӻ�����������"O���9�>6<`q�+�����^�%�`v��bK�&��#��;�Iay�A�>I�	NN��l�-����M�ϔj~XE�0��;���c��UV_cr��,��3k7Cvgw l:� �	2�'D[*�>�g�����j�!\>�/�^V���W�<�_�	̛Eq^����`阖���䇆B��r��ך|.6.t=îyg��a%�I�(�k��Uţf��UyX�^S��&Sꅏ�aUj�R�%޳���u����|�YЊd,Lʦ���6󵺸jk��C�ןa�dnv���?)��	��
Or�P�=;��]Y뢛2��[f��;N�׆Z坠b�|�J|�0}^!��O5y�	L�1�N���6V�>���iW"�,Y���k�?d�;�W����^�����<� �B`�E�x8��=�+��5�o�R:'^[M˥��3�(�,W�T��(GE��0����y�f��NY�6�m��������������K�Uc\�g��ԗ4�����Kz�I��pU��GL�f�ȴ��J�y�n�H����6�Zr��4]B�VN}@�xQ���vt�\e��5�E<Ƒ�KL��z䲱0T蜉�*�M6�Tݦ�|�����&�"'Y�:Ή����� ��� ��o��1I���jVx���ʽ�ӷQ�NZ��mxw����li���Ff'T����*ժ5��6 3M
W㴡�Q�].��?7���j�R����������{�c2�$ޟ'��1�^�m�1:������Z�����uV��sז@����w��"���T��t"'ӌ.��@�4�Ź��l5�-l��Mk
'�s��r^�ʸ�gƭ2�յ�v��-�L���|:
���#�;សEA�� h��2�[+�T��x�}�.L[^��1�+Ǻñ��Y�׮��k.�fXXgc>���DQ^�&�<*g��n&I���Y.��X�L��h]��:�<��^=%���� �b�:�;xw����\_�T�vr���p�����{�G�(���h7�	a�����݂zT`�t5,�Z=/U/�u���R���1K(|b����{Y�CZwqS4fs�,	������ -W�^��e}�$EE��f'������}F�W_S�7���l�0�j��ԑ����yz||�����s���}��o����}��o��������|���^�����#ڟ"��q�I���F�J�:wd����bd�����wm�ǉ�]6MF��a%�)����*wah%<�ŋm�=�sB����z�.��J��F8�4�x�t��Ww
�A�n���"%��Ps�v�f^��.V�&��7���@`VL�Y�F�C:��l���}̽ۈC�\���0P�n�匣��nu�%A��/�h�((t�[Wc�ѝݵڑ��vDS#x���U��4_=4V�xygtH��K���Ї1J	+���cox̺��3��v4r
1F�4��Ֆ�5y��+֊�>�l�5��WR�jS.>hHs\8�zR�A�d�8�o(e�a�
s�/ɝ3�w;���Ð���M����L�ywi�����T�*�]�RK�Ď�U��n���v��q$�����j�����/m�T�1X֫�&u��d�|gnHֆ���L$��eS�Ňw6�hu�����;NlE��3rr��eӹʇ�ƍ?b��R��ȕ�Q��'R�n�a�3��`�#[D��[�}�s���tpm�yX�;s�2�k����t<�
�n�*u>a]Q��QC�Ч��w����D�W7��nh�ѹt��u�zR�c1֕|�t�;r�M����r�,�����j�C��P^���J۷݁���x��[=׎3E�.6v��0�Y��
һ�q7l7Luh�'Czf� �Yd������A������x��oj�q�j���(O���6�/b6���%���yx�m�m�ˌ�8y[��sIE�QD�$(݃�
p�0�o��h-A2���I'�YڵaT,1�-ZcqX��弆*6#u$L㇛{�GM�����+�J��9��p��0R�6�����f�<p����\U�Ç��:3-�v���e��F��.��	/�u�W9�ײJ�q�yo�Q]�.\Ne�7�0mP�̌���(UV�:"aaT��L=�k`��W>�ʮV����Hkso�Sr���3ҔӦ/P�J�sǷa���+�up47�lQ����[�cv��n�X�+s��KV�9֓�(���]GxB�)������y�.,=������F;=;�uܢ7pMe��jH�����L�������K�[�YRV��:=p��͚$+Wy;N�R�oSv��ziE�q���bH�&뺕�]��!� n�f��h�ۭ�3YA�� 8��_h��n�%�@ix[}�PB�/Fa��u<�Ŧ,,��%B���7c:*���8�g�-z��O�lf�bs�q�enWeu<Kko�i��vgUQװ8k�f���On,��4��kڰ
n���[g�P�,:3y����	�8��7n.�IZE�3��@L�]q#��{���,�Ū�	���FP����W$Xڻ걃����ǯ�MKl�SQ��8P �A LE������[:�1��6f�"*�b���UQuF*61&�r�h�h�QUM�4E%TE�D:ε3LV�E�q�)�ưD�1�Fơ��}���Uv�"&��"��Ʊ��m�M��E�b�уcE[j�C�lU4�d��:���5Vڍ����#c5�m%[b(�b�mEMEF��ժ"jh�ޮ�"H*�*��DE�kTX�j�VѣQA5�j�0ƌQA��
#F�����6�[|�]CV3��mJ�((����F	+�d� ���X���h-�`�(��V-F���Dl�t`�`�@��Q�OO/J�f���_����qiڕc^fS�3�����wg �}՝r��8{�E��:���#L;��T�dY�$U���>�8u$I��������`K���h�{GZ��	F����Mk���s�w{]RX�ݽ�[�b� g�9��6�}�|w��0D����+ںA��E�����il=Dg��݉=ݛ�X�D�O`�4��)W��Nզ�eo�:�()��>L��+���X��x5gou�8-�E��$�O�9�N�@�E-L�Q��|��\�� �ŊМ�e���u��x�QA�@�,�vA�;��O�b��:����wV�>c���J��^�[�{�S�DkuL�{�_A�0�s�M���Z���dz�5Kt�4�Ց֮��I=�˘ ;"F@a�K�i�#�H��Z���M�;Us]��^iez���~��0ܧdd,�/����t��C�8�z�?C��ܣG��H&��.2^C��u5�f�~HV�|���o��̊�V�p�� �H��Ż�l���?0?t�Ж=�S,��`Ǖ��e;$w!�)�,����N�U�%���GPh��ACB⟾����^^�w׏�fZ��Sڹm���×3�ٛ|�#��Кtl�]h��Y_P�[!̃���z�3�1S昪��#����r�,j4�f��4�ثwu��ZT�vS]�^�h��9�����k(�s�AAM^�*�,SO�n1����A"w^�p�O�
n?"#��7�m.�kG�Xb�"|XS�X��޹)�A?M0$89���j/��=u���y�璁$1���]��i�T���Q���B՗
_�wPny;��]��nc��:���;B6SO;ySsWs��ё.�0v�N�����58�o��>��4"��$�P*m�h!�u�Z��Mq��Ka�ӛI�r�\�m���d!���|W>���Z�1BA��7�F��K��nwty��r�A�I�jf�2�a��zw�$`���1��܂X��zP�m3T� o{:�2�0�}k�'�P%�Fm�}��3�+hv���G�6�*�AV=R�C"��'ح�l	��'6����w��V<��]B��*�
j�q��.[�:�L�|�5Y�',�ࡽo�51��E�!=�[���&I��1)դhZ�):�YgXb�,p.'CC���9�u�<�
Sz �q�"�؆V+e��N�L4��T��1I�E'l�)�%�*��FVf����zz0:�<;�D\�|�EA��3qNB~�&���˰�7\�Q���<�5��s�R��Z4�'���ژ�
�-�wv+����ɲ���_[�d�Y5�3�ʐ`k{�n�l���[Y4у3��}ں���Q�&]-��Ϥgv�K2i���_qk3�V�B��b��N���8����J˿L��G:R���� }�)��)kڼ���r�I�Ԕ��W6�9k?��0�{��g;�0!��f��#�\P��c#��������^��*�k������2��Q˔���Ic\�����q���|ɻ}qvtFU����ͣ��i�u�ĭqd�,
Ι���Ͻ��:w�� R1=���!}�l(���zq��"�~��Rm��ޫ�ҹ�r^�K���'[���oj�W���;oY�v;���3�Q�>���>�f뜺���-�����>�MKspSjJL��4f�16N�O�{@t�gA@x��L�-���2O9�͓��E�Q��j	�<笿#}��O�%�UQ��-��l��y�q�C�y�<����n�-y3sQ��N�լJ����m֭g�x:&>�e�A�ӯ��C 3:�eĈ�I�$�m�M�+*�P�z�f�w�@�3 �xj�o�,�)O�E�۞��y��ֆz#�v�J���}�ߜ�K�yp�Ey�v"�Q˝j��� ʅ���%'>l[����_���5�8%�Q�x����2�\r�)�IV�}�}qݺ��M����$�+j��v�ˬD�i��Z�;(���7X���z��áb�2��a>�B�;;s]�g{:a��rm���W��f�p��:�.-e����Nr��_2'��Th4���d8͝��� j'p�q;�[>��
H��|1F2W;R�GM��G���'d&T�B�ؔr����%8̥��p�6<ty��Sx6D�8l�Ղ "%ux���<���%5y���8:��=��e_6Gog^���:�F�[������\Ll�p�@4#�5�GE�=�XHK��{��Nrׯ[^�|A�K$���,ʁJ�
�\ᮢ�� f��L�z_�!َ�W.�m�rY�W���{l!��a׏EL/�Ԣ���P�hu6�;��f�A;0y���\��v+iu�^�ސ���hХgiC���=/^F-?5�����S�2a}�q�h@�{Ỿ�.�uU+�~�;#����!�ǣ�V�0��.�Te�dk)���5_J�vA�Q�G
!�6��}��b>/�>�:��بmP�U�Ռ+��W=�����t%�A��U�vvk��Rʹ2-�����C�w��3��i�f�y��]
GY[�Q���7��zҰ�m{x7����v��d�ʁ_�V�L�G0���|��㚪#�a����׃_�U!���s���&;=Ct"�r��9ҳM�Kg2���M��ܔ�r�ޙ�2�L8�]��oN3�A6RF� ���K�H>��E>].�Z�+�N��������T-�J I��	ؗ7��U`�M\-nF:���ޗ��ޣ�.f�+]�b|C{����W��������m��?'��ǥ�!��g���.^@�B�}�7��5Qy�����s���=z<r��X��vq����� M;H/���U�|j�/��f˳�VF��s�CF��t�^�T^=��uz3,�4Wt���PFL<�ش�9#5�O�{r'r"�7V��ֆu�DkKJ������z��5�#,�fcEM�L�8��Wu.�pǸ��'3�=��<2��,=�0qm����Q�-����!�ѰD����ڭh1�����@j�J,$�XPF3���ջ3� �]��~��ϵl�� �x��fQ�f�Z�=��Թ����1,��J<Z�\�B�(�|j�t�On��	�ȇk�4{�=�x��-r�Na��|��+�!	����~�Jt�	e�*Ml�P3�.s��pgގ�z}�OR]FQ��%dY�gl�ղ����48�);M���>�Ú�1���0Dܳ�+ֳ�eSs�w��#��#�a���={"S�(��,��z/�� oG���s3�Ƈ��"`���֏��Ht��`θ����I.&�/�������~՟!�D_U�˸_*�R˃M_ �'�Na��!�^�����iS��s��J����	Ѳ\w�8�Vd���K�Z�Q�����e5�\އi4��������ъN�o��8�0�w�DD��`��(ָr��̹�r%�Gj�G!s˔�k�
40��)�7G���o��-��0S�?����4�+(���`p���?�}��MuC�E7/^�2�J�ګ����ֱ�q��W�t�zU�T��l[�4v�!����0�]䭹N��Uufov'{q��r����Xu�������i�a�3�!�u�5�F.H����'�ms�)��>c"Ġm����86���P�hb���c���8�ݒ&��ͽA��v�P0!�2���{��u��'��79�&;Qs�v�tdMr�`��S>(�e������lvs��=�<�e�A׹�p���S]��յx�i�S�Q>��9i�T9KO�`���~�a[���bV�ِM����XW�4��J�+o'<T ɒ�A��E��*�Ο�]�X0"ä��o,�(U�����l���m�Pb��t��0�"�	�ui�r��`�~�ځ?��(�=~^�G官�ݷs�T�%�LT�������Y�骿�Y�K��]+;.�巌mN$�w�;!�%��bZ���G�:����k�j�6�aBݭ�l�NS�@]���
��3w��!'�%����MB�w��C[�Z�����Z��_/�Qcs3�'-�T�.W���*�0f���އ�v��8ɟ���e�`	�Z4)\�,)���8�z��r����.������{�sz�H����i�8vBnmЙ'�1)�FB0�'2Ӹ� �e�k�����akOMl�z=!�$X�!���7�����J�,`&K��%�^N�S�3�j�k�:wy	�C����/���"n1ޟ_�.h}u>g��l�wP�+^������P����tع�n����^������"�.z�wE�m���Y�v�vU�Z���
9�[�\���5�J�����#r\?��M���)��{6�TpT��t6�EM`��7��#��qvJ�t�*��������9���1(\=b�Oz��ˎR�02bc�e~��wVbN��$�/���C��{�}�.�����:�m5����G��	��j��^D;2�ۭ`��)��w�w�7��hL�;7��I���6���Z�<tm�״Ba}3�탵�^G�!�'�������O2Q�E[Es����s�蹊��sP�{�%R��=��ې`F�c�u�nk��d3UA3(�G:�}ƛ�|�+�xlͣYڎ��hdq�����9��ͮtի���0f��`���������QNm3ٔ�&2��حY{c��Cۿں�I;So�.<CuP����4��}�?�E#��ճ�ہW#f���Jg�y�N��:^7����,0��n�<����7�ʫ�/�;8T�8{#�?��!\%��a'5p�o�ιñ��\ �NFk�|m̎A���K�W!
�k齥���eB�b�W!z�I���O'�K�y�x��7j�1�Qk˝�O�-{��2�WARRq��g]vS-��j�DRډ\�� 9ם��@ƌ��q�0�2W;R���D��&BcV�
O3D�C���+��N�RLf=[ռ4�S�;G��\K\�B����y���Ji��F��i6���Fg_k����9�e�IP��l�=k�:yV�2E�-��0y���|��.�5�[S�]�{���myfW9�rE2�R���\��8������ f��B`�����Q��˲�nv�o���� ����Ǣ���jQu��L����-^w����E!���lQG{��`��Ļ��	�6��R%��q'�T@ŧ洠��y8�K�����7���U�-�[�i��Z5c�t��]��I�s.�V5�-�N�x5l��pI��ٰ��[kC�˕�;�>'t�c�M��9�ܹ��c�u:�T��d*��� ���;�ɛ�F�/QmfI��`Q���u����Ju��k�^�����o2�x�k���z��2i�5�ў��7��ݪ�V����Y�h%C�Ѵ�w�;�p�9���G��U �����>�s�/������{T)��6�q���J�wp�6�һ�4��o~�[K��~Q������P��<g�>e�H������cв��Lb݆��#����C�xE������&9���4�T
=�J9������ʛ���}�5�Q8��^�l�`��]!�$���|�������=��;<hu����ڠ?XT���g��i�6m��x,�
&�2��wPn�����	Hptq4� ��Z���W|��L��hb�[y���e�g@�^ii�1��K��ǳ�>��,�}�%����a	J�����Qp���<�.���=+K��xi/,�b5����ӛ��O={r2C�ԕ3U�A��|g�}|:�DZ�$S�L9����I�������RN�_�/�Q�����>����Y�7��#=]ո5 T�ɨZ�N���߹�+2��`��E���08E��p@?g��YE|��P��|�钫�z
���]W{
���]ەs4,�e�J�����<2C�:jJ�j*ݛ �VѴ00u��ͤ&7t���.�{��Q����ml����j>ǵ����uf�ӹ�I�,L��]�r�lJpB�#2�p�����
�Aq��%��?>��v��=�՟�9Qj�BqHĲOa*�e	H�Pq񨽳���{�`mOS�LdL�'駘WK�FY��Խ0�d��vI�nt�?0�V��eE*Ml�".�j����|<��!t�U�2~�	����yyp�	��3X�A�l3�ܞ�ҥ'��m��-�,9�k�n��,ڹ�����N�uu���y�#��%	�A�l?��$�b�m�zŮ�2���|y��˃��w��\�HTzi��@~��<�+ H� ���G�����^��B�ӆ�{�g<�R)z	Gs�,gûFE���!�6@`�a�q�2']-ݯ_1��&��n|�wv�D�C��f���<�,����=�0-�wf�1�3����!��w�E��I���k��U�jrhx�^�-�㊅��Xp�c�z}Tڛal�dP��Ę����N1�U�ži�"}`T����X���"��O�L(��<e瘶ۖ�1\���x4�������c;:���І���o�0$Gu瓸hQ1%ځ2�X��O�����yx�|���w����{�~�w����{���O��������d�{�e�x\�c9M�ю�"]��f���q��+y���^&�� f:/!@�$�Wz0mF%�1��lo�B�:vAIZ�;�Sp�������#��y�eh�]���3C��	�,,m�fuH�<7z�b���/��k��Hz�e��=�<�Z4����;�j�ئpM�9�Xc�k��v��]�-�#�j�}%nM������*�4��$�A��4���v2�$�ڱ�.(��jӶ�P�l�.	X �˼��*o}�ǔF��jn�����-�z��ڮ�L�Sq]��.Pz��n^�ԙ��p�c�Y$�t)�-�܄�`�M1�Q�3nq>��^s��V�t3
�x�u�4����!��Nl�펠��Z�3%���]��t1Msv-E�T:A���^m�J-����摚�n�r�3	����9�J�i+a�&��-+p�U�a��c2>�	�C5$3V��LR�{����SJ���u���GI��k�U2��7��̛W�k�)��i���Λ:���i�hlj��v�ӌu�
�;P>&���x�bZ��'V��K��0�[�`�T2���ʙ{�u������3Z�/����u��|rn+u'1��G���.E��kE���]�k��d)�ow�;�S�^Ӭ��̦�1�q�<�f�f',�n�a��i��`3[F�N%	`[$'���Y�*a��=A�<��҇�}y��O�/�U���I�
�I�1���r����p��<�)�57��e�M��8�f��9X�n�,c�l 6�]��hC�l}�hL���y;#��fEy��9a���vm\;0 ��:���(�/x�W4y�3�b���U�]�٧�_�0��"؀��/\E�3Z�dvfJ��f�T��v][�&­���8ݺ^��]ǋ_=Kd�O��cU7h�z�����2�9������O8�b�Ls�ʥrTm�
޳��yͱ0��"!*���T�wMӛ|X��/��
�Ϫ�]���m$�m�b�9K	���s[2�u;Qp�\�쒻�{��
���yݼBvA�p�M<�ⷍT�Io4�Q�V#\�:��\�g7�ƣ1�5d���>�� ݸ�:����AIƤ����]`�j2��:I#$be��.or뛾��f��_G���2�:}��{V+7��y�����m˱�;fڷG:�M�4̼������V�Yc��`���u��FP����D��$ND�ڤ��F5�k)c���!�j�S\���S;G(t���� ��v4�2�:'j�Ȋ���%���R�k���w/���+0��7��<�9W�������x����I���� ���+�_;�oEܛ��� ���<�C^%��j�$�8#l�|4,�]�OQ�:�6/d���.���ٴ�e�\Qy�wt{s�wu��>@����j	�m����h��S8�14SDm�lN�����kZ���-�F��CF˃F6�U1U�S4m��R�U��� �ձ�F-E���3TTUTE��D��:�F���8h���ح�[��=ƫ��V�&�ح����kIZ�AV�h"m�[�6u7��*�""��i�������*���n�:�n#�(�~���Z�EmZ���u�Z{:*������(&����7GN����۞)�QV��5Q��5Rtm�E�
6;�4��`Ѫh��������.�]�Rh��^�Z�c[�k]k��mj'�/��]�����������aL8� ��9	Ӓ$��T �cGa�~?N�9��.�ъm�ʻ�K](3Wg���C"X��kF�2��Y]�ֺ#�	v�zW��Nbe���@�J���%�A����6S%���)"bCM�	,� ���C%�A���]w`ϳ;k�*4�IW��/�+��T5Y]�=�w�$1ю�q���l�K9��]�Q�dPr}Tpۮ�j%�ݢQ�C/e�A}kO\�o��f|�s�g�^m�����ẝ���P��[y�����W(2D�3轜e�)�>�x'W�v�(c�X�':t�|`�)Ȭ�L��0�	�֠K$��>��q"�*��݆�Z�;�t�:��s�_oo0hB׆��q>��أ�Ddv�!���	�F�+�����l�i�Bv5�Ɋ�P�;ť�U�C��g%�C7�(S~f�0�����=������r��w�%b��]5�0��o#gV�pP�8�|�-�W�q�!��:A�Ð�L����n�~�j�>�m_���^�[}܁k�`IuĚ�������@���"'�pG=s�e^����Q�����Sq�1!�1K#U)\7(�%�7@M8�H�=5�N����<�~��(�0�A�? 7����N�~T�b��+;I�P9+�Z�˔���5�J��gw�X�#O����~ϸ��n�j)7텯�����aؘy����D3,yt��Տ��5�i����q2m=F齳��'[vH!"��������P�h AYf�W�>[r�8��&qs��֏�f�s�"��:aHec���vhs�ݘ���Ö�I���*��{}�Uf�{��r?a޽�公��o��6|�E��U<h�m�h�*�
:w����0���ťõ姼���NmF�-�5y�>`�^suϯWfhˊ'�s�PK�Z��zs^2�s ӑ=i�)gl����V�@7���~%A��ag�!��\�.��nԤ�����B�q�Fe��v��Y�j~��]I�Cu�8o�����|�z�M�h�ߖ��NT�F�'�
����z��C�Ir]����� �c]��Ϲ��046v���Wmr�ʬ&5u���l��-ؼM3�dYSv������4p}�ٚ�&{&���Ts��g5�U�[:dk �%��SГ�m����28����%�r�r5�q�髦.��T^�Z�O����K��u�1�,2./�w5��˸T7*Z�J��� ʽj�*�Rq�ٖ�iJboc�j��YG��a����}�{�@��>g`��1F2W;R�{��Rl&eB����`5b6���t;�#z�u8��x�f=zޭ�S�;@ Ŵ���	W�n�1��1�xݣ6p_f�Ì�ܓ}]�����G�ɒ$[U��^�m�aW��w�ǹ�Ե��;�v=��0Tw(X�)Y�r���/�^�p�����"Y�{P����2wfc\���{k-)u�K�֑�8�Ѡ��S�j���h<ڧaG�ܾҝ,��B%�C���qՕ)�j��ocg1���>
{w�!Ŵx'D>W�N�k[>˰�u'1���pZUzA钝`c�=�.�eE*L(?Es����'��@0�ansLE��y�Y��}yS�B]�А�òL=��(�a�T�u��)�b4:�r��]���ϯ0�W ڻ4�*e���}n�&m��t�(q S��'���5�S�2t�l�U\]޺��;܇2��"��O���Z��ΝF�0��Ք.�*�Ş��5���:k,Q�H���}��[�Ti��\�� ��!�G�ך_����l[2%���c���Q(Q*�x����ԏ?��N��T�ek���`����>�W掯�4NZ7���0�d�.;�;'��J�h�z5>�?OLU�|g����;�5�V�a?���(��Kb2�e���崛���,;���n��}�)��g��~=��׻B��:�;F�D����᤽0����r�x�P�Xz�"zo^�{s��ɠ���l�C�$@28�v���G�֘v<s�f~@����NY�ﰠAY�fQ��o��7�ۍ;�`�f��s�F��L楪�.�j�ԣ���Z8�1Ӧn�9b���`bؔ��Evͼuf�9xkx�U��wmM��ib�̹}t�k�l��{C�l=0r���X�+�Y�(�+ئU�w�ݴI?tWI��>2�i�C�I�/�wW�fY�h��,x����7�d��g�R⽴!1�{���F<���	��<���S���{l��h<\��+:�w9���1!��-�l�f��^�ʙ7(фJ?�.�_��̷<�A���xGUf!�:����������4Jt�[�}�{ǌz��;�&�F�qT�䛼u����v�s�rת�B|3ͯ�Bq^F"]'���er�
����f�t������l�F'���9�t>09z$!#�O;z��	�{s�_��L��*Mmb:�f�ٕj�b���Dcv��:�b�5�~~b��Ƹ�l$~�ܜО�Ғxa����E.]�d;C��q[�]��=��c	e�1e�>@�G��tc"�zz�O�.%-W��UJf�}`e�X���޻�8�~�4�r�i��Qӭ�A@����E��Q�0�s���^��y-�+�%W�����L����i�1(��^�����������q���<�7��<��"tʽw�!�T��`[�b����f�e,=|�gׂ�W�rFV۶��MX��{��X�����Jgy�[ݭì=\t�[*��Q+��MW�*_j�K1�D5e8(�4�r�A�@o^e���g�:�/`�޴�0�q���q��x��Q�M*7`����j�t۷��ﵰ�e;����K������j݂\}೧�Ҩ�U#+c@��"bG@S t��u5�Hy���=�yס�]�7��y��d�Y�: ��U3�#�l?�C�jBY�͆�+QV�{o�C�q"sL>7�.��F᡽���|����b��-x��O^�^���� ֽ2���q���&v��@��V�yR%}��A�4(bK�[��V�������ohv�#)��>�Ux;��ʇ++�I�2������kT؜�t�R���6IZ������#�qv^JB#��b�ԟ=�6�v6�4!��["�C�v�F�7�gU�r&q��8�}1j*�����ٶT���	���@��y,�'zx�55��g;���ُ,H!�X��ғ�^���ӈe�#X�=�q71P��~\���6'��٭=��vB���)Ĉx.�c��B�?A��	��"W	TXH�'��'��Gp��>���.0l��oA�"�a'i�8ok�LY����9�N������{��ci�F�w���5Cob��C.1��Z���E�Y��U�?�h���~���mW\���仚2�V���iްWi�R��CI���M��oq=�Na��9j�MY�����sw�q��sm�h�s�"��J����.��w����mu�v�W[ri�kS��+��F�Ԭ�Z5�Mџ��ր] �D9��Z�>�H����f]Ujº�M�wm�-lL�&J�n�I�&G�\�%v�1��������uF>�Z�9g�[��u�6��tl���r���)��P�]�����e���y�����Ǫ�����[BǾ�q}���*�]��K�����������;kus�#r������0v't�G�9�9܊���MyV�{\�zI�ݯ�����Z�u��=�0�`�H��;��$���{�.��I�e�|ٝ�v�1S%=���K��zDt'P ��{7�����N�^�o����M�k��n���4{�!��0"ϗ�U
�E7��c1s����_�_wGj��?5�>�X��G��Y�$ㆾW�)�=�	s|z��G�-�n�	�H�q��?j���� ���^�ܥ7��_�Z�Qe�K.�2�cu�EW�T��+7�rg`���{0Rf`��Go�m�& �]wf�!U���;X)�������J�AE�n���m�5�-�5��X"�@Ct�����B�`�vwf����$�u��Ў�5�Y�J[=��:����'�foW�f��K�oc�#O&��Pû��PF&r�"�V��u��8b@�{�4&c�e�O�"�
��x
��$q'S�%i<Nd�{�T��O�ǟ��%^���a�{]^�	�:b�.M^1���������ȩ�3V΁�Y7!���}���hw�SK��q����~�-l���<�zT�U��%�u%��U��'��3Z=9��s��;��p;g�
�1���d�U��t�w<=ڋ�ۺT_j�=��v�L��P"�:�c�v}�9��K��JI�06�d*�m�-j�;��&��v�1��/zU���؟��՞I(��j�>�4=Uv��ڝ��J������.�x�m�5�y=��)����"�I��7����k�|�;&ڄ!��������C���z|�P���nvaS���~
�4,=���ec��qNy�ֽ�v=Ҩ�N��H���q+1�tKggrǤ��j�;BtLF Uƺ-��wJ��m+�6�d�.�������5򍫇X:����w:�!�h�S�U�ܔ�5���zp�w��_踬&�O�����qG�"����dE��O����#��n3;�-��GHp#�ة����>oֳ��C��w���\>���$���I�b�Ӯos��@<�-վ�p������fۥmF��Y/LV]��L�Uc͞��m���:��bO��?�{o�+�U�$<ڸԍ+#F��O^�����R#�tc���J�sh�����<��:��ׂ�^���E�)ڏE��q��VY�:!�T�z&=��70N�L8�O�5�X��n����q���sD�VX�����l������]�_C��8�ں�n�޼�1Ѐ�x�������G�.%̌AV�{7�9tTM�}��(V0�ǳ�o��B�*	U�ګ��iȹ�q�uծ馽/�<�z!�#c�7��غ[R9��'��T
J�����(�l|�-���Ϸ;��s5ޔ�)L��T[��[KDL�S��n��t��:P�OJ����.Di�t�eWX ���7،�O;:�eu�v撵ı[��`0�XI�o27^�=�e='X��U���^�oTR�dk6vQ/�av3�FȌ4���5';��*^)�&���@�v3�k�v[���[?��D�][�[����/Ϫ
�袺���{;��{�do��2 Ǎ��\9dG�[]p���eU�Q�ҥ��m�>׍��졪�6m�l��S����X��H���I3ׇ<�y�m�n�����׾�	wN�g��C��k�7�����uo]���E�G70�WU=�qs��c�����JE��4���O��>z���WHc��omvpԸWC��co-J��Ǩէ�yԳ��5��C�:����^iD�7;#,%¾�9#�.��*�d ���ؿk�Q�Y��y���Τ(rTh\�K�w�r���\,5?�cg��ۯ;y��3�$%��7��2���k����w����,�2��牤��f�!��w$����9m��@��X1Q�>-�ތ1��/"���C.�*ވ�J�S�e�Ջ���j🠋1��:�]]�!Oi��'
$�n�s��ha�pU�9�ӺL�|0}����\L��qI��t�F�����7zP���w_Ρ8�RO{��&sf�	'Yu
�M�,ӊh��m��Qu�s�9��|biUȾ�:���h�B}��VR�V�GKw>��=+a�]K^����*�"���#IY^� �4T�	i��3��S�3�t�c�&^�b:�Y�v1t���(�ot���,:&�9���}�zwi=�2|f�i���؄�z���y60��)-��s�ы���$��,c/wl���\�T-nS��"�$�z���c�Q�*�j��9��wov����䒿7J�
&[gg�X8��t��??N<F;�m"R��m9��������9�aE���f��T���M�]�]'A�S*:�JMǍ��L��j�#��Ī���*�*K�F�B��q۹tg6��y�1դ��=�#����	���F�a'�d��r�K�Ub�w��dd����2+s�uNC�L{ty���P��;��j��O-��{}ޯg������w����{���g�����{���OOOOOw���E�y@����j����MB%�b��zTQ���T鲩�X�;o:�kZ���NBv�r��A1`w�ǯfFr'�H:i�u�D�A�.]��Z!fܘ
�)_Uj������s�v�0�a��oH#wI�E�ވ���A��:��K���Y�뽐T���J�:�z�5e�9��&�\YI�3��Tݑp�ۋ��O]L���ms���W�u>����%+.�i|����h�n���*\|�j�L�݆T���nm�ض2�GR��*-��Z�Ie �T4�.8u.�S�U�L��	n��W6��*��e�e�J�HۧY{�,��(��J�����љk�Į7or��a��Ev�֝��vQ���K #	8�0����6�FQ�VP/jW��F�@ݧ<��B`Ĭw�b�WE�����y���WSbk�%󨻊mi���{�zX�UC�%ѽ��^EvR�W�v�ӣ&Xab5P�Z�����F!X��'f����\�˺R�9�flU�g{�H/e΄<w��Q��[�pj^�G:QE�u��BC���#qF�}o�\w�wHl�pA}���sq;�jQk����ވN��׃���X�7�����a�H����`�B�}�o\�b��� �[!f�\spv�5I0!+�Kǻ�$���ֺDJ�+V��x����pP�T�C4q����*�w���I�e�}���H��6K��m�����72��yW��s�\Q�؊�w1�:�L���I��Uu�oW^�h��;����8J��B�mć!йAt���ҩu;����+mne�<ٖۜEL9e��i�s��Sb�51�f����0�k~Wj�^+�{��]��̴�,�r��y���]�M}�L�\K1:�{p���T&�س�w�T�mn���wK��ug;f�{=��2L9|�n�;���ݽp޾FwV��E��Sp�˒;��u͂����c�<�Z�ą�[n��,�����u/��YBd��_;��C�4��k�
P�]Y�%��B�1Y���p��u���|��6���s��m��mq5�:���0��D
˺�j]v�`םT�[0�kR�,����q��2��M1U�}��{xF�N��oh:�6	i��S��L�$�h��A7���5d��Z����8��v���B��j��U��C����_<y��"q���1܉�/I;��*<��=2���8e��ͼ����"�X�:9��\a�l����:&��PlVf#���jxZ9z��:U�[��8�B.\+I����ׇ"=] ;<{@�^�ƈ� .1���`��Rv_�-	��XnD�iGp��*�����I�حT�R:-ʷ���8L^4!�5�3ٷ��2���[���9ޥ8�s@���������`�GE֫�N'AIVب�.1����V�&���z�1>��U֭���cP�V�֝��th�#��j
�v6��&�l:
��RIv\LTu�"h���6�k5�֨�6MU�D���]j��"�����%T�LUS1v�SEECTTNÉ�"���-�E �ѡ���T�Q���*�b("h�v�CZq��b-b�(�c-?Y�X����X�U�T:�(���Ӫ(t��5���:��LIݺf�*h�)v�%�i�th-�nڵ���b"&b*�v/�Ӝ���Ϫ<�2��̬��Վ�v�v1*�ġ�T���$A�vm�A��.�����eS�2T���b8K�s��'���VK�$��*���<�K�P�z��#�[�����p���G�/�9)���ً�c�q�-�~kǳ�'��a�/�|��!�(���Z{�^2]}=H2�*��Q��b;v�s���ua�Wkc���8V?c�>������[�a#�#�l:*=�/̬!=��yY���2��\�@�����ѝ�Ѻ�z=��TF�MM�B��͔��e�ќz)�t5TAP�rhL�G�.nq"��(��g�2�J�¥�`�g^�b�i��
�9笋S7N�F���{�s@bī�2-�+���ݼ��U�׸6O�UZ2�9U�4�j��@�ȻH�\H�g
-
ڙ�������	����R��oܕ�WT�w#i�	�xwL�Ov�a���5u����7Dp���Gt��1�JK��ĕO���u�oG�ܓ]���my=�ǹ�Rߤ�̉�U�S`ca�a����̾y��G+�o����	�$�_�lU��{��k�+w�8|e)���kAH�kr��&�M�4&B�p*˳���S�VG�5�"��W��s�k����Ӕ�O&W,���Vy�}�T�Y}��<(��J
pP:����W�[Ԋ��R=kv���k'�6�f+37�͹F=8>������t��S�G���'��<���R�M3M�o=��/a<Վ_��mJ����j�{>��Ϛ��c-g��L�E	������M�u���o�:qLی������w�i��/��X�0H��>�$����o�>���vD̩��"�)>��fpA�j�����6y��n9��;���B�U�A�`���+��<�Q+>.kNM�C��1��K���vn��'O��ȁזl���#�������n����X�S�y����h�ey(��$|�=~���Wt}�oe��w$X��$�0��c��J'�y%E�ΰ;5=]�?{���h��@̳^hT�ñ4wC��wr�4B�����s9,��D ���x���z<�أ8����r�3��0�e%9�t D���*�i��nL{#޷$^m.�o^`�UA���I������Y_r��ef�;B��'j��t�TZ����8Di3[�p��kJΗ M8r5���s��,	O^;�yV&�g.U�Vz�Eȉ�� ��+|��o|�u��.���ا	C�w�hH�H͵r�a��L������4��#vw��!S���`�B�����=k9�q���2����u�A�<��:�p,؅����K��mAJFR���P��۸�-&C�� ͎�����;�9s��L�}r*`�7����R:��T�4�a��М���ȅ��n�����t�G(
���P��ۜ�;�%$S�R����Jy^���}=}p�|��#�d��6� �Ð���g\�в��
|��kH9��޸!�W�L��-�\�=��7.�7��=	��*N��+6��r��ug�zMv�;֒�K�uc@.��[\3W��ܝ��G<s��{�G�z�m�eHW�d��U�6�u�5���{+�r�Fa��P]7��ی�K��p/�h��_���|⟠�{v�q���r�n���<�����y�즶nk��ۤY�ڄ��)^"5�$�6��_-
�̛�0��x˼�W�X�0������5�sF�m��&^_h�`TXy��E��ul���;�����"��vS����e ���z�I��6�5x�I��vv�_���k�w�/0����2odm���$M�~Y�ex>����Y�jq��Q�����GC89�)��[�[�"������<Y���7���5���9Lc!���1FSLN	��Ǹ�묫]�2v�h���^}�H�����9m���ϴ5�<벓U�U���S�i������%Q5uY������HHx=�_�h���Oi�d��� :Z7+WoS`���`z|�r�'	�#{|��z��^H�t�[M
�
�&��//h��i���}��������V��.��
�Q���p���Fwl���f���UW���0=�3��gIʄ�q�֦27�wS�_#��M^���5�RTQR�T=��W׎��H����݌K���Ƚ��8!�Glq7���JۯԊ5����̌���{|����x{��"�F�XC��+�b�'�SB�m䳸7v�Yi�Ka�,6ڂu\R�[�A(��i��t::�4L0s	�{sH�[Q8n����L���P��¨[ʓuef:ݳKkvj�u�κ�\z��_^�Ԥu���N5���J�*�-g]4�/WF����ʽ�^:���t�6R�[t�Ϻ�du�1 Ա}���gl�8+�#y�p�3�ؕ qtr���a"sK*[��;K�����j��l������D%#�y*�ӵ@��K;���7u�f6��p�W׻θ�C�`�f�5�%�#�O�.�w��\�m���[e�i4؍���j�<P��Sto�h�#z�b`�Mji�iU�W�nt�@iIPO����ӝ��zp�6�!��0#����.(�Q�u�OkŘ�ظ/�P$	2	��b;Ews�׏=[䨜��Ңq�͸�{!g��}��:��ٯ�&��t>r�]����|swo+Q�n�k�k�z�����2"�ȍ��ԕD���~Όꎷͬ�y���nn��L�2b� �g��	@{�539qX�X�>�?�ގܹ�Nu���Ç��P\V�"-�c\���D��\f�zh���5�8E�(����@|�O�O��:h�Qk�֔��?!�Q���sQX%���Sz��^�_?�xǭ_�Pt#�&���ݦJ�
�S���c!�f^N��@��y�R���W����my_TK�,�!Tn~�k������&�Un=�r�2�4|!���ܒ�a:� ��D��k@��z�C4as������w����M�$���B���Y�`���"���g|���][���B�T�$���xe���W6������x���~��>�X���44\�)7u��y���T��S��p]e�c�^F�V�<��3���:�7��2l�dOi�>��}@2n�������t^��8�<mlX�cdc\�ح��j�y���j*@���f;[`0��!�k1�E�뮗0��y����6�G���1^���k����os��tx̄ǵ{+ms�i�����'_������'�o��p炴��D�#��d)��}Igm�pTƾ�A�:��NO��7�{5�d��#�6w�����f�ruTձ��Y6�g~;�'s^��9��ĝ��;7u�26W���c7�s.��BV"�A^�^J���`=X4��_d���\/�di�;��/C��L8&[��v���-��ِR��Z`�kf�|Z<�L�͝kz�!J꒭e��}ؙ�jn�TRPl	úQ��}�yo�+��;�O���pv�=-�`�0:�H�u��#�2rCc1�
�l�U�6 ��;�r���ZoVZ�����ۛ���ih�����2
��;ӝ�Y����ǩ�RoP^�{��ȶ
�S�Ng�,��D �5R&2*%=Ӵ@����U�{�n�.+��.(H�C��%A#�#6ԋ�P�?��ю���]pm߸�V^Â��v�}쭣p��e"��Pd��G�&��;j3f*@L�ӛ7������D"#Ǵσ��m@��2�y#*��g	�=v3�3z(��Un�s�����cĂ�/b�B*}{^n�������-AGP{�;E���U��7�����#�_���/Z(Q=ӱYu�J����H�<uiٖ�x�۠�Ð�c���=�"���R�TI������n�.���#��N+p���-�5m��ˬ&e,�V��u�>SF���NԕC]��	�L�����H\ٺ-u`������YB�l�GP&%�+��R2�R�N[w0G�-�vw8���()�e�D_N��bk7��{����m4�i��q�B�S�� 0��/h�0ֿM�m̳{���҈W ��P�g�F�Z)J}��լ� (`���k��w	9͊I�����T?a��vUutvU�{�L�3e�S�qmw#��s1��u���V$dD�o0ʷ�y�_V��:�<�F�jt�c}wݽdi��C+�6�������bzs���L���ĹJ��E[���Hrd��l��Pc���SH��3��
��)���3��/{1s��Mk���9��wAR	-E�Sʈ�G1��������i+C���8O� ��i���(�.9�`f
�j�������o�者��&vzӕ�ye�|A��	Ix�z���vW����������;��G��� f[ȫ�\�w�Iga�f����g�̺�����\�����Yc��lfc����w2l{���G�{yR�%�jjMX��!͚w=@��	ov����q����]�q:�\�-��z���f'x��݈͐��k�;�ō�$L�eb��X�U����`��O\�U�%̫�g�nÚ߄V�F.��Wq��X9�4��D��k1��oٜɷx*i� s�>Rq���=t{m���u>�v^�Gyy�%I>rMS�ܷ]���i!pe:��+֨�w_n�vV�K��=�{\���Kt�(�m���Ng3ǝ������?<s�:Z��qSKxz0�r\vg�G�$��]ŵ)m=~��mؕ >��E���4�!%où�_���ؕP8�'��*	w?H{w6�w�0k��}�K�����D��ʮ���,�K~~���S���3�(�9����7:�����̀�|as��}h�{�VhNzf���]���!�OS�r;��z�����]/�9	Ё��>�b�T�S!�kա�jĮ��*�(�~��z2Gtl�v����bD���������|���]H� L���*1s� �e�����(ೆ��"_��^6*�#/���Y]��U��#b�n}�Ꮔۂ�])�kD���D�m������f͢P�-�)��q1����ƥ:�.�E�ݖ݆�&�b��
�wK��2N˂��[�/o{�$,���q�e��$�b;t�M�̱8R�,�f�kygW��,��'Y��EY=�:ez�|7z����t�ڟi�D�um�L�5{��N��K�_������x�<E��t�6������o����=�8	Y"ĝ����"����ޝXˬ�r����g*����FuQp���Y�ss7����WR ��)K�y�ٹW��Y��8���ㇳ�"�LU����ٽy��tGoty%BѕB7'n��4歮}33��Б|��KQqL=q�=7Y�;9m/:�n!�{Cr
OB5�O%�JJ�♃k�{-��,=��g��ѽ�<�x+�0�Ʉk��=В���-�>�J���&4J�L��l���9�����
�)m	�u��/{��XF�@�͊�0qֳ{���d�dwW�mH!!�,�#V��煎����������x������{���w�����{���w�������w�3�������MӿY��ڻ�yX�� �wWGWy��^|	���=�3��=��7+V���ȻI�6s�����{
�6ӝ���%�C�X��</�t�Z��f�d]�!�p`J�����*mr���p�K������e�V��Ƶv�t4B�;8T�w�n룴R`��#k7��jN:��fݭ�H�U-�q�z���M�uG]輎ޤn��z���TM%*�Te��M�AKl�٦h܉�c&��P���_F��ȳ���C�6���u�u�(�*�[��v�ϾH�]G4��r�N��%�R^Ϯօ��vN��Z�Z�7E��r��ozc��Y�.k�f�\ۇ��&ge�[�;O�י�.���`�T���ܕ���F����Yjg��ʆ�p�]��޽���Viś����b���#��އ�V9�[Um�bs0SU��������Ʈov�4���F�L���Gwsn7����{|gW\�Ŭ����8h�M�e6�!u�X���z^73����Os3l��fWeM|F۪Za���+��薱�؜��h��	�۴Eom+���͞NL�j���"�3s�����w'
Yyu��yv��Ŏ����ng Da�猊�\;Z���v'[�b���V��5�+�n�k����]N�;Y������Qݧʜ���] j��� �N��x����1Y��Y����X�lHc1Y�@����.�n'�4o&�y�Km��L���M��ٷ:0�d,�ڼ��8�r�QB�ڪH�ee�Ԉ#B{�W{7u�n�K�,��6���W4뻛GO=�$�1/��i��pb>���N0c���BX�^�f$�)O7�h7�����'�;�J��]خ��(�Si�v�gQVF�{ug:fM࢕��Ѽ%3rݮP����
7a#]��F���Tb��3�Q�\�M����6���m�ӗ9,�o�}�l_^��RR�x��&�ůo�y_]���!xu����2s��k�S�4)Y̔���50Q����:Q4*�v�H}{��V��p5!kk�ܫ.&�������j0�	Ip*
#n��t&B5lÄ%f^���-��(ī�U��=��Z���,o2�V��>�n�+)�ǣ)oCq��b�YS�b�"s"b�`��mA�e<�u��Iwv��(j|�V�p9����]َ����*�U�>l>���icYyGE3M��zCe�֎���6�+_
��Uj�;<��Y��=����m�Ԙ��'Fګ�vj#��T���)z��7�;GI�fr���)kb�W�ʞmj���10�z�-���B�]o�\�����^����8�MJ˃���+1
ea�6�'Y� ���{�3�z����i�۽<5ͷ�Ϩ�b��H(g��*�ڃ[n�UI���A�X�ڽ�$�$�Q�J�z�;S��`�V����UGm@h�b:8�ݺb�(��D�k��WN�v�뻣�JM$��i�5ݦ�(�Vإ4�4fmlX�&�v�ۮb(
*��z�Ez�յV��jm�i-�aq1I���L�U��Z��l[�&�E#Z�m��v4v)�Q��cDTUj�lX3:��`��ќl����f.�t���5-��[j4i�j6�Zĕ�d��#mM�Z֝0E�[�.��y=G�m��&ձ�;�b�P��bhֶv��������>*����nu��h�SiF"nF�!I)�:�q��|�*V������KFco�x�Vu�w�:�.�̍�|�<�L��gw1�6�	J�,w�l�99-�Ǵ0�A""�6YL�e`B"E��mD��DIE�T,D�
�Kʏ��\��Ts�.���;2@�ͣ�iB��s_���^��ukR��A���`>z
Ղ"�6��U�j��z��x���ڵ�jYT8���K�B��,+q��h��T���R*0�tCN
��U�]ݞh�1�����]�o��S`;��~��Y"+���n+o�����Bvv�\e�4:Ϲ�ew)�x솭gf�o��dE���gUng>tfث����+�gg��y�0`��W��e��ywc�nAw=(��i���'�LTz�����^`hJ��ītoe�]n��ݠ�z��n���t���=�)N�?H�g��u?$�+$��D�1�:V�5�1���owyZ9�+)O��9��qc�Bި]?LvS����̹�Yü������y�f�C+���IRG6�Z����eR)��c��h�ƚ������SUA�:����PE>�����ex���8�nS��7�3*rb32��At�5��oiE���r�;��������2�}ʾ��悔s�|E�r�����fDѪ5��r�C�*t�f��ľ��p�ҝ[�i-	�1����ɼ�� u%-��m:k�e�wM��r�&/	L��'35Iڟ�
�˲�r��Q#�TP��@��p�R���P+B2�$eT����aw8�q�����ݮ:n�ܭԊ�q �r*D0*oG���#�Wu�6�c��&�������ϴ�E���s
��. d�y�(��bĕű:�h�ܞ��i�Ě��n<F��ǗQ6C�1���!p�-n���`^J��������o ��<�Tב��-�\�>�#���n7����grT3ѱvN�M#R�F)�ɞ��=kcz��(���V4p�����t�}��Q�k�ۘ��GB4�(�'=(�A��Jv��`�P<T�{�L���&���c�c"�;g$���#7��
3���2���Q}["+��􋩭��Ш�f�%�-쑻#'h6�~a^�o� n<��h@Yg|�-L�[��E4F���ޝ���eh&:Nّ���tǄ�c��l^�~��*��Ι�dJ���M/
�ΚS�$O�ӽb�Gf'<t"�z�n��w}�%�I
����>�e�{Hd�9�܋ou�Tɳn\ݔ�w5Wb�^��:"�ORp�{�q7aL�7��22�ˡg2�ӂ��):b-^Z�Z���m�o�u��;�$�x�>�"n=VS��d�Cv�G}H��G�ot�&����2�=ĉ�S�4�r�Dź��|�*�+��w���H)��s�5uC3#�Ȏ�_d�BB\�iV���wkV�㍂װ/}�;�;��̞x�7ŴFE�ԖU�����ݩ��>I��eC'�����v�U�Y�A]X���@���긙VZ�?V�򧍽[
�>��}��ّ̗V+~����Q�0��45wj/�w�m�qנ�n��ڊ�+��I.�䚯>Z��uٙ��4ۺ�Ս<�]��9��9�� m�n�F�ܒV�*J&|�;-T��g��T)9Mͱ�خ�a� p�X�X�6�B�/��\���Թyg�aO�؈�o4s*����J�%�}�Ia.4�u��!ut&`ʎ�ժ�qtJ�K�oD��`��������v�2Q�K�K��v�H���"=�R�_M+��z�� �;�[F1(�ݸ�xB�XC�[7<ıX�������ʍ��U�M)1M����^���ގ�/B�1r�ԛ��N(��v.�:�U��n��#[K^�ѽ����>ߘw�%�oW�
��I{k�|�f��G�|Y�i�oޏ��)�[��xt�|�Fl0��y�S1؋�*蹫�/Ή^ZTqI͡�D*�m.Y��mG<�qҡȎ��0�w.ʲyJ������:�U�Q�'���y�>�8h�c����GK�������!'�x�z�°e�h�$�y��P�cׅJ�x�Ǚ�U�3�/ѵ*�} <*5�^�Gp�̶���#�^>C@C�.�}��v�<O+,E��Мb_&�pO��0�ڹ1�_P�ӧs1 �N�U��S񘺪��(��]�����见��C�<�Mw�c�����Ȋ�9Y�il�ι���|A�%%�ה��s;,���PFB��Y&�3�{��܍����W:��}�+�$�ѕP�ώݿ0��y��^2 ���{��9���b3X�b��f����Y����	_?���
ն7u�.�7��3�n%q�|��ss[c7��=�*u�f�ba��Ro2���!}3e�6m��C�uBE2��V�^���`�!�3eB�����;���l�
,->�C���������p��Y7x��).s7(Y��kP����6��߃���]��#Ύ��P��*p�v�������d�:vڈ�g�H�D�@��#�RV�Tɳ��ow.ӑz*���ݵ�M��Ԟ��k�2��*��'����)�/۞J����
Er��ݵ��o����G�����g�~��� �9>�J�S�� ���2L�:�(ַ���U0ݱY���&$a��i�7j3��WC�<��p�t��wh��g������q�QGVUx�bP�1 �mv��q�s��C��[��F�'�)'9���j���⑳=>����+�$MJ����m�v'�s���O.܉�ڷ���x���u�j�y}':�>,�ܧk��v�yc3O��Σ�s��a��4E�>�\��΂1��.���t��7�v�D�kU�Vj���{���S�-vz��6+��1�f��ƥ~���oc��$I������"v�ݸ�c=��b�O��6��N�>�������
{z|�����u��k�טX���ɭ�P����kT
��B����Y[�rPL',�3��!�V�7x�yvy��F.AR�&�A�ca�)lT,q��(4.m6d3��bn��v�4�lG?>��;���i��F}�O��H;�]�vIbS�
>R(F�S6��pM���w۸�ZO�ޤ9sVRח62YŎ�� �3�ol�p�욉R���H`�C�q����f��^���%-��������ۜ��/�	c�̃6ME�j���%4��'������r���=�D��A���(L&�`{Z5��y��s=�[z��Y;^l�Lj�}v������3dEG8NE:+����)�[7Zw�O��h��v]ws�8�6��&��TIUy����H���t�?���;0&kc�Q���]��aj�iWL�V���28��=�!�{�a3���I4���/���>�
�~Co��*Q��������[���Q1�6)8�l�{���$UG��O�L���Ӵ;���i)��p��
����ϙz?����Z=K���7�m����X�]��W���	�-1�M��LĘ�&V�.eU*�c��)�G�T�3��>5�����E	���p���P<D^����@�J<�������
�2��:�.�'r����0����K#��Q ��d�̋�=��}𰾀ú<�q���Fɮ��s��ڗX<껨����iZp�/7y.U�T��y��f��`�|��)tq�*��1�=��݆SkL��:�Wb������:wb'��E^U����};8s�4���Lt�� u	�&�9=x3�w�[�����*�v�UB����:�3���A ��%���1����҇=F����+El<�6*ʽ��_�|H҈��h�ҩt����W����%�P�
�Fz��vU��|s#։W� �@����k���S�5���G��*�?h�S����Ne=��`�^��c)k}h@�T�i�XM�����*Ux�Ɠ��}��vӿ8�;����y�b1�YL�^�}r�=&� ��'��q�U��3�0����{�*?�����S�."/c�I�-�����F~TT�_n�$M��
�Q��� ~��"aΝ���72��nc7�)�7�m�%l��E
���R�ƺV[�2U���3��&ff�@9����w��j5���Nt�)YUQ�Lӊi5Zު�wV�V�z�c��ޅ�^�{g�*"��;��S��u ���c�k����1�Ξn�)�
=Z�����rIXn�%-��2��Yݣ'���os[�wBA�'���U��pV.��j���P���Fi�7&�.of�;w�8#���atz��WbUGF����3�hDjl�4l�����>��F�P���&<���yU޷}ǁ�c76���[�˿ӄ�go���}��_�+��S���ف�U}0��y�k0�15C��yݻ��[�ɴ:՛�{�Z���6GT��}*�nV�ڪ9z�x�YX�ל�C�0��.�wiD��q��Y�2��{M�A����*���uzZs;��-�A�,נq�v.Z&�L� �r|L3+�v��N5ԛ�ǚӲ2qS��_�������F�o/��H�̶����7�E�ju.��>�-���U�m��OL0����L�HI��n��gu� zI�����]=uEIF��eF���hneIM�nV
&�#��_y���f�o��76�2$��_k�Δ��G�`���fY{��HUu`��;�+t>xE#�vٝ��	������ݶ�G�($�\m�����S���0A�^C�S�ں�ܛ2��k!Ukڗe&��>���վ�u������-�绒A��!K�����^�6oV���Ǌ��()��HK������Z���*��B�Qx��*:�k�_b4#";PW@�dQ�4 ����
�rB����p_�e�ʃ}���} 0y�C��[$1<�dn*A�'�y'D��V��[��F���^�E�Lc�L��H��p"���#�RV�M���������稤֧k��/d��'pu�s������]RGG[(e�=���/������wm�bCU$�7J�V�'���jA{��ՙ���b��F�ܽm�Y�����x���D����}�cݬ�cDLl3�y�셣J������:��W���,�'r$�N��������x�{+���%A���Y�W������-N�S��	�F���*��̥-�� �!��R;M�X2�b�^��1VK�MLL��3[f��H��gK���)�o��W� ]*�aQv�wd�lk�Q������G�]A�v\eL��N�2���F�͵��\�1���^���W} lm�互&�M��2"٘�6���3]U�s	�j}^�6�p�P�E�]��/�#���y�Z��VM�oM^��GQ���At���&p6قx!�����2����,gX\h�����݃�O���ѳ��q�:�8�gC�`<+5
ϼ|Ӽ��Z���R��Wp�Ψ=��r"A ƞn�&�)�FC8A�!\��eA5��zsv�g$	��o�z�o܄E� ����eb�g�e)ا22[^ݥL�t���EnO���30�#��+J���3@)�wKBG6��74�e�pm�!��\�_+��G�c����v�ѯE�O���AM'��o.a��NP��1 @��Y�e���9��>&����#���B:�u'�R�!�l��U�^͐��q?�׽���9�w�5W�"���
�)b�^� �/���z}~�//w���{���w����{�����{�ޞ�����;f�[q��Ϣ�M���g��Ϊ�OLwY;S�{@ģ�[����x�0vI�m��53x�X��p\�䆧�R��#��,
��'WĐ�B�vG�ž��<�uy�Pv<�wY:KZ"8J8[�h�vq)�F�3��Jou��gY��EF��-9~�gjښf���m��Y9��v�G}7[O�G�A�\8UL�	�day���I�Ckf�����m�֯)�Àa���p�������wq5�&���	�3�N]5.?Un6�uf����=���5�' ^vE�n�˔vOK5�֮a��6��wVpWo7^6�u����óhd�E<A��Ӫ����I�C"3rpUqI���l�b�J.���z֦:g�u6;/�R�Z��J��]�V�w+{E���ٳ]z��h�Y�@�J�b���PA,]geE����$4���`t�I�w_\��Q��X�G�&�]�v�T��;���u�u4�ew:�B�c�:V4�q�i�)3F��:��,��&�a��h�b0hҹT2�*ۊȨ9��z(���n�۪oBf�`���Ѣa��3�4�P���3z��^��F�R*��cT[ȑ��v���l�,[l��7&�R������(��:�P��7:�����a>�C&��>�_/5Y��Y��N��Vtp�,�&�u��K5P{i��:[��mg}2�p{�f1Rn�ͥ�ѳ�Lq]���k2���B�!��e�"��(�;ӻM�*��0�x"�BUm�f�����{Na(������ cHp=�J�2���:�K�|�z���*m��A�c�h���vm�Zg:�u��.u��ڗ��ʜ䧦�&��kP2Д-��;d�Ѵ�8I���o5�-��8��ˏ8��CI��`{�g9���{���s�5@� wS�*DW��r@쎶�w�M�v{����N�h��Qmk9���s����x�t�T�%�Zo0���ZMȊ����d>[U�8�n�Ȓ�8O[�M٫d��,��;Oe�e��r�9�����8�֪����B������Q��"�X�c�{ ��z,��e��v�wo��9v��]Z2l�=�(�Sw\��\d�7-��a�9����Avɻ�J7Cl:/qX�`��W��b���Q+�AN�nT�'�]k��@�mXx�M��e4ULk���*�z���|����?XXjM�l�$"�w�g]d� �-p �EG�#(`�zٕ�9c�T�lu�vF9�5+�mju�p���Lڄ�!1b�iU[KQݻ�-v��ow_N+5��݅�0]o�]�浼S�c�Yy����D-���}�9=׬�F�a�������s0-���T�r�p�؁ʛ׼�	�q�ˍx��T��ns6�spe�d�n�K��R^�GtFdOs{�����$���CT�Y��æ��QL�F�}r�9\ȧѭ�)����N�}�=��z�bΓ��U��wϮ�X�6�\i��vΌm�bj�[�wv����������tX����7w�VɋF����4DGl�]��Ng�5Ӡ)�;e�����D�l骢�;��j�j{����f5������ɱ���bz�5Q��)v�Pk��g�ਸ਼-�C���݌kQC�*�R���K�c]8�;j�:�l;o���ֺ�;h�5�.�5����ާ��]����z�
/X���'W5���t�Z"��Z�i+Zě՞�+8�����Q��i�h5v8��^�]��gV�RS�F��h0M&�[k�&-��z�]����z�]�EU���B�0��H����֧�K߯;�%x��{�z�2�j�;���n-�L��U��+�����9w�h�Ӄ˭�y+��������="6�i7)9dF���q���'�U��=뎺u:`�HL��إ�0��Nv�Õ�0�����.4dϸ��&̆�x�%�F�����ؑQs5		�w!V���^6�SH�yr�3���m(�f��ٖ
�����ؕ�#� (^��M��{�J�����p�.+.nӭ���ǭ���G�'"+�L]*���x9�ʺ�u_21�xn�6�� �e/อi�7�=P�F��~�3���f�ħ���� e�X�����}��gsy�j��7�,�U���;��1ۍʺ��������ٞ�=^/��ă��a�3�1�h��Q�]�3V2�o?0k���ҵ+�p�9����3�q�IhELV��o,�"����}q5��c�DP[x�>ث&�����/$�$D{O2��T�~72c#r�Zww空m""���T9���|'Ր�\��a3!>馥I�!����t����\'q�>M�7�E�w�ݣ8�Q�;�B��fXT�I���A�gg$��ެ�u����Ӕ�t��[e���Ћ)��A���ͬ����,�Q��oX0�v�WU��-:�|A�S��9�⪺��<f���t��}YW�5c�Ył2=��f[ʽ������1�u�2�鞮���#�}EJ�$q����3��ň0�=_!��Zڦ��sٵ٩G#-�+%��hA�U�ٓ�xL��e1a�N��j��g���"{A}�RHK�H�$�>ZܧY0��,Zm�:��+-vw2D(�.1`��#o�]#��$��QD��܊��Xϳ�q��
�pӎ@n�S���.�mi�������0j+B�D���SEuݿ^�v���2=�1�	 VO��]0�+��v%\i�2�fo�k.����콄4�4Ot�-[�b��̷x�a��oW�]Tr+�w�0hC׍�h�oOA�9���}��4n�7���-���6����"���?��f�R�ɹ�om!�:I���eR������	�&��Ye<(y��]��o�x��� ��>�[�E�p}���-�me�<�J�֪�>٪�\��<���B�z�Vʛhl���`��)GQ�j��lwݱ˺�*}��o�;:c��}ôn�ݧv�c>�?_O�*0rA�[@��Vq��ݠo�j���uY��\��pL�N�:������^�H�~��ђ;�dv�;<�!֥c���VY�{�$46�g#��C��q�=v.Z&�2I�%����:i�m�gai<��5{bWG(�����ޟsp�̏[�0���[;�CvgOgf�)y��E7�b_����Bͼ�`֕�Y��)��l������SE�'��_���؝<�omO�E<�qC� A"q�d3����l}t��m���{��U	��k�Y�s l��^���ڦ4�V����pGH��hFGi
�$W�N�g��w=Ys*d�����R�OJ�2�"��2v����MG�Ǣ��܂��J$�J����t<TNY�ٝ��9���14�ZDfBx�z�F� ������6)h��*,>L�H��`����?�A���;5>g0���[�W�`oiKټ�*�i�����F�{��t�S=�����xْ"����RQ���h(t�6����xhĢ�)��+����`��q�eM��c%cC�t�ܘ�٭E.sԵ��y��q'��t���B�C8.�:+c��U���ʮ7
��q(�I��'���V	�U�J�]�������|��P7�<0Mɨ
'�"rn��N���4ʠ+�J�PzN��D�ԛ����
&$p�{B��n���3Y|�ۆ�Q�� ��6�|i�ֳi�Z�v{l���/�c�B���w�Tv�rߗ%�&��L��MCP�{kz+p���2����o9�Xb^Y#r7mt-�Ϟ&�T����:k��)��G�7�P�3h�����A}��]��ئ�g�#\��>��v�1�]���!�k��;�"Ψ���c5��������\I��V�*��~�F�A�4�v	7�O�c%�k��.�������f�oh�.����:m��7x��9sYJF�?Ug���}�~b�zm��B�;Kk�Xӥ빺v5�/����E)j'1��`�Z�e�(o���
I�ˢ��w��!�N�b���a3�=+��,sg���`���ySd|��Y���7�S���km9�Wp���Y��t���{Sp���0�i���O��_�Q��?zgp��N�V�@Ґ�\�q�J[䎲d��&;^�9��]�|z�c��PW�T=�ϔ�5>�B�PTӺ({+���;E4�2��}��c}�lD�*��Nxb�	�ֵ�g+�4�=M��W۽]ݛcRIT
2���1��n�U��.�
tVC�ȢOgv�ݕ��o?[���gY�M�&�*�IO��*���W_J����Q����ۼX�z�"��;|���EA�q�M�lǔ�*2C �c�n+�λ������ �oO���Z���T�F�+��To�ѧhJ�[�"���q�m���6G�t;X��[�����3ֶ��U�i�c�Nm�k^n���Y���2ڬ��Z�q��S�]C����∺��-u��x̝�� i�3F��͖3�f���ǵ���{��[=IkX��m�a�4�҇&DZ�WN�����i�S|ٌ�rC���b��w��g��wdf΍��[)!Ӆ��u�TKra!y`�,���F��Y���ٴ��6[��4��C���ۣ�,A�y�J.���{K&�r
׳C5c;����:�%��(�V���G��ݸ�T�A��*����8.P�1�C9�bv+��ۍ=�r �k'ð�-���vA1��3��CXu��b���QqQ�ums�>�N�Ք.Wr��8���#��2	- �J���j+�,��yu���������F�
�Y�乓�-���w�Ț��\�u�7�w1��p�G�ϵ5��F�	У`=�5WU����`�x��#�x�'�����r-��.΋m�}�:�^��w;x��S�g�S��C�S\������9ᚨ��W�+}+�Y�z�Q.�u�Wa�!����yU{S;�{݊vp�X5XUF���(��^yU̟t�Ŀ�̤��̾<���;�/�f0��,m��6����%A"�9&�)?oR��N<o��mʫ�9��������le)#\�:ѷ�7`�a���V�*��6�'�?:K����J�� U�gY�X^5�P�+|�%u�
�!8�L�X��9J A�[92��`�Sƨ��z�7���C��2&�����kK����3{M`���<4%��]���gn��a�j��50�h#��4Bڊ�,�A�Ì9n��SroS�Յv�����$�U�S����ٓ�WV�1Дb����W�ދ���,�kq�����-�7���e�S���==��]�]ǝ�W�F>��n��g-q-X�^�p�}j{�B�*�]�+	eJ�[ 0�T��=�U�ֹ�+Sy[�f#�W��+�n���ύ�{���z#6"Z�tS�Ƙ��Ո�e�J��c�{$���{�)�'��b�Y���	����q|���H��]y[��C^�g���G:-���g�{��]�a�Tow�V�Pk\�����	]��A2q�4��2-b���[y²m�`��W���b�,�xTr+���f��)�*Q\Y�}M�s�T�&������p��=8X@�h~�� g�#�Y����VT��k�3�M��#3��R�g�q����ɬ��i�xna� g���l�/���s���^�[� �9M�9�Q�ǔ�:仓0��-*v�0��o'��}�s��vӎ|M�̼&Y8���	�^*N3+$�M��ouX�R`Ks`=)֠δ2��8���SS�a�d7����T�C�c2o�j�6j�9��N���n�tn����^�\\�Җ�A)R��[^R�\Ӟ6*jjƶd�I��F�3!]v��b4s��0��ĨF;W�k��+F�����5�N�h�[�u�\9��dS�*�����"5Yظr�Fi�[��g���9׼됂����F�t�W�����FW�����@�Z�����m���������[7ܯ��*��t�ӭ�TEmzx#G���[Amh��u��/7�[��c�FW�H�� wWHb�O�ǘ��(cdZ���Pu����!+�hʠq<x��='W��I�V��ƶ��!NM\]¼�����W����L���ՔJ1�^�wd]�6�"�T�,~ȵݺ��C��.�3�-�̭}��w%�&���e��`���]���a��:df7�B��!�q����p6�m�\�O�ɂ6"GF�8�,����nBV�3�Q:X�q�&Vu������Q�
����'�i��Q�(��e��qO�&D˰�I=�5�R����>�ԁ�&a㍃N���׼7�*��f��\���E�[t��K&�!�i�e�5)���l)�;2��דOn֕U�S:݆S~��H�(x��������E���W��h�n�&�9�o�{�߆���_�}�;'�Ѳh��C]�|;�4F��2��zVk�e�-\Ь�I�g|'��Xi��(��?H�>{R�j�"�m�*'5���T<W:�~M��7x�-�E�VR��v�["�Y�zb*��a{a�. j�j'���si􂣅r��IB�5Hs�x�MJ�r8�(��s'��{��Ȍ�mF�u@?T�	{|�H,V^����UC6�k�p1�ݼ(�#��Q�ɹ�3�U�r+�//0����Վ�➼O����I#��fA۽>W��h@NE�qmQiUỜ�ͻ޻��f�og�J#���T�UO����y�71T���99��K��/\���9�JV�m�<yux�(��<s'��mXY�;v.(i�_���܉Z�
Lw4�ұ
)��X��fv��p
��Q�1����K7���Sѵ]�wK,Q)۬���Y*(0�Y:���v���Z�F'�ܗ�tѪ�IF�h۠���UL\crж�	)�Rsk+T��#�]�')q]�����;_�w�aH�O�J�ei^e��u��*K�)��ȓ���ޕ ��-�[F��==]� ��Z��e��m�s3o��y��O�l�ވ^3\&��C6.k����9]��Ȟ����K9ͭ��x��L�4��d�i�z�F��{�f�ʰ.���Ua!ߞ�o�l������=�}m;��3d6��o�8��������M�S���_B+�l��o��@��_��1�/l�5)XT��U���W��z�Z�#!��q��w��7��ңR������ꢙ�􌞊:�#�D]�'���=�(�h�΍lU����[�G�ߺ���+���)��=4����΍�b��h�M]Vfp+������	��[�9�����"A��rg�y�� ���N������?��k���O� x�{���AP_���� ��T_�P�G��|����
d%�fE�d�f�V``V`Y��`Lȳ̣02,³�J�"�0,�3
�2�����ȳ(̋0,��̋2�ȳ���̫2,��*̣0���(�*� L0,ȳ̋0,�� �L L�2,��(�#2,�3(̋L L�0,ȳ�2��"̫�3"�0,ȳ̣2,ȳ(���"�0,��(�+0,��"þ>Ѐ��dY�f�`Y�f� �FdX`I�f�dY�f�e�fU��X2�³(�0,��"�2�2!2�ȳ(̋0,��̋0,�0��ȳ�0��3�0,�2,��(̋2,�3�#0,ʳ"�(̣0,ȳ�0,ʳ"�2�0ȳ"̣0,���3̋2�200�2
�>��(�*!(!�! !������|ʜ����ʪ��ܞ�r��ʪ�  C
�� � ��2����  UXd ` eUa�U� �UVU_Xz@ �  �UVUXeUa� ��K�a�a�a�a�a�a�a�a�a�{C�0,0,0,22,0,0,0,0,:0���̫2,�� �0��_1�|}A����*$�  Ҁ(Q�}���?����o��g����~����9��|�?���z`瓧�����k��$W��������������!W�_���@�?�?��������@��?�y���$;�?ޟA�_������?� �v+�0�*
@��@*�D*�J�"�@H(�( !@ !"* B,"�(�( ! ���J� ! B����) �C�I
 I�A" D  I" 蒈�� ���Ǐڟ�*
�Р�@�P �%���7�����0����`z����?������������������=$~�=�#��o�O����  *�؇���=�����C�������D����=�����O����_��������=��4��1�o�?���؇��gǡW��=��;��>�������q���߰��� ��O� � ��H@@U�}��#��X����������}!��}~��������?w�������}~��W�>B��~�ޙ��?_���k�r{�5QW�����TD��_�}�_�� �~����d�Mg��5��wf�A@��̟\�o|��$�EB�%QR��EJ�THJ��J�D�
�E"*HPRT)�
��U*���BH�Q�T���)UR�! (�T!D�"���"�
B�QT�J���mD��EAU
6ФTP��@�!QBB�"�3�J@TQ �EJ����(�%)Q��*BRH�RUP�����$���	URT�T��BEQ)J�U"��R�D�D�  ,�v؛���8WNk�eJՔ���-UX��ٻf�#����`u���Zv)����A�X�n�T�;��+m+P�[[���]Y�UJH"���E	R^   هC�ЪP�Clhnz7C�clhhi�^�C����Ѷ�s�p�z�S��K6Uj��AݤNE�[f�`A�Z���*�Jj�W3;���gN�bw*�SN�JP��J"*���"x  3�o[�*�wsb�vi��M�h�v��ݦ��1��V��c �ۦ��%uݺ�*��U��4�Y�V�ۖ�-�q��
V�,�tk�:��t�AP%� ْ$ �   &;ֺ92�[�wm��]����vn�+��%���)�k��sN��.�-��Z��vgfw;��V�j�U0U]0�H��)D�A �Q/   ꧦ���e��vr`Ӑ�]Z[�1l��;C�Q]���T(C(�@�cF�Kmk���Q!HUE*!UBJ��  �Pz�%��:�cQB���kU])Lt������5��G[�(WTk�:��jW*ݰ-e+�p��5F9(�R�	JEH�(�  �*JZ�(=QvbՍ�jp�r�� Z&�� �ٸ:� �,�
�X �Υ�h tw;i)J�BP�)UI�  ��  �� ���:h���  Z+  ��s р 4C: �n 
 ̖  :pp$(��	IIO   3� �Z��=��� 4[�� 
v�W@:`��a�P�m�w]n� �k��m��` k�\�*���$�UH�H   Z�� 7C���0����: �`M:��@��'p  �` 5���à�u�VP <���U*��h�B)�IIJ� �T���Q��  �~%)Tz   ��*J�4 2�JD2�@ 4�i5R4q<V���r�$ ��,H"�^daE@[s�}Vrɝ��3�x ���������L co݀6���1��~ 1�����8�m�6?��~|�����������x]b!�Y��{&��Aջ�R�'�k5����]"Ό�՜���:q�̊��]<��N=�S,�r`nȉ� � �SL��Z���n`Z��,��2,��QHT��C��V��wK�V�^���X�"mٶ�!�V��Ф7m�� Hf�(��6��ä�3`uq5t0�b�z�&��[E&q27pxƯ-��E�M�0EQ	K��f��f����2�N�P.� ە����g�luj�W.���^6K�eQQ�̳��]�F�Xl�c	�U����m��k4�ݘ���R�gʷ�[��2�LD<h��T��.��H+�qˑ��^EZ�7�p���fcbmRn+�ƲVsj8�+q�ŗ��IZ*�ƌ��E�E�����rI��3dJ;ⵋU`�d���0Dj�Ѣ�KU5��C�(2���{{(�WV���lV*�J��Y�tKljn1��Բ��[ze�$*��dظULH�=�%�2�ε�ѧ[��?��W�X*�#]P��c-�f��n��t^����ݤ�)+�aA��&���{�ˁ�e��2�kn���c�y��of���Gv��48���ٶ�E�yb��t�����ӺX��dҷ.��)��,VY.��Jm ��-�cv�Q��)�[d�d(2�S��^��'Hc�T��L ){��X)�0i���jL!df]�&q��N�z� �P݋c� ښ����� �9ML�ؼ�(Ы��I�Ena��v]��q� ��D�jX��d7M̠
+5�YYPj.�ں-��M�*���I6�ʲ
�C�]d�N�։j�9�C�iG"ub���������L�/X7�Y�в�9)Z��%�Kf�O-K���C1з��E<�h;��o��9b����Ep�Xioݢ;@({�)Ć�N�[��j���������;���j��T�����["����X��n�8+
d ,*��
�\R^���ad��Y��*Ul̋��uJӌIy�°1�`���{��J��m*nԽ�s,�hݹ2��m����i��B�$��B��X�E�X��vS�Ỽ@n+K8b�El���j�׸eL�*^�3[C5�U0 �hmG�1@Bb[
�^^(�QO��9�tX7rua�kV�e�tܽ�&�:�%��W�������Ma��ŭ���np��^"�?X�1	�٩n7��u!l�� �顆�B[ܙ�kQ�Բ���&��3M���\����$ݻ~�5��Vuf-Z�]n�:)�=�y�[L=�P��vaT��@SM��ɵw�{�طߡA�b��,���eF�Fި�\�wD����z~�1��j<f�ù�����(�Vfi�Z�vm�
J��0�5�i��1nTJ=�嗂h����I��>�&Щ��k��{D��*@��gB�+C��,[1Va��Z�&����4�#n�ʘR�0ɻ�-�{Y�[$U��6�e�T�P�.��7j�0�M�"ƛ5���ů�:�jk G7Pt.!��l��ygG؄�NNz0J�ٔ�<�
\�-Yh�LI+���i f�t�`Q�k�g�
�]�j��;�6!�K�Y�KV,l*�R����r���9�[<���eV����S�Z�hn����P�b���H���f�(�0j�U�ko
:�˛�) �L�x᫬�e�>�ѭ���0���зGtCcf6���ZtoZ]յ��J���ێ��r�+u�M�fǎ�-'{�øݚ����#�KH�b�3Z�)��-i��}�Ad 	�1�ʳ�t6h�����+bi�Х�2Su`�(]0FU���7�����Ĩ�5�3	7V���fH�i嬪ؕ�Y� Y�j܁�)R������n)mLق��u�.��6M�t���H�0Ue�QjA9[�s ��O!��lӢ4H��%֚�.��΍�R��N�st޸�_���f5�!MYc隥����%��{V�x�8�Ս�4�=�7V}H=9�[Z~bĽ�V����ͼ��U�ݚ�G$�weU��3	1,�
���5*�
Ѕ��5��86�"n������&�����t��������L� �-�7q��th��X��i⼩V-YP�6��# �QT��@ (l(�w�*l��\r+8�L\9b�v��J��jM��g9��Uܞɶ�;��Â`u���ݚp������a���P*�f� ѣj�X��$ r;VE�;� ՛�U�*�b�Gtc�11n7#��T��
`���e�ǻyE����)ՐhV����h�aFʥ��"�Kr��sV��wZ�xW���O[�#����Z��ɹt��7[T�q`��B�m�y����3��n�����дt"�,	��J�&�ÆV�(�8�2��T�'��wa���!gj#�`�IRy{7& ��A�1c��{f� ��2|��e<[��hbtD��yZ�����O㗙m^Sh��~X	%XW�.�$��wEd>*���	�*R�]�� Jܦ��W�2Ί�r���/6 ��6�R�[�����]ټ,8+V%��K��ʴ�Q��R#u}$��W{j��tV
���f�YջtV��ԐEQ��ҩDf��v��;�:���m��)+)sv �f ��L�h��s7��\��,��P�F��㆐(DV��<O���3�^�k+#v($�D�5���,�3�Z�2�yе�d_��wk��N[���i�U��в�al��J���9��B	O4�CYkE+hh���ܶptD|����t�q�H�6����}t��*���t��	�Tmm4]+ƤMV���[Ae#M,�8J��j���"pV�Ô�^����񖤒
Csb��ڄJ��RB5T��-�Nn��C+!���`�C>�w@n��(���,�u�l	1�Ѓn��u,F�v���?�t�W�/#%T�Kw,+I��Kn�*��k��-:�*+q��k�CS �QU����ո��[Vβ&��`�ӛ��l9�U4�LN�-[iF�[�6LT�r��ڂQ��T�e���������z��ۗ��Hi�DH�Zi�a��*G�B�m#����C!Vb�6�]�c�2��e�2�����gg�ߍ+ܡb��H�MF������	����뫤4�^!tu���J�8n�t�|��S2!G �B�	S0���V��]`hm]�	�X�2B[���&XX>p�o@�ɕm�W���#�5q��ָ�m�*X��9c2��e�n����Ll��Or��A�\(iCM"��sfs�@��b�����Y�i��â��ֆN�	xw��䥉b�m<�4=N��1\AH4�ӵj��D����)������k���T���t<ӓq��]2�ڎ�[���7T�%�B�_��#�q�X�MAw��x�5ӌ3�)	:�"�T�l��4��Ψ�1[t&�ح�a[U�KL�[���y�՝��
�:l` N,F`y���"Xp�P���b��Ĳ�B�B���Sm�
<���TR��)�*�[���c�T�	hh˷t�56�.���CY .`��m�9v����B�O@e����Rf�(j�'��`w�f��'� ���2n-�\Ҩ,���ٚ�[H]:�cЦ`�PnJf���U�Qܶ�$�Pˉ�4�#.��fPum#	� �k.Ļ��u���0�ݖ�i)^IM',�˛B��V6E�D�z�	.��3�7/p���Q�a��5�7�+Q�An���ݣ���mww�&sB��Y��v�4Hxih"V���ed�����J5��L�Z����6�n���N���,f�M6��!&M�����A(�I���9��4�`�&HMִA��ѕ���K% kNd�� Y�+jf����VqZ1�%�hF$%��ۦ�/R��Ӥ軂�	7
������bG������C�YGf����0�2�L����:��(:t-�f��$�Y��ݫ�'�c��vݤem��mlX���$�2�9�&U�m�f������� �L@�
,-�	�J��^:���(Ym*ӵw��oh�{R�Y�	f^��>C�.�{W5��{h� YM.�G��D��j���gC�Wd�R��0D�^̺965��l]M(�q;{����M�͒�X��\�R׸V�r�jWJ�յ�1n�)n1���`c{cpI��qe���wNJx�o�D�g��ƌB
^
YQ䘀V�)�̅nSƬTˬF�4n
dZ�j7�̠��F�
ˊE�QR����m��b(6��F;��ԩ��x\d������&)�L��ub+��X�*��$��n��
V���@�/r(�f<"��
�R�.fL�[)f�5�i��	P��F@6��U�%���PM�f�� ����t"P�j��0<"�Y��bUz(�ɁY���1��)���-�fJۥa�HV�f�@��-��ZF���4�
��S�k(��DZ͋�qFq�`9AV�2���9M���SڸjMe ��t�W{�R�
�;�K���V҄�2弫h�Vav2�n�L3>E���ɛ(5��?��$�T��2�Y������Ǜ�Q��u
��u6S'�3ш��lұQ�f=���n�����M˭YT�ш�y��-�]�4K�m��"�eS�U{�\]nޢ�HÃ$��I�5 �[��Q!BK�&������%���e���;5�c)K�����ތ��ng�^xr�=	r�e,e7��zi���]dj�LK°ʉ��1B(R�>yZ��2妴d�Z�3Fj���z�m��@-y���\�ɸ(퓎�:%�Y�-m�X�h���mj�ע�g�X;4�J�|�g*� ����������P���i0�sF3��k&�UL�K�X�{Hj�Y��O"yx ���Q:�ʰ�̒:�BBm��3�EX�fC�g�޷V�ii^ �V�hMX� F���!�e��"<�D�ƲPv�v1��ݶ�Z<�AP��m	�2:$y{���B�2�����Uzf#��޿�0 �s
��uJ�n�y��b��A�̗@��EZ�h�z�S'�i�h�wF� U#X�L/36�<��Ք�EN<7�
�`r&"�:nZ*T
�xS�U�ѱ���ˍ�:ͱ*aݣ[��D^�Uь�1��#v8En��h�;�
:B�'b^�sr�!m�D����+Iת�Ŷ���4\j��-9�b��J{IL�V���F�Z�9Mu+FbC%ͫ[��-.�DI6�j�,��-�M[L�Б�X��D/.8�m�h��2$Rc2��f�j���0[�bˇ*1�k.�,�ʻSM��X����rU\���x��T�&���+i�*���*�|\h��Y�(�AQ%^�{��,�c�G魦泮�����nڣZY(��4�e�u�Myn�Ħ$�M��P_Y�>Kk4�b*T1�ty`�b�GrU����
�Ol^�.�R=��l�̎+��� &F��] "4(��F\�����PtZ#-��h���`J5u�IF���s�;�˽�V��kdj�SiG��<y�U�,'�6�A��˓F��(���;LPp�cMё�0جu��im�rVGPd{V�mÒ]!�b�]��E��V��6q���Ky��[	��u�s5�IV,;k&,�L#@2T�#�w]�7h�Y5ޜ�q�v'�Zd�I=si�	ڼ�]2F�D� 5�w�Xŧ&	ZP�κu�����i�U�kvC6c�vS2�	9Ln�ڄkN<ˈX�ǳZO,L9��ۉ�d�ܵn��mJ�7�%�򬇖ա��5��wXkt3\u2�����p�m�h;��`��Ɉ]�fuw��Y��hrk2&��2A��6�T�X )�p�`pH{�F��jδ.�|r��t�:�*�0Ţ�$U:j�=�6���2�DY���P��8���֞�AI��30jD�������i7)�nBcz�n}���Uʘ��'ڢFn[�SI��g& ���ͫ��*4�zckr��ۇ|*:Ğ7���M�f[[���̸["�*̗��Xҹ�S�D����2�R���c5He�WV�i!�f�2�l�iޛ0���������zuD$���,����H1���m텍�x�f�Ж�	Kwc幣i����ĝ����$�үY�Q�)��]�btĳ��Am���[�bXM�����������2C�3#��Z)X����I��z+u�:دxҙ�R��(��:`�	�e�Q�͉�
s�S�22*Uy�r^�[�^Ʋ�()Q��j���m��-*��n�KK&Ɖ��.:җA��L�	�A�+*e���4�!MT.���c
��gk%;�qQa��L�r���6X�9�#XRn���p��`.R�(&%9�ҳ*${:�>2V������7!M�����
�i��y���5[���k�m������@�z��A ��V
5�/c9�*%	�aYSBF��,6��++f��os�ۗZ4�dXX	+�w��[.�-&^B�<�m�on%2Z��-E�º�Y�a �:�dVbt褱�Fj��[Ca.%3k('`� �:{��;�P�t��Ƙ�j�Z�w��?G��^aӨF�ݶp��7Nλ�q�wi�GEFp�0�Jxg.��;�����K8�A�e��J����/�9l@ף;�v	�MI)��	
L96�
��fd�܂b bMS�)���me�5jV,�VJ�!���6�����ڔi�X�օYP�`�Tcq=Z��Qڰ 3n���d�҉,'x�=d��GB�!����wnE�;egMh[�w�E��y������Ch��;�ʎ�N��{V�Tw�@��;�4VL:��mt���άkq���7��B�����[��oV����jn}$��e����i��X#u���jI�*bn6"�,�y�+�����S�5r�z���u��P��v��N�cM�[�pS�@���DX͒t��ҧ����b�K�ɞd�<����t��;�e.8��ܺ�`���[ٔ[4�偁��Sh��
2���C�E�D}w;����8i��wt�y�_t��q<77��w��t��}-��c�Yu�{�X͝��dkYט^�M3��-����y<���ᏰVb�P&��z�=λU�Εh˖�l��q��Om�b�/v��n+H9�(��bו.a��ݛ}���U����S���Kz��f��Z1��s�bc���v��}VU��B����q��^&��T,P�, �_p%�sj����9\̒F9n�vJ���/�iLq_wU��x���ŏ6.ٍA�-I�|e��|k���Wvd-�S���@�ֺN5 �Uδ7X���	x�.s���թ·v��eI�a�׸1���W�!��y6`����K��)����i��6�l��86���x�+.d�.@��F[�w��J������1�-�[� ;��T�_r먌�[yƠ�Vy@�Eݶf+쏬^�Y͊b�v|�ހk�oc�#�9�wm�*r𨚧r��<� 1R��$s]�k���:T��B���e���Ƕ�R�&��KmΥ�Y�CC����2����g=�C ���J�Q�6�X�|gp���ew,�ugn�C�A`3r����0��:P^��r���B
�|[�ٜ�.��r��/`���:�FZ��\+[/43�:z����'����+}�þ��@�]�2W�Y]����Ř��������5�.��^�Xm�$�[ާ"�l־z�������C6&������bWNL�9�)����Z���� �l�L�f��4;vr�[t��F(� b��r������wk���Ί��ܧ�l�S�K5��:�.�><r�e�<��{n,�+qQ�^3:��cy �Bu�bs;�k�n�]�|+;{�մ8crގR�Tm�n7|i�ʙ��Ѷ��ՙwI�"�rU�V�Q���WZ�6��T-��"�K�{mp݋��Ⱦ: ��D��ƌ��
����c�i��rdWԩJM�:��.c��u9X��nU�{V�+k��eū2>\Cz�%��;��-��)Wrm\�uk�ַ"��V�Q�!�{�d-NgV��2Z�Fu�{�]�"i��΢��6\˕{uw�]v���.h�u:� �:2;�ц��μ��屍���1"������Y)�U�O���{*!��zp��۱���W�ڸ�To'h��ol㯐ځT�f*�湱o.��׷�;	�y8h��ڝ��;�i��G;r�vӁ�7�8����VQV��eoG�t�o�1S
+7�PUy�L��3v��'s�BWV������k\�M�C���v�Z��6���HA��>6����Z\,G�ǎ�+�/�r��	�o����0(�,���îk�T��qv��Wn�pX�ʂ��3�A=��0��x,�AQ|'j2�rORO��(2u��5(��k4L%T���F��l���0rK��3�pu��F�a>�15v�L�bN��vh
������}m�v���4��l�a4@n� �g`�LN���ɝ�Xg;�g�������K&^v�j(��������c�]�=��f[��N{��� �tE�P4�,���	Tզ�� �����\{�38�3}�����f'���3:u@��9�w�>3loA���Ȱ6�P���i�:�wo�J��-�&�u:oq��Ә����K��wV҃~cF�uv�.�_V��kl��o'@���v�P�Zc�m]^Ҿ+����m<�Y��u����c"�C��+lN{}n��e7�֜�ӹ�ע[I��'��TN�)�^] /��ea�|xm��殺/*���p B���[B)��ofB�$=��pW�FK���$��Ϊ��7�h���0�+8��+��D�sI�7٤]GY|�j,�\;1�l�L�6&�o>P�O�;{wq��8����;#��]�x��T��k([]�eR{s�������o��w�{!ێg���z�j�*	���Ty�w�3Vu8Z,t���J�]go�¶���v�I&!�y	Ƶ�z���%-��z;����b]C�؛5Z�lU�F,�:I�����E���d:\H��x3��:�0��v[���A���E�ɣ-��[����fVJ��3�����$�f6`�B�E���{�a���0]�cI~�EL/�SD3E��]'����c#f����딳Y���H&�.�鶔�5��-��y���
��ݝ�*^>,�E('R�0P�s:v*</c��m�8�Vvc���*��4?.RS�5��wWy@n�+��Ձ��Zӻmu�IK�KMr"U�,- a��hA��]�l�%m!��l�Im
٣�P�*<�n2���pX� ݥ:B���[��uvE6���FW{�D�EgB�[��ھ�D��l�d���d�;�;tm�ʁ.�iS3D}��\0o(]ړ�.�\��$��uęz1J�Wc��`
nH���.�AH��M7�{:�����'V�h��u�Y:���:́�|��p��s�;h���&�X�;�GE�_H�iF�T��XνE�<S��U'd]��w�K)>�e3,)�P
�
DA�ۣ IR�d�fd!>�N�n۱)λ�����au�>�P��I�]��q�W;vF�u�fեkw&���s�R;j��h���gu
��=F.h4�wTӋ�h���rZR7�`N��d�Ɏ�v�ʲIw�Q�5yۣ�J42�%��-j9м�z)��G��R����.�#�n����y��8��K`G0�Q�)� ����[s8Sn�_
�.�P	�73c����
j!�u��&Z��SZg�W�r��g���|�f�KM�'�V4�ƝH�;���ӱg�&$=�)a��j2��ݨf�5t}��j�ˆOx[�t��gd��`�]1�;p�U���	sU�~��P~@�י������CS�LM�\o��;�t�U���cv��$@8:���A��XG/32�������z��=Ii*� �����WdH.�ʷ��9A����DE��[7�G� j֋�W��AJN-�̑�.T��jk�b�ﮭ�Yx�*F�����[y�x�:��l��7	��K:#Dp�:��࡬��s6��"�]���Z��2��z��k1t�ϫ�Κ��b���^^|�m���8����ˡtR��v$s�xC]�B�j���T�*�hݠ�	��Iӑ�;3�(e�E���Ca���4��݊�ޠ!�G)�7{���V�A��sg]��>��ˢ_9��s���,�OU�)�Ѻ��fKU�`Kٗ�Βf;��/�Tpe���MW
��I7{��6a��<��е��ba*�+yQ:�u��[�9�(}��a�ͩ�i���ޭNj��B��n����v-q�v	fe	��hsD�hC����u�fp^�rZ�Κł�2B��,�6���NS!��ҭ�r�#�@J��>o���T�͵�)��V�"��P�;79���چ]�ކU�S��V3���s�7Z�
Y�FE���S��霅���1Z1\�U[�$M2�p�tP��ۗ��Q(�(�Y(�Fgrzfe�42�.�F��R�K�H�,�[�N-Ve�sZ�`��2��g&��!Ùk;�Q�M�z�h��.���s(�뚜ծ�� �=)��C�f���y���8�+-\Y-U���JI̛"���{��m�1�5�]sF���Y�i�S��V#\�-}�C�oj!��Z�V;��ji�������K�� @C1�N��廎V%W0a�Z��rLŸ@��GqncQ;9N�eg>�6�,X��4�n��X����KZ��qu�I� !Gj�[<�'�LDS�Z^������M<��^��뭖sG<QCz5^�gnpEp��K����v����S�7'�;|JV\y�޺j��T�P����|-�GS�s*�W�!o�;�Y4I��DqmZ�\]�H���ڝJ����U;;!RYN��b�LC�e\Z�;$�=����V ]tx��6M(��k
*�rv���WR^mr�5m�%���s-�uk�]W����X����u<���bd���V�ğe�x�Z���;4�fu6�ݬ�%=3L�� WK�^�>d�kب�5�F���E�p1F��3ݝF�̼����ûǈ�0D���Ok:A'N��^�7�^t�x�gobN'e�2�F�}#�%n�Ɩֶ���H�Y
�٥�Vt=�����VZ�����OOV�-���8�l��RU�#��K�k�ռ՞���v����(���t�ԊMG �(���;���]6�y\�)j��"\�nL�4g)�k�iG��%�/n��҇�z1��G������K�͘�V�T��%�l��M�Dg;%ł�ƥ3�YK��i|��1q0�ޏ:�%�z�3�X�1��Hkڞ�^�����8�)�\;w�5��`2:�����ؒ�⋺��޺���<S�5��۩�u�jv+�ßw.4җ�
�eЫ��(�e�Y4of�L.m3Ǟc��pݔI�Y� 8�;��` �X�NC�!2����j�p��T�Ż�H�^�TN�Y�J쎧(��sN<�D(�����*�s�W�V[l=c-�����x&N�\����C+t��?�W�$1�����pK�����{��� ,QLX��M�_nAd)ȭ/�z{�f(�U[Xu��'���O��4��Msu5["mаC�:�7E,��"�ԡ�u�.u���@��8f&��w���Mw�[�s"BhV��u���Pw�g��n�㔩j��
7�e28�rK�=:p�:�pl�;�����T��4�[�wf���D�V�MqA��y���J�
��٫�m)YI�y|&��bM�n�Iov[]p'�u6�+�u�n�a}|x�
��c�K�E��wi�r��+�v�ȭ-A�9O-���|�j����9u�RTO{��b*�P�������5����$x���n�@a2�8�R�6�ً�Xn,h��3��#�֪�X��F��u�ś.oRn���6��b��.�n�pv��6oXs�+\��r0"��CA��Yx���[�މWy+�}`<�T]Q��*�U& �3-�	r�v\�',PF,�ut��t*�59��s��5at뤉U�	��K͟r1I��Ju��B�^^L�D38��ԍ�q&���$����ƚ�8@�b٘�ւ�Ճ�	��ܻ6�5K����O�K�QU$�Et�̱��� ?_�o�m��y.�zv'��Q�T*w/��K',�ML5�'R���j�nwt�Y�]��Q�#q뛚ƒtqfNF�3M0�v�q�B�=�gy#ס��y}�T��r���U��Ck F﨑ơ���U+�i;[�.�O軇^p��.<�:�aT��ou��;�:���b���u�@u�ZL��TO����>J>��f���m:_B!�2��.�R�����rX�ōj�tH��]C��w¤�=GG��2��}�*��j��u��1	�`��S���A�^�� ��i�Ǡ�\����e�G3&49�&� K9Y��ݸ��ڧ��ư�a��r�醭N=����H��"}��*GYTK:��N}��a[���t��$�������ř�Q�e
�@`�|�[��v��u�le6�ŗ�"�eX�6C�ǵ.�B'���`άn�i}ƶ ��ˮ��6��t.���=�.[��8���y�e;��9d_]t������(��Þ�N��_[4Gv�5*"�0Qoor��i�V�/�i6��_r�t��L�
�J+urS��;V�"�tHӍ�?=�u����B�ڨzE���#Pw�8i=��J0�'�$������.r�RJ �lQ%���A��-���;\8�Ub8z�<���v���7�rʮ��.��S�Dh��A�o�]�Zr�~�0qzQ��G0C.��gn�w�+�'4_�X��h��ĝ+��IT��k��V��c2����.M��Y�lP�]V�;��e�N�9�?qv���E�Ŕ-�������Ds鴫/
 ]JЎs]�P��҆�uُoo�<�vrg��j����t��X���d�uu�B\|je! ����D�Y��Z}Z�dl��뻕*/�b�K�EwVf�<;�%4*��GX�o4��Yv�5!0�Kh�o$��X���igvU�;R�U��$������-� +hU�ɖr�#\�7dksM�������Jޚ��Z��"�w��uhq�3f�h*�\fpT�kPBc�D�[�C�8�N����+��	��&��Q��)�&�����NM��P*e'Wt�;�N@^�˱g����\ꋧ���ww3��Y�}�R�nv�݁uu(�c�"�[�IY��spѭ��F�8���*I�rvr?��\��VOfuѱ\����h�j���U�-�6��J�QͶUS{�m�[bR���	Qk��YD�N�K�*�F�Z����� �cŲf��e��x�Y�vVr��K�R�Ⱦ͔�6����u�|E����jˮr�rN��7�m+��ۆ�eR)��ҶH�t���_M��9���+�Y���u�����R�ۮ�!CQ;��U��Ó9�|�!�*��Xd;�yS�:勤7�՚��wt�&˧j�3��Uͮ�z�]K����{|0v��;��dO�����L2�%��yO��gR��S��t3j���(f�%��u"n�K	����{����� {�`J	??���P�U��9T��oS��c7{b�<����hX�f����M�;���5����_4\Wr��{)R�;ڑ� QRd�2�g+�[.+E����K��^�YɍS�����J�ͼh��{�2�b�縆��F���_!.�SaɁ+hT�D��ޑ��6�|@���ik6,���<[2�A�;^��ы;��l�f%o�x�ԩA�Z�"|�l�6&�Q��l�L��wkK���\����)
�������֍�9�}z4v�{@��E�Wk��uϯD�lJ
m�\��Jd�Z8� ���n	F�L`�n��k�a4Rc�w�4o����kl���K����0O;�fb�ƺʼ��e���00��)}�7��w1#5��M�ޡ�Ed�^���v��O1Z���1��nX1��M�r������]�`���O��������
�J C�G��������B�v��hR��s@P�����^��]as�/���S�WEo��;t3���+d��
fX�\��j��D6Y1���k&��_U�s�d������uۼ˲
W�4����(w�RU�ʹ]h$��ᴧP�tɈg ,��'=`�.����{�h&R��<W�ks�u�E,"R��c��-8M��i��Xt�
��yK�CJKwm�&�l��B�+>p0�-ټ��t�a��˾����"��1u{��Y�k�i,)��C6��=9�Mpف.S:�gSKF8E�͠�0���Fִ0ԃP��4eʽ���esu<���V�]&��\�Q:`�wW�e<H�k��l������n�mjU�H]J�S��X��kI��z22�Qlu��3X�H�
]J^VU�Y9��oi��"z�.�F�^�ogZ��Gv�N��V�w;��%k��A�x
t�2M���9+(Ζ_4wPꂯ���_m�
Y���1�	�,N����7�mrא9���sZ	�0��{#�.ç]�;��e$6�^C�1�fu��RU��Ґ�y����O^����򋤝�Dk�"�Q��W��@;��o�#5���T��,�V�E\V6�2���ja*T�uqg1.ܑ�핳���/�����#�h>}��OV��r3�k�����:���eYﷀd�2�QFHF\Nާ��-�9�$����k6���մ��rw]+�����93g�W�fD����\�V��Y4�u��D:�Յ4®�]���{:ś��� Ap�^um
I�
k��a�v�ȃ�հ�M�da얫$P��N%ag���:�7[����\�����<I�O�Z�h��eeu��Fc��{a֡n�Mi44Փ})��@Ƶ�X��3N��l���̓/�X�t%�R�k�����Zr�j�y�:Mձ�
�in���Y�5�F먻��W��Wq���BG�����A>kh�,���+\z5|:�y�)wׇ��uw��ں�"�˾8�Zxwl��:�31��2c�Wx����Cz]��`���sY)7#�|��� �grd�����տ9J�?�3@�8�9��D��*6��]
��.�Ѵ��]�x���C�D�w�1*j},+
�)۲��sd�Z۷{ĬH��Ke�jwJ��\�e�W���o$u���+�Nm;��L�pn���[\��ܡ+�bi���Z�X*���ǡ�Y �H a��:�,�wjʤj�[��![P�
��2.Mf}`j��z`x�f�l$3��r�u��#�|�h���դ]c�Z�O�RB��f�e�Kcn4k)q�y�8�.��gT����/�jG2cS�s���#�J�c6�<3��S&�
۶�u����|ݻ=���c���eV�N�6��:�U�s��<�R`l����z�\ "����WQ�J��qb�/��w*)΅���������%���\�ŝ�]\ai��R��p�ķ���:vGm��ݣ9�ڝ�ۚ�_<��4�!h]�,�����Uz;��$��Cޭ�v4�ۉ�� 
��-7�*���8*����ňr2=ija<����T����٨\�W���5���y�����e-%^:��n=�R���FV���f��i����|������64MÌ��ܸgH-���pT��ci���ʼ�oN�HL�lN��n�QA
�\���VG�ظ<�Ucx/����)hBf�|�wf���$����x3�L�Q�S�њnTͺ4���G)�6�<u|�u���ȟ�\3k
$a�uƣV$�4oB�Q�v͋��,<�C�����m�m�V����QÊ��_6R��핓���z��w�henLr����`]\Ł�e�
�-�����sm曽s���P�Ն�v}��u(o�%��n�� Q��:!������.��y_<f�,�^Yo0�]��'k���٭��u(�A;Q�e'�p�R������i\�(Qҗ�i˩St���u�!`S�64m�R���8���uv�H�M�\�*خ���۔���U��J�ܝ@ӮÂ7���Z��cf	�v�\��R����չ�O���V��Åu�f�z��`�7�S���ݬ��ӨZ����N_m��گ���oX�gC%e��CǶ_�0Y��P�a��b���4j+�y��qb]nD�ڔ�.o.@2طnu�C�}�*Ы�<*j\�Y1�mi��.pZ���n+�y]����D��#���[3'%�H'*Q <��[�Ǜ�D%���k��0������n�ww[�)m�=�9�6���w�&F�ܙ�̥�[V�����J���봆�i����~ȩ�Z}��iD̈́��M��+��8�_'MX��ג�c�6É�W�u+6R[S���S]�@3oUw{u�KgT�U����1�ւ�?m�����Lc��O3�֩J�4Ѣ)w׫��YH�ˆ��-踱�o�v�&�z{;�Գr���u6�fa��)}��1
-�N;})p�1�W���E�S�v_R�r�v��=��J����uve�}3Q�9a�mt;�+�K9Z�J@���][�܏m'c�Q�G��|�K{�Н]�����Ħ�X��]jX��v��9r����
-�h�Ҹ��!�ݠ�9�)���P\���u���n*$.h���y�vvҬ\���A��ѝA��/i[fe����,�uo]�n����wZ���ک��� ���l?dx	����y�ڛyJ��h��a.��v�7d�J��Sݾ!A�U��,�2�����ܔ��^6��� ��&;�U�5�!��(��D�v�a���Яh��g�x�dcb��9d����T����kz�'hn!�/� �v��&�O�р�I5�~�,>��9�Mb�Q�i�wo�.pu �N�{�������UQ��^�9��}x��Tk-j����:�Ǳ���Q[��h���b���ʙ��)�.̆澮�x�ۮF��6˗[s�Lؚ��w*��G����y;n�a�1!��&h��~+tj�i�d�_s�!����or��w���g5����[� ��;yMD=D��-L������z����py�i�\7�qA�ˆ�Zl������1���n��F����͌x.���03�zvg]�K���r�T♡h�h�u'�E��덪ٔ���.��*!����+{��V�ovԵ��o�֨}�"�cr�uu�<�+�;���*��aWWg8�Wh{ �	Wb+Y�d��w$�[
}t:�Y[
A[���N�I�swJ_-�h�P���{S����Z�\�1%�{tb2�S=��$\�J���^��ΐK�1n���(��A��|�n��Ӊ85�>L��s��+���]7�2Q�Ck\2�!��Q�P�8k-9-s�|�2�u�Ū�$v@kv����Z�{\3�ITc�Ow,���a
*��w�V8�/���\j3PS$Y6V�mE���0V��(�9�yR����c�/a�92����܅C#��u	$��\0Q�/���"Z5�k6��G2C@Yg���Z�t�{���ٸ�!Uú�ۼ"V��wT��mF�����-&VJʋtjG��K4sq��{Fv5�.@�-d�ݳ��<(J��ΓQ�����&ɲ�gs�s_Zr֊�{�|�*i�i�'��W��Cv�D[�$q&�*����qn�^�n���	PY�vK�<mu�[��uX\v�.�8]�
a�OsR|<�El�?���t���7&��5�"��Y��JG��)$�:�ŀ.۰l_XB5��{�B��Ju��t� �H޻y���y��{M_9��J�F�l|��_r5��.K^o��k��`��0�Lub�f9Ky��غ�b�!�e:�r�M>܊XU�)@r���Ve}GM�J�{n��Z|�e�S3�*��1�Yo�6v�*�s�D�[�m0��@�U�W�RVWc�̊�p���S��B�Qۇ�yм���ׅX�]7pr��ɺ���w������_Z�Vnrə!�]);�&�n*Ka�M�3�U��h�w��ki֩WЬ�SZ�lM��@�eAQ\"�ɔ��G_c5òB����@-U�.i�\EvS��̥-+A�(67\T`y�>����Xq�yު���n�N��.��z�]Z���3�=����g-R%Fb���<��k���O�\�,N#�b�֗D:�%WIvݑF�,�űJu�|g x�x�"�t!�W�r�嫕oj!)�����4m����L�\�re�+��o-;c9�Hd��Ӊ&qz�"����� )c�Y��sչ�t�z�������Ժ�!or�nvf<���VWaȤTQh�a{ΐd(R��+n�TRK=��F�Ng|�]`�e�12����K�H)Һ�'�=��g5���]�s�<(���맄���wDN�s]�������
Vڶ5�,��B�z֪0t�g��u���>����G���Y��N:`+��ՠS5�Q�Xr�[���4�u[h�3�b;��vډq��5�29+$�� �Ǌ���2�����<C���$��E�Y��R�02W|�gʗ0�ng�z��gZv������"�:���Օ���.Gb�ę��R�G�	�ô���v���Ы�nÕ7��Zm����ͱs`���nj�Zϴ;Ô�x91�J��n�9L�,� �SZ-�v��<��Η��3r��� V�u�.��հG�,���v�2�T:�S�vk\;�h*9�c������->�ˣs����L��'Y�"/Hcyr��p7ZoN�����I�g��Ni倊XS�]}r����鷔��}����Ww�[bi�Ӻ�۟]֭e].���Y�{/%rWK3A�S��am�+u,���gN���f�)�c�iƩ�
����8�H��i�㲦pyEk�����֎f�D�I��^��d���osa�qEW��w�#p���Zq�"�-̓2���99N\WD݊�هl��^�υ`!d�D������0���p[������"��k70tW�Ud��$<��Z
*��G{���'j݊L[Z��	';!B�,u�uc���E�U��)�fK7���
5׹9Y�b:��;%@xe�Wql,����H
��b�z�
 ������S�5̺M�']�FNı���"�Lu:Z�V��X���s�$�(���sY=D�dЗ�FU��ZĻ��Qf��J�PH���%t�^�*� �WngI׻P����R��w����Z�;٥��蟠ǘ�:�]9%�tm��m�T�s�)xL�P��%��4oK[�U����[w������+X�u�n�{�oG��rby{Nе�Z���l�	��H�cgNq�h�zj�T�F��1hq�{���K.�nLǏ�
���]�)rOh��07����Ev���G'ד+RO9�1Ҩ��4���݌��l3N���L��Ո�q\����f��xM���:
$@�+$��XLi�jY�U�j4���"�:h�����g�m���7��4s��=�.ijgH�f�uM܅\Dվ4�L�z��C��N^Ȃ[��K^$ph4ӗhر�N�ۯ+kx��R�$���'Ӌ�4�	W���+)=B�s���+��
�����p�2�"@��^��<&+�w4�-��I��s��)]�;4,{��{	����*K,��@h�sm7�ˍMSQG����.�3�񣜵�{y��WX�u����֠.Nu�rvq�:'-3FڱV,[A.C�M���t���s^B��[м��}Q���ЯxK��mle���NB�A���У7��/�ػ�qԀ�:٫���SNb��5�΅M� �,�8ZC[���zD�n�r�HB�eƺ�\��%ϰ�N�"i�ne�Du𼮱��Vkn�rN�W);>g��s;���|��e�p�5��o������Ǐs���k�:��WooR��Ov��)�GVKD ��Xq܇��xٲ"���vx`z�˓Vt�+V�p�7F����Au�i�n���nm�����jX��U3���B{/Y�-/������䥔y;&��ܮARʈBd��uԁ��Np�e�2v;
����žn�+�r��I(S��I����@mjKP�ΏP�*Lm,���S������խ���w�R̔��Gr�,&o�������>��Flw��mc}�[A��H"V�{{��nثݠ�t�뱕�A�w%����F�n��b�J#�� ҰK�Λ]���}G���8G:���iح
�#p�9�֮�+%I%芕M+q�[��9�E��ծ�]��F�WN�2'h6j�e�=�n��iS���B�h���I���k6���_F�����N�b�7�Ui�Ip-Ҭ=7�S:��]�w"���(�G��g��l� ����Y`iX�7���I2|k/^�9����]�rz�Ow�� {��v����B�����{sKRYI��V�b��=*-U)�f�畍b��;s`7]b^�3�x4GȚ��s�[���#%]���A�`ۡ�yuXV-0,I��L6z�ӹ���h�[	(�쾷]]�S5��&g�M�ݔ�U���8"vʬ��V&�U����	�G��j ����l�{8,zgKwXV.Q�)�Q��3C��l���㸵�6V��l��u]o
b�t�V؎K��S��y��"�ZΌ��%4���-�Y��Sp��]+�8��:��Q�o�C�EnU���;F�B��r:T�� �7�U��N�,�����f�����=N��v�V�}��Io����|C꽃,��Lcz��>��f�v<�J�Q��qVA��
v>��-�aw�FWYK^� 9�|\�f:���7F*`k\yP�ѻXOӇټ��ۅ�_ �V�T�G1Z�*޹Q3��5:&Սuyd��,d*��Z2��(6R�d��Wv���t�p�*���%���[BxX���²�d���.�q���Z�+9�W��*ƾ�u�'0���uڡ����Yv��Y�e	��v���\���\�TX��Oc��vKD�	K�:1�����&�(�l�3��5�S������N8%�YC�:^n2:�u�ѳFm�h�Q�K��lq+)��z�������]������K�{+;�Q����ֱow����&\+�dG�r(��܏��C�U�%�J��+WE�;��G�r�UȈ����R̢��!*��9�^Br""(��WQ
�Rd���8Dy�E�,
=ݹȂ��̖Dr��d�p��%D�Ԅ�G"��'�D(ul�QQ�eT{�O9�ԫD��<�d�4�Dy�
/K��9�%�)�UP%�D���܏*�$kB>0��aH�������$���Bs]�.E�p�U��9�8UDDW*򻸔^��!Ap�k+^<�97>u�-�+;�숉$ ���%G*�^��E\�'=$�ӹ�HY$S�Up�][�aWp����ZD�`EW"MANU5-�Ze�®'Z�> W��������䋇k(;ȗSX��]�rP���S��q�V�w/�a,���b�z�J;�����B�^1�w�91�3��"����2�ZCj���� �WZ�HԺړ��:h��:����3ͪ5�٩�G<�>Y�7��uC��0�9tۄYcn��`��t��F�7Qx�G����stuC��׆���D960�8a��4zҘk´#��k�1xK���� ۠Ob�-��T��g�c{�v-:=�u����<"���عؕbv3ME��@iD��92r�^
;���1�<�ne+ֶ�M�otEn5��r�;��`~�i����Qin0~�v����2d~�����s�ܥ����i�@�x���� ��h ���Y�;���ʯ{+�皊��t�
p�����_Y�\I;P.'���!!�0�p[&+�g���-Ӏ��ˎ�S��.y�W͖zñ�z����cC%UE��/�Gx���^�I��Bu��9��N]=����!��}2y;�lŵ�W�������������0�t��϶���]�U�&3�6/o<d2U����C�����6��>�t4I<��A�a쥻��y�H\[�B���.>���O���ܻ�W�˔��K�e*�5�*�nk�鷹���V��Z��T�\ҹ���7�Քf�Y�'k��|T�Au^"�5��uq����}�]�h���V0�e���+j�u5����k�-�86��0��o�|PH]@�OOn�Y'��;��n�4��FBX�q|Ny.=�d(b�^�b7�M����{Rv:_��wD[C�b�[Әp)k������.7u�M�n��q,��u�oM*Ǵ	�+�Y}�u`K���D�"D�b��y|h%k�Dl$�(_)U��a
����WQ���q�����TCV�Mxx�&6Vӣb��c����6�Pd����N�O���6��&��4�/@'�<,��:x�����/�b���l�j�/S:��{p����]_-ި"��&N�$�^
�e�j�IU���\>�c������w�d4������7}�܎�A����i\��Bܱm��68�3��Dv�.B���Ӳ��	gWbC1u�#���xr(m��E�vT; ���>��S��u���*͟���C]Yn��F�1��� ��Ϝ�a`T��� �{:�DW����!K��a��E�t�f����*=Ö�ר�|���8���ܲk� l����j�Sr2(���$(����`��9���[M�wd�����UN�"V3�K뺚��
&T�[�L]�}v�gKj���f�tBo�����iw��u�^�2�&����������%����진u��^�祽ٜ����\��W>��3�z/^�����	������զ�E�LW]��^�.�{����i�ω�q.��+l~o��*������}C�f��^+sc�G��ZV�n��[���|�(��7'b��DG_�}չ��RW�"����uD��}u�ڳ�bH����U87�"xm�L�s��ʦ�U�E.�� �< ۚs���<���%�{��8��Ԕz'�k�V܊��N�z��t�1Ȇv�Vg��g�B
�V(l�6^g�v�+D����ϕ{L������z�ׅ�^즈�I�������W����D֧�fL�N2N�<5I��O�U��s*��׺)k����F�������"���}�����+�0Wʩ	���_i "'��ĥ[���	0�ފ��#6"�eu-<��I��Yg��Ź��6W�#b��I�Q�=��& 09R{��E|@��)�|'f��(kp� �[���s8�y
�!D¢2���V�ԂSsG��ޡ�}9��g�W�;�XҴ�ra�_�)��ɴ�w
�
�vd�Q<gb�n�/��f[N��JxR�0Cr��Oj����$:x�{�7Q�d���n���[;=��H�L��{G����A�Rm������u�w6`@�o�܇y^��h�Ƣp��۫x���r�Om˜���ݞ��bj��{u�P>��;c��Ko��f9�����i��V��3~88c��O�M�H��&a��r�	��r<��;ڃ�Է����(�Ƀ�IN2Gu��}^�0���u8�Xk�	U8��3�Of*l����q�wj�`�!�=��hS���\�!��Ş��+�f���4��כ�^5�`@��n�i���D����[V�l��֨��W�l��a��r���w�<R>�z��Y�\���Q;UbT�2ɘ����]7���#"��Ä��3�@��kC�a�OR��;�T'8vTB!�H�*�2���n�a�a���ԍ�g_�=���U�0y�c�<z�&6|/��:�ls�]��9ޏG��ML�Jp�^��͍�Zג�j�,Y$r0z\X3�lU#����w�%x=D�Y$/QJti�@}�h�U�������k15��",�<IT��U�2���bY��}E*xn'+b�ȪÃ���-F�gd��(��ym���[ �=] ٯ��;+�[W]�o�i���΅�MA��]/8@k�������LS���V׹��w��C�6����kgv�i�j��Q>�(���-襑)Q�Ѣ�t�e��r4�Y��f�g@�u��_\��2�f]�M�B�l<0��*7�CA��i��+'Q�2��J�'���)�[QT���r��)�üṁ��Ef���<�� Em�m =ܾ|�u�D�qE����ۯW
��6\]N�#=6Z8�F@���v�S3�� �L��\B���4J/�FZl-�0Ĕ�j.�����T+S��[����-��xHR�IBsse�:F���L<�֫/d�$rb%���&l�"���([�B��wR%y@jY��Rέ�Ɠ=����!�P0'��;B��e�
WV���6�۶
���UraaӲm^�^���w�

#�p;cɇC��ؼN0~�.��6?<�>Ⱥpwe;���nno��ܴeN�g���f������Y>��A>��J�xV���tG��wֹH{ڦ"e���XX<X�g:�{�����+Y[�ī���H��f��2�
,��D9t�EpTޤ���(��*]P,�9y��+ۍ`q�];	s��'W���"���:r4��dIB��J�f��N��Ft�¯ǂ�Y�/�	��)�4wy�;ҩ#��u��Jvۻf�+�Nva��~s}���	앚��"��L
��J���Z����L�y�1�s�V�^fn��q�Er�qZGV5+�:Ƶ��p�6�f`d��<ے�}r�s�Ǚ
��&��ƺ�g�Q��T�um�IW|f��2/�c���}�Rw�ynA��wH3��0G_�	ӕ�td�B;�"EvN�d�Ǟ�s��Θ�]o��\U�W���6�t����f��^�$�Ɔ��<]vt��R�M���+Q�.�I��w+�ݥ��,=��T�����$(�$�* =���2�q�8wQ����]f�,����bb[j�Ie��S�6�� �H����}���J���F���T� �W��l�s��.:2,%��:ԝ*����A�_����%�2w��6<���ܩ ��� Ǹ�����ثF�B����֧����^��bf3�[ⷱ.�_���DFf7^��D�<������ƂV��F� �V��D���KV\�W���9ܸ�1����Cx�Mx��l���F}=���ӕ�_!��*0u�O�K}Ѿ�s����;{8� d?B�����(�"1��[Y`����o?d�Fo����,A��͵@Ţ�2y�Q�C����,�=!�%@�qp�%�:O�����N�.�� ���v�;ϋwuۘ� >6n��.~$�7Y��$l[���q�o5e��Q++ ٨�j�z{�ǣ#�M�����h�0��廲��஬��6q��+m����i�v�ƨoX[ƃgy5�'w�[��z���λą�����[;��>�6̲�y	У\������>d�,A��(���7�"#���а����f8b�iO�! Ga���	�̞d�wJ˅��i��ث�緑p�NUD�%�U:R}���hY��G�Ɉ9�9!��J���3�DE�A�E�A�5Z�ŽTT�#�W�&���]��1���ȝ�&g ١��_�>�Xe.�;F��{a
ź݃,o��o�s�w&%&�;�&�vˣ�[,��3�tY=�V:�O��U{���*�D�������u��wv�L��e��w�
���tvtܝ���D�����\5�
�mT�B���Ł�ډ"��^W��dC.� ܦV;w���SK�:(�<D<��a���۞�v�
�����$k�Y��v�ϡʋdB8����<Uc>�Jݘ���6d��{s�#�.�d�@�DO��&(�.7�t%ڵ��\d_��h���8z;V�ɠj��RwOa��"2����J:#�zB(�ZM�y���~������=�/8�Y�b~��y�
k:�&K-2�$Z��V����'׊[�S]���f�T%�z�(Z3;.p��hbMh�uK�#��������
Eʚ��|�(��0�TK/�����ڂ2m_f7�+�xԔ�f��>��}���u��],ݞ��G����G����T�k�d��1��z�R��pV��&�>쓝�w����O��������s;��r��J�S�zd��=�ɀG@�Y��>����ݧ��j�#�f�0��6#z�	u�-�� �q���4���L9�`�b6.̽�|�=�I�]+!��Șǰ�ޗ��\�ð_�N��N@�p�`��fI/؉�&�:�c���3������t��}+��]�p��w"9�v�#��F���|���m��D>�n[@ҖOP�X��>�s�o�T�;����CP��fz�6��f���3�'���W��[�L?�F�?�Γn��|Fb�Q{HF��:�w�k�2��ǝzף��Z��͆$�na�p8�О����vh�z�g�3�c�����tRGم�ݜ>���W�zN��'��Xe�Y(Tӛ����0��T��o��Z\,��I���o)w*|�X����K���ذmB�*!(���ps��2�T����3�O��p���p(�Q4�	��{H_#t�-l�A`�6���:���ڷz�l���ȋ5]���O�=�)�]�&��.�1r.�<�F����V��Ov�u\�#e!
�\�����.&�\̓v����ݧ(���ۇU���I�1�\�;�}u�Q��#�i�\)�>c�X��υ��E�T�Zr��w]eY!�w�E�wx�m^FI7�,�D@���S;��U#����Z!aF���e9�OG9�MDY�7�C�{N��D��$�3�a�
��G���K6R��~V�Vs��̹�M-Û����6��dvW�dd��'ހ�y� jh�)@H�[e�cEљ鱒�sS�v���U��=�;N7&U�f2y>)�$�[Di֐�Ȃ�{�F�bz�Wz���a���ޮ��Jv��Z8�F@M�9��30�(�'bzR3�����b��nȩ�ȅ�;����e�2�_��{h%��F-Yg	�G���S=5���A�)b��Is�5Vz��G���w�[f�8<��i���{��8��Q��2^�6���.�K��wov�Rx�
�z�Έ����;>�N�k�7Oxc���S��d�E܃�w�5�3V0�z�Ԯj��Ih�D(l��/hra��?X�N0~�.��6?<Ì��@*λ��[��q.�E[Pա�ݗ:����A���ڼ�����葶T����gKy�Q���1�Ͷ8�5�U����uk��qg����P2��x����U��A�ʾLa��{��P&裺�]H�4�in�f�,U��OhS�[��^�]�����{��R� +i���N����m�����f�
Ќ^*����Y63}�p�ڼ�ⴷ1Ba].'��l�R�qRm:y��E��5�S��P?ץ6����s�{�]���d�w����Ң;ۍ`q���p2\�=�:���>/�-��<�������0�xU�V+�P����N̢���V8��A��O���8z5FA+�O�����Ե��u˞˙�����.	�:r�@������a.�9��Ne\>�ŎZ�{���}5�WO7��o�w>vƆJ�	8h	<�U�C�^���1�m��p��0U�kt��%KNxF�p���	��/�]sGP����'%�/���4;�Z����6�b�5Ͻ#����0�ȡBk��i\J+
��ʵ�,��+
���w,=�#��[�q��+�8���j�B�_J(h��د��Rt��K�c�
��m嫎�S�M%B�U@�;	N��{L���;_W���� {֣I݈9�
���˜��+4�;t���>�Vo��:���a8��7k��8dFH�F���Jw_1ʅ-̻��J�آx-���e-3z�ъ����*�l�1U�î�S-�{i���;�ԯ�j3��0�\l��	�POZ&�=j�
���S���n�[����Yݭe˜�/n�O��� knt!��;�b�R��b3����v6�橆�n�i�����ׁ+���.�OA�r)��S�LD`"v��u)�$�\1`
�vq[�Z�Tlǻ�U�O1\��o5Ȼ淚�����g��U�ge�ז����]�'�;
�#�@����ͣ��d_B�2k�ںT��G	�L�ُZHx�r�&(�C�!�IN�����2v��)KN`�sha�`]`�mZқʊtf�WgiA��ar�g��+�Zeޑ�gwoK�[Z��t�����^M�|z�X���Z*7����GQ�eL���i1�\�)�C�6m^fR&�&PĞ�:���T\].AvG�4V��mi��"�y#�iQ�R��U�VZ���Ɩ�%x��s�ی&��3:��}2���;;��h0u�.ؗ(�r�%WW/JWx��#�\�����Y��Τ��:o+��s_G�M�T�WoPwϣ�{ֈCP�K[��I/i�Gko8u͘3e�@H��[W�)*Kz4����_1xS`�r��λ�.��6��{��h88pX5\{Jy�ۖ�D,<=�r2s������yV*�9�S��\�!=�:�$��`�7u���ö:R�%=��`
��`v��7#��8�@���*��q���!�3Q9*�]_R5�:���ME����D(^p�SV-�1Z�	;]�ٝ�ef-pdur�p�V�@bEřU��9V���	ϔg1�eq�Z����O�3b�؆��_W|Ԧ�ٵƇv��Z�SbVB��5h��0pͣz::��j�N�INLvrU;%^�o1D>��]�G��Lz��@�l[�|f�[�xj;��r��=��`�ԭ�uf�������ʐ�em4[����ԭ��ޤ�h�z!P�{Clo �*bf�3;��ʋ�&�,M�ӹ%?_���Fg�],+U���0{k���K���nD���҈�2��]3<�&� �&�Y��s�ciX���7�*iܬǼ����`�>�G�k�S��Ʌٔ��Z���x���t�*�F9K�:=���Pe�V��Zۺ5D .���	{g�;�+:�#ڶ[T���Κd�=x�>�&��Quɗ���L|�7'ȑҺ�!�"z�s',�ڼ���pN����>�87�S�j�Z�L�n�a�:!�]
4����t�Iz�M�M�w��Y�����Ԫ�tRV4]Z�˨��4��xzfi��OV�&:��&���o�Ҿ%�$��M �W�#S��<�id�����e��Ma�*̝�� I;g�DS~x�*�r"�$"��2se�QZS�f�z���ī�P�Qĕ+C����� s�d��lIS�Te�u���"�Y�U�Gr�t�5
*�0*�\#B�Y�u;��8P^qT�̺�)3�(��$'s�R9QQ9!�s͕:�\�*��UEh��'Bj�t�s� ���C9EkB������R8��bfX��(��d]�!m+�ܓ8YaN4u�$���GIQ��m"�hJ��k�9Eģ#TB9w&��F��;
"�騄\���鴄�+ ��Z�WD�Qp��+ �ɹ*V벜�eG\�U]M�U
��(�eI�d��p��"����RB�g*(���9r9��I�\Ѕ�V��*������=��y��ʖ�#wc���G(V�G&��b��n%��U۽G���p����4�n�j�]G�|��N��9N ��Њ���y��?��Ǵ��6<~!ɅS��E	>!ɼ?���t��=?�ܜ�_<��޿�zC���7*~�_c~{?�I��|v�|�����@�I-���q���,�C;5��n��������������v��M�YM�	�v���<1���w�?��0�����Ѿ���������d�v�N��|��Ǥ���ro��?�r~!�ߤwO�} ��
���ܔ���b�:�,�A#�b���#�}��,G�;]o��7��I��:v����M����>A���1;��w |y���;I�'��z:?\x�ǇN@�`x� g��iG�c}�o3�̿߿�}'{C�܇�='?~��;���}�����
������7!8=�����P���n}�~��SӉğ���_xޓzBC�����_vܜ����x�~\�Tv=��Dx]]���~��q|���?}���~�:w�i7����}��w+�/մ<��� 8}��}�8��j����aw�����n=��ra~�l����9޾�w�eӹ�O� ��;zNp#1���D{`	�ز�(�7�3^�vw{~�w�%I�����0�G���]�� '�#����v�����z]�9P��{&���v�߾�;�1;����^���'�aw����ͽQ��r���Q�"�=��:��z��n�z���x�{�O���O���߉�{�cs��8��C�ٻ��®��g����~G��<L�S�ې�>$��k���������;^����N7�$������<z`����˝�VO}���߽�������Oϼx�N�o��N����q�~[�{OHx����;��C��x�<L.��㹓�!�aW~y��7�o[w�|��N�|$�AAA}�}�Y��x[W9U��]���8� ��G�#���LL}��i0�_���>��;z@�HO~v?���ӏ��~[x�Wo[�ro��!~^��xw���������a���XB"G�
�=LP�M�^��z���]�P�Ohs����y��tﯾ���ܜ������m�c;�����U>�_#����$�������ڻ�����O۷�;����yۓ�4I��� c� ��e��F.���y�8`��b1Ӕ3��=��y>���Ȗ2�V�ۓWl�gF��a�;ɛ��F�²N*���.碚�ڰ6�*T���Z���t�du�%ں�wk�ͼW
���A�@bz��I5�>}��,X�j����û�t�f�!�R��owM�ԣ�(�1�����l}����ި�<�ޏ��|��aM��?�|N��u����]'��S~'>Ͽ{���\r|O��>��0���{睗ۏ�9�����I���"_�����ߟ>���������~��NӼO����V��|Cã�������כnSz���x�r~�|� ?,I�7�oN�|�0�{`Rr{�p@Nt/�e����W{����_~;۽!Ʌ>��$�����cr��Bw }I���w��&�$���7��o��ޯHx�|��~��x~;��@�����;�w��y��DE���}">ܼ�}�J�k�wS[�oh�ֶ��*�=q0=p>����1��ǟ[��n������A��8��������;ï�e�xu��������{:7;��|���|�ޓ��+]G�",G�,�z�y ͺ�)�cRn�Kp��lDz��1���O�����L{������|B��;����&�����Ǥ��1;�|C�۟����s�j���/�}v�
t|��~�]�#�#G�"��3���Uʳ>�뺉:>�����#�G���[�p<" ��߾����9��}󷟰I��}v��~'���t~�~��oi���'��ǟ��7'���n{�b}������ǝ��1#��>���]��8%�{�<�ez}���w��9����&�O��?_��������r���NL.�C�����۾��9�����7�o�I�����������v= ~��O�����ɹ\��=Q1�t	��y�g¡���t����C�����V����� z���o����׾��;������ݷ��;����}�=tbw���}��zw�Ʌ�}���Sێ|C���7 (���W���}�w
/�Ch���o��wM;�����9>���~u�}���raw����7�90��}��v���v��͟�}�Dǲ���0<����10����|��zO^F'_>��V�_�8U�Y!��������ΝQ>��ēs�����;��L/�폿�zw��A����9�'���O�'�w�~���&�ySx�8�C�{?��<��~�����=�}I߮׿�כ�ۓ}B����d�X�4�����f�	c��4��7%�,�U��o늃;2�ަ�|�/�}��.�" �G�KD�Eq���������f�r�Br��	I�ڴ��_ۇ�`���W�u�
� ��)J���4x9��2��:�#nյӖY<���!�9�k�Q�[Q:;��/�h����P=$��� =��'zv�9�y�|����N������ӏJ���&�NNC�Ǣ��bw�������]���ߎ����;{;�o��o�/^���*�'��2��Jq�
�=p���������N?���I��v�ܞ����SK���wߜoHx�|�S�}������&����nt�N=�ǉ��u��}�97�{y]P��1;�}/��]&f���'���]��>�h�D2����9��'ӿx�E�x�C�a�m�y��7�?Ss�ۓ�OW]��ۿ�������
��{����7����{v�w����>���ߏ;�ׯ��_P�b~=U���r�[���<�<!99\
o�}<��'~F'�z����m��O�cs�;To�����]��T_>w�������ty��|O�9?��ם��L.�O������?P��&�����q�����}�Q�����>"G�B"G��? �/��O[�x������Gyo�nM�	��<v��8~�o�x��ǾF�/���@�_ϝ�����;|ON>8�����7��'��?���?Η����mWU����>�i<����!�������zw���8��Wo���)��o�w�Ǐ��;ߨ�ǉ��;s�e�!�}M/�o=�����a�~��6�����;�I/��}�5Tޝ~���|G�,0x���m��Ͻ�\
o��y���c����?�����;�s����8���w�׉�]�S�>���~X�艏TyÁ�����#�������W�y�,�o3E/`'ٜ��\}�"�} ����޿�~!ɿ7ߜt}v�w�x��'�oןg��?��&�'��ϟx=��p)��}�rw���������O����ڠ�Q��˾�J��V��<U����7��=T@��G����^�����9>�������'ü��9?��C�=���SO��;����te�O[�߾m��w㽟`�վ;ro��;�k���XP䝿����e��oޠ+ޭl�6�_k�����">~���Ӆ��7��7�~�8�q+�� {�
���R#�Ǻ B���>��90��!���������q���������0��=��I����0{��\�h9�9r�Ш�]��e�f�j���7V��ݚ\�ks����q��b˷�[��8��;1��ت
��K���:+u�\9����Ͱ	�Ӈ\ٚ�`���W|�k��yڤ�Y|��
�1;�wCz+z�Z�����E�+
�*�4���o��?���O��ri~��G�x���9/���x�N������{hܛ���Ϟy�p)�]���zM��bO�|M��q�����waw㏩��!	�T��ޏf��R�H�� >�~�px���|��'s�_s���NL.����<����&��v���w���m���v�w�{�����$�����zw;I��?o����p(z����߇�e�}��ܮ��)�n�)_�(�����nw�[~���]�aw�G��_N]�ҡ��c�|�9ߨ.�1;�~��>���&~�|��Ǥ�C�q��~�<W}M?�='��zL? �+�W�q	`/��[8TW}�̞���UV*w���m�ݼv������k� z���M�	'o׾��;�i҃�������7����z�W��?S��G�o=�''��]��?S����J�FE�~�g�{�]?�|�G��w�;���xc�q���X����I��Г������#�N�rn0�b2Ἳ��τ!2��i^Уyg�w�=�Q]�b]de���x绥3�J��HxE��k+CWbU�v3J�Ph�Q���۪+��#�"�[�@����+���W�x�r�u(��`q�];z\�<��i�4ݪ׭��͙�{���t�^�]��W�vp�+�x:q;2����}w�q�,�~�v���J�W�ܞ<��Lf}L�Ƀ]�ˋrG��4�5��-/'0;���<)!�9�v�G+�S\��Γ-��{E�p�U���{B멍��$�1�猪�I�tK����p�
o(kzb!�k{e�v3�YC��R�9l����-����xt����s{����W��\�N�.�Y����Q�ݻ�5
���FE5��'����<�P�u,ܕ�f�J�uu�].8��|�/7���]ŁǼ�_RJ:M�纻6�^*�}Z�}ķ����{p�K֮����õ�5+ϟ��ˮh�l�\pq��w�7�+�������E\�b�Q�Af�QQ5�kO�IEi��eZێEl�x	ފ�6�9���$a����/��˂!#�s)��צ��	c�� ԝ+�Z7�^��u^��;�&�|VdȮ��#e��̠9]��N�U�i\)�y����xK<,-��o��7:�&�6�	�T���F����D� 󞣔F���	.��_��e���;{"�5xs.8��!�FC&�n�!ۡ:,�����12��W�������1nkz����~j�&�n��i 4G��\l�?L9�����j�6�k�gv�={�m��´�O��j�P��L�6ۨ�y��4�2�
�2�>��^Vd���vƯ�Ƈ�G�f<�czk�N�0g̔�b�YFim:�4VO�ٻitR��gKDD9r;�Hxr(u��E��P��r_���0juBw�q�N�0� ֔{n�\����*�GW2��ƒ�5W{YY鳗�pF͵q�6To$��/��,����ԛKt!n�ҭ� ��W*vٚ(��fbJr���]��=�7��W7xp�We��J8��`�5&��
P��Ǘ�tk��ֵ=2>�_^z�*͟$ՙ�I̔Wܨ�\�{ 3og ^���p�6�|�� ·)N��α���U�i���ډܲjg ٪\����U����\��9iq�$<l��(�cW;1~�T'<\])���WB����-�XyR��g�a��l�8]��]g���3P���&�Jy��n��3�/4s������_�d�*���J�*r�&f[�k�G0"eFX���Xj�H�-u�5˃�D2�ߛ���n���"��
Ú�s&�������S� �+ �¼	գ*�F��\���9�q��ҌdC9x�,�űtͷ瓩�_Gg�����A�~����\�wI��v�[#��ӯC��/�O6g�����1�NY�H���.�����8k�۰�FIf�xoO��"�����pߥ���Z8�n;�� v�}�v�1��:�|q���m�:��'Z@i��x����%���VI��x�ҽGn�'&F��W�'IN@l�;Y�w�� I*/�R�(:��n���^�v��r�Q���W/p�s�}y:�ީΙ5�Y�XepBM�m\���=�2�˲�[���(l�œ^��\uQ)많�Iԉ�B�Kpվ�&3�z� ��͖�]�V[��=u#���oUC�W�ٔ��N�b���U߬����i1���zԺ���/�g/*؊SH��S�4K��vB�U��27�*B��l��{Ҵߗ:0�5$SIٓa9^J��Ż��\�֮=����Nْh3��>ڂ삺E�	�OM��u�'�%V��A�DOSS�׃���նCKۋ %��V>y�h>'j
�/n{G]yϤ>�w�/kL�F�}���NL�w&c���m�a������0�$hS�Γl7��U���9�
]J�nH�i蟊4�_pp�z��!�6���]	����TA�����GÜ9@�]��7͹�W^���`?ƉG<v@�}A���e��F#�W�jo�����!d�u�g,fA3Wю��;���X��Z^fĢ�ǵY��t���2�N�+=S�3v�,]X���M�bW[�0��p����@��
�|����� �ls�\q�}���r\�>������_Ve�+z&��hG��Ek���8>���]^؅){5��nWlU9�2��W�0@T�55��Ϲ�S�^��#T��V���@
n�77+(���x��~�ה��%v��	%�u�2���U|�X���*�c4�q���:��S%�D*��)��{6�v�Q_�Enn��8���^�cOn�Jm_���#��{F��w��]t!d��I)x����+��o���z��]g�S�����w:�"w����h�F<���Ɍ~N���O:� �Mo�	7�N/l�7V���k�*�q�mX�2�q��q�s�Ɂ�mٌ�摚S0`B"
��R崋Z��ݕ�^�=ƴ#<��6���/�\ioWG`��2�q̌��n�엎�8��T\����6P�$p�4Ey�D/�����^A��8=�.�
1�VY�of�v����H6M8���M{�e��H�'������k�7��ӈ�[�fM����!4�ț�if>ab�%c2�9�!:*_ ���ymmgMl-y^��n��ou�Q3Ԅ�y�wP�ܻmF6�����	J
����J'(�A���8Lc�/(�.I��Rk;R/�{�GBR6+׹AZN�Nju���P�m���/�ٜ��tw+
69����\�l�b��MҌ��O���S/:����4�k+CWbU�v3Oe���c��.wN���7k4�	�����l���]2���[[@3�`\w�2��wA���$Ҝ�]5��p���,O�=�F�U�������"��%������s������C7{0k{+��1�fHm��y�Ո$�N�{L_������ V<���W�`C ���2�P�FNB����ɼ�u(��`q�];z\��kY�0�����x�{�\~ݙ�S.��+�v���{OT�ve����!u��S��]E���rc�8���Ǿ��~L��ˋrDx�~�g&:��:k/��8OJץw�w�K�k�**��LP{<����1]<ޏ�ݍ!{Up�w��\�2U����a���i^�[���"0A�A�s��#`8y~{a2-ҧ�V_B�
ϸ; =^Oj�J�Ԑ(ߢ>������6�xp�=�ִ�%�@�eZێM��m�=�D���[�w��G<�P@Bb	�&���>�uI��^�r�"��ijN�Q5��t����s��e�k&c��V@v"��{D�P���C'}�����E���y�C)�8�q��֏V��~���݃��K>���d0! t�by�h:)ߑ��k�u��M�]�4՞��fT��2�%*���F<5�J�j�
5�����A�^f)��ۋ"k̥kw�A�뼱Y܊�Jm,ܺ�4h�Sn�peE�)������˝����Jw5
S;�F��X.����dѐ�)-�F[�4�겴�&�ʹz�rպ�p]��gO�p<����Ѝ޾ݦ@��(�@^-l�r���r3���{�Y����^4fl�|��B�����IV��� ����O�U���#H�Y[ޜ��4�Ƶp��8�"���loJ�i>�X	�1B��&M�J���(�aV�U�-nv����(iR�.zظuS�}^�m���Myu兀rw|Fk�2m� �B�z{��-��T��nJj���~G��#��r\H�TCÑ]j���T43c�w?m������j ��Yyy��	�}U�\߹�f�%��c�l�Ͻ�VƷ+�o�u�҇����XLqo�E��%Oz"�߾�����L�L.�~ߑ;�L��2��g�A���i�z����D��P	B�����g����b��tk+���9$P���@q�ۋ����b����g���S�<_\�ѿ�!D2�ԧ�}���¿9���vPΛ��)+l�}��ĭs�/v�ph�@!��%��=��g0�5���F�po�D2��nS+�~�n�wd�nH�nZpnSJ�d�
Fp�9`(�xG
��ѕS:snb��T�ڴ*���U�W�����p�#��*�b��'�v�;�;re�דm�o��u`���HR��6�v�Em.�u�SIV1�1�o
静�ٕ��I���)t�7��9{Сw�Wrw�%]k�g��]�X�9]�1)���G�wkg	pu�1h��+�F�E�7[4�����$+M���F���ˊ˘���m��\d�,����dbi2�3pL��!�*����d@{����+�lT` j��l���R����5�1��Î-p����C�d��+t�y�ͭ}���=�:w*����]�2��[���Gl	�:�vJjoê�i�;m��U�R�a+�66�N��d"�qo�7��6Mk�,�z2owVlҎ�M�;Z�V(��IP�\���â��������G���瑥7�_�+�$�Z�w+�9Z�g:�+��)Vz�=�2�#�g.f3Yt�C��>�0Kcp��`�El[�'������	����뜴���]�@ӁG�қRp �E���͝,W��؄�z������[u(�k�\T쪜�r:yR�&i����;�4�F��Y��L��U7��1�k�:�Y;�w���ؐɮq$Է�aL�����ϘU�-��8nv=��`�Xy!��JɩkAZ�o:'L��Y�+���H޹q�r5o�1�[*�m���CK^8Q� lm�fRt-���9k7��;��V�iV�������ѭ�R+Lky�q�f#ʳW;&23{��
|�Z����#s��О|�V뒮۩Ք5���n3�JHQ�T����eц�Њ��O�����N�M<�^�]P��n�CB��m����仁o*Zm����Ǐu����;}�k���Q@�����{���yV����ջxx=�%:ᝐ&��3	��G��v�mb��of����Ȍ7�l�T�t��b�YG����|�Ζ���mM$���Y���;���ײù�,w}t
��ͫ�VR�u ���s����\�%gRg���Mx;�*X�� �ng-,q��n�+-�!uM�O��J��qH�]�ůns{I�v���Ю�.k5�b�u����_Zvx&�_::�ۼV�̹E�`���l�R�:�q`\�&��V`,�,���ӄ���>���2���o]FvK,3�r d��R�+t."��Vc��J)PM�`kp̾������w��C���v��\��a�S��*�K��j�v��T lN%n&e�Ӎh��1ns�=Dޅ���5�<�+y�l�TX��b�������!��Մf��htI���-���qֽ��4P�����3y
��ΰ�j�V����ʛ�}�{�O��Q\��f����)��e.b�oI����&_V��-�wt��ˌ��&-��g ����lghI^�V'^8����9��Of<��N�^�K4TtO%$�Վ�L9���9&:2:�A�Vɬ`I��r�G�G�4%�:��}�f�`Y;��@UCE �$N��S��-
�՜�Z49)@U�jE�"&��G��b��1RP�$�nN�!E",�ZHTFF�,�t�*4�,4"Q�'K���T	��B�&Z%�D(�B�QfeV"��P����J!R��q
âaA�(�"�ұB�'Vr*�P���H�����U��H͑		W5i�t�-�b$��,�Zp��ē���J�8P\%N�(L�"�B5	�sHEbH��)22.��THq&�B��j�ar���Į�$�T˔QHWe\��C�&uX��r��Y�ȓf���L�S�i!U���EYR(�Kh�JfY�Shj��T)��AUt!+�i���II$ȣPL9'
����d��%a�"�9�etP��Ƈ�w6�/H�ĕn���:�K�H&�yc�6x��>�Z.��]�\Vʻ����D����f_ġ�Y�.3;����Xds�'ޚj�g�Q�� .��X�\��z��"q1^>U�f��zt��įeu��A\��˚��^���ܝ�����A�I۰�FIf��zA��IJ���e^Ӆ��_-8#�O'�?t����}��g�o��J�i>F ��=2zt 8ǂ
�Dܻ{��� ��)��:u�U�b%���^z+�t���vg<�k ��b:��Q\�<4��Ѡ;���-�����
4.����뭬aZLd�5nXIu�6܎��Ù�K�U�2�a�_Nn�%�+��c����3#��:�*\��{H��+M��ч~/�I�d`8�In��qp����Q��3UVh��fI�qd���Ђ삺E�	ž`���B~�|��cV�^"������>���#�j!)@Z���W2N��$.�D�r�uʀ�!���Y��ڝ��՞��^:-uR�R�(P>/yS�F�X�e�0o����{Ex��QI��n�-3�ky��F�ߩ{=�mu8B<&����H���s���.���!��)����ٗ*"8TF�/:���D���y�*έe2_�����i[E(���=(�����q[����2��-���h5���o;�#r1��S&�b�V��&��h��A�b<�dw�Vl�x�2��Wnf��q��ɑ�!y���꯾�����q���G�\�u�Ui�R�(�; H�}a�g�d�Db=i��[U�l@��Y�Kū�ka�=�����%���/��J���da�;�eB]Ө�}�*�SNj���}I��̊�J��;���0��#b����2���gJ�%�ͤ�������	����һ���w���ld��Z=�롬1|E�R��d�̀g�E���6"����$C�Jл���>�]هlE��ׂZ&���m;��`*��B�GB<IU�>��X��)R���o�n-�zm�]���}E*xp5%���ai��c;����Ϋ�5U��^g5�ݶ5l�ձP��;*���mX�,��;Ny�0:��1��3B6��y�����Zw�ӉH�D.�U2�7U|* G`X��ޮ��)�d`�{-H��U.��;;�8�n�T�`�j���s%��\�b ���-���xt���u���F_����ZQ�>�k�;$�3I�^�\eI�29��F	;MU��*��(y��p.o��a�\].�AS��L-�'j�8�n2>X`�ٲo�Z2�m�|�M4�q�2b�3f���m'�Rx�o�
Gљ��@x��i���u��^\���)���U��a�nM�+Au-��V���È[&N�؞�U��_��xA�r��ݼ1Q�=G�T�x2�9�!:�(��A��/�)}�5_d����W{�C�%;�J���Ֆ����rn<P
�����5�t}�N�v����!�*E�-�};~�;��Rmm�ۭ�ސJ��#(!­�6��k+1�Ց��/��3���z~ꉺ��\N��͌�W�*C�,4�k)��<��w$��,�5�ۦ��
6�V�h�-X�ճ��->&�U��_���\�l-���p��<�K��Y�R���8�H�g�h	�W��t�vg���P��f��4Y(c�Ɲ��IrŅ�~�gop�������{,�� $"{���'�pG�_!xN,�~��<.�9�����1@-�n{mӁҼޏ��s��"�N���{�)Fdж�{a��J;3��E���L�Z����OH���"åN8����$RC�H�WA e%�����\nA&�D�Dc��C��QP�bp.V��K9֮���.���Bu��ÕO<��v�5{��Ws�
��W=ܻ����B������r�{�z��)��2Pɔ���� \	��B����g��].�)�\�8���Lҡ[��ۍ���M;����z?�+Y�.p 6�je�{ӆX�mԕq�ƛ��w�V`,5|'����=��=|�f]�AF�#�@%�Lt�{����9��צ���i�gl���Y�!��lޛ4�J�ey�^�Dx�� f�( k�������*yk���"����%f��7I��r���iQ��w��:z%�O����W�
ϫ'�h?h�~Q��c!V��5e������:�FC�jr��%%9�;@����$k�d����UQ����Ջ�ݹhˈ-]�K�^Q�N�D�$�A^�i 4\z����'�TWݎLђI��Iج�����^�7�Q�͞�qܶ��]PE��L��@�BTk��&�Y���a��C�sS��<j^�k: �����+��WaR�� ����g̘�,�v�Yt$ӄx������]X�|�d��������ʼ�}�+�+ߡ�`Qo:�~B�^��q34�W�������\�[=T��\��*͟�-��p��{>����^`�vLd`�'���Y�{�r {|�(��-K�!���o��W��.�K'v̅��j��JB�][Л�u��ӂb*��o�
Ⱥ�����k[~�~j[ug�c=��s:��ξ8q���o�+�pu�w8�d���y�n�)��n-n�T]���D�}��=��fa�	�hۃG'[t
�0��m��I��gQ��WdV���xMh���KZ������%�H舑|��X�t'<����U�-����rF�,��O�o�S�M͹�kJE�T6�j����~;,B�K,�Jy��-ߜ&z�����N�;v�%,���Srj)H`���D�ú�}#�LI�����9��~nS(4��絔�T[�u�	��ަH�.:gkd���2�&�pt�����֩�������){D7��2
}Y�5*����l�[Dq���z���,GI��$�E1�n#dt�g=�k����Of{�xf=V֋�ki�g{��A�A;v�,��x9�+��wk$���Y/m�}���ޥwTk���tP_X�t�tX
r���Gc����J$���")���V��b��ǵ��{�>p��Ȋ|V�O�'IN@l�;Y�n�"Ü�F����v�:�vqʷ"�*�&a���o��D&zIZr3�L�oA^K�ɰ܎����2Z��AP�;������Ѵ���ć^��R��C]�ƼV|#\�`�Oh��78 ��`��P�X��̾.%�۽�\~C-��ˬt�V{�YD_z�9p��[�b5����_s>y�v�o6�T^Y�Kv��>{w���CE��W	�L��!Ģ�c+�MM�%���s�9��M綋費V&�!�ob�f����uPĞ�������8c��W>�ɯF�U��ut�zK���k�`�k�Ճ}�@��ߖA7y*/�`^�`��y��PQ��r,r!L�R�&�O���Rv������W�%�S�.x�χEyڮ� g0�0�UN�u�|��+���[#B�Y�m�x��Wm�c�Ӧ.{:�J>���Pܥt�����콴 d��B�18�z�%�-%�?��[��]y8�>�1^�8�u�Ui�SȔp�&�������N�#�5~��U�`O;���?/�<G͚���F��K�A/���l�{V�\A��)�ܷ���J�վ�A�&��];]f�N�Ϳ'z��i�:hu g�u@�<>x��=t11����P��ښI�㾈kci@�ܦ{�G��Mvĸ�4`��e��'t�[~�x[׺ۋ�p�S��7^Uo�]�K��-�{~N�����]%�<IT�"��2������ij+O�ea�.ģqKg�R�����h��x��m�w�b��P�zfcב�V1���tAW��"8��4��u{�:u�Z�$}x'����U3�SF�^:n����.&�m�-#t����u�뤮t��c�6��C���x�T�G���\l�GkG�"{��d0�K�:u	{G)��	����\�d���Q=;�xx{7i��[� ��t-W
b����i���L��)���r`u�F,�>��l�{I߷O�$W��"�z��Β��@�z��\V��oJv���Z"�ͺo��޴���q�.�b�;a�#0�<o�"��D*G}��T�W��+ø��ߵn���CzH��u��¶.�������y�K�:OJ�r�}�4���0����VU�"{OekVg�󙂗��dpCd��.�D�B2���"<�YU ��_0G��D2�G�H\���y�����WH��ݠ�w�=�Urla@(dx*?���'�y��R�C��-2^��i`��S��wn{�GR��B�r��ޜ��QM������&�P�tit���V�zJ�]r,�u.�0n\u�O�zn�e����=�)��u���!�����&��b;swS�������k6`�xQ�F��R�]~�X���[5GO��Uz��t��Q�?���xj��mf�����{uq��^�S�k
K���W��8��E���2��t��V�}��L��A*�z�������ۇ�<����Td�8ǭ,\*/�c��Or�����.�y�v�v�!�;&s�9�ueL�S�����_�evuY=I��q7vC:f!��8���-�+[����4;K�U�2Ү���H_{�����Zk�G�W[�'�y��.�+:�i���Aqn@H��>ۻw]���X�U�J�Jֻc��6�9�������1^[<��'��t�z<6����vƆH�������<9�[1xl>>���W�_1�~ߤ�G`p�΅��,�t���{a2/��늳���/ G3�֒������5Á&z���^�.5�>ب�|xTJ�OO����l�y�(sٓ�c{p]ƅ�xT����I�& l�4
�yJ~��7�X*ʻ�]Y:�l�g�Vq\Nc%ǲ��
A��h����+��>'}���+��=9W�b���+q-�>��FWu���Q���/�݃�}��Fx����E��]F��<{nԄiQ����if�"�S�J�X�ؠ�V��(�����F�v&�,��A�Fv7i�oJ7��[pgW0�lÜu�o�W��u��.QCyHd�Ӏ��� �,uW��+��G���=Րu�=�K�'�8�UGq�p��9Gx�<������R�2m�Q�>S�h{W��e��k��]F��O���|���X.��J-d�k�#wl�����E	�E�j��3=1�U�*c�#��A��	Q�{T}�Q�ź�]��SE�&�S]bΉ�����f�wsP����j�3P"�N���-��6����Wg"{�{� l���SWuW�t�$�G���Q�*{�N-���F�(�/�x�*��x^�
S_�_j\����{�:�ϸ�A�1]̲��|X�F�f��g<&�b��*�|�;��*m�O6ʍ��ݰ�:�!`���_]�fa�s!_yvk��W��X��C��Z�Wݚ�.6?7j"+qPqp����5O���SQ�q�רe�L]����+$.rI��u{���Ź�3'��~3+���HQ|��l��0�Z���碧��z%�j�9�E�C����n��NBs9���
�N�rF��b��&�S̾�n��Xs�3}��s����i�{�����8%T�I��<:�L�+���,u��"������"h,���c�����	��.���~���x�x�8����W�Z�ckϗ,�Q5d�_@��1/i���7��:�f"�	��XϬ�
i'�����b�.B�݌�6��y}�Uf��H�c/qEE�R�!���^}'Yq�p�N݆,�v<7��B+�����L��r=���8m�y�Avh�����R�X]Ve;S{�T0�������9�4��3+�|po4��s��Vgvd�Ukq�xz��R��B�Ԭ��71p�X��sw����+ 2����}�ą����p>�� %�J�Ӓk�%]}j��G| � 
�Y���OUʴO�����tW���V���F/i��y��e�P��ĞN��n�PU���)���H��񃞮��bҖ�W��:H����s��m�}v���#�rg�bRbXG.yn�}�$�S�)���D6zzJӑ�2�#z�.�&���!�&�+gg'�
����v��=<M���Fx�j�4��6==0����͞�}��T��ʾ[�;w�ܮK0����d�@�Ш`��B�i�u�_c�}�PZ�~�:B�]긕����/v��
Wr,r!L�r�	�n=�^T���O!v��+�r�p芄���'n�-5�R/�s�;���lX�X\_��p,N�����̈́�m��ˣ�y����Bsg�@��#"Q~�b��6jF@ȼ�L�m���0�M.�!q�ˮ�v�_��(h�ݻ(�tX��+�	v,A�EA�%٣Ӑ�&t�O2Q� W=�ߥMs,�����v���s!k�|�6^5�����3b�y7).�_k�/3b�{U�qp�p$yG�d�{n��4�a]�{r�(ހpH\Re
LL}8c9�0�|�wq��B�[���b\r��oW#{q�{C J��®������ꗗ��Uw����ި;4CS��%�~��f���K�P�:{0��φ	�]��[w�2�����`��6�T�̍�O�u�g�a�J���Inw\�F<͗g����
��a��I�icٴ{]��Kl� ��r��X���k.���13���n��c�ή��0�d�u�q6֣���]�����3d�����T7���/�h���jTy���H)VX9;;hC���j�vj���
���.����}J���W@dQ4�����񫒨��lbM��o������4fnɮ���b�v��_YGG:՗|��k�W�zAq��ՅkV 	؝�8)V��1���k�ȕ.Յ'S9��N�}ϋ6���=mg>�o�+�G^�sVl�:��C���X�xkh[�uԠɻU%�kN��ό{���QN�C�j��a�.���U8f����oJ G�
�9]�R{0���\��`��֩oq��Ai���p*nތ=Q��hu�jQ�&2/h3��j���9t4'N&\ћ:r�۫����*wWb�wȊX��9�$�*�!X��h���iŬ|�j8�M}{��J<�T��:�:��������-���u칋\	ج�!V����IR�K���{�o��Z��i�(���ee�#e�+"�����]NK������N\+��|9f��n�E�ݣ��tT&R���U��l:`с�7�������tܦn,.�>���ًhW9e;��gQ}� ��n��M�3'��J\��d��͎��E��c�����`���|*R囮W�i�_]�4��\F�$��P�J�9)�P0f���k�:u�������]ZMwM�׋"�Yw�xi��P�9���&�7�ِv��.p�x�U�b��mb�Ofmr�C���&ev�sp����ȦV}nN����UL�Qeg"�H��ObR!v;�+�P7yՐ�t8`ac!�ry��t�j��W*�{�ŝt �ݵ���5+q�`���Ŕ���c.�j��ϥ�2���9�)��M��us�����W�ɚ_Y��v��t������Z�r�bpn�^Bn�i���.�ɏ��eq�yR^�_^L�v���M����P
�}�h�W�N.�q��=��u����{5_Soa2V��AѾ��n���$�-eF��=�����:�+�\������u���b�أ���Q)��W�:D����orK����9�pgw7Ur��,�>�5��Eu5�\U����(��Pp֙���:�>Y^u!�����%`�-�)�5 �9�T	���q6��ku|�7�{�c��|�I�vt]Pj[���t
�gٍ͎7�w�V���۩Y��I!�����FP�s�}:�n���ᦣ�0<��7��X��@��*EZI"��ʂ�D�G,*D$����fY)ڬD�+i'B���
�K�{A.PREғ4�A$E
3D���3�E�]4�$ΩT��*�Fh���"(�h�h��EBi%���A��\L��$�DL���#K��t�1+ib�EiE�Nu1Eba$%IRi���RI�	��(jG
Ε�d�W*��ww6������L���Ҫ��TKRDčVPi�rP��$�j�X��WK�Y&�(RW4�Vp�W+9sA*�+�ubE�H�.j�S8Y��V-L�Z���$[Mfr�DH��]"ȹ%DXET�H�AʨEfd^�̊�1$��TQAR��3�Ț�H��)&�d](�QL�.\�I��9�T��ʊ,�K.i����N�%�L"&�D�U҉+V��	Q�rnL�J$���
NA�(�&��H@|�
�
əy��{��Z�����_D�l�n�R�iƠ�"�J⌟fu �����xʄ�v�$¢� >݆��������[Z's�rn1,l�xv	tS�x�X6tЀ�wQ� �Q��\�0���
s�33�{�*D�{˳*�Z��_,
�ܦ{�CY3�.��w�D@�ə�ɽ}�ʡ���yG׽g֧&��q��7Xv��,�n�1�Hq�ч�������/��yZǥy7J׽��Ļ<��0{�h���-�R�OD�1y�zq���	������.&3=���)�'s�IQ!Hp+�=[��z�TWGt�t�!�R$FU��
��5�I%�Q�뙲-t�D�#`;�1%>�	���B�^[���)�dD�o�\���N���m�U�v_�����	�^o�\���"��1�G}��O�x\�J��P���@�r61�^Лמ�c�ݭ��WQE�F2Uï	
U	�2��	V�U�i�#�ȥ����Rn�=�뵙��&p�~n��>Vaų�}A�L��@b�"���PDLi�r�Ga�����YU�c�I�]7���[�=[#�j���ڽHoܺ�MǊ !_%(+�:hd>�������>Yort���D?���Ybt�������w$E�k�r�dR���Zk(���{�4�2����j㛬c��1!�
����	h;�>��+�L�$Y��FE��ѓrf�-U��S��R�/�1��\0#�S=��mlZ9�l��8����z�wt4����N�~�4}66�f˕�q����b������0<��<*܇"�ܵ�Qm^𦮬�GF�Ͳ�7*:�'Ȝ��P�@ U&w�P���������j31�u[j�q涧�bӌs��N�iuƠ0�<M[5��Z��歟�Z|M�Sz���L>���5I���w��K�G���{�D^�T�P".��{Oq;5j���,4	���םy����DH���ŉ�z2]6V
u���ӣ~��T頉���Rΰ}����o7���ؔhu�D5�:���0��s�[�9���V_�ˮ�7���y:���v�z�Tmh�6�.�RB�ZBQZ����ONz6���!ʗl-�-r�p���I3}가��v d���B�S(�:�i�S���9������Y�3{�)I9��o5���Ƹ�|���'���l�5 ���je3�v�Ӻ��!bq��N��K4�FC[�i����%ǲ��
J8勿�\���zbur�Sl�kpM>���S����h�C�>�@:g����r��q$�y��N N=����M�Q��z5*�>������W:�ۋeN�G�<�a����z����-�Ngu��V|��eq�����m�R�Y�v][����f�S �n,���o������5�(����U�>�.����sK��븛��6=ϥ���$ff�;'��n���[�֫������l�J���F� �V��D�dd2h6�b-�4Adp��:s��u#���5���E�,%�F_0��!��ӄǳz�I*�R�4p��1$�W�y{98�U�no&@��p�H/k"�����+O ������d�s۱�k�Ox&�y7=0�w��e�W��**�����N��mm�����.�Wav�k�����K�_�:j����Ʈ��|ɫr�n��C�6W�"�.������"��i!=��X0���Uf�vE9ԕgdS��9��3S����ox6U�<�����3�g�ڦ��~��ʱԏL�����Ǩ	j�4�eݵ�:��-K�!��/϶�C.�b�t�������J�����F�yB|=����<+I܁1��� �\J�����F��e�жZ3�v��c��&8��3�h;A�:�oî@hߎ���&��e�ۿ8X=�ܪ"�-��7�^EӘ�rk��Τ��3��F����Y'V]3f���R�SZ�2�T���׾�-�#�|.�S���K+�̍�
�Up��7�j�š̮P�>cj�����V�p�X3�y�}ժq�k������8�&�c)��Tkh�V`�2^�B�X��vO�UUU}��ˉM�����R�U)��^ + ����i{UJ���4������?��У}��!�ع^h�;���Z+��Z�zxh��)� 㢸�p'V�����lea�k�l�ZR�7��b���d2�>}�c"�	��M��pHGI=T3���w_pJsY�]��y�\b���GJ�����uv��S����aޮ�����G�l�!W����ѢN�(��X�{��Z��[�c���)���Q��"#4:�mh��;*u'�����3-����Q�[�iy��q�����$Y9��M�Ք��@b�Q�w��⼏M�XlAP�I�_mI}6	Bg�T��#6
ez7���%����{IZ�'���/;q)R:GxN�(y��>$>��Mo����*�A������^\����5�h�V�x�s�sݻ1O�xԐ�td�N@�b˲�O����Ӫ]��}�$"V������o3;\��qѴ]�E�N�E��B�H�	�l}��RFJ'hzc��g\�Y�
-����Yt�#��wr=SM�'&��>Ur�q��,�[��z��n6�Ӵ:�LB�I�y[��Vw�,T��ү�WjR������Pd ���$	%�zn�z��ӗ*�9�m���������	SuuJ,3���k�(^Y�xx  ��x���Q�>�K��{r�>��n6,a�.-*��'C�<�gyS�dhT��+��۽p^;j5I�G3gv���Hߨ���C:S7�}n0I�xKR�>/�D�>�Oٍ����s�W]�>�����>0Q��!X���f��%d	�}a䩮e�z��#��P��e�}<���]7�����ٲxK����K�؟�{U��t�h[�����Y���ޙ���a�|�Ĵ�����gQ�q��\�:�K�%T���í��ٽ�J��ۇ)߰��y~m��s�S}K�����)����u��=�wt�}�B�bM�U����!���jߞ����M�O+���M���@�{�V�R�@���J����ER��JS��km�=�}.��.�en����̩LE�s�����vJ�T�|='Y�X�ۭ=��8oB��/I�8�e �ھ��^K��[}վ⺀[���,��� �Ú8K��2i���fl�u�ifG)ו��g��t�!73���j�"Й3���;$Պ���;��t����l��ܡNЮA٥��2�Uc��(vñ�ik��|�`u�8�Zb6�&v^�Vy���3{p��'s"�WI_�����Cs�M�M^���7�`gr)�v��eS�J�`���Z�Lm�h$���c-�4�1�ѵ湫���\;�(�v��g'c6R��{�k2�U\��̥�0�C���I�L����)ى�lκ���f#c{��5sܧo+�ܳ|��n���ZjM&IOЧ(��%o�v�����h�al{>���V�ER�~���^�5��f�z�,Bl|��� 5ڦ��L��)g���\�>���y��U7�/'�nt]a,݇�S�$�N����������7CP�t{�w��(���]�r�i�/���˙�Jt����T��[�:ͷ���9\�2�W>�]
�\��N�XƢֺ��ls��/�E|�`�ڱ/�Sν��)�tOs�])!��nm^cZ���9+g�\l�x[�y��m�uϑ����P�\�7y�­2��9��I��Bf����Cѧ؂څ{�5q�q����g�WN�W[).z6�Э��Q�қ^�宵Cs�>����t���,pooF2��٩�(s��� .���;���{d3�ŏ��J$�`]��.��rF�@���W�ެ�ܬ��5�8���#��}��Z�R��{������A��w��!�����M�EC�-��(�II�Fy�>i�o{-ak�^��8��[�#sVGe-�~.� ^ސP1�!��P�z[�_���>�Y�`H��0��Vֵ�Fun2�uI\\)�{zA��3�>�N.�"��Ks)oI���v������׹�7�m��Y�aH�$'wiC�rtF��um�::�P���S��=��ť��I�l��l��oE;d��H�ޡa�k8nE�u�y�)סA�z�����t�F��x6��X�"�E=��Y2��/:���J�u�hAhuX+rh]'�`o-��]���6{�6fx�R�=^}�]��'\�����2�=�������)�e<����3u97N�'�j�\�o�b3@o*�ὧ�g�ե۞K��[|���矪L���&�ۘ�ƹ���!_q�z5[z���u{�0R�̠]]8�H3 ��ڂF�[Z�Č�Y�M���Q�l������,��J���;_0��{@xv�b�E��4𾖦�i=�ܹإvwOEjӮ��&6��Xᢧc#�}���������Ǚ[����c����cZ�1��T��ױFex�H+�,Go���+��9�:���{��+EOVR>�#��ϻ����碚��͞܃nv��T$7s�8����#˪n}P'��������R�u�5�C�r9٫�����r��~n��(��D��`�A��o�����k�{��MZ�LU ���h��=1��-i��JP���=�nM��C�g� ��]�B>Յ�j��x�y���޴�m����M�mȬ$�����+Z5�*��o7��ݳ�2��g<���=��Ol�lT,�؎������2GgJ����8r��Wn	��皥<k�Fuo�('M؋����6\����������f(�B]w�u ��ӗ�`#�����n6B�al�;r���.���1r�s
	Kb�-wйf� �J��n��eZ��Z���dcU�/����U��4��S劽9g�F(�uP=��vH�n��G�<�[�k�.T��&�V��I��o=��k3ޗ��DnпQ�3�Ў�A�^W�r	Ї+�Ur؅͎�2$)M��Mt�Go��KRf��JN+�_��{� ��IB��ƍ��`UǢ'�ݶ���̕T�{~�-�Y�p���xM�rY�_ls�b	�+_`���y?���y5�~v�[ɜ����m��T�5䓃A65�,��r�ȵ�Ť�_��n�S��Sym��I���u�.�\���f�lF��-~"���:����<��$t��X��OfWR�����c����L3V��X3���M)�sq�[�r�\���d�-:���@M��J�����s�T�����lS���vn���	�<����C�F�fQv>Ş�����������;�`���d���Хy����5!�s���-Ч����n{�^uzt�&�PB���n�l���Q7v\�_��gD�{ϵB����ƭ�1]��[SBE��S�v����0�\%-����|}���a�Ў�wmu)�,xQ����RK���C�݊S������Oϐ�j�+F�+�:����oҼy)��O�b]l_-���u$w�_rM��$@��5ǁ��̅;.�ݳ�v�A�mT2�Y��	�p��aS'���G��%��v��Wn�)�z�J�]�T���{��ױΊYmr߽n�꡵].µJ�kyoa����4��'�oC���Z����ts9��B���\�IK�î�R�QN�P���{���[1Y	N��팋�N.���������]j�M9}ۧ��ê�+gZ=[z��Ϋn1̩�aO{z|C"بNK��E��ht(wX�6o�I�x�r�3z�3��;A�3�aOL$6,����K-ʉo�Ea���#ܟ��W��j\�e�;���(�Qڃ��և}i%��]��_��a�^XE�Nt�C��4N��5�G��*�k<ż��������]��U�Q�|H���j�����5'�-0�lc�Y[7ІJ�[<�=�{���V�0�������)k��[{6�'Z��UK�U�u����7�OX��֝���xn���o�����M�l�}��������c[	��7W�2���0�Ʒv`�Ź��s�Jq��l��;z�ٽ}Ah5�ݳuo!Ǻ�c��W�Ag��BA&nqq�'
yd�Z��O-Ӥ�U���kl�H����bm
���r�]�hfō����8�:U�r�ԱΙ���Ko	c[߇iY�3�j��\�拑NvӶ�n:��C9��e��pb"�j���9��>�A�� z/�23s�Ef��bvc����7sx����GQ�\gN�i|A��s��oC��r�I�h}�s��Ao]ť�B��::9<Y%��=e�ZǇ}���N`�a��!<1��#��Ԕ����Ք��VC�<�7���P�Y!�p�+�+�}���"��Ī����L�3( u<��7]���g�/2=����rr-^w�V�{�Cv�����~��� ��l��1����CJ-T�X���z8�Ղ�xώ����v���5�ϲY���T���P[�Y�IY}�Mٔ�e[U����:�6l����h㨟��ƴjb��Ѐ��(g]�����r�>ɠ�(��\�i�^�v�<<��A�Nl]�9<�]$U�U�+�F����	�ZCsp��n���;�{O7;�Y�XS6���m�h2>�;�ʨ�ήv�j+�����<�n����-Eo�����D\5L��ZB�N�]'�x�yQ9Ӊ�8�k�ɧ  �E�d�0)�y��Β��LX��c�̷J�ʡ��z,��\	���̉�5̧�Hk]�x�:ج(�1����n�9��Ө��x$��/��gZe���c=8'�M�W�^�n��	�:o�.�V� j�1SJ�\|v�M�#�b�gv�0�L1��b���;�:���G�էEF��fTV��h.�}�}�ӭԻ��KF檛�{�7,�W��4t�W�*��c�]�БxE';cvN9}s�.��\���U�F�W=���+`�Z�D$�,��Y�'N��Z�h-��w�0�`�:�T���B���wKc��"����۩,k�t�_U��]H-��E��'BR�E��D\�ӾX�k��N�˽n��7�Q�R#
�tu�ǏQ��������B�����+]G��`��da��:J���i8]�2me�W;�et}�� �w,�D�yi$�i{}�0p���l[��MGK�9rH̊[=� ��M��y��
����I�
�f6�"���B�l��u{m�����wiU���u�#��K�_�T�΢�I�;5�+h�=)4]%��%\<����)b��$�x�nѰ)E�X
*�.
��J����Wt�GfC9p핲kr���܁{�؂��)����R�]��u+Y�L�5��B�6X��^Y���5���˃�[;����-s7�u��Z7ش��/�Il�o��e�s;*����Z����t��h��P�3�֧f�^��d>
��&_;B���]o�;�n nN�p���EUDQ&J
p��+B���a�Y*�츨ʪ)D��Z�a�˄UHF����3eV�VJHEpNhtF���BPI���4�P��At����NbAp92�A2�ÔTQU��.RW)L���!�lȌ$�Vr�(*��S��U��i�
��8�(��UQ�	*�
��#�"$��R��r�"4
L��ER�t�d���u�"��p�*��uUI*�L(E��v�2�AUUBE�z�.\�C�{��s]N谈�'Q�,��;��EC��\ᒪ�u �.U�Ӯ�
g8�30��t��2S,��p��̹J��Nf���Hs=� �.^Ek1 �����Y\JԎ%q�Y��˴�ġ2u���fE�fr�E�t�H�JB֕'L�3�UJ�˜��N���I���O$V�N�+��U�Y/��j��M��gn,��d��e*���h���ݖ8��˙(Gح����TJ~�������m��=;�����M~�Ox�u����Ip�C�$�%"#-�j]�j�n����B|2�;*S8�;
u]�D�:�_9Z�󛙷MW��[�b���p�:X�_.� ���=-�_^'����M�l��8�Ob�)ng�T�v��k+��0���^[��M����w��1U�r���ZTq��#g�)�ʤ���
�����Uy߼��̵tݏ]����LSwԵ��9�Ba,���(|��R��=]]S�.�/�)i��6u����Qۋ�p����.۱	{{
GtO����N̢�X����]�,s=��F�������m�S�HT,�{zA2t;0�v\��s9j�]m�+�k�9iXg5�7��f�f@FHVV�y��X�f�k�Q��%���I4����qA����^���:*{[lOt�z7kj�H��h���Е��W�e�ȍ��$C�R-�����-..�&���S4t}6U��7)v�3-�V�
�Ζ+R,l�0Քu�XuةV��ܒ��\��W8*o^����
ĝ���1+/6�B����W�{c�sɣ�ٖyЍ�^��+rhn�F���כ}������h�~U�zf:��[U�엕5��)Ў�nM�y9��=yY
n������B�Sj�����lk�!NV�1#�tŭ�z{2��}GsA��a��,;�k6�o�i����6،��^��E��H]H�J�y�m�N�U�T�_|���]��7Z�^�;�R��&5߆9��Kw�H;�Y��LT�nq�x	�ܡ1eM���/3�����R�,4��j�5�nY;��/��8��^�_0�^��C���M�TJq��_.�<���x��)�Ǐx�Ow2�1�)OVF�an::������.z��j�k
��mD�
�-��|�ܜP��=^ؙ�]��}�sG���>�\;����%WDj�OZ�ٓhn����m���{K��� �>Xt*���yuw$�G�+�����
�6���/7v�g�W���r������Ȣ����S:5�8&ݩZ;y�Ծ�=D6�>�����w,�/du�gP�a]�Qvwz�뮣M|;Y��Ac�84�K��w��Kʻ)��g50@�Ӄx���Ю����{�Mk��if�]��*����Tז����^{i4��VبX؎��29wr��VR�k�?C؟����ʖ�)O,5�s��[��N� ��lK�avT�)�����ǁ�{#�]�+�-}5���u�E�5{�� u�鎈�D�D��s1K��#���[-w~�oFhI��R�8��5��+wq9U�}p����Dq;#��`'��Og����9xMua������CW��ҒА��v	�Ԏ�c���/s�\�/F;&1�[�k2�N^]4�����4N&ƻ�N�1#�h���;#u�eZM>p�n-]�';��Vr��|�L2��s��Ɠ�X#&l6^��T�v�B�1�������S�������cH���,[�w����W=�ݖ�xZ�w7�F�����P���܁=����C���%�6�'��y�S���n�3���R�91���5x�^��X}�O�	����"xR4_e{uyf̫;�|��� ��P��D�����C�)Y*rtAU��*C���^��r�����];���Pќ�^���r���J�yo�YJ�%�f�磌ﾨ�{2.M-����I���P��ֱ�QW0����nZ����WJ����\;3S�D[�9��1���{����z���*ÛY�M��R�;�Ӎuyk<�S����W��!=ڔ�{һ6�oUgYڧ�U��<�Yb��V}1_��Ep�E�sO��{z�5b6Z������[m���XS}^�{���7<�u�mZ�+;s��*(ܕ�6�JT�p�o-�7�a�&��R�'����;��6�r��N*��r<X0���ݩ+g}=�O/Z�`�F��-�|[��Ȝ��~��=Tc����Ƭ�ey{z|P0�����K�S�"��F�q����n*�j��4sV盌��ey�)�aO{z|C>��+П\��c�_G]*pf涗]����W�oZ���P���t�CbvLk��h?D��ګs�r��=���͋�o�e�;�<q^NĩG��y�9��cqtj-��,�@������󢫬+Z[�sb����;d��Z����D��q�̖!��]� �8ز�o��H��o����Ru�Sz�7S�q���<V���#a�4s�8�L��}{l�V���b��N�ܻ,�ړKc�z�E��W�}_|���s�}|�n|!�O>������-f�Iÿ2ƻG�K�}�粡8�rUF1Յ�E���=i�=�i�9�R��8oϼ�n?cU��>����ױ1Ӛ�۷���g[��}����*ǈЯD�Թ��f�M�h[q���Uxn��/n.����u-��z�����3�YO����oUt�]>ۛ�ev��]ih��g׹-�]F��!~��בZ+ҳ�}<Gg�~���O���Hʝd�׸��^O;{�����5����/_.�����7כ����L�
��������Y���e@�s2�X����P	s{-�݈�B�06����ڽ|\����մq��l�B�����s��V��mJ��6�e�;c{��W���\��nu��&Ax�����	0a���]�|���w֖ڳm2� &����A�hP ��B���ׂd��t���kEG��w�o_�Z���Z���sbZ���ݛ�r�^R���4k&i�\C�3�u>��p�`��}�@�Ќج��t5��}t������9Gsv쮳cx������`���t��}ݶ�����]�qp�7��c��zϰ�s<��^�xR��^|�n��:�9{5�)儵�}�� �%qp�����:�:�����;X�؄�ޭ_P_8}�-�Kr)(�Ď[�i�U�u�a�՗��b|��,	磟����ލ��J�:ݳ�Ls�F�nL����;�zn�6��0��yM�=���[\彮��h���3�`�!���)覎�a:���R�sWI�������d%�i��r�sݹy�F�Nlc�B���1�7<"��;��y���Y�N�Soj�3�N_e0�my�b���؍��k�:�-0�svI���c/U����y���ln�^��w�����1��*�]��>�JG8�r�Գ�j1�k�}S}��E��R[�`/b�OZ��u�s}�#[Ή���q��S���O��r_˹�+���zL�";�x�X��M6Q�}ks�u�l��㨳�����O7lfYQ�9ݜ�5��;���ޮK���n��%��()َ�-lE�;ݵ�w��P��,%S��Ԯ�7Ү�k�on)|'��UU�͝,)һ��vm�]�=sH57^���g�OOz�`��I��n>��'S���Ρ�<㲊���^�3���V������fc�#3�y7[�����V��o�;T7dsUzK�h��O�U��0�~|�����������O�������g��#gŬ�6�˭V�_whԱ-E^?I���]�UAky~{彇����ZȞU�*"�>2�F��֤�Sz��X��*[4Rh׻���j��7%n�#̣Y��/2e8�>~� �c�E���غ���N_u��>�S#�+�z��V�����_��m,�F��y�dg�sw|WR�Մ�B}ef\D�B�8����9MԳ��E6���g��HlCӢ{72pS�{7Rŉ��z�F��.��5Λ}�8�\<�HH�A�B6�����J�gx�k�,:�4� P��R��W�b9�m';��$�o������l�D���G�*1�D3FˆO��\y۪!}�����pXi�;�ͫ9B�O6��]*��AR�/D��DR��jV`+�51Z��C���g����X��7�QV��B+0�_x{���=|�VRj����d�jT8u��QI8�cXV��C���>�2���D�#��s�O��os/'7��۹=�'&���>r����B5ǹ�hO[Gp�d&"�j1IWu���w-�^�P�oo��'�6�T���.zd,o�{��ܥ���{m.ʦr�y�н�j!����i�TO*ڞ	�Ӊ��KQ��k�Ѻ�w ��	��u��Rc�Q:OW(�x}=���Fv������o�k����9Z�2�C��޴J�OPB��.ֺ����g�b{�(�+�\��o+$�Ӎ�r�U�8����x�t�䘃�o�mpj�-X��PZ�[m�uϬ)���{��HL�;U���Ei~�r��w%��U�������o-�ٮ9rdda�S3����}Ld�10�lA����{���EҤerx�Bш�=YlK��/)��Do� ����}-e�*�܎VJ�-uf]�ү�s����+����{�2��זc٘���X9��u�&��ivLX+L���� Bs�m��F�Q�{\o�2�TB�<s�:�g+�<��!P��z��si+�=�Q�ӕ<�59��߂�[o�S���p����}n�{syU���6��w{�g�s�A�}�q�V�eT�(;~ͳ^4;�*i�Fm�g�R��v,��d�+���SJٽv��Pm�����J��!�C+���;�����ݛܟ?2�����J�&U��C,�!�\�5mOjbU�����������Z�$�7cZp��96V�Gq�W6CA�`����@�`g-�=vj�!v�7�p���p������e�ѽb���O�h���;U/2����5��9��Bv���^kY���ʶ�&�m��o*���1z.������΢j_<�67���[쭎m��t��cZ�uOr|��b��<� �47p�)�����֟�x����T�e#�����k];S�d�H\���f�����E�ٌ�p��$��ڬ���L]���:�J�A�+�GmJ�x��ZUkʹ/���S�Qw�X������F�]*�ȩN�$�.Ă݃�b���2����H��.M��wX*8)��s5ۘ��ui�g42��j̤�	�<u�R{�mL����>���s�><=�i���g��J[p=�1{��Ht��^�M��o����h�o�����GH�B3�;�\�֫�[���[8tl���b�{�<��މc����k{]�(.���؍��D �����k�rBs�E�b��I_��a���'֦��B��oP��N߰L�i�ϥ��f���H���������|�˶��p��(-��W��-T�&��|�J�`CY��yJ٥)�X֯ѝ^�.@N�::yZIB����,�?z�ۿq]Ak����7��lU��i�VVm�ik���DS~n}
<���v8��-��I�l�bЫ��4֩�T�#�ύ��Ţ��(���B2	�愭���:z6�k��b[�:�;Q7<��8XB�^��"��R;B�ړ�殓�~`�=0��������3g�;o-�4hN<�t�3)��������.�
�x\u�jj�v�y�n�¾�Ŷv7V��7f�_4�[�|nDa���}���7�����v�VV�f��/��7w��,����X�nT.�j�:�]ڐ�Le���i���ɷOj1uf8O��ڗB�*T3�:�d[����Y�,�a.2����*�e���|�VƸz�СBu�v��Z]*.Go1P�u7*Xa���aXɫ]ga��p�d�%TO�q��7�۽ob<���1���]�G���������۽��{z�7����&��V�m��/��HU��:H���>��kx�ԭ���C�G���͇.��j��t����D��>�zlv��&ۈP��g�@SM�֒#eе0t�  �V�}�e�j�F++2�F�њZ��aQ5ѧ�	|k���>�ED�����<����>��X��WzN�\Р$�7K���vfa'�Sx5�I�J�b��5��� _q㬕z�#��78ŷ�X��҈��"Jgu�ꋬol�a��y�nmH�^��/)-�s9�����YX�{�t��C��a�Ttb�oj��uw|�e]����7˺���N�A(�#�M�}�:�uJ�{���`S�8����K���*e%:n��C����	pmrK�ԙ�擤C��4�E��hN �>���9X�c���j�>���T���Q��_^�(��16��lըJ��]�5h���O_]t�����{o.�����z��mY%�9�Z	���֩��b9j��u�u3B�M	�kY��{3���tP��3tD����k"��Gy�Y��dsi��X���0��V�Ջ.���4jKkw�Ap��j����[�qel�Y;��7���	 �J<��[����,�E�x+V�p�Y�QY׭�le4h�3�4S�2��Q`����i,L-����������+d�xk�}�����)+\[i�!AbF����/��XL�7���Z �nw(��uo�KE�7/��u���Q�ĭRN��wF����
��W1�ga��]nK��T #���76��
't�`�Xc&��i1���w�l��Έ,G�6t`p2*Q�xb������t6�h��V�a����<n�[���_ѫ�c(_���$��M�f��`]M8WT�U>�c�tuv��md[r�,��M�HvPPξ��v��wI��q��l�&�$�x�*<�ܹ�ߵ�ӗB.�1ט�����6�`�O�%���{�J-���µ'z]D������E)J��i�WD>jT_�׺&��e�P��(�yåMJ����o�����7NS��Ok	Ԧ\f��Ds��I���ʻo��eH��S�wI��JW:Y���z��^�VBP�t]VVR+�+�8!]���L��+��C+%�H�e�ԑ%L1��2L-J�HZ�,�L���t��@�4�-�)"T$J(M�^"r�b��TNʕ#rq�Y�[����C;�E�:��Vb!�.�$]�"�sq($��B�B��K�aZX�Vj^J��*t�r�ۙz�D�B�'7u̪�D�ܓ�s�*u5B�At:r��)p��ZiB&��-i蹁�]eDE�ZW(�!
�Ą)��99	�D�z���v�E�G�L�$r҉Vt��AAAww=�rU�����4��""C.V�PG3�!Q�9MөxEx����˺���=�bQIX��e$P"��9T�g�EA�E�G#Uj���%��G,�ܧQg"ZI30������7+�uP�g�9fTDb�Qe�K�{��������)��ڙ��[+�˜a�T�Xy����m�c�����X��;[�tIM��W7�4�
�.���dޣ���諭�j�)��������ʃ}E���lk�Y�L_�F�[���;=�LR�ZU7���I��ޫ�h.�W�զ�؍��^���r�:�k�'\F>V���6��{2����W���R��&z��r�w�s�=��9��trša�FL&.٧�"{#/9�[�eKذ�ֆ#���?f�VH��[�mx�vu���{�÷<�oќ/�
�1D��~��YWE>�i1�cR�s��"�Y=qh���b�^:�b�s��]g%�F���k�/��*��ogY���F.V��6)`���;Iv�0`�{<-���ϖ�Ox��Q��s��Ya�0��j�^[]��I�[U��Z�[���o-�=��{~=}y; j̛�낯4j>��������R٠Rx�X�;T���U�=B�W[�	�+�'tw*��-�Ѩ*��t�R	λ(j�ܼ�=|�������6��u<�����{�}�;v�ǌ�Ji�xFU���x-BM�J�A�Y�Y�a�NX&�]971_[�鳩���H��n�]I�7-/��h��Q��`�ۜ�����d�yëݸ./�-�v"㽛~<����R��^s� ���JO=���y&y��	��ˤ���!S�� G�vE������UX�՛+����+�7����B�$܊m�y�*!_�a*�Azu�ۘ�����wj�"jSGz���i.t��w�q±�J�Ԏ�z��	Z���y�l.�`�ɡ7�47S\����4�qI���`���,��6����(�wVѾ�Jv9Ź����7�+2����д�-��y���1{���>�cֻ�92��8�oE�:�K_`�[B�����4ҝSg�6�^�c9D��!�=�Xs�&^E�ŧ�3��\_g&an�2��ų��r�S�0��>�?w�=��׏����bɹ�F���-�FԪjox:���y{�;k��T��=�x��ͧ׵�6��/�{�!�ي�;[מ��.��?Vz^��qJx+�&
�r��K��MW��ߝ�t��F�v/�ǍШ1g&�m���{��\D�o3�]��VS��P����rV��w�PHUlݱ�*��n`i��U+��HH�#���{�=���ʟ�|���i(̟�;;Q:C{��J.W.�*&}��}x��9|>�״��y����f�D�R���A!��qK[��m�<�WR���39�z��:��e0ݙ���J�z���,��y����� ���g �ގ��ә	��V������L,[a!�P�����T�[}��]B��ݡ9�橴������{h[��]�*/oB#�v�Y���@�wӊ'f��ۙ;�ܾ�	k\�/i���{����^�0^-^��iO>9��|��۽�v�]�V/j[��^G*��p��!WoIB��\���( �)�/Vt%�z6�M+�/��<qI�����q�Z�G<�/��b9��K�5<�j�ܛ����m�37���(���ϻ�L�cN	�'��f
cj�ܚ|��۽����C���`Uw�	#�:�b�cr���)�qp���T�^i˹�bEU��<nJ(W[C��H�Xzs ��Qxv}�V����3�&aFN����j�N�I����uU8��Z8��h�OO>5j�,��&52j2�J��U�[KZڹ=v(b������y��Rj����A���Ч(vby��^~ߖݻ}�O���¹nc[8���5Պ�N��B1��Z�޸��j��C��B�CNɹ峹��S��ou���i����]GSܥTk]���ܝ�!��u�ͯ��_z���@D���B��eKذ�.]7��;l�1�ym�=m������KG�I��TS��_.��7�]����*Q���y�o:=�O���O���0mJ���k�k
����B\`f��B��k7���Z�sל�u��V�l��`�/�P=�s�"�m�'V�U��f�7t/�SO��}~S}Au�U� �}�v�0o�+�-������Q�.g97�CYa�Y\�e������N���΋8<��)�W�v!���-yR٠�<�5�s��-�br�TEj=�o��@����k���7E>��~Q���x�Z\��y\y����4pM-ھ����w�z�7D�=�=ӨwD9Y��9,�F)�6�M���wM�]�[U����ߍ]*^�'�kd��=�T-#9<��\�}�ϸ^L���B���%����Q~��j����L�7�T[w�����_u������2�0�y/��7������qc���q	l_�k�⺂ލ�$ғ�§R����%'2�=��*���Ȧފ�e\R�F��Nf�4��`����KpuK���*�����G1�����g;��R;Pg�i����[��o�鋏$����{�m���4�M�v,��H��yŶ8��������g��o��������������i�y�#y��0���z'�}ܯ�e�����R�+2����w=���a){c��3�w/q�H.x����w6�:��y�̳;m.��r�~S��l��w'�`����]{��ti�L��]�������\] �!79^��q�On =��!���l�����	o�zz�՞];ܜ�-w!��n�Dk��g�}᫺����ux�Wp�##�(F��=ǲ;7��H^9���tk�GZ���mY�����_Ti>�r��n������5�=����B4�m��Ϗ��<���=P�ة�+/����V��h�v�RC)�:�����wCx�T�Qfۇ�L��Chd//�7��y[��捿�4��|�7->S׍�^��)�ub�C��<t3ˡ�G�sO��{f���=QiGd%|�}a�>�7Ժʜ��g����S�׸�N��P=��XߗO��V#[ǰݧ��4���L�7����|���9�`��^��_��+ghwy{�ܷ|��=uq]���$��M�?_le7M�����(!'	wd��O�}c��W�e<�/���D�ށ8�Q{�eWdp?��}#�����Y��1���[K��Is-$�kX;�M�?��&_u;��!�ԡ4�
��fu�E)sٹl�Kz6��>���
���o�;��x��ceJ|��}\�n���o���:�|���t$�;�,b����`��)uz�p޿Q
:wj:��^Ns��Y˞�MQ�L3������)]�`��v���\�,��*9��Y�|]�v�:�s0�r��@�ί�����Ivky�\.A�-�MS<�}�ͼ��%�n�����F��CTH��w3�P�h��(r��b=')Jm�1H��O?�돉�{Jf�A1�aѫǳ������F���V��3=�/)���գ7<���~�N{_��n罷.kz¾�څ�f�M�j�3�������1o�Fb�M��Զ5��F�^�g��{i%9r�SV
��1����=^�]#X9�e��^3э��שvv��~�H�|�M�	y����Ϣ��gZB+?{jq��c7լ��ǘ�����8%�����F!>���{R��ˬ]�m�12���=e�1SuN���=�f_�C���UK����F�W������m�42j&�s,��s�4�V���ބ=�wo�����N�*��C[�N�C��5j�K��������vڮ[Ʒ��F|�I�W�E9�Ϧ0�T���2OcK�MK��ۅ�v_�ʵ��ZV,t��f��#t^�'�*��&����k&gzs[��N_bX֯>���eT��.���Ll���rxa�"�8tB��p�9r��ɭ�ťo�Kh�2�ֵ�:�vbW:ɼ�!��Z�;�QcǛH���iK�襙�7
���.Ď���z=����7��L��$��W��ln�M��x͗*ð���8�����OH0�<�)�{��q��:��¾�'qP��������m+�7�[܎xβɞz�_{�j}ѻ�y�X
��T��ɩ�^�ݽ�2��V��v<q�]o	��r�螫{+���amq��Ӵ
�b���ܫ��t�F��.g3n����N��ܼ��r���GF��J$r��:��nJܚ|��9�qYy�42�W����9wy��ꓴW�'�1�)���1 r��E��v�Ofm]�t���J��v+��K�ܧ���Y��W����xn���k�s�bk�5z�>�Y���zѮ�/2���߆�u{X�){cֹ�yr�ټ/k�ث�gpܜ�[�v_��%�=��V�ꔏ��^F���uf�l�FȬ3�s�'��_�H>�%r��;p�޸�ug�t�����N�C�	�X|ը�E��>���}�~kz��ge�\*�z��=[H5b5��]�Rg��S�<o,���V��))��r���B��ג�i�md�ǈ� �:��K�y���FZ@�э���N��+Y��d})��r)j�*�ܕh8R�\�}̪�'t���՗��`�X,�i�P�^V���Y:9VL���#�_�� ]F������Vصd���V�5_o��TV�u@θ�����<4�ؽ	��u�?)(5�:�P��o/ͧ��I�����ʠ+b6)��n.�u�o_%���&��Qu��<����k,=��OaSb�Eq��u9|u���N�&"�"�L6��]^T�iJya�k�>���F^��r��u�	���̙B��~�%y-�ϫ����\����`ͭ���py�'Q�s�_^��R���v������Wz{j9�o�Ƿcj���¥�����ʓ�Co�fQ��,�	�ؕ����VGz�w�J8:c6-�5Ɵ�tm����l/_�_*��3�v'�n�2=�j�{ǋ��&��U\��kwf���\��O��I�����rc�F�9���U�y�g�����l.���i�Nzi�{]5q���V�e�#7��G^�UX��ZJ����(U�X��\��#|r��2uu�G���`���ў���8"��c�6���M�"b�qv*�*.w5(cX�p�^��S��N���3�[��.̧���]�{�E5%�dӬ��f;���H)�h�ښce�Jb�쟪��\�.W�˭��_��{V�Fg/>��~/S���L3������T����>���RKv�ă�Z�3���>�Uy�ҝ�q���o�_:�+VS�����r�v��^i�q �����yp�hO[�ƣ���1�Ҷ�]D?\�#��w�˱���o�"B��Khq�V[�2�TFZ�}�u�0"lsÅ�ڔ?KO��N��ڡ=rP�;���&�(�gx�tZ����=�iE�	bi��|�v��6Qឬv��꾕N�q#�t��R{��r�Z�q��=���{xZ�Y~�=خ����]�n�GתŅ>[�⁇ʤ��:��@��m��<���r+ke�GV.��kE�ܩ+�\){zA@�N]�+jK����f=���˳�˹��gn7��^��3�aH�wO�ilg�k9�qdɸ��̊f����|+X����#�0a�(k��N�D�D�H`��
�^YR����:�oB�.��;�&���b�ǋN�����F���9a����zTF%�:��c7��y�7l3l�b�e�[ù��*���
��:��Q�%�q��bY0�&���e]Յj �e�����e�`֎s�U��^�|>�Hw��}��d����oM�j�g��������C)�����=�+��c�\:T�Ѱ�W�I�}��6���]@����!ocokYW��)�g:v�k2��z%LE�����V晗y��>��PM��+��n�?aQӣ�XE�
�Ϋ��S���Ժ�U��[�=���roU��̈:}�s�|(*ج�Ah��!AQ�n�]s�块���9�R���3��;���w%��[��۬��i��!s6��]�j��p�_44L;2���p���q�ťyD���c�ӁQ[ݷgo��[1'C���vx�2�Q͕���KC&0@��ঘ�����2[� ��]i�h���Zu��&�َcDsͭ�ο�[�7��I��[���k�3R�Q�;49���Ev|�S2���3C�8NᙛK�.���3\�P�TU�'�:��3�6�Ҳlco8r�m�@~R��.�&1-�r�v�_g>���ט��:Ii�Õm*�u�fw�b����u�;O��=��k4�u�w�I`�Rj'C9Ei�ٟ��'3��B�6�߮��v;��utav.�d��P7�u����K�%��Z�)��cƝ��ݛ��e"�Xa�����Ba�Rf�Ե�d�Ⱥ)�������i�U������a��3#��*:��0P�y�e�V�Ց�߰V夒p��\��*�s�25ܒb쭘�]�jل����'敔�n���ɶMeF�G@�oi$��^h9c8)k�U�jMI�(�ܴ�5�mu!(KWK�ak`8����˥�ޣH`�C����� P3���U�Ykh����v`�4�YI��Ѹ:=J�8���>���`[�MVN�+��x;\J���)�B�T�eB-����l�]�7�^�?n;�]D�����jn�FXR�.��'7q�6u�͊��J�l�9yK�֍�J�-��
��3tPJ��S�#2X���,�D��-4�ZJk�V�i�7�7�ր�i�J��-pU�b4Ռ̋"���2����hL֜�P�0�<$+s�:�U��h3�1�q��\�Wl���#�坸�_>aK���ۭ��RoK�
��b�V%}��g[I�X�/����S���K����c�e����b�k�k�K��ʝ{P�!޾[K�qU�����wd�fO���	x���!�[O�Ɩ���
�rŬ�e�QI�3;Z���ӛ�2'wS�LXw��*�]�Ȕ���j��)w1�x��bX��W��#��B����N�}��9,�
�+�)^�P�J�*P�8^w<��)"�VE\��9Y��&Yҫ�P��E��hgKSC@�s���E�����a�DZ%P(��P�˔h�"8\,U����9� �)�g;��! ����:Th�T0�J��eS4�9t�U.]�u�Ȇ��<��\̠�3\��SYU-�e��ZY�49W4�W9I�2PDQg*���')��SE�VjU£�%�DW
�H5���\�:p�TU%BƕXeT���.�Q(�e+)P��)&��bErNYHQAg-D�T�Ke%Q�"#�q9L��h�ȩ�b�T�EUª��Ȏr��a���r"�*��r��$�D��
 
�V�·&_e�VgPĂbf�Q��:�����{��Ax�C]6�;f�����r��#���;̫�]fa;���(s���������"]��j� "�y�w"�qx��w!�sC�d#
}�	ٗ���2��3��[0�w%o^�qJ��m����p�±�����
E9�Q_)�LJ�ު��J�&�eh�M����	�2ƺ�����@A^c���W�"���u�#�G���O����݂�zFa�c���"��V�W7N�����~��ǿZ0y����Nj �\�g�eN�g��ʶ�&�t��{U����>�}Q��m��\OP��W��6�v뼽�m�/k��/c'�z��fӴn��ex��.��� r�$��D�7�s���{�祥<;�-�)��x�Ӭ��u�g��1c۬{cx7�iB���b1�g3�'��j�VE���}�~ΝlO��sv��)��/gR��m�ڮ��.�A�R���-X��R�oU�S�Q�H�ڝ��	@8ᓹ�\��9ԏhniν�lw���x�n��Փ�����vp����V�Wtz�_M�s+���e���PG'S���Q$�@vR��C�Vޑw|;(���w`�ם;wJ�*�tѕ�4�s0��7�ӉcS+_Xs}^��
؍�y�T$��@��{�P�WDojvv^6�QS����ֳ��I�5ˀ��>[�P C�R{�]�B���{L
sCbkܻ��*��i��kB�-���v݈�K��⽹�X�jS��5r�=}}ϔ��x���t�hy�촵��>����A�%qp�O2��*k����61��֧Ơh��qˮ����m$����#��wTpX`o�f{�jB�-�=���#��^������B]�-�ԚH2�x(��]�vf=+;�7�h��E��!�\�˶��O�n��3�P����\�a����L#�U(�Q��ېV���=����ѬYM�z��y�w���ڣB�pi�5ߡNP�f'�tŭ�2�t�~�zi>�
��gw��0��V+�m�ж�m�^��;�[^��gl���+��\j�Ws׷Ҭ-u���;�/�ͬ���񼋩%rcWtf|o��_Y�n�`�y�
�X�m�׷h�k��qӛ�r�Jbr������V[��1"`;�&8`PuV�9��ir�bB�I��+���,�;�mv��s�i��ά\�_R�ǔ���	�Η��7S��z�����k��%\V��Qgj[�Yy��-���^9��m�D����'-��Xb���+ۯ3���Q{�\Z=�H;S�[=���El.��/�M��@*��~{�D��rb'~Ƥ?{���9�R�=�����k�^>�s��Dw�"]�����#���7��m�uٷ��;U�><��uA�Oi��nBH�W���c
�������Cx�z�'��WB;~�v�Y�������x�q����N�ڢ뫪y7�CYa�=�Oo�[y�r�2X�\r���O#�ID&�atH���]�l���ֻFq*��M>�C#!��W���E�����H^ސP0���գ��Z�h/��9�}���J�c>}x����Y~����|�R�<^��!݂���Oo��InǦ�w͕0�	ym:�X�଎@�u��d���c�ӭi�N�]�t���V,V񎐔���ꚴP��-�on�Z�ȍ�^�*���yy��IЖ�U��D�Po.u�k�E�6*�k������P�jZo��l��)b�y|�:^S�A������G�<�N���܊m�t�#
@�HlX)�����'��7�n��DԦ��=��K���C��8w*/����[[C�޼�5g1��NM�q���d��{^\��	��I����	�F+�n�S�1�徚n��N�8Z�՞�˜Oj�V����|���4����O��j�F䤮�F��z�Y��Jmg�ک���y�z�iK�:{2�p�ʷ;�V,֔��,-�o}m�Hc���1wΔ����ʽ�);+��hJ�&iO]+�$�ט��`�i�X���6�Wf�\fW���P���qZ��V���o�U��k��E��ʞn2^.�&���m����U��e�OU�k�Q�,N�Љ��bщ�%�ŉi��Wf�x�:Ϋե�s������z�J�����U w�$��WGu����*#���i��\���ۓs��!kS�����\�zQ9S0͋�z%�W�%R�[*��u�|&��>�� U���,�s2p%����"�rQ�� ��iE�"3=�I[(b�EnT��v����m�5v��)�&`}�>�{��Vr�aөM5��u�LR���2�m���[���{އ��x#�@�1݃j��
�+5����8b�uNi�.J���v��4�����C�q�}���I@��BJ]~�ԭ�"�t�˸;knju%�w]�����19o�\)����$�%�r��*jn�E���}9�����SA��#�����e(�F;'�e
3��-7�c+��J�i'�F��W@��a����jZV�kX܊���(���'`DN��(K����8�Z�Q��ǵMz^��Ū[Ѵ�̾��AІ*�)�B*��-��&��b9���mvՁܝ�����"�v/{B�%�$��Ż�uV	��8%�1�7 ��w �̹�{W�յ��^M�f+gb��)ދ�|����hF�cZ���p�>��}^��^�Z��ָq��zz�ms��T�5[r���4�;ۖsB{U����1o�bԈ����md�1��ٷ]c�`��љ�{���+��L�LPB�%��~39&݂���FmdPN���W�=A3 ��d�kP>wPC%��7�8f�;r.�6�9	z�hmp�F�U,��Z��8�Ε���=�4�"�v�8�F�"�G���}Z�vEiQ�-ko�-Ę���j�u�k���d�fם�B�,IBP�ua
�M-�2��r��Bnr�WFX�BF[�~*Sq��u�:Ϳ>���Zh�f��*��K�����qv��T7}�'���*���V/�vzp"Oj��)W#��ѳၥ�2r�}씳��g�҃��N�����A��R�x�ڠ��.�-��Ŕ�~���B	��C��U�����}L%��;ʽ|.!����\�'�	+�@ʠ�Q����,D�����U;�m���UwwfQnuv|�K/<��>�C�Lw�z�/d�tw&P�aNwF��wK��/�9�k]���^͎��������\.V��Iei��,�ǟ\-�u�_��(�( o_,���c�v�.׀8x�{���Ͼ�n�Uç|0y-v��>���<��ˈwv�(�O��ye7�ѯ�8�i�= ��:~���<�}�2�Z�|8z[V��s�7��c��튍K%�r�^��t�l��R����(�q�:Ls�}Eiy��P����F�I�@��:�K�Y�G}���\��[�kr��|�>�9�ws.�:�����s�Ya@'��{�
�Z��bOuK����j��põ�R�Zxn7����ν#+&NJ�G_*($V'4F�d)b��U˪.��S����x��t�D�V'|�g_f�Ж]mt��죞�����&�%�su�[�q4�\�@!#�d������\�;^���5��EȻ�z�u�+٫2Îy��M�n��i�5��k �WH(�e3pv|*%m`�W��\����N�}����9�}�������5w&��?|L���\)���~�50�M|}(m��=�mǽ�w�4�}����b��/��+�n��k�.'U�:#�r|��QZ^���W�;���^�|3�$�
cd��+�â:�i;�(;ʯ%O}��s�#]X=��h�.�G9B`Nvlf��W]��S�2�̳1ʾ�aO���4��gZ Tg�[�N�F�8A�U�{��tw��?t3ؘ�3ڴ:����'2�d,4}A_�*�ė���
�<�wޔ�9�	�ߪ�ږ��!�u>rr�F.�Cj�w����_ѝ>����'����G]:�*=85��4bxt�S��Cՙ�W��7ŗ(<
Y:��/r-�6W���o��B���q�I�x3]}�v�9�T��׽í�wv<�}���K��k��t���Yx}�r��C�p��k�P�2�WJD踨��Y[ZUrbm�(�R��m��"�{F*@_A�?�7cj�Dyly\{���dQpْ�Yq��9�r�m�����3��t�U�I�8����wQoCZ3uu���b�U�U�j4���I���銆d�P�wI��-25d�ܾ�=�}Ĳ�p�b�*Upک�9�_U���������v�M\=�uR�xjշ��N5+S'�� p�_3��FXq"���z�b^µ��^d�;\����z���VG�d�6i��A��:��If�D@ި�0��I�<�{�jZ��-�`cx"��MfI����+�9Z��Cu�I��tF�:�&�L�5�R �:�+K��|��W�6��PK�^c�����1��iO��T9��nw�_����B�%
��R$L�;L�H��OV/ݹ?z���=�{�e�p��F�]nM�r��}g>'��"49�LR�sә�I�[��s�����gw��7XU�t�43֫�׾ޥ��:!��RcZN̛�����2�l���.����꼉��T��Ih��C��'�`���)xo�i��x�'w"��32�[��]t�f.�נ{=�ŷ� �l�z����su�:�7�+K�����~��a�����.���RwC]x^��{���ά7��_��T�\d�9Ñ����>6jV�.����v@�*��; T4��0k�����{9��8�dn�<r�H�z� 7B�	%�z�S�t+��s8\�&\�ϲ��$s����ܼ�q���팠j�ȹK
����+�$��W�����KՄ=��3��&e�LWpm�Vu����3;`�J]�l�C3��������d�'~j�֥�����
�ɿl�p�*Ϣ���r=�oveS����"N��_�'�{�T>�T�2ɖ|������k��g2|}l�.)Y�u����w��]��L��S�pY���}%�1[�J����g���3}�7x����X�vNwj����O[�.,�/A�~��Ē���j�+�f�X������t���oʘE�GS^��yF�<o���/�ީf��'h�&j�!qS=��6�B�n�.��b�)���Mvi�x����]a�n>�^R���Y��Ux�b$��R
G��Y񵃡�
/�	&ނw�v�8�y[��-N�����}De�'v���R ��(	��0y����e�S�O���(��V7��v��Ӿ��3�������<ݑ�iD��@{;n� �پ���YO���|��`���q����p�D*v��|�6�9gp�����êf@;яm{-Nx������2Z�#�t��<�h_ԧY�Ga_�z��K��<���C>d�Y��8ԙ�1L�)Ss��δۧ�o��ScO�$���TM�/zI��_*��4�7��fa��V��ܨp�sw����pS�]X��wi�j�r�M2Mۓh�{D��,L٣��_r�f>V�Ņ\�a��=�2kg��s��7��7q�F�J��~t���f��c�J�tn+һf��u �*!��[A��m�Dq���#�w�݋���h΁��n0
�?\�Q҉ڀd-!�ǢV�a�VO3��P�����/��߮�|x��{f_;;�\����n���f���Ѳ�ڀ|;H�c��f]s{�>���f�â*>'����1��R��$��9Iq�t���X���3��e�ƾ��c�}>뼱}Xaצ�sY[�>q�OIӺS+�}p�����=�N+YX��'���7��
<�x���~���^w��������ᓃ��N=(�{e �<���R��TS�G��X͇]�*>�hܽr�5��K�������N�Q9�¸?��6gǠҠz e +�_.{U�y�3&��_+����^����}f��u�4���s:h2wz���B�3�iH�ڠ�o���?��,VTz�E������È�µNR�8�w����Z��f;���O�2�;g�rs�i�=kz���/vk��Ƶw�U</Ie�}n��Lw�W���d�tt�}�x�ı�,\P��dvME�N�-���2��u|����s��q�{��;�5��ǔ׼�x���'��agY<�;TT�36	���a��9Ab�P:+U�g6P��ҡ]���^���]ux����(7.��G�!Bp�oq�k7���3:K�5��2���QsB������v���9�k�VT�����u��r�a�V� �s"��e-�A�+��r�͹s��=d�d
n|v%����9�N��)��(�!JRu�*�l�������}�	5�eg}�'B��G=;IPՂ�����0�w�K�kV:r��X)m��v(f��!4[�>"��N�3l�ؕ.��X�2�jEMe�)��:8�Wî�ǵ�z��6�յ���Y7d�z��V����"�=���@q��ZtA��	��$l�����Ӌd��S�;��]��Sȳ��ɱk~]m�.�}���4���Q���3�������];��P<���7{Z��(�ѡFQf�VPYx8~ܮӓB�]x��2����P���c6�5&8�U��<�	-�_vW�uf�Dϰ��YDe�zgV���1}�$����i_Á�o�j[|l�U�9���u0��9��3a%�t���:v�����٨Zy
<��f�����zrGl�wj	\y��᎒ܩH�� �Z��(H�6a�d*�\�o�]cX�����P����Mh��D�Q���x*�n��d|�S.<.]���?.oI8`J���w4�M6a�S��QѪd��n�Vg XV��v��>�d�Sa!Av[��Wʑ�s�����墑��9Z&�Yi=Z�g������:*�qT�������MI��T�M���A����"���p���5U�R�I�e�)�opf"����pKS\1!.7�p����ƺ�U�⌍�ȋ�f��z�VU��������p黨)n�|���bYa����:yY���lᙬ�"��\���@�3B<��ʖoQ�G�v�)������A��p+6<�8��Y�Q嘃?Uыfg_3��`��l��.��H
�C����]�I���"��W���#�B[�3���h����J�G��]��m�߭nT7��9��V�79m���]����kb�� :^�ǉ�ufʾ��\H�&�=����LUk��>!��c���o:�3!/�Ne���ש���ј�E�� e���fe=Ư�i��nck4��z�-����բrek�>P`HlNq�u�˘�4�.�3�iM�9ݔ!�r�R�v�{nln&d9�D��Y�Zo�i�e�,"���ܨ�󃁗�öo�V_P.���N��Vg�:|��پAG�v���Xg��ރl�ts�0��%�Α��ۂ��Z��&: U����Z:��t㍙�6���,<2���Z	s-�K��]�ݽm�&Z���}K�4�ᴟp���UX4�f�\�PJ�8\�R�v�Yˑf��I#�UR�J�i�21G.�2�Y�$r��,�p�B �J+�iU��E�!6�1"��eq4J�)P�VZ�R�:M4ƒU�h����t�+���͹���VZ�zSL��b��(�u����]�\D�l�G"9y9NLw˶UQvLp�/R*3��F�U�dQy9ܝ~��S��7�*(��"���_:� ��	��H��*�rO���v���9�nTr�����5;"��8U\�r�D�We�!ʉ��
H�>R��ϑ�m�y|O:���9�<t��;s��.��t�/�����o)�����ՔݔJ6,��v�O`��WR�x�;���w+�r�}��UpV��چ�[���k�4� �c�g��_��ے�tz����V��\B�oO�Iei��,����}י~��s�⣠�_�2��La�Ý�	���'��`�)�.��t���ҡ��=�����[:�u���Mgn��:�
,��������R� }7�eZ놎�[V���m�;�7J����K�cf}١�w�ӟ��W��*���d�Q�@J��13ζ��Eiy�5	-�#}���x2�qI�&�y��|�8R��LJnp��J%��=d������u�㴔Z�N�۪�W�{;�TM���F��u�6ۮ��`~�k ����Q:(̦F���>�v.�o�]V{M{֟UkB�mn����+M�.{p����~R�2o����P�.�NGL#��^��.�6�kɾ��9�z�5�>
�p���+ѻKM����ruXc��✛� ��7yg6c:��veϯ��'�������"�t=1�p2�)/�R�';��A�G������bt5��х5s�Y��9ی��m�f�ߒ�@��6FWz�b��?1(o���Fu�g�[�{���φ`�b�4yɬWm��{�O,-v�6PqWc�l��E�Ufh>���^C�7�c{��"��w-	ӵ�F�gv��3H�J�a�e�����h�v�Y����~�q����6����$P����t ���[y����Tp_T���ے����mm =y��p�ˣ���a��ok�|��7�Y*�T�"���d<4~T�ʭ7�2{'Q�͋,�/J��vҐv�!��nNE:�]-���m������*3f^z�.�PB��q\wk���2{;�x���	�A�P�atɴ��{��)�T{69琼�����t��ɱ���[�d�*��hl��T�)�����Z�r��Yx}�g��\>�G�W*l���,��k�i^q��A��rA�tqb⧫���O��W��<�:C=��;��#gE����1����W�Ë%��$�}P;�\����]D��V���¤� �&߫��6�'rq��[�u=q�\���?}�Y@@��0�L�I��߸�.(�ĳq��>Y�wN8���p�9�|w"�M��#\��d��� Jj �"e*�N�y4�dݏe�>�z���U٥�c�����I�G��sKg�`7��-ϙ�I({�R5�ˍ_3�]�E��s��d9�
���83Ѧy��o
��K�ɶ��,��2_���M"E��4��]�������qH��1�@�n^
ݳϲ�3�}k$

Wu%Ɓ�&�2���E�{�;�G�Eҭ*�!sBwgpChc��k6���I$p�˳�'u�w�˄�]�Gp�@j<�o��ݔ N��3:�_���A%�g���o�c,�:���bk�CqN��OH&91��Q*uz�v���-6���O����Iٓiˁ��Y����G}��|sʗ]Ӊ�Ӗd���'c����vW�V*zo�����z#���Yx�Iz�<x_/f���2�g@;q{��yRl�z���	�1�N��\�/������PR�=���W�W���p�R�_�Ϧ��O&�̩�҉����̨W�|}��%�魎`ݽ��[������#�o+i��Ա��CWQ�k�jY�,X�g�3��^޽�*{����ޗٞ�hS���M��|O���s�A�Q=��ބ������7}�q �%��ߺJ�����O���	�:��tp\tH���iW2��S��y_\f��r��YGλ7�۬]t��7�7x��P�@3���_�T^��C���Hq�!��Y�5i������3ޜ���m�և���2�������&A�C�3�n6�]Os '�Ys���"�6�V�ק��<�y��ӷq�/)CK:�U!���{�Ցy��8��n�@�ʵT������[�Ҏ� v�}қ|�p>wo���1����,�%�,r��ɋ`�/līA�� 9�E���g���;�˦!��yCZ���x�P?&)�ճ�:�c�o$�g����k@�{��C�k���?�ƍ|�959�8�/�WKV������!a�>�2�N��|J�R ޒr�Ԯ:T�|�_��T�@�V��U��Э��_Ν�O��-����ni�2
5�{��W.�[q�+�{�1&�L�{2�0</c��7�ޮ�N�1�s�ms;��6�']�3��ڲ��{�n��ά��O��RBv6��<�h])�s�e�p����K��=���q�3���/�i�r�n��s���mG�S����2���	��bw�+�[N�ץv��z�v�Yt.��S�n/mD��������N����#q�'u ��� �Zl�TT������v���PjdX��v��//ػu��|�mCj�MǓ��L/���� �d�@>��O�o��jb��2�s�u�}�֑{s�{�Gt�7����$��F'@97�t��yt68�L�K�s��d�w�{8q�y���]�r�9cn+Ԇ_�t��;�2��}p�����=ӊ�V|��'����#A�<<"e~�~�"��z�VU�5o��֙��Ó�(8Á��>���u2s�Ԁ���C�T��9N�um[u����*�&�f�l��v����H�f!�c����-�/D�g�Y�m�x��K0P�]�DdR}t�t.N���9�&m�M�	�>!m�,Z�{KL鲝6W�|��HN�;\J���&�-��OV�u�<�8�k��(%F����56���9�+��]�(�Kq�\9�az��(]zk��@>��@Wb�];*Z�yಎc���o���i�Χ����г�S��'�L��3�
\���� �H~�0�:����o�vyС�Ǻȸ{<��[��;�w�z�_˽R6��t�}'�����c¸Bه�x����aq
� Oz��xk����K/=�ۄ�}�1ޅ^�����:	:q��k���`Tթ����x����S=���w���V��.T�%����g|��g^eկw,�L:���\��ǔ�kx�������@���3�n�S�\<5-v���8z�5�)DK�)�N������pm»�0��x�Az����H�M�q�:�����-�C���}ݢ���j�+5�~�uv�p��N�t�&���q����:�7Eiy��P�ÿ1�EJ��^/�^�g,�dpq����9uĶ�'a7Z�Q9
e���&��B���1w{�-�1%��N��?���m�˩���p/�� k�#XB�@�t�tS9��<��"<j�1�֖R��k���<�C��7idhk��i��UٜVhc>]yl��Ԋ`"��;un�O�ވg ۊ��F_q}.	Kq�»u�X����r�N�Dۦ�o%�f� ��B	j�����+5+�ʀ��4�L[`���һxmYdS#�iX��}3�Տ��չ��Q�/J����ܛ�)L�6۠5������x0������N1�h��q���:i������[�b����B�˅�N�Lbq.J�� ��[���>�{�����ϋ�g��OG�>�O�ةxp\u��wѻH;���a)yq,v�dj�f�#��R���};l,�8}V_�vlג�@��42���{~b��>>���#�`��o�������/�J����:�V �\okiE�eLe�K'v�����PwYU��AOR}�o]^��[������ TG�� �nJ�u�}���ko��t�N��'���B8�uax����U����<�mR7�\����.��M���/r��e:�g?_i�8e�aL��	�Y�%i�L�u&x+���JD�X�(��K/ų�ꮨ[K'�Nڶ1��U�d��͕���(�e��7��v��$�������u<n:��U�ݱ���:C"�{�3�b�q��^ճf���=�^f���I�P;I\����]D��k�(.��]�g���[�����+ڋ���u\���x\Ӻ��R�}�c7v3a(C�.m���ߞ��tc&:��e`��I0�o'���)��Y₋euo�\�X������b�}���á�Pv�S5?�de���ᰁػe1�a![3W1�d���˪���aǁ��G�Q����p8n�p�=%��a@ҕi6O3���un���'j*�r}���3��b�qW���z�>;��p�o��n�	�2T�q %5��LסwU?d��:��=�}�j[£m'iO��T9��nw�3l�$�+}��xd��%y�X�x��I;��\T�83A�z���.�%���Y>D��U�V�&}s:�w����O��o[�$8W>�6fc���
�s�и���5��Zn:!�'�rb�N̟7���dU]����-�g=�y���Ȩr��5œ��L-��/�*We��b��������@W�k)Ep{��Bu��9m3m� �;�� �l�z��酶'0�]:�7�+K���u�2_�R�5uc���ח�����6?��W{�h\�\N0lw�9�	G�cO���u��:���ϴ�S�N}�Z7�=*��-K�_T��{��/O���e��2&�SO��sW�r�c<B:1�z���q<}��P*=Ϯ�β��R��&�3y��3�uo�k%y��U�s�༩pή6`RP�@�{}�KH��O��$�S�%�3��-B[�N��ٗL	W3\-��N��@Vbr@�X]i�x6�!�vv�wֈ���w�`x˅R��ӻ�,�3�G6Z�;�fU��^F �P�H.0��NM��d^�»fh6����gG� L�r\���0�;�+`��W2��)�]w�T�������u,Y�w�w����N����2��҅�T��{j�+��qʐ T�<�޵5�k���޿`�эu4{���)�q��w�Q�:�	�A��.�{���t�.�}������4��vav"��z%��d��������E�#����1�}P�zoH49�ٽ�io��]a��w���ۊ�����5%��|��Z|�H��vÁd�@ҽ.~���SP�����ՀG)�X=ǯ��>2�a�}�Цq�ӟ7'\y�#.�3����GҼ揳��}8Կ%d�Q��A�S<=���kz�w�S��z��E��{�ls讨��<�yzu7��=\��H�Z�άD]R;⃨��GB�ٶF\wu��p��X�Vc��9�^-�r��6~�s�JH�:ARv��s��;����J�ޔ�F�(j�7���ՙl�3z�E�ҦK`�1�Q������Q; �����k��QLU�uJw�>_���>�^�~u�m�MT���Tѩ/7�[)d��c�F�H8'gn��q°d�Z�/U�K��`oٕz���O�����i����g�R��������}��P����i=���@��X��l�䅕A,���z��u��ݯ�n���}�{zq����p��Ϟ�	��6����v������s ��N���Tݼ�-���ƨ�Y�۸=��.ſ��a�˝Ҹ�Gt�7����y'w�����������f�(�3�E��K��_1�YK*x;8�W���ZN�F�n=��Ҧ��N+YO��v�z<�O��l����x���N������rr�eC'���Q�pk��9��@W��ކ=*������z-��zP�w��֬��V3}�8�]�������0��C+�Xn*��e #&����G���ԇW~5^\�m�!�=���w�]p�>�����4=�2����^;�w�wL�����w�kk��X�PA�0�d\-�nw"�0ס��c�����]ꑴt��"O3�K^.�cmz4R�+j�P����q���;QkU�/@�O��^=�OeC�Lw����Y+��=0e�[�'�/���q2����P�*e�c�޺�n!Z�k��>}%���d��}p�,�'��vy���宝�y���(�8 k�c�����wI�NxWC�|0y-v���L��LyT!�f
7Y�CD{��s�J�q͵�����ǀYx�ºi��t�K�Q�魼ȧu��� �Ȉb����/�w�Z�@��.6�̹)vC��.��J���pw\v�զ�T���j�!������}�n�Gohb=��sKTW�y�.38�r9I��7�.���m�^��}�@ޣ 9�R�"����}�P�Z�����>F�G�ǌ5�&�vx��jsm�n�I�7ptۧQ4��k���&.'�m�+K�l����U�n�ۓ��r2��w8�z���p�V����_���ɿ�u�[�q5
e���!#gd������9<�i�T���T�T^ܭ;^����Lf�˭ɶ�p-�`hO�_+�N�{=r���V�ry��ޜ~�ʟ
���W�Gh���ZW<�i�T��)�&�@k�T2����/;�Qѷ�Vzd���4}:6�t�+��8.2����Zn^\.N�v'��gF *I�u{�,�u�ݳ�`�W���f�'X���X�R���U��iqۼO��Iw4!9B�L�_:��/���8p��j��h緂ůz���̳1΄�W�zD��}���U&z:��ܙܽ]8� �s�=�ރ�j��.��,�s*c/�Y;�����Pt�ģ�>�Ƅ�Tv���}���S�K�����yε%�:�]-������rwb���W��V0ǝ�A,�i��Oo+e5Xb�������ڼ�m��D�8\Fu6��_wY+MB�ʺα�x,xz��y�C��*jc��r��;����.�3���}����E@������Y���ut����eT���ub��ʾ����f�t�E{���<���.1Q�6r�z�-�y�F�VWZ��u�x��R��ʹZ�T'J͈n��4,Nw{B8s[1�pI2�r�_Lu�x�N�F�����e7Ҋ�옕`{�Cwf�&J+.�%4�C�����:�����'�vu�S�o��EG��M���Le�/cSd|��v���X�����P/�	�b��o���wZ�q�;�5���2��|�6��Egk�&��^�Jθ-�ܷ*?��}\9�N�>�����j�(�x�VN���u����+�ٙ�k���&�n�M>�k2m��.�O-��n��ߢ�O�t >�.��R��3b������p�ڝ�&�9��U"�+��eAC/�,�K4���#����GdZ��i!oM�m���8oFݶ���-�ĦKn�:�ͥ���l��¯@�:1Ҟ���q'N��u�i�+[1��{`�7�L0;�EӦz�� �����t�u.�z��*�
u<^��r�:#�κ҂��W/x�8	�63�"޷���1//�b��{#��j|�R/k�(�Y���ȉ���Ϳd��@z{�d�^���T�缜�p"��4�ش�=�TW�7�a���we�f���կ����)�Re��QԾ�97�����z��B��#])����Jߝ��PE���f�H�78-$oM�i)oa�j�b�4QZ[��1ua�MW�յ ���n���YD�)#��@lRЈY�b���n���`�F9��A^h-+r��51ٷ�yS6�N��G(��j��c]�v[�:gv`U�}ѦX�y��2WfJ<ta��]X3FzC�`��Lg1Me��__�ֺ�d�&�U$n�id�ϠN�8��A�IB��;�HmsyWr��/�@*�8s�P����vm��́9u⳹�x�v�,U�x�\ʨ79�2uW8(C��7�Z�#� }j�T�je-��]y��qۈ}ڬ�7y�pW �;�͉�|���u-�פWM��bx{C��Ӱ�����ܻ.���'hEt�a��u}
�S���}�uJ�+f��v�CO�޴�̃�ۮR��޻�N����f't�|ҮN��BZ�RA����-nf�nU���W�ɩ�nB���������L(�����mG��Bdͷ}���J�k�yX�f-�.�s��:9Z���o�wbי�c��j�dՔ�6�}��q)�8���2�2���qr��{F���t�2�k�-�o(�82�����S�͠-q��a���{x����'���)�T�ɪ��<�|^�i2��HQ�t�4�GS��m�X�ǻ��nf�
������*�igW`�^���
1�����G��UI��Z��Syݲu;
=��|C��F�<�{��ī���ʫ��Z�r��ǎzY'�	U]�(����� �<W����G$����.�Ng��.<yʹ(�DE˲�U_�y�G�r��g��U��ܒdEP�-��u�r.�ú�+̊��� ǈNU=�)��\�5�U�z����9G/uɗ.\I�,�
���Ȋ.���Nq"���p�|�+�q<� ��$�Dr��"��yҧ:�$�2�EM�GX�E<�T�lXTPQUʞV\��*�Wg��u�s�̈�*�=Μt�$�|���IHC^-p��*���T����iQ�Zr�uG32�$�*��`Y��UE�>yǞP+����tB�T\�xw�/[�; ��uUUD%w����Ԩ��=hr�B/	U��E$���9��$�p���>'��
��	REʫ�e<HQ��7D9Tz;���4;�β�"yK���T�
�0Y��O��g����`Y�{��r���f(�^�xdp�"9��;̇p�MR��۩�}\6����l�ރ9tH�^v3��(�?�xP�mCQYT������ˀ����p��/i�6yC����s� Ҏ��u{kkV_��}���l;rIʙ��&t;��}1{j���Z�r��Qe��r��*��bf.S쫬�z�|%�_��6̢��H:
�|P���wS�㯪�\svƏw�-Fs;�f�ju�gU`ǃ��;p��{��Ë%�t��e �+��.���� �s�۠��վ´Pz���ki������
t�@��P7��(*�i�r�>7�]�yY�Ԧ�sF����_\Uç���S���|�p�n<���	�S%Mq %=���|*y�ǎ�W'!R�{i��:�7�=���5���q	;H����9>bw�3l�Ez����e���3��U<&CU<���&%:�W+N���mo
���ܖ��Yd����ذ����Xs�]�t�3Ć�vvl��V:�
:��=���ޥ��:!�}w&7��Z��~��=���Л�yb읬fK[;{�Q�[.̓\Q;C�`�1��x'�7�(eo?���ѻ�F��oR�I��&��{�� K��^ܸ��ea�Di�Ǚk��Cf9���frv���N�{�;�Z�QO�EH{R�Sd	�cv�t2������4�ʿ�@�YB���F�uw[bZ�qk�)rh�p}�y^T�X��(�����w"��3m� ��?`�z������j�]���nM�z����#��۝�~Ӝ�p�y^�BUOO���2�_��޴�Vݴ.b�q�����g�k�_�^��ϻ+xV8�S�"J�>.3�3q�=*��>���jr��羽
�ɷ�nn�葵'��/3��1�9Šp�^5'O�p���'��P3���(�2�_S�G�U���[*3�μ��Q�����(]��?���	b��%���J����X�l���`�wS1�=���?*����� ��a�{�~~|�t��e��
�t�qS/��ڠ���d䲕M]�(}u�F��{K�CZ6��7I����>���ީF�Βv��{���SK��X��.N��={�w�;7����
��Gyz�?@����l��n��|���x\�j!$��XE���b�����r+>�(����]�f�V��%+x}Ijw�h������N��|J:1tk�g�C�K.� ����be `${�4����[�}�Цq�ӟCrp�Ǜ�3��������U�n��՗�vfh];�}�.�fRDt Ho��+���y�_�:c��ǝ��Eτ���{L��t���Ku�����z�9)�� .����Y���6 ��*t1����r�V3�F ��[���9��|��r��u��܉�gi�~�2���pB*�@?$�A�3���+�����z;Hǜ��G�)�pez=֞��n�4����A�ꑑP�J5�$%ch��Ϧ��)�s�e�p���������ܫ1��D�g.���a�Y�~����>��+Ν	P\���;d/g���~�Y�|���7���:�'&�^cY�G�ں�B��)d�
F� �O� �J'j���~����H���O/t���uֵ�tʎ��=�=�j�O���v����45��>�e��'���p�`f^�Of��3K���]mf���+�wJ�}�^I���'@97�t��=������pS����kG{��gZ�4},u�����uJ�p����\?D���<ӊ�T��s�x���{�>{��q���׌�~>F|n8�98K�Nu>���5�����Ԁ��>�1Y!�+��~���X�c�?
��V?��{�X�^�S���s.��	|P��Ma���˦/HS�.������Wm9��`��'���R�G�
�i�y\/;�:n�'����@�O}���[�R�Q��Go`k�(P�wV�G��y���5�fգ�Ds�-�~�Y���������V��[aA�%�����i�i�ǻ�ٹ�
b���w����@u���м]@�W�YP�
�C�W�J���u�4Y"�4�Q�z�v�vF���{{D�wn>��y@s��j��[�-l�s���a�U���^��R6�t����ೊz�����ԕ޾�kK�;Q�:���@�o���k����K/<��>�D;T�u�f`S�<�y�v��p�^��I��g@��uC��JX�z�Q�V��\.V��%��=���p��1)��ͩ�ᱽ�<��r����|4���Pex�{���t�t�9u��O�z+K��Ld��d�gk���p����[��a{��(�Ax���O>�p(v��K��Ն� 1�;��wK���wZs�ln7]���n��t�&�(�G*����s�Ūf���ד���/[�gVi8F�'�d`Ԛ�=�����d�n�v�%�{>BF���#��I���`�cq�,�>u�7�+�׻�7�������n� ��k �WH���F��jݍ������K������>8�:[��x�7[��g˞�4�T���S&M�n���"yLLH�Jr�k��.���O�}2i�q��Co����T���دF�-7��˅�N�Lᝰ�˽6{/��o��{w�l�퇨 �k��v6�~cz��� ��L]��� ��ڽۊ�ʪE�m���k��V����r|Mó��Km�H�e�l��R<J)V*����S}�ی(��Zؠ4'D����t������R��d3x�j޵�~8?zN�;q^Y�/�ޖOTL.��Vu/�:Nln��d�^�u����ys�[CC�����N��Y���z�{x,\$�4ǀl�2���6+Ƶo� �ّ��uq}��ѕ{��~���U�_m �%W��p|�YY��x���neLe����pf���˲UT�����~y{��qN��M�����R T{�Yι�9�1t�U�������:a�y^d_�v���3�D�DݖeT+�U����h��
��JG�x�-�6S���`.,�+����Y�s=�z��7>���d����&t)%��m��ֺ��]0m�^u�/D���]�s5����y{p��k�m�^2j �+�*�	�\�J��ϓ�B��s;]�q�t/z��w.�/F�R�{E�����^f���P��z��$�E|\��}K���������mNױ�w8�z��Pn��ki������θ6�����,�B"�A�P�6��*�~\3=���\K%a�z�\n���t��=
r��놓qn��2��*VR$v��}�����o�L�0���z��v��{56,���"�/3+��U��唖��
@���]�< :��k9փݱj��x�rc}���On�=c��D�0e��th����U���;�((��)���u��=!���aǰ�.}�q"�n�1��uwMy=ŀ2��zH�ܤ���{�B�kxTm��#�3�[9��X(�p4��.5�[�vh��Ve��pWΥ24��n�Uԭ83Ѧy��[£n�ro���,���g�]#˯k#��ٗ:M���T9�$TG\�ٿ���;���Q�hg��i�F�-+����Q/�}U+�Yw9]蛜k���L8X�̖ˁ��
�"�eْh"�ꌐ���^���3ծ��r�w�#�wݵ蕷���<һ��n�G}��9�nXo�~�b�ו ��'���[p'0�-s��4cb��=��z�S�&�g���۝�ݝ�Ƌ��[����}��fn�8��2��r�q9o?R�c�y��۠���-���Q�^��IxO���W����D�����5�Ʈ�z������p{=Wѯ}ގ['\9`���e�����+�Xn	�O��P*=�\?DJ��Y9��-ꉅw���^��{˼1��l��a�Kx�7�x[	h��_��>����9(��+`�ҵT)��Q���K%w����G�O�3}�w���gz�M�e��peP3�	%�͵A�6�,!�[y�T�"���e�(��=��.��&�m�m��X�W�"U�w!3z����b�7z�����yF�����gK%�{��յ3-ΰ�
��-|9s�SOV�ӑ��1��#�P�j��MY�n��z��v��l��4����@\�o���Wݽb�({�:L���p|��؅ީF�Βv��f�3ԇg����{�1Ͻ�]���wX+���!xkw��D�s�C�!������W���(�:I��g�X�����'��5Vw����Xe"��	gU��������Iju쐰��Q'vè�n]D�(˫z=��z}+z_�� �ĞG:`�)��*���o�)ˮ�Цq���>;��j�wq�ms��W�G��e�mMa��̃ƺ��2iV��*3���T�`u��Gكl����uI��;�槫�Z��&�wm�3"�L�j:����'�M	GY��(��k��K0w�^���}��)����_Yd3�J���)R���*Nؙ�w&![���D��R,�5�j#3�/c8[u�\>VC�]ȶ�2_���#q�'u �D��yN{bv@>5�&�X�P|��.+'���v��\�O����� �۶���wR���%����Z^^�C�|{:Y'������'î)�a�/��P	K�`g^�x�����M����������o��c_��G��3���s��9y�y�詒]�ڙh:����ޚAX��6�[3n�Ү�찫���3�tZ���Bc�vc���u����ϟ
ٓ&�[�Cqu�ѓF���.�T��W��ڡ�F�_VR��+��w
wZ�����z(��<b4�7�{������}3�X<E�6<|��1��t��=��_��X��?a�{K��w��{޹�o����k�ت�u�ךm�"�������_��X=�pB��	ˬ�����Ƭ\V�wNk�ݾ�Q�쭴��{�?��{>W���S��d��2P���׈c��'{��^Z�|S�w$)��|��V��ԫ��S��[��Y�rD~��2���$W�<��>����N)��#u� ׆��0�d\-�nw"�0ס��c�
�|-w�F���uq����W�����D�E��P��#nT	Ej���]<>{%����	��R��o7���siǦ����n�p�Utt��]P������u(ڵV*���ޟ>��ӑj���v,��y��.ڶl��T,^e��( oTA����k�{���wI�NxV��{75.lRu�T����`qw�q|O���n��û�axzJ5�2�-�,�}>q��7j��&�(�ý��=�mp��5h3�3���o��6��MD#%�� %_	�c�D?�y��P=��s� ]��/�F��0�]��� �pGZʙ�~�̋@m#e�f��\ԝه��=���:��c� ����:˰�i��=k�`՜�:��RE_C��t�E��u589~�-=%���FWEk��=����9��G44oz��t�kRW�ʷ3�������+On{�A�|��E�ڴ=]q/��M��@�v�&�˙���ݚF��Z���{���T�3�J�Qcӛ�	�И�����lJ bp�`�8;pr׵��t��;cz��<l��di���`���3�}���6���]2�G��L���������B�wdm�b�v���2<ܯL���g�x��σ������[LWF�-+������vc'��WT�K���0�bT��.ۆ�,�ixg���z<av�
��xp_Z�'Nm��Z�H��	�r}Z��޼�;���)�����5O}��k������C!zڳ���
��ꂼ5�ߵ��f�N�F�N+����D��8�| ����c�*��?9�y��x�kiE���1��N�o�����*����ܯ`OZ�px��F�W���/��HQ�]d\�nNS����mV��5�����a-���X��ϴw��I~�uI`UGy�7�VE�<&P��.�6���A����w�,���Oz��_Oxc�{޾:}'Ei$�D�BgB����j��Z�`�3�`؂/���h�z�߂�ov̴ �Կ�l�I�'3�71�c�xZ�Y�W���S�?/\y��q/�t�y��Os��/�=}k�u��5,!e�`�I8�0>pŤ����P�hDS�Sv��� J"y�^*,�e�q�sD�_U��Y��{ݹl�wRo'�1���~G����f��#�2���k�(	��	=<6�g�0�;�ßu�}y�s
�W�Z07���{E���5p��Uy�qd���'��~����u�+1��{-g{]]˅먝�v�����;�膶�=�>�����N�BIf�zz/Z��j�}�1��k���u�n ����a���t����9�7\4��7DmêBe��h�L��ʪ�|��^Շ�9�/˄@�I��0�z&���v���-�s����h��� ���r��⼏M���#5d�:O�r�)�
��V���<��F���o5f�H]5GnNyg���q6_�g4��u�WЦ�#��Յ*��s�ꗖ�,J����{��n��{��Vj%�7;�k2��z�L4�=�?���C���O�d��z�d���d`����U�v���%�����Μ��m�u�o��x�rwr/��s-�͎~�c_�l:����B�+�0���,M���&�.���-�:�7�+K��4_����%T��=���J���}��۶��U-��Z?:"��+X�l���T�� ?@�avV��f�>�c��'gu[�'�gG�t��r".҃��^�iǟK�L��u�����\; �i����<���\����7No�e'�b�r���1��nCce�3o
�.	ҙ*dt��n2nZJ��ΰ�*�z|�G�#;�<�z�򲕃z�J���>'/8��"s�����6j1}���4e�!`rʳ�8<�.Һ�s)�:��F�A�y���S2���.�#Uck��1�ruh�g�"���ޥ���$u��"�Z��际n�q =�}�5-#	.�;o�7�?�fkڮu�(��*����k���v�̢m�L�5�
��;[˴���ٵ��1��Q���3ݚ�DX�\�l�\�f�Y� higZ�6w|D�ք@�O�2�P䦖0`����EmXJ'�`%]wñ����{q���\5+�hԍ�V��R�"3�T����us������=t�}�?X��:5���-.�������O�m�h ����Ŧ�h#��G����&rcs����7~�x�h���0�CYLQ��Ie in F�#�q%��U�	�m���Yf��-�˜�S��Gz�	P��]t�S��NE�48�.rSug�B�I�����D+\�r7�����}��k/3)����\�
q�[�{�/nr����QU��.��#���ԗ��<Ғ�"����u�YyT]�5t�*�0�.��Բ�+�Vh��؏b2������=Ն��F|-�y�g���.����w�SV�>�n���)&�����щ�-i����Y��S/@��͖U�����>���ZXnQ����;���.��dIZ-.���c���]8�eۭf�oj2lpo��� um,��q^�� 8ZS��D�\�А�xs��о�p֫e�X��m���w|�]Q�upp��x�V������$ݞ��v�w��Oh�N�ֻ)hR��]n��]�3t�\�=�j���{n�m4^!�7x1�;�Š.W;���u�����6�cS i�Y%���a
;z:��ms��f������4fܔ����ާ�nD.���T�ptؼ�x �h����]&�\"�kf��K_6�X�����TܺΫ:u���1�}���F���ݜ�F���ku��l��J��[� W�� w�*tP���-���C���aM�'!r!cksk;��f`0�\�+��.��<��}����ߞ*k��QD������E9Y��Cһs���nҏ��ք���ʆKU�����2��f�[7jS�w��T�`�U�����յ*$�Է�8f���y	+�t��gLRD�
.�Se,���3��+6X#�j�ܧ[���§mv*��o,K*�HcVG+z�l*;"=(�K D�d�gDg��t4s�*%#��:��XygT�\s�Pm�wf��FL$�*�$�5q��nY���gW_-�;{���Wj78��7��>
��v�m��Ryzu�sn�)�9�q�C֑E�0�$ʉyc�ā^eUn��Ε�HR� �w)Ը9� �*�FV�Yvh�m2V����&vJ$PQȹ�D&Q �l�H�X�H\��PT��q瑔�Ҧ�*�ʥ�kp��w
�&���Q:'	6^���nI	�YEsև>\�as2�������UMD��U(-P���˗E�\*#3�]�)tp�(��"9P|�DȮDF�=z��9��\�:W9\�Y���
����Rek�<�y�Ȩ���er/��ם*L�E_D��$Qz�&�{�s� ���AAr�$��E\��<���+�A�W"��yJ�����S;8RH<dQGUʊ��(��PW(�
��Ȭ����;�vUQA!P�W� 71X��/Wwpȋr�ww j�2چmj�]*�f�i��W3��ۀ�l�d���|�Ѣ�!L�c��N	�'�v6�Z�vz)�� _\���+��.6jV�ѝ)���[L��S��Ώ�Е����krh|'$��	ai]�x��|t�˜
��ZD�d�Ӓ�W����J��Y>��s���~���v�%f�>��j�ǰ��8/�rp�̡�'Gz*]T�ӧ%� ���o�PY��5�}{oAki�`˔��ڏcU�c�s8h"w\A�=@Δ/�|Z�9=l�R{��˽yu��{u�8Ú�������'I�����
k�aụ�Y�N��϶E`�W���{G_nw�����q�w\)�����5��臢[9致C���MΎQ�����E��%�Cks+��$���(|��l�]TK;�q��-�⇴B�y��5�\���G�{��M{����L��5�D�%,|
G�&��Э��[�}��g�9#�b]�.��Ƿu�|i��VF[�fj�(�ǉU�����q���ʔ%��2�&+�_ےn�Kp���Wqngp��7pv�uL�D�}�$%ch�9�Дu�T��2K�A�Y��ڇ����~�q9��Ѯ��֜FҾ�!܂��t�p
�]�Y�m�' 2}���2��g9����Zo�cQfʝ���1
��9:��+mC`���|��T��{[��2-[��r�l�6wE���Tμ�`��$���ޣ�t�ഛ��e���"�b�#n�a9}e�ϙ+���**��T��3��JP���v�nr>�V��֨����7�Tø|���t�S��`k�7B~��Q;��Ǎ��\�ܿN�\������ED��a�d�;~�v�i�\���j�MǓ��L.��^�Fm��MT�����Z�'�Gq��C�S��{r��������\$�V' )7y�b29M���Օݗ��vމ�̺~���l�x�Kp2p)��쎺ZN�}�����\9� .���:�l��eOu}X^��Ej+]���ךo�|���Grr�e��2p+��Q�f����əRR1"�����Ӯ@q���D�O�s�u9��>��w3�8�s.��	|P�W�d�Iw����wm���ר~���Wc�_�ڭ*y�u�4�����7Y=��fH�o��U?n�WK1.�6~�C�յH��}@52][��nqE�a�C���yW���w\�����{�w,���N��C�2��QX���t���Yx��=�����M�9�V�'��q����.2��@�{�u"�
�3�m��*�h�"݃���eetr�j�K�Z���P
�LNn�J�y@Q9���,-�4z��R���0�m�Υ۩�05��voAdRSr���%�F�W�m��E�6yY��1�k �::�D�T����d#��V@�`�q2����_�2���S(�V*�r����s ;=8����&��ǵV3��_�d����C�e��QP���Pe0:x�{���wI�^�=7�7Y/^P�^un����z��`�5��}'_��9n�хJ9�@�p
[$Q<-�lvg�Y��Ǟ��.j��3í�<�C�9Ͷ7"��n<���C�Q5�F�F7o(�᝷���T6,���T��Ƀ�n���i��G�����p�V��ˮ%���ɸ��h���M_��L38eټ�R�</��3�	�����{J���*�v㙸\�F�r�rm�\bX�$�eU�;~��/�K���3����:-D��pVG�����ޕ��sۆ����y3T3� 2M
�	O�ػ']�2\-�{��������P�|��Ki���ZC�qY2�@�w[F�_����ſ�+�1�Ĺ+�\����l�id�L.���\T�86�Z�����N�M���OI�Bq��ǒ���bt5��u`����X���S�qY;��!}u��TbDDӨ�eA�$�.ov�NX���/Vk�i�w�=�q�����m�*��΢�x�h��i�����ٷ�T�iad��͋��{���`�l��dIL�y����'��f�X�ve�Q�.�o+���a��;[S����՚D��}� ��>�=�ނ��[43KkiE�̩���"ğ�W��תs�D�83Ơ�W^��pjS'�% 6=ˬ��u��ϩ�b�MN݁���3@���~3����mϤ���<2�e��ڎ��u\o�P>���+�.�6��/s���_4��Y�Nj��~���4��^r�tJ����.��z4�r���//k���*����/��/
�˯K�Z�:V7)��C�p�Ц����F�d����DT�p�U��T$�W�k��k��p���pڶ4y�t�y�v�W|Uy�~��(�#���(E��F	���=�de������͟C��J�k�()N�5���>���\N���Ielw��o/:�x5`���	�c�I̤M�)���B�-}qN__S���|�p�o��F>v��T��Z�3��ԝ���>B\9��` ��RD�)V�iw�aiQxTm������il��7Z3�ʷ����Exد@fќ�2JR��;$�z�i���<����/x����+@�UXϻt��ΐ��d:ۣ��n�Y���=i@��&���-J%\�󱑡�����{EN(�4_��T~��*xbǗ��5O������A��k��B�Cwv�xp�M�6�G���v��
��B�3��δ�%÷��=6���ul�'c*�&�w��/$����}��K�U�#(��S���6
:��[��J^4z�Hy���zeOfwf��j�![}w&-��ɴ���ȯ�]�&��v���vaM)sG�m���Ww]o$��]��e���x�ܝ܋��tͷ,���,\kʐj6Y=�s1�9�r�-���Kf�]Y����Z_gu�����[J���bt��:�p�,��ޙ�3��+�]{�;�F���r��L��2�ϥ��5+	���L����c�*��>���jn�1�
�;X���}k'�����=�,X��3C�`���W���<��rT
�=Ϯ�j��w�K��G}�/�t��V�q��FoCW�ea�K����|%��tk�8!~c�,ث�ک)�c
z���n@���j����&{Ժ�7�ޣ�w�t�Yd�X2�(A�.5<���0e�?N���yC���f�G��F�`T�y:L����S^���(��N�Q�&�����Ӷ;h�z�k�����on�?B���^���C�-���!�h=>U���ߴlW����Y7���f��ߣ�@�70/`W�h�m=��j������* h�n,{ӓ����ҥ�;�s���R�f�LN�g��L
�톻��R�g��7{j�����";5�K;�T4���yx+��K����������&$�ɺ�͓{�x���J:����)몉gU����?jKS�������SQȫ1�ͳgJ�
n2<�[w�� �HzH@\@J�7 �z㲬.>�o�*�Ӿ�ׯϮT��ٳR:o��9��>��]'\y�#.�2�tǪ&@iN��S<=�!�z㞉dgӁ�	y�;r^�q]|�z��G>�3�M���;n��
d�Q�$%p6���Ϧ�yVL��m��.���%��Ftu�������a_Qd3�J�G�0EN��2����_%����m��de���u�'e��+�o�ԃ|��9>��pҦK���_���)?\���"p���Z�xM�5��}�/I� ��7��TT��a�d�;{�.{l&���r��v����4��/_c���]wO��mԃP哴��0��s���Z_	K�YA��V��:r>������5/3ٯgm�r\-��:�]�/&}{,4},u��
�LgT�'aL�B<ؚr��M�׫ͯm�s�[�q8�'�q=p��4���U����K��1��5l���v׳�C��J���F7�����7���t��w"�	8m��g�}��\i�9�f�n�;���rv�m�l�9Ӌw�vm�M�Or6�B�i�n>��������2IVjY�H�h��5�nw|�p���<��g7���A ZCc<��,௻1__�JnTG�q�{�T��9�:�y9��{^��{�8o�'2����z�g�Z��啼a��kM���]�R��_j���;�:=�|�W��T��W� N��1O/	}��'-�f=�_ꎕ3�#mP	F̆an�Zy���[��;�s�<���=��r����+���I:jJF��B��/��ʁ(��U�/t���Yy~��c�Ug�g3�g�;�.2���DK��^Ī�S����!��ة���}޺�o�j�T��(���B_tT�1�z�j���/p�]'����gn<��o��2��>�Az��$t�4q�;��TiWBn��'ν������R:w��-v��Ϥ��7pr�ݣ��Q����/�ʃ^�V=P�깳�������t�Hq�����:�Z�C��C��c[��z<�����N|��S��+ؙʏcwoXݬ��(@˃�Ý�Tn(�+=ơ+[�#E�MZ�ˮ%���ɸMց�Ƿ�9d����������Ϧ]�29�;$L��F��+NU���3p�
���u�6ۮ�ܢ�:1�zn&kcd�0=T�=��y�qX��G1��0D�V7�Yr1ħ}2*柗��8s��3f��*�^�8u�{���%�1��GqC�^	y/4�X-��s6܃+���}Yڧ�V�o�V��Y�݊%��'S��a� >[OMMk$��oq%������.�fe^�����@V/ �WQ���PfS6v|*V�
�]s;G�Ҵ�.{p��t��Hbn��7~�����VI,��ɸ����U��_�MDt�=#������=���b�l/s��@�L�=^��c���+˄Ӫ���9>e�8�z���ώ�Oh�������c[������S'��T�����(el�8�v�Wۼy*{���c�Q����C>^�O��Nd�y�M�g�}�p�>��_���]���J��gZ Tg�[�N�CU���]V3O�ep��W���޿m�ey�v���r5�Y9��~#�a���7�2z2P�m��srr)�b��Wۮ)ڬ��׽�䧖w�4/�ܶ/��������^4gj:�W��4zˀ���_�u�{�/�[[m��ܟ�c��0�E{�}q��y�/����{$�'��t-���U>���˺�߫�\4��$�ݘ]F��.Qe��7)������|�����F�d���,��w�F�Ve�Ƿ��;wV���t�C�V*���|!�d����{肫�Ë%0����?8�V{E�O'�A4�C[y�+���e˘5�CSJ��������+��SX�|Zuϫ��wMb�ȷ��җ�4敾�-G�$�`�S+i�È���/$���wL�yY���T�U�׊�PA;y������Syou/&��H��0�&fh��eg.����wk�/Iǻ�c�u��h��:�ֶ�<�O��y���;w�Er߹Mm�n���f����3`�&��{��P��-}qW�{�>��9���R�/���宫��/?}��'�#��� ��H)N��
����P���p����m��}�h͊���;ٞ�<x��۽�ϙ��S$�Q�)���𮊕�{L�3��1�/i���@�Y��(8�_I���,��2_����$PW.zl̅�Sq�K���[<���^wo޽�����-6���O���IѓМ��Lz4�2OGN�����`c�*�������k5�^0|�^����졝��!����_���n����/^T����2#Gg�3u�vt�N����0�m*�7�/K��cE�o-�|�SӉ���U�p1u]�?tt���2L�u��뮻��s"��Y9P�#g2�\W��R��>Δ���
�~'Ӯ���^�9��Vr����%��~;Y�ѩg�_Ѳ�×�^2\�W�6jy���%@ߪ����NX�d�O�Ra���r�xG	��fcU݆���	�6v���\F��uc�~n]�~R��8�����ɜ�s�+J��d�ðp����\.�wi,ɠ]��" =��[/�ީzq�=X/y�q�%�T��1{����'��˯M{��׎5�;4�G"��<����8�zg�/�=BgG\T����f;�h���嬯�S�ş���c�m*�X>�t��R��|��1qީ�qe��fP�-����9z�n�s�.���g��u�Ti��ʐ"�*C<�&y��{�)�q�]�\�>�O'�|��g{��M31l��T��{wHR����^��zg�$�������z}1�~�g_��zV�z݄��rQ�gI.�ÀL/ECn6�Ĳ�mEl�o��-Nϕ�Ոɥ7N}}��f�U�.��m�ݰ��U��Ԕ���p
G���.>V��"�N��9sU�5�v�/�3�=�!�8z�ݑ�摚�L��}�G��d*�l�Nn�S<����3�Gгؗs����C�i�9Ͷ�9��Su5�3"��F����m�����T�T��,U����r��uӚq���[�F���	��,���J�u�_:t&��@��J�&�ݟ�w��p���Tn�Z��*�9:��:��/������ 1���`��`�� ��01��S co��1��# co�01��� 1�����m��cm�� �6�0�m� co{ �����m�� �����m�� ���p�m��`cm�`cm���e5�I� SK� ?�s2}p$���������Zc[Z֛V1Y�X�V��Э��Ѭ�l�kMR�ְ1��ͳ[UZ)l���E�X�ki��mV��m�j���	U�[Z�Ze�[["o�I�`(!�8��[Y��e����&k7\�ۓ���ku�n���j�mgݺإYZZtt�m����-�Mm`m�R�����>�٫i�jk�f֣Z�m�f�[f%k+F���[d�d��JSF*���i-,Z�R��2kQl�ޙu��5T�l#R�e*mZȵf����W�W7�  6��:�]��w��:ݔ�볞�z�Iڙ]�zǯk`^�מ�kVܺ�u ��ރ ��kk�w^m�ZmĞ�A�+ojӧUl��^R��V�Q�iI���_  >�b���[{{GV����
���t��th��r��z�4h�E�    ��   PۚqѣE }畀zF�(��  �
�{V�b�[�t;VȌD���  n��ǡ�6�.��[v������V=�ocפ��:Ͷ�Z���X�m�lzu���x#�V�Y��C7U�5J�Tz��lk-��m�Z� |   UP�>����m+a��t������{�^�M��ڻ���7m۹[v��R�ny�w��T�Q{p�^�����*l[��n�ت�fUjkd��2�gl>   ��/��*�:��
[=�T�L�+Y�{����eBv���r�Y��q��l
����{V��E;���6���n�UNչ�-�fUJތmLV�,i��Z[e�l��   Z��!�o�m��J���[ާ��R�ʥ�������7�ν�f�SN��r��.:�if�:w��g�:;�Y�u��j)u�U��cYw��5m��m��Xccj`V�/�  s���M\�f�:�C+}�=t�J�j�Q�iRុ�Ŭ�M���on�]��n7t��-�]�Uv���v��SSm���v��gl�iF��b�Vj��ط��m�)|   c�� ����_l�㮨�]�\֫��j޶��E%���{ox݇��+��]4��{kw�+�[9`���\Xn䥦�vK::�tӧs���j֝�f��Cl�j�B����  ���ښ��v�Ν�N�m��/���q�n��ސZ��Ѭ��ʝ���f������i��h�������w+UIo^p����q��^�[Xg�휧�*i�54���[Z|  �﫴���m��=^^�u��g^��6ԥP�v���cT��qX�P��[�Jn�=4.�ۃ�p�U+�7l�K-�M��l��f�{����]e;|���ʥ* �S�0������T�LSUQ=@ �JU  5O�Lj�T�0  	4���U)�L�hx������~����E��j/����H��lywڠ�=Þu��n�j�޻������K���$ I0�		脐�$�BB����$�$ �w������o�|��j?�vo�r��5<�l��v�X�jn%e]�/d�:Fk� �d�(c��	�hʷ������2�����Y��`E���O-�B�܏�b���-�$�E�đ-,���2i���~.<�ܞ�bE�qP�=	�dv�.x�@,�� 3-A�Z��鄔����y��Y��Wb��P��H��N����䬆���b�,F�u���6M���3>H�:�l|�	����ّ�Ev݈A���Wdk'�vB��D��{!��3 �F�g4
��Ce�ʼ����rP����V���G	�m���%�/kAPY-��c-/%ϝّQ����In��K$ڌo�md�����T��Y�(�ֺ�����Ѵ0i��(f[��t��L1cQ�v�6�����;��Z͡X��v�����-�/.T.�w�-�]�w�s"q��\n�]M� U൚�b�B^mh1L`e��8���EL6?�u�Ýt��ZX��u%M��i�0<*���2�k��ȃ�������Sc�!�4l��>�� ��X�ND�3rOn�3m�4��&�bCң�72�h��ט���b�/��a�u��Eΐ���/~4�o��:+M�"a
`ۘ���vDyRmb�n1f���`�dMZ��R��uc�6+q=�V�u^�Z5�-�5�m�x�M֣�ʭ����0��4��L�0a�f��Ώd����a�u�,y�,���&{��1C�me�P�7̝�S7pm�`�,���ÄޓM¾�M����p;���cR�R�D��Fg��~��k[ɍe��؞n<���[�uAo"�$�Đ7�>7���f����{�5�qVe:7��,�o�a��GY�˓�|���zGX�؈D���+ovm=;��yG �9���h��4�5�ɪ�:������N��t��`Jz��6	�Ʋ*ʹ⥓1���Ff�1��a�{c4}������!\�Y�&�B�`yN�J��h�)P3��J��j�x�����sc:��m����g�ov o ��3�*��v��Ɉ��ţ2�=�b��� ��M����f�@�c鶦��$�l�A�F���!��~��Xݾ�Ofk̶K�!D�pf=�J0q]��t��c1�������x�]Z�v��D�>t��2,���IM�I� �e���]��l��Q膅�,^:�V�#]�����O�=��q��5��Ʊ�5�*�F��4�k,*��b�Y���P�r�oIՇm!�(�.��AR��:�xۗA
ݦ��T��J�c�M9w��&���WF�����Z�՚�5R|�@o��Db˺�xe�����Y���ޭ+!���ʍ�2�\ߔ�t�/���3��׊]�Z���VXnEĖ�4@�9oqmmfkG.�aB��y�� h@<.��n�J�tIs4���l�˕M�:�
@�Ɔ?� ���s17뻾*����ٸ=J��Q4D�����i�x]�	-z�mlN2Ru\�u��ad�P��AN���-�Aal� ��U������L�KШM��dQ��'Z�ҮR7��f���)t�'u7t������F
P�P8�U�J=Z*$V�ۆm�V�N��t����"ݼT�1�q�.F(<v��բ��M:�+f�1�X�L��$�{B�`ф�lVO�;)'�ܑ-��;��<���DE�F����j�j!�Ub��Ђh*߮Z�-��\��4^ݩ �\�����l|��=T����N3��q]˦u��m�
tU��
�EXZct.=m����r@|$��U�zh;�D�=V����[Y����n1���[�l+sf&�J���v&�O8j�k˴�jdZV,�eC�Q4&nl�U�nV����z��-d���N�ʚ$f�ۆ,���CU�]B��_�݊�L��܀�Ȋ��3Z�Wd�+]���p�r!Jƈ��c.�����۫m)
���͡	A)Y,P�``�UӠ
Y��V�S���j�Ķf����E����֊�����դ����R��B\�f�z�7�6�&�T�'K�kdOI�S6j�i0�u)ٰ���އ���OV��ů��9�FỽP%�&>x��3!�K2�.�K� E�1L�콱���7e�d5�sf�	h.�}�r ����ǺH/��w{A�6���$_j��	��85�ƤAbh1�X3Wui��-2lk�K^�wby
Ӫ�dd�q>BYR��PIn���Y1�K��M�����6.b�RI4+d�����j;�j���,��Y���HnB��e���r�˫�t��R�/H���o�}э�sv)7�l���a�B�F�9���0J��U��Η�\Ahgۨɢ��M�F���˧�7h�K�^0M��5.)C��Ѝ��舭Qr�Y-�S��+Ul:퍆����KyLe��WYF�H��(�x�ڂ�lwW�aH!3L5����CK�֮�����ۆɣ�a�g�f<
u�E��.���Y�Lt����1QШ���@/�^`@a�Ŝ�i�x���z�u��`;y���n޵*ق����)Ej�d� ~��3��,T�6Ql�k6�_���=���)�ؑˬ��z ���:��1�M�u�@*�%n� ՠ]"- 'B���iU��p�w!N��s��ق�	�.��~І�|���w!�I�x.֡������L��%�3E8$-R�u3�`0/��7��Dk�{��a�(��r�̢I�ZkvZ�O��i��z)�Yi�@],�thm�N�ؤ�@ٹ���/A.rࢦ*�'�y VnC�\��0�R��:҈��A: v1A6B�����Wn&.P���WWgPǭY9{/r%n�-;f�V����NV�P�N}f\;��*�7V�TH�1���6��CY�.4�U��N5�<o�5�m�7��3үQ����;�Q�ଷ�m�:h8�i��˰z���h�DM�JL��Fl�\Qı�Y�� �Q���8R�����������f��/rB�ʵ%FT�[bTF�.�^A6�E��Ֆi *,Ϸq���-$I��р@u=���J'�eo��ږ	/B�T�30<���rFJ��7Vm�ԫh��6��ZשE���y[z�BZ�����RK.�˃2�Y@'���E8�3���,�M���شc���S;{��FwRJ�ݡ�v�3�-�e�JN&�Z�4@ʶj��Sǈ�����B�S�(В�'��F�/��'�ږ�c�uPl����]0s����0�q�VtR/����֒v�U�Q�+	3��)���^�I+�9M����F�8I��5�`dOh����������O�Ԟz�y��&���]�bN�4%��@i�6��6P�	��h)Q��r�r�-	������ǂ4��ه�w���J�/F㾺X[p@��$��y#Y�} ��s��[u��[�J��=�MD��
�zP�,�b��ұ�+8�d���)�h�%J7qڶDٷ�����O=���m[�h@��ty��P��A�(d�w����!�,!H]fZ�i��2�޿���1��&�#p@q�wgIy5�&-�ff2�!� ^�qV��nMܫ_;	�a+4M$��l��������3�^B��cX&hBŽF�%J�f�㴖�`*ОdJ,���0��x�+�}Qǀ�h3[QQ�G��q�$�f�/�v[���cC�6L�˭��jtmՊ�Ulׅ^TԶ�qֽ�QR�P���aa�hK!XjMJ�u��	����n	C.��Z��xb���5[�%---91�cnasrÉ`6�L��C4:gtj�'V�K��īV�1�Zڥ`=�a}��^�kt&�Ya]m	#�K�(栘 �S#�[x�"x`��z=tE��f "Ք7D:v��]\�chQ`E 9�f�p7fj�+nB��j�u�*!vn�5�u5^�r�����S��D�t��jr���!ڲ�u�Xj=}2J�-�����hq��(M����G�6Rn�n�n�{�AcL�̌Z�,�������ے�l���B�<��͎�;���)�X�&��}��A:�^O*̪�l��u1P�vH�F�ە�,,�36	�K9��(U��:˔���<�s{zd�4�[.������e��7�HVSzrLR����1�)ks*cܭ�;�b1��;���M����y�J�}#�/+�5��:5���'le,��C�5k*6ݡX�ɲ"�Q۫�Y���X�3s�H� �U7&�3����zM���I|XW��c����5m?A�=���p��&T�����x66��[t2��ZԠ����%�Z��	�.�û7b{�!wf�02k&玧��l�(��=�t�~���a+�-�� f�����ri;�:��2Ù���>��bz�\Л�W��ɡM4$�0:x��'Fi����ؓN�&�3�FI�d�:��GTJ7~"�h�KsO�	���l��^?+�r�
�E\p�Ӫxc�������k(odQ�rdj4���
�x�؄���nŪ٤��)%)0�m�Wx�����R9b)5K����juӵ6���Ǜl]��X�q�6J�����tK�Y�&R�aQ[%60e��M�vKZ��KqffB�W�<Sn�	k��6��Ql�t�37iVlj�nQYV)��K��Nn��ʟ6�6Հ����Q�_#�vLZ�s_�:ߚ��wa*K0Cay3 ��t���[uIFf�F��xk�w�H̖�j��_ۧ'��:\��N��u\�њ.o��h��A�z�.����+҅K��&廗�'�v�cu�Y%�+-�uB�f�U�����ǣi�"6�u�I��j5`�����J��q�P!we�5�=h�M���ܫ߯�v,<�����n�3m�?Ji���豩��)9S���Dؖ�6aɞ�NM���ȜM?3�vIG%ܫ�[�4)��t+��56���y�a�7RZl��n��Z)�
���B�ov<�MҤ�f��-۳m�!݈S@��@"�݈���=���'�^���{5�0�5��$5ջ��s[;��F�,֫sv�(fVZwV�5iS)n�n��$���IKp�^fQ��W�\�xLOm��352Gt��w��3T�U%�/XhE�v^P�m	��rj�5[U�l|*��ow-:�Q޳$5��p;�M�2�1��ۻTdY��Q]�#5�F��Ք$�h�/Z�(nFͨ-O]^�
��E3Xң[�\��փ�O^T�80

�w�c�[���H�
���QJ	���	��|��'�#�w���M��e����;ϕMԂ2ݙ0�J���qb,PI��IB�;��^�Ěe�����b`!П)���ꕶK̗`�{���T��OX��3Z3q��Tʱ۵	�`�V�f�YA� %X.���m,u>�!=h��(c�Ȑj���xd����r\_M����i����fs��%d&eԪ9�uvj�Yƌ��CZtr�8���kƐ�Żv�/H�N��,�M����EI�h�f�7�ⶮ<�)Gj�,N�Y�81�u�H�㡻�P�>E�����͓����F��݄�[j��ac�FCv�dtjMSJ`�/kt��j�A��z**ʮ�hl�϶ ��������5��(խ��Ԕ�`����Ū���*�54H���ջ8�a�bE��ͤ���
(r]~��K��v*���24�2)&��eIn�Ԝx��%�3��M�Ԧ,���R��h��y�I��ˋV�������خ}'D��v�V)�\`��<&���Y��R��XQ��U0^�$�*4��{��M�V�1b[+C^l&�Dč�w�]��Op�5"�fZ�j�kŮS�Q���l���f�T~�/f"�8M�*�'��8[1�"x��5&м����+s-�4��^��ol�-9b�X�a��ⲩ��Bw]����$�^7j�d��me�Nز.h[HlT�����R�P\gF�2���b�D�G��.�$��x]�v��l�U9*�E��t�S"=�.T_f$`b���VV�1�n���I%��9��KKPB�h$jK��D��'~GI����7���U�gS��
����p�B����X�	 &%���%91�1��l�dݞh\2\9�ի +�{/"-hw���ql��/�b�y%���6��1ͭ�2��"�Me�ܠ�+/^/�mַ!�`x�'bMN��BWsQks���pT֪�l�]���W2ڄRz#�Գ��j�~I��	W�fD�Ͱ�aˋl��Qe���5�	���]&c�ܩ����Vj��X"�٫��Rn��.�/N:�.�EU������<CT�m*T]a���S]���fϭƳS&'Y��Jv�)���ָֈr=�D�N�Z���s%i-<LZ�rPj4���2�#�Qш�L��7h�ڼ4�Ɛ�)
5�#�p�*��r�c�m�Ø�i3,�%�nhT4�a�0X{O�V���զ�����Rv(ƚ����մ�*)�y�n��ɷf dO&ꖷn4��	�K��:����yY1��VPK)ˠ���m7�|�'^A1i�nz�GS�J���z������6��ۧ�K��K���vL�<a�b�GW3-���W[�"Ԇ�Zeu����F0�wu������Y��M\_�V�_U�q�dFLc�o3�b��.�)�N��Z������wH����*�m�H�a)�]�bp�齌���s��7%'Q��W\��o��k{�A�:��"vN�+��&���2n�
�s��m��]�Gaô��[uϤ�/�ʚ�t��,Z{�9x����\�;�Ç.����:T���49��4�f�\���,c�d��#1绬y�{�Lkdڐ�5���A�k�6r�AL�d���Օ+�RQ�ɬm�#��y�q��^�+�+T%��O�{i�*��-c��^E�;�g�mh�'��ջ��#A��l��pg(��}�Y�7H�掫��n�H�ա_&+�d/F!d����3�^]x��@烐��A�Κ��s�����E�o�̹�vv���	���j���7#��1܆[�s[X��(�؍�gI{���<e�����Ho�}4D��9���t�Q�ؐ�7 �b٫6�W�����2,�{�s���U��J�Mٰƙ^c�{�1�N���v��C�s�9���4!�Ľ�^�^�0�S ��{Ǆ�Z�>��`�Z��ȭ��T���w���;��7��u�廉�[�YP�����[�)�t��K��!,���ہ�V�������<�Yb����J�`��ޭA����L-�w9t'[[pP]C+Pղ�!b����ӝ�!�8�h�ヶ�Ϲ��̷�[	�RˋJ"�v���k5�&�v��D:Fa�{��ϳX]��(#n𮼨�o���H3;��l�{Əo>��hu�)����F���$x;j��5��6������uî�>��"����rt�OU����C��D�,[�;v6qۚ{�s�hV���T����xfv:=�f��n���Yx�=p;�	 I���w�]s.���3{^�1L�qI�)MWӰ_w��+L�[�N��ݜn�i�����m��r�n9C�)�S"�'n�5G���9��6i}�����h#]��X�B�R�ܛoo8�i��f�D���(Tu�ep���U�n�m���>hԑ�,�, ��c�3�:��YAQ�#��o` |�T�K��j>�����*tf�ia��ni�`�י:ŌBp�\���Q��[@^ʝ�7ϹM�ع�*�2�!ϸͬW�Z�w�._�1���=q�L����F�n
��:����]:�h���qVC�c�XmR���O1=�.p����t�V�!O��m�:J��Eh�,�/e\]��W�m�]Vz��\
����kxt�2�R��]�v��Z����-g����놯w�|Fv��96�ru����L>S*�\� �v7��}�e�V��u�=\�}d���u��ij�ߣ�*��x�P���n�]	a /$�{�/�yS�f�bZ�%��g䲋�t�WMԘ͸0qT�t�3��!wӟ!��Â3s��*��;�����Xռd��׹8lY��B�;�E�h�/�������շ�l[ワ4��2�_��[�B�_ �(��t��'F�4^<mc��H};�e$,��v��F�I��!{��g�v��-`{�w�Gd�{^�Fb�J�m�$s.����e�5�V�!0�[]��� ���I^�S���j��;-٬��L7��Z�go�m��c��<��Cw�����1eP�e�PfkFj���u�Rq9#Z�ЇF�t�l�q�:��S,��^�ƸJ���/�$Qd�w,��e�՝��WY�ދ�3o~���k�4�8��r�;u��Ͳ���ía�W����Ҥ�	�r��
����&V�N�n�d�y��M� ����{��C�nr�Luv����h�nP���D���H��|׏�'M;�%����M��UI��Nu�{C7j����"��t��肍����UpC.`I8��fv����O)�r��IZѽM��ݘ�%�gƣP�nK}κV��kK�D�wn�qmXljcMɛx�ݮ���wXUc+n�H��n9)qkF�/�����	I>�j���GI֩�"��*]��sn���y�^q4]'�yX���(`���W9eGӴ9�X�3��M���uy��g������}�΋�y0.=��o��ӰEϫS|����C�zr�!�W�%��g+`��}M��LjV_4����^qZ�	�w����0���� kjM�8d�33i|�WS�C�81��	��5�/f�0#�������e�s�X��8+�Q��ͺ|tΝm`�ՈbԻӽ��l�=�a�(���zR�ǥ�����#�GAg-�D��.��-���pa��e��5ՇE��D�)�J�/�iU�>�]��X��T��5ob;y�Cs�(���'ٖ�Xnr�ɷ'����5��[ҥ�gfpEj�C�:0�hGu�M.�Ξ@�w��$td9D�,Jo�|�ve_[rPr΄��]��������g����Y<O�<�"SһN50gRt��C
�&����F��E�V�F^�yH�iop��^��ӓܜ�M�yυ:�``������dݛH�d�8H�A�j�}W��N���v���:3������\U�>�{k	r�S<: }o�6Y����)��vj�
ܺj�r/N���*?�*g�R�v���=L)�'����!ΥVfe�)�q�������`�1k}��ԣd�&1�9�w�	ۗ��T��yv�!�u>����V���c�0�����fގ_YL�8Ë-�q�ζ�VbJڶ�B�f�ے��#��F�J��'n�������p �xr4����n[�^}͊Lp��wW���f����F$�쾙�	vY��R:u]�0�=�*nT7���p���"���N���p!Y��*�νtn�������}9n���w�]�Ld�nRel���B��J�Q/�h�	��F�y�ת֔x]��������x�<�����Ն�v)$;/!�D����N��*�[��@7�^h�e��O�M��gf��{����F=j�bH���xv��ȝ>),�.C��ts�����in.�or�B���U��8(��·N:C]�0N� Z&�2�Tb&>A�A�NU�'e�:�*���K�r��U$���(���b�\21�:�{�E���O;�5�z<|1��Y�l��u&�t�%n-�ls��t�ږ�pV��1�!�T�,�r�i}��9Be08�U���p�����U��Z�}�Z�R>�Z{n�l[�=%��"�S��X�-T*����f��������o�7=�z�����d�#��÷���Զ8Se�_vL�6\��3v���YqJ��@V��g�Ԝz�ŭ��Fҫ�0`�`��.=�!'�s�n\QSt:�=J�q��%u�(DV�f^����������8r�<K.����AW_-"���oR���yw���o�ޮgc�Z��������v��w=/}:.��r�"���ϻNSd���I���n�.��*�Й�:�Z��	�\:���<�iR�]=�ꯖ�xd�퉊��[���m�㈁&���$Z�Z<��̵,⨴����p�9Vͼ\��\��"�b����y�;����X�j�5��Z�t����.jOq��3z��՗+��v�N39�@л�ӈh���:�q������ĝc�}zetў�	�0�������mQV��(����Eq�fְ�Vf���涖t�kT;���ı6t�y�d�v��nk��k��k�yw���K��ޱ������BI`���*kX��.n0�"�}�[5bz���:�������z l��zu_7.2�9RU���|t��D��䷋�F�%k�l���S��������ۗ�v�'�^�#��^Y� /y[&��ͨ�����&�f�܅�d�q��kp���=�ˣy�(�����Rɯ��+��9��s����곶&PZ�VOrɋ2��{1x�H��U�%�us�sje�-�y�aC=�%$�o�J�;�c)��rY�s�m]�d���� �nVc ���]3jo7�����%��{�k�|
�� q�!`����[8�Xm.��L�Oo�v�$���䶟VV�u�(Y�6Ŋ��ܻ�_6v��>����<��Q��f��P"����j�n_h���y���յ湾�;�YC�ޱ�/utq����1�]s�<��ݜ��c�5����۫��ܦ+�8�5ָ9�ӏP�^��qĠ쎓��Q[i��yv�K�n��w��.��'_[7����m�%\�jc���{Z��DsY�(S)L��>J��,V�w)��j�3^�B�Y��J�魿y#�mb�7��\&"w�~ �%���q���ԧ*ۇ��m��C�6U��3M&�lʻ���-\|��a@TEK��wDp\�Yﴛ�Q�7s���4��
ED!�]wu�.��<�S���rk�ʺ�\�]��]�U�z��JT�B��}�[�M��*!��2:�E��ew4�3���Y�L˛U�;<Ԥl{y\�s�1)�|�u����`N��Κr7x�5��zX��oso�ݠ$�5�%��iA	��%��S'�3�Цb��%��9-����8�SN�t�G�X���y��3-R]
W7
w���:���;�q���Jn�;�j�t�qE���)i�p9l�0�Q�$=�j���@*��|�\�aa�n���3i��x�v�.������3[5p]�u��4}N��T3��b�ʬ�����C���\3U����2����&�;Y��9]��S��X����pr�>�{�c�5C/�;��;"�^�=8>�J��뻘����u��7a]��S*®r��$��a׽j#1�M�7�{k��;�Z�q_p�.t�%0_\�׹�WL�,U�j���ovFBD��a�1�}n(-T���(ͧ�n��u�z�����N�����*\n�nS�QדJz�^������=ť,�Ob�������\j�A*���B^��AO2�P�x�F9t2u� [���U��Q������J�	��Pa�;x7�3��Tuu�$v#֗T ��	*k����$�}��ԏG��9u|4\�~M��o 0�׹��Wws_-��w����x���ƒ��4$a���L�Ca����ed�����xcNn)�f%0e6�_���0�Qد���U��Z�^�S^�)m+�t���lXb�!;���m�"Txit��k3o#�y���ٝ�Hf���|x[�w]2k��W�8v�0�ʽNi�y@��N�!3�7��M�.=��_���fQ�3m�d�dق�'(U�wvlՆv��nM2�f�5(Ζ:�w�_?��}��7���G:A-Ӊ�{���V/
�5����G�:�3�MbZ'!��"��w^Ø�k5ºp l��������z���0������!\[�@wX��l!����Ղfݓ�x\��껋�9n��`㠡�]���..��Ⱥb�Zd��Iڭ`�e�l��M
w���w���qh��g�u�F��+k�wh���o�+�h�z�Wn=d���s�t�����*��f:3J���M���N�u��Ρ��M�Վ�\�O�^��b���Mѳ�>[p�1�<qڣ|�4��Y�u��4��@nG��a�>�1��:1s;w9a��$2t�8x�0�wls���ONٷ�5sh��{�S��C����\T��{���W'	4��F�v/\�Bx�ؘH��{��:5K��"�Vn�.q��u���E�}��;q��R/��WZ)K�39�VC�^�)��P��W+�y�f�/[�j7 c�ǘ��rxVwOe�cb�𒮥� �7ݛ��PZ+*;ﰄ��5,W>;/�CB=r����x����%����0�e��4zѲS��������G����M+�:.��vP���A�P��og(�X���.Z�'6ѧ`��*^�J�^�Ns���I��(��$7��S'm9)Vf����4��r.љ5� ��E4ohy`]��+燻�=�n�Mf��+П)Om;7׵z���T�1)�K�,�ӷ�o �p��\�s�Nv��+��҆\�w��z��ː����H�v ��X�.s�Nc�\-���8/����QԮt�Sx��r�4˒�����uY��A�<�ec����,��Ih�;r��B�ü*��+��ZP���Zv�2�҆�s"��|��������H9pm;�7)�)I��J�s���rco���ut�;����!NZ���lwi��u�3��=ԲV�ƶ���Ɣ��Z
����݃Fu�ݾHK7���ձ}Z@�aK���|���LɎ�b��k��"�d��laƹ��{w&N%^��ܖ^��ݻ<1���]���׶r\V�Q��̗D�s�;�9���F$UءrR]�.��w���p���ғ��ئkd8:�"jrҰc�_6�����3������c���H�t�|��Ӻ��xo�3%x4h�� '�vz�>}�Н��|۽��Q��oJY�!;9�Kz���}��N�pj��s$��-vgz�gS��9�*�>z뒫6��
��4�9��Z�P}��K`z���4:��ݻ�ǰ_[}X��0�,��s5�VӐ�4�/6��;+&uYw�v)�U9��̣�v�y�E�,Q�O^�Nwi�9({���rﹽ=��>��@���h���z��Yκ\�]����or�zQ�/����e�L=Ǐm�o�7m���{9�׸d�˻��
X{�雟Dzw�S�+��0q��S���W���y9&�´�S��y��v�	�u��^wo�B!!��IL���Z�th{znMU��KV�V��ۨ�c��b�B���u̓�p�5z��=�;jh�����n��j�ۺN�l5����ض���a�Q�wG�3�>�����ו�u��#L<c��v˜�����ۻ1�C7�ۢ�C��[r�L�:�VM��`|�5��cC�0c����3sD[ٗ��n�����\�wo�[���t�N�Ɗ�-��ta^��h��+3/swZ{�,����uchAQa�s����<�˔��Jܷ��1P�������g3��	)�����4g1�?^^a��%���9��R���oW�
тɗ`�J���i���
�g)��g,3vp�{�Jn���T�z��l鬳�ir���������~Z|:H��껂����:w�!�%���(��[S�/���Rdv{Õ��1���d]CFxJ=�k2qǺ���f�z���S<���ΝɳF�:�DD,%X^�S�uM��=��4@��R��)�885��N���������۲��T�}1���`�3U���.�f��%�g!��m��Q���뷃�F�c%: �� �����Kv�6�݋.���4�V��J�͵�ˆ�n�%�k�'�ek�U�'<bؙ�ܺ9i*h��J���$M�OC�<Y�-��U�X{OT�zňѮ�9]�ک��<�y�F����B.uq�:�Ig�k�۴��@��;����\�^7u�]�0�D�����ٸ]Nz�Tl�)ҝ��6ꁾ���/�t��!{���f��9:���G��,�Ɨ�D6�Z���,=(��ݽ���"��;�7�m�|�;CU\��m��w�Ø{�7�=��6���c9�G�s�S�,)�+`����`�&�4�d�l�[�T�)<�&މ׍Gh�|�Q�9.��jM��I��:8�@=ܭ�06�+H#v�{@IM���R��� ��&�2�oR��V����m�F��Fgc����2�@���$�3�K��Z�Y�U�
;oY�wY��Sy�2�[�d��q[;I�-W2��\8C�ً3�H)�oL���U��s,
�YT�)̔�##(|�EDn>8�����}�%�C�9f`�:��vOhڛpRѵ�6��M�+�W�a]ot���E!�(w�`Dc�E����O�ً�'�x'PY�\�O;=�{7��Q��5�l��z�L���U��\�!_r��Cso���Q��X�H�P�����	ǻ��M�'si |9��3
Р�/,�Ԩ�(wt;��P��&�nK�=f1D�&�5p�-��˗�U�yxt=t6.O�#�A��]��g�*&�z/-�h�y���C=U{&^�[e�Z�f�Ιuv��6�wOocæ&�ݺ�ڝ}6nʷ�jv��;Z����c�u9��R�kD�1S��VM���֝ɭ"��S��لr)!�71I�E��{;rx����xЛˤ�SSS�+�	��ν9�p���=�=sz,�C�vg'7w(� >�f�*>��K\�eX��[f����Z�	��@�{�p��J��r�67*;K��)P^����`LP����jD�-����o%J�h�W�/4���C����|n-7va��guB]ܓ0u�5��Y�.Q
�nP��e��i�ʜU�Y�RS����;F�<��{wR��ڎ��-5���17)|�Ԥ6��ٓ:��,:��h�����ޤ(I;�Ρ��N�#*u`��fh,�9Rܺ��N)f���D��D({��j�s��>�J�N�SK`Z%2�܆D��8p)v�}�!��]���Ô�o4~��\��#7�LQ(=��^��:��cP`������y15)�Y�.��{9����J�KkD����m�)��.p�L�[%�dz-G���.U���0���:�R�'5��@������s���#�굔��@�;�	�̸8���Y�:�z*ͮ�2�zc�m�0Ci{���#���7q�y�
˹O���^��Y�KU�I�1V���%Ɩ�*`��b���&bU}c�/���L�2�>�r���Ǖ�qW��Bi��� �M��|+�}�����f���b����4��im�Z��eEA`}�xk��=;6�zCJl��:�&;�G{>�J&-��`���$�n�7�m���C��Ł�[I\ZGX������؀)���j�W�Ū��s�[F��"����it�sg�{m�����k���"���O\Ք�N��;��ڡ�m�p�q�0p�Z)F�1(�E��\#{��X�)��2!E��f'�; ��Z~��,f�&����[Vr�hD�۔ԥ�o�MU�̉�Z��.���DQȝ��ͤA#銸H4�Ք�U��N��{-{[D�;�����]�9�Y��k!e�4�9��*D[�&CNv����kj|��W}C7�9$S�+�-��f��!a Q�"J]]�(�S����OQ��gxV+ټ�cu`�$�t-����ڵE僷���=a����?�Ak�z����V���ZKm�	R�Z�D.nR�@�3Z��=V��W�묻vC�k[T��d�A"Q6��^=��n����VV�$�\*���(��ט;�mrYK�@x�}�v\)��͙ݜE�bD���+�ԅn���Vf\�Y�QMF���]�^���:2�O���jn�k$���
Ho(�Y�������.��j��\jn�����_5R�d�4�������5�p꽥bP%�%�Nm�q��?vt���ǬqA��}Gu�%j��՗�Z2�x���Y�v!�Т�&�lb�����]����9���b���\ϦH+�/o�&�:yХ8vV0�4�e���Һ���м��S�0�T��-l�M�n��5��(I����ә��r`�%�s�g1�rZ��y��v>�j�89�ڍ��ƞ�s�{d���!Z�$3��;��[���+�B���򲚊�V�-���;j��;�*=��a!о���X�4o/dߞ���6�/�<"�}�֥��]ն$�Ǌ5�A��x��7��Wj֎��T:�OmꔉˊMb�£��f��Kn]Z�?�N��4�,l��0b�o1�VRftWCQ�{��}�0X��^!�ɱ�� :$�s�u��v��5��9,���KoS?+ΝM���t���7��!Q���k�gʾ�h�V�O�.� �U��Z�o2�Kŝ��apP�`KF^m_Q6�ގL�����cfۜ4[$Q���];��������O4;*�{ �pgˀ0Cy�3��
)����}\��ɘz�n,�	k���2\� J��n�D'���=K���VwL��a�g^�\�Tَ���笍��X5��tt�R�e.�ᙴ;s "�vNk�{x��k_5m�^+�w�	ȶ,&��Նr�2��0���R���6�2@��1�����'R]Utz�Al�ı�/)�M���R�;�Bȱ��0@|��)F���8�4h��c7��[�Kw@�M]�5��9$0��3�m1a����];���*4����|=7��kE�X������5C��՜�,:��͇���mg6���+�{-V�M@�ٗB��l�!*�B݋䴶+w2^��Zn @�����jQ��yo�I�|l��n&Pw`&h�/*j�JX-CZq�X7��9ۇf{-P�f4ԧ:�U�P�DҤ/崛�T>�r�
��7���"����X�P:�^AOO��O.�%����W^�u�qwX^*WX5�e���e�.oV��\|l���K1�������D����u�,aW�X:!�z���s���66� �yg,���N��>�%���;����{:�ٹ(%�i�o>�Xf�.�J������X�u��I�%�V�E��ʴ���#��DRg]�#���U��]Ůe�s8��Y�r�2���^f&�88�=� ��͋�+�[1�Sv�b,��޸v%�e^ �;˾�pE���鎨rP�By���������4Zg7xrQ嵜���*��W`z�y�1���sy��٬�����D�;�N�vs����6]:�ی��x�o��Vk�f� �#�V�8`��e���=�&}׷1�A7,^�ևC�����X��)$�>��0!K�c�}��K�oB��R��S@J��[�fU������o.��%X��k2>�.�CX��p�0P|�.H�ե�Û�NB�f.Ә�R����s��Cg=K�"�-�۠�o	���W��i�V�����.��3�kE�1z(����V�+$k�Mgf����o�^-n)��{՗\�{K��=�E� �����ce򡯫^^MF�Y���;�:�� ��N�z����/k��SO8�:�4�� _\}����\Y��:�Â��<+7��k+�N�}ݰ`�Ɍz���o�����t�S�;N�0��գ�{���йb�Z#rܫ���R��yr��k--6����_ݱ��T-Ww���������g>��7�d㢛7}S��4�zp��X��oePm��[��l�r�mR�3޳��Tj�N��I\͊.��{c(wg�r��.i��V�7�y�l��f��Y'�����o? �(oi�w��Iv\f���)�h]�Qɒ寃E3w�*	Qu�ؔ\4+Yڏ�:];(�QY�X��FVmđ�&�c��� �N՜�8�
�9x�^v'ʚ6�)3965A��+�޼�r������ן��&c7Ղ��ʙB���Y׻#�ug�����c�.T�/�%�ir�"��nn���I��Q�F�����98�p��E���F���;:i�k7 ,�ҩ�_L��pe��9W4����c�v<tfpp���]B�%���j�Yκ���b_#;~]F!��Ml��W̮q�\�{P�ھtp7���Ѻ�Ɇ)
���*Һᬯ*tg=��wm�|��2=o�z�х:�꼻�E�]szeD�osL�U�(�3^�Sd�uv�ZC+0�Kd|������fi����I̜�C�����j���3�T�ݝ�ݕ�LW��a�Q
tE�ۚ����1N#t�:�=g_+ƗQ<]<�R��h��;���z��@;����8fU��r��n�
�H>8FN��S���]�a�T��֛*�(���iV����(�ͮ��ٳiZA�*&�<��\/!�XV�
��L��7f��X�0�C��<�dc�;�����z�������p�6�X=��)t�%dQS���ҽ"�w����=��ᓳd�pT����Ot�d�1���hĬ�,�'Td+8%ʗ���#Ò��7pn�4��r�%;)��O<�o�R������=}�=ڂ7n�[��hU.n�o��QMI��4��ժY�C\���7(��#!��� ��-�i.������P�c@��9}҆��|3�]cx!��X�_�5�����n�Ӡ�G�\	����'C�W��3�+�����ܩ*�q�*Z��O/z�h������C	����M��Wˉ�\kj�h��r����]6G���� 3x�]�fM]�jie��D��5x�T[�f�g�6��ي�tjK*��!����qp���CW�J�W&��n�[�e�yĤL���+�����\��^k���3z����tї*'2[K�>��� �v�tRT���;&)�۴H��S^��0���Z2=��'um���[������԰�gOh����w6��쥛t�c�l�[omi����A���ە۸AHA���.w���vǡ���a�3
�$ڳ4-Dg<<��R�q=d�e�{��2&�;o9�L�n�p�L�;EWX^����+~�ν���̤�Np�F�ng]�f�僺�j�����˫-�i.e��ѷq��t��]�z�- �q�p�U>�h�����+���0f�wy��h6Y�Zݺ�G�S�\95R���1 ���V�rݰ���X]%��d�r-�ه�>�Thn���D�Hm�Z�+Bv��9a�*P����X/j��_�no��t4��\�=�z���.���XA}n8@����չ�����9��W�T=�V=��MO=>mg�.y-f^�:�PȺ��;a����{jP���P�޳/m(K�B��	Ǥ�@n�Q��� ޼��z;^5#U���;��B��&�L<�ְ�:p�_
 �!6aާ��Y�x��mb2���y�
�l�ú�k�J=؀/Y�B}M'��քc.�	���fk�|����o�1uMG
sl>
6w{��K���n�Ӻ���<�:ض�s��̾�s�C۳��e���L�w����
�̓ �a��;emLsa��|�xS���/�ƌ��fB��	������b�O��oR=4�F��L�:+������J���̷���Ejͬ!�}6)M�2i?(������2!���[���!4�4���@�y'n�v�z��u�W�(�;h��C�Tw��6�Dn̂�_:V�Y��H�P��y����L��l@s�_=�΄WCwA��x�u��4o�W�iZe���2����O����f��+ˀt���B�j.Uu�(���iU����w����=���k���*�.R���7��nHM�n�^Q�PS�k�l�i��[H�өv�]�����R۾�FB�U�T�=�k'@ԣN*�����_�yx��g6ya���ټ��E�uy��
�_\�N{�vP��x�]�C}Z�t8�/��r5yٵ���}���W�}|o���DF�>؉�#�>��E���÷--��Sc�U$����_�(Ès}Se�j%�=۬&����Ev�W&	5񬛛�Գ<Ӟog,�U��R���s�����eZ�JS�&�}�t�e�Xޮ[e;��®��4�l=�Kn��+�r�vs��U��\�����<�Q}�GCFTl�>�d/6{e,;صȄq2-��n�T���Ŗf*8k���e��E�ӏ�)��p�k�d�k˕δjK�����W ��_��ls��82�V�s]����0�E׵��K���X��H��s����ѥ��u�[S��yu����tHg�[s���?V���A���HϑRyg�+i�hB�1M�uyZGQz�9F��2��-��-.�{�<���}M��E�+�z�\tg�;�t�fS��u.SM �u���b~�uu:��^L2��Y�N?t�+��b�f�j�ׂ}fK�q��\t�����Vg��8r�J:���9Ǟ�ګ���7HU��f����� ��%�R9�<�9��AV{-}y�^��J��u��}�ٯ;��y��K���M�N)s��k�U ��PI*����<
q�sN�l�K�H>2a��{c]^2-�ߏ%=���YƉ�2u5q�dцٷr9��\�D���sHF[Yw|��7I\�[�^�����@|>�_"�1b�UU;�DTD��`���"(�t�H���X��b�5(
��mb����(��ьm�cR��"��V�m�T�Z�*R1TDJ�`�ֈ1m�hb�֊ԙ�DEƊ,���QC)QEQil
[\�+b�eV�V5,,Q��S��.a���ڷ2���3Ȫ((V��lr�[D���j̶,SRЪ�F,��l�4Q@��6�ҋ"!�QV�e�+*�R��∰F���-��mQ+*+�q���EQd�B��Q�(��fZc*�iJ�b��#m��R�����E�-�b�(�P�����m�|�"�
,QADq
+[l
��jֈ�X��U�V(�֥�,����"�1h�KmV0Ģ�TPE��U�XԴk���e�Oc��~}�������u�U�u��C���S��N���*�+ 
1�����:�j\1�xN�ʛ%�o��{�#)�� m���ωs���8��2.+'hC���h,�@�<5��4�J�������v�1��p��C�o�;P<��I���^j8EJN���j\T|E�s�5^��gޏ�g\�n����R�Ԧp���fJ�c�D�؍��9Q�!z&ҏ��aj�sʯw��t�'��?Yt�i��>7�Z*J��H�?q@F��o��X�|�{��YǪ�/Ҥ��"z�`Vs�=i�T�	gG�˗�y��c6PԬv�A��F��cD���-Ђa���#B���a��/N�������{Q�%���sE���y�~���r5�$��G��y�~����T�<Ƈ�nmR�c�����p�j�t����b7�����x;"U-L8Fu��HV��56E�]C�UG�E��T$h�<Ĕ??-����2��+���!�\]f�U�L{�:|f�K���!�%Mד��T,��b��j���ͷ��}݅��B��"�����J�����P�+��A��}�D�sS6A�� �O8��${��=6{t�-J{P��kN"�E���1l\�E�ar쮇�![��{rS���MrZt��zl��Q���7"����%q���js����m�y܂��1���MI˰�Z�YW�Tv`����Wn.��]>}#�M�j�8b����)m1�P|��o(�2!��X/��`q���|�<=�i���>�4��^O�f0�W�y���@��{��.��+�$�7�c!�q��i_M>�WH�����	Ѧ}��on�Z)ֻ
��G���GR����Qb*��ou$����Eg��+饲�&jQ�\�� ����ϭ��#��El��^l�Zx������q_Y��L
�d9��Ozzv�26?2yWbb�_��xwK�&��%ޚ��+��szvy��9~!�qJ�/Ik���5��9U����Ƶ�Vt2�S1$+H���7ۙ�Z�}�9G��dY�`�U���`;�wk�N�[3�Ƽ��i���6Nd2գ��3�IS^����Q�Ƶ��E1Z�}��y���:���|d���M�?�Ë[�W����!A��ؗ/	>2]T&�`C�e����g��(�ʾ�ЯXG�j��3w���|&�iM��э3|p��~:Um����.��f�_�+�uq*�x{���=��+I�\�Lo�NV�%�҂�y[X���+uXѨV]��,t��<h�b�p�J�,�i�P%�E�\; �Wh�g9WdF�
����h��W^&���4:7�(2���։�{�����/]��J�tm&�iD�Ӝ��[�N����+dq��K�� *K��c;�V�=mZ��{=���#��H��{��+X�<�5
���Z�-�4]=�͟���a}��K���5ӵ�`ʰ��l�m�6F[{��,C�
�U���[�^buSJY��O��+Kٹ�umOl�p�ZF�.��.��s0�=a��/��Ī�b�!��^��+|GD�ó�jww��d���Z��+�J���ʆ7�e��U���|Y8<�'Dj �^ .���mC�%:`�rn�r0	��f*�5�|�v,���HNq:P�Eh�+�ݷH�+R��7�{��{]9֏FL�ro����Vo�psV�,v�����{o�:��V-���v_c��� ��K����5AY�V����AM�aCEl�G>�oO��˻J����s�@����]׫��U�E��釨�Pk�h�NNKmQ���ܝ���,���;��;>tO�,�64I`����On^�Y�0���g,�^]gyZ�=�V垔�d��2d����I!��_E��W��\f!���(�f�^�J�Z��9jH�>ڵGW+Rަ�Vr�N�;�&Ȥ��\�0�l_��ɛ�Pbט����	���ޛ��U�������&n�.�u��0}^���.�b��{=)H�EO����=;��n�t�Q���W����'y��	�������HU�I�%��C8���>��}'�C<�.W^��[<��8�D�Y�}F>��C�S�d��`�U����s>��)����^͉�'��ռ��O��=�}�:R�}Q��^���>��'X�͸w���pܕR���V����y-��R��4*}(��6Lz	o�>�m�5}'�������[_u�E�Ui��G�y:�)�%o���z#�W�ˊ^;�6	�*<�ܩ;��-Y���"�yG�ڝ�)@
�x��!J����f��=�����I���v�v3ك�}G"_��I֘xm:��w���/{��5S5�/S����7�$�s�\�E��/�y���2��m��/�wQ�:�`l+n*~�/��z
�_KQ���y�%��o�1<��Z@��P_�C�p2�;���A�V�:'m:y�s��]�uu��eQ�X��.T\���F+�󑺁��\��V�A�p�P|ৠ�mK��g��Z�(G��"ޗ=���箝wn��[j�3Bl躹��5Ĕ;����w���!��Lkιsci�2T�Rlbsܕy�	j�c��k�86�&l��9Ӂ���[�{Z��}���eOR������l> _�٭F�n���ꚫe�O¹���5��.�]�r�=��yd�-��FH���}�����{]����2٦���=�%I6lx�U/J���8��NPݾ���3d��+��;Y�t����� ��t-C4���s�t��[֦Ӟr��`�����[��%�Q-����L�x��^���#�nG�T��K��3�ˎ�u�H;*I�wf�ޖ��}E,赵|�����f�{�����.�y��2纽K]�j�ڮ�{zV��xJ�1�ˮ�m}�/ūU��]�y[ܥ��Ӝ�R��ƾy^�l�U�o6�`��}�U{��w�_l�mK��qrq{�v��o�����xd��{�0j�^G4塝VGʠo��tff�8�W�ѕ�T�ϝ�7I���%�/�a>�A�:�	������,��S|�-���*���
ot%Cd-5���ā�IX��Ԯ��[�Y�\��x1�jb�5��X�;���\\�e�W���J�Oc��/�7UV�����7�|^H��.ɝ��$���C�����~�F��ʺE��0�d��T�u5���xnv�u��Χ�בngd��9���uy����qS�Y�<u��;s�s>�u�v5(z�9�����4s�|g'^ڒ����Ν�1�n�3��ռ:��n1��d���5��y��+λ˜�@�L�13/������7��[}�+7bo�(w���cω־��/�͊�����L'#��y{���o�<�]QJ|N��ΰx�g:R�8���a��k�-,]���M�<�r^L�f�:Nu��il�""���/��ߥ?u�a�V���׽��[�\'���ӷ|�{�'�E��9?S�~��y�G4N��;bB�%������l�s]�����.��k�u�}�R�5ʛ�U�Uf�2��v�8����>�7�	�r�o4�EDm��o�yu��g�sHI��2M\%�;�:�i�A���9"N1�"�!��r�Y��g��;��;b�������i=|
��S�8j�kyn����F^_d��h	�Ɨs�^���ӟb��j��xp�'yW����ުZ1*���Iq�H8=r�z8�6�M�rf�^�uZ�Z��x���N���'\���[KK����>����c�ʌ^S^j�ŵ�,>Y��,PG��k��w9�x���7�OeWH�I�E����-���%���O�	D�.~7���xﲖ�uz�'ҏ�N���uS��)X[�d3�g7y�$���������i��j��ޕ�R}�-����39��q����pjI�Os�5�J�ؑ�<��˫Ηf�WZ�O�c��5oB��Nc��s�עO}�wF�Ŷ}g��]��.�W�N��^6�4!���0���������=a����{O���c��G:�s��X��5#�$�SB}�Nr����lǙ)^�Im�
��9�k�D����\����}�����Uώ�H��G��fa�Z�o�r�K�)/݆l.���Fo�wVE�~޺N��%�<%��Z�f^�@�єvY��s�fWj���ղ���Y����<��9���Ll(�����u)ot���$*k�����o=���~���z��$��AH��<�+��_�ͪ칻M.��)��Ǵ�r?^y�z��h���r��yNܾ�S�o?zo/uH�쨙��ׁ�ͭ���Sጅ�p3�W�o:��5���˔����7QOω)�k�#��:_�oѪ�hQ�xA�ϑ�<�?}�۷C����u�m�u�;���}7L`�9�e��V7#�C��Y�Kf�}�\<U[�k�͵�ݓbaW���ъ;ݗ��JI�*�h�u��{���_��+C��n�w���y��;U숱�'Y��Hb���ev�l7|�~&�v�rQ�����z���X��Oo�h͈��'	Y���
Q�mu���t��y�\�v/�S��|yZ���䷔�T���
�z�r��2��:y]��ɧ�=��~�`�n���=�����U*rߺ����9�;l{�Q��i�wu�:gs�K�8B��>�d���H�$<A:�L�U��1�����ݐ�oct`}d�z��})X�+d[��]Ϗh�w�t�W���k��:
�3���t��n �Ւr]�J�˹K!wl�Y�����xg�w9�a�#�m��H��8�*y��&�rؾ�ð,�Qx=J?|�S�Y�����;W���^��'��j?N�^ח�ڮ-�\m%c���q_�E�p�/�QOl�/��O��.͌o����$�������.�]]ث�d��|����t�w(�)F��`l'�S��uLǗY*�UIn-�*����&-�y�6)�P�܌�f}�5�[�k������%���<���:ET]��mf�7X�!�������O5���w����S�^�
s��F�vH�~�E��uNSղ�'�\����ƹ�w�������'P������}��M��7Ԧ���}~��*h6E-�[�Hl����J�r�U:Y�&s¥N{c��~Y[�^�)��H�EM�R�%��=�\0wcg�N�7���3Յe1��fi�8E��J�nOP�:$�T�*!o�Л�ٔ�Rp�׊���7j��~��e�GՏ��n�(��{�h�ݗ�d+� Wg�i��,�&Ϲ
���,��mӌg#�+s��]��r�ժY{�^�tG�a�Pf��Z�R�c�{W�En=� k�h��s�i����w~�v�{+�}k#���f�9q�P�t���O:[�㙉�?-ٍ�jE�U���]�Z--G�ٞ�7���z�R�M:��o�����d���,J�1����oj,-_y⻖���Qk~�qou@p�'=i����D��Ib{�P�݆�������-�,�����K}s���[K|�\��;��z�_�2*}+S�©��$��d�P|h�����fVD.v?å�{��i�=R����]j��{6���7Z�}�|oM�Ԯ]J~�@�g�����o�:�/��ߩuyҮ�p]jqS�Yz�g�ޏ��kJ�#�^�1k��w���7<4���)y�
iu��AW����h�N�=Y�=��w[�i��6o%I�W3���5���'b��˜
�ԁ�1�Hx)��
>���~��蟫7bo���}D�^��_>��#���	�OMN�}C�1R�ۻ�*���mۼF}FFٽBƫ�6=Rcҳ��&�����}Ɖ���X�\jg�����*q�1#�.�+6&-;��dls,�|>#�R�Ӧs��RٶiᾹK�7E����<b�¬�F(oep/��:e %��OT� 7d�SwM��C`�	1�V#��u�Z��ήX�M̔�4[Wb���-�#��q0]抃�q���ý};�MKC��f��dY���Ȝ����� .�R56Zs(Iή<7�U;�a=��;�)�@�����C��:�y�ze�Bt����au%s���]��C�Kt��#�X����2���̐r�Ũr�珚�xIR�G ����umj��K�5�(W[M���c�.d3ky����Vjh�����wN�"gj�ܺc�����.��}$[��#�{8iʵ�PM����u�Y�9���n�؁���Iwv��Q�^W}�f�1K,_*��ls{h=���89�i����]�u�����ƭ��Q�iS��D�Az�
me�vMvm�5g�IR!d��%rㆎ�l�}�)�8����Fc��d���X���A}9����Ǣd��l�!�N�*�,<��B�2��T��˚�R�r_":�,3V&��6�N�is]o��pR��l{�s�`��_+���lwX����s�'��U޽�F�<dZ:ծg]�[��v�\�̩V�!O�,��
�$����V=w�^gje0�+޺����������-�:d�Uf7��M����{(��4>TfO��C����B�q�\����9p���Ht;*ut��z,���-��2_����BN�I��C9��vFc2�駞�O��@f�&%�g���嶉�H��펺��|Vr��Ą�"���-�<�p�eǳ@�F�u���^�ᮏ�7�A��Y��jS�W�'e���s�Bp��^�f,�4�[U6��#�]�j��U U���nb��;��u�����r	WݣJ�ӫv�W�u�c�T�����;	_p֓�$�釂@�pP8�^�X��O�uG�Z	-/:��_oa�gJ�qg��T\�J؊bҦ-��]/4T�fu����� xo|���z=�U13��b��죯R+��������tw#�9h�!�u���oq{3�m���ً�un�[�k�'8oE��f�y�m��f���_�q�A�\)�2���7�_%r=nE��-���QG���}8,��w�Eu,���әpA�RF��s�Q#��I��*k5r��K:�gRRr)��4`��طv��-s-܋�|�_q
𠐱֮��7��=1�*p��k��rԬ��(H���h{�1����b��`e�Pd��V��Ib�R+�:au��a���f.��J�d�Rw��^ɝ\�
$�_���j���,P1��Z�����UT[]�����Y�j���Z�[j�+lYR�UeKq�TTF1m�*��j
.e�jR�hZ�DQg�OE|ERZX#�"�4U�&&"�*��T��X�h*�F2���kQZ�9B�fd�l�
cP�UZ����+R.Zb,El�D��R�����V�Ҫ�Q�������*6�іԶ\���(�h��LE��Օ
1e��k�Ym�R�cc+Ke-��a���ZZV[�Um�e�6�F�%����ʹQUP��"����j�R�m�hҪZ��5�����F��ҩJ���m�he�0hR�
1��R�-��f`�UV���������*�%��{�.�>�����n�V͋e�mt���c:�uBQ�v��oY��7S�W�$+ ��m��Z��ٱ�5g�|�I��W0��8o!&�=�Q�Jv��M�uڵ��G`ck�5�*�]9�%��aףϮ��j���5�s,<s2�o�=���:�#�l�O
�}���֚e�bv�W`����5�ԸOW_M�ps9�w����9NXvw7�O}����W��6?�e���\������᳜��W������{���M�ݴ#��X�d��:_˦��QW5��I��7�s�]�~�g|�	Ǵ8�τ����{*I��r�h��^f��2r��t�y��m̽�؈�y�J�B�N��j��_ �TA�}�,�-b�I�ma8�u��|�M�Nx_���ғ���fx���͉�y5@7�/J��ͣ�>Ҽ}�gT��ϥ<�I�Eǻ���s7%��q��r?sW��.5��y�s�ż�_ڮ.�m��0��c�˺�{	GD#�G�����X:�2�<C�K���m�wU���fC�7y�={!�@�|(g<��A�Ac{�*�4Q����_T�4y�M_�o^*���c8��Wekʄ�s����K�]�e`%\��kRf�6��e6��p�smx��9�7��&'��$�U%y�������egVŒ�����مѮj�C���=��Y�p���u��Yoh-v�L[�B��Y�x<:��]~�}������7�OE/T�XI��%�e�6��y��/	�x�~v���[��O��0��1n�I���d��R[vP�Pѯ��������������@�Q=��܌���������1��������eםv�X�#��6z/�s(�k��_w�˪�����s�}�p�EƼ5_d�:-���r����-��{Q��`�JCy�Z����o�(���;��]s+��5vd�����c��Ҝ�5O�
5� �ǟ#O����cs���d~�J��)����n�k$��r�*��� �N�W����7ޞ�X��f���r�TK�OG�'�.A�$��U=M kX�z���OR�[#��}4>��ʻ:>p���\���d'%��w*
Ǧ��9�MF����J������ńn�z<��GCw]��Y�����`�w������ˈ�9֢/]��;N��˚	�Hۍ4:���Ѭ?kP���n��;��boM��Yڝp�.��y�������;T=�7��1��P�����kQ������m&���>��^8(��RX�vE�oB=OeWH�H J�2�2��v�ޗ��5�J�^�l\�ŔyZ���䷔�T��4'ҊǛ�|�=�����&v��g�dU�-��A�����)o'R��f`��1#�6JR.�W���=����|�m{�L~R(l<�Q��._�J��]�=�}��s^}b<�NQ�oi�	�3=�����>~��Z�I����<�9}{9'~�uެ����g�q��RIے�*>�PN�7\��G���e�*=uz��Uv«n'����c��W�)���*�{�}̺�}�ҳR���ED�U^�ޥ͇�K�TRl���Lǁ���d�n������V��~�k�c��-z����^F�n�: �;�����8wi�mgç:DN��+s���u���u>��x"c��t����wh�>]:���і1.z�׊�k��[����e�m���-�+-)����\�fLeض��.ԛx��P��g�S�D5::��S��˫��&+�1o�#wB4�w�\o5�3��W�\����̅�p3�)����Sm�Y�n��-[�c>iφ�<϶o�޿y�^��6�?�23L6���ީ��]��OJ�����2�e������^9��RTc�qڅ_'�+%]�w.fӬ}���~�1��^��7�u�*u��䕁In��I�9fG6�˦j�S�r ��h����^:<��@�?3��N�q���Wl�CA��8�bu��w�:�q{Ld���s�{���|�3/5��������m��s�	�=dߔ�I�9�$�XN�nȲo���Rq��O_P�d2���&�6��߰��O�~>�q�bW������%qſ�嬜���~��������d����d*d�+��=d�sXx�8�[��W�$揲E���(q�i��݆�8�y������A_=���b(����oqn�~G��\*��m��:�m�C]�Ad��s�:ɴ��Rq'̨~�0�I�'���$�dެ��$��M?�:�2é'���?͵�~���x�o��61����������N0�Ou�@�4���>�z�P����>��u��P���'�6��T?N� |��'�_�N�|{�!����AY0~��h��p�	3���.d��W�8ɤ����M�S�$��o��N1@��'�u��/�����CF����I�?�a�N%Bw���{�&�k�}�9�%/�I?Lq?%�%�̔�b��^�"�Y�7���DI�fѓǳkF2%ڵ,�1#�>�u�"�ʮ�������^�+���k�-��X 1zڊ���� �_6�O\�\1�2�@�CCd;� 6�g0��˾��i�uf���n�t�2md|�ڳ�Iڰ�}�����|���xT�Rx��іC�u�I�,�$�+4�Rq	�kx��'Y5�rO��'R���X�:�2Χ���=��u���'6�y���w7�?V��>����k�g�$��<�+&���Rx���P����J�0�aS٪Ad�y��N��h��"��8ʚ��q'Xy��߾��\��y��ݹ�?Y'�:w0�&�XO��p�'|�����:�|������!�h|���!�,���'YLd�!���XM���:���]p��c�˓��o��J��?������:oy �q���î�N��9�:�o6���L�z�ɯ���8�q?f�J�i�Y>b����u���)���=t��_�۴?~[V?~�ѼZ^/����z��>d�V}��d��=>�H,�a���jo��i?2~���M��Ms����i��d�&�Kg���@}Ao�\����Қ��~����O��I�OS�VO&�o��q��yC�';����=I8�|��'���s 봟�x��p���Mw���}���bO�yZKu؃�9~�����
��
������I�k
I��OV�I�y��d��!���N$���u��g;�x����u�>�>���>�:�O�O�u�p��+�c��p���'�PY'�voXJ���봕��Y<�m'm��XN2|�jíI8���m�~d���a�I��/G�|o���\�_���Vo����������{���'�Y�y�	�=d�I�=9���a>N0��J���N u�~SG���'��Z�m}�w_����;{�W�?`$��/���_e��9�?0��w��<d�OP?w�
�����]�Hu�5;�<d�I���J�$���
ɷ�d�'̝�Y!�W���e��[�#�4������ �!�}�y��S뫒�?�m�Ǭ���s�5y�1Qy]M����n	Kb�E��{�����v�W'�ڑ�b�[���kO���&���p�#�����9�G �Z�,͌,=ܴL�܏﷗��33[�����i�'��C�s�!^��O~�2LJÜ�Xu���9ܚI���܅C����S��'�<�x�q&��$�����N�@������߹���Ow�5�_�{���ɦM���1�̜d:k�OϬ��m'۰>g��C�o:�1+9�Ad��u'R�ORq��?��=I���	�N~q��s������{����wvJ��z�vȰ���iXq�i�4��N�����O�8�ٯ���'���z�Xh���$��9�d�VC]��8��Vo���~�O��l�y.��m�J��UX>��_}��M{�$����v��M3YC�'��j~��0��&�:��=��&��'P}�	?!����SL��=�~����2��o{od�VC���������y�6ɶM��Bz����ֲx���XO���4e�d��O&�:Ì'��d<I�oܓ�:����������y�y��\����k~^�m'�w�a�i$�ӝÌ���w�u���>�����O�|�VJ����'�d��2�z�:�2�2OR��VAI=�D�߷t~��_������5�P�M �{킓�N%g}��N���0�4�u��ì�}a?�u�>v��~�:�=w��+'���|��Ĝf����N&�;����s�u����ߗY�������2O��<���>��u+G��d�Vh?s(C��'wd�a��a�N>����L�~}I����q��?L�IXm��w���mߗy���]�;���R�q'��RC�OSS)�'P�1&2M����8���y�Xu���~=�H,�C]��XLd�o���?2~��2I��~�~������q���o�����~ٞp��~N��d���O�T� ���!�N���0�I��6�I6�,:���A�̛d���w$N���s�l�d�&�/oNj����-fƛ�o~��K����f�Q��m� u�g�N����
�]DM9Wgi�S�M��[[}z��ǳuk�f\H_'\�K�9�w�'�:��5�і(��z�ŵ|Y�;�+A̜=���L׺�j�[;��n��ϯ�ZkZ*�4�܎�>�O��c�UV�}c�B��~�N�L�����d�Ms̒��6�!R|����M��'SP��6���m�0�f��:�H}/0=@�]�чS[�޷�u�y��{���\���<I;;���'�O~��I��'�?�܄�4��,Y'�sY%ABd�͡Y:��̠m�6���q���I�g1{������������:d�ćB���I����L'���2i����$�i��?���:��5�`)'��*T��+&Ҳ~�m�Y6��o��6߻���o���5���zɴ������~��&����:�:����I:�9��2m����a�? ���u�;���ONk	YXO9�}�z���{�����>�����%d�C)6��'_N2m=��i����C���'�6{�<�c*�N��$��c'RN�!P�OPY��T��<��D���Oܾas���߹�m�q'{�	YXNxw$Y8�@��N�|���?P�'&�i��L�C���Y4�o:�c*�'X�LO7�:���=��?����'{�˯�oןr��*d�*�!Xz���a�	��d���sG�"�����$����hi�����a�:���{5�@�4����u��
�y�ܛ)�,�<V�;��~���¿o�W���*S}��N2|��������=d�d��d����4n���ɤ�e�'穩���q��k���:É��s���s�k�u��ۮI�I��RM!��p�	�5ϲu'Y�'�6���ON� �&�5�g̓��=����O�:���'��M&��2OYSӿt��}�m���_=5�w_sw���'y�>M2q����u'_��8��6s�:�d����2u'YC���N�|���s���>N~�+'�Rz�Ld�h�^�Y���߰;��Za��q[}�a�o�xh'�n���E/۸&�-�+̎T���� �7���D�5��T���
��Wn Jʙh�ѩ:�\n'o�s�\x;[�b.�_1-;Ԓ�p|��8�����n�iiخ��.�2*r&j0&�m�t��(�}��_��eRM�����I�ό�q�~�>C��J��a6ì7��x�m�f�'Y7��i�N�|���d�d���`�~�~-��˔}��5�������W�=ed�Ь����egM�Sz��
I��d�T����T�d�T��d'u���v�:���ì���}�K�w�ϯ�7�O߼}������5�}.I��k	Rm ��+'�8��Xa�N3F\d�!�זAa6�vI�V��!Ru�����rAd�����̠�(-S�jZ����zW����G�	�+�6��N��RO_�5>��!Y&٣�d�����|��H|�Rq��'�8�<��x�6�ȯq����q�׸��<��޹J��v��^}c��P q��|퓌�2~5��l��~�qa8�2k���$�4s̒�a0�8�d�����2u5��m�������Ja���G��-��oҩ����������������d���s |�xk�|�'�O?���'�'���O9�%a8�9�IPP���+'R�}r���=���_�WW�{���m'6�0�O�|�&�m�����d6�Ϭ���:�?;a��a�O�&���^����uܓ��O�x�v�u��;��q����xg3n��u}����~�T'$�=eIܠu'Y9�5��'���C�d�O�d6��2u��N��<a��4ì�����l=@�l�O=Af��ٿ}�<�=w�vj�Lٜ� �<G߂[ ���G�7���I3봕&�Y*N�|�����	�����}d�'~w�+�M!��q������u$��oϗ�^�o����m�gw���?1Ht��
�̞��\��2h��u�5d�XN��Ȳo����N2|����l�CT<$�&�~��|β~Cߵ�x[��\���D��(��ׂ1��KlKb��[������pYs�4�Y�@"{��B�ugz;i��R�t��Kݸ�a�k9Y���ià�c�q���ЙRv���:,V;lQ���C4r�5tK���o
������
o��B�L�,9��x��~�ֹ�>�ϙ&%a��p�O�LM�d�]�B��OR���0�I�'�5����5��%2Nh>�N��<�d�&�x��C㟹�o߼z<﮽sc�����s���=I�N���'P�}��	�No��LO'=ì�A`w�?$�OYP���'��{�|�u�[��W�$��E'��N���~Ϻ���0z�;�������}^��4}����a<��=f�:�i=����'_�I?!�9�:��z�y�d�T'}��M����܁�'̚>�|�u_k��������{����}��2m��ve����IXm��:Ϗ�4��O5�>f�8����!�N����~C�o�u<d�����u��P����}�%��sM~3�z�!Ozw1揄���\r_��`h��֤�i�,���&����Ԭ�����o<d�&���>C��J���`N$�9�N��'���Z8&Q�_�MZ��;�<��>l_���������6�����쓬��Fy�VM06�mI�8�L�=O:��8�m�OP�$�>0:��OۤRq'R�� G��bv����v�۞?���_p�����:���ì�}a?�Ì�I�O{��$�I��f�J�l���̬�0��!�x���S'�u4yC�,#���Z����`*���~�~���Q:}�IĝeM~�H,�a���i'Xr��x��'>�O_�5�y'N'�5�T�Hyh|����K`|�o�u��{-��q���O�����m�;��ya��qѿ08�Ԭ{�P:�ߨz}ܐY:��]�o�&$�l���&�ᐛg̟sY
�6��%I�B��L��v��j�����g���HVN ��>C�O�FI��M0�c$��ߘd��!�^`z��N�C��r�'���;d���'�\�:�'�?��$�i�y�7�c��("^��4}��
z\�6k5�owa[����a�7�x��bJ�`�x]���m	io�"Lw�T��>+U�B�X�%7Ҹ5�H\xI��>�c�ʳ��ڍ˶}��KG[�F����S����⣊{�s:��gq�<R�'���gA����UeZ�پk�p�_�V���a*
&��
���:�l�
I��O5a�d�f�P�'_Y����I�=�d�'�&�;�x�����~�~��v����߳{�����}�8Ͳ~a��{��M2s�$��5��(L>�IY:�����q&�F��'���RN3��a_�:��a�I��/�ߩ�w��wY�u�۾g�o��|og��0�9N2x��ܤ�<d��;�p'P��S��Y'��J�����aY6����N u�~S^XO��O�?V>��U;��*��/����Ͽ~߻�^�WĜa�}��&3l4w�~a�I��p�=@�l*���N�$:�̚��u&�~�*T�>�aY6�@��d���Su߽�{�o������k^~��{!�	���̚d������M0����I�Xy9�:ì&&�ܚI����!P�'�,�y�*ORy�d�$�MM��/�$��{�����ko?m���ݛ׺��ϺE���+'?$���2|�w_�~}d�É=�o m�d���βLJ��}�PY&;�I��{g�d�+?$�n{~����{�[���;�~k�l'�N��I_�&�rȰ�����Xq�~}O�<d�!��:ɤ�a���^O��������$�Jo����(���u�h�q��ڽ[���]���߹���~�~a�OR���� |ɣ�}�l���I_�'S[���Ri��P�	�:�?Xi�O5�>M2u'R{��M��N���i�˽��s�<��s=�r����ow:b~d�!��p�'����'��=7܁�M�kz��OX=����2q5��4�e�d��OXu�Wʭ׾�+�*����kg���{��?^�\�5�y�~ۮ���|��w^Bq'P�;�f�OP��a�N}a;�:��O�RwV�������%d�Ԟ��q
�~f2u>2�2OR�I��;3��w�_�i���E�L�89(Gڵ��OA]ufV҃/n֍�ZjG����CÁ6t]t�=kv�Tmq9o�k8�]#\�-Xk�ѮZ�Ħ
x	{3���:7L�R�.���W��=EХ.��ݷgP3E`X�U�pM=0t%!Ws+޲p}E�la!9S����;��R{yh+�7�e(L]WϷ�19Ow=뛛��m'�Rv�v�q2�����i�'f�u���ӫ�:���N�4E[���h�י�g�0c �Ƥ���Tyg1z66����;����;pGyZ�])e^#��-[�����6-�O������eSѮ����%]Gڎ qR�;�@��ӱ2��{8��N"�Z �ͻe��ՍPn����VQԊ{ی�*��d�f������}�>)�K'pը��^>#�_)��[�B&�5�iYr�=�Z�kBw�v�����:�+k�.5*q��q��R女�0eb$v�֪
&�w�EY���FLc`G5�n�{���&��:yy(��=��������Jˣh��-�ϒ�/�D���-������=ٽo���%v�	�6c����ƻ-��Tav��.�k����W���ϙ�&�V��o,���tS��������T9�XGl���
�'��� Ul�0���5RJoI�"s�'�v�u���	�e�6�J����2�|��r��>݂!Ǔ�����!�wX�un�Y��ާ.l�$�Q�u�)*wݽ/t<��V廚S�dj��*��ͺ�^����0�t.SB�m�MLν�۪��IR١��#Cv���]�!j��u��]��xd�.D��owx��W�.]��=Ik� ��ʣ`��bWwo=
�T��VA2�ǯG�;�Fc��-��W=�*��Jv�lͬ��L�����כ寁�=ǰ����p�pWb0ⷥGB��ɷDj�'����_J���Ǩ���{(������I�6n�^�L9xtX%�Õ�����w��֥푕���t�\����̏�ڜ)WY]{�	Y��U���������s��VO�p���ΰ�VjQ<�Y��LUKz0���[j�	���k���Z��v������R��KJ�k��u�Ӊ�qa�ୀ��8��!��Y9��*|�jg�b�Wۦ�x�u�~f���1(x�mL�IitwS�7+��x�_oM���=ɀ�9�,��_r�� ���_a���z��^��9�%�]FcI��=���"������n��,su�յL��v�b�,�=&�R��}�#����B;{PtތW�[kIj�;f矱ubs�m��������O�
��gs���"]���q�a.��7@϶kJ�̊�'ܴm�W��bj�W%.��/�㭽�mg_b�q��D,q(1dh�}�
����U�m���s]��v\�������k���5.Z�N��٫�̀aN��\UN2�'gW]��q��^K�wݶ�l��y�8�W�]H"G�~$�$F�ѫTj�m���Z�[E��DF-iD���)QcJ,�*������ԉj��
5(T���Ԩ"�ʖ"��EJ5W�\Z��X�ԴAmK,e�UV����Z�VUh��ʕQ�Q�iU�Q��lPh�e��6�m�Z6Ѭ+�
��JU*�J�[E-JYmj�JDl�V�m�iJ4U��V��h%�"-�ڈ������X�6�jZ6�ZTJ�Q-k)m%E��[J�V�%kV5*����ikV�J���fGZ�m+b�R���)m-����X�V�X"��[kaX�jS��֊�,UV[*V6�imF���ֈ�+E(�ƥkTKe�cYDYh�KT����-*�(�D�EU�1`�+5*��elET�ҫi\��U�(�-(�[V�YF��F�m��F��"1��3
*�R��%��h�ĵ��k*����Z�B����C�;���ry,`1��������ngU�pAkv`Q��o�h	1�+���9���{���^Q]͸9n��  xe�[������#�Q im�~�AI�N%f���N���0�4�u��y�Y6��~��u�>v��{�d�?��IY?0<���x����\�ƻ�{�+������쇬�'��&���<���<�:�ĬO��,8�Ĭ��a�x�N��:��3�q����L�~}I����q��/�~�Ͻ�=��}���7߾�o|��k���Vd:Z�d�M�YHu:��LI>C��yC��$۬�C��J�׼�,:���=�Y:��w'~��ɭ� ��~��������Y?Au��l5��^"�y��{��z9�[*J+4?A=�[E�q��ދ{��N4�e�T�+�߹�5�ԦtƑ�c�{| �B2g�� ������ޑ�zo�T�M
?o=G�
s7�s�/Ե#�I����JﮋW��ײE��"_TT�M�p�_i�(BE�/U��k�|��d��ޭ�ĳ[��;���c$�BP�����f���T�؟�Iw���nt�:��J\��_8�}Byԃ��[��[��f﷫m��[��\kۨͩ~�6�����;e�͈�� Y~���/ɰ�Y����EI"u0�x�0�%R����`���b���k_{#p�.'�(����ꎖ�����q^�U�v&{���>-�|]�9
�ʓ�Թ��?��yl�ǆ��q�D2���E���6����A��!�!�}����1�������}�W�g��b�7'+�Q����5��'��qq�����맘�:����:� 
�ڎ��ۑ��Ib{�Ԟ�6'Z�^�9�9��>��"�u�p;t���g��}��:�����J��0�gn���S_���zrq�Еc�Ѡ�Sg�h�螩W��\���_��$����B�+u�=wvs/9ُw�=�w���'F��MҪ���qS�N���$ܰ}2�z�w&��M����(/8{O�t~�
�a}m�gB���p߫ݞw촴��m�7�:�T�:�k��j�ثҹsci�+��Y7���yf��L��M�,E7� �h,�#�8s�G>�OpOn��k}��ϳ����HSBL��{ ��o;��v$�K;_s!��h��3�x{�(�<̻{|��s��F��D�<���8k{��鏶��#��d!�oP�3Vky猙����ňR���74p��ӣXM�uc���V��p�u&vU��d�S%f�h=��U\;t����&�R�B����X�͈%���oef��'W۷f�mn�����<Fr���Q�r�
��өd�Ir3�~�ꯪ������\�8~+9|k��2��m�r��V�����¤�nG���7g�b�4�e<Ώ�s�B�F��x�\�|6]9�����vE��ϼn	��nM�τy]X^SUڀ^�
��'T�Gz�`��^�߳F�ש�2��ᓋ{��Vþ$ʔ�u���g�=B�֍�
)���[�/r޽��rt#��H�q:_HQ��5�Ž���y�=�� 鷻]~�O�;�'���8*}(��N�-�ڌg�d��=-�{,ۃ;u��f>�j�Ujy^.��S�בS�Z�1.��M۷Fi��O��������;�\�e���%�yZ~Y�J�yo��qm���]�Y��.X���;Aq��P�Kݭ%c��/����W�.�p_ڜ<�㕦�IW�S�c�t�=�&�s�`�r��c�z�ߍBwc�x���x�b�=ý�g!C{���i+�
��%��0��N�k5�
l��1��[���e	������n�
kc]BLJ���q�g,+ ��j�dp�:�RW�K�1I�x�� �P�|4IK�e���t��_W�U��}g)��i`�M�U=:]S1�����y6��Z9��V�fB-���,n�]w-tgivo	��
�O}]'F'=u��V�n��2���7��	P{G��n��@2-Y���r{FA¦�ٛW�=�:��r��8 �#�d���r��BH�s��r�G��������s��C�3z.os;�E��u����T�(�A��ϑ�������m;w�\�:F�쀾�M�ݱ�~��w��NK���u�<y�OT+�e�;���QX�F�,ȸ��6J��"ڿI����h����E����u�}O�ZS��*�E���Iq�P�yH=���I���h�c�\g5+����R?f��g���c��T�������t�)}�5�=�p�f��I��-�z�p8Q��iռܛ���v@��'
�݇K�|��d�a�|lc�[�i*�mV}-�H�,������Z�NtM�!�Ps������ Lw["�Ta�۫+��]��~T��;�PC��P�N�{��9�k�r���%7cRf����F��Ǳ�B��ڵ�hʕ�B�q��z�W�W�}_qY닻g����ӐS6��V��+Ǖk{���Ut�
8լv���[���w{�	}ū�Ib�R6zj�y��]�L[�W�7v����=��h���2x�I"۩��S1��N����]�%P]��ND���8%zz��{���Vkr��N'��{u6Nس3e�Was6����}�����]c�˛�=�a�=��w�҇9R�M��$��/&���j�Gr���ȷ�s}#���Dƾ�m82���t��3]d��}Pz'KB[x���S���Qz�-�������=ǛI����I�-��M�L��݋n�	�r�K;\γ�>�<ޠ��}�w��OCء~*˻O���Vƹ�r{��{�_��Fu��yQ�~]�Z��s�(�Ǡ�}�ރ�9C=��&W�7��I��׃�s�!�t�Y���1z�5��~�<��4Y�t��;�(���j�e�pf+<���g	+{��oK�&�t�����B���^��A
1�V��{Ђ$�=���u�靬ྜv��1�GD��87�u�b�I���*���O@�B��Z�$T�'~������(����~�i����u�߯͡��W���$�zR�(��s���&NzVw/pz�ۃ�S��c���,z���-J�f=���{�Q(�`����c["�r� �c��}��yK�Ws�+��ި�&�hx��&v��I��j_�d��-��~�:�����Z{lޛ��`Sb�vfP���t��xF3��^��ok|yZ�&�"yBe�T����{V7'x�_@�t�tЧJ>y8*�1躌g�d�μH����N�Tݼ���+�m��v{�[��֫��J��0�gn��'r�����:�w����L�mO�A��jux�J�9�?E�#d��N�w�wgo)_��:�{������)��pA��*�5�z�O�>���u��{���z�ei����^��y�������]������%/��}���.��i�X�V�f���V��[1���N� ]��e7F$.�v�
B>��fV�>��:�n�L@�3��)���'+�d��aY>Žq�����O����󭵜W	d̎_w;+(��i�j3&,���U}U�_����{��:%��ߤ��`ѭ�f}�]�\ؓMK����h��=c�fJn��g39�Ul������w�h���cD�8�{�V��������=�'��a}�$��eO)��j8}��)���ˡ�N�M���ޏN0���ƻ��'��g���'�7�8w�b�>����ֈ���:�c�����?��h�5���}6×��f����[�={�p���e{{{c�5O�
5�8{�ϼ���z�ds��Q��32�ޖ'b�s ������{_����#� �����o���9y��s�,�]ۏ�8z9{.�� �$�Qz*v�T9��J�iU��Gٚ<=\0D���x����G}�2�o� xc<ן ���=E��Z��J�9�ۍߠ����+{S�������u/����f{!�4&��F��E�+���X�$�ˌ��׷�M�y>�bX�:��Yռ7��>�W�W�����|���yLr�k<���O.�v�s}�iћכ{#�پ{�������[�
����|�W�M�;�z�p1�������oj�3�C��2�����UU}D�y�������s�x�5y����uu�"}+W�c
fv����K��h��K��]�[^wF�*��_�R�N�ٲU�j��E��6��s�w2����T}۹T�uS[�0y���)G���J�5�V�j��z����5�mɮ�;��\�ۛ'nT�����<��E��'K���}Ʋ��,��]���5Sv��s����g���/�yqU�}��V��.2�d�r�7�BԚ��y��S���R�6�N��3�f��U���W���kv��v��OB�R��2�uw��L�RR��Ut޻�]�������)Zɹ�;7��p��;�o0+^ֹ�}/FL�ͧ����B�"̯g��o-��O�īe���6�T9���l�<���6� =��E>�֙+ң�{��[�9*j���A|���&�1e3KiB3��Y~�)�ʘ��c�٘%�֯%���>�=\�.I�ZH�l�7�[���D�5��-Y�f�ooUe�(��j:2�F�{���sƊ&�.�f��0�hWK|���T<إ�� ���c�Ou��PE���V|�����������^�̍A��;�ي��J���k�����u���M~�z�,Cn\j�wt݂�U�Vl.E	� �T�6/E�/&֣fׅ���5�H�������ʽƗ�K�z"Y��}�O'�R�����f�q��Z���w$w�%�ꃭ��߭��]��7�s��eO{�wz�+���RvZj>ؔ7�󵔷&�6y֯1��ZW�]<�՝<�'O0զA����IQ���Lz#��[1��K��_�.� ������+V�nNb�uH�*r-�{��K�_OI�Zԯ;C��P�n�̤(9������=�)�y�f�O�N*~�/���s$���̱,��+�~�sБr��k\�33�'r�p�k�Q��������I��x�F\{�m�{�a�3�������i���6-�ޓ���yD{]���.^깋�O6�9�ߗ�N��u���ʛ3��YN�-�ʽ�X�7����Y�kd��p)�-�c�ז�0$3��.�N^nص���i���i�Mt��ŏ�wrt
�#��sǻC7
��T뇮�iL���+�z\��� ��<�r&����6����Z=�־�Or<���'��y�1��@\x�J�[{��2ou�d���F�N�Ȩ�j��hk���2��Qz�[=�ۜҮ�6S��o?Z��둥[,r��G������w�������ef����;?|�y�g3��~�#�]R��T��B���n-y��"K��ۍwl��El�M�VŮ�W�C�˒-����;��{+=���0�v��%���pb��_f�,)S�[x$~uB8l̼>n����9V��@o�g����dw�9,�=�9q�x�ǆ�y��$�A0��|�P`=����yIZy�����*m�2��Ww��'H�C�����5���_��[WN}�<��Ð5���7�ٝ�/�C�Gj�N_I�E�c=�,��_�U� ݨ`f�vNy��f6�e�V=^�,�8��sf9]�O]l�.&�WR{]P�{����V��[�d
��i�+��~��ol�l�� t4U�SZ��nk�ǻ�e��W4�,j�/���Ѧ���՜����A9��"��ヴEb}.�8m^Zh�
��q�o��\ݷ��d�ؙ.	*�G-�3,N��0r��4;[������a������Μ�+�[� ���ޙ�Z˹��D)kY퓫8E�t]����Eiτ��k���0��7{]���i���,�Ha��n�meZ��n�Y%t��TRN��뛦H{d7�Xf�H����.ER�9u�ח��uB�r_,�A�W.�iL�v�&�q���r�q�ᒶ���]�<"�ƷA�Ʊ+{�ڵ�l�%N`*A�2�w&�]~��h^�b��˷�����
�g:%,�F����o�	��0\`�dz�`,�W4B�\���e�c6�
kZ*��ҲV��jC�9\�;$�A*��9�ի�h��[ZB�)]w�ݰ�v�V���2ZI,�l�m�N�F*7��*�Xs����\��:���v��k�/��}[�O-�<|P3�����t�g��ސv\wƹ���tZ��Q�<��MD�w@�cn�,5ٽ:�r���p���}E#z�4�c� ��qcEuwdnCMLS|�ul����7�8�jCZ�;v�Vm����:ث���'��I�ءR��Y�A�L=���p���BJ/e$mБ����t�����A��#FT�uk���j��7�'N��%]>Η�L��u	)��5�M+�*k6���%�8I�	��i	d���y]�@�Fr�.�]d��z�ufn��b�#��r96�~ 
�WT��j���Mw0U�d7:�7O�ڹ�D��I��qj�����9vm�й;����.�Л�}W��PV�:�IA۠�l�%�u��f㸋��"�[��1FQì��@ŕ���q����:U����ǻ9�Y�eug}#�+"5q;K�%ܻ�ٯ��X�T{�z�A�v�=��$���v����w}8�v�y�c5ۘ!�mX��.:L�����Db.���j�����5G�ڬiwX�f<1��k}*�Zqp{-
�^���e;6r�a�ӲF;m�O�ku1. �B H�7[F���s��C����÷M���j���Uo:R<Uj�H;�99г��,�t��s�������S�n�xu��yP'��7�u�-;]���k71DG�ͥ;J���ݽ3C���фP��cu*��R@�T:ZZ�ּ�P�����V�9��L�k���hV}y���ٛ�ͭk]�D�2�}�[�n^tq�:��ъoP�ML/�m��;�m����ÓF�����`�T�5]p��֘o���i�.^�}k��.^�˾�u����-�p��3�ʊ�PQ����a��S�R�X9���W7�������Z�Z�1X��Z�h��R�����J�ň[UTb(�EU+(�kQ*��b"�ҍ�J-(�������5�F�+W�YZV�V�b*(�Z�DQEEDX)�QAL���Z
ZQ�(�k�Z�"*,jU3��6���Q��B�KZU����*U�K(���ZP���RTF�[E�
-F�mF[UjPV*����Զ�(�2��ZZ�YQ�Z�Db��(�b%��K)-�l�PZ�eQ�"#�QAE`��,H���DV,U�Ub�,�J���`�����KeQb-�cR�`֑��JؤUX2ҢPQJ�U"��X�*�JF*)X�8�\VATm����"ʬPm*1Ec-+kE�խ���F��ZUB�ԭ�V"�h�VV�+[kZ6*#"5�Ҡ��������Q+R�*�UF�bֈ��"QF1Ab������aV&0�Q���R]Z^�ۮ�B������u&�ֳ*+�ۂЩ��mj��]{�x:��Q�ͬB
W#Tx(h�ulA���)�w�U}��}[����|���L��Nʥ�t�Β�i�a}S3���uV��V�x��wމ>������>�n�3ԛ]�u�b�*�T�WH���_L�w�^�B�H���nN�5y�&�Z�*3���{j:]�ອN*~�R�sP��1.Ş�Y#��ȓ��^���~{�R�0v��uA�]��F\zv�yE��"�sǯ��~;�����]d�R[�ëF>%����:�u�=[5R}fK9�@�/6�_�48�T��&˦g>͕��v���[�Yo��`�W��ds�ȹ'1�d��k��:�̕"�ʧ7�ꤧ��9? ڿf6�?A�x�s1��� ��i=�T�ٙLt&�I����z7��Gŏ,�Ech�������
=�i��]˦0֪=-}�%�>�w0�Ko}��I9gm�+͌c��!i��͠�(����s�wK�����k�	=��'����X9(��$4<0�/pd�J�*��+,��ɲ��tm�3E�-�0x��Y팶G^5�-��˜̔�]j:���x�M�������)�R�����u�t���'�g0Ke&:��B�>���Lb.��� ���O�{B�~&z��+�'�JY+�i��������t�v=��(���]���D'&��R\uکeI3hJs���S[���C����|��n�.V���lK5��n2�N���b���X��� �=~�Z�엱N��w������f�L�4v@��4P�݆q��w^�MEc54�o1�z�;N��^�T_�V�����u��S�^y8T#��}�Ax����ѷ�?���Æ�/��=����4���V�)�ܯD���m����*��/�ꦷك�Q��wy[��%:�^�R���^�n���߽���s���A2M�K�#4�K���-����
*������J}\�U�Fcq|�"�:�F��^M����k�!���n�.���s/ڱ�y������(��*��·S�t�-����W����m�V/zne�Ͼ)ǂ��s�h5�*���ċc}�V���hǞ3!5'
j#^��
6�z�U��([��Ē�U���x����د�=��]-��v�ju�ݟ��� ;���4؅�����TOz��V��V<�/]̱2SR֍�;���LU���}UU��J"���qx?�{�TN�gy��K��Q9�F�۱��yW�V|��zH,.�w��6�������]����36e�uDU���>��;1��zR������1�F��VU��=�:㞚|A�"yZ���|�	�a�s�S�=���5O�4+j���<��f�)	��9����b���9��W�Y$�-��4�X�2�����U\��6��y-�Y�Ѿ�n�/�y�w�캩��I5E3�k/��ZN,E�y��w>��Z9��^�M�=*�d{���:R�O�c��/]�Θ˞��#\��j�յ��˯F�b���7��P8��n�Mk��i�'� ��Wz�}�y��NyW�yȺ���ۧ��R�[k��%�;��"~������I(��>
���>�Z�~{��=�{*��aO[�ۦ���_��n��W�Q*���6�*�Τ�9uĘ�S��E����(e���l�V�^�U�|2<���+�/:RnT�PJa9˰m���KUC����G.�Ϣ{I�X�-�"hS�6��T�6K�(���1����w������� ����c�����ީW���&m=�)�۹'r�[��cTv%~�[wB�2%����̹�M���;6zWf�N�8��ˮq��&�Y��N�x �����9դ����wͽ(k�^|�m7]���~��q����v�T��;=}�m�����g)��ڠ��1���W1�;��������@zB娤[��:oR��C�}Cr;�UD�3�saԋ��κG���s�U�vM���Ѫ����SUl���w�e��'yW���p_-a��<����Ц��s�l���M��Sz�y�l���~�m_�ɗ�[���*{S]��s�����L������;��)���i��K���Ϲi�k^�o%uch1(��F�����6�;�կ��˒-����c~>�<�Ok���@��.w�ܫ����*�nY�;�=^�z�oe�!�#>ol:(�&`�_=�^�t�e�!��n��ϟ܄9o
���Cۇ�Mw|E���\f��
�}�wY8up��l^-|�$�������lu׫���i&z^�����o�*L<X��%[�86!͌Z��ˢR�X�떾����_}��_Y�-M��a��~�c��G�7�c�A����}j���ѭ�n� �7;{%��Ԗ��}����w�s}Cl��g����Zy*�ݩ��݆�\��]'DX�'
���}8���^��Y�{�y�C|E�X��6��ꕗ뵳�y9��S���������]F3Ջ"�a�o�S���7ۏn�p���u�pпe�����o��l��`��+r��Ņ�EkgL�%8���+e�v=U���zQ�[M<�U�K�D�r�N�ągOF{����׆<#�C$g�ric�lM � ��n�	u�N����>��+ˮ0��2>aY~�B;�d�-z���!}%Mן	�D�>��Z6�3���[B�c�9�*��ns��/�x�����ޭD�|9�7�������x;�x�Z^�a�b��բ����%�xtK�Q���p�J�cQK��a�1C�<�&@ǳ%���b_|&,9��x'ͪ��93��x��ǽ
��fj�@y�J���7W�Q$Ѡ��AJ���ۣ�w]ʔ� cჁ�sb�������G"LI7�ZŊ]s��q�ZM� �%��m��8)d�r.4�հ\f���qgG���ʺ�o~�ꪯ��U�6��r������xW*ԧuC�34�"W�7o�)S�XU�f� S7]�7�WdO�����C�}�,EVҸM�E����Ϸ�*�|{e��\���������>����j�/&G��4X�W�LUO�3�^�j����~�~0R��6Gr�ْ��Xj\�!6ưA{K�W�l[a�;__�0'�5�f	7�s���������)v%��,"D����\�'�I��@5�Jlv��c�>^�w����<���%�+d��T�yB$��<�՘ �-!���=C�F��#�m`wA�#��ڽ)=Uk��ɋ�ޗ^&B�r�к�ŝ��DhU-(<>Vuݧ�;{��q�q�x
��^�sP,̗��Wz�/z �J���]BCl�2���qRLXߟ���=P�h=�	f��ʥ������n��]j�O��|{����隰���q�{�
�9lv��Pͯ�\�5��N{iټ��9J�eCż��l����X�dڋ�5W���8V����Bly�^�ݙw�.��>aӷ��)k7�q{h��\���"&�<���}�*_^���] ��yٱ�n}Ī��]8em��$�G` ��.Ipr4���³������]:<˥�os�_UW�W��x����O���z4]M�Ob��+|�d��+�	��%�ϕZ�4�Pƺ�ٽ�j����{��{���M�{i�uM)gFS0=7U6(+rZc*��L���R�<�r=Ѩʽ�v^f��x�7C�1�xήV�WT�o�r���q��'�B12�<�
T>�5�
������qg����I�m(�u�h^�{��s1W�MbX�+��5�����y���#��z){2�&����Xር=�*�sr$t�O+��[������x��="o:��<.�8<42Y���I԰r)�7���"ŵӆj��Ǘzpo�u�cɯl��1�u>��qC*�w�g����O��<K5Ka���֞4sr��6W)(����]��~c������b���YT�O�S�(�X�� �h���}�z>�����g�f�wM�W凷��c;�)W�;��+��r�8���,8k�,�W���z����]�8�v�.J7�K�>��C�g��CL:�,w��C��j���BjC�z��׽��x�K:�Ë��j���q7�b�)�&h�{Q��:�_4��.=�g� X�n��[Y��6�N�'{�p7�E��H6V�/n{��Ҵ�n�3G�z�Xm��ǒ�r����zFm�^��,�B�kt����Y��磌��s(�n-q]���~$�$u��
�U{�j�
t�l]o5�U3
�IЁ�{���^����7��ݝ�Ez�����{���G�}�yh��n�*qK��<�\3e2�Gf4I�kz�wy�ĸ1����y�&����t%��/!ס�1^�Q�eԟ���+��;q���b���˔x`��(x<��C���^���պ�-�J�xd��x3tй&��h�r�wF��p_Y�\����E��U��	��̞���트pᢳ�p!��.u1?wYSw�\����j/E����Bm�6�R���p�WZ�8_�T���/g��������J{��u�t���*�f��67^��W���uzB-� X�Ŀ����1=6�u���gg����z[<�R�
������Z�שu�����}�zBr{�z^໫)Iz۫J]�j�d>�c�dجk�ib�8o�k^}IA�U�4s<,wD?.ڄ����x�C�7`K����Wi�u���"ĈaQ��<N�k�Eo�'�.G����k�沴�e7Y��q��n/H��k�]�b�"軩���ovj���h�zi���>��'q��$v�u���ͮ7;�wkŕ�H]��|�-���2�'3�2ˁkopT���b�va�hf��십&+e��������o�UW�_}X�b:�W����ᕷ��/g��Ɇ�����m�����G��,�:5���PW;^�.9v��g��1<}K�Wy`\�SM*s��9s�U�Ժ�7N��n;}lp�ϳo=ۜ�g����9`a|�g�J:�^��A�x;2���i�-���2"��y$����(%�%.�k��������g���\65�ץ�Xڵ�9P��pw)�<l#�>������뤐`g���U�U�K�iL�I*�[�Tdt�Nn�%��
E�X<�7!}�����6G�%���� �j�nD3�t��]͡����l��]��	�w������BB�)��uQ�5<+�B5ʼ���;��5�;�U[�N�i���*�j����5u�*�m��^{&4�vF����vA�N�<���*&���1���0��۸&�|��/g�WI^�y���g�,�k2�c;��8�$pj�1+s��N�׋���W
��L����B3�QS�
�y�p��cݭƳ�J8�7!w�Yλ&X��3)/7޼hp3+'3P>����rΩqf�v�7uc���l.9�&��[�M��N��ùΰupΙ.����v]�d��R�uaѾ@,��Ё6�cx�5�V&��"���m[������}_}��GXT�0��~�F�d��V������+aKH�
�<�����#�y��x�.�G��͸�Ӑ}*]�����ISu��p庤l���Tש
Z�*cA��v��g-������C������!�S��K����~�|��I���#��Zf6̱�!���:��y3r���S�%�0ɑfi���.f�Q��ٙ\�\7@�r�BCPD��t�/�X�L$���Fc{�a��S�3�Q�Fj�~�%��D͝�I��W���t{ͣ �h�V�������������g�?���o8U��~����o���fu��мd5�
yM#CG�)R��Qq>u��V	G�C�j��hs\Ѵ,K�/\��0SB	��4e�w�g�*��5�����ض��-Ġ��:��OW���sL{��R�r�y�cl󜰉�:*T9b],���A^=X���:H�!ƹ�>Wy�վ[�}���W�(3��8F�萾8/�9)�YH��X,R���2���j�o1J�)p���|Ol�A���������Ҋ�=�|H�R�s[�)����Rj�2<���YF�=��;*�.Ji���� ��^˫Z��n�љ�sT�g_ڌ��|�q�T�GYj1ou����}}�wV��$Ė��Q��.]nڛ��u7�d��o=�M�1e�������/M��ne�ռR���=*��e���T.(]�R��:Ӹ̋t��|��D��}SUtf>�3p` P���D�ZT�mQ&Y|o��xi�+@�wh��+����B�dq��Wm�\�e��Ќ�`*w�E����w	U1A[u�4��,��$h���8#�Uf�:u��t��f��٨X8��w�F�����/Bl��vv�ū"W��S�S`\�ެΛ*i��S��ne�9�A]0vM��G/�EǒQkUKbL�Ӗ��q!�.�ݶN�<���бN=�Y妇˝��A�-xn\�.
�8���Ю;�r}�(��ls39���i�h˺��}�RcBN����[F��W^==���&dz���Oh�Nq��j�\���gv��oiK:�ͩև^��b��;x�7�T�]�����(ؚt�����V�1	l�
�Y�w��7�����2��W7-¶;Y}��ެ�:oU����CO1��Wrg5xRt��sF��W�Gׯ{�=y
��*�ư_'Gp��t
�ɽ�M�UH&�q�.wc��S��=�|�G����1).׻��q;$����.[�����l�P�|\ZemDU����o�FW�a����<��b��CB���뮰�,}���;���.��ˋ%�����%\�f���g�x,��WRSN��Ru��u�xN�r4�[�1U�\4�����F�R�{G��o��2�y���)h�h�[���esI5yt�����,#����D��!C�4b��)��=O���0�̘L���R�L$�k'�Jot��������c®ֹh�xA��}����n]�ڷ��tu�۝�_G}f�� 6�]U3�}���c�s�d����V��'�9ª���5vd��[y�!e0�����z=�@�o��t��h�2t����Zj�"#�
�3Dт���Ö�:�$�5λ��G�c��st�y��>7�<��&6�HE]/T��������9+u��#9u^�+@$�ۡ�8$���fãU��c��@w��J���ҡ�e4No]���#tm?$h�s��@�}�$�؍�}����]��x=�����u����ٕ�o,���0�r�"t��N6�p�L�%��ܮ}l ��ݫ�f���$0��˾��W�C��Ռ����P�/]=G��]oG�D"�U��[u�{�.7�Zm�/m�=�t+Rp��R�uY��>{���Q��#ۨ���׷��qNP�C@ޗiK=z����4�6�1*n�x���U��`��V-EIX�c|�����Ak*���%iQmicR��J�ZTK
(,TE�F+X�D�[TQ����VҊEDFV����jU�6�TX��S��QA�,R��Rڭ�QP[e�2�صm*�d��V�`Ķ�(�"Ķ��щ[�UU�V+l�J\l���j�F1Qb�kADJՊ��b��AYZ�1 �ʔF"*��j#l�F�kEADF"�QF1A�Z���"����U�QjTQ-�V"�փ�h5����U�����X��Pe���Qm�
�UX��R�AV#QJѴ�EdJ�X�AU���"�iQJ�UUJ�UU� ��* �(�m��(,b#��V(V��TG)Z��Tr��EkV�U1XTUX����(�*��R���b�T�A2�JʱV1Q�)JUUQ�T`�J%5*��E��AU�
��KX�j*�#Z��B�-1�*��_/����������^�k�l�s3e�V�1A�)l9{eV��Ũ�ӡ])�'��ȩ�Z)��̌���#��n�]�U�}��i�ے�&C;��Ō�֎�Z�a�����ҡ�T:]�7#\�����n�P����Ȫ�'׃sy��<חX��e�kQ��i�ˊ��Y�ވҽ^�qWP�Mȩ���;�<���i�}�G����>�Z��48Ӳ�Zq�ǆT�s��c�����v4x\N��]�퍶L���+g�p�#�V6���h�Z>j��Ǣ�
��(p�`֥wWdU�6�9�w�߼tA.�e�4p�d�F�1�+�lz6��֋�A���V}�`΃V,����bӷ��X���t.����y��Җtc0=76(+b�]��=�Wh�ΙNǪ0͒/�6��n�y����z�Ѯ���Y���8SQA}���7�Єz�xn������e�����tI�Yw�hP߽��@.0���o�BMbo)\v:'����u�������]����u��çȭ)��ҹ)	��T�u��A��/�/z0��F<s��,;����γCJ#�KR�h%�����}K�8�W훬6��0�\�Qަ�O��ݢg������c3��ֵ�u��j߈z/�f�%9z�����"�zr=��8G��.6}�}������|��e�M|�7ۮ�[��o���͕��TΝwt䫰�>���,QZc��p���y�߃����v�8��r4������U\��PϮs��
��hW�p���w���^���b���j�d~\<&NOHy�1�1V�s��u)�뉋���� @� ў�O|s#^�lI��W؃�W��_+Շ���c;�U�gjOK;��0t��m�!ݠ�=|�b�ݳpY��g���Lg��r�qWc��J�;L�6�R�UڜW���f"�ԫ���� �`�@�
�5�G��wU��6/��J�� f�cQ]��dq�|�I�"����8S��m�8m3k�E��u���*��}�y5���`�\�/yڻ�g�,�*I,�)�l�!`��E���T��pӿ���Η�K��i�G<h�N�7��{��{γ�O�fa�UO���{�p�zL�?��u�+l[��Z���e�!���Zwa&��G��y3J���i�]:�U��|$:ؙ77S�QW4S�vߎ��C�gA�Ȼ�<kv����r{�߽������{�*�*p�SR�8Xu2(;I�Q��o�m=����j��v"JH��oa
��A���3a��W\}OB�hV#7mn�<um���-�ó��u`(RHa:֬}� �����6_)��>����6�#g:�7�Ϊ��;�[�8�f��FTg*��I��着��ЩEr?OB4�7�F�}H!�����
�����]=U �~b]5��8��	�/	��=&�Ŗق����s�Kʈ��z���([�_�e�H�z=!8މ3�F]X����.*�ɬ�}��O��c W�%-%���0���kh4�u�U����l^L�z.ل��6��D��17b:��E*����`�W�ԏF�������X�Ȼ���n����qWA}�v����4׏��L5����o������Z]D<��؏<���^�c7��YdP���ƓS|���/���i�9��g��g�����65V��[�<���}�֥_7�r@�a�cq�x�u���U���(��|u���&Z���ϵey�a���H�7�<��r����� �XM���x��rkW���웚\١�.���I�)UE^�׉5�_�EiA�=zi�dvR� q�--��ݑ6���Ҍ���،__��8��d�����Y�.X.��ނ.�rŪ��&(�?L��PB�z�#
�=-���[��wbbcxb�o����A����Y�D3�h���LN�HBU�c���/U���܍廒q�p:�A]��� r���&�먾����ٛ�.��.�����n����w �t�'U}U�$�/`'}=���qzXT�K��m`�ϯ/L���$/�+�H�eX�!�57���*�y����[��F�}��
�+���k�a1��^Oe�t&4ƈ�l Y^0qa��'yڷ�Yc�
�i����~a}y�pM�HJ��)WIJ��L�ȇR�װ��o�a���C��uY-�k�J��-��0y����Z�	u֪x�5[c�u��ݮ����ҧ&IY���{�Ķ��yy*�!�"�UB�`p�5�����y���]�q�1zoI���b�z�\�N�o��M�G�Qg�z���b�)s����3/<�)v�H�m
�Z�&/�zo�T�M)�~��_�=�w$ۃ��h�����	w�.�q��׫ٹ&���h�(�e����C/"L�0]|�3Y�1��v4�A�i���Z���ξ�Wib3�譶%��>�b���W9Ʒ��W�Ƌ�f�����^���XB��Qcq��(��@����?�6:su�ht]�Z<0?����nC}튻y�xw�/ޑ���Vv��X�`t�)��y�_ru�{�@�9�8s��${�b�1I�N���4IW���{Ͻ0�~��`]G�`��$Ȼh����]I�'�Ү;�ڹ�ģ�mX�~]Yάn��wo7��Y�̻
�M��Z��=�`7���_}�,!v�vH�?6����rh�@�=�Ai�e��0���"�2c�1X��LC��ظ�f�M�,�Z%	��4e\�|���Vh��8�TJ��[a��oݶ�.�U+��Iy��ô�'�0���x;����i��n��Th�s֓�I����8.�͙�=˗�W�}�h�f���x8S5҄Iꐦ|7ࡇ*]Q��|���p����6K���H�)�B�F��cn�-��JD���[�h:�GM����;�Ř��Ӟ�6v����)k$Y`ör�Q@�3o��V��oE�Wϥ*�X�����:W���t��g�G�X�D�m���֍�J��Ɲ�c�r߬�Ϧ�F�o��e�D�R]�s���I,�1�$d��r�纯�,�/�<sM���e3�l��k~�mzw���l�5��o���%^ڂ]S�h���f���aT�K�fҴ�e�̞�m��)�C<1vjr��Lj����JƵ�2���^0r��X%B3�]a�Rʱ�]\�lb�:�J��g�Wy���3��p�.�4��=�
���}9��喕��x{	�W_�\Ie��')ֲ�&�^��^J'�2��vΝ��󂦜+0
�NT/n�g/tf�H�/;&v�ˍ�]��L�y{���;���w����C������kuߜ��A�߼��[|q*�1Z�h^��+|GEC��������3YK��K���]5��`�)2����)mᨒZf}R�u��M^�{��s1P2k73�v����O�������!�ק?T��x�T7K��q�:N�x�2�H;�����jYG����a鹋$I�\]�W��V�9�́�j��ƇZdia.K'"�^>�,��\��]�(5z��S�f|{S�U�\��P˜��04V�Du��
����'��v�T�U���}�*�;h�MM9Fj�X���s�AI�e;����A�ǀ���I���mU��ͧY92 ���c"�zX��Vb����c�C��+�C��.�t����,{7n-me<�`D.�t�|+Q��p�૯-�2b��r�س�:��q�����?^���q*��O���D�А��ޞ�^IpЅ��*��0f�D��i=���Em-��ܾ�y�t�2����<Hח4���I��h��^Z/.��qp�Zm�m:�1��RV�D����r\ՙ���7|��μ�*K��S<7q2��J˘B�泥�����s��
VG��[s�Ux6�]l6�T|rՓ��ի��3��b(-\9 �XZuFf�Fixl�nV���|�������7(Zy'w�ꪀ��|��OiҸ��t^UN����T�� ���2���B��X���m'/��bx��ɴ��7 =��s�WR�m��\:
��P�T�;"���n4E{*��-����z��S�3˥���i����~˱��V=��)��L�a��+�����ߢ�0�peɢ�q���_���)�oخۇ�����ZD�N���hp�tNє�ÿf�im�~k�p�Lz��ˈ�y� ��b�C�_2}Z��ei��)�/�<�ɦ�?Z��*�d-=9B	i��Vj���E6������_�u�.�#=ԗ{0��U�D��f���Io�)�����c�dد�-q���(,,q�5���*�����Z�٢<��{"~�����&w�,	sբf�Ӯ�i���D0�u�fe'���:�6���y���
�3��Ww�d��ɲ��}sz�7Q���	�6z���w���_�uߙ/�rr~���/Ő���F�pc���r��q��D�I�+E2�/mY�r�����u��w�<w�����8"��җ�/�{�Wy�D�;[2my�n��k?[��n�(��V+�Т0�[P�˻�����;O���}ӿ�xvr�Y�|�	����m)��@5n�s��8���w����ݓ��7����_U�ҽ��X��t�@���J�|g+.!���W���a�/�y���}�*B1�-A����׼��}h3b���Ku�@���<J��{�v����"��� m�q�K�Q�Bp�2�-h�"Ln}S��n��P��:�$qz��L���M�L�11�Rt�aV��Ӗ��8��Է~�L�R�=G\��!}�،C�l�k��&����r��n^T��E�/`{���Z����j~����e�t��I����}�V)e���Og��)p�8.^��㞽��/�`ϭ�ǒ߻`��vK�D���NOz�nn�+pg��}�Gyd!+������Y�g�0�u�)���3a�S٢��J�����ri��g6�;Ķ���b�YyP�����k���.>`\DjǼFcl�g޹�2�m�s�pl�![7̓S[���2����ŉTV֑T��&*�[��k5W�m�j�R�&.�gd��>j]���xi�اw�g���DXlC�x�5����ɪ7��vET���jѼ>w`��{����[�{��w��8+���N�������l�����bu�+9ًz_i8J۲x��$%mP��n��r�O(���jC��䑇xkz�'���v��\�i�S�YMS���J����g�����iu*�tO�Ⱥ���*�SۊP�����LEM)���������	�w�;�x��5�#�x�u�[����_%�c�������o(�{��+��a�5C��o!�1�^u�)e��v��U�ۓ7������ֵtȳ�{�%���w{̓���i�D*v��r���ѧ�����u�Do:��?ږ�<C$ue��u�,E�����T���^'7��s=Zh�reǈ̾�y	J���%<ٴ\4�U'�h-<L�9q���P�)]���y!Yy�IP��S�'�菉Bs��
D�.��� �#��#8������V�Η�����zϕ��b����O���W�*�"V4r��a�V"����'�d�F<����0ŷ���'n��1]%O���p��5��oK���!�Uv/H]0�[k��G��V�VIW�<`�-��[��3�}�:�Y�}+ĩ=�n���Ʈ�U�/�����t����F�F�%u�g�P6�������x����; sn%�K���R^y��A�E]�#����{C�]��zw5[L��؏��^Ȏ��Ԛ޸��¯�WD��b�o's�g+���8���$��,�����n�2˵�t��_P��44wM]���7vۅ	�� 9�خ�fAO���u`]�z{3*V?m:����{�1�S;��>��C�8P��9o�xr���Mʹ�ŷ={����|C5aʝ,'�	"����W�纬m�	�խ���Թ*�z�W)0e>/���~��z;�4��P�ƻ={n�?q~�{M�S�.a�g��6�et��4��(ѵmnc�ٌ��ڪj��R�Iп���*��LK��,��`znlPV��֍҉~�y����[��v`���Rۇ�p0��c���Y��#���w��=7�#MQ:6�G�S,in�Y����a|�6��>�U��l���f�x���.���=][�s킆j��[S	bY������$��$~��C�}�\��=v��~4��߀�']xA�Pc�N=,�ڙXK��i,�"��b�`����]��k8&�ONQz��͈��m�(e�w��V�Du��
�b��g�M�On������|�O�^����ZjiϨ�Pk�1V�Ns�C*�O
���<����6,!.��{v�Q�=�,�xQ��k6���
��/�r+Vo��][a��d�xl!Zu�䚄��A�r#g��0���/{j��u�[����MKN�#e��ބ�_�9��O�d�.8@�4�����q5}(�	}����k��ϸ��1���S��A���i#.�>N�bgj��l'u+eXd��Q�m���r�gp��o�עy��8DW,�tS/��_Ob�*�rF
�~u�����]X <}EQ��Pi_ZdolL�2��_)��j�#��i�����		�﷪�Y�ά�X����8�o�/r���x[G<��\u�����sm3F]I-L�2�ɶ_f7�Y%�+r)�2��n�H򻟏fC�~mV�1���>�������@��ms��k����sGZᱶ=�q�̩��s��#���.����#.��5"^xTCsj��\��'��Ix5* P���7��L(}�vK��.!��C���Ų�eK֬�m�Y�}��3�5�8v�Z�r�7�Ӵ�W�P�m�il�8Z�T�1>�yd�+�g(yt�I0� � ����L�
>���A���4&K}*�,��cu`�kP�e��,�.���Y,d[vr�gw�Iˇ�����M�T�1�j�A21�zgI�|km2�jhqVM��c�s�����u��k!�f��d�.��Zo��w�gy��+���`=�����Alrf�T�fĮJ���Ә��n�vn��2m�����ެ��OC����y}��n��Ԡ�n��^ⷦ*�إwT�˛e��6�䮑:�%�TL�W0*���<]3�*�0;��U���s�T���Lo���r1d=�}.���G�1$sg�VN�b�
�U��_c�ʺ�g�<�m%��&hsc�=�r�	^���U]�mh%���9f��͚��w_n���DW;��R�ұc.��Z�E>%w]Xf�2ە�oWLל��
;����$�{O�Y�I89����m��d�u^��$�G��K[��;\�y��
y�x�h�c��Ⱥ��w���gD�o�W�+�S�S$Y�L���:ngQ�y���c�Ui�ݽ�;y_em���2�#N���fΔ ����;�z�s^�J��MHX��v�}���؉���Xť�w�oz�h��?/�ˢ$봻(�UN�7֮�{�LU�k+��܉��`�S)�}Ư���WxLF�P���dnc6&|����SZ�y�^Wm���^w��w/��=���jGV�R�Wan2�w���	pձDa�r�G�r�bQ��7/kB6��Ķ�Jʳ4��������գ�n�����zFM��%o�*$7vS���>��{����c\����5(#�_]|��yƜ<��:�}}��C���i��>6�W,�����V,"��Fڱ������l�TQ[J����b#�V,KB�DX��,LJ�*�Z6�V(����UJ؍���[(Ȋ"�����b�"�VZTb��F"���[X�Zآ((0cR����F)SF,X��6()V�`�"�#Z�2T*��X��#�0�6�X�
�1Tb���EDEF	�(*(�1m��ԨT��,1+-L 1T���DrՋl��b*�U����FPE`�U�X�&5EQQfZ�� �eH���Uc(�J���+
(�JQW)Eb�QEPETDF,R,X��X���H��m� [jPDB#�����*�DX �#�Z�b����E�m�(�J�,���c1b�" ��eQ+TUE#UcS�������.Q����l����DX����UDYiUQe򺏨�����A�3��t����v羰��7�b��t�ޓ��*�GL�H�M���q�i�%��6�P�ʯ��x)nvĆ � �
�5�U�c�z��},gyJ�!� �+��r�T�~��ovҞ�M���3�s��fu�ƺ�E��*����C�<���L8]z\�`����yN�6�a+`��/�LZ%�	m$�Əy(���7�K>�g���>������U��΄��24K�4���VP��9��v"K��3
���3q*c�DO	�^"������9?m����,��^|�XO�} � FH���uv#��Ԭh{����NU�q���Ľ��6��v�4��U_[�����U>R��{�~
����t֭�\��W�(>l���4���9��~���r�D4_��qx��j�Qо��2f��}�1m﷖���{��=��嵇���2|����Uo��[�*�ԩ�tԻ�{}W�[��bF.77��&T|�w��.f
���k���Og0�^�� U��*n�;~z�m��*)V'��Wb�E��=����t���>N��}�����xN�Au��M6�x&h�G�h�io#nbG4\�z��5�)܊�uf+L=�-�����9=��Z�be� �|��u.=z�n�D���]d.���b�`u��E�k�;w�p���^ۧ,Z2��:�u�e�k�X]��s�ꮻZJn���#��_D�ҡ�К99�ǆ@���2���C�k�5��g7M�Hz���{�kɺ�d�����=�nUl�"��D�:���^�7]1�$CZu��vߟ��L�WN�p��T+����;dޜM͖��-Oog����r8��O`���v}+�˽��F�E��Z�k��H!����7�c��������d�����]{��_N[�E�+�%��\5�S@��T���aq��چ�<�>�E�>��δ����żUm�Y���㖃6����^����C�!�����J_c�}�͏��Ӯ�zJ��|�;�Y1z�$��OTGh_�z
_E^�׉53��_˖�1��I]ֶ(u^쐧&7���zkG���6/"0>�<�ą�#`F!ʍ��K{b�v_m��7�U���ԝ��x�1]RM�U�����p���u��e�AT��I��cj�^�a��G�%G��80�F�O	�!��*��«̗��yu�i6�R�'���B�Ǿ
�[�Y�W���-��e-�}Q_!;�q��O���jǃ�i�O�1����S�zQ���L��M�y�l�����l���\��͉���m��b.�qŽ�5e���l��Ҍ���tq�VW��[Y���v��\8�]vU#��a�K��+N'F8���ﾐ�Y���obBZ�ȷ{�/e�����}i�X�ͻ�m��2�WG��k�s0���;����9�<6��#_y�� U~a��/}e�x+���7;��Za}gBd+�&Vm��Z��j��=艱|D��K�ąm��5u6K�;1��XŉTV�*���
^�w��ص���c�����7���Ի9���&J�� �p�m6;���-��U���ݾ�w����@��A�YF'B�G�f��LEM)�g��di���w
Y��v[//��M1x�;m�.���)�cio(�{��+��a�^����8U���^cM_f���a�L��{L>��|h-kQ�V����/�l����7�c!�v
�/p�a��^�Gn8ǎ^�!���l�LR��aW]4�G�:(���|��T;�Y�����.�%����s���Ǿ� ��Sz�,�ꜽK��_DH��J�-|z���Q�o������i>����0����uBs��r]�Jy��P�﹂Y�ħ�h���:�[o�~�BUĦ�/ht�P13��2�{q�W��t�M���3s��d~4b��p����b����k{��ħv��a��?�f��#�E�u���"eL���7L'�ɛ��E��E�^[���D���{h���ݩTy�%w=1�HT���k��6�^�{�^�`�~�`O<k��c.�tr��tȫq��D�Y1�����z��\����v��z�(&��k�U�=!�O��]x'=p�ʡzd��x�z(S��\<0������B�@H��u� ؽ���X�<|�7{���{��C���;9�*�n5mow��'5��ґ�Rꡱ�k�X�H��<vלp��ϵ���1G@A�ӲM�ܙV�{Y;�$����N��=��7��/#~	�٨�O�ʥ�Lp" �_��y�ڥ�z�?{���-�Fw�O����� ���c;���T��БxU�%,g$�³�+أ�����`cQ��^�++�`�O�!���"�y��©�C;��f>�Þ�Ӱ֛���r�*�C�Up\ka�m�%�4���3�u6(+e�U<��S2���T�,,0&"X���8�\=��W��q��]��a�2�ñ@;�K��#sxʆ7�e����]v�����I<#��@*{K�5�
xs�g.l9��3�]��MV��&Lf��I=C|f:�~D��ޒ�T��f���L.��
�{�p��C��!��V!V�由��v�O�y'L����:ȭKeG�z��:��+Eۇ�E�ESy�LP��ܶ�Rй�]n:�[��ĝߪ��`+��;�X��F�Rꡉ����0&i�����X�D�3ȭ<�gf�>Z�ޛ���=�EW֑�u��O@/��3j������C�|�I�,�]Ҵ�OI�b|��t�2NͿ;H_��xO�54ᚠ�ʭ��m�()�XB�1��4*<��XVA<��v�պ|�0`J�m����j�꘽�P�b�0�9ݠ��YR�b�a���/`>��Yؤ��u:����M��Y/u�K#��A�������Sϥ��)W�;��+���:��œڽ�v�9͜R�ذ�"����U�1]����T��oM0����%�M�zݽ�T��%X:$Ռ�JU�a�B[I1���VzCU�1ʊ������oF����6#���K1҄IА�WCd�©�T��$�u�}d��6�7NA�y�W~mά����>ӢY�~�/b�i�H<�
����L�G>�w�������O�>�{JZ`��V���p�tޔ<5�vD��)W�	�Lj��K�xo++׊f"����R�������m��oVun9w�d�I,]_v�o9v�	x�M=ڤH�|���K�����5��ri�+ig9�`ul�hUj�s�YhK����Y˸�6r(x�-=p�DܫrnZ���-�����������K��6K/�W�So�ˬ�U�Ԕpkؙ7�u�lM�:��C̮�F	�i���.^��W-�>���2%�	O/�N���z�n�xX�.��� �,��Ԋ���Ǌt�g�v���9p��X�g�{�`�o��
���.�HE򸻞�g�W����р	�^bOO*}L���$=�>��ih�b�R��g�y�3��J��w��1m�Z����=̑oG�&�T"�ͱ8��c��BR�)<CV8��-�ڭ�*����U@�A��0�Z5K��g�prք�(u>Z.]��j����<�Z��C���`��$WB���|��o�8��,.sU���R��ݼ���l,��*&���8F���<B�x@���Q�j�Kl!��s��_m"���*�5�������V��Q�ǘMx��L'+�b30��ic��cf6�^��{��������/x�(�׍���z㖃6*9f�ש�v�s��������*�^���Y�׼�2�����ڠ��ނ>�ꂔ�����[��/�xhİp^�ò�h���{Ѕd�a�%���y���F^��:}�wS�]��YŶr�C�9X5(��N&Ҝs���%A��W���[��߫�}�/d�t=@�&��Hq�^��y�\sщK�*8EJJ���A��^��_
.�K*�R��jG���7պ�%X��>�w�lȥ�xD�![�b}#dBs�m�Z}�.�l����ۤ��?!�s;"��*s%�4���s>e�t$� e�;�FGX�sY��]�d(xhUZE�k���Xy;��K�X;�Z�(bW�l<o���-/{-�}�^ q�l�&n��4-�~�A���!�B�/��*^I���.�oz�ֵv����o'�`�$�[5�K���x��M:�z���o�;��x�Y�7�ũ�.�
Oqu���������ȝkDs��OT`�͒����z_/i�:J���T�q��yR�C��S��oW<�ZcM�}^BP��f�
��\g9T}�l�؄��c��XuH�����=[+:��f>�����B�11	�������ssT<�����@H�:E]����H�I�dSGZ^�7��(i�cN�g����K&���5��o
��Ӯ��`.�e@�ISI���M-��6��O/FT3����k8�?1+�h�s|�����	'v{�U+��ť�ݷ��j�ާ�9��K-^�W�'\��O��n%�����GY�w�%�3��p��a�z_o��[�m[�{��ꪪY�����߼ �EW���??%�֫�^��@�xM^�U�6�2���Um���7����Gy7����9-��s7`d8�,��mj��V���e�A��h����U'�V�gΓ5(�.{�h���^��6��i���
��8�Cy�Mݞ��M<�.ƺz��<������ל�9���w�)�PT)���P��Պ�|֜v���w��VNь�=^����&�Ʈ��Z����GH}�O�Pk��v�3�S)Mُ=���0�pH�<��*|Vh����r��9놞��܎�9��Fʝ[���l*��� �x<E1\�l^�E�}k��h�%��+3��n�zvhAh�>찧{V�oHS��{�r�bJG���Jפ˺7]sB[���^��B��z�g)��ysg4kQ���Ľu��?WP�{�=�!*������i���E9㉞���:�)��~s��s��`ھ�l�c�P�K�p�0I��*r�Z�Ж3Լ�)�s	G���{���Z��X"���>�ƋHN�٧_��Vڄr���K���䚗p��
���/�A�9����_�=YZk�X�Xg�m�Y��]���#�%�R�cd���y��G��-8椩Ä��W!�R�T�l�`M�����z���h������&׮ǡ�5^�++�`�O�!��{�M�[��ѵ+�Pu�e���-��S=خÔ1W�C�b�Up7���e_ն��M)gF3Ӏw�����+��I�,�u=���l*�W������)D�Ī4m�8�yE�>#�~��Wҭ���F<o�I螜� �ɗPVO���=��Ė�G���� ���ʋ&c������9�wH��k�}���\B_̓��K"�փ��}���o�"����������]9֏�2�m�a�*=��9�e�S��\=D�v�޿&r���̸\��f�L��O�}�o��T�SN�
͞:��|���w�e+혈��]� �{�_vzo��@���`Kyu��5V�-���3T��U���s�C.D��]g��W�b�W��͌z.;@q�:�%��~����}zX�
�f*�;Ɵ*҅si��#w쳰gK�������]�1����Æ����Z\+Qb�b�������n�-!Q�%ދ� v޻tcO���%_Bm��Y:�Q�����P)/���j�Ed���˹�� �]m���,,�dN�S��2�Mx�RT	<�!Q�W��咱�\�[$
p��r�4��u�M�Ջ�x�����'\B�u�0�wﾪ�v���d������9�fD���P��XpԶ�lh��������'���V����ǧ�x\|�6/��JfЉ:'���!6r��N��D�:���ʇH%_;�=�2v?%�6%Py��3��gz{���q��	R0��F4}S����{G����zt���q,R�z��C���Z|+J{G��׌�!�:
��P�{#�����U��{��7��]�-�^�]��b�t�W�D�_���ZS&�ּ�u/��^���;~�W=y7����^8��	\L�W�����嵇��/ᄹ�����z�ä@�U� �Ҭ�)?^{6�T7�]�ጲW�"����h�6+��^d���y�AUm���<p�ν-߫����<x9�Q]<�bzj	ᗍ�z�f��(�F��w�Y37C�ͬ@O9��e�|��z�ǜ$[��	�ȡ�m��Nv1��Ve�2���=[�J���{x��.c�Z�~Ԯ|��$�pVXd���M��`EWh���u�'�&3�6,->��Տ��.�y���C���#nÛ�YK�jܟ#�Ѱ�I4��l���'�ݹ
�˕�KW��,����f,�+���Q�b�&9J��R�S��vM�uȥ��\-���ffK�Ey5^���l��{����D
�kt��4֒���ޟZ�X�.��z\���\�c�A4�֚��b�}X�^�i�u`��%ց�J�����H�n���-ۉ)d�8��/�%Plwd�]�B��Ұv��g��3��þ����7��띢��u�p}���n��1f�d��
}�ҝG�;j��0��3Y�w����.��G*�������Ko"�ʱ6mѩ��U�<�^�b�����4�U����f#y����������Z=Qn*����it[F�]2ʵ˵'=�������Cm���{�����ta�7����.�z��5�n����B�I�Bsb\0p��;{L�$y�]�G1F�ҳ4T��]�iy�6%�*<��F��(b��w�z����/��]�`�Εׯ�v*Nw� ���I��n�N�Z�N�mm��WG�`��c1=ka\�y`ڻ�;��ͷ)���[��}�k��4��7��q~�u�e:�IΕ�,%ua��ܺ���;K��cܕ��O;���l�'Lvg�@�
Y�A�˹Dwj���}.bl�$��.q��h��*��DE�¨�� �wZN���^=��xQ�Xdڔ�&:�l�Cr�h�C��sێ���/!��Az�l��J\w�v���p�]�:��������z-�t�Ƕ5;�Ws���|�yV,*Ħ�v����ހQ͔'�� @d�s���7u�]$�ŝj��̭�B8 �����̹��s#��.��s�f�]���!!�vmh��QiQh����x7�EsG.�+�bjz����ʏv����K�����'��.�T:�LՐ�+f�w��)TC]�#Ր`���oM�.7������%Ү�3q�3��t��45�3��_.�E��2�S	��1^H;p���v�Jo��i�u�*��C|�@���
��e�ia���w9���@�Dw+g*\_s��w��"if����E�}�~����9�M$R7�3�כ۷��xC��p0S,Ɩ7��վ-�6+��6{��ew;;;IG���*�/�kr����,| �#Q�7��2�z5���:�0v���)�hɦY�f�yQ���*O_D���;�rC�gcµ�-� ���,�@d<�H�F{��\q�(��3<Մ棫V���:k�ohV� ��G]���'G�5Ɓo�sηЭ��\�w'�|�]VU�ҡ�CЩ�aDG`X�8�n'�ȩ_1�.�w���N���J�wT�۴�`5�gV���ْI[s]ܻN�g���]-,}�N�Uj����Wn�J�2-��=8or3H ��`ϳ��E#mb&�("���"��Z�*�R�Ԫ�X��+AF",Lk��(��6EEUX�1TF%�*TUUPTUUQPUQV�
�ŌX"����[E�UkQ
��X�j����յc�*�*��Tb�TEQs,0��R�Q�ETDX��Q��PUUb+&YEUS�VPDR�\�A�DU�b�TjV*�hX#Z0`�j1,,TDL���EDQDUF9k�jQ"�UL��UDE���4X��R"("��1�\T��ZTm
���b(�Q(�j������b�S �*���\��"�EQQ"��,Q���4��`�h�+�B�H�Uk�TX�PTZ�ĦV�1��`�b��U��T�+�hX��AKLe��`�"����4A31�,����P|w���$����)��'@,Z7rN�\oG@SȻ7^f��)�4gwڳ�!�J�s��㭦i�Хʔڈ7�w���qw�֒�����`�ˋ�I�!$o'�k����ǌ�d�~���Yd�ݵ!��CNE��S}똕��;l���2��#�i��A-�Kzr��������X�ݫ�j/3s:�TЂvK�/�n�Kj���kƇ2a$�48S\=Oʲ�;{�z�Zl��ؘ�4�(�g�o���-lTrԠ�`��y��.P�3u�O
�`��-͙���*v.K9�ڧ�]C�7��#�b��P��:�$2�S~���g�0�mm��ӴL�:&Z\9g�MA�O/^?xHe�z���`H_b7�=^t���'��}�W�;�ԯ<+�q�t����>
��t\���m�`�mzF��a��뜳����V���=�᷆��(c3΀k��m.9����|;�����a/�3���4Y����_wO{ԫҫ$����7�vF����X�}�����p��qϯ�wh�<��3��EK2->\\�e2%_�ݎ�~��m3\�x珄U_�w���Y��x+�P���g�+�D��5Hj�9�~�A�uu􊝯
��
�7�"��.�=�^��1���h
����K��b����^�yz�d\���9�Z�����ƃ�ur����-��O6K�mބ��N�v��e���v��jB�I�[9f�wF�nw�I��D�{�`��:"�-��ְG=�Y�=Q�Sd[��3�������N��ڋ7Ϛ�̋:1�o�s&Nv)�$�__W�t.�ip���Ŀ��cr�*zj��;��=ڔ�ӵk7m^Mk�-#G0|�� Q�T��*{���c(q���U?EX-\`[!뗙��d�?C�{�~�y8m���4�K�EV�k�V�:�%c���/D�P�RV��M$یx���{�ԭ��Ϳ�f0�@���y��2+��]6F�}��p�l�v���7�.�oc������p�3w[)S��aW[H�T_��@�p�z�_�8ߪ��K(y�-�9�b�Ⱥߦ��j�/�������V�g���T T�D�L����O+������c���5_���x��^'����_�N~��H���\N��
~��@��e{v��{{۝��W�����;V�P�oF=�����R�'�\*�ր�8�-z�9��ld�h!�֕A�����*E��֫���Y{]�>��k��� y�Ȓ�4���!J'!�{:s�5��w��e�Zo��I�a����w4(9�<ƄԇΪv��c�HJdE�\���{j<��ڹS��aI���\k�,�O@.�w�4D)���Φ�˵�k�fd�h��:*<�bo�˅RY;���Z�itpXPÒ�0����m�qؽ��Z�a�ϑ���x�W���4+�ѕ�]����J}#�	.���"4E�A�<pˮ�b��s>Q@�w��]�= ���Ly;��k<X��x�O�*�Cd�3��~:Um��l� K4,��������o_>�v�=I�+�����V���`����@)1=����3k׾3=��-کGW���8{��n��W����p�d+{�J}k���CE�=�ȹ��t掜E���� ��oN���гN�w�p�Or*ҭS�RN��ƶW���ވ�We�X3���KT�]�6,��*F����}����atz��Rۇ����AU��0�_-B�Q��o<n���+tȥ�O�=9og�.��� �-Ʃu���+�1�I�wVh^]~#��O��9~�0a�3�ԝ��2��{Eq	m����%�_�]>�FD	�ߌ�R���6c�>*�$�6��F�'��FL����;C��������u��sDlU�ҙ{o`�Aם����?��\Ϻ��CD��=گ䋊��Mk�2><7�@�ח�ű�-��ME���}]~�,�=W.�!�]���w�� ��Hϯp�R[Xm�o�7(�\��s�El.}�Z˛(uRt=SVi�Ĕrvn�����{�K�(����|ĵ��SN�
��� "���2��Մ ��}����r�Go�+�.rF�z�������z�߻ōi��>3T��U��w�%�5p^�B���&)����7Vp\��� ���S�_SF�y˭t	�*{)ݷ��zu��ɺz��9𞥆�zYԢ��^� H���J��5�#�;��5��r>+]S]���	\���Fn�.]<*�u'�^11h�5-��=�n=!��FF�{��ݾ�c(���w�3_�Kf���uRx��g�N�#��Ќ���΁/K-�g�#���{)*��V_���Y��
����~����.�'J���`����t�G�rЅN������f��
�)�w�fap�+��P�{!�Uxf�S��pi�;Ǳ�}����f�+[^3�gZ�{��+^B:�;K�zb��˓<b˜��S�q7�=��w<�F�����ZW�JK�꧗���z�6	�MvFV�B����c��X3X���;�e�³/=t}��Xfu�q)��å+�����۾o7;!�{��:]�hxi���+�Z#��Z�<�>&F7z�d7//���}R�P�Z���v*���/OfeEwN���r+�N�'�w2s��-��	`��Q*p�R�(�Y+�A�r�����Auf�])+�.X���5ϙ���)K��%>�s"�p���%�Q]<f'��/"�����U
�^g9����֦�5�$Ō�+J�p�\��.D��J�P�6��';��i����4�ƝO��/�D+�E�nf�y�racO�)��,
�e�J���M͖Wh��~�o�NQ!!-����O5���T�}^�dt��C
�uO
k�Es)D���2z����L,�Dc�J�Ai�R���5�C2�����|v���G��,�:5�*�Ѯ�KzG�d�%m��^;������ϙ|j�5h�\�~�R�X�/���,o5K��.# ���j�k�Kp�g<<�7��Z��W�}u�cT��z㖃6*9jİ�W] _?�Qݱ��WJ.�^X�ْ���)/��e֥��z,�8xF��!�x*8Da	A�75f�S��g�W�2n�&�^����G\��Z�k��Gb��Жe�ОL�u��HٖA�^��j�Y�g�vo�l-��y*�N	�|��[%Z���J�$���/oc{«���S�Ey
�Z���>�]ES����r<��.�� �+_>jw>F�M�Q֕f��ωL]ynT��M_.��:;|�k�J^p�R����Ohj��m���S��
���>��r�gWT���^��>��
���u��e�=sL����[d��$cۤ����aH����z�G��+b��]�_���EY6EN[�7=�Ǌ�c�Y���沇���Âd�K\|�u���^T6`�9֡��xe�¤^7C�=���C�)MN-~���ү�Y�2�{E'ҕm��l����x�N��ި6���+��J_i}�q��W�H�Ѽ��YС�hp���X%��B����"lx�ǫ�n1Z�n�m��Y�m�ɓ����Lp�6�qu6�B��&}��-�v7:*zj��;�:v�'e��y'l�[F��F�}�]Eme b��Bj)B�:��7U����8���}GF�34�o�6��4��dA��ɟ\U�Q�AizbX�E#C�Ɲ�Ͻ���n_0����C<N����_\��=3Y��Y�.�`�x?�x��2�6F��]ǵm݃�~�g*޲�ќ^���
���9�5����T�*�aW]4�_��
����N�c�˫�֛��4���7a��%�#�^���<��n���V�>�{q��P�Xf�%���=R��o���n�Z�xn6�;�Q\�� �;�������5�|��v���.��u��ż�5��F���l��-��<C�K��6$T�' Z��Lg�kE�|���SYx��m4{��X��jq�X���BH�J��J�XZU����}��.��]z����&*�����t�PO����h]��셞}�-Bs�	�|�gs�"��#p�J����ո�;�r�Q��ʨx�r�{B�ɨ�~
�O�O5���C��"|�p��@0�� Q�����p��Y�������^��7o�ˤ��|[�Z���5�D�NS��m] �����#�UW���c�Z�F�Ý�����^�I�o�A�����bF�`�%#�Sp��<je����w�X����J7i����~��ޭ��<��YO� �}YY;*Pl�%�f�a���r��ھ��2\&k��f�[>�睘�!��}�z���bzT~�40��v����>�D}Jv�����w櫂��f�o�����bVUu��<0m=����ex���;�@L�Ǿ��skhx��tb[`r��c�z�tj��LM�x�W�`�x3Jlde��y��h���\ݫ���I&�.JZ�j1{�N�}%ؗK�[[����8xE���5�Tm�u������xD���:L`�GW������wu�\�y�ȶQ�q�v(�7�V�F����8I@cȜ���)��ͬb��dzT�5޵��=����;��+'�֍�,�]��JK���,p#`���ɼm\�},��fTR���ON}0�ˡ��F���R��I-3�a�5+M]۵:�'ϫ�|A�V����2k�}�6
��W�����O%��`�qǠ�a���[<}�n�4���R/ez��	��U���p+�=��{\([��_K/|B�9�i
b|J%�D�e������SNQ���϶ "���2�\�x�:uw�-^�m֌�}~#gܑ�^��I�S��7��\y�G���`
P��:�ӛ�\���lc�j;�eJ���ˢa�,�X�h��#Om �^�WmP06=�kk̯EaV=�Ke#<�+c8�Ca�W��R�mˆ͉a�B@�U�G�ip�G�W͑{{szy�4���x]9�n�}LHo���τJ�lH�/	��XpЖ�OcG�����.6ן��o��٫��՘m���(�[�x�L��t.OYAI�WF�J�����8��#��3`��|��W�������g6T��z����tu>+��/h�~J�غ��vЏ�4a5����2{=�õOI��rr
�-89oq|r)��c&U�m����,Ӏ&�d�	ի;oz혻z��@��)�w'���yV�n�q(��@�^��7�ǒ�̮��Qε�f���/���Q�H<���T��������B���׏ܴ!^5R��⢬��pҫ�Ul�-�٘\:�J<5fL�:C����*��H��U�u�+l[����p�O�������ԇ՗<���&'`�Lz�ޣ�Mi�M��v�E\8.: _e����%xd��a3���"�M�+��|��Or�]�*U�T�j]և&[��Uu�ѷ�/��k�V=��Х������^eo{Յn�`��F�ݕ�q�#���ON$=�&l��l���^|��-[�{���@Wa�#�ܪZ��|e�H���J�*_s�bxrs�R~�L�dG�o;�S~��Ԙ���!AabkR�1��:l����r�XU�Z ���֪���v�\�~�&��{�����^�ע^J����W]rvɺӁ���U��I�}���o:�3}DѓrXf���|� |v�z��bQd��j4V�h�Ύ�\2R���B(Y>r\+r�W�a��啂�i�;�/�����MD� ���ev�5�Wh�pw
b��l[{a_�&Ρ��]e�K����[�������]���@�4���ᫎ�v���Ĺ� o)��9�uBg#w�Y�'s����˦u�C��<�1`�5
7�Խq�-�Ci`�/�S^4=��K�n�;O}��j�=���դW�p�j��W~�]��8��ck��a��^������JU��л�m�h\�O)�sp��nZ<��WU�k�0L�m�'a�f�-@�I�ϧ�#�-OAKnWzF�B�����K跚��r��H9��T-3�ù�x�ֶ߳��e��'� `#5F�T��|z������##r�6D4:�bV��T�jʿ�T�z��^ՄV���5i�����M��ژ�C�\|%P��\Ǟ�q�5Qa�"�z�G����ʗ~��_�4Y��b���f�'��=�jT諉��JU�Oe�&4�Gdh[z��)z�7��^��`�=)7�Y!���<���Z���lM�]fPΞ�I��[=�ɹ��x�N�[z��������b�S�|=�̘ͭ��k���:�-@��L��V��x΍���P�2K�Y���7�Y��5-�'@����ի>��_������N�EB�:<��]���9ʣ�o���O\�{f`�0�7��/iYu�Dw��Z�֥�ai����K�������%�Y|���_��ʕ`2�<ֱd�m����Z����Dt�Rw�����Ь�H���;s��p6���+��@T�����U�R���g���^����܉n�b�T�T���V{�o�_G�8�Q�]\�C(
5�Nl���ssx(�V�ݖ6(�o%�����p��t�$yYx*�U	��2��p�{Ţ�[�-˭� I�㨁���٬�\7�=��-���r��:�2D9I�� �j�؎�s)ʇXlX&�Y�x������g`76����X�F9�	���)j��+"��f�����G}v�Y	�5��Rrmt���%]�!�iN�ɜX=�� �M��:C&F:;��=��t�w�%bήm���iG�U�d,�PY�����L����x�ا�rS3[�����:���Jl<�ۡ�k�M]#W�s��w��̜5�l\�S����r�"[�)��8q/3�,�c˙RŞW�$q�#�>�l�ש.�Q�ƴQ�.Xt2�Rp@�>��f�������2�gga�������|������-�4f��Ꭵ6{e������_����֡�ӑH��fQ+I��j��4���3�-�&h�7(���陬^�����*#�Q���8�4���7o�5��������6�@:��+�#
�Η1�eZ�:��&s��D;$`��uh������9�E�Jz(��AI}� ��j�r�,�A�mbc����%'�oB�C�VܱYO�t�y��;p��N�{ƀk���4�
����vXD}�	�ॊp�*�:�k�]`la����N=~=XZ�޹���طE[���B�@��v���.��� wx��m���S���+Z�>�\�z�� ��އ��ݧ�ӭ��/�f�C���˰�&�'Z��8,�CŎ��	�0��k�ݺ����@��><2n�^"6c"���ȥ,۰��i���
��-��1�n�����Ù}����^<h�bw4�� �.Bl���l�xgU�[�9LRcdH.����]�LC}��h��3C��>:$��4�3�كx���n[jKCޛ� �$�о)�Ε�b95V����頭�1^�2�&��]�+��^��c��(Lv7;����U�3���}�o�c.Ԕ��y�5�ȫ�{Z�ُM�N׀a�\��
�n#(�-�[���Eqgk��F�XY��/p�C��Ŏ��t������/w�#k$�	�規=��b
L���OU0��i\=�KL����\���e��4���� k����G�S�2ayn�;��iknI�������377�Qm�+�Ġ�l[�� �[g�()��L�����{M]&�qh��M�s�6�q޼��C�{��K9���F��s�6>�4�vڻ�e>��ۄ�@ (U@A_��T ��F8��"�E̦�
*�D[h-j,Y��+Y��[6���V#UF2�-A�A#B�Ơ�Z�,�j)Z����AU��Ɗ

 �cZ���\�X���Y2�+���E*V
����X�,QAEr�8�\r(*�c%��V#kFڢ[F �D��lAX���Q��V

�)�V �Z�ETR�Q��Lj1TdUDY�kV��*���E���X���1�`�b ���9�E�m�,E�`��E���QV �%j�J*��0H֪
+XU�����R�E��X,��cm��J���[J��J	PEQ*4-QEq���ң�5��Ҋ(�dE"��,A+Ar­�Q�
�ʬQP�VV�bZ��j��e�ƈ�Ƶ����`#djE"�����3���޷�O�~߿k칇�|�0�;��&m�\��H=��i"n�S�c���r����[�,#z㳄��o{/�9Cn�.+����}��yÖꑳ�S�YHW˘�Lp!�T���Ǖ���oy����`�k�l{޳�O5X.�#OOmLۃ��h�k��cSLi����[�%^�\��oq���J�9���2�� U��E���5y���a|{ǈ@�xAf��sd���^O��{��p���0n�ӟV�U��ʆ����R�)}�®���#�:�`s�b����T[��8��W���W�4��/��h�{ׁe[Q�G*h�@��
�7�V��w��_�=B�%���W�Ly�+�^'��������2��.�$��u_�՚f������0*^�A���T���a��Q(s�Ե�w��!�U���Z��d�Q��؂k+H��u- �G_�C��es;�x]�/����-�Z�	+{b^���!�[�($.�CW�[c�u�B�¶H��5)�
%Z8zg��M���q�W�n�ʦl�ү�p����t$%���KJ��u������͓�D�hH��l��`$_f�ș����BT��]N#�K1�~�BeE%b��>A,Rm�me� H��tfh;��c�U�{mK U��jU�p�[�����5�����;��Y�ɹ�F�����7f��\��!\+N�KKͰ\�K#��}q��j�C���s�Eٷ~پ�I2�:�OGYsۀWݰPt:P�hH����e7M�T��΋�a�I��^��v�*�V��pz�^)����V�ϻՂ'�����
Rbz�Y�94wjH��[�Ѽ��3�|�^�8z/J3գ��e��/yA꽎ǧ/0)7׾P$}�;`�:`�DI5V��ޮ���n� ��iF<�]!��U�ޡ�AL�+�0g_:�c�G�}�-�|6}�t@�����	u�1zx�9�3��Q(q,��!F�}k ������*�|8�`�|Ի�;�=9oKUgyc����hL�V�Kyc٠Ot�왭�2eh|I�D���bk�{�`�������գ�ul��*����z�|��PΎ[NT�<�ȑѐ1<�ѓ(�|�j�~��S��Wb����3x:4.&F�İK"�i���y�ŵӆj��6 "��|�Nd�>�$��;��z��R���و��uH���KyKa���]m.<��-
f��G~�G�g5Wr�L���+�Pn!������oxάѻՐ�i���]��3�k��5\m�/B��|�s�����g���Z����3���4�gT�.��!��/Wm*K4sR�fjo�V�!��G����w^�r��B�!�ʓx�"U�&���#�ܘtl��&J�
׎�Ĺ��Z,xd�,W��^�
��z���-V9��̚��=C�<�j2�s��Z��xi�	�XnOK:�P!�d�2��+�G%�g���Ք�spV�B���ҷ�C"�.X�T<dI�%	����$?X����!r��̫��ۚGb�Ǥ:��;J��OkZ����iP��Iк��VP��7���h���{^w{�՝*���i-2�Tz}���qR+/�eP�2��E�U>��?Td��>�s��B=��L˓w/��'���sj�BƥcC�}����E=��-�ٙEà�3�o*���n��{ڨxcz��3��1��߱b�:������	��^4��QOv�ߵ�{�F=:Tҳ�{���=Mz��$��Sؙ77S���h��Ӄ�ܶ���J��Ip�nze��i��۫��ўx$}w({O
t�R��.�p�Y*dPw{��,��|gWm�ƹlIN��!�K�v�VHE�\ �W���WO>f'�ӞOơg���^?䯫�`��F�����ZB��ݰ�қ<Ҧ]��]=��i>����tzK�G�w>Lڊ��͚;|����s7a�8�ݛ�v�����3��4���J�q��cPٳ�;�SK�����/l,����k��A*GX�!�bt�ʵݺt^9Ϟ��8}�����z.z���/�`]6�9��P��؞��c���_.�ydM�9Op��tB�x���k\�=�TM�<��\3<2Y0�U��]�}1b��͏��O7o��ҽ�o�"�H����+�_(�wy�If�]�r�z{}�J�k�IwN�O����\Y��� |v��Z<c$sǈ@��5�Й�)��$p����������s5��b�s���^��3�����^��ܡ����4:���K3Vv�s���������XC�,E]�羿��ĵ�$+
e�^OK>tk��J{.���P�w۹�ɡ��Di+��5�A۞�߸���f�-@��ca����ӟq�y`������#y�RH?�KԨ8�ʿ���������������0=&yv� j7J���o�N���Vy#�FȆ�Y,J�W��ՕUH��E��H��~{����3�����d�W�i��".���'cDj(x1�#OH��/���Q�tf+����=�f bqs����ƣ�E�r�z�`�أ�:������Y��vsč]�yL��qSL�f�83V�ű��(�-\<T�G�c�n�S��{x���(�o�����b�+\�M$�U�6`H�wG�e�	���\ʣ�7y�>�_{��7]٪	Z��K~��y=��]	��7��mꂐ���#�}Y�A��i�N{|3O#�}W�w߯�Y�3��R})V��e�no��&����2�֓#s}��aIs����A��T�X����8p>";x=�.�;�HV��`�������'���]���oK�1�/i�Ӥ�H�^U���+�������7���_5.ƣ;��'~W���k�Ԓ'��fu䈰��������j��O��.<�)]^�b��W�e�L��ÒUNP�G(xߧWbܞˇU4x�Z^�m�)m1�P|2����#g��-7�Y]]�8h���"fq�ߢ�k>�^�ݗl0���ƾZ֣@�E0�Wk�,��׏{}���j>^�'��ӕ��W\F
�VJ�p�hz�SH񗽤_�^H��_��r$:���7�<�iu�J���{�<���YmFq��-cr@�R��&�6[�
�\���R�|8z�>2��S����]��^�3y��CmX��r���=�NJ�[�g@$~^��2<�b��2.���YN$��N
 ��0Z՜��.�t�A���4`pw�(����t���5�����;���>�\�V��cb�w�3[���'+.Vg*B�?�����xU��m[�*h�oZ���oq�ܰݮf�
�4(W��KG���y�W�L
�4x��s����`�}����s���>H9�	�gF|$+H�r� �k_�C���T���G�;�o�� [����7Z��E�}�^>'�*A�6�������x<E1\�׋����_�M������9`���ϟ#�oK��OAE|�ۡH�,$�p�n�k�mf(Ez���8ÜT�/�Ӯ�o��Dx�l�{�^����2�7�l��}�юEz���p��G��WMM������x=�F�J���<�YC�qz7\�.�Ղ'��� +�~���)	��o�y�}^�M�]Є�U�0N{j^�)�C��![�BS���*՞�\-�<��F|E��#�.��ӝ=î��������[�'�ΰ��'��P7)�tV;�O9z�w���]f�U-1/蔳��鿦�n}-h�9�����2s�h��q!��D k�:���n��6,'ϫ��+�Y�1NMK�2��=9P�o��B2ãVhn5K���^�,^n��&������[Ӕ�z�b�7����r֤�s!jSf7��#�Z91���u��Xln;���(]���}8����W�e!��ܫ�t�D��;5�Q���5&��j>(>��s��hĲ���Ժ}k��u��)#�8�n�vŮu�X���Ih�O��BO��'�����BMbo)]�s킆i�n�犩͖�ɝ���� Y;�8��i�6{�#c byX�d����a�TB��A�}�;�q׶����Rg���ZQ,�Y����)�-�����PVel@K�g|$����>��vd�'��������U���B���m|O3�Z�X�i���ͥ~z��yҪ��/w#I�Ο)C�z��}r'�e��ܴ
���~ 
��P���v�d�,�o��{��|�������K�R��w��W��嬯���4%��Ĺ-x��u��*o���8k����+�eP��૖�n��Sr��2�x܍R�(MW���h��,δ���<m��S�� }����~�^_{�r(d2�96/y��>�D�		t/�p=���Eٷ��\��Q�_��'��>��yh��n�&]���nC+7����+Gηgze�����4p�� O�x�T�ʥ�#���{P��}��Z|(���&�dxWՍK���E`���wEmv���"eh��ܧ��5�5�ln�a�����֭39};T��\������D���b������3O�3�ael����/Hr���s㇄�yt�j�^Q.��]��۽[Wv`6���ߎ�1lw�lN�6_��V�r��,�xXrv��{	l{�:
��d]C��7"�X�T�1S�zQ,\�(ke������֨#�Y�G���^-���C�Y�,4;%rV&=��NݻW��V�Y��o�	q�.F�K���~sz��%�Zk2������R���K���d���^r��
7c<�
l��-V�Y�Ia�h�{�q�W�"ޮj����k�]A!�3�'o�5\)�}Ӆ�ʹ�G�B���R��*��/l���9�蠤�:�_���n�����E���=��w�'Ӄ�+��\b��,,q�F���,
����K��g�V`�=�������ۜ���u0�so�`�[-���D08���̪��5�m��1�@�J�~�B�������0`ܺ΀ps5��+�;�h��u�4J�a�a0p�,H���
�'d�utE�*�V-��Q~�^�M:�����)cm_ì�<����/-�^z=:�rQ�9��z��5�x��x>��R+��Z��%���F_��qV�32�v%	���#��Ͷi�����]�`�O���՗���-,Ӭ�r~�K��TWIן�K��x_Q̑TĐwU�̽���F�������ӽ=sݽ�)��X'jN��'nw3��d<*X�*�F�"u��gS�,�|��:���[��%�^�����˭K"�賕�.����(GC����|JK��g)�T"�p�������&��{�,��i(;
�L_��U��-W^Q�n�#U'��6�n��Ӱ�X�����n1P��}�K�=�A�տ%!�Yz��Т�:��k2��O�&�W���&lK��$/�+�u#��x����1��@5���D��Oʝ��oH�+�m�<�#Y�դ�u*[|��t:,��,z�c��
��������%��v�c�]����^$�uWˬ��Oh��R�{%����	��;��� Ћ�y��{�o�3��ס�[Mr��W�Go�E�v'F��y�( Q�ނ��~�k�ʶ�K�ȚX�yd���n0~a���ݡ�H�Hr����c4�M�!��,�f.U �u6N-z�Ϥ�؅̕7^|'�8�F����+e!K�ԇ/��J���e��@��7��4kli��p�%8���`�����3nϽh�����cH~����������]Ł�xn[=�r�,lh^]H�`А�@Mm�����#V��,Sld@��7���0f9	V!���rpN��Zo-�����])u��D跬Tyҳt�ӿ�Hw$ώ�`� ��ݜ,���I���%��ԣ����L�a�X*�g/�蹚�F�2]���7�z&-^8g�~�m�@a%�ɃؒZ}6F�s��x�)��df+��p�3{+��v�
��| �f;ڊ��ܢ�Y�o�:T�Qb*��vҧ���9��=I�^�mFq��5yo�wdWY ����ʶ}��+V�h,,�A��^b+�&<��;��_.@V��-γ;#��'׮�S�- �#�0A�D�淖�����P�Ə������ȼ�̄�r������Z��h+�
_V�	cpw��U�]�C�n��a����s<3>��0���^	�\4��zr�Cj���i-���r>���ӂt;`�޾Rƽ�>������}Y��ҡ#�*���bF�`���p�n�c�P�M+d��5w��eɻ�VH�r��!����&U�OG����6�z�:��E|��U�ֽ��O�.��.�l���J�FϦ�/4��y^)����l��V� =>��|��@�K���D#�Rꕉk�kE�5k�Jx��U��Z#��n��51N�7| ���mqo�P�\���4�Ŕ>�Mj�ۛ�%�k��k��R����"�C��gTջ�7�ݬ�	��I�E���ٱ>.%�;���k	<�k5�0�]�m�/Q�TY�œH���Q�nF��tS�_[��Q}JK�ρ��;�� e���\��8��zV�詊�ˠ�n��
@\��"X�3��x]��Ϛ{�BpqE���,��v��8Xe��%׺��m�Y�2(wϪ�nx��-�|��5	(�V��M�����G_d�iX�:9�7�m�r,gn��k˨Q��Ӌm<0N: ��,�WnCѝ����� �Kq��8]�����Ei��EƣΣڅ<ښ���cu�c[�s��7-WY�a���Z��fh��֋�W0\��7����FP紩�&ʽ"�����X��خ�]�#{�;�X������z�?N4��1�Dw����f�^Rwm������d�j|7&��n�� +���g��v�G��"��k���{�.�5�|�����>��L�]-KpS��Q�q�9���6��c�9{Wf'2��$X��I��覝;��8�({iN��3 �;r>������.*wp�܊�s8�I\�n����)��q�c��� � uK���Y��⽜�U[���O�(̓I�391_F�Y�E�#/ (@��5d,�fVE�;WQ�(��U�;��^�>)Ҹ��	���V�s���Xw]�7�.��(���wNl	rS.�r��'�WQ�T�}ݘ�W<���t�!`˜�f���V�"��@���X�[���E�y�%��4Q�V�{%��si�A9m���P�Z�D|�Z܅X�'w�ww6.��v}xk�]��ɺ�R�	���e�s�Pw&� h��Y.� 9;�cәC{�{eT���ܹ��4)-��f���鴾
�wd�ν�9d�Pce���2fF�"��]h�������#��}z�f��{dK#[�CZ9�c��t�.fI��L�cB����Rf�NAǑ;cj���
�͵x��	�nծ:�9J�pU�(G}9���NG�;b6�rnM;Cv���w8��R��[xtm�6��^�9x�q���Wr�|�+b���9w�X�XdR��<.�e�3�D�3B�F�m^�ε3�s��UF{+�ܽ��M��;jg��ȯ�1��NӬz�����:[r���ԅӃLD>N��q6���~��Yg��bi�;�����1\̦8�:�k���6�{�;���O��"k�B���u+�2e�u�p	F�t�cX{+���s{5�21��"��Д �u;n�w^n���c��e:ɾ3eZ�K��mC�q�{�7�r���y��%;/�Z�Y\�wu^�i[v��â���&�UEBںmj$�R�U�,Eh�5(���e��L�UcX�(+R#r�"�1���X��UAU��F
 ��+�kQV�QTDq
�P���PcU1����֎fb��TDDcPB�
�TQ�Z�e0*TDF1�EX��E�c(�Eģ�J�iV2"-kDYZcej�Z�L����P(���lTQ��DDUEq.4QTZX�b�UU\��"

DD`������*�U"�V#ČQZִUdVe*��P�TE��҂��ň��b�C
D�%jT\B��a��J(�DRڪ�Eb)Z� �ib�R�E���eR�̢��cF*�E��
�h�����O--+"�5��-F��yj*[
�U�.[<�2DX�#�*	m�,�b �*�A��?�w�k����Ɔ�yG�;:4����9��5{�(k�3��o�y��DsX�f�qOC�N�2�6\4�%6uM,g	�Ǝ�wp:���r��/����^g�`L�ڗ�YL��FC�^�)�{���uJ;E���.��yj���E����bx;rF������c]"��.�qe=�S�1l����O2��M�W[i�m)k{˦J�d���,�/�]�ޣ��e�'�hTc��s&7^�Ru�/�f��S�5.���ONW���}�k�Le��s:���z9��w\$��ZI0M�D�W����=���^<=��sմ�^�hՋޚ5��YHz6�Բ+]m==u*�.r$w by_�&W�&�=��:Q�+�o�+�/_3����>�SW%��;���k�.�j)��`���Ƿf�d��K{�6ʝ�ANj�u�u�ruR0x�����ޯ��;��g�;"a�e���9�=�L��hΆ*�J��c>��<+.&.�!����{�X#Ok�����7�e��d�+���;���w�>_iB�����9k+���fİ�,�}���3���u�B+�Հ�6�1�{�h�n���%7�L̗�w%lm��`M�z�s3��������G_�7e����st��e��Z�f���.�ُ�g]!�#�iȈ��7���؝��k��fb������ӯ!Ȗ�$1�vn��o�tz8՘n��j���U����4����&(���V����T���A�~�o(�y�\WV�������h��4��G�OkZ���M�;'A���)c�Y�oZ}�߿Wot?�����8W�iW��D�Q�Uz-�T�pL�����>�7�@�$8��n>�k2�&�o�pbb&��|I��4}]n��j�����8��z�!V������h��(������׽�ŅMppvN�l�{�Ԉ�����5S�u�]wC����4�֡�Bkֵ�#�3��_�A�?c'��c�j��,�^�+_�����_�9l��֗/M<�1߀���ߏK���zDU������rT'�K�:�6\mu�r��cZ��rWF��o�o�Z�xU�&�)�<0��+�Kj+�����Y��M�^=v��]h(=���UXt!��V�����E�/l���"W�P��2�`�w���Y���6<n�d>o}Y���lK,K�t�
XX�@�u|����\y%���]F�rZ<��.�lw͚ۅ
�#p�҂���6	�=Ajh��zn^���G���.,����H�U�/q�s��%{GR^�%�^_/�o_&��},ho%eȞ�sw�J�	d�	ޡT�J�e�����s\��Acs[!xr.k����8���*�wV��ۻ�zǁCr7`K��35v�tsL���z6�iz|���#y{ٱ���k�5�5{��?kU��\L�	���&��a���|�$����G��E����*YS��׫�/,߻w:^�4iZ߃�]�7ǘT;a��(�v����E�l2�§:�+��g-6w�r;h-�J�oL�l.!֖:����.p�R�vs�R+��Z�"��1���;Lb�q�g9�.�QKF�2C'<�V���z���,8u��KP<���N��c`��h�COQ�wFI��pZK\�y��5ژk��Gó]�rr���w{'Bs�:gD�_"rB���9B6D5�Y,Mmy�Ք܈zZ��!��-5{��v�)#�/7�5�{�rdF�ؕ�:��TY�3]x��w�w�2z��W{���=\s׿QK�����E=� 5]=[^{��P�X�u��m��]�Z�pfȆq�|��{����{,�C�δ��[�~ʨg��PlxGl{;%�W1�<H��My�n{�����K���5���ɤ�L��/Y�;���-V䒰�W�Al޻GǷ�w��6��Bev�j�e	�9jҎ�}�31,���mN���]����@6e�n�����ε��������7�c~[I�E�B�}�n.�D����h7�ﭐ��o��m?�+��Jv�{�^�b[�
�XK�e�Z�.3i��{}���N��X'��/i⿱bU�֑T
�ꤤ*������)�{Z���'���=}�^�[��:6}��=569��O8q6��Z�B��5W�p#ٯ��i$���9IV��=��e�>����g75C�1f�^�d�p�wH���Xo)K��0�^ţG�����o���DG�����U��3W�d�A��~����^��٘���ل�;4o3}�����(h�}T������lb�r
}��!�f�e*b�#5fk�$K[흞�W)y�&��Qb*��vҧ������D2��*�B����� �M>�������].#����*�,bԠ5��Ǯ�^b+�&'�������I�����f��y{�wK`���6zƌ�.�,���_Ɓ��#8�������ո�1���}�^j�V�&�L{��R�r�yF]���,��!ZEҊ��h@
�Ou��䇎X-*	�{�i����!����KnĄ�ݒ���>�p����1�~��i&��T\��������J.��>B��L���=4įo��ЂH��b<	���gk}М�is�yg־E�wc���Wnb���`�x��x!ܠc)Y�d�h��n��������� �S�k�S��i��=9R!�uF5KH@�<�-��9B��uu�d�3�S�<X�M�>��Y��E\3e����t��d%����f{ ]w�t����ɉS<p�@�0A�r�E�36�=��Z���O�*���T�Z.+]��6xso{��M���s%��`C�]�)�좎 ǩ^)������3�X'*t1��z9����cm��ޕ��@l�v�9bzڵ�s^�j1���GNR��썻�JvN�i���.��T�k���\��Y�{M�U=��a�g��6��Os�Lx�F�ͿD�S�5%����u�|kau{i�m)gC<.lPV䷃0�z���c��{u��JL�}�nOzOg�z|�J�Cա��Y��:-j]��މ��`�{&]A[;s.Tv�B���~ݚw��'�|Qw�{�VzeԢkB��}z��*���@ɬKf'��o�_����I�<�|�u��PEx�[`�%�g+]Ei���Q��D�����艘zq�Y�E{��W�[��cb�ۖ���#�)���w����A�����M��L*�n��ZM.=��� /[�w�Y}�L����)�|�珷�ַ���<����L��+���2.�M*�ׄ�*�d�ʹ��,�ʕ�"x��=.�r��KS�3p����m`�YFL�:lvG���>��w5Y���cg�(�>�.K'"�z��E�j)��p�s��Y�~g'v��V��.m�(e\�x*�b#��h|�e'���s=(S}�V�m�c9?^{�O.e����c:Q��R��e�'���&./��s� h��� �)��ؾ2Ϸ=�COlA��(LW�1w����Z��+��r�W�\6e�Eic5�GSo�n"}3ǉ&
~^"w�3����_�\��2�x܈�u�H���J��4��ݜ����S�_u���h���Hiq���'���67��)� r~+[C����4{�糣d�*����	�)�TXU�e���^]Su�|˸�_�p����[����z���2I`zl��0���^1hB��+?V�i3KO�K���mw�k���y��ڞ�R��
�ps�u�qx�%N�G��������������J+���^�.5/6�g±�L\Z�a��+��3+��c\����f�����F-�X�'��2r���q!>~�x�=�ȋ�x1�#Z�
���\z�&�:[^�g�]��/u��wmksTK����.tA��\����:�VW����6��{�����Z���b�f++�v�6���뻵�:a0U�ٸc�x����=^J�TnJ������ip�T�j]��%}2(;��ו��Wl�ϧB4�>�n��|���+��=�����˫�t�p��^b[Q]7=�kM�i��g����v�Ŗٔa�����c|�>H����iUo�{e�H���+&�9������#�ꊯw�9/i9�'�s��}�?b����*kP���k\�=U�.TF�xz�Y��
yy+�y�L�bnl�"���AS��|zQ�/�"Ĉ`p=C �\1}����I�䮂��S��;������`@�s���;��_L���xϯ3�行��z�1���+,�T�Ѯ��-�����;\gW9�#�\�~�UȜ��FI�;�������4'w���br����(w������j]N�j�^-�d�U� YN{r�<�g<�ׄY�}u�i�49�%�%,� �[k��p8u��w��W_{���^��L��0��>�9���R��]$�qZ�g�M(9}��4�r�h$}N1IU�<����%�j��;�0U�é�ǖ�4q�os�毢��6/	�dnV娼R�����Z�RΔ3���>�6�U'JWLoA�p��7
����2��'���t%������YD�M����WPC˨���Pz�{�5o1�cG�=�xt2��O&@���b1Tl�z�Bxh{�j�N��N8\��8	���ъ��^�9��8�j3��"�H�v4F�(x0���Oiނ׭u,�����l�}�:/#�q�oM}~��E�y��c6Pԯ�
�d���ƛ���~&���:��򼃻�,�� �1�ߥ��ˋ��y'������c�(�(e�K�z����������z9�Y���M~����N?^/pM�-0���2-b�!ְAu7�i��k��	�o6Ǌ������@��������k���RR�>��2r�U۫{֮I��Ki��%K���C�%MןO8r�",*�ǔ7����W������]k��͈`"�6���+C���;��G�e�cg��<=�,�^G��FM�yO��ؽ���1�(���^?a���g.���k6W�6�f0����־g,w�H�I�E�X�<u �z+�1�F�}�q��,���;nR��c��7�����S��3���y�ze��%�Dd�I���`���;��g�ٹ��ӝ�������C�8g)�bti]x�uȪ�&U��D�d��;�<�S)k'��sH�f���n�*����������&��9�::30s�bӝv۫�HT�aS�H�Tg��@�pߨ�-���z��e�s}� ч�\s1�q����.ѝ��oͅ>�M�G*��� TϢF���2�����y���2bx��/��Z�����`��q���J�.}����2���vn���B�kG3��z��vɤ���,�v���y���{��O�Y��*�"V;�?K:0HV�(�ۖ�a �d� t�%O��Ȍ&�Q6\���	��v�	������x"ONH<�՘ ����=�=m�[�S��+{�7$���M^87���X��V|�oz*�2(�K�J�ŝ�Ѿ髷O��7����c���E�z7�}[h���P�xl7)��:��ʾu2��Y��n��Y[��->�� j�����`��%�b�n�jϦ�/?�*�>LpN[�����U*v*�����d�"��M����v�XU�$��\ZЄ���vS���
�G^L��-e,Qv����x��U�R�U��g�m���"��oi���\5P�X%f�J���ze1w�W�'��wV�-���#�x�FV�G�6�B)��6	�g����½�(.|iS|��Ƽ�)�k�MQOv�m����hq�@n�Y�>�� _a�:{�lm�NT=��
����y���%Ʀ�בQ}�l���<���g-��M�]i��1^�Ԕ�q�fU�#��86��麛����t���	���L�65r9y��b\�fM�g[h�a���W��q�K�|5��^A�'V�a>/�����9�>��)�5g1&�7���zeԢ]hp�B���7��$�T�r��&{�W����[7�"ŷ�ߒ
�����`�a,K"������t�Aߚ��{+�0�ҝ{
��{�r$�ypv���U�z���ɪ�x��	����,�K"��OO]>��VjzQdHo��U�.1<7����+3b*��̠�5a3E}�m#B���3'��:)z�����-Oo�����<.��SNQ��״b����e���<+.&.� �0w)�/.+Ȟ���8zmr$�(�k��W�	�+՘���c;�U��W��嬯r��5&��w�(�\�h^����w]c�E�ֵ*n�Qq�p���8���:���x��+��+]I�l��}Q��1_Vt�rΕRj���w^�"I���q��㥟E3�KU��7��G���	*B�R�l��6'B�����2�8{U�]!6�1u����l����$��5=i>���rV�x�G�]]1B#=�S��[�أ�	�+���P	N���+U4��;�p����!J�Aڪ�����{I�.'����8c�*�J;n�P�4��%{/3D��v�P^>���w~����F�I]���P���:]/m�vYW�F+�`�\<�rT/�d�iq:�A��_Y�9C���h���4X��AM�Wd
%ُ�k�ݴ�^�;��ٙI9�
�xH��nix!.J�V�p��ս���o7�����`�j)f45]9^��Qrͨl�$˯=�-�4ƍ��ɕ�:�1�mҹH}�o9������yEmJ`�&��K5��#�Y�=��Ε$����E`u`16�I��k��&oa}�u|,���_Ұw�w1�
��vL�g����έ�(�>?8^��7S����;�{Mebͨ
8K�������,�dmo���ˣٷro��|�4:p�0��s�V���Xp�ne$vu�Ǎ���%�5���_G�z��-���5�s�G.�{��w���5����I���2��
8���s�:��b��=��mE\�Š��ܳ�k]{��b��w�DY'��l{��b!$#s�An!�[�)�`2q�W-��ҋsX�c���ʠ�йI �yMTz?M9�Z� 4�*�$�F���X�� [��lv��R�v�&IB�������_N���i�;>o:��>R�ʝ)�l�Ћ㤬�7Sf���H�7�obat�n&'H��H�`�[�ɮ��^�9��xl���h⩻@�ou�8�ʘ��pYе��|�P��c��IP�����2������IajM�5�iWG�tqM{Cl�;{�5��s~o���F,ά��LjZH@��ت��cO��+�Wb8�)�ý�6��Z*��ͶE:���:p�|�v!e4�>M�	|٫;��D>��\�.Tyc�@�3c�_�[���M�t�Y��VI�Pn�\�E]�.�ռw��<���p�].�����#]\���֋��*MS6Ɛ����5�u�h\P����K��j�l1��r�n�q�#��<Z���6,�fy��;�a��A��gA�tr���i�U��ܖ�P�[�ŔN�bݷ]�cюwT�8��07�ޥl���cAf��]:8x?(=8j����g��h�����r�V��6���+@w��;V�ˠp]bN+�o ��f��j/��n�vS�P�|��j0�9�7���#1HGW_6���i�{��F�~����������Z.�=k����R���m���mLqP�h^ t��F)5��N���jҖ��X��s��ٚ4j޺]m���ж���:� wu^���sqM|z��n��D
$�(��T�.EU��TJ�"��YEE�*��� ��ĕ�0J�������
*�Rʕ\�`��A�UQq��Q"(>R��2*��J"��V[�0Q�����#��0|aTQDQ��G�W�EU"yj�����-*"
�E�aUV)YEAP���,b��"�be|�ADTR,E�����V�E-)�U�ʦ4T<h8�T����h��PUQ�E�EU�(�5AX�,DQEAU��b�UQSƊ����(���"�1�(��[h(�
*��Ĵ**��Ȋ�YQAA����UQ�_-Y�V
�"�#1C�`����D�T�E����+<J�(�Z�ePbcq+C��P�(�� (�hS$�}y�i�(ֺ�\#3ld��KFKs�l���J��D�b���yp��%�&M�j�]8ޱW��)�÷۪F�۝�y$8w��U��VPRx�UNҧu؉,/�)�@8��r�z��V����%�$7�}��+���S����Q��!|I��W�n��7Լ�^��Q�/j١�"�����b�y[�����
�U>R���{�C��7�h��b�P_+[]��-uf͹iz��lc1t��@vQ͂�E2k�k�GR�v���z��~�'��c�j*����h�u� ˳./cOvwV�[6`۔�O�����Ī�U���2���J�J�7�R��������/��x��z�i�/�t�)���%�΂������z�@֯1
�~{��@����֤��u��Zzr�0ȷ��K��^#H|�5�R�r����*�x��+ڸ�=9n�^�z)/����I�H��=:�0c�S�^�6%�"�� ��ƈֺ�c'z竼9��������Ӑ��b3����A7+���tso�lػ힤z6�K���oz\��t�c��ޜE_��Y�|�U��[&��bnV�Us�ׅ��|��v�Z<t^)�*�ͽ7���^����)�w�Z�K��y%a�s�=X}�G�@���Ϫ��&Eaa���E�Я�[�E���Wp�ϔ�M{���s���x��e�pd��ff�a�f���]P.wa۶ $��%`���ɣM87��LU��� q�����T�B� Th�8�}���0�A[GӊЏ��G%8����U�-�k����X���{���C�0�����z���5���.p�W�]x�YSr�����C==8�5�)x��f�OK7.�M;F����+��5uIAʭP��&�o��c�f�X:d����6圣�X`�����������h�^�X����"���ʺӝ{[k��紽�}O]�Lv�צl^̳�uș
�#�1Tl�z�Bh[in$p�ӝ�Ln�	�yv^��ۯ¶�yW�ٯH��A�ꚙփ��%9��TP�aնA���8��j��4�J�<�ŋ�;��̗��<�?���&�JU�:&4��{9����-ɱ7yc�[5�JTz�7�Ex^WQ2}~fl#�j{��OV���ޓ���4��F�;�ʓ���&���o�k���m:��ǥ���8�����K�8��f���5���$HV��e�%��y�ZߖbĪ+iAqN�D�ѭ3/��Æ{	�����;��I��gz�b��3��ȃf�M�&����k�+�,��Ԣh0�VkH�Z���u�jX�xh��2@�f�k�n��Q���;ښ,��u�h釗n����tV��s����''�6B�m�����ʜ�s�$x�ߟrhט�k.{i����S�&G3}<���4o����YHw�m�;�ol�P�c���^
P4���C���P�9���N}�=��;D1���]Kn��qz�}' ��^�#�^>�(�5Ù��2�X&g-�)�QH�8ƪK����uk͵~����Z֣Ei�Xm�"7�mWqC��0��W�\E*��Yכ[��ܹ�W&^vŢ�W`cH�d�Cy��4t x8o�X��itҧ���No�{r�}�/Q�sw����^�Wgʄu*"WҩƮK���=a��W��L��mE�%i*����o�{�S��x^פ���cF\�|U���T>`��Ĩ5����=#ܝZ߯x �x�O<�48t~d�]�5|�xeߎ���Z����>ϥ�<C$��4��%7�z��'n��|b���U�<�~<n�˯
��|"ONH<�՘ ����Zϕ�oݔufŽ�'���Ȑ���X��VS�a���l����F2J��F1`�����f�%z1��w���K�3c��ghh�\����JF��Irxc����>�XI���qz��*h���ʺ7w��ǐo���͕����iv�=�u���uRKdƔ佝�[�����Zy&�Pf��V`X@���5 }|W�ok{��<UJ��Н����,k$Yg����e��}�m(lf�i_��V���PP��s^�ro6ƇJ�p<��w}g�X��e�b��j� ǾW�a`)y��xO�q�Ż:�z��x�l�]ʄ�%��S�b��MhBx,	�s�R�W�R�G����֜�����\9W��~���`�o�!��h�7Un���u��Z/tyc��˗�a��+�x��9�fZ�)u{Ώ��2(,e�}U-a��=�dp�p��n�`�~Ii��l�h��@�5�y���)����,�Ī�b�!����P��b�*��pew�zbw�ĕ�)\Q��so�V��vL��[yaWo�.�or��oLq����&��'����s13@�.`�z���$�ձ�Eո� �(f����S,K"���_�����A�y�	x:Cm�+fj�]�k��(w����.M��C��߸9���Q�K'h"vA��;��Y�-o�s��pJ�����AY��U;e����04V�Ds��
σ�3+
�R���PW�t�Z&��/���h��xqV<R�z�#v�׳�
m�����4,F�妹�홛��5t'����Ug�s����e╓2�2�/�N�����[P�dv�y,�>�n���
ƫa|ʩ��q��B��b�=f��s��3����Ui���SH��1�h�Rs̱�"xVU\L]�@@8NvX�xjlq!�r����4I`#L�A�^�:��Y�x>�3���4�OR�u'��]7�U���g/>6gX|hu���rT�5�q�._g���8�V�,t4$�Zݾ��t,��{�X�|QʺqT�0Ki'���VzC��㥟E3�KU�>�ߛ��^=JOx]���䳚R(p���2$E��5�]uC��K�
yP=>���W����_�bkd��}������
},/��� /�`�����-W�V4<bSn\�u�uc\�vﱧ��6���+�S�0cGJ��|�Oc�.I����T��[��b	��'�O=��n���/j�:׊��[E2k�V��u*gixW�A[�~��n�;��͛~�wF��뚺7��0M8<�-�=i^��]O/S�OP�[�+}�p��K��ai1g�J����z��.@��6\_t�Z���վxU�'աȍ���	.�s����������Y��b���%�n,�n6���X�r8���z�+�nzźN&/J1Fw�,U��:���3{%mע��[}���j]�evc�f���:�x9o�_��}�ST��؎C}W�|v���/%��|9k�o��r!�j��	'l�Mgq���߾��My�v/�qK�y6�o�a�>jy��W��A���@���ӹ�%t���ZH�a}�p��؜T�1��+2�n�j
|ֹm��xB.K��,;wٳꥒ��Xb�&c@9��Xa�so�`�j���z6����ȵ��j�~�8�®)��4���;d���ܭ�
�s��=������lp���4����#���� ���x�ƍpc�����!�e�q�^Oz�h�/�V��f�H�km���ˆ���5���H!�4��]7��/�i���!ٻ�g��n��1��+�F�"��n�]z�v�s�����j҃�z�y����!��.g�ys�|����`�:���j�$��O	K�Q�#O�I �qz�|�镔�����Fi>}�]�v)�S8k6/	fby2�<􋞨6*p^�I�| iY��U�_m>����δ�~u��k�.�oXj��\�͙K����u#ep�iPB��i9-�GnV�L/��av���%��s�"j�:�
���K����<��/+Jׯ�������m�D��=v��U�k��Tq��',��-O6�\�3��1lB�͘�Z����|/'M�ݫP'��
t�c��T� ��lm�璄�FJ+w��?X�ĄY����//���W�/�f��B�l��v��߇d���}�͔O���r�M��Ą�=�E��^�6n���y�����^�L�_���Z��tN��L� ���t��K�v`�Rwl�x�@_�w�2��~k
�>+ppW��}gBda����+�ծ͛�#b��R�	t�B���6�L���K���*���IQb��)�{�BC:�Z��'l�}^Aк�2o�ĺ����|6P�B�J��'�9n�=�8�5�������~�9籚�s��}^�A���ߴ><�e2��j�Ü������Ln�w㻌�G�����0����#yK�CH\Ӝ�S��Q_��r����V� �xu�3ؽ�n�*M�ƌ���i����_-kQ��ȭ��X���\�`���<!�Gm��5G�oz��\��׭��Cu]�ACH΢��k��H��X�����O-s��C��>+Y�������h�)�x[Q����Y"d�@�5rX|������=/\�4�Ug�s��2�X�{�8p��C�t����N^i��Ch� z�\����.��f���m]ji&�*H��Rfbx_M�Y)E3��x��2F���u!�U���s�}rί4���@�ud@7��{�t�.H�<M���;;ڭ���k��B.�PL���t{���/��'?Xї%��r�՚s�#8����k[�p�8#��ی��'	���oh�׼�Du�*ןw������*��i��nZ��r���{r�k�L��;_`��-)j�lv-��_�b����;���Ӓ!��b�\/�<'�ϦF�0�ѱ�}�h����iD�ev�����+�=�V�x�������d�����t�#B�iAo<l�}�
�Uϟ���y,vV��|>~^<�m��-ə�߽7"X�RH(>�p2+��	�b��]T7�k�^�}�Q�R�c���*�qw8Y�L���y$���G�9��<��� �Rbz
�vH�ͯ�!�<�w]�S����V�7㕢U2�T�c9W��Jκ��8l�֍�3(f/�N����3y5�{���˷��n7�p���!��U�U�b�K�'B���*��LK�����|�y�}tϽ�kJ=GԽ��0�"�xk�����)mÉW�����X�|Ի�����{2����ѳP�U�ޘr���Ő��w.�s%n��R]���q�J�|��<%�چ�Z���н����*���<�u�S�.
arTtu
v����bl��q��˖�e^Kꂒ�kb�S-i�͝�3�{�7��g;�p͓.��� �*��E����ޙu(�hp�z��)�X��������+1��Ki��9P���W����i_���1ґZ:?6;@7�h]do~��^z	-��#hbyz"fܛ��j��
bݞ48�4�%�:������:�0���Ց�^+2׎��W&��3�U�l@Eso�C*�;�����_l�G[HЮC�q���]r�˷�ۧ�S�	Vv�����#���&zo�h�9�����O
Ϯ&-�z�;�oH9=��˵'����ǀcu�K#���zX��^��kz���.҅J�XA|b�rvnƃ�pS�-�w�͎��%����%A�#Z�8�v�~km�i�u���j�d��uK��C1���<�Ûg���#���Llh����A�;J���O?����P�<R�3����$�J�`�؉:U'������
v�;�D�Q�L��^�˧ηۅ�'}���W�Q�j��w��؀�~��
�`���D����W��8�h�V��f�,<�x�쿻��6֪�&�K�V�S�G������sX4&%�F�=�NÛ�7�5��l<�����#G!��:�E-Ɵ;�8X^�m�����2��(ΛڷKcѻ���X�]����8�b����3"�f�oVm�\8k|zS�=�(ɛ?�{G��^2=}���)C��h���n�DWgs��H��̍I��rR�r����Lm�|~z|iU����Ⱥ��e	(�_=��Mqû8�=MS����ވ���y֍�����ma����.K�����]���*U֥N�yf#0���)�J2J�dPwyˇg��`�V-tJǡ<p�����F�Z�9� ���=j���/4`5�%���f'���qzzP��Z�\�שE�Jߝ_J���a��.לg�BVp�d�z�X���2�i]�c��Va�)�(*Պ��)���t]^��<Yņ)�W�cLg����<�v�}�ɗ��o��ҽ�o�"d �A�sq�v[^��GG��&
��]
�D���;���3�,�h\ްˋ6�Q����Ѿ�^󬬰��#�hxS�<B��Ѯ�Kzr�����u��'�8��L����=1|��X��`zu��5qii�H#�V6��7���!I��B��!	!I�bB���$�䄐�$�$�	'��IO�H@�����$���B��$�	'�!$ I:BH@�XB�Є��$��$�	'�!$ I?�	!I�IO�BH@��	!I�	!I���e5������ ?�s2}p$��.z��P�(P(QT���� I@@ �@B�%P  PQJP  �$  
�B�@�$�$�
��	T�T�BURP�$Q! R�R�Q%�J��"��U*�%T�$�*�R��AD�j=4�AAR�!((�Q%H$
D�%P)PETT��P� �*)"EUP ��"T�HA*@:�D�J|   i� @ @�@iX�MeV��(��&ʕM�����PJR��6�UR�5m��� �Դ���)AJ$�)Q�  c�lBZJ���QV���m����P��`eZ��Y����ՃT�46��hPSAia)T��f��5�j�k[`�J$E(P%�   ��CB�
�� �
(P�nN��@(P�B��
(P�B��;� P� 
���B�B��K�P�B�   �p��J�����CT�[(��)��f)AR�QBI��w�  �ڡ��X1MU*�������B�jjU[h-��f�	��KFhjT�l�
[l6��J�0�[
i�4X6ضP�m$P���QUH��=�  �{j��l�����T&�e l�c-� �ƕT-�5���S[�Y�#U�X��M�, )055Jj�&����������   �=���j��� ��b��4J��4U���h֚hV�j���И1��6�F04,�4�h�4jڭ�*D�*��P�T�� 1�m�JUkjh4�̌� �cj��[jʨ�PZRڊ�l��YCM�+l�kil F6̪ئа��@��QI(�IUIJ��\ ��� &	�7b�C
��,�
�bcT �р�j
 j�Ԡ*��4j�U�PLJ�R%$��C�  C� �֪�� 5��( �P*�ڌ ,�  mT�(��YT�0 �0P�B�TP�H�8   68F����X�E���� S`��UѬ�Z�BDi�Ui,Q / 50�*P)႔�@  M�)3(� "��	QTd#Mh4�*UeC@  ��L*U=&��i����܌�C.1w���B�r���
L�K��ܳV~�1��K���!$ I>�r܄��$�@$$?����$���B����$�!$ I?	!R�,�U�j�u47Bp�n�L<4K�r���I��]m�h�5��i�V�qn_זR
�zq%��ݺ�zx���-'R|;hy3o/-��7����ba��i|nf]]BƎM�H����٬�+�H�)��r�Uy�d�X�w&�caaT��4��s,��	I�X����w�0)�գ��o�ԢlT��w-c��(RWI�V��s/�H�ݽ��_8���)4���ᔫg5t� f�?2��]��V��oϯ�#���K��ә3(���!Ȓ��`㥭[��:�u4�T�Ŵ���h9�2�d�J���Ƒl`�ĵ��.,���q�����54w�2���Ew�� iµ�Lk��D��3H�"�U�py�XzW��Uf�P/1�ԅon���xv�U�7A=��%A���ZP�0��q7bS�hvw��Y 
6xƠ���ܤ)�u`�z�t��.�h�)�U+>����utda��vI1V2cv������32��<�K�h�.�8�J��+��Ua�f��
�,A���'���h��0�vj���ʵ����H�e��U(�9����R�8Ud�5���L�.�m�+{>����z^*��'S+Mʛk1:����=w4�n����2��UK�`{d�&�m��*���X���MZ���4M�B����Wf�]tv��[���-�n��4s�Ǻj'�A4�*��B�:�MX�f�⚄��@^��f�+R�lWV(i�6��ۖ��ˌ���Hgslʎm�� �VulB��;�e��]�TU�Z�K������H��Y�c�+u�xE�z���w=,n�(=��+��^���tR+�t�L��2�0���x����� e��J	���k+BZD�� �t�U���H�d�����¬�qIyl�9����x�
Z�V����LnWv��UE�4���U	$�͗z�,�P��gr�r�em�*:����:��&,�P	C�ř�Y���j�ʒ�횄8�CEMe�72]��vhLq�i<3r9Vf��4�u�e��ܽ�V���6 �����&���.�)i�u��nɖ���S4�(�J��� Z���Y�5�c4d�����|�/l�n��MLی'E���-�!j�<S�=�8=m�tE2�����Q��,�Ǚ����z��(|����4�ڀ�Yב���ߝidS;�c,f�2V� �6V�hY`��m[ZEY�����jw�㙰+c
f�CrMu�]�[cn���Y�FE�SX�LfM��N�!=�d� :8���ۢ�"2n��
�R4�0K�܅���V��cl�5f�mba���U��H�ͽV_f�f��O.�{�*;t��K���n�U�[��0��ӻ�nȤ*���i��"Gh鶥<{�J���A��aWf��k����Y��N�$ �-�[��ѡ�YddM�;8�Y
賙zF�ڭͥ�V='�,f�S0�@�tq-�Kt&^��I��Ԇ�e��ĕU1�Hݸ��&�u�6x�����]:�׷���1�nc+�;�Ld�
j��AZM�9�T��6k�U�_7�X�e� �r�jߊ��O�/�j�]��-�����R:O�}�����t��+0M����X�V�c��D��a�E�貋�'i)miv���m=�U6�,��3K�����wRj�b�������.��cx�k�|²�V�ivC�4�К�e����J�% ��Ou	�Q�HVqX�@�\�d'�i�%��[���E�k�V�
/s%(]k��4'�)Kl�j�h�;z��v�哧s8q�A�6�����v��J��j���*��X]u�*�ߊח��6u�t�sRy`��mx(�x�AV��cC�y�*�vm�M�����X�@���xCʻA7GC4�;�ր����ŠÁ&؁�i����H�M��ءF�Os\�[�A����ֱze�,
��ݢ�,U�P(�%�sC��,��Z�yhP����Ѣ Q��jӤ�dP)�ek���n�T��b��%!>"R!�i���o۷{�mA�l�ׅn��D��
K-��hL�l^bd���6�Q ٰY�x��_\�3=`m_���wWq��HL��/�c�R�	`��8����$�e^) �kYZ�»�O1���Wp <%�pA�P���,=-b�1譅��F�$^'w��F^��GM�W�ۧ�lz���9tA�"�}Y�H�Me�]�+����(<�Q�K��n�˶ķu1զ�{�P�&��J�yw�ʫ6δ�@���,���,��P��qꊔ�b��Y�!�̊��e�4�40b�QRm����.��nM�!("$�{e2�``Y�Xv�L�jTz���e�p���W���&�[��F���SB�o6��z�f��Юe8I�/(<)Ջ]n;á���gko)��E1��3+e���ȝ��������-�P�ӂ<W#�S0d����r=	����t��e��n�oPF�0�v�'p*צ��i2�҈���W��7\��Y�Ӿ[�mm��k���/�D���i��%��۽�F�qk�
�w/M����)d�9�T�ݻ	��Av
�u����H�PǣF:{�$��4��N�T�a�N,�7�W���%ͬGP��L:G��+cF�Urk��1��{�o	E(u╪�K�,�8�5�2���%�6��& bh���	'GB���0�T��ؽ6.��ʸ���Lຘ�!u3&ִwwZkij���ې��c�Qo+�+[wP�v�4Tt�H8�����D"i��͛z��o&J���^h,mڭsUӸ�]�
�Y8�Qr`y�,Mߌn (�sl��-uy���lfM�ytWE�����j����{ٚU�������V���c l
٩�2n��M�1�6!Lm��ւ��	�[�+����ZL�WA3X�ijOy�,�0�DŻ۶�C<[7�41mܛ�aܑ�{� ]\�u^���+2��LIӊ�ފl��nRJ�l�FBUc�n�u ���v{ xHŭ��[��tS/tض���(��r	gE��{]pyC_[`����T/eD�o7-ԧ��&f��:@�n���@r�EW��I;��Q��a��U�+)}�*�WB���R���%6*�R�V�v3/fV|&m�G�j���ln��7Y{�����ɗ(�VI��_,�4,� ��Ί@�8�[t)����Cjm�^荻�x����h�o�R�#[K^ ݤ���yeM�4�ic7SKVc3(V���[l��{�$)��:�m�JTw�b;�VU,��̦���Ff��nv� �b�Y&��}xE�{�]u6PЖSf�5���P���Zܛ55�#���=!�6��/""�X�l�e��k,�An^�<C�"�|�lS$��ނb�cj�֭�
�S69�$t>˼v��ECYj�S�ݤoS���bB�PE����Vš�!A5�K�Q���Zٵ
g2���P
���)u���z����!m�c6��,�ЩK�`)f����U�a�
\u�f�D�Tu�E��5��U��.��v�+�kI�0��xE���w�꧲�X��T~	����1��Ǭ�/�s�	j����.��e�DaU��k[�s�m�J�s�c�z����&@�ժ���jax�.A�lm:ܢw2�ST�,����L/��ǔ����L�d=}���eo"Z�X��`1O���8m�	5v�t�т�7[B+�9[�XC�4�����n��X�VE��TE��Ij�	���Gc.��p�t�G��.5n�]�G,��2�%V�La�48�
��J�T蠘52����K ��o�3[U���1��b�v~u�J�^by�(�Z<�"�%[��ol�wwyʚ��-���Z�K+x��0ZPTܳ�
j���s%N L�vH��Y��&\[�3��$���Z��%�3o(h���х���"]6j�2�wu��se��x��0+ V�^�n��^���	clfcwo5�ebw���-�]�!j�M����te8����v��t2`�;��[M-#usJ����76�A��V-?03k/��7f��	��Ӌu���-˲���z�B�%]�A7rԻ�0]�D\ו`��
r�]��쫭NX�%�j��tn���ODŹ@�+e�H��O��V,��F�y0� ч7S�ur���qM�AM �֨ކ�+[	�*��Y��\C	f��ʖ8�37qJШ�+Ec1�BU���-����xD4�頾I��mſ��ޡ�evs��A���#���=9�� ��%�4�� ��b�Լ(�^z�cT�$)-��;��;�r�r�E��vM�_Z�-��]k����̬�j��c1�S)GN��&�&�߶�d�Z�T5e�t31@�#�{j��.�Lz���q��W��˫�2�ڱf��xoX�=R�f*�v�F�72(4`���
���}��̖B�Wɧ�%���Z)"�S��l�"��(�ѩ��e�2����.�<̇oI��wkcNغ�鿪$�Y�Vm�xA�(A,�V�V{j:��6��ۢ��k�h���������ɢ�2�eJ��zr�����l����:
�]:elf4��0�d.e`㧹���r˼��oB毞]e�b��]C�F��DN���b�<��V�y/4�@8�0��ќx����p��D�w���c^������N%4��r�;�l^(�����f-Ћ\w%쵔�5V�J��cy��b�PK]��g������X*]��vaE�dU�
T�����1v�V�1�rwQz9P<8�Qn�a��)9�f�u�3n��4�_�ج-����tEX�Z��IL7S�6����b1Ѽ8�����U��і�!�ل0㑓�%[���Z%�4tErT��r�&A/IRĄ���cx/v���\�lJ�}a��W���f"�9R���;W��wW��ʼ�*Z76�xs%�*��ԫ�ەb�B�s�����{[c(�7n��n��Ʌc$�T�:���V����ʺ��$��WV!�ѵ��l-Pն�����:-���8���rf��.�^Q��`6����E��RV1���j��aBmT�쫻0ĨIQ��\�m��E���P*}�q��{wNa�)���#F�Yz�q!�4��j�u+-��N�f��C묶�%��M�)�MVDz���t�V�Utt�D�.�av�@'�ZG{2�v�w�YՔ�
t�<ڷ�h��%��ַ�B�(�Mc�˫b�a6�����R����ڵ�y�2�G����)�F�����j� dC4��[XJ�LQ�y�i�ҥj�o/�kwy��L��:��熷���.�!]��8j]խkB{[g�����WH���w�-[�2VH��[��+v}����&���,eZuufVfRź���["JP�3e�wX,�{����0���n��D6��4�uVĸ�|(��x�Z�:3t4�1���l��"��Y� )��r�@]����-`�����_m��(K�m�����k��-��,㭥�I�ֱ�^QQ�w�2���ȥ�Ecsf�F�9M��{*�{-Mf�b�p���<;�h�6r�j�{z~�,�,d:����#�:��"�N$2�մ��hƉ�P�o�T�t��*K�l�I;�Z���m�v*Q��7J�)�&]�!��Y�^����'5
�,[�͝�E]��r�� ��ZO5��̿��e�Ќr�؀L�	��C�,�b*�3%����cv��I�$�f	���u�(�3���7�r£f6�kژlf�YAx60�5q�oj�'.3{us4嬚�ڗ�͕�&(�bu;O�.*�_ms�:
�O�(��]�/緎I'&�E�������c.��V��qn�P�1��v`��*)����R�-n� �r=�>Up��4� M��|e��R�����4�z4�uas.޵�]��y�V���y��hat\(����)���7"���+�Cen�9U���Շ;n�uܲ�����P ��/_bD�6�ޜ�L� ō��(3t2������M邲�
wv�*bJ�Ӓ�EM��Y�#G4Պc7J��@Tc*�
��5r��gU�3(�e��;�5d�F��/��=.�%�7󵃰]��mh�ۖ������o,�XP�E)��4+ �bZ�-˽M�������Ɠ�<GsT	�c��4�Z�z)�]����3��j`r�Rӵf�ۥ�03�������t���q�o��ExT�m�u��^�i����4�(J9��K��z��g�ye#�r����ŷhҪl������Ic@�Ov�զ7-�M�JN�~V�ŭ�|���vdic�8�5r��{��{�h����W��.�*۶u�QVf�m���]@3r�A���3�l��[��y�kƨ���[� hT0-Ϟ��Xtl����.f�f�˄JM�z*lP�iH�Ǌ%�IWX�'���f�V��ۻ�8�����n�t C(��ܝ��j��V4su*]�N�<�u����Eҫ-��p8JZ]�"�Uu��Z��	�%�Kެ�Ɗ�p%��^�.�DI�h18��D$�훰��7B[�]$��Ȭ0*��͏_#�͌SD���Vl�QKr�Bİ�Z�q���Ife��ڦm0n����4RG��o�;Uk���d<*�@J�m�Q3��$Z�ckY�����Va�#�u��b駵*Q����[;Z���Պ�h�O��#���O>o�s*JK�78�tMv���'
䘨�a�2!|���"�oJ/4��g�EV�g'�.�)X�(����[�y�����,�x�2�wk�+pZ�VR��;����f�#v�Jk8@J�lgX5��hqc���K�剚�j��̚��DJ���V�1޺��A*ݔJ�Ss]t�����v �(��T�XZ��N��[K���ms������=K5��"��7DQV������^7%p����˾cE7��@�ꩥ�6Z]B0u��n��;_-����◫yg��kᩛ�עtT�h�inB�o���JQ�%����_)mP����t��[O��eM�2���b�Ѽ�O]ن
��a�'n�!��z�K�tYW���یA��v����r��2`S���UugZgtwgҫ�M�T��7��ݒ��9����W����͖�;�Վ1I�LrH�Fٵ� �B�ʧ'mY�΀��(΂��%�!�@mm�+iP�V���Y��V�2���\����XQe}ǅ�G� b鼌�ŐVoҎ�+��GF�Ӎ��[��wR�(��y��7h�-
z{O��N7S�V'�rW��r�#at�n��S��ct���g~;�^�W^��ʑ�:M:8:'p���p�ǅS���;�rD����m�=��]M3vst'��EjˀK�5N6Mp��k���u�c��k%���8���]��f:�tE]l��)rι.�&a��"��-oS��b=��G�s����YTX}.ѫ�P�T�����j§�gi�A��v�2v������р��,�>jY֧u��*����m�ٙ��m�x��j�O>a�L_u� �Hj���G'2���Aj���yC��Jè�f?�ڦ5qux��A'gf�'F[mEZ��6�����k���{2:�t,�2�|`�'Cs2jL�+�f��s�.r�Q��BƲ�o3t3dF���:b�-#tK�S�Ϥ�k�;�d�1n������X��1�B���[�Y� �����y��T�RCWPˎhw���	�����ݼ����o�12K58�cAt���
���ab��ꕢK�+{j1���Co!�k��n�vh�-�k��yR��;�21Kw���i1�M8��k�\�te>��$)�yX�ӣ�H����k�Y4��j��q��X���rF�nB�1 f�8;帪l�L��H���t�Ɖ�w����Ggk�:d��8H�Y�i$�2)L:��sF���]B��Q��vi�DΙ[�zA����`�[�o�Q��`0Wi��vʁ�u��rwq�+gM�mD�b�I�$Z$Ǌ,�D����ە.�3hp��\&ﮍ�;n��A+4h��g^�~�[vU�Z�E���\w�:��;���c�Uo;���V6D䞇���"���ˉ�M�����o�q��V�(�_	ЉpY�`#�iT��a��(��Ӝ����ŏuv��:�y$ǡ�� 8�k��zۘo��C��[9�odbݘ,va�g���E�ӻ�H,��ӎ��>KH�-�P<5�-�`�5�����d町�B^�Y�4��熕4V.�ݚ�f.r��	���n��d�-�E�YoA�gE8Sfj��S�,���P��K�Csq�;}����V�1!ڕ!�.�7����}nje����;�W=�[�d�4n. ����chqfq��ֵ��o1��f�G�=���Ӝ���3A�vu0B��;�r���ǩL��`���	��J�4��Y��	�	dT�k�n^2�H�$��
��ԏP�����x�=�/�
���B�Y���̻Zem��X��rV�[`
�z�5,-S{�U��$�tx�����n�w{v�L�Uo�Yɉ���%��Ud!O嬼���e�}���K8n�LF3x�}8Jޫ�T�s��\��Z����}Rl*ʔM�x�r3X����e#�H�/���p�,�@��Z$<���7��ɗ�R�:e}̤5��MU�Qx��܉�7^=�u�w�d���P�a���'7�ݘ��rK�J和�[���|�m��l��5v:�\F��|��f�9R��\i�l�cI�Z��]]@$�<�f���킕�K��b��ᩎ��Y��m��.�Dũjѧ3k�b�.<(8H}j��#!�F�t��Ʃ�ɸH]��#/��]h'x�P�_B���n�e�[v����[�&��Z�����X
u�ܕq�a[������V.����:� ��-��X�g�Y�U@Fb���gB�V �ܪ�ɂ�jR	;�j�÷��`IؓrV�]fgqȺ�nS��v��M����z\ri˲�Hm�Ch[+cΧ��)�n�Mǚ�o.������<3�uR�N�;�^�d������\ұ�ҫ4�r|���r�>�-�e]�ɧ�BF֓|0ɺrzsGwu��]0oG_"{5��
t.�ŪMӧo1R��u���傷�BoTl�Y٠���^��/N萑{�%���r�j�C��*.�k��K��]سFV���e��ee���B���yv�YŚ�����g8�wAvh#*n����'}wЌ:��w5��u� A��\V�wwaNX�x���:k��L��Qy�9��J�3*hi�團��Z�8iޕ}�l�=���ʝBQ�Y,��dt:�;G^Ѡ��J㫗}2uk���ڻ6�C��̩���S�it�ӥ��B^���}� �#��B�+0'��_l�0Q	�P	A����/*�>�:���b�L����d��V�)8Xմ�S"NIm@Kk]�Ҁ^��`J��:ֽ��CkK�uq;��N����ʹ�GU�[�,���B�v�U�I��w��C۟E��j&v���c�;�*�8s�y�X�%���:���r\Dۺ���Vr\��yI[�AM�[5�i]��s�4-��p�r,����u����
2�\����SH�WC{/06��W��7nѐ�����N�4e	�`F�X���L�kb}H�μ�hAL�]����=0�L`����V��RZ�<�w�*��3���w�X���KkUꔵ�m��fwS�\p��j��F�в^�C�K�J[�/x�ښ�Y�z-��C4��@a�]����/o#ƆJE�J4�8tb�6F<	3��^Qj���z{LiM�(��^�}� �շ�� �K�5�nT���(۫���f����VRn�:�;YהUC�9P�yE�wY�W]����t�eҮf����F�˙}���7)�1����Z+�F�����K;�g3�c�]�&�u�΍��c��%��f�-�$�v�v;�"yZ�դi� N<SL�<s+%+����*t�����)v��V*���2x��s�-c�o����Θ�zy�m�y�C�����Xl9��L�[�*�c9RhXܓ�p��������1*"	p�wR�΍�M�F�]8#N.4�wa����p��w��XQů0R�U$��׎@�o`E-�r sT��p��8n�X��^RP���)Q���U���;̏�VMV���ˈ���;�	��X,U�R�t��֬U���]�5�wjt��RU�C�Sܸ0Va��}�)<7Y��u��4�3�6�,�o�<��ͼ��� ��c)��-�N(ؘ.�{�`}�N���rG;��l�����6�A�V��:�^])��a֜���u��v�d/����Gt�^-6D��K^ܶ���]Nm��Յ��76'�d2ί�E_E����c2��b��4n`@����ǎq�~�u��P֮�sͶ��9������t�Ms���<�w��k�"��U����[M�ׄ]AiS�#�0l^�?p���`_�Ýxhe��fI.�
�W���Bޕ��OL�E�#����t(=��.o+��1n����tL�����O(��RE>�C��g@ܩ�5�vh8L �p��ϟtO�}9�ph�Ӷ�){�nh��+T��HokAj����y����D��|t�r�a�>Z�]��6���;��z3lJY��Ƹ�T�%7zD��("�X�mZ�m�:�c�2��V��ܫ��4>�ӗ�&��5���ҝ�rd��Z�-u,=��7YC-�P�Ns��GD�:�n�F���������yh�C�Z^�l	͑��}��MQӰ����e���G�t��M����C0Xo�2��qe8��V�X�Μ"j�a�A��I�5�\�D5c�m,׬c��Q��J[}��Lf�'�̗9���Л��R�wQb��|t]=�t5�dÄ�oFm�jV�;YM-ߖ*�U���]&V�������B鞏4�(���s"͓ �nR�s�.���o�#E`��/f2����a���*��]�Π���3��b롑74����`�uJ��ݍF�Qe�	��o�&L��.��J�d�G��t�݋��P�|�\*�ԭ�o'o�^^�!ܤY�VhO�0�g�\�2.�/��M;z���Xp��+��e�e����|��I Ƌ�w�Y*d��ZhQBһĺͫ�d�#-ۇ0_T�>������6�&���.Ť(I�%���4J�ޫ$�+�+��e�^�ǭ��t�g3َ��M�B�oΗN��9|xeY/���e6�
�%P{N���V�w�1��{�Y.�_u�.�t��g���u�4����[��&Wh�mv��`�C��Zk6*�˾M�W5C�4wZJr%+���{I����U�؍s���8y���ډ���R���4'RQVk2�fP�X�:�1Wo6�xȾ9*�gͤ󄎛�;����*Օ�s����[���4 ����t��vcLo�}z]Lgh�!�v�j���p�4�mc�D�G�N����ü�U��K��.�FN0���[2oZ�em��R���M�����\78��PBJW�f�%��9v�R��TmS=��݈N�\� �L���l�ѥ�my�b�.Y�>:�uhP��E��Ӝ�;u���U�,�_u���O9��S��`ޕ�W���H�{������kv�����ɹ��-鲹�Q�;���a��61,��8������V(d���f��JUpX��J3�7xs��1?�э�V����[#���nD^�{�q< ��;��\
����,�
vtB>�F�WX�����J��S�Ƨ����[�o�R�]����X�+{
�R���IM���髄=��=x�'�mL�;@�bTF�P��`lx�՘�eM���)�8��R���������)l����q��H�_}�u�xDΆ7O&5|칊��-T�!?2���^�jn��ż&{��2�E }��k�[i�����$+z�1���$�zf!\ �<l�Ɲ<�����jѾ}j�����Y:f��X��텫�C9�1��x�ӋaE�f�4��3�ϡɮ'���(;�n�U������,Ϻ��d��t�)���װ�݈��J���x��&�kf��Ӥ��Z˧I^�B�S���=�u{�lM|*��`ܟKl��En����j��*�:.�w��ɓ9S��)D�K5�����;��:�bem�x���b��ւ���c��홡�5�Ln�2��ge\�8���7r����b�O���X�E�����3V�&�{���9M�k
��|��Z���F`���ۧ�d��Y�T
�7d�X����s����ḙ3�4�hs�=aڨ��Bkv�k軝����+;\�:r+�Th�8�9�+��k�R�7�67�ToREh�2����ҋ���Z6G�[jf�K:N^�C�.�m�Ϯ[�7\�jįw�_SS���0N������t,�<ثEm�+��K�c���/����zW�/F��n�,ky�8��m��[յǭ��9�u��B�ͪ��]� �uҙF�8jl��@��U��
�5�U�'Z��rjW<�GB���Kb��y`;��R�:mK�t:���|R��s2P�G)��^��e�F�Y�.���#�X�͜��IsO(���V����*[�V�J�F���}z��ؑW��f�txK�A˚�k���
����d<n�
����� �M��u�2���[q���-J}�l[%�{�*�g6�,D�6ˈ�[ضn\�z޴�u�]��0/,�.�S�� �ű9:3sd0R��g�=�Դ�B�d�2�nڰ����{��`���IF����4����ڀ��u%�]ghi�p��#��hћ��w��Q<���`є���`[Bl���DLu.�mTr ����w��TR^������kka��Q��-���Գn��;�o�5H�ٴ�$)׭5��j�5��/���R�h	�
�{��-*��]�"�7��u2���ž��[���	��8��N�u��w@�[��ɹD�Hg�_�-Y2*b�N �M=yt��w|�$*�m�J�6��C/k��Y�Yޭ%�
��L�I�ܵ��ʛ.�)o�V�]��j^��M2�۵�88�ٽl�N����^�I*z'9-�ޓ\�qˬn=�|��|b	ΣQ,֩:b��(����3a��̋�GJ۱Q=��,e�݉%�;z�Z�b�r���8LD�"rZ�kr���R��O�]�ׂ��(d��c�;�lt��b��z̫�Μ�F��:���U�e0��C�Wf���+Ef�����o�}fՅy�������C��͗SN��0V%e�[�ɂ�f|	ޝz��s� k0�bRxJ� jGRT�7�>��Y�f�(b�&!��F�Bf����5�^�t��RP�U-�$�ňP����0Ś�EG.�����JVZq���ud\pwN���KzOt�"��.(%(Y�o�m<s�����Hd�y�:�����HH~@ H�	@���v�?��9V�KO�%ݟ��0���TWjd
^<��'��E�=A��|K)�a�"��q��mh�p�y/NN��V�^'˫w�M)c)ڂ�hT�k(3�dûqji�C�m��J�r&�U��iPQ��1�N�a��4u*ܥҒU��L��A�3�p�[��p

�6�Z�:��r�K�4�����ܫ���8�ڹ.M3s�:��G(Z�"���9R�68(X.��ًv�_^^^�mZM��Љ��X��1�w�0�h�9�I8u
{9�ԺoM��yf�Ye�=�R�� ��tVa=�����)ˀ��,Z��g1���j���o�����Ji��"�]�'u�v�q��־-v�ԕ�\W}�u�{�f��=�ݢ���(��5���۔���Cd0VIfdK�h�2�G��^�Oz�_m�up��Ȩ*�J{��z�l0���[1+4��,t�8*3OW\�j^���l%ўww��t�A&E�@t�-_lA�#��2y=�n�������m�K���:�}2�}.�5�yko�U;���'fY�H}���ƀ%�[Ш��q��S��b�E�h_*����Aݻ����.�<��q��*�Pk�+Bݔ�Uʲ��'�\��h��.osU�{�I�髼�v�g{�Q�m��/c�"��0J�7i���̋�`ב�̭7UL��z�Ċ��TH%tN����`�iU����X÷M>�4�dwu�fj	Vs�d8]dPW0�1����͊��cK����(�泈^G��	^�T�g1�[��sR���2�S�l��;6Tyf��wvnt��׍�f�KY�C�;��YbA;������٥o�F�*�j��֪=j�Z|3D<a���;�F+��"�\����D���o���\��3��t; �R�>77���T�S6����ܖ�3�%�ɧ{��{��SiS%�P�Z�y#�
��[�8���5�� ���d���%����cEf�R�U��R����V�m����
p�̵�Q3�}YmڥM���.k��Qej��8���k=�)[Аf��R%&wSW,Ta�p��3'}u���v���Hh	>[�/K�.b-|�nR�[��L�2�\2�J
�%�Ԯ)Іi��s�/`�hT"��%��!�)���r�
:��7��q�f��i%��nL,_\�%�nN�e���\�2�]�M�*{��0�!�6�q40�|�+zy�|���,���9n�N�9��2���b�\�N�U���棾����t��Y�]C��Y�5F(0�3�2�[���=�>5�Բ�H���7�T�b^�n
����tm*�ʾ�M��I�G��j�ol%�\f�+k���m��x.���Z�Ŭ��n�5���\��x|�^�/�A:�<���C@��L `�V.���WJ�U�Bv4(���̾��j�n�]C���Hv�u���[9�f�P�k�Zx/���qc0��FS(����:��Ǹu�d�(m�i�dա ��xΛ-�YNFU:�Z��)��D�:��q`a8��Z5y�}�m�N]���w�v��fҧ8VLt��(A��7k��DQ�ɪ�R��"�}+f��]��V��f�ā���30���q^�f�ŖFכ�gX�L_6tgg^�{bԢ�2�8kNHPt${K���M*�J-˺��s�R���ϰs����<�IZ��>�v�pAy�^-8b�M�[)������}�Յ#�l鋕�o.�0]��-n����pK*23�q^S;)�xw8a5�s2�Ĥ<V�]�|�ŢH�^v��Ϧ���텒�b� =�8��1ʉ#yd��ٚ�%�l��jP�[>�Զ��\x��wֲ�<�q��K�����gc���uȷ]]�s۸���ݸ�w�Y���;t]k��ٓ`AMԥvB�r���(����W0�F�*�R���cc[��K���Zrc3d���E���C�(�ݝ��ek8��s�������*�o�p@���=0V��V�[���uf�U)V:(��i��{N[э�{һ��pRF��4�ؕYG:���+uZ㻷9;AXx/��$�T��[�KSA�&K�%��d7���ókM9Ƹ�����=��]�Ž��sN��N��o�n;=��rD>��w+��E\Rk�tp�*�A6ML)��;N����U�9@�g���Y��w)��t���1����U��nT��D7�6�alS���Vs`K�&ѶV�ѷV���؝�[�݈�X��Vl�ݔ���d�qf:AP�+��ݠ�f��yWD�b<^7Y+6Y�����`4�v'�:��"�l�3u�`=���R��g6�N$U�g#.P֠2�c��M��#���FG����D���e�B���F�����,�aB��Pja�lt��v���r5$ۻ���z��uj��ceJ����PH���;Le2�	\ȴ����#F؛3�M�L2}�1CE���iXE+_��U� 5g`ŏ�]�9��i��&�tL�-G;��ʝ�N�ѹ>*=��KS=�"׸�{�B���x�@o:�b�+f�
y;^h�N]L�Zc ���Eo(e��j�_��d�-���t��m��F�"��v�sa�ɮ|��+��)����1*�� ��ΚF�v��\����䐘A��F�1�F>�r��PbF+W\�,��o: i�;NC:���X�;���坍��/�av�"�
��+�U��\ϊ�r�g��'UJR�j����^
+p�n�v���dz&�ĝuCj+7��i�ڀ��I���[u���e�c{ ����r��Fd�H�uv�Y�I;uǱ���l�鐆�t�ˬ�9��J�����D�Y��L;���Ӵ{'��Y��G�ѥ:�+�q�Z���������na�6�|��<����F�Vu�1֮����
�z�&3��G�is2򦮙*�M�䲎S���Vpը<3p�JֲŲLu$|�VM	�Fa[F_���r�F*Îjai
;:�y|_Jiq�ӌr��!	0E#f���E�OP�[˧KӑQ�k�a��K����k U��T����5�En��:Ų8��ђ�n��YJ;��,+;Ye�؋/VJ����Wm�Y[Au#��s��	\���[�e>����Wr�qs�nYƺ䗵6p�[��"B)Mb;R�k:�f����n�9]�1�TWq3`;����ta{Y9eA2�2�)H@tu��^�M�����R��*���g7�_n�dy\�Z�WY[3�3;�]K�,���)M�*{���F<K+j�=��RG|�9���>-^b�e2^���nH�ݕp�\�`��H��Ǳ�{��%]'�o鮀�S�4�ʵ3Y��csBU����L��m�q�
ܾ�,����+pqZ2� �0��fց֕��_-T.uu�C �y��V&T��T���ũn�F��49�w��J���u����4r���H��F<*�q=�5v�Z1�J7k�!�����MM�b����v���-l�Jm`قAB󆇒��jϪ�@(r��.�(��5>5:��Į#j�&��;�5wq]Z�u��+��D�*��0��&sb�?a��NU��ۭ���Ƴ�\mp	:k{������������c��Z8�8��jC���o)�8�cu�AV ���a��}�,Vn&Iַd��p#�otVm�nuwz�P���a91���b�'6]��Pm��Lsp>�� N�-
3{�ᠩ`���	��9�Զ��:�d��|�l�.���0>=�;7z��k.ሊV�.`�K�+�Od��dϦ6Vp+��'d.�wbW�׼A�[0ݸ��v%������Q� h˃��v(rC���Oj������Wc{Y�2��&m0,Gy������tXe�ó-�ܲ��Ի�s�b8(uc��m�L�(�۩�2eḛ;�}S;�a8R%�Л�A��f���h`�K�r�%�j��x���d��w��:V�1�Ҫ骽S�r�2g�r�,gf;��b�w��.MDc���ȷQջoP+rұ��Ω��ڃ
%���3�q���F��N���yl�sk3�}�� �F��@#u7�B��v�����2ճ8�7��H����+*˳|pn8ú��ܤ��գ��b�Yӭsn�:JQ1��ݖ���fc�]�8��$匡1����W��V�5�sap7���2� �L{@�į�*���Ur�E�
|�S���|�܃�p��T��l'n�X	�<rn:��Zj�26o.r�G;F��'A^3���s����ؘ��"�a�r�I*ܓ.,�Gu[(v�2���<��9�����g!��mX��ka�hڭ��"��YL�$�MXŚ&�J�:2u�9V�-��}�K�M�9��,j�T@nٴ�2�7��l
��d�!�dɣ*���X
��WY|}�.<&�6%lZ�H��ݹv(�-�a��ݲ�S�.�|U`�����5��B�z�`S2�ƭ���\�۹9�	�1�Ņ��m']�D��^�K>��Vp�r>��Xi+�z�̫��YA<m�GYs����=�x'\2���)�Q��]tb��;Ei�����������^lQgG���m6�����sc��ΖX�3f��٦��Db��}i��N�^Ft,���wY�d�]��M�5.�oh���q�Z�CLH����t���fȎ"������B�x&7Y��vn�MLԺ���e��єC�c+q�L9ť���jl7��B,w�v�����+)������`ӻ��7#9.l��[u���ڰ܍�����X(�r�<�cٻ�t9�ͼ��mCN��Fԡ"��^�W���-:-RF����H�6	]�;[��CY
���AK�U���D e	:���o� ����fA\�#E;z��񤾾3�`�V�(惋7+(�pU{�N=��y�ˮ��$ck�TS�W{�~Ϋ/o`�m��
��.�9+�V'���l�gQZ�f�i��N���G}�D�z�ح3+^rGt����2^i�{:��f�^�&���f��iZ|�]�i.���N�ރA��Ȍ:<aP�PcW���Wsp�=�8����>#M�a����F��[n�����|V�L%wq��֛<�
�wP�}������VA���˸��9ݫ����̴N=k\�T��.3����[�f�Wc���`�8�N��M���S���/;��q��2��{]���[�gMgjE�N��8�4�����hV��1��6�5�з*"����,s��۾�bb�9Tsv���l�3A�e�_7F�\]ϑ̺ -�}�OW�I,����o�hP3::$M��I-ݩr��Ɖ���	YF-�yۛz����u��ޕ�n��wDڹl����]Z壌*�5ga�Z^�%S�u�qc�Տ/Q�̻+a��WR����
���Q�瓏4��:6ZkzDk(ؼLv��hur!�p��S�ɕ�l ]��xr��$���0 �ֽ�|wN��1�$3����W��nr<@i�`�'��EW�&����	��8)B@���ˬ������z����9A�o//�x�i��wq<�˒�CʹE�5_�v�z�vS�/Lv�qtU��h�8��TN3M�8d����	;�񃨱E�
��=�e��{�4{-ܘ�ނ=���,�̮��]@'v��!c�����$�9TuL��ۦjΣ*�'+a�2���{��L�w��N���Go3`�yB��ÛCZ�X�.�T��̛�Z��tF6 �h�yC��Ј㌬˘ye]���t*k�f^�/(���G�[�y}}`U�+
�:mXp�К��X�e�r�[y=�9y���ڴN��f��%nL�wd�����A����/�����ծ;��d6���ݥ�a���A��d��_6��ʋELvcϭn9�>'���`��@��E]j6,.o��6��J�6�]�-�0��q��s�����:���cU��3�*wc�].;W�K�����c�X&Ьt(5MP̼Ư��UE[����*�4w�{�VI�f������O�9D�-��>�<!���=�e��<Zoi��f�{i�j�xl0�Zc�Ǖ��v��a?3��zcǭ�xhpo�qCD��A=���fnGGL4��J�ǪCB�Pz�����e�ʸc�Պ)�G��ia��q�g#u,��r����k��a�0�N�(�Ok�)]�kr�AS��NTP[��0S��+%بk�i=�9X�e�j��'s�p�k�\�f)O�Cr�����.�g^�D���Vv�{ �됩��k��)��r�\ǡ�Q�D����r��4�}L*�Z�4���<"�R�g�AZ(�`����ւee\E���3�N�z�!V4��ҍgd�L4�4���X�\S�U��%�0�v�BЉ_wh�kr��hu_<��%����[IWxD�LkB�J��
��]!�G2m����f�;��i��tKv�dx�Z����b�)l��!�.�$">ۼՈ�`)��^��^�d�-*�ݭ�Y�E>U��{uv�Zy�>����i`
7�oT,�����3&���hn�u	=��M���Pk��^bەk�Eւ�R޹l� vV��R��q�oJٴ����65�|b��}�+Y�n͍��!ImJ��n��;V��L��+�t�Zx��ݔ�u�c�e_4�T^����B=z�DE1s�`�\:�"&�J�0N�5��h���`�Ҳe�*�hpڔ�B�nI����7��V�._T���^����Z\�8e�$ѫ�L�N��7HYB�;M�Rv���+}4c]��ѡ�m�K�����eZ	-�P���I��*�x�Z"ef���������=� �}0�P�z�������ד	D��R5�F��ǒ� zy�K�v��̳y�B�V�GmT�uj7���Z\�v�O�����+�M�5[$�M�i�㺺���r�����H��&�� �F^|�eS�.�JL���5�����q��{��j�"퇮��@����lw�b�F��WU�N[�����DYkP�s�D�c�Y���`lF�����F�}�2�V�T�;�E�!E7�im-�6�K�2dw�h���Ǯ�=�F��ew�u������3F��p�ܰ��	�{Z�>�ߖM1�4����W�����JsF�Р�u�m���	�E�1Dn]k@3�ꅜ/ge�73:�"�x�!N;����m������u�U��A�w����0Z��[����s6�s����`"`[��}���K�a�&�Y̾�����q#י9*��Ļ�`=N�.��B�R���(�*uC��̧��u���}����TQ���;\tw���K�a�KY�۶���o�ͪ�X`�!�Y��%�ZY�y���!��f_unp@Y܃P�ʻ8��E��vs m��7���Z��yӠ��!V���r,�Gnbש']��:�����k���&��>c�
j7����:�6���s󏋣:��vd�*Q���'*���z1=��!�FA^<�w����~�o������H߇�ofEj��5�z���<��\���t�y�e�KJ�����N�kX�l�֧���֮3��z'Y1�3�L��=={�����Ջ �{�or�"ʺ��[CE%9eP׽��,֓YK�jr���u�"֗\*s:�ՙ�*�ӵ9"�{�m{GNUh�N8Z�α{ӛ�gZՓU��WzX���z�
饝8�MM4֭*k\��Yٙ\XɭS'9��Lb����e��2�ՠ�.3J,as\rcV�8�p��ZصԫZ�M�
�CU��S�*r֚�kYb�eKS)�J�,�]r��Z�/7��H���ɽ�z���,#���&6�Z��ʵԔ٪h�R�5k:�Ze�΋g5��Q��T渴�&�fbU���X��uɪJ�s*����+q�R�[ZҮ�V5s9�%�U6Z�s�e�YREe+4egSA*5�ڶ����1)Ane.��6Exڐ�1�y��[��8�<�Y:�
��[�6�n�6��W�8;�"m	���&��XtLnuC����S�����wV�w�s���M}೩�������ߊ:�nIKݏQ=�8�l��ׄ������I+,r�H4WyM[D�5��[@���ǽ{6�H��j����W`t��r�ѻ�幋��97���J�9�wr���Z� ��^�ڬPsz�wn�Tf%���ZF��Pk�8vq5v%��!��*��Q<�:�+��SMNd���RDMj����m�<�Jhc�u�|�HS�lҨF]���u#�T�&��Vm�4��y����s�{�j�b��\D�o�W1��NWb-B�cA��;��f��[~Ͷ�;���}�޽��̳-�&���~��$h[CCq�KEk�Ƿ��gIa���(V�N[�i��h�B7���[��t���Md��3sҐ���,��5�\z�k�j��^�w���w��ξ~KE�>�Q��XbcN��C�s^ށ�c>��T/N^��Cb}�}�R�);�y\,_c�z���Ҩ��,���kV�B�p�+BU��>�CU�y�89��lw �J>�|�=������GSnH����!�=��.�����y��� �;�ej},�'��CZ�+
U�L�Κk<�Ǟv��䲋��y[H� �qW��M�H���U!bO+��UcU������i���d9;=="�[�968��Ť��0Y�,e��W{�X9�Xlk0U&V	���Y��L�7u��{d����J�S����>È�z�3W0b��۪�9&�Ss̾����n���!{�K	L�	j�	[��W3���T�%n��?\�S$�ڰs��j���/r�$4�{)f-b�#9��˶{^�i*��JO(-aieS,��8����!��c%�\V���Y���n�����s�����8(vq5v�����*��/*4Iǫ1�b+��,�2�fT�׀PW�p�b�����4-��A�.�ӗr"�¸�A�D`�aa����dk�����9��S�&Q��u�lv���1c/��3k�&�&V�M�'-���dW(��Q�J�YV��+�j}��!�Ӯ��p,F/0��cB��QN��FfuBsuRx	�\5rI#ڿ��ê�k���f�77�j������&��'m��`�s�g�^4w�㜦�үU��u��hf-�3^;p2������o5%�Ds����x��Ѩ�
�6k	�*��q��l�S��^�Y���%~;��4o������V��{^�Kj��F���Kn_;E+F�����6Pg&���y���os��6��y��W��vkK�i+Lp�J�V�ʖ{e���M�Nӷ:w��l������4v�QI��8Ċh�Q��2�%�i1�M�1iUsv�۳�+/!6Ih�*��\�14;`6�B}h�ƪ���x�9�S.��n�Y�c{�+�\���cQ�a�����:'�q�A���J�jS��K��4�"R˪d�u���a+���F2�w�/@�1+�ah�B�/j�4��vk6�E�����`h�Ć��1Ԅ�stE��hh����.�A>{k}����S���W��p^Wn�%{ʚm۱j�B�"ٔ5N�u�2;zj̻�n4��z1�����&ff�["c�s��w-=i�NW��8�X�&�^��7V�%�� �+L�ɉ�6��ӎT
rL�@c�bӮ�Q�Y��]"��!J6&-�9T�3m*8X�I�`l�1Br�
��.��6aF��X��HJr0z��:�y�S��l���W�r�Xo1&W-�A����lT�:x�@����̸��(�*�=u�!E��k4^�K7%I�\Z�~�X"m�QB, �M
 ᾿���-���\+��M*�+{S(Ti)�-e%qU1�<ӷ��T �x��)���e,�B��WH�.��QJ����pɮ�yxa�H�WR-Mj�e�p*��TZt�K&.��ix7�ұ��o�6��g�Ԯ[�8�c$y�V\��^��j�`^wf71�����y�_N��V���	p���!1oBG��2\�k�`�^��aX�F���mg�a�d`�U���0��^�k�����~���U���C4��F�>�݆������:���%`;;n1μ6b%*����sy�Ly���|�i�Äd�ו[���ӌz.�P�*���mR
N�y�8f\�'���޺X3UzY3�1��5=v
o�Ρռ��	����f��쭭[���\F0���C�[5��&qw:N�M̀w*bf#a�{�7C�8G�jv8Y�#Z2�1ȝD��K|3�OF�t��z�%eӎ�>�ݎ�[��d���VG����bja[U�qy�
:K��ͥ\
�}⎪�O�J�;��ru�+�VOM�j�u���n3Ψ���T�
�M�X��>6*��S=�e�{r���֛��#�*�\�r�#"ܮb��9�P�ݨ�.ddJ1]^"�:9���ͬ2�i�ͭ�\�"��'t�q=.T8���U�^�P	X�dt-I�{��n��D	���Kon�j����|=Q
gGէQC�PQ���q�=�^�צ~�`nTty_Us8�{Z�5� 坾����Ő���U]��@�n�:>| �tp�!�.\(Y7f����M�ޚ�巩-i+�������н�ki�������3O���+�|�O����h����v��OaY�U�\vK�8�.T���M�p���@����'aL�N�70�q|���z�N��*�zZ+��`WI�S�7ޟ6|:��|��o&?p��Ñ���w��Q�"�j�׾�BN���Wqxg���}�7�R��q75��UpW��(454)*��}ӓ�P���W��02o�<��S��L�pճG�t������:S�z��t=�!��o���yr���cv>��DԷE2��Tէ`�l��l���
r�`�CkJ��G5qWkV����3�Z��&j8�E��Y�V�3�v�<OK��׫Fh^9]t1�ۊ�����-�A�	t~��}��ٖV���ƛ�iW�,{қ���e��9Y�uw�
X��Z�obr��H�+i����Fv��=�P��~�WK�.��O�Ԫǂ�߬a�A���܊q7D��J�I^{B���5*3Al���ޚ�ͬ���wQB��ߍp�#l��69��yC;=mN&R�5Pe��0s�n[��x��}��X4_�V���t�/H\��3�fmM�Wt��<R�Ua9!ԨW�Un��b�UnV�����NE�ZptiJ�l?R�+�u�L�hR�L)[�$۴xyT\�����¶�pC/��������ŌX�X���§�<�boy�*�6�b�c��"HRp]+��A���5Wx��yߏY��О��3�^�ˉjX�G6yH{!��V�!���84ix���躬���*��w��Cl�	�4oE�d�P_E����x���`k��Mˋ��^��a/P���ח�t�7:�,��<���-��;�Ae{r�;;�AW��W��WFd��$��=gw�z�R��s*ȩ�{!�-�X���Ể���I�g:Q��$M�of�^�b��Ӵ�^^��(k�q�A�{ݖ&�i_L��픺���s#&�� {{�2f����T�%��j�Q�ٳ�c�^yg���;(>�q��>��������j�:5�j�0�����w([*�S&Y�](X-ᇔ�}���9�.�B�Mm�{S=y�'es�ei^D���憕R�	>'�jgpT�G�'adষ!Ήu�%UʼF���uy�d������Ȟ�m]��@s}n*,�n(1���S� N���F��e(�tJ��]Ř�1�5�&�v.�ПUp�S1NB�U���h���9�q�r�P�K��Se�_t����/�7u��{b���l��S`�B�
����lR���񝣽�AG�����։�F�� e�l1�Ӊ�r��W5	Utx7WK�$f)m�t�M���<��a4R�7/���Ø���a�v����t��Zڸ}�&(ϣ�����c���wos��Yǋ��qk�r�iptr�!��o�1��|����(�6�1.����9m��LKڃ>��kK�Z~=5�����'�`��w��s�E�A��˨QYUױ%{��!��9�D�G4A~7�؍6F2;z�6�U���zeQ7�KHb���쮾�R�D{wq�X�v��صnd���5J�2gi���gPzy�W��CUp�}��Z��m���S����e��Z�@���	��:��"����@ޕ�E���(9��Dۛ�H�B��f�z�(3T�5��g]����G�(4=$�˰�Ǯ�W��rke���k�K�#g��uU9|ONfYF�(������~��I�j���hO��Ln���L���Q����l����K���'�F��g)6��9&Lk���Z�`	�P����c]ʜm�T�'��Q�����D���X�%6�@��]N&�j¤h��*9&|ߝ`�ya<%�]��iR��w{K	o�Sk��L�!@z*�С�g����zs�}w#��|X�Q�cf�.j'��A֑)o��S�Bè�D��t��.D
���i��Y��|=~��{90z��,B9m�Q*hlk�����|���E}԰R%a��n���TLW�u�+{E�E�N_G&|]��Lr�sg�v�&P���@��� �@��B�D8I�/-�*�b���c��Y&���Q�C�0�f�t�O�B
y��[K���V8qn�7�SӅ���Oz9��#�'\4x��%8Fͻ]h�ҡ��:�ƼC�����{��k���,g�n�H�,2��p6�wRpn; ����\g��O�1�S��"నN���<���u���]h�Y���u�T\�h{�6��۵�3V�wf71��d�p)�_N��/���v �]'��)q�}~���s"�:��,b��Ӥb5�n�j���4�>�� �]!�Y���J��k[)�W)�n)�f���ϥ�������b�-㎎6��M+ߎیr+��0zvM�S�R�_���x��Y��Y*��U�?.)Z�o�9�K�D��eLfF�TT�p�23�=��8�a���c��1��<��S�&f�{H5�(U��Mk�5�J�+(�7Վe�9��-V�2(�zM�j��`c�n<Ml<7��Gn����ֺƐ��}0�H���f��Ew$�%["�B�gj��5�\2-��s1`�(Xڍs���XWD����c["�\Bתb\���P�CEX.��t�z\(��aņ�AU�^�+�dt-H؞��Y=}1��y-�H���.+ЦK���'.��Q������qz3��?^���0���Ƶ�5�ݨ�
=�v���k�[
E{�:)<{�7O�/R��g*�O����I-;f�d.���u#7.�2��ǎoJ����u�MU����y������ԉ59[��x��Eܤ�l�!��}��\��57��s{38�ƧD�:kY�C[����GjA5��=7������Z���`_���}�!�Ɍ�"�%c�ucy��&9B՜��c�=����qB��<��`ˉ�8/U��y���ZQ��p��jt�(�.T���M�p��~5K��Ԭs���i�%�3~��z4j�RF"e�����8ܕ3�H����͟�|!�%��a:?p�2��s��,����;�`��ǃ-��N���lz�����|��I	��3��k�8�x��g��t�\�+U������R˩��ݵ� ��#<]t1�ۊ����(�c��j7&KQî�Y�N_2��4�Ү
���o�
�Nv,S�}�x�����L�Ԏ�����d��u^�zr��A�`���u�U�t��E�]j�xI���YyY'?��ʞ���ݝ�d�y�'r�t:�[=����^���!��*�Dk����)v!��U�Z�8R�7"w�:_��1
3ܨ[��ӁoŽ�͎���'=��5b�o�GZ�w:f�_rU��������*z�P��0�79�V�jw�x�'"í8:4��.��3<r��sQs��8�;s�]��֣m��ĥ:e����U�����2�n��=N��Z���n����1�{8��
��Du+.�Z�|��X%Au/(˹*Δi�uX��.�a/J�9VE��g��kp�G�fp�A��޻R��<6/�["��n�*�!�>�0(,��Zk�W��fц��W�B�!���9�wX�[r�P�6��]y,f��� k�dYTk.r˳vh %��ıP�E𻮦#�Ʀ�yس^-w7N�E��;데c͎����W��W��#_AŹY�jS��jݧ.�i�Ģ���+��AkAq{���V�	��D։\*�c�Qb�d�|li�����l?�]���Nkx�?]ȵ8��B��j��IP��us [7+�$����4��7��i^���U�Sι��;������Z����jl�N=�a�g$�c()yr��`V��2'�sVϸ�k˻%d�)�2�:q�����-d�+�pYͥd�)�yv��jD�u�ivȺ��D-�.	�XS++&v�8�լ7ii4�i�qLz4�o��ծ�d�y�nFhPCQO&v�L\��e0�[�t��U� �k���ь>u������5�r�tusκ[h@���m�d���풬�m�[t%��e.ڹ���e�)y�@��̮�B�ۮ�9vS	c�#�Ð儲�^S���O#�	�z񴸜�iL���z]�-a0K+Y�i����ܺ\��mcn�����j��pН����*�� 5o�H#zLl��MaL�YC�|���q�d˚[�Z�S�4)IZ���v��AY��(D�v�A��p�P��ked��yO��,��<v��i����;��MlE"p�z�.Y]3�r� ������j+��w�I��(�G�V����}�� ���3;��<�Z�SV�?n�;��[^��\��k��3i-�	z���g���O��>��\�9wSJX��Y+n�VpUp�N�z�Ř_i������P�����ı�6��-$�w������GF:I��|�JȮ�����Wg\22�T@���N��5��ʔ�}	���8D[�*j�f��N�:�]f�BV��f�L՜�h�6GoP%��I\n0�Y{1�v��
u����X���5���k7|S����SI��Ms=�Y�}J�f�~n"��s��s�	���E��w/	���PL{q���0MP���T�wi<B��ԘM�+���-^��}7͉�M��^�Ri-��.F�	�+p� �U����t<���v��ob���l�����S;Y�`���x�$��-��z>��ʰ����6��Y�����uzKV�f�+h��+f���l̙X3����ǜ�-R����J젷ᶲ
F�O�@*SV^BL��v���o7ɤ��Eؐ�@f`x56���EF b�m�k&,��K/�ʷl��]^[�w�8q����}|����w�h��5P�i��9��Ϭ���;�J�]��d�8,�֤�TU�Za�t��j��S.�RsVMhl�6m3RT�J�cR�R�6�٩ej�:�i��Uu���#�l�L[���V����)��cD�fv��,�c4�U�`ld5"kkUz���N�%�$�kδ����WW:qkK0�4f
Iv����T����VU���2�&�Ʋ�k-jֲ�M�:�"ƕ�Y���7Z���H�Z�S5���S��y�oq�M3d�Q4֑�Fd%���V�Z��Ç&\K �6��F��.�4٬͝5�2�p-5�{y�L�km\:ΙgYK])�J�M�*�͘�l;��U�N�̧5Yʵ�ٖ���AWY5�uU�1�n�v�rv�	ffN^_�E�ē]�w�	�M�q��z����w�բ�%.��R�)�l.����4uYλ�}+5�I��$*�Q����F�Zb�8����1�UJ'����J���8|&b���,b��ǒ�c`E9F�)�ȣIsF�+%��8����c���a�ˠ�xb���E�4��w�V/R3;=K�-�ORQq�,&����́�C�Ea;VF�����KŮ�E�סּ�����V��AE��﫧}�f�	}3]���8ʑ�@q+��fX��]�2E#Q{���7��Fw.v���k ɲ�G*�"�-�0����'}�����j-j��8�
��kI0�e�M�)Q1�qu5���V0¥ ��I��K�*��f��ϰ7w���A�ݭ��o �V��ݻ�7=��pD@�}�|�seE�z[��\ʥ�)�W&�܆ia4�6��<dOw���9�>��8�2���(Վ�U��	��8h�˳ȇ�a"�1���}���nQ�=t�m��t��M�Q�*�Wą�]t������\���6�ms��Ċ��2����/ɫ���{b��ɭ�qu6��"nϼn��]U]{Q�6 ��S�=^�+j�H�W�弶F��_n�=8i�|�u��=m��"��i��wvc��>�o�'�X�_�T�5�oJھǘrF]ag�
pP�z�j�*�`Gyjl�q�}z-q
\R-�y��8Wt}���*=�Y'�mV���.e<I"nEy�~�O�	o\�����O/�<����,���e���}��̓��u�,���kԭ��K��A�-Y�W*�#�s8#�WKb����u��v�m�^�3Aٞ�����3��]<�������=C�6���zr-��1��Y�NU�uhװ7Sǧ<ۗ��E$Ȯ���>cf��m[�����p�f|�lM9l'n1�˕�V�ɜ��K�kd�����#4�
�@��c�su"�	t`.�=Ki����X�j���^g7���~ZU�_K�j�J�_�J8�?`�4}�7~n����Yԫ�#����Br^>��<䇷�=Uʰ�}ল��1^W�����l�0ciVzg�h^0����2i�E��|	�nv�ZOk/�K�Pz&>�&�e
�R���L��B�m�yR�8�ٻ��u-����W�b����p$�S�`v�*F��r�S�e�ǀ��:�������,D=[���d�z��qGN��J�ގ�*$B���^���ߺM�Q�j���ν�Rx*n�o"q�˽�a�[E�����x�����PGJ�kZ�FA=e�:�%�F�dmϳ�ި��:B�!t�5s�,��e�B�Ȱ%�s
;��[.�bK�n�s#R���}�lCܦ��Y��t����u����\��g�'^3&�ޭƸR�Y��9
�����t�~���+�@�.D@��=,ˌ�(��]8��<��sp��9��HZ0���QOԎy�6"K�! �M+�P���[v!�B���ÛvD͎1D��(�I��,C���;��<� ��w��P⑛G�YK8�_�
lFVl�A�݋��{_"�'.^�b�۶1�q��p*�6��Ӥ:^��Q�/�zk�S��In��B.��-(��ttMeq���~ݯnj��^��s�������7�SR�	X���rv8<�-ں�wJ�䳧H��78�+�7����B�І��*��+��t��q�LW�1L)�u
�����X}�����*�uO��u^��JAԐn�~h�RU�rs�~�	�c
�W�^Uc��|�xO%��/؆WKZxDȤ�V�`��p3ϝ�睬q���A���S�fM���{f[�8�D ��-(.�),%T�a*�:E9ozl[U����[��<.�k�v�堧Z�;=���1 "�V�d�}��z�[��2T���z�����Qc��3T�"ҁ��y��3�1��9k�ރv�A$ {ޠl;�����`�*����I���lo#r�ܮ���õϥ��j; #�!{l�Mwdh�I ��v3�
�N�2��].�M��&��w�cP	�:���f1A��vi\�R�3"ܬŌ\�(Iݨ�:�Ĭ�;R']��yq���k�t��k�xvSUO�1xpBk�IU�^�+�d��h�9��ʙ��{�[��V;n��B��h�q��d(�v�4~{�8�ϯL�w�g�G]����}���*�(��lyװ�	��G&��8�D���t�ypcI�±��:���ȩ����+7E����ɻuЈL���н�ki��%E/O)�S\_�Dt��������+ET,a�r�0��.��[N\�y���5#\�HK������)�ӵ��h�i�4_L�/�0��W����%T��9�)��y�K�2\`�Z&lW���x������w����C���Ǒ^��ӛ����s5/O�˩���(eb�8U>�ZI(�~�b�ȳ�U��5�>�����A���Խ�<F롎���;��G��WX�����gr�T��*��n��pBŏzSXRs�,��<{<Ƀ&�uw��*n�NE�XG�겐;��A����^64�9ڽY4>��|��03�cK�h�Wt�#p�;մ}��=�%g�����?]&l�p=|`z]�j�L��F���w�:�q?aU��G[*�4���C��df^�G�n���&9ֵ%�4D��n�m��}f�1�_MZV2f�	�״Ss~����Ä��mi��l�e�O%g�Eo����y6��-;-�g��٨�6�f�t:�U������O������7'�*��&6��(��9�HB��*����z�U��U��X	�|5�(J������j܃�Mr|j#�����P�3JK;�<v�n���۠�#�����~��v��Ok��V�b}D���Tj�n��r����j��8O`����Eƛ����0�X�������%'�C��uب�!9��P�H_(z&'��p*c�z��a�(��lr�y:d��3��B]H�7IX��-�����fӜ����.;a�`�~fk������Ust�*@p���LBA�z�DώV�`��<��L���2���ʵȨ�lهv�ħh�5��9����+%�ŧ�W���%w+ ��I�SF]s��eځ��Re�.T�wИ�}��詪#�#T��u̝`iMf+&���nW1K���`���˘2L!�� ��������q��')m��nCúO�݌�d|����Qj��}�,	,���Σ8*�[q^	О��H����sU�;`11�WTU�K]����������0{&W.�#D�O�j 8��<顥T��Bp�Ʀp�J�Gƶw�p�R1e�5�s�􈤗8��8*��7�kP񢲼�j�Y��x�Y/Ӆ���M�7�{F_U���%+�鎹iךB�C�6�u6��xN���r
��������cE�9)��w���=�zh�L*��j�,'^ذ�^M`�qu7����S9�3TI緇��CI摛��]�`�3�F�nK�'N&(=���_�d�L��*-�^�'M+;�~���o/��!����Ί��d����`��'Ke��ʸ>}�&)�q��x��,��8�U�����ڃ*,V��[s�yN��!�!��r-�y�>7��n�Ǟ��lV��MK4�E`��8�t������<8]b_pw����8�4T[RU��E	*
�\h0�N`��y`;)}b�*���Ѥ<מ����,%���� ��<�)�%��ڍ��My��b�M[�k������LD��x��������5�!v��3ԓx��+�\Q�Uّh���W)��M?Um������\3�%���0��x�0��L�}p�\�a3�aF�m�fc<۴��x�����J�3{A�NZ��s�O��@q�Ygj��N�j́8J��j|Gb9���]_���fou�-�rU�6�pj�n���
5��~�p�]/D��U�g�h^�uFЀ�Zr�T�e�ܴ�B�l�!�.��9P8a��=ʵ���(X9ڙ���y�}R���C����E�RV����*�Q�j�]�Oq�ǅs�t:���']2�ZΈ��QS�i����4o �����+���W�
;���cx���HJr_%-Z�ۦ,�V�-i+�r����6�;�yWQ�-�]��O��Mg��,,0M���A0���B����o�R������It�p:����]v!�:�]rt����^Dʦ���b*�D��EZS��(����nN����HFC�t �(��tUt�����;R�zϘޕ��ץNgN@���dث����6�\�a�YQi�,@��9פw����M�Fz��_V�EF=���ե:.w��k�/��NcsY��8p:�uY�>��7Ӆ��O o���7}CC�8T�"�#��MX���`�^O�[*��\�$B.e��1�.����7<ݣV�f�e#Wy}V�{l���v޴���Q�����F�4�ͨpQV1��1ʒS;�.-w[���\YY[��(�I��ݘ��=|;.�]vkV��ohDeGCa�H�G��v��-�_8�eHb��5�ϼ�u�)S���Փ�[Y ��M|����-�ԍ��U�����F{N!�.-oD
9۫�I椯4�v/�6c��i�� ~���ˊV�'[!�FH���]�}�˜,��jL?�����O��㵂�|s��Y�Fv:e� (7�@X\�J�ӑKy9EPΛ2��V�� ��8o=�bڭM���j�ey*�57��;�A�{tVғN{<|ұ�𪍟Dp���h���.��b�,	�P�ݨ�3S����)��\��{ܒ��8�"�:.��`�}j�W���γn�Z��T�U'�����7�t��Z�S#�V0�yS���֡�A\w)�<Ү,��S���E�󨾡}|w:_�Hd��܍�m��1a94���`W�\%T+�쾵���&G�3���^~N=�}o���C����B��hfEd�[BDQ`�4Ί�r�������WW!0�;c3�U��(�S��
3%��b�̓�n��r!",�3=�0&Ҽ�f4#�ln�Vj��V��ܠ��7D����`��M@)tE4����Gp��^����[��]�����bA�V$xu5$t�FA3�;L���3݊K,���O���AEի"�8�* 0o���4"��L���_W��^��4�f��UF�S�0�����ζ��
�#�S�)ߪ�	u�g�J���	ECݶ�SٱO��zaȠ&���]B�݊Zo#�]�M��O.�ߝY��ƹ�;���в�X`�K�O���5�-#�y�B_�J���9�}W�ήT��z�Y��-�a�߂��x̯yL*Uj��<i��\�cލ�a}"�_��$@���w4y���-��1lq�bV�f �۱oo�c45xJ|��uYG�R��Z0S� n�[��(���s �(�ZT?w�����y�6n�}�Z�WY��,��j��x�j����>�x���\�tV�T�e����=�HC��*x:p-���ٱ�l�y�,���2�K|�YC��^z�h��=T�b~5�O�ۢGP�8M9E;�A9zto_n����4p�r��v��`��X����/�>����
�V��阧-���(�w��ּI(�Cy��=jLb�U]{<l��c��$KrjB�Vbb��b��U�\ �fϬ�6�,z'p%S�q�,˷b;��_z�������'d��Ver�3w4���>��n_�P����a%�4J �Dfۨ��
�rl�uD9g(۽%>�e,��Q�t�P��f2����o�)%��o>�<�|����[1Cu�������*qt>K2Et���/e�E��f,���+�U�>ʴ0��<.��bf{\S��(ju��w�TJ�Kn5eJ��_��%��7�vv�t�*F�����V�IyݧV�(V#���joz��;ʵȨ�hûw�*��f��:���?Bo�8����<�"�p��0���u{6(�aҁ�z�Z�QO�������ִ]�F��Џ ��{���">��F�R�*�\*��"0�q;3��e-�S=t���e�&`n YH�7ú]>܃0�J�A5
D�t�j�X�U劈�<�=��v�ں��O%e*���LS�<�z�B�í^��E�Q�(_�v%�h	q�*�+GM���y,��=�y�zҗ��E16ں�N�����t������t��`�������C��{��@l��#u\7:Y��:q1A�_@��W�1S)^�U򻫨j�Μ�l�'���U�#�`��υI���a�:�����'k�=�"�������v�R�2�-�u� ����E�]N����ǛN���������ur]�i٪�{͒Q�\.�.s~�KM �gQ���j򯸰,��p��Բa1���),�Y��'*8uiK;���jk�ylK��.cw\ػ\��f��d��R:�N���,LkN!���-�-�������n�:@���7Y@�U
k��Y�V�a�1���#�F�����\�]S��1h���l�6�h#��l�h�4ﲖպҰ
�ф���R�%�0��ձ�ft����|�A��^͂V�MH��/�!Q����w����׼��e=��b9��;]J�r���6�m��"rYMZ�W��5T��v�.�v�b�1h�z��ƑVس���cr��BV�,�}�����G{T7�ݳQ�\*���V��o�
�G�Pӏ,ෳ���ׯ^=���Muk]ܳ��>�̡P�p����Qt�:��j�Vrg�b娖���!� r��ԬU�Fm���t��XW�p����ۋ^��z��Cm����37�(���W�����^�ʕ3�^h����9b�+SW����2r%:���ٛF�>YܐU��n��;ޱ��u����r�+`�Rs�+y#����#��"��.�7%K�ows��V�l*��H���*���o����yr4M5�\i7rԸ�S;��f�-���[��s�	,r�.b�n�+�퀷3iv�>c����(���ln���
�kq�ذ����2�� �Yf.�;���.vv��Y�n��v@:�QK9:�JF��B�� �JS���U��Y$����jh^\��}����쫚��aP;��%kv��/Z��6�{y���ٙ��<B��n�4յ2����RwVn+���c�nw)"���͐�M_��oU�ǻk�&��ַ�F�x�1���
�Y��_b���Xy��p|����� I��hOo��`G��|5����#o2P�U�*�]e��Y<q���|^�]z�س�\�z��o��l�B�I�3�5��uرAZr����9V:m`�K�EV�OD zE*����]�J���iu�Zauw��-���*�$��)���\�{�*��e��|��F*�.���i,B�8X19�m^&hT��i�۶������� �,Ѭ��v!p��I������CE%�{���J��'_7RK����	�M����D�(�;h�s�{Nv xt\^U�8*�5�12=R���`dj���Ks��7��g�z^ҽo��MN-����Y�7�K��%yۻ�qs1�bN���[e�VF*k����r(���˧�vv�����ں���8�>�m4 ��3]r��	�TCP�=�wTw��khg+����)h������q����Q��v5� ��r�Vuuᓺs��6�~���'�>4m�:��H�MV+��V(�+Y+5SB��:��.��V��fM5����W�mkcT��e���C�U2r�[Dᐃ��u�Κ,*̹�5Q�5N�Zհ�f��YԨ�-2ٯ{ݱ�{���YmW$Z��a��u-%��@�n��T�&�WR��-
�Ъ�R�BUYeJ\d��]jV����l���r�����s;+j��SI.���R�(�#4�cb�9ٍ� �L3ԗ06r��b�c7K6*a�͙G���L�iM5�jv�;;&�KU�b�cٙ�sE3+e8��0��v���KU��t�ojqL�T��a�0�����k]�t�S���޺�]Z�8`ff�z�oc�k�N�jf�T2��E�m�G�J�T�/V�{X�nk��Ȯ�69�Vl��f�dW3�Np�2h��\hԭ)��;�fU�͆sn��&�Z�fl��a���������?___�z!�`M�c΋��A�Ro/�C!�{_�v�wyz�f*����&��;N�/�m\49=}J����k�� �ç��h�*�+�W�G
C*��V��[s�w췞�a�!��LC�R)�u!HW��<��U<��(���N���+b~�?�^����������ON�1nfI{ƭo%����v��N��ӝ�؞>�l	�[�jlT��t���rg����O٦���_���aHzwL�d�Y�>���@Q|�����Ri��C�Ǩ�0�U��sO��h�-�I��a)N�`SL��~B���1B�|>�|*����q��_p��*RU���)�*KE ��s��B�5>��j�Y=����v�JHv��߭d��u��zÎ�
N:=�N�m�Q
������ԖͲSwT�qd�6/���VS����ֲ������4��^�@�*�k��R-����-�aH�35�����B�����0�S����u)���̽Kd���hq%9`T�
�3��ɯ��?vj�|�2<c޺7UB�y�2���(��)�dɌX
�N�LY��6�!�\1�!L-�����3�i��٦KC�R,�g�&6�Cɍ�I�%%��dʨ]�5��G�(�Q�P �)��\8�Y�*KC]݆a��a�[I�)��jꅓm��
L∥�d�YԶ���E��H)0�>��2m��!L�o�|�ڢy<��;�PMA��_|k䔥�0<��{`M�- �6��ݰä) �Sް�i�بZR���i �
í��H�����èZ���=��SS50�II3�1:�H
)ͷ�gj�.���f����j���*�G�)���'[��z̰�
|�����VAgY)�g�sT)&g�a��VR�y�3�!L0�S��,<�H,�hP�6I��a��!�r�ܸ�w�ǣ\��
?D�`�r_e*(�k#���T}�ٍ��D�u#��0�M�jq�����sZ����9����fSU�>��"�a�9�)�WU�B1�qL��rֈ�R;u�ݛ.]˻ʈa��e��K}np XƔ�qW7%b�G���ɼY�fH� ���h���}�7��A��Z~��R�!����e�y��>��"�RS�~�pKB��O_,���2��)�Mc:�Q4�3�4�0����+�B�a��6�
����ܼ!�<����g��3�9~��Ih1E�,>KChR-�)��Rg�y�T��e:��0���O!LתKOW���0��3=��I�)�'}s�d�l<��,%:d�Y�ǻ�Ӹ��1�����ǝ�H
-��)���	��qRi���&(2Ù�u<�ϳR[>I��d��0�A``ν��^�I5�*L�X{�JM��i��Ϋ+�)q�L�_���xڎ����b֒���)��i�n�ƪm��j�p��2`�F�u���˲�>m �SHa4���P��C>aO�2}�pi �l���zĞ�
Af�RZN�)!��!��b�k?vΖ�|�	��g�}ygXq- �+ve�C��"�wD�0��0��L�T-�u� |��>�Io�̖�&*Z(|����*a&��y�:�}��l)�h����Cl_ѓ��ܖKKr~���y�S:�w�@URy2s�2�Re�m�}a���4{צy4�l�ZM�,)�a��0�9�ZAd�Rq��uA��,Y��d�+��O!L�>�4��bɉ�P߾�Op�G�@�����q��B�}u�'[a�o�a)O�)�s��@Qz��nM$���9���V�{�e��9tL'Rߦ���-�1��R
G]���<����a��������DlxD�*��Ka�T-1tM�:�}�`�z�H�jn�(y%>a�57y�5<��Q��\��|��بw<�H�1�N2|�A����C)�L7ʟ2-Gv��>��R��eg��ǁ�	���C�H,���2v�R�����C�%n�S�����2����xf��-�aH�ܻa��f�JH9�u6w�4�::����}�*�������٣}�$m|@��@���'���P�%6�{P�M�L�9C��
a��,<��<�3��ɄU%��
Jf��S0�Q
u����fR����0Ϙy-2����#O��*.7n��r{jP7�KI�=쇑}m]���_����̼f�������r�v�o����y,�ד��)��:��'k4�j`����; �jN�&�U�꼛}�S&=��YM,B�ϰv�.�+$�k;J\�s�������ȤN';XC�- ��,�q����.y2��)���H,)��1e2m��B��T��N�Ø�Z�2]г���]��1'�I��;Y���a������p=�Y*��@����b�.<6<�:�}�^�<�ͺ;w�Ik��`��2d9�����ҫ	I:��S�R[�0��-$��:�f�Rjm��&��U����;������a��n�M��L�r��N2���d�9�|���;a��I�ku2i��sW �aa��I/t�=��c�/��_L�Y�\��z������жi���,��l)1��u�T57}�2�:57��!Ĕ�:�N{0�RS�Կ\���S<��3�!L8���e�a�n��)~�̖�b �T�+��}�r(�@�����\0�
�@��S6��l�Zo4��y-n�i�[��2���ZC}��)�0�ai���I��B��Q�}p�Aa�f_���&�I�+�������V�����w�s���3�Km�>��0���2]
,�% Y�-�N%��0��Ri��$���D�k�y2�Y��;�1��!I7ʓ�/����]H Tx|d;�O}Y,?��9_9�s=�.�:�$�ZC�~�&�%;`S4W.JCI)�0n��Rja�g(sP�
@�R�>��d�}1RZy���d1Ai2�&�2kמ�
a���\���#���Ww?/��"x��ڽ1��9��9�8ᓩl���a ��g}yC�+B�'}s��Y�Ka�޸a�fжa���\�,�<�����E�aL0UO���%>O��rF@���zb�<���N���ܲo���|��4�3���I�퐦u��e�a�n��wՆm��
�����e ��}fY�L>aZ�>�ne��Ķf]v��Y�����Ii�ꅖ��@��F��~���i�K�.*߷ڒ��)�(�$��k^ęH,2k��2�d�i8�9���O6�s��eIOS��E�d����d�[�U���������ǅT�����;�#�Kut�#&�1���T�w�Sm���(:N��Ϛ��vR�����
���O ��u��݇�4#���|�fS�("��7�{�N����v͗�-S�t�uh�Xl��fV�	�oAvx�Ud���3��k9+������+�Vҿ�@�e�иI��R��Ƙ/P��(����؆�m-WE����2Rt�q�
IO�^��!I5<�{V�����{�2��T�$�WBϮ̹��:m$RO�p"D����q
KC����!��dǨ�AO��L9d�Сi) ����(y%r�|mê�3�:���نygS��̢�Xy�/�)18&�lc����%���@P�*�Ǳ��l4�6��:�Ci)�q��PP�,�i�I4�8�'��!Hfb����tMLz��% .y�0���S'ݰ�<釘W��3l��FͺŽ�,Ef1��Զ'�z��Af�q=��y
E �]Ì�4�B�h�.�ILYi�h�@�RKB�f�u&Y��XZy�ͤ�l0�{BɃ]����0 ���!��*~�⦺�ĥ���p,�%!�|��/<�ɿT��C�Ru+�UD)�r��h6��H,�{ް�%"ɯ]Ł��/P�Wd�Kf&�~�a)&��fb�l⧦>�z~S1�&�|���᜾2�V�@�P�����C)�fo��O}P�
I��l�2��T�Mg���'u�\$��MB�p�wD)�3�\��O�F���%:d�Ц��Rks�0Ӽ)̭r��*�����VjKe�ʡL��S�9�2�!l�T-��y��	�:��vo�cꇘZ,�
q꓉�8��&{�bM (���}a�l
I�j�t�2}x���}5	��S�\��~C��>k��(���e��r�f�)�J�M�I�%3���
���g�l3�\�e �L5����)��}�$�)'P�}9��)�4�u�Xi��p4�q��Q_9X�kOw�G�#�g��]}A�M2a�<z���n�v��XR���4�H�����Q]�y-�ZJCwRgU/�B�e���Ղy<��SS}�I�)4��ଇ	}<%��n|�~IR��G�Ƙ.�Ӿ�)����!ϪJI�|_�L3�IM��Z)
C\�0��n��Of���f(2�H}U:�K�PS̖gw����Q��^,֤52D�����5�8��K�ŭ6�-�>ʾ%���Y�ܾ7qfD�o�=��v��w+Ǖ�ؘ�/VԵ)�Ư�f{菇��?V��U���lCy�$h.�#F��1me=z^��U8��StV�5ѧ�Q;��v7ycBY7�x��{H�����{wGrE�H������0�}U,)�&{F5�\�-���z���c��;��2��W��|�S-�y�2�Y�a�E�"�Y�t,->C�ZL��P�E�B��^�EM�����C��i� `�鏤��$�13�`�t���u��e�d���}�ZS0�����:�Y�Ja��\ªO��L�z�e�m�kx�S�	l��y0�Y���z�˼�X�UcY��o�k���C�)
Jd�)�h[�5�RS`5�:�(%$�_wlתK@]M���,)<��ߎz��2�}B�����0�Ƀ�^�.�)e&�v����܏��|�8UW|�\�ϊQ���*����,�Q
a��7Q��䴆L]ͤ�i4��4b��Za����ITf��a�T-)'݅r�S:�)�d����P�d�2��ж6"j��
���җ}��eφG���׽�e!uSRZ�S�m ��kS'��!I�>a�̚�a񚅳l��&��dR
C&����C�+�>7ۓ,<�S<�W53��ǻ�oW�s~ַ���w|+�R�8�'sFY��A}�Xu�S�6���9�i���;����H[n��y��SP��
B�H[<���ɳ50�l)�a�������S:�I��Gj߯m�8���������ҪM�L5ʅ��:�3�����g��T:�&9�}�q4�ФR{���)M�&(R�%1o)�@�)�Сl�jKI��-aI�M;����W}�w_o����׭'�RA��ܜrÌ)sL�d�Y�7U-E�'S���Ri��f}D)�_\9�&��h��3�8�L%#��`SL��������>���������
S�iI:�f��Y�INr��)�L=a�-�\�y��Ob��9UhJHr��ZɄ�>���y�\�u�m��}.ۇTt{��\y�muW-�����Ȯ�ޘ�d���5Q�
A@��I�e!�����yP�jk�&R-���[<`o\�0�
N!�-Ѿ�}P�E5�Z�JC���s/R���.�m�z����n�cN4�E��oM@�(w	y��1�Vz�J*	��`g���WS���=WZ�	�m<#X8�j+��mp��_�b��z9��"�TtJ*��$S��%��4�O.��2u.�]Ӯ���Y�l�W�D0U��*��W&�+^g"l�������I|Ƶ���9�sx��Jr����,8�Y�L_nP�aL�0v�qD�βd�,U'P�,�Jg�a|�_(�0�}>�x4���ZA~�٦KC�R,�}ra�l�<�������{��v�����{97�*��0<"�ޘ��m-��y)�ݸq��T����"�,)0�'h\$���ں�d�l80�K|�H����C
.�1~��
L!���s&�\��{x����Q��s���w%y����#��P=�۰YĞm&���`�A`u����(RA��z�I�b�iHk��ɤ��+��d�R
_hR[��hd���=��SY��
JH{�>�;����99�ҭQ��=�@�N��i�O�t�l�o���a����Q�ꬂβS�ɏ\9���ޠ��VR������T)�,<��YoQB��
E&}n�c7WN�����s��ǡ�aI�>g�k)�ai�����iHcz�	���Kd�Wn�C�)�'��	hS<������aL�h�.u�i
g�>��T��r�RKe���Z�q�g��z�9�1��8���o�ÿQ
ao����Ĵ�fXu-�H��@�O�H`3�<�R*L���,�u��a��/)<�3�T�����aI�r{�t�S&g}s�d�l<�w�H������o+~�_$�� `Ll{�"{|�0���9QL$�M�u&�^�����h�O%��Ԗϒm��>��"�X�ױ��) �}˓I��Bғ��Xq4�Y�f��＜��O�w٭�k��W_zaǽ0"<�z���)��P���,j��1����2�Ƀu��J@S�)���)�B�L�o���a��)�&~��4�Y�J~�nOf� �^����1�:�sW�{��;�s�Ϥ�N+)��z�;�Ê�Oz��0�ZAu[�,�g�)4{vL0�
KC�������(��)���)-�y��[)>INk0�HS<�\�k�7�g��}��s����sN/�)��)�>�#�'P�u�;��*�<��>�)&Y�����1�!Hs޽3ɦg�n�aL����)Ϊ�%2�Ô)�0�uA���a:��5��gX��	��i�B+��&�k˒zy��u
�Ef�2�e����x�`�:�����H��쌼�j��N�K�&�zO�N_����
C#*VFe��SX;�Z�ƺ)�ۆ����P�7q��s�✧Ih�cX�Z�j��<=�g
擴U~�� �����g6�0��o��ͤ���_hY:��}�J|�H���<ɔɣٸu4�Rf���I�W(���a�]	Է��g[h}��6�­��;��*�~J��D��*-�^!LB�����B�Fqd�e �����	�̔�&ꢇ�S�C������d�(��y�P>Ja�f����% h=�`S��6�{��R_��yQph�]e$�|=P���\V���I�aM���(�Af�Z[L����]@��VR�Y+tB�u���,���5�^�yg�R)�.�Xy�'Y�~��T:��2g3@��S�q
iO!���?(��G�xL �z{9�m%?'-�N��P�%6�{P�M�L�P�vB�m�9���'��wFnL *�3�H))�_��q�b�S�[��8�a�e. ٨�EwB=ys��Js��Q��T�x�-E �u1�o(q-H;�G�p�i:��kع��O��c�S
,)�.�d�i8�3S%������p�R�2d�,Y�J@Qk�<���y=w�����)U}�d�#�)�P�jO2�DϨ0�L=tO&^N���Y�m�T6��ACz��nX-�L�z�;@i-�{A���RN����U%�d�XS
C�)��ǹڲ�����뿽�g�iu0�[�Ì))L��\��O2S����d�h��)'��'��k^�a����9�>H,�>�,,�]=��RZ���)/�B���q\�:ُ����{9����>�<�g�8���T�S4���).��Ì)5��<�R���bE�aH7��!Ĕ�:�N{ a:��%z���B��_�7�Y
a�w޳,��tL!N��~5��֯�����3�d�UMСi%}Qm��W��VS>Ka�u-4f��S���n��L��2���ZC��%1fS�-5��I��B��Q�}p���:�c��V���j��W9�g�o�|Rq�-��Z��Km����0���3t(�̔��ݖ�'������jM2�A�&S]��L�a&N��i'�H�Ѿ\�r�|� �M߾�uY՞���|(%e��{�Wb���#�����d�6��9���
f϶6��/�Jn��VS�8�)~�d�7���\Ѝ��b��
i��IǬ�	�ȫZ9&N!�nY�o��0�#k�7�&�vDg,qa���"=p��BRܕ�D~����2�jx���?]H�TC;���i2�	iz�yRS�%"�׮JCI)�0�!����a�P�����5P>��d�cE<��i-
I�)4ɩ�^{D)�S�s�v+��k�U��B�z~K*~���l�l|l�t��d�=s	'�3�^P�J���qP�>a��=�1��9Q�G�-	4F���)��P'�*���i�C��y<���u�Ӯ�mر�y,K����W:��������F�E���%�U�ޗ꜁{������c�rx�l��B��b٠�q�f�E�^`X7�hTK֕��~Ш�p"S�7��:pmQ㔇:p-��ڙm�2{�n��޾퍱��f��\6
���ޠ�S�X��JF�|�?�$uリ��w�Un���]bh��P�����OU�ܰ-���5I���k�9N�;AG�^v�.7����<S(��k/����+1c'�<�ũ�*X(�נ�X~=�T�uBǗf^��@�f첟g%Q�&�J�E�T��X�o��E���f,�����$l�p�0�'r炑�M�<}ܲP��k��!;�ֶ�VQ�6���r�!-L��5��R��^�`����2 	��t�-�,��E�d�ϴn�ù�gq�J%��]�pN�h%eI�q�,��uM��uh��Ǖ�$���r[����w;A�l���}�c%�{
(��Tj�E9�#/z����=�kc섮�����굼����>�g����/=v-�ӯWa��yV�lه{�<o��G*	/zq����wٽ�#(z�q�Fm�U��#�Fʦ��K��M>|*)��0��ˡ�2�٠�j��g�N�c�;;>�U���E)D׼� (���©ŢJ��x�d��@9��z����*�.���)�W$S;��}.�D��`5
D�t�E]l,�Ԏ0n��Nr�Kz�"�$L3��3��s��r���h^C�u�&�v.����:����=4C籥	�ϋ�����t\�o>5�vE�Rr�
�E1-����{a�������5Zo���?��|㢨�V���L�9��`�s�F�nK�'N&(=�����eK�2!��i�J*�d��,��x<��H�,V#ਫ਼&6��Iavߐ�,1��,�;�O{����>{%9�Ⱦڸ��nb�ƽ�2�T{%���7lޡ�p{*�mشg#����)^���Yǘc�ڽ���f�P�7X��ʮ�
�^�����y߷�<�g�z�ǟ��4�f��Zpgb��Pt��s��L��{q�r]�-ij��\zi9{]}���bEX�Q�;�R��{�
*�XU��Z{0m9{��4L̾�~%��x�B�L}�j�	^�/No>�j�T|K�=͗��
r�I1F�"�F���Q�"6�eAP?x <;{;z\�|��̃U�朢��bӡn��@��N^�(:ؾjM8���AĢu��X:-ҵ`�Oi���k�s�jHM[���Z�B�&j)��[셙�p�7R�ً<�J��O��:7]AO/�r�s�S���T'��^W��-��s;;�9q��J97��-�b��V���+hp�MuSu���/(589V��E�v�f�=�JQ�d0��20$�^�$���V*�pT(���Awy=Ư��Z�y�Q9�;{TT��h��C+T�����Tg��ڜ�\R� R��S�����
�U���\�>�T��g���#�Ǻ͈'�/�!)ȧ#������f��ys�B�DzB�Ꙉ�I�֬J�Uz\����=E�b#6n<��\���(�Z��z�B��L�7z"mm��t&\�#c�k�՝��pW�$C���}N��a@Qg<9d��:��̪B2rC�5tU�gp�qn�e�&���@��t�����m�|U��>���ʎ;6�Crbn+{n���Zmr%۱�ͤv�l�+�}9g��t��6����ugV�θ7�;�%�X����<�u�x�rބ��s�5�m�M����]��:�\��[��B�b�g�4<�gZ��5I�H�>���I0rnL���#�ᓾ�̹�u�Q�y��q�{�V���j��K�v�N�جGc��Q��s���R�3p�$�pc�9�t��	��=��.���7�	����$��ٔ�c@���(^up�5�n�1����Ԃ��c}NmnP]i��W*����ؚ��tP�M�������s�a��:��lP��ui\][fYv-,��>�m�����7��`ԏ�CG�:���8��[Vԭ��'9uf.�3���mK���]��p0z����İ
�[؆vc����)���̘��p7
ÍI���:n�X2,C�����M.A��0�^�.ʻ5��ėR�]ֈ*:�'`+̩�z���x���6�m5��JW��i4{�<�#��8pL�(m�hu�ܧa].��b��m��":�ǯ>���7~y� x5 �2a��{�f��{D��1���{ps�媄u���[��H���3Ԏ�e�ާ'M����|z�5�w[�o���]�D�J|+�c܁*���^h�A̔ +z�m�BOӸ#�����t���	K���[���)Į�K������ےP5�2ʣN��Iӳ!tXD*}�>;��U��Y��G�]6&�"�n�V1,�Khw��$k���nA��"򶯕M�;c����7��[X�@wi��t-*�b�jK��p�[�n�+>W:�oM�m���>㵜�^(�QN�կ]f�U��e*�ݧjmn��,����v]�MB����b }y����S��Y�֖��S�E!�Еn�5z���

d)E[�Ԛ�'ڎ�|kp�;����АљY�J1cO�j�	�c,��ef2M�Y3��B���t5;���Z���&V%��-�R>��*sr���b�Ż__mj;�(���n�!uݻD�oe��Uh	��o3�JWj����B�0uR<��:�٠����鮌�hճ�U�R��+�ABV�۹-u%M
�6�w%H�A��qg�<����:���-����87�v��:����at��j�A�\w� [G�<ثwuwP]>1��q�Rh�+N�x���18�l��9\P��8G����V3�,|	̫��.�f�Sc7-ӫ�1��ko�98)��b�#�w[V�X�%Ov�ۮӖ3�t+޾�hYWf8)L�n�ڽ��j�{H��r�kyW�usĢ��S����;qG�ﻵ7SQ�h��@Ea�:���K�ҡ{cvP9[�'�(NTS����ǂ<�ٵEor�	Յ��-�*�V��	 �S:���HW��澫�|�3��劙��*S(Z�s6kZim:�#��Bh�f�s��Q��\[VZK���K6��9gwY��&`�cM�;�&�[9.�&V�pffm,�،:;K�Y�g,�p�N�0�����ml郱�����0�͍Ke�c�نE�;@`�1��f�����U\�hbukZ��3lcYQ�Ml�0�1�	�f̹9�MPq�vga���+u��UVl���Tf����6�$�����7R��lẶ��֫��h���3���ʆ��]Zi�VMƙ�@'I4���30s0&�i�ʳ�4�fWi��Ma��p»U�K��\�f��Zi���5mq��Z��`l�4ū���Wv��m3���3bk2+��գ6%��1����V�Vf�Q���ڐi0v�*ꮲ�3���J����U�*�T^�"��2�ooc)O�W@��:�bd�=/4�\�tH|s��|Q�K�Q�2��9��4Ǉ���{x�mb�Y��s�QW�r�����{J���x�0�]���.�|��_n��쫺{�BC��!6FP`5��6��꬇�	px]R�~>���c���XcO��)�pM=-uȴ�g��!aw��t�A�X���<)ϫ]B~�b�{�i��о�q9�;x�2�K9E�#j:0X�8IP���S�5j05�8�A�騼�s5��1�'��5����{.�(ŷ~�������L);�!��;��;X�O8�����>�xM;���K�;���ޙ�����6���4i�p3�!�o:l[T�����n;*�F�18�a��g�7b�v�5+z�MX6:�U}Bv����;4�{�c� ��(`gq����S�Չ%,o`�~wj5΀����AUN�WR���Q���p�pA�U�u`̍��;M��fM^ܿr�rԁD��27c�t�b����b�J
N	�m-h=�+6��|�@��Iˌ���Qz1��*���ʎ�}ba'O&ވ�r+��`[����F�M��5��,�L�L�o4Cɛ{Jcm.��\n��y{܄�(��%�ḆOrH^�����N��11Be�B��w�im�sБ��'%n�3��ܧW��F�m�I<���x���6��z�ɴ֎u�$�ELS+oC��ۛw���-�x���=���b6��`Ӌ�2aB�A����sy����h�,-�"�vU�35�Uu��B��qT�>�3.�;�ە�0ͮ4��R҉0̢�(��paߩ�l�of�3S4����f��Ks�MC��
K��+aX�}�>dqU1|�~��$Rõ����_LF�l.�y�4J��k�pOFI�w�
�?p�ǄO]��hx���\���VEb��x9O
Uq<2�nQ��ѣ�>�b����Ug�4������#V b��4�\;Ư:�)d*��8�z3AW�F�a�n�T_�B�� ��¦��XǍ=�\ak>����v<Z��
/ߜfudd;�Gu��'f*�{�hz�;=�iNW:�ՓBq��QM�SPkEp�s"�������^�7m�=�^a͝��[��fBɽ�/o�M�6z��i��ʹ��k&x9�p���B��ۑ-�ɔ!��A�x8��f���
w�HY+ajC�z�F������ꢰv��^ �S�b~4E�ʍ[��0�%5m�q~;-]�m,��@%ί��Oi�d���F�Ro �{�W�	gwwSkcwk�8@a��/(
���ts�9!�w�Lt��
��2P��z��0�7����V� BT�B�R�9,6�]EB�0��E��[�	F[��'V�ө��& �Q؈�x{��w��;�|��ڞ*�G�;	ȷZptkj�R���UC��"������Jn��7��;��\�\��
�8��r󘱋x��4�)>T�Q��A
�b�Q��Q�� ��R������%HH`�q0uP��a���k��"�޳6�`8$#:f��O� ��]ڕ�!N*�=[��^]:��X����j�+-_��ĨK���������(DEџy���[�n������įOC�T�%T)ΊU��6T��=O��y���R:G6�N9�l���p�M��!C�ɺ9�x/�VIsV�������SC�L���ԩ:�A��;<�RTa�N�8x+�`�w{TxxQ�����w����F�-p��=�9#[͇b�2�.֖�j�Ԇ�y9�r:
�_eØS�%�W�H�H���Dԍ���*�/�Ƽ3�.i$@��y�ۄ�![�s1NO�������=�Z{�M]G��iن�M���<�yy#&PG=��)�tY�����ޘ'oe�LM���Zu퇞�W�LxD��^�dB�Jn�p��]-�Κ�+� k��';y�P�0�,]4����ŕ��%�;�D�S|9�{6tW��c�Q]�3-�u�� ��S=���df�ւ�rtX�u4��� *����ݫ�a�=�I�p��sf؅�ŷ�{�����e�e��S�SyK*�T=�3b�I���_��Y�Ġ6N&5�o`���������z�JU�^ٟ����+|Es��Oq��#<\<*�����ӃGP�IZr�,ȍO6WF�g�2���r�9v�!:�_Ut�[�C���Y9]3���>���L��K���ȝ��{�!
���`��w7,�(�5U�q�U�k�9;���$�1*j5���/�YX�F��(�UnQیs�-:�NtU��a[t��EW��<���U������Ɩ{�˩๾���Q�T�&���x�\����IUD�@۾���X5�����Ie�Ϫ?P����V:�;4�pͧI�5�`�+�Ƴ�J�7����P�u�jU��7�s�fm*�N�~�Tk�<5�*w:,��jsaSO�����%�$B?G%���]2�F1N�w�/bLJ��Z*�P`K��J&��q�
gH���KBu��$8)i|y�:ќl������4���ptZ��\��0�v}huI~��zh���5.b��b.��$��+k0�"w]��f\�����^���wks5�Wu�.Woj���(��y�Y��e���(^6ooO,]��e��vPE ���ɛ4�C�l���3c��師���B�Ș�=6�ݾ��#r�"���<=}�Ӽ�;ITEF�dمc������e��9�]�T�s�B�������vc�gyn{s�i��&��z�J2�9E):p�U�1N��ވ���P�:\���9�a�Qh��J
 q�%C�C��U��lp�y\ù❸̪B2��o4��)���T���E�e-�!q�Dn���m�|VVk��={:�}�dx��7�ӷy�h_�9�i)�/��\��c�O�<P�s��T�p��Z%ח���y:�Ȭ���6p!�\8g�eΆ�:� ���\��}[Z��[�m���ǯ���BS�'"��ߔ}�Ԅ>u��T�C��[꾚�B�}^Voh�{���k���<�Rt�|}�r�`nێ�qp�%`;;{�5FY�kC���L��fcر{����(����-�bt[�١]F1o��Q@\�$�mR
N��!������Ό	��n�Cf�5�{��p�o<l��I$pf��ə�b}��(8�R��6i�p0t�!��mV���z�8!sD-/��pޏ\�q��t㬻�M�c;Q�*�]����oɯ�7BT�Dw	����^���+���������Oj��GE>f�c\U�b�TS�2jŰgt�5ܦK�0{����{2�s�~�AaT�:�o�ﬥirWR�!�r��W�� z�ar�$�d�P힄�uI^�16ڨsꝤ"���~;V�sܫ��s�gN�Tw'{���"���0�x'T�����砯�����Q��j���n����Nڛ�[�]�4�"Rˊ��8��s���/Uf����N�)j8c�ܕ1�|k�v�,�89R)��p(�*��P�����x��c��U��s�S��~�pLZt�m�T9�v�1���ɨ4�%W� DP�N�Y�%ڌ��R�B\.o=����hн��8=��փ׉�\��`�أ��3�D����j��:]��QF�.���pa�W������o ���'%�-z��6�5K��*���t�����/�^���E=+E�310�Oz�ܺ��4��bT,�=.�L�5�|�tC�)�����I�����D�vV紬Iu����p�(�3R��<��	���"w���"�\X�����e*b6���f�A����̋cz�T_�^��^9u0���QQi�}s��Κ3��i�^߽�������v�P�)��������Z��9���Om�c����֟6̫�\�s��b��0��ǡ��+q��{���YO=Vbm��Rd	$vX8q�n����ǹ�1��q'Z���n�e�6�t[|H��p�y:���2�)V83��=��3���&x{��ϟ-��R��#��� �����{핒���	z���wQ~{�����5k��nw2��i)��,h�Uh��Ǫv�6W���ݶ$�0��d�=���ٯ�!��3� ;�G��/�n�������I�x�"�-�t��Bg*C�%+7ٷ1�3���z�!*��z46:f�L�N�����!r����Ԥls����lw,o�'��#q�6�ܤ��Ӱ������՘����"��_��qb��	�ｏ"b�e�(��UM�
��GM;p�1N^s1`Oyƙ�$*�N+11V:����y�xZE>��RU���P�f&���r��c���"��1@��lr�V��}>S0 �GawFN��FELع��R����W�+~�/n3V�1X-_��ĨK����'o�0ƶw�N���{��F�a�ѯ
�k~8��!*�NtR�Ev*yN9
ٳ��y�v5����W+���\��+闂xl(:���x}X6$<xt��T��>y:]4�Csw�9\�o,ͳ���w�����2��k����j�f�gn���}��yV��Ǜ��Q���:�&V���m��hY��;aJ6ݺ�m�����Y���gx��@�kg�v�J�=�\��sndݴs^�;C�#�˻$LM�փ�M�F_q�
���������xu}�	c{�U��=?c\*(�4t^yg�y(��W
4��� �{����\`�7!2zO/U��ʔ�g(7�0r��-�ad�3�v|��|��q���W��vYW�nS�5r6�J��q�@3f�T�nS��u1nS��p؇Z"l�R�C���f�Iy��ﷶ��Ҕ��zk�(,1�}^���9�m�P��&�ں����T����N��\�H��I��!H��t��nj2�1^��6��lN��a�Q�4ݪ�ܙjd�ͫ�Ee(�~//`^a/yD^Q�o�-�Dg���]��70e�D߬�}u�&�7����X�w�����Yڸ��bb�^��sP��kNWL�~��;�ybCgT����Ij��a�!A`�bk�L�����^񩆔6����x�Mz�Z)V�/|[�ы������in�-��^9z6��Zt-֜���gM�{�й��q=kL��T'4&��	��\ـ�ʵ5N~�5��ƹv��	�i��=O%J�r�~���;�����M���e=��Lv��Q{7�z6�Y�1! }Z<�9,�-�wn�����i��I��o�$����M��v�(����cM��z����\�O^Vd�+h�9Y��w
1CE3�i�:�^`ԪvE��b�!]N��ϼ����M���|:T�k�(����!����j��5��ল��+�C�xJ��D�4ߥ��{�w5��[�O��v��u5�'r�tg�
a�Rn]��s��N^�Yj�)��!��8y�v�F�1j\�ڔ�bk��aL���s^�J$�۪{�X*�j��֧
+�U[�!�8e��7�직E��Tf�{S+�S�</��:Ԩ�WQIÙx��$�������En�X�b�*p���x����t9Js�癵0�ؠB��Uͥ�Y��	��d��,�剾Q}{N=�̨��IT�b��]���ވ��4+E7�ٙo��GN6V$��eq���Č7ѺW��!d��u/��_�9����N���6	�>*3EſGP�T�"\M�6��`���݊��1Mgq�cg��֩66�-��x�q:+�N���t�K&,U�y|Um.���p+�<s�o���TMp�;��Y{i�.���ʜ߹f51�,�c%ÁOk�m�5Y�Y.p��f6T_�k\�T��ޘ�3]��ok��2�NҼ��Rqٽ���|q��b��6�y�q#�E\�;q�c�uh�)�|Ĥ%q���{n�̓��fH��PV�T�&n�Q�Y��9�NQ@4�)g3ݢ�sH� �=����v��}UU���Kp�Eё_��ѽn�dwZ�}7O�F=V+�U��]B��,{�x���60��d����s~�Y��W�w}�<�X�Ġ�%@6<v�1N�ը��<�=�1�5q)2Z�q�r�p�d�*�t��C���sU��W�6�&6e<G���;�����=�TH6�>�F;���8�\pi;��[J�/�Z>�5��^��X��
f��fμYX��ug[�-(�z�FU@��h)Y�]&$�6:�*���muC�G:�O������PVh������a����N^s1g�x,�F��T6'�Y����!	p���r�Xjiջ���8Ŀ*0���c�r\���65�<݌s�ӽ�{�Ƕ��@)�ͺ;ܼ	d�I��g��*AǨv5��;Qk�үC�s�)��5��<�y�{�ʽ�ozk�E�#}�2�'T+�]���TaG)M/K���;0S;�ֶ.Nwa��Sx�0�n���îCk��XJ�^���<��+�RV:��i��Я�)ǔè��oo2.�	� tft�u-�ޔ��S����@o��XNi��mm��1}��T��Z���umt��P˝��:��RL0Z��ŔM9Q�ӭऍZ۝��P����9er���S"�n��vQꗮe�����Հ�9֪O�vRٖ�Ӌ�k�T����h��"߆D�]���YX3O#FWr�5��;f*�i�Q�z3T7��{ζ�0��^�6���
��kR nzӜ�Y8ޑ)ۮ3�!�����D8����٧�Uʲ�	�k��#`uEH�ҳ���e�Ds^Aӱ�K7�G)�Õ��ܭ�3\�M힫�Z��d`{-�	����6�o$�)tX	I.�38���JQي�cb�������rqb�X;;�X��u�N9[]ȉ�vK}q�
eD��l��0�����p6&�ؤu)}H;�jU��zm^��j�I���� �z��B3��7�&�p��qӋ/~Y��v4�1WY��d��0R�PI��m��Mz����'�֪�)m08;����K�[�jC�����u;���)��_�sxC���3N�C{Z]���Kp�������TA�v�rזZס���ە)4`�L�Gd��������1[��<Y��F9:"*��l8
�vc�]v}���wO�gۦ�d�w]ĔV!���5&��!����v���U��
��I��ᤌZ`ڄ�Y�<Z��
E�k
�� �Ck*	�*�C�"]�w�������ٻ�#�e��fYۘ���ْ������di�_GX�ÇX�e�b���O��=��y�N$�Cf&q��H�9g�`�.�^o,]]x��N޾(+�ů���G\ m^j�(m':�qy��w����GPW����P&����=o�p
FRO2����:�q9P�ùQB��ΘoVj��(�\/,	�GVfȈ�ՍE{T8�5��6	���ż�瀴mrcW|:����)cX�O��C(53՝+v�	{SM���ms��ɴc�մb�C�3��o�t���	쮸yF[��OI�}p�O�a��Y�E�ź�W�)p/�.]���7׈�wpr_G�A�Q��U�ގ��e.<эN#ܫ1^�|*
i����]D�y� PN*��#���Cc����"8h�R���ͮ�O�o5�
�їg��ɐ/{�z	r��$��m�ҎT����'"����t/GLw6`��t����;O�Ϋ#��9���s0���� *���t��������AL	��R	���m�{�T�������1Z/Ž��n�Z����2�e�)WV�`m�VL�e��Ux�^^�÷�Ŋ,;w�	)�']������Ɲ�1u�l(ibnL-���V �N��R��1��=��T�95;@�u��T7��E!]xf�Q�F  �:vV��b���͔d�9�c���8����QD*��47MbX�Y1����֜�9���f8`��cfs8��4�gK�Tr�Wf���K��r�Ҙֆ�l�k+-������3\�3�T+�g9�`cfN�Ff�٘�F�Fΐ��4�vqJ�q����JUM`�fsg�RfZ3����ʘ�6:�մ��K�XզZ�GYV����c3��l��;V��5YƩɧZ�Fƫ�
�l�lƬ�T��6gfm4g3����f����ە�)v�v�*��3WL�V�1�Xv3��lcq'ab�SI��8w6���pfl�fZ���q�[�5�ui�����M�8Mi��i��fer��0�1��N�M�R&;37�v8�b���S@�.�8޷�������<�6�t�BL�+fR�U�`�{hS'�����O�D�y���]��H����6R��y��G�}U��ld�s��Wq���-͇���Q��@����'c�!��1��a�JÏ�0&k/�eU��W%�*����E8à'�����9D��a3�
8G���4<H�u�D;�(��,���L�͏gv`�SrίF����(xJg�4��>���zL�Nۙ��/��{����<��B�6b��iգ4��.�n�Trh_\�u�5�תX�kLJ(����U�YFcMO]*о,n�o��9ؖ}���uKN� !�u�;:2-�Cz��W,�i��=�V�62f��`���S�-`���b�a�lO^a͝��Ub�JDe��"�>)z����G8T\Vm�z	_er�uYI�TL��e��!�̡8*!hf�$WZx�i<�J�����<;с�c��26f��ؚS���ʚ��j#c�������{��_vwj��Nf��=�V�jw�x�'"�i�ѭ�1K}��Uv�q�Kc'�S�ڌ�k3lK�N��(Ϋx��r���Oz��S�UU�sc2����.�+�
�ܳݥ-k9ˇ���zEj�%�i��9B���j�C'���iĻ3���n�u��g,���5�5��ܔ��T�cg�nr��]w�e�����S����i8��V�*�*ha��=�Z:�m���yP�� ��E��%��H�BUHB�� �Qxh'/A��+e�E��f,���P���X�2W�XW�R3X2���@��su(C���`��OiypF��b�W����(H���F�����v��q#=�yiM���B���֗P�J�������s)��[d<Z
�����7�U4��3�Fݫ�a�镞�&�����8e
��Hx���O	��;�����]q'�q�q���UY�2���HTQ�h�����n�\|(Ҫ�\�9ʗ7XxT%(n�笢���ޭ�ɓ-��Po g*.B�vNS;��D��j�A�R'��W!o,�i�X�0��(���QQ~;�h
b��9�Ź��(�KB��u�%��eR�z1�7�7۽ò�����J��_�Aa�x����8���}��=G��4&�Y�r�i���w�3�'��'
�˃F�!P�W@�L�Ks�;��sjA�pؖ.��Y4E����v�HN!��\U�
r���K�򈼣��մ����a����P�ĸ�� �����U�v�uP�6�V���5�+��-�Y`�C�W6�C���@ǸO�� M�/�	�E���2��gky>�`�ʐj�|.��9��ε%�j����V4̭~���� '}�ժ��s��}ӯ�8;j4��$���	�E{�������i-��3B�!���	��p+��}�&(ϣ4R��v���X�h�9����J����/������b-��uȷ�0Ǭ7k7����W9|j�OX�ً�ҥ�Z�)_�t�)��z�E���oUyA�W�^�m�9��:o`p�tќ9S��	�4`��QY��J/�&�ة�͘L�P����k�g<q�u���̚�DlO�޸�\��wuy/Ʃ���=3%��E�B+y��W8fӤ�
: ���q�Q6���J(o���({�v�^����Q�"��!po�HEbV&��P#W���.���7M�J����Uk���P����z��)�N���1=��0���S���mG
ծ�%>W�TUD�I¤o�qʁ���;�J���	�>�k�{ �E.f;2^��#��E��e�[���ڿEgJ�
7�k���%7
�R����*a���N3�����i�yLGޟDv�F��N���}���8-���v���
.�����(ME�2x�!�����{lm[�b���Y�sS�Ηt��rd����	����c����0�	ӫ�S�Dإǲ&M�ӧ�T�ǹSC��\�Yͮ���j�l����np�s���׭[�G���0�Q����qB/�*�����UB�TLP��nvs�L<�6�'�M\��HM��ފ׷MX�-�U�ӛ�v�yK�-�,���'[n��gfj`L�i���F�/RU{Q�_���=�:ʋ�t�K�D���c�zhJ,��Q4�\�f�)�!���j&�7��-lO��x�P/��4���p�w��ۜ�U�����*�>�H��+��C˳:�j�ڜ����ѽj�d{�Ї�}`nّ�:�l}W�W���᥮r�`�}���-��ظ|':l
��}��a_�m�F8�8\����E��V��w�39Lu�em����n�;�ح4W!̡��>��t~ZR��:�o�>�=�H):U�8;�5^�1b�2�u��q�Nd?6�\�3Jw��؏fx�
*Է9�a`�V�gHbtm+�*��gqj��+rE��W�*p]P;=
VjV���mT9�zv�����j-���f��k�[}�,X���"��ŌX�<��k�uCb{<��؞���)��� u޽�w��9*�(gX�#}w�mmg�����ҠG��ɩSٛ�l�q�p,��"� am�(Dn��i�]��,�r�����b}�ݗ|䵡k��(/�V��x
o��f	��b�k��R^F������}uK���P�{��n�o�pJ����Q�m[�%ֹz�:�̂|݌r��E3^���ѓ��չ��]�Y��Ǒ�g�4�\>Ǿlo�_��������➏�pLs��n�(]Ua���o��i3|⣤W����2�%�b��>O�-'�ʽ�J>7ſ-q�"��͎Y��j`�P���\P�!F�/O"<x?���Ҿu&:��i�u�Bw�%q$^�R�B�;��'2�b��h�*��H�Ƃ�|�?{49����Ti��IkJ5Y�J��]/��aN�DK��\d��2T�V�>P'�0�E՛�Wn��Ue֫�z̠�2�=/�]�:�#�aPp�:��S��!:t0T�xJg�5��!���ا�}|g��]7�ܠ�nu�_z����9��3�EE����s{5�J�gBi#�hO<�ѿC�4�yJ�*,w���F*��w./�^!/Bv`�THy]]E��kJQ�|t��v�c&��^y�ɚ�	�V
nf6-���b�X�vؓ�טsFm��{H,��嶭I�;S�N��r�]�����r5k�w��v]���I���E�b�����b ^�F=�j���H՞�;{�:�r7gf��yT}ne�ʆ�(�TK��b�I4�����pACx"�nZH+�P�A,:�o[�pf+�l����u�XA��𵻩��G���� ���������	Y^U������\mH��:js(�*���Ř�e%ٺ �*��:p-�xw�<ٱ�cY��5������|���?L��z��YQ���V�z5�]Y�BS�4��[t�|�N�mY�[�D���J12.v(��9+��z�åV��Q�gh(Q���8}阧/1cy<q�tΩ�%Q�F8`����Q
�X��m%�q0ƌ�@�D���Vb`�QfBr�&Ԗ%�E��f,�5�m�V�o7J��F�.@Y �3�f:_�K�`1-+c���ՔQ����v����g�^ci��Xڎ��0X�gj��R��|0l���tn�����^��a^��f*��ަ�+w�$TQ�P��y�i�L��aA�󎌪�<����t���:2��NEMB4䔹ZJ� _��p3�a��ܨJ�R�}���	�.�%^L��c�{�yokH��֔R�C7�]��C6�fL�.F{��*.B�vN�<l�]�±��aJ����`O�_X�BJ	�)��,�)��ԡ�]�XH���w�b�5DY��r���fd�����*�����d�U�"��i3����Zw��ñm������M#��|��+�ޚ����he6����VS����n	x+6\�&����{Α��x�(����F�����y +�QQ�;�(�T�\�R���Ĵ/!��z��u5�Z�{��J�e�H�(�2��ϑ~5�(,W�~O�/��� �c�{+�-~�F7;�홟^�{�5	����X)U���S|�υ��"�gL��/��ɻ��-˸<%�̈́���=���{f{��T��..��f9g]��J"��`4���1��"�u�i��0g���א��t�gj��P��>���n�9q9��Y��cz��;e+Ib�.L]����hC����N��ޓGν����L4�V
�V<h��W�v{��h#�����-�������r��xr�r٧刴�9�{�q�弗����m2�Ib٭����M���P�E���(�Wn�5��b�ђ{���T�X�kXƣnG�K��Y��������x@�T)����a�{���ޝ����ɼ�&������Oq%x����+�qB���K�L���R��m/�|k�xkk�*�Ήm�Y��]�� 3R��N���}ke4 [����N��Z��Wu����;|���T:Fu�nTҩ�B�Tngċ6�����]ln�SX�^k�+pR���ֲ��쫩ǲ-]�ݒ���0�iS��*�"wp������y�Ec%,��x��.�}ε�,J��ڙ�ũr�jP��>���T�ar��w���,e`�]J&άnF���Q�L>w]�\���~�hϻ0�J�ӯ�X�����I�`l�1Br��
+��lk��BS���r�N���3jbz�ӅK�Wn�w�y��T��z��~.����]�<>��r�.V�;p��d�X�'�2{3�or�osj�skJ�1B�t&��*f:w�t<UC��Y1�ƸW�+�5��(�wv�-RSs�;q�*����[ɢ�h�+){ą�!�~��g2�!v�֥�"��.�j��T>��*,'Ht��H��9צ��dVn���k%��S�F�///H��>��Ԯ��9��h,�c%Á@=��8�gUd8�!�ʶ3�P��OO�)P������*�#�۫Foc�^�B}cv��k�t���Y�̭�LSJg}�ǖ�ByªϾ����Z5a�7c���`���z�:��L�2zk��7�(;�}
G5�E�ơ��Z(���ڒB'Vy�mq|oV�V=g5��)>0�k/S�n����[��س���h���Z���t��R����\m�+��2wf�&��zG�ՓgK��tQFfQ	��r���������<gx�����=s0����k�O��0��J��O�MVӌ[�TP-�1�ڤ��W��B1V�7�I<r�BQ�?;9�QW�Pj��)ޓ3B�����np]��wkp�ܧo���ľ��8��bڤ�d�q����)Y�Z:�M�Lßg��!�����d�z�9�TF�0UZ��r�r��/s1g���:�亡�<��Н���}��a�:[u����XޅR�F'�B��6�ܰ]k��Po^�q��;اI�&��TZEO��ʋ�u,8.�������^\`����w�J�`np)��{�r�0^����ZJ���d/l!�J�㢕�Ѻxϟ'ڨ�A����Y�N���ť�gx�I]�G>G�=�{"�Ҋ�(^�S1L*�]6+U��:]�z(b�q4WA�kx�����|�8��paا��t7s(�(_�R�����V9�C�g̎.��%oU�Ƶ�ET/kR�)�ʦ��r�q�S�]�\,����U\Uϔǃ]��m�^�
g�  �c�5@�И�#4.�ٜGT��nZu���u�q��Ѡf����ֶ�Co�8Z��ų�r�OM:���&�@�˂�q�Z���J@�/�;	�^l�v��N;�(P+[�4�\7��>������.U�4��w+�_}��[o�y3T�-��uoB���w��j_��o�:b:q�'�
��؂m�rNL}R�6ʃ�㎴X�Uѵ{��ˬ��V��iգ4��#��-�QQi�}s3;5������O��/�+������8��5�,X��X��g��/=�x��������6���6���T]�{��ɂw'�>T�ﲏ�J^�t��k(l8�U��vؓ�'n��8�ݥ%�Y�+�hR�Uƿ����x���V�NW�e����L��m�,ϝoD����e-SU_U3�!�8�<;ўl��1��3W쭉�)�_U��<.�a����I=�����k�eո;3BS����������NE�Zr��zs����Y�o��M�Q��b&T0�ҋ��'=N���
gU�p�f)���XŁ<q�g�\^f��$��V���Օ��q1V:�
v� �=:��&��v�<zπ�Lw���D��c:���ǉjX�9�0 셑#�h��3~�BL"��=�^�K�u��wIw=^�+���n����I���J��㜹�����b��s�+�#R�Q��թ��{iʁyg t�S\K����3�Qc%6ZЧR��QeL�ü��[���9��2���]����t�J@��y�v��n��S-*���L9���bV.m�z���Z��ut�+ =nbSg9��
��p�P�$�Q+|���	l�I��Yd�F����xe�Si�p6m&b�pV+�	���s9������o�N%Yx����if�fnK�mZ��͢�w-�[���kٮ&�.4��3rPbJ���x��'��1�x��� : ���K�%v��s��c5<�jv��h������.�]����"ol]���;������\,V���ãHaCcJ�]g-}�SR�O{�.���Z��L���QoAB�f#�A���_ݕΒ˘:�_��V� F���b�Nޢ&�r�	��)�t��7�c�,��Ւ��b����:��^_E4���*��*����n��3�f�U��WB�߇eDS�#�����aW�m�"�@V\Őu�����1�
���M�q\����Y
,���I̗"�g=f�:ۢ/c0�c��"����֌��9(�����l���h3@���W���
.f �� �Dv�W�8|��F�q#�v��ݼK��[�=ޫSo���NʼF�r�Ke�M�K��Qqj�̽/rME]e�mNޒ�޽Pۡ�(�{ׄY�<-�V\�g�f��^�@��&䮄V��g��CC�v�*�0��]-��ղ�`�]鲩d��E l�6;d;ۨݑ֡��mi��F���f��S�x� �������2f[ഭ��n��Gk���uN� VPp���C8�jQ�Ԩ�x�ާBeh�9�rdpx�X�9Z�;㵨��^Q��Hš��X����S��)��6��i���N��L���X�8E��t7��a>�����5׻�3:M�g���q`�9��P����K�g�6�y�V�陼��i�yw��f�l���c:��t�2�>?j'Z�I: N��)�:u���]�,W3k���Q�L�3���z�(�7�p�-7/��%�7��B)�]g+ a�[�����o>�1@�ڎ�vugP��Wt2���_��es5b4��n�y+����Rˬ�ox�G�ۣCn^����@e�i̝G�h�Uv�H��Lâ��`�X$⩸*]�}ʏDJ��\Ƞ��,u�[��);�֘������EJ6���P� ��uJ��ˌ�=@a���W}m#�F%�05�ЌY[L��	���VF���۸WR��OsI�o5�v�1B��j�@�6���z���ef>��L%�9��O�fx*�E4�U�hZ4��/9.�Tq ����#r�!|i��[Ҟ�������KN�GF_c��WX#�kg%�Ej�/n��5xg/1SW�{���������9���:������b�]��f�
]�@�8��M��c��;Y�����F��bֶ01�a�Ա�4�خ�g�٭F���t�kCFժҺ�n�
�86nl
f:�Lf9��G7:X��w���ͷ�=nV����Z�枢��F�4�8�a���Z���b�Vٍ����n�g31�ltר9�����7���D�N��µ�5��1��9�g���n�8نg`6f�9��W��i�g6%�������+iٝ�co]�fm�n���`�<����39��g��fs`v6��n1���{1ޮ:��X�έw��u������ٙIUD�"�1{�co��Y�9�b�f���6Tu����-׼�>��)�!Sk��R��/����J#�H���Y�'f;Y��������UA9;�����J�~����;U�ӌ��A���Iu��?�|7S����������Rܖ�R*)�0�y�t�"X�Pu��:=C�
��<:wm���/�]v�4V�����4�>U�Z��@��[�
]vO�7w�'�+�
Q4ə��yl����q��U%������+�|���4�>����g-񮿟�t3��<G��OD��Z�u��[��Ս���F��)DԌ� ������ƅ1
�g:��8�3�/Zu������1�5�&۱u6�D��j�6�,�VF�n}��x�4q��洼�Cj#`N�V�j�]���%�7u���'
������J��
_���Q�'��)w���['��|}���񫆄�,�aˉ��ܾ�mW�g��E���Y���0VV���,��μ�F�mrK��^�@���f`�0�6v���;].�����Y�D�3�q�,�mN˝���H3��-����{>��ЇI�!��oa�[v�zy�ΑJ{��������)��i��<.
x#M\�1�:����T{4�n�`�IB��3h�*0���q����=�vW��6���m�����V"�]{���(��]�|/��aCx��ͭ�43`�#f
�o��7I���k-Z"�qۍA،4Wٽ�K����3��Z~YEx������k�qO:��{���8�,��Y��7}��,��Z�4n��Κ3��PU�`��6H�o͘=��(�Wn��^i��ٗ}AB�M'�v4�T��-�|(^�ǉ�(Wq�~�Vh��u��
����w�f�\KP*�ɬ�Ԩ�2�"h4���9��>�qBuKe��1���D�>�B�ԡAP�r(�8��۔��|�D�$Ɂ~�V���V��g�ڙ�ũ.��KؓK�aNtd����X�%6�0$R��N&�^'#}ӎT�Y��S���������ī�߸r�G"$s����)�l@��b��R�E��6aF���!)��n�)��`-�е��z&�'��5�.�,�P�Q^�S��9�˨�{*=�̨C�Qr��V-�5�y)�޵��J�'/ɂ�DM��"�t&���RF�M��UP�!VL~�>��={ ���N�Up&;,�y'S��HFC��T��M�xU�����J�E�]�D�[L�[s��=p}�ԙGU�*�*�GW��R�e�=r�<������e[�k�ũ�������� mǀE�r�ޙӺ�m�����-�%.�ri#B:7�S����q���V
���h�*��6�_dv��2h�1< RR�G�{;{��3�dO
��f�q��8Ku�	�,@�����D��"�@�';�l^k����8x��xg��s�5�
�\)0=�%�C����Fܵ7�\!����ST./�׍W-e{���1b����u�׺�tf�<��u�����u���R:�=�j�2QW�5o�dϔl`%)��]�;����8�8\�����b�����eG�=9�yĆ��B-�]x|4L(:��;\j���╯	�T��/\�$�mR
OBb�^�8M��[��:�@i����gF&VMVtє:L�X�ex�
=�-�٠�r(i�n��gZj���Z��"Λ�h	���q����R��;=��c���w��R�s��u�72I��];v����=��.RŌY��8X��k��lO`Vbc	�*vU��A�k��y
���,@M�17ԡEE�8���u�^�͍�r7c�F""��w�;�{�;����CTp�*XRr��ت
=�]�p��Ӄ����׿%{��0KI����t�鿏�sb���1��
��2N���C[�]�>A�t�0�h�?^�kVm���h��42�%�Ī�5��vr�t��˓�!K�5��9P���G;x�3d��t7�^������Vo`�Vk���i�`Q7�:,� ս['o/����G��݂b�U�M�./I��%T+�K�Q�ʃSE�M
t�RP��Y6�;P�����u�
��<|s��G�H���_:����	쳗H�Qa��w����q�.����×��[��5F���HVº��nW5pm+����[y��Qe��}^�&۞S0+��QN0�O=v'å|���(+?p�6b����
ye���\GI�*��v�����U��6=��;3�M�:�LPN������HWR{�RUE�Ӳ����P�cE����H�Y�MAn���R���]o9�R���,7j*4Vɪ'��Z�S�8p�QX��n��N_"��8�u���X��%���`�z�-�Y�:|��">��0��⎹*��W��m�Є�Rpy�6�9C㒗�_�اҕX�×PV׌�K�w\��[��D�y�'r� �����˞�xPsT'+Ʋ�)1K�g�K0:Yg�a����#M/�ש��bg*C�������͎��%:���>���[٣`8��p�٬�BRr����ή�˵�}��,b`�іv�g+��Z'E��$1�#�� ͭ4��{���DHNh�Q+y�yN�+�֙�� vM�0��E����ɻt��3/_S�������Κ3���d�)��w�:Ft�����Tё1�X�]Z����!)���+@N�m�NC��	�f)T�\�5 L��X_.9���\X�t��u[��J���GM;p��S������wos�V�a7sf�\��ݭ�����Kes�Bu��DKbN]+���uب�!9}nM-죂P<���m�kN��(��ޖQa�M��� 셑#�h��J��Hb-M�(��^��K�-�,�h��G �J)�W�� LR�L�#]�����T�Xo�����t��~=�p-��¥��bK���'��I§G*�"�-�0�F<��Vz\��Z�,Ny	Q��p���ұ� A$��Fe���Wo,�S�a�jr�2��:P2��X)�l�<��МR�H1.bgt�֍��R�,e@��t�hiU-p����ᩊ�徐�݅����pB��9���1���\�D�7�j��Fڋt6	Ⱦ����![��:��/kk��21O������Wx6���3�$�R��D�Wą�]t�x���8Ϫ�U��o&ܡ\���]�v��=d@\`Ĭ�D���m�4r̙�Q;�~���~��{�fv�(L�WL������f��&�|!ۚ�6dj\p�g,�'7�+���=X��.�Q=y;"��Hø,��#ه56�1�Tׁ\��;DU�ځ�r�ol��o��yPh�	�����!����Sd:�����n��O��W���ݷ�����`.��8�)�W	��Y��yӉ�r�������>�,��G�Oa�ۼV�>�y���� :�S��f��&;�agk�rv�qȳ�p�+�ƽOm^Q�]L�&���8j;,b�j�=��_p�>%��M�'\�n�ǹ�Y�:��D�̫kc#e>�x��S��f� �4��m<���]�ە�tϔq�x��6����A鵽���j;$�@J��]�aR��(�VQz]#HwF_��-�k7eԯ<�k�G$}V4�#�w��<Q�]�p�t֩�TL�3�@��
nN]"�:�*̂'."���&�Im�ܾU���)��_��񱋰�uKe���k��p���k�xo�cN�Y�ޗ+��RJ���U��8e��5jM΁ʵ��X�;S#\��'Ν�Kؓ�rr�_e��8V�kx���lS@lfT�����8�@�u�.�<
,��5�uU{Նee�����&x�tT�^�w�V�R�gǅ����t�ib˃t+@�'^,�ދf�N�����+�D��¶��&n�L]���W�,E�m+W�˗a��Go�i�sVLG���Eq�7��a����Y]�> ڵ;ݕ;���b�)RH�bq���:Th�*��uK�c�م��s�$%9n�)�f"ң�wV��%�U�fԮT(�#���.��Ѡ(�\>x}����ǰ?VbtM<]zR���M1�]���m���*�ʊ�X(���*���ed�T�8��ęx�7=�X�({3ЏC����.��*��h��<&�Ss1Jzأ���4�����1S|�Slc��J1��T>��eBr��&.�^� �Qt�����e������T����ʝ;�cv�5x�8����`K����s�VuV�7�'�8J��p^eђ�G@`h��Ll�]mj���c�u`���y���Bu��o���e�%w����9$ȷ����)�u	���WG�.���v<���`�N!������˛��'���mhElv�Mڌkq���Q�*g<t,|x�>���L��t$��f�D��ٵ�i)#���q���w��΄ʾ��W�iN����>�$(�Rܾ�!�t�L�B��X�)�zb��8^�$|�i�bT}o�f�xX�rŧ�*�/:��#+���N@p��Sۥյ�[8+�t�ZM"�3�p��E:.z(IS8٣�\w�;���P㨉�)�56�IuzT�ƭ��-�4�A,�,/)H��y�R%aJ�ư�Z��1�P�i��`:Tຠvz4�f�oQ��hs�����=��s
IX1��%R~�
�v�\�*�.��`�,b��8X��k��lO�ٕVKj�M��RIq��4VB����16:�(��8��rԁG+\���r���[��I8�]�i�Y,�^�^�5$�Ԡ���=�
=C���ϖ�Q{�c��U�xX���l��=2M�Z���:��*b���o}�P^�!�KEؾ�v�#Q��d�u=B�Ž��Vn���q��ݺ0Jg�=4/dXiE�%E/J�չ~�yu�S>�u��"��$ۂ��*ÎQ&���+)��b�����8MFz5��A
�\��B��QtuP`͙~��5��}EΩ�҇(�S�Q�`�%։����gcT ������=��oo�W��W+Ƈ�b�i͏`�Ì�SrΧ��1e��P�hW�\�I#"Xޱu|/���6�=�Sq�5ۊ��:�f�x�`��,�(:��q]�ۺ�쩳��}�"�w�r��ӕmi�(���~���n��*-�an7�<k�ė)���0�ۖ�f�/{>�݈X=�[�4���$[SU㬎\cꔵ���S痃��a�8�x��Ǵz�}bmȭ1ù��f�.�����`��0���V1�M�m*����_Xo�
�xg����R��+���$i�E�4D�n�m��{}{����V0��~R��H�����̮���Lw��s���{�0��x�l��BN�A�[7���ME�5�5����W���p1q�B'�ĕI2:��]�Bg*C�����xw�<ٱ�cC4:f�+bMK��<��P���q�y�N��^�Ԫԉ���eո;�B����N�Ma9�ZptnU�ڷN�,�������6m5��O���m���b~��B���S��!Z6�7��<Z3�<×ӦaI�\��a^��:.�+11~:�T^	�r�%T5�OZ�kq%y���3���6�lA�H�u�Bh�E�Buf��.�f��oNs�RYw�������&)B�jf복Y���T�ѧ��n�Kz���'�@�+53��g7;ʵȨ�f�;�y�a;镀K��Qaj��2��~�+hQ�sUy��uڹ�3�2c ���[�8�۾9��I6�0@t��g9㤂�t�cu�ɡ�[�w�.��gPN�V��t�H�jB\]�kv�v,Q]L76!��%�%�Q�1�Q�-���� ٮ�z��74�-n�b7�G��s�TԐga�Vf��U�*�-M�P.���
w�>���ЕWV��L^�Ru�ѯwogX�^�Ph
�_P�<|��%�L�.FPo g*.B�-�Y=�$\ves�����Q�����
�!�OV��_�P
�Ȓ6�ht6	�֢�����]������pK��D-�N�Yk���8�%!y}�D�B�t!>�+T�S���Y���}ê��z�jJ�{�.���B"�������9��ы�������X(�ee��C���5��#7���̃�W��Y������\x)�s�	{�yG��5���;���1��K�+=[���w@������`���l�r,�\g�m���TT����%z���O�ՆϾ[o%�OZ���o=��Ї|M�'\�x<�����#�`��}NA�㕾��
�<~UtWT�z#�v�qOU�yA�V判l�魄��l�.<�e	*
�U:o`77�]>��p�2�H�o.l�X4��=&�ڞl2�2v���n�g�h'B�w��T�]pD�KEi�V���l�wC��v�����Q�㋃�k�/��߅�n�][W7i��+QǄdG��ԫ��L�����.:�=�V:p�9.*�3*�/.Wv��J�.����(�^�N��ۭDvmNoc㴪!M�@�백8��ח�u
#_<E��1Q���l��S�J���09u��j��E��%�UH���Sq^��c��vk�ƣ���L�U�e�hT���7t��A�jq��9M�8r�ԣw�uɕ�*Gj\��`1�<�w8Yj��hܜh<���̂����{˜Q*Q٦'UƵb�)u ��s�ݣܺ j��'����޹yK(����x��唘�u�5���v�j^_M�̖��Z{aϑt}���S�Ԑ�][����yf<X7!� +H�[�l�^^QO�=q��d�#���p�9\aܷ'uLU���^6�]B�'	%��������w[A��se_9<����3^�am�"6�ҏ�ldsx:�2(�{+`�����Z;V,����A��ѻ|�9��yPDC�6^��{,�ݍY���{b��9��e�=f��6z�%�d-5��=yX�5�nF�h႞�ث�l�6�u�y��:������w.�k-+�)�nS,V�t�����Mn�X��b}�d��UeJ(�q�2 �{�p�9�8�惷�ۉ%�^��n��2�j��{JN;%�s:���:�e��&'��*\!�DX��S��p�u�f�����ý���*˧R�@QrZs���V�y�d��:�6	�tG�KL<�w �]�-0w{h{4S���zz{�I�t�X^u��-t��u�m��`�)0�3yfu�n֋�m�l	�E�.����sP�G�Mb�����:�V�-M���f�$�+]젃�|�����
��U���Z��u؍����J�X�Ƶ��.^���F�.;F4m�v1u��yO\��sW&q@�n�o�!���j05�hs����U�;�=�x�P,���d-\�T(	�2����%�m�
*�-��z�'9̈A����!��B(�)G �ϡˢ��k��{:�n�άՂ�KL}����\Sbѹ�kYGe��h8�9�'Z%wpu���f��H̋^���v]�=��m,��N:X�י1�n<"���k��M��R�]�5Юk��Z�6�uaiu��2�1	�wX���A!± m�2�9xٶ-J�(gE�K�h�y�7WQ�꽩�6�D'�v�-4�jgsi�#�R��GM�DT�o�q's�{��xQ�1�P]�T.)�1F��
N�:n�{�Yc����c�I��ַM	[�Q0���븚���Էv��}kx���VgG!x#�(�Yfc����gc��/&�GDR�'p�z�'L-[�� K\��e���}r���_P=``�D��W����c7o���W��a#��SL)F�A�n��'�ⱶ;y�wlv�.�;����9Z������f���fv�lq�Ӄ�&�V7w���QwDQV[l�l�KI�\lq��m�9���i7���mr�6<�㱦�̓0��c����i��8�^��޷=mgq��fs1�6�0�T0b=�{Fn���lp���ެ���M�'M;9�F�ձ�A�c��\v�lj[k�oz<���ͫ[��ukzќV�n�{�lj�9����:t�lfy�Λ��`��Xfc��Zmz��n&��u����F�7��6�w�L����1���;8�2����lmz�fw8w�Ck;D�6d�l�lo������Z-�wM��%�t��O<�U���9U����f�.E�c�o���%ڼOH)��o/�G�V���:x��]����<q�w����_�Kt�\0���R���WP����¶��&��׼��m|=T�Z�����}�5�g1^W�g'T�Z$h��Q8
���ڵ�����ռ��#�1t�at'D��թ7;�U�F)B�Jd5ьS�Ӿ�n���	=6�B4�Eq/���7T�~�Jh
T�o��r:-ʀ�n��ބ�(�]tʊ.���۶��ww6�9f�9�K��+	��)�t8QHt�0�J׍����j�(�f��=U���I+���*�*���{<�V� >5���Dg�F��N�G��,ʋ���NRj�ca�gW�8ʵ]w�B��L�7z"l-�"�W����#�n���:�n���ڞ"�L4U�:!@Qg �$�N�Bz���7y4v�u�����d�Y��o,�'ks�����Sk�M��v�9��q�w��T>nn����:^Ċ��|��mb���t�-U��D�|+�Eի�;s�7�^��x�8�7:Y��.
{\#n\c���<��r�hWL�DwUO\�s,-�)��4��Jp��e�& ή J��g��<��w�@[�5����Y�۷\l��?q=N�j2N���s@�x���S�{X�_rTn\�0�nݚ��tr:�T;�s��D�ɦ���W*+��6J�,i7��d����n��[O,�vu�7[~�X:3{z�wZ˭���d�l�0ͅ�æ�U���������������j��ݏ;����78�qދ��Vq7��I^h	��ba�{�	^��r���2UmyU���Vӌ[w��vF�at4U�x㞜h��hI�j�rt��p1�<�	�}�B�xmfm_��u�.[XZ��#m�S���J*�tٖ-PV5U���mV�����ڷ�����ԭF'�޽�����\��T�$�w�Tl���",C��ҹ�U�\2)���Xĝ�	;��Y5�e��}	'��-��3կ��t�`5�xv5T��3�G���u�^�P\�Y�������ǉJ%L�~j��*w�ODW�MG	1b�v4ǟԕp�}�}�~u�p}�@���;9�}J�2��	$2yOYV�����������ob�
^��X��]���FDɨvnl�{~��n6Wj�.��\�K���;0p&{C2+$piE�%E/O)��r�q�sӧh���,���]��3��ݜ���t�WιЭ��x-��l�z7Vҫ�ZRY4���/R�q�|krag+���x\3Ժq�Jܘ�o8y�ۊ��8r�3�,����̺�yR�){��\��BM���q��LPr��-��k���c�(*%dN8e-�Ck��uK
^���(�^��{�[��5�
J�k*+&�,���ZӕL��+��HY�(7S����n������k�z���`��u�d���S������j�v����b����U��{uk�]�����0�8�3R�;�woz(��}ƭ��Y�����^J�Ղ-����Q0��]dm���TX�:�f�x���V�q=�<�]Ƿ��#�,4��E��/�s��t� k�4:�Ȼ�"�����W���N7�ȷ�(��oݧ��Î�����;0��u�;:3|�3W��L��>���v�J��'NU�'o`�(�ZT>�~�a�hI�k�9��yBvXf�ټ�zj,���:b�_g\<��z�)_� ?Lِc*v�O1�(C�9Pb:p-��l���!�3A��svo�_8��K��1��h]u[�1��.����!)C���N�M�*E�ؕ�ޤm����U��s�sF��to%�o��66��ŉ��³mW�?Oa!x�=����i��*��V���#2�L���EP���#}�w��xR�pe����Mw`���ҧXgE�O���d�GJ[ypv�'�=�U_A_t��Nv�-����@U�K��s�uD�4���h�٢�Ϻ�7ʐn佚�NڧV�x�"9{[A9f<��S
L
��Ŏ�`�-�8.���/oΐ>�1�Y="�F.���f�:Z̑}%�����."-N�	�o6��k�U��X��<-��6`�Ca���J�P��ۍY@�j���b�,��`޻;U�7N2�� �z�)�Ï4�,IZ�b:�b�z(v,*tr�r*0f�;�~%;镞�&�֫�[�W1Xڍ��K����Hq�����w�I��
�Vr�}�'�
�-ᅔ�}i��7\�%ɸ���R��>�>iu/���|>�m*��C��Po r���C%L�R�h��%M��;���*�Dߓ�HSD�j,U��X��EF���t������a<U���'�r��2��Ы��~�:h���5YJ���k�䠰�gԩLӺ�o��נ�ϽE>����,I�j�-:��j�u8��!лA`�9D��)iu�c�~�Yze� �3:�25N);��;�͆������_Y9�Qχ̾�7�j�s��O. X��IM��ᾝ�2��ו-�F�ZT1����lg���#<(�m��π��6i<>�k9�]5q	��,[)�$%3E����Am��LPU��i�ЅJ˟f��N��3��ݪ���t���}�N�G�2p�㎱]��^3C�C�V������=����-���Om1�0��~���u��n�o:!{�_��]���>X�r�p7�� �hC��&؇��E��m؈ܳw����Kf�y���oJ�{"�V�ѨS�<g�ס��XK�xp�~��C{P9�q6���Y�jy�n1Ȥ��Nt��k��t	��bțSu"���͘�<�."�MW�l�KU�P�]��|��ƹv��'Mj��&j���hP���5yݙ��֧xVrNRU�D2���ӹ�4�'O���
3��+�qB�;���H�k�'̆����_����S��tt�P��M�qʁxjԛ�S�G1$o�ω�~Z'��]	���^��;9#�{S�%���w��T���m�}8�@�u�.�<
*l����F0��%�*ga�ojuH��`R�S�Ĉp�U�p��t�0�AZ�x����]+ձ��㮛JR�g!�t���=%�;<�S���2��ȁJ̿����E<��'�XҺ��"�l5�d7�ص��.�;�4��y�O1l܅v��i�v�'�%6����
�%���0;� �	d�-���f}���-� ��Y��,w�p"���<�'Kb�n��r�Iܦa�x����Z5e�^fVu�ds�
$7!q�\�oD����z�B��g<p7z"o�o�P}^TWR�H�����2h�{Ӄ�����-��:"��d�LnnH�E���;}��'�u=>U@-��{G��7�53�cA�k�m���K!�.�
����y�{n�+5�_���=��j;��,@���ƵB�{t���+�ܽ��ӷ�:|}�����J��g�S7�ݯ���P/��侠����㴝�u�N�y���A��]���YG�-"���Y[��lv�<��ք1pfC�v����rU�^��(U�zn��oaOU3k�]x�V[v<�߆H���]F#��e��8��N�gk"��j�g�ǜd����s4C��'Գz��[F������4��rk�a�<D�ͪaIү!�����+����}����+f�՟	�`�}�iO�,���T�9}Ai�P8�b�MQ�n��N�을R�R�M��aؗb���VgD�`�T)�N�p�°v�\�r� dS��P�S��;�����ˊU�Դ�1�F�qdV�a�~��E򦰝�����Oƒ�M�����Tǚ~�7 �u�s[8�%"5+�gݙfjYx��A5-���׺s��m���XNVI4�Y�]L<�µ����J���B�ư���μ���L�B3I6Xx,���rcjEϯ�z��̜�GU�^)��������T}m�s�_a�	]8�yT39��KSԔXJ�2T-K��S��Q�L]J�.iW�M�c���H��{���s�L��34���w�Oׯ�ʎ��������������b۱|�̦�9�����i*���f���A��p`����	���н�~[J(E������3�^d[
�)[�I=���wk��+T�*��XQ��Q��|]R��"�����8MF� �E���{�2��Q�z�w�}L�3�a����E=!K�Xs��߭�g�}D��J�'N[1��J��**��*�âRx�m�8�$O��X�
UM�>h��{�n.n��������x`�
�K]m>:c�F�g�P[���B^Ε/m%1�]'Ó��Yj����,'j*,&�����¥V��U�x�u���,{қ�ǎU��ɝ|\H`�OExE��1��u�Ӯ�n�,=�Όj����3YG�/x�]�n��lP�f�{ȴ�Ť��]����W�`mk^wF�2�t�^��� B�ܺ7��˾�8\s|Z9Ֆ1�(sROwIq��n�������xb�K�1��9S��Pӵ��2��!0A��JA��F�vp�G9n�٠]v�2��M��@W���C���u�V���r�\2�����bO^a͝��Zv_�4��|�
j������M�o:��B��2eN܉.�d��r��<t�[vsc�f�A�u)>9kM��6R)$.f��h+ixc��5��Ԥls�?�GP�-��C=�w��x�ع�.0��̆d)[ca��f)o_�}Uv�q���	�S��;AB�귎f5��B�sP�;�,����VdZ�`&,a��8���:�D�0(畘��^��:.��������싽���sN�%-�q�\�nT8��,f,m�������#�h�b�J�n�r�-9�U;���,�r$Gq�/ݩ��j�+-_��	�P�KS0o���Vy�q�# t"/6S�]Ƒ��*�[�U�9�
3.}�ÅN�r*2ٳ�߉�w�*��|��¹E��qer6lK"z* �4T)P�]_M�n�`U�9Vj{(Y�xaj}uj��^����h��|����3ǅUԸ�
����ΚUK\ ����
��F�M��uM7�4;��M���e{�N�8� W3��-��wFϳl�27����V�h�^��)q�F��V��z�>��!�J�s��p zs��4�n
�ID[nb��ΐ�܂V	mY��FF���)��p�G+9-S��;��%"7�L�{���9���a��$����u<��#��@�Z"m;�UD�j.����HE���w��)B��SYM�%�#seB��F�:��8��p���DIt*�P�D�S1NB�3s����Ĥ�\\S�V�ml��T")��6�����=(y8V�Vו9�=N��m#���<�2��}����a�߀�lY��FwU�bwśc�ܾ�x���A�V��j.��kj
5,��V���a��|X�Q��ヾ���y������a�V �^n��:�"�^50yK�m)���1J}4R�ه.'gmQ�8��뗯�xv��y��{��v�͈8W�mP� �y�=e�����N+j?]���>ְ>�W��a���Tm�ƭyy9+^S�����c��N���Nt�t��
�@��,��6H�o�"::�����V��8Ik8����J�(�Wnޚ�Y�k�x��*�3�7[ͺ1fmҺ.1�A��Vunam+�Y�R��5�~;V�sMbt�Md��c�0S�]/D��U��r(�tE���fy���Z�y6jQ��,٨����L�m�u�m����?�6א�Șc�W�}�Kƍ�v���o� Vߴ�Z5��"4nc����e7�IQ�n�.^��i�D8s��Z��C|}�۴�c���V��T�	/3D}�KP*uX_˯��k���I
訟�W� $1�鈬J�����&�G*�#<X�9ڙ��J]�L�>I#g"�Y�}R�D��^�
�P
�E9�J�M���r:-ʀ��t�SY��
���Z���$�U�f�~�3��L�)pU�V��u�_b��po叝��ھ�6o�������H�g����C��99�mN.v()��/N��S�e�@LM:�1S�E�3ϵ+ETb�0�)q��Qr��<���S9�*��t���?������`��\�یݑ�>}��}������ҡ�FL[�8W�̏3��y�H�P����T�MIȗ@���Ĭx�[(�Ľ�n���	���.�X�������:8��*-:C���S��իy��D�RC��08צ��dVÉ�\����ϧo�q�nt͇��{�b͉����̫�P.�F��&���\
�	pF��Z�#e]���'��6�/��lgi:��,�"9���!�} ��5�'�<)�u
���,*�>�hՇѻ����Y^wuv��̯Y]�v�]�^G����������l��T!Q�V��%ՄۓUJ��z�7a�dÙ\�{����喩��I>'�s��iH��:"��N<I1���.�E���A=W�-:#��v���q[IV>E�\�t�r����'ꆰ+��$�,,�%��G�;c��P�Y��-Z���n���w�o�,�l>ˣ�^��^���h	�2��--�i��mk�5�@�5eN�o�n�I}F>��e�}��r�ϱ�:�[!v�
���k�6�Lq�F�M�pOE���
�:���y6s���V�Ә�M(m*l�x�v5c��*��v� ����+k��ꅜ����1�̚��K7�|t�\n�(�\8+z������;�H9�˱sܕ�_k&�v��L�=��U�K
�T��2f���2�zv:�A�ڊ���"p�����x��gg'�yAje�57�tq\�;X��^��۱Vv�GJ�%j/v���~|�����P��Y�;�L�-�(�opS�)�����z���Gn��4Aڈ<4K����Ƭ�/n��[����t�5�[��'nø+8�p��D�3M)f���W07��������o��qc����KQ�uGN�"Wa�1S;+>u-����n��M�ajWc>ۯ�=��|C�\��Ղ��7�M�wv,>�3�V��%�֩Z�KV+2�9J�uʵ�����ҋV�!�`��o]d�p����h��z��T�N����bL4kjB;R<kvż�����;\C7R�议��Z�6�W=nU�6w�]j���\q��o6b����k�7���spׯ^��g�FJ�����/U2�Y���J��!y�1y���;�|��1���Dn��s����}��!CzR��juک8��q����ʩ��ʇH5��[��8�tM�Z��m�'-e���^&S'j�t�
tx��:��x2[Z��m4EA��ҝ���]3$;�!v���4g̹�������&T�8�+�t\	;�:�V�w�,h�,ː�37��b�aڢ�[voZ<��GDzC���=��1ȋ&f�`-݊V�v��*�g"3.�ƶ�(���L;ڻ�� ��И�j��T�&*f�=}Jﯥ1�t#�^���Z�]����LU�Nzqc����h<Ѵ��@)CaE���s�Kn�mt�G+�C�+r���\�)b6����Kg�6Բc�Aťc&���ycڕr�&k*�s����7푂�_���1Н�����׸V2k9���`T^�C3OF�u5D�K�8�[��&��F�LLD������'��V38�$�+F�ՙxRJֿ�YN��q\�sEr�n�M!�3(�ĹU������x���S@���x�Y��,�׵�FY����RV5W\��SG�4��kT£��ק�WKQ� n�ɝ�����
� ��"�
��ʳ��ڠ�6f�clc�\벱���s��32���ޭ�ه��'M��iӴ�MӘs:�ɬ͙��x�����Ӈ�Ʃ�f���v�gz�޺��yc���f�349<��g�36;�	v���Vp;�X�M�m//V=u���oz�q�Y����N��ӌ�3�-��U�v�6;�hp�c\��Sc0�ձ��4�V�`�v�����bn�{�]s�5\y�m �1�[ގl;�3��9�قM��\�1�c,ʻ���@�Xzh�\le�<j;�FP�Ej�
ɲY�����TD�)]��}X���'�=�K�a6�-�Of�{-���<IrEy�o�aЗ$گ{�oc���kq���Qc$\��m�}Jf�J������GSV����/�~��,I��� ��*�|��ҽ�L�7��0�y�o��k��d�4G�:���#��5%M�����7�tض�|����ո�T�Av�y]u&�8�o{�NDg�p*�k�i?/����9��S�mˀ��NW1B��}y��f��EF�r[�k���e�̡xUNw��V��Ү��Ѫ��堺���	�����5����SEcZ�+�T�t�Նd�v1�N�)�W�@5$Ŋ����wT޻��vu�/vq���u}q��n/����W�����=:͉�N�M�N�0"��gMT�Pf����A�Vp�rmFFyU8q����K����f
gp5�B�B�QB8!*:j-�L��Z}���K����JlV���vg(�N��(ʗ���A��P���4�
��G���6V.�4EĿh��3}�UL_<��Ȋzeg�6���]�� dd�U����7/�'�{��J*d��4}�1�ѽ�.%�r����׽�	u�K���^K�ҵ��D����Ob��7����+�*�͚�v-utY�4�����:�e�:�6C7��\�����V6���+���:,xں%�����X�	�z�u�M�T�k�ǌ;=�e��`����)�پg;�{���5���pb�_uO.C�Y묍�v�p�l�<z�1�[z���'7������a�ڊ�	�}s��)�i���cƛ�U�|,X��k�8z�8��Oѩ#��@�����c�%��{���ۺ��ױ��3V�\��T�q��z���^��~���(l�5���Ğ�0����-N��f�ټ������V}�S_��tY�5ӭ�Z�ڡt��l��&]�����ƞ�z��zc�gю�^�0�A�N���J����ժ����]4�UnVx�S"�A}�#�BW�
t�kh��oD�k�S�;H_��`�$6!MS�X�9:x��Y���Y�bՄӰ�N��z�y��!�e}=��#�q��K���0�QU~�m��ū�ճ�'e�N���UY��"7��x���C=WH	N���`�Q"	9 ���5���+�մ9SE�to֛�"��
�ͨ�"Hw �;���n���n�K��_�6ڔG]�!����]AQ;��t@���V�h�S@��6�C��_$H��I�E���Y��]�U�8�`���a+�����n���R�,mݫ����Q)j�[rb�ԕ;	Y���u�ɴ����L�j����._��аC�/q�ҙ��u|��)@�zA��1�6��W���V���l��W�/�\�AD��5�q��<�v��MK�e.���QpH��}o�x�j�K8��[�^Ađ����fW���������,q�j�K�E%��V�s�g<��x!����ͧR�Q�7��HϠ>.g.>��U�&kם���h��S�Mx!�M�u5�Ds�*/o���a-֝E��Ѧ������}��_u6��,y�4��o�D@��ꎬT�%�;�,��F��k �u����m�%`�b�N�̣����{)�����>Κ��>����zwmg�j��iA�=���ˣS�%*Ra\9s�W%wk;O�&ŝ$e�f�d�6��qQ:�N���ٵ��%`%vt5,��m����dn�';U�����[)>��T'R��Q9b���q�B��*�]�� v���:��Dd�#�*nc
���Ü�e�5[�+��ڳ�vz�v�����C���U:��m+9��p�ط���Z��2C8;o�o�nt�ho:NoD���"���<��ǒ�a��˔UgYb�,R�����Y�oiߜ�Ԡ���]�c�%����l�J�&$bV6ʳ����o|f���Z�e'�{O�_qݝ5t���<R�*����y�iEƪ��5��5����&�R�s���������{yK�c�O�Ԡ���R�P�-熬j�6�M�u��O5	$3�QIr�8��ɩ>,/q�#�w۫~�N$��:��������q�e�_"���XO�g��ͅ�B	{VR�����as[w��t]���_�ä�����-��6x7�)c�A�.���F�䕍,H�lP7�z��
�g�:�Wr�ǂO�mh�k��1��>؂����qv����s���������v֙*Z��k��MP�d�Wz��\�z�7*e�*�3t�8�\w���U��%g�:,�A�>�"`��B*��+�i�a��A�`yX�$�=���n3w�������b}���:���s��b����}���V��Q�1�mr�xyc�[Ւ�΂Q�i��Vmf)��'
O��g��9,�W���d����54��Մ�f�;�px�T'u���+n�e�#�3s�5��ܐ��O��84��������B����wmoK��B7ƍ�BP��S<v�a%�`���Ѷmohg:k*0���Q
�	�o]�(�~�rլ�rP=��89[o�4�r|��g:K܎�j��΅��E_CP�F6Z�(���Ma��Mg�x�i������ھ�j���ްK2�oD�C�x�l��Jlj�ޙ������x��&�1�8�QCy����k����#�C�� ͊BE����^Ӝ�Z)��1�3V���>,Y�����7%��#��J߅S�Wt����iXǅ�^�u3�x����lX�te�,�{��.<�������R���U>��H��^飣:�	��yC�@Q1�m���V��gBx��/����R��G���v�Z�%���Un�ϑ�fT˖��f�\)��/q�I�S+kI��NRm���o{�ϕg�o>5�M#�A#��M�7t��qmp�Pz&)��g�fowbkTP�uF�<��Ҋ�rƫ-���S�G���Z�;[O��ԳzLu7�.���!u]S�凌�������}/p��(�ͨmC�Q��Kzľ.E �X$sw@��<�r�g=����Y����J�ŢT���d@��(�pj$�����UIH4�Rb޿C��Ə��aJ�'�(����h[�x#�����U	��=Y���v��n�3���<�D��Y����Sjh&F���ٱΦ����9Z�W����|����=� �}Y��u��a�<��o j�j����h�#���K+�s#n�N.�c�m�Ia�eFٵ����+����lJ���;-�\��@���Q��k+j��g6Pg&��o��qTE�=��ݾ���n��Ȋ&n_�;�4���
�ѻ�1ɷ���߇]I�Fdm�+��]go2�Q���nTE�zΔN�w%Ř���.�xkOn��G�gQ)`%�\i��È���iu#9�ӮC)ô�a�#�Rl�~m�:Κ��C��J�i���T�Y*M�X�7d�O���9��b�MZ��;s�y��V�O�="^xN�=,���+"0����z�͕�.�L����x9�I�|�N��#�p#C��6ؗ���L�b�*U����auxm7�͵�����-�x��:��'�E���p����W���A�xF�ֱ�0���A�g&7�����}�,��!r�<�����k��K	L�Tv��j���d����ʕ�͍;�Yjc���:��䆔�`�G,-Nl�;���Ar��i����9N�P��7{"��"���5d�j��Wgu�Ʋ�`�*�f�)iF���p��.��ܳ�<!�� �"�$5T�j霛��Z���2P+�I,gd��M�P����h�h[�s�!D��r0W6���yѴ���̬҉��[|��&��1���*���ոO���;���(��#�f���.�;��Ϩtl��ֳrY�a�.Vl��z�ٽ�W�qv�9Q#�c�/k��7�@Y���l��c`�z{�4��������0)6��hHV��{4%g��eİCjSCC���ٝ�X)T����.�ƞꢷ4O@��	y�m����ѽ�}����k�Ҕn����n���F���X+b��o�%�+��藓h�~�dW���蹞Y�c4-���-�WM�*���ξ�y���'J��[�g�7k{|�t�l����o�F��/fTP}�MXR�Z��86XG9[x;y�i۝;����
D%������W$��`��*yX�ItKm�k7�<�;s�V�='��D7v���l�M�,� �t��D1��k�R΍J��nP�{������Q���Y%�A�,3t��;��>�B���A�ޡ��?�k�Eo������:'��jPF�zR��an]d��ɳ�s�;�n�[C�l�Qv[���U��VTt��� �7��*e.Tim_AKJ�7J��++#<k8���U��EδY����c�n�	�YZ��˵s���%I�ZN��\w��Ob瑳3o7�˗A��
I��j�l����i=N7o�{G��Y}Y���O����ұUѡ���V�A�5xߔk�$���7�H~�H7=o��>՞�{+\�A/jV(eb�S�6���(��N�H�W}(�������%�-����!ž[�*k}�V�e����k���Mvsx
�g=��M]�Ci�k��_S���WJ)$�P��U5âG�h��P���':�w��|j��|�K���ǉc%]�wW�j��"��-��W��K_I��>|g�bp9�Y5m"�%s�|E���ڰ���;��T�^��z�N�4��؜��7��.��4�+�A�^�~j.�.g��,׶C�����_rWR㏒�o_��c�mtXgr���>����k���8I;��w� Q�bkD�6�V��`��PG9[x;y^躧�O]K+������R�� 9�%N]bH�ހ���_f��G����wc
�A�]c��ɋ8�gԭ�=V�����֙�6I��˼i�`��%��gd@D�Q{I�o�nF)]�L�+l]Z˵e�]���cf>�"C��9NN�З��GY�f�y�$�N��1A�N��7%pi�XoM5�	�qO�Vk
�8�|�uĥ�Kr�{G�FVoE��:�[*�Sz��o�j#u^�xǒxG �}��s������،P��3b��Z0��nf�kU�f��JYu[�ʘ��7����7%�#�@#��J��]XV,`�fQ*�X�QC�:��5Y�y�4���r��O�ĄS}j��m�U{i͎wTjZ�$��Vd��IO�
^�8�L�S��J���G��C{]HE�WF������XZYX-��"�"�83N'G�>^��tV{�el���܃��_G6yA���k�mڪ���֒�.sM݉K�3�B�4u`�|��֙��O�n��kL�Iuͦ�+Y�qL�NB���9Ԑ�U4�H�te�Û���*���Y����j
��b�CR�Ҡ��NYլ6C:��]27]���nVԔ�$�2����)�t���ŀ:|x6sWL_�lR����=O��ΝlVg#�n�ܓ^�ڸH�X�?J�qbT(4�r<�@y]^�f�^G]ҕ2�j:��<�z� �Ytkp���WJz��]�0i���%���a��ϟMʼP�4�)�{k��x���68�NS�5�,������&!�|y��h�^��l��ni0�xR�Fv^ ʙ�ˣ�nd�r�r�0gXyҎ�I�w���]��1�i�SnΗw1�hվ��a��lfEcxٹ|����>/��Q
�����S %��Fn��۵zR��dl�57rj�T��\mF��}!܉�m�"�n���,�n�]���a�����v*7�N��|�=�����P]�ջ�K�H±q���J�P�%m��{�k�bG/K��ɲ�N�ۗ!��T�#����B�]�}O�[��!y�H�^*�Ks�ۡm�z[�ᴹ���ڔ�t�r�ٽ�*h�q�6�"\�Ǣ�+s[�x���wn*�e̦�e�[,Ku)�'dX��8]��K�ᡍ��)G0�O��Y�j�!��ۄ��J��{�#�NT�*�eC0�Z$ۮ�K���T>k3�0�M�C��o��m�F���5J��t��I��Mq��q�mX��k0AA�'Ώ�z˱իm���4��d����C��J��L7#�rwQ��dX�.n�)�,�֭x�R��6г C�e�]B���E4n�ܣB�sh��y˦�'2����8+��ӊ�@'��s� ���Z�dnG,�y�v�/��U�wF
@i9C�\R�W��0Wk��AX��RseC̍�ǰٻ���������]���q��L�}�nq��hUs=:��P�w��Nu$�q��Lmͫ���]$ޖ�����hZ��:[�pA�ں�5�[�{c�Y �s�Nn����o�kR5�z+iӕ�̦4b� XSM�B�GR�����M��X��S��7���\Vi�gb,�0Y�
Q�Å��f=�t�Ƹ��h&���v��i�� ��B�\�f�ɖM�le���v#C��t��TL�� T�I������� �h���W,9���us���騪l^���ͣ{Ld�v�̂�4����q]��W����,��%�9[Ǖٶn��R�תM���]b���˅�/c;9�[� �g�P�-��p�1A�yђ@/��#������Ǔ0�{����]8�k�B�ʭ5,�a�HV�c�y{/X��,�{n���ɭch���wv���7�٧r�:�0�qUjs��`ܛKw%;�1����g��.���M�[m�d�1;SV�X�;ib˾D�)3&�9]���\�)�:����u���|��%�f����r������������L����i�Ի��7���3���{Z'\�&���30�3׷�F��{z�;1����-W��\Xz�7�����ɚZ�f��D�����{T'���Y,�j�FN�����­^��y��7���kU���;����-�*�;]�oz���S;.�9Ʈ�6���\<��M�SO����p]Gq��k�؝���j�s���{{+i���y�֜y���F��f���g,�:l�c=ky%7���fg1�^��5f�kZ&��z�z�{G%����-[�ou�����)�h�)Yt��i��f˥��ޖ��7Lʠ���u�ِ�O�7��*A�)=;�܄��r�g$�sv���i*yt�a��@����p�FJ��(ޙ���x�jݤ��>�3?W�］p$e��ڰ�������Ъ��8�^b(��D{8&4r[+ҟ�����m�W�O��嗮�#�nT����:�%��V��o��Xgr�ѕ*�|,Ux����I#*��of�W��{E*�㵞��M�epra���ӕ)NN"��=o��q�=`�\u��͉=���N�x+UeS3|z��27mcpe���f;�M��i۝;��2�����Bv��Lf�}�$W.�ۼ-��UNc*���M��󘴚eΝ[�c��;E�،�Xk���ZU�!:B�FĪ��o|f���Z����6�㓲�/^'Q+5B��F���/�K�-(�.�8�e�ga.j���4]�%md��)���_w\���Д�U:����J�����]hZr�"��luC
�B�(I�1�7A��9s���ٷKv��5�Ρʝ���I^|�Y�L'z�U�F3��-ά1:�7�	ʆ�J�����ꇟ6���3%�9�g-�o�#\%�N���0ԝ�2K�I��;�ȯ�X�dt��!7`uY����F[�0�*ȉ=�d��%W<�t;���aj�
W��W�U��gI*h�[*L��r����y*���-��L�%��ȵ�Ey�R9���j�#�����ԱP��I`���E��j�a؎nC�$�R��}WE�-��%/�F�iS]z�@Ȳ��ry�T+x9�3�4�{����g��$J�[�3�*�S�Ǽ�#!��4u�6���fv*�/Ŷ�����W�-�ϓ��&�RqI"��L�����@��	[c<_1�KtDMUv�h��e])`�ݹ���eey-��7o�)�Ru�m�5(8{�V�%�AK46�X}gm���O��&��XOA��xt����\�x��MsԃG�i뷎�Xn����� ۯY-[�ͺ�+O��G4.~�Zo.�͔���|�;NÝ;�Γ���W�_�Ś��hj�v[��ݳ�2���dybn��ӝ��V�ܨU��1r���K�;����Q�:�X�8��	�7�<nAkT�B4��v�^�OWpk�F�`�kV�]�q�Ȱ	��˭�d:�a¯�t�|�u�o$Fھ;��JĦ�^�E�J�4�t�ozi��<�v��8��F9K���q��H��slr���R
7HH�]��W�6��6�b�`v(:��#SG�J	��⓲�F��^��B@�����Y1|�v�%9h��M_%9�_�߹�7���/e磢O�ץn�ץ(�lEA�nۇT��rk�UWl��[�t�\�.�c�Y�
B�QJ`��N�J4�mB�`�Vl�<�̦�ܱ����V|��G��f��"�B���E�i%Ģ�.W��S�o]gK+=�E�ej�YÁ��왝QbzR��aEb25��ڤ*�;z�*������pk� ��W�y�]��(#SD8�ĝ[Cdnh�����g������B%%,��_t��Ӽ ���#M��9��s��B�#UM=yY���,f�W]�:_��n�C����7]�ˡŸ;=2�5m�z�������;U+�9�����!fkI����viG��m<g$JVwJg_d����r�N���Qa��Ohi#q�k���S�U�]�@4�f��Ԩq�l�G=�yK 50n-����eD¢���;U�IeNm�V�z����6��^����<F���J/0M��@��6o��<�7Lf��Ͷor�c�]o���5�B�'��Y��aE��������3�Ҽ�7�w�khߙ������Y��vD'�6ֲ����K��km\�B���|��ǭ̧��Ol#�{�e�z�˻����7�h,"VN�y�*��Xe��{���حjq��+��a�z�J%i~v��ӽ����C���P�U��q����7��܊}�d�K]�|v%'�Z��NV2���bhv�f��AlK�X����M�rUEU��Y�x�ś�`ߛX�9{,th#�!�GMf��]�s���ǎZUcy��Aq���5T��Gɥg�cY�M�1�V�N�Q�Ҵn�t��%����wU�%��:IX9cU��K�d��j�_H��lc����Y�=h���s���m�o��5}�3,Z�K�9��)zro�/�9�ZR�c�mc��*�1Xx�~�)a\1v��q4�Z������q"�q�I�60���jV�H~�Z��f��J�N�Z�Bv�:j����e>��M�X��p�F8��vr�N��j�He]WF�ΖW(,�&땣�¬v��d���}�B<*��Y��)�5T�n��]ܻ����A�%rK
Uq=o�;8Wr����(��(��zh��Pb$;�/'��n�䶵SE\\�8p0��8�s�Ā����EΤ�<1F#B)/y����YU}|�b�a3W��󍷀6�|�V�Kۘ6����J�7xt6���u��Ѧ�;��f�b��xﺐh�Xm���=:#��9~���y����|��ScT'v�V�Ś0�`����ژW�P�8j��{��J�����:j�n$h[Z)F:ZmP�l��؇Ϋv�mubcRY�+�	�����ś٣�=���N�s����rK:!�<�ͷ�j�,��馱7o��Noy�eg��h=�)�K��xؾ��9U1#�+1�����o����\�柶�����}p4,]���;\��-����V	y6c`!d��r�Vx8�L%Wg:i݃�Gc��hS�.G��[Z�i�OU�ιס��Ֆ����x�m`&�7`ǁn�`ڹ�W�%JJ��|%|�-�� :i�����)&Ss�V��F2ݺ(pw*G�t[)�V1@��'��WbU��}ΡE�0m��H�B��3�V�k��-��b�%lS-(����F��3���̩�Œ誽��7�ĵ9nܰw/<#���	A+N�%Ev�jƩ���u�D�mB(g-�m+�+���aj����4$4�Uuz[�j�q૎����c�KҍV[�kE���[*Ľ��d�\�(�!��s]�ZMp�w[
y�Î��"���-�Pl�"�m�w�,��C�[�@ �_9]�K�T�ݖ5�c�X�P3|��s��T+x9�3�5B�C�[7\3/�ַv^����d9�N�3a��A��`��^<�0ڑ��uw�'�Qٳ��f8U����h�T���f�,�v���lB��B׵]b5�u,��;LV4�}ۺg����ʸ�¢ÆJ��	���ʢfȄ�pg%Rt�c�pekśB+��ʜ��cȐ�6ɯ��e�O�8�J�E�Ě��w.>����cpͰ
��"��4��+N��(�9bS�\���W��rD�Ą�jV�e�J�l�����S�jm��Zҷ�pTI��ȩݷ
��ݜ%��v����r��t���O�-�Н�XknN6C�}�G��L��,%��޻x��t�_^�؟x��ZS��������Ie+��թ�7R�!��i����;N��N�w��)h��ɫ�f��QY���J��ȩ*��]�C����;Lr���-��ff�Nr�t�$n��/���C��6l
B�zv�i��3mbѳV(N �:_��kN$�P�a4�x:Z���C���A���J(v5Yx�.[Q��TI 봉Y�{Lr��ń���`k8���y�p	A��ו"����=��"Z��J�a�%j��[�u�&��Ьg&�%r�@K�V
6�Ale��U�Y���h�[N�ק��"���M+�zJ����;=~5���7l�̵[o�E�XW���JR���v�h�σ��S�!���3M\�n@	nH|��ݿJm��Y;Yb[��k����{|[��sjμ�*�n՚i��7�Q��"�٥�1ۛ�2�_�d���@We�=@��۝f�k�$U�Y�k�c=����z����9�K�Wr����TB4�m�ʈ�I��P�7�����v�=z��� �VyC��|��Z�ߛ������^ӛ��\����:��6ۜ9ة�6��-3�;��2�W<�qK��Ԧ�0��Φ�T���g����c�I˅"8N#~�&szͱ����Xm��6�5{7�w5�pu@�6�;����V��uصI^1X�f=�f�W܃@�b�\��_ֳ{�׃EKGg�$��1�oC��T{�3�ӻ}:�Ƿ��gIaߎ��M�޽��b�4o����i�n8=�ju��ګ��͔�M����˹�eÅT5|����l�a�x��Iގ��E(�oEXi�2�h��Q#k��ߔ�|c�t>�z=�޲�q�`܍�$7�[*G�	yص�����f4VJ�������נ6���H}��s�	DI��i���Tw����X&-�RAP���r�c3o��T���gHC�1�lq���뀬�	a�Ic�^��ה�F�2���N�nn�Z��Z��b:��⥽Wt`]�^������WtW%��X�e�i��1j�Mc����F:�mHA�Et��<%*���!|�p������6�c�lsר�M[!��yT���gr�����E9��d�Q��Տ�5Yo>4�H��r2�cٙ�M�qi��[\��ϹB	mWT�v:IY�X�S%ҿ7ܼ�8�j����m�\��+�w�����P[U�'U�2�����Z���2�yJN�!����?{Ed��R
'�j�#��kUU�B��'513�r洣Ui��+89ó�5v%� ��(S@�����:�u���z��x̤����6��ރo9E2�pMyW��׈Tǂ}��.��2�:uv��׀O�er����Kd�.T�*�T6=u�\�L��O�������K<�����՛��Fk�y��A��s\�7�w�z�e�Eb���܅e#�87�0p���>���)W�.A7���!t��r��di�qլV�K��L�ig��B�B��zZ4rܬQ�oe�-JW�}���r�ۣ��c�J�/����[��(������n����ejIJ�_M[��
�u;��ծ����l%�����QY���h�B7��ͣko<gMX7�U8�N��6e]F��w��w��#Iiv`=�����g�7ˎ��5y� ��4R�;M�j��8�_B�sIc	�
U�����,%�-ݷI�:w���ef�M�H�z,�s�&ғ�JK=e�T���gi,4��t�y�Z�Ӱ�N��z����K7�Dd���-$�T?`���tţ�ƪ��oG��X9�Z���"����Ѷjz�e��e�:��7�LH�-�T�GA�g���l�S���iE��_B�j96۹y ��J	]S��}H7&�ZMs��˿��-��G-��S�M�Я��M���X)�k�CJ�6A�'dA�g�|�%P��)����t����n�E��E �P�>4frgX�z�π����+�'�K5t��v��W(�p��5�\��`:pn�|���AbU��B,R�g4�y����N��dc4��E��b���Uf�[�էUVsN\Wυ�����}�����K���*A�)V�[%��$��2��uN��m���H��Ϝdqz��G�b��]�WWs�*�<�N���'F�(�F�ݨe��Vf�^*V�q0.k�.f����t{aV���o7�ѴM�|:�$4�bV*�x%x��EB��0��ܓ'�)ƭ�)_�.�i2D�5]]��\�_��`��Gp��w>�	��������9*�mv�4aݱ��(M@ɑkX+^�Z}�������'P�w�1]�;�VŇk?�\0�^�!��)!�_f�7o���R7����HLB�\��A�7���S3�a����аN	f�x4+NY
ۮ��,W�&�wc/���yv�r�q���Y��r�H��]Ǯ�(f�.� �XӪ֟e��m��H�@+GF�t
@� �4ڣ{lv��Ь����Ƣ�O=j�l���������6侽�:h����/%�]=�G�z�d��݃��wD[X�lw[X�tb��J`����������K�h�8�'Z0Q�b�Z_a���Y�N�Q#ݳӕ�ӥ.�1z&D��f]��u�<�[V��ãG�y*\o$]ro-%���r%�C[�5��8�ے�=�n�a�#.t�j�Nv3�{C���>G���Y��e��I�G���M�w��|�@�:���g�=��i��9��z��`\��Ùu>�z�T6�agg+u@��F��͢��:a�V^���7�ݶv�9�l�6�4��C5��j����P]d��L_=)�ޱ����Y�O��M���LP�f����#8�㙒Kmm%|u�ˏ�M�ѓF�8�r�*\�쬔��p�y[��V�>L3O��z/<�\Q�t>�G�|QPԱ��ۺ5in�h�J�Cy:�^)��Ϟ%\p� ^I�`�h��Sܺ��b�&U6��M`#z��-���tl���ٝ�]�*h<E���#hZ��N��iX�F^;��2��[��p�KB�3v���)л//.U;ۙ�J�U�dR]<���2ӵ�-��d�O/v��nc�h� �ⵀf���7)x�gI���[���b�u�ШUĢ��CN�U���!�vo
z)���&�
�I7ۉCm�U���Lj@��F���F��t�2��oR�vM�_u�&�\9U�c�>Ht�6��e�L<�t���GDZ��1�>������G(�=pi�GR�zaJ�Oh��o����k3��dD~s��Z�lI����A膧��QY�)\�j�� U	O;������6Sf��S(�?� �>�Ծ�ó�ueA�N#hJ�s_j�&5w�b:���s<s#�u��]y+%�ޑ��{��/�ܤM���%��������R���f��i�9Y)*��&,��_��oi�z�����y�{{5��֕��6�mk]��ƅ.������ї-����
�!k�]瞮ުf��L:+���f�fV��i�s!k�Vf��64q��uh�U�2���%X!d���:��9���-4�������``��%̴�MT5�1{�z�����皹��Ѳ�.�G���R҈ժ�imVVY�YR�V֥�]�i���mLl���ٖcUs[Zi�i��L�YV]b��V�SZ����i8���y�gK�Uٙ���ʵu
�TT֪�&�z��3�W�	��Y�2�e��VZ�f�,�r�Y���-���KF���-&s�]��^�b�#9V�T���������F+�MKW���͌����6r�KVV�Z�z�Θ�Ջy�Nz���<X�/Zr$�(|
&���Dѣ�nl�Ӹ;,fԥ(�5�� p�\5�m�O���hL�-�bͥP��ok��n��t�Wy{!��@���c�R�0RSZ�K����_*�ҋ���E��j�K8������Uw+S��k��Qe	��B�/����*����z�@Y"5ѹ75ǚ��%���z��Fp�SOVVn7;���X8�y��ښ����]��V"U�K�=A���RC�j��=�Z��;}��V;,��h�!���+2O����=���y��.�G�N��	�+G�}/i_�[)xd	I��i�GIA��B�\��_y�tՃq:�/�f�y13ڞ��h�h�b��]�4��a��m���v�����y����m2[�8�x��w:+Ք�OY[K*Y�Ar�+o;n�.t�u����٨��f�I$��08��[DS���¤�2�����������7��R���9��$�d����RzJ���!�~�-�rU��n�b�d�Qq{W�g*��	�}����|-?-���5�"Pimi=YQt����Lʴ��yD)W�ZRuu�g�9wl
�+A��K��F�Ƭ�N|�#�t��-���{F���4*nn�41��"�DJGAے��8̾m<�*+�'W7wct����
/UOW>1�=��{�-[�mM!>��\v(�ueӜ�榛�JYuLe�sư�����z�'%���4��ș��tKU�=ͱڑ�J��'�W�bo�j�[�u�M+/�X�rlbW+r��>Sq�����^�~�|�Եw�VX��-����Z}��d��gF���kW��\�C2G{]H��v^��t����ť�E�o�9�"���Pks_�^��A�AA�YH�����9sP�������C��x�{��H\曻��1�b7�T׈Q pn������2�++�Km���,��bK�mS�XqO���	��=�ls��B���i��-���A�)#t�����m�|ņܽᕭ^����%M�,�F��U��S�*�xNY�3�m�y܃�����\�.Y�O���4 ���Ĭ>���k����h4%A�Ѣ2`��.[��],u5�ֻ��+�cV|yC+�Ƨ�1�'��n0#��V��{�.���%�jM�㧵�u�c��(Ws36#@:r͑�;��Fk\2��<���f�]y��JQe��.�9����0����G0߅%���&�z���{c�Βðwm`MWps�hFŉʭUe㜲��m]�of�\ItJ�N�X+j��a�ܭ���s7��J�vѵ��2��\�����/��9�sz(<�)W�i�U4уGhLL҃p�t��%v`���4�����No����>�����f*���n{.�M��7J�ߵ[lĴ��Vi������:w^Tfz:o���Ǹ���,�u�D6�`�g�oY�~mc�/e��NNW<�=ɢ�C�c�X&��p�`�.�|���o>4�H�
��>���y��٦RI]Կwu�B���U�%���Vrƪ�.���<Ә�n�n3l�Ԓ��|�_*�X� ���T$2�Uu	�w�ʓ)������T�rķ����|���l���[���^A�|��{�V�꛱']�$U�7���li�����ط����F�g��y���_�.���k�����uu:�7u�ч��9��[3�f�j��_	�P<;4p�J�;�S�v�a�=�c��V�܏�p5x�L�҅���N]�X�M]򩵲��i�0�#�sX
RX9A���;8WXa؂
��O�*�\�(ӆE<�K[8�J���d�x�c���S9��SCC���{���d���KÛ��죯f�'5���y�������ڥS�E�b�-j�I�H��|jHS��q��
͡����x� ��^�Rt���T䣃fy����|�^أ^��v�V�1nlu��bw�ؐ�VjJ�B~oo�6��km���q��\㵕��F�Ν;#�G��6R�4_I��÷�ۣ���YΚ��C�)`��}�O.�����N�U�e��,��A.�h�7m�d9ӽ��+�`3�M����R���֒�)��*h�ʿ��%��M7�ūM;t�u��*��y�k+T�[��� �n��ccU��h͵��-6��IW��i����!�fy0Gڛ���v�ork��]L�W����,J
b��A�z�,ǧ*�S�W\θ�KEء(�"�q�Z\�+�M7�=�f�;�{��s��L�/�!Jmo&{�휇��P������cq8T�\$��i�U&�'����8���tH#� ��-(��]a�jW nC;&�J9��J�Q����v5Ƴ�۩d��9(%uN�%Du��[%��b��9z�/�UY}�ʝ�]S%=���Z�t-+�h	.��t�����e���.{.�SY�XZ�-���ʹ{�w�-k����7������e�9��~�f��C,��9ȼZ-��gx#3UE�E��^u�5�+�����]�()�SG9��*��8�q5�m�<ёѕ�
�Q�o�0E��"��Mㆬ�z�
ͬnk�3�VqxɮT)�e�����<d���74��C���hꃣ/�t^I��č�g޲�䲧:��m/��ۚo���_Iu;�k��XOL5��IڳsO���5$]�f���<@%c�u�k����}�5f�}�n��0wF)e�b5����:�!t��������M�VʝA[w�٢SQ���%lw��sx�揁Jnt�e��Nܼ�(�d���ۚ��!3�sf�N�����۰�N�,�w���*N{OkL�F)�I�;u� A�x@�uxY��d�M����1�v�����av*O��[v��3�4F>���"�h�|��f����uZ�VҼ�g���m�|��v�Q��ig%I���4r���Γ�z$P[@J�;M�IV0�]�ؖj*�v�om��ʬ���J%iTKS�V�='<�&�m	��!��~�vn��P��Mj�r���m�ū�X�k���:��!lR�*�[��OZ}|�D��Ư�Y�,$�5��NK1�}�LpYʧsJ8�JJ�o1T�IqC���ڥ�yγɥe�+�ro�^q\d3�9]E�$�M2�D7�hHI��	j�t���4��t��'ڳc�f�tLѪ����|R�~��W�r�P9�Z��K+9Ah���4S�mE��Ƿ��D���9k�`���A�!��#�X����A{�I���է�N�.��S�9T�;����	�v�5yNU��a�&�h�V�vd;KL���7�q���ŻK�p����6 �Σ�Q�J$���^��ȥ�nrMyn�ܵe��ā�p�[�͒�56��d�aL�!��.Ƚ�Y���)���&���9C����KCC�
��O�h��PХ:e�23�0#�/s�U�K�q�Y����g���&���&�9��*te΋���>��x�f�Ӳ�C�4.�+Λ�j��m��ۚ{�jڽ�^�~������ϜtG�4]���w��m�xu��b�m����y0-�Ƌ��w�i$J+ni����m{BU;��կ1�6�:	a�ݴ�"fn�����kU�ȴ���2w�{�G���b�BD��v�
ګ�����*�V�˚������8���^QOɫN��	�㡜��x*�[K�^�[�����ms�Q��-Wi�$7�4�y7��d:w��ef�M����[O0�Y�5HIԜ��6����u�U��KHbզ���o���B;��}�FsI�g��P�,qt��1ؕY���ư�gY�ٴ�B�E�r�ck�='L����^ �1����B���3RV���
�*����e����Ǜmf��t�/shQ�um��Ԯ ���ƛ�4��3)�rǔ�ZոC�"4m��-J�ԅ��̕��b�6�y��v��a�qW	��v���6�R2N/U�%��o�N���]|��"�|kKp�^Qer5��'�?���Hg9������	mWP����G,j�3p�����[}:�/�QIIC9e?[J��j�s��Z����,�ҙ�V8"���G4	�KҍV^�r/ť�L�/p�n�J�#�Q>CU	ٺ�юe�.�F�z�(�c{.��[�Pl�(vSTD����E9��:�A����'F&yIԟ�D�E�;{�;y�qL�q>Mx!���9��+^�7h��l�4��z�4�ef�74/;��qL[jTe�1�oOS��Ŧq�D�*�u��U<�#U{	����P>�W�t��oxmv��
e������!�:M9��^|jn�n�v�
�Y�f�f�8���p�k��ZI-ٲ0����&��mm���7�T'���t�oj"�q����\�w{��>� �u�W"�R,R�լ��кɨ�o3��ns�
�-P��@������!�3�X����T�R6w��ai�:y��Ȧ;�v6ї�eΉ۩ÏP��֫�"�VP·X&%wS)P<4���羪z�=H�&�L�g����g:j�lI}JW���Yy{���J�}
Iu��.�͖�:i��nۤ�gf��2�-�{�Z��otV�K+6���*���*��Y�M����E4�d%�\ilS�y#ww��8���BC`ؤ&ъ�U���ʹ���<��U*5y�SԔX�(�(�a��X#�|G��͊bE��}��JaY���y.���o�x}<�j�sͻ��GA���T���o��k���e+��ע���I&G�[%�d�Ј�rmj�-�z,��یc��Q)�[,ꁙLU��Dr����YX-�~��p7{!k�n�Ӯˮ�ǽE�3+���Ȥ?`̩��7��t��89���%�|�EA؞�2��kM$��?�"�1>#U	�ՀPs|��6J�o=�)��*BS w���86�GM�n�����*C���'��R+���c���e�F��J��)�pV(/�յ�s*�,o�7J�m�2�q�P�K;���tqvs��3���ա��m��9G��zsy�w
��w!kc���ݱY�ʨ�>=D��p�51����h�r�u�ч ���p���M=S{m���U�,!���r:f�AD�IU�&�"���Ma�Ύu4u@�U�nouUF;���c�e�����R��oϽ��L`/��ۚ�{}�����hpu@�3k1��t�U�5�i^M��Ƕ3l�J�����X}go<�:h�OJ�dg�qG7T�Ԩ-�	�+N�v�E��B�^�'A9���1�V��G�5���R�t�%]K���r���Z��'gKiS��l�×���t�މ���E*���
ᆒ�t�o�JQ� �f���^"�-kMb��7q'��](vԆ͊BE������ssۄ��-����zf��)c�S�� rvP��;hHA��ݓ\��ⲡ���kT����RoP}�R�Z����5�O�$�	'���$�Ԑ�$��!$ I*BH@�~�B����$��BH@�~�B���IO�!$ I?����$��$�	'd$�	%HIMB����$�����$�d$�	'�!$ I?y	!I�HIO�$�	'�����)����L����8(���1&m��J�I��R$��%����R�N�H�P�J�IEBH�B*�T(�)BP$�B�T�E"(H�JT�fL��P2�����l�4-YQ��M�Z�Xf���̕cSm��m�-jiSJ�f�mm)T�2ةL�UV̭j�Te��{���jYl�R65��T�*m���,����el��`SSm&�֚Rm�$
M)�ɘŅ��5�f��MfԖ�i�֫M]�9��F�lW�  vOSѻiK\�n�˦��*�:�v�ws7IJ%ԝ�YԺ��V��8P]n�tۤ� !v�����[�	���Z��\p�:t�S7M�4Yk*�KRQ�DҖ�   ǽ�h
m�n��[�Vu�r9m�v++]:���u�Q�F�j����K��Vܡ�AL˸i]��-i� �5t�뭦�P6G"�e6��m[h��j���   =�=]��:V؝]�rQ���sv��݅5��Uۥ�m�ت�Hi��+�K�λql5�Tps�(P�B�
-ɸ( (P�@�6��СB�
(=��Ռ��[Y--�ڳkff��   =(P��(P�z�(P�B�
(wx��� P�B�;�xQB�(P�CΞ𦴩:��tb�c��YH�t5gu3�\]�4�rbP5F���s�j���u;�f�24TUU"��J���   ��+��m���i�h;� st����n�t\� �+��Uu��� �NQҨ�M���B���LT3f"ͱ�%f�   x
^��n�N�j7vۃF�FtU�wC� ���їTlw��GwPPun�E����A�U]�d�V�Y5Umk5�kl��  �EyӀ%�'r�T6��(��v�kRc 
a�.�u�4e�\ QI�����3�hmH!�6`�Ͳ<  <k@���h��s�U[�erTWln���ZT�n��QC��J�Ó���U���WKm���7v��wY�M-�IN��hd�
�ZFj��Z2mm��0���  ��z]��.���6�J ݷ;8ӮڒP��⚩uvN3�U�B�n��t�q�Λ��v�m]]�:H��CZ
�ݶݦ�R���7Xkk[+6��I�-Hdժo   �=km��w5�5m%�,ꮭ�N�wU�v��wrӍ(�N�u\]�ڭ��*nt��l�j�f��
�Ӭ���:���q�i�;(nx��T��  Oh�JRSDa0 �ښd�@ �J�OQ�0��)R� &L	4�eR�� C�!�v�Ģ
(f��� 13Uʠ)+&k��;��9�v,��j����}����C��?���$�B		�H@����$��$�	"B		��L���KM%v��@Z��;�jk�jL,���r*������{�d&��zݜ�ۼKrdԨaA감wc8%Z��f��u�P�^n�F�ZS���.��sk0o��fH�8���FV4V�5���nl�8�����hu5
�jTp+�ö�B�����
M��8f��b�2t���ţ~R��&4C���`S�i���C0=�7[6�� �p�v�-������Z��L��$��h�~*L��5P�V�F��u>ۨ��f��ͼL��̖V�A�k1M�5���*K��sv����hgNS����s�A��ڲE
�h*��F�)�l����BRCJ)Kswi�E�.�O@��F�ө'�B�h���׺�Ѣ�%�����pAgzc���H�[P��*�=� l��$7l�)֚Ҩ6�=X�)X�7�d֫�v�*���@��	`�����t5-Y�eLЕ�[!H�l�a��.婦)��R�f#�N���EK%��YV�C�3c���*dۛb\[XN�LЮ�k��j
YA�kc5�#$��O6�
I⤆�ŷd=Y�Y�;�-AKĞ:� �`X�&�	�^��R�Y@��WCj$�Ӳm9E=@� �0�����^�̉Ke�������Z�d��.-QH���2 J��QʛFg�*���8.ƀ�(�n�i��զ�I{�m�MǯhƆ�wvn
�����#%�Qkmeֶ�a_���@n�qi���,F�:q3`��4[mPQ*D���ĵ��e�YeXX���t��B.�Y�a��5tqf�t�u�wpP)��,�o#�WxUb�(��U[Sb F��î����3V�Уx*�(7�Iܣ�U �ff��M-�ܼ��Yęݎ��\�_����X�Uت��7����U��F���<f��RA[�K���C��q��X7z��V�eYi�HfX�-�9NeZw>�F��#kj�ă63�.��Pؽ7e�u�E"N�&��M[ר�-�ނm�A����
�#�@�%��nV@�W��]�J-���X��s��2QV�1X�ɶ.#R�e��=jὢ��qj�)#�2��ǹD���]��*�`0!V��6�m����L,+��oc����]n!T��{���ئjcq<q�AR�C0�8�U�f��\[P#bX֫@4�]�r9D�[�H�$O��WC��+�3S8)��om]�߃�SR�Q-��(��n�q�\&�5,(����[�դ 5�ʴ�+l-3r;w+R��ƓF��A���n�ժ��E�dL�U6![FE5���El�J+[�Si[i���m1�*@��,T��-K��ٕ����[Vܴ	L[�n쬆� ����uDfZԴVmW>D�q�r�K�O�Q�YqʱL ��ۥ"	�����
I��4T��@��K �w��+�j���i���	*���v�˱Ej�e�(�ՆNX,��VwFQQ�Q�����c�.�S���/Z���<�h�u
vh!{R��X�F�V~���.�k�*���G�ˠL:0�����&$�TV��_	��']�Uu#�t����Aٳu�HfKw`�zÆ�i���y���Qg�F����n] ��9�FV۴�4�e�;+,x��uvڧyvsW}Ϯ�k�e��¡U)�3^mj7c��-�Z�����Ϭ����o]�D��rEPݳ�!xޑ�|�L�CM��i�y1CJ�mn�c�͂�˫C2:'j9z����&��I�CT9�e�,�U2$r� қ�O2W�aNV=�4�Q,\�U�%��q���ch�WU�*l����l#0a�f��HV�zkDѫ3�3F�Z\
�]<ͧ�CYm�6�!1$�,���*g$*�,(�L�N� sA����AE�c5�Ov2��A  +���Z��*�l՗�����M�F�5�,c����#7"!��:J�l��+7f͸+B�H�
N�m�*�Y�[gI#U
��3v��Ъ�@LN°.�췆�{�*��DS�yL*��;�|J�2�:�Gi���3KjQVG�Xǁ`�B����nn�j��Yh FB�Դ����nS�7[RF�o��ƫ�%x�۫t��[:�j��kXD'6[��f%Gh+	 ���\�40�r͝b�k]��jRmZX���p�6*�m�{shX��4&PE��3�ʗ�ȎfL�&h���%Dk[ ��ݗ��cД ���;(���qT�� �H�2�#W˽xp����^�ts� �f;��mѲRy>J ��pZ��e��[�YR�u(E��n`y�j�n�����U`:���#f�(�&������^�f�ז�E:#2�P��\�'fD�wf�,i-�)��x��1V���3��SWL��ae�y`���ט��koqU�4����L,{��!'���e��"�]"Mmm7�jPzgQ�P�[�ԇ0ŗ�#;���e�U��4�$�BĄ�ݧ��i܌!E�h���eK��f�J�#(X�t��1�hPVN�ZCV�tfu֦��r�~Ǣ�<l���xօPAņ�n��l�f���Y���Q_C��b$Ǧ§z�6�u�R'w�v�x����U�nn�{"ە���/`V.�7p�L�4v�H�LR36Ң�6��y�BR���G�=����<�B�d��G�m��XڼCU�mAt2������ �%��J�z�J�a��7P�"����h��4^�V�u�&����sD��a�P��.��'�Ѵ6��/Z�z��հ�	�J��l��^Ih�P 4]�q5�f�!���Xa �+�u�iB]$�6�ͶF��#�JTdOr7Y���K��+FU�Yz[tt�2�[��X�":�1+q�E�,��s"�O,��U�~T*T�2��A��e��l'eVZ$S3t^K��-%d��^�ʍ�\B�H��N^؉kzP8�GfCPE��N���l��h-i+��;N�`k�@zh��s4��(�kh�h��@۽yK� �	�r�ּR�2��00��m�\9
�n��M��B�&�9��K� �Xr����8`Vm`%j��?��,�Aӗ�(ǩQ5�M�3����k7吔�V�ǸP�5�U�yzEM���4L��/�`�e,�F"�۩Eǅ���c)n\�����e�6���j8/(��i�u��K0}���F�M����v�	��
�T�����]l�l�(���P�@�7���a���m�n�2����ʖ��j�\.�`y.��q�'�Z්U�v�a��ڷv�K�h*T�ڑa�z/q-f:ɕ�����ͼŒ��ˬ�Ju)8,@Gʘ�&�D��ڒ�n+ijb�xC��I����@-�4�ۭ��{V��&�YWW�*���Yt�����f�Ʉ,��<J��V�1N��5[{x�iۦ�"��S�!�������t�� �)�i��V�y�a�;�\!�f�#�Ф�Pр�Fn�M(6I%6�2*���b�C7��M*`�z�mk�w�B���2c�]�(��h=��Z�[�s@ h�z4���)Z%�ST����R��i����3n��w��P��B�[m��;/o>�J��V� �Z��T�����"�����ʺ�+OɃ��Ws%S**ۍ�t �e�Z��"�AjU�a�&R���ض�`;�"�6Rݖ�(Q�s(�+J��$s <� �bq���t���3h�+)���C�v�h�O*�7rj�9q��Z1 ,R��p���sj�
�8%���nu{�L���Z櫔qG�qQ�mKxn�+9��V���U�S2��G$pM���潭��P�A�5.�-�kZ[�n��N��#U������9wyZeYi%C)Օ�]_$Lq#��J�"��	�Co(k�sV`ēSZ�`,ɄJ��@h��y�^��}�[� o�i{�E)���&�効[F�ԥSYz�@巁֚h���՛�S�!�> �5�V���+ٰИ�l���x-�KD�ySv�L�YR�T�'���J6��ķX�id����H�o���H�xŬƴڽ+ D@ej��1�h'�3iGAi�+p]Ad���e��P T��ɒ�؂�Q�C.$��[?�+�vtdY�,�*6pj����%'�rW��2�mq�N=�@#Gr,��ǂ�d�;�W�#���(��WM�b�x���K*��Xԫn�Y5"-aV�ڛ��+�0� ��Շ7d��Fb���ӣ2�$N�Y�Hc��98eoڎP�K�e�h�(^�KQ.�ͬ�$Ct�>i�J�vw�T4:
`qF��`�1�𨥨�bl�W�Le<�$�J�{Ec�4��1^E��m��p���oԳ��J�ҁr�Z�
�Śhco.��#H�2[�tf�W�CIͺű�f�kk����(�v�p<S4T�2�\�SӔvQ��E+��R`�@�tl���St�"i�LVy��M�t�V�S�͙%��,��c�2-*]�Q��L���6n��)�6$�E�t*fe�U�&�B[����m5	�f���{B��6�m�c�5V��U��d����iҢ�L8>�ە5��mg�ô�X��oJ�Skos(�M�µ��]�*B�a��a�{{� ����ը髠i��["B-iV�1�p��\�.ӭ�]���o)�!����ai�s)5�r��B�(�Jx0��Ӭ�vS"�Ğ����͕�O�/
s��dT�n͠�P��%l[fUbr��Hk)9��O:FP���ʻ4�+�y��N9W$����$��{z6y�T��Bx,Жu�%JVX��?���n�4�0AONmlյrVlT�S-ޭ�p��[I�:VV���g2f`�:X�n�h�U�ۺ�)[z��M2t^ּ!8t�Sbި,Y�����J��Z1�(�s\�[%ٕ1`�"���m��hP��7��0���ԳE`U�R�u�(3�;�S�+B!��`N�vWm"r%,���2m��"tS[Z0�%�£/sZ���z���܍�O*�Xrӑѡ��D#q�yw��X��n��J�nj�Z�cET���3B+����+���<����U�Ԕ���Y�J�b�ڧ��& +t�.�3�4�\��P�;a7��D����M$콧��ƕZ���R��/!v���
j�Y����`D�H�y�ۻt�ɭ�)�/.u���"ؽ"E/U�(2��)�*؅��
�ፈ�lزd�,K"�=7P�#NQ��(}e$�����kn�,��$�R�L�Uw�cIrM�L�W�b���d?���V��5*���x�7R����zؔ�V��I��J�q-�u/v�L]�M�2ѣ�6=̅����Ú�-sf��)�41���d`k2�5�mn�<P�Ԝ6�
�����4���Ba�,g�^ۇ�E7Rf�{a��[Wz�[ãi�c�[	��mC$ی�Q٣{�Qk#Y���x������nf���6�E�k�BH�x�ˠc�Ò���4%�If6��C�f���Ih��!+q�ˤ���e,<�+5��	�lr��ٓm%��<Ѻ���6�̠�9�P9�.k�P;���Ue�ܢ��b�i�����A6�P;�p�z0��e�Gn�����{0b@�<����i�
׶m�Bvj��ͥAD�j�!��)Vj�e�Cf�,BU]��:t������TyW��(�R�~
��ovBf����vQB:i���Jk�6��a�"���^[5��%kJ�3/�YVX���SR�ʔZԕi�]�vhEW,���i���f�F|V9`��yb��-m��bL'N,�V�&|N`�iU`z�S[O�/�M�d���p��*Hű�.��p2btl+�:P��C�bʍ%��=�&�ޚYU1�)�F�C��312������B4��ݫ�N�.�V��Y0Q�Mڤ��mٳ���
�;�̀Q7h�n��J�%��ۄ�E4�4or�R��b�9r<h@��}/*M
�ذ2V����Ӣ�W��l��O��P%��x*���Rm�v�V���T����w%�f�=l픩+iP�V��%
�_n3ET�&��E��0R�%V�����աt�*r�ݽ�^&�� ņSl6�8���hCX�Ə��IR��6�`/�+V2�Ǌ���ܬ��h�n��3i+�В��j�&�3\���$�f6�H��m�T�ۼ�
�T2��!�Ĵ�3$�o4��*n��Ѯ,mdMXh�ՠ�q��a �(R�R�Y59B���&Cz�1aY��&g#y 6�Y@�[ݔ���[�b��T�.�<�.�(%q��U+L4ޱ�R5OV��1I�a��fh���*��j�C���hj�,�f��I�pӕ�a�)��X���� 5�X4)2%���|`���c�T�Ib����r]��	PÛGN�'�=�y+�_1�`X�Z�6V-����ճz�v�@�)Id1Q���^��#4L�$���wm�w3ex�k7 �%���y��L�q��P�Vc�L,��t�cl��#u	Pڻ��\�a,rJ݅V�`�CLۻ��v	�*�ֆ�32���"���ҭ��S��Zq�tCô���-Qg,���M}����DkZ�
������ò1^e��E���� זbF�?��ћ���Q9��F���+�5Yr=U���5����`*�V
,�X��i��U��Rz�V�v�;z�h�6�u���
�%+�F�N��0�rn$f(��VG�]�)/uL�n�O�P��*�롻�ʵ�Ws��Ru��e̥�6���s�幐����wc�p�Xe�]n�
Qq�9k���I%u�1Y����x9e�t^eZ�/ )u��8�4��������1�9e��m�
�GA�Rb�
�XΙܪ�b͠�w��>4��p�3����Z����V�e�u:��\�]T��*���u��:w����<m�������n����o�#����B��oIL����1lq��sV�ӹ3���r>��)μ .Qڵg�V�2�lݠ~�tm�X׳���y3���	х���|4c!��x���'\�B:�����K�۱��m�r�#�,5��P:�e���n(���J9���ֆ��L�E�*�2��/��K+�w=�7Cv�Xý�v�3'��*'] ���al�y�R�`w˂n��Oi�0d���y���ݫH\�Nf�1�t��]����wq���j��W�U��Ǖ��pn�>�Ȧa�Ѯ�Vݺt�Vr���Ì4���V�	�[��<��a��$9���MC�f���rB�� {W����Й�j� �&J�����}��s����4��>��A��К�Gİ����k��J�����L�u��m���2�&�T�n���b�f;�`wy"�;��p(�z�6(�5�Լ'�2�v���G����&�o&+(�Tް:���l���ʛTxU��8��,��G)�Ugu�n��4c��x	ސ'#��0$97gY��FɅ^�i�,��F����l�^��J$)Kzː`5o�YIa�;"H����d�2�Ϝi��t�vQ$݀�м�n�<z2]�bէ��5鷀@��{
c{��LÎ���eN����-7,��9�r���x�h����ָ�!'�:�V'�q=�bu�TOr�u��kా�985[w��<�Qjk.��b�ŵ`U��Nv���=�w7O��EA�$�+.$�.mk�im蟓��D���_Y���#����Q0�2�c<�A���|!��+�����C՚��Y�*0r�_�X�44�Mo6`���E-R{wpNլ�P�>K���@0!���S�n��O�\��U�O�V��/���8��>H�����r��-�vԋܥ�0^*}ZQ�G%��֚�Z��f��tE�	�Lg��b.�	yIo[�F�
@\�]m4���K�fk�9�y@��uM�ث�X��%7��,�\n�+����-ʃ"�@Vh�/h��Es���D_T@�g|�Ծ;u�!]���Vݻ��5��WιH�1�f���x[�F���,����R�@8vr�M�i�)ֶ���Ц��T�9]�fu^
	nTJN�^�*;������f���=����'|�++Z��ɒ�f'�Ȼ��-�äq�<&�.��8mrR��W��������u;Z����/G�c*���M��i�X2��K��KqA�3F�2���T7�jꄫ���n�1͹r!oFV�a����C������;�8��ql��$N��������|���a��Jأ�����VwJ��kw��I�g���-�qS�|˅�Z��V�u�,&8���T��N�C�������f�����ܶ3�	Qq}�G�ਜ਼/�R�5�pwה䑽wW�]Ͱ��|� 1V ��	�U�dWd�K����s�E�c��|��=�.�'%v%��ٸ�(*n�=,K4w�)SPl�*��f+<����`2��1�n���h��S䮳����8;�5�-�,%y+{�[6�)��U����e�A|�Lw˳�3�Ax���PVԦ變�(�}�ݺ�3��;��M��M.�S,��,���1t;/kS��Kt��E_9��6�/�l{N����������q<b-"3bJ���|����J�gf6wz�%_%g��{�}ٳ�>Dn^�����
wP|��͍<���B�Y<Ǯ��.�Y��,u:��2E��k�e�.�y�l���e� ����p��yM���P1�[��zcVVm��%f�J�h�c��E�SYVc�������rޗn[�J�� W{2I���x�U�4e��Y�t�u3�h骓}��u��
�N��w
,���-!ep��B��<��Ւ��r���"Wt�1Sm`��k�a�D�9�I���Y�����
9�[0�.��Yx��:��Tc&�Ƣ��S뎜��;;��ƱK�qg`��G��9{Ҡ�c��$�Ĭbo%�)��᝺�
KX�^f����U�Qڹf+:��=3s�h����ui����f`Z���k���n}gZ}3e�m��b�pw��c\����}�wd����&���,ΰ�5��n��R�h�b��7b"�O_Q|��辖8]�9�S������3(Y���tI>��Z�����Pұ5�E�[���Ya����C�^sGj�nD~�,��kA�[��.�������Y�-uPQ����K�����]%eΉ�����9�2��}���绢Z(1.[�6�Z��r�qt���M%�/���
⒬�]p[l�����#�U�ٛ"�Sz�W)sQ�T��0s]�3D��e��TTݸ��|��p���O���A�l��˝��oِ���8�ԃ�ިw��� �j�P-9D���-ɒ��V��Lb���c�����m����q����FQ��H�w��jR{���my�Vw�����e37��Fm?x�˩����a�P�rr�|�\v1s�U�Xݍ��t� *ݲ��O�2�!+=�wP��9�A}zN
G�2�VL�&M[F�Ƶws9[�����M�m�I(����M�eD�+�Z6�����D��s8f �Z@�HF�r�]:A��p�.+��1j�L1ZN��u�$W%1�0r]��dz�}��V��s��4A�N�0�)�;��ˮ�gJ�#b�R�n],o*q*b��&���7U�<�o(ю�XSC�$h��yS�)�U�+��ߙ��)��`�YMr7���h�e��d��lb�
(Ps^,��(������8�u|Lb�m�6T��:$C;�4p�RZ�y���'�{��u��-m���k^U��i��[+�H�=e���F3/{y-'��2�M�z혔�N��y�Nu�gIyB�aP��a�W]x�]�@\ul��FgN��i�qw����;1� �ӊ�E[d��QoRꚫUZ~ó��,�֎�}"�W��HNnбG��Mq��z!�j�� {k����%̇6ո�o���u-�G�(���M��{��R�z=���gf2d�dVV覜�_<5���0�:L����Ӫ�B>�t2��6Z�9��@��Dt�풮a *��Ш���R���Y�%2\��K�)8v<`��-���.�,��,rvm�.?]k�Fu��E�Ot6ə���*��V-t�${�k)�e�s��%�9�2di����9�}P�����V.�[�F^V<;f2�,Թ�0O(E�*���͗��j���׆�)6��V�-$^��>;.�ܩ0���<Qj�]�B��뵺��Ծs`������y���[:����b��i���#�v�;b"�3�1o�'+��ұݣzHW	����b���~xf5Q�*$B�J*�l1�܂�)��[�j�`ל���-������M՘��C�;��{��2۾j]onG����|���x+�o�1p�,qW��d�ҵN����C�8Y-�#B@��З&}y�1k�%�q���X�m�t1�}�ճBՋ�K�Z�xxĝ���m���v�",q�FfܟT?@��X�X�M�����BSU�z�"�'c%pd`�܍
0��k �I��K�Z�HJ1Q�9��yvL\���)RtML�ɮ�k6��F�8����/ʐ&���9:w�d��!�j������m�=π���Rs�bnuѲ��X��`_a9�/0�m�V'F�%�)N���fWpB�T����	4�1�4�t�,���x2�u�ѥ�M�雀p�G6�*U�,5Sܤ�:�4���8��]�9��.7�nJ]WhY}n�"Q]�5f
lts �\��C�z����;6�o��U�P��2�o�q�0Q��-��X�l�ծ���2�[��uVl7�\���\����st��5�\A{B;���$K��{����j�:�
���h7��8Hf���h�^���"LJ�Î������k���nnr��I���ɝ�a���̥O�**2u	�x�2=����-+�ըm<�^�2��p����wi�{�8m�[��%�Z��ASԩS��1��Y�GN.0ė���B�K��8	Q5�s�TKY�����:��.u�q8�.���'ahWZ�믜9�v�r��GC�c{��	Z(���6�=�0!Ի%���p ̇�;�`:Vj
��+H!�Q�[��miܑ	!�����A��Ҭ�%� �<V0��Q,�V+�8�>�/.t�X!\~����\P��1���� �+��J���\;3:+3�q]�ĞK�
1r[��_B�n�D���m��gN�� ��ۓ*U��uouSɨ�|�<����oܬ)[���<ē��ຳ`�(�vy�,�zh��Ý���C�"�l����pf�g~ҝ	[�o���U�C����G��vP�̢�*�̬�P�9�U��\mb�t�&\[�5��ѭ˵�);��gO�m�������m��d��d�m�2u��K��'vJl]� F��S��vN m��6�ޅ����]Y*D�f%�H8��#���<�Ӽ�h��L�.!,,�'�k5�K��wn� '́dA�XX�������lߤWO�4���2ζ샂c�R�7J�l�R6y6U��.���4�ڈ�>fV4���y}������]��ޤ~t���^��Z���3��Z�tp�K�C�k�=}bq��HU�h��]m���ٜmD���{9�s���$��X��v�)]kΠT��S�)m���G�9iܽ�[B���y�B�m����B����`h�{nnđE.O����ʂ�٦�vB�%(��M����ͽ��{�W����r��l���1K��[��Yՠv9��.q�VqWpǩt%�c@��c+�6�&��o[Ws��-��=�`	3uvnȬ�)�sE��8��zKȭ*�5�V�@�Rj�m�Y�����5��R��ލ�j�S�s9&Z�n��&��xg9J�u��O�;�Z:G8����I���&�Z65��U ��w}2�a�];��ٚo�w���o^%6����q�b�k�Wܽr�,��m�0�G5(�W���C2�n<ȉA�J�K�q�0��p�g+������f��o;1p��QSv��0����ɺ��- �!w,���צ�^��c�����������lwh�$ƗR/�n� �\[�v8x�p��²Y��e�h�kk�բ/;�2�ȱ��Q�y��=��6��kV��1�QXC;];Q%��m=ʒ���E���|�S����K]9�TD��pVrT����i���\��*��T5�.������_�ym��t=��_�{�)l��NYPX�E�XWm��0֣�+�lUm�)Q��]���.t�Œma�N�M�}b�:�p��ո����CDs��M���lcl:�9>�%A�L=��t'k�Ȩ�&���HySOUu�9k�"�F.������b�^1�֍�s�v�:��8/������˦��-�fSG�E����ne�F�\+�/��2tff�٬�{�+�8���lk��0uؾ�ð��Ag
�v�6�w�м��tw�|�y�{��o}i�{�_��
�G�P��.��g03��/*mG���XK=�:E\	����a�ąX���{f����Tcl&�vw�th����r���}`5�&qJ�W���Mǎ�uS�0�"f�\������ݺ���郧*Gn ��ܥ�v+���ӸF���n�"�HCϩ+��ݭs�[g�{��f�؊9O�*>�]�G�Y+�.�q�u����J�Nԇ..��C�]���&���{���jCjy��ɺ��-e�zj�wN�vkn����A�A��j��e��`�&�աh�!�����C2��ؼ���Tj�#DWL�r�V����,�����F!6��]���ڨ�n�5hs(���'	��Vr��b�mi�r�Ԇ��yR�Z��o��<�X�K���Ƙ�,N�k�ǧ��R��SH_2J�ݯ"2}m�:���m\��-5
� ʏ��č��W�����P�����Xk��I3X\�<,sz���h�P��vv�#���Zi��
�wN�p�ځvi�@���y$@A�2�vv���.�8EY�u�cB2��ns�uf�{\��g,�<1<�K���b-��yc�+�w��wB�A��8� +R�a��;��n�<,T�We��a�W}ԝ[�m7�Z��J�k���Jx��U��=��>�H��]s�	����ݙ}.���tL�֓ʕ}���Ik�)��"+mp�M�sW�go+��"��u�9�c�����.ǰ �]X�JY�s�I#B�w�7e�Z���b�8��˘��;v_;�{
�;�7�Ԯ���/�8�Q�qn���Y-��[*r�U�q.��p�jN� ���	�\�M���!�S0�!��U�-]����8�њ#���^U���A��[�;3���#LA�Dg%(�F�,6�0��hZJ�q�����s��J�-�6��ntU���otUƕ���_hY�����Vu'YƟ(t�:tÃ\���� =Ge��N����3A2�����U�E�Ś	y�|�����Q�ʇ�������T��:��Z������7��.��! ����	!I�����[�L�J��hVZټ�F�q[oY��,���y��jh�mD�����h-�x+&�5���C+,�F�8�
���:�I[�f��;aiB����x�Uc�W���J��XZ��{��4�:���j�����2�M��j���k8u�� �o5�]�H1=�%�1�u���<��8���X�	YwO-�����DIb�㌗�8���,�W'v+F�[$����{�
���0��w�U��աP04]���� }���1٫7v������� �U��TJƣ0���V
v%JB��j�)>{g$��A_w-��b<ot��ߧdmjӔhu���I���y�]iS��]��MK���r4'�n�cnu���!�L]�ua�	�f�׽�����]���YdH��[:��l/y�s��-mf��튳K6C	��t�/zŋqI���4;�b�����.����q��hʷ#1cc���Mv���j�l�)o>�<E܎V6�.�v�z�$�N�.�Ga�F��ݕ�輼�8;x�Ev夅Fp��L�W��G�YX���4�Ck.�+�:lRC[���뱎�ֺ��,dv_o�Lͩ
���jЌV.����"�Z���laZcJ�u�mۛ�֡ݝ2u�ī�V�q��D7��S)̫�F:c��M�WW|�
p����������νO�(��[98Qn�+������.ݖ�qںԢ�.��y\9nfe`�Pµ�^���u��l�F��=�<�d�h$g�*F��vn��zjYB��S�:�9���/7�|]�옗-��������X�u+�����P��M8j):�k�f�]�[V�7c#qH`z��[��y̾�����%&�e�O�lP�.��ݣ5�q��[艏�70��8�5"���Փ���*�+͛9�Wu��F�-�{�i�1� ��ڃ��Y\fM)��nG4	[���0c������0���w��b���v�!i,�Io�lT�AZ��zT7j��W3�P�����Kܽ|��Ԑ���b�
<7�buy��j�'��)ޓa��mh2I]]�d���fa�5gU�`4R���'72�:L�[w��:�w[�5��%>�&�^���X.��xH;-+4��־v��d���Zr��Ȯ�B}ܐ�W�+w͆M�Ť�g�kZ3�4�G[[�v�^g&ӄ^sӧ"�S�:�]+�uc���� �^��|n�����l��9�CM����o]�cК�I�����Í�nb�@�ds��,1��q�o8v���_s��0��Hp>�ۧ�3�$D��_a�8S��S�����DL2Z���V��8�1�yI7c�в�Vi�wV!����V�1[f��y�>�R]�]�V^�4���= �cM�V��	ΫKΓ�bY]t�f=U�0�g�8�>��f>ܳ���I}�}��ʾ�����/j�/)�(<�Oh1B��ę��9|T�i��Onr�=9d�
�1iȡ�/xn�����1�aκy�G����g�2Z�"�9��2���v�
n`��ъ�1S��Ħ̫����N:�d=��(WT�&��ݽ3� �wŨ�7��-۱����ؖT.f�{�&�}΂�Y:�ݳ�t�7��͜]�\��eU�˨H�|r�J!H�˲�vVv-��7��gt�� t؂�'�e�Vv�fQ��\���`j+�I"+Ei����cLY�D�x.�]^�ݫ�$6��v��r�w�ǂ;�Tx�V}���u�o�I}ʘ�~�`f�d��J�o94:B�i.B��:���-�Ӥ�ä�Ѭ躠�r��zv��L|{:HO:�Nkw���+m쪮2���~�\x��d��&ˠ��������/#$B�0ǹ�;/2XւT�3m��Fl����Ɛ�l�I.\�%ji��{���r�gaXyݺzn�7����IWL��)�1�T�ۭ-.v��;�Kމ�n1����
B�(�B=⻯��4�c]=̵���a����E��q4�tcrA�p�lE�����v9�S�XBy�剜Ѯ���=m���]v��յ3&�8�QkD�P�Mm�FTD���r�s�S�x�����AIB�ӄ����Q�qZ_\����"';�F�;pԐ��R�h�%��z⭹sGB �������B2�k�G]�̱�ˮY�A��>�7�ə�z��8�卩")kHK�S�5ή��!����>Ÿ��璌D�ѥ��Y4�������mR����bލ�F^5p�ƍc��H!�R��3z��Ye�Y�Tu�DV۽瘟n�Ş�K]u�ܻ�v�t��`�g�'roC�&ކ�r]f;`���-�l�uun�Z���0�b��:LvWe"Zӆ��e�}E��l�}����B"�{ԵP?^N&�c+z��`����!��g�(����g�G2��3ʝ���\�;lHF���k�2�dN�C΂��2�p��v�֋ER��Q�ֲ\#Z:m*m�)��[��Z�jl�G,ͽ�j�����/%�M������.N�♫Zt�9o�mZ��w�M���l+r��,f�=��[���xr��Ԋ�ꝟ+f���2u�n��S^ա�}q7oyn�2��nɿr�Z�w�i���E>�G8���Mlh�J�Sv��xu���NY�ƭu�eQ�+l�- W�e\�àF�^uis �αml/9B�,��d����7�#���An�>�u�NP%ll��`M�pW��:*&V�ƞ�Xu��"��e]=c��ؑ��e,k��6lc:Q��*ō���J�̸�rm�����p+�w*Ն6�����]�m.lp�3���U��{4��}Y��,�[X�П-�m�����%��\�u9[�'��t���Lc�Z���D^iu���O��-4`��
��f�9{!����5V���'b�)S����yܻ��8bΠr�%
i�=Q nVV�@Ңo; ��ԯj���n�X������E9��f*���ûeŲ��Yγl`#h��ڎ��t�d�)�]�s�Ya��<޽ҕ�˭;�b-=�@���#xu��&H;w5���.�8�.�C�`����-�,�(Z]b��\���W(�6�<;a㠍�YOEvh�\��D�WT�o����i]̰�gi���O~6$P����.�bA)2u������������yU��*�}�*�3t�w}��i���j�*�x�grd���
�X���[����ʂ�iM%��d�$���}�B�k��,M�*�%S�vNA,�:��0�]r�ws;�������M>Y��U��̽0MТ��t)N����Ȩ��F�+���|�&T؅��}����jڜ4�NP\�G��M��9R,�������ݒ���9؇O^
��\p
�x��1k^������\jRŴg]�X;r�Q:\�I)%�����䷙�J�o5�YwR�8M�͠S��s0�k/���d�\��o	A� ��V�Ët�{d���7|p��!��i�ZP�q�Cں��7�|�sӛk�!K�#�4�rivl��-�u.݌�0+�:��K �W$8)uݩZI,�4�����΍l����I
.X��MɅӪ,�p��;������3`R9`����ޓ�JB��쓀b��֛��)S�_ZW.t�ȗׯF����v��h[�uՎS'���kq��ЇI���	�|��n��b\�2��ѲQɆ�)k���t^�H���^Q�1Ԯ�:S�)U�I�RY����	xR*)xyfn� ��͚oL]�}5\�e]�'.��}l`�R4^��tU	a�..]=���o�iL��ӵ�2ty����v�V����1�wcs�X��
�R����c;L8a��J�v�`ʬ淨��%�ϙٔwzuB���$�����w>tH���(;*�\�����joh�&XȰ�����0�3���Z7��֧ik ])8mZ��PN��6���4�Yr�niD�N��+y9'Xf,�ޝb�w�V[��K&T��B����{O{i
v�ze^cu#�±j���VEF�b�f�$�
�����ŤK5���l5��F���v�w/2h�Q5�(�ϏM=*bw����850�^���K�x��C�;��ܤ4���Xޫ�	1�D�C}sn`�I��,��M�c+e˭4�"\�7��SYz[pܫ[UL�6�H{{���vS�!�ҟl
:��4J��k�XV2���v��v
sZU7R�9=�U:O��t�u��M�4��K'�t�Y,�7#���!H\�N]��D��um���0c���쬺�$�J�T\5ǻ���!����[� �UU�Lp�v浮�l��X�EB���c�v]��bh��-A��1��r��;��z��a����c�bo}V�d�+��Mu��K0`/Z��oΞ��)��!���qh�ˮm��V��]<Ó#u�0��R����T��|T[k���F��M�5���l����C�#u����xk��J�DܘA"N`=$m��p�{�(N�aU<U�K�d#"�ʆ�sit�W{��A�Am�̖��')<���o�c^E\�T���Es_J� �#����Wǫ�D�����ے��v2�:�v�捂���ivowP�B�把��[���tv�r*��i��0[S:�\��><^��f��r'*�x7,�"#s�Q/8l��:@�l��ee�&J���uˎ�x:iw�&�f&�ޒi0�j�v�v�t*��: ��:ϕe�94�N[P�:SV�p9.�u$�ū��5��JJ��d��e��`���]�0FiY�� �K�u]̲qF/��]�.��.�1p�G4�20N�:s�*�[�7X�k�S+0륳�F��T�kȍ1O;'G��F���PjtC�$׏6�Ja��K>zi:
��Ml9T))A���"Mޮ�L:s7B��o_UeqD�����h��6�2:�tஎT��D��0�a\�gZ�6���N2i�t��E˦��&�kH҅��x[����GG6�w)V���DGh�]�"��!��6��s�۵A�r�Y���Ch�g��(�謶��Z�}i��/���K��)��WH��9;�0�/�6,�:��PI�zH7�ؼ�[��VXz��Eڜ�L��yv�6���l���I��5s!��T��x���wa\����9�̵��RT=Xl�����9��ވ+l��N�k�jy
�2cؔz'(�JĽ��;>�ozՎdwm�X+,v�K��uހ���2<���H����x��R��v	���&�� ��7w��SYV��@i��c��źE
��㏸��;��a�oY�\P[V.�IU�̴N��֪���\%��G����C2��g�0�ȕ��,�v9�4�)�k�R�4�OTXj��6���xW<�nj�쪈]T�u�muv����;-J���fpT�,N���`�д��ҷ�ݹ�Z�؆���1�f�����-b���{MT��,�BU��m��{	b��T�^u��:���0��3��!�B��Al�N�Y�XT6r�/��	���gu�f�+�z�p9���]�pS䆁�r�%�w����ҝ2�\��m�6���'d�he�f�
*�;՘6�r1���`�"ҏǲq�L�˔��ͬ��3{a��IA��@dR���<�*�㬹y�'�u�4K�E�v����-�X��o�Ϻ�F���d* �\yhA9SE���e�#R�Ϫ�bB�&�E,�ސQ(E��z*�Cˢ��x��waFA�〝��^qe�

syۺ.�������!�0�Z���1���� �&�KK}����ʂ{�V�}�����"6�����h���D��]�}3���ݫF=���w;m�K�YYO��,.Ve�ٓdK�]�>U\��*�YiN{�	B�e����-�ۉ,�	��Mk�<��AU��}{��SZ�xn�f�Q���C(�*X�s�C���q�J�ݻzrU��z�lX����n�Pfh{���\u\�;r�L��ƪOd�MF�i�K�u1��n��f�g�F�����ӧ	���4�5��P��v�]]
�ͥ0��fY�
����j�rV,�pfȟJԳm�:�sus�r��O뼾!���&��<t=.�ȳ���P�{��e�G ����7�u����\8�d3��ߕ�4	?t�fe
�3�kj����R�b/��h�=,
�7K5Q�n�u��Y(�m�!�r�s!X����%sr�H >}J�ۡz,��u�%�`��j�����
�pM�����<ǐ��)jJ��Ul-�~fU����0X; ��aWZ�F�u3�9�Wڃu�*�g'@�����w³l&>5x�E��G�n�X��n;y�єi�@�za޵��AcU���e�B:��N�f*Ml*�Xj�ك��
�� �9��,wL�$�a���iRc�j+y�t�_��x㊗SI��k����pg�.);Z���*�G�qVͮ���5b����b�i z��Q�tˌ%�����!t�M��]��t�*�u�n�{�,�|�5����+��ԃ(�3n7:۲���7?�\ܫ?>����{��B�kPإ�o��q�57���b�+j���Ui�5{l�͛3tp�������\z�M^�'��ݛYĚ��g*P��L�}Ii3S+#G���{��\��9Y�-�E����j�������_<�Z=�t��Q���V��ۨ2��W��?�y��C�>�y�2vZ�+5�U��a�a�����@�����ՠ�;��[�3�q8~�0�
lT�D�����<L���~��{���,!�*�2����X�u�ʠQAϮ��aXoK3z^�l�t�u,n6�nm��]�T�땴�Y]�<�;to|�a.�]�o�ͩV2�i@S'+�+���ט.;�_u��aI6=3ǐ��or����1�e<!�*���A��)0WSvzg]�y֢�e^_$����H��7Zx�QQ�˽����̀f`$)�[H6����u�q�}9u�G�X�ntK"YoU��O_-�]s���[�΍���W
��K�jA0��¹_�:�ƺ�J]N�o	p,H	跱M�+�켳����3oGHl�N��o�]��0b=�]�W6֣����X^�l_�V�]9&K�������Q�x���Dk�O�s2a�ˏ{-���-5[�cWwu�껓�0��e�ֈZ���龑'���v��a�n��L��%�b��Z�.��X�FfWu��ȋ
��7����n$5_+�v*�ǵ�*��q(��u��ާ����Y2k��[^|��)�N;m���2�7ȶ��o�n��_m���ЩL���u��u�n�WFڬNA�5>#i[c���tK��d�Cb|j���o��������U�������.b�Y�ufY����4�˾�#��;�9RƝ_[Ȓ2��
n��0��6[�8ɏ��3����Y����"�\_!�0wh����s��8�tб�u=��"!;�=�Ts
+�R�T+YF%Դ�ն�Z��Z(�-
m�KE�l��1��R�(V��R�U[M6M2����iV�\Mh�kJ�Z*�GY�	Z�kV��B���[)Z�ъ�Z]5�&5R��-�b��X�i\�����TmE�-�F��[e[Tab�k-�j֫�-�U�h�Q+TTUm�6����Z%%iKj-jX�m�J���4�p�nR�q��kQ���#iUZ5*�-J�kT��ƶ(��R�Q0kU-.\Ȩ����jV�kJ����)��R�Y�������[[Fأm�KA[(�҃��kYmR�*6�(�jZ�V�E�q�B�F��U-��D0J&\n"�)U0��e[j���X[V��E"�Zŵ����V��������spDbd�-(�ڗ��xz6�r�ܮ���+���Ì��.{���lU�gz���ތS���:;��Bvs:���.ָ� L֫�����������ď�풶ֿ��IP	�`�r�`��k���E{��<��9����@��q��3AL�
���-��Vh��&�>�f}uD2(�&-ӁyS���p�k*���p��Ǐ��E���<�V(��,=�Ȏ�P�!Q8�;S�dʏ���p������NtX3��RX�N,��\y�tv(\q�(��"�ӕ=g`�)�;ow92�wI �8��F�hF�q�,HFo�i�G�L^լ	�e��3Ɗ���ن����L������9��u~�
�
R�`at��"����s�!�t3;�+5���>�����.����fڽ8&n��a�!(�Jv ��:f�{a߶I��U�{NP�=�qM9� ��:Z�0��ǋ�i��p�,��0|�x�zGc�Ӹ�Z6����\/����`
޸}ʠ���&��S�7��M����`a5�u��p!��H��Ꭳ;tMO6�ig�,���%������ݾ#n�ϔ�p�k��SpR	���^�Ǫ`GhL���ˢ�1Ԉe*���;�Y���K���7�G�i<��2uq�MX�;�`�t�N�[&�/Y��l�\�m�Qf�{S����m��N.ܓ�[��{�H��ҩ�J:��Q��K���],1Q.��~n}�%�*v�.�{�!R�Wϼ�G��c;g�*�8i�{�E�o���+�SV	շc�і�9�x�|��Tܣ^M/_�i��B��C��"ZY`�O,�K3���{?_~Kdy�/����vn�����Mb��	�mF`�'$��x�QV����@����{b��rܙ%��K�WF,Q�6��l�н��Q�XC~(׃��=�ʯA%�ʶKvD�-N[��3�RA����������`��}yꚯV��R�C7�W!���������9�]��5�����|�8��r�9S�0��t'Ra'<�L�	B�X����A�k���4Й�qb��T����׌KQ�2����B�(��p��o-j�U�0�>��T
�ǲ�RP�p�h����������W��/qh��;C�m��;�G�R"F�1��=�uC5���X�j�PG=N3��dܐo��U0�bs���㠏��\S�iy��$�( 9,{˸�_''6`������i[���f����z��=&�O3gد%�z(M(�H��.�hW���?���B��P��Sͱ��~��|'�tɘC��(�wS�*�jUݡ���8y��:5k|�Wl�.'�6��ES�N�1�2�M����7���w���3�����ۯ�PN��d#���Zv�M�}vE�I�&@�C�P��d�+�������FU�B8ύ�AU��l���.)Bu"�nks���
f
Q5C�.�}��=��2@!�Ƚ�����b�5�(o)q K]-�� ذ��!n�޺��B��!����רD7h�y��d"����(��N�,b�D]�-�E����X6�F�1G�C6s�a�Ȓ�zHW:*�+�� ��m��SSV�N�^F%�d���p(0:�j��o��_�Ta՝�hf����-����d��W��&;#�0C)�S5nx�n,��!�MD`�i��g�`����N�s����>�*N�s����%�K�q���a��l}���v�W//e%X�{f6��n%q���U�qQ�&��5��"�N_9U5��Y��iӎ0�F�cxN��Towr��p�
~����z=lS�$���t���sr2���Ε�3��^�ڽPʍ�}:�a�e;N�G3!U �k��K`Lި�?]����}�.%(�y=q%M���%�ŨP���s>{��]���PK`q>s�l�f3A����e�]3����ǭg{:�x�F&���-�Z���՚������*��t�7Y{�	G��!TĽ��Ϊ,� �\������A���<�=��n�������!�;�
T�~hM�L�*�mo؅X&i��V_��m�7��wgdڇ�%@�nAQI�XL�����T*L�C"���5�J5o)�*V,y����ʤ�'6l�N���A���rH��#{v��؂$��$h�pU�wq�}�z�sm�G���:�~g����Y&�qƝ5�rȊu�ds�2�Ŝs��E���ٞ�,�.@1}lL"�������Z�W��8`�+S�g�.�B�b�(���s
��j�UR]���%r��+�Z����<�B`Q�Bnx�u�������]�!�.Muk��;�W�g%<ւ����Kq�9U!���A[���<Wq�45�.:���y��6|,n�;���qu��.�W�q��t<�8lDw��d�/�-��Ui�:1�}����s�TVC�,�D����T�Q�<v*Bѓ�Z!�qj����u�k�	7�U��s^9�ǆ�+]�ȇ�d�U�p�{��m
�X��YA�]�P'��hrf��#��Y�Zߛ7�!o�V��3$��u���ۮr� �}�q��6��K�6r�5f�ͩS��s֢�A($����[ ���\�{�\\]��� ��n��Z
��6Qu{w�Xސ��%��iE\>�e�aE�8��"5f��S�n��n��IGp����)ߦ�\۬<�=r�MoU��#�6܅[x6S����M;҆٠%C\=B�W�mٔ�������j}�ϼO����ÿ]��y`�/�Lr��'��_��ޜ׵'l)ĥ��a����G(��`ޠ�7���DLLC[˘�F��v\k��4�_���{�o�}k�(�'P��#E!�B�[�@��M�i�Fm���@�O���S�C�j�9�آ���hq�r��	�vw瓭�K�{���0F^O�d��'l�xk����)�P\E�ܰ� ��ќ��O���~��O�SMH��s.MR�Xx6�`�E��<E7���b��P�����AN͘���A�aP�_&�y�`�Ⱦu�\+]��
�{���׌\v���ԯWŴ�/���,�z} �0D��h�A	k:�S���u{�2�m��š}�7�IҒ�%�u��׸�C�b���!��/J=w�0�`$�RbI�����h�s-��K}���6��D�o�}\�E8{5y�ɮ������Y�1���B���\/�^��zj�[�#\��'-��'u�j������r��8�dq~<p�7nň}���@)�Jj ���3^��{$�I��p���k^V��UZ.�y�ND4]Qe�4��<�Q`>Hl��)��q7�L,魊��\}�"!�_����:�t�:)N �r��QC�N{�au��g,ᦞT㴗r
/� �ba=�\���̑����J��g�b�r���Mu�@3�O�O��9��6	�����J.��C�gO�P7٭�=�u�Y�f�)-K_��Gl}+��d�%�h/yx�`حt٦�W�̘r����ԳS���+�+�Ȼ���̡u����]M����r���$������/��C�Z���Q�Ϫ�����%35vb�c�ښl0ΨM���ŉW��h��uF�G��������3���u��TU�hP�F�� ��w�3Ҧ�Ep15^~�dVF\dFс�w�CE>�7��g���ᩉ���[�H��D�W���k��8Fm:n,:t��s��rȒ@��su�f�8{v�޽��	n�d��ż4�쾮L`Nu��r��.<#X�u��u����ElD�i���Z�׊���S3�!���\�ͦ�Ԇfe�uv�I�gs�r�*�TzA�S�$Y[����M���]��䚌�-i�����*΋�.����Q��CY��$)�TG����T"���-An|�j32����\�^e[w��ޭ���	^}��:|Y����`%�ډh	�g�V��WL��s��A��}��<�֭1ȝ�$���(y��g<���+��D�c��0TIק[�&^X�W9�����o^S�݅
���~y����9[T �/b�Zs�ÒI
D���ܛ�v��b�N5��fw,��^m2,Ct�g���q�	ӡ,K�,I��$�4�[�9$,��]�jIf�fX�R�G�0:o"�7����.G�qJ��sX�c�$����)��vi� ���E���0ѰG�jơ�kyF��FÒ����=��������=�5�J����\��*"ֆT��ҞY�a{��BĒ�������ؕb��9�jަT�7%i,gP���B}���@��G��|.�g�yڮ�ڼBqX�ۤ���6��W{�L!�ޢ][�#VMy􈹑Ca��l�8c���R,�.UZ*�ԺѲf0�.M�ȷE����뱨��݂�Z��b|��_;��exu2Y��G	/:�0'�\��#b��	(r���\�pm�����r�]�ڀ�|�l��+`՛��z���f����<����X���$�t+#ޙk���m�-�;\h{�1K2�e�q�&��{!�Mz 3�rp��c����O���}u�%����GT�"ʗ:��"�*�����gswkBp�w��*��1�e��gbKQ���T8�����UMF��Zn��;'����9|L�'�ɥF�ϨT��D٭�~lSZ���n������P9�
����3,��b+{��#�.g���`�<l&���z� !tP)W?�^�*������/�δ[miA��<���f	�w�7����7৲��jNĨR�L�_4%�j�Ey6�/Z�f����zr�`�n��,w�'�
�[�TR}�y­"ޙ�~
�P�8�zŇn��'Fq�O�k�:z�gHb�{b�M�Ўr���c�C��W�{v��؂$���)�7�U�5�Sb��[�@�r����;�R(�����i�nYN��ޕ�t�v[���v����'h�*� �&	���TB,�����\��G!�8x�wƥ�" V�����*d�4�MU:<� �iK^��P�����ݍ���p�R%>RU��ٝb+��H�!%S����ǽ�;}Ortn&P��ܨD�2�a���ueU�-U�Ԙ��c��\׍�	WQV�:=[.e`|Cd��pΊ���d�{�=x릱sRα��:��O)MZQ;����Ⱥ���/�B{�!�5�^<g�ޥ׸1J`�a��6G?9��y��ȿ)�t��P:]Q��[���j�-��\(�G�sp����T�����uE8�I�$�iE
�q�2{��4O��.l���&��� ����V��,��$a�Gos�6�X*�2���h�S�g��!nT�݈�ɇ�Ⱳ�.�b3�#�7�����K%]8+�W/Vu�"����Y�	\`Ţ����Ǖ����)	g�e-P�n�S�M9)tr����E��d�r�zR����vͽz��.yP����xW*M�'��Z�v���~���Z�~m懺8��wÐpX�u>��������ד'�JY\Fx�|Q�J�A��h-ۉ(�^�^����� ��W��`�!,�К���u����Ҋ��"�Gy�ۢ��+o��g�b��,fMlcA��y�A�sO�W��:��CUe�b��O�&5���@b�gX�黹��]H���̹b��s^e5|�;��m��.8-��	�jU��*�O/��/��%B{z�v�at��L�C쮣	�;I�a;qDvtq��� (�u����_e,�,v�Fa�tǛP��=�8��3����F�b2�1S$q�099�[��9�k����<�V0�Y1qTh*�Jw��{���G�'@Ti�����}��,�P�a��N�t\U�!�)��JzӚ���Z��ƣ��[�C�|Pd����Zо���.<��2Ƙ�n��<}v��3�̡E�T��&6�N}+�*L�1�@׌Z�P
+3nbi袢����gKMݙWp�l�p��
t�h��l�@�|�ɒ*��6��{�9K�����Y�yC����D�34���f����x]Q~.�Y���)�.���{v
��S�mwD��y�Y�A����.y�r�#���I�	�nX-��e�'��PE,�V�����SQ"�<h��|�	]'��wo��5�v��^�%����B���{��q�#�O)�/�d�셶�'Q~�Y����x����c;��E�Ѹ��D�����w;&}��z�I��3c�� p��c2J�ϔ�U�qW�C����[0��5�ԗ�n-<%)�x�W�9������k�ٝ�9ؤY݉�YG���4�yҩh��ج�w��[p�o�թ�f;&0�5���n�;2��*ӫߢ3��	he��
��Wks:/4-!��Άf�#��@��IPJ��=Mr��x:���}5�׫u��Y��.&r���;7�s��я1882Y�}�Tq�s�����J�F��u|��<�יz$� ��c�B Q��ֲ:��m�(,�c�N�F�Ĕf�J�N溾�+�6҃�($+�J��!��@��C�_>��m��X���l"��8�d��vX2*�q��='o1��cj���3��8�Q�_s�G�{bqJ��#�s�@����+C,Sۺ�kX�B*�:�t�������b���x;���5���i]�j�*]Iq�{��g�����"�+�6��P7�.��A,�Q���Za/��զn8�`潁	P�����r�i���\p���k��2ٛ��.*�2��vû*�����NUt�;�����6��
�Z�n�N	�Dy�w[@N��<����4��|Pܑ��1es%��`��;]�粑��ٌ�	S�Y�,��,se��jڷ�R���]�]ܴœ�6�<������G!s�kL$�8G3��ŕFehr�PK{��,�K4	o�uٖ`����a bû�(�k9(9n�MFU��I-�0Q�h��B����W�Nݩ�s�4u.�I�m�Gm�ظ!�C��e�����[�W$w�=u� �Ac+�w5c)U໾���f���_�9��2G���\͵��
^9ӆ�_R<��R��9�BZݑ}��v�$�F*����|��3���L�.s�z�+l���]ˏ3��B�r�s��5HzAJ�������m��p��N���R|^^��������.�bPL�Ye�u}N�'��ώP&֖��9����2-yMN���{�2���/�hV�����;[�)���ѷ�B�i��=pb}�)p7ڪCW��=#p�<ѵ(��$m�<���J�[��s���M=���6��d����lƸ,�n� ��7ՌH��c͍�H�bezk�-��<
�]0LP�=�V����VPy{��IK`ڦ6���� 2mȀ� �o6w1��]՚:�nV7��C+��</�cջ�HC&���C]\��zp��k�3��d7����)�m�1HOօ�M*�;V��#���� b��|��~�7��jʒLv9��+�Z��*�w�᩺��E�G�f�䪴���L��c���:���9�[���S
v�[�� N�����=B�X�
ż$ݭSmQ��U�ή�r��F�����Z�s�2ܠ�'&3ƚbaC��<w!�y�!M���>��ޢW)u��us����8��CU���
�b5�~�ŵ����o;�;U��̦e����
�z<XA����@�H%��>�q��*�6�ڵb�-���"VW��ժQkU�����R墘�b��TU*�֭([)J�e�����F6�R�������ˊ�73-�%ʊ�h��6�hYFTCR�ˍ�l�A���C"�)U����Kj!Q�KQ-�R���Z�օ��+lDJ֊�\�G+i�&�U��V�
�)DZ"֪�D�X�1�(�����؅m�Z��m���c�K�Q�TZ���F"*V�-���)V�J1�5F6��`��cUk����¥QQ-�[J�����VV�ƊX�Km��2��Rնִj��kEV2��-��X0Z"�J��k(ڴdKj#��V���Qs+����iF�T�cQ��1�\�Q��*5[j�Ҷ�m(�QVQ�
1s(am�VՈ��m�1�������U��-)e��e�Ym��<[���~��I�A�N8Wa��黻�6>��̥�%�W&]*Z�4%r���̓�4!t���wn�F��.��2�i�)��@��]9�Q�t����O��Ź��r��t��F�i,�U��;�oU�fգw'��9U�.�&{����a9��S�9Kj�7�s�R8ً���u��O���$^s�;yYy*)��5�d0g��;���J�!�Q����nVEd`�ȍ�)���J��s3N�6l?LwC69$u{"|��+�N�	�qaӤD,�\靬�U"�3�wG�,�7,�GI*�*܁!^�^���ъu}%����fC(��Dk��;Ӯ:��F���_�/_G!�"� F�k�c��G��y���Y�ƶv�R����ʲ�l��$��8��}������)#A��|\�E��!�eGK���`ާ˛ٙ��S��^߯���	�;mP�E�R��&9$�� �*u.�1��X�v�z���b��ء��p�%�p�l';�i۱6%���IQX$̗����0n<�H2�uŌ�A��=����r8�K�Q�'t1��p�)���quz�EޛO����=MS�x�.�8M�ip�f_,^�맀��P�ic*M��W�����j[���H��慗v	�=.�}Ａ��U]�콍����$T9rʭ��S5��,�0��î���cr�㽄uH3�>�U/�:����۲�>T�l_�r���L�ѰBܚ�@E�w\���MrT� ?x{f�a���^�NhB��O5]Y���htV�_'��.+6C��!��m��S�`k3���ovr��=�Ct�Q{�[�ٯNX7�ӑF(�ٖp�g.0xW���n�^��nO��^n{��E�9f����.�μ�Jjɯ�"�C���AA��mXR�?��i����S����)��Ե|Ǌ;^4&@�)`�c�k��"Csf
��d����w�Mf��������DN���q� D��:��T���"�*�����KLi�W��"g��P{����2ٔC��5�u�X(��C�=��UT�`-ŞL�R�����
j�7��~���:XKP{~�"�:'�l��:��hr��Ƞ����9��ʛ�����:���E�=����r	Dj�P��r�L@gS>+;E�ƽքt7�\�Pbn��W����7~r���m�G$ؕ
Ti�(��/�Tʊy{���&N���ȥ��9�����1�}��ةM������������w�dR�N�&1�aU��>�gQ�E!^�l���m��^�'˦�ޕ��ܓ��4'���@F#�xN�y�7�^uJ������9�3��Ɗ�'q�[���������Æj��4�Q�#���=�K�B܂���u��p�H�=�X;9���-ki�|��}���e�LW�WMT饞2��>%��w���FrH�}B(7�j0'1�WV��^�|�w���"I�b$93`я7�c����;�aJ�QȌp�瓡���"䞏J��U66���\Fn��^��%�����-(|n'X��,9~��5����7���UKTt�D!������O��4�Q;�����ݩ�_ڄ���:��&��q�mw�*�����X]A�6[���Su��aB-��ѯ	�y�,j�'���Q��8��PVu�E��q�r�4��������-��XX�k|����_�{�O���������Yk)Z��]���C��(!5DןuNE��x�;�j&؍:�wfVRјʯL9ydӌѳ������Z�3of�U�|*��E�Mr�#۫ގW���X��1x>UU�#g��e� V;�UC�U��.KӍ�-�����V�*E>���:;c�L�Wy�ڬ#:u$��<hd:bH�:�;��[��O9J�/�g�'kWL���-�l���wz%�Y]OgKL!қOM�MĈ�@�ˣ�m��5�C��F���5b'�'��n"�q�wm����}�*�Rz�<�zp��oT�r|rBW�qiYC|Hʳ�M^�N5��އ%�-ѫ��N�{Vy���~|���ʣ�V�,�#���xѡJ�ݾ�2�96��ğw)��"A�,��n��(��d[	��cs��\��":QF�%�K�#�+�)���RN�sr��X�t͹���<O��i�n,:�:���,u3��r"h�}���"E?8vbg�iM��%V'l�.̏qa4�<
$a�T��P�Nx��&ݛJ%�ÓIK��3��H�#����P*�8��ΝC]�V.����W������F� ��s���=9H�[��p��$��?,�4/�~ s�r{o�F/;�unx���0�=�j��-�fL�GBs�qA�I�r'��@�0t�N*&;nt�s�x�m��Y�9�ʹ����QgN݋�-�.	
���)��vAs�n��Vp�ԼFj�SMw���N���>�˺����ʃ4��9��u�y��q�g�`(�%1������gQ���|�F��)�����9��K��W*_'U�V'���r���0��
6�zr�ז�z?q���*�����conq�ܝ��̴71ӐЭ`�6nF�S'	��轼��{�;f�	|����TT]X��E}f�ۋe��g9y�����7�B��V*Q�C.[��s�"�u	5�S�6r��6��X�00�(�Z6h�r�N5�Ѕ+5��F���F|&;r}r��e�������QA��LW��	"Ս��
��}YS�꩸�9��N�@ ��X-M^893��Z7��ga�63�n�;a��xW+�^הכX	�Yrf�\B�c�s g�Hf�
�.���#!��:��F���]˦&�\P��}T�07?����k��w��7u�F�ig�5`����^�4������P�efc��X�{�הܠ�Q��k�ڲ��ڑc�dP���}G�³�.}���W����RE�]�j��P�C���mJ�!ȟ��Mߪܬ��*�BgB�J�9hH�\%����+���x菐�޹�҃�G��鸷N�Έ�)�W��0Ԑ��9�E!�GI+ኽ����%�6*KUI��>xĵ�n�m�8���<!�r��Y����*҈�dqG� `�ht�pL�<���TĪQ̹����,Ai��8��w���l	�� 錺��)�h����W�RQ�+e�o��r�5�!¶^�ɽ�X���LO�,cx���[�J%���\�{
�v��:T�sf�d��$,�]�d�ݮ^�[���\�vl3M���[�
˳�e7���c��G@7�l��;��Z"F�1����tQh����7晏�u���7[~��ѡ��a�S�;����mH�D�I�؇a�$�@ӓG�L���{��s2�p �S��щ���%�p���nG�݉��D#D�Q���gY7���{�D�3D�����=�`䌷=��>��3~�6�ӷctԼ�ܗ7��9�ք1�Q˶��BM3+�t�̛-ɬ���꒻�G8�^	���-�ǽۮ#�'@b��N'�-�Z(W:!�� ���+��ٓ¸V+53�Bd�G)����VY���28�D�,�j�Hק,�N)��b��2��Ĵ�_]{re/^��2���H�U[���;�/�]�à�1!5d�}"/2��X��ᾂ�w��7�eh��/ޞ�s�E.���7J��ߊ(א�<Ņ����f��g�͘*��q�x�3�jƛls�^�#��T��҇���6����4�x�s�0>�"�*�W$�����jƊp�=�v��Dr�7{���A_t��B�zŞ�^<���mX�ʛ��kӵjG��@���($�8��<7�m�
�2{�ـٝz/]j_7�q�t���g�*����/�s�V'0g_�9So!r�����ЌQ�����9������6M՚���y��/��L�"���e�I�����yI�R��'�μ�|x��;GH���%��S�b���P��:��8�Y�������cO����2.�D�i�+㥨�7�G�\�Dx���"v��Q/��!]�T��q�kzڤ�"��q��GQ41�<]�A�U��uǂ�z��
A2||ЏQ�ݖ����>[���-{�V�5��X���G�d�}`�bzL�<��Ⱖ����/
�:���i��Ө�%���F�H��\�-*�L�f�s��tf�$H��bl����=6k�؂��j$G�"}�"t� �Pk�=Ϧϑ��ZuM�E�F�ө��Q��nNO>BV�Rķ;C�"6Ȇ6��@��T�d���; J	�D"�-���/��U����'q�z)*��tk �Ô��>�m����LX"���@�׋�v�!hBx_nNu�i�fe��O.������yCM�x]av�4�PdZ��S�%'b�-^���'�b�J��O�o=a���F�J7�]ژݗڀֲ�-:Y�\�VV��<;Z��'<��@��k�T�Rtz'��əN�����b5 ����7|-lfi��޽y��}��=�b��=�iY���~�}{Ϝdv]�3�]"��AX]�uQN �r�4QXY���Ή�;�y�lq�ۍ��"#K��N��orFΜ!_s���-�
���4���3pv��}�x4SE���b~��ާ�}�'g+�
VF�vt��{w�^�/�k�-�ڊ�;[zmP�v����p�v����>&����n���Y�@r��Eн�� ��a�A�@��ӆ�?
ޯuf^{���G�r��s<rB5�@U꺭�<���L;f^��`�U+�������UMF	u^Չ����ӯv�� �b6��"�Di</�sͳkvO,����Ky���\{ 2L�y�8�*�#~S����߭�Z�a�|&u���<�s�a<��y_r2��9�#��V6���%���m:���h��G��Q�.j������҂\64�hh�w(Q��b����.ݏ#�M+j�Mۗ��oyg��p�7�2#���A!Q8�xF�q�/����1����~�X���a
��Im�'���������˕��mu�i �{�<f����v��d9"5Mٵ�s�.`��h�0exZ�2�^�j��{eL(�r��޷�q�.�Vf�*B˚ycS1ʲ��L��ɉ���\7u��W��b�;j��y7ٚx&Nѣ��x��C!ṍ�R���LI�R��L�hN�dtB���L���WQF������]�ٻ�;��ܓ�-�fM�mB6s�qN)`� �εU��1't�־jfgrŌ�3l2:��z�B9��5��ܛ��l��B�>)Mz �qo�'lĠ�lf����^eu�4�WB��H�>��A��A��r�!�"�p.�Y���yNQ.��֞�
���b1ta��פF�QS��Jqi�DF�Q�*y/#��}�f&���;�ى[����M��U9��6g�r}~�/"�%�7��m˨��ϔ�P��v�tk٫[��7F�ւ��qB,	��P%����C���X-,�ll#�2E\"�k���5���*5Wf+�~�tH�y^SA5��iF]���@t��n��ſ1-���y�D˓I�\�)��P���F�꯶1����{�>�x�=i�mF`�qt�:C�>��Ȭ��T�}��G%e��!���YApSA ��uF �P�[XY��7�F�+v�����-H�����M�*�ؙ�՝>��3#/_����q�[�Q�q�Ɋ�{-ޚm3A���L���Wbm�ww!j�9;xL5�N5&�<�Ro�A��e;�嚺��{zv��fl\nr�WǂD��B�޵��<��B��g2�*�ѵ�V�]�x �Z�nf�ܞÁB=�ʎ�.��_ڠ,Ƃ������Y������`����'P�����>a����:��Pg/⫔˯Zf�$>�_z�10�)9f��pY��"v�p�'d�ap�}�^�������g�!\K�e5$�cU���>|պw�OZ��.��9�FU��n4��H�
iG�#��U�.�|�N�Cb��dZ/�y�����F��4b'�ސ�n��佑�	�y�a�S���+R���T8	�	���Vȩ�Ijzzz�3��Ik�۱~�j��\ws�r)�,�)E�gb�$�]x���-%���oV^7�n���:����X�q�Js8D�<�S�g�R�!�O)yB�1�u�A��5ĘPƈ'��@odo���E؂�ܝ��#�f�!ͨR��W�x�f��rɝ�	��p1�
k�f
V��d�rk "�;�J�#�IxmT�V]�ڴ�%+���{�Dc= O��v��0Yn�!i��Mv:A��7(�]U(���W�00��a�aFk��2j�15bB=�����(���}���k������3�0�W��:���������Ft�f��XD�
9��{H�V�*�!A��H5ϩ�וu����m��	RBu�m!�pRY��[%���~xe���0>ַ'|����W-��i��A6�'����
f^�.(�Xܹ��j���Va]�4|��E�v'2R���Gb����Hgv .�2���S�]��fR�՛Ti[I7Wy�t�Dv��j-N�#D�+�K;"!=�ˍ��7>meaٝ>A5��Ϻ�uFe�eSa��2W��iҲtk���6�˂	�<ɣ��ɶ�yIb���J*=]K�:���v�N��F.��J7]2����z���̝�����]��iOF�+���&�v�Y�+�D'��8_�Vv.�o��[A��Z��*�)�
,��QTiZ�g(��̉v�����?h
;�#��y�浚N�,u�]֜s�ᆢU}�r�
�G�a��Ҙԫ��TÅq�y��Ln���%�/�p/�n�h�[n�+%�[Ga+�*��6oM*,�iF��+.՜�o*�7���lY���D(Zx�ya4� ��oy�0oM�Yk�
6a���gt���c�x[{$y�p�
c�4�_.&w<ݮ�DqEb핕h4OY6��>5�)U&f^�ay�Q1,�Z���$-i�x�}��^8��k�Y���������d0��! �� �,�t�W�ݦ��ճ�jt�0˿��Q�\}�����⋛c#@��M�XF��J��0���px�9��udQ�;hB���2�ڍ]�ǣ9Ǒ���Z�yٮ�p3��)�,]{;E�f��-̝0��*�w���@��Χ��/�����'F��e*�}t�u����7�s5��趐��J�������V�q�X�%�z&]�Fsx�-r����ܲ;�fP|ey �9Йí��,Sd�gX�_���B�2E�$��3�&,ǇE� A��0J�T�cky�K�(�s�+��h {���1Xo���7�u)��aN��X�\���:L�uj�;Y�$y?�<	&���ΰw2Lc((�NeP���h��*�.�*U42*�=ӰnB�V��������仄���v�]�Ⳝ�ju6m��N�X���W���(ڒ�z��H�a���An;��Ej�J`�� *^+x�w'���N�n�C#G&A�Uԓ����A�f�*]��Vax*�DuKZ��l�c+E@�^�}�[��,Zw	���밺�8�f"b��-h����M���!}eB��bF�:e���o+��8��՛�fG|{��3����:���P��(޹RMoQE�p�����`�^v|�˱1 ��3r�[��-��\D�Ƭ������h�� �"�c
[A�DUF4��h��KOl3��T�e`�QQkb-,����QPVQ�)jԢ�[� ��Dh�،Ecj�mTTJ¥������EVR�b�mT��*-�Tmcj"%��(,Rҕ�m�E�5�X�-�iV���#R���(�Um,�j",b(���"�j.["�U*fTb�4����DQ-�1��h�[h����cUPU%kA1%�+X��E�c)
*��PFZQE`�
6��T�E�f4Kj֭e�J��j�����%F�TTQUEc��*�,UE[j�J�&R��VV�2҂��ڥ"�(�fH,YmX�"�֢"���(���R�)j�J�E�kdQ-�ƥ��#l�j�jµE�*�(�ED�`�m[e�
1EXQ�c`�9aQL���)Z�T��ۖTb�1���m�ET��Q1���"��PZ��V���Eq(�*�T���ʕ������Re(��J�
��EQ-��DQb�`�JX�|�}c�,��}ŋ��o�a���K�%���2fǺ���i�YѷW���>j7x�L���rC��;�Y�t�����J�k�����GٽWQjq��Z��zr���S=`Ř��â�;�=Vsq]�Kv����u�E1�A�X.�G_s�"���.�:��	�����oܼSj������>�S+&��A�Y��-���:��_����=�C"�ڦj��2�0yvژ܌�����)�g��Hn]ѹD�N�'�P�]�@*�v	��\�4~��<�h�ʥ�ٝ��Sk�lڌ͸|�rpyj[ghM�^"%��T^K�T&}��z9غQ�Y�0��G�����Qg�����\靋"��$+�R�[>~lS��l�o��b�{;a���������E]3��	))�.��_-FP����z� ����:S+�}Α�F����7�Ǌv�P�`fU7�:&�)'���ۅ^g��c;�P�)j��?�ңU=鬟B�	f�̭҂��;�4��j����5���QA4�<�ZE��1ܓ���b�ͻ�M�3�nLD\G�"H��P���8-*�~���9���4��Na��J>O.���Kb�f�,ݤ�c
��l���	74��Fp9�Ni�<)��+9���Uw9��T�6��ϱa4�AO�<T`JUs,^zn�����L(`����2tct+m��^��#5j�嗎�//���[SL�kDWi͉+QY1sY��߇�� 
V��(cz�΋��\�����'>*DA������pJɐ��.��Ӷ��ޙ@�%R��5��Yf>�W��Ȇ��.���9�vL%��8��է��j�l
��3;׫kԜ�\0x����[���C�<jr����
�:|5*��̾��-���)$�L��:�m����>�E�q��.��sF��uC§ܔ�R��{���S#n��s�^zy����n3fT�F��F�ʐ����aw]�_�)��nY&�QXY�9ל�'� �$���Lp�}�6�Sf�i�Of��W�)��I�ts��,!�D�O1էFL��fg)(vLuOA~�iF}!h��R�0�N8�(�z����!�X�Q�L�=@���P�f�ꧤ��Q� ���Y��������dAY����~�Eׯn���5h�8ny4��1#K�l��sϦ��z���7bN_H'$x�k�<�����Z'��0��/�W�K�|��}��f	~��P����z]W�`M�ߟ=�;�o,��W%�W��!�:3�^f���b��^���Tm�@�v7��w�׌�j}�ۚ�Q/ϲh�D��T���d0��M�W��X��ѕ�4ud�9�T���]�;#5��3v��U�>]��:��|����4*]��,c������T��opyڌ�Q���XU���������4$�U��$�8�;A�D2L�Z�'��7�=L�M����<g.��t�u�*�v<��n�%s�t%�xR����W�����3�Ӱ�9�!��{ �jm�j��,�te�vo,т�U��T"H�(��(�1�p��1C�̎�Ԫ�K5��I��]���Ω��P<K<88�xO�]�4��G�:�xؗ��L�!��t�.P�ʲ'4��T\U�,������v�YKT���_/gp5���ԣЋũTH�)�繛�e�g���7tNյlɰ&6����R����dF��=B���q��hd.�kDǎƐ�ҝ��s��g�Ԙ{T��HR��)�u�WeE�s�*�a
�+{��px�$q�٦��!�P��< ��9�E��Q��{"nZ`�m��F�ɺ�j���k��@��q�ڞY�E��Q��G�9`��m�♙�I�=�V��j5`:�;fUjU��`�|�e����32Q����n��u.�4a��q���!=J���۫n��K~������v�t��4��n�'I��η᛻:?�m��d�c���+�f�|����fa{��w�Z��g7g;]
Ɛo
�j'�3��<�l`b��NK�7�g.���*��{xj��fm}�{�� %��w�#�Ƕc��@�mEk�rP	ѐ dY�q�*C7��W1�'�'(6��^���Ue�=X�w��D����4X	��eѫ�� p��c2J����۬�%!�LS(0"��<Y����e�po�%}�������_�<�Q�#W�,�@��)��k�
�+��=�2����텝SA�S��F����x%��<M3~��R���]��o]�-�9�]x�.���t��5@i��V���d���(�n����#�.m�)��̦=���u������Xz|י�)I#�"|���X'�NY���y��bw�Ѩ�px_f��U�X΋NY�a�$���g�!\K�c�t���g�I0X���w7۳�&�0�Y_f������.lR�ç����T]�М��X��:�b\��5���۾f�ۢ1Բ�k��E�Q}Q���:<�rS�IJ�{��Gg7�G�Ӝ���ZQ�P�c(W��n��ϝA��\ws�r��A�^�(����om����o��uӴe�ֺoD74�E���;�@ۺ�C�T�P�����ZL>�W1n���V�۰O��EJr��p� �) �����Q��^��lȰ8K�t@�K5ɗ�X'�u�e�ԍo�1tԆ�E�>㎮b.�nʻX*q�SIa��xxx �>e���$�_z p�@Ʒ=�$���'\E�Ct�c���'=�`c�beJ�)v��jT�e�(7-<�=�,$��L�h���L#�/�!tQ͈*�'h�.GΔԫݱ��Os�(��m����{բ�S0R�$ǶfO���.��䧗Y���H���޻�&�h������	k��ߛ��1V[��B�p!l�X��&�eŞŷ1y5;l&e��|��ߚUu��'��2h5B�kӖ	�b��l�~������h����׳����Қ�H�rUh�u��;\����+�s�"��D��AbSVM>�2(l3�ZVFP�g7���;�F�9F�-֝�E���兂:a�Z�`�m�S5~x�c7�w;�::���kd]S��Pkj�.�;Zl
��N�8��f��Y�4�Ny���;kl)��{s_k	�J��Eb��n�6�����]p/
�|�N���/��h��9�9����i[�[�U�Jr�=���:[�*�|����;�8\B# wS�(���3����^�:E���2�f�����>��ʵ���UX-��/g���}P�#N��UΧ9d�%L*N�jg��w��s�ܛ��͖�������!	�YtvQ��Z�BNe�x4ɉ̉���T������xn{�����l}1M{�����ow��3��I�fQ�%8܄)�-ʮ9�CQ��]ːO���b'h,�M=v�w�Ԫt��7�����Uq$�)'���7aʿ3j{/�(G�Ur�ϏC�1='�2Р�Wj�uęp�u��"�YN0k��e�c�TW�J��
��ݸ��6yoSQˮ7�M�6j��e$EE G��U3��-*�L�f�Ý{��'ܪĲ������`�P����`}1�0I��Uă"8
��������ˆ���ihp���)����l�|�R�g��u�jz&\2A	����PM�Y�!n�*�������k*��\�s��P�y\�遇('vϬsn�*5ED%fA1��L��/�U��ֹ��;�4ڮ� '��^M�x�.�уe���Цm���	Kj���\���**�S�AGe��.S�5u!����f�����,�q��I�4��ߜI����8�l��cs�WY��`בtvl��Zw*[�7��k�ӄ+��wu�TX,�D��E�U|�%K�	���0�r��ނB��0#�L��ܡ��m:����Ҁ�ʿ�L�2�7��J�
2n���1�9��Wn��z�x���\Bk�������F�L����)���8��]:�]�s���tr�c�jHr��7q_| ���i�=LÞʍ�~�u9�y�3!m��z@�/#����/^���G��w�8:m��Y����u�W�z }(YQh���<��H�^53��K:��8Zr�-��Q�z`�4C��&dY|�>s���������v$厐NO�HF�yM��9�iN1��8�#�-���^MN��&Ծ�yURqgع7��o�ޜ���b���4�7��y�^q��Ma�s�D_��Z�_Y�!sy�8�UA�F�M�}/�x�e�*ǔw~�p�`��<�&�=�Y3N,g@�>g��a��S�9����;P�bk��q����Y�P��^/S3.��n���`�%V ��t\3�C�/t����'p���g7�x��0'RԚ�I	q2>�n�R���=��ֶcsQX����u���UQ�˄^�Uǳ]�!����=9QЉ.$p�I�R�8`Mp�r�e����NeT�,Nm",C���+!�n'D�[V̘;0��9�8u�(w:*�FR�4���J��wsDUۤXIQ!e�����w����3N�-�cm�u�|�J;<��߱���Di����<�T��9�.�ޛ���ǅv݃lK��0���f���6�
r�9��=�LS��y��XcȻ�|2���*mst��U,u���#�b�S�	ͭ�u˦Յ��{���=8�\ӛ�̥Z��Ď��C��
����gN�@�[��Ց/B�u�G/o�Wk��b �'#WR��d��}ٿ�dxY�Ϲ�lY�Ld�����!��uow��!��^�F$P<JÜ�V����q�ݕ)/��u���2bO�RW��3��b"�ݰ��AH��S���N��n�@�}�O̯��r�q�q}N!�>9�O��Y���s4�0�$�I��I��t	�3#������q�����_̊T:{��1�ԗ��|��=>��'���옟$�Ă�*~��'�TJ�������8�N�z�<}�4�į�~��|N�}��O˟�Ue�������_=�#'�I�w��i�dm���bi �����^$���Z�9@�
T*|ş�8��жi�%H:oԘ���1�d��Lz�s�l|pʼU�}�:1�xY a}g���ݞ2b䯇{�Y<������u%d������q&�w��Aed����i�����ԚI���8��f>�*>Mۈz���?o�0�A�b����3�W>���>���0�1�m��c1���I����?h�6�@�Vx}�0����Ɍ=;ܟ��%y��zϰ�&Ш)]�I�m"�g;��7�&ٌ���CH�&c��3�r��o�uf�����:�����8�!��A���g�Y1���|����UH/��o��<H/���m����Z1�����&{�����xs��'��|@�=�-�߅mF�Ϸ+w��TeMt1��&� ���1ԩ����2��i�_Y�>M?0*Ny�>�m1��� �FN�&&��c8���2q�1 ��o�$��1!���� �Hd#*{���x��g�5��X��<LH,��=���������3Ԙ퇨f�
��I����(J��C5g�L@��L�&�����vCIY*�3g���
E:��QY�<	��}۟NR���,��_��8fo䏟l{ݡ\{��][E�ܺT�H3E-t�{{:}��YD�)K��^܊�0uåb7zc��z\�-4�u��o����Z��fȚ���ݖF�q���,�/7��H޷X��ݵ[�;scw6��{��X���u���O7M0�»�~�6���bw}�6�PY�s9�P���:�b�0����c�C��~CI���i��T��Y0�u���&��+�X>�~���Oپ������:�1�~H� A �>ݑF:=�F�R/����l�f3����u;�N�56�Ru��g5����Ԭ<k�%a��0����1 ��)y�O��Ax�w�w�y�;��y��>��k����Jú�I�O�Y����<@�T����4m����V~����H)�hbJ�2t3�k�%@�Wú�R~O�*��*2bcĞe�
Dd��5��f��o���s���:�u{ĂͲ6����m ���C�I9���ݘ�PS�]����N���L�8��Rz���s!��:��|����������jm"��Y��ړ7g1&�����O�泾�������b��}�d�H� �d���2��OɅ�׎�*�c����L>C�.���8�&&�y�Rm��P_�f��Ld��ɦz�b�0����膟�~C����}Ꝍ�\�P�_vLo��#��>R���<J�@���aS2c��LB��9f�I��
��-��Oɤ��%�d�1<=�& q>��~f8��8�>�|I�+��~ך�����Xv>@�Y�'�}�Azz@i�0�c��N������F��:�$N�^�Y�RVo�M2c+9�<�4�R�g�cĬ���B�-��2z���@�T�s���oʭ���~��UUm��&Ϩ��@��/�N&:`T�hu?2bc�r�	����}��H,�'{�Ԟ�LH.<��O_wt1��,1���J��m1 �k'���IY�߹��{]���_�%6��z�q����'$#��3�6w�=eH�q+�9�7�d�<��%gY3.�s�i'P�Y?N�z\`T�k�h��� ����}d橦'��|`T�O�ϝ��}ޭ�<�3��{�˯�]�4�����q�P�1�wa��
ŝa��0�Ax��1�����H/���:���T�O9���V:�'uT%B��~9�n�*���s�&�H,��{�UP�G���X�㓥Z�P�AA9�7����<��WP���@�y.�����٦E�cc*�an��F�mxϲ��־�� ;h\ɽZL�<;2M��H��%�'%�����3^!�}�N��}�l�����c�ґ6�nV�uo�x{��kJ�������@DL{�G�n��J���R���0+ڼg���$�ݚAa�X,�.��Ϙu1��{���<H/�>ɤ�:���9�=H�����N��6�d�+7�W9��6�^�|����_��]U�����4���-'Y�ۤ���O];�1"�ԩ�n�z鞲VM��M>�u1�N$��_���R#y�_��Ag�Vf��}LH8L#}KwF�p~g� 
4G��	3���&��*
o��A��'S=�`��~a���+��Y�1��z�$��=�4��"��f���%ݟ�1<7I��:ə~g䘓�T�=�j���Nv7�%��]��l� =��5�ԝ~t�S��d��OyM0{̆>0*O����<C���}��i��P���l�<B�g��i�i �a�yi�i��Ă�ἇP�m*En�m͡S�Z-��b�&TM�|#��0���t��6��T+��6����Sg��I��:�A�}�4�Խ�w\ɶ|�P=O��.����S���?;I�+����}/�T�>g�9��?}��9�W�k.+v>�Y�� �'wa��>N!�<����T�߼�hJ��W�y��&�*T7�0�jVO�'y�$�Y8w\׈)�O'5����2V�̜"z�������jm�q9���~��B�ɉ��6��)���?'�v�'_�4��I�P�v�\`Vo���>I�Ğ�2�b)<{�si��Lw9�jC�<	��]�dV�.,���X�|��A]�t�xʑd���SL���$����3/�P4��*Vj��~`T,S�8��A��M2i����L��a�0+��q1����v�@'�A�D�ٯ��o�>�螗�P��ޞ���
ŝ<��C�� �a�{���xΡ��q����R/ݲ)�+
�x��M ~J�f���$�ݸ��~���(�P8���b���q���Ш}�������ʋvo��^�=e}`^�p���?!_���4��ְ�wZ�J�Y�7�����Ă�s�jE6���b�ƤYP{MZ�R�~M�9�& T��(�+'mBy����v��w�
L�u��gnn���wE��ό�-W�x뭲�������C�m�-��3~�*��UF^=�M]��[|6����L���*�a�D�x�"�wܔi�
�]smh�Co�Tm)�*��V3�t
K;��6�]�ٯ�c݌����U�M�]�)�q�L��:�/L��w�Ն�Λս���ucE�I�3V|\��r4Ne�XW�l�!W�U�4��C�卾,�!��5�<������֋2�f�f�yP�$˶KR�.�@�eD��I��֗�t��n��x,K7�������n�V���톎6��_eƪ,���p�&���V�F=��'ZV�\�X��6�!��Rv�IU�\�FlM ���[�:��L�n��%�F��Ն;��v�"�Wm��ւ��������qZ�N>}�J�Zom�y��e��A�l�'��rC��نG����ݹ76S�N�Xz����Q��3MI��z����:�T�O�q�P჋(��j�Ohn��<��^�w7Q�G�
�
[,=�&��L0�1u��8���l>�)��|ګ�����7��}pNh��O�e����4ދ�qp�"�
��եj̇[�5�Ds{�[;�˟!F�r�I��Smg����b�g;�!o9�W��T�T�Y����;�DL[�u���ѵ��ؒ0�vv.�R:�7����%]��$���m0��Ie����M�7uɴ޻6�s�>8R���#��Tҳ�8x�ͮT��ӛ����T"2�A��Z4[&�<��"�j�E���s%xh��"��.[sdcu�%\ꕇ!�
�A'��n�1��QX����a�ȭ�����+�vI��Mf���E�I�&P7;x�d��2�e�A�!+m��g���oY���;�$�㖲��˴�n�F:fv��i��u����e�t����NMC�m��:8��Ve�0* :�3�l�Z}��lu�xtUI���cAQq5�[)����:k�^� ۚ�er� �H����/\Ҍ�t���n���,�Q�t��B�;��*��n:TT�xpE��xؽـ餪.��7"8�"�p�j� ��2��ko�HycB�z�C���v�P��k��\�YC�/c���/�r�����[��l|ϊ��A�h%L��R�F��V��c�/��5��*�=���Șm���N�5��<���1�#x1�ޮ�����2(�okmI9cGU��t�Q����W�n���7R�7D��a�w����+xge�HZ�w3.9���q�5���6R��[����&c�V��M���lL���@�i]S�$��O�;���-�}���&�fv[X�M:(չ����A���s)����z�v�-���N�*t����;G�ė�}}i6�<���测��9���D���(���SL#.�c+9�]k���9�.�}��ù0*M�,SR}/5)�Ni���8����X��*J���T�>j�m���UkDA�PDcR� V6�T�T�Z1Z�Z-jXʔUm(�,PUV�X(�cT\�f�F�",����Uh�
2�V�((�(�cڰPb* �(��"E"��ZJ�ň���A���,�EkJ�J�1�FTEU�%b�F��h�DRE��U�E��%DX�*ڠ�!X.0�����EF$�KmE,A+FG)L�	P�c
��AVE"��kF�����PXVU-b��ł�l)QccX���b�X*�EDPA+EE")��Aȶ�"�,PTF(���cD�X�m("�-(�Q�QV,PFDLJ�LF�DPTQPb"1�#F6���ʹJ�,X�j"�3���h-��5A�*
�(��"��"��dq�X���X�m�cF�J��@�~��]��y��r�r������͗q���I�.)m�r�ˌo�۽e�M�����]}ףvR���.���  7W��s3;��H/��Ow�栤P?&�{�d��%Os�OSo̝Lz��s ��
�ɹ���Ǭ
���gsRx�1 �Ú�R;�i�bOP�h�Nr�Zh�`�7/�*�Nc*�v}�y��DYN$�bIY�z�v�LH/����0�1 �~�a�LzʑCg;���>d�gP��&�=Jβy�m�0*O���z�j��P_k!��']�@׽?;���u�nw���]���Y�%q���հ�v�����M�ĕ���>eC�=�4�Y�+�߰�
�H/�ϰ��6�$���uLJ�}�i�XV6|�I���4� kDE���tGòc�I\��ĕ��4��y�'��H�u/�nZ��x�XoVq>ݓ�+����I8θ���偈,<k==�3ԩ�g���x��m1�����"� I�g���U}fb��s������eA���vM�T��w�M�^�1�C*�^�d�ҡ�H/�����
E�F^&�����Y/�����'S���&�q
�C��Yp� j-��Y�˖5�%
����~LH/C��q�ݓ���d�|@�7{�$�~�3h)�1'�3��1KCĩ�>b�}a����ǌ�&=eH���������`��`�'�ߩ�����V��-6�L�m���A��>�t�2�G���F�6��
���H�R|��{�CL�%zɿ'sg�>a_�
�w2��bI_SϬ�AeeC��Zz�H,�6Z��=LH/<��~�kᒓ�J7�U���8��YHG���HbbVw�1�XV>ގ�2bR���ᴛy�{5��AH��d�{��)�xw��O��+=?w!�}�l��=������$������[�(��f��L�;��2|	���0�%H,��(|����1&��Ǭ�T8�1�t�^$YS�G���C���N�l��Ld�\ͦ�Ĭ�s_od� ��g;�I��
E�oÑ�NZ�39[χ��B!�z̟a���@�+��L�gXI�+�ya�����!FN�& zZ,�#l�?&>偎�:�}G�4�Z�̠��P��'^��x�Y��N�kp�}e�����`ղ�k�v��������橴���7�4"ݕ:��	p��@�(L��r�fM�DM	tj}�O=�*Q�5*
P�R��M ���%�ճ*M�i��澽X$'�ğ0J�ð�J��R�d��<��Twmv~���ҟiJ\���z��<	����;�m���c';f=g��&���K��[�&�:��'��֯�
�����J��
�*E:��1��Y����=�i������_}լ.�����7�B��"�ʲ��AD�z�����@PY�T;�`q6�Y�>9��Y��N~�8��1�ϐ��x��Į����XTճ�̘�ľ��M<偌�ݚCH���/o�DȊ������5]e�H�
E��z3�'�����"�ݓ�W���ܓi+:�M��h+����~�0Yԩ�w����ϓ��&5�J��f$�yn ��)nf}�!7� |%:��ևt���{��tݚM$Ԩnk�;�N�R�s^<d��"�K̇���O�3�zs��T��M�w�<z��4�r��4��Y���$FLz��s�}�1�,���N��*>�����E�۽��q�a���Ak6ZLAO�T��U4�Y���g�y�?%H/\é<xÈcs�>���op��g��|d�IY��U�fG��A���1K���$����J�U�'O��
E*O��w�2�W�5hw���Wl<�$�|��Xy��
�ϙS_{��*m ���s&س�8��{f=a��gP8��x���$���8�`�����>�y��Ċ����O2b3�4�I^n��%B��_��Ka�6��I���k����m��8�e��W��r�q�q}N!�>9�O��}DA��}1y������j<����3�c<LK���w��Ci�'��jb�����I�+;�&'�11 �J���'�Tj��������8�N�z�<�ܓH����\�G9��y�U5bآ8�Rq���ͼd�1��N�ɤ���I�l�p�gYd�y�bm ����>׉5��$�r���T���~M$q?'�� x� �Ԙ��aO��c�Lsn1r�|��7���Ϭ�&>2��a�J�X{�uf�1���M��`Vrs�CiY*�a�hi"�I��;�z�YY+��sRg���Wl���I:����ُ��"��VA�j���d��6�[Ut�U�s�sh� 1)cV��3�ͪ�[x���Q.�rf����_����匱��ưN�l�49�ۻ�؜gc:��g7�2G��"뀺�.Q�[)j�]\;x�;[�\��!:�j��Q;&�zeb4�Z������{�Y��}��x�����SP�,������/Xx�3��H/�8�l���i%g���'_Y1������%~�����6�AH���y�?'�)s����m�������ϯ�s~r��_6�? z��M�In?0*O�㏁�����Pw����,���a�1�0�cg��UH/���é��=�xi�A�%@�֌}��{Ӡ?�dY�����[|��QY�HÚʍ���� A��<ɷH(y;L@�*c'�;���@�W�(u1��Rs�>�m1��wH)��ɉ��3��������Ă�M��:����ć���x�@K��qp~.��� �H��K�䘐Y�;��6��T�{��3�Lv���CY�1�7q"�Ĭ�,�Ɉ�7���M���_7a�4����7�a4��N���o�}{Ϲ��?p�ޞ���*N�_Y9�i�Wo��p��u1;��x��,��sR��&$<��:�b�0���n���1f&�~CI��LLJ�@�_Md4�I��Lg�߇�ݠ�E�f�]��p�k+�F� �A���~��&Ш({�c{d�i"��rE5�'���;��N�}�56�Ru���ki?!^0*{aXz�>J�g,1�a��15oɤ��dR�U�p:η��Q��߀�0�Dx��p3H<��6j�&�>eg��s6� ���4����B����4׬�� ����i�N2o;���2T%|��ړ�x��P���T4�d�ǉ<�9}��]} �[��6T���ĀH�ޓ��t�Y�F�FX~~M�ܖ�Βw�1�L�0*
u���N���g<�� z��ܰ��u&?�~NO�������w��H�bVa���;5?.��}nLw���y�zH���Ag�L�����R�Uy�f@PR)�2Zx� ���f?�>�4��=.���8�&&��I��A|���m!��O{��g�V,�ɇ�O��'�F����
P����� I���O��Atæ�����*E�g�+
¦<dǌ�T*J�~-&�T*
e��v��4��p��%�d�1<=�& q>�����q�Rq5�}ޱ?)���+��}�7ծ�xƣoM�U���ʸ8� pX��͇�H��ƺ���x-ZcE�^�Cgӱ-?v�b9y��&��ꋷ�XZ�w��wy�KG�I|5��ѱV�ֲ4�V�s_�\��g���.�a�X�.�Q���ͥ"Χ��LQt���'�}��� �M)L����t�a vg���>J��gp3�La�s�ju<H/�OMwZ6���1 ��kԋ6��Vnr�I�Leg9g���*T����v�i
�[x�d�����a��If�k���f��ȀE�>ޟ#�4�P>|��/̝Lt���w�m����&$���}�M�x���u����bAq���=|I���a\|�GD	#��$x��!���/>���&�� i+1��g�1�L������a��@�WÜÌ��Ͳb�8��d̺I�;�i:�Jɾ�z\`T�����%}|H,����>�|<=���G�O�8��؊���]}��|�<OC�M�*�6��1 �����y	����i�2O��d�M��>�2,�t�|�>H�\��nO �u�L��,yB��)#�u��R�p��Y4�d�b�d�l-�<d�O��e��i���75xλI�
�I�cm`�ľ�p�3�Lg��l�6�^!�>ɤ�:���9�=G��>#�aS�>j�G����ꧤ��Q��+7��wrT
�&��>%d�I�y�� �q��N����O�e���=d��5x�}d�c����N!_Y11��?P4�Fk�:�O8�a�~�iK~�U�����F��ޛ�z�G�m��}��N��i�����m=I��{�,���b�_9`c�1&>�OPĂ�'����
��g��V~d���'L�&e��=C���"b^��sY��b7m�a�;�m^0*CfwZ:�箒
zNo6ɷ���M0�{�CX'�w��%0/���O��C�c<�ȳ�+|�Zz�H/x�Zi�g�1 �f�ܲ{nf���3s���� �$LaXT��;��:�
�g�f��T*o�a���l�M!��bR���3�J��=�.����S���u�>$��O,4��`���T��l}u}���1J�>G�>g���|i�M���݆&��:�$���R,�q�y��6������`�ɴ
�yI�J������i��O;�kĂ�ԩ�s_jO_�%a�|�:����v\Y�f�W	�r���:�2�ӟ��gyKg� <S���@��ū�'HcIown�(������!!���t�yP��A�Jǘld]���ʁ�z^��i�k@�ۺL5#�k�����!Y�'+�
<y��G�rVL�a��J�lZ7ew�MNvr��������o���Tk��">����F"L����¢{��+�J3��I�/��`���@����#�T^c��l6�^��t���8c�R))b��dIB�}�$�8����N�:
�Vֺ��/���g��Q��)�X����}1�PA)P��d\E�ڲ��2�b16�C:e罌��.�qY\x��4�'CM[�D9ڥ|��,� �O_�H�ְ����,oJ��2;���| fםi�T�#�W8z`a�N�X���Sb�E���c>�a��;n3�0Mv��kW���� "�u���4`ٯ7T<E�('y|�ɳ��
�of]{��bu��G~7�]v�ܱ�;�lL��A�y�d�p�$��FҾh�.��~ؓ��9���P;6at��)óMe+ߔ�u�O��.G�g�\�i�P����v���$6���� ߣ���򹚵�e� �W�ؼ$h��'�au����鉬�<�`XZ�:�f�U�jjEQ��q����ȩ�����1�����`&��w�%�-��imм���y��Ŵ��z��M���P4Z�����NЉO/���'�
b�W��(�~�jaєd:[㮺:Yo�Ea\��{���J
UQI���	¯I����Z������:k�r����OO�IG��������/Oo�E ��T��7�ɗ�]����)���.�u����v$厐NO�HF��ĺ2�����^ˊ�21N������Y������8�3�I������S�nm�NÚ��f����� �E�c��@D2B3�%��A���;ι�J��S��܅��D6j���~��ǳI��'k���b��Wי�L�D {��LӋ�P5��y�-:�F0-�'����&<��q�h��5g-B���ń��uD3b�����FR`��Eq�ΐ����=�;>^=�_CBzL�jjX�(Q$hp
���zm�sJrg�xqN��MM�����9�a�������"�����: �(��)�x�02_Pg�9�_nm�d�/WEI;].�)��
��brN;jٓsP�q�q�2�	�8���|[3�p�6`ѝ@р���ν!Bt�������ܝSz/��5M����e�٧�b$8�2W$OP/��ຍ{:���Bs�='/�8'zݶ���*�F�VĈ�v�\۸h��4yao�Sz}˶G�	u������Ep�'z����ͬ{۶,�3|* R'P����m��`|6��M�S%0p�ύ䶴+mun���lH�y���E�5(�&oS�3�gMZk�1��%��	ݵ}� xt�oD6Mɐ�>j�N�(�%�q����zaN��+�M�nJqk�A�,{���k��]��t����I�K�QC.��hs�.��L�h6dLvZ�R��4�W�!e�Lo����7�O`n��M˨�����A�!���T�zA�l͑Y20�qՌ�-?l~�arD! ��!�?1ֶ�V���t��D�y>R�X%4�.�_K�]��N�^���r��]Z#�5��yC����E��F�e�XI�<�����Y~�Ln��Q%�r��Ҧ����.k3�9��9C��ł���4w��_u�Wj2��ջo�i��Tܙc��X<%�,ƪq�l��k��Z9Gr���Hu^}AAP� &;�o	�J=o��m��eԿW��������k��B�����L��(�����O6�ӻ��\�f��K�`ס���Yn���P��jyx��G�C��>5DC����r�ʼ�������RN��wDV)-Ϭc�ae�N�"�B�(�:p�4�DDOD�jz��[y\���^>�t5pKݷY1��n�N;m�Y�֝��)��ד��5�l��9��F(�Vs>"�W)��>��[��%wx������R��_F���f��;[7{q���5��9l�{��x;.�k1ٰ�biz��Q�h��o�ҥVn�U�+�.����<��SN�0P?YC�z�G�E-��Ωe��%��$��>�(ߜ��*hn�c^S���r&���o�_��M�V}R*(���� ��Z���G<j��(���WW��n�u�tZfv!�I$)�)P �9�V��!�t��{�f��*A��e	�.��Q���;v&�����*(	2p4H�C)C�Zim/NҨ��=��{�yuU�� ��h�.G͈sj,'n�乬p08(IQRN����1�9&��>ى.��3Nfz
EV>�.Ԏq&�u�r�5�Bۉ�8Yn�ǔI
�tD[�9�K�m���R�^]惤w��z�fO
�;��o�qI�&����zr�131Z�n�*��P�m�U3o�,�fQ��\`�d:tE�Ւs�#��%պ����n���y�|��ת�J�x�aA�������v�nQ�W�!<6�(�/��{E�ʐ�6�cX�u��F�7���x�!��^�q�Q��N�8��u�܀��F��U��>Z��|��שUx��s ���u����,��R6���Z�Pڪҧt�Ff���ζ��)B�IV����š��u
Շ���@��<��+�tW�iV��Kuc.K�h�u}��r`"Q�D�-}���ҋ�wy���ꪪ�����o�&�\Vɉ܁�T�`}4E���y�݌6dFQ�,d(�3�X�w���Ny�^�}�V��$ߗ��։/��
���ŞA�<s\靋"��$+�$�X�.ro��팙��
uDT����D�u���T�aҾ;��(�������5E�Ù���H`��Q*��D��(�ت�7�:&��I��:�U�b�Sj*w7�0T{�^����v�H.?	�:+�Q���"��q���<���;��s',�u^wX~��{��RN|*�4��H!�"b;��Zj���Y�"����aB���Ŕ��#��I)�X�o��g�LlAJU�&@0�}=2��U��f;Pɍ�S݀bG�y䝣nm�(��w���2#]mځ�>.,8 �&	֍�,Nne������eڸ$�8P#q��O�T�#����`a�N��j�*/'.n�f�(W�Ǆv�jO=�O�2�Z�+Є���HL��Ƞ��0����L5PT������`��K/�UӀ6n���.s@ْz��3:Ϻ���g�\��G����E�cZ0\��v��Bw3;��P�R�(;j��U��>�b���qE���/�"TK�x�h罫ïwϮ���#�0����Ê��ξ����+y�Fܨ�FDR���a)=pJ�f��q̩���4�.��8w�	�[d;7+�n�K�1�Iy�+�����p5�z�ٳR���)���ӭa�^��# 1��9����u�<��UE��KJ��>꜂|�8��}B�ʏ/Y�o���4�x�ۈc�V��ky�Gu�cv���=�~X�F{��q��Π<g�|J�W��vtۛۡ|�X=�7=���%�Cl-��^��GU69H|�<�h���g8nĜ��N3��f�ڊ����jUIu݆��8�7�Vx5�O�$���g��&��m����!I�]�i>d�e�F'����P?��Z��,.��xz���!'���:�b��ˆ�f��N���L������CG�.8d"=��D��W�1(�ᛷsy�o�*a�B��;O6�(s�Y�<�����(�׋�j��.��Q��Fغ�����j�3�O~�h�.�6|�����D�谶c":-B�B���<|���u�x��޹^M����Rp���-oV-��Gn��Ut�����CVv���T��î���T܀�-�$���ڝ�2����4�7km�9���]R����(�L�7f�+����,�ݎ�	�f������-v�㺳&1�ks��k�G��@�+l]h�D�l�e��ky�4_]�z:�t�N��uS�A�*T�)z�����YԞ�ڰ���Os��B����0#��6��������(���K�X#���`0���L�1�%֌n �k�ٓ#�A�wE�l��R��(�#Y4��C�����k)��7n�i�H΄�t]Y�j��:�X����j�k��>����)R�74�h ���n��
v����$�}�OQ��+J���/u�����r��_�y-��u�{1s���]7Z�i���M�>�V���w�΂���S-�Jʋ�4)*�0U���X�
0�Y�	�K0�<��E<�U�����od�9�\�_:wL
k�n+�&���Be�7co����L��N�3ֱ H�����P�O�Ǖ�f�m�V�8nH�6��\�5hL��C�[ؤ�f�)e���0�%S��w�݊Zu̫�5�S�p*�ga������*w���/([�8^�yݻ�C�V��/`����|9TFDδs�c�U���m)�9l����4�:=����W�Y��&�� 28��坽�QW:�jk{��fS7k(3}��)�R�7��U���!j�C�KԸ��=�oK:0�Jˋβv�̮��&��z��yփNV�םol��7�j�
���|6���t���2mU��*��Jx�
oxMΰ�A���l]�.y�8͹��P���(�_i&���*�s��1�ݭ���`+Hin��§k�j0j���m�S����wY����� ��{v��H����v7]f�7n��B�ޝK�Tl�p���g=�Ѱ�O��ҽ5kL޽YIf���)�=vhq��jZ�&ё�<ar��(��n��Άe
Z �Utiv�d��N�� �O�Ȧ.��i���;@���	���tH�88��M��\�b�B���ꯗr��N�y����pO��*��z�����uj����Ӧ��hqC��axZ}V�u1�֪�����c�
XOUv0����_NꎁpHZ�Va�;������{ۍ��\�u�7�VN��	R��}��1�E@���PSq�|�kS��j�D�1�Xen�Y��ۏXvU��ތZ��pMO/,s�(l�Dr��&Q�����J�N��>�vVO4]����u��*V���a��1Xf�k}J5L}��L�1��
�:��ئ�B��@Vfbss7$�T�e���]Gp)���9���q��ظ������������;��X�}Oq>�3���_.��xڸ6KT0�A���+`�(�*
��Ԩ���jQ2�*���TE�m��R�"����TkE���Q��V%�`�dPT`�0jVTQV�J�m"
T�TX��E���iF+�Z��1�h�QAb�a�QEVڊ�X���#iDEb8��X��c-YQA(���J�h,�A��
��P�Em�"" �be�������LlA�(�Qk,����X���A�m����
�"�4ZУD��U�����QH�����k�QZR�bV�UX���Ub
�����Q�h�b�ib�P�b�s3nZ�2(���B�Q�	-(�&4KqȰDr�Z��娨[D����*�`�Ee�b
���T,T�b`�*Ȋ��X6�Q�TDS�A�.aR*�E��U�����PP[J+R�I��)Y)�E���*��+"1Q(�#E����JZ�(�\���Q�������i�{@.�J����;9�)����Gy�(��Z���`�t�����guQ�c �p}w&;߀����O[��o�:���L��[�iU	�aΝC]qǍ���g�����;���U����3w-P�7��^`�N��ݞ+�y1�����J!���G��>n'R�m�:���Siy=��پ�W	�`�԰��y��b%�;s� �5�p��ۋ�))P#�~u`T�X��A�n?N�6{+9[�2�8�̎�@�Y�6�ڠ��nqߔXs]!�p��	]����2,>�v���\�����pu�mMI�~-��)����O/f���P斚Ӧ�� Z*qX�>|�d�]�<��Z�XIT�XÚM����|�_���=;�{�'K3����I{'�ޮ�#������N{aZ×��>4��S��g."��gU�s�l�+l٦^:2c��ʳ���Y:��Oڟ�~^�g鹗TtdE@鬚�Lڌ��̛m��q��Bnv�'���"����p�9��0��ب�x��%a���L�"ٰ���B�݇����-Jۤ�F�2�K~�����N;֜�^7f�Zm��Ѭ�3�u%�G����]����Yz�^d���(���Y�<SiN��`�`������P�X�ql�hbU����k3]��| �	:�Ø(1��s~ӵ��ݝ�,9'��f�jP}�k�Ⱥ���	(��QE��j�'N��{�m{�)ZnT�6�k�R�*���u�r�ʉ��&��;A��i��)�A�抾�{;b���j����bT�U�Pc�+������M�0�{�� ��0�X�� �'`(���Ӈ�d1�F�¥�Qs9f	fxI��)�V)����X{���}�c��7f�m���w'�G?%�7�ƋJ�0�w=�T�3���YF��]dξ�����#�9�zҰ���?$F�)	;Ϯ��|g��w�{2��Z�9��$��@���r�|�;
0B����́+\Q�������33�c%�3N�m�~-�v�I�ˇ6�(����T��[��t6b������&iK���ν���.�4���Ć�.��fr��s��P�k|"�۞�t)��J�Sո�6�p��F��]�Y7�����'GL��]��/q]ܧ�
�k'ED��O:-�KZpWw�u�%�o-̘��ޕ����� �"�������v�Q66Wr�Da��p�ev(��LZ��V�.�xxc��1�e�����M	�쵕��XIT�2�Pz
$�J�w8��a�<��1/C��2�[����X���XZØ&69������k��y���Ŷ�x�Vw�9���zm�����g�ڴ�h��/���U]�c5v�\����+�pc�9�![���8���l5J#����&{n�^%a̼�r��<�z�ō�d^�9 V&�S�
$�t�Y٪�]؋�G�.��+��ƣ�5�&�����kgf�R�pitܺ�U���Ҹ*��bzU	a��_0o.npSn���|֭l�K���z�B��4뉏�^1������]bO����sy��X�U��>�'$�k:��l�D�=�A|�LwT�J�)��i���y6T���qreY��hS��h���Ӈ������-*�#Hnͳ݊�\�e�9�/<���Θ��(�5L,�.Љ`V�'����)^' 9����O�ǰed����p٫��0^f�l��p��v��=*���[A
��%'|Ɋ�TP��y�ђ�[BtK%���0A%�������iN/���g�?� .W�6�bk����,�9���/��E������?%1�
B��o���z�[�v�]�k�m��
�݀�wݡn�P������5Yd�5)M����ԄV��,bM�g�J�ɤkh����m��'�D�����w%Q��'����BV�`NGf�\��o�@�q^*J�J�}5Kb9\��czq�m����O�k�}yᖲ�YTuN�������
��)zu����e��$6����
�9�/��nave�S��>|{���ޯ��x��M䞪Nn,aO؆�����k='V�̄��>W�+�P��Էُ�B�鮮z�i�ޕ��9���45��Z͊z�\��n�v��L������|�]�����Y~�O��r�-��"�L8}NFm,��Σ,���t{M�ק���z��3̎�>U]�)���i�D���9��@!&��,�`���O0tＢpU��]�NZGN�s�3���-y���t��e+�vp`�q�l��6-�M�q�:��������e�%Ø�X�4ǱH�'[{�z��̮\����4�3I��n��	n&���}_}]�sϼ�Q�ꍼf�,��߳��P}@��|�|ΓON�z��O[�Ǡ����l���W�������1�pz�!�F��83�7�o7����ʺ"�X���m�\��;:���wH�����;��ޞÐ��^{�x�m�~v������5����vvu�8z�D����>����Q�6���y\j�}z����٧s:	ݝ;���0N:[yf�l'=ї�̹�����z$n
̝l)]�V=����"k/��Q��l��l��O�����!�>��&����*�!�T�9矛���r�]�xfҊ���(�
�����>�Z�=�٥b��w��f��͖s�r߅掔=j����s��XsC��Gh�s�W`���K�u6M�K-����g_u1�Щ�T�$˰[�E�s+������>5t��O ��׎͓�aB'����T
l��A�/K�d�	:=������;���`�S4�KgR�z�Ҧn���lvq��Z1a�H��F�u������Y�5��3ggq�/8���,���9WB��M[h)9�
M���>;�+��=�=/��s%�]gt,���Wk�~IT���Ɔ��0s=���*���oy�T��vʲ�\u,�heի�u�േ/%N�4*F�;��8Qo��N1�:���r��]���y�w�_;y�ߧ�þ����b>m�;u��:��3��^��g/��I��b���O3��G�����o�q���4��ы�q؟�����{���$��l�� �);�]3ݭ>s1�p^#P�2�� �=����[;~�= V��2ob�5 ��յQ��|�s���+��Y֛�ۮ&̈�Ɩ��^&�b��+�'(%^�*��7v0�X��y�N�vr1`떦�9����Th�����J�S	P�i])������ݱ�*5��g0�ثf�u�|�^����������6l|}"3�M�̸���r����-�|ݤ	��e�y�Q���sb1��V�z��TBg�͗��Z+��S���y+S?��i벞������$��v�����p�٭;ف�m�t^R�'[.�}K�J,��1[��s�LEYr��{�p欴��>���s���,D�;|��S�=�~L�t����){y􅔳}�L��o&��k���ԭ���O��ӊs��(�
��R\��Qu�*ܽ��v�<���Kd<ҫܚV[��j��<.)�Qa�!}���К��e<�"���Y'�NvW�Ҭ�K���`�%��n-�b���Tf�3�|�B�U/!:l�����Z�׋�J��&f���mЩ</��be&�O��z���GQ��]��p��+YՊ�s��Uo	�2V5��(u�,^�����hk<-p���G8�ߔ�zezm��j}��{5Q^Ggb�B��uP�Y�8��̑
�"=C9��7���.���}��ƪf,�ʟ7ѼŎ����f�V���)�-i�f0璶�W��z�y�c`Cd���e���+|�q������0�c��ӯ��2`+&uèT�P�̏�wԪ��J��U�NĖy�:<��u�8�YV���֫|��o��7��ye���EbFpY�y��Sn��\�e�^�l-Rp$F+�D1��r�+�����Ҍ�d�-u�](^��b
5%������'��uq����nt0�Z_$o.ns�ۧ+��Fb.s*nި��x��9��������X<�Y0�KF)u�A�As��6�qL9��3Al��x�{���gZղ�R&�_(=�%JlJ����5nN4��%�XBn���cx-��vv;�Ӈ�%lh��gť}�V�/�N��Ɩ�TMeWM:��.���=}�������Ӆ��S'��5X�7�/)W�v�C�@�[@�]�
ǻ��պq^���<�ut�����[V�-�>�~1|(�T���f�@ri_��l;�N�Q� �E=B=�6�f�.0��Gn1�b:���CS�[��>�+G.r���in���z�\��D0��\�mE�Ω�5�R�ԁ\���2�P�eu>��i7��S�&���M^閛�]>��C�9��Qg(tH�w����5V_ކO9�{�6�^��9��m��B����v�8��f̨�v,Ȇ-p?�n��.a:�<��	���y�iN|U��ӟGyQK��pj�{W���ms�՜2`�%_(��h�/!�AS�]��Z%
�]׫�'��w}��5�5�n�g_e|3k9��)�����Ƴ��=���mt͢��};��y,]=�x�깹����ְ���&����X�q��.�]���W���R�`�]��%���' VV��L��r��K��V���Ff���#�Ě��Z{�<w�1���	�{�z�S<��D+Y�N�3��6� �T�;z�����9 Yes^\��?��C�+���?{�9�F��]8��ny��^7����y]�=~U-�bVd�-b���������=/0h�l.v�n>�δ�˺D���c�b��y��5���S���fا/n�k1��raGgZӇ�$Jt�e�)3Yp����O̯�Y��{��K(I�a���>��7����$�:YU���E~�vȍ
BAiW�P�n��݅c��&0��0$[s�L�1�q�Au�=\�����S~���WL-����`���^�̱�]ȣM��zh[�wn�I��TF=�u���)�bni��n���y��I�-��u4��Pe���|��l3�a��b�#���Q���cŵӯ��l���xxv*��a�l��F���C��� ��\��F���z�A7Z6�r�n��ʳ�����ӊ����,BPR�6>����u���Z�.m�me�W��y��|]��Ru�[ТÚ����/-����܁_����nf��J��ЗtΎI�e�-t]�0s����Љ�*GA�Ѩ�x@~�W�o+�밒�XÞM���b2�Q�̺�š[f�?�x唲�]���2��Akk�)I�s�cFQ�UW�(q�Q��EL��O���Ʌo,J��J{V>s������3Q��4�z���-~Ҧ�v��g,s9>8��9���k���@ʊ����=��W6ڙ��1V�eu��X��̜^Xr|+��T��W�o���Ono6TU�h�~��Z���J{a7�c��g�W#�$�א�D�Sc��Tl�v�3yf��ū�'�]pU�X}m� Tyu�|�c&Z��Qc]6�,r�����q��5�s.��u�ұ�Z.�Mon1��Й��Վ���d<T�n�$�rSLH~#J�1�����������z^L�/Q]��; ݖ���� �7PKQ���]5�����o�Y������u9�Kq��U�+Z���6�[��_c<&]��m��4��W��l��k3*[���'H6eժ}�.��8T�l�wOa62���|0�_k���,1����_pZ���y.�5A-�CM(]�D[�x2X�'&�6rH�=q�h�ul���a�(��&%�Ģ�g
ʴ�`]����[�\3�Ħ\�Ԗ)�[�B{fv�<aڰ����I�]6y'��\��*n���!��'=����R'4u֪�,JB]���N�ÌT��F��;���,r�|©Q�j��]���_1��JA�:���u��E�>���'��]�!��e�T�cSu�ݰ-(Gz<��ׄD�ˤ,�F��Ȩd�]r코�f#�vn�IE�4�m�ª��g�@�۶����	�P��S�t��ݳu[>L�:��VfY.�k,ܐҲe���P����9���KF(�Ʒ�W]��t���h���qi�S������p��^�����#�^z����J��l�k���[��իzNGd��9��ʜ�0�1�)j�1�v޳V�ו�`�D3r��N�ҭ������J�zJPN�n���Y���2TT�(���PG�p�WPe"�e���ͬhhщ)e�u�
�0�[Y1cLӝ���3�m�nb��e�X��2�������� ݻ��y*ۻ�"�.T���P�ԫ��Wv�]�Q>Jm�7��ͪ���� 	;��cѽ��g`sqV�g�hI�6l&������)��Lf��N]�\�l���=�^:�=��Y˾f�i���-��w!5X����bwb˚���Z}�[i�2[�i�*r��:J��i��G�6U,#q��c[׹��k�D�tn���{�E�V�U��ޢy{�fD��!GE'�k�G��+�zS��gKxFQ�ou��Y5�я���=35Er5���te��:��Ļ���9�|���2Eױ��in�Yf�ܩi�t�aW@Q�o�L]��wb��r���-��[��Z��s5IuNϴ����V��ՙ�A���a�1����kk���y�&h���5)���k'�;{*PդP�W�w.�v
���j܅��ιf݋�X6]�%AiA�n�гܢ����qwwP�ja����{�����r���Q�'"̖Nâ�3@��G|���A�j�����X���+u��z/�����web�6yU��m���f��y�+�U��\�v��6�9�W3���f9�X�$!Q$�	 �QV����h"�)��(�U�eV,*��ʨ��Z��0����E�*����-
��"�Eb�5b9j ��+e��+��A�1�DU�Y�˙c��&Z3*
�m�b������UB�jQb��+�̲��i�3ۗ2[DKLpW3
���R҂��Y��+13
�0�(�eeJ��EAQjJ��((cH��̬DDr�U1�ChTb�DF*EE-V��UF�(�F9l�J"��B��DbEVckTE�±��Ŋ"*�e���h�"�����Ecl���(�(�b���E�"�X ������b�1+QX"��5�KJ-�DX�
�J
���KUP�X#YUU�+�JbQ8�bX��Eb*����e���AV�KeF �ff)�Jʙh����*UQ33Um(���R��E\l�(�?oF�KR.�ŝ���z�Ti�m�D�I}A-�b��N;�$7�7I`�����f����@�5x�u�4y���<�u���\�N��2%_+�52�nW;P��7��9U+o��;�n�;\9�2K3�F;k��	A*�*������6��R|{�\��J�t;�����:�M�a"Go�()!0ұJg������+Eᦪ)�'h�~��W������4G�q��L'S��Lq��Z	����+��M�=�H��eo��{I3e��L������{T��s2��N�S��ܱ�����Ci[�ո�m[��4lB�佪s	��]��S��̾�.Wu`�٥�&���~ڠ�<�sn�Xsz0Nb�ŗ�JL/d��C������/R�{wI�wB����o���F�*{c�Ȧ����<ʁ����ܲ���rhJyC-eת�U+3vO9�^��p���Z�����^�_����^�Q�ihup�2�[�쵕�X���ȵ��Z���M89%������X��c�%��>�+�Ŝ���*�w��Q��]�� N�����-�����d�/n�R���Iں���z�g6����eT��A�}�j����9K{Yt⼗�'P@%9D+�N}]�Nΐ�k����]�ݷ�ﾮ��I��u�_�
i�!4tT�k= ����)俗At���k�>l��fo0wdR'���{kX����p�7w
���>����
���齛�-��f���Xy󙜌�����=����l#�+Z��~1뱸ST�M�-�\nzy��2�q���S/n�>{�t��G(�n7&]^>dܳw*�x]��W5����v
��}����m��I�[8��T�C�s=Go_���o':�� ��ug�T��(z �v�!gN�q㲷sk���dF��r�R{O\�%�C�`�ˤ�^���X{����f��z�"�/���/�raGc����H�tQ�5�+r;#�9yt���	&{��oy)���,���Szl���:Hu;GX��_0њu3�A��V(=�|�)]�X�p'�n\h�����'�R���Ҥ�qfJ�Xds�z)F,�4%W�+T�7D�Ax�LXp쮺;e+�KN�i�;6v�i�rʹf�M�0f�|��n�PǠdml��ZPc�dG�kYۥ�;��{c�����+�u���D*�R=}ٗ��(���	�)^�n�ɞ���f��m'h���rF�o�8_l*�J�w��/2�Z}�q�D���f�Byd��~�nË��JU�4'�r�+}�V�\���oA+Twf<.Rz�ٱ�ͺ�n-�Snx���j}\Ծ�}/�Q�����=�wB�ʄg��N�&e�44��DX����O��l���gs�{ʥv4�d�]�02�P�Y��g�0���>i�3Y�V�Or3c|�;r��0��G!�/�}Z���W6�yJk�4$4�&s�-٭R&p����tr͙e㣙 G[�To19��]�}ʟ<��rD�B�n)��,G)V�sY�M�(�G�+Y��;~]������u;S<�8�ِ���i�@�C����a�ݱ�vv�ÃX1�7��b<'���G��+5�I�� 1W�	r�{~M�={`U��y]�Ba�Y�lJ��:
��4j@�cg:�j��S/Ep�jhq
�iq�"ת+M�/PE�X�>bq��c��b�-ݖg^q׹W�Ľb9]m�S����#]��M��DG��;�l!2Y��9|1�cC��|X�}��s��Q=�^O]�)���.�l���Bk��a��_K	�A��`(��	��b�0y�P���������Rn��s���U�A���1�!4�����i��7��N:�����\�a�h�~;���R�Ry�sv�0��t,P����ٔn�V"yڎ�ƣ��?%"4AHIiP(	��]�
ǻa������]��TE���[I;���H��◵>�Al��uuQ���b�֭�aZ�>���3T�_s��^N�P��ѡT�v�:��s����n��zyN�4��%��o���W�����4�=��Fn��]��g�w���=K0��6����]�<�,4lS�s+�9�ʩ��pg�b��W��r-��yAs��Nnܼ�z�$�V0�l4���_Sާ4��\��1����!+p��^	V�U��:Vo�ʮ�W����'�[^b�?��y7�@ա�gqR��CIRu��&:n�]�RT���s*�J�=vM���V�v6��X�P3��	�WM�y����ח�V�qI����Nݚn%��f�k�ޙ�(k[*�jGg:��]|�f���лmq���>�%n��L��/X�����5����S�L;c_�k�EQ��V;��.����UK��;�l�4�/���X�rN>�s	����9Y�[�
�loS���O���W���y�';K;�gma����9�T�	�Q�=;z7[*��K��c�����ޅ-<r�oɽ�ƶvh��p�%�Y�7�u��f��+f;jzUK�2%��Bo�npSn�r���������UUX�w0��5*i��`�F9�}��X�n �߱���6�����S
�3��N*2����`=8z�D��_*��U0�G�M{�\�Z��[9�Y�<��)_1��O�X;�8z��� �%�^���qx��7��eu����u���,�z��X�|�a�+�g�?%06H<h�1W�1����l��v�PͶ��6�����O�ܸ��i�b�y$=(7�Gf��Uv1Ն|�B�8\H.g�k=�(.{�3����`�TL..��L�@[��M��}�c[��	j�Y1�s'aS��i�����c�u}�����:]���9�e�o
W�X��m��\E}�]ЖUu>�quڰ���jh]��<��.`��y1��=�٥ri [��j�N���qspU]9���bU�R��uP �k����-:�	w9MiL�;/8b��lrT�-�B9���czq��|�ڑrh	O(e���gN�kl&���gn�v7Gz��2�B[Pg^�IuKh�/��ҭ�Zλ#$���)v'�&*���<ޮ�-a�<B$&��蹚�zG����S��듴;HC�U6zi��x�=�^�NkA�N�SX�.��sN�]�v�n{�s�A����ܻ9X�M�W�Y~�O��|���W�am�Qy%�
����w����y����L�!��q<��x�ɼM����RUq��|�I�>xΛ�i�އ�J����KԌ��oC6z�^g�A�w��ܶ֫��v뉏\��}$���yo0㙑����&zn�Ĕ(�׮T'�%8v�ԉ�Ag?���7k�s;���^G9z=:��S��Rl]b46E�O>�����`����[��I]z��J�?���]�Ǐ$�\@}w!J��z"t�,ͲGX��[ܢ�^�F���{��֘�&47w��t�&�_,�^�L�>Y1ݮatV�ٗ���(�ʮ�`VN�;o0kr�!4�����6{�%ӆ���5�۬�T8�؊,������*����g���}�M�7�˅4!޸��d�V�2�wO��1 މ������E����U|��y)G���N�f�}<�`��wD!�Qژ��
��rF�)	�X� �}}���J�w����.ݲn;����jn��B�"�~ͥ�m߂��))Q�[��9�U�pfgz/��"b�����`�u�.��fs^�)P���/<�^��ieR��N�)-x�=�*��䙞m�iE��0W<s�k�j������x?����ig�:����*�Y^άW��hyc
h&�H!>}�b���V4t�]�y:վ��yJ픦̹V���$VU�������SA46�mײew��G74��Y^nU<g�*A��yK[��M2u�S������f^�1�,�o���mg�%���������p��� �<�e����Gp�hg�<�b�"r�#�-܌-F3��u_#�:�IX瓛�8C=Y�S8TV�Wo3{x{��m �E������9&�P9��y�g4l��鎪n �������s(��J�zL�z�-����$W@�U7;S��B=|��9�#f#as�bU�1t�'u�o:�=��=���Òq]އ=�\#��!���n�s1�.���!7��JV���	�W�co�g�Ǧ_�t�
�
���*a
T���OHzݮ�<5�D���b���mӕ��vro%�H��ْ/F�kۗ�t94�![���e�t�bհ�߱�!4�=|u��A��H���&��q��N�o���	��b���T�g���`c�6n�k]��rѹ�;��'��p^JDh���ZPVd�t
��kr�/�1l�ݻ���*��,�n�8�{J���"3A}�v���&e�1��23a����A֤�y�ˍ����,B���6(o�`K�{+����w�M�Ph�n
�'����*6���ou�&[��c{��鷺k�gbP�Ӝ��y։��|(ݥLHJ@>H����z�H�&W3�5�@���r��dU\IN�K�����Z=�������5���/�N�V��v��}��}U_S�O�|�N��W�Hy���o���:���x��׳j�Ղ�F���x@~���zue{-���TrL��-t]y���9�4��*�z�.�)Q��c!1�b;s.[̥xk�a%SAch���㊲W;�$)ܼ뇦�/�_��k��im�S��*�ެ���{κՉv��p����AqPP�06]�)��J.f���m�Ʌo!Q��[���A��mt������m����K���7��8��9���]�8'��r�y����f�O]��+S/Vy9�X��ǻ;u��.։;W i�u����W��o09r�t>��Gb�QϙP�N]��&�o��b��6n|Lz}���^׼#�0kn��㣳҇u{"]z�!7�79�~�׳���\��Fq&�3��;	!E�l��<��r���(%C������ȳ�!�J5���7��z����.AF#���/mv��B*�ugZC���ʊ��cU�Y��ޗٕ2��CT��V��][�:r�9U�}$hU�ɔ3j�Vea��gR=�p,�k銰�['�6��腋�,��)�:5(t�Bf�{���k3{�(ӱv� �}���&Nټ�'�Xq��M��$H�_()d�J�I��۝"��뼦���A
���i��o�S�W��ޜ=K�Lh��CJ��"����k����݌�g���J�7݃X�|༕��L��T��퉁S�ۮO�zmfR�,�b�l�-w�~qz�<�mt��i�b��U�,�Q�ե=��,� �tЕ��.�ҹ>�o��]�	�Ί��T�w�V�w��P<��tؕ	o���N�]Nݹ��*]�h&��+���u���O%c؆�:*�SNq�
m�����&��/���n�wQ�%�8z�t�4�y�&Ā҃:��u�����ٖ%[��C�q!�Ѿ��|����s�~�ey�)�/�.f���mp̩��PB�vs�Qm��^Et�q����j�����/e�<�-���n��[�'TVM9�	Z�4��c���S0��c4����'��KXt�����O�G ��>������5F�@���!n)!��zfٙ�ihoYE���׶��\嫫f����ۄ���h}�9�ѻ[�j0%��5�z�Vr�l�eL/���c鏶Q�6`V@++���)��OsU���,8����=(��|뢻�n�SF�;�T\���xյ]ز.��M�+\S��qg1�u҂�����eY�j�;kT���=��w��կp��0�1��d�7xIӇs �&����=#cI얌�WhUԧ��-�S �٣�x냭��lu2o}\��n��=�e�|5F��e��[�^T�}5��PN�V�)�N[��`��y�w�XU��=��C����A�]��R@�.C�Eӥl[������� �b��A.P�W4^<�����3:���U�36��ɴ.s��Wq�6�K��%q�3n���XfV%/�N���t�
)J��um��m0��o�Ht�����f$�N�'�+{����̩Yh�W%χX�#�TF�(�yC��jq�0��+�$IX������5!�9�8�sϵ�x��Γ��˘��8�O��	tI���'�x�6Z��`�ŧH�"�H�'=��-b�j��4v�R�P��ȹ�7:�b�
��7����u�,ƒܻ�����R#��0��b�5K��v,6#�r��~N���Ե�:�+;�-�]c�����n��2����2��i6	��c��)XY�
�m^l�X����{Q�eP�'U��v+�ݲ���k����@Vs�g�Fѩ���65]��ۛ�L�cf���̎�46�C&�t��z�|X�h)��lCeGmD�󙺲݆�Nn��:�BԖ���#y"F��{�q�ꔜ'�{��������eS-���,��i�%�z.�'���9����M�K�C,`��ז$��L͔�$��+T�&�?rKgoc�X���_PHI�ĽƉ�
bf�na���[F�J����%�5���AZ�r�酅L�lAu�M��:Z���l=ΜiL�d��m�R��Q��P��k�f>��b��R��am��煷��\�+\zbK�WXڜsCd�����wR��[U��v'u2�Ҟ)�J�*�����d�%��C$�VmX��F\a�����2�;���]�����pTb�s��0��`�9�w�����!�$��%:���4Nkc�b#ʓ!̛��.�)��y'9`9ku�',���+^Vc�h%;o+�{�G\ř*�K�)���t�u�"&�'B3��C;25��mwCRdS�w[�"V�ޛ�w}gV��"��t:"̝��d�%fL�X>k�f�K���%�&/�V��ԔKb�-[#/Jt��*��{9E�kH��G�����C��J���������٢��Kr�����SFc�k�	��OęK�HD"
6**��.%1���
J��3���\��c�Q�W.8��rܭ-kZcW-S��T2�(&%m��*"6ՙbª�(�DJ%�����W.&%jc���3�J9e��2�X���Uƙ[(��ع�2کF�V[�.\��m��-��1X1Jʀ�bU�%*�LlL��r�TX��b*5r�⭵#lr�
�(�(��b(�&X�\��J*�U�+-*�Q[��I[[�X��m�%�cs+c�(�Ѷ�QQ��D�V�Ymb�2�C2�S���l�EDQ�ƱD2�EV�H�m,G�Ģ�-Z���Qĥ�D1
(�!*@TG)*(ƥ���6�e�DEL���˩x�rpd�����u���l�й��op��YԺ����#;`�(.���%���Ҷ�n���]D�̂N���K�'U���]>�k�	Vr�!6�tB�9S珥�^���}c5lTr�ϛ+*g:9��rN;������B�i:��R�����7yaokq0�T�=z���o�٣�+�ޯ	s�(>�_F�H�}Q��R��c��1u��o*We�Z���������PI��Kr�!�b���#�z������}l.w��p�GoRղ�R&��xW�(�q�9���S��w6�)��M�kr�0�I�
;��RD����0$�v���®Z��n�(�}Iex�O0s�ݬ\��A����;�%z��a	�4QO|�} �$��(-���wg�Ǻ�a�	��s�ף��ȍ�q�������6HIX�[]����g"�ʘs�3CbaY��g�(7O.۵!()i ��BV�`LdZ/��b�����vĩ�
\&fu5|J��cK$:�Ohr*�bT�^��X����[��Af e�8-�<�u���E�F]�ogU��[�+9�3k[;��$!z��m�欇l۫��!.���n�u
�|O-���s�w�����R˪����=j��78ͩ�5�R��V���!f���yfZW���Ge��������wܓ3M�-(����������F5׉��ܹ�2�Vub��SKSI�!��E���H7fk;��1�VٳO���Ʉ�,	v�Ƭ�ʵ�9kh��F]��6�^ �FmF�z�&m��m��"��F�؜���X镇o�8Ĭg��N�;�=P�bi���.h�w��k-q�.u����5uE^��=c���G�ֹ�S3Wf*�ɕ�
^�	������Y:Ū��9���08�4����xtM�h���N��~�)Z�{a7�޽��VzO+�;%�ň��u1"y�^��8�؈Ps\�}�_$_"��M�r�ߔvu�&�ZåB�V�"
�Kx$f��/��u��2��JUA��cf0��4��#�L윇"�^L��Fh�{G��6��P�"�_a�C�i�|���i�����y�c��y�بnu18a�Y��f�����G0]���%*�G��Ҭ�e�ǀN]�m[k���`lIL?�Ŀ�z^>����Gdw��Z�9�c�Q�A���{f6�zN(���M��$J�F�/�L%S�R��;|����ހ՛���9�FU��[)��W��:+�/4��*u�`���<a�_E�{�P��;7o��v��H��{I;��)��R��������Q��SKc�nfgr�K��Ŵ���`��N�P���(�
�����4�����y7���}j_����ݚ]r�ž,:Z�E�s���×J�x�NO������=�m���#R���Yi�wB��SC�eߋbZ��Xдeu[�����z����C�N����*�XÖz�Zڮ�V'��Tn�z���4���Z9T;��'T�gڴ���ͧ%J��U��*5Yf)1��^J�M	�J.gY�Ox���ʳ���'�#׭�.��#��X̤���pO��_���^v^��g/���~�R$���W@��
,�ӮN1��}֓��sq�oH��\ָ��zeyd�Ǯ���3����VI��:���v���#���.�ђ.���#�qff'��*�x��&��|�l���b���;�$9g%kV�M��$U՘�cl�s�qmI��=��]�%��@��,��bs�W�����5%2��	�PX��y�f�Za�!����~k��f�nY,�.7���!�\O>|�O<��XM�Q=�(M�����l�Tj��g��^5C��JՑ.���7(Sng�f��S��v�J\�Q��2u��v뉀.�L>�A*�+n����ejV��Xr��8�|������g�RD��^/�	����b��5��s}�b���=w9ۈ,�0��&v��gZ�S �b���l�<69�v�!��Y�c�n��R��u{X�|༔�g~J^u	\:��Mɍ�����6�D�LI��b��範6���[�>�r��K��sq�؊K��RNѮ�����of�k��}٥P�Ұ[���ڨ�c��L����B9d��;�,9������-�����
�s�]k��7<n�S�ŚDJyw?'Qf��]x�ڞ� a�=�oz�j���&��7��^���ٵ������K.EY���xyέ��+b��\vs��Bm�8�j��8n�瘳�d�(�n��r�Úq}���.q�-=�aU�<��öm��Ho���l)�5��c���M���o�3�=�`8�o}�̥X.{�oT�L� �J�zpP�Q�����a�a���������پ��c-������_��������3~~�G�׮uc����r]�aY�lK������Xޗ����˗�4��g���0�"W��}��/�t.����Vr�	��GL��T��KTmMp6^Y\�K��ǳV���(�G��Z�~�Bnv=��_.5�Б��9�����!�z��㟧yC�y��X���k��pxEY�鶻�<ʜlj�y�Zy�����4��Ĕ�6���kU�ogo���<��cUL>�������ɭi��k)��;^��h.i����(��%O�hǼ�S�.UU�C�#Y���������+o3X{�1�!4�������[L&��)|���x��_RF�r����J'g�=%��E��x�����]����nu��5�c[�����	�%�hp4�܃^B_H)1k�.9kh��7���;؊�Нd��n�s,KՍN���o��.3&���Un#����Ŗm�SSpu~���7E>�}ֵ3�`��G��#���ש,
S���g���)�G%�LFAP�#4�Ln�v���S�R#D R���-�|��T���{���bťZx�e��=�6����<ߛ����f�a^�bN\�!�l��,!7vf�]n�̯'O/����E�J
ZF�O��n�U���޻n7��3�6n�����]�j�����l)�5�R���B�*�w��S��2�:ae������.�I��ؖ�] �c;s�Nf�,��|��T���	��_d�ߑ�j�R{s~SI��(MR�6r)+����1���'V��	V�Ƭ��Y�/mkE[�V��%W٨�U;&r]��̙�k9 }@�H�o�U����N���:#�iN7��j�YF'^m.x�\מ-�Ov2�H8���Ss���{|g-	�=�oh^�fW�N�N�D���Y�JB� dI����=W�pz���"f>��~+&GO�݌��<��8�|���{L�X�tVz��湃��tea��_Wa9�V��6)��z���&�k8��Pᕙ�p�}�iᾛLY���j�[�Lw\x�3��t�i���������f�mZ�*ѸQ�\:��?z���K���X�z�1����)_���	�Vױ��ù���0WjW���uzc�K�a��BE�-M��9\��;:�j�=r�@���SH)<�J�b��)u�Bc���J��+n���Y�,,mb�����u�}Z��~C�;E܄�\>r�)o�rm�.{r��Z��_<\5�peY��)[���w�R�R#D���L,~WƓ'�*�;�J���w�l�ߠ�*tV�[ɂT��CP-�%���^�u1�Un{����;���-��V]�X̯'N�z��%"gl����F�z�W��<���viZ9sA�,:���.�nq�S�r*-��X�$�J�\*_��jc��	]�Iﳺ��I�e��Hn�[�O4��O�yX�H��g�W�d8���
�'{�Pr�t����[p��8  ��q֥x��욙Bé[�J�,�E"�ʛ��b"
��OWi��]�2F��?o��g'��[NW.i3Q���I���n�{�,� ��!��J�������{������>���)����׭%3YH���jfki�1f˽BCj��(u��{�jѾ�+8��ȓ��ƍ��;�'�V.{��oV�Z×��|�ҋ��g�}G2D+x&̮ �L�W٩�=9�{��'��^��߾��U�_�=��f��j��wS��+t$TV���P��r��@�z�t�+
e����,X�cݝ���ݼ�"�(���W�4g,�e�<�znv�,>�+��ϝ�2��.��tr��#%u~5�����$7���3Znev��J�2%оM�Mɳudd�a����w����gXM���c��S�K�A'�+�~)^��=�:td�ݑ��	e�m�r���kN��0{D��P�J'M^�t����5�58Q5�]4�&}n�y�a�߱�4�����7;�;��~Õ�s�{���z��I�0�@�M�
����ssZ�g[�k\t�X�L�T�'��m�ΞĎ�0N�O)�(J�F�p92�vom�4ª���Qɋ=��1)\4�`4���'G�������c�����HG�.8�Ɵ&ҡ���/9����߻7�7������`RYER���_vc'8�iZgUs�,ٸ�����I6ʙ�>�p�u��d_=e���ո�t��\�QH�>A7]���5ۏcuyy/m{5+]�t��J�M+-�}�0������-����r�]�6��(�����s^��^�N��О�Ng�f��9���[&*��K��*�lHk���l)�<KZԈ[�	�[�7 ��9]s�˚��F3o���j�ҩ����ؐ҃�M�j:�-���I�4n�_�Z�'���$B�՟�m#�L<������׈D�4$>蹚��!�T�*�#����
�ҫ`�[��K���沭^�����v�\�y�r�ݫh�9G2�-�h4��PD��ץ$�q�9�����Ϡ{ʟ8�(�3��.�ۻ˶�*�Rgu��`=݌��䃊��s��z��t�G��qx|sn?^�cm�}��̎����K���k���8�%�h�mDmn��y��ŏ�୛�&���ސ�ȷ�U��Y���]���!
����bӳ8��ݧ�����Q$,WbZY�]�������÷�[�)9�ٚ|+�Y���������)u�Qt�'qco:�=�ƶv�VzN+��W��8!F_QP��ӳtEx�����Sn����cy9:O]@�+7�r}��{/��Bw�z���m{���As�ۧ);
;:��l��"r��n�̼��?2]z��4s�/wG˝Z��5��x�h������p�wBI�\ɮ�E{��� ��iA�z),�U'��_vk�{���:)u�M���g:V��t�:(����B��.7���]�`=몹�'�Sc�jݷ.4C�V���ܑ�!@�����i58�����Gsa��>�~/�y�˽ۿ(�	AK|F�)�� �i������C'z�����C�9��=T]78ʊsĮ�R#��R���Z�q{qyd�'�V[��eR9&f�bZQt�cx	�K���ӷNk�%
���r�IVj/�ђif��{�q���)�eF�eЌN�T���fۭ�Q"�MH8�`G
H��y���rxy�o��]|�C^�T���rTui���B��o���*���L��%���t��fM�=��u�
]۶v���(]�1lx�1B(*�1����Pw[�����n\y�srԒ��<�m'�~�{Ք�U���JN�}���=��T��%՛�[5��|�� 濲��m1�lE�M�ˤ5s��V�E�zd:�T׏&��rL���Aal�	�Z�fn[�`::�Y�a��е��v(��Q�yh�[W��6V�uM���h}Ӄ��U��)�����M=c:���5p)R��Dʃe�J�,�Јzъ�B!���ɂ�@�����k���EE3�^l��M��"�/ӬڻY����'�o3%J�+P؟)��]_k� '��W,w���P��[Dm}���T�)��v��u�/��W<�$��b�V��I=��t��m=[��,���½��Sf�]\��V8���r�b^�0�;�󸹘��$���gV��@u�L���oSW	�[�,O�k����JU[:�zj�T(u�I��
ͳ��Ya�ZM�q ��ǐ�����Gg<Z�ʴWD�����b������'�=w��gVϻr) @�{r�.��י,�7"���ZG(�ni����#6y*F����S�NQ��l����N͢OʃQ͟Gخ_[�_R�q�=����gc4VCRmu��ٮfw���X�?M�v���I�=�6@궷�#����ip��P#�*W6OYW�o%���8<�!R�ݱZ��H1R��jo�}�u��7�h����Z]���c�7U�1]����!�x�6x�58PƢ �VJE��Y��u��tAn��oj���2�Xm�9����쬨�Đ�Қ�t�&u�O��1�q��f�_^ A�޽v�pё�#���9Y�o��`��x�&�1��Dn���kV3$�W�'�jZ�iȣ����6�gtw�=��$�Q�2��a^��LʘWeEۛ��Rv�-���JY�'���i�4h}�
�1��_���`[!�bZ4�"� <1nZ�.]K��S2L�Qmu��=w�l�V�4=X�q号%�yP�w��r��� ��K��Ϋ�ÑwsP��z �i�Z�jv�Q���{c���k�p��tu(�@C�2������T5S4:��L�3���d��ic�IXQ����0.����@8�_C���i'�),�����ְ.cD�i�g�l-o)�&Z4���v�s�p�#wX�D�n��8�j��w(6���:�:�Ѯ��y�E�Nu=�9k(,�|(,����λ�'�D_	����e���&ोi[�	Hl�[��uT���N�1��*����z�2��� �'@�I�W-VfbU
�c��a�Ģ"e�,E,�&F��K�b��f5-,��QPEfXb�LJ�زR���
�be��°T�U3&*���33�lLJ6�Dq����Q�PUDH��֥h��R��C"1M6(�� ��5J���X�Um(�(��
#j� �P�隶LekZ*��q�������cT���"�@J�ֈ�X���R�Ubj�EQr�[t��,r�֪* �DT\n6D��ܥq��ZZ�Qq��EA"��]f���#F+2�5J*���[&%�˔+���-�%E���Ɋ5iUcneU-.�f�DPPX��Z���UJSN&e1L�qĹGZ��,ƙQF;�$�EJu�G8�yO� ��O���2�C��Pv�_m��@��s:]L㫖SJ��\*K*��\Uj��Աt!J�*�������o2��ub��SKSA6"�	{_lK؞��\aueN�z���O���;���̬����]l�LTj�T2f��>f˽�-��]̭g$}@�o�J�Z�Ǵ'���$�����$};}<�%�<[��E�a�8���Bnvp��r��V�z/&4���i�)�w
^������O'5a�8��&�%����,��b\���B/�7�;�)Z�{a7��ױ�Y��1ջ���8r7Wi�[t��&P�;�"]_$_"��m�W��������e�i�XI
I�8�"G>��^��2ҕ}�7v0�,��y�q�ڹ���l����#�rg��8z		���9�R��7�6�W�B.s��a
���i��x}�^o�߃Ӈ��� �$����3�ч��s�3Ү^-G����4����;�&�P^�0�`̱��(y��0OJ-�~^&��j�K�1�j��]7k��\WHӖsn�#���8lz�H@te�8�k9�������Ϋ�\\�,ksqjT�^�	��9�K��'BT}ױ9uYL	�T�݅c���ɧ�*ұ=�zǾ��a�ǅpJ��z53�v�yok�l�}��H:Ԑ/2��=�aE�]hT�������{����MK�C��+��~-�v]��)�R���/�v΁x<��}������Z���i���K�g@�wJM�1<��/r����:*�W(�s�5�6�χ4�w���c��c����������x����?s�>U��r����Xc��R��Y��G�<�����gDvN<[ʌo\��yp5�TG��t�IFt&��jD\ȡ��u6_E���[w�`%9��vy����)u�V�0�N6�����c�N~|l}�_�9�gy`B��O�Ž��`Mk����<Ш'��j6�cZ8��Uj{%v��@@̹���ۂd���{ph�v�{�i��LX��|-W�����l�qH�3�����*�m��y.�A��;Tj��˵}iR���04��ʼ�ћ-"�� �͙���[f�x"���Z�Ԟ�9C��
�zUu�C�!u|_�A�p<��R,@r��β��� q���h]F0��;5`!�]�֔Qe3��KV�"�78�4w���,�ln���亩E�=�5�g��֦F�\��~�!DK}����1�G�"!hy,��m�P�o(�����=R��J-,���ye���Y�
��&F���nt�w�,˧ݤ��^��4X�K#\��t�*�ͅOq���Iؕ
A3��Bt�@�������-;S�����d#����>C��*:�u��i�p�_�T-����z=U��}jg�F*�d��dQ����ഫM�R�9��A����IO���K۵ze��<ߋ���!=F�AD��I;>0�}ϧO����/�l��1{(�r0��ֳ�ujH0��#l�{J����EJ��@��c�mE�P�5���V�*�MB9۽�~i��L��=����^n�X�9�E	u�B����V�E��i�U�w��c|�wt�>YUU�ffq��M�x�M{�A{�W�g%<ԭ(r�Tv�}��۔J�sRNr&��Gj]my��XWu�8�A9d�iEA��# �/������u�r��\Ǐ:�Xy�)t�D�B?�!��:͠���ͼ���5�����:��c\�Sv���;>��gw��u�q�;�i;�F�+��yzzA�v�vGP+]���ֈJy����x3�E����m������М�V4R��:qث��R��69��|W� �.�k#��e+�S
����0.��P#Bj��uNEV���(�ݭL&+l��9	���*jӢ�j]ɟ^��t=�`��oя��P�y�5r�ڴ� �����iP�^�7f��>(�|x�8U#4iʉ�bp�s�����hNl��4R��8�û�'/�H'$��i�n7�3�$:��S�G��5��cJ�]��,Nm5.�ذ&��l>{|w�Y{��@x�8��x�P���d^kě*&򷁫ghp5��3��:�A��W�9��cs�޹���<���X�}� �|��D"7����)�5@ײ|�;	�n,R�v;ֶ:�YK�N���R�ry���p�(�I��]B��f��$��h�V<gy�q�2=Ǘuj�'�*�Ή���Gϱ0��%���$�%��)��z�L���K=ET's�;Ec�y��!Z��7���4r,��}A��9K�Ă�
���I�S�z0P��
��;���˭�;��*�/b�i��$�"�k_w����Mo��0j�s�I��,�4�i�(*-��cŘ��uz'T��(_w(g�b� ̓u���g��s�h�4]�\�Ҥ���K�@a�D�w�d��i�3�����\6�'�y'��V�m�?{�j;cp7\z���7鍨FӟC�H-�4*
K�|���{��Ymu��*��,Xʼ�c�J3އ9��p��ޕ���`�D��J���g{�'�3yr{�y�5h���6��!��2��(��C�CYU�7U�#VQ9��TV�hر�}ih��0�m�^�F̊�F���9`oֈ��v(�r����nX-��{:�:f�7=��,vLt%��P���24ѱ0�'�*^E�J;{�zVy*wl=�)������᛭U]��a*7F�y�����@= ����ʫw��l��	���T��>/+���>���X��1\��tH���:��O���7�ג�i�[�X�C�`"bK+��T�֖���'��`�KG�����^E�WL�j��]�_�d�ſt�F�\f�^�!�f�>�2zE�񙸘��lG9�/�XjbC<T�:�ol,8p���H�c!ޞ�+<{����W���|W�˩i�5�j�����n��(�ࣜ�������43��M�ȴU�_YIB��Ό����$�k��yݾ��cXy2	ux��Ӂ�Q�0lɐ��)K�h���a/qi{�}��m OK}x��v�x�j���=��Ul�u6s�-�X:W5�3�W<]�R�$.�>�C�nD�F^w>��N.T6O0kD`�>�/��ǟz�+�P��'M�^hsMj���{��\5'(�a��E�9dK��B��=!����3=�3�֮��b����昪�'ppn��6��+��*ȉȶ�b�z\>��0�ǎ���R¡���(���e��>��<t5�+|���x��u����t�NK��IT!�q�^o������+��D�D%@�0Ͳ�0]X;�Ϻ��HPz�eҽ���b�Z��)�����V�!�J��{FaےI������6���ݫ�%�t���7�|��v��=r-դH�/U��?:Z��
�ʙ��)�8�I=���\I�1SI��&��E؂�ܺ�A��.+����9g�$���� NmW+yV�=��b���d�k�X���yZ5}���j���vo�]b�%��kۆuzOO=K|]-�P��g �=�Qj$�j�+ha�Jyn�M��u�u�h+���˪��}Dqc7��-C%��t�jD`�2�σ��S�|qҏ��紏�-[��z�h˛a��'p�U!�u�a��|n3j��zn:�X�
�+ɲ��g�0^?Vݺ@���d�0���eM�:=ܟS�SBJ������Gt�Cq(ꊃ|��ľ��y��;�3%da^�`��ٚ�nl6�)�:��cNZO�Ŏ���cx��J�΋�'�k�̊�g�אۊ�{��Z�ND�gBjɦ�Eʧ��렠��~���5�;Ghӌv�:��E�����c���G�����s�r-9�'3Sor )4���������^�j�:�t����Mh�v����z��@�2�\'AeF�ѯ5=���*��ob�<{��yj[@䅖�zf�l]).:��DϱP�*:_9��56��Ja0���j��_�E��޾<X�W��:И�'_��rvYlz
w�u3����VD��b*�٘%��	)�r˱�J���(��=�=h���ؙ���K1@ڮcf�\�Ks(Q5�P"_�*��a˸��RQ��_��_I���(��rh(ʐQ�9s���4\8�{b�/�Dڋ����`�d_O�g��p6�:E[S�w���ά.$Wf���H���d��be�(�Ȫ��� ��M��Q�0r��t`�$��������[���٨������o/��`q0IKDI:
Po�ǹ�ߏ�پw��t�,��w�R��.g�"�TD�ͻW���6��n�*�N��v�H�H�񋹦��fu/�zۣ��
�I	KN��ӭ$X"k�̾�Ό|:1����3WS�{���q��7J���Xgq0�9=�7�2Y�t���B�.����	�ܻr�g���1è,3�P�z�3�E��&D�_O����j�B����D*�NFa���<ɚ�*�,�ޥ�RuL��sn	X/ְEII�@��\}Jũ�U�u���kۯ��Km��6���6�D�0׋�M9��7T
"�N��0�؎�;�A��+\��(�uyS�u#V]EYAX�뺁�8��9d�iC!��d=_q�ho���EEm�uz�{�6ʛ4%�ӹS��ܑ���]Ϋc�K�Y����\�[��**�.9Όi;���+�0�YB1��ذ���?<��,�t�!S��g��������D����֠U��4w�@xϹy!@�vn��5x��a[�m�iߦ���W�|-��+=�3Xv�_8k5��*1Θ0���F�h�PfȜ��
�(j�ڮ�{~�缉܀��+A�n�����b��{��{zsZ��u�@x�8����xT�˾�ç�w��T1Q�보���3��\��:�2������V�֙Iz�l���]��|���%�j^Bn�^���z�qD)��J�z��M3���W��d�;2�:6(�X��qX���\�qsmsMn�f%��T��c��{��/�Ǫ�m_X�A]�^���p
Y��e��]�䵮���ofo$Z��GG�8�C(��i��Pt{'���7��Q���:q��2���g�1�8���tUX�y!�(d���;���F�b�Nd��j�-�yO�����9�H�b-&�i#�Am"|�L]W��.M�̴�a�}o��=]���*�=[�>tv,��7��E��ʇ�������	4����!S��V���G����{�+�nf�W���߻�F���Dr�N})��Aؑ	P23��V7�;y��R�Gc����;B���Q��9��p�N�a�u���J|R�h��p��!�0a��@�ی&YN��ƨ��$# vi��r��)9}����U@�M�c��7t��<����Lu.a��P#��Cʎ��q�i����Π�]�$��)�T7�[M;9��֫��{�]V�v Y/��Q��^`�#�k�z̻\2fɃ���aT�}���}�˞<��|F�~�}SPTV ҹ��A='d-0�8���V|&���Bbs�3nһ�<��t.K"F{Z˿�w�ҿxG��_�۝�)ws[����Ƒהڪ9��ڊlq6Z�c;��vQ�;%��w��zu�L\w��_G����oH��4�0�u}�+L%�q<�Ziw�WFs��3�����j$GF�J��rH�s�]`����5�^K��!�����<֐\��ad�u�#�#��F�s��}�{t�tIY�Y����yr?w�,��+�t��nF�hL��Q�9r�0�G_�����SA������͝��H��䘩�R�V����ʸ�1p�#��X3,��K����C!><#y�8���\O�r��2�L�v���m)W���� �NW�~ũ;�Ur���<.Q#�ǝpT��4����Z��*
������l=�\E�s��rȗ�Q%E��	
I����K�D����6\L9�c'<���L��Fn|�h��1x��OK���R��8���JZ���:E��	�9rX����s�*���5o׷� ��l��E�'���%��l��;�<04v;�}V�dP���\�V�R���TI�0��V.�J�q��;bڑA{���јqG%1q.C��^lrU6Q$���:�����%tP���X��(�3�%�s�	ӡ7US[�0�z"�f0d��'[��"�uWR|	���5.��v��}FD׭�	�W�]�{�NjLm��sv���:��]xPM*8�X����rz��*�-E{��q�Y�<(0pq&.���q;v�[����IqW,�y��כ_��5҂�rڙ�mv�A]�v_<#y8T����L�/8na���_C"�]LC�Ь��"��+P�l�M�r��:qE�֨���4R�8V�]K�!,�mV���I�M=�H�;�j�����k9^ຑ#���R�;i�4N86dU�ћ�� ̠�z�|��)N��s�:� ����/��;s����,C�x�U����
�Y��]�8��R�,ո:IGn�ְ�-���E����k�xV�����u����R)o!�Lں׆�,"t�uu2�+0�Z��Yt{��lrh:ͼOx��WX�,��358]�'�
\���o*��(�,��c��+�*5��j���[:�v�ĥ�/{���m+xs�m�a�C�S��Y���&��IF���A<�_��I蒀�������T��}|ف�l��nT���Z����R
�3w`]UC.M[{�%a���'f��}e*k���N�fpX���(����Q����a���C��J�\ъ|9U��Ȳ��
��?Z�̕њs�8Ko�S�=MM��]W,�f�I��j���
=�X'x��u��s��Vw���p��Yn�DfGy+�h^�D��l������e���D7��,��@������s%Fw�.����p�'��̌�xc�`f�)�-BR��)+�;�˔r��s�(t��?b�[�\�T�!dF��V�uF�;Q�J���5_^�|��^s����v�8��Gj4��*�H����g�����h�êYY*��4�1 �"����l��fM��a�pJ��ܰ��{��Zz�D����-��n�}���7->��i[}���ܧy`���ԝ��]4ᵜ��H'��� �1�v�ݮ�/%�,ԩ�=f�8F������ଙ0�+pM��U[8ӧ�����4����f��x�H��/yT�`�\�Ŵ��G��y�$|V�͎]Ln�x˗c&TKl;9��j:�q�g,��u��8��k�JM�����U��(�Q���j�O)���W�n��xd*bW"m8&g6H�X��вw��q�&�DK�{խ�X9��c�	�9��s�㿹��@����}w|��{n�6��v�X��2�u!3[S6]���j��,p�,ay�g+\�Ϸ98�;Qo����ϫ6������f�R��%�&����ߟQ��@��;Eo;@I�u�C�x�=���;�MwI���j��nf��b�X�w,_c����8�/
�R��Q'�]�����K���;�{raR
U�\�a�����������'�qĢ*1���PZ�J\q�(�X`�TժkS�eXƹ�C�k)���MP�MYVj�f��T4ᅬZ:L�9���k����-U�Y5�%�\QUjc.J\l��3&EE�*�10(�*�M8V�Z�r����i�)D���۬0ƴS.8WUB�L1���WWYa�ˆ�B�Z�cLʋ�m*+X��R�j�,��RҤQ���e�8�m�b"%.d��r�V��#mS���X��n��Q ��٤�]Lb�"�ՔbE"����[Z��)uV��1AX"8[[��U��ʅb��"������"%��)-���U�Y1Ӛ�r("�M4P�V	����
i*�]ekc�Q�5�Gtj�m�Tb�J.�Y4"(��1��4ʱX���t�X�ʃ���(�a���AL5q��T�fSY����~��gV;�{M1U�V=��YXz�$DZ�4���C�`��!t�ޮ�M��\q[�ˬ�Y�MC �'6T��q�����t��΅��u��>��V��e�fڨ���Ϳ>6��U���y26���k�^�,Qi#'�H��G����o(�y�8��uㄑ57dED�/6�! k]��y5����O3+����˱ՉJ�Ɖ�<�}U��q�1�|GS���ߚUu2\M�MP��^��&��[���«󨃻�!~y9���$B��z�{\���W<M���V
(�y5d�jD\ȡ��q}F36��ik��P���*8�K�gr�Yp���G�lXN~|o��Շ<wWz��DcL����_����|Q~�U��&�5еcѫg��o+Q�Oe��� ̹��VI5���ol��2����Q���mFD`�
�2	�5�b��{(��q�Qx3��f֮K:�֊S�#&gyH�u�&�,mi�r�%��?6)�����$>Y����I#����/}�{pY��BnFz���Ε�y�x߂o��Z�,��N�HI2а,��[�M��0�tЦ)�ޮ�� ѯom�7�q��Р��r$j5q��_��N���n�j�NEeR�"\�}^��hn��~��R��K���V�G;}ڬ�"�aJK�|�KX6fKL�UҖ͝ua�h�a5M�M��e�q����'V9�&�h�t�{v�eu{|�nIG/��7nU�����	Ȏ�(�uC��^�9L|}_�U=�X�M��D�J3�L�O� �%��r
�{�9��#t2�Dȶ�a7�1�&��F7ì�ӱTɢ�"���.��nI|qE(�ʃ=ў�$���U�UZ�C�|�e�[.�xOR䈱����x��W��پw��t�pM��8��h����<S�CM�dF�[v�b�Q`��% Q=E?.�����Dy��Z���N��p��O.��\�s���Ct�Uy;�}bہaM�u�b� �:\������s"�%��w1�gzr�c���u�L�s����ȵ3n��D�jH}�kکT�Pq�f+Lr�4���{.�#u��%wQ~8S�4�IiD�����5�7��,��P�m��~����f�uiهp�nH�C:p�}�� ],Q~�ª�>�"����))�rǲ=]����-��4a��`����0[�d�Z<�Id^����D7U��ّ61F��׮��U�;���x��}��R�ICi�,v`�+#�������u �Ƃmb�Β�D��$l����wt�{xHU������l m��*bRN�]}�l�O-8N(P�\��U���)�N7���s��P��s���)�t-г
,l8� ���s"
�dh�6c,e"A��CFM,Y���4��鉫gڪy@z��E��q�xs
9P�Z�W��?�o�.�|��z��v ��X��A��I�K��,�o=�����ֶ����D*1�Y\�?^#���k�0犹�"/�ƚ��h/��@�@D�ʹí�3NUq�{���{^�����Q����+�N��*)/+�<�h�<��E^P��{'�󰝆��J!��F��僙"E��N�	M�[O��՜�EW��`��T�hL��*�c�w@�E���D���l�S�;�����9��~����MT7�����I	q4
m"|�\.���7�ŝ��*���b���O�B���M�/�ܭ���Y��k}A���Î�
T"G	 �D���;�W��L�U�G*ݰ��n��.��`+!�n'\z��v̛�ڄo�ϡ�8 �FA�SbU�e��K����vfZ����;k�� �C���9Άpp�'n���[8\�T�QX�2�e횚ׅ��I��C-�^ @N>}G���r��v�9��{9꡻1mxSJ�f��̿s���d�&�NU�;�J�Y����m�ei�-��<�ISf���NZ�|�g�	�#�)���%����3:��y�?vEb�!��C+�+"N����oY�;k~=R��%ώ�F�T����Hf{4�W�T�p�!��c�T/s.�ҦQ����fۨ��~�.���zD)�0�Ӹ��߭q�o�*y+C�f�8eJM��b�����X�00��X]Ga�׎�0Wd�;����޻ҒܼwC���08l};�F�6��������Vy�s��xl���ING!��Z�������9��M�E\q���s�D���Ղt4�r�`�
XWS~����"Į�w/ߦ�{�J��}u	eOE���U_ ~��z�>��Ź��rb�t�F���\�.�ɮi!�Q��O�`#x�?uϬ<��� za�<��<�i��Xb�vuJX���{���:2��U�6���oƫ�Ϯ�i��jƨb y��4B)!i��m��$7�L�;p5�;��/b�(�G�c!LC�/Ԥ��c�/��vT��|�����
j�13��mr��"�}�D���*��	
��[�6�;�ч���ǉ;/�0<���fq�p��kI�[z�9��z�c��e�[�Ty��mm�/��/*�L9�R��¢�;6���[��<�ػa���#��H=��Xپ2"��)z�4���Fh�w��z�nQ&mʊ45��h��!���s�f��),�)��G�}�|+�i�1O:fz)|a�x���(���h2>��ղ%P����k�:�&g�vv��
�9�K����G-��qZ��|$�^��2lvm�ǚ#7n�
ź��J.�H�Bu;�V�q*-�btC��A��)@/nv�Z�����	�4��'�I#d@��cW��Dƶ:d0��E�z�H�j�v�w��)�3U9��b�ɍ�%��vE��LEr�0$ C�b�=����N���%�;E'l{�y�7F���`75��$�D�ۊ�E�4+�ӳ\<���f-����[m�������*q<\�!���L����E�D���p*V����[$���$�&���[�#���!�J��K���M�A��Ӗ��s=f,�ѵ�GA��W�s��혆R>f|Ί�Lu�]B�cyݑ~Z�ND�e>�_@��
�(�7c�5�1[dيfY�#gM	�v`Qs#�U��~��!8�����֕
���Zs�Ã:6f�6�cq�M5���cM��+͋�6��[���3��n�+h��Cv����A>>����f�H�'�;�sX�kz�iK$!���%M1�Md1��%9ֻV��֬��X;�ݧ�:u�1��o(yN�ٯB���S�F���a!�ƭ3���]I�%��P
�݂hS\�I��&�1I� �pP�53�u1O���n��a���lZ���q0-����(����;���s�|�)��0(�8Ԍ��r!����<s\靋"��=!]�3��uG� e3uF�KǩYKI��2v�J�X�!7#)�.Ǯc>߂Qig��Y{�	�#W��rx�÷�o���5��D�*!���8��p��$��1�nܫ�6�_���>j�6,��*�Z����\E/|j�4:�T򢼤LB�t��	�/�U����K;@��e���}��G��kJy������4PdW�zJ.��V�����+���������"2�+7�@�$1y���ڥ�=K�"ǂ&KTOQR#`���`?C���z(k��ke�v{�uI*�ţ0�i�rȊu�n)�R��B����8ڋ�E���c)�L��ԛ��ܱ#)�+O��j^��D<0,���Ûp')O��(��T ��չկ��$�k1���!�N�D�]R��|sr��+6{���;#!���f���KD"ܜo��i���Bk��nwۥݥňz<�}�d�aq�����Ŭ2�9�N#w�k
:�8����7��n"�/�e�
�F�2&���8i�[�\\�O�|��K3o�{Cb��ps����t297\a�.�4�f���S6�E�č���k�u���p�j�"�(�x5�F��]��w}��8�p�h�k�(�.���o�{���PP����8ty��\٩s]�[������T�uƤ�0.��h�"����{�]K��x��&y�b���<g�r_�W�Х�a�)NDm�g���7F��5�07���un��[y>��0>�qW���0�K����F��=t8m�{���b/{�dq��r{k$����8U69H|�M�;�]ʎ�	��C��	]}�t]K�\ݓwgp�p�3��$;>}5�I�N���U�Xy�6=�9�k��g�rc��X�{
�k�篷5&�."�[�TW�/����27�s�[�v�9U�fk��{�4��Gj�%�
Tj�T[��1>�fg��L��
Q��4���C'��'a���urɅG�������5�!�tc�]d�0�&�s�_�d�5�қ*�,{�ޞ�Auv��z��\�\���I�X5"F�yÍ���GD���9��{6	�c!�؏f���^
���߭�u��Nט�р�`\��}��j����1uc{�>H��Jkv�,ԃ9�'[.�:��L�r�f�S�Ԯ���y�{ݜ�'��lV��ܫ6j0���3�Ұ�(��,=�Ȏ�T2��(n��qD����<69�o/=؊{UM�o�Ӈeo���Ѣ�}A�~zr����*�$�D����L+�U��R��s��bF���ZAT���+!�n'\z�ݳ&�6�N}(8 �x�v����r����3)� �+ �!�gX�NҌ�9�� YÆ��zpK��Uf�w6���h!=F�		���~�	��f�F���G��lLPs���x��+N��H���sɝ��ު���au%^;^�
u�_�����>oֈ��G��!��ya��i�]�Z�L"���:CI��z}k�܆h�vO�T�����Y=:�jc{���*���2�O�Ԯ(��)�	�i�`ךW9 ����p��$��8��MC͢*+��B�������H��w�V�s�D���	���.�h�q^1�p��S�P��%|T��t^#ؖ����vX�>j�Վe�����駋s��ڌ�;�n�����-��)�]�E%=�M<>���vya�#r&��}�c}�So<|0��^m�N�y]�"{�*�1E��ok{D�w��]t��C.|��a�9��iOh�`�lPΤa�E�39�k:�<�c�M�FZd���zKշEwAN���E%���+�P��R����F����>@���=1!��j17���"薮��NOn����ǫqf4,y�Ȩ�g,�=b��u��х8D�����U��m�O���F�6@�m�F��ح���Du `#tN¿
�q��I#�"|�asiW2o%o�<��� ����Ƭ7MŇN���t_��D��P��zC�d�jf{�<�6{(n����q����❷88�^�"����%���Q�5H�P�J8t�Q�)ʇC�OvG���}�{�Q^�W#��$q��)�k`R͝�9/dX�$��8ɠ�]����B6&;�5�R�Nk[|��\����q!1{@��n$�s���P�Чn�vŵ"^��5�8̧I�v�ܘ���&c��I
P�������cW��# S�"��!(���US��-���Eѿ���)N�#�XIF��E�4HDtB�gb�
ؓyyO}m���m[�L���9f��B6!ͨ�����ָ�&��0R�0�2|�����X�l��Q*�26�87e�}w]�yDMW���3$X��h���YJ�s�C�����[10�b`F�[V>�̺/uC���nQ�6�LW&J��\�Yy��^5AB!x.�k�$�a�h���s���8��-K��ʉv���Y��p�3{��oJr�����g�t����O�	k��ߛ���ls�uI@��ٸ�y٤����ѷ�,⎩R��0�E���	*��P�q5��Ԉ>׆��s:�%�<��P����J��wB��(wUD��U���	���B�$�N�e5D������׶_�ݝ����:�z�΂��eX�~nE���9��m�>��a8�񯣸�ܨ)��L��l7U=&o\#��Θ9}!�N��bՎ�5l���'&*�J{%s,�̿\�s\����1Wp��S�3���M��@Q�G$,�e��J��>C�i2gW��q��wf�y#{w$���9|�`UT۝ ˋ=i���{�ƹaC�]	�W!;��[(%D��|��ʉ���u�ʢ��.	�1H��e9e�t��%E�)��:��$p�3�eo*�\��7�\G��tcqu�UE����\��c��x����-=g��Q��$s��m����������j�TW���huŸ�r\�t
��ڭړ]o"��X=�i[yѺ�0�Ȅ�!����3;[�;��u���2◸w9��20)F(��ɷCtܗ֦��2V�8�]��<����^�pv��EI�NM�ژt\�\�1�`�u%V�ӏv$�nҘ��h�ޗ��L�=0=S5X�;Z���>[y,�U�n��Xyቛ�Dj;���׊�C��(sy���C�Bn���0���Y��KV)�����(����[�""��hr�lYÄt�ut9�p�2��!��no(7/c��Lj��eu-.LK�ku�N������j؃�܎
3!�:�k���M:bg.�D�'b�':�Yj�1i��4:�6�����q6�iUa��U���'�
�T/�	N$Ҩ/s�9bL��*�1�*�>�b���no+���s�rp��J8\�3���,*8e���0����ig��Vj��T��tN��@�c*�]i�W�L�+WZ�cs-ބ�'В܎�EB�%ٽ'l�o��k-�k���&n���WË���[�K.b�ך����)�z^��"<w�E�nWR&��U�ų��a�7(�z���v��v�2�)k� �o��R���9x��ù��s8�<t<֮Ҽ2x����.D�du�wZ^;>�DW]FAXF�1De��_#��S��l-Y.N �Nt�k�h+�Kr]�J��:�;�fX�.2��US�][80�ٺPJ�>-�i��R�n���U^��(�a �Ox�>=����B�}[Ǩ&�ޞ��Ve��ᥐ�MQ
���%��I�T�4�5AC]X˜�Ǚv��=.���V6RAe�}i�[]�������Dm�s(�������+��K�:<'1�X�-�K��|�x�	���PS�:���-`q���c�Q��L�d(���Œqǃ��qٴB�1e��{����
���s�`�ƭo)c[�5�-�w�����'W�/�M.äͼ�l̨�f]�-�Y�{��K���nH�d�Y�D]zs����p3�zT���n:����6����;�.d�%ֻ���r3w�&��6�Rͼ���N�h�ص8��P�tR��d�Vɒa�X���NV^f��ܽ� mv��V��3:��Ù�Ʊ7B��*�����AG6��]t4lYSl�4�;j�K@���y�m��Bn��� rb|�;J�F>����V�s�Ԛ�U�\�c@ݡ�+��*��R�����v"���o��ʔ���&�(q�7E]^ip����.֭8P�-�Ǥ�ۙV~�Չ9oX�O��;�U�gA�7�."���lw=�^,L�E5SRI_5�,V����3|�j��U⤝,�u�8wΆ
`F�==������͵f�Zr�d�.K�=�)��[Cs!��i'n�\����y���O�vf��K�f�+�d�En���̂>T�� �_U��Z���pV
�f�"���X���
��J�VE4�Eu���I�k$X����EPJ�c����6�R,c�J�1Sq*�EY��#�W-լUX,���@a�\4SV�JX8�WV���M6(�u�MunR�1�e�(�-��U�]YPQB�Q1��]�fPED���QV)u�kCCYb�e��E�1�iV�R�h�b* �������c��J�V0]\pE��,b��Eq��0�-*������R�����Q��*�cmD�q(��պ���E[h�ZX������UJ-��U��eh��YX��ET�K�q���rʚM:tT�ŋkU"�KV���i�mb�b1m��L���R�������Kjc�JV��*(���%n8�+m*[R�QA��f[J
�j�Vҹj�2�F�r�X����V��0S���%e"�UJ�TQs(-��el�X,��u��﹅c�n!/��{5]�aiЦu��К�kiD�𳃆G�	=$[S+\ҷ�̊�f<{�:�*��E�;��f��Gq��M+
�ϥ�b�2p�ȯ���)'=\2K�\L�򨴙�a���w�\������4�؛���Q�Ncb� ��$��	A�c��`��e��K'�[}��d)���X�p�3e��5nYN���Q�eG(�z�O˭Pq"���=�w>�jo4_��Z|�KP��(��U'w����<k���x{^���|�����ؘ'�Z��WkZhI������L���.�.8�����ȩ|�P��Βr��=O�wѯ}��S�:�k���Ԇr��A����E�)�NY'IԼT�:�'0\�.��}��l
|���ב��sf���;�+!�ܑ�:,��� �f�F8�]z�n�Y�j%�K��Ȫ�3�b�.�r�>R��ME�o}�ώ�/+ꏛ�U�����!lZ�s���s��Q�
���@�G]Y����(�wx�\S��B��ώ˻s��?V�E����^�݉8�y����u��o�<nn��e�WM� ���:���-"�;t�`���n��:w�!���nVdzv��vߣ����C{\Q�7�ۻ��B�����;�ȍ�ӖD52�.��1��Ş��R�g2z<U�,�Cy�.��Xu�#ި����]Sa٣#svt��%|�I
�2�J؃g�b��D�S��ϱro=��=�:���X�ݗ�x�����n�/b,"��d:�g��C���8B$��p�}n�4�W��EM�옽�{r�f7��HM|�šhv �:灙� ���
P�)�5@�yn��x�ҋl�]N��w�L,�z�&�9��̵
*�.�� ���uD3b���~+cE87�L�Y�5��������W����o�_C=%�8�o��,I�Ix�[H�^�b��~�k'y��^�����7=E�7y�<�Ύ��<E��"�ӕ/�)'w5T(Kfq4Ծ�ۂ�>^���A���#���i���=/�x!>G�;�������♞���\H��aH@Y�:�����9ΆC6l�v�H����U7}y��Cn���\:���$��S�5b�tm���4�r�����Ù��Q	rd.��������f>�cʨ������c~�F�ז��Eo��w�s.c�3`�����e*��T�kB3��=�+tNӾg6�X��~<	ZV�~���zh��O��vos�����S*[�Ѥ���5�����I+kl�uJk�Ud*��t1LK�.N���=��0�s�]2N��&��^��=�w���n(e�遄�:��;���fD����!7�+�ޢ���m��
�ٷz{<�;�6�|�)9`�x4�+�@�	|z��44�:�k���'UI��K�!	�yYc�mR��=e�񖫧��4W��M`&�[�F���lVw9��[��K��%u���5�����2��q{R�\!��mT�Jx�=�c`�Aic���\��@�4OL`:�~1��:EM��@����*��S�Õ ��z�ZНT�;hs�Ztʫ��j��l"�	a,�;>j��l�t"���.�ĩ�\p��۲�q9٢������8y�F�7�n�Xz4�tG�
�wy}52��}|�9�ͳޛ��ˇ(��:n�D#��NY��D����\�P�qWu�_�1=�;�UJ;�n�P[�[�-�d�MJ-�<F#JP�!,%�=�n;���Ө�@�!]��D#�V�U,���K��IU���o����C8�-�Aա���׼/�{
M��y#�_���3µ��[Ws<>��Z	\���`��vZ��oV�Lӊ3UW8e��;���
v'�
�j��*j��b����u1�ZPe��h��>�,۸N%�t�
�[�$�7�~�n&F�i�Ǯ1�EW\���ꓣ�۳f�Z~��KϪE����{ҥ�+@�<n�΅�.�p����Z�Y��+`�,�+�<�0�9$�( 9%�`����DƯc�F)�um���=��95�^��Y�G]�"�DIr�xW�aTV%�2H�C�b�=�h^h��鍃��J���ۗW�� ��h��q�C�Qa;�a��p3�pP�^�)X3�QfL�I�.��jf��V�:��2��<�0JԚ��<.@��([q3��{n��I���L��I޲��F�i��;�S����(ˋ!�{���J��K���MP���僘�uD^ARqZ�o>�b�ͬ��YN��8jaȿT2��YqWX�wd-rK��QFW8��u�ˉ�V&�)��K�t����1���;߳���
ۣi	�k����9����ؓw�$8Gì�4��T�_��܋�s�X!�I!�Ó�X�ʍ��x�����wq�=�a>r�yW�i�˝q�Nh�c���l(Ȍ�v���D��7�cgfB~�އ��Ppy�� .l;V����d�\ZE���n!��}\ӥ���Ԋb���P��C�:�FPZ�8�GHT$V��G��`�=]ǲu��]#\l��b`觘�e:q3�#��[�Q��ݕ�6޷��gP*]��ʹ$�Y���%ogE��O��iZ���O%�/h�C�#�U6�A�z�n���s�v,�#��u�mb��Bƞ���n�L���uDW�d��Uy�TX�sr0S�`��gڔZY��<��*�8��]�<����3vd2FlP��&D�KQF��:y�rJ9�Ciʿ3U}�~×��\��������:��*����TJQb�\%�\	3}<[�p\G�Z͂�C�5˴hl�� �?^wXL��9�1��D�
�x���H!������w</ ]{�����u9 �`Oz�=њ�"�;b^ݨ��6 �b	��{>H���~u�7�8aܣ��_n�1�~�,ʹy˦Y~3e��i�rȊ�p`�P�p$��m
�VQnre$w���r�P�6n�:�*j�n�C�ʠ�g�m��X/֟�hm����w� �Ry�YELI{r�'y��\wC"�n���_��S(�Rn�v�a�6�o�Pv�{V+ՉO5<P>�(����uq�"���&�&e��y#xJ�V1۟[���Y�i�� I��n�/^x�hą����sLַ���������.�Y8�W�x�k�|A�i]綅[8�;V���g1���#����Q�7��[���&�c�Vi��������f�[�&�]7�oDn����&Ǩ���K����G��x�`�8���;|k�� \��{^��φCP]U�\���E!��g715�Yf:�f���4�^}�YnR��B��]�[�Q��6-�s�m�y�Ƴ�L��E?>�B��l�ua�`_��\�M8����aFl8��W^���AΏD���7�b�7�y+ʎ"2(ű�ɑX��8����H|���������i��Z=�v������M����7�^h:���Y�q�2���&E�.�=.S�s>�a7��o�ޜ�47݉{td�&u�������Ed�����|S[�����Bk����m�g_d����9S=Gj��շ�1��]i��������ZDE{*���A�9�2�F��l��\�+>���lr�J��N���:�Y�P����G�3���n���:��`�#��V�鞪V�j�����E��l�M+��E�l(�H��.&�)��>���k�Au?��O:�Lu��C�L��[��qe�ϝ�������S}A���ÎpAI�Ob��vF}���@�+y�$Njԗ���}��ݭq]G:�L.�*Xc����n��)	�h�C��9\�#kb�X���� ����vZ�N2��9���ua� ����f�
My3���Z�MN����k�1>R�q����Y�Xx�-@B��W1�R��{s)�Ns+^�ܴ�!&���4<k��CӶ�Y��=~o�G୻�n��r�����KУ	P�r7@׌.�����bU��Q�C��g8p��r�i,���8W<���,J��p�@�W/�rtH�y�r��91^
����A/+�۴�m�U�5J�vRȌ~=CX.�Y���b���,���1���,�h�M����v���^�㓳7z�o*"��H{yw�fW��A���O9��5 nC4tّ0�'�F���Ւ��|��$�=Mg���YX�;�6�|�(',�4��M�;�	�;!ki�Xi���\Wd@��f3�|&��8xf�<�o��޷�M`&����55Of�'�|�=g��0��¼��N����+�6��x���<`���t�=j��d`Ywu��0������z�%�`=��?c��9N�x	��_5a�Mp��ݖ�/$Z�ap,1��$���[a58pیʐ�a�������c�T��+!�t�����^?M"ۖ�ZW�
�JeZȜʶ7����-c� :_Sn��m��u��� Ź#N��V�֮ǇW��;��N���2����f�܊�FMlKP�*�{t�R�$��λ���.%4ޓdv*q`=J��wx���:�j	#b�@,U��HG�s��x!��{��ыRv
傫����I�:rw���.���ʉ��$�~ȟm���qp��鸷N��s�ӖD�����oU�&�zu�i�5�$q���b�x�J��P[�<bZ�,�	��O�iG<t�x�JCxo&^�N��*�t�IaA����(��US/ۓ'!�]3�9�{"�9%W��q��rw<M;�k����Gw"����#��čD%@�r�]D��5��V�q�S�7tT+M�	���Z��tx���A��J/��K�D�' d�l���h����F`��M�f�=JoGLA��Wf/J�o��,�;�ґ��++� /�#��d�9�G\�m͛Z�P�cv�mC�͈;M�����C7�sj/��P��sZ�g��'� ����H�U�n��x�i�ܸ�K7n^_��Y�T�mR����y)qx�Z�w��`��C�W:�q�p.��q4�J+�bb+��9IŸ6�g���$����^N�4T ��{���UVt�s�8I8L��G�M��V���d̤"��K�:�>��,�0�2�X�1sC(�
K�����&����]�0�bR񹖶�z"hZ�l�]�Z���&���#��e�4��ڳ�dlHs�"mf+sj���{�[u�#dum��]ϭ^%�;`X,�p�½��5^+�&~�#�Y>�lZ�GL�0)��j�e���"�w�ɤ�E̍,�ǰ�XZ�j������̕Ԯ��E<�j5
���-G�zX#����k��܋��/ä8ɠ"=@��V*r�Oے��'k���^rq�����U�)XX�k�z!�8����V8�Y݁���mZ��C�]�z\�wóf���8�˹*�v�=�L����B����yax'������\��1B��U��F�_734�#B��P:T����*�Β���#�����W�a���)�i˜/�ba�Tj�ѷr	Q�c�90�:����ct�0k�Q��:��8u��g`\�c$�{K�y|w�"u'J�*4��B]��g֫�Cp�N�x��q�.�˭�At��u��u��ZC�c�ʉ*	�&��#�P���u�V�ʗ'���R�vf��"+!�s��tf�$H����ڤ����x"d�D� T����K�kg�ٿKIVr�>5�]wdœ�t�D�j�|��ZtS�i�"�4Q���YE,�E�\9�t���0 z��3���A+q��j�ϥ�WӘ�V2�ff�/J�E�����Zg����S��ye7~��f��+e��5�i�R�S]]�ۯe�8�=��uG���y���[��~�N�gFl#����nYN�����E�Y�D/��(���Vvy�}�&�1n6��Q����ui�T�#��(���Iݳ����Et��L�v�J�K�{I��(�� ~ӃȶxR��N��逬Gt2)7\a�,�݋����{A�^pb9�Θ(�7��!�S���WP5��8�x[��<�d������Ӟ�SCV��+p{�,�\$K8 �҈�`�=��:���:P:^׃.��>��W+O��ӆ�|�9�@�&�]B�����`��
O�TM�S�Us�x��������oJ<\-�|���LS�O<��{��9��Q�~��
�&�U�΀d�Y��ϰ��9~c#��x�pt�:v �!�\ٌ�e2f��p*�o���_D��>y�NlnĜ�
s�hj��НFY�L�zF#�N7�|�x���
k�$j��侽�{��,:���b��=��U��x`s��`�%�+O��ԡ�V-0f���A�w�g�v��$��B���B�� IKH@��B����$��H@��B���$�	'� IO��$ I?�	!I�B���B����$��$�	'��$ I?�	!I��IO�H@�XB��B���(+$�k0  �@3��B,�������0����ꊢ����ʪUD��[��� VCT�$U%��ͨ�R��ER�Ų	K���H^�*,���(�n���*i�i��f��F
0�mk��)U0��n՚�����縯3km����KY�jkf&�����6ƵJՍ4�[@U�V�M��kF�j�k&m�Ͼ��U�v�  �
��]���@�u` �kf��к0Z5Kv�(3�� �ufU�5�fڃ� �@=��s �uh[�AU�w f(�ۮ
Q�� �w\��f��Nλ-4� �B�uSv��ݚk v�����΁۸ln0 �n�`�l�)�f�jem���JL� c�K�Xh�j�� �����  )w��  ;�r� )@��� ���ʔ]��Y���*׀oU+mZ���;k�vv6���ڬ��#n�ݖݖ��Z����k��6��v���k����t�[���մ�����3[Q4�m� ���tѻ]�77]թ�a�v;�weB�ۭ�w9ݹ��k[���J��\��v��v�Y��v�������j�f��ki��� ;˯wn�wV����U�ݫ�n�s+k�;���͚�G[�r۬�j�j�n�dE��ŕۮw�IS��ꭇ+���d���̧� w[c�3��ڸk�-�s5]]��۳�q���;]��m�;k���������V���Y�f�p�m&��&Sm���ږf� ��u�ZY��WTm���v�nwlnպ��ҭm]��k��
������L�k��Y�m-�wn��� � 3�[��t���t�1��� V�p v7@jwp����P   �T��@� #@ )�)J�F       ���%RTa0 �2h�L4рA���%TJ �a0 M0�dD�dɒdɩ��S�Q�=@0'���PI��b�Q1h&&�S�d�ɀ&6��T��^\p�|o|"���-�bq���8�b  	�����
�u��� Tw�� �S�
�PX�����#C��Fx�V N� J��BB� 	�#)@�b��^K���j��=|�`��B޸KK?��a��&Tr���*�$�Dg�D�G;ԋR�2�5��������u�,il��2� $���`X*nXдV� �Ǘc*�	�Q��XС!3/�nH�#WiXշ��v A��(�6F&�tq�^��ں��9��S��+TKR�lV�ݽ4,XuS`kq�Zv��z�93]J ���@��B�֘i��2�\�)|tSm��v��VVM0�˺A;;����Ô0& �Z�c��GM�	�`R���7b�Y*Ȍ�j�t�FbT��mf�GH+bT����ի�2�������MXF#YF��L�	�Ǐm�YlY�v�ki:�c6nJ�him]©Қ+FD���.�ͭ[
l�ǈ�����2���2<rj�MꌌϯV�2�*U� �V �ݦ�݀������yp4U �]�Z�&���fJ�&Zb<�呌���x�(B��4�c���oڝa�1
pR��#�1�7v��i��`���H�kN*WFxBFśI˚a�2����Bh�N�L���Y�ۖ��7��u
R1��.�̀<��dȆ���7A�N+�i��m��ѩ�h9�2�@�6�P���C$��e/U�7�4P�0d���JҚ�5}3&�u7GB���cm`cQV�x�U 0@+$�i?���(,�1�[��W�vfɎ��v���8�e�Y����,T�0���g.�������yVa���'HIKCOi��.�dP�+U�c*FcsV�غ[eF-&��a�k\h[��ӑV��g�^#�%���g�7�m����L�M���U��Z�k!�u�ճm%B=�sej�M�SIm�J�{�	J�`2ҐQ��Yj��Mݳ�Ⱥ�6�<�]���/��t��R�[�l���.�IAK5�:�j�|�iӫYl��zi���3	ٗ�Zm,ٕ�/D�e����1Sī���P&��6�%eË�?�㵚�Q� B77��E�8�c���ǹdE�kLa�EL����û)Rhv�t��Zp������ohcRh^�Y��3*���x�׆2r:F�l��$�����/��x*�G��3N:��:9޼Q��ÉUD�d�܃n����XJV�-]EtbLճ$U�iL�n�ScǛ�4�fTj��j��ch��&�ƍdYTU:ƶ��4���p��:�n�V�Z!���u����ig!�6�l�5ClV
�S����^�4$i����ժM;c6�F@�b�,� 
h��4�t����㱴+&}�ybb�����L��F�!R�PXT쪙tr��`ѵr��U�ҥL �K�B��Vi5,���i0ă ә{R�"��vq�!ǐ-�-_�8��YB���%n|3D4��#����)����u���Y�M�p�/ZG]mB�9q|���Z�v����>SiXi-[�y.6���
��]��	�t۳+v]���Q{�G#B�/N���vbܠ՗���؏�,ll��=K0�a��0�WJ� �t���(���86܋H1�	ô��^JD�Xue��"���t�Z�R�:�+���cS^-j��ht�J�Qd	+
�xowH:Z�lK�u|�A5�(Ы"Q1���[[J�,�f���2,��j�kn]����Z�n�hI���,T4�rj|���j������i�wFl�TrhU����-\v&�u�8����+y�Qv��'$�m⧠�H� �7.�Y.�*�Ê`�/d]L� i��
��)`[�m���V��)qq�W�e#�B��2�n���Q��W�,e���)���ۉ&�	b�4V��Lm��E&��!��Kz�e���XTYc�ܻJ��E�{Y-��-�d�M��)Y�:n���B\T@S[U�+$�ު��q�aL�z]^�\F:	=&�ɐ�Cf�5�+=�r��}gZ�r-����Q�Mk��ŭm��řR���Z�)���'F����^M�]jY��GPX���`�;5\y{�����kb�*�2�nK��"���D�Be�PZ��T�]ؔp�4en0 �u2�5J��yl�̖��wjy˧m���b7�B	z/(�0�4$e;Ͳ�Í����r+�۸��ҫ�nrTeJ��J{�	�3\v�NH��nf�k(2�ڴ�7��7��o&P.eeٷ bKEKa�"���q�J�jDҹHٷI�1*�LH-��aǩ�j����Œ�҆c���q&kB[r")uz�����f�pa
fJ���cH4���v�!�/����霑�员�<O	�ל����k���+o���F�Ir! �C��8��5ۣ9jWƛD�z~h�.�7��S�m���P'@Ve=͵���C�Sn��0ųD�lX�[q�ۃkF��e<ǒ��b�)4]���.���ʢ�#Q��b�U�l�0�)l/7d�D�*�$>sV�f�!B��*���+L��6�+.��X2���̍*y�\�������&�X�h��l�n-����S�sv�;��.SЅ\w�P���[w&���ͫa%GiՖ��"�<9�72[��ô6KǍ�G@���n]�n��M�0���%�� �
��qӱm����F����֭�K�C.��ȑ�ף&�n��+)���s -�̵�RW#͚ZOu�$���d��X*�ܲ��F�t�j$XʱLI7��*��$��hҊg����˃NȯLn�i��e�R�sr;xi�O���#��V��%]����̧���1Җ�\���L��S.|��ݶ"��JI��A�-ԔM+W�Y�����,=��ŧ6Q�8.dDPb��j*ж�̍F�g	�Ƙ%N��ͼ8+r2,�`[$�tV5�\�2�]Bd�Qմ3t�M��!b�(e�R5j�i,AZ7�x\:�ʳ횘�Z��Ed !w� ��a�u��A��@�]��+0�Y��DƲ����Ьa�!��,Ŧ+�����P�p#�ZH��2�kZxN�0����]1x�;jcƲ�d,�ȍ�S$�7C��D�Ǧ�Yb<�Ӧ����۴�l��+�6)�JD3.��c�i
q��Z�r�Ѻ��]��GUa�ZۮX�5���7ŢXB�M���!ҫ��T�=j�݂T���r�X6;rT�{���a���a��1�lǯF�-T���D�NsB��Oh��J�*��C��=z���l�si��dXhЫ�md���h�=He��M��)r�ݶW���E�Nk�a<n4��MX�{j�"����I�qǚ�D����(f���
G�a�&�����8/Y�K�q1+xQ�v��8�]�H�<S�i_o&�.�b�n5l�V�E&��X�]��	�@��}׹jՠUrXk�O��Vr	�9`�fEh�K�X+��iUl��=OI�w��^�c&�e�a#*b��ۼݧU������
FV w6�l�A��tު�&����gvF��T暉XfZdM��H��0����F���^����+�Ez�M
<��vϵ��G;�
N���5^�,m�J�3��{P�$,��n���FT.�;F �mB�A�^��F�ѕ��g@8F]�J"6��o׭H��*�낲Q4��b�Mba�-jY`ޫ��S�2���d�hMM9�T��9���,-�t[�CB�Q(��4�T���ڻ�+a�j`X*Tn��R݅�,A.�X�u�7�X��l����P��w�q� H%[�W3o-�35���*��,�^�=�JOq&v�V�;tlEb1�jn�VM��m=k�`;�a�B|R�.[���x%^e(�k ��#p�4�sXp[�˥Sdk~hPvCSU�˸˽�Q�_�l�ˈ��'lb6�ڎ�"m��\���hh[�4���4N[�Owf"���c8ʼ��aY-d�QS�U���V�!�@n��F��v���4� ��YI3N��P�E|ܴ��𕲵��(eB�{��x(R���u�̫�7���`�3n�Id]nC�̧Y>�;�`Ӎ��d0�-�(����0Ԋ�̼�%j3b���e[H:���X���˧����Y��t��$Z���>%�R���Ċ��� �)S�2�0sZJ�b�jȵ��]d��IAHW-Ӫ��gB��C�qTqD2r�i`�t�ڮ��<��+9��	����lY��4�ʗ$D�K%���`N$���*3N^R.�7��
�`['�ر�?�gU�:�gnR��M���B��#��ɡ����꿷"� ˉ��4kU�[�U(n�bV�s,��q���2�k����uS�A��*I27+
�.��@\l�Vt��:�RXM�OI�
��YP�F�i���¬�u+)�b�-j%�;�%���MI�w���nh��G�ӽ��j	�h�AR"�����ۘ4@V�ͧ���UDe���4n�ۨD՚i�:��e�y5�D٥�]�
Hǈ �Pa�]��7{�m�vRű�9����X��(;4B�eњ^
��۲b��i�Uf�+Y���jǍJ�wF*�BMBnj'I�UFB�Z��ҥ+5�h{xC�=�2�R�L���Vf?U�.:?QUW���߻�E���])b(��������wFe]��NFiL�AIJ��׎��E�-�P��A��ie꼾��d�;��I�B^�⾮c��[��om��)�_fK����"��_]�L�g[��X�c���E�����*P��:ٙ��4�]�x����k�%�˃iޝca�0���]�:��T푧�+�a��B�ɒ����h��C��a�Xb�=iY=m��Fr՜��J��3�-���7�xY�1�v�5����o2�TR�X%qͩD�w:�N;`�1-k�i�r9�mh|��Z���a�	����Iw�]'��5�#�ҙ���.�*e`���u�eD�=�3vq����k��>����@Ȼ�G2��,��z�Li��s�t�Zj�`�dִ��	���^�U����|����֮fY�?dݧ/c��d5/z,��A)���Z���@T����
��ȣr���0��]�p��2�<
b�5/\�,N�T �$��R��g���usr�m�W7b��\t�m �����|��+A�(b#Q2�x�n�Φ�y�1��wQ{-ݸJ����7b�
\���X��2��Fg �Ν-,��3U*Ҙ��w���
� �6ʓ{�Bc��wy��v:��طsFޛT��8��Z�K&w>�Q&�θ:�T�;��\听V���\4�E�g~[�&�`��#�9�Ξ����5�]U� ���� G-�U�ƯqW}�Cw�9�(�)���G�a՜�,�ݜi��"e��1��;���äԵm�6@�a\!��M�*�Z��Kc����$w�^ᖅ�3����`���� ����GA0�{J���@ţGr�9���y��Hb3r,����~�B�V��S�Vh}���u������U�%��{���-�f��b�����#f��Ks�m`+���Q��qE�\_*Y����7>r�/fM��u��N�Y�Ͱ��'�[��e�����(КuJ�Eu�*���+v�
N�
B�>I]���|Lmet�V����մ�(SLf_ euY���L�S
ae����D�j�X$����>�����C(������9�i�#�Vg��{+�[W:����+/�q�o]�t��7��v��aQ���83���T�W3V��}�����B6$���QN��@��;O|��0����p����y;�g���F�`��m���[1��C:��k7`|%�t���y�6�]Վ��X�uf6f����/pP�dvt(C	)!G����em]�ݻ皴�=e1]¦���Q�̋XI���Ҝ�"K�+k��52es&ؽ���.'�j9i5[΋惎��ȹF�м|�O
<�����	�N�Vq�f��嬌�_wDr��J��sr6�N瓁J���9�R1�$�j���K�W}�Tɢl�ݥ�O!�k��y�Vr�6���'h�YC�D��#.��2�e>��=}Q��*SN��x�o�q\����g�.
B򳙻Kj�������iI�=�O{�
��AY}V��M|��1�����kyp��"3�z~Tz�D�sMؼlQ�rӒ���i��+w�@�We��.�Yq{;����Zsc����bv��]__g/��}a�)�\t���,.���K��]&r��z$� ۈ`�At]��LV�y� u���F�a4��@E�:���k�����M�[ى�i��	�ݷR�׫V*c��LD��*_!W|���&��+ؽ�����w�i��y���YT.�"�Jt�[��9!�Z��΢�W��v%Z��W1�5���]�q2�Mjy�
�*���]X��-���[[ص��;9�v�����S��W{bJ�(�)V[�]���*Z���A(���k��D��y��Mb3��eq�^ɫ$�t���d�,]Y
>Όڭ�М���)n�n�S���$�ܙ\ݶ�e�D�E{�fG�'o5S�K��i�7j(���z$�v����bx������V�ܙ�O�.��3uC%�Y}���}B�]���v8*pUêu���A6ܷk&�Yٶ-�|4Q+�:�ۛBE0�-�2�,�
�zu(g6.�����K J1oi��;�M���D�-֏�\���DY��B�ȱb�s\�z��-�/��F�)�^g����WoS�3k��;n����m*�7�+�܁��rI	�Z�LG���gu=�w��`lǶ��C�&E�xHV+�ĳ9w,qá&��v��j�a��J�
ڶ��*�v�c��x�I��5�n�nZ�)��Y�X��%��Xכ2���-]䝰*6I��71�m��D/[�����\��Ն��?Gvθ9�%�����j����Z�Z�um��wӎ�����r��_	;Th��P���X�k���d�z�+��WQ6�(�,8�Ba�!GՂXDU���33J%�l�5�e!m�?>�ļc)�������-l�P�R�H�ڻ���	�A:�{\8���&7��u�=
�tIYٛa��X��X�/	�97�J���lRqF�6�c�.wi�C����ۇk��f;�$ ,]�YYv,�yl��b_a�@L��qA�n�[ƦA�\D�۳V;!��p����9�t�nñA���#}t�@b����&����Ǯ�g{iP�������J���Tz��st3W�҈����4y�+cp�bV��7�st�SZ�n=� n�����`y�b˺��l�q�ܑ,�G;
����T�F/ot����m���\�N�.���DW-�9�Jm�c!HA�\W��5|3ZS7��<ޗ��*&�1���=���Y�U��q䩕�lńr�l�y��8������2pܳZbO;YJ*J͸?V����\KXL�}�Z�x(6�Q���z���(Wr�:d�θS\���p��6F��Eu�2f6N y���R�7P��i�e+؉[	�}O���B��m�T�en\U0�a"QZoNl���n����K`���&��9(����Ѯ���/{R� ��%R��F�q�w/-ܙ�1���v�ئ�!p�F��O�������xU��ݑcݶ��FF�N���ɘ����C��(�Dl$�
΄n�1H����>�}ʵ�����݌k�����r.��d��t��R֥L�]�t�ű��9*�o.�������ʵ��4��A߄J�Z8#-�;Z��NY��պ)_B#uԍ�-��u�;Ǜ-�{[�@).� �tbۏ�K�w�zL5�66�bpt����Oz��]d�Kf3[����]�-l�Tyc9]��v�\��D���J�bӕ�έU/yV[��9j</A�.S�U�Ü��M��g]
�P�2ہ�\%8� �7�b�=��Yjr�{��T���mX��(NH��b˕5�i������������d�:F��RG-n&��فQ����u357p�G��2E݇��	�y�})�
��M���WM��2sNQ�ȵ�+0 �),;V%���`K5��(�Mn����@�̸h��]�8���/%5�Ν�kf��1��A|��)����^l�����v�Z<so%�N�l�I��4��^�` �.	߭gj�z�sq�pOngAi)��b��i޹/�l�`���PJ�#]�s��+6�����;n3pDl��ۣ1�ϡ�oeһ���Z��| Ң��G$��A�\�k�#�^Co4�ۧk����M���(�3fe�a`�S���Iӭ<Uja�.�.*�X�6�F�o[O[
��jV����,;y�]��,�V��J��VФ��U%ZG/s��`�N�zHVd���u�t^"��0*�vGQ�f��6��itft"�ɏ�e��Tw�5��H�6�__U��lOuu�S�{���8p�rkS;5�N+��t�e][��j�eS(]qs5�"t�A"�mk�/���=���[����Yf������P�Y|��Y��c��&�>�K����e;�-'�V�9���3gV���:+R��[4*eg%���ȵ��%��u�	�tm>k��e���k"��L_&��=�3l�-�%&��\�J�'\�[ל�K\7�|{"սv��f�c��y���C�q��Mo��w��5˸��彞�W4z���R1�r��qzÚpEnG6�GM�g3e���Ø]�K�[��w�+)fl�(�e�]®��3!ge�hȶ�U�r��d�T�D�M�+���$����aݹ�H7]³�H�ޕ!�ࣔ��J)ê]�J�s���7�ryNN�+d���6�$�=Ӧe�W&��ͭ��eImM��;��Jl�7js�nHg���[��s�$��'Q�MfǢ��v�ѱiNBt�bNt��	̰'^n�ʆ�t����-�q݄��c�N�o�|���	W��ɛ.�]R��$eM�X����<�ɪ-�2�_@#�D��,��u��L����&�a���&Ց���:���t�k"6\/yt��� �҆չR�����v� [o\ZQ��uծ�J�[�xmF���.�R`6��n���St��Hme
n�b�t3Rs+oj�r��=�������D�+7��� n�N����mK��Rv;3{�_�������~�~[{���"�jАh�2��	�� oN�Ȣ��	��9�3vgB��KŋڔB]���gLs^�P���m���4�e)�t� �������jY�[�d6x7G.��m7y��n���胷�_mN/s.	��+k�w:����򼦋�w0k˾�'��c�������C�mƀ��a�:v�e-�`�l(!��%��m�
��H�^�(�DoB��Τ�z{P[лM��.f�ߞ�d�*����Ls<����w2�RꙌҭ@����H�\���@Y��w{]%%����w ʵ0ajj�dK%��T0�K��7�s����t�Ԇ��#��Z����(�z������k�=D�Nհ�-e,<b��� ����`:��d�Ю^�pE+]��C|+����$�Ȭ�Hu>/%���R�=]CyK�u�Pi����݆IKwTIgB�M��.�]���xl	�^�+
�K)>� %�m+�}y�c{�G� �R���K�)gLȉ��'A,�Ԗ!g��쮥���������6ۥ�nhv]��szw}%vN�R�v��h:�+��T����wv���Q�lj�
���^�69M��>�]9;q��4��U�^L�@Kbˆ\��u?�]5�m����uvda(�wM�ج���d�!�����A\��oC5
]P�o^c���M� B��дb�2����ӫQ����2�&��Gb2��|"������vГ�S���˩Ӳ��]$��֧<ͼ�J|�3>���3Ab�64��/��3�H+�S)��X-<���|EՊ�b���7v�v����HE1}ZFnQ��n�^��N�P��.�%4���u���+r��X�W
�j��m��g9il�tz5�g�i�w;9*:�V6q�tJ�;zۤh)�BC�]�� �,����0F�U�Fd����RTw�72�]޹�|i+�`�p�Ë[jgj7O/�\����$s���e|:����jLU�&����u�Z6����8�J�>5s���۸��;z����;��6��F�+��z����X������-����`�*>1�T��l�W�V��U��*�5� ݛd�H��"�݅�qګ��J�k�.����\����Uxa���[ZJ����`C�.�B� ���͠X1b��سh��'���:3.lY��iR�9X�8 ���YZSҳS�OG+ʎ�O�=5������f���u�%��8��k4�b)�AҦ�C�s~����A���m����Z:ن�oEr7��5]�u�s����.���P<�ţ�J��
/�b §Y�����̅�{�W{st�����@t�k0T�v����]\n��ʲ��`�Q�e���Ф��[���%]E�؜.gJ˴1r�Շ_j!s�m�q��2G5�fN�s|�(�b�Q�b�[ ^V]܈::p	�|���wxS�|�'���=-=ʀ����K�G�a*(�����30N��n��BTl ���u��E(R����z��P*�S2nF����h�ru�؞K���Ҽ�3S�gFJ������:� �^�i�y�k[5 �O�bjvTceMŒ�7�ТUo x����r��#�s%_C�w�:5/T��N^�S/i�E���w�nt���V������л�F�h�LB�<��+n\WQ�Gs��n_=�(J�3T0��L@\:��X�w	Ț/-]p�T�*�R�P,��L�Y5�R��M��h_�N9�G�M:+0��i�E1��+���X�C��=֌��]�jm��e��s�{ݖ�r;Лk&��c����L�ʝ��9��t#�D�4~5D�_6�s�[��}kL�[�ݪ�}¥�Ht��x�E[e��N�c��JΎ�9K�>����	';���j�C+V��hE�u�n��[ƶD�)3��(��� ,�"�GbQ��_rt�꘩jb���� �Ŭb���Ք_w(� �֦�(��kf�/k/6VB�Ts�]R��wW1�k�+�ʎ��ۥw�3�ф脐2��TM�������J4Խ 6n����YݣlgmDH� ��5)a*��3n��j���B��wf��L>H*2����k7�Ӑ��ٲ<a�K;P@���;L��;25LE���ͩ���t���VC��M:ۧ��S��/Sͧ��_uӡ�I�2��wy>�
'��*\y�k��W:޸�o-P�
��'3���i�0^q��)N�.dﻁ�v�D����^�T�;��P��K���EL\����U�U5F)
�Z637�+"[ث&�րv��¸Ơ}�U�[�YC^���X;��Fi,a��F��:�4��祑y)�%+
kXqeb�Ctd��nm+h\[V�a�)��:�*,qR���l���5R��޷�s�����ݼ�W���)��E4��� G�-9�7D���Vs��5m'n��I[�AKm�X�����D��V�L���n��V}��ݎ&q��QL�Zӳu�K��Iq�Ar��n��Y+0�r�hC�T���1�i���{aM�Gn=�o�A*�4yY-ܕ�\��2vH2�ܶ1�g�sL!����q��J��'[X޹6�4�o%uv鐭sm��څ�B^�u�M-�%ч��*f� wr��yX��_=�M��#)ؙ�\t#,���Z�(�2&��c��<�W��+�k�i��H����wf�Ơ�ꂬ���յ�uwE�)�U�X��˗��t�@�w\[߭cM���ŗE�J�6�ڕ�z^L�IX�� ڕeS	wnJ�
��󔼱)��R�Λ'9YF����m�v;-9Z�Nf�fuh���S�
���֍ޑK�M�S2M��0材���ݸ��3Q��
�\os��l�!��A����v�7a�\��m�E�&�Í�Q808byȸ͝�����ĕ9Q,�����s����>�,;F���V[X��7���Ք�3�V����K7��}��v�>2V�r�g2u��(�f�������ڜ����uS)�m��͍'.s���[w�r�TC���PWv�Cj�d/��V7�lr[U��C�.��]�n>W���"�17ݳ�
�*FJ�rV�Mquէ���I�ӛ�t	���U�ݗ�(��n�g���L.7{HeA��bh����7���z!���:��b��e�R�9�-�2�7�m�'
������pQ{O��f��d��g��oX�Z#j��W���;Y}b�j���5?���a;����Ԧ7b�Zjۡ�2RP����]x�ȶ���IL3�J%>���M�X"J�Q�qh�%�}�'ڝZN��وu�;�
Wt�=�78�����j�&�-���v�r���b6�������{��iw�'7u��j�W���đ�[u$�2�밓�tov�Q��sEj3��:�u>��3%ƛ�]M1hr�{ۂ��@�uK���7�Kw�4乏�JG^eC�ɈU�/��r��)^��L��:dd����O&��z��" �1sBv-�:
��37�P+��/�ʏzb��D�˺Wi!�j)�J��W%�l,��3�5���%1N]��:�M��L`�ڭ���w\��w_(�(�����Ue
�B�hu[�E䩖����lwA���P�G�;����g���)f�"��}h`@�S&F�u��yY1M�� :�u���V:ˡ���Ѕ��F�L����9�dm5v"¸(+�0>�*���j��ܫGЋ�U⡴�L���\��{w�2k·K�\��vƖjy��z旕u�iq�ػ(#}�x���g�Tc�5����^�Ⱥ���5P��.�m��b�ʓ�M�cΙv�p��Loe�워[��}�=�N�<�s�i�i
۫�(0�T��w�)�yA��j�Nw��6#:rAcD��=��^��3����]�|3�Gr�Vc��,�'�C�2�6�m��Ҧ�5�.��W��O�峞�zX}��J슠�CbW�V�f]t����a�BD�6���s.��ֽR0�r��[��S�V^�/{E7�:e��L�Y]x���3���Tr�̘�y�vl�99W�݄��zu8jtW{5Go�,���pR���ۡl+�ũ8���S���4[ 3[+C�׼or�u[���uZ:���+Ӊ�RӗW�8���H�gcuu�f��ˈ���:��_�əYT�uݫ�CIm;��i|͎Iu;[Y�EIW:���-�Ɨm�1{}V��֐HЎg[J%2��/o:aܧ���s�2�*�[̛+:�y�s:H�78�7���@n�Җ�n1�=�3'>�]c��+����ڼ�dN�NJ]�¡=GU�����{RJwe��cxj�ղ�����߃�L43S$wO��(ţ����v�3)/Xa.JJ'w�9�p0̄tݹ�S��8�[����S,ƝWp嫢s�k�h6��@H��iY�����7*	�2���B��7&N�·��<��j��E,Lv�˵N��ˮ�f[:��K��i������e�|��p�4E�}z������~ AR/��&G�(_�:�D���?8}��hdM�Zʳ�tS�O�W+]\&��Gd�Gm����]R��uÎ_H�o"�s'm���M{���(|�<]1ɛ1��Ρ}l�����Nwgw$�+Ю>Ȳ@�c1�O`���B���N�pXu]�p�,;�Bk���&���j`�j'T��P�QWmTw��ݶ)��ݵY����S8��n�SU��XVR5�ǃ�p�Ğ�. c<�#4��VsyAN���[%]���]GTF2k&ru�Ȩ�/���6U�ۓ6����@���Dp> K���XP���)>�z�d�I���;�s��ʲ/E0pRuҪQ�x�<�M�PL���Ds\������V����pÕˁ��J�2K�`��K��K=��_h{�����ar0:+p�G��0�{ǎ%�Nn�y�%�ݭ����w%6��{x�:{o.���[rIF�1MJ�GRQ���Pn��s�(%+;��>t� ڪ���fQDEDd�)X�QD�G���PQSR�F
�6$R��KkN�UY&YDQV޲�J"�Kj�E�+P��UDeQAD�*�TU��F*e��B�U��mj�ph��k`��`���`�Z
,EV�"�F**+*QU����"�RVڨ��#"1AU�*�(�R��1���UQTD@�*��Z�T�AA�mr�h"���"""��"�#����*�b�UU�0��(������D��AJ�H���Z �TUĶ�+(�Q�Q`��h��*�Q�y�5}�{��T�?��k���7�ػ�haF���d17DGY�ѪE8�J��懫�N������|�߱��i{i���4�$B�_j�mMOc��v��,#�e�Id5nj���0ѻԪ���Y:�}��ӑ�-R<K
L���^��́W�s0P�[�2M�eU��)��f�pά�*��'��ц������y6�{֞hm�"�׮Qk&5vI̩��=�qT��)R�u��O5Ƌ���ደ纬Ϸ�Y�Sn�\Kˈ�!�1{�"�]$�i��g)g��В��������:c�8�DWoy@��n�Tl8(͟L�$�J��yʾ[`ʶ���? ��N���n���y���8R�r��OpfNX��7:��4� dT��G�K��:ㅈ����Q�L�|)�rb߯�v�!�m��������~�wI]00C�\����[-�SM�H�;m�16�WP�/�rGl�|���˷���Q玽�f��{h��ڇ�P�2WT��8�2O"�o���b��v��j**P&����B`�q���H�}��ݥ��?M������y��k�'�d`vǍ�/��W|���$�쾼è�C����c_P`ĭ��7T�#�vO.o��mq�q��`�	>vj��))�/�
��<��}��t�gj������H�@��a���R"��e6�]�SѬ�i��s|]���$��Ou]˼6�nLi��9J�/��<�b�V�*���joa��y1ܳk��7z���Y�j�bg�)�+-m*0�}V�G\��#��⻻�MrArK{`�:団R\6i�����I������G��i���_
dN��#�������GF.����U��/UFP�=�挦�%5f����-r𛤯��l�n��\LL�Ӣ��%|��E���b�@N��*�"QS.�gU�@k֐.�ò�����ǢNyҰU�:�U�U���`	Mxr�ϕr�_{�;��+y���[��*����LGw�lF�$��G%]-���[�Qm�rs�ɹG3ժ�uv�e�۽);��M���_�|�x��);{�eޛ3ǂ
�7��Q����
�7o��!�4��P�ͬN���O�Ǌ'����ݯ?�k���W�T絝e����R��{��kg9�;��OM���i�Lt+�ٕ2�jj%���'�=��E�ק�,1�.j:�|�TC�RZ{Yz��%���3���m9�b���z��[N�9B���W����H��}�QO��O�m��~��B2�q���r8��f6��7�jM�zZ;=9q�Q ]:��#��w0�Td�Z�`o=�_���=t� ⥥>`�����E>�;��d �Uz3���oLnTn5m[L'K�'%<�l�T��eTb!I�܆����u����Y�����Rc��{�51Db��F��3	�,Pu];��\�l#n�Bx�V�h��&�=���`L���i��it�Q�ٟ%C7KG���j��� M�5�Bk��i�әq�_^�˝�®�\."[}D	z�}9��@����Y96��B���9�s��U�ssլph(�p���B���측��F�j�c����/K�F> zН��U8A(�Yg^��'4�H�I���qM�m�x`A�&k�N\���4j�a	d��^?8C�������ti\W6�����8��D��}����Z����^N���5��I6R�E�D�����ՀAˡ:�>w�أѓ�G���=E2�җkg�ʺ�<�O-�e��x1Q;��A�Kq��D��9M�%3���g�Kǃ�z��k��eAGS�!�-d��r�F���z:�ո�{��V�"����T�JԤ��!�OǛi��(ں��w������I�ܾ��}�P��J�YTg0�!X�+kkU� D�O��-\�]��>��[�"��$޶*��#k��!=��)�g17�y�#\g`S�Eٔp��B�иJj9���(���Qڇl��cG���HM:ا̗<|d��.�����*����$��N�����`t:=|�طQڷ�5ϸzH'��������Bu}[�Er��$����I���x���U�L-\��5n��c�)H���qZ扷�� ��YEA�&8�ދ��%�t\�r�~�s+cP�ygZ�+�h�ZE�+�ͯ1�
�6��ӕ�1d��b�aU�� ��u�yl4�|�	��?�_>�LVb]+wu��N�Q5�-:s;�S�ӻ%H�t���Qz�\�#�.9Y��[�[֞�S;c�^;�`������ 3wm���ѵz6�>E+�N3E��\i�'�rM^uč����� g2��I�j����ԓ�����kZ��a��k�A�|.2�l��.�=��Ok�Ę�h���q.k�\�/$l!E��r�4��P+Mmc�چ�{vG\�1 ����W��t�&�N�iZ�OG)��ZFSq<�P�ۡR�q֓�V��_�Н��>]�3g�0���z�z��(6��*R�*b��1�5XieU�+O���:���99ek4)\�{(p��޿���̓<O�i�<丬��3֫87����K�H�rȵ[]7^�/{��l�v���(��XS����9����<[�L�kVţdqh���HU�\Jo+�E�c�V��5&\��
fƧ��VX��Z"��ϳr��a����D����ah���§T9J���7��Yї��(��y�2��pm;q�Q*��y�SK�8��ԙ	��^JMU�{k�P�p�k�4�8oub�L��J��۪V�^�&�5w$���:�J��f�NiS��w���k'��V$�,�
��\���w
�gB4�֚�3��m,���U�L�B��p8f�37�U \R��&�܅{�Z-��|��=�s��Q+�:UZ.�[	��G��P/�W���m�ʾ�:68!L����ru���<$PY�a륳`�*�u*Y�@󹮤H�5D�����ı�vl��!p.;wRJyZ�J�L�Oc��
�1��9O\�\�{V�H<y��S�"��Ȓ{�<3	��X���7��y��\���g>�KΓ��ؾ�3���H�~�֌�Ab�$����t�c���
��E�������}u�.4)���ز�sݰթ���r�l�]R��C
�	�WX[���͂+i�:3�I�k�3P�(P�A�uC��
N��������$���9�m���. A�f�	�r�\�k �1��7s�cJ�Qg} �V1v�+��a2ڱL9�'67u�۵��X���΂��ez���N�t�5����tcG)R}�N�X����Z:�Z�c#Fu,ES�b��� ��N��IL�G,�-'�cb4Y��n�p\.=��:�⡕X�sŦ_N[�s��)39=޶v��^1rw+'P����s��@��i-%���
�N��W�!P�B���o�g��By��ep�����kF"�h�٪�K��8�����_��*
:� ��zr�3�,@E�E_k��1Q ��mf�q��BO_n�+w����G���o�x�>B$���x�Yу����ے��ᐙYa��-<p�nC�靔��ݒ���A�%:];����%�c_�j��>븠n�@��R���^���ڱ�6�v��h|�'�%~]2:7�\~�ʯ�}	���x�Wm�����ђK�7n�J�L�2�H������o�(��j���cyr�7R�V�9x��s85R\�v����w��M�{Q�����K��f�3/`�͗k�d��M�K�kPa��T��a-���G���J��Q�[R��q��wB�OZ}v���خ�y5 �Tp�����Y��x`ԭ0r�M�RV��"�Z�8�i�]GCV�q����ڈ`jS�i�z�a���6�\���m)6�L!��t���[Rmd�<��5q\��z��(��9J�oz�.�+S���"QV�#�rp0�r �3TD�����e���ҺN%rn�� �o�e����[�(��.��g@Z3���Xj-%�����s����)��c�����5�h�!cfd��
*ٚ�s�a�&�9��\7�y�Mr󃂆Q�9^�2�<iT�[5��3����݂,UhA B���sJ��4%�ڌ��\T4�47���}���xq'g�[�%9�}bN���ƛ˃�ȱ\$��W�=r�����ߓ����/���^X"-��U�7WfVu.}�\)Pn2����i�G��k}��w6�����i;q��FdT-:�n_E��
Ү�������p�\�36���m������n&2�BS<$�)ZCmX�Գ�-3�E�T�A;��7wڕ��(B�Ԣ{Q����6�yR\̭DW-<��Y����\�ŸN����d����a-���\�tRu̕��r`*W����38�0;��%(:�Ǯ֢��D��|�l�œ6wcR�d�Y�h�s���k4n�C��}fڴ�{E�
�Mն)�%�t0k��v����P.wTE�]�yo�#��c�޲C]��V�A�ֲ�j��{�R��%ܜ���ջ��Q\[��}�4�&��.ٻ��b�Z�'.�wu-O0)����1�Mq��ͽ"9�$�2����y�,d�}�,L~��Gk��?��<�+�*��X�"�1hV��YYE
��V	�J*�V"#&%UQU�DF" ��*���,+*(1b���b"1EL(Y����"��-)X*��h�EVҨ�EQTAb�+�U
�X�bE-�P[kb"Ԩ���YPF
�EEb��TX�F1Qb��1Jڥa�-Qb��V� ��-�)mP�ZQ�R�TQ�F
��j�֭-h��YTQ��+m���AD������m�kR��m��-aDZ�Tb(0T@RAER�T���@icl*#�s:�ys��9�OX���OFK�������Q5��mnº��U��wU���L��'���/��n]���=&��j�k�@B���6�e�p�Vev]k��X����=���> m׷Y���#\O�����[�]Q=��w���s���/�i-�"���3M��d)��U����\��h����v�8�����������q.��z�7�2�xx�jO{��خ��n��hOq�5�]ؒP�8��µ�d�YáBm���H��(�����s���+�vU���=\�:��Ü�ЎүH1m��E�����vS۩D`�J���
�Q#�H��FCE��!:�\S[>�Y�g�VX�~W����E���*�j�kӷhSӣ:;�Lwi<�u��u�����VzK�$����#�Wx�i�O�Hb)Υ�DU�uy��\�Y��ra���9�����Qg� �}�jÑ�M�]���*�<@�%r��<���	�.;ݸ�_6�m�8��r0�o �^߀�+b����WG�/�am�s1��Z��W�oJ�5\�P�̾��mq�#=����Ѹ��=�j��b�f�1v-�g<����:��ˡ4u�~�@�EMH�l����J�oˠ�Jb<8���n�ǃ/^��V�=�e���,*%U�;b3`��+a� w�m���8��@�N���Pv� Ú��դ̥�]�^�5'ws�t=r�	���t�u �']7ps���]7����u�^�˺�`÷�=UN��!�?A0cD��Gu�>N�u/z^���yl�:s�n�S	e��
)m�Hg9/��f�����ޱ5�瞇<�j�I^o-$�K%�����0^\L�v�R��j2��]9�"֭]��Fsf�7=9}U ](�fjӍ�]�Y%oZx�7� �����Y1��
�X�/��JM�g�����<��}]���q~y͠U�u�*J9C����T�>�+��s~�U-�J�	�ǋo^ý��+� ���%"̇xl�\��B䫠���v��s�/��fIY��iq��ںd�
@B��Ɯ�L�9=��Q	�)ڣ�=��c��F�?ߚ�N?����=���g�){�S$��u�(k��o2l��u%�R�8����et��m
�7�v�H�{�"�'9*���������+*]a����`��ݑ��s�r����.\��+���\��gP�]c���e�J�w�����l+�6�y��$����� 䞝DN�ō��s��x��I�O������7ڨ�U��XM�ț�,:o�gM�D8�ݏM�'���񋓹Y�>q�1����D
F��O�iN�Qyp�-b�Z�$95��w��<VsZ1pC�gn�{"�uo2��Y��}��)��9��(�jz,��Mn`'�+���\���B4��j�	;�����ѧyv�����D�PC�u� �����T��Z r�h[��t��9�eEK�P�����W�����w���.�>���������e�¨���Ƕ��Ok��8� ߡ��L]微L��8$R5�^��5Q�/��pl=ȑ��z����y�[�n)+�8	��H=
t��{���H�; ��,��߈��;�����u�����
]��'Ya�G=jz���r���	\�� �)e��SNcq�t+�xm34�Dm0���0c��F���=s�9Ζ:�j>�K���7�� 7��Ďrs���rv1�ʻ"Z���=V�(׭�עp�(3pC[�4���;	�/���mU��K͎Q^���1��3ҵ�y��<��~&]M{ˑ�֭��'���S/�X�����®��Zg��{,�aB��U���&e�n�:w�j���D��*�r�z-�z�țT+S:|q��FE$փ�ftU������R�s�.``�Nq[��������G��5�˻�%�#��4�Y�L�m!y�q������(����s�ʭ�	��&��v�Ll��]�:�)�h!b.Z�szЍT��l蝯�C�28n,���`��>W��"�<����7��{�(ӒEJL�!�[%'��l��Rٰp�=���t�录�l���LO����<�l
�*Rw�ty����f@��|����Ɨ|k�mҽJ�nvib��ǚy9!��{���٣qK�{��d<0�s���n�f��
�H�"4�����V���1[�,�AF�)s�p�L+)�ұә�=@�`�ٳa,�9���q�IV��,G�{�HWJ�eU�F�-���Q3�/��u��,z�����U�T��o>��[䤜@�X�_eyҧ��]RL!f�I����|�/7O1��C�i*��ہ��l9u%����߾K�Fn���迱�ڈ�,�����:a�g"�����^��_���7�I����@�����y�'n�3�VW����I��-�(�}��3�zm�@�l��ރJ�c���q��W{VTj=2��$&x�8�vv�ĭ�5�7�7�=\�k۱+�/!YR��il�#aĞ`�y��z�:�љs���4�IKzz1�#%��$<��-�}1S�̢�Wd�q�q.�N�N��^l��*�r��7l���:���[|��C;0 ��6�]�h�(�9R���F��C�K��t����Wu�*�R�ܑi_lYM�jrn1�r	qy֔�=e
9��=/:N�QQ|rS,��P�����ʘ�(\�tWN�Z����eV���z]@�T-�+ �H\"^,��/v�.{y� �IJf������G>����Iך�9�]o{ⱻ��T�a�>u<��J�0vLa&�Nk�ˊ�%��Q�)'�kr����nYs�ћr�TN��*ͭ�ӭA�h��(�=��yC�m(3r���.����`�z����Ƚ$^B3����ь\I�ˍ@�r����n���7ZC��L��񍼬�)�
�u�st��2����z��ڦh��Y����x��.�k:�_��	���?`�k��,[�]�.��e1y{��il@T��y��Чٴ���{}1��^t}$�cA*��O��9�⵬4C�Fv[�X�2K�q:d�ъ���\�XQ�jz6�+$���Cdԟp����cV_��J:WQ]ϓ[X���=qE�y��\���9�L�F�ȚG�XS�\�e����|g����s.��]�sOB�u��s���)E@H�=�>�zL�N��
i�F���=��uH2;�p��c(R��ؚo)�أ�Z����ܺ&�%`��(�X��e���WW4fV���|~ps�%s̭�q����ʞq:'�����.ؼw�(/b8��&�g���A�Su�����Y�n���4��K������@+�H:��Gzɒ�&q)]�]LMj�N��ڵe�K�U�6݉s����*e�l�.u���e���ѯTS���)YH�G2��u��<�To��ť���)��m�������l�=bj���~R~m?����ﳌr�_1��1{��v������Z�{�M�i�	>�j�,K@�-M*��$W�)�4�W,�I0����Yg�(�x��̓�W��le+m�=*n2����4E�գY�&�zyv�2�A����Ϩ\�U�� ��˾Ao`N5T!c"cj$u��
����.m�"�7�+4�\�cU{(�)��O&{�����p]�%�����-<lU~����u~9����b��-Y~G��1v<춟T�jM��][s5Z��d�xf'Ыq�s(Y�im��9���M�:v���*g3.%��w�L��"�&k\i��.��GsrXs#�Iuj*5�C����%��kz6���~��-��+��J*�fo��0��35 �K�s7�$^7��6�ݚ�a�u��n�ݔ��,Q�i?
-��)�[2B���qe��0et�'��E���۴~8�uYP
v�Z�ޝ���OxD&<�!�1�[��ُrs�f����^r���D:��3��Y/S���G@�so�%��<I�z�_fo.����^�#:�\�]��n�jU1�y٬:ǩ��n�;%��G��)j%�K�4ҲFv=F�j����*'k%�����t��u���l�.L=�NR�T]��k~Y��X{�pcv_c�y��;�B(r��|�M���DT��{Mv#ksv�E����mo�����FE�kx��y��^�Sm^^�X��u;s�G5oH�A}����Ҩy���B=ج�u� ���Pz���3��:�0�6^�}z�WV�Τ��R���֪���n��\FH^E���D�v�Z�*�$a��q}��L�+.�Tg�KX��.���1ᾩe«�
|�݆�t:[L��,Cyc�v!� �|�����u���]�(,���w������Ya5ʝ�Z�f[#���Z�����AD�;E�E=�;Y��h��PV��c��>����Z��7�T�[�	xrN�^�
�� ���G3�,<R�f���z_ӭ!AeN�ˏ����}Gl�����Ky6��tXɸ1v�Q�N3��곜UI�ŧ����a��}����̺�ѻ�%��"
���Pc�#.��r�4�jY���3�W�gA5���"r鹎`�!��q��Rf�3V��^h���$l�:����n�p�צ�m�Nn^��(��W��S��>��I��QEE��J�kH�T���PYm��QT��QE-�1Ub+(�
�UE"�"ł�*ńX�PY����`����(�Q`��X�E���E"�`��(�D�)TT�P�6��0�(("8�����T-�����ŋkX������+D�V0X���
�1��0XT��R��Q`(|H���.�㿉�Ѱ0�wpK?�7P�l���&�퇡�|���rq���4*�$uR]����sۉ�|��=O8��?}�&�q��|V�x�Ag��4f@�Z���/�D��
x�5,�}������z䋗�]�7إ��"�MkQz�)�[R��ãr�)�Dq�x'\����BIO0&jH9�xA�C��
L#t`��s����2C9w���Z�x�"U&vv��Op������e�@�/��L�;����Z<x�����S&t��k7Tm��xVj��F��oiP�ED��ѻ͝���q��5�O"�eq����:�G�Z����`���ð����H���;��soҟ�.;F�;�C�:v=��U��s)�=��z���S/il�-Ύ������(��*�CU�i4Ș�^^���\��mlYy/t��y�ԋh RY��y��q]��"��1�Q B�b`T�kz�*��p���"��x��״���D�ׯ-�U�K*�c\��H6Koc����\ߵv��]�`���D���Lm-,�!�rvx,�o�S��Ad�KM�xj0 �A0X����%�dQ�P�#y�K�rcd�*`��U�uwӤX���ͷm���j�tEJ�U�ʶr���[�w�>�դ�q�ɼ���N5�lP�vr2A��츔&x��7�{�y�JƧ�{���~0�tt�) oH%����nP��O#)��mr�*��^f�|�f<�yy��iIlM0Rћx����5G�8o�c�l�ٶ��r���G���*E}�X%*�6���u��,>�t��S�:=!ũ�Y�!�wz���Dxr{Ŧ#>��ޜ��ۖvTc=#�qd7�2Rǭ��T[�p���5NnDN��۸z�gŹσ:n����F�2ij���Eh;�i�k%;��j	�z�<3Lm^\��@X�Y�'w��+��O.�M�[�hE�!�No7F�l��M�R��Wb�_&�e�OD��М��}y��n�)z,�>�4t�Ʊ]�V��%�Vf�Ǡ�����^۝w�o~����vE���o���5��!�����ܶEIy�&^O�9i@KISq>l���pK^Y����h{�[�9�:���GZ��룹��W,��\ts�Aը|�1���j�l3s\�:8���j�k��K�� 7w��)Y��XN�N���j��%/�����)'c����sz'}���]�tk�NV�6���r+��\��2�ïg���i�@�k�{Û]�R3�F\��n�i�XfZ�!�s�6on��!�����G9�r3"�.�I�V���D�WUa�ᨸ�`R!��N�/��Ъ�N{��;�ح�Ώ�U��:�*ڊ�+��m�@j�q[gG{���+���c_Tb����Se&��z�,]S:�GM���[�*����՚[a$�O����^�Fr�B��U��Ҟ�D��&��^�p�Y3�kd�jTd_�0����V�.��k.b���M�f�MɁb�/����չ_..S��!�vō��Xvw2,��h����R�z3nJ�')/�B������6"�[�H �Q:AԾ�{���z�w��R����OMr�'iԃ�
�B��{����~�W���4����2&6�G_�c��j�V��a�^��+G�4��xnC�=��y�R.��a�{I���3�<:(9[; �9�v]�;Q���_\�n�����P�}M�Q��ֵ"�q�+(�s�E���W�oK�-���C�_s(�����m\P�8�A��Yu٢Դ�uF�;'�G����2�΍�\�gQ<k�cS����I�;�)�s�NB1BC��W&����W���IVo]Ѳ���d�\���޺���16빭���%��|�AF�rV���1�޲j�]�FXp=4�ݴ�3�)�/r��(��`RMOq5��c�M�J*�5#Qy۠���DG�}��x���XF84��md�o*E���=8�fw{SNz��\��艋��}ih�=�l�����"Eܴ��_VotzF۸�u�u�]���;��6�1�h�xv������V�A�[u�٠7���l3�_s�����M*z�\0riw']^�"�GHoP<3ѥ��V�OT�+�WsO#\JۗS�Q<���#q�Y|1:���Ug4�i�ZS�=�"���C�L�]�c�b���F�6\7Q��:��B������u!Á��2�`R�D�*b�V���)VA�]	Y�*2�:>~FwWsnW{VV���n��Q��k�Pbx޽��q$��+F�k�ɳK���
�k�^'��¦��wFfs���i�"J���X�wQK�z=�^�[*O�>{SRp�I�1�JQf��{���>�y�}pu��:��Tަ|U��Y��v�ߎb�<�w�O��z:��Q
�g�	%�-9Iܡ�Ze�yw�8�m���I^����8�چ&�
U�C5���~��a��<È,�
G<�[Zn���l@*�L�9����m�M�%:�m���u��QQ�#��>��x��,\j�֒�����A�Z�|^�N�1�ֳ�{�:9�]q���!�|V�Z1�ӹ��9�$�x�ہP�ޣ����f�g&9^��r�h�i)�<�%����L�}]u�r��j�^�� �{��)J�3hI�\AV(N�8hQ�/��iN��];vi{�Va��Hu���(/�=�;<�-�j�����c�����hiPr�Z�4�	�[�9�o^�w�A��r��u�����ʽ{�-Q]$�P��5���j��(7Hu�^vE%~�"T�Q]�[SY���uĊR����ڞ���AD�wK5\���K�B�#1^]�E�9n{S�B��R1�r�ki�����֌�C�>w/����Hu{܊y���]�ÃN�q��#2+�tI�V���W��$k��#<�Y
$r��H��s"��S3�<�� ���۸�v��\�P�aAx�j����N~/|bz��\���
&����}�[:�Յ�v�);y�엫(�x�ƶ��O�Y�K9�[����j��NM���.� /5���]x��g/��\�&�YA~{�����Ŕ�3vv�7E�=x��`"�i�6"���6�)�c[	��X�����-y�
��i�Z��{��;�Hc���P��R�kΣ�d��B��>L�aG�ɝ��rkͫ��n��
9�SL�����#SѰ�&�zyt,o2R�P��X�\)j�BǷbGVr�*)^��M�mw�-�8T^��BV�Q���S=.^h�A����s���Lo(���ݜ���E�n�����bAto�G'�Pn�@ټ3x�I��Z/�'�Nf�j�<O�s�|��I��0ٞ��J��㵍���պԀ��\�����=(��UB0�u���Z��J8N��7�^��MWQ!�FWZ�1W���A�u�����	�og�ޏG�����D��B�l��g�.^]vhl3I9�e&ZR��T%�99!r��D*lY:�3&z��h��V�X�(ao#�J����$8v�s�����toʌ����{|���l!,� x�m^�)΋��u�s���'���˒�H xtfj��XS�7u������@��RzHy�����3���7�$m��F��|�>�^*���	l|���co+$<���ǣ�tC��0�6�9��G=�B1�of�a�N����^da��A�!����i|�TG��.qqU�`�����s�=��ݹ36��o&�U����FW��<�I>r��.�����J �	N6�\ȶ��B��:�[ۗ���ԩm�q�hF�gr����4�͗7E�h��Xp��5��H��`#��ll��Ǚf;�ezM��uyq�y�6��M�;!�!����]�4J͢�y��Y[jĩG)��������</��s4�.�c0զw�w�v��+V�w�&511��\[�pJ!������.�X֏4�7$n���u����������eZ˾#h_]s�=��eJ��~�%�.��g�m�˫�u�Rie�}X;^|��U�Ƶ��G�"��2X��eL_8��������1n�2�����Z�	S���avu�����8�\yHu
��ަ��u�u�����)�D�3�Ju�;�W�Hځpq:��뤵���3���I>W%`��!��Y�Y�|m�B<c��iҬ뽷�Uǜ

�7N�P�#1ud�i����37G����Ӄ�I~=R��}Bxj#Ok�^�d��ն:�t�q��q�+7rq�l����R}��Z,ĩ\��y�������Ʋ҄����;>�b��R��{IH��rq���8erk������-4R�2,���j��pn( ɍn)ԯ��W�|VN�}�:�u�t�yԢ�+�h��%��W���{�6ԇrXG-P�{�Y���;.�ovgu.�j�)3wK-2xe�_M���q<��5�.�Gn�n�AD����;�geκ��y�1B#s[�� ���;/�H����8�xP�;B�ٖ8D& �s#����o@X�[��x�V�rZp��tz8�v��ꐻ��^c�*Z]^����7c(��yz�^e%�bm�&�!��rvCj�Ԛ؃׼"�Ǽ�}{n�|ц�)Pӻw����r��.:K��f�nv���������ǋ6�.��k��8�r͋j,�O�'=�W�@�X-m���`�}�eaRdEVc*D`,X,Z£�%���PD1��cQEE�!�-b�d+Q�#�1Z�U�PX�F
����"�E �Z��ԬX(
9VUH+�T�(���DQLk"�UC2�*�����AT��PD�em`�+��e���"(���Qm�#�T��2�e����X�q*�"5�Ur�G-b�����Ό���^�u��7�79���FNq��`=4#��FEGnG9�C����=�������"\�E6y���Lf��ծ3�#���k)!�G'��v'�x�w\Z�:Z�FG�
r3�)5�u�9�Ы'_� V�����eL7�T�꛷��	�UFS�\��������(��Վع�`5���:Sݰ�M{b�A7 ӡ�Ȥ����	!W,��]r��[��A�e'����p��EXG�����	�Ee����V�M�M�S�X�����[�Ṕ7�� �E:��D�hטH ���3�U��d�N�
�7���-1�=�ϝ�rM��2JA��=I�w��L�*$��Lǈ��tt.��W���l��]��PL��:�	�F���jA���M�ZݡpU��e:�&��&hOn�E~{ޏG�&�֛y+��_:�1��#��1����ݰs�*m6V��YE��w-\�8�&��Ṧr�l�|P	�c����W+��9��+Z����ۈ���p\�������1^�Y˛i�sO���KD[�գZ-l��zLTO���]Ώm�[Ae������.Þ�6z���_s�@ �D9ַ���9n��'$dq���5�Y���R�QZ�}��ŕ�/�(��C4��$J��N�۱U�&�u�Y�Y��f�OF�CY��I��';F�)��ȋ�f*A�\�9�OK���{�6nm�z��޽��$/��+(PV�.Gy
���d�'].���J
��S�ھ��L}F�(�
X4ijص�J�5��t�T�[͹��';��_�F`�W��b���G��CId��3�o�Υ)�9,y��x�� wn{ݗ���%�*A��:�T#��={���k���ˋj{�
q�SQ�aR��V�"�V�j_p,�w/��o��Y;W���6�޹Jm'�=כ�>&�����;���{�)`J���'s�B)��8$�݈�7T-�o7�Y�xՂ�����h|)p܂�^h��tW5����,�7�xe���z��j�L��&v��m_�C`��ݲ�7�����^�������]��4[-�Ӣ��ZE�i���aHX������f��td��c1W�R�D�(����|���X�����#v�á�v�ğ,J�n�W�軫�V�{��$R:�eaWݎ�����q���yZ��Fk8 �ޏDG�>��w����B��x�h1��$�K&��GBM����7��Dr`�����<4�ktKÁo��8u���s���2U-�F�N��o/s�2]�dIt��`�
=|��1��/C ��۲"yæ
�`񞸉"�/:��ukrx�'��Y��F���a+)�Ȑ���/�=�Ф������>�����n|�,��]o7��u� ��\���PM�k�te�f+�]iڅ3f�> 2�։�3a�j�l�UX���2�� �"*��zn�`��8�;�����U,z�?��:�/��τQ�Uvڝ�lD��r�f���yYՌ�<&�	�S��5��SI���.�V���{i�}�<z�*��'(����F�)}�z=趰��E~��1��T������@�hz��'�ɻ!�&�u�i$�)Ğ��u�$�=dR|�x���ލ(��߻w5�}ꘇ>��}
����ݲOXq<�Ɉwa��v�q�4��4�6����ROY4�P���t�����;L�y�=����C�{�d:2ϐ� ���M0:;�q8�猓I��I��C��!Ğ?!���O~��M s�u��z����߼�rO��:y� �E2M!~������ ���6ɤ��'��r�XS�$����@�O0�t<��}{������$9���	��`,��P���E2�쀤�� ��i�l�x���&��t>I6�w������~��߾����M���P&�x���ÿrt�:��q
�z΋@=I�Œx�_X
Iݲi'�w-�L�2q5w|�Q׺˓����ѵUG�f#r��!���Ԭ4�~;�l��0�$��CI>IձB[�>q�h���{�5�{�k���m&��9I8��i�P�d3�a6�����t�WLa�r�l�i�ShC�P�
�P�Cs3����^�;���W���{�W�q�I�VM���q�<v�e���q��OY
�oϲI�m�YI��Sl����u�:�]{���aXT���̞2;�$�d�ORM�}Y8���:�R�O!;<��H}d��S�B�~�B���¹��Oj̖*m��h�v{��*hh�K̂��x�,V�ʻ�}�S�;w�_����zԋ���v�ib�7JU�L�U��mf�Oe �]®�R���Fx�h)Z��z"#��v���o��6�1���8�Y������2z���i��ה�i��$�'vm�T��Ht�Cl��;���z����{�w�;Bs�I�Xb@ϽÌ��	���d�4���(�;o��L
��&��'I�ٶ ���6Q�3��λ�����:I8uzC����N�|�S�E&��՚d��}O�+�	�퀤��'V���x�g2He��q��=�~6u߼�5�^z���$�gg(I>a���&0���!�&����;I1�^SL�$Ϸ�*N�wl!�y�u����y�9Ϸ�߹	�C�P�2N�Hx��ӌ����Ld��a���	��v�̇l�0�)ē�=�O�.��D�ku|���0���>�Ű�$�:﬒l��0�Ձ�`u�|�I�����>v���4���h� q���fr��u���k�v��v����x��v��ݰ� �����e����X|��'�4���$�:���&���o<�]|��￷�w��$��R@��\�;B�i+	�Ѫ��hm�m��ChJɦ�����;I=d�_;�~w��9���u�w�C�i'��>d�!זm���?!�HzoXq����V�hM��'E��@�� ,&�����}Q��/&� /��y�x˘����>�ͯI8�Z��O~�;�6�q��q�s�c|ÈVC�P�C�O��z�}����;S�Z����;N������:`�{"��?]���;R=&�&����([r�w�v��I���}��j����IQ���:�?q��ԙ�;�������%��G���)������l�d���L�I���{BL:���I�;��m	�l�Ԩy��'iY�����4s�5����\��~���Xx��lRN$���2Nw:�>d��r�O�v��	�'�P��@�,��N��(d�ɶI�����>;����k_w��B�4�Xj��Yl�哎$�u�'̞�=a�v��e���a6ÿlY�!�[���u_\�޽׻�:�%C��N��Y>`,�G�8°>�����i����8�i;꓌���@8��Hm���}w��\�[�Z�[� s���:�q��,��0�d�d=`,�=$�,�=H�����$�O;��`;��zr���޹��d�*s�Cl&���̝r���C'�a�aRO���&�+	���d��=��&=�[Q���B�ϲ�N���_�a�=��YӉ��lL�ē<�3l��8�m����������i�J�	���%d��ϳ����{��}�ܟ0:I�|��-���	�;��xΘw@;Ci��OXi��8�m�����ϩ�l�s7��Ϲ�u��[xc%a8{v�Y;Ցd� ��i���:@<Hx��'�'hm5�Hx�톘>�dӶ]{���u�o^��u�x�N��;t�8yM$����I�N�&�'��P�d<2��tr��0<d�����Y1$����9�k}	x)�������1��|SR�2~z�ѫl���*��H�<��-�����M:mV.����6�R.��d�m��"���J��r�u��ۗ���6���z=��Ģ�?z��>�d������HC��z��x�Iğ8�t�v��)4�5���:�g��!�1�)�A��b�Z�?����G~��������9��4�!�(|ɶM0�l!��=~Bd�V�L'lċ ir�i	u����3���[�rm�����8w�m8��2M'�4��Cg�m��}a��O�g�@��=J�g�&��'�g~Gw�g�����o�CԓHs=�!�ݤ���tr�m��g��L�'hq� |�x��k�4�6ã��&o�:B|��9������s�r�x�ZHxȰ�wϰ��e�$�'�$�&�8���|�uC�ԓHw�$��!�������{�����7����1+!�I4��x� 񓖋$���d��̓��x���&�>O�`q>C�ԁ��{���Z�^���*c!S���T9�q3�q������Ol��=d�XB��'d����'��+��">�{�{�)&0����?{�'�9Շ�O�u������Hq
ɴ�i浆�CL�J�P�� ��/����S�n�}7>��3��W�T��>,��9%t��Ն�&�״���lS�I�,�2z��i��P����H,���J��Om��O�<��|�߻�{�sz����;t�|�ݓI+�G���ٓ�ChOVCL�ꀳl��$��,1�i�_��o������/�9�X�@�%���S�*R9�F\���΄��^�]#�gK7�"���J
g�u1ü2nMP[,����DgZ��	:��<��L���H]t�P�k�}� B��������>d��>0�Y=d|��`~������i�Gt4�VTϬ��y��CL���L��,4�>�ˮ}�o�7���������q%~a>M�VM2,�@���L�M�+'�C����:`u݀v�ӯl$����s\�]sf���θM$�I�O]2LC�|�����X
N�M2M��m!Xv�����L`gT��v��{���W�u��[����C��P� �g):I�M!����M����I�'_]�T�:d�!�d�	��d���o;��{�W�y�y��C�m!�n�I��&2N޼��@�hzɶM�f�6��SI'��yN$����'��"���<�g�����_�Hr��d6�i&�[$�����}������c�TҞx�+94���0��p�9��<]b� !2����UO9y���9�\7� ��g�{�M�i�H�鍩]q&�DT�E6c���*p�)�yo��ސ��^�Y�}X�+M5D?I*�'Ӷ���ݦ����zsM�"VM���U'�#)�]�.��z�E�"Y^dp��k���u��KY�f7˙Ķɖ����z�9�K��\{�ߕW��Cw�oI[�F��1���+�
h��/o��:F��'�ﺕsV�Q�������wwcY�M"�n��(���_�ë�D��3dk2�#Ů�o�E\8�f��8��8���u��B	���S̷YIi$��*z7��Gd��E<վ�X�k�*zH��m��[ݐT,r��2t練t!��z�n4�-.�wC�� M�^lH;+Ϫ�gZO%!.�<���K bWi���4LN�[�	��ݺ�:m��Yzc�\t�z��\��q6�I��N5�u��d.z��&�x r�&���&V]	[���9V;ye�dH��[�Ҥi��� ����R��v��t�4��E�&������+^Wf��G�5�2��ͣ\�6c)j��̹�B@훩����(�L	�wGW|��H?��������[YYk̡���0_3D���xK`�;U�9��Y���r>ƚG���J�-yh����
��M���,kU.��K�&uhV���n0��Z��ۨ��{*sI`R61��.)�oSp��;���٘_+�SA�l��yJ�`]��/��������r���*�:�V�.)��-�6����̬̆�biqGec�!S���x�Ok��f-��廌�U�F,�/6�}գn��ԮV����Z��J�7Pw9j��� ���8�R#�hc��tv)�(D^Q����"�&�q���v�S�\�?E���A gS[7)����,�;.O+��:�h�k��ʡ[C/YM�j�`��C���bRl<b���u����Y/���ڷ�.&6�Ér�n9�7�����Y.C�����Ǻ����jjp�|9>ۘܓ8a����X�y�t7FLP�6Θ��g�Ŏ�;^�R�Դ�����qw���[K�*�����7\�Y�-}a��o��U"�����1�Q��{�yʽ���.5�u���q>h}�7%5m���4���6�![��MI���Hm�n+
�jf�h���"��\)˽�Q�2��'Y5X��X��y]��tm	s-�k�$f yږ�����B�u�<�]�sOH7�S4�F�Q��+����oP�.?���h�V�k��͔֡�GA5(�BC���* ��\�B3��ۡە�'S�T7
�����c	^np�Z�x!fYt�V��]I�y��]CN�8K�1�fJǑS���
��z�f�w
�r�h'O���;�yf%���Bn�.5E�������,���--��B�ĩ#%h���Lh
�,��`�cij��Z���RbB��J���YP����%��(Led�Z�F,�QA)J�T
!B)j�c����UR�VAIF��"�Q��T�S#�Dm�`�)DR���0+d�DF
�VVDJ�CU�VVlYR� �R��T%j��Ę��AL�
����hE>�(�B���[�_t�B�`���8.�Svy*�:�v�:[���9v�Jv2�V�8��!-��z=��	�%�U����ÂU���҃J|X�����<Њl�-�T.V�K1甚�́C�Y��M���G��u�w�+vs+��"\j���E$��
���e+��s>f�P��e���L�S	��,ۂ�t �^߇������@��F���.j�I2"���LĊT�5��TU���8֜�PQ������oye��{��&��@=���u�O��������=j�de���3���Q����@�}�
`����J��;�0!�:ǗZ��V�X5u+iظ�^ "
��Mx/��^�F K�CZ���2*�Lφó+"�@73"��&�>�O�iك5y��Yo�R�t�RJ�Z\l1(A��ćH�iR��V�m��ȍ�ݣf��/��)`Qb[��$���e\n�^�<��v�L�9l��:��[�쉾��ojY�:�o[7-���$>×�猨C�]�k:��,�k8jH~G��Dz�a��S��"�����m˃� �!�˹2.��ϭ�{��C�,F%��{v�)�|U4��W��T�V�nI�X���Q��9pk
XP�7�]tX��[+G��˓��&}½ڪ
���օG�����Vlo�83���;K[�9�@��5�����*#z����h��p��]JVh[.��!�Z*�T���u�d�b������o̓Z+	�i�4z�^�z��.�3Eyy ��]�Q�W���/���
���"/����՗&���:sx+�+��J����;t2�����ᩥ��Ɖ�7��u�  �!��_� >F��R�����#E[��x-���柵��kշp!	J��.���Q������M�kXXr�-]Y�wP6�3�=8�6�R����G3��;y���M$�W}���&��t�vS���\nHi�¨���U�:b�p;�Y��x��'�[�o'��꯾��$�1�_��Ʋ��0T� ��pѣ�9tC����#X������^�����v� � �\)�`\(Yy�h0�d����NL�٫!�Y���F�?�TҨ���[�{� !͌u|�K:�ߧ�=�w�=�KM]nA�0!�ԕ� ���n`�eOF�7���w�p �������|sL�f�˃E0#�
��Sޑl��i�Z6&���������0����ش^h���%��q���raK��]H�B��F*�Z3kU hp�/:�)�˔뎸�V�d�5]
�Nz�T^������=>�׆eA����i��S*�u�H�5[�	%LBg޸8eOaT���ӷ�.O5{'w%c|l|~2( �V��jȮ�uy[�pxdOªl���..ڮ���뺻�g=��X�?�Y���w�`����yU�Zï't'pF�%�*��Y�!Y��I��dVL��2J���#���S��ﾯ��>o� â�P5��)7
g#n�K.�r���{D�ܕ%�`��`�S���U <`�^T4�/�Z8�ɐ�de�w}��qmog�uC�|,�1]���Q����\=�pdu�%��2m��d�t]t������C	@P���n��K/h���~J
C�o�mW\�����@�Q����+�Ev�b��8�+���ucN l��2�Xxpt+Q_(�/.Cw����N�ڼ1�*�3�V3����'�8��|N�#���F��VՁH}�`C܂�A����C��`�껭A^ᥧ=9���iXkG��g�
)����L�5�>�^{���ejȪ�S"Tʧ
�.yU"��;	[�Ƌ�>6����{� %o�:.8�ֱ�E&��cz�0M�ˇ�;��w���B3E����%9ʻs^�xGgIi�ʎ��l���⮥��%�8� ��jE���Y4 ���DJ��-����\M·=t�5��s)+�4k.:shEQ�߯`�����I���1�����E_����T�����db7}��v��&��&+�5&�h�q*�⡩+�
��+���L�,�'�����ҡ�n]?/G�ͫ��}y��ʳ��ޛ�6�}�q1�f��&�̡����&�b��u������o������.��9��0���r�L�NP�v�^Z�MΪF�����~�}^5'����i2!�s�D�O��͊�P�X1S�l->*~�keL=�:���K�rW�@�m ���!�@�z�Uy^8.��*�i���{/Bv�z8�P�vEЯt?m�e+�KdҊ��,���σ�����O�k=�]��2��@G���Z�]uA��(h�����1[����E��3sD�����Z��:�B_k7c�y�tΨi�{*W�*�q�5�Ɛh�z" k�	os�f�}�T����l}b�~>�0��\�}f���	T!����V�?V߰�}fC��n`L�@_C��`����8[�u��U�f���ܬ������"�f�	����9��¾>j�B��6=M�L���:`���e���<��l�<Hz�YJY}r�n�=�z{���m��}h�_Å�
��&A�0@�(
���C��O8����Q`����RE�اƸU��|GͿ�=��h|���{!�G���"�l�𫞾
�Z
�)t��S7vg�M&f���?:�Y	��ꎪ^4���ncf����"�6��`l���/��+�\���/�^��f�caݩI���rzz��Z�J��T��R�N��+Pw�\:�p����G�+o���F�
@�)ezʗG*H[��%��m�du�����+0��Ϋlu������<|v��EM�}*�0+ r�[T�	Y�����Ā#V,�?DDD �0���݆c,\�H��nẇ&Gs���jO�aʞ���(�O�(����Q �
��(����;���da��Zjn�r�$[x�l���&�� ��pe
�� �_�����#O9eL휎M|�nF\5�4������x���,�B��=�0!�H��{Ck���!��*�u�\j��� H�r�p����ǥ����{�P��~��4x{*(#<9��S�� �������y�ɫ����,��W3P!��&��s��U�X�ܒ�/Ƅ�,�lX��]l��4={�U��D1���̬-8盁||��HׅxhgT� �X�I�՞\� ~w�=�L|�W��Vz��4)qp#æ�0�gy�j��<ܼ<�SdGuD�kyK�j*;t��\��Y$׊*�s{g�u:���y����H�m']��Q��*Ek�œ��n��릹����W��� ��YoQ��3/g"i��)ߤ�I��*��>��F#p����^SǪR��5�� .�\�:h}w\��5��f���nys�.����O]r���%�r���{���	5�L�祗tr�R��W>��v�����Yb�����C�{y+E���ww�=�� c6�^
��x]2��ۺ�<��7�S<��t��ot�7�G�ߗe�Q�=�(�F��팿]YV�%OFP��x��O>E)�հ��w���kN�|,�1P5�_�*F �U����4������,K�l�T]g�Ve!�PD�th�q���GW�#��r  E������`�>Sցf�m���;1q�-�Iqq+��5=��M���`�<8}��heyp���N����G|p�:�]X�+A	���
�_	���_��Z��HK��6	��Y=���}��!6$������ٮj�Wm�u�f�.K[[�1I*{��v�Ϣ#ހ�6������NGD�9�]d\��C��+ǃ��T֩P�_�i$�s�3��)5��x|kO���D�N��u��y��*��)���8ʕ]��\+P��u�
a-r�=�p�'�l8q�=F��\�v;�2&Y�w�Ba�a/�՟�Ά=grWB��Є�n�+#]�ߝ��1�mL��J�G��W*w��cku��	���U���҂��W�/
ڜ�Q��!�g=���iN����IY~&���\Ī��8�:�B��`h�]u�U3��w�z{c=x�<�QuqT`���G�륊�5b�(NUou� nul�G����v �]T��:xe�e�5�����p�Z'k''���-7�z�?�Z����<��/?�̬X{k^�c*s���9֯ܭ_�N�&�k]>j�Ӆi�p���1��#D��s�)�!̥���Y`_PuUu�plGLփ�	�օq�Q�7/��C�u$��z(<h�����}�%:N��RB�^�Y�F�����KO���M�~L��)����B�v)��fFFە9�i��|=�r#�U�nN�P}<�B��`R��l��٪��PJg���L��g^��vy��DW������P�W5o�Ptmd)yg����C�On�#�M�_]~W^Ďd U��1�廥�b@�/M�W�ػ���@�qp.5�/3M��r�'0<Hh �2�p�f����+|׽�S�S�����L+k"��3�ip>W�����wW^�iâ�p4�yp�(1����vPWd�M�^Œ/x.2Y�U�u_ά��A��k�K���fuq�^�$�tr�/Y�P��ўU�]�L��
56��U_�[�v���.���`�{���)��Nkɋ)�:Pi�VM�ݵن���q��zk��b� KWb�7K��Z_*�$���5�D����95+���`ݻSLʻ[S��U�t,�����lr�BG|�"�Fʎ�<� �k�ܨƚ�@+�7��� �{L+�L��ci��e�ge\X�U��˙9QCY9-O�0}z�U�X��z�aC:Qt�ء�z<WhNK��j�ƈ]@;dfe)�WZ]R��X��
�=/��W����1��1��D�lV�H�׷�h�2�)c��P�g���'�M���Rʗ�D��;���ԭq�W�]����Ș�F�Z�8��
)�f��c�Gj��ݦ�����Zt�W-yCJ�{¬9Zw �T{++F�Oi`"y٫)��	'7�3�-Շ%K��W+ѻ�͕��Wb�;ړ�����}[v���,�R[1VHf����.���:v���z�X*ؙ��}�*�"f�&��u˓��5�i�٦ŷ)-��$��ͧ�s��25ʍ�KJ jB[�:\]�h�}��J�$^a��rYR�kb����r)-F�K�{�����A+{!Ǐ�QV��;L��t:>O�!�儢`r��Z5�Q(+1�l�3�8��S
F�ˮ��[ӎu�v'%��h�������\ʜ^:q� �`P�ZʺV�8�G�D�T���ȯT��	���ɽN[{v�6���X�㇟T���V�K)sTa�/d�p��ZV��%���ȥ���!��5�2ޑw_l�#h�9�kqU�f�Q#xUB
t�ȸ����e�
��鮇���4=緖��'F
��2�J��%�������f���5��7�d�U���*A�}v�{�D�]4�����619�h��*C�"��K2+8ue��N�ÊUl�FuY9V�wX*�~tD55�t��~��Y�VJ˖�8�[B�PXVLT1����$��,� �*()AI.X
c�8�X
��D�1��Y![l
"� ��RbE�ib�Tk`��X%a*Y1���-1Z�B�P������3�(LIR��2�j�#s���2��H�(�UEPY�(� 1+�Ԙ�H���P\B�R\����La\IZ�}�·~�E,%��.6@]~�+��`Ǝ*��E� ����s�nN���"=�4Kygjm��Jjo��M�VC�_
�����è`�G�vߋ�Ot^��qY3.L�Nt�b��GUXw]U�ہ���wK1\�g�w��1������u��HJǡT&F�>��&�X�t6����gx选ǃ=��J�0HUy�TO���5��C�?7��l�޺�@���QdaL�m�O�cM9�Nt7�m�j**������t��t)�XS�3��κ���,�+�0�^��۞�Y�~�����D��
� ,A��#N^M��l��b��7��Yj�
��W[v�#	X	���7��aK~�R�o+Ke5�����y<�e��U���f��� h�on����~}1��<2������S�0eY���ky8x�ß�b�iw��\���7ރ�J�3����7��'q��&���C\����(�!�ڦ|����^���g[ە��Q-�ƻ�3��)r��8����/�==�v~�́f��/���u��
c�%��bb�!4����(̙Ϳ#zD�T0<�7>�[�O��Mh��+������Fײ�w)�������"�ɪ��P�I�5�\>���ܽ"����@z�C�i*���ݫ�,�L�z0Vq�-����fP�9jqֺ�ȘSD�I��*��b��\=�׽Y�O73g�<{�R	�c�5y� "<.���q����P�48FF���t^���nhʳb;�O]v�5RK��+�^�jPg��}柁�V��h#�Q�c-����\ƪ�/��KJo;(����vp��h��A ����*���]B;��v�JH)pS��i�xf,;3�B�^�AU�<jΨ�֎W��]���O��ֻ�a��g�uk��f�)�Fi4n�v!w�n�s�#���Y��E�W�H�p�n�ƈw�����E��ٳN�E'a]���nM�'a�֏���Ii�6s��0oc�Ka(8�2�v��#J96����Ψqm�}�rr��6��R]l�λ�)��U���h*�����YJb�N���4��k��>��<P,�{0�<x�>������|�Q�G�ݚ���Q?g�� �J�f��*G�O5w�s��P������P?����(����Q>�t;S�x:Y�߳�����گ�W3�D��F2���7�V�ܿy\hx���x�u⥯D���ՕwPWz�R�	�
)
� �ї��겟�� Iﻻ�h�$yQ�����
�%J�q<r���;g��P�m�I��Y�gp�49_��\�ۀ2�tF]d;��}�\�|����tw�Эf��q�ۘ\�����d��t�'e�"��]����\:_IPJ׾]�׽J�h�)�v,r���
�W�E+�-�,5�nm=륓�6�{�L��]�z ���҄#W�g��R�ߑ膂�e4ޔ?�!H��&�Vs���Ы���"�M@V�qs��r{ܣ�v����t#]��S�ۗ��륏W���+7v�����3m
�tU1N|+f&4 �h�5����� ��ys��z��{v$χ{lz��JZ7�&�$���P�m���E�GD��37������j��V�_:����U��Gc.���ƽTe�A�a𩥄��r��keL;�srz��3ڗ��l�x\݁Z}j#>�K*��cX`��e��/>󛦡��
9w2G�r�@Bx�%{�(�z��A��w<5�nff���c~�>��W@O� ` �S
��t���1�I�)K[���6Vu��U멕J��.m70! s( C-����^�b��xs����4b-kUmխ�V_-�L��|���snm]�.r9��B�B���u�A����Z��ɏ����'Bҫ�n�/�p9w�7��ɚ۫�_G���oZ)�=�.��ו+�F�� }-[.�]��(�stġw^�ݞ}���!��Y�g��p/ʉ_y��D��U�7~��3=���d�}f��u�>�5����.�AK�|�]x�_�ְS�=�
"��Y�ٶF����(�*׷U��%L�v�\#/w�XC�nlԷu�6HJY�`��\��+3��lOӺ7�u�G��1������XN�0����GܓY�C�g�ᾨ���ז����ܷ�r�GV+�~ϑp��w�"ݞ�W��t���<91����*b���-�됄;jcix�"���PV.T��]ZU�5����WU����WtKэX@BG���hT]˫<��馊�ye*�x\��:�G�ҫ�ի��R���a���p��Z�@��~廴Xu�(�ܡZYg����Z�˕�\�H�u�{���N䊞::@G�3S[v���?U}�ն�~���xsƻ�_��1����� '���.��;6�wݜ�,Uxwp��Ϯ����<L@��>���d}�Fe��H��/G��p{"{DxT��U3Se�́H4py����Z��S�\���jpY�A��C�~���#��5��*߻���!��Y�a���]��?h��D�V�5U��p�]�~��nY�+OҌj���i�鯍��,�ג���$�du��y!��b� ����W�:h�]R<	7\��|�NOM��w�Ц<(x�i*JYX��+>��<x����ȃ�����P?�l@�@dTUn�g�Vn��k�tیlN�w�T6V�6�J�;��� Z����gVa5_`(軋�t�AU�o�d6f�P@����Ek4�sNzd��R�����\5���AFZu���-*ż�Q6���J��-�����������N��Dur�J^��7-�Z�3Y�>��{֘sW]^��N��KK�{u��a�T����T7��eǔǜ���� ��*�gB'������_�>
�l�E]g*�pu{�qH���Kle��\�=��%�������b�3
��օ~9M�){���3|�*~qt/���^pR��J&�j��k�*&���~49.��9V8z�1{�t����q�
���m�5��/t����#t�ˊˈ�JS�2[�i�pU9�r��$|J>U�yv��r�G����0C�k³J��t�Y��˫�����ԙb�&�0�}[U��p�8ߚ���.'����V�VB :��@��]6w��O�M+Y6���m �R����Uv��| �E`g����H׎�@%�x;ǝOkq� *0a7�LLƼY;��ؖJBT��j�C��_7�GT���jE�V
�T���o�LLy66r���ϧ�w�j�s3�t�!/�=�u���mX��D׀g������ V
Ӿ�~���Y@;�y�%���8ۇ7,�~�5���m"�5��#�%a*$�d���G��c�pW�*��m��h�ۗ�o���xZ�V
'D���4*��zPLӏυS:��;-O^ڦQ��/]\�u'�R����ւ��|V��>�@l��'�%"FL��S��d�'q���:�}4��7.&|2쾐lUc͵�'ͤ}vQ5��Z<6Y�~�jb 2����T��̵�C�YerMd�j�WK��Vْ�ƣ0A���Y:3�lvf�ӊi�|[��)ˣ38+ە��tf����QI�#����sz�hMe��~���H��;�¹ը6υo��Rt�|3�ygE�%�؝7��w���j�(7�&)T5�/I1k ��'ow��0�����{C���I �䩰p�YL�o6��y�v^��ө>�-��G����@m�s��o&2b6��z�]�`P��~=�UVҼp-	84c�I��Ӑ����uM-9���@
�5I�PF&��0�z�$�[[��/*EA �b��l>F0�\�%^�kAeREZ��@uE�4C��]7.�����W{�`x��/l��� �>�]DX@�^5Rձ��P���r!���;�O
<NYg���������ς�G��k��H�d�k���_��)B^�ʇ]9�[��M��I��^���bX�C9�����+�x�k'���=dj���/��K�V���_^�D6��_!E����pP�"BF�����\,LV(���o�b�_O'�C�u�X ��Z^v]d5	�5�
T�~6���S�� 9�hۼ\�2�����k(���k |�r��b�S�zu؛���].U&]��q)���pz4�V}��vP��*Q�����ʜ
9��_{��s;�'E)����R:�����1�=)+�P��͊�����:1�X�N���H��'��چ۴+�ma�C�X�5��m ;�S�Lϼ���� W���ʕ3��J�וx@�/�]�K4}h�����{��>��=d_��>49XP���[Ӡ�fs�s�ά!���g_�Kc���a`5H 8�g* .a�R{�����Y^g���Y��������b�j4`�����]/8�R�DM�r�9g���s��W�k��ഁ^�n���O8����ύ<xA�+�86��b�Y����S�,��F�L6��n	�P�_��#A�{u�~�:���~g�t2�6y��q���3��H�'��z�\�M:�C׸�*�a��{�c�2�fa�0t��;�ɮ��llx�d���N4뎫�]R�%e�mˮ*�U�zm_ʪ�C��۫ث��+V���꽷W�4�'�Bܭ݋��r��R��y���p+M*��Qr���ۋ�t(*��V�;@�c���s���-»�j�1W�[ŗ�A�j�8�]�"�s��&WM{;����:��$�˒���\��F��Fڢ��:u!���k5�re�j�]Èɦ��8��ƞ���kЯ�T#�b��yz���<���jr۫���P�˂�0��% �`�&2�_hbi%A2��Y�w��c<�uh_�R�nC[�ì,���tc-q�6�n2�ٯ�̝��1.J��Qk��3�J	:N9�sk��͚�����Ȁ�I%�q��=�@xM��n�z*�h[���^pz��]XRd���2M�+󝄾��?0R!wR�D�U��v��̝��9�lD�������BJr�{�Kv;o\��"���
�����ޤ�p�����.]+w{����-��Kz���ӓ�e���:Q:Y����n�6�Z:ѱ����u����o%R�B��YR�m�ˊ�|��;p
r�hv�Z,�X\�l��C;�����c�&n*:ӽƍ�I���+e�Y�L���Jw/U`�{�0�S"wiif<�;.�RI����3c�����l�\Mج��=���7�ؙ�~�qj#�P�j��Y+:8vv�1�:�Dq�e]�q�XM���r�cf>\v�:�(a�Ժ�Du�_�.h�h�2X��-�_N�3���	���ǯU�՘��/P���Ua�&�"T���<bvm��Z�AH��巏(*��qf��Eef��U�K�)4�\�k7�L]�k��t��Fs#����n�J>b�>[�SPB��Eԙ���W���H�nc��Ѣ)ⱺŝ����>=rZ�Bu�1�u�p���
��b�� 
�I+1��d���
�0�$�*$*L #�
�@�RT�LB��H���`V�T��mX�5Ĺ`b��1U
���Lpf�B����L�J�-��&e�c�f[�ܩJc3,1��L���EkaZ�Ă+Q��I�.e�\�d�ĭq��S32L@Q�V�+��AB���q����E0�(K��+*(b�5���,Z��%dSm�b��k�U`�1�2��e)^��/�+b��oA3{���4t'ĭ��|\�hӵ��;5���4�+�=GrI&L~]J��p-�ɜ�~�ꙉ|o��|㦏��8y���ByH���`�b�N��|�#A��ut�)dm
�n���9�f.d���{�����ŏ���у��ШH���l�T�X)���,_��~����mD�mwTT�ՂC_� V`�GD�.�R��I��=�4�,׾]��h�K�o��S|��j�<;��oM�{M�cA��/�aU�P�%�|6Z
�|.��yK,U��C�qq;�{�uV�	�*��B3aP��hCL���Y�j7���[�=�����W�ڲ�1V���F������ʹ��%=�31��礢��k=����������V֌%�ߒ����.u��E�re�pd^[���7�Nm��bU��Fye 2��jۮ����yFTD�2�lW��:��v��|u�I�	���|/�G��Q�����ۧ��xŴ�əƏ7ԯ#�����,K;ݺ�z��5�Z�<�#�m�ȧ�U	��WM�AF�f\FĽ농^<��3��Q�z��{M���T>?o^�����Y?(�7�<i���lV�I��If���x:�  :�Pc�S�]6w�<=��Yn����K\W����W1V��ŀrf�`Ttߩ���&�ؓf���ɶ�C/�A���k�D1���ʓ�8W0'fX]Ou,OW�n'j�s��)�7RUr�V~����Uy*T2��+���(���?`��C���Av\�0�`E������&��<�����OH�]��_B���][ j�:��po��F�
�z	��*�yOƠ�m�|S�]	ڝ�Ǘf���8�ɗ&as��8�ƺ��w&��umPn$cam�|{�/6ւ�͛i�o�3��@㻐��V�Vx�����S���u��G�����S;������n�c����4�="��[�ut�M"����v�L����iJ8��=����4���U�4�3�ޙhh}f�(���-إ\�`�$˳nvaM�l����R^��Q��50���.�
�b��2l��W`��3;��Z�;Pe������x@�#���"�xW�1�����OZ�]�
[�F��͕��=̊VP����_6�����v�ϡ���eP{V6���yA����u�Y�(��<��>�r���y4��Ĭ���xOA��7 ��3�Te���aR (}���ǼJk���h節p�P{"�F�ƽz��h�'�I.�S0�]_m��SSٖ=D�B����Ӭ�JصF���KV�&��[�R	��;{�n[CG��#Uӫ4���WH����6��D|���f�~X�3g���{]�����j�4���f��f�-�c�Q�Ƒa�m6e�3й�t���H�}zm�ݩ���Z�z[����V4m��(��;1g>f�H=����8�m��[�/l��%օ�������CW�}9��&�Jo{�H����0��^.�aJY�:�=t���o���)U&��K�Ӊ�S�?���.DB���˃���Z}�'&���c�kz� Xc)�G=W
�yK�.���TԼ�}]��<2�˰��t ��t������<��D��)W�@�����ї*F݉���R�,�ܬb�=,���6`N<]�ȁuu~������q�eT ��U�7�OeLI,�#�}Z`��c����0��`t06��;�t��1�OK��Q´�1~�1�HA�B� =Vl�U}��S��#��F��ʘ����r�i��|@Y��{��O1�������P�[0S���G��lU�miÈ��U�RWˇh���4��<4kb_�~�-��MR�˷�KٞB�*@�n��YR����;cJ��G��"l�qǛ�㎶ǩ������F8��Y𫞾%��[2Z��
K�v��o{�^��E
U^ˢ"8<2�x<e@����y��~��^7y�zt��~��_qо1W5��Պv��x}�D,'X���싺H�{�^O�rky�O	^k른�#�k,����o)��r��8W�F����?^1�+F|�<����j�Y���!�X$ߍ��A�Pe��P��Ha<@������<4��0<��1c���������$4v�Y�ǜ%�:ײ7=Wakծ���b4E��?]XY�i�v���j�i(�-�>&�+:k�vb��p�9U�����G\ET�'k�v���n���#t�J 1�����Zi:a�K�˸�Ư�;K�e�b^����0\W�^N�4zG�8��$_g�k���/0�OSM�(��
.�<��k��+JC�o(��\=�G�ܞ2޴�.�ˤ�xkD�f��ϖp`e����`�f�p�a��s�o6�S۸��㋫]{B�0@�����⍙�n�� �]���GIA��󥧴����x�o��$��~y����wƽE���g���
τG�.�7��z���J�X�$���q�: �� �pp{�W���g��;e����3YP���<j�c�
Ȫ5<X�Ջ=���b��t�C&�$��h���4=��f
�@[�L[�*�#��,��+ k�6L�L�9|O�^0^*��E[���VTy�7)r�W^{۳�3�5����X|RT�f�����`��w�^���044�{�j�_�Ʋ��}���U�0{�W��:��� {��U6�q�I>�m$�lE�I����/ ��Js��jn�r���{<�7��M�l�P��ՊI�e�{Xz�F�k
�vwi�����4c�bS.rR3d�3��$|�H�W��|hej��^  Q��;���H�ꬺ�2����h��
�����s˅\�~����7��a3w^n�ڶ�䚩*�6�TV��5���!G�x	���)��F8��ߗ�Lϕ���_�#�54�B���n���^ؗ�^�B�3U��@���ܳC W���oc�^�j��f�"`�G�i�w[��+�/�Ω����7�o��+���h�l���0B�#"�J�+:�㽷ko`)��H���^�4�<�_##�¹�1�
�O��f#��RF������[��vZՁZ]����u�7|���K�<Ύ�5kKCȈ��{�Hh�r�c���'#՘��]Cf��hɔ����F謗�uz�e��ݹE:����U%����eM�����3:�]��H[G�鎣��Mgm9iĳF^KWK+�vI9��DcVE�LOM*'|Z�@h�f�@�h�2w��j���k�Y���v̬�n_���^È�#8�ʔ���Cf_N�=�6(p�0x;/늹��[E
��2�
M<�`��M���nf����¨�TE[8 �P���4X��L�~��Yc�կ$#�+|L���j�������P��)���������n  S��K�uK!�0M�=�~���$�Q��pAF��ׅ�5]At�]7d �ж(o�Ύ?w���V l���H�1.���@L@��{�R�j��١��L�) )�jЬ����
�$^S�b�ƹ ��$��WLWC���#�Bh�}��U���CHp�9v|g
��e0V�)��`�D����;�j$�f�0��V36ط{TM̤DԚNm�NY,�;�5!�������*����N�ZA�,�ַ��b�p�{6��)٦����򂲗�1�c����uN��=i�3���<=�::��b�h�Ճ�A�'��-�-���Hq�i�p<j8VF���~��0 �������`��ԗ 7pe}
zЦ�eLw�j
^*�]i5�a=ٜti�}zKU�P��H�E1ah�-�.��u�]�uɥ�(�`�اc�q�C�.�3ʈ����^P,<:�pڸw�l�y9��9�����\uy�hYWy������zG�E8qc���{.�-�����_�[g��w~�^l�ݒP�%��*��i���$A_`���>P{���9�{�Ɍͯa�0|+L�>��_���*�R�w�8��R��}�2(-h�1p��D����o%4��o���zp�c�+)����Wl�N�Z�jn���Ծ9�4���cvfN�'*m���V���n(��Q9j�i���z��
������CG֑�=�R����>�Ub7E]]7t��3M���5�`}�p��-t�3�=�v���fK�٧T>�堊�s�����]T�p{�6H��3��t���{J�0����~>*-׆Parm���1q��FY�p�� <�l$Ƹ���+��D��gy���V�ͻ�9�nG]N}�,3Ti�N�D;�W^ރ/vy����WVJ�p�S8<��]:��vx{xVt���Eo\��& <�N9G�A5[���L+����b���e��dW��=	�PBp�
�G��PP��Y�����^��;���x�^T��Vr!a�"�8j���������~ք��qz��_@�V�����;�w�U�(i.75MIm�;S���Ԗ��]�o$��ɥ�2��Κ�!F�h◒�V��f��!'o(i*�}���zr,F�}/�CASN�P��+{.�j�N�3e{̅r�6�s�ted[ʔ%M�J�V,D�B��c��i3k]�{I����VcO�����p=A�y�j�]�F���̃n(%)�u4v!�mb�X`n��%1ρ5{�r��RQ�7G��{LJU�*��&��U���YB�G䬬�M��:��\(�j��wW7u�-G�H���a��m]��t�d�-2�O��\�2ީϡ�FX+��"K��%�n5�N��8cW�q�̦��
{�����|� �|�ص�����J��R�n�뚤���}9���5�ȏ��
�2�*��8������b����F޽O�x���"���6�^-���v��k��I�Qᔥo%!���l{17�=�k�V�� ��7ع��F�(�f��Y������2)窂[ T�j	�h�Z�:oG ���xy�A�.��rLm�q�E-�Zb���
��zb���ީ{����@�z�c��豵:�E^^q�mW^ҭ�TyK�(�ζP�Otw�LM��x���,6M�y�(85H7K4��D��W.PXm���l�I��<}����;)S�|Bz����̈aڙ�*\�����]G ��rCB���N�y+��z�����M�z���i�8:����Z�s;'{���J�ݒ�������e��kW��]M��Gn������t·uPY҆䍙\��RM�ƺ)���}�Gsv�v�c�m�ۼ����S��kav:e<�b�Gq�1Di��Z�l��8�x�l��:K�]{��:m�:#J���6%���.��}ۆ��+#��0����)R�EA��HԹR��7c{Cҷy��_�>�c�������P^'��@���S#�B����6�s1+YX�����b�b
�l�qQ�9J�F-Er�V(Q��-+�(�1���bĭ��1k0r�q�ĸZ1.\R�WE�����%k-m�J-mT��a�1��j�i�����Hбh���S�)J��E�Y�$��B�Ĩ#1�UX�Q���"��Z���q̳h��V��*�E��E!���.%F��QƢj�ۘUC*�J6�PYX�E��V�Z��l�6ڪW)V��(ۉ����Ĉ��*�H�C2�(�dKX�k!��ֈ�j�mm�-3
�Z���Z")���g^:��2/��f�8��ۑ�J�ɳ
�!Y��ʊNч5�K�}������,UHO�`�*|� �c�Sx�VW���s��e&�>�e�x|�,�$�����k���3�;�C� ��/��u`��<�IR�q�k����@�P���vL�!�40�f}j�+���N��D��g���l׾ċ�0��l��BxW���4;/E�|(�#�y,��}��`5�@�~<�����?B��wy:�H������y�����Z��"ӑ�@S�5[u�ޠ�\8�%��w�-S�p]{9\��B��9�k���0`ắU�\��w?x�@|���������k(w�)�ǡ���hߙ��=�[�y4��4�k���WV�c	�ۆIsƣ0A��ϰ����ܝ���n>�k�|jW��z�
�vsGN(m�
5��^�	\׸W��p��H�ոLa���;�����j����Jt�`���$d �+��;��f.�b���3�t0F�^�����������ǆ���V_r�s�OtW�k��߁�k�D3���ɜt�ё��76p`Z���W�K���xW3��Z�S?P8"�������ٍ�r{|��3���ۏ�g:�PQihu��e 0Y�+whi���v����c;!�"�2�*V���/�����І�fy+͘��륻}(R����W��b��w��L5���}oړ���H�� � �>N�^J�T𪞵L�I�Q�l#	�IX�Txˢ*𠪅x�Bz��>��E����P����K���j�[��Z�ma�5�"�p����R~�E~�+y�|X�YP�rr<^u��Ŀ�WL�ܫ�(u��y�� f7eF2�:�noi֮uH�'A*�2�}�f�-��ٌ��w��%�Rxo�,�һ����P�.`��ݑ��I&N�ꗸsM_�xU�EJ�_�UpUH�U���o��ίgf��
L�떄?��`��o (��3����3J/���������O��]A�[��!ã�E.$^*K~�!���f�"��ˬ����3K�wWD��^0i(W
S�����m��T�}P����1Q�Tɭ���ʘ�[k[�
Y���V�w�K�l�=�^<��>�q��B�!w.�fg#:绹���!�m�G+�YLW"��u8�Դ h!Ϸ�z�1���>�=32k�"	-ؘ'B4�R�^;v���F���������
�*zL��9k&̉{Դ@�s	�U]�Fߢ^�V^_B!�tѢ��+.+�@tAáy�0�+վ��m�#��yפK�3�%Y�x/O$�MB�%�]oMIW���`5lV:�h=������r�U�q;��M�8���6-��-��1t[���7-R'c�~����	
E�L���YXhi�kǣ�ը�͏�_�$#�7��2s�"���ַI�_�ɗ�l�~s��k��w��]* ��u�3��Z0��=+h���=V��ma��Ib��a
��4�5��P-;LY� ��nn��H�az�� �ڳ�-^7T7�!��,��2��"�����DT�މ�\� (��^}����s���8�MN%�k��A���zko�S� ֚2m�92���]����+#6��Q�ʹ�V�۵Y����/���)�3W�DVC^ڠ��	��gЁ��V��^[�^��C����ꭻ�<��V�:��f`*�hUn�Kx�*.�ߟ��Bv/Հ>��� ���e�dH�k�Q;�����X�ή-�^��h��x�WXmX��������eG=�%�q�\:L30�s�H�l��9�`3�Ԣ� �0v{޺u3�i�
̏	�^�M�H�� ��if*F UJ���]*�S^�/lU�W�|�4ృ�{ٕ��P�P��0<+���a�7Sה��I�(Y���Ǒ@�����H�)B�,T��3ώ��ݵ�9=�y��p_
���������,v�L/6J�y�~��]�BRu�B_TϷ�ڞ���j�A ��I����q�T7/��^\\�V�	��[\u:�^8^RT�ǜU«c���}I,�~����*Ǆ.�����2�WqUyQ�?EQ�)��k�,����|����E�:N2���Y���<seеl"y��f��8�Sq
����	�C),�]k! x���A-X��$s|�,�w��c��aU�V;H�Xx���hZ�
:����FR�d�Xy{ݙ�Ci����2�W��:�ّ��s���#�ud[��sh�}'1�Ϥ���)'e<��� <��Mr�S���x���~�3�9	Y�L�!�����5����}y��w ��K��wƤw��v���~�c,ר��: �QJ<9���W��Dm�eb!�S.6�����5��٨K���]^5�űt�����t�Y�.�'|j�f7�r�L�
��.v���V$8&�	�y��_�*���\"!�?:)���S���j���Rh�(R�x�=��x+(Ui�P��X{�����y�DǸ�I��ۋE�	��/��R'�DG=P�
���&f���Ȼ��T��y���^9r�)��q������x7�3/�Ϯ'������`Z���.�����V�N��fR4���^�}���N)/E�Q+����f���ʚzC`T�/��2��tt땍FU��yXsQ��z<��o;����\�ij)�v�#��]�%�ɸ���{��Y * �
���6]U�^z�U�P�W{�|8D�NvUw���;.��S ��Q�d�|�*�4���x!C���ǯI٩���^ �!�k���ä`�	[n�+�B�������b��k=��f!���1;�����:���A0L&̔�<%�M���{�Y�Yt�<+��G��׎B1]At�6H���/������h�BةǄ�h(~5g�u.� �thU��ԣM��r{7��[��kĩ@蚵O��^X<0T�Bg�<�G<�^�/b��O4���iGu�F���Ǌ��4B��IB��驾���a��%u1FR�R���a���ʬ��٘�q� �<c'^���֕G�^d<,x<壾�G�V�y�ץ� �<뾽A��t��d�`��n��=Wi*ͥE�p<�t6���Is�<�3o\U��^�Mn�}�
,�Ҷ9���Fn�l��4���9G�,^�ۦ�y��5+MB������y�Z,�ݬC� 'T�����Q�>�^���u+q)����/W%$�Φ8��k����ꉇ)dّ/E�h�t���&��q�m�������[�@�:h�~��9����o��҉y���l���'+��~����S���v���l�g�L7[���&l�����i���c�X��԰"�E��e�o�ʶj)~���=��a5�_[���C��$Af/�1��/p4׳s��xڥF;���,`������S(#�.��B=�e��N�P�=1΁��~��0���hvxJ�z@��m�I�~]���C�n�ޢ��*���Nr�M��4FS��_�p*�/ݴ}5'�{��f<��nIln�d��
�}5�
���RJ�2{�"]A�/E�Z�����KgD�n+������t�F ���o;��`
]�oo�C��	8VjMH���2��{Ƙ��q,�N_���(R�����wh-��Q�6�w�t�h��0��Oy��%�ύ����S�>�����5�zХ������ʼ�x.1�.�[�u�8�͞K�+G�f��W
q���8��� ��`*�_h��F��4������Ҋ��
��)����u�����Җe�^.<������2@��T��52(\C�-�"���uk�o\nH�ͺ���`��2���(e��5�� AP"�u���<�{�zt|k��a�z�9�5��9�8.+�F�z[��пE�G$d�����
��TTW�p��@�A�3 jnx�O{�+�7^G�P�z>r�|6,}�N���ւ^^ĝt����C�*[%
T�r��&�,i�q�櫕��Y.-��V��贌t�n��C�l]>|yOr���Y5���J��P9$}�ˣ��U�Q��_9V+�����}��*���,����O�H��!�0/�T�'fe��p�_��?m�_�̎���n�0�!��֩|3ą���>VlhT��p^7��.����\=��9�`�8+а<@�49,�]m2�o��+X(d�_y����Gl@/���Mr�8��D*��z����g�'G�K�̌��X�D;��*a*��C�}uM.=<�ĭ̿wp7N����V<�٥jT�-♜z����S��7��;G��<"��)j���	���ٖ��&{in��'��˭ӂ��}t�'CmN��0x���Qa���=~Nl
��e�W�4jz�`<M_�b8]�����/���L���}	��6,��۔�v46���Q��ƫ�|�]!�"	U�$0����V�_@[�8,+;�c��5�w$�ܢ]��h��:�`e,�9)055_vr����S�k���d.�Ra>iwn	��&)K=ϵn�E�X@�O����[��pc�t\�Ԉ�y�cZ�3b��#�ʒZM��k���޽��u9!mv歚̨j�b���gb���J��ڦѳ�0jX��D�
��VI.K�(1��-������ח�R�>�p5[�^�U�9�|�F�)8N�8���r@����-�"�1=�f�|}��;P�O�H`�\Nnj��ˮ|b����]�̮�et�Sf�4z�v%%��}�v�I�f�Sz�E{YS���:��¦�q,m�-bW��wS�z��k]ݣ�ʒ������q���ʻb��ie�w��Y�\�F�>Y\�f��hR	�W/3�9�[fJA�)k[�<\�k����)�/7V���y0��[�jc9���W�EO�G�t�&mf���$��77.�+���0�_�F*25S�(�(i�L�X��;8���ڨ�E����v�M�=�m�o[�7��o9�[��=�\]�.>I`�k�|x�Ms����٣���9�5QӤG�������-fA�V 8��C71��l7D�Nmi �X0<�y+_R9m�k
�e
�6�<S�p! )bIab�Kf���Ĝجղ��u��x:�Mc��8%zb����j��C9�ζ��C<R�n(T�}:��W7�T�6�.�I7���M�X9J'wى�����v��s�Ik�W�n.cp�֕fYWH����6[�XwsVE}{�w[q���zoMخ�-��V�7�y���c�q��k�=+H�*@��0���F��,M����L��9�d�6�3M�ooS�d��Y�m��w=��r4�_�X5B�X5`
 �A����+X�jLʎ&[Tm�Z
��\q�1*�ʶ��\�m�AU���*���2V�
%�" �ZL`��E�9�Z-�V�bYR��*2�F���r�.%� ��-KW2�n65�ְ�\+J*�%cm\���32�0�ZT�E.U�*�R�[e,,e�k���2�V,�EB�Z帊+�6�"�S#r�[2���
A`����ȅTc#�-r�"̴��V9�Vb
�)��`��i-�2�F�L��fZ��%%V�}v@&�$�@|���؇���G�"�p
�Q@�{z�]V[p�ݙ�EZ��fv抛O7Z�Y��y��?շ��y�0�+���-
UB��pD5+S��fC�.�L��+s����2"����5��AE���Dg[�����Ne+�D̩q����j�`��
^������9�`=4yo''� z��Wʷ��˫X<�p�E���=Z�.�����d�{;�>V�tU���: !����|�f���x�ƶ�m��4�~����U�l`S�8 �G5YHӲ'�ge]@�ָ�e�6�ګ�.%O\���j�O��f+F����*��j�ww}9��z�~,p���1A�`耧>�YJ�+�(u��.��E�|':z�<iz���[(�K��o��  �Y�*�0W����#��Y�*3^&�:�*�t t�cR�v2,x�N�����W�����QSȎ�P�Bc`����x�ނ��#��:ooe�{"�P�}�>��ݰcu���|7�,�����-������������s;�&Sۦ)��ۭ�v�h ���ᢛWc,+t��K{_�|����j�+��p�4��ud�:<8���<�JH��V
��`L�5�񉌘��U�3d��I���i�5�;���;��>���T&s����uj׍�i��GI�ڇ�2g���^���k��ji�SS *��ozL�u6�V��=�ǽ�B�ŕ�4���Hh��������e�]C	�� U��+ùP�<��yvk���u�4�=�sI���*���k�&fcEpѧ���x}�}0v�����R~M�����~�#WJpXP�e�L����9�k��i�p�"��&��"r�!?7,������{w��a���u���K��-�^B�N�ȢU�M-ě�חA,�V�=L�7�N��
7w�mvj�#��@��q�R�9�d�"�Mö�������5b�]�)P"�i�53�$ ��!r&�3���ӆw�+F�F/��ˤ<,@IT���h�
4��="~mי�ĉ�hn��#�<XB���
��绍9x��s{�K |ǽ���,�
�eT��/��u��T����@uG�����?]d���3��NQU��V��5���ZJ��OfM�L7��:�W��U.��<;��7���=�Re �z�dܞI�X�ǽ�A�4��+k��E�9u�o�p`��e�˝�ӻ�8?�
���>FaT��B�m�͵�{B�0.�v�U�i�,�3!�u[������*D�`�t�~����s�"�Ğܛ��о5b��� ,T��T��5PA�ꮘT�}@׎�DU�.��[j�媍^��:�t��<8���e�v���A������øJw/��g��o��#(��f��5�vAn���B�N��M�Ot����Q.rNk�a��|/�2��("P�&��� �����9��R{����i��0{4����.��pѥz`�N|��o�M�\�\���1S�� �Z �X�un�����s|;��N3��W{H.�\�L�7�:��E��,k)1Vf\���K�<\%����U���J�Ў=��I�>n�&�H�^�\��
�&s�f2n��H�;3-W��� ���mn[x���zyN�l�ǼC>&�s$pd�$}p�����j6Ѻ�����owCt,��YlVx�-���A+�]08�&��Y�gtu�n���y�H���ݹ�h#�
��qAȈS��\C�L9��{�Rf����*����y�����+����`��/��`Ie��V}{O�u�u������J�	�Eu�7V�5���n�7�MIC8O����������sSr��_6y�dou�T�}��'����)Rϻ�^���S>��
�qq���:�T>��߷��_yu� "��<�TJ������{�2�;b�[�K#�قiå/
Ϯ�d�`�&��p �炥�K�{��%�w\���.uS�a�'P��]Uԅe��~�yΫ|����]2�1^���Y�/F������J[A�J�q;�h������-N}H��."�lˬ0]3]1[�h2�~��jM�#��4v��/{�
����zj�� NL�B��~�bƆ ����
F����}J^�WPC*����mH׾G�N���Μ<H
�о%��e�mo��>�B0g`�ijΗ�W7
�5yA������[G&ij��΃)}�I}�76w�vTx���JBې���m�!�s�oX�Yک��J7ʱ�3[���[�+5��Q��I�N�<ۚ�Q��ٔ�j�#�o��S�h+�!��7�F�jx���
�.�^�@�o�ˠӷ�s��	��	v7<�|X�CO��� (�����o.e���^��I�x��ſ*1W��X�ǃk�ׅ�5]A����t������#@
��S��bc֎�:��G@�:.����Y�{ܵ�&}��PT'��3;���Q�����swG&P�<�C�|S	1x_U�7�9��D�m��L�����0�������e��R�^�XG2�N�\e���/]�₞��Xz�}����5 ��ct7�+W31�uR���< l0=�!�|C��fF��Vu�ڡV�l�ۡS
�j�b!�d���b���G%Jt�u���|��n�
�^�B�x֋wf�f�G��u�S�|�7���2�a�1�Ɛq��_%&�����'D���D��u%(!�ca)fj��j<�Xg]'�)Y�\LH*�{9��VZ�N�օX�:����~*b�@(�a�焍����4�Խ��J�7 �3��V.�s�4�M9ܸ��=fV���T �\��V��]�o+
$�V�*`����4��9-zo<U�fG9��eK��FD&M���b�&����1���m��(���&�:3nEAq��uvR��6���q}k��2�΅8#v5��q��pֲ�&5a|�/ڪ9%�Ky�j�*9ț׵�^�.���q�D�k[�kg7���#�w�������Eg(s,ߩv=HcJ�yvs:[��/T�Ϸ2��kk�N#�
�3o1m�V$���n(�f������iTg�I0YN�ohi`�� S���q��~��n�nCz+f���zH���\���ȥ/ϕ�+�܎�&uN�*|�In3V�r�Y�$Ԉ��)5�����Z�A+�]���~�\z]��,B���k��݊^N��ӭds��r-Ӿ6G��r6���פ7���+!^�Q�]�}F[�.]z�SN��K<�ۉTë�����Lt5ӑ��U�t��9�QL�"њRl�"-�k�iؒ2Pi�����Ԓ]׍���nF��U�ca�~m�݇5��|��rZeX���]b�±�0G����Z�
y�b}bln�Wm.��yR�3�7
��xS��0��뚐�z�*��M�nv�,v�L&���vj�����j�f��23=]�Z%~o�n�|�|~�ކ�m�`A;�����W_a6u�}�.�\%�2��U�U'&7n�v2=�����E����U�w�;�K	�$����M[��ҷ*x���q���-\=�ӻ��.�bj��!H��x*�H�A�uM����z����d\2�2g	��M�0�S�7�h2�v'd�SѮ|�����!{W-�U�}�)�:�,�f�&Ȏ*ڰ�V����.m_l&TJ�$=��W�r�DFSC}}qfgc�F�P���(������1�*��L-X��jQ��X�sb��W����7�Gb�������[�n��[��GI��t�v��+�.����
IS���Y8듷�g�	�=Q1��6�w{K�="��ܚovY��O�ŭ��s��N�d6�"Gq) ���w�J�A�����s��r�WnH�6�1L��T�63�uļ,cg�N���G���,n�h�T�{��B�#5�wC-�u�o]��$�`�5�j�^�y0��P�nBF͟�v�iSqW��>]^\�K<�<�VkD���3;Y��1d=��"�Gw�����k��O�WPG�-���zì�66�k-#U4�|I��/��zC����qC�k衜�霉�ߊ����L���ΜUe��+>�Z����)�]���:hBt���4��=[��Ob�.wr4�;�|���滹Ig6!�t�.�}Ք�RչJ�FM���[��u[ͧ���4ZtVs{�EjC_uĤ=�ٻ�{/�Hж���^�5��۹��p�P�|�E**����ݹ}u6Э�؃.�;|��$�����%�Rv��J�
�ʜ���(�ΰ�pԜ�WV����P̇k1�R��\�X��G6iϚ`��}ԫ9�餇,���IR����ݝh�#�[\e�;��7�Ի�+����*1����G�p!*�"G~J��
&j#s�;�٩�Z#wڭ��Yð8���N��*������Onh$^�b�S}���v�,�2Eĭs�u! �ʹEѾa.�ڱ��M�ھ#���e�@������&�vv�)���Ufb�����N�U �����ϓ�mU��zN��'��2�O:�X��H`�3�#ޚ��m�Ů=�qm�Н[���0��u~�t5�����E�|>�s���-u*�0�__e�)�ZZ�&p��iQC]��Tol<#Jt�.��.9L�K��
���A%��us��� :����5�������Z��b;��
����*)E�rq��]��M�����B�}o�y&#�=���v��)
��3�����l�;��:oK[Z��˒qԥ���w���T�fbS"�[��x.�j��!�6�tܩ\��+U��N���=Xv���im��m���R/���R��mLF_oa(՗o�{t���+�T^^� j�]ښ��N��*�EU�v��vpWp�Af4��(X�+���(�+�dWyb��w\��t�%�{�O%�^ݭ�4z��ܛG�ґ�y	������u˙�vۮak�1�ygX��[3F}τG+�I˝N\x��>�(���z�t��[��dj����y��v��ګli��2�*�be��ѩ�Yp*��-U�����-()bP�T�$U��Ԣ�����r�رeeb�1b"��QR6څDb�*�AG-DUT���QQUV
,Q���bUE�PF1�����X(�%`����B�""��UX���2����I�V*���Eb�1"��(�QSc-�*"����$UEX�"*,UTEEb�AA���EEQUPDDH�UD\�AX��,kX�bT�lTU��Q1�*�,AG�(
�O�E��o�@�w�8������ke���#�=*nӧw&��j�4'�u"��j$��?����R/�ĝ�/Y���j�����)�7��s�]��@�b�\lͥK{�O�9bFDO�H`�o��#J�P�7d��6ˬÞ�ڞ�"6'�)�*�������Ah���YZ�vv�1�MIj{����僓d�[�&��{6Fb8vL������k�E��q�[F�D�*`�J�^ݖٛ<XN�HT�N޳};ۤ
詀w5��@����)���7;�ŹwNm'A��[�ӥji"��}r��w�n��И� ��D.��e�����r�UǗ8\ʏ���QW�V�}�
�O�����{E�N��]�x5�#��㍒eZ�Q���+^l<�}�����|gH��S7x\��Kq��T:��r`T��b���b��[t7d���_Ch�ob�"����4�\^��}ɧCU��u���()����.9ܷI�ȥD:���scUG$����ݐ6�n]g.n����;թ.`����2������ͫ���Jb���y϶],�����{��8j���NHN�D.[��S����j�6F�k&'W\��<W��Z�Z	� �o,o��	�]]�S�����&��>�_`	�P�)�{�|���hLU�u�[+�y�x_eb��U^ŀXo�4Qw=�bFv�.˥����}���V������.��&Ղ�5�2"�����t�g�.y���kqѬ�������E?n�C�d�^������P��*�mz����踯4�v����,�8���U��J�"�ά�Z��,d���N:�D=�%ٮdE��zL�%êo&�j��
9���v�c#�r�C�UDJ�;�b�tb�e�|���G�f���UC��={Z;��w{ɥ�Rx����p�T&;��8�5�J<�n���Ⴊ.ե\!�H�GjL:��HkM�K��S����}t���'��w�r����/mF�]	A�� PwZ2������ [�4�f�������+��r�J�T����.�*�����Y���X�����;O���]rh�א�
��_5�Va�\ؐ�֬�ɵy�(5�e�ޒܘ;x)0�iJ��)������ω��U%��	{�v��e�Ye��v��*e�X��>�f����,&�,�m{T�HظA,�1�� �z��lvdM��Y���"�_\2�:��H�3$[{b�w&�;�iMGuzc�7ہݥ�g�x�@�������îfts9�rza�{�Im�\Wru���1C�]����Ǭ���R_�Wƺ*�@�A�����9nQ��K�ɧ[n���^�4�m0��B�<i���r����5:.����Q�'�NV�d~��<7��j=.�4��f��rc'
�44��z�Yم(���I�swpD�����:ډT��r�#S i� �L������Sz�stN��-�Wd��
�)�U���9N��8}\º�U�J�q�Y���f)��oE�ؼ~{�H�I����i_���^�ܠgB\�zq��*.�Z5u\c)���\8�zv�W��'���I�����{��ٕ�i�{@	�s�d%��c�X��I�cN�p�yy�SnֿD����r�y�s��|�Sc��(Xr�"y�:������=�N*^�Ol���[��ɍ����\�E7�N%���e�u�"��ruN��LmRZ{�;Ypd���i�+\i/�Q���i��n�r�6�߽��gb�t��)�.�7�!y}vZ)%e�942�}],S/̙^os�ZỈm�.��9�腮Y���n��ʴ�F4_���U�b��KN�p[����-��F��|ﺕs@Vѯ4�ELm��|E��Y�t\Q�3��vl"�h*�8��j$�W��"���v��.�{MF���>���T|���戞�L����EG��� ;�Y.�
�]�:{z��S���r��.���/+d���A5�Z�Y�<Q~��9�{�+�`=�4��`fkd��W���s�:�vWi��ñ#Bo�nˌݺ�8o�Y~�\��:m�T�����Š�Ҭ���wS�d'Y���5%��fN���5F�4����Fo���$���8\e@.���Ѧ�eL�^�%�J�u���Y8��RN�����"b<œ��d��Xz�U��f�ʳ�\��\M��f�򾫭�D7Q��zF3;��u�@R�ܙɭ�}\ۙErR9���y^f���)!U9\R앱ܮ]EU��Ywɖ/
׮a��`�Cށ<��%���"��x���;KkTꞶ�⵽�U�$�NEzx�!cx��+��Y
y30��y|1�����1,��r%�I��]���=����������zC�8S��±��i��\�����_
�����:��9}��s��W�') z���@�!Q ��n\P�
��8F�Yl��h? �br����+��af��F�N����nt��)X��ujيLw4��A�F��Xª�v~�~�푆�J����@���η����彵:ے�P۵�wVSӆj�Y�.�I%�ɎĬ�S1i�$�Y1�t��s��%1qWr�Bv쵱"��*3��&ұL9�sb��˸Z��<�i�C-V�y�y��[5����;q�Q([׼�K�Oq/Iw��X��Lm^��B�u�]s��SV�i^'Zti/!�h������9&Jؕ��l�w2S���E�`�m��x�&nve���j�Q��p	_k���R_������=�P��vڐ,=3I�����I��*_Z!�1{Ɩ�Ԑm�Ij����w}�	���H�����]�L��
o�=�tzc�\���svbлzɆUs<*r��Ҟ�$�{�YI��vp۹����\7��.1"`�-�l��LP-]�_׋*c]��sH��ܢ[�s�Q_A��T�{�ԐMԤ��^����w�wE0�j�1EuBɣ����J]�s��M Q� �u;�f)ə���@�������*��1�aP5�@-�Y�K�j�I��:�[��qb�d���b�ٝ}�Bm!]�<��r�N�����2�fo7xE�a��j-��i3B/ �Em�/w�\S\�f?' �ca�������E�3u�!�Z�
�_M_��I��/��7�ˢ:��R�Ɍ���Y�I>-��|���x ��ûͷ�G��v8��T_�V�<^;��W7�P�|2�;Y�Դ���\�'��=Êp���4�D����R�9��n,|F}�Ri�ᅄ7�(ɘ�̏�ʚ(��J���r�\��b���u=��nE;;�ՈS���U�-�x:��$�|i�[H��xnC۾��3{�y��8ŋ��t2�Uv0x�0�ڲn5Nߧ}�Mv�'.�10�D?D�I��N�ٰp�&@�TY%�y$o�L��zg���9A�.�1i�q�$g�n�=䚹�c*��zỮ]pڏ�js����.��Fy��]�"ܽ�����¬Za�w})K\2�z�D2:۪<����MU�O{-�f��Sp9J
Lu
�t����P^N��|����[t�E�
}�μ:������?��?�j~�+UUU�4@�I��DP<|\� �"�/���K3+��S;��z0�>���O𽧶��	 
!a�H�ؒ�2-B���!�p�w�%"3�!2�Y������:SkM9>���kn�7�:g�O���s釚���	�6w=��d(�|�G��,�q}�^(* '� rAP?$�F!%hr4��^����l���뢗�P7�e��^�	8w�( ��@�ߌ1:l4�ą�'Y0;-�kЍ�1����5�3�K�7ٸ}m����^tl�'����F5��+�'UO7�W�0P*����+�&���Jt�p�*���Mj"�	��^�����i��o�'~�")G?(vi#U��
�=�k'�˶���<DP90�$io�g�?�Øj��'���2�Gǯ�#��������^���B��}~�a�@���c��b����c�g�z�0A� 	F:ވ� '���h��-�����#�Nu'#�"��/�}TP.��H���4hDϙ��A Ham#c�u7q2�"֘�%��.!g!���z�@L��KW	yQE "���s��]���W��х#[�X�Bz~i��ۘ#p=I�h)Ӗ�Me��l8��<�zc�<T;͉O���C���P7�
��#�)��;A N�P�0(�D�2פ�8�c��4�nj�ᰱB[ƥ
%#t���^<��_�������0��9����P7�J8p�v�S9�R�0fY;�?���Nݥ���x��5@���}�Gʞ���lx�Z��ߚ
�	�v�Qp�����ݵ��+�l)/)��2�}AȕrЦZ˟�]��BBs5v�