BZh91AY&SY�k���~_�`q���"� ����  bE�� >�         �Ԓ�iB���� UR�͌�P��TJ�Zj��)�H��R�
B� ͌R-��QT����TQQh�[b#ci����B�+[A�Щ!������CA�B� 
J�f�Ke�(����4$V�D��5ى	J�Mx �v��U���� N�J��w6�m�$i�*�Z�T�U�AH�a�Bm���-�IEU ֆ�B�U6ңm� #M*�  �%$�(U#�i�(4�(̪���v��ק�nƚU3����hj�i���ѥ���)Ӑu�W{�{J�6ֶ���kX7���Pe�A1�)@��E ��w�% M{����փ=��]��	\��<�jT���zU�m��/uo{N�J�^9z�P����r�=*z�)R��{��j�=� �P�W��ԢT�����(�O�JP C��R����V�=à=P=������5��<ޞ�Ԩ
x�鼠�R��^�5h4��<==�P��^Pz���]��y嶴�uʻ���g�^�*��)E l�礤 =ϟTsf�[S��ʔ({e��v�J��`-��������˗��*T�4=�����ڕY��ޡi��sOn��T0=����a{�v��ゔ���J)F��>�H �����QV�7�m�P(ίs�餫mO;���[�u���M+;��D^�U�G �][*�n����)�n��斠�Zj�9)�aP�*�m	
{� �B�_sm�*����9T�T���Y�jP�J�N�\�M(q}�]�G�(;�+�@R�u�ҭ�R�-���lmS4Z�A��J��66b��
��@�� k�m�:'p .N� zxmm�F��ZP1� K�nà;��� S��
���b��!M�x��(� z1�4}9�}���GA��t ��{T(�G��� u����ݜ zt]� �@q�H�)N���6ٌ)��J@ a���kz;�� 6WpI�.�f�� F5`+��@�m.� ��\��� ��ED��LƊ�(RWϤ� σ�[]}� �
�Qj��=���@ lw��Aq�� ��)�g�p=�ί���� J�� -
 � L�)RL&L&&"yJJJ���	�M�d4фbT���U4�4 �  ��L��J��      ��% ��� � @� "&jI$bd��OSSL��2== OQ����'����?���术��C����V^L�Y��X�����>ʠ�/Q��( *�@EO�@@U������?��K?3���������?�* *�B��O�4* *�����S�" ������<���F1�b�ضŶ-�m�l[b�6�� �-�b��-�lb�#��m�l[b�ضŶ-��b���b[�6Ŷl#إ�`�-�[ �cl�%�`�-�lش�`Ŷ!l[`�-�[��%�`�-�[�lB�L؅0b��!lB��س5{*g�oe^�^�{5{&M�b� �-�b�Ŷ!lc��b�-�[�lB�S؅0b�-�[�!lB؅�i��
b�-�^U�٫٫�W��g��Z�-�b�-�[ ��[�lB��b�#m-�`��-�[ �l؅��[`�-�[�!l[a%�`��-�lB؅�bS�0b�m�[ ��BشŶ	lB��`��0`�Ŷl[`�-�hb���`���m�l�[1m�l[b�ضŶ�`��4��1b�ض�-�0-�L[`��-�m�[ؑ�l��m�l`�-�[c�Ŷ�m�l[b�ضĶ��6���lKb���b���m��lBضŶ%�`����b[؅�`Ŷ%�m�1�1-�l[`��6�-�l
clb�ضĶ-�-�lK`�ؑ���-�m�l[`�ضŶ�m�lcL`���-�lb��6Ŷ-�m�ĶL�6�-�[ضŶ$al[b���m�[ �m���[��`�bF�i��-1m�l`��6�-�le��-�l[`�ضŶ-�m��c �l[b� �	l[`�-�[��l[b�-�[ �l��)���m�[��[�lB�%�Kb�0Kb��-�[�	lc%�Kb�-�[��#� [�lR�%�Kb6�-���c�l � �#�6���m�l[`Ŷ�[`�V������U� �E�"� � �U� �� �@-���@-�$`��P-�	lblb�[[b�[B�
�
b�lEi���-�	l `�lDb�[B�L m��1E� �� ���"�� ��
�F0ت�� �V�*�V�"� [b+lDm���� �6�Fآ� [b�lm�lUm�-�-�����1���V�
� ت�[`+lb�[�-1T�*��؀�@�"�-�l@b�[Jb��@)��lb�[ � �V� ������ ��Q-�-�U�*�� �*�@-�l�*����T-�	lUb [B�"�ؠ�-�!L@b+lP`�lB��m�l
alZb���m�l[b[ �Ķ1m�lض��l[b�
b��-�m�[ضŶ-�1m�[�6Ķ-�b��6ŶSش�-�l[b�ض�-���[b� �%�b�ض��`[ ��m�l[b�ضĶF�-�l[`��6Ŷ!l[c��-�m�[ض���-��ض��l؅�m�lm�`�ؖ��%�b[ضŶal[b��6Ŷ%�m�l`��i#�6���-�[ضŶ%�0m�l[b[ؖŶ-�-�lcb��6Ŷ�o��@����3�>ڻ���]e:��Oq'���^˗yb�S�]p3�Tv��ت��Y�68����I�X豻���A����.�MG��H�wq���,X����Aa��V�ި�C'5��U)���H1x6C��������h٤�^Q*��Tɬ!�Ä����[�Qȭ��"�C�)��*�ܒ*���À���r�λ5�+q��  $zh��9���mQn�ۼB�d�>y#Z����X����V�:E����L}n���5w"�I>�E�ug/V+byvn�˳�blˆ��
�wq]�yY�F*ҫ;vb�R�z���7Zqr
�Ie'�5��ds٤��I�X$+6laP{,�ɪS.�&�w`λ@�>��aFR2�.�ܦ��7{SZ
�=zf�!�i,˛�n�ܼT�:T{KE7�5��Q �%�do^VQu��2� K�ʽ���:��yZQ�5[��x��l*;,XM9Etv��/Y��R6�o�0�T�Z�۫�]��n�)F�7s]�@���3aӹ�fc!�N"l%� b[���� ��ױmml�a;��t���n�h�u	HT��]��m��k������ʺ�z��� u	t��76�r�MTF�w1�]�/w]�#%IH�pm�+X0����f=�m=�#9V��#tŗ��
�A�5P�wP;���Oޘ�V��Rs��L��ɬL��0��.�V��x��[*a�1�j�G�2�^+Y�&����F�+{n�b��t�u-�t4�xj�<\Yc8�ʫKf7i3׆f>�]�Jؚ�9����P��H�Ekd͒����'Tjf�ce=ҁ�)��r�+�X��%�mo+��4"��US�S>N�;{>Lg�f�0�F�r��SS����ÁM�]�!jK��5b���xU��x�֋j)P��YX��7����D��T"-D۫w��UyV���F����+�nbY��-%*�$Y��R;uy2Y4���7r��J�d[TG5i�����b��t%hآ�ڍ�˖��t��
:��fĄw�̨�Gb��t�Y�ĉ���&eO%4�R�^$�/i��Q�-v8r�"�Gv���&ފ�I�-��oe�3%^,8��i�ҹ��ƙ����`�nf[���U�<�0X5Jy4]�#i��[�3v�Q�u�\�ӡ�t�=����.�!lݹ�U�y��٫�+y���K�&�ޥ`�+c�RZ��6jL�y5L��"ڃJ\ײ�˻�-n���wp9����J�UM�j���yXVR��6&�(Z�f�ږ���W����Bbr����d;�P媇oʐh<:��n��7f#Jͪ�2G���%i�NԱH�D�m�n�݆�o*|�����ޔrU�y�&��ǲ�UE8J��C2��#�V[����v�"7�\�1̛eI�=�6��:WYP�d�-$��n�h����C3����t¸l��P�.U�U75e���%UXR�����E����n�7�S0�O3N�2�q�$Ӱ$��OHϘ�5�R����k/ֽh�Or{eER�j���AYVU^]��ݪ�"ìAT˳��iՋ>;�bEۥ��V,٬�M�b<Jef4J�+6�E�I=��w��lv�U ��v�DVe�J�G��7i#�Ď�΋�r��Ѱ�r�U(�OH�{��Kpٺ��-��wRhT��+���dh�X�2��M#�̣U� �v�]�f5)�4�dRM�qZ�F�T9 l�F�\�6m�l��i�Q�ԭ�wcv�qm��i(�sX��Vc	=�+��C&���b�b�PQF���f�]W����n6�d�v���4�6��z��a�hVPm�]݄J��%�ݗ&AG\	�6�ʘ��in�-�lM;�ܦ�ڤs�@�d�7tJ�2��Mf��ێ*8s��Z�K;t���s�I��Mn����Q�]oqe���QYR�MڪV8�.�a���`H
�jז�ao.Ǉ��hm\�Σm��Ę�`��UJߍT�^�(!BeH2�SE~q8F�z%�x������E]m���Q(�MZChj����[n�Ҳ��3IEbN��h�YuE�*�YN���rTP���-�]
`K;�+�he��E7V�������.*[mK�康)[2]��1[��mҫ�T�m/)���h��۽@=���T*���؄�h��[\�Bi2\�	�[N�w�Z�1�{	������,c5a*�D׹�e�5͑퇋q����%�k*+Ք�)@��^�I+!깴�B7a�/a�f��0�1^
�z1ܹE���9FkZ�^І�w�݋q�6^+�%5�� �x�ZL]��Z���5V/K��ՙA&��"�ʦ�����ȓ�](����W3q�ib4��`�cÏL�QZ�b��Zjf9W�h'rPU�mѩ-��f���I�m<"<��\�4ވ��J)�J���,ۏ���=:J�ϝؔ��^jz4T��%K-��U��Cv���q�k)��&��՛*C�f�k5�9������mFV;�*H"���8=eh�����mm�۹go�8�E�e�������_�Ǖ�t]52�nTAAt(ؘ��FJ��1�iǙhD�57	�2�����UCx��,fz��0 �m1�=mÚ�x����D�洰�D�,,A�=�p��^�mr[�ڕ�+�J��k&beL:�C�Ī^:�X�yO+�VqL�L��&����Ѯ�:˝�����ŎJp!Nk����R��Lq�fV��6ȧ3+u*0�ݥ2ԗ���뷹7+"˱��[
����(J#����]`ܳ!�����L[����kt�cM+��yN��O-Y�R֐�9wV��Ȓ-Z٨A�5�2ԫ4fVqĹ��Dq�nt1,Ed�8fv�̅�4l +��V)rFf�*(wB��Rm֝[��儢�7<������w��և{bd�B�Qe<l� ja��Ylh��b��VK����t��t����%`�1�ě��Ӣ��r:E����ohR����R��;vM�eV�۔�%(�iW��3x�Ar�ÃN5�$�����^V62��V�l��ˈ��P�2���8N���4<�*&t!�E����Up[���+�X��<w�D[x��G���N�&Ii�+!�Vr�Y�mw*��r�РA"!OIU�e��5��=��m�[�/ �*V2����ݺ��e��ъ7�ںwR�@�f�7���S]cM�xP�.�ٌ�	�{nl����ŷ&n��4&�"��F�c)8��i�.Zw��m�y)[�{{tk=�fҬ5����+!��.���([�q	Ŗ��_k�H���*�l���2$t����U)/��\��v4�{�P�f�,�&D�F���6��6�;7&�TF���ӭ�ݨ�cA̎��;��E13K�$�Ƿ�.��<�[6e��{rj�dܔ�^�B�7-�-�'�]�5l���N��ؠ����B���"��ȯv�<��&�B67P�/R�50-�*�ڡd֙�%��J��kn&#ML�Q��-E��)AEe�l��ˬ"���b��p���naB|t���X����N�)�[��#�wh)M%��A�	�ՠH�i�����FEE<՝��^�*j�X&Ex�f�۳�kn�ܐ�)�iՍj�q`S/,SOq�^�� 鬽Rj�EZ�	�n'p5�$��nfR�X�)�t���4�w��	K�����(آ�EtpB��5S������Jy,�v\aP��D�����hs��J���o4#�َ�Ѵ��yu�qJ� T�S�ڐ@���E^7��1v�`[u����*�[~"k����תe�o�9���YLv�d�I f��XV��9u"��2���-��{�l��;��Ԉ�GC˔��T[����
�4q��%ܭn�a���+5b�z�Sy�J+\ȪX�򑣖`~;�*6���T�f[�V&���g^3�D8�~�b-�7B�@�X�̭ٸЙ�!ih8��̆�@Z��	Gx��>��YٸNN���Q�2�n��%'*R�+�X�60 n`�hC�tlZ.��wPY��#���ŻN?���eN��z�SQ��b��z�]����i�>��#���m�
�2����'WX7i���l�Xi��f�U(2D,4M`>ѭZs$b���f�b�t�e:Z�\���#*���̐Yx)A�3cn�ͽ�5A�!Ak����.�YZ��.�%��/)�X�#�a�ɇcV�U:8�kP�J�vM&�էX�wF�jٔ�m�;��V��M��uLڙ���7��t�X�X���v�h�"�X�i��Z�2ػ��Z-��Y6�p�(7"{�Cu7[�����p��7
Ƿ �n�e?\��`l�SPɑ���a+�k����,�܁f��Q�a�rd"+�mKw� ����Q9�k�Ŕ0\�ܲ�݋N�@5�c:�b ������O�=k2�$E�����:�[P�BTGo��٘�kmj.���{mZ�e�{��-m�&�
Jx��q&�x�n������fZ�v0q�c�X��QِD4VVC��wQL�+=7F\���fnX:p�8 -�Gʠr[J\U��ͩ7]�q�osbSv�m@ͭ����a`�.����L7���ޡ�&'���2��mJ�:�`30�LLRͲ�j�ll�'����0\�2ڷYQ��zMe���RR�r� ��%i��FD.�ݻ�y)$M������D�V��<�.��SVҸ=5�L���ym�ڱ7&��ѳ6��t ��2�P�,����6iܼڥ�6����Z%c�i�V�}��Q��h�t�)����ƱO �d<v���V�MV�B����bο\EICT�
H���I�dx^9�]A=2��Ą�e;��+���*lݒ�m����	�C.�BU4^��Lg-J�j��G�fhuum�R�d�k3M�X���@��
�ǆL�t��Sm�j\��R��$�1�wy,�r\��RXݙV�Ȫ���0l�*ʺ#�ຶ���<7+YD^;�#��M��T�L�s���[̹(n`
휖��������J�����O4��(+�ڴ]�7�3T�-k���<�\��T��%8UurUӅ��D��m����
�a;7"�������N�]9F�ʊ��Î�NP�Ji�Ch���i�N�X(L�t�Q�ѵ�J�7�KA��	���(D����������e,zu�.� ��m�f�L�U%]"(��[����&��F�������{ B�6�5�wSl5P�őm��\)bD��2lU�E*m�� �0P͢���3"�Z�"Ƽ@F�F���5AU�b�2�;:03jUC,ںO6ȗ!Cn��X4y���	�bfƷO ��3.^e�s2�SLfTn3vkbeM0L̥�˸�m�����[��⽪sKɇd���V�C�-=|�h�F,����3%ь�q4jdEh�b�B��61�,h�4�z+P�o,4
�e-��XDĲ\ɒķV�Y<-�	��N�1��5�H����VǗ��e\������Ĥ���c��-w|�E�{r��ʚ��snV���ejUO&��N�U�{�] U�Z��vn�c6 ��MA��s�J�[���J2wa�L@T�%�V��܇n!��.:��Ҧݚ���z��f�j�*G���Z�`�Y,3�upa8�B�}-C�-a9��ʕ{���csV�U h<,a�Y�A�����s���p��Yh�5m��V�֓5裻)�gj�
�UL$YEaU+`�VL@��eZ슡J�O���P9$�n)��t�v��}X:ޱwzܕ��y��	6w_��*XX^�q5�-hJ�a�/e<�k��0���o���7��D��$C����֤qIxO\�(7�Z��噇R���K� �Tj�X�3eul�x�)�w\��+������,�ӌ�]�v]"�ڤ�-���S�D�mi
�����Y|R8��("�a�o�����n���d�t���5�{�[�h�n��$#zE�Ӑ�#'-H�il�bR���IOq6�@Ȉߖ�3��[�Vt;��wI����.�D�I~4E��ah�M)�x�>W�2�0�*�g����iL�mghQ7���\�.�V&��6ib際j�x�Kfq�+�Q|W��/H䚙x(�:�ⶈ0C��6�G�j֍�g���N%�—�'Sk�J���:&�N,�-*Q-��Rhb��Y��Y�.�����Y�D+N�QV(����J�I�A`�E#��)p�fYp�;@�����iG:gRXfC(.(��a��=�ac��]F�M�e��6��YL�7@�6F�E��*�%��'�5�\T�1;_Zm8�9�̔l�v��H��YZ_ż���H���5��:M��X�=��jY��T�(���@���-]�E-u�J�N���N���$����@�]E��)d2x�&i�b"������%i%V����%�D�@������m�V�Ķjn*{h�5]��MV��!�u��0�	��4.$q�	n�q�	UJ�0�e��+�����G��G�0�#K�9��,�%��$ŀ�k�5c�⴪>R֔J�F��!��D�MdJ��%�%\EV4y<�ٜ�Q��b��j!��$yq.'��l�%��$�A�ah�UR�D�S2Ѹw
��AK¶��b�gaM�vWbx�I%*t�Iډ&�,	�@�h����q"	i4�P2)��=yv-�YB�ʥ��&���Q@k�*S�Dͤ�E�=Uh�mV��`�7Chv7��x��D�z]���A"'vrlR��AV�F'�Q�f�n���6u�E#,�ӄ�qBlQ�e�4�F�׳m�q��V�	dP�=fAIJJ���]�T�fM�Ū��	ܵ%�� ����$ޓ	���o���!uq���?v偏�������J|B*����]�tH刃���+�_^��/����}yI��u(R|��=�'�B��c��[º�=b��|��e�^ʱ�9���Tj��8�1W��ybV�b�[d�P��'{Gt��.#��һn���nJ�5�U���эk�m`�����Z�6�Ũ���W��ֈ��Dun��-a�X�pe�3�F�q[���Y���XBcha��0M4��B\&:13�j�S/�;>���#t�h�NئE��8m�!؛=��Fu�Qukm]��m�g<��n��v
��.h��:*Z���w�_ǃ�Nʅ.�A��b��g*Ӹ�[��k�{����������9��ޮ[��w���;�t/��s-.�I�dJ��b�*�w>�w[V��φ5T9p��;�r<\_T��/�צ�3î��N�V+�R��Ǒ綰P��9�����ѵ��s��@I�N�˲㬲Y����؟7=7!����[r�4oku۝}z�8�Y�`:�����e�I;L�Xvt��}N�֦�x�5s`�lZ�Գ]�N| ��`٭��pb��R� �c�J��d�Մ���8��݁+��	U�vV�=O^e�OmH�ګ�s9�Vk�Mk��L��W�R��J:�\���[͋l��&+�i��,��7��3�V��{�1n�ȧ.t+u� ��2�v��]�w0�8��u�ĻA��w��ru�%2��T�ay2�s���x�B�vm�
��9�]�S������GGh<sdJYЦ�=�M�g$R�$7R��`���t�pΓ��,)���C�/U)u�ם�Tr�ୗ���L�V�y�њxI�����95�6�V�ۣ�ؑk�1��:>݉�ٸ��^T�2T�n�p]���}{�v�t�yl�'#H��:�D���&��uw�p�mod�Nd㊻��^!�O-�w
�z������ˌ�:���/�����gc��v*�uݥV"u���	,�;Krad�K��о�ixHYMu�K��,���C���8l)�]�.�9ڇQ�U���ɫ���i�|9����&Z�VK�٤��x�J�%y��R5^\�J#E��3I�m�b�1�F����7ڼpv6��f�v6n�3f�^Yr�3p��9|S���V�y]�݂>�\nP������Z���ae��:�;2wWY�^�9��������	�r�I�Ζ.;���Jq���۬��a�����Y���^x�ϟ**��T���zm�kk��6��׽x�:�ôEJ�Ȍm��҂���ѓ�U�#=d�@�Z�yj���mi���Uc������$g��r��M �Jv�Lu;�U��}����GiY&_�n0�/s��#9C
�m���C�Z�Ps�&u�tIz�c<�4R�ޔ��^	�_#�[��!�Þ臢��u�W`E/mڐd{��5ؚ�+p�u���[ͤ���6�r�J�}Tm��ܝ��u�6�k�Ƿ˫��b$X�s9V�Xor�f�R/����l�4<ڻ����h#����;��yp]ڵ�:�EÇ��x�h�6_8�6�H3�YݼВn*]m�~��iopWWj/����l]�y�d�������
���Ta�5�K0;���k3�X������P��"�N�TM$��A�^�3wʕm���U�0�εq<1Js/-�.|��A��.�_4��y�����d�wZ/X���졘�sST�^L��T��I�������μ�����F[coa���3!r��w-m��6]��8Z����2k�2u�t�`�Y���j�\�/zL�x8���M�Bu��iYʚ�K�i��{�]��V��ӗ�&C:����Kt��7�H"wt�X8�MwVY|V��b��o�t���"�2�G�d������p�s*�m5+����%x�C	pѭ~�H�۝�G�X�v
mݱ��LSx�no�Q��X�j�޸� r���I��ܑ`QP���9�ɹ�KUtV���"��<�Do.ۼ�u��gb,�Sδvef@�o�z�RU}��u��h���6������u\�`����j�<vƦ/�Vy���"���`<�,	Z����Vn�o�����!Y3b��é�P�E�,B�:Y��ٸ�J94�޽M���[�˕Yd�\��9�;ff��+eb\��ʆY�`c�7S��y����ũ��1���}S����C[�����#�r��v�<ӳ����M�jTe��\4M=�Ţ�kNفn�t%譫u�(l����Cq��SJ�1�[i}���L6��'.˶Jq9�ʌ8�ᝇs�
�_3`�Y�v�P���n��c��cʹ�l��ǨŤ�(V-7 �'6��7�����*���y�л]m����6��X��8�C�M��[
ˇ7k[:aJG�j�J�op���Ʉ���7��sN��Fm[��:rQ�l k�$w��v�ӸBs��Sb�ܳ:Z��`|�ǝ�yj[Te�3�JK2��û�a�j�.5o�W�Os��5�c#{$w�_�������?����w<������0yx���N'��GA��2�ᕛ3v֘����Q�n�ŗ�+s�l����oP�Fe-"�G����nX}[���v[$Ǝ���G�ˉ���׼��$�2�G�)�`�܁�� ��N_�[�܆�)b�1񤢶����-�g �U���G`�*`�uܦ�(���ӎV+2}��묷�S�Kp+x\J��YyP�[}���ȨXgv���P;B���`��g9b�v�A��*��V�ᷥ���n��*�*��C�.��hLԯz��llǔ ݹ\�-��-����ᆷ6�#��7��{�*�݄&m��h�V�)�u]���e��+W!���ob���G�`����xO6wN��\���l������#Qp�WwK/v]�µ*�`#��o�boWQ4�������;� s{��dwd�y��a�5F�7:s�utr�Vr=�ԽZ��P���Я3U�6;+xNd*L��z�J̢q��J�-����&٦�էd���o-��l'���

h�����3JҖ0��N(Y�Zv��x΃z�������ٝ[ot
�@�u�});�f�}sG!gELԔ5Q�g�[�X�렔���,�B�!lm͑���*e����k���<�+!�p�˻�n�NQ'u2�=kR0��˩e8�0埖�Ed�fCz$f��{s]�0^��y�MkZ-�5W�0du�1�-�TOU�(�T��r3��Y����v�v�7 04����n�7}�.k��t�����]h�˫]�A]*3���Z��Gb�oA���\�K��2ͩ�D}�}�/P��yX�b�3�X�w�3��g�hv��ԏ[v�*۽�h,�z�E����9󕻧e����_Z�0�6���w>��B�z�ofE����Ә��h���Z�&��nl�+���z���+�-��ES�[�쁔�0͔BC��7'!kS��ҭi��Nu��w�(=Z[hXU�z��B=�&f@B3Wgn���n��ٽ���cI7�(p�%�g'E5����6.���ݤ�MtӦWD`U�J�#b��ҍ��7�_l��d\�N��3w��ET��FH�w;3N�8]�<*2��̚5�0w`����Ӎ���S�3[]YR*�D�����;��!�8kK�����辯�	��}Fd8����Mw{;�aF�øM� R�*�jP��2�����c��"[|a8v����5k����VT9x�sCnJ���O�n�Sq\[Yu���\��Rvڽp���Py�nmɉJ�Y)^*2��RS��KqGm�6
��i��/���;c6.%��ME=�O0�%�e�ॻ��-�#�hwW��b�m�YV�˧���W*���d�H°�7��4�!�ټ1���7�7|��
������2ӷ�G,w�5���z��o�����Y��Fe�N8�u-�y��J��;�Y�ie��j܇v�[���9Qˇ��,�:���}y��Moh�����w$��uf��+wG��voR|��Z�oP
C��kz��;ͮF��9ݫ{v���;��%����x;�hI�S9Y�V��̉��C�����+*�3whlW��1\E�Y�uM)��$��Vel�U�t��n�7���-����q.nnc�Ђ|�͕(�w�b�e�G����e^�y�,lw�Ǻ�f����[4M�0����xP�ڝ'f;;�ts����6�͵����WR��n�$�fݴC�b[�2���w�ۄ���|m����nM��w��
�Ց���o��X���މ�E�f����NN��i��]]��9Q�7{F݀/��^���@�]����ٺ���*�v�/:���˝W�؎��m^�x�����6��a^u'S�I(/�8+�U̘.�%���g���J7�i�圹M�]ὐ�����i�	{��V.ɹZ�	�I�ֆM̻}���ogi�a>��7��vd7��Y�ǳ���Q�2.��>���[\�)�����A�c
1wT��Uj�ӻ��:�S�GB>R��v��o'I�[�O<pa�1v�y¯�KH���$W	�5]��3Hr�.5����N��V��_t�����;����J���⪬bj�t8J�Poopm-�q�y��LUn,��&��e�I�};���vo`�ո���xb78V܋V�锩��j	��q�8��e��@��g�53-��`'�w��b���qk[�qI�f����$��M!����M�`9y&'�d�m��}GY�e.ݲR��woS����[�5��VuwY��O�-#[�G����c�,��ׇdX�.�zڰ{�:��OҞ�æ�q̚��*cެIIۻ8��OJ�K�v�=�����{Es#S�F�<{=kc]��f�H��U�ם�S}ӹeFe��7ThX��7�531�R�VJ���x�N�����͋���ث�i<%<ŐM��WW��9m
�b�[)nS�;Iu*E�����U8+/�>�tu(ά�V�+ˉZ�Q�"E���}UMF}��nq���T�IŠ�gv�k��W,�c�;��Z�\�Է:�,Q�&�s��M�|� ��{0����L���96D۾�"n�9J�(Հ_t�v�_T��V��]�7J�[�(r� oU,=ٶ @�V�2�긵�4�u���ُF^��6�u"����\�˜s���utpR�
L�Q���b��e`X&�j�	�՝4jL'v9�(;��m������ZR��w�{��1Uجډ5�=�'S�$��)$�f=��%����C#�o��o����rCR��pYn4q�j��hf��>>�аs�6�[Y�&�V�J�]wN\��v���;��Bo�uz�'�Wi�;$�;4�9T�}�Ju-���rm����9g@��<���˽)c�g�9\λLG �렴�`jH&n�΃ ����=E�y4�m��<��ҒN���_'o���r���FevJ���PN���Qw%�Ne�cF��7����)����\n&���ǉ�}Q���F�M��V�}Yi�XEm�:�!�1(��@��ض�L�{Ղ�:�+�
g���i��t���M���t�UqW)d�=�:Cs+�.�/��.6m�k7Lɂ֋8�uG��pKze���J�0V�C��vű�C�jϴ�⫤����q�t�¬�*�Μ����_\�a�dM�v[�+�HMSw�ə
���u���1�(S��u�7D9ݏ�/��U��b�=�9�s8���S0g.��'n�{,�P�`��;û�%�vE��DZ�s�r��wz�����/eIl��V��Vr���5ʌ���`�����k9-���{۠����;�28�W't}�n�f1�"9=�;��j�P�|��x�U��Ƭglw����^�J�rΡ�2�����\��X�������=������"	�ՙ5	�NJ�����|�5�
��2"�Y��`*��n
r\���p��I7�9���%r�=��5���P���� ���Fk}�/��9�Py	]#؅@2�55 <��<���sT��V��2=��O!���P%A��k�v"r��� yQOJ㡒ġ�b���b�ZG��8pՀrv�kJ��R���&�zC�C�O�rv	� v�;�5j��' ���k(^�]�j���j!7@T�^�V��D|���О��� ���H���<�CPS����;� �<�9���&��.��A@G����~:�}C���?�~'�����#����h�����~%~_�ti����p��oΒ贫eH����f=��7C�ՂfSJ��-�bj�ⓕ���P1wY ����+x��k).�
y9���0�70�陦�c�R+4z�����P<N\eq��y*�,�������l'�ޙg)fSW�#�l�r����]�ܻV���&���VRIcGڬ�p�[��GR�F�l;�	�.֕ ����M��v�*V��Z�=
�j�rp)X���ǦX� �m��Y��>�
�GV�V�H9SEI� �:(�Ѭs�`��J�Y ƣz:�W$�]*-"t����ŧ$Ι1Td{s������N�eΛyӹ']m�i��˂�)k�(�#%�%c�ݕ̸7h����y�q���m8�[6�S�N��c�̓��)���}Y�*.&��Yq��cmᣘ��bJ�s�o��.��7�x��ͮ��̓8��[}ʸ�M�\Uk���)��H�<6)!����-�X�u��1�yT�ڸ���h�-[Ѭ�ͮ�P ��{�^���vn�X�Uu����y8�윍g!$�R�H�:���6J���P��<�]j*SM)�9���D��%f��K]:���<�2sz�_z�맮<qӎ8��qƜq�qǎ8�8��8ێ8�;q�t�8ێ8ӎ8���q�x�8�8�q�N8�8��qӎ8㎜q�v�8�>8㍸�8��q�n8�:q�qۃ�8��q�8��8�8��q�n8�8��qӎ8�;q�v�ӧN�q�q�z�q�q�>8�n:q�q��m�q���:q�q�n8����/���v�^w/�5�h��-M�Z�e��q̜N��͋N�� m0(P�GVN�#��;� J�;�{�״s�V�۫��6`5�T�9�]n�.*�6�sgjO���L���@7Y�<-�r�_pͤ�WK@��)�9�;G-��[��$.Ȉ�9�E{��f�ѧ^��+�9���we��֘A�b����\��d]�NlmRH]\��eP�N�wvJD!����W!��6���:����j*{��]��*IHt��\�o�U�z�p�{k{b*�����l6�D�ǭ�,*Ń-Ss4���̶@HU�!]T�`��,a��(I"<y�i�G����OD�W�l([̭P˧��go#��W��q���@���Kڮ}r�k37f�fu#/���q6���2�x[/kno%j�^���'֬����m�zE(�]hM�dpr^�t����K�#����*).e���@r
���L�V�W���˳���v���êmr���o[>�9�65[y����kh�E8��,q>Uձnn�N5�&�Hի�h�B�e�Q���ڜ�S_p�D����kh�w@�`*f$�W��x��}W�Iv�Du��g
��<q�Ǐ\q�4�8�q���q�q��8�8�<qƜq�t�8�c�8�8��c�8�8�1�i�q�c�8�8�\c�8�8�88�8�<qƜq�q��q�c�8�<q�q�1�4�8�8��q�q�q�q�q�q�ݻv�ێ8ӎ8�8���8�8���q�q�q�q�z�q�q��ʭcS���9Sh��Wc���z�u�AÚ�X^��=n�Logdǻ�۫�Г��;���`��B�I��jlAG�b�8�2��l��Q��*`�9e��E���w����f��h���j�����ɳMέ�b���R};�zuQ�c�0�ČR͛yjf�Ǩ����v���ľ�3"�|"T(�+�>Q5K��׉�ӵ����r�^��EP�vެZ����r�]�hP(�L91q��-<�H2"�'9��=z�	��	����V)�\��]=	���Eʹsw�Ł/}Ğ�+ �;�ީ�.��A�"��.��{Y�^�U�LҺ�u(���.�⼹8���	|��_v����U=�+"˻a�qs�Y�ڸ�VSr�H�ѠB������ �ڍ�pؾB��{U�%B��e*�V��+s� Blt�sۆ0�ݧw� �<�Z�ǽ`�gQ\!S6�䆹y�8pԅI/�eu�a�.G� ���7�i]�{�)*B��^�Vw[��:��y�`��We.�`�L%�A�Y�̛�]��;��C��44�몃
���)v�]��V*�q��DY�ZZb�=fgd�QV��VΏJ�:>�f�i�Ҧ�����z�%[���ةW%�Z�w�2f��nu۷Ǭq�Ǯ8�\q�q�8�N8��;qӎ8��i�q�x��8�8��q�qӎ8��q�q�q��q�q�q�1�q�q�8ӎ8�8����q�8���q�qǮ1�q�q���cq��8�8���8�8��i�q�x�ӎݻm�q���:q�qӎ8��q�q�q��c�8�8��c�8�3G.N�W+��k|�y��]�V���Q�cEX����-ȭqd�Z&^�2���m���۝{�^X�P7���f�db�f7�:�3�)a�)��_>���nӬ�Q�i�˖!��ә�SF�H�27��:MB�Y�s+nT�]��Z����h��sW9���;�;e�.yu�ݱ�A%��\������=έ��ۙm�:Ԡ��v�ō�y��]ĴK���Q�om:�EiP�C��s��E���x�)ˤ�Ȃҟrk�:�4�ٵ�2�ɧ�Di�Z/�23;�<��엒)��ة�	J9}K{�p���tn#zEIu�Ԥt�5#�k�vl뙔/k�;��1yhj�m�
�;��W�Yӳ�;�����)���y�NF��°9���L'y��_/�r��	-Z��9J���4	�]�i��{v<|��)c:��⭂��r��\9K�.5R��ʗ�]s{k6>K������f��
�J�#Sޗ������:�B��ߕ�Xɠ+�Y�.|�pk�e�[�-
�Ư�6��J�ں\j�+`�$�:*."������s���ɲ���6�S��${���\V�����n�B���:z�4�K.�,��'H>��VuB{�=v��jW>�+�^�w*)x��ٍ�V:K�����Jź�,��X���Jĥ❱�#��(����6u�M�-.�S��_A����{l�%��,�[�;��j�+&w.���S��֭
�t*p�Z8���H��E�����X�7f��姬�+�΋h;;����,��U�hO����oL#S��VѼ1,ZD"�1>�a,���٘�f�ے�����g�lG�i⎳�v*�w���T�Y������n��*�gF<+T=/訹��c�n��T�W��'{$��F4)c�vAaЖ���L�8o��\�{�U�}�n�֦���A'�e#�D�c`����x�r��k�k��%���-o��.)��#�[}\�uGyv�A[{Y��^⏞�5��n��9.����;��u�W�\�{73��҂�h���B�*�m��S1�Ȃ���u�F���T�Z���c{�K�1VHW^�2Gf�%�hVA�G�O'�@�L�=U����f�q�!�ШgS�$uw!JV��=�}����*���ڻ��]��n��nk�,��ڵ��p̔��s��(3Ƃ=ڨƕ+�w�2�r���ͯ;�����������C��߅fl�I�ylZ��O���T�v[EX�&ǆ�%�.|{:YT� ˗���{/�R��:��]DG	����K*���w���i��U�>�g+rK-aD��
��A��U�Gc,u�������7^������X���0!ȯ/��i˹���:
fG�_uV
�M}��*��
��s��h���5��V*Cn�1K�$�����4g�;�l�Wj�F-r�t���`���U�k�}ۉ�J5���Ϊ�c��B$A�Ii�8d�L�
�*熮�W8����EP�ࣺюc�j�$��OR��@���B�֢�Q��f�u�����y����,�<�d�2�n��ѱ�8�幗�78��抇-nj�s��vCĳ	`�M��:7�"���86������7�v�:�*�xlM�x+-�P3R͉�Tø��CW�J��Ө�;��n�߾�x׽��9�2�P5���ބ'ܳ��ĽΕ�w'F���lT	�kote�a�7��j9��p�:��UB2{B�;؈�<���5\n���ε��qv��kvd�ZCe˘-2�2�����껩D3��ЇU���|���%X����g�>v��t�.��w!;�W�Z���d�[}A��`�e%��%��,�� u���sm��ܫ(�Y�w���Om&^<���*.�*�U��x�_v�Rqᶧ��Ը���c��M��0$C9nT��S�V��4�X��n�
G�.�2r&�-
wєw����ިY���R�{���j�k�E�F��C.�R�4��kZx���qrm��U7���He����M��*�Y=1M�����T�\�ݽ#�h�_U�E�����nj4 ��P����]�G.�0Xk�R���{����9���;T�t�bUb��e�4f8�#�MR�#84�tOb&�i�͜�"G
IƮ�'�C3a 6��s��jW.������FLY`��m�{y|�����F�P�j�He��fA\�l��L��<��;ܻuk:�X~��!�}��o�w���T�1��Fu�2���ϣ"�M��m�#����d� WLJ���I;��'
�6x)�1*i�>���;q-Ś��꺈����]{w���_u��SojzP�]]T'��x"E���+�b��zu���C��,�v�=(p�Vcs�GW�|����E�V2�<I]���`,w�f� �S��5�9+�;P�V~=�4fs� ���ꒊ��=�cbQ�ŧ�wEUO{*�qо����Y1e�w��8��6��W��خ��U�4Dއ�	:�'x�W��p�w<ݕl&� �۷�0��V^��H���[U�o*v��m��f�)-�U]��1�/yۮׁ�:"Mn��c7�a�.<U�+��Ȳ�����^fS7�0��+���t�
ڡVTuj	j����p�u[���%�h��xJ��xd����%������㶭t4:٦�ұ���h�┣�>�&�CH����f� ��cp	����.��1^>����+��ZA�����pZޤ�%��p}�c�l@��q�7/a��w�C�qa��{3�3K��"�&�-��Z��B��o.��l��l�u޲��Rf�ܰ�S��RlE������y��)�h[��/to�?��./����B�FQ[F(n-˺:�'pgu�����m�ŝ,	�����*��W��Ӧ6"N,
ro;���LF���L��\�ˣC�aV���;��b��7���@�b�uY�M����hL!)�tx��0��mnIû,vj�uݎ�B��X��γ#0j��;8u�(�&8��K˘��YDAmے%��C8=v6�G��u�3�,mz�p�e�-Xj��.*/��`h��k'e��ଋU�nf���A�I��w��W��
�
���
�̬f�4� ��fԅ�is~�o/OBq�qB�����#�^u�MM�.p5���YsD9�%M���9�_]]n�t%���u�^u3r�=���������88Dw����J�3�X�&z���N�x�)nf���׎Z�Vt��x�G�E;1[w���� T�����=��ԉ��� �i���u4K��|�wio:}���HW���[�W����VM��_a<�Q�D���m���!%��	ָ:���j*6�E�!X����%���y@�yq���e��KG{WA+X���P�F���_0X][����K����B�Kl�ߺ_?f��+�����{J�:��h���ʚ��m�ņַ���Z���/�ƅs*�u!��;i�1�� a�Uz2�7oC�S��(��Ŕ�҃#���U���]-��̺0�4�JaغN�{�:��45���r��c"ͩ��gy:��ߜD��*�z�;7s����N�p���x�#��!�N�uN�r��N��b�%WX��2&��������At��]�ZKp�[�yK��L��sys�/]�޷�2��K �5�oOwu��qb��&2ʷ �]��hǔ�R�ڐV��Q��vf���܅�'J�vsSnm��Q�#���r�6 �����Cm�1�u��D�U'{N���l��q��s�9��.�*��c�	Q$�8�r_Ɵq�*Mh�;#�UxI�x�YU(��[9��	�r���j�۝9�k���;W�"'Je��۞YR-�$aߪhM�#t�,uMӝ��z.j��$e�%���V�Y�
ޱ��\�����rc��="g����ѷ�IwQk];�xh�S��v�\�K�*fa��O*��,�np�������2��ַ~nV��bX-��aH�w��x��]�ОO�fUٰ*k5%R{����`M`�t�9���iu�e�li�i`.f�B��2��Q%���*:&�Se;\���m���l���Z�=*�<0Ő���UG޷`���@_��t�E>�9
���y�ީO�Թ2ռ7��vpW%O�c-Eܴ���aJ鹕+mWUL�lh��Ę':*�jݤ�1��j���
���6�x%�T�@�Q��Uy6�%��ٚdu��f9�p�Sq~�h6��������r���ywen���k=��>W�=@%Ǧ��<͆3���ċx+{��6^�t2�����SM9�ǈK�K]�ux�°<0�%�P;��ЅJ�yyx�u���CX22�Ϋ�G�Y؃�anqO5WhX���������RtZd��쾥�.�5��Q����*��=:�%-V4�ƫs"�l�[��o+��W���19{wա�Yo0���,���t�{����w��֊ *�2������_濚����W���0�)T&$��IE!*!�NGRFRn#&AF� �?�vh"T5�!��bNS�8!�A@j@�A9�7A����@��&"��H�(��,6�<j�a�b�#�@�(�%�Z�F��SNPEaH�H�)E�Y	�bh�a��5J����p��Bq�x
�D�N1|1��BB`�M�D&8�(�P#�R���zx��:�X$�� ��I$Jr"��"�g�&Kd2B"�($���qB�1&cp�L�����H�"!Ȕ�V�Ю4�h�������+��%��Ɋ;��S��S6��XL��������M�3a��5���w���:���^��u�+����擎�Q�V��\�Z��ed�ǋ8��r�[ݰ-��x���A�A���F#��b��w�R�xem�E�%󍯓Z��K���wN���]�v0����6����M�z�`��̜�0�B���"k6����88-u������TqTI�)Mq����}�^R��j`J�H�e�4��yXo&� qIc4@|�L�=��'O���F�ݵ�;J��o@S�'��-ۚ+;-l �}x ��r���Z���b���*��\�_&���.];�:�Yʇ�CU#��t���]�v�g#�A����jgl��#�F�Ij�EVZ�$���936͍-=���k68nnP�2�ЃZ<*�uض��v��Re>�\�+���jӽy�[wwzcO,�ә̋�>�Var�YglQ���J�-)����Į���/�<�:�������R���y]$Ũ*ý|wc�����e�-�N�^(�]}Q�u��׃{jl������E�ۥ�����,sݭ�6r�uc���j�쌙I QJE��b"؍. �	�m�����R�!�E�\.(��qHD.�
1��i�`�Xm�M
"&#1ƚ��s� �B4�,(�h'( (��A�
��,*��Nq�`RA
��2���x�F4�eF��$6\�D�\���I)�I8�0����-QL��4$̑#\d8R	3 pEP�A3.r�-�0Ah	2�bW;$F�Be���#12�i"l�8�p0ZR8Y`E!0"�"E�R��È@�!Ĝ,6�%���BPFc�5�)h%!`�Xm�M>4ˁq��B�R�n���!2
��p!!q LH�Z\�!@��q�n"��ĠP0�(Ba,�c(6�����p�e4 -"J�h�&D�r3D���&YE��+�H���BLe��Rr")�2@�*��A2�I�̑#P��h1@�2�c%�H���J�E"R����JEȂ,��F6���J�#)�K)�r8T�@Y�I
'�,2��
�� A�N{��h��sX	�Q�}�G��Rouқ���J�&U�U*�o������8�ׯ^�q�Nݷ�B7�H����S��r܌SNQs0���B2�{��o��o���8�8�8���N;i۶k7#��{���˦�qs�0��5�S��뢄��J�.�ddf���1�8�8�ׯ]8��n�@��!����d]˹2wPt�N�竤M��ط�{�&ɦGҡ�ې�v�c�ǽsy�Hwu�M�.��/q�u��=��7���Ww��u�;�ww:��q��Nt�w��m�s��[��9�q�\���t�w\�V{�z������y^�����.;���  ��%��S�����d�Qa܄�wk\������k�Ik|w���[��ξ'��V��w�yys�BE�޽z��:��=��T#~��ξt�s���ִ�R��unώzt�qȹs����o^9��{P��Y�˻N圝�����5�U��O�p�6 oK�4�� I)"�wwu�;�[�^��$�r.O�����N��-9�Ww9ֺ{�z�w\��z{����x����vs�׳N��HR �,[o���lG�+�������O���_?��ڎOC/��@)��<)q��^�e�E�w]�ԣ�W���t��]��"�z�'�u,2���I m�	q9q��f�pNI)��$Si��'�D!�8Xn�Qx'֞��E;���UT��ZG3Ow����`�ح�hKჃ��M"q�wd�g������Rl6���!�@��$H�)��&BP���@��6I�(FHɑ�8\|�6�eH�@m�$�[.5r���R&�|���|��<� ��<t����ݙ�<#���h�p�Ӭ�ZP�]W\�h%E]�04E�vW/>f�<��v�	�1o�,�22i�ł�2���;{vO��=3�;���z^{
��+��|��8�|>@���]uX���5[�}��� V9��s_�~��|�f��n󙪫y׷�'cg��ȷg��Z��&(�˶���40˖N[Q|/Z��]o}�("M��W��f�z��>�}OB��>�����6�W�%��W3��u������瞞�{�k�@b�������V�̺�����}�^��g��w�X�z�
�C��5�S^͏�}�6u�$��ї�Ŝ>6��O7��^�4|ޏO�l\��PW�e�ހ�o�S���{Y,��D!�~�t��޸��B���9����|g�i�gy�����s�93Z8�����1A���2��b8��=���o'��� ��9=P�]�"pe�Hvr���j�l� ��	����mЖ��9�5�U�R�{gn;�o�>��x��D���x�~B�������K�en��x��Ѯ�:m�'��W���st������ʰ�v]YnTr^��7N){��[���T<<<=w�w"��z��S����y؟�eR��7�2�4�/p��[b�`��U��T�8�܃=���	���{!����>�o�\�ɾ�WWN��-A��̪��T�������!����|�@��hZ�����L�x�0EU���A�7�^O��w}Wc�kA[��ש�ch�|U��,���Q]����8���{�犽{ Leh�5��fGM�^v)��z�c�e����_���U���	گmsz�G9��d>���I�:S�*w��i6�:����eȩp2�B0јr�������}y}�y�l�~�����V3������y��آr'':o��;L�d�Oذ0wU�8�V�F�}�@\��Ih�l[Oh��<G�:�����'O5�F�I�L-�܏}�0@h�5�V�e�T�uߡ��mYS yJ\;�r}���J�!�&�&�%U��o�2ǫT��Z��)��}����bĜE�����(>�YW�z���E���Nn��5k�nF�1rtz��^*��c	Gw��9��Q$מ���[����c��a�|{<�Ne�9�)�|^�����\b��������� �)�N�U�~����rv�FXz耏i�Iw's�Ҿ���b���t>�Wӑ{T���ԧsϦ�����x�x�@��f7�Y�-c@�>Uc����z��{_TΆ������a�o�ΩI(�~���{#�ݵ�a�����XG>_p��Y��l�/���T�a�;=<v�'FO5S���{Ѝ�${����k��G��ܼ�}����7��gL����=�I�x�E�~��=Þ��Y�3y<�`P��v������[��@�Ͻ�6[���'�J��n^�y��L�I�&ﶏcr7��D����~�[)ϳX��,vgj�<��Z��x����d��b�U�]�����jhw1�]A6lua_t���;��C���K)����ާ;4b<�uq��%tGFUϹ8RYiǶ�(�ɨ3r��ҢE��]j5�%�>�Ub�n������]O��;�s���I�a�q���u���֏+��ڤ��� ;3y�˝\9�z=c3iLs�v>=�o�.
o�=�ڣ
7Z���ۮ�W���s��k�fR�~���nP�&�u0��wڼ;�w,*x���1����'N�5s>�o����.���ޞ~���[���y7��x��wq�7�l�w�"q�v��������'��z��x�_�|�c/�{��i��Q�l˗���|"�٠g�deu��7a��W��VϷ �܎���U��.��zN晴�0Ƕ�Q'XϪ-�[\C�L��țى�ƭ��<��t��0��׏W���>��_�UF��)�Z��t�`��ަ�a�G��;�S3��������og�_����5�t��c��rʫ����ҍM;�h��G�� ��{س�黵�F��t��A5�8��Uw�&�a���B��]�+�[��6�M��W�p��>����$SCVu�1�r�J�b�ܨ��)U��
�����u�o$����7�y�Mm_Rͽ������Yp�3'�[X��rT=�S���s56t9��p۾Zp8<(
ڬ���
�)'�g>!;F�&<�qU~��w�:V�ͣ6�ÛE�1�țEo ���,��+��"�t#�#_�����}���[;��UVz��j*ﾄ�Y�EgR�>9���b����5�M��*��7]7�3���5~������+����U^�u}�b�v�.v4$5����Jϧ���*�w�[S��hce��蠺�4�C�ٰ�[�E,���ڎo��M_�vT�]>�/Ӵ�y,ta9џ���9����ܡ;0&z8�����L���n\4���ී��r����@�x�~i �l7mH 魠\�Dt���;�;k\�"������l�W#�=�{����A����{{p��Xw��Y|r�>�W&�f���ۏ��Y�%y����gd��_L���7��4wyv��ϴ_�<����	���Q��뷑� C=@���a6��3�k�TWC�]JY�J�Fڊ���J��5c��hS�=R�g��1�/^�|~��/���k�slz��@#��������(Gt�d9�cM��(�ݥ%���+n����j��]�˄GAr��p^�éYs04Zn�h�xxxxx{v���p�4����7�o���D����o\����u؅|�ԫkW�.�6ݯ�j�D�2t=����|���.Ym��9���-�(1g��קm%@��o��h�|w:}y`r��ݲ�|KhffӖ`޷v����z{:��e{�2�
�=����|���^�������>��Z���w���v�ސe�'~������..�K��+��3���O^�s�e����_t��LN�l`�� E�����c��k����d]i�z++Jm]Y0G=�����(��raa7օ�7CƸ�Pj���}:�,Ϭw��]��U�vmy�h�}��M�Kg| ߢ܅�{W��_�o~�+0������p�|�|������<���io}M��0�m.��:Y�}�13���sǴ�q��z���2��.��rw�}�q��ނ	krZ����S�A���X�e�7J�����*��دy����&�e}��Q!Q����Cbo.�KۜO_�,��u�{��S���L�Uٱ�lt��EG��
�x��;����'޿���I���O��@��
�[#O��+ޓ���6/:�M�����e�`�8����b�V0��{�=��@ =�j����ɨ�[�/8c�����T��Ww����z��;�>�b�,�Y���z��s<����O��#x<u��l�q��$�U��5�j���9㭯^oD{\�g9���>~��Q�,M,������h�-�'�&`�S�^��`��_p�yܶ���\6G�♟�ՙ�^zý-d��{q���E�lF�g��
��f�`�}�����U�0���%y�76�d=e�3C��m`��;�Y��7��cM��~���=�^��jp[��a�=�$��U�� �M������r?w}��fP���ְ �oܨ{��NX�h0_�a�]�ydj �˚�l~��~�/�!a1���S��k��mvR�z�/�]�\Q
l��\�g.�=������2���Q���NȭuotVK;9��'�~��/.�j�W ��B�p1��-�x54 k2jȥ�Z�R��7�`s-�{�%��*6���Gϱ��/@>����^��VtS4�
����!��}�_`ν��N�u�o{��D�xǖo��V��,Y�s�s ��ڞWa[����y�u~8�^}�&D�������&�]�嫻��fc��[�A��j^��5��Y*b��M$���z�oS�Fx��/�=� l	/���Q�W���q�n��ڗj-1:�T�O�}�K��>|3{���:K���[�u�>�����[=���wzۿZU��#�f{8M�IM����_z{*@RI'�'��:t���p��������57g�C�ѻk��X	�ףO��M~�-� ��>�|D	�>�:��f��z��m&5��6��7���y��rx_��eъ��[����g��p�V�ɏlʿp��p�s"��S�6��/�5M[W����U�îk���{���������d�U�)ۏ,;������z�k�ˬάЫdrw0VS�;k%Goj�BŎ<�"i�at�H �	�� I$�U%$�et�k3^i��5�W]Ji."�N���_ZΪ�Dհ�Bj�\��\{�6��u��I���^��C��0�F���%�cQ)̊^�oe��g0�U��[[Z�2�Z�SE�f�j���l��l����CEyϯ�s�N�;\[�E��de6��ˀ��k9�R��'������&i��޻�ww�������W�3�yoK�]\�xL����� �z=S^���]�'y_�voý���Q�8f�L_����� $D��$`-^�4"7g��j�>����c�.\�zN�u�}�}�~�0B(�3}N������7�ʥ립;�5�'����;�jZ�Hn�=�u��(�{�d1-~�ǰ��lz���J�]��R߸8�;�ә>㾣C	ﰙgܨT�ǝ_z6�/q���wT�g�}GKf���&}��8φ��A���'#�e���O��\���^�bB�������$������J脿*|����h�yt�2T�/��?z��2��b3�3Y�%��x����͋h���uf�����*�: TN�ELI���Qg�m]f��Pn�� Y[�0i�۟h�Y�Z�����f�joٗ��GLxw5����$o Qf,���8����P:�������v3��wë��n_��]�4�9{� � �+63uqn�=K�!��T/e]���>���~��~�m�욄ꖧ&�#��O/\�O,Ī���@�K==�~�����#�.�+��f#�V�K��}�D߆E�&�G9���5>�|�sp+k�\�=]ͻqx�� L�On�����������9YZ�u:�]�݇�>�y�-"����6=/�kN�M�9��b�t�	mO��f�$&���C}s�}d<�P'�*����K��|�&��\�K|���"B^�\޿�u%ٯ�Y<��ݞ!{�̜n�Lp��N�a���Z����]��|�ҩҽn�׽�����{pw�S��v�,�ip�O�c}+x��xhf���(�v����~�-G��\&Zߟ��]��'�v��l+;Y]�_(�IFG���4
����|.������1��^~��8qq�¡ơK�{��Վ����θ�X�uH�+��H���sҋ�eA��t<�ewl:t �*v���.1B�����)��4�q����P;s.�鋍��;)A�/�P�݃$������8�]����pã�GA)�$��[lmy���6��ҥ+.�q�Vԝd�n

ܮk'>�J���ʧ�ֆI��m�YKZF�q�ńր�*5wV�$��M[��y�V-��s�S��ju�nf�X�n�L9ݥ�^�49ٷS��"�&����{�su��w29��7W=��[I�H�V0nV�B�|z�..��˧v�8v���H1]�6�.cL����m��1�l�KU0���qMf��WFMڽZw�e���V�@�!�nԽ��ȳ��&�}�b��f��G:��D9�JY�;'u�����6_"����������K�\6Y��޶�9�KWA�`un]SU�n���}g���|X��򊶭i�G��NwTo��o��j�I��1��`�����e#4ۈ__;�r�iR�D�Gs$�w!�Ov,���s��hno1cQt��ِ
u�v�v�E��t�-���4��0qS%���I"��A���_����c�#ڢl�n��^�j�B��a�(l��.�3�ț%�S[cIi�],B��%_��`+��f2!e=9Wcj>���%Ղ�V'j�x�����*�ɭȱ"�&%�"�O��F�љ�+�OF�Zw�F�i������kFd�w
c��\�6�kOD���K|��	Ua�	[�ɯ/�b��5������	��U�<��yн�{_l�d���:U0'��+��]7c��{{"�2w��̬,C��z�u٢�lt��/��K�bX6V����w�-T{n��q�*1X���d=�]f��7[�T�m�-��V���7�^k���|e��k9�+T\m�X�7Ζ��]K�`��pv�/euEpu<݆y&n��X =i��̮��V\ݢ�7�H���2�I�B;
�� :\�a�mBr��v�S/*߯��ԉκLvf�X��{��8��d�	$Ua���fV3�y4T�^L���t�9-��3l*u�۵��9+�л�3�Z�p�w�"5��!ņ0�T�#�k˖��'2A4Tbt͔�ffC�;�r�.�fN\C6-݁�tʙ��eU�ǯ�Qe�a�R��΅��OOv��gm��Ƥ|�Z[D�;�ʼ�T�d�Һ�źɢ���u�2�I���3FZa����'n��^`��r�˺@�\xw[�h�Z@d�]�f��XBl'ͺ����ElT*�C	cp�r>��=�V��.�*GM]|/��@IZp��A��^���]y���G����w5���%,��{�ە��$I
��<z�����_\q�z�����֟>1ޒ&�jT���)��N9�u3G��A'8!�W�����ׯ>�z�\q�z��������߽�LO�F%��Ɠ2ff�~u����w����3�b��{r�=��|�e����__^=q�����z�������������t���$�uݗ������ȿ����D�����?:�k_WO����A��������r ��{g\���<��z�AK�/NBg.�;��L���{��u��9������^��wuB>+�L�:�N]�t��8��ng]��Jfwb����\��组JL	\�C˹pܝ��wEyėv�gs�i����t��ݦ������z�$�벎����ӎ���1�$d�y��&���& A �SL"
�
��"� ��$�E{���	{��9��K�C{�H����.�˛ :��}+������Ct��]�rw/�u{����)_ϯ��6��]Kl��$�Cu�fU�mvq�5y���=���*����o���
<���%����4M=}i���������;��$���|����O��i���Ǽ���X�}*�4>n��1����6u�[a���`65���A/V����fN5=�� �c�a���9>X� ��ic����/�]7�������"(��^b���s����7	 #�)b�t1� ��h9���.�h��>�ނ�ʶ��%��a]]S�`�i�	��)��e;@W�D�Ӊ�����Z�'&r�x2}'���ɋĨ���F_����V���0�5��yn]���m���MYa.}�)[�U���Yss�{O�/��G�$��GH�O�o{cV��SF�C������]��+�`2��P�]꬇�����ey�czDÙ
�en3Z���vƻ,>��� ���_��j�,���Qu~�>�_��U��`��q6��vg����6���*�_b���<c�s/C��4���b��:T�{J LM�L(^ժ��֮Y/��&�sBi�̔˳7����e�p�5*Jb+����.oO�ҽG�F3G��3@Ĥj㑇1�sJ��<v�%��D^l�:�]�����NP���^�Ӝ3�ǟ��t�G�j�ƴ_)#�Qr|�ِ�E�ٻvm��a��,�N,姥M���w�b]�[c�i�������UW��s^�Y��7Ue�U�w�"�\ͷ�Kb��V>�2�N�0T��ɝ�aX���j�l�~���kD���<,J���\m�����բ����j��馆0b��s9�3���G2��}==|Y��e�ԑ�4ҷ���s��L�z���e�n���=�Dզu7+4� �7��
'=��g�/��o��������f�\@|@�ZN���*���q#o�_K=�4��ü�!��P�:�]��	��Ϭ���zաɡ��~��a��]so��]U���PgB�ۭ�|��2a���Ʃ,n�x��7"�	��sRkZG�r�����L���v[e*�}Η��36 ϶����0�qΌ��Kg�Y�Ԏ�~9L[s �p�Fv�%�{�Oz_I&�����W�����������ixl�x%����$ܵR����3H��#�j �/c�{	��[��c�@�'�!5g|�'s�rT�;�܌Q�S���/tVRx;p���έ��f®�a�q^��TN�c��t�!MQ_�xk��<�Nг�|�{1y9�Ś��k'�6Q|?z��B�	u�WZV�5��/�w������Κҵ�� {!��W��ߢ�5�@���3�π'2�d���dJ��fԧ6��o��X���t�5��`�;���3��iw�A�:�:$�6h�����r�[X5B�^osJ�a�Zëf�1s����ۡZ�;�/�]T.����4�jT���(��ǰz�2�����t�[r%�ȸZ��6�jAM����j��W]z-�C�����/0�n_GD��q��p�8xxx���˨޷���Ϯ螰�;�c��;��,��\��*m���±�[[lP�!XV'W��	�+�!�8��*��WO�?tV�|V&8�/���nO�jSx����뭓P>�Fo���� +#�����'��RpE�`Tc����p�I��o��]1"�B��`f{��.�W��n������K]K���ps۵8/\�B�?�˦?�����C��^廃����Cb�+.�3O�z|okrym�Ԓ�����	��u!q0��e��KA<����=�g�?Ee�x%{������)��q~*Sתy��T�qA��d	s%Ĉ�/�Lx%i^��pC�^S��"�qpMG�sx%��J;��(kΚ�ěB�f��zO�j�RG%�/�Bb1û�潞���a2*�I.�j ��' ��q|
��kLk;�S"�0�ۦ[��(x3 ���^�oC0f���v�����E�0��J�Y3�q^����K��]Plsz1v�4�+8���}:h��`g���(u�� t����>0?�H�|�ѥW�+#!��Q����Ģ=���<#Mʇw��p��š}�e
�z�ʢ=@t�R���Nѝ��	І���+��|��t���ge�����u	��̣D㉱�IX��9�b��Zeή�B�wQJǰ- ��"G�x��v�r����9��#��vjs��c[&�l��k&0xc�]ǅs�٠�|%eA��`�c�g��;��]�J��
�9Zu������T��#�� �3�e�v��#�
#�p;E��Lt�aQ%�w�p|y�^���h�_j�w��Ct��/��36Y*���sI(�폏�>��v;gF2�%����/e����W��M��5�eXL�`�Y�P�>Ntͻ�<�7Pâo2��l1=ܹx.�9���WHU��di�N��O��߂�w�d&TNW�c�B��Zv��d�����Ap������v6�1+ XJ͓��8�"n|�/�s�_��}�>@eglY��R��q.�� ���h�k{�^P��:[]:��)ƻ�M,�kC̟�=y��V�{�L;��M��X�cm�fgi,[,%29�UM��<��ec
*3&�uqN�ᦤ]�������Fjq6��j^��a�Eg�
&(�4L5(�2n��Um�jq��n��`.-�Y�bsVfV|�Ǔ��1eW �_t��2��4q�.�}�����h#@,~k��әY���n:��v�{�Myxxj�c�b7��S�▙���0FD����p9��x�
�=[��@�Һ�?%�@^���Î��ly��nWW/��}t����������c1>���J8���i�Mjj9�6��g�l�W�Rm���Z�q�{��9��b��ۡ���"
q�B{K%��\�<�w�w���o����`�0M���]������g�T�?1�ºG��zB<G�66s/�C+�4�\ޱ���ʬ��;v]6u���+�C�7^BS�g�s�1�CA����0�~����QC�����\>��ސf�//e��h� }�l@��<�#���5�KT� ���cc����??z���L �i��G]�&.&���e�Zj2�5�Bi<��:�f�c� ?+z3K�0pG�6��{E��5f�6��F�)��v�*�qY}���(�g:�]������?BX�*k`#^�G^u-3f�bP�n:���G2���1��IO�w�'����L|g7K �K��j�a��Uk�[F���9ռ��Og�z�e��2STw�;9�����0O�ȝPC)q�c�r_j������ϻ�0)�]=]�H�2g��4GM��ȼ�C��Dv{Ӊv/ky�~R���^�i5WPE��>�s�x��lt��m�� �;<mi�_ǈ�=_z
<�lQ��iz�:���G,���p* �����(Ĳc`q˻`7�Z�����e]|g,�T����^븭S�e9K���0�_<��{ς�Dv�/ʶ��im�R�ۏ�}wYh�H �y`@ū�ukI�nc�-�:�=YF�]u��}��]o,�Tō�pHpp)�@��-�ܾ��E�w-�yt8��n��c#1��^��7�	���>wBkos�x�z�Lu�֢���@���R����X0Z�J��#�q�[y���nz���x	o.���tc�-�4zLcO�s�*@�.��%8���^׭V7��7=*�*�0��{� ����W��7�v����]<�x���,�zK���<�[O��;�>d��C�haL�G,��K�k/i7S�R{�R�D�ལ|�t��:(�0�>5��Q��-�F���܄#I���3�olW�m����1��cO��3j`��7듄��J��_�g�m{�{��>�<��2f���H�`/����!��?�����%mw�y7۩_����l_ �]�F[�y�;0
�}���y�Wf����n{���r����{)Z���Z�V��%b�.�|}~}�-�2oa�x��dϓ����y�kIw�۱���-��H=B��H�ũ@p|�<���kO��
$�Mx���Y���-��-��N*�dOwzM��PXm����e+�׌ZA3��<9o
x�]�jC�lMk�E������G�ɲ�~�}�������C�S?��Z�oLLVѾ�$��))���B5�j.�cr=��܍l�C��<���D�kS������h�$;M
�e]�6h���]=��Ѧﴃa��~oh�ݑ-�Z��й������=�4c(���P�H������v�ߟ'���;��I��p�ہ�Fk�9v���u����D7� ��b�wc���������������ZϠrzt�,� ���~����h�sI�w�,"���xfn����1y%��O���if��wy8�θ�<���@^yK��|s)�9n;Cg��c�`\W��6]�����>���83��<�7'ܪc];�z�(��Ŏ�0 �[p��b8�m�.7��l5ž��t1N�(O���1�6ܱ�s>f�5V7�6+�����t�i��m��`�.^˻R�g,O�ο��KRp
}޼ݠ3���t�{1�낼���Q�:���M��W(��!�-�;L0B�W,%��6���.�Ĺ��񭎟u	�hMt��N���T�g�J��V�_��՜�(G��̾[��SxS�����
?���ZrӸO�Y�򺻜)��2�q�@�"��S.~Ĥ{���Gv����x�z�%e��zصB��Y����~�Ӈ�nf��l���
���i0�r�\;�I>���*}��A��Bqc��.Xlۅ1=_o�S���&�{`#�E�B��iN�y�I7�e��<�65 �;�&�4v��C�Եu���2�l�6�^OZ���k-�Jq���;ƌ������Sy�(���<����z�8H����_i>��>/w,��q�����yW�z*dZ,���@��4-��}��eKH�L=@����s|���ܜ��!��;cLi���cH��=��K���k�`2���Gs��m�4Z�AN�i
�c\
��2ʒ��"���f��?o�F�}h�y9	¾<�_K��rz�YLVW7��1��; E��SA��u��&�yx�qS,�+������_|���sЂ�� �Qw�	��� >5�\��Q��b�Tg����hM߸x�!���{�J���~��@�������^����D|�FV
�|�j�1޾�|�o��~�H���>�t;���h믍��Z���^�z<����E��������t��=-�ʸ;�k��`"�W�]5����ty�X��m���Ŵ'L����$mv�]��l�گo�m��h9F�x<[��	N�n�W�.l�Q��z	oh�G��I�\8xjy���<)�F����.�G�0�=�%�4s���d�: +��t? ����������u0.��a�D�^"�v��h˔[_�����d�:6І��7��r��*'ʭ���bU���&㮶�[x�oc1t9D��Sl=�Uֵ�و{f`:J�RH���*�>c��k�����^cf#7��n��̚q]02�/k}��/]�Tp-Xv�Y�Ѣ�hv�W5��y���k���+<�d��78TC�,S^�ɫ2&A���x��|"O�����oL��(�B�<,ӱ%��DU��S��F>o;:�<�u�U��x�x�cJF�ңL�}���}�=�G�% ���ZxD�� glo�L[ɯ9M�Z�c[��``����لz���Tm11�\[�
�[�	x�e�~]�,.�=OEL-b�1:�����e��!���e�z��y.�O/sk'�x?�cK��]�^�z�PT��F��Ns!9mJ�4�-�����8�^����M@�^h2���qQh�=4 /���,�;�����g�Ƚ�ͫ��O�( �pFZ�sX�@�Bj��0yT��2$�����^;��99w�'(~�����r���^d��oA�M��ü���>,��|�d���Q ��(�ШQ����t�^[�dgM+����T��i��K�c��!��F���[�� F�� S]��f��qm��C�g�d������N����t�������˵�9go_��W3c-i�� z��x�g�qX�J��wn�h+�v���5����s�B�O����7Pm����]�\�Q���S>1;�[���m�Vk~�~� X�{�����p�9=�@c]8EF367����R��fxk�L�=m;���qz��k��7Gʾ�Mͱ)�x{��Z&[���8��kZ�����z��L���R�l��7����Ae���E����V+�+�8d޼k]���ݧ��8���y�Ts9�J�s+Vw}��vyW�;]����P�}c@44M��׷滏ϟ<�����U;.֖�O�$�����?Ր7��^�wj�3���K��[��6:��^��kAv�wY�4�!�׸�Br�3ohvp�*Q�0;~�@J|�
w�Cus֌(���Т�"c��so3"C�G���6<H��,���Q-���0Ó�D� ;�w��!ʑT"�SY࡜Vc������|7�AP#ݑL��d�����[
YB�E7���pˢ]�mR��)sf
���	�;�
��9��'è� �Z���CqM��,����M�� ʠ5���[���ֵs��̺s׮��6.hҠ���+�_|�:$�:n劋��Ok/��)�u��/�p��R��>����Sura]8b�>7��'۸�f��@f�RS�M�I�Z�sy��\�-y\�x��{����^�~9c?v�9���f�ny��Z<S&��ٔ�Ƣ�%�f{�Ex5�:������}l�Q��v�ce�kj�oc��}��K���p�(N�w\�W��n��,�t�~�,������u�34���n�Ur��V�WbD����;^��V��R���fw/�^�Cqo<�i�2� �(N��C�Җ�<�~�����}�@ݱium`�ʵ�,��f�X.��ln��'��= ���̕Ý"7�O�Lc!�V�/�P��S����+�9FC��댎��=�˧E�*gEG
���g�p��B�rT��R)�Sq��B��}�T���D��nL]��޻��:o�u��.�����37eΥ��N���yi)�1�5� �RgWˍ-�Ԧ��ܖ�r�<9�r�(;U����c&�y����7X���!�t��U��RCY�eVՠMAصv�`���[��u���͕=�o��P��.|t�t]�۔-�c���d�%o<�eK�����?n�	OJ�B����|�����+�y�Y�w�B�u���g�r����&�T��k�q<֪ss���0�(]���X��*W�s��,Z�F�,��T,����)C%���yyl=��v-x6ݨ�OES-�x�kIq5�V\q�Up�n�f�L1����N�(pI�2AŽ�d��r�� *WS�"��E���dY.�ȧM��uv�v�/_\Ѽ�s�_##��z�ܷ�Mۗ�<���
�j磒�_0vv�ldBEi�IX}�*�a��˰���k�_Xc6�ǵ�1{!#.υ-��Q]���5C��$`��I���:d&.f{x�yM������7�,�f��;��fAD�� ��"�����q霑��&U��/\�b����(Y/�Z����3�pk&eV�T�RUg;2Y�a�vV��e�R���A�A?j�Ox���T�#�Sq������������ħ�����4����6awv7�{tk�㚹^�c��V�[�-7�okʻ��"���2r��>����倫֝��7W�ڪ�jv5)��;$V3&\}ì���T�H.س&1�R_f�԰F�����O�u��ݚ�8пr�3� ]mۗK��ʢ�=�F|�2�h�g,Й�w9m���T�oP'��M�i�ouk=v�ÒK��k�Vus9����a��%�j��ұy|r��N��#���A�5�ա�S���)��[��9ێ_	���R��3�������7n\�.A;)K�Cl=o���B��@n��+�s��U�]�q��� t�.�2	.XEX�[��,�R�Է�Vv],1��̕�3N\�h���!�����m�h�xkE�bCۇ_=X�m5��>-F��t��YYGp|������2
�[�?�q��ʕ�z��:�U�6g�G���Bm{N3��ы��\�@�:ȳ�����!���5RsstE���H�+���.�B��j{`�B��#�jtuݚ�:�M��%K��7�_\���R����FK�MV~|$aH�u�û����^�#����ni�K�'j�]���Uz�ǯ_^=q������ׯ^<q������n���Cr�F�!n���J�������w�D���� }���߻�w��ǯ���������ǎ>��>>6�TQ%�;|]��ə_wq:�&F�v�	/ּ���Bi��_]<x㍸�����8��������x���Q&,#!0H��?�;Й$��RH�ޮ'�J$F2��?�� Dώ����В5��Q"M �&S�۔$~w>�fI����H���fIJ!|qAa�H$���0�t�)KI_]�&c4D��R���Sѐ�%���&)�b1�_��;�G��L��$���Xf�LQ��v��v	#�0���1��@E�A�B`2���Abe���J�,���Í�o��T(0�B�n2��֌�Z��p���Tw������N�v�j�Lh���	���3��42l��	r��1`��a:�U*S��M�T�j4�$Ƹ�-�Y.I����&�I��%��8�*G� E(���H�"jr"�E|!��'��R�BJ�A#%��2B�D���(���j^��z���[�iD���hi)"��ó�I_=��y�ך�,��o7#�̑��eJ� [���G3�+����֚�S�V)��͂���{��ք��;>�&@�r����Y��t��-�c�oc����4�h�t�C�4c�w��*�\�b���Q��N;aNl@af�U��Mm�tW�IQ�d��q[E?��E��>��kh\x���j
r��~Y���=��}�f��$�<]zF&�{��0q5���gu0~><�h� }/Ӕ��6�{�f�4����|�ffg� cރ4����h�RZ�`�@Ɣ�˿e&0���~�� �Cݝ<�9�b�$g.L;،��/�K�7�y0���	���d�}�7��~���|�P�LW�S;53njHƦ>s�4��]���G;�]��`��@�TH��t�3�iZ|EUZ�j����m������Y�X��n�P�br���F_�y2��; &Vț�j�aL����43y��7�����&��唍{�YϨ���1-U� ���m��<���c�M���:�N�1�F;kb�7��r����V�{��Ⱦ����K��m;(�NY�ҧ�lG��q�
�Y9�������*�~m���_x�M��o�n�ԇ�Uݐ�+�`)�-v�2ȹ�����oyv!!r�zbO�ﻅP��=B�U��j�Q��h9��,̺�9]�rm�\��} �;}A=A��<2sVCǻv.�!	��ն9{�U	� ~��ZhiD)��@�WZc�:K�=>��0=��k<����a�߁Y/���)��½���Λ����f�*5s(k��)�c�y��2&0�x� K׉�e�ؔ�u#t#ۦ�.#�l�%f�k��?�W��u�#���߶�*-�d^�,�#L���qr�	��`6�p�顔d\��k��\�E�s�溂'ֵ�ط��d���=��
/��$�36,,6�x��Xby��lSk ^mFGh{M"�O��o��Z�0��[���������uG��[���_�g�[��c��M��0VZ�j�������$��ɰ/�>Y�P����ެEP���W0�ʋY*S��CD1o�yz��0jn�þP�@��{�w��x��yЛ�D�q,��SL��{f�9�pq�N�������̸�Ba��w�;kx����z0�u
c��nuG^�Uzh��4idS���ŵ^�4�
k�q���F�P+(�\�<�xg�T"���Z	�:e�V�kP�/?CV|��q���G=��I�T=򃮅�ߝ�X�v@�-�/�=w�	��e��R��a�[�鬣����h�l#W(�1)��\�Ff/�
7�����03:#�I#�*vj��+�ț�l�k��N�eu !F�nΖ]��xd������D,�y	�Rӷ�z�x��$�Auw��F�}"��j��J����Q��"�V��䙟>H�|�W�UΌ\~�z�5=u�:���%׊?���pi�3w<�{�;y�No���z�o�=*����s��q���X��ha��S�������o�=��8*na��C��{}�L\��� 2��a��ٟ4!���a�;-��-S���k�;KV�ؼK� U�Mޖ󎴷,]�ݨ�d�=��<�Ԩٍg�����z����!$_pG��F������N��]�ޏ �|�E����S��-��8j/_��1\����fE�jqx'qm�}o���'�B0y�K��)��Ul20������}M����e٨E�ǆ�M�ǝ��5,�s�A�npE�O�Ωs�~3ƽ�zkG7i���9z�U�R�h;[��_3�H/�#���p�b��c��Of���F����݈�=^��7V�0Q���8�~�L{{]�>:�<�/](��Ҹc^ f��S=��pm�x�rG���3�o!�8<����N�y���L���|��g `���$ �\?8	�_U�|��ˌ�n?���q�hh���������ea|���2]q����]�#�'ڽ�!�~
F5<�A���M|鐪����\6$�c��؈	(�E,���,���;�m�tU.͚AU�q��%[x�.��W{�E�����8�844"��
��w����S��'�?\���^����9W��7���@ ��G�0-�'���c�?
�]�Ŏ��ˀ��c�^Ǯy���!�8�~���:)�n����U ��E�}: ��vSͳ�s}�Cp��Ѱ�`T����62]�4�l
lm؎/Ǡl�́^/��E���Q�;�k�2���TC��&OX]p� �NUi�I�������ED�W��`ןH,���6>���CX���s��|���Tޯj���%�
�L�/;;��W %����wþ��NϹ;co�v���6i�on4�q�~T5���LQ[f���R�)�g�c�C�l��{��wf\���G�d�(�fO^&%�U˷��."$s҈��cc��U���<�$Hc
�Od��	c8ǡ\@<��-�n`&�%�VU6��敓7>��ܞ����>�4�#Ν��T�/ /;�qU�#�FLxl�k·�,q�֢�z�R-����5�lrd��3����Y�+�e�0��٧�Ag� ��ӌ1?S��R��LL��nڝ��m�(��d�����̳T�^D{�S���w�5����<.��Ԙ����L�WeMf�_����͗w@�<B���"�
K�%�aɼ��FS�h%��v�7�Z�)��S��Nf��u�ao��R���Qi��z����x����
�44��PD9�pЀ��n��ѥ���5Y�g0����ԉ"�����55Z�i�g]�{���䈯�7��>4=�����%d_�>��}� 3WG�5��׍��~�1P�4� ����gD����H��n���Z�~��+�L|��1C��On-l�Y9����XB�r��0��Aq�!�f4������cH{���<�6m�W�sD�xx0���m��C,���}|��B��s�ː5�ZFK%�0ޟ,g�����;��M��z�=���f8D�B��^O-�]-7�7�M�a}���)���;͖�Qh-�f��_�M��D���q+F������E�p��ū��I�}����;����zE4�Q�1�7�ʁ�R�4|�s:���MD$�`�6����[k��ô�9/���N;�:�Ćɭ�h^���w�﨑9�j�d��a�aw���Ǐ������oW���=��Fc�2r�&]��	xm�~.K��_�����~]-,�q1���ON�/�r<3a��f\�*l�\�SS8�Q����현S��@��{���:�iwiU�N
��)=�w��S�	c&.#'4wl<]�J���ãrLx'��\�w��x<�X�BslF�̏~�z��Y���_������M~d����V��mA�֞�Ԇ[�9~Us���ˏ4�+��V?C@M*44�h��ˬτ��#���Ty�}���a�k�v��1��%��ͻy�}�nUK�)1��y�乞>�*���(E���D>}�F΃�)`�<}{ �;4����9��=������ݞ�䦋�N���\�5CS��*塸W�:/�?�}t�[�U�{���B�8�$����#ɦҢ��^-�"r���g�."~�����^�?�D��S;Я�d7�Gs�1�ykؽz����wV�bB�a��4�M���:�?�;��툰�\3.�;^��rz&)�?ޥ~-a���U��C�\�5�5���q��Fh>��e6TVt<��LEQ�,Yy��1����2�O��Kq|��cT�m�c�O�a88x�;��w������k�,]|4_�On/��y�FD�b�K�&�zy�%�4�<s0j�:�!�+�YFSS!n�a�d�u��B_$�*z��X��b��
��x��ل���Z�B:["�lM�7��u����Zc[vn�����4������}zx��K�}���3��hX<�]p�v�9��<͝#b�Lyj�ә�<��@���k�����W�L���4���YvqNu�Pt�V;/}�hm��E�}[$��w9���Xv�u'��MԐ�z�h_7RSj�a���ڗۮ�O���4(��SCH�Ƞ���ϙ�V��̮ʔJל���v2(Z�g��CZx�1j��C��n0�a0����A��"��$����1���-;ѭ����Ba��6v�>�`r��%��?nc�t��}-2mi��,+?A{:bB�:��U����j.ZY�g�d՚`2T����az�i���8��E걄>=��J�e��ʍ��]Ƈߝ��+�6SȾ;��t��wnE +�o�*^I����P*j,�^8��-�;F-��cPX�8��w3ʟb��fB��6�w����u�]CmX} S`}�&����F�Ը-SQM�T��f����廮��S��D�{-))�A��^�,h��!i�Y���1o���B�c~�wش�_|.������� c%暶=���=�XV7��U勰/�C�Ւ̹٫�魢�Fξ銰Q5�z��p��P@��u��^D9�WlS���A�+QQy0*񢓩�o^K��*Λ�C�P#VH�p[-�7O��D����L&��7v%]�w�S���!fL2�C4���e�vʝcgbXt8���|'�xU9�G[v*ٲ�ځV=�{	+e�\�d/]���/�ϭ�0���4�5��&�*���kw'J�n�Hv��۹j�a��Co��9)�R�L��}F�c�̺��>��#�p|hhQ)��T^��e�>|fs�n/�C��W�PS�᧡�j����O�ީR�G��^S�*���td�
�r���e�3��Lh=���� LG���qAi��u�����<}~q�b�����5sn�t��j�u������6�@*-���L��e����5���2'�)��Cm{��y�mK2낓\1ЦB<�SK (P��r�P�ycL��6}�s�C2���X]� ��VakQ�팼�iY�f�W�ά+����c|����b�y�63ﮱ����� ������߉�L~�w�]��*�K�N�wӲ���1�-��z9�5�4f6>i��;�v�DVB;��4>���S03��õ�kU�g����\!��n'�@�>Za����KAdNW�E�vB��[��ˀ�ɢ�ٵH̯@�r1p%�sm��~���f�
|0��^,X�~�5
�q�iia%�*�2��vw�;95o�yv�Ԭ�go?m,�mԉ;׉�a�%z�k˼��[_���o��}CM?I���A�9O��/���tA׫�U7rX�X�ǫb������-�����<�ӽʗ^���=,�A��:,Iު�ѪEW�}ѴNb� �3n̥�����`4�zyz��U�|fR�USpd�)��)�y�K(=UU�~��F�ThhQ�w�3U}��C��~�6q;<�'����G)5��e��m�$��I�3cn��Ҩl��1&[�C'}Ͽs�����G���O�_}�J9ck���m�7�;k�����z܀_:�&���܇/FȦ�R7���E4ە�r�f%�+ ��m�%�*��֙pd75�;K�=�����&�~ra��Ǩx�Ct�E��}�_���fҡm��>�O4eU�8y��9��v3.��϶�X�ߝ+<�@����� ��:,{���㤬���roD�w��E���� {�}�KM�F�ǍA�5,��=�O��2}�s�Y�gHf�y�L��v�n4��>�d�TP�Si���F�Om�^�|$��Vh�
����_d�ٍ`:tUa�멣�s�{��~��
�h����x1�.Q}�������(�TE�j�(���O�z~�$�N<67r�^E�����z�)�_�^U��о�~�t{X��};^������bW�z��P>�@��@��E>_|�R�^�W���{sf[S՝��&�4ˋ%,���^�mߟ��^V�@�]�}$j!��K��qZ�޽���"w`\a="�]zme/ՙ<W�N��ObW�sq�sJ��3���O��OFK�V.�g�b�������L9��ΗnǽPx��3)����j��K���Mbllv���p���D+�p즭��֧]��9�{v���/Yݥي�7��z�^�C@M �44��w^|�wZ�������m�g��v|k�2
-"m��$��H[�\C0bhT5����3���Nlg]qg�Ai�N�����rd��0���M�������z�@�>R�g3)��L�_B��WS��(hlFϫ��}#j:'߸���UJb�M	�]�S�ր�gvB9B_�K�(�v�4���O�����P�j
��^I�<�b�Cq��G�9�3��46��i�晣	,�A��H�y���}�-�f@F�Y�3��1�rI�a�o�vm������λB�V2T?z���>�C������s�/���1�҂���:2փ�Sm�~���wvqq]�}}��BbY���$��j0������5��mA�4p7`��0�1Mu� -{���t���Lܛ~�g�1�ɥ�.hw2�:�aSe��Ҧ���瑑�n՟���g��K����j[��4��r���j��mĎ�`�b͎>�D�`�����a�{k2�Y'j/��kFx�����c*����?@�o��1��a��a�̬���q����l����ѿ���ﹽs�}.��o�mA�7�vsР���(6	nf�x�֬t�rf�-�ǉ+5�ҝ��
��;��Ė�&j�&*��*�p������J��Jﶦ� ��Ym:��!u��K<�>��:8��Onb��0mU����d��%8-���ueE/�WAq�
����mJ7϶�(����Y����޴3&̌m3�UX�:�S�܀�h�V�%e��=��W�7�r�s2�i�c�F�S�@�.�M"�R��iv7�T��ӽW��n�=�WV#��]��Dд�:�"�����n0���v�yE���w������p��Ɔ�0����b��+�Um?n>�0]8�r�m�(�n���/������3:-�ī�.��q���n�ކWR��C�{�8,T"�l���W���W�� ��}]�S�"�.Wbe�!��}�P�l4�1̔��-P"�&CZz���ᣮD�)amG*��Ⱥ��V������4�,p��]�pj`�h��q���ڴ2�xx�di��}K	=�a�:`�W7q@kD��a��i�pd�kՈ�u�ol�f����:ħ�P���8���oEh���9��Qͮ�:�v�֩ �LS�50P;+z]�
��,�Ucsn�>�ܥ�s]lT�c����1Z����kKo/���8W'�alTA"-��஖.��hŚ4yV�h:�E��Hm�7�t
$U��<jJ)����!v��P�B�����5i��7#�`D��$JAt4j���]����u�(��ţ&p��1��+�����Wdz.��kٽ��v��UK�88L�Llx)��{���|�_bz�
��t�G7# "�	]����j�'����%A;����=����ͨ���ӆ��[�U�j�.Lj�^�]8#�3��V�k��;�8r�"^%�l��uqǝp�[�{.�清��g!�\�ވ�(X�M���l�ث��;��Z"4X8�x4�����)�I ;GDf�ӻ�'.2�.��t���X]4�W
&�`�ʶ=#�[K,݃C-Ej��e�m_�:�N�8ȹ{E`8�{R�����&��:��)w3�^�˜Uc�5m����2$�F�)�$k��peft��ڬ�46��p��^�=c`���9�腆L4�u2��}Y�6���#k2����7������t.
��ʗF���y8�y���o������'�l�0gX�c���,��E����v/S���tEI*Aud��<������:��Yv��Q��S]�no$f�Y:t��kC�n<Yu:�=c]h�۝�#�Ћ�O�ԭ��t�Ս��\�f��|c�Ε�^�����Ҝ�vc�!�ee��D�r&�u����ٵ��4-w�	�IEp�	 �|WKB/��\�)��p���F��JI���^�|x���q���q�������z� F�"I��^�HĄל�_�s$�B2BI׏��^:|x���q�}q��}}|||n�2)	#!�t~:�]&1F�댌�#�HI�O_\m�Ǯ8��q��8������V1���B7M+3dْ���~.��DJQ1��H��ﷂS#���w	A&f�����|q�7��o�z�+%�\ƙ�A�/���;�]"2Ad�ѡ4_���(&S�WL�3)(�!�&$'�]&��u1����rM�~��A���W��}u��(S`���&Ɖwr��rl���p0Dȿ�w�\PbL�4�?{�)
�1J`<�i�B��8=g���������������.j"������j�l�b���7�!�c2\� �鷯r��w9rrn�����4��A�
�44  H�;����k������ϓP����h�b`�E_*�����)���6�R��n(��V�j�f���D&YT�/�0��44��S��( �3�Ś�\�#�N�&�UgW\�����b����?�IZ�b��I�O�*=�-�K��<\H�=������S�C�s���׊��kLk`.���E3�h��/u1��^YYd��~[01C����T��$�3��߷��w:�<�{�a�z��D7��&�P[�W�Gh6s�Z��y���j�%��ϓ��F�N	�Bjҧ���Ơ"!��6�v׾H3�*#��ՙ8�(���] ~�V"?��`�ܿ<$�n�P�Pw@�i�tX�CC܅b�0Udc�L���l>��v>w�����m��"3:�,3j�_�ƿϦl�Ak��#�����+��2[aS���j�Iy��zGx׾�+�y�5�����G�܍���O���jfk6{���O���;��t��w�Qc�s��L�?�*�W�Ú8
�be�$���M+-ѽ���r��w3jA���8\�7�e<�&ɮ�@�b��Լ�N¿����9-c"�]�I��Ӡ=\�ߡ+DI�~�P�9_-����Ä�ȹ�ϵ�S9W��Q���Qӧ�3�� {�o�� SC@�"*כ�f2&Sϑ��"1�s��¹o@jƑ;덯�+6��l��Y��4��s6�2���{u|>�zs���F�Y�q�*m���,]�[O�g�-ٗ;5���{�%����W]A�q���Q�	��*[�t�Y ϶��
���9L�N{T�u��XM�,�hm-���[��N�H!{PZCONY����'�k�<�L)*��ؕ[r�w9F����Y�������1�5��3�����	���Md�y�ƙ\�%����]P/0�ӓ�ʹ�����@��r�б�zy�_���I�\o�Mg�~��4�������ll�T�.�``#exB�T��Qˬč�)鹴�;Ǆl�|f�t�}XTD&�^nʜj�JִX������KO�u�Qk�aE��أ�@X�<:�=�h3���� ��9�a��uW���5�S���8m�ҍ_G�O>+���;ɖ�a��j��ŪD�lmZ�qi�Z���،d�R'��>������Z�S���������G�{�q�n��q��Ֆ3Ⱦޙ���.�g#�ܙYC+��2��ݹ��_�����"��k�����:7�,��b��\kP�r�fqR��xEV�c���km�._6�ꮾ�:�O�0D)?v]��R�f��מ�3=7^���&`�ҫM �@s����v3����T~�ܦgvv�1D�95��`��v��Pm3�n���wf�c���0*B�/�������,��\���$��O���ZB��n��~|;�vO���F$��Й=ô�W<���'!�C��$��C�.��b���.n�	ׁ̀UĎS|�7����ę�*�39>~)�\[���j�,ˀ
��l�m2�2ii���������Y����~ZI�gV�_[��8au��0o:T�j=R+��༜�|���?/|����흑ٔ�^%�V(��e�V����,���,��"�g�.�
ߝ�/�r����!����
{DxK:��}>�~��	}m3w������n��*� 9�x�_��>�Y��v�6�א)Ek�y���'��OK�?6�;���j�Ƕ���(V�[�����AR-�5�Tc	�(�p�(�C�똺�/8��
�y��,N%B��ol1�G�v���T��w���`�?X� 3QR^�eWRfrt>j~!�vm�tz&-�R|�P�ԍH�J�`�m�c��q���"�,7���ݯ�=��'�k6�|�h��q���qT�:ZO�\V�>�eޝ�5��Wk�q�R�3ygd{�zUKՈQ�n<J�֐w�:�,��Y�v]K��
�*�e;����5xRG]��fu0N]k���=�v�p~ s�~��Zhh���Q,�Ϝ����)������X��&�9�1�$c�G6�r�C�7Cȇ����Q�i�Ǜ�E/^D���e��%�_�Eto=v\�Mi,�9�,g���[|7���{�#�[ ���(zNΘP!�yh.�ת=^�j�2*����П����P9�p\��ӏ��Y{������\��`%d��X+4��crv�hgP��]����u�p��զf�h�����[��ᙶ^���� �|H�>H�Y����[�����4���~Y�����[����~*����:�u�y�(�N��PE`
��n���@j"�7���f�����3��+`O<`XiT�.�П���:kd]�`��^�.��;��d�#ug9^�����|�{ư�=��9�np-���jnl�f�ۤ�4d/Cΐ������Ϩ�������0��?��!�tk:���Q������֎~�O�R��ϫ;,�	�g��[��"ڦ{�DX�����~k�ff��|�t�i-�~ǴD�o�~�Gu^S�$��6�̒i�"��F4{�I�ƴm��:Ce��Ƨ����y��mxv��Uv�4ѾuX5Ն-<�Z8�9]��wr�6��˚!���Xc��r3m�����~f��Ms���>�� ��ЋM
) �/����_<����Uww){J����b�����mn�Z�Vl���:Erod��8�yT�X %�v�j��b[X�7c�1EՌYCJ��k&o�!�p{o_���}ƽ�
fkx�;���,f1��tL�H؂�S�<}���լ��"�=u���5=@OL$^�r�aF�n�gz2�ph����Iξ���ދ��E�(��r�ߍNdB��+�Rx�ߥZ}�޴��_��a�c�̛,���uIn�)��zi�kWv���U۶��
��������Yej����O�՝O���0Y�.(j���=0�<�%��oC�-7�9� �?�j��� 5&H�Ö$F�wt_����5�FO<�������ݭu��x���;�e�T�֩��D��02��_�|�G�^�����5�f��l������2��zFoq���-������ި||H;�
��M��1R���	]��"���/W��@��\p�W���=��7\ߦ�#���7�;w���~�q���t�i��f2���E����A%e.�P�܏zC�2�z{�^�l�R�U��uÜ��Ҽ`�~$,�4��x�lj��OC{�]l��rI�3Ґw�ݻy|�_	��m�,��]B��E37��LŊn��d~ p_>��JhiP����Oy���k覲��_��>,VU'�l>Rh=X�;��tf�ʨ�H�td&�j&�M��=�iM�O��B#��"'�g��)��G�uF��,,mW�@��������'��e�L�����l��Wv���C7�M��#��
Qg"���s$;'m��-�V�M�c�>�@q����d�L�Ao��7�qw���v\񲺷�b�5]�m�,��+����ysJ[>���L�A9B��V���s�]�4��ȳ�lCulH���d��7P�1JSs�lL �5�ǟW@�YKխ�W�.�-����N�G~;Y����t��Ӛ@��%��L�Uy>׼&OH�o��lo��Oc�m��GoX��~TJ�}S8H~��W�����,\C���`�}���sϾ��)*���M�B��f��r��w�-mC��*���|j�k]�}hw��-�~9V��K��g�����!އ���61t�+_Z��g����Zvy�_��`\��c^Xt�����
���6(�J��hq��`6��6�����戱�AL)
��!S���r�6x�z_��t���ex������$ol��;�.�܋=���	�,��v����+}go�.˾��f�m����^gj�'a��/ O�uڣt?����� SCJ4�Ъ�ٯ<��y�>��Uq
줠���o5.��@��������/Ghv�On��Gi�
m����z<��P�k�ڈ�\]H�~Om�>��#�l+��lOH@k���[��]������-�f����5�!�-�ݎ()��� �,i��@f�C[���i��9
��-��#-�?446���5l����d�B�Y�3W��-R+9f����|AF�}�}�AÏ~T"��,g�����!���`��2�|+�6�,�]��%��}�{�����3�����(5���?N����Oa� m�m��kc%�P�M[�u����Ы_<@�2��|g��,����Q7�|�/���\�)�*+�(�\�D����w���O��'1��Ǝ�)�q]0^��ZIG ��ʋ~����z��G驪���(@��i����c�X K{ۏQ�<�V�!�q��4�V��L'^.Ͱ�#�>]$�d��_|�K�����om8�4E03��	�s�x��S2z���W.� ���>���g�;�s�s�t�-�A�n��]0��-|���,X�[K`�B�9wͺOa�Q�#2bb�����s;�g|����Ec���}��[�}�^=j]Ǝ|��.ӳ/v/T�<\p�H�w��]��h�&�[�9�����޲����a��8�u���<�q[�p���K��oe��u��{o�Ҵ��%44"�����>|��9����Li�`��J����[��	�Pdk���,q֙;\j���m��B�����tZ�R)����{m�a����y������Дǚm�c�g+�&�4�wv��qt'F=�v�al�p��+]'1�1V6m�Ma��XsX�s����3�
T�C�d�P�Тo:��\�Y�)��֡�9�1I�p��)��'*�ew].�lT7>d�_3��9����la�W�zc;kh��N���ȐM��9��(���u��0��=}�N.7+Wyǖ���{�k�5�ޘ��u��Ś���z�S&����c����F)v�l���οl��k��R��־���_��(t��}B��H�^�C�ղ��.r
��mn!��X�Z{!�ǧ��2�Nu�P�
9��s��!�|�uW��!�q����q���ۥ��Ů3�����Us�ɰ'`���vk�}.�/�C�V��\:զ�e��\��kU�"ԉ�O��1�=�}M��"�	^|�J����w{�	�%��&=++��+ꩵ���񪖫-�\5&n�b��AaYӵL7X��t<&��P�>���j/�_.|@~�%���OU�U�hgԉ�!7M�u&��G�y+i�۵�#Z��|�ԁ�Oê����};|+7�Q��}#��i���ǜ�z�Nҩ
ަ���9a����o�w�Vcݦ-�Y�~.��25�y�J3�Q,���[=eݢ_Px"���BX��:���-�V0���\�ѕ��Gs�bً�%����F�w�{e|�سF�T.�2���6���"����ؗ�qmB�͙v�r�Ѫc�s-<�Dl���-[�2׆)�@�Y;��D{P&�=8r�_�����'�)��������fgv�f�V}��<��5"@�5V���1d�<��v�g���x0�����
7آ�q�95i�PxT*;�w0��K!ϭ�������Q���T0��v]@4[F�[3�����ފ��s�h�:�հdN���c	��D��+�9d�o��Ð����޽ʜ8ڳ*ti��C	Au췹�r�"��]�'K���4������ɑ�[����ؕ!oOu�5�=������cs�>�g�օ�8�_=D?4�������&w�L;��%��T��ݚ�_"\�m�wa^g��B
��9��$t3������@c�y�dM�����4ܻ�g�ů:�w���lf�)K��xd)��z%�8����P�*e�o\�YJw���$��e�`��ֺѬڀ��,lH���P�6��lB)f>�gU��'ox!�t(���m��+Z�}R��,��V�M�rjф>�6���9�����44�M�'��)�H0�`׋�|Q��a���)�������X>x{Q�A%�����{y��/}F�D[�l�e^u��%w*)��z98����RXH[�{�b�݃�h�~`���9�aת���}A�n�����^Y>�7�>lfs�ӱx`5O��֞1LZ��>�����Z�Kᬶ{37N��\*�t�	����ıg/l������g��2��Ba���=F�8�u�9Zqf�V/�3j/d�O=�Q&+)QC�}�a5�e3u8�]w��K��qZ��2��nG]�^- �3����_�@����P�yt��T����,6.�g�	�S��w��Z]a*G�i�e�}�dl���c����@_�F��b�Qw��Bk�\F����?9Nש�/}�ҋ��!���0vg��߮���I��W��N�;i�rhХ��|ɩ b��z}��d� �	�x��X���n+���W=��f�v��L��n�d��\y�=akVW�HbZӱ|}4�(�
9U��F���=��R�w��8ȣ�#O�de�h�c1%�
�-��WKUC��x��F��WCF�a�w1���Lj V�:��C��&�TC1X�ى4��T�^*��$]���8t�=vb�z�l޷nU�Ŝr.�0��� 
*Μ,ȷ3��e�	���[�e��-QT��b��N��1>w{he�M	-`�&�+wGl�(sh�ҳ`�YS�.�9;����{o(ޙVE��KQ�Nk51�%��on��BV<uu	���y���|/�� �����;�y�<SWE};����Y*Y�y�2��kY�uv�@��NՍ�{����Ȍ���<��0�x�+�����WZz���lsC��'+W}L�y�y��w�S�de뛌��|]�b��'�`Cv��}�\�Ӆ�n��7���R��n+֓�n��p�;gG�1��w��8��l�G���j��R�i��r�u��e�m���mr��+,�xfY�2����t�)�=�F'��Yޝ���)�{��w�a�ܱ���#�z��֨h�R��=t�����˂T��iuc��Zv�KaC�P�yͪ�r�V��w�hm1�T�r���]�!C V!Bf��=��5�H=ϒ'��4���뮈j0�ss�=fƶ4�U,ܥ�H�v�z�E:�g���燞Q�����w4ɒ�hQ���.���}QW/m�{`�WN����&��uF�������^A)�:4u��u������`({��rs�;�����68^��LI���ᩈ�hc���њE9�H:���a����H��(Չo�+��h�ò�+7�u����W��=cK���P=���&M̘g,����7ǂ.�̛��������\]uWPKB�V���vp��ª_h�9С�)L��N��u]dAocՓK��c�km�8���WͱA��_s+�`�� յRL�vmgDv��ꤲJ�f�T�ט�I�P$i��9G�JWY�S%��nM�=�'q�\�H����N����B��k�wA{o��y�i�=Ō��)�LE����j1UyT�QK���d1���B��Օ��Ò�=O2���A��$�=cnt#v�Վt�GkB��A��Z ��X���kr�w#Z#��"�`�+|�Dvid��z�#�^#t��]��,;�Js/(��\���]|n�2	�K!�d�q��c�2�!6���е�\���%
Y�%jI�G���w�4%����XEC�v��8�Ҥٽ�e�(PR!��T����3�_ʙ�b���y�3�:wۀ0'vYR�6���2���S<�wW�<717���v]�n�ö��:�ɌsGNhA�~~�O�� H�6����C?�t��C����|$���^6���:q�z��6�����ךMf���y�2�$�BP�C|�I$� �[��׏��x�:q�z��6�����Ւ��	A�h��la$��U�>7F��K�*#1$$�����x���q�n8�ׯ�8�돏��[$��$�=݈�
Rō���r�h�(b����4b�,/��_�DP�CDF�&��1��\b~S�m��nF�h���KPF�wF���@��cO���BS�F#�IcI``$EL�&
��,d$"�1�Ɍ�{�2������f�H��H�L�KHK��,��Rb���=��+�F5�����k�$0��;�&��b��߫�Q�$���c�|~;�W��mE\���CH��0�c���m2�jGȃ$�X1�RI"ˠ,��X��k��S
']�:6G���2�y
�Xv�=��iN����uP]V�����W�6v�;jU�^�*(Ij4�E���
�I�!�XlG	�@�M�
�"�8�I$�L�a(�&B���,�$I6ʌ" i�!l�f�i�T&&�K�F��6����fU���������CH�C@�}��u��=k�*戋��Ჱ�/��+�o(=�-�[����C
d�zzU�ٳߗ��?��'BfM��_]|�\�S'��循b�m�6Υ��kS;̓uͭ���}dxwϽ�_R�<	�.�c��6� X��Z��M���N���S����KW!����[oi�l�0��4�S�~�h^�fj�L��d<�[�(�3������q�v9�3��R|n/ͽ	R����A0+i��]��X���Y�\wBT܄Ѷ�,�ŦSzn��eO'��N;�uP���5�2��'�}�H��4��խWw�R�DF;���_H��Gg����Gԧ<��ձ�S�X�o�3l\��&�L�t��=l���T"�/���vQ�w�ǵ��_�Y�3T��u���/0���g��тOl�B��~����χ�L|��8_�<��~n�.��K�<���"��V|�����ۜ��+fbY���d��� ��=�-|{����=|8���������gz5�S�� ��8���39U+E�,�ks.��z�H�3%��5ûYǆl�J����b\aP��-��v�_�1dS���fY��h��ff�3���+EW�����L���H�:>�m/��GV��	���QA$D��D��-~��9[�����in��{��jgNͶ���P��ɰ_�ƛ���-%����wA�s���\C� �q���5�#B)�3]�*�V���c�f�,M�_�V��奥��W=��xi�%�Y�ѐϔOWsGi�L[O,�O���сX��H��U����(���vmG��:�x�t��ާ���&�]��a�Y�uNW'�J���;����2zL��;N���U.|��J�H���e�|�Ż�w>}lr�]��B`q{�T����tK��0�l��͒W7.YB����s�oy�o.nC7C�N`�6F�v��(N��e$���5re�u�QE��P��Un硛4][G�@��p�����t؟z	����&6X�C��+����>���!��ӰGF��2
��{�LM�{V�.`�H/@�z�[
§�4�e�]�\�sW��RiyC��G��f��ζ��M�)>�� Z�܍�ȶ�v����"IS���ꃲ�]>2�1i	�Wt<y��"{�Q~,�K����:�A#�ʈ�o��2�^�[:M��ᐇp���f.
g%ᱷ���"�0�M|�׾���M�}��~+�'��[���S�a�:�sr^�bW��/����~�\G^U
W};k�ֺ.��h�N�k������t����c�Cy�f`X���yx�|o/�8���[:-�ý��d}�8�`��Ԭ�W�I�5�����ӝ�������[�Vg9��]I�O���CM44��=���9w�F��)?q"���|�Pa.�qt����_���R�y�&��HŌ!���m�OJu��.���)�z�'� ��OV%D��}��q] ��c�s�\ �B�hL�&��f�0B����{�~�Ͻ&����M$M�>�o;�␃�3���]뵣�G!�]#:��jɏ6�8��5�љ,
��W�D��8�i}J� <F#��E0>��F��ԇLf.Y��yG��5�<qr#ީv]L������p��Z��^[��K��cY�ON����]��P�)��3������&��O�Z�3��J�c����hǛz�4M�k����UZk������4|l����{U*n�0�Z�����ۻ��K��T��3�~c/꬞�^jCv"��o��E��^=�e�;�$�Dz5�y�c\r�f��ۋ& �U���v����_yp.���e�>ݩ+�L<%��,���]��ϛ'��<����X������(my-�n������5��-���=҄�ڿﮄ�÷Y�wfe�JV��Ǵ��pʅ�+������/�Z+��F�j�]��44:���F�����8�@#�$�5�j1J�unη8Pp�v��4v�(o��hu�5�%�(X��>�f����*��e�<ow71Y�����\C��Uo9ұ-�Z�z+е�r�s�Z��,:�tBO����X�~�"}���&Z�FI	<�mƛ��GyL8,�@�0��;�q�<ᛁ@A���rro�L�璟r����dOo^�f|�GOM5F�-���q��5��ݗ��OH�}���4���{�L3��%��<�1���V3�wu�hi���R��B�hg��{�,��m�y ��2����mWl�ݔκ\!���J�d�(\O0�-�m4�I�,��_N�q_?�Vvh�6���w�����ֵ]
��a\\X�0�&~�)���x-l�2��f���,�����.ɠ�Z�ƹ���z���y��L:��/BW���6i�8��0����<~�����{�7�D^꽍���VE���2��<���qB_�xd�����}n~�N3I�l��|y�9ُ�4*�a�+���Ƴ4�3��Nb�4q���ߖ��H�³��:`HQ�g��n�R�����\�x2̯�_�p��1º�����@=3��'�+ߖ��e]�W�_z��u�ؚ��<�}ΙZ���k�lc�{�5�ܚ칑�v�u��-����z��gk΍vf�f�ڄ����k�����}}�+lӽ�E���F����oJ���O��!�Jٗ���M�휚���y7�y����T�D���N���B�^�؏M�o���_V�:˼��Zt�Խ��E��y��^��},�9�-q?���t$͋ZB?}�7���E���be��[�{��K�;ck9�����I���"s#G��Κ��*�)�_$L�Ǉ.�R�ME6�=>�a�	��i+o[�,1\�<��N����}�ESJn����SC/^E������q�kQ^Um`J�.�D�VUc{k�^X��0q���v���q�e���N����o��>Y�+l�,dzg�3��T��9���:_&p�7:u�kj������x�f4;��R.����_��r���بzҮ(L�W=�QP��׋s�
��Ԡ	�E��\b����1�"���ߧ���Zz]�,�>Ӫ�3���9Ui��к!�S��O��{pXE'�)����R�-~�އ�;@]��G�F�����g�=��������P�I�MD�2����IP�%W'��9�?��Ǣ�ۚ��GCȍ���.�\�-�O9}�����l�~�>�o�޺����
i�~��p�D��m;f,i��6���}k.*}�W�.^iww%�L��[�X�~�7��uI!w�w:�R�_g9�JS.mu��������� �;��~�}�;��,_rV�+�]b̓�u�(u��	}{Å^I��R���\=��΋���ެ�}�9��m҇�D���\C�.!� �P��3D�k�<�Aaw�G����ԛ%嵤Ft�^%#,�5�,U�wŕ�Z�ܯ�{>U;�9�+���jp=D��آ֩!�$���_|1�;��v�1�=���v\D6��\��!���/s-]"9L���P���{\0�G����|�O�}3�[9{�n0��q�A@-�*!'��0�&"�C	������xf�������f5t��]"
�B�㙘�o���lw
l��b��֡���h�I�ΨW�z�t�>6z��;�:��/�
b�眩��ֈÂ��}y>|&�ͭ˱�9�|p�چn�JS��sG�U�Px���1f<����J�l�@��K�N3'�	�l�́�������S�ӹ��q��ȏW��#��x��+��F�p�3�R�|��o���Ql���&�u,�ꧼ�Z6���*�l%�*�)�x`'��C��ߘ܆e�J�/��Nvw���"P��U�;���L��	�zb���"�h��{�0�9w��}��qϚ6fy�۪]/�Q1�̛�jSꕪ���L��ۺ�Z�sH����ǯQ�u����E���eE��*�4��Wi5����T`6Bz7�����6��l!NwW٫�]����v�^(wh<��:����q�G��J+��./v�`������ׇ���9K���I��N�~
K
.y�t�Z��И��M漡j���rɌz;����R�kQ�!ͽC��V5�s���Y��h�S��9b� �dk!H��rE�b���r��6_m���y<&'�]��i�H��v���͞��T�ǒ1c�O6�y7l�5Ѕt�!y��^�P���}	��>@�O���ux��.v���?��I�u�O~�<d���|{��|\�ˆ�kԃt�}!yo<4E���sg�5W�D�֋tt���&u�) M�֏���c�@9O���8�Ig,��ő���K��h����ם�=��빸�	q�OP���ric��Y�D$xQ8y �p��x�����1�(/H{/�}������� ���k����7��r�j'���N�O_f����V��q ��"�9�Hr�ݚӝ�������y&<i]RZ;'�\���<-t�TZ]�Z���8N��d����7�
�v��q�����wB��r�eذ����Wu��ԙ ���C3�gF�74^E/���?{�3���Ѫ)�2�{f>t���p_[c;��U�^�jҾ�l��l���:Q������WBuj�r3:���יSs5A[5�ޱ����ko�y���.����o0���5m���PPf6�}R὞����w�55Ez����ʹu5v�K2�Ӑ���c�ZD��v�}y�!�i�w�q��L>9��dr�Mz"���K�;��]�`햾�+�����4�!���'"�f���1w��s�T�۞g��ܟ���"���9���u��S�^ׂ��n��о�N�\��o�U8��`��[P�E�9��f=���se�6>�Ƀ-��3�N9�6�&��Cc�N�$�~&|Q�1Jvgf|��}��7\A��v�F«fe�'.♭��9m�p84
�ДzَNK�.}��;�n{�Z��I�׏�	ι#um��������j��9i�������K��A:j�d9t K[:�fj)v�F3$�ޖ��@T+�n���^Q'W�����mz]�D�&ʘ	�����	](*bj&��ڶ�o ��q>F�k$�d��&�9C�,ᱫRa�d���ݍ�����+�m�o[���.�,�̓1�8�����}��9�Z�:���۰H�P��Bl~��rv�F�#���B�A�I�v<>�ڡ�����sY��Q�[].���%ٗ�1��17}����F}_+���p��D�v��m�W��]�km��fy������*^�Imur�����N\��ڳ�vgrAzN~<#��q ��#g��'��}	X�^K)�����uq⏶�1{�NM��a�*���n�Ê���B	)}k􏸪^[�2SzF"�e�=^��.x�|��$űj5B��� �2���&��>��1,���C"��\���}(.�yE��LMT8� ��(���2^:�P�w!R�0�C֤39}hw�\f��vN�*s����`
!�����g���Ɩ�&�1���n�W�\�>����dg���t���)����<"\O1��w��";�3�ia����\���{�$��kK�p��H|?}�4�5���[M5J��'���]t�Qp#?.��X���;H.�tF�F���m|�a>ݙ�W���t˚E��lv�	q�SQLT���!4I�	�r�cޭi1\�;r�nu'�nM�u%ޙ;��|6͵0���G�����f�]�_��olnx~����FY�����e��rbD��Q*9ΪO+�1��u�´��D9ra�6	F�w��L���q�/-�U�E�Ow0(g��!ƚ�n�0���y�������gEK�.jk+_��:����.�C\��l�(8*�`�FL&��4i�ku�ʃ�׭�Jև�-*�<��d����OE��#��
0<e%��fAn��ȓ��g���-q�;k22�Y���r��f^�PSb�����9�q?����E%�����yAacR��'B�9z�D��gOZ��h/��} �����/&욶�m��C�)�4Q�¯�qz/�b��_��n��Ե�`�;"�x?�]ځ&0u�o-�Ν�y������z=���R�ޛ��p��M�*����̴��>*-��s��s�E��x.UgY�@Wÿ�zbzDm�ͺ����v���k	�>��ɇ	ڃ�RiZ��v�r&�)\n�l���>ڊ.��幤F��oVt���hY�
�,ث�����y����+���M��bRmo�(k���qiϕuW�x�IZ�S�<�C�����/}��و�`D�4����!�)�o~������CM����ͯ!�!�װś�;�%D��6f���m��^����)�q�FO��@Y��Ol0���θ��Y�7��������1���e	�M��Cȯ�4������j��׉D���?}�w�X ��8�Y��4�0�B�Tcc;��/X��2̍NC-F]�4���;��
fk���_�$^X8�眷k�f̾{���u�r���]U�Z��ھt��pkafw;���ttv
��P�Y�����[��9o�D�t�Rk��Cu�N�ܠ;�he����.�j۹݊麻�S9k���v"ewt��ӹ�C�h_7�vc��G�;f:��3�V
r!;�G���*�a"�T<r�i>S J��M1��4.�){/�Vt�Բ-qw�4����|3���d�	7J��̶��a�RO\��w��(�߃jIMP��J�|u'������6��T �v٢_['�o��Wl�G3{�������v�-��v���]�'*��8�����{�w:J�+��M�a����>~w�ܽ�6�B����iv��+UË�)/:�MsT�-Wo�n��n�a`�2ຐ˱a��9���ܶ�&ƽ2*�f^�fˉ�N�{�Ǫ��ĭW_!��H����.���xn�J�a���8A7���s�����Z��v���Vu�KՐJ�0,H��=�Z��l�W��E� �o^ƕ��&v䳖��&zY9��A�}�F\�i��(�3�Yl��ø.�iҢ�x��f7Ӊ�/.�wkޖ�l��s�tY�gcxj�*եֵ�6�[����˔�)@�q�� �7�w2�;*�[C-��!��ЃW��n����Q�Id�m�Q�!���A���&�邥u1Y�P��X���j�j��	���U�/!b�)~Tw���9J������jZ݄4��*�:a{+��j�<	�k����m[���.rz(w,�Sʯ�v��مm*��&j��_D���l�$�9��Ҕ���ϟx@��wd�Vc�y6��"���cG`p_'uq��L�Ӽ�<n�ӻL�r�����+ �v�WVt�f���	w;��SgM�WPg:m�h��x�\5�)Zw�/\I��Cq�;��:�3{m���'��<�%�y���h�+�;I
�eZ6���Ef�Z�W\�����uO.��f��I�)C�)��[���V��`�%gtC�rؽ��/6:��/�}���'�+�8�l륐�;N��I}!:8�y��C��b�{�Wf5�(�	]�WW�Ҹ��;�t%��V�G� N��Q�9ww%,�i�8#Tä/S�-t�[�̺u����Waor%)����uQ�w�Lѹ-nf�莓���8�c	D��%fwi�Bp�L+��fs=��IJ�c7!2JՊ�nN)M$'�<�>�����ǌ��щ��hK%����"��l�����t�B�cm�[Ձ΢�1�5��1�$�(-:�/M��;�+"����9�Ւ���Χ��wu�F�#P�N���o���u�����ۙ9n�ގ��E�Z�-� �H��t�#1�R}�Q�#$��T��I�)��<qǎ=m��8�q����}q����(KI�(�"I%&2i���}���F����>�����qێ8���4��7���{�i����H�RJ�W��Y$�c�^����ׯ_Zx��q��z���}z����Jź뤤(~��0���\ƒNn^���������ݏ��34;��}}�K�.��������l_�_BI'�D��K�
!#}6�:�7�ׯ!HT�ۥ�>�3��7�Er-�֗�\���F��?]�F6�]p�QW�/����>�wE�d3��+r��1��vW4��X��w�t>�G����/�]����n\�PB���Y���o\d^-��l1i+�c;�WV���ƻ�D����3S��m�1]����
��5��uܑHRZ��<������(��o�ʀ��U<��FG�:�H�)L��si��+��s=ݭw=�Ǜ�[n�����^��]�Wx��\}���cqK���kЖ�5��Һ�Z�7ypOeF���0s-�
��9/-�)tHw����>}�uFy�8�ܾ�����m]����r��r���E�@-�M���p/Tn<4��v���o΍�����]���g���I�v��t�G0���p��}Jr����Z�a�C�mm=�6<��wkz.�2o��h��흜��|��ok�A{2��������ڕi�Pۊ��2ͬCY�����.}]o���`t���|kA�ɟ[���4�D�u������J$etT�}�߯��½or�p�,a$�-t�w�m�NE��߯� ��/�C8�fj��.�b9^4.f���2�)����ݹ%���}cE6V��@v�`zu�L*Tu�/%�{���yt��&�/�j�K�Я�Hr�a�ru��xY���擐�sA=Y��	,ϙ����
(j�^l�/�C��j�6~�����e謑E/��d����y�����EZ:Ty���j3���x劺��xp����a����	�vтW�qRzbY��z�۩۵�Rp���
{k� ��=:����Raj]�
����]����p>�D/��Éq..8��Z��~�!spZK㷨0`�����d$�-.��^��h�i�ŋ0ml��m��/P+�b��^;��"DV��x��k6���%꜁�9�ׁ����1Bc���k�N]��}&���ݜ���LO���o��Z}h�;�~��o�F��/�ņQ-;ձI�����l���҅���w}�Ŗ����"8�w�ǀ�a!֙ƍ�t�p��	�y�ͼ�Q��'Y����i���;{��:�n֒x�+���ʄUhQ�v��tެ�V���s/�߰��sX����W�)�ֻ�v���[B��Tx������*�ݫ�r��dj����&�^���t{a�)��[����{�^7�v�m�"�����G�}��}�ڄ��J���d���4�޺�_=&����z�ފNo��%V��n˰�MH�5KPZ�v/BvT��/L���Ir�T�g���
�	>�⍌V/^���g��+n҆쥞d5����ks��ѱ�&O�M5���]k�g��d{�s>i���������j������w�N!�;�#�ʦh��UN!�)�[ڙ{ѵX+�	,�c l:L��ƴP�Kxc�j'�U�]�\w��u��K�创�s��[ԡ����ו��Vj��e>Vf+Uk��9/��W��!�9�
Dj�'�%�}���م�Z��ݡ�Ӂ��]̠.��,b���[�f������RuD�K��6�����ϫ{챷cz�f���#�f/�L�~�#���u��L�`���!��1N�as�S��
��*�hgל{HV�Jx�F<wG�O�y��������.�jS�|�8�M��`��W�0T���b������,�|�~�{�O_�����m��We���B"-9�X��Fr�T/�������i8�weI`���Y�����~���GF|�/H4:��� ��=L�sЗ��u�[�eH��F=Y�H{�#����o��xr��61`6a�����P������\��]6���P�ִ[RR�q�j��&$2,��.3��P�	����՞]��"��m֣X���q��5r��\�n]�#9��@>�gU)��ht�ώ�#��?}L�N��e?���#=�s�e)~o����E�\�n����-5�uaЗƇ�B��vk�s���G�a���MN&ʭ9Ht
G�@SQ{��܄���k��p>�w3}Q,��{�dd|3ꈻx��v�^����2Ť�^�cl\��!j[�EӪ�w`�d	��g��p�J	��=�Z��;e�&g������!��r��o�6��iȽ�݄?�\	�K�7���Jjn�ݎ�t��.;U��LJ\隑m�P�q��]�D(������Aq.�p���}>����V�0>�a�� �D�𧻓��ሟ{�=~"�Z�ˁYB��j֐�	���zO��}2�6��h��Q_�Q+-(j��K(�e?N��Wg4�==Vo�9�2I�[�?�M�(�3;����[�.�.EX���b��(٠�y~Cǵ�xw��`��Ae�	#Sw^fBƮ敬uTȽ�3m���T_L
��:���@�3�lx��Xʷ]Ƒ_Y�^�o��y�jzO)�?���@7v$[un*������gw���)�w�.WH��=1��@;B- ����(������}mG7
ߛ���@�c/��S^ץV��l��AI%����ņ����юl`��Њ%W'N��x�Plz>vt�u����_`���h�%����w�L��f-�����5z�g�1>�م�F8�L��wu�c;�'�W��q~�����ݡA�������988���5����}q�ϋs�7��֕$t.i+�|�1�q��Z�Iv��0�s~�x�<�������P���l�d��~�4�ɢ�b��ŋ��+3��)ww�	�����)a.��w$6�����#=��0Y�}�ݘ)%JP�Z[v8���0�'$���b4���TH��']�vS�Lv{��
�m�8/��y��<�a�W=_.-統9o� ���o�^��^�����wj�քz�H����SY�T*�7���L{��>��ܲh�|u������ʹ�l\I�G�7B(F$��A2{��{������-���O����qmm~�Ny�AD筌��x��_",>�l�b�'Tu���M���;�Y����ؓ>�L�+ؙ�S�����9����F{��l� �L;gR��5uǢYDB(84>@O���N[�Y���j��~�b�К�]�Ͱ�cٮ��{���I��{���ٵ}�3S�x�C�K��1q�)_˼e���Aܢ.��b����R�g���lV�����ڗ`��^c.xnc��X�r&��d<2��M|l�w�Mo�)��Zo��'ߞ����^��-�02}�����~c�B�Qux�Sm9�w�T�8��v]A���6��0^pCc�>��o^kwf�͌��n�Lҭa@j�^�iJ素�8�VR�a�ܲr^�:���v��-��*�Vo���6�->G�~��d��̆h�u�k�F(���P�y�h�wûҼ�=���ii�+���2�k�8ؠh�����厪��e�g�U���}�$��o�'�����'�H���|F���;��+��6ݞ����P�B.�oA.�ڊd�M�:e�GnNݭ9�^�D�Md�fg�|�yVw}�~���������;�XϹ����~��}�l��xC��ƴ	��H��گ�S��P���*�(D���ˣy��3���k�t?6$�X�5���(zPK�FO'�~��5_�g~KW��vJ�����Y�.�V�Ld^�f
�x��sZ�#r[m�r2Y,s>X�-��ԃk����}�C���P����t�۷�f}�tD�V>��Z�$U��0�����d��ߣԇ�j� Ѝs�(7	`�2ʞi��i�6agg?M�[oL��=�z/q�F�S�[��1���!���g�r��;�p�=�嚄��M������~��Ƒ��/ @ծ���f@M�f=�\�`dC'
�~���Ϫ����#R��P��D�
�:�|}u��,�f��i�^�v�׎/W:��(�n\�{]�`�d,2*KWDSG>s�O� 5����'��N8��.U%.ñ\织��gjk��Xp��
/��Y훍Hd�d��g�b$C�<���SԽ7�����3�V]���ᜤ6!Ga�坷��q��i��w�+��tdy�$�.��=L�++"�-^@��t���c��)p丽��=*��<e�F'��M��MǋQoz����\�^qټw�䋱������M�}�1�Yn���L�1Q�v�����Wnlӑ`�'[�n�M]��YT�k����Hi9��� �F���Z�)��h�}~ﻛطgm7(�������1�v�.��㛢Ԋ����?R�-QuC\���,k��P��U�-M�"!�].����a�ܥX��6��_���<��e�txM]�tӯW�O�H�*sX�l�~��s�*�WoavP
�ּ�ǫ��<<�3t�0�nm~�����8Ǌ��kd[,�u��u�P����r�eS0;��\�6���+a��ӥ�4��(:�"pbnN�ۓ{U1����
a�*)���)�H�r�٩̈�Ϟl�����Z[tɍ��߅e��l�O]vět�����R[�z�&{R���,q#У��}�a�tz^hFzw5�&�V�ֽ�Bю�9��^ʡi��㶫�X��K^9�ǝ��`�.�4,���}��e'Qf�d���{�xp��2���;"oT�q@��'I��YQ̙�֩֗������Yw5�P�6�z/ܶ;�dD�����>Ud�ޱ�*dކ}[\�������b��9��9ІB�ScW�����f�w���aa���~1��*c�!�B#���%zX�D��-�*e����H�E��P9�~4�<ْ�҃n`�;�n������g&��͚�d(�PaR��O�����m��x��yf��ˑ�c��C&U7��f�o2oU��ؠ�K�-�'bt�R�H��Qr헜�+�y����������s-������L=��ghk��8�W�z�9�/R�~P�,5=�%p������`�ۤ�v2�meC
�/��9�E�y�x����!��+f�CS+�+����2��)Ts���e������;�3��ux���E��˦�7�t��������f���KSJ�e'��v�XwGa�3�0P�zzj/r#����^y面Uzx1�摳��m�950�A|\l��Ӥ���{༎�ɨ��5�o=N���>*D3"��-�	��&�V=���і�"�B���W1�.�m+.�~�h4U�����<�(�!C�w	����՛[
��;�-�f4C���ql=���n���!��DC��w�%F�kخ�<ǋ���}�����3���.y�%�QݖKz��{��Az��[�,}�̨,w�<t�C>�.�a63��L�
z֓�5e�o3�&��<�Ƽ �o>�)�S��R��<�[uS���q�#�@�����K���R�[����]y�C�>,�� �U�A����w�=힫O͉��|
�yحHu��9W30�>�g؛���ܻ�h-��/h��?d��x��`�s�F�;kzѕq�#���|ewÏjn��b�,|�q�M't�S1�P��im��:���)���N��.X�K!4��:�Z.	�UN�&��F��|���< �����������t�ե��<�עe�Ū��.�*����e�bF��H�U[{l�`�c�u��ވ�`�CA�=�O�#obϩ��s�(�^ɦ�/:��'y��L��hk�Ŗ����u�^B͟�i�н�������+�b�/-�1�4��]ɬ���o��c��^+�ȿ�y�c�1�9r���ώ�0�|�����RGV[�����|z��U}�����~�Q�c�+����3�y}ʱ__ߤ ��Rc����n�/���c]��Y��.�j�q�S<�5��,�mWyN�1�����2���;Y�{8�	��z$��o'kA��xE��P��͔k+�jk8-���X�˩����&o�����74��P�Xg\*gT3��;q�~Z6|[/� ]���7cB��C��>�Kj�F������3��cd%sHS�r�ꡨ��LLP+b�v�ʄ�ʕ�Q�\6~.�6FY�sʤ�A�ؘ�"�����l�YN�⁈���zw��>��D٘�7Ho��A�e������ǅwk�3������J�V�¹����+��6��uZ�38�e%&F[']1s�2��}���\Q�xj��x�+*k;e;�Ru1K��9ô˜+���x
6�N�T�J�Bf>���=�}�T���I��Ç�s��ދ�P�<�ß�kH�ɏ%�G4z��_�����p/��z���ub�Y���K��`&�Yg\��	̴ޒ�b���]׽��<ն*ƹ͍f���"<���w՟	�3�xewg����g��sH�ΑЖW�$M���4�.u� �v�ش}�0h�XU�k���a�x���r��V�{��ll{��%�u�I�_O��ж�6t
��y6�l�m97O���3]gib��ݐ��r�>N��u��e�xN����&d���f�����fS�l�\�L���cQ�U�L�_�ߟg�:¿j/�f�4�i�������ٮ�Qݺs�'Z��>��@ֈ�F���1*۶�sc忄${'�qư;�^�r��l��l�F�"��i�X`e������ힶhd�85����[��s��z���{��ݹDmk�/Sz.E��Y}΂؇N��n��	��B6Af��m�wsy5�q:����ׇr`�O�#��-{���&�ԩkҼo��y�f<U�{�U�x_�<�8(R�>�Z�I���ծ��K�C;,MOi��x�ǆ��M��OGk�l/��]�k.ge�9t����o����Y�kj����S��4eN�P�w,������\�7[Sn�I�k�����+�����Z��e���3�C�`�>�A��
(�IvV�\������M9��@G
�CP��ԑ�֬�W�oN��E����Wz�!
��Bnhk�-І*��d��l�|�I�\�_k��ە։:*��E�	nP/�v�C3#�֫�eAN�=���E�_KW]}�^�����=�5��ʔ�]����*ml\u7ʤ������Գ{u��G��"�.B����z1�:�ͷ��<�b6�\9Qa�<gK��o��@�[9���e�v�T-3/30�����ֺ�Ո��LZen��mp۶�B�ZpY�\�t}:j���6#]�ˢ�F�O9��f���f뭸.���`��Y�UH�j������*u3�MÛM�0H�/�Pݺ��`�-'�h����]Vto�ܼ���1o�4�dQM�nN�Ͷ&�ǍdY�&�t�W�S���4�V�n� ��u�&M���Y
��#�Șӷ��#���]� Q �Ƿ[�s�a��?M�}�e���[8�f���x��V��tV52f�6���C��4G��j]���`�a�� y���.҇)z��ɬ�ĵv3לiam��}��!Gy,��싛b�m�]L��f9�T�ehxv�0�3}���r���eL�mQ2K2[؝�Y�����Els�bdy����
���}����l�\�a�����Qf��;t
q�uj�� �n�������@]�t�S����oTV(.�M��v�劶m�=K'm��)���K���&�wj+�;F���C���|�v���%��&g]�wْ�$s��tʾF�[�%��6�������ˎ>ySj���u7�r�F���9�Y��YOcy|�:
��R�ʾ��+eF����>��aoWk#���\S���E��S�P�%uٺ�Y���D�P�mdWm��{m�L�w��R�D�n�zb�;�ы��ՙ�Q�r��ʵ+_q�����3�b���J�ٵ��n��W.N���#�ob ��G�)�f���:�]��":ȯ�m�d��q�Ƽ�N��);.�v�3�����6r���}�E�f�����c�sv�C�Cb5���&$V�n^�ٓ��$A$�O� A��"��$M�]\��.������ǎ>�㏎8������n۸� {�[�"UPH���#�PI"Hx�����O���>8�ׯ_G׎ݻtkP��T	*�jo�n2��hH��#h��o���|x�8��=z��}x����k��]?:��u�5���y\R��s�����r��V�V|���n����z��$�R�{%�+�� By6��HB����E����~��Ǜ�nM�t �+�n�4&���n���c~������A�t��\�깿;��vߞ�A>��������_����}9���h���ȱ���K���e
����x����A+���	g�@y*#��J
L��Lca��dFT��������n7f�t�r�8E�ۇ��A��ݙϯ2�iP����|,��-�<��̺�rw�;��� (��`��E4�B ����r �\�1	���b&AQ%�6c	�A1��-�1dn�CĂ,8"- �(Ă��i��E���[��J#
&Hb%(�FȌE��$��xG �@���Rz���bDv]��wַv���="�eM�ѠE�����;�!�|$
��������;�{l}�+��֯0c/�Y�.ǳFB����؍gO\@�$�F�&��|�U�ڤ>�>�X��6wE	]�p�Q����Z���Gx�� �ʟdM�^6Yk+m�.��@U��;�_��]j�����vI�=�[_�}��'��_�,�S����E���I��׈��|#�ƤF���U���³��qs�޵U��C�ް�sqb���~y>m0���Nf���t���v��W�:��u�%ٞ*%��6�j�Y%�뵮�j��Z"���l�t3�5���EDI��7��!u����]����.h`�Zº�ռ�v��a�<�θ���l��\�0p��R1�1T��>=�W�?nû��^Y��
�9���U�x�c*q���F��g��?��|�:'�x�yD͉�-�����LI���Q�]��/�m̺��������@�]��9���")�fk��걼h��N�h٩V�=�A��A��MV]s��͞���A嬛��l/�Qu3u��vFu��Q�����:\�u<������y��*���Yz6/�[}��\b���u-VD�ť�wyg�r��}i�&���v��ZR��*_�a�%���3#W7�Ы�wfYE�8�6�܆�q�<R��f{��on:�����N.@7����=���Bg@�Z��p��O=�!�ێ���lS�n!�S�n�n�4���ی`،���aճ�3-g�
�;���o3Τ8��l�eƕ��l���O��}�FQ{�%�����Mwv<U�9[�c�׍x���)��e�繈�7����4���O"w:p?�Hn��K'װgj���N���k���"�6@ne[PE�nΘC6��S^�ꆙ�;��$���/�=>�t3К��ZF�jtW[��۩��g��a���t�W%B�O�)��;2͛���u�1��cG���3-_5�����q���g�2u� ͵��7�q��f�U���Y�fR��N{.�MY�{�
���U1�r��Nͬ��%�e��;@�r���w��L� ��Tjb�]�sgQ��!�ڹ:m�h��Ubws�JmJ������U�wG9�ם����b�?o�ެ5�ԓ��wh탾����a��X�n�� ��d�V*�7UϞ}�a�0U�YK�@���*�f�z8�`6�/H�u��%U��&�W�^ݚ�w��4y���
T�uM���w���ffUJ�q7�;�����RP������C�6Oz�'�gD�q���ۯ�D�NC_�;B���恥t���޶�\�WW��tb�vtlV�-xs}�����������$t
u���7�T��a�0�n�b��s�2����W?�#��β���>��.9�\u��wR�rLvWnEK�9��:��J�gN���l�>�����C�k�)��jl�LKŕz�j�y�h���x�=i�G�qi��{6C�CoC����x:UdٻrX��υ���_i��i�t��ٽ��x�鏠4�4��
����@�ݟE���6�_�]nF{���qѯ!�s]
M�a�1c�a��ulsMGrDu���)�3Uֹ]�wK��5�=��F#�C�/&Z��,�n��>�Z���uWn���m�vK:�BX�.޳��cO!��]�G�КO:6Y���3��(�y�[���
��{�0c5����{�#ʮ�D�Uf��_υW�{]d��� o7�B��l�����Ӝ�oO|��ŀ<H�~������	������QSa�^k��=ۏ�7;ad˵+v�L�ٕƊ6<1��r1�ɚ��h#%�lh`�s�c���̃<��ˆTzw��x��m�V��k2�1S!���IfU�a��0~�<��i�0zQ*�E����V�|�m��7q��6���N?1x�o�\գyJyU����pU<x�]��k����%�W��f�5
�p�+:uos��X���,�k��¹�v�wlZ�fCv�]�-��j��nb��܍a�
v��:�z����dotI7�ԣ/��x���Fe�<祽2�����
,�͝��y�^��|���0x�b���F܄��׷�����G��53���y�oK�-��\j����n5<0%���7��w�Ug{��Uq�����ҙ��LY�C�xط�����ú�{מ(�@�C�if��Z9�(�{7LL�.^��g�C6辎�)�1[��i�e'���!��k����v���T0~~{���y����G�w�گ����ah��V;�x}��:S�'l��ڑ�h�vV��C�"O�ʙ��|:�K���XӒ5y�?�8o [b�<6�#^��Sמ�j�[��ݨ�a�ue�u��1|z�4��ch�(�Oq-�q�+�=��)���w+�~|03
�n�g[	�\ճR!�6bknd�yS�M���a�*��FF-��n{MG��Ķ>����a�ۋ~}a�?����h�R���K�_@�N�7���ۯ�F�,��u�ݼ��q�͂��,�7�}0\K��!a�D�$���Rf�ur{�o2��9�	������tz_S>�95�59���P�4A-��j��_0���������^�����y�hP͹pv��t�ܚv2�f���^�{ [;����7���Q-�����,T�*������Թ����<��.f�XO33e5e�fR2_����65��F����l�k�tй���*b�r�6��Y�;/��as��1�$�N�ZPN�;����{�X���O����ձtwY��扙�D$���<ͽ�:GyB�x4!w���uvf+�9Yw֫�t]B@r*���.�ȮN���+�p��"��G��k�{빬��ϱ�𫜫��B"V��h�ڢ˳["��a���9���ӼWk�ZE�õQ4�q����C���z�XS9E�^&�&ݰ��^&�}8Jݲ]u#�b����O�9Mx�B��N����7y�P^���=-���-Ӫ{���V�-����+�p �+�����b�1�o���z�﬍z���yX�1h�n��D�d3����d��Uh�z�{�������Ԕ���~7�t�����B���i�Xl;Av�ۮ���~��v�n���8�K����ѝ���΅Þ#���Y��ݞE[
X�˞R�z;{��x>>�xN��fl����۾n�c�qimI�٪��J�vQJ0�]t�͞�y$af;�@<�A<�&g��4gKia���[p�I�r��B��x��!�tU��U�>��h���[�E�љ��7�
���qt�]-���w�{Yyf�c=�+���U�\���8��۝oZƝ8�:��e�M���� �8�s|]أ��8)\�{(�pzy�ySx�1�k�U�r��
a�[�$0��wF,�2�����z�������;,�'D)���0�>m�|��������֡ j������lfP���7Y�9g-��Ց���;������U�x�b�dw5�W}�蚍y����&ӾoK?\w��E����ĝ��"|?*�s)FU����L�=|%ڨ��}�#�m�:Z���1T�[��<�؜t%�e��\م���;O�LoW[C�ͻ��u�����q����q�r27\9���>=���X�=��J�jrI�TV>M�)��<D�ٍ�:������c,4.8G���##I�9���H�q����GEpa"�3y�\��7v���i2q�O ��+L_sF���;áo�qS��3�o�ƙ�Mٚ0�zx.툱.`C�9<x����2ݎ�ĭ�`�p4�J���p�z�f�_:6��=7{^���y�"��>��-�^���R����f��6�X��I_kIP;WU�7��b��k��L��^�*�yA�к�캵fڜH:�� �D�A�3I�e��S�eWK�x�����%U���Jꩶ�,ά�׹�fț��`�H�]QEא�=�D=�P8�k$C��o\\K��"0f*��$]��6~?(44�V�;T��5g_�S0Q��\]��|2��9��]���F.ۦokۼ�/�6�$��-1�^�c��j�n6Ʉї�:��vi1���ww�f��YK%����.鲹j�+�z����Ɵ�����<J�yj@l��E����P������6�&}��tǞ�N��e��q�j���v\c��8u] G"�`��Ś����a��e�-�*e��4��������hl6�����ފV��g6w���B��>2ԿQBo����O�,�J�n2�͋���k���_(�NU�U�����m������[�]�|���-����nV�-e�Y�YM�x��U�2{N����&T
�="���t<n@�edϱw�"e �˛&�E���RqWD�� �{�\�=y��犑e�R�TT教Z\�U6(�ب6�:� i��c�ۭt.x�in�7q�ظpB�(�K�w��bיTRCv^���4�����>�W���Y\��Kˋl���u�^:��]����>��v�k��p�[�1��-�U�X܋���H� ��..%��?_��\}������G�*��3�^kɍj�53L�'Q�����G7*
���6��?��˙�s��u�p�������K
Y�5�Ǟ���˗���˝�9�f�����ex�̵���bϲ�=_	a�R�bF[�������:��Ϋ��,q�[W^=�+��5�+��}�(�ܬ3Ÿ�3�!��Mbؕc��<��ٷ�ԑ��ԍ`s��/q>�53}ݽ���I�8�膈xx�/A�PUSn��K|�r��r}z�0h��� ����C{�1#;�A5w1���^��_c%ǽ�q��2�m�OtJ�f�nF��`�^õ�m�u�K�Jw�|ޝ�WC�M��u/���k��5��X��(�H��(�Й��+�&ql�t���?e��~_�<��v>���$S����<Z�a�8�z##�@*(R(k����j�ȷ���v#��N�6������aV��ڛFߌ@VU�B�����W���G�诞��P{�8�5�U���)!��f��/.0���ϫ��.��S�P�w�}�g�r����u-+.���6�5�
M�1�]���
|r��)�*��͔�B+���$����]}�rO��X�1����<�������]>�U3�=s���K���l�8ө�>~T:
�i'���yxDլ�T[|/�_g��æ�N��^�T�U+��Q`" �v3A��O�q�������:`L�]��^Y�ܲ����y!�GX�v�^�"�f��l���@���S��1�H>����aK��(�|�k��0��eGF�޲j�ټ�[Vؤ����[�)d���[�Qȳ0m���l� _j)f�G�WO+�������>�+�pt��y?:HR3�S/ky��PJ|{�����z�WM#�Fm�{ne�<x�z��N��x�ڇ���3��ǘ��Ż����]	ͨE�Uvf�bU�3���&;z�13��hǲ�M���]�Y��qG��\S5��^�J㥨����+��p������#3���o�53`�R%����#>?[NXl�67+Y�x{��i\��eOnF���EӅ���rW�%fV2zJv*�MX��Wtu����d�o���VU'TS�/1��>��A�����b�r�G߄U�j櫫+�q�_ �f�=/,���r��%J@�˾�ԛƠ�2�Z����u9z�5����E��$���6<�m��4��˄��{YY�vS�{J\������]i�H_n�[��[�q܅�����al�r��r�,7�8I���so��$���sI���f[ar�2��Gm�����%���i����y9e\\MQH����6���~����J_�c֪�	[6d5b����	��ţ�{�CS�/)�2@[b�Ro��rЪ���q��wx�+��Y�nL,=��K[N�u]s�grJ����+�y�rL$\Rg.Y�k<z�ŔrƊ����[@�+n�]�%��١�fqS��%[��wff��bcy�6U��R���	�-1����۷Q��f�B�������Κ��[���n'4��j).PMvc:Au�1`F&{�L{[;9Ԗl	�Ii���L��)e�'X��1���r�Y+v�U[���G�(�6U=��6
��ƚ��/iK����������|�B^�Ք
��)���S����8�ep�M5���.g>ٴEv"{ Z(Y�X<�(�j-�Y���"P��y�\�T4�튭Hs7��[�ݖ;��>�Z�L��uw7��<9�h�
[t^�z��K�N#RG���A��l�T0�t&&n���5ٺ��*E�1��M�̝q��mֻ&�=�hb+-���o�՜����eoc��0�' O�[P�Op�%Y��ڃ���"b*�ǹ�j�t�s&��Ev{A�[�Բ�*X
{�k���8P���m�.�F&���b��ԭ�.[pvR�O��R��źѬG�Ջ�}UQ�=��fna��O�Y�O�w,���.��|����޺����"���auu���Іb��ݬ�9��ȫU�l`:=X�pGԊ
�`�vf>Y��0D�ԣ��Ql��+@���4��iq��6������Kܙ��j>{ݻc��g5愳���F뤘*��hD�Ϲ@�*�<�����Em_:��'՜�ʦ�VeFΔ/�����y��X���pV"j<�t8�|�X��n�)5b����W%ݞ��2��O��[S��Y�o�N�<��N[��9�,�mv�VǛ�.o]�|�oN���vo��������`�.�e̬����'-����,<ˋ{/����dʉ���8�r�R�朡3M�,����ْel+�j�zc�W2��}�K�r��)�tb{qp�t��Է8d�$��%�j����i˱d<�7�^Gp��LY	E�j! Hy�P��-@�o�x�ǎ8�>8�ׯ_���n��#�RFLM�W1�Uy�yj{�W>��|}c��q�x�ׯ_G��n߭��Q_��O-���7����p�#�����׏ǎ8�8�ǯ^����ݻl�j I$�**�V���o��<ڊ?�C�﮾T�n�����wm����k���6*��m���c����k��y]Q�����%���/������N���P:�B&�\�ϋ�I���Ew�{}*�[ʮ\�����p�~Oǲ�%����F��[�t��������n��j���W#\�������yߎ��\��7-���yk������ߟZ"�}�X��v��vwRx^�)�T��^n���Hu��(=g��1�s�	l�t�3.��ۊ�.,J��_��CƏ��Ɖ�f<���D4@g�{?>�:ѷ�\V�>�!��291����8�ka?�����n*�g���z"�����Th�z���~-�ϽoU^��M�Um�Bq-���A��V�*�=�b��}Bt��7=wW�Y�b���gj�+"��_)�f�)��{y{k�iX�=�H.���*�'[Ku��^6�K���Fa>�8��y�M�0��}��ZF�,Y�EĲ����5��P���5j�AI��]���?���b�^fs����0��/�$�g���0q��:0ر�7��}S�R#��U{�vK>V3�/�*�,�]����E�.�Oy��-��FC��r>����בV*�|�['ET�[��B��]	U���U�W�,w�`5T[��ɜ��
�(񺊎 q���������*���&�4afM>[��M�n�_��fU��'N��8z�*����6�FQ.�]n��9f��'Y��}O������F�a�8b�b��0��s�zj�˹�>e��W!���Nr��E��t���Cx�x�,E[*��ͬٺkbg��=��>��������8k2��w���#���,XeGW��a?��Fi�%[4��Z�eT�䊼��0�/*���A�����:�Q�gg��6��+9/�2��޾m�R8�y�r���I/#:��2Ȏ��wW"��$�S��ׇM���h�CgY�};@�>�s\+���^��	��~.�{�6�(�{����ކ�LT�Wg�<�&҄�����w*�J�.�6��}At8��3�v�]���gvݥ2��m?o����lQv���ٺ��;�e��-pr!@-���]����b���}�]X�����C�o5�:�)�sk�s8o:�a2��z
|�~�0.q;�oz���P��<z2�ޜmǹ��N��<@�����b��i��u���0g���O��c(�WE�u�=��e������]�k�sӭv��c�l��1�"&�/X�l����=b;O���͔�*�u:�M�3�Ե�h�x�VT۝��y��=/�������|y���L���5դ�H]bJ��Yj\S�)<�B��]����dǎ���/n����Uĺ�䲲���<��JS2�b��5C�m��a��+���4�1�_k+.���.�>�\���I���+q��<T��ggh�S�ѽ�$Ӌ�{�ݯ_s�K��N�gylN�k�{��-4���ܹvS����ڪ>��p/�A^&}7C{P��e�e���ƴ�����D�u���ꫡ:j%�Y�\�C��QK*�ڽ�`:��Q�]e�xnM��������}M���ڽsSd�ҞT*�襚�7M->|���u�˼ �"v��$���9x~����|��������J����Ү]��mk`7�'s�c,iW>|o���Ts�<I�WW�]|�:�$U�[�u��*�=��C�{�I>T����S=�f7#n����C8�V���w8��)�r��rZ��)�q���^����u��u?*n�{�rT��xߺƌ���ui��;Z5ח;h!���rwD���@�3:�r�6"����׻���.����Ky�B[t�=�����r����;�k��҆�����]F<�]�l��C��gsE�m6<�We6*����
#.8��{���L�j�r�AQ�4��pL��.�����U��6�8�r������,h^�7��y���_t��J�-���"����&�@�*�N,��5
�O5M����^�o2��y�p�<�Ü�w�Ud3�r�5m�	�r�c]j��p��g;n�ڴ���Ec�E�C�/���[��n�S�Jǽ�.{�c�)�unPb��<9I,�;]��e؎�xke@�u4U�t�'�(���2&sˮ1p��lA1�O��aL�*���c.��<�T��Ӓ[y���[�r����/���1xi���B�gm�fΌ�}X�"�]�����!֍3^{U1�cӴ����~�Fn���Ը3��f�4�8���G�n�<M3���H���e5��;��*�z{��Z<����:��fһ�m�zE�.������n�˶p3�vzG=,m�=��Ǉ?u�r(�'�zW|�fo�<
�����<�������'�P��T���1_\�E�d�$�A�_V�mR�PG��\>�畣�$��1,u��������ݙU����Ul�9��Z�;��%7�u"�+h�[G4�ѻ�opH쭇&���4|1�F2��y�'%���y$�R���|�����5��27�n�+� )� ���V��z�v�)��ջ<�����xO:��-����G��)�e'qnh����I�񵾿o_qT�ĵ�����H�QIo�_q�K@�rD���е�D_{r����*%/b�F�e�c�>���V��T�3UGwTd\2�����wwww�ӄ��(�֝����ۺA`���#��m�������V�9]�+�k�Bӛh��tݑ��鮣���Š6#=�a���Hf�>lL�@���D�0oO6]�§��W��m���{y��Cw�n�~��Np�%~u�6�h������R�kU��ޙ�q�9I�^���^S���*/�������� �a��Ό1׋��������U������5�O~����:]�op�|LJ��P��)p���F���L⸾�-����)?`�V37Ff�F^]&�Rv/��K�&vf�f��f���S`t�^����a��iڼ�~<u~@$���Ӷ/�Q'�nc��mh�����ؓ�E���E�AIon7�
�o�rR V�A�� �o7�{�E��_e��E5��5y����ᰳ�Rԋ�F��zp���lFj�ֶ��,�r ��o92cC�I��-S�h�d=�7*k�����&���x��٦,Y�����e�j�E��4���P�
+����Ur}��P[T�-�z��Utq���㒻S���񉳍�yvr����n�Wq�.9�X37[tҴl�.jg��+��Όe�+#���EUZ��i_6�Uk[C���*������5��=ۘ��]י����rkT_s@վM!s�#�2�N�uQ�f�'�Kvz�<�W���E����{��pا9��K�F��ͱ�i=ސ�s��-�s�'��_q,�_�|�c��\���J���Q�{K��s�7|�7�E���@��V:���M>����vBf��s`����{�岔Rz�w���BӚ�UETm[������LxWy�k��N\��v	].�-K��(��%�3��E̵�cŸ,w'њ�%4�
k�����duoR{\�H1��*e��=�=��P��m�R��YI�g������Wʠ�{)
v�<��$�mZ���d0lě�;�rK;Ӵ<0� =�� ����b2�0�맏�$�·����2As�
�zq�*�v�dXv��I�8/F���9Y7��~Ň$E��S���u����I���x��{2빚���}k�~ww�>�p����h��l7�����vfg�����3H`�g#���VC9̆���#�T3��3"�*�흻x��Z����FAMb9g�hj��\�s
�z�y�:�Y�:���=rˈֿ����;:�N)$������J< ���KB�v�ES��3(�j�K�ŵvh仍v?l�򻣇�O`qAI1x��V����0�FB�Jd�m�z�^�\]X��oD�Ti��WI5�7+ڞ�zr/#i>�i�L������=)�j��:�yEf���t��ގN�^	�Ͷ=�F�X�xvu܀��f=x�<
�;,�=�3>̋P/���Y�5�R̄4C�^ULa��M���ͼ{��f��-�w�Ԁ��Ě��-�������2\W�-����Ij/\sX_u��qY�<W][ڶc���{��!|-�u�V��yA	W��0c�
v�m��Z��oY5`L�]R<Ȣ�p\��}��Sq�ʸg���v����KchԑQ�|�<��sgt'+u^p��ō~��o7���9D�·�"i���g#�M1��h׶Em߲�lĮ��6BΦs��L5ċuB��&0t�EC��wioX��G�%��_|'N4^Z��a���;��r"ɟ��EL���M�t����,��E�p�t��*�H�]=vp|���5��X�x6z�=��Db1ҵ��:��]I̢;^1�FR*�e�Y��8�V�t�?��i�,Cu����*�=�����*�]E��gc��z*0=�)t���*q�C;3����V-��� ���d�$�u3�s>YGw�f��I���a|�#�"��qCқvp��Ž�7u*���<,��e���=Q3WX�]�i��������7�x�s�8Ӻ�`߶���Z+�8Sƾ��:�X�s����\�`�/���:-`�e�eٚ�����Ŧ������c5�=�x����wP��2���A������7/�_���]���{Y1У�����>U�n� �k�R�;�h�V*xbO6��=�i;y��-a����v������x-"��B}0nU�`ֽ��gd�ڪ�8�9���G]��=���c�ӵ��̀�ᦗG�ow����	�#0#��j��d���@�槢�u͋���n�R��A����d���,�Dn�e�����X\e=�U�n��gC_�u��TT���ܟ�y���ós˯n��Ǝd U]P���/t������n��g�y�]�m���A�j=����~7^ȣ�s@�w=�P�V��"��T��w`\]�ŉ�,���`W;I�������K!w��w��h�|��ejՆ��ƾ�{�1xTg�Gl��h��J;��[t��b��ۺ�Uwq��8����O����z��9q��zFE	,4��Z����q�B���gy߶�� %����l5g@��k1�#�T�]/�И��5z��U�ޘkɘ�w�s7��{uY�!kN�ݱ����L�j<p+g�~$��Kq/vC�]�����^��';,oz{=���$p�Gn�� r��Z9��룹�f�/o���p���\5�*���{�L׻�'�/���&�u�O� ��]�i%{ α��\/!�ʡH�-��7��*�s9�鉆4k2�2�����#V�m�tn�ދ9��ᬭ�]�J���b3���Ƀ=�=u:۾��g���l�q�C��t���t�xDV���i��r�σe@z��mH�h��p�T}��~3�=���~j�_�d������Gw0�o��2C�b�s3鲤X�滟<���sԨ���/�͗�ճ�Y�N�e�ߧ��s��c�ޟJ��
�Ť�$��L��oUc}�iђ7��3G����Ki���'i�%������ǔB�.�:�ÞJ�Xޭ��}s�K�&Z�+��da�9�^{�Z�á���6o'I�go�P*����@���J�R�,Wcq�M+#^32��c��tQ�����i�con���d�ic����y�м�b��"#r�>D!�ʹ�5s��%�0�Z�捎H�]��ʼss"�A�y=���{�5���Ϲ\��AA��e��}�z� 4#YƧ	�m��n%-�PՆ���B���y����//^p����`�o,�(C̼��
\[�9��+�`Mؽ��X�{�'���5��{^�oX֡\.�jU�Ʊ_Gn������f]jco�N��bᖮ���Ȝg�n�=;BR\�]�khֹt�5������̺��w4^��$U�q�DP�̫���,<hu��x뻰cJ_n5�e�S+mlۣ��R�e�sA�/w�+6�9^ɻi0��b�Fa�٧�Zv�T�*����Xp4+�g&��C�IkG�(<|�����u���ꁺ?vwn��Af
����oO{���xL��P����.z����=K���	[��D�G�b������6�6횴.�w^����e.go,�&�5��+\J������C.f#�&4xv�n��9��sa��Wy`���\u��y�#ȝ����70>��o37#��r�X�|�r�_,N�ۥT.�o��!�wip���tj�곙;cG[w����|l�$>9]����E�N�ۥX��{-u��W�A��[��F��k��dC���va�ûw���W�|�[J��g��r�E��gw����ܺbs,nܾ�" �ѭ>��*f�(T%������D�P�a�sN3X*�C����fɯ��sa*�y��$�*�|��W�����Ze�!y�Љ��v��w=�Uݒ�v�9_w����#'���(���Ey�2��؏�g^W7�����.�F�.*%�wY]�Dg*t�JG��-w�Gm[]7w"�%�p�q'�\��#E"�Ach��(�<�&n��.�}�u�c߫_3�^+�UQ�T�嗙]��:q��Es]|�;R0gf.4�;�trT�Z�]��.c�4�f����]B�-�ڨ1��.�=��y�yi�w[];��#C�[�K�d��;D�A)�y��y��A��W�$#EM;i�Eќ7:e��gU��A;��B1��X�Ђnv"�k����k����s4ۃ��+5�'X.��*-n�k6��6>��%e�#���n���Y�
3g)-ed��L����5��A����b�+5�r�<2���ɧ's�-��%Â*�+R����Ô ����-`]`V�[p��Vr��㝷��3^�)����YN�v�C9���m�w�����.���[��zkY�uv�AgU_\l-�o���s�1�{Պ�87���}�GyĞœj�w8���N�U+����.�}�Nk��zY&�-u�x�6��"<�(0����\��v�S��Z�5��t��}��*�Op�;`Y�۪��}�`���gvt��A��j ���3�������ns�a���fwm(ffv]�Ս|tMs�e��t�t���ט��K��{�<�Yq}ɛ�ܷ1��oG��=��!������W����� yҟQ����sͧv-�n��ުJ�@���׏Ǐ_�8�z���}|v��w�J!##T�S��h��ɼ;�r��wv��{.#�5t��>�x�><q�qǎ=z�����ݻm.3t��p���:�{��^�m�Z���|w:;��v�������q�8�����>;v��J�5U�Q�Q�%H��/��|W4t��U�q�lh�v�i�u���r���\ؽӍr6�wTb�{�u����O]\�\)"w}�m��ޛ����Q���>z�cs�o�r���{�lnk�t�����"źq,wvg9�k�q�|�ǎ܌��s��1\�Q��W�I���ڹh�󮍿;���|���z<.c`�K���N��sz\�so9�wurc�]_ϝ󯷦��{������	�;_�v3ݺ�Ʈ;�����_^�y_M�k�\�÷n(�]*� �p��A�=��[q4�#�1 &\��q�Q0�I�!�@��Q� ��X���1�08����b�GѢ�]�	���y��s�#{�k&ӂ�G���⻭�Ep�-�Tsm��Σؘ��y3p�e��k�p�n�*�,���JQNC�Ri6�1��ɐ0�-��h�ِ�d��@�A0\A"	H���Q*�`�3D�Q&�$�PPE )HD!q�SR2�h9�1�0�$* p ��!�[$�h�.�U��c�{���zn�׿S�3,��� �Ϙ)�f�L�͔vx��X����wL}]�wެ� ���+�_����p%ֿoX�(yȳ�3�S�-�d旹!�!��z3�ʂ}�F-�W�3��5�'��3�z^�.�}��xtK����%k�Ό������9a��bֽ�V�t%�2d�.������Ԑ���TF��L�W�:����x�+.좝���a��wI�vvg(�T3�m�1�d\J��j[��{���^�wl=�����J��5��{C�v������0-d|9��L;_UQV�z)w9�}�O��wg�ذ�}p�̮��V.��QbE�ཱུ��<����}����l��B�Q>~��q�$��Q�+����I�|���h��D��g�a��xӼ�,�e�
�h�N�6�K=�<��hMfR�u����d_M��)�׌�T���f�S�)ez�ݸ���!���nKG��Y o/	>�xB������W�׺��q��tTZ׷T6I%�5�2�9�h�j��SrUڔ���֔|ns<o�`훊���)�&�%�˖��2Ss�<S�&qWkw;���݂�IZ$[���� ���sw���9ئwW����dgX��(o�/}�3tu��n�so]�k��{��1�!ͻ����2 eC]�_�feo��|r��̞�L�q�8��7{�T�t�P��O�g�^I��ϑȔ��LܺQ��p�R��B����OD���/�_��ĝ4fϨ��Wps$V�V�-��i�؜�7j8��!�wr��eb��=+�2:�o����;�E#+4Y[�w-#Uǣ�-\{�ҷ�şJco˶�9u�z6D4]ߚ�+���i��x�w�.2V?��.�O��J$�w��*�]�ߺ����Ρ�����۲f�Umc�4Z�F�(ϧ^���Ӕ;5�L�TP���E���7��ՠ��oL��;ٰ=��.�Ƀ�J�j�զ�]�U^Y�k���;�eZ��l�k{�q��1i��:��i��%�&]�E��t�;�wW��[ �YLI;��
��|)��4��V/^V_{��:�*�(�fR�wJ|�~���T��x�+�n�6��IO��7�����d���G����]W)q<N�m���hz6�w,�����x@o0�m��$��xb0u#��t=�\�p����f����;5"��MMv�V/"��C��(W@�Q������S����ER��.rB���ѱ�fvc�M�]����v���V;'��x'فԆ��6L�Cjy�Wc�,��D�ڨ<P�^{JDMu���YgY��rL��N����nN�	 �}��NR>ߟ-�7�� 1G�Q�S3��fK�T޴dL4�k����Q*�n����|�f�
���)�5�s�"�P�"�/S#����K/
��q��2���6�a0�E�t�����G\S��<���1�r���W�[{�ٙSʺ&����6���};?T�|{�������{�������YٔH(�?,�n���H��Օ�g$�7En�k����.j�S�9�}�J'ν�T��<l1��B���&�ΕYU��LY���e-c���ᚵ��ݫ4.o>Vr�f����ZN=�ĕ�i�r}g8!i���"� ]pu}yL;��X�Y��zBu�tƱ\ܓo�X���K���*;�vT�'��/C���5��@��������^����L�[;��8��z5�g$7C7�P�[�2
F=vt�r�1x�'��hӜ��<�uu�S�k8|�e�>��漺뀧����6b�.{PWf��C�6lɼs$�-i��m�og�'*wZ�"����5��î�_����ex�{�DLof��{�>�Ș�^��5�º�޻uݰ�J�7&�5�4/��k�8`>r.լ.��L��[��^U�]|��<���Qcګ'?N�K�Hb�%��.�S��;ђ6A;���:�&��X	�ז
���M�ҚL+#��^�nr�����4^ҕx�Y��i���gK;h��R�f�����SO�o��t?k[�ϐP�3��R�[��v[�a���4KU��lከ�a԰7΍.�����w�/�*&�+V4[q��dB�UQ��V�45�>>�^Pv��O(L)�Ԛ6�WU���h�W1:�S��Z��`��9ǺSΌ7����v�����gq��{􆭴*%8���zw�vCʙ�o�ٮ�����7M=�%b�fwco�u�N�����_%fO;�C���1�������ͳ}�+Z>2���f)�{vb±:��q��c��Fz���t6�ۣp���h:���P��}hg�z��*�+;�&�d��ܼ�e;��٪���H�8\4ƣ̪�z�����oV���RU�����zڷ&�����#�����W�2����[�:��I��Lh��<�j���4��A�Z��u+�h��x������Y=�/����w�>���V<�p�{"Dxo;��N��|Wt���Ћ��!��ƘS0`�E�	�v�U�me�����#8��*<}4�I��G>/e%7�s6��nѮO"��x�W��w�w��&: ��9�\�$��2T�Z16��,Q���9+��H�Z���y������	��l�T��x�,=f�z�%Uy��Oq���%_�I�h�|E���8��:̋��%����ېӼ	�P!�����=g����D�V
�dy���"��[vb�{w��v�Ž���P��΋�)2��Ē#����_ۗ�g�ռz�M��u5䊵���8�;ޛyD��:�c����q��&���<�H�	����U�7���2˴��r��ǫz�i<�a��);t޳���y�Fm!�� �@?7�� �Bgq�0�_:x�K��xg�b<�k�0��K�M����8��F�r�Zb�J�饥��\�#y�G H�3��Y����Vk��ZϚשnt��>17}X��֋z����ɤl��T�1Bnv��wSSy�L�6���"&�EQ�X���Q�;2~-�u�뙾yn�{�iU����� ��}o�G�)DzEhޚ��)T�3�m��3xˤ�@s>�3듗�����H�,�L��K�c$�c��H�r�����">��F��
�^U��U��b�M\�Q\+/#�t�y��VN�\�xpa���{��S+)#�fo(��Wq�v����L`���\R�ݨ�?o<���pW����0.�4%�+�{`��_wc"Z/��e��}�׃��AW���+��,��os����z���n��c���Q����US�%�7�e:�]X����W��8���Y�����ϣU����ϘW��Z�e���9=�������rw%�ؒ*Z�a�'-�zzĆv�n�L�۶��s5޻�	
Y�k-�X��y�o0�63;����/!�)��l�܁���ȫ~�7}�޹I�!-�]�A������8u�+�����F?������@Iޘ���m�=V�������xuM]�:;�>(�;��h˾�l`f��Q��F�T�1b����ɚX^(�y>9�=ز��i��5�����6��0���2���'�_q���  ��kQ��~J}Yͦ��p���\�G&h�+�;�[ca���e�X�d��V�fd�]R9�HG�NÎ5�pE���N�;8��	���}/nׯ,;z�����m�x�Mc���9��!Y�m��E{����B�qE=WU��YgYZ�
��{N��ך�o���*�UJ�����z��q����*;e�S\:&7��F�����N��7�_ޚ�����;��qS�qq��}ma1�!�2ئUoE}.Z�f?�nL�R��ܡ�����k�T�]K�V��ҥ��!f����
�:���]Ʀ:�Ya�o���E6Ki<�9Z���6
��d���9����ㅚ�,�̓fv�3^Q�z�T.�&߸xxxxx@|��Ϗ��C���l���fQ���U]P���Y�Z�(ރ�G��S\^����ڡ]O��í�1�J뻼��iU/`/w��/A�;���)mJ��~(PC����檧�+y��ݎG�ni%���Hg�F�b�q�6�i�`����C�-K,�wQ�L�ه|ܛ�N�&�ݎ����#�Z�<ܦ��<ydj����}&�iZq��zr�a�y3�>i<��i7�K�哕��_�ѻ�����v��|�m|���n�Weɗ��x�h���g t�:�	ݵeZvGq�6�m�[�(TԷ�*2!DW;�z��N�[@�8<1��)�g��Dǻw��>�������{x�}�b��BY�W��o)�O����:��e���3��Cd^�C��{�Zn�L��.���Y�1���x�3#��?�ZX�;c�TR���Ԕ��cὑw�?xƑ���M�V�{޿F%�W:���9�sY�w�n岹��R�u��| �$Fz�Uw�]ٖ������i'��vo#�lX�e��I��)P�W�g�⮃��x/qfj�;X���~C��Uw�>�W>��j��>�r���'r�!}d�,A�6e�V�vN���D���s��ط�ȸ!a���_y�����/���۫��ivq���>z:i6u9�l���+���G/�R��)pDZu��h�?��J�ϧ����L��9���g�� 2�T�G<sKvY��v<�56фj���qVB~(�pQ�Cj�=f��)j/
��+��_�~�������&o��������W�o�ژ:��<�gZ�\��VKHY���~
���6;��>e�h���<ϯ�zF�ܯr�~Z�06�m���׮��ç1Q8�"񌈰���7���oB�,9>_��lU@�z̺]q[���9�iVI��%U����>>��P��J���`J<��*:tnʭw�����slڮ5����F�=;mf%�M2k�5��{��?x��������河c/��ѥ��a����ە�b����[���ڡ�^�O��3�A�k.\�l���tɣu[�`�݃���4pG+OI����_��vQAv�:W|�*��w((u���!v�GLZى�>�Y�R�lh�D mgvv�5�ƀ?��o0� �]٨�ļ�yS�B&�����iYռ�%�o�g��q��\wf����$�Ԅ�`�ȁ��T�jQ`>t�J�q�	�N&�m���=J��E�<3>��^��6������շ��^�Ly��6��U_S��5e�\����3.Ïjo@~��������D��%��mZ6'��cs�1�aʶ��#�Ǉt06̾3:�a�#��r�=�+�Ly��2������o4S�8=9���gϞ�u�'P�[��-,3��g2<�y��ݵ��B��Y �f�q��.��:�"�Y���o	���eR�{���s�u0��\��^5�.k.Su>��
��h��mv AV�2׭T�U�1fؐ�O(�#zSf$ƪ��)V�&��6,���I��i�ڥ��@g鐷����X�_b�>>�?8w^A��C�X�K
�Q4Eoo�ܻ��*-y�s�[�m�o9��uٲ�J�g�nR�ǫE�׼W[�{$K	Onc����b�Xw�s��a�paY�\e�n�*$!��զ��U��t<���ܼ�7hخ|�k�}�L��K��.fή�a�}��%1ʗnEW�*�5%�����R�6��e�p(�×�B�7)m����)<������YY����-�8U���O,B��z=���Ue��	w#N�%vVr;��M»��s;|�p�0G�2�̾s&�vT�Lm��Z4�.��O���Η�fk�Un�����*�����w!��������3�'U��l2S������- ؇7�\�Z6������r
�u�]���/���K]���Y�I���}�o.؀�X-��2�a���F�#�`��s��:pTsf���*�*o������9|n��;�f��k�*nBj(h�R[�!y�7[֟rںr7xY]����%�메te��+�.���'gXk�����wYHN�cqp��nà���u�����t��`٘s.%�l��n�.3r�	�}u�7���b��}�Ƿ^�L���)���� ��g��U�m^��0�R`Β�K�iڐ�9]�Y�l)#ř���8ϙ>Y�WO� ƗԹ�nI��84�+R3Hr�đ�!9�B��
�x�л�qc�wD�2ܻpynP������7��`ӡ���tƋ�[���9�u֞FK��q�ޭ�Q��?�Y��Og��ݖ-h��l��Nt�Y��MT��s���;+g�z:S���\z���g
������5��7�h�XY���_1��+���o�Ξٜ�jkN�D��[����FU�5d��u�j���CoyK�`���Wf,Ŏl�:���S5�즜��PS�R��HM]��F�@�f�@�Wp\.�d�udz&+���.�]p��$7�؊������T���f`T�7�]�Efu�w)\yVޫ��u�d��WĞfe]f�t�}� ��2��	��	Z%��Z�;]��fL`Ժ�sx�_,�v
��#}��Ҽ��1�C'#t�I��]L��kR�,�/�e�h��])��v��Äs�"gM�L��m�ih�H�|̷�����f*�-pXF>�v��.#XR�	\�����$a�����Z��"������\�)ի�(a�=��Pp%hh�kU����ZX���SU�Cr�JƎ¶2i��y'Uά��t�y���)�W(TX_C���Z��1r���g&In������^��㑽�v*��5�цFj�4����ݹr�7������n�|[�v�\(����;��h��{|ߛ�~o���8�8��ׯ���v�M}��k�(��bܔwF�F1�L�g:.����K����������q�z�����m;v��pwR�B��n��T�#K���?��뾜-���r�/(�*IQ�����ףǮ8�8�ׯ^���i۷Z�,�P�R��iy��7�sE��ܒwt�-{ݷwm�k��,TX<�)9�f��x�b����4�Q�C���<��W�w��������������v�ݮW�������4P���q�BRb��^%cEy�F����!�DZL��J�t�~v�(�^�wu�ɗ�r�tkswv�W�K�{�IL�����K�o��w-��;�ጛ�y���ъ��F�+��(��;>��K��	�q�y���9ǯt��8I�#ޔJ�euA��rLX��f�\�[�S����U{ӭ5kFP%��C�v݉�k��?S^�+P+��p1p4���
E'�\��ƻ���E�i<����=B ��.�k$Q�b�+_enȴ�,5٢�Еwڳ+$����T0�C��d�r4�V�+����}�ju�z�귘>��|�z�����S�%�,�z��ޫr���ʎ��^unEe�w�[9c���x޼e.�N�^@/�0�ȸ��ݒÉ�嬆Kn6,���3�����DGm�0��NH�gaǘ޺��Dk���l'բf,�=y�����v��n�\S���t��9=���g�P��R#����j-����JX�{��ni���t,�������a�c�s!jm�g��7_�;ٚ���0�Kwط�lg`ˬA����Lx�z�w,Z�lѝվ��� {��^F>����y�>7�9�����!�y�#Z[R}��hԲH�[:���i���kk*���� kr8j�r����O%,�L��Wئ���ʊ�}{�O�Ց�ʐxx�/��ز�om��d�˭��Ɗ����]��:���w!���(L����y��U�/�G1�gUG��6dD�*���T�+z�b�sa���=oά�����A�z�lG�����_�����Y^��4�{HE�H4����J��a�5�����c����4�5�.���o<��=�j�%��Ƶp=��.��/��;R��5���j��n���j�\�ܧ;Nj��V/
��WN�O z���ϒ1=	W+Ħ�Ǭ�B��M�Cjjq��K�+�`�
���������k�J{ùf/�lYf1@�}�|w�&NwLTTD�>5�,�X��_s�"�=���9~�W���6�u�K�ʻ���6ӎ�p���kML�<��נ>�2���h���VOH�f���Oe`�澲�N�������	M�6L��ľ��-�s�N:2jkh1ܛj�Ix��^f.�#�@�{t���׬d1x�s{Zif�_�@]�ml��@-���*�{M^��ћ��s����)��sT6L���g0.{�!J��v��R�nX�CR �~$y|�����oOU�����e��)ؘ��u-}�[���նZ���R�tQ7�7z˚�;����Q�^;���浏�wC�T�C�eA^mj����	��=����-;ꈃ��L��a��؉@�տ����A�z��]p�VX£�Z6x��toZ$�����F�Vm�1�@ ��0.���|��J�]M1���A63%���ɧ6�6����7e���G-�ړ����~}��"��"�C���Y��ݤ�8�{�����8�b����}����[�q^^����˿��u���$�ۼH���.5�9�9f�o�K��Tع��M)]M�yLr���T��{#j�{z����Ex�����g�]� ��X���z�9�23Sm�ψ�z��=�>�H)%�� �f�4�F���5Z5$���DoWa�raV��Q�#^��=���/{�J���6\W1����A ��%��@=MHz*�Sh�����/ћ��M��s!a����]��v�*���I��"=��8N3A�j��M�nÞ7&m��9w���4�]�$(w.� �Uq]��H}quX	lܻ�1M�8|���!��u2�Y� �4�<�Υhn��Khn��F�痨�f)
��u�;��lUB��q5�;:�6Gv�n�r<`F1����+��y���մ��QX�/�����R���h�	8�D��ض��S;<�og_?j^J�0f�Jsk/'U�H�0�eSpY�i=�^�Gm��~�L��ɐ�!��c9p���\
�]~7�_���ul��������m�j��̋1c��cӺ�ٜZyi����Ua��Tť��u���6�P/=���q�������#�w�7��)�O4������R�[��ۡ��<��1*�+:g���v;[ܞ���sN�q�"(��}|�o5�z�)�;f5�o��LY���-WA��zG��;Xک�@�c�׷��{��as��=+����mV���ڐ��j�0���c�� q&\���t6�1��|���t�� �j���|ogP���J��җ�+�3���yS��j�>]an
iX���lG����x�Hד�2���>���_n�v��b~�m���]��L���{�z�͗�e��+�w>�
E�Z^�d�ȃ���9�9�]��;�FI}J7�77e���4�u��<J.v��y�[��� ���ʡ�~[�Hf�5}��w��x��ja]�x��Q��?����8�Iw�`�������V�s;d�&�lD�H��TrI��%�]��`>�[UPz��ï{��F}��eƞv�z���\=�>�%G�T�w9��2�V�ZMKV�Q�^��*�߹1]�h1��!r�t۶tۡ6�e	��35�^}�[��ey%��
��+�#Ч_�(Z�7wz��h���5�������N�ң]+$��6|R9]�fN1���{�v�%s瓳i����W�+��	R������o=�Nz#;���]�gn�v�p�P�UW��!�����5Z�޾z�\&�f��s�a�N���ʙxN����6�9-�����[��Z�,x�e��!�VU�Xi(4n�f��򐶶{Y���fz�SH��皳�cل�=��~�J�<�;��ugn(�ea�j	�3ܕ�P�����_�ݺ�
�m��Ax.�uc+.���=c� ��w+��cW��)�Ԫun㸃����b�Q��&����s��^v����ٳ��ČU��F���B�h�3�v�{��Vp�7<�͡�Ly�u�|f�q�Qoc�86Qr�5�H�VW��e#8�`Tω>��̩�H٭kr���$��sp�l.˃]>�`_`�W�jF���/�C��^s��O�뛝Ʒ�2>[��֜�B�=r�O�3���u��,܄�޹��g2���޻=n�.۾���x�Hx����<�l7��.���OaϷnw����O�����Py�} �|+����ILMuU��{�r�v����Q{{�0D��s�e�����l�%�Ԙ�k�����qU�j��:��ֱ
�A�~�Ҡn8��܌�nn���V����@k�Ҳ�s$�L��W�<���["��U�[��:�ig��'<��cX�kn�S����ʽ�<)��6߳��x�H�ڝ~�~�XM}~�麟�����Zù�M9y�j�1�����<�[���s�{l�%5EK	����=� 080e�*�Q���3vVJ��:��4��n��d�wn�X��zR�=�.�5�;e��3�-�2.�s�Y������%��g��_�ʰ�c� p���vM�|׼�W�������_/E�ѕyg�VMm�3&�0�1��s{V]Ґ$7�N�ʳ��2��d��$��I)���a@�����]vo=�˻�Qº|)^H�v��KK�Ưh.��3�M5Q�n�25�w��^Ҋ�R��W6�)WP��m����:�ե���)ߣ��2��jy��^��58ꔵ*�J��^���e���-��jyt��7m����]�G.����;�stXn���б���z+ۑ��,�0�J��g� ��ߺ�\S���t�T��N�Qrۥ�i�>m�J�1��}xԼܘ$n6�Eɇ�����=��ң�'�7gLM�܍�75��|� r��7�ό�	pp��}�D�^۬�uj�w����^Ǭ�{rAI�i1��]�2�[<�}>�T�c	[�7��S��p�7,��O�Z�	4@�i�dږx�g��2���}�?'/�W���䷪X�m���C�S ���0���95gKp�-�Z���tV����$��_����,tw2VQ��iٜ����!��mU���F%J����/���������TաS�X���� 9i7��[�>]uY�G���h�!`�k�4ͽ.kסά��U�5=�uNP�/w��Q1'�&����#*2u[o����^�sW����u�m��x��=�1���\`U�Z�l	�K��G������b�W6��!�a5
���h�P������Xw�1{��;L�@���E���ca� v�Wӓ��P(z���3y��O�=h�[�"�tC�U��r��Q�y� �������$q�S��^�o*�nعY�:t��ކ��g�䬋A𭑕�]�ҹ�dx��5�v� {o�V���<U^�Fl�@eΨ� �[�I�6O��%r�j8���cA*��3rq*����'����hc�zE��z�dm�T�w*֊v�vQg�כ�bq����$�'��>�n����vN��9z��
�Hs�OV�,�U�5�#�e^<(�4�e��<�l�/!,�u�;u{}��9:d�������L�
�\D�j�8���8�3%����u9}��~~��0TR���$����+;���y�=�&k�[�##ʱ��u�n��wM^����֍of���������Km�����<��fa����z���E��&:"XwU�Cɬ�h�Hw.1��q�~���/�8���p�{��8���XK�f8Dls̲ߊ>��:���%����~�p	�=������q��U���j�q����/�v:+�^4k�c�I-/�w}�s�7��4PR#7pu<��H��*��CW���\x�-��pt�}p1p3��9��Z�ȧ�|�9xUp��@�����=�U5Y�%�����n��7�XM����}��r�<*�d�z���|��ߡZ!U�E����s�O?�<*T���7�_z�ZO>YTN���l}�/�q����3am%��fY篢�ܦTql�WT�"��n�SK^&�8��Nas�NگϹ�J*�w�Yᳰ%VH�s%{К:2��n趬�;4,ŭ��u��JN��a9�xm`Ht�Im�q�k��v����YD$�d��w�hvqT�����wZ���"R#��;�%�go�vS
��t�غ�)�.�V%C�Y{�A ��3�e�����ϧ�c���g̾O����k�Y�;�	��M %�3�HҷPY���+w����3N�����O�����]+���l�S����ˍsbɱ����	���q2�B�9 ����r_=��d�[�pcԒ���!���ffR�&�$�d���;����Oc5��[ܮ����쎎:	�������u��]�ޯqv��]�m�2|�������kА��U,���B�"ק�ϳ�U��Ӕ,���^5Q�3�9�8�O;$�/o6�����6�7�T4nP6�E"�/͜�v���ts$�BV�z�'1t=�5�C�vC�5zY�P�F�U�~;TV��Z��H�:u�Ƴa��	y�fb�H�3͗m���N��QklUќ�-�؉=��|�$q��Nn{}�p�h�Vg�^��7�}?��_��^�ڤ~�PV��U����?�J"������W�Ȉ �蔧�0W�mn�SU���Lc-�Y���SZ���Y���c5�Ŗ������f�������f,�K����SR�55���jjmS��ԵLYj��jj[SR�5-��j��f�,��թ��MKT�֦��jUMJ��ڦ��me�jkSR�5-��j��lԭMJ�ԵMJ���T�ڦ��jkSSj���Ԫ���ԵMKT��jjj���5*�SU5-��mMMjjV���6�j��jjkSSj����֦��jU���55����Զ���jU���56������55i�Z�Y�MMZjZ��ZjU��jjm��V������m� (D !�SSV���ԵMMjjmSR֚����je�ZZ��B�"�$��m����u�V�Z�j�jU� �E �P�� �MZ�jm����U-MZ�jm��������T�6�R�f�Uݭ]m���6� �� ���RԫU-KmT�5j�� ���A �ڪZ�j��mU-MZ�Y,�����T�+j��kU+UWv�t��-M�+Z��[K���*�Sj���ԫMJ��z��6�ԭ����3V�Zek1f�LY��S[fLf�K��շmY�f���Uf����k1f���m�ԫe����m��z����Ykf1��bʬ�j̶��5jjkTŖ�1���j��g���__�������� *�F"*�BH���O�,�����`~��/�q�C����l?����pq_��G�J���_u������A�s�"�
��������F�D_���
�
��s�����3��1���/�����އ���
��t{�7�~�W�n�H�����~�����?�?0����JDTaH�@����ڦ�-5��-R�kR�Z�Kjm��fڕeZij�6�Y�I��M�-�Kj�kT�j�[X��mQ��mEZ�صZ� 	D?���j�[kU��Q�U3kU)�UZ�*�EU3mE��J��Z�ڋT�jKjSZ�kR�Դ���T���m5ST��i�KMT�*�YmKMjZU���m�ijkRٵJ�ZZ��ښԪU�imJkR�mi����MZj��@B*��v~�������Y�'��D@Yd�T@g�?`��o��?o�ϼ,����~�H��A��[4W�o��͛�`�ω������i���/�* *��	��0��N�W� U�ă��#����D_(?p�P@p?��66���i,��&��:6`lT U�����_}����
���'�*���?��>�A�~��L=�?P>������*�
���~D!��PW`ka��Àx'�]�!)�@�Oփ���A�5�=�"s�lT U�	�F=?��K��yË���?dϋ�""���t�*��OD[�t1������B�������e5�n�� �m� ?�s2}p$-�Ϟ�`�m�ٍ�T�Q�ŵ����ʛf���l�-��f��$V�[KSmTͶVX�mZ���ؚ�(-�M������ѥSlM`�����l�h��ɵ[lVmf1RڛY�}d���&�ͫCW��eB�j�Ί����ٱ��Zd�e#[+6�Z�Yִ�ؔ��T���m��2H�Y�:���Hk���U���5�Z0m*��[�4�`�jh���ʳZ�����kR�1����%Zg'.5�mT��m���J`T�WZ�m=i;4�i�  �y�f��]�ڮ���T�p˺�N���nܚUt��X�iJ�6֮��7m��v�5�]*�Wrﻷ5��ݝ�,�<{R�n�.�k�M+m���z��֛a�ݗL�
�c�  ��>�
����M3a��.V�鬛clm�XȖ����BD�lH�i��w��[hiӻ�������t�:3�wm���68;J�E��V�i�����zw�έ�[+���-R���ݜ���۹��[k;uq�ٶ�ݵ�  �+��l�����:�$f��-�l7\m�4�jڮ�;����e۫l4�+m�.�va�Ҹ��\�mvҭ����N�j` ���3Z�L��2֊-��|  ����P{�ޯ
]jڣ����[Y̧.��s��	"��� �s\�$۫n��%v��U����J��;QZ��UM0Kfc�  �����p �Y���5J
8��]���nj���5���V�Tp� $�T� �gg�@+�lST�6��V��5��Ӿ   9�v*�]n(:Y�p�5�K��kU�۩���Ъ�;����Ӷ�vgGn�th�˶����ڵԠP;(�@ �j�5bE����-26���  �  y  _w  9`[`ݭ�  .�� �݇ ht�J  ���t  �9\ A�-�4Y[�X)JU����w�  =π  ��� ���:  ���@�\  � P�;;n h Ki� h[����Ԭ  Q���B̭Y���&ڬ�-�V�  � 4�	� �Ӱ  F  �+  m  L�  6 m��fn�wf�Ӡd��)��%�*��D��b�   �wƵ@ ��� v�]�  �nۃ�
 �� @۵� 
����  8���A��� Ͷ`  ��O��)P  E=�	)*�=A��T�<&UU10 a�JR�  T��hJT��  OT�D�UI� hf�{�������_�d��s.h���P����u{������;S6l�Ҵ�TUʄ|������ϝ����km��UU���kkZ��kkZ��Vֵ�kj��׿������ԍF)L��[Q��Id	.�ݩZkr�.�JH��4�h�@���}�mFo2,K�W�9�\�*aM�d �ZMKӒ`!�u��ࣘ�;�C�㛶@ƌw1BN�v�b��(�X0�Lf�n#O+ �@�Y�e��J������3wi�ɩMxKŠ�ۙ7)�tK�{��*���8��jf�$*Vŀ���uf}�Jۛ&d�j\�i�"�4Y݄���6	���[�.���d(���Gb$��f�O�6�4b�a��.���r�EwZG*�"�7�F���b��6Yׁ%�B��I�y���y������;"�[����V�6�CL�s%m;�GY�XqJ�j�i�Iࡇjz�-ف�eML���(���XI8�eL©,n��KQب���mU������f�D�r�u p�Pj�G�70��M*���Sq"]&����ɪ�TkhT
�	�v�0�m��b��	�N�f����D��pӥS�Xe��82c���ִp��Y�z��K�7SOv�Sԋ7�LV`�&V��m�H�i���.)�P�')<��oom�1,��VYQ�o2D�h�N�0�2�5Cv���n�$����cu�7�2�@cy3�y
t��9󺽗�ӎ��m^��i\@6݉�0��$�A����X�c��t���F6���qRr&�^3X���ژ��D��@��;���h�!�mZ�۸bܕY+K�-e/U�L�
��/,�1xN��Z35�����VT�x��P'�ùi�a!Ymɕ�f�L
�(Q�[�I���4(����j�a۹��h�P%D2�5��R�P�J�b�$m�7Bcc����*���w]��P$�
�MwD�53PsM2�j��ޡR���lGj8 m�rZ5�����.�R�A�B�t&B\�c�7Z�Jx�י.:�J��o�mXsU�5��"�4��a��eͼ�Pd%��x$�U5���w,\�7�fꕻ[tE	�������
�bH3%�d��Q�v�9hR�7Pc�0K
B�T�����e�0|DY�l���dJn�D��%�r�ћ�c�Yd�(;�;������n��jH�,W�O�^�^��i㆙��)q�te?F�g����]YD`�OA�[���1�[�㼃(�٘�Q�9���W��"]��K�v�ҠN[���f;�X*�,�mLq�d�f�V4�ɛ6Sp�N������WKV�٦�u2�A�e�ҝ��#d�$�oo M*"�]h̔,�Z0;3^���&򌵧�t��#Dh` ���z62*���Y�	ledц'��ɬ�0#	^��l��7Tw�Bm��-a�P�e㛺5�2b�$}�-T��V�Bs.�l���UPʖ�%B�h��o��Y-���G���� �Cui7X���ā�P�f�D��+51���X�j	ڨf�,�',���D6t����6�9W��5�F,B�Ø15��,J�M�
b���N*9�X�S�b�٬-Yz^�S��w&=y��v�N2�ӓ���kzޖ��ɉ�ה�f���m�IU�a�:�ƪ��CӖE=��G�����XXXܬT��L���<F�O3q+$�2�<	���\/H���{s5�xe�,���t�a���ՅR�,�EԸ��%nݕYre�N��f��ٙP����Y�Ͷf�ւ�A������K!�v1Հ�AZa&E���b"6�6-���.�F�\,,�$�Em �5��A����	�дe��K4��̽a��Ռ�$��a4p��SAnQ����`�U��GoTNYT6X�t@�htTڼ�[>�	H���A9���V�Z���*(l�X�������L��\-��B�+���Qr�N��-��HN8f�ʓ�c��iܥV��Z���P�I�X��^��uZ�֕5@��8Ve����Q��6�b��0-"��x�����ͧ1^��7��:�_E���y�c&FҰq6�bj�LޣY�B%�SB��6l%��Q����R����Q�.�I����Q�ʱd�˂�Z&����`&�^�E5a�dh��7-ܽ�:U��dB��|C��#V�Dm�v4�[+fG"Vsd�|A�Ts[t*�!n�
�/�n*�QmJ�MU�(-��Y�#c����02�/&�1U� �jۚ��OU�����L��:V���u�[��BЬ�E�bD���Ѡ
*�G[s��;�9�[�)�;"���ҝj����l�7J���Iԧ��y�^�̫��1�*�v��FQ�#'.Ŋ�r�Qj�ɪ�ɩI��v:lkŸA �iQ94`�#צ��Jk�����P�c7n�(�0�f��2ee۽�TGR7��l��)�,���JU}0��^�z��
�Ջ{>�^8�vWr�&6�m��Օxגif�Kxd�{�齨P�DbۋRД#rٽ�%ЙZ^����@�� .Y��&���q2hfn'�%4���Ȗ4��z�a����R��;Xຕy��ly`O���o/u�˪"֊��CV��0��H���,�p ,����W��ٌ<P�����إ�dhkw�7!�I��ő��.�F�{4���ȧP�}����:ޢ��-��b�@�A��6��7)&�+��V��ELś.h�X��ݙFV���Ԥ;�cw^��j�%��4+A�
�v\t+E1�:(�_��V��5���-pC0�o��i.�նlV sr��mL��o�]
Y#�HaF�b]n�FX�)�[NU�b_o))rYn����g)�D�)mlne˭T�5k0l9[U�,���WF��5LvM	�;�2�r]��bѥ�T�ߞ�銯]]%V�����/(��j�N��l��.�5�� �-Q�w��pJ��4T��U��Wt�\(o+�E�6�V4��5�-n8�j�x�TM���735�X�J��M�ؘ���9�.�e'�&ҷE^�Yd�MMn��@�&�,�6@/R�m�BշR�o(ǔw�гM`)V@ɹ��� 5����Ť������rhTs�˘+Em3�ˠ���M�o[�sv KV3%�SZ{�e7�a�j5jږ��7�S2}a=��%W��AW�-}l���fm�]欬N]=�q�˹[ ����R���������C!����oCĆ�le��a��lU�m�"	<F�x��S9w4
�2�<�Z�W���^CtZ��8�aW�ᵬ��H�)���
�UҍC���%�K2^%x��]2�Nb̄	�:���Q<F�8wr�xp�ђ�Nk�]�v���R���Q�#�XX.F�sN"oz�e^�2بN�u�� hڈM:��'*�B��f�9�;>��j�Ok\6��R�!�нR윹�R��6E�"���\�uؙ[��.Z)�����$��PET����Ȱ�KA�v�iHҼ�Q�v��ĴS��؄�D�0tQ���=͗�Z�p^�Ytp%�U-��kR��hR���ye,
�]".���kk���%���� �����K�r���UrWEe���ԫv֜P?��0�Z�B��(�J��=��
�05��˚��*XBV������B�++,�2�z�+p��G2,^]�d1���wR��]�J�u�������v	g[�t�;--T�
3�DY[�XX�{ga�j�ƒ7�b(8�J̠E�-��J�@�!��u��`
'g�E�^9��J�WqLpϰf�-���A�1��pM�1�otC���ܐi���l̫F�}v�"*՗%F�a��**��؛Kaq֭�мݕ5�1�o0�Rv��[bCD�wCM3r��2��7���=hu�䥗Ƹ���8�h�ϋ�ٚ���s�N,"˸ڬ̘en!��I�h���6╯sYH���2�嵩�hU�dSt9):��iʳX�8V��q(�r�Dre7df^�H�6�j�S1e�g�nfV9jh{pRkl�+wԉ9[��@�t�Q��WI\�d	�yv:O��ٖ������ֵK��A�U�)2c���{%��0�%�zX�Y��u�����8��٢�M��r���uoU�op�zZ3�f'v�J�rۨҔ�;�P�=[{���oTXq"��/m��ThVkVl�/���%ԭ�Q�z�)*l�vL�~p�� ��"\�pҷu�TZ��=l�o��k���@M�&�{�L62���ґD�0�lku�WY@����A�)Y��x��0�]�w���k[�nb�@��D̴������e�̚��U��bf�Z^�p���h�ct5����]C��Lv�d��o_����/�6�ĥ#"� 8"B.��t��N"L �7�:{��A��n�9�ܠ%�K0��ҫE@l�0X�Yko�a9JR����1�YX�C�u vŚy�MU��1��N`�lݭd����T�2�	����vebC+S�q�i�J�dj�r�c7+R;��n�f]&�5/v��Z�^V)���!ǧx%X_f�Xؠ�&bj�
���
��1��(oc����řY��)��g*��?� ���4��&A�[Wnm`���r-lmTW�-Qx��:,��ð7��Ou+��=B�T�@�f^eLNkC)�,@�o%�!\�@�6Z1S���u�`���:,eݸ
R3O@$�Y���-Ɋ@�Ļ���f,�1P�F�CFdt^�y��4������%���KF}����\��-ԣhB�v1�5��a���j�]ѷ%�lá�Z{Nan�z�(ID�&�#cA7x,J��d�\�uU�Y48 m��q(_�0��A��Z�Y$��B���ÍLϾ	�h��^�.�%ʭjk6'4�NX��R�u��e��V-�ɶ����	/&����khSx����̣hif��"�!ną7O&͹I��ֺ���*�s4-�ZPY�jG'nP�/a�q%{{R���%�e�Vp�`���ƬM9H�v�\T��m��F�*�&�V�@˭�m�4n��K"���xUm�w*T��x~?6��[&E��Đ��-e��TXS6�A���S
^XZ�R��n�+\oe[7��3xp��xҖ�߂��X6��x*+F�ɬma�	����kz없� ěɷL�fH���hr�˄�M%07$X5�㒣�W[SIL+�'k&�6�����֛0���i $T+��eG�b��X"�"�XE�97@�o�#o&\u$��t]&U�坼��*�*;�PJ��JV���4�������i^�aͻGp�����;3#&��AJT���4ͩ����u�#��U�0�7�����u����A75���jMغ����%��V�9�ʭ�Q�v�U�k��N&�d�A�N�oV��+	5�If����c-��>� 5F��&��݌�P|����[�똁Os�r�$�Y�Q���V+�ym���$Ku��,�
=�Ѳ�j�TaJ���	lܦ�,b*@K`7���onU�jP�;��Os��8�_A�T�$<$G]c:t�����B�1[8���9z�:j`�F�EQ�YqT'mjLg�� �˚��2�k�"�J��#>���d�V��L����\��Xĥ�g0�fK��.V ��0�KW�Px�[�^Ӱ��V
1���֗�dJn$�ժ�t�fMBn�B����X�ӹa�P��&ѩss-d��w�%X���Y�������!��cw��(�EHʛ����iUxͱ�K�����lQ�B��r��v��1#G1�=�%+�	�F�('{��!>4��)ҧ��*RM��dv+E���m�-�q����,�ZFj�L<���3�k>ݎZYQ,4٨"y���l���e�*it�(͘��ڌ��mJ`^�0��s�7���ȉJP8
֑�`}�
w�+l2nJ1���9b�V
���0B�Y�Q��m�y���5ب�3�I�j�*�g84T�X��;W��V�`aSt-̭3DZ�헳*�i���uxA�f6�$���ڽ	ҫ�BK�Xl��Fq��
�7r��J��BC�6�71%IY�������%6W<����P5�)�P��3K5+Y3v��B��aј�朚�)J�R��5�L�~a�E	!An��y0�ǉJ��4��3e�e��-S@�M�Q���J����b�%I��u��*L�q�r�h̩� ف ���Slebn��.�����Ɲ��[��Y���I��#��<۽"T�U�s���={3K�� �@�2�]'F3��8j�&2�۫�u�B\r�`H�߲QtNYb�2J�!4������w�����r��ťD�B���U�C�^Q)9���КjB�Jԃ�4G���r��t,=����`�Ih��.<6B� ��^��Z4b�ĄR�b� �n�L5��P���1��&�k�i�Z�$�gf��q�pZ��,�����!�b	f���W��Q��xY�+76!>w6�@�0\�S�c��9�!�i��80-ןm����V��)�P;��|�/��9Q`�����P>�k-�#̡ì�ݒT��GJQ����Tm8�*8�U̨ݭY5�^*:���Tr�[�'wk`
T6I.�ǃTh&c.�`T���Mj�D�/:u-G	�ZI�|YI�\{`�v��vM�Af�ma;�˄/�kjjJ�70��-��մ����d^�Q;����-Jl�i��5�E�S] �9p]n�s(GTÔ�TR#`ddӀ�OD�z�oov]]���6\]ʨZ
f�����h�$k�-[�ob���U��.��4Ӕ�Y��2�3^��SP�s�����%���Vk��ݵGҷ��Hs	T_S]ȕ��h}�9.�${��.>�e��v)M|I(�NϜl�E�@u�w�N��n�4�yiJܲ��xl�+:wc��
%�R��A�J�tq*k��y�-f='�Y>��޼.���>�c�&)>��s)�3f+�[Y!�a�Ѯ���y,#����r�ft<J{��Mݯ�J��{����ɱ��7�I�HF$�e՜�yI���j�w�/:�>�� ���&�Σ���A��R_D��h^�'��O��n�ܮ�WCz��Po��{B�ϓ��ᣲLNGk0o^v��k@D��z'eB��=���R�9��Z��QD&^���خ�q �c����[��~ސ�8�3�l��N��;�X1�/a��ت�ӺՅ�$VL�ɩ;�d;�х�[��� �MP>�Y�����n|�e�#���C>���*�R+�s�+��-����+Nݸx5jgM4�cg��|��N}3�RʂV�Yz��E����+�_N�H�;gj���y9��֡�>pQo*,�h���8��*��N���U�F-Riӛ��VL8/��T�U��::�;B8A�CI�nA��f�R��'�7mg�B�J�z�D*��Đ�y��b�{�@�_:��TFv�Ւ{Q���)��1������nS��})��W'ɳ����:�&���8z�;y��_*۩�FN�8�z���t�{�6}17Ke�Y�I�n5t����L �m�g'�,ޮp:!����#��j�2�{��\����mA/�\�M��~J������椮`��;Fcܨa����GK�L,*Qʈ��j���g;(���Y}ݻ�L���sUv������d}[h-y�$�x	WAa&��2X�
�}k+4���,gh�������HqNdE��<�nesAx�$���%{=��ޤ���V�-��3@��;ka��F3������T{���H���1��Pֹ�$U��-��^_a$�!qJ�[]�b]3L��T���M��5�dh�4֛�W9�ߵ�����)�����twkk)��l�7:]Щ�N8nX:Dڕ��xٖͬ��Rк��ۅ-c���+x4�b�(q�����
�s�Ӹ�vws����Z{7K6��$�mw73����/k1�ev����5��Lr��u�:��6�f�Q��s�D��]�{�B���dCqթ�]��X�N��B��A��!���yt���k}Y���ݽ��]�$-��r���Ϻ��Z��gg\��њ����8i�\m^1_G�&13e2��U���j��9Ț2�m��0�Foc|7�%u�n�ɷ�'���#Dвv[h��y�We����f��ȹ����s�I�J�P��7\�>�m'll(�����ϩfwר���eT�;�=P�ړ��tTƬ̐��e���j�˸��j��V�*�E'��S��i�J�n�]�:(:�,-Q5e��f"ns�2��p��ǳ��]3��P�q��%uk��R{%�l�$.�|��9]Y� f73bBM��	�D�)��(<�b�\�6��Q�]�x+<����l`Uu;t,��mJ���`��5��8��R�U%�>f'P:��n��w�ȷ��\�-Ь���
���k���6�K�s��]�ul��-jMm�6�M[k��%��QE�	�u�l��b�w0�(\.mL��&���Ұ�,��[Ϧ��JA�����"��$^�f�����n2���v��
e-����2~�3S��T�[`ಅUlc0�HlXk"$`)a���|�z��)t7��6c��WQ���%xj���\��F��h�S���O5֊ENs��('��,�g��&*�%ĝ��OeeUY�4q�*h�N�V`��uؓ/Y��h"���o:T�&>J�UMX�v���*D�lϟX���)-�<�6;aS��W0`��Wr�F��*ɏT���*U���E�,+i�vj�:� s��,�]ns42�QG��;����N�`ܱ��R��a���"�F��wC�WgUPy>.����Qê��#�ʼ�˴_]c�����]`�AN��bҪɣ�+��Al�+t:| ��mޘ��:�b-���t[����\��(s�[Y�iDVf�#��#r�;N[��7����:>$����zj}�����F����Vp�Q��rtO�,��!��U��
:�I���/(��f�m�
O�*�c�We�c����Dp�.�F���5�Uю�I3����g�\���m=�"w���jو�o�.�o�w��s�:Pgw(qR�T��q}�kҁ�
�l�̝M�$:��ٹ����S�j�U�-�����r��o��]Al����X�&�v���ѽ�ZHϜ���ƺ�ٹ*�wr�o*]��[u��"RZ��MB�w���{��^��>b�r�Y�tx��l������Wg^���R��a'&]�QQ8`��|u	�fv!�1'Ƴ8IXj�[g�<���p<uWf�����A�˻>�<�IZ���;���v�	9u�hZ�23�u$�Sh��N-a�f�W%s�h����˔��ys�u�M�n͆���bЧ��E{`wg	��ݚ�A��AW�Y�O��������޲wi�C�P�X��ȳ8Ҽc%� |z�a2��z�0�yM�\��3�"I�Maz�7�SZe+N�`����M��"�� �Ir�s6ڗ+N�0�ϯ�Ge�V���@q��t1�WH��:�N{y�m��5�-�x���=R��\��ʹ�i�9�M�[Q�;���R�0�+Ox�	��u�.i|٩O������/[ΙN�i�M��c�}l��r�us���qW,��uĖSd��O�:���N�������:��:�.����UtV%4*L=7��]���A�]B�&�¬��6���B�8d��/-�"LQm��|�`{�K��§+\�;)����v�n��,�`���Ma<+�5�(�;ᔱ��iĢГ]g+q��U3�&L�@��"Z�O&tO��Y�:e���#�N��F���X�����
օ�����z��M�*.�O%7���z��8��QU\�M�%ț7]�pZr�r������Z9�(���C0��C_%Viv��w�W�"�T=J�[��|B�'hq��
J(ĝ-����;'7�n�IJG`��>ꝝHH��m>��ieY��u���4�	d�Q�.��՚o�s����V*Cvs�螎ih��HLMB��5̺��I��^���ޡ�4k,��,����죽]��f���E���giO��W�=9u��[�"����Ի�xK��"tE`7聭!���)�"ڹ��V9kJ�a�#gD�0�y؇RLu��9���Q��y�"����ҠV��l�2НI��� ���<c��Ηo�b�zz�D]�v���>L�+N\�\�w^5äP�8&,SE�IS�6��z'죴�@�n�4e����Z�>����䃶Т�\�5^��ã��	�y����v�v�^o.�T�:V�R����k�ms�t�hvF�[��Zγ�е�����l.\f�im"9��B����BV���ْ]�ȍ���e=����Tgk�fNi[ӊ���q��"2��� ��h�����b0$����ҫ�9ūl6����k3����i�t,��W)���<�)\/�#XV%���&"��5���\�Ѷ�����o��l]G׮f��B�[�ޭ3��9۫.�Cji���٢�ǳ�anV�����l�����vp���%�L樋���ۚ�U�,V��n˜��V;5�U/�{xӺ�<��gWPY�:���꒠���D�2��=���i6]c��/�"��U���8$��[F�.�tUv��I���9��\����Ms�Z�\ݒ�Z�r��jй�uh�-��ڨG�ꎕ�o��1;�W��̌�`��"$^<+����8��Ϻ���]h<^�~-���̰�XN�N�}�vQ�|��@����&es"���(��a����v`��k�-$�3��ɦM�]j�Lv�L͝iE��ݜ����dҎ�\�y�fn��Gif����v���o��q�N� ��-���VM,������KLR�2�2�yo����5-n��&����/���Jl�{���u֎��Đ��p�]FP�=h.����H�YSZ��h�vF��]�B�m�v���[l.�A<�2��>���陣�[t��z�ek���og^�������m�_^�9���[�`����6uad�t��w)�r���A���C;�} Z)��]��u�b�sq�Ԣ�W�o[���w�ۼw2}+q�C0���s���;/�(⼐'ۻ��g<:���L�1I�Ʊ�a����[*�P�sxz�yL'�R�Xf�z���Sg$�X�Kf#ף/3ls�P��&+��c:�$����;�o�z����_oe�gwiGzi�b�0�QU���uڕ\!�lG�pD��f}�]�Å�@��
�٬wbĞZ��/x�����DEo:k��� �Y<+����w,鋋�{N�����s2f�$�MG��G���a�Q�8k�IdBS�ܰ�*���g^��fc/Y@�s8#Pꬳ�il�9N�!"{p�@��(cWj�r���ےI[��>�+�b����GKa�e�Ʒ^�J;�A�Rx��嘮�#�o8>A\dU��Xz=Z��V���W��ow�i�z2Y�j�ǧv�M)���ѥ��Ŵ��ef|_�WV�8Qٌ�\�9'M^�wN��5�A<�_p�2�L�٘l[�Rk�9�ճW,����r�:DNJy�T��߬s��tkz����;P� ��W(���ئ����J�E�G��c����I�2e�����cx�.��p
�ng:�B�:����	�g|��.��� �U��l��7 &V��庡TFÔ�0�ԡƠl���{�]���lC��ĭ��C��O�Q��S�@���Z�Y�;D�#)MJ<�8x�n�C�uzv�u��S�^�@�PLtv��d�ҦU�x�vQ���/xj9�O4+�V+�	J��6!ٶ�&��M����̮�su�=h��l���O��[ή}��Ky,s�MI��h�ohj	К9�k��`8nZӄ��1��bZ�X+�[aϠG5W:���
�'�;�+0wt����I�׃�t4�����[n�ʽS���A��m�'u�
L:gH���3t,6qt�4�}�c���^�0��dl�9�&�٥[v�А��P=f-ۗJ`�E�h�|�v��2�Ӵgrb���=%�>��Y��n�ك�h��]�=j]���\�:�z�7�jG&Ȟ_���sa�R��o�{�h��\yAI���^�M�a} !v��Co��4��F�t�q7�:d������w%ȫT�U�r:{T�7�fn?��� ��X�E�+2������5>��7O ��+�}][��N�Pk�L林��Zq^uU���
=�.j���u��F��K��H��T�/����+�y��Ķ��Z-[�;Plb����L�q��<�����������"C��ÝS�Δ$�D��NR	�7_6��a#���̮�7��M��si�S��w�܆��f�&��5$�#�Z��8ze�����=in͜Ⱦ�5��2�_������<��1m��d��w�}���GU��xi����<;[�!��S�6RΦ�d]�C!wm����Gɠ-��:o0�E��]����\WHfD_�H����Ah��|@��^<����_-N�D]NXo�,秜���o[�B��U젴+:Z};���ȇ��ѥ_�IY]q��h+<ӣƘ���b���s�inEN�K�ڤ��܃���mf�ņ�����M����N���er��ˬͱ�t+���y'i`#ַ�üč
��6z�P�}*��u{qaNTy�� �;�ic�p����+�L�4��@v�PB���G���٪h:՗�7Ψ�X�*��y�S���wV�>�t��c\��q��Vw<��ʀ0-���LM���]2�0�D���wj&���sz���^$�4���|��u�.�4z��Tоw���;���2���(�>�V�LY��������dd�EtT�X֋�4i�<����f�,�p�t<S�u�]�?H,[��U��#��&�Hб�y)�({9I*<Kes��nm� ��A|�<���[}�0
���"�e���q֥��͕�
i��@g`�PhT�.����k<�<��WCl�F��e��V�6����j*5�mM�J8nಬgb��}���g�d���o��{��t�w��dư�\*�N�c���%n���6g.B���޻r#,j�G��?6@O
�!/�Q��}�a��b����ۤ�w���3-Լ5�Ͼr�)o�#/�c�c.d����wQs}("�.l�t�%������$N�P�; t�|�	�;	����*��T��1+
�6���;ol�沘x"�,95ݎ֙o�Y���,nrʩ��[v�'���r�������u����u�w֨XZɖ�-��v��Y��1v�O�Z0[5}��x�Z���җ�sB�k�m<� 7�91��E%}��=���Gj���I����-ŏ1U�=/9Ӷ�[lI��w\�g�j�W/1�{J�e��#,�k�j\+��k�1���C`�d��4t�2�텰���Tx�Oz��M�8X4��A�7WdG'Z�,��R��S�6��yK6�Vٮ�)l��Ш�X�E��igu��6��Z���i;�M��-v"���Y��P�����s����� ��G�菾����g���K͞>��#0@��j�����\fc��4�5�Gm�e�
�L\�o�*v�q\k����׸�|1�'"�r��ʡR6L��ϳY��>I|c}(S"_%g.��ǳ�m�2�hƵ;"�����)��ܚ7ۻv�].u�S���O�]�,P�[�D'5�,��F���Ƞ�z�9.���1�*�,`��JK{�ބ�M��syž%��N�G���;��qȣXⶍ�9��	%�oB��͟��&:�+݆�Ŕ���2OPY��٨�ū���N�����ca`{�%l=�K|ղٶ]ӭ5��d��j�f���Y��\��T�Xe6	�����C��؉Θ�nb�7�Hm�%��Z�}�0�We6:�m�)�v.�h	Kjf�\_�u�I�=���_Q+���A�j�)����8N��3�	WH��/��+;E�޾&��2�,2�H�=��#ѐ��/��|������mukKB��f�x7Unk�H���fF�z�bQ8Nnݘ�wOQR�x���	�ج��fiWحah��|�4uJuf�j���#y\�d�
g�8qua뭏G0�9��p�;��SK��2��f�;��.]��p��R�EMr�J(��3�
�ʲ���u�;&×�B.0]��[I/�K�uBi~~�F�r�H�i�5�n�u��u�9YZ����o��Œ��"j��B�K����$�R�um��έt��2�)��o.Ŷ3�N�1��r=�jz5���S�t�hi-�u��ȴ��Wi�)9ޮ]ʪ]�,��x�&�C�t�vj�ԈȂ�D���z� ���/V��->�ոV�nʧ���Is�R�3���s� �8ɶK	�ڐwu�O{)Zp�C�L���ɛ��������X�,X!r��b���ś��m��Tip�r���Ԕ�0cș�{�2��+ފ!]��఩S[Lo	�R��O�W�(n�ږc�z1#9�\I&b�R��WY����K�os5��D+���z/C��Ծ<�8�X�v!�'_L��;w��+��1C*⃸�{'��^�i޷�Ȉ���;8�ww���0�0�3��>� *��;�v֝)é���'=����2�������5١�s�v��p\Z�mH�Vu���Zz���5h&����G3�!�����x��jt�c&j�el�qF���t�%ǵ��o]�
Fn+���+��spwO�>�[fX9\vR�܊�Tt󩺃��%p������ �M�|hv�b�<�gg7��H�:h��� ��t���(tVg&#}�@6����jZp�.U󦔥�aܣ]@�3;��s�[ۼ��I:�j;Q̦�N�,:�Xۜks��l��$" �3����l�]�ـ�������1�U��)[y`%�������UŢ�n#���r�yH7�c\9�P���<�JU���v���$�Q�����P��4b�o)���;]�bǁ钣���b�lo�ڀMm?��ٮ�K"��̶'̎`���+d}}��鲎��!��3f1g�B��;hu�}����'c�"����W��Po >�U����4Rg��I@���^�ۦ�-n֐�k&n;�v-��.�w1l�����F
M>��:�ɵڛ��
��w���}N,��K�x�>Zt_��0҉v��ÙyM[�&���GU�V���[Ɋ������9i8:BGI�9�"]t3���������3#�,�.��P�8��j5�ݼ�}�ٔ���t�R��l�q�`-��eh�o�ǝYiuv�K�W,��4�0��p���{`O:U�������shS�i\�iT4Fo"8��Q�:�К���ʶ�fn� �O6E�Kw���!���U�p��K7q�D\SU��eͩ%��nk{C��>ϒ�_G��Q�fMxr��D�&u��rf�d�0��%�\��g�0����]��ְ�ӗR��:�=�jl�t����V@:�m)�[�tͅna��=u���q��C[e2�>OMCǟn��iְ'Y��&�sf��+��3D��d&.��<(u
���!�>	�����1q��Ɍ>5�a�t��M���s{Xc���Afm�1����-�Mz�G7Zx�Q���z�-�MsT�mCSZ�d��ͮ�Eo��<��8l��c�z�P+��(��/�U�A�kbnb|ŊN�)u �y�{V /i�pp�t��6>�i�
3�Wm|�q�ɕvS��M�?���X�0(��F�������Lk�z��T���sG�b��!��Y}���Р�Ჲ-9�K�Z6��q͠�u";���������@�M��ϧi%.dT�o�}TL"��r�F��?9q��q|9�f�y�J��z'k
��X�B,���7� QUq��r�O�]�w(uK��LN��<P4+qv�ʴr�T_Q��h����k��W��ό�-��JZ�{�Dl�0�6x�9����$d�;Fq��غ�hv��N��"�'���9����6��Sy܋΂��a�&E؋Z����i̕��x���X�݄D���u�GsQ�V���޾��E��<\Y`�Х'F2Մ�)J�q�IE�+K�=VB[4L�\t�<�\6�mʔ�\e]��9����:#����\�Q{C�m�G:�qK�t�c{�vяwG�7�!F}�Y���L�b%l����fq������p�&�;�kj:����0j�:���9���h�U���f���5�_R��,9��2�$k��+'eq�l
���d��7Z��vB���\vs����$q�"��8��[�F��h�ؗ�m
��e��m�e���iT8��j���v8fG�U�A���>L�/��\��-���2"K�$��kv��9�y%0����ۊ�-s�0λ�y��l��`pS��.�sw��-��Sv��ڭ7I�*��)F��Z����hp�oU�pf����� �줴�n��� �eMLm��gmqb�\��m�o��Ee*�ʜ�r�J�C����������󠩑��9��fm�Pv�*�eCCd+�&���
h���h�z��HKnʵk�ܹ$��4�
�������X7�����ayh+޴�v$)�{�a�:�=��u�R��m|6q�~���=,�7w�>���Zwp���.�����Fk�G�����)!
7;:������5D��I�
T(��6-P�8Z����%+	
.�������G��\:�aM�M��YǸ ��7���4���[l���q�
��D��Jgo�cg�`��Q �.ѽ�\��m��g4:��*�`��m�/��Å��aܳ�uMե8`x���+�܎S����VF]�Zا���z^!k�a�V�Pg�v�z�J�V(i[�f����9ձ�by��.)���;Or��㗝���<�y�ޮ����qT*K�d�!p�G��U���4�em;�8J]��
F�>�:Vٜ�_!9���x�F����
��=����Տ���@����0lv���4w��.Y�g��i�<�Q�=o�j2#,�gg�0݁�����*r�U3M��%s���݈��'t��cf%ܪ`�B;�Z��ܵΥ����v��y�}8��p�����#6��](����٨e;N�aE��j���{Z(�[�1��#���l�a�Vp��⮨�U�3!Agoj#�����0v̘.���\�Npf��oJuoU���
�Օlh��Ż�n��v>��B`�[e䇛�!�W�N»),��lt���g�z�gs٫Q�U&oʞ��Rh�:f�����"�uj�k�ZN��\lv�6���x�є�����t%*������/P����'���\q��YD�����a����t~	���{W"��c[��3z:�|U��p�8{�φN�m�,e�Jug}4���� �lţTκr�ӳ�p�+#W͛�!ز�Ɯ��W�Ζ.�Y���d�wT���'��f+C2:��ەZ�8�	��"J8�.�-	d �è	�"���yK>��	6�r@7��\A�B��kQ54�l�:��`Aң���h��u�U��)Mc���o�(�7kh]�s���֐���!u��A5H�`K̭��+�ΟE.w����e��ƶR���<K�q�c}�$1��ں��rV�q�5���j<xa�o��G�(t(Z8+%خ�
V���&�NZmV����U15�HnӼ�*,��]I�/��<��ר)j�mG�]_Y0|뽪қ��t`��ˋk�r��57����*/Z�[:}�b��� �z��FIY͞$
sv���!]���ܛ;�9�zA�������
�@Vt���|X+�2�$T���d�Ý	˼�*V��kMY��ָ��M��UWsc�TX�Ҧ��5&Z�u$tcb򢬛��880��
�0s�[d�Qb���V5����c�
f�m-MnML�v��m`�	a�p��6�W)R�J���S�yR!I����QPʽ�r,ʲ�m�p­���;ۮlr�i�pV]5 Y��z�V�1p�8��9�,����gj<��,%tc�//�e5N����;}�zhl��%b��!g�\�Gj]6�Z����3�c'�����cC�MF��kjު;.��r��cVU�v��g8`Ų���C�I��R%r��a�Y��f��F��b��3���Vwk��Ki^G�}�POr��s9H���"�C,L�_gE𭦛��Y�t���3��I,;�4����tܑ����ᗸ�j��;������]f��dm���m���wͶ4�Vp��xX͙7�p0n��⻖�^j��D�w��n�6��Xw]N��F��wVde|�u�],>eU�	���C�[Ƅ��Ш�X��b�$�����e�AMd�,v�/�����Н���,���\�{;���8(_	O��v�(�+�����T�w�����ZkV��3�]ʒ�$��;&`�����*�6����B�%��Oɤ@ӽ\	6JLՋ�[;6'X�7�Vb�����թ�I�/<�1� u���b��b��.Q���2� ��C1Tv��!�k�\�W�f6y p,K�a�ö{I��j����,���T���:���ﮇ;A_]���?$��W���O��(�;��+4*����:�zaDqXq��P��(\�w����BOMI����N���^��+{(E��E��*��;.�o�w۪AuA��6��L1�3A�A"��̇Hkf���n�6-�L}������{�� �%��Q�{�ky�u�z\��
MMY�&��8h`ö�޻�ݭ�.
8 ��`P�[b����Lh���;�X�WX�[KB5���Z�j���<��l��6db�QƏJc��Tgo1N���Kp���ڃIu���r�:��i7E,tϛ�J�M�*p.�N`�N}��q�m�(wv����Ǚ4k�Ҵ&�Tmb���{���6�j�bǻ5�\�h��#k�U��ݵ�A�V�_fZŀ��r8�u0t�5\�F0r���ʠr�:Hvp��Wi�	��c�{G9&ywZ�f=|�(�f��MÐ�\���q�إ͜��@+�1���K�%*����ef�0!�Ne�Y�3��7f.^֧�ãX�&�CX:���vS�5��C�����ȸ����,��U���=�Ű=���纯�^�%=�I���i�Q��1��ӼY֫G� ޸�T\�-��d�.�gR��Kۦ��"��q���M�,U�����;��|qE�|;�S��7�(�iR��W^dy��&T����4Ȧd��^��;�9qL����e浽|���G.k�$�WQd�%�1�۶���"�8�BW>����R�����5��wܠsm�f�{e�X��c�J#Z����}��mت�L�i쁩�Mt�Mug`�d�9/�]o�S���lJnH.�C�t�G/z�8��^�l8���iU@:�4v��Z�͖��)�3J~��ض�(
�J�+w�jY��F���;��ܬ;�:�r3ê�;�24�.�/5'��R�@t���m�7�!Z`��+_#r�ae����0!nBЦ����h0rg���/qU*�)+��a�7�0��֩����sAS�E�ˋhԨ�˞����\hQ�jh��,�}Q��f̡lc�3.�t��Y�A�Y�(���w,'��m�!vӂf1���6���;��*���*h٬5Z�X�����R��^�}׫���v�z/�Z�G ���):yAN��S�Pu����h���p�.���.��μ̐�&�*]k�Ὂ.�챩�����n�gl9��б%���=qQ���z�5t.��p}��ا;mW9���/
V��=���mm��x¼S�\'"�d����:�,�ӊg!2���Ӟ֨Ȉ��r�߸e�H<xs[�B*>�	�*�h��5+���N�h����چ#V%���s�òd��A�}�|����kZѧ6Jy��!b����XI�3c�k��"�p�>�[�S��r��(�\�t=�|C��2�̡+w�KV��m[qm��e���N�/2E"��Igg=�17�C�����T]�Gm�xB���L��D��.t�$�oE��-��2X}xv�;-S���ty`�b���t���Y����7�q���#�B�$]sƉ;�9T%�Ƹ�+H�\��������Џ_wZj=C,�#�,seqL�9��%�i�ʾ��8�}��F�v�y�Z*�L��u�,����B\sY0��'X�ۻ��/9���٦'���
�1�;��(h��uE���4En��u�m:(�=o:P��s;�G����p�E��l����ol�Q3V��}yj��>|>��}���?S��}��7=��Nގe��2R��Cݔ���L���p�ܛ5�-�[���ɠe��Vj���ʜ؄ֺ}��٧y��	aO�+�+]�)��K=�����#-Q��J�/xq�u�,��2�8�q�Yv1:��@k6�\��T;Y��լ,P��<�_��M	Ut�:G����ܻP���\/_.]�h��j�)���[�/�^rZ����]�zL�Yk�E-z���#	^��.�5���3��JgV���C��0{ ߝ4�z�	귉<a塲� "�5��x��D�7�4Q��b�mrc
�w#KD 0��T�'��1�(D���n`�����L���S:4��$ms���h��=��8f�I�CxG2,s�wV�*����
�U�+z۳Q�G�=���f\\YY0D���䐭��s�C$4r�h�F��Y<,7�4ԥr*ۅ�aR�kJ��Q�E�L3�ܥp���喭T�8v�DJ�{��8��s��2���5�V9#Hmj��(1i�|h��������5.����U���R/û;'��Z��Ժ�Ǖu�a��1��J��4���V5��`����[C�Q�6�a�S�{�n��o|��	,i5��L�z�z8:�20Z�|���� L�;Zz���Sk!����{�1O}t5�w5�;�������A.��.:���\nA˝�&���R:�]�;��nk��s.�9��黷4W79S�����s�'9����:������9�:��]���t�77@�5�ct�����������"A���L���%���8�ݝv7Nk�� 9�r��ˑr'v�	a,nW7�$�!���L0�s�ws��w;rwR�̢;�6w]��]�eݻH)�s��݊���$��L�ҙ.t�;4�WYs�]�]�1��9��4��Ԯp�93s���rL���"79��I�s�"���\�9]Gv�u��Z$�f
Q�b�jN����E$���9ۦ�1&M�Df���2H\���q�$|~+�4�]Y��ǙjtKz�'��!��u�v)�4U+�D>|��������m�m'�]���s̈L�b��}�ݚ�]��sr\�G/n���z����AV�@��%�E^qb��x�P�1{�iu���*Jն���q��j���c�˯�ܩ!�ׯuX{����Hѵ�Z���1�]'t�u�IN�{3Y=�8���t~G]я°Ar�����p�2ll�cgk���4��yџ�9��TBq8*7������j~a!��c�.�]}u����<�&�{��Dz�ˁN߀�μ/9�T�yb�w��kܜ1s�=����%�-�*�����RUI�7b�F�b�	È�vP�M"o[�`kuuFu}��=7��D�R��^��z�s���ν�{�Yh3�~��S��> �:��/�9 �O	�����D��L�i;&�"���{�o�C2����[Xs�X��Y��y>p�������?�̑�M��_�)ՙI�|�FfV�7���i�/zO����`�����L���ZX~�����9����'���puG�6��9L�.ЇA�%�y����E�]u�,L�f�8.|H�o���ubz��$�_m��d����_Afq=|�C΀�P�3\�؈�[c��e�͗��y�S����-CEΝ���]����4�B91�-����h�e�$�=�1���&����]�`2]�֨�ׯ��2��� K�ǫ�nΕ�\A�6,�CwU}/��p�a���Rm���b;!ĺ!t������U=�1�iYu8�1�	��IMiB:)�/�u�q�%��,����3�
����h�RI�����p;r�E���
��ho&u�hB�W;H�(h�@�ok �5���C��q$m��>��<+���2��w�AP���z����\��ȱ[������=|�Em y�0S�~��9D=�><!���J0|~\����	 \�� ���%lNVg��?���,��e�6@�mY�[��t��"��
�q�����3A�l�e��N]�)E�٣� 2�Ш|�Ә�>_{�O`?u�"�FJ*�eNGuB&�(#f���cG8s�Ɏ�l}����h�*Hs	:�=?[�����=��cW4	Ee���&�����H����P�LgVHq�mXcI�B0��	�`�i��c-�ˋH��SN,�W�A(�R4�]p��d���+
gge 7�,��f ukUu�3���QTn�*Ac%������5:o��`U����Ml��B��a�.ndu@�V��W���z�ϖQ`����(d�D�E���\԰KS����Xv#�l����#���,�����d�U�#FT�l�F�m�����u�ۈ����r��y��^@������5�f0ٜ/qg��r�2J��Ԍ/��K>D�]�b<����<� _�1�h��!�
Ԑ�����w�k�b���qp��n����4T7�#t�H���vzZY��K	�y�ypY��0(Y�u���t�ˣ��鯓�~/�r}j���V"���b�ߩ��Nt88`�{ɗ�gL�ڍ]m��TK��a�=��T���	�5�|����[~�9%�r��P�-{��
��i�d�2�<�XP��c�>��2)��p�+�����8�]»�A�,J���L&=�>�tb��`Ws&����*���F�1�ԉc2�c����ۼ�u��2���s8;%�p���`#'�=Ƃk{˝���n?�z,�[w.��ײ���=&]��@ۯ#ǅז:#��Gq�H�'�!K��jP�9�����.z��\R��. 6��/����B��8{>wD	�);d��x*���tݒ�W�+�իs7ԥw���>�)Y������կ�h&�=-�����թ�$��JE��a>�����K�Ĩ�::�u��Q��k����n��Ȯ�$���'Y��`�Ρn��˕��N�h5����r�����s�J��Ԇv�3��ŖU
K���K�"O.�լaJ�&IҟtS��:7�p��}=���e
0OR�%�C������:Bw�G�̶>��3wǗ�������dK�mG]�����Gj�
�x�Xu�.�1#!'@>*Ŋ��������s����%�R�nEM`zw2atf�R�!
	C���v���u��O�2�u�:�#&�βp����K���?ECO���ETǇ]͇g'g3"�qh�:��bn>U����.g��W���{��'S�4����7�!��x�o�&V�z�:;(>��u���WE� `�.7dk����U1�/���Ҝ��j�}�vأ����{.�B�3%�6Ĉ����Q:f ���C4č� b��o� %\�l�gF�ѯ����1�(tݛ�{��]��k�����0u�.g�r*ِ�^�K|��n��q�I��1���==Cm��G������7��4����θ�r%�7Z�ʪΟy���o0d�틼Э|��z�ῼ�����<�}c�ω�,���L�y|w�2,�U�ۛ*f�3�[y(��u��vs���v%�/�wd(r}�=i:��5�7�B5�k�������{�Vi�墟�Gn�gh� 5��0�4��f����Q�{�Ʊ�}�5Cpʝ��ã/raT����'NΖ�.����!��.��|E�é����Ge.�i|1F>.���<!��2ȡվ�6�\�ֈe��d�@�c;z��r�"�؁��G�v����8*����sv���
��F��&X�����a[����1�PVh��8xf�
�L�Å�!w(u^�ʠ���o'���`��U�d�QZ�#mr�\�����׎���ڬ%ڄ����=��b(;8_�ހ��כ�5�y��a�;����S�"~nJSprH��VP���(2X48���oc�Y���=Kл�t�\\N�. u'p��者
�(����#�k�]aZ_�b�	Q�%�m:#i^�:qBd���͖���"�Y:�'�M�
�>F.�����U��ϯ�0W��jN�g�QA��u���P�O��SX��x}�2t�N�z��X���&<���l���nS�6z�)�A�԰��
�'��/���UM��}�d�����{4�s��Xq-�)S��՞�����q�D��x��WCf�����#q�|D>�w�]�u���ziNv�:೒Cm\��Emcn����h[�6�i�U7='���(��e���<fN�/�ub?UC��X�5кU�����y��	�G�O�XU;xl�|���R��p���sw���9;�`�)�yP̔�8as�Տ`�M����2��hp�Gm�	G���P%���O�dYÓ��8#��u����X3T��Q�] �I��5oF�k�=�����ָ1���_oqx3�X��Y����Z����+(��#sy6y��;�=t:1�0�&8ks�a��=�i����*�+���L���W3�!:yCk̌֋��^����u����¾׵.�1���Z�Q)Jvf�q��f5�H�i<�(� GHnW.2f8+�_*�2���3�m9|Tگ���B6�����Z"�[��N�i/��vM|�i&�kys������}<�}�l=;�9U�w	hN�-ǖ��}���n������Y*���F����
����u�h@�;�7�	��r�K����Soy�����K������b��ا����M�d��߽yZ��W-#s�&x�����B<1e�^�X4E��$7R���0AlJ:��/���@!�.4�\j(+
��h����^�!eM��r7t@w�	5��'�E�~#�E���9��{L]N�	0��E�1�}b�i�F)�M">\(y�J�@����!��e冖��/}���|��*�Ȱ��H�Qm���}��wDalR�u`�n}}H��y��Y���w���֞��%��Q����劎�lqy��i�vb��qGy�)Nt��oWq����5)PT!�~{Ӻw �&Dr�nc ���T� <gh
���AQ�yZ�Pn�^�;���4T��LX�(l���*4���D�C�9���c�LŇp������Of締�sY����s�Z�5�j��8�+p�[�#�T)�Ob���8�LҙNq�ą���D�c��딕SVX{cؠ�3��\F��� h�X�^��fӦozr��T��D���'L;��������3��'b����,G�6���x��F���gb�r�qT�ĥ��9�4�	�V:��_a�}��V�^�:9�^���E�aQ����L�e��ju�c�nW��b�����>5yP�Og�;6��_n���a��YX�}:	Fq�4�\�6F?��s8����L���M���<���3�^�Kk�A�8YqK�+7�����HQ!�ʛ��&*w�Ү%�}uY��	���b}~��5t��p?	73�[p�RV����B��Ƃ	�=�>��E�+����V�W�_���]+:ѱ�a�WY��XҨ�^�M'�8:Ϟ�>˾����]N����%�\�׏ ��G�`�l�'%l�j��З�e>�]�_�U�d��i��1)W4�[Yz2�B�ns�i���^ Z�Y8��& �sW���ܬ�����,S7w�	:�#��>��V�����S4�wn�
o:����hY�>=t���pj#�_�A|���<U���ǆ���h�.Kն��;y�5n'|���g&Qd��A r;Tȉ=/�l��ڝz�����lE�E=�f���N�Ǿnc�!od�W=-�o�q�Ƈ
��!f,ӗ�UqR4��0Xz�8�C�jC�(u)����S��*uPo�SNH ����)�v�r�hUqptO�P�ɉ��1�36��X��[4�NC�rb��S�|��ڝ�
�G���>�*��-P��U'%{/��~V���c�b���\y������khY	��j���P�7@楂�Y�c�>����Pfc`L~��!Q�
����*\�/���Ɯ��[^0g���:�I��{�0�\������ˈ����+f=
�p��w+V�}���`�2�C��cp�ȝ��Z���1ގr�p�1����\7a�D���ԫ�$�MO
�F9��UTD�K�0K�[��Jb�l��|��$sK%r5c���^V�&��]���&ՙ/eKL�>�Qr��N�E�5�;�(,"Y륙��Ҫy�Ư�ȃ�X%5h�O�\�jzK�����V�YR���ͫ�|3��;��a'�F��b�Y�%b\h�2������eu�9�u�������=��HKgf������[;T�o�9����md*�{Ӳ_()#X���k�U<�z��ʣ�X�>����<s6�ȃ��y{+ӧ�ޞ���Mq��a�ۅ��3�|�F;)?��u�7��%�7Z�÷�W4Lt9���`��\n��dk�8\�V	^�l"�bs<��޺�=���]�y�:�u=��Z3Sꨩ����z�pr����¡9b*۶+:�#ֺ���X�M�;��etЙ;!������6c�#��Qݤc9®㑪~�V�q��C��.3!�gFdc�d��ݥ�	直��]�<n�q����U�A��7��N>����#����Q��/q�-a0�A�\�����|n	\c.A�Oq@�b���7:<Rc.�Ԧ���i�w��	�܉_S��ܚ�G}�4+���	�D��K��t�l�U���^e-�ޠ����w)7� u7�Z�r��m�]|��e������izA/�:ya�}A�cwV�aT+������'�_rP���Έ	�uª���6�8�S��P��>/9�u�����&�7���5t����Ӯ��<��ّ�>;���T�<���8&��)v�hj���X�蕼�uĥM�˕��HDY@��w`ΧYշ�+:��D���OTC�>�@l���������P���2{��6�2��[�z���K�:Fu�I��<����ŧ�2����c���+���c%���:�K��}N���@}��0uh�$\��ՅS����3��X��}��!�=��Cݖ�>-6��>��H/uxR��0+2Ǎ��0�LN� �l�'����{l����/wD�<�m��Қ��M��~�OuO��œ��Cb�yk5�	���/��MPy3��$عܵ�e��ض���U�*~�e����9n0���	�G[X��DF3XTF�jrZ�u8#k��[�UQ�Iu �����u9CF�3â1m!�rV,����=+�>�=#�<Yi�`w�q�jo��!��˳')��^Lh���������c�%�YHAf�x��Hș���~L�`i�G�-��pwZ�������q�E�W���R�7ז���CC�9�y�xf�<=By���	��=[�����c�j�LQ/N� ��}�m1�b�A�ʓ���[5��پPZ5qô�v�|�v�c�j��f73��;�:�;�K9WV9�m���1�^;���P2��:�E΂��qBOr�n��d��r��J����E�ntˬ�-6��0=���4�y�6F�o��u��N��L���[Oz[�z��x��^8�{�S�</r�][D3�3	�U�ܛ�E�+�� �IO��no�'�+��y�t�ɽ4B������n\�uZC(�B2���*����.�Ԗr��4�/��=�;ǖO�@���jIf��j��"#g����_DJAry�m�4�0V�����P��g��Q���!e��MPVa��^(�Vw4v�C7���))�_���  �)ș���Br-weK,�;`[ݒ�)�8^ee}}V�ݻ[�Yug_�m�=\A�x)ܮ��Ke�e*V3TU�ȳ�����_F�ߎ-�E���]k�;@�"ɬ�S���X#�r�v"q��Ӻ��B�ܥ����z���u��Fm�Ȇwy7��,p�Ml�����fVK�C:13�e5],��c�%_Fw%�q�V;sש	V�3:�2^��A���\�N�n�%��쪽���lrho\��)�j1�s�؜��Nu�r���"w+���dk/s!�h�\-}��.Oq��j9{s{�n«�0��A�_@�u�v�{Q :�ly�eʕ�gB�a�Z�J6�i�3�����ޥ�,�5DF�2�!�b9���0B�}]2� �f}��nugN�B35ܸ��e陼�&�2�޲��
4��2�3�C/һk_=���}��죖��>�fv����޳{L!��08X�G�/�E���nr|�Uȣ9��|���з�=��LT볚�u���� �O(0���O{�CN�݀�;���Ȱ=�"(d���W9�陖�.L�!����g���c��+i�WydT�Zά�ʄ��o{X͂�e����.�4Uhĺ� �#�hP5�r_	�dY�=T�\TD}[�h�i�x����xÛ��w2ML�k�mMӗ��T+�i[o���/-�sX�g�D+]{�T_v5�0�u-�-P\&����s�a��op�Q�o���ڜ�#|D�զ��Ns�J�����ƹ���[P����6���F7ς:�]쿃DЀb�U�)��.4��v��tTv��{�H�|�2��;�4�٢�˵�q�7Z�w�M���4���o�`�]KmWc��*s�2��W�)�VQA�R%����txr�#��f�j�ź1�+jdA�?k7٫l�X�6T�Դ��Y�s�]��IE�q}����,�\��*����z�A�6(�8��X���	�h;�J�3'P�Ά'ֶh��Ěc��lb6�6�`�yAE�e<bѭ�6�����w��t��zrE�����[��e��5e35�$�˔�/J�]�/�8�l3�X�LTi�`+N�,!�+���ܭ��v�8��������u�.�$:��4�M6C�ts��d�����h�t�&`&H�K�(3��wnhr�(��2M�q"�b\���C1r�JL���ewp�u��@@	��r8i�e�7ws
���]wv�v4DIADD��I.���ngvWw;��IId\�wuΉwrc;����H2)�����κ�F\�(nu;���NGbg.`���4b�7s�X뮝ۻ���`��]1.rL�r�L�����FĔ̻����4LQ����. �v�#.�)wv�n3�s	 ]v�$(J��&��&':9r���su,� �I �R @?RJ9]s��L�Ũ=�Ɗ]CR�@��������k
��"���A�Q��}&��������F�|}�-�`����������/?��߭���h/}���-��[ߟ|�O�G+��/�{�گK���z��|W�\�^�η���r������i���{��[�|\�����oo���D-�Eo���T�Z-H��i�+⿗��w�<ſU��۾���W��ۛ���~����h���ץ��
��p�5�~�OM\�׏�����o��ܮo�7��W���h/�>!缶� �&n_F_�u�^��H�+��������F�}[�ߞ}��{[��^?������s~����>�z���+���=z׏��W�����ҼW���Wwx��.������y�(�?}��}^q�>�P�����p�^�����<[�/|�^7�o׍������^փ^�u�^���j���|������W��^?o�m�^�ss|>��ޕ~.m�}���7�r�޾z�[�����y��}�U�Q��]aCu[�翞��ww����6��n����������������^?���o�n~�������o�{�����m���-�}��R[���>��_|� Q�/��� D#�������" �"'ؼ5Q�J����w������_���r���z��W�G�1}d���� i�|����Q�����[��+��-�\�m��O]�W���W�����>�����z\�׀���"�D���X=Y[�����H2	]�2>� �F�+�@��x��_}u�o���+��/~����[�~o�����������ҍ���x��/�+��J�^�|\�ֻ���j ��� ��]?X�,S?DH�"����_��1ݳ���Nf�}u {�!��!��������w��_���F���� 8������d~h������!�o��?o�k�����o�_��ߪ���x���x��ҿ7������1�{��I�qz�g���G�H��DBU��~��ߍ�7չn~�~����\���yu{[�_����Ͼ����ۚ����2(���$�����>D|~�H���| i#�L_�!~�����Y��"N�������3���W1w1� } F�zo�W���W￾_U�W.m��|xߍ�^*�����kA_�{߿?=W�~-�����Z�o������?W�z[���m�ﯾ�/J�[����v�-�?B��A��|���*��;֢�u#����Z����k�ا#>�� pJ�GM�oe���eLsfo��؝b8�#Ì���9�#|k�3��D2̏VJ6z�s��'����f`u+0�;e3y"����jP5=��m�ۄ�ޖ�5�n`�3i�I��{C�ϯ������(��ÐmU���h�/��\�������ţ�_�������r�U�����W��}[ڣ�Տ���~��c�B>��ޯ�+�����|������&���Y��n��~������UR���_+�m6�W���m��mrߟ:�芈�x��� A�G���s?}�>����6�7�~�?<����ow���ͷ��~�u{ޙ��[*fo{d�1���H������r���^��|�?|^7��~^�{U���7��כ�����._��k�2�����������;�O 4��k�+����\߭��~������ǂ>�b�DtRK7��,����8}�Sڌ�A#�<^��_�X���߼b �6���[��~W�������ţ�Q����+Ү\����צ�o��剐�����W�??,��>*3�d�*���\��>�GЀp���;O�x����Z���~*��_�w����^���o�=���>yk�|_��nk��үw�|�7�ܹo��\�zn_�QQ�h�<G����<~�/�Ň��n��7ʨǬG��",}"=�c�b�^�}��}o�}_U�o������Q�ϋy����E�o�r�}����⯋��~��׵ʹo����/Mx�>|�^?<�QH"����g�~�	��ȭY�ח�NWzz,E���>��G��#�����x���+�_�������o������徯��W�߾zU��o������?}�Q����! Q���[���P��DCv'���}B!����O����vto��ȁd}�p�#������*�{�yzF��o�����K�������-�\�ׯ�������o���=��~|�����ޯ��}�|^��}�x� �������""�[I��q�;^)u�A^�b(DH�� ���~��!��D����7/KF�W���[�x�����_潍�no���Ҿ����/��zU�r�U���r�U���������|j�"\�G�>#��B�|�\`~{ʼ��P=��n�8�+� }�#�=	e@�z���־/����{�\����^5�c��B>�����!��>���������^5�{^>5�>��{�� ��
�P���2 ���`��6w��jC��/����-t��*Xz3b`��6z(�D��p��N�l0���ڞ2P��T�����'��t�׬�}Ë��WQ�a�ꅓ�T�nN�%k[����yX�jV]aQo
ͅA�6T]^թR�J� z$} B"��ڪ"��G�CG��u DX�����6���^��r�}���}]�m�����z[����/�߯=�Z�_Z�<_�~���h�����{[���m�������i.T�;��i�Α��x�Sf���^�������~�����o�zoM�����.�}�xۛ��-����V��k~��W���Z��_�r�Qr6�s{kϽzU�r�m���{��֢�U���߽F����"���k�盋^��;�u�@��>���Dz������B(E�U�ԕ��u��V�߿�^���_�]�|��W׶�������ޗ�A^��=k����x������;^+�Dh���=1�|F��.��謏Aܕ}�o�`�����D!���G����;�~��}����}m�u_��J����7�ܹ�[�����h*������ZG�Q�� ���<C?7����G���}�ȁD"���/j�����\^��M"|�}#�"�>�)��&ܣ~��h��r��������m⯋���_Z�=����{|W���~��~o�W�z[��_����W76���~y�D`����H�鏨G�D~�to���7B��PZ�$�h��A}MVz_W�E��矫x�o���k��5�m��o��ޖ�:������׊�.o��^7���5��W���o���d|���@G&k��O/����T�+�/�s"�O��ة�} C���}c�_~�^�._Ϳ>����[�\�_߾�ȋ:~;7�}f��_�g�N�G�~�|�?/]�h5%�����֏����+�|W��ߞ��5}s7�y�G��ԧnn��Ύ�_4$�!f=F���k��U��o�|�O��׃+�޽*��_�sϟ�_���~�W��sd��$}�������V�@�V@��75����o}W��ۗ/j�z� ��权 GM��~�6G����b��-'5s�����/���7��/ţ�#`�c�Dh�FF����~�!�z�Ӳx���"�An�Z���n�$�P��'+ ��a#�,`u�7i�
wJ��	�7P�S��Փp�id��t,���Dz�ռW�~���J����BG��Z�S��8����O'�c���D��Q������-��.\�|S�ru��j�1N6�e�+���By�f-Sk����:c^����qVa���zd��nÃ��RZ��Z�-�⋨�<*��]�aϠ��.�P�ο��([s�M�ڑ�E-�uI��Fc�Wj�M���8���.��P֞����եڄ����lu�龺	!HX�\��E�jߜ]B@ҁ���=܉��F"�����J;��A���C�K48�*��hF��u��e�U���A�< �^X
�HɆ�3�Q{D;��.��BnѶ�n�E_ދPI��&���bÁ
��͛�'@4s�Y@E@V@�j���@ﮝ��o�9��Ѝ͡�4}����>^�U�k%�35��ҡ_Nt�f*-'<S��]�TF�����7;�s)�u+/|R���^���m��:���
g�5H	�i�1z�TB��'a9������R�.H�R�6�J�G�/"^�1��~0�LN����k�Ȝ�G�y��R�[��̣���Y����ͯ���̘/�^B�O�?�r�l��i -�� ��4��kR���d'��.7��zC}oM���cz:Őy�u!���O���Gʼ�Q��U
ZH�f�#���3o�N�u2ևTj���`�ڗ8��![���!^�Z�=;�p|���H[i�01J��,��l�{��c��p�ǈʮ��DЧV��)J�]2v����}�+}�i�����[������qȐ��Ƣ�Bo;���)
�#�XeC.��a.~�+�NP�kڞ9�j��lX=uZL�UX7�[=zƀ�-��?U�|���!+�K.ͧ)��~�����hK��>[O4_(��x��W	��2�U��/
�K^�`[���L�z��_i����9�8��J����"zy\$�7��](�<(Bm
�!��[�&��	��w��/���{_Ӡ�9��Ҥ'+#��(�v�!�S�����	��@{�U"�JT��eB꺍v`�wCi=nR���H��M�.;�P��:�b��n��TZ��<?h�;U��@w�za�	\n��*���f9�YwXd'dh�������K(i�0��u�v%�uU�gQ��;z��[�1O��O}�����.
�e�ϥ���Y�`�� X�x���ܚt{|�(��#޺F�8w��֍���u��%N�a��=���-�پ��`�1��r�,� 5BG�_ʚ,F!�u㔙���m4�:��?��Ǐ����ږ1������]rU{�+���@��@p{u�Q憗m(k	641���e9 �&��dPӬ�T���1[w� V��0�u�1h*�p���v�Թ�\���@l��Ͷpq���8T˾���O��N��[�F����S��l��2h�ٕ�I���,{�S֬W�ܶ��,I�0�&��:�A�Λ[e�Sw��JQ�S���}QR!q�|N��B�r����H�y�9>��^×k��Z�XS;$�!˨y��)�∥$���%���WS��<ɑI�+�I��w�Yt��� jq8�<�<�jJ�� '���d�9~��`��h��.*Έ�?6�t��q848�|�����ke{lg�0��e}��kynt��v�y��a�Mf{Һު�$[,L'��^{2��N�{\p�F�����F�e�IL����ם-���վ����OONo�&������ל��Q����7 T�x�puᾼk
2�o&�Of�x��B���e#�X�7\�ALb�:4��T�-?T	��`:��e�´<V�7�޲��5:)�nግ��7v!�+�Y�a�<]�s��X�D��`�`;3�Ȣ'm���	9mNV�r.�k�����F�$g+¡~���V0���ZD����g���H`�5�m�i�́��1-�WӰk��p_�()����f���cKG��)]���,��i����O`���N�q"��w��+ͻ[˨�\���/c�h���+VCv?��B*��`/���Cos0TLχHK9�p��S�UUw�Oz>�Z{u��ƅ���Vz�&��o���`i�+��Mݹ(#�eljÉ>���h�tjǨ��/R��s`�*{_�3�l�w��Lg��g����lGX9s\���8�\HA�9��Z+'�Bi>�H?���e�\-���&9mZ$��mP�w-��ҤŁ��y�J�<][�ŷ�%U�'�OӒk
�eJ����ܾ�/��J(h1�b�Cn�}���c8N %�`�jX�ȩ�Nn�B��i��s�xJ���=�s݃��(X�<��Ik����):��6S�Y,u�St�*�[���,��� Ӣ��p������v]C��D��J7��8"�^[��0J�Mr�{ϖ������ĺ7�c�ї�,��;2��Ѐ�U�2���-)�on%i7��W �H�w=��xI@�Ԑ�ܩ3�a��8P�s1-nԇ��R +41�սȊ�K�t좜�_Y���;#}�q����j�J��j<.%~2��
���k{ˆ͋���YR�ok���B<��Ab�3��k�NV�R�s�Ϊ�]ۗ��<���8 4�I�v�@�d띃]0�Իe]�k"�b§M�Gz�.�F�g��5����2�K���7󌟜Q�k�����vz#��I�	聝��v��5;����a�4=�������O�/<�$w��7��ǲ��V�J2,K��E�r��ϝ�.U�輎Tu}��}=� ��x�)��`�7�k�� lC��!�7��_�U-9~ct�',B*��؎ɤ{>]DE��`,v��<=��Ѷ+���..Q�Ƈp��F1�K�q����ghUe���B��Ku[�%f�@p:��eP��B4��l�U�%�������to�{\T�6\�ژ�۷�"{��2^ �rC��{�´�hn�.�Z��P�>+���)q�g8m���o=��\!�W�	��H�3�"�9-U��#�ځ�B��y�|��zW��e�4����Lh��N
���+)�7 u|�X�; !��.�co.�rroS�1���k9�r6fK�9�������!�n��ßjtG$�&;d	N�N�~�}u3���A�%���z�K9����]��	]�Rx���e�5�3�T��3��{@@-o��yˣ�*fwi]��0��bq��Tv���3Z��U��Ⱁh�*���=6o�gS�بwm�S��hj, �:�KZ��`Gfw&p�v�z1`Xx��Ṍ�h�%�t��{k�'�f��������#䞍;3���Y|���ﾌ�KB�����}����3��@������VN>&�_���*�Λ�~p��~[��Vv�.�#�m����R��KC�k�oP뗂p�,A��@�D�oc�����W)�@����m}�/�)<5����k�Y�K�?����O=�P��Ú}�s�Z��y��!���u���u{�41uY�|���E�s�Y��έ���I�����_Q"�C���M
˕0=;�q �2�]=j�8���I��d�dݘ�X����[��9��h����뎸ɝ?TYc���2�,�7�j�+��s��_�Q��[�VV��[.������k+ R\M�1���&*w����&8>��_*�)�3���z !�h���l;���?��b������m�7 _5\ OV��ͤ"i�8�����u�Una	�UFZӍ� m�w
~P�h�.��h`R�`:��G��]��X*vd	�Y1}���X��q�qϓ�C��=D�Ǔ�E��?+>9K�~�ʰ̋��ﰃ�.<�Y�yb�	��4"��W.l���^�g��{\4�֑�R�I�K*o��m���uq��3T P��ͫ5q/�	1�+�1Tڳ�X�+8K
eK��y�D�k�=�ձ<�s���/;:�u�����>Z��Z��f�0�]g)_������X�SxRi{k�'��L6x�ZdBvF����R(7R�C(t*(#w�#P0*���J�<>Xk��9��K�\�����Bʛe�.���ȷ3��0�8���j�t).�Z{�nh�q�6�����/�zΠGM�OP'�E԰c�Y��N�F���wt�2VmbD�2��Sc���C΢��]<z�<�P���Oy	�HE�a��֡�@���f//qԣ�C!�ʫU�9�X����Yjcg�1�,��88YU,��u��2+���K����tȼƜ�粽��3Υ���W�6���%�������#ke  �������6d�L�c#�#���	�DJ�H[^V��YW��~J�x8_���@NO�\o2h�l�����ݘ���*#�T�ұw5AX��Y��U^�n>R�n�Ų��U3��X+�^gJ.�/37z��Wq�H.��	���-%�Mx�{�ǜp������r�*���ڢ3j�o�>>}����C>^�7�Q���+�uH4c*�D�|¤��u�]�e��2D�I���2,?�Hp��l��XT�s�7�6��Z]p7��Dd��\Q��a3{8T��eA��Ӎ�]@�㪍ש�A&g#�^T��`�s Wt����J.�cEq0]wj*V�Sc��AE����¤�r56WΆ����8^
I��OHJ��M�Hk����x�����[g�L��C1��koN�TZ�4�ۺZLSGIlҙ�n���\��̵�GV�6������=+����P��*o	2�"�u���B�]˹���|�=V��qtbx!jD!��
X�gq=�A��w��������´@������i��ҍQ�ۻ�6+ݬ[�O��L�;�
����t�%�����bZ�cJ3����/�Kz�H�>�l\��X�z�8U	x���YT��tuI5�E.n���h=P����)�k�9)n���Sۖv��z�\$Xϑ�6\�n.S�v�V+)$n��B�7���nj.� ���z��A�N�^��I|�_>�Z�f刺�.�w��;H �|vԩ�_J2��i���_r�)�*�#�Ϻ4�"66�f������[�p;c3��;�����+�8"�.Bx���Vg41�2�˸셔�u
�$��b�x��s�
��^tPoV]��½܇7�Zeb��М>�+�M���8r���������D��j�����d�	\Ms�殣M��j$$4"�$7�v��Xk#�,�v�j2.91W䪏WI����Pn�Ҫ��O����(�f����"%=�4���nXð��z���,gkX�EA�Z�H��NCp�N��VN*μs�"Ԉ�	��J�#afv�kp�?��C���i� ֋����RI�Z�N5,gV���Jr��Q;�l�}���^B5�uQ���~G�h+�V�]���KZ鏞1��B�j�C�UᏧ#ʢ��V�S]1��C��x�1J�s]�Қ�]�usƜ嵙
oRy�Q�ZS����pD'kF��7���MV8<0�fV�]mܹx�X�V�s�M���au30k��[������ݳ�M+)ԉO�O	�Ph�&t`����MMh�v�s�J�5y���/�ba�z��;F.+�jۛ��6T�T2��'JM��Z���3��WDܜ~J�Z�V��H���%��k=]��9��c�ᛋz�r��|x.u�����й�M h����ō�N}�:��?��WT������bo�m�V.�Š5Hq/p�Y��R�b�-Y����ז7r� �A>T���E��cXp\K2��o��H�|!C%�]h��� ���ް�KԦؾd3,?�&�"�TX�b��X y��g��{��-&��]�%2��bYJ�ɸ����~F��3�U�\�.s�Oi��7,�skӂ�+t;_P���Z5+�9e�XT���H�8u��Ҿ�+r��A�A�?Y_$1wsA10Ѕ�ӻp�I���H���wM��L�d���`�Ha&I,̛�4�"���&"R�G9$�7t�s�7$��`����*��D�(�ݺh����(�����	�]�9�2l��f�ѠD�H�ܸI1�2�۝!���ĸna����v��eFR$�"��%ݺ�a2`��S1t�@]�9�I�&Ҕ
&�)wp�4bP�L%� �0�.�3wq)��n��λ��	�S�
�D]݀���M%3H�e�FT��u�JJ,@��b(K�i%��#��T����W&>�$�/t�W]�ee�V1��B_-��o��A!�6�0Ži����ЅMq�������s���vL��JՃP��Z���_\W�yO���k<xJ����]W��..���ͪ&ġ����D�C�g����F$0�Uބ3�lt���ѥ*LB͟��R�+�s���ζ�R�|ޱ���w��P�D3�3��^/1��	cw5�-��17=Ep�������פ�{�ߤ�%�:�
���7�Oa�Q}��GJv�l�ˌ��멆n`��H�/Y�:�����]�,穤)AR���3w�K�Q}���Cs!�{'
�yd^)�������=M^H+2�Ƈ�
���F�P��V�,Bo��4zT�
�=&L��NY�ܚ}��mGu]��I\W"��ϗ�x��Ui
}�Q��¸��#���0����5�ky��"��x,�>ڔ�_z}J�OBkgڶ�9+������rMaB���{�r��:�������ȱ 7Н]���07Q��>���uY��e��rM��G���:����>�b��B�P��.n�a�"�'TÅ�h���j"}^LY���OuǦ'F��;�)s�7��7S��|���0G��N��z2�!��e�����2c]�y�8v⚥�Aq����N�kVڥ��0
�1�Π�b���_k��;o���ER	H�	Y}�(Xw�\��:"6 n�f�)��Sr˛G�+:X���}��W���2w��wem��j�icׅ��`�����˨w�vU� o�2Q�������r�t*{�-��&z���I>����X����t\�7�F����U;������Y3I]j��<�b����+~��o��&���t��bz�/��L��( ����zR�!ܣ;O��Y�Aq�K��cyhw)(��|s�1b:�f�K�Q+��v��~�=R��m���ێ����12$&�<7��P��;������m�2�@�vRQ��u�o^�����Ҿ[{�РБ��bV=�"IB*5K�p��c��tƋ��gmWY��*�RﰄT�8�Z��_�Ux���Q�;��♸�YP�)Xz4��鿓�"�M�c":r�=Uf�Ot�u�W��˦f��A��@=Ȫ�e�.c�F/�(uAc杶a��]�"4��lZ�)�{�'|�پ�}I����='�SX�� T�I'|v�ʼ$�����W�ǅ�"Fi�Ǜnry�S�����rF��#M�&��-:'��,g�t;7�1��(9�!�6sv��5uB�8���Ì!���.wh�;�k������S?-Ӟ�v:O�-��X<"+��F�fU� ٯ��Z�����v0�Nۊ�͢���czl�;�;��!�x]�H�_bU7�Ӹ�u��g�]N���J��o菣��8�q��EK���N�B.Y<
�Z��"EY�b+����I�r�LM.�yDȩѭ�B�aApb�8hJ�i��� �(��y`U�w \��?�s� ׃�v�R�-v���#åm&"تhD����;�D�-�$2�(�� ���9���Լ��k'8q+,WR0h���gl����
O�)�]f���ų�N*t��ΫC�Օ�ӻ�U�G{�͍z�R����O�:5�uv��W�$]j��aT��r�ǆr
�;T����9V��[��W�r�n&1{�5�o�(��[^�^����5��&2��;d���Z�g/d�'�2�����b�<y_'��\scd
��h0��B���4_:�y�=�㮤��۬�� ���6�	�([.�x+<�;����z�ÞJŝ[T��+s�ƃ�\��#��z�?{�*pߐ�f�1�n���9���P���t�-�2������ܧ5�$���h=3�RU	�dΟ��>Sze˳i�gF;��;1n���4�I����n�.72�\�"�Ζ�H�=W5(@"�+���]Њ59Ǽ\L���GV��os^M۷Z����P�#N�$���.I_ 3:��:8�S%۴�}|�G/��)�wj�*>�Z̙�R�����U�O�m�ͿF��^���R-/-����ܬ�z'żG���| ��ON�����Y��{����|(�I����*��B�f8;�+U���S6!��t�R:f��]sֈ�n�L�_سo�!��w���|�큻&�t8��o��\B�8�ɃW�1VaN��.f���%i���'o!��:t+��!#Eʀ�*�BK���r�B������{�F�K��p��:H�VX:�+�M�� #,}���ȱr�b#��Vm����PR���ً�,Ւc�����^�}�ބ`���4�y��e���M�pD̅R����P�Ѭ���f��H�%�07��k�lq�uT�rm����8�g%(2�xl�f։������,N���F�<v/��u{]P<-�����<��>_{�4�b��&��$��D�
��+�$T&4`(�H�ȼ1��~4���o�L�zj;��$�ݥh�ڭnɀGL7ڬ3^'���@*��XS��G�rSr}��خB���b�)>y-��ٱ!<�e��
�4�N�x�S����ũÿm?V	�m��{a�0���v=Ӯb�L6�X���6k�H�x��уQ/�t]WA�E��ڜ��o҆Fõ��V'���v�3���������'����!R���:4����*����Y��m��=�}�h�^N��6	P�H��
���s0�5Re ��d����>����=���n1�B㓒����}ʪ��bt����`�u���ڼ��/��u�>fK���D����*w���1�F�*9P��BR�h�יq!ٍh=z�f*�ƽj0cH=�"ܞ���Q84_�莢v}*��*��a�X~��=(:����i���,�S�&�fww�-������Ⴝ�j(�o�]Z�8:���2����[?jܽ��jW`�5�,<�	�H�YO��/۞?b�b�S�&�Ǆ����p�_����a�_����b���Ӂ��.1�S���P���@�ʳ���\�Wd_J���գ����Sc��8�
���
�_���Lp�K��k�89��6]J*�3�q��w�<sMN��|O["��v���N��1����?���r��$g+������լ#��ls[~�����RVE�A =;u2"J��/�s7����5
·ų!��p�C�3�/e����4�`�ܫIb�W��[3d�)�0YS�b}����WZ����!@��u����+9wn�����cL[;��=i8�]Z�vj�t!��>�`UI�GF�2Fg0������|6r���j�v�[C��L)8c:7#{#��Yw����g(����w�T�{)�Y�/w�����u7�
b\0^>�����h�p�6ps��� �뭞������ǧ��w����e���|X�#nj�cg/0�Ƶ����o���$G�]����&,�N���x��l�V��u�c�~T���;�Wo��/ ���'�u�|a~f����b�D$��̋g���,b�Աە5��֞T[��qY"�s^9)�ˍq�ɭ1�l�ne��3��L�+�2ÿ��6o�މ�3���H�<s=�"ep�J�3��mV����X�J��⓪�~�u�:kQ'3����������Im�.��Qi�&0Pp8e:�g ��:�5jN����j�k��M~�P�^�L9�tꧺ1����.��iϱH�9�D7�9W��6�7B���㘡Q�@�mHz֧�m��sU��ue!��H���19���<��jQ�V��yЄjC�C�q����o�m�vթ��m7@�q�!���iϵL1��xmל�[3ݏG^��:��:W�S�~�׾���(��!&D�㚱-#G��c\;�4\J���H��tE,�RERw�MQ�ѵ}�I�5XQ�u�T���r�_ZjQ�U�1��_St��rUg���73�<z��?N��P+ Mvg�Q��
�]���ᷕ��U�]X��nIː��4����E)Bm�������ᢱ�?F�I���Q�:�L��:ww\�k?��  S��/w�P�/�0OΩ3��P�;����P�����ڦ�8�0����i7W�֔cn�J���F�q��/��$n}*���ph��C����7k�)��\+�!]L�4�:����z�Ӎ�G�����^|��[�n�*��sݞY�+6ʥ��{V����C��}l���
1��&G�f���	eT�'C�d�1�Ӯ�G6�gyͽ�u��|�/�}LE�gA�N��.$���d�:rH�ӑX&բI;9������{���=�-#W��N�,r٤x�� �G 
ٺ�k��.�0�����/#V.�Qڊ��p��V�d��^��	��S��l���|�(�
�x��׋M+��=�K���#
,���b�ة�%q�3_iA�,�Tq��$�e`NoC��!u���	�ۣc�@�hA%�|b����b.wP��z��b>&�?X����9rvSk��究EB��=9-��)��-Y����?h����,<<4XV]������?js�h��ђM�W`7�p�c���g�5@;ye^�%��]�Mt��B��t	�a޵D���)��\��CXJ��=B��V�\h�<Q�X���n�CI��W!�//WA��M|��:<{OY��;���$�?����d�:3W`��܁�8�D�v����!9p�w"%�T��������6�W�gО�|���k�Yȱ��lV��%�]�nOd�n�ͣ �q����qB�u�7z+|ք2����
�~JŜQ�	���O7����U#<<��v��qp;��G�1�d���8����Šyq���u������׉7wy����ԇ&{��	�P��?o�a�2��˳i�eqva_fi��J=��}@�ܩ~�sv ���|(���f����Mh��?��L��{Y�Yљp�
b��+ޗ�y���ث�d��~�Q�`v�p�p���s�c��K]JNJ�lsg{�J(�A��W�Â����\1�m�Y�����B���y�Z��X�`\9ƻ�V�9p,�/j9\Ɔ6"S��7�� `�i�3p�IF�X�{;�┠�{�����,�� 6r�6�bc/MB�U�����B%�h?�#���g���V'�E���}T�5��-40�g�+՜�{Vb�.���}_T|V�!eM��传;@D�7�i<�x<xZ�P�k��X��qع�ɡQ�]�t�����3���h^��E�8��Բ�����Ƅ�G׷����z����|)�O���\�۳B���[�x]�c`=���T�#��P�#�i��.��e�R�%-�Mv~������5n�
b'6�'�����K�%�4x�_9��Y
���n����amS��;9л��qr��������%s
�d)����C���8���/O�%�D9��xK�Һ��P�'!�Sj�1p�bÅs s�gZ^^՞��K�T�u���y)�����[���2c�1̈́/fq|�=g��>>�>��2R�rUyﲵ�uz"p�����JKr��AmK�(��-���zk�Pc���8��3��<�P���յ����[J�
��=�'_4g�Y߮q_�Q��Td���'����fm�����KG�Y��ݽS9�!.#��W�<�qv�B��<�'Ծ��������^�����Qi-�Ϙ�G�wxpx�3{j�]�Dzs�Pi��x���	��g�='����v�F��{��[<�킦
䉘��Z��<��O�T��j/�dR��Sf��]�+x��dS{Jo��L-L���Q���Օg6�:l��\Px��nS����ӱ��]�|���������m��I��!�\��x֡&__�RYx�s�s��ss>-XɗS�T+��ۋ�O@�f�EU����.#j�
��]d��,��}Y�e<IL�p{�#�*�nV:C��������qٞ��� ;��c�Q�wb�������n����ܴ��<Pڃm�Ë�삜��⹵7��qo&�Ƹ�W�'�t���_`�ّŶ�܀V�18����Vy��\��Lu�+���m�Ei�+�*�S����Ys��H��-8�b��+�59-��Z���/���ۯ\�1���M%����e�֞B�BQf;P�t<7�>P�i�{1�E�Gqv����gG)�o��1>�\=��:����rN�Y_^�YqT�}}�6سMf)q�����U	8})�p�1�eM����϶n��6��x�/��0{5�<�Qx���g��Y�F�jn��m^�W��.3_m�4Ѭ� ���'}{��/'*1x�e�ΜP���B\�k�GS���s�#{e�a��07pz����b�G8O1����������e���;�c'���jb�@Q����J�U�V����U%ׯ��>�&�Ї�4;� ��ph�ζӽ�::�5���"rřv��\%S/�����As���X�.��9�����x����s���u��[�'%�_k">r]Uz�z��m�O�(��BPG]}E���)&�C��-��<���=w�OVlrZ��J<g@x���
%@���fd;L*#ki���"����uZ.�mN�d���P`l+UU�S�]��c��v^u7�TnY�1������a�SQ�� �E��oo�<�X��Ɯ��=CN�(��{M����Ve!�%𨋭�������;����M�Z1ĵ�-�|;�G��z0�� ��0�G����ji�Hּ���ǽt�j���e'����覣	ƃ�gw�-m�ڕ�1[��=r�"�}��'�%��7���5�SK�m�!Ҁu޽ve�Z�{i��[c';���v#�ky]AWE'�y�p��j�V�
��ȉ���n���7�VY�$-c�_U�9B��<I�L����`�s�P&!DhԴQ%���*�׫�n�疴v[��
�t4J0�c`Ŵ/2Y�{0��]�+0��x��f�5�Szq�]�r9�G�p�
����z��RZ#�%2I�̱-[Υ�	}kkT��󨤭]�� �0ݤ����5����b��Y�z���qNg�	j^]��.`¬�%��a��%*�2�a�Qq�����,8��݉J���)����+�)4J�̛��E����ǂ�U:Q֗	�2mԦ9�N�9��:�� ��,ӻ��4b�[��_�sV��̕^�������%����Y���lt�R�Y���̬̀�f�t�[Pk.	�6v!���goJ��p�T��] :&Pf�����������T����e�G�}M�6��`���
�`v�3`��n6�U��^WNal-��t�-�:���t�R��]�d���n���{��{1���Nכu��9X�?��{ɼٯ�Ay48��J���	�
��lзx�n7*D,L��=IZ�;QYm�F�
U^֔�T��B.�sy]��H]'��f�؎�׃��[Mu#o��*��&�:2�,ȗp�k���z���En�C���e̮w{U�#S�N�'�(���ݽ�CY_F ͎:]Fml캈�PѢ̔�*3>S>�3sM�{l9�&t�(7H�&����`�O\��;5�:py�d��a���qlr��o�I<at*b���s7��(+����2�M�('����u�2�������ֆIZ%^yҗ`�͡�Wwj�t"t'�)�wy������H�MF1�nF$�E�!&jc;��M��
ɑ3(B3I4�Jd� ��"c�BJ��$!
L�2L�Bd�$�"ntH��
H�la�F!��JJ4f2��*!2�Ć�c,IR�	0e)IYΑQ�b�bK#
 u $b��2�fPH�s��L�D�BB���h�	�30�
L�FFL��%9�H;����w4C���DE�(	$�a�E$��0ғh�D̤F2��P�/=�_��ˤ�;�5�:�h�n糍���.���F]gٔ��V���R�<�M�T��Ùv�7؆�)�|�V�����>��[]MBq"M�����^a�y�Q<�g�����qv�=ߗR���΃|`�hM�%4�@��Q4�9�Mus��xd��s>Į�FgyQڿn*��K��~����K�]Nr{��v�j����nB��o\��P}�3RIȽZk��؋+��R����}����޸աp�.tV�'+5�&�AK:�����r���i�/�m1����W{��tDSɫ�U���9}:c1`R�>��M�J'��jo�]4��t���U�]��Z����4M����9n����Z��g���x�]&yͬ�oǂ&�(�r�r�����o8'��Җ�*,>P0rۓs�Z���	2[�{rs5��d��ޗK[��hI�8���������������+�S���̸ٗ��~崯�
�6U�SwJ����XI�m��&f)�V������˺��_7WS����`�.^!k�'4��:weӎ<����x�����9��p Y&a��;�%��D󾆭��rvV�ɟunt�wA��h3ƺ����)�
Z�D�'�����I��犓���u�����_UU}�Zb�iSBux���e���n�w�_l��̯�8n����t�"W_WCكz�zo*J���@wpWmD�>���V��b�g��
~ΐ�uc�N��������=Mb���e?m�����5���K��{�A����+��w�y��f�oq������2����α������u{��ńtm#��_{uԞ�wD����k�<,v�c��>�Q��Y���{*��ۦ�zn.�i��^�k}];v��{~n3Tt�nU7�pݩ����6����_ȉS{ˆgW��w=���溧m0�\���D;ݨN����I�Iȗ��Ed�Q��Rns\M��j�*V��Q��i�0 �6�����2��w���Z��*JI��;�1O�}es�W�4N|е�y��^�W�����o��5������uP��b�(�榌REr�^�]P-G���} �Ԭ��y�;݂�	Ǖ{ʣ�Jq�8�M��-��ybj��Qȳ/],ʼl�b�+ԣծ�J�C�zf�ј莲���;�Oaز�*��湇ҥ��e٢���+�il��yn�b�� ��Y�9h>���'M���c[[ioR��&G�����*P��Ψ��Db�c�Km��c����	w��n�C��N�DÁ�ai�.r{��v��zvg)�}1[����m�j�q���rʸ�3X���G��{춘��!7����n���g��<�-�/���b�kpk�s�VZ9E�X�l�V���2kƊ�V�S�|�7ch��	ܗ���Zv�^3���6��,/_�3+�Sw�5|`����=���vn���Qcg-���{���������';�(�͔�Fԡ;��)��o�S�8��)�서>�3n� O8T[�yy���:���:U�e���\u��ɍ=�q�窟i*6���{�#��5��.;6�� �26'3�թm���*���7��3��~�����=9�="}�2��y��dǔ�ǻ<9�A��z0��s�hݨ�ڣ&9A�v��}��,�����`�P;q��E-5-����̔{�"�yzWa���Y����A)�Yx��#�rƊ[neI��O���9Z[� wE�Ѻ��p��}(��|�������;�^���K��n�_�J=��G�}g�[zM���*��:��n�̅��u.w⩾�[��9���f��$.������vv����+��z殸o�>�Kѣ��RX��b^�iFW����{��?���OOt����J���p�������y===H��W�q):E\lM��og\�GJ��SY����-�*s0c'!]���+	wF�UWu⇻x���i���R;���T%��WB���n$�j/����_.�|G�ޥ�~=��U��y�e1Z�\7�Hʙ�ΗU��֋���Ϯ��w�kuT�����w�k��Ⳇ����BQGa��c{��.�И�sm:cz���(�O���o�o +a\5
b;�,ķE��O*tJܚ�:�9�lfok�Qa��m��el��U����*f*:C�U��_N�_0_�Gl>�̐
���<�&��Jtm�C����($����jj�g	i��~�1ZE�򫤠9�	rDI�Q���>���P\��b�Uw��;ҥ�����6ֺyo\{��x�k/���2G��M�nc��4��ZA�{L�㇝�lRs.I����'���o�քAŝ{�1�pk�'gr�����> |>���`��zi�ΝՓ����W�����B�-;N���ۍ�o%�췲1�;�Ne�1��_	Щރ[�6����L�����q��E7�uˊ��?އ�>�ۉ��^f:����w�[�6�ޕF���>}[��R������h�moݞ�d?-���iu/m>�%�/������xKXa�V�on�y�������7E󯧱��R���
�R��rԞN�U�v��e�*nv�Q��n#^�x��v:�u۫j�:kԺ;/�@��+��rЯ#Z�Y��|�v�j��C�׈J���������Q�N&wG8��Ҩ�<�,�z�ҝ�&��7�n�N�B4���jǏz��
N�P��6�9Y��q��O��:%��u!7�-s�ʫ�aˎQ�o�7������T��M�J'��jqwG���t��
s;�"�4�d/�]K�:fj�}�:w1�;�p�W�R<A̾�t�A�ط��^d�i�ܧݒ|��`s;Z�[w�@jgs7M�����9��ʏc2�e�k:��<�7��'8,G�L��,t�{w@��7��e�n�r{:����}߾��>��k-N&ȲOo�an�Gk����_q�U�0%Xz�I�<��.wS�
����[�څ^y>}�6�����t�*aW�T0j��$�ʋ���Z��^lm	J�]x�ne�J~��PV�aގN�t<�4����=_��е�P�sbsr�%�
�3Xt�Q�\ٯ����'������ș�+o�m����������,9��8���W�-�es��;UM�6��B����2�Å�9Q���F�g0�).��3���R�dz9mC�ɮ�]��x�ɝۭ̊J��ޥQx�5_m�3�o3��נ�Z��%+5�v-*��e�Q�sNOE-e�{�#_��ߩ����Q|{l񬞵�;�)泥O�*gVSS�Ԅ�g�K7�K9=g��*]�&��1�s�����L��*ݗ�8�Q�&5A��[r�o���
�l{� L�
���>���|9���������$���#�Ŗ�X��X�c�G��,�VWq�ve��S︚�hp6�>��Wc�#��˨l��N�T�b��7�Mm!Y�{i�w[����bA�Z��fV���~ER}8��dd�BDsC�S/�3������o&Ή~������!�7��� ��į�"�8��D/m.��LymSn&)rsi���.r�w.�G;v�,e�{}���f��j'Z�j��zR�-�f��AJI'���V���������PU�n&���LS�as�y�-}wYؚ�{©�r�.X�c��o��;:-0��8Xv.%(�Z��|֫�z�3S{��X��⻯=�����p%p0%A�z�w��"38�A��
9[�}��b�8��uTAO��asϣNe9Fa˦R㛒�Bf�2��������cC�"�]ve�}����;�֘��H\��U�h>�6��9h���Q�Vl�?JזfXW1�]D���t��9��[��LN����aՠ�g��Y�T^�]����{
lA�f�-������v^W���V<���r��P���'�.���L��wwqt������n�I����I��͘cWH=0;�ٳ��s���y�Ë��٣�:X��w�0�)l��,�s;�v�
�Gr�8KJ���Ed�3����Y�l�K��Km�[�6d"������G�}Z��ǜ���Nu���$ễ3n�Ș��J��ɗ��o�Vm�2�)h����c�� �K8ՠ�y�U:��J�Z����;�pָW�d��.-Ʈ3Z�e�D�b{/��1^�m�}Bg����Wz�>�^�1ս3�8Ejk�%�*�[gr�.s���(���2~�N�o�h�,�E��__I �	���,M��������oե�o�;S�r�m7�z��M�����]/A4�ƽ�\5�YFom�;��3��ک�=�|�#V����\=O��΂�����J
�����4�f��=����� w{�Y�;�V��+�q���=�>��\9���:���J[1��׻�bA�{퓷�;��9t��ݕmmC�Ms9���c��ow�Er�!Lh�_�mɩ)D�\����[��>鞭��k�^o5�Qo֑�'u�WW�pL�;i������iɻ2�B�ek�/��/F�<{��.�&6����"+:̎�v39��5º�6if�'u.�a�N�z'0��!�5��Ȭ"a;5r7�+�F�귚�Ѕ��Vg%�HNn�[<m�����烈��P�a��}�Z�E_�Q��lI�<����ize"�sg:�y�.��OE�;^AP�JקV�*t.)Opj0r͉�Vs�5W�*I���5��#]t��̧�9����W[p�B��b&)1�P��3U���C�>��y�S�����f��*ȎA�.��N[��P��f+d5��	뺣VE�Ã�gld>	Ԙ�^�V�,3�֬���Y��=)�p�'w"[�-v^�i��d������K�P��s�'̯�\�e.�Td�`�{��%�lBBq���~�iҍ���?��|}��c3^NTb�8���n2 �[<dֻĔ��3��s��7�nW��-�c�E�+��^��oЖ4��i���0��E|�ꋍz��ovo��r�Sݐeͱ]t.�PЍ1����������Fy�Z���>�.��U<c~BJ��s>��R9X�^�5ՠ���X�$n��q>�?Y�i�J�0	��ut�ُ9up|��4�V��������s�5����m\ �;�����f��9$�8��Գ�_4P�И�օ����㗊6�RѺ�m)|��ʑ�݅�GyCO�����&}�r� Y�������y�c�Ǻ᥏VV'��b�;�G͑ܯ+��_�a��v�;~�=�iKBu��}��n��6d��;s9R�����n��.����J�~ͬr�o�o�Rz�ti]�,�dM��ggJ4&c�Z�����އw�ʏ���J&+�����aV����n�F^���i���������8�*��B�*�7���\k�6��ksr��f��������p�d��4��+5"�%r�t���Yj�qV������e��;u��z:��U0�(�s[�=M&�9&�l$)LОp4>ۛV�\�/�cXs˺�l��tr�]6c-�X0u�-�]�������vD�T^�?Waŏ!Wt��̊ʎR.�jB�hLZ��7	�����O��f�\fbOaW�
�������.�>Z��a?-�Rq�R�V�"kra�^��Et�a�ܫ:��B�Y,Q��Jpɪ����ٷ��s	Y#�s�X{cJ��d�=�v8�Gw�n�'��X���1Y��mY�yu��a�i�N9�B���=qJ�C	�L��q�U�}#�훣i���X�JEV���x�`R�z���ʚRKcӻC6�����)ޡ�RfS��F�.���j�n�,<ܮC�Ib��*o�h,������l���6��c!�S����K;R�9�s�w��n9t������j��i��;fe
���I��g3�?��LzVp�/pN��g$٭5�`\Fњ%g<��u��t��h����%JkM�I�4���&V%nZXn��L3�%�Hf�]�-h}:���C�B�v���D��q��^��y���D�Z� �ֶo%)Vu4#j©³o{L0PCR�M2�77�!�"�����s�ڣ�P�V�,�ǯ��ŷ]RhNI�Ykǈ�³�`���>��Vj�
��v���Z�/X]q1�ҹlx�e��}W�v�} �T��ů��v�b�;����PZw><y޼��I�K��(�a�}��N��9���%�͟i�d3�ʚ��7��o=4K�5�H���ivdͨ徨�$���E}����禭�N2�̘����s��7�l2�wfv��ۦ���[խ8��	t��G�GZT;u����T�5��J��t���ݥ����u䘉�lt�E��`u��i�݇�t;i�0lS�#�'#�檕��4�������+��%vo,��(c��Tx�r̃e��x6����[��^SeT��p�O��>��[2��}pa�F��$�Nq�V�to�6�}o2�7�\8�0e�և
�T���Zr�ӧ�Xܹ��mMj�jېܮ�E�,���}�t�n��������*k�2��v��>��޵��� 2��#/zS�lZa�' ֻ�G��E5�Vն\�˰�lݳ؆;i����p�j1�]
��U�#��Ϛy1�|E[�m�Em�㵢u����7�W��S�N��Wu�ؓUq�z�ƻD��<�.�oU�)KJ�]Q���gMެ�t�:)��#��&�.��m�:��[h`xt�ވ���Y�j��dPM
�����{ϝ�2]����x-62��V��7 �¥��)wZ�O����s��Pu�����2��u�%GYI���u���!���i5�p�{ǡ�\wj��9Aْ\�)�R^fp�&�e��Q��uoMn>Օh�"p��A�CUp u8�:E��z]`��I*�K��=��t��W"�P���bS������J���Y��U,�	�1���j��/���z�F�����,�Wݫ���0fYx^T�a/gy�&m�tT��HV�[�
ܐ�sgtA.!�v7�f���
<��07yƵ�Ͷ	��ZYtN�%��l��M�,�<�hX-LδG
�#�LS-�ԣ!Ls�b_N�a�X8A����I�E]����/��&�8� ⵻�z��V5wJ�7��$�@L�ZI �L�d�$�F$�(�_�FF2)M�K&1 �D����i�Fr��a�n�;�"S%����Q�!%"B�L)2R	�u�$���,���e�&1���2�0�:R$	D@e0���(Q0�&�b6#3 d1&$ɂ�͆����5�DlX�F���H͊R4ј�5 I�1K"�9t$f124�S$ٓQlcD�q&(M�Ý3�����@������I��9p��dA���I�1�j&0����2T30H3 �����r��bH�{�J�5'���J2��l=�/XX��C%gf�^(��m�tV;��ol�Ә�|;��C]��U}}�֫j����}i�=l۠�&���ͯg�5����.Ҽ�
/n�V^��S����E\s����%EB�v�Np���޸A��x�@!y#2�����q��F�<���cT�Q;�_˙ڌkvnfW������yB���֠����<���Kg�c���O٪)K)nb�J��P��ε�I����G�ޙ}Tqv����v�1��>�ӽ��g�e;	��K{K�:����wkqƭ=V��js��֪�+�F����7-؁][���1�vɅ�*efj[�)��*��=/��bPT�ؚ���D�>D�mg(;�yo�Pz�M�����-�8y�	����)�6��Zf*eBT܃��f�7:��T�����mLΑWu��Ǻ�{��W�uTRe9ڭ=(hJ���ɠ�.��7����TS�οT�\�KNnm�m7<eD�����4�bVT�O�4���j��/�7|C�o(�N��`G�;��c�)E,OF�z��U��3Y�4F�(��c�W-�I�m�-���40���%�^�WS�i
�ǫZct�か�.��k;rt���c$VG�}�sz��'�qi��`������]�]�bs�e�U[��hLe+����W\XWN�x�N�t�'j�1<����o�bV���2¹�^��=K�v�6g��iv��|n>.㛡����C�iX?J���xu�TvE��R��v�gtr�0�󣔹�N�R���NOC�3Kr��,�{Ap��u��޷�i�1����5����Hu	8}q
f�+�r��pu"��;�7�I�ێ!�*�ŵ�A�O�]��J���0���n�uKe�W��ٓ��s7�\��c�3A��k��[�.���=����O��󐛅���@�D��U���.n��-]K�O�N�e���yY�MB�&M�}:���ɨ�<��샒�|�*���~���`�!p�b�ܴ{��T�@)����s��i;�zz����bWVye�:��W�g�x�k�B3���Z��Y��i}�-�y!�J:��O�����L�\S/F�y�,X;���K������_:|�n��v�Z�3���9eL�$���g2?������PΓ�c��,���a)�k����_-t��W��������[�hwO�ӭ_t��n��7���|R��n.Q�T�W$o'�<0�Q�;ڹ޻�r�ڋ-�Y|�����>}�M�5��7��GI� ��z����fm���p���ĵ�>UR��j�O$�#o͟>{'�`�*��b��0������uin�Bʓ�(������Uɤ]��P�٤���DL-�dúI�g�֯�~�s��4'�5}<O���PC�3��\m��i�.�����m�C)J=�9m��+_]��]�WO{!_60��8�)����Z���y
���R�Tt����*6�Enc�ǝ!}E������;���-����Ҳ����·uB.a��*�ӆܝc6�FXي�8����&;h�וI8}jf��3D酏8�,�@|�;�6f�e���f1`3�'�*�ΐک���F#��(������fo�L�u*�wt)�ort�'D���f��Q�^7�����/M�r��:�������GV�H�-V�1:W��l�^pv��┤4[�(2gje�{v�#C��F�iv�Y��/iv�pٸ$���n⍿}�Gd�������vN(w?��y����/��uy9X���q�ږ�J��}HR�g*`���:��b������]�~�W��I�@�[�)�LFJ3;Y���������������z�&�Q��>�u�d�=�����ޛQi�����6�[s��\�*1�ڵ�n��*����s�⼝�4�"gt'�1n��{n9TiYZ�z���w�QZ�)�]R���+N�9�(J{�UC�C�E�Z�E�Ue�ҕF��>O�h�[�g�97���w�%4g�ͽ���lOQ�o�1;�1O���*��Hsw/��o*�\�'72;1��څ6��hS��ZD�J&"���q7;��x���ϕQ�;����J�q�+�lm|�9��a}�b�B�64
�T�qŎ�f�������Mn���u�7��ѓ�Ke��05@*��*uѳ��{����ìP*�;���w!�JͭUϦ��]	�@��/:�CRMC0cY�U���M�ΚC��k��L=���)�loVwHi��֬�q�$�y�����J��x��f�M����q!˯j���+�G�����8پ�s;���ˈ	�v�+��8+��O�ݑ;���Հ��Ŵ����XaÝ)��:ҷ2�y��W:Ø崡Sfxۊ��:lC�[\�"��Y�)R1_t����݇5�qc�
�%�N�w#5IN[yT�� �5ꆃ�`����q���bI����B��Ӛ9�L-��2�g�Ys>��Ϥ�	�<��ϟU�ڡ�nb�������Y�滗Q�8�y�ρ�pvS�%F������n֍El�g����S�&{���ՠ=~��^NTbzkTqQ[�Z�v�a��Ý�6z��3`~Q>��Õ���ݝ��oǦ��^��X�V}8�or������B�8��\L������!���*�l��:}jy�8o<^���%V:��_M�j�Nj��Q�)K�^�|���zzՔ�%p����<�#ӽl�=F�؋�F��_'zt�]�b�F�̀7��l�Iq�&�J�����L�
�R��5˪�ݤ*�� C���wz�!�����H=��IG�d9\ٱ�C�ڙR��m_��ޣq����1��[�wevP��A���|pu_d�6U�菵�[��p�5�:����+�-=/�1�ARGbj'z8�޵ �6�*7����aMmW���:����,O�i��7˅��a�@J�z r��nt}=�7�Nc�}�F��w�Ǜ�v�!�������׳ޗ/�<h5Z�P��Y[��S�o��nܚ	E�.sx�r��O����W�2���U��-�!b�R�Hۘա1��5m�&��]��w��En�+[&tݝq'��=|�Ej�CG���)F*9��`���2��>��
����h���mĨ�i}sx�tj�j���e)f+�.�.�X?J��\.4���T\�>*4�a\��)�T��	�ۅ7�����f+��n����s�ۥѓ[:�=ln��_���^Om_n�;�I��E:
�y�=3W��w'�� ˘����h�^�nrN_���n<�*�}2���*����E��FDՙz���p�
'�R��ۘKp.���<'���-|�k��N�������/m�m�+�*�F�z���ձ�ouW3l���gP�<"v������#h�}gVU����e�1�Bphq�U��h�����7���}�%/��Qz�"��]|TvT9ח��������֨=-�G.�qТ�v��#Sx��٪
y��ٗæ9@̨.#��"�:ٻQo�FoLԍ�:���L����p���vZ�~�A�C�T5�s㋴��~�󗵿<�;Byu�6`E�Ҳ�����'���D}��m{9\0��h�1fW�.�&��<�� v8⺬�WV�F���{8z��.{,w�n�Ӎu �L�U�G�^gO^�]՘ޏa���h��Dt�[�����������%�[�&=��Wd��	L�YQ�)E�S�VR�t��:C���cE@<�,o>1u���R�S���p�� `J�5H�)Erj{Mk]'X~μ|�y�|�yk� ���]�)S��V�"�%rn`�밹�EP��Y�GRoJ��:�O�T^��o8+z1U�?RC�0�|0j��lv4M�!�v,��>I�㷯��ˑ��8R3��Y�����VmZΘ^5��j"���SP�d��M.H\��٧f`�Yʈu��t9($���^�gq�h5g��^[l��u��[9�;�'��j�cx�JWQ�嗳�+An�Η������M�p!*�@�̸��n����*c�7��fZ�9/z���T�*8�b�w���s��nMF5�@W?sc�Ұ�=�*㩻�%v*ɷ.�&P�o
IedF��l�v^XT�ڷ=�����`�N{jFL�s���w:-����'�݂���}y��/ŀ�}�U-Tfs�ְ�\�Y@ޝU���@!=�[6�ಪ?zۈ>�ۙ�e����/'1x��B�/��F���L�b&KU�gBc]��vi�>q:��a��ɠ�f7Jv�ΞkcF�=*'g�����?�jy����L���I��/�76�x����c�_P��|�>���vV><C���%�o7r0�?��Od�S��m�*�Jʍu1׼�G�`�>� ��7��N�of�\�X����q5+Z��l�wR��)�9\�'��tݬ�����[є�K���)�e���"��3E�H^It@�9��8��o\�����P��h�&�Y:�μ춳n�̰�Fc]X*0���J�;���s�oU�0�o�o�._>����Cx�d�۶X���7��u��QY����;�9�n�L����m|ZŽ����U�J����|�$�)����#yM�Ym�EPQ`俶R�p�y�6�����hUA�ZD�J-D��Rᙽ�d>-$�ը��j{zzӎm+���/~N��l���жnpm��}� a3ow��f��.J�t�e�T��C9�[�]R�nQz��gq�B����R5bv,,�n~/U�ٗ9��PV��wByqe0�e�yw�яV,O;(�8�_p�J�{q6�̰�e�W:Ø��[1�:a)64�&3`=\�n����9
��J�cHK8�{e�5�g=��t�9՘��:��y����j�,5������|��Fs"��>b"����,ń��)�9�`�����=�rN'�}�n�S�_m�L�ҖE����N�5��n��-��h3�K}����'8y٬�\��(T�D������T��Em ����<=�Z2�/�wgQ��MAuL�7��+�k}2J�L��$�&^	*�MI|�7������	9EE�>sO
�Ep�ط�v�Ev*�n���3���լ�XG.};���H�&��Nh�ǩ}�1#�q�ӎ�97R�;���7yMF/A��eꨋ�ʌoM}�m(��^��׊���u7���x藱��S���('WK샗���s���'	�8X���|/�R����L4�M'���O/����l�cõU9�%p�����5�;X�Õ�������v�-0!�Rat���4��ֳ��ϗX�T�y�C}��Bu�4a�Ū�-��i��z��0���
�D�X���H&0�h 2.ͫ/��ZS�p�9&6�g+�h[V�wV��q��O���q�� �)����]��_l�6�8���w^��7�t��v��-[���)85���Ě�)Er�6�}�܃���Z�s"�`u���x�!¢��l����,rW&�
}%ے����q�n�M��y��c͇@���2��lb�yfiJ1\�T0rg��~U�O��%U���<��§n�� j*�h�]�X����nme��;O=w�h�4#Y)�u��WشWs�`Ҍ{ݸ%�X�J0W�������)X=9V9�̜�.gU�<�ӽ�rMm�n�k�7�a5&�us�ӳ,��vi��DtX�j��8���pX�����]\�#yN������v)�+�0rw#˻ytb{��z3��B�b]0@r����Fb�2�QE�夎v��k.�X4�b��c��Q��[�}�Ul:�E��N��s]Y�}7U�֒���%u�1������n�����!S�|��'=���Ӊl$�v���x+�iT�Xk�˧:����f��7G�ڮ�eD^����a���Io4��Ɖ�$�u$ld�(ޚΐ%l�B�m�-�6�}9Yr�����Frb����űs�gU��y7�Xd����/y��4���n�������C%����_\r�Kf�*�:�ܒT����1i�1L�Y�͂��=�����ק:�%���`�]B��2�P�3xifS�$�8(l]6g7wÏy�14e�y��Sbd������&�u	�ns���5Id�V�x_R,����u�;O�w2��rXYh�A1�����k�w5N�[Y�i�7sk���u��/Go|�$� �:ח�⇶�}��~C�a͛H�"��M��@�V�J[k�I���P��8ӗ;�M.�Q�J�vJw�A��{�&AwM��Jʹ�͹N�y�¹��ю-;��	�宩�x ��Z�h�۝����8r�AX�I��{���SikCD�&�
�x��٩Ĵ��Gne��\|NB��G� ���:+T�vP\�.���]�{z�gS=n�Ө0>�	�1r�G���|�����c#MD`{����F�sf�Z���9�k.���z�(ekcq\ు�=��X�����we�r�Ƹ���o�oo��tu�&֑c��뾼�N�}��wn
)���Js.�:�J���}�fc��t���ȗ_X�Or��X���t�RM]jC�.�[!'0 �>��:�rSA�C�w�\�g.r�|H �l�{˗[��1�9��`9@[�Qֱ\C��':S�V�M�s璷��ǯ]�<�U�K-
5ݔ���1�m��W]R
x�7X�8mH�:��|C�Sc:󲒋9M���؟s<ϔ{a\��t�y��9�ӂ���F��9v�&�Ӿ�868�ۉ����x]�gvj��At�Jj�:�N�[n�npi���5.���9�"ult���W�:��]a�������p���u��v�[a>�5��BF*�z���u���[�;�t���n�A��l�$������X�>�P�Y��6�0���l��c�\
�r6%�ב��Wb;��-f�I[���Q��ҳ {���k�*��ۇ�ot\�N���o/�dw����a����A���:k+\.���']YA����g}�ŝ���aef7Gx���G�)�������������~$S&f RLP�Wa3FI0�h�Q0P���e(e��E%ERf33&��̝�`�ܻFI�3�FBbD@B$I���!�qIbbf�H��d������$�I,ĄcI��Ȋ!+����D]�b$�QA"wW ��	�H"676�JB�&Q&�vb$$d��,�%���	� �"P�&fL�(�.��$`ɀ�IC!F��\��s2f��s��AD�	��큈�j!0��$ ��l�baQ2�H�hD$��R���tt�d	B�3I�ha�	��	�꺏�����ڷ�A@Y����/�������v
�m�9��8ow9{|
 ��N(:6{�����^��1�\=2�Ί���:co�֍}K�Sd>�n�(�LD�:-\	w�;sJ���p��v��v.�yݻY��:W8{jnC7�V�TGH}�npsՑיb8ڴ��Q��7f�v��Zg9�לB��.��p����a:E�QM�JT�� 4C��՘|�K�Ey�����ޙ�1��ڮ~p쩵nj�15��[q��׏�8j���u�C�yy���r�=5��1���ӓ����X9�w�T���A<�����Փ�ت��ڿT+���SO�m.����c��Q7���p��Ù10�tJ���Mu��Ciy�<�g��*�qu^�b�w�%u���j��̗��J��Tu.n{������h��ܙ�\�-︧��6�q�Y�a��ҷQn��kr)�*���ܡn=���&1=���YVjB�U>�p��;h��GO{1	�^��Uo�����{}K2��{0c4[���d�tx $�tW7f�EG�|3ed�ɨE�mh�>�n�����!�`ԯX��*C;��<;F�u�y��x��e�����ɦ�9Y�H.�C3���Ψ�:�q8ź��c�����P�DR�'+����hoR�fN�<��W���b��^��-�ȥ]��9����y�%g��>N�gE�n�W?�]m'�y��u�у�>��jJQ\�����|�1����R�Jӈ�I^��W�2]�W�2��*9mɹ��㎚�Efۭ^���}�r�l��7�GKZ������uu�<U|}C[�^*���z��}�*��<�P��6�u����:�<�V�LR�c�Ҿq\�*��	�S4'���+nw�ov�+��a�ܺ�8m�q�Un�[�^Wa��B;ս��)h>����#=��)��Ƭ��
{Y���H�s�3#Z�f-E��\�Ȗ��7��M;��W��F,c�9sj�-k�����K6���<WE�4��2�|˿���n����ʻ�9j��_���ٲ�E�}�8v�d�}Q�8�s:�ܨO�C�7*��垳@>�{�T��Sƪ�+'�YS�'knO���s�e6�Ԥ0��S�Ad�f�0��&�clӼc����e֍`&�-���jL�y��c�N�鬮��R҆A��u�;L?�'�˾��9���[���ER�i��]gh�'[������v�)��ޭ�<�ui3��Mt�c�U�J��x�����o2j3E���Ub���U���JND����ss��mTF(�Z^j���m�|�uG;����bz�s�;B3̎^���~�Xf����}S��9k��������ƵuϦ�K1q]t�ԉ���ݚ�iv��l!�cb+Z��<�,�w�+f�F5���L��[��A*��}�M�AW�z�.�
�-���ދ�|��5�oe����O�MFi�Zy���{��&���spx-�����t,�:�|2Y�y#gc�*7wz^>�x�9��5�n�F8�N��㌫ƻ�`t�ZdW�l>�C��bo�'Av1��l�{�J}��OPy�1�N���:�&1�ꬽ-����C�XՏ�7%k����^q����?_��BE�����hg��h��p�Gn�����9��6%n\������ڶ�g�h� �vyk�-,4la�y��nD��wb�Sn��_N��v���L@�HJ�3&� $KH��q��z���]{|(n,�u~4��*���x�2�y���l�!�J.@y�`�c��L͙��?<���m.�έSZ�( ���ZDs�\�%O! �=�|�0K>��)��o:�Zr->�
��C��
�d[�o*�I��&����z�f�3�y��'���|K]��Vj�;���*���z�oOHS�!����9�qdLk�zj���9\j��4N�?�b���mF�\mSw�TV<��G<7�0�^�w5;�8s9���o������;nT`N�'�8��v�k8�*�S�z-ZY7�g�zf^�?�� ���(s��?�?�u/k�,�5}�ب�Q�p�T���L	�_>��v�R� ١�����B�����;�����sO��$��:|����i;[kӮu��\�ƗQ��Ez:r���������lwN�\�KU[���5��t�w�����=Pz�4��7�w�ae+I��4FC]qZ��|�R���p�m7�W�cU��XF�sDF��cQ^Si��J��,��A>�l��qU��fBd�Ez�4"�ס~��pvv�Z�4��Im���6���[�S� h�F���7�#N�uM�#��}����0�]�LpJv�|��k�WP��N<���l�8����a�4��[��{������MEķ���}����t����8���&�m��-Pf�K��w����˜�.��U>�v/��<���T.����7,��s��o�5_DJ�9q��_sJ���.��T��Ӄ����p��٨G�/�x�g»���g��ӣ?[O=C�Op:��3� e��`���6x��n���S/�{<rn`7e��m�<���$�!�l�Fkݸ��zB�r�Ӈ����i�034��ӕ˹��X-�&/S3[��^m_i�x�ד!v��'�Lۓ2�~�uQ�<O)EAP�@uE.�Y���%�W���c)w�g�����}ks�M\u<ȧ�u�B)��kȀ�n����s!����U.���I�����E،����<�'_ϙ�{fS�'��t=QpcW�>Wμ:�� ��+���f�t[���S�OM�]
dM�)2�웎�ٺ���)%O���Z+a�s% �^Cմ�z]��]��Lcjs1l�bvU�v,f�]���d�P��8 ��81bv��(q4�UTNr�$Jվ��"���0�V���>�O-^�5"��n@�7WZ}:���8I�(�y������{���īȝڬ���/0���vOr�s�y�^�S�7���ԝWx�_��G���h�b�L5����b�>�q��X�#���m�Y|�J�M�|�C���`��[䊽�삄S�
���,q��76���1:�H��t�{1	�^���+Pd%�a�
z9�a�q�x�n�J��7R�|�,����F>Z���uzi�k�Y$&n)���w�hv��Rt���\���KP�V������hU�Ś�s��q�2b�T���XCzr1�پw�OW�Z�=Bl�P��q��"�U|V�n�'���JQ�a���rWC��O{Ө\o�V���$o��&�uk�;<u���������������1ҫ��*�<��G��[q6ҷ&�ݿ�����-�p��)�b]Eȁ�.,���*d����A���K��G�����*5WE��x����L�
��lrs5DT����.z��=C��� /:�_�+{�=C$wR*���3��ǫ��-����j�	�S��N}�y�ҲٕK~"n�����Is�o�T��������Uc}�b�z�i��v�+�c������'�u�#��
6�^�S����=��5�)¨����7C}�I�W�.V$��]�܇���KʧP܆���Nq��eT{Ж�A���L��1�e)�r��rQu�����s@㋍��qG|y�6nv
�|eAp�D��`����ObS|���I�^NT�y�mp��O�ݿ�zD���my��&���3{݌nk��J+Ǣ�������;��J�����ysk�j�B�nu����ms��#,,�s�!�9g�f��G�;~c��l�s:,k�H��)�)[�{��͇�;���C�&����<��/�89��<�{��(�4���5�M�W{�B���ur߱�9N��{��fF��Ɖ�b��ڭW�Wf(y�	�F���V�-
��]w��7���ȱ#�\�������rp�N�s�ʛt2�M��:�|"��%��ֻ��(lމ[�8o	R��`+Av���氞�G�w�'�^��9Mύ�g_>�̋�E�]��7$qia=y�^uԝdV�ЪZ��.��R!�9�4�f��w0�z\�:��;J}�{ls��&���)�]4��i(����׺�{�6ʫ��{��ӻҝ�(�*'q�rjJUP�q���PO�������;`�̻K�'UE{w[�r�{}���p�:`�tZ��.̿�s۪��o��oTڼuH�G:7�m�+P��Oa���E���]�uK]�uޒ�נ
�V���z�S��+�1�n�w�vٲ�:����L�GH��}=��ʞ�A^���4�j�;�E���m�W/h����I�h�4*9���}�3K��92Mҭ�������s�󞐦3�4��s��,��@�Ӌ0��47�D������2�o���[�A�[q�u*-1�	�=�;�2�@1��WV�u�l뺽�_^NTbzk�P~�Q��ă؜��ʆ���Y�̒=�AmNA�=Eh�gN)�}5p�O9�+[[��ޢ���邯���ڛX|[t��x�rSe��B��!Ս"���Wc|\2��#�cWţ����s�����Лz�R����Z���Q�+�/���Ҩ�䴛�<0c�ݲ��;�<#��~��g���=��g���qv����l�\&�K��9�3O
ʆ�w{=�wx�4����w��k�guf)t�nP"n�^�:W:�q[V_;�ҕin�!��q����kr���%N�p<c[��$��
܉����m
�J��:��wܲt�{��P��5��Ш�)hLqt;"�:�M� �6[*����b���혦�q]׊����=j�wfGRRLż�n�GV0%A�{rjJQ?W.sx�c/J��{�6��&z��:��1%cF֬�ŗT���E��0%J�'��ý	���ݬ�����XdI�(E�ݨ/[��G\&1T<�I�a��`շ6��H69bw.ґs�%V��e�s�]A��7����	E���	d�_?��8:5"�A��A��MF7�p�HS��\|�����C7�ȼ�s���4:nU>�I�ٞ�u�^X�alø>Kե�^#ה�UJI0�]`���
�,ܮ�OR�NM$��\\O'8 #�),���a��4,�[G�p�(�V(�Mx��c��q����Y�f,.�� �n���8��7o�7j	w}c���^Q/�V�+���5}�����3�R�zg9�ד�mZm�$�N�����Å�������\���g��3c�v7v��ϴ���}�ƣ�w^˳]�0��34=�W�.�>�G����7�V�g��P��H�0;���y���x�a��L�N��~ۉ8;(�^�/�TT��湐2;Ӭ����ǟ�I�&���\���kJC��G	O}#}W����ǸJ+H�>��6�;��}~�ג��n�M��/a����u@g5�Yx����������</&u�d}R=���
����?O��|�)^�!8�4|�<GO(��ݟGT�쪅��]1dγ��&��1��?_��{�y��W�z���b�2����wL��ë}��³��'�_��4����Nrj0	���ÿ��f�e��s
�J�x�:��
�<��Q��7;�c�/۪��=%���"�2�{7���>Nn0�mN{ow�5���o$^V���|3ў�飑����}���ߩ�|VT������@>Ϫ�]}.���f�����������^ �@�5���g#}�"$�T�����"|S��Sa<>M�[6J���8k.����X�#J�V-�����FR2�>/�r�����ShWu��7R}�͌��p�CO"��[���2�\n�q���j>�_Y˶7lL�DL�(�>�[m*�xޤ�j��r��0��p��1�0�%��v] �=��\���X�:�k��Nm}�U�=L̔��:���d�5R��^�Ů�*U9�\���f��E��nc�g>�Wu�
	�e7�`����:�7B�Cu��!�����֯*�
f��>����2<Κq�3����g��b��3�bˢ�A��b�粢	$D�4E��M�����{�r�Rﴘ7�9�;���o7M�fLs�:f�w�x��:e8E�E�Wl4��	��)ub�×����miRԭf��v���s���>����_pvn�+e<�V5KQ�.��R?&3c\��!��/d�9t��]�Z�!�	Fj	#'oN3�.��j2������dU����G�غݐ��ɖ��ֺ5����i��B����vV��p��͝��ot��rit���B�R���%R�tlk�QR���ݡ0v���X��tT��6�ě���%�i���(84م��J9C+�3���p�9t�+z��.2�6Y$���6�|���v�t7�`�fd��ē������s��o,�C��:��� c�e�,a睍p8j:���Wf��Ʋn��!��J�v9H:���b�˫� R���g(�J|H'E�2g\��r*��Rٜ0�ҝq���ٔƃ�sv���� �(9�-��<��a7oT�;��{���u|�Hvn�٩n8o=����e*��^u�Ht0��&�+;5%�;�P�X�B�t�qWv{�;̃SBE�nk�ɨ���wH�n�v�[ �>�!�m���s��V0U%Rا0��H�51��o[T�ї���U8�ֽ���1wF�c�)�hi���|5ZT�n��ښ
H�w�WxJFwvt��a:��2)N�!��^��O]�:�sD�1n^I{Si�{�I��"-@�ֽU{�yXa	{�H�Txb�������zw��*�݂�RM������<���vX�2�֍Β���6[�����%���Tm�/$�SCU��)�"�p���oU�]��|���{��ܰN��؟w�A�H�ޚN��FݪǪ�38��)�j��T��	ǧ�wqŹ�x�o>)�wF��"���i�8� �wԝ��8����ΙF��i��i,���LS�! ��m����v��"(s�y�}���j� (�5��ɱ�S0,��e[P�g���C�jĚޕ}�De#X7X���s3�����1g���c#@��gc�!j8^�֯Dj�;:�#>�����*��Bu����Խ��F�4#�ue��x��䮮�S_Fb�]Ib�mC�"�Y�t��(��7cx7.�P���a�����X��mM�DA��Z�r��v���CL�,��Y|�uʳﮯ�b�ʉ0�0����1L�o�5�j@�b�A!4��&�Ay�DO;�03 B1��L� �n�3"x�C7H�˘،A�)L�RL�2m2)�##1L$�d�2d(�F<��7��/;nF4��2��B�)EA�F��DeݷIDQA��;�-	��ݍ��RF�d���4gu⼁��ٷ��2�*D�%d�!� ot��I#2�"��0lP��&��Q9ѻ���;���۔�S#��X���u2��)��D����.�H���2h�GwT�@)ݸJd�O��H"$�I�)��m
.oY�J�C��o��5.쩺��8˥�Y,>�x��$��q�S+�W;��3��kU�K	���5�:Pt�_?Kfo�����F��e���ꝿI`@l��������7y��e��:5g�o�w�g0���S9��௧�.wǇ�O>�I�3ِE[�n��L%��atk�E���Տ_D�ݕ@A�u4p���D	cԺ�x\���9>?S���84��^�1�])��Aɱp<ꥹ�$���	��}[F���/	�O���_�Ѫ3���ްoњ��8����M�9;�)S�Ъ���5V��r�w��;����o��s>�>$��E��~�N(�~��\�����$���>�+���]a��\r*��77kC���xS)�s��Zke[��(��3>�(z�wp�UQs�<m��G����_��_���ǲ*�����a��gi�{�;��z�>Hߜ�Zn5O���`O�^���Z�5^�7�uc�#�{�/�	�+�����{�w�Z��xi[.�s�mo/�͚�k�7�L	[V��^���Q���#�q9Ц�d�4ݜ��'ӹ ����yi�qϥ�ë*��j2���z��ƹ]�H����*�g��_j�_�3��j��ۿ�N/�8,G@�L���o��6�/y���L���P��V9|Ȧ��U�K���7֫�oj�1GD'w�����5�W�i=�`�ϳ8=�v�$�bR8��t�v��6�ǋ��/3��6�`Ƴ�}ٶ�ΰR�]�_VK�[9�g����ѥL�3q]ü��N@L��6���ԉ�'�M����D��X�S�_�.�Y���lg�QEk�%��L�ިk�Nb}$n�q��7�����}�2<�z�g�~�⑯iR�\m�s�ʿ��E3r� �*��ט/��FO���+��>��}ΰ;�����hz����J��=
�Y�υ;*�({3��O���5���о�`S�UH�|��2�>�aU��x/y�;�+�f�����G�z���g�gbǳѕ����n&%i�?@R{�ge@�L�C"W������P��t�;��Hߧ�|�ɳ�_T����;Ά�V����W�=(�8�|����NE_W��Ĵws�0�iwT9�3
�ȃ�ɴ�R��|�� �S{Հ�ʐ��9"�^����W��eL���_��϶b�Y���ҽ:c݇�߅G_�j�M�+��n=^��޺ �{�I�H���_���#��*�(z����Ή�+&Q��Ξ����B��ʽ70ߤ{�C���r������
��ؽ��/����C��a*q��ȵ�YP?�d�DT\9���0����(V�F���e^�B���B���P�B_�!��ߓ��4��b4V�HѫGVy��+�'xmTa�u�[�YG��rwT�=��z�K��c��k�ki�#$����{#!�P�,}�=�#1��N�ǵ,Ay�r�'ʏ�=1��������<�� OW���UK!��N��={՚�>�\/C$�a��:l�s�>�iȍΨw�mV���zo��`	�N��̐FOW@���Q��Cr"O���i�����n��BpW���"��њn_Q���2|�o�,����,ܗ�w|�ґ�?%@O޿V38�Gq�y뉿��o��{R;��N��������j����f�������ǗTǣ�G�7���@U/�����Oq���Gj�gE��N�h)�y��=��U��{��UY/@�ޕ������-�d7qƽ�=�^G�=��o�v�7>~�Y���eJ��<�v_��r�������9V�� T[�����x�����:ϴ�����# @{���R�:M�17�E�l��7�ϲp�ۉ���7@U�^3y0�����E�G��to������Q�|wЕ�����d)�,��[�},t�"�[�r��V}�x}��p^͙���<���1��Łν2C(��AŸ֎��u�9��S��k#AH,.��E\��l�O��w��ƥ4��Ȇ�&Vt��]|�^MK�Ӿa�C�XкV�r���:���y�E�T��g�B��]{�j�k�_q~���q��Y^=���P~�W���Ce���*das�o.+�U��@{�W��+��4^�g��Q��__�r�8�r��w�ˑV꜐/��>f�:%΢���g��ڋ�^o�9��O�Ӻta�Zv��z�z�]u��s��L�J�p"=wV�$��&6w+ۯ�C�}�ۨ[�bZ��������[W%��,�����T���4+v�rb�k'ҽ��L;�$��%��5Q�荬��3��kK�꾯�����
B��Y���P�otI��W0){����	�k~�W����W��M�����K�#���ġ�_��a�:�/*^�����al�ù$��l���?Uh�3G~�D�r�}@-7��ܜ�NK�S�w,��T�^��RM�Q��>��%׮=i�o�תx߻*%��Q�|Oi��D��� ^��Y�ލ��-�2�ۦ��
�{�������s���{}01������*7}�<c���q�ݓ�|_�u�3�J�i��c+&����=��]�H��GS J���5����u�e�چ8����zd��|��zy�MͮO/������Q����m�qm�7	��j�t�dC*��,�e��r�(_9)����V�u�����V����oWm.G���@I�C�d�Y�R20y�*&襛�U� !�]�ss�n���GC���3��8�-�<�����ЬY�F=妽���V}U�Q�鋌��n2g�<��u�?_��;�*�~��WM�\�zTV27ܲ�p�!(+��F�U8�1`g�޸w�S8K�G\�#3��=���nѮp�A>X}�>�Kb�~ڦ9NQg���w�`>���1M�
��s6+�P���>������Tc�U\���U�W�#���Zm����O��"�M2� �g�@72E �!y���K�K�Olr��|���k#g�TE�hv���ޅ\�o�i��[�y��,d٬F9�N��k"vC��oz*�a-�g~>���ς����^,o�i9��e���+���&������*�̒���R4�p�c�2\��3�KGw"��=����[!���{@w�'��sz�Oq� ���[�n��o�>��f��}9G�K��τ�¼�vS�Q�r±�&3w���T Z������� ;�&)��#����vܐ���l��/O���Z~���٢j�\�]ς�1�gʄ�R��l�����9��zH|�ļ�u����fd�{��Tj�򘷷��-���yV綤tA�'?�Ȕ�Ѹ4T@�^�x��[��/z[Y���y��^5��b�)����k �*�H���
ޒ�E_s�e�qڡd������%$�yKe;�����Vh�}�R��[�x�jJ�ː;��͜�([�]Ai6�ܕ�5m.Q��0ǺL�gÌ�}x*Ww�5UL_Ͻ<m�]����U����l�L��k�{{"�r<�N������Ѿ��d�7��5L	��������Ң=�Zj��np�}��-��zc�ٲ��q{b��`~�d���S��1�?����`J�@������qn'/վ�>������
�H�j�Z/��>6��;�VET<9;0�=]gYuH���@Wxn�G��K���C�'��ך���;�ƐǓ,�z�F�2��w�&w�q��=�&=~������.����:��"���Gq�6�}�Y���e�
ʫo�p�}H׆swޗ�)�1V<��=����!��߰�?K�H��}ĻU���+7�E3q-���UB�B먺�����?�����=/H�����ɟ��9�Gh���ҡ�Q�o=Q��Y�ڦ8+>W|bfZ��|�G��� �"�E�Dϙ�ԯY��
�s���#�t��{�dk�7j�r=ތ�Ś�L��(n���������҆#��QŴ=��4�V/�_{6���븱K�$O�Uz
/s؝����]?�C/k��ܽ�֓ȋG��S��Ϻ�M�٫s�s�U�S/xY���[�w*�5�imfhI3�F�E-�gQ:Tuzm�e��\T��c/Zۤ-F�{ԍ��=z�l�gN���z]�J��A�y�P�O/,־�V�2�e�u��I4������W��Ϡl�9HOfA����>%���+1�;�-ݱ�8}!�
�E�׭��<
~� /G�nE[�rE��/�W�g�YDLS�ӾH,?@5=�k��Ma,�/|�������W���E��I
d���]xi\��מI�*�����-0I^!z#Өȭ��{>��V.�.�vLd7�M�������+�d�R�l9��I���q~n�v_��ʵ�Qy倧X�?:���x�z���	�顾y��K�FLϮ����}�N*
�|�	���R���ٵ�a�f׸����f��z�^�]� ���+����5���Q�~VV)��\q�;�J&���{,{ɬu��ⱋ��@k�;�_D��/vΐ�����[�<��Ҿ�n܋~�Z.���H�e�Ek5�埸皩�x����}&��]�l� ^O3��Xno�m�p��W�ϗ��y$v��_�Lcе��ٌ݀��<�}���nc|B���#�}뀮Zs�*=��_��oG{�Q��;%����cyJ���$R��ڋ���d�Gb�Q�:��r�9OM_0��i����I^����\��1���c����w���m��䮭3A�oz���[N���s绵7Jc��KDX����'ž�ݨʳ�̈́���,�et���W�C1$$�r����X���/�����/��S~�ѾN��mϼj%�C�
歿+������+���l��?1w�&�\��\�O"_�3y2��u<,\GK����O��Z�׶D���,���ˎQ�}�}Yz<1�\v|�+�m̰d�d	���
�R�g.=~�C�5l�]�@9�L_�پ�`���������|8_���x\J��ʀ�JޙV}-�
�MO���ýi��-7|��яA��j�\O�i��#���'E{-�q�x�Hl�Y�$\&,������D�y��򳞀tv���Q}�����>>��Q��G���h�s.H
�k��^sS>qQ�r}�ѻ�z#�oz�I��H��9���ޮ�u��2�{�'��v��r��raqT��g/ߖ�b�~h��t%x���P�͓�m�s�݂X��RX��l�P�����5�%��xM-����V}`_�������蚻��7�Fz�MF�����U	b�B�x������wgt��U2 >�}ڨ��T3� ��*�T�G�෪k����<������%R�^�����h��V���,I;{fS&%�Q�@��ԉ�{(Z�y�Q�� �&WZ�^9ػG�˚S����ٗ�B���(+�!=�n��]��Հ�oTt�wLֹ�d��eI�\��!V������!��N�ڰ�Bө#����6S#=%�_��~�b߲���񯟪��D3��_�蒎\:��������uhp����٢◔H8J�#�f��.�؜����y�3��n��߮.3�����j^g�ui��9S�����x��X�7��F�o�j�
����׻��sojt���r뛺��՞-���w�Hed֟����r���G���5[W��ep�g8��������oQn��2F���ږcў�M��T*��qT���:��ς}$1��^ç��B�'9�%�����Ge!��c7ݴ��tiͺ�ɘ�2����n2e�⢽�� ��W�|�`.�Q"�OORG�+��}~�
�_�)�,���-LӑF������&��'7���kwxy�O��#R�������r<{�{��Y��²���d����j��<�k��q7ո<�H�p�NVQs��k#e�Q�|C~�x�GNu�;�#���<��'��H��<���z�E�T=z}��ݟUHʙl�9�����U���=⇽��K�F%|8��{Y�7ܡ��z)_=�肌M��Sۉ�}��Yqë��A8�e�= C�ך��ځ��ޥ-���
�Ñ񻤅n_rE7}���Z�HA����U�x�ڊ��6>�����C��Ί���hq�I]o�K�'m�˘�Zp�����u�r��*�3S�Ts�h~�>����F���EP~�}^G"	h��cܧ��Z��,��$|�	��Gd��[�
�3Z�+�'�u�p.Qno��!{�"�LS��8��T��un�k'��4��2�#�=ί��@{��� ޺�z�
����Ua���!���Ml{�C��^�_�}��ÌRn�������C�u�n~�
-L�������K�S���VW���
ځ��:y 5�^�W��φ�����Ww��T}1o�<n��zM�~�����݊l�/g�)�L���Uz��9��N��{��3Q�����G�D%\�GO����V:�ґ����H��^�}.���z>~d׸�h��>�nmg.3f�� g������/m�U��77��E�z�w�N��Gߣݷ�E��Ѯ�y����]*�k�,y^R���O����G��Ys��=xw5�����{o޽eW?[�:CF�l���,���*r�Q�����vr���Y���V�яg��,mǽV)d�>�ǲ��y��!�$JX+"*�"�Sn�0=<� �L�N�\�y����N
.L�N�۬��<��v�딥���>�.9��@�
�[ڷ�3n���vK��b���h�*� ���ۗ��L���㫞L���퓤c��%�i��'���t�����s4�愡��g?[��N';%�4SfJ�U��F"n%�u2�;�)B^(zu3�p�;��,['K<�ep�wK��"�/+zr:���C�.ќ ��nEmH4�6lsQs�;+-�Fj�Y��;����FѬ]��l56�'���:ޤ��)6��Z�Z�hP��m���vV+�9IJ�'w5]�����1������α��k���aܨ'=j�k�Cd��B��5�G�@
�	���$���>t˔���n#3o��4�� �ےV4y;u+/6�(т�@Fy��w�%A����y&�V�՜�]/]�ę�����0���`��+F�l<��	ֹ�u�u�<�N�Z��8Ҿ���P�;���W1pt"�
9���U��>��B���1@��B��w�F�C.�ebu���>V(�:��r�fda��t�|w�k�1��+`}{����J�(+���7�^��駢q��d��|)靸;���vr�o'.��}[�ԏ\|��P?������w�H@�C1֊<^n�6̝������jg2�d�����VvG�����s����*x�ZY��ڭ�Sa@�,vq�uVl!�2W�)k�H��٨��Ώ]u�>�=��*�B��8��]�.����������G+�;�Mn����ԕe���%C}�q��P�\uxN���_�`�7z��bWׁ�`��8��bw�C�e�Gݗ�����6k��bl[m@o� u���\��`wK���T4c�6�u�	�A��WKBAK�pNҪ�X}v���j$�K�Rt��C�̐���[��ZWWn>�36�+�3��t)*FO���0�l��rt ���Rݎ�zr����5�h%�����,JV���EGr:ч8:�i}���\�i}ʅ��i�*m��@0g�%݊;%'X��ɳ0�e���f�8�Mŵ���f�*�^\U�z�ξ��=�]v(��H=�R�T�*PTv�Ңh������/�VX��U��D9D��'�-,8--�,�&�둤s:�5��1��+Oz���(z��u�Jf-KP�3J�w��c=��w��0�I*��L'�<�/s�.k��ȯ>�#,Q1��������TU����Лi;�Q�u�U���Â�w;j�eΠ'�ΥhV�I%WRQ��z�z͘ę�o`�ޡ�Z�~)�=H-�}ͪ���Y§����4�ہC����7�Ļ�R=m�ʁ��� ��[�,�IV�{]jzze�F��nG�6���ot)My���Vi�g��S4i�qy���s5:ʶmj뤘�c`­����ݡ�C+��&��Iy�(5&�
S5�%O:����QRT��Fe�H�ƂM�&�	o;���nnQL�,jM�F5���B4�ė�җv����e$���(�*�$iO9��(�QcJ2��d����FM���h��MQA��,A��J$s�&* �<q��1�aΛ
j2%x�ђ�ǝt`B����̩'wDm�;�),y�c@��4�flj���EE!�E��Cxڹ�����u�/!� 4S&k�A"�!�e���n�\�Dh�O���A4i$D���F���o�{�����T��
��5u�:�f�UآR�f=��6u+�ڵ��;��+��W3\vN�A\p��A���K�$�zr�� w���)�鋌��s�q��^��?K�H�<�O{���ʽ�Y�L^^��l��e_�7���ު�'�"+딋Kg�9�q��������7��Yw��u�b7�j4�hNI^�0��R�g΀}�R.�[ U�^.�XIg���?:b��=��<6�R̈́;�E��(����#8��z�A�PȊ�
��ω|}써j縰z;nt�U鮍ݽ���H�(�����L���4{)�������>s��E�K���Z;�x+G֦���ګ8�>^u��c�ӓ�������ݹ��$T*�ϋ��;=$x׸���]u��k̜�-�f����;�	xk���B}v�As�>���^���$Z�!��7����f��9����c�(�e鑞���J�C��U鹋z�c�H�cd�(�W�%<iz-z��Ty��V\-�ݽ�|:Mk�vX�%��U\[~�=>z�Ǣ�>�e���|#6�����z��G�}�UW\{�s>ͯq�z#i�:}>�f���]1Goi�˥��s��`ݫ:qc��|-�M�xܫ=�zlN�֫�N,�m���mqWC@
;��_��Z� ���w���l��SU�M#��m�:��C>o�Kh5�f��z]K4/CgH�WҶK��h�"C��l:�ȃ�b�������NZ���$�Yݧ'���Wc��2loz$�˟PGO���{s���i��v}�9���x���Ц'�z�����q�N".W��4�6r���k�ߞ�g�L��h�f���Q�`1��ֿG�6}ǀ�M�p6�� ������w�y뉸�m��g���mh*׈S=}�Ͷ�:�g�4�\dι��!9�2=����[M9�����+����COڣ�o���Gdb�� �wv�J2G��gʶ�g�X�E�'��/���׼pg����ǲ���������w"�?>�m頋� ���8~�\�.fh��@���p��S���S�húTp�)8���a�*dy��n�8�CÔ�w>~���̰g�Q�'�n���+�o&�{;�#d?]��/���
WpX��@`����2!N�e��-͟K�2�������x����\��X���jr��	���Q�~���}C�3�����_�FG�\�X�!�ptKg�Nξ5�ó�W�;ҫ8�|Ni����_W�W�ӜJ8�'K��H�2䁍n�tu^�״2m�kGW����b�#K��%��wR�5�Ν.��
�=m=�G��y�0_b�9F��]v^�ڜb���p�M�3��꼠��*����Rv�|�X��Ϟo-�a׋V.ޤt��VA��e��V;�X��{��Ȋ��q��t��Ly����	�g �Xq|�]ޤ=�.�����L����/wX�_���<���Q�A��D�=�����ݟ*�bb���q�|;���R�%�^�f}�cQo�G�*�[딅įS�S�;�ˀ+�<�Y����,�k�|�1^+��ǘ����h㘶�
����~��E=�ݪ�r<�@n�?�O���YR�\:��]���7���k�Q��WR. �J6g����gʡ��G����Rȷ��<n��zI��蒎\O������7g�p*%X�fw�O0��{��ޔ=�<
}Q�	�o��>ҽ쨚�~�'��ި�=Q�=aL�뉕�/B��^�y5��d�Zn5��M�`m'p%]{=02�%9�ۉ�u�5s0Fc�k�+��4��я}����#��c0Ζ7��� k����`	�m_�j����*������^��;ܯ3ö<��1��[7ꗤ���i�WLa:�FL�'�R�>9ީ��J��Zú�q�G��:�]�2��#]sp�p79Q�LWz��a��yc=�5�Y&u�x��8�B��{0
�ue\rﳋ���KmeAҢ41�������,i-LJ��\��U� `���=�8�����q�4��{��S�_W{֗tc���M�}�%Tz�ĸ4N�$��N5ˑX1�Αv]쵇��{�<���⺽^	�+b�Pg������̎���뒶���d�+�A��3���0����{*�t��G��Q�|o՞�������+ܷ-y�.�=�9k�:�.64wx�Vx
~��E���W+��֖������c#���x��>�u	~S"k�W>1���ǜ�����u�}��쪑�+�a��x������]�G����\�����+Ξ,����>#�}�U���Y��#AA������������=��/x��|�{�W���v�����^石��EfJ���(Nl��?��U�
���g�ݪ�r`Ӆ(D����i!�*&u�r��l�P����~� �YL��j�1��D>�ɚ��_���:n7�'�a�>�|V��Bc���\�o���uU���@������n�\��P('��s}������=/I���j�̇�d�aDo�u~���y4=B�M9�/Օ�x�F���:{�EW_ồ�ݓ���Ѯ5��c���^@j}==?t�!	(�wR�Q����i�b���r�ɬ�vI��K�u�F�
�k��|�.b�
,[7|u���j�Y
�	<-�:�çE�(vLʷ�}x�=$V*���ݰt�K�)7��B.���,e򆥽;�T6=H�PRu�Z82���[7ۦv�9�1��-������HGo��\{r6���p�}q����l�q5�9ɛF��;U���fOy��N����X4\o�֋^�]�"}#���xj2���z����@���v]RVO6'ٺ��"<E�J������S�p佖��q�1��;ުѥNQcqUCy����{)��S�hy*�G������b�f�#�w��"�n�7���H)��B|��r0�[�^�ud�@}u�ɗ鋌�R��2�.��!�_�Go��%ڨ���Ye;>�]���.�[ݳ\�ψt}=��UXSȊ���2��$�E\uSGF8��7�?W��J'X�<ߊO)n��D��kԮ��g�}F���o*�]D�d
�ԯ[,%~���l$!������:�dv��B7�<����#��hl���;*숪�b�z� ���j��1�?edϜ[���8lN�,��)�y�3�C"=,�z'&|��	��v}/��v�r$��(@��Q��Mo�Ƴ_{����{�z�A��?^��v�U��$/I�aA�+Ƿ�{�δ����:���5��s7��yP��*>��(��x׋��+�U�R �л~����h���*M	�܊�A}�+��\g5�j�t{��t{H��M�75��ef�zN�ur�Ew��kT9���f�I*c��b/�s��v��K�Ư\�бբ~#����<��Ȃ}���&=P�]�Nx�K��m �<�	����H���<���3�C�
O��_����m�
��#<s�`+>�Ba�*��ŷ�S��r�`�1��e��m��緛�Y�Nd�4�}�V\{r6�K��|:N������SD�_j�댟�#�Ɏ.���=��������{`>��Y�F���Q��vN�ћ^�qޞki�0��[���O}Y���y�T���W����P�6���_z$�G������~a76��b'�EK�N�Xd�!�듓�W����`Zs�!��K9�ʐߴք��H�����Fk�u��징��D�/D�=���کٽ>}7}j9�
�g��7Q�n9�&�|�@{�r��+���.f�+8~Z�<�Ȳ����^����kJ�ɝs�Bs|g�n;�_S.}G�t�%Q�Q�����meo��J��xrKg�z���U�L\���:��^�q�x��yב��n��J��=�W{�،ڥS�+���螽����[�2ʗ8˜����ȁ�_�3y2��K��c��uN��>�2(�Mv+<ُ��5���uM�l;�V�B0-�W�u@�笢�U�^��Q��*�%F���Yq��n]���2�ۏUkD��C�h`�=f�g��YYj�MD���;pG��eҷ�$�'WR���7Jbbޭ��=o�v�� �z7�}Ǳ{�#��r�㟤��9��1p2)��^2���<���G[�̅Q�>���y���q����v��z�~���.�l��ϥ2/�����j��S��Zp=ʵYQ�j���/֑���#��Ѿ���T7��Iq���+�j�Y��do����G����ފ�vR7�a�/ơbW>���n#��(�?I���D	�Y���Wۇ���A^� {�K�P�M��t�82��������W�o��k��;����^=-b���"xw��Y�k�sNH
A�=�]G�"a14�m�\��d�-��ƺ��c�b�g����\�{�->)�=7��x��w�P7�T|��j��mf�y��=���F�f�<>�����Xwx�)�bǺ��O�R��ߨ,sT3�<��/El�|��SX=�s&EZ�t��N��;~���c\���3�^4����r��FBU���?Uh�j����IG.}@-!o�d���:�]����
�'kf��zM���Ǯ��3�>�~쨚~˔T}:�9���=�ز�sd@�	��XUwHR2����ޗtL�n�l�O4�y�m���wQ��,yV8S��ɤ�Eٛ�����s�&x�cYeR��z���\���GIg8�7쨞k�����՚�^��Zx0��H��v}+�3���C�*̕��Z���&s����W�C��+?[56���ү�+M둾����څ� T\�=0.w�9/0?y`�����!KKI���^�֣�`��s�RϢ��������;㬁���G���ާΧ7����9ױ��2e�i\��?e��]e�zi��8ُaQ�����o&|��b�ƨ�N�bE��ϥߴ�G��3�>�~�A��	An�4�I�ܙ�>���2z8:f�:�����yp69�tΏ#�sB�x���^)o����n�[
r�<�$KPg���Ξ	�Wޝ�N�U��{2�T\���,�Tw����s���'��q�>�r�^�,��2�NǠԾ�.ř�>�g�S>�ޠ<�E���\�|�g�,*����?[f3�
������g��c�$�����=��l��G[��|O�84pu�h[���	��2φ�΅R�Y�זlS��_G���a�?	��������Y�V+Ƽ�,=��%���%���)6�����{*6��T��8tz'�W�ex�XQ�܉���'���(";���~׌�u\P>�����%L?������Ʒj]���s¯�[�Y#�Ϋ\��'y0qoU����v�uf5���߳v�5Ybw FZB����HwNw��沸����cL�鸌mN�1�.�g����8;+�w:�T����VYu��.M3��l ��_���R<W	�v�J��d���.�O��+�=��>��U��L5ީ�ߤq�:���y y��J��@PjE�*�c��א�����x��Y�ʵ�S�fkK��C�uS鎇�Ɵ���Me(ڑun�o�䷜����㟫�O�dR��-f���VyO�U����Vuk�
v-GY�k�Ђ
��W��鎘�#�\��ڸ~ܜ1p��O�G7��\{r#k8�y�Zo\������sazD��z�j��ʟ9 {q���R����V	�2��!�����Z��yZ��i~�A݋��i]g���r3y�e��^U!����no���?Z
ײ����([ɔu��F�9E������9��Ϛ��\l8���6�V*O#�l{.;���x���Ek�%�3�ۗ^�ٹ�IP��{�b���L�L_�3��H�5���}/��ȋ���V�3��N����v�-�˹x�~�Έ�O����*�	��EEϑc	l�s���GFF��w"��\^�gxh��J7��B�OSp���d����c�P-��2�\���Xc�:��Q��x�;1�;�pvsu*�i�� ꥺZ���x�[��F(e\����������Ś�R��8�ˈ�n���9tŎp�f��K�	Y۹I|��1�l�^�{��Դ�4�:��=��O�v>���΀}�R.�[ Z+�il��#s����S�=F�,S��8נٓ���NS���1��q�:�ǰl���ʀ�>��`�M%���<��W����sGۏ�M������)�m ^o�������ñ�|����d~�����r��s��NWzoz���㻂a�P���*k=g<��/�@�ʈ��T䋎�S���Y���9H_ݞ�VQ[=�r �����	�TB}v�9��%܀������j�zۉ~�Sj� �\��HL�}��g۔G�.V��|{c1P�h�*a4�bT���iTWT����e��ܿl��P�&C������{��_FO�I��:���SD����LE	A��SY������r�=>��n ��X4��O�ު�vDmn�y��;��$���/׻��� {]��2<ꥑ��W|����w��Vd
Vb�g��~a76�L���W8���ݾ�u�`�(�3�ux*�Q�վ#!��7�ݹ�kE���<{"'�i��B{0G�6�W��"<���̲��ݕ�o\U��,T�(�S�W$���Τ�Q:cT��V�馳t�ϯ�	�NZge��Jz/��X���hC�w�<!]�dT����R��V��5Q�ԼԻ4��$$��_Mc��M�����x��^��4��>�P'�b��3��}H.޳wx���W(���E�re�y��B��x��d�W:��
����!Tɪ�[��N���9n��n:�`�v*r�u�4�Ź���9ƒ�sv봔ic�Bm���Ң���g�B�h���,��}�l�� ���h���Y¶�D�������?���O|����b� ��./�=�3r��Z����v�v�:�M)x-�������J�n֞�\��JI����N���st�7{�Aai�����qK�<73����.��b`5i�u.��:_d�ufޜ�T�d�Ε9��EF��e`7�H�B�T�ݶ�^��}�gᬌ~�5�t����M�)�vr,Y	6�w���vb�_g-�W�͒�v�a��y��#g
�^
}���(�Ў�ބ��]�C�PQ,}O�e����]��p��Lj�/#w}���E���΅�~�����lA�؛�ճ��J���ޝKu�ֶY�#�^j�i�p�Ka�:U�٧{uL}��8��e���X:�{13�%��5=R���#/�9�����X �E�ƎLr�&"LH_m������v�����Wp�S+f�J
ˢ�6���1ํ�=�t���.ý&����g���F{æ,)��7�\�D���dt��$�*� ����RΊpo�;�
V77�ķ��Ź��k�
ڋ��ޘ�F�H�N�\��dc����\;.�bD��+&��nV�,�f������rl�Fl���Ě�Əu�1�@(�n�VX�U�V�	��	�֡�.qX�u>ytVK�d�{����Z��J'D���'e�]�46^��K��:��gt�xu��R��G2��X[7�Ƈv���3��ʊb�D��t+0�h)g2 k6L����e��.d+�|���9�p�'���\_vӉ�/I�o�L��ӧ'TU�M%1�z�-�_����b7E�-��a�{�V�ol�z(KM5u�b�����+,�1�18���vz��{:���/x��(v&���S�R\2Ჷ��Ll��V���2,a�6N��^v��sP4�[ޙ8���ޱ}ۂ�3����fu��7���2s���A��7�BIP/`t�q$��r�{T.� ���X%Y��r>�Hk��b�SV�]R`��efg]-��
��Sw�n8)*x�|�����)�՘6��e&��y&W-��=�k��e��dz�%�xu����pm���W��,<��[��i#��H�,��˻��2�y�r�TS����LTWwUr����t���*4��yx����M����W+������f�k�\��)+�;:��tj]���[�s%�v�ܺ3��.�nt�wqE�!�s]�.Eˡ�Ü�Yw\��\7wl��V����Weu:Qlr�7w�]:�v�s��뮧�n[���r�MNu;�4t�W��h�\�9͹�.�U�;\�X�`�ӷu"�2���wqs�9�Qk��]9���7wV5\��wD�<nk��n:�NnPQ��s�5��x���S�w];�ѽ�����j��/�ɤ�,a����U�\��!�<���'5�1kη[b�uUc�%p�&f^�"���m-S���뮅@��G~u�^KW:=<z8��:U��n�#q��q�ݔ��g�_�Ko�9k|1��w�>>�Vփ�C0Οld��b��!9������뀮Zs�*=��r�)����o�f��eP~��uύ�d�\��+�� ���/��o&|�Ι��k�8&�:=�a��]�}�Im��B{r��{��;#ʏ�+���r$�.n*�
<��L��2�����^X��E�u�+�N}ҝ���D��c�{���A�S��v?Q��Ù`>ɨ�O�	�gڂl:���m�����=��>ل�}��U�t���j�X*��ᒫl���|}(z[��J�[�7��7|���ޝˁW:ܺن���w/֑��GY�A���[��Ϥ����r�z���j7� ��~#4����E���h�D�ә����q-,����J7���]Mw�ם����򃬁�N� z|e����W?S��чҴ�/~�Wҗ��*�u�XR�ν���W�$A��>�:~���nk�@RDz�=�l�SU�u���d��B�F�������Q�YV˺]��h��h��i,���.�RJ�I�9׼�t1�H'ϔs'�%wP#��G�2c����4�"�X����qWaSG7�"����N��Vh��WX���p��mk���,V7Q�s*J��rb�'V� b�sa:��O���s3�������/�)ߤ����*<���)��;�M]�܍����WI�iJfr|=qި��6�Rj��cEG�J��Yo��9���K�*Q��}^�*k��i����a��]ܚQ��~���o��f���4���t̲:W���w��g,�z$����"�ONz��2�3�5�GW�ϷkCó�����3q�1|�q�fs��ީ��|K��B�����O�a�Ͼ���7>�Co��#0Ε�d�V�dg���6�;��}~��vN �,{|3|Gk�����ʉ��nx�xg���FS,^�֖/&w��� k�#��j�hDG��{r��x`�@��F����/yu�b��l�ީ�%g�Q�5��ɝg��2�$A�k�R��sF�^zH��~�i�9����v������]r��Nz&� �Q���>��{//U^d~�ߘ o���3�o&�s
�jU���#�:�����)W���ϟ��q'��E������e�ǰ(�}�WO���?SW�Rs����a8��#����+K�=Y��^����J�4=8tO��u����a����j�P�Ue�'A;�ve���Q�G� ���u(�*"��� 0���|�ֽ�XR���F��l�h��*Ĥ#ܹ(�]qW]2��O�8��N�w���hM;��|�� ��qܼ���]�od��l5tm�/�5�Z���8Û�m�����J����>t쪑u�_\�|�f�
�:�<~��\l�:���zq��{8z���He߆�%j���IaA�-0X{�R2��^++�3g�TE�psH��3m���\�W��C�xn䢥�#��fAn��Y�|͝��K��8KGv=��z�`��ڞCN-��i֘��7��C*�6��l��� lW�����A���S�X&9���tv�|}�/;sdW�A�����G���I�����/��>.� ��6����T|WzϤ@�����B升�\H>B�;���l��O����zT�����~��2Ǽ=���NE͝Csg�z��\2B��U�9r=�>����ͭ����cL�F�=P���>��ފ�.�
����ɼW���ݢg��!d����Z}?���dUu��l�a�8q���K�z����P�G���[B��]�~`V�@/i�O�页~Vl�}��k��l�Ϻ�۳|XY�Zo\��y::���|ô��$��}��4���}W�]�;}��\/i���ueT<9;0�9�s� >�uW�Z�Z�W�f�s���$�|v���2��#�4{e��8N�tn�Ti�eԺa�;L5��W_�]m��5�*Ri.R�$U��V��J�qu���������g7��7#{�: /��m��i@���������m�%[���o�ւ^��4r��c#pKz�*o�nF��z/|���yT�ψ�Dk�����M�ap7�,m�ޫ#�8�\w;u���R���M���Ǫ���)eP�����4_+�q�)�a>^��C|��aQ/Ǹ׏�Y�o�s*U������g'B�ЯЕ�U�s�-��Rٞ*yW>E�ɖϹ͇��8/b�th�T}[388���b�F��Mi�r�q�Vz��eK1��S�<��U"�����t��P�/_}�9Q�Lee5��eB��`�kv�w�)���t�W�<;�;�p�l���ʀ�"�E���4;˅��|Z��A��k�J,z���N�����/ԑ��P/=@`���t/ޯ����7vHO���{�mË���=|�ߘ�D�Ñ�w`ǼzuC�}~�Ϗ����@{����9#�^���t�Ĭ$+�5�E�{+(��Oi��;�>%��
�\>�f�.s��rVP��wv^��������$W��H�D���ܢ&(���w��R&)���g��$��64�׷A����g�,S��	Z෇,���<�h��ѐP�	'@�f&�+(s����W'ls}C��*�0��	���ε��ʗ�^��j�1噱e�M�H����ر+fM�F����T�Y���/5%�jn�<�N��M`J�]3���RU�ڎ^��C�S��LΝ��7� ���lÝM��H\Z��?�T��ry�zL)>G{ꬸ{��_d�t�=;�Ǳ���)_��ݥ�3���%C��Hf�^��쀶�
��To�>G�f=�7fDf׸�ܶ��vJ;R{7��p�r��xL:�!k���o��z�~�.�Վ���������������b��yN���h���5U����=7Ԁ��)�߈P�xJ7��_����p�'���
�}��F�麿H����}+�F^V�;�tk=7\� d+�g�71�o�y뉤;���VA굾�^!P��ԇ�%�YLed֗-,��g��xP�s=(/�d���2��f�d2V��|y��~\}	�G_��xթ�)�mh*f/.{ŋ�&u�'ȵt�w������6���S�=����4{}��n%ڸ����Du��U"Q�T�U�5=��Lա�}�W�Ѿ��o��^����}��^���;q����e�4n!z�q���$�Цx�j2���+����_��T�l�� �JR7c�j5���"�#����Th�����dB�����[����e]��7+�6i#ȺauJǢA2��ܹ9�P����"��Q��b��Y���7t5q��p�>�&��S��[�<\+�fN�c(m7��!�z��̾s��e�n�=�f�r.U�\����^)QV����ӧ�B�(�gd��On�贡}^���dUDKW�W�>�چ�_L:�M{;��qg~��f{#}lb~���s���3��V���+�%�:��9
����GTϸ��(w�i~*/��ܾ�x���n��z=1>y�9���[1=|t�j�"��JL\&'���슬&�� u����w���z�\������^�����1�m���ޞߕ���ޫ� \(-���ud����7�ùbeG&�x�5���:c�~��8){�l�A~��8�T	9~�Q�Ϣj��m`��|�]9#TM��r��8�HY����F�꿢:��J���v����PYU����O��5�\�^b��[��ܩ�}u\oQ�S�-v�C�ͦ+K�f�2���]���|m��O���h�T�{����/���\��X�� �ҽ*��n:��77kCó��X�4��j3��o�R�����^����p}yw:}�"JҢrPۇ]q���V	ñ�o����
�WK�+�h���n>��A�=8��SJs��p�~ȅ>�e���oR�!Vk�埌� 5�u�L>΋K՝�:E��
r�p(1��W���%U�,�-^�����w�rԈ��1�U��<��I��Hgt��S��_�C�Q�2�㗛���,m��br�]F���w�!��uEX��9Π��!S6s�^\
]k�Ė���[eK�G{��i�zwsZC�S�m ��O�WޞO���.��^=4��g0�Ȫ������nX"��X���[�}�Y#_QA��#�n9���>�:�=�������
Af�T��:��]dm-�WgM9��䇣 �����>�9�U��~�⓿\�	⨮}E�=Y���Ǎn��i/��������J`I|����9}�y��x�^�q/�����.�^�z�Z�w�+Ъ����fϕ �"�E�D�`U�Fn2PꈿV�p���遑�5퇷���Ys��"&�z���޷p��k�Xel��H�W�����c��GG#9�53�p����g�יc�(�~�:o�0FD?S7"���:%��W�_W��������fv��ч�Mo��u��1_������z��č�t*GxSF��H^�c�F������}
(�p��FG2;>��
�iU��>����*-߮@��i�^�ށ�[�U�Ԡ���	� ����nQ
���O��pvT�G/\�o���u8=�n}h�@����^�$����iy��`�����d�����1��l����Yxh�.-����;<HkHcgf�#�V��66We<&M��WLJ�y:U��ĳ��!��d�ƙ�˜��H*I��Yٸ���rl;�s�Q����|O�T���VTe�e`W��f�6X�3ZX�|���w+�鋅�	g��^���$*�z��>��^S��^������ʮ��s��Qg�:��g��'r0GH�߮���}{�U�~������Zf߶�\y<�Fϲ���Y��٭#3�1e����雸|��G���?g��@���j�G�^���!���s�U��;=��Ρ���5w��k�@�q~j���H����� ����]�R
ײЋ�}��Zos�S(���|,'�����҆Sՙ�\�S<1շ\�W�,���~4�t�g���.�Q��k��Z�"�e�7�E;�z���C�<ҩ���WU�M����,�\Ϲ�}�BW���8�/���K���Y=7��h�f�~L~�I�k���Vo��f�\��*�	��DT\�/&X�ƪ��s����]��R��e��{�������z}��Tï�,�p\��9?����x��r���v���H��"�#��������Z"��+C5���do��~���Cs�\ţܡ�����B����0��Eep���-�-V��辂�8�1c��Ʃw,�\�C4>��(,W��3��H�o"��z)Zq�g�J�S^e���Ԩl�U ��WPs)&��b��Y]��Ht�ƴ`�)���e��[�[��ݫ��G_q����1�T�W�t�P;�Ҏ��Ὢ���)�+�G�q�6�ʾ��,\K�$s�zP瑯��߯Fz|j����~�w>��Cz��Ѯ:4(��+�d����Xp���~5��w/��9��W����=�D�o�����Mi��ʍ��_+�$z1�g�h(f�7DLR�����s�^��G��S7�+��QP�
.��w3��c��/od�_O޸����ϗ럇_Ֆ�cl�u�}�� ��
�C�/6^-��V�=�����A0G��nt�l�7��(
�<�I�'����<Q��]��t��NKFan=r�����4+�4O���U�}�H�_/M��=��/@�f���m��m]fhuԈ���gT/[9��(3ҏ���5��xt���]U,���zO\?U���w��l�G����E�L��9ڼ�;�/w�*���M�R OʽQQ�վ#!ҿ
��ʑQ�և��i.�uגi�k{h�#��d�C�Y��Q[�����P�aP2�z���X�Cs��ܬ�r�5�eVy��ii46}��(�=��"}85eSQ�Z]��;��!��
�VzP�����~�C%�)$����u����G4��*�
w���~�ѕ^��r���B[�5�!�lYc�B�W���"D�H��7HCA��I�7�����c��?]������g�9m��������JťJٝ:�[��$�����y�Υ):���_�ɝWСQ��NU��{��?^\n{k8�b����Vւ�*�&.{ŋ���p�"� ���K�ȩ�j��١��T���}㞹zOWTg����R%EOUX�Ox��cڬ�WO�M�=s��i6{�Gѳ:<���b�_�FF�}ǲ�îe�®�~5=��/��qA'<��D�+����J�%���{2���l��aq����@N�9���ݿ:��z�7���Ƃ/ڸb�?��z��	��C����E���p,�s�Q���t��#��y���N���W'ċ�\���#o�^^�O��G�����{>��S>�w ��9�l���w�� �����Y3*�U{��ܑڜ
�s%�\旟���uNL_��>�
{�&��Oa�xY���������Z���`�OW���^&�ޜ������չ�I�T%�p}1�sD�E>��sY�V�����ǋTW��zEg�������.�f�~�=9����p=�D��蚻���5vGg�>kwx|�/}�Q�����cB�c��>*���l_�c�~�qYU@}6k}^�M�C�\"t���v㋮��������|�GS�$����]n9÷��︽�|Y��tCP�����V�)�B
�sT�дp,���)Ҡ�F����k�(�v����+�n�m,�k��g:x�����H�:�m&�r�n^>Xv�Y����T�	��ӴQ�}f���1���-`)�r�ٙW�_i5~Tu+i�fegG�(�z��.�X��1�٫�R�Iz4�,t7����L1ټ?o'gN߆:���Z*ዬ�y��0(p��5�:u̙ؤ�!P��:���>�	[�#.�ZgfYQ��t � ��tb���Nb
&Ւ�3�X�-���x���w8ή8Ԥ3(֨��'����ީ�_wlEǁ��t�bXU�՜�����U]�������J��)Gs�k;h�Og+hp� �t�ܔM�"w2�K��d\��M�����J���μ�[9����V���ǋy�/t
aJ�f��u�z&^ f=�f�$Z�݃��d<�r���r��M�lg��e�r�h1�Y�[��K��WD�0e�aQ��C�����Yܡgz�&�V���4v[CH����1	Ġ3�շo1l.t��<��㧭�#N��cQXw�'�Q>���v�6Ѱf��eu��m��Ү���r���&C��a����ڈ�l�Nb�&>��(�lU'E��R�Pv.�2޸�p֮+��1�l�K{%2G-�9|�zѺ��|�{�x���e��>IR}�2IS�.���۾������s���捑����*� nn�j����H��U��q-�RTl��Üf�%ݙ�N�54V��]f�������I��5<&h����_QC۩�������&Wb���|����X�U,q_#��D���vJ0G�CfX��u���1-5��3�_,�M�8c�#����ӌ�:��*�7�I.X8-�2m����\d\j�jV��B��C;,��F��)���)��rx������<�Y�]�JwԤ9c��KI�8��]�F���t/w��]W|����{�H�Mt{�0C��!rB$���v�mK���e"�n1�Ϩ�+��]��SI])]w;45򃑵��W�&_Y��x/�u��_��;��8c>��-E������{���S>:+�@Y����1Zr�5��f]D�L
��S��af�̖tJ��\���F^����A�s.]��71��,��{����V\�۶iCݛՓ؄i�[ �l��v/i��Sxjh+�ű���������8�;%������k�v|�aZ�h[�y&vaRr�����s�v�n_�Ӱҩ����}���Dkз�kq��4�������&շhʾ�dw��L�p"%.��Ím�.;�Kn;!0�Ȧ�ڻ5���adMƨi8��^:ݪ%L�c����&���-}�O#:�A�M�|���;��`}���F�����KO��i�"(��j-@f%x��u����~�wEȸ^���4��s�m�N���s\��J��Y7"��L��wuc��&�s��!�����1�����s�w���\����pq:�\܊9��p�<��%�Awvፄ��f2���]5wu����wG ����w$nh��%s����eˬnWD�ݲ�������5��U��˥������!�k����;��qӧv-�tT.�wu;��s�uܹ	]������Ά�]+"K�λ��Ee��\�]s��X�����u&��;�r�һ�ݤ���;�t:fu�Jh��q$��K��r���]wd.�N�N��ruv����H�u�������s���r��b����t0\Ms]��m˻�\�"p��Lh�.��3�j�L{�]��*y�9���A��ͯn��6������V��Ȥ®�1��1��9ca��㏹f��8����v7�f8��B�K�g&��f[�US�i��n��
�����wdg�ԮTQA��5��܉�Xkյ��{9]7��_iwyS�gf��|V�	�?$�1o�~�����p/K>���~��y�zpt/Ըd��e\�W��Z��C?)Z|�q3�.����Qn�߯�遱�^ns�v�%g�m�R��3��;��ui�?N��Xu��6��.3v�M�~Uf���T��� 9�����u��Z�]e�zi�vOmT=&��P=J�A�q�OT<� �h�h��Hc7�O�T�{a�n:߮�ё�%q��ڛ�}�k��]�c]~��(�p�\��c@���X3ѓ,/�0�4���?J�Kb�~.b��p>��^EFW�_o��5b��Έ�g��}9l
S�}�o��9�^ۊ�t�c���ng����S����o<>�>������>d�A�Ϫ�]D�`T\��f��C�/ա�x��^?W�5���sS�U�dY���=��_��k��w<v�%��:%�q2�슩S+�a�>]���ܞ��k`�U��6(�fOÎfʨ��+�H^�,ı��ˡdd��cGa���T�R��^����U9J<�t�.nK$�c�w�����3�+���;:c�{up<��P�d�ᅾv���A{�8$���.l�t�r�՟��l�b__�c}�����$:�����B�^5�s��۪�ט�M�zB>���q�.�z}���G�����C��)���n�H�"`gz�S�/v�9�;ym�����}X&&��E�����a��
�>�dk�s3`�*T-�Fn��x���J� ���TY�g�Ձ���#�j�MF���r	xj	�_r�͛��@yTU.A����r�Å�9�26�B�Ӓ�>7L.9U���nևq��Q�ƙ�{U
��v'��u��ܘ�oNur���IS�&t��Z� O��l�O���el?��<l~+�A?	c�>`�g~_��=����ѽ~�c=8��������ٵ�����n"}!��\{s��ǳ���S^�V��QL����^d�^���zO^�oD�~�Z.��q>"�9�~��]� �{�t��+�:}�Q�t��o��O��]P������W]�.7�k�`�Ӽ�!r�\v��,���{Ъ�i��QCk��ۏa;����&o��ێ�0�y{c�q�Q��N.�~tWj'����\%����n�3�w�s��Î�vr�9�vq[Q9R��Ĩ�[y�j�\�`&���8�ٙ!�.z��x��moXq��5���""�u����.�o�;��p�1�w|�@Y�B`W4H��R�:Tg0�i'���V���[�
�p�ɖ}�ڐ�Z43@Wz��ɝs�>Nr8�o����yԉ�ɒ�
!
��Z�2�/�<�Ȕ�/~��ϋϷ�E3K�a�UXSȊ���,^L�}�^��D}s޸�yi������L���G�������U�,�f;�z�n@{�UX[ &ǳ�၆�¾�������y�h8W��׺�u��1���B�Ƕ=�j/���<G�`���O�{���oH:�c��lp7r��E�چ�.���I�z%y����^�wCޟ� 
�ޣg8�v���&���|zH�t�Q��>v�����~5�Į:W�7�<
�����������9�_j�QGY�$�.=!�̮��&����>Gt���{�=r��}��nb�n�����0_#�}+(q�dT[���j���]xo}�E2���~���J]�G�h�V��A�{ϭ�6��l�����Ϥ�_{�S�d�C��6�;���;oG���ע�纋��.�����(dj���t��u43���z��F�'��{*��痽�x�
�����*5�\k#���q��>x33� Ȣ�&� u�Zx�J�Ȣ��Zt�;��L��'0��kugf:kؽ������U9��뤀��z­Ζ:��T��yөV�+`r����{1���y����{�7���Ky�Y�E������7f��<��0��Ө�3����Wu�.��E�W�+ޙ%�45�&Qȭ��U��>�T��fZ��fr�;��ڇ�3�t�Ǧ�:�aW���:���U�<n7۷#4e�Cw��������s ��yD�����2��d\�y+�����3�Z}j�%_�<C���w�o�������n�Gm�Ȭ����d����	L�vg����ʧ՞C<��P���]ͦ-x�ʜ�emNvU8��1 ��ܯyʣ���7خ;;�r���vKg>�mh*g�62U�/&u���r'�x�g�t�e�KƊ���t��_~�ѿyϸ�}⾗j�o>~��)�6���)����c����%e�gk��9Ÿ>:pz�q���O:�/��ё�^El_�îe��B���Ӝ�W=������ϖ��f$��@��MF@���R��aq��z���]$s�lW�],`S��𿦵zl�E۬�>�z+��͗��{�<XfA������.�a�[���l����3�Wi�?Q����$��΅�C���%��Cf���I"�UyϠ�g�>F����?���vs�1G��í�6_4���@׷u�?v��xfu oI����'�/��Œ-<�f-�Q�Maǂ�O!P���7����#�SS��6 ��#Qfu�y8�[|�Xo�I�0����ܖX�:���k�����\�ӈ�}�������uNJ|'��A�(>Ȫ�f)�x��8����t������J�ǻ��OS�����S��N���pcm׉�T%�<{7�XLlҶ����3�kԠ��]j�;� KP���P�U��_�{��`.�~̀*-����Q�Yt��xS�G}��:�twq�H=��z��u�d֟i�\GS*Y�.9z����޷5C<r
�v�4B��~��z��M�v}SX=�7v���mzN����C�Wt��.��}�x�:�l{E��zڕ������[F���%��������gd�u�\n4��3����~���~�'ݱ:Gz���D��2NOl�e}�s�� ����7����X�X??e��d������6��S�����s��t��۷o��L/a��|E��.��Cͣ��:vہc_Q������n:�a^��x�E��W�Z�%Vѧ�#�;��<
~��~�Y�}��}��^L���!�߻����OǶ=�ï�-��^��f�GxОn����T�捧������Ns�Z.6-J����N�	Hj�h}ԟ�X�^װF�:g��ҧ�A��	-�hL���;-TX:�61T�S:e��;���)C����)�-�>kE�ذ~�My�q�q�ށ�@7�x;ٽי��5��j���ӌ~�W��o��^9	UD������7=�z�'S��ڷ3���z{э�u��-)�W��	t]p�Q�&�\
��&o��9�����Ӕ����1��w�Vf��eq�r�q��g���{!���:�UH�偑r��5���h�z{Dx_2V��i2⽢޷m���q_q��]�=�큲��_�8)���n*�uL��{`{%3���3ٱѕkyNs�l_���t�꾮�u�PϽ�\�{�������W���'��A�(>�;:�]$.w}���M��S���[�܀|<�qc��{�����h�������F���؟�BA��3�>Q�=A�=��V	��}[�	���G�a��	�O���/+�ӟX V�c>��uG�,��^�����>��钊͂��m��U�t=>���T&r�͚;�t̫��a�������ee ��|�}*j�Yr9��6�6�;��q��zL��,{.�L/?I�~���ő.+�	�w�ު>�~q3��^��������C/I�3�*��ܜ��w����اiB���Td4�M�����Fi�z�(��¬��S��G�:�;�0RJ�R�(��_v��Hf��/8u����]'pg����n�#UM3�S�]������+����������ԡI?[i,�W��"�$V!��~S�;�K'l�&��t�>����l)�S���~22v!{rp���-9q���\{V<�����骞����K�6;L��,l���`O�i�+�^���U�=���!��P��������:��܌�i�O���}�Y�� o�� 6��?+�{���R
��Б�ٶT��Yy����,�}C��,�|�iS!�ܭ�w�;鿣K�������;���Gޓ�G:�A��|F����.>K����(�=�e��K�
��3��\;ɝs��L��d7!O�O{������%�>�x�;�S�ݪ�������"�.�=U`Q�E"���^y��L\�y���h�s�+�`P6=��Wqϗ��m�+�XUc��z��Z�g�V^���^Θ��^
v<�G�<��]dFׂ�N�:�hf��q�����p:���nf�4�齁�7�є;��l^��*[�+�>���u�q`�JG����=@`�e�����]kú{n\+����yd����>��B}9FFTK��9�w2#j�E�T2����+�Qp?~��e
��W������t�ئ�usR��5�=
}�C��3�o�a����V�5�b�s��݁e��ߒ�D�*D�zC�kٗ����3Z�w�q�5�hN��v�>Q��,N���6�=b��w�����5�f�"����+%�.�ͣ�zա	��`����gp=ő��5e�Vꔑ'Gŋ���dVQ�x��wH���ǌ�������W�7ΞMwP_L�a�:��� .��Ȩ�U�"������ܢ&��4.5ϸ�������=��ۅ����9N���T&2�����l�u9���P_y׉�~��ۨךz��i�~�;y��l�|�-!f=�d�3�����CQ�XȎ�c��#�/�T�ʵ� L{�*7>�#�>Mi�5�V*��#�ws�0{Ѻ�0��ٴ��s�vX�US��3,���'���o�|� �hKcߛ�(_�"��3�~�~<Q�纺��s�ݨy�8p?�����~�s�\6��l�R��Y��FV��5[>����|=����¢_Qem¸�Ui���7�q���N����$T�-����Z�>��g�W�|G�7������@k�=ː*�Պ�/�}kif�댙�L\F��ަ�i�{��_�.<p�:`{��ד�Q؋:�|��Y[%��9>�ߧ'S>
ʢ�ğ��ȑ+lΨ��;�K���Tx�e{�G����Fo�y�ey�v�7>~�af�T�Ĺ�\�$b�zW�?�͕����v ��5�u��Ѻ:�T�x��^,��ptt�̚��uLe�Zc3[�h��td���o�C{����͈8h����kx�S%L��]V���WM�2��5+y�8kNk
����xpS�2eD���S�F��v�w�����>��^�vXQ��z7�'�y�z�ĪA�^��� i4=(z����7��f���ڟ}u>����^rx�l��*7ިw��G>��ݾ�4r�3}0���ҹ���j�A��~���d�����N}FE��E�~.�6��}��?[g��������֢�G��Q:=�_��Iw���S#��U�r��l�V�i�?a˜�y��P�}o�^���sޝD���{,��T�<�_����Ș�=�g��=��������==�s��ג�L�9��|T����� �E��s$��<{��(�g^�#=y���>dǽ�[F�z}ǰ�����i�/�=�Y�?f@���X�����]g$��jY�����
�Vɯ��O����J��_.�]aȇ�ə��lʳ!:z�tX�b��L��x��ώc������dü�IZ^�5P�j�1k���2Ŝ�xMzf3�v�k�K=�8��6n;�%��}^�}U����Տ:�ީ�߉E��UA��w�JExW`ћ�F�[��=�wI�ߖI� �m@�oea(�b�I�{�ޤ�5�Y���BoU:vLv9�~~P��ѮGe�qS�*�[�tYڒ����w �:�����a���]c��h�\������i�6�:v�1�B��]YҺXaB�٭��9��`�����H'��O�P��u�n}�\�d�>)���N��+�&�mb���!��p9K�L���NG{v�w�S����_O�aՕLb�.��V�*�swx]z����Ի7��7�R=���
�_�ka��V�y�vǺ��Ǧ����zWb9o<d��Dϻ�s1�}��b�g|n#= 'qR��{���ڥ��{+î<�����S�3UQ�|�Z��P~�ʍ9�T�ed�`}�q�P�s�s�ahS���~)]��yOt�z73�7���/�hټ��K=��N˦�Ϩ��r�s�����k�T<U&E���������~^L�,>�q��/MB�w��䣽����@>ʩ_K�}r��5a��\ݟe���M�\��2+Ѯ�u�{޶�gzw��5��^)���[==@>�"���7��oK�@��4 cx�*i8�F����9���/���N���K>�A����q"����YD�z"�.��v阘��+�h������7�-��L9��(\J���wZd'z?��w��j�ֶ����ֶ��ڶ����ֶ���Z�ֶ��kZ��Vֵ����ֵ���[Z����[Z����[Z����[Z���ڶ����[Z�ۭmk[o�Vֵ�����km������umk[o�j�ֶ��kZ��Vֵ��յ�m��1AY&SYɊ�1�Y�`P��3'� bI[㞕ET*(H�QJ�"�%R�BB�
�J�)JQTI)(U�(U	EJ"R�TP
��DT�UUIZR���*T��kX�eEP)"	RHH"�UJ�(��	JU(ERE)UQ"E%�`EH%�D��U�Ԃ�%T�*AT�*�)��IH@��P�(J"I�@"�(*�l�@�H(�% �P��U4jJ��T�V�  Ө���9Y�:]�\�IP�wv�H��]�+�5M��TsR�mu�U�wT�nev"�;��tV��B�QP@T�T*    �u^5֎32hw(�4�]o46���(��(��袍(��;�X�(�����X)B�QD��s�I$�(��9���E �v���(�K��ᤅ-�*����E@<   ΥR�yYsB��n�Tv�J��*IN��SQMv�\���iݭtX���vUWXqm۪Δ�B��u�v��U"4E
��B
�  ��n�a��l����gv0���uUn�ۻ;v�mv��H�m�wh�ݷ�S�ݥ6��ݶ�.�N�������u�h��wku�e[Gr�*j�N�:pUU$�%DB�Hx   9w�ۮ�n��WV����L�j,�v�*�ʭ7n�m�mգC]�m�u�e�]��4��wkeY�n�v5�m�aӭ�����s����m�����)$�*J�U%P��  sy���m�j[��(�Ws),u�fλ�w�e���ݻ��nw4-wn�l�w;[.�SK�3wYˬv����;6�t-��vֹ�Λwk4ۮ�)���GM$� U��  ������ݙn��)��n����t�;sm��[���T��@�n�r(�GdV���c�ỷWwn�'wrqSkn曶��鴶wKu�gh��6�.�kN��UQUI
�@�   m8�Ͱ����k
s���Ε�N�5[m�*˝ùlmuu�m�٧s��wm�b��v�nHUS]j�Nnn��[�]�[Q��KmssC;kk��è�UB�"H�)   ozZ������W]۷f�a�We�����[��b��\Gj��;v���.�Ν�]�9v�]v���t��Mۚ��V鮻36ΕIX�6�eu��]ê)R
ђ*J��@�  ����GV�֜�Wv�[���7(����n�ۈ5�n6����7-���[���].��ݨZ��V���WC��̦�wa�ݥZ�	< ��*JT � Oh�JR�  Sa2A�@ �JU@4` T�I���h&F@	4�e6UTڀ��\��F�7L�I��+�H�����h+�P?{���l�������$��Є��$���HH$�	'���$��BH@�2H@$$?�����wY�g�WZ5��_2�ܬt��d-:w���Ь���E�����1ûr��a�����9WwK9��س7A���~r�*���~�F-3㺥�yiiup�n%�T�$QwEW��,���V��P!���F�%b�L*�搌�@�P�<N�b�b�Fa��2��cA�pL�/�˚ڌ���)�eO��w#r�Tn�BJ2'��#6^:]ɉ�b��0�����ySvb�	k����俉v@�˦浻kf�5P��#m]���w�6��ۉ-�Y�N�Hܚ݉xm�5�k,"��+���+�( �+7)��X�f���aT偊�Ǉæ=5�v�n�L�o,�5q�f�b�M�V���4�)�����5��ֺ�*�'�Z�I ^��Du�@kwv,h��шە��{��́B�5�i���YG7�Y+FS{�24�-��˙���8޼�)�VF�Һ���Œ��L'��sj<Z��n܈�� h}����@�)!V����;�Ȥ�X�q��H:ư%�&5�z�� ,�$�j֚_*w��l�u��4X`�!.e9h�՘iA�4�l5)���q5;�%��W�E�h�r�m�ۘ�(����Nm4��Em�Ϭ�S0[���ʁAz��X���M[�j�)S�'":�r��[L9���8�6ذUZz�EP_��ˤNM$1��:�K
8�;��<��qIO��P��fU�T&asS�A�ua�ݡv��%�٢��E�NG�C�z�U�h\]p�6x���B�+:L.�.�iAzЎ� >T�3��82�*>�	Q�Z��D,�E Q�;B�-mi����Y���M�wvu,�i_�&��Vp赔v��9�uT����Ԭ�5����6���*v��Xtj�f�m�l����B�ސ-Tpҳ���䁛��NQ:���s�pL��P��H�����^�ǰ276���TE��VP��:�7*�ʒ�˘b�ֆ>wf��.�I�4qJ��k�ӳRYrSa��=X�[[�֢ji'.�bj��W}��WM6٘�[H����w��g8(��í�z��u�k*�*�]G�Rz��Z�#�%�-n��F����TSt(�b=�R�K-�n��R�O]Է��%L����h[�3�m��"���1 K2�����[�K)���	(j�c5����YQQ�PXb��ӹ���j���T������ �CF5�����)����PIQu."���V:�&�)�:�1�ܻ��\�"ʺU��+1��[GLEL�YadD��fa�4<#:��ѕ[k.�kbc�,����E;�#p�*9���.&����w��"ԫki6�IN�)+Ԧ�(��͌ұ��FR�+k�7JU��[z��[p���L{ �pJsP�bxe�����HI���[	e��M�q#JZjb�Bm�Á-r
�LZ�2�eV�w��N��)8k!�X��&��	FRsvi�v�yr�7�|���XSL��,;cu�`�[��\�i=;�MK79Q��f�Fk�D�懠L3hR�L`��� �۔ �8�pm��h7k2��ݑmSq�`5u��IOJ:������s+h;r�B}y�R���	��tr*�Z[���H࠙0IRf*���a�DM��WoU8o.7��9�w�&H��m#q���9zl	�F�'����Yuyvq��bGgK8Ϋ�%����.d��aln=na'
BɎ�x�]*�P�_�eT�X��jQ��NQ�FV`6S�U�]�t�c�D��[Q�4�aJb�o�i�X�!h��nkU**O5�Mbf���u���т+,#�'J�tk�`+Or:.٫6m�MA�.Ʃ�)�r�
5x�ېEO)]�d*̳[�\K,�K9x�VRRT�ӺkR��7���5�3��Z�on��V��٬	h�ʱr�\�jƊ�i{pCb�ͨBѐ%i�[h��h�L!f�E>�B�YoN:�V�bw��_E�@d�~�V�T�Ō
$-C[�MeXe���4��6�J��T�p^۽�D$�*M׹�f��"��h��]��tC�V� ��A���mk�5�T��Klk��h�"�n��v�JW�ˊ3ܒ�K^T�f���)'a��)rۃ12���Cb��h�+E�>+����
t���:�&�5.��u�icbH��a]��
	���
L:𙛄���z�ĺ)m�@u����&hPmӠܬ���+��Nġo.^:§�m��TF�lhT�L��*Z�:�1k�4��-���6d:��)@�dJ���{{Rh��Q�,@� Z�Ә�R��Wbx��iiR��femE0�B=�Q͸&�n%I�ۺuj��ϑ�R�X%C�J�Ǣh���ʼ�6jQ� %�(e[W�f��
l��[�X����n���`"��-�!.�a`e,y�Ee�C�� M-"R��N�`]!�8$�� ��:� �Wt����6�����k`#[�++tJ�]X�&ݺ�v��VT"Vƥ��:���'���u��3�E�wy�RQFRZ���:Z���m��,��u�Z7+*F�E@.�5$����r��6(j�%M��e��Ta��1Fjˠ�MSw��f���!�S/b���BVѡ��۸���k��#s����-[�c	��Y9a{���.�n#n�uM1V����8�r�ۂc�(�SD��ہ��ْ�%j�Jp�V%����ڎ��fr�o �!��'��bTܽʲM�ؑb9p�Sr�i�H3n���ĝպëXã6�lti�%R�M� �f�l*-�U�DK��SZ�\�Z��]^�F�(5�`=��eS[�� b4���ib&8B(Y��]a*L�!��y�5NL�d3B�+����hȕ�eһ
.�ئ���2xu�L��6�ޚ���ՂhY�&�5#wa�u�l;����U
/oa��Z�AH��&�t�t�Z0�l�mYӡ����_�ᅔ�ǫ-<��E���j���J���dk�yR�7��ZM���ot�[X�B��Jݯ���#CkS!\���-:����2�v�0��^H�-&�CN;A��^K���H]-�S��?��$�G��_��Etބ#[p�2���ъ�o�z�\�w6�e�L][�)f�V��%	A�n�d���eX�ڊi8��Ueh�E�
�$�R��N����kq�!�4��(a�*A���-`�2Š����J]^`˺E�s"��z���}p�vR�Al81�Z�`���	en��f����6J;$�4��a�*3U��4�eh���p��4;$aZ�e m��mC���)%�Tͦ��������Ut��n�6�-���<�HZ�N��bk-���H�m��n�`a�u'uF\��fc�B��ńmb����@lݼ��͸���0�i&&�j�h��G2ה����ޕ�!���lL��V��r���YH���	�7m��K��qۉ(�hrV;@l`ZPm!����\�)37#��o�n�Kaca͠&n�"�̙J�����״�&a{4j��6��.�J3�P4)��]�c�zܵo\Ԇз�� �x�:	Q�٨�5����P-�e��Y��T+�k4�"��J�h�;)k�@L's~x��v�cn��/��Nc������v�Ƴf��[E�z�GMU����� �π���>L
��6�
��ZE��j��;@��FaΓ�ey[��Du��2`�n�������0ؼ��_��Iu���4H.5 ˸�[���Ĝ@�B����8r�Z덌��:���4Y��J�zE�~�Dc�qV���m��t��µ6�F�z��x(f)�^e@۸�0'ͬ�Qr�u��諳��h�4(��-^!R
HJ���J���UaNG�a�����i�(��wQ��Tkq#�\CT��E�-����1��8�����j���^��V,}��*�2�����@��%�Z�H3wl$B���pI�l-,
n++�v�Q�q����O5j��\�[��V5�k�kv��0����e[L�c.������Z ���q �I6*Zn��f�)Z���E�C6���L�$e� �B"�㖍�ٸsZ�/r'��ك�!Ime])��`+�)�O6�S6�IC�wt��`U�!z�[lhZ�f�0�
�$�ʈ�t�3����)l�ܦ.�����.��	��uy��!d۵D�hV��rq�-O�k�-Y��$����;��j�ӭ|˙��oj�wV�+N�/-�c�%MV������6l��jQ8�8�ͼٔEe �6���U��4�:��i��Dd�J��^*�)�+e[؂�^et��O�%Iy��h!sik۴�d�֍LؒqPu-�hQ�n��{RQ4��%�2]�e����g]ݬ�E��n]鹪�����F�R�˽�.�$���ŋI��NMWs]a��KD�)�S̨�26�[2��a{��b4�n�ǩ�8�6A��WgwY��4@��A�ժl�3,v�ߎm�`X��/��؅ʴYŐ޽���Z�d�Z�]h�7En
�u)�?�;��0�R�JH�Z^ev��Bi%����.������jZ����ܶ��u`�"OF��'D��1�l��寅�u�PF��W6���D�ı��hص-�p�in�pb�IskP!6J�Z�	ҭu�J〨VR/	�@�ۡ+Q�5f�MRH`z)-"�e�u(TTl9�`�����2T�J�dra��o	wt��Ռ�B̗��r����&(w�%���P�0\VP�%���Z��qI70����@h�u�Em5cE�{�cl]�Ј�L4^����{u�Z��ڷ��"�V7���`ī>X�w�ZՅ8�Ӹ��Мە���@:�S�j藸Yy1�m袰+o&�7N���gYр�&��4������CA�GE���K�ی҂�~��f�(�>�wzV�h�%�U{���p����슝��z��Ŋ{Y>GC.ctѺQ�U�ƾWu�]E#�94n;1P՛v��ӫ.�ܙZ��ʰM�����V]4�I)÷.��]h+L�C�1V�e\B�I�t����Yp&���F�ڲ*��R�����JT�m@V��V+# `V|�R4sr�0섅2j�L�NӸ�x�P/2ej*�f9�[qk���X��b���1OU������X!�j�a���ek#�Z��DV�K/Z�%0��#7͗OU�WZ���s
X��ђ�i[R���Sm����.Z��1+"���X���H4*��r��D��cn�@k6�E� b�*X��A�����!f�N�+o6�6�(�#@����iT�KR��")m�Nl݊a�Šm[�&h-.�u޻W4�S,���lm!0���q�ѴY���ǭ���) �R�*�S{6/q���ˇie����f��t#.Bf���'�i�������(����ƶ+tstց�.�Tl"���#7M*�Ťe�֧������ {M�CKN��:	���4#-�D+46�fF� .-r�V^M��oQ��Q����D{��{[,[k��T�B�(�@qYD�v��ZU�1�e0ƺ�02�h]ʓJ�BZ�7�l;�-�������֔�Ŧ�v� ��xΪv�"�ɤ��1�+�T�6�ڳw�G�U��U\3�aF��V��U�Y�P
Ѽs+F�B��V�V�g����j��PQ&���PQj�)D�F��(VY����+O�w.�i)�3++�d�b���'a���p�*(��Qaˡ��C�5�t��:��-�kwQ"\�n�݊O'1�r�FU��5��v���+c���@@$��e��nG��V��lt>��r,2�'tu]�.ZTs
 ì(��ři֢.�`�JTͣ��l����.'XN0V�w[��.�� :j��$�OrJ$�bh��Sr�h��=��Z5;^�^�)k���X#��ݺޣ��*ý�Gs&3Ch�J
Q�F㖥l�)|�$3W�n��<r[��t	0�x�a)	�ٔ%���E�s)(�:���YpGX��?V��z4���zےZq`շ�i��kz	3\��_Ҵ22�:�ЧWJ�\���%Y�j�dY�&&Ž�؆�)�Ze�b�YWYA+0���^���J��L��S�j��b�xSz"9T�M	�&�fL?mcbʠ�d20b�����_3J^=��F��e�M�{�f�^M�뙴���!��:6n�P�d3ym�N��j�Q#x���Մ��J4�Q3j��^]�{����Į[F��S2�*+@�����9�֝ı�hf[�R"P[k���J� �Z����jVڔ�L�����[�����%�R"�A����R#3T��f���-��Y�Ly7yHb2�n�i�Z���*�/n��ٕ��7E���V|r*4cZ��tDb��Z�k-�&Y�y���9���EW�[����n٧Y[x��b˰�WJ��,�����R������v��[H�:1V;��s,��2H0J�oe�/
��m�,��d`�4C��խ�,d��Dk!�	��[�`�EJ&maC��R�:�d�b��A�U��O�:rK_Ϊ������T�ti��t�f�]4��VZ��ǆa��{hk�r��-Aջ��y�0Ս�����L�4k�uH��4݊ÓKq���*��K�kB�)ۍ�9����r��A+�_�����B���m�W���J"�`��G����'�c��nu���7mu3A]¹_o0��t�b�sN��V'a���m�[�>ە]�F�9֢��]mu�h�$^GX�C9��.��S�鄜Eѡ[7��7*n�L�[] ���v8��\�����\n�<�D�}�̫/������[{S�b�������ps�8Vf�ỵk/����(�ḺC��Y��ps��	"HL����K���zF��ŕ)K�.�E�N1���dބ�F����e���C�z���\��P��e�*<�덌9��tuY�5����zrs��V���r���UA	]j�fΫS�o>��i�r��N,W6��څ�&w��g)a��E>=1��Pu�BH�m:�/n�MA@=����Hk��c9B�������m�]�ecں!Ź�"kn�K��!����_=C�v��x�r��9�%3%��'�^�3��h���wdA�w,7�M��']�(N�u}C���/I�0^�7�=���Z���
��\@�A��O�*W�4j�d{K�ZxiLU��S�M�}��(ڣ�x�AF:���:]0�B�,�q��)a;�ܠ��aw<�b��;�ݦ+�s�mv�A��}&���VlU�������*�'q��ۖ뱙Ʀ1��\ښQS�XW�Sf�f�j��T����%on����I�p�Ԑ�kY�f� �(^к����xV��wG�Q!�(�F��L�/m*X�ī��r���IQ�,Ton�gb�{Nc�����#H��̫Uꆞ����X�T9�f+ݖ��|o�
;Yq�K�i��%l'��o�u����bҜ�Ll����鮑��0-jS�åEoU+�4�5d�]��y.��7݃O3�o_�Sp�y�]��K����y](srLu����M�6oe���&D��KU*�퉪�31ss/�U��u���_��]��x����[����̗WB���<xT���T��r�tQ��[��[�)|uR��Nvy�-�(�q7%�Æcn�hc���Q���[���Kb�}���M}�s�hp�cp��:*�E�!�v��s(:/h�Q�<�����׺��̂�2���J\�0��J�-��9���7�Y�'��1���J̇D�r���ю':v9����lᇢ��E�TC�X��M�[�Ϟ�6a0�3jKT:l�G�fV��3Jf�Q��I<Zf�b(���K��=�X�w�;��Ƅ���sx�Bc�W8#�� h�٨b���
�١�����
�oF� �F���vCVI�u�S)������v��°��+)�v��ӊ�XZB��WF���9ʱ,�����t�|���Z5^����K�u|:f�D#B[v���V�y��d��{[J��.K�'�$>5���@�\�v��]Ơ
�d��b���n,sI���i�Fjl쫻�\�]��f�n��)�K
C���s\��d{X6澕+�|�O3k��שЮw��*J?�.��h�rk5�GKT;+2��B�?m`'g�ee+�0�8��3�[���:;�s��6,G�x+���4�\� aƵ�;�5`v�ͫ��dX���$�6ѳś��w��W�;Ǡ�b]v�>�P�ד�:�m�6�-++4�s�u(���(W�zOc�!Y�Py����A��s�sTc"8�\�oU�aY,�4雺��P\����ga0)��V�;t�����1�A�L���)[�ݞ��QmN�j��2�a˫D���C4ZZ�)}�#?.�OD���
M�4�}m�Ɖ�6+�ےd&>@���n���ѐc;�>�q�nT�๷nŗ����h�Z��ib��zӒ����a�\�+���P����^��b��r��)�d�%Q�V]�1�&�;��-P����U���ɖn��ϹoU���E
=�q�rj�G˭VQc �G�o	@�kI�Z�E*�Γx�T=a%�P�z�:��`�6���P��}���� ��_�N"�){]�-���TK\��9۔��\;v+%�J��m�]��z���1���:�_qs��)wu�u7t�n�.��\�P�V��ˁ�-���e�T�BQ�����y��݆/��c��IRy���)���]7�3{k�w�p,��[C�u�].�d�2�S�KҜ��ښqg*�pE�ym��O�<����pc�73����+h:�����E�����V��1�r�ٽ-�=��[�Nn�ܕf@�-�=���Wظu�o��iե�����X��=�3��w1�v�4RX�u��Ӛ�0��ֆ*��B�si��dګ��1-ӵӸ!�b��*ŧ�i������E��k[��
�Fr�WVE6@�5c%fZ�Gv�v���-�Vs J�rv:�<��F)��l�U�;z�u�Vtg�����"j��C�^GN����K&h����\(_p�t���q,4g_,�',ffH:�#��a�J�V@�K�Z���*�N���9�E�'�N�rW�s��d���$<$;����W[}��|)�i�d�m��H/N؂�X��A��C����*�Xʎ���q�-�w,�U�H�>�����!����k��k�"݆����^t��w�}�w^jǇPgN�It{Τ8Z��u�wIb=��}��ڂ����fJ@�K�w\�����l�EQ�ɜX��6ֱf�5Wq[��Ճe��hN��:�݁�:�u�-���+N
U,������t.,��ݴ'Gl�"ʴ�7l�5�¥�L�u�w-��ؔ�V,�����t��Ү�X`u��}{>y��,���4���W' ��\�Z�#qVen��}Q-�Wn�,8�Eu�
�4��e���Zw��F���Yw�5 �2E� �1�i���Y�Fmp�6tCZ9(��J�z(��P�E�:���������C�MYX��S�wQ�ӪѮ�r�,�Y[ۭ��g�f�p4�FC(x8m:��ˬ���{��c���+i!��^v4��5����{j]�S�!t�ܲ��*Ӓ�^���f�W!�B��gȳW��v��ܮ�[�\���˱lo�<�{Rb.T�ˆ�R�C,����y��]c)�O&�m>���v�������v�.(q�;kit��k��ӳ��_r�hK�!r۴�c#f_���H��n���x5�,�G(�˱�Ѵ�	��-�G�,�m�0l���l��E�7��hCg)�{�&ng㮴�oG|Fs�Yʕ��A{�L�OY�].��]�՞�F�r���8�c��fJ���.Ʈ����ˢ��hX.�/Cԡ��u#�M�*T���Y�/�*�6���ʴ5:�\���>��.���4+EۃZ�*�6s����(s�Y�ɖa���������G��܇F���m��Ƽhr�sh��U�̭���ܸ�b�iBU��y�ʽ��2��/�0]�Ԩλ�m�E�IK'3�!���b���C4a��2�ga�i֥a�d�4��M*��#Sv��V�54E�<"���`8���s:gWJ\ڙ,r�Ȟ�v��� ��^�#��^�{j��odV)��h�\�
#9꧵.ewu<��t(�؀;m��D+B��r�̅0r��|J \c��^�s��������c)(�ںŉ��Q\�0V�Xk���@����x��1��ί0RR:����7�N��|V�7~D,���B	
]6�C��;���92u��"Kf`����Z��&���O��f���+��`�tm�� ����t���f�ܠ��yWq�Ղ�z�8d�km��l��B�G]1WY��i�':�d��tz<ʹ���vObÝ]{Z�.}�N�Qt&Z��u�8r���Sٝ�ޕ�&U����9�ߴ�v4H�Q��j�K��}[���#t�6]=.���]O�!����كs1˫{\z�B�^�+3Zg딀��սO�"`�]4s���I8dR��M�N������2���򋝺!f���޷��s�Y�@��iE�p��6m�txB
VNN��H�4і�w�|������h�����8��O0�sԫ�ȓӇ�}��Et�%:Ȯ�Q�պ��n���Cu�'S����ԽS"f�P�crT�C8���5�J4$�̜��x{�{jHN.�8��]����(�����Y��c�$
����P��5���+Y��w~�.C5��˂�e\�躱t���s]$�VsP��9�L�Ý��Rv�G��Gv�S��V��	!����TS"�7�V㫰R��W�.��M&���nn�(��-��iU�YuO�f4�0٢�{p�6���6�Ii_qw)}2C���O-#���޷+��f�����
�����b�X��RG.n�8�2�U���w+��ջcR5����y�VN�OU��k���{�X����s]s 'QSF�[`e[���j�r��H��{{Qh��p�fh)�����5v�<��]gc�3�������q�(}�7o�7X��}ȇ|�b勪GT5`�9n�N�c����)�X
V�s�����r16���oa�6��ٻ�����U�n�1�w]����c�6��qش8�71��L�*��U���c�n����˸�hqs�<�\�� ����dE>���m^*�����s"�q�y
Ǘw΍���i���(�"c��
n�d2����s�\�Z�-"���lh��R�i����a����1`q���r�I�p��t^d.���M1��;���e�ߡ5��u֟����N���!�]���e��vP`�����f��wG*�`Q	�����h�Y��Ջ�b>���8-q�F-�ܟ�~�O��U!��+K8���YŠ�`�l�L��&;�.�V������<gPi�<���]ً j�-yj�UǷ+�]}03����i����e�j6�-��v�Dygj�
�o �9G��ܭ��R�qI{r����;��N7YN�*"�c�+��Gs&lT��j�ʾ�����j��n�1Q���9g�/�������%+qY�,+ܬy͂���p�ۘ�<�����.���'b�}ǩ��u��I+��]x�YjZA��Z�S�k��h�p�)֎��rm���Mr��[+��l�������lR=C����ʻ�)Wp
����R�� �r%�t�_��U�F]͓��#s~�Xo�2a�R�+d�SG�yN��o�,�w��y#�4yAfsK;�4�����f�/��r��\6�.i_;ɗC�<�1��C(S(�Z��jfE�1N�T�_K��2ѻ�J���H�j��Hi������q��;�9�r�N���Kiv*�c	Mm���HK��䏵̗+̩���=��oV��en��N_mKZqe,���K��n!�]YF��y]�p�2ȭ���Ю<4�.�wm��u]��Ϥ��C@[����y+C���켆�
�������QÙE��vY�Tdܗ��&��h�[�&�=�w�V��o�'�����n=aøPa@��}Q�Y�+�ko���&������7�įEG���ĵq\0(�V�ѧ�����b��wT�M�V+���3*L�������m��.��=}�D6"�b�u�Y=�jiV��]�{�	bڬ�I;bC���t�G�79W*�H"M���
U����b��|T={��:�R|�~8���MF,+tѕv�f"X�s+9�5j�.��tm��<;�t�IU�^鐽wo���ٮ�.���Ѡ�Ϋ��k�*� ��N�AE.+(թVw��w*�GJ���B���v�a�e����v�I$v�ꄺFV�9Y�ϑ��+�k�[��ѓ_"�.��h���x#���B�ox]�i��ZT�%M3.�&���R�)i�=mc�Nl��
}v8p���V��%�e+�@`85��m��>0
Z-��n�if����dj 5Q�6��11|�#9!v�p�E�,��S�F�Tp,�q�yO���+��	��[M���w�LLf[q�Z�m_ۨ]>+�@��b�E�uy�7��%��T����R�>��2��Kp��3�M�[j�2,�IS�a��Lj�H�δ�u������Vt�QIf�M6�i���fR����;"�X��\9�%(�*��.L��Ѵ*��[z׬�ʲB��}�,�r��YwY����]S�>��@��`��깑
�ʕ��rN�:�0&�;Gund *�
��GA��H�(��j�d�����K���%Epɜ�N5��3��j�cj�2��k1Kc-�4K����Jtq���Vҽ�w|��譛�A�����n҃VX�(%8�찧T�x�b��8P�x�o��3�W%�+ۆ!v/����BJ�Y�K(A%sͻeZ��d�s��s�U4s�w>㡛:�n��$�{ XͳG���.��ķ����(*t샼��ٮ�1�d�u��0�҅��н질�8;i[�������wM`YU��QЯI�a����/h�pZ�QbV�"�1��.H@K���3]�@��\шg%�j�t͚w;O
h 2�|�мW���d� ������Y��]�N�e�����6&�#��m@8�ݝ���.>��d��D����w��������O4P +Z	�����x7�D�ȳ_S�Mu��E��՚�j��B�����6Bz�Lͷ��x�dٛ�,v�N��Yyڡ�zӂq������f�	b��Q}�x���Ә���:�~���N�:�v:���A6����]pʧ��]b��^1ѡ��ںƫ�V͕y�V:y%�,�a��u��g���N���%h͕����B�h��hul�lw���� �î�Z9>��Y��xL��y�yZԨ�Lq�(d�#��4�\���V�������=��x{����t���W��~���UU4�-\rh7@oCZ�2���� �TR�A�lǣ	�e�%@w֬��*%&��-��4C���dBM�_v>�o�r��y���d$#�;ט�m�$*�A�ێک�Es�7sk$H��ͬo1p�	��7��\�9�Գt�&���!bV��ٻ}
��a�����G1L9�v�}���K	�Ι�MK�mݙM��]�Ρ����M�w���\3���|�ؖ��l�nixDt]I�Ay�1l{��1Z���+js�#���uum)�Au�[�ݩ���ѓQ9|�ւOK��]�iv���Ry4>׆�/���kU�N��^�
��J+�r�ͅ�c��L����	;��"�Y}[��0��j�藖����� ���R��X��P?e��V��ˊ�$*G($��2��c��u��^n�R��<,V:yq�w�R�]���6����m�2F�B�eiޜ�
OM^�������G3�ntާ�FҬ��bƜ4B/N�Yʬ�c�:]A���#$_H��s���0�@�rk�4�*m:����a�C����sҫ!� FEJj��·9>�dI���Y{��D�|��DU��)
=[����g���}H�S�9�:�Ƿt{x�c��ښ^V����S���r��
ȑ�����J��
�Z��\kp��-��:�;�6�v�;sk�kU4�b��4B����(�����Y��RŜ�x��+����]:e�[Z$tS��u֚en,hr�T�х��9�J�����Q����u�ŒO��`9���zH.��ך���Th�5s:��̔��
�u��l�W�6�,�+�!���e�OK�2�]]L��.����0Ƴ;*-����I�^p2H�Y���^�uj��$I��}���\��:YT{^�[F�ngl��]hb��)N�aj��b�t�o>QT��"�H;v�&�p@�rX|"�Rv����ZE�aȩ�ĝ�2(��\�'U��h��s[A�t{]ٍ�ѣ'm7B"M�)���w��uCh���,]��b�xt���u��5loS��Xҩ���G��D��'p�Y(ɷB.�ѣa\���c(G����l9����Z�.�vS��0gm�R{p��q�W'8�nBy��-����p��Ŏ6���w�i=�Bؠ�V�1�Ԩ�u��u�(�ĩk�+e�<;�,wl��!�:�sRW,�O����B]��Yv�X��^����t��'��Eleo'	�V�����m��N�I��V�I��Ϸ ����ҏ#A�
h���_PQ�b�<s�q�|��Z엔$��<@�
aSZ&���
�ť;��Z䢹�V�fq���(@o2��y�\�}�c��{�eG������H�I�w<�#iѭ��2�+�3ԉH�7.�:|���˛��N�⾡]N���c��oEΏ^J��Nqd��xR�ж����)x;v�F>�x*�ᇙ�M1�u�S�7�G��kӧ�����1}L�K��5�YGk�;-:#������4
�﷫���WMR��ȡ�
���em^J�섮���{Hr��&��]l;�&Χ|�H��"h�ee]�]��[��܌f|�ܐ*�|��4݈s���I] �V�.��$.7ƺ1�r�}��5���9ZH��@��2t˭\k�.h/K�a�=Cy��wh��W�����@��}���(�����gT�-E|Yi���{Ż���{۸
��	�D��;��fm�ԡ��j���YiJI�칑��˼�7�6�aλN%\¾b%G��M-[�X���J�������rm�n���M��˭���$ػ�~EhЯlֲ͝��_]�����JUXk���*BL��|�N���p��o]^��&�|w�r;� %�c{9�o6����Wbc&��x�${-�.��;o��{�=έ�O
]�o!6�/����^f��w���QH��t�9�4.�1_�����QVoPYdm��*�l���I�8�v��o7�i}��U����V�"C�^��L!�.��2v����,,q��6Y���u����oEX�	�u���۪A��৓ud�o��N)dy��2�ද
�j:R�/y��˻7��G ��і�dMU���Dv
�*�G�
X,ଆ�R[8�,��8��0-���܄��w�f�k
�B)l��E�fJ����M�nw+�|і���Q���W[+f݉�vAX�2M-A$[q�qD�ռƯ����uc	=O3�EHކM�랽�<(���7��1vsII{�m���;2�-S9ju_B5u}��L=��=�YHaS`4o%.�D:t�����N�c,�R#cZ�"�6݋h���waMn��4�!C��ʻp��5�ڊ��iVg�p��L������ ��r�3�ھ�JvL�f�P�z�S<�d���#���e�0szYUɝ��82^���z���]p�q�H<�N��G���\�ل�	"ޜOxg<�;v��i����M���.a�E뤆G��=�c�?1�  �!�z�g^�O�!*&�㛛J�!czi�E�^�ә.�iQG��zk6�n!����v�(]#��P���[��@fR5����X�I���]��.��GNY���9j����\�u�v��(�Λ�8ZXb0�j�tR�Ev�kd={Ǒ�v����WBv`�I��6���+2S�6�3@��g�k������HR�M�L�Z��r���f���ZM']��]�����W��r
ܔtΦ�4��t�frt����)=q�u7��!\����b�V4X+�97b�K�]um�d�jk�n�Qv�oer0��b�����n�N�3yc
�:o��@֚�l]MK���Wm\	ͣW+2v^��f˟_7y�e�j������vG��R��Ĉ�mm��=�;�����Ch�E�,��L��!�wT��M�g;������n!i�=�ցc�1[|5�{j��ʽ%��tv���s��{�Xv�4��=�r�6t�{X!��L	+����U��~��٬���mh����.۱ϝ<�0LH�.�$eL[8��
�o4�W,��[�;'U�M6]]�B[&MaѢ+�������+��X��������fG� �/7>C��)w!�3��
ZC���:�٣�aΩ�>u}���Z���`�vs����7��b� ���
��F��˺X����sq^Z^����t7��%�m�`}��N�4_*�姇]t�w̷��1�tx���pEX��ZeLdCt#ȃo��Wf�ø�z��n�;�u����$9��[���f��ʥ�Y/Nv�}�`�SfV���+x� v�6�����k-r)-3#Q����`#��d�vBN�z�j�H��p��X�;V�Nłuu6�cit~9����u�Cr\
�r�҅]�5t3��)N�n���!��G��I-p��ҷ�%�e/�Χ�@
���J�'�dNǛ�VӢ�h㵌.U�Q���x��]�����e��p�'Y����;P��S1��2Wwp">����qXbV��0��t��.��Ou�C�����\-�=0]tyw�����{o�����o�������M_P�eA�ૺွ��7�qp9u�U7�\A�?7���sE�S1��m'�g|��v] �s}{��[�f�N���W��2���@h�`��;pWI@Zpм�I�����Q<�œv�҈���i���^P���֖�܏7��7	R� �
(OR���<�V@�KV w�������w��ϠV�$����=�G)�{����1k��ڭ�Dn���� ������+魪ol�+��v{J�)�mbԡ��2�lqi}�ݔ�Nnf�k�-;��:3����Y�0�P� �D˥(�7������e�_.�T�C
9!oKJ�+��QR��}u]���q\�Xݛ]��+�Xl�pU�:lzZ�X�e�][�J[�f�3R��@�Գ"C{8t�e���c2Rn�����
7�Qp�M�a���ƻ�5GЫz��܉���\lvqNm�$v����뭆�](�d�L<8O�M*�Aɳ�	�j�n��-�����,�*u;}a��s�:&�2E�6�>�RPΆ�,��򕷔+r.烎:����%��e`z�|�r=��t��[�ZÕ��RyGR�rsʻ`�&�p��v����-N��ʱ�+���}WWQ��O���uŔΰz�_�ؓ�w`�i;��v1�[�\ɥ��G�ܬ5�XK;�;we�x�qjuGg�NR�qi�ެ��4�{OS
n�����7!�)a�|ŭ�|{F�\Y=T+X��k�}���nA�I��T� �qᲝ���&�˔�B�m�N��F%o����Ae��Wg����)���/���
��4�����)�B��W�p(�]��u͡M+�z��u�1]5��Q�����ͺ�ݽ����lGP� �ckjt�
�+�U����BP�I�����U��1tt����Esi��E}ѽg�������}]�j���i[|�C\����Һ34�w���^rͬ�o]�s$��N^����b<�zim�+�$���R�����콹�$��g����[4	�0��u٣^��v��R�2�Y#��C��wE����F��KNP�ы�Wb�Ȼ����䘥������Y�����/�A1ƹ��ƻ	�+�K��h��حI�ШԐx6�*.��ł8��GKwvՠ):(S�Hv��>��T����jf��(#rU����\��n�b�@�א�ʱ�/*�M�vu:}FZ<�W	�i���ھ7S��J�#x�F��>n��'����c��Vfa�ySO<��(6�����K��M��[�+�d$ц�Xw�%�qN4�9���N3Hw���Y*61�*sL͎�@��H�}�~�F�}�O��������R`UΛ9��1�ld|���Y
E}Vl�t�$�m��`�1�T���Ա��7=�"��{��-�Kj���㹣;�պok*�Y��ww05�o�]���K˩�_f1�l�Y�f�&�]Oy�a�%f]\��'u�Ѻ�T�Y�B��U)q�daH����R������9h�rQH�0�WX6���4�r#�.yh{@SZ`�������ki��+2hn�e]��Z.[��BV�Q,r����������W���b�L/z����O��Q�^���ic�����t�uM��s�h=�şs�qz^ͬ��|�����.U�k�W5�j�T���υ]dݬ|����;��G7��
��^ۼ��@�)��±�Ug�*b��4�T�Qk*-R��8#r5�=Wbъ93�U��f#�>t����y�r�G+��
�w׏����'��/3�ut[L�)�I�	Ԑ�}Hv0OjK@֎]�t*�)�����t&fپ`�2�S�M��¸˦�,es����unұR�� Mv�N]t�J�E�����)�*��0)v*)d�������UnCpT�+73�5�8�Z�<����o[�vonY�;�[�Kx�1j��l<X�V�F��1�6�n�p��܋�=T�*9���dg:��"���6Hv�SNA���AK�I�ɵ|��U׻�S�4.����һ���Ev�Н��t�R�6�*G�jK%���N�0S�x��n����L)�Zxs�y�Y��L��g>���C`���u2�_H�=�N�����%�jN'�.�P��&+���+z��� ��i��ץp�Yn� �9��.���yUb�X��p���]�J�}��fܓ�2`�Ւd�W���;�n�ѼvA-쇹�P���Mw�IȬ�'��u����݂��vZ�BkLH�@��;�ll�ZGP�(_]�ϭ����We��q8-b��^]ӪB���*�7��L�7�,���������.转�����,a]`M�]	�9�K�Y���Z���[��)�vjy:Z�� x��{��^��I6��}9��s�H�ҺJ|��R�*�%�
�@.m���8f�2�Ng$%��4N:���V���9�k5�`!������$�bZ���s�4坽��kku�� ����H�/�F_U�>�c��w3��>�Z �Q��v��nS�˨��om+H%C9evZgi��*��.�����BλZ�)��������gWj��v�KR,��;t�������}[�*s��=+C��!�TN��/W$M_7�M$�[ݸyUՌ�i1x�@q%:�L�M�L|�e3T��s�ׯ�DL������b҈��[X(f�5�V�)Vok��`�8�]���oYE�j��f\z��L� =��FqA�zS�4g�p8a:�mm�V�-���f��78�Ӱ`���#-������*�)|��z��(�XP�V֧��w�7\���}P]�U�����'��\i�4�WZs9�S�B҂�m���17iʵ[�[��Q�W�@�-�+)�"�I�Ԝ:���;4G��i�\��	I�Ec[�Uτ��.v��<+iWq��-��>�رݒL,^�J�E%(q�w��=w�ru��ʧ���[�l��G�c�h>IV=F�m��\jo�k9�
�d���J�U㬻#mPcS
�Է�7JS�ʶ�:�������	8�g{�d׏�w�����3���{b�5Hڛ�-�����C������;���o���6���P�p����3;@ �>g�MU�۹΁�];[rv�i�].����8���˝�����ö��U͆w�2@�`i�M^&��:��;/I��-݇r�;S�>��q�j�
�]a[�-
�)a�bV-h��K`�匁ݹ������xx{��3u*.2�/#�L¬11<�,���wU�n��c�Ŋ���4[�8���r�y�m����l�([`\O1<�r�]ꅘ���]�hXܬ�h0q\��ےR)��2b�M{���4{]�3�N\{��w"ڶ3��=}t
#2b�p�d�s�]�[贺ʺ.���޾+��Ǩ��2L<9nwv���c��֣z(�W'df[�lCaɑ+i]���h�u�\\�<����F�.ess��s�놛�3��:�v�{�j��}��_:}i -�MQ]����	�}*V�� Mh]���;8K35���1訬��ݺ�����j�`����櫸���TJ���tk:�[�i���X�=<�ؖ���3���"���S<ʬں��&ze=�c�@��ٚ`�!�
����ٕ��v�]t�}/q�(i�����_f��z��r��;��	�-O�c�����y:�Na�����|{X��IO;�}��D���.�ޞ��Z��\��f���K�6oG,��)Ws�T�k����̧��َ�=��]���fgkXʠ7���Y�N4�ҚnQ�������l��{wh���s��R��f��ߛ8����v(��km[N�qQd�8P�	w�� ����\���i��i�m�;x�.�ް�]�����;	'V.�Y��@Gh�CE"3�}�^�T���ǮAI`K��M_(�&efs��ᄕd*���1��N��Ӕ��(Ru��+w%k�;+s!i+2��������D�"$�je0�r�������k�D��L��iB��3��[h��\��j�[l��*ֶ�ժԬA)\�#��[Ymm
5���h�E��l�)e2ʙZ��+Z��J6�*��*����m("�Y��QJYmR�mR�Th�A��	Z��V4��B��#Vд�h�ee)m�����EPm�S\(T3.��#Z4e�h��R�Y��TV�UF(��U�JյTe[A�Z�ʶ�j,�F6��J�jV�8(�ZS-h�ڥlX�-�eF����V�J�i��r҈6Զ���ʭk��K�����D�T��+m���j�ZYk�k*�*�i��DKl�j)LqQ1�X���Z��jPZ��T��5�Z"%h��m��m�R�*6ѵ�KZX�,S.L��ޗ����PD�[wˠ�'��0"�庑���wnG��=Z�w��=h	�vN�	�V�����$��6��8��=�0��8����u�N}�;m��Q�L�V�*��}qcnh7�U�5Ev��7m*ө�ۘj��V�Պ}P(rq =��V��m�V��]<���k'��2S����i�;�J׾SM%9[M����̻ݢ���^"rou/e�e�eQ�>�8��x]��-�q8)7�%r���Ʋ�3˵泥#�/������8�\���u�0d�Ƹ:��0[��%�+��x�x�>�drB$!GA�W�lʸ�j�X��@�ػ��g$����aڵ=ol\,k��5�m:��۰�P��V�{%'ޱ6��B�i��r�9��Q@$��F�hk<ݸ�3]Põla[X��˞�;|��v��Rݎ������o+�u�[s`s�(a�U��ڄ�n7������,�r��4+53Jܴ�/ΰ�7g��:��������Ẑ�:�]v���>��ҭG3G��w]�s��������!�º�#M�����h��0/���W��xM��R�27<3����:7��I�-o`[�f�`}V%��0Ս�ﰡ�Q�VN���JkmQ��1��KC㭛1խއ�.�Ǻ593�Ci���65"�;j���_o,7y��I��kkV�ܯR[I����o��4��&z�#"��#���q�k�a+��#_m�}����K+�Eann��C�z���qX����̥~�b��������гz�t� �S^a���'R�p�e
�ww[)n�W<��b+-�u�-���a�;��C��A�ʆ�����Q�kK׊.��W&�\�OVW�<�S� $�h;ꝲ�s��QՙA��b�q�ܒ�F�����o����:[�%�����F��`�냶��[��ܨmdO���a�>Kg<��N�OU��x�ǽ���D}�5M��zX��Z,[|�ĩ3�
gK�<nD���"��c��R�,n'�k��zc=��pJ�,N��8�'ڍ_yMYO�������L%���M7�z�:�ǴGK�|�:��s�&���3kF�R�<��X��ؠ��,Ԓw�j�H�LE��5H��R���rr�
�r�M/)�����*FK@b�e�A�v�4;:-�Ӄ���rN����ep��ݬ]?-�MY)"efWD󞸷3�ƣ��]J�Waw��N~��y5���[��|���q+�t�1}�f<��@���q�S9�7������_e�6+.�BZ��wv��g�϶��x�Yղ���OF�sX3P�*��1�.Z]ܳ61�������&�P�n�\�C-�]��k��,zl��3�b̙�[E5�^��I�i�N��h5�SȎ���uj=�ڇ�byº������S<�V�K����ͧ���d���sbrg��U���idFL���Z�Ư-"�׹T秢�پQ�5[]�?�Lʭ�{Ya+�)��D}؝/wX�._%0���i=y�]^�VT>��e����wfH�:�.��g����*eoz�H�+k�Y��S�����^Re��=�V��������n�k��C�%ڴ��ar\��{K��417��S���w��ˆ7N:��xI��l��]=@C�Bg��(k��J{zϽ5���N��˛W�79g3����Luu["�'��ER��)F^D��'���e;�X��=�W�J�Kwr�d�E�I(֙��]X�����tu���������p����+wz�;�y���~J΋�fEP+i����T�t:�^!������X����WcnC�YV)u@��=#ʫ����j��ݿu4-Ÿ�b�LR>G���])�I*�bS��D�qN�\V�r��؛n4��y�{��˶<��}V#b��#��D�h�TO�e�-{�}���[��R'8���a�B3We^J�s�d��aR���p]����q��@)��DW�n��<#��2�y���&������	���s��r:9p+9���~ܸ27���!��9����JɧN�\�C-��+�F>H.<�sS=�����j��{�rK?U�\@���>�������l�pu/$��䦵ڃ	b�b�򘰱��O�/�r1��+��a�o�"f	���˴�f1���p�f�k�[�ֽ�n���N��������+�/n��\�,lJp��;	+m��rmt�Uۯ�́h��]�։�i>���IP�@e�;h�'���#��*Gxs����P�)���C:�F����9��{���E:��wucC]6-T��=ϖ����T�OP�Cxm��l9{�u�e�|� �kC�ZgGmr��}���vk��5�y[��j%��~H�*�"ޭ�I�Ď�i۰�|��\)��v\���U��71�fk��2���l�|��=^�\z�)���d��F�䎃�=8�gq���7c�hڍ��V�t�s˶e>wTΫ}��sf&7�u���y��a�P�t,! =�}g
��0��T�rV�n�{�g�M�wx=��k�����c��,�c��yX�,t�e�������:���̪<���_��סk���$�j�'P(*Qm:&�F%י7��y��/���}`Kʢ��U��wyN��T<�lWG�s26��`�ܝJ�*�b'�9�뼞;FU�,�R�0C�zy���P�9&��7w�.�Y�.Wb��6�މ�̹CQ��|��y���O��9��$����mV����(���}�W������c�`�,�s�\�-��]+���Y-Z�L�g������>�[}]b5/���1�p�F�q���Wp}�Y��pf�o�YkoV�5�e���"he�z�!<�M�ws�wR��#�+�M�����	<�uy��14�-�<�����{��Dm��R��*���&�|�&W���9�y����_:�'��F�u���"y��ٚz���������Ջĭ�����?��bڣ����[P��������U�(�K���l�=�4<�ʥiS�[���\�BƦd.m9���uQv�f����:��3W�p�� j�n����S�	��ԏ����]�9S]]y3��wiVnְ����Y���@C�ɰ'�E!�WC��R���=^�˅��3su̸���}�����a��V2���!�U����2���{�(���:�t>�|�s���r�y_���+tJ�\	B�9Gk���C�]����%;�=�ێ�$T��t1vr���yy��VwbC��8�%-AW�t���Xgֲ�.���T:�~ո����ua�T�H�[��M��MO#�/^�����L�L���1�N�U�b*Y�[���KFl\p<x�]n[�^q���w�bZ�chO�u�k�,�E.<�B�r�*����nś���0�ӮeY����EbV�&u��5����Q�:ҩg�i����VL[��2���;���j5����Jq�n��A#$ݣ���]�#���kps�q�=R]{:;�P���@�T�o�J�}��C�#;q�lܞ�+��ۨ���w�r��
��V8��g�-r�{@��f�t��vb�\5j�8�)����*q*L��t�|�g��p�J7^���ޅd����;n�;U�P��Wڥ��m�P�\�F���.�`�7���\�jK��G�ٺT��&L�*)�Ѹ3�ą9U];N���Ŵ�!��5�g1�����u9�[��(P�q���h��O���V�����5c�%}�YS�-��=~rP�>/�
�s����['�%C+���3͉�߾q%������o&����������~�/�4ܬ۷U�Õs��j��Q��k���=��#/u�V����Qu {��qm.+_�_^�v���n_k�n����6)de/	l�]�KV���Z^��uG��na}��>��Bم������x>չ��BF�9�ϲ��w�oI��Xr�k�M*�)ͨ�.�A��<�2M����Q0e��,��̓�4�erV-��èe$k]%�c�����~K7��Ǵ%�^x�N��ѯ.6e=皷�t��l�H���˄-�j�;���>���J��~J�%���D/�:��\Uv�%]�A�oylc�����2�8홹�̼�<��F����P�`�u�ޭZ��T�s�u?��Zq�\YN�^2\�r-���u��!O�â\>�~+*�*�jni�څ�;���+)^.��}���;��x�٪j�W5fC���l��N��ٕ��U���ǎ��-(�ci:ǛP��SM%84J{�(�̺������AD;iU(��W�o\��>~�P;Ρ����qI3���h��)��vw/��}���XZmv�U�v���FBW۰ur��]�����«���}�4���'����3���m˸�[k*Ѣ���M]y��^[���$ ��.�]�`�},��Y�lm�-5��D3{b��vKU|��26���R�if����J�ϡ�s��҇��<q2�k����{����u�v�pF�A���)u�����NCW]k�fc�����,'�j���-��%[d߻�!snx�J������˭�{Y�Bb�������ՎnwjiUQ{KC��1i=4�fN�uq'�?yǔV7.��/G9t������^�C�S�r�NsgMN��(�֙�]�nf��w�o�Ԑ��{մ�#C7����=��k"ě�͚�:^��[�p�?Fud��ϩ�LubfG�Z4#��m.�;ړ�Z��C�6�o��-�fC=�w�DL5�#��z;�H�'n�)\��\ڶ�R�	c�k��=��4�C�P�six��[�jy.$�et�m�y�)�*|�'~;�P��N�r�
�x;�:�1NT���[:�v���Ꝼ+�K���W�m�<<V�&X�ϰ��=«���qk�kr�4i۞���O^�'{~	V�תm![�?����{�M�ۇ���tǯ�-�!m�Pc˕%�)��K?0v�ӎr���yzof-��b���9����],�=����r�>�N�M1�^q�ys��4�|1�;�eǛ��ތ5���d��)��5�,��O&��ð�/gc��{�٥�Q�8�����]����C�ђ��T�%YV):�'��e% �5˔,�|�se�Ӿ8X�ڭw��δ�U��x9�듦�-���mɍ|\�<�T�r��D�2�s7��O�W��Ҽ�q�g���Vh��GaT�a}��k�	H��dO�T�E_R�y�y1Y��*8)W"�5�}�F��p4��js�<������ҧQv���ǟ���vK�R��y���Qz�+y�6]�k'm��������Z9p]9j�;ʛYq���e�:��V�kv�$+�B�_.���-U��c8����us�>���xм�ʦӔ1%��ptn�U9w�s��{�7i���bޫ��>�6E4&�3Y�칅�����ɸ���T�/\c���^v�K535���nzi�L��'']7�Vp%u�9m�T��rD���P"����\�Z�X���H3W���GB�f�uI2K,��'B�!j�r�dZ��DRr��DB������I�aM���Z��uGo@ɼ���*/��{\8��r��W���g�^�oNG��m��	jE׽A2�~2��i�<b�'��:�U�^p��_J�qa۬U����a�Y���>X�R���-"��V�09k�;�-�`��;��-=b�{pt݂�
�b�϶Y��vV]3��WBu���S�Έ����g:��P󎬎iĵb��b��|j�����4�����l���՛���F�˩k8c�M��e>\^Ϣy�]w��:�A�,[�X[+��N]ф��0�Vwe&б�m���4o;/���b��m%J�n�{9�X������1{.2���h:�p�sk�g�jG8�gj#�Hw���R}4�gv;��U��k�ˎ:=]�>�ٗ���b�E�	��/%��v�}���͋��x�d\U�ɡ���Y�/Ү"�諐�9�27�rv�ݹ�j����>~V�M��V{xr㵋�}�e�%S�;g`C:��]�扗B��P��8~X/w��<����P�	��tF��`s咹2�H�wq=��V�x9ip�n��m xNo2�i���J&�7�^�����.ڒ�	��(u2�<�w+��.�Z/M9Wa�9���š�Q��I��Ce'�A|���o��F*ɂ�f4j�����+e�ۡ�c�-_cw�+i��d[f`a-�CO]Q�q���b�3�7~��'�Kpl���e�G��*`���,Iͣ\uō٤$/t�t�c�۽mU�FKk���v�|tw;��՜@�*���3ZT��v�b��s��X�UӜ]�_S���*=�*��Q=�R�z�Y����}�Y4ӼߙyA-�%7���o��&J�^m���&h��\���i'l�	����32)����ݣ��_075������f��H]6���iw>��ò�+�n��%���wU�KR��Za���z��^}}��+/B���fem���'XN�V-�j,���n��8�$1�+���,�j���H0o�֒ЄQKcr��Fh!��-�Bl�����˛W%�f�7[�ҭly�R�66U��u?��t�e\?P&�H�����w#��n�]X�VVkۛ ��<	!�M�vEyY�/c�lё��T�b'�%��0;�Y���W�wuhr,�O�@b�n�JJ6]�C'�U�7n�'��m䆄�VD�'�9 �+T���f�ϥA�k�̬����JGc�c�L��C�(ݐ��Q�fX!x��#)�k N�&@<���f(C�3��Yi�R۩C.AB�b�QV��=�*��V\�m�� Y�vf�7R��VAV.�Đ�E�4T))�����$�S��y+�v�6�����}�x>VV�Ki]9ʥ*֢��K,�m�R���h���kEm�\n6شe-��V�8##
,R#iDh��ŨVڵ1+��*��YAq�L�d��2�U�����Y�-��L�1em�\�CU���m�TeV���2�ƭk���VE�mA��[QE��ҴAKj[X�(�DYXT�ijQX�U�m���J�V(�DV�D2���������h�e�Dj���,m)DYQmmE�����,W)G�Vڍ�ƶ��Q*rʹhĴ��j�J�jڢ[QKJ�-*�*����ʪ�KYr�Wn[ �p[���X�+m"�U*E*[k*-j�hR�jԶ������E�h��j���V�mH�-���("��*��(�[cV���F���8�L^�{�~;t-�M�ԅoi��3�༌צP��^���q[����mv]S��{%�R�o3M��g��ɋM'!\ܣ��t�Ż�N��.�i��g��
����_}��-�r�/���Kŕ'�{~�͙�7�[�����=[�3r���U9�Î��*	��M�U��`g)�-�피{�S/��OD�Z�)�>�9Vk�WJ�751�aºQ��Hg[�K:�!=�����E��	R�ll�.����.��/f�U�yX����l.0�u}I��"n{���罍����Wy>�~��dwMaӎ_a���R+i����-���Rzd�WǗS�ާẫj됨	L�=c�/�\���rz/�<S+efރ�+�+�Uy���]�����h�K��8��}���Z�W����h�j��k7!S+p8����y��s��Q���k�r��8P�$�ߜ�Ҩ���S}.�ic��X;4��	�(
���Źojq.�y��긍��Q.��6��(W����.O�D����T�s���%z��u��[GpYx�  ��cOj� ����R�q��#�;�V ��<5�3�=G-6������	z��k�|�`����k���Odohs������1��.��N����k&)�@Du剥�uMظBE�c�W�Mf����zu��9�	ͥ�g��v�Q�S�����"a�9:���G���ZE��n�k��v��{^�Lz�u��rg�;q��T�z_j��ىf�2q#{���������g�vMRQ����C�ɂۙ�͑��J�g/�T�ϫ��H�]��·�������+�tS�JL�ܳ���U�^��A�l�I�щK�yN���a���Ӟc����r�)�Α��+��s�!qT;T1s��=Js��ޕ�w��i��u��³��yP�xO�.�g�tu\��p�͡h�y*��MOFv���n�X<�^�����l��<�N����%�n�r�oV[Yz�Rp�턱�s���R�'0���8_��,�75 ��W��mkmm��0SN�M���yO.��{�J._�,")LoX�"���]b��ʝ�]���,�]eW[����as�{_�#�"�^U_IC��x��S$���Y��$����ߚީ����X#�Y�0�l.w�b�ܸwQRT�WX��w3�������;W�cΚz�NO`O�(�&e!ڪk�,�к]�����<TqY�ʣq����F�Yc�ߜN
=�o3U鬥5�1���ۑ�c�z�tf�wb�^J��������>,�L��<��};���������W�lK���U�-�(Qy|�f�7@���.�s��{U��A�`�Y��/:���O���{*�RU���Χ]�ؔb��Y���7A'�������鞴�v���8���=��6��Χ{<+-�C�Hʡc���v��1^Bjp�|���ѩ�~N�_C�0��9ّ\��r��xدf�k�[|��sپ\�纐����r�vk���~���^���S����?$����'a>t2q����R~d�'->d8��_��u������`j���R��+r����t?!�=d;?}�2���׽�6�~g����i!�w!��m2��0<=�
I�'��v�'��'9lP��4�2��o3�ק�^�������Gov�ο��uI�����x����t��˦J+U(!c.`ck�\�Y�:�e�y"z�g{R�V�v���00�9�Xy׉�����Cy|���%g.1t�dN�U��r��(l��jƕ���'Q���3��s{DBW��>��z}��Ï���u3�C��a8��ҡ�I���Y8�2g�u�ԛE�H|��O;�=�@��y#�F��SJ��=�l8�ڼ浟k�����O��D>`q'����
�u?�<I:�S���3�O�~��0�>��Jΰ�C����P��I�M��Y@��5��3�w�t]kY����I���!��I�k�'�=x���2q&��5ϲd:�N����l�S��:����]�y	�<I��O��@����D��;G�}�[]����~�u�x��MZKh@���a8��~�z�a8�<�~CL�����C�i�'ܰ��!�OY���~C�L �w�@��zH��{>��߄��U�Ǽ��ʊI�;��@�i'��3�2n�5i:��O_K�q���l�bN��6��gO�:���P�$���Y������9��_$4���'X���_�̞��Y���i1�����g�I�X����8�����&���&�=}.w��d>C�m���t� i��"O���!|}��X�53�ff~�4ΰ�'�1�H�;?}��M��Y�)�c���q��w%a��I���$��OO)8��1�C��N2� ��>�2<{lG�^��}�w��C��M��'�;�̇U�u=9�u��X��l�hy>�Hu�s)r�u�S���Xi?0���z�>��}��	>;v�a�5���9gn�W��y��8ɦm�z�d�/��E'S�XuY'a�s��'�Bq�@��-�܀�VL�w6�I�O~�+��D��	����v�3c1$����`c0�a�߰������C�N3�5�ɶOu��H��f��w�$�s�I����%@�'�~퀰(�������.�ĕ44�r�d���W�<��ڼ!��'�9ф��쪳q�q��x4���_G�ӕě4$�ёu��>�y�o<x&�~xF���i&�hǆ.���N�u��]�c�*�M^�}����렼��փ{:��P�\�J��rI�~��U1��_�&��	�Y�hi�dמ��$�e������<`qOu�i:���'�L��{d��No!�<@�j)O�_D}?FEʨ��[�^W��OϨ~`i!Y���
��>���&��1	�1�g���I��̓��<����E��t��q��N0���n��j��u��B��U�K�����|t>�C�O�������k��?2����%d+5��|ɦx��,����s�$��ӶN"�`{�'�<�������o�K�ǰ����?Y�?3�fޤ�C����&��!����C�?3�s�&�O�㥁�Hy3�����<C2bM���~O���.M��j7���{�ﾀ}���UA��N[�R~@������C��s&��:�S��u��!��Τ?!�����p��$�=3�+'���ܝI�&�O�CS�;3�j�ﮯr����>��>�����$�O�2q��C�$��~7d8��yy�?3�'6�P���<g�~Cx}�*I�}c+�[v�>�';{&�{{��τ�z�Bt-�I��H��(@���s$�2o;�}l'��|����t8��gɮ}�+!������I�M�'X~g���:3��J���W�k��>��{�@����TY'P�~���Y%�'|ɻdԴ i��~��N0/i<~I8�yd�����q�Ԛg��ԅa7�>3â�|x���6�O۹��#�@� ��s�8��=g	�+'�¢�8�7J��a7�0��6Ԛ-�a�?XN06{�	��'P���4���$w���1RI�b�O�*߬�@��3�i�d�;��C�O��^�!Ԟ�b,��!�LC��E��M�m��$�=� ~a�MY8��O_or�+{�����y��;?�t�.K?u�$���e�&(`���AZ�{��+8ʻp���i�|�:t���^d����g{ I>�������{���-�sټ��!e��Z;���G���T��K������QPe:�;�*���_8g��vw�L�������kz���Wi'�w���m�d�o��I�V~�P�I<��|���T�ré6Ɉ��}�C���N0�����x{�²|>F��^>��u�o��{�����m�I1��	���{�Y�C�{7`,���n��m
��`qI�ә��&�`{;̇R~d�a��C�	 S��Tx{��e:�U�rU����U�G`�z�v�G�������#�$q������=��!��Rx�l� ���O9z�VJ��}�uI�{�u��d;�Ԙ�=��]������z�=@����x�c'�(�����[`~C�m�~Xu!�1��rOY�bi�2u�I�O�1����$�N�����|=_@OQ����yN�~׻��·̚�C��*�i�ܰJɲ}�ӌ'Y=�d��?!:���!�ly�N2M���:�P����x��@4��G�>����������5��y���%@�;����LC��߼2}l��)���i<C��r��i��0�J���rM��!��e���l��gY=�����{���FB}�S�ݯ���7���<����08�'A�I>d�i����ῲ��m�?P�M?������O�s�'�C����J���0>a�M!�5�	�<d��_]�O_o�?s����'���|�I��~d�=���Ì5=�	���~��:�~a��p:�O�M}�d8�ϩ7�l�_� ��|��%���k�}_Ͼӵ�7��̛g�x��(�O�7�p�E���ݓ���������x͌��&�^��a��é8�!4w��xq���C}11[_c{��-Y�f}+=d�N��?!�����zɵa�e!�M2x����y�v�'۲q�����Hq����Y�g����<��}�}G�>��8m�Z`̭M��[qNX��x��'#cD�j8r����˖��nS�Y}՛��¥�r�� p�"���������X;L���WB*�;B��-��+hJ6f��o�h�ɼ8S,`�zZ�_'ҳ�{Se�V�Gˢ.��q�A^��U&o��H}g���T'x������$�5�Y>E	��'R~d�Rh2��0<�:�$��Y>���t�I�����'��w�>��~w�w�<���zΟ��'r�:�I1?��$��0���+>a:��ܕ'ȡ</�8��M�&��qI<=SD{Ȁ,O��d#��}w\;]g>ن�ŉnf.`i ag�}��}��O�5ϰ�Hm�C���Xg�9ܓ�=d�u/��1����E�q�N�����"��Om�e�q�_y��}���i��쯶��ڿ��'�T�AG��}�'�~`Vq�Ԟ�i��d6βOy߯��'�=@��N0���	�1��`A�y��>�}���	畿S�u���o����M�j�;i6��S����`{��fМC��Cl�������d=gY'����'�R<�C�?2b)��p'c?>p7�+�����͚Y��y�����،����Y^1�'��'a�z]�̇���I8��z��Rz�c�I�*~�����s>G��G���7w-L�����z���e��C��y���:��}�+'N�����d��04���N$=�
βx�$�J��pt||=z����z$b���6#~Z~]Y�o��I����m&�H{ϲT�e����C����6�I�O~�*O�'��i�d�/��C���q��쁤
>����a��}m�Q�c�{����o�2q_ߩ"�L��E��<;̝`n�{�
ɦL��� �C×iXN�}iP�6��~���G����i�e���S���f�Uo7��oϽ�>G��{�a���'޽�4��'Q��$Ru���;�c=�2d�l����l���~�@Y*L7��c!�'�¡�~Bu3�����{��S���_���^�io��5�J����A�-�K�s�h�f��t��+d>�Λ��c����nl��X�� \'V޹�X=��"1B���Lu���󶍲|�C�z�U���b�)>��v:����,� ���5�Q*N�N�,���ˮ��fT�Q_�xz��mo��F��@G���,e�{�3�G�&$�,�MP6������	���}��ԓ�va���}�q��=fχ/����	 i�Z��4����׺���޿}�5���)4Ͳz͡���c'����O��I�ROo����n��9i��	��yg�&�����}��΢�b�󆖃�9O|����H���}G�����}�$6~��L�Cٜ�|���C�h<�a�'��$����8�	��~�d�=G��||����Ȼ�)\�>��2j`�݉�_����!�Y��t��~z�iyd���a?3�s
��4��gr!�&�a��>I�O'��I?$����D{�GO�ϼ�<ם�>�i��5fFc[�1���q�����#�?O��2d��aԟ3�CG;�a8��=�w
�Y'��>r��!�}�Y=I�_��a��_�^�� m�}�(✜WFL]^[�ۖ��=����:=�|0�|t8��O^����s��?!>Iә��3�O����Bq��{�u���+'ȡ<��q'm��s��.��[���2�U�H���������̇�N&��'䞽`{7C�3l������S�����L����:����W�	�C���*�N!��G���d��G�y�8g�v~}� �=��N�|ɻI�@�L��2�����	��ya�M3�ܳ��P�?&��<��'��N�=g���$�Y1~��\�T蚁\¹��I�.�$��"���N���O�Ȥ�I<ys�	8���l�~�i�`{�3��>aԁd���Җgw�}�v�v�������̞��?X|��LE���	�1��w�u�7eI��'�=� |���&�)8��O_e��!�`Vm��wI�6βi7�x���[���Z���"%K����1��x�<�ɖ�4�b�3�;�x�GU���q�ۼ�X�Ђ�m�j�*V�R�W��BEC#��_bJ�r������d����]�1�oVa��	��d̽�`%B��n���W�*��]H�5�����<��K�a��?;�3�{O��S���y��������,NRu'䘋9�!�a����d�0��i��wy�>I]�bN$>f3^�q��][���~��ߞk{������w��L3�C?'��I��M��C��8��0:ɴX��l�hy�rC���Þa|��d�3�>F�<���"�q��u�5U%>/��;�}��d�t�2C�����<g�7�L`q�RE'S}��N#�dա7��Ɉd�C�_�ӦH��>�w3��K�!m73��5�Ėc|,�>��>3�4���}����	��I�Bo�4���gRj��~d�'Qd���o_d;�c=9�:���CӼ�P4�I�����}������}��5����Xt��ӈL`o��m���6�C�i���:�6�ٯ2N��OM��<d�,�@�'Ru�>�� ������W=���g���HP��������V����� {��q�G���|�Y1&�g�(M02}�*g�M3�jyBm<`y�w��I�2��d��E�I>@�'m7��k�nzy��7���]��L���a6��~�|�i���w�`~C�<a��6�b��䬅`f����4�זChx���0�{���}�A#ޯ�#CO���������������I���Zq����g�6�$��ra����s����k�d�a?'�9�&$�Hh��Q���H� ��Dzg;~	:n.���^��>��4����$��'Ι8�����O�:ɤ�h��q��y�9���'Rn�u�����s��~}d׼³����L�J��m!����߻>�޻����οy��~}�wى6ɤXw)�i'�Qa>@߼�>�I���a��Ct8��O^��vC��9�������O����q��	>C~�yӧ�{\?yv���V1{����X;��HU�8���h�f��B)ٛ�+�M��m��LL�3�k���4�NE�mC����h�)���Y��qwP��fL���	���;���\�Yu��bģ}
���=��tej��������ֳ�g�A����q���=��>��|ɴXk(@�'���$�2{��>���ߙ'�4�`hC�!�|��~�}��lqx|}�.1�2���ٹ�Z}�߽�8�L�3�B����Qd�C���Y:�!�d�O�7l���Ě`y=��!8��;���$�h<�|����,l}��O��b�6��^��SG{���t�a7����P;�Y'P���|�/0'Y1��E�q������w�:��M�#h@�M�XN>o�z��|@0�>��k�L8Q_^/��^���i=g�y����|͜��u�w}�Ć����d8��LE��!�O�v�,'Rd氬��$�� |(���£�g�i�ws��u����?y�����=����N���Cl�ɤ���$��g��`u����|����!�9��O̘�=�C�1'��%���υ��>�Dx{��]��N�Z���<�̶�}�0�IG�����0�'�u���d=���?2C�vì�&޲M�Y���|��1��d�,�!ԛd�a�=�@�<��~��o7��|�w��畟zj<=G��`��#����&��{�Y!����N2O��$+'S�/XJ�S�P�,���2���K��쪽ۑ��^�nڟ����LBmAx�j�e�#}�����xf�x}���m�Λ����7��ZKt�e�֠y�<Ncz��:�6��r���w��b[�,�0Dk{����B���=4�fM��<�k9{���Vk��V��*]:�@�:a\)�)Q�x���2��0Z�Vr�4T�����]���8�]Ncd{���V��N�լN�+���W��_k�-*�c^>�R�I[��M��%���j��8�Y�#-q'@���1R��f���IJ��.VjT,�`��4���k�QۡK� ��Q�.�f6F� �ٙ�,p{I>+��_��
��� #SH�*Z(�LD֫A��U��j�sOJauk%���E�$Qk+Z�f

M�Pef_P`�+���V+â����vnq���~��r��u�a��*}��*�B�I�W*��d�����xW�M[&>�gfKCF�x�b�e=}�������H�������T�ew	%dGC��G[�Ȭ5]�D���ޤ8����9b��^��ŧ�.�$Vr�J�u�J�;�@`ÄR��Ůt�X�C��T��o� ��V��������u{[��0w7R�bB���kG�*�
iz�)']��{v�WP��d�o/j>���3������G� Ȇ ��{�;���.���y�X�qoNA�P5X;��XH��j�S:420�ٜ:��qnMV�䥊5����p.��\��vc���Ю[b[yٝ��>�G�<�l.,Pg^��8v_m��%�U×Ư�h��\����6��*���Y����cJ��32�*�*�vt���^�˧��>��ᖖ㏙�����LB�׶�m����ũ#����q���t:��=èvu��Y	Њ�[]��a=t�뺉Sw���j��cg�� �f�X��;5tt��b-�[&��2k����V�V�B>�һ��Sw��t3���	�����v��8Ed/��jo:Yk�Vct`�k-������˧�6�+i+�'˫��p�����Ďm��(�;WZ3�0���ZU��D�����8	�����޶�2���I�#K�pr$'����T�z�'år���+V74JǦ��:Ό	\��ü���^����0�S�v�L�����.���]C8ƕ;��o,.{�7F�mũT[-���E�ӛ]�A�u�>�6t�)j�����!�o!��<��a�e�@��� x��q�#
@5e�˾��h�+L�Ӎu�,�)��|]QH�������E��n���
��gm@�c�I�э{{��ۦjf0`�����=P��u
TU�]۷���|۸;Et[�]U�_��؈УyG��d��F��B���s*S!G�c);hS�neC��yth:M��y*Ⳏ��ƐѨʔ�����U�f���kc�G�t�&��f*b�a�@iY�0:9m:�WI����S
�����PJ���,�!nd��(!P�.�ɂ�]?��L�
�]Q��yj�+�P/.Z�T1�P����q����k�׾��f6���������Ze�R�Z�--k+Tm.\"�QF��ih�m���[Z��E��h�[*ڕ�R���m)��J4�1�KRԔ�b±kU*Q�UEV�VV#T+[j�YU*Z��*T�X ���U�ը�R�ڵlQ���R��jVV�b�J�j�m��KVƫQ*Q-�"�Z��	J�U-�Z�Ң��e��b�-(R���Z5Q��B�U,ieTZ�ZŭZR�ڵ�B��6���mҫ*��iZ�ʶ���VҴED����Zխ��U*��aR֕��V�V6��حh�i-(��J5��U�FmA�ETl�D+hب��R��KV�%)i+*ҵTl�X�j�UJTm@QB�EaU����UYU����Ō�me�
�������m��EEPR��*�Tb��m���񍝪G�ˡn��Kk�gM�y�ݛm �վ�ư���������r�Hf&��S[�j���Y��zwO����N9��2���2W�S�k|(��~��b}�x�s�d��R����;ϵX��ݾɬie03�����ԍ+s���/�3Ϛɼ��Y���]�Dk�h޻�鵇dհ#z�lN�!�)1Չ�J֥�Vl�\"cBǮ�GJ���pH����j��g��3k��\�1Y�a���<�t�	�^����������<��G\�s�qZ1�ײ�WbC�W>/�_l�>X�<�:2$n�gp�WY���8��b�R�9�o#�����+����ǡ^�k9?-5�Ի �HK�a��W\.���V�VWO8�c	c�����R-���֮���T���m#�s��<U堲�W,�5�e���M:�]Z,J{W�-�n��>b&zz6=%�ڊًڼ��z����n��9#ͻv��1��BXi�]��+����pm�8b�����5��r ��w6�z�׉H�UӮR{Zk�P��ȳ*�-�Py�X��]�ym�=��M�W=�`��j���`��L[�N�͈}�@Sc���\�Py�jط�gj�d���'z�÷:�0�~��ﾯ�Z*J�(+6�.������[�!�)��v#:4B��Ue����Ӄ��6Mt��,_�S�b���/���C��>tfܻ���f����3Ou�(Xb��]�}�F�z#D��0y;<9u���W�f���ēQ�!gEP�qk�.�q���z����cGs�ŧ�CK2oX03����������C�Ӓ�߀�f��a�L�<�U�6��v�=��x��}G\^|g���J]���V,���ڹB}s����.s����SQ�s$��*yk|�Ŭ߻���L91f�4)�Չ�5�c�:ad����z;/�=*�����asJ޽ٗ{�H��>�jާ�޹��Օ�+4�`��^��<㗝z��=
����m��ݎ=���X,G^<�q���V;r����{����bT��K��;q�Ұ萙n��ޘ�c�-��1�Gn}bڵ<�����l�}:d�aa<�!W��T+׭�i5+w�y$�Kj�:���{�mRW����=�œ�Aa�����,4��)�l�X�#H�!˷*P�cYI�3osM�����;��g)��ʡ*������#/.2�i��E��!\�]A�*��CgX
z=��n�X=�A�;��1w���k\g��P��N���r�s]*�m5[���=\Q�7�p�綂��qC��4WSB������l���cM�����Q��K4��+w����mr��J$̪��P�.�mQj}\qN�M�[X���_n��j�%�8��}�S�!]Q>e��Y7�zr���etO9@�Ǟ���<���q^2���T�tk��T�C�,F�B��0��F�u�S��N���t�4�U�w+��*w�����s
�OF��0o�*�`w,r���^�C�z�a����Cה�W\�{����� ��+L��"��^+��urPz�s�!�nG�M��/7��{����[P�R1��֪7�����J1K���5�ʝ�7���sn�b�����E{�6zy�a$=-^; )$��\�q�陣o�<S��U�#�97������i��0�:]f�@!����w)���E�"$�R�05)خ�X�V_�*�w7�
�櫝1����Ք��ãf���K7o���)����HX.vǥ�}ٜ�զa��\:k�x{�{�6Tl�Q���Go7{�\����0�x[�&��3z��-��pQ�Mحq�{Tٶ�l2��T��(��^������M�_���7K6�f���d�E�Zy�w�a�OUl�7��/Ǻ.�m��&YZ3N3nw��.��#��O.��Xj�c�jX����j�Y�3�9χ���'A�N˫% ����H�Sv����˝���t���%�k�%<�"d�/���)fv�����aB�V���P��'R�J�+�:�q��-Ј}L
���"�*�o�wճ,'=!JæC��l����\]K��-���%Z�!e�,t��תJB�W'��HJ0��U)*�cwuت{s]v�5A�<W���ϻi�ntT��+�N'�L���oc:�1�,[}Y3w���^���uq�C�V#\���(x)��gC�*�&��P.zy���GWe>��4_
ˇ`��ͬgp�B�Z�\Pnm
��f�|�s
_�=k��p+�Zh]��x�:`�X��w���Q�q��+ 3��f��)_U�Ck����������H�@��0�ޑ��G���X���着�F�=4>��,O�I�_�	k>�A����4�Qz�+�Z�zLM6b�,ݘ�W���y(Q���u�p�4S���%
|��.dT	��]�����׺�Յ#U:��Pڃ��#�"U��b;c� �:�͇<�;�A��;���_:�cw���oUTVW]�Y^�� ��x�	[)eS��J���xM��Ym�nFN����͝� ]?]�g����DB�\����|��ِk�X�#�i�����z���z�g\��nWVּK�^�����ºzs��HnSc�#�f�V�>.�o}.xZ=�Ku����
euB++���\u�!�R��	�����W�MK9ݗ�U5}z�Oovx�����c7�i�l���~:;G:l��_<�P�W��Χ����󮵥���p�O s�e �����>��b���؟?CX��h�]Ak�:�ܣ��(+f���5���]�R���1�Y+϶��l9R�m��O麶^K��;���ݮW�<Sz1���S�.ǈz~}}Q��|�j&y
{}H�+��f�#W7�,f���K��t:�r�c/�B]4�������F�����==�U;V��-9ٮ�[�t���aa@�ޤ����<��u��5�wg���V�Qջ	��X޹ʖ�M��_s��f�кѻ<�E�i#��x�=�Ζ�N-nB��S���E�<��&��=�g�������2�e\�tz��C�^Wνf+�ғ���ɼ�Ĭ��v����Av�<�ѽ8y�累.��f;0�r���%jbq<�`sq*^�p�[�lK��ҭ,,��Y��꫗��T���.���l��fq�9ݖ�j7��n�e�4�DF�|��T�H��C�P�e�(
/�EI�+�����S]z�\��{�����9��Y�<�缱�V����<�`U\��w1�n�P�nE� ^��U�d��m��ri��r����ԍ+v����yՌ��s��C��$bZ����=y\-�����}]6�+��\�ʮ��1
��5�H&�o�
����]~M�8�(����n�n����3�`�@�q�p�b��2P�Բ(�ph���о\��wdİr���7A����� �RRJf��V�;=u���q7���^�4zj��ާ�ꎗz�r�R7�T�.�i���p!ZV�I�̞׏�8��]ԣ��f��dL"��ڵ9���k4�Ԍ�V�.S
�X�}֛�N���5������l��P�=S����_4�_BH��s�����|�8��XtHL���n%����Z�gk�������op\;�s��(�hbY�>7��ͺ��v�E���YA�c2֬}�q�Bcq�
/�׊ٮ�Q:Z�׈��ϻ@\�ыe!��t|�aǞR��A��cz&&�Y��g�˪��'��������5�.�땹�r��l��+E'P��̺��R�˕�@�р��Xc�̮���v%�e�ޘ-�q8($����&Us6��d���ݞ��	�G�����r#�����7�^�:�K8�,l��.q�Uw���zO"���l"��/=�fw)��\��c��Dj#Y�;����8����Ȉ6�OV1�C��ӳ�l�lO�V�Ne���������O8��3��D���]��Z�V��Q&u�ؗQ�����������4��Hf'r��W1(B�["m�^�vjh9]���T�8"�!X�T�l������{�g��}�=�^�6���?a�z|�ug�h9L))�|jlhB�;���fw2���~�+I���G^\��+=�-��\_:�r탖iP�.�ow5J��/x��r+����r�%^�Sv6�^6"3<t�����<�{U�}�.����p���"�^U�m���χ��KQT�g�f7Uԯ�����5�n@i�^7�ksvm=��k&=o��25���Éè��T��B�4?\��'1���7�V�𤶓5c���R!��g_c\�V�*f�٦�P��z�.]�Vݎ��~M���O�-������7}�3I��q�!��q�>�:E.=^�j��>S�Nn����a�Kv?���<��B<$�X/�
�⸤3m�ĳ��L>�T C����%�G$5��x�؞���	�a���C�P�T`WGؤ�Z�=�^ߕ�V:mM�(b�7���!a��t�L��N�;n�����ܻ���
8;/�U�V�]���Y�+�۩	����]�w����m:���0�|�L�2]������wv���}����yOD��K��М'�PCLy��6YA򱕓b�%��������~�N��P���%�뜭�@��D�CXt�{��r�R;	��UM�YA,�8�mؗ���i��~O`J����˨8p*��]�5ݘ�m�=bx�������Y��l\����9d8z��1۔�,e��y^�M�#,�4:��1W_�ϖ���L~����'��y�x��
�����<y��ؼ��e�U�&v�z��(��4<& ގ�WdnT��B��`nUY��Tͽo:���Ń�C�;�)=�_N.�ײx�P�5�됷��H�������'�vߣew'���oP,+�V��7�=���V%��Y�Y8�o��Z�k��T��5wV���h�ݬ0P.�Qb�p�M}���rb�ܼ}���󸰅f��Sj���U���~̞"�=�)ui�Ӏм|bY��J���X+�u藧Wy7/�	2"�9��k�>�[���Һ��]M�[�]��e�4uQ�`�����.Z�S|y@ۘN��o6�m���j���#��۴+4t�D���נQ��:V���}wW�Zö@�ixx�u�X���Y��R�`���;U���m;�K|0}U_}_R�|5N^~)(�o�����Zb�dݥw1��>�v��Ft3oB�]^m*�ʉY6���i;��^�;z��,w:Fg<�z=���r�X|֚������4S0:�R��i=ʸ���G#[�\�;4�`uqF��V�y̎�ʑ��P��2��N�тe��8�q�3��k
co\��um��p&"K�!=<��g��:#�B�XĞ�ڇ���4J��۪�٘�����/�A�jgO�QWS��VGZꃫy�\qe�o���+�H��˥;u�.�J����*�~կF���^ꚠ���Â��w�Y���鼷H܈������)�ruz{}h�s����T�T�t;�z���<��p�L5x].X=9��
�� �[h��Or.����y��O��(P�u��׷�oV)�<.@q�^��'�I0�+/���<r��Mb���uL���YA�񰋮��w�L�|��o�7���Xn���ι��K��>�>�ZIn��i�����bn��~��t��m���SH1+C�q�bL�
#������v,��b�I���e����K���wv���Z�0w;a�]�O%bRJ{|��ga�CqhŷK(�6�U�枨�:~���[uu`����K3��� ��N1�P��b�Elo|��e���K�O@'����T�c�m;�u�l���DÝ��`��k�곈�;�]�^*o���
��Em_m	Z��H�AjʾO"��F��V��*�+3�<�f��W;���q�+���ɧ*�� fA�gzXzS�zX��z��H���yΛW����Hf튾n��R����V��5���!A7}1w�c�|n����'b����Z�7�ΙM���2x5�2��\R�56����2uM��o3�H^�K�=���y�"����Q
di�{�f��q(��S(��e���>�gj�ڻu١�뺙��ǣ��m!xo��>�㋦�$ƺ���O��ٖr'/��r�,Ow~��`A�-o���"f��:`cz����:�� N˾ȡ�Opʆ�J�!�u�1�qZ���鴍�&�e��*��ދUrj����,���X��f2�_T�f���}Ѯ�E����U��&[NN޶�k2��X��kz�����)FdE���s�V���ְ!��u�/G�����u�aa�K/HR�������]�����bvm��r�%p}қ�́�m�46��'�Y�'}��OX{��f.�����Ǩ<�ya�$w���9������7[��;x�����h����:y$�����i%Fu+���=u�'wL%;���}��Q�	��O��e��ѧI+�Ww4���p���iz��6bW�U�V��"#c&��d��kh\k�\�[y��+-)ޞf���$����� �o���~,����
x�,$|m�s,C�{z��Rk��JjV|�Z ���ʁ�@Ҩ%��$;�&���Jpo��
n=3M8���[��o%o+C)�����K}o�b�,�"GW].}DYM��Ui̠X$������}�R\�O�V�$�[�������ݩVBu&p᧳����QY����V�!�k(�y,Ko6B�@��L��LXo��i,L��Q��5Qy)t���E3tV�R�o5V�&˖wf��>�˔R�n�VV�W�w�����w���5�����+Xot�\�3P}H��|(ܮ���N�V�6�[mݬ'1RB�n��v~i��X�N���q��.�
��9�ӯke��:ݦ��`M��˩��=W�n�,
vI�&+5#t"���@"l٦O�x�Kv���%�V���)��$C 3"̩RH݄F�����XY)Rɶ�E��֗�����:�X�n��i�U���EB$�1f1*࿥��0���Ĩ�K%AUZX5��jUHR�R�Z��Z�R�-����F"�IZ4T�%�TejV�e`�R�XUhµ��m�R�R-�����
�Uh��F�X��m-��-ZZ5�AeF�Z����+���+X-Q���V�U�R��Q��5V�Z��l�em����U����
�V؊����1XT*6�(Z%�B�dX�AJ�R�iKZ#-T�Qm+֕�����X����1�J+Y(ԩiPj�����V�XR�Q���ڶҫm��iAe�mPm-�jFږ��l���*���UV���*%j�Z�-Bҕ�D[-m)h��mB��V���dPF��X�Qk���jF"�hЩmZ[mEE�h(-aXX�P��ŕ*[j֕�#l�,
��UB+kkj�X�*�o�J��c:ዝelqS�뢫�ʒ�*�&����G9��}�������5�K�zv�T�=��JG%~����{����1�t���)o*�LV��"Gl/}�ޚU�Y��[ր��E����ם����g0}�����<v:��X��J���b��ć���x6��et�p�qm���@���ٸ��@�=>��VT�~3"�L�9y��+~1��Lpn�����۪0iܾs��'�d���X��u�\`QW���Î5�(��h��{*F�Y�;k�;%�3�=���R�����d�Cg�{����7<(i����o-�&<��_U��W{'U(�Z����f��6���׶o��4��!�R�YយG���h(^u����[�6�d���:E�F+#�b�qS�W؎�iN�"(	e�����q��n�n�1u�KE�S����D+"�8�T>��u�vM(^�zձ3�1(�R�.�g��]{.�#�'����x�ϧ7�'�x��)}|��]4_�����93���`���M�T�C����i%�C[+l�K������~>������#5T����s�7oq.w�I�7�T��6�V.��5
#�XFwQ�e�JrV���`�{\�N����l�بG]�e��r�\��6�	�5�n<��z�������t�[��Pص>�ڬ-�4�:�Wn�Rڬ]��J�����&���ֱn]h�;������	m�V��.�'9T9 |d.�X'-��着��)�c��5��=�ẫ�\g�9Ŗ=��R�aD�����7��ƽ׶�;��Rr
�����m_'��:@e���C�j�ʺ:,O��Q��5��-��{k-]kF����YR�o�J�K�Qw���0S���Y	����"ջ&M12� {�e^�K.�r.�:4���6/�p+��>�dyd��nJEWABB���eWGΆ�:=�O]�I���[��6]��g�vҭ�?/�x�0ǃ�tP�|�sX*��I��]�n1���}�ݞ��Þef"Tgk���ָ|oo�^{({���Xp��x����=�+<��=}[���ͽ�����X�t.Q)ο2�ÏL�^7Q��uB���U�J��3\[�~g�\�x�8u@����<��ݒ�U������+��H����^��<5����I�|d��}�v�5�8d�����C�2�,��w�7�t�X�Q�k3�N��w�aY��ԯ�j�KM�5	�j;��d��ґ�P��Z�ny�w�oU������J9������G�Nk��Uf�ީW;�g6��Y�U:�챜5<�WƎ˗J�Wێm�3Aݩe.��[��4�x����y�ۼ��u֎�YU�9v��FGo��)W:�n�X���ٷ����Z'�X�<N���W�/�����A�î�9�EQjB#����m^^E��6B�K4�˨�lLvE�tR��5�8�k�l߲8�����,:�5��:��y���t��)ڨzT��Ig�UG#�����T7Þ�Ɔs���/�'*�\��3!�*���~r�O��z�p������ Â����I>K��kC�u���B]@�ޛKN�[{c�)~�!�j����CԼ'��V�p��HpИ^�Z|���2wJz����j��,C�4\*w��7q�;q���a�1�������\��^�s����~8��q6rp�P���O���X�k�r�
���|���\�\/>}L�`��R�&��_{I�abT�	�_S����>8-��h�j���U0Q:�U'�ù�w}��
�,��'HO�U�7^�Q���y���Zs'�:G+x������Q��t��A�u��Z����j�p�;�a��x:�[g.��jy�����!����{����]�)��#w��HS�J��kB��ut���N��V�Thyг����[_E���^_PB7{��A�B��Jq�b]���sDĮ�Qו#З% ޡ7�gCۻN s^T�e���w��mN�"FGz�]ꨰ������{����.��j5?WK�((��٣�ZU����x�d��ૐ�ǯ�V��|��^�˷��{C��t�L�����*Y��#M����Ps��g��]��%�D�2 o��b�6c\�8k�iɆ��e�8Y&�,��Uc{�b��˘�����`�'����>�w/i�u�`�ES�#�.Ύ%����k��[�nD�N�-�Z�{�uS7j/o65E���������풐��/��+���s�5�s^�=���V6��xf�œ�19L�;ɻGTnE0-�G�R��kMXH��t�(n����ns�{��tG4��F;z�ndwE�ʑ�s8��(�#��81�ҧ+m��W]�$q��#H�R�BQ}���Y��Y��Q~���zY�Ϟ��2�޸{}�r��%�7�2���cGF�J���5�}��lxs�4&{Tm(�o=�����4�畊ʿ^��/>M�,P���+�ZC���B*�W�߼���0@��%s�s-��1���OX=(-/1�Su�;�1���@j��4�������b��Z,Nki�P�`�T�.�n���(r��u}���6�L�"O�Ҳ��¤��M 9��=� Ζq3��8B���9�1���5��^�V�b��x�;*��b��7">:0V�4����i|�l�n�,|���ǮS��9�5���y.��_�*^Ξ�cT��o�ʴȰ����3$:Rp��=x)q�|F}�r����]�u��nc]���Ȑ��6i�e��]�a�<��<%�ZZM��j,H��zc2�3��Qy�q�~[��j���KF�;��{A�1�k���e�MA1]��N�a��پ�w�_wp�^�ᶨ{n���7�d�D��loT§%i��ES��IVkKTW{�&�l�Ĭϭ�x��i��BE�nM3g,-�UDE%OL��$�m�s�z�l����+sK9��~@���x����++�_�fEW������\�y�m�*lz,l-]�xo�هx绶��?O=h�w�}<E��^�
!V��Ay�5.X>�K��C��9y���*W���cu�Xr�b��;F��:hKUj+N��$q㕹�kQ����i.��k4��e#F�8S�{]��2�=s��xt�Fo"��W�k��|��=7��6�s"iV<�ۓ*&v��
����� F-ɬLv!p�lL��h�w<w|���4f��G����j����`�b�M�#l�g>��$U�T�ȍ�؟�+�;->{�M��f|�k��w8�F����Ү�̠����ёV�l�T�ͫyN���\�L���`(��2oرL.a��0Ĭ��x{��ӯ�]���Ə�4OƅҢGX���E�"�],�D��C�C���9w;ht���wbB1Nn{B�8e�۽��~�*!^Ȳ�xb�p��At�����t҈��'�*�b���bB�a�2��ͦ�8l��h4����|���Uq��=��f���!��MxG����0+�}���^�ǁ�G�K;c�(D*;��OYuS[�>Z����4��0券�mw�^�<9b���O�\�b�r��:�X��!Ne x�H���+�(o�PD��r�i�L�Wmޮ��j�U�*9��BM(��W{qI��t!uj��,~��`��=�/۶����ֻ��}<A��e�3�^���N�DR�d+qU��j_D�
�5�F��/��n�����kz���>�c����˯.*�cҫ﷽��b����W� ��;��1�d�z�y�r�ҁc�64�/
��K�E�&xW�ɇL�;���ʹ��a�vcS��FaTʛI�����&�\)-����W�b�V�ϼj=IoQ:,�v��V��Ѐgt�Jv�šXA>j:N���~�T�=�E�r���yg~�ڀ�=�l�-��Z佻����bd�OM��wg̕GvA�rN҈u��ؤ�9�_����X�@��u�r�u1rN}x�%f�L��T	�o\A[�:zʬƞ��V�z��׬�{��"[x��^9�����J�J�9��q�M�U�@]_�!}�1�t����n�Pƌˬ�ܴ�v�,m!C6���{�\U�R����.ɕ�}>c�b�]�X���;��*Oon��� ���nX43e�kד�#Qr%c���7�j��jMØ��/1�����$/�ͮ��N��fަөh�|On/�ΑeXS�B�e��uS9��k��qak�c0{�:3�<zW]*Uxy�FÆخ(��mŸcT�f�y"7�V����M�R�ѳ�KR����J3NIgh>���ǁ���*:��\k7{49�fuA�7��6��V�9K:��\���q�����;Z]�@�C��SĚ�B;x�E5���٪��ʹ殠3i���V����D1&��<�%�"Q��z!%pn��]\�T�[����As�c\fS�Y����g�:{=%1��U�W"oL��n_o*���b!���Ǵ��}�H��vte���;�]WլtX��	K��$˓z�n3v@�1۱��5%���4�ժ�>�+d�2\�k�'�Bq46�f:{�l&��<,bL#��j�,���zo9ml��ͤ{�
����� ^��}�7�b��סi.�����?,\Ьw��g�8V��D��*ˇ���d*�̬�6�I�]"3�j��t;x�J}O�Geײ����8�Յl�+ތ���t{��ZG�����g��aB:I�*���Tf����S�qN�N�#odR�ci]���*���/m{�<ut�]�V(<��SJ��""������V��k�����l�:!Er�1���E�N�G�̫�SՀ�P�DSFp�^�&����)9Z]�;���+�Ǖ�/k��td����M��v�dKYC�en���b(�T_������Ɂ��Os�V/#�ֺ�vp�볟]8��fx�y����]OT���ثɛ>�����#�u���z��qں�S��y__=#�{�-�RV�k�ˬ�1-0��JD)�JXPk��i�ޥ���9[Sbܳ;~���@K�&��TW�lӧW,���<�Y�\�Ȱnnܯy�$�E����s�Y���G:]��2��g�c�`�<F
BG�,��*��D�wAYF]Q���\��]#vk�Cp��2C���2X�J\U���Stx�7�����xnܭ2��ʭ)��]7
�w ��=TjƇP�ʥ'�{�rGx��Z��K��ۃ�Y*��P�k�e��If�yiW���� gvs�J���03᪔E�H��%dK޾69���6OC�Zu�|	�᱗9zq�'k�;�x���Y�Ry�Ż^�Ɩ�4'������҄35�7Pc�n�rnc�x�ɹ/��N��ht��JE����5��vW=�d��^TX,���A��,H�U�b�R1��]�k.�c����%�<>�}P��TB�3�nT���)��N1M���$��<�^[�g��Q���{�Dl�;а��f�=l�z��Rbq���7��z��Ru��"���Ø'���y"̓����}ޮ.����x����Sg��1���N̗�����J�U��������P�����<�l����ͻ�ų��<����H�O�����a�����=^���Z#	&7`���+��%��P���T/;h�˨���{q���OrV������䵀��h��H���`�����K�sX�Lx�Y?͈������}ܝ!~�b
�����Y�?)�+m1Ն7�2��яMt���95��˸
�U���j�b�c�(C�$˩���ף,�(��⪇�絯Gq�R��2uor�������(��2xgM��R���Wރ�dY�@�&��:^>3�c����ƈͥs�u�hvn;f��jj��Dzc�B{q骿��x㊕T�Y�^bX`|9mn��r�U�]���p��x��j��nE_^��J.+^i$;����&uVOI���й�V�=hS�/�x���nB���i��wz��:vL
���ʶi�kY��~�=��G\i�n�יĆ���x�Ӽ��c��n;�NqF�F�gK�n��ZJƌ91��~��H#\(�u"�zR�t�QC�{f�J��ћ�X�3PDs]ǻq���T������<jܒ:�JF0���8��}��.��-���Wz�W�󮭭�����Y��J��`7�ϣ|p8�!^�(�P���Ӟ(�*�Qq��`��ɞ~E3~􄲰���ʿ_��D�Lк0Qf��.mCʔl��!&<�e�W��d����F.{�`ھ���V��C�����Z��Ƨ��3���*u�q��VA2��mby����C�{;�c��3�o�̋l����<X�,�⇬���:���S=�]�n�櫭�J�I���]CΛ�:x�S6�[n�2۫2,;�f���ia�%UQ��\#)E��ΓV���+�YT{��X�̗e^.M�f��{Y��&�f�_jZA�1>wm�k9�-P�]MW��;�r�;6���ۻ���_n^�8�Î�C�t�O�1�k����M
�Y �v(
�G�g4;����w�hm��Ņ��u��w�<]��Ւ��x�:�E�2�puͧO�0��9W&�t���a�:g9���lWJ�n��ge�e���陣I��wniK�]��]!�u���xp�x^����Jn*7�ul�Ш!����TGP䲒��Y˺��h�I4���ML���,i�R�G�}�UA�w��	�]���Why�ҳB<�qX<U$/�i��F��y+��ً����@�˶�j���.�7���UDr���P��B����Wh�fC��偛m�Y����uG�2��B�I�6��H)wt��{$#����߮bv�sU��*Y�y�=h� 1���یQ��u����y���;��|��N�����t&uc�KL�]jvʹk#��<�n̉����󙔜��t�`���5)�:�v⻬��8�Tw+���`�qP�5�UvhʝDu�����g������S��m-�т�6��7����g������%�/�u�[W�sR��B����U�&v����.^7���S&U�����:.)W��m��iA��s����ٝY���τD�O_5�.��<��`�m+vm��6��R�>��v��U��wP�\�t�����˜��b��3��7��S�����'�͝�y#Xq�X�j�����1}g��յ�y�x¤�)]H�+�]���שN�i�T[�ŏ��vv�E��.V���X:Va�D(tΝ�:A���k58m�(]���e��W*��Iuhr�Z)��fƓ86BQ�ʸp����Ze�5k\NvԦ�O�{Zw��mS������6�65܎7�օ�0����Ʃ�҅�I�81�?��Z�5�۲e^��6:ʛ���:/GdI��uk��F�ˆH��bok7��j[V9���;@��:�����"1�"z5�K��.� �-A'9]X�����Zݖy�����~�;�t���8�bm�D�1��jQ|�]�W:pf'��p(�j�ˮ٩pb��n�*��J�݊�$Ts���6"���(p�\Z�p����>C��WZo4�k:���6�Ҝq-�z	%�]���l��N�v�3���.���;""������ք`��tajI*����pd�ڸi�J�!�^�����[�J	fwq��r�t�Q}��J{�j��唲Hy(<�Ǹ�y��J]Ą���q/�C�ui�C�ڇ��WA��s��6
�����w9���ip�K��n:Ƹ�_V��l�r�`ޜ�7��h{�x�L*q��Nv�5�gn¢��R��0��K���sN�n;K#����4���[��ڇ�b��Sʓ�����wuww�(1��֢��҈�Z"�jQ�5[ikb���bR��T�lD-iKB��VصK��V�T�KJ��V�KJZ���F2���+F���҈��"�)XUVDAeE[�*��"���TT�VE�J�X(��TQRն���X�ED��j�Q�J�jZb++X�c
�E��b��F�X�TQij��)[e�Tm�QU5(1K[FЭ��"��-����YQm((��YYV�[T�ZҊ
�i[����ZZ����U�ʅDU��!U�F�UDb�PD�Y,V�ضѥ�*�4kKUEDkQ��1J[YPU�Q�R�[�ZիV��+Z�-�YR�j���R�����b6ңJR��Eh*��m-�Q��h�V�-�bV��-*"�B�k[T�[Z�[J��ȫF"Z�e��QE�YX�RR�j"��-
b�ED[m�mT�-QX��`Ԫ"���EX"�%eEZ%@���U�"����jQKA���F�D����"��E�X��R�-�
���o8�h
f ^�$ft��L�@�=s�>7Vp��Mn�%[ѝ�
�f��/7r�j�}W�L���i
�J3�� �6�-��x�,l�71�'���+cq��:Au�"m�`-G��|wח-���,S-��<㜊�z��;ih"���#V8_��bx�ZW8(N(x����#�ň�ҎQ�5eO��j2��s/إ�4�'��`VW.�>��3Ñ0�cn��m��>�Zʄ��6ߙT�Jcf/	�-e?*̕n�Uf3���"em	�pR��}t�
(>�rF:wYg�P���Jcz��;=3�yx����b��h`�Ŧs�����]#�*�F���/����gòVj���6o����D*���Y��g9O�7����1���/#N2��Y�8t�xu�׍ܕ���+Nոp�epЕ]���e����:�����0��KC�y0hf�$�F��_�J.�]��!�ɉͽy�l�Q�Ie.���k{՟j��N�=L:3��|OY��9~UNZ:�$�q=�ތ����O�c̬�r}8�ڛ���u�(��@��0�����.K��w�}�K9����8�귾���L�K��ȣ�$Z��C5^�e#�ǲo�+��y*�=�=m��`�sw��Oj�Bf�ڜ£X3�ʰ�gU�짰��y�����G4c��;p�����3sKݣΘi�נL5a6��N�	������ �s�A�����5p��\�ĳ�n�+�G�=WOs�:!�ꇇ���%������)�r���!�*JJ�z�dY|��X���j��C��G�\e�W�� ��<�\I������l�<�5;�W'5J��J���^r��Z#*c���y��0d="Y�t��Ś%��y�/{�n�
՟(�(�\���P���r~R�_�:�t��~^�U����<�oxܺ͝��Z�x�Ɔ�z�9�῟�	(���c��k�r��u;gT�PT��تb��}��B�WO�_0�Q5�[�='�|��(�;@��V5���+^>ؒ��/e��*}n����6I�B����UZ�z��F-��z��$����o^=y����в���u'�C�s�ixN/T�1�g���S����{uL��7����;8D�x[b��R�����o`h�GiT���x�%�Bǥ�`��mU-�5�o^zvm�1WH��L�ܚb,la=U:��g��(u�Ϝ:��������po1�T�l�tM
�(f$��Z��W��5uz��9=g����V�Isw�w��e���PE��y�rMt�р]]�R�@0�p����e�X�7~,�����0��u��c��*��%��I��oqoc[��c*s���R����x{��.��,X��;��5J#6F�87i��@���e�fsV�{΅�K��������U=�L��w�z�pdjx�"�g�!_#��2���G� �|��%������q88Tc��w�?m���T�|�+��ay5�,9��g�m*<��J��]�s��ڧٻN�*����sQs.��oϚ�_'K��%�R�3bc�`�E5�LU�8Ǉ6��%B�,����Dn)GH��3�̎谹R5b�C�6%@���N�w�ɤ��S��u�[ZhU�ק+5��҃c����i�+<z�Lq��*[f��w>\���Y�/"��$G0�qQ��ӛ�*�cG#��xu��D^vo�"U	�ܦ,����ڻU�M`�C� ��[�!�e�;�r��W��y�^��uƄ!��vy�4q?X�Y��g�Ss�L��^��\[C�c�t���T'(�� ��u5>�M��W/5ݳ�O�v%b�?J�w�iF���l'8X�|]�Y-�(M��x�K���fJ��A��=��{x �@�C�lԡ�d�[��{ٔQ��^�����G�n�.�	t{4�S�;x<�f�N�Z�+cWYV���R_Z�ri�ֻu?��Ӻ��힏��n�ѝ!䦄z��С���R���"q�\�o#]�e���l������U��UZԒ/oϸ�c�|U3crv`]��#�SU��-�����Use�xA�Ǯ�?xDns�sn3��5��vץ8m�����b-20�n�C��)X�/U�!Gl���@l{P���v�3}�&+�F�x)��u��.�k%����Hc�uo?`(pGUhus�{'t��O�u��,�45�x����ּ
�f�Un:(X����Ӻ$��\����6-���!n������N���O얼�o;�n���d[x��1���ʞ�6�Gs�ȥ��'�ϵ���?B��Kw�wv�5T���jw��n��A�z4���?\۾'(�B��<�Vu��k6YQj���#�4�sdw��n�g��3��a�}��p�"U����ۓ�����ƅ�ud�c��F�\Q�=���Z��}�^�h�Sܽ�kNNoWr�+2 y����f��zhz2F���3��#����w�ZS424)��anG"���J� U�`V���̬���:0L����0�Dr�Q�b�p�>�/ ;�v�����NNn���^8�A�I@W�Y�e�}��c���{E%�X��W�<��1cFX�f]#� �p�=���i㌣�E�^k�S�
�)��{l(�"꺢�T{�E�|^b
���J5+�S�ͮaZێ
�>[��9�Z�!J̍�s�x�l��T%�o0��cV�j�˥J_B"��&�j�R��Û⢮��<l�u=x��-�K�oJEt�����FLr�ۋ�NM�1a|;H���p#�u���/�Q��F.t�9�ISX���ؽ�X�8�Ĺ�턮���ˌ�Y��3��(ߐ�D8gz.��%�h��uf������6�ߌ��u��җ���3Wk~�h��ixzJ�c����*�J�ǠV��ǌ��r�����H�"�<+�
��O���Y���:�_5��*Pv�ªY^k[��F�{�1�n���gok'إ���=hY�~��-v��[��
�'%f�j��A�z3��|<�f�T7�5]F�	\��}%Z/���>1��e�C�uvś��m���k������)�Ӡ���"��^U���b�0r.�Cm��ž�Meo	��n��=����v��6Y�K�b���<a��DǍMvV�Ӽ�=oe�Vi�oz������1li{��E�mPdP�\�c�.�#:�ě���^ݛ?Oe�!z����tI�����%��I�,k����2���]$rS�t��Y�sñ)�g��ŕ��&����em�Q��2�+׀��ښ��W��ܬ�=c�v[�o���<�7v�����>�n��`�k��k=�sU��+T�p.�8E���}��T�+B�o��\��[���,��bE��)�U�qM�a�n����\��_�6|��}�t3�#o��t�U;^�wM�a�:��S��������B.��x7%��8�Kj E���ʳ��8P���Cv�Kl���^[�t�1:������>%T�PtH�(GWoT���'��c+L5m�9��ct"���J���T=�_{����:��`�����F�4.s=d�GR����Z�P��Fh9%��1��C��ٴ�*�9�筍yW-��	�T���X��qX������i�#LvL��X7���:��j��ѳZ9|�{VYv �<#<�h>z��=}:�<I��6��P�E. �fH���E�שf\�.<7Ԩ�Zmx�EZ��9J�{k<2���x�K���-BV� R(�J\�c�{n$1��k3���/XZKSσ���5��6z�����
��V�<`�����&��ͺ"�;

�� hu8]uC���u;���a9����Cd�ⓢ�J�/��ų��/�E�e�L�.�rh�Z�϶��2O
w!�e[���:v̘�=�$�gdh��ܵ�Y��gs5M��z"�{t��Jv>Ok^\������}����fM �|����'Y�M�O�y�/
7���;��X�÷�U�	)����W�W���T���W����G~�(��z�*�w衲M}��u�ʼ+Q�c�z񸇚��\vR��COn���B�G�,*� <yG����j����3��U�wY�:g�P6Nv�y�x�[w��ɯ+�kv�n��*��`�Zl��']�Dq��������f���*��7�g�6ǫ)7��yv�C�8�άM��� 8���!�`����uz���Pn����i�<E�a��M�*P5�,��e�w�^k\����F;s��+w�`%KT�{.pLa]�ȱ|֡�^"�b��>�|}o:�ǻ�r�OWG��3�|<�Y.��*Z�bl��V=+�ɯ!���I�����u�r���'��f9k�����p��TF�#o�"�]ao��V�>t�+=mE��L�k�k�*z0�v��M;ޫ���J"�~L���DV)G>�Y�<����ar�j��xKҹ���$��C{��ڮ�<�]y-	��huҏ����æ��Є3y�ȃ�mSd�Ūw^�66$͓� ,lY]�g2o�U'S��y�ѭX벺u:�Y�\[߷�91�@�W�&$���ec$Y���f�T�g��n�P�?o4V���Qp�M�]-�[���ջ'xWX̭�n�.�=�@������dd�3�.O�W�_rj:ޏ��'K����?�=�h�s|
 h��W��~�db���N�O�&�n�[�g�7.�sC� �ƫ��6��ZQ�VkO8k��G%�w������dӬ�4Or<�9T��,��W�x-�7",Y����&����&�,P���S��Ti���v�U�_�$itU�G��>����
#����/ի0͇O�ε���:Ҟ�U�]z��ŉ
���*�k�6#��GEe���}yك^�|��:frG�y9��Y�<���kظ��fW����\a��IC��Ft�l'��,�B�e�R�����������zQ��rS^��u��e��X�K�P��0�uVoT���s���n����X�T7�E򴡠5�x��O�Z��e��W��%
���Y[�:Wr�Y��e�B�ǶP��Y��c%1�[l�����+�R��W
�'�|e�.��Bj��s�י��O�Ǣ�au���ߞ�+vk��CT���=�ŵ�p���j�s�8�:�oFv��F���]��)O�o��Z�{�i!��bj�^�w��D�+�����;jsД>׸�@��t�niᗥvk����kV���4�Kc���{�%���tG0C�5
��Fn;�*��W�Pӕ�����vTHv�"}}�]�����k۱+MV�{j�F)�wa��H���Ӽ�anw"��g5�\aA�z'{S�ڢ����͜\V�.اSƭ�w��	��5U���zYet<S�wǭP47{kr�<l��_�-����7��z��;rR1@�E� �R��Ef�¥���۷X�ۛW/ǚ��Pr:��>��*�\,J�\�ي����U�@��Oj���۾ŧ��<��ǎ�Ow]r�Ϛ�0�A�Z	�ڬ���7�|��kr' ��O�;�^U��BˎRx��Ҳ;u�v+�F�[T�x����(M_h!��J��W�����Ly���K��Pqj�R�ذ%ϯm+��K7q�ګ2,yHf%�@(ז���fN���%�GA������,���nmu酞���)���>k��&��ёA�33W���$`Q�bubٷ�پ�@��-/	�ʈ��xc/���ǧ%p�����a/Z����5f�ㆅ�\��c;��eTk���+�����S^�����/<�J�
/)� �o������!�R׻17Y^Ç��AA�O��t:�׳ ���q󙝪uy{��5t}���5��8Tj��݉��z%�_5R���E��8���g-�y�H�OO���^��k:߱��v%�����B]sc��܄��D���Jt��ڕ'Ү����< ��9؊]R�xH��bF^IT����HTj���6�Hi���'�eq�F��s������Nr]�v���AŜ�#��R�"��U����^ÓU�m��q��Ie4y�{5{�y?D�{�8=�0iv+�0P�L�r�7�J�<^N�3�eA�C����*����_R���m�Ik�6V]%Z)Ko�%Y�T�V; mW?k�}��ٹ�v4+E����n��59+b���h[���u�t��B��c��Xzc�`�)Jυ�Y�V�ez�ռ��m��J	\�W�-��~��:�բe��өhq������9rZx�K�	�\��r�Vܶ�ll��G�L�a���ԛ�����=u�,�Hm������Z��zb��'aɶ�v��S�������࢘���/-��%�E�s*x[*�\�Cx]F~��7���g6��gnN;��y��^��;*mB(�~��{o�9�t�*��0�10�=��[�,�P-��ŋ�w�[�U���0�n�u�T���qƸgj����#�ˮ2��q���Y��8FtLRӔ�]���ܨr���Z�����t�	��5�z!H"��v���F�#-a-�]�c@�SV��hRĵ���e�`g�jY6e���'�m���VjQ��9�u�M���W^5�=�()MsOK=�"�zL΢'T�q�T4"�ޓq�;�V2�����Š]�2���is�Z/��ڔ�gkU���H�XS;'ruzA�8 �\ʕ��VI�G���"���*t��.�Jyw8V7�%�REmF�<���9�6uE��;�@S�5K�=��'�6��.�p�<$t325�n����.��.H-,]��
:��^�{2�����s�WF�6�ܜ6����o`̏l�D����s7�BR�}��c��3�S���3�m��s�ʺ;�&�V�w�A�Ո�]V���ۙ����e!0[�'����9��U�2*��nPڮ���I�s���T6��;�##z�\u��ek��g�޶��j�[U&�<Nt�V���@�+-�n=�1'ٛ�4��ۊr$~/��8���u=�4Q�k]��C��R���'�S���6d\��;pR8�(�<� ��ԓwb��'����!�%'ou����[�|��=�LRWfWR���e����3�)o�Q��U"﷔����1��7��٢��U��hH�]n�T��y���GӍ��痶x���il3��4t��զ�[�۔���ӥ��를"����s�!=�]V��<`�֩�7��I���%��2��@��|��L%L��.�Ȼ���_Iy��9n&�4�0�U�E��Z��|!��k��"�_fv���kz_V�c��Y�]u�w�'r��87��N�k��2���VIj�t�����=�b���@�������'�9��f�R��/��"�sn������Ɲf�v:L�d�yt����Cz�jU���:� 0K+l7��F�7 D�1_�uo]�\W�����G2�PX����S\� ����jj;��@��l�����hLhe���J��m����KQ�*_T��&��-���h#��&�ɗ�y��RW��rN����AJe%������  ��i���o��ˇ����I֐�u,S�e����:�ۮ�n$%�� S�훸e��=����o��y}F�)�(3a&�f5�$�cR�<{���v���(���:�;��i�W���uɛ��#	��ç�m���E��p�oT�(��ڕׯsϮ�N�U89��;��w���#��x��o]mJyd"fWc(�������e�yvL℁3��|���U*����ϝ*5z�'�̎���+��4w��egn���r	��#��8�Rx�9oYUɺ���\OI<�ݛ����I�=F�b�9e�����GzkO�j�
h�-�+��4�l�2�I�	�:��6����Q\�xQ�=��FP��(�<�O�q�u�e̵P)7�0=Vػ��݊`�`�f�h��ׯZu��b!�����9]mYC�}��٘E��TF��sr:�mY�M��i�m���##w��S�8�|40���)������ӿ~ן���jȱ��Z�D�ڣl�eH���F%-D
�֋"Ŷ���X)U
�*,*,�X�Z���Z6�XҶ��ԬD��Pe�KJ��
�eEQh�,J�,�U��iZ��(QZ�Q�+%�F�*�-X�U�+6�YP��[Z���aD�h�(�T���ѩPikm��m��5)m��IKB�����YR�T4*�4�TJł%���Q�#
�"��µEdR�k-UkVШ��K+U+-������Z�U�+F(,V�T���V	[F,*V�#i�ZځD���@R�ڪ�
TP�VPU�QV���m�cl�,jڢ)Z�(6� �FH�kF"�YEAU��-��[b�Ad�R���T+%E�R6��EXڵRQ��[QDTF)Z�����^dF�:t
B�q�{9I���+�_E�l��5n v�7{F�%�&՚A�S��ƨ1eN�^M����}�ˌ~[�{î�m����XL��ю��`�f��$#R�,�}*Cĝ�2@x�eC��7�,)ے��S�$�u�7��.���헩P..6����񣔡���x7�.;=q�b���\�^����w�m�ꮜ�]t��:�9�	�,׃����z��@�pkV:������R�`�>4��v�a�yo8�ftE
�@�Ӆ��yW���=J�o�
���>/-���J[w϶��_v������Up3Ó��P�&�S��Qt&���r��3L�����u�};2˾xD����mL�c����r�,�xZ�!�f�v=��}�('���X�\�P�'gՙgr[ͣ�xQ��jWK��b�{#C�6��}^�PT�wKVq�s��D�rkY��,��lԣ�}�����c6t�."���b\�F���!���uH��%�9㼇��/�"�*Y��K���[]A��e��,�����]m�m��QSFr:�p��ni��<�s�K���wA?^�K�h���J���k�w-�������œ��H�v����N��8in�d��s�t2�H����w���S�mGGmB�eRFpn)�(RJ�b������ϓ�AQ�zf��e�l桛TNrF�h_Vm"�W�B�<�]�����ԈuF��#G�A�����}�QH�7x�m>Ş�&�|�L�Ꮀ�{,�t�8�|�tVz�3��^E?��JBR:�n �ә~���~�qA�z4/\J��7.W��<o鳽����P�{�r�Xr�
���j���O5�	�E! �`ub�C��<�k)��tDإ�\kvNW+lڟU���]�՚�.*bR�@ߡ�8����Mv�;�{��=Z�v�!��׸���5E��������c�Y<
��)�T��2��	�;��Z�F�(�WS��U�j*�=�ʁ�2��)��� =�����W��<��r�(�H�Aq���P��!E��l�Yo`x���fZ���G��֧4�]鼷H܈����L
�]{��l��1ȭ�:����}�e��1I�yF�^UV�4t�'ZdXV횸C�u`1s>�x�)M��Bܬ��ٸ����^-X�+_
S��Äә�H�kn�5X��i���2�^<�~�2B槊����Q�0lV��ׅ����xez+�ZIxn�C��V��q�-�"�6�禜.T��n!�p9R�n+�62�Q�L�7v4̏��,�q:�Ưj�Xа#�4�0_yc�֕��_u5jۅ1��vwT�f�SVm�!sm��G]FX�+{,XPۨ�k��׮
Okw2� ����)/���6��Vi(���l�9Nk1��,�0-yt���J̔�JT%i��2�߾�_����m���ׁ�{�!6���m��ׅ�����S�c-@kQ"�Jv�}JU��n�r>����YT'5i�C h�iCk.�u���ևE�m��q��qY�u�{�܂�$�uDEN�Ą�wt�ld��י��,�G�5x+~��KN��hr�#�ߣgϕ����e�1P��+:��ٴ,��/R��K�;�q��ˊ{Ӛ�v	����/[��G\�a�����.�a���ڮ��$5�v�Ƶ�U���N����4��y�o�qޞ��l�U����l�\��+nWCܦ�W���B��qՏq�ܼ�*b�
436����Ό(�bxз$��d�b�Bq�0P�Y��4A���r�G����jp�j�b�t:ģKb�<�Έf��~���(�[z޿I#O���g,�c�����'���b���5���]�A��Ϲ�(]��D���������ks6�K6Eb���TOz�ŜEMO u�}�1ءal������dF���|譺�^u���tg�����*kQ�O5Ԡv���辳�}F��:T5k=Bܒ+��R[��p6�e`��:�{����f7=�{ܡ�R�;���e\Y�h��sg%���q̗��h���
����B/'b�o���E��s�2�:K�=���XF�[��\<s�k;�b��6�'�.�t���G �9��p��n�a���V��:O����3��bAuV��:�	3U!.�ׅ�<x_�B��-���5�>"dX��=�I�\�S��@��R��(Qϥ�|9�R�҈ϗ(�X�s�d=bx��Vv]t�"��T��BI��)��0��XVH�k�L@���/�o�Ur
a��IV��)���\�����d��KQ��fvXk�5{�hL��H�B��@M/̗�{̄��>(�^������ܱ����/uw����O�,�9X6Y���:�y�/����T	�o\A��̛�^.B�G�����߫4�i�yT�T��21��\�7z�D���L��vo��pQ��SΜ����`���C�Ű嵁��?ߩՊ����h\TR����C��*t�+�x�yN{.j����k��>�/+<*�ѡhO�^��424�`LrO�_���+��vΩ�VSa$Q��v�j]��s��[/(�$c:�W$����� ��K�}g�gs����w;�,=��u�W��9wK�,.Bm>:c�̷�	Τ�vV�*���t�	��z��x��R�G9Px��"N|�WkG�s���z�]��6��8���0�Ӎ`�R��R;jnҡ=��/-�ٺz�u:���N^'��4ً�T=柽.c�d׾<���zbۨf�Nr�b(s)�<���42�Ջ�j����y٠��J��;;��[T��uŸ�Y����+o�8�j��R� �3�%Tp����(��V-\����0fo{��	�S�Lj�R�z��tέ�>��6��*��<g6%
�R�&!WU�Wo,̀p��N�0�q$�h�@G�.���*z�oT��Yk�B�7$"5�]���n��[�긮`���m ��Ԃ�N���"���ƥ����X:��A�nS�'�
�@ξݮ�y��z�fV��ci�kB50�$�-�S�� 5�=
�xb:,�*fn�b��ƅ�%�Q��v͖�t����������az�=�sV������=*EȎ��g�S�-�=d�{�!��ʨ{y�:��X�q��5B@K�]�$9ڞ.�?N�{���^��U�����ˡ�jW�)����KӋ��"�fV�fV�������C�t&qmA �8�2�OA����ƶ���l]msYɶ������5��fK)/xl���9�����.p�s���E��m�Ù�A
�������\=��0(󻭡`�ػ�H��[���[]�=m���}�9s3y���+�͙��U��4��X�����y�oHQ�ϔ�h��������=��'E�	k�w;gkg]�F���/<��98�`���2Pϰ�^����&��������%f�8�K���m�u/I�Խ��,�#��8�,�/�xl��;ӂa7�����%�j[֛�:I�5��f�2U�ё���b��a_#��0U����^�\��#�ٕI�n����k/A{�����Eź�l��5��G�K����L�&�>�o�f5��<�ز\�W7V�WB��X��ڂ�gZ�����nG���͐n�돒Jf�u
�ɛ��fݾ������\i)	h��*#qJ8�Α����6#cux�_m�����ۆ�����#��ދ�#�.2��J�V�w��q&�ˢf�'��^g;:�ޡ[��=Z|�p�q�e�e�o�h�ka�6{j*�.Ԣ�G������v�9[�/<���5Sc��փB9\q+Q���8w�v�n�u�9��-x�e��x���lEYc<��v|sU���h���N|d��!l���:+F�����g��{�{I���=��tk:vM�.�ۣOp�ٯ/����f��$��wG��0���r�P���!��HW@� �����x���+��Klwo��+�Hs�����z;3�fvN��И��+qoo�n�Vv���|��{�w���Z�GƘ\g�"���z�(Wo�(���_.O�k� }�MG	���Un�'�N�Ȱ���̐Ǝ̋�wt�k�'X��u��G����-��o۳Ut6+��m��u:���u���X���������t��0y���u�Ǐ���<n���I=�(v���xOV�,����=}�t�-A�8��ӇQL����MxZ.e��������=6��mV(�n�i&�>��u���hmSp��֬�s��R!}���u[̼�/侖X���u{Z�=z��nu<��+:tW2c�D*�S
���N�2S�k�� o>��&F{Q�yɝ���.�*��I��4xܖ\)��j�q7�V0w{Y��A�Y�A��b��ܩx�C�u�=����*��uHG0hz��Tf|��\rG�4L��T����;~�脼������0�՚%�ܞELa���C�\ Gd&cA�EyWk��������D;�*Xr�MN�+X�����1��Tek���ݕJ_!t���n��g���'ە�J�g>�w�3����ʹ��W`�J[17�Am v�s�R�&o�.ZS�]�f��{��7O�O���Y�e4"خ6:�#�/���:�
�#l�>��V�=9�a��ߌ�g!`S.�X�ilX�UgFL����;.TGM{��_=�v���5鴯��g���q�o!4D�u�,�4!�L��^�|�i��-�NEu�g�g�y}[�q��S�u.]aCD;�ֲ�m#()�����t��׭P�!���#A����2���Z�{�̗�벉�*��ǯ�C��:/��׶�2�S9q�ګ2,)ŮKT't<���͎Ae�9~�f��4 ��@R����2�����l���^:��f��O��I�ٱ:=���j�^�L2{,w������Y|�?uoƸ[,�psB��r����&�#�ua�M{���[�3.t��V{KwBWr�*�G���K���0�[z����FE�;p��V���N��nİ�)]��4m�]%���U�xX�̩i��� ���<Z�(��f|h�^0P�Z`=_p�*q~eP��[118���.{�7Z-u����]cW ���kb]�}tJ���X��Ni\�B����0ifٵ�#9�V�j�M�l<�� j�`��wL�����.D��D5���2�,$�Lve՝&!c�,��*�!5l<��]�sy�Ra.����R�i��L����=@r���L�I�,x��D�cRa=+h�i�����SX�o-R��1.�U��N���\�\PFX��L�Gx��N-~���雓bGMc%y^�����m�]<5^�p1��(p>9�.cb���&qR�����^��37���_(�;'NՁ,��f�����g��ѡhO��`�l�Kή;�mpbG�N�)c�OT�x7�}��9k->���7��éԴ
=ܒ�y��q����K�� �� �si_�G>�v��	GyF�˰�uJ4�Aa�"1Y��V��u
���x�Q���GR����Rժ�#.���s��љ�$�4'�7��'j#hW�c���܊sC�]tB65N8�5�:�>�?L��(�k��/e񭙷:�l�5�@�Z���i$�5�5=�:S[1L���dU�ex����=/�Wk���T�y�m��3HP��Ԩ�e\�|<�Ý�6�ga��(����}�r`>vD�hU�J����n�!e����Yڄ���1`�S��p�II:�2�o��5�Qz���Y9WǃB��gkE���
�]h)�c���gK�5>�L=+_40�9P��v��]�(�p=���;DX��d��+T�V9��.�p�1��5Ѕǂ�kR�K���XP�g	@�������v��C�5��b���`�EҖD^U,�*3A_3�Y�]����x����[7�Z]ܲ˾vg��8��0�P�O*�=�NDM�s�)��]�Fר���0Ǻ�1m0���x�rG1=]=7JFMz��yt=���j��vS� <k��KӋ��_r�s9䬧�ܺSfa� ��g����qV�<g�^ZݯY�����2�ќ���>3z6�ڵ�Ovܫ�n!��+�z �Ђ�r��e������5�4�i��u��� l���˪��t3۝�KǭY�YG�3�"��fñ3�n:�yR���b->u����w�*�v�х:p�&�Yu�����z�S�K��t����1pV�n���
/��p�f�j�.�U�����������e#<��g��.�z���=j]�5�(W� L�jX_{z�|���|В�@@��N�<oT������<�^�XF|գ���U�%[S�|ٮc�f�t�v������F�i>m����BS����\�}��9�*�>)m�h�]n����-_��C�F޶f�ʷ��ϸ�5�t��ՒKY@�U�1g6�:�b���oN˥�x��W���
Xm*v���皥�-�ͫȍ����:���t���X���f�Ǵ6�\���)���,n���u��h��`R�S�e�F���#�˭����uh]h\���b�>f��s ͢������Qh]�����;�:���ܺ����$���w4�r]�E@]��qU��f��;
ˤ�`����㛅�H�_;�glڜ#�;j�=��*�զ�IP޴�O���1�9/�QJ�C��ѽ� �f�� �׻ÆB��y��Md�F/p��<��cQm@�%��ۻʄ�:��C��]��WD���eS����ΦdC^�f�J�S�[}V����ANwF��SI#kv�^t�Z'����.�⭥EW*8d��Ak\�w@��ﳷ���9��UɊ��w-0`�3��`����j��gc��^lsL�I:0��&ϓT��xCO���V��տu3]]]����E3�r��Gws9�*E�f�W�hV-�.��n:��R�֖��D�C��꠆N����c0���P�o�5��i`9QvF�"���@��[ǧ�j��r����d��L|V��6�y�C0�����wӣ��Ah;3�R���h���T3�m�)�.�Z̲k�Z/�U|�_9&�ϵi�+V�e��4pKU۝&f����`�,rYӟZP��t$��O�Ied���il�e#[k)XRn˔���vm�W ycU�����yݲn�eI�Hk"�׆�4�\U�kxJhx�T ��σ�����,�Ö��O��+��e�#J�ȴI�V:_l��0Ô��YX*��L�7����B��7�WZc+.��5nRʏ[�ס�o�;]ɒ_��ȧ���m���N��<�]p��y�L�!���Z���SHfD,U�A�����V�峹V�ۻ������DhA�akR�:j��s��Wx�l]&�:�a
��ج;J�Nj)�(B�Qۘ-S����A��.��m;�0M$�����
�o������[���Ժ�HT�I�;c�۴>�v��{+�&��p��ܺ]��6��J�a��Y�����g����͙�#d1��.�����ѯ�s�i��j�e�3ջ6�e�5�3�T:µttβˇ�dA�9���2��YV8��Va�h�o��X�imYʐ����Y�TE!$F��]7%뉛��(;)��e���"�.\-KYt��BI,c
���a���L:�x�˸Xw�_��PiArИ�E��l��x�f�X�sS���<�Ӂۻu����6��&Uݖ">s3-`�	)ҬIb�J�#����,`�*��T-�Z�X�-�Xڱk=q9E-̘$��DR,QX[
�"��V�q���"V��Z��[�-�"�nY1U`Җ2�`�ZȦ5PX"�cĨ�*�Z��( ����+\�0�*Kl���dY"�TQR�F(�mDeAQQUJ�PPYB�U��2�X�
�EƱ�e�� )P*��
�b[DR��Ԣ1�e�TP����*UE�
����R�PEV"��*VUV,b(XQ��3�-�"���((��FL+J����P*1�*-lU��cmEX���VEdD�b��DJ�6�-�j�X���`�R�dV"�R85TDV0\KJ֪�Q-m2ڌVZ�V���������T@F*�,��h�UQ��hQK`��$�L@������j�&o�Dݬ�D����sFIw�B݃R{RdI������3�&���v�1���/�f��)%�ж�l<�.�j<_f����C�Q���_�i�&pO���>J��Y/e�8%�~��&��ƼS0:�R��4�:E����:B*�́��5���bm談��Ÿ�Xq�|Ҹ�����i���4+ǳi�3�9
���g�uxi;pS�62��O���85�k{W�it�8�������T�U2aݬ��k`L��R��}y=~Y�C�|��)z|�>�ZQ�i��S˭���;%�?ks��5T�l�����ا4����(Ԉ�0���J���m�Q�p��?wE�Px�����|&�-r���&'����P��i�a]#6�Td��l��,+�hew[F��%
�]-&��H��C�v1�S�>�!T2P�_u"��uX�>�]�/M�����x�g��xA�֖�yO��^�Ʈ�O\Xq����J��>����T��ꗛ�F?���ų�b�;/�{�pW���n���]L��}�4��t�&�R���v���C��"3����K�sX�[F�ZP��]��?���V5��J�C����d�ŷ2X+.���
�
Y2��<ng��9v<D�}c,�a0�8ȯ!�{V�>�K��֢��c�a7VP���{z ?vl|%fD_կu�N�O:m��(�1�5 �Lp����o������~ʾ�!WuL(xN���<�$�Z�k�7���fo�]���o��֧��7��L�orQqaVCU;�{"��[[�X9�t���o��ބ-��栱eY�!���.��Z�7��_��:�\8�;3PȬ��VF�U�c����[��K��9|_��8=�����m`lOS��:E�f+�'
)Wk"j�Y��F.Ȟ��wie��>�>��)�6��Ȱ���K��SԴ?����p+]�1<C�8P��a�̝;j_���t��l"��H����	SGB<w�ꕵ���,e��g���iN�r ����>�������募5FDP���ڰjw$�Z������zU�[H��uHÊp�T�dW�J��]PeL�v/>������E`�*W>����G{ۛ��*%������*�nzm�8.�OE��J���f�֛�٤�˩���	��y�.��kZ,n�$"�Y��g.���V�2]�>X4NJx���(���^��t�+�	S��6wom�,��g�>��} ̠�B�f��ٱ����.Ӿ�7�С�H�e���/pPs�O���toEaR�����a��O���]f�����駏)rqe�"�4u�C��������ѝЉ�]���<�D▽���5A��ɨ��;M�;^��=k�E�T���8�T"��+`Ǚ�{[�D��y�0�Z�1l"V�r��S�� ��~��-V|�Dh(��ѓ	���n>�Ĵ�#�I3�]��
"b���4m�[j���gè<K,xΧ�m��j61r�w�������	�+�d�Z`.��H�U2�"Vl��3���۽Z=�;���w�&�`V{�ٔ���|�xa���뽩�χ(q*N,x��f�����=6c�n�yDr�����,����2����{����4�{]�Η~ǌ�Ofө�1o;����f����_\-'��汬�z8p�]AT��U�,`����ç���)w�_^�m>Z֡�a�VT�p.�e�Y�w�k3=o��VUi�hG���~۽*��2:j�fq'v8�0�.;C��W�y��]1Qּ*qk�a�m�c�M�ц�I��0O[��\�ϳ�����5IR�*�)���p��M�*�B2,��߈5��Gs�%D��t���˜=kKX�a�n�@xl���_n���
�Y�=��_S�:�zZvG�����=��{�7=$��ΰ2�r�7�OT��=/9ձ3]��|�v\ȷV�p��� ���H��c	y܂��2�y����ꜥ��ӪS���!(z��,ͧ�q�x?���fr��ţ��}s��C4z�u��cV�5�}W���-#�ч��������
�C�J��F��8���:��\K��D���ZO���{Y�f�����@�B"t��I>	w�hqN��ֺ�9���.����I/0�����o���.��v���JO�eB�	�>4�V�AǢ��0����c>9=���n��r�w_7���2�9�^t�x�W���F�9�L{��k�
ebZ=R��V*<>�zuA��qW��f���Y~F��^1,��XSS���U�xWJD x��̮~��z�W�g��S�Z	�\N£��{kM@ↅ�l�U�N�(p��B��^p_�}���s���y��EY��3<(�,��~Mm{��-J�E>p49ʴ����Ϲ�e^�������� VBF!+A�+��O���!�lC���bӽg^s���R�L��]���-ٲ��V-���kÈ�Ƕ�[g.�|0J���2��gϧ���r�3G����օ^��C_5�Uq*��oY�5�
�&����"t2��3fm�&1�v�&a a`G	�ts;u뗡v5#{��Y��pD��)��s�l��]����n�1i2<�:�l���"�\`̈�����$ޗwݘ��Zq��*f���\�T��su��8�"tY���L�#�����ˎ�U{עj�r�t����z��b�t�M�.�N�Mt�>�O�.#��ش�x-|�t���:�zv���5���Z=�a���j��f�b�VD�p��������[�gt���"0�[au'[�p�����f��e�~��}��>��n�t��8E�ϫ�d�2U���1{�5�5�6�<7�e�9��V	z��,R8�)�@b�C��"�a���S$ݽ�}�3u^�a���7����O��N��i�H�>�C���7��r	ם��E�~�f����s���(�h���Hߥ�@�'H�a�pеT��y�z�V�Ck%<};im�)��p��Yk���yq��؎q���P�Ac��i���^L�#܂���]����m�t��B����r��r����*�n��~�D��H}�N^ �eV1�-���r�Vr���n�&��`����p�`��>\�zss�d�:):�#u݇j��
�-�B���Te��ؘ���oN�o�;sf�/�Tk�e寳��<F���D����Lr�,/B�_^��b�E�r�Ы8��˞�� ��-�o[��J��z��8������<g�[��tc`*]f�Cʀ�rt�J*<:\�a i�:4�=B^]M����W�@^R����z �!U��*�E\�n����ݜ"��`��{�g'C�V�������se���KoI��J����+�X�A�]��q�[��t֒��c>9�b7\R��)X�Yk:�(��j�����P�j5e�
��V��@V�k�=Ẏ�3�v�����0�$����H��P��˼\��g�Zͭ���D��=;�q-Or�,_M���G���e�RK�UDE���efS����Z�&�@�Q|�:�ޛ��wy�y��/��U�tx���=�A���+v~�z�� �(��{����ٌ;ӝKrʁ��u�Z;חvb�#{�T��8`�͔TZ�,��}��^<���kQK�Iu�kcUo=%o��������_�ԫDG�V��&c��ET���S;�Q*�᳥��k8�WB{f�+æ�n+60J�8,L�ƭ��n	K�ћ3S�����M�rS�z��4���m�ԧk�dCTˡ��F�ŉ�Vtd�8o�jʕ8|�o���GP��6�9�����)�Ejm-ա�/�uY�r��m@�c���c�Ӱ�Ȼ6o���\�Mǭ�m���J�x��À	��:	���}h:g9%J�yINY�LL�1��Kg>�)q1�pm�VD���C���.r\B��Q�(U��*="qo2ߵhJ$!�r��3٣QV[�,o7����r��+�7�)yN>�R��C��͔] ��lY����/#�̓�Ù�<�zS>s���>��S�����H؞�p�
S�']yE�v>���D�!�uy'\�hǽ�F�g_�_�Z�0���EY^mz˕��*�2p����/*�%=�dxެSKY��S�Ԯ��0ZufE�=P�����^%O�A��n�����\�z��P9��:+��蒙 ���y���js���p�M��E�;U���Ss�6ۗ}mD��ܖ�L5�X֋��\^r�^��N��J����ˑt��{������w<Ϋƒj�s讔pEqcIB��Y��YЩ�E��rb�9&%ժih��ܝ���0���M<�<5��y�t=�Ȧ�^(��Y<�jy3�P�Z܊�U&�2�Y�fߤ�+�۬�*L��v�F6�w�n���dnmR�F8b�.��ޒ�P�n�l#9��Uv����h�+C��N�"thS�w쬴3"�44��:������]��H��Q�w���͖4��y��>�x�O�qFL]`WmǯN$��\c;��x��Q��GՍ\ݮ���.CW��rȹ�o��\Ѱ�=����V��������_�vnq�au~��a���y�`��N�u����w�.��P���~�,w+a��P�����b�=P�^�f���u���Ւ��D�����/rL��D�y�������y����N��8|�>:�3�l!�;</yl�+L)Owq�%c�|#��0V�3��3ܜզ��e?}�z���?1��;/����e���`6&7"��<hZ���s�/�\�f���T��(电kG�L�o��w� xM\��KM�fصS���"���Ӊ�J�!Qn1�9��>9��2d�5n'�B��K��<VCv�0Ј����O�����5����]5�Q��o kXJiFa��Wy�9����ʇP�)�fM!�0�Kqi���(�\y���jt����v��E?UӈҎ۞+���v(ߩ�7-HQ	��L��N��	��-^�����u���9Z�eB��!׏�£µʇ�V�\��p�E��vj�+ٝ]��26��n:~��ϸ�秅쾬�mU�{����[�Z*:ߡ�r՛p�%<`rq�SɊ��̕y���Ā����ۑ�>Z��旎�F��\�=m��sg`јe�bV�l\+�e��H�&��JYf�!�D&!-��=��x�x�"�G'k@w�fhb��oS�Y��:�
��+�T>~C����Ӭ�&w�\�0C��s��5�	v�������^�B+�ˡ�W��24U�*��C+3�L��)�^�=0��+hxO��u�+o��Ө�/Ʈ�*�� �uzlhl֗eIyt^�֪��4g��Ү���d�Qό��5�����O��8�k��Dً�w��T�ۜ��8l�t�.������}`��9Qz�y�c¯�X,N;�h�xiZ���*�Yz7`ڸ�/jP5������2:8��Ucs���x�ʩ����n��z�s���Y��
�U=ע���\b^�p��*�`Mʇ29姾�+�W^����rE�/t/�;x��۲�nt&���m*��J���ϒ���|c��d�/���z)���������Y�]]���R��Մ���!�A�Uk�|K����!<j�w���
7/)�W݇�{z�����#V:�lJ2�)�8"��#OJ�A]�*��w��ދ4ѭ��Y4�yzyV<]�H�r�_<1	u��H&A�F�E�Wvy�6�����7���O����Z01[㨥z���nyⴧ Q�E���枴 Ӷ*uY����nST��e�kB��XK�6�B,6�*|�"�ն��gT�vL��:صm���鶸y�~3/��T'��%�1�o�j���\�qP!�/ec8����6[Ɔ,���\j,(���+��dr郚�͸�����-q��!�;h:��;D_i�>���k\ḏ�Λ�����!X��6�y�p�I�U�^9F�EY
Ղ�g�����䮅O}f^�(�zj �����=[O6G�0�ٚ�E�.4]]��
�Z�\gl��-#y^��v����k�Uq��)��%\)�<1ÇJ�?vo��!���#{39�r������;�at8S�K���Ç�[zNF������<�P���ꥵu��W>���РQޡ!>�Z
�Yk���.�]�
��������}؛�U��~E�E>��ŕ�@9ݰP�R�ϧ5������,�I�*ތ�I��'Wk�3J�W(l�z��3qن�D�����E{�9����X!�}���q{����L�D�.)+"���ə}x��9��9ٕ�S��e8X��	����ZiX��ů f��n�]4��ۺ2��8м[��Y|=�L[(�U7��]E7+%���:DȓX6j�p[;疬�ەp&��}�*�;V�[(��V�὜�������s�;��]�V���m�U�l�����G��ռ��r��=XBT5[a�1��&P�i���Che)�
����f���]Bs�V��N
���ջj�V%D�n����Q��K�`�5�oł/�h㷨f讧'�-Ttt���Y�~FQ�M��:���#C1\WU�sY���Q��N<���]�51�31�M[��g+��[�{`�-�c���)>�GۃU>�4�Qi��1��,�r��u6N�t�a�(�ʇ-t P�]��<�V��9�r���cA⌷���J��J�-z����+�����ܞ�A{�Ш�+4��<GY�=�w`��4�u�k�M>��D�������qU�]lfl�ly8�1#b�W[���ق��cM*be������C;MK�ry]N�Γ'Z[ _["�;�Xv��f��k4	ص�_P3$X���.{�gr�Դ��ѧ����C_@�޴�vl6���W>b��B�Y׮�d�p�v��[;��6��|�w�"!Q�gf��6;Z�t���Lb�]�Hc��Ih�:):�N�h֊��4V����M�*�M��zk�5Ƞ�X�c!���.���yq��)z�0�{"~\���<N��<�z�V���%�U�y������ނ�S7�%���y0�Λ�P�D/�J�nV�"s�Ev3"�Z�Z��/B�qI�� A������J�͋�S��]�*�>��0��D�A9%�x|���B�A2�d�yۦu�5L�ݽl��PC
2��X�8wq�x��@�5f�ڋ̏��wG���v���R�m��J���`������n�$�Et��9Fp�evw+]�9sU�:0.��D�+��ep�!Ն���b�Ҵ�md�=G6�oV�.�׈�I�*�.U�P��uЛI����*����sAo��w*��`��&o���|(�s5��HTe�"�U_>�y�n��[}Hd�u4����U���7�l���1Ӟ��a�vqj��!�t(�kl��"��0
2]�L�]�	��d(����:M.!X����`Wt�p�n���-��#%5i3�d�wj����U�ׇ+L4�+�7;�<5Ҋ���:o׸J�$�����H�sBZr���#���yq!�0�<GS���Ѷ�Z�nf�¡�s!Y��X��o�����qcT�O�b��Z*����-3��"�I^�Ĺ.�&EԬ�O')�i*�a�%�WA�.VJ4k*	+��0J�\�͓B]����;D��3d�����뱖��Tp�1i�r�0�v&�����6�z�@+7�Ã[dV7��:�ֵ��㪳X������V-�TR�D����*�m�L�,%�[eE*e��V�\��T�Ҷ�T��TĨ��PKlb��
"
c1��1E1�D��UD�DL-B�U1���� �T���6�(bfS��F�e��Q�V�\Lʪ����(�(�m�L��cmB�hY�%F�Ub�����R�+n3¨*ֆZ��(�bX���,r�����dDC-T��
�"�c2�ʱjW-QQUq��j�hԢ�2��(���U�&+�����ֱ�Ub��XTFc�X*9j8[��m-��mDƖʋ-��UER����(������S+PKlUU���f`���33r�F("2�8�T���P���-̵��#Z�زۖ�-�`ܳ�8&ap�c�Q�-R�B�Eˉ��T�,E�����a��be� �5�j�YYJ[��\���kiX��jb9r8�Q��q�bS&\G(uf�/Mv�x�:�(ճ�Ӷ�
���H�˵P`��V��{s�+;��ee%M+�{a�G�7�����}��t��\�JA����_ye��S��&q�0���<�\^=1{��-�'���Qչ���\�b����׵��y�w�<�9���Oz4��F�{���3�d�<�����ٗ��v�خ��W0��Y҃�^ɕVt�1V�9���4�zGN�6ؖ%��}������_G��Xy�|o_T��0V
KÝ\�`}�R�82��&�E}u��bs{n�e��4^t�V��+�Q�R�K�9�xt��9��|��U���$�U��.�36��^�U���y�X
Q���*.3=>"�>����1�/6��3��+�:�M]z����D��g��l?gʼ�>�)[�Q;��蔼�������n�+�<Bt�.����ګ*�ZufmHf'�jF��$��=�/�Qݰ�����zΏ'���j�w��s�G��U�$o)T���\]��_κ�9���_(ũavb�u����q�9b�tۧC�(*�Cs6P�$ ���^tj���uu\`����3�'�k��Ҩ�};*f�D�+�v"r;Y�C����p!�'��Z0߅j��ݚ��$x���ʺ�R�޴_�]SM,af��ӷt:����[bJ�@%]�d�J���ӭ�:��$�Y��^'��ډݏ;{�򴎜�ӥn`���59v�R�gJ��n�z���{*ڀ����r��`�P�ǥWT�܇�Llq�F���_:�>��ӫ0�k�a��8�Un ц�xXL�D�L��_N/̭�h+�t�{s����]���Y��[�/�>V<�JE��<7����Q�z\ޫ+�b%ʺ��/#�z|��<js���$W3����y:*���A�Y2��qn��qiE8���-�݊U`'��y
�9�lX�<@,��D/�|1휘Ӷ�:S�B���	�ͦ��;�k� _@�4z�PJ������\fx����`�+KJǞ�=H<�G"��onN�MA�;AL\ Y�'�{=���C����S��К�E\)�ΚI��քzk;0�o^>�t��`��׭�*�Yq�"ʰ������5m�;�8�m�I������Y��(],�B4k-W�<5�ډq����G��Њ�+o�1�6Q�P�/+6�}�+ԧs��L;��-�<�E���%��#����޴���-/�<���j�}]��h3�:��y���ܫ$���Z�l��N�����
 ]`[�Kz�ɦ�WJ�f�#�j�xRw�{T�|���	A�춡�����zVR�s��(�֎5�c�Cx k��qa�����*Ζ��0��XO�U��6f:qq����e��>2���X��	0z�����־jVxkǙ��A)���=�%�$�z�W���}�SV$}�]fT,КC���^�*-6h���Do�߼����sg�$<6�w����ˎ��P�=�G�(l����(X�Լ�C�U ��sH�6����j�N蝭5p�Zg
!��X/�[*"~
��p�JaR�j�4%T�Fk�ֺɓ6]�ý��Z}ZթQ١�|hyk�
����UB�(�t����`�aQ{�u��4Ivׂ{��S�!⮋�W)O��q�𩆗�!;� ��NzC��n���h,̷g�������3��U��(��_�p�<�eV[u��c{r�J��1��m,��U�S�WX6��#�M������z�{���--���Bz��39��g$r�k?!�;�ua�l�R�[�t�2��g��Q��wo�$w�_wL�c�mx?���I��e�r��yӁ9��r���,U�7�Ihb�g�ҝ����O,�h�w��_N�S���w��_8�q�-XO0��"��գ%sֶ�}��&[:dW{���g]\y�7h�j����d�m�>�r�̾霧,�U�y6��*�-����	��ӣX��EΧ���]]��ds�!d6��9����%�ѯ6f�XDH�
��}��k��l���K.�d��]<�z�U٫��q��IJ�ɡ٘���u(��:c(&�Mv�HO�A|:�[��2�W�u��q�F�[@��s;���F�ui��Nz6��5��/���.�:3L�#ӎ_��������ĞI�m1��f�K* e�{��j�>�p�H�f�P�F��2G�,b�:��][��m�Ӂ��Jk�z��\d2�K<�
��ي�2�̠kН#���br��~ky~�w�y�^���W�艢a�|�����+��FooK�.F�4����``���t�M��b��M�><�9����t��r���V)u��MӔjDUG�0ax�i�{�]��kp�n�����v�<��|c���9HY���/Ci/x��J�32���זtџWq�,{\)��dJt��^��Ԧt\�υO^U�5	���{��FX��3���2k#�
j��`\ׂ�l��P����������:9V�D�tVQق{�r;�b�������v���"��p3HR�����c�-�-T������m�m�LvV<z�<\�q�b��3ƍl5f��b��9ͺ]o�=7���N #(U��3i����eN��oqr.��撚)wSq\�)]��t���.P&�:�J�|$/U*Qc��GI�!X�dj�H1�@���os�����+�qt�Z��"Glo)el氢_��D/��>yR�d����k�k0����fˮ�Qc�h�8Yb�ۜأ}�d��+���y�z����;׏]�f�}km$x�D���W�R�{:���/��靣�;~���U[�6�Ѝ��kr+ N�ek���C��.�����������6]�(l�5T�݄�w���ڳ~NqwJ��hi����=��cݼ˶�9�U�>��SL�8�Gw��턼w��N����8�b���^��zp�<U���f*��8��8y�q]��T��My�P����J��]��Y�cP�ڋ �="z�#��ZS�-9E�R6��wE�s��Y��.xtFWl����-8#O��r�Qr]hQӡ�WZ��.vp����{��pҫ`�m�f�~�{�a
����:�P����7�R��鋄�vrWM�󇘦u`܄��s˿T�n�y�Z�-z����م���8̌K�F�dm�t�����	{f|��-�q7����*�>pS�I^˥�W�(�
���4�g4n*���X��wf�	��%�N������;t�; T9��S�f2zNښܺ�(d|�"��ݗ�v��xj��w��G�CM�0���f�W��3t�Ms�ܰ��gQ�nw��J�Xj�g:.k�2�<k��C��a5�c�d��~���������q^���s�=1j��9��ۻ���X����&�;U�x>a�e�
�ypn����Ε�O'��Y^�E4����"��2T��s�	���M���Бyim>�̴�U�!�Ϛ�,z�^�L�������B����Z*�8ՕY�W�}yU�����޻+l�V�Ɯ*/����!�_+�3E�Yr#�QR�"�Z�De�ra����������ׇiI�[{x���a�4���3���a��[���U��vQ�-CiV�c��J%?�_��Õ�_��׎��xe�!��8��s�H�&r��b���dp��{)[�y�lN�=�ň%g���ʬ�ao�=�C���}n��w�#���m�#+ܝJ��{ s5�n)B�É�lr�3b��uW�ȝ�Da_���9�
�p��؝�W[Yy.D��Fb���bPʻ�5%�C�����A�V�n�?�EkI۵5NNLu{�l�K[O���uO)Q�� ��q3�n�/���}42��R=���t�&-
�YGLS\x`b�<7��Ժ2>[ٽ�)�9s��r�^��j)Lwa�Ƿ��]*`�d���ⴉ�>��\s��&u�u��^K&��^��#�\������^�W:4/��[�U�e�CzE�~S�P�����s�"�S\�j�ؾ{�u�U5����f���A��px}�%�FT�}4hZx��[�s=Q7D�_'�b���}��/��.I�0���B�ޡ`��t1kĴ���s�w��7�h���z�,��t��ҘJ��S޴p9u��kK�hÂ"t���a.>����/`+B-��oc��Kolt¥/i�z�=<�5�e*��CG�|�r��\|��M1�M�-��[5�xښ� �g�҆��[�Ze���	��}Q�B�P櫡Ѩ�Au�E,����o��g8�`���@k��lv���S6<�}. ư�p�	�&	�A;�w\�<ϧ��=��k�����3��8���5ACe?��	z/��(��Ы+t��;�N�����k�|á�*�;\�z�*1n��Њ�W/Z-x�ԹQ����U�fӗ�JY�b\�p���gc�|u�Ͼ%V�.��Vc��j�N��U�-=EL�&�w*�]H�8;��)�&�s�X)wl��BJa�~�����X��W�7��;nRU�|��g+�$�|X���GFWP�\�;@�-[��H�nZ��0�C���x0!����>�Kl�FQ|�U�%�¸��++Őc�R05��W� [:f(K,�
r��a�7|r!ι�G�xV`�������\��}��^�(��0b쁣qCiN+���(�Y�BF�ߚ{kh�UF�uo76�U�nN��rV��S67&��C�}�o��;�4�C��C{����e严k4�:-���0��؍6X�U���(�l���6��H��_M
�c���h��G]_��_�:�gLB�L�Đڟ��Ұ�맠���]*ȋe�ɒ�9�|,�nN�)�a���_)�O�]��B���|�$�"��l�t��P�R��WZ4�4�IR�2�뙄x�l�i�6V������5��/	�"i	􂙁�<*�w=UTᕹ���ۓ�q-&�^��s�p�gM����p�~��z��-�(H ��/�	u
�d�`�#��sg�)Gyq��[��	i��t-��z������̔�'s6���w�W<P�ۙgZ�F��:5����D{�=.
�k��EZ�v�eG*�q苍�w�z���P�&�e�;�G�:=wQ�^�]��b�a�6�)paU`
�������h��u��k�A�{b�B%�M�ڼڻ�ZS�H>�0={Ǯ���Ql13��m��F�yƸR���s���f����Ij82����+��Y�¼�܎����WnL����G(C#H���
���i���&���� ��sV	��K�l��l����Վx��㡌|�*Ώ�W����k�E��y��[�\
e��	��ϣ>������R.>�X>���zx�C�k�f����?nQg1�hsŉ��^n5kK�]_Fl��7��jh6�xZ��
,u��vU���}�d�:}u=�����2�᪌~�g&(],���ا�2\
��E��B��,��y4�l��ϗR����e���Zq���қQ�^E�XAI/�iS�+0_pjma&��k���+��I�S-y���p�6�O�x�"�[���C.���M����(��0���]ҷ�rI�M��~Uᲂ���6$9��gu�2z��Ǩ����&��un����8A;���~��=o���Rج��T�C���ˬ��F�y�L��CwD��\�2-4�r�C/�R�+��Bt��V�ig)j��\�\֛7��R3;��v� #][Qp�N�3�����3����=#�b�^Ҧ�N�'e���ܷ
�r9@�����BV
�3�7������*_S�wu��$����ܖ<E&<�/י�8[�4��k=U�O3�e����CW��7��U�嶵/xO��Ւ�T-	�~#�������s�"E|��3�yWyo<,b|��V�vm��d�h[�h[��l�(�P��>R��a���w�Y��Ϧ!���>��Fj�)���m`6�'�>8"�1q�3�Gg�TS���B��U ��O�ffw���-k�u�U��!���#Ak��'au1����mS�Ãӷ:��<��i����s������ئr�SE�1
��:o��$P0�$[��}��9Gf\�7ٳ's����ɯ*�����w�-��"��3^r	fV�-Nt���e�%aL�t�5�w���!��0�B�������J��p�����JZ���
,J5PםSl�^���ss6{	��n�"�����м���m�ZSPxOLX4:1h�W��͡��G�B���`��ow����ǖeKv��xU��/��L�Dæ�}^\X���c�vV�z�j��P8�K=��/V��(�H�Ȫ�{œ��)r����jb�"�K��N�X(h'ܤ&@GbtXn>,�u+�S#v������Hy�F��������K�ٙ}�.̪kv�לelC�6l@&���\��HĶ�_Z+�-�y��H����ہK��ֆ����.�p�:7GE���R��p��;��Ï���5�|�Ք������Ю��A��f����jy2��T@����T}���܇
���tgv�];�U�mu�9u9]L�.o]	V1(�G�O)R�omKt,����¦RG0U��k.�����xoT�W�K2&0���8���@�oôH�`�0���0up6,`&�0Ԃ��o*��ć�V�w����Ȫn�|���U7����������ā���Z��+����ɘ�J3;�����n�9����.��e���zр�N��U�Է��x''b�r��N�6by�Ѻ� ]d
�Ю��s��;�5;���wF��*M(���+uK��i+�iM��V��}f)�bV9;5��,���'�����ӛ�A�t�.;;����*�h�)_,�o��S+T	%ȭ�{���AOr|���d�m��wuv���uk�S,Wu=�J�p�d*Њnٗ&�ՕC�
���+bط4�%8b��cl+���Q�x��֓�����gWc�6����^�)�ө;�q�����=9] ��'d�G�I˲���>���v�3�\t z4�<8�=�z�� ޓ2�ҭq�����_�{���!���x{/�� :�QCR��B�DVɮ�`h��\C�WV�@�#������낗F�ὲ�3����i�t�Y����,�Fk�ɥxɽ֭'��o<�Q�Z����;�֘�� ��W n�j������ӘJA+)����[ˎ9���%�j�̱N�Ts˾�:!�f���.�y\7h̳�]کZ�2�hQv%.�PG�D-��v�@���p�,��Ư೰s2�Ğ�p��a����ɜEb�\N�l*�fa�3�S�l۾P,�kw/�:��\�1.���(7�[s5��X-��4!�=�@9�78-�qK��/��-���μ'mc��>�¬{8Lq�\�e�Y����e�2R��U�[�`R��z+��.D:�j9-g:��K�%����-����r����6���NV�͝���`&�ʬ)c7Z�շ�Z6�%�M�cV���TE<t�z�1�[�)iq��V�I�d���`ݹo�wN;Wj���tC�-a�֯Uf���i[f�N�֛+4�4�P1�b����%V���s�i��',�tGO3�2fe(�5r��c.�����1_
!@�@�-D�DZ�YEXօe��-*12��%c�1-�Y\k�iR�%\n1U�ԣ�sA�UU�31q�E1��-�DHۖ�*��̶�KGs	��.4q*�q1�����m��و."ʭjSe�F�[���F��`�Z�JT(*�Lʫ*+mI��b�jڲe[Z�7����-
�Kmm*es&�JܵL�0D�f-*�P���[j�̕5�Kk��#pfA�����*�l���(ʬU�R��-"%Z؍˂\��KIm�3
"&[�����+X��cq�[F�kP��F��-�E��֬X�V�QBۙ��Q-V�R�-Je���Ke�̭��,Y*fJ�m
()X噖�l�mm�Z��V*V�(T�m��0��Q-�em�
cQEĥh\���mEr����q,U�⊍m��ekP�`\�����T�����A�����b��r�S�!�T�R�*�AĬ\Kfa�[b�-��( ]�T/��'ujd,����9��.��	B-��'k��Vwq����Q�f�nͬv&l�zi�s�¦D��1�Jn�#�v�_�t(�o��������^;T�~�ʍ�i�%y�s�dv��jΕU�O02pٯ��6�w<^FJ�����q����u�C=uBRk���Shf�X����mm����Ѣ�˜�wmk�,AU�@]_�Y��>F�B͘'�e1و�weC(�6`0d\"��S����x�;��B�|,}�2��wH�����1�M�я�ކ��K�e�k#JF|ּ�Y��z�w5�q���������}���=��!&N�f3牉�td����x��i�9Ҟ*��[ ����O-�	�W�z�#�@���/�̧P���f�,�k<�{��@{\K��74}�(�=���m�c��6�]�����jQ����Z���X>P��{X��y�D�<u�1un�}J�N	���mUq����҂Y���Dj�I���>&�+l&������?{�em��_M�Rάj������Rr�)at̚��%���<J�s+og6	�ED��g�G41Y&0q*��`ׯ���9i�^����lb�q��eG�&̠b��L�z���,��M�O#�ӧkGA��N�������}~����=���o�U2ľhP�i�e���9�C��W݈:Θ��`��x�kVy�{ٓ���_��?����6�a�mfm+ީ�lC��)��>S�A���G��({�*�4*:(dcZҸ�K)V��9��3���Bԩ�ѣ>\�HpO��׬�1����^��^��Ŕ�1�G$��!>�ad)W_���>����9��F����C8cg�.��/o��i����R��(�aX2�� .k�OXN�oy��^ĸ��
�E�]&+8y��6���V<����3�WM�E1�@a�r��qxZ��>V��7�-����Q7��Ӣ����}}�m^o@cr�i��4X"\.b`����H���(��!�|��[�tC8�MM0��HJ��F�g���Y����cGO��:�7��E��0�E�(jv�1/�;2g{�9f��y
�3�e�a�ӆ��p��1ل���/���lŊ[7:ƍ�Wn��Y�&��s�Nh~6�DSTG�`*��m�֡�3�������Q���ޕ�I|�dq��q��y��}hS��|�,�"ة\f��;��u0���9��x.��/��z\;�ʧR^��9���K�V],�ZZ�^�-=8��m��|�e��`+�u��|
��� }P1�����vLv1^�iI�k�8��Ѹ��k]�rܽҶ0��HӁ�H�S�H�ֹ.6V'���!���I�(�+V���{{�}��z�(=ύ�P�NuC�͌�ᳫ�8�Zu�|OG�ļ[�g�[\���䷊{2C4%�B�U�V��X�������%���Ǯ�yU��P����]W5�ʰ��g���K���y�4t����TkaǹH��/<�脤!pu��Ӛ��+�ly�Lι�m�th5�9\q+
</����PWD�r����X��ԟ� td�mB�r�r���Κ�
�dP~�ԕ�#�K~o�z8X��0���:������7Y%>�P�2l��'Zf�z>	��B����iư�CDwT<�U���.M���S�;+�dWZ)��k(���C�"�v�at;��U5�"��WU�YE��s.��X2!e*f¾�Q���9�ŊNp�Y�J�0d*2�K\��l0�fJዔ�gn�����-`������2� U�"B�P��+�Ӛ���ҳرKMv��;Vo��ޢ�ʓ��fR�I�v��T�
5r��J�T�SE.��g^a|�	KX�SS+%-#o[ `����p%���	v�){������yA�}Wx�e�>80v�l��b��`���J���s٘�^w ���r4���n�����\Ѳ��A�(ّNmE��Yf�,(%��TD`�D9�[[%�M�C4��2��n�(�n���Oe�f����vA\�dY�͚<�K,�oq����+�:����a�i[����CT��[T�E����T7T�2�
UM.�Q᜷�+��u���Wږd {�x�9��E�q��6�������V�M���w�D��v�<���+˴�_�8eq�c�����	�w�n8��^ɕVt﹙��ެlb��n/����B�X��N�xn7����D�cϸ��'���õ6��=��-�� [��[嗱Lj�=�Sʬ��(��*!l
(څP߶BQ���sJ/t����e㲟um[�S[��!���5�Ǹ�����;�H����Ԭ���`]��u�;د�`��V�N6a��3Aqp�RYE��Ӯ?E�7�R�b�]�r~I.�.�����˷ֈG�^/��e x��,��P��ߕr�<d��W}�-����g�U�ΛO��6wmgd�/=BX�yra�0n�9eh����ۦ�ud�l���An*=Y���vY'�R�WFp���l`�Fs9����.^�$ĴV��g@Dӕ����:��u�9���uoj|"�������JA���3�z�S��W}qM��#����XeD:�.Iv0l�d�rͥ�r�&߄9QQҍ_Ҭl��̧C�(*�E6���bc{�=<W��e�&t~��������@����)�Q�T��_�2��h�	B&<
���ˆ��/���L�o�G�ԗ\��|Hҭb���|E�_/��:R*����н��ŭ{�v.}zt��H���ʡ��tV/	�ɪ�
K}o*1n��T���}�4�P\�F=��q���c&�ܞ���>I�8�������[N�Z=]x������4 ��q��ҽz�v֩�C��\gC+��P��zL�bĬ� ��!Uk;]����Y�9��qy��~Ξ:o)���4S::�8��Q��S�Q���5Y���0��y/����Ml����#�z�[��1;����V���r�*v�cX�֩�B}��跧(�$��n{��3�z衵����lth{��C��{�1,�(�s��c^��c�U��.��mΘ�a�\��>���:��\�N�����f�M��ڊ�(Q�'k���WY݃kj,����`iQ��#����wڶ���a<W>��l ��v_v���$��b�hS}�hq/�_����s9��1�e'����k����եM�fܩ���UuvMu���8:�n5r���,�%_tJԧv�~J��F�;�+���d#�����ȫBx����_����WXȂf��$<�d�=2�����ժ��N���I,�	F�Qʆ`�74����V��g�9<m�)z�l�~���_��y}�E����7�.Y���sҹC���Zޭ��r�����>����<]{�m;=nlr�r�H��*cS�qKR9{�u��K��5V=���㾏�q�n��Â��.ã˃���t���9).�WC�ʟ��S�t*�]�oL�V��u�ݙ�Z�x�Ɩ�K�Ǧ��>Z$�*�p�=2�����)���C�;H���ծg0q��G��5A_���le����8ll#D�z�^�%=�FN��v��nݎ;�UQ�}8I���������9�s�⣊�>�œ+��S�ͽ/������!
M\�Lk49ʰd��kC�^Hxa	h�^}�jgNTMsg\3���2�nX�x�Xܪ���c�๊�@�V�N.�T2x�_�Z��#پ!�(6r�ؼ�˳�YD������M�W�����`�e^U�n���S͝�_
�G��[.>z.�ZK�$�e�E�R�o.\��j����n�aC�-_�-�w����3Ԋ�9aǣךf����6C3��sC-'}edaZ'�צ\��Sͮ7�~�׊���c�7��e�a��[����ل��W���z�Sv7�5�Sk4ܪ���a�w���F�W^8����p�g�M�y�#�}�(`7��:V���r��չ�/o6c;��������������o�{T,�mY�F1R�+Y�F��<|v5�(����z����k��۝��ڮ)���i��\i�1ưE����/&,�m�g�Ǿ�N����)Z��۰�kұ[8�A(�U)E��K�X_wY繶�]f�͖���`L���̑ƥq��jh�W����Jo8bפ>���Ѥ�֝�|vs Y�ܻ���<�+�3���#����s|",h�u�8t9܀�^m�4�=�\wrmo�+���w�]C\k�%'+��V�#��������֝dշu.�*��{c�/Ѫ�˖i�,���$**4��4X
�{���fac�%�]�Ѻ���Ȁ���C��1�R:b�J��]a�ۮ���CD'Gn�p��$���B��5�|�+U{RL��
�"��g���Vta�1�c�}����C�龘E�jXu��t�����A��a�&��s��R�}���2,��	k�L�<wf��>���U��L�+��C��bՌ�e\j��gq�Y��x�{��uꇪY�{�P�C]H��uX�=+��:��< ����֓�/o���}{w�3�����U�zk�k�X�Zĵ��p�s��e���������OA7��fOts����U�oUԺ��R�LU�R7���2�R�B�$,�U��fo���lOb�=;��^M)�H�Xl��A<> ��,/���+m1�_��1�r��H�^�vN�p�O{���n�q[�8�LJy&��s���٨�:��C�.�1�%���c+��tw�]b�J�b�A����t�&��ÂW{YwU�`u��]�.��e��rS9Z�U�$�o�Ð[���ں���l�qaVP���x�i�+v+ M�5��5�j�Eus������N�F\h�B�7����lǹB�j�f5͝�n/b޺��Ҽ:`��V�Z����o���>�g81�zOR�����^���N8��o�:e�4=|z1A|VM�Z�kie9휰L�i�[�+�r�W@p'�����,�	a*\M��/oh�Y��X��:����˰r�ވ��V���tF�ok\j�W^tA�� ؊����<��嶐�׉TU�.�C���W٦ز1ə�I�]��s��+`�l��ü7�J�f�2���(ׅӥ���ڕp�W�ż�p��h>�a�:h��o�bLu���J�0�\^�ak�X��١�T�˕�l��[�u40i�c���]��*��>���x�W���i�#�ҡ;b���6���Õ����)1�s�~��j����s"��$x���С]m�vHqC�WG�t=�U~��u/׳��P�C���إׯ��2�(������mՙ�3NA�4A�{���=�8�������d[Xo�!��E��V��f������\�J�b��Ln$Go�(X���,l�tV�^ �{$z�T��.�XЧ��{1�������ැ��
�Q�޽b�l��y�\�p�2��[cJ��/�j�L�>7@�]|-�v��h^��]�Ԋ�N���`-��C9�z�T��u'��9-Gʊ��zv<��W��P�ucޛ7�۝OZ��g"e�ڀ�C�6�	ŏY(����0�8�{�Eu�>}IPu#"�d�R�w��sn,Q�z��4��N����C;~�i���Q�6O}x�a�����k�A/��d#�՝k5Q�Łv�����^:�̑EӅ�8��T<{�eu�|d�F]�
�su�0G�t�]��Me!k��q�f�4J���2�衙ҹN�+f(����4[T�w|�i��_�C{|��Ax�Y��� }֖�4wT�����xyvG1R�fK8w�LP���Ȳ����(l*�61:ގ���Gx��7���C8����x/�;^�w�xs��Kk����X;��e�Z�>Ӻ�bj.÷Z��BY�z�os�ؽS�>4�^[�oSu-4=�1���Ǐ'���$L��Afb�wI�W�g\�;�Sp��7jl[*�X�ha�Y���dW�	�jB0=r�����+�&^�r����K�[<]��⍩}}Q��L���ep�2�\�V��Y[�Y��
�`��U�m�8W����������l؎V�,�������F��PǕMէ�v�_ '�gQ��鲹-��dbg\�DeI�c<����ʅ���4�E��|�����fX�{C�-�Q����{����o��c}ٞ��;�8[���)L�n�;��LޅW��k]�(raz��zm,Q��#��e\�6n��c��������ܜ�}71_�>�V���]ރ>R���ţL�u�} +�s�˖0wT� ��gYBQ<��"%�<����N�*$=�B��	��b�
��b%��[��T�Ӯݽv��NhNއ!	�l���0)9V�*��0YO��3�m_W:ec����t�Q�+xX�3 7VjQ�AN�p;��
y�N%�cn*��.�r�~�����	�e��vI���.Za�p�/^EZ&Ȝ��mJ�P����w��۫v���:�.�[��#"�,3�����j}�b��-ջ���=V��¦;�vn�ь��G�uwR�EڗIםo�-L��k����P���ʆ6������v!5IӦ�޺fG�{8�w�yE.u�AՓ4��0��p�Jݾ��:������|B�Õ�k �)s�,Qu��R��R^���;��!X)��2E')H�vFT	�	 6V���v�4��o?�=�Y�j�`���ɳ�N��y�Z�gM�\�&J����د]�.�fm�,��Cq�f��5'WZ����Uۧӣ'T��V��"+sR0kݛR>�4�\{Z�k�ƕ�c�wv5v�E�PjC�0Χ���K-@:�~�M-˴&Ot���(����S֑ƣ��9���6F'uA��4��y.�{xY�m�퉚�Txc�t\q�ܠ�Rr\�AnU�Spf�cP]��Ǎ����sT�ȤU���Y�3��i �w������V=�.����)�ټ4�+�$&hܶ^��s#T4t̩Y�YZ0�.!�Z�:�(	��%v� ��^�YZ�]Shv� ����og*>��U(����j�j����k;��c{������Y�ט�իY6˗���D�:XYғM��Æ�W-ix�Fw����i��|#�[:q\x��A39��m"��j��5tt��T-ɘ巜���U֍�m}c��m�Lq`4�y�y^����X3y]\��uU�1����A�ڻ�p!�e��Rq�����G�3���9�F�	�G�gDӨ��3fq�.�ٻ�ñ��5f���B�o#��n�C�H�w�o�9f��R��&���,�-�����	Y�f�E�.Ȕj=Ы����Ю��ǜ�2Wd�c�d;g�N���ݫ�yt|�G��5�py8���_)w��>�(����OO�_n�A�.�cw-��;�<���ۼR`�B�ҫ��JM����XY�t!��0�&�÷w���gEpסk:k�^q㦣�X���xq��Qw�,�So:�Z��n
/lu�΂�H�����s�|px�Ą���x��e������!9!Y+i��]�BS���v��ևO�@�mӰ�rNW�nv��X�ήn�"��E\۲)d1v`��+�CĢ
�*�L�[��<J���S�w^��p�Qý��';<@���]k�����MQ����KZK�RXج���em(+V�Qƣ-�T��pj�-,[[i�0*V�Z�,�ֱ�p�\l�X�Lh"*��+�Q+DmD��Lh�+�VR��iqE�[U�Z�c3)%ʋj��Q�E���d�ZU�[in&&+pk\�pʴQ��\��f5��.1.L��-��ĦXZ-��m��m�+[j����qU�2�r��X�Qknpm�"���-QmT��p��E�PR�\�R�
5+Ls��r�*V�bS3m���ƙUb�mQ���L�KYl\d��fe)E�0V�ٌ�LAJ�-pL�\D�2�%� Ԗ5�6a�cEj��(T�"�ʭ�2֍�JƣjR��
���E���+���*�[Z	q�+bQ�l2̩���[�[b6��aAG)Ls-�崪Zcqj�����U��-�F"(�J��V���e~D��%�_Pe�������gi���ki9��v��6A����vqKUa�.W:|��9F�����@��o��!��)K`��vї$����?QZ"R�"С���i���U�s���^�!%�{L)�oe��u���%�r�N�5MÆ0 ������#5W�c�S�Q�Z@9����~D��o��c�r���b�xZ-L抱�@x�9V⬵�9�wYU���e�화]4�	qx(� �鷮�yT!�"��X@���*�]��Q(��e�^�6�eI�ۻ�.�0[7Xy�W�W�7)�~n�cc���Չ�$���f�Y�Ԏ�\/���z���St4_ٳ��MN7��M���� �����k�˅|g�PTdc���$$G��ğ:�{z�(s�z9a
�F��k�/-����J�l���U��lFPY��-��!�"G-�w�y��݊�7\go���h�[�.��]�Y�C7�m�\�e�]ݖ�N���Q�Ћ�(�դYΒ{���T.��VcZjvZ(���#���yi)D<�#MFV*Q�R�<�f*eD�A7H�Өq����aM�U�.͹jb��X��(��q龏+����U��x�r�l�:�:7�@��ʔ��n�Ӿ�qN����o��n��*7��,�-ɇ�޾}�1����M8�D�K�+sW���D�f��{�Lluk>�:��dZ�/gd���0��YZ���Y����>�w�V��p�Z.��G��a��8 B?��|y-��fs��y�˱��Ճ�
Q�(���3�&Y�V���X�Қ�}(������6���������6����˸~P@D�tƅ�HT4��.�؂�ܣL��L��P������`P���r�l&��ɯr�qWn��e�D���]5j#!Λ���uB��G���5ow�m������,���ǃ̝��]<�_�l�4�>z�v���z���=��,�eΑWN6�ù���cH����z+,m8^���g�Ê��~�,���nu�y{l�nu�=��]E��A�c���`>w�,�^z�F��:��::V/��|%b

���l���E�2�	����LE�"<��
�͋�O5�b����˥�����kJ&}ֈ\l��'�����>.*�L�6�џ]0}}z6�t^1���'��j������Tߺ2S-y���P��v����~	��4���-���:ɔ�FB��?w;���p�z1vJ������'�s*��<C�U��m��z{�¼�ڙԂ���&f���G/jm�J��e�7�2d�gh\���mv�F`ߍ��!}Wn�_r�Ψ�[�h��v�Q�
:�x�QwL��~��\�]5ߌ�hF��i[��z��;���v�+�nFQ��У�M	�z��kR̾P���H6����e��VBuo�"��+v+�3���"L�~)�=�Ե\,͍���b��U�C�����w��EyR,�\�Ok��ίl���5��,c�����ɾɗ�x���^+|��窑�V��]:$qH�.���GS�w+�o��s���o�6�F���ʡ�%[�-՝&Q�lB:-ʈV�����|�θ����>����T��9���u�~K�a�����`6;5�U�E�D�z�t.���{[��9a�4��kj���K;�:aߏO����8yNَ�Bȑ	t�c��7��ð`�"o��R�<x[�eg�׶����L��y�4�͖f��
2��!e����I�$�_��vm�m,x�֎S{*!8
߼�K#{�o*x��u`���Z�Ӹ��{7�(P��%@?J߾B�_(��N1�1��w�JJ��۪�e������nr��ԃ�lHrP�:n�u<8��X�&��+_�vS�j��;�<	�>�޺�ysF���Z�u�c�꼂N�fR�&orΜv�^�v�S�Zg��ݥ>�}WZ"������GH�@�Gm��>Քz+�δޅv��i8,��[z�wK6ʯU����K-p��p�9�)��t��C�X����A��"Į+��J��>�gمߜ����X��0	J9&,+�1@*5Lړ7���%Z�|S���<��g�l��f��|.R)���2�8I����{���������jr��Go��X�f�Eyi�t]�v�l'��=]ʜ�(��Wi�5.��(���K�lx���z��jN��)�-U��C1�_o�M<��_r���U�ɑ�h˪`���X�eO�u;�+\�C6l�^�$��6s6�8}��Dv&k���jY�1l_����z����g�4�8����6�Vy�81:ކ��
��v��74��>�Ј}kD~��0��Kk�U����<��o��:�)eu�Lv4��߇7��z�T3>ړqQ経箊Y�-S4�<;��1)%+�^��q�[��࢘����g,s�� g�cR{OJ�T���Д��u:��նo}��-���1�ܺ ����+��*���(▭T`i�5b��3�i��WA}hI3����E�-[M���;VjI�x3����e�R�t��N���S��Vm#|WL�)�;�s�8Mô����3p�R�v�]�p�e:&�_J�^���@���T��-�b��Vn�̮xd�.aV�Q,�Σճs��ӇQ.^w#���,IP���+�v��8���}p}!�޸LX\㕅�ݥ�woh+�~�~�gz�M͕V��	5�P�T�����n,k��`k ����eE���S0�i�/x<��o��E�_�K���bU����x_���#�rQ���\c:�n���8"{v'2.���FV�u�1�B���=R��Vx|G=Zg
� <��ɪ
�k�3��� �����WE1�v����E��� �E?��:�`ZO�;氯a�wÓ��Vg�m��\�3�^\QX���'F��$�D�����J�����x`�W��3�3e����.�YA�v�R�JE=c��C���qxZ�!�NT�W�-�E"x^�W��K0�i�������ע2�8J\0k'���"w����XE>��O�G}��.^��}���3v.�YB������62�[82%���!����4&�e�G��8�����g%�ΏN�:�dB=jkO��V�"�k��+ q�_��/_ִV���8e�/c���ݴY}��2�sU$� ��G���%��qyU��r���=�A��(�����!�o�Ӿ�6�s5�=��e���+]¸�G��ՠƇ�Ը�%�V�@>˽�j�aw�SN�7�3�ߙά�Dε.��ѐ#Nu�����n�X�]OzW�i۩��Z������*�T��[]C;Z��pa|I��V�:i��S���Њ����;y*Z�bnV꫒����>�(7��s��Ҏ�f���b�*n����p<lj����H�S�Y��V���W4p�7Qp�j&�K��+-76�77��ZZC��1��;
__W%��hzQfD��G:dwE��#D�ֈ�Hud�;��V�V����_�L��[�:"�2G�Ƈ_�ڜ(�s�|d:��Y�\�+�wQΧwr��;P'X�sT;"���\]+O�l�r|p����G�º��jo����Z��qi��<^�y����-#�`Z��� �&i��9��ULߧ��KC��[����,�.rw!�Li��[�>ax0�0�:L��s���O��Rˊ��Ok���G����8z��c3��Un/�I4v�Ӛ2+��,�	��X�Hi�&<
ؚk��tx���o��+�qʇZ�Pũȸ莫�谱�x(ꐻ�?�De��嗵c0��Dݥ{�P�k��*��Rڔ��PS�6<p�f�^�Ԅ�=8�E���'q�V�;6�M5�r{�!�	�S��p��H�1�
@��ݐ�5�l�� v+���0�;�Qt�w�uM��QS`��W.h��g�y&��(�`�[zNF�Z3��E��C"�j
�;�u]ފ�/�ʹ�&�D�G���o�j

��Y�|m��ƾ�9�/jQ0�0������Z��q���9<§%i��E��҆���_�?�k�%��EJ;bKu9Χw��������ܒ�7D�$EN�i�]�?��u�j�B��Y��HP�� C�R�g�q�6y�;����@��ŋS�֪woha�m=hj�۰����޷
!	�َ��D˪|�/[�lqW4X"�t�sa�d[�ya���|��tx]�.�EF5~��s���s!V��յ/h�c���˕uq����"�^X��y��yר��P��c{���/�ׅ�T�){���Þ��x�[��p2�x�K���b�ݻ>�g�=���lL��FZc1���%x࿛�f����qyF�����tVV�6$�Rm.�zz�o��'7]r���Ta�Au�ϮtTG�Y��<��#uӒ��Ŗg��ՈL�>��1�l�I���wƁx���>7���ݨ�6[�71��:�O�1g��"@��}4o�C��3�|�ע�-��tњ�1�c�z��/��r�+�Ǌ��G�rG�Y/�1�>��GxN��8���ɂunN��J|���K9�w��8[ml�y�g���a�u����r�/���-`�����.1�i�Xw�=`��uʗ���]`�q7�8������+*�R��n�hB�v�c��f[��Lu�缼�S����z6<抒�����lJʠa���Cmܽ2:[4�a��sQP5z�N�{��yl
�P�¿s:]��*�k:E���9�{��c��A���v�K2pu�Z/�<�*�O��(tg�,-6�}��W��Fŗ�U�n���J�1q�d�a`)ᦍ��sp�!�uXybβ�����۷Q�䛷^�S�ǩ�ڎO�ղ�c�O�fU���:����t�rɽ:�.�k6-��壩���F{F���$�c�9��{��x�j����ƣ��������L�[���x�z9��ey�<*,w��@_u]�oۅ��L~}]���v_�D���ƺ4Q��n�6 k}9m����`ܡZm�힨��w	�l�o+#�N�N��j��M�`�!�G�\�lMwiRN�x�1s�a=w�|���WٹH9���SU�9���N���;C7�j�{��R���o�mͦ�v�\]�793�M��B*ӽ�N��s���A+jYò���^o��;�z�f�,����C�ɱ=3Hl�c��U4���ދ��ƴ��ar�
�X�W�vo]^����M����W�1"b�bzu�aN��%A<��[F ��߹)���X_m-��������GVj�r�':�k��j�e���t�B��J{�a�oM�b�1B�T;+����=�gX�vR]�{ZS o�R�ݶ'âz�zyo��݀�� ��f��d+��;ifN�Gm�ԭ�]oV_�aV'�a��@򭖣�8Bw�b2��K��ޣQ�Ů�]�OuV��:�I���9����P�~�k�̪܌f��Z{qE�4�J��ԒSc��)�s^b�gK���qׇ�p�^T��|�-<��Xw���ܲ��$�x\���2��	�W����Iا��{芺�9��N�/N�P{��� L�'Ƿ����>wS8�Ԏ�(l��I|q˺���C�V�X3yv�t���RG)��ӽ�;B�w�o$+"��LҶ�&�::�@�2=�3-������FTջ:׸{���aI���h>������o\Ϭ(��M��磊8��ȇ:�����瘽#�H�U�m��%�O�mV\��������)<9R�:�IxF��K�/�7V)y	�Z~ B���/U�m��Ҟ�S�is8�o%�(�I�ߪ���T�V)q>��sHj}����t3e{6�T�����M�e�)_��b��o/&g6t��	��Q�L�ř��#�(s���Mw)#K�:&J�Nz͸��1+�{{��r1���nk�t2z�*����3�ȮC�23Z4)�Ǘ��J޽ٗ{qƲ�.��d�{eK�]��ݸά#ni�L�bFE�n�t�v���zﮡ'����/����s����J�9W��Ƽyt�G�ׁ|���ۇh�;��+O^gc��Ұ�D����oP��N�ׄ*޹�_��x{� I?섐�$�p���$�rB���$��$��BH@�2B���$��!$ I?����$��	!I�d$�	'IJBH@�j�$��BH@�i	!I�$$�	'���$��BH@�$�	&�$�	'�����)���b���o�9,����������0�_�w�$QDJ �� H�UPHTE J�  �Q@T P( PRRݜP��D�%(�(�$
AT�%
�U*T�AT��	TUA�TIG�� ��(R�REQRJ*!
�R�R��� �*H�EITDQP�D�E��%(G�W  ��ږ�LLڬ�hf��T��2�FZ��B+%EVB��0�ڶ�S#��SeUY���UF�UT�  3u m�cf�*�@mR�6�Z�VT[-�ZmZ�ڪ�ѩ���V����,DՇ
(c���%"Q� '`��E
(��Q@(P�E��B�(�(s�:@(�P�;�P 72��Pj��R��KR�b��F��dڵ���[P��IERRC� wU*��3f���L�H�V6��Y��j�ڶڵ��Ue�j�ѶE���X�lXf�aVT�(��)��� ���V+���j��EZ������hL+J�kh٦�M����d+3* *A-i4�*�T�
��� tRJ����!-��e5��b�C3HFŘYZ*�,��(T��UT�AV�*�Q�  ЀN�Z�Ձ@��*L*�Y1B�S��L��� ��"�HB
��U�  -�m���0(R����Q"��
e�@Z��j��"�1Z5m����J�)J�*@*�   w'T5V��ʒUddEV3U@�)K&R�L�I�$TeT�kj��$JH� g	@0
mE��h�Uk40�F�%C,AU+EU��ia���hl&��HP 
  j`1R�T b  @ ����@      i��&�&	��0`��E?�Q  �     D�h�5<��i�I��FM� �E$1T�y!�mM� L ëln�ǯ�N����c)�_*R������BԜ��d�F&�3%������=�(��:((���Uj�(DPR����,�(��P��S�~A���:�E���2�@ $!	P� �� �!�@�@�Ud�XQ/��}���Xc��χ".oԄ HZ�b�e���
D����ֲN��U$�#-ߵ�]����q����DZ�0�>;f�K��z���ݾb���Ѹ���m��v6ء�/X��­�skt5�%y�^����[��h�˥lkt�l!���"���D���o^��"��^� ��;�Q�+
�Y�m!��f:��� kܼ��v�ь�*�Ԋ��oCh�+�kK���Ra�@�;t�{�(��fA�b+F�f�{z7�`�m��e�wA���mY�'i��vq���[I�դ�
��
����㵻�E��ZN��o���lȳm51�f��·0��
���(��1Pa��l�X���l]���eZ�r��^�f��@j
�I
x�~�U���xl=�GQ��Y7#v2�z4�JU���iw�,���,,2�4&M���|Eb���ڽ�F�b����S�uuU�j��[zs���7YIk8��f��`e�t�ofr��f�M�2H�$��)��ڈ��-�c
�Y̴H����PG�¶�֛����d�D���K�vm��A�}�᧫��T�^�k����
�u[�v�m�kq{�;J���[R=�z�b�4肮���n�V̗C$.hJl�i�gSڕ*��aD����f='���6��+)��ww׵��My�����E�h�ٶ�}��A�a�c�ι �Z9V�,kr��Ԅ]H��U�F��[Բ��/+v� ���d��T۪B1��#^��;��Ve�n���]�2}c)�1x�Ϧȩ����M9X���D��Y�1�)/��ӗ�����O�(���0�oc�����sv&��P���f�̈́��&���:���!�|��I�W�f��@
��l�]��ׯIӥ�;O6�Q���خ4���\n9EOhl���gm�e��$;/X�u�tL�Y֮�e;U.�ŀ�ɯ�{�\(�s�*�a���c����V]jZ�R��x�Uq]�`X�����`Ha%o�*<&���N�h�h���ܻ�.���K�6)�JE��)'q\�WZ/��Y�|���CS�X09���>Sn��7��C�:e�3]�ڼ���Y�u�l�l��<��@G�S����;6Y�����hl�͵�޴WV�h�YJ��$U�`�B\�����:DL�Fj.�s�	���G6��˓k&��y�ĄK-n���-&0u02f^�{:C%R��C���;������
X���^�e��c8bF���x�Y�7"�X��z����ƅ��4n�+)-��i�7j�ᆲ��\Xະ�	u��5i�����j�@��n<tH8�D{�����eñcd,�����^�c *a�R%�`��SGR�"S�gz�+7in�'}���iY'��,�i���Y��n����S)����#d��:������+��cX�k�+4��nm�y�cD�n �V�Ķ�㭕v��^�	Tޕw-dS��l�<�7iP+�VV�!� Z�����ф��X�׺�ە��ZV�����Jk�]��hB���k.�Yb��mc߷Rͽ��(���8��gnS�VΊL�����D`��^Qe &���g�~�D�	H*��,\nw����=&�\�wOj|aҕ^��k{/6�m]7t�æ��W@7�s60wNl�WC+[��ur��P��5g(9�dǴö�s��ŭ��L>E���[[�P::�/����k@��;W��U����=�л�i�x�۰�f�J�� ����!�>�� ���
�skp����%�r�չp�:%�:;�ݵ��
ʺtw&��*�Ab�_�]b�Fh3p�Z�M���ڋ5f���K�t�͓4�2����Yf�F�:��2�����ce�y3,03��]B�$Z�*�8�Q����]�b�ڗ*լKŖ�UF�ts�6��Z��)W�ַ��)+�r�w`į����ͭ.����x�v��V�ې����uj�aA���+�O�ޮG����y�%�,���݌��m:�xr�cA��V��Aۚ�`��Z�/��u��X��&��ٯt��8-����w�)dx6�i�6&�ރXoV����ɆK�Q`Ď�i�v�܃F-"Le�鋔���d��R��q���7���Z���TIaI&��NYw�]���aǁX��g&Q@K���(m���ϷM�
�fʑ����A����7�۬GW-�Ei���YK���tU���Pf)���G�E��4�//7ie�-|�A���=VVn (�gwD�j$�oVcG,˥�@X2�پ��ڏ�p�ʸ�N��kr���7
ś(�ʻD]9��c�v-�]#��֊��r��h�m�N��k{��,�6B�)m�KP(�E��eU���-DYb��+F+��`�r�8����v�Tm�OZb;����HXb����9�a��#l3�yHZ�i���"l��PU�L,�
�f3[������hF-7Se���nQ]-�X潔����fAt6�r&r�V�1]��Mo �68�vV\خv����AQW�SѤ�f��U�V��A�����$���Ɗ���f����V��¦{���M04$��+$�)b)�C0օ�w���1ѿ��vJ�WM�M��P��ւ�+w��89-
g�(��w�n��٣n^ٺ�vVi�Zel�����ST�'�<�f�p椳.���s����D/�n�A+S�d�Uۊ�pUEtB��rD�V����r����p���k,<Ңg�El�y����,�D�w�wFM���v ���b��m}sS�!�V-˺�A���A7ib�ܺ�2���P^��(�O]�d�fL�ct��+b�*�X�eXL
b�4��[��<xk�����-�x,���ERާZ��oiku�')kģ�tk	�@#�:�x�`w�!/ b��[kf�Wj�hC0�h��+
j��(&,�5�d�7rK�F�nQ�a��BG����0�zqS���.jhؚ0�l��i��w��p�a�4�D,x.��
X�Jۨ�f�☓�z$�wDD�κ�A�JX��4���vX{�R��*�1��D��Fvq�f`?e*IΗ{��G2e�b��q�r܇70��2DH!X���2Pe�#�J��Ѷ�M�R�U��Qә%F���iZ.G0]�������556N;ndY:2�G��hv��4F�d�5c�YA����u2�(�!��X� ��_Wf{8��W�����YK*�oE7�m��V�*���+r�a�t�+jd�����@�:ݻ�Ya-'v� y��SĠ��!J�qYN�ikNmXF�qU���V`�R>�r�ZI&6�j�}y]i�w���/,�X��Sb�w��I��Vb��K���,��R�D��s3.��Ku�S�m�w4Ѕ%��TaM�X� 2�@^Ǭ��z�xk��n��9^��j�uԣ�ຉ�s)����݂�#j��Y�&�Mx����bC�ES-Zh�x��M��v	EU��8���1x��n��n�@�p��ˢ�Ú�N�����[�aN+�t��D:2�M<�&�����_ �DЖ�`�ԥ5��d�����)K[��Y��M�6j�\�eꬬ̡R<�gEl�e�5fޣ{��J�#��4'��:CF(@ޜ$�'l�U]�����Z�HϞ؅��ZzDZ&�ݦՄv��Y� ^�ذL�*�-COdh�0N%�5:�����&,aU�@�ӌ���
�K�Ɲ�Ǜ����f�V�G��j�PT����DE��*��Y�ؽ��-K�#l�,�7�KL���e�1جEHL�ǔ���Pi� �Glm�:�*C���I��(@f�H �*m��N�إe��pv���qGq��MK�O��QX$���7g4�Ƭ:��kPZ{���!�v�U�l���\N��VFRU�P���l��Z&����I�F�"��[��y��Vƚ(�md��s
���e�8�	j�[v[1[�܄/��)M��KX�x��D'^^<olLZH[��[WD�����6X��+����f��6<��ѳb�`�^�Y��G��j�eյR��GkoZdm*����e�p;ˉY$�p��Xkv튔�1K���j��Sd�m�+�dݬb�/FVA6b�p;��6�{Cc֠v]+KٷM�Ŷ2���)8m�$��M���n�-jAkJ�@8��Xxݮu��e;�]�l���Q����(�m�V×K�)����\(Ժ��*W{���vy.���:�6�۶�.¹|�����@J3EfX@�'AF�1�)K�F
8cn�	���h�r���,�E%�k��:+h�:��gi�s�����x�fY����$D^�O��C3~dT���Ս��Yi��&��lܹv���茌�d�\�A�L��zu�vҰ�GGp�B�wM"w)T!��&Q����@Y �̧a��e܋���MlI�!b�k!h��0t�GQ���GV2(��Gh.��ܬ�{�r4�RZ �p,�cV�ق��uYQ�0<KR�d�'@�Q�u��"$6I`����Ӷ��`)=قɠ�^b�#���c�4��w޳�o�2�hu��lgC�oU���ͺո��ڱ���,��l����0q@Zȴha��Y�i5l:ةCysf��k2h
+:.����kzNҠ�����s���h��$�=єޱ���oq�:���4A!��˥@ZN�52��7D�|rLܙ����r��Ii��:���ۜ��cs���o/E��y���ge������xW��J�q��V�W,y[�݋��A7�a�	�t6����ۗ3C���fƉ�e��@dW5p�M�4���&����.�1���XU�Õune/e_ׯ@T�XE�:�� 7ĥĽ���mf�p"GлX��h�ɔ^�j�핸~�el�-��܍r�XlK6k41���S�ki��)�I��H�jԄ ���㥡Z/��8{�c��S���9���~�?��:�WݼΛat]'.����D�>�����zE��Ww,e39N7�Ef�U���p�C7�B�n�Wơ� �sZa�,r�aal7o�����т�3nWd���g�5�4�]���"�SU%��ohe%���)˸��w�����i�'[��:r5:\���)����
`�	����͙Ɠ�WBn��S�ҕ�D�o�Jy�P/0񼽫�9��Bu#��R��E��(�-K����;��Y1IS_X��Tܭ�dx�hW�jyҬ��Bb�4vC��,Ol��og�J��3���x�h�ӕ$��x�;���ۼ�U��4E�|�������>k�vA�4,�R��.��F�����<s��^�1��v9o�)�%d����K\d��y�Y�:�U�ҙf�X}�>�Pܤ�X�A19�˗E�R�����1û�>ZQ�U�e�$��U;��s�[s&�t��3)C�E�Rӄ�0$U��h���� ��8kCd��qA.�ž��a�[���(<����91����:SQʵ��H-���Ύw��.��@YX��Fq��k`�]0��j�%���ܠo0�a
��k��79o5z_t��VoE�9!�&���]e��I�I�ΐ�k� ���0��׍M��(r.���L��	m���p�U����^@�	*7G����$�%r�E�+��OQS\S������oxR��܀�����7�p*�_6^Q�'{�ͳzc4�,��Luda���"o+����^n1�Mj�#tY���/��x)�䡙�i�7y�keꗕ3L�$>���;[n�-ؖ�v�t�r �1*���^���;�nl�<Iӻ�"�#7�m9׹3���&T,����s�{yr�=Bo���)���X�w��W(�T��rX�19jt+�:"�Vw�t�VIҸ�;��#��!\�o�PN�_-7�j��z[����ط�`u.���ս�B�g[����-r�d�c�(�iWnSw8�,����g
�Aԃ�8�N�	�k)d��뵹��H��m�ꔸn��wc��;sC�F��b�/7��L�矕fC��C9�Yܭq�@��󺦍�=IJt�iw�~��ɧ�#+H��=�.���sXUۢ x�*T"�5��HfBgM�PvS�ɛTWIS�ĸ��2n�U:D_�D�{^񼠹&p�hb�g;M���Ln�O6.�VV�'�(����өX2�����PH��mSՐ�!��T-�O��.9J�J<1)rt5����ɶ\jt\�,�Meʇ]�3ز�y��;ptrw+uK{5��Sǹ|��3�f��Z�����5�C����_�0_p���25V��V�Z�E����+)�`���]�6��3OM<o�������,���;�����)λ�a������xxT�)e3v�˒Ѓi�޽w�eQ�[G(��)N�}�q�%�/&��5G]�S�s8��m."c�7t���ҧ&u|E�˩y}���N��ܺHMW�9"N��{��7'#A�������j�GF����u_f=���+�г�#��<AJ��������&D5V��,���s� ���M`��htA:�^i���=O�=�-����(��T &щ$�G����*���GI+!�<"`$�Cx�as��;�Y�4�{M�)e&��:�NXw@_E���S��������S]�\m�d��vjם+�q��ķx%Yƴ.ң7y���xְ��mu]v�ɣ)���}P���V	�hh5m��aӦ.���]�(�C1��Za��چS�ͪ�ə�-0X�w*�l�`0�$���樣�A!�]nS�-]�j���4�D����m�+|�<��W��h�jf��'�.�#�6Ҡ�}��ʌ���>���x
�r�@�$4ܩ�%+8bw������576t��ٺӷ�:ܢi���ݏw����ض�e������]>^7r�M�3#�^m��	�-#��`E,�1��q�@Y.e��o[3��NҫN�h{nn�F6�\S��m%�c�oy��:2b���M�t@ښl�-)}xY'���*��d��Skg`��՘�E�NRn�9Wcw+I��5�/�0S2�����t�S4���7j"kTy\�V��ʺ��]8ͫn��2wC����!ҷ�7�(���1��7�0�U�G����Y��[.)I�W���+R�E-���}�vx��kJ$c���ǐ����Y�_b<�J���j�F�S�s[��)�}u}uЌ�u���!�pr�H$��Z/�K����*_oe:��m<�׺&`�l���o�F��L���Yl��Ęf+�T���ҭ�Z8�Y�,�N�S.$�g�^��p�K��Ww���4�����6� Z��qu1Ӕ�{���@|������w$N-�H��K��P��/.���F+����=�u�di����B"�Gg��)��Z�N<2JW`���������p!��ɼ�lkh��'1��u��:�m\l]0�dT�%��5���e���	�c��^M��#��d�j���xW������B����4�d��	�M�9T��5[��Q���+V�ѣ����y�-F�h��j�!�ɭ��!R4�N�,�"�n��[	����BLW�_V;�T6�֭�#gc���M�x��&"�����·3�÷�,�og�!m/Bc����kiBR̳D��gU_Ӯ�ݖ�	79A[�q_���Çϒ6�P�6#:"h����yN�5�fq�����s4X�S�%��6�b�8K�r���]Iv���n�G��)P\1����6pK��9���L�ĕ�0N2M'gN\��?�7Q��po1�r�f�E�BB�b�ȇ�K�j�Vi�GS̎�MH��M\��|�|�'oky��w"d���"���E<}��1c�.s�tD�n- ��V(1�4�[b��#qI�ґ���V�ݱ$�,vwR59��a�[�9�*����e��`Iw�r���M���VA�6䦙];ye�*��5�t���މ]�n�*Z�G���f��D���xw}RɥTQ���4�� �m�j8�5���F���8�ѽ��V�v�V �C-��JZ�P��+tv	<OՎ�E�T&n��J�Pl��u;<�MK��]�"�m�A�xE�YZq��{��7(�6<4I��{n�Ak+����"�*v�*��1�j�n���ʤ�s7sl��L����:\����(v)����"Ś�+��V�/N��ku^�:I�oVL�5P���]��x�j�]�u�m6Ї6�@=hݴ�6��S��������ù���d��	,�}QΛ.n����S)��A��&LkL�Gh-9����fV�� H�V�XT26�^Q�r{���ኋP�w�.��[E;"�\��{wʚv��^j\i_cd%kyl��q����E���AW���l��[��oVk�~�H�LIt�V�^ݶ��n�f�/oHZ��8����M�:;+l<���e�3'�����Ԥ��c��I�.؍�<6k3	�[X�Ֆ�K}ҷ�۪�@�q��]]��nl�e�]�su#Ѓ�t��f��.�a�8��Qq�q,�V:�F��ez�;�5�+������*��n����&�:-���v�|Ge�%�`Oޭ
�3O��D�7�\Gw����/Y�Y��3��B7ܕ�:I]���ԛ��cF�E��.�Ǒ��n޷�fC����ꙇvM
�Cƶw�N�o-Vp��mg;�A]ZL�1����έ��JcL�:��2(��x�\1����)�n�}A]2�U������f�P�r����r�}��@�)Qc�����Oe\K�Yz��^H0<{c �J�iJ�T�Aݗ��8���'5�'�6��ݴ�I��]�Md'$�����/)�=��T5�%�`Jk]�Ss;y�gI��b�b���*�N����M*��z�{+���u�9)�}}�1��'(ok7�QS)�b8�o;+_b\r񁉟�����k~T2f3��i�;/�*�_H��˯5L�u���5-�g�_?���R��H��i���� �>�|\�Ê�8�v�)��PF�u83��KXJ�85*��oa���0*^�����>u�gI)�e�Z}0��9K���E�V�e�I�1+j���Y�u-]gR�H�О���7]
�������u�sJq<���s�y58�CƲ���\�S:�mۗP����z�Hv����׻�x$�w
�|Q�P�IZ�$39[O�/c;�X:~��Q��o��.M\��W�[!�
;%��YOn���L���f:�J�۹�*���|�mA�{.�}���{��$S�j�,�F��ܣ%����p���m��Ib͊�=R���9�p�Kdَ������^�,�L�R��l�*�3�T�VV%�U솅nṱE�l������AN�,t�[�Dk+�����Ʀ¶ժ�H���c�'����5�����S��>��%1�(27��-IժQ�B8��:�)} �T!�u2�-ǴF��O%z���f#�TQ۽

�������T�2%9ۯ��C��7Vj�[�M�
+J�k5J�C4��[������*�zh(N��n��po:�.�y����$�r<�8�)�Ԋ��u��Pz/�6�7|�K�<��/�:����t�#�9��n\ˣ�X�c�	=9�rB�{@M&��`|�S����Q̚ӑ�%Խ�R�ymqҍ��K�r]p�V��)�m�Пй`��y�ԙ�9�Qu쒺���׷���6���8�$�I��%J`�a�'(�k��\jm��tmu��o.l��M�:#��L�>��k��	�r��t9=]�]��k,CQU�׬���8�m@���We��|H��ܤ.�J�Z�r.�wm���kb�\�|.e�etf��Yw�%7!�wj�'��5}w������h��+�>����{_n���A�#��JϋU{���֢� #��.t���)��n��:�ĕ�I�Hx�Yrj����f�|�Y������9��M�����)\�ޯ�L�}�"�s$y	�6�**"
r>�����4N�/h��Y�8�k�n�ݣL�r][|�껜�U]��'G���nĳ��s�����S��3��]�4��H\��0T�%+8)]񊥌��FLk����ۼg���pt`�5��mk�P��km�5�����B��=��H��brX� k�M���;�Eh���Յ�)-�K�Õ��o �c{��Y��oJ�DR��� �CE��K��R�˝��Y�^��p�
H�uu��h���n*�;����H� tC嚲��!}�_F��sn�oA����w k-�Nm���>X�$`��;���CZν�w��"
I�z�s�z����u��%�LRc�m�]��ڬ���i�d��n�m���}��w'{>]�&�:6�Ηccn��)pT�����@l�߭�+9V�0c���#�N���c�1�	����T���6B'VM]�y�9S�cc�:ӫO�ÁҤ(����vW���<=W�t�Nƶ�՛��n�5=D����mP���Ldc
\�|IDr�y����0ꮹ��"�{ĪaR��Y��b��K
�>�ܫ�%�;Sr�u
����0��pI�Ht)���}��
 F����v�{�Fd�!F�	�� �i:^�Z#0�EY5����{e��P�za�g�Ѻ��r�����U�bv�^hC�p�|y+�t'*ء|��yN�6��m�P3l@MX�e;��=|ݙC-���em���du�n���-�(��
?1�����g,��� �I�9a�@�����ݙH�1)D�)���y��m�r��q*��JٔI��]& <ͱ�]���f
4�^K�������3{r��R3���v��Z�R��I��r[=�ʐ���)і���
=��^��*�^�'�� -,U�ŁǕ����E��h���<`�5�)�/2δ��BG��$0��wj����C6����:�wZ�<&�sf#X�op':��̔��Ec�2"���Y}/�0gqP�e��v��-�c�.L�=����٘x�ͤ�F�����7L��VY�
2��W؎�����`H=кXg��j{y|й& ��2*T=G�i�Էx(�U��n)wYrl*�)��|�]1qc�v�������i��*��R�N��7jD�4�/���7��է0R63Aq�6ns�U���Q|ҧ�r�PY��yV�\����
���C��T�Ԉv@�-�k��鈪�'p���:;;:Jh�-ue:I� �vۼb�]�tF�.��.���Pie�RQ�����w�innʄ�b�� �ʳ�c4_�@�^*HU�:�T��i�S��حJ�W`����3f��ġ�v�QE�ل�CWLZ@.�vظM�B��Äg/�E���D�R�Ui)1��-��l3���\/�zK�[�V;X�s��3���l�dXa�gt��J"�r�1��v�U'3��--d^<Ö��E8a�؄^pō<�5��6�lU�M�3C�+t�7lܨ#]�H��+N�wX�1w5�����#��B��S��SN>��9}'9�����ٮ|3;E�iV��cC��aT{t�Y��oos���z�Ք�	������jn'K6Bq;��lWh�'fT��R�,�3'72����]�l둘xg�K�0^]0��49B��f����۠iMce�h��x	�A˩�ݐ��l���N�a����݂�a@l�ُI�����C�o��:���d1�X��ac��+��6%%ګC�/����EI]M�̬�˵U�q:�t����wi,��n��g���(j3�R��<��Xϑ�wK�X��ݿ'�t�>�C8�s\���݄Q;yXd��]]
��dH�Mà
4�ŊZ�v*I�N�7qd1��D|�=Ɲ`�ӓ3�;�~�6�6]���;�K�=sq�å[�[�n�1C��2���-E[�ۈq��2��	a�R���r�c���=��@�k��f�;�B�e؈*L
��Nv�e�Scu��C�����rq�O��{/���	Z���MiZ�`K�>S�&��*��d��]���M��|YJ��͹�e�;��=W��v�g���#E�Nr��Nfku-3��M�nta̹4��c1;��s���d5g1�anH&�J��=�,`�od�R�{q莗1iE��\8۸�;h�v,�V�Jm�M�}�gVdڈ,٪�=��ʻ���[eh� ���L�g�c�f^�5=x\�1�
�jj�a(�����Z0w���˷�y��Żs�Z��jtX�_.�%�+9�}�qnT��1P��9��q�Tm:d��.���Sb��)JɯWn�a$4l���'5��G0t��c?
y���%�izd���ޡ�] ���W$e�U
��7�P�*���y/:�\ǒL˫��σ36��ڍq���|%��9�5c��tn_lXM�6^���!�pK�m��n�p�3~��� 0�3M�ͤj�O��&m��1wA&��ē��yؒ�〔�r��[+Ui�Q�r��F*�d��(��h��km�h��E��O������L�\fgYYJ�7�>�n�Yzx;T��@�����6��Abt�j��\��ǖ���t�J�J6�n��2�鷧U��]����ԗD�F���ަ�?i�<��������^��he�h^%˝^=W���ww�)�R�ej��yy�o(��imq�7�PGX�&Gf�zuӭ�$�R䢰��%� n��e
w�f��=�v�v']p�+*�`�������F��8-ގXy�k�����fnc��Pҏ�v7��։�-����\���Cn�J�wb��,�g:������׎��v���.���2v��jU��#vb,V1r�/���̗��V�����@��FTT���7�&a���򞥐��]�]ܢ���o3\ơ�p'�ۗ4��6�-��u�U�#G��h��@:�����2ֻ�V�a�Ʋ*���f����QqB��+Q@���<�+�
��]��Ԯ���r�=.�%(erZ�}zȬ�������˩��<}��B�*��̇����s�;�nfE
�D��p��������>�Z�7��fa���z:a�/@�Gv�N���pܣV�Ij��:����ST7����-,z�[���;T6�6i rY�Y��i�z��Z�v�����Fk�R��+����6Iopd�̭�}Iq9�'��m�Т�]؆�f$��R?�����QY���*�j[����R�<]mWОUM�:�R���d��YY��e��Mm�Q�I^����r�Gh�m'��x]k�01�S�w���m�����p��@G�S�ƌí�r[�Y��Jb<ݜ34Bp�`�.��3[ �3{�L��!P+#��n���i˔�$Q:���231�2���s��*�{���gI�;θ�]����e��n��g�t�����|�WxJ�^vK�6��/�B��קm-:�3�p�:���W75�!�[������g\`���|5�e��u,]�ww���J<X�{f^�g�xBý`(VM��)�oV�4�'V��v��b��e]���6/�T�M;}|�Һ�.���m\�פ0I�,�m���E�
�1W�t��q��bUs\�G�M9�]cU(O�^p;O/Y���oj,�k��@�,ma��{;��,WV��ڗ�mu��07�Kl�L����Y7�>5�-\�S8����'�Fz�t{>},]�ґ���tfdF�T�[�.
ۮ/׺�r͢c��u��eqx���K[�_�8��Z̛Pրu��Y"�:��oh�yՔ>��O�{k�Ԭ�3�Š>�{J^Sɂ���+a�� ���ktj�t�!%7j�J:�]�Wr�Qj@�"\��z��գ�Ή�':� ���T�c�ynm!|K���0���8�����u���1ހ'sGl�/�����+=��4\�rȭ3�k�f�q��сs�N�]l�فPO6�	d�~چ�R�����n*1�fҐ�n�j�ˢe�dgm�h��9��9��{��b˜�cqf�6��D���;�P�v� �we�2Ly���JA1j_$��6V��&�1k���8����;�8�[י��VͫB�/-��ƀ��1�Er}Z��z�<�$�͵�v���4.�X�Vf�n�#Ǎ�ص\��X��Ѹ�Z�X��]���t�k���=���Ԃ�M��W**e�;�p2j�3\�tqQ��ё��w�i��c������&��V.Ӻޭ)
��6�VY\z����=�`����o4#���Lz���U���,��z��q��0ԃh�#]]wc�6�[�P�9V�"�&�j�`�΢;��b�>ܮ�x�i=�t��,��"h�6`=j�x��u;�����n��q�CuK���g��ד9��'ǵba���[ڲl��`ַY��_b�ζW�(�b��b�\���Z��� B���4�r�\�&f*r�v���Ǒ5��&Ӄ�P�t>�m�Vq_QX"��B�D���D�V.�'�_7�9�\�9c:����&�v��R�<��]��:�4�'Bp;�8iz<�5o�:)��|u�]r4�
�Kv��K��_IE�W7{�����y{����_s��q�/�r�wX;��LGJڽE<y�hOU�����t_KЍF��'j*�E�.�/t-JE���P�²n["=Ĩ���%ի5�/]�Ɛ�Z�������f�	G�U�
M� #�'6��\Q!�}�y�������v�g2��gE$:MY��f�a#}@H�
��(.㽶��Մ�9j��B9�ү�4wg3�7�:S�E�Жi+ѧM�%�F�ܱ���# ѓYє��wc��	�F_mv+ڏ��7U��[=��#{3�{Ap՗�Q�Ss2�cmVP���J!����ge�!�O��#��=���U�MA���$<�-�՗R���V�[�bR��q�VYw�W��D!f��k�(Ė�6t�e*�C
�E{���1]hނ�<<r�c�u��m�y�[dݓ�����A�_l��ʕ�:�DAH">�4�AӉ�M���:ꈒs���y�Yɷ��u���{�����13b�]�pq�hw�2L��G��ݱ��X~Yy+��8j̺��\{������V03rk�YD{Q}m�@�;�]�����)�̕�3��Mt�]e�ˍ�GM��A�s���=:��Ź�R�	�0��MZ�F�Jo���;�7yc�ʕ`� �9d��0<V��v8�d��r&^.����c���:�:A�0� ^��ȸ�7m��{���dap�:�HL��l%�o������umcsFV�\�M�v[M)w���,#V�B��������n��2����ʸ��]�i�-a�"�e�z֞]��zơ�h�RY�T��\��=�}/�;��F�s�+�^���J�p��"H�KJ��e|�ϴܒ
�Wh�k�D��+e��si�i��-C|nz�7�oB�b�%�}{=G���7�8B\ů:m��5�y���!ӈ��	s���:�WR���/��x��r��7Q����;�:�c���w�p/s�V; �ʜ[Ⱦ냂�@��kv�\��;N\��
yy;���*�|�+V�?5���J^Z��kV�֬���Q�+vsF�K���5k4��*9�ʨۗ�`X�W��X�Z�e)m>Zd��A���i�����+��MJ�YM�PVj\��J�U[J�����j-7,ܲ��6[Eh�*Qm�9�4�kKmaDu�l�r�Qm�h��:���-��)m[c�V=;*2��v˹���ckkKVm&��E�җ�f����9�J%�[��U͕ijgj�e�6�3o9�*��˩ǜ���k��5���je��f�iE��ul��9��]+R�ce�X��k[m-��kUFڨ��^]�ζ�(�o.Qu-��5p�Z뛶E��Z����1�g�w�D�w %+$͸������1��E���=M-���4��W72�l�w�䖱�ү��[�c�Rdv��������f�С��2��5���5Cc��sP�B��̸�2�D�q���}y])r�ʋ_�A�5���J��"��
6��/6���J��Xc�g`W6z0��PaB����;f�I�}	l˒�\rǱ���!K�e<�[�B�Ppu�^=5�T僉�#��OT'��w�0e@�9r�_�_��)��B������SX�B��b%�{}̬٘�#&'�@�����j��)��r���я
���d�٬��S{�*<��"�R���2��]*�=�U��3WK�83�蟙ϋ_�<�^�٪���*x�������J�ւ���{@˱u5!��tN��1�mP����:6(��g����u��x���V�M�؎�Ȑ|��(Ď�q5�ko���>�X��0t�:�
�b��TR��VB��H@B8���*㻭��Vɶ�;WHi�$�ېR����B�t�ֵ��T�;�y�Y=�@K]Ȥ$�9��Sn���}p��hJ�v"*8��~Ӄ��yo���h����9u���X�lx�m�7��'����)���&$\���+�J�-I��^�򚜐��0x��=ou'y�L�u�pl�w��Y�^��oG��*��E	tR�917Ս@w6����G�;�KM�(�=D��Y�����M�yu.�0n� iio}�`��lh�5��㭢��Exu��W{U��|�g��(N�ha�zDJ�Su�N��^sСC�]!!U�&�Bsu��`�.r/�z��΍-Z�Y99�|<��1-�֯X�./��Э��%���n������Ն�%�5��^���-���+�Gl%gؖ�k�ڰ��Ů��I�X������EcO{n��B�33.-�wj\���g�����G�4kE��fyh�M`�ו`��\7ީ�5 )������Xg(�8��2s���p�B%���oӖ*2�S����!t(g��l}zI���#qb�n+ʾ���+k����#�"}mi��o�[���bU��>еs���I)��9�Xu^7�=b��\��Uz���Y��H���ݠQB�(
���A�ʫ�:-�6|ʠ��|��6�
�B�t�A�7�:�ƣۼ�p�Y&�q^�C�����qX�Pc� ����j^�'��C���t>��ZU->��(������ڱ�k9��PJ�y&n9An��@��ĳ!P� O�v-MB1�����''g�%�{jԇ��Yf\�v%�_��	���jq��$ϖ�#d^�f1\󑂗��H��f�ޖ�vT��^��1F�����J!=��nMB#c�6��N'ݮ�"v�*���p�l��.{}���-Ĳ����g^�ʙ,�#�לс�*�@�GCBo$)=;���&���|��5��'�(�=�;�6xzݞ��]�V�7U�!>W�>'2+���y��א��|�W�c�<���^GR%>����63�^�ߙ�&�EԱ��I'�a��|���a���*aV������=�vX�ԌC;_Cxx�l�q�H��GE?|��>TFxo�)�R����s�_M��֊�v��7���/34FC���>;�0cj\8q������^�
�t*�V���3�����'�����e�1�Lz㓧�dtF]i���%�[P48p؞&�M�_��;s0%NWP�=����q��#=/�~ж��Uּ:υR�Y�+��+$3�¸�����<
~�q9��;�jL-��t����\1��]"�v���0fOS��Y{�����q*=�����Æ *��>����L$V���)�gzN1p�M�xDumdLj���W�n�bS��[�Ed����A�k�G�Vׂb��@�$q��T��J����oG��4�X�J�Ƶ}���Ltq�©�u����O��V�}��:�D#��떽�6�M93R�4�C�6-�sv-8{= =���⫨#=6��R�.i��0���������!G�c�YxKs7f�ݾn�
f�s0���=��+WI"�>��ȅ��↎,b�y��ު�P�O�oWI�^�i���CG)�50�
�ւi�V��R*���z�'��®ZצJ,�[^�tmx}c��K9��O*�WZ��vpJU}��:m�a�O�۩j�0�<1�>�U��,�r�wӡQل�����^��4+XC���Rcc���\;�4P��~�j�����WqˋԒJ�\lvo�S�/�>���(k�Z1�U���!kf���j��n��aI��̨V!�b�v�\����R��ײ�� ��JZr5�򎷶*-��Y
-ʇ�eG@�*��f��b��6͠����?5��\���z�O)9C2����0���p�]���Q�j�b(N��j��v�xK�	�"s:��3AX�n!*y�7j���T�<��¬�"�R֞��Bȥ��QK70�o��Obo4Q��g-ʂ�:���u�m�u�:JV��D� \F�O��ϝȳ�2��reEB6���=u�+�T/��C+�IɈ3q��Ń=��.[�*o� ���I�/�������D����v&�٨���#L�5�-�E�ldD\s&:�
�U��*�.��T��>GrxvhD�a����1Ħ��1�D�jb����H�"&7<�F����S�^0����m���W�B�xu�\�̅\~ �B�ҍ��n�6�9�i��MYx��d}C��I	 '4g·+�U
J�ZǞ��t�w�"6h^"ʅ��Ə}g�ˌ��=P�J��ȴ�mw��Eb�[�*?�ܛVc,m5�~8a��ʵUj��u	=Sa�/S�2�lo�6
p���㣃���y�):W�P�A�]��j5K��x�ߌ ��#]��Xy`��x�;MsJ�T�w����ͽb�ofn��2|Rs)��l���<�V����zZ=���qm?�������,�\�߁î	��p��H�N^
ݑ�u]CL�K��NR�d�;2N3�g>�����勎��NT��_��[C���C��o�U��{j��|.AKw.)U�yYi�Mb�FD��?�+>>���)˰�9��+��aYÑ"��d����FA��O��[�E��q�*�to���6�A��V��)5�����9���������眘�uТ���Ǻgj�Qz�잀p����ZK��Ux�Hg]Z�9|�X�7��d����
��+w26�Ӌ�yW&�p�L�;'�hY�yV�ٞ�}�ռ-��/��:C�
���C�f�2xu�N�X�V������	o,w�;�l�[	k�,��Bf�<]�B q�iU��<3�~�ָ�
��{Rg����S2 ޫ����^�z��Mr��7C�2�(⹾���h�П�jc�wK���+�Xg�QX��ؘ�h{�޻�]���fa�f�톑5�2�8{��36V��:�BvqG��T���N�=���9�I� j����v<�tv�t\U�R��k����4Z��:_^�e�^]Ľp�j�nFޟ�P�/�p����Y���c}j���ʁ�g��ؾ����c�{3}�u�Q��#��X��W�����I����.C�5�>A������p�b���<��ؼ�φٔ+��IT�`�Q�o*7$c7�K�ߜs���7�C�wF�6xw��z�k����߼���u\��w� bv�/�aB�%�����Ҝ������2;�+l��y��|��wH'�y�Cخ����}�t}�DG���ǽ������q�m�zq��e7[���S�#95�>u^��3����e��ϊ=[��R���AC���T��X�ɡR)M����B�\�
ͦ�.)w���am�Xi����
hź��{T���)��
�~�+�V(��)Pv\
�WLA��(�>;SF-W,9�9�*�CQN1>ɢ�5e[xM�@�U'Pȝ@ �m�)W�b��C�O�w�9ؓV��$�̓*,�t�֋
�і��5�;�-��uK��4 H�ɼ�W0�*d8�W+'P��;�r��@V�j�+�gWu�Tf�Im�s[�ڣCQJ9��_���n���~�I��w�5�@���n|`O\��m��g���U��b��7�6�&5K���f!��-ߧ1�q���!2G���
��箈��
�}J��`�|��H��K�F��˪��AkC�a���)�{P���n|E��G�#��_sw�֏W5��D*�<4p�`���M��W�
C��۾]�	�vƾ{���|������4�
�D�0uZ�c��hl�5��{�.��O^>��PԸG*`N�s�g��Yɉ���`��X�G�(p���޸s���yp��a3�h�x�/�_?�⩧�k5����w}�A�/��׊�(;5��*�-��z�Ç��}9�ð�-��t}F=V�ఎR�|Z�����<`�kFf�(n{^)o����%�O&e���d�x�����k9��n��NT��;� 
�{�y�šL�}�ӄ'z`x���×΢;7���őn?!F���z��X��xx>:+��<9�=��lӢ�nt1��0_��L�>g��÷��gi��J��q��p���i`���Br_t&!��.��@gX�08�\�V_�<���F�hi@���z���[,���X�P�ʆ|lxR�^ѱ����y9b:8XSt�dY�ė��.�z)�b���{M7���aB�ZpUz]=��n�����lq�%�S^ۜ%#:�U{?z?�P�A�o�7�ܟj��t�
��
�|���J�LVz�p4:��]���e랑7���W*�/�T��)[ڱ�w�)���}�o��\E�t�úL��0�G��bl�b/�"�c�"A����s�^�~�a'�ɧ;��bb�N@~r.��,@NLyr�p4���RbH�	?~�x~�1_T�&��G~�eэs�2XU�Q�c7�yb����3�m���c+^q��8wrk)b9���t�n����zY���O4��{��-B �Ʉoo�i���V0q˄H��b���i<�����e(���VQ��p2�Jن�=��V��$�^lW܇9��p�U�����feI6��,e#Ѳ��[e�D��帜Z�pݲ���n3�(�- �?�m�Op�yX:���PݍKq�3�1El��K��1�',f�mu�'f�����_i�:�z"�'hǝv4v���/��]��ҍ̵����q�R�6Q��I07�@)����#F��]���/Ve�X�:A��Kt0��φܷA>Y1Gn����0C6'��`8N�a�x՜L��ͬz�L��f�h5o��"�/=sc4+[8v�(bv��e�w*MЙ���.Cz7�zE�ne.��A�r��{�̺fR�x��`�Zv��0ݭ3��ƃ�v:LZvQ�Y��&�h�HN�I4�#qGxy��U�}`Z%�����?
ީ��S�LpS��S:�Yp{���Pe��[���'�;���o�%l��@�HOupyv�X�!�s��
B�QL��Y���6�n������HuIh�;�2H1m�l�f
>R�S��v�[WK�d�2̤ �^�z���4���n�N�N��`1�A� �vQ�SE�C����!�.��C��{B��d�Sy��,��2�ј9�¹�y�]́�.�Q����w�7	��2���Z��L� ��勥h]uٔoW�ZT��9Һ�����q�V��`�[*�~8Jˎ���\��U��
Iaܵ����JS����N�����|��7��6_D��-�6Q5���Z+!�M;���p�YI	�껜���ҟg$đ���f�	���9�|�Rـ:�E"tR\dGs,���m_�L�j�Z�i����u(CeÒ����L�/]�D�|^9�˦�% ��|�m�IZK�e����L�aDq�?o� <h�s���SU��&e��R�%���Եk9�-Njp�ntg���Q�+TjX��%D�m*�kjPc����J�p�[�9¨ԫ�[�ٔKbsb�u����]W2�"f��
�-VsQ�]����J��feL�"+m����rl�]ZѴ�Q���elJ���l�GR��[V���Wb�ZV�j�klmZ"Qh��z�(֖X2ڋA������X�lm�S	�s�b�Sһ6�	[[*T�3�UR�U��m�E�ҍ��Q�J������9�9�kb��ݲdΈ��93JT�ib��Jֺ�2�2�2h�Yj�U��Ѷ�����=���O�|��}���=�l���/w��JSpjܝײM�=H�$�t�O��gl��Zi�_�WS��w�=�ɸ��dY�qT,t64�����L>�j�o�lJ��:b�AK�.±�y;�qICl����?~�.�xb�����{���+�b�L�ldX��p���GA^�V�UH���w>��髌����u�-.�S�W�P[A��}#�+κ�����WU�&�R�Ơ��]��l�����8�=Ҡ�W�uv�Pvr:.�J�>��*-ó�Ŭ򋎎yB�ת%H�)0;U�t��*q����!0Yz�+v?r������LR�}j�`�P�ƽ�Cx;f��
���E�N-U����~�Ϟ���}������]�3�E�k�*�>0�̽ʀg����)�jFC�J��e4':B'<~�^8� �ٯƪGƵ���^\�Dݮ| kW�U�k��5C:߸L�H�l��к�:�+����E��
�b<p�͈�Ʋm7��5�W����ԃ��6�k��1�R�����x꡵�Oo��w{�e_�D�vW+֋���Ј�:��^g;�\���m��8����.�^�e܋�PTߺn��O���ܫR�����g��s<�g-�g!cF� gE�?E�j�б�_aT�BA�:���vAeZ����=����SW9���T	>���bL��	M��k���Ĵ����1�51�v�O����g��;��V&8^A��k~�����#�g��Y~5�4��0�f��Z�7>��v|-^���	���d�YB����t]
�c�<;����Xm"PB<�]FGX�h��sq���Ӹh	��Y�����φ�4��X�J���5ͼ¬QY��7�D��k:����xjYJti��^�w�e�<Ӗ��k�wNČ�uY P��lI��@[������)���|�;�d�I5|6:�اP!ƈ�=>w&6A�y/��V���⹗�a�-�f��So��.���v��a���6q�5������.{f#Ǐ什�FY��l����;��J�vk-,����tGw-�l��\�P=��$�N.�B/%��y��ثj�,e��Uzc������{�H�z%jͦ%��!����Q��k���i]
<R���"�l3q[��⡹`�(T��z�륯
�OUo��Hg�$�Y3�[�'��ޗ��葪ll�{8�X����z��U���m���5N�~��G��*0#�8W_���:���4� `R��@������\ͩԣ;dz҃D�X�J�]�"}|�+ �(�Cf+��rz��������1KSK<
�����4�Ɏ���,/�������WŖ�o�b�S�ƹ�"�ӳX��ROz���_�1:'_d
eu;�e�|_on��h(�u��b��A���
:"6!]�;�N-{N%��\����^&P�����C�\tLu�����V�^{�����`�G�՗�a�����u:� `R����ᢿ7�k�C���Ǽʽ��y$�e��J&i�Y%���v�zf��������C��6M��w�56w�X�E��y2��Ӽ��x)
*�c�
������iu������Ɗ�V�(6i+W;=��]겝�-yh�����G��0������������t�6}�����<5(�(2��O����;8��v��zh����D�P��0:�c{����f)@��\x)T5�D����T��I��W&Pf�9K�I�-ܸ�ζ����C���bw��l'������p�hu�`�([=ʲXj�zɠ���Bڣ�a�薓��P�Mt�zm�9��yܧ!z*�f�L�J�yjl�o���㣣��~VB����PB6>��~�EN�����z��v.b;j�i��Z!ǎ����T$U!�K�@�x:ӂ�ˠ^�緾)�D��%p�jR�|Պ��K;�2�tj�?=��{��t�VW����-�]����QX���LY�%��^V���o��mn�-F
��Xd�uʀ>����~x<|�ڻճ/$z�v�k7t3v�f�4M��2oHA����I�E�흲㓑ĸ��G��)�߮�׮�[_U�n
���DW�K�*Z�������55��!�6�^��[��́�n6�&�^F�lb��WV���t���W�ศBl�b/�*�w7�}v*��olWJ󵌂q{x��]['g o���6�rc��W�s@�dǓ�����w`���/��(׬�n��:Z����J��,��?�2�����G�@y[aB�=����U{�SUP���0VI��w��ub��7���g��[5�p:s�`�p�Ñ�TY��B�G�!�T��uZ�	��o����a�t>����-:.���
3�LyLtX����~!_��5�o�����~y\����=oig�Ai���+��T�8��GM[Җf�o�덓Fș��4�Xr�u�X�t�T�?�3�~/������W���n��v��������=�חNH�p2���=���m�r�ݝ���Q���(�|mh�ߚ��/�^aٵ��n�\Qf7:2�C'���Z!�T�L�Y���i΍�x����k�_�
��r���#塅��V�X�3�ε}�/�!z�7=ҫ,���B�ngdŊ���
t��_t�*t��]�q���AŇ.�e6&�HFl3w��""d�PqX�҆7鉸[��;к_��[��dK�%�ǕB�B����˳�2�
���#��KT@ee��d��P��2Ǟ���<9����XA�Em�*؝�í+�1*,Ȱ�#�}2�t:��@�
��DG�ghp���[�jM-�'VU�fǬ�`���W��W�>��!C�*$��1mTWY�|Q�4M)Bo�#��m��e�v�j/<���\V���ֺ-ZF�.O�ϛ�3jB�AM�YA�2�-����FuƎ��۠f*cU�SP��R��
7�_��V׺�t:v�*��c~R��nAf�l�s^�&[ߣt�A��P?��U��x��s/a�BV.U�Iʅ��:��ɡ_Rݹ�Nqmv�PG����2���3r�T���{��6�nщ�U�^�Q��ܽ�����G�0u�̑�����ʡ�Y�'�n��Se�<��D��Ď��;�vGG�;���;x�b�!�$(���~`�����}���v���^��q#c��`
�Aؑ�k�e��C�2��*1Nbm�������B_�鯼q�)����-
�`�h�`r�a0d:w��QK�l|��Kmo:������t�F�c�ܴK~ڑ�zU�]ŵ�#1��B�}F/]8f�g�z��[�Y��H��Q���s�3Ϸ���l�7#a�����a�1ҭxU/�k���m�����m:X�or�<\bg�M�@.{e���"�X�h�[���ٟ6�q�d)�<KP;cʌ��<+W��}>�-viU^@ۅ�][�v�,�n��:�̇�Cz�Ղ��ׂ�H�5x<bЯZ
�6������[�zȯ�����:ɻ3QS�˓��ٱY�eE��T?s_��]lN~��Ǥ�:�e��!&��^��k�d$�6�ԏ���Y5���澽0ws$ȃ3k���[*�#J7�7B3���{
�:[d�{OW���r+��m@�3��`TQΰ�n���r�N����r]�E�f��B�x.A-�b��Ͻ�N<���e�/���4\w#N���;A��h���Z5��D-:
�cC��d����Z����1�3��z�)���.����6*Xi���Z`7�Ft\F����ϳw��/�V�ҷX ��@�;��7�f�bY���9+<��h�2�b�:��8p`�X�>p�T���ћ��kNn�iש:�Ԩ��?�iXjQI�t�W�kG�����F��X٘���-�ߢ�
��Ӂ�O�'�F�����G�bt��ǃ��˥jz	���]�\¡��a�9CHT�u-S�ߝmhEeb@u-����+�g	2U}n,d�6{`ߎدB���mH�ǌ�T��}���u�U���Z���k�M��DY}��5:�����qV����_q��\�tL;ԛ|7M���me4�tџ��,���rv9q�2���+�� 
��g(��%��
�麟Uy�랁�j.=~y)��B!�DTg*˓e���~ɥ�X�B���j�||+*���^uY��VmX�YEvI"=�$C�\R��{�x:���B�x�r:��$z=�f�Mjކ�$h����琱a�SaϚ�Tǡ��S��Hr��xJzD�:����LD�;�
2P�@�J��,/�K�2�J%
��[���V�#��`(~�P7ENt�!@�U0`("A5C�gWn�� f��-+�1���}�gJt�c��0Wn���}v�oމ�`��qfE���:���+0p��'*�}�5]��fk����ȋ�;}��om0W/��E���-ڃ�pp��'�>�֍��c��f�KgNr,祈vx:V/�\	��b�^�&Քں��*�X�|�I������Ƞ�M��3l�⟼�����G�s9��b��S9=ס;1�"B��:�Y��5MS����H��i%�-��T��S�y����SvS��Q�Ml��ނ��?~�����kJs�J���t\X��U�aÇ�)Ã=4+y�:�����{�ZE2�h�	�=���;hR��+D���]
g���b�Q�n���%�o����A���ߛF��V�Z#����ĶE+�g3wQ̼}���2�5Z>C|��h�?�2�+|%�/+`�>>嚝z�g2Lrj������჆R4Ƴ���7��J�+*8zu��p�6���&z�ф�m�a�P��5�s;&.�ƺ��\(	�஘s=//5�K��2�aC�t8pe6&�B2�|\h�EI=C�{���>��N_�}|����> (��i�
ϽY3'l�<B��=x��
æ;�3�J��fEX;C�d������a�ݟ����8���򀢀eV�='輫�jK��L8��Z�U�����$����>yd��@�Y�z�=w`fN�_Y�����VN�fg���$Z��Q�L=��:=[�~�.�c�V��ꐬ2zs�:O�!�}�9:d��K�� ��%}C��8�Ak&�Nya�z�$���Y�+
,Z�Y�������}OY3U��S�	�����k�3�V���_F��y�J�Y]���T�E������2��+*�z6+��3g�J�$gf]���f�|-�l�ӷ}ԂJ�aR���{�I&�Y�2��u��pC�k
�Mͧz�^��a�G1l�+�l�\�3���q�u�$�F�����^���ש�/t��5_�U���6+,�n���5hJe֒�c� �gדkж�C���C]:�m�+7*��eڔ�[���*�me�Kfr����i�T_>�/�8퍐�A�a��ӱ�%�8�Kˆ*��"As����=9��u=���/p�Ѧp{]Z꒯��,0u�z98M�P+������R��k%�4�"v�W7q�¦Y����$Ю����MʹS8[��7��=��S1,�U)V�v�!�7�m��у��f!���}1Ef֪wz�ـ��2��Ub�K�{	�uk��.�Z�u�m�c���_��q��ۊOV�!,�抴9�;��J�t�Y"�L�����8:���Cie���9�ЬS}����/Ș�%�/�c��Cǣ�^�����sm�ei����+�Ib�5eH��]a���cl�9:��ȩ:�@k�*�jR��O�mپ����Z��ije�:/���ۺv��R���p�8wmZ����ڽ�U��^Ť�2�6��G�jO��چ���ٮ�G�����V�k(��B�l5����Kz)����D��9+�m�������M�ݼk֝�[Rr�ʅ�������fJcP((�X����f�N�N�D�͐�Kn�s����B2�eh/�N��|�L�LC�Kƅ���}sN�	�ݢ;`��h:a[U�B�w�:��}ٕ�z>���u��T�q���������pJ�H�)}�{Me%]܁X�C'-6E[ޏA�2�/ ��j� E�QF�6\��'��Y�����n�t6���9uC��C�n�~�\$Y�C���b4Z�XC@Pݳ�@�$�X��+O_w-
�ݘ��2�v�cV���W�F��f]��~�\�R����B�J{F:���b��v�yE�czqU�\�NQ�������+�~�߿����бK,��>�S%m�(ڝ�����E�KP��*-F�-��Uֲ�F�U��tp��KZB���	h�%��m�-����9�Vۚ2�T،F�mA��U��+�J�V�Ҕsu[mT���%��4F��ҕZ��L��l�m��e2�Z�-�Z�Z�M���e�[KZZԶ��Z��%�h�+R�eF�)ml����iF���d�nśf�ΥʻQղ֖��m��DikZ��&�fkKZ��o9WR��ʩF�ZѩF�KZ%`��mR�m��մX�h��m��)���`~XB������V(�ʇ���q)�ay�Z)��Ó!�K
�b�W\بF38��~  �E4r�=��P<t�*�'��8�Y+�}�C�J������>0�R_�>�q�Y+<I�}�- �2p��,�� �8}�q=g�.I�t2Ag�?_y�<��~�����o�E �����+�~fa��hd���9��fd�
)���}C�y�ɐ�:��>��_|����+�>��V|d���z�"��8w����߿wϜ�翽���x�^2{�8���=az���Ag.�w�
)8{C3�;r��A|@����C$?n�}N�����TȡPQp�ª��_P}�pRi̘}��V����^{�_��0�{�&g�JϨu�@Qg��;�2T�����
þXd��}�Y�%~�_Խb�2W���dR���y��a��9."���b�4<����������l��g篿q�:H)�<d�>!�� ���&@Qa��Ι+'}ِ���R�T;Iz��D{�ޘ�����W�)��w�(2<!�Xz	�d�Ԃ�}�*x��\ξY2Ag����X>���v� ���<fC����'�,��`�j� ��l���Z�-��U�~�|�O�w�Hzl8��
ä����Y�&�YQV��ɒ����`V���s�B���q��Tu�əĞ9'_(d�����O��h�����_Dx0@���ϼ�\x���C���IY�;O���Ad�8{��RV����X3�%gi�@Qg�:L��*C�S�
�`V_H�� �;8�L+��.�x��y����>2W�%�<�É�2W��i8�A3ԛ��q'~P��� �n@Q`v���ߘ��AC�Rg���?'�՜H):�~d�
)�Oϭɻ/�=�����J�`��J����t���/]��3�JΏ��{������'�@�+����ϧ|�8�Y�����@QIPL{c� Tx�����@����#��wOh�[J��f�ٓD�cY5��L�t�d��k	���k�v?Q�]OG�;����<��Iu�I��Q�c)`��\4�<6Ф��V�s���DnF�+��xx݇�Mn��<"��1�aR
����+'���R}B���O�)'�Wǝ��t��
�߶=@��g�q�����~�퓤���=�c�G3&�'��П�/���0�����@Qy݁�ğ\�IR�E*����`~�r�Y�}a�ԕ%g����T�ɧ�i����
<H���zc�rW���7���|���E���6��%@����~@��
���O���VVJ�a��p��Afd���������q��d�V�P뽧X���ϝ_|�|���߽���Y�*AO~�3��hfO=��Ad���E��T-��³�Jϳ�L�I+ߔ>wa�
¡�������>���E ����h��0<e����sW�e>/��L@���!��$��=��=N�P��,񇉙=eH.I�=��<aR
~�>���Jé�2):B���>�� ��y� faY�>z}}R~̊8��ݿ@c��9��2����ed��偵!P��s�B��wC3�����YR}r|��$�y�4a������Vx�|�κ�o�~��ן�Eĩ�w��ä����3����2Ag����t��~�ə�*O�t2v�\��{N0�N�+�偙�!>�*������|�~'}�?~�G-BVr�I`Tt{�#�}SQ��'g���>����^O�fqE���x�B�:?lA{a�;gL2Aa���gL����ö���HT>$�]!�'텟
"!�7}�}�tx(��v�����s?0����>�qOZ�_�
�3ǳ�H,��x���
)����a���^@�s��	����b4��G�tU�%/��?2������Ȥ�
��:���Ă��iǧ�a��~r�L8�+:��'xʊ���g�J��_X����C��B���&g;�D'���u��$S���m7m�3?_o{��P�Aݧz������ʶ�s0`c�Ff`��-�OM��xt��pw��)�%hY��:�M��@���������չ���Q����	���w������� �������AH/��L��>0�>��d��|O��t�P:N^���~a�*�����}��Ag�:=����%H,���G�1�F�F�����K_��6 �=��T񓇗���W���x�$z�򓏬�Nwf0/�~���AHkOǜ�:H,:C�����$���'|��~Q���;Ͽ����!ā��C�w@��'��O�|ĝ�7��>0�Y�'��0?���v�πQ��<��p�e����+�fx���y��0�2|@��|Ꭓ��T�S2x���:<� ���g}w��t�R>P�����?yN0�§���x�������c��G�:�&=������
<��0�/�B�H�����T�̇;��I!í�@����>u@�%g�����
=��'��� ����_m���?vt�Ŀzc�
==1�G�8�Y��Z��T��+>�Vv�\���
�ϝ�q�L*x�C$v��n~�z� ���L��QC'�6<�>&������~�����'�T�Χt��g���X)�N����L<aR��������dXt³�n�q ����_X��P=Y#�c����>8�_ښ=��k'�d핟�*,��7��F�OP^��������:���=a��R
Ar{��里+��̟Y�
�AI�
�w����׿����w��N�=�����0�P�8§��������|;���*ԙ�^�,�<a{�>�x�Y�Oڝy��xDz`I�:*�G�ǷZ"���|�����U��{� �x���{��$�<}d�S2q��J�AaR>O�i8��Rv�g�����nH)���Za�>���}�s�vș�����U��W5�]�Y�T��B.)	��e�`�������ٻ,_t�Q.�k���ѻ,�@	�.��V�+1�&�i�y�s{�S��̸j��իjR��D��ku8�~���������~}���q ��?��q���Htsi���*)�򁟌��i�:H(�9l��O��������*A|a���0�*)�+%~T���U5u��/��JF߽p"<6<&=���$>'=�8�a����/�B������}aS�C�Jό�a�H/��OY��
~-g�=LÇvdR=a���w}��u����z}H)��9'�tÌ+:�Y3'�Vfs�@QI�9���Y2Az7y��@�>��8��I��Y+^�ܬ�*s�>�+�=?S���x������;Ob��yG��	�'�� �2c��p����$�� ��¾�Ua���q �~J��1�}a�E�9��t�'�'��e{bç0�¤�9��_�{�ξ�~��x�P�{C"�Y+>���H)�'n0+0��`*Ag���?Y/t��ٙ�%}d����g�6>'l��X|�Ü��*������Q�Z�9��_��1��`xD_��}C�>��>!R>�����XW�����Rg��a�wb��>&`sۙ����<��� TyG�0"=��^��ޘ�]��π���'����> �!� ���3������Ӥ����3Ğ�0�¿?X��Vw��I����8��l���Rx�{~ g�9����{ξ���������°������L��+��{�V�Y(�^0/t����0��uϺ$tè��@QHc�N$���{d�XXv��
���|�����ܟ��t ��S�bq���RVN2�1O��8�l+�ng�J�*d�q����R
}a����a���=@�:\{���"c�e��M|�s%���}��=+���9� ��/>y�v���Ag϶N�g�,�=J�Ƴ�)�H)�޺P�;aP��&H,��C�
,<B�;d�>��������\�{�l�#ߢni��*a�'����~ը�̬���>M��A�%s��7	T� �͏f7wK{����C���8���,Ë���ݪCm�r�_�:kRZr"������(�RL��0=P��2�0�v����8�̕����؂�̕>�mYR�O�OY��>%H,�i�{��R;����
AjN30����w�������}���|��'�W���'P姈V~�ə:�fI��������VT��3<d�/�dU���;<������0+^����q ��k��sG���f�ظ�� � �H��'�^}�3P*�r����AI�z�����J���Y8����&a�
�޳3�J�un@Qgl��s�|�����AO���紅a��y�I��:�y�N�+��JϬ��Y+��9���`�N{a�z�$����x��έ���>��}S T��@�5���3a����X �Ǘ�'XT���2V�}�C�
��`d�ug�C�K����a�}d��_y�m �2p��,=eH.Nl�OY��u<�G~����￿=��X_)PR�퇉�ACԕ�;fa���2Ad��<ی̕E9<��:g�l��T�'�+���>���+�*z�Y�%G�<�ׯ��z��{��^�����d��$�OS<`V����2Ag�v��@QI���Iې:� � Uy��p3�����fO�2N��E���=C��u�/����{�8�Y;ez~�I�t¡�%gl���~��
,��|�<���o�c��֡�sed'">���+/S,mPՏ]�V;��_���P=6/�ڃ�\p��Mv>E`�,l��Y꯺�*�¦w��"1J��0+��f�ͱgbMV�6�vG���k�ΥWj��\g�ݣr��%^��̆��;a8 �(���fӦ��|����ӵ��
��1D����j��3*IE�;3w����ۏ���.zč�s�����s��f����kIL������|=�{����K�d�1Jrn|�˙��iX�Gs��_yp�kά�;��I�0��xTs9�t/���ክؽ����~� ����u��Ij��eÍrp�^�TӬ
n����_`Gr�U�\4����
7�NN�D�m����c\��6'�P;^Al%F�]T=m$�8�������t�����v�˅��f����*�iXؔ�<��u�0h�	���tҙ����ll�[8��t�����K��̫�_[�EhW�`��#>�<=�薝`3p���+���m��i,��1.�p�7�*TMp��04@���.�j��'z���/7�u]���f!��m߮R�O8����0u�ѝw�MF�1K��(!��pOW��(�"����4����U���as�r�4J��z^��s��ݫ:K�D��^��9N�\޷#��7bD&q���Յ�N�G�V�n����v�2FN��Yy���Yv����F[|�k�Ծ@��N��x]V5��D*ӱ.jb��꓆���or:ڣ�؞�b��Χ��:�[��*XXU����M��~�Lsݾ病z�u�lHtl��������(l'>�FH2)<�~zL����}�ɈAb}Ƭ���g��t�p���φ
Ѡ����s=�+������ܰg�Hߝ�2�Ff���xh�JV��,/_fY�#|�=ٜNC�d8�����6�₣�����J���B}��R�Z��Y.(�c�P���
��੹��PaB��f�u�<z�;[�4D�ǪB3�'�W�%�����.�ιu��f���q�1��Չ��"àp���*����%Ƴ��a�Q#~&��>�p�C�yCݜ���K��!�P��*�����xWv�����;<7�A,o�,��^�v�R���zw��5�D�sx�V�_�cGW�ξ/+���p�^���ܫ��Q�vc�Z1����:�J�x'nʪ�����a��획߭࠲��7,@�sjR�
�EbS�
p�£!vil�f�8�-�@�tCb���9�V+�}ڋ��D�6&v0B-f�����-*Zv�9��
ZkB'�����K�K�(Dd([�Q����	��������t��]ac�<�Yć��m
��C��]7}����O��$�F����y� l8b!Qw1YX�QX��Ꚉ�yvl4���΁���9+��`��(����^�bE�	��+B-�9�o������A���Q���,��
��p�Z��ޣ����q�
�����U?�s�+���NO����e��6�b����f>J�`=�QnC�r�踸P*�1`9p�Ñ�TY��D��ҞO���0:8C���룠nmx��T�q�Xy`���s<+����IF���]��{�gL�{�2��U6Py��O?)\"u�����̛�!=!B:��i�Y�wum�rofRӥC��k��qZJ��uO���Y�F��{�{���i�d�hu��pM��/���l@mR��υyg �-[^\2��Z��Q�L�W����Pt�f���ѐW�]'�GiF��%4U#>U)IsP�����]q
0@�4'�rb�ӁݼN,o�#39&�ݽ��S�ƞۤ"Ð��gdŊ5�݉[����f��r/Ƿ���`�K�С�H����˙���Nٸ���f����)NB��^�ȧ6˃���E�t��uPUt�A�[�ob��4��%��.��DL���(�a:{#
����;�1�[�����7�9��x�m�����!����*.�*��Pc�C����p��{��rFGl�bd:��ErШڱ�S2 ܵ�GxQ�z���x�Sq�׺K���= �P��b2�R?A�����V�p��}Wx z<{i�%����$ɲ|������v_��y.:�z����Ѱ�J�r��='V07NE�ӝa�#���+t&%S����Ï�=��q��5�r���}2	%{��s���� {�h�'S�6}� b�]�5R�t��t��؉4�m/�L��
���ɺ��6.:�k"�H�X���)��P=k��\,`�Û��d�M�2$~(S�Ѷ���z��ee�7+�1}�X�l^/Y^�6B�_��^� 8U�4`v
�d
�JBo$,u�e���R������Vk��%���B��/�C X�`�Ӌ�Ь�¥�GxX(� �ڱ�<VB<�<�����3l�4��t׊�"0i����J�#���z��.��*:5Hq�}�YT�ە�I����U��J�0Q�%=' ��z�iǲ8�q��=k� ��Cbp�j([;��G6��12�n�Vͫv(ޑ�s+����\#���*3NxK�v{�wh�Z^c?,+�F��G9��g��~���H��8�L^X��{�6<7h�+��a��:�f<�(�k4,���&0�F�bC��m����d�X�tV�)Hn��{V��u��OA���3|��J#P��U�(AarJڦ1���U����7�V�fq�m�*s��pste��v�V�4��d�765��o���`F(�6�
݈�'���f!8�P�:Kxj�_`�S����F����Y9�b��;;���1P����Q�K��3mg�yJH�;�ej���U�\�F�6�KVh�Κi��v��֡{��T H���#Zd�P����Q|E^t��tB|���n�ô���<P�Lܵ�h��*�֫{	�t,�s7ķu�TI���-
���IC�+��,r������e��*z7$�^:��Qiu���+"�����$�&�m�㠴N�j�5��@��kM����"9�7>VrLn�u(W��lml��;|�@����9�]��B���I��y	�+��Z;�&�����E��v09�r���:��X�$o��j��q��Eek�Q�!!�g�N���xIp���;ת��-��V�������;oP/�׵���k��A��)��B�
�1�l�rfa�4�����K� rɲ����,xͽ�uݹ�	d�&�������ƨpEf�G�;p��T^�\X.
�%�W�(M��r;ġ-�g�P���Zq���
r����uf���%r
+=�`+���<��ūMY���+�a'�%�W�Ol(�b{{��\9%|rd;��h�H����c�WB�]H*̋�N����Wu���Ǻ����^;�d�x�:���y�]G*Z}�G}/���7lՎ�Y�]�ˈ�p$f�Y�{6�Z�XL���b�	�f![\ӧw5�yX��
�)Z9�\R�̺WaD���^4A�5j 5���eЂ� ��@��r�r�)���S�^|�	g�1�癶�[b���������om b����5�$��@�Qd�+�ot�a)�f��kX��ف�ژ�5����.�m,h8K�Щu�)wg)`� �A!�ł��k2
ȓ���(�7w��O�|��Þ��`��J�EV�ѬN�QG��(��B�m�����Q�36R�����[Z��QY���؋mqi�Q����-��m�+Z��.B��1CZĸ���Z%����eEkR�R�U��b"��WZ0Q�^;+m��L��ZZʪ",���\���Jݮ�EU9h���m\[��v*h�<�s�n�QDF&El�kkƂ�a-��283��9�;�h����"�j��C����֬�sn�9�q��q8��.�,U��غ��ъF--J��U�����s�Y]��˅�h�*U��Ѩ���7�iJ�ԙ�k^V�T4Akm�r�)(��Ep�w��9�:�k��v��:��{�����N��|���60m���3gu�4��im�;������"
�ͷ��U&A�ط^7SZ;N���	>kµ����}�S��Ɍ۵ӝ��a��-Ks耠a��mX޿���`�M���}��_^�����7`���n�bR�O`_
d��Ѧ6ZgS��kB��w;=�+�����ظ'��� ��F��եi�>74P6�TGZNA�5j.���bE�ӓ�3�b=AmZ���5��>(h'+w�7��_kE鼉��9��@���.��!�����[���L���E	~���Z�:������*�b��^X�m+F���U���'���R���{��n���8�`��X�����]J=y=:̧t�X]Q��z�B�)f�Pg��ay����6�%��6�P5V"�h<��f�בj�����W�>5��� ���p������E���WJ��=&{o�>�Js�&�Sݢ�Y�>Ӣ\y�<I͡�лU���J��%�'��8�d�L�r��P��z]<ޖ`o�ة��/*d\��9��Usy��(i�Z��}_ <N��[k!!'� tg�C��CcǇ�V3�����\/27���rw�z�{NS�-���ap�O���/��9F�p���C�J[<}$�Vo�2_��^
�,�a�H�c�}�I��e3в���YP�JI�oz��j��dT��E�p� ���7
��m)��w^&O��`:��sְ<�#��"�ym@��=�T
�����g_rs��*�n��
t���KSaϚ��E=���5��dvYG��W�)�{��PDL4D8�)�-�X��ebV;�f!g�ͯN��2(L�pu���6�9Λ�"�
P�b���\�V��UX����Ȏ����q��O=0��F�Nf-�F򇈶Nd�G����D���9>��X8g�Ag�ʣ��Q��ecy(������2���_���<e첶vԅV��T5h'㻗ZLٮ�0_V^B$�ͅ�E�L�v���̤�lj��S�N���M�[l�uJ�I�b�h��'~}���U����e4a�˹����㠮_E�i��a�[��G�N<����4@��ß�閬
4�t(�N�w��U�d�lf�'�!�gg/In����NgWE�n�3�PʴȰ�Ër:,`�݊�g�CV-� ��`����me�����k�+����*���n����ZRLX�5곃�m����,}��mY\pJB[�Y��n�"<�\X؝�����1�l��^\9�����<6�Rx��sJE`)u�د�.��4/d���tx�:�4/��	A
�]�և�S�G{sv�%���U��.\;5�����!�!B'�fvLX�����i���r	ήS�����C��C�Ը
����ǚ�����G#JOs�?���h�(X�]C��<�@�.ƫLʓ��]ɬ-Gq�XB�K��X�v5Y�v�9��L��wu�[���|�飆���z���-}%��t��BS0�l������:��9���u�)ûNK�����z�u"�&g^��\�9H�uu'7N����꯱t���L��*���$#J��G��=��]e����k�w�E��Mol�%�{��>���R_����_U!�W�-��签�l'�T�w��(��C�t�=�lm���b���O{��1�v��,�$f��u	�*`�T�v��r��g�d��`O���$�m��6��xQ�r�j�1��1�AR� �)�o9���
���9��O�R���<�Ac����S�U�f�E������Ƌ���+' ���^*�i=BC\9�eR�;�sQ̯q���27v[����K	��Уs�:4`vU�Q=-	���w��]"�8d�����CE8�����f���FNZQ#�J�P�^�s�.9��":��>)i��D����r�eQ��"ᩔ=`۱{i����W����[������ȋ�p��n��
��}�5��^�n��K2�;�&r�Ί�A@b�9I�m���ŝv��SZ�x�:�{�l���r�r_���Ks�ɷy�ؠn�8QюB�s�2���!|o���6e�f
-�:z<\��S�>w=NLl�n�t�����AC���dp��U�W<������~�:;g�X�w�cY��dV;��\��g(� ��f���,���ʰ�.���seB���\&�!��8����TDzyV���Ehuڰp��H�
�ʔMQX��Ot�x��nn��P�=B�qu�/���(4Kj����ǔX츪Ӹ���J� (1�_��/�W��b�]y�,p��h@)��wj�ڲQTJ٨�4)�8�1�����+j�#��Y�zj���T�?����5�������Z�}���߽)�j��l߈v�,Wx�&��+�Hr������R#oT���O6s��*�j/��Z��\}�αHČ���ݴ�LzŉWE��Y����u�]}4TI�q��o
t%�N��[�X�^�sq��v�V��)��s�P�Lٔ�����3VM���&�߼ �c� �t{�����1a�?W��?�e0X�J�xAcݴ�B�vY6y�;����U)P%�א�FY��W�vp_�Ұ��6���ӫ}$I�����^A�m!��2���
34~�f�F	��'��J�|�����G�utX��V?*��4Wƾ���X]��i�fP��,�i�h�GM�sTO@ۑ�Y!��:r�E3[�À�X���L��g@�cd�8"���H��rE[���Pm׶��Y�Q�����ޭPpu�/�W��jX,:Eak����@p�V��J�x�ez%�ߩ�#T!�n]J�c'`��C�ss)�
ǈt�,���Y�%ˤ��1�����S�N�����j���#��wE9��R�<p,]�NA�lP�-K�51�y��k&�k��7���6���d{,ut�|Ǡ���W�0~$���]M���:�-rU�}erU�k��;��ѕ%��L峍��;�3g]�����%��p��D�A�+���{���4��g� ��Y��=�"����2��PD�c�H���L섥�W��vDD�烬(��2���p�X"D�ܺ�ηZ{h~�s�5�]�F JT��>v6*�[.���׆&2��k��1��*���X9�QV�l��[�b,V<%Y��]LOw�}xY[��$8�ǟ:�j����N(�Cmn��=�룐��j͉�wf[�_�n��>�ڦ&R�t[Wo�w�o���^i?w>�>�X�u�S�
�/�j�X��T�`Źp��H���|$�h4�Y�:7���L؆*A�"�H5����B�+w(��'�fMiYx��~�}P;�:�3O����F@��	n$u�_b�����9��/$�z:*�P�Hg�j�\5ڤ��:�/��p9�
�%:)s;S{1&]
�-:-��#���z�d$I�(p)M���ژ������x�2m�/,X1p���y���yzh,�/��EY�����U#Q���!ة��|���q{x�����)p:ƻ�t�T��������@�}#7��<���y�+Ѿ墟��r�ٯtV4�g���h(�a׍L�Q�#+<Ng���jϹ�C ߤ���g1�=;��t(p���g.�c�<$>E��G��-��/C�[^����ˇ�\�=:\�:>UZ�����L�yNvʱ���1R2"��bۥ��s��Å;�⢝�p|�������W�V��c��A���"�ʣ���>��kӧ���>�|>>��	��}o���ݰ4 ��ӫ��kjdl��V���;��_SBl
���=��b��/��'���OS&w��3��K8 ��TUV*��٪�������\)E/�e�-�v�}pa�Q�f�J��Hlī>�}�P��P=k��40f���M�z�G}�:�:b���cYˠ�OTݳ���\� }�br|�1Y�4Gv6/� �i�a� �Zw89�rtfr�v�}c�.�f��7U��yuT�E����{�XQmX�Α�ʎq>�t:v�*�xu�R��ܬUY���I�>�90��I�e��g�֯W�a�#�]+���ʛ����j��E7���JN��W��V��8���&�S����
V�!,��{5s���g��n���ę��dYTrpȸӞV.��1���?����u}WFzү��B��1�ˎ�rp�^�T۬
j�k�����d���/�^��㦾c���(T�J6;g���P�P�^�R!�����rYT=�̥�B߮΁tR��z�}�����@�������~�.�`�~�\6�������b���g��/�VNH�[pb�����r�+�!k���j�n��Z5ТD\`3�t�l4��;u���[l�t{�o*~sp�O�1�q{��D�
`�h��ˠ� ���Oej#g֬�w`�Q døD�Hh�U`m��K�m�c�Nv�z�����[������S���&d��o'wO[Ρ"�*�,JjW�LS�8��{��J����Wv�E�ۈ_	��&T��oA�����54��ͻP+I��z���y�y�<�0�W:�V��"��K=e1wB�L�d�a��ہk����}/�T�X}8 d<��\d��e�&�x�ʳ�A�n;�y�u��=�F:8�ϖ
D�}�����������q��Ի�"W,�y�e��V�c¸���Z/���(`�F�x]p7 ������j>r+�>��/�
K9�����5����lbt�:���gl̂��ʵP�z���O����o�a�Tn�]5}#����֞I|����m�*=!:���?��h�q_�ث��-\�8�5}����
��?�.�&�ذS�
�ʬc5��^oGN�܆��ڽ��~���EpdX�m�h��p�O�~_X��������WS0�)��h�o��N�;��R��K;�*����d�Cz�=���n��L��wW\o��r���Q�o�W���,����t!\�
�.�3.�f냐�5���/.��nZ�ݓ]�W�eM�aWV1HA	T�A�C%ޭ�p���L�}���X7gK9�#ʽp��S'���q6W�_0,�F#����V��5S�#u��D�,@Zc6�k�v�u�r���v��;�;8Q��1�Z�J�Hᤇ���ș��W��)[c5��յ2�^A�E�+��r��Cy=�,�ie��ZR�ތ���@6��֪���B�q��nV����V5}aN�R��6L��Q��c����F��[#���
W�4�L���ij�%����Rԇ�;��t��dYj���+$-�oFܚV7{�X�V*D�u���me����ԅq�F.����2��fcލ��[̎��V,��!��~�	+���xڋ.����m˭R���trӚ��Y��k@��zݮ;vx�_�6S���/>���Uj�#�U��n��1��Ü��/��}[��6-���:�X+(���+oKz���U'>�EWQB��ܬ4"���|�!���ל��~s�$����c.�+�QnY�yQF�.z�����J=���W�E3�1�]u��$�5�~��XnBZZ.>+i�q��&��R��<�Z��P���&\%��j;3(���5�L7�G*�H`�թ,ӫ�ܹ jj�;-��7hL�J�F�e]٘�^�5����}�y3�B���Zb`�yr�d���2���U�$E�� �YU=(�)T�s�a_� ���l���k�`E
���o��ނ����	��JV8R�r�	�f�t��1J���ى��*]�M��X�m�ʭ��/,�,f&���a���L��%uE�9�Π���/1��EDq�E�N��_n��J|3�=3b�\�m��Y�)ͥ��%)�.�^i�T��Hm

���Wv��8oA*��F���>��{��x�J?X���ն���Z�J̴��Sk�eKZ,ɱA6���-��E�Z���ث���kG�Dr	h�QV�m�k�Qr^c���-�����SjUւ�h�.�;gR��FҨ*�J��ت�����#j�bV+h)X��k��\� �v��R��Ջ��-�b�֢s`ʔ�+[m9�j�lC4�[E2&ڕ�&.\��YG���9*�y�isso4� ���3R��[x���QS4�7+-Z�����XZ�֔���X��U-��!��/��V�Ͷ���R���QE7.��r���94��UP�ԣj*��b�)�e+sh�Uj�aK��<�{�YO;S�a�NbCsI�g]�u�;%�8�\Zui3zR�Ս%�e�6a�z%�~���ܺ��I�i5ި&O�V)��!Eb�����b�Mt˟S��Ά��'��ɁNP��v��K)9E3@�i@�͘���5p��'��z/��\������T�%��,�#���F��P-���q����G0�����܉P���r`�ŅOyϚ��*g�в뷹�[��cWc����-��t�H��f!�FA��@�
��ҽ-3��d��~u^������-�mJs�P�"$gs[)򇸡�6��#�k0k�r���բ�"��Pv'b���j��e����?t�As#������T4�����X�lRY\!���wϜ��Z�D��񟼳���\�|t����j�au���5#�8�R���
FVу�f�2�r�'��}��2I�K)g|�@d��b�X��ک:�ty.��Ne7/��nXWz���v�Z`p�a;~�Yz+�yme�����2��[�+I��1釤��])�peBl�
�X�e\��]�q��i]��� �$��w�}�3�QQ����p^��Z�`a�ʹX��b�̿l�r��� �X�W��P�(\:��=��,t���^1]�J��+��+��ai�x�C��:�̢�w�g��k># W�,d�O'
޾�Rϛ�\��ڽ���2�h�m�-����0��\ �>{�Ez��KL��诏Ӓ�3�:�'�`�>F��3.�7 ���tNz���u�w�/�׺1�c��HC2H�^/l�S��;������u>�>��=�5WF`��Qb��r�+M��7�N���1��(,8O��8� ��U྇��5:y`c�:QX�t�q���K�4��;�vS���j )���)Ƨ�*X��� �%���c��D(b<a��hĜV,��@���k�>�!f�fyl��"e�E��)����5�;;q�o��ùT�b	���=J��s���ӷ�u[���%��a����#IG�o3^ԗ�;[T��t	q��!5������Dj
u䮾���ˤZ����=��y($�O��sh~t�_��*ҫG�xa?r�~��hf큡���Ѵ���ܝ��b�S+�@���K�%7b2�$u51���J�~���/�f��jó��UF����Fq�A�[�3W�߲'S\K�0T��a�*c<h�ʅXvx[�_ux���5Y��JUױ{�Q���4h��W��]yV�2�P��:Po�]@&�9e�P�g(ƣ��sqё�:qѐ6;�с�"��		"����Ϣ�=�
������pt�V/c����NO)1]�Q0c`���Rt$�ť�����N��bT�H4R
��`Tg*���"*GK6�*��U�S�c)E@pcj\8q���(����ZtT� o��h��:�z�b7�Sr��������4�;k�R��N,�#�<�93J�G�HGSD�'�eܫ)����i�@;���c�ڣ�im�:1Ō�����}X���o��t������?����?}�g毆��J��q��-���C��,�xK(Q���p�4h�U��=xL�6�T�=T��Ӏ,�:�p������G��+<o���kt��iu�-����]�qPQW��.�лV� tx*|��-L[����~�c�b%�X�;��z1��6�D:n9���9�f����/*�t1��E�^�����W���5:�W?+�gz���En��2����k�mx��Y����=b���t����q�ʽm3sY!�=9.d�X`�:E�w�?����b��{\�^�+�b�kp_��lA���,���٫����� L*ɯW��a�*!
�N�s��f:��슕i��B�U�E������9!�;	;�;�飏
z`=;g��tQ�g��𱢬����l<�6���vׯ�];��5�fy�|p� )z����=�S�QG�R�oQM�X��;R��%OѾ�E�~9��5���Z��*���,ç�i��j �7��M��(q�˟�UU�5���=���oז�__�_�0��Lߚ��s�_���(-3�7#��~��R>��?H���=_:1~&��\;���?@����mbA�L��G��"�qw�V^S�[��Ј����S�XY���Ɗ��3r������ّ�Ό8p`(�ƔU��b"ѧH��p�T�����Ws��8����)|l�S�V����dʬB���{�n�yW�y
Hc���E��n2�������{^Sr0D�L�6ҏf�01�A� �Og���,g���
Y�ca���d�NX� ���-�ѡ^8\[��PE�he���Q��A�R��-���Q
d\`��I�)�iu1���1�# ؟dY����P� <)i�j���hih��{#�=@���t�u��f�(V{p��~Um{�Vr�]�L�1v��M���5�-`���D���]��f�M��Y��CgZVV�=�;�\����<4���Pb�qUΧ]m�5�N\V[�+��gWKi�9���[Ğ��{��nC��bp�a3���1�=�H�w~*���A����^9����ܝ<P4+G���<����5�]Qm�Q�tdN�ÁR.�#��I>jҀΪ��z�1^����s�O$'r�.(�H�<����_���L1����6��'>7���>����p|F���w������N��Ӧ�����*r��x
l�Ur�e��,8xg�z���'Z�A��k��(�Dkè:��O<:}�>0��ꋦg7�}�����쑶Ux�Ѣq�Hv���.�U�0}���_u��^q=NjݯU,��"���-���>�hKs9�o�Z1q�C�ı�~�sJC����W�R��`p?�Z��LW.|	b?u��r����4W/(<#<<�}�T�zT�k�?9
�z��v�Y���T��Gf&,�)ڄ&���<���G�\nL�yk�}�=�Վ�sUb�Q��!YMMt5���<���=Z�V�Дw�f�<�y��V��b|�hcTF_Q�m)�<=�N��{ݾ����c������j����Q*F�r�&��-�e����e�'��j�Hg_ث�UN_!cYvxv�	�b�VS�$�K�r �	�F*�B���r�`D�ѳ$W;��
�\��x$a~�V���nmA���	sj��.�X�Z�c�x`�$Q�+�8M��Z�k��˨uI�����X��A��6�KyIj�Vf9��T&'a�Q�5�N�Bt!T�BnŅ4e�u�D��,��1�_l������a�QX��&8f������#�%�
�J���u�]zB�f��C}��A���y�/�V�>�����k�ƣc�X�v���_�a��,uz�Яl�:�g�6ֺ�T�����H�ƾ[�'���Ea4��;��Z�Չ�`�t9�q}+3���Z�j����>��E/!t��l�﷭n�g���p�0vv�c�����}m+�}|����.�fa],^=syKmƿ}Y}UM�:E¬9YW�J���l�Y)�O~��hVA�m��wF�6xzݞS]��TL��#�7���06;��=��X٧7�\�R4Xd����ū�r�<z�g�It �#:����}�D��=:1�P���XTӠ�=Ǯ�o�/*��}��u�_X�U*$Y�G�0|��C6���f���F��p����'93i��q=e��;�	�ze_s�6�+��@���4�FfS�������xG�����Z'k{�P����@��=jZ�	J�:+h��BEGC��2:�[�|��П��hM��d��&��@L�s��D
5�\4U�TQ"�ܰ[�u��SA���N�4�����Or���ǜ��xeJb�(�|0�/`0�I���"�_R��wk�,�/w�(��>�棶��"j6������Mjmj�sw�	�ls���T������Jo���e�ҥG�� 8찳rԸs$��a�.,��{�l�� D�E&rM�?�;NMyvV,�ˬO�	�PZ�}o^�˻x��=,{HrOjb�O�n�g�-�e������_I�q��9͂��g�禅4ӓ[����ƍ��z�)�o|�����>�SY������x��r [��YH�|[G_�o6����^�6K�OoDH�.�z�5���:�?s��kF�������w�*�<�9��%������檒X���k���m�hҰRp}�/��PɑK�6�;D`�Z��?r]oq-�I4ذeb�ޞ�gq�ۭ2we_oD�ʴ������B�4�3M�W: ʁa��nLJ�:+7�uC%�Y��P��M�7��i�
��F�A8��V
��P���é��zRͬ���U���%3�B�q�v�;"=�s�n������ܩ��G�燀7�i>�~�,�����R���6lZ=@�2��v�_�n���ċG)��|!a�ԳB���>+#�wեg*d�/�
�=W4�xemމ}��:�"pc�9N��2�_T5�9q���U���Pt�ry*+�����[�nѯ7bH��ʰs�ġ_f�mwK)s촞j��^�q����� �J/Vkl����,u�D�O����]3"woR��6딙SA��⬈еc�>���N�v�=#�����%<�V}�[�JJ�:�칫�Ubv��-�o-d���=�Ͷ[�a%��ׄ���R�{�QʕL)6�7]D���:�ӭ��/S�І�5g�8D7:���rhb����B���$��72��-iS�'h�{����U9��gohޜ
�e��gD����� �Hr֖�S����ʆu-F�%E}�]��u�����\��cђ�{�Q�*|;"]��l�6�,܏�fK��	B�I&�z� 5�6���`5�7nswGy��
�a.�M��[���%��L���}�7���:l���E.�|���G�X�Ԩ��樐��&Z�/j����ww�����}H��՛W}Sv谰��w%m#���f���]s�I9'�e���N�oT��7�v���pF��M�T�rpݴ�c�����,R_B����!�aH�}w\�R}5>,�YՋg9	���ϕ��i
���z+���Ï.��R�����=\����sE�a39��GZ�����Qb�Dq��Q�}f��{	��7�2�ea�X�����*�s!*�7I/S6��se�k˵e�(�6��� �ռs�9dڣo�É��`e�1�u���_�0)&/��Ţ�z��Y���4��p"�"�x�ڀ���C#s�j۵��)TR�C�����zIc�#���(��4��n}إÃK ��I�8k���]�X��Z�2Tvy���`Xs�^O��k��3@h�g
���x[���ZUs� ��&1(�p���ԓ�V�nT���He��P�+,��q�g]3��*qAs�Ѥa�+b��˟&�@����ڡo��\���ǭP��*�N��i�����M����$��3{niBm�v�P�謡�j`�3�l��Ů�i�p�ﲦ��]Zcv-�/����gn�|��fF�hh�G ��I*�7�I3�bWj1c(3���iWf�@Q��*_[�S�WV�����ջ�y���M�D�:7\<']7yҁkP���g{��լ���f�@�	�p¡��D@�hv[�X��Sv5Ir���f]�2���*��_au�IT��^��IHd[�����	�0b�d�xp�)�G;�^�Ƈ)����K�W����ٗ��2�Ye
Um⭷P�l��oʶ�Յ&�]Cr_7v5t6vC"�J��p,��Ք0*�1mol�������P2��uJsRrִY�Q��3U3Vq�.eAj%�Q��a� eJ���]�/���R�0���[r�U/,mG
֨�-cLҸ�kNb�]jQ�J���┪���-Q�UN[���KFŔm�s#j2�g��K˵(��VҫkNbŉZ�EW6Ӛ���9j)�%��Z\����h�Q��Llh׌��ư�F��l�L�QQ^]�m�Z#��*᪈k(��G�]v�֏kZ�kDsQ
�b�m����^Z����h�5���p�[�DQ��9�:֏5k`�Pe�GZ(�ƩY�Pv�r��Z��r�U[l�j��^�{����y��|L��� ��c۩���tj�қE��P�܊���v��%%����]'br�zk�EK{�%�*MQ_������vS��E_�{<����Ӂ�	�9]b{SV��;�����-���-�ǺֽR:��:�fh|���������ʞ+L�
U6M�	YH=�b	�.%D�E��y�\�6+�Zv�U��N�+;��]���C�����&?
�s���B ǌ���t{�Eb�ޔ����Y<X%
�h9F���"ѡF�+�v.�h�[�m���#�-����.����7��!�5G��eiT���L<��<�]�߂갼�Y�����%�L��d03��CHn��-�V��@�~�ًK*(�y�f흆�+<�	R�	�
J�P��97V�r0x�Lٮ@�g":�ΈW�K�r7�{���U��XR���+Ph����э��Nf��z��t��'�u���veQ1{��{R����#y��/P��f�ٵz3/�'�J�8ڝ��b�m��=U��C����q��}��^��uVk���sk��t���pISڎ}�HW�Z��B�f�U��|�k�S����=�R�W���))p���^zO���O��һpj�gw��.�xø��1��2�%�oM#A9=״�a|��Q�@{�'�?.����Դl)�Ȳk�M��֫^�A܌}:yы���\��	���/ʲ��Èz<�k�ƨ�WW�f��Od�|�͵A���'M�e2��ͬ�]	��[��%ݻ�[4�<j�^�h(�NЁ]Ҫn�B7����⦌�ܕj�.��nd�$浵���,9}�V�s�M�z;�R�U����[��0.Be���m�x���(�������q)+$��Ee_u���úJs�ᛩ{HӐ��a*H�h߂�#��S�A�[�����w��'f�4!�A5M���L�����(������5�*�a��K!��h�k�+g/�aZ�3���p�;B�Vn�)�-��:�$A[v�Q�}n->(���aO;:���Me���1:�Bb9᢬��͖��ٮ��J�C1c��C�Z{Sm zx��8^��x�~��U�ʵ�ֱi[�r���#�6k<���.�.G��u��z�tVW-�j�J�Z��OH�=7�tG����-�<�!+�M�'zzOM���{��Ѝ5��&�T띪����<�s:l�[Rǻ�R�yܟ7��.�{|^�f/|�ϸ];�Q�y�y�8C���7�m����)��HA��)�6���p�i�ʜ�\�J�HcMvA�uc�@�od?�U}Z��'��Ի�>ȡ��N`�.�</���v�S�W]7�Iw��Ͼ�2Ϳ|��mYJ��+&/�ӣ�^��r�S��稟H^�"�tPD�b̪�G]Ew����S�ar���Vt��9mQ�x�e ����魲T�FL�U͢�6=�M���_���?QЛ�յ~*��ɬ��c
�Z$o�dj��m�6����J��^.q���}ƓJ�G=Z&�mk��%�_��Q��ev�O�.�&	Q�ы����>]�f7���%���J��9#b8�N�8r��^f����1vv�-aLz��&��9`.�<E��ˍ����f��6��z�H}WIi�\�9�YwY��f������HE���e��+y�B�N:�y�)����f>Μ���Q" okoO\h������x�q-<�;独f�c�Lrhۯr�*Q���̧�[�^a{1�v*n��4������ ̆���x��"ؙ^�s�p�ޞn�.W&m���pS���L*;q�W�;�i:z��wo�)�q6(N�,a�o��,�7Y��Ů�c�R����I�g�bv�'RE{Vm�������~�h�Q"��ֽR��X ��ُ������-�(��HT�{%N�ўV��^p������9�3���|-3�m�gt��Җɬ��aɬ����8�v���.�WK�)uv�4*�p���I�H��z��A��:�#��L����:D:�D;���K�I����&M�bb^��¹|i,6[�7����rF԰b0�D�̥�Qy��cޤ6��o�:����!�NB,[{7;ܒπ s��-M�v+�#u)�����#�aw׆�r�{���Y4�V[���=�a�u�]���ʰ������E �#g�
!�2[[TN��TO`�otI[�;�&���%��浱EIp�Τ���%�u��1��V]Z����k"k�J`_s)9��{1����ϸ}���d]e�gl�fh��q��<�S{�[$��|���C}<{�:�i%�����i4���m��x-�[Zt���e)�/����t1���j5�^�j�`��v�u���"v��S��Q<�qK#Om,8����8B���ngM����I굺�5w��_(x�'���jE٭��Qwz��敋�,���
L/Dy��z,��,��sPȟ�N5�%�hI��m\%3*��� ���ڽ޼���+�K����\�֧-h��Z+NsK�yoia��ׄ>#+�i�\}W��TE���ur����1���m4��j(f��BeP���hD*v����~L��i��lU�NQ�2v�W.sv�w(��������թ�֮��l�RF`��|Ţ�t��<����\�$n�L��&��I��p-E&K]�b."�Yx�����w�U��׽��̥�1XZtN�ێ5�=Aˡ���굓c-��>u��+lv��g!P��>a:��#QugN��Ξ��$1�i�m�"��]C�˧^�L96���:����&r�pv���_�n=��[=cHǵrg"jh<ⷍ"zlǛ+Wt�XZP�o��"�=Ic0w-f�r�(zEpi��wI��Ƌ�e���2���F&mRۅ�%v"t��s�ꩉcQ�wM���ܬ2g�K�{j���qr�P�*�c�n󣾧j�o=���Q�3���Ѝ�d��ẻ??s���}\N�zVa�}痽����W)�����谑��Vf�^�M~"O�BW��Ż£�I>Ӫ�X�Z����/=}i ����:Rt���!��Qcˋ�mX)S�+&/�ǶeDb�8���V��ʞ-�]!S"�9�N�^�5�%�C��Ӵ��z���sG9�Gz�x���^mJ9��S"Gp��i-����VY�X�jZ�˭#���X{^��n��_Jz�J�V��k.	V��h\s�kTخ�쫢��в���r���0�C(C�s�1�7�+j�xU�r�����ݭn�w���V���-�3u6���r����r��5��b���p.W�8��g���F��ӆ��0U�X92�����w���5��'�m���U�*2m�n��L·s4��%���d4��"Q���v���|�^��+;,f�!^"=�'�6q������\��=�C劷��)�����'5�C�����d�X��A�
7�1�����{�"�V�+��m��)�ܖ;�ם���E�"����/�՘��+I1�i�Eu]��F�l��78NN�=��\��Im=.�� ��H'��5�[Sږ_6�2aWDЯ	օ�]�)���i�h�0������ ��*�惿y�d��������y�|CG˟��Nkh5U$�7Ś�Υ"^W�m���I
�yiN�l�]�����(L��+s9[;Sw�<b����m�5�H߯ԛcv�|$Ӡҕ-v�]ERn@ͨÕ�
s�8�{�����!������Э0}�1�qu������[g�I��~�>י<>���i�ެ�OQ��F��w����Q�B�}e�֪����a��>�X��d���دZ4���F�ϭɡ�#��ZQl�"�+,>��C`�SI���л�D@���]
~�SӃ��U��pB�#KTT��I��sA4ڼ���;./}(�3%�b
�����2���/�kydc��sWv7f%W�y^�� �cnMw�q�o&�I~�J�g�y���r5=_���=�}Z��^�\��/Do����+��&YL���j�O�/
���W�&����6Zә��Œ�kuZ%�c8�Һ���,��u�&�����^�M-d{�Vk+z��g��~���&�kZq�G�w��:�GF&wjm�M����{��5���1�G��f�-�zze��0<zt�%qX�k-}�K�)�s3LU��3B��bGɯ��ɺW��R��Sn��j�^�§�RÞN��|h�m�'d!�iW�LTOQ�޻Q�37b�d�ەdvS�/:-��AHа�]`:�s =��b���*jpu�A��;���n`�4kzZ�B��C"���2!2]�������tV5����M�LڝE!x:>u�-��b�%df�Ǽ]�ov[�W��F�� :�1a�L���@'bi(�w}����4��ܹ�1|�'l𽹄&�m���������N��l{��`&�D����u�Go:���zr��tj��F��P��{)�����+#ò�h9[�Li�p�!9�eD��Ҿk���+D�yJ޽×�a�o1�MF�cz^֖9vn�`B��!�F�Pvz�㌨�ƕ��M˘�P��X��w�z_h��v�c*hV� ��j��Vu��
�b�����z�����T�n��X��.$onZ�������/��6�m�r���r	R�C�m���	q�j��6�p��/:�T��a�d�SUEp� ���j+��ޡԞlȻ���E8g9�8���lIFR�xs>OK�Z��5dv�-���a}�NB�&N���#�k���T��^���*�����F��!@�0�z{�zb���X��LҸ�o�̐�&ݒo-��[�dy�3,QS��(����iqϦɎHz�/E�/��:� {si�{j7��������՗��h�564���*��>�b`�J�+N�_X���]�V���Plr� Y�z�V2�?��,�Y7[}z%�v�q�XF��G/h��x�����1P��2IXCg&%#�̂�R���ϧ���J�V5(�>k����ADcǘ��NR�:��:"�0˫���ȹ�b��)��,Ff̕G^b��cyIDUDu�4V&�E�-(���H�5(����UNP���s)D�T@V+"�R����m�-��i�TX�V�.j��6�DUa��nv���T֨93Ssc-F�Ĩ�*�ImMJ�����lfJ�5�Y�R�-Eb��
(����-�ڛZ�L��+bcm�����h]]W%T�R&����[.,�9h����U��neכ36ч�)��4eb��T�D�Zi�QR��ʊJm3��l���+l���m�������-�Nkκr����u�ǬJ���L=%U�Z�幭��*䠋PmP�lV�i[��m��X��ֽ8V/M�/-��V�T�g�x�U�����e���������ӻL�$�ιN���-Ǘi��_8��'b�Sl͝j�mE�5�&��d��t���;s�:�ܵfQY��IPs�~}v�J���uw��-�P
���E$5>�g�8YY�V��Ċ��i����U��7�y�������d��U��o�����h=��&���!�+�;�zc�G��I+��4��yА��.�͓����ƨUV��s�I�令�̛	��M|*2�w �nю�k;B�i&�1�O7F"�m�i�~2r4܈SmpWՑדع�Gxo4�s-���h;&��3oq�`��#ef��qb��9s^�\�ԵL���1��i��I��E�`����4̽Hlw-���۞��
@�T����iP�z���Ч!�+0V@���ӳ�L]L׮���<q&�j�gp����N�y9ys�D���z�^��c��UՒ\�킱o��I$��߽�je�	�6&�{�M�HI>�E2٥9Z���&��s�ڼqW�*|�oe,��Ikĸ.���1V3i��Ƈ�a$c����5Vt�ܜ� �[l�k*���0q�|LK�^KiLq�����y����-��/S��6JT��i[��}a�M�ul�,=��A�K[�8��Э��K �O4ǌ)�Np��ٴ9^��M�Y�Ú��W�=�^m��i.d��1���F����[ӊ��}F+{�"Ƽ�oSf��談���ߞ-���yj�R���N`�Iu}\ww���PZvK]���5�C\�ٶQH�(�䊌��f�۾��9%��gP\ՙ�]�a^����r5j8t�1P�64��U�#�;u�5�wr�ώJ\���
H��]:P����8�C�ݽ�\�E�<���-M?{А�.��V��ų�qsS)�(eE��;�������Ĭ�3������r�J�ޠ�;HH�{9��+9�����7�iѥ^Z�N���j�`�ނm�_d�=�;&�����)P96�l�A+�'N�kv^V����
"�S�.J�e���W��zc_m_r�D��О�{��\yq� w����x7��Ǜ�nUqަ(�����^��H��X⺸�w�zj���](N6"��Pg�d�p_8
or�_2�\G<�˙�/F���[93O'���Yy�X�u��ٛ�j�S�_�-߳Q���y�'Q��n�;Y��vu��Zs�6�vi���zC�{�un9�(%��
�����j�ڎa��(�����kz!]���l��2����wv�����)�q^�^-G��Ͼ��s�RL�}�ܦ�w�.'7���TD^c��H;��Mu��k�S�o���[wϏ)��:��nu�s��X��S+;t�7�Իp.�v�=:p#a�t;j�M��"9���&V���yi��#���Mk�����ǆ���iΛ��=��V�:tY0'�e�"K~����k���3�gCs�Y�=i��J0�b����k��8:>rV׃�.�z�4�ʘ5c]�������v6*�CG@sޓ~��wd䫪Q; �.jgf�F����B�SI"F�-��# Kg*�ᲷT�b%;�S��ˏ.9�>DQ\��u��[eٴXmx�b{U�����Q�F��5N�1�u�Ӥ�A֔(m�z(�O��jnJl �[��[�jm�.�4&�l�A�S�r����keO�<q�zS��OL]w`��ّ�=Hَ-�`���5��J��I��q7N]���p�5�憶
��c��v:�>*{x�1�ht��LZpJ��V>>�4]v���o�ީ�.���&���;7u�^ɭtZ�u�쵝�<%���^�f���	T�>�+k؁c���B�̶�R���Ƴ{GuP�o<�ݝ�d��g�Tv$���؛bZ"�;��!�16{Ng�d����o,�����`S��B;�d��i��P�=�Kӟ�}�q�]Xx:�ɮ�/��L�ZB<Ӯ�K{�YJ�o_�MJ8��*��@����suz�L��sS'�X�D	Dj����3�h>�M�l��N��R6��M�}�n��5VeYku�;c���<ɥSouoE��+��F],^���o�O
�w:>2	:r"�����=�'qSL3���=�ⶇf�$��i�������:`��mWk�T�#��7<޽7M#�O�lW�����Yڒ���f���~}0���4�N�Ū�5lI@��{���&�g�U�ܯ�ez�}I�vvi�2C�JQQvy�rxf�\℺�óg�e�JM��ܳ����ɍvJ+�j~�e0��^r�8����L�x�<&�v�3�"�#*W�8��6��彝1>�B��!��gV��5Ƌ���G)m��}!�-8"y�R�ɐ���g=C�.#��zz�~Y�n,c)���:gI3�2ڞߕ_p��&��m����Cv��z����z{�o�%U�'U��,�{hV���7�:�.���8ۚٻ�K1]��7�gהݻ�\���^@� ���8p'���N�r���F���{��M���^���sY������3t[���NHȒ��Yh��z��;mm�]tf��M��{�٠�<�$����?�:g�����<��r���N`�%�lS�0�Xܘd�Ee����/�,}q��8�x:��<�5K룼�v��F��P��RZ��-���~��nb���=��qd����e����.��^;���+=WQ�̽�W���h�����t��o6�h]4n�m��eWm'�N��!Ea��=�U�"ѯF��A�|�3N��i<j��ڱR'��J��E1@�<���Wr�qK�zdЄj�;JLW�����U�!'`/�������g �1�hU�yW�r뚖5��f����z&L߶���K)e���Bᳬka܆fZ�y�h��a\s&�\^�8Ԩ#;M��[8^fR�t8�
&cz�
o�79rGo�3��`R�~�_W�*�Y-<�V�
-��'�$Q�9#�ƽ�u�}Y�g�{��]�*�,f:��'[�q>J#c�;�9[�Z���n�Ű�3�`N�Y���Y����XU�F5���y;+c��0���w�����y�#&׭���p.? R[�&|�kt���L�Ki95,�q�^y�n�w�y謁�a)2���{|Q�r|6�{��"�qa5o�{�V{�Wq��A�ӈ�u�:z�~������kT?syi���lr�<�꺺U����������4GD����DH�M�)��~\9O=S�.�c�M�y�b�7��x�_w�?
o����%��--�c�����i�^�:�
l�I=��2�v�oέ0�]�a{�g>�{�[�Gn��u	ٵ�%�t���}_/n������S����D8瓦�َ�W,��Ɍ[��;ɦn��]O���G@}J_o�I�U�^o>/{�������Cc�T�����ks��˹�kuv.=p%���'���N��4!�	��8i��m* ���-`�s#{(pi�'��1�2;iRl��m�J�v����Sv����W�R�g~x�L´��[/�_��+�5D�pEZʜ��E��`s��+��K*]:�)L�8����gf�VYw[��nmC�o[vi���[y�RnSɟ8B�&}�W]�W;����܂W����G�
��=���[����^��Yx)-�����+{5RS��{���E��ƌ����YX�9��o!&���_z"(�	Uד�3��ɥ��S��*,@�nej��kc��V"i ���9=�R�Vu�V���I��/G�oU���E��>�,1�1=���#�+!2zrVY�a��˯��;{iZ����u#���%0�	tx�.t9���.��l��5r����>��������&��C�GFWN�Y8`=�s�7��{u�*k{7F"�m�i�`�N�=}z"�k�!8��6�i�����M��bɍj�)pg/J<�����"���H��7�_Z�j�1yp��U���H�&��r-T����};=h��LlIq�'�(��!p����\�b^�U�6ri��\dem�Y:���K�d2����4�̻FXǪ�O�؞�V�T�]wQlޅ�˕��Y�̽�uF��Źj�!�ʓ;��
]�Tur\�ee���e�=:cT��܌3�f�#�/Vѫ�V�U����E��9-d��8z�v��Gz�Pv�!�
4I���gs��y��Iƺ�C�,�Ss���]1f��W���E��oH��i�4^t����*#k�VSMIX���i�Un��S��2;��c�*he���O4Z�e!��6	�ƾ7�X��>�2b�l�N���0-�94W3V��V[yا��ŭ�N�/1����غǨ���������2�1�5�ޗ��<Ɍ9X �X�[ˇN�Wǟc��X,]��łԆ=�2��5Ӄf�S�9���=oiӄ��X�����D��ڮ8 ���D ���l�5*�¼2���k�%pD�k]j�C{@d�6�5����i�V���9�<�h9�Pm�Zl^t�OA~2�����/N��� B^d
��Q���$����U|�?	Gx�fW|�";jm,%R؂3ۖ"7�%�ڠ㢕<n�Y��a&��O�Z�u!�}x�J[���
�R�j�<|���G8��^p�Nq��zuĖ��C],;�΂=�>��!0]O�^��^v\m�;��ؖ/z����� Hn���ж�c��bڂ��N�^HΚ�j"�a����.�wD�;3L�����'�D�̶ /E��4�&D�����&Z�/�v��*ڛ8bV�]NyPI�8�� �VR���V-�$�>�k�kaT.������O��kb�5�4g�j/;D���D�G�ڎ�:���Ej=�(L�9�=��I�vQ�]���V�S
��[�h�@���w2k+mή���]�6�� ��F�k�v������u�)^�7i��λ80�-y���y(�ɀ��ۜk,���z���b�5R�k�/�v������GW���ɺ��}:^4�7���9AÄ܊�[�4��3�ʙ�\&ʕ��Ќ�5�"�
/�����~�F���� ��4�_B��WeV"Nv�
���=���OGT�H]R4v�m�}/8U#�T�\�#���k�V�e���oQ�h�~�_V5��QDo)t�(檨d��q*kb�<�fVjE-��C���hTQWZ:ʈ���r<i�Z�Z�,DͶ��F�m�ʃ�[�l�����`�DQZ��Ѵ���l�'9�o.-���5���gj���kJ��FJr�Z�+��7r�TzJǔ���b��M�(���F���&���67Z��^Z��E�X�8ԩDFjs�u�W�[o6uJ	�U`��֕VFЧV�)�����겶ݱ�QgL2��"�c9M�6Ӎؙj��ܦA�h��b�ڪ#�t��4DR�x�u���Qs�ʪ2�*��Ml���`���䭴��D��X�r����[��6�ԗ%Zδ���Ӧ�!��C*j��9Æ�(��,(�Xj�L��i�b�9�UrQF5��������]V�jez�����y��̣)�x���/uh����X�n��sY8��IMoX�w$Y|{o;4'���7L��m���K;~6��
G�`ڪ�Z�:�uc��16���s�����%+�2�7~u\%��f�No���Yl������ۮY@�-�h�bͻ�����y��ϲ�uk��4��<T���
��F��#�q�#�v����93g�Է�� ��0���u���6�R/{p��Q
l؉��u�gR�Y�V��OL�I�9_�����ϩ yjrc��U;b�ȡ�3��W�:ߢy�ز=E�H�68�98��s��ա��6w�$��'=�/��>̋�GH����j�`���ie^M�������4WT����:M��|} u?!��l��}h����$�J��N�
.��h�0�
�w����u��7׃�{n��dSzĈ+|�)�[ۓ�f4�ױ1\,��o���[7.�ێ��&���x��)���ﺈ����zh�4�JU�>���V��5j�i�V���w���(۞w�1^R2�L�P�%���q���BY�l�m]H��Uȥ���W��B/�����IgdSdK�d�#BJz`���NP�/r�����V1A)'�s�+%c��I#q�˨�!��"q6���7V1W�y���$�[T�,���*��$��3rK��#�g�fe]�!����'���#��Sj�1F�ʚ�ג��&����������bW�|E�fM̤�EoU����9�ɔ,�zM��+�]�E+�`l��5���b��[7���A�,
V/cY�G�3�r�y�5S�W4��t�T�e]L��I�����2�ޭQ����;�(��e
���w�	V2�S\���*�w@fdea��{C.��=�=�4�lVk��ܡ��jbH���W��n���1�$h$�����h�
�N"�ء�a�p�����po��t7H��E�+Ϛ[^�\��cRMIq�1�M�i�o>�@&ޮ���%wJ~��t�	T
d5�Y�kמ�[��u��Cγ��~��q��ƙ;h4�1�'Lm���p*�K�.(�5���Q~�#^<�z��;i��+\�c��6��KWt��@]�jV��z����"�+(�Un�����0���>.i�b��N�d� ��~���sT]��1��>��k��p�72,bO�)
7�j��v�N��Z'|Z��XY�)c1�a�[�y�Vc�F�g�e2uzhAfX�z�*�{��s�{n�b���J:�ۦ��C�����qo��i��.3VKMr��]*aböK�04��q�y&��!�t$��%���nשW���yIV"v��5˖����.�告b<f�����e�hz�K"v��c�,�9)����i&�uKN��t�7���ʞY:N�צOZ��	$�b�ݺ��;u�Df�b�lj5�j�YH���T�,�h���`礙���7����L��R+n�����z���"Z��Q�Gq�i�㞚�S����`�w0r�m�H����d%��kQ�\�
x���:�x��e�\Wq���.$rzw�4���/�ʼ9�(\w�9'Z��>�/�=<�ķ�+TlY�P�����qܛ���ez&6��Ts�ZG{^'��iS�t��R.���h}�6a��
�Ղ�8�WY^��{*Y2��
_j�����<��++=C��[v�lRƔ��v�i޸�#3�2�Ⱥq�/����� ������M?��d6Ͻog�/勑�&��z�A]������/�xP��pqW�����vw�s+d�����G�#�lM��3�*m��M*�,���\�TzK�z`�k�^IOŇQ�\y����Sp�r՝��0{d�[ԅx��9"8��r{��4��ի��g4U��חB�k�˥	�0�PL_�q�r>�Щ�iV��vv�,��t,���f�{�q����\�7fo��a�eb�o�ǟpG��[NCk/U�������ܬ����sT�抢(^O����j#�L]ݾ�,�M�P���m�5W�J���G_�A���K�Sѓ�}�d̕�G��r@W��Z�yr�L��r
z�T��#�N։1�!ڵQ�ig�u�^���pX�KSx���L����e]��ʮ��Ѹp~z�L��1:�x2��::��.u��Y��%቙���=�C<�%z�u�]i2��놠镪ety�c��5�.j��q�:Z��+���pİxסZgN�t�I]]~����-�i�@�{/w�<k"�q�3m�Wa%��(2E=^�Ή�F��Z�Q��;4��^4y�ݸ뙺]O��Z.�=�(�q�tNC��}6�3�2�#���Y����Ԧ�S�H�˭��Orv:�p7k�%3/L��F�]��i�E���ֹ�'a�L�wV�c�
!O�g�2eM�bn�5g��\��+}�l�wvk����S��S�h쮖9�+�-@j�����氊Z"�*�f�n�(js;��U���ҝ��I{��>�f�٨.��ɾ����2hq��{z��?*̻{Q�{;f�vU{1�B�.��s�zl�K�_S���F��Ҙ�tE���"�U����p�����G���UI3���bצae����L�H���&q��>���y㽶�Z�k�=�-�w5�{\�W�Z#�S숡1bl������F�s��[���Uy.8�<���kc�epõ�Wp����+��=����\�1]�\a�L���굗n�p��ʍj�<n��U�z�N�!]Ɵ	�������P{�����~M����6��U���:'rfy�r��I\SY��ӧ2ڣ�A�W��T�W�i��ק[~��fc��%ѩ˯^����s�5�Q�Cw���R��H�x�L呻[��k#�r�����$���ܢvr���F9�\���,�ZA����,EFT۲���;�[�VP5�lFq֯������S���nƔ�̂�U���X8]$tC��i�z��gb�Tx۞:�8C�)�C��$may�9����9u:�>|K���W�	S��(v�����b��z�Ŝ�\aa-���/ǘ�#ܢL�L'�U��)w$�w_y���Jm�������;]\bI�tV(CKP�]-']���=��.7^�'yW\�u��>�Ԟ���{���I���^� ���qyݙ�Ѳ^���
去{�ޅ�1�o�p�p�c�F�ȶ~�o+P�K���M�wm���>]f+�&��ߝ罕�ɱon�g��ԯ#P��h`M%j}q�����+���ujǣm�<�v^�(���^e�ܢh�] ���Wj�d֐��K��ep��m	���֟ �ۗL�}{5i7��&�r�|�G�䧺�{��xO��62�QqC2�B��H���f�[ޡ�Pgz�ME!�q�NjW,�Jؤk&i��Ж���K{�A����.�����呹�߂�:����2Ҡw�<nv�t��O-���Q�z�ի�Q�Bo���W{��=� �J{Yk��D;dO�� ��ˤZ��|��^�S}{�j�4�l��a�N��^MPm���H�����E��	��~�͘��A��Oc��Y�ݢh��w#fE�*���=��� � �
G��U� ��(>�'���&{��)#����V����zs���K��mGoӴl\M��'a�C�Q��'��߶ވ/��^|��X5�/@��kH�/��;��`~iҽ2°�|G��wY9u2�p�k�lȑ�Fs\���|���y�u��.;�T��ֶ�H�e��s����+7n��kc�4��G���9F3q�g��%��k)L`;7^#�}z(�$���xߘ�!��7���M�T�B��ÏT�����l�⊛D-z���KV���|iM�6�La�[|���!�}��������mvWܵc6�"���bw�&M�efh���'������V�!�iF���j��-֭i�j����^��h�^�i�,�S�;%�nNr~7������{(�7"�s��N\�6��x�1����C���~��F���g�)y�=����˭j_jƱ�K�q������rS����ҦsJ��n��D���t��/q$���R�q�-u �77��-;��L�!���U��F�Ž؎�L��t��V*���e�ڏ�f��^��C�i�j�����-�ޱ �b�A�$�.dF��x���f�z����W��oBH�:uLU�"L	/����۝�[egY�D��P�QN����l=pg�R:��*��Sr�g4����:_YV[�D��_Oq&"��)e�i��+��
����ڮ� ^�
4Z��y�Y}�equ���Į�o{)on�_j+��CC�m3D�kH���\r�a�ɇ��{���nc���r3�#�3������@U��Z�n�t�9x�	�r��o@���f7t�.ꃶ����uvo'-��&�JݾT�'������G���.��Qd\��B���n����f��燧K�o����帀�ը��e��J,��Fa��ɺz�1�ܧ ��;�2�gU�j�3)mv�u3)�t�{6��{;�v�������{r�!��6y�p�7.g�\�3p�͇��G{M�׍��)��.�W9Y�y1p�6^J���E���M�r�w��j�^A}�j���8@�R��a�(���1�c,�ٸ�����ή����0�����kR��څ�2j|���"�wv;����+{"08�6��Ɋ`��]�}J���ˊVS�x!�۴�:jː�y�yt:&�yr���e�QG2l�9,���]����+Aξm���h_H@��=O�Ճ|�gVK��)}�Wz��Gx�j�TYB�f>��l�K�g��+<�LV�u��p/+hN��Z{%�D!��@�yYz�q}�ӗj�N`:;L��[�s���X0�-!z��' ���0�门�Oz���P��9%��}�qR��M��vl�k�e���n��(��:���k��e��Y����d2��S�b*������u��v���G�0 �]����q�{�(�Mp���8H�Lel ��Y����.kjj����e<�"H	��1,n�Tx0���J�6-3�����k ��x�[�Cj(h�)P�>%D]l9��v�\�ʚ+5(�U]�Ռ����Nc��F�򖔳�9C�"f�̊]r,��Rڋ�1���8�Ff\Y�pԜm�u��re3Ī�V"���q,J�ˌ�5����:��1
�:�D@y��y�7nh��[�\��W�m���Fػsq��j��P�[y�����mV�U�Lr���+�ɥJ�rל��������nR�#J�QE�faQrG3s���\ڬiMK�]y�a]J��ٵv�5���m�%e�b9���kU8��y˃�.��1^:.Z�"*��
[������sP�V7p���^%��i��Uyl����9J6��ֺՊ�(�\�������VaQyh��ʢ7�]i��#��Ԧj�-(Ѹi������fAK[bR���vE�حd����ZYhX-J��l��m8� ����ڈfc�ho�&�����R�
3���T/��} �s.��&\zN�ǎ�=g����.�jnq��&�����iMjS1#f�#I�e�D�R*t\�S-;��Rvi�9�r��G,%[���v��Q0	%��V��>�B�)�NJ�)%�yR5��9&؎�������7������rvf�O�}��ĆU9,n)�H�ܬY�Y�$��u3��v	��:��L�tR����>�-i�^	ڮ�-Y��eei&�+2���.w�MBL�s�^�����[�<I�K�ڕz.��2�͊�ā/��}7�x&QcS]B#�&�Nڸ�c�ݾ����	�<���kc��P!T�|õ�	�>\��'~�u�*l��7h���͟q�XP�u�d�yHиC�fͯz\��Loa�y���r~�����:���OA�Ƚ}=��]���K),���#fG��ƈe8��/r����9�?Ohj��|���b�GQ{��-X�}c[׽ɧaR8�]�}:zGr�;��);'�X�J�}Gz��s�i��&�t͵]΋��wx�|b5�6�a�-*;�5~�ŒT���y�%����$/ ��ף�!W�����"���V�S7�o�}i�[0s�(²�7�4�����I�6q9�M�x�`�yW� ��94/qژ���z�(o�ǋ��ʮ�`��Xm���j}��՜�j�Q*i5�ǚ��`Қ(�"=�$�c���&��˜���\m�^{.Τ��~��I�6������wG����@��֫�D��y���0RQ�����w2�x^���@�3Φ{�V�.�� �b��F��A�8ࣖ����S��l�ƹ7,<&r�<�N��(��)�������}[��B\n@�n2�1��+Ѽ����2{��f��mR��x���Xuӷ[o5����Ʃ��ց拲y{Ѯ��#w�X��C(j"�d[�&�f�t�B�4���m��<Q��z,,j���}�W��nNy�^�O����5�0*{Ci�����;Kn��B�K�@�y$����i�m�+�J�P�b7.�n��u�{�4w�=d�w�b��!@���;~&^!�ܓл 9S��=S�6xË���7Ao�k�o����$h>�7��{O%���M�=�����ax�î��A[B�b��(�ͦ��#��`g��%��Ֆ���U,Y�R��/+c��� ����܊<D
�CbZ�A����zY�gx�ٯg>��I�@��������K���kk�-t�Q� u�`��S=�d�Y���a�|��@;��W�)^������9f��A4�\*C:��u�]�d�	���Y���t����[#���r��yU������J.����{i�2/�_I�sw�o�/.������Q�@�/^��W�#q�P�go=;���ױ�lW'ݍە!o*Q�ͳͮȷ�\�f�f�ج�bsQ��Gb����im��je�"u(Vm7��e��t묹ʬWؗ�W,n���=<��m�����Kˋ�����$���{�Ug�E=�ԇ�J�|�[d}�VfP������S/mdf�Д���6�^U�^Ͻ�"�
a*�<Ϥ�h�l���T6��,Y�[x2���q4`��s���M��_�.g���(�˺��x��}3J�b�l�PZ����dmI5%�o����Y�w�5ݞ�T��r�x(�l�e3��&�I�uy�������p��q���TY)
����[t����e!O��s�F���c�۱�){3})���*�uycW����A�.:j�EU��E�K�V4d[1Ciֵv\2)#ņ��c)q�p}�૦�5�%>�yq�J�l�m����-�>G��z�.Ϭb���'�d��Q��VGC%;��)����/ tM>��[�+��+s��Ҹ�4n�)�]��R�Kn��q���f�Ov�n�,�pgT���==�m�C� ��1���9�Ak-��q�3�S��^ɏ�w*�* 4У���� n���Py"U��/%��mV7�§3W���:�����vKȄ��=\�lɦc�#�����!�Tr���mY��:.�%�o[�bKTe�׫���h���fej��\�a��k��4�ЕI[����w��cp�W�����k�RX��<�����k�j^~�����o���T�Q���cj:�����'վ(�}�د)��կv����&�M�� �{��y?
M�q��Z_*q���V�C���p�f�i�6®���>��4ԡ�e���6�xx�z�k;�o�m>;ۍ3��htt ���e��p�~�;(�<+�g��'x�SƯ�%m�o6sQ�G��{/���"�h�!Uz�c��j�ܱyb`�	SD�=cKsZ����ދ�(�n�j��éೢ�]��xo2��4]7}A`�YY��Ҧ�l��S�m=�g�f�wf�OXA7ī ��G1'&���m��sՔ�ܱ�mM[��L�.N9g6����\���3�a9#p��E"&yT�6�۽��.��2�����k��y��L7Fd��j����r�VFH���޵^+����!�d�ujX�&0��9^E�G4F�)<ü��oٕ���5H�49D��roT9�w5�y�ye�e��{_�ݓ�7�:��=�\&�#'�u�ṉ�6��s�j�v�m߳Z��O,j/�^��ε̳�����i���5�q��)�yZ:(M��%
��L'�ڭ.�pߚ��Q��6#^KM��%���X�œ)A���{��;Δp;(
9�ʩ����|&���yx��ˋ�5��|j�1��K�n<��{�;�q�IS�Y'[��
6*��kt�E�n�OV���/Wa��N�������)�ӇRZ�F;U�����ܴ��l�[ý�
lӵS�
���Σ\ډbH��J|��<?pV�z�t�3I#S��j:ٯW���G\F�KhQ�X-)[�hEa�'Yg�����(�d�r���NPF;÷�*���}{V{5�k�rus�!����G�I�y@�nA���U�9rRnUs��p�=[,І�&�6���HgT�Qꥯt�k���wD���$#���{�(f9�FeB��'^S�f��v:���y"��Vv,�O6����弜��'w�Q�R�)�nÁWz9H���z��Ī�0�g.2�^ݪ�<�lNc����ewe0:��)�b|�p�ڏ�_h������K����]fXK�3hr�.�6+k�'(��ٞ�
��jlN�T��{��auϻ ��g3δ��͗b;��#���\3
�w�g3:v��(���L�\�x^vh*L��Rp��y�u <�LP���e֪��$����O&�����ݭgY�6u;�m;���	d-���o4��8�%�r�P����ö}�6�v�����*o~1�R.��r����<�n.1�N�����O'��Z�'y�
�6yɚ�cH&7�'7ٔ�o{�YS��:(�B�I��GY��Kݖ"v�hnE^>,�2��[t�m��>n���F�b��~��(߉V�iӷ8���5���h9E�c,�[sJʞm���s��G�QnP�*�&�v�:�"{������q4���Z>�罊��������-"���Yz�^1����N#�k('�bP�"�7�F˵]Y�7��"����;��a�x���Y��6�
v[�;9���_ �jq2��)P4�喥+}���Ø�=rnq�p;t��7�I�q��i>�2�;2&��,ȿbn�҆�9sP��Z-���L�.���:&�z���P�38�/bj�e9�����%�n���6T�GVp�X�dҨ����f��CzT�rP4�LM��rn�Lr�qC{P~�wȯ��GJ��V���Ty�E8�.���#q8�s���b�fz������)f'�msh��v�慕���;y����l�T�B�)mFj������H�%�"}T��a���b�!�r�/jg�r�׍��������U�W������x*z5�4��2{�
>��|IǓХG���jP�2�{�Z�M􍽍�aL�F��9m�zt*�3up��`(�YQ�D`;�Nh�`n�'X�Gi�����Bj�+���6�w��49�"e�b��n�V��J�tt9 �\�ܘ��pI�����Q��/��NM��"�Ӂ�)��������3Vb�G[ַ���Nv���W:dU%:j�8�[ǵ�^G��Uw]mv��
�f]��o
O��Q oW�O7a���3�4�:��׵�+a�ý��c����7J:QW���..soj[�K$�X�^�*b�J��%���(�vZ�w;u5�k���:Iȇgg`7̷);�5#n^c�wVe��R�w����K��)��N�T�u}��W�}�
�*�dh�i�M�wݜ.�4�@��gb��25��Fռ8c&���W����xTN�݋{:1��C�0��(���}x�\�2̧���7B��a"���f��)VfC�݄�m�4m��W�P�%��=NЃ�0f���`�I�]C��2���ՔT:��xaע�z^�}R�M
�#Z������^\#7:<��ǋe�̻*2Pp�w�@SX���i�S�dÁ����fcx��1��bXŦ:ȗ�%��hU���'v���	˙�:���u�e�/)�lwpγ�ʔ���^މ�k&Gf�A�N�{q��em����i�9(Ӯ+ٻ��)�&��S&�Y��Zލ�za?v�c�]huN���5�t֍�o��L9زUb"��jR�AV�Ǧ�F��Y;�`ͦ���3� ��A�z9�L�f�k�3����4%�c�)��8�-�x]���1�A����%��1I�f�^r@�o�M����V9���L �寍L���nm[�(A�&�p=.6�ۋ�����B%!J�{X��69{E�Aܡ}:�	5��n��7`+�їn�{%G�@��Dl���+��VH�����c(�p��r��ܶ���>�þ�-i[v�Z�$��4�
X�^8�1�Z32���������8����d-efF}0b�'wc��WJ^D��O[���������-J�KT>s`Q����9v-�����5"B�TSR��%U�r̊�eԻ���-m��V���Z%e���˜�N9��F�R��b��ڍ��kiG��j�6ª[�P�!����*�"��m���mm(�%ֹٷZ(̋�eN<5��-�Uk-�j�j����B��F��feeV�����-3����*6.���T3jЯS�mg�"�^]U�p��^5�T^�TE��ܰU�'.�������^/(�9^2�l���%F�P�Uv6���5��֚�"^^<g*U#h���:-����յ���xp�8ٰ�Q��V��*�Q�H���I[/���D���n�H(��鍃�^'H<��ހ�efEILL�Q2#��`�8`��nM��}҆�o�Q+��wN�X�Ϟ1�ټ-���es�ڦ��9��,u�2^�Z�<d�m�����k5i�K�ާ�XU��T.^i��n�8���zu�=
�g;�>��{:�
Ӓ�muY��f�)8��)���~u���v#�4�ZP���?A�B�yR+�hk#���v����L�i|�T�ɸ�\1`��Z���5^ͩ��$J���k�{mN�4��JF8���������M��w�2��Bud��	��u�Ƈ�������K�}��� �������u(Z�F�9c�X&]�{�z�����|T���oM ��=�`�Y���m����_R@��-�����+��b��k�����7nF���0�����T7�Չ�����NK��;��k���<ySx��m�^H��y��6�L����1��iIĻ=H
��#��Я��;> �DB��q�����<�Ƌ��s(ǈ���3:+���Mx��r��-d��$�;��>�˶yj�Y�g��j�iaIފ��6�[ө3�Bi��ҍ7�����Y��cOT3�]Tz�f�P��i999�st�/oI/rs�Qm�,ʬ\���S;S�M��F��¦1q2�.Z���&�&��b3M�Y�S�/H��Q��ѹ��瑵�&R��kR�[�(�F��@{�V�a�Y�������4���R�lRj�mL	�)�֐;�+Φ&�!�JO4K��MD"T=���c�Ծ�U�m���)Z��%�

���tV��7i����˧t�ed�� ��^�<��k����hM���n�R�\���?o��e龊�Q��]�ŪKQׇ"5̳�#�k�8���i�rrHd��MX^T�N2�y��ھܴj��Ա^o{d�p��pV��W���f'`JZ�lY�\v�f3��یr��Q.�\d��3�w*v�ܭǒ�����e�evǕ;|�)�bBYJc(Aػ���j�����-����!�o�3^EI�^Ǘ�7�&���Ϭ�xMAՓohk{l�=U�R�7��c�Ҧ��ǋ1%�W8�'H�_7�7��]�>��,Y�
�'�}�g�h>KӶ(�9������,��������g��J����J<�+��EƎb�h��nC9H}GºB��k���2��#C���5��Ǔx���E�ݏe3�;[���y�~��vxK�q9��:`Y��l�b���	{-\B.�P���a�Ա@�ֲ�}
⹾B�g�Ir椙��*I�i�;���+̑�f��ch��9x�G2�*����|��V�b�PX��b��w�c"n�y�{�ϧ��9�hF��K,>�g=���h�Qѵ�$s�"I�90�
�5��W*m�dRf_�ftn�V	zz���Pk�d�v�t#�1&'s��J�x��o��>$t��<Y,���z]�B��y�N���y�Q�q!6���BB;>x}��)q%�2r[��=�:�=J��L��襰�VEn�6x���hf.̥oh���W�����\z�*�p�e5w�OW<�籜*��7�����l��;�j��2���Y:�7�U]��uY��j,`� -��]�,�w-�8��R�؜�D�K��g�iE�e����l�;�onN�/w-6�G{����9:���R�n��������5��yl����k�v�[�n�FJ�<{��:��I�
�{Y=��|���9�q�t�+]]ot�R�.��̜2m��ln��ҧ\�1]�R� ���Ch�o{ZǚSmB�c�j]^���Y���2���M���y�I�<���@��^�&!^�Ep+Gu�߂�/�푕�2��{��.	��Y[W�{U���C�򌛹g� ��,��)�A_�����+�H��t_2�\�+�0�|���qŹz��G��Ն�\W�{��Z���J$7^3 ��N5¨ub`ݎ�ɭ��G�o%k�x��7m�*��s9���e�xq���&;χW$�Zh�YI�$*�a��M�Kʷ	ü�M�*�rY3�:Do>�V�-�xsZ�]b���嗨�R�Wˎ��];�8�v��օ:�R��La0�g����_O��]U�3.���Bhj�69B��N����r�QF�;�^Ki�q�]�&w�R.v��C�F�ؚ�9:������v��+��K��,�[1{{��F�����p�3��N�5���㜡�g�3��:լ�fH�����aZXz�j���nkr�px����f"<�~ԫ����y��,�{���P<�D�O�L��Y+S�Sz(N��}�6�X[�5&w��T�lt��o��zx��|��}��G�dϩuZ�������ut��q��6/�U{&r"lau�fTw'�m��+�v�O�PYB�X�-���mײ�~6jJ>P��3��J�ø�Vej�t���\��&m�u�Fczq�4�(&�өv�n��8+���,�&z
RN+�Iȉ'�lyP�t��^o�o"1Cb,ػ�qw'8/-��]jR�[��/�5�k�O4���n�����c�:g�D��m�.�t+%Kt=\��f��ǉ���pj��^�jRE)�x�s\Y��NS�qs�\�w�l�&VJ�j��J���}|��Z�}`��r�̿f*����`�8v�6�nה���K<N���)�ZO?o\ѫ�Ǫ�D���5�gp�x0[�n��&`��N�/��f� ��.�שY%S~���Fv���<��[Z'r�Pm��ޮ%�woMN?
��(�pq�A�ب
)Ɇݨ0G�nYo�k(q7^�����.3�r�,��7�N�~��'��X� �Z���Oa�����^T�#��>۲y��P;�\�樗)�'3B8�4削�E�(�r�:"���w<��b�<u┠Ep�j�x`�~��#�?9�#�~���6��H|kD\�p�<tR����W(�]�j/���F@o�*>N�C�ޟ��o_�)��<D~6�U��/ƫ��nbᮭR���������3]"Ԩz�V*�>����DA�g`©峪NA��KY�z�@��`�OU��j����ҭ#��Xs^;X������=�h��ǹύ�0%�'89Q��u���:
Ƚ�.�_�j��z].;�}����:�\NUV5:o����&=��՞S�>
��O�kգ*�E�Yu�	�ŷX�`�0����؇Oo�X�V�����w*��"���tMEÌ1
���2%�u�Ӓ�BÝ�v��@ԡ<�њ��*����:�n���Dp
��a�Y�Ȯ���ܶ�oVK�S}.����&W٠,f�J9�c�\��9a?g&��&O���G�I]7�N�E�|�Oά�ەh��ꡑ���a'E�������p�s�5Hp'e�$�P��	DUϦ]���;�X��[�=;�P�߭XvxAg*��W*���j�@��4e�^e׆�l��7������!��aB��EHl�A\'b��bb���"(�s:�K��x���Ƕl0eB�U�=9[sp�^Hp�$g�K����^���zg[�S%��mxc�]�Y���9[�6�"7�U�R]�d34��*Y�Eh���oyht+ڶR���TK�W�V�X���T���+���t��2��c#�b�˙X|1U�)�!f��LZ�y+��x��Q^���{n�8qюB�5׺���J*��NL�'%���6pPs9���w���ɏ\j���A�1���čʊ^���j�l\7G�^����&�t�/��{ˆ
��3�s���E孯|d�cp`֍z' Ot�L����,�-����4�/�E��ڷ��u��n��>vv��!�7�򬷎�o�|���g�I�o�M��`dlè�t8�	�"���d�q�]V�L��ٰ�z>V �ŕyB��6k_�����[�jE���J�����]M(�#��NE��5�
�=3F��P��~���37Ā��-Ks�
��1���rb�N��!��ؘ�kW�Ȑ⁘�����w�����;1Pd� ���}�w�W��bѦ2�T]eW�����:�*T
��ǜ�_nk'�.Xu@�x@�Y����X�B&����Y�q�����ƈ�C`�L`~<0����XM��$(��~3����:Ӏ����h�쬦+n];�lqg���SV���cݽ��7�F�;f{�`?;>�e�0'9�E�Q�fF�١��vpZj���3(���k�o��h��jŇ��
�Ʀ��ժ�/�:.M7���?�?�@����O�iR�(*�ԅ�D�I��"
z�D�5SI9O��~�e�%&�_��M�������u�秔��y5���= HCDPc���X�TP �P �AEqbB�����r:����B�XegD��m�����F�1 gcvV�o��p�D�4ʄt�Ъ��*�	nR~�t����?}�����>w���7 Ŋ���\f
"
~h�&z���Ǵq@C�
����Q?@x����;M_�*w�#������0P��fZ?�P`nv|��ٰz
D��J" �|��A�� ��q���*�_sBs-�1�J������!B�f{it m�Ho����r�eN���̇�,J��)V�k�'eI�uYAD��*��'�Ӡ��<U �S���a.������L�m�*���DAMmļ!<���8��8����؁T����.`X6�axlV�@�m��󤷘��h�g��
c�o�ɫ�C*" ���萊	�=��������6wѹVOq��:�$p���=�}���"�n����vd:����^��86��DAM��@�1�������d6�DjI�Ձ ��T� 

Xb�ܢ"
{~��@�8-�8���@k��'UC�s2,��	��tUQ.6�" �@4hF����@E !lJ0B���\0\y�SE�g�Z�����xC@���ae3�kʋ!�j�"
f�a���=Z8%�DAH����V6=� 8@�ݩ}�M�@|�?�Ձ(s�5VX�T@P��b=Zy=�b�<�<�O��Q�+����8��m7F�#�I�Dy�}a�Gx��)+�X.��d��}�3�<5����h�����<8D�tȁ�$Q"H.��C�vO-��D����&��́���Dyx�fT0�w��:�l0""
v����@�.�`�S��2$�l�:7#�8�HRc��"�TIJP���F AO�:y�Cp���7��78�ٱTD�C���p���_\���b�+�[�Ҕ�p5�D u��%C��H������H�
����