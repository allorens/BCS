BZh91AY&SY��Ƌsgߔpy����߰����  `���>���  @ 
�N�[���@Z,z@�� "(� � " �o�@P�<>�$x @   �   .;u �� >��E�7�;�޷4}:{�n�w��k�Zd��4װ:�m��
җg.��n�'c�֔�95:�O@i��};� ����ݠ�����Z6;Ct�U�i����pι) ��j�#����aف�ItuA������N���9"駀|�� �{�袎�R����E(5 ������C��pҝt�w h^�ttv�MWG��8� 
t/�vd��a�v϶R��&��p�7z��tZ
4R��c�(ѻj�E< ��7=� ��9���`�z)��;��h)�7@t�a�$�l
���[                      J���T�M b`@b��)*ROS �#�����!�F��UJTڍ�4h    4z	*�L��	���` #	����� &�!��M4�����LS�ɡ驦�m H�aJR���hh�bh����b>����'W:��9̜�*�V��:~g����[��gٛm��zt���~�ٌof�3q�c~L?��6��7m�κ�������o�o�������>��?�>�
�����cm��ݣ��v�䫅gݼ���a�?���kY���۶UUFv�~���c������o��_����3��s��c��mtA��ؽ�9�\�q�lQj4q��R&���u<��$���%�R���<��A��f��V�9�:씝���9��O	�gh��h��/ƓW�u=��ٯ	����=#t9'���I����'q#��Ox���X\`�g,~]��!d��X3�|�ĉ���l.���	��<�Gg���{�zIgH�A:�Aę��lp�����og�-�&����h4H��B�!�IϓC]��7'��i��8�P��Y6Jd�ɽI4ɡ5����C�G�zN�I�$G�	<��'��8��K=�J��	�H�Ad�D�ו<8���7x�j��vU^<{�Ğ/ŞДs�D��dO���~����%�4�&�^�"{i<t�xJ���;'��P�6"s�;����>ׄ�	ݤM�"x�I��vO���\"%�'S�I�D��DJDGŔj$����C��D�Y�BlH�'����'�i/�<p�H�Bp7I9Ĉ���<'_��vO��%�+I+�)I�E}[6�����e�A����C����DK�e��J:�>Ft�h~ؑ�D��&�o��$K��$KN�M�f�g�(�'7����"i:y�>Rl�wAZ4j�$KX�HwB�k�"lN�nN,N�f�9�5Bn$N'6%'GЉ�u'�O	�H�-$�Z4vw��GӢx�Dd�(��Qh>�\�J=��}bz�>��tx��(w��c��7b/jP���"'{4>�%��6p��*�6I��w�~�q�d���{�&ٳ�6V�؍Dz�H�>��p�QR|�KN'S��' �EoC{*��(/v�w?i~Ə��������q��@�a��G�G�"���a�i�q����,'���l]�>�����5���Q=s�=֧�r�d<h�:2�#|��"rғ��Խ�u7|��K�S�Y��
�������M�<X��D[*�	�[jlJ'�"�tl�f� �b"�D����Q�D�ԣ�F���",�N��SB;jY��FO:���bX���DG���7�(�>���Q�j'��J���b&�ԡʈ�ڞ8RI�&�'���"<$Dd����"/j'���;֥�Y�pz]n��8#�TN��R�2|��U6��TD�ږAg�FUN��7ʉc�TD캛 �|��U���ꈝ�R�,�8i�J��:"V�Q;�MJ ��#�TD�ʔ#=Q�jY=�CF��}Z��]D{ʉ�N�į	�z�z�N��%qZXB�L��'C�|�Ã)�Tl���7�
�KJ'"u(���� ��[Gɟp�H���ñ#Ã��Tpu��7[#.�>�OjP���N�'Kn���Eh��_$��!�f�g.�p�~��`b:�Py����b	Ԍ3ӑ�C��Ge�M�)91Z=;Q::�Dz�'ue#i^�QDo�,��pյ(��Nu��vt�v���z$%@�<ʩ�K�nl"ŞF�wȽ�tCh�D�LEs��y�^f{�{�{�w�x�0������L<�����k����Z�jC�k3z3�0�L�M�r3m�
���{v��#xz��F؊�F�*�����<�Fv�,��SQ(N�<y!�D�;b��فJ�<�{���EQ�=����p����y�G-G���Kd+ݨ��հ�F��}s�dBjC�7.��TF�QgijV��S�G+��9|�i�7�sb�F&�&����b;����w�J�ZNr*��#�r��z!�C5��R(�Z<R=F{�#�y�=�'y��g"���P��{�3�A��.���R���|b#4z�a�������5��h�o�B�� �G8h�'�I�f��͑�J�C�0~2���7=]Vg���Yg�MU���.�X�m�Q5�ODN������lM��+d����;R���I�ץ|��U�DN2N؉�I,���DKY\4u�%��+��J4��Q�%|�Ț�UDG�Y_?v�lM;���r�r�h��H�R%���G_�#�J�،4Q�&��H�bP����jR&��D��D]J�c�J���MwR�M���둩I�ze}_;�����9�WM~�,u�_?,�4i�"[�H�w+Ƈ_O��R�4�U�D��Nu+Ŏ�+�粑5�J�6�R&�Rpޙ_W��&��=x�/��|��[��H�>�%��܂B�JN��U�:5ҳFU�4�t7�(A����g�K�j�p��ü��ƥ��9Sf���D�O�$,���&���W
"�}i������oeAxOy��[���x�Mvy'�(� �#��}��T楍D��%'�;��ѾU&��N��UI�쓧�����l����G�<k�Uq���Y� �N-�*"0���J���Xz�2�<��l�O�麯<�qv�i�L�:غ�|&����OA��TWj�+�EjRRO�'ԓ�+��rWZ��$�$�$���J��Jv���Jw��i+"i.I.��#���}�_rV����0�=FQ�q���k	d�"���"����ᰨ�H�t=Fu����hޜ�K������n6������x�����>I�)�������
�C~�_�5 C������>w��}}u��ף�U�t�Һs�9������,���e:��
���Z�$���B$V4]7FaTUƎf?��"\{#uO7^m�(�g��)M�ݎ|)kݬ����4I����U���hُcރsss���~��������t9XΒΒz����h�̔l��L�v��AB;q�/�ѕnc~���0���ة�����M�)�f����C&V/��j�y�e�f����Y�c�uBl����߅�Vc�8~���Cᆳ�F�v]s�>Q)�4�kF2�dIm-�Gf,���/2�M�n3E�s�<߫���r@!�&���[�H���Lg�7�j}d� o0�	�:4af�,�m��-����q�r_͟�|�t�����Z����@�__;4oB#�S�	��H�o����p��[Es��*���Z_��d=���2I���,�0���|4����_nTϚ?Lw�ϵ�YK��!
g{�	N��Vc�S�N=W�x*����17���K`$7�!�t�J$7o��V��6K>k��)�t�N��;�kr� و{�krkӦ�C��������r���f�U�L�4��nYX�����܏(���$h	��D�����O�8|��°��B,8b١��ԧ�& �æ���e<�7S�� ��t�!���g@٣��9��;��:%�:h�ٳ9�O�l��Æ�k}� C�QAp��t���t��'�F-63��S����jp�;�AW�c�@��%+��C�4h	l�@(�4n4�@td6h
pቚ������>>4sC���Vb�B�rv���lJm�C4�b\C13ll�Ğ�n'lŲ���5ɋ�M*�v=��K4(�1^��|~83,�-�	�VEI>�����َj%t�֑s���2�^I�UОp��]0�F@<%�r<�}10����}tůzbd���LLf��](��	^�&�1l:5zY�F��ݺb4��!���Y���yH3��I�ìv�08����t��h�Q��cT@;�xa��	,5x3����Q^Q�aң�w�� Vi~aB	D��[[h�����IYG�e;j"$v֬�4@<����؄�Z\w�of.K�t�J%��=����d<x��g����]1t�W��r��1�ӦC��l���M����[:d��2�kn�|ۨ�~{�D�m��M]�|	���?/���?6q�Gȭ�d�g^�\��oYM��*W}����d#b�Z��Zݪ|YU��p�m�t�J$��Y��ݍH譹,K��eS��O������l�����t��!�O���k�|ɧ��Y����!d���+�u
>4:I��|8�t�<��V8IX٣ƈ(Sm��H�8t�:����=���(h�
p�њ6@Uã�ٳH��F+��1�p6	� Ͼ��>8C8Cf�l&��p���d)ks��8u7�뻤yzݚ�zB�8x�)ag2��,��ó����ف�tz"h���MU|;�; ���/�	�LK�Sf�&�(�s��g�͚[Z(5ǉ�|fV�q��7��g�a�d�����>x@��3:���6�(  Hㆆh������  �be'94xٲ��N�!���<C�Æ�l�Қ4p����}1t��!���l�6pѣZ��4bm�p飧^�
3�)@|����ލ�3g �2�<YeV6�Ӽ�l�M�6us�Ξ8tZUݕ���b5��ѵn�$o�����<bf�o���p��g{)<p����p����tt��J���u�SF�{�f�C�����є񹹣d!���!t�l�/��`W&�����p �&J&��ݛ%�g,����U%r�L��W��Vw��Q�y���^["�L�I�tg9�φ$�MJ��vt;������h�O���H~x𭯲�%�2�:>\©_2aZݝ)Ӈ���v|6�uΪ|x�ʎ�6t�s�N��K9Aq&��0��0ϭу��+S#��ƍ�����!�.�!�:tK|l��j2ߧ������Vѣ��Ky}XQ��:]cF�q�f@�%g#]4��X�&�Z��/��"b�n�� �F�:MD�!���)UsOBo#9�*�o{kw0���n2\�,^[�N�?s'	$��FT�AH�GSv�f���TVb2�k�͖t���R`�Wk�����am6O6v���匐� �D��;���(e�0;�>n���F��PU��Fن��y�o]�39�yզ�ژhѣ�PJ:K��GHi�Ⲃ�������yM�l�>yl�@U��h���f�3�����8lwSsr�n��<;¾j��&��'��h���nBa�@xc:k�������*�0�k��K<Uk(-:Yg�7�\l����U�.r�&c�G*�O�e�,�#� Ҧ+g�&4"F��0�5M7��qS��6l��F�6Ie�<8IϣdV��<z�vp��\t�|Q�k�
,�ѣT�+�o6l�Bj����Ac�B��@�\eϕQ�,���Z�R6��I(��+z�X+��l��ΊUk(*,�#�+9�캹�{S���G��Y���A���&G��?O���?���w�:���}�����{�F?��D��Ϗ�#DP�ut���G�C�\u��|�p\b�s=��ۥU:ԄB@�Sf1*�II�ٻ=w#�g�qɔ=���&�b_�S3C����D�WQ�F(%�Jƒ�kU�SCR&�w+�N�Jd�Y3��Zzšc�1��ԉ�е]kP�'m���hZ��P�h��4,�lX��B��ZnQ�J������uuqV�҂5��'Z�LI��hT��I�d��8��<j)n4�I�˂oJ������L���e� ��l��&a+q.Gi�m�ݙ
(c��t�i�DBe"��qh�$�f�j
K(����,�;4�z�
Q&4+;2�����'����Jy��w��.oZ�Hj�*0���1)��sǀ�x���G\���ٻ>�p'�����:�=zz��'nP�HOq�2����#��n7|[��8���^�0��%-J���k���T�u�-mhR`44�R�G_��"�! c�P
+L�Ţ����������@7�橄���SI�O�L���'�!�ܚ�.vPƅ�/05/l�6�u�pݠt��l�y�<X^y����a;v�1�\���:�9{���=[�uo���ǎy��x�&n��.�՞㩽�gV<۵���:��;_V�S�n��ly��5 ��ʶ��d0M��16�`U��:���g��{��3��Վ���՞m�OW�՚�s�ǻ�V��k��~E�������__d�g;�lo��ݼ='�oǻ���}����o���~�e�m�-�����Ww����ϙj��*��b���*��t��U����X���iU^�UU�+U}U|���]*�Ux��j�X����EEUUEUUV�U괪�V*��UW������V����,+m%3rm̔6���I[���o���O�� 55�U��U_,UU�+�V�UU|�U�]��Ux��U�Wj���Ux�*��]*�*��Uv��*��iWJ��,��UWʺU^*�UmUګj�U^+J����z�Q�sfp�em�LkXS=Y�f�P)�D��e3h������'ć� ��I��֗j���Ux��U⮕W�Ҫ�Ex���*���U^+�Ux��V�v����U�]��Ux���]+J�����V�dUWj����t��եUx��U�U}���߿[<ٞ�Xq�[P�H�[dXKejڨ�|���V�39��U^+�U�]����UګjҪ�EU^�*��Q^*�b��V�U_1UW�J�j�X����t��EUx��>�:UU�Ҫ�����������*��}����mʼMֶ��o\�%�PK�ܶژն�6)�A���][l��b����L�ՙ�m�nMɷ&r�Eہՙ՛��jn��m�{[�:[}ϻ�3~}��%UIo����_��?�a�������_���zw~w���x{vy{y{v{x��<'��<t��A(D؉�gH �M	���O��-&�m�Ĳ �$,DD�(A��<X��%�blM�BP�d4FA���6AD���tN��E	�	�NDDN��AD�,D���t�,�DCB �'H"I��"�?�DP��!G����G:�[���;grŐ����s���[ۓc��v��v묏2�u�=�����=�!5rD�b!�������]�f�K<��j��k�ٝ�p=(����O^�]=w/a���j8�=	��x�H�^
|/���[]	ۚ��a�� �OU�:���c�]e�gsFw�^�ˎi8y��`�瘚9,=�S���r������n��d��z��w<�n���mù=�q3�8&}�>��̈́�w��;^-�ڛ("!1!Z;#v1kJ�볾�8�v��v�Nwd���n^��nWT8���V�v���V���փO0+&���ne�A���I�9�N����<I۽������ϵ���sb���;*z{z�v�8esZ:p�Gk�S]���v饆�]7(W�5t�Ƕz�u�YM��eM��t���`��9z��>9�p��K��&`���a��A�Ǝ͎��n.�g:��8����O����m{QV_Vh�=]n��]�݅���UvpdYb�n:v�X�j��v�%�M��6Nz�޵pV���G�6��{u/JvS�9O7�E�[��ttɸ`�y�\�[���'�9猏n��j���wϟ.��/f�|J��6����.:^�v�۝"slJj�G���ɦ3
��7U/	��;���ƪv�'�y�Lq"���y�jM:9r�<ls�g���u�ζ� )N7���p�ˎ1���5;b8���=y�n<���E�uө��v;�.+���Y赮��)�\zx����Zp��r�S��1N^̩q��"���uHmq��ަ���p��)��mk�;h�c��OcqW>�{S�X�"/ca�<�M�.m.��[��Mh�9��6)L,x*�r+Kb�ilJ,9������V�����1bfε�������j �úyӺǹ9׫C�M��S�ۿ��۾ntp��b�wW=�msָ�g�����s�/N۠���3������7imӠ��4##��K����͍�h�9��<��w%Am�6�v�����AW[�r�v�Ky����mtZ�tk;g<�k�V�!8����{�{�ϻn7&.����Y�<2�ӻ@<��9�6ذ��G)��;>){ �uCi83���xL�g�7]�j�GNys/\�8���<�\�m��z�z��]�n�:z�^ƻj㞾|���/�	�6#��۬��b�0noa�+�:�Mɝ�{\g{v:q*���qڹ�&0b�tvն+�厝FݳΧ�չz�{R�t��5��ܝFN�v�=g ��v�F�m�2�M۱��ju՗�k�n��[��ٞ�c�N�S��cCV�/]�zsi�q��]�UۍH-ۮy��˸O%�C�K��k���̼r�8�g7��{tؔ������՝�I�z���u�oqG �C';�v�#*��h�+n-�)����b����ݹ��||a�������wwn|}��|�fffb����ݹ���ffff**���ۇ��}��Y��Q�ƚm���Q���2��xζ����Uj
F*�r�"�6��.�7�V��C��Th,^I�b�B�4�[����h�Ȏ��ng9m�y�a
�.-�5��ԙU3,��Rq��*����3��b�-�ˮy��N�5ռ#��ʲ�w��$5���Ѵ����	����X�
�烾�y�`�)ֽ+�J��{[;�����(u��x=���#3g����Nܤ�l��U�2���wgۖ�`��Nf�:��69Rj��n�]<�v��1�:Ƙ������{C�ڗ7y9mfK���%ނ(�f*G2�l�gGyx�
0�-ͭUxۻKc�k(��m��i��cv���M�(�h��E$����g���on=��'<��;��.jC"��>��t:2M8I��D7�p��!��D��x�ln"��F��{ѓ�#ƴ�E"����H��!8d�N�%+:��5~�$�x�O�0�
0���Q�K�GI�6�l��(�բΒ�#˄W����B�6���J8i.�"H.'\6��xb �྘��j(��Q��)�������V�r�iw�:x�ˉ�����<A
*�:uXYrϵ��g�6lN��aae��ĜL$=���L#�&�&E�0 z|�qY"��T�1�b��b�Z1 ġ��|��t��֙C�p���B$���f�")����yt���w���ڥ."�"4����+�o���f5������ruY����I ��J��|{���@�ƶ�W;������@��b!A>�ag�ӧ<a��0�0�,e$�)/��9K��m��:�Zꃤ"�D���kY�iLpM��nE!כ卅
��o��Ɗ����'�&6���p�CD�"ާ�:J-x�dt�w����.�8�Ba�#�8>�6�B%�E(�OY��Y�XYc(�+���>�<8�y�SY��[֪�Dn�SL��Qk]�G��ˌlQ�9����$�E��N3�pr{�2��i�J��5��w;e�d�j&*��ʕ+���1:�f�%�*�w0�����ښ|o�Պ�fn���b� ���clm.1J��!&�#�ސ`_�}
����g�|B��1s5�M�F���r�Q�x�	G�
E��<�0�A�I ��" ��J ���
�pڨ���lB��D�$r86.�F�Tf���\�1��0\,��xO	�:'�ǈt᣼�%�4�<���� K{[@�Ky�φ�{��,W�@�QƠc=�mu\8t�E����(
<�N�:��tcL(�/��������7LU|q��>�:�Q�'ؼ�wF>u���G[m�;(I�5�AH��(��\$�(��afaFX�<JR�`��G'-����3ۻ������U���K��,!���6��mJ�A�.�C=��c����@�p�)��}�[-$a�,p�|�`�|��O��_��y@�����	���"�;g���VA��%u3I\�e����xO	�<<C��[Ԏ(���k� b1p��F`�I�࠽֤�Ͷ��̫�...by�G�<�"��E�q)D�������td"1�j�t�#ē�V4j�8u��n����M�-��C�ܩ�d	F�D�bx�ç���F�0XaK�.��(B2��5u��6�{�lPK[�2'B@�n*�EaH�� ��TWSU�=z�O��j��7j����)����`���h$+,u-�Or�\���S���5B�xq[W�(U�v��z����V�w�b���]]1k����f#L�ߋ�竝�YӘݶ��yxw֕];g��Z��(����*8q�c��D��lTj�1B����gĄ3��� �B���DP�6�~�l�N�	T��B1Vw��G���FaE�Q�<'�����:pѫ%�~��6�m��b+����^���k����V��UIU'�:p}�P�
~��w��ms[<3���t�A�����*�֣C΄�N7��װ�b��:�1&�0�Ӽ�"%J�BZxm��7ċ�DfC�$�";�I�.겈4f�ќ>!`�kp�t?�Q�+����h�4���i�<�I��O�>������=�I#M ��h�z=�DGĐ��|9> ���gǈ�lz=0�m��,��4�<B��k�����hF�IBRL&;%a0�DÆ�L	��a���L8Q��`��
I�h���<=<BӤi�#����(�'���>�6�#�	�4�F3a��4f��Ti�p�x2�!H�96����I=<F��5��¸UL*V�T¸aXORa�L�=Rp¸Bɩ&3FΛ-��65����C^њ>ӄ�]h����;S0sZ�w���&OQ���?��$m�AD'b�Л 6�<N�z|�����*QO�ȫ�LٯN��T)�|!L��0T�Sa:L�E$��;嵃�<�&�6���ű��Ld�H��ۆ�i�V:ǳU׭�ؗ�O��}�6\��a��y��QU����Ϗ�32f�3�U����}�}��39��������Ͼ��̙���c�ffo{����g8p�0��xN���򫊦����m�������>��˸QŴ�̇�:M�������rܶ}\�vo�*��zxĚ���Kk��:�޴x�o]9��G~�9rr�Y�;,��QJCD�80���s�(���G'�I�b�!(ag$�"��84K�[���=,z��ywα��q�I%��)@�PҌ�pJ�V�@����<R�SKɍ�%pb"^crB�<�T,ͦ�I{�@P
��q�@ѣ!!&�i��x�J,��`i��J8�m{������smgg���u�^u�sg�۳���bf}e��)�H�F�
��E��(�Pp���Y���N�:T��=�gIo>;m�X�������9g9���se�7q3�g��m�v���7{�����s8|�i�x[;e�2VyG�kx�;oN6�O�ۉ��͸��>=�;�|�;��yOV�	�Nwst���[|����3ζ�OZ��On��3ŷ�j&Pא�|t��4�Ř|Y��0p�>8���̾1�EL��"�"ϲU�peѪ Q�,�6̳��z[���Em�;82�5D��v��I$�H +�]{����p}��kv��o�f9�:Ζܕىp��<v�Ȳl��<9`I����m�U]�F!�)m	UW+�I���j���f��v�,h�]��r��v�W|=7�&y���#�R���E�� X>;瓇���f����8���mo���߀\��cþ�w�V�V��J��6y�=e��{�s=���c��3�yY�F���;�]n�N�/�e������:�v���m#��x�'��Ne�Ώ�g���g}d��ӏR�K���[����Q��hc`��Ã
���g��s��K93'���V#J����z�U����q4��)�!�Z���4��afaaf���*��RqR)�.�)�Is��8�im�Nr����H��=:������� ��3�CH�/'�soV��|���M��k��X��������};�,;'�m�I�g�jo�ә�D��w�o|�:��q�|N'V�s�#��x�1i	~����Y5߸
FV@��ݫndv��A�=�+�����z�n��g�xO9m�{�0KE�4`B:�KL��i�!�w���;;�Z3��K�vM�c��*8Q��O�i�faFY�k��*��	/F�L�L~כm��Mb9P��YQ��33�M~\yf��s<;q��s"��l���vG|��Y��yX�G���n���e���m[=ۧn�:ϖ9���ì���w�m���f�ŕ	i	>��*�v>�+rZ��۝s�߭�o�mշZ{������l� ��A��R�B�YCgSR�����t�Mr�<[�I�o��5m�����yG�����|��<EHH���E�4��b+��nI�s=g����N�y�{���m�mճ�x�x����3~ێ������i�Y�Q���i�p�B��śB�R
��E6�I%�8�i�['Yç\�ϥߒ�Y;�Yf��:q��+�ݜN9��P�x%0J�M%�%�����p�[v�Wt��)A{i.�4bBK��;.md�:O�í�(�˙�X�q�,:�C�I�S��m�:�t��=d����L���wN�-��:�n���w[nM�3�n�=u�S�4����$aE2@��:�!��6����k�T,O1��p�À�Uz1�IF"��Aф&)$ ������>�j�Ծ�������q��֝#�px��D�Y��g�4��0�,�(�W}�*"�ۦO�����rM����b���O.���W���C�0� ��uwrI$�A�
��PZK�-͛�f��Tr�X˽��9��[�U�[�M��℗t�^�vʥA�M�ل�c�m�W�v��՗�c����q2�i~Q�!�Fpa�k�B�i�v�LC���qF	ځQN��u�m�\sc�-��l�����x�I�����
G#�=pz�u�Y˾�mm�y���rq���\������:�e!�6lo�0����v@�F���	��L���mn�>5���>,�|�nm�u�v[<&wL�v�mߧ
Γ�wͯ�#*i{�yG"*�|�ϭ�l�����}�)C!���d�"��F������<HƐ����Z5R�6�0��G��<|i�faC���G� ��}8�RYj:
Y2�"""" �:����x�D}��I��wv��o�6w��'N��o=>k9��x �Β_�jF��>y��_�6���W]�����t��7n����Q?"Hixa���"�x�^<w�ov�rvvp�ŷ4��̺��s��i�>z�\���w�;p����0��\1�"	j=�:xGr;s��N�n��:_Y�x���s<���[շ<����7��𳈚AI�׼@֗ë��0"��,��i�faFX�,����=um�52v��9�s���7ȥ��z�POeC �֍5�����q�gHY���-����v�#Lxpz[���Z�
no��Zc{ŽeBWY� ��&nGR)ڛ�A�Z�Us>���1�F4�)������+w�wl�s��^�s9�vݳ��:۳��7�g���=h�w�y���SGFy�w��D(p�<���}���st�2|z����[���׆���n ��sC�H�e�Q��||Y�Q���3K(�9�XyP*�q$�I$<Gh�����8��D#�u�4pk��hS�rqF�ɼ�n)��+����8�6�i�WWBhc)x�]ܑ��K��$Gl��ך�޷no^�q՞���= ��8cl�4B^GQ�e�7���"AG��$}]8Km��R�y�/������*<J;q�Q'~�o���9��t���},�]�����v��rS�g4v�۷�]%�>D
�	x�)/!h��4��|8X:�(��0��A��0�4`��&x�0��aH��Q4�=�I4��#Fh�z<�Ѧi�#Fp�4�t|GͿ���"�n�Y��tz?�pj�٤h�[�4������i� zG��&���������i�Ɛ|G��<=<BӤi�A���f�M"�A�7�/��]֗Ҫ�N�r�_I�s�7њ3Gѫ���4z2�!H�9���xڢ(zL=#M��Y������(�!+	���°�0�&I�G����A�H��G�cѱ��z�g�!������F�xgF�z��A�Y=ʾ;��U}�\�lҺ��ʡ�A#K�{t�V7R�-�YV�$#wZ�Ė�+�']w3���j�']4���V���v��4��v��bg�&�`.�x���҂Y�Ț7Z7����23����E|�/Ym�E���g�W*^K]X�"��-�v��tu��=�h�i/ ����+s,H|˕��Ȯ\W��;��Q��#N�¶�L���B3�e�LX�
�*P.J���]!q*�TN���<oM��K��/�|�Ͷ�u�ւ�y�r�lX��t��7π��4�y-�SC�h�N��JH��,Ex�Z�%��Tq����*�{��3�y���s������7ww��9��32�33����o{�ff4��V+�˻�g~�̬��ǫs�wy����e�8a�0������:a�gNM�96v�n�v:�j���J`S�f٬U/`���93���N���;!��|�t']��u��:.9��;2m5�G\Hz��V#m����خ�����ٝ�;[q���n�m`�m��#�4���&��c�-��ݣ7>v��ɝ���݆�QWA�x��q�;;�N�덮��]��1m;���ɀU�v����R�oI��n��hU�[�Y��稜s�'��WX5�q�q�F�U�,[n�^d�{�L�ö�q���v����\����䡝p����׫�ۃ������Tl'�����z���q�^k��a�ҷv���m��HZ�׾��k��!���u��x�;�����M�ɎEw�+3jT2jQ�2���������J�cq��jޕ�-���2�Y��GmZ����Q������7r\�;�����ηt�g���nq��[;N�,tH��P��r��!�J�DP�2�(E��!��T4KK=�����+i���Ӷ[��⹟S���<gIF��{�em�ĝg���^9�M��n�/nv�#��ی�g���	�%+>�����>U��~��9:v����8�3F�J���OIBd��P�Q��_&4H�w���"b9��o�Sz	%^0W%�B�O2�qi�(A4@t넏у���a��$�߇H��h!�JP�gO>,ҍ>?��<<C�6WQ+T�<�s��9�&|���s<��mN�}m�:�\.���F�VJ&Z���<����8�*]c�9�t��ͥ�>���>�nd�s>z��Wgv[{t���z�n'K!�gH8�k9=�s��D|�ݓ�}ǅ�w��xN�r����^�ݑ�ړ��׭u�SY�_���3:/#*�b��ƉcJ!6��Ό���:��X�}߇{n��Kt9����G]ms^<�R5ᣪH@�A��A6x��4����4�
0���Q�;�y�ĺf�S��,��T`Ƴ��Sm���9�:��<��n�˛��=�����sR[:�}��=���Y�[����َ8z��o���[�+�uRvy,�󾳬��:s>;9�4|�s���Վd^��Ź:�͹9�mv�q��M�p���I���Cp�U)����kG���Օ�����n�3����J��<#��7��d}<q�/���A�e�D�%S_#�v����"�<������h�b�`�X0"��s."z�h}�C�[r������1Bh��:d���&Kh�����L8Q��i�f�aFX�4��m�.1�#Qi�z6�m����B]�v};<[ñ;�e�ㇽ���t�~�Ff��[B^�i;+�I_�T��']yw�Y�����˺�:VQ���|pCF���Z���{�%�T*ȳ�<mYۧG��s$�s4�vNv_;������8��g7��쏑�8���{ugY�:�V��'1U��)Q���!\�gy��D���u�.��%�:�GK����c��P6�Fb�J<Y��||i��aFX�4����H��v����!ζ �F[��bFS81�SS)���rF'��î*3��~��I$� w�U����bW�r�ڨL���N�X���b��\�>��=aQŧ�1V�wV:�J�f.'o=]�W@��a�T$��V�幗y,�6�t�#�wçM��Zn����h�����ݜ��Y�x�N���Ŝ㙻����!��4;%p���0ϫ�ǒ�fJ80�KCf"!�jID�F/#j$�_�Ȝcd� 5��O��\��E#�O����#��h��	.�D�x����JÑ)�@�Ԛ8ID�:�	�A���q�=H����1\�U�24���E��i�Lr��ME$��"j����3�����4G��;�>HkZ!C(��J ��L>8x��J4��0,,��iG�Z2�s�ܑ6��6�m����b�?%TX��+Ԣ�ӠCFO��.�g����h�ˈ|��WBM	vp�#��A��o?d[\���No���z��Vb:�8P��{�v�n8{��g~�gyxx�|���:uG���4xJ$juDN�=31��x�M<`�_oT��b���jV��T��%
A�J1�Pw;;��[�N��w��3�����wr%)EL�=l�Ƹȏ|x���(����M4�,e4�^.��m��BK����S�k�0�"���R0��J<qI�HHͦ��UL�4��n\����kx�IV�p�u@r���CXa1��A���s��m�(�©f'�TPG�F�
HR|����5��ڥ235�))B�0��D��V�P0%��"�}8�4�%E���Ðu�ˆJ���ޤR(�]��"#��CZ,dO�.)C���A�~]e�x�Οa��i��`��=Q)&y���$�Q4����d�"<�.��B�.e�-�t�q�xݜu�.e�ÿ��Ւ �Ai��u�t*�m���(�v`�����:���%
�!B(h�;�nM���B�L(D.��H���"H�ā:��*N(D4@@W���(�!��s���
�N/��9�t����N��ǵ�Y�'��%#ҨÈ�iuI�@�f��K!!M��u@��GNi񧏊>0��M4�K,e$m�Yy�K��z-#D6M��\54�P����**J|���$�I$������l�z�"�q���l��tb�;���#�ǻҕ&���-��E�%t=B�j��#vzZ�CU1V��ʹ����mo���uܿv�;݈����>���8��1Y�Hs$+�ב(��[�Q�q���Y׎i�{�Z���n��ݺr%qO/�V��7�N�!��$��n cmcl\9�s<��U�CɼW&/wKW&g����ገr��|;,(Hh�mL���4AD��!�H�5GN���/��G�~i�U��j��[n�����jgk�ɢ:q�G%�%�Y�F>(�O�4�J4���Q�GK;"fU3 �/J�"�F�[w��m�щ5�ȿ#cƶ�Fb��>�RgQ(�РW܈�PZ:Ȫ}y��a�ީ!�ĞB�A�NU�G�N*�JZ#�l!qB�up���\��YE�I�,���$�qs�m����2��)$.=Ρ�x��r�R�8�!��<��$=0�>�}�硸�\�V�Ti�|;����á��4��h�kƘI�4J�$0��aE0�0�"`����=�M"M#G�����f��@�p=$�FI�h�:F�[z:���?BњQ��Ğá�������$���N�G��n
aeQ0&VF�Åa�0�&h�(�ep�l��h�aei�G����F�,�-��Ë���I}*�����\�q�|[�|^���|_���e����eC��zl�#G����!��`�YTaXeMh�t�0�&L�`����x�<3���oa�h����a!a(�¡��
&�|>��I	|tٗWQw�KrT��MM��Y�nj�]�Գ�nq�3��6n�c��۽���9F��7�V][t�-��cI����u�0�i��ڂ��΂5�{��Ge��>:W E�uNsN�U�*Q�1��$�2�yi��hﲶ��k��s[k�����Պ�˻���]*�*�]��ff:U^,U������t��V�����p6C��p�f4�L4�J4���Q�Nsb""""��1�)� � ��O͍�x����><�%�.���{Ͷϑ�W#�JX���� �8�����}��0>�Z�E�䝣W�A!�T:���s>��>�!m_�`�^VI��I��y�8� gC�G~m����~3���5f�k�O;����t���!��@[B���Ldx�<�J�����28�TZ8sO4�O�<Q�i��iae��đ�rLPQ��U���m�%�#���D��>�,��Rv�I\ ,��9��~���[mVZԚ]�!}��tC5�qQДK@��%{����G��t�0������:|�8HQ��D@���D�G>$��?H�u��Y�ep��_�Y$HK�\k������(���|i��iF�X�<I$��g����}V�1�Pu��v��M�0"�/$�"Ҋ')|�I$� :��3;녓�RBjZa��6�HkF�&�޹i�q�i���W]��J�e�:��A�c�VI�a�	d������Aɨ�ls}޶�t���I!#�"N�k��x�#�qb%/�����R;<QЮ66�wŢ)��G���.����"*A���9�8�2�&��W��\+���dع���m��%x��1y��w;/�Mު���ӻ�\�O�N�_ o��
����p�8��tH�A�^�q]�����h#>R���n�[�,��ƟQ��i��i���ǈj�@C#��������"�:1Ĝ
>)]!H�
9�ou�L�(c�<�_R����|2Ѣ_3 ����)t��+U|j-�ּD���#��U���(c,����%��=N8�T������)R���8xD���G��5��p��#�6Ψ�+���L<igƟ||ifi��`a��)��j��A/STi?�I$��#��m�r��Ȇ����883�!$#�!t�����Q�Ky��^!�3>�x�o��ȈG���?~��ZB��ƅ�R&lP�A�|)���i��qK8P�.����3;�w;��>���ۖ�.yvN������\ ҩ�E3��K~-(3����a�d�w&�g*IY����v���>(�,���,�M4�L0e�=��%f&2�6����m��
g�D"���:1�����ᚮ�B�f��`8?ϱ~,b,��.�^Ɍ���J�b$�:5���:3�-#IG~:�����6��1���e�z˰�ۜGLE�W���@Ƽ��h�\<3��������壩pdꦵu|���<Q(��>0�a�!ㆮ�����>��q���[ݪ�li�nL������Q`I��m��4.k�}��>2UO�����f�E�����otX�5̃V�(�ֱ֡d�2�[Ƕr��!����.�,��S�)�;���E#��,�$�ю�#��p7��ha'��wO�����cc�z<���}GFt�1��G�����:D�3�}�KGPӣ�׎
�@�C/����J�8b�3���
T�Fs��L7����RkԠS H��3������ƚ��T�hWg���yZ-xãl�"Q9<#�*3��~:"x�&a��D��n���D����TuB�=�$��s��K>|�o�w}��:��']뵜
ç����<�u��cz�G���F
I���aӣ�3��|���}CPp����Tf�^# ��?1���⮪�J��HJ�h��V��td"qq�dA#-����-GMb�I��^5I��T:i�Q�&a��D��}B��kUG��km��ƅ̀�j�P�� _��P�>E7�)���o�,����N�}����h��b�&l1z"!x:2�j<��ys6�#��I��j ���pcLߑh�VyxcJB��jga0h��y�1����F��V�#��I�x�>?~���i��XYc(�^��nx-h����ۊ��W����m��1�2CƮ����<�x�N"Qd/�5�]���p������q��.���A���>>m��b�1��yw�zL/�U������61���Qaf���4�!DBp�O�È�Ȯ��Ç|@΄L"N�$�ϱ�7� ��^�<��m�A|:�VV7�Zj��2�|3C�e@Y�3G�4�0��"C�W�a��`��ROd��&	�%a0�XL&Gc<iz3H#GÄh������(���?Bў4��H]�ɲa6B���a�h¸aXL&	�XD�YTC
�a4aXL8a�!�VI��$8a\0ٮ�
�ON�p�8=�0��~8A������]�O����-���8h֏�(f�eh�0�896�$�,���.>'��3K#M�dp¡0�Q��VV	�LԆ��F��MǛ�<5�����jm����C�d���[���B��=����hQ��}�Mr
���I'9�E��b�UK,��4�AZ	�F�2P�U@鳚8\*���"����\d@h�:|������8��{v�"5jM���Rt&�v���pu�sgz�=��K�Pr�ޱ���!��ڧ�j��.��F�2v�ϭ��Ta<7)u[��n�u!�W3Jl��S��n	e�#eqیL�����aB���v�U�*���4M☦�%ǎ<�c�AaD��G[d�h6������+P�6Mk$���DL�r][��gn�q�u�)B�X��1��k�-�u�\�=�绫�����<V��˻����*��n���331ګjҷywy����U�i[���Λ:YgN�0�&	��@Ѡ�(|�Lל�	��#��꺮��b��vp��TxrAa�gq�����n�y��Iٞ�K����	����G
�suk���c�����b�z�Vv�wM���@&�7�=�5ٓm���'R�M�8�r70UF�9e#�	�����s�ֵ��m�"W/`܎�{Uۓn<N^.�Y��<ܦ;v�]���o��O��u{��Wcs,۫uۻ e�N����\�[����=b�����즞�Y�P��k+���v��խ�\+��:䗌7a��L�\m�y�F�֖�ղ�b�CY�;F\�8��Ϩy<�8��vܽ�	o;�@]��/TFPz�$�Iy�?~R�t�t�Ӊ���W^mUc�kK��HZ�r���f���t���{wor�!h��Y͙ܽ�[�z��l�YtHH��m�O�+#�@�F�?4|D#��{N$�������7d�{�R�zwv5s�Fx��Z_"����5RSC"���.[m��WU1�"��p�س�_���LB��O~B0[Ň�5��Ch>:�T�GԏF2���<Q��ܟ#8Q'Ş4��4�L4��,e3m���{��'�дb�Ͷ�oVk`aqyw6r=v�҆1|G���PΣuӗ8 讓�ҋ[�R�A2o���qR�<�c5-fۃ�E	{�T+Ϳ�9&FӒ2/���T�����N3H4��J���-��0v��H�3��O�c���p���,ҍ4�,�K,,��t�XT
��pTpԒI%�aqJ"4|ah�;Ѳ�$��1r�����:u�	(��۴Y�#�qZP�Ҵ"�Z�B���"G�ڍH7���e񶳩pd��&��2b>8�N�-q2F4�F��������$jJ8�W_��	l��C��L��4�ǆ?���a9Dck��h��M0�ϊ4��(�K,,��i]��/�Kcm(�F��m��x�D"��<D��U3L͇h@�A�@���DY,n�����=�x�_����q c8�j����3P3x��g�ǒ�3�!�%����3ȃ�o5��.&D�΢K�H̝8�~ �۾/��0���
4�L4���Ѡh�F
�ڦ~n�b�I�7BM�L#{{Tz{�hv�"��JRHD`�';�$�K��n�ޟ�W�g���aV�R�!O��?oZј����5e��;�zS�R����mq}����ٚ0<v���/��u�ö���(yJ�'�軫pT��(�r�v�E���w����I���1��G	>���,ПH�����$$e*G���gѸ�:��ss�rV뮼�;�g�����oH� �5 �I�J3����}g���te���C�<x�d�.��褉�XIkk����C,�(NJg@�d���PōOŢP��6i��|ig�|i��i��X�:rNd��9���_"pUY��m��	i5���eB9(�M��<JgFe�p�"�����9���/��cm��<�F��sXq|b�#Čg�A n���|.-�
+��b�$P �84�.�>*��B�rH��#Q'W�߂���%yѷ�8@ƾ ��(� ���>0��4�M,��,#��v�!�@�UP�$�I/ G.��u{K��^<3�%���pgq����G���X��@t�Bu�(��uL+j�ڴ��Uu�7�È�%#�w�����G�t�[�^2��D&3�2��q=��8��w�q��b%�)b8�|0����#�#��vPL,&�d4>�p�Y�p�
:QF�Q��a��Y�Ժ��ŵM&e�1�b{m��g�(�\�J|Z��"M+ȋ��R��1E�/o_&��h��q����~��y�U
<M\Qb����yD`��:n������[Nk"#���<�."R�pt�y�)�B:xc*��\5�GN�3�L�Q4�ȧQDA0J�Ea����x|p�M4�J4�L4�,h4��㱠�8B)u!T~t�7rKD  �֕���rjh+����q�$�Iya��}&Ӭ��j�p�t"��K9�Z��f^ڣC�
�Giƽfݺ����v(N�L��h&����E	��6�(�94]HM��j�0�I�'WD�}^��2Id�lpu|Œ�:Ng7�^=s�x�I�;*vx޷}�vI����r�N\�/9gY���1��h���:�Q�>:I�+GgN������tgB�/Ww]J-qy��V�H(��'?u#z����'�;E�/G��!>����g�,�/�q�#C���|Y�Gƚa��Ye�2�(�؆���M�Ɓ�p�{興��P2׊ќ:���2�s�tc�kU����9L��6���"JE��	�MJ<�#$�m�Ylah�\&H1���$��/��h�=n���y��I�h�(��g�>�㧎��t��CD#��GQё����:t���,�&Ν?�gD�0���xO	�O	�<'��<'��<lB�DЈ�H��B�Dѱ�D��<'���&�؛4&� ��""xO'�2|��܈�$D����ı,M�A,K4&���Q�>�A�6&�K8'�����l�:a��a�0æ�H"&�D���8"'��,K6P� �'�%	A\O���X~"���̺A�]їE�����[c*�U�6�WvU_'�SC��Ib�4�k���^18���I@@�g�ePi�g+�癯�Y��z��L������Q%�T� �Z�+J��6n��n�-���m��;P�����o��[r0��؆��>�������+jҷ{˼���ͪ����������ګj�[�˼���ͪ����������<x�K(�M0�L,��І����I$��]-�UR�4�U\�$y2������G��#�AQ(�~d8'ȤuL1�:"O�ގY6+3��h�r:�&_'��1�s��j-/�GJ>G��tae)7D����s:��xΎ|}�Nn�,eM��-F����)�T}�ȓM<|ae,��L4�
,��YR��4���"
6X�o|m��xЍf���fTA`��@Ң$��x�g�L��\+Q� ����Ky��� ��y.���5t�߇�����B�iX�����2�k������Bx�_�J㲵-f�[]�\�-�z��Dd���l1���p��q|>8�<�25����qp�2�(��<i��a��Qe�2�0X���RfښS�٪T�S>@�J�ƍ�iC#I&��A�:� �$�)i�$�I/ E����׸���wlˮ�Ԡ��.C�<մ�����k:��q{���ڣK(ܢU�4�#\%6��b�wV������X�6�.�P������^A#�x�⢏c, �t����X��`���/�x�Č�=�p� ���4p�gF���)��L���s5y|j9���0jp�Xu�S���jV��T"�.!k���=��Wm>"�Q:|t�i��i�,��Y)�-�1."s^��m��	\x��}���6�pQ6��R�|��$��j"Dw���Q)2F��tg)�m��"N��uNgϖ�9�^���|�*���[p��de��Ll������)qA �D~Q��o���O��F��r��#������|�\D�*��F���H�D����$|�4����:�Ŧ}�Z���͉�0���	�	�ƍhC�� ^�MTK��!V
� Z�Pz�I$��&��H���Ru�<�v�Ӊ%�O��n���� �G�cA�n&�m�0C"fG��qG0�e���7����ͳ�fK����'�@�J$cW���xQ��V��lgD�%�i[]c��c0h�忈ll}ߋ\:u>#�>,��ǌ>4�4�ŖX� ��q�2 �C����������P2�G��a�n�.ΌԋjX��<?#˄B:�\Ӆ�w��ӑ8�0ҏ�n�
��x1<:1�YM��d��8�kF@�U�yth��Y��pG�����e)��p8p�p�����|�G�������ג��~$����>><|x�4�O�
4h#B6�0�o��R]e0ʽ�D-�����nKcV�hʚ~>��l�I%�����⫯�jLe��	�q��]6�y��*�ͦ���n�]I�˝&VG�:�dy]��1��}�ݏ�w��U�ׅ�ݗ[�%�)�B	��y��g��ႀ��d�����A�I˵�H��P����zϛ��;����<��r�g��o�$�H@����/+L:����d�h��@q���1���fc�2@Ș�I�ui����ғ($��n"O��
 �i��>0�ƞ,�M0�L:Ye��
)-x� hlM�w�9�s��3�Zγ���'|x��G�A�>x1��� 5�b�j�ׇ�33-�9�&���ć�_HRp�|D���R�t �q^豣�$�謅�hPԹn��;�V��\,�1��;�S8�uI'�Ϙ�⃊����cp�\���ui�ĘY���i�i�K,���-`J���4/I$�� !�}� ���ב�V�2-&�����8�� ��y�E^:���|/f�N ��e���a(�����"I��6�ۜ����g͎og[ʖ��ݶ��;�C$����Ҏ����><i��0�4Å�X� �5c��9���pLQ���m�k�c�H^B�"����hm(�T;WZ4)j��ն�Im�N�Nf�K��y*���J6�,�b�Aŏ��&��#�/ߺ�������ߤP�ډ��-qXt�q�j��9��됳ˈ��i��ȣ���3���Y����Nx�����><a�:'����xN�� ��:'K(D�"l:"tЂ$4"lN��4'���؛f��4""tD�M"A6xD�����bX�,K4lM�BQ҄�$d��9�&�N'�����h�d��4a�"xL<h��a�0�8"xN��|%�f�AA��3p�7^��a�K�NԽR�2�)��K`�l�P��J�ē�l�taU�1զ�qV��iY}�F֕�W�9�:�C�d�`�
)˼
��U��ɒ��O����;�D��WvؗT��D�M�Ui�^�/�9�	�<Ъ�œ��t��B��	/%R��+~Z��Tp,9Y��]��R˚v��L�u��J��f�+��l�e����w��f�8���O�����*��\�5��ۡ�1�CN��+��$E���랷kۉ�5~.o��������]j�s[�������$q���cul�[p���^.�<�[�.�t�w�����̵]��n�yy����j�U�����3332�v���̳��8p�0L����u5����"m� I#n��f����	�j�2ö�OS�7&<8�x����C&=���A���ʛ����XV��8zz���lԊxl�m�;��U�9�ݵ�n�^9ڷn�5v�]F� �k�&����l�v���\���:�rOWT�����YWo,����\�����qE���K���X�����okX�g��\x[�㈗�w)�S�M�u��Яk;��mŶZ�1��5Wg��
�g�tq�yS���7Fۮ�(Ù^�W� ����b[��pɸ�ܑa��z��YUU�"�3�4���}��I�d��r�Ŋ�Ż��e�),_6u%=rŽh)(�WB�ʷ����ei�T�ZA��Lr!����8_Y��yԙ�M�BQ糖����qp:���<'�o����"�em����󸁑��Q#f��7��O��8R;M��Hx�Ã����Ȥ3#	�\!��j�.�j*aإ*�zx���#HM@t��ͮY��x�Śa�i�,��AF1ǭ
t����������m��5�S�WQ)w�{�8)7��Ȃ��l��(��"���T�-6
/'�&.������o[��m(a�	�"��W���1Z�� �0����#Q�&#�q|�k;�xt���ۛ�~�Ug�4w=gǌ��i�vn���E3K:Qf�x��4�M0��hC����+�/RI$��
i�m�[e�Y{�kx��6�7�$�t8�җ�A���h�~m�Ա�(�P�CGp|	>��2r9�\}����''�!e�#�R� V�E��d��Ӥ����h�P�Oz	�������3a	UJ֑��<���� àp���><i�af�i��Yc,��8��9$��(�M�om��oZ��mU��d\�ҋ�#PnE9Ё��#�1�/Bmp��R-�<��+m��3�؎�+WǞ�`x��f��k4�Z��d�fք�٘xH4�.�A��f~/��y������t���#R�&�t��YF�Y��p��hC ��M�*���ѻSZ���ٱ�5�4�u$�Ȥ��I$�^h����ю���b��u~��Q�}\���g��K�u����/h�����\���X��t�h�ZY�c�YH��y�X����G�&��/X���XD�$TJ$bx_��xqǡ���F|WG�p(��)#�&�p�K�0�8�>����q��cժ���D�A�B�iϔ!�$��lxpj��.��!EȄ��߆�Hy�G"�aϖ�y�X2�KL�xx��N�i��(�0�L(��dB�r�P�2ZIȇ�M��oF�IJT���/��W��D�G�c�H2�BL]h%v���#�<v���[�zμ�|ϛ�:_[����6��!{���z95��b�.u4x�������J��z�y��(İ���A^4��.)\!eɟYE�8p��DO	�	�G��k��||��#��ʩ����m�u�c""AߋE���d�D�/|7��:h|�ݬ����B�����kt�\�gȀ!���@��+I�2�d-J�A�9F*^G���
Fy�Q��Ά&)|cnU���H��Bd��s���T�B�K��D=J��Q�:i���(���>4,��ADy�ɂ\I� �{�m���ы�ȴ��f��aҁ�v��|�'�3��2�U��u��M�6�UP��7	��PA,��6�LCP��t�&��0����C�>M�=�q*I\�xC&bb�<��j,���gN�0}M$�O����#��t �5$7�_"t�O�<|x��4��4�
$��Y<���u�j��S\r:P;C��m��h�)�J�~F�E��l��5[�$�K��r�<Cp��E�>X�E�"������6/��M.���v
#j�Gh�����&�����j��=g��X ��W��^ui���QƇ2e�个wo�R�<�2O9��B��Lū/L��H�cU������}R<����rN�� 4��q\[O��r�PQľD&�$��p��ld�\G�lc.�Jj��1yQ���^=�f�(��k�"\��LA.\�&��&���ќߺ|�8�E*å�0�L<||Q�i�Ie��
^~�q2��1�|�[m��&���$j�-&�'�L�*��G�d�E<��6��C8R�A#<�$�cm���a).��k5�L�m�CH4���G�Ky��\��R�@�8������!�;K���s(�4�up%b�O\:������^j�#�n����TP3�9e�8p�?p�㌝�xO	�<'���"'���
!�b"'K(Ђ$4"lDN�'���؛f��4""tD���DM�"pD����ı,M��L�,�6%P�A!;"B"%�p�:'N�f�4`'�x��a�'��B�DL,�:a�a�xO4X�h�AAC�{�*�{�g�$�0�N+1:�@�̪�����u�u��y��8�Sg-�l�e�5_-��ܗ��ѦlF\��&x`�u*��u%�oU;hd4�6��.A�e�{>���bꊵ!�s*�[b�v�H(㽽�������ffffgҫ���y�Y�����t���fffff=ZUv���3zQ�<x�i��i�Ie��8��m��v�=)mq���ƽ�ŧ���y�%�����,�w���ˬ�b���is��U�ҿ���Le(BG��t�u*S}���À[
� ������3���xHz���h�jV|��p��%d�G�阈~�r�<���2���OC�n���'N�d�d�8Y�4�,�M0�K,e�M���[W6}Yۮn^���9�s��|�b�=j��%�+�ǧ�C���}-�8!�����t>�H�VZi���3K��X����<yi�ߑ��Ii�shM�Ts���n#
 <�:a#�A��/x��,������UJ�USL]H���ȸ�m��z�"�\*z<m��|�P#�o����&P�GQڲ�4����L(���>4,��E6�9�p�N�%�Bܳۦl���,�
i��!�e����M덶�o��ޒT0B�K�c��:f:ZOU�v��9s���g��"Dn�ܻ-د�}N���]��+���܀�DR?�7�%��"�&]Jp�F}�.��G�v�6�\��ͺ�ls���8,����'�Ph�Eo�]D*[�>AJ�p@�$|<r�S�8B>RRlm�O���CDMPJ��>(E�t��Ϩ(<3Ŝ<�G�$�WzuuZ���8D*h|��3��	�"�"aY�J0�,�L,�M0�K,e�M���3`|��	SbڄnrI$��+>A���m2���A�����H<�:�v5Ƴ����`�76�#��
�{��7�
:I(�`���od��||�e��~�uo8���Q�AH�z�l�G��K~oȼ�x>PA!&.N��E��x�c���\m7��d�a���YF�Y��aD�X�"�s��$M�]6�m�^�Ͷ��X�.����U1���])<���Zp��E��)|���C�7a%��1��~"bjF8�q��P %�갓�CP4HA�Y���B!qp4��'|,�=� |H�ݯ��]�?���U�b䙪<]��2@�K��7�jTt<Ag�4��Q�a��Q%�2Ȧ�������%��"""!���yx(�Lf#��di�����gy��í��qR2�]*���U�����ia��s��IKJ��(�0yt�Ͷ�yv�J�T�&JG|s�ab�����"CsC���F�x4��ǌ4�,��L(��dSv���' �Ȅ�{uQl��b�i�!q�M֜ٳKDb�m�+n@�W�i$�^�]�gf�T��R�C�
K������T�0�ER�m�Y��քgj7G!�r�3�a�4���aH��J%���*��g߉Ŕ�	�%����؉�%�ɢH�s/�[����IhŁ�ؚ��4����DO���"Q�c|r,R��Ո�������/~�%��v|ܔ�ǝ�z���x�!/-����M���l`���J01�$�f(��4�H<i�ǌ,�,��L(��dSntؙ��c|m��x���+�z�L�b ~��q���{�QDx4/��?[�X��\4�q]��A+�G���ܪ�����;�[M�qF�T�>gg}��7S;��Ϋ�_.��qϙ��^�H��2#9��2Q�#֍D�E�|6�lf�Q��4�E�x�J>0�4,��E7ڊ�)�Jҹ�1�A���+����m��ܑ9
�$�q9�E�Do�Q���Qh��-:]�gқo��y0��^�s*_?�Æ8��O�m\_{4���h���|�>�}�p�bg��$R	�����}^�16�(�*���V<I2�	9��ƌ�G�xWQJѰY��,0��0�N��u>"N��c ��m��o��(Ò�#��D��kQua�t�2G3/�]��w��zj>-t��.b ����T�C�M�p)��>9h�丮{�.~z�u�����1���M��#�\��pq��/"�����"���C�驶ܑ�R<+A�p�<p�:a�:pN��<'����xN���D�e(�b"""t�"AB&��<'�b[%�lК �"&�DD�(A	���<""t�,KblК;dM�F�#'�ܒ�Q@��BX��:lЛ0�<C�af"xN �D؈��<a�aӆC(�A�(�=򫻥{�o���,v�����q��$i�m�!Tb�����5l����DY6B�Hl�ֶ]�D�5�]�G�m��/��+K�$jAF#[�t6�Ci!fؖEX�E��:��¦a!SS�Q�X�?]���P�s��|�����ϦV��L8�:�˳Y"��rgC�l4_Q=�k���9���//Mҭ�!�<�SY���P�Ÿ��zq,�ܞ���W.�kbؘVUIQ4	���g�>��Q�-���\V��S֞�Ԉ�3
r��D�,e1�!�N[��a3N5bm�]Y�xr���GG�e�y�ݟr����US��33333�J�ۻ��fffffuiU�ww�33333:���wwn}���8p�ƚQ�a��Q�2�$��'�;����cRvEx��lg�s���J�sC�ms�^�����t�u��b��l:7��]$BH6�!ۋ/�Y�#z�>oo]G�c��93��S�'���c/ny��Y���>�u���p�١4���ʊ[�t��J�]�W|~rd��G���;'b��{�68�VN�]��	ö���TUnOi�͢��v��9M��]���sN�.��`"�i��Q�Dq �T
J��e�e��A�f�ĥ1�����ڈ�w8Od��!���;qrgn,�X�%�+���#���m�����m��ߒiE��*�WJ;����PJÙ�o�'k6��к=O+�@@=c]�/�7�Gc#�i IH#�g����_�,x���H1����D0:p)V���z>�Es�q8m�M�+�{�����C!1E�F4u2���S��R80�A`�i��|E��^�m�]��_e�b��J�^o�Z�
0��,�ŘQ�a��Q�2�$�/�ָ�D7����6�&L�Z�㹮#�WM���HN������s�pLy��M�;�Ȥy8��Qc+W��Zisa��)rc�(���Z���v����iMw�7�5+�������TZ,����$��g�>:"xᇎ��<a�<C�M�q1-~kbJ��{� ����dPA�|<o���.�;�
y����Ѩ�V�����}<Ͼ��N�;<��	��ޜG�b��r�U���Zw�2bG>l�x�����F��1P}��C�8�%�C����e"��o��W���K(���iFY�iC,��Q#�0zT7�\rA�6�h�Oc]�66��C3���S������+k�����/��X�^]�t�69�4��;A��0��>��8o#����ذ����K�-��6i0lg%�7�@Тх���g���^w��h�BŧNp���(�0�ϊe���7~Z�LH����IZ�քM4MZ�q��-L+�@�vz��f�N*�v/$�;bS#^Pڲ�0�5MUtw2�9x�'��P�SX;#��ƭ�q��U@qS6�
��g���R���JԉF�I�
G@鈱�.&0��5�qb9��^�icf�ϑ*ь%bǱ	�I�����h�[�������}���[J��m�ی��ډ��Y�U��M��C�q�9]<|Ie�x��Y�|P�,e�I�=]�r���ݮ�<�Vz��cƷ|�]�{�nk����;.ff����ش�h�X@Z��:�p�GQG�3�<�
�G��m���n��j=13ɓ#bc��r�rݻ{�����p����r.N��T�����lg�tupa�W��,��Q�a��P�,gW_|��K&�6�6��>��i8�OoHp���h���h��J�:������G�����i}:ߦ2y��26��`���y	���)i�Z+�U����{��
m�.*f��p^����oa�YA�e1{�I0�4�'�:Cǈx��S5�7	2Q7\�m�ј>"�/�k���C�D+$����@��	}��۝TiFM*h9#���h�}�B�tR�aa<d�Slt�8�Á�e7sG�AQ�l�YV�o�(;��vk:��}zUx�ɼg:�j�8ܶ|��w;m�p���{�����p�OQ�a��2�eV@���>>�>d��b��@����T�x�2'7"m����]��!bi���I�?��;��j�@��enrfw�F����5�C,�b9����Ow�#C���y)A�sy;<PB��1n���P���Uհ2Rr1����p�\G5?��8yv�Z�`�)�B�M�RqBJ8p���DVIH�<��N:��G
��"�0���W���S[>͍�<n�+@�y�>�f����=����ˊ:x<|aG�a��P�,e�I�Ɍr��L�m���j).�N���*,'ڏ��$�dk}�3b"g!�P��!��
���������oR����6�d����g~���l��#>��$dl�si�ˋ�/)�b1�J���֑�
/˃K�X���c[�Śp����:q��tO	�<'���xDD��:YB""lDDDN� ���M��gD}""tKblD�4P�$�<'
D�"lA�'�DN�%�blM�BQg��E�����B"%�:pН�&�!�af"xN ��"%��<"xN�pÆp� �M	�F��c����z�l8�ξ��q���������5|�@�+]�(۞���C,�����	*;�xs[�Si%��Ļ{�d����p4�S�\�U���&	x�^9�l�u5V��]�t�p����>�]�h4�u=�6X�u�ID��o!ck}�L�K��w/[�_�o�����1Un���33333<�U���\������V���s33333�U[����,��ƞ4ҍ0�,҆Yc,�JG:�-��h(⾞�_m{�y+D����5cm����e̘�s������:a�áS��2b3[�L����}�F<��a�}����J�|�������D��p"��l�s����*�{�y�,��Y�x�
0��0�Je���3V%[m����|���	K�#�!ƭ���^���ʛ�XI��T�����FVx�G��(���8iqB�L�hӇWk:�/g�ڦ�T�������I՚̢�@�t�usJ���$Q�� M����m8E�,醟x�
0��0��Yc,�M9E9�K��h�ɭE�c
��f)F�h������khL�k����U�,O�|��#��[��I���ߏ����n��_ۃR����X~�������X?˽��&gܱ�u�\�����7}��[ԇ{��W�թ��h'P��~���<;!��^5�p�͌c�%��J����v�8�I�#��ߐբ�<��<��C-_�)�����u#>Z�\��X�K.��r�g�m�/_Np���F�+�)��Ic�D|i��<QeY�|P�,e�I�nnB)Z| ]MbO��.D��U-慽6�F��پ�9���|	D/!�F"�.@�e�Cp�:a(��D�!��{	�$N#���I*����[W4EV�|i�H�\1B�HG�L>O��_� ������چ�z��|���6h�8'�:"xD��:p���<̢@��o���|�`��\-�C��=��4�i��<E���6�(�t<X�J��Æ|�z%˘"��L�4�HdH�m���i�x�WQ�:1�D��D�����E~�s��Ls��وh���쀓�Ye��,�M:Y���0�,�,��yL�|��
�������U`l 3�	hL�↏��P�����Iu�6�YL`M�14`�[������Ti���5�6�:�Cpz�Q�����g�-��X��Qh�GO�MW�8��jY����4�ą��b��O��Ē�C�zy�U#���k�t��<xN�'�O:C��z��N^��V�!�ZӕT90�f=56�����Qh�h*��IS6�Dh���I'ٟNϷ��gK�7�uݣZh�2g^V�D%O���"��ͩ{F̝.��S�qL��԰m��6��>΁��U��;:nE`�A�u	ܾ�v��d��I��m>�:8�"�ό1�6����X����m�))
a�BD��j�E���R�g
E�Z(��9��Ʒ��T���FV<<O7$."a��S�_��ݛz��٧[-��b1uAg�uJ�����x���<i�afa�e�ĒL�I���j�{�f#� =M��I��w0�q(ϳ����:4)f)(��K���[l�+��^~��8b�?��S�cgp�:cY����L���y�OZX��Q1GLD�Q��!\z>K������:x��YFY�|P�<I�(b6Y0l�U"��[J�E�  [����pjG���D��Q3'��Gض�aTWs�!U��8��Ÿ�h9��%�(
��3��wI�Ab/��N3�S����Cq���`R�Q�)x���<|�"&Y����<Y��ƘQ�aFP�<I�qF	��cր U�Uob�o˭qw5�~�F�&�}�8H�޶�6���v��9�˽q�4�p�F�B �ĺ�K�0����p�Y�6ˁ�cd8���k�K ��(FMv�,]�^;�Ç�������o���~M)e~Z���i�m���ߣ#�m�oN����
����n�/|q����6�i�;�����l�N�k��l�+cV�Sb=Ls&��F�k"�OS�6�Y(��d�E�ɭe�Z-5��d֚ȴkK&�Y5�Id�Ki�7E�H�--M�MdZl�Ii��M��M5�h�d�E�Z-2K"�Y�4�dZ-$k"�d֑,�h�--"Y�Y�,�F�kh�-i"ȴYi%�Z,�i"Ț,�L�ȴ�E��d֋"i#Y�"�E��$�kE�kKK&��kI�ZD�$�I-"Y-��%�F�,�I-$�yAĴ��E�KL�E�%�KH�dId�i%�L���KI-$��Ih�h��$ZD�H���"Y"Y-��ȴ�-$��ɬ�F�Id��KF��I-$��d�du�tK$��,�I6�I%�I�I2�Id�K$K$�e�%�I,�Id��I,��K$�[L��m$��%�$��%��Y-��$��I-$��$�$�I$��K$�id���$�Ig �[I,�Id�K&D��Id��I$&D��%��K$F��Y$��M6���$�I-6�I%���$�i�$�ZD��$���I,�,�$����%�,�Ih��%���ۈ��IIȲZH����,�Z$�iI--1hZi-$k$��H���$��Ih��%��"Y$ZI%��h��"i%%��:�����XЛ!cBf�d-�5��q��	��hA	�[d-��F�f���87m�B���,��ۯ.�rKVŝM��؅�!0���F!6�F!6��:��̅�!c!����!���k96�b4-�L�M�&гBb�7B̅�Bm	�mmh[#���BƄ�	�d ����	�dB2�B�Bb�LB2h ��BY�ad-�,!f�؄�#Bb�hLBAY�؋mȶE�LD"��ȶE����"ȑh���DF�s!"�"�"Ȉ�D�"E�"Ȉ�$kB�!h(֍h�Y�DE�h����D�dH�$[D�4YE�H�MB#Z",�-�E�"F�$B",�-�E�DY$[D�"E�H�h�"�"E���i�dH�H�d$kh�m-�D�""Ѣ,��"D�h�mF��E�H�"--�F��,�,��"#YD��h��"��D��"�$[D�dDY-�E�H�di,��h�m!�F�$[DE�dH�mE�z��$[D�h�m5�H������"ȑh�dH����DBȑdY�!D��E��D�m-��dDYD��E��d--��!d$Z",�H9�h��$YB#YD�DE�H�DD�DE�"�h�B��F��h��H�e��BF�D,��""�Dk""�DY�Б4HZ$Z$��BE�Sk#Y��DAdZ$YD�A"�!h�h�Z$-�FZ
5�,���sp�F�2�Ѝdk#,�dk#,���dk&�ہ�F�$Ydk �2в#Y������"B��F���dH[D���F��#-��FYC�5�Z2ѭ�h]p�h֍h�F�kCZ5��B�!d-1d֒-�Z,�!5�Y5��"�k"�Y6���-5�,�YD�E��[Q���z����5�}�sg��{����6��Q��e����{>s9�����������y�������~���~�[�=�~g�~_������/��o���_��]?ٿ���}�ۂ���}��}�_k��}����7_;~��g�^�������9����m��<��3m���o��=|���1�Ӈ�����3���������fq��翝�k~߻�߻�?ŏ���o���6}�m����ݿ���}���;?Gڟ��?�cm����������L����q�~��қ��-��3��'Z�ўv��鳙��|��}�nn���}o1���O��9x�����۾v��!�ם�?]���c1ϳ�Ff����1�雙��k6ح���o�͇Sm��6K6e6��}�[�nk��z�ι��������;��cwo�	h�l�L�(�l��2�a�(��lk�����������L�=o�x������{y��M���{�x�k�����n������:�o��4Fm����py��o������m�Cx������o���6���;c뻞��E���߾�?x���������?����߼?���ݿ[��~����r����l7�o�m���~���������y{\�C�o�6n��{cm����N��~�����㮇����:���zW������8���w0�g}�n~Z��u�[�v-�o��1��h�?���Y��wh���;72�q?��n��g<&����n?N�Ku��ۛw��=[zg�7�m������U}�+�����f�;x��~�����#_�?&�>��v��������������3��e�M�_���r���73�7��W�_�ߎM����[�7�o�o��3�;o6���>��>������m�g����l7�~��������7��~�ݟk�O�����a�_�����r�w�)'���۳���K��vk�~��?T~��M�?O��`}z폷�vt���۶빻7^������?�~F������~���s���v�'��~F�o��~ǭ�>l��,~x�<�v9�l�����7�g�Ϸ���1c���g�u�c����l����?�����c>����Ϯ����6��<^\����Ϲ�?������Y�1�F��������]��BB"�,