BZh91AY&SY��W��a߀`p���"� ����bI��           �/F"T�ڵJ��aKl�
$��UJ����0UB��)T�i��[m��e�����L�R�R��6-�RZ3X2�l�)UTY�0{7l̚Ւ�j�٤��!����-�X��A�,f�Ml�ڥ�F̫[&��4���6�Il��j�YF��U��   ���M���׀mv�2���� �\��[6�N�]��d[\g5���Ui��%�k%�#le!��$���$j���mf����KYûj�eVش@>y)D� �ak�kbغ�X���iN�mY��!�ٵ�����l�K��5I�r����n�F�GcJ�n��lk"�KY3Z�����T�oo���J omկs)A�E�i/@:t<���KjP[�{Ɣ�֔�oS��$�(e��� :A�Aꚦ�Wy�vR���y��r�Y3[35X͓m+lZ��)@����%@z/)�AR�G�<���A�:�T�뼼P:����`
ܯ<�3R�3^ox=�S=�yxP �^�����3tV�����Z�f����QC��|�]�zy�<�5�=��O)TU;y����^�5F���Cӥ)Q���z
h7���4[��z��[m4g�q��{K	J�iZ#��������i[m�խJ���m�Fzu�j�I[��@(I���z=(Y��Mpme+�k:]�x����=Î�m�(,�{�z��<��P��m�7mR�H�s� ��(L�-iZkmP)�$4l��ϥR 7��V������V�ly��SCG4�:��P�ˮox�� ��p�ҕAد{�I���t�@��U��Ji5uà��tʳR1�ն���MVVl>|�� ��� u�ϧ��t&��4���w� t����9Ӹ�B:{� ;���<G@'�ۀ���  ���TŚEMR�eil|}$����hda@h;+�浠�}�]	�����V�׹� y#  ;��C�th��Zt����m��UUV2�44��|�)J �u� �.h j�0 5{�� y�3p�Z�� V��\@:���� 9�{Ǡ(�Ox4=hov� 6�e,���U5�[Y���J� ޻���K����#]�k���9�� �g{Ύ��@ζ�� ���²�ݥ���8� �� �R�UB � � ʔ�#` i�`��ъR��      j��������m@hh    �*jR�0 	�  ��E4�T��` !�  M14$�f�RF�	��I���z�h����5?���E|����@��?�_�n��w�'��|�n�2���D�y��~@Z���D|S�X ����	�����6��TPV��$�O�� ���B*� _?���?O������lKi��%�4Ķ%�-�l`�٦�)�lb[����t�b�ؖ��%�m�l[a�6Ħ%�m�l`�ؖ��bSضĶ�m�lKf�����m�lضō�6��%�m�lK`���ClKbi�lb[ؖ���4�`SؖĶ%�-�lK`[-�Ķ%�-�l`�ؖ�����%�-�lb[��Ķ�-�lKb[ؖĶSؖ��ؖĶ�-�hm�lb[���%�-���%�4���-�[ �1�lK`[ضĶ%�-�lK`Sb[LK`��6��%�-�l�b[�Ķ%�-�l`[�ؖ���-�lK`���Ķ%�m�lK`[ؖ���ؖ������-�la��)�lKb[ض���-���K`�ضĶ%�-�l����m�lb���0-�lK`[��ؖ��%���ؚb[ؖ���-�lKcl�K`[������-�l�6Ķ�Ķ%�-�lb[
alKdbi�lKb[ؖĶ%�-�i-�l`[ؖ���-�l2��ؖĶ%�-�lKclK`[)��-�����-�lm�l`[#ؖĶl-���Q� 6�F�(� b#lm���0� 6�F��blPm���`�lAm��l@K`l@m���K`lAt�Fت[`�lm���@� [`+�6��(�`�l m�-��-�0A�*��F��Kbl@m���li���A�
��� �ؠ�4�[`�L-�����؀� [b#��A�"��F� �b#lPm���Q�(6�#Kb#lDm���� ��� �ء+lPm��Q���� �`lPm��L� 4�ؠ�b�l-��A� 6�[b���� 6�R؀�`�lm�� �V؊�[b+l@m�-�E�*�b�@�*���*�� -�-�@�� ��؈��"�؈�؀�%�����*�b�l ` [0-��lPb�lm���E�(��؁��[b[[b�lm���SLU�
4�Vب�blQm���Q��al 
b [[b�l`�lUm���LA-��1U���V��؂�)���m�i�l[`[ؖ0m�l[b�ض��:cl`��6Ķ-�m�M���t�-�[ؖı�lK`[ؖĶ%�-�lcL�%�4Ķ%�-��-�lb[m`[�Ķ�-�lKb[2�Ķ�-�lb[ؖĶi��)�lK`[���%�-�l�m�lK`[���%�-�lc�[�Ķ�-�lb��6�0m�lb[ض��`[����%�-�lb[L�1-�lb�ؖĶ%��F�-�lK`[ؖĶ�-�L�!l]1-�lb[����-�l`�ض1-�lK`�ض�-��6Ŧ%�-�lb[ؖ��m%1-�lKb[ض���l
b[ؖ��������^�� mg�J����/��+IF�K&��5���<�L��b�1f�ɉ�a٢Լ������n�,Q���m@j�*����,����̫�8D��&R5T���LLf�r�f�2$���(B�0ʉ]�"Ν#f��v[�_�gu�!�XG՜t��Hc�`Z2��D�	K��P�i��I�UI��:1n⫵5��t��El,M�bE*ýí�E�d��qCG+*h{��-7��6��˖�⌠R.�Rd2T��_�����{���45�zf��V<x�;�坙Tˀ�ٶ���cwC�`�WF'�6���BR�țgpaX�b�![Cm�Un��0��nU��S�ҩAnm7TA�W����[�e�Qc����[�7y��)jʍ�9��哭҄jl+�ao2�T�ҼN5�IVJ[�+M�T�V)\'7҅�-9GM�B/]�f�(�;��N�8�ˣ�u�aI�SEX�&k#E��з�jU��j�'B���V�i�����[��["�婧���L�کy�h抌g� �lUj�F�J�]�2�LF[���:ֲ,$�V�Զ���mIi�r�+s]cj,,����u
�]��'a����^"hɺdc��"$��B~�B\��#\Xoj�bY�.G�y�|�������M�FQ���
ɍ�"�`��2�cQڊG����f<,X�%������V]d	�)Kҡ*��4Q0:�*��F���w\��!L��PƤ!h@���PL�{
bSU�
��3�O�u%B^��:�ݤm���d�4�6h��ז�d9XE�{M-��d�x�u	[[��d,�ζ(������j��f�YS�6�U��T��~Ք�ɶ�3j����i��PRlV�rkM��ŏ^d��1ʰi�TA�u��6�ݙ�*�%$���![�Z1B�������3d��S�.޺��ضHK�Ȇr�UH�]mm-n&PШ����ʘ-��]���Q�Zt�hW-�/�b�����׸��}��D�yZ��Jj'�dI���9�d�V����YѪ�<z��mS�$u����>�=]0M��C>{���n��YZ���ie�7���ɺ��[�X]c�p^Y&;��avƫ*��b�R'&A��+32�������v���$,��z��t���o2���J�N�6�o!�ͼ�_gФE�L�`EE��=���N��Um]J��3oVxV�(5�`�lw�5���0[O��u(��F�o���Xڵ�5�۵x�
�('��FȰdŵ�����Y��*��X�7l�e�晹w�!SM=Ie��<?>���Z��՚ᴅm�OX�
�C��Ś�;H�Z�J�0�R��fűaM�0L�����&�I/[�hj�R;�B����ۍ,�4��t��kc��o-�5�h�K�/FBe�[vt݋sr�T����&���*�͕:!�%���۴��h]�k��o��qi�w3t�@��q	w�A���P�'w�����r��,F�;����gY����+BX�3E<N����#mȂ�nU)G6�5�d�e�V4�-ZwX��US"dHA����n`îQ%Vj!�XEʽo)y"����]�샮3X�cձ+��9�	��S�qf�p8���n	[�5�im�cNU\a����[-iԇ*[
�Ԕv�^�����3*�m	��r�1=P˴����Ԁ�3en�CN�TN��iwW�䧆'��L`u�*���R��ʐS�B���$l5z�n����t�͑�\��$��8�M�(�VX��;X*��7��Go�"ʬ��E�!2E1=z��C��J=RXwnʎ������H���o��h]����J�Ṻ�YTc�s*9*��0�Y�����n꟧�^7�s\2�HN�cZ�X�Q�y�֔�Z��V(�x)��$�4T�Z0n`2R�1Q�k6�1ɳ2
i�-Ĕ�,!��N�ܦ�؇uMWV����hT�鳢n��d��٘�P�ô������˰�i�8,[����=mV"��X4�$#p17e���ybӛM�CZ؁w�Ti�mY�x�ި�R�i�r�u��;��Mۃr�`BT4�f�h�ݐ��ܑ[Q�Kf-Ӳ�C*T&Q�^�Z���,B���ӊ�L�5Z��K�RPEn�����X�3�1)�T�m_�mE�����6&�i֝��{�m�y��&�˫w�J�����͎�el׫5'f�$�L�*I��C�Hm;�Iژ�Ptwdw��.�4�{śm�����,^.8���ēG5�'�7C�+M*
PSZv	^^���|k/p�7,Z��rm#HwΛ'C�5֝!������R9*�]��TPG�*/&V�!.���,7�����A��[����hmb���xV���7Zҷ��>���*��3�D�M_�QC�z���ر��w�b��Sm`2�M+R��1M��y�x�F&e��Jx�=�x�q%x��{�����!yt���-+շ�͖��kT`X���&�Ө@ݺ7lm:;�K�f�ғVC6T�Ȩ�5J��V�[�C�4�h!���w(쪴؆����V��ɛ�*xm�l��̷���E�;��j�%�@hA�#�pkP�E�Ge!y��Ű&���Q-�(K���M�Ӣ84�E��U�Z���"�Q�p+�8F�s]����yB�d�z\�ueyn�)��9P�=� �f=�i�5B�H�B,yu��0����Y����<��d��5nD�*�0�ꅅm�Ҳ2,`�ZAk7,̺ٵ�r��Z��=:tV�	)wN�c���Se3�T���6)��Z�ٵ3m˭��o5�b��6̭u�W���J�V��U����^JfX���j�8����*�X�4L�guS��k���|��ͧ�*���y����N��O�uG����$L�����Y՗62j�uz+ed/.{M�U�sw*�;ݩ��(c?;U3>�6�Spe�7	�����1�ۡU���5FF�z�]��Uk����y��̖�ȳr����U%#)��kd%f7��ԛ��6`�ّ�X�nE��tԦ���pQyl�m��`X��j�҆�:�w�
��`*2.L�1�%ߡ7�(��bhYT�ͅ��I�d��-YleF71O���M�MG3�V��*,RJƔ�U�Uz�ބ�6�-{�O;J����ۘ,�9-����58����׫j݌o-�t$-���YZ��-�\��ڶ�H�z7��N�N\�(���)b��2��p���20�YU���kW��%[�;7*�IZf�n$�Ԙ���8�Jzf�7X�+.�Qy���i�d�>K�RKr�s��t���æ9ad�l[�٘[�wẻ�X��W��V6��j��&��6Y��x��y-���9q[v3�O1��ƶ�
j�BLG �Y�b3x�E�"�-
����S�qn�C�mS�a2��B6m�{��Nȇoen�9(妊U�I2��L&T��txU��`w�/,�:2�n�$�ol,C$Ym������<���{��07Z�]�X�q�l`���b+4�ù�9*�ܗv,ӧp;����6NnB� �"��Tm����+(��>!��Y����[tvcSt0�f�KZ��F�M��TeG�Q�m�i,w�P*�g�N�&:�MfV��m-t���,�X^k�кhD�P�Ӧ��sU��/4GbM�'4�-�ӌ�l ^l-%��Y���ːeXKݥ�U#�m�f�pE��[wE�́]��՝��8r�U����k2���V��vȆ���1�����9�J+r�� �~�X��ܴ&h��f�����S���D1ۄ�z'U[-�fM�{[�F*��,e�50�����R�iӀ��q�
�d��d:���ʲ�4b�h;/A�t�e�����Hc	" �Dě�:�[t�YZ�J`��v�v�*!���DݸN�e�ȩ�0k��˄����b�,��_U��g*\H�Vwq�r6R�:t9pid����J�ܢ�T�[v햲ͤ�=�X|��zM`:k\fvmjG7tS-�e<ja��$U-�c��o^���(,l-���Ҹr��c��������,7W�5�J[��Z�e�y�����^�3����b��x�U�,�T����E�E�#�J��N"�n�9B�kUKv�@�ߪ�Vk�W��+�T�k�L��gC�1��ɓ1X$�ڥ�庰�c�wi=��V�J�n�TN�2�:���l�O��m�J��$����YI� �]��[�PU���P�v��1`t����QI?m'+M�~�H�^�%
t��!7[��l�c`{��9�7�iY�"O�7��34��[�	�W��������DMͺw{���]� �޷�m��1�M�?-�Ԗ/�֠֨�G)�*����ǯl��(����	&�٫��0����ќ=x����̹3d�ͺ.��Jō�Mʩ��2mH�U� ��zޯb�Ԣʫ�r���x23���٦�{����rn��I���)�V�ح��db�zr𽷗l\E�t"©��J����2Ua���V�(�δq��ݛ��И���j��2+�*�i+5��Xj�M1f�X���Ƒ�c������T�w����*�9RKmky���8�#��������ۂ=V���ĭ�C��լZ��m�E7tN���̨hX́!�)�k%ۨ]J�%�k1�6���V���k'����V 6� ���yÎ�[��ZX��4r�����C�uh[��1o!,��/��^�.� �1�D�C��A���ʭ�w�C�m�M�cf��ޚ���2�]nc^�2��%ڙ�N�
�dZ̦�M�Xj+V-�g����yW�d�ًE���Paf�k'mܺܫ8��a!n,{�M:���]AmYp���дb�̺4��Y�����7�/Fi�EL�;t��Ť����E�,!�������!M���3��f3,0�i��7#�~?Fv�,�yo�ap"�UX�i�'�1Mu,��OkB���(��)�,��̍���+WE���P%�Ȧ�f��RS��C*�n��U!�X׮����lHoD-�V����zt8Z���c82CnMj�6��i����fn��ʩ��w^��i�A��bF�	�"Ym���yAV"�2E�HL��Dڔ�E��(�D�ꕛ_F-�t����-6��i�m�v� pޕ��Z++%�yO.]�uFɔ�R�,:�Ȧx��i�F���j�Nh{�ň�-e�d�� V��=�Z��I�G��jC:.�1^��R�i�M��Y�FcF�����ݍ�T�h���XI�u�Fd���������dY2:)R�7�Om�H�+b8���Yb{���M��ZO�7�=:�\%�"�ܭݵW���#kK�)ەx��X�2�n��f$�>ņ�r2����]�K"�`Ջ7l:sc	;�R��N�lrB��2���KԊ01H�
'���wwcw��WYeJ���Y����@COVc�8w���v%E���x�M`�0m��J҉�M"�K#��9b�j���<��Fє���2�3��N^�MB��ٲ]:����;x���M5����mU*tt&��zR��2�`o�z�&�k��^M��8DD7I�Yl�R�V��[r�2v�k��)��S��Wy{f�$�["^&�gj�[tu歶�+�T΢�&�lJ�E/m*Ih��-���wN�e��Kv6���4��0c���F�X�O[*�9Vd.�Ǻ^�ޥu`�a�9��[KJ��k�.5�1�֚Ks�����U|͠�gVa\Cz�ei*�`��I	h���/Y�j�pS�aأ��x�B�ov�^p���1�nӧ����V�V�Q�N�Ф�t6j�vIa�u}X����D"J,�A�[�������km�C�;x�Rչlf ��y���zNZB��v&*L�Q��{(Tk'o=�s~��p��c�D�":Ә��ɇj�NwA�������Ud��&\�X"��۩��Art���mk�[�J�n��-�&�7Q�س(��Ҹ�ME�(AL��*U�Kە�+DɉK�[�tR�)$4o�7��wZ'v4�޺�E-e�5EL�V��[���n����f�]�y����kAH�*9z�^�#/m���)�6��
,�]��z�id�jH�ɲ�-T�ޝ�ܭ>�CgEM�V�R���K׵jvb��^�c���PuT�,k������w�C5�\�Ls��k.�!<�+�:qK�W�h���'Bo�=�7�,Sc���R�+v��>jJTG�K������8K[�EF7�d^nJ"f۴r�P�;q��A '$ޫ�s-U��fr	}R1�)4�IdV�%E��E�{m��ɬ��Ŵ�sD�f]	����o%J;9 ��-��{���c�)���)�-��Jr�yZ�з9�ojw��\z�I����-bsJD�c�[�7,�ܖ����[�-ґ
M��d[�yK�7�'��r�9f臄lW	֎T�L��VGxÏU�.�
�QJA���r�7-wv���U��{��6�2�D�V�F7HѬĚZ�$��V-��mw-�D���$�7��Z�+�}J�M]���]I4A�HI4R�m����T\���h��R@�F��uY�q(�r���<�qb���/uLL�R�+I��JWK�.\��x�`�Im-|�ݨ%MJF*���KuKȚ��ښ��0�#�P&�ͨ6����ԫ8����!�W�$�=�W��,S��嫊�Uj��	b�3+��H�� Kk��ݬ<��N,�kS�ϕl�צ������c��z�^���,�!C��F�g�x��8�J��T�H���Xv��}t�u�r%l��;��Ĭ_T{��ve�6�7g��]>�� M����^5Y�ee��˯�����7-q�&�Փ'�i���M�a-�T�Kim�ھ����+�Y���굯�ĕ����F�L�s̡)�#d��Z:�:��Ř�grU�j�[zC6��{��X}|�y~����ޕ���#�h>���?�I$�H&M�&�
d<�]�`�0&v��s^��yn�{�)k%�x\x�e��K����l�)���Zױ��Jܺ/���n��Ř���W�ҋ�e]B:լ�h^n ���έ|ևU�wm,�˺;��6Kf@;��Q���ǻs`�x���F��)i��1r���3���Ry@{$T�Ib�=�̻9U�*o-���	��5�a�R�RkhʛZ��ߓ��S���Ӥ6�k��y92uc$�t�c����Q��wuq]4v[�	21O���{z�J���:��q�ӹUH�dT���-�z枣����P_Wr��wݸ���e�!�.�K���Qp����V�v�棕5���`�(�i-��mAK^ʱGf�&���{�y��U8�*V�_ע�b�.�.oeI�L��Q-�2<�(�wu�kP꡸��޵%>�kŻWPtk);<�`ޚ1M��,&�4;�r��ŽBJ�{V��T���-�6�ϻ�c�On95k��7v�=Dv�^��BI�v�W[D��@@<c�l`F����n��]"Ԋ��e��\|�;�DF���q�S�C���}V=J3^�ݠD�k��͇*���^�)�*���J��j�	��
vռ�	��'�ةoGv-�2�YB�\���T�aX�&5�:mv�j`���b�GZ��ޫ���̧��[��VoVe��
X�˷[��)�%H*�fi����pZq�ݩ.I���[0�J��� %}]30��6�v����
4	�v�춣�,��o5=
�G[m��;�^\7�U��' Oc��k3tf�E�X���o+Q����������ӝ7X���n�[��{��s�*�w��M*1�}�2NK�)�����+�
�i2��s�= ����K2�N�6�<��b�$5ly�����Ε�J�]�������sf=M��]n�0ٓs�n��@����p[���6{ss�[NA�p+4�(���YJ�bpt���w��dO���NA�u��c�<۝z�AQ�c��W���ʻ�tdc�����27��:=�ҟ*�}F����M�����YB1/r
7�Ӌ>����'e�8\�O�^�{y�G��ME�I.u�xe����2�K1.D����:�����ފ�2eK[����uu��U��*�L�IԤ%�A����[l�t��ޣ[ʷ�nkz�LY�M3��2�M&`9��XwD*��V	}uf&����Hn�����-��� �Oi�d�[׆M��uƻ8�e��9Fѳ"�X����5c��nP�z��.�8�s�L��v{f��+���/�ծX�NW��wtES޳@��#ue]��fk'�z�,Sc�����*c*�Y�������J�9}�4-@�c�#w�Y���S����n�!*oD'��g)��i��V�66V�
�&8ܖ�,�������u3vf:`�k���I�����'����i1�\�ח���Nuܭ�l��h���Jtw�qP#h��&���zZ{�����v6�����%����`��&�j��6������۾�,���Z�{k��ۛGO�]�r��{O�s�B�[핕7���&[�j��u�]�}�xqq����-m��\DR5Ӷ[(fb��bw�؉v��=y[&�iI@`W���k2��޳�9�G8ˢ-�g[a[�j>���Lu�M[�|Re��{�Zw� p|�+|3e�n�D�����L�B����׻�$m�����nR�b�����z�����O����eJi��<��%N��]=ˀ�9��mq=�7F�m�g(��,��Or�>-A�W��Sp-֬%��/�㏫fǚ�Z��F���-.;�X���Q`�˄!W�r}*�Y�E�^*�ںt�RD�4y����������U�B�,���`��6e�\�X��%�p�LE.���$�'��%A�i1��eR�|���MLkl>�N3v���:�J��P�(e�ůmc)�7�p��9��"�q1�|����f=�X�m�Fqǖ2W8���k'][�z+/��Zš�����Q{��^��Ig#�!�m���1��;Lj�gR���)9-h��ia\�f;���˶�:+np��fL8�KR2�Mt.���^�X��ձ�r��xY���[�e�2���f���	"*�+om�o�z�� �5���r+
JU��n�X���4��к�&�"j��v�����n�s�}��iq�ae6�b�W^W��n�^��Q�m"�c��|�K`t3������"v\k(����pD�P��q�L
O�ڗӉSY��a�����Y���"X1��)(�Mkޠ��	v���f�U#	]��p�_j�L��",{���hL��L˒)���*��z�x��}��/x��nlTsZ�ԯ�A���P�:��i�Wr���ʛ����D��n:�)2u��n�7�Ε���NRB����w=�dSC.(s$�,�fR��t-�r�|s/Me�(mrKku�.�}V���tj�8���l����붞o׌�m8�]�a����.	6�����>�/^�ћS3{t}8��7��j�t�6���c�{,�6�FMޔ�:����S�J���I�	���j�u��=*Q-uI%j�4��=E�!m�x�M�ub�c�U�-�]8:oNW.l�X;^.'ȝ`L�z��0��~���h�}���^��(�y��h�[�m�j�Z�åY��u1�\jE�+o��tjH� �0��+6�:���	��<�h�����͓̽n'�Ֆ�igiU��6�8o�(��S6��\2y�e�+�NNٗ^�L��-j�yǔ�C]\S�"�3wv��+��B�L{J�ྐ<-brРs�� ��n^KkI�ExxQ:'Σ�2�a-�g^�XέD���u'����h��U�*�Mĕ̺d���;�Lrǟ:`�;��Rϊů�;�Set�pُuIWEjH��a��0���l��l�� �}Z%��bҝ���ِ��vV��2#ثc�jQqܭ�4�	(�N���ʴ�K����
���ֶ���bRa�2�־�I�M�̖8Jn�#�z�Y�r�ʹ������Z�g2�&�BuUѧ��3��ەӯ.TZT�<��;�Og��Rk2��LmV��[S�`�z�s��*v`��;DuI�v����eĵ���%R�.^�Wc�����בLX�"�R3!��5��jrFl�Е^���n��w�rؖS(��ن��&e�u��3L� �opn �p�Y-�̡�����ԝ�9O����|#�ځ;�����P�2���7z�5t!N��͘%��Ϭk1���u����2�W�7օ/]��]������=J�GFA��^��,o���K5��X9S�DN&}�����y*���㻮[8a抶�|L!�HtU1��Ԑ��w�R;���y�_dgt�o��f^���
��߻r*��-3&f+}G�����S,3Av�v�P�[���涞��.m��s5�^��{(�r@���L��;�Í���n����e��=[zFr�d)ˠ�Kv��	T�p��zw1r+F$�Q{�;a?�c7,u]Zɳ��U���hߙD���r��g���A�ã�/z�}^����X7�
�:�8BOT�7���s*���s9�;x�+��\q�ǹ�{wo!��(u�g����8��㭡�P�
�9�}���f���7�'��u�$��fsJ1��k���������W5�gA|Z��a������p� ��К����a�(�9i�:�0��#�B3-uGA*�ʹf��/}A�͵�ntJ,�u+	�x�7�ۦ��L%2)�9f���d�W��;O�C�s�A��\�}P�UH����V4GJ�����^�K2�G����نyy�
)�	�&��G��1�Z�b�-��oc3F�of|��#�$�M�(ޒ�̢��{Y�k��_1���
���B��>/S'-7'���)��	�Y��1V��5��D�S��Jd���h��c�O������Jv$��w�Y�&��s#<��%>�=j����,�;{u*od�@,^�A�fv��$��w,U���i��������+H�C�m<=����\�����9o7a�2ӷ�㹔f�'t���㵯��,�K;<k�\����J�ch^��-�T�yI�|1;0��ȾI�d�	����A�s6ݲ��Wf�7z�W$�e�����\)�����2
��l�
_P�2�'�(鼗�`�䰔x�r<�ӣĂx�z�R��K�A��U��vMF�Qt\\4D�_U������7WF�ΚK��U�.��
PK�����˖��̾�pj�"�] 6WuA*<���}�\���
�H�v��KT�L�y��G�c׉+�m���%�uq�vrY��=����)m}�f���,��N���3�]W�1���E%�7�gA���j�b�-�xT�{�iY_8�r��]��<��7�m��6�{o+���B"���#t;#�@���4��W�d��$�uۋ(
df�j���sp�8s�ڡ.����.GU}��A8,Yܕ�+1;�d���57��	29�:N_+�D����p!����Id�\����]+ڴ1p������fj�9S/q���H{N%}�bn��X�-��{�sN��h�)ՠZO�)T��]��؛3�Mt�7YJ�坳%��k��=���u�� �}��M�+/fu��1>��N�I�R��d�u\섙��v-��[ʅ���<�Q<�E��#�S��b��NQ�\.oD���u���jT��:�/�ȩ{�%�X�4,�NV�eb4/d�fvPƲ4R�o�8�u>���q���Y3(��l�{wm���H���МS7�w���Jee,�9���`D�a�����1��K�9j,����!�pC5� �}��.y\3mf�O0�T/0�r�Y
Ja���[Ӊ{�����0�HܡAnuM���p�:�3+kA��
)��t�(�muRN��8�V[1��J����o�-���2s�WH��ݳ[CEM��I�ΐw�Y�-���XI.k*���i	1�⍷&[�M�9�׹���W���e�+�r��n�=uV���::�m$��
�[:Ï+���h�fG�ڬ�o�M��5w�i�n;x��̬��$�h��%������%eGW3N��6̤^xu�EUv6k��T�"i���Jr
�ne��W%Fx����'�7�nR'�Zj�X��$�� Z;p���P���4�I[\j=a�fTl=�ʜS�9�pҤT��Z��D�N{:V�[�Id�Ġe�����PIuK;�X�U��GN�k[��ܧ��wV�.1���8�uGujCXq#��ӥ�[ŋ�G`"8�[(vN;��Ïfq����:E˔^*��^њ!�*�q�*ж��s�m���&5�v]'r��p�)��E���!��0�̀m�]aT�/�6;9�����07�N�������XӖF�}K�T]�p�\]M�y�^H����-�����l�[��.���R��F<��v������t����[Be}z1<�C�M�iD9�����z��ͦ:�,��n��dz�l{8�~�c�B����|�,dK����+�.K�;�6�nw|���_����d��/	��>��4��t��95�����a���e�uVt)f˙!%�w��.�v{���cc��]Y��`.��:���-��R��Jw��ڝ�f�XpT�C;�Vg�+�i��i?t����'5�kLW�L�nH����&�L�f��V8��o�l�:�����xw��C��L�sA�����缺ֹ/&���^O�&9����D�&g#�o>gA�����y��qV��7��J� �$�xv]�N[��£n͆�kw>���I"j9$��I�!*9$�����6ɫ��u�.���]�P��e�,@|Z5��*NإJ�?*����dK$�]&G�/Ye/�y��,,>��U�,@�P��,SDe�Z
x���PH�@��\(�b��dB0��h���M�$�"~f7�i6���μ�0��}l@����)���mG ��� �8�ah$�uƼݨL�?
5!D���U!xԖ���2D�jKF8����N�!M�QIy0� P�H�iI����8��������O��LH�d"�-PQ��H�#~�	��
�@�1�08ψE�XD��h~����
l�E$���ȩC=T���.	0�d"(A�� $�4E�n�~�B6�H��L����&EPI���Ң�u��[R)"1�GP���Ad�T2�`��e�P!�aD�����P��X��$�>��!����R�j������� [��M��b�I��<˺d��Q0��@�IV,�|�lOʶ\Jx=X�D�$ע�V��B�6��~r�4U(@�P�#�T#�L��0ƙ6�Ԑ�@d�Kʛtu�?%nQU3�1_���H�T�yr��ڛf�&��f2"�	C0��00�e&�����������;E�zϿ�碘����7�������?S��/��~ECDd���}/v
sV�2������Y�˺�;2u9m58���O*휘�7�f��U;�b�>�N�HD�k�*�f̧Q�s�)�A�2�'V�E�ސ������Mv��9Tۦ�s�ei/�d�K��$15���{�����5��Rm	Y��H�T�H���E�*g�m30�:;BV��t�"Ů9��w��DAݷL;Т��������Λ8�v6���ӽZ�SmD�ą��ѫۃ������5�2۲&�yؘ��t��*�m��S��D�$fq�gR�UT�sbU�p�֭�����fr=Bɋ�n���[�`p0ը�@�i齼���7^M}Q�:f�yn;#A�RT��Q�Ε7K�����n�x݋�"#z�����@�!�r���*=�qjC��O���`��u�2��H4n� �>YLWb� Ⱥ�f6��{є��õ�4&�ʙN�s�ԇ�`�}sj��&�Z��;��GP�ޒ�����셃S��Xj ��F�ߜh����KiI\M�E������y�c��G%Œi�\���I��ib��iJp���w>C�I]%�q�{���H�'����zʡY���(4����x�8��8��q��q�|q�t�8㏮8�q�qǎ8�8�8��8�6�88��8�ݻv�۷n>�㎜q�m�q��q�N8�8��q�q�q�8�8��8�n8㎜q�q��qӎ8�>��q�q�88�8��54���4��m��q��-�m/2;��pr��˕����,i���wU�*,��M��,�iL��� $������3N� ��V*뺙6��$��Ů9�W]�nǽ=����.��R�K"��-�Ɍ�
ٻvU�Bq��%̓�w��ŧp���M�\�7��k�0�c����*ݶ�Gu��
ߩ_u�u���qUG.q+v/*Q2ěj����S'M<w,K����;{{:�jW��!���t�u��D���xn���!v�A�uI�R�w�oe��-��p��f�Is�`��t�y&�=�%^
�;����{Z^9�4��8VIǝ<m[x�� ���V2d��F���̤q��� [���mT�S��ð9�p�;���Y� tiH෫�ΐ53O/��S0s#j}w]JS9*��G3��t]�Y��au�2�Q�&�&&�6�C;�9�鸢Z�YN�w��s�nߪi�ƪ��=�0�.!�%Pav
��̸hP&��]*Ө���c�Z�l�T�8*E�	ե��V��Xy4M�ZfU=xr�3��n�n�D�7q^雬���M�F�ʔ�cv��b�����3GM��;(���x�[g#�U5���xv���(h����� {K0!q*���%gs=�ں�{�t��ǃǎ8�8���8�8��q�q��q��q�m�q��q�q�qێ1�q�q�1�q�x�v�۷n�qǎ1�q�qێ4�8㏎8㍸�:q�q��q�q�n8ӎ8�8��:q�q��q��q�m�q��c�8�2�����_#p"H���n�o
��3Fk������q����xՁz``���2��;3d϶��p�� r�.x:�Ϩ���.�^g�)�͂l��Yxf�d!h���om�a�8�@ͪ�#��wKT!>��9�Jj��IU�3s]%�͚��r����uQ	�k�Qvµ��Ɩ��d̈�X���UkT��6�ZF�3n,�r��Wd�U��/%k/N��2���$&վ�[�q-X��� ۭξ��� .���XZ��O�����.Fێ����k���W��g#��LBcл��C6��>S-2TՔ/��T	gX�23�G�5�l��c�v���u�2������E̴	r����~�}FT�z�����C��ށ�sIX���`�f*��)+ ����l��n�W]�����6��-��Ǹ���p1C�����fg0�r��w����!.r��|��ۛ�#�;�[k�EJ��^r��нSzÜ����Z�ňt;��>�M�S�Q=�mvŔZ��y�"��{�� 3:4��O�oP�H[�.F������`��*wq�FB�p۽Ai?d\(J	E�Wgb�8�a�����/�^�%�����׍8�8��q�q�q��q�qێ4�8�>�㎜q�m�q��q�q�q��q��q�<x�nݻq��8�8�8ノ8�8�i�q��q�|q�q�q��8�8�8��8�8�;qƜq�q��qӎ8�}*��=���,�\J�&�v�;�m�[��n����E��� ���-���1x;�mFP�U9���b3�6�Ni��uG�\7.��c*3:�RdUX�΅�}ݒ�t��V��d��Md�gYW���1#��4���V�n-sr�J=�`pu�韕��-ƺ��
��gnh����o;Z�dX�uݞR���gU�8gtFC`����;�I�] 臰�ݡC\���R�C%#2��;:������L)�ľ�37$�a��ͤ9ua�ۄ�h&�U�������z�7�v]�őϑWmd�^ G:us�X�݂.�v��w_+�i�����4��2�]���gg6���]>C��zi��y�kuiɼ+�hn��,)��c\����rn��e$8+��)�KC��묬3.Wp}µ$$������s@�lki-b�ˌ�=��m��Q�2A��ד��+	Z��θ3!ø자�`���d�	�$�5��� X��|虃�v"0Px��s�4�v��`�s��w}�ټ����On�)�e�A��p����ڬ�T���$��tVaϨ|��5;8[���ɽ�����׊SŎ$,@;eq�g[I�x�WS�V�l	��[wZR��X�=�00H{1ʓ��x��촳6���)�~��3ٺ��m��n�<x���q�|q�q�q���q�q�88�8�8��8�8㏮8�q�q��t�8�>��Ǐ<x۷n8��8ӎ8�8���8�8���q�}q�8�:q�q��c�8�8��c�8�8��q�q�8�s���z�V�vu�C��1P��%W��o��+-�or�P��U��Z�z�ZbP&�oR1TwCq�{��ʀ �U��P[�Ū|��3QT��컏������n��}N��-+�YCK��SԑV��������2�k�y@��.m�A��JA����˫����<�WsF�lUE:��3�2�b.�N=��}�� 	����|�굚r����G5�˩�U�#�4n�@!8�%=�Ӭ|=�������cV<5�+2�\s���R�8Ԍq(i��+��D�(�L���Y���WJ��W�ng(�Xɳ���s�r�ײ=^,xWBPܚ�*̹�a��P��ɕ)������|==^��|K�ާ����Y�9aF��)����QW�9�z��-ڙ�&�K�c;�[�+*�l \Y�}L�A�!|�Ø��X̩ӀɁ�7(>ک^�ڢ�v�iڻd.X���V����v�ݷ���u��������m��>�_|�ue�����:���0����U�U���Sw���b�|���Z��[V��YF�ᜤ���Ñ�9o�\�B��,0�^ؖ����p���:;+��@	2�EI!ܮ.������G��b�O�LM��� 
0NJ��m�B�b�>��3�wuc�m�m8lVv{��w�B5���VrX�D�jB�\�4̪�}| ī ��\�gf+�����U�/�#��w:�.�A�د�A|�M	d��׫:�Px�C��Ը�>�[��^�;�X���
=�����a{]�͌|�0�NT)�S���F�d��;��������$j��j�Z_rO�}�>��sU,`
�'�Ҙ�BPY{)��u�nd�]7�r��Z�_��Ju>��$�.�����J�#�p�t;���� eܭ�P�{$38����oib�m$:�=�:M���-����VqN���CóW.vM:�R��TeSBĶ1Ww���Q�+C�b�T�-阹U����t�����z���v<��V�v=�K"l����9ͮw�����rf�	�>ĉ{�����J�s���ĝ��QO,fp�� aNi�5F3���? 6_.�F�6u���>hzV��N(a�T�&��Ύ�����Ბ4���)Z�K����ƞ�.����5�����17v��m<��4=#UiB���Js���X��b�9L5)�@��A�\,s^���UY��c�1��Kw%7J��)�΅������o_f��:�ch�N����]=y�)�tt~b�ȼ��M��,���]�s�$��}���Gspؕr�ϱ�f��l]o37�nv�u���C����'�B��XťB}��T��E�3R��w%�Ur��!��.���t�>5��.�8h��W�ϯ6kKyF���ͺ��å|D���Λ�p��o�1�����GY�&����� kŹ}J�a��:[���j��\���u��Q�$��
I�.(�ȫo:s踐,�ԣ־d���s���5��X3ӻ��g_,%a��y��|�����*�(���v��k�Eܠ =�+J�D4���:����\f��j�4i�"�z�u�����I�Z\����_u�cc�Ohr
�3��uԶ�F��)�l��E� �X�2�uy��39rz��i��&t</<���{z�3B�!vۜMO�V�6�}���βvT̉��Vpw$
�����WL�Qyu�!���u�&;��h�g"c5����j|��CW��<97o^9������Ց����V`��:�� ����B�S��˸օ{�x}Z��U�w+�����76|"�Ħޒ����N�2�ø�P��W3^��py�&�$��o��,J.���.b�9ܻ��l�O*A:X�s�m�#%��q��܇^����0T�ش�Ak��)�z�Zck���7���F9ך���=��ITx&T22LF�f�_h�Ǔmϵ��q��"�M\�X2�����U}к��z*x�(�hz�۶58h���+�W��#�a���a��4]�*Q��X5��;���5�2�_r+���L�Gn�b�L�e���B����RR�����#���կ��̥���ޗ��s�����Ø�`�:��r���͎�s#��s�wD���5d�7Wެ� [J��.�Z2�lN�K;�:���|{#��sw"��m����n�̾���:,��]��Lܙ,�t�����p�"� �+l�SDW�y���싘[}��M�9���6�u���#E����[Δ��:����6�����ø�++�e��gf*jA�}����9�����#�{/�|mF�d�ʛ�a6�.�R���`����y�D���/Y�@�Z��A �a�c�w�Z�5�@ܓH�w�ԭQ:{R"�u�K'��P圙�Ce�c5�/����;
�����j�}t5��ҽ���-���&;:�v���y��=]�vv��iΧ�!6�4�m���SI2�M���7���!Z@�;��f�A]^��񩁬-���et�Z'a3��g���(��.��j�	�@7��%�,X�Wo^�	���k�H�8�us��`��2}_$q )��ƦHd�����.��ISP�6SX�n�bY�Ϊ��
�3/�Ca#���]ہ��%W�I�<��Xt�w��e��M�s컗�>�Y��S��T��.ҝ�L���b��wRmJ���T,m�m�P�T�jYFÌ3�J���+]�pz8R�wb�(=�rc]��n��.�)J崭�i������5�8�'o��U�&�u)�*�T��ʣ�d�{"�T��d��T�n�J.|�V�"D���q�vA�:d����i��<���A�j��t���Er�6΅1o*3��7�
,P����xRUk��y�yL��8��0��lx4;f��m)ӊׯ�5Q���媨X�p\f���ʖ�� ��&�����`pWYu�*Q���'n��a|;3�ۑ�	H#x
��x�a��6������ȅ���3�^�[���!]�\�칒
��c��J�{���޾�%�$k0�.zo]���+8Qx�%p��ڲin��̧U�:�kKa﬎���H$�ۑQ7�v�V522]��L���tU˙��(���ݞ��~Je\����:].�Шɔ3�ǔ�^�h❱K���5x"(�#�I�-��r\��]OF<b���g,K����|0>��mc����{yC�;�{4��NP�˖3h^nSRc����v��ښ�"�d0w)6��y��>�%E�l[�{�k��c��޻�o��M$}U��1K��)�f9M]T.,*gfi�W��N0��IB�SWc�K� �Q��R�U�fBDt�qwK�9�.�!
��	nX�#�;dN�bNv��,�\�]���f�ΧXZ�W��2jl��WU�CF]�Go�I��^O�}Ԩ��馌�3+�̩�"������\ he+Q����S<��t��{(�[(`�j��M|����-��ٺ�i�0��yz/\H�G�Q��	����Ǩ�l�
57u�A�G�L���Z�*$�wzp�!ńA{q��՚�Y� �A��Ǹ�����n�Zӫ)k^�rc޲�sj]���Դ���C�5a��]�p��!a�14��Z���[xr(�M�firfn2o锯�e�x9բ�]v���)6���/8��7���Ԇ'޽���],��f�����iW$�)�g(s�T]�d���jU�v�t��7]�5�Cf�J���)lLlF��e.�ǈu��To�:󖼩V&�Imh;��˷O��TeΨX�3/[XNSW��&޼��wV���c��
�&�Y$h��բ�n���Yr
�İ�MK�^�� �i,��9p�l2,�W��XW�N@�m�󅧒ྸ^^Q�n���g����������@_�@�����_ԧ��c�'�p��R�?�漽UI(��5��0K�E��Q �f�d�[�����LPTq2�"2RHA�MD�1'$����2?%(�e6\e$�)ߠ/͉�HCe������Ϋ�S����b}�*t�������[�˲ w�����O�t�Q�����{�L�����g���17�p�����`��D���c�բ21AN��m�_99��G��$q���yF�Z�S�Ph&��ck�UHۖ%n�uGے�yI_8kk�^NT+��8	��s����!Y�݂�4Y�&�1Z�9�{��f��O�	wQ4_A{;���D%�è�-G}Of�XC��K�t���v�(�V��b,f�}LR���p�]TRf>����^3%��ݒ����U\Ύ��wb�Qׅ`hAͩ)ʬͭ��J7TL�{+�	�ڨ����'�+9�6{bvN�>[t�B��c��/n��Š�g�3�����0MTj���"ܵ�+�Y��X�
ʀ:*��!���3�T)�(I���,7huV�R�f�U��Lܳǥu-\F=�&)ı�C��%�
�i�7b�e����(�Kz��h6��7���	F�wa�v�e�y� ��t�
��[s��!Ҫ��P1]IU�S-/rX{Cuvt+KҬ���T8�r=�γ2+]�*F�ƭ�{��NI�m!W�`�p���A'Q��pH�P"q
&B��8�(�	!��!"~H�4A�P/EQ�$&�@�y m"��0���A��7#GͲ�e���@�R�I%Lё�al��BZ�(��H���4U���Dm8ABG�H�����$�Q�."`e0P�<**i��4�L�DL9 �D������o��1&j���E��&�=sd	$�I	uR,t����v�۷nݸ�q� B0��*20E#O�o�M�z��("K�̚J�؊��m���ݻv�۷n88�A�H�Q��ƍ`��]w��2_�� �@��T$t��v�۷nݻx���-��!aO��#&4E�U٘��\.tK�t��k�N����r�DZ]�UR��$�B��U��׮޻v�۷nݽz=S��$�	T�#R7wj��.��m���Z�N��sZ�t�B��w\�㚧�\���nUs�I�ռU�Ϊwr�ͣm�C�C��w:�lVB6��I�v�$�����wWM�h��m��\�Y%�ks��ݷwC��M��k�qi�ѷtn��Y]�~u嗎�����v�n�L����s�Y��y/3L����!ιu���U�ywW.gwN����Z����<Ѻt�ld����is�΍�S��;�wG]��$�H���L����u��h�d_��&i�M#lW�v!B,�Rh�n��_������<K�Ȉ8�6�	@T(]z���YJ9��E���E;C�eOb�svVBۦ�Ǩ�ce����ݞ�7VY��,���S� ��f�L�	p?F��PD����	�p W� �tb�"�Z�R~!!�ViY��A�s':E�Qx���d٣��}<zF�ۉCk=D��_g������:�'����^|������}�M�Dh
�Bz�zo��8�=�ꋟI6�]>�=�9�����s!��܏S��j<���r��k�{��6#�3)��X�>����3�v���d�����S�������6����9��=,�1z����[├k��7;�ד�t{,?y���MIPC�aWi�>��>��y'zy��y��ܮ'8,v/}�h=�o����q�ެ�H�r��!��~όy�������/_�x����I�:,��LZ-e`:��9��ï;�~ڻ�/�U8�>�sf��φ�߉}�>�h��,��n�t�O<�@'��#�A�o?����{vة�ב�������Yǹa3��n�ᢵ�4t��qnO�U5�e�nE\Y�CMg^��x��K�~�ݼ��g�Kl��Z֏w� �D�<$��f�^|����ݫܙ�6��>Q���:4�e͂"v�v�9e��.:�ܝzH��ێp�_US�KkrJ;~�Ί�2�#���t��㑗7�tU��9���'L$ncUܷ>Y�hW���B������ݠyvHGp�Rx�{��^�|<���9C^�����+]uxe_��<�v��ۼ)1n�O/N P�嫎�?�`���>���T;p
�
�[U�;�b�0ߪ7~��?;縦O�s���?J�}:�g������<��)�qG�y�º���&�h>~�	TwY��]L?{�3��a�>޽��|��<�%�S�!B�U�/�~�OǺ���-�����>�n�nd��z77f���<�{��g�+���X֢9�+��'3�:�e�J��ꓦ缾���g��j{�+xy�C�{�f%s֗����{>�~�����_���Oyj5��S�ڭ�#���g�`��qVH%S���'ѨH��s��(�0�Z�[n��a��rWGⲏ���>G�׮8�-�~��൥crjހ��umj�\$U�Y�R��en�S�;UB4'�^v:��ݥ�ce�wm��}�jj�p��������Z���"?u�M�Y�.�{̂��(]TM}���r9���,�WO�0�q^�EA.S�alek�ϓ�R��k/;j�ck׎�&o�轳���<�� ��=�_Ec�^M��ޓ�gw�W6�m:�w#Oi��}�C��l((=�����ҵL���nO�������࣒�,%�#�!�ߧW��/������3}2,�$B=��p˞�OQo��~�q魏������]a1��Kv��5����}t�{����TP��l������oMC�}��I�^I��~��՟�����2>�ɕ��I�v���;��~-�����֬w�>��T=^pټ����8+!�������Hש�p�^�ߊ?�jx|�ڣ���_��r9i`_w���FS�?h渽e<�u��Dn��[P�bb^T���̵�Y1W<Ρ��b(Ӷ.��"�7��ၛ`��y�������������.�$�M�tK�y���_lr*=��x0�5���4j���[�p���߷u�n�e�?��#z(�Xs�������=뿓涑�,��z���{��^�8q���8sW�yp�d,�;��;�݉�/JݞFg�w�z���UXvV}��X㙣ׂ�I�q���MU	�^��p^�v��Y����W��G�� �}x�5���=�Uȣ~���#�����P	O����s��y9g���>
{�
�`޿f�^3A��gyz��;�vMb�)k�-^��_{6E���=�o�>�&�X�'cR���K�Q�y�
�|=�|EAV>d��"�֫�%.\g}d$
��k}p����=Gx�>��99=���"�r��������&�x�=͌���>�<�^p�C��;�C�6��7��ù�\���+�Ҽ�c����c^���ʡce\��C�3;q5�n�wy�[�J�P�������/L���13��rEo�ov�f��F�U��K~��3�����$\I5���Cd���]�ʭMn�T��u�f��+y��N��s�a�����%�w��綋<�>9>�ݜ쉛��&�4��Q.�{YyVrA	'"R6��$q���xo��xaQH����($F��#ߋ��a���e��o�6���yjG��0���F\%��W�!�_����r��{Z�o�]�t*+E��g�#��TM�&k���0к]�l��y��}<���枽w�O<��g�Õ���xf�(�F}��L=�+z׬m�{�)Q�E�*f�h�A/9݄T��3gD��n�Gu;(F��[�6���u,�X:��"A�A'�Rv|��1�n�r���{}�sm��y��C�y՝S_�rٔ|�Q�W 5�3���3�����9�\r;+|��UT�����`)��)�y�;:3i�8�A=�:���1W1P"�?o����vw�>'����x�q��g�ü
C��������[^�@n�Zy�֝��{�A|�������){��k���%~�A�w�,�}ۧf���t.ckwe���v�g�wL���z:�����Y)u�%� id2�+*=�G)j2-�7t���/c��^���+���'ބ��N��|`�VI�5x���=��Ч�*ݷF�T-j�Cs[]`�gG�=��:�+	�{�c���4�3�]�q�p7���}��:�}��&��������pvS�]c��fp��g_z�t$"���zy�{�`(���`�Q�ol��K����{;�sԲ�}
��*��VG�)�8��ק�����������b$+�A��rn�7�v����#�Xuzg����C~.qk�v!4�j�|���C�{�[�?���8]o�*|,�H��4�{ݛ��5\fZ���n�*^3��Ev�����c�򭟟�b�>�y^�Q���Z���N�����~�]�|��Q��Da�w@��y����&t���̼��yp�vn�61�J/`]٠,(�L��[>���|b��0�ܶ�������e^k�l�:��ҽ��d��A�w���/���.��{�eD?�3N��qzk����R>�BǦ���l�I�!�ً�c=H)�j��K�71�3�U�p�o=,�{7���q�⹛���Qn+Z�ts�����T����,�%�dWp�UO3`B}/h�L�k��B�U�06.�j1Ώ)ϖ�vsB۬���� �>�G{�[��o�����!������Ib���[�A�y�lO�@��}7�6����os������W���a}���Qߵ?M���h8v��w5�#�����8�Sp&��p�_ ��]]��/?O���W�'g?2�'��{ޛ�Z��Q�뤎�o*�a��4��R��g��o��o�R��g�O���[>�t{�H?GRϹw����@oW���X�o��j>�hxw�Y��uxl{Y�Lo����s��\pQ��U������7fZ���/8����d��{W��6���4��H�X���u�Sn���\�����`��S+���sɚ�Ͼ.].r�;�UV+�}����~���|_>�Ϸ����L��ϗ�P�҇����<�vȬw�Sɾgٹ���lq�"���O����$wh��Bτ�D�L�wF�;����ft�E����߼�	<�nV��u��>��=*�=�J@��^B��m	�X��0�i^[�7�;l�5�bO�ؒeِ��3)Xp��@�1�U�f*�g=�.���Y᷐�:Pf�	��EB���K���w>��)�9����%�[�͝���xN\��_��W�f���lg~�q�D��\�~�`P�bQp�N;��ob{�7�gM��r�ڿnZ^������-27ҁ�7���x��u>����X>=҄�7�6�z����د}ޟuc�<N���S*���'=ۅ����s����m�3[FtE���\��W����UUxT���b�|�lT��A�^Qr4��q��|�}h�*h5p�'6��'��wi����_���[$�s���O5.nߩ��~Fc��+�����C[���O�4��Ry�.���������,�o	 ���9݆����N�C�A=�מ؜��|�{��C�v�[[Y���9=��٩/}'�>97������?>9�J�{�0�X�f벯�fhe��� �#[f��w�Q1�ï:�3�w�8�=y���*�>wc/A�;]`L巒�w- �8�k����Ҋ��Df�Q��j�R;�]g���س;�n�(�'y�������p��]'m]ޅ�w֮ S�r\�E&n�MR�a*�eH#_���uV������IH�U��}�֬ރ~ܒNK�x����� s��9����P�g��\������OvV�9�{=#�Kx������i�*��
��J�q�˪���+��q_��{T]넯8v!���}�OL�JL�Rovf�"��W3ޚl[��Kף��a�鱘{r�n\죒!�^���W9��"9/��_#��z
^�Z|=�bu��������{���$�K̘�W2��YW���L��t�rt={��L����}^�����}Қ�S��f�Xs��}���)������+;�S����U^G���H6��K�~�<�YC�.��Lۧ�A�߳����IA�;�_F����u	�{c$о40t��g 8��̕<��F��܏������T7���ޏ���{#��=�#�ڃ��oxc5s��8�[�B�!%�p^�K�}�̊GSx��E�vFJS���cF��0����ە�u��X+j!�#yF�5AD�s�F�bK���]+1��r+=]�����6)��\}K,�����Jm �BL]�{��-��ګ�ާ�>�õ�y�[׈!�y��������-K��5D��u�>�S~���0y筶t�/y?ט��_���{c���&�z0N����T ���b��g���1{�-�>�^+�=�f�����;����1���m^b�����+}�l��O_۲��3��H����zIͭ��z�X�G0�Ⱥc����to7[g��޾���~9��i�����O���X�{<�,�,�'��ҁ�I���)���5^��]7#�?Yl��s�t{��5�w��Ǚ��׾^�)����󛘽w�U|��>�kYyOks��79,2��+�=�8��(���U]}a1�'�����g���M�����so}���p�^�+Vm��D��pGhǀ����K��[�oc�cLF���S���b\�8z��3,�뺌�ײacu�
�6�+�Z�[cE�P�vuC|ڎ�Y4��r�T��úi���MzQÃ�f�{�ռ�sf����#(JP�~�Z�ʍww�e��y|�;t��U�j��؝9�B5�1�'�1ٛ��׷6��W@��@moZ�h���9M�0a�SN���y����UI�*�:����̧��fL��ob��xF��I�5��0`|hA�^�=��A��;C��Ab���\�+kA�S���uv�o����ʅ��
ai��i˨���VU�b��M�kC6�'Vuj� ���X]��vm��U���+�KqGg�Z�����x������������RT��R�۾�
������W})s�R���+n�ZΩJo�W�����p�g^�7N�,��E�v̝��6�6�$(�J�w l��t��|��^Z)?�p�˘�9]�V��K��󬠜����,V�>�Zi��a�φ��<�Adv�o�p3df��L��=���T�\�&�:ysV�޲�,�0�̏uݘL�z'6�%�,iZ�[�CR���HE�������4�䓙�kP���%sܢɠmkĠ/J�+5WM߷�ʖ_лB�5Nj
㵒��>�ŉR�/�u4Q�X�c��h��/i�:ķj��iwŕ�$��Q�Gt�C�\�NB��/)�d��BdBN,R)Q&6�{�X�ޯ6TB�gqf����ە~�;�o[�����4
�pD��t^ᣳTͥ���fDm��H��Q��R�o9BۉMY�T��կ6iw~�T����1y�%f�+״�Ҕ��d�6Uv6T����ϻiun�p�%3�����Tm�r�G[���l��&7��Ic�gL�	k��n�G�!f0�G1si���(m��<��rƌ�bY�Ds��Y-֭9�j���>Ls�{ղձN]0�6n�U0��its��u��Z{L �B�p�&u�Zۙ�0t��e�<!��]�1��{�!�hD�[ë� p>H��x�m�Y���dPV��bV�k��P`���)�T����Z��$܇%�7ͼ=���f����c�2�q�Ԕ���9(�

^�xX\V���T��P�/x�c���1X���1�i��ɓȥ��ͭ���zb�Ce��;D�ݜv�f�?)b��^՞�h@�Q��D��ٕ��&�5�,�`�0خ1��RY�G;)*�m���x]�˭�(Ӧ���ع/�!�gj5V�
.�i<[E5eϐ��嵺�=�\��b:]���.���$��{����a���#�%�ͮ��j�8����;^αL�� �e��(�	!@�j*TH����Ǐ<x��ǎ�z8a	E� A��(.����#!(I$��$#$d$�q�q�׏<x��ף�&�P�����A
�4�2��d)F�FD�8�8��Ǐ<x�7����~"!y�dR78F��ܒ�h�Nv)#	$��(	�
��-��q�q�׏<x��ׯrB I	!$�&�������n_nA��I5�}v�	�$�K��#I�4ԮX̍�u)JI����&�^�}/����$Ơ��2i��i�h�4�|��-4_J)�Q=��w]���@j��F�H}�[_nD���0D���j2F20�zW���z��2`I�ە���խEd�s��s;sn�[���ty)J����Tfy�U����o�1�F1��\߷�ٱ�)�&_m�L�ف��`[cP}�N�{o��`� O���@�'3�#���#'����}�������ܧ����yo�7hy�\5 ��,X�ߥ�i/4���k���xz/My����`9.5;$�Ϥ�N�jY�4�p�¼k>ɟs@����"w� ���.��ٶ&��Ug�!�|�)h�	]Ap+����^PV�"�(�o��/G��F|6~�G���Ţ*�o��j�]shCG�%�*tEs3̄ p���V�_�ו�˰���
ϛ���<l��At�Q���]@%���3-����}�|�Ni��п8	�dK|�+�!���*�NC� Ʉ�.�w����=��y�Tg�ES�����o��s����-ᬺ������2c�� 
�V��|��1�����*��k��0�Z��$(�����>�����[�}���������;�WDϾe��Bn+g³E���35ʽ���7]'��g4����O���<sxG��O�9������}�+��hm��E������	��w,��}����S[�"�J�,�|�x�d�����0��T규o	��xb�-��4�t�H�|w�s� �M��gf��Lj���F��seE�Ti9�,�D���3e�Oh)[\�CG6�1�4��ڜ;;.����|',>I{�T�u��<OӋʶ�Vۉ���ݙ]|���,�|��<��k�H���)��4R�[Mд���e����@<||G��6%xVy�ɽ����d��y�<�+ȁ�s!auc����ߕ����>�P%���kd�2�fjgy��Ls�>�#�������_/�Y�稐�0��3^�眰�Q�����˭��g���!����Ϧ��g��v'������_ힺ��3�5U��/�b�oޢE�gv?����e��۷�������_E�I�~����>=>��Bʠ9���t�����۶��s\�pr���������Hy�m̀�Id�cp}7B���6��c���bL�M�g�꘴��,8�x����	���6��G��|�(�~_)����z��ۨa��܋l�� qu�6.��%�F%��B ��%Ɔ����)�8�.���cH?0�L>8����.�5�J����c�ɘ�&��lOMEtpCM�{����=���>�۳~N�>}p3H�]����}>>�)x��5���/� ;�:�!ȅJ�I��J�/7i��<�`��mG����~dކ���2�Xg�ߕNC��6�v��:���Dd*E<c1�j掭��>ű���K�<�Qm�4b�}A�y��ȳ�^�u�Y�m��������P�O��s�q�8�K�bZ���N���wr�C�=��^ ��0pڔ���%��<gʙ�y�*҇��[�ӤĦkݱ��h�GJ�i:a]@hyc���i��O�i���
�Sqm��y'�b�s�#05,T�b�Nէ5A:[�˙hS�KL�}�}*\W�h+oQB��7�a�&U:Fl�OU��0#�l�MQ��{�6w��C�$(�=[�J%�|��{�߈��_F?�F�Ikk� ��5�I���`�HҢ��+)�aC�^J�USL33���=���~ֈ�]�H:�Q��7�fWl'�_��ׅt�����7�m�ق}Mu�9�N�y;��뎷^�-�W���,�K1x3=d�`i��_~��~/�%��>�۝��+�l��e��� /�:ܥɽ��)��\�a�7�O��iC_Z�p���}���@�Dڄ�m�z:����hC��YשN����-���Jmo^��|q
ϣÄ�-��P�X�>���9gs��)��*k�� =�k�M��τ��q�c� (`Q�ː1<��)��k���ac7u��vf˄i�Yx`1LBq1X{X�G�<��b[��8�Y�v�j*}>�s��T�|�5�6�b��ڏq���E��7���Q�L���Z0�V�$��\�j��M>��S<���IP�g��
���ķJ���.t��3�xE�>�w����x�H�� _���OƇȃ����n�p��C���0�����ޛ�}��\�_���L�-�!�r���Qk��@xn����}g�2����t�f���w�Q����>z]��3["v�Ữ�QUX8G:������7���d��s�:I˶�yyZ^�lj�R.�`�Ĥ�Ƭ�x�vn����I> �� *�!��k���혮�j�A�Ч(�|�	Z&0�[tv�.�m�����9��W�%Ȯ5���h����!M4B��M4
H$ r�~�==��=���� ��J� l�j32���I��-^1R��i�xg�.��~dg��B���:i�b��hl��*|�@���Z���j�K�u�����a-^(%6���(�@P�֨�8}PrV�u@g��n��y�{�_�/p(�Mw��k��w>|��i���;�FO�7��Ի#'s��ͬTP��w��goC�����sKz�=7JR=���`�6��Pa�e�es������G�>�T�biB�0ߨ�ߞHY\��E��4(SMj��Ş/:Dg{��-�5P�<��{]�����e
�-O���"ݛ �EL�>��!���e;���_w�c�3ל��������
֞�@j7���b�Mc�)��UE���;��^4}���B���<3<��邫�聓J�m�@@x`e��O�ϧ���xN�w��_�\�8T�U�����i��2d	��˓����L��5��O��_c�?1��X���޵.,�7�o����O�c�k�R��*<�u��x�c�7�zYD��xn*}��{`z��W������2�J@���2#�y6�J#�m��|7}��l̈/�n��v\���U}�r7z���TZ�A�L[3)�Y�ˡ�ϠD�V�n�X\ܪ��Q�"��\�>��䶏�nL�1���_��Mkv�e$���1�(ӗ�uvK&	cI��Gp�-�QT�]EV���Oϭ[���4{�// ���4�H-4�+"�� k�w�$#�	{�������މ~��t�����m쩖ٵ>�m��-x`cyӮ�Qt;����b����|��GG������?wP�h%�ڄ�ߐ�_�>����jd:���xf�hc[/��kI���~i��q���@�������}� A����L��ު�u��*P@�\�G�ӭ0��{q�OW?�7k�
<9��:O�K���[���A���-t��a 	����~쟯�p���p�v��u�+��(s���G�f>K� w�oF��ٵ��==�D��{i�7ۑ�hh4�y;����!�/� 7 ǹ���6�ԚǩƷ��Q8���>����`�|<o��b���0��2єMҵ4�A7j֢� m�F:�C���A&v���2�.9�����^��j��`7��� 2os�̇�������ҝ��f> ^���[�qƐ�2%������w�h���UhYa�����T�oJ1��y�!�(�ei�Y%���<=x�O�-��@�Ji�����(���4�� C�Xr��3P]����]Tӌ�:�����z�>;�y�@|9�2i�2���������!ထ����Pk�B��o�.!��=��b´z^~�^�a�_%޶��A.������6XV��)$2tԖo�M!�-���_���x7NO#�9��TN�������{49+�	Bn8g��<$b<�0i� �J���<5Ow��kR��y����y%}"�֚T��)��$�hRA@ Q�=��Y��������*���n��@W�G�u�lSx۬S"�
�*ް�Ɔ�p]O\v�n���M���Cyܠ���P�Y�G�G���Q��6�����*@Z��P����]��Ś���V5��lk?�N��[ΟL�b�h��i�d�e��c�+���<����%�8�/f������C�O��b):����[Fۦ��5�x�/{¹�)��H�'�����^�#x�0׌��@V���652�z��#"�O��!l!�"�6�+���t�<3����-�ǡ ��VW�����>7�4��,� \�ɸ�7 O����x*T[��wn���-���Ʋ@�V9��d���<�i��X�M�ю�8F7��Q����8��kS���� �[��2�5�Yt�US�2��[�u~�r���ߠg�j��/qlo	���Ս���lB�(��nj�����2�>�MR�<T�Qw��l�N��/�g���@{� cp��^ws-�j��lj�&J `72�wf��jwi�@տW���21P�z�f|7���,1�n���qs+��1]�i�Cގr��^3Ba�M�͋|������F@��&�[�[tڐ	؋lEW�c'[+���ϲǳ�XD6�9��&�Ƥl.�roS����j�W/E_B�K�CF�86�1�jc���s"��µ���Y��|JM�iU2�͋�����MX+39�V��3ع�[����s�c�����X\b�S���P�ʫ9\��9�N$��|�PA�j�.�CZ*�V��Ƞ|i� ��$�h��$II1@�U/����~w�>y����H�׀y݃?�����-@9�g>��ť�j�O%~g��Џ�!5g�@`ӭf������W�֞�Ə7��(�qC�� ���4�t�L8G�T;��4&��:�M��x�f��o���
g��J�m�v�8�<�`
��p�!�󰞘{�A�D^a��(��8�"�/r�2��Q��q\��4�r5���)��c���np��Yz�k�[Zݗ���^�U;�m�� 2]�P�[d��?���t�]�)��pu���^厽_E'<�l�Ձ�w�u�q;��`'.P�{hOý����G�����P߰~����@�8ɵ�s	�D�E���=���-x{K���^�q���
��Z�Z�P|�N�3�eے`"�n��K��1�Ӄgf:���_��Q2����?�k�%>�F�nɜɊ���C�5��M�ġ��˂�zn��0<�����gIH&��|<������,��^�1R�ި��JVG�P��%�(z�y��K�?t
��n��@�ǆL�L�ױ������6�XX�{�e���FdScP��>6�̪q��יl�͖wm�:�r�~�_h���==���2<{�I��4��Ӻg��������̵<2N�}r�5o����H������8u�ٸ�2J�ӛF�id�}�۹Z�	QS]��!�x����̝�򄆲��?ZE
i��#iD)�� ��*Db"�~g3浗�໌-���.�5�T{b����������z�e�%�[mAO�jL����e4�2�p�ϐ��(y`����Ƨ��WS���TW�_x־�Pm"4$���Zɪ��7�e����m[�9�=2l�
�2W~a	���9��r���ױ�-�ؕ�ٱ��s�S0�y��AMt9O3�q�DCv�f����:R&60�3'�X�3�teJ�d =a���M�a�[Jm����{�1����T Z%�z(v�_�eՍ�3�e��z��]-U��_���M^P�c�$Hÿ�'�rM4���4�3M	�t���j雼,��,�;��#�>���X��)r�
��b��q&}r���4��O1��Q��}�GH��j.�x�x]�<���4GߣGr��.~d�F�~W�O���J}�4q���{���IT���W�{z1z��}�3�o�u����f,�Y�x�KW�8�Ϲ�F���c�s{SIJ�[P�v�^7خ�0vaA�[��8�����]R�������f+�:&��8M��G!%D��ǃM�>=5c��ׯ�J*��r����ŭT����V����tn�9\g>�K0���Y};�����e6�E��݃ku�O��{g��Lu���Γ`ٳשni���EZ�]�3����<<=���@5X�@)M4�TI#M 5BA`�$P&|���>	]�@z� �x�4���8̱NB=6۾�u�$f^C��v/�̀.��)�0�5]f3G<�SC/k����@����>�ax�Rc�߭�����Ӎ��q6��Z�ɧ ,�l[
�o%ʼ�:m�2N	fo3A�W8�0��zg�g��d�+Z�8�kW����w:����e*m4K>��}`(J��>��e"�y� �)X�mr{Qض�q珟�_~���Co�c��5]�,f� �D����d��}�<8@�|�&����pK�6y�L�j�m�R%�Զyy��~GL���q����ր��7\�9B���Pes��4��ﶅ?�~U�M]QM�B&����>"��fONw>�=oq��)-�ᑭ��י�xηz����P�`p��,+��9�`��W�,��2��X�S���G����zOj]ٔ�mw�J�oA�2���N��}!k�{�8�E�g9�m�X�
���)�iy`��d�Q�����#�^��-���nr�J�B�v�3��X�5ʪ�"�E��u|�$z|���-����'����s'הde6�-#y�Qf��Ry�Ȳ_�~ꍗ�8�>כcP3���I��\���Us�[ʦ��۷55��ޑ�x̡Į[�H:��-߽�{� !�Ί��-�A0+����i�-��%xcR�m��VsoK����3�}�xo�9̩=���)�֐F�h)����ƚU���"��>��Vu�Jļk����樂�;�`w��Oȋ�ơ��W��AǇr�y���F�����*�FF"o��v�����.���h|n�|��ٵ?�N�[�g�E�MG�EE0��=:jz.�М��e���40t�����S7:3薼������\�����&)CA{���Xf+B������BH���렪'4�1�b�ĲeemM�钞f�S����j�ۻ�C6ޣM�_Oh%��;y�����ʐ�3�y�ME�E�]8]k�j�Se���X������\���1պ;�-���<_�)��t
n�3��8�3tE�(LM��{���Bt�GV���1��1@x���%��~��G�60�j2�":>��3E�Pf�]��+v��
Q�/��)L{c#*�s'��O���y��
&�m�p-�r݂Z��|��
;S�����������t�!������z^��Gs�c�
|v{��M���~�YԛXF���'�'�7���A�&�B��0z�Z���<я��2��I.e�&�{�����yl_����3��|���<_fFJ�M�&�K�m�����Mb�|Z�����|;%Qc����j@��pYÙ��9:�L���Cd��0��š�:[���!�L��%�ՍL�䴃��Da�fp79.��n	�]�qnemw.l-�j�P#]��ǈ��d��*c��J�y�4�A6��c�%}|ѩJrC�CY�\�X����U	��MӨ\����ٝk�)գX����c��9�$���c��ST��8�tqc���F�N�$.;x7�j�E]�Y|�a�v2���ڿZ�[��V�;��3^�+:���q.Y\_nf�����3x ���{�l�C�[n�7�)<�r��{��M��!��8Y�k���N�yfOa��}�u{^�Y�RVڮ���{;A=�J���pU�W�FҪ��[,*�m�KL�������5o*��������y���fn$�\3�Z��=�EVB7β� ��7(��{B3�c���4�׻�D�%�t��
��;K
�Rd��Ƀ}�9ǔ�p��H���!Kv�	��Tq�׽l)�;�3����,�XVA�:Â��*�9�dIr�v� ��\�	���� f]Y$e��3;i��K�r�Jж�����'������JkKX�XQiKr��{u&���ՙ5�GW�teb5O���{ʬ�+uamU�A���31�h�Z�ݱ�����0��}c��n��G�7�Yp!�l��N��V�t��"��mqxj��8Y ��g��4V���܎��|�g��Ą��5uA�V����3U�v~���;j6�����.Y��g/Fz�FU:��htQpv�@��l,O��t[��.��M��K/�8��r�'Y[�a��2TN���Gy��^kov�Dj�VUkTtm�Mr�����*,j�c*�Mr�����t�T�Jʷ�6�I_�-#����k�3GR�w|��H_)�-	m}���а.��*�H\��2J�X��������^��Cs{bKe��r�q.�2�
�v�d����uԙ�"��8&�+X�b7#W�f�� �[���.��^��>Rn�x�<�I9��9�mN�N��
Z��t� {�q{�ZGn5�C�N�qZ���K9f,[���S#Ļ�`T���̳q��|$xA��r���Mwr�.l�uR�VO0�N=["�%|sv\�p��>��V6.�k��:�j�x�P�[����ET/���{r�y�U���2֍�;[<]ǃ�ڎ�u���Yy.�{��!D��s��F�ŎktŽKf��WS(Sg�Ӥ��d
hbfR�v����w���Egm�"�p�sE+#�C%�gTl�@�Ռmq�緜�޼��Kmo�`�W�1,ɹ:��olcf�=o]8q�ˀ����x��6��P����ƚY9GYb�hS�qdُ���"�nvˮ������:�$	�a6�B`�a
E���
��USc��T$E([4�$@�e� e�L��HD��R u��,��e�8��4EH�(�b^'�䨆ݙM�$�"�(`-5N#���$�
��`ך뱴�f2'!��3����|x��׮޼x��Ǐ�z�!.�d#FLb��
H����^$*3�
��8��x��Ǐ<����w��lL�؂�DcY �NQ���0���q��x��Ǐ<x��B,F�yݞv��ѐ-6FD�"�v�ߛ�~o�;z��Ǐ=z�N�A	$F@c?.� �_;�o)z�6�%����b��y9DPT��M��$Q���Y�&��$(���PIF"�۴h�*J��9L���+"�� E��QIb���p���F7����H��1�F�㖈̱���Qi���ʹ�ŭ����Pl��U$�	��5.�v���/z:��I�;tF��/�n�<�n�x6U��sy	q�pMm����ǐ�q*�G�Q���\�y�GA��P��y2��e�"!nBb��.FJ/����� $$~4���JM4�5cM"�QP! �>���6�_W��>�52zD6`�x�G�:_��~W�*�c��ނ��"���t�v=[�y������k��"�ٝ��hs
{O3 �����.4��zN�~݂��/�Pƫ=!�ֳ�9�h��wv�h�I�64�vx
��h�`@�V�B���*ͧ$`ރnA'[�ʵ����ޜ�l9Fΰ��ޑʇ"s�@꠾a�� ���2�6z�~�S�v�]��s�>No�tom��Jk�^�Q^kI\���)�=����g���9��H�D����j�qF�����)U=epGi�� ;����|�9���l�T��RC�mQ0��`��D�D9~y�T�u��R�J����-��l��yGeW��>]6;��,�>9��o5�����t��tF�c�t�w2`g�Լ�za(��~`�W�XߍH��P�8��x��c{N���۝��u��aިI��0�*~��:F����Jr�l?hׄ��Ɏ=s�u��4��F��5[em��д�o^u�0�wc�/|�j�C3�	�1����b���JG�y�P���5\2h5J�v�3>����T'^�)������[�*���4�Q��~��=W�AӡKz�.��r7Fuڠ�]^ �˔#̗��u���zoڔ�P�v&oU�Wc6��y6>�/��h蝲>">̖su�\�'��9�}~���B�Q4Ҁ�M#Q@$I REdEd I b��o�;�j"�n������oJ�Gr��{lw�50��iF6C��Q�e;���vW��ĵR�imt���OC�S.~J=���g�?L��ܧ����
^b��?���)V��hs6��t1����,�S	ީ-���&�Ԩ�_�,q*[��>����Z������N�/��!i<&� �Ƃ��FDَ.+�o|��_����G 1 s	b�X��T��kdS-<����C	~:��F�	!�������*����5�]/�ח�K�}[N~��~�ͬ�Xc߅g�G��O�w�1�<A�*9�6��(~�'LϿ}c_�Z�o)a6���u���f�ݞ_�#5 ,0�44����'�?2�	�-w��G_�O0���昧i�ʺ���*��{]fis1~��c��<ώe���بn��wf�����Ґ�cщ��v�釬���Fֻh4��,�hbƌ['qMr�K���fD������z���<92�b^����W\�gM۩y�R�+P�2<c�?y��=�E�>l��z"��$��4�hN�+	F���L�5w�����A�Kc����u]nV��=xI��i�z�J޼ǉ�t��u���RCO�VK���ZŻ6��2 ��7Gn�:�}Il}��`_0��I�Rٚ��e���/D���)��\��y��޼�߅y�{���O֔R�iAi����i�A�  ?/�G�]R�O�����!�0"^��ˎہ-���ҏ��<WsH�&�vtU�F�դ�<H�3q�v�L;f�x���|��9���6���cx�Mc�iu�iM(l�{��)�o]
ǝ�hѻ�%o�hن�w�HY|�Z��q������C�V�u��]ƪmm�ᝉZi7����w�j!홗;5P�-L��@v�v}.fYOf�$���Űa~��{<�C�eḎ�(�`]8�~�u�+aM�@l{S�;)��i����B s������H�`��DIt��'I��9�߳�����/S=j]�	�˭a�h��ݹ��$�Bۓ9h����a�C&������s�s����Qͻh��ޗ�r]ʮ�:g�em�e*��x��x��;'�,��O 7RoG7�^�B+��/����C6�XV����j��f�@����vx��$�������#�"_m_ć��2���P�'�-��l&x���1��䣛V�P!cT����6����CzP�/-�v����4�t�7ٛ��4�f�v�r�/Tu�Å�#��uv��v|�]�<�K�����v,Zi[ܧ��S�\$���j��Y\�����즢�/.���[Fi֪�X�7�,n�S��ץr�[`͚�yY�xs�}�5U���� ��54ЍET�4	Q#M#D��3{���<��M�K�ɀ%��6}�y���z���cZI"y����ͭ~{�u����i�C.v:�S�.���~P?xc�X���ޞ�C��O��:g����:�w~u I1m$�l��t�&F���e���kK�~9��^��k�~�9�65�t��z���O<�k315Hg`]ݳY٭1���q�b\"��XW�O
��ٯP��lt�;���X�F�Lk���`͊���H,$�|����MY�������x����p��ݼ���#��.�����,,��O�\�ߠ	��+b�v���Ӑo\4�D��e��-�C��oC'��3'�L-�5];OQc���a��V"�.]�4=Mj�#���0|ܞ�\Kf�-�7�tȕ���ʹ>�6ކ����7ai¨�,�֬X�yCzD�Ƹ���x�c^�r�]c�t���%7�u��1���d���1SC#�����-M��"���������8?J���*})���+?K���7�9����g�~�}nk#Ʋ����\����v�c��yTZyc�w�^��%��,�Tl_�>�4Q�Z����Ǆ;	������P٭vgp��TO���Bt���;fD���]����=|��w�oK�G��ǵB�t���q��\���$��%/,����ЫK�B�M4PE@�4�5!�6Uz<[����O>�u�M��j��H�]b�a�D��=x�zq�������0��ߙ��3]%0�D֍�p�Wۏ�hvTD����x���H��9B<��.�\1}ZE���^|)`:`���1J�Z����W;֞��nA|N�r��:�^<�GC�^�r���!�4����A<"���; ����=V�۪�b2%=�ҟy���k�FK#�gб���ô���m��K�$�q�>�ڒ�T�10�З�Q����Z�`N���Ӭ���v}f¤R� =_�&����m��j����V9�H���T/M�Keɨ	pp���״���#se'z�Qٿ7M9|k�<�&�ܵ��Q�v��(���6�yݛ 5z4��)P�6�o�j�`8i�+2Xk�x�:�a�˩��D~Q���w��+�=O��a�U��u7֜��w�f�S�t/�����;<8��O��]'E���-A�S:z�}T�/]����@�Zq���D��$=T�w�_קN'�����dlғz�4�]�;���=;ݬ���?�Hb�z���T�Rz�qu��ޙ+o[��%L���T�İ�v��lTZ1y*���-㰼>!}�\E�����(?L]��tI�}���ո�w[�N���f+8F��|�����1�\Gij�tVJ@��>A�֑�1��J#hE��UV� �B ����LùҼ�9_Kո��w��lb��0�G�2!������WM��[��2���l�杠n @9~w��6 dUDZ��/u^�a	E4�߃y���fc(�
ٚ�N(@� 3�����Іw�*_��F��r��x�0���L�^!L���ѳ��UNt���6T�#vb�3emv�-���m�n+=�*M�;j��oG���ؗr�J1�6��h�P�m��OUO�z�j߹��$mm�ǧ�O��_�l���>;�l|�h�cK&n�^�����c��Ŗ��E�\`3as��(���)��bS�n���ȡ�.^|�le�ޮ6#���揮{5�eݵ��}���"�ra��ퟘHީ-�="gj�m�T�p��Q�:Vl�r�N��rj���_��>oS�m�[�y�dN��.(q�\��2Y��1Q���0�[�q��ЮT�2/���٤2�n����2��zn�ݘdO{��qga��VX2�UlvutL� #�oٳ��܂��s�&7ǈ&/��~-��dP�N>K�u�����*��M��eE5β�D-ƮO��O��� �C��nZ��;��L��=�U{vu�Dn��tuX�Z�jj�=��;JJwO��3}X��mw�9Հ�"���/�2�{����RH��7����)��y=�_�_ !�#PA4� SM�4ХD �$}��=�{��-E3}:�}�_"��j�hkH�ųǽ#@x��gCE{��]٘7z�?��@��śjz۝&��\��@}d�������p q�0�ޯs�l/0���[X���;�A��vg�.��b�#��,;\���A��v����ޠ�e�ŏS�K�+���Q�ߵ��}��x+]� �r"6-!�^W��#��IrWy��}~������������9G.���D4������\p��K	>E��`��i�_~�j�	3�o���|�Jy�;�?]�õn������el��N0�f�;ծo�E��Wߺ[AA�t��lh�Ԝ80ԥ�I��q�R*)�|��[�Z���3qC�M֞�Lޅ�Y�̨r��{�3�m��*J��Y� �讀���55ҀVj1���H�W�d����2�Y4��w���zTK`����WB������	?r/ʩ`	Y�r�]��v�)�f�hsK@"��d)t�\�Xk�e|fX�8�^{�s���7�6`P:Þn_.�N�X�j1-":�n?��F�c[hd0[�	A��]7��ީt����xq�?\:�*��U��>�v�RX�9q8�:�J�WS
#ʷ":�h��d�ϏJ�_$�tU��.�OMQ��	�j:�O��6gN%���l�c�yJtr�ۂ�;��;�;�N�����$�Oer5��h6�vp���Al��,nMӻ���s8>�2�ƞ��!����^��x)M4%�@	M4��!< f��f \ݩ(c���_�\[Pkjs��B%6�4^t�����L*
�E���؀������;�T"ucR�'��0��
�h�03Q�����l{gcu*��^��;I��Z��Z]��7���ѡ�7i�~Z�;<���(e9O@66���\��O0���'�Q�3�R����%ҟg�o��yl&�] ���/ܶ0B��02�\½Bk`XfY��z�K%���a���r��K�&������l��gS]^f�'���2*E�gm# 3pV��S��c��k�rS�&����U�=~b�ߕ�����aS���L�?5=�"�.�z,���nt��&�u�HQ��y��}i��0���>�W�@̎�Y�t����O۽-�נ+.��v�3"�p�o+~��)�*5�|�tNW���#Ψ�t�3=�S��!l��B{f��=D'�X��Zi&v��0	��#��~���׻������xs�-F�ۮ�2[�'װCue�[N��^F���;6)*�	j�ߖz�ޜ�/|g��"�Ia��^l��P���X;�h�M���n���ڛ�����V�����Y�'b�+��c١�����I�L$�"DU�D�ެ�B�(q�Jܮ=��x������iktuM�WHM�A	M���gޫ���>w�Axg�I��-�����_P]?i$i�F�h��h�"@`��OY^ѯ{���|w�(I^0�@�O���vE��y�g�K��̟��^WNÓ�D_=g�0��!���[5��
��&݊�]�bӞkh�*h?<�G� �+|d���L�+k�o�VЪ������k�۬⁶���5�������O�|]c������]c�u�����s���:���@;�Q��8�^����g�T��h����#T����_^(�q]*��d�sN'��}� \Q]��|�������Y"���G���Թ��ǰ<[§��>ۖl���`�Ia�o�uot�7Uj�.���i���ڤcD��r!����g�&�_=	r��*�*�KoT�
�{y�e��C[�Ѹv��3jW:��F�d{��u��v��>s�½OA�p_P�`�u��Ǹ�Gb�u/̕d�O6`K\�Ϸ�)�`���3�X�M���.�V
���Sۆ��~��L�TJ��z��
����/7�
[�/L�����m�kbzt	���qE�1�؋&"� 漬���^;c�#���~t�U8�c5��}�D�F�|z�0
�\5U�۹U�+�����z��{:�;��㎃��y%��4�H(��Պƺ$�u����_,!�oX�~Ĭwb�\��V�T��Y�ٙ����4l��\�U8�7�Ч��wY���\D4�r�&;xu�p�9�5��=����F�i�ƚ i��J�$���� ���6�d�3�߄�kI覄�6�;�d3�wi�D�uo��#>�@�����ig����w]�Gj�\O ��V��\K0�d��&9띛8mz�;Dd_=	Y�f7����t�m}a�͍(��R��\�0D}���2yg���.��� ��|�U	W����ۭ�=3f����v���q@�3�Z4�tG�uC�ͪ'n�2�<�MF�t;}�r��a~^�?`�q|}��V��6�?���<�� ʑ�-���߹�yg��
݆&r<�#0��m��ly��N�j	~����S�Q��Cl>z�����fR���7	����e�V��c�j�.��=I��U뀾��8j��P^0C&���	�+բ�R�Ͻ3�kZų��7γ�r2R�..�bˆ652�v��Sw��\����?l�3nY?�}o�s�Eaۗ6+o�ɀlq����<W-�x���g,����q-�p#9N3��f2��w�1�pj�T���A���^�D]�.��>�E3��{:��{F�f.��Y����xj.���{.��GۼV���`��z������vT�O��WݗO�B�h��f�	��v�	�)���:�5�fH%�u4s�w'��>�R����8��)�g��g�i�C98iǊ�,���� �q�+t��V[�Z�̻��`0���Ԏa��
�np�.J��y2�Iv��nY��u�n�q7�U��� �w
��CϏ+4{f�QT��
!.��o4Ճ�EF�V��6�rS�͆c�N�]���Mm4�7E,%>�'��^݃2��<Fk��S{���9|�Bg;Ţ�lL���ͮ=��ի�ǆ�w�M�=<Y�:�W}}hЦ!�au�5�UQ�O��@�,YԖU��wgI�7�����2d�O^�\ؠ��:�C7�\K{��Lڳ����gi��s#��n�yn�2�r���IJ�3_<�]L�wl[�:jr�2M�d��z�im5�vX��6h��J�����k�A�Z�]�XA�r���nV�����v��X�f��9���B9mZ2��C+��F����m�/[�ӄۮBn\��X�8�M!Ky��wis��}��I��;���sTXu[h�F�%�ꗷ�sx3�7�Gه����J�dw9��t�1�k"�L�e�X�In�8�^�]E�\�],��4/5�O`����WM�d\^ⶆ�Uy�^��!��a�ܥuF���r=C*�XU��B ��{���
��2R7��M�]��-�w�5y�;��6a��
_/��@igkr8�����K1W�rF-롃Gb;z��e��hLk�.7��N9a;�mon5�jѲ�i�k���:&�=�j���m�*��F����Z3m�:c�Y��\r���w�B��U��j�Y5*^bΆ�z�eZCqcm��GmNg][��0f_W;�|��g]#��A���f���S���o�*n��Y�uuo;!n���C/n��d�p�&Ǧ�(���S�1�F�'*F�/ ��I�v��.F��ם�P�e��Ӝ�G:��R[v��֝�wצsC����(ܶ
�^��i_h���@j9k���h�2���rW�3;wd]�Q..�����IW}-�ػ9cT8��ՠ�l�2��{����p��jX�G�Z��-���z��Mڱ"��%�:�^�<(V�*\Z%�Ѣ�͢k/�Y�f>��F;����ܤ�oz��I�f����>�|h�N���;�Lxi��(e�O�����ܡ��^�ƛne���ζ�M���㧰�3�=K%Y�M�w��Q���Vw	�̽�2D�<8�/���o9n�N���=){"ֳq�M�n-N����ϻ�I$X���da���D��
�A�o���w��ߛ��x��Ǐ�z�$�\*'r�d{�pґ��ٵ�f4��;x��׏<x��׫ءS�T|\����W��W����@n4�}qǏ�x�������w�ߨ�Y1;�r�:�_M꼴�h�k��%58㏮<x��׏<x���A;	�|�Ǝn��|�/��]�1��(�#O{s����x��o���S�ۆ���t-w�^�B\]�kEơ{*�7.T���1\�k����6.�x��J5�۞B�\���+���^/��`+�qs�;�1n7�^BFyD�	�UU
y�K�X��\����ܣr�F���J�����hw.�DuN@�5��o~���E���_K����W��]�Q��(J)#�Q�;;�����6�(�OZr��=�	&��5��r�����]�=��c���<�y���}���n�.�a~ߧ�B�~�"SMK�@TE#M5C�����.��m��ϭ�H����:b�,��4P�4�P3�^�T��L�jP��VΠP��u�7�3�ZB��f
���m�h	���<����6+6��z����m푘ϑos�ܶ��aZ@Ư2�ɫ~e'�@�&�{}-�j����{0ZT*�O"��z�̔Sfw&��/��e�%���S�^��~�q�n`���	߾p��s��@��I?=����.��������]*c�S�г���^���|ϽY�C�&>kT�Y�)���S���=-�R���@�2g/�~|�Y���-�"���9���/ba�p�����B��F�S$�Ɏ���� �������(=��L3�
7�7�o1l��j�Q����z]$��on>��"�3�҈��k��\����ՐS�yߟ��ݷk�P}�Ɖi;[2ig�T�Os���~��^-ij%�o��xע���;u3*b=��,���f��V�_�i��O5^[�-�ԋ��ݻ�v�� Kc�CŦmS�KP��>��'O~��eM8�
���ɓ�RIǕ�R;t��!��r���ʬ������I���v���k���J��V��ܤ����鎋z:�E��G���>��8`��܆S�='��K*��55ɩ�[��&{���d�~ y���F�P�"i�B�ƚTj��;b����J��Z#Z$O��q�LM@��o~CSk�T�ɬ���	iӫ��~��E�0�y�vU7n�C�ԧɠ��j��b�o�S���uB��m��/�s�����^k�g���n|�<�Q%�Ȣ�_qG��z�yzŚ�c�+��>c�	�o�j����ئ�*�P@&�,9�`73 ���򻿹�g|��?�QR.�@�Ƒo������I��WE�&��ǰV�m{�"^9�Y'��Z��k�^��>g��J3��Лj�&�_t���W8��<^"��p�dSUU�*Λ���*����-�
qQ��r�;@=Cх_u����}DP�}���K���M�b�֣N�y�%��t�̳�H�z��ƿ.I�c!_j�!>"���`�G:#�W>�v�
�+�^�����F*1��:@�ƙ�:CW�gc�CC���w�/-��g69�����Z�s/)��@mi�i�n�I�_�U���c�0;��cobW�EL�D�9�̀���!�2��^��>�z��k�#�僼�l��?�Cz�ǰo9.��U�2��/»���1���&�pI¯���5�6����+1��X���e�L�rGD����ߛ��h �i;�T˕q^K�~�f{�=+�cM�UVh���q��᫸5�UU��"�V�mP\��d�2��.���~z�JN�*��ٖ՜���XfB$Rx��mM[/VkZ�W5�p�V������jF�U��P2F�U�b�$�x+3�s���S�P&,�JDHH�A�_�▟���&�:������~��	�u>���#e��5>��pc;��5�?I=/�d�n&�r��Ƨ���F��~���0��G�_��>�������0Nw�O3+��ɤJ���8��k#�+���(�P,H&o\s�A|�^�j�v��2|���Ҧ����m�xj�����Sv���\�7_8�A'��@&]�c� X]�G��N}�15Eoʻ:�nNJ���mT��V� ?�uͰ1f}�;��b��^�Q8��B�n�;3�X񏑲�&m�,n7��$q��5l��*F�<iOc� ō<2e���6�r&�lI���xu�p��r�C�{|ȸc�%� 9pȦ�!p ��c+\�~��,u�ҭ�޺)s7$n��0m�wQ�x���jg5�l�E׾�����=5��*D��h�b~�
�u�)_O�]��x+Csk{�lu��=l'��t���ź�c:�ɶܪ�=Ne�:�y����_�~]x���֤턳�t��Frj���[ �F,�O��*���7ClI����2+ь �<U9��1ow��ދ����g7&����A�#�3v��"�A��K
j]b�`��I��Q�]��{�6��
=y�yfF����R�Ok��[�ܲra��a9#Ω��׭:��F��nt5�®�9�o7�W���G�B�@�4�4�R�Ҧ�ګ�iYV+��.�e�����ŧ� v���Ry�f��%�Dtkm�;g�m-��=�5�?`�pS�����E�c٦vg�Cq�o֠KH�ol�=�Bd�QK#�s>X�-�|�C6�bf��g�_6t;��]�h,k/�ැ���ʽO�L����:�+�Ӭ���z�')'g♤�=E����g�~j�^���"l�q��W~\k�����q����E��,���C�q��?�h)w燼��3����K�-���t����5˫~��$���(�3׽71���8,�d.�AwIǲ���`^z�T�	������[�|��ٿv-�D7<���#�ѹm!�%KQvbدg�3��5���1�a��5�r�|���m�w?iP�y��b�T��b[�P��,&}���ɢU��A׵�1A��e+��įL:�j�Ȯ�gu�gR�wB��V���"�r:��B��sր1NX��(A�dKfE,��ɣKD��w\gČ�^�7�2R*�.�ZK�<�z`��U�0𺫂�R�hȑa��7�fmwd�D3+���&:Kxֆ��m��(\Wy�>!�X9��Z��1Yz� }�ے�Rr�ptn�;9�	��I]6T��[��	���n9�PR�p���S�~6k�Gg��s������!��H�KP�JSM%0Y	 ��Lϝ�|���|��N]��~�D3�\MtK��=u���g����j	���S=vo��j{7buZ�',u��b��[�6���y�be#���~����]�=3k`,�Ɩ����Z�.�bӱ�$lBO��]�x��]b��׷�B�,����;�f;�ߚ�EŚzv	uRtn��S7������f������rzb�s���>�����れj��Aw��W6���^=���ç~h������hL��2��9�`�_���۪:|�d�L�n�����ǧ�h|��f>t�J_�ż��
����ה��c���j���K�m�J��s�cwq�7}k����:k�ԘhY#凚Z�6�|��Oڼ�������y��s&{�]�Ye]"\ �K��$���@�*y����];W��WFƆ
�	~_=������0�9>ԡ�\�aIoHYܬn c����&F�1lX�Ӡ/Cg�k1Q���DbW_|3���̏�-?}B]#�;����8��-t3���&�}!�˗�O�E����r��LdZ����_������%@������r^]�ԉ�N�U&����e۶�g�bw���I2�ip�}��e,��׭M�`lb�(i۸:>�N�w|�����պf�I��:���V����H  �y �hi�)`H;��U�s����>�o�ʢ<�����̢_���!��w1d��QgÐF6��.�wk�mBhtvV/������O�qx`�~�Y6��\l8�6>�c̝�q�����ʧ�d�"X�j:S%��]������PQ��`슁bj,�^8�ϧ^ �
��9Y{zu��v� nz�ήy�\����z4F�G=�������)}�ߓ�j�ó��-��w\�1)�g�p��y��BeG��c�Ս>�"��)�<��,J~}U͢vl�8��!,�W����_�X/_�����v��:�S���U]xQ�Cȷf�磊e����L�����7˗���t��1���[4�����Be�8�1Obָ�m*���b��M7
͌I�X~�s�U�@����Nn�M���!��v��������
�DOL!L&�]�,؝,=\��kZ��7�v�g!���kY�8aޝk*<]�6����iS����,��MZ�橻�[��)<c��J��*��=��G����K�\���둞��D>^+��ƷޖEB0D.�^�Ou����	��f�|��б�v`F��D��[�j(ES�}:���KWoZ2u���:�T���2���}���pn#Q]#�����FN�tZ�`��6l��K�X,��N��\��E5�%c�glzF��Z�8$���)���	����:ZH�IM4�MP�X�$@O ��$����>f�"�������g�F�:_��#�m�
�k��	����%�������Rp�OV換4z��,�e��[B�YM�^zu���}�0���7-�T^�!���K[$e��be�3����-Og��Ȏ6���|�>9.�/)��^[Y�[�����:�5���Odxi�����H�~��9���BQZ"a�9<76�Ҟ�ޝ��6�޺��ψu���_3ٞ/zeF�W��Z�|��*���!��]ٶפ���0 '���|c�\�Ͼ�� ck6�bK�U�p���vx�@���
i=QA��I��l~A�� 1��΀�NQ���ݨ�W���א��C,4�,y�p�zE�C��q�����.��С�5D�g���*1�V�4x88�iֳ e�6�Wm�f�/��]2�.�ح�����*ɋ3ohx��5i��=ѹ���S��qQo���ꂝ�w�����G�T�2}b[+UӰ��."Oj��e��RiK�s���H����l���P#�l,���64�Ĳ`������ߖ8�|����/�Ƌa�TM�^خ,��lDM9�[t!h��oJʕ�V�k�/֧���ȕy��I� u,��ES7L}�*�4^���� �zB�=���{[ƒmQ�@�����y_=ƇW���&V��NA��Z�=��~���0#M	#L��5P�f�0���=�[S.�C�1�3�����Ĭ���'�L1�u��i���׮����oE��R��SYWė�
�M���&�Xp~�c2�]O���*6m�����)F0;�1���Z��X��"��ap���:�t��-�k�����������g��3_��_��'5�p����b��7�:-S1�!��e�^�J�b)>�x���F�l�o�/��0!��E��=����ƾ��{�=N���<74��j�7���z�k���]���BG,Pc.���F�Q�o7F�k�4'���&,ǽ���ֆ?���<�5�)�X��G��sq�(K2%��9b��`����Iz~�=�}5 �k����Hh_������A�\k�&��.�(����e��r�FX�4OƔ_�NM缿{>�O�J/X���%k Γ��z���q��k�y� �f�3dTT���5�z5MѮqH41��zc�A��ަk�ă�'(�V$~�u�~�����Qt�^�?q��ζX7�С�����A��p^D���>46��N�0vBDh3P]<\��h<��V-i�Ն��b��g ��F,��T�0����R/�j���9k��{ךY�ka�O�e��6�i����|o�ܔ��8���5C b�h�GhGWI��]��ֹX� �S
e����W���y�>�~�L�4RS5P���<��ZM4B��H~�:�fƜ��g=�clq~.�j�+���M�C�<��L9�/#�����Zhs�R"D�L&&,�(0/���	A��3���\O��M������[�k�s<oK�R�lȞ�t��+�*2 ̒�؞�r���+�І��	A�9塐�U�Vc��BZ�c�C�Ʊ�w�N���|���U��~��OM^iJ-�"��iYn(�.��'L�����4á�ʹ]
��/�-�-�x~�v�g{{����憚PS��-\�kٶ5�]T/��J�1v|ie��u�Z�+�����^�~��|�%+DW��;�-�j-�����|������-��L�&p��P3`�l������#�U{"�>dd�[�0��zh�2KA��H%�KWKL���2i�O��}-�xlL�~��_��{��Wv2�S�F�R��=ttZ��n�US���y��<�64Ð�^���&C��)�ގwf�-%��\�5��3m�����Pd�ՍK��p�.C��I �z��Z�����"E�������hf�����[����33
Y�y}ՙ�\��l���9J����h���v����b�����u-iXߵ9�/-7ܷ%ZLB�X�l���WC�Y��X�����C����+�T��������'���x�;������=V8������cg����k9��%lSkQ}w�-�(����k��]�
~��l���@�\�M$y����qQ.ٱi� w8�Ia -j�j�rw���ǁE��ʘ�]�[Q�M�O��l;�A=�w���4�����b�%��%�*��J�ͭ��n;ށ1��kw�g>�?������b�� a�^�Z��x?����P����qX�&2&�P�6" L��$WQD1ؾh�kﾛ�\G�K
��{0��fY�ɍ� F�Rw>�e�ߞ���z�����4��3�����|i}Y�;"!F�<�v��v������ڰIx���nӚֲ�KVk@+�6��]�Q*�$O�(����o�1B��Ñ��sK�6>�*��:S\=u��:��v��2��Ũd�MÇ�MӰ��v�IÐ�<����᣿N�M��O��{�4Sl�O���<d&\jq��l���.�_&�6P�㐕��h�I�D��n����l��[�p+eex��9�jʆ/>�ɝ��U�:���ؼ��0��x9���<<}7�T3��_l���r����;�v�B���2H�C��;1�u��x"�#V ���;z��X�޵�rӍ]l�=}ɳ�\{��N���5+��6��A���<+%��ћ}j9r���Xk�� �.����ܖ�<�^=�,�c蔭���Fo�$М4�����f_�������YCK�F,�����JyH�)�7\��l�&�~�Q8����Jx�x��]��	�t���=����,2�x���bȊ��,,"Z��a8.�e��}2
�,�LX%r���]��1��C���%�z���Ү5���8x�@��-�t�pւ7WHQ�wd*>ǌҪ�b]<r�^�.aW ���5�*C�����{���ؽ핵�
�m���G47��L=h��W�����©�[[-�dڪNe��X��r�1P�tz���a6���}��8=�s�C6��ԩ���U����gD��;��p�xb[���Mxv��]a.sHK�i�>�,�����;õ� O�����RU�Y�1
#s!џ�`��*�fP}A,����}r�7�:V��zFGZ��0川���U��5,�T՛�\ 6�����6��&�g�f�7d�I�v^��\��m���c��Un�����4s���1X혨��{���5�zb�8~���|�n���[2�-��$+ġ
h8��K �c	�Va�/:Ě��t�[6�G)�̬�!��e<�F�۶ek�U	G-�.M�}�T�&��2n;�֨h��9N�0�0!�'P���� �������z��9'�AD01�21��t��2�e�pn�[n���׎r�V�eDV[��w�Y�3�-9}Ju��i9p�>q��QpNǎ�/�i���<��H�{A��V[��v�*�Wx2i�3���_4��ZѮ\��D����Kr1��v;ۚR�J'�L�T�ruc�I�d㲒��x�����о!ۢ�>w�U9�x��Ւ��m�y��CA�����}�wns�ocW��Km�F�7;z�WT�>36Z��_� .�~�E���L�n�)���uݝ���|����#��*��H��n�__�vowX.T]ٗ�u2�m ��	eIt0�k�3#R����觼�m`{C8&+������nu}�q�Z��B��b��(�j��u����v%.�ӷd��(K�R���*�V7u�=��ژ�e2_-w��J�Ղ ����:����oC�r��O��=}8��E�Y�}�X�dn�ĉzK�z�遦y��=X�n����'��)&q�#�<���$�m��uvZ��?7U<�Я��Ր[�������U�Q����z^؋�����0�3ye�D3��س�-����Gg:�k�ph����U��쓹�ws��A0�F���E�j�md�	A��L��D�JA�!m�J�4ځ�SM�cByB�m��/H#%�JjZ�B`�C�FK��WH9��2ـ��R(�p��d �~,&'������㘣o��H���w�=��z�OM>wםp�wm��ݼ�}}v�ǎ߯<x��פ� �;/'|�v�h�{�[;��6� HT**��Ap�T�i�}v�ǎ޼x��ǯ^���$�ơUSE$��>#!I bC��=sDn�ۘ��Νܮݿw���v�ǎ޼x��ǯ^�Hw�)*�o�������������X�Rʢ�Gؚ�G���Ǐ<x��Ǐ=z�yN�(�'cRJ�'�������>{���h��x����P>����{��/������[���{�=m�h�w%t9�w5����ד�\�u�x���������	6>�����`��^6���<��x������޼��k�@ԩ��UJu����N,j%�
%rv�\"��stD��=n`��{�_@׊�79�������sW~\���~;מ�wyD�r?pI��Mn�p|�0�\���n�b�\}��f��v���.OD�n+M�F�덞�o-<��&�|V����P�T`^�����	&�!�@�
i$1ȉ ؂H�$V�J�:Ō�1�=+�׻��e��E�L"�n����L4�����?*��.��u��S��)�M��)!���b`7^ʦ��z����>�2�|���ͣ���֒L ��T/�����aOϾ��9���岯t��텍z������>�S�Xf����_b�C����l���u���EڻKy5FenJ-�d�n�s�T��z���q�m��e>(O�E��+k�������꯻���i�VF���0�ܡ�z-�5��!<�;�_�,e�|����lz�`����'�d3����-C8��v
#���'Ϸ�!�`���`њ`k��Q�7-�S4�ŦC3��´3�|�x#��,��:��ɗ��a�O9�+>�_N�8�.�~w�1MgS2g����.�ZA;���|�Ё����76�o_(�1c��?Q�d�3i'_����o��Lu~~�A{�  ��E�7�D�d���D>#�(��1��8�F��혣UY)����@�d��;�*���?K��^���ԑ��x�0���EF�;�(Ʀ��!�K�[�2�E�^E�7߯+�ˊ3ܪ������x�#���\�d��շ�ɜ'���ٿ�=ƴ�y1<���y��K6;[���哆:���=��!̐h���e�U���g�;�g&Yy�������  ���Y�,Ɛ*���5�W��b�ߝbΣ��r�i�&`�'}g��Z'�*�E���z�P�&5�Y���f�`�n�v޷R; Ƚ0�*�A�ޅ�����4ᙦ�s��b�i�(���
i����MG�j)��|�:�b2���},�Au�0��q"�S&E1��n�q���#a�|���P����y��x
���|d�q,�T��)4�E�J��$^Z���+:@�xn`ǣ�Ŵ�\%�@k�ȒX�ׯX�+�V'�Ce�a,��_]��17�>�]� �QugdSe�f�6x,�`*��v4{9��ll��[گ����9�&CC�Ͳ��a���2�Dp�l5���&\0��t��m��V�Z��'%��z���aQ������ǵD�i����Y�a��;�y��Q�1�4�>��F�tnE���<#�Ŗ��8Me"7_��v���;�c�s��ᠵü9h}.�/����x�y.�׌Z���T��?{K�매����UB[�r��r�dO�2b�$O<ف-\�Ϣ��2k<�Dv�(�ݶ�S����o����΄�R9��*5/�z�53|��N3���za��9pGw�O
�B�ѝ�e�fYC+Y�6H/������E+�O��\�}�B!�N7Û����t��К���}|��'��
�wAi�"� /���l��q��V���U���c�}����k����%�v���f���D(�z����ݿ4t���w�\v��o6ؒx��8�)��\K�.c��9�\q��r��8;c숌f���\m�#�ӶL��En���
h��k}����\e��a���b��	$ޙިk��kQ$��ϥݥ�HW���m��+�:Pp����g����s�m�o^���e�Q"#��ٵHx���1���Yjh�������\��(�U/��>�i�s.�.]4y�0�5�^K{� J��M	ȋ���Kva�{��w3���0ś</ҫ��X{��0?1EB��܅y?3��Y�����g�����m�zc�0��G�LH���c����ljz�o  ��wlY�`X��m#☲�β��1[�V�����!�5�������Ƈ퍵��j?t�H+ �S���Yi� �SqZw�����~N������ ��o�����/�ÿ����j��9�m�{k�v�d���&�>�ӽSB(c�w�7���b��'
D����^�����-`T�w�f	շ���cZ���{"9��3���eU?"�.��s�WvkKH�zK�Ҹv �j�˹��GO���t����w����NIW����[U��\'�~4�db�uy�~J򼑻�mu*�î�o�3�N��1��};j�gd��c`�ɹ+e�dZ��RA��}��{�����u��S����?e����Qe��6j� ��=>(�K�f������VT���b�=�T̪:�qT޳dm-^ o�Bi�"�����`��LC?��f�Pu׬��@\ �SJ���-������ T؁ja=�0�j��3���1!���?��nlc�K���8X:���|X��j˖
�4�OY�<lW�N����݋��wG��l}_j��yCBk�aU�9xM��\&�|h��Sc��h5���5j�rY��a y���U�,$e�j"���'����jO�$�Xx���źmM0��n���>�
T*� $�vw���=�LSϋ�Z�6�]�zCנ�
�&ojK�[���y����Υ��O4�`1C9�s�p.��M� G�B��D%�:���T��b�i�Z;��]���(E��<>����2OR��!�c��ޟ�_�>*�"~c�ʥ'W!+����xYP4��9��a��~�k�)h�ZD�?]bIg��S�����Mv��l�3O��nʜkة�Ҋ���������L���C���R��7ٍᝆ�_|/�״��ojwk)��)/_a�K���Еx�n�m����G>ɂ:o���DG]9��$W˲�iY�^i��Y�`�T!�d]!�:Z�T���ӶoG87��dCj��t%��]]{yE��f��}VV�����;���L����()Uxye�Th�kE�_ʚc�%�!U����߾7�-
�0�E��,i �|o�a7.h�`��i�=t��˼6K\s	�Q�X Bjϧ_ �f[3儞�h�ʃK޴8�xv��|�����.OKh)���[#�G�s�a_+$��'X30�o5+N��iЗ����umI��F��D�2*���k׎���H�s��zw�WwzՈ蓔�v�����q��<3ω$�F�|�e�q���*��ؼ���Jѭa�n��lZ�ݡ���,��ezϞ��� 9ٱ�;�<��S�z+޷[}��\�Vg�N��E�"N�i��
��h.��E�@�y�+�����[y�&Ʀ���9"m)�P��U.�]Wvt��lG��>0^�R[o�ǩ��[,K�fɿE��,���R�`�6��M�N5��H*�e�J�h#^��3@�=�)B�/~"��Q�G3�k�T+�iTh=�?���O�
뵱8sW�[ͯ໯77�t��
M�{>8ݐ_*٧���ЊUH��9�ߌN����n}/�-�>�U1p|VJ��͏D��e~�!�o��݀]Sv�)l����QEF6��`@�X�#,~E��!����J�-Qb�t+���V����Y��3��cbɭ!ӯ@@漕kN)��N㬓�����a��|��!�w�pgc��rTU:��y��k�ߦ��7'9�����.�ƻ�,�v��q���oS��.�����Jܺ��	o���>>>>>>38�]Z>K�h-o����|�+�:c�`J(f}��cZ���ԕ��h����,�z9�٩�*�6�Z`'�g0t�laao@����|����>T�6��S��uی�6��U�����6�o/k"vC�	5�fZ�����<���,�C�1^f��/C,��a�̸��:�`ͻ6v�����ss6>���'�)��?�X)��#��8N0�6�� X9�D��R���W-� �P���@����O\��73�fHMZZ1\�9��r�2�Uq=�C>������,��s�)0���fO�@��h�R�i]2&|⚇��jA�t�v��+�y�1&u}S8?���8P?3��X���!�Eץs�\z���l�>�0��|�ߓ�{b[*��0���	r{�R�]��;���$�m�O�i!��ͫ}�e�+����C7�����C�đ����f�ޗ�\�ם�-���
�b���v�D��=�cr%�9�PP��א6P{:I�|ersft����9c��Y`�4Ro8	l
k+��쨶��ȋ��꧑�i��k�2��ϧ:�jr�H&'0et�̽����'>��5أ������Џ4�M�I�v`���F��d���hd�P��yN�z��=R�,R��JҌ�a�Y�r�'&l?Hﰍ�C��l��6wU�~VA�=|%�2��ʿaA�`F1�u�s��;[�HmC�@��s��<&�>[B���m�Le{��c�!��2��h�e�����\�n`tj�w��^ȿs��6�N�{�b#�V��Z
��4���9"۱�-s��t�'v�inĮ�+P�'���74
��]��u#EuJ�8^<�E��<�a����r��߂O7���;�P��:F��:���ܝ�Ǽ�^|_'����cy�&l��dL��e���q=��.����3�&���8���}���່�>�:�a0b��E�zoE�Fy�9����T�WRU��J�k�R��W'���ӽ\}��p�Եs�������T��,��Q�����]�u(�<����%"|Trq�zE7Y�g[8�4��Zٰ6����BD�YR�ݻ�(��]�|{L�m~9^\��c�eA����v��3a�����5�+�(��K��GF �|��������?+����?���D�w����E�q��/�xd�{�|e�'�}#Y�@�#�B����SB����܅��\J��<h�x���&�f��bu�Ǔ�i۱f�si�r	|N�����%M/d�ˏrw5��]	��FT(�W���ͫ��$~��VqV��JIjOd�:-4&�qY��m^�.�މ����9�ZGV�:b�.�G�^\��mvԮ{�����5�0���s[#��c�&��$n1zvC��7m�	��?�T`�ēO�=b�mg�ŧ��%?��S�y��<�,V��õ���ufe\dKb�w�f��C�9Ȁ�68b�UDY�k��-N�����WY������N'��^vȇ�Uy�7�H���iAcC�Э��_VF����iA���l݂�����M��s�g��ͳ����O����2��-�1�3���{N�'�C��}�*͗nZN�V[��*����y�F�[0`������}�`i2��l��čo�_�F�۵�ld]ȸcM��5,�*�g��UK9.]Ĵ���Q����7�!�C;>�2�6`��1L��{u�P���6Ա��Y�<'
�?,���1��<�e٭��局�}qՇMwE����Ȏ�dI�a�c��es�ֺ-�梥&}pc�$�>�+�O�,���@�O����P���Y�ba���s�l*��~�����\�<�敱m�[݅3`e���b �#gr���⍡���l�K����.�(����]��n����Z��Q+�b(M��i}���r/��XΝ[5f�'����P�+���9��ߝ�3{闪�;Y�C�Y���޴���Ց��(W�'֪C�!Qs�
"�BDR?�v�צ߼)qoK���	�w�'m��|f�)�Z�"&��S��U0��f��J�]8NJ$̫�d:�9gM�!B0��ː�4����u~��`F1��]��ɼ;ﶝ�k;/?BOBf,�	yn|�ޱ��T2x�>E0��>&���,¦��:��q�>m� �{~/��W��~|D-9���_eW�@5k�Y�<`�����p\�!*��r�Gs>*�!ʄ�̐���j�1��Ԁ���~VE�g���I<�!�BȮ�� ����iU�^�[�1��B��������k�+W���M{h����\�q�=�[�v���~�J�T�7{[e��2O������KK�!r�`��~O�]�=����*�5��~���J�ݎLc����)uZa'r�[�vZ��4sY�p��M���5��Ķl���l���P卬��W���֪yn��O�lߚ%52�VP�{Ս"q\�����X�;�]__�+�M�:�:?
���|�P^-Y 
i��s�<c�*�����^�}��������J�C\Zd������6���<��W4{ز.�e}�֐-t�E�XO�!2�uv��4U�a]�z#*�c��y�y]s
E���ƊOB>�g��c�M��d ��ֶ͇%d��?`m��lXMqIG�S+���;]̬��v�JZq��K\Zo��I�L��f�{�?#�X��B�Uw��U�<���T3]��.��]+J���v�,��w��:9��[�"����9���EG��nh���T)�'[g�c��c�>f��N��ϗ���j���>��=����/�[6�]Ӎ��/Hכ[kX����	���o^�K��Q7�i�{8���C��ffcF\W��f"�����J��ĨǜN����q��[�l#6�	���il�'i�d���b����_#B+���(O�Z���ͬ*"C��X���xzʥ���w�ZCY��g�e�[xLDsvL�{,�P!�Ik`mG���%L�;�y��d��\���b4	^#�h5�W�a�i~7�Py�N/ƚ� �34���+�Y�M��s\^�lz�[��O��L�z4e�;�Cm�VG��ɞ9�h�*���Vp�=(]
��l{�o��È�

� F�D����OY������F�e�48#��l�Ϟ`ߜT�#���n���0n�G����\��5�
�F�����&�����/΁DjH��	����Ř��}�i�!ԥ�?&s��K}.;�����_2c�+1o���8- o4o4��7�(��>�z�tS���R�ֲ��LM����m���o"uH���z9�ݙ��+��T�DY��N�~���5!S�*�W��c��Er���e��*��w>)���kk�*I�A(�J}���E��\Ȼ���mh9�}r�eN"T}ֲ�]t�����UE�Y��!4�����Ip���|�{�m�����Ό�$��5.������3���R�F�_[�)�0f��EĲ���Į�C����Mٳ-s����N���*�a�����v�oc������!E����Y�3&���f��V)����;�ǁh��}�TQ�Ƨt�][|���P�a���Z�q�3�h�V�O��׊�If�Y��Q
�p�����Ť��M�7�v�!pqСb�Ģr��{�����z�J�1m�4����[ʜ�����Sgn���%ʹ#.��Z���G>ki��Y�fp��|�@��Z�,�R��q��1iR��3���ۉ:��]ۏ2D��G�h.8��0��c���]	٘�)f v�X�a���="\*vTY��T��Ŷye�o��.CUѧ�:�޶��i�:�_S����n�{W�5Ր��� �U���w���s���p�����Q9��]ZX�!4r�d����=��@�̦���8gf4����:���:|�i��f�cH�t
ۣ��vW�ভT�q��y:�������'Tү���������N�,{��w`������'л8yR�iD^!|+��ڷr�R����J(jw3�wTc�:��f��cT!�6b��vT���i�8.��VУC�^l#��|��)�"c7��A�7�)����"�#y��T��`3�穹�_��{.�~�/�.9v�-XO���iFB�nf�Yk�3r�|j�Vk���F�"�4cAQ3!�qr��j�%�7��]��E�έ����˴�>��ejOK�i^�85��nfӽZ��6_ �^��Lc:�O��{�d��c��t�	�$�4AG2�
̊CVQ���تª6���>D4��T�s�����x��]�p��� �Z1�ݲT�o��}�G���:b���+7z��q�V*V��U��E��ZQ��ܳ9���Xa�ꝵ,Lk�B%Ҡw7�g4��q�YV��y����E��p��x]�B���[�v� �6m�0�)>,Z��m�ǐI�*�qlk�"���@�t�ُ�z�u�|�)�+�Wdh�,b�o(�*�ӇaV7&���3����l=�a
�R�zq�%Y�ܰ(�HI!y�r�FU�5�ͺ�ܝ��<TL�֎����cW�lM"���ky6��p���z�>�C.�kPj�d��PJ�|�Cu��@����6�.�)��))+/���ք�3$��C�0SQѭ�Un�5uvԺ
>g�������Md`�s�ftf|���'�e�g���e�"RJ�^�ϴ�!�y@D�H>)B�G��/DcR�NJ�%FIyEG��N8���Ǐ���Ǐ^��踤�'E;��|����y֎c�����F��T\��z����n<x��׏<z���I<��k&�!$�|�H1�vK\�0J��O]>8��<v��Ǐ�uѩ���:\��;'�т	�Td(� I S�O\}v�Ǐ�x��ǯC�B2I�*�$�(L �Ǔg��׽����s$��n�Lx�^Ll�y��ur�;t��޺�TH�m˚�dČa���]�GwP��\��5�_'�F����S�F{��t��uˡ��.�[9N�0I_�SI(&fm=\�fhǽ��0��"eLe#}�͑�{�o�Pdx0�
u�G���&�n8c��儶��qr���;��������PJXj��˔��o��������rZ��gk�o���O�n��V�k����6�)�x78J}a�����vO�z�g�d�X컅Y������{����|O^���]"��r)�izU?�S�l�P�r�aChͭ�|�m[sf�-�
��T
�yn-�u�|p,;�yjs3��,���b�����oծAA���s.}Yoа`��i*�|�x�4��x4y��5�Sm��ay��������f�T��`�^�� �꺜aW��C��^��&�amڵV�Z����^�`W�2�2*�6�P���t��Å�}>u�Us���#��#J�kw�W��EH��F�k�Z��̵�Se�N�ez�C"�@k���ϱT_�xZg�+�#*��:?�~�ǖ�cԅ���V�ɝ��mj^D�赱��Ŕ��_�c�}�E����A5\�B�䴎���z_���+<D7�߫{�޹1�G��u���4K�:1ߓ0g�~�5��qxhNK�?5 �<���+�\�O�Ԇ���ʾ�gOB΁>��ߧؔ^��[��hh`�~g���F��^�l��7���3~�*�^���˪���x�,�o��b�w3�	�i�h%��G�wT9��k|(U=׻����A�s�\sYR��V��;�mt��Z��
�b�/N֛ׄxՌ�d�g���BѮ6J ��7oX�1�`7���ܝ5�=o�§������!���!tr�,,b���c�L׀Oȃ���-~	r��w=?:�T�mF]�>t���ߪ��g�=�M����}\F:�����b뒄{��'cE���+I�LL���/��_���xψ���^�����M����+��_~O��"�@[[�W2����]��� Y(�g��D��
mg��G��^<�Ct�;�_��tޠo�{������МtųO��o���:�c����/f[����%)�Wy�ِ.N֢'��w��笳$���. 5��1�c�ed�;�36� W�C��j#�T���7�<Z��gOQ�(���_ٰZ�!�)�[����5�X��Yz�SRܗ�%�*!� g��4�F7t��h֜����� �|���^�n����LǭyJ��������h�鮹�3���.^ ֓��P��BW��$��b]��c+�H<�kԥ� �>)�j�yB��i�ڔ�2�c�2�''%�[㸦�D\����ֹtЋ���A�3ap;�vby>���k�ݿY/i�OyՎQ�]"���F~�:�Q�U�E�hjd���s:���u�̨��c���UI�J�� �Q��%|n�V�P�o��	�G�Q�vv�v��-�����O%���m�{R���.]]�+,�Xj��%��Q�%�N{�}&�$�"j"Qr��$XV)�Hua��>>>>>>H�Y��O�;�^Cc
? �#�=�W���>=|r�\��3E��ȇƉt����� ]4&C�d˙���ۻܢ��LKԦ�|0�t��υA�_�|��	�(��U��C��(�Eb�U�~���m�3��1�,�7�K��j��F;��H/<�|�)�����@ƗfQ�A�Ɩ�Y�8au��/���N�XG��ȝ�⮧f�'�Tw8 �൪u��ٷ�6��3�yCnX�e��O�hA�^J+|�G|�(~�<����g���U�&-��fpu�0ɠ�]ol���s���A�P�@/��@u�D�_\D�l��z|�N(_AkV�UV���WpἭ��J��#ˤL6�l���(��^	���^����� �7J�k�ƭ|��ښ����u�M@<�� �����~/��=�"T�s��+bS�~-:�-��nі����`�8���{/�ͭ�Ĵ�%)��}�/�ѭS�3�|F����\��E�5	��ȼ��*r)�1je���s@��M��<Y.2�d�4b�:ފ�P��������cj#�>Ȩ~��6��e+'د�:h��.WKa9Sx�B�`J�WD�R����Ljun�����MJxa�����w�nR��Z�� �w�^$m۸�ͺd���ֱ�Q�Ց⠒�W�vP�@�]�XG��c�Ƴ[���y�ϟ<��J�Ƙ�%�]y���o�U��{�t�iH�T�P�{Ս7�9ep�����t�w��u|��~T���<�٥��fP�<w�~�S
i���b���7V���5xm���s��ᾙ��u��h��[Q �,R���&�-�o�	���뙷xb�Kj�{:��km�<����>]6�j��?|�x�}��C����c�ZC,2�δ���MU�b�;�P��^\��Ӽ?��U)����mֺm��cd<�0|���j�<�t89,v8=�V��`,h]��@{ޓ�(t��a�"��IQ͵�|�!�Th=o��G2F!O5nOQ�!7�3�B��)�� �=?%�a��d�|gcb�y�7�ЊUW�F̺�čǠT[1�300�Ƴ\������K4�9�]�(�6k;���{Xze1M�Sl��^v[�/�'QEG7fyLX�dΰ�����#��'Sf�z����X̯K�7�~�^����A)���;��p�t�iZ�}�&�#�u���,���h|�l���,��|��}#Y��{j��5�ao֫�I���6�b�1密������7nJo �ɞ�L�No�E
�ͺ]Kw���IW;�Xs�����e+}��igԶ� �q\K3K���۾���CV�5b-Sw�E��h�]t�x���!$y��ʽ9�{��8��c�!���y}��:d�J?_��>a�g�=̚�q�h}�b�����)��XH��`E7[=��D�t~/�t��[�_b������qz��1�zd�/Tcj��5D���uz��T���xjh��LS!.x��vm��{��l�Z}���BB3|�*`�s~u7�S�X?ӫ�KO�I��}ə���<�.�.�[ṗh��$.�Q2�-���ʭB�C�x�A-oݻW�(�<�]�=%�(�K6�=*g�ܩ�������b�s��z���g��3�����l��U��j̳�^2�V0o��O�Q���Q,i҆��'���}[l�b�g�����%CC��{���*cP��(��gd�AYT�`�*�b����pˡ���ȟ;�qNh�SA�bh���y��#[��-0�N=�Ǔ�{ۀ(���)���ǻNC��캚<֛X75�͓s*�w��\��Д��!�z1�⎗ҥP��N��[B��7���#��ʧ%���u�4�F�.��ח�^��rÒ��l�C'���;E�h�%:ձ��,�'ͰUf��-�ww�.U��YZ�P�/emlBKx�w�w��IJ�)z�Q��Y_}�v�b�=㗪����I�W\��}�Gƶ��D �_P��[6���鹡�%�!���Ga��Ƕ�{8�;ab[�R]ӣ�lsڔ*f�bZ��9\;s��euo>hbȄ�� ����J�[YS�F�YBG(�ь I��R�0��Mu�.��{z�s��[�*�-af�۾�Y�5�W��aA��~�{~v�wl�8��� '��R����Q�,�Ë�	��D��}�G���U�&�'����/䌖G��,h����p큥�c	�� 0��MY��p�ƽz���v�5濕�)H��U�62#������3�>èGk��]zH�~+GߖDli�>���ٜ[M7�!�)�i�UxV�N/�ȶ��|$ַ�r��;�p�=��������V�?o�h77� qA��,��v{G�Neh�����χ�3�ϊ	�%Ҟ^11Z��`(�Iٳ�<ׄᕊ�0~?m�l�W��g :��ʃ�#ny�t�Qd6���u�s���<��㟤I����Q{�O��v{�c��U� Uo��x�g�`f��r'�;��ţ��`wvf>��X��z���ڑ1���M��"���k4"��\��=�e���q�h.YC����0�*��ͻ��eLC�gI�\[���_Mc�p��*)|.�@�ǭe��)Q�WN��)��1M^[����ULkU��-d1��FK�e�?T��dC�\���ܷ���hԲ&�J�ަ� �7c3�_Y������வ���g��<�iB=׍��+��`B�.UU��u��(��=c�1�^�<����f�:c~Q�F���(~����S߱�c Q�ʁWB�����O��<?K���X�jh�Fs���C.̵;ٯ�6EQ�^F8�ׄ����B��-�:ŹM�i)�qj�`EV����g��a�c�n�E��52���ħ,ʣ���=�dH؂�	��-�7y=OFn��xE���+�'����r����Z|�9t�T9e��CE���Pu��y���Q����7���\��}EO�i��&o����\Pcxe|��~8�|�<�︒�*�d��{[�t9O0��Jn/�1R�oR��j8�
9��2+���;=O	���.uR���6�^��B���*-����{�n��2Yrx�E65��f`[ �w�^!���o6]ʨ����LDsu�݊dM�S��Y�t�
��iIa+Z�Z3��f�q����Xl��w��D��[�͎�yO��W�EK���W<ޑ�*|g��ˊL��6�)9�����ۺ�&3A�!�F)�����?,.��_�AZo����B|�]�k;J!D����������j/���#�������n�YK۠�!Rgݼ�t�"+E�䞼˕�%(�ݏ,X��×
���h> +YNH!��]�j��=e54Prk��$�:Fuj�d��I+��͙KwBjuR����^�Ǜ����������U}��w����wFU��x�@��1���xtd>��h�a�����n�L�a�=����V��_�KC3����c?*�cI��^�O�-#^��D{���"$	S��]�kK㒵��=m#}q��W:�\@ô�@������i.�
Uެ7��E�^���W$�A����%�vJ�OÆ�L����\��`��<=ۦv��+���޿>��v#�U{~ܟ��/<�;�ʬ���@f�H]q}l g��-�R�@D&��L��P�xE6_j��>�Բ��C�=7���䡀{�HYv=C�����_��1Ck��y�ܐ�m��zUa�fvo݃ȗԮu���W�pfxmư���vmN�v��zki�^�G�h��	.*�)�p��لD��	D8zv�'Z�ـ��`S��)~�M�O���*���C:���^{��b���`c�H�U����醕R��U����8�CL�>5��d3�g,��]P�{����t�y� ���	�
8����3��>h�\H�S����6�Y75��JC�F�tû[J���xɍ�;����-WR6���r�y�_ރD�N`����\�Zu!���~��S��!E�`@vV *m��I�t&أ\ΰm���j�3*M*lcv��7��)47�˛p[�Z���ܷL}[d�wS*������y��`3	��Lmu�Z�y�j!>�M�kͼ2��\ޯr2"GZ^�G2�s#q�`^��	c��b�������>��t�C�+��
#��˟P~�K�`+�'Q�G;t�秈�Ԟ;��G��>ta��W��'g�"X_.���w�i�8��׻����XG�����v�f�5,����5�j��֒_��G3��zCϘ�@=Q>/��VVƼs����PL��f�yߝ�G�k�P1�_���z/F
�N�?oHZ�|K12��>"�vt����	GWٟ�d\#`����Α����F�'�<	@��@~�T����Q��#��f��2��۬�Zf��� �R��Ɠ�͔r}~�R1���s8�؍d�ɉ󥞳���~�f�}������bu�l��(���Κ"�ث�O��� w�H�.�D�U?m�SOx��2��C���r'~�����v��R����R���Ն��zF�Y{��UަׄIfOC�S�70�N��G4��|���I�U�F�g�/ќ�����o�7�8����a�e��J��c}U��D��s[���*��~��������ֆ�C9�Z>1Y�t��K�#{g�KX)��ݶ��m�����&��s@�Ί�w�tU�K�1�Rݗ�` �y��:H��.Xȹ�I�?�|~?����X���7�9�U��gYR�d��s�,��Lڛ��,�`w�����^$��!NiZ��q׎��R4z�N�+|b�F��,���&�쒛O{2��%�]d���ϟ}�,�q֕��><r�SP�^A(�r�!�ȁnCE(��;�sY�Je��j���c��3���멶΍�s*UK���l3z=��6�GXȦh�a��R�`(t@)AiOy=sµ�%n��~�;P�C�]��x`��o4�9��ʄ_�����WtF�~`�L����u5��=�w���ѭ���Yԑ�0�Cp����=��A9?���"]���,��v��CYS�yEg���H_�lz�u��<�]���ߥ_M�j�X�ۧT?D�u�i^���Օ}��Q�=�u����G{u���6N�[�k"l�ل�d�g��*ꯜ6�������̼����AR�j�	���/s텠2�t�#�w^�{8���L��g��.@���lvgm͇m�]h+n�gh:���D�ov��4vX�yɪhRj����x��{��>ת���[:��&٪n�RM|�e�1S=�z��d6iMYJ���)���Q,U�\��{��*{��Z��Oc�Y�b�ۂP5��|��^ۏ�]C2V�:�d��:�2�Vj���*R�Q����L�{��@sղi�Y{��iC��n�}/�3j���Kֈ��GT�B�3)�.f,�xM�n��#`����q[r�gV_��)�澒[�}Tn�a�Y3l��7*ԌvTtA�+���'uݻ�S����"h�|�2�묺�u]щ���<�X{sr��kNW*Z�lX�i�a�+&"�rv]�p�X.�'cn�Z��%
lmr�@�.�󶯚&��5���g��֊��:��u��v��嵢��<䓉�o��<v���z�ơz��Y4�.םj
,��.4Xqqk7/_tɃ^q�#�)r:��ԉ�{�[Xx�#��=]��aer46�%���S�L�FZupU�r�o����t|sIe��禳en�|�;RBJ��٭A�a�-�����Y.m�k�)���a����M-�w�5a��&t`��\n���E���}bv=�r��;1Wb	K����mt�h��b��q|�1TKfbx&*V���Xmc�9�*z�a?Ye�,��b�����ڲK
��*TohKY�M&����q���y"�5��łȭ@�d6�ە�A�&%i��?��.e��f�/�t�*c�"]Q?Jl��z��J���ة9�<S9�:�cwA՝�e���fL��/����c�M׽z�>� :$0u�:`�Td��B�X�s�i.)�����������m��N9�}P��J��:��Z�~Wa��|GQ��Mx��;;��:%op�?..mX�Yg6$4��FTM�x�񬖝�����69ST�rý�j�H��1Cd�#�{�Y�V��x&����N��a��Q�E�l;bp�d귢�{9�<ky�#j���\i���\�a��v2p�홻Hh����C�^�
i�^ll#�`�U|���ox�����4:첹�Ss9�{qu����}vh�X4i�y�t��U��7�e�-�00B���0,V�f9ݍLB�#�θ��������/es!.�.Q�;���9��5���^Y ��mϩ�M1��)���w-�]�``縉I�7�s{[B�WE�+��f��o�,��j�î�TFe:9�Y]Q+�d���2���n�;S�;.����6<���`
�ZwQd��}/>�)�ӳC�X��:c͗ǜ�&܅��MꙎ$�n�ǈ�°���eӚ��k�NK��E.i��9F��,H�̐�/��%@���W���?�&��؆8a8�M("�2�Sl��\��i$Y���F��5A�E��H�B�P2y�'��=���{�%��u�(��Dk�<�&��/{��\)13 I	��� S�v��Ǐ<~<x��ׯd�!�$!$a!��u�κ@��u��;���f�)�0O:�����\q�Ǐ�x��ס�(��*Bd��	�H��R|����I��{��Ξ����<x��׏=z�$�
&���;�2�fM�Ӆ�w��{w�:�F�~��۷��޻v��Ǐ�x��ׯHI		!$���\9�l��Y�]ܰb"��Ę����|���Yq�\�|�ɣ�Ġd��Wwi:���'�<��2d�U�]~�y�}w��	��S.�urdQ�%��^y$��vL�� .�q$�ݝܱ�>��1�]�r�z�}5��˘I��w[�@��ݐ�O������<��s���DB�^v�% !�d�;�����s�H�CD���P��1F $�q��"�Akɉ1��XM�f�nkX���|��<F�^t��b� �kJ��[�q*)e(�&�T�lm䮌�Kvr�����L.�(�Rh3��4kUu�*�VccǷePLo~�͜���I�$���������(a��7|��� ��]��^^�39�^�;=���ᷓg4�Ξ�uP�t6����/�+�b��K9m�X6�:j�����9�@�#�i�F�u#P�^6���[F:N�Z6��>���R�k`��ԇw(Y�מC�i����˝���S؍�Q[�:v��-ݹ'ѻr"�=&��{�^����������4>	砖�R�z� �����en_Zp/S��ïG;tw��a]���Qھ��e�[;�
o�v�{jo�w���k�>k�}gޫ��K;-� b�f}�ȍd���e��;��?վ�~���	��>[�$^j��}䟶�z-�{��-�讀�<O������=�V�Xu�s�	���<���s(A���L�:��1���<�Mu-UX Fua;�g+:X��*+���0��)88��&S=�
v���B3Ր���Q��n�"e>��1l	������tV�1�VC1����>�2��z��ӂ���b"����J���P+�*��]9ϛ���7ʯQ�4�4j���/?��륕e׈�G�K8ϐ�(���;�����n+v�u}�����y��bj��,b�>�G�dt
*(���޺�e`�Q���l�����&Z$�Ѓi劢!��0;����^��tq�Gq�W�)������=,��玩h��Dxǻ|�C�l2T�z�:�3��4W��]��]��ܺ�6֞|�U�r����Q�g�!��X���T���ʼ�ݫH�3s:�H��;�s�*+�w��/���ߜ[�e�ӗ�_N�4��uQI+.Gv��F��4�i2�ؔh�y�x]��~�d^���~Q�7/|�-߳�hn���RI�J&V��������{�@����?>tE����Y
b1�S0�=w�%/�g�6j��ե�F���ڇ��Ί�k�
���E�_�S$e�{Ӱ-�MH{�~�y����Y	���,O�oSj��f��7\d�w��h����4
��t5���}r{=�&&��1VS)��;��j��͘�����6��tf0v��Ǚ����u�\/ueaB�s�3߬V�gD�?5B���{יP5>S��me��
4�{�CI#9��.��ZUF�ܙږ���.w:�&��c�Y����񬂛�ډ����y���y��o~N��H�b����k{>�,۽Ƴ��V1���)���5f�Vt��n��q/�?+�M%Rɹ�V��țƏ*��7w-�_:.{����s4�r���A�w}'�s9Z����y�/og�^8ΑG�ؑ�_"c�o��nM./��j]>�;��*ե�>?}�[�>5Ck���vi��ƭ��_U#���b�~�L�[�Ⱦ���I�{Pz���j�D!uSܯ�#�͹} ޘ��Bcc�W���k�ͬ�)��}yČ���G�>+h���� w~�<~�������]\iͽ̷}5
��nq�j����b�^�\w���*a'ٰ��1E�4)�rr�T^�F�#�=]�|τ��������8�]�si�k���:�.�M3V7!1Ҕr���׸�����sM�׼h�Ɂ� ��>���h��}oq�&}$q�b$`@Es����m�)H��oj���A� ��0�zew��r���+�_*�Yɨ�9�}�վ��rWN��mL!���k�ܕ�8���(lظͨ�)۳���S���>�W�fu&��F�����|��cǵ��{�w����6ni���0d�h-fE�ܛ�Ӽ�����'k殝^//�>�Ş/���z��@�J�H��傭�T�nI�?L��t�`��9�o���~����3 ��	�j�X����Swm���a^`�ZϗW�Y�r>C�T{z�H&)l�����G/[���&^�
�9ڟpT�ы���FvL��OI44��s"�f�b��^���שȵ}���7�R���]T�h��\�'���MC����20u��Ѳ��M�f�ʽ^K�����"�V.��XIo�Ʀ���&��[o7t�vԢ��dO�6��z3�]ǯ��-��ZY�܌��=#i�;�fg��+�ٶg����d��h�[ޘ#fzWsESS�A�	��ڽ���O����t�_��7�gY���/�6g��e��10`�nFF@�i�v�昑[]��Wq�\:xT�%1�/4�EV1����c�~�/{���'�U
]�M��O�X�U�-U�nI�}l2%ݟ�������SQ��������օ�(��5;��%��/7Z߄�"�kc�Қ��p�z+d��v�����%������B0�~n$"d��N�54Ԯ/�1�c��77&sW����Ά��7���<��-���G�k�*+�H���W�yVOqR�g*�Ϲ�_,޷�x1ڽb��9�Ӫ:��e>�b3wA��4���n��bcV[;����O�C`zv'�AqS��aU��o���}& {��M��^l�@�'���A ��b�R���ߞ�T} V>�~�m9;~��o�4^��Eߺ:�?��ĨB�U����vE�2��V
�u����ԛ
�ש�oN�qdΚL��^�mM��z&VS��|�l�̗N�.��K/f��F0O��E3�3ؐ%P��u#Sj����@5L���*�rl�Gwl]ϳ:c�K�Q|�lDva��z݉��:y�q�V/�}��	w'��<3x�I�-�H~�~�"�:>��꫺~���p1>��u���U�|��/@���h��~-Q��Q��	��jI]a�0�u2(��ЕYO.�F)����i���6�*]��^~d�q�%eVf$m?e+1�b^�E�i{��5��M�C�\�Mͽ���zr+Hu����0��:oR��8�e��TF<h���e+�ݩ�eD�	5sivz6a��!{bS7'\�/��ڛo78;�X+}���������n]�jkԂ7��Nv�ݍ���r��Y�7�s�IQ���]w�gfn3(������B���*��U��t3�K����p��<��b���/��2��J�+L+��i�n�GT�j�Y,x�q�U��MD�rhs�6��6y�Ω�x�yYC����P��>ײ�5�mv�8���F/b	�=;�b��:g�z������ېö�k �-��GW1u�f���C�YS��fF��yKG�V�-`�����ު[���%
w�	��=pj������"!4�v"�9�	�Q�O�ŏ_����
�q5'��K�	�P�g���.6���)��9[�3-�Z#Fw
�3�����.Q�|=�ÿ�KY�8��m��;P�5�Pع����p*31�}�g��ģE��zۆ����e���~rx�����qc`�RZ�e��X�	.��N�q1\��O���������=�ټ�M�䕣�\B+n��>�4���L��7(r��r˷��R�eu�\ح�:���o����l8Y6��.��sa|'.�1�c�9�xw�N��������͏��l��$6�.�b��e���DCV-��͗��b'���E��^%�(�\���T����Gs]i�w���.kOb�g5ݑ޶U�N�9,EO�r��st�gΜ ��:f�+Oq�^2�ef�r=m�;�5v9M�&�.5|��ds���!�b�f���޽gg;�
�p�N�Y����n�(��H����ʅ�5�7j��ow���1��جd�ܙ*�M�iaV�>�`�_��W���6�/��wmv�G]�zm�=��s���� ;n�$mQ����� ;�i،���z�G�\�Q�އmK�k���j�����B���K��|��2�'+����~3��K���ƥoO�vy�6��عu]��ݺf���wHsPy^�-"=}��/��d�ooW�5�K}$����'�:/~���:�:^�/Ǌ2���jA�R�*���|�嗸w�nn\c֡�>�[�+2�"N.���m"(���*� AT��&=���[�m�*�u͗��,�w�ƣ��U�LԨ`y��ݭ�5@�<)P=M_�)���0����ѷ��1��9��o���y��6����J��[���� �pݰ닾�:P��ћyy{����#vӓ3�n��)}�#�L޽��o@}�A�lo�f�uH�~Dv���&Ա%�b@��\�
��/�,��H:�;_���>�.�7�.�w��&
B����=�_`S4�%�r��n��7cא�O;�]Z<���N�2�"������k�TK�@tv:\`L����	�V5U�V3MsKj�sV������A�&�Vm��ׯ��]=�/��C����΋��,Y��=��`�n�o_|���ƶT���u#�(����DMЪ/����]J��Q-D{yo蠷��D.���~��~zv*f�K��4��J�;sw�W(�t��p�+1Fx���dZ��D�mY���y��;Z\�-����l��2W�ͷ�c\��9*�T�����qi�eF�����
��]K���*^�g�rRWSb�^���[���90�Q:4�s��4Qfs��ak��ED>8U�%� ���=���nƫ5�45��v��krb�[^�^Z���,����
�8��@�T�I��ޮ���h������]��*���)�1פ=������?W���d�A$%��>v�>��u���x@�s�P+����á,���;[3����ѳ��mgR�4������[�*�!�A�o��p���;.&�{+�6/��Nt��;�Rou�]�آ��0l5�ׅ���zWTr��j�ZvG:��^t;\	Zs_�6��%�Q�h}�ɗ���a��2���@v��"�UPe�=%H~N7W7.XՇ����0v��GfZ�I�;�ܫ�=���Պ)�j��e I��5oqƌ��Pm�Uj�Sr��z��C�v�vuT�`�Q��ݵ���[�@�{�r��X��ە[»�S�F���<y��Y�?�*���gWA��soA���*W�}mʞ� ��Ě�9�~�������N
�=��vR�}"T)�=z.�K�M6p�3�����Iu\��$��f;�:�L]���4��q�!Y��d��a�������_,0Mt1��Q�<�(�u<c�rs�m�x��l;B��ݬ�l�a��y�1�}U<2�����?*���wm�|+�-l�r��s-lYk�&�N�(BfeC�y]�q��u�U�R�4��ط����1����w�|>]_�����%���l{��Z�!*�]O�6��/ǎ�-�~i�M����H~ˑJ�,�דױr7L����	���Ox���x��ƞ�pݬ�ׁV�=^�����/Ax������C��'��{3���eR��%����dz|��S��e'��]y��7�Ceu�ٜ��������^Ͷ����W��_���5p�M�!�kM����X�����-ds���E,ٸ���W[Y�%�?���ܻ}/���͝w7��u�0q���f�v��COl���y��@�ok�m��ѕ�R��m��%��NoIڞ[�!���x��oQ�d;�[ckw��Lp>�t�3Y�q���۱�6�y�m]�@d(�U�4:V�+���I�~����Pn�����g�p�������'�^��W�qE^2^@~��ݓ�J���dt����*ԥ�+6��.�ؒbl�V��I���p]����,ͭ�.����k���p�ǒ�A��1'�l�a�ͬ�U��Cǀz��-�j����ѱ"��#͝S�}�l]�t���,�jd�9r�Ox�^�����;�|�/����=�V\�D���+nh���o���zL����2ިc��9�oiL�U�y�b|oV�#�z-ڱ�!;��P-�p�ཪm=��(��ǚ��!���gW0��B����dL�;,��b�l�������sĪە�g�C�j��SɈ+/;]�3�Q�7�%���[���0>�IR��[i�!�!6��OG}]�v-�T҇t��k�)���lj��N�۱���e�jp3GulEj'4V�[����]��=B��j2f��D���<=ʕĬ�7��ml7�x(�ۃ�&/�g3X�p�t��'M�H*������*�-t�s�`�oGk���-�ʡ�NY���k���N�`egs�d�M>7�\��AX��y�6�:�rVe��,����%��6����q�,�w,��v!�$|�N�,T�ܺ����z.�����mۆn�H�\YM�����ɩ⻛�Cr��0]��k\�z�5䡄�U<b,���w��÷lҭ�ʵ�jd�op��՜Ź���h-0�O%�7v�$�\7#�����LԶ�����[�T�z6���-�]�-Ʌ]T(�� //m6g6u�B����~h{W���R����߹�ܭp>!������iS1L� ,.�o��jҡ|�����)�#�n�E��'t�U>�sc�֧/v�0^��l�]��E�CC����wAv���<�f\��wM�.P5���pGa�u��f�M��3��ln>�f_G��^˺b���x5R7�}��%���7��n�qFz[�]T�r��^���5>�jNBV�u��	�Ƒ �5`�[�N���ub���MZ�����X܂�鋄ռY�qP��'PU}]&۸c]0���v@�.�Q�8ڥ������nir�_��c�,�5�۹B��4��Y�f87-f(N����g�1ś�K�#aF�v�1藏.�>�us�ch5拗����$�6�$U��Z}w+��:�a��r�{xesE��`FZ��l�e1K�E1u)݂�t;�7n^�9/��ޥ��FW<"�c��5��-9ټ��egN5 ,����n�M�c wj���soR�|�g-!k�/kw��ۮ�5�����p��ӻ����nv����k�fЕ��<ׅ,hc�:k��M���iwT2���|/��<z;t�ᙂ�u36�v�7W@��̶0^9�*:�����jQ�_(`����E�ȳw����_64�qξ͑8�sS/k��9�_=�����0��/��i��3w\4�uُ�a (�()�L3v��{��\x��Ǐx���;$���O*��n���H��׋�$��B��5��aa�@�PI	Bn!#6�����<x��׏={ԓ�RI"BB�@ӻ��9�rIC&�!��Ɲ��O��ѧ�^�8�Ǐ<x��Ǐ\zFB@/�8Q@)Nr1~�@#4םu�M*I ��$��<��t�ׯ�8��Ǐ;z���;v���2T�!L�b�&Rw;pd%�t���wn"�r�G�\�;q�HK��@�&A�e�1��h�̡?<�1!��@2sv��)���D�
=/��`�����七D|��Ȥ�!�HC���[��؉��Dْ��$c�R�i3H��# D����R(�JG�W%���_\��w�<��ڻ�񾃚����[���w�C���HQ�[���B����-w�:V����������ͯ��G��ߺ����V�����2��3
�B��J����	�W�������K>�(8�	���F���>�n;��@���0�m�f��u'��'�m���LD7_*�5<z�`�p����0#���H���=���SH��fE�yM�ؾ��6^���y���*�g�?U,*g�����S�y����g�M���S�lW�����q��v���o��K�R�ϡV>��N��{�l>��l���x�V/�U3֗���xT=]��C^�c>�V�F�;@��a�c�C)������ٟ �]�d��l�7�Ͳ��Z1�iq^��'+ҭ��ڱߢs0>d�R�=Ang[=�7-��x�P���w
�-V��U䑫��U���ܐ��Ó������>mK����5{LV9;(�*��Z�
�[)�˺��g/�ߟ�Rȏl��nY�(�	%1g���x����Љ�S�����u:d��x������!�\W�b�������yW�Ld˿�op�L5�B�0=�>�36+��qc���ض]�9cn�k4����:�n>{r�j�Lyy��o7���H�Z8����?�M��n�˲�.��yPJ=KV]4�&�n���3E�cu'&\�L��u-q���"|��Wsw�R�w�sʴ����T�_����	Bn�}�[�VT�+3//"�������ֺ]���pا0%w|��z ?kJŵ�ׯ�{�K��ex9;�Vt�����ɷ�!oT�즈���q딺l��:�wd
�kЬ8�o]���
kFNkl�:�q{d���g���R�ɷa��w�W�k�W�qi����7�]LFb�;�����-d�T�22L��l��F+x���i�����e�N�ݸ?I���u�v{Kq��Jb����CevPm�ǧ���m��Z�z���+a���x�Hu#��K�wv�?WLq++͇D�czp�Cf��cL��֧�wk3L��7��3���ֻY���w+}~��T3'���U7�O.���7Bb�4����{�8��*DПM�2S��]��"*��I3����͎OӐn�}V8�m4��Yp���E��8!��4(/{?;��P���n�ɧ�R��]X�e�t�x丞�����ֹL7Ja��͓�Y�Z�e� �JV�W�& E쏕��&�t�L���F�~m��M6�.GR��3��>>>�����L�Ϯ��oo�_kK�I-�"zP)m��y�������[�<;��#w2�=�֝y�,X�Sz�ZY6��#�Ax�+<ʽ�.}+�7�5k����列�`��G���\�>�z�U\n�])�7��I���p��ն�O�ߦ�(�2��Y�}Q������������������؛ۍsR-��ySyQ[?Go�i�K?H?O="zR�^o���5r�WU�[��ɺ��,��K�-[9�.�٦M����gڲ���1!nԆ�ĭ�[��\/1ژ����bo�va��c�0b�]�^Vm������3ך2�D����!f�c����үwѧ���n]�Gz�wf���t�[v�rL~ڠcn1�`D�7��rs�v��`ᇣH�&�'��Z�7�.R�V��y,f֬�aM����ݞ1U�B���^�#�w�s��+Ⱥ�p���w2�+��鿿:#:�5��Vm�K,u�I�dT�왓v�O\����D�[xuY�3�;=Ьt��m��bd�<����f�DNM�Z����6�rZ�"��'��_�2Q�wx+K`���sOI�����U�W|���k�fK���?Ji��iY�}��V��|�M}��m�g��7*�?�cQ���ս��QfD�<��3)K�����5�w����&��6��]5���^ݫa���XDꛉ�ن�ݫ$A�
3�!��ϛy�T�V�Ͱl
�6@g6���m�bU�A)�u,�����<yT��_�5��h�e�ԍui��u��y�/b�f��h#'���h
`�@�dv'~�s�⛂
�A�cϛ�"iU��l�b"9�H��۷ZC=�/��u�k��~��p~g�w[)4���7L)�Fv����$ީ��L���QW�+�IH.��Q�R�r��K~��n����9�_8�s�t7�y��-�q��U�?;�����Λ[��R[�^
jdQ�S��]-wW~7(��0)��"�sn�T���ގ9b�l�����Wq5���~~����lU�=�wY��ׄ�.��B�{�F;WsH��JuȺ��ܫ�6��W��#����?_����4����-P�*F9��ԟR�]��.�_ι�X��Kc=Z3�8Z�ۄބ��qIN��S����֧/5:w�������^���hd���|�gI_5?��{�MϜ�x�CL��ͱ�u.�ւ��ht\ěn�ꊌw���*o3K��.=oḂ.(��X���7�KB�Ź#�������Z�t�;�%��sǌ�cL+ו��]{����]�F�-V
'�y�wr��sj��D.� 9/[>CFX�7gH��b����~U��[B�8j5��'G��i�';�K���-%�Ϭm�[�m���\Н�|j5G��e�-�M6f�s������k�D8޸ƻ����a�il�08S_>WL�T�5����Dn{=f��콕�W�p.8�0�����n��!�#{Eno3n�gQʧp��:��N}��'S�����2��V���y�����f�.�5��oZ��WOO�k��ߧ����ͻ��F�6g3Vk�#SS{ga��Qu�IOj�=�=���
��@�Q��?l[�h��sJ�Ү������{K3#r�3v���б� �1�M��7'h�6�v���u�<��~Azj�{]B`���E���{�Ә�rf{�I7ZWӷ�v\��>�\$�Pa7/_ E>��\y���怦�)��i�y���
�y��ϡ���y.����ac�띫��<=o��I �M��5�Rcz����t`��ur^��
�~iP�/֤�{�-��w�����S(�i���L�b�@(/�6��gî��{J��Վ��UPZ沋�ƺ��%�G.��r3�mcoX�G*P,ᨫW��o2���8r�UƄd�l�[��#��4�{��-�~�裱�v�����-�*���b���:x��Q���w=A��p��5��ߙdʭ��:��>;���7�v6���3��=9i�BK+�Qs{MG�َ�\3�{����os	��.�l�=~�&�w_��e?b�RM9�3n�O� D-�gx�e;���z����sH�]ݠZX���q	�m7>��w�U��S�̷�&߭�yyS
*�g��UV���e\Zpq�Zb�͏z��-����qWR5���^;*�
n1S���mJ�a�"�bX�F�W��w�Ȱ�!�Yn�ٌ̼v���]m��C�O6��T���u��;��4Mv&8�f��-��c�qAt�<�)��O����:wiA`f�ܼ��F�:Ӗ-�ʗ ̶���		��� ���^^K���S5H���9b�����h܉9�\$��w��,����>�.K�rod���>����OT�Y9�e����\�ϕ!�[�{auLa3gM��n�Xo$X >��>�������x�{���DfS8uU����E�������0Ǯ�=<��]�
x���=�݀�3��Zё���3g�s˝vÁ��X�\�ߛ_7��(�����sJ��o(���ZnR�nR����0�y�s>��.t�4&�7M{�j3��*�Vd � ���7��B6���\H���7p�l�S0�s�Ӌ��󙹹E�0^��U Zf��C��QQ� F��H�����_��É�p��v�=��vB%/�����&�IF�*�����ngHa���ٙ�~��
��M�{���ݷ��aZu���tJ�G+*�L�WVl��ݲ�9W"�-�w2t40`������@i�u�{�t����ն��E����=�$#���W�I����f���NCu�dܙ��D-�5X0AR#*��^:����[�o*�%��f��G-:�[.��q��jwN1�j��h�K]s��[������^���o7���)�)Вj���O�N��f�9��}���Cc��v�|���Ty�g~���y�QP3d#�%�R�ʲ8_�'*���5bQ8�����n��>�����]�>�����Ε�_0�Ɔ���~��µ���{B��D1�XfF-Y}��Qݹl	�al�u3����+s�[��h�F���M�}��g{nr���q��;��y�n�Z�Ѷ8�O{\��4��ؘ*۫��4���m+73���[�,r��v�����H��؍A0^�5��a�}�S^��D3(�X�K��pn��n������k�sz�XB{�^t�GЩN��t��Df��ۮ���]X2���܃��Z��G�˧��ُ��n�\��&��w ���b[\Mm���k-h��grG�т��5��"e��ndZ��j`mt
Hky�f���t܏�Pr��7���9�O����e��a�i]:.譅:!�N�s*eҺ\q\��D��Ld����	�e���2�t7�ol���;�6�x}����y�?�� `��t�ھ!W[�>�7��C����٧�L�j`�qȨ�dfVì�۽��u׾�ډ]����6	��r�~�V��k�5�Hc����n�D�
�����9)PY��8���I�W��'�ۦ�^�����t�_>����&�w"��md�U|��i�c^��U�;���H?��Ӽvz��@��1q@��y��$�iGc^9o��q�.ȕה���(1Nck76$�a�.����D��(ޣ���%�ؼ�F�N��t+��}���Mt �s~�-� �Fhϴ��Z�v��M\�N�Շ_D���?%����K6^�p����e@=;h͸*����\�zb�kQ��^I8��
��$�s_M���j�gfZ]�S��5��O���F�7�Wn�e��z�r�$�Mpѽ�;�}^s��lP�te���8c�g�xݝ�zJ���{g�̸s �?	 �p\���_Psvk��H����YK��q:��;Z>��{3��R����ǜ�����7g��I��Bq]�M�W����:m%a��;�+��\�+/�9ai�ݘ���{=����w������i��4r���T��?\7c����YƘ�[�⪮b���*p��sK�ɶ�����b��n��R��x��7z�gS]�c��Ւ�uQ�fa��*�:��
 �Q����7����;�"��X�{�]��Ӓ�էu�3Mn���k?d.䪜7�S�M>�ꂽ�3nÃ�6��*Xp�������C'��eֱ̪�Ŷ���V�?m#���:��<�����}ӒM1ҏ6h�՛��=��z����K�~
�+99�Y�1[�t��w� �6�Ju�}~�7��{��a���ڠU�T�@���V�)Z�^��k�	]C/u��[l�������ou_�p*�1�� ����
�[���Q]�e��t���}�|�~ͷc0�D���>�ޱ5�W�s9K��[�-��'�@���u�\Fmi�ݧ�U�pW_��ɭQ}�R�����U�Haf����Ά��U�gQ"`�|�S���Yy.Y39=�^��_c*e͠;�^_�/c�&�����K���o-H����w�����7�-Q��]=��-8���ά�3�z#�cC�c%���B�M���F�gdl���ZI���)2�N��\���� �-�d�C���nY@����f�[*R����*�J]]񐆵�DF<B89-�ϭ.�x����{V��m����md�7&�:\,�i%�8��䵷}�|-uh9�V6SD�l���L�E^�
�i�f��\��<ЌZ{@P��,`�!�׶(�u�:�0&�F��#7�5y@�m�[�
�G�(Z�2jUpf�������V{��W,K�`����]���Kئ[��*�A�+�t�8���YS�f���c3v����#PsQ�\[���#�.�s��ǹ�l:MY�6�e��5jK"��]�X�u%�:�2=�OS�p�B�^*��Ԕ�qÕƏ��;(v�iU�J ���U��λ�vr�8'\�q�Y.�s*�_=8��4�	sC�eC���Hf�]���L0��W�]�f�C���%9�G�Ϧ��4�{j�޴�T��UP]u�u�pֲX�f�fu�plx˔q�y�^}[r�Yl80��W� ÷H�K2���;B�)%�Rh�)U[�xj��p e�o��PD�C0�	�S{v�����aRמ.Mf�F�V1N^�f�*�7O-�Lg)�d�͛%Ѻ�̰Wq�M�+A�liU&����g/�3R^�+8BdF�5!E�E� O�b�&D�
���
���5��bvз�@�^4��u���c�Ww�1>�/MEA��1��w�Q�C8�
/N�&���vn����88�Ђ=N�DZ��9�B�`�1S���X]x�P�j�M`f�j�{�:�;�7;[V�
��r[|J��)��Z�n�VEj+w���qU9�z^�:���v��X�I������6N�$Ԟ�lI&�8'U��Wp`���f�D�,���Q��a�4����o/���%[{z#M7��q��j�䁗+\o��m�ޠ������'yF�:��ˡڅoo`'5����c5ӓM��ǵ��� I6����:��M]t��>m���.j.�mE�d�^�f嵚.P|�<-�r���j�� �i�z�hBete�u�h�6�f�`�tu>ݵ��
,�/6-K�i▝�����q���U&Z�^r�Ւ��C��!Da;z�:W�#Y���_+<���������J�
��md�SSz���Ǽә����{��=O)��9\q�	5.�1��-�ڗam෮�\�����)�!5`��w�#z�Ў#���UC�:�˙���v���C�����.���J�d�DC�	��%�ԅ��(*���%0�`�ۨ��^�B[p���Q�1p�$�@��E#Rz@��(D��U\f*j�h��yF���,�iQR�|H���.���I0F	��0R���df�@�#F@�c���v�۷o����ѿ�7��"��](�L��FM��I�_:��^y�Y����\ĳF�z���nݻv�뷯\�!�P�43�!��6��d��qW.`��:z����nݻv�뷯^���`�I4i2�h�뤇��WM�B3@�u�bA�E�����z���nݻv�߻�~��~��NFe?{�Q�]���!H���I�4���0�`�2d/�:>��IcF
DB��17�ndȃL�μe�W&h����.�xf�"$��HF�(�Xk���\�f'���@Y%�˸Ĕ�t�C�w{��آIY�L��̘�)��\��0�_]u��$��K�$LW��D�3O;�h0(�#=]K�\@���1��q@���߇��y�|\� OŠ�l\�ظ�X�lĴo^u�J�k#�V��v�x)�oUT}�3��vw��]��&(xm4sE���o��������t�"IE5.�uR�j�
�j�S[z�i��������Oy��}E3@�C-HRO���.��'��R��Bǭ-Z-yw�㜍�.�J� �5g�����]�j1.����HO�ן��u�m���33C>'x؛�ؗ�'P��{+�yT��%oH���]�,:�Zո91����$���Os���z����k��a�3ͦ1uh��Uŧ�O�q��z����g�u��@e���\�|9!����]��Yk��*�����D����!̜�X�=���EًYm�4ioU�d�i֑�n��lϟ�9�:>����K�2�<B�{%h��x��x�B2	�×�o�,�ڟ5�"�7{d����l,�/���;�G��	��u����϶�����R1v���K�S��ҧn2�b��c��=R9-��;��ֵFꘛ�WfV8��/ f#=��O`^˫�6=��pdb����死P"��͸�Z��kk.��E��K�FȞ��x�f�ˁnș�2���+�gG(4��l��]���i�s�<%�*�En�A�^��rSGiCϒy�c��/-��%�"�����y��o7��T��nT������-w5~�a�m\z�}NF��~$�\Yߢ���"��G����8���}��Q�!��@l�MR��}W�4��7��2���i�v�5S]�Do*���.�.�֘������um�yV@�.�D2�Ȗ�y�__�0鞠۵����j�����2��Y�k���-�gΗ�54&.�Q�z9@�x?����"h71g`��Wf�'��{z��Rx�e��Q�x�U^��M�^�Y�������ZC��r<cX�9QV()�Ƕw-��o��[>ot�3;�6.�}S=S�gtRS[��WRT
�<�~QmN��6����c&��k;߳��1Hް�L7�朓:�y�c�����KF	�]���K��}��t��ٸ<���2#���!`}<��"�谊����||f�}����#������Q�y]��W��M���y�R�ӕ.�s��jә�j�.Y!�7�`m�ux��j�;2l��4�ʚf�)�5{�e���TW�\9�U�H������ǉ��J'{J=1�=��jŭBӲ��y��YP�jڌ�FY|K�|n��2�3�T� �o7�����kR%ZM��T� Q�ƌ����Lx�$_fԻ�>�b�G\w3�rTN���s���E�`P��Z��m�)@�a��WB�V�:��y����Y�d�D�*�}��4+z�,��j�RS�z�݇Z���C�K�Jn��eH���{YŖ�GMlf�z%�����r5��N��an�)Ď;A�h�kR�z���S��&v����m�R�K��\Mr8�4��{��g��x�m���r�K��)۷f\��3���Ϋ~� ���崲J�� �J��Y�S��]>k�a>��騡���]�^j~vu�Q� �;����g+�����r���i3gˊD[i��[؉}�F���"�<�hH��^9i�y��ym#{;-M6�Ie���`��a�]�e�,(���H��&��Jļ��XX������P��t�y\w2}ĤR4�`K'���m��,^�^_�kz����Uҁ330h�����F�ԤŴ�3i9>	o,��*������kf�f�N�R̀�ښ��֕{^{[�=ɿh��{�73�#���4�ƱotԥHM��m/����g,7<:���-�)�:_2�c"�m��;�^�^�@�V�`:|�vN����2Θ}ߧ�
��i�����ܰ�9�i���%��K�C���lgS�^�T�Ե���Y~H�i�:<���h�-+�\���LFs̥�L/�;��b�H�VWk�Dqg�{w�uz��X��^W��GV��Z���-���z�:�����<��%p�ܬ?Th���p�+/��[Lд�K�7C0�Te�6^��o�c���,oo\{��SU�ٺQ�swZD�}�>d/<���Hz�bv!i{��z�wq�!ܴM�;��y�y��R��/W�x�f�j�e}���0R�f���������7�;u�����2b�n��e�N�:텛�xʚ�F]V���4E��+9[�g� �x��rr��m���b\૏;�r��7�J��H����������C� ��_~�s"YF׋�ɝB���l��7}-��{�Mq���|���z��UU�0�T.��+6h]Yr���d�d+(6�����w��q<�u�]��T!�n%��=�x]��v�O�R"�j=�dS:�C\θ���X}<����щʩ/4�d�P/����////��/���rQ�Wv{��l&p$DDf?Ҥ�l${	ux�����-�&E�w3	T�6�}S�+	�x+�U��^6j'�O�Gh.��eyz�����2��~]f��m̥��%�bF?��W+�z���Ru�>؎Jp�{Q���'�su��?f�e���l�/�?�zf��M��=P���Z�_s;�ԭ�����uώÑ}�e����d�uzx���󽙗`�xoK�`c�Ϯ��0�C��h�a�b)���'?Ez"�=�oӪ�R�?���[1�q���,�� �~�N�y	���i`��ݝI�r�X�������͎�d����ޅ�=����cͼ�L�=��%tی��;���~!���Ry멻�Q�3F�?#Z�����o@tZ���n����U��x<yj����Ǝ�h8���Z��©z9A����q�;$ee;�|y8���ϻ���;_���J�ر�}e�'-L�ߩu�4K��ü�t�c|e��x4δ�c�yV��[����Q�?"!~ hz���s;���a:H8;�W�f�x/�Ө
��9o4�J���Ӽs���:�m�#������������M�p�;W���"WO�@�`�<�{�q��Lʺ�q(u�U���v��αp}�{�sQ��8��9�λa�}8/��Qѻ��Iژl��Sx�<eKn�ɠ��V%n�e������
/�M����G�\-K�s�B�Q�8�3���̷�2��q�V&v�H!�a��S>�]4���!�֯/�F*])�Q�Y��Y��MBl4��N��jw4Fuz����j�=M�c[����J���5��(a��F�V�~�����^?�$6C;�3�fY�5��(%yES��l�q������<�8f�=.��?4�}c�z��U:\<Q꧂�%�6�����vq��}���S��}).��zE�p�p����>K<���dJ�ʎ��ٗ�/�$ƌ��B�]��>��78r�
(��=6V�1Kc�;rG�96�s�P#�g=q�������67_셺A�[B;��->�2������f��`�4t��vzϞ�hPfy���]��z��GR*�/��}�46z������u[�|��j��u���b٥�5ެ�[|%�n��_��S������������[��,,�+��[��q�.6))��ޠ.�IW��=Y�����8�,�x�}��F8k��}��� �踻ܪPYl�z��uB�`����}�gt��=D������m>h�:-��n�:���D��\�q�no�d�qe�^}����gؠyŸm-lY��|.�;?&mG��'�f,[�*�*��aX='ܱf&�W�f���&�~����l�J&7p\�͋�
��Ϧ�C�-��tQ1�1��:!��b�Q<�ӱ��m�{��!C	�v�!״o=9r"o�`�L��r��x�h�5f�c���b�r0��'��=u1�L�,��\QQ]w[�O6{�mb�v�ٱk5��ѵ�b�Ufj��]�-�1�z�!d1������v*%�ק�����r*�~�$����g�jZ�W7�E�w��ؗ�߿x���o��9L`�+��1-A�����Ԏ���v«��Cf<�)]��Ė��1���G�#+x��ک�+��67��o�F=	��Iv�u�e��(�E�V�nĴT�oY�ʉ���kt!H�4��KNSX��*�u�_�4�1�|�����o�y{����K{!.fd��ꅛu61�K]�43Wl�r����gkz_�/"{�h�]��y[y"�\򻉽�O�f:�*�����g�t"�o9��8���;�+��#^yP�+6�$���	�B�%��y��|��h��M���{�B�l3�E��,�ޝ�7���m���٫=�f$���8�Mߔ��<���(F��� �i͟f��`��1�0�q��Z��)�d�i%ed�~N�b�A�t��1]�U蚧g�����}\���Jl 1#��H�j�F<��H�gcy���d�)�WD�[þj���ެO�G��pEO����F�>�v��Y����e�Nil���Sl�̥^�>k�P��L`͏�X.i��x���*�6t��^F|��Dy"Łֲ�*�{�U�[^��q__��k�~�Y�ɘ��s(�YǴ~��4�^��ڒN�||�
�(S��65R��]j�B(��T��s1�[;孒�d''(������+�{�.I��˲T��Nk���u���2.��0���3�2>wECu6-+��^F�X����eu&]n󳷔�JIZ�GŶ\i2��ԄԜ~?i�1�j�zouS5����2J�=��i>��p�{��l���;Yn�K�k�vc���,��iNPk�hյ�>B�thΓ}������2���B3�״u�"+/�=�=�S��b�3[Y�*:��s3�\񧁑�� �h��9���/�d�!��hCt�fbξ���"T�0�R�$���J��N�h��w����F�R����a8�/%�JW�F�w^�/����ój�f��S�=���g7�f^�˗}^m��qur�\�7�1��ɼ�T5���ޕ�$Z����k������y�[��&�8��>O���]&}��Y�������zh��3Hwvd��\*��O�Vx	�)�ڴ1/��e�s��]��y.Ky��ճ�9կ4��>�s�A/�����{�:�Z6��f�/1B�#a��	`�y�Lv+(�������$����P�5|~�zIl����E�q��<ʛ�N�l*�v�;f����BV��2��ƛ�V��h)�a�.�H��&�5
xIb����Eɽ��;ĝ,f�C������\ӄ�J,�o�-:�>0���;�,�{�b�S�pdA���^��n��O_�c��c�3�����|�_R�;�7�ccԢNm��H+w|w 0�1�;U�z��cH��i��݉��@,5��Hb��x�A��q�h����-�]{r��k�8�~��˖�������ju
�CKMg�/֛G �R�fEʎ�v�iW�n�7��ߛ�S�E�~�D:��\3��y�
�v�&��q]ͶHxޞ����7�����&`�d2Ά� d~耯�<����Y���_J݂*�@�����6i�i�s�K�v��i�ͲO{�o>�z;�@}���_�}��Y�hݵ丅�̮BV�� �D��ޖ?w(3����^<�/�W�i��t	�.3�u�,@�+5��"����ϛ�v8U�+m�2Z�UFZ�j�LT�S����a�7�Vf�>ԭͼ �\�r�e��+�3{�_0�i��l���~:��y]�R3����\��+�����l�b�T�cy���ՠ�L�A+�*X�WWsoK:��Թ�i���f]懌�З�Ym�uӂJ�{��ͬ�K�|/@e�����m\N�0�m]-�{K��)gg&�rX�e�7W�����-���2Cݩ��,�G'^�X�%���,0�k�kf:	c�,�@{vG�d�.^�꒔���?e:�g]N)6�tۜ��Y����a�G9�itz��X��R��=�]v毫3�c���Nto��	-غ�f�ç��˵�O��@KC��ɔk3����eM�t���(�R��L���޺�v��R��ڽM6�����d!�r��brv�(%n��n�A���V�U�TΣ�$���W��w$�6�htf�"�ll�kk��5E��O0�t�SWٹZ�]���fmlu׊�DG�fj�l��$s�o4^L1rգ1��B�*�tKp��L@���K;�Es-+���#�Yyt�K��t��:���+Ӻ���lVE#����;׭�+un�B)��PX�-K��K���%+���*��6���K��ګe�LM��(a)U�e�	�7uV�C��	GTE1}3�vm���x��f;Nd�x�-kv�ۭ�Jz�V�\����(neF(X��Gm���2���&��ы�6U1]�t[	Z���U��>C:]�H�*�=��I�83�o\د�;���h��0Xc����P`�N�˨��������Z=�3��ʕ���TT�SU�*:�1�N[bC�@����v����o�%Β�"#����{�ؿ�3�rs�I��Z7 ��i�&�S�y]+�:��"��
�h!����M숥�U3�0v;v-�Nu%��,��v`��7�)��c�;�nbhit�&dZ����z1o�#%V"	�,������i�M�v��hËt�w�zrZ��eWׅ��r[���!�M�b��M��6���=���C�Zc8خ��mt�Xu�^�}�T�J�l����Êa}vt��·��eD1��u�F���e�S�T�\�"�s*"�m�'�s��7wDVW����:�2VKj��w�2ơ�s��j�r42�#9S�\,����M7��vݬk�u7)R��4��)ՠ�c���2�Sui����[��HZSKnZ�ܕ2�s2�d��9}�TW�r�FDc�\9�4<�V]����f>�xT7%[��aͫ�2ҭ��Y���'"�#Yx�T���AZ���V<5i`}�y��2��/v3�!�ٲ�l�JT6z0V<��;�ӆ9q�Oyt��L�����#%"[Ńd�H$���@ �K̑1<rRN�wtg������ S���_\v�۷n�_�^��H�'�[��r�HJ@	�͙�h����"&33{�w���7���{�۷nݽq����uOe�#F�{�%7�� ��"F	I�$!����߻o�v�۷n޽z�:@�I�T��V�� ��塿zᦃ*x4��D�H�@���z��nݻv��ׯ\�$I�*H�1�Bz��W2H��Ѵ[�r�<<}y�ҹ��0EfX�޺Sî�y��\e;�����34� 5%�6�h��s�����S�s�#AhH�f
� DWw`�ٻsn����z�cx�_M�c�Q=�@;��y�������l�c# b �(�c1I�x	 ���!ݘܫ�n��]��ʜh2jD���O3z�����Yͺ�-��Bʇ�3UR�^ӫϱ���<���2��_�c����V�]y������7+�Ϣ��Y�[�l�@b㫙�v�����"iS�W��[�%�0a��P��	e�[�ӊ��k(r��;�,��c7�\���˪y�'��aV,���"Z愲���j2+vŪ|g�6sFdrۜ�׍�ъ�(��W��U����H�nD��9k�;��Y�h��C��4�k��:nCa����.2����<{�k�pr��<D�ۜ7����c�?~��}c���@���|	(�yF��^����;k��^��k�6q��V�@�?U��fq��';ٸ�6�Q��EÚ�S���^�wJ~������{Uг���{�t��������-�k>>�x��x�u��1����4�Y�gc��+���\�g��k総ZhM�׺�'�X�i��8ޱB����1��ę2_Oo����0����ju���%ͧ�UY8��3k�N���g���e��8�Sx��n"-�^�{�����^~S3{G�.���\V�I���`����w�O��tJ���UL|J8A65�gܒ�_��������&�>I��~y��o7�����{�4,�1��;����ǡ&��U�����l�7>;�Ō�2�?4trm;yַ8+�3��k��V�Y�=��SVr��}!?���T3�p�f�.�ӷ���B�<�b&��r{��ݠ�4e�Xb�^�g��ؗm˖�]��UsKk�5c�]~�g�5=X�Uz��䟺b��{�ڟ�Z9=;�������rGvE�@�e#�p����sR���d+���-/Me��H�|[�K�}]�oVWxI�:�C%[Ȥ�nLѦo3���w�Ť�����8��}����
Gu;.ޝ0��S4�UϹ���j�-��l�>w�ZޞM�}e'ų�3]`�p�j�+3���] ^NPǶ�7#�TcRq�M>]�s�d�-� �R����]T�^N��фq�s�Q]�X�A��G����w���)�����Y&������p��v�jgAG	�M���0"Afk��n��跆�>~�<g��i�_���(�Q�5YJ�hQD�
��u"]��I�<�6v���ntoe�����96��+ٽ��\����R�d	A�Ǽ�˾��waE��IM˚E�)��Q��(��Q�L)(Ͼ������������_�r��;�yߙ�l�}?\]3���GO��I�yk^�cư�sE	�s��1V��WɂmJ}�DG@{��#�~�P��B޲�fr��H�x��l��|�n=�H��4��*���53ӭ~'����7���&�W)߲�@l�S)�����2�*:�:qlڹřؔ��[7r����+��er�������۵��݆I�FaP�勞�iz���h�����tg��u� 7����o�^޷3p��]� �����6�l�n^o��U2�[��xք�,����Hw�	����zT`���d-l�y��ׄ>a�j��'Bx�)P�s������^����h���Z��X!٩�'��A�jB�V��0k�v�Qw	W�ã'"��T1�:[�n���a��Cv�<ʭ�U��M�}��#���������[��@�[�G]���RZ���'[�R��u.��̳���U��o]cQ�R�2��v��(��z0gd}$���8XGu3�/��U���[7��|b�メB�'�L^c�acm0c�P������Ow� �����yx9�7��j�������(���Y��*CϜb�\��'n����#�ot5�����*�����K�B⳺�/�n��
�XwK�w�L���{8�q��˓��ޡ�*�W�n)_7�xXG�=�0�	�X�M䌲b;�5��9x[�5��E���&�u���,�ͥ򙪘��j����'������P�S�P
Y�[����'�v��y�%�V��T�Ǔ��!�g�g���2����kC�L�?" #�^7�]��L80qP�>�ލ����}�I?Y˔ر�By��s���WN税}YG��Ǵ�}��;/_�Ѵ*~��4u3M�0.�r�����f���8�'\�{����Y�|=u���vdEв����M��Y��61���s�<���p���zg9�gƢ�XǷ%��PAіU� P���fԫp��ܷ虽Ύ�rS�MT����׋�}w��ԋ<�{%%{y`�
4N�2��	��ǣ����:��5ӕ��6K���s�/ Q̧��c���_6��.����c1�����V}����������3���E�r�.!eIS�NĊ�n��7_�����6d����"��M�NڣY]�c�䮜G<�W���}v���KuzM�Ƨ�?\���3^xQ����ʚ�`��;x��36e�����n
�=�;ڗ�g�VڸW,�Ƀ�*{��G��W#���Mu�T�_ߡ�K��&�%��I��2��Z+�l�}�bqM�W&J<Vc��2Z�{f�9m膌}ݮDG6��;B4��]<�VX)oW����6��̉t
zjrǠ1�j�#y�ώ�.���|�YYc�7��m,=+�{F�Е�6�K��ۻ\Э�I�.Tq�f�F3���-�@;Ը�[��OY�X0Ùf�ޥ$�	۞=�!�h���ls��}�L�oO<��zI�~��y"KV>�R	���rG8����m�r��
�+vo�]�Z��)��<R�˱���ޝ�.�9�i�/��eX�$�s���*��>C�줐��T	�D����ٔ*�A����3�:S4��n��[��)�PF+Y��fSB�!r_s7�|�ߤUװuf~U=�O���y��o7����U�`��`����R��c�Qݺ��"��;�0��#����o8X�1w����%�I��NM�{�o�g�$�n{=|tϻ�mo�j<����w�����	<y H$����c��XΟz=�;�K@~�H��Dw1&��qc��Q��4�L���z��/*XWoZX8٪e��ok���k��\�����+�L��tbE��
���qmnȬ֐s�F���ڛ=�f�x�,`��1�9�īSf��k^,��ܤ�u�@&�=��X�Ӱ��jY�"��l4�N�,��Zo2��@����7C��X�-�=v�����Å{ԫw�0�ړ���)>:�(��J��ؕLݛt��"�%��o *��tzm�>j�}���ֈ�Zy����Bⶲ:UK��g�sN�:���p�zy�g1QX�LC9�s���q�g|�w%�@�W�����=����=�c#���[&�d�ݐ�6dD,Oh6F���Wp���۸gz������纰������8t��egKȪ��ыC���9.������F1�תkB�Nd�]BY3�$��$՗.���o�1���=�UY�^w�>Q�=�4�m�x�'����/��/P��#��"�?�y�#��x��B����%����k��:Km^X~���,~��{91݂�C���Y�8*W�<;�j�����c:�3��7UrJ�s�����+��JӦ���>�e�#W#V�Zݲ����ކ����1w���;�"��t�wd��#m�����3gH���/B�~�N�cǬR�]��ޏO&Zv��%'f"���dkV��`s5�:4>��6��1��;�Ȋ"t๮��1��_/_Lb���0��ȴ*�m�\�I���u����v.�j˽h:sI�ͦ�#�f�5�'�"ڱ£�װ��{��ؕV�n���$��E��j#.D�%F�Ns�Y��}����%a��g�qT��H��w,�ދ�p�$4kK���zY��hf��z�An�D�^D>�_q�����(L5��lUy���vB�O
b���^�e��JKo�w^�޲��w(�~'∄Q>7��=����V.��ir-��f���b��L0��u���c�л�OZ���]-ߪ7��Jz�tp��u}�1���feo7�����������|����k�\U3��ȷ�P���l��h�NO��6��B��۽��7���*�ݛ{�>zd܁�|Ƣ�# j�����t2�a����U+"[D��:(g����>�"������ ��uJM�93�<%�~��I��p�*Cs��G�λu��7jn���߻Kϕ�,g�aelQ�W�5s=��ƻ&��ժ�L���0����� �?��7�Zg�kiѓ/Q�������%	�o RΡu�9V���ʣ�o��&0�iu��5���CGy��zE��z�|��{GlRŀ*�z��mF��=�8�(�#y�o Jn�y�6��E?J��_&�����ˎ*옼��^3�b�{Z_���5��6���c�Z���R�>��[.�S[z�٫���͗�Ei���{���~U�_l���k����;��Y ���^�S�p���\��f8�k-	�כ���BbT-�v�Z��zo5�E��W@��ٓc�]G�Q�+���	�b��21��2���'PS�M\t�]Ң|ٓ��z�6�l�O��W7�,��V�S��rݱ.�U����i���x�}��|�濽ڳ׽�(���lo�yqL5�ޜ���9���c���	G��ډ�m~���#����Lb�{s:2")�֞����!/s�+9����qǏ^�;��� ։0�su�Bb�Ɯ�9�}4�m
����=^��`�ޡ�q����@�n��M9Of���ϭ�ل���@3��ǟ� �\�XT�݋x�����1o�͵E�K5�p}�/�0ag�j\���f�U��zل��L8���g�õ�{��E�	9����<M��k2��T�z���ix�#jw2��F^-����7�ָ3�^5s�U̬����'��n�[k�ڎ3��vO$�LR����iU	qd�WUR<
��C2��d)��Jz �a�.���b����=�C�g��U�Б�aK��0^q뉥Wܮ�xjjMՅ�B4K\p)ۍ��U��#���j:%\��o�I�0g�m]w��N��\���r�O?�?{W}�Q���j� ��\TS6���"��ϸ�ղ�h
HG�0����p'�B��n�\�l#k;/^&�"����xyo,��vR��=_i��`Up@+#�wB�Ա��y�]�y�aws�VWA>�6X_hg�1�{�2y)��6������d��2�Y��jN�O{we�j��6�7# �����S�*zE��Ja��N�iiJ�)[��QؼN�x��([;#s<��^���(��Ĳ�LUZռ�ӝ��!��W���Vovx�M{[�w{<��ؖ�u��b�O�4��:�W�;=8���N�m
Զ9WH�i���_�}r��\�1k1�]4���᳔��k�36��d�d�ͱ
��n������iðz��:�%b���ʸ�vC]��ȸr�15U���ה�k���"!�����N|�Ÿ�c�/��ꢸ Ftظ]��4��Ў�;ﵽ��Ni��k�y�?�����וH�b���((#��Ȉ�� Q�AE_�EP"T�j&��L�Ҳ��������f�+6�VkiY��K2�-M,��,ԶҲ��K6��eVj2Ֆ,ֲśk1c5Y���Vf�5��e[5�ٌc+i�,�[i��em2jkk�[u��ՙ������V���l�UfL�c*�fjٔ�i��f�YU�T��flԪ�fLe[32c5l�Z�[iX�b��54�m����Y����J�ZX�[f,e�2�[iYZͲjm���ef֙i�[J�k1�-iYZ�ʴ��ee�-M,�iYkL�Sm�b��$!�(��0����]-�e����>u�VVkef��������VZ���VU���Y�++eel���ʲ�[+-ef�U���[+5eel���b�(�`,`�w����@`� � V���J�mT���J�Z�Ym� 1@.�hD@ 1P@ 1D��JͭT��j�e�T�
�kZ҈(�@`)R�֪Vj�J�mT��UJ�کYV�Vmj��[�j�f��VU����R���Vmj�eZ�Y���0ִ�BHY�Jʴ�֥e�+5�Q 1��R��H����iY�J�m1�J@`)���(�րt(J�m1�mJ��VZҲ����VU�e�+-k��ڴ�եe�1����5iYV�����Y�J�m4�#O����@�p(�~��"�� �
��I������7��6}������O��O���_�G�������>O�
 *��?����TU��E a �C�H �������`���~����V��
�~��M����NX�����
k�4(+��֔�MM���JU�5��kM*Ҧ�,�K-i��+5�i�J�Zm6��V�lզ��5�i��ҩ�M6��J��Z�ٶ�R�M�mM�[J��֕��m��5iU*�ٵ���KY[J�mMR��YV�i���ZU�Z[KjY��ԫJ�֖m�l��T#HTH�Q"��M6֔��U����ZRT	dA�DdT��U *
��*H�� �c��6�kQ���I���i*�U�U��L֢�2ڙ���jM�)[]y�j�C���O�
Ƞ"� �H (�<�����А3�?�-L�7�+� �����������y�z0?ߌ?������( �����O����br  
�� U�(~l�C��DQT�u�AW� ��(?������PP�W�x�G^G����- U���C�~����@_��$�o�|�����a����Љ�����PW�ڟ�������4'濱!� �������\S���u3�$��E |BH?����B��ہ��}�_��_�TE��l
�Z���S���>����
C�O��PVI��k>����` �������G�>� �T)IE���P 5��QIJHKZ[bU�;j�H�T�cUJUT��H�QV��Rɪ�U)*��R)�,n۵�j�i�U��w���5�Tk�3��GW�1Pm���n�wk���C�ij�T�f�pk#�N�m����J���m�ZM����vb�Y�����c����Cm�WQ��]a���l�������5a3���ݦ���f�]t�Ð�Wm&C��ݝl̛f�(wwkZ���m�ʄ繗E<J麚�  ��&���U�����R�R�N��9��h5Y��m�)��uڔ�!���r�b�Lݺ��v��z;�����i�*��+[�8
�MU۷U]�f��(�+�  ���P�B������|��HH���}d�;<�P�Q텱�Mv�^�Ϛ�l�m�'��։HT�V4е����I(�Gj�����ݽ�������NpSM-m����C-��)��zpv�5  n�T�V��ʭ�(+F˾�z:ʪ]��l��N�� �B�a�bY�ܒ@.��kB@�^��U�%��۷ ��f�!�V���4U���wwk� �>%E�q��AUP�����*���J*���p�()rjQR4X��
с��+@�� �/^K�n�j̍��εm��8U�| Ͼ�H*��y� �z �)�8t
Q9�»1$w��TUꁨ��۰�U�N �kJ�u�[�kj�6ݷ+Jض�m���  }���wv�xh��հP�PQm��T��քW�(�ASUXP
�+`j��n��@H#{׼T��/a�B-"M�����ak�u��  <
��4Bgۀ �v��4 ��  ]  �` m����  vJ�  Z�p (5׻)��6ӣUM��M+w�   �>  �ۨ  ;]k�j����   ���  �`�� [w`  .��  �0@j�p  #�zݫ�iu��J����g��   ;_  ��ܽ����� (6{�  �^��
F��E�g  ږ
 �X  *˛� �Bj�ٹ4k���)s�:9F�  ��  g��� �]��x: q�@�Wg  ���  �� ��� �v\v�  |���R�  E=�	)*B4��5M��USH �O��Jh� �T�I�U%�P  $�J�U �������?��c�{��N�Dj'�����R���"�=��2�"e{^���|>��}������ֵ���UU���mkZ��mkZ���ֵ�kUUm����N���% 𔰓�R���(3�m���;����տ��h�{��}�Vv��b�jt���e���V�X.����V�K��n-X2��E[0&U��کD
.\�ã{��ZGn�7hU�N�����\�`ݖڸ�f��֮z+�_Q/��E��3n`���f�H��n�^Sٷ�q2��[I t��\�K6k0�wA�3JLYu�M�?m���lȑٲ��y���ƀ ̙�u\j�[<�ܢ�r^�E6)�m ̅BQQ���;�7�����x�4�ل��/V�oD?I�.�Q�t)��*��a�nR�a�1L��en9�d@�`*��h�Ie��V8%ܲ1��J2�
�F��,Y[�4�%+E,�V�5�桮�����!JVO�k-��� ���J��&��+�D����aHb��)RV���hn,�~ݒ��6��L}%�B���lf`+��Չ�-[��Y�����nC���3X0#4ExJ�~E�<�Y�ܼ�.�u!7�Fr�C�x��l�Х����;J��x
5�ɛ��X�]�f�l��1i�7����ŵux�Ҋf򜻷�Y��X�D��#���`�
�5�Z"�G�T�c��Pi�wX�N9�p;YkrV
��AX�P�B=���VR��o/*�6�r�q���.eEHe#i�qk�[��2n���������M�IInE��d�Ʋ��5����ʳyaR�[I)D�hkK/m���`#����5�Y���"_�bY4���5�$����ݷS�3p�ݵ,I=h�^�89����x��ĝ�|K[��ㆈY4�.�	]f���V��(�b�j��F�ՎA�"�o7��[�p8+-�h4K��TPݵh��U4c��׃jM/��ҭ��,�xB�G�x`�%x^9X�J�3x�,Yw�JjS�Xv�a�*��7#��j�����ŋ��]��X^Nv�YV��ݡz��6�C��Kӆ����&�nՅ��Ԍ����T.T�-z�j+��:Ǜ�M�d���ϵR��MPJ͛�1��%:l�,��lĵE��P`��j��L/S�Й��T
��ek@4�{3 ?h��U��,�.�0^2�H�A"J�.���&���̒�m�)]h{S&Gը3D����C��kjÊ��y{V��)�LHD�0Y���c%c�H;����i[���L�(#����(e)���(�&L�ۀ#7�-�V�;P��R��#(8o\X(�j�������������;�M��WB�Y�-�jn<ͦ��ۉ�����-�m��VD�-:R"X�]d�ɒD���7[.�$a]�Uz*+��`�wpm�V��ݙ"�"$"ᛶ�`�U�X!�l2�Rf(��S>�nC[b�lMӂ����(�Ni9yNk)W2�Hɵ��ۣ��å�k��,��b��7[��Ʉ��d�X�5f�1����+��f�$aR�z7.�)�M��jm� ̶ab��Ջi�2�K�nbڈ�������[1�;�5�=�	�q�z.���B��I6f�n�|Y��&�ί C6�Xv*Ikv44l�F��1 V$IC�S.�X!*��w���r��h�j�Ȯ��v��h�I蠘n��Fn��X��5u-�$;��$@˽7&���2�Uvۻ���m�]+�~�M9�M�pV^�4�,��ݸn�7jB6�e���\Á)��:J���� q8�3#�z�f�L˓qn�v X�.�5����w@���8�����+ۢ�\�jL&XVUM$CX�5��ڛnf/��IwF]�׮�g���)�]��Vi���32�[+K�afe��l�w��ne^�u����sϺ�]�i�S]p(w+Ts/�m���坠�W2���M: T���2����n`j�Ȳ�i�fe�@4�Rm��{��F�ENS�X��0���hD�D��������[�7a
'��`�c�)�cv��y�$!9j�d�zbI,���� �]ꙭ��ygo�"�Q�Y���d�R�t�	�A7�����(�i���іr���R�i�� ��[��6(�S*J�v��Nk���.����e��F�IVNF��܍�밝�e��3$X�RvǸ0H�#Aj��jR6��;
^Q�O�d��8)�lk4����I�L3l;��<�\��b���C/U��?���*�"�k�
�慗xC��j�;E�b\��EZ#S�i�Ք���ڊE�u���/%,�7��U�9�4W��d�D<���.�@/ҷ&[g4U�vR=4�pˣii7��QoH���;(<[EL MH֐-�����o,�u�\	(6�>_)�.6����kECJ�I�sH��{�Ԃ����1�"�,���"��ܙt� �k�~�f�t�[�չj��`��4���Ye�b2滼b��+U ��m��n[�^���4'
�qu-��U1��.J�H�
��3�A^��>F��/'C��{��v�%���)��k��@ .Z��
5x�Ui*�0AyM:�ծ����x3I7��D�b���Y�-m��t�%CKL�r��=�U5��Ue���w1ӟ!{Or<\N^�`� �U���3Ǚ�y�����02�^� �hK$�a=k�WLT�6�"� Jt3Ytrm+��2�0#s$ަi��j�ƦX��l����2��t66��%h�kR7,� �i�&H�ֽWnX�����a��,p=��{4r"���p��]��7j`�1kf1f�S�^�I�hْ���y�.XʇX�)����u���'U-�0���.e�)��%mSR@�;Cn�c�:PJ�MK���zF�kC5L�Ԗ�]_��H���$��k�ɢ�-�2D@��&ȺxB�n2Ю�P1��8�o�25Y��V\l����n��H7��%��>wQ�%�҅���Ԗ�D����w�9��|�ݗ	��{f�y����[he�Bj��fX��nL���*�)e�#;u-0W���j�Wod��v�L�H4�Z��mɇb��A�]�;��[j�@�M��/Q65؈����m����޵V�)U��ٱ�\�)��1�h%�B+"VaOvn%Dڒ},��/>���2^bzFY0�N�V!x�e�����bS/L`�f�P�&J:BN�3ks5��θ[�Q (lfk�E�Q���\��hi	Q���&��2Uݠ�g�\�᫠^P�i�/�A(���!�wb�i�,ă�Q�Pԙ�]�=2!&��������P�bX�v+-S�>w�&�+!����v1� �K`
1��-ZU����2k� b���)Y��-��a�[/��^U�x�ӑU��u�"�6�+Nѫ�ymd&(��E+�XK)�T	�VfB��Z��cY �FIWF���!�P��kX/	�ON�{�u$�L4�$Ū��-:��Y���J](�4ԤM&kߕe�E���l;e�h��J��E���� �=�PꗙZ�vɠ,��u��wPۢc�{��O�S"�߱��l�9u;�6�pf6�1���oI�w��L�+)l;0	x�dܤ+t�F͹Yh�Z�iӨpM�W z�)m`;Mh�_�X�9a�`���a$9R���1�[�5��ɂ�Kw�{�������Ē�<x�L[�0mm����2�X������z��&ډ��T�C�x0-������1I��ᗓ3kM��Xa�R�[��	>��*��LH0M{�A��4��b#+* �e�9�ҕ��m�V�^���F���NԅM[y�����ɟ#��|��H8@X��%J^ۘ)�I�&�U�Y�j�԰�T�ӭ��d*ʓrͧ�1If��X�"�	�T�����X�$+,�~m:j��[�b�	�&�0ѡ�^�t���F��������u��/fb�76�1�z"�s-�ݦü��Y��n2-YZ�l[�S:[`V�Hf	Bщ�x��Su�P� h��)ʛ�,t˺���b(���֕E�rI��v�ǃA[�B��V&��06��Aj3� �t,̥���i��ـ���י�Z=��$�k�r��e[�l��J�C��4�l�X(*5�SU�	 ���fڭ�	��ɒ��ݹ�ER��ْ��5L" ���X�[wc�̳j�MY�Rx��k/s#В3K�a^��l7,[��,7�w��)�:��w��	��"��v�0�T��w�N^�����z1k-ilV-`�$�N����gە-�-3VjUjʕv�5,�8�Д0j(XS�X�$��u{���Gl5i��Wr-�ж���e���%h��l�i�R@�7nKX�
�<4!DZEm=��lߦ��ux/ d���%4]�_I�I[6L6��l�z���P:�)�M���K2J8�6��K��pcvi��@�K][ݠ�f+	�5��`u�3S�V���]��t�ϵ(�o=~�u�-��i�wn�`� ]&��V����{�2�*ۑ�)�г^�HMS-�ɼ�-1��-���1��'�A�5���I�����4U�85ck®��P�YE�S5��4����df�Ś�v�11aE�[��ҳ7�8�x�T*f�{���>ٗ���~��BH�M��A�.Z�����f���3e��7Uf�;D��������E�΄��ib�t�Es.�f�&3u ,e��X�n�,w`��jeK�f�2�os\��S)9J��p�a�cIYe�-�C^)E��i�%Ek&��U�)��YVrM�
6��I���;Z��$�
!-i�6�U0ZߤR=$#z�v�Gf�`h��l�e�Uh5X�Z���
���%"��ܒ���׮�-����	Kpa[kr����6B�z
���B���U�����&M*#���{��U�V�	j �V�l�%Jt����m�P,�hLǮk� �޻ݎ�4�Z�Ta�ͻr��L`��u&:˖B(��0>���a��� ز����AL0��1��f̧SRt�����a�z4|2�:����\R�t�^���	��i��H>�{YB2��;��$k`��[0��r��L%s6Њ���R(�F]�Ua��X�Ȓ�;��B�m�v���b��e��Q�x�go�EQ�5�Z��(�i{b�)�V �(���nS�t�����&��U��ob,���ˤU={�43=ut�Q�U�wX�I&��U��ɺv7G"0���AVH[ҙ��;��`V��Z��n �b���t*��y�E��0#P�]REw-M۵��ے�MA���:aM�L� �8�df]�V��9��^�e��s=ݽnݭV�`�@�z�q(����/�=&��wH$'/��q����T94C�Ã�P�����·c�E
C6�Qne=�Ǣ���,Z��vs��b�`�iJ4�v���ʼ�zB�Ԑ�KX���.�"zP�$�C-��!:�0�͂��Ze,��b����[rɫK�,��1�;`0�f�׵3pn,G���&XOh����ɚ� ���CjP��Cq������p����V��&[xHe�r�Dz-��A��ڈ�k��`ؕD��be�w$�B��]��D�΀���l���R9�,U��LQz񇱼��Z@�(ġ )��n!n;���rf�y�ˈ+�Y@a�?6w&|r����P��Zyz#�c)եyVt/+|�#.�G&
�i2^Y��X/(!5[�YB�J; T�^���ލƵ�n���"Rlu � [��	����/:Xk)���܈o�ctR��̑i���@GAM-ʒi�Bf��˻�.�<[�H��a*���f)�ُc�Z��jƼ
�-��X%�I���h��Ԭ��+&�J�iё�,6���,c�1��L��)^��D�0®U�m+�ݔcp�h�v�U����U�K�k*MH���q�O1'�Ei�-f^Rr�ի1Ax�B� [�ccV[�:y�j��R�k��O� ۥ1[S.�6V�mB�Ocu�u9R�ňj�ʏn�L��sVf�-F�l�����+��y�2�^*�- m�j�p�#-*P�H^}�����xLư��:��m�E��×qlT칐d#5xq%HÀ�3w1D�-�wAz��a��cv�r���l���~ۘ9hO{�ac��ȸI;%��H�{��i@��lB��b�V���UB�ǐ&��x����[sotRGLu�Rг5�Ғ'�ik�	k)���f��!�f�0��C�[��֠pX��1�D��J;zb4�ڃD��wW����XE�ZXN�4^��Ьc?Y���[�ph�����&b4$�ѠU*pçp\��lQ|nlI'3;������*���"Oj;����死b�jJ��$^8�11Ʈ���Ka�w �k��H�C�n�����6Ҡ�b�16-�)�R��XM�IHr�杠��iK-U,�M���9u�Q܏5֍.V����MҎC���:�Dȵ�\X)��VFn��u���zP;��F��Ĩ�um�YS5̻��,G7kZܙ�(��}�6��b�*q�`��l�Ď�x;Yl�Xҷ�=�Tqm����5bڦ�m7Hl����������ね݃!�M��%��(N��]��+hĖ��B�4��v���QfJ����Er�W�C�(��H��ͩM��i ���{��^JɁK�Ow>%�֐
N��a.����<U2��*j�2�uaVq��u�ɎŜ��5m��� ����� [�ڪ���j1B��}=U���%F�6��ɵ
;�ϩ�{b>P��5�Y{�v��Hx`��Ȁ��Ӯ*e�NXY����p�0�u#�M�-��������+������^v�$�����àR��*�yA�o�����{ڕ�oE�ˆ2�]�.2�W4W�?h�WR5�R;���s�6�=�_��蹛h�$�j����{0���p&rҏ>;*]$<eq�ƚ8��c���𮡭���fMW��s�0>Heݼ����%�턱�{����RWM`�D�.9uvj��u��	��&�ͬ��q9����w"Ҟ���gIS6�D�%c����t���2hŰ�qv�2� ��`�:5�Gy*۩m$+�kF�>����N��ӆ`�m�Vsm@�Y�K%��]8���X	l3�]��h9d�&���0g%H\�x�04�}��dӃ7{�N�A]+���}r@�-S��,b��[z7Uk]/��\�/�ς�P}g{[b�6���Fw(�XPbɸ�벞����>E�b��73��Dt�֔�L&-c���'��}��
����^N���5��Qû���;�*	���U�v����ۺd&9%�Z�}�[<��.A5�ۉ/T}�ӽ�F)��NYŶ5��;�\ƅ|R�0H���Z[���r{�9f�i�����V��Nq����&��Ѐq^Վ�VW����Yu�����4�[������;��=�m���(�hv��Os��4#�eț����K��o�]���8�N��Z���%�!LL�Μ	u;�fh�kT���U�j�kAX��KViM���J�"�� ���!j�K3�/��G��Y�:�@��H���N�O���[�{16q�*�����,fW}�RzaD�n��.���]\�\9��ſYr�5�C���٩.Y:��e][�X��ts�F���/.��g�L	 �E]�P����K=�=�1�3"�ձ�缴���W�9v�*��},�]di�Y��	���a��珺��\̻��CR���EVͭl�� E�
$To��Pe��je����th���v1S-ٛj��z�:E��@��%�x�VoP�v^��T*�7;h�׼�Gp���!j�R� ���f�>�ގ��ه�c��8��$���F��K�L��܂������}Ο6��:�펜e��nc�o9��z���̺�����5'���<H<����6R��qy�2Iw�;���y�u��1���}q��˻#�A��=B�G�� ٵ��t�	M����f�����X̮ ��lR$g,ޗ�q�ގn��u����]������� �';+�U�Ynݱ�ə�,��Y���7�K�GNCV��C��@6n���V�����W'm
��+��r�vh��r�te����Z�����Ők��W@&T�nG��a����oz�߳�J2]�Ι5�w0WfcR�M%Zב)���E�ԛ3�����9x&m�=�������+�T�nK��`o��<S�X2����h6J����&k��*B0�;V��h��_;�<ܧ�Ը)h�}�K��<�����-ٔz�w8�[7˧��8X��B���zGA�����Ǝ�{�b��]��	X��tu@:�&�X���+4F��� ��h�J/C>�=���(��$�Ո�b��n�T ζ���Rsc��f�ݛFU���L�ɳD���{B�� ��qm+@���a ������ԯ���PYIl
���]���)����;7sJ��rv ���[��e��&�W��T�8��/gAWȾ���"U
'����n!�w.�L�R��k~AA�����α}�{��G�dr�,»X���{8Qj���b�}�y1�y_&�r$���)Z��o`��V|a5ҹ���j�2nn#��͆�Cn��k��L�W6��M�������[G+�$�6N�����CX����Qx��=��;��A�����v�]	�vG ����P�Tv��fJЯz����|­��w���wj\��WI:xܕ�2�Vy�������#+��,Qդ/u>��>��V�l{Krb�Gk�d����J��(�K_
�n.�υdJ'p���/�
��15#�F����C	V�E�?I�]���<�nӅ���M�jӑ��)|]�G�Q�ǂA�e�=��TXE�+�@#�kF�b�fu���,�������)�tǼM;�)��?<+D�(ֆ�		��X�7��/tv	n�QSW�)��q�q��dБ~	���[�-���'�_�����O{�����-[��T��Ṵ�M-n��WZ�\�eՔ���.09�	�2+��ƷJ�)*4EJ�8��id��]���*Li�+0`���U���]tfﱒV�\�ub!Ӳ�^����Zc���*��z��=�/��}�sO<!�X�;q���R��V?dߺx�Ɔ�!&��%��8r�#��I��x�s^njD+3r�׬=�$�L�f�oO;
��R��5��K��fg%,\�y4.V�"v��A�}�z��k�/ �۬-�uj/j�u�]��>�%j6}����!�|��]��Nܝ-�^���\��P�1#u��N��=�]B�^��>�ͯo�>���ɼ�+v�}9h\u]�0(Mh�/JhW��SŴxW�M���f�qAK��K>&(�_fC�d���v�DӜu$�=ǷKW�A�mf�������AC�'G���Uwa�F�钻�N�W1�}0!s�(4���G���
�Ūݩ�]��9P��u�ީ^��#Yk���Б�y]�V��(�݀�����k#�w��gIw���9��5x	�Ŏݐ�ne���o9�ؓ�b�X�:�{������|tiR�Pu1�]��C�S�|2��s�-=e��E]	ڢ0O���/��)W�"�5hX:Z�#�⢮�M�Og�k4�xC�њs��N!xj���BlJ���Qmx���n{��vR�:�1T)��e�&�g�d��0tYeq`�W%A�OxQ�2�MwI�r���������Qָ�J�T�W���]7��+nU0d>������h��IÝus���1�p�rt����*Vd��l+Mxǚ��]3���휣x��+��`P�h�Cs�p.=�d�I+w�oqx�;|��]7{Ɗ�IcĴ�F�eNk��M�1�隸e�� Vm|�̠��GL:%���=����.y�fʂ~���',?$�V!ݣki�����=I�;E̎�{��Οds�މ�X]S��2 G3xz]-8�3) �J�͙`A����z���&�aS�]��e�*ꏻ@ ��i"a�g�]��og�#�;���KWۻ��ۭP�iݍF��̖�}Zٸ���-�l�;��RtUj.�2���G������\:v�B=/:�3m�97����x�=p`@e��ڱ��7���Hx��Ӷ1}��e2�.��鉉G���4���J)&z-h��wLTӻ��*�y�x��A���b�3�Jv�74n�g>�h�/l�^ {� hp
Q8F��fq��)��w(Jw�Q�5	%�H���V��ם>�OS�����
���e��]�\��yN'��B�Sx���[�P0³�q@UX��w|�����eeI�݊/!S,��r�����q73��\�4Xčl��IfN� ��ͤv�E�7�
�����
hb�N�8	�Ӏ�0S�V%�ծ�oo����wGؼ�外�TN���O�M�J��QE.��A�yu����4�^��������6
�.-S�<;D7�	1�.%b�s���.�]�n%�,�O��wB�{j�I��g`em��n����S&;��i���n�[�M���G:e.7�o_LK%�}|Wb�.v ƞj�[��P�T��ٵu�K����@q��h=�%Z[�������Kӷx���z �`��s����l���G�[�k�kdܯ-�{!�՛���Sיs{T݀(� 1qT��y�t9�w��(�B�oM9����m�;OI �U��F�`�Q������n�#��lj��	R�*e<�u�Pm��4`qC�{Fs�-�s/��)����I��k5a�
�Zr�K�5�a������m��s�����<1���F���C�s�j�3�޳���<ػ���-zkw�Bkz��Ό��W��-:��p����{H��Pyeڶo#�{@Է,��+/R�K�������6Mj�vn�ԖV�=�U��η�1$e����8�$��@����Q����1_��۞A�-������o��j8�R������.F��ݶ��u�
#�Ҥ{8�Z�"�_E��*��&m�1����pl��[�m&�#�s�Wf��;O��R�K�v+Ӑ�Hp��p�z{�Uz��v�˸�-:�	�\�ɷ,.��o ԕ,K�5���[w�M��,�
;WQ��Y%`�y����<*���9l;7�#���vgoE��o��0XSy�$��W�髾�u���;�������Q�N\Uu��Jm7|yә��V��-�z��녑홅�ӷܳ�%Ӓ�&��C�Q�W|L�Q��p���]������tm<h�v�An�pga���:T��m+�E#N��Fe��;�	I���uyFP�3>4�W)O�r��ã�Ơ��~�0LU���4q�V'T|2ڽ�ɫ��
g���1��meM�5���h �� ~�	k���Z���W_B�X�%����$wQ`��贶�u❜'Jʛ!��Ƞ�^g/��pbQOo��ȴ]׸�T���Q��^ε���<ka���d��-;Й���&݋,V�s��wf�Pk��������3��\$��[�������n���"����ewn7|VN���l0��G���}[���1�%��UD�ǻ¹`n5oeϥՏE�V�&�[�a�.�0	"��sܺ��r[LG���+홉t+bg�����xd�fŧJ5��J;�D2@|p�&���s��"f`�M�ty���:�Y�9q�A2�5�Q�["�,�#�s;k��*ucu�r�b���a�E�% �g$;�O�!����̖%6& ���g��mv�����z�T�zf^�ø�������w~6���U�*-�
]L��k4���Ư����gKA)xtgV�;3�Ӡ�vʦ�m$9��e�5)M�(�vs�R��uZOrˡ�^�Tq�:���\�7��d�4�_���UV��ի�ms�cH�p��û"erc��Z�N��*��>1��Muo`���z��T�θl�
�7�Q#z�9oR޽(Y���,�ƭ�)2Em�o4:��YL�Gf�ڛ��p'�T>{�Rü�r]��`^��+M[�P<'e�E��.;�����ʱ �qI����x�D����Nwܩ�BFx�̝��Z�4C��� ?_��(dp�w�����R�ټ�^�u�O�ʈ�wf�Zכ���f�m�c@�B�W����;��m���Z�*�g��%�y�D��<ۋ��m����<���b�hy&�L��Өxu����=)���V7���f�־3~��>����/!�΅�Шq��]	���N��������U�n��C�j襬<��U�[>~�Nh�.YS�v�I�Aw̎e;�fFmU�j�CuF^P=*3.�Nbʶ�5Ğ��J���]o��x�MX��&�=��d�0��0U��ۧ�nk��}ӁA�h~��K��i�e�#��C�_�5g�R�g��NUN۽WR��7B�Pam��b�nu�ne7������R>���=V��A�+���ء����6S��Ǻ�r���
��{��G�.�z����7�r4^�|j���d.�t�8�Vs���b�Xnзب����u�������ܫ˅6�:�.�\됭8
Sl:��Ύ-����X87:s)i��P��$w��t.�}A/o�n9Rd�W;ժ%Ϊ� ^�ɽJDilr�Cp#�k׈mNޭ���,&xVf�̄Z��a��{�.�e��׳Y�MƬd7G����غP�p��9���Zo:���9��)1]pR�&tH��"$Q�\�j��-r�@�Ej.�}u��jCeN��n)�Ux+�p�Π�N�Mo�j��[�^[1Pi��U�TN�_'}��%]F��|�5>��,��3,~���\/ZƊ�����%ԧn0L��D*���F�yt�=s�s��o�@0�cY�&��I���]`iv���@�/������[y�Nh��,���M!ѱr�7%ӂ����!t�%N=І���e������S
̤\�ne�W����rF|Wgf�	]�f��\嘻n��f��9	������F��g�x#{��|x�gc�k8-���Õh�Xܻ4k!a�c&ʀ��0����b/��_'c�k�!>@嫶�y˝)��}�5"��,-'v������7�T��u�8�(s�hVo=�.�pғ>��j&��;fЗc�OnP\�`�IM�pa�7��q�����u7��]`w���5�i���^Qr��4;�>R,�2u�haec뭶��[��w���.F{�6SW}nJ����ݕ�r�؞rs���aN�ce��~.������G�Ğ�Y���qf���/!����^͜{)9��nm��#��6��a�y�������.�Ƶ]G5��1WL���t5uí�u�Dfk��W�0[㎤��n�}v�H/�[ۭL�)L
�&.��������侦V�^K�)a���m�Cz��ݺu�"��=yv ��gj�L\����:2��p����B2���3w�W��?�����UU���mkZ�}��|��x`��8$�c�T��-ܻ<�+޸:�1��T�
�i���:'gv�o�Or�-��rf�:�";EF��	���y;B�V.���9L��W+ږ�7�b�v���geMp�,�ކvhm\,�]X��y������rbxtNB��7��|��z��Lw8��O��n��0�B�V�r�\l�މw�˳$�񵄯�Ng�"�JUt��Ζ�v���YV31�Pm��J����H!a�nIW!}r�M�*���	4��Mnd��1>3���%����1-���H���=�'(VK��u�K%�-g���I�=r	`�ʕ�t���A�hU��K5M'�,���.o�xnW5�1��(���Gv��Z���8�لm�b�}���h��)�N�OVF�J��Py�P�r�Pt\O�����\��ly�v,_ɢ��ok�-bvr���r��]uR��`�\��ڽ�C�:��	����؂0����!��f-��Т��R�ю�m�c
˙�>�<�G� �޳x�����ك�Jݻn�.�N
Bby���~����rq4�eՒ���ˑY�dR������ؙ9[��n�oF�U�cm�]�;P�E�D�&6I���2�7W����,��T��}�ةX#�m-xx+[�G[���
1�̀2F�Ja�zΩr��i��$n��##K/l�ƃ�O.����V4U��V�e��gq�J�-l�ѽq��#�0��`Rc�`�*r7�^#re���E�s>ʦ�Uwkݳ�������E�[��Lk�m1�޴��]X;;j�(+��i���lU��۴���N�/�7��8e��NZ�'m��o8G�3j�L[���\Aƺ���pc��4Y=*i� ܖ.cs�m����;	(U�B���׼��S7,.�%-i��n��ZD�j=åy�o*�Z-�N�i�z9:�8Js"�ܯ:LB�n���7öv���ĆD
ք������Mj�i��HS��s��������#��owq���/}Ԣ�Ȋ�Ô��+�.>�,�|nz>�J���E��hw)�aa�LT�k�E��H��6+ wǑCz�^��d1wv0�r���&Q��u��ʹ �1fnNW�5X�;��/�);.P4Nd�\[���@� ��buD�YSf�ݘ	�}�1�f��y}���J�t�I�����pU�L]�[*���5g���cai����ݢL�=Xj�n1,M��7�-����뎧rqS��u�aё�}��W�1�|	.���,��[��_�Ӫ�_��6��9e�=�E���n9�b����>;6V�K-�}hsś��3ݷ4m6�6Ѣժ��jb�L��VhU�5\� Z�k�����T.���x1�"p���Dm��{��mL�z�\��է���D����}mq��^ފ�Yy�w"��b�]��C�o�ad�V!-*<�o{j r�I:��F=�CoY�t��C�7mi��ylF�Y����s,ع���B���� �_fU�G+,Z�8)�&�Sn2����aB�w5%(��]9���qQ���אý��r�h٣�,��+���SK��dW�*]��A�ୠ����i�ރh[̴&�"r>t��X�X��;1Ԅr���Iz���T5�nXw ���9@���.��!�9o\�ѿ�9q�GRk,:l$o�� A��P��فVQ�e�ވ�\=��H_N���h^<ME�y�Ma;t�ˏ��V���PF�m�駳N�$@�5�O=�ql�ݑ4,�hzrI���*�P�+^2���L��%�`�F��\�w�h��qp�t�����yb4g�'�� ^�y򽫥�Y�[e��:���J��eQڶ���<R��t�Vb6����n�GB��r�Fky+���X�5պ)�9o,�F	 ����8�[�����;�kC[)�M�՚Փ��ƚ��_����%�!�sS1  ���W[�Ȼ��V��þ�&b��/3�2jٿZ�"�9�aB{/x�S'��lއ�#{b;ǙYg�Z�}yh�Ũ��7���e��P�(3V.�!B��tعKdZ5}��X���|L\��[o�zk����u{i��v�e�RWb�ܝL���.t�mei�Y�^0�KLE�0����f#�;st<��H����}����T�^���B�Eɻ�nyix/��1��FM��Y>ǈL�����q�)��Ҋ��6f輦�S�cVh���\:�T%�r�Տx(48��.j����-p�|&�@�g�v���ޝ�L�0�`�hZ���17�p��7ۦRb���eȔ;�ff�=�7nX-
����e
��+i��uv]�lV��m�l����%l�V��$����7ٻ��|�CF?پ��'ɏ1�{�<�/"��]\C�r�5��T� 550�kd��xV}4%�
v�RnS�Vk]
1h�d��0Μ��^�����Q�uB�$: ��n����ˉ�we]��ܵskM3��U���M�Zp��^!,Լ#�)��]Z��K�ؕj�q����c�I� ���%`��X{�B�t��,[�˼����t�bU���!��T˽�资�`��1�	��Ԁ�\q�F��ow$���7\���(�ͺ1k?v�t�5g-k�>BT�8��<�6+��R��%ۡA��3)�)�x`7Z�P������n(�Nږ-f96��Z�D��fRY�\_cٌ�df�@;����o$]敱�Ð��ň����f��͓Z�Q��ɡK���_��xy�^�T�_�m��r�%����+��\�dtx�Ia$�|c�n1K]��}N*�8�mԊuM35��`!&��7b�� ���E�ԓ�FZ�N���;�����=�,/_��{���8��;)����M-wͨq���D��m����˰�KӮ$6��p�l��:Q;Y��{W�U{�SS~�+�10�R�=���h�:��d�xI6:%e8ԃ�GY)>i��?��<���=��R�ܵ��C-qܗ�7���g����R��w� �U�d���{m���|%d����7��bWEX�qZ��ʛ\�[��J��X֚�y^�G���q�<|���d�����$��9�MMʹ.�{����A�|X�}9�#(d�$�cݚ�Z�c�e��綤[��

��{�[��4]>}d�.�h�
P��1��o���hgQ�,��Fec`Y�X(.{�~�l%9R�k5jᙙBm�܂�tD�w̗�z����\$����V�
»�V�&q���|�	J���n:��չY,���Z+�-.�	��c��Z�/�<�������{�d`�ۖ�;�+Fq�]26��-�[�����\M��5�]��C/o�l�o��>�
��]��+��;J�KkƝ��$�` ����x��7�N��v,r���.�b1W9�����M�ŵ���Ēvz�8iri��&j��!{(&���>�eAY��l�dD��w��+k;Ô��4{/5�ۭ�s6@�8�S���E��s3l�13�pӋ���7D1�ѵb�%f�(h������S<M�������>C}�o�ˏ������Q}-\C'��Z����H �0ݎ�m�?����iS�5����[�=)U���G�"��_n�ƽ��N�䭁�(��Wco����7/���uB5��T������t�A���8˜���`��tM���s�Ap"����H۾���Way������4�*:^��������D��F�3¾w�+p{I��fe�\��Z
'�9V���T޳����1s��`?iY�kKVj�ڹ�Wi[KM٨�V�1YŋF�����oj*�²�eK��ٜ�����7�}�E�n��r, '\���'m�x��呗Ʊ4�D�_+�a�Ο �ͮ�V()A�q� ��X�ꎀ��Xÿ��$;����8���r�+�&��+Ӫv�.����\����wf���n��vy�Z�h��l��Y�;	{��f��]W�"��%H��Q��%�仙S����i,��I�Ah�(�k淃��njГZZ]ۺ�繐���K/���{��Ŵ8,C{o�
�s��Đ�!��q�l�l˹�����}ʘP-����Rf�&���=2V;gy�؉Ύm~�ʄ�c�l-�Ř�ͤ\�5�&: /}+zE�����Epѩ=�q��x�'����I�K��Ʉ9�7�y@k�z�q|~�E��f� �%��$�6ȫ��v�5�X���H�	B��ڞ��ʺ|/�"�7�א=�}�~nމ�������ٓ��Â��Ք�w3 �fn�7i;�.J�r�ʐQ0�nZyN�*:G������r���uƯ�Э�F�޽���@�9����4$Jz(S����n��;��|J�LX�b�q^�J���4sb��@��}�����Xz�p�{�T9���޸Jw�_ZN�C�L�Ю���:��Z;/r�j��F��KV�����C*�6��K�to!����o���Ac�����p���Ά)���J=�M�ҽFpچ�\p��#���B"LшeɈ�� 뾁J��������u����������B=ҕ�2�ė �\K�����s�Q��y����x�
'���|�cO,G�oS��F_i�b���{`a��	8�������V��'�q_DgoVKrk�Ŝ�<ݤ�����H�k�5(J#�̹4���1^�&x�E�*N�|��^-���<��oi�����TYJ�z���t�̮ː�n籏4����ږ�i�Iλ�ƾ�W����uk0@��5)	ݕ�h�Dw��kO'j{�:8���eh��m�>�[�4�Xw	�VC��҅}+t����M��h�W��P��OLA�Qta��fsεtP,�1�������qHMx˨I�D݉���cF�w\�xM��|)F�v��{M�����G�U������/njp3*8�"�6;+S7,	cu�q�轞;�`ܣvZ�r�Y��X���
���A	�[A�O�H�x�ǭ�2d��d�ck<K��;�
~u�׆i�h��|[98�mW`��,І�h4ѻ�`*�,o���$�c/�	{�9��V�f�f�WvQgӄ����}4{�B,��sč�WN	�'�(��FUrrm���.L�t%�dq[�t�dWׅu��܍�-�p�*u����s1ŪY{�"^�^ƶ���	��Զ��(¹��y+��J��N��<���K�/��w��V1��4�v��j�n��W�wB�*�lqPOq���B�o�O��ǜ.�˩o�۰���jr*V�`έ4�Eu�4�!�]���D�/s�����jǛä�#�T�tϠ:�1��b�L	.�6
ޓ.?rHb�7����,��^޾�tH�6%��Y7}��#Y�Պ8@{j!�c.������	N75
��0Ƈ�j��AO�s��(ʮ���ps7B�ik�#�	�^�Q;w���1�����7˩��2��b$��Hg�C�޴=�3Bo%�"�������c`�)(�n���4��(���V�Rn��P�6i�i��RB.�Y�yK�wO�9����2��veem���Q�ő� /���Y��#7��Y[V�a�K��7��	]F��le�w��f��魟B6�P9��{�P��/�]Ԡ��Ӫ��4D�#N�sm7[�ﯓ7u��%����N��iK7�:���qb��*�ߍ�W�z!n���e���f�Q͘�AK8x�ʸ3����m�:�_mj�U�z�2��O.8��h^����6�i6P���%�b6T���xg�y��z��
a}{�V*�$�yӼ����=BXcS��{{!���Q�,��J������Z2���_Y�J�̽q7�ڷ;N��i��sB�b����}j��b�r�-Tɕ{vMYu.���4*7�����q9�)LE/�9m��.����gk:��gǖ�\�977:N%7Ja�-5ukV��i��y/2�1��9w%�;���eI�����a�,{d̨ͮ�.��݌`k�jx]�J=�v�uQ�kF��lJ*H$�����ju�;�[&t�w�/O�2�ܹDn�����[m���w��`#�V�eAwA���<s.�t ���,�t�*+�h[0����ƀ�X��t�r���v�x )���F\ܫ[�6fk�'9kN����ۙ��tM9,��p ��hleI5+'.�fk�l8�粒y�T~�o��:�3q�=-��˚(���p���,<�g��V/&<P')C7�����e�xþ�[F�څ�{%�c�
��{�cL�6:��c�"��[Ap��]�"��d�*�U�>��s T��8`��w���b��ڽ5t䷸�Aq����\j�պT���|���o[�U1�.�s]���H]D�6�E-5�)az���r�3���׺f���L�����V͍�|�>D>��Z6����隌�mj�;��fL�,V��,���w.��@�5+$��e͗.�nZ7�8���h�.=$`�U�ݠ��b�q���;�{vNK���������h�A�VX:�=D��c�.���#���hO6:6\�*R�[dlkjj��(����J�e����}�J:��Vc�o��`���s�(N��uj��*�^�/�:�����Ӧ�tx�ֱdy[Wa=�+C:�ٲ�
�t�(���r=s�vF�pr ���*���5�����ZG:��2T<��I��4Ψ%* �S$AG͌YJ�ΆL��aDŨ$�f���y�iX/VC]Oq���}�ԍ�C��`��C��-�{�������_���|>G�|"#X�#(���VS�H�N��DE���y"�e���7r�5Չ����7���$���*	�<����^l�[]�\d�A���{��Ǵ��{��a%��.BN)��z˹��˭�j ���`���S��� ���7N&�����{g��e�M>0'�,�Q��2��y!�];%u�v`s���2ٵb)� �\�ƀ��k(=��:�e�:��e���)<�}3a�V�aN��Z6��23(��:4;��bl]uշ+NL���x��\}�'��C������	x����{�祽��ɪ�9tݓ�ĽAb�����^$�g+K5��z��ix�4��Â�sE��f�����3^ښl�b���v�8���\�3�^,�qiwC�kB�n|_Z�5ֽ��Tr�G	���o�~���9�E��d����ۖ0��	�����+��u��w�`)�Wva�{ђ�Z�:��>5���&㶷F�����Nܰ;�SqjƖ���[l�D��0ݱz�.��&빝KK��:��e�V���Pu�Nt|M��"o�q�^����A����rOc ��es�	ݍ�2��7'Vif�A�v�\ [dqu0�_=o���1h�	�ǣ�ZU���]R�q���gfCX �����1��^��k�:�H$A
B�I)��2(��b����Ib��F��JjhFɈؒ��ؠ�wv�,�`�Lh�!Q���"DC6(�&S%%)(�	��d��Y���6�QAAX�,m0��Hh�L����"�H�1����a%�1�(�(ѱ��A��"�4b������Ɠ&j��$���6�ȓD@	�(�V����wp�`�4�wth��ALH��BR#`��\�6
�@�������r�I$ �!��`�ɨƣQ�ĄQD�5Ja�����lR�Q]ݴ0"4E�\�$�4l%b�6���> P��jlX5����#qD�+3�^C�7{�;�����F�����s'��m��i�*Ψ�T��,E�y]���&(���т�s�ຣ����|q�d4��tMp��AV�_L�����3�m���cΥ��;����ɓ Ն�������T|���q��5�/a�����i���~+��I�^e_(�׷y���n 7I�@W�� *�G�u�D�+��u-��/aN�pc2�z���3+P{�=\0ԼM}Q�`3	������(��+9%��c�]�M[�����s����s����:�z�~��3�uN���)�&1��e�5��vV�}��F]q��䣜L+�!e�'b� �@gM"}��q����1W�y5�Lm$���v{�S���^ˌ�}�-q����j�� ��`�Rr6�R��Ov���^�+��qn�GӮ�ν���ޯr�a��k�&*�kV��^�:�^�e.v�dl��;u���Ȑ�����+��4J�GK��z8]b�`S=+�|ȯN�[��=O���?d}� �����4m�#�_�&8R5�2Ẁ�^6C�>]o�P�k4����?]qA��׈��d���*�,�/��{<�3[����T���2��^JS��\�5�]��.QѲi��|����yκ�or�ƽ|S�)h�����s:��l�%u�+vp��l����͊�
�hI:��S��⩽P���Y4�SĦ�
]m�1u[gM�݅�8=X�p鼯�Q���a�=�ۗ���?5sF��q�ۉ�:�������C��=�U 竻���p�O��	��}��� ���1����S���*x���|�OԋS*n}U#n@�1��ʅ�Q�
�n�;�.1�6�آ��Ou��X�2����m�b�F��mħ}� ���m|�n�%3��� Y{5��z���]P8����U��RFGz�(i�f��N�� �;�g9՜�؊H�'4�z���]���G��Z˓��W�۲)�TH0����"���"`!�~
{t=�����;<u��t*BT��2~zzT�t}��́)r�b��}���Vpꞻ�
Ý���%�C��K]4J�9���b�꯱�@��%�&���M��$]��Ӧ��D�iNj�켛�
�ai�S��L ��l�b�fm;M�c��V�8I�E������W�pJ4�����v��{_U��
ٽ� ����S0�.si��VRs���0�v���+F_BՈE�y�� �(U�'<j�V���tPN�s��
�ʄʼg�R{�����ɘ3�)V�{bN�����6�7D=L!Bj����g�6��=}��o�O���6eI&.��l͙�4�Pnuо���M�*�;���ǪY��������&X��o�a�R8i�"6ɳ�En�my╆��*VV��{8ޗ����#�4�s�	���*���P�T�Ӓ�l`�#�?�'g���T�=W�s�P_�E}�܍�I����8��eB��}I9�;f3MCy����(�H�s`��T�o�ن(IХ�ڲJ}����.�!�Jp+2A������P�����E}��t�*�*�얼�jy�O����~��x��n ϴ�ʴ��ĸo�Y�:e����w/M«�i�=D���nnWz���g�z�5U�ҁ]�
�-�#q�?h�n�B1��L���=��,��34,��q7.a��<U�ru����4[�\��q���J��c|_V�b��;����.7���q��*zt�~V莖P�Cx䦐�u{�\C���X�u&��{�8/�.��ų!
��Q�خ�	�,d5��M�,�/�T��w.Q����2�F�zV����WZ��'=7��*�����N��)`�e=��gA�c3�(Fl��m���ۇ�,�t"����6�t���9o�vy�o��NE3K�nq�G�v�j��*)�$|xm�!����:�5s�0�U�����g�!�o��N��iW�x��)�o9͑Yd'�}dfL-�e�Ł_b �'l��S3���	C1dF%׈��:��B�����'i���2�o�2z2w;&�m��KU�귄������'���U�.��;ߧ{n�'v��uٝ62Tl�=�Or� k(cje����Xzs�ͨW��5b��]��d|7l�c]OhR�A*����s;�˄S G���6���^�T1��;=���U6���҇��AWz��D��k����ߏ��M�N�y���5�aC�]�֙�@����վ*�YST]'xf�}qc��q�F�����&;����)�t�r,;)
|.���u%�v��oMf���[`��*i.1�P� Z�!�gZ W֦��	Ύj��[ey��X�Ί=��e!�ݥ��	T\NL`�s0��@�(U��7�c�!Tl�C.4�oN�s2��z��T�4����코�RߺK��.3��|�v'�y�]>$o�I�g:g�<0yK5R#��ŝ��z�KkE�O�}����~d>������]Q)�BNy��ۮ�<jT�jR���y���ݨ:��,@N�GJ�H@�c�\�`�w,�9�]f�:qF�#9���]�|���y��p�ƨ��qG�Mz�cU�2�ī6Q��Rӳ��f���G U���U�a��9����S����Ң�)E�9M��|�w���a}{��,1�v�}ӔQ�]DE
��@-ʩR��5�T�Ƨ$B�yѹ�%��8(`u;H�CAR�~��b�'�ىH�RfY��*�1�b"�	�P�����Y����&�u�^��|xs{\T�k�j.��T'.L+���6��'FkaR�r`��6`���@�]�d!k���l`<�`
u���R����Χn�uA��?k����5��`��][�	�3/�0�N�,W�mZ5�Ů��A��k�{ݫ9Ӹ�}ʠo� �z0%%�\f�{~��H�i��o�s�Pl�J:��/21�m1ک��h�"�����T�l
i`�z?#��'�X(��IϹ����J�<&g�xVxߚ��I�iѵ�_O����N(鶪�8w o��.K�3���c�Y�H��ۋ:��4��b+zt���;�6+�����x|2���k���w�FHN��6�UA�1��e�B�	�X��5����D
����u u=��G:��w�����|=�t��;\�����A��vJ9��j�a���x���X�[�>R�۝��b��E��T0֗:��wlxcɽ���.]�Vlb�ۉ��\ǋ_u�K���m�/��v&G�|OV���%��S<$��}�Dh*��B�D�é��Y݌gIؕ�U��lo�,���lں��u���i�"cqP9gjؾ/K����oN�(K�S�e�c��b�Լ�a�t�uV�}_�C8�#�񫩰/����@��'��D�ژ�~f�.'���*����q��06/]��t���Lº��А���ҚW:��q�V���-�F4\5:�͐�_
1&Ŷ�ա��gnx�����6q�0��5W�AL�߃�wM�/�«W���F�Ɋvk\s�ǚ�к��E���-@>�v��@����R�s���K>�:��r0�y�!���Ky ʟ�D�QX�>��q�~L�*ɒ4dJTY��eB�І�u�q1<8i�ڞ�X���\�{�F�V���/J|�eu�C�X�޵��˽6͓�r��x'��c�WLuVܘ�ju*'��S����/�RD���rE��LL ��c�*u����3m�x1FVN���I�17��㯙ل6�2䗒t7�@��	���^[t��L��7�O����Z�ui�E7-o֬�����w˸�ٸ5wa���eX[����T�h>�ô&�y"F> �R�+�;�+b�v��nHF��ze��q;z����C6lFB�����v���ŃZ��v�2p�}wӰ����oind�*K�*p�z��;� 5��p�]��e��Î��P�U	S�1�g���R�����˒G���R(MbFt�\���nI�uF��Cd����t�(G�1'A��*bøF� ��Ns�c�>���;C��~�'�iaB�U�����W[R<C���;�-eg����,�lH{|�Z`Fޮ���ry��
6��x��e�uq2F��EXZ�g5T�,�p:exݔya�4��f}J�����g���������q!}Z��� X�7�8S�	Y����Q�*F��q84\�.��\e�t�������5
L���ia�����d�I�Q_I��yC�E�
�7]�g����
�o��sùZ�X.�'�(!d�;�=�q"3~�M����v;nq������~Y9i�/�{��j?B�TN8�7 _5�xKJ�8���K&��b����w,l�ԯ���.�f�7e���B�્f��+���K�@��`:�[�Z_`w�:��G{����x�����HUg�=�¨���r��d�y*g(`����$t.n�t�s3a=<q#j�҄�Ѹ����Q�$��pOoRt�tG3J��'���4�g���K�u6����6r-��{m�m%��n>,��}���d�8n"��f�e�9-��A.η~��5�j,ڮ���*MC�_a��_�s��V�3��+q�9�m���]��I��!#n������r������`r;qY�X&z
��7������H� �z��O?�w�D_uC�3���8B�c��Oe�u���ʕpZ���I��\ڊ�['�3�.�WY���U�މ��P�S�)�8�B������t@9�T
���"�+a�$����\�S�&&+��F2�f��2�1)mZ!9���o#A�溳-�)��ePvUR��/������~V��<+������.��Ķ�&UC2���OW/Ǜ��` �/ƣK�r�p{��B��rtF9�	�ن��*k\��0iX�z7yY[�5TQ��(���+f��ԫ�ϫ����5�c��V�)�iv���j`Ue���`P�2�A���4΢��bx�k�����s���Ӕ�r�K���`=�X������7�7��UTD��/����N>l֗���=��)�5y���~+c��;����۳�Y���L�v��`�<>��)�[ż8�Mn�)�x��N��v�Ze)/R�;��־�����&3T ��Ъ�B�p=���8�F��|��Ʈ�񻐳6�����Kuw<[0	��="��W�Q;<'ת��@���!��t� ^����}��#��N�No��u}
\�3KD����m���%^�Z��_�����x��yΞ�G�x�%Uԭ*j8���p��N�����tW��~���Q��}��+�$r5s,s93�o���Z��u���¸�i�F;>}L!s�Z9��!� �4��9�b��&(�S�,�;<9��3.XU�;X%��Mt�ܨWU-9��n�nX�e��T��u*�nET����$9�S���\��J����cQ��,uAc�i�F2
��S���,C����e�R�h���,?]�{OU�s���)���RHBo����1w(u^�ʔ���Ὦ*r5���Gʪ��ɰq^���t˴k=^4��V*Z;m�)��a=��|=׺xZ��O���õס#.c2Cu��� ��vd�K���_�5���1K�p�]�B5��h�H�����V���{+���A�1`���YN����>xd�������OTQ\�d�j��"�?_��Ҩ�`�)ZnV݇�༘{����&�(w[G��\����1����2�S��&x��̚�4_yPN�m}�0]C���Z{����2b��p���V�0%���I���7{@�3�]��F�nm"���s
��<�:��l�ߤ-�2{z�L<]9��6���^q�P�i2~��)��ԁ! ��d�g�.���Kv�6x��f�3�=ӷ�oL�Wf_�PU�_Nt�f*98������r��?�\��8��[�\���9���@Z���j.p1�A��m;�/y�T꯵�j��?�����)K�d'�5c�T�3 �0D!f�48����e�/
/���-O�w�<�P`�V���6��Q���Ej�Fm����]�א���?���nUO=�P�������@9�Z�j]H�j.{��=[5�~�&�.�ُ�����/���8I�~K�_U���¨��N.]�T�NVY��_-4ܡ����ض�!eN�*�	��p�]�f�#q��ތ��0�jo�2�,;-��i�cC�o�e��z�����B�kkk�� ���v��@7+����1�Ʃ�?q�;�]r�6'��߻L?��ifٌ���~�}Z��e-����U7`3^ Jz�ǝ�>����.��h��p��>ӧ6ŏ�ܫ�؈�)�]w.=�ٕ!�c���a��3e�_e���y����;��J$s�h�(��Y�Y��iG�n�RJa�N�dQĘ���x��d_m�!�M�Z��/<�FM��Dv/D�A�zgQ[\�W��wqSC�aZ�� $:�`�G�ȴ�4ú��<e�%r�X�1�d9���M�C.�Kn� ��[Ѓ÷Ŋ��KT�HɣugD;�D_A�J��5�7�*�V�øV�[a�!�7k�*�֫_f����p4��՚7:0�~��Ф���U��mա�;Q{��1�3&�+	�6��ײ������;pjj�� 3g^һ���g���ÒO�d�)�흧4�_5S5��_s��e�R�jV�X͊�]^+���D�B#f��s�=�h�<��5/OC�m�	�����j�wZGi
�r�/��cZ�P}���#:7�J�^#��������PU��c^<71���\S/��Bi	�tr⭙�+ds�`�ұ��il9]���2=:�Յ�Z��AqT2ED����&ڇm>7����,�_��pi:3�����!%o�[PZ��mb� v���N8umq�u��l�aրK�N����G�@��oG6��>�c_�Օ<�=�(�Ȉ"�E����pk̛�.x?atj�o�E�m-;���=���LU�=���YB�w<���犈�g�t���^����� ��g��u��GC������v�fU����7*뵀X]H�]�4�4�����:�8צNX,�7,���m[��X@�9�t�K
��㨨����}w�2�!�z)�۴5��7�5{Rtad�+y��Ip��;�=�ES��m�;"�L���@��=̀u*��\Pͨx�۲�$Y�9��Q�w6蝆3<�z	����i��)��+�=B`w�AW�������x;�K�@�Ð[X�&R�+[��B�W�Rd=b|�7>�]�ݰTI�Ɯ��qPl�ׇ�A�xu�����.6��xj4��G[ck���
�^^�n��

��)�v.yN�f��]�[෧��A>&ou�3��6�5��ۄ,�%�Q8zc�vX/���ضZ��{@7\ţDej�Ж%G� A�z��-���p��C�h�*n����Uγ���тV":v􄝺ء�>�1����mnfGK[�-�[�ņ/zH6��Qr��@gf\������ /tUׂRs(���{�M�à�b��Ti��x�|���ȁ�vg4jEX���M-�qѮ�GE��VqxSb��H�9Ql��f�|{$��U퍶"�����Z��=υ`$�;��G�(-{�_[��f��#M��1@�+!��fL�:�Q��i<�{ˏ�}yM"x�Vf����r�)ǲ����+ �dn=��gy� 6��n��-T{-(�:�j�:1�&��=��*�J`�C�v��[�O���q��]c�)��&{>�C��M�Amᒮfn#�\�o<N�
�>�
��3ӆ�r�3$�2E�F1&"��J�2b���愌d
M��F�d�܁� ��]ܢ�ȓ1�0�FƂ
K&wW!�bݷB.�4�Ɉ�b��$�(���r�%�7R0�gu�f��"
,f�aH�۪J�(4AcL�,h
2I��CQJQ��*)E�h"J1��QF�#E�II�
-�*D(��RD�d�h��AI��L幍2c���Bm�ѣ`�IQi1Y9���K�ō�bR�� E�C0F $(���*(�O���	��$��Ez�V�z���k�,�pFz$|�J}X��&_9�{��X�,su������B�[��B�/z�����QzR�?�)~�׵���}y���-����d�����ϊ��Tr�����]zU�sW����*�r�-¿Z��_~~x�KO���z�ކ�[�|\��z�}[���>�DG��q�/��N�>V�[�ވ"9^���}��1o�s~6�_=y��鼶����:����o���Ǎy\�ǁW�� �5�~�/~�W���{^���}^��o��nW7�|o
�W���� ���9�{!�	2Eנ{6���>>���yZ{���ו��o�x�k�ߊ�������ǵ\���p��׊���\����\��xW7����zW�}^���8�ʊ������׶�j5�y�"�����4}��
�l�O6�}�z4DS^^�_���v�����z���|^��ׯ�~�+|W5|��ǟ}W��^�Z�������ۛ������ͽ*�\������7��no;�r����x����������@qT|�coE�w�{g����_�nl{\�6��5=��U����?��+���W����u�h����������~_|��-���ߟ�6��Tr��|{�^�r���yo��DH�� ��΃���s�>�h�*{�_�����}����\�+�{�;z�nU�z�~|WŹ����w[��~-�{����x[��������]�¾-޿��Ms��ѽ�Ͼ6�o��>�DX�4}#� �s���dd��hnC7�����>���7z~" ���1���_o=o�_¿W�>�^׵������U�~+�������}��+����y[�\�<�מ�_5����yDA��A��C�,�" �Zކ���J��-�/�QHU!HX��ي���(���|z��5�~x�y��������}x�J����߫�����h��x{��}_���o^�����z�����"#���6"!�#�����}O�l�e�9>�%���#�B������oչn~|�-�\�x�>x�kxU��z���[ys~�����y^~�����>di��!���0��G����0R������1U����[U%ߪl����4n�`�����P�>c��=�x~*9_���/����6�׋��{o���<zZ
�k����ߚ��kG�{�|�y���6���וy[����?|�^U��~�/�o����Q�{q�h����8u�{Vk�@M.#��u^]�呁���e�+��Hg\���]ٮ�㵀h��BI� ֌�� �27��Պ�/m.F��[*ʽ�׮k⻂w�0�X̌���@i_]�
R�,��]�U���� ���l	�VE���w�T����}v��;�?�����"���U��b�} ~���.[��o����}k��������U����7�}^W�ޗ���5�_��_/�|���h�����x_���������D|��j��{|�������*��=/���������W��o:�����+������6�kUC|�}�����c�}�퇓��������X��o�ǔo�䳉{R̿1�~�G߿|m������|[��|^�����W�͹����~���W����k�yWŹ�o
��s�}k����{�����^W{��/���sz�>�������bD}S�ږn��mY^��6�0G�D�ﶞTb1�B> <���b�} }��/�?�����⼭%����G�G/��/����+�_^��+�o����k�:����|x����|4H�٥���Jz��O�>� }�>#��}��yW���_�~~��{U�r����W�}�U����E�_R^������Ǖ^�}�yo��r���Z<��㯋��s^m���|k�������[����N���-�1������zW��=�������Ͼw�����6��ݼ?����o�|T^��_�����m�W���~}��^�*�/W����|�ڼ=��xW�/��z?}C�|D@�<!u:�r-)w�g�^�~|}�/;oM���[�]���o�����R�P�R<G�����!d}�"�^���U.[�~}�9����DP�>���}c�,G�"!�;���>��|G�C{�_t�'�ks����_�+�����k��W��*�~���o�o����W�����~�l[���!"����>�w6��f(G�̪���>���~_z�o�7���w��$DD����r�QY���SU\�(�Dr��
�r�y��c�~��xkߏ�7/+F������xW�����ּ��nom|^�n~/��wkʯ����O�k���~o�<_��{�^���V������ۏH��	zhxU���9��@o�ܹoo���%�����ם|^W���޼�x��_U��5��y�K�Ѿ+�o�^+�^��������yW��_���r���_�ʯ�������P��UW��,���ӯS�0�fK�,�z���㔶��t���0����y���nv
�K �lΚܤ�4	���/��"�S��Ԫwo..-Y�Wp�ح;|Ⱦ���vFs/�ҝIL�=��>�-er�Q.�\��C� 
\��_~~��Ms\�����+�ܯ�}^�xnm����Ϛ���m�{�^|W�����o��{��W+�_��~�~/��h�������W�ᷯ��߈��DC�W3�Og=>��
>��	Bx_o߾/��^�~�k��ז�ߏ�xU��|\ۛ��[�~��oJ����~w��:��^����m���ׯ��^�}\�6�xx��[��߷������DCu&�zl�_�2��p�>����R��W߽Ίw�m��y^��U�jJ��(x}b>�<#��1B�Gb"DD[�_^��|W���ǋy\��}��^��+¯{���v�+��Ż���UȈ�#�4FӇ}G�{L�Ut���a{����r��߽^{��}oUＷ�n�ߍ^�:���u_��*�[��n\�����Š����>����+G?�z�/��?���ՙ�#H���3��@d">�+=��']��8���G�D5�^��y�������h��彯k���m�W��j�ׁ�W7��o���5�ϝ��^��nW�~��x����͹���ʽ���~���/�|[�ߪ�~���߭zVA;�:���}a��G�o?�"���?C��>e����~���5�m��o����z^?_�MxU�sz�ז������_���-��o���ו�����~{�~z���������ضw׎����_t��w��"D�`���}��+ү���o~x�5�W%~�|EA��*�+|�����L}�'�7�����~�{��jKǮ�����|W��W�+�|W�^���yj���o�&%���alٽյPD#� �����k��W�x[����y|WּH��<@���:?=�)�� B '�DP�#�[ꈱ�6X��u6">-��|<��]W��m˗��W�о� ��먮�P��u��Pp��h�K_z�\��U�y_��|o��h��u���^�����-��_��^>}�k��\�|��*�\�����y^}�Y� �ޠS7���2EߖH�,�m�w�ɪ�h�u�j�����i�F3悥�#O�s�˓,Ӷ���[]Jkʗ����j�����{}��j��J�:��V�p�h���6�ٽ��.ú淃WL�>��ފ��<��:b"q���!�Ǖ�H�Ȕ/7pwp���	*u�F��u"%rq��v(��:��C��K&ٓv��W�\���`y�S�a�_ꤐ�/x���	g��ݟu���O7�����}w,����Rq�78��?C��p��#Q��)� OA+�d�;��WS8)�!����*d�}��|��X~����\� �\����=�Q�F�UӰ�����ׅ剄!�ڒ��u�6�	�������AE ;by`Z�RK��K ��l�G��E;��&���o����>���\&s�͛���9/h���
���w�O°@��r����2�\bl��/!&V�-�p�,i�ߴ�:�T+��:`3����tO5@O�O�,ǐT=Oy��wgW�
�ٞ�mP�g΢��O<����~��+��S���ͷ46�y�[&M4�����#��6$G90�YzP��}�X�Q(2��)�P�)��ɝ����y �)�}�9-W��BV{-8��zVT>�GB c�`B�׆�QW�B��Úv�;���
pOܮg(�Z4��QC++o�1���S�%�ب�g�lj*6��a��k�p!����ٯQw$DX��:���KƒΫ��u�^�Hu���Vp�I����j{���P`X��TR+oW�����{�G̊�jt���4I%�B�u�[�ts���Y���mtq�Y��U����G�v���@8c&��F��X�0��?_���O�]�A ,P=3�_���+vZ q+ܛ~k�y���q�َ�7��	_�Xvm�L�;nc�D#|c��"x�
�í=JC�hW;*H�B����2._/&c��?.�)�k���d�xy���?>��΅�l�7N,ű6hG7�r��6�@���S�µ�X�+Wl�}���2e�/�M�z��6 �u�?��W���,���T�),Ɔ�#*U�hB�9\�Ӭ�X�ʍ��̭�.���%P\`u^���U�5b�z�W̡.��6Oq� Ŕ���c�oR�����X*0��su��t���*�$/�����F�^>
���4vy�ؓ��o;Õ����9�0�>����r��B��\��{@u�yd<��#� \utѹ��2��-(� ��*$?����783AC+��¸�N�b�g��D����&�(�"���&(g^�h��Gkh���1�&+�>�V<���1��c����ަO
!�TBN�1���d�J���r���uuDF��\���ɗBMpq�;��SF+���Oh�
{�%m�[��6\��u5�˅��C���}���e46aщ��5����K��\���Cy�Ì]���L�t����s����2^�x��q��U��V. ��C����S?W�}�}X�9�}=�>K�0M]��es^�I��ʫR�t�^���p�����_-pO{���떧N,"/����y!^�P�����<��y��]f}�k����3����j�rFq�S,r�Q':� 	��9�@lj����!2E��q'LS�#��(^�m�1�3�¸����
�zOoX��©A�ī[Q����F*��RX�*�:#D�j�N��q84u-׊���o64�1��>��yT��0Ӫ�����ꦾ�.g!����}���ٹ窔���c�c,.'2��T�a�Q6��L�+9U��l�b��d9���N��I��y�e<�q]P��u�?_�	o7N ����J�?�\7׏��Z���e�I�*B\�dv�l����B��p��M,9VJ��|���_J�s��z2g�
*�4&�(E6o��ae�mʸC>��cw]!���\0,�/�f`>P�ƚ?b=ƅ����i�S|ZU{�[VI�U=Y0����$rI��F8��Zr������Qȑ���3����V�۾�X§V�Uٴ�Km�R��/t�a�k�%��J�У��W�/�0]D��6vESUK�tf]ݽ�P�bw�ԧ��%�k��e�<��JW+Ml9���aI�M�����__j��U6�ڲ����_����}�M5C�.V��1s5�/��L.�:_M� ƓXS�!7�n���;O<��[�����ŇR��JoUp�-�PWx��X=+��S�8��!(�|�v�I��%�8j�H�Z!���M��bF}�Xݺ��[5�^���A?.����n����ʙ�1yg�_Ծ��t-�'Wd�Bܝ'�9&�9��0rg+�6�ޮ�]:������5@>
dc=�0���/Ƨ�/�-��7Yx�^?#B�����j�.{��X��ؐ\l�a����>钎 ��7U��YF��q0�\D��T�8v;j��w��b���3��oRڬ5F�yץ^��@�IԣO؝��r	�ig:�R5a�U(n���r�_�,B��pVdc��(3;�ۘ
^��yQWϯ�B�S9�F������pÅ�C�}RE^�\"���*����_ /�cC�7' *��z`AX�j<+��lT��[�!}ܲ�vB[e�d�;.c
�}��W3��9F̄2�����0w7������y̩�d#��b��]V�rBڸf[]��]1��D^H1'�_#�`��.���Z����b�-�n]>K	��5�(���P�B�.��,���KB�_}e�Y�>ٟN�r���x,Tg�J�;D�Z��i�����������}�}��| Em^C�Q�]:��+��=�\;T�R�$Ŏg�u�k��p�W�y�V-b+p�����c-�nS1��������!��O@�H@2�w��˾Ib�(��?͕KD�����U>[\c����ct�r�QJ�Hϻf��]DC�x"�V��Oyy_-���w��.�iQs1xP���|��F1�K�q��	����4�ṣ7��J}�EV#��ʗx��^RHGIo�ٺ�ʼ$��s��{N�z֞Mn���w�A5`�l��N~.���+�H_A�U�9�۪m
��Q=������	�{#�$�=P�Gи.Ŕ!�q���t�O��!��U?��=�UDo�];
�>ט@�	�ڵI����&l��ux��6�����N�l�����+M����"=�z����u�!��C���֯
S%�9Ǹ�3��xp��@4rN #��i�9��꘍k/:5v�������`YA7�����5���5�iAҡ_Nt�f*#��:n����6λ�Q�v�"΄Q˰�+���Y|�.�>t�]�1�h�8�p�/34��4FtY�d�C����)�r�����W=�j=h�����NoU��-�Ғ�w4��X���,��;&��7�+V���2o���]���C�VG��WB(veې}��}��}��N�Sֆ;ȟ�H�jy�����g�k�k);����ʈ��L��bv�fWcZiL�
�܋��m-
�a��
�m[��a�>���G>��-O���I����%�)n�^\o�W~~ڱ��s�Wz˱7�^�^B�JX���Q��� [T�x�V\�r���5: �n���u�'�Me𡑸'�ۺ����xs��O�ӾѐQ���1���#c��E@h�^|���ax���_7(h�}�x�ض��*p`=-�<�m���};�@n�F�����9�!"tv5��Wja
��2��p|<�5�s�f�W�u��� ��=��Q��SY�C�xm�Z=���»���p����*5,��uy��-��/��+�?C+��;n��5\ T�o�4����_\��F�#��%AE�e�'�e3f�DYNᎃ�W��~l�.ˊ�+�J�����]�Surp�=T�R�uB*(`n���BbPC�������
i٪�ā����,���״];�0q�ʟs$�$���v�I�E�t�G^�{�[�?0�nj��p�����U�5:�,
��{A��=��AQa�Y����������󉦇	z�*��=<Kr�=iXa���Zv�8�m`�V�!=�{ ����#��Sl$8�3'{�_p��뇑3����n��惒-He
���A{�Y��X�be���ў+4��{�����S��&�r{�{@swDkʨ� �2��)æԣ)S� 	E?�e��˒$p�?c/o��5�P�X�;s |�=t�3�ύ�+�\aӾ~�����u� 5���)WK�V:G<%�d�t50+���}$隊Ils��l�a�k鲼d�u���#�8SH\5�V��k�S��L �9���2���z�]��C�{Tt����=9�R�5��'�k�0򸆼����V�S���3K�z�e��-������S0���L7�9�E'$`�q'LW�d��NJ��*�Wn�)��ot��Y��o�5W�֕*#��21*�B�L�l<����F���{ �$T۹w��x B�'g%ZYʥg!��U�y��3������mW���"���N�n��:x�uџCw�MAw|�݃�xL�T��J�˙|Vtȍ��M���zs� ET�e��1���9}ʎ�����.=�T���:��ؠ	 ��dPh��-ԓP�L�q|�n�m�۬|�7˦K( h�Y�m��J��Z�=o�Ǭh�l�I@a�7[���*��t������ir��/A��������S����.�4f��Q��;6��{f��x�E�����}���yS��J��*���J'q띖��C��&�:	��S���xu�+��s��=-�) �O]��ʳt;��!��$fl\;9#�zϟoE�	���u��B/C�LQ�>�ֹ������*�B8E��	�Hp�4�Y�Ӹ:�'Tyn�tWd�}Ұ�����z�d����%���z��0����ԉOe��i��p���4���Z����L�̹�����<��AWH���gs®r���'v���Y@�o^ņ[ƹ+wE����Y���w1��v���&T�w;N(�q�[�J$d˨�H��}�*���ۨЩr�w�oS:,#��iC��Q��qQ�WY˜�/���T�v���'{32�퍐�-�g7s6�9��8�u�m9FL�v2�5����|��W'���M��ź�LuI�ݗf���V� �J�ǔ]�� 뵾�q��6�}��ZH�a��y��c�&�lNY��� ��%�x�L|�_h<Ee.�p7�F��(��d�jP/��glK�⩋���U�5���\"���]��D_9��W�-0�e>����i�ɿm�ris��Gk;;e5��<�9w�kkz��gpl���V/[vMX�`@�f�ٰ3F���D����}WtK ��:r>RQ�ؙ|L���e�|���E���/`N�'���7R�{,g�gn.���
9J������|_����R]����C����ӑ��v�2uA��Q�{��k}	��շή-�g2�dN�rL��ɂ#���Z���Λ}!��з�.g��E���S/�<�Wu���v^�8��}�D�ޛD"�����Z�{���խs���G�Pr�{��-���V��-�*��1�no�NVwZo�.0��,�Y����Ջ���FQ&A�5�[�p�79�3pp��v �ڻ�P�I�GMݸ8���Ì�]c _��H�ֻ���W�?>�����-=K!2	��,Mc㘱VBn�Lw�YZL�|�ܨƐ�����wp�;�a��]B9����5�X�8�l������V����8{ڢ��O	Bt,�ܝQi�m�"�n�kf����v4F�k׋�kŸ�5���a�jOW��[������}y�ԭ��}7i;��;k����Se�����s�w�:��6�H�������rk"pn�a�i�-��2��'F����h��OU�Ѻ�6�w=x����V{�Cm��{��1Z�����tY{�19.�5`Xt�u�v5n�r�U��Q��OK�Y%<z-
����/F(����W2IQ�`�4U����ƹ�REE*(��*4��6H�hѣb6v�E��L��PF���sE���F�ŋ\�JExW�����*(�D�F�،a4h�A�*��5����"Ѣ��r�@m������m�KJ`Ԛ1h�\�*�E�#<v�[<unF�lF-�FH��LE�.�C6����J64%��nr-sb���D��A
����
���V������nq)�m�r��`*�uX�v�N[�ƽ�
��b� D�Y�խ������y�M͍��o��>����lf��4n��S�����0a�!h����(�(Y0�������Iﺐr��CKv���+V4?��|bC�Uބ01�Х3���/���`?���Aq���-L�s�C
~��6���]G��cw5�%/G^V�8��rg�@�R���CM9�h�V<[�̒���=YP����~R��[$G3f�Å]L[��!` w�E98x�)���E*�y�)}G�b��3w/�}}�
��|n��\c������6-/��&=�󷏻e�j3�M��R�أ"����5psٶC���)���T��X�3X�rR���<8��S�a����y.��ab~�sd��ډ�Ú
F��6�f&O��8�/���;��.L�V
65׽>��G�(JZǵm�'%vb������!��#f0�;=�`!\d���i�B;Â#a9���v6N|,�L�F.	c��5V�ڄQ��ȏ��I�qAw�0z�*]YR��[�%����a��+�G_�0�_���o��Դ�xu���b}s�݋ܩ�x�`w��Sf�ue^ueC3�m��rz�.��^��Ӟ�A�G|��������̦��ł�t�T��d�Ce�;}�r�-�XV�d�����٬�Դs�Ձ5rnu0M�
��������i�r0�뾣l�7X�ѧ�2tD\l��qY�z�0t�?k�o�Cˏ���wV�3=OŢiT xY��_ׯ�qXveU��4�
������]O��%bt�F#����jاӀኄ������3e�b�"��tv� Z�kVЇ֐yˆʾf�
�<����#�b��.K�DP�٘\jQB��q��r"��D��&�����x�֝ncF(wX6�����z6곙|�5+��λ��Ӂ\wR���<��1��Id�	'�Ζ��r���t�T�gO��,��%#(R�V���t.w�\a�;R����`{΢&(�z~�Օ
㊥�4C���"�M;c>����g,�U�ꭋ��ٯ��3��M����:��{�\aC�4�#r��#O��<!��a�V[ˮ�,���;[��2�i$i<�Y����:����0��2y���Z���U���� m�1�L.�1-0x-�" ���%q�����^�Cft�˕���}��g\��(���_�'9{[���/b`�؋{���%�l��Lbf��E�8o0�)PO.��p.��b�.�-F�<=n��]���W��Z��q��_���G�3f�������#��vP�R"�E��_W�U[���V�_�u��[HC���@UmdP.T�{��-6��j�aR}��zL��L�N�rp�<��f8"_	B�ڴr�1�
 �o,
Yn������1�A��њĖ�l-�]v��+�&��<>l2�#�u�9��6-w���!qD�gQ 㜛��z��8�=���3��/�"�*�)f�}���a��O{������TRUY���;yˍ���~��/�lL�1��ª�[倧���x^s���y���� 5�X���n_���Ysf9�4Äp���P�	B²��xQb�T��J�s�6%�șX�g"��րΘП�˟ ��Yv7�V�>"�X���6+\��K7c�\��;g>)+�^�ﺰ�P9�gk!����
�E}���Ug�����z�.�4�Jš�4��ȸ��9��]� ��Ө�.C|�(�œ!	�]*صт�܉Z)�8���X�m�;ɝ?W�a��4�*�e�l�p/��h�Zb�J�E����<�f�K�C J�5�
'f��9�q���Gv�w2+�v��nzD��O=��V�Pr�:!VX{,[c;c�0ƣ�|*�����GOsX��+;3����ܕ"���ĉ��]oT/7�Մ55ܚ��.>N�S�#���q�}�W�G�ik7C*���@�߾�@W�YHA��`/��!��<%ZU���>�x�*�A�q�{'m��9��WrS��gP��o��`����������p=\��F�4���L���j�̎�c;7��Y��=�r d�v�Ν
��?w���Ĉ��s�`��b7y)�jr�>@A����T�"�pA}n`���xJ�q�U��L�7�|�=���&bt=kFwko�>{�^��϶��p^V��݁�*-�P��$W:,�L!�A�\���v����6>1��s|wN��>��OT!�)�f��CR0�7N�Զ�ͪ��+�u�Ӏ�g�&鈽$Bg�R���t����;sg�ė��G�s��RP5��0��~d	��Z0�+�պ�΢��]U��
�cַ�\˯8�-���D�SZ&cR��.~�Kn M�4��Ih�M���k��W���X
+��Q� ϖ{��,H��:�����'i��Z�5�k�<m̞9�;P��=���9�tg����ĉ��pmӵKk(x���tB!�N��r�\8qvm��=�7���3wI�=���^*���nVN���.O��?7�y��~V\�i���2��Kےj�Ok}k� �g�v��p)�9�V����`h�_������Jj6u.q�Q����mpD��BUP���S��+vh\7:4Z�:a�GY�'RI컆N�ϙ
�!���ع5�5W��P�[�A��E�_h���*���v�o^�}�Y���g�,�c����V�yVqkcO�*�V@ⓞ���qR�
��������K����>YE����F�튦:�ɊU��7�L�+>�Q��?9�ӫ���!��ў���P�}�}�E�����&�);Ve���,�9����zM�A�K�ֶ��Zx8ٞ/E>1��5
��!�aLkr%O*�����2�"��<��'?��w9��;h��f~��F�Q�։cw]!�K��.#�(���`%5��]�t���:��N/k�\�w�g,����ҫ6�#W�_TBN�9��"9�N+E�*B��A
6�*�%��l>�V Z/�`.;Tȉ�._�s7d�5{¡Y���s!�#J����\�NV8�J$m��c�|%r�\�j��n�O�xX��٩B�yV������Q>o��t{������W��]H��f�����݅ۤrB5�j�b;��Er�=|dN�z��6�R�R,�o��Tj�N�yі����Go }z���{�VIf�)�/r\d�����s�n�V 0�b
����E�kpNb��hË9�������0'�=��*V���UV��%�Z~d��q��}|Y5c���̣�{3���
���e�;[Ç
���n8̯yyO����������jۤ�����b��;���.��W��ޣQ��D\���)Ж4!3��dT5���>Mw�/ˢ��N̶��u�y�53��F��W��b��ʥ��E�f�`��a�YF���&������BާҥT��̘я2�,;9;Pff��16]C�3�����p6O˰�ap�}�æ�D�gn>2�9��Ͻ�V�4[V�.Z�u�fU��>��rUNn�g��'fҋ�9�o�I�^��gyg�hVjz������DU��vxO�ʘ� N�Ƈ��*��T��=���Z;Glapa�0��9��5�ñ���^%i��\�뉘Vhu+��Ok:8�P2SO�	�T4os���c1�!�󫿲�ǻ��Arh�:Wԡ�t�3u�^�s�I�2������%�x�j_*��7�f;!�1��_^������C��դ��s�E�c�W˽]$3�]
���.,f��5�Ƶa�a�QEn�.C!�� /w6��{�x�x����jѷC��yt�l�������TM���{��f�ġw��ӭ�8:�{���K�n.cK��Z�u$6�����O)كjP����G�|^�l���jEi�D�|�����YP�+B�;�׏�.Rz�<;�WǦ�_�@��,���u4���Ц6{���K� ꢭ�(u0:��i�h*\r����Ә�5����4�;G)�C#f%#{*������;f�*�p�U1��wx�9R�A�r�Ҟ�>��r0z�{g-&�q�b$�L�Yf�ɉЖUH�'C�q�1�Bwz=ɘ���h:�J�@�������,h<�`�Ǚ
�h�4CS�rH�ӟV	�3��"�*�^A�i��UV�0�e��B5��%�h�)�b�H�[9@-s l����ޝ��3c5<�^���<�:��l����� E B��f��tG>��R4 Q�����q�ն�-�
��*�X*ǂg����΢���)`�����0����?%B����Z&�Z6�,�q�(
J~i�/����*��!k�k��m;�:Ddo%�X����/���Q��i���8b��v�V�j�pp�
�a����F��O;u�2t��0O�mv����t�Y̩��;Ꞗ�7k�ڴ���Q3_E������{��TCd'��:|��x���Om|@�e���*�]���2�/�E�G
w��,W�����U���8h������G�f�k�T�S��䱧�.�Vjx���T�������V��}U_W�5^��+����Zv@$��~�0�U��<5���=��t��~7�B����J��͙O�?>��6����� Fڐ8r8��Cw�*!�z�}���oYx0�X���m	,������ 2�H��U��j0�� ���`W�&ןCW�q�e�=�<sOn�&Fm�J�mCP3u�!���������u���z�Di���-�g��5�7������[�����|G��!��*�`&�Hq{O	iV�^��V�L�۴�G[�в�[��Yݗ�W�Sh��a�ĺ-J�L�S5�̪ͤ!�9&�ڦ�F���L�P9O	wz�p���ΕCp*�@�	J��j�`)H.�IXJ�a6ű���N�ڄ��40��q�LJc X�i�3p��v�[2�Z������*�H]!�'r�����Dm|��Y��_˪!��+� �O���*f4]e�^������;�__����G_�VT�h�d��+����6�����u������.�,R��Loi��׺�[U�*S˫̩p1�ٲ3vpY�F�Q�s��8!��.Vj�,�,Ghi
Ox��6.�Tw�^uх���������M4�'M!�1��v�����g��.��3r����w ��}���m��mvB�}_W�W��������ɂ��0�/-����"B��W��r��oXuγ�z�o��8�6��`�%�vK���q:noh	���d	K�hȓ�*�X�U�"��+g��X���G�4�1P���J<�N1��d�g���jr}rԳJ�a��]��X�ͤ�u�2����a�F����|����+�zG��G��/m����+"w�k��췦zԯB�~o&0W�R;7H"Ya)�`b������W�=X��E�`��1��1�����.�tD[;�iP3��3Kȿ���V,y�Jr(���Q�l�<��_�Hv�  ڷX:Μ�9 ��e�[�ymʯh���v�V3�Om��UĞM&�E�k�o���<a��v�K�e�c��_i{O^�+zwk/��5\l,B�F�"��p���v��S�Q���G����&���1�m;�b�����i��S��[���~��^>}��
k��t�ڈn%W�z�]���z�th��=jъ��lK�zwϞ�1�o���v�8y�p�(k�N��/��*P��2hE(#z�N��M�7ݚ�u�!��#�:��o)��M;vx$�;��r���^xWF�s[YJ%�m��'b�35����̘S�xv�;)˷	5��K�3�������N��l2mG��,����Di]�Cݸ�ck�v�hK��������凉OD��H���I�7�kqRM+�ù\c���t��V�>�4\Z��URz�u�7��0������s�{;����MpB�Tn9ǩ��1R���$n*�F���`��"�jW`�ח�]�p��u����&k�+=�_r���w
��\�A�]A���~��5��:ؿ��m�׺��N�c��:d#z���'֡���5��ճy��Yx�sE���+��]�<�bc���y��ɁLg1\�=��75l���ۆ/g��e(Wi:��p`U�y���b�g���TFt�K�a�4�u��׎��w���u�~���'^lfg�"�r��^qA�n�ΜQp��ګ��I���9�e=Z�{ҭ���qZ�G϶�ĺ������ߖ�G��2�l8��Lr�G�N�7���wF�O;s�s��f2��cڣ7�=z[6k"ǋ��	��,:]b�Ո�Yۏk��:b#"n��`���ݚ�u���J���#�GC�F�����go�'[�$��þ1���k�F�o%'8�`�z��ܨ^F��r�4%��¦%(�d��;:��뗬̺��J�;cG��{Q��u�wBu��ī�tE��LHf�;�-�^�ᛗ{Y��W'X\��O.V���G��HP$�<�ȏr���o�PÕK�a������A�VA�ݤ^j��*)hU�K�`���f�5֧	�7$�ms�Vy,1ʽ���s�-�rui����A����mWSC� a��Qʾ�G��of�,�ޢxI9�|�.������fpIs�������wG&r�5Vs��ޕ�tC��qȨ��y���cU�wA����r�	f��kƞ��o<X^�[�θ����&T3-qXp�Π�/-��1Q�� \���YKlI����x��uk]��R���YĶMc{���kBY�'�91���+��S_K��˱W�3�N�7��ڌkpDm�󝎴3j�	��@�\�,�|�����m���U�����Y�{���$���ʲ�簾]O�4��=�kطd�:�0Ԙ�_e���#�s0��[d���LS�J˜�p�ax�<[�2�9�w���)�Q����E�v*FjW5�{qP�I\�������-�/4%� �F�>89�}��D/�R�e� ��&N�56�ٲ�Lv\��G
���;�4��X�P����5�&*z�A�V�;Tl"�e�{!c0����]v��`:���=O��dr� 9,�I�)�}��eGS A��<��Z�f����b�#��u��z�ҽ���ݓ�I��fm[da�oR�������ݽ:G����vf D<N�&��O��{���%ѧؗ=�A|Գ�b�⻬�]b���� Nڄ�����6��gc4+�>[Y?X��J��g��r��!륕y��Nul��A\��RO��έ-@�� ��$�.ڭ�\e��R�7kv=|�rc|A
S�c��zm�i�J�{���A��O��#�Bu�����,oGL�M�ؕ�R��Q��(
m]�7�<d�u��E�]B���z�'�F*���9P�0J/��oY��5�@mgf�������@�%h���:/:h+5�<�.�lR+,/n��s�Y]�8���n�|낊"Fn��'7e�g�J�·���;�r�4�ĞY��t��,�F6�MpEW����.�K�h�9�)X��@g]��d:�.�5j�Nz�)�Q�������#�͜�V�Ր�I����R��lg �c_G����⦟wpy�V�X������O����W*�ʌ&��lmTX�A�4h�!bۻ�H%ckr��&#ưh�c\�6��5����Q�#`cF�ncZ0��Ѷ��j�s�6M�.���f���
ōF�X��s��ф�Qb�lj���A�ZM�F(�5%�nb6,h�
"(�*�(7������e��߽	�hI�
��d��i�ݑ��A�{��P=��6�2�V��*�{*MI. mٗr>�yťw� �睊E�d��)<w�����p��i�$���l�QP�q�8�O��.��o�]`��X㱙ש��j/J�Ϣb��)�}[���XV�v;bU�E�-��:St����U����25�Jr������/*57��/w�U^)����n9��ξ޹s4�=sA��OV�Q��TGO����<�&�"��S[��.�+u�[�x��>q���4�6���Sg��C�}Y�;~�);�V�4��Z�o%<y���la���Z�zT��[P�*��ܚ��Mw57�i�j�SJpbT�lL[�:���oT�7/����{~��q�
����f�ܞ}v;��P�Tc%����ǡn��2��ox+��T�r��tF�L��=faUJ�>ʹW�ڃy�x��_-n�9�!��B��q�nF�jI�V�g<� �;ou�wٳ.��ݙ
�5�)m$-��VGSwK��hCC�u	oʻ+�vPp�B�o��tǁ7{d���Ү4��*�
-�a�<,ʏҹŘhOi칝��cN��M`cܭH xs[J��3NC.u�^k��be����qeMLf�A��R�<q�i�=5*��dj;����9V\ཀྵ�>��/1	y�M���&V71y:�k:�bt��>������z�Ȝ^��m�XS]�c=��c:���*�N	�aZ�;�Q�oz���Y��T�Z�̼U��3�ذO":B�ΐ�
�*V+��u�*�o�џ���%�y/+uA�A��iT_urk�z\���q	3����=������ώ+��ު���\ml��5����dc�2Qq��Lw,qq���{�5	�ʎxwmȼ�8��U��/NN�_.����W�ы\^F≮X�q�޿�˂v�O{�&1l�2o��R�sռ�9y1s�Qgb�U��B�
�k�{��ȱ]x���O���|3��n;�����jkUqU���7��[�m>oO�Z�.�;�wD�]�s���n=ϓ�k` �������S�W;�V��<�RU����XE9��of����w���6q�������V7��Η��-N��=���:��vEnFL[H�6�\��t;���w-�V߱R��.�-$r�n\��fyjg.�#�j�mA���N>t/��wXV����HK�(�Z�ܞ>o�](d��ê� Pt��Sx�	 :%<w��lm��^E�0�]d�9�j���[���}UUQ�8�pC�'}��Q�RY�v�d�t�\GL%L�n�*N�S��L.�Vf��R���7Wv.�Ĕ���jX�&Қ��xa-�NF	���˪��A���N$ܜn���.�19��UB�n�[�g��[�!�8���	�/z��t�a�N���������s�5W葾8����:��	Z!�X���z����`���Oe��.T�ܔ}=���m;�n�|BҦ�<�}|�.�8�����/U�Ԇ�w*�e�쭡=�f�4���ڷ'';���ӂOoTʇ�}���F�rp��ƅA�h�r�A�y�^*=P��g��ke��k8��6��N@�g.�y�(�LmD78�5Z�u�q�w�`��O&Ϻ7+�'}�B�T��mj��Mީ��U=̚OwY�fc!�y�t�s޽ʾ���8��ŵX�Dj��.�w�n�|g����q�E��[.o'�tj���<ǉ��\f!0�P]���w��T�T��Z{��co/
��0�AN�ę��g]�1z�:$׷k�m׫���y�Iy��"�,�&����K}�� ���JU��߽��6�w ����9��*���F*���5B ��I]�2xB{袗P_�z�t��E�jޞC���W��f���=:�'g��x4;�����[���#�Ɩ_�S��v��Mv_����%TAV���3����@�뛾RR���6�3X��):E���Ό�A�*өn�H6�^���eu��w\�Y�mh]��q�mM�q���A�ڗ�&�X��ץ��Sf�nz��w�
�[#����JHGFf�Yq�^m����݋h0w��ٹr�߾�ۣ�}�������+�>��{�$5@�tVj�չ���g�7�:��fa\��k��-��bV���2/\���
]ApG��k���c	�]EؤY�-��C�z%nNU�ґ�K�뭝���Nc�e�>
b�W�NQ��/��T�;^܅>�I攕7̷�gX�f�l	�4+.��v���<��[�׳(���'%�o��q&�|(s�<�]0�j�۵ =�ε�JL��R!��v���^</��~���'���'*֎�2�l���Pύ�Z��)�3҆�]5�ڲ�s7�r~O
��9�����r�W�VYƹ���O��U}��b���v�>v����5�'�,�'>���M-�	���emTMe8�X+Z��c�?��nU����X'�uR�!�bp6��j�f4�Z0��w1t->*M����T��g��c��$��b�]���?<o8ڊ=��,n���C	��[u5�.?Cmm{.-��>(����P[�ެ�m��N�˩���N�zs��,^�y������_Үb�[�a�k5���'E5]"z1���,=�,{6���'�my����TԎ7����xVi���7��O*��9TiY����q�ͨ�km����c�Q6��3��m ��D��#������E�ue����P�g����{�]_*)*}�
���Sy�kEs��y6nӽ�TYK���c��~H�b�M�'B�㌑<x(�sJ�M'h�[p�*��P��ML|R��jmj�x�p�7�b���1<��J�0;��ΰFD[�/_x*z�f����]�WU`R^��{�cy�o��� ̗�j6�HZ[���({Ⱥ��ʗŝ���*��K�3��Y��h*�Wr��<bU��c�y|,�M���ԑ��V�}}=egb��3Ӟ|$eOS���@�8��w+���9T'�5}��"c�s�x��gM�x�bq�����<Я�q��LSl*�0�Fշ'6�]Gk��n$٘mNw猓�)2}A��[�n����.�v'�r�+桠@ӱ�ϓ��1=�o��'���6Ky��������\٢�:���>	5�2��{�k�ro���q���V8=on2ß��,y�����1U�r�zw�K�QL������ER7��Ǆ����F�]�|�R�c{*��٨'[[�D�"��K�r�y�yunS��6�M
���_m�3�n31U��z	Vs3�v2�;���{5�	�QX����s�3�1�y�o���j��}�������=5�������Η�p���ώ�"�>�8���_n>RfIAN��J�-�TF(Ǯ/#qD�rǳ��T{��^��r /{�,wgp3�Nb�T}��'Xr��}��f-�Ԍ9�9���e�8�n]��c�utFJY9��kDی�c�Nr�}���ʷW>r�P �q�#�7���$���gE�R56��f�_yvy���{<�(F��C6�˜fc�����/:��u�ؿ}�}�59�×w�h]�^����s��=�Q;jL�?I��}�5]�����Iݪ>8��j�֌s�ѾF���p��C_�H]�zq��;��=�L�&N�}y]��<�-no�����UU�nj'z%򠵹ؑ5J�k��Z����KsW>��Mެ;j-0�+��2�+5r�У��3�Уd�kS�,U�wZ��od�M�	X��2���5ִ�q�=c�����{��t��/��e'�F�ʇ(�n�GZ�ws�}6lu�9�B�{�њ�s�:��D��g��of��w7��;sVvg�&q�I�nm/�D?�#���Fզ�ĭyٖνh�l=@�������u#&��=��F�f&0��4����Wd�'�`
���<fro
����!����Ъ�j&9ۘ�<�n�̫[oH�mz��犱��u�Gqmr��\��ǻq�����~�;z�ڎ�^@���W�P��:\�]`Fz���X!xf����D�gZ٭Ju �G�D�[���쭳z�&c�������KeE-��ܧ#��s�ܜ7pT�n&xJ����3O�����Nͼ��cۨp�w`rwi�ǵ��7�/8����;�5Z�u�9�U�Ӌf:[=.��C��[�W���������d&6^,�Y=P�ncQ(,�t:�:ou�k�kV��r��ߦ\[�\v�)�b�Ԟ��Q����5�	�p�^�_S޽�Q�9�P�q!v���u.�<��ʗ5]����V�e�[��:��(y+��<r��ڢ ��7����)�\-NÄ*R��֞\=O�����ذ׽Ro��;hq�m%�ώ�Nq͜�;��FUw땾�}�>�j�J�^>}Ξ#��G\����X�Gs&�7�����N&�s��)r�=��ٯ�������t���7�u�R��O��<���:�5n$��J&�57�kqT$Ҹ|;��!���Ȭ���Z��&�3Wܹ�g����ƛG
]�n�����z�E(7��;Vm��R��A�Ӏ!���`ga�˪A�VM���U�{�յk�:�v#t,�rӮ��G��KVj�
��Rp���/�Q"8(w̝�k���}���u�T~�Y�'~�Ï�Wv�S���Л��~��1Y�	��[:��n8����V��١�K�ٞ��W�0�Da�[q6%k���-s��=��Z��p��+�5齏z����}n�J�bOB�<��3���4��sS!d���s�Ժ�ak���B����U9���ֈx�j�U��&0f2, 3�P�K��:�>�
c9���>�؄n�o�ą��o%��q铋��x��ŀ�؜�m��N�8qŨ��fiv՜���3��W_���Ϟ��;�1���/����}m��*+0է�9�ˇ�ꇲg���o����\Z����R��x�K��խ���'��p��*1�(�k��ݫj�{��"����|qs��_!z�*����8��JSX������*�9���W4����̔B��z{�9x�3��EXP���袹�{f�� ĵFo]+�ه8����E��6j���-�ƶ/U��=t�tvz�L���/2��sM[Q`v�Ol<�J�n��R�9}��M5a �-5Ѹc��ή��o���1l��Y�dN^O|{/`G�| ����Ȼ����_{�Qʾ�++Syy��~s}ܶ����|}F��s�5�J�n	�	�A�n��������i��v��^�nS�è��z�����p���Jz��pgz&�*�);�U��+��˸�;Ʀ�k=<�¹e�$�K�]��hY���w�p��	F�WsSq���iqn�iΨZ�%s8�+u����|;��br���X!.�=nM�ǟ]M��]��m���Ȟ�����Ok�]]����mpW�2]Қ��2�CSf5(An���d�u�i�Zb��I�ٗ��[
u������.�݅eLR3i��Lj��q�IS�����s`�nd7w�\��9�K�`��|R�LM�,��v;eP��M�N@qt��y�[�i�E�s�f1c��+��P��=�G׽��bީ�r̷�b�\4�^Y�|&��FFo"���.V{�R��g-bN�Mb�-�Eǋ	Kǵbh�������Сg��++w]I;��ܾ�O1��p
�AI���;�{����p�����%Δs�����}Y���T>O- �L��=�����ͽ�mn�-�Y齽ܪ����d�x�8�<���9ܭ\ln���ր�h�t;==�(�����,�}�6�
���vw���`r��KycѼ+�Ѩ�h"����>���*��c�6syǱa�oAGf�]�9:�$ed��ܩ�F3ч�J��4��9�����Q5c��ǛE���uk#�va7�_h�Al����ګap���y��� �����%k�k���-`S��9fү�p�#��f�,�y ��t͸Α�nzW�Q�iУ��4#6��>�ĕwf3b*�⾤�QV�T����w!\�̕��yt@W���XY%���Tͩ}�t]��HP�{���*�@ww��z4�R����Θw�C��dٽ�F�3L�'�rښOv�+�V!�O={������o�to=Ф���*���l�6E�S�'p]�=��L�S�l��#<�b�o�-���8���"��k���hi��k�; ��i��H�ʌs��e��r�� 1Ԥ��Q�At*-o����{ޏ:��������8e��l�Κu��"y�����F�#����jXW��&�>׼ה��/mT]B�X�ܾ���l\�(���\��v��o��c����YCǣ�<���a�z� Ǘ4���V�U��vg�^�.W�oֆ��;�PN*���z+���Y���
M�=x��4�/���`�2�3D͠����]O@��Ń�ҁ����o���򝛒�r[ɚqA�d��N�1�Yժ�l˖y]�`�"
������S��=��ڻS�N��6��s�Tr�%/�&�1z5fء��U\Swlv��$Y׽ǎ�;]g���wh���،���˵�h�bp����#O���E8ay�����^o<8�3��z9 ����{R�Us7B�b7��u٦��2+-Q[�W��Un�D3|����)�>��'�(K��ٍT��s��n�J�Ym͹��
rg��N������N�L� }�x^<�P�R�a����y��$a�h	��׺ż�JV�:b��t� �f`�Y+�HVi��l��FR[:�T�����ꮸhf�5�F:M�X�Is�W�+�E\�������b��ޠ�f�(�f���+ډH�J�qQU���W�0�ܙ9�����R�I{ų	B�ө�R;�fH��6�yY!��w���ݫ�r���Ki�\�1c�$��[b����0O�I=���2��b�'�v�0o��պ�"�h%�>w�)�t���]@/���HR�.�L����<`�Ֆ>��OB�Kg�t�J30�B@��(��ə33S1U�Wᯎ�Wݥf��n�;m�Q���g���I+T���=��)��S���fd�J�,TnV��!l��;Pޚ=~�y߭zm�W5�k��BQ*�lT�66��t��ݹ�6����%n��775��\ڒ�.�j5��\�[�k���r�7����(�3��ub�DZ1���ܭˎ�[s\�[�M�t�����*��m˻���r�-�nW+r�ʝ�-'8W79�sswv���\���\�ι���]��Q��i�\�\�ɣDl%%n�9vXœ���J����[��c���;A�(���ۨ�Ku- ��n��Q�1j�n�8K��R�/g��v�pn�z�}��o&��V���y#)�pz��Q�S�\+���ُ̤�J�y����]��m��G�"���TgHQ_bc['O v����l��ɒ^g$���*���K�K<qq�,[�}B�ud�^���SջV�2���mL�β�e�v�LECU;�Uk���:��2��Q1����W�_KTY�_�z9�^!�9\^u�;��y�]�/m.��Ly>�v�>���6I�WnD%��b��}e�C�`귅 ��l��j������iJ1�/*�-��el\��+�(����&��}
kz�����EZF�j�D��Y=q��V�����Y���F�N!m��-�ㇻp��S\�pY��U�-�����c�*�K�>�z��]醗�o�m	�"�A��=�R�G	X�ɋT���um�������=�
Vo>�]3[��}	��q�2~wJ`�l	��dЭ���mw�n%�1��e+C˶B>U�7�Mj?WAy�WG[�Z�5ܬ�)C p�gC�}r�Q ����vl!{8'�^ �8�Y�K�g������p�R�k��W����9uZ�Ŷ�����%/je�zk�&e����/���or��N�s�*�}wv]�sY�W�[�	愜^*�*�9\����5c��ʍ�l��}Q�ۉ�~��,>̿��3��֌�[�2�_=j��l��
���J�szm�on2���5���]���j��Ί��:��j�����p��C�d���V�Z���i�13����s�Q/�{�_od�CϹ8|����TOK/r��f�qf�V�r�f8W�x�cV�8��S�Π��I��e:��d��fk��[��Sq!'rW�:�-c������j��Kt����^�OG`�r�4b�t@��s�+T��2U����\v�)�GؗQ��2�W���;A�{��V���zmz����/f�o*{��T?g/�^ڥԺU�1J�K}U9��Wk��m>���{U�Ϣ��y��7�Q���]c^�t R#�ڸ���M[���k���l�G���R�*ĭS�!O��P?~����b�s��=�^Bh��/L�4m�y���P��K������vo:ϛ�e��MFG�P��tXt뵟D-���$<]��]�JP�k��S�z"ǋs����SW������5��4����f�����s��*0�+��Y�ިɅ�U[�+�ƫUS��>�v���+�anrqh榗j�m��+ј���-���c�~��wJK"7^��Zi��u��`��f[�*��&��^�ق�MrjoMn$�Eŵ{un�����=�5��x�Td����U�J�rۉ71�\.u�����')�8k<�{�*����m�#o�9�T���5_a�[M�Z�&"j{E�V�h�'������Jxs�?lu��B�C˘�к��P���
F�<V�ʍX������wn��_0�䶕����K!_��c���[����\�췒�&Lo'���b�x�a���v��ݪ���#�{9d��D�c}!�g�J�M߉�Ό���Zy��.V'�O�U�H{�L�̜n��I]�,�,�-����ݓ�τ�k���DJ��)CGW��&&�s�7L�W6���naۍ�� ϽRK����/mC��������K2����G�&\ѓLOL~#����V�Ų���aB�ָ���<Ys}v\����79�͚��+�������3E��Db�8�֞�c��3<�v��a�Z@�������t=�)���q��-V�oUE��ƭ�k�,p�3�C�d�L-}�b�ʓ������ͪ^AmO ١�*�^c��..��W&'�b����/*75E_-}96�r�6Օ�j鼊s��E^B���Ƞ�QT�ҫ8��qʾҲ�SycO���f�ud�!٢Ayc�+�c�Ī��C�&��V�VyTY|�OO�3��Z�iC��9%� 
���8�S��񇧥�}y6�us8k���YI�j�����g��|���ݸM�|����ajЧ�5n$�J.+��p�!tg����z�w�r�y*_t��k�N1��S�[rH�ً�f��*we����U̕8�j���[��K�
�d��5�7,��_�XT�U�x:ד��5�5�|!�fy�dnm2ǵ�����*nCa#|�����2�g�ս�u�7̥�@|¬�o�XJi�_��[N��1[{����/�U���[��јD2�.��x��7+7_"�[y.�Gn����O�ɴo����ps+*oz�^�\ٗ��uTF��ؾ	7
b�9#(As��!�nJՕ�a�T1��9�}:�+s.y��W1����[J�l��`ӓ�Ì�-�:�B�-�\O��LQ�\�x���߳�e.^f�����'Lm�ԍJ��}c�]�	o�BY�	��Rw3�n:)�۝��W�}`��яV2�;�m���u��T��1�:YO��ef.�L�~��2K��i^����@���p3�v[��
+_7յm����6��#���V�nr����օq����v��Pb:TOs������Q	��hv���<�Z�d~t7޽�8�e�k�|qC�Q�?Rhu*������0ז�����B+T�������7c�WM�*��<Q˴���㽺�3����y�oC�L=︷�����mQ�;�J�͡U��ms�=;.d�nW�7�"�ER�r�Øm�|�S���N�ɸ�3�.���6����S��}�]�C�'�͛W+j��3��67dN�ۯ�{N���ע���\�r��E2(�|�e-Ӽ��%J}qoJ��v|$��qQ뻝����f[��`v��������$&��=��aOv\7���������އې��1V���[�y3\��C�����j�Jyx���ͽ�5˅��.P�������6�B�:-1i�
m��X���1t��\Wu��=��9���[�:�v�B&����.�'S2+�Y�[ql7K[��t�f�P�u&7V8�)T�-\9ؚm���6f��5XcV��|;П��+�5����Lu��v�I���֐�ur3�ѝ__�+*c#�����ʽ	u|L��v�v^fJ���=��p�jj>|��.㩻�s��c���63���A|=n�	�XG}+�d?��c.\�1ܩXN_�\:�yӘ�϶�����)Ìl�ލ�Y��ۖ��;ּ��vq�N ���ĵd����&�>�Qۉ!�`g�C5��U�j5h3���O8������x��U֘)��6_$uz�$�v���4�Eb#�gG��uФF����f�ݗL_e\�C�^�[�L1��/͔&nO+����_�T��l57�e�qi��3k%��l���s6e�mrYY��� o��g�$�_w��)
����5�kf+�Q^aX�["�z���z��ڙqo�x�tV%�AuJ��m.�~�u��U��lk��qt�:�ԛY��g'���e�и��>ſ.��}K%�TE77����|�CN�"����sP���!��is8���D/d��s\Ú�E�2�Gn��J�w3��kz)ssО.���e��טX��V�ĸ�����u*Ml�ޡ��4��M�O��G!���9�q��%��㦫|}+���9Y3�ʾ�ά�w��F�����q�º�S]Lp�	�G�U�0���q�+��Xv/�J&�+���һ���wѷ�:��!�yk�8���4����-6�6��&ֱ�������x���V���g�S��zm������W/��eg�9LY�J�M�}ws��*�Tk�u�p��c�N�ξ���
��q��Y�V�1la�[q6(-c4g�Vߝ�3u�-�(( ���J/	�O:L{�S���-^����i�H>�zw+p˙.��޾j``^@��!]�R�=�&7Ə�/5*f��oI��[M�R(���˘�!֒M
C���B��yǧw\Km�uxC!���j4`�V��n�C�)d�i<������:�r̰�n�+i\lu�ͽ���>E��V6U�j��rf����9�-$G%A�<�k3`+�a�[J�p�૎��/�{���*�2�Ӑ�eN�Â�^�����O,s��&"���Drp�u�f���8�Qs.x��ss��8��G�P��(�Ҽ+
�{&�=�ᵵ��YϪ�S�k�jf��$n�~�]���?y��'I/
]����K�p����ƻk��P�E�)�8�Lk�o��Z�n2:���-�uO�wճ�g��j���Fu}�c���<qk���,���O ������^�}6we�O7u�*n:��-mWأF����b+�=��7�����R��Su[f���9UYV.�q�q}J�=�-�*�J��SycO�>w�d�v��"�B�q���K�����BUAWï�1ZՎ[e�ê���U/E׀�t���^1rEi�Kܘ�W}���d���wQ֕��#Gڠ�݁"��;eL�ŕ��@|3O��`�x�~z2:Ɗ�k������ �Pݨm���ס����n]W\�zC�vݧ=zp�<me�Wu�eE��L'���������y������VV�v����c�C��S��z�޸�\AĲ�>�����I�~ZW��[I���SۃM`ˁ�W3��\�D]�KmM,u4�����0�7��]a*��е��;�r���+�TbK��87�w��LVhZ�J�	��uJ[(�{v3����퍹���bt�va��c�t.�М�n��S��9���Q���\.�|M,�)#L=H�넰F�؛"V�\�,+���.���/c3�{_V}/+�vz��'�{�m>��*�1Pzۂ���1]�b1c���w4o:��8�ݾ�Lp��mC���D�����}�ie�^*������&��m˱�����{G��6�5'�p�l�͈̾�׳`��ȧ"��b�'r�����1�l�Q�!EF&6�nrk���m�D��Ãh9�Y�k[�N��5�)Ew#aQ�Y;�`������R�_l��J��U��Ī6���]����oZ�`�7�(A���ʔ66�Ѝj�U���c��G^ڧu�S'Ah��Qwp�;�$}b��}�ܼ��:&�e��L��:�bWu�T��92���z��r����Q�VҞ~������f�OH�)�Z����ӴbC����߂�B��u/mk���\��Ԇe���c*��V�����͹�%�<��ڪ�.�!{WTU���Q�\"�[kh��M�gg��T4������ ��ؚ��W�gND`��a��س��I����m����F����Ī*��j�6��<��ȶ�1���u�����-T�4�����͸څ��4,شÛ"��V<=͠��غ�q[O��+ؿ��%7���*�+���v��L'M����"���qU�ӤB��S��r�{�	D�-n�t�_r��1�F�(�Ⴏ���s��v�A�L��ٍJ����B~���]����^���)���A�*}(��M�4;N1[���LW0�a��ᱜ��П}K��XU����{��Y���3�6|� �����|��1��^<ѧ�O�Ԉ���(^��5�30���w�N���9��=ՃP��,�  �,�7�W[\wP鶲;��EӴ��
�Q.Ąz�<Xo0�a�|��:��/LQeggH�m�u���i�:��7�ʍ�a���a{�Q�4l��'�Xy2�5���w��5PU��l��NQ"6����ˈ�fwu�ރi�e��f�g}ڸ)\������"�2u�/�Xgc<�2�A�Yz������Ib�IB�{ /���IZ���"��ȓgQvpRdI��V���]����{�+T��Z�� �iM�0-��ݥ�#T�Z��p��m ���z���E�n�W}���dݫ�s[�7�V�e�o�	����73W�J�'j��r���aiI�MZ�/t&�9��Ve�b�lgr��*�����ȡ}oU�eG��L&�ؓ�G��XS��06��K�-�B>�f�G��$9!h�`s-xZ��O�Z �O�]��xӵ}i:�]&E��u�s���[�/���a f)[�W��X�U�.��}�72�4B�s}C>���� ˋ��m43-�wV��S�wi�Νe��3b�F�W�#ų�{������hP(Іqo������n2�n�����,��fhו����7F2g��`�!.{�C��c,�]�ǁiŕ�%�8:��V�=7�t��(��� cj�ʤ�Y	�p��{dt�#�gbf�����0J�V�����%©�.AT{�����7��p���T�^���nRG��Lm���AG*�8vWs{7�	꼮�w�ϡF��Sr���v��+H���S/d4��ó`���Oy����0c�gV���ǻ��x�٦�s�![O,��~��7��չl\�[�o�X���(�2nI��5m����6�DY��Lhyk��Wv㴵�}F�J�B�fl]S2h�S�`�]����c;�L�����2|vv�np�̫����;����؈��ש��9�	�i�6�Kl����&i5۽A�.6��q'�9+�r=���rE�����x�w�p�k�VK`�&Ҕu�Qp�A5K��!gZ�Q�U�J˰,l/p:A@V���T�m�G9��ݖ֯�9��/e���[0��LGb��̽�b���(�Q셋n^�x�� �����Ǚ��N��آ\/2ᷡɤ�.%+'v�'L�(�sz%��/�A����i��O�2,�^	�ᆖ.�m�ӂY�w�x-��_fz��ZU�dӍJa�ǫ���+����gJ�蘷Ӕ���5���8�Ø<�`�]r�T0�״E��t���*L�.��ܫl*�n�}�م
�u��ލ��q��o��r��ʾ�kNn���e��Frq�n�d�@������z9͒��i�]W���P�vԵ���Hp L?K�ni5�����B�Aup���5F�k��jwss\-9�;�wvwt�ۜ��C�nt���RcC��$�nZd�;34���"��d���.���s;�bww;��:�,���tŋ�ww.��H���I�s�]��n����ȑnN�g;K��r.�98�\��u���]���wU��$;����v��ΐ�ݫ�ē$�ݧ9��&!1��wf4��]����]n��L� �݉��h��7u��s��)�h��sv(�u�C��[�;��л�{���s׾�붝�!�ʣZ:�ؔ���x��P���m�H=`[�1��1|b�r/ǎQ���3��{W\�I�^]�Ga_��M��l<�ϼ4���V�a��4���U�%ӳ�ΐ3�+]��eL���a��t�=Ε���UC��t�>�5��7v�����Hh���*�w��M�<�U//f�(/�!�-p�A8�߲���k��,Ev��5{ ��d�#6#H�ߊ��|�b�gҩ�t��&6���������3��]�B^�ݩ*��p�������ū��j�-���tuͫͻi>��7�k9�n�5��	����3�hʯeŴ��[7��1��o,��\Mj�j�j+c���z��=���/���6~���8�])޿���Q(�{�p�O=^����Օ���=�:�x�k�\��w�n�c/\�4��W&���R���TY\�,�)��|�nE70�����fȮ���m�}�za���\T�ol�:Y�p�+�ƫZ���Ϲ�ɹ�e��@PkϏ����͎5?Y�2[��n�5V_�g;Yl;�S{���d�����U���os��W8ʉy�R��Q?x��8y<j,�x��\mwO��:��۔�:I���a�[��+u�$E�F�8z�s[�q�Q�\��Z��_�ы�?��w���JQO�����A�]��LK���+``����YIf�Y�#ymo��>9Pjܚ���Mrjn>��#�!B��W2�5�_χr���K�J��U���1ɋ��Z�W�[p⺚�=^�`w8�ޘ���k��hY�u��qZ�>��	oA+��M�p!-��n����yqvd7��譥lu��B�v'�r�rZ�m��Zf��z��ކ�>�2z��1ۓX��s�>]2�4�y
�)[mgd�-��ƙ���^�uFl-�U�ʟ����y־�9U�'�"h�Jd��1�I����uu]�ǔ��Fhf�Ev�ᔹX��π��N{Z3s�3Xޗ���7jN�y7~�k߰yZ�����+����e߫H�Ck���^�;՝8��s=_=�1	��p2�W���Щ�0�^/9eI��scovLv��ީ��n�i���^�3/L��e�8*G�FQ�+%��ƃ�n��F��ĦywdBC1�mz73ژ�������=�;X3�w����t�*t�diG�7MA����n� f���_k��R�)2�ܢ��N��O7�g��𒔢�.s�����,Iы�TΩ<}O���^�X����{�K�o��jy�����nv�<p���.��Lyo�ul������n�Q7}6�u����%�z9��/nf.��u�un9V���뭦�^8��1�PL^0� ��귩�.���C�Q���'i�w6��j��bq%z��ʡ���v�v��Mv_ڰ.�bU|�Bӆ��?o�.�?-��F�)'*�?W������Kr7^�����4��L-����:�uW�*&�p�崍�*Z}7�����Ҹ|;v��OН7|q�xa(����
����)���tR"��w�v.��T��[o�yy?;�.�]���%�Q�y��9t��T�pW?E}�	��؅:ݳ�;�Vh��O@}�nH볰Қ���f~w.b��j�sۉ�bV�XO2�
���+{�w���!J�4�-�=�5�O�gs�z���Ɵ%�N�_Y�=�o7=�bJz� ~;����xѠ��X�󐍧[��b����t��q[O��O�}�����@M��'�mv���fe��Ѫ_Z�G�����W��oujv1w-<g)��aka_���1_��p]����"��,zh�����dOUl�',����dV)8�ʯ�8}ed:�j6z�*_m���"�&�����׆+i>�����{�#�,�BN�58��n%�����L�^re��~��ܔ�+�~kA�Pcj��!E�֍���t���m�\�^]n@���V3b`W;��u��ד����P~�Q=�_ژ�0.�f��zg�{�������{�l�첶�.:qM>���y��i�hc\�q�1���p�!�_K��W.ʈ{�j9aݸ/0uī����!{iuN.�iB�u�Ln7�{o��>�|����v����Wְ���1��!���z���yoTk�)qSW�*�-���&�b�l�w����[�z�&l�i�`偡�n�m��P�j�i7VW=T�4�����oj�.@�jE����<��ڷ����a5b��_U_m">��-fc5رr��e<�E��T��Ü�����_G}����m���D7���b�b�x+E,�q�C2�"#f���f�N�q�3�;hXG�[A�$���&N��T��*�Dy�EG�{����,��٨-��sSq���鯏.�P�-8��cfʬ��L��s�	؄��j�ܔ�b��q��+uT)}�K����yϕ�u ��&�3M�*��U�9m�&��]�]��Έ*�.][�����qK�*��Z�3��jE;8�|��c�`+��8}=Ǟ�^d�`ŕ�ŉ9�\��P�i_��f�/#����\Ɖ]���[C���	�m^Z�(|1�-�wfhw1!Os�ak��������tjO&C�[�]���s�7�3��2�TZ�?c�:�#�,�'\8�8��DѾ�o*\��uc���q|�P��(�+���aw��w���7�Nȭ�g��>����H���w�qh\w���Eb�]�P���Ʋ��Ә�I��<Q�O瓛�.g��Jvo9�ܧ#��ą�!�*�����z��������c>V�$Ař{��٢���9�&2��V��t����):�f%�U��7�7�K'����]��BeOf��X=
�+�bt-�`}m���r�܅�K�L�yI�^ao%B��`���HO]uqvq����릗�����\(�u����%d��ڜ��5�ߗ�{S�y"�s�Vs��~�:l3��rR���tZ�/+���<�w���=�5γ��"tk���Vº��P\)��ͺV1�z�vg5m�۟7���-]��T����k��N5Ī.�75u���+�j�ZS�|�zXW;|�>��ue�f�Y�N��ḕ_�3U�C;�>�N7�����b6;Y|⹣IV<��w�.6iN��gvU0�Cj�t����	+5���7M{�ӝu��G�!����޸m*�z7z��O��*e�ц��1�n$ݱwG)�������b��)�]w���U|�_\7��8�O,�*{~f�_b���l)�z�1��M��� ≯	������Z�TCyO��j�ݷ�"���������t90�=ーV�ɨ�Ov¾a����'z.�W���ۋ^��$��3��IQ�:��ˮ9]�R���&�`��ݽOyv�T����J�5v���9s(	Ĝa.WS"�f�ۋ�Y/�0��R|:�UYeѹ&[=��g��XKt=r9�}�G]�w�T� ����U�ӥ�Z�i�:4kZ�����
����D�>��eh����F��"�ŎkVOݴPī.
��'v�6��l�n�UO���'��KVʛ�}�˼��Q��,�H�rk+T�0�$Mv�4�	�VTs���N�78�5�Gq�~��g1�e%�_�tF��=��qq��(���0��7z�FGK�l�������r�cQ�<zC�[O�an+I�^NTb�u��J��n���2k���HU�@���fGE�qS�[9���j�OF(Ť���Q1Jڛ�&���L^ѵ�2T:�g�[���W�T�:�U�_R�8��,
�jo3[뛪3"3���j��_t�1=6������;{�C�\G�~����Dz{�a��]�L�ySj ����&�R�����hN��-��C�H$��h��8Ş>�mg�M\j�ZWe���n{Ji��ajЧ����_��++�����ֈ1�Ʒ�I<޻R��)�[��Z%v]j�>;1�U�Ѷ�oFڲ�^�5��G�N�'a�'���R�oN֢Vd�R�8;��$t]�q	��z���<ASOm�^s4��Y���=�z��,7�V>ʺ�R�hwK5��a{��̐Wk/+�W\�-J��m�;��%*��ܥ��~�8�ҷ̮�y�広�l����
����d��-?��s���.wb��U��p��W�8��v\��"�$��n(l�8���}�����I_\ٗ9��T�[z�!�֞ꄲ�!z�FH�ˡX˺�Q����'�:g4�_y#W�M�-;���CN����
q�)[6�
��n�UӘ�b�����؀��T��٣Jޡ�@v8s�*�Bf98n�+!�5�ɞR��q��e:�j	՝�x�Z�]�zǧr|���g<��q�BN�59���W��P�t�+Oy�b�;�1�np;�̾���Qx���3�l�s�(ߓ?7*s�]ᬩ[y��uc�m�T�eŴ����+��O�L�ʓ��^/Te�|k�<
\�OF9^ ^z�D�~�ڜ�f��V��h�G�WQ��(���GSn�ј�LO��ۈ0*y%��A���Ps}!"�.+޳
��/:k{�1T�g�V�y�;JҲ�N��Yͣ2�v�F�-�@��,L���S(�g��'�Kg4uJ���B!�����PV.NY��I8��ϫ����^��I�_w�����'o~��f��E����+�*{5z���+~�.��s*p���w�Q��}����&�ڝ!n:w�X�1p^��6�Wh����r���_in�!4�e�]7��ּbS�ݬ���J��n�G+&aħ�.ues��Xj �yne6����Ĭ�Ftt����yڅ��)��0�f�7R���tS�Q�w\b���
���r���Y��k���;�p%�T="��K[�]Y�lQ�Q��Fg+�6��n��Yؽq7��QY��{���ݨT�/M�&�"~�V�8��96V8��_9���4sqk�؉�V�O0�Fզ����;�{�㊺��\Ѭ2�\Y��#^��U�W��l���E�\��\&�z�������
���3�&�ݿ���
c�Ұ�>��@u���m�Lݓ�,�x�<�t>Ҁw�e�V4���K��N}z�P�nhT�C;�wy�!!���]z�h˧K:�U�3���(n��H�.�Z�+8�`
1��v3^���Cϵ_b�_hc����m��ͽ�1�{H+�L)����o���6v�i9
f�?^o����t����#�$h��Gva�^��4𢽴|�W˗�~~Q��{�'z�a���Ng�U��As��%�f��3����<��+�i�.�}7}�饆ߌ�ɛ��]U���5�S6�5Q�]C��Aq><�Z��V7z�v���
͛�'*�v���θ��z��ݫ��I�ݸ6��+��s����#��OS�����oW�r{�{6��{<�dz��W���b�jOn��W��9��U�'P����4���Q5���O7��k�pӚ��b�ʞD��v�<��Z+o��T{b���u�ɟ����\s��N}�u�{}��΢�t�|zP�p;��S�B){����D��P�7�s�Q`LWz��FL�d�ǝ�5�״��Y�b1�������d��G{���=%����@�O}G���Eϓ���!q�kYc���ٛ�	�y�>�P���$s�t�㑾����_��!N�eƒ+��@>�mꗟ�ʪ[�6���B�&����K�U^�M�`�HH��-��j1w���;F��ݜ(	5�Oj�la��D�{	p�%�3�0h����6ƶ����EJ��8�P6�ɘ�K���4nK[;:�n�6�+#�u�NjwS�S���}��^
;�l�p]W˗�Vv
��|��<\�z�L��^`l�l7�G:Z�=ճhC2�����0��Y��Xtj�W=="���Hab�hX�m���_5N���q�v,v͝��"�)���gX F���*�`�B�껝� �����5����]��8���w���������[��y���-�����bT���v��s}�GgV�K���-�$�j�X�VP�/�޺�P�n"pk���4IZ;5�T9�'��
��gnY�)i���Q���[�.�y���5���G^-�lgm�F���t�p�+d5\�(kt�Վ|���5\e�c��� u��vbά�Y��WON>��JZ���[;��U�z����'C9VL]�V@�3J+d��+3`�2���ǽhL��q�.#�9S�oY��9�5��D�����d�^�v��:pP��vK�&2;L�u��:ݨ�	2d���n��7���`�`�G���������o��y�g�pD'��SN�7��>�Ѭ{y㫱Cg��ǔ�#yP)���ڻ�;m�>f1:4X�K������uy'b�"�bn��tI�L�\wv[�u2�'�T�<�Y�WU�m����N�[��%���#h�yW�&�'o]]N,���{��g����mS�OIp�{�{�ƪ�p>��TI�%�(���h4:�F���$�w6.���oq�YSY>���0�6��'34s�&e�W��{�vm%�Lcv�����G�.��ޞj�Y� f��+H�{�]�J�;��[�E�.2w��	�Z��*�_�Ɯ@Ԣ%p;G�^�O5\�`��*m�o�X�(��Y]a���&B�0��쁻�����N`y%����!�!�X�\4��0ʻ!܉Ι�pW#���4#c(���W���Ն��q�P]�Y�$Ү�$!�ٿ)*K��(]���B2���;���d!����g�T1a`F���(�ݖ��!a�B���CG���^E�ڼ���WJ]������)��&�}��9�2���b
�#q��\�%k�����B�ߦ=�n�b�c�7���'J�:L�puԠ�2Ý꛶�����$��8ۺ�_UJ�6��'0�A[�����2(���MƯEa�rv�=�x`5��*li�3�KW��(Ҷ�DԐ�I��e��u�JgQ�6�<�3��h���w*=��Ԡ\a`E�^���a�yڽ�E��o䘒���F�Wg�VwT���t�qz4�_ݸ����K��{)j	�����n�떔�Bb�:�lK�^u(yH��}0��Q>������1PH���=�\�`�$:�İp�,eTܨ��㟿޽������h�;v�.\I�)���۷-��q�\��nr� r�P��@��DwUĘ�)+���]�J�R.n�n!I4k��llQQL�w[�1L�ܗ: �u�P��"���,Q��s��$(�k�9����:�		2�(1%��L7wq�s!�1�#.�d9�HhSL
6��tJk����fI�C �2�W.�;H�K&�;���2� �.nd�r顙�B�D���)\��̻�FDR$��	n뱌���0����@�\�@;��]�rB$�]� � a�)��SR��1�� �$�$ H<�{Ff��yW}$�+V��m�d~vwng�P�@l0�oF�9Qb�$�څ9�ų:�e��ߨ�.��@X��i����Ҿ��lǸt�s�a����ȟNߤ� 6VLO�B�)�s���l�gZ4�~��+|})����U}\���C=�\���q#�^��+���k��7qį �;�)Pa�}��ݟUa11K���%���%�T.�M^2(����r[�=�Pʺ�XV����=�7�|���A {M.�>��i~=�aᯗ��7�L��<0����D��g}��s|�� :׶��y~��P�\&h1��C���['C��=��z��q]���R����k��P���l����3�3���P��.�ς��W^����N���F%8Sؤ󻶮�8o��߬B����J����ƿE>��s9Sf��?He���?�{>���;���~�/X�����4=�{���Zn5�vX^��V����zT߹Պ�eb1qށ=��H�K�ͻ��v�5����e���,_ٳZn#} o�:����/��q�̬���C�>�f�f����7O�9�� ��43�~��e��}UFV�<��d{$xf�=i��M����K��Y���M��X��yghn�.��ŵ��t�E���ģ��M�"�Z24MǷۛs�z-a[�r�-�\ӕ�{}�.�z�v���BN�(Rh�.(}Ð�{��5R*\�������-�FmZ+U�f�
�}n� '8��mɜ�
��j��c��SN���st�	�?����#.Z���!y�4�N*z�Q���L���&o�c}��	su�㚦��z\����>�>�]�Q�4�����(��]L9��]U`M���d�s:d��5�=�z۞?�{�>~����d����q�΃<�}DS7�@>ʬ}R�<c!x�nн��G�3��=Ӟ>�/����_OM4tkC��}��<�=ಥ�Y�;"V[?��{��!��&)�)w���y"䵐+�r�u�L*�V��{������F�����G���
�,[��P���dU�B�3!�ofTvUH�R�K��l�K���X�~���9\N߰Wj�x��n��s�P�u�ё�����72}9FFT��a���	��K��Ԯ�Ƽ�\x�=E��\��a�A���~� ;��ȧ�N�������J�쬢'�s�w �oW;C��
U�:<�n���&;�Lw����W���K��>�P}칒*��۟e�,ܢ=����u&��G�k�B͖������=�_*�����C�r%��������W��9S�{�U�m� �,}{jP?�JC�:F$�����d�}5��gaB ��U��j��p<4M�a~쬭^�;����N&��FT�a����`gS�6�Q��I�iUMO��ą5���٨s��ZS�:3��B�vT�I�*�������,t�gA��<��,V���?P*o�fY��� Bu��V�]7��`�>tw�e��OT.����6������F� OW���UE��;/����8+7�ŹGѝ��ZQ'�\z���;P��a�ͪӡ���S OЩ�e?/f�\�)m���:��T��G���G=�ۡy	�Pߝ�+ftf��vX��ۅq��si`o�j��u��\�b��E��^�u�~u�=^�F�^x�*�ݢ�Z{R;�D�kAS,]���{H:[�g�~�X��'ڮaqO�����������=���Ǒ�}|�F�%�[�Q�۩��V��mw�U�0=��,^L�7�L�^Dt�n�{�C�#����u��s��?
�8���u���s���Ug!���,�;34�DE�L��2��:���O��{g�{#ޯxNb���釣k#;���ht}��������t	��Ex�Q�����I=���p��u��5r���EG�{]���_�)�,��[���r�����\��ճ���~�%F��~d�Z��d��(���rQ>⸅v{���Q� �=ػ�t�R<X� Mʚmlp�۫l�WxaH� ��Ht�s��3VK��\Ie*;'[J�l޶���$%�mj�|�X��[���BM<-�*���˥�1�>��P�<j���o���	�PÝo��oB*��V�G"�R�����Q�w"�ު���dΘ)��_K�#�����Qt8o��.0z��^�O#}��u����3�J9�.�=�ECʧD��>gL�
ȟ����c�e�)>d��s�F+N�>Qޮ�U�����T�� ��e�W��k�@��c�Y�~��n=L�D�.dF�����݂Ÿ[W%���C�l�J���{��T�F���¦���}{��u��ǹe�rW���3��t=>�����J��Q���D�ѷ�%6���7�<�>_�����܁���j��^��X���sj�m{����mC��~��Z��y��mR��L�G�e�F���g*l��蒎\z����b�Ӂ��v�GG�W�t����� �JgЎ�1�Wۚ����ۉ~ʜ;������c; ]��*�����G��yΊӼF)︰5s��^�Ln��9�*6��s�-{Mw֖Fո�	�Vlϻ@�J(x"�e��d֞�:���@�q�#�q�l_Zn�ƽs�{�{-�q�1��{�%�A�����=���9�d*p ���ter��]�ݩt%��'�]�c�����.�1vj��C�ovw	����嬢���Y[���9����������;b���W��ұГHN)w[�u��'B�Ai�7%�"�Qt	~+����>�;����a�R��γy3��Io}���>�����LY����ׇ�X=���ﻲ��^تD�a�蚋k�p���)���ax�<�w�6�UJ����I��ή>�B�٧���)z��B�իc�{>��
w�t�}9�~�n�Y�r-�k$)g��*��pǐ�Sۉ��i�G��q�������U�*�\ =�@7�UH�{���Q��}���S7$����Ѭ�aU�hm��0��*L�o�i��[�y��,g�1-���)8^��<�8�:�}Q�)��FTD�x��^6�6|E�pv���cO��s��<]G�e�
�̘p�^|o�/K���}�	�|`��긘����9�wpK�����u[8^ׁX2:d��%�z��g!'5�=ِE{)���QM>��r�LS��;_�v	���xO�O�|�=<6c�uwOK��X|}�`6=8 j<�	��&�R<_\�vDnQ�ղt=>�q���~��3��%Ä|Q�u	�~th�~�<�K���r���μK�3��M]xn��z�3����_��͢��U�Ny5τ�tx��A;��ɴv���J��)R�Aev�Q=�� ��{W_�
�&C�U�ͪ;�U����̥nrꖝMv�c|j��k�<`�r��:s2t����M�C�J���<��ϥ-qa�;-������A�>�:RJw@������.�a�_B��w���/_��������9�2��{�����0����?��f��'���5��������;,�����א3�u��gl?m�
�h��Q�~���=�*���������o���NkM�7�,�V��>�W��q]�����O����=�֋~�M�H�8�"��ڇy��:��H���@]j�1���܎n�l׹�w��ן���CGDyh�.1�K=��ѥNQc1UC�s�c�9���/��u������pG�x��jC=��F�^n�w��Af�"��X+*�	���j��d��v�N��j��Lz6g������8����{��d��ëW�}�l��7�E2��{b\k<7h������7�m!��~���}���?��s���-�����n���uK1ǔ[�*gq	��,9�}�lz���슩_L��Ex�[L*�������1q��{#}@o�eEUy'�Z3&w�3�I,�s:}g�m!Q��!�����H���K��l�J븱:�$LDm@�9^y�^d�ʾ��1�`�	�҂��9lכ�;a��Y>h%�g�v� XbH�FK����g)���`�:�m�.NHS@|9<�˕�%�nd�OFp�)�G��]:Y*
%����.qH�ڵO7*��}�rW\}��MO���T����꼕{�9��9A^�w���]z|j�2<����>��22���A-�0�j<�t<��#׻6U����=���z��3����z w�{r�SʧDy��alį��"~�=�N�}�,'�}���~:wO�'p��Ba�ж��2�}'"^�޺�O�������5�p�*~�>��W�
u�,�2=�j�G� ��ٸw�j�vLdC~�zm�<�H���.����*��ѹ���.K�_���nmf�d��k\�3Q�Ǫ!M�F�����	�9����2�Ui����ҧ�M���c�O��}eI�;�]q����0�6���;���� gW�����d���(9%�;��e�׾L���Ƴ��$�����[\���Ɠ�a߭?�u��E!��o&v*��B��7���[�ds��ǻv�?a��3�Tz���s��^V�+�'��&�r���>���j<= >�}�F�ϕ�V�<}^~��.Z�܏>�G"����+��c:m�
��;���s�!Q��ZJs�T������?d����+�=�޷Q�[e�1��l�|�����_��璞�|�>�r�w�]`{�7x��\�e֙C)�Z��3\=m�v�t�,ҍ(=t�
��3�9��2�)]��K�=��u{����h4��@�~/��w%���zi�z�$\Y;�ۏ�&�qձ/91������#��y�L�t.5�m`�/]egu�[��;�����MϼX����'Ƚ$4������u�{b.}�Q�^,���ќ z��8˿m猘^��h��m�3<EO"}~���L���O/ף7�>��-��~�=��e��S~b����p;���^�qe��&� O��V�x��چ�_�����К�Z�񥬙�^�G{K~�������wҫ,���BsQ�@{ӑFFW�����MO�#�h�~�cw�xz)F���ԑ_?IE3����Q~�r��W�z��f'�쩑�/�M5�D̡{98w�ﴻ��:;����l���}��㞙�%{�x�2�Ç2�Q�kȯH�=WS�3�g�����Ǹ[��XL�ϼtdJӹ�,ew����S�g'ޙ,�����W`�����Ye�۞�Pq��Jˏvma1?SU�n#\�wAb�!u\�.!zi��#ޚ�O�^�W{W��z��{@�@˸�y3p.O��5P�v�L;�WI������EB�,Y�gH��3���u�ޅW��y�>�>��>��r����ԣW��j�{NnmC�����S}��χ�-j+��c�j5�Y�s�d��s�"�4ؕ�i��)p�w)�,\ҳ9F�.��쌎����~,��g�T�2�el���*�Ya�\;�uB�K ���Nkkb���w�5a�nD��&�G\�'�p,���B㸷����P޵�3|����}��֋�����ρ�Q�U1�gX���%��TB�q;,e�C��KlO�*}#�}gv:})jw��\�Ň�7ŀ��{�����ݸ���nt�>=:/�%���k�*�����d����e��;�F�o�,N�J�_�N�ܧcݕ_g��[�;}P��{|�^�;>��w�>fp�td��޹]�H��v� U���k}�����S�W�8�}4^fI}=��=��c�-�>��VUG��b�b�&u����O��7����T�n;��ѹ&�1����筜����z�c7�n�!�
sr�s�5�z��L�d�����UO�M9���yR[p;��>��oN}�_g���q
�_�B���g�@S�����67P<_���&$�Y��;�1��i��9ȎyP�>���r7���O���)�,��Ce:���'])�����T�?D�`���L�l�������~�����>�}�w<v��8ݹ������=�O=i��3�bX]�R2�g�+D+�4�%���Ϋ�PϽ�\��7�T}J�
������5yԧ�kW���X���7k������tJ]Pc;��i�:^N�m��}Z�t��+/}�[}ZB˭$^�@��>m��wz˛x����(��-���s�5%�:Ox��&١w�!�z������-��W�	�d���6p���9iE�LG���Z1-������	����9�-��KG��']We+��,+���;��;1�����#Z��w>����77�B�NE`��Ӵv4��0�������Ù��>�C��{ݵl�z���sX W�m�O/�@\J��>5V܍�!ߧd�䲽+R�o�v'�}钨�8��u�s���?X�S:<���O�����H��׆��8�%�	�%����;��;���^[(i��>�Ww��T}1k�Q�q�Uh��l��2���7����G��U)Uˋ�Uz���gt����Zn#\�����~���:���s�w��ޞF�C�Kï&���}�K���ү@,�O��io��y�Zo\��������/m��I��V{?Fw?}�Օ���ZkE�zk��g�;++j竬޹]�uH�ؾޏI�x^d�{<B�����=^�޾�:C�ǹ�7	g:'Ԇ�9�2��<'}5�ݘ��J�/p�JzB�=0>���ۈ^w�9��}���{��ʂ*��Û�V����Ňc0_�t=�tA��7�����b�z�ᖲ�w[_Y�(`����9_��3#}���=��[ͷ_�QY�53�>�ݣU���8�0�U����R�D�eg]㹅I�j�N�'�=w6MV�:�ݭ�.��q��op]�]�IJ�ی�[��[��q�^�fn�_I�K-gS]ciu�7�av��p����;Z�kj�2;�H�i�Pm=�n-�n,t;��v��fL�kn�|��uH>e:��H�xz�7y��1�,)8�g-]憵�G���ȟm�\"���WՌ�����%G��(�.C:�m�ss��}fH�,����,�XB�`z��G�O!��ڠ���0)�p���������^*f�ͭ 3x�	�UǙp����]g�9����<�	k�_8Ֆ�_>c*�������l�Ӣ�/-��e�'�G�z�$��$��9�ᥝ�|QW6���U��7��S��_G\2ӱ%�\��1��W��
֤��yȫ�՘B�{wT�&^�W���/���D�q��x)�v�Vջ�n�j��v���t<�q4ru$#�����;B�uc?_�o69��:��hGEYw4\�3@����	:_�4k�v>�sW"D�{X2[3��U������u����6�mm*5�x,�-��Ś��^Lڊ�$�{�ds���97Mh�*�6�y�4���2�L�z{�¸�s]�f47�*C�;�#OO9���bG]�|Iyt��x�GlW/�6�@�⩰sB�tܞ)Y�+G�^�p�s�mC��w]��t���ޙ��,�&uV�7�͔ (�����գ����:u!��x�7�:5�3k�Fs��.7��XKW�寫!lZ��;c��ҰQW�.�F.�C�L^�d��d�Ai��=z�	���,a�F�u�] �Cy��l%���j�zҕ���`��V{����y�1e��pPv�awZ��Lo%�K��84E����S�b�w�5<B����Y׀�<��iO��`�A�|�����a���n����޾ۈ�S��z��Q	���T����[K3��R*U��O*=������rK��
�A�׋�eg�
I�a�ˋ��󤆕�AYx�3o�^	:�Z��Yz���2��ݽڍ��/8wj�n�S�u&�y����r�5�����Г���4�Ց���X	p����{�H�:�dY���y��{/S.��)����[y���f��c1RG���W���	`>%q�`����u��$7OA�I%A�5�g- t�3��+0�&�,�d�x悵K�PR"EҟwoN7�o��k#Z*��j�rg�2�e��IV�"��8/��&����� U;w�wRi�*�@�����P&�t�Â�n�1����r��ӹ�.u�GH�A�`��:�Tm�@Ҿ���y�f��\�uL�6<�+�H�_h�}����m�ƕ�W����zr"&G9I�bĄ�w]
$�4D����A9t��(×&�#,CDL�-���r��;��%0�EI�q�$�.W	�wwd�7Jd#2,�ܔBIR"$�22�wn�J"���%��J$��"�;�\�Q(Sw]]�3��,c��r܄Fi���ɡGuvL$c�� @���P�d͉���r2���2��\Ffc.���fl��� ȋ&�$a�w;�!�QːbN�1G9"L��34��%(�ٔ\��6nv$�(��ҋ����	��p��9vD$\��2DВD˻���a�ƛ20�Jsp#B\���De�P�R��d�f�;)%�Pwn# =�y�߯~�o����t��&	�.���^�O09��5���5���#Q������Y��3��T�v�ͅ����ǅk䌩���_��zb�e'9��u�=��R;���x�<WԖun�ȴr_nQ�R����m{pV�ʒ��EV1S�EEϑ�e���X���zwK�ޟq�W�zc��f�ؘ�o�����צ�?G��fϝ �d�Ϧ[ Z+���aU�_�,{A�w��}k�����Qw��M�+��y.��!�-�ɞ��UH�Q+԰�-fF�5s�X>�hY�$b�z��2�a��˩���X*=�����p��2<��f@O�"������9�w}���"����ѵ��ǣt��������\G�~ ;�n\�_<�$y����u�ra��Y����;�s3�n��ͻ��Q�9�}�Ǔ�y�珤�D����`S˯Q��h��2=ˋ�W����Nz2 � ���v^�����^�)�����9ؓ�=L�q������Q���W�)�{E�����dM]Ƿ>ܽ���_k�k�<��Ʃ�k�'f�am�2��ܭ���u��r;}�. �xM*7��=3�ܜ�Fm{������`	�:�^���KS��xK���/X���F�)U��{����m�*�r�8����1-r�46�u]�靔��О�l5������ƪ���S���(��e��.5�CD�:�
p�ry�G�Nլ�0׺�ı�do[�P�K�MG�t�����z�)�f��u�z��]������5?V��83X���_�׏��~c߇K��@�y~�ۭ;e�W�t$3� �W@{�)�E���۷B���Z.���zd�ñ;,e�m�@_8��%�t���&��j|πޛ�*�G:i:�V�������v��'�<xd�kAU�uO�n��� 2��5E�8�=�Bsq�G��� [����;u��\<��(��h����'Y}���^�/O�v�g�V������dϑ|Hmq�x��~u�z�>�{V'\m��k�kb��)J_R�
��0�X�f�%�"�"����D
�Jg	a{e�A������h9���oU�Sي�Zwܩ��T��)��?Q�͹�욌�1M��x��چ�x�x4|�m��b�.Ǔ/\���=I�}�ݑ��4S����,���-ω`{g����n�KP��|=S�H@�ָT�=�R��PѨ��Q�~����Ogb=�:+����g�e���7�����Y����5��z��ρ�Zs6}�}��u��>���(�G�#����Ȩ��N�����^N�h���k�|TÛ
���ˋ$.ʞ*3qT�E����Д�z�v/�y�3��{(K܇S|���`Y���*���T��n��HG�&c1��h�nn��<�E\,+�}N��0t����F��=q��]��Eg	�+XS)ŻCq-50Mu����@�~?�R�;n�	�S����Zw>������]L_�O�3s�V�ѩ�r78I���%�wg��ǯ�s$@�9���ͬ&&"���z�ú�)�X��V�Ų쩛�Ԏ��U�J{q_�Q�K�X��_'~��D�S�5wvo;��^�U���{X��Wx\�Q]��'�gP���Wg�D/z����ϲ�o.��z�������׍'����?���{	�����^��DϺ�t��PϵUE������yW�� �Ճ�?�E�z�;���߭[:��V�(����{j��iAt��Ł*�q�nk|@Ϻ�^G"=�ۊ�򣆛�{�n^���1|�����pu�C�?}>�����8w����q`ju"�{=02�r��.ۊ��m?dX�����k�`-�.��x��2��T�:�*�2�kK3�7�w�����`	�M_�iV�
҄z6Fv��~M�
�����	��1��[7�zJȪ�a�R��γq�>	�uHc���z��y���f�n"9��٧���4{}����=��/��
rY��Z�@=�+Ҭ��I5�{Ż��D�ͤ�I��d�<�Q������R��m87_՟�^`8�]{�y�W�QK8v��"Q�\$4�/muBx���̭��:�����"riF���X;co#v+C$�-�2#e���*C)�xc��G[��m�:,������כ\dp��!n�͓�!��������z��b8�����ujجUA����yPf���H�Oa%��_�b��T��D�ˢ�в�����=�z��O�q��K�s���#�Yj l��e7[�B�B7�۵Y�u�7�[�T���`T\�3Y��
�t>��m��/o�x��[�}>M�'�����V-��ܯl���K��oDUH��ex�9\����U��pv���{�<�o���gv}�w0�Ű��9�w�fD��W��g�O���U���O��r ��w =_B����Q٩��Շ7�M:�N�����u7��HjG�홰a�����~=޳��a���*�}w�-f=���R�C���5�p���y�
��`�Xcr7(���dY^ox'�}��|V��Ba��)�@�D��b���+����t)k�r^_�sX\L
��<�q��3��2wK�Y���Q����'Q����zɣ݌��p]?
=�=Ok˕������/�슮��ݭ�2tV���?���uz���V�����Kt��bϩ�֏ӱW�ٗK��������fB
O��>0/C�T���ܣ�»|щIU\H������lüuBxS7gn�COL�c��v-��|b|�z�}��3��G]͝�WuS��\v�Zy��be7H�(:�G��|��ש�}���bk�W��_�q�y������X�� o���0���=¢�!��L
Gy�J��_%��L�s�/}��\/i��>��VUC�Q���=]f�� k�����θS�P+��/k��ޭ��������C�G��B��K=�>�T�b�UC�=�{��p�j�U��>�s���GL���?_�������p����߆G)(��)YU����Mm��c6��ޜ���V0eB�L����x��d7|]�?K�H�{'�\Ҩ��Y\�3
�b��[K�z���^!���N��ʬjy�Qr�b�e����D��4tc�J��t�!q����X�D7>��-D�^��Vݳ�z%Ѩ����H������^.�i�~��vý;�D��}�ɮW@zpߵ�P��#����2��fT�R0TJ�,9�-fmCC�8�Z�c����gG�^������@����ǯ�챟zY���\��$�n���}~��uש]�]��xjd(�铻�1�k���u����p+#޾ ;��ȨyT苏:,i��v-��I�����혾J�U|`Y�\z�h�/�ϬSsu�ε�v�,iOz��0�-zdշ��э<��;��Ǧ��!�Dܔ�[2ڛ��۶�^#Uo<�]q��`R7�NK��i4؉R�7�\}�r�W�j����w���'.+���|ƫF{�{�l����wND�5����Y��I>�{�*�˪�)���U���J3�NO��YW\7۔C���Eo�|{ ��	����Ʒ�S�K����^��}�v�=��p�Q@�����.Ͼ���n����X����Qu�X
u����D�Z�z�f/��߲�Yy�;�B>s���s�. ��Y�F���Q��ތ���6���<���>�Qyu�̦�to:&N��׉�z�m�3c{т~��83�=� i~�^5I�%�l91���(��Qs�u�	��Z�-9�q��7�ݺ���[~�V���7;,f����z�(��tr��Pœ��y�z��@o����9�S�޸H��x�*��g��{R;��N��p&D��;:���=��D���U�5��2gT�ƹ	���|v���Q��z����j#�n㺷6�1P��{5�K.�t���>�ϧ�Z
Ȋ��x��dγy3�_\k�8������'tR�Mי��V��V�}�}X�7��0��e�͢��UX<��L�d��u<,mϥ�N�`�Ls��CU��s�F�,�H�$�����U�1�����@��>�����o=	��]�7u3)h)�[ۘ����x�8}s�;$���N���f�N����9���N�,�4<4]�2�p�<�PZB�xV�T�ڽz+zˎg�[<&���J���n�mnHMW���J������wH0�Q��}sne��"j27 dE�^.��}/^�q�J��݇Ř�Wy�
�>�q>پ�4{���UA�cd�>%힣#2�O*�!9[��Jԍ�@�mw����h�_uC�^��|�%�o�t_�ԍ��z��^i�-����y���H�V�p[�&��20�����4�i+�����Ǌ�Q�zF�{r�����U�g��<���QИ�񽘔dVYN{�F}Ҵ��Tw����u���;^�ήo��xX��UfO�y����̃O&�.TKG���\{��&)��;��{ 2�[W%�{�����p��v��W�/V����(P��K���yOdM]�܍�����kK���چ4�y��-q�p�����^�,�~�<�����(	�Q��Ux.Ϡ�X���sj�j�"�����s������ڏ2���;��ddr���3�z!�6k��IG/�D-8}��)�v�	���mhw;[7[=&�8�&z�������ޟ#q�ݸ���nt��p��r��4��ݲ?)���.�js�=Xq輥�Qҍd�͏�,�\�8n:�=/ �?^pf��a�۶��c����9y�0L+"!��^�j2J:�Gs���Du�+�iv�7y�:[���VA�-��S�j$w�UǶ�З�O��1��H�l�N������J�f|	v}B|4�{�ZV'ƹ�����s�>�L�{�}�Z�':+�=���ޯE�eo�=�O���ESQ�ZX�wǵ��H�nu�Z�n��1�e����}�)z�׾yZ:��-ϼ��1x��d��f=eb�c	�{&|�\�I�Q�`t�-*����i��ϸ�����]��{��z�)Rp775�z��)��	>ꜿSq�я��������qu�;�{���89�Lt)�,���-At�}>[���s�u�X�v{8�Pc�{r�U�����eC�t��|�|Z;�����U�Yj�E9���W�m�UmO��G����R.���+�ϙ�,*���~��y<��Ht!��:u7~�r�tT�~�K`�z���'ǖ��>�g��x�w��dco�zssӖ���#�~�9��6�0[�j����9�x�Ȋ}^ӄ�wpKxk!yF���W��Ew|����j�'�����=�T<�M���A��>��s��14���/1k�3��2�'�5q�۵Zv���i���G��ƒN��+�n��7{�餏��][՘�R�rC�����Yŏ[��;r;W�m��$�f���踊��;̪�qf�PwX�e�V��LIC��yҎ���
�.�q BU���R=2w`�Y��P�>�f�P�C���{l{nj��#�u����8ԺjٵQqf�����]�'�{)I�+J�q��j	���h���J�����s�.�>
��>������9>ጙ�ў�����3��3+K�wP���v}1��t��,z�`JUW��S�s�ԅ�}��#�N}�]O�g���u��_ѓ���?�����ǁ�����k�O�!���v���zO���7f����[��/��	�>�Q͉ڇ�^����i�r���`6��u��������I��D�+��y]�+c�X$Tg�֋^�]���8�a�Q�����{��;0��f�W�b�,��R4m�v�9����y�!���R�jY�V�<���3����JArc��.�R��}T���,m�?_��_����q�W�����:���DS����NI����RBCa�s4����FL�L_�3��Ȅ����w�>��~���V�6.�D�v3�k�̅������5�6S�"x�R�EV5<���|��-�ds�㌴tg�����g���±zR��T�𩋢�nnJ]�9���Mn�ww��p��"#�+��gN�7]܆m��0(G9���DM���&�¸�����)r1;q�}~����+��v8���}qƆ$�4ُ�k�M�i�+]Z��;�A�΅�"�+��[�mr�n�r�Qئ۳�w�*Y�ϟ
vn� �"�E��d
�ԯ9�,%�﯇���V��ۂc@�3Xw�-	R��Чk���@�~�dxq�j<�L��IP̑c�W�a����HOY�9OFڍ�B+��lxz})�{}`p�e��/�{����dyΒ=���#*Oq�Е{�z�:�v�v��2�\}�;�c��.��+��ԁ~��TDú�Dy����_X�hp�� �;��`C�_����>Ӛ��9���xLz�>�g�x�ND���t>���qy~�k)Fvn�w�DzQ��+/ó��#�+L��;����C�S�o�+�(��Z���U$d�Y;�϶���@T=�%Q���"�j���ѓ��k\�3�Ƕ�,	���|�7n��;35Mh��^��o�C}���XM*>��w���ݳxa�m{�x�3Ap�|Z��i]�W���G��Ѯ��dw��"�g�Uǽ��q�ע�&�͉ڇ�=�}�^#"`��,�6����^�>��#�}H?*�_%���s����;f���v{�܂/ۢ��Rt`�Z��hE�ȋ*f�%,���\k��N�����ܕ�a��9�;�l`I�b,׭��O���7�E��05��hY��V{���h1÷LW.�ȉades�om�M��޶)E@#�,*A�ԍQè\����H��;��wKe�}+GF^�u,��B��5��;q!,2v3�<�/z��6-@ǋ	��W6�}cKErDf��T[���	z'L>��v+���c#P"��8FR�*Ŋ��k�2�n������`u�̅\�ۆQ�� |j}MR��boTwj���<�E��2�:f\�����٨o�]���u��1@9p��v,�N���>$Y���n
r��B���L[��$k�]ȃd��\2V�����5�q֡�{%BGV>�ǹP����f.#l�uk�4�J�W�K*b���p&š���l�H��1ό�q�.uٴ�խ��]c�r��e['-]���]CP�P�g4u-Bó�>����z4Y&^�#�w;����m��u���"d�:wQdu'������ث�z�טۆ���wi���Uk���\ê���`���L"��eޒc��9�Dn��Z��2��OZ����V��b�p:��w\Q����*�����t}���3L��<��稔�Ƿ�n8wz������>B��}uv��.�b[1��H*fv�M*�9����n���zH�df�v���
C�1��޳�n�,�E�xb�����/�<�v�c)�Y�R�%GF'�+'@���)�-�3��L8<��NV���Z�Um�cU$\q�9p���ɩ����qbu��hɼQ�4����a���$DȖ�<-�¼��4�=K��L�K������Op�H���Mkۙ$|J��=7�^��<_���Ԙ�ԇM��F�6�=��A,;�8@<���X��vu6#�Ut3��m�6�X���#�*��C�fP�[oq�� #�T�N��m06.�Ρ��(�A����!�+Z�؝NG�H��������S� -������{��Ťئ��Ή;�s��I�VM��i`*�E=��Z���b��Ѷ��|�0��s1�yR�����qЕ.��Pӄ!���3���E+�(zNgqԂ�_f5��3V_Z��\����� 'e���c��:��ʂ�����ވ�2���3����/�b�T��9v,#��<IF��.��t6�k����=�pU�k��LS��rr
�#��4_zh9܂&��l��y}I��qvby�gE�8)�s8��z��Ŝ����/V�<u;�5W�d4��d.x��I�/���(����Or\t-1�xI	��,Wk��.��}y�Fd�^;�!]�H���1%�+����&E(bK�P�%A���ҩ&)%i�u�rIbP�
&f�2�����;���,&�)�pF���R)�$�J0Cb�$F�Ȍ� ��&�IL���F2'uѻ���13�D�HFA3,I˂'8���d�n\�&�!!4%��4�d����4IL��wt��wp�J434�;�&��"(�1FiFE�(�C2�"@���6���L,�1�4҉	 ı�1�wvi �&1I�%$E"P�M �&)��w0��4ĘH����0J�� A1�&\�B"c(2����$#L4�X7+��#1�2��E��ׇ�ö�'�REK}��:9�]:�5���{���Ѓv����Ի��[�q�)����\v��g9r&�b��*(+�
���0�H�.�Y}S��.��q���@b�Y��Q�\$o��F�y��w_�V�nw�W��	�����_��3�vNzc��Nx�����|�;EE�{�Eq�9�&����3*
�/������c����{Z
ʫn{Ō'Y�}��!-�l=���{8(wazv*�<�V��)��a~��m�]�dyQ񎿷|.��6˙�O"_�3q�,/w�P,���5���V�7�l�z27�>����^�p��1Nq��P��%���j2�7@L��K�b�(̻�w9��u��5�\Jr��÷Ѿ�4T?_��>�[e��nk�(zo�ׅ����wgT`��s3�O�/D�\
�缥�mCF���ïZG�����D询�n�_�U�-�f���!�ٛ~����>0�옖�g�22�U4sai�/Ʒf�v��;�9ģ~��k�4�o=9����Fz@�yӒG���"�\L�9����;���p��si��7���{�2gs�N⨝�dϾ�8\/fA��Mz��Z=�O��ݳdĵ9EF���τ���������F��i�$[[�C��弈�����й�i
�;��[3��:}OG3�[�
_n�1sOh��3(������o;5unN�=�M��1ǌ֗����3k��Z�[� z e�c�.�u;> Wp���\V�2��c�v�y�P���6��n�g,pDK���ݨݪ��Q����g���F��������'˘��n������ü�t�xEڣ���Tn/WGd_��QU�\4zAC#UQ�O��AuC|q�PxjQ��W��Uc�C�n����Ɍ�E{�^�|}��F�{ƕ�x^��Ƚu��߸��Z�A���-g��[��WX�Ez�v\���5��������2v�oK��^��<@�z���n'j�[�~�jF{R���p� ��ʄ��;Le�֕y>����M�Ł����{=0&qH��7錡�E�ȵ���W>��qF�3�Q�� ���}��Hc�K1����G��u!��GL�Č�X�Ā�X��`C���knp*�����<��1x��g>�N�*f=g~�t��L�-�'�z�}��a�Elu�H��Po��G�����|��w�,w�]��}�(r��)�f�s�5�W��zg�^�FW����g��y2���yP�z]�ӱ�#�=�����*�F��!����S��ꍸ���ܣ������>�6j�rӛ�!�9�w�I�}'Ǹ��_����*��*�"������ �hA:��Pӆ~м�'�����e�7�cI�5��n��:��v1�Q�ȇ3��v���i��QN�z}��B�]u �Hd�i �ԕ�gqZ
E��F��oyb�:��n0��uN*���f�2�"Ϧ�pu䝇mɱt�:Q9Q��н�4(�Bg�΀}2EdK��ϙ�,+ޮC�6cǏV�\{np��P2�Ա�7��irX�LKf�bX}�R2�ex�9�����W����s�n�q}�σ���r�Gӑ��5�n�F��sp���3q�����	�����9�waAQ��V�߮�����h�}�o���ҫ�>���נ<�]�~�����nG�c��Foš�]�����S+�G��=�a��>�}V�~�=��`_���+�@l�+��({|=v'�rJ
��`A��e��l���=^��Ba�Y���	��2Ǯ���]=�q{�d��]���\���r&���6�<;�=��ft1�wp�5ULk�IӪ,�n���h�����%1e��D�6o���U_۟߄U[��\T���w�~���X��	�+�M{}�������խ��G�v�O�dmw��0נOi"�Ó�W��q�5��� o��Lb��V��<��&�¼��6@�?-�D5^��oE���н�{OO�aՑUN�:�:�-M�V��IkZn��?)C�:��R�\:1�֝�2�oe�dT��n�.;�����-����I`��߆�&[��vӤ9���C8�-ϝ��3�M�h��y�j��=.j�pg��`SP�.3-�Q(߶���5\A꠆�:~��<}Oգ��w���>�c7D�����ҧ��ǻ�r�)���w�.W7��/r���람.f�X�k��>��V��e�q�^�|2<��)����΋�YZ�yGv��9��-x�``�*�	�����Nb�&|�<m}�<�����}�;��.}k2�~}�D�z{��+��ʕ =��2"���ϑb�ɖϲ9�qe����B� H��7f3��f��+����t�;��u~��+�f7�|)ٳ�@>Ȫ�u2��J�u�L+��sA���o�ƪ��3�4%ʐ�yx�Eo�;����
w���i���̨�H���K�X5ϣӱWY;cA`C�9ޅP�E�q�s�H�l�+�����P������i��72}2E�3�De��9l?D�o�s�Z;�c�4����x�N���� ��Ƽ�tD��.%��t��t���L,z6b|�dVQJ{N��ӐKÝ�1�}T�&�}'�V�
�8}2��y����׫֪x�ղEG���:}u��G��27\�@b�
�P�x�����r}�Ѽ��^p�L̑[ҽ_��r5r�F��G�͔�od�C:��V���eCxB"%E����I^��]%CB�<�ڻ%��%�L]|��4�8e׆RL�U�W���rH,{Kns�
n���Y/yi^�PF~sV�>!ϳ�ݛ�@�I+��,U�w�a�j*܁PW�9�X����l^��.v���*!<�QTr�|�dD��=ͬ��2|:MF��f�i�Ý�\zst<]�+R-�Al���{�5���i�0�a4�ߪ|�dMuǻf���ͯqJ"�j�M7��HE�}X ������#\������Ѹ��X.;�'�\z����	�Ty{پ~��*	��wos�ɮ�w��ZoJG�㩀&۰.W�|F|�xO�k�_�1��~{�E���@Ñ����|Bg���ˌ��w�d�sq��o����\�	V�<}^�Gq򾨫�����s���U��=��㒶��Uxf��&w��'<�o?d}^~���8���W���&f�F��W��>���>�E�K��ȗ����������b�&u����/:d7O�����|��/����D6-E{���F������^�n�\n{�g�F�U3r�s�U`Q�@���K��T�U�~�E�d���C]����D����Fz�����Y>�bh�ת��Tә�Ț���(��g/ߥiE9|sz��VW����"�#��'�{#}@h~�W�)�,��l�禺�[&���c��Q�J���ұ�(���B�4�7҃8�)=WN��C�۞�z7��<w%H��k��/2s���������v�����c�/���K����j&��|����9o�O�+*�J�,��_gc&��V�{{�/��~eN��T\�)�dmCF���|���ߏ��L�G��z�tGF�|�Ϸ;Һ�_�Oy���@~;�28��7�Ndl��}�:���zgx�]3c2���a��4�3vJFX�~��ʧD��7����f������Zv�w���_JB�� �ѯ��y�Lx��i���t~W}쫪 (���\yf�MVѿ�χu��8dK%q3A����<|G{f��P�����C�r%����M/x�
�T<�L�C���0���L<k����s�W�O��8�t��H>�'����,<��x�\����Q����]�ޒ����@2�Y7���Օ�[��ѽ�i=��= ͈ڇ�J�5L�Gk����ϙʛ3ּ���>��ݮ�`�6_L��</��G�읭�{fx0v�dy�� s�T�uW/� ����}�������O�c�q{ޠJ�l��;Le�֕q��Zn5��M��w�,�[N�D�E�ϫr.3�^�LF��)�ܨ��T�����O�aՑT�Td֖/&w�Yb�o_��N@�F'4��'8Q�s�<W�5�]�͝<��yԹ��w�DG�՜Vgb*���J��(E��n��z�v^����^���&�x��N���]���Ɗ�ވ�^�vb��0v��&�h�h��j<��5#�K	x	�y�\-*�(�hu�twt���/Z TE��o���tu}�;#�l���g"};����a��]11^
^�++��+��p$纏�2ǽ�C��~ӟo�y�χ(uv���{E �ES7.p7;ڪh���j5�y���ۨ�a�3dς��squ�;�{�{ۄpt���=E���4��/U"N��T����C��tȠ2��_\�9�Cjv��	�)������7W�&E�	:8q���|���1^�j�>�$6n� �d�.XS>F������6�M���9d0N��ݓ\��>�>�9���P�2}%1-�ىA�UH�W���+�26|�sԧ��z��;��/`^�W2�}�(���w��.$W���,��3lĠ�"�1/����l:R�(��tE�T��87ޞ�Þ�g��x��_ �#=�T<�M�*%��}$/t���������Qʠ^&�]�:=��z�Ɣ�v|&���^�5V�� � \��<�] ����Tc��Q�� �SE�V�(�)��Ua��!۝��}��o�Ҥz�F���@y�pyˈ��v�S��������a�Xɒ�~��w"��״d(��m�KS�pu����:��ovr�,����Qu�N��|�}���F��+S�kNv%��e�D�N�R��o+�b�[7fYn.Ǔa��پ��
�a>��'��o���3"���u,i���Ǫ�ÿ����¸��9Y��T�4fz�3�cՇ��\&���~�_�S�ǲ*��͝�댝����f��`MF\T�E.��v��s.*lR΍�E�G���s�7�4��6cc�{MǪJ:qW�U��|%�x[��<�@�%��rWxi��}�U�O��-=�p�߼Z��;���=>��,��x^lw��\7S�����Ӑ���/-�Y��H�H������o�ka��/;�4{�Oy2����Ǚ'm����(Y�<�7>�>Q���y3����	��6�����S/�u�_7�y�T�4�hU����FRμ���\�`��+��	��\;��Nc	���2���_���>���y(d��w>"�mF}�}�j�r��+#}DS7� �>��(�#.|�Kg˝`~���%���䊿+:=��v���q�^��
�Y���]� '�U"�&[ TZ��뼎�ҽ�w'���
���hb��;c#�J�پ�6�����9
�*��ϱ-��H�3��V����܄�ެ>3�c����	��d��A�Bj��S>΋3������/�+6�s���,vق9��#o^WRv#��[p�(����\��u�E����g oϤ�Q�:�G.�XT{Gyf��-K��{�v͚p���G�A�oP���wRr9"4��R3vok�)�%~���y��a�]ŋu�H��R����g�ף=>5�.hy�^�<��"��ɘ���C��
����:��t���L?��C�u���ӵ���z� �3�d~v��<x��92��М���ic�1+ǲ�����i���%��
�_Ϫ��W����{"���o��$+X�ܰ*ܺ�.��눟e�-�#����#Y��Xʏ�
�Zo�Ԡ�����ٌ>��Ӈ����wu),�t3t�Ϩ�إ>G�&���}��]����j5΃7�څ�����,א�#t�:<��FD?H=>fC�C9p$� Uz��P���FV�F[����Mg��w�}���f��� ���x\F��Ƚu�z�ު<�M�D�r�TQ��Y�+��(V�מj���0��Xn0�zo� ��z���o�Ϲ��J9ܩ��hDm��l�߽�e�k�0��NJs�pT��(k
���G[�e��Ns;
����7r�1��^Kl��47M��+�߅�O�U���L�֙����vzs�s{1�y�@����Aؕ��_ï����HI[��=o^�̊�꠿:JY�<�u��2-��lJl�����>����h��vC7�Ց�6���N`۠W�^vu[��{I�4���׌B��oV��;�۝v>��[Z�=~ݳU�.����=�c���f��	K���=�������X�u�'�\���K�FgԲ�;����R6=����r"�^��F?e���n%N"�*�	���c/�J;��EM��B���e��]�4�Ve��G�^�:�w��EP�S(��:�!�7="���Y��<���}�\ks޸x��Μ���F	�޿_�t�}V=~�x���{��u�+L��%��d]DO�p*.yz}Y���ߩ"��J)���N��J�*��̽@�������"}q�@�7��O3�S#*"g�n�}�������yZ�I>����U�WZᶨ�����i_�H�wT����+f%�U��=�I�9��b��<׽�-J<���{9��1���O�n����y5� \J�h���ۇVLS��'۞ޟ
>�w+���4H��	��e),ZsL��@���Ϊ ���_K��+"j����k�q����%ܹ>´����4T*�w����܋����yE����{�ǁ�c6�FA�*��*!ťc3wU^�(���π�n�&��� 5��}I��O�`N�ޑnU��������9�]�t3Wb��v�V0u�%)ͻ�w^������>*u�#�A�$�y݀���rU����qkۡj�u��-���Ӯ���:�639�ɴ�h��޽��SV�:yh��(|��=�f�oHQk<�ti�%�r�#A�g9-��U����P�� v2�zy��7h� Q���|�&α��F8Q�n�d��YI�ͭh큝�
�9�+���c�em�\�*�X��Wv<%�s�/�Ad7�v�b�����L���mK�k�`L�p˼86�Ԯ�(�)+Ԫ�6R�W�f�!9�� �����2�a�U�-��r�'k���*��N��!�ӶL�+c����VaiF`��m�ÃKމ�`Ŭ[���+WOX<��x{0j;�a��M�V#ka��>�p)�;�w�,D0u�ܔ��Ɏ���v̙E��o���o�e���yՄ)���!�p@�a�wض�R�,�� &L�Ҕ� �7�<ۙ]/��3��,�Ou�hJ�Y�fT�	�5z��F�4^�s�jN��`��9�YER�h]z�β���psX2��<�]��-�k˳0;ȡ�Hޢ�vp4<����g2Ύ�dʖ��ʅN�h�aÔn���h�`�o �lS�/���R����%��.�$��݆�}��-p�g+�	[�@��id���T�c6���է�w�p:��/x�iV�.�A���m�"�������о�����5`���7;o[LH���rȞ�ڥ܋���������1��z]�ҤUog+:(���(����>����M_45J�8��g����k[|-X9�m�]�[VhoE h�}��,������V����R�ή��v���s�նXI����Ţ51���:�>�4���N��[�u��[l�(��K1N�I���G}II��۬s��Gk-I@Ջ��0'o�k��)D��oײoW��ꡥ\��%��S���ӟ0����ܴ��y	W6�E�I�sV�]��hm���C��׼&��9A�\cǤ�E�$��� ��V@S����7���qV�(��o���G2g�:hN��&}g$��1�k#��J彷N�ܥX��o7��" 8关�L�m���j���D�i����b��.��Gh���������i'��%c�����T��u=P�7�'�^	����>��R���(SR0�����@��=�K0�)Z���lSػ/����6��wp���@!�<��cm
�Qc��]�NN����Z6j��{���-���V]�3%��u;Rk�o��I%�:b�G<�S��WZ8���ף����cZ�/l���y^V!�B+"���띢#���w�� �ݻ��\��+�wd�V��5��0avMfWj�u�;�|?$�$#�A�RD�i�(F#�ʁ�(Z���
���1� �)�3��f��&R��M4��КB��Ĳ�i%��X���IH�Np���!"J�L�FXa(�.k���%�	��@3,e��*2��IF&Mf&$a�";�
e� ���Mk���يa�L�Ai��Ŏ]i�L!7w0�)6(�M��f�
�3	@�d��*�DF�&
�TSI,D�c2if�1�K!�H�$��$уd���!fc"�1�T�P�4AnW(�Q0��1�BJb��2M	��1����Ȍh�Q����Qd�Q�(�R������ѾV6�Z[ck 1Y�(%�v�N3�wW	|Q֩���!�;�[�j:8A]�Q�y�6��@��[�v�L��i�ʅ*O����v�a�f�^�5�ƻ3-��T|oO��~���OTّ4�{�5���"��:�WE&�g�|l7s��zX�5����d%5���~�Lڪ�>=4�ɋ���dM�}�Wr�2N��%;1Y�ϴ���7��������ٻ����v���?e���������F��ݔ"�x'p�z���ʤ2�&������Go����>��U�%��%�ꑻ=� �N��q��w�t��ym�b��b��s	쪇�Ќ��>�mJ�m��I��t�f��Hco�~�i��:�=��\+���c�G��;Tҝ}���������@T%](��>��X^w�'ütG`��)�g��{/Å��p��Iv�^#�4����ҋ��&�z��*"�2�{=p	�P(���!/K����n9���>=�3�����.���a�z�<���d�A��"�%��P�3���h}��;�o�:��1�ٓp�x���������4�n��פ��eF̠�*�e}2�V�.W�hb�8���l�S���c���䗭Â�h0�
RחP�xL�Cu���4��;��R�eֻ ��;�q'(
��68�E�l���E��6~�j���s��ZN@��?'�݄��VLۮ��yZ$n�a?���]匚)�b�Һ�x���s{���Ԋ>��e�	�W�a��7�z@�G��&|��B�\�y���늯�j���\3n׆a��������Oq��;^g�x����ِE<�P+ʃR�;P�\Ħ��j��99�V	��N�g1@�xk�'�p��0l �=�`+��zj�����]cֲ�s�R�AUc�r7(�U��M}���/*���6��"0o��BS�^�L_�o���[�<��i�㫗����	���3:�ª�A��ݼ�*���m���q���$�O��8���C-��S��Ȫ��;>��5p~�z��3�F
�vx�>u���G�g�28g���x���FVǽ�8c� ��L�r�*^W����э��zcng�[�>��E"�<}��WԀF|@�K�~9ׂ�v�
���Z���9��Fδ��#ڰi7}�m1�8|�T+�WY�R�����`\ru�*�=ZG�_�v
�~�(�������g����zYÓ��Q��ʨvNzv0���׮)�{�ˎ����l9�&�;] g�����܏h����f^�rqH1n�,W�hq��OZ�+`�e~�<ks�1^0��J�eF�o7r.F��FɴqobX7\Xs1�5u���u����>��r�e�}����dꖛ%�n��=��L؁�Y�{�УK2����ǻ�E�d����
��3��ÿ�e����9ϴ�J��=����<}Bs��;2r�����	87���ꍸol����L۩a�}U�LT�"ϑc�e�d�1�ura�~��Un���)��w�z}��L=u(���f����b���U^�������l���^���� �L�N����dxd�#�\��b��f�5N��f}��1�>��4�븱p�ԑϟ��#}`p������W�åi�ɺ�+��{Q��h����22�y�ß�ۈه�_rJ��Ε����<
�zn4>��}��},��w��o�N��������}1::��G|s~����?��eOڶ2e~�Vº_����3pz�Y�}/h�~ˊyu�"�U���_�dnQ;�������G��j�ȹ�u����E�W�c�	�\T}���I��~��Ϧ��fއq���l��?:|2wC�瓱OW�!O��mDzh�5H�F��o�hg���6<�To�>G�j�ڷ�^��6��u�� P���%�����W�~�����.����5giA^��b�qw�[o�����M'1.t�U��wM+t��v\��|�׼��й��"��ַi�{x�8��O�
s������[�G�w�A����f��k��\�E�ۜ�����[�ءI�q�������3Q�O�^��TY�zO/z�p��B��QgP�W�)F�v��ER��t|t�D��a��0���~=7H0��	z��ds����n�'R~��9T�7=��4�G������#�ʥ���[�]-~e���J���@U��'8�F�<���D�5�|��dZ{Z���x�>6�c*2kK�ɝ�����3Zd{=�lΛG�QZ2��%[�3�B�B��)�;~���d�l{���S�R9�g�Qs��x�y3��F�Kޏ�T2���s��{4�L���_�tl}�>�����p���G�`GV�h�\T���,��zn%�g���T��#e��ɔ�vX]/ף7��=�{�����a�{ޡF�+�4s<Ҭļ�}�[�MF@���3xaq��ިw�H�>f�����~=r�����l	ģw9wa�EF���=2��rd]JW�yz}YPѨ��u��9�QL�g�c������~!G(�Sp�{=j�ײ�%� 6TlĦ{>���3�7`��9���k��q�,�~�?�c^��m=+{�%���qܣ��UwR7?MUv��[	<�K|l�Hv�p��+Ǵ2�m�)f:��]��l��������¥u����>;�����5^e��N\��~�\QV�m������`�^��pA��l��]��xI�B��:_\�P�.��|_�'��m�
��N�\y���X�p��vJ~[��a�7?'�Z�E��鼎Qg������jB���9�/+�����
��̃'�@ؕ�1�ߕY0*��*��!��_0�&W����vW���,R^�g�),��]����yO,\��ggq�=V�~����
��l����4W֬TTF����=��E���9@���Q쬼���d��+�f}�vA������<����Q�ƾ�b�U�s�x�.rN˷b��`	'1g�7�r����D�r�T-7���zp:�ʮ7X�:��N��T���ht����9���D{Χ���������	�3��E�����k�xfy���x0���c
��j��q^@{2�L?R�01��)�̨��mȊ�{n��Iý�U!�T�X��T����?~}2���ds՜��R��nu�F�w�g|�G_����%VѦ,�s	궽Wh�վ�｝���z�C�ɝg	��m����9��ב�eG/U!�c��H(X��'&�?Rs۰)�K�Y�:nJ]�+�f�����
4�0�[;��ʅj2�N�7�gG\˧���v��c�c�����zoz�Z4�f'6V�J�f����GZ�kw���<��y�Ik��x!l�4� ��k��DZ����y��c������ۊƨw!7qd�#����y>�������+]C��<��L��q)�1���9�_f�s�؞��˻���;��g�J]���y�
Fx��G ��P&�\���B^���5] �ٲ���nv���޿^�r��N��^�G��~
r�7d�͟:�ET���L(y��C���&���63��/v�N/h~���1�W+C#�Y����z6\�˨��D��;>�^+ݎ�r�'��*+��vzX.Q^�L*���2�x8���s� gD{.�E/S���1>f�bP}�v�M��mh��]כu~B���S .��|����S��Y[^����pD�{�f�e/L��le.�-_�K����G�N}X&&)uh��΁0��w��S}V�As����8���:�|�1�mm�� sv�O�˂����C��l��K��|^�P�u	z͙����+$�ʹ��>�K�pyPO�Mu׬�M�e}��\d��ke�2kK�Ɵrk�����=�{��L{�$��ު��w1���^���O�{#ꮿóv�U�����SU�xU���a��tQ�4����m�X��O>����o�.T�P�^h��oKr]x�M�b���?>	�a]ke�P�ǁ�my�s�h=7�o�Se����LLP<��U������)T{F���;:��C0(�$��7���;�؁�I���u�ٰ=�Yb�P+�u��页oۓ�-�@�,�G.'*u�{l(��2�{qO����ǣ�5��4��u0'�4�	{+�w:�*�=�z(_��kB��"�tg������4��"�.��n2�����Y�3�> b�����w�*�85y;B�?B0/7N*�$����/��[S��*�iS#��쭸w�;�.f�|6���P�S=�{r�J3���xz�_���5g��C[E�mK/%֍eU�}ꇱ�:�0�S+�2���:~��J.�Eo�O��̮;��mڨۏyY�Y��)���Ü��&��s�X�[1hw��;��s	ZF�1��_�Yף��p\g���sޟq�V�%���>��T�'*^O�˩��3Vf�7'��e3�ﶼ_�C��C"	�ȍ�����:��2�5��E���`��s�qwEן���=;���/��mCUj�,d:�6s�x7y�E<�t6��u�@7�_8@x��s�ׄ�Gy�Ӥ����FFTK��8KGs"6���t��u���'�]��N�8yJ��I��$��ժ����GwOBq�ᦞ�J�0��P�a�}�,�w]@���ve�M/U�R2�0�����JM+����V`u�r�j.��T���3���6�D�wm�$[ͬ�A����'v��	+�[�C�&�]��Ԧ��GvYɟQ�Gŋ����dEe1N{�r�;�	xj#;ƣ�c�c�r�\��r�^�>�L�5&��Q�e��g�Fê!����/ór���+Mg�w$9�ᗖפ�u��H�YG�Bcj�ۘ�s�S�.v���4�^�J�#�5ws���u�<���(�K�['��WHmD)�X��c��C�O���]p�Y4��ީ�=b:�o_�]7޿@��Sxc}��7灚�i�U>�����>'}鑞>��b���sSY&�&9/]9���e{�>:vaYߣ�{6g㲢:�mz�9��~�z���'k�9��	(��<o�wHe�,3U�t_0~Ǟ���t^��zX���f�@*},c!׷gt������[S�e��Nct��vz�ݶx�d��=��'��c+&��'}1��k�ŧ�qˆ6�ެ��W�=�s���7�Tv"Σ_/{VG�QF����x�D��*�FJ��Vߘ�I�*`�זvg�z+�϶e������w��u�{~�W���Q��m�adkL��.q�6j7����o�бu�������QG�~;����s;�õPG��z��駽:d^3�Z�\7ۄ��ڷ��.��.'y��.���{�1��2Ƽ�P��BN�����웜ukv�e�\��D�!�{��ܶ-�L�m�{�|�����ͻP@Wa^_v�ɏ0=���c	��FL���O�K�����+cʼĪA��δ{!����D��~U��8�J�c�}R��3"����)�ɘ\o����I��|;�����^y�=5��go����cO�^L�\a)K'�[>�#+�n�U�~.�#j5}��[e{k������|�H�����x���z}%���g��GT��9��x}Ʊn#��xMf9K�L�=;k���e�3ޭ��C��%��H��ۗ"�U:(dG�'���~��{�?o�R�(&�d����wТ��w����+A���: �^*sޝ�{2{�WT@���	�t��TRq�/m����z�ɇ�*��5J��J|O�7�l�~��9.pq�f@��7�f]#K���{[5��_���������u�j4�O���
Aan�Y��@�"��]~�\��W���nnd�ꝝ�R��]�~	ċ���k+�=��j�zL��P�i]������u�'�.��%�	��^�~Y�p l�=U��<r���8��_�����a��WMƗ�d�`e}Wg}Q�k�۴�mE�r��r�Y���S�CV���Iʢ�\.
`�6-�M��A�>\�)m�~��.�0�qT]�b�s\ �A=Du��:���[�n�o�\��0�*��T�0%==�^Q���u��&q�x��tp��~��E��r���
zi���>���Q;�~��h�Ư�H�`�?u�=�	�=��E��������X+k�l�˳���Ά���#�K�p)*{遍W�J��͚����1]��Oہ�wֿc0痫P�b����nwe�
O��;��H�G��*-<�q����#�����Z�\c�O�jw�ÏTU�NǺ=
�E6M�*��j3�L\d���z@N��t섽~Ӛ��;��c�{-��>N�{�����L��n�{���sD�p2���}�q�P�s�s�aTiU���~)>�꩗x�e�}��k(j��ߘ�ﶭތ�����Q��4�}9�Q�&+����'7�e����y}gT>�,>O6��EZ���3�{�}���*�~ӔQ�t���@>Ϣ�E�,��#�j+ḋ�м����<�+C�~��c�)�+}#M?_�=x��K1-��g��U#"�ٽ����g�؊��K5�ǧ�����;�2���u3�϶g�:W*=���<�1>���b�?JS�;�����)?��D�q��KGv=��t�j���΃�ց�z������Zֶ���Zֶ���ֵ���vֵ��m�k[o񶵭m��mkZ��mkZ����km��km�͵�km�}��km��kZ����ֵ��km��Zֶ�붵�m���ֵ��]��km��kZ���m�k[o��ZֶߛkZ����(+$�k ��	`���B �������+G����H�� J��HH)T($��))I	UT)R�J� T�<t�P�P�(� **UAR[5*!��)HJ�T$�(%Jj��@�%�H(��P"R��J���% @�QUIEEJ W��Q
7 w9�)�Xdl)�ADU��&��-m�dT�(Յ	�����
8 &�hL�`i��ƀ ;   ���  wX   ��v�;7�uhD���E� [�d��+k5&V6�AkH�e%c(�P�@ER�,��5�"�I"5�P�whԅ4[V����Ma�ЭkSbJ�)��k
i�UBM4U��m�m�"IKM
� �V�j�CJVՋZ�MM���Mj&�[e�15������� h-�6�j�U��-T�p ]� �ʥ!U�d�m��B@�ѕ@յ�ST6�B���&�U5@2I	%�Р� TS�+���J�`
�6�-)TЛ(4�Sj�Ui�fiZ�հ�m��R�6 � �hI ��3�-�$�����TS Pم�*i"IT(� n8J���*4�H2�*d�6�j�VE ��� ,J"6�dU�`��(*�SM���30����
Y��dڨ�c�J�" &%EQ�� M1���$�RQ�      i��&�&	��0`��5O��I L	��`LQ&�F#"2d���d���ԂMDR�'���F� `�F&5p6p�=u��n&׶8�pȋV���iZ�����: ���Tj  �=H����"@A
��S��������x�3�#�3$� @JC���R >I.��`���9w_t�k`���˞�@eq�	���P��&�;#��
2�$0�
{������7�6�p� �t��{1�(�BE櫭�[3m�yy/k6�G�YR�<�B@˔�l[��3�1�ۇjm�Zn���We��IP���v�bn��
��]#R�;&���hh ��J܂�� 9xt٣m�!f�K��jM���ʶ#�z�X530��+5��l�C0�U�(FݫE�ț���F"D�1��6��� �PZ�[v�e���(�� Z�]e�kicm��w��TĲ%��lF*�aV6�N�:��"�ZN��(�,�B���y������K��,6�PT�`,�r]b��w[���Z��ޣn\��9/Z��ŶF��D�qةY�E"�S�7��dy%�u�	uN�Ͷi���h��2�Ի��蛶v+�5b��Q8��n��/�K�d�.����!�^�4oP�����e��[$"����J2�U�!�e\2�ܴ��MU���3f۶ۼ�j�����@�VP`�!1n�/
��v�9{���ɸ3h,;�l�
*T���'.���MM�uI���"��n�J��fŶ�-7H�#v�Tz�+e�Ӑ��T�Z��l%��J±)�Uي͠%�L��ѣ;�@�����F�Qe5S,n<�[-�u��C��Q�a��t7.�a̍K41iR�dI)�Y�����A��EeҘ7H�ƚe�m�����ݼ�kW��M�MFj`�tM�,�C�ۆL�X9-m^��Op�&��*������4Sia�n��-��d�f7��i��A:m�ߥRQ`NJ%��-�P�)n��SN]֌Ћy+b�c�Y�������FV�6)P
�a�?cYh��v48�5�V"���+fU��z�S�j�ӄ�H;Yj����.�F�H))ͣ+#����i2�f=�7��	�����xJ�Y�Y��2�5/*��5�,ZrMb��s�F;K�v��{�E�5�{�3m�Or�aQ[��Q`(0%�ʽ���j���P��#7#�1�����sv��l��F�x�-� 6i))Ud�B��*�+�;���5�ݚ�T�[-g�[3KT���o%������K4�x�b��ͼ"�V]����q1�q뢣� �7R2(e��m,�Ǣɖ��K4M��zor�5DUȤ�4��J�*݃���-�L8 i`��=�($�k/A��v�Q���)���!D2蝦 ����Z*���,�P=�R��\;��S('n[r�s)��:��0�0Z�byz�׎�� W�n�!\��0d��H���AM�{0 �Xr^��
X���V�<��p2��/ohMzIK:*�m�GH��×u��r�N���9��wcG~�QTx�&�]U{"N��Z`����L��Y�b�4]:#�6��`䔔)$�އ����;j87E�*_�+5�J.�؏>��1������ܡ)2�f�ܷ�[�U�kE�Yr��#�x��C[�n �|B)Z���������q�0657����LRbG����Ss$��2�D�Cy 8,��]b71��n���Z��W��Dvֈ��%���Sq\�m+�E6"�O�խ�*V]1h�@��4���6��R��ױ�v�L�1�Dr^\!��:-g��((�&]�D6i�����ӎ��з�>��z����z�]A����t[�Y+5�;S�Y�VF1V���Q��ca�ե��Z����!�.ĎʽJ@d�ӮW[m�Q��.�6�WW�!�f4�^YRP�*3�X4���u�H�rd���.馂�kua���ӛfc�� �՘����I���56� �F�֘�X���5�i�7S�Д5@o6��U�٨C�0̒�2T�ͽh�{E���5����Mn�0[�ޡs���v�W��k�7fIpU3jf�owv�^fS�� 3�X�'��i<&�	de���ӟ�9YDU�R���:�n��M��Z:kq8�C(�h���F�g������qT�9H܋
Zc���|,b�v���TP�/C���~[�ڹr������-4��������(��]]n�R���G�.��6�AB]K�6p�+(�R�ē6�V����vv�6�u���"�(��D�h$�&�0=yj��p�e�z��i��������E��pCrݢnJ�+۫+��T
rE�/0mϲ�*rȠ�f2mpP�ϖe��m��1YX16����ކ��M��̖@�qR5�,�h�iJqັ��&�*��v�X�JxDŨ5���U� N��������@�pՂ�͓b+�!�r��₲��	d��e%�T��������2�Q�	@(��.�MQ"�CN�C�ȣ�6��/�8ux�oMڍ|n���J$E3PW�uM:�޷��I1���N�D=�N��,�n����%�����_�VAϘ�cTr�o���t3�9�=qo�V�P�j�oe���`��2���yQQ!W;��^JnA��mH��چk�u�H�m'A&�hs+A�RXvU-`�Ln�T�pѽ�Uo#�0;�%Չ��E�Vn��dqW�{#��B�)f�m�0�z)�j��j�łzv��X��%H�<�]�O'�v�,�k	��$�lM.ء��Ѕ+�+`a��S�!k�ջ�W�.�:�9�ux�Ƶ��˥?��em��k]���͢�`j-�kv��u�`V�aVQ$�%��2+W�U��gG�q�pj�l�� �d+����� m��ѵr]M�O�-�E�Jb��~�zH�j�,eZj��t�e��dV�%�.䆛Q��ޔ��WPe�t6�2#��'j��R���U�<GB�`��'[;Ebw[��#A��ÛYQ�7��� ��4�z�ܫ�#)�)��E������gԾ����{�����N��zsh���ƃ$�O�wr��j*OH�����.b�f�=�B�)YA4,��mX1�$b9���㨔י����7Qd�A�ô���i�EȨ�Ik�m�v�wC��r����̈́���V![���/VINf"0�!ݨkS��V����z��r�Z�������ь���"
A֤n3e̫YN)&��9p0�%
.�f�a��Y�IF��-�e^˛Q�a�ًvU<�"�	=ݑ�,��EI��[N2l+1����]�[�[���x�[u�d]�4B�2�Ix0,�Z,�)[�E�ܬ�ךV�o�:5�V�ʛY�,ҧ�x���2�MeAwH��5(�Oj+YMhV� ;�Jg�7o!��[7�p�Q)�i3k�#^�����+7��X��
�%�`O/qY[xM�`b'�P�wM�'��ӽb��:����J�N�H�$ ���{eD�6#�r��淗x��o(�b��Y�Be*�3zlL�̫Eг�'2QM[��Z���25ݤ-l����v1�[Ha�R6�
��Qi�fU5���Q�w���En�*��Y����Ԭ]M� ?l4S�V���W�o��'2�u��elL^�X�ME�i^�s*%�oV2�����aRH�.��+�������ء��wа�S���7l�dˀ�Q$뭧�E÷q�r���c�U6Am���^J��EJ-�UQ�Y��U����=R:U�4��޴ދ��Yy[�Y2�!��Tcf͓�͑�������Ytuw��H��r�^�)�34+so�n`%TEI�k)��)nk5����պ�p�& `ƣ�ڤ)2h�5��+ĝ�X�,�ó��P]�rЂFG)���nl�W��-Wcj� �!�/50˩D�ɖ��m���ಳq=ǔuDmKݛ[t6�ǔ�ųs5�j�61LŐ(rR�ZF�԰6�hlS�,I�e��&���(/iQ`���l<�����]�[yEm*2e�[ج]&�w++e��mӉR���A\�٬
b�JN��x_Υ[�Fh�[��XѮٺ��{�ּ�>1$x��B
�����ޓ�+bؗM
��;���y�F����.@�C\FX�@�fMr��T�;6kٖ@� bI4���đI$�I$�I$�I$�I$�P�4A�Zh�ٔN#�&�Owoe*4r���I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I%�jI$�i$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�C�\p]  �x���6Ɏ����
$�{�[kGG�0v�y��k��WuR�-c�c��n��f��'Cx�2�;��PH�V�WH�"�C|U����@Efph\-V��V=nu��m˲z�UID�V���S��Σ
�
��ͫ�~��n����|7�a�ީԚc �n^e��/�2����m�AIv�72鼴�
M���۲FG[�.�#^[�grj��&�4X�'f�#�/����f,ݼ�w�+� f�H��h���W�AQ]p�����n92�T����ղf��2��ұ��j,�`��Ύ��<���y������73nm�2��6(X��\j���ݿ�8%�M�r�.Jx.s7O���k�!��/M۩k(�!�v(�x0d�!c'B�`�{Nq��#�~��6��d��x$���3 �W�_ȗ�7��X� RNeƞ	�W^b��wP)�aʊ�s���� -U�����+�պ�$+�y���Cx��k�9��b�|м�NZ�B����{���+Y��kxr��P�5�`����`v��/�o�ID�����o0���8M�j�������ƫ{y��beF�z�u�U뙵�Q�r��2��(�Z
�;i�LrQ�	��V�M���u*����JSA�{%-5�]��7�ܺȸ��P�;sS2��#�ӭ{:��n��Y}�*�}�q�҆��{E���C��|��:`��I�����'@�9�rg[u�(�۝V����)\jnL*��9by0��&w1��m�vV�u��9GA[�Ḥ�b<��7�����
ᇡ3so$�o���epS)��*��.��4�DT����N�h6���y���Kȥ��$��f�ڴ�����d���Fܷ�e�)mt��A}���,w���J5��UmT����:�p)��[��M���mg^��݌z������p-�E>��l�ͻ�[A�r
��W�t<v��t�M6n�]�V���+�p�+�[�o;G<T!�h�6!��Sڵ��\�!}KcG��S7��\Y��fr�Հ�����W{�M	LJ�-���:�L.޺��YYVe�s�|#���qh�[�@��[N�sgU�diY�9%jv�c����'.h��~�ˣ&��S4�Y��J�v�pe��On��T�nfQ9�d�W�I�>��<P=�̺!��c���n]e>޳\�"ܮ`.��P�>f�އ�Q����w;ֹ͝}w�C�]��L �2�n͡x�క��m����|]d���e�pf��6tn�/��-�:�;��(��Y��и�T$ohܯo��9jnf΍_V��H���l舌��ӱ���1v�/&�C�K�f�ÂX�:��zE�*��ĩQ�"�XqS7�t��*q��ɥ�;ٖ�[�Exi�����������'�k�^�l�{p��ɥ:K����=������j5�3z�`�|MfNLVs7��h9�G��ý����U/�Ë����c���qK�� :�6š:���yں��.ߦ�&Oa��7�sCz_.�}]e�g���m��ZPM�W\r3Pc>��;S�vxv��AkMI�}:�����T좡Gd��+N�2Z�F��9ү��eɠy�h�7Y�㙕��X_+��&��|�y��Κ^`��ᙃ��%�$Ե��|��ɳo]�we�?C���qӦ�hL�K\mR�ñn\�4�CM־�y��8�e-.c���y��@�Q$TI�S�9��&��'{(P�2 �N*��k�3��畖�X�Afi��X5Z}���.���d4���9j
�f㻻�%�ݠ��zouH��v�����ڡ���ɷ��v>]0͜u����B�d�h(�3�ƽ���2T���yA<���B�]�@��A�V�m�r��n�q\�[M=���{������@'�>@9�h[�?;�X�Wy���TS"ڰ�[��;�q���q�����^���;;Cw�}�s�f�M��������O��F�q��c}�e̜�# ǐ��|/پ���UU�7����K�Xц'�z K���Mew^�2�&���V�E�&:��>κ���k-#�>˲ݰ��U���&��}%��ά����ǬQ��#�.�����d��,�F�]�Xr�4���ȁ��,�������S�d6���O�A��;�aKԴv�gSG����2�:{���I�xj�4�B�b�j�*6��q��o�s.-9��J���}��i&��h]�I%h��ŗ����Wl��nM<�W���S�v���ǐ��V��uzΞ�f�;�ɖ;T�)|��:U]쭹�
=+R<�q.��\��:j�;f;/Y�qhU��;Y�3�B��hZ�-�^�s��tM�-����.�s]JӼ�c�ٛ�5����ܜ��W�Z��<P���vح7nc{ؤ��*T;��T�w:@Nf��\����>9�����=�V1��8��ƍ���E7�s��V�ddû-�e�-���p��S��� nI;��ɆlW�c��Ť���'�vʲ#�Fۧ��c����cu-�����ze�jh�Z.�x-MB%od����t���"�\f��S7V�Ÿ�qu��Wr��;_V(��Pe\��v�,���t1�q�9�΍e��E�R5S�]A����,��KuP����֩���|9u���F�(j�Re�A0�-��Ҽ�ە��\����2V��,�rh���˅�wL�3��e��Yt�ӝ����h�8u=�W6�njX�35=,>˵.��d"F2Tn��EY����YQ�L)�~T\F-�����s@�M��t=��;��oi�?�d�{����&���(�IAW[�iĂ�S��9#kQ2���߃�`��q颊�S.R�p[�LØ�ݖ-��y��IU�C�U��˖������OS�TM���e�u3;���em�x�iC�v^#ǅ�Uf�;����6�R��H���׷�;�D�ą��t�+��B��a�}�c�	�8�� �.^�}սkY`��|���OLލ��M职yy���MJ�e�-��+PЗX:�Gn�̘�u���5z�7z���8^�*mJ�W/n��	w�I�\&:�����n�4X��wm���H!�g�S0��wu�bLV+��`�L��-�fUK2�NW��3c`�E:U�Ct��'E�p�yt�m@�b�L�H�=G�{m� ��9�/��v�bm+gv��E�����rj����u�J�t
���K�Ά'u�՚��<��9��vu�a�7�Юs���%rc(�����ڳ�.QՉ8֕t��NM��/���4ަ4�M��歍�G�Xv�I��H��mɟ	�v aTp�E`W���nq���sj�&���%j�h9�+#���D�s�Ҧq5�Z�52�!��7��d\'v��v�(�jP2���:��J&V�
��Ǐ�^��z4Z��S`��c�XW����/�*�Ǘ[A/w��I�����F�7�Լ}D��N�5|�bx���.mM�}`����ت0�qu�ILpDV�>��ы]���V��V(u��l	S.�ٽ������c�p%u�@�E7�(�tY�7��]�C;x=�{���`f�1�щ�+oz�\/��Χj`�VSWas�8�W��m��_f�{��Y'<�s ��$��-����X��7�{��ְi�i�LMY{�/�C�)��l�J�d�-��J��('��ۮ׍������:�MIѬ�\�$��$� ` �$���L �$���$���PH'k�I��D՝aN��9A  "I)($�y�W������A�i��}�[�¸5����*�0M=}��1$B`�/'h�.��
��{k���s���خ��H��<��knw�Yӟ8��8ڛ��m�]G���Bq��t�)�;�6
[y��QX�I$�I$�I$�I%�v�ݧL1#^�9���(������6@5_* �X������Nf3Y��$_n�2bVq���Ͷ�8`d����l�"�}PQ���	bT)��eQ8�#E��'M��dJ���]�y٫�l�o�p�8��Ӿ�S ��z���x9��tW&`5�S��et�F�3�Qh���Vk@q��ŉ*��rV��9�D��WO^^*�/K�f��&����T�·���P�5�y��8`/]7A���7��@Z�������w��PZ&�ǱF�=;dwX�i��q��P��C/�s�:����Y�,e���q=��$r�sy��7E�{L�;66�	3�Q��a���ڤ�Uۑ\A�m�v���l�:X;��P��377���ˎQ�.n��0Y�A��*����:�sRՔU����2���l	�lw���2m��z"��]d8�;"�:�0��t���\�C� ���Ȋǥ݌�̹��.BE8F	��؜*�:�{�j�<4h�6Jt�NRA|�fuF���ۛ����׆��|�i�qp�0��6�U
4�xpSW�*3!ۍl�2�ՙ��)��wNf>��I��ֻ)0L�*��,��M�=�Gv�B^�pG��F�Z�QL�y&�^�ϲ�i����Wv���!��g�7׺��|��ݪ�[��,�Vx�p�m*/�h&��0�yf^�K8"�C(��4������V9���`�����$�5'n��g��q�W�}�ܓ�P�����$�ͬ���(%l���-�
d���y[2�tg���i���#f����/�6�4��S�/� %`	rN�	�fӨ�+!๲�HM]�5ڝ׋*��	�1�ӡ7���VvK�U³�i�V任�zJՁ�&��LFn�9�z�
^]�����{�<�^8��ds�%j=�K��������V���doo����9ܬC�Ho �I��sl�Pԥ] 5��I�5���[A�,��<��;2��Z�L�:�ř[8�ɫj��t�OC0���b�n��/P�ʳYd�/p��k6�i��V�J�6�n�����	QZ�K�6�d�K�N�j ^��'}o7U}TE��9�n��:�E��M��,t��foE�_^��b��;2*�A��&쁕�k��f�E�#�eZ�wl+���[���Ҫ���Gq�v-��.mJ��"<��n�S�/�:� WC�u0���v@����8�m��=�k�-�0�ŭ�یI�ȼ��YJ
g�)�*�ua�Z���ɣD�C\����Ԑ�Nawڥ��gb;���5s ǂ�&�wK �(�Fg*��q+j9�������R�'Lň��ZJ*��е�r�y���,��v6���}C ����a'����R���(�l�[��3���B��.R���SlX����t
�.:�q�Zh�[q�t�D��8�i}E}�:EuΛc�\,K��S���ʱ��8�Χ�b�r6lvdk����fr�d��TZ8��&X�w���꙱W��{�g|Aa�:{K�|c�@C����{/���0z�d��+GmKh�֛Ӧ�[��u��*p�y�W]�GΑI����-�*����Z�1�g��ٕ��҆v�����X�z��Y� .�H��3
QG���bv�έ6C�^�^�W0YR�����ݸ�S[֔�*�t�����HdЫmHI���I��j,]Zݣz%*��69u�7�9@:͖/��W\�t���c0ʶ-�}VHٸ�80��
ze^�,��Rw ��S��`�	ŭ7�Ն�O]��zt�i�/�^�h��@ʻ��ov�B���^J0��$�� �fh�ˣP�����ԫ�����ֲ�:U��6W[�M�}��Z�֜�r+?S��#�p�e�Ƙ̎�<,�Tx����x�YKd��̕s��ݨ-��r����u�8����VWE��@��F�m<Y��<�1Ѿ�����r䅣$kf�񉥽Wyx�_وɖ�WMM���ѭ����YZF����C^�+2Xh�K�G�H�8��L��\K{�
�'��T_^p��;4���s�:���}�\_6AL
;or��z�������|T��oG
�|����gWF�.�9����vQ����q������ǂ�hbb�����)�qj�G�s�wI_H--9����%p$��P����Ʋ�+�1�fM7�h�sVT풣�"` �5o+�b�u���k*|u͕��".��d`u:B���Oe���%�S�s �t��֑|.&5v��犚Ю���m��VHj�Ǥ�;%uK6�#��N���w��A�kc��R�c�bK��Qu����BP7c�-�쵁d_vEv��=�"��_X5���_ �ƪ�S�d�v���D(�l�����^R̴�p��!��	�.��I����d�wa�Ť�[�D�����c��F+̏-5�+���@��3�r�Z!I����=���>CK����4������I�3L(�Hѷ�4�S'wN�q�j�϶�ȩ�[�N����L�ǁD���|�ݻ�,WrW�Fn�r��u�k��e ���H��+o=Ƌ��S��r|DmQi�f��1�B�'�͕�z.��y7�{�n5�	$�k���g0\�W:�J��b�w�t(�Vz���7wl�M��U��RNOqe�}!�&��ˬws��Nxz�*d�Fѳ֢tUɥl²˕n�e垹�5o��pɘ6]��ݦ퓍=�kHP���m�[W5��5�i`؞�)�lvQf�7�yRj�l�=���wFP���\�]�;أmR��zk)O�*�����*���o�Jl�?gL.��N��{�[��s֍�ݙ1��_=U�WCP�͒>�헝Ug��J4��9k���;J���:d��&]�2��wfjN!�����wo�Lu4�q/%թ��n����
/;��.Z.N���������T�>3MK�0��gkщt*B���y�n�KLs �8z�\F�M}Os�7����k�ŧb��Z�W���3�q*tozE�����du�]�����;%��CF��m0G��Ռbr��	t3�����gw��Edfnŷ+i��#M�Vu歭5��<è��*�Xd!*��*K��h�C2t�8GZ��m��e>��Պ��Z`�2I�J���*j�X�wZ�,���|r�E����ˑ(p�����]ҮLq��oo/%������c'V��x�Z��S���ks�vc��cx���<���>�����of�ׄ5/����mPB�q�gR�ɚ�����)[̾C1��z�J�Ɂ��Vk�͏��h��N�u�������]H��&�P���Y�ukz��ӳvd��+r�pWwc!w���3���VY��|��k\(�T�ڭ�q&.颦AvY�� ��,�Os���x\�0�	�c ?
���#�I2�#bpc9�j�r"0^^$hFs1�U��<9�T���V��{y�b]_bT�*�.����/�Nn�\�=8k��4�MPS��XX�L��ê���n�fc���=Z8��+J����=���W��u�pG�w�UXzf����z{��:��λ��W�}�1Ѡ���t:�6.�$��z1����v˽&3y������Y(v�%5ź��Lbd6�V�-,a%�u�Y��}�a�"�I?�O����MVJH�I��n7]����u����]H��ܩƪ�� kSGJh�TU��G�`v��<-ͻ�.�R%�˘m������6��Ml�K+F{����WK3��	�Y����/�NO~�6�M),��C&����9������.���(�QDL]*�푚�{Gu���d
�%�2��H'���K�e\F��S�x�p�I��V�*7E��L�K^8�k:ҏ�(8��͍�<�{&Ѥ�{kyU�}֤�E\&�}���/~ׯb�aE��;vi���w�͜ܔ�wlJ��<���X	�E�f`W�c��I��f����&=��M<�iH�q;��:ᬷ���w�]�0u���?bI$ ��)��? �N�$��dbcqv��ߨ\M�I$�I$�I%w�YV6�t1Y�*�ĭ�y�q�H�+&��
��n�&S��%W]u���P^aPX���b��i��}�/!('J�!��7�6)Vm��s�J��mC����*6$�yy[���7�N�;ƹ����_3D�����Vjbg� ��k8��=�]^��M+�� �\F�q�}7;�ޑf3*l<F�b}�M�8�D����׳[M��t��N_�	C�9���a|��������˽OE'F�bX�Ls+5�;�bK4���i�!��A0SP���i����-�<�Ȫ;�]�uc:�oWo ƾ��L%tH�����3�Y���[c�����e�*`u�56��E����۸.��H�C���eaH`ތz��L�s���fb�`�(1�b��7v�,�jV&�4J#Z�`���i1]PNq� � a�[��ל�]�*��,���Ư�齈b<���P�ԒB�bNj;���J@�9�τ������TN�`a�
�H���e ��Ad�ł��&Ӊ<�IVP�JM$YHN�)dRM�ZL�+ �R��IL)�)*�
Q"�b�T)8��%����4�0R껇R�E��)��̔Ȍ����\T`��)���US�DQ.��L!I!!�[��?�� O!�.ߥ
�k��������Ew��Q"e�س���U����)t����U���^cw$;F�X�pQ�2��{R��7�Į��kgb{%��8����F�[�N\[�.�`�} �\'�+����{-��:���xVd��K�'6���0��н3z�
0�Pf�;�������$�$C|�!�5W�݊ESrk�7�IS$����P��"ND����߬W��~�My��ί
^������5��r���׺�j�D:��J;��'��	q<F0m�fP�1:*:��6�}��៣�_���P_��J�-�{�D�
���I�R�nۋ^7�F�d�� ���TtgI�yh邷�"�b�o�˛�I2w�V�ts*]����b�{���s4c�?v��ap�[�^ݧ�' ����Inљ��V�=<3j�)�a��}o����Y���G;cY=��j�.��Iv]�9m��;�[V����<�P7�DGuڔ8ܲ����NpG��j���;W�Bs�.{�v3z��+���<�}�IP���ʴs\��5'od(�G{[UځW`�w��:�s*Ĺfʜ%�ۭx&�v*T*1y�6�έN��Ngoh/�-2�ɖ�c;��%�񍼴Ϭ���}|��2��ט��tP�V�>z���j��߬4��R�zl��#�y5=�e��uQ��7M�1��=M�F[T�U���S��w���|ϔ����k�;���)c�r�����u�|Qy�����Cu!�-fl���do[�=�^��
Z���^p�>��g�ѕ�������%��nkm��{���ͫ�B��3�kWr�5uw3��
dv�
a׻0(�Ekk^
̾m���86ZԵ	��xr��h<�}<u��du�K�v��$NF��w�M7"��aZ��0����Won�w?T�Ǉ��By�4*�_�EF"�@\mu��q~�嬽�����쪬՗8�<P��I��+X#��v����j�RȬ[�qg��4�y��H��s��M�%�	#�M[Zrh�̘�f��Ȼ�F����;Q�/r�Gg���
��F�{7ル;8�	2�s�c��dnԞ!���n܂|@qD�4n�[C^��#�q���.���G�^�ϯ���T[~����6�i̼�fE��~5�z���Mg����$�����HVn���B{J�KuqŔ�#��,[��h��}P.��S0v8�b�p'a}�.�Ć��Y�^w8;�k�Ź�[ѨlW��H� ������b�5f��n��6��&�a.�.9��ю-q�oh(��u�E�@��ﶽ�7{	9]D�6sښ5��}�U��0��Q�������T���Ƈ<��k�3���z�m�:>�T�o���F�egEΠ���!��Z)E���DV�޾*@Ot��Eݑٽ�W��(�&~���v���4�O2���ψ�|�\�vgd��]R�6��4����7�v�".
��y�ͼ�.�w�ױ+�Nd�Yq�|t����]�P�._�*��it=ң�b�6���)@��MY`����U��'�Qw���0��:�ʖ�_v�dDZ��u�e���	��;N��[�wR;䗯�v[L�2����D���[Ywd�7{��s����Nv�X�Ƿ��3װxxn����x��bU8��e�w	��w->Ѫ��V��ҺgEȑ��;�������+�IJ-��a�i4���^S�
�Y�p9�8�ڞ�y�8��?ϭ��~��v>"gZH��Fj�oG{'ڲ��֡�_+�W#L�>`f�H�[#N���Ud�.����\j�n0^��F]���.8��Pc@�U�],�ढ��Ej�\����vz�v�͑C(6��ɪ}'��Oe��I�5
�#��经�S�rmV��s���*K3���&�n%�}��ְM���q�yr�=�)�e�F	opa�V�ʬ�J�μ�P!Ld�彩c0��cTg`Z�"��[_cu�U��o��2����P̮T��dWV��C64x�ҝ#�����[�;Zw��������#��`z))�{YՎ���ن��z{3�X{���3������Jy�]�;��"8i橭��ěT�'�Uڞ��d�X�"���ќ�8����R:�Y2
N��.����N(H�vf�J����^W��>=2�S��	KeH�^�Vz�7}�����C��^�L �ka����WչG^R�b�.�hE$���A �I<��2yTB����g2��űP�>�Ѣ�m�q;	m�k������n]���z+�߷)"O;8���/��=c�e�.��ۯ
�S�&\5k��fAӅ޿�,�RÙ�_#\���X��|��k+�n�]>Q}K"����.qyʏX�`��|W��r�қ)�'�X>�uf�Άz���6Nck�4���gv��]v��쎒GG��*#��֢�W�Ӹ��Ѣ��;�Z�J�=�B�U��	�m���Ws�s���Usd���Q-�8b�#�y�Ψ��J%�+\��:�5׻]��Ka)vb���|�F��x��E�����߽~����w�_ѕ�o�V���3��`��]��N�F(;2�b�;E�1�U��+�,��;�a'�g�����:2�����g��]:��֝�{ϵ��f��S�=A��p�u�� ��yT�x��::>��p�W��#%��@��P�K;�����Uɻh ���,�c:��Nh���\H��4E-Ş�o�8�ն��#wswC'�]�`����ʸ尣��l��'������R�mAi
���F٨]ڶS�O��Z�B�gv9b��W5Ѩ�����/X	R҃���r�A3�+V���V�j�Zpm�L����4����Wp��k&Ѧ<��sˈ^=��ovs�k��{���h׬1 ��)幛����e! �;s�^T4ں�4�>�$�h�w���׀P��M>�8@�:z t�Yn�Y}���вEkl_o,�徂�'9�_��Xt;��{R�.Omsz7�����t+��9�3[��μ��qH���X ̤-�b���z�Tu3�:���G"��a����C�n����1�Ps(�Ů�7����J�^ԡ1��Ƕ�2blsÔN�=�"�h�����@"�5nm���Ud�¦��	VUI��V��H�V�Fǩ�z��-WWڪ% y����F�I�9O����b��ZE���d�Z1�5K���1�b���=�W�O���0��y�3�� t�<��p���lw����[p?S{<�<V���l�X���l���ݓ�gj��f��[�i;�ӹ���n��s>ޢ���{9d�])�4Y����>Y��\��"C7L�R�(����ty�`C��<�|]u�C�]Q��\��|Q��I�J����W�+]�û���T��"6ء ��*��SZ[�Wf���r����4�z�f�#�,X��x[�]��0��D�W4�mح�,eY��C/t�Ѣ$������*'w�� �Έ�E�I;ow��k~���������:�>�;4ǳ�.�[�)a�ˋ\��K�:�F��--�9N��H0���'s)�vp7ت��d|���:Ϩ�o�uV��VM�Z)M�2{�f$:J���*��
7���,�=�qoJ����K�~��.�33���`��+�K��ٽ���P����\M%�$�I$�I]��Qy�/Q
�_ʄ7���긅��SJ��`�]�*�0P�T�jP�>81٤��-'PU����.��0D��'b���M1����cp@E���T�j��N:I+ʍ��@��d0��R�Yt�2e��8~��d�*H�r՚��1Hi��b�8,q۔՘F���C�[9R��Pd2AM�2�زY�K5m���k"聕yL�$�Ѧ�$�d.�~Q�ZW����mRY�̕H�%%�u�8B�����e""h�C$Th�o�.�j�����̱��K�*��E��6n�z�W�U$�u*�lU���f`)��Q�wS ʻ�]��%�YqB�X�	��W��;��yM�N⧌�5f�f�`6��^���ݑ���H��sZ�>?9_��
O2�# �YI
b�!L-��,�Q@�a*�DV+ul���SL
d����`,�ЬeT�'��"1��Jb�T�Q�����M4�&��a�0,L2�w�L� Y�T��!Icl�^��P�Vd���-:���.*�AUH(�@�E�YV�Ƞ�����
At�HK�G��t/YLP��EduE%���Pa-��HT)��h��Æ���Ȫc
a���+x9g}[���6�c�7&�bѱ���x<�����C�֑z�Q<]b���
\�aa,S�}�M�jI�tf(K� ᢓ|w�whԄ�Ll`���G����}���V�me}U
�iTg�w�J_w^B��|ހ	������/G�_��gwo�)��(+��FQ�~h�?k�w�f�nc���#����W�����^���
R&w^��3�%l�т�E�����R���`5�}Ž����=5V�h�������p��f��B�����*�n�'"�_���L��_lgHy�>��i�I����y�wBW��6���'X�2
��TS�m)�V̓�	d/���;��U�}�����i������G�`p�w�#3h	' �}���^AH�52;y���Z8~�y���C�O[�N�P��0ѭ��ዔ�
~����=����I���h?���4�O�˯o���ӗ��I��m�XlRX/�ߖ�_ue�2:��E/�Tx���D��G��\I�U=�$�O�U�i�k�u�>�Z���4�j��������- -[�Oop�FWО�}�c���1�2�j/�����p8�n��k��L+��	�U�W��AU�Y���f��k@%���������uW�G�U�N�F4S�m��������F��e~����pL_n��H��! ٬C�.�V�om��w/��Y�1qR7d�F~�!-}�C0�����t��vU�ݩ�3WIc��Gh�/<��y��,��g=Ƶ�y���������w˄�y��
t�ŉlXӇA7��m�U�ѫ�]�s��o����ݑ���#열�w�U���*�%���}p	����\.p̭D�룕q�X�DԴ�'M�If9�
�J R;j�Ű�݂(�_�Á��˸��`�$Y4��݋����O��9 �nx��b�8��n)��hv�o�_75�]8h#��,GDs�܈���@Bj�B�ll<e՘ω�ẝd�a������������&�!2��6ɔ��ԆR���0�`I0��q$�L��Hm����� �|>�����Z����F���$����5��t��4�K^�u{}��X��Gq\��ೱ�	G-$���ɇؼ�t���C�H$�vz���X��Ū���������|�=��'��u:�;���:�vR���2�N�0�y�Hd�I�M⤅�RK)����������o�G�~ i�I�8�<�f�N$�CL��&�u}D� �ScU<�Ha28s���I-7�$/��:��h8���ΪY���q |�|�q�p�fRd�W��hG~���n���u���@��UI
+w2N%2i����I�g���C� c�&����c;{y��o�v�q���� m�d��a��Q'�\8�@)'�a�`n�u |�d��A䐦">��{� ���c�$��\�EϹ	ĝa˨l�	﫨Bd��]ܐ�T�d6�Q:����@a�7�z��݁�@R�>I���(����8�T��I6�q!��7���!��XS6�W�����V��u����l�G�M0��uu�!��d6z�:���-s�a�I�T2i��6�3>�iOV�߷���^�M$6�#(ZB�!�Q<�:��2�a�� d�h��m�Sl'��V�T}\+;�����C.1P�@Ǩ�Ϫa$<�:�K@�Q"�ɶHc�YB�Q@�!}�l3��y�:���6^]��¡��'[;��UwZnܷ[��r����+=b�rts��i!��\�ғ�Q��1�u���u��8V���Be!! s9���{?m$7ʁ�'���4Ƀ@�����*�1�@a'�<�u8%2��y d��������������=!ԝa�)!|��J`_��f�I�L���I�����D���L�<�p��0��d�^9���*����s����a��e��N�Ϩ��3�\�!L;P6��-���u��06�d�6O �g��|�1��������)�PC��HB��m���!��!�4�0���&�&=RB�T6�����d�I��������{�v�I2u"��&P:���Hm��q�2��u�l�]�<�Y��8�g�H|����c�:��^����2�L���c�H�M�<�Q���N���8����d����8�c�@����I�V��W�}��9�hC��&�a�L�]I4�f>��(>@�!�8��'ɖ�mˤ�l�2Hq��5o�]��߹�ma�He8��!�q&�O�8��K��!ev�&�rm�S���e�L�a7�{]ůy�~�x淭���2�3��Hy!���0�'���qy!�E&P8��K5P�`c�N��l�`cX��{��u�����0��f��(��z��C��R'*C��Ch:��@RN�@�	-&]ʨM�?o�׵�~�?ͥ������íN����y�wNh�q�삏��͎K7.�BYN��u�ͭ��F�Op��u3]z�7{�si����0�X�u����`/��u����I'�'�8��PC�C�'��0�)�Ru��o��P�@����I�T��k���V{���&Y0��$;XS2�q!>d4��4�2�C�ꇘ`q��y	I�u�z�#�H:�5��o`"xۊ�G�_�9�Si3� ��1�	�C�O�%��
0,����r��II�����-��o�p�P-���$XI�I�T2i��y!�-��>Đ�L0�!ęa)��H��7�'X�����W��~���S"�{T
� d�ԓ�E�I�'Y!�,�
��C�M�Z�ԙI��}�c���9�����C���"�|��$��`q���!�Ri�d<�2��T�$���5�e��u����v�Z�:�u��ɔ�`_*hL�Z@�Pu�/�a��N��@�y�8����&�M^�v��hCu@m$�դ�@0�$��:�Ha��I��T��q'2�u��a��\��������s��y���'ڨ�ct�MNԝdX��4��	<�C�&�|�`y	�ԇP�6��d�kV�y���o�C�{p�Hi��Hm&7�<�����3rq�`e$�������H������n�ݷ����M�x�\ ��YpT�N.�)��Za�;�ryUUу$(���432��ص�r�:M���'wk��9�m�u�7ݺ�?!$$RHI��Z�{��v�\޿!�8̲��d0��\:�8��B�ʁ�$��e�u��i�E �Q:�^*`i��۾r��kw�>g3�O�y	�CZ�M!����gjZЛgRm$������h�q���+�߷�k~���4�iv�:���C���V�!�:�䇞n���R�~�Πq�6Ȳi�I��=��O~�9O���u�}����JI:��M�>5S��i�M}RB���$�aL��('P�&5A�@�u^�9�5���}�v�a���'��K����:�h�I�f��HM��$�(-�2]Hu�����:����ﾖ^5����zi5ʀ��b�e$�N00�H�������C�N�&P�R'�)�k�}Mv���;�z�l���V�I�L}G�٨I��a��PN$1�
g���	��y�ޱ��//9��uｭo���!j�HH}7RdXY�!����!_Q��I:����d��y��g5RB�(�2aX}�������c;��w�0>Ǭ�I�b$� �T��P,�dXY����12O2]Q�M2Cl�0��q x�{�s�޺�Z�w���4�}�2�f�6���H��4n���C��!�C�L��,�e󽿻�{�����۽p�n����^@8s#f���?��o��Ό����X�F�j��T$����2�����:��yv�̽�SM���{���1N���=��	$<�I���9��vu~9�Dd?y�r��x/Q}Ȋdu�z����#�"�ھ�G$jk���Y��͗{g�Jb����U����.��Q��ӌ߾5�6���4�]z"��MkA�Zo�qv��U��y
�]*�Q�Ԡڠ�-��(�Q�$xh��OOlw�����夷������x[f�n�'��������Q"��WU�ȮW�Y��$���d�zR�w1 \hr�v(���eb����P�N�z؂t��z�9�}}�^H.�v&�f�qṢ�Jq%"MK-��v��V�6�*�{3_4�����d1��߼�P��x��s�]�`��/�o�^oڽ�8�￁l �( ��ﾤ����1�g�`U�~(4��{O[l%��e1OO19�7�p@=����ȡ���R;s�D��\��@�MfE�����з6�X4Ѝ�9��KҝN�h���L�/{j��,ѣͱ��ѱib�U�ÞWo �޼���3kЭ��:5��h�eI�7ܽ�����}��+l����=�v�Z��bM��P@���ˊ´c����o�yۼ���{��X�V<<�x���R�&��k}O�v�c��9b:�����#�>O{��e�öo]�YMv�^�i�${)��"g�S�Ӑ���neV��ݕ��U�y�M�h���7s����d��D�b�b*�u����RD��37���}/}��$�ABHH�$ 
@�E  
Xd�`,�


(*(,���|�u˶�v�*Z9 ;���	�{i�&�p*Q����Q$.,G=��f��j�|>��M��0�+X�~��}�%�6@浮}˪�ru#8kGT�p���]=��n{i�{N�*M!�mi�=nb:���N���Y��K��J�� ,|��P�3דz1\ �j0�*n��5$��y�LhY�.�9�b4C�X����S	4�z�Cx�b�2���L5���=��@���)$+5�B%(��D����~��\�wǅ}��4b�ϊ�]�:
g�a��KG	�.��I��u��G��n}.�oA�,�{��w�Ɖ�p��f��X��y�KS��S�6�UCԷȝʹ�0����ʬ�7]���f���քiU�T�c�!Z� d���}���":ػ�ƣ��0sE`�0m��9{��s�ԸVn�jp0P�������Ŷ����e���S��Ӕu��]�n��W3&]��6�i��(݌�؊�Gv7,N���g��G ����Ʌݔ��.�7��Xm�[�&ȸ�yh����/reChd�����f�Q���ո���K4�I���<q�[أ�nA������N�ָ���쓸[8@��P�V�좈�ڈ�7��1G0U�'n��n�u���M����Ջ4%	$ᙹ/���!��i�gp��I{C�7@���Ԑܳ#�Pg|�1��3����2��͟�����I$�I$��.�̑�1u9C2U��5�Z���#�w>��R�A���["Ҥo�j}�H�:0@��y��ݖ,,6����h�:�56t�TM����p`� �oZ�/��g�cddv�(� ��S�Ŭ�@(1��C����PB^U
����C��i�I#�ZtU��	&���4�zA!��T�sx��5x[�Kk)*!n�4��32n������E ���$ه,^9J��Ta�^\B�
�b�d��%^WQ	]��a�`�c��%�Yv�4�b��1*��]�v�(0��ëq���ſ]����ϛe$�n�(�[&�0n$,�5�c�l;z��m<M�kO��Hux�.��ՙT0)aa	�V �{��"����[I�h:�G�]�����:��R�?*�&��U�?�B��D�wU�5@S%9�[l���hPqQ#�+�Ra&�J`�Im"��uwFh0��qB��RZa-�)��u"��a��f��-���b�ԙو�SIhf躪p�6b���i��T��.�B�x����lah��j�K�b�W�c[�3�e��L��T&Y����aL�o4Z^�*J(}����,C�S�\��ٙ�f�fM�淥�D	����s�A���n��G���z=�ĳx�S�1��ք�?ŏ�SN|�͛w{y%tMN��:�{q���c ],v,h���+j5m�p�f��S
7�]�lㄪ��q��t%p�N�0>i�zS�
<)e�����a�V^7KHE�.vaF�o��T�S�]��݃���;7m�Ƿ�`c�,��U�8�L(�i�|��x�\��Y�^{�s�2bz��A��{��F*��>�8-���|�\�b�G���O�a��Y��֧Fk��tBiB�������eY�q��y]k��;���|�Kn�~���1)����z�n ;-mu,�jM��Ip!�-�u0�R�p�P�����z#v듢�T`bE�Õ�01�q�]vh�,l8Y��>�r���r��~]7������ٻ �}o���R\ � ���ys7`N�]�!H�ݹVȇ��łcA*������|���^�kq���;�]�qS�}Z�AG%ɉ"^����WP��ʋ�gwN��K�c����l[u��}q��
��:/Pmg`�G/Ϯ�c@���X�5@�݁y��)�A��j,��Z5�}�iʚ}�ݽ*��<��j�z�b��wd:�R��X`��ry���wM微�gw�^B��-B�s�ܱ������4�� 	�i�|̜+�9]p�Z��Ԛ�2w��M��G�=���η2�Dԛ�9oc�gcv��sn:�_F��U`�zĪ�䞪�YT�g��X����DEދ�ҫv��!�E$�lVI>��{*i�U�U���/�E������I��T��X��Hg�#�l�aI��kf����3:�Z��೷3Jcm�ͧ��ĥ��nU@��L���EU���ʮ ��r���?t���;飸U�b��b�t�0����ѓzQ�XK+�^�Tg<��f�̺U��#��Wھ�����ʌ�-�.AYXҾ����^�B���6�i�y!ȃ�5���tV�e\�il�:h�[�k��!�դ-��U�Y����DG�p�xh}��:W˧���SFT|b�kz�w7��^�w���x,�:v����@���F�ыxֺ�Z����`�;�O&����J�����鏓Xԥ���nԳ�Ӷ*���oI{�LI~O�#�\�88@f1�Gٙ"ޗSw�Iq�{��Z�A���_��ѕI��9]�c�5S��GDٚ�_ZY͹)hpV���uTQ',QL֬�Vw�sp;�Np�QǦnW)u�&~��p>��c��a}b�؎��/I��ӄ&kyuۯ�D�U�'��̫��i��b��s���8IH�!��u�7{�A�"y��y%����z��ܯ���O�I��c�.�9�ui��E�qy�!���"h�`�tG�����W�ZF9�p�琢��G���0kݰ��n$C�3K~�o"0Q5�w���z��A�"���n�^��-b�O
&��?>
���En��t��gXps3zF���� ���i�f3V���a���s�����{��66+��t0Y1#�+���f�����5hGx�_ec�R�\�aS��e9��Q993�Z�QflanIE�幬�9+�$Sv�+΅���Y�럕͸�>߀�ꯤ#��q��+��3	��M�	7����2xBf�ߞs�/{�\��Pw�Z�v����z(n��z��W����]L��p����A��X뀞=��}mZX�+{pw���n�SϨE|���[Ν,B�-,r�+
j�V<V�֧F��N��cx6E�e8ޕ��5B�9ýW�7�e�5J`�֭��J8�z`�+ț�w\��륕z�Wi	ֹId��; ��	ƪ�U1�+�/�w�Ȯї����H�Ѭ�y61�i�p$��Oz��r�J�Wjn,/{��a��kQ�+
�S���ׇ��w��]�F��O��CM�ga�ʱ����ݻ32��r�p�e�;V��t�h��2OP��Lo3�'l=��z�M��Ou+���z"=��4Hhi��	}��9i8o�����}xN^�㩇egA��c��f�8�8�kOU��o#3b�|��|CWY�;wD�ָ>�	T�k�Fi8��p�r՞�����{V�kE���w=�U��3~�iVx6Uѡ��T�\�[C��oW���gu7�sI��mObb��]$"�V}K8eޞ[�&Aux��5'�*�l�&���G|�.�Z]2�	������G-OA�A�i��;QO6Z�>/fDAd���0�<ffx��+n2��F�S}��e��f�"������`P���û���X [�a�<��Z�r��k��[��ݸ�ޓ*Q�Ee`<��|8\<��h��iAl7K�5oI�XL�Z�g !�ډ�\~�DG�J�A��������|2%[ Īu*�Y��2sl��3�q�ZC��d�!WF�`� ���[�v���ʶfT��6���r�a(�����y$1{��3%�
��x[��A�Z�]'�2�'x��
{5��s��n��J�f�����ƛf�I�{NgG^��� Yӫ
;:�X��ۥ}N���uW]k�j�K�@G��]�������Ӕ
�2���E����	���q~]�����(�=0.2�G���f�^�c�d�n_����Ԑ�w�Ĺ��vgv 5�0t����{����zT������,ﻡ�A�>��'�[���ڤ3��I�'1a*�@�8=:t�Ɇ�8z{�A��y$U�׺��BG��Xz�U���a�G�_[��V��\��켚�Ѫ��kT7�~�e9��K�,�[]���2U5�9��V�ǩH�w�0j�{�9{.SⰥS����&�M׼7��
AA�0�j��M�ݍ攉.9;�7�FK2���#q���k\Rbj�O����8ߌo��������څ���8���cZ�At����cL�XW�i;��y�D
�[Yp���NYo(��:�,Qs4�=U�Q�4oIv�{\�������NH�~���b�l�W/��G���� ��O����K�ƈ�'��ty}��۳�9kj������I��^ȗ1�2d�:�Al�ӫ�Q���bkq�=8`��2��Q�2{ݩ�5#S�.vPw���uN��4�ʎ�v'<�QB�f�ߵ|�3�QG���>��6��LΡ?.�񡉚#ځqs;��z���6I��ˮ�W�W��%������೚�7��A���dن�X\��x�j�7�����w$�90��[]WG��^#@{~߼V�W�Ԟ�_#���/��'��Ŵ-�:h���Mr�ݺ^�ήw���2o�j��>�9�ώ�&�ӥ��������T�g�x~ҙ�+o4�V=�bIY��w��YsPx���e��#��Q�.����R��'���c��w�K��+"�M�Fm�;'TGLްy��@`IRy����`�µ�E�ϝ'>=I�����
.e��vgVw<�s�-��Oa����f����*��՛]J%W���s�h�uҶ��g��^�U%{�f�#�j��"��@�S A޼��m9�n��!;���<���_v����͡�E���K�P�y���頊`��ev��*���6���*�٥��Å�.�/��:���Y��֓3���n��g"o�!]eav�.�z���`a��Wv�_u�*ҺԖ��q`"uqĊ�+PʎH;�'��$,H��Pm��톤Lu�{9�*k�R��v�pޞ�T4�\���E:6jł��gv��i�@ڷIb���u)h�:�n��{�Yu��W�w������O��V�� ǾT��=�Nb���I$�I$���vp��3;�bt��0k	˱y��2���Q�Z��.�ղ��$�]K#Y�)�VmJ�"d�WG*��5���x���wbЗm���7fP�S��q�YX�!F�[��[�mc �%c�X1<��U�R^VFw[ND�@��%�Zyp������7YF���+1�6S����1,ܽYt�,l���-<9tU&m��d9X�UN���-�i����$FL�AɦɁ-ҏ%AŖ�}f��M�n��f�����̓"�,�3ټD�˗�ޛ�f�6��E��:��cV��I������ޓ�����z��T�Ja[�i'1�4�E��K�F����ػ�F�Rѫ��^�M��,�l�m)*b˖��(S��U��m[@���QH��UV�V�Sl�Z-*#�8�L*����(e%]�m2e��tTq�Fa1CEU.҄�R�V*�.���@�*�B�nU\1Z��RS)R���Dk�]�c����r��.RV��_H.G�n���2�B�*Q9��'��Z?�G��P�7u���j�ԩ��+P������#��2qC�ϝ�uC_]Y�2�]rk'����&�*e���}�����d���2��ߏ�DkǍ�p�S��tkeN��,��3����Y���_����6��9w��䉘��z_&�Ԗ/�/�L�zz�����p���Liqa�eS���zX[�#��r�K�[,ҕ>�#6`M���ɽI�喔��3�D�P]>�@�7y�_�^�u�s�������M�yn��E�A�&� �v���p��o��1K	�����}� �mY��J�?1g�5��[��Ǥzi�J�s�k��z�NlTQ�t���-zt�^4~t�w�?%MKN��"LާE��OnfkX��`�f���cY�03�|%���/v3����x���M}�2]s��'*P�㏻�]`���-���;w�@�-w'��mM{W�/+:����w�����=��}�¨��Xsjԟ_��߮xm��~5���^u���/c�MRK��>�T:�]zie�ǻ�x��_Q�-6pG�7y;�QY���+���[�P%*F1`�N�:F����׷ڨ����Ƅ����ZFh����R�y�����>�����b�Q�C�~-Ɇ���:�}jNM)�2*j����7bY�AX4���n��B��̿.0�u�d�]Ijė�����b�*k$߹�r��eGc�1��r��uw2�W��+�U_��<\zs'K�h���0��颹4#���'GS�0�#��/���i���`F:�/�X{x�=�y�n�>A�a���l��t��!{�jy��,��}�Yh�ڪ΀%�KGL�NeJ�`�#�.�ŋp>���/g�g�}�����7���-��*ޙ\�����Cg�̓���$m��_��,ש��zq�ɐϢ�B��p�\�+��5nG^Ԡ�3�=,�uӛ��4ŸC��0��b�+��{Sv��K�/y�K:y�ͮ��I&�O�
��]�$~�tm߮��Ou沇Z�y�b��g����@�3S+,�/�*]+�{!h�]��Z��#Nz]W�+�hJ�n`��v&��#[	\N)M>�--�����f̓����:+(�v>,fH�4�9oaBp�/b��-
�ۺ����T^y�"��)6U6	���tx��x`;ɶǎ����"�u�>�ʗWA��;���39.)�1�Ic��H�oX�F��4�z��u�J;:	����r�Mt�rR�{A�]�X�ҹi:��� {��v�.��\�.�n&|ʏr��7I��/"��7�Q��k6�f�Ժ�T:�������D{���E݁���)��e�]k�]��B	��_l�)�_Q蜞X��f�gԨ�����`�t%�8�|7X�I~��q�َ�4,��P��-���B��5�����[���Qc�g.�&���p�_BVڙ���*yjz��\~�݌�QG�~zE{Y,U�/j�w�}����=����[Ӧv�x���[\���4YD�`q�{sS.�NeK�+�O@Wcz�TBzQ�?�Y���~ʙ*�������)���.�p��
=��+�]��P�>����n�DC�qm}���B���J�:Nv\͍n]�����4�@�Κf�$��!yq�o��~���-z�ڠ�,g���=�(j����Vˡ�Q�-=�7�)�y�oZ������7t�8h�&�܍T�̻�ں|fX�в�ͅb��n���*x%��J���8j�)sp��r�O���-C�}<U{��zX��L�՛����9�&�gL���<ni��~�R��w������<!�za�����|��
�",銁So���+8�5�ߘ&���qM��K�|v��/W-�w:�^{t�iQ�xW0�.;H�kᨑ��ʑ2jeȔ�r��hhm���]*~q3���=N�8�g��ρ�i�EC��'�� -�<-ɟ��S�=5"wv��:�;���e1�4�.#��Қp++ܙ�m&Q�|%������j�Ç�}��gSû�g׏�6W([�4�gj��G=٤��ő\��ƅ�џ{_�/��v�}i��$��(�R+�ԋ�[ʻ�2-��l$��e�i�/�w.�wp�P�@�U��F0��+[���-B�����-A)l���
�]��]1�`?\�jod�+Q9N=B[�wo%�Zx- X2�l�\o)e/^.��|�6���?�����+����F��yQ�9�T���U�����N��L6h�A>dޠ�տyj��o����*ˋi��H�ݍ�tEC7q~�6��4Sn��)y��Z���d�ԧG�E��*i�C�#"b�k�3B��MF��b��^��oiɜ�7�hG�L��ܴE���Vn�B꛷���7\���>��.�ie�{���]�I�{��z��G�sO�7�=uy�Gk���43�yHa�Z���ޞ;�n�荋N9Q<_��v���vR�
�5�Pf8�j:j�Eiۥg2�b*�5�MÄq�G�z�0�_���m���$J�bh!q���f�r��yq��T�\h����K��믃���CF�������D)9]���z�/ql���Dp&v�h�OX�����O�L�ֹ�s�8�R��l�I*=�}�����"�w�c���ܑ�u�4EeX�;:��3��wlq�R�y	�E�Ӿ��� �TE��>}3k/<�J�Ŗ-��u���A�9c՝�qyy�Əz��L}u�>�C.���<2��$Д��٬l��&L��y�h�55桚�９��E��N�CǠT��k�����/�dM��'a�9�;�n܄?4��.5Z�G���[���;kOR�;>�����6l8�K�3�����fT�
L�C֙{.����B�	~�RP)����N����#5J�Jx}|�FM��e�;R�t�;�<�"B���[����̃F�N�|�uj��y#c1^�l3y��,m �6��j�z��Lṩ`�s��2U��Uo�r4����㯂����#}<nR���+�,���P�+�+�^8��T1z�Iվ��-���ǽ���Ӧ�8���R�gM�/�U���W�w��G�a���=L?,#yf��������Kμ|x�r^f�q6�9q�񠹌:Mg�!�F��U�KL|��V1L���;���f�7�Lr��&\�H�V�M	X&N�OsI�{UH�"�|��EDd��g�\���x��Y�i��V�3}T�x���!eg;4г�b��*=�
�š�3��iW��,�yfe?|~�܈��1��4�z�b��]0�������ט�"V�S�M���ύ[�1��̆���B���)�}�{Wk��gk����/��!��,!}x��^��0�XOZ��[�l�kfǫNa��)�8޳��
U�{,,�����j��}��;����Gf۰j�r��T�3�.�OS��j�V����ׇW�f4���5Z�"L��.ЫPg탩i����妳�5�JH�Ҭ���~�F{�0� #Ŝ7���y�mq�����t�������`��ƾ������r�)R4\�qR���v�9�Vt�'>Z���R��\�TxM�jCl�ܬ���)�\i��m��eab[�<C�b�S��[F���^��-�x��r%�Ν~|w��ȟ��t�?��z���<板?Q��+���,41�g_k��Vؙ��+wU��z�邴�O�yr��y�P�X�,]i�5��G�jM���S�os:�PU��/��a�!Zǹ
��o�+.y��{�v��	�G���4�����ᔇ��'����'m�T�eߖ[���i�h�{p@�Je�кݤ��δ�h[U.3w�=^��o
�[��:]�R��Q�h���*V�C�:i�P��Y�"��L|)�
�IT@͵*}0k�n��u\���R枴yۻH �<���#�o5W!�k���)8+ �Opv�'�����yO6����t�-�+|�sX��l�M�ռ�xb%9�G�c�����x糥�<s�Ҡ�Dw(z�k�]��=/3��g�Cz�Эc �bva����_���5�J�&ks'�`���}(����"猛��kuGPf:AQ�=I���
�.��l�� ��&VUp��0K����{�G\�zG�㮝<�rF0�D�Z����$�o�[g{�m{�3��Jr"���I��n�ޘ���)�;�1�����V5���W}4���q�@<D��
p��#y��<��6��'h�c�����U�:��r����Y%���d[n9�@&U���g��}���6�
�>R�a=�� �IR�ⵔ4�4q�E�DE�/UrT�5��:�5FaV��iÕl�mZq��<�`��r�x��������q��G��¼�n�N��p+[��--m+�6~.�8��'fЂ��@��wj�K���2(0پ����7��y}d��أ��v��`��m�$}�+��X	������Ҍ���9č�#��Q���2���:��L�&����PbY�k��bP4r�ʳ}�(�\s8H{�i�,�x�n�嚊��.x`-ee�	E��p�]�c�g�����S���;�-&�V��̸�;�M�Q�"2ov�J���^�{wR=��}�)X�p�m�G[�P7�L2��mQa��iDQM�T�QZ2�K�n���T�C{�oe��ѳ,�X9%>�7i$�I$�I$��)	��nZ���б�� V����`�0to��y0����݁m�.W�':-K��B�uٜLuZ���o*f��u]��W����u�[��q6&��;�r,��`@�]���y�M̸ �ѺX8���o�gcCHy��.�|�(i��M�<��ͱ�>��!�3M��dD�	cA:�:b�۶����F�5�BS�L�3)	[�twf�֣7ߢ�uqd/������ެ���1J��4�҇j��;PL�1�ҍm��\`��q�B_!����T����$�)̭�ᲊ\A��go%^���,N����;�a���uS������;�\}���u���*�=+{��©r��`@D,�*��E{8��A.S�x�ׄ JI"�0��we�<B��;�J���(]�0S��ҩi�%U�#ʴ��keP�B4ԭ�[B���Zm)Q7E�m2"�uQb*4��D)9vU�AK�B�UT0��b"m�Ǖ����
���tZZ��������i�a�"]J%ܨ�UP�c��FUJV��*�Ve�"�bj���Ub�EEH6UU����+�����[(�T"+TTEQ��T�X�Te-UVfYB���Q��7E*��.���X�IS���;gc��V���N\S���ril�ӏ�����S�>�Տ�f{��ߎ�jأG����y+�	)Q��+K.�A�Z5;����H�quG�h:\�%���벣cYCN|��]F�����91��ݤ �K�tQ���8��L��=ps���&l���C>��5�c�Y���N�������V����{�!�s'�}s%����7�0�Zәt{rڐh����v��Hz!1z��1����Ǹ*:X�h�����=�Q�_kY��Yr�9��n\.���<��D+�m<;^`Oy�R9�J4Q��z����Xt�8��^�~�{fﷲ	��[��~�t��� �U&flW�ʺSu�h2��[G��>0���_j�p��,D�sY8k�(At���^W�eY�~I��1���{(n��Y=ݏ���^I��F��);��6}�*�-�j�
��=K	��^�&�ʼ�;�|n��iq~��T�|�*�����6�I�,�:�uv�m}�C@�M�щ����I��Z}HSek������g�ݫP+s���W~K��W�vG�;+�b��^��s��=��?m����	�������	�5K�:�
g��(��w������^��\��,?3W�Xe���R�C�jT#jFS�_���>{?E�L	Ŗg&3��D����g��1i��p��u�]�e�w���!�<}�y�=cؾ��u�/}�W�f17|\���{��z��<O!-%��k���f�oڣ���4U�v���񢎐|����"���%R��R�-X�P���!:'�b�������ᔨ����+�	`�<j���xk�a�~�K�1ELUڗ��UC���\� ^>&,��9=jaM�]��Օ�F����_u���)�$�7�'AJrb���f�j#mE�_�oV�o��sP�-
��C���ö��G����P<��v^l��{���X숿 �9�8ݙ���kI֕Au}�~���L85{l�)2��ԧ�I˘����d�򴎥�Y|[�$n���]y�"u�s���SΜ����3�,m��M�l�O_�����	t�{�87�x��PC�"s�/ʡ�q��9�`������Q)�5���Ǧl�>��+Va�}�W�nv�����va������U��=�%pa�q4+=�K�K��MYҌ#7�$�T/CgFv�	s|���a�c�k�H��iLh�FFn2Y�`�[�K�f^��������^~c�C:u����m.TTr���Dd�s�\􂷵��of�tw�u�0�J͢�S��wQ��vh���6��/�L]�	�Wo7c]���6��W�	N��D��VX4%�K���޻���"�����ƻ�3�Ot���p�/���`��;�T�w��/4!w熼y��|��	�4r㧉���0���c+]����ڶy��H����P��Ծ��
�=Y����O t񳆖; &�X��֙�x�d��=,�UU_{ެ,Q��D��B����F�x�i�%!�Yz<,Z�Ǝ�]"o���a�M�TGm[�`f��}x�5�^y�]�q񂖓ɞ��I�S���Ū3Q.w�����F���������j��z��k�����0����ʫ��W.
��\�S�U����"��/�/f�H�x|Q{޾�FV8t��xD"o�Kux�c��r��s�嗣1�|TNa�狖�t\�9�2�q���M�ң��A�`���-�K����u>x��٠�a��Jt���ID�����h�?|{��9�}e;��:3��ӱU�3�J�])S�y���]o��N�jW���t���)ќ�rE�"��m��Z�\�����9g����k�pt���Ǐjf���fT��	Y�f�P[�}}t��3�q5�n�~e����e��ǈ}YT�~[=�������<a���U��uX)�J�\��f@��s7[sM C�j6p٠|t��f��TU65��B��vΐS�2�0�J5UQ�Z�@!��k���@�.�d��F���k0�L�:�ÉS��ڸP)
��޻5����ֹ����*U�	}^f�z����\��bĝ��|�^n����#)�Ծ�H��C�N�8�jb�Ɔ��LZ�a���8i��Zu����/]2I��Oy�q�l�yQ�e�F��>�I�8��<��:�m��B��lt�v7�����N��z����E!i�A���G�4_=;��_�k;��=j�j�4B��Ը���:GX� �nY�ӯ�u�ĎF���;���s�;�rf�qa��:IN�ћ:��9ȸ����l����,S�{M��*��VAv�M�8��5�d��I�g��t�mʒř.�ߨa�L��!�%�Uוp9ޭ�{����$;y4����WW0�.:l���9���v��1Ʊ3��VpK����I���׌[�\G���V_�i�;��ʎ��s�9,�]WN�2��/�O����m�>�cyqQ9���aG��������.�y�>�p��0Ϛ�gk$d��L9�-.��eV���w��f&�'�>V��w����$�y��z:�T�\=\pZ�^@���s��*>2�,�|��d�_Ecv#E����/_Z�ꢫ)�U+s�y�h�l~<t�k���8F�y��s��f�$�~>Ou�"d�	3.���T�㑮E�zH���a�^�X��ƅ�t��������)��Z(����B��U	���[����Y���6n���VU�e�g%Q*������ay�qk����Шõ�r6�T㭕�-mF<�����l�GH���;#��#^_��Vo�����]}�,�����w�B���xR�%�(z���廱�Q|G����q*��s���R&s��۔i���n_�f�ʝ�khʟ�7Q׋&vL���$��T	��"��fD�;�M��y798���B�N�"��s�!�;6��/�^��	����`�e�	]ZD.�E����H"�_]Ͷ����/���$xU:��_�����,w�;���X�뒌
����N��f#���ݎ���L:p�V7�?��=���1��f����{��9g,4Q�os��XIz�lTZ�&�K�j�Al���\�^��v;0��&��c�w!��V���_J���;dy��<��f�!�q��o������%��;0:C��8��|�
�OH�\G8�ǭ�+���ouU��Y���b�أ-abi�����)�4�e���)�{5>~̽w�����K�e2Yz�������+7)��y�|-D��a|ic�j!=��T�q˛}C;l��0���.<I�]�a�\x����n��7�d��Efφ�Äz�������c�]-S#a3Dgn�I�9�?O�f.q�K9N�{��iuQ�z��H���G\�wO��6���7N�,���˄�ȩ�d�m�O��N�{E-�ۏ����w��-K���O�|��x/�)�2�C�+���x7�Ȏ�^�,�/�./Ǐ�Q�8��=����K�/N�X���p�o���f[�]/��7{�H�j]���n��c��{,�&h0�,d��ź�v���'��w��"̥Ռxyo)�a�a���4���=�Y��Zzvm�(�ｏO�2q�fχ�E�ct!�,TYȻ9��Ƅ4h�z�����i�ǏjgOڄxt�W݇;��Wv_jk�"�0�-�G�/�1�*�e�<:������y��<~��v�AK�k����/!��W���[]�ܼ�{�HA�6f*,��8�4|F^�+��]0_D�~��f��G�����c9��2;6\������U\��ަ&6��螺���˼���ǝ�6lv�v�͘��.m��&�*���m 6�c>��9�C����a��0�m|\xh�'x�;Ћa�����R\Ҙ&%�
�_��=�yn̵�ִpmL��R��B>z��_Ok'A�ƎM{����{��R�2���~!���S˭}��g���\z̝(7jqLX.z�}F��ݘk�)}o�Q���#���	��=>���?BM�Y�~�Vlؽ�(CǆzT���S"aQ\���<	�k��.�<#kR?i�L�e�=\���ʰ�1n��ZJ�<g$�j����Z�`�K6\���KʾW��i!�$K��v�yJ�;�8-ʒ��*a�@�ڹ���Z��X������B��Hw�L�zy
���gî0�8UmW�A��I�G�׎��?���T�h �;x����S������I��i�ǘN�v�<�a��iM؃���v�V�Y��gg·a�����_�FCG#�Q���wH]��Wr]�Wd���oH[l"��<X{�͎ݽ��	�DV�҄������+�_n�
��q�io�|K�6��&��3z�ƏA�{%��}�B�^����[9�tfa�g�[�kjF3jLf��w�M�\L�3�҅�e�;�9]g�Ý�;��X��Y�u�'2�r��ܣ�&^�n^��>֗N\::�K����xm>.lTۺY�ck�4���s,p�lR�3�e*t�����K�T[����ӽ�$�c�iΒ�˫}oYO7L�']���Kf�x��:����P�Hܱ��I�+ef:}}�n��t�r���M�]����l�l-ua��j�\О�f�aaie�g3k�/.�ѵ��F4B�y�RI$�I$�Y�7s<74�+�M��؁������	=��(�C�ڳQߙ���M.gH���˼��<�15�]vJIcSP�9I7f��twCf�k%�#F�^�xx���!���R�pX8"!�.�'�d[#�Z4]hKU����B��_<��[��,|�3��.�n��J/�gN�CEvд��גsg1����r�m��W���-�>�/wFt;1vʴ.��}St��=Z��:T���}r���[Yݳ"��M���.���"ww�JG� ���5�P+zX�`��PӹA��6\	��p�u�����g7B����{xz��(�l\�.�S'l�h:7G]#!ۖ0Q���-t�߭���^�έr�<�������Z��éGm���:Q�h�Z����Bb�Ђ��Y���k��H��x�ڍ`����$/�����;k�'z;��j�V�)�Q���ٹ��F��sK}!}�9��9�6��ZJ7ϝ�9�̆�5)�`��杶�A��hEbm(Q�.�m1DQ��*��uB�"��i)U��H�]SHTb��#�H1�Xb�st��e�*�b�0DQUvԊ���
#(0DDW�R����EA�R+��2��EX�1Ԥc1T�څ
�ˬ�ġV(��&
��$p�EEFA`�4�a���E\�
�DH�Km0��*1`�TUX�E4*(�Y�R*�1��n��	�)@Q��������*����o~���	��3w[!w�/����\2�P��֨���噥�dO�>���S�>�P7���+�-�Z>�MY�c=��`gO�<F���ᇵl�Xv������5�W���'76njY�ew!5ܬ�0�+�t���{"���Lc6Y��mqQ���$k��j�����f%�N�ǀY1"��&�ֶ.<s�x�(p��6y���o��5=Ss�ճHV�^]���.�A����CI��Tŭ�R�^�8�U�6i����?=4Q�@�;��I+�%nz�=\��Ȫ�?-93ʈ�_r�����
�ə�ӥ�=���k��5Qʌ;^;J=u��W���{i���õ���w<?uvDk�i��˾�մ���b�����%�
z��J��X��^T��	�=���n�H,�!̹�^
�*���j���3K�}���e�3W�U�Jm]%�������=��f?37sf2c#PdO
sG��O�u�	|xI���;1�X��k�%3ns���|�)Ӝ�z�dV��e�4E�X��:E���)x�xt�ނWWz��!\�bZ근�*X��Ӳ'�����O����V��@�qHYǴ{��dv�m���Շ�cxQ�+�}�O���%����T�G!ٶ��L�T;c�3�k&�EZ�&OP�����D,6}�Լ~^C�Qg~ŤV�Qan�&o}����]ݹ�C�1�����|Y��mi�k��w��=�eN�͏L8c�M6�ݯ��`��+�7�q�5i�QK�$�Cg%
�5S9�����%�����]���ϋ�zw�{l_��@�C+2j�I�W�ثK*eǻi���IȔe�r�f�N뱵�CGi����cډ;)^����Wg$�'Y���ޭ�s�!R2�c��VR�(u�(NM\6wC /l&�˔��#2	��VE�ޞ	]�o��õ���g#|i�R���\e��݆��Ci:����@�53j�;B�b*��:�L��Ѧȵ���������
�$1��r������!�2�D0+3<I�gO�-/�C�"�GUY�Y�56�����=ͬ��i}�9x�XO&z�?�s�:�����SF���W��Q��0�CM���0�5��8�׆{_Nx����'�#����L�ޭ3�̷���6W�d=��f4�jRO\1\��W�7c�l������N���a�q+��V���g-�~�0$,��� �iY�VOM�:%��)H����)k�LC��ogBB��aZ�DVo�n�z�Y|x��hA�y�.]rfe����$�TTY!�_��y�a���V�/���t��}��YǍjd���x����8X����n��0��HT�Z��a�g��Իe�ї�=4������N����-D��F�N�n�S��R���\.�0�]:;CJ��"���b�ώ�'f}hx������~�����(x�k�u$��{#~6���ݪ�m�į���,����b���x�4.���B덑�}ڎt�~�6�O�C2����ɉ��s�\��{k�$��]V�_}2x�5��S��<�g��q�i$�um�L�xelg�a�1[�=u�0�� �FmXzovo�~>�~=Z��m�e(��z�8t��$�%a����.�.˱�.�Am.cWfvZ��#���$Z�M�r\��-q��^��9X^��ҹ���3H��w����ZFx{�6�+���T�-<{ѽ|-���\e������l�*��pHe��7z��jy=wv����:2&:V+�ZY���|�aRH����#��L�N^;pە%�2}.\܉��ɍ�Q�Y�]v�J�#C�2D�=2��<@�������xf�c�4�yݹ>�<l�z�æ�	��p1�{�P��S>�mM�O��5w��_½��_rd����=���y_$;-s��x
�{�h�6Q�P���aֲ_s�'�ea��w���EyL�����ϚŽ9��x�8��c�a"}K�g��U_ow��u����E$$��O{�Hp^#P�7�[�o{�ܻq�"{<E����-:X\�Ť�="��c�N���*����菻}j����ȃk�]u�f*����;�`~�#��&��G�.5�q��g ���{�T�k��Z�
�w@ʚ8��1A/�a�i�F��c��f��c�^���馅�����fds,޼�#D��R�e�P�믶��-�F�?��������s8b�O�x�>�<D��C��YDP�㧧�ơ����QC���T7��#��|~)5���J'fo����f�i��'"�t9��5i�<������t]�b������t�o^���#gM�n��Y�;���Jw���va�l�W��t��ɇN��xt��0������:���懍kMD,�_�7�AVèb̅]�:�Ь]/�4-�_��k��3��ܲ�נ�YUω�l�nN�2'NtU��6o�OI:5C�U�<]�^UyFM^Z1������Y�`���ܘm���6���%�j6�EGjV?Tsb�mq}�ȉqӪ���4t�+vs�o�]t������)��^
wټ�t��-}�;�R=sAN�� ���pQ�����*�ܣ�)�Zb\p��԰��x�+,�x�"����Mb�3v�T�5q!ҾC�q�e������g1�#
�cj�����7�w��#�Qg�X��O�j��Ez���8�E��[���l���CƁ��7x�ŗ0��� �|���]��b����UW�}֞�r�$x�DP��;C���к^;)����}����G�{o�=D�ܴ�ǋX���a?<;��o��y�U+�w���-�堈5x�'+{�@F�>4�26��\���47��e�g�E�~C^�S��;��F-vQ	Te�Zi��J������9���z�P�JNP����^�]< 3��^���V��.��Qayx�+Qb��z��)κ�j���uY�x̫�[�F:��V����)C���kn��wy�d��f�k���J#?��p���zx�߶�N�)&xr1�'7
	��� �pi�?r��{(�FR�E��M����_p/�!�`֊�=07�r��EVCW��Y��ר�jfoy����K�f_R�+�O����p���0�dc�͞[ds^�ac㦃��Z�\�].<Q�����Z��ݾ	�ԉ�Pó��uļ�8�����JG�Z��>N�aä;d�c��2�!R��my�hg�ʞ��7��vR�u�^�;�;�-�oH�(5F�8h���ٖ�o�g�
;�Ȋ�E17�ZCظ�h���x�b]t���FY�"��(&x���t�#A�|t���4��G�z˴�m^ܓ4�j���q�0�O��Y�)"����b�gO� �u�^��`�vM>��ѝ(�fM�Gh���Ŧ��;z	�侈:�plwe������_.3��D�_���JоZ���c:�����<ò{����`�ʎ�ǆc#[�]k�C(���sh�P�'��4_��0�-i�40y�h�C�_-�i17����c��� u�X�e5E�"?<=k�w@㔪�a�^��w-���!؃�Ϲ@5�u�c��7I�M�<"�a�� ���X<9x���s��f���R�����;�E;�g�_���ٹ�9�����BH6�Ib̹�1Ӝ����wD���a�Rzy镶e�����I�&j۶����n)O��.�ٟ4�D��g��zE���	��<�u¢��E�Ʈ#�dO�D��	�����v��E�#ʴ��4e;V2�&V���γ��K3��m� �Jg�#hN�7u�R����d�sE/�I��x3nX����
�2�֧?Q����m���m�u��b
�;���O?Q�l�A˥�3��s64��-������8Q�4�35�c�	�uR�;ٵ6���>�a�,4|G���.<{J���`��O5ݙw�|���m�!J\�,Z�r^T9G'��XH�o�ru^�$Y�΂Vn|ޚr�_:��hZe�@�;��ɝ����$��hY�����[V�_x鼧��L�y��v�S�<]Fk�����P�j�m)�����W6w�riad�B��J5q��w0:o{m���8�b�T�N��Ra��C�t[�1^b��A��P*=t��\��g?\d��/��"n�][�b�}�~0v�Z���h���|��]*�b�Ò�P0��K/wY�k�����o�8昄+'wn�2b��o�I�"K���[�2�G�o�/I6؜�˨�\r�&BJ݃9�{��X{z��J��wP�;7���E#9��y�`��
�Mf"-�C���g:�:���B_S�P�8���_,�1��uLߚX�݆u���
��f�Nysz��Y�E]��:d#�-,7]��oG��Wwe�o_��v齪I�݆�-営u+�����������0����f��;�sla;l���L�*W��� ��'}V4]vL`YW#
��B��Ox���&k�Ֆn&~�-늫i���jݞN����_KZݼ&���3x:��)o���%)X�t����!ޜ��%���i!yr�_f����<�Fɭ���_T	u:�g�nfN��T�`�Q�U�I$�I$�I.����/�����6Y�t�ۆ��r�"��ՁV�"�dpA��g�Xm��Vu������*���+6��X���UV�bc�6k-ؖM�B�X��h����%��2���V��i�EP��ئE&���.�U�-�^E�ƙ� D�l
pPX,��YK-F��m�V6rEs4^��T�
,ݦ�H���_É��Ma�J
���t��C!f �@j%�'(4����2�4-�xM�� �%&�d�DLL$�9/%XƘ���q�HU�XF]���.�˧K�)g��*�B�w/c>Uv��M�F.�X�p�褤�b9tRUu(U]!qU]ɒ�5f�'%R7c��4s-�d�@���V�v��V��7x޷�{|�1��u�Q�%(�5H�`�:���),��0�J`"�����(�"�d�T����5U��J�U����B���b�ġTL%!L
Da��,������T�ADV]R��ر"H��QB,A`�b�uJ

D�1TF"AZ���H�a�R��.��T`��4�B"���E�*�U��:��"("��B1"$X��PYX�����-�)���T�JJX��L]KdyE1H
�'� �H���,����)Umb��!�{u]|1+�ђt��t�E����ާ%���/�\�������ۿ}��lp� ��={�om�����n�۾�?��B,�@����-L��ӯ��0g1�B��������n,#uY�m�Qi������y�k}\���^Y�8%2OR�>�̻?A�����c��Y�%��#�^.�$Q�Z}��,-��x��=�vx�'K;͐��KŔ�pB�����ɜ�o�Ϫ\�[6xb�k�.;wW;���'�'�K�#�qc�:c^&C�;�&����v��5������	��~�暵�+��<�iso��0�;�����F�.��֞�F�����չ�Á�G�E����T)3wQQ�N<p�|�j��㧭��_+����	��O���ٵ�/�'^��/Yx�i�/8G�+�{5B���iʃ,�9Z��f�C��"�yr�Ԉ��ӽ��%#�]�}��_^v>z��o�rt��@�h#ٯ�x�{����|Q��"���&tʧ��m�e=`+oux��>�Y8�x�;���(٣��
5��_�͡3q�6T�*R�i��qg7g:�aܰ�8QeCH�0yx���c�Udc��? Qݹ�ѿ_ӆ��/&5���e�2^��hJ�zV���W��%����X�,�ڀ�B�zQ��?�,Eݶ�+n�Ș�}h�¨Q�/�g���pj�:�WK~�OX��4��fݕ�(b�Ƶi�.>�d�:aV9�;�=�(8��v�#�Ʃ ua��2)����3���5s�����5�=/�K9�X�=-2^��>��/��_x{�v5��&��&Ž�P�a75C;��<x\��l���֓���2{��Ĳh�!n9sH�BV*�Sz��,�!�����1���ܾ��lO��~�{w��2�M�H�(˕�^�S6M����_@�ѿ-�<wЩ���� 6��Ha�[���7�i�f�Qg�N{6�=w^����,��cYCN���R�b�q�0��I?Xꢃo����M��,����=x����x<��{]�*˳���6ڬc�չ9�~�����D�/����~>�ظ�ݛђ��Պ������=�B��/��(���z�+/ޔ��;�d�}�=�D6tßTa������ vcH�cj$��WEm?MLUs���0#q��4Q�R�^o��N�)Q&aP�U�p���s��S0��c��3ݾG��!�i%�O�6}c6<��zs��cҏ��S��~�RweM��n�7��+��{A��Wq�Zj��5F�p�b� a���g��h]�@��^��:����	��S�lb��Y�QG�@Ի�{7?SFcI��~b��_�a�ǎ��������]����+��,����,��b��E}�=5�O��*���q����ᚾ�p�w��9I�~\��{�-^���UX]�-7��h�\�A�T�Q�-T\OLȟ_��ܣQVt^�<�|�ov�7���=!�>>2��܄�Out��n��� ��]�/����܋��a�ָ��p���4ÅC=��q����=���"�>7��e$<x��JUҔ8�9m���P&�x�^�!I�.��k�O/ �:O!���/V�Y˯���ɘ�O���͢��C��/�ML��mo�/M���x�&��9/���-xx�T�����L�<�J��C�L��W�3��H.�6��
��ۺ�ixwe���6�4^lX�D���&��!V��
�q)֋�CĻ1�=J�늉s�ՅH��=����`g@��<�}�
�����E�s�Nܾ�;Ż�p�ɼ��9�[>��cW,�s�G�h�����˖�{����*7KH����p�HJ��_�����.��ނ�g�˜������#��\^!��>��-�h���;��r�W��W�0,�t�x�g�[��7�d�&oA%V�F%�{Ȥp�����8�Àla��P���OMy���+ǃ@j�)�o��a�k�1��[sxsV"��/�_�?E�}����؀�^��:��/�ˮc�k����� �";�3�q9|W[�߬��ɐ��ϝ�p�+X�Uz�q+}��V��r>0��%��;V��A��8Y��y�5��>�r�����5(�b9®�u�
Њ��nL�I5�;����#�9woXݾ2�YO���d�j��u#�(9�J�I���C��z9�f���Q��Oҧ�>�n[��6~�'����p��׳���[X|-x��1͜>?kU�>hCv��>b���[� kEK��8e�	��*:�M��:S3�Dz��xq.1�h-��Q��z#dW!z���M�#�k��K��Ut������_��j���5��@�>i�C�9��n�X�Fj�׻p�dZ�<~6Q�"�w�4��V����(^���)�gvV�U6��m~a��`�L���3��?���=˕���������3���i�}KH����'S�2My����:�˟^���n�P��l�"5\��
�7�S&cg�����'�^�}��*���p�����Xi��}���	1'����k����U)�����p:ky��2]9Cn�ۺ�5�v�{Q��뼹�5��]�)�����N�$<ĻNt�Y�Fr�<7l����\�g�dGHt�	������=�1��}+k�e^�dB��a�|T��2��K�0�C���j�mwM��`��q#ج��;l-:o珌�?��T���Pb���׽5>2$I�Q9[>3\^EKγj���������v}95��,n�4�D�t���i��Rw�ݛ�����(�$O�{�Wэ<Q�_jѳ��x?�
̙�V��ǆRoU���F#��I!؆�h�e^v
,�����Dx�t<GU�' U��������o/LwI�$U�'�q�yq��'�����i b�B��e�a>��U2���T9��9PoسH�[)���M�mp5�F��O.���tJ����k��yvh��)Z�~Xuoe�J�j��SXFk���Fl��4�pc�wc{��lJ�j��s:)�	�8D�����m H-����..�.a�c����0�"�������0�W밦�{w��� �2�C���Xw<��m4U�,�A�.d}w��]�o��<�݌F��5�}�c�n�8C��i���;bW�FJ��啲�C�;*%��=�\����G���_�B��{u��^�r_[�{-�D���;}4/|���p��!��b�Y	�Lէ�[�ͮ��r�6Ϗ�ڲ��6g�9�S����!��F�&��߂�j�q��+嚂7X��s�8~��7�G������k������Pv�|�%Q�S%a�!kґ:Ҵs��<��!ՌF��q��
:F�h8)ݮ����7^rVY
��3�im�E��ݼq��1��.f�b���)AR�U}� ���1���@f�P�M��^������:���8����O���W}��:H�����FƠ�1i��MH�@�q�3�������r[E�8Z�=�m���Q�b>O��a:q/�nس�i����Z��M�GLb6���ɩ�Q����0Km��|��<��t�C�7�:p�,�m|���H�!JΞ	e����=^l\KW3�*z�[�+<(��[gx(�%bǗ��'�<�(�B���>���P�\ts��Ӯ"�$yLU3^�8�LU��^��KZN&E�ϵ5i�Zȧ=]���]px~C7c �����MU�8Gb����WO�]�o�j��#��ǈ��!^0<E��!,RӬHZ/�쾯_������cH�^�7|��և2��LF,�����a�n�fLwv�)*���o+�gv��\+T��S�!N�Bq������;�*��ݻ�5�4T�۳="���N�Mgr�f-�S����Y��-'�Dz-8'�0gg��*����F��	ac5لC��O����=�!}.|�*ȟt��x�r�9�;P��;j���֜�3.n_TX�'��J�C�IC�{��!^^1.��ex0p������f�����,�ij����b�F� ��6�,��p��L\��I��~��=�v:����4�$�a��g܉��A͜>?kU����}Z}]Z+ޢ�y:����k�O�g�1i,!�K�|w����W��y�����pu�7)���HU�>\^#��|L�P6�r2�y��2�-��"���Jً�k�i�b��Sޮ��+�e�x��߿���o�UB�3�-
���Hh�b��|������
Sdo����`�w7��l���s�Y8�xإ�����5��mp��]aȷI��q��SB�����ξd���+:���t	�X,�'
��R(-N��������F�bY�Q��$��a8��>���hv����Ɩ�vtF��5����}�e������Sv�H4�B�+N��̻b<��I"PV�����/��W^j�u2v��S�/�H8}���n���DW��:����V�o����J���i؆n�{;�u��@�%�Ӗ�ۤ�4�p��<�s��¶w�F8�� �� �5����|�a�G�>��';[�ML�Zr�2��z��!v�	Wc��emnw����z.T�i���\]�򧆵]ʮ �LiF*m��n�����u�إ��F���pod��u0�gw.I$�I$�Wf��ۙY����v����-�y1�j�����F������p"ɸt�Y�
U�8�ʱ�Ջ�lR���x.��P��+&[�l+6����A��Ke6Tg`4�e]�)��3p�;�f�,����k�B��-�h�H#���,���j]\B���t��Ab���`"��ѱtJ��V��cp�j�
�ˌ�v���H ���ȣT�D�EQxJ�jY��V	�o�q;j�CI5.dl�[�
2�XF�tk8��v!X*�ˣ#�c�	F�nP32�՗�6$�Qe1v�,Ʈ���G-0ٲ�T+(#>�%�hB�&�ZA�wi�;����4�4�w0�)ݡAZT�9�e�B�I����gHܝ��#'>?�I-�FM�.���I֙-%2#E`�,P�Ħ��"�z��*��!L-�U��0YDRaH�����*�)���`�U�(Ԥ�aH
*�MU`R,��)��Y��lX� ��dX����
�IJ"�y����e0RCM$,Y0��UL"�$0�F�
]T
IĥAb�!��R�X,\SR�H

�B�)���) ��'� ?|m d�rvN��`ӕs�ҳrT��*J��e�����u�9'��}�i��g �a(U����W��c8#]�z��H�L��:��(�����n	�ˢz�5E�A�6�}�/'k�=m�Y��e��z��oRe�����l�h���-S�4�n9g�/�$�&2���,��2-��܎d����=<J�D�R]�6�>�+��	�� L�
��5��)ۙ�q�ߩf�m�S< f��*�7Zfnׄ�s�E��@|J��T�O_��������p��_��ۧ�����I.Gh.d_�wB_1��P針˽hX�vY�O9�¸+�(��!Dѝ:�o")o��b]�r��7/����`U+�Gl���h��DE����x�n����n�@����Uȧ7Y������=2�:�=�E���&/w������x�M!�r]����H��;�U�v�l_�U�(5��92�1�
�e���ї�����	nw}m��&�t��ONNva��n2��}չ���U�(�O�e�;a���?LƎ��"��̣�uj�W����Pn7V��\k���d�@DM������!�TF�]y�܌�����M�NCHC@��������ø���㳣�v�,;�3E�2���w4�.M�����KB�6��.]�r�Q�u��f��r��h��-W8�ﾯ����0�Bo� ;��Qe=wQ�m8Zސ_;̢:�Y�e@�2W�f�E�2�b�\��C��F�xٰ�F ��:8mS۳�#�ᓪ���a|{����K.H�V���d�p�a��\�Ξ�Uze��93����w�p�W|�ד7�a\;j3':y]�Z�l5Tdh�	9��m��:�cQ�1Xʽ��WW8iR-A��IE,aJ�q�͹�z�b�2�l�D�1iT(c[ʪ
+�d�Ҟa�Xn����P�(�ث��ֱ
y�2���r�U9b�`�{�NH+I]X-�W�ʤ�hY�0
sq����<��u��Y��YC�pasy0�e֚����A��_Wݰ���w�������Y�.��
$}]�xͫ�\Gb�ǭX���-������֍�x��z�&!���s�̿��<s&��p��E�|+�Ki$�C��q�r���J͸W�íjaj��gx�J�U�Ǻ�S����a~����B���v���e����ӻ8�O�u�$2��X����k2��ǹ�M֗i����R�wAt���q�ȡ����P�`������gF����L�U󧲱5q@�`��5}�Q��չ�-P�CuJ�N7�����F+܍�]v��١Z#�T����U�]]�X��U�F1����w���կY��Φ���ԕ9i	��sw�{Q���� '�=�GGn}	��(|�!��ajl��e_<�·��b�)3/f깴st��.�Ū��g.���0�Jk���%@�X�!�3�z��3r�/xH8 {[D�PzY����sk�	^���%%�kl`�BD��`�E�P��L��zlk�m�egd@�m�u��3��L4�j�����V��V{g���ꊋ/^��-Odtn�x�G��i�˦06YJ'�� a;���}�5�i���=bξ��{H:9m�7����L��ݡDo
|^m(ta��ur������z�#�)�fS��y������.W@�DD�&<��֟~���S/��}m."�m�$���z����^̡�x�-n& u��l�"�E^�>�����%v[QI�����pOt]sed1-��<�W��z����y�������d��+S�=ڪ6��#��Z܊�;����򇵵b�4^��k\�Q�Jp��M��w���3S�f?-+ ����+�Qh^�ޡPc�cN�E`b�P�0%�)��f�j��	 ���w�٣�OB�l���f!�����t�-_.���*�˩s1�w4��P���@X�ԭp���5�cRV&Ï�����q;�/��RQp�\�G����3y��Il�Ǆ\����\���WՐ��Փ�v<�\���jt��ܥ;*q^�o���5U�3��^ˠz�-苭5jւ��cd�r��8IFVF�h۳���s�)�c/n���ɭ��$���z�J�r7�G���ǅ�FП�������`ͣ�Ѡy�F'S�T0���GZ�4�n�`Z�E��.�J�4m�y���.�#}pV=�]��:B�$�̠^c�n+�%X�3~������38Al�ƈ-��HuT�W=z5�C��9�7j�9�3����dtɽ���L<�j�^;��O3�Gܫ���\�sRBeU6_57C����ص��}Éf��ڠ{��YB����{"�@͈�+����hh�V��%��S�@_R)�\�m@�S1�)/�=��Q-�����1��=rn1�����A�;wY�^택\<�q�j,����m�
s��9Gs-���[Q�+Nu�k�J $D���g7����B��p,N8'���s
�	�%�ec��:u�������(>�6�GWj$W��Y�
xVp�i��X�e��J���A��o���X{xb���!W	�J(TRtO���˙4C�5ܛvw�Q�Q؅]Q�q�u�НnVIT�5z:�+�����E,��'ȟYv=�1Ǧ�a]N�x%+ ��s�=�37/�����yF���{��p�
�+�&�|]���֨R����dGbJ��
�c��c�/SW�_���YLc�[r֖m����)Ҝ*��sL��d�����`H��%��K3;�y�
����$�d�S�Gu�:C��)�u�#$�<�����]�vٴ�8�]��Y���f�B�f��U*Fre ��3X���Gz�[�T;u�1_W`m!�y΃C|zZ���U�e�Tw̦��
�f��P�&��M���\�������q��X�>�KFv����^h3�t�u�=d̮��7�=�6.�8�����5,�.���l����'8(L-����5oZ?F%��9��*����³�F�#!��@����H�^<o^�³����A�;�B��^M8�Yח4�B�$��|+��h����];c� F����2�
�xv����Q���n��9����a��{Aw��'������F�kX*���7�B+o���{H�nN���E�@z�{+�.���yM��wm��Yu��N�����QJ���'�ܨ9�"����o9ýh�7o>�2�T���~�i?8�:jn�^��8ޢ�:1˽޾��,Ʌ������6y.j���̔T������]����v\�����]n�%5*|w�l����q�fJ�Oe
������Lmfl�ae��	]�O	�C��U2Bo�fm�Z���s4T�un8bԐ����C7;]!í�Ia�Y��t|�r�L�9L�����B1�Y
v��T$7)۹�QSQ�np���;w)�!dEr�X�۫����*R[�{)@�2r�J�T�Np[��.蔓����0J��2��TH�����v�o��ӕ9D=î<YhE2IOt�0c�X�u�c����n5*�P��y�8��g-��F�����i�Y�m^�E��ZBDutG&���M��Q�N�|�8Fœ��[ΓaU"{oqt�X��NV/6����s
:��AHhCn�co*u�,k�����
V�Kɵ�X�J�4AYif��������7www����Q��Θ�t��!���M������*˻��E�I��UW�n@�?0Y�<M����ljn�^X�,S��
�]%wF�)��^K�!�m�ּ�����n���"��8l���K��V4�^f&���F|i�
!2��I��L6�*��`��Rj�YQc�����|�^}��\Q$ʲ��s1�AQ�*;����61Zcwc�t�k G̠6���L�m�S�&�2�� V(3Ղ�[�WF�'��rK��%�U�}����U+W�qA��	�喬fs-[�U`.��zJ[-��I+]��o����l�HH�RU	HES)*0Y"��Q�
fP�`(�	�^(��Q`�Xu
HeJQ��TR�

 ()Qi�8�)l�$��j,"�����!V
E�`�E�E�X��S�Yʩ	��) ���r�)�6�BH��$� �E�KaJ�E��-%�Ud��X���*�UPB�`�q��@4��B��˩��^3����=
�2���z=�h��sw5.w���*1q��)QZMꄺxѫA���>�$^mѷ���'-�2�![�&��8�
A�@�!�;6�m�j�M�}8mV.+0I�aw������wS5=��ޱo�i�k�)�gbY��s}ۜ��b�'���g��_0r���t�X+�c�����;gH�e��g���뭆!�!����N�;�8 I����#��U騱q�	�g�˵�M#���̡�v�PT�{w�9�n�!i�C�(��抎C2!� X=(.
�..���0�Qy8�w���h����pv�$����ښ�<{�:���7�i��Ӹ#z1V�Ii�e�k�c�f��X0*ZL�A�v��c�`�r��� �Uxe����5\����^�W�su.�(ܽ>Jg(#c+E���k���8��8c�����DN�*�=�'\����X��uXsy��WGV0�/B��pqX�p��j�6c�y�3�R�/K��d�e�D��8�.�n���9*�k�^�����h�֛j9�Q�l�)�tjx�ݺ9EEK�S��je��ꮈ���a)G�k�Z�-�%�����[QA+P7t���Y[/��e�.9��錀\^�`ȥp��s��ͳ��y"9�"�·��7�{�ąM�{�Ia�==*���ĳ��?�vh=ys�(�^��*�˩���m��t.\���":�kM���$VhU���M�Ν��J)淭�.�%<G-�E���Ӂ�8=V₨�ᐐ�	�^z[�
�gc��O0��zX���aw.�e�盆,��#���=p�_LQ#+��Z5�f��\CMoj��!�*IXvº����T���W�J�58U�^�x+rkYb��������<�=]dA^��(9���8����_��\�UBANW����ы3ˤ�[Ԓ�4i�7�{L�`ѯ����&��q�N��ΙW!['p���oڇM���+�1Rk�=k���Ɩ�L�`/7�5,�����dc/0��d�d�K[���Z��|v�o%�޶8�_Ov~�׷�2"�K3��6&Iop��*�8#4l(B9-�����ў��>����S�D��9梱�R͎u�Țm���p��w#��[�9��`\$F@��>��w���^S<�vdtߐ�֬����=,�Y�`��U7���� ��׷Q��Wӆ�\�th[��#�+T�k5�v@H�*�n�T��%dՀ�k�e���^����j��î#�	��� �����P�l�$"������l��u+��vb�����y|G�)uE,�}��7wnb��A����:�`�wY����7Җ+��G"#����2����Z �敭L�n�����)&�w��2镓�-�>�$%7ѐ����˫.t]n$�r���=-끙�Ӭ��-�7�{^��N��z;����o��\S�WW���تl�U˝�6����!��O��i��TQ��'i��K9�F��c�]�okdkAR3U�&���&Z	 ��w�T��a|Ԣs+;S�*�uTo#���¹Mfi��ߖ��+G{C>���8+��p&�3��~~W�t����L	�c�����&�m��{�ن�$�-�lT�Aq�%�?w]�.�^ˀ��g���nbzE���1R!�ęuE�!+�l�m!�vՕ�:	��1n5h�rM�G�̦c�MB�n���_W2^a���E�%�ݹ�۔W��@�)�¾�x�+�J��z�u��^t+�zYtx�~�.w�e㸁�75N�X��=5�m�`��=�z���ť�5e�(y<>��m�3��5Q��1M٤�I\�C�,����uo���y�6���p�=����V%��f�:Sٔ�A��1:��`�,>ό^p��jt�g��Say{M����y�2�O*'b�l*�O�������_�s1�L��v�	
�ȫ{��U8&���b4�y��Dٲ/��s��n�����+n��#���Rz7�3���l�b�����w�p�v���s8�.���ܺ�����.9dt.WR�PH�� o8g�0i�pF^�v��A�K}[UX8�[[D�9~=5���-P�x#Wc�mIgv�Gm�܄��3����7��%���%wC#��<�aYF��V������;���쳓�Ug�qk���f��(-���z�̽�*,EBw�9���-��b�_�}�O0�K-~g��!�|��f1�U��ū������H�ץ`u]����m��7pQ�80���m:��ox]e=UW�41G3ݭ_T�����8��4I¹�w_��q�v.Qɢ˻WA��.�uS�B�L�뤣�x�i�{۷�V�_m-s��P�ĦI况˅I9VnMe@��ջZ]V�'�����A.�dcՒF�ȍ�t���Vo{%�5���"M�~���(c���z�CƩ<�i���u���ynp�t�����&R;W\�yx�W�aW_]v�I��}�'=17=
��Ǟi���{�+��q^��532JS��PGW�}��v�����G#~8	z�@��;\��1�x ،/�Yʆ�Y�21tѱ��s\)�����"�=�����%: N4���Bz0(E�'jRWB�OU�P�t����j�Ur���V�$BYY.����U�[�ʺѪ�K�к�O���09���]�_Ѕ@Kb����#������4�۶��٘~�w� t��U{V�FMV��D�L�.����W��̐H�/!X뽢-a�P&�UR�ZC�A6k�䈋�*2��f���R-�Y<SrYH�ЯX��%���[OO���uk��
����)#*�����=ؑ��t�Z�+�%����:ٗ�yt�q�m��ze^�yW��wN��C�Ju�I��;��Ȍ{9(�.�!�jK�u5�
iRpds�U��ߦ�y+�v�ÞS.���Dm�s�m{��+f��|�	�t{~����OOm��委��]$�k�/����]��#�Oq�A]܂r{wj������b�P��o�bL��Þ�۬��7�E��KpQ7�}6zwf��N�/7�dY1]�IU�I�v��ׇ:ATbB1���rE�y��Q-�1�b�ZJ�>�Y\j�v�l�u]���o<�h-�E^�'�8�hZ��n7���Px(�wZ�:�T�����m�j��NI���
�Z[sAL���,�6\��J�t�2�G����sǆ����Xy�qw���/�9~U�@�{x�
�!iӫ�h��Qy��3'd��`���{�ܫu�]���ǡ�D�Xi7�l�fc�f,TN&v���#�L����
�{��{>�E���'�V���[}�豥��2Q��#Q1�zH7��:N�!�T�*ZN�`6M^A�5��׵�o'P�������+#����#QNU񡶣#v�;�e�>"�j�Ҿ܁!"Ρ��ͧ�؜��5|:r��U$����P�Օ{2�[���,��h�n�F�rj�HssM��mڛ]D�m�&��4��S�&c�˃rw/_cr�b���J>X��|4.(�jďm��i&�nU����(�F���{��b�SS�KrrYʺ��K�����	�3�.��N@��ʋ�np��=l�#�]Z7�2�F�u���F�N�)K{GV��g�ċ+x���5�u����>�8N����d�W��͵��Iw�o�Լ�m��e��$�I$�I$��M\Ob�꽫��0���ni����Vx��HNNC�]�B��T)	������ˮ��[��&��5��MY�#��	�cb���/=4��	��V�꽬��G���豯���+B%�S��z�Ө2�륷�ժBl�Ӄ2�YVF�L�(��<�:�LY7��GW��i���iq�$˨��A��i��i�z�6>7���	:�]�0v�D�Xf�L@��҅ңZ+,�0�ht�ep��U6dә�fw�Gn��ȮP�
�6�p{�B�	���+�&A��u!-W`�r,ϖ�7rr[������+�����,��zӒ�V�r��6M`��j��!�rl�]nǹ�	�\p�L:����fr��b��]֧^�nΤI2��Z-�w5�II����,x�)$)$�!HTi�� �d�J�� ����*�rIh�([HR%P,��`�2Sԅ
�,-�S X�RJhHn��Pc�
H��d��,P:�dAE�Y�H(�y�Ͱ�0���JJB�E(Q&�.��B�b�R�ZI)��AH�@�B(,b�[(at�Kd�I)R�%%$S�$-� �Y�s<�ֳ�.�W�)Q��v�sqƕ�2K�1�u\�˼���tp1?��O{�3�2�E�*���V�K+��-{�$5�"�G������56�,ыy��]���)��nR*4�K=<��ΞHL���f�U�'!��*J���n���r��s�n�["�#1�
�5vD��A��Ȓ�v����F�( �D�4lZ��е��=4��5%c5X��u��4�@�q�Pٳ�oy� �0�,,�Ͻv����p�^kx,M%���V5�v6ڦ��b��%���L>"6�{e�BY�|!Q�r���}Nv�S�Ŗx�`>���|Nq�����B�c�{aT�	h��f��n�J�YE9�&��ky<�&��a�t�|�C��ä������b���t���:*zZ��v�DV�bv|y���!%Ѥ�ҟ�XX�y���c��#U2F���$O$�1z���Y�ӫ��l��V�Ga!2E>�ٺ����B��qKRvg.�E�*���ӆ�Nu]��,���8����{S|�,�Ǣ�����O^�ӳ�B�I��vf�1�o�J��-��t"3M�7�n�֣�L�u҆.��eE����f�ٷ���G�Nsg��hf�L�l<qQ
�vi>մ�i|����!���t���P9�hve=T�Z��� 壻���ԯڇ<��1�kͻĒ�[-�DI������\1��P�j��'��"C����W�����g7�^�g�{�����Ϊ�M��V�!6�̓'q�M��[����,*��N���M��@Q�zn�<�|�:͞mI��h�c�ȓZRV9�thF�a��'���U� ev�|��3��.G4�P�e�4��I����\Fp8,�k���F� ls=�h�|�l�z�IoVq�X���=lf���m�R���Y[�f�@�_9(�@��D��w:!k냝q"�Cyƹ�R��z�I�D!}�Φ��Ż�0���P#1ñ���<�%	,.���^ި�=�=<W�Zz_:�;9Cefk|	��\
������r��`gYR����5&K��U���[�2:��s��ӷnZ��	��y	��N��� yt�q�m�� �G�N����d�U�=S&L^l�I�� ��SǗ���b�v[SZ�Ï��p��e�qm�<���Y�?(��ʸi
.`<��Gv�+��;[���>1hM�������y�C�ӌ�ea��5R��V���O�Ky=[[]� 7w�cU`ᖭVn�Uf8�܎l#�JѰQ������=�XD��뱮�%Tƴ��	���"�{��}�Ml7���?.��qRrB�͙�a{��_UM�(PpzˇU��;ro-H��l�W����S;Z�L]��IV
��1=nfV�v�vr��eΑp1-&���!���a��ۯ�W�ZU`���,fQF��t�����h7�`�t���;B����r�O4eS]�l�L!p�T��Qi��V�3ӎ��8�}�ˋB�u���tg�譎��3�h95+/�q}�"����Y��E�y�3���lN��kd��;ϵ�٘T�B�����f��I��FU"p��}�4��Jʆ�ҁ����ı�Ggqwt��ۦ2'��h�@��>yG�I�0M��ͿY��g#*����T=�H.$��\�A)3��ϏS������ʡCg��MvY<����A��18&���ʷ]w��g��$�ZɶT�ǅV�������Y�v)o�U�SD�!v�V���y�'z	�����QX�&��0J�y�˶�%���>��l��zw�Md���&��C��6GQw�eEFi�[�Xyh1���՚}VT<����1X����> ��}m�[��q�j�s��Ê�G�ΏJS1o�� ��I��[��F�9ofEO\��;u<�ŸN��;�G����{ܐTd��T�|�����X3p5m.�R�)r�"�v������.��rt���M��B�WuU'ss���e,�/T�l�O\딺��IQP��i��kfoC���d�V��^U�4��I�膪{���|2K։P�%5C�/p���l�΍of�z�Kj���A���9�t.ou����L�x{����2~�;6�������`:��R��Q\��5s����ڔ���Y;OPL��A�B$!��wE������s
'�Y	,�U\#	��F����U�aOm���-�y��ff���ǥ�用��I�U$w:�1�0�gu��:Ŕe0��R�*2�0TZwy���a>��a������T�@+-�-����'a@�|�g�	\��p\:�Y^�Q#�0�y6T���ʥŰH!o���u˷2�W�z�X�7{�`]���ѵ�O&�:�V�[F���A���{��M���w���RQ\L+���A}a�+&B]3�ĭ�]#'sV���,��:�������tw�Cm�l3܈��q��l�b����+S�M���f���'�GXi+�z��ײ �5R������fb�^�_�U�:e��qm��M��Z�X�Bي���^�qO!�`f茸�����Y^�5$�UT0��Eؚ�2l�b��)#��r�ƥ�J��թ��ܯr�=�1)��0{|�ܔ�����f�Y7��҃�s�9��Ⱥ��(2"Z�D��l�D�'�Ӝ���P�Z�بyhT���2t���X�Шk2�^�R�u����ud���ϩ{~�X��x����	���2��.���>�1ŋ�M��L�;�r(N���?F��Qy_{�$���ї�>�=����	���s�D��YW#��f��s��M\N��N`��_4fyN���5/���h�w/����(�y*{FŴ������֑q92��Q����T#a;�6x*�H�:/*�ɫ�`9
���s�.�X:�.5;��iT���*�!#�흨c�bp-�I���Lʩ�(�rTv��z�fc���y� �'�p���y����S�`a���r���E{���I�sY�=��Ǻ[��׮؋��PW�%E:bĳme���X~k;�M m�#*��C�E��8"��[�z�<��Ki�WgM���4"��w퓟���u8�8�6�������IX�+4Y�)�^mF1�8!iƆ���:�|���PUw��WCbЗvȄ�7)1�7PrK"�a�D��#퓖�Hs�fq�Lki����Gz�C�M3���y���ַI.�o(���Tzb�s{:W���C�	,��R�m�i�\m��ٝ��c�)��Kx�b��^o�h�E���za+ڲ%[c*&�7�%����wQ䭾e��
Av�Ö]8w��������@~��
���iQU_��d �I�� x�� �����D�Ԗp�8�V�箧�K\���u�� 	! ���I $?�z���qAB��0�D��]0�ڨ-�̬�!�vCHUP=dF�$r��Yݕ��?���`��4�Z��E�#/9�o�5�����ܘ5ߗa��
��@�A`��5�  @C��Zk�ŏ��t@C���	+C�����M���/��=��bO�M1�h>�B�O1���  !��)����Dv{V���Ѐ����d���>�mHV*�&{)t!���H��!�5W�G���s ~�� ��Dr����#��Tg�p�p��%VEm���W��qd՘}*fw�[��I�_�mm��WK�z5I�G��\����ݨKfl���A_ �}�/����94�d �k.�b��<�U���y������A��f���%�o)�Ù~�ǉdڶC�y:�T҇B��^���檠kx�;�:�!�x�K&8�q�D�EǼ����@B�Q� =�܌�}���LJ���Nu'#�"�K�\�h�\.l�Q�<K�?�@���?C�$ ɒ��c$��CA�c��/ރ������܁��\j��[
�wfrc��b d�;7��~J�M� �W��х#[۬�ߤ~�6�@������Ѡ�>[�Me��u��q^��=��'�x�z��O��&_��J��!�tv�a�6��x� �^��#�U@���_��Z��=��}�?f��:]�����{&7V(�x��@��H�<�@��y��Z��ȇ��n�����h`�6���겪�!ˀo\���)��5.��w�A�'V�4=Pl!�&/;�,VCؖW�4�B  !��/�<Ɔ�]�����:��D8��kH�t�8p��k1vW��Ҕ�t�A� ��J��Ҏ{\�.�p� �$�,