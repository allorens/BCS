BZh91AY&SY�����_�`q���#� ����bG�@              }��`����))	E*
R�T�̊�HTB�$�*H�R")J���EPUI@�lى��Jh�5-6Б-�s bT����J�T��N�*�T�I@UQ P�TP��I*�	UR�PUA$� 4k@ (�:QQH�p�R�D��2�
UJ`5#�`BpgFF�[hb��4���jR�l���-1(T$�
�RJ��P��R�%X�B���_���>�U%6zk��Nܡ@8�7	P+m;���� �S�t�PvW���W8J�� �������(R�%U+m�G9�ڔ�G��ݛ�44R��o=�Kх0wr�ZU)J�����J)Uǧ�5!�9�w���I[j�;��)E�U�^��J��IEQ%��E" *�>��@7�ޟ*T���X�}�(�M>�:�Wzz�f��)m�y��m5()Xy�#U)J��>���҂Bؗό�j���t������B�
^��>|t}hyB��BhdJU���R��q�v�H��S�t��*��{Y��PC�7�=**T�{y�T�Es�y��ATz��y�5Uѣ=�T�K�����PW��4{���P)g�*%@*�J�TU)J6���E$ yx}U@�Kp���T�+ݭ�*�B�rwUR�Sf̈cZ�����]�UD�]�r�R
�����Oa����Z�TlQ�M�nUJ�+�p�"�YC�jUK��I( ��@�T&�n�%T�%�6uJ��3k�9ҡE
\�wU�J	�uU ��3�(�p�N��;����(�TH%P�D�UW��)( 7=����r��n۵ a��*�l� �� ��p �!�@;�ݗ �. ��(QI+�UT�Io>�I@ ��| wl�P 9���D��l��� �` ���[�غ�� ��r� 2Q)͔�$"J�y� ���., t  A�� n쵎 �`1� ���@t�\ 9��P s��ITR
�(UU��ϩT�n���t�p�p
1�� +�}�����R�0 OY�P�`9 9�8t�<�  � T� Z�* ��d�*Q�)���	���O�bT�J @  hh �� ���� �  C@ 4�5*U=OM �    '�JDeT�� �@�Tڐ�J)�)���A�=F� ƆFD�>����?]~��1�c��9�>���l�^/����y����$�3���	$�D�$$�?��S�I ~��K�������?�����Z���_�����$�>�O�T�bO�ܤD$=o���ù�œ�X�Z�k�b�*b�*b�,�1�b�1S1S1c1cLX�N�1S�������b�*cET�LX�LT�LX�LXȲb�*b�,b�*b�,�S�L^,��Ҧ*b�,b�*b�,b�,�t�����LX�LX�LS1cLYT�LXŌXŌTŌTŌWK1c8������,�I�I1S���b�*b�,b�:S1c1Rb�1S1qd�������b�)�U1c1LXŌS1LTœ����qS1c1S1Su�Ҧ*b�*b�*b�*b�,������&)������S1c1LXŌSLT�������������%Y�qS1SŌXŌZ�������$�LX�LZ��b�)�b�1bb�œ:XŌX�LX�LSŘ���,b�,b�)���b�W1c1LY&,b�1���b�)����*b��*b��b�)���&,�&*b�,b�*b�)���������S1c�LTŌTŌTŌY1c1c�b�J�1cLXŌTŌY8�:Xœ1dŌT�LT�Ŋ�����&,b�,b�,bɊ�����S1dŌT�LT�LTŌTœ���*b�*b�,b�,bɊdY&,b�,�����,b�*�ŌTŌTŌY1S1St�T�N,���&,bɋ���J�������&,bɊ��dœ1S1S1SLXŌ^,��t��&,bɊ�f*b��LT�L^���qdŌY1S1SLTŌZ�Tœ1d�LTœ1S:\Y1S����&*b�*b�,b���:TŌT��*b�,b�*bɋ'�*b���b�)�����N�1c1S1S1S1j�,�I�����LS�J�*b�,b�*b�*b��X��LXŌSŌS1S���*qLS1c1X���LXŌS�1d��,�S&,�1Rb�1cœI��)�b�)����LS�LXŒb�)���1d���b�)�$œUI�b�,�1LX�qc8��b�,b��,b�,��J���b��LT�N�b�1N)�$�1LV,�b�,b�)��,b�-X�LX�1dŌS1SU�������*b�d��*b��,b�,cETŌYұc8�����c1c1cLXŌX�1ӨŌX��,b���1c1c1c1SLYV1c1S1S1S1SұS�,b�)�b�U�b�1LS1LT��,�&,b���$��c1bqI��T����"b�`b�#���H�Db�1d���ŒF,��$b�#���X�F(�PbĒb�I�I���IY1Q,��C$bČY!���$b�1Db�1Bb��bF*$b�1RF*H�	���DbȌTF)#�#AҤ1a�Pb��$b�1Db�1bF*#u1d�ҡ1R��X&,�1d��$�b�1Bb�J��Hő�#$b�1Bb��T��1Q�#$b�1I�*D�$t��T���I�#Db�#I�1`��#�Œb�:Y$bČY$b�Y$b�1H��LP��#I��XF)�1D�,��Hb�1bF*#�H���Y"b���e��X�,��LY,��Hb�LUX�LS1S1cLS1cqdŎ�ŌXœ1gK&,b�1S��X�N,b�,b���b�,�V,t�LX�1LXŌY&,b�,bΖ1S��*b���$Œb�ұRb�S&,�I���LX�qd�:T�1c1LS�LV*�b���b�,b���b�)�$�1d�ŌS�LS1LT�U�1c�LXŌY&,b��t��)�1LTŌT�1S8�Q��)�����,��c1LTŌTŌWK1LX��*b�*b�)���,����,b�,��*b�1S�u,b�,b�)������S1c1c1S1S�LX�b��������*bɊ���(#[��UDB�����q�;����m�p�`�Oj�{e:�u;�H;&m���ԓ����a�,�ZY4O*����u� �� =�������n����Z�7T2�T�P4wGe��m��̭��u��V�|�2��ؾɹwذ����س'�  ��P"&�ܮ�O�h������k��;G���������/��2n��$��xč28${����+�Ћo8�9Ų��m���1��=LO�]�4*Q�_\�jݴ��$��4!���!���c�hG^�ִ
� �vf��=�_g�I%��2����Y�$!K��tn�}��F�vb$���74(,�a��m�#��Cz���|H�՝4Z�ؠsl=����Ǣ��*y��K�����)YSg�+tm:�/����ź���χ�׹�^�<a��*51F���f,ڬ�cZ��̅�5�ȼ�����栖�N`���f���j	�� nǮZ�ܪ1�H:�T�}tkn�q�l-[�������[y�A���z�nk�L�T��X�0�TDW��5[f��*'6V��q{FJ^&���3^ �ǌ⡠�}~�1"�F䘽�C~�%�5,��4j�U�q-7s^h[�V��pY��hHH:Ϝ�{�~�ʗW�r�a�����z�x�V�0�C
l�g�z��/������4�j�љ�<3�N�Q�<�mIaΪ���wzRmGt(�bdH���T1��vbb��q�A1v2�ǫuLb�R��?���3��y�u�3	�l���2k��J�GG�qVAr�)^�&�n�ݪ�k#��A䕸#Á��~e����鹓�aZ�+�� �����8s[�9L>�3�"��bj�-�E���ֽ,z�^>9k�LF�u��2qDfAa�5D�ZAhP"�f�8�۬
�7^%S	`Żr+���*Ƌ�mɷhL�T�^��1L���A��b�Ⲗ&sN?<��B�c�-Ďy�`�<[zdI
��r޺��L:W�ZoH5�nk����VE�b�o���܎��NȾ{�a���^k�}f1��q�.����fb��j��3�%a��!��9
ͤd�R�ir�q��Ō�~�JKsA�R�k����'�u�^QZ��(���jݐE�e���̩��X3(VH\�J��#��$ǰ��s��knf�c�aU�.���N���.�wb�H�ٺ�]e�!��V�\�^�rg��\F&n�zz�d�3|���$����¨B6��n_���,"�T�&��K�F"���J,�^0��k{C��	a�4/7���1���6��,�Fj9u%Yo٘͹�c2<�~��PFy�6��5�y3��y�s�+�X[�虱h�^�d�ܠ8�"G�rEJH����0�6XkjΉ�{�H�U�B��9��9���m���E��k]�<�f��ȟ�ʌ�&f�(.!�a����ou�ef�4����պU^�wHD^���Z�mLH:El{Yơ�)��$�(/S��Bk�{�6�C0$e���$٘q�P���^�{��������L�Z�]AFmX�ncvУ��PC5	ky�ݑ�^�`F�����h`�T�)ԫμ0`��b�x�C|žW�=s@6�l���9��̚>g-��wcD��V��*��uF�ka��0�"�|���m�B��l������y�,�|��U��C���Ǎ�n��JxR������ceE0�+]ֱt��������)׳Xs�'ѕ��Ր		��]�a:�����>�Aw
���+�T
g���v��*y�_1c�۲��hs�j��ڋ=a�[����b���͢Q��sW��8�����I���ؼLW#0
O����xӲ�#�z�ԛՂ�:71���Ml؇���n���������6*�����|��U��]�����sP��\���LY̖�����&7)���#%�D~J"=w&,��b����e�R�@אݤ(�a=��m�b�(&���F���anA���9WEJ����V5%�. ֮k!�><i���2�֥�nQ�LŎB�ʪ^kv��mU�x��Å+ɰ��YD���3i��0$,�K��m�+�EG�r��lމNU�TRV$#�y5#[�#2x�}�"U���:�#�d�2���%Tm.��n"��瘼Q�!��[BM���t2��sK���LN���Jɘ�	�ٹ��)�F�)\��1�����ә+74l�Pǎ��6]�ôj�A��i��F⌶K"��S8wPwz��M�=Kڜ����7|�1ۧn�.��@@c>^���s�+Bњ��=��U�+U�K.D���c��˳�a_Lb�7�#4�4�MV�<�ܙ��^��dkH����[��<��	}v�Ko�2Z�6}~k�|�c�Xn9�֍��8�
�_�Z�]�d(��pmAT-�2�uD<�,ު����^�ׇ�I}��kү�w�D�|��h^�Ѹ!�"��.bx���`ʄ�0��9!~J��6湏��[6e'۾O^Тȴ�z���-w�r����kR7o�<%����݄��{J�D9��� $6���5��:��5��2��۞�g��}�<���'���Y�/g�j
%���2�l�#`Af�U��D�3MU�zUE-��?jۖ+��S�����H�{��+5	�.��a���q���Geһn�S`V�;V���ؙ�+�����摚E��w������A`�^+�P�?,9��j0��l�
�0�d\�0���z,j"ρ�<%�ǋ�]�B�a˩PKN���,zrVP�aف�f�^��<zQ5 �ķ�c����5sb��CcX����e�h���%�U����/fA.[���W��C#�k5��U�3Q�/n���!�{W�swC�jBȽ��V������;�`�s�d>�4M����K��h�>��jȎ�y�I��cCMO��n<?`�fb;)���^��m��j>~�~Z�\u�*����i�եf��VѬ9,��v�0��o[�<�5�T�x��3|��:�%AY��D��L�~JzBj/G��~�v	Q�����	5i�Z=�L���bZ�#�2y�Q`�P<e;>u�b����� �Ed���-��u2���~��scǞ	s0|�ߔV�U��OD'sP8Iա�֞��p�ܗ�4䷢�"F#l��p���мwH^�*����8�Mf�a�~J����@nc/5ff�!���X���<��=�V�Lj�� ��4�ErX,I-m\�]<4�����mi� g�=��-�y�w�C_��P���Tܖ1�e8Sͱ��� �j-,�6�`�&��V�@ɧ����Rۘ2��,n{���ԖkF_�Z��B��*��Q��jC��g���{/kpd9�^�93w���t5���[�5�rn��S*L�Af�LTn
�n��7M1��M�a̡�1R�,��\��K�n+�N���NI~��E<�tbeF�wfE�P��k��LnЛ׫1���ݻY0�'m��y����y���k[�{f�L��q���1h��.ژ�[0�i��jk�Tv���[�qN鹾�%#��l4<Z��i溭���y���a�G�V�j~�
�MӾ��c�\W����]�+IJW���軫��m�t[�vރ��lA��!�/d�����L.H�i���Hv�M���#v��-��������ic.�ak2��-k��q1rc����b�j��f{}�4Ϡ�fKu�߲��&�j�.�h����U��jF�%�5̅R����ɱ
!I{d`V��w0��z���׸|��&
���V&}!��3���ݘ;T�݌44k2�o	kk���On8
�p�l3�	�j�R[u6��Mg]o�ە�.�Ai��{X׮P)���+F^��\��D1�%�ح�/���P<v*|�GA2��}�ض�潠�� o�V��m��@�<���Y��C"����.�Q��ܱW���v.�a�":�%%Xsq�e��UIc��>ѳ�D��l�����P�Ax��h�[Y��)�,�_Ve<�+��<۩�3wt��ٲ�d�j��I�&���,6/D�j�"n{u���.�ՠ��d!{}���[�;���"��l��L�E[��r�.�F��|��L@_F���U�-�Ҕ��o�|2=�sEZ��Vd36�R��cQg�������i0a�zqL�R�D^d��q�7c�L�l�ʂ�l:r_k�3N��
��aur��ɳfct�`tj:it�@ZS%���MG�褞*s�G�꧲�h��Eݖ0ɹ��)�z�i>�<��^�y+H��j��<����w6nJ4���\��]���4:�{��J4�f++[�o��dnR�y���l[�Dý��ChY�0B��o�G�/]��un�T�������b��tl%L���dV�ȉ���6���3\���gu�XY��4�lQ�62^��*mh�*5RW�*�z�kY�+����N�W�`'4�!.��8*�ܶ�TL�Lt˷YR?:��o�?nG�yPηM��S��0b���f�K��r��]�^���.�����1;����(���@H�m�v�0��O��9�j���s^�s]���C��S Bo��d�sb�w��
[^�&�g�rX=�Q�V��&^��$EFI�{Q�51Y��݃=6`:&3]��G�Y��1<�2�3I�����f-���R�v��B������ȄfE
���a����F���ؾ������E*��iZ��XF��,�s 	�}�xV41�byW��,8��u��{U&��k�\���τ��H�����5 �/g��ܽ���#v�;y[,F�W���IV�������X�!���	x�1]�G�Sl
o���N�]?������
ê',�f�Z,R=ݙ����m��.����I�Ҳ��ѳqffke(�kys'�
=�=C	e[礳p�fVՆ��
t71���&^��lt�u�7�@v��>Ym5ǻ�)��&�y(kv8,�-�a���+lGZ�=�nוh��>�Q�Y�jE���"ތGk˷����s	��y���ˣ5]�:�p��{^n�y\�M��W�MĜ�jj�t���KBX�ؖ������`�:BU�w^(Y�Т���,�c��|̭o��%)�UP��=��`���~q�"���Y4�X��r�Uۅ���&�`2�E�����4�Y"(�	[�ӫ ��Э:�Z8s@
�#�^ܞ�m�����5�a�����	�y��G4�0,����Y�u%�=�}��K�B���k2
Uܞ�"	Q�!cH�>4w0l��H��$~Rm��7$Z��H��XZ����I���O���"�Wp{"�Y�iط;��,����m�J5�-5�f��Ī��%�`�`��7_��	ŀ��6H�l���jMR��A�%a�Pn,��A2�Ix1ʆ�3J�M�.�^+��)�H,��ݗ��<����JL���!���\��ъ�x��nC�ć�<���.rjw���$�<��YI��N�4�l��&��-��U��	W�!ĊTEQ+����m�L�C!�e�HD��V�Z'�����9�a�:_�T�|xy	��d�$����j��KI�	��I�%81�hT�NZ���6(%�Z7�p�n��.X��.]�L*X�J%iE�����,��]:��fqf��E)�N����I�0Hr%��Ӧ�n��G��������]���O�4�-&��FbOP6�F�1|��T��e� e)]�$��ar��׸'���,�z$�#Y�%�x�oT�v��2�ӄ4��lv�C�6�ԑ�`�a��:%�����xA�G��JRd��=��w�YR���p�J�)w7�8[�diB.'b0i�<�q�T�P^m�{J!.Cx�6�-�c��UŤ���*c˰lJ�w#��J	"`��%*m�������J��?^��$�+��"y�,�v�_��W�����ܪ��6�-��H~���T�a�hF��*!��"���H��d�J�yU�M-�������T&��F ���23���F#NƺIr;GL��ql#n�����~CƏhGA�4�a0�Jh��,0�K$tڼCői��kI!U�J����Y��������J��nC��X�N�)m�F�iO�G;,�����v���X�M���r�lx8��%cP�0�)�#vT�)���� �nS-0J�F1�m4�AԬ/<��7��]��F��_�,6�J�֘ë	�	s�f0�~K?8�������L9��漃ݣ<�Ms]�?s|q)��C4y�Z�ۙq�!ʇa�^>���klP�ާ{ֆXD�L�T-0�ũ<*��1�6�IY�R�e5�}�ռ�۫�b�&�63:�ZU,��u��G�o�,� �CN�4�bXK$��L�r������dQ�������p�WlB	��\��\��0�Gh���[M�a4̓R�d���n K��쪪6!h�>EI�;�٢g�"
D���lj;y�M��&�$E���wt6�����	�՚HK�$�&<Y��B>u�:�K1`������|K(��Ѷ`�強s���k����	�N)Rno���ng�,�V�G�jQƖ+J�(�G$�	KҒJ��j$�ؚ�G]S!a��m��������s���è� ��6א�{UgYe{EZ�$�<W�3'���tf�[���T��+��| ��Z����P��I1A�Z(�A$RH��I"�d[�i��n�h����'ztgw�{��xs�jW�p��Kɹt��l�R�i)4��*����r�89��V-�)U$�eAz��S6i�wc��G���}�7��@��áz�3��;_�T�����I$�I$�I$�N��r�>����Z�0�g�׬�B�#�oZu�>׋u�-B�iL�`�9ү���.+�#}r�*���8��/e׈�qS*�z�4z;�'v:�WV�3�sשI6������uƚx�̛����ɣE~�僀Sݝ�6�@'*~m�s�Skdq���lZ��3���l��)�6���ag�No%.�`Qŝ��t�O��2��	Ͱ�&��OҎ�~�4p�7߻�Z=r_A�[��1��sÍ�oF}t�9X��	��.��;�sܵ�o;D>�M��6s!�+Xc(U' ��6\�'Dْ�wIy��Gc�]\�ʎ�Ĵ���h�^�z�J�yG�'S�&�%=��Z�g�z�Sܼ�<�g�698��ۙ�\��޼�������1+&U�InY� +#z��՗±��F��rظǆ-�\F�2�C7�4p�fc�k�^�eZ�cjoӱ�{�ݓeU��{���
AK�v�D�<�U�۫#��!�9m��#���_f��ڪg۹����\9�3E�r��ϟ���uk���u�����P��'�Vl �2��;��5�d��Us�)�w<���=qp�i��dx=j/b8��e�4��i��ˋeJ�PG��#�=m's�7��	4]rT�-�冻��u��she��\Ba��R�����j���	��r�2��`y�,�r�*NƣV8��n><Ι�N<W~j�D��g7\��&�/���1�D���b}��Q��V��Fz��Ï�C���y{�c��c���r�K�q�0Նh���;��*�n車����R=b6Ҝz�9?'�c���-�O:�z�,�kh3n���ü^��w�dC������tPϫ�����)�eZ7,%eLf*�3���u�7M��K�h��М+����-8�=r���UY:�߷`<h�m�B�|���k1�L1,Wi���)͜��;�ʮ�M׏ ���!�Ѵǩ��ϧXjɦ��C|��۪���z^��_����4*�ٌb�kY���i��۠�6�N�[jR�o��N;�Ftk�`W��c4��;�\��)Zʭ��Z�]�n}���՚�Iհ��k7��勢�.��uR��ܣ��s3#���p�7����qs��/!��8�{ٳ纻2b��gúx���Yʜb�
[�nl��R������$o
TQ#AƘ��J��Be�r�{IJ'��|����27�v�s�\{�JUL"�F]�	��ڽ�眫s�ޝRfa�^�r�[�vU����|{��1�X�'�y��Z��@��⤌�q�=�Z}J�v�s��k�s�wfJ���/���ky���ރ82�k|�0!���"ĵ��J՝@�2��Y��m��o������x�h��٭n8p�=ٽV��$@���2�ڸ��GMa�8������*�=v��e�`xo�)i_ofy�}�=���.�@ާ��{8�Rc3�z֟
����.��M��6;�+*Qe�=��4��[�Ҋ$�Lx����d^X�r�%�rY�������1j���g�U:Bɷ�+:<�Oe�t:p�wC9�YO73��X�0�އ2���I��=jF�}��r�[4f��*ͼp�v�"9�b=_����Z���
���h���Ռn�W���<��j��?4��9�wؙȅt*�]�}p��Y���,W��̇�䰘��>���+����>f��J���|�䳞w��o��7�ܲ�M�{��=�[�\���-�hģv�z�ss9�-��y��s�3<�\����{�e�����ݙՇ_P��:�uk6��$��m�=;��vVe�r�����xƂ�	�>Z�F������&$^6�C���|!pŶ3�5�ʩ��|����ҝ�Y��sU:�M՝���uP8zK���ػ��`�^:G�'y��MV��0;�z+������l��v3��%�Z�H��=���jeȰ��ze}�'2����wr�%�k={0��)���w��I[=�z���,�{k4�:F�S�!7O�}�=ڞ�n/�s�%���@�
Ww�K�%����9�F��f>��F=>���C�ժ���?,�N�̇�K:�C0[R���N�m%X������5��|,m���b5�+��7�k�v���޹��{�7��
4�j���E�-k
��� ��Y�w����#���g��\X���G\;&4�� �O!���;�Mιٺ��L��a;���m.M�S�&�}M[�
�ֈlۊ�� ���8�^仼� 6x�������?�>J�K�j%�v��4��x=:��ͽ�x����6؏��,�ï8�v�?g�r^X��?�����9�7�q�g�ԒۤD7��g�a�%kT���7O.����=��x��o��5A�)��n�2(�SӖ9G����eI~3�[]!n��'��z�2��粞��/Y��>�s�kడq׻z���#�`�!�=f�y��M!v=1��l����s7��d�6�k�Gok�;H���X��ň�>Z3��ݞ5�=���R-��t���*�b�ޥD�8�xT�˲����ׇ�os�5����Gj�;���Q-�Nr%N;(d���g8�&��;��ܮ��"��j�Q�v����K�m�Q���)�m�2��J�V�����gR��i�_�]�Qʡ�rJ5�{^�n7R�n���9�_�1A�W}��n����%fɌ��o
�=s�Ӑ�z�	�T�^�?&S���uKܽӱ/.�������O����ѵ�x��0�g'����||=wo3�on��[�$��q���pL��wSS�Xu�w{k�\�r���SK���G�`�{�h������z�k|9���6�q����c咮���&��a�2I"^�(�WY�qgr�;�wf�V}�gW���NޞFu�Wɇ�#iz�>3�œ�wVX�\s<	yԁ��AeH�~�� �=�t/3�f�	X0)�����:޼�^�}U#6�gL�s2U��38C�}�l�ǖ��xo3]Zܴ�^���X�>��vη,��,�6gs�G�i��v�",~�����Y��$����8V��9�Y�h**u0�E�);)*]Y������M��ܻ����yˀ�%��d:!�r�g[�׍PO��[E�6�^̭�b徘��GR���Z0nN��ٙ��`�'f���]��"�9Х���Q�_'��3V* 0 ��2����-z41TX�L�q��9�M>? �S ���y!45��V^+��&.�n�R�b-��}�D�q�5's6n�3��L<�7�;�Y���G
)���r�y;
0K޼ �3l]�Yw0+JEq���*��pE����X���qo��lfj�Jc�%l�'W����CWΕV�W9'��pS��^�n�#���,U��uUn��9y�h@��IT�wNV�Q��B�	��qh���(c������d:g�-JG���c�M;XVUU�7sp<ߐ>́�B� I3�i�u���28	٘�c_�J�X��i�Jy��u*�U��r��	��!�]�y�:Q�+VxD �Ǖ����`�cQ���/6���%�;�����ZW�ˬWE+��{�7�oSsN�p��_ bkrx툣&��Ywo��++������=}�k������ä��}h�J��YW�GfaW�dw�.UNN���ɇ�/�n�$Z��4��,�AK4.����i�-��Zާ�ڜ@uq�=�J�Ȗ�S�����~�&� ���Z�&Q��L�绬*��m�Z�w����ہ���h*\�$�J�v�2��'G�O^%��'��[���jM닄�O$��z�c+
�����B��:7�/H�*�����gK������uu�g\WǸ�ѽft��e��O�"P�p�B���\JyrQ�}3=h�,��2	\y�Bb��+���Z���Bs�0�\��ڐ�j�:�=�1��>]���gTP�FE��̣�a�O_nҞ�˚ߋ׌@�X�9�ۼ|�]Rﻜ��<%���[;j=�-�ݭ���|WN�!�Ŏ��#}]�	3M����K�Q�7]��Kj>�"Uþ��R�m� �v���8��$�m�A��t<���c��M�������{���\#�4㩒��e��]]�䦖�5�y�Av��@���y3�p�XTC�6+v������i"��Q���xxB�%g^���U���}\�ީz�u��&m9f������'=+"�}^ ���;c$�3g5��1z�9�,��Csݸ���2�LWӮ.9��6�(�8�B��mLW�g���6<��xh��;Ԣ��oo��=T�u^�pܪ��w�r̹t%�'E<��gdY�PBNf���� ���ɼ��Gl��;�����y�c㸃�n�Uf7�wt���*�s$v5�`�����g�sıM����H)h}1:�\���R~n��c���6��ƶ�Z��v����dL=��D�D�u�V����c�;��o�B	��m�LA��h���L7
vú�Y�����Q�9s_�N�ݺ<]�q�пf��>i�n<嘬>�+�Ws��&;%�)g�;���+�M�i|�#ۯW�O[:f�ކ��D�xw-�X츺@|��s��u�ʋ������P=�tݝ���ҡ��rU���\���s�2�_Q�a ?N�O,�.ı?^��}�:
�%�vq��k5L��:�>���z3voIw7x=��ʹ0��^���&�X�Abvm�U:�4���&�G�K/�3^!�x��VwG���ԭCbU���k˳�0���f��bO�BrDu."�ޡީ���M���9�M�mVU��^��6�&���iq�)�b+�j�܏��=Ϧ��lOQ���A�v�w�uL�(�,�J�#�,�O��4{���������퐼�P�v��6�o��w�ZiQ�\�w*���P�(��y�i��E�_x��®h����B���[��DoSF��/xx��U��b�é� NgԺ[c�=Б����yp���I${�[�}��:���4e����k}��o���2��S_*p[6�O]���_��'�U�����[�,����Y[CvR�OU��A��s�_p��y�_���aGË���*��p�-�ff�Ĳf�gE�ZiI=z��0������3(.��v��4Hi��v;���S�Նt�^cޮ_4vұ���S1��K�f�n݋M`z�����؎���}� ��)�'\�N.�զ�U�7�	Y*�J*�������v���]fr�6�G��P/�w�Ԉt(y�*+�ﷆ*�3����9ÁI��r�����z�&˪}y�(wlǷ]��n���c�/9�OPR-m�B��y���x{�.f�łN����M�sM\��j���;�eX^m��زxr�G{�.�`�r��ì$.��_�ME�v��{�wq~�>�򋷦ի�w���.���S����p���������k���	�䉸
�@�l)��#HY�H0�R$�A���e4��CA�a��,�͘h�I8Ds4��M���b,R�$�$Ha���AZ%���:Dc��nLjB
����D9��6�nԑA�)�����*�h��e"���E;�|w��c@�d��c����Z���(A)h�X�-�˳��I�	2�I"�f�И�U�� K�	H�N�}6S�X�ā4 d}.\��J$�	m|��.�R8AJw��!��/R��P���b'���4T4��l��k��<iH&I�#�c#����l�&�L	2�=�p��P�d�
 �bNEZR6�ƭĩ%[ѝ��Hq�ˁ��a���.HIED8��(�a��D��0�:Ÿ۶t�7 ��<�l�1�+.m���#�9�ĵ�����N�rQQ�j"d��q�ˁµ�v�J�T�CP��)���l�a�\����#���� �	c��Ѧ3	�����(�M��#��SVH���a1"��N��l��P�K�w��k�G")M�q��*Q$�D@V��H�
��Ё����gF�ց*�%#��,�7#-�E��DL���H�ل���W����JJFZ*]��C�Y��h8�N�#����0^�*6�m&��#	#v&Lͺ�Ki��(�*�2��+��7��SI�&5!IPMx�뭐�u�(�#r�	&$0��S,��2�`p㵖2��S8Y�$���.ɰ�)�$��w,B̐2`-ơ��V�¸��J[�&���՝Aش�n�J|�j��v�	)���d�M��tK�]HC�Rl�\��Me�>�RAca�Xf�&$b8�e"3�"�U@_����o�$I"'�������O�>�	$#_��������R��1�I��6��Ip����y�fY�����+����/��Z�������%ܑ7���cG��Ī��}�ﯺ4J{�^��I�<�4�2-I���{��C�5�����[6N1l��`­m�;قw>w�j2����7��`��L�.<��%t�x��obpz{|g�{�/%�]�|B�g���RVTs��?,�M=Ǹ���ǘ��9�/v{�7�ʅ����>ֶm1d��Mr�eShV[�}���t�ܦpU��L��}kx�ȇ5�z=�M����^�IGei:��&/Nni��������
�#�D��h,v�RaU�e(���]��Ș1wB�f��t��exW=s��vZ/��  �m����ݺBE=oUc�{"�� ��K���hd�AJm�������8��|<uk�ε��p�̫���g	��ww"�%������z���;^�`�x�-��Hh�A=5�p�'c�&�e�I��r�Oˬ��_h��]���LP�t�'��)8��U�����X���H��f�j[�b�3{����Kk�i]kٛ3��#�w����f��������zv�Ƕ�5�lkZֵ�k[ֵ�kZ��kZֵ�{k]5�kZ�kXֵ�Zֵ�{kZ��ֵ�MkZ�Zֵ�Mk]5�kZ׶��q�kZצ���ֵ�k�Z�kZֵ�j��kZ�kXֵ�5�kZ�֫Zֵ�k�cZ�On8ֱ�kZֽ5�q�kZֵ��V��kZֵ��Mk\kZֶ5�kZֵ��kZֵ�kcZֵ�k^�_Ef�t%Z̹6_��z]�H�s����5k;s�2;�����b�y3��-.�cˣ����)��U޳��M�D+��j��﫳^�ؽ1Y�Wym܁Zu� ��D,5���l�����i�@�������q-K���p%�eᬋw����ç<�Ӌ3�����<�J�S���na]��\O�;0k�&��G�Q��SF��?�Ů���b�N*]�ݒ�%[�daي��#��ҋ1q9~b���]޻��6Rڔ�{z�7y�d�I�fT�z^�� \ƠL;���/9$o��}v��e���ye?/GٙC�V0�f�ê�f�:dфdv
�!bޝҟM�ns�h�'�Hs�bH×7�q��;�� O��HZ�}W�Ld�)��k�Hʩu�rq�|�s;{��.��H��w-��8Sqh�,�
'�b�i�L�I�5TD����خ�p���ꤼ]�0��|��I�1<�؃�X�1�-�v�XR��h]�nNv��y�qAVFr���U�sB���������\��1ou�����gs&=2����k�~�\j���(����z �ˠ��/��n��־5�ֵ�kZ�֫Zֵ�k�cZֵ�kZ�ֵ�k^�ֵָ�cZֵ�Zֵ��ֵ�kZֻkZ�5�kZ�k^ݵ�5�vֵ�kZֵ�Zֱ�k\kZֵ鱭kZֵ�tֵ�cZֵ�Zֵָ�k�cZ�N�5�ֵ�kZֶ5�kZֵ�k]5�kZ׶���ֵ�k�Z�kZֵ��j��k���|kU�kZ֕�`uAY	�+'k�����X�y���K�s�ֲ���;.X�7�{7�P*1���|�z-�J4Ob"�ۼ���}�i�ZƇ�����UaQ���ޝ�X��B�k�uYz�_����Or���p*�_�y�&bז���q��oMZ����+�|/w�Բ8w�xm�m��w�toxl6�P�L��<:�;�C�A�,�g<p#(��1�<0�5���oK��IޏS�\ɑ�8Ǘ#��n�>�&���ЇB��/2�p�{\�i����y����>�H���'���3|/'��{U�-��j��w�����ZnA��u��x�3�����[G�k5�2��w�����|!�t>}�F~e�Îc+����>��3R�_MvT8��5q���!	��+�#�Hhc�����ݦ�H�Y��J��ST����#�,�ح.��g��{wZFo*��w:���gi#o�.~*���Nɲ�vj�-D��3����Q�(tX2�ر�ny�2`�%T�gl =�v{���5Gk2a���8�y���֟'��-�#	��1��SE螿g������kZ�kXֵ�vֵ�5�kZ�ֵ�Zֵ�{kU�kZֵ�V��kZ׶��Zֵ�k�Z�kZֵ��V��kZ׶��Zֵ�k_�kZֵ�k�k]5�q�kX֫Zֵ�kZ�kZֵ�k�kZ�5�k]��t�tֶ5�kZֵ�k]5�kZ׶��kֵ��ֵ�kZֻkZ�ֵ�zkZ�ֵ�zkZ�ֵ�{���]�B,wFl�t�Zr�X�Ӫ�4���z㽺
�������]E�݉`H`B�Yu��	���{���;��>�>W���I�̵,q�yY�6��.=Ti#(�N�9̝�.��n�'{8S�^�7��Q�9�;ȋ��J:�ݖ�=�ZģɌo��[�sUS�F��%r7�T�.�s���ڶGxw0�ɢ�`��]�e9S���A�GU���P��L}��w4]����gF�[��!d�����-��Hc93�R�Ԙ �O��FW@� V�f�5<��e��ǅ��:�\O&yt�;����k��g���{�����h�����˽�q幏�AU5N2����������Q��`�]LV7K�kVt�A{�4(�P��*';#a��t������w�2�1��CT�lR��K��^E`jFkH#\n��ܦ-�z뭢�!JaK�=�׻��C˫�x郬Ǫ�q\ķ�d�G��}�AP�p�`�I'�C�	�
��w�>�G�4ط���j�y�C��%��=�������F%;�x���)��c���6�JԺ�ٱ;�Ԓ����:�OX�n����ֵƵ�kZ�ֵƵ�k]��kֵ�kZֻkXֱ�k�Z�֫Zֵ�k�cZֵ�kZ�ֵ�kZֶ5�kZֵ��kZֵ�kcZֵ�kZ�ֵ�k^�ֵָ�5�kZ�֫Zֵ��kU�kZֵ�tֵ�8�kZֵָ�k�Zֵ��ֵ�kZֵ�k�kZֵ�mk���kZ׶��Zֵ�k�Z�kZ֯���z�� ����v��0��'�wdD�^��۷���*�(���+�EM�.^�P%/G�-Q~!}���|c���Iӱ�63*��/f6�3mS���<��*���O��I閈�3Q|��#�}Dդ�ߎ��m>͙�4����g���I�����Uׇ�y��w*e���ק5e�
��ѻG�Uv_'Ns�|��Sx���l����cg���B���ۋ��ֲI-����uL[������_��Oӫ��3׳`c��˨��3��}��36��X�ԃi�y�K�X��Dlp��W�uʰ��3��Y��c@ Q�]��]7 ��1�Uݶ�ͮe:Q�U/3�[�&���Q����[z�a*�FxxV^dj,޻l��	E��3�R�p#P	g��F��7�dB�:M2���U�S\��r�ACeAE&| ��y�+������oJ�9od4č����u@��5-�95��:+����}�����V\���S\�L���-� "-u�*��_MF�6!+��Ŗ����7�v@����ڕ�CN�Ը�[{[p�������S�Q�&G��A.q�9
$V�w$M�������uŤku�������j sn�F�f�xo��'}�N���Au�E�iQ&��ME���ʬ���������}�Z�S_q�'^��9�|`#�m�����r�+�����9K19�tWM�(�0/�s�G}�嵳=����|Ġ~5��(w�0,�9�F�6�U.�����[���#^������ˬ8v��s���
��c�؍���sJ�S�:e�z;�ԇ�P�,s�/&V��U�*C��]򔉛f�'W��D��9oRb�����x��Ecs�̍#��,��'h�x�k�8�S���'[��\��r�N�Au�9@e����:�pkMD�&f�<ڙ��$sGX��Cm.�z���8$�`{�Qb��&����lGT��֐a�gZ{U����#Ԇ9ڈ�����fDv�|�b����k�sr\=f];�Uɺ��i{�vGG.VfP�Pv+�6:.b�NT���T�*ô�!}�w(W���l����x�!�����fg_J�ڴ����������ͻ
�xʈ��=�et���D�U�֥9h��� Gt�ga��e�������֯�k!%Y��I����ޗ�F�eCU�����0Wp�fV��2���5�E�޾����i�:�4T�<)�w���܆E&���Q����pɗD��	��d^n�Oy{5���e�Y4op�_G�-WW����"Z���wS.x�J;��?c'�m�<��tUKYhu�*�u����+��]鼐l���.̢2}�$�7����U!�D��-�e��]+صs�	�ΰ0;��s���]�=`�y�v�q�L�p����J[�+���_:�� s��[�!�|�)�r���3��#z���/�/}�6�U�
;���]Ӥ�v�\�L��"R���<�{�zsM��{u�غ ��U�1��u�Z�%\z]\�Gv��p���6[,V�D�{N��jC�Y���/�����Q����PnJ�7��17�sYr��E�Uܠ�brK����*Y��Ja���6A�q	Y�tw{�l��b�ȌK�g��4ԗ�}�N�³�校<7�m�Xڞǲ1c)gXP��θ�c�uuNuG{T�]y��;gv0K��z_:�ܥ��+;�m�[b����l /���b��ȝ���6�Ʀ�)]Q�}zEd��7P;=������V�Ⱖ2e��P� ���r�i�U�|�=C�\�|�E�a�勱���ۈW[	�b���u�c���X���!U����+�����G��*x�l��~���'�ua��y�겗�w���-�Rݘf�Rc����	-�Ϭ9զ���[���CP�ӷ4���xB��2%
���<����|;g�<�Jv��W����D�E�2�#��w��+�δ�T7�t
R���,"Ѽ��,Úp�B)���0{��V��T��m#��[��fX��q���q��v+zڠ��NU;����u���7ؒ�����	.��Z��=��Q�;V�@>��~��>�,��6���S�j�t?^^̔o-=q���/g���)\�+'I��u	�C���o�maIf��ں92]�VPB��9繆�ܹ����a�sw�����=^�y{E��@/"�5Vm�8�/���:*�b���sF:���Nsfæ�b$�����s�-.n�-hʚ�."v-�"���Ղo%ۇDy����/A��*����vUv��<w�co�n������-��i��Y��Vxk��^�q�c���*��i���`���E�#u�����sogD��U�Z��S�Ҷ�R����
��ݻZ"�Q!f�8̲*\���5�]�ΟN�߱A��
cv�M:�Y��̣�q�J"�#۠��dt�o2X��6�v	�Ҽk�Y3���&��#�%k���k� �ƐR�[��K��i���>��#�5�춫��G�r�~S�/M���Q��޲^�u�]b�μ���6T����V�(m6@זvo,]�/<S�o��x�Ǿ@��=y�^K�����⏚�����1��f�L]�f6��~�?b�S���9���_]E��eֳp�N�j]@�:��x̇�c�;q����Ү���ҽ���G��vަ���盋l�V�/��Y�x<�D�Xtа����Q�vj�Ac���wW7���V3��Q�Qf������C���_�٘�R�d�C�#{�.�yY�|���9��n�YWTI�L�;��K��cɽ҄�WV��Ø��fx`�2�K��0�>�Ux`�W jO�^�*~�e��3ܪ�*���`#�'	]�r	�50ۓ3�^~=��>��B�yqY��Q��5u�
L]Vܕ��HK���x��	��,֛o���<Lr�5C�a,���%�f�`�{���U�Ļi�o8�:q�ӽ��M�=>���Y�v��FEb��q�ܼ.�K�4VG���%Sع�/ �U�w_gW�3�'ό��gN�;
x=Ć��Tj+U	��k3B�nK��ڔ1�}�oi�wf���ݝ͎&ķq�y�T��p���,˭9w۶�&��`)�Z�3(l���i��9�Yx3��ͥ�J���!L5U��!G�Z;�f-��ݖ����yz��Lؔ��;�2l��
T��p�^��}��<���.�E+҆oP�6����o�߻�]x�U��+��g����wU�G�gT$�}PP���nv�d��J�F���P֞�v�fVRG�2���}�+}č�k,t[���گ�����US�&����l�}��{��<�7JX�;)�g�Ue������CUD�k�_p�he�nT�7n��U�J�b �:�8\����W�;Fi�����b�����*��Vx�w=�ײ���[��S��{�኎�M��ƹn���Ƥ�z�d��s�2�]���0x{��%��gcW�����	G�5Q�2byi2.��7��� �a���;}�6�h������o$H�7=��������	.w~%m<PV�D����]�O'��ƌ���a��+�=Y&��mIG�+v���==�4�բ�
��w���$��l����?���g�3�?�����������xr�iƓl��&��a�Xh$mJi�FAc0�6���$����Y�@4�3ªԸm��a��4�mB��2�eF�&�	%;�ܿW����w����i�[cp6; � ɤ���Oѹ\��Op��9��hp�VxJ���G=�����1p��q��+A�
��V���9;�8�]�9;7���
)Ƒ��y!7@��;h)vo�|�qHZ�nў�듣&�غ�y�p��O�Վ>K
�����(߆�}fG�{������Ҫ�f�����v��GA���$���S��]�L����\2`�=���tԭf[�m�U��Zt�37��"�g��z�ռ�m6i����
y��E�q\B����r��m��\��8��v�ⷦ�բ��LbއOc�8��r�l�,3���]�0S��{t�{���2��-�LC~�g�V�l���0nf���>�8�c�`��W!tc�@�r�E��r3�˶��-�R��647���xr��i2��F篐G�w��.���q�M��N�u��Z�(���}��8�˃1��oUՍ;�������rY�g���J����s�[;���sk�31]�+u�s��<z[ωr�޴I{p����y��d�Y��I�!��A5,6{#TI0ZI�!�\�KWp��0�D(4�	�S@�*�;����F̓/�L�mă7eSVi�I)�N�P��MD�p�MP$��L(-�RJa�L�p�����0# a�"a@�r1��+�@˶\��$�S���q�W��v�$ȑjG�-��h�@��[ghU���h�z���z�[Km|�t��Ƶ��kZ�nݻv�{��:r���[s_��k_����[P�S#��c_�ֶ5�kZ�۷nݵ�(��R�[,�oVNX�oR%��WW��N1�kZ�Ƶ�k]�v�۶����&Ԝ�[!gVU��-6�~�G���|߻�~�׏�ֵ�k�nݻvּ��ɷ�Z�Eژ,�un��[Z�mgv��I���	m�"[]�NtF��5`�Eks���[R���ۖ���E����wu���u�m��ҬY"J�ݹ��2I��l�2-�@Kk��-F��ݸ~�^���-�^v"�O�[u�s�����\z��m��y�x�󶞝���̷�M.Wn����򧩚�bRQ2� Q���h�H�E�𮻣]�^�����,Y�����5�ݮ���V���ﾾ5F�[�����(�mr7�|���*�$�K�'ȍ]r�
� gKj�_V�nxAu&{J�U�g>EZ}�������f!k-Piĕ//9�7��q!ׅ�xs�rٜ�Q��u墼�8q4>U*�0�\5ܳTIi�J�F� B��9�;��חD��~�����q�E͜���,^]Jkr�l���l�%���.�3R�#q;�ea�mdDe�G�1�D%����Ӑ����%f�niU�l!az�\a�*�6�E]����CcvQE �(���:7��0�I�wF��m�;�x-�ٹ��� N�tv�#U�j�Xf�Nt�5j���f�$��ϱ�q[����~XQ��a�s��kȔ��ɻX	qk����5��k�I�;c�����	�|-���-����Ȕ�:5��9��$��	D-Cc*�_�)�ٮ����i4)Y4sqY�"����ҟ�UV���a/��?��	J̈���5(3�IU^���fg�P
�Z�E숅{>�ĕ,&���!u��H=�|�� 0��n��7|�@�h$q;�Ҧ�2���ѯC��C���I��p�����5�"c�#K������7]Ef�Њz��E��*�p�۔vS�ã7,����ML=�ܾ9�&ny"+� }��M;�<��r��J��!~�N�o�;L)�����_��⪪*���ߝ�����6{����A�F����%J{�T>�蹁}��j�Ln���Gf5,{��2�cu�Y�\F��{vp�{a�ѡ���(��D�ŇS�Hl@����Z��C�l:��Fz� �xp�/D�7�`��;�ww���Sײ�u�-��>��!;}��p׌�9{�&�5֣��h���y���-�����M����l�y}��1���S�:��̶�����L����5y�A�
~���Xs����K�J��}�^�nk0�"��B���A��>��Oub)��,,U�/��O�G��Y�eY[�R��F�s���E[8�o3y�sN�l��O�*_}�y/_Z�M��'����T���}�ۧS���$^��d>�c�D��r|�p�o���L\o��:�I3� �i �Ow���hޱ�3�c��mf�{Xt��t1����t&WB.%@��i���I=�:1��GhA���	����c*��~n��E�\/{"G�OZ�;�j;�Y��3�Yw��:Vwܯ�[ʻ^��!���7�V%���������v�N�ѣF��D�Ι}����X�$�/���>�I�W^E)�Qe�G�aֆ�ld*��Yok��C�ޫ������������iD���a�����oeZ)�]��e��Pv�T�p1h�FC��bL����R��\�w����ٛ���EϘ85���1S��y"��5�)6i˔���r�uf�H��8y ��_;��������6���q^C�>8~#�,��mɼ��IYѸ��V,�|��$�4`��q�CVg��/+�	أl6�[+T���13����۟X��Y����`6��6������/.wdu��xZ�T����H�3:������]���5j����
�Y�8�6 �p�H��F	I/��s�ZRg/�&.������ �f�VV�ǩԍ�q`��=V+g��O}p����g��s�0,渫���9U��;ۘ������W|����q%Q�n��ŕ��s�NW�����צ�+�Y���>Q=ю����q\��sg�ǵveLf���o?[�on�]�n�s��{�}˫��4h�@� u�v�:g�d��ou�8���)�~����m}liK���/r�0����kgԶK����9��<SW�U�v�U�בwח��m��U�k��<>���aaU��d�K�x���U^|�˧��{�v�լЩ;��e�5(�+ׂ�J`��f�M��"o�7
�`����k4飴����m�,c����53҄w;��u�����G]e�A���v}{!V���s"h��m������FC�%��J�%J7+f�U�\a�i3�5��ͩYk&���.|�!��	u�Z�"
��g����Q�[���h	9`�<������5��{��N>�`�֣�)Q�6,e�՛�Tf	xhw}O~KR�;9��7�4p��Fi���B:������q~Z�n���j35�Ms���x�N�S�9�u��B��_I�3�I�^iU�n/�l�c�v1����CU�ť�4딞&׊m=�ű�>މ6$�$�u'���QmQ'`�Qx�M%%S��:#-xէ�{��-�����\���kZn	 �66Q]F�U�2���W�(��1�|���fN[��=�o>eP0pq�G������{尸�ܽ�5G<s�E�J	�I��M�!�!,�I��lpȂ�@�i�"g�@4hѣF�(!D��f���e%�q"o�~ayh����⪲�TP�D��:Y��vM�Sz��Y��sO�ظ,q�P>Q����]��+�2�N�Ё�kEL��#oU=�,G�1�ioH���D��3�" �-I7�S�����uWۜ�6r�cg�'r�T�1�ƹ�c��>cj*�*\>�6m]Li�B}+'U��c��M��8��݆\���L����e���6����X}�;�m{��gku���Nѫ�v�LT�9���I��#m�����爟U�P��dQFNg�7���[�nf\IA�e�K\
���G'%T`�:�ll��q;L �3�����0����2�k	ho<n;�mV�RKNͿ@���:W��r�~@sD��n\�[��v�N�)�j�Hm���l�a��>]6k��ov�+_�|��1j`m��#1��2���Ռ��l_!�8%�(K�L�ʹ�U�+"��|�n6�c�"��z]��L�/�V"�{�\�w��"�9~��<�}Υ���/���_g���ۉм��߻�%Y*�s�|�����ߝz��|���� 3�%���7�N�l�7�N[ƾ�㪴�0r�m��C:��jEk&��x�-�lH`�&����4ffV��0������]P*XN܈��*�Pn 
�I����
��� �^
؛V�(��WFO�>�iƨqu����=�t"��6m�2�PUUBӰ7jk
� >g���!w�^Ѐ��R R�j8V���_o!�$F��^�cw��Q��a�Q	{��ݧh�Z@Ù��Q��MBi
uE�>�Ob�����}�0-��ݨd�ŗ.��z�f��'E���DMI�a0�eǒ���@�O�%�:�ҕ��݂N��T$&!X���zQ��7d��Յ]FR ���IQ�7Oj��y���D�b�X9��ʳSL��2�m�[-k1�Xۋ�&������{�Ǒ�2\����B�.[��-Vl�5��Õh���'�V��جL��ܫhڊ�Ĳ�Z�M2a��8_���^�.�����Z{���|�����Z��mu��<gc�<:��S������[\�h�hѣUC�g5���f�#�u��M�v10�>�Um[��eF7#ib�:&mi�aoL�&�FQ����3V��9^�!�cԱ�!��9W�
'H6wr��'M�I)��l
u���U1[����rr2�p�a9nD�N�����Y�J4�9�|�{�T�Y6 �ҡ��6m�7#,H��"$4��2S�<|.F:�*�py�Z�̶ʰ�6�B�ޯs5w�Kh��nH�wY>�oFO�O�݃,��J,��]-���sU^I�$[3��g�;e4��d��Ȉ�d=읖�)��F����Pﷹ�A��I/h�1�8!}��6�΁S0\�Q;��+_\k'm��3pJ�C��N��H�+rV1��>�B քv�
�t�g5]�ɳ6���2=J�,����ہqϠ+��K�u�֔��}���sR�ü�(�8A�����L�t����s}��ڝ���q��9E��>x.���g��?[Oz[�W�fu{N^�����~r��}8�*�w/���L�vwQ����t>�wz��VJ�U#���{�����=]��o~w�iX������ Hq��և۳7�&4c���Ԧn��8�������6���/��;�u?���ShL�0i��#v�6��,�1R�@�-2� ��׬mE�?`����I��ɛ$
�1�a�^^��lFh���4VJ�m��,�M5�v�>~��>aTl)~�l��:��WuVF��,j�
t�i;QQ.pR
�����V�-jX���f�hf��nf���ew9�ۙ��Y�4�}��{;��w
[[ԃ�E?��&��s%�	(�|�����'Z�I�j�W�&o}�G)�l Q&��E����-��Dl,ġ�"&r�P��mEঊA����/W�6`:��*�ب�� q�-�u5y��
�fb��/���YEϮ�#!�#�ƶDl��j%�1�I���MF��`?n�I'�^|�s�����)I�=39��W�YߍE<��3C�b��B�h�J�`�*Sn�3�ad�ј�㓆���!��|F{�������t��1ys�#��+2qݾWVn�<�I�B��,0!*�	�!�%�ѣF��R8��|�9��v�&D41`����ۢ�$�I�����^�Dߛ=����B��-�Ù,����x�Q�{3�w@7��N+@[�g�y��ת�vY��<z6���Lꅑ��M�Ȝ�J>L�ҍõ^�۟nm������֪�f��|9Y�QE*D�RrTc�3+��}���W�h?��E��K>��;�� ����J�v�j��&q���od��Yb�J1��4a��ǻ����wd�5FnX�햯"�/��P�m�׊+#��A���W��5��R�\ig���t�C��X6il��^�mW��Ͼد��ǯ%��)(���'�^�y"p�YG^_؃@�.aο��F��])��ݳ��Y(h���<w)u���13E=|=��q�XG��W��Iy������rC��;�J����?���5[[����?$�V�2E%{_���P����б�EE��w�3��}�U�gi��B��z*A=����W+���b}�G��� |I��C�o���%�7�>�����2���\:�|zL��\�cԨn?Is,�S:�h����� ѣDDP���w�}ݏ~�iݚ+F����o�;�Q���Qٺ牸O�5�q�YB;uV�f������P�cL�?��S�*v/gҲQN^MbwJֹ:�@�	%-���Q���\/���ε�v�
���c9�:�i��A+�H�&A3��#j��R�v������2�v�xa'T�Zj�p����C�5��H�c�p�:W�Ta��-���8�l����VA9v�9�kwڽK�x0�g�v+�kPNb
�EBk�x�љ]�Z������CL�#B�YT
U��¸�K�Q�!C���$ML3ө��f�N���5�⚝ɟG������C�f�/��FL|���>�u�*w���L�{D����Fg!|�oO������X�f^�Ť�9	�cP3�;���!��w�D�<��z�@�d3�v} �D������}�_jj~�_�fHxn�Q��ǝ��^�JZ�y[*�vc���:�N�'y�PVWK��Y4^��_����ս�/c��'��ڳ}W�f%^g!s���$zv%��n����{:h�h^���y�yp�VA�yv;���Ý�ʲi��v���.xw++p�1�N_a�xo^�0j�s�6)�q�bS���\��YjhC]�+�t�rm���ӽ�oM���L��ϼ�Dgl
r���:V��<�\��3ə�j�����ʬ�N� s{};^ϡ��{x���.�Y�Da c�$�Q;<;�u��3������sv'Q0q>��e�MUR��{�D()��f�Rڎ>F������O��Wu���AX�+�n�+�9&>B}ݫ;�O�ς�����ڬ��{/6Ъ��CteQT��]2��q��HMي����wR�/s�v�r���v��Q
��;����.����s�=W�I�y�On�:c��֗*��A׷�7:��m�n�
Łvz�R���t�z��kي.��go(_�ὗ����꺽�e]�ٸs:�{>�n��u���z�xE���Y�!�*��wb�ADm�F���k.���ȑ�6+GF�j��;�{v����k��Hgg.2'He�KC����T�}��tn��@��e*��f��z��������9���E����t�/"eh]ِ����}m�Md�0�YSܷnU�&�RW�T��Ap[����������??��ywU��_U��}-5W�q: :(���ڶ���w4N:O�)ۢ{+�-CgB��f{6m�[�=k�*�"T�������ye����{V*d�Ikal\]U�W���I���W{�e��LGF���u�]!d���s��������J���(�{��g�{"�>��к�S�O{P�-�o���cY�����T��5�̞�:t�<�����ۓ3;���1��G�vޙ� �t��V]b�:H�����2�o��-dL�r"�����k)K�d�E�5t�"��a{���<�c�ս�g��QCeM���u��m���P��-��n�݉����8�u�e�w �3�lڵ��ͼΐ3b��(9�`�L��{����}�6u�˩,H{Ft�W�o�ӛ����$w��ʍ��4�˾�9���{DZHUWsvyW�����:3{'.�.�pN�W����ܳI�%s��b�'q��E��i����g^�R�mM��D �c��_s�6�;�����
�Q6YՖ�qӏo�kǍlkZֱ�c�o<t��KdڝKl��[�W��m�z��7.nG"��GN+��mk�cZֵ�cּx��>Ro:���K��-�Y��N�rYo���8�o<x���kZֱ�cֽ�ޛy�RuW�N�gSY'Uy���_?;}5������\����v���Ǐ�<x�c�5�{|�ԶK��N�YmM���6�J��ׁ�����3sEo���K�澧+>u����{;�V/�-5�T���.G9n{�g�oM����3��~+�y�|^mzm'�t���ܴb>��E^Q�yr<�h��j�b�s�B>����x��3:�Up�d�����9G�d"�<d���>�n��}R�����&�H�h���q(�������Ө�ӨԿ=�ϝ￙�rx��MϮ{��� ����f��j�u��O%}�t>�̕Yנ�5�F����~��΂{�}�;�o��xXч���]=��������e����6�K�}לp-�m��]����oI5��.�7������3���i��AS ����;�s����n)�`�ع;�fj�o"n�� M��������2-&0*^��b �����P�)����s�]c���!O���,�q(�!�ߪ�l@`<9����~���C�᥸���I�t&�������q���"cn��Ded��< ֶ��ǠH��8���t�65]�he ;X��oI��1��T3��+ݵǶwg� 1��q����رi��l��_��9�Yz��g��t6�5�^�j����5]�'��&��Y�|����7ގ~�%p_wdq���?��C��-��B?JN��Lg�1^��:��J1?@�bb�;��xO�h���HC y��.�]
�D��/,���	���+��8j�u���M/,�Q3/�
��׽��ϡ�d�=u��}�yݙ��'[:=Y�~�����4�qX�y�bT����7�G:}+-�=��m���j���:��˫�]5�N�.�p����.Ӿ�sл�D�s��~�C���x�5Iv�}@������e�m���[�_�}%�&<�ɜ6��n��_�l�������.�� ��O  �ʕ*UJ�*��s�f���9����z���}�|�@NB�	< �0{B4s��0|�_��X��}��}�;rov̓}��'��������y�lz�F2���������@z�<�/g3�������ԙ��k�>}�Q �MxUPH�P���[�OM�Z}�Ͼ�����ؼ�in��+B�[�"0D���}�n	3� |�x`b��|!��b#��=����B��!���/Gz��P垾�H�M̚C�權q��E�q���>Ϫ�~5T>0��>
>�t�&�a��j�󽀚����	�9�ɳ�䥘X���iΗ������6�~?���?�������A��P�P�<� Xv���ٳ� 3p���k��|=Y�F݃b�ݤN)�����O�.�_T��v�q�V��a�+�XA����,<��.���8��37�unw���d����(�0�����RFCM�հ��CT�i,1,�����U�46X��2��'�0�f�����snߺi�s��M5���{��w��JU�� Pm�&�*P��?à^��ݨc;^|߯>����l�YP��n�r}��w�V-8f- :�� Y���i�� �}B�XOM����-�������Vz�Q�=;z{{3]}�k#��y��� c�v��=svM<���+}�W�]�z���ƨn��t�D��X*+Y-��*�4��#���h�=J����X�}�L�/�+]����/I�s��f͜�S&;�˸N�b��ù�p2������H���(Hh��W�#ܶۆ,��*f�)�ҡ���J�J�J�*�$XA7;��}�}z`'A![A��!�T*�+�}t�Å�k=�_b5��|�0��ǜ@Z�ڮ��wPڎ�osG�Ϟ������Tq{«�Y�<,�.���,,y}�B���>�D������V�t�:}���cxKEE�N�n�{�/\@N����N)t�Ϋ	a�,��3�����ysIR���!�iJj,:��5�����.���ɸwE2/ٻ 5xsr��H$ts� u��(@�����yi�;�ܡNfq~U� {%ĞRo	�P@�Lr���Ǻ*��v<;�G�ר�/��A��,5�s�t
�T�3Me��4��`����_�vB��O�U�z��:}W��yD�i���Pj�A+ӳ��Z;3�
U��,�<�!� ?�Ae�=�[�Q����k�&=��\�;�����j L0��Y?O;�E�y|�H�� ��]ĉ4��c���>��hn��Ú���0�٤��	O�in�%L�tv�.oUi��������p� �0``�N�|B�^"�7������ݚ�Sxn�`��u���o(�^ ��~����/aTZ &��Ο�a�p����]�9�^��p�֩SebdZs�����:���}��x�3|>�qЫܬ�B�j���E��\�e����"v��K�p�������ە"�u�(�����.aP]�4R��يp�ďvڟ8��t�5�Wfl�W_Ltt�ԝ:t�ӤO}u߯^|�<��|�������M�N�}t�R�7�[ɾ�+��W|S=�0J��Г��Z���0�k�Cqk;o�{ڜ��z/MBE�� [6�;T������t>߮��|���m���;s�ޫ����ٹ�x{��[xp��� y��t�!�d��|��a� �3
�&67�5f��*��Q��em���V�+� 
Op� �x ��9���^B{`;�'τ@���@LhY4)8���o�Հ0�����;��%nl�UU���1�W��ZQ�5�U�>0���G�v���L5��x�Hiٕ�yͻ��p��|o:�0,�)�d����� %�I�> {���Jα�q�c>����^ԭ�������I��K� PΠ�	J&����f���>����{����-�����c�C#~#N�Fy!�}�3�{���z�����&�S�|�yN4���~0��[�5��S�r�'�^�0P�����~Ɲ��k�� ���� d�x�0!e�'���'�}d�Ƿ���幼!�rۮ��xx�r���y��\H/���I�B/!�W,���t9a�\�Kyzcŝcǵ��Ǻ�|�2qlWt�0�غ���
iǃ-]�óZ�]�@�g�������gp@N���h{��wG��1!�|�#��P$�Z������G��#�mؤc%gF�S���\w�o{�R�ڬ�}6��/1��',�����}:t�Ӥ�ө:t���g��o�:���
��B���I��a:���|�R��-U4��,8��w�����z��Gl�Uuڬ�]�=���O��G�T����98�0@���s�4z�cL�޶�1M�p��onr���68{�?�``ˀ׬oS+�>�zJ ,�`ZA<������A���sx�TF��}����OU풇�6x��5��>k8�G�}�(t�wO�ah���=�)+%_M��yW�Ҹ�3�������a~IX�Q)�ߐ�Ց����Q}��oh�����zSޠ�>�/�*mIì��Zq3��������0�_|{�ڊ�el�W���!����/iy�[�u�3m���Ni�<Ϡ�q=Yt�@7Hqmbj��:l���0���u<��w@�[ ���vf����1�uZ���4����wf�\8W��9�*g`>�Sv�Nz2��p���鼫{n�<�Y���Y�8n�k� "y�(�j0cս[��� Jj�ˡ��0�$"�>�_��1(h2���e�� ��׶��.�ib��ɬ.R}o�+��7�s�|j/l��Zp|���������vʾb�݇���ih"��n�m�û�X����f��uA���}�4�W���/-��iH裛��<����wZ�F�9JN�4G��Ɛ�ٹχ��1V=�f�]d���r4�}��%�8�{t�:t�Ө�Ӣ|�����7�={���X�g��V��j�Yc>!�@�V�%Հ�E7WwW0��9"Ok	�x������<�[��!x��{��,��N,C�3�|o�y��p����8چ���z�4:}p�F�fc2|UG�1����o���X�m�]՟�U�կ,cK5ӤtyW�(����R��`���3ߒ�/��}Y�zw�A����������zˌ`:���>
��aC������X<���@���Ԩ���g��a5
��Ag���{����f���O���t�~���Q�*�&��,(�`{X��ۛ��2 �~�Ul��.�l�ly��a�`�7�sUyH���C����#��^w`�3��B��!�����[D|˪��i���޼�\��^�ɺ\���*�� k�|nO�H��TF6�S� 8������U-T��6㞳���W�z�Xk�,��L�,5������8Y��,0�m%K���C�M�m��j���iY�ڮx[Ho;_����@�	�v����A�'ھ�wX:�_٤ҿ
ۉ.K�&|f�H���ɮ��z��� �C��8`��k��J�
�.�c��s��^���};��"4��	�fmT�o~n�y��i��a���������PWF�)����f�vθ֔���?]T�����&�
�!�K�_zM�B��/��)��v�M�����؆<8zC�8m�6_u��ut��V��Χ8���^l�ƽD�Ka�Q�
KM�e�M�U� R�J��J�*UN������o�pN} $���<jS��?1�`��=:@��գ��?�vP�I�|�D_Df�X���n;�3�t��}�ξ��bg����'6�uh=�;��|L}�/]����Wˌ��A8����lN�ِ��o3U�=����K�dUr�����W��y5P%��J�A9� <ík��`kVp]tk�^5f,<�K���%?���gf�/c���m��CK���ѡJ���ǐ:�>��f.��K{k���'��2k+Á�E??�ˏ�@:��x����x>Ġ�k�����GL�ry�թfg��▇�n��'u�]w�`pԪ����?L�|p��`�<������җ�3�z�^�WI�=e�c��"���p�Ʌ��/W;���ˌ��n�	�L��@!��<���~LQoI$�V��<c��c��tSq~�1�>^�[�~ ���	�����3��@�߇���f;O�:uĵ};�=�ꄑa&4��V�C���	�������NBʝ��	�T7����xw�������;�JU�vD�~�æ:�Xae�2.4'o:�n= ky0��=Z �WT�	�֟�y�Z=��<Tq����w)ǔ4�1�5��ݵw�GcV�t<��z�b���T�U�W�j�2p��Vd�J&��'t^Uڶ�v��0��3:[ݨ�s�_r����_o0J���c�u.fw���'y�ӝk��oÎ8�:t�:t�#{����}|�y�*Z���{`��ae�z�>������x��v;���p)�ê�{��F��=�۷�?W�=m� Y��X�z
�ï��|�M�[����{·8:�)9��/^s���B(]��qPH=t> g���m�-�_��~ �Gqq�2t�ݚ�B�X�P���=���<S�xp���ݖ:O�p8(ǅ3��yw�p&4?{TP��p-������d����Ҁ�-�ԘP�ڙ�!y��~��a���X��,�~�y�K��(�S!��i�7�N#�y� ��j���Nj�����Lޠ<���ply�dt����	m��S�!�I��]�_��ޡ5R+�+���`��h΅���B�P���	;y���TȦ�Ĵ�ӳ |�	R�^h᩷v/i�W_/��[��b����1L��p���F'T�`p��u��:���c�����nH[�:�����ޔr	ﺳԵE���_������������䯁v�÷�y��І�	�H���<Pt�^��	�&�jN/ԘsgMu���x��
5�@�d<jXḄPy{����\710$�a�Stv�l�[i��;.���-9_�����*��5���6��ݯ��+$ޡ�I�qs�C{��fo��8V|������r�_����"7�����-�콭��L	�Ÿy}{}=�׫) �R��R�J�
̋�K�PM���#|���b5�t������~"�XՕ�M�q.�1�����]�3x�/�Zg��``:�����4.:�W��E7���-�]/1�)��Mޤ�30mp4�y%u��{���׾x1�����Gf�_e�_�?�w���_d���o�c����TU��^��<��5��3� ���h44�>�|*�(��>����t�p��/K"�����_�4�
��j�v)�f�vw�<v��4����x&��N��������m[�L��P��FJ>pV��"��{�EU���\�ה����9=�ߍǇT�� [xr0A��=�"���h�����Ogz����OU�j
x\�	��)�N��F>�( ��r!��lk���`�u��V�]�E���+��0	�x'Wެt	�V��m�1P�peCG�����
��9z�b�������b�~x�o��8h`-�p}�M|��܎O��ݘMr���U�t�����)d8)�7��v���/Evj�@{!�8��p����|{d��MŦ�߰l�R��$n7��j��A����ޒ+q�[ۯߖ��h�iv���\�<3ţc������{���8(�z��xx�!�HH"�$�J���CoeT�)\J0��[�Ţ��/��r1}t�hh�nl�^l{�p�F�|���Ovo������ө:t�N�:��>z�����ߛ䏝D��R����̭@B�xQ*x��>�Ky}��}PZ��^�{
��vn"'��f6��_|C���7rYK����}Z�p����i<
�m-�-��T�xF�yĵ�a> �p��.֏zw�z�m�Z>��"X��B�;����y�<��&���si�����<93���-�%d�Ƅ���Tޚ$`d��˯VG�ᑭ�A� nAd�r��y����]j/l���{o;-��{=���T�j�����q�s�J���Y $T[7���j}�.��)���jb#�������sZ�Χ�^�=����H�������|�#yEB�*�|�������݋�'P�̰��u9�8zkz���<ӎ"X&����f���A?������;<��K��b��-��_4,���@���x�@�=i�782���H���R�o�Ԇ��	Y5��-��1�.ۖ�r�nl���ī�pI�7��_/��^�^�A.�s��1>Kæ:�4%lc���^=��X���NJL֖�z�nt����G��U{u���A�s��Y��g�AyH�M�H�ˤ�(
�s�p7̙��=�;-?�`f�G���N�ЮP�#i�·���� ��#�^���8�����A��4��f�z�[w������}����o���.f�܍J�+��w���IiNVl�Wuˣ��nӰn�l���M�ֶ�	(���I��}/�y���T���{
�<6�<49M��ߔ�r�;s{(/�=�v��Sv�g���܀l������_v���bysN�~�?J�0Un��<;ۏ�?A�������mZ�5{������i�(@�(>���ֶ����s�F�guM9�����P������h�pn9[V��>��C�#�������n�]\8LӻE�;���W��lfG��Ժȩ�1q�������G�v��GgR�=�y��ʘ癃C̓��﷥8�2���g��k��<�k��P&�
�qiOOK�v����
�{m�4s���NԻڮ�U��;=�>�ǾM�;{OfM͛�	ӥvIԬ"6M�b]^N^,��X�:]7�O���?uA���B� zgv]����f�3�����ڏ�T����&L�1ˇa�t����Mmu��םs3w5��������t�\9&n�꩘/���n퉃�����闥A�Ӽ��{w82K���"7H�1��t�= }{\�P��㣩�H��C(&]]�E�db;k"	F��Y��V,7��*��	Hf�32;�x���`h���P�&2V^��_;ߒj�}&*|q�)!��#�eV��Sf첣$��R;��{��i}�W{�����U��I��k����v�ަ�ഁ{����� �����)�h+�3�Gr�e�`��b)Ōq4 ����!�8`��oS�Ci��������j�Dυ�K���]S���T����;�����!C�;�\�s���)�ˑ�Âm�^b;3rg�l��ٝ96�o�:��������:��u-x�^�F9����"{%�G��5+펚�Q�BL�n��Dn�.���r�3o�T���3����2c�u���>Sƀ�_��������t~�617-#�+K2��6
����b�*8p���<cM���g,���B��3AX��b������ٷC���
��<�F��w<��ʞ��@Bv�ԓ�&��p�����d�Rz�1���n�엝��2�ww-�OL���UgN��}d�x��a�zhu��l��Ӿ�>6W-ӥ[�������8z�4v����HO��z�Y?�k������tL��f���_
k&�=�o�n�����h@��\��r}�e�5�i����g!�<O��N%ͷT"tj��I1S�I��6�����p�Y����$̈6B��n�o�0�I�,c��V�i�$xŰB#U�Iwe�Je���l�-4����#$����dCMB�q5c.C.͒�2pi���q0��d�BbZ�&�`�2�	
���P��a��� �+��.����s�A�+��4k�\���Elv�ݽ���~���Ƽx�<x�cֽ��س�Јߋ�(y׻�	]mKz���t�Ƶ�k^><x�<x�c<x��-�gUl���Kd�n���[/:v���$κ�ӧLkZ�ƽ��<x����<x����Yg�6��D�Z�_*��S�|m�{��t�Ƶ�k^��kZ��ӷn�7��߻��$���M~�b�ђ�w�����l�����"�r�c�\bo8�e1��۟'9�H�������t���F!ˍ��$@E��l��ѰW��P��Bn�ƛ�r�n�&\�����?���a��eS7A-#�N��=x{�q� ���m�{ѕ���W0��
�Wp̯B�#�^����p8ܱs�c�[��!��r+�Q�S�E*B�������!����`��m&�59���~Z�r�u%t��j��h������s��\(��]	k�� ������V=����i�;}N0�#��@�-����S�I^f.ী�������,��b^sץ�&�vg�l�(�6��T�������@]=��!,t�`9�.�R��l���N0I���_��D�u����km���	�:3k>���_]��uLL`�nFwk�]8��]�py,᲼̛8��q�i_��X�@��\��$n�_�n����9/��E�o{�U]���W��=�\�ÃI�f�_��հ[����OGX���f�ק�@{ٿ|��/YY{\PO������� "���0�j�H0	 `1�6ʂ�m�:y/N�aG�+�i����~l�ŻD�A��C�=7�ی�,�L���+ ���(3�V���t���&ְ��#��yF�
����C@���i%��ώ��}�3�V��Ƽ)\�L)��L���A#���[2�7�omta!J�U#IU|��nN�=B��R�E1л+~$Y^˃,F��b'����qj�__^�"��W�io�ʁYf=�+�f��qY}ށ4�u���@�=�1�>8u��i�Q��\s���c��n�
�b�eZ=$�Ψ*�mq��l0�r�/ҫ�`�U�0�$t��I�8����r�-�;{�D�+����m-�KBg.پ���8��d���>ob�f�zw���5�~� ��I�t�i���oJ6j�6�chu��.�_p0���S���5����+�������Of��&��>z`�si�.$0m(NR�cۺؖ�M�,y)�����.�qHy���2c��P��s�������}����L֜]�\��`5�r�l8.y�&EA�-^�˞osX��z=��᫘/H.)r�e��U.v��C�Tۜk����}Z����1�̯06����Aُ���P'��XZ�6�ޫs�'��m��5���~�>̴���Z~;��>��1����j|+��S�'k����	��m�ڵ�ɗu�u��+*7��-�՗)�ua��BU�D��G�Mx�O���u,H����OYݨ-��r�L������bt�[�wv1�z����8�
5j�o�׵��{�y�Kd���d�l�՜u�{�-���7'K��e���=�����f<���<��0��%�
G��5���Һ����Ȁ��c�vz{���y��+�|��o���E$mZ�r�$|���A��f��)y���6�^s{��{�j�i��/<�Y�=a�l!�q�A
 ��o,k5C-Y��� ~`Cc�q��ςό�m��#�.C���gf�����^�E=�dF����%��(H���[�\��1�`�T}Y-vD�s�`��z������Ɯ���q𬕰��D'��[������sM��^�i0������い�rr�TΎ�n��K��h�k�:��:N��:nC�8��-��']]�_^z�~����f���X~�*�~B�/�!}����΅�>�6��1��Scr��Wx���<K�� �7NG�\�5� .��T0�h��@D.�XUO{7Q~i�5�;q�Q9���N8-d��±=�k��Wh'ؑ/1Cx�F�um6�@����v��)MI�fvp���K�㺾>�}<G��:����5|Xn���Ҁ�����ٵ��A�~4�"���6s����IT���!�%�8�Δsm�,{}�#��`:���
s\P{�9�k���|�-���g�pО|Ž���Y���7	<�^S� (grxfe���a��|�Q8��'c(y��V��0b�s�h;�5�J�����7��~�=�Z�Nīy���L��>��.��]���aD�3�8[�À�C\k�e"u����ކ?��G�R� �Ǔм�Q������Q�&)Q���Ҁ��8�mu*^�@,iw��ϭ��^f[�^��R�Ԃc��V�}C�E`<	�9e�Y�<��xw��R{��uק�|���ccT�x0gFS�`4x�x=���w�Y�[1E��7G1ܲ��[z��:�
WZ��i��gk�m�0�n�KM����d�Cɵ�����_ԡ�s�����2z!�y�Fuӓ�	�����(���C��9u�gu.�Ε9���}�WH ��4$�n')%�[��,�Wp吮8�(-B-��I�ן]����y30� �ڍ��f��:��H�ż��3m�9_���m`�~���}/�y���O��k�׀>�q-�+���_�Y=���tP����+Ë�(m8�-��xѓ�[���f�g��*H|4��� j��>Y=>��O�L�s2��=�^D|��Mo�Ӭ L���7����t^��l��F�G|1����^���
W|[���MAϴ	�!km����ʺ��6ʞ�n3��,����#��	�xY@p`} C��1c�tކ󗖖i�,��îg*;Mj�<[�>y�Lpi=�&�k}�h=3��cv�?p����C�]6�LT���a߶����i@x��2�R<��	܎X��
J�cxZ1����x�x��n7
�扒�O'U�����<���j�%�r<6E�61�Crr{\������{�U���E�~~��=s��5
�o���=�n��A���<�!�S��#]�c�P�1/A�y�ӏ
�P����5��̺���z7��l�d�V�f#G(pٸ��rj�*c�a��J�n-#�lq	����]0[���՛m��hh�ڧ按Yh��|B�ԧ%iVR"��S*�)g�mm<mZB����t��DĶLܙ���<G�b�zP@�!EzD,�՚A2��\E�y}�c<`��(�ޕ���-����W6|����^}���/�j�iR��D~���hv�љ�yx���
"QH6!��L�P6[�Ĉ@b1ʋ�P��UI��',�$Wp�8�r�l�q��$Q%�!-$��  �5B�$Pw����o�x���� ���Q� ������|��kv�3Pmq��%xyӤ���\}�@B��=����lN:xk��K�p�L���/E�����Q�[�S����M�@u8a�5kxW- [��Lk���~rEd�|d�K����я�Pq�����k��� �W�B\+h�xk�\(�,{]!��FcV;#,�U�Q5e����M����ia~�L�DzY5nGs�/*yf��[S��$_���8� �mx�'S�7e�k�i�g8��n�v�)�K�ɵ>��2u���a#>��N(�P sz����*3�J�6��IW|H|@}��OJ i��b>[�:��� 1m�o�k���N���������\��8t�)0��'��g���1���n�Ʊ�vH��WHDь�J!��6ڷz���c���C1iԤ����HVY��q����>�NA�\��Ϋ�1:��=�'�m���#3�v�<s��JQz �t3�@��2c��R<.��pu�$�^�g�u��`Ǻ������{!�Z�O��TM\��e��<'�&�FP<y,���+��\�myvd��{O#.��Q�.q�'�ثF	��[����w)J����v��B�t�uD؍�;.b�{/��۳��/tHo��m�b�D�� ��3�q��������M���9ݗ��x�>G�Y�N���y�={��߾�߄�wd�W�ӒY	\q�I�
�D��BJ���[b��m��E��mbEg7�o}���~$�A� ?�mZ�MǇmz��74���!�\Z�&�t��y��r��O�t��IZ�Ԝ���P����I#�\��O��g}�bӤ��Zz���}����c�����a+sxy`��rs<�_��֦-)����%��-�� 4D:1���!��`7^+efWM�6�5�z����^
�t����6q��ȶ��G���/Q�e���A�gO߾���؞���K Q���9=�{�pP�2��wc)�zI���v,�\k��ǲD���1���bo�k�������Qp��p��ղ���ʅ�%�]cݩ�k{B1E�;���L< �	�K��~�Qm�F'����h�u�GE��
H�ɖBNP����?׏}��.y�Ȩ8倠r���zy��z��9����T�sfNJ�ӊxk���p���7�	��%��РV�37���)��
�a�ʯ����Z��
;O��������S�U�@g���mMB��PJ	c��!w� �:�"�1����K���N�sᖲ�K1��]���S7�)�\�fnE���ϔY�j� c$ᅨ�3�a4���!ٕ�	��*��	6��;tK�H�:t<Y8i1ok#M�n�_����ɕ����_A�݊et�����k�٫���k"Q�ПH�aڴ2����&^��ۼ�N=�M��r�^ݛ�wgUw�)�����^�����=�뽟h�Q$��$�}�$�ʮ8�I',�i+�8rĕ��')�$�ȓ߿>��[�׭��瞹<��$�ܠN�J����%�Bz��fpA����P����L�i��+2��Rř��'fȣ<�w`	��^�e��D��4@Eĳ���.�8�]hOp��U�l-�=����M�����ђ�4*�xgxǱw�c���'��0���3�RS�TXQ{�{5��=���� �����+�F���襫0�ʋ�����o��kYi�B���rw�8�nьR��@5T�'��چ<�&B�
�M��Z�#Dy㶵���S�v-I�J�]��xs���+�@4�[^�
�!lm�t@�8���m�C'��;GF���/O���Ub�<Pq|3g|ɎI�)̥�P���U�L�k
/��yr7�~�g{.z�f�ógx�f�ɼCp/MX֝؞uat����F��|^���׏�@�сų忞[]�C�j�����Li�����8#/}>��iͶı簌Su�aA噃���2c�'.��΅��t��ø[z��0-0����	8�)��#R���a��j�g�}W<�b��pu����<nF�0�K���l|��H��v,�r ��9��3	~���H��͓5g�OA��o㝏��7ouQ@�3ό��Wzl>a�������Ň�g�/g��U� ʚ9/��Et�rB9R��q��-�H�8��X	l� YR{yu�=-�o�0��ٲ<���UD�G6#Gc�O��J/���|�w5��3���������Ν�F��B����!P�%?t>P�]B`�֟_)��6�:�
����8ob!��;�p|.�>',g�P%�0|�&9�'��t{d*]֮�;�~^���[h#<��e�g�O���=�BOt�O�`]�wfoN0r�J{��m���'s��tv�d�=l����vlO"�S*����&7�O�]'-�nD�1a��������',-]|�[ߚY��<�dŶ�2�r{�,ju8�!y�D@Mq|�v��C>��j�@z�H�|�Z�_B��G>��ȴ�װ�l��b�����Z]x�?�l�-�o9~�s�W:�u�VP;DQ��eo��F���G���"���#E����{J$�-����,7ݽt4PJY�V;�t�z��+�NV�ӕk�W������ީ���	\��ӎ� ��zi���<�#��j�OE0Ơ��Y�ծ�V=��E;�amV����
�VI�ȩ�2he]e9L��-Q�ğ%Y*��q�������y,����ڪ�^\�]��}j:U��'�Y	��,�����@�u�(H*�߷%l��m=G;-*́����[$����0;����vP�2Z���U�I�u��]�.�	)R�fB؀�LL"�!�L�&4HiB�.՛0��UOM}�q��r�I\q��+�8�I�"y������w��z���yح�r]Q��O���p��|}��ڽ��^j܂�[�rLY�@^�1�[պ��Ϩ�l����]��x�da½"\_�#%�x����c��q|�{�%Rio&��4�;�M{zOx�j�۷���ҹ�g����A�<�]d0�j-�s�%��$���/��ͬe8���4�l欫��2n�nH����K��ǜ@��0?z@�6"�>�� ��==�N���\nb��Ngx��Q~j�J��k��+]'Ǆ1��L/��ej�	���:��Iv�Ʋ�֜%&���^���rct��ڞw�Ԍ�W����e�OZ=�CD�6ö�c�6{���e7���~#@M��ˠ���xwֶv�\�J��&�g:�
}`?'���T+�C�������D����c���#����ٌw��j[��ھ!;���\dr����=�g��돿,�� �"��5�H׌nO`$g�^S;�{zy
��18�/��R�vP��ڽ.�?�NUǧ�D2^@r���?y_W%��ݠ�k�*ʇ���op�Y/:�طyl[
�;6�������a8�])����a墖mu�9��S�[H}�?�A�󛝔yٟߞ�ˀ� ���2U2};_.]��:�Ŵ�t�vm���yw���7�:��1����*���{<+����s�^T����nAI-q� 8���+�99B�	-��w���}ԧ���3�Z���|�a�>x���0twV�w���P�K�VYQ��5i�|:�W�b���v�0�!h��6�P����K�B0ZJ�ߖ�۬�Q��EQ�ʼ�I`=M���T�;����ўn@%��>�-V�^m�*.�Cf�n����9���o��	�3��u�H%����-�b�W�)���#��s�hws�W�|1��(��Ya���uN��z���w�������ð��#��'��Z�d����y$ެhBm�co�k��xy]꾨qީ��Z��Ƀ)^�N�t�����)�Xj-�ǴM��j�Y���ެ��V�#-��
�Ja-�٧�S�M�Ҙ�vk��3#��N��p1��熝���+��}��c� �s��%C�GOs�}�a���ď	��H{h��&x5��f�?(��a�7I�ã��[lܬ2+��rU���W����� ́�46d����j;Ӽ�:#|�4��*���71��<LSb0�̠~/7����9�y u`�<��n��L�t����28�������c��u�h�ږ[��Ui[��M��{���r��gC��ڑ� ήuC�(ٖݞ�y��Q>Cƅ�g���qx=@��F��o���6�yRf���{-iѕwoXS)T�oG�(���yn>o�-�\՚�m���|C]�4��H̟�x1�o��B��S �+�^g[�.��j<d�p��1o���p�b=�*d5����g����b��pv�^�<��+��-�������^���K�ܾN3�j=+�x�m�K�op�zK�n.�!K�Y��s��;Ӄ�{���kG]s�Xj���,����`�"��'i3��3;�0��9���[���U���;��[jl�{-�$����HR�A};�h���=c��w{�4Kv_X����.k��巊Ǻ �/�������lR���z�� t.��Z,�wkZ�T���]�)���ޛ֕�D�on�ɱ�[��� &�4P��T��m4��z�c�9+�]-�ٓʪ��`�3c��=���_z����C�$����4�$���8��fO��d����ޭ�͸�ۘ�"N� �L�c�k�fX�y��G���5P��{���ݱ�И��*>���
 ��7OM�9�gԥ����Ջ���s��ߢu�]�߼�>|�7=���u�a��̨^�|�9��^�xN��۴��n5|&\j�J���qa�X��*eQ܌p���Nd2J=�MK�Uqէ�Ќ:9�2������J0X�G_2��6�NQ�S�n�U�ѐ����*�)�kv�dC=j�9�4�2�LI�u-��"��&˨��{ǞU�Wc��Z�'S�n�8��ѹ5��p>΂�•��M5�\3ʓ��o���X7�Ã�<�9�2��{�m'	Hm�$9���X
��:Y	Q7�Zܜ�I;�"f��;�g"�Q�P���3H��)\�ʡ]),�k�{Ʊ�y��uδʴ��Y�3��Ǯ������
s�7�]��ŝ�8	a�'h+`L2z�(Xy�s��D�s��}�6����Aյ|���������89�m��2@V`����F�x�7�p�z�9��^Pj�é�FLg 9��O׳���#���w�)��za�0r��u3v�`�v�:��u�\����ݸ�����̫Sa��[�m��P��݊�]˅��������l�ƃÝ/^�W�x�Ɛ̓D� �h��%�[n�E3)�G�nݸ�������Z�kZ��۷n�<x�=������e������޹��Jk�����؃��ݽ���kZ�ֵ�Z׏ONݻx��_"�#󫻪�h��V�d��]8�Zֵ�Mk]5�v��۷o<n�{�նիe��-��)#}+���{u�9���]Ye�]8�Z��ֽ5�tֵ�ǧnݼx��m�KV�*_�u.u:�d�K���~�do���4D��|qL�B��\8H^�������t��]�sp����)�b�9rH�˦ 1p�+�30��u��/�u�����B�)(H�.be2a&H#$�����S�A{���O�|E$I�t<�+��Iu4��d�$k�ff.F�[7��җp��n�����r��9�n���=����N��"��ۉ"q�8�H��rD��jċA-i
Ib%�Bl����ל���{:�>��ǂ6t�b���:���O%���9s�����f��ou;���E[h�3��T�{��G蓣����W>YI�������K�?T�1���I�����[��U��[�x֘�}�VM�OlZF�$�H&>�d��C�<�{q�>�>���x���o[�c�8u�ݽ�O��9O����3���uY�@��	$�A��a��Q�}����������:hY������D�!I�r�;	��3��T[!�*9*�Z����M!��f�
ƈ��ME��-�|���pɶ�O�0ͼ�>wk�R�NlIza�k�w<Kg�@�(~��Y�S�#��=�7)p���^���v�5i�'��V�ѯ�8EE���f��v�� ��p�h*���kF�;�b~Ļ�oo]_���:�;�a#X^����:���������*/�w�c����)�R��������޸�\v������ ��#�/yP�2_S!wE�Ae��Y�W6L�����p�8��0/���^͜a��5dG�xe?0�X��������/��i���V�	}�f�h�w��͐bWv��-`��e���I����#�2�MW���U�|_6�K��O��|9n�)���x�<����7���g�%�5���N+ˑWz�8kk�*��Un�t���� �� zI�q$��8�'qă�D�3��
|���T�uy��@q�dc*�	�X�p�$��ع��1QqQ�+ ��:1��5���6��)/c����_��G��4��E��It�e��B��f��¼���!��}�|𝎱�����8r)�9+�4�B?0�ޘ�[�����Q��׊��A
�ۻ�y��3���	����a�U��ߋ�X�7�c\�1��꿚e��FjQu�Z���ޙ�ۤ�󼨑�ښ��j⣂��-.�����h���t"��W2����2{�=�y����/c)=��7�oI}nG2�b��=G8��0�(>�C��!õ�V	���a톷%�۬�����eb;d�2�V)�uo���u_��mON����pf�ٞ|CO�`ּ��ƥ�u����=�y�33�c�J�O}Г�\E8�*�ޭ{a�6Eái���vŸ́��dG.�����>������"�x�ueO�]'-�m�-!���x�qH5[]�(3p"X_�W^���+-�(����._�f��=�=g�`#~����������&�m�Ͱ��<�#r�"��wo����ڑ�\:1߫f��&�|�F�\|dG� ��N���Z�#�ٰ���B���Q�/s~qW}�Ƥ���}�%y�{��,p�ӯ��c�<���ڙ�M�'s����7n���%�m�$��!�l��T!iFCl�� �W�b�EN�prĊ��8I9d��EP��ũ���׫���$�1�aY=C���6u4���eh]�G6�|��t<_��	�sM�hm�*}-�K"�|wr_�(�|n��f�_z �P������/�v|Q�-^+�+e�[;�]��p�7z8���'�v��U#���$^���)�S��H�4>�`�z=ŗF3{Z#nl��6kkS� -�'����"kc��^X&���C6q=c�:0%޽aŶ(Ÿ�3Wۥ^��\������ݱ>q� N�Ŷ�JzIN7�IN�l=��<c��v�[Tt�a=;��v��_�mM~l���ָ��=��܉�t�'��i��͊=B�CtF9r�Q5���/�ML��{��P��xN2���Y ���-���=1)���b�M���i赗|g�i_�����ȸu@�p|��� k�ä}�o�AwF{�5��&�/�̚x=�� �I G��>�2�[�Ҙ��{�<�a:���$mz ��:�vNQZ=�֕�M�_��i���S��ww�mԎ�X����İ�`9�����=?�������/;F:� ����⩠�ݮ&��{�vRR-�j]�$I��q���F����Y���de�" ����U�W��b\v��K0�·I���*�ܽ]b��S�k����rL�csv�;>�;�� <��}��9`�8��8I�I+�9$I��D��7�7ϯ_]�v}y,������G�L�3�L���' st�t㱜&w}׶�]�۟8�diq�n$�7��#�qz-�\Ȓ�~�R��bi�&�ݓ�(nW�{ι�0�w"�����@xۮ�M�K��`��!�y�lQ��K�������kק��O�Y��v���[���9���^�]�_�iT��BtS�����k�#�ɹ�s넜lW^N�^5�h�+)��"0�a~8!�ќTY1d؞�WjӃ��E���4߱wc��Z��=��tv�H�gW���D�y���!��D���}2�۫��݂$�Ѓ/F>���K����M�hY{������LP�h��W�#����t��d�����81�f-m<��6�hl�󹍲���~�y�߰`�	��H{�;P��	8�Z�F�J���>�y�֭n��8�ػ���<�jg�lr{w�<0.��Y�L�`<s����d���M���[ �D�r�A�w]��7�v3��C��@��Sz�*�c0'�2�}S����O���}���㽵������?����P�R'������pVp����C�s�h=��	�t��nr�<��w�j]���h�	�0��&� ���`��<@�!���I�l��r��ٸ�(�u�Z�3c"�ѲT�(�����;�����'�yZ���7׫�3���{z��ǧۈ8�"rI%�-H�8�#�8�!�$� �ٽOʛ�96�R'~�I�27�}6�*;�ZW <&�c���0�S����;	(*�=��n4���:��$��.�ǭ�{ަ7D��w���*�L"�?s��Yь��7�t��Knx�8nOl�Ml�9����`��oXM׭R+_���z,�{��q��5�,h���Y;gD��_X�@���u��s�I�n.�1��m#4_��-�L�����Pe��g7���h��d�Z�[f�^��9����ӗ�������S��-��j��l绉Y��ʨ�a�E��y�\t���!j;+�o�E]�!�:�p[�RX2��{��}�ɭ�̓�yō/we�		��;���>�Bt��ǭ>����Ou�}n���{&���.�@����\����:=o�=��,=�`�]t��,xq�T�~�k�m���=gS1��ۅ�J�Nf��q�ߛY0&��狻5i#�>�\/d7����v*��'�E���Y��Td��b'�O+�4�P9֌�a'���33t�g�N��fe���[G��ѿ(���8z/�ͼ�D{�l]ק��7�v�u, [���%$?~���UU�ݞ='���=�W�?{b�y��ϰ�/���u]X6b���r[�4�)Ǧx_)���Do���G�����5�A�N�]f���xa� ���߃�8�A�Eq�"'q��I�D�"��s�����Ͽ����_��;�b�(���,v��W�2F�P�9�B��a�� �3��ԛm����b��y�b��8w8�(��bO�AÕ�>Z�^�X5��/u3/_���:�$�������qe�&���<0s]]������8�XJ�u�����3T H��c�4�cw0�N������g�����\���E�}�)�ׄ1n���g���F 3`�L�^�U6�,&��:�ǥ��S�A;�9�&�'�K+*R��_-:ԭ3��+����f)��o��Z�Oi�	�O����V��,��F�Juat���+cf��|���K�,�����;˗�h����vC�A�����_a�i/���a>�J��r�o9�ފn��afY����G-���y��5�Tq1������,{�}-��yO����"�$�\��U={���95����3s�}��H1s�v�	^�<�с�1�9P&>68К�������2��#�a�_�9c��j=�wBe\�����'�v���[@�#Y���+��mL��WzV�C_�ѻ���û��}�ߎY�.(�D�i#+H��&MVz.�3�ΌW6��H���fv��D#��(ξ�y"|K�Vi�PyM����G�G+\z�8��χj�	�o�E��2���^#3�V/^��;�'?<^�%�l��<��5AU ���R �e�D���K7Q�1�
�k���I�%���Iq� �+�8���B̾���y�>��y<���,��ע	�ko��EV.�/K#�;�3�{κ	;�f�[Bzw�p�:7<�ט8�2�Ƨ�5��]{]��q�\&%��L�e1�XH����{���6,�^���g{��c��B���p�ʮ8C��g���-�Suz:FO��9Օ>�t����0U��3���U
C���<���4�!}k\;�q^;+'-{��i�0s��i��z%�k�x��4z�w��b���/SI���R�C\ﯜL��1�����}Q��W^lU製O}���P�:;J�s^5�&Q�3��� k��<4۷�R*�q�s1W��\ίn��3�1��#ߕtDn��O=��jz<M�ֿS��ĆA"�^m���o��G<��B��B��l��5$r���� b|jgXdS�����v��<ilD�!�&,)��i��}Oӎ�u򸇻�>XF�-���ӽy%81����GF�sd��s��p���ٟG@���V	�1���n���7��Ad�r�M2w�-�ݍ���'��a�n�[��I�V\=DeC�q�����2�+s׿\�<�'�H_0�Ϩem�'�u��ά5���ĭ����FK��e�$qj�=��*�Z*p�z"5ON�,�0.Zr*��ozk��:̓vª� x||����"q���q�$'q�C �` o{��������������V-bLA��,�Z��!���\cF:b_s���=f9��kv-�5����>c�i{�|Q>�+�®ٍ{��L'�� �r9k��(����3Եs�-�n�k�NrN(I�9m<�}bz�]_|��W'ׄ>x�h�">��������ma�hĽ�uVt�
#���]6[׋�t��Z���ڞF�3M�j(�=,�Nf�&� 껽Γ���C�2ׂ�ۂ�DϪ;����]�f���q.��Jk��>s� ���8ɝ�>x`���`壟X����&��d��+۳���'���|��k"	��7nw����p��xB��	�ש���i� �8>i�~�kZq��O�VלG����rp �<7_6��0ܞ��V�us.�Xx ��AV+�]Nd����PE;S��y�oU����j��y[��X��hp���Qdœ&��pu��%��G@�<l�:��"W#�ҺۮKx�0i�)��y���a�dg�d�;���»�4�G+�վ�4&; i?b���eh$[;C��PA9V�m;�N�XZ�K&Z�3�R����T-�����eW��'EݷX����SV2�9k�O�����:�z�7��t�m��b�h�T��W�~�n����;�~u�~�۷Ӓ$�9	�%q�!�+�8IʒIjI-����R�83�}�a9/�t���2"F��z�pi=��`�֚{לx#4�6�}�����5��y�-���ק�oM���m�y�!���ZK�ϙ�Vc�QhU��g��l��_�/N�aFѝ��}�"�k�9�;8W��z�!���ȝ�*s�9=�3�����g�q	���*��%1��iاTZ|eb�`�z�����d�U�97�kyV&��8�6��5��
��)�Rx>��7�x՜�O+��i�}q�_�Q�t�}R��/w��x��b�_ }��K����u�����vfe��h�S����gf��]z��iÅq�C��ɴ4����6� �+��]�Pb�_��-����v?%�^�	^�����b��t���#<�	�n�	�Oy��Ï#[ͭ���z�K�����D/�/� uPAC��3�.�5���M����$�dN����2{�9�-|��D��?o��*=-�۴�$�q�KQ �in���K��Z�/\�A�S��ALw�@z�c�|H������5Y�?���l�ۏ�����T���Y=�N�g7�6�ey����*�<3�G��`8d�ǣx�@�K�F�d�mF��x� ��M^���s{!p�h��o���[��z���N]��m�A���=�[C�7ˎ�WQ]'�R���~	�qq�$��8� �7��'W���o�&.2�S����S�ks��MӖ�Y*q	�~c�[�C����3r��8���	w�8���wBOm}PXH��Q{e�JCT7���������l��E����Ϗt���[L����ԉ<�^<h?%_O#k���'���'R�[V�M)�2�lf�mS��n�^��/������:�f��n�q])���i=������@��#��t?T��wt��Ϗ����#C������HeKxy���V"4�SB�#538g��P81�*OvgR���f��䀹�+?s����~��O]�X��魳��ȹ���[�uB|̮��옴[�uH�Hπ3q��ne� |ז|XR����̫��.!7��k�02�Ɩ������bk��rX5z���(5u@o"dۇ��`��T9זp,!�f�	�p�'/�߫�I�B%�>6��^?�a3�K�n֏���O�������'���ӅX�,�d=���]j��0#���K\� nʟ �OmDkH݉N�˥ Ú�O�c1�f�P 
/75�]�䳋�</�ku}+����KM���F�7}��D+;E����*f�>�"'q(9�h��g�����s�Vh���rN�>3X/f��j�R�S��2s�ɖ�3FL���V�<��R.�������̪������w4�Z��i&�v���n(�/�9�8������nJ�ͧ�K�q$7=]sD�!N�/���M�0�`�gmxƦgS���R�H�r]C91��F�T�}|�]:�ܮ��h��2��w��񌁈��<*��U#��3w�ͳ�w<}�aP]�p�<�5�E����j�澨1�3�U�s7�%*·d�vg����#�_� �n����8�4y���ߗ�GN���(j����?�cP�V��q5#�
Qㆪ;S[��/�+�&��ɀ�>��$�ق��g�A�O�j�?����Ȣ9L�ך�NhW \{����s�W�����=��c�潹i�n1x�Yc�B�f�`�:�D!a�U!���F����&�vu��>#�'~~}o�w��ب����h�}ܝ�w��e[��9�{�>�
Ub �c�#%�v_L�gX�b��,�2��[#��%��"������^� �$�6�S{Ӥ�55��
͑u[M���e.�����ĳ Y
4���kΟ�]�MǕ�Eʤ�7�l4	%C)��ߌc#�Iv( ��B�ɶ��N��<��QH�M;�З{8q�U��o�N�rn�I�)�RgV����]��7�U���|d���ء���(u#ğM��E�4��oe�"��`c<V�J�|4����<���毵m�c��<�if��PGx�u��f�����ׄ�X�]Q�~4'�[[�8aw H���F,�Ȟ�^���Wt|�|FV��55�!�0�}�\�z�b[��
������節�]�[ݼ)��֩Ax�
���(;����;�o2�cQ<< �"-��8�u�gg-��vlC_nS̏;��ʨ�7{{1N3�=޽fIi���^�6iWf����D]9;���r�O�td��`��i�ׯͰ9fz�%�c9��B�e~s<�5V{��1��_���]4(�܉�Q�h���7��}��W�H$����2��G����B�����L��w�g�դ
�Ɩl�$C��ɘ6+�*�#r��tzs��V���w^�?�N��	�t�F�˳#���Mʸ%N��f�R,����3�롴w�<�(���S��2p�����p�	C���1m1AGB�Xc)*o8�H,��C�p#u��3w���[����/��V��ӧyyT�qv��0��t>��+�Z6�r��hv��kdZ��f>�3n��&f�����&K�N����'s:�{13+�g��+5<��b�S��`�x[�9��l�h�ئ�;��m���s�8��/P�t��ޖO��z�[Uz��\Jz��:���}��q�dX�=G������=̥�u��<����l�Y�7�ǥS&�\��.�FV�<{�sx���>����]��0%��� �*6!'l���
�(�Ŧ�4I� �]7OlDNӦm�28M��^7DX�F[���!㎂�xR
;qC.��I�L �n�m�qE"-�&l��2$\0pJ%H�1D2E�Y6���zڀe��N8l���S�Kn���	����ZQAٹ����}�A�y�j^sݷt�w7~.HyҪ��κ���x��{{||k^�ֺkZ����۷�6l��Z�_�/,o9� #! ��>:%&	b$I(Ax���Zֵ�Mk]5�v��۷o���w��������_�Ȋ�B""Lou��2`�^v$Nnb{7o5�kZ�mk]5�v��n�<x�~Rb����+�u�HR��m)��f�ݓ��8�5�k]��k�k�o��x��dޒu��,�[lmu��K,�r���>��|\@D� W�\B	4����n�*�a7���7`�I$��$��u�A���3,��fDƄL�I"h��@��0d9�LID��}wW��Q|r	��4���u�\L|n e{��$�p����@��$��71�d�L%(|�#�t��ۅ{�=)�u�"�(>��Ȥ�D���A! ����۾>��=���#E)Q���R�W��7/�������5w�sGu^#��}�����^%��<�,����FGh�����Vn�j�D+K��J)I��
f%-�,��_�����`N�0)ӧN�:t��P�D����n���Y�Qm:D{�ө*_˟-���fF��]�C��յ�)��,��S�%��e�N��79L9�/\5�A}`����a�`�Q3�����Y�S�Ƃ߼dfl�z�;���ka}��Ɩ�:��� x���<�B������^���wsG�l��UVuR8y'���~N2��t�����=������K�\�]u�|�cH� Θ-5|�W�-l���^d�1���PҳO~[�5���1/c�i�b}��"9�p�
���.���1v�5i������:�ULS��n�%��w9�t(򋇾�
�X��q���{;�Dꘒu4��}�`W����7dr�<ŝP���l�Q�ጬO���29��r�Ut��<5X#�����~�F�w��G�ec�|N���ϔ�m�e�y�=����'�gQ�ѭ�T�����n��x 鼰�|M'�\!�ʺ�zg�%�$6e�Ʉ�z�ۚcoS#��&�\������3&�ޭ��s^����f_��tqp�k��} s���~���HatJ��ɼ��=?�Zt��)�F����X!��'-�(�%��+���ppoƠ���5D��k���go��z�0gA�0����,r�ŞN,8��^^f?uŗ=�����`;"��ĳ�i�J��r$�9$�88�H��bU�I}����o��oԜ�����d�Е����F{~�| ߙ^[�z���T��ֆ~�M-g��+���q�K3���Y��B�>N�a�{ 5|dWB�T!6$r���"�ր���}��Jww�k}�j�L�B�a��z�<���4dzS�[s��q��q��Z�k���)N0�����喎���krzm馮$�vg\��d�uA�#�z�k�|Z4������`�Fz[���v����������}XW���x�VCVpA�?'�2�u�^�����?Aρ����\K�Z�U�X��%9�@���)���n,�����
�׻�d9Xd�T͵A�De�t��ٙ�ŀR����::98�	�ԘԔbz|�<l[W��?�۝����A�n�M)�U����8gDg�uB`Az�-�[�I�z�<�Ўq�{5�����g���'�c���O����[��� ��8<�{��w�&*;׎H��}\�{��5�D^��?��}��ۏ�.�ʑ#�_!��.���ͺT�'���Sl��j����0Xa:]X'�ql�;�5cW
�+��]��|�gV��Θ)�L��7o�O�a���YMNZIԒˊfؐ��Κ�赶,���GY���,'�n�dݬ�����h�X��r�=��v��s.��خt���y�}65�W�/��iW�t:t�ӧLN�:�d������r_<+���ۮ<H�z�?�yՠ4|��g�n� ��Eq�0͈=��������0?O�~N��.O��5�'�{��f6������c��~ ����D|��ng���v��{Q
j;���q���C����6HӃ�f�+ieA���Ə@��C
�Nbc�6܀�� �*���Ky�۱%���2d��ف�<��C���Զ�;�ʩv�6��G9L!�x&���}�VŃ���M����H�B5k<� �H\�W6}���;�Qէ.������ӹ��o��{{j[���1'C��Ňﾧ���}�M��Z���k�������i�d����ջ]��3+��gO��z.@��E�n�Cݽ0���?54+���6�/�կPg8�� ��r����A�2;k����ɁϐEu_��>=�a���s�]dN�8���ϡ��� Ʋ�|�4)X�I�2ۋf2}7.m�'�4�z}ФfFV�<pΝ۝�F���p�Tkbݮ��*�ʄ��oGOs��8�w"�8�7��g�W�1�WA��T�7�Gа^�dEٽܛ��(Y���}���p@�/�9o)c��P�ᤘ=�8�q�{��u�7h���4�gvΡ�M�-���R��aM����n��S;/�{}�a��2�z�N�:t��tiӨ�� � FKr:��?ßeā����dq���x�(� �����_�=�='����\:f�i�cs8�*�g��jD�#�1��ӻr��:|����y����8&)����<9��`֣�<\�m�����٢�a;i�s�Q���}WI/��d�6��t�<�I�����=�˕�C�3\z�aVO����~��q^M!�KVRC�F�4|y�@NWι���n��4��}���U��*q\-u&;ǟ�:luְMm���;Ǳ�M�;���G1���m�km6�){49#g����dV�����N��v� C���&��_LW���Q�;�1/����5U>��w;K��V>��^Bwfe]R�&�}�-�_f��J�%ZŲS;3y��[jz�ݬ�n���ۙ��� ��L�|Ht�T�Wv2}�*�"q���d&����= /HO�'�,ᒻh�s�Nq�+�L��5�܎qZ�<�E��?��$dN�,�;�F�����Ɠ�5w�_�M~�����������}����O�!��)±
���;��3b�KH�ｊj�+a�Z�}9+/��r����B�����Sh�+H�h�75�ssti�l�IW/e�+9i�g.X��C*>��.)m���a�PȲ6��-�´��y|��G�A��Y�>3��WW�c:�vK����]�_^
bl��jr�ݸ�`:u
���u1��VCԹ��2
gΉ4i*�m�Qe�E�j0�E+,�ME��V��aӧLN�:t���µy������+��M?}��
�~0{��$��(����W�<ju(���C�%�0�̖��z��Z��M�-�yg)���J�{̎⮤M�@�ݝa#�1LK��8>�ؼ�g,ΡW+��[�o�(����^�#�����Ps�rǠ��"xJ�-{�"ޭ���F�&c��	&�a���χU��IA�R�+Ҿ��;��Ƚd"�,ħ��ҘsP�wX���Q~�?��G��sv�����jCS.+J�,�[�)�����x�����p�Gu�]>�x�]�kq�l*�6v��a@.��"�u�Ӿ8��3�@�G~��cæ��gټ/|�Och+�'L
�G��-{>��뛿6�I��+>����a�xuӥ���Jlx� 4w@�}�N��������,Ƨ���ݞ�l��S�B�O�gs��Yutk����f��'��1F���W�ݜ8������1�_Bwf��]z#[��A/��Y'�x��gR������Z��bެ�#�!W�A^���[q5Ϡ�h���d0���@w�p3ܣS�=��x
�Fdsգ$�`��T�"�y<�Fեzv����,�ٌq��s�Ow�E�,����J�4+��[5�2�$M.֨��;��j���Vb�FK��u��D\wl�5v6���n<I��ދ�Ʃ��o��&0�>��jL��*��7N�0�Ӧ�Ӧ��:�������ėA�C��ͯ�~�f�z/t�#�d�^3�X*}:��t�,7sۦɝqx�u�ȑ[ulg&�MH��(�X����.s�f�� X��� ķF+4��=���o��� �ZA��5e?�Bн�(U�H��ߖ¸��^�ێJ
c�:^����.S���J�О��q�@r�\i� ��c���kŧ����Oo&��GSܽ�`�R��`��`���	4X�w�|Slhgxu�3����d�V.X�u�2����?����˺��!���b��XJ�����8�;^��:j�M�q���o��9��e�öI��/�Am��8y�{S]_�H��+��? Ĝ��z�zc�}>�/�4���㛺����v�-=V]%�P`P����PI	_l��h�=���OS+ζo#��c�{�<��[�&�xצ�{�|�Н��b@���4w1���ڍ�5{=�:[��t^@u�Z��w�Ww�8vn<�Һ�S6p����������D_��������'2�m�-���Ф�K�V��O���m^ܷͅ�؞��J��_n�����m�{��k�Ǫq�s��G��~��>p�z�����ut3ѷ�<���6�.&/_z��\���:t�R��ӧW'o8Ԯ�p�'�
�S�
T�{a1W�2+����=��P�}��1�>i�V2�}���/=�wƈ+�R	!�7`�W��'�t�Ź:J/���t.p􍠶i�hi�X�U}���sBXN�ւ�0�G�"v�����G6-��q��Tgǡ�]	=Ξ�>�1QW��y\3�����}�C�\,uy����S���Ѷ/��N��}���j�4<æ�h���˞|r�����f�3D��Q���×pr�� �����C�.J뺈����HkR+���ݧr�S%D�`��9�{�g�)��7�u����m����p�C�y���v�?��ʸ�̔�\�u��/�r22E���k�٦	�%�ly�$�@ǖw�X���ć,�9��*�/�0o�&�}Q���`:�_���9�f��̙'f�I�jg<h�!������XG���� ��y�[6w�8�S�JD�O=��81Q�U�7#�jg���/���h��g���kg�����a��$���ßc"c��><�  `��!S8��y�����.Xi��g;�t�˄�XT��h��,nq5Q.�x��(���43u
-�/mRh�z��?�@��w�w���D$�:	��}�g~֪��/͐������}Ӟ�8׋,4���N��w�q/m����á�n����3w��)W�T�R�J�*@�O�qA��1]a��d4�m�xl�:�S��E�54|�нĎb�`x�Ʈ@�U�ϱ��i�:o�oV-��݆�(5��^s
%*�t��`1P�\3g��?U�#O�u�>���`+�aO���n]�;��Dgq�#aN��>��tf�q�/�Fg����l��c�:U�qY~�{������3�UU�q�9=�o0Kȷ Th�w�b"%:�m�ᕎ�=�.�'H}��x���\�����{vt�X�����M��؆���!�^<Ǧ��.�7]w^�v3w���J7[�p���=�}�_yV�qx%�L�k��Ώ>�P� ��2�2ZE�z�1M��=쓰q�(�ʎ�C�ϝ�!:9W�0�
�t�S��^_�5��=������l�5�T�1��ݡ�t�u��}ia�y�~�{ֈ�I�n�Ƣ�~D�ʹ�=���K�~��	,kgO����3��8�]%�̯c[��^�ل�P�ZVz�% �&�_ 0��
�\u�����]�*eޗ�Sku�0����Y��g��wBOm�冣q:�^��0mgl�տb?<�8S��cޮ�mw�TA��B�4�X�L�?K�䕍9�g,��x.5�)���H��u]z�W�� MC��Z��EX�7�Y4체^�I��tb}7��O��*������G���u��m�ON?�;�q�^����X�o_l�qP�L+uQ#RUL��W
��_��~�:t�R��ӧB� �G��h�������->������n�L8L���4�ħ��	Ԥ��.��v�^�4��]����4p
G�0&A����\����ä"NHw|�#8_�z$�i�e�jsphz���������k��(�~�:>^d[�ZDx�� 8��6�+>�Gڠ}�L���mgü[���c�V:ø��v����=,_��>
|����֥�~��)��YE�uSp.m�ǣ[z�$�1O����La�.5����
?s�TD�i�f���f�[Z�9���ޔ	m�qDc��;��B��xC�R�je_��mgEY]��d-����^{:�X�נfPLkن�'�)e
���9����9��ySy�'�xgТ۱f]=�{����9b���7C�\�/��Ûtp�ff�d��� �J��\�2!����He��N�:~��[l�a_)kp!����V�yG�8�F�n���#��.��]�E���Ӓg�Vp~�˕�u�z�ר����R܏U�YD�����8=lz�����O��	R�++����M̾ˎ�'~#6����a�oG�}P~�ZL�=�/1՛>'�!n�0�! �"�\�z�dŲ{�&gz�u�s�E9.\���U����>��ӁY���[�|(��T�l���s��g v�J�*�:t�G�� 4O%մ�XrO�<�a���MyZ�)��M���B׶��^<�Lp��!0�7\廼�V�����L�E��4�8�����}nЙW�t�5s�Kp�A����90�;��#+������v^�z֘,5�_:�POR��k���z�G�X��I��uR�Ł��{~��(����0���PHfe;��3��� ��A�=�"s��^������"\Cl2��%Զ����7�&*!	p��=+�Wz������<^��wU�d�K=�I��!��_]KT�ٜ���`���K1oq�^�1�V������������Z-n!n�����mlo���­��p������0�V�o�>]<�`�hC���3�8Y^��MK�=6z�V�+�Qg�j�;ŷz��d�{��WΖ��w�O�G�D�}�c���KD0��.IrM7ϕ6�GFrn�9�?k�V<���2'j9���|9�$J�w��x9P���g��[Ȁ��d����wЯ|{J��y S@(�a|�Lz�=3���H�x!��/8fH��l���b��|�Xǂ>�aq�ٚOsb#����qE^�V�����8,�|���k^���:�c�o�Xl�vK4�ƅ�5K�g+\�}ZD�{w$�y.��Z�{w�c�����rB���|L���$VwĬ��,�.��uZ�u����(ٚO@�3\��j�&ܹ��K�����9;xe=�sD6D�*Q8��f�F�-oz��7Q�Ev^���z��Џ.�
��1�:��׺������Oo5�E���N�E�;�*&̒���_�eeJ+]J۾�v-c�7�yL�L���4;�x�5η�QV+G8�zI�{b��N�q�3�Y3�[�����<t��ȱ�7�r�<��Ӹ�A���Xs���i>AZ�kS��8�{{�l��z�����L��{��;��+�OEe��෽�H�r�.�:�Vrjmx���ż����{�ҍ�3�=N>l�dr�L12�+�r}��DKئ�.��i�5ol�Gז����GX\|yQ�0�z�3�� C���:RÆ�.実o7����kww�}�kh��̱8㳑�ql���L��T�*���6GYI���p㳷 �hlPZ�����a�:����F�˝�2i^�{z;=���Szrf�`ō�U�����N��*��bt�woq�Ν�V�X1r��ZY�S���Y��'^Z���\�U(��H��L��Y��a���Bq��w�b6�^E�(�kIK7$��o���":��ӯ�m�O���%�~S�Ị�`,S�ć�w��/%��	�!��`��JjXb|��hw��+������v��]��i�ރ.X�|��c�*|�f��Y��q���g��^�X=�-y�՜x5�'��V_�m�7Y��~+W�X��^`K���w�_9�Z���RID0.���U5����7���,��Qq��#Ǽ؏y��7����i�<V{+t��FvL��C���5��l��I'�T��'"�q�Y�f�Իڹ�m\��i���)�P\;ӻ�s�8Qx���a��}G@D���L�fLg�.� {���ӝ<V�\�h�"q;'��!�S�����n�����Ls�)��ЌQ��B#�ݯ�V���yoi�܋�q��F��9ܾ�g��&�݇;�LsvI��3,7gy���EK5��3�>g����XunO��.6*J�Z�ûw��T�&��}�t���u��/��M��>v��fc�w�E>���z�u�RŖ�>�����a�w곷O;�!w(�ڇe�/���({\�6oj���h�=�s^����wL�����w�w�w{�ϯ��z�aLQi�YLd0Fb�%��4D�i1D����oo�����^;kZ��n�=;v����� ��wr$,�A1=�d�fh1i2��έ�YՖ�k�N���N�k־5�Zָֻv��o<l�l�g69�F�4��s&
614��d�"��oR�,�Y�N�Ƶ�k���q�v���n�<x���өb���m��+���>.Qb��b$(����v��w��kXֵ�5�ݻx��Ǐ$�I��~����hĖ��0|\��n�bMv�rf{��	6M���*F��錐Tzs"�|�B_6�s%���*#f�9�����&MI1�)��)��k���U�D�4E2�l��c@�n���t��6K/��d��n)�+�>w|�0�JF�4m�i53M�^�EE)��ݺi%�Q̡$��o�W9Ml�n,_^Q��C1vw��{5r�x]u�d���Et*C� ��F���/pƯ�Ύ�y6�����ӧN�������u&����1����3P�0!���|�(ӊ�y�r�J�б6W�rʧ��,�v7W{�Y�v8�����W�>q]b�O��Rl����9���_����4dIu��W���V`o �}ٳ���(���"x	�Iǆ�^��逷{��G<'S��"�f��<�ڳ��!��g�vׂ������P���涱��kca��0�G�tCc*č�|̉�;�7m�ub��n���#���>T�p[鮑;==�+�(d	�Ԙ��ӿ����퉦AЯ2��=y���
p�\z��$7��Cey@��z�->�a�;������O���^�e�ۊ�Kw"��7{�n�P����i/�%��c�\7y��Tv9��9�_+y�K��}}�':|o���A����.+��D0=�;G�e//�[ʀ���0%��e5ss�A��E���6g9'^f[�*�pUR3^���gO�!���!�?'�}lM�6upr��N��������pc�w=�3,)�δ��*��r<������.w�����ne�������I|�_C���(��N[��%�x9���1���*�s�J�Y�.U��M����Qx��<]�C����(�$��ƝZ�Š���U��}Cj��Z�,ޛ�P�_�:tçN��N�3@����g���Q��ާ��Mc�
�O�{�]{�8+׌0B8�Inm:bм<��Y���Ǎ�K�gR��3�p��WQ�遳�]�}^xwі�Y�LJ�`L3&���>�}*�����+���L�5A�0����{��>����~¹`#�j��������ִ���T�[���z��x��������f�/MQ��<*��'G�s������4���S��<#�!;�%�KnvM^p;
/�a�:�R&C_�oX¾S��8AU�4~м�2���\;Vy�r<u��3G<�&k�����'�~�g�=A�BDLc��_}��M�ϷZŸ������J|�� ������l|����_E9�3�&�o��A��r�{�B�ʤ��S:1�lj�9n(p�yB��>}����
��>���s^@�"�}�|j�MV��.R;:g���l�/7-Һ�*W�w:��Z.}ʵ�!�&t�h��W���i`GD{�����ω�m�V���qɹȞ�|��"r���%0�G\(�ysCb��W�+�����(�|�/�^���EN�gas���4�����;�j���C-yڦ�"L�u&F/��.�^�-u��#n\��I��#3�V�\\$O>�LOrfK�3���g�h�1蘵�D~9�9��Z���K��"$ݽ�e�YsL�ª5��
��%1�h�A��N�IH�*M(�$�k��T�R�J�*U��9���wwټ~̇�}��32��?k*t���2Q��Q���̥���A��x�	�>����Yݢp�^q�辵�w���%��DI�K"�ζ�\��$J�9^c��3AÉ="s�������ѓӏT����,+�"=�5���X`	����J-5(�XB���,���ٻ����(v�an���6����TN��o9�xI�_��3��^�oSfKl��xY�.O^$A���a�@������ĉvn�]<��/�d��q���uw<�kPP��T�u�w.��ܬ��J��M��;�s lw]a1���B5�q�~��YI&/��9�r�^r�����]�܌�ʊ�猨�*D�2u�(�{��^Z��9��7�>k��Ur�;Mռ��٪��#y3�@:�w���J��8�3��n�`1�t<�����
�s�ֻߣ:bQ9���M�N��y��w�o6��L�t�qD��+?��J֘ c�=�F>o���Y�J�Z_��b���L�I�P�ŝ�����1�E*D���ꬿ5�/�R���u5p��Un���~�F��1�"���w�6]���*�ƪ����q������E�8�/�&�)�d<���x���z^���'��ӲJWғ�D�]��oP0V��V����7����p]���8Is�݁���؍�վs:��뮨�N�vww�[���Ё���*T�R�J�*�=��y�Ͻ��5�<5��"Ҕ�͵�dE�c�B�^�L�@��4�UT
��!β�G���}�����]?��fwbSS��˯���Ǿ��^,\���>�s�n<���S��3���f�cq�����V8���k��XT���.1����
'��w�s�<g��QZ�
��:z�R�6��}�7D��I��tWW�C�=�p��&�[�`(1�f�ۘEf5���S�,�rI���=�:{^ByɄ���aW��	��=����WĐM��^yF*E�ռ]afn����GR��8g��Y�7s���N�	<��Z�tCYa�
Z�ǚX	�J�w{h�fd�X�4�u>����G�#�갃/N�o��W�|GO3 L�ޮ񨵱l���1/���Q1[,VLw�e>�������Q�����?�@a[�LKgUS
�fꌒ����ϩA�Tt>k"_�Z�7��y��u �����
�6z:�/񪾷k��7��m[@�ɳ�p�=�O]�>����I�j�����wgq�By=}l�Uu����ϙ�;:�j|g7q��X��%t��9��`�5ʂ��ʿպ�BZ(���R���}Yu[G|�t�]���;��a��Q ��^S�)����]�Z�FcK�5���r�f�a��������o�N�g[}s����'�'s�����שR�J�*T�^��E~4���F��}`|��i$@X���v�x�	 p����\C������'����U�����%�*$�3(����>��G�<F��cEWkf���)�)��ug�p�B���>��Ե��6Uΰ�sg�9�h� �А���F�ϡ�@�{������χ]1)��0��a���>|�&�Q���+#D�oE0M�W���a�q�\�-/%��o{��i�l2�d���9�|'&Ϛ������z*����Q�|`�\���L�����UD��4�9�67oD�גS�(#�)�׵ـqO<�IG�P<@p*p������C��(ȗ��{����%I��n~�&Ux�2�)P��'�/l��{�fi3�3D�/<��1�T��+�a��B8�;5cP��j�mxN�G����<�Ϲq���qV��E��5t֓';>��r
�k�����]#:�纏O���hߞ�x�}[�2��F{�[� =���v+��u�ÈQ�z�H�'�s�9jb��=���f�������]�5��L�В}�ƈ7�Qy�-m��v���R�҉ko����;+D��w#���sx[vc��/�g{gb���V��;U�eUa�k�
I����9����q�;):��G0J���F���Nv﫷¦l�^�J��:T�Sf���d�:	���b�O����E0����{@��q���3=�����o��D<ͨ�W*��6g;�䣋�qg	�)\XQb�>!p�O���9W���~j�my��ym�Ĉ`]�f�a�N0f�
m�MW\}�v�{=^���t9
�`�����G�u��UĊjq}�l�nq�T���g5f���1h��v=Ɂ�����ޞ�pf��˒Μ)�SC?Ww�ܫ��/�d�ο��R�o�A���������I��+��e�k(G%6.H2�dfg�c�S1TF� f�f�+��s�{i��+���B�q�0�>��.�ݪ�u՛&r$Y�< �����D@�I�9��5sr��fU4��gۮ�Ƽ�Ӥ�\w)��Ǜj033Z�e���fHt��{v�����u�ޯ&}�T{v�p��z˚���|Mz�\���gP��Sܐ�n���}�����7������[�*5[���K"���Շ4���R8!Բh��͸tqt�?k�	o��Y�	��h�";�%�8�D��w$��>\�ܫ��^>Vz;�;���]V��j��썓�Z2�=�ӡժlίM�V��]������� Q@���G!f"dF�
�D�R�)��E�Ce�^�J�*T�R�E��0#�h�9�C3L6��v�3�u�xUoO�y���gٝS]��	H�U`�o�[Z��n�k�#��e�!t}o����QV���η�6�\���*��څT����^J�ǎ�kڥ"�Wq�'4N�������w�Qk�j�՛� 1i���>�������K�GD�Mn�K��k�gk,X䠔�C{�j�h�o�nc����Q��ζ��Wni�~U"�Q'�a�^���;��3y��m��`���K��W�f�����La�Q{���oD���W����7��L��n乯5V��j�
p���3p�Ϫ�;��,��s\��۳�����m������s{�ff\M�
�+�K|��l׋���O�u����5��{�E���g1�R��Dm�Ed+�eN����z�lv��<������G�J����� ��)�e�;��sCӶaQEB��#\�0��UΨ�s�˗�=��lY�_�<L�K.g�digߓ�@�=�>�e��$4U�63�2���U<f^��v�p�LK�K9��C{�u%�ºy��m���c |����~?������%j�JǼ��{�����m�vF�W�G(x�Q�|�J��ηo�ɉ�ۭ��WQC<pH�/R/s�Лo=[,�#Q�Kz�zgg�����$��1tVR@RXU��4'���l�{
�ར�n�L�� n�|N�H���fp��jS���d�W=�*�������G�ޕ�P��3{/Q�1�^2D��˛�ӹ��h^]�K�!R��������F�"�`�8W�?0����g�Ҿrp8��L��Z�Ү�^�٫��tM3����w�͞�^ճ����tVZ=V�_q'd1�U���J=� Ǧ|]��~�)�}�*f�J�V9���c#���`�]@�%@c t���%�&}�J���p��y�ie��X�ga�(sϔ�l9a���*;�;�j{�f��m��v"84\C=�X�Ƿ6I�'��}9L�df�͡��CG����ϯ�L�����#��L��z�e�-HNuQ��{~S8]�o��N;/(5����;=�{gc�뛪	{�U�}-�����a����כy`/~�J�:t�T�Tߧ����z��y�����Caߓ�34��9;}��}큇���Kr��yYm؞NQ���K�
��-b�u�Vg��R"3�==�ԍ��1���xud�ͼ���0�u�7#+�Amo;y��@��N;MF �(��Oq.�f3�%��J�O�45t�F<��l��3Y���2�Ƿ�d���a��C��̥��_A���D��hk=J�]���wxN�О��y�c��"��C�oWn��7-��zY��v�9�<��Cط���g�I�vf�B���x(}~���:�5��MGdD�duC����"���}<Ii��-��hǰo!^�n6�}�V�{�g]���Lw�Q(�#��\����(����l��=�x�γ����螾���i�6�*l��/AH��W0�T/POV�����gi����aHIY�r*%֎2��h\�=��Y�����zhC(�.m#�f�{u@n�)�\�`�]�"u�ٓ7�lJ�[M+֏���#߁�Ш�	 ���T>l���lަ>ʕy7>�����������{�^4ȶ_k��V�ٽ�NQ�����گ�;��'�kԩR�J�*T���o>���9��q��x�,��h�gz�7_���7s�o4�)ݰ
����(杙@��Rx�nR9!�
=�|ùD�B�YOPn��p6K���*�wy�����d&A�@�I>�a��������\k͇�6߫��Ww���ep\�8�b�J��� ��/��3(=����dA�p��]�����Ua���f�X�nT��L+�M�[|qc��#=!O�C��'�.���3Yq~�� ־�����Ir=��H�M���q�5�K��k����މ;@�mu<[��Q}�=˛�T,&ү7���/��;�_�����(�*�lӧ�%*ݔ�9Q��>�4�۷� &��7�C�@ق��`�1��Q1����M��n��/�*o���1K�\��#),�0�M11�]n�{���fݕ��*�q�3��s[^�����dW-�L���4����b���R�pI�#�J{_Og`�b���ǂ;���ro�*5蹲]]��*p�G4��AY��+�xc��Վ7�,dv�ܺ�8q�9yQ�]����s/��ǳz�͘�v!������s��*o �v�AO�I��ns�ú��N�j��c!3�`�o{L����$5 �/�8���;�N��8V�ݛvk�P�ܦ�1�W7�7�����jB��:櫬꺳r�PD��|��.�ۛA�|���Vѝ���(��ݾ��L n�8ma4:qw^�ݶ�oB͸&> ���LKΆ���{#7��+'=U���=";z���pɯ(��9�xtO��������CL�j�?b��U*��J�G��B�V)p[�¥Z�	��
9�3v;7��7,��QQ�0��+䯛���t<�K��m:]9��=��$��o%��]z�:��R�z���q3�h��U-*��W�-E�����i�`��@v)��|�yb��$ ���=�.]Z��P�);Bڄ��S�eX<)�m����*V&�e�7��J�zCŴ��e�%s݈SFk��;��i�r���q����F7Svm��7*���q�F���y�\��Mx�̿�W\��I�#d V�_>�\�jSN�;w�7�Y�8���k��,�0����(sa�CF����2
�B����U�~��\�o��w�,�$��B�\�����j�F�[CK,!I��.�%�'�P�P>��/H�T�8(�E�#2�!x�-�y1����`�}}�g28�RO�In��v�-���N�[�����;{�:;�y�Xyf�b�l3a��w�z��e��g6�����Y�L��U:m��זsb�K
W(z�
���jCu�g
m����wp$�u�{��r\��;��[g�~����@����������w����=#�����_\���ʩ��J_]�g^�	�74�2���29�,��s���$t���NG�v<O�/�6����v.��]뽂��.❍�|�X(�Ԩn����Y}�4e'�Ĵjy~��8�ө�L ��d�v���Z�1sz3$�9��0��b�A�.ګ�)��r��6��]�}���M����]�y���)M(����m�J�;{R��쫓��K;��nuK7��M/6�}��[L^R��W��<T����X����8�Sq���T۬rV:}��j9��t�O����#�k��'�X��(����e�_eC�Ch��R	y�'{�^Q��c���׵�=�7B�6C�z�w)�+oY�{�*-�[�3��L.#�����w^�[�G��/�|�!a�Ep��M���E����d4��&Yj7E�I8�A��+�x0+��%��-��( ҂&nJQ�:�l�[i��$�"�hcXlKk� ֢Y"�iABA�	��6���Y�{�%6X�daEL8He�%������,��$���A"����$тM���ڢ
(���(���VLWN1㷦�<cZֵ�v�����Ǐ6�,��e��,�e!F|����_=� ��@Bl@�s/.���a%��]8���ֱ�kZƻv���o<|��]-���Z�Y|�Զ[`l��np��
�e�UU�oJ��ǎ�ֵ�kZ�5۷n�;x��[d��[l��HH�����D�"	ѷ�n��<vֵ�kZֱ�ݻv��Ǐ?���E�&;��H�6wn�X<�ɐ�&2jM=�69�#W�����D1&�$HDJ>��h1Id�d���R`(�� *Q��Hd�4Yb5)�d��HQo�rF#}�2B��Z"33_]m���IRj$�2�wL؅,b�-�Ta(Ɇ H$�$
4@&�^o�ّ�4�Q�Q	�"��A��٧:V�\rE8R�2��[�%�A���Ί�j�uöcOMd�i}u �[��B{�=Ȉ+A'�*E�Y�0\ ��B#i
��m(Ҍ$���kk�T�R�J�*UvF�����s��J<���\d��p�tཇ��j��7w� � m�3$q��`ޚ{ܳ�7�q����!J�H���0Z���ȕ�M7)���7SGw�Ka�)V�x�g�{��ٲ�:46�3�٦�s���\c; �`P*�tXy���;�aC��2�"�g~��~�E���=�r6��(���#ǽi�]�x�^���3{���;�i9��}2�Uk�ԙtm��������r�����[;���ۯJ��Mxr��ѹ4W�k��G��aB:������P����rtyI �
V�2vMoǧRK[kh���[�\ ����1z�#"����9ʶ��;;;O�h��$6ǻ�UhG}��a���n8�0��U�2��N����R�-}[�鵪BU�ݞ ��p��0wS>��@lk��0��^8���I�Gz�T�����L�է��o0"����T���'c;O�R]�?U�h��"J3��fL%�V�ͺ�
1�1�9�������Y*���0?fK�{7ԣ��+`��;��K@boq�z.�O�������?�������[ؾw["�(�n�ǯ��Ǧz���^�d^2�1�yx5�`����C;y�;{�Ѓ�"����`Vtw8K|Z��W3���b2%W^1QS��ϼ�7���T풧Xv��e#e��Ey^]1���i��CN��W�=��gql�7��8$.�UG�D���z��ZcX�Z��&\�_pw��o�X���:��w���|ǎ̫�[��:a��c�wB����A���y�l�p�q{G��#s��E�foC˽Q@��u���2z�)_�6f�����|��V�Yy{a6�Y�l�Wo-�rx���᪷����G��� /Hӳ�I�dI��g�n�����u+��X�6��W�G���� ����޼�� �/�Þ;���v��8m��d��
�@�u��tz�j�M���1<�xV�NED닻��Z��9I�]�g��� 5��\c
}�S��z%M_^�>�U"���jL2>ɱX��C��*h�S�G[S���O&��̘�h�Cg@��1�Oo\��T����ۛy�{W_�R�J�*T�R\;�I�ZA�װ��d��u���q���>�ۼ(1�A~A=�1�2G��Is���$�!&�Gh4��{讞�bK��n��p��c&�۪�aΒz=Ѕ���9ó4����>nzew�K;�;c^iG�p�6�#D&C�-?O<�5���`v��.���Td˳<ت��f�c2( U�H&��_Y�P9��;�Ɨ�n���t@�������v�����U��3E�]��ϗ^x��8�ô�F�$OK�0��1�=�r�}��UY���)�QZL�U��U�={�Z��,���o]���]QO(��AMA-wMz� ;ϳi}2���X�L���]S>�z��U2��`���_d
K5�;�H�H������b��Z��N�Y9G��p��WTou��I�D��@��V�h_�{C4���y�讎��� #o�Ƃ��A�ZN1>7׾W��!�VL��"ꈳ�<�]6�ޓC��-Mj�Bu�f-�t.�츧��}������x��ݏ#7��rI��#iשR�J�*T�S_)|��}&3���x/���`=P8�9�^��âF_��C�8�\���YݼҮ��dL����dy��A^j�@g��f*_�Y�i���K�F�у�g<�;��]�@��sciP(ʷ�y���e��A �(��L��# �s[�պMh���áetq&����8Q�.{�F^�0� ݽ��M3�[�����hCl�н�߫����)��܃���ke]4Z�2E�Ub��2#��}�d*��Q�j�TwOws��w;�a"�lN�]�{M���y��F���o7q�-����zm��=�����9����1s�����1O��ށ�d<�>���j�آx����gn�(4`������W&�̧:�=�ۣj�������?k��o<M�윣צ��oҜ�O��������*�:������=������$���Uf�ʩ{찣����6�.�3#����8P<�z��U����a�k������]A�A(ٍ"��l«^1%&s�ޢ2:>;:�e2I3
W�7	v7q�:��1�^j�1���2���k�v��7_{ݘ�H�2@�I�,�0�E&��۫��R�J�*T�R��a�&�QU�5����;4�=G�B������_�}�^ۖ�O�+�"���]�N�fq�kUM	���ѐ!���M��|��&�N���݃��=����D>�� ��{<�#��q�r@t�N��VjD>vB�
ӵf���53���I�3�	�����K�X�帽x	�i�*����eU"��8l����3�;�����.��`�؈j�K�mʞ��ʱ�#H��i}���B�y�=ɘ�!���FoV��~F�*ܛ�ׁ��p/ׂ�P��S�V��>�Xr��eu�D�����|X*_�boDNi�M�����T,!���ge���TnX�Þ��=�V��,�v������r���.��;grc&%�[36\[w;�g# �zճ�	^�����|�ָ���X#~�>���3��4�2��1���_ܴs�W���҄16���{t7���66�I���y���o��L6���rjo�wz_V����7�uC����t��̜���y�]*�*T�R�J��ߝ�{����w7�y��3�}#i�wE��ǜ��(��
����1���d���!�oJ.+���{��t�;�����Ml��,�ֶ��ǒ���'c�Kj��j�h���Q�����v�a�:��OD\�v��ocǽ�"��� $�v�_�ԛ�C��^|Ţ,�N��=X�����`�W)��D,މ��W��P�7�-���駆^�g<a�o;��| �H���^����EyW��ćX�Z����YiF���Wtgj���kCL�㏮�����~2��BޛV�wYJ��{;(j���w�Z���r׫�(=�ƇȈg���q�cP;��^k&���s���9��`�h�`�J��~��ٻ�JV1�|;ј��~��ʙ۞�o����,�����V��p����~���T��8�/^�6�o
�������D�{�Q�����nM<���;�[���$�{1�<���p�G�4x�^�?/M�}Ҹ��`��w)1�r����=���)6��}�4�ޝ���`��k7��9���w:���_�J�*T�R�J�����s��OR��T��_qg��$aP+)X���c)N�� +���]����B� Dx��}R�C�=�@	��xuWC�^T�۵��ڲ}�6�­�}p�ce��a��%`�T���j�g�>l)����8j�2�r�ދ�rW��U^�un��p�*���r`u����t��g�ҶZ
2!�;��^1ᑛh��C�<'�{j�m7M3�c�^�>���y͜�S�U$�<���Q��K��lܿX��66r�� ;o6�鱸|�x���uq��Rt�1��0V��~'6j�&�fv��y�N��3�4���v|��Ə,�o_q��������ʲj��y�����>H��A݋a�{�bY�Z��[� 	�����Ղ�v6�#}
Y�_�;fk�i�ro��z�/a�x'/�����f�[|�vF��t���#0Ș�k�ŵ�\�'2[!��jxq��=1�jpN�Uá���?�#\�����݇{�ޚ�I��&� ��;�p���7�ky�?/_��o�ꆣI�/l6x��?�������?���L�f�������Q=4:�ֻ���z�6����CN{���ys�r���r��kn->^5��{j�Elё�[}|ٛ��忤�ϑ��{��͋ �D�	�d��p�4����Z�wA�'`�d0(s�>^�Y��,��:�]gToގ�ka��ַٛy,܄u]�]Ըrrw#gJ|XiM��2Z�!�C��VߤF����OY�z�}�^[�%���{���Z���������d��
�l!ޙ���L�=u�+e�H��Q��ݳ����i�@WRD@��ƙh�c���9�|�&m���֦�fV���7��D��z;i� ��S�8r��6�m���37w	D��3�>�{W^/�ᇶw'�hR��2۽T��QQo����ǉ�W+��
��&#ա�ӗ�nt�꯮��{���3�ff+{�oē�|vY��d��(6��i��Mo�c�>�}�"*�����yk*D�"!ִ:}��V.:���f@UcL�[��v��B�ۓ��y�k�O�y�V c��mۈ�۝kL%N�L:,�1��E����G�U��&(�#M"Z�D%	h@!U��*T�R�J�*Wv�I�o������J	���RQ)x����0��S���x�U���i��w����jӛW��س�2�o�^AW�� /u`c`S�ios���'��hǜ���|Y�%>��̗�_䅲��j�rO�����,[��՘�Uֆf���b��1l���ao����O�z�;9ƨ��狥�;�?i��Z�q���Ex�u�zV�Яw����Y��O~��ol���_��cw3z����k�g��%E�|�ܟ�*5Jv�k�B��|�#Y���Wq��0G���a�t��]׍��h�ؗ�l�t�cn�v�n���;{�6��08���������͓�'k�ᓸ��;��f�E\�$�D�@�������倁�2��3������o���;�]Lj�������Ҽ���5d��v�
��{ХT_۞o�&Vֆq���{ %p�ro���a�R\����7��cC��MZ8����ָ�i�5" ��$�L�!I0&�TA�R<*R-Iݵ\0<%��Ve|9d�v}X`/�]�e.t!��9�d���P���x���ݺ���/*T�R�J�e���;��{5?��U���x�oJ����U����a�u<�|r�[��b�Y��Cc�9,͕O�0�0�+oG�J����}�әF2�iZmd�r��h���}1W)���w/�>ws�8+����zb�iKsw#���4�LB�E2U�M�թ�"7�srl�5
��o�3{���;���Y2p����2$[���s�o�<�8�rQ��6u�uy��g��-f���u|��zڹ�u��k{Zs&t���	wޠ��VX02v{M����ճ�l�+�-T����wh�;�J�0sؾ�g�\��p�5�u�dbM����SZ��=5"���{L�1A��`������<9���uA5���,މ��O�T��2bB�}�;�=�[B�SB($h׌��̏Wk��+��m@n�u{���v�Z��6�A0 �9����������;l�˖%$�Vr�����W2��6�6;^�B��X7Y��f���ɰ�S.��ڵJ�Z��Ŝ���hmΘ,�9�	���M����A�!������\�Az�l >��X���B����byr�/[�:[ї��F�-�P�ڳA�x�'{��mk�l�ݎ�||d��?d_6v!��dHYu��m��R9����n��S"�x.������i	��I쭉��W}��Bk�}�
Cyz�Rz@��x1b��x�Yj��1�|�&=W�q��Ѣ�^y<�';"�Wt��g�y��E����
�Z���d�k_*3]�������IWH�g����8�	b�&�[�N{I��`ͮb�=׽��n]�ˮ��p��ݚa���?�v��/���'�+V�vA�kFt�<���PX���[ĝ�Yoq�ӓ��f�f>���oEy^��p��RnO/gNY�Ou]g	&�۷|3���'��������twfMV�8m���MYZv�*v3~�NcK<�;���f���L��ɕ����.�=���\Y/7�mD����6h�[n���=�H����F�-��F�ӢOExw�؟��>}�v��Y�*����@�B�m���8
0H��m��:��q�Z9�V��I6ݚ9�1]����jR�_���?��"�����w����/��7ZoX��M��wSYw�7VI���u��d�O���jl�kY;������R"��Q�����0��Ʈp�Z�!#��=�Lc�3*���æ��wWq����v��|,Y8fd�[<��$����n��.a\<C^�XD�S����Es�AP$�
��{G/��器wP������E���ڲ�aG�=��u�ңw�R^�F�-��<�;�������ܼ�/g������]���kO�MՀ[�o�,��1v<��ޤ���ܤ�-�ss�snŦ`�Vg�=׮p�giv��i	�e�c�|G�]}������w�����~�·�sA��z�˅�+�N$[�E����eM�;~��1�x_.׏!�>���.��"���ZWg(ȣկe�]�ɗ;�⑋��p�ýv�7z����ؤ��4�)���k���q��о^6���_��+���G<e���ٝh�Ë�$lb����֞q�pU�Ѡ��f�-�MV�쪫�I���v�������Nq�'7�v{W��^���q�l'p#�g��n�wً̘W�	&� �	&0QC3AR�$�fQb4o��F�ꭾ+������ֵ�k�n�����w��ߜ�H�LX�B���^Acbɡ,��e�e�ղt��<x���Ƹֵ�k�nݻv��Ǎ�d�Ye��"�1o.P�e�$I!�ۆ#��F+�'U-�ӧO<x�ֵƵ�k]�v�۷�<j�6���-K,����3�߽���4G5ʒ����0�D��)�t��Ǐomk���k]�v�۷����w�~4i
0oƹ���6�1'�۰�$J�"A�ܾ]�V�Y�)��2�1f�M3�I������ܫDb幓W��d�b-��\�N��ر`řX/�r�QPb�TP��� [}u���W�_}��Ph$�I&�]�LA�-΢��B!E%��i�ך�����QK���@�'�⾊)����h�\ܽ�ĩ+:�_l��v��Y��a9�rj�����w�pL���5��8M���N�*T�R�����z�s�fs���>���Lη�3��E�I�H��u��:ҵ_������6li�7��'p�A���A�(Yl�n�ə���g*�3o�-6{�����8�F��iq�X�K}��T�n�8�A#���t٫ܭ;a�cY����{���5���=���� ��C�n5�˱����s�����U��	�%q&RU��i���|;q5&��_F⁝(HUu�.hGTvd��駺yu����,j��+�aj��D�6\w'j��J������o=>w���=��T����IMB\2lѧ�5��w���Vs�jzId�6�ji���S��2������dC3��XM��g�b5�#�=���;���L-�A�/�tU9��L��ͺ�¯N̨�"z�	��*�J��s9�,.�6"�m���PZ�Aze7-�?��Pg�񳿱���~�2<_N�y���\kv��;��@���V�mކ�����W�g�s�[vN)^��[zwr�Np�g�F��ગy_�������:w��mݍ�y�U��*T�R�J�*ǽ��ҳ8��u��g@��Q����z�����<�r�R���,%�q��z�u��S�O-��퍺������f��O۽��>��0HBBL�D�Gw����樔-���=�����&��q��wv5l�N��[��} )f��-��}�ݪ}�Σmp�j��j�b�NWq�ٙH���T��&�6n���7<b9m���{w���^)42y����N����a��(���9 P�nwvm�-�c�WX�&�܄�Z��6���Y>�ɝ�p�t(��h��C�j4��z����nhw�?'g��<B3�����s渉]��*BC�e���������C��S����"a�l��_=oL
"^�S���������� �=��Q6��5=r����+:�p��m����ci���4�h.U%H���)7�I��:(��oxmY�Gw�{��ht��.�u+�M�ʅ�ū1�h�R�
ؙ�=�j��ֳGL�Y��z���ȶ���
%����p��AwQ�g3���sIU:f��+���(a�J�1T�*�A%��!��1�U4Ґ�n��˶G)שR�J�*T�V��\�H��r��U40�ֈ��3읏M�b��-��R[�e�X��[�2!��S�M�y��ۣ�f���.��)O�1.����D�"���L�[ɧ��Z$O{;��>y��YdW���1<eP�~7��b�ۗ�vɣ%���Rͣs����<
cUbR��X���v[#U��3,�brmT���.Yw9Z�<��Ϸ����9��Y� ?�����8ZO����VQ�[�������F�{�a6�HVܽ�8%���~��\ʲ9*���ZsIG�H��oa|�����5�ez<8gFie��x38���K/Q��~����˩q9ɻ�C?�6G� 3j}��%�l,�Mk��ߵt����A3�e'|����2=��!^�J��'����"v�۹~'s�0|�OhO�����'z ��N�V�����j�3�����à�
OW\�v<�Ykl0�5on�!���P�I�h�]c��j<2�ou���h6,D�X�.%��IM^�>��0L�y�9��t��읡j�0�;�xK��Oڼ�~��ho�CË��]�6�x]z�*T�R��R��~�w����ȩ�+Ի����(�-�ٔUv�k��l��ո����[��Tf�N��i�:5��ѭ��t�Ʈ����mwۭ�/s�s}]���:o�F3�R6����	�/b��ɡ�"�TEFVm�<_s6=��-۝s��VV4�xm�a���Jj*VVN�I�;OT���vn[���ޤ'������낞�J2_���`�,�k�U=B8��p�f�\�����������U�|���e���>�Q1(K��h�
w�v��c|S����c��н鑖wn�z�>[�mֆ�;�{���������xL��݈�
Uj�gEԸ�=e���[9�ُ���m&mo%�c���������F�t�-����Uv�p5�o����(&C���6�Hק��\�ֿ������J��|z�z�Ϟ������C/	ܳ�,�鷳v�5'#w��ƃ�Dv�h�be����[<W�o_u���z�> p�����Ƞ|.7�*U�A��yi�5�s�J��r�e�u�}J�)�f���x{fc}����5���E��W�R�J�*T��w�߹Ϸ��`!��6���Oltj�P/=��WOj�>,q�m>ƻe�Շ��9��p2w�0��S�B$zzϻ���r�U�L�K�����da��^I�6�aN���"��S#w�,ދ�|���tSE��ǭ�gi�f2���a�\�gVTK�	�c3j_w9�L����6l�Lȇx�M�-&����lϲ�X/i�P橿?��n7���d;��z�~���Xt�G�	� ��c$�����L�x��J~�����'�uI�8�b�
�gݙ:6�d���2�k�Lj�SlZ_w{��9�H�?���Ѩ���hݑs淖���7��'`���l��5�95���}��o������j���V'���.�7����F�bN-7H��L��)��i;`�5W,��]38wsB)�ݼ�Lҧ]S)�O�<���[�A̛�]Pw4k���`�;˭
��j͵M�N��₅޵���9��č)�LmS�{%�+z����d�c̾]��E]�<��r�=�����}֋�s�,�wz�78��=����������t(�7
3Gz��ݦ��>"���<�c�.�TT�i	g��gMp��ݞ��X�}���~ԕ�۹�M8
h7P:�<zT0���A�	�+x��htnG �����5ƙ��V��u���oZU*+íX��8�V�GSk�.z8�{��2u�ا;�5�N*�����Lz�ƃ���'��HߖL�˲��c�֘��+�����6�v��œ΢{|f�C�׊&V��[��yj}F7[5���#����'g�V�
.��g]GL�ʹs���p�{��'�=�" W����6wi��=�W�͸�Vۧ�r�؀��|= �RJ�hfrG0��u3RWH�2ؽ4��g%SB����}J��٭��˷�+��V��u�;�7m�eHǡnq��s��h��X���=?֚7ٓԾwcy`.�>��O����4]�����D�4�6e�3�$�kYG���l�g\�4o�aΘ/�n�S�;��n���;�<'��}��y>�u�ϼܯz���)���9QZ=���xb��R�	$�B��"�EW�R�J�*T��X"���ow��q[�B`�@gSx< ��ˬ�:��,ָ�n��N�U�(&���nwFuZ�D����(3�z�o�˹x`�<X����i������3�k�}t&o�'��>�]J��u�w�K��=��&5���b9�I�z�prp8�+_l`kޙ?�z^﹢3Z�Ygm��z�O`{c!e�4���Š�������{>�F�[0ff�4�	D=Yٸ'
�^�����y����X	7^V�Ǯ%z�%q���찛L�,Fv�B�GG��\�;� �GG}Jĥ3�P\��[���~��M6��PP�@��D��V��H�^�Tg��7V������fww�q�탦P�Y(��>Q"=pJ��Uf{v�y�F���6�`'+��ێ�y:�T�*@H�4q�޽#n�I����J~�>���}rK����;Hb�OU�*��vm[���%�5�oOc?Wx�,�d�K]�U�ݤ�E�gZ��c1��"�XC
=\�wٻo���6��E1-L�ǣ�� �����`X�=̶������!�uh��g/����+�*T�R�J� .�h�t������d�4ǡf�v�`���\�͆s�/V�*�l�l�h��<�p�J�tD�^O�Ou���q&'`��eg=�U?]Zw���عV"��z��};b���q���zhub�oy���M7��՜T�C/�{5t�)��}��zmOK�@p������"%ȗ
5m֣�z�f=���q��m`���{�\�c���@\W,�w��/3�Rv_w:�^�r���� <���`,�8�Z����euӕ�̫�h����&�ơM,��Dǆ�T r�ґ�w���ݧ�q��{����<Á�������_i�ݕ~����v������)~oW�\�}�j���v�T+��%���i�o�^MM���R�(JZ"���f�d7V>�'��)3=O���w�MUϫ�aG��l�;��ʚ������X���˲RX6}�(�7�T=l�s�C�5�㼺����qh��<����;�p]�$�״����KX�۽���)��{�"6B3Z�f����y�[�L�ܶ�����*T�R��R�����Xsb۪��%�9�>�((!׷һ�Y{��d��0�˱�)�(��T�p�ħj	�j��<M7^�6�P�Vþ<��Q�ʞ�7�Ӿ����˜ک�gp���|v۫ҫ�sv��h6	-���q'9���o�>��t�z:�6Ԍ�r[���R�/^�N�����niݝ��A�3�F3�s��\���I1��췻M���8��#fw5flg��gt�#��j�=��ٙ�1�ݖ0�J#8`Y�7+[�$���]Z���Z�mL�ѣD��Rݏ֛��;�Z��bet��n�vQ��h\T�D�����嗑�W���5�;y���ʶ|j��5�`�ȃ����wWΠ���oJH��+Ԓ)�n��r}���l!�����|b��=m�xU�澝�Ѷ���9���������P�p��t7��:��Y�Yq���*u�R��N|�k9wV<�o+v��0�??h��y]���l����.th����2��<"��M����V���X�,��t�<&�|��&'���sr�f�����n��'��ǏO{�sl�p��W�R�J�*T��o;�A����f��ؾ�wff����4M����j}�hL8Gu���;��^>�c��i��O�:�(Cj��cv�1�4H�ڑ�{�˄���aLu��m���͜��Z�R�a��^������$YW��M\����ؑ��\�\"�'��ܔ�)1T/;�+gb�CW�߶�v��oP�--��
�9/';7n-mi���aB=�Q;Q��y��C,��A�p8S�C���ֻd�D������#�o=�L��r�P���r��Kz����'�L8s�{���lm+�%n�6�d��pwQWdmnBTɭMЬVʜ�uT��Y�����WuZ"t�:1��z8��<�9sϳ�q���^�
�!�(���j'�λ�V*�f�۳� ��y�)�5���@#dwC0h���,E����@�9���O�QN�s���g�l����;V,�W����lΣ#���po�.1�v�Pś������|nm�f��˵�N�y��d��=���n>�m�q�ݠe��ZVF��3�����gB6�i	��������f򸓸OU4wd����`c�J
�C!z՜��%*����<Y����A���g���{3����Ǒ�$s�k6,c�\�YFw[�Tv/�2��BG�:�-7�WN��z�d�k�*s���]��	xJ�NɚV�n��&�#�
�|�rHu&:��\��^��#��Dxy�D*��	�{�'�rvl�\���^Q�;ˇ#O��<ޅf�2�
������\�7A+{�or����Bi���q�Ź������|�ȉ���GY�->��!�U��f�c9&�
&��U񪞬���wj���?h�Qۆ�Oj*G!���� �˗�$��\;���˛K#t���sw ���}��v&�g5�`zǧ���u���F�]�s��|�wرi}��/��a�>s�1ա�A�Qh�k�\���PUH� ��e��\E'�1�eܤSν��@3}|TK=��,f\��i0��hԃt���P���4�������.�S%�Α�QD�|R%�J8f�w-ABuf[w�e��LJ!d2�2S�����3$�[h�y��x/ap��'5�Fd|�p�k�q$F��r42��b�Ñ���S�V(=|�s.4�qmu�������"l�ɯi�z��~NlY��ǐ*%ȟH�p�5գ;�8�m���O l���fЫ���ê�s(	
�7��VK���
c� `G`�;^����'hn��]իC�F�F-;Ld�4�ʋ�vÝ+P��t�O��#Ӕ��˷��=7� ��[�j's�T��K�9'��G׼3:�M���>�ޫ�L��<��
�.�=�wS��e��W#�B��4VS�X{Eٹ;s��r��Ǹ�b�2±Ҙ(�|낈wA��mݾ �^�9�˅���aÇO�J�Q<��-�z{.�-��w��Ͻ��p�% Dwڭ��.A�)��D[3�Ѧ�d<;��fh�Ш��L��튬p�rg��q����H��3��4�1��p�h�r�M��>y�5�2����]'>�fi.���z���$꺚�60���b�
����.��2��v��o�|�����)�,��'|f��J����Ꚁ�����֭N@ԵWC˭��z��@pe:�޾�܃T�w�u=q���-�V���q���3�eXó�o���/�v�k��iz���n��j�V�b5-CD�9�	�X� �10�A )1$E#�:!��8�c�Pwb�rY�i��r�P�$���q��a��$(�KD�PMZ��p��V�5dH�7T�m��4eQUI�*�KWQԢg��Ϟ��|��_j1���Bh�c���DX��r��g�$�O:v�=���ֵ�v�۷n�o<l|�Ԗ�����m� i(��lk?\�t�%�l�q�Ǎ{k]5�kZ�۷nݵ�ǍI�Kb��]KmU���h*��(�X��m�ܳ��t��Ǐ��kZ�nݻv�<k}N���9z��[zd�X��m�bKe�K(�:��vǏ�m|j��kZ�۷nݵ�Ǐ<�ʖ��KU�g�}j�F���&ѽݣk-�]��ƾ��^F(�^n@cc1n\ۚ��E��ME�Tgu_�ѱ�h�#Ee/*��Г�k���j[��ҹ����EQ�-�S�k��W��Z5�F)*#k��/�4&O���WN�>��� `d�I8�E�ug�ɋX~�ޗ-��q�7�x��O��͝7�ΊI�ɮ�gOV�����/Q\+ԡ��"��E� >|��%�"�Q4�'$�*�-��%�yJ���R�J�*T�� �>_��߬	}	@�����-gZ�ڟp#;�����F�� .�����d�Uq�̔\w�֫���u_D���M%�6�/�pu�|���y겞�6��tcIB#�{5��{��=4:��f�evx���19��ƭ���g`�z�.�u �����J��<{�����e�{�5�M�w1���?�y��������+0`���f�h:������}��&�7���	lЁ�����F�ba�X1��Ӹ���"n�u,�i�3|��0�c�F��������&��=q���'y�f����wvOL�dw���'�<4:�*A�phho`19����*Y�Vh%����,.���'�L{}X| ���mW�-d�.�����gn���T9
���N���ui.iO��j�7�e��O����o!����$t/l�6�����`�=�(��7i�=�oz�>0?;��n�S���v�Qs��ᗂ�Bk7�u௽Fmi� Y��f��|�k^��S�.�� ��n���+l���'b�����R�����7�����)-�k$Ӟ!�������z7p�`{dM�Q�t���G4�ndyw;���S�s��+����m�������W�K���P�/v��tχwuW�on_��L����r/V֓	��˾\�d�-�}�A��A�RG�֊�9n8+���P+�2���xvj:�B8��_g����ff���=�_$�O$��y��\:b��W�Ҳ�/Ba�}��^��^���&��w.'92fq;8�ߺ��4yo���t�H��.N�򟷞�%[�~�[���omb�����M*�p��c�X�s��y�ur�/͗�A[ùX���
S���s�����M�ۗ���r�*�{8�;9{[���a�so\�d�/E�;vjXd٠c��	u=�n5%���}�c�է���*��~ȿ��Y�c��H��T!u������v�6�nj���ٯ9�f���n>wGE���N>����WZs�\�SW:�o���p��� ��ope��'��E	���I\�dX��B������y��o0�g�+Q��6@�ۏ׺��6X�M����%w�^mKwm�8d�Y��y��P��@�g�쑼�iŲw��g��^�:��\��tp7�dw�O�Yα�ݝ�+2��d���K��>KF�y�|�I�j��[	^���]o��z�����-���tǄ޿��0�\Ճ�{y]�Ή�%��G�C8�q��7F&���+�Gf�q�9�<:��25�kmI����äR����oEIwf����xffQ�xia����I�E�ϵ��,�VNꥧol-�dn�*\�T%T�]��f=w�������=w׫t���	��"&���������S�3���mM���N�A��ɺ�.3q�N`�`��o��;��g���ɏT���l6��[�5{��{Xz��'a�y�5H��z�"!��q���|�jt����u�rLa�.6X�1��NYܸM����ؼ�|;4��T5	Y���{����� �z��o����b
xۆ2�H��*�o��=,�?�;I��U��jY���{�߅C�9n�s�V_��n���#//���F�շ�w��?��Ä G����=W��}�o4��F)�l���}�����g�5�`��c��8q�3��b{�����l��,�l�\\�O-�ׇ�x�↲w���<�`�R���U %y�C-EZY�o���`i�~��e�53��vUޛ�*���Q'����}�rZ}����>��4���Y��8�S��E�n��*�[=�u}"��O��ɨ31�ۍ�7$Ƿ��Uq]��c������^jlw��ݚ�A`��y�/}�*a����Rq��c�q��J�6<�����EDM�:���/�S�ז�Zx���*9�wpf�e�vK��@J>��Eet�S��ݏ«���r§�6���T�VF�F���Kx-�ٸ�鑆�)�]�M8�͵xxA����n�8,���'�9z��y�-	,�POy�]�����ry���{n�lo"�q/%�}�W�%��wW�g+e��/:�	� ��yl�,t�e��-#�da�M	y�p��%��j����R;W!�i�~���%��R�r̮['P�9(�7�<t�n=#���e�򾯏B@V�6j�qtYWk����������(2e4J�P�h�b6Td��!�R��F�4h��r��S{ﯜ��o�`��ͳ��� �T�_~��石חY���~�����{j���`�eK�o^m+�i�e�Ђ90�ӱ����m���G����*�ۍIf�s�=�>g��[��|Y��Z�$v(�7c�����6
�[]z�se9�]�1��73��9�\>,�9�<dDVu]���f��V�J�a%j9)O�֟��|��o=�ō��S���F�g�K�P���8�;�je���Ni�ѾKvB�&i�i���9��٫7RS4;��N�v�GDL���vU ����ԮzZ���f�����Xe��O=}zA����4�O�:,6M�w�{�J����;f��a��bɽ�w��$��a>
�,!_���u3�8��)]r��ɮ��1
N��L>�Y�[=T;�<U
���n�	����g�څ~�X1��g����d̀���b�,%Ƥ�����p,�0:�޾��vP�X�����r�O2�_ݴ^�Lc&���i|χ��x�b�W��O?]�����|]�9�b�gfr����L��[w;�9���5tV�zvw+߼|||||}�&�p�Zt���h)	��m�f�g!���`9\C����o
�ryFnj�S	g��ڐ��>粕{b��X>0/@a긕�h�/�*6��﫺'�*�Cu4��n�6�O�'nRwR�m9��x���'a���v5TR�3V��p��Q�$媒.)�ZZ\�ֹ�[���GW�^���vvg�`�*�jő� �HE��q;��	�0sw[a֭���f@;w o[Ǧ��	�G�P#�
����_M�K����J?v`�+o�̈́�%yq��f'E�j����W���rF=?O�0*{���՗Ԗ�bQUx`�����#>l+F�!���ffc�f?{N<޹���,��륕�7�:4��C����9몏W$�w�7I�>��2�&w�;
V���r��=[7-�x��;��1���g�/gn|{�û}��ަ�ن%wGmeq��X_��G��t��ӟ��ƾ	팪�v񇗗��5;��W-7�=]�^qkWj��W��ܑ�nw^���Yj�(ë�K��p��[�u�����1��<�y�hre����Y2�@ѣF��7s{��dl�����>^�Ž���0�a����u@zC��D��Ν[5��f6Z�
��wr�ـ)O6-{���*˕���>�7�
9�ƯQ���o��{|�!{��:ڗk�Z=:��w��o��b�|��e�3O�߂F*�cg���N�hp�q�-��{�jx̬�(��h�S~�Bx�ط���9��H�46X��`<s����.�#;NX�B��7s�-*�T�筀G=[�G��/�P��M�ADTB8�]xMż=�ha2�Z�=%";�uWv�X�P7�y4��FNd�T�*�O�hLΡ�o��"�!�OUT�ؔ����Ny�bƙ����9����/m�iF���q3�)�r��S�Xo f��<�X���4�7[&����܃4�4��E��N�NZ��"]:u<��x�N�أ}xB[��Flq�]y�fⅻ�*�<<��'g���dѷ�u�!Bq����}�OgMN���;j�l*�o�@��Oe��4<�!�@/�A#:��������ʤ&>�רѣDDS�|���~½�]�� ��. 0�?�e�Wݲ-�|�:F�tw>���3TҾPs�b
�O�t�
���h�c�k����n�kj�j��e��O���/|A% ���R%�+�2��!�: tN�t;��������-ٛ7�׽WRނ�/g�1�K���F^MS�;:~�X=\�R�r���.omv�6/$ݳ�Kw{����mv����u�u����R5��U��̪սO��Ǫ�]��	g�g[�h�o;�����6��V���Tz��p��gѨW	�za�f�v�<�(u�f����WW�TзN%0U�}}����R3t<I�� ȯ6��WO^v�V�q�����fZ�ݙ���0c���Gb��7 ��N�1*��>a74
>�D�]�9Ƌ�=wQ|��Դ�ώϜ���9΁�v���3�;�l�슆�{+��;�0B�3,<�۞V�]ȥ���59qm�"{G���5S[|EꗾF�?�Μ����OS���
&�(�T�����ye���K=�k�;�#/8VV_S��-oW]o\�o���N���\1f��P�9���q��)��)$Uh"��!d�̈́Fez���oՌb1v�������涓�H�,�{�d7��
�/7��;����&�Չ�.zN��h�|$���R4�C)#a�+)H���J�0�8Uj/��qy��d�*Ӹm)��\�ʬ�l��y�7�Pe��)���Laȴw{t����{�xv{exֺ�ĸ7Ane/MD,��k\�����aU�2|��)��l:$wcȼ|#`nBU�#�����8%�fMNR��j܈ɖ��P9`_��Nh���#����-�Dd��͋YV�7g7����ۢ��6H{���|�3N�<��j�k�a�my�u�-ŮH�wLg�w�%�c,����8b���<��2�<���׶X9޾_V�Ŵ �O�����H��-X_p���k�߽�0m�ɨ��u���6��oZ�"������}�2ɾ负۪��>���!��\�C�,C��w���Uר?U���y뽁���t��Yx�L�<�M$3X�F�_\��q|�HiA>B`�GǏ���(uv�s7���V>;݀͊��!�ی̄���˹K��
 ]:�+=g>m��Fn�3�G�����F�4j���i�>����]z_�s�vTG@{'w�BD��߃�����Õ��D��w���%��`��
�
�~��Pm��q�|��15�����o;��N�o�/ꃖ��(�ў�=��k���=�q��CU�M6n���{��3ٛ���n�����x7Q�]���lؓ#w7�z�2�ͨг:A!C�wD � ��4.!���<��;���j�z���i��h��y/1qB	�W�Nd|a��M��E8"�on��N.ݫZd<D�D��l����ˏ{�bBJވ��U�Fٽ��p�:����o���c�2�h�vww�c�v_ү��c`��>6��K�<3�2�n%kM��{����qOZ(�P(Adz�=V��n�T[]4�8�_�2�5�bc�]��'���4����T���k����3K��s#LWKV�$�m��Y��U�t[��r�Y\&���o��0�ۨ4����+�f[U`�J�֚>1�y�9s��#ո��Is7�K��HS9��>���������K��w�^���.<�,�B�'�O��Z ����'�O�럎��������?_�q��S���RNeG�Ak�ǅxoNW8dP�Kyjaf�n�e��*.'�>�R��'�&_IR�<18O=��MS�C��q���:f`��i4E��l�����zH���G�r��z�/�7L.�~jh����\����\�^+歱:	�j5�\��k{y#�iM�{�p҅����n�U��V�u鞝݉��{M[�F:�y�_l��s�Թn��Z�}�k��P�8�t~|�X�V{8'9e�W���wOZ��N=�a�����V�ܭ�է��^{( ���\u�m���r�!����y�5�t,�� �8�5��Y.h����ׁ��u�h�:P�˜2Y�K/'j�Ez*7i*n���J��.dAx��:
a����4�w.E����G	����;z �*N��@�jMKVc��Р�Q������"�d�u�۹�z	��N�����VmGY�ϲ��W8�¬�꿄[�2r Yuq>P�.#��P�hW FV,v`͔iY��t�Q�����`�uNG������ޣ�ؠ���}�΅�����B�4����]�Qt
�	5�u׳CɻD̀����^�e�[���5f�)�2�Hm1K��wf��Ƌ��}s�Z���}�C��3\�8���1�PO#��y���M2�F��3�	������t}N��Psa�m�ӀP��>�f,�����}-��|]%�ެ�l�P��5�؏m�3d?d�� j(Cˉ#�oT2f�Gg�����Nŷ��G��w�rU����Z��w:�����D����~���U��$���q:i�>��jF�K�����vmA��㩀�9e�z��}��g�.QD��g����s\2�i'ݚ���s�܊Ogq�(Ŗ�)�9����N�ȧ=\	�j�N3���/�N ��w�A�l����Sw}�����+[�}�AC'�S,4q������:�x&����[/f�����E�`��
PL]���C�����%T�o_r�*W�I�ߓ�<g���8�����y#�e}�.����*��ݳ��_<ÆU�+�[�s�\�P���g���䳥�8��w�g�רa�����w��b%c�o�y��s[k�exD��t5���������l%\��vb��h�o>Ղ���NN<n�z5䖰n6�=τ���=���!���Uyo��oT�8�.u�U�Zʽ��nY���X�j<�w���A�M�5���үK��2���7�n��e�+1�U97D1<���y���Ƕ�#�A2����m^���x�gD<�v>�bwl��dr��wgw]s�Fq�0�ݍ7]~����Е���F�ɣO���e&�Q�Qg�{{{|v־5�ֵ�k�nݻv����=����~�/��%$�l�Y"Yx�<x��V��k]�v�۶����%�-1���Ջ�r�U幱��|�8Ǐ<x��kZֵ۷nݻk_����PT5E~+�--N���9N;t㷏<k[ֵ�v�۷n�׏�Y'�-��:�Qk�nh������m��p��W.~6�k^m��\-"���tۛsMf���U��ѱcZ4F�+�1ͯR�ך+����gu�J���Y����ל�6���^m{����sz�o5��ז-��Ou�9$m����׮�Л��ޜ2����3m�i����������[��+s��;��|�eLh��ۦܽ�/}��y��o0<V���g�\~ۖ��EwH��}��~�ipv��>w���"o�����S����r�`_����b�A�y#ڍ�v�2�Ԡ����i<YA�&kw��������aT���=�E�Ǉ%z��g��"��ݹY=�tՍ��iA� #5�׳�{���X��&0t���a-1���VSM��,��{��t�>-���}� 2"�+�V��>K-�]!�se�e�̒��ٻ[<e�}�M~������t
S�R;Vۗ4(�'*$�WrUȚ��`����H�0#�z�� B!��t^d�m�u��P�u�z�+R��
06��?;4�vw>����fŸ�P7 �����Xh�<^g'���XK��zB227����GD��W���J�:�,���do!H��ΝQ�u��JA� �˳ǻ�݄�����Xp!�c��~[���Hb(k}�s��~@2~�>>5��m���a�o���{�����@��û2��)��{��}L�{4�0�]�'>�Z����7����y��2�:ն�du�=�B�H�|r}�ː}��C�ݮ�g}���C{!t�GB&��V�-밆��$^Z�PO�v5)j�
��^����:��M�g�G+֙��e�9�c��f/�"��b��I�c�yQ.�S8 �\z�L;�]9�������-#�#/�+�S��Г&vv�̥6�6���&��<
`7�Ƀ���9�v��z��ur@t��*����nM��lְ3VNgi���B��0`��0^sD	���A�F}/�ܓyګ������k	Tr�`c+���K�t�p1��z�_H�i��t��{Ke����������Y��إ�禔� �]m�QԼX�[�+�o
B�Z��M��H���t��3����e�����.甘T}=�Rj�3pN�V���=۲醜��c�4�&3r�d�fW��D���|\8���a<�%N��X2l�ؐ��y�/e^���c��Y�U:�dpm�-����8)&�N^v,��J��A�W��t�z��}9ʣ��f;�8,�1�Cw2��ya1ۧھ���u����]�\^��wh��l��cf�b�)�RD	����L��	ā�B-!pW�� 4h�)��c��ߟg52�D4��gqe�Ȯ�Pr7u$Ozۥd^�ny������ʜ�]�x�l8�85��H��Í�o_)�KaoT335�v��;��˷+[�����B��7�4���9���\�7g�����p���ԫ��U�զ�5�P3u��8�����l[�l)�:wl����8dV�
��{��/2����A��>��}�-��E��*Ή�.�W!�a���6�vy���>@17��}����A5`�}�#V3=��K�8��a���Q��D屬P�bt��͒N�e囖7�ɦrE���k�7H^�<��.��r��^�IE�Q̜�������~�a��w���8��-�a.4�hj �w�=���h�m��ّWdh������N�p��Ӌ{4��\yW;Lbi�r�X �37W�|F�x�m���-����#)�7.i�P�o8fW"d��o���	�;e$�ׄ����I=���Ky���O��b���YK�i��SƩb����ĳ}���͙S��AYz�4�����Mjo/{��N�k���>ThF�4hz&�[&Ue�p]F}��h9���`z���C�m���]�bd�q����M�7tC7��u��z{���s/��Aq��3�װ�V��~�.��]��:I���c�v��
�y��{��3��ky�u5�׹�',Wx��=�w:#o��B��^�iNT_B������Ƀ%���#�Ҹ��a9���gw�BD��޷�S�{�L�:���33*���6<�-�t�FZ�n�j�"n��ok>l3	�7nQ4vk�������g���� `>q�t��U�֮��zU�ke�8-�e���7��k�������=�P�Ni���kk5��%n��S����$(H7�l(-{=��
����MOxa�SGJ�t)��p2�����nr�r���C�>�;�vzgP��}����
�{�&ž�f�j�1�|I����
������/�w��+	�g���Q3u��}�g��CHd���Q��!Ǻ�ӧ{�s��]X�﫲��y�+�c:nc罈c�};�=����:��|ﬨ�;���by���-������|�{�}��o���|��;���ya���|�p=��l
��h�;���[�4f(���s�zf�Ч�=�=��z��K�z���s34s���Mem=wDtj���g�cs ���\TK���\X��{���,1�����%S�*��wՒI�AK�v�F�>��>�pZ ������2���eEԏ$���5��K�$���-Qi"4}���>�`��{�yt����u���4�;@9 �4eT��4LTæN��=g7���8��5�����bOl"JBԵ�ǻo��,U\�O��!$��=�0h�O�<|f���=�.���a���3��EV��Z��m���k��qs��?oc��+�"z�p�s\#]�Mn�#�wwedu���mf�j���.�iɅ��!�[��fjv���C���>)�,Lڜ��������*�,���r�{����J7oa�<5e�Y+B�bz�--��k��c��dK&"y_s�k,��g��Ѕ���k�&U\�geXՑ����G��dh�b��Y��u֭�7)T�M����#��k'ZNn��c5hy��r�b60�o}������o0������:`\��&7��iU⍛�T��v�v�4y����(�fl�ޓh�����{�@�ҿG�.3ݐ�����#�F_%Y�Ө�U="g �h�?�!��{��J;��y �KRs���l��l�f����H��<^���P�Lta�^�N�R��gU\gh��C���*���X�����3���p2��־X&�g=ܰ�U�l6�`�o���?<�՟Lj���Iu�Ms��TxxP�(';�
�.���_����l�oS#Y�� J�$�c�/��>!"/�2=����y�
�UD���$�[B7�"��"��vil�J��Ϯ}RX\��2}�IE�3���G'�}�HFS8l�`�TK���(J�ϕ�s�ԕ:5*�;:桃�9�#�Y1j+tD׽1��{����Fz#�3�u���ʁm�u���9��^�SF��W�eX�����UKu�a73��߯+'�*�ː�?8����C�I���yy�P�2�"b�*\X-Ë��V�H�7[�T�;k���[��l��-���Zf+c,�}n��B���mk�ѣ.Y�p��"�A��6�k�hѣF���Fi6���gy��Ι�fYük����e�h5β0".�$ǲ��cS-eR[�aV��/2�+V�Gxc�����{��[C���R�C{kR4�0'�Tx�muw>�M�н:h2���v.P�]��z�7��-  ��xi�&��,މ���PX@��%��<���̿�-���S450�f��B�����\t�l&�|h�7,V����MFY��������8�q�(�Z���H��'lt��^[�v9gmN��끽��pGG�K0F|�:�t皳���vM�B��:z�'t��煥�X1��x�g����=��b�nkv�:#;���&Ce�'d�E8&=�/���pt(�ߗ��2�_z-c��)"���7�n�;K��M0�T6-�a�P���w%��_����F,e�:βEt�/��}0eOi�ؽ����'Z�9�.�g��m�}���vmN�)>�5f�/�_��(��u>8�C�Sf��Z�e�1\�c]❴�}�;�=ؤK�7�^��[2�A�fa��St������sU�M"F&���R�;lD�'j<�pw�L]�!��8�蜵�I�mS��������T�9�ln��X��J����n�;������+/VY��0��s���WC�_dU�7^�������PD�p��si�6�֊g91�Rۚ���J�/9\8�U��7�%E���ފ.���ǵ�mV�'�B�JL���������>.H~P�3ػ�M���xy�5��'@+�\l��QT�{��l�&}�w{<� 1�M�� |��6���[K
l!��;vh������^�es�9�@��3�p��o8�y��a���V� ��(�]�N���A�Æ�»蒷e_f�P�j�/n�{�wMS�w�gW���a�8�W"#:}:<�L��JD��̞7�\��*Kf�|�����F�vvg^�+�-O���DWB3(°����͗c`��we	�=8ޛ�M�q1֮�9�\^��E�խ9��#NO���zˏP������̏��咼=s'�e�^�.!w(�oقwo�kth�u\s�ݒ���>9j�%�����`����'su	+�	�+�R� �ddf���8�;�q�s��Hp���}ߍ8/��3ﹲpm��	��b`6[�w4}le��6Z^3�%M�gV��9�R�υ�z������\$���d�۴��M]���gyդr���z<�/۲�IW��1�{�Ӽ�{Pq�)������>5D�4H�mo{�}�z:1�e$`����*Vf{�ކ�\Y���O��2�|�oFt�-��xE�%��ݣ�AMQ���l�5��!�z�ȁW=�E�.�*�ŕ�f'�S��k^�:M�#l=��z�^+C*��#�ܮ��uwעT�˯�S��S��;w:�}��,�:���Q��Q�﹒vw��?qA����l�����Tn�k�3zc�|]�i��Ȁ''1^N��^�O�R�<dv�bn�m�}�6݁#��{x�ρ��K��g���>]�î�K[���ڶ|ӭU����&�+VR���P�	|�o�Dk>��_�>e�z$M�ٻ�f�7MU*-��v��,�XqNdܒB[ ���(�"p&�=l=�%m���*IAq��A!	��x7%ܹ��u�M5��;���d��,��k�T�fǼw/�i��]6�{+d����y��o{��l��)b�)������B{b��;P�7U�j;��Nɨr�d�6�Vz�F�u�8��=�^�=��7mM�+��g���j��u�� �f��R"�x��W���"��C;8��>Olw1�v���P1I���YD�̪(�W�I�W�,�f�Y��1�>mP��Ğ�;7�ZJ#	VE0����^�vx��NM7�n�s���a��n�sw�s��[���d �}3�E%�%��f=�GjԴBʕZSì����t捐���e�kj9t��͐*Vzvk,%��e҃�3��F�;��[���~c(h����k���NOwXڲ��񫦲Ū:k+��*�9���ۃU�{������k�A�ij��n�UM 	ay�.h<�{����a9�w�j�e	��\�o"D5�AZ����������~h�I��$�I#����r���"$��_�'S���K'u���wī��kMKL��SZf�LY�2֘�ֳ�mlɋ6�jL�l�f����U6�33U���S5Y�&j���)�6�,��U2Y�U��2Y����Z��YV�ŕ�����1����2ե�*���3[L�L�S�j��Lem1dͶ��Zf�c*Ҭ��f�1�*�Ō���T�֖,�S%��Ҳ���ZVZ����f�����e�+*ҳm�fڕ�Ԭ�Jʴ�VU�f֕�֮��J�ZVkR�V��iY�Jͭ*�ZVV�em+5�Y��f�J�jVmiY��f�*�ZVm�Y��f�+6���Jʴ�֥f�+*Ҭ�R�m�f�+6����f֕�jVVҳm�e�*ʴ�եe���iY��fڕ���֒ȲD�*D���d�1"YIk5�Y[J�jVU�f�+-�YkJͪU�iY�Jͭ+-�Y�J�jVZ�fڕ��YV��wVV�eZVm�YZ��Ԭ�J�jVjҳZ��ԫ5�Y�J�Ԭ��eZVU�eZVjҲ�++R�եem+*Ҳ�+-iY��+ueZVU�eZVjҬ֥e�+-�YmJ�Ԭ֥e�+5�Yj���Y��eYY[+5�����Y�+6�Y�+5��VVmeYk+5���������[+*���Yk+6������ȱI�I	$�E��K!kU++j�e��VZ�J)IdY	$�(�IdX$����$�ȰI%�d$�Ȩ�J�V�Y����کYBI,�D�Y�$뤎�$��-j�e��Vm��f�T�ִ��Jʴ�f�++k��[�jV[R��+5�Y�J�ZVkR�Z��Ԭ�]ڷ[R��+-��2֕�Ԭ֥fژ��SRejVV׽���5&[R�ژ�����Ҳ֙55i�ͭ5V���mwU�U����K-i�jZ��iY������3m��5Y�Y���w���__�u�/��ZD
��$��'��{�gg���?X�����ՙ�����������i���?��?������$�@��I������D$;��$�@��?������,��w?�
��O��Rq$�@�����y�O�w8���O_�=����O����N��'��ޥ���"""�K"��Y	R*$��K	V�ҭ*ʴ�����ZjZҭ6��J�՚��%D�IP��R%DY��6�U��Kjl֥Z�D���)(��K$K!D��Mi�KYmI���jқZmSZ��V�զԵ����kQV�ʴ�ZZj������J�U�ե�$O�(�I#�D����Z5��E�%�%j6��ԚԚԕiJ���2�)V��ԫMJ��jYV��ZSZ�J�l֒ĢJK$J*D�O�%���?����k�ʫmU��V�U���R�I���u�����?	-����2d��~����D�HI��'��;��'��g��|���K?t�?�e���2~�܉$�>I���R~�9�Sݒ$��I$�?�O�X�?�'���D�Hg�'��%H�H$�I�����O����Q�_�$�Id�l�}v�?dd꾙�d�$I$���I�'��?.�D�H�O�j~S�I>s���?��ϛ'�'�I>����'�$�~RȒIg��O����I$��d��I���>$�%�����NO�$�I�?��?�����#>I>���*{�{�$�i��,{{��t�T�$�}�9'�~����~}D$?œ�>��$BC����7����N�~����d�Mgqs� yf�A@��̟\����}�SY���UK3"�3����kZ�9:͚�ՠ�͵I��4��2Fkfm��V���R��ۻ��V�m���ի-m����L�0ib�lfm�b��1*�������<�gk7M��W��ݗc�mʹ�V����ۙt�j�3�\�]��۹�k��n�]��w56��u�up��wu���m.��v�4\Gu�]׼�;ݻgwmu�i�`Ϋs�[;���T�77uL���Z�۝ֺ��˻Wu5+;m���κ�n�ssn�-�u��۶�w[ek��[ZskZlRUK���g
�r����Wwwv
Q�o� 禾�2�H�>����6�{u�ԗw�պ�ڝO�o]նR�s�woi*�ӭ���n��VӬ�9�.��jW��\��׽�V�y������v��������Kյ�۱����ܣ�n�wT�9Q�]�   ���Pё�F�m5vм��g��!B�C�h�O��^�m��'��w}Ƿ��t�׷�f�����zT�ܽm�٢�ˏ[[�����ݶ�U�-����ۇ��ݦ�����ʶ�ՏNn4綻j�9�����7s��۝�֦��5]���  y���w`��<����dS=4;��'7��۽�y�g�ԗWw�v����oWh���Cn�^���Q��a뺩齀����@�G�=ޝWZ�8�j�;v���rMqΕ��خ�  =�j�P�_y=�=wZ�Uwm�����V޽oh�E��=��;�w�P���]{.r{^�\��cM{i��וv����օw���ڻ;j�7���.-�s��M�   ��Σ�<w����Yz�{j��u�{A�{j��{��-�kݮ^��=-�mUR��^���j��{��x�����oz�^�v�ݗWI�v廛X�Cu�㏀  w|4�Я��]ޭOl�ޯ^k��v��m��u���Ӗ��z���B��Ӏ PU` �z\� uۚ�  ;�z�]Mӻ����v;n��kM{��|  ��>� sp  ��x=  {=��  W�� zh<�m�� ۽��Ч�޻^� M�e�  w�m� 4���8vM��w.��n�Jmn��   �| @���  ��o �^  =s@ Ӽ�4( ���  �޸ S{��  ���  ��t�u��ζ��ˮ�kk��n�n�  ��� >V�  x����<׽�  ��^�  �z׀  �  =�p�@ 7������^�  ����6�������j`�Wwm�չ�  =���  ���� ���@ ,�p נ=���  $�@�uǠ�� :����  ��"m����Oi�$�*   "��	J� @S�����   jl���	� 4 $�JDU  ���W�G����R�����ώ����}����\�l�N��B���;zS�?�����������J�����[j�m��mkm��Z����*�ֶʶ�V���/��� 4G��&�6,�k��1ӹ��eV��N�T;Q*����¥���ތ�KiçC�z؊Q�6�d5�l��1��p]J3e��h����y[�M	���8��5rS�`K�m�&1c�yp�n��xRtLFM�'�)c�c2�항bͦ�4(��Z �M��6f ��H7���sA��r+آ8���]�i9R�ཌྷ�b��]�,H�La ʽ]:E�n��Ɖ	�bX�5�RT�V��
q�(�hA��K��ޤ�: ywd����:a�4|uy@^0��֟���@n棭���̴ "%�ՀFn^�o�0+�B2�MV���6�:�'NMB���J�r[v�%n�k���ذJ���v�z��~���jc�b��D�j���v�:���Rg{YǊ��3b�e�sN�e�&VIb�mVMv�S$ߍ��j˔��*-Vl�Q���H�m$�G1Б�n-S �ڪv�V��S6����W�4���1Q�2��j�m;hm���]��!J\ũ����ϱK)S�E�,=�׀�z�Ӆ٢���X�:,ـ�sN�h�j��YyzL�0V�ld쩥 1ӿ����R�o~����Z��{ ����
aU��*Emѓp$�I��;���+V%��1Ec�Q�r�Tܓ[c�X�v#٦��lM��W��wJ*��+ ���u�46��P�)���U�,�4��(K�ש�݃m��?��&ո�+eڈ��f3����QRT�ס���i�>RɃԷD�[���*�-91Zِ`٫�hL��IM�6M�:(��&-����Y��r��̫J��^c�&�Glް�"�Q5W[��-�Jn��w��]����d�omb��,��/R�\�0���AUӢзS(�Kr�EX=Ͷ����.��f���Үav�
����\�7�,VH(�/,� 䴕+Il��QVX��i��&A�]�JMt��]J���ge<e��@
2�7��޷�ۗTU�����DU�B���/(�n���S�1V���0�D�b��hڻنH��Y"��K/���V��a��Q�B�X�ss��}j5��ݤ-�VR�V���#4C�8���í��,'�Р�efEz�*�vk^��.����
*2@���s�7��Ÿ�L�+x������M��0n˗J�H㡺d���l\Ini�o~1�/Y��O"Ȯ����P;,�{]}���i�d�y�,7�݋�^H".���ѻ��8�x-[���T׊&��f�;6�v7t-W�-���r��I�h\�J�BR�oU]�I�	��v�e�M�yii��rn�qIl�
��vdՋ
{�O_��7yPZ���u�tJ�7:U��Q��[QT��=5�ݶ�h�����^�`[!����Ix*�i�oӲ��ú��D���K7�����eP��uu�]6���/����7C�v&��m�RH��Hi����AT����X�Y2���ZˆB�)���m�Dw��SW��#�p��aAEv�H1��dEGS5>.�:��傦��n潲[pn�q��u�;���4��ɦ䰆%�k��$�+]�t('^�2���'t�#ڕl�;��"<oƯ*Ƭf����J,[��P����%��1-��pȁ��:m]�#O�Fj���2SD�&��x���,Ɍ�VY�
�`4b�J�S"v$��!�n�]�\_U�4�f����"�*�*	dejG�^I���B���B�g���	�b���BPg��Q偃SO+&ˎ��E�����aCs+9��b�aDj�bU�F���h�,�ց����������E�\�;U�_H)D��}GR��Ylk ^�³V���j<	SY%փcIp��H�l�]YGV��ݬ�b�9p�+U%��76�+B�e2 'U ,��=Բ� �Y�PeT�[���V]�
QJ�^e"��I4�&!Vk(f|�y���;�t�RY9�"�b�aӗ�,+c�r\Qe���mԩ��.�b��j�Z��(J#.�͑1��(i���/I��Ê��nlMf��M[2K�h
05��TfK���	��;�-��$J��&��7qմڋ���,81����Qh� 2�w�v�h��2�� !O�:���+)	�Ȕoi�A��(`��ToH��{J����h��P%���ߞd�\��m�Jo�Y���c��6����
��(�L�e��i
[m�晛aQ�+X�%�H��;yW�r`�U\���=b�X��)Z
���FY�JHkH��u�VY�PF��ݤFj�ԆO��[�x�˟�^'F�R�$}��"Tqm6>E����r�Eӭ�+~�Rl	B3V7J��ղ��aF�$Q�a�9O���n�B�ؘӔ*�c)2�+�fP�P*�c�e���gڷ��$�e`�ux�*=	PfSxv�\�!ŕ(	VtᕬZWQ�b�ǀ�6�|���r�b)[�+ksl�Y����8��o,#�Bv"Q�dF�SV��	���� ލe�f��ۧP��� �`ћcI��%��QXy>p��P@Zܦ�&n�m�uqMC�X0d�44�daԔF*�*����È�>A]���1�Vb4M�L4�mdzg��,k�diT�i�X��O�Qubf^!R^�j��hS�wu.%)wx��:�Url��B���Q7t�k��0�K3w*�=	2�j(��z�V�gop�;��ۖ�xT��k���4n����miU��x���Ů+�W[ª���:ۺ�nϰ�5��L�WX����X�̽�e�K6�4ک�yv��y�����4�;�7Rgv��H�67�K���� ��љ����&匤)��U�J�5l1F��'-]�j�ҫ���O�-Uv�0�go�V��X�-�U�擘X�ș���+��ǅR�K�*'3&�SU�;������J��	n�F��lk�ɧ���T "�ïD�m5,V��� nSl,�5}�,����+ki�h�]�pf0m�:�Z�9�HC�.��`H�lݻy3
&�bj��^�<
����R�٠�\G3TI�e��5 ���iǀ�jݖN�N�$�#n:i� M��f��?��)�7Y(�Ha�JK�.�n�,Փ1�� A�-����b��	�zY��m'�a�H���Խ۹�, ��Z�]�h`O)j�P���͟�'����a )�H �; $�6�*9���6cv���X��w/r�&S�w*5,%E�jPq r����eؽ�@��*ԣ D�bz��劙��H�cN�6)��	�O!y�Z̼��Q[Q��EdM�^q�ƴ�e�e�b<�h䬛���R
������fG[FFe�cʲ�#��P�v�u����T;f�iD��;���1�u�(�v��Ԧ\��\�/.D�0R���Y�(Y8�56�%��CY�JaWhL���d ���6+`�t1GX�A���;�u3dqȬ�Ed�QSY��N$��$g*B�����B*H-����˓I��I�`�x�흳�¥R��=:�]���jeY \�x��V��j��9[X5l#r�R)[�{Q��Mj�b�9Zti�@,SP4�HJˏu��+b�M����U���:#�E-:8�%U���`m�4���]�%�d���O([َ�ً��p�ff���DEj�W�U�;�z1���j��գ�C[ou}wX̤j����Kq,���j��C��*黺ŦIjӔ���V(6��\�B�*(���"�(����)(�Î�ݎբb�vKm�@1��Ẑ����2�|2��Ōяi�5嘥ʻ�݇WYK5�s\�pa�Nɶ�k#w�1;�v�Y.�F�YQJג��6�nɔ��j�bT�R!��]����%�'nś�P�CCv2��gsf�M��ި��T@IЧ�w1�R�K�$B�A,iK�R�[3E�!��(������$�Z�@�r�����M �-��:�(:[U�3!Iո�m6�t���<��E�fֻ��Q
�e^*�i� �4m����.�me��e'��!1!{��T�Bauw �bָs)�"��v],J؎�E0��C��!:�t�f��A�L�B��T4a��YmM��fmQˢ��V%��u"��N��]@a���e+.�#.�O�nɷ�cMekY�R���rl��%L��i�H����[(4��{H���x�n��m��1�����w���-9�F�hd��ر�CI,V�U(�]�L�'�����f	CC����)�m)Xŧ�aQ�u��S��n�:r��L�YR�M�n��ts.���oI��j��Q�0�t�=x"� ���A$�� Y�R�)�ML76�U�)��D�f|��w��fD�:�2.���R,��0Xd{z*Q�J:^�ܻ����h�
�hj꒖=�&����`�ܼwnռ�ynu�ؐ��:�X� G�fiz�3)ԏj���j��G#
]2�R�V#̴�Z�Bm��D�H�xr�TI
U���@i�yb�kX-n�4嶵$�P^L� S�F�U��v�3CFM���
!%�.H�ۨ��=�[0:��մc�X�݃ #D�1`Z����[�M���v
�yw�c�eݚ���e��J�h�M2+�wD�w��qMg6�"�i��j�!LT�s=�M<p�GjZ��2�٫t�9M�X��M��Q�U����� ��(--Ø6���	�&B�������J���)-���Iށ��eo����H�
�e�Yx�¨�ؕm5\�.��[=bƢ�J�yV�sC�Qq�5�#ѡA����ϵPH��́א��&�@�����<+a��Ee���tC܃5x�Ԕ�,��E-{
�u76�%j�(�q(cE�w��WY�T�U��wu���6)+���(��z�`T�hu��E�
IQln���m"F�w�8NQ�٥��( ���r�1	3^��+4m2<,�-4��f!wb�uhP.	sA�x�&F#���d�V[�bӘ~+?�@hE�<!R�L� v�:��+a��5f�%��2Q�U��!&,-L�i��T��r�v(�EV,Т��G��F�ܴ�`��L�3̷J�t1U���,����ځ�5�@jݚ�mA3e��V�>��hV[�ƽj.<�ڤ���#����	Z�BF�Ĳ���fՋ�K*���m�D��ͤ�x�($*M�v���' 
�^��G
n�4��2��Tn��.�j�Ȱ�t�sSb�PWt��n�G4�WQ��Y�I|
{�hr2�l���`ʐS�K:2=�i������iV�mD��t@����q��N���԰��s�ؠY������Ȳ���̧�2&Ɏ�ʚyQVR��t⫭�.\f�tPf�6ݪ���ՠHJ��7%��Y��m�P�x����aQ��Ly`QDm��н��H��b��M�
�f2�4�/Tv�)�'�*���X�-�Ad�U/pDlh�Υ��hL�/
o@
�w�ZMY�F�b�nƯ��CX�A5^�h�v�8�$$�e �����A�oɪ�ի�&:�,�h�ܼ
�ʽ�c ��0Twgre��x�3�������hm]m�\يݓ��(a�K��J�]��.\DBA�.�R�\aJeL7tZ���1+sv*�.KB�n2��ݚ	�:�(�H����;�Mp��^}����l�������М�hڪʽ�e@���A�74���q�A�A�g)`=��݂�(�VQ�3��i$*1Q�-���v�vi�A��҃���DLk3�ޤ)� uc�rk��Z�JR�I�oi�Jh�l���#���{�<[+*a!�j*Lf`ڹz :p��#U�b�e�u�k��kwF7F���s+!yjӏ�#�
ú��)�;A����T`�&c�0��Mm���̔�ͩA��lU)��^Ǹ���F�K2�.�|��m�%V�P*������s5;���w��m;GH�x���& �֙���-l������8�n8��Ь��hA@�R�Շ����(`ڸ)�DV(���ڷ�w`7 ֖�)5{tv'Y{X�i�ڏ+S]+��=:�خ���#6Ԇ��L,��$X�,X�F�8��̀�3��\�m$�1[�>��v0F�hRk�W�ܠp;f�mM��`&�.����̕4��Bs-ԧ�@b�m������2�3��%U����Wv)",���Vtc�(��ż��[bZ�	��݃a��g!�&R7bV;$��A1���6�$�HQҕ�&)r�H�̙6-K�[�s~�+ݩt�&�VP(+iSdꌤ�� 
̑�w�m�ɡP��z�U�jW{�̘�kb�_ݻX)
�P M��	N,t�C�2�X��vU!BSYIjE��c.��XP�r�JM7f���*}���⊯s^2�	f rn�a�W-V�t���Pd[D�5v��I5i6��.h#u>����mi�BJd�%�Cf�x�"��V2�Y�7j�^�Z6!O@*#��˓�,�mT�51�>�"�Z����J�X����]쒔`U�_�-q)�	IY�N?��&ݖ ;aܡ�MY6( ,��Ӱi��xN��c@R���ҵbe۸WRԺ7�G�����:�hl�j6oM%�C,	y��v%�d��.[�W�sp&�x����I��a�һ���e�-�)�+UZЛÑS�a&�*ɤӠ 1��/c��,3%$�]�5v���#k�����nat�2�t�b�X �u��KP���H��N€�R�m��¸*)T߱dKt��Q�y�'GP[k/(-{;�qb쒆����f>��.h�禐b�)��>���YvxD{U�b�\�G��=zEh�g�u|V�v���5)IK.�*����.��glD�S.SW	�������5�=�Ի#QL��ܰ��$=�e��Z���<�E�,˨���6N<]�D�w��ۙ�b��:G�<(+�U⠶�^E�r�����Q�:�����w&�s�U2�b�9�cR�0��Ѽ���],S�3l���2_F͒��,�D��"�jB��(��6�$�
�q�r�^����PeY݂^8c�7%<T3����9��LF��L|2�,�%������{o�o��{���w;�uu�dtB���z�r�t�W{�� =wj�q��lzx^����ڨ��̫����ue��b���l��Q�٨uv5͗j�eB�z=!�e��h˾�1^���-��c7�g%f�s�v.��:b�ħ�lK޺K�]�YB�X:7�tS�2��v�=�Jty�P�+�=���H��#���<O`�	�v�v�p����^ͮ�:f��n�U�gZ�-�	�;&�헛 ��q�����V����7նk"����ӬR�+��HH�N-�^���N�Q%�v.�wB��c��%*�v��.��qN�-��=�y�ye*o%>� �l)�L�z�t�i�7+���{���cn#\S��X��/�F���LݵR�ّ�a�1<8��Wl�fe��6�v���</��툾����Ү��0�kT��$^u�|�b�ga�\{�7;�PHh��v�s6GQL����n'PCz-��F��	�d9L�J콵��Z��T9� �ţ���ܴ�C	�����t��`���e��r_p_��Jg�}2�./��U�Y�&���<������� m: 1`���N=Jo$RYC�G2�mv����TG��Rǚ�C�E�TK}ݕ�J7�m��Z���U�M�jDRP���u��X����='���9��r���rJ�.�)ő��[�'�oq]L��Ը����	S��(pV�R䙔,������.R9�(z��}�,�f���U>L,��)�$�P����Et���!���s9�Q2����h&Y�՛[����$d�|Ewf �X��ƀ��e���+s�F*�WVN��j���.��2�\�]6��Ʈ����_,jC���Y���}MՌ
١�J��; ��c�q�6�r�W/n|�������W���v�s$���6���2^���ǐ �X�HENMΞ��^�Q��v77Ԇ��K��'��S��1(Ջϻ�l�gP�zۭp3���Q-�P�4����p��F��K�M �lbn�ν��	b��d7{|��6lJ���%��[խ:jp]|����ăV3�3�8Z��3.e�T5�~������%��n��J���:�8�m����E��ia+3L�tIYLc��澂�kb:�=3�Ͱ���X��ު�K��E�Ww�R,��0�vM6 .@��6��V������k3K}��.�7�m�ٍN6n�e�]=ݥ��Fv�ft�f����oc�v�;��Į��oΖ0O����iͭ�F>v����m����e�=d^�,�Cev�zP���W��`��ڄ
������yd��۠��n趠�-w5�Ee4;�'��AS������wKǗ�~�����f9���	`ޒ#F�T,���S;sΝR��'<Zjsb�XF\�Դ�̊�Bΰ��T��sC簪=�_4	|�c�NY����v���^���p)c�z�Gp͘C|sC�oM�p��z%��X��+"�'�A�:�S2^S���&e�P#]O����z]�he�l���9��ܔv���Q�k7��-�ж-��Me�i�2�/�E� �C��p�Xo�{*�I&A��܄���w%g�;4%R$Õ�е�6H��)�h��ˢhp�J���
{v4��cW�Y3�O�t����3qe�V.��g3cv��GzV$6��*��wUM�goY�-wC�6���lHԄ�m�ѕ�X�|m�RR��f�G���U˷����>�����E7g������uw��܋á)�,bHM缮�Y���[!��%�f�8U�!�������,u�q�ͣ�墹=��׷�泚z�HB���s^R\&07�e�ܪ���u�JM���/r���Ë��	̤+���Ψ���q(�nC���[�l��6��]|�\�\NL"B�� bN_v���%����UJ9WpD:;��!��겦�Pe�z�qń����(1v�iR"*+X�����
ӯ.�VWgU��\g�f��9���;6�z84�A��a�f��b���K1T�Jr&��Y5�h-8��tWȵm؜��+<d�*lׂ����S6-���N�<rq��w��<�m0�+�R��ܳp��J�'ܵ�f��R��o{��u� z��]l�*^�����O,J�����5.��wnL]׵��b�A(�Uq��۷ML��,���
�Y�n��V�saL.��7:`).���T�5����*��īl��x�S�W��n0)@���FgA���c�=�;}p�����%�'}�CW��J�ꊺ֠�h���\����T��460�������B�s�y�8�%��
j{���ñ]n���ꮫ�˼vz+�]��I��Ҡ�u���'D�.ݧn����H�A�s��K��{����e���cT̈IPF�A4�Y��]#�f�-[�E���]���+9�ǫ��w�=�!�$������Cl�z��x���t�F"î��9��N[�aξ���w�|dV�I�����6华+V��l��;u��V�����s�E�+Q��x��WV�]"zq�ќk\"���֪
C�>�m�S�����EIb��ň��E��f΅*�����1Kjx��g����Ui��#=��m�N��w$�,U�W^�E��spZ� �N�gEҭ��
ns������Ȯ�u˹goN��Zq�Qj�n�`c"��1�I��Ou���乵�{�����ڲ�,��@�:u�Q�x�wC0r��>�¹�f��;�Pe-՜1%��$����\�m2/E�V��O��0�+7#��1�ǰ�ۈѣ�z��>�T7,���[&�7��+�Y�G4�0���V�Ytժr�ճ���v:#�u~����(a�A�E��zC�IV���A#��UoҌ}���v`7[G�M���g��TM2�ͥ��`�%��e����N�N����}�7ܩ�$\)�\!�˧fKf�=�N�F�;`Iz�S�qeYy�X���fuI��O^���&�gt䌠]����z-8.h����l+/�3�M�v�Y�Ѽ�>Z.q�VD&�E��1�C���os�#[˵_f�0D5 �˨�g� h�q9�nrB�W��J�\�x�|	;��ͽb=m�����ʱN���XA.�E�a�ŖN��[����,%)�dޫXl f�鵽��]l��\R����̬�V�Eh�\�K�+��h�5&:�5��sz�jU�®��Y��C/��D�Ջ��PfLS^�j���; R�UY($�[��[��1I�}�*B��軡vM"�Q�/�t%:�HBmb���@RtȨ�i���ʝp�����I��ݮ����[Tv�v��b�.|�,��[���2;������*@�C,٢eK�
���(S�T)�i������lBgco�´f��8h3��<���5G&��H.e����אu�Wh�C16~��u͔& ���9k)�XD���h�Oc��tz,�`�ò%0C*Rz���v�Sxp!T��Nay�*�����=*=�%�����T�I���PbM���A��xi۸z0���P�
��"�ءC(�ɥ�$������|�ice��z�U:��9t+��*���>�D>B7)��IӖPY�Vc�r7�2ӻ�����ث�WA\�Af�����a6�je��ۛ&��<�Yat5�x�ɕ��*��CF��եٜ�1�0����)��\kkYȬ��N5ݨ���{/c��@*�ɹ3M%�U3��t"�Xu��C�ͬ�D:�Z�����^�����Rѝ�n������t3KN�tq����`ywC�<�Q�0�^�=:R�+-S��7Y�xyqݲ�eP��"n^���-�X���ۧ��ۊ��$���\���zd��^�TS=�	�{m��ͦ[�6�H���.�%�~��܄o���p�}T*m�+8fr�V�sP�pkq�+���hRK�mؐH)+V���:$���`�2 �[ب�t�s��9�nV���7�0k7b�����ӆʩ�k晆^n�p@b��lc!�"ZKN����ѕ��;�H���m�Ԕ��7Wb�Gr���m!�;��$�!�x��]�g<n�i��L7�K��o��WSpb9�vdY�b�h6:�
qԍd��Q"a�uP��C��Q�0��ō�7DW𜴸]�(@���$56�a���^;��t�c�(�#{k	��u��n>�`fu��	J�ͮ	��U�ؙ�
P*��֨2v;��7�a��_MW�Y��Q���K��;�uy���29�����[��Z۬�l��Gu�>&w�vs�*[:��;)d9�y]ĺ���n��[t5����R�l��u�;�W:�ޚ����%e�I����(���9ŚV(\��x�D[����)L�0�/���/���
� �Ge���k�]�*[m좹�]w���̩��rU�h�����*��}����7&�eGq��xJ��^R>8���)�%���"���W�9�X);�z`�]E�v�m<�z��f�y2F�G��K��Ƭ_6u�}^a��`��H �*�#e��V�7�����6��2;V�w��m%G��hr�;��=�5s�m�����˧K�FS��%c���c��s�;E�.�p�ׁ���Ӹqz�Z�vpy�Om3����G`��.m�w^R�+M��)R;#�1��J��67�5d�(.>��wS^<�깻]۫hZ]���@����e�!`ǀv���T�ml���;���-)����Զ]N����Ι�R�uY!��Rǵ�k�fą�T"�u�\�[M�aG�����S�����E��rL(��<�v:�e�c�ene������{�TK��;s;��u�\�y�>�>9"��َ�BL��@��-:���ƱS��0!�Pv�N]����ς!h�˴����h6�TDL&T����X�k��L&��E�v۶����#{�p}��Ԣ�w��GW��;4r
�<8�C;��.�5jf@mƷp���A$3.�T��9i�X�!��wk촛����0V��{&�+F�\�׍]T���
�0����q������4�`�)]�Ⅽ�_w�^�&Z"��Ǹ�&D�K���%b�f��)k���d۵r�ק�bQ��P��bZ�g	l-lQ��@osݘ�Ә��	���Ԙ��k�������-*�Vn$�6�#��"��C7ä� ��k�>�zIN	p�;�|�'\X���Sȣ����r�����m]�kq��7�Wc��Ψ�6eӐ�Cn�P��BSv�\�L�W�l�/)�lWm�ӽM��iGbߝ[*
L�Ɣ�O 8nrDO�������T1����ޭm���8���XIo��.ʲ�T���̕�[Z8o��%lO�J����%�U��j��y�&^�F��6�u.���E�0pۜ���c.G��/trCM�!N�nCW�U�Eܲ8�a�Hk��@؛ZM@8_l�0�u��{.�kpiv��\�ٗ���{w+)�ٛ!��s�e[lV.q���`4���KE��j�YՊb�K}Ҽ�M�H�+�#/�A,ZG�ɶ�P���P2ҙV�������Ʈ���c.q"".gh"�����K1y��uow*C!���[�)�N�D�.ԙ����LwH;��+=P��+w���17lf��Uca�PU�)�C,�S�0Yѹ!��B)N���?���`}���T�s];�#�RfIk�h���s���!�lā���Be+q$s����cd�:8չ�A<� Nwm����'�ۭv�W �au�<���,��!�%tsKr�n�eY2�uÖ�-<3�aC,'A��nэ ���a,{̄�h�]tN�#Ntu�G2=��<����˹�M���ɷ�Pw��2��2cі|i���Iy�f�6�����c�}f�hPf�%�ᳲ6uur����"�t��b�O�\��,TZ��@jlԞ�;��9��3�f�MQ������K�����]�<dJ7E���p�Ylfh�F�6���k.�׉#�ym��n�s�]\��C���<�<3ֳvH���D.���E����#��')��X)M}\x�8��J�B��;b�˷�Vr���5!�G/��2H�.W-�f�v���[X��Zw�H�{)B��Gg65^6˄N��t��3�-_b'���]�;�sN;�ޥR=�J�ʈ�4��'X� ,|����L��'qQ<uN8C�PS�Ώ��vatu�Jas-��6�֪]�P�R�V���&�O���T�=���.�;����&�A�\ ު����
؏"�H�t�)�{s��guo_;� xfw�'Sɲ�Ix=���z�1m�c�'w�m�/�Ӓ����WBCLq�a�P
�kӹ��b(���gd�[R��yV8�7�"�����h�V�l��8v8*sW�jK讧��� ��:���RB�I�s6i�]��,d���\�*IϜ�I2I�rN�Y.G����� ����oy����H�����k�c�M@�����:�ݎm�V���y��:Wr��v,��Y����$�@n��лY���{VҀ'�
��WU��٢��=nլ��]�V���N6��f"(�T.�Q�*��5��ݮ�>0�����6p��"�qv����,S��lW=Փ��J�����ŝ���욛�V�ýSe^��Q�v�˱�5
ݝ7��N0Jy\�#m
fp�׍�{���Hsh��^����޳���At��J2��"�]��E��dh�L�	d��ݰ���R�P�F�w*�]�-ۓ���6r�������Q�%]5n�m�������M��t���'^�" �V�����YP�S"��& �Xy�7X�MSrs�����.�
`υ:��r'rnn�*�;�LHk�M�y�=��B:B�.�=[�oU֕�0_݄����V�"8)�a�� �&�9���P��Vhv��<��)T��GZ��(Z͂��p>�XuPyJ��(dU*�A]�B���ɔ(���h������8�C��;s%"7����H�,it'uR���~{x�u>�Oh����ܙ.��5T��Խ��AY8�� d�ohs��wY�KWgm���{�u�E�WO��K����Xl���K�)��6]Y�Н �1�
MԂy)fǴ��͙Jmڡ�T��1-�&D���s�J鵨��X�ړ�fo���>�r���Kn�HM�z�f�;�l���&p9�c�f:�*�GҹĠ�wbWgD���x��53��k�r�k��ԗ*n��\��ڻwfK��mA�էUI�����4<՛ZE �Q>��u�|6���2��1JM+��l3�1%0U�*p����J+���LO뼏/��sz�*� �0��Q
b���GDyәs(��(K����e/��s��F�Щ9wޮ���\ՠ�cpl�U��4o�+�4".u�E�⊫�ˢ'%Q]�Ҕ�́������*K�z��(��gEŅ�$�Y���̼�*0A�dɲj���S�+,mk�p-=e��f]�A�2p�e{�d�ۭ���Jc*��qU�95�Gnn]6�dX.�h�M�ɢ�{�}���(�:q�/:�����b�⍅�4T�bȓ�Ǜ{l��5�lw�WuÖ���U�j�l���n�Uh,���M/U�ՄYD�ʃ
+U>��K����p�N{I��'Y&_}�	�T��;�7���1F�-�ڏ�V��YA0w�
�(9�GBڽ��Ȧh`؉��Iּ4��_I�+e�qS.�1;�E�05�sbTY2� �\�H�������+��^�j«J6��D��Y��\_5�>�V����_V�}&	�������o�)��Y�Y���4�U�u9�j�M��e�2�G�`@��8o�F��e����Pt�wʄ�M��	�u��m��첦��+`��t��г��NS�V���\h+C��ٚRY�D�ޮ}Ƙ���X
0��}��A�p�PUٝ�R�k':鏟�X,5�(	0m֢و��;Ķ��s�v��!�E7�+�L�~x��&2�M]�A��@�t\|6-P�� ��66iP�����}v�^j/e�-RW���6ƶ�%΢��Q�����I��4�Cw4mӱ��N5Jc�#v�-��	8r�C�N�n���_�5ȕČ��b�߲�J��<��{E���vY��mU ���<bU�����+s�k�b��
4&	;�,�{;[�T���V]�m���jyje�Hos���bl�0�]�R�ػ�}��:9�O������vEX4G�:y�U)w 8ެ�s%δ\����DIz	�r;`D;r��&�Mz:9W|�X����ZvS��<쾣{ϩw,"�Q�a��a���1�O�헳��c`�c��k-��Z���fC�[� u5գ"����8М:�zA��Y�]Z�k	��i�p�usv��-F����ų|h�ۘlW	��d�q�O5�W����ݔ.�L����_�Ԅq�קu��A����w��T�C��5��ϙ씰*�N����_u��'iR0m�v�(#����ɶ*9ۉ����ھi�#pW]�,�&��ʛ!zݘcו�V�y_>�]Y/�@���#�*�K��(T�.gpۢ�g�%y��:��]\�2�f\|�v񱉽��;#+��)3�;67w/��=<U�3U]��b:�P2�g^U7�VSJMK�0=�R�Uj�n1Ȃ�W+�M���y5�ݴ�����ں�^I`��D����	��]���oM�\e <�����7���y�E!�*6���ir;��V����JWN|rn����t!#���Lb��p"2
��MZ���!Q�{.�vWGv2S�f�F�l* a�Ot���\�;T=�yةĭv�e,��tg-\�M���$����M��\��5bf�C:Ρ���,O�Ja�-�|�E� ���ԛvO0="R]5a")�r+����!�s�F��II!H"6�6���J�<�,F&������Z�ˡÈL���RT��.S�E����x�oMBe�qÖ^�̽��6�����䒔%ڠ�����\��%Y�V�%�nM�[dN�VIV4���x"��J7݁7A��@R45�������/hQ!I}zىv4Y�R�ɌU�"*M!�ɂi��ͬD�N�n�0��*�9t7����JU�6��f�mG݈�2^���5Xf՜�<ޖ�ט&�$�;#zS�t��\�L����^�&��{SN��8��l���VЋQXʴN�'�)Yk���t�k�gI�0��K� �,��b�����e'	�h�
�q�� 5��ӑF���޳�"mH�&��M��n�*
Nĸʟ U����W���m�9�P�T����l�WN��;B,nk�1ُ�g�Mx���BV��t��YZ���>��T�ʂV�4(���Fvv�m�x��7vi�kNɴ3�Yq���n�vM��5mQQ���x4�7H3+y�Db���]Ž��^�&k��/�"�mu��P���A1�)_`���Y��9��
�[Ҵҙ2����Ϟ.�j�q�;�<G	[a���mk����pK��;xs�w6ɗ�9��G:�5�v��2u'Z8Ð0�X{w[Z����nޭ=H�Q[s�G-K��]n�L��f�m���^��A�h�`^���h#,��`�z�����G�DU)�ʘ2���2�	��6V�����F����KGx����}8 {��deu��UӔ���y7iu辔����؅��T�ŗS_v�iN���"��Fd_VH���z��
`B���u{��᫏j%-c�m���Ϯ��|�ç�7��+
wC�c&mP&��4ڻ�*T�mc�2�gٖ�Cn�<�5���L�bMՄ1�;�<�8X����̡ڣ�J��#�e5�AZ�v������K"�f�jo1,�S����񜔥����v{;���7M�`1��rtfY��n�N�P�${Fq�L��6�2"J�l���M�D�Y߆�{Y*`�om�� Uf�����*p�����ySgF%�����.2��򲷘̊�̇9��<��j�g �6Qm�G$���A�J46���a	[{�J��a�v�t��ߝ;��%�*�dՌ��{3��(�K��ǧ�T(����6�(����t�k#l�R�FEs�C ��N��@��wN;�Kp���7�U}"�.E;�C��"�2:+��]��1d�Kz�@^E�{N�|��wCQ�����/.c��TT�����`3�����9�ڥO711��O::*K.	3��]^mgdWr�KhR���HfUڦ��"JȺ�F���r��8_k��B� fk�$��e��J'g��ײ����U���ķ��]���f��-��+�Q��Ό����u����0Ga�����K#��b����u�aw�Ȑ1Ǹ+*��7v
����k5k�GI�ҭY��-k]H�-�̼�]�h���;e���6To��N�Q�;Wuv8P�I�GV�,4��-��So z�¬oj��LF����Ħ�����]ZM�2c.�Zd�S�u��#4��ԙf$�7�[T�7�\��`N�
B����M�͚�H��f���LC�9H�uN�[svZ��BqdX��v�Oj�Ƿ�B��M����W�X��E&k�Vu�;��K{��\�n��m�E�$�7ܹ��Թ�]PY'5&h�p�U1�f���l$K�K�:�k�����V��WJ���/{�֣�S,�� 696��lm�o#�rmnp��C77�д+��sc��,��4������!���t��FxvJi�b���F�9B�*o#�v$�����*���m^KW	��Y-v�WO�q�B*�C����V�@�R��i5�;���0ۼ!��R��ptḽ���V�u>��$oa��Ph�fB1p��=�K�]Ѥ�$:��%-���oEMJ��Lǂ��i� �R����
Rw�y�宬�.��H���(�T�^V̕�{3�=cI��4o��d]'��9��V��+��.yA�)컐�1�;)���9B�K�h;�\!%�����M�L�Ss\o�*G� ����l�*�In������X��)$D�����;J�Vw�)�P���'�'r�#���ډސ_X�\�zϱ�v"V�ޓ��-�x�m)y�>)�c/E4.��Q�J���Cw �HPYW���#) �c�B�git����v1�Zt�{v`1v�����ӄ�/L%Q�'�]~ٸH�l���v�dWGx�Gc��Q��:V��ZL����3�k�����Yx7(k��K�Y0շv5_lF���� ����sz:�uW�����h�GjT�ÛVP�b�G�P��`��+��F;	��1a��Q=���|�J��D��˻޴�f :*���b첰�bȆ�������������׎��EHfֶ�-&�vU:�S��P�'�(�.Tx�ە�o,+��]"��ӽخYS�̜%j��̫��m,\��m�έ�;PV*u��U�r��,����Wmֆ�h�V3ks�l�-�8�i4�/^����\���ad����X]������A�):��>1�v�ҋ�u�������yt!��G�[\�0w��ǁ��V�Ӵ2s�5�X�;�hܼ��[�~�N-*՗��+�͙{u e���;���͘�k,�ۤ�NT�r]ܺy|�c�.=[��`;�>��k���c��jtm�v�A؛ݝ��HuI-۫�&v�!��8A��w��c�,X�n�+����H���gk'>��s��g��Z�2a���<~����ν�5��ʅ=������y+Q�_e���ˁ��%�a����Vq�MM����9\�uhd���Wmև����/LY�".��I������H�l�e���ڏ�;�s�0��v��v1.�$���O+�WL�N�Q��Urn�e 0�Π�&à�m\�$�vk���9@��2�B���D�]�u����Ŕj_N�ϴa���ť��xE���7|�c[�J�7l(c"�#���y�\��ʏ3��33jP�8��7ŵȔ������䖔���U��]u����c禲Ns���4�\YT.�X���2N����f�?�An�d�9E��/���C8XwzB�m�Z���/L�Ӊ�
�^�fe!���^�Ⱥ�����x�����uM�VZ��_&�$�W}o�}R��{���tB�u.=���7jtL�+u��h`���Z��3hk03y�\�i49+4���ӕ_+{�7}�ƱRo%v|E�����q8{�i��e&�"Tj�v'e[�C*u`��&�ATM��@��[u0%&�t.�v�yS�>�	U�)��ހ�uop9C�D��!��z�5��$�8��>%�vX��c�gE�kuf a��h!�%Q�mi˹��$�W�e��AX�A-�d��Φv3d���^��!w4t���˃ѣnV�񸚊�tr�u��]'u}�>{���y�sWe�o� ºt�;�ͪ�l�|)�e��.�p�9U��*4\�4&*vI�A��4(p�R�޽��t�@�.M�c�Ճ�KXJ��'^]'�@�d	H�ۍ����r�P�+��A�X;RϞ�5F�=I��48�:�I�e.8��ܹ(kÝ����Ί��N�U�I�,���r'~��*eT�!�䐍�X+�)�n!�q&e���&e�ӧ"{��m�+�'���9VaȞ_&�rk��6��rSWA6!5�ܭ9+�Ok�x��-P{ye��ͤ�N��ghc�,��
�H�0���Ȭ}�\���@ �a�_٦���t~�]%{��:�8%ɮKJ_^��-�a�
��3�t��2F��r�Ք��J��Q����*�tp��c�[��`�\ey{�b���2����l6r��d�z�R����,���뒴#3p��X��w��M<'Ck�V�::�t8�vI��d���-� S;����� i�j7��'cЍ�I�d����5%J.��X'r�e���AZ�n`��n�Q�
ȏ�P5`a�@Q�:J`ГE���b��+�Z7S�+��U�w�9b��Q�G�2pޱ���*m��s��R�m,@�;�[W�k�Y�I�B�:[m��|T�Bcj�"�a��w��k�����zP�p��ԹX];];����O31�E�4,�t�@���],��4H���9WF�{��hV���j)�\�.I+2�v��m,:�� ��n�[m��cx�d�k��ǜO+��,qx��.�*��e��&�m	7v���M��*��/�=r5Q�Ut��2�"o����o+��C�}!��nꫛ���Jڢ�5 xx{ޞ����28k�ks~��J�Ê&-�H
�/zQa�1X��S���u�尳���Y�']$���s �p5������j�J��s0u��ݵv���WN�={�:Wt�x���fΎ�Q �n�q�X�m]�b���V�` ܣ�غ������l���y`p�]X���9n���q���sKmb%h{h�'e��r��N�W$�:��q���0��"+�hU'J.\6�M���!���I�R�AW��=rU�y���WKC�W��"��{5�qYޮ����u�æ`�zT�깈�P?T���ͱ[t�H������2'��\�)�vzcn�3�!ej�A��ӣj��7
ґ0 S,�;Fp���j�Ѧ�#�s��%�`�&Rԓ]j��ʾ%�u1^me0�0���]�^W&��8�8@잜Ĺc�΃��r�-�NqȀW
U����\:dR:�Q�c_<���u~5��k[�GܮV�@˜�����݊� �m�t�d=�ԙW�`J֒�KJUǣ�]d�i"�`�:�E��V�M(T�:!�L�6V��N��swl� i�X�4q^�F,��F�փS9����nK���Y9;',�Xd�p�w6.��ћq�#��r�vJ��e������k%�̻Q+vq����ܖ4�6ѽl��0�o�˺�˩ #��v|�Ӄ@~r�UQAIM�.����o�˽����w]cns\��9u�[�M�!\75�ѹ\�x���;r�����F7;��d�ru��x�%�^���n�n�(���bK1�q
�sr؁˭r�f�i65]��s�u�&Ƣ�ם��yֺ��7(����u���q���\뻕NsI�%ЊLs�=y�4[��H9vXܽy]0�͏N[�,�w.���v��qH.�^.����]�����h�6����]ݨ�̘2�v��:R	[�ؠwzxɉ�"�%6Ld��t�H���n��? �����}�\W�b����'^Y���3q�s�B�SN)W:Gպx�v��\�bN�,f��%����wN����Dp�ڷ*?��ˑr���Z�op?��#�D�[2*۩�ә�Zco�\^�ݦ�l�p�Y��{�S����Jcx�4'*�=�|}]��Y����<,���V�i=~!�YOz���1pkbT������q��W���?
�C�z�U�����V;�׮^l�{X̥^Ew��F7|���MzZq�ʔ�m�%��jy{�T�(g|���*D���N�w$�9�Ǻ>��C�fn��u�)=�-��7�|�����,>�y��U��J�*ʤ�����@[N�Bx�.L'6
��!ֿN����߼��ŕS��u�n��R��ێ�����Y�1P��0�+���t��u��
U��Rs�+>\��]�lr�6���|�wh�x�`�{��n߫���ѫ�O�8\%��Hסt+�@��������k4v���
B�{�I�ѫ�]Hj�G�gk��.f�?.�����]4��G�q��E[�;�LF�"sHl�ifպ��������d�E �ϑ�1����{n��pe�Z?wQ��۱Z�v�&7Y��X�=E[9%ȉ8��T�T �E �A���O�����i7�Z-���9nR}%�������]����i�Z��*d��>f�� �����=��7�4<�y��t��N5P�;^j˴�|
�w&{��R�|Ff�i�0ɦ!���ON���	�C�4��z�)d쩛HB��<;�/��73����3�ӊ�(V <q{�[�CK5(�/Ld�z��5�ҝ�)b���1�Ӓu�5e�;����sH��5j7��Q��5��S-Po��G|c'PkA��	�S13:iA�=S�Ę��Gq���y2� �9Q��!Ϗ���R��x�z�o۲�%�Y�'���<�����̄�뇤���U' �(���tS�9)���M��E&�����.�}�p]ϽQCB�{=�0w���ux�������3Kƶ�h`��� NO�N��,�Ѫ�,M�ʸX2%Wf�]�W���.���o��cg��Q�n�5�44ׇ�w�%�or};:�O�8�,����f$���Voy�^iC'^J�pW�^U�l���w����%s�6�(����b����_Æ��xn�\T+�u#�����=}��
����6������=ݩN-Gv|y�����ҵX��-W �_��J��]��s'-`�K˩YlS؟���U��U��-à�$f�w��D�h���{�$fD�V���xK�r;�y!,�?{u�eug^ֶ�w�K��6uLg9;��'Fm���.��9�d:���d�Rr��l�[,{7�39��
�E��'5��{�G��/- ��b���*���Y�i�^%��2��c.��4:�n�"f��������@���F/>�u����`���V���# 1mh'��"}���	C��8�g="l�w,7n۱}MjY��!�PP�Ү����蒏]K܍���D��"�w�կ6{���ԗ8.�^�Y��*<�U3�_���d�i��3�z��a�Ԣӑ�O&�w�x�ܗ9L�D��P�2�U�}���i�5	���CS,�� ��i�4��%�΃��������GN{O�}`8UMUY���(:˴:�ծ��3�%s�T��ꏔ�?Tz1��f��}�TF:�&8']�ו�  ���r�,��8�:)�.};�IK�YI�ɽ�lz����	�X~����*�����<��)� Q��L�^�\�%Ϧ��S�#�'pxǧ�֪�k�	�kn�/�%�'���>��.�ۤ����&5u.����ĺ��9��_m@��X�"��lkF��e"7�}���`�Ƈ�c��~g�J���{�V��^�iWpt����n�vHx4״G�Y�@��h�H��P�i��[�7 �_M������K'�!*��\�r������@�9�a�o8�}E�B��SG]���Ҍ��}�����۩���}b����eeC�)�Uvv��t�q��q���FFa�q�҅������bBp1{��>O9�U�C���wr��[�	��nt�ž���n���2�3�!�>
Y��Y�����x]I�b��x߆�zR�8}���$�r��Ot��Q|��	�Xvt`�UΔ^�Хt����(���6n[�'�0u߹i��636�]5����V�K�����8i�"G���B~'X;;�z��t�@��5E�^Me+e�2����m��߼߅M�bf�\���s���?u��y����=Ɇ�ϽO�����c�z�{Qd3��4P�@�Ox�冟o���8`����o%=�=��t�A�~q�XP�^C�^&=/z��<~�]�9*mѿ4Cޏ>���[�.L��۽i�x}qQ�����K��>@Wa"	~LI�]x+���|�rg�T}éө�1�DA�L/�!y�\��`!,R������"*2����%(X�^\���r��>��*g#�����	�����/m���h��* NM�`�P��.�P����(�u����~�2�;n�%�Rj��4c_|�]{�W��upU�Ⱥm��b�w�	o�s:���Qj�Gӻ�/�5��֚��O[�`��[���,Y�q�Sފ�L��:n�����j��T�N1R�t�[aw��GT�{��g��ӄ��|^�lS%�走�YZ�2�n��W��E?��z� %v�nK�uӌ���wgnI�,��E:0gt1qy��ҭKFR��%��c�/Ⱥ��SN{�M�od��7��:�T8M�8>�Rz��������2J��J�����c��l��D�SZ=]������l��@�~'A	����^@r���*4�|'E�TK���#���7/�� lV>�ֳ�4z-@�j�!^�UE]tg��f�d_�E]�M��jL�c��(�cˇG#�+����4'�y�k�膖=�^�{O��ln�DME-�(d��x�����Ě��˺�^k	��%��{�b��U����d{O������U���<��y�V�Qi��	0�E�ǖ�1����ӈ_���.��Hk�:�b��V��ׯ�)n=I�����><]���x|k& ��,���uͼ_�y��'�:y؃��xU�e��>�Z���?I�����#³O�<6�x��ʾzz�;(gԹ�x{��L1�׵�9��g	9� ���}��u]�ܝn�/U�*�w1���
R��^��n,1b(��jڎ�(��_t���X�qnۗ\�X��)��k�,9b�l��,v��X�I`|OW���f;�:����	�ȭR�}�;vtL�]�s�b���%�Q�:v�߫�u�	� �x���&
�G�q�~��g$�*���1Md9W;�b��Y㶭�zoγݖ���Ȟ$>9EG�F��'�%�)�c{�pͷ��7�����\���x���>)v�]9�jߗOZP
ȫ�"
޺���Q^�a:��Ȭ�'K�|�����[�Q)n��2F�=01h+g�ǂ+�p�8y��v�X݁Z�7˓��N������T����2]=�yTH�P�0��JY;-cH��.zU�z��W��Ӝ�w,�� �S����i�_��\�_��-|��t
X��D!J��b�5q7�������P��!C��{X�Z�?��o����A�v�S�4��Μ�c���=��,�~S�+ �Sʈ�$B���a�q����5���Jrv���'w�&�F,4 �o$�V��D5�Ǌ�N�Q�!���7ؽh�h�CFs>��O�ʷjW<�sg��|����r/x�n��`Ox,j/�<�y��^5�41D�bnL���T�5�q�(���/t�>v-ٰ+�r}���e{�k�i�`&d��*i^:ȣZ�(h:��ە�{{��t��G�X/ �VK8���%X���Q��O�;��I1���Ʃ��ȍ7��CXv��8ŉ��5Zg+�������ݼ&t}ǋ���m�,�dL2�f��Vc�	fJ8������/��}����M�]bQ���lJxb�4* ��{�mSh�v���>����i�׬c��,d8�C���g.�[ͼ��+��z�єvɳ���k��zC���|<V�\T+�u#�򘴻˘�>y�����|��\�./w�#iO8��GΆ���j�<L�U�~��su�_��{�'_�ʕ�x���{��=
����dV����;k�ر2��=oJ^�wm$��}ZEvL�S����3��N�5)���vN�M[M�p���7��|6���V�w�U�䒗;��N����������(�w��rU׶���kJ3ᜡD��5�}�=�Ӯ��|
a��8.�GLK�mƵ,��dO6���H�-�g�Ǎa4�IͅM�-�5 4:̅ *C!�M*��POe[�8�>7�s�!�d2V]T�j���
֌8���,�E���R�e ���
Fm�X?)��V�mTq˭���纶�b�HM=n�k�=�c�V�~}~�y��̗��bu�w���j_��t��,l��.W5�/
�w�3;.^��(pF�[��Պ�|�W:�I�^��+�yf��3-���0��y��U��n�e�3[�,��T�R�]t%r�җ��=�wF^�iΊu��
c��w7�׵Q��w�^W�r ����,퀡�\�XɄڗ������E8HM�s�[(�vD[(ɷ�*��0�,�<<O[^�H~��7�7���B#e�0TE�̳(�FY�y^q�O��ጱ;H��(��d��- m��w�b�<X�J��I��R���(n�-}��;�!��hC�P��4����8M)�*A	�C6*"Z�|T��z�'v�E���z`����g˛"��u�]`�^^��p������h_�qI���^��o���-
OuL�ݒo��Uw���`�U��t��|�8d��<]rՔx:����R���%˱6�A���J��i��T�ߟ�
\����ƛBp(���W[i	��.���hV+J���.�x� ��.��Bx�n���-8������b�p�%.�\?w��<��P�~� �;��V��~���먟�ٿY�J�y�a��7j���8^��7'����%��&#ԡ���'{��S�3�F�(_�K����p56|�.<{N���ŭ|��qt�1�2P�+�\V��л��<�B����J8�-�6]\�oy�T,R�Qݚe�u������J�\�_ɼ���Fk����W�M��)|�f$gXcW�r�]�/yaj۱Ӥ{Z�]���NxƢC�CZ#(LJ=�DoA6��8�wv�*X����V�.�&)�C��ަw85��*mѽ�rnΘ���ܹ�%�x��JJ;���%�җ����
�%睇7���zA��UY�5�/����ַ�G��A�g��4�&�(��
�5�D�*B����%f�fS����~�?NL�����;5��}r�|�=�SZ�����р `�������M��s�2K��¤���U����)��Nt_��v�ej�e׭���Z�WԄ=t�³�8	�eUn��[���5�3���;%�>jQn���$5���X-(lvV���UW���Np�_�NJ����[�̞��/@��*���yׂ�xFp}�y�d�=�%%^lO��\��T��+��NZwi�y?#t��� A��!#0ҕ��Hr��шzIS�,gs[0�(�<=.���]`��S"������+~f�Q2}Qj�k;�5����,�\���6.�5J�����ΒE�1�r��	����/�=}P�c1�(���n�8,�~����
��m�]Ukċ�ڴ}�t�� })�������v�j��������l�{�SW[���{�Y�;�7lJ݁�%_:��:x�n����#v[j��8;�ܺ`Z���V�<v��0�!��G�u�,�+��5a�u,Z�Ӕ�qi�r����jF����ړ�:W��L��Y��#���k���Cߏ�P3�i;G��ynnc"�n*wI��zM0�k�gO�L�1[Jz��T�O�9���U-۬�)�ݖ@�z�緱��Ws�Uᗭ��� s�z�����|������P�lQ(i��V��6�I���XՏb�NW��~�4��Z�)aXr�/�h#W���R�[�xQ��VJ���J��;ټ�sƪ1d[�6wK|r�a=�^O� A]�
���
����G��=O���[�7�%�O�/p��G�ܼ�����{�W���H�b���:+�N Y��yM^�7�=��K4��sy��.'��iMd�=�	�Nq��~\=i@���Ip��q;���g�Ѕz��
<|���� ȿ>;'��F�;�H-|�x �̱j}<5ҦT���w������ߪ�k�{J=1�SH�����#��ڡ��
���z����b#�y�ꕲE�8م�tx� 3�e8����0v|^�Ǵ�N��7��>��"�少q��VK��5�*.�$��fފ��9�֭�]Lܙ�3^Yr�F\둘�Yv��l��V�	QaurX�3�q��n�y4kכtu�֓�hV����9o�9A���c�6iӇ �Ӟ��Ƒ��)��B�Cf� V��oOES��0�X�ё�7�]D�S�E�;}f��u�Y�(�u�*�l�k��(�e��9�/��%��ڮ���M�Ƀ����+;K;���J���6P�V��YM�����+�Ժ�gt���qit�����[��;z�ʰ�V��`���)-�v�h�2��LF;QS/d���DS�6�vSt4��H��('�����e�ʻ����8٣�f�m�������F%Ƶٮ6�R�3ur��\�\�4s�{��V����Bp��S{0]�s2�8Pc	r[r���ݤ�o)�f��\�4#��-���>f�1/j��o9ǎ��:&3��d�ܲF�r�tr�l�	
��#�)Z��+�n�^��b=�<�yDanV5_���6���ہ`���ڤ-�b�ݚI�>�,F�g���b\͌�j�n��M`�2+�-���iԨ��{r�cz·&5WB�Q���Ӧp��&�{D�;9¹��4�]�c'U5b�4d��J��o�^ô����L�{H�z��Yy��\�6�<>Ʒ�u/�塤�6�㈣U�jt�D���{lZr�iV<9)	m����\m>Qi�4�,��7Q�Q�<t+�X�7�$��^����R�j	���I-���[����cKH˽#�f��n�ga�����Ww�#:���7�6N�c�ڦ>X��o�4�0�lAX���*Ȃ�O��Ĩ^����𩕵���^�2�!z�YBIӄ��< �^���#�Ii�n�"�mG���Ȳ�%V�;rQ,���W������d���Y.���kxBH5�ȽMsx6���^Jowp�}"��]�5ͅ[]p\��s�Ps/,�a�1�p4�Ff����5�gU9�r�2��Y*��3��z�n�,Tj�aԸ)s{�R݀�s@�.d9o+�����hb�]ʃ�k�ݮ����_\��6�t��1tk��L��ܻ�f:Qh�i��jԪ$���YJ�*�����i��K�����ڛ�#fY�ƺo#����"��S6	}v�c����-�h�au�^����M�Х)Э�*͉Φ�c]eZy���j82:_ƒ)���da���Ź6Q嘯^n�Ѫ��sc��	R�"���r��sd��)�62-ܨ]ܩ��<�.��s�f=�]�Ѡ �+8b�J�1�5�]����&_B�{uL�� ��g:��7)t�e�m{4#O������aB�YRD���|vwQ˂ԓ�d��K537E��]}:��\/�w3g�q�W�r"����U�(���VU��A]םu�ȩA��i����͙�O��=�~z���J���h(ɢ��1Cv�EF�/  DW���11�42&Nu'wZ�#
(���1ˆ�(����4x�a"��׎DX�"%��fKמo#!���e#;��\�#�p �u�������PQ�I��K���ܴwu�]+"`�Iy�=u� �fJ��1`��<l�۹uzx񨠀�wp�%)�y/M��ђ.]'vܢ���q�����\�w\�w\܍b�S�Wx��wu��WM3��n#wp��1�WM�t�����H�<�&�v��Ɉ[������i(�w"!!&���wn�˹ƀr�TU�QKu5��H
����9æ���E�8g<���Y2���·6o��uӊ�q#��N�Qvv�ռ$���(���Ly��:�Qn�ڻ��ݾ���%
�]z���,�潷������5���^-�����ݱ��?��w^�r�߭�W�~v��r�r�W��m�y+���}6��^�76�_������[~����&�GF���2*���3C��?�]����b<���f��C�W�u7�������P����֍�w������_w��/B������ڿ^7���/ƽ���o���^/���;�-��>��}�~v}���s���w�;5;y�C7nT�?���m�|���߭�����y�_���n��y�E��˛����}>�u�o�����}����i㷍�m��׍͸j>��w/��_�}W�={���|�Һ�����2A������@e�~	ڼo�~7�����zZz�?=W��W5{���=u�+���o_�<����5������-�W��s{�}y��j����f�o�f�k5��?�����k�|DI���Y*8�d��x?��)�H��o������o�w��[����x׿�~o��h��}~~��}5�ޗ�G�����b+��^7��<������?�~���P5�u��+Ǐ�� hG��V�ox�Ѽd�s4;0wv����sn׵��_�}�^��mʿ��������m����z}����~v�[�\�{��j��`�O�&���.���w�j���x<;oS_C4��3s�oF�}��-}e��ԘȈc��r���5;y�3S���gC��h ��ϐ�W��C�	y}/�~��wx�k�^-?���X��[x����\�m���j���{U������v]׀���42+�{�L�^T9����Y0��s>�i��^;����ץ_��xޛp��μ���z��j?�����t�<Y���uu�@u�y���hܯ���ο�^փ{��ҽ-��[߮�?z������늿�3�kΫ��v��ı�Q٤?c��ٛ�r�{�������s�y����[�;�T[wO���s���3��1S�������~�����^�+�>a
�
��~�m������M�������������3���Ԩ���h�Y��w���ݯK�^>o��������~|�ܫ�6������߿;os��������ܾ�|�ŧ�_m����}�ۛ{����{_��<o���}z��{zm��ן�m�o�s�{���íbx�ɩ��D6�0v^.wr����dC�hnvG����?!��^!�����ȹ�|��a�[��l��0WS�i^-g����Wȍ=L:J�|���8/��N-�([�g#��)Ҽ/k��`q��/D��4:�H�>�4�
/խL�Y[�E�qr{�"��PL�^��	zS�t<)��_z�۟���}��59o߿�+�ӻW��sx�5�K�����|^��|`�}C�� �m
�%{W�ƝxJW�Ϻ%`��yv��������|��2*�r�����=+�W�k�C���2�%Y>T ���U�J���]��uJ� ^��~^����~
���z��>#¨��t/�/�y;6�\=#�Շ��ɭ������-~/������W+�������������W�湯��<�߭�U��z^-������w�zW����{^�����_̝��\O���������G�;Oy?���:�F�#3�d���dp�������ok�|����\�-��������Ѿ�_k�^��x��}�\���_���KO��ܽo;����\�^�;|oM���x���z^��W7�n���oj��9X*[1n;����5o{5�Z�H�����s_?�y�׵����~5����گ?/>���V�-����=y�k���7����������*������ݷ?�?{��\�<����Ӻ����������ٚ^�iE�5Q��6vx��{��Q~�_����k�����^�����|�ooֿU�o��^o_�\��6�����_��}�������ٚ]���_���V��.��ץ鷏?��=�ߞ_M��K|=7��m��?����n�m)�C�Uf���'^�ţW�;��_K�zWŻ���U��+�_�W/KF�W������o�/��z��ߪ�+����ʽ}��+���}���{U���^�����|m�k�z�����T/�U�ԝs^h%�S������u�[�;�_;�齶��i�דo���۟}�|]��}�����o���o{�����Z��[ߟ���k�z^-����������_{�-�Q��?�����{���`ȑ��ly�əw���hJ/�򷊹r����}�����_�ok��+��_]�Ž+���>z�{�7����^���o���U�������/kN��v`�ͤϽn�!���l
�z ����]���lʍSilKΝ�켂q㙡�����s����ѫ�ϗ���}�{ZwW���u��B��W���:@�kߔ>��~���Z/~��[��x�����W,|_�~/J��7�n��鷊��>h��A����K�%f����K����{�;��4V;���F�3��芾尛F`�Q�9T��{�s|�#�X��B.�׎��H�#(ʹen�G~�$N&Ʈ8�ޤ��í_`6���oJ�[tf]�,D3����/����;Y+R��x�N�W���k�Uw~�^�6�y��y�˛�n_��z}_>y��{m�{�~yO����>ux�k��@J��ĭ��k�@J򡨎�:�U�>��o����^6����k�\�;0-$�٘P��"N�[E�i�i��E��������oj�.k��^�k���m�f%CK�o~f	���N�N����6���s}��ξ����������/j�
>�*��~�yW�*!���5���^ëd�TU�N�d�7�/O�/��_=�����^7��}_�W�b)lC���_zZ^��W�<� h��|noϝ������{^�������潭��U�yw���x7�n���_k������+�۹����O������������z�|ow���m�y�ֹ�{��o]�|~�J��:�7�n�����\�}y��׵�?��Zw_~�|������^5�v��W�����������V�^-=�Q������ڢj�qՄ�u��������x�;�ͻ𥳐?W���z�^�}�o����=v�m⯋�[�_��{�j7���O�m�%�ױS;���"�fl���z��&d���x�sJ!�Ki9S��F9F����t��+��H�eg��6����ڑW�X^��N���F�^z�_D}�z
m�M'I���"f����,�
'����,�;.Q�#.]�Z٧XZ�M�l|&/m�롫��@	ɣ �/�/A�˃�+a�QO�����3����ap�q�_h��.������TA�B1ô�h}M�XgP�LN��;��w��Y,��H���9J-�1�D��qy�P���4^*�B\ �B��n�m��.m�t�j1�X��t�}�`6�P�:{���˖[{�I{ҳ���ﾴk*�n.R�:��ܥ�Dd�뙚t.d�y��/甪4Eb��Vy��Lͮ:[c'�s���L��%��T�b��*�S�@�Sk�N[;i�TЀ�t�(�^
��r�����g�(�$a��;~�IL�n��P��{�����DLH�t�  D�!#0�u��γY'F!�/ㆌ�+X�m�Ƌ*�q�@ZbT{�*�����+~d�0�=��xZ��\(d�u>�Oj̞�t�	t�M@���8y�%	��x���fQZE.����|~��Z�� �m�U�M�9���ք��l�&GXk{�ƚ�U`��L#x| ����C��	���"i���^�(���Ш�KMQ�G=��g�o���c�:~5Rey��=E�*~o�vk�5�y�u�NX�0{=3�d������W{�e��3����$w�=�\/�m����9[��gWOI.uo �l�Ʌ�zZj�����6�����h^]d<��¸����U|���vP
¯D�ݮ�j�i���?ni�o�e��v��S �x��ފ�%�
��k�g�wN�bk˗X�C�~[�����'.�b���t>N���k�Otj�>\@��!�T��^��C�+Ks�{{��G7yk�f$尚m��4��o6�i��ÜF�a��5yNU��8cy5��Ld�F8��P�w�������8xOQ�hG�"
Գ�ز�v�����nü�7te��PꝪ�Fd�j�ݲ���W�N����qhD�DK�G��3�k8q�H��~����uCa��c��\��(�������2v��,G����e�I���Xv��H���tQ��y�sy�<���{��{C�xz�W�l��uڻ���������[J������>.�TH�P�x^�Y�P�ɡN	���?+��rF
��M��� '��|`S�]8ӿ+/�K���nfp��l6��ƛ�dh�M)�eG�(a���F����`kA��:�@G��������Fo]�ؕ���i�(�D5�ǰQn��6���<9}A����D(�Z�C��5uθ,�7�U�'0���MIᰨb1*u´'8z!��
�N*ڈ`����`=������1���u��#��0_^|��jL��{��x��ɏ2�3����r�k�s�ny>Ӣ�_^Z�x�3�R�����5\�7͑Nq��/��걏|���)�We���ڵ�.�A���"�k����AԠ��mſ��[c�n���V}��������Kڇb��Yb�Z��P�G@�5�ȧ*��l�;M���>q	hn�ь!Q^C`|n��+���+�R�A���Ol�bW�C6�ۀj�iT���ɠ�)	bN��m<O�j���X��{`��+�Tެ8!�Y����&�k*H��c��2���^�,mw��j���g��0�#^�hp�q�c��������[���N��N��}��+�s=S�n���>��7���0H���Z�g㛊��0�#�6W .��z{�h]�S�~^m��7�޵�5'��y�z�w�Zu�[��k�k,ܻ�\b~L��I�Ѻ�d��,�>`]�n���z����S�����1�Нt�EN��:e�}�q��7�U���'�i�������3��p�<���q�U׶�5�i<^�r���d�gn�E�L����z���x4���^����Q�T�<���lK#���Fia���wz��S��+�����DO�
��;�R$A�('��v'g��3[���>3�-ݚF�C/��+�\X�J�_�r`����
^3n��~R���V5Y�&��K7�Մ���흦OL������#xߵQ����Wy��g  �U���m���E=����\��{��c�RU�h�q��׀�W��B]z݊L�D�u=m{��~�G��vP6ՓA*u#���z�Y����kQ&���[-��:=��eF&����H��gxu�-�"աY���t��N6�&	OV����}�k`-����J��4�`��A��fQa���oR�{	�[8q_s,�6\��V���ޕ̓8hy���rHeW�>�n)W���oϘ��E���OL�- o�N;�6�����M�|�8
e�j�:aȑ:�	��5�&x{��٨�N`�'{G��fU?9L�'�]!�l}$�`9J�!d}�3t��*X(V�������\/3����v�,	��<^Ë5� 7�������V�=~+�}X�:�F[���Y�>G��u�u��\j*�Y�kѺ.�Ĳ�|�3N���c�<�o���SՏ�[�)u�-�k����n�l��L�}֟�r���D;c�	f��ׯ<@6+۪]�=Zo�L��ƺ�e�<�6k~�F^�=2wW��T��ՆL[����!�c03���=�R>�u�7�S|��<���M5��I�s��ݞI�ݥz���j���peS���O ����o|h�E�.��5�\K�r�区G_f�����u��e�
���z���9bm�grr5CRQz���
�B��,���:�L���_�sE*�v5�>TG�6T|.���n� +���
�g2���/�n�-Ɵr �ut�V�*#nrN�[���`s&B����oA��}g!_:�;I[��ĉJt|��A:�T��d�th�1���*�w+�y�4�p�]D	xU�p4�P>hf�ќ��t{i�=��� ^d�5�(����_� �}o�#���_Wl(c�,��oҫ�@5�@�� 4�=D\5Ι]�? �����Μ
�}�JP��b4a5�f�����)�G�� '&�J�<�/v����n��7��^r�� P�UF��$m�&9�>��u����y�åx�t��r�����92۽Rds�]3�%UGb��Í�ҋt`�!��^B�iCc�2�-M��O��ڶ_G���Z�=͵�x+��[μ�0}���� ��g�)~��G�EF<�QSOo��'�g���ΞR�����>:H�5���~?&E������Ǫ��ʭ�^�1b�m��	�T;�;�	��aH���_Ո:�+���e���ۭG5-�ɨ���[5�:p��'|�)��hg�μ�#��C��Y�k̙/���`�=���:�R�F��?n����w���x�Z�m���@0/Y�qS�o���w7�/��{����2�m��bxt�d���z��O���3Yo֏�2}�m�j�d�gv��[�������T����e��r�w~h�Y����[-���9Mun�Mk�zn�6���O"����yL��S�'�U�hq�B�z.=z_c�9�wjԵW�~��>�d�ղ���|�����!Q��QsLۦ'��/�������+b�Qؚh}~[T�5w����T���0��������J_���-�d�����١��{9��.C3�O^��}�TF3�Y�<7O��8����z�e��\�}C�},����G[���ز��Ѿ�o�S �~+�hi�BYЩq��(���%�H;�LT;�&����~�+º'r�Uo���{�W���k��>�S���Z��P��֛Zkh&fv�r��A}�2�d1q,L�(5�2��B��u[�q���б�K6Q���6���u���� ����(�γ���3���[�d��Znv �e��3�J�:M�z�g�'� �j�L4 ڄ?��%���8�������Ը�� s�������|wN�o�48�h@N�+�U@� ���g�8mq�w�e*���Z��J��o����r���劚44A�ZP΄��΍<;���tb���j��~���ԵF�o�:H�7��):��IE��'��w_�<h�q i�}�d�н�^�xد_W�J�M5i"�xӾ��&U�;�}��0�U�{{J���0������A��C�s���`�(��ު�T�U����Qn;x��:�^��mwgiy"α���z�Tg:!ZB���}$Cv�ꭷ��l��:��QN>79��{���9�m�2�5�#g�����we��J�p��N:p��C[�T��R��"�N*����������q�g����Gx�8;�|�f���J7��{>��:����ezX��n�5�=;��,C��.�tՍ%���{��\�ɩc��`6ُ 	�Y�^��??D�g�7�o@W�cH�lQ
u�=0*��Tja��|�ƴx]��	#�U8��D��H�v��֧��K�~�2�������z�UOB0=�4}*���k�_\�]~��7� ��\_��'���B��{˷˪y1F��/��wM��x�!�V����yz����N{wv��{�%��*� ��\%E�k���Xul�׭\䆢c c�[�X��{H=,=}=�oT����m3U!��~< 5Ry�yxW�P�>��{k����"[)�윶�X^�I�nچ���	h�iH��|����<lCωRP0�}��:����*b>�%GLâ��>��X�
��Q��>�3�`�j�yU�9�׾�%v	<�{:�]٦U��ǲ��θ/�S)H�Z�:�j0�6�,�q'��i�mk��L5d��Zڝk���cc2�Ob}� �)��En�#�7e��eR�/a�Ȯ|ƅmfov#��ue9�L�z��#;&Eng*�ޮ�n�5�/L����R^{%��c�x����bt�J]`̊��N�Cw>{)���W��+���ڐ1b�t���qvU_h9s{�[��I)*�io&����R}y������u�'eh��2�)V�ְj�b$��!�[Q��]vfl�/{�Ppu�x�|j�ox����S8��s�l`�	tǝ�MfRT�5Т��]�#����C]=U��e�F�R��$��+]��
�T�9/���L$ɭa��o:eԵ��s�&�A�1�kU]��n�S�^�1�|�R�\�
��(�^V�[z���-����<L��s�b�"����s�(��C���:��-s���	Zܱ�uk�I�)ݍK��Ua�LTZt��ƳWǜ�n
�ҧ���
�ʍ�]��9 ۦ�jW/8�.�WRB�B��H�_6�6��{����&��RL����ԣdѺ�ҷ(Ķp�W��
�0i��Ejj\Cn�@2:K%j����ԁ��5���C,���
OX�b��V�]��NS�2�L������̔k���u�^H�X�y��c��]�5.�I��J�MV���0��q�(�>�Q
���%<�9p��#�h㏩_&�{�d둲�u�Ģ,S�����Z���v���sq�Й�m�Zr���YF�V����*���\4ֵ�7xo�����eA|P�v� \�E=(���׷0.2W�OT7b�O]s�&�j�Х�"�J
�����K����W9�H��Z@k�ߍ�Q�3GY.���m;��L΁�!�"#��q��-e����4��`��D6�	�T#%էy�����sr��[CL�^�+]��j�Ҩn��	Ԟ�r���|t�����K�1���l�ͥ�{�����F��b2s�C�b�l��	Nԡqt3��:�]�V�E�u����%�{Xf*�;+y�/t/�Z�T��YŚi�%���={9�h��7���N�U��\c�M�1cH�ڳGW&J�N,o;a�iN�hd"�˜�a^q�.�Cv"��ufk�kuC{�{g�p�X""�cwU�Y�c�c�X�b8�tZx#tԒu�q,�����Ld�.4�k锐��wR��jEZw�ݪ���ioMB�9}�ԋ{(.v#�!���/7D�Y���x'e�!�;!�$k�(�&��w�	�8U�`��]����3#�8�.�k3Gk�r:���ǯ�`8J�nvp��Z�;*Η�{�gS]ڌ�r�sU��>��,R�f ��d�39�ё�H9�,nH.�	SmRPM�uH;���n�Qh[�S��<0&�9��*�Mu��!�1����2�;T.���6��fv���\9ߟ�wv�6B��-����$^u۹����b6��F�utɓwp��q�;��\܎�ƺ������JS��(��(�.t�ݫ���:]��.cr��#���������û�D����A�K�w<�sx�RS�)!���6JD�P���3���I�b���WJ�E�&+���仹%�m�n�^.�����$���u��t"�c4�F)K���H���,#��)6��%���ۮ�@2wY�ؘΔME���$�y�`�]ݣ�P\�L �4]IQ��0��4.�5�:�"�ИS�q9���r<�wsSx�d��b,E&/;���؊�%�p�� �ka�w;\zo�	� �����b�xrݔR�ٌ�����+�nt�;�� (赔� ��V�7�=S�	Ci{����y��45� ��=��-�;l��x��\;Ǒ>� @�</�iWL������q*��v{y�sgGu�Բ^P��ĕJ�6�AN̈́��
@�U`��*c���n�b�ߙwL��VU�]���͕-�EB�k̔��>�D^�1�>�k�� p�͵�����&yp[=�~�f��:l*����?�x�Wf;�p^�U�{�-ʯi�
�e"esz(�y]�����9;�-��H~��'�x=к�
��t�qϼ�A^&�OJ�zE�[T,!��@���{ݝ9lZX��t��ȑ��cX�`��GC4�jN�>5´�M[N��=��Qz��K�*���� 9�yy!u�b���R����T����j���zd>�uyXT��u��wq�j�D������f���u=�Qs���ʯ&��<Hiu�M��@MA���x匝݆	�w����x���ǖ^�WJ�����;�xgE��#���=��g�Sy�۾����v�hfF�g�N�vO^�2�6��u[�2릇�=.�ǭ�њg��aޙ�Fs?Қ��>����Lڸe�w��>�E��k��e�K�	_�1��c�=�^e�B�ӑ��"h�ۢ�l�C�)*��UgS.�oM���<E�K;0n�D�!Ñ�g:ɳ�x�v��H莾#sfT�p�#oP�1�$�{�������G�� .}��K�7���U
~�][18C��|B��N�x��R��7�\�6{|��q6�R�H�0�g�L}�3I��\U�,ʥ�א/�p���'Ŵ�7ҕ���O�'�7�,]���4���hP�+����a�ש�<G�bc���;��x������ZclyFB%G�^�К�!��y|w"��}|P+�R'�*�f*٢���f��oU����%��2�.��*��SA��.��4��3ֆ*h��m���=Z�`�˒9�#�TBv�5�4��qL �~]f�?>_S�|��e5��EUt\�d��R�Ś��ݢ�$�ۺq��zt�8@��U��H���':-lmV��̪k�!�;����3�=��=�{8�@��JCǯ䀈{]O�
���l{y��
�&`�^��7P����>�o�[�Qޤ�^��X����n��\�*�{
��`�����I�ෳ��}��ma�\m఼�� �)W�	�x�#l������M6xy�Ul =��R�;6ŕ;��v�t�y|��*[��EC���yk�7Y<�s�zi�P�n���V�Ԡ!Il����Ր��DxI1�l�w_��/���*k���MJ_M�&O�E�3����ɷO,m����(���u��*�lG��!�2vQ7u���Ȏ>�ӿ�{��w�.ﾝģJ�;��)��	�U�v�xb�?��R/��>-@��h!xD1�^��vwWW��X�CZ�O^�٨�`�p�'|
؈��ea�=�Y@�1���ʫ6����6���e�`�,�3ZLV*A*+λ����grB�9/�z��R[�O�~�ǖX��v�qU���2�i�`1���xs�y
����O����-M(���ĭ�Z۝�R��-oO[��q��5W�#<>T|`�]�^�]{ĕS.V1�_�Wճ���J��������u����xйx�쇆;O�^:��iK�
�K���'A�K4���\�6�~�-�S%Y���O�4�Z)�}��f��\h+�2���!�(#�d��zyn���� �U�@)����\��](�;������Otj�>\I� G!yZ�	����_/���Ƈ`�g:�'��.��d1q>&S��Oʳ�e�
3�E�V���q�x�.󮶐��R>�У<����qB�W��t����T�u�B2��WlP>���G���,f�p��6���bg#��]X�ܽ;���}�*��m�4����o{h�{�AdkXN�<��;�J��NQ��V�>�g���:����vM��� �+@ �4R��`Y��]��جT�m�:e�qi>fd�W��x\��߰ܛ�J.3��:\r9j�_��!j��r�iT�C���>.���$8�E��Q��Ɣm �+�h���
�֛g���	�Ep
�� 3�c�!���S�e��P��}Pf�ѪJ��S�zяk�N��SF�g�1�:؍u�@@�k��A5Wa��t}��G9��àW�t��	\�����IN;қV��×�P����^ښ���o�j�}_��@ʫϺ�<1�n� 	Q�d'8r�N�URpW�*�[�e�1k�-Cڼ��eӃ��ԫ�jqv]M/��^A�j����p���^/@o�D��� �J�ob��߽�ߐQ�
w�����>g���P�W*s۸+Wg������|�ڇ�W��^���~��cn����B�z���U���Á�Y�WZ|3c��_�<7��ã��f3�ӎ'�^��;����,Oj;n�����j��B�NW�c���1���ў�����>�;3��j�<6T���O&(�y����^c��#&||�a����^�p���XҠ(P���*,Y�8U�0FP���;�A����{�GyW�5�z#}��7:��z�;�^�-���6�,�wԚ�<���:��1͕�ؕ{m��T�b8��!��a����:�;��W�Y�=���w+�EKC$[�_l��y����Q�{%�#��[_��41wq[����&��D����>���mʥ�]��D�t�Y>�|�B>��n-�(���+�z޷�隯B���� ��<E��d�Τ'�JX�Je���[#f�*�w�7�x��縏
t<e�d�H�i�O�<5�s���|P}�}�ʣ��f3{��J����{�µ����h�*�t
���Q�m�NYUe
��U�^�^݆
V;)�e7�7z�0ϣ%#L���#�ϖ���0�a���pi('��n�(�#�U�WmnDYrp�2�iUm�N�W�:��>b�*g�|m�L�k6�b�zˊ��N��Ĳ0�b
�����$Zܴ��U�r�LIPi����D��¤�*�b6oQvƋd��K:9,�te��z�K!���!��2��M[���E��ے0Ӷ��,4�u�nwma!k����vW�DMײIޚ��^�N�Q?��=�I�Q��Nճ�5�^|��/$�|�J���#S�y�@Ķ�OW�x�5yg���M�@ײ�]���ݚ�V-(�����SA֣i\[��
���坕��J1r4�b�6wL�FP �����n�/z}R�˗�D*bn+���B����g����T��a|^b������}�.}�J.�:�l��B ���*-�í���9w^��&͗V������:����W��� �k)���lMm�\V�i�%�f(��DU�bkE�-�K���\5ę�S�z�
P��{���K�xh�W��YC�4��jH���8d榍7-or֍�:�u6+A����QLH��`�ո^�a�gҼ��3��T\��e��`Պ����u6�b�jl���ڎqsQ�U�P��x~7�6sG�u�#�~pX�"u�/��Vw���-5�z"��&��;�����uQ��_C������U�6�H���i��ɚ���)8�^�qK}�s������>��c�)�A�nS9X�Q�K�	�Sd���hEm	�1��>��1�X���Ϙ,��5�&����g��}8�MI��Z�'���ꇧ������]Յ���ٺ�j�m��Z =���:�c����0��,t�..�@+`�6N�+��m�P�=� �0�����)�h;�����@�,�������� �Un�B"2,a3D��B��c��@��i�����CZG�c��"�ޡ�*&�v
��~��7���^}#��`���L�ҪgL�;tN#��{>V��t;�N L�<�����q]�{�==Zm������߳P����jT�;�E�����Z)����C���[��^�F(� wڝ��ml@Ê�ӔӪf���8�˦19��ԉ�FU�-<�KTW�<�D#��
���#ݶ�w�#�/�k��$e&��+�V��A6*���Rr%E��[L�H^�c;��g%,�0w��
4�O�n�U�nȖ�)ĲI�Vz��?_�ۿD����S[�G={��_i��W,����&�W�����J.sj��j���>���S#n6P�i��m�����t+�Mi�jzN��/���u��E�f��%5�¦�ߝ���s*���f������>],R
�9R@���|VM�tt�P�oثf�\S�`�u�n��A�=��E׹唨m�Xz������q�d"��G҅}�H*����q�V&�j_�y!.Uy`~�*�ٔ�42��n���8o� �{�������M�2��ƶo!Cʾ$R{��ۭ���S�D-��ju=®e3W��+xAAϜq0�}��33y�+�xӨ�ҵ�B�g�i)7���?/sɿC���;�{�Vr�oeR�$���L�L��Ym�-�u V�P�=�|W�d�=��ݿUϔ9�؞ҧT�LL��u�	�KX[6[l�,�V�"�0W�����Ĝ�F�N8+V�0���2��h��������S8�]����|���cZz�T�iay+��4�a��F����3uW�t�1�����^���"K�	���>��׽}��}6�Jc�hB�|GF�n&M �S;�SX�m8Hi�3U2�--Ǖhb�1l�:6쎻hsmYG%��܀�VQ0��#Ll��Tչ�;�E�I�<�,ie�L@(â*ܹ[2��ڨ�Q!�g��P�kU��n�J�T�ZuLE�I�e��M��	�@�9�Pм���a��p��ۉ�qi�6nH�ҜII�l�)�[��'�u����l�Ţ�,��p��&�Wp!:�1>�cr��[$T�����R;��߼,W=���Q�.DܺRabR��ě��:W�h[�V��k�2st��w,lf�9���^3ӎD*VmL��۠:z'z,X�.�t����d�̵zzo7˟9s#�����j�s���:$>?G<�`����?�z�}
� ���)�s�q����}%$4�'1N��l?���E�c��3ʎȏOfy�r­���)�Yd>V`�V�!-JP��Q����8�f��).f�E2�WH5���������6[b�{uj��Se����X34��L��q:�ӡ	��Ŧ���2щ�l���Xlaj��j���~շ6���Snl���ȕ��jF��.����	��Ym�Ya��5��
U��U���=S���u���L�w!R��t�ƥD{U��P�T�����z�{J��Z9�{/��NG�ϵ��5QF�B!ΰ��e�nϢ���n�!U��+^�
Kx�g�ϻ�OE���~e"���5��k`��`/�w�_ae���Յ��^�;&R�E��e��U財-g�X۶�a��F-%���n�U�>���_r��o�x�}�v���*�.�|��g��gȢ��4�զx�:d��q�1�>6�ӕ2����3s,k��I�I\-���	���i�������/L�A}.�zq`��N4�j������+8o���=�zu��$��?���sX,ƙD���-n[$���йe'���{ȝ��pujbC����|ϨW6�K�B|�r|�te��x��m�I�Q������h�Ԙ�����C���H=
��iFv�X�W��I��=�%֏j6S�k+KO�B�r�Ŵ2Tbj�/!�j�Mt��;�4w��j�� �2��I e^�.Zν2)���RW������)���d��㹹�h��=�F��Q��+dO�K!)&�\U�&����T��K�����-� ʹ3'��]5ݤњ��6���T^^�B�!x�d��"��"�y]���[�Y����4��h�>閊W-
���G�0΅r۩�S5�Ck�kM�+d��7�����Y��}Uiq��G'���*�Ϡ����Vxy�t�zW�͊wZ�w�=�q�o���?�o�-����ldu�Kaf�q����=7ln��y���P�t�8���]
ޛ���t/0+�bd�;D����a6ᩆ���e��{�<���ĴM��n�,�ݤ�,�,&5W!7{EGp��=)���+�^tkpt��Vl�)0���K����B�ܸ)�:*0��D��:��֔�cۃpM�ycɌ�*B�y"k{A����"��3tX4�2�G.b��8-�DԎ`�fFU�)3[Սk�J\Uj#`N��s^XUC{`��K�+y�$�EGoUz"�oeg.݉�q\�1����i�C��`T����AY�u�F�ͅf�����	���V�C�b�v�q.^L���.!�H�x�����Ѳ��S��0bD�Z�fuF��mQ�X�P��\T��noݎ6+sƔ�k%̛���Į��g]�wq���H2��^�<��5j�h���"P�����:W�ˎd�&6Y����co���h�Z�R�'MaG^�&ͯ�phIXu���;H��ꄞ3��4�F3d��]��]����.*��o���$y�n�&\u�T�$����8T��U��� ��Oģ��R�Q�m�(���X�3�"�K���	�1��ʱ��<&$4\�0+�K;ZNn��e-���C9m��ͬ��h�.�/�tW�2݆^��<��x��66:y�h��
�7\i+���b$�&9R����nN݁��1�xs�����3R��|�u��ZS;�5ه���R��-��D��ê��8됆rEf*;��S�
vh�PM��{��ꌞލ�簚��7�&ģ;Q�Uv*NX��)k�v�W�������N%�jŅ�cs���Ъ��6�鶠F���sr<���ih�^�W��6�����!t��#qr�s��D�����$ח���-�G(C"P@
�B�<��E�o�Cq�dл��Ps�Ǌ��޾���o%�7d���`�`I��B�A�_6�'����S��˗�WM��4/gGF��K�+�����˂(���3����Vq�f�vm�[+�M���1��ۚw1�\ aA�>��ݮsF\4��qL��y��9�N̥0�Fk���7���2�8���QY��T��X�Ƈ=�:��h���*: �;�j�r�Q�&s-n)ܼ�ou�+�9�(�#�ԓ8�A��H�Q��u������mz�(��$Hi��-�z��&�Gw9�i���(ܩ������Vު��d����E���:нXn�>in)_�_[��{�Qy�V�6'�WT���q�Yz�����{R�I�o9�/E
Yd� ɕ��'3����U�3�g.�^ٮ��u�[����������]ZW/5����w&)�ӎ�2��Z��ɑ�@vs�j�������)ٜ�ʳ�t�Q�����Zx-���ޅ�03u��K�&(4Q9�:pM4²�X���;ա���n8uy����6���.6^9��9ǽ�v���ׁ��P^�P�H,#4$�r���7N!���v���Nn�uӕt�]�]�wnp�&L�\��iD4L��-��9�9�y�7a��LfK$`4d0�Oe��y�#���"�G����30��뻼bm�;������r��	�]�O��H�H�% h�Ԓ2�w]���I��P�.]�$k��l1��F#<w+�4���0�wvL�M΄��r����4��ݐ�d�2g:`y�xFH�!4!�r�Y�S"H4F��&�'w	K�dP+��Έ%�&���FIQ1����n�#�h�혒)�%���B���� |>I��8���G_M���� ��U��E��jd �����zWT��M4���;q觲VDJ�{]Hm9�;?��xx����|�d�o��]A��Knm��6	�Qw?X�?b�k:�w�ȝ�W��������55�+ZFz
(�*ZEnn6����@̫��O*z��^G��~���8��M�z��1l�d�m4"��i��nd��ws0�Y8Uj4I��ܨ	K@ZjF�8h��Z�%^�uIb�4�����>��M���},Vu!RK��3�L���8��׽0�E�bi1�nΓo>ހ��-v��'�Xq��
�BY��)X`����3��5SQ�ͬе��(���+CB� ;��gmsbQNv�8��aWi������$��6U� ��2�RXҢ�H0��s�WN������(��O'Z�l�z��f�J�T�lU�-��O,�)C�D�y.��m��2��y�u����Q���_�Q����ҜJI�W�����5�~�`���)1w���ܣ��Ն;�o9L�e��
��*�xCE�\�^dޞ��Ӟ���/U��"5������֟V����G^��[�m�<6����īn9�U�}��������-�7��o����Q�(1��[$>���3{��d��-�h�4�!����䊏���*ʦyc�����Z�
�d��%�RH�,vzz�5�C�}�m��dHr�������j^1ޞ� �{�U��]�y宻ڷi��K�㪴�����+Euuzon��d��d�Zaf�{űnQ�hŊ�}<�}�$�f�o/�0?b�T�d��1E(�X����,��ǲ7S8��RqT�E{�M<�=�bBc�6�x;����:�e����w,��Y`ۧP�^mO>^��w�Hr��<>���'B���9��`n��6�m��ZqB(�d��k�ymqk"aJD@��;�i���|5���?�����!;s�T�=��zk�,)T[m�q��$��K_,zap/������_#�=�z�����Q����̋)�b;~�ת�V3%)S6
u>8*p�c��P��R�~kB~4��@�7�=���ُ~�@�I~��~�0��z�ɰ�\Fos㜌ĮM��W7XSs���c i:)�-<�k/b�s�0�s�.�db����Y�a����)9�=�Wv�����A�vx��ڼ�C� �Q�	a:��fwfw�o37��g[�eQr+�f�}��i���in<�Z�[%��#�v���vY%�xΛ�\��\L��gU�?I�J����4��� �-�3���5��~{��y��l�
�C���C�����!�J�T��TE�\HU3��E���<(�`�L!,9���2�mF����<
N��f]M$0�ݍyN[���(���Wu*o?CU�]}x���B�C�+���������r{��0 ��h���Y�E�jlR���Ϙ��n������QS�^RS���=M�F��z�T��ܦk��R�/(�oj��Ŗ"���W'u���2���vg077���%�z�Ǯ0��zmիC6�aSQ7S�7Y�/biB���|Q}�)z��І�����K�-CM��%K6�m�j�h�{�0g�����^b��0��bF��b�e�[+X����������
͊3�u��h���M��}���c�uei�C�x�>��K]q��:�N�c�;׋Xt�>�U/q0iJ��girx�����3�u尤����r��5+��r����F�`���:q�F��r�S�m����ͽ�������x��Q��l�7��� =��gZ]+gR�UǴͥ�����ˍ�he���h��^�y�XI��Þ���c��84z��'oЩm��n"�f��!�m���\�I�֩��N�z�U�To�c����`oM{��b�u,7դ7�C�~��_^_��7�zs�w�Ǘ\��9��ٌގ�&
ze��:nL�l�̙�͔��b�4��)�r�Q�&N��R�޵W��5�{6�*\��^5��h9��U�F|C�h|(K>��6Ͱ�5�Ot�)�S�"�Щ��h��|��7�0G1�ȑ��L:���0ӊ6��U��7]��ұ�>���wX�{/6��O��`D�V*��*?��N�6T��ƒm4Wi�棺���RN�ب�b�Z�R�m�i�2��@�SM-.$��iF�,LBj7�NnȭL���1r͉���S�Rة����v'$(��lXIV�]Ž+�����Uv�n�f�X�drr9ex��5�=.�ΩZ纉2�B|Cc�e�R����7p�97ʶI5���̫�Wmd;��)뮜���[.e)r�v�w��6�F�nv�t�s����ﾯ�Վ7�>=9q���5�G����O����R�2�(�MQ���[e,����K�E��C)����Tz\U7ƪ�4�=�ت�!�2ՇQt�#K��j;�~ˎ*��]�r/�ojN��7��:��r�':�9[���M�Z�;V���i��\_�^�E`�t�oz��Q`�����[mJ�ј��Ti�!��\Z�"S�5x�m�7��0|�Ew�嫅�6���g����4R�Fm0�:�4Q�T��b�|Q�ڒC��ע��%�]\l��H����-cv�[6�B°�Z���v�T��.乯��!�=D_�������5,qr���O���y��U2�%��[�)Z$@�L�c6ݵo�����3J�L�;u�q�q�F�jPiN!3$Eʙ&��T}�Ck�j����ִ���9�v��B���r�K:bQף9OM!��=�^�x�bk�U}oIPT�.����n�6���:�$�;
P�p��9Zנ ���ou����(I=��`t��F���V��BM��U���b�+�^Φ�&�o ���3��P
�[�;��­��w������4��`ڭW�Ԋ��w-��ǖW��x�a��Ƨ����W C��[N<Y9��-hWi4d��E���mKt��E���+le�A�%�Ý�l�Z����,"�ȧ�k�>��z}������$�u^A6*���*�όR�a[н{We�<ν>\�%���^<��a��
�y|�#gzǽԻ��'n*���f'��>�Y�+ޛ�~�"Jy�C����!�����:�+�qY{a�W�=	���
�'��]Տz��Өn���c�v*{�n�{2Ky�H����[�ya^�-���!�j2J��Ŏ.��Z�W�����E׼�C����z
�/o�W����:{_��'�{Vn��ok�{��,��A�́泝�}\��)'�<����+N<6B���N*d�f�jۛG#k�l������]�l4�w��ޭ����;����m6�Y`ۧP��U�6�0 ZL��O�P��/O��vCe�ZW=!�QՋEE�	6"�w�Js���'ML=r�z�u�]��sT��S��R90:×�1�f��pY���ml���]t����]E�\ؼ��\U(��&��t��Y�X�������"A�e�����������iW4�e��y�)��`����l�� �f%���AϜ)݃�jd����Y��d�}t��s�(�.qg�zu�39��y��i�Bl5�7x�Qf�{���Ⲽ��@�_Z��]�!�U�3�y���XH���sm+G-5bW�҄��:�v�,5�9��YW{Z�B��E�lA	�Եm�DZܴ�Z���?y:��^�jxX�:/�[�7=�K�L�xD���j�;�wX�ĭ��yIc!**=���"��S+$��p^Cާmc���Cj�Ƿq	�+]'�~�2?>w{0�4M�{��z�j���zhZ�o����b�U�Y�z�hh�;MIZ{g���n����)�������XgòG��C9ò�˜�M�7o(�AҲ�|�I�H�	{Z��]�w�{]^g���x' ��4��3�2���ٞ�;�n�ķV��>�'��t�Y���qz�ho�rWd��T��l��ݪܳ���֤�'Qr�DmJ���w�˕�l��oZ�{]:��[�m�-έ=��֖�Y��J�h̼Gu�6ɣY�33y��U���#�K�޵p��۰r��2JP�d�'ڪ���U�uQ
vݝ����Ϗ>OUd��kJ.0��z�n�Tء�7�U\T��ݤ�C�jz����������3rr,�Y޸�����}W;}�y7>�fe�� ����\>{�3x�W�(�C�Ѯ����I���I�)<�L�|SҲ{�1���N+�y6����V!賫��,�N��}�~Z�=��-�Λ�S�B(��Щm3��(�(D9�	�q�>�m��>���q2��_E�TS,u�̑YL�ޚ�nJ!ְ��=�z!Ȗs��S�wy��Q��5:d�WL���厱^��)6P �cM���YJ��KNk���3�hf}�>�9�{�9�{滯_��Œ���E44m",l#�6��;c��	�NO��϶>�����9v��gѫj�+�"Ee:��Wi�d�P|���,��ӽ�G���閬v�3a��ʪ��u0�j9�nB^ۓ�|��9���3LS%�l�׊�-�&\��o��amn�5�Jۂ�6y�)�� �2����:Ax��Rc&���œ�K�oe�������Z«I�[����F(�9�R�v�W���u��O�_8_��x��*	�Z�P�LFT��4��x�Q>1
'�aΰ�g8���ң�V*�JZ�)U>5�����Ԟ���:,�lT�E�w��UO_�����o�V�C�z���X���	�ݙW��%�K �kZ�B~���`G�$�sH�o^�~������5�"篒���/iOW���^�7,��A���aWMU��Q�L5ym��f��Z^9�C��Sر�3�d�?r���6����/;�W�Y,��*�Ǚ����rr,�w���N�O��J>w���L���ʮM�hȪ�O������X��$ǩ����Qf*=^�0I����޵�kZ1j���tk`�U&��-�kG#k�lL��\j���X�U2�D媰�I�kv�E22�f�m�C
(�*[F/O�Ԕ����)ў���4�P��Xj��P��B���^wQ��
�h�4/9 ū���w�q:��]m-��w_WQ��v��c8\����{\�5�nY�qc��7!�l���b�ol�K&x����ԜQ
Ŝ3"j���w{W'n�j����6�JFR�DоgR�d��>��-ja��*�Њ���[+ZV;^"�I�R[�`^�Aԍ`��Z!֜id�8�8�իԱn�������cgS�@�-�1����4.��s�gz�ܺ\g<��b��+9��Nm��XҘ��ϕ�j ���}��8� TЅ>�߫�J�>FR��z�{��a D-��^d/%�ꐴ̦|�ܑ�S½�T#��Y� ��!��r�&���L�G�����]S!i�X��)D�K0�s��a��Rr���tf�Z�/*暒��0ٸ����yب�hb�8�pr屰�
�R���t�1E�PZ��M{؞v,���\��kCM��Fl�l��ZN���Wz�v�2���������⾝ЮU�{���~h���Z�w^e!�U�x��MQ~�n6P�i�1O�n��ܵ�^�x�m�v>������蔗a�ژZ4�2�pt�7�&.���<��ޒ�8�2Tݽ����qV�ޏb���fdt�ᛪ��6���:�T���٘��ÙϊکW��[2�'���]1hÛQqfa@<�sk�b<f�(M����=�%��b���m�z� >��|rZ�H�hڸ���-��uWW���A�a�(dy+yv�oL)%^q�^a��	��JaT�FR���]J�_9���%IN)R�ҍ�`2n-9����e�f����6�>%��fʹ:�o^��m�c��"�$a��|������(m9i�Q}��֎�wĊ�k�Q��m�E�NjFm.=�d)tv�UƇc�KSguZ��GnEX��i<��c�T�π�ZN`TB�x�3s���ݭ�[!�����N�*��^���u�uv� ؽon��9۹@�����&����ެ�eN5ˤ��t��zyf�ƥ&Tʷ�O۱ꤕ�4X��h�d�J��������U��������v��ow�ȇ.VA��P����F�"��n��j���o��:�QC����%�kv��E��h.�̘�k7.�
E��)���H����hݘ#
Ip�� O��+.���X��pee��+e�Y0��G
wк��6�����+彥jiE�`��Y��vx2���2�s��VS��2�6��R�B�����H��3[҄�d�{'(��m����H�lr=6 nu>@y���֫���u�� A?bR�t�&�yw�\�l�3K�R���#1]�8���"�J�ݝm�^�]ڽ'��w4Dc��{+��R�[�3��Z-\��lT �gw���Sۙ����J6s1��ă��vmőw����e8t(��*�+���^�'�9�>j������4�os���n�iF'9d��Z���q×J����j��f�s�0�]�a�.Z#B;�\tnK���y��٩��J}#lv	�⼽3��R���sաvD���&a�W��|1oi�E	Q^�'���C�^��,ɇ�,i��6l�n/��ڮkj�75��8�xMKC�ʐN�æ�S��k��U\�3K�ԬGhoC��8�7��-j���Jj�a4 )읃cC�!��P��!Z{�Y��KF��)�����:h�@T��嬸����f�S4��m����T�6��ė����z��n����s�`{"��o5_VU��4&㬦ˑ��%�6y%�#X��z����<0�ѭM ^2jv���
�j�qIܩMg;�<-��8�e�͢��jw�Η[��r�kc����ʁ�L.���n�����e�EK�l�O�N䈧�����gfb�}GZ����f�%�-��}J5�\A�����/蜎8熇-)�Z�a��h5}e��Ӂ �>����ie��9�1�ɸ�����k�T=RlRf��>�#�݄$dHH�R,��"A;�h�#!�n�N�LɄL���J@��\�lP��$�T� # �F0JD�L�P!��]�:\1Aw�y�\!1�'u\f�&Y�D�ݸA�fI4䑅4N��A�$��.QF7v��A��ۜIi e$�'.�ܮ×�3�fs��A\�3�� %x�#2�#%2SM���X��PI$�ƉdHĒ3#��.r-��'u�Y����鄅ΣnWL	"��"�L��8�tL#$�2���svi�D��X��2�NuEs�2wt�wc���e	I�B32��t��q�C a�F9rI9ӻ�$H�10 '+��7��R�X���.X�j���o�;�Pb�;���<U4�T��<�����lc� fe_@�gX2h,�V�w��Y�"�;;N~���Q��G��7v6{w��Z�6��d����X���a��Ϣ�4�-��K6+�-'�1�E�R͝��{U'����<�~�W�f����Vn��![�e��'M�F�F'ٲ>>�Bs����OD��"{��,���a�y�"w�ؑ��,���z��e.�Rt����{�g�2f�jqF�c���&c�����1z�����qP;Α�t��=
�G�珵��v���XC�� �/A�k�^�Z�w�5�=i�qMH�U��'pc��BM�Za�(�����O�+�Z�`ɽdkzׇD�=!�ʅ�i����e��^�;>c)]#��&�W��)J��v�,5�������$0�\�N�7������{���FL�f"���-ǟ+CA�fJ1u���'+*!#�u�1;�6��V	�V�7�x�{�Ė6d��*�><���5f��(-Í�יwu=Q?�T�t��}��b�gfհo�x_Xs�bdާc#�7
�1��[���v��I�m̤$+�}��=z�GCAn8�r�,�uz���|iT��2R��u*��k���C���r���憎٤�Y�cG2��9>�V6�����M�}ރ�`���Y}E�����U�hJ�ɊQ,6�3�G�‶���zә��70 �]1��H�2�\"�g�	Y�T���W�2�d���}͐��g�Oi#yj�j[R�-ZY	d�>Kj�����T�U�Ϙ�`��w�w�E��`�'q�B��N,�Xxɞ{�ԥH^6���Ŏ.��q�d�X��̺�#F/>ᖊZ�]�e���ub��֫	�qr�z��#Iؚ�)�����K�f�?d�º�V�����D��k�{oۗ�l�j���)����X����ؑ�8��s��uGK��M�3ڟ6a�I�t�i�1G �=��
U�Zf���T	�n��̴�����us�,+$(:�H��׌ZI(���KH��(�*�C�a:Ϧ�\Ɗ��2�׎N�[DS��M�qҮ]�WWU�x���Y<.7�v��jw�4�K6K1O#4a^Y]�;��C���}�Ƕ��et��ɝN��Lܮj�ł�����[Y_`R���"|&h�7�ﺬ��;��tR���1Y�'rgm�����aJ�T��4E�R�Y��
�n��6��X-̱D:���+Qz4��1ɻ[GQ�f�W!�Mi���,d��]�,u��E�	0l%��1+_))Э��+�T�f;#,5�:��tL�Ӕ�(�1��^���'�Wi�c����f�~�=GJ�Z��y�}9��v}��v��[ƦzN���s� o����,�h�y)�S*%��2ڤ#N��qezM�E�o��fz�����vw�=-R����1T����l9�x�fs�(f�/��X�Q�S��)����߱�D��M���h)���R�؀��(��&
�al��Jp��.��ĵ��T�v�d�M����Ml���"�M*������cӴ)��Ƒ��/=��+�e�T�z�2ԥ
��Ô\�-:��)���=H�Eb%%��Gm�)��N_�/�{b�����̣��1z4�}��]wD�H(��}�s��v�j�]��}`�}S8��(�L�"��"�����_u�t;fjM�A�d�}��L�u�5n:4U������$�����{��Q�i�E���ȣS�S�P�������v�qkH��f�1�i�ud��G���c�wȳ��T���VB�?y����w��� ���*fJn)͵WE`̥Mz��NE�kĈ�q'�X��4j���c�F�j��S�5x���9M&�4�.�1��A��f��1-F���1����KBmٸ;6[l��n-"�
7�6�7��NOE���s�T}@����g�L�ݛSd�hEa��f���Ԧpn>�vz�����#��Q�9��sG�,���\��30+uJ��L�m����$��x+J���6�|5�3�{��3�m�Uu�����xۑ��Gn��ǬJеN3!n��N������0J��^�[���>��u���9D^,��|���S*$�>�쌳��6SD\$�(��j�e`L6�E3���[�wHZ�O),ifQJ'������?z8��c��K���o:e��o�8���"����݌�WK�S�[�}�����6�6����X}pX'V���wR��ˉF���R����m�ްn+���l��w2G_[�B��T�,�,ZamA]�ި��\�����1�t��(-��]\ŕ�9EG����V��A6"�ֵ֢�b,Pv�Ñb�(�C�ax�.U���O>U��*{ޱ�6U�0�{�=� ޖe�wS��/yW=��y|rEG����Ю��w���uF����7���RL�)E�j��n6P�i�1K4m���uUR�W�ihp��L�~���%r�1���ǆ��&�N�$|lS{k؎�M\��x����d~�z��U���Ԟ���󊟶�Y��a��Sdb� �/�HKΊ�EE��h��x�XY���J�m��@:WVM�����ﳹ�L�,�q�X�Ta�G�ڪy��S6��*
(ʆ9n3lNZ�:-A4s/�>}~#\�58�Ng����A�z*ޢͶ�]Z�~�+�}|ߨ�����Q��f��5(�2�X=i�qK
��Δ�����X:y�7f�T���F^�&�,���?\5�굮����/n�H�D�(2��c9TG��\p7����
�XE�a`P6����tMu�6��y1��@�[�H�(Y�;���{�5�X3��|N�Mb}�XI�<�х\�9�)�k�C$Q����ۢ{�px�&s������+(ťL�@ɽe��z�'1ix����[�3U6AM
����J�E���My@�x��m�t�<r��^}zk�5�-#�-�=cG�ҘG&��kr�+�ehb�1��N�V��N�i2��glu^�"���՝Ż�E�6�e���m���*��1uI�G��؀e���^v����]�Z����]��|�G�
�*S{�K����/R�U)��FÝa��q@�Z��1����u4�#��}[{"JI��&�^�ئ���JYn>Lwn�{e�H�W:Xк�-8m��&�Ԥϯ���o�M��Qx��T��T���S8�J�R�) �鳯�*2�+خ�Kf%�z�	jR�S%��`D� S�iL����I�pj�CZ�碶����g�qT��ߪOO/��&�Y��^I֥�q��{0�dԮMf[�2D��*��#�i`@>����q����n�kf�T��}(:}%s̾G+���k}�Ѧtq۹�N�����Y���(�\̣v���Hv�B�\�:jTK_+wz ��=/L�בI���1�n�����,կuM\U{u���g����Tw�i�
^��sk�!l��m=�c��f�;�1/N�?-t��������9G�ڧR�������k���ՙ�2�$�0D�P����#q�&���<��0I/:�.�J�׻���W�m��ui�Щm1��b������B1�{���ܽ�?}���w+�����
��Œ�[L�ޚ�nl��܊c��Y�)&�>}�H/�W�>��j�>8��N��®�tqc��W�S�Q[!z2wĬ1Op�%-�Eu<D�{�������Q�2t�[z�
�h�`�*[GUc�¤8|��*d�aKQ����o�׵n-����=V�.���p�#�]>$�K)��ÙmN���C��CV�<��h�95"�Lj�DBiOq�H���3!i�+h*�K1�Q>v��' �>M�� g�k����b�I^]�呚C�b�7CE"�7�z���vG���ۮ�\ w;��Cr�E�x.,��$��Wk*RyFʩO+������#A���������R���+y�850�m��e�����2R������*oQ��n%�6/�ж��_���<�J5�tw�ĥ\����$ֻ�?j!O^<���8���/o!g��lTD[�M@�j��7Mpq���L-ѓ��m�5�#Y��v����Z�^/<�<���9 ��,���U�Q*Ζ'��V�~G9Z*y����GG&�� �>#�\M���i�B�^.�[��~֖�����GѾ�%f�/�����+T��i�8��(Y�͊�Z�^� ��/i>sx��r��FK}�6H���-G�!ajRPj�ۖ�r6�ɪ�;��Gbr����
���Ym,�,t��QF�VO�^��/)�i���w���M+��|G2��{n����>�f�l���+a���>Hl�+��X Ʀ����ܰ������`l �ڢ5�Xn�w�mDΓ�D94�v�G�&�D��o�:�+
d�
��n��q�������	Þu��]K�;�B1�*�!�P�ẖ��[��0U{�7#�D�s5&��
��F�7��MA��5ZbXv�0u����+����F>f��1���H�ۯ�)j�`�*��m���V�"r��F��nhW� N��g��,$LZ��m�X��-{�o6�Ou�x���s0��Fp��KRe�Q�ݳ��/9�,յ73^��d�Z�S"T���"r,�8�Q��z��L���Cʷ1�ջLF%L��I[g�R����jP�ڵ�Y��A�f��;c	˦���V�7q	%k��OzҭTi�kӤh�N�LلL�l���O�l��@>vK��(]��J��Y�gQx�p�cb�.SF�Q5�k��Dm���<m�G��t�=����5x�3�E��$��!X���S�|7�j���'k������x��Q��(�������ʽL�/��*��[�N��J���wj�*r�l#���f���7�Xg�m�V�Af���W���h�2���}^"K{��v��)� ���d.*��t��c{G"�bT��[c4�`���{���:��u�|z������/|~A�������cb����^*X{�١�ͤ��|�/��͍��7o@/����b�>�|�iٮA�z^A�X��Ko7��Z��њ����=G��	��)�Z��,����鵬�R��8�H^j���kؕ���+�n��-H>w쁠7���������C%�+TQsV/�@�Zb�ͣ��χs.*y���WX��!7D^�@��`�6l���H䆩ѡJ��%��k���� ��q� ���׈^0�ӥ����6V�0q��++�,Ϟ�CS�_��f���g�U�����?l>FZ�M3�L�u�Qʴ�e��E�)U[@������ȷ%��~ɽ9˨}C�|��t�i�Rs��z[z�������^����Y�p���Q`�6}�n�v��_)�_��]��ڮ	������g ���BPai=�z6�5�Z8�� ��B5�,�����r�&�W�'Hͧ�gS9��Q���!i�!mU)"�>��ʳ��<Q�;�j�2=�j<A����f�y̫y2�XR��؅o�-��x�;[��<����,I��6�P�Z�k[�[�j��M��fĭ[Wk2.R�t�3*S���*K۳���UK�A�/�b��f7�tM4�w^\JB�aռn����թk-�x�Κ��ނ�����&�VE��gI[g1&��Ӓ<��B@�o��鶵dF��)<�u![c,��}YR�]�Zv���1�ko�	�ؗQ��Y�Za�ͥ:��P8���J:��M���&�v#�͇����/�e�ɹ�H�3��T�RK�,�x�v�
��>Sb��^Q���I��4��]��lvZ����כZ��kxҩo�6ӧ�TD%�Cip
�'f��0��u�L!):�|#I�	@�6�V�69ݹJt5��E�l�H�b�j��4B�O"Bn[r)���&��)]vۂ-��}%L�����93���)���%2�Iۗw�V��A}�t���\�S����O.�1�g_mJ�K���kX�A���䎔Ij����t���3n�]��ܴ�E����U�W��i�x�%++qm�����A*�N�3*�꘣�$����^�.J|�h�#i�8k��A�e�I*�B���3�#.��3k��y�DnW�;l�b�(v@�0�q�E.[�jjɳ@B�I1���=tH�G\�GZ�-�k�W%���&Y��ohخzq���2�8m��"8@+D�iF�at�<u�@����p.-z��܋%[&;��l`�G>u]�M.�#qI�8
2��Y�Q���*}�78�u�>��h-)����j�D��ϰY��0�AQb��n^��ǅYb��;s�)0��"%�iHM��l�����̠��ź�Κ$e8�=(�8��\�]�/W{elH���#j�4�QU�wۙ��f�!�ͨ�%A��I��7��V��ݹGjwN��
f�|����$M^������,�J�.��ʥ����gQQl��N8����IV�7�]��P�k�g;z�K�V��
w��"��}�}J�u�+�ʭ����+�qeD�.L�k^ⱻF��Һ��OP���&���k'����B�1'�ɏ)���eGznWc�h�$�gB��;�fKC��7��J��dE^���9�2�wQѢ�.:���	�7�t�@F�僀��_N�Z�#Piq�"����np@$���F@��wջ��Z15R\̴�Ʋ�̆;ͤ�-$>(���֎,�U�T޿s��Y�f���ks����7��)X����̭,R�͗�X���7;�Q�w�]�����ֺ�*ۖ��5l1�Ѝ�W�a<�;D�)Vz��Or���+��6��m0��p�����=V��u���N���d�2��tH$�4�v9c��.������J�x���0��]KN��|�}�;p�q�l�k1k��w�ok}�����^�f���1L3C�h����I�R���Il���Ƕ�)���܆�$��)�@H+Ϋ�@�Q��HP�I�FN�L����ҦD�e�BI�4mi$6M�p�i(2�20$I,5%�%Bd��(a�\a	�b)�1�%��
)�Lȃ2�ML�S2tA@��D�ɘ�4�4�2fE��1ACT���$&"$��XB	�<됈��ۅ��0�
H�@m��L^v�DHfRQ��̡Q���(� �D�x�E"b(�Ő3�����,20�1��#5%��"e�&����U.�7OlqQm�� �%s�tYI�q²�w��h����.�����,��YT�ofkVt�9e�N@KɄ��;�>o�d�X�g+����%�Ry)6*��SSC6�Q#Ykd���P�"�
�q9��Mĵ�j�Sx�KV�A$׍�.[[C6�q0}��膋�D�Mν����[ӹ=��?7�=Z�	jR�S%���o:���Ñ�*i���j94�8ą�g�B��ORޭP���'��
�͊�'�����<G����^���]�u��V��9b�B��T%�l�ɧ�l�gFQz��A��')��T���0ނ*��U��j-�m�Y����2�>6�զ)L1,֦a��
U��-�F�*M���w.5<<f��告u>�i[��mz-������e=��7
�ыҍFA���3�w��IȦ��ϻB�������$+�*YE2œ����Mw���m[5KFؓ�f�d/n��6�{2:���s�e�ꝹG쪻�}��"��>�:x�|*�zt�z(��s�%^i�ڗ�i!��ݲq:{u���ЗV��YJnk���YnyVPV���EF���KPIr�\�U��Z{0+
.�9e�@p�0.�+3dͨ�ԟ
�|#2A�J�C�ä�aHmi.T��
3}�DcJ�n��L.9��4�aI�+�
�}݀"�侏��o���gJjIZ�1��9��{�V�ʙ3�'}��j�e!�lʻ��̓�?o>#ցXHb�'�Z�e���J�Q,9�N���C�~�����@��9���cgay����6f����!i��[AT�|bO�Ý���T�wYwL����IC^8k�Ct�Eة��*Z�+4ED��"�l��w����NX&{��Uƍ�&��5�3��&�!)&ŕ)ޖ0�pb�sBB���ӎ&)���Ѝ2�B�9"�=<��3L�_fygk�U�,��Z�����j�ᾧ�D�+�l?Z�-�}���9��((HM��{����C�m�ۦ(�*�m}ђ��o3��t;�K�f�~�N]eﮠG_��w`v�I0��>؃o[�Ub��m����M�X3�ڊ�# ���h,�&����I�T	���A6dƼ��,�&��wm����Yӻ;w�p��\}C�U���3D�rȍ���9`x9��E�Bc�D�܄�E7�(��,����םx�5�E�AS��z����5�w0�>s�Gp����Ŋ����,�῾𧳺�$�FMg4(3�e�0j8��qS%K6��nѸ�rl��k�a�s
��9��;�č�ƫC��EꎗP��:x�Ц��M	)bi��wru�S�.F?t�w�&/[����w�U#��T�l�a�A.鞡�X7f�-�/��v�])����E�##�/N�������55����a��d��1L��JEexJ��`ύ�s,7կ.����eq�.��Ud�x9k�'e��t��;~Z����\��J���Q���m���'/|��Qb�gGn����o�g���ΛDZܴ�Z�dĕ@l;�f�7 �����'>��A��B	��O��+�^W/4�K�$Y�I[k�|apZm��^C=�Cފ�jZZcB`��rw��`���o���E�'��I��B�<�`��1�{R�_\�ɘ�KW�;}慷f�ӛH�N�$�nf(���[�%kla)�O�<���z��T+f�h���5A�UF3����U�c��+����f����1���=\�>d����=��`a�}շ�z��*nҲ�Ee�������g+�	�%;Q���&�P2�: h�G7z��/4�}��7M��D�1b{s�b�b/M������UiC����3ޅؚ�]w	{��L�)�7�"%6�"}ZY�=�6�����ة�y�����lg����+����z2!��d�V>�sZ��L��=^����x��8�g�Ė@8ōV�[oEkK���R4b}�1KgЭ��Ƹ�539\�~�����^���Q��{������YV��Bz�]C��񙏪�ڗ���#]��n��k7�ݚ����*����v�^2+ʌ1�j�զ���fg�I�)��#4H�������a��pH����g�i�<b\5�hQ��fpڒn�1,�2[&eh>%�Щmz���Qe��yƛ�C��UV��P����E�RϬ��B�VN�^1zi�(�D:0����ܚ���U��L�/=�K@JZ�^��`��"�����g��f�*U�j���kY݂��du�*ة��Y}p:U��H��L���^���rt������i���R�p���K��]�F</@Y-�-�z�Z�;<*�b�"� +.�av6��޻�"^	�{��lec��7
i�5-�H*�G����o(�F�i�y�����[C:&Z��d���zԭ2�&.��\���e}.�[��͡��EM���ty櫣;t�`�Ȋ*iPO� *��H����e�HZ�PX��;�m�0ӊ+ε���n�yW
5��D�&l�*��-uL��4��R��B�a��i�2�(+)�6iBՑV�kM�ͨ^�Q��Pٹ"wJu^A6*"�
jh�J$l:�4��]`(�,�g���y�yn�s�S�Z���'K �$ة�������;�%f�ȕJ���ɸ�н�>I�˹hV��YK��ꞯ�>�4�e�2�W8�����w�����\k7��+W���B���D^�X8�e3�EK�u�Y���]O<]�{�V�����z�ꗜ�������:Ci�g9��L6	gF��P�m�Tz��]3j��@�=�uJ���먻��x�h�k8�x�n��M�V�304�wO�nL�C>ީ>����_�#[x�^;�Å���w���o�ړ�x/Hδ(�\���o�l]h���T�2;�+���Xx��h���G�EX�}g9��l���_N��ib -�Q��=�9��V��R���v5�y�0��7W������'�=�u���C�g������ehg��r2Σz��L&ݟ\�׶u
��!J�c����,�!vv�"$՜�ܚ˭���}�p��%�t����Dpw*�9}��u�J�6��)��OR~!�En��y�Ʃ�D��{FH�LT(Sb�e�4�HW�#��u]-SO��`#��GC�����^��� �!-���u�}���d�r���xf{2�_�!L� ���U����:;�s�Qv.ok;jG[�9�ш=��j��MH[�����z!�P�t3ƋU��U�����-��q���q��nTt�����tΖ����/LЦBy�ߕ3ù��������ѝ�G:�C�4��6����bz���QƇ��wSk=7M�4��F3S�����Gy�d^"w����4ˉ������ꇦK����9�z�
lwh�u���_,��9�n�E2������)�.4�,�Nu�zm�L�;����M�G�ٲ�+QD��ʚ��(X�kX'm\
�z��`��;l�m/��2K�^u:y	C~\i#�Et��JJ�l�����w��Wk��ʇ�1��e�kY���-$���֖��Ɍ1�+�=�.h�����T����]��!W)̧�٧���<��f��K,��%���B��%�&�g*+�3�b�8����?T��
􅃤V�"a�^�M�܆�͇�sP��X8�.�5�K���|�oK�fޜ���t�5��������0J����b��\��2;�sR�L�$�kw��L����������og�qqt���}�|�u��C��`�}K�Un��Y:M� � @�f�N�gi�׌��ad��8f�M>�l�ʛ�6���y\�D��ru8���s�M�ক��Jw��:��g�[=�����o�c�|�֌f�'m׵�B���f*:luld��-�e�92D ��['���b�x�*O�S�r��R�S/��2��$�u����͉eK��R�  H�,�Dq�9B�#��b�q�u�3:�<�T���{+�z��`;��r ��hYE�i����< ��s�,�� �ji����QA������MP�٤v���5o������)n�Q|3�c��ÅB�3=�q���P*.�zNb��q�ޘ�]��R�|{n[Ԉ�00f�4є˪�7^��¼��ܨ�����{Z��Y�3�틬<e�6�#���Og����>��Sz�rʜ�Mu��xhIQ�0]����XY�%��Fuy4�RC�%�iOy�,dȞ>���#j��;UGU�fZ'^���IԶ�T&q�,Gy(�q��f��6˙��5C�o�}W}~���������DG�q�m_M�u�r�3���t�����E{��4����GX8�f�W{I��nD���������w�DS�95t��{��;ñ��k����v��mcU!��wv�0Ηst���3!E1QP9�Dه�h0�d�<2�7������*�+h�ܞ�4ޛE�u�����:ۄ㼮��
"�a��d#�%�Y��<���)�,ʫC�*�{~6�b$�~c��0
	 �����w�ޗ����o�)���l���Q�1�b�&�Y��G�����/?z�KdԲ�ު����=��������{���y\�t��<����k���C�La���"]9&{m��K�E5�W��h���*�
��y9��^.�����t8@<�\���Tңe{%?<�'e=�X����M��'��5sS�{Pz�&��կ}o<�[FҜf	W��@�lױf0��k)���g��F�����M�p�X�w�7:��U��Ol۟g\䍴�`k�t�`�YFD`�	���	��ͅs=6�)�)3���O��Fz�}��<F�;nO���/7�phP%���d��_�6B���n��(=���f�C�L^/�0�N�y��6�M-k�X[�U��t�!��-���,Z$<���\�/���ޫxxgpW+�]N��@{���93�ÛV��ϖZ�)�>w�يRqҝp0�y���%; ��,�A[D[����1a�_{A�]�
w!�"�����g9���U�,�qTp��K�p1�-�X)�)��h���0�P�s�<�/X�\��I�y�	��5�aIzi��ڄ99���q\�m�#��r��Q8C+gۘ@uaԋ�zt\�����ͣ��`
�]��x ���\��M9B�.�~N9Y��5��]gUmi�t�r���iZWO�"�}ɍr9���,��]�t$<=f����3��q��"an)M�T�Z��u8�� ���e<���GB�ʃ�u���g.�&��eL� ��݊����5#��2�������}���L�f`'��1���,��h��9�v_�'�Ԙ���x�{-�C�|��+���#�/�3�V�'�t�	zS3�)��to��/�ud�Vu��-�;�h��/�7�F���y��T%t�����᭱t��y���`n���H��������[���T���p�<��tS�級�z���"�����
i�7�ʱ�hР!$�����	�R�0{%�a��!/��0T�5�hIkr3|B��k^�c,���}��zЈoS�`���L���O�˶����S�m�_;붂b:<q9��"
����e)79��e�m��(B�6極|Ú��|�ϼ�Ԧ�:����q�%�\ÓoA�N�`���v��||���OMh�a�~J��̘���v���3�y����K�)�z,D��E0̖U7=��B�0V�#a9�ڹ�CT' v�u�M�u`�0�sgL��Κ|�.��g��`��t�ᑎ��0d��`G��FRň���Mt3�q���4�}h*s��t�>�m귖����{=�6�!=��;�רd�A'/k_�Ă��p�ю��ֶ����Rxw��y�s���Y2A�$��$�
��{�Motʍ�a�^��!x�G�!�l�;����\��б��ߊd5
������5pof���ձ��aDH�<���!r����G��m�e?{z댭��}X!F������m#�yt(Sb��a�8Hl�s�$�V���.��5B���"��aj�10�j#!Ίn�)�㲹��\�$;��]��0�~��H���k�S�e��|�m8H�/�9;c�toFq���gT>WT�
��1�5��!TC��3��{��%M�N���[�1��X�xΜ�V�ǧ#�Tv��u_�u�6/.9����¹+oqI�̈��'e����Frl.:���N�Qt�⠘�;��l���1�sZ}α^��H��M��#�U3hI���-o9!��7bi+�x_��6�b�&���eAe4���uw��xP�.�������G�Et?f��R<��h��U���r��y�xz�m�h�)}�^��`C�Ŏ��]� ������Y,�e�΢�u i�4
��U0]�eK�~'.�^���r�r����,�镨�Hˋ]�}ES���y	pc]��ϖm
�3czO���fa�1��|0f����:��k��#��0]���K��e��mc�y�0���KT!Y�����Ɗ�������{���[���.��͋6��V�:���UV`M"�ΉD.5� ���u����A�dB�%�����"ٵ���%Mg��s��b�_��	���sFNM�mQ��g���:!�<�}1
*�e�>�OE��k��ۛ;Cy7)r�m��t5��,��rβ�gZk�qf���tl��C��6�g��Ws����=F_�?�N��I�"�۲��y�k���AoJ)r��4Ʌ����D�U4K��{yW^�����1Һ��0�n%�[Xj�H������ͪ�Iu��³O.��hoB�fT+��S>���y�f���g��X ٕ��Cjm����bV�cuayP���֡:�[hf0����i`��g��wS˾��������pq��/��bƦ�u_d�u�iUݛՑ��zR\�hL���s����@��3��Z��� %����D�\�(�N�۝��ZŲ�1a��L���=�����t����rO_t�1����6��ĉ���yi��O[��m0����Ut���m؟[\�+0v��x]��/kI�t�R�Yc&�h����/F�p��B6Z@�\)	���v[�y�r�o��9��z��	HLvc�zܩĎ��\�Y�Y�C�pJ����&%�2XbT��&�r*WV,	G��x��3��K[z+)�nr�	Aw9��A<�������W�Y�2�p��bmD����y0�ښ��q�(�����=��4���.�P6��^�<�]�s0O��ͷ�2@��J���O����At�/nP��F$�	M�&ޔvWP���wj�84�r�C���9҆F�s��Uruχh��B�p�@\�j��:�`)��ʻkN��[��!��Bh9�ow7�z7�2��}�ϔ�BL��K��㛨+d�`p�|)�Ww϶Ƒ.pn]����.�"�4��O�f%ݭ���ـ%�Q�ݴIrq�b}νL�Z�c��؜3pi�mE��'�dkv�B���ޝ����U�Z.�u�6	1�.]��n��K�̍��b�uA.����at�NK�l�;���AP����]2�g �;}�ux� ݳJ@�V�v����������מ�f(�jJ����@A�r��0�$"$�	���z�2Tar�D�2E��(5�`�K
l`0��L�64DHI0�ĔD'��0E0�F��
 �"cF��#Tx�$d̊H�,�wt�Q��\�ccHP�Q�e0�(,����y۳F� �Lh�Ɣ4RT�H�E)�1I��&���a�M&1`$�2�
$�$�`FI)�W1��bLb7�撢�b�d(�F������%&�c&-+ьb�0�H
5	�Ϸ�}~_�Hp� ��Дo�H!��
I�Wt�if�1�x�v���o ��͸y��r�Ê��=����Y~�*I�E�!����lҔi�(P���,���fR������;������zfxK�)��xw��W���)�W�<��59�w�Q��L�	�	���C�bz���QƇn�����Y�o�����8���%��W�u��Y1"'~F��{q;�/?O�d:};���I��#���ض���SU�1�tswws+�sC���a�3td��c^|�H��Md��9�)��L��L��\�+�{P�Ix���k]�u��|�o6S<���S��D�kN�`���t���p���)�~�hN<�r�|�$����]��C���uK�oK�fޜ���uo���c�ި�'5tM\�TR�i�9������rjX�1+C[a���[��/��W
}c�8���d>ݬ��o�T�e� ��'��L.��1�e6Bw��Nb�zw�6�O;�O�s�*l~���0v�s��W7D���>M�ক��6Jw���g�[=�����o�`j��;�p#�����mݍ��װ���ݩ�mJ2�n�l�L �*��"�C��ws���<J����t�¢�?;#r6�g.�y'r�'���U����9�ʬI^J$�@�J;MǾ�Y�kݴ��5Y�6�gb��Y�>q��ce��<�,�Z{�#��u���Ͻm*��9W���8���|��[�(5a<�e9;xҘ)�T���.�{���q`�I�H�~����{�S��YR��J��D���T�#��L��f�oi�O-}����0���m��K��l_�Nm�e�Zgd+j�O *�Aw�{2ʽ1�g�{�.���.7�5@ז�[�ޘ�_lMܩ�m�)��-�{�&]���m(;�a��j��1n��q��5LG��
r�R�|{n[Ԉ��-�i�)�uW�m#�l꾖�7���xL���GNk�}�f����� �B)�Ck��n���Q��_I|=�t
nΦ��9mptm����8�`<��ܢ`�e�ҧ�r��]�B���M]/;�h�����kF�Fl4Q�:2�,3�z��@��S���6���L�Ǣ�r�9;f}���k^<2c5�;wM}Yٌ�g��06����'�u���y�)�醨3!w��Y��\�d��I[�1y�<ҟ�k��3Zxl�]�P)��� R�}�fBq�z���~�X�Lp7�اqv�)Js��B2�/n�2{PǍ1o=�pO�j[��7��55���;�3��=R�^ޗ��;�"�T�즚���w���<jǂ���7�ƢP��7*�F͹^���\�Z�J�[���m�[�g��(�U�v��9wo
��k˴o�i�ڹ܎��̅�{}�����R
떵v�d�eڸ��7/v�:]Hr����*�'�=2�wh����$ff@�$��bߥFp�m��>ɚt���m���芾��}�Ӡ�lG�_=	�ƍ�j���MG�� g=CAǌ��M7<EJ�q����rvSט̪����w���y΋�[3��'/x��rY�Y���^�2+��-#vW�Ay��Y0d��l����󐨇�������h���F�}"�u�h8x�>uE��d�`k���`�e�NL�HL�E�7`��m���Zwt��޾�xc�%�Sθ\uK^Z[e�(��RɄ�[ܼF��7�梼��EJs���Mv����~QX%^�,��|K�p1�-�Y��"��h�\�)�+�c�]�j�L�4��F�z�R^�aB��u5<��s����ܩ�l)�D��<�M���u�-;�jGD���� ��8�צ!!S\�ĹCYR�ǶnO��t�Ƽ��rS�;�z����ˡץ�cĎb�S+gܘ�L�9U�Y�d;���4�Z-����;z�+fS�6��mF5O]�c�؂�d>]�0�^�O5�2:+� ;�Ȇ`�Y�B��֎֭��ղ���n��\u�O,ސ�ˉ��QE@-��f\����ż5���묤��Z/dN{k�}��Y�^t���Jõ�h�7��5Ƨβ�.�Q�s`�F��(��;5q�#���ܢ#i�
�5�Zo�kx����x-�r��d�.K�-�f��0����3��-�#4rѳ�;�a�z��M2��	�T�(��-����������}{H�,���p�p�	��/�#�/�3�V�'�Ep�Q�A���rկ�+"���u�8Mt:�z�D�4����nlS�j�51+�p���}�B[Yt��}�Z�N��g��8z�m���G4)����]��N�c��;��%��ߞ�I������#�s�s��LF�<A�z����u�e#��d��q�%�����d7l��
in�{}l���OMh�O�P�	�.q��0��^c�s#4��%��y����zpD��E0̖T�s�!�c=��y���d�\/T���32p.P���y��u[�yu�H�c��0e4t��g��p-�&�x��e���ӑ�d�� `�����[,A�;�A���3ϧ6i�G\�=�ٍp���:�_^�j��4D��gz�`���Ɋl�ke��7�PgJ�:a=�7u��d�:�=&*�!E�+t��\}G���C������<z�1�����
�#��r��Bƞ�~/�^�-l�)�$B��D��C�t(롟��/���^�����ǰL��Ѯq����沺mʽv�K���ϔ@��̾VE��q�r��,��GD
U�l�34��S��l������+,>u����3LW��X���_J���|��P���gvg���6�P殅 *�D�2��#��J�r�&��駓�J�=�A5�F�6���4"��B�s��;$��ђ�]
 T!�;نW"�1�����>�os�Y�#-&zY�+L����`q��[!֊��)�㲹�ٟc *e�ʊhݬ�
~���V�2�٫Y���U�BlsUB}��8-�������Ψ|�uM ��1ㅦB�i۰�?E̢-�.�i��5V���+�h������D��Q�]�;����Ѵ�U\%U�{w�d�x6����j�##��������0zw�ۄ�o$:�z���QƇ��+����Ό�r�F�[v����|����ͯ6G��mѠ��N�/�팺yӽP�t8��m+FC�Y{0���y\�)�ߕ*a���Q��E��y`�de��E�^`����R�P���������jn��I�P;�vS��e���:��K�6�e3���e1Ob�6)�62�4���;l��s;F�x�Ym�c]�S�D�nk����]U��
�~�M}��6��_+z_oE�o�.yվƿF�rp��;Ng+�&/�9t���I���"�)	99�fE.��mŀ�%�M��1�W^j�˩�"���C
��	�
�t�H�滗�̥d�U�q��p�X��j��ʶ�ыv:X�d����V ��eI����h�K�2r���x��2�a��(^�{�nEi�ѝ'v��k��߀cX�%�&��11=��4�Ι���}���[��\[|����$t��h���%��QP8>s>�9����ң �l��k�Nb�zw�oD�ӽ4��^�3�F�j΋��rk4�;3��dc`nߺ%���o�i^?��U��*�8uQ����΄uūrE��[�*6�g��7q���q�9mIJ2���2�NL�;����w3�]�I���nk9=1f���-0��N� �OU�>��O��e�jR�*�a�Ȏ"�!3�:�h��<?�[孺��sHΗ]�.���E%,VŴ�)ʹ,���L�uҞ T�ݬ�)�h�|�F���8#9��r�z>�0�zg%|%��z����"�`p��Tݷ�8u��cXb'���-~�Y��V�$��w����/��#�E�
r�����H� X��i�)�uW�f�L@��mn�'+LPBGxw�B�8���6g(n�M�zR��Q�E�=�'@��ט8��zG"�?P~�#�F�ﻰ�מ
~T���,�wдC;ں^[{���wh�=��ؚ���i�J�����ϊ|@>"�L������N��}�2��[�׶�L�#��LۜW2H0�c"�j�'m���\2�vQ�m��h*�/7�'��c
�/v�l��ʮ�{jT.� r7�|$��:uU�bʹ��=���X:�ϗu��Ⱦ"5�
]Ӯ���@PX�TB�r!�lÂ��g�\6��Nu�����@?4sm�(˺K���8�㭐�w��_���y���\��,%�ǣ���3&`r�]Dtj$�,�#�,����L.�|��n����|zm�E1� Jk�_���>���'MN$n�~��y����Rʙ�z�SYM=�s�=0����;�uE��z�<N�j0n�#O��/�G9�{G�?�/�z�d�����m���芾���7�)�������׷�^9��f]yV�Nȁ��\�g��ʚnx���+�)��6�ʬp=�بX��+���z��x�̈́D>�šO�U^��N���6k��X߈��K:����,}���&&xgBY�=��3l̤�:S�n��q�Ǭ뜑���}�7%���'����a����u���Lqg��9��:]�Px8Q�xw��Z���/IF^ږL ��-�+hB�z��7ѳ��Lb�ޘ�a�z����R�8�8C�]+��O]7�S�.�}�^��/n�j1��� �B�ɎT�#�|�fM�$��+�]3B�JB��8�if>���w֭N����6
�	��Z9�������o�Ѩ�i�v��>F����u��T���@K`U$�1�4�.�|\�	�8������f�m�E�v(ή���T�����3o��8��%�c��j��KK�AO<�7l�Mܩ�z���gf�z��yY1��Lh�*��ݞ�Om�HSLAs��eK���C5�cf!4Ϊ�Y,�>ގ�9�O3wIx��z[�>��� 3�^Ş�w�	
f���E�Cw��瞷�>�M>d�mo�]O�2Q��>]�0�]UI滦GB�ʃȏ����3��Wo1.{&�Ù劋��P澹c^S�H�Q���tl��|��)L��z�9E�s"��F%t�z�a$�Փ����l�<�8$K^<2���Z���[�㼳.��/JfzC�������7��r���VG��9�j��؜�B�-�ԳiڨLJ�-�#���	ll�m�wh}�X���g�;�s�w��s����ĻC6��cߥG`�f�O��6��L�=��w�z�=YB��^F�x�w��)�$�,�⮄	c����W�E~ߌ-��<����4Ο\��k׋�zk4��qՃtÑ�������Ǜ)���A��F0̖U7=������y� ��+�Z�׆�Ǐ���pe�U�1צJ�VRk1����\6u��\����~��P]P�o�y+��XtH(["��M��5ji
�1w��՛d�oBmY,SV,X��D�L� ףM�+8`��������=��e����9G1����R:��=7L��~%K��m�3�ٳ��kˮ�E��w2�.D��uS�s˺/��6T��Me7�tsH�`,��vY#Pw�=9ú#�4�l��(�Ƕ=�6@��V���.ͬ�;�w�|��S#�z�V���K4oV��pU.��|�n�8�&��Me����	���8.�Qo|� �x�d�t~6�����4A�T�[B%��=D��{�+��%��w�'45x��$_�B���/�����"�C�U�\׳���f���V��S�����:Г���OR~"�d�Z�eР^ŞY�T�!!M1�0�e@�'3g�5���1K�͚~f퀌b��e�S�vW?[>�@T�$;���̰��\^��[Q;�;��r3�6�!4ZU�2�G���``5�Ψ|���p��֚�<�7je9����Y�׼_������.0�h��)��ߩJ�CZ����pݝMM�U�_�`,�;e��R��4�H�p�3��1�w�ۄ�o$:�'��{ehp����=�Vˑ#/v�/[#gZp.�l����4���e�����>�O'j���-K�L��tv�;2��;K��G�ݯ}G� +��gs�֥�E�P9���ܑ4譜���Gs_�z�"�yu�x\�rV��9t�S
��[�����<w�#�G+���1��;���y��;�2y"?u4:ȇ>�r�k�?Kf�t�w��f���]]N�ܖ�Λ%�u|�k���!M���J��?�>E����X�C߆'���b�D�te6����-SP/�9�wW;��d"_)��)�Y�M��)�x��b��c,=Rn�-����P悬�nHL���'&��3f�V�����)��]��uK�oK�� ������Q;4�+���;�&�=�y��|�Ln����Șed����<Ӽ3�9�O�_k���o������Va/zp�'t�u>|�~��C^�=Sd'x��d�!]0�bz���O<א�̺N�M�ܽ�x�.z�_���xr�(��^N�:x�[�����ׯ��F�{��j�s�MdW���_0^v��$^:o#��s�1�Ǭ�$](�xC]�e�NL�R�ߍd󻖍�϶]��M�ޝ����jJ	*z����{i=g,�st�@T
"|#e�4��;]�[m��M���S>��1ş,w�!:��w��aJ��(�sp����;!]t���3&�� N��MEtP'��U��'
x�@3܍2�nd4��^u�'�r�(~���؇@p�>k�j\0җ�s�Z�8���gPc�!�*:����};f�F&e]�G�> ��L�sa�!F�ibq��ل=G{�d��6-�Y�z�.�97S�u�e����B�����춽���R�2\�&o�w;�T�a8�ηV��#z��b:���F�sD�v�_�&����p�V(&(3����VڪՏ�q]uN���M�%��=q]�����S����oN�,Fˢ1�$L��ժ�F��+�����Ox;�f����m�s&����Q��Φ.�w,��m���z���p���ʗ�lW"��z��Oe'��혜	v��Vḁ��[R�.��Ř�;�#6�QNf+6�dʶ.^ƈ�̭w�SQ�î��������|��Aw@\�z��;�X��pҔ���:m�=YACc2TU���!�H��Y:9uZ �o6���u+���L��ö���@@�sX���T�#B�F���̚פӗQ��ջ�j=ī��m��I�����Nu�x�3[��&JQ��:�}�sӡb�Ww$d� v����Gm���5l3u�aq��sz�1��-vq���׸Kb�u}�
U;���q��f�0�+��p���}��W"#��e��oPyi�H��]�w
��n=!�+w����;]���Q�E8����!���7{���'1.�G%���*湺��6����	z���Zj�����&�����9{f�Q9�:�ī��^f�,�NRc1�ָX�{�<�{,%Vݰ6�ˢA��m����Z}X���Xz�Bo���U��v'FL�w`�1Ef����%��O�*��� ��"R�X�t-m�=&�[���ʔKI'ndJ��r�ӻ�a	v:��g�gD���h���,|��.wY�n�L�����ݣ#v�G=�\M�k��A�V�������c�����@i� �)oJ(�k�M��u�ٹyl҅1/��̽x���tgs����v>@��`�wK#�ҝ.�]��Y���̏n�e�wm�eu���$P�N�����.(E,�՗܆�)XI!�:*U�V)V���.xᤇ=5R�)�p�Uu��=�a99ҁ��n�]i�jdx�:�/(��r7N���ü��!�+�9�v��/l���;��xW]������p9�}E2�80��U(�-�'�\��Ɔ�8���� �;�Z�M��A�m�=���'K�Q�N�p��T�q��e�}����YcE1��\�q�z[W��V�l�sA�m+y4"�7��[��ONfPl�.a���rjﯹ��$.I/�g�R@މ}tK�}�awcP�9��͋�f����}�4�P�i�=٬����{8�g�߿߼E���،Pb�����I�M�cF(�c�r(�4\�E��&���!��X��k��E�n] 4X�d�b��0��wuE�a�IF�z��XB�đ�<��1�A�E�mM6(75r �4�/M�h�:�Y̒�F���HFH��=y�f6(ܮn](��X�Y ��������#!wN������k���niz����b�(�gu�+&M���,rܳ6
 �)	6�r0XA-�BS�r�p6.U�*$�6 �75��5b.���W��X�m�J�r޻�EzV9\�a,I��Q_P'�4�*]�T�l�m��R��W��ST��y�lb2<dP���Ǟ�X�
�G����/!&���cW�G-,᭥�v��&3�;�Z_|�]�O!.Z���oDpR�`p��Tݶ��}�xBr.���6+���9[�i�އ�]��8��ji�'��S��W=��-�DgvhΥ��4��{�9"LWZ$GAy�d�)�<;���,���S8(m3_M�z�h����/�YS�n'�k�0Π��x� w��4h���i��1@g��ܻ��|DS8c��t���8Ũ5�-"��Ů%e�jD�?2��Gs�{{�u޽�}m5
d(��P9w#v�<���%g�]��g&]��#����|��,˶�
�]%�sſ8�㼲�qL�f�a���F,	}Y��b���/�lV^��&�"�H��	l/�vf10���!8�;��X���Z٢C���Pf�:�7�~P��Xt����,V�iu��z��ު���)��Wts8�c�/�8��j�E*ָ�s�pRx��nD	fF剷��U郃��Fp�	�rf�=x��a�~��w�@�k���i�q���]�M:)u�[�6�ȁ��.Z3�`eM7<E4��M���['e=�@ye��y�h�-�,_X	YQ�
��f�{�wZ�ޥ-�{j�x$�hHq��=d0��G�;>]H��Wti�ރ�n"A�c�SE����j:�����r�c�|���n�V���I��P�!�^im�6=��AoR���\�=��6��;(�&���4"V8;Lb�6;:-��^\�����~�$fK(����3�ZR�l���w]���5�����S�Lΐ�y�����<k�:�$m�;_o�3�(A�]��u��a�wDV��&�N֢G3H�~�^����xbzO�Sθ[4uK^%�^ь���d�lR�Ռ�1�9.����Lt=�<B{���^������b�s�c�>%Ҹ��,���6E6��s\�0���4:��u�2��`�zf8����KK��sͷl�p��_�^x�h�XZm�
sC}Ɏˡ@��8���$+�\�ĹCU.�y�S���}�ϣD�1]�F�؁��9�$�`����lϹ0�,��Ub�K���HT�Z2�n��һܐ�Ŋ�D�f�m'B���e��vt��3uU'����X�P`9K<���)a�x�83�Ti�b��>�˖F�(���pȷ�����S\&�L����r�vOL1�4�e]��j$'u�JZ& ��yg�*�2,N�j#�/�3�W�q�|�o���uC&���V�z��9�Mi�
� |������9u+l.Z�h
YZ��%l��L���|o���.�RL��^	b��*>q�L��Ʋ��K̍��K�\��G��f��.%�R�]*R��j-��Lw�/7_j�odTM�Ѣ��1YF�=)�%F��ǥvδs?�y�;�P�<���^�\3@u�ӵP���8_�#�����j��U�j����m�hm0���nL�b���.ڷ&�%G`�	�3�ߞ�;�Ў�	@��٬s�?��/K�c�.�M8+y�Y�T�z����h7T��
􅃷a=���I��j~�ZhXR�!��JkE�9K����~����y�����A�p�x"�3%�4��О�ݘ��;p�\u��h�j��GX\26ᙕ��OK��y�<�o:�����$Y�w/|�2���z*�:�2{�J�B�#x�<5�� �wƍ���3ϧzi��U�cԢ�@u`ú���Y�N�ɪ�!����.F<p~1��;�Z�a1�Z�=�
��t�=�A9��Hs�I���k�D��2�ڞ�J2Vç+� �z��"�C�k"_�)g|8�[F^�?8N�#3U	��V�K�N�_3J�tm�'je�*H�P�L���S�FzT;���&�K�Uw	Xp���<D�l��m=I��hY%ն���.� +���*9μ�����6b��V/�/��'�TBc{�2�m%�6��LCIQ4���F�kj�]4_yma"N��1�罦�>���oFQX���������!2�9�GL���X����Cm-}e��*ʖ�!���Ϛ\.S��O+p�d��`�"hd,(�E�:j]�UdU�n^��'��Ni�oU�y��F1lX,2�m������2�Y!ܨ��]�"��c�f�꫰��+��E`�$&F��J��pZvuC�LJ|��h���E�5�Nݞ�)a�n}��<�%�\����[}�JU��6�F7t����pH��N�lV�^���^�1�0K��:dh���S<;�u��T�	�p���R��/l�8��w��kO0X�h��A��6��M�i�1="�̇E�����p��$��?Nl�O���f]�29_cS\M����6Pm�9�z�
lw�.��
*zF3���<|g$SzB��/z��>����չ��1�F�߼��@���#�S�\C�׹g���S��-��?k��-�9W^��ۨ�q��#H��	ɩn�f�V�¥ߠ_t;��n���{�ޜ����O�K`z�X�yY�����'����ʘ�9�5,��p�N�Έ�?}R��q��E�0�
��^`��bz�'ZTWt��Z?]5��O�Iۭ^g�u�|߷(�~s��x��QV���,+%���AÌN�'�������Qղ~�\	�)9v�@"��9�[��v��M�;�n���M0�ez&,J>]�@���G�`�LD%�O�;���n�M��W��PCqX�ŷ�f�pܾ�o6��u>������
I+�����_��O�n_�������nW�4���,m�ײS�Z�p�':�KG[M�?k`�9"6�8�9�ˢߴ��r��jH�.���t�ʽ���7�S���J z��?k)�N1���ײ�������z����Jr͜���ҕ !M�q��5��kn���/kZo	�F�=��;"�lR��IK��}-(�yi����< ���j���zY�ӛG��k�ݫ!� ;ޙRP�-[�o^[����k�Sv߂����ș~�U"�.'wOCĎ��
�x{��\$��b	�P�*�R�|{�H�n00̽y-M���p[s�.+oK�⪈e~ђ�X��U.��`w�a�xEy�Co��>�F�������m���C����\���:�4tʖ�])d~T��^<K��Z#1��иޭ�Q��&����KI������?��ɸF�]�:�]7��M
d(<& @r!�v�8�r9�=�s��`�ˣگ�3�xK5��)�;]�.�㭸N?8��n����@[��MF�����Fk�\)ԗX�-��໲D0�� ��uΜ��ȿ�a�4���-�,� �*��:�
9R��o�%y�'�f�*�Sn�� z7�E�3^��_u-����l��Ӳ
���+�����ܪ�ڍM9�f�Қ���][ӋaNx�͙�5�람��y�5���fs�)fӵP)���@�.�w޴'�ͽ/a�sv�������Ň��(�l;F�ԃcy�b�`��Ƕ��ǚf�X%�jYVoU@jk)��S7ts8�E�'Ug�������î9<��|���@��[���u��0pc�J���[y��j���Ơh���jf�_6�ļ�s�LV��f]M:)�^U��@�{���<fT�s�W�F8��O�Pف�g��Zגϻ�QS�d��.����d�8�2�G�xC�l΋}�]yr�g�`n����{J%��-v���^\��]��	1Ѡf��w�_l��3:��O�/��<k��rF�S�5��g0#"� K�^��żb����!����9��)w'��}�<녴uK^Z[e�)����q��np��wV�WA��,��jb	��P��`��K<U!��t�'���cVk�2�6��5��L�N�#�G2�:$�jJa¦Ne���������\9;�MNq<�^�̊���u��1�:����ӄ2m��5t(�vz!>�BB�1�]M9@��6t=]��O�s�㄂�X�����r"�W)Bvv��ٓM���@cg�f���ͱm��p�rs�L�[�4@�<=�����M�ڔ�<���w,���4r���pm���}�ʹ����1f���]����!JRy|�|�"�,�mc��L��9�I����x�6۶G�vIx��z[��L!K 3�L!�;��z�����ڇ������{Vz��'�!�!ec�F�H|"���+��<�.������Ez��˴���]G��UU�?9������.[���-�Df�C:6q�wL>o���M4)���t�Ԛ���؞�;��;��fu��-{c�o�㈖kǆRN�l�#�/�3�\�n�L�6�N��g#��%�D)
d:6�/��Ѽ%�Ҡ�����iڨD��°�;ܴܟW;�d��&�nAT�ŞW`�Ɵr���%\�h3!��<K�jܬ���������~)�
F7BV ?���kx�'����sLˣ��������,���B�~,2Cqi���c�e���]�m�(��湩��+��[6���/ё��/�y�����A��C��(܌g��<��_]���5�pt��0S`�'�;)�Du�z�����V�Lˮ�E��w3O�S��ؑ
z���i����<�
{g��U��;�oOp��}8��oɣ7p�U��5
�N9�!��l��u��Jso���щO��8���3׏�rS{����r��Q�*RC�i&p�Uug�
��~�7U��\D��iv8����� c̺�st���_�H��ssM�9$5�v�Ȇ*'�'(�}S���P��H���ѵ��tj��t5s����Ǧ��+����ը3��p�h�l!���Wr�&x�"�\^�Q����jH�.Dt��8#�&�H�P�ȗ�Y��m��=:�u]����co�:vy(X��o��NԹeI�J���D�2��b8�Aܭ՚�/p
��ݺGkˮ�l��g	\&۶S��O�[B�.�FHApP,�!�<0�,�(�ocUe���w���1I1��B~�Z��hş-��E2�)������S,��Tړ��Ug���st�ac�>l��=�p�j�.��R���(����Ψ|�uM �%l���z�>�pc��^9����G� ���,��z+�
ؾ��U��3k�ww�m�lM�hGE��8Vț-�D���fCΗ@~렀���(?�-�o����t[F|i��c�n��h���c��3@]��B~y���y�������Hu#ۉ��П����.m걡_4q�w@���Vf������)��Yu���e7]"�đ����ڡ�X�&�[�{�<��\=R�X�#�5<&c�#������2�X���lA`�.���u�� ����jd�H��f�;�n�߲ə����H�Pp"܇�����X#��=E���x�!��f7)_QN�h�י�Ӄ�ئ�C��(�l�G��R>�r��E�d�HL�d���Qό�L�*9���}hD�q{�|c�}0�bSWC���a�coo �:h�sޕ+zA�dS`��5,��z�E�R��/��ouK�6��
���x���]É��7 F�e8�����>SL,`<'&��11=��4��x���3e����Lj�a�p�N�߫�y������d>��c�����zT`M��᯶�=x̬���cbe5�|�qV/Ď*$�8��n^��*l[.����V<a	��`�Q�B��B_��˕%F��8{�o�X�{�����oE�t[���<g��ԑlԣ -��l�B���"p�r�i�|v��\`Y�D�s���ws����J��.T�����d�M���͵)P�D�d+J�sU#����$e�o4�DSH�~B�#��)w�SE2R�l_�Nm�e�-3��EK^�U<wr�I�v�������},�b8�T�IB�A
��z��oLpR;@ᇹSv�ˆ�p6!��v�fP��J^P��hP�o4�x���[M"z.�9Tʕ���rޤC�Đ����U�����Ŧ\��g�l�j˄�o�rW��zv���i ɻzU�d� ���R�\�<��vw�����e �F��^	rW+��:zv�]�+`�f�.��.L�mg':��P}Vq!��l�^_�B��6��.�LN��me��ƚ1t��$pX�ܢ ��8X�l^pPھ�t���MS����[U�[ƤWS�T_sˤ���ѣ�T��tLp�,��ʙ�ܼ����&Ah���T��;��]A��Ǹ�{Q��;8F�^���zf龶���L�Ǣ�r��M�?svA���ma8w���E��~xmBZ�ᔱ;]�.�㯄��'强�SB����L!�+ޫ��S�{zj�0���e<�D\���O��N���LL.�|��n�x�t�t-�{�lGn+���u#�MLm�)��o��K6B�95,��z�YMnӣ�;1�1\eVd�l�{֪_))|��@��r�m�g_��<!�3v�d�:t�����3���l?i�.&��L9�����M:U�>�@�e�\�g��ʦ爄1���Ƶ�b}���n��arJ�|�_���=tɬqd�=��/�c8S殼�{�Ӱ7_����d�z�_T潞���ܝm�N��#�G`��ޖG933�=����s�5�Y�9#m)��>f~v���Y�ɏvX�1Ж^iͅ�%rk�����+s��\a�,��뻩Vp�r%���H��gfVx\q��x������-X8b�_�Z�8�QR�ocz��lC�B�gS�w+{2��z9����t�1��5�-u�2K�OQc'Z��r�r�u�e��_ӱ�k������e5_N6�q�z�.�9����]�6�>#t��P�Qr�r�=�:���i��П��kk7�C�Z&eMV;�,Q�i��j�ͬ௎c������<3�	{!A؍!��9V&�F��Qj�[�v�]��t��3���;�����Gd�9�'k�tCX�K�SS-�G���gL����m�T��嗜�;��9����'�*;�SޙD��9������|�hުkU������x-����b�_H�$s|n�Z5���rq�͡mk��.���mH��ʡ�k]Z�;[œ�xb�Nk�&JQ���q)	�^n���`b�Ő�x�;M�Cr�k���۠�Ê�C�r�k��� �\v��J9�e�(v�
�+ Y���İ:0�[C���7���H��i]�zk���t�iv��!�+�q���3rk�h�S ��75������:�M
��O�ꢺ�G�i�nS� 6�P��<xzbߣ��`�����U�G�s�����,���z��F�ve╀u�:�إB�BZFX�u,+4�+�0�J�΀�q,��p�X�y>}�
)S����ӨU6z�i�n-Ov���p�U��CP��[��P>�ou�đ��[Ԫ�d0ݫ�颚WcX�Ǣ��\5lD�-��N�E!/om^�7S�|�C-����|����J���bm�A���p�v���I�:Ӭ��WQ�K����q�
���0I�<�AmZ.e��M����e��S+�f]J����6"��}��gt�6)6."����vs��B�a�GCN�d`�N��a�8>ڬ$�����n�"�R�v[Y����+�4�2���Bb�3;���Đ7����]8M��򹻌�-:V�����0ɗsB��n�B�Z�/Lֆ:��ҢgKP�9Һd�H���d�ݛ���eC���Bf3� �.�0���*6h:f�ΞB�[9�+��ȫF�:m� �]������ۡ��]cD�T����;�P6�G+�䍫�6�� Rgbњ0�z*X�H�|D�e��;�N�
jYN�g}Ҟ��8�|��_P[3O]�[h\��VD㷍�hn��(�[�YU�^��!��
�/v��Fyn^�+��
y+���Y���r=̚MmN��Ǫ�xq��j��!�/�3��]�q�Nu]jf�*U�I����*��v�ވr�[}; ��=nea�IS�;�tզ~���E}ν�8�>�o%�|��[+��ݵ�<!+{G_muwA��$΄Ǚ�_v\V�Dt�#��Os�/��R��ۜ�͵�gZ̚�.����1�q�
2㼝Ӛfn1D���#b��5;���\�X��4c�9k�n��7��o;���M��)��5�s]5�I�-���U�ڙ\�wnmwQn��$s�*�,��c[���N�E\�sZ6�\�B\�$�F�湨Ӻ�W@��Y/]׃��-͝û[�	���͹�s����.�sh�`ԗ7o:�r"�k��%�r��W-ʇq��[����J�<�n�rK&��vX��平�b���Ź\�7/w&���wr��r�q�\ۥq5�s���$���+���\��b�(��w+��������Uq9o49���&�����gRF1Փ�e���:��EΦj�cV1�Q�8b��p4��wS{;pԃ)��	1gK����!Ku4��~g�5�&s8��	�<�Ч�p���k�d����z����n%7$sMEtȷ�V��mor���1a�ҡъl��)g�U!��\7���*Y���Ι%�o��U�9����x[W)�
�S�pB{i�%�f8��`�s�Ν�����c�i��8Z�ۚ4��I<���9��7m�8C+}Ʉ)�B�9�w�qd'��HSzb�xŵ�R��"b�M�{�ǂ]$t��S�6����m�l�M�%�yuu7[�L!Mj��Y��w�{�#�w�33r3��P�4��U��}1��n3.��Evt��3uU'�e�1�L��P7�`�5�hEtg��7��99���W�s�yrʙ��-�Fh�3�gwt���Mp��]ƃ��l���4��_vb0�0��e�b
���"��,'k��Q@�m��t�{h˧�m�79{��5)�C�7�^���̞H��>	��S�bߗiwZ���؈�.ѦOM���z.���V糸�;�#Y����ƕ���Tt�b��LR�鷣��.�xj�@+R�w�[�fkJ�:�i�~������k)����+j7�w6Y��x=͕]�LLѠ���}�O���	G3e�1qb�"Y46vܠ�3��d����v�|]�_p���I�����u�kE7	���x�o Vr�B�4��+����M�
qH�N�ӂ�w���=��:�~|�T=z�K�E{�9�z�
i�[͒�>c�B����oA�62�β��j�k����/Y5���K����{~l�����֋f���"�}4����y�Zq��8"3p�x#k4�J^v��Mv-�G��]�+H�6BrvS���OK��m�3��:���u�H�y
����u�efk�i�T����!	a��jng.�z�g��2ʠ����zs��L��4r��M]L��
��Gm�z�rD��}9��z�|��b�c�J���;��alѽZ�:��n��1�`)ث�ڛ�K�-���:��˨�j�[RD�p,:q�A�b�9�e%ӹ��N�j�C�)���`s;�e����zR�Y=6�o�'e��H4�@
����S�LGJ�&K��G>��}߷��7�}ϛ&?������%p��Oڧ�?p�K�m!�@�C{���˥��f�j2�ެ�m���xkTAuL�U�-��e���Eya��m����nTYp+n7/)l*�sx;��h	�籠��+� ��dZʕ�F�Dq�����:vu�ta���C�f?�n'�N�+@��$�ۭ�D��8i�7SMױ���o�v��.������+I�E3�Np �#2�M��w��[i��L�y�G�W\ة�����쮎M^jꞇ[��Ʉ�h�hT�k�ɹ��Osp�).�MUn�+��ϱ�SZhr:���3:�g�8���N
د5�[�)THkQ�]�❌8�P�V4�Q���o*h��B^�L�8w���O�,��xK:s��M�+��,�'�C��g[D�aF�u=9d!���+�����o����'�W�sd{�� ��"=���ճ����W�-{kc{��׾����UC��@��#���
lw]]LT�f&�5���oPr��[���dt��M6K�7<��L�
���Gt�N!��Y���LF^�k�(SF��=�9�hrpLpQO�;9��
E6�"a���V�*�f��w�0��(�_*�C�]�uf:ո+���)� �n���k����� �nx��U�b{C_��N��q���"%���V�J��ċ���W{�_{���⢓}2g��Ꙧ/�`�	�/��>��m)j�_,L	QVǬ�7�9�TP��w��_S���=�<Ͽa���x�z��+|�ʜU�������Jt����G�=����eoGp���><g�9mIJ2������*r�ޑ7�2��{��ǿ���Yo�;^=p\����W�k�u��1��W�B
M�y6�\;U�޽i�V��L]�c7[N�S|3?���C��g�a�:��@N)ti���rv��$���;aW�[��v�������J��'���i��!���t�ߎ��ߕd�w8�ܕ�J�C�t������|�s.K5)P"�!�V�+r�P��NԔLt`�
Z�Dq��xo�#��)w8��d��؄a>�YE�s\&��L��k�'���ȩ�O .�Dv���1�W�zJBKzi�oLpR/ݰ8l���F˴"�l�6�aF����0S�+}�x��8E�v�\W�rP��'�څ9Tʕ���ń�9�3�#���fp��_97a���]U���d���ܧ��,��`��r��[��L]�jڳ�p?^�XH/��t�=�gQ}��gSF�n�T�^])�C��xw/�d��p����QW�QJ����=�G3�ޫ���y/j2w�s�{{�uߢ��sЦB��`r�oS<A��X�f�&��b�.6��/2�bv�2]%�_�N?8����y�q\:{�Z51�"�Ct)�T[0��a<�c�����GN�@�ap)�t��K�a�Z�TU���8�C�1R�X�ۙ�50�J�.���pe�^�����
�5^u���("/�����A�E��6�4��%Q��Nq��S'�y[��%y�������(��1s�S:'��,R��\��z�rB����)W����_�}��ņ��2�Io��%��CV]����cC�e��ˢ�
(��5D��o%�S�␃�]�.&⬧�u٪�%j�[�YG�m�%��7�q���z_���ȁ,ܮ[��οT���Lң8n��y���Ge`#&%��{Ec�ՖC���x�[ml��_�*�+�m�u4�=yV����4i��`eSs�[_�tnԷe��꽫i�7�b;\o{�)��vKљU�-��=��-���WUԽ�����)�(�d%��5�^���so3J�Bx��N�}�Ϟ33�80�8��q�Ǭ뜑�����Zv���9�&��J"�s�eM93��#���l	��b�x�='���醫��	��)��0֥��s�{_k���	���a[�<Az���:1��<6)g����8���b��Յ�9�1[��oļG�*鑱ӄS.��x]r�p�E9�Bz�2^�c��oP�'Ft<tjA�#r��v���~b�h)מ��{��a`�eo�0�2�P8.��B}oLBBZ��cm:N�s���F�,.9>�z��J����Cv�ὐ^,o�WSu��L!V���pŝ�Q�́~]��'bn���κ�w�Ȧ��~�2ᓷ�E�#
��Svt��y����yt�tv�[1�џ�n9~��*��0�_r����e�D�b�7�!S1�D�a��2[Q<&��q��2Q�kzT�K����*��w3kC3i8C��Oݳ�x�B�'�6�����W6�x\�|���;��-Q�:�r0���,Wq�:��Ai�Ļ��������c�v#�F8.�^T2��$ /G �6q�7wT>ۤ�D��UmNE�#Ѣz:ds�� �Yl4TA[�~q�O�K1;\E�� p��7˸g�C\��( +x�~�B^�L�H��2g�}�:��/���Kf�u�a�&�c:Q\Zv����H�����C��Ͻl�KcK.���,ǮzEA���%�5nV<!�&�u���ԉ���i��7��Sە�0��T�DWts���ӂ���,�D��~,6Cr���M��Y[��can�;��y�i���&������m���E_M?F�p���rқzpDx��ٚ��֫T36�tu��^4p&YT��
f��
��Y�vSљ��~bz]�Ι�~Ϋ}��Yݸ�ػX7��ҙ�w2��A21�4��
fs�`�L�|e�zN��~�Ӝ+��pe{y�8;�f]�Em�/{���Ǫ�К���=�6�
]�Y� ��p1�T?�N�ֶ���ƚ��	����:(��r����!mSϛ��Gg,� �(�	[�|�G=zn$���Ksp�W���{3��&&�1�������j�f
ޥ�n�ۨҠ$���lj�'\�v�ݧk�:�������U�^���ս��ﻁ9�|�uNBj�z�{uwZw �4�JΛ�w�q��.�ת�(gu���Tr���T1SP�cNIX�L!��s��ג����*�/ҧ�Bƞ�~6�p��.YRD���A��)�6�6�%���i�����29�!�udç5�SNq\'����z��$�׸k.� -��NG<c�&��[ʱ#��63��k��½1���ꖪ����[����h�~�5�/�b���y�����m��\ͻ!ߔT��e� ��B�l�P]W�*8�h\``*G@c%��Q8ӗ�u[ZXb��U5��3�Ǆ-0r�Y�d����h�pV�5�[�$��j�X�sl�L1�7��u�Ũs#@�vu4oL��>=߂�� 9�(5<����K�.����I���t��hp���)���Y��7��^�������^ه{�%��S�/rl���v�̠�f�t��z��.�_�}����+���2���^3��=��Cκٰ%�o:��3����(�ȩ�Md��9�)鴙�eO8�f�w���D�W���3�m�TQ�w.{+o5�l���1�
)���g0T���)�,�5,�ٽU��w���.�^z+k��r�n��ǅ��0A�����c�4+ؼ�J��jL΃����ʼ�fxQ�M+.�%ŝx��u[�^�W�L]��md�	\(�M\:Kz�T���*5G�kW�pg٦��
f.&/&�og�XR��ɼ�!s�ub�����t�3;�ӆ�{�+r�[Me���^>O?y�K�n3�A��_�c_�L��4��0W�욖TLOhmY>�Z�Y���5n��/0ݤs%2^��T��7}7���TV�2[:ɋ�k��0���O��ߙ?�~�5NL�:�y��̜��Q�~މ�7�ܽg^Tص�Hݟ~*�_Y��J�z��?z���e���'`-p{'��F�{���l��Ύ�N�c���Y2A�m�KfY�!�V�b�{��_1���zɦl���;�����<�,i��������.e$��V�ㆴN�յ|`
�8�cm"	�9B�#��|8���R�l[J2���x������:ׇ6&:u��ld��)�Q�̲���a�ޙ�(K��ޫz�ޘ���������4n��7Y!b{��-�Ӝ:��1��!�>]��p\O�rP�1�_�S��\�6"dب4�2358̳Ө̎�O̷z����{��F.���[FH�ùN5ܸX��`�����86VHv+v��*�CZ4_��gM��1�4]�/���t
nΦ��T����$p�kP��������OOh7�_��M�+��)gP��*�1�ݙ��d�aZ�,��.O�
L�C��v]�YG�7��)�`u����r�0��J(�y�T$��gU�nM�m����-T�[�6o#<�_�L�j���gt��,�w��#C7V�1�*�)m��ӳoMM�x#�p�%��:y��/j2w�s�{����o���L��yv�kf�S�Ȫ��'s����p[0�У��.�����	t�N?8��n��)�+�t����qi���㣦�!��L�b�����<��.F`X'����&H�&�we�?9x+0��7c��s��n@u�1�>�����v������ߕ��B�-�R��/lz9ք�f�Qر��F��.�gG�_+z_��@�|�[���u��ziQ�6���&6p�F67T�H�k�DK��]'m�K�E5�W�n�i�Lz��{d>Sp�h,/+��HM(n٬�8sx����=�+�:��6�U�-��=��-���i�^\�����yݎ�S\V��^��\s>f��Ss8)��N��33�=�O�/��<k��8��eR�t�����~�	��{�Vj���Q(`�:���`)<��*�̹�D/F)�Ωz	q\�Eek��; ��h2�)��4�q����<6)g�Z%�4Ό�Ϊ|$-!�1�ᐄ�7n[@�oqc���;������Ѥ�ح��J�l╤ek�j4Q�Ǖ&���f�9vL9�Ee�[��Z9��o��Z�����I�zQ*ި>���$V3�s]I��e��fQ�ty�;0�8ol��y*s ��Zc��ޔ��O]7Qdk2�Z'����Ä�\ۈ!=4�����O�.�1��M�ҪNi^W{6�����y-�#��r��8C&ۈCWB�:�Aw�qd'���쉖[����ͭ��T�҇LF:�j�uR�ǾO��7l���Ʈ���gܘB�vr�Կ?��'�	�����]�BB�#�h�p��׶c(��.��E7gL>SuU'�E�\륹�]�f��j:"c�@w�܇�|g�\"��Z)���x�Q!z9��<�f���z�U��~U5�A�>x���E���l�O�
��q�K^<2�v�����*]���J�y��l�l�3@��8�>]7�^�����谇�u�^�TY��f�3���Ѽ�������n]�C��Ds>��!-�>]/a�O\����m�%�>����Exa��@� �ѼT_���yH��:m��I�������9�8�ӂ���,�Ǯ�	o���Y�P�w�� M��0d鴨1�RpSH8�l���MJzbzkF���.�#��%��6SV������ɡB*Z��RN����z�ϸ&�N�q���N5t�0���X���X
[��@�W�EGU3�&Ñ�)�]ᣥ���1��7�5�F�b+,p.f�d���=�O#tj$�����|�ȁ���:�s��c��/�n�﷊*Q���e���V�Ǹ�:�y&���}}ӡS�(�Vs���ۇ���M���*J7x��,ga�e�T���.Z�9�w�1�!s�j��Q�D�-j���mcՐ���^�Ym��F�0�WuhM<�f� ����Y�8Э3cz�rN�3M�dy2�(5>|7�y�A)A���w�k����6cҰ�m\.��G��U�}��O�R&*���3�+���:C�C\��:X�S������knK��n�F�S��B�&��cl�1tF�XV\��TgK�2�fj��i0OeuQW��sv�Z��hT_p�1Y��gu̙|�lT��
����z�rf]��mQg.�wJ��)e5Qk'jd��;������-�2�u�s��JA��[��Ft�S�aiJ�A�3��BHhqIG-��q攅�R�Qe;��Զ��1�E��<��J+�{��$��P�N����H�TR�}�U�Q�֧$�_E8����]�`��I��E�|��+P��M:(>9�9��j�m�[n��-<w���h��zէ��*݁�0l뎭�+�!#��m�8�[`E��"rc֍w�rU���/��������o-����γ�vw��*��*e��=q킸��.�K�%Vz��YN�X���/\q��b���	�����}�lp!�n��~ywD�}an��!��B\}�Pc��].�Ūr4�i!��njua��18Xl���b�1��0h��b{N����eX����s�Ō�dh�6��F�we�ٽ1��>;d<�5�,R%�Hae�4��k[�#˱�*;�ذDb������K���NB�jݙ{:�C6��~��q2��҂�Nd�w�+�d�q�8�;�RX�=���h�Pm=����֫��t`�In5\����;�J:\ܷH��*�k�!�A�x+N��۳���1��&Y)���ŋ<��@�o��hPv���fZ�Q�[
C&WL��s��%�w:grƪK��t���#uۇ���3QxAH�Ҫ���}[4N��N�Zf�ge��z�;pY�Ʃ^����ǃ9t��n����N�ǃ,TM^[�m��D��N���)�̥�wq��̘ ]ݝ���_:(�nWw"u�}��j�l���H�g]����n8�cd���wAT��K���h�pD��P�]��ȁb��BŐA�7�!M��ܻ��A�aTj�����=^�x�.���UP�ك��7���t���r8��2����Mɚ9��nU�W�U����!Ë2J����\G����֤���"P����>6kV�z�c�b}{�׀��+�z7����_���\��u�;���\3��:.\�%�¸b��Ҽn���pwV��ȱs��]�nwv�+�N�]�$R]�W+�+sd�s�s�ss�k��I[��+s���������Ѷ�ܮr�ۻ�v
�Z#�"�����c�����5��C�m�F���"��7����Qw�m�y�\�nnc;����wmzx�^�5�;\�h��#\7.b��[�,\ۆ������:���6�ʹ�E���h"�����E\�Z674n��ܸ���x�Bn�N��u�C�x;���f�H(-�w�(�uH)wx2���m��7s��5�X^M��d��:A]r�50;7�D�}ա �9�s��d���S�|V҇n��&�� �^�xKd짦c3=�؞�s�:#�7�W�3ّ�F�^����u��U�H�be�`�����Qq1�A�0W�g�_l��A���֪Pb3n�M��ث�E�;0qS%�緪��MLc��j��������3�ߐ��G��?y���r�_9DOm(J�`,�!��9R�mSϛ����jH�Q���|�gG<X�������X*o`^vc9�_dK�Φw����B�]4����52�$_�B�j"�KRM�++��&�N�$���������t��a˚Κyc�J�6ݲ����'�.Iul�2B� ����+������xC&xa},�D1�j�.��U[�-��b��Xe>�-~#M�����9|����3�d���Ezwk0�А��. �R�l$�x",��+X^O_�Z�ۭF���ʡ򺦐W��ǎ�9�;�gY,��OCE3��)��ߍ���v썘q�(���j]����]@���h�n���ЦBǞ�S<;�g<����f��~�~nI���'�	'��l}�w���\��=�0Э�S~��*K� ��ts�.�#Pwo���Ŋ=��i�7��i�Z��9]Qk�̣��w"�U�I��iT�ꇹ�׺���yV�c��[$� ������u���.��\��H��~V�"�=�\���C��Dg]�M���7����@u���\ٮ�nK�\�g�)d�ѻX��~h����l��}�z��� rn����)��Yu���7] ���LI�U'��U���8Lk���+�
4�,�O��S֓5ʎq����u��˭�/��*�e��l�P������c�.~�FƑ�?�y��+�~%��T����[��k��j�c*�q/4����K�P�'TX���u~}�~���ʘX
�xNMK)�5j��R�*"�ܗ"�9iX��M:��t�<o��}��o��������!�|��b���Q�d���*-5����\�6�߽\i�� �0�����4�z���U���]w�0�g�!:����(��݃��d�����$B�w�S�5��>��V�mV�[wE�i�<g�9mI�Q���̰v����tUdɌ�X&��
[��&H��u�y��(w�%I�*yX��o��Ƕ���Y��m	�-܎a���{�� tp���E4��P���4إ��B�Պ6s�xN�ˎ��K��\4��!Kά�FY����"�@i%��/`��0*�b�CT`l/x� ��˻W	c��_���&�u�7]���ZGmU��t�@� � ��=�4���Rk�w�3����cn:�26$v��*���z[}��2s���GoQ��o���m�v�쎿WJxS4Aw�=�e �3�P�P�yoU��v0.m�+��SSg4aa*,)�6��Sv�����1��!�, �����4 OFu��+��GTv���'	O9ƶ���woR#x=�-�i�L�n:2G��>]��|�r�jGql�����Z6ǡ�U��O^e(�{Q�E��7 -�Φ��J�i��G
�����"�L�U���XzK�~�.�ᑨE3�9W!��oq���'xvp�|���]���Xk�w�ۊ\s�A�l'X曅1��@(XC��zh0�d�e­�#�v�y.�㯄��R�Jzǳ(4�=�SLMf�˩,;�u�*وj�28��	}�:��i�#$V�[:�yokdƻvK���0�!U���^z��m�n˾��8�;���S�c5+�쯄V�t/~X�W�����<��5��y�|��r�|�$��޾M=�s8�=R�[��差D	�+����f{�g�xC�M�=��R/�9�rf�=x�[ml�z_�*�+�m�u4�=W4����4oQ�t�"��^��L�f!{��zkx���#�b�g�����"�+��T�{ss���s{��񡫗�^j�5ތLJ�)^�P����$ή& ��d�Z��	�j�t5�Z�\������`�V�/�{+$|�s CK:�]�sj9�Cy"�ݓ���2�L�F8���眝���eV8�g�E�D�A�f΋}�2�˗�R4���lΩ��vњ�S�g��3%�4��
��Y)����<��3:��A�����{AX�^�O	�h��vֽ��;Qr1S�%������5��cj��_�Ǫ��rz�כF�Y]�4����nr�$^:_ttuK^.�.{T��K&W
q��^�0�ҡьx�kq�ZKT":a���0��g�3C�`���Yk��ˡh���0�W�S�q'��2_q�p��񉰲s�C�y�K�;���!үgSS�AW<�l�]ʛ��)�[>���Р��=XܥE��q��7�wMq���1�4�s����(R�Տ|�9���k�K����|��=ql^���D��vGQӻ��k��2g��]�(T�Z.�ɓ��E�#@{ЭD=�����=x&�)��՜����y��1^��~��E�Y,���S��E�C-�E����v�{Ҡ�C�a���Z��.;9T>�ġ!D �zb8�3 �Yl4 V�<�q�K5��{ց���~�k���뜎��mK��+@������k�����dNy�s�u7�)q
�`���S��ɷ�\�7fc��ecG��-c�f���R���wT������8-�
�6�%�|�¸p,�Kʠ0��ff��i\1�@��l/-Ό�����W����rE���̢5�ۢ3�V�'�˦�Kҙ��@tu�_Y�/�*	l�[��M��e�am� =��0u)wDs>�xkl]/a�O\�f�2��K��j��|x`�a��]�|���7��L,M��%�M�>�3����"��9�y<�X�6�d����z�Cc>W5�
���5=�I��˧g0T��m��|yl����zkF��	����c�C�:�.�U�Q�c\_w�
a�{���<���n�������짯���z]�q�����q�.��j��E�j/;��M>Sr+�K�����h�`�#� ��������oa�O^l�{�'Y��/Q��3F��-~o�?;���Z2��j��cW#�c�J��U���jkq���m�Դ鎇yY,9�;�Hg���p������wQ�՜���B�$���4s��6����^�Z{I�ペn����w�8�[D(��SOM�Q8C.W2D�`��w����tჄ�4`qqO��W�T;�Y0��gM<�BW	����]h慒]1T�c�O���h��Vwc=�j3l�6L7{�������%v���gG�K��axK\e[��,���K�}~�A}v��f�\�`
�U�b�+�����9Z�bݖ�Q�j
uлI��7N9�p9����WENWj*HԨ6dgz��̱�wM⏋7�ȟ~*��9Ε3H���P���U�-��e���u��%qr��nqk[�t6u0�׮�,�����@w*�V���HS4�!p����R�������{h��ż�1F���y3vuC�uM ��F8�V��M�a�d�ϙƞ��pV��WCGsٺɓ�*��#�K�1����ћ]�;����ѵ�U�^�
d yÿ&�\,�"a^��0ʑ93qy}�o��c|��g	�Z�C�T�.Tq�����wt�3�M�4�B���fC��WDL? �:�g�K	�wO�-L8u�}�,ٲ<��ꇯ%�@�q����Sc����U�S�[�]��T��R���� Y��H���2i�Y`����&jzʞq���;Zm�d1��#*�G_-�Վ9<���)�Q�S�b�8ō�~�����M�`���U��Z:����R��6P/�q���\^#��7�q�˪_)���V�XF���M�_�4���L,`<.".Ck���{ݘC�6n�8��N�Έ�?}R�L���{c�8��o�C�F:�k?����[��f�����%�?YF݈4��+�n>"I)��r�6�}|v靧�C��SB���<���1�c-�
gp��ا���l֒���X���uJ8n��e7P#;��+�4�^����J�)'}�F(/\�YKA�ϰ�s'c���,�RsI$-9�9�=}���B�a�����N{z���U���]w�0�彭��n�6D�t�V5���P���Jw��:��g�[=�[��)�6	�8���$F�����n�Iu�3 ��I�Y5� �n�l�L#e�NL���s��lR�J��5�O!�z������,�&�4n�\�:v�-~dNT�]t�
�DH��U"8����9��.��a������Weͭ��5�e���Ge��vB��V@�'��q�DOq�I~]�>�:*��oH`F�+����dr~�ޘ�_�`p�n�M�aNp�}�xB���
�Aw�=�q,㒆�y��f�l尬���^9fGP�F������z����7a���n���.G
X��S��$eЦ5��]u��n+����V��i��mӨFK�(΢���t
nΦ�2��;�GՐ���Z#4�D-8sy��y��ǂ�w���E38c�WA���/~Q��;�c��� ��B�`j=��W��2,�1�9��fc"��T���G�l��Z2X2�x�ȝ���t���6-x{���8�����R�?+�<����Y%wk���%��v�%"��pJ�Cǰ��N��s�y���L���c�]V���7� *M	3���=wJ{2�rח��Ύ;�a��0Z�.<ɻ2�u�6��|�kw`�ی�y�f��r�w�㼷+���D54��X�.�y�r3�-��������6���nE�07 w�t��Z����a�<����_�e�:��4��~��OKrݾB��^#)gͧ��o�\Ե��VSO@��0���ޗ��P r�n���������'Fѭ�p�;��x�oޝ��o��[&i��3�m���!_Ep�ǯ*�{ @����K��ai2�)���t2���"��e{%?<�짯�X�ɞ=��-���nS=v�K�i�Q�1j�;q����å���C,i����5���}��LfgP{h2�x87l�����k;����������D��%�_�lo�8״�X��_�-�>�R�즻�g��۹�0$_2جM��l�H[GT��[e閩��L ���<Az�i��M*�g\�t�7s�� ��G%�Gl�ٲ���C�2]+����l�N�,��)�
�S��!;�	�F���z�s�=���~��]�!ѬT��q\���we����&�.� sE��cJ��Ss�`�=P`?�?I�zg�����낆�B[W��ݵ�	[X�f�KH��h�SB���E�v*541�P����5��Ɲ�`
V
�Z�8ٰe7��*�ovbvH�\��vX��/-������Fr���!W8�������]ӏf��ݰ:Ֆ"���p��w��ަ#�T�s�l�4�
T���8�1{�G���uu7O`wBw�Zg�`d����^���C��a��W�1g���,:1֋��2d��ٌ�F�.��A��ݩ��J��+�,3���ͼ����jܨ�D3��>}��)�Z+ח,���{����<��o��l-qуls1��qK������HQ '���Ql��u��1ls�?��V��3�����L4�$����m��À���+�8�>]7�^�L�H�3!Ѷx��u�^q��*�/���lF����,ٰ���T�%u�Ͻl�KcO�K�w�=s���m�Hs)�}��Q�K+`�5��vm�Ӱ�M{!>Nt��֓UeC�A�w޶d)�o6K<?],��ok��w��2n�#��^M�0�2�1�ϡ��?3����z�R�u[U�F�HT�[��YݽZ����e5W�S�x#d����!`+�9;)���`�����Ɇṅ{ez�Iy�w�	�׍�gU��묑vz]���!�c�i��� �)�&}o����H��}��z��^[����V��g.�Ug"&�S&eö�M��r�.�b��%kL�C�Ez���^Ԓ�_���sa�a��Eb�7��}��!�}��@��a{���DH�uՉ��:���N�!�Jk ����w�Ѭ!{�s
��1:r�F~��������wL���귛諘�=�3W���z��t����Ӗ���ٽ�jy1�9��i��4֠�l�U.Sϛ��9mI��I�-�R�u�P*Ȍ�q�׻�;p�J��M=A�ȗF�3�1�z�-�O.��=6�o�'jf\���.ʣ�.�څ{�k�)�N�
��")��ܪɇ.i���X��M�l��sԟ�y��xg]e��*��Q�b�<�2F�o
 T�!�<xY�T�!<r��AuL�U�-��cd�n�j��뜷��7�ۄ�wq��q�\�~}����$;���=�`��. ����n�﷜V�3�˫C�dgFq���vuC�LJ[�c�i��T���K<��=v��0Lb��mY4_�.;��n�����6�FwA�+���i���K�4)��xw��ܶ����/:�J�6��N+�6��q�f�C��=E��(�C��DgM����]7��P�yὊ�<���o��������<�h4}����^U�×��!�Q�"�Bw�N�37��o7���j�ֶ���kk[o�U��m��mkm�*�ֶ��V�����Z����Um[[����j��V�����Z���ʵ����խ�m���ֶ�V������ֶ��V����kk[o��[Z��Z����U��m��V�����[Z���d�Md�2���f�A@��̟\����B;�j٨�*�*K�ΰJ%Bm��TT�*P ɡF���U�WY*!R�;UJ!D����՚t�(R*"�wX�j�f��[U�iue��մղ�g���UZkX�l����Y"�m��FfiV�Z�;d�n�F3SkcS{�n�f��m�*��;Y�mwe̽�{�[`ږ��ڐɥ*�fRͶejͦ��if�µV���i�M}t�34�M�ɬ�V���]�wv퉍��&���ʙ�jR��Q��5(��ڶ�x ��}@����nU���ph�T`���wmp������g'����P1n�q@gk���RM���-,Yٺɵ5}��ݩ�0� |Eyӝ@�mWt�UQEQoQ�@QEQEu\: PP ����EQ@y�}��@QEQ���q袊(��(�{ۼQEB� ���x���y]��f�]�+X�f�U� x z5��woD��ջ����`**��0ݵMR�P�hn�Whh�s��׮���
�6n�6�)��ր���]5]X�����s]k�]���s�  ��ֵ@,d�G t��6��h��l<Ν4��M���l��S[w:�iU5���j��;�C�Q�`Ҫښ���մ�e^��,��ֲ�յZ��{�  =ݫڟ]�
KowGRZ�\:�u��k!i����C��)��l5A+�Nt(V��u��4��A���m`Pj������Cت�T�^����k�-�ݶ�  ]���l6՜.�kA>��m�G�Jt5�{��m�
�:�4�Ͱ���Nt�+*U���B��v�W5��mR�u����g=�:l�e(���e�:��O� ݾ U�:s��/�S��T�=�l��;��j�el((�e���[ ;�wv�^�]���Zl�C�t��R՚�A��p(领���k4��kT�f�7� wO��$�[U�p֔�t]��KaB�s�� 6��u�m��.�:l���3��� 1��iГ{wk'��.��pr��
��[J��6jU��6�Ĝ��� ν/��F�Lҳ��lH�;n v�F[��t�(�mm�S�Ju*垝�PaU��ݵ���uY��5�rhhMW�*�SL�j�ݠ�vZ��l֑֛jV�%lYm+� M���5F�����f��«<���Q��s�:��l�4���\UU�L����Ljѣwm��
Uwptv2R|��*D� �S�0���   �?Sb5U)��  E?�(z�� Oڍ���2dd �(�T�@ �����/~`����O�ٯ��w�����9���>��{翾��﮽���!W}���+Ш����"�
�1W����(�������뙇���Y�_˳t�,��b�CV�$�R` ��L��X)R�1��hTK+2�{{�fȩm00�L��ɵ,�/1}�]��W*f��K+������B�u:+bJ����w�����Ot$���!^CrRB��Z��m7d����n�M���2��R�E4�h�+P����ʵL�M�v]��i�Ӈj��h���r��.V��(kd���PLڻ����5�z��	e���ʠ2����"��`�-��i��i-�u#��U��K2)�v���Y�KD���E	���7�)��<؞��GL�C�\�D�ӏ痲\y��w�v#�}b�{X�hS�%��2�4��+.�ًisQ�ql��9�5V�c/]c0Z��`�����`hčօ{j��vNW`��۴alkӸ�yU�̦�*�F�u7q EVZ����JXG�s������?&F�����,�am�zƨ�{��*8(���-����{�RH�i�%U� o�Sb�B�H&��k��m���+f�7 �GoÕ B�	� �x��i4������n�kL=Tެ�%:Zi����5���kp���:.������Fk,-9�����NI���h�l9�ba,�nTo^V"�ҫt�{b�$����h� �ʣ�[��ۭ��P@���,��6WH����jR2�V\ٕ��%�-)6����+"ܩ��"�E����Ҁ9S2�����:�J��d��Cu7C�vjmjajz��.����6�@���޺W�ԪJn5��Ď�7��umc��ڻ���ܧ����Ơh1���Q%A�"��,2�ו*���{�8��b�T�� �7V�5����� 8_�a�Y���H���܃0㢵�֠�H�AY��i��l՛a�E[en�d�)i�Cq��x�{H&>�I�7amǆ�m`v� �AQ���]�c�
7����$��
�C�����qx�v��!�`�K�ka��Kw�Z��&;�,=WVгz%���}$\��#F��])3.�a�O5��~�!�����p�*�T��h�4�X3sM7J �^GL�:\�1ˤ��W�0ŝGF9bo& ^\�]�/V{����`�fp!D�D�K� �4��Jv+1t�8J�q-Xƛ�L]n\��[.�^*i��e��%9z�xU�yE�ȫr�\ƌgh|�.;A���;�B�y�)�h,�&���z]�[ ���VB�5�"��t2`�����!1kKf:D����kj���g�#m���������մ��F�]��E�7ZS7�K&���b�kq5bݢu=�����v��nq��ܲ����DAt~��8���Tr䶌��Ws\9�k5��7,��蠉t\��Р�T�ɵ��:�ŲRdQ�fY�B�Tǘ��V��C#��V�!�eK�kw,�9#_*х���M�+\kaӸ�3#����Ei<��O6Fu$��n�;@6R9T8+*�I��q����k˲9��A`o�C*�EQ���V+Eɶ�gs%�F
Å��r[�{�e�[@�r�Ҿp�m���7�r�ED8�C��:��7�,��o\tj�U]Xu6ؠf�kSB6ifV����,Y��+u�vS�VX���즅�$��$��[����
��	���/�6��1�i:�]7߱ۈ����� �����ڠ/"!�]�&�U�6%�����J����5���A32� �%����a�q8�t�c�w+n�KNY�޵��]'�N�KB�J�r�ӧ�ȼ��D�DIS����t�Cedifକ�t�;�wއ�0\���a͕�H�P�*ޭA��gEB���2 N��שX�n� ZX���X�P�v��Tga�sh��=eJb��O�����R�v�s*|����-��� �{*T���M�9�a����MD�6#b��n���[Qò-��6����H,�b^BS 3k6�-	Wً&�2$18K�ӯ'="?9Ì/g&V��{0��AC�n��!M�kt^S�,�fZ��B�uR�b)Q�a$*䌆�Ss܌߱��DƸ��=���!M�u5�&^���H��n���hjƫ:��Y*6�E4��V+M����yZ(ķl�m걃� S��;����[�sK�Un��Q=��ؤ����5���
�XÅ���9�F��	��0�-&�:v֬3.|��µ(�U�*jF��Eꈨ��F�������$�Ǭf�-�`�,�'ђ��ǓKc�!�
��¶;®����LVun�J�)�"��[�G��^l���Kܡ�Dm��z���,0��m�+<FA��nj=xpc�bLǣ!D�C2)-��� �vl'��4�mY9�1�@
�࿙��� �Gh���3)]xu<�*�)	��h�u�2�R�m�q�e[��3eQdf��"5�-�S)n�Z�\.m�"��Hg؍��oo[���)��� ҖU��r��F��R��M��%���&������x�	g�^�n�(i+�o�m a��޲�w��V�Y*;��j��%���KI�AcTU�]7O//�u&��#�p�W���ZZ)�m8%�
v.�����d���	��Ǔlk�-Yȣd��iљ����i!�z jH��$��{qc�����(&�5�fERnf=��槆�XrӒnR�H�溘�M�&�����hф_�ѭ1�"6��"�ct�-����bb2:��N i�T0�`�J��olݑ%Y)0�\�vXZ]aF�{�F��%:��#.�f�Q�Ԓ�Z�1Mu�Q��(��.��k0lr��p�Q-�Э����b; 뚨eHn)�Rz��d�z��l�iu��U�噩!Ǟp�#X����+X��3&m��׈w���x$�\tr���L�q�����m`��Jsݱ��7Y��(�!Sf$�����aM=t���ܭ�EQǫ��j<ǟ�G1b�j�6��*	>���I �UeEU�M����{�t�n�k�k�µZe���F��Y���7����@Z�N�ŲjΫ*��1h-
B�0�p�B^n��S4D��n.�f�H=u�J��彅�y�[���J��'dt�X��Pj���Vm�r�	*V �q��FBۑ��[iLvT�ö�!���X��k`�2ؽ�D��nsv��7�$Ѝ]��B�ʰt

�Гt]�Ph�nb۲h�	q�.� q�7��am��2�^ a5h67����
�{��T�m��6��D@���Za���㽻����(�(S�C``��	�E"/�xM� ��D�ss�'�><u�b�9 G����z��#�&5�jV���
�̅�$�aV�F]��orã�%M��{Ct�l:a�TH\����yv�1*6���
�+�tGV�M����*�D KH������y��]�"m
���R�Ҋ������/#-���I��v�f�(�t�y���ahb�WH��%-���.U��7&�k!ḓ�%8�-��L*3�mmܭ�^�L��X��m�+������6V$�Вsl�tE-�2 �v	&�V%e ͊yE�u�q�ZgdL'M�!��0���[�u� �=r��gp�#l�e��'pcF�0J����1B������T��Ū,��ԋuQ��7JgV���`�X����2���׷���էyL�vu[(�Xn[0+xj�;�D۸/f^j�.����f�uv�ƨ���pcË��ٹ��Jb�H�Ir�I��-"���̙���@����Dӽb����kJ�T����7K����@�-)��.�$��)��Q�0<`փS(h���D�N^�u�)X�4=�D�3d��i)$Y:kP���C�6;3�w�w�6@�ZK�T���@sR�ӏF�U3j����F�ӆ��u&��5�W���ks�]�j���t�z�.��ɱ)�kF��[�}�طn�ɇ#Īu�ԭƫ$��tJ���R��C�J�`�V��V�Fƀշ.
4�Yr!3Z��#4M��Z�`W�&]��[��nA���
�'j��l�.�H���j�h��#o���+�i�躒��V�/)Q���-�6(��0�ʁ��8�]����>*c���E���@�@q�J�����('0�4�kBL;��oT�RVI`Ջ{r��M��0������V& V4���p7,^��Ɯ�$�دPov�v.�3vSV2�m;�c-Sϰ@!�/%������6�F��J�u���ؐ¨҇�!��KE,`���K/]8�����8���΅L��F9��sbgFeJTB��0�ƍ
��
Ʋ���-Y�@X�b����H̖�"�+-̛�Ō�W��*Ś���6Tv��H��]D*!aE��!���,�w G%�5��v	�E�lK�Bk.��`�$ԃkR�ˬe4c��#Z�TRʄ�-�ډeZ��C�t�����v`�r��`�.Sql�#ZMn@^�'(KȐ.�K�lS�R�ƞ��4��dթ{�Sы"��bS����f���v���$d��t=ma�B���4}t���.fnP���W+�Gh����3��-��v��ڙAw�l�j�*:5t����ɺ5�Cf�\�7E7)�P	ZX�1Io�t]&��C�
a�t�e�%��Ŷ��l@�E�A�mJ�r�%��.k��dU�F���O��巏^c��P�v��.P�V-8���	�f�HL�6���l����J�qyҴ�D���]���#U�)'G/gұP�3(8�`�&�,EJ�[�V֬�d5w8M�X5�@�O~�6n��@�mb� WX��a0JR�]����[Q�H���Բc�W�m��hj
GPЬ�k��X�okhu��6���/
K�"JË/
tV�Ӹ��ag�^f�2QGT���&�t�³u�b�B��~'[6Ag�խW���q<�X�m�u�_̀��T�e�����+��5`�!��hN��/*	��b�(�Y�$��+J܌�`<�Xutb0 �X@��e[ƛh�%��7i�lm
�%YWv�^��h�V݂��dؐ$�bͣf����L��"���:N�z�˷�^��!ь�d�tg�Ż�C^����>"�f���GD9l�8^�t��]J��ƌb�[Q���[�j
L4�'PK*�ۛm�"����X+CwZ�#�6�Ŗ�vR�4N�V�N)��h8f*r;`8oSJ��ct��cc`�a��j��n s
K*ј%��4�v��xZ�i���)�Hn��V��yt�Sh��m�F������C����cV���w�R�-�i��J7j�t�e��z)�f$3C\�2�̗3vM�v�x�ٶB��GP��c���%&'��9���t�=�*q����NM����^C�i{���MeaH�g�x�Y��8�Cܦ�9N`��F��J�ьn�x���d��PK4���ƩmH�	Wl��k�wrA[��3�A#����8uWu{X�
f�'��0�;w��8_a(�OR�_����SV��Z[[.Ј,U��{gF���q�l�㄰a��K������/c�J=���ŮZ�W{���a-V�a61�s*u�N��0^B�KV0T��\�j�jttk�Y$$�r�X\�*bNЛ6����%��ۈ�#E��ɸ�IL�cf��lT�X�;�q40���藨��"�t�������\y�%E�Uj〻+��B&B��K�y��/u����Ĵ�j��n$�҄W%֝5#�Fޱca�t��5A�A�:.�zr�\-����,2K	N��6y#d�z�['t5x�%@T�ؗ[P��V�Ù
���`�Դ�%�@��QfQ����mL���m�cu��d{m�K[��ԫ�L��Э����X��ں݇q�ђ��ˠ����^�ͽ:QyI3�f��[�-j�*6j��v�f��v�k&VvDR��Zص�E�����z��.�w��Ԥ��sT-S6��M�n�Nը�9H�B��f0��Pߡvh15��� V�eoS��+6+n7Ewi�3m��,�r�{�j�]�
m�������R��5*Jֻ��4�I�Q�j��+fŸԼ���%An\q�+����Ih6-hhTܩ	x��.<���TIy�8�"|�*˴M*dn�]�j�ms[9��@���:#�m��4]���U�jP<�J���xQ�٣u 8雳�,i�ۇEe�����mRx[	�5�������TM��R����aj��@b�]��x6I�	�a^�)�6�X]�e8��Jyrͦ��M��Lm&];�_f�B[k^U�����h9"��b(ܺ�.#gcaڠ�^�zq^Psf���q�E�&�K#j,��U�h_�=W��%˖�njJ1+vE�6Y�i�ȃ�K�۫&��QKn�m���]�q���m�j�(��Ç&M��B�iV4�;v���3�%}�Y��,�A��ψ��M]�NTǛ���XI$e�GEe�b�;4�4�o5��uU$�
9Y�T���`4�fЂ=	HC!�%�8�ۨ���;I]�g��Z%�����L$M̠����1�2!x�jkdHR=���d�+j'0�1���)B7)<�J���I�hT�\�Z��v����h�%�wH�cV������Kx������۲BDy�{�FNz�Ye�m�f�+ss��ޅ=�cw˃�
;۵+�s{Z����>�ݍwJ쒱�7{t��C�#V�f.�L�>��4������wc$�]��B�[���V[�_c˥%&�}��[7��qp5�킕%�n��/�9Ol�by�s���Ѥ�� %5C���+\����e>ͳj�\9b�a�k�vsy��� �3�*r��z��p����Co^�mB�Q\��e/
��/��x]�ĳ]��/�.��|#��og��o�㸪n�UBt+":�}zmF|���lt?p����$��rʙ�Y�������ӎ�]�z+�A4�뵜�8u�u��&(a�#�Rzivcy��Xj�վ�B@.4w��y�q@�$WM� \�3��vVt�&<�ޫ�D��L�N�fkk���#w*��H�ݙiժQ9أ7[ú�,��'�4�QNg,�&���%PZ0*f��O�-u��I����;�I�bP!�Hg�.,�t��K�K�䭑���39Уك�sD��ʕ1K���v)�����#��[�U�"�%و�����7W�YޞZ�}('�v�n|I� ivf;���5�����j矸��&x{L� ����K� ���/�~�O:���}�k]�f��H�&�]�*5�u50W�[�9r� ��A*4.��n��V=��9ԃ�@�ճ�g3k�AI;	����-[����v6
W{s���o�筟>�xxX�o�:����-�����u��v�cl��]���x���n�X�����38�GhfŦ��i{*�[��s�/^���/T�3L\���6r�Ş�:�Yw�l`0�K�V���UL��0��2�ƴ��{K�݃/��2��kE*}��'YC�Hs�$(��OCGE����,��U���*�RY���S�}��7>��uE'Z%�GvJʚ�m���&qˬ�ٝ�[���ou[ZU]�'����1-5�`hgS��5�(�hRֶw'i�ǋ-���hQq�����P��5�T3��%އ$%�����2'�u��P��W�[�.$�묮�DY� ��7�6�6ݛJ'��mۻ�\�����C�>od%s�0Z��2����0��1Ytݹ��:��Aq<(T���U��tؑp�s�,��'��x�.�i͎���T�o	��.��ے�u�87z��L��t/��Z�������Q�(c;�.����H�T��1\i�RT��.�z�v�/k�'���n�ib�/q�i�ƹ�^;_e��oG�jF0LN�z���6��]�+�\�:�Q�]�85h7�+K�y������vZ��}����F�+�E��V��nS�qKyܹs�A��J���ՐS9}����]	1�.��ܽk�s�YH�PR��ߡ�����u�4u�J�Z�2hqوa&����S�.2ëˈ���}�w�1K:u5�a{ω�Z�9s����� iv�$43��������Z�5���&Wh��Yٌ�q�@���vyAp��ͪ4���t#�^N�l��p��Y{���J�J7\���i;mf�Rk/��Uؠ�Z&��+l	75-�);����Sj�oL=s�Ѳ��#�I����8%�M�VʌL��T�|��0t�(+��FܬwW�K�'�]v�p^^���4�������FV"��J���+)$������#޾U>T��V������/������/-
Y�yqɤ#���Iǘ�6ϥkS��n��-�������� ����q�ubXvn�mLlgt�40�&me�f.:�e��ݥ+���L��Yc��lQw��,e�L�B-�KÕ����z���Y��k�K����;02�ҠZ�10'��9��t�Yټ�R��wsxt��J7�u����vv��zҨ;��i��06ޯ1a�e��Z=��Ү���"��W��ſ�	̙�:�}S�9�����ִ�G3�k�y�7�#��9��P%r����)�N~ܩ���{�<��x1�6��3�bE���7��\09ݷ�a�V�x�k���[�<�����;՜O��WC��X�."�#������H��N]W�[/��3�F�r7�B��Af]����u{�ly�	��jƝL#p�:��]�uD�;7��:{|�Vs��Np�q[t��o����F�C��ۼrz2��9�6��u('B�X��gn���V�^׭9�(n��Q]Ƣ*D6\ۻ|7�]|��i�k�,,W(<���F�e���z��AT3K�:飒b��%c����utȹ���J[B��g����5}ԔE��yX� wQsy�r�On��R�=2�V-b�Z�ښ/�۲�LD}q����Z=��F�a��lV�zk�β��[�"^���y��'	j�B1���K��!�m��\ո�
���GP�L��� ������i5�I9�9��b��w}��F��n�ǁ���Π�������_0O9�i�Y�l8��޵ʎʅ�-��vî���=7�����z��tf�{|��-�Ff<�tm�]:�;g'*�Q`���uʅ��}Eh���i\Q�OͶ�oVH·�v��ߡ��|�A�J$����݇��[C���J;_�a3�,�i�꾿�u�PN⩨�Yk��Ե�"MNi@r���ҷ'��d��ohh�\�S-��@t�uC�UUm+���{SXGk*���b@��)�J	��;���42��$�՗�tTDXD_e��Zu��;3�ZM���eRVn3�Z[��X-�W�;�lݢI��gd!�;��%�;�Nq�Ǧ���p��Ӣ�A�-,��`�t�'6��*���;���}��C;�SA��ѯr[��곫U"���μ���W:�'��y���Mh���������Î�ǚtj�}g�����P$���Z1U��Ӱjާ���LPE:lq���Ki�P�Vڭ�[6v��7�$��zQ��5Xh����{��O7���}�c���f���%1z�gz��.~0f�?�.����z�W��hWj��y����*��T��S+s����#�<x��.TD:�{	�����}u����5��/��^����F��/�]���n���{�,�z:�c|+/.Yԩ��/�/Ӻ�ϲ�����ڮ]Uo�ݣ;���e�LƯ�)"|_Dx�*��g��-����$���B�`�%ٶ�Gi��Q�tn�Z�2e?j^\/@�޼�As��½N�s��Z�M� VjZ�b����"��|�$ �wg'9ڮ2���۽Ԉ;�)��[F��_������ԛ.��ۥXWc'\��8�<�OemwC�Kk�AwӄkJmK�7h����v+���v nN`�W�ǪJf�q�	!�hR�V@�.H&�
�6����e�x{;s=�~���]���qSWO0n�f�t͓�g1Jw�
���(
�m��|�%m$B��β⹭�pm/Lϵo�6*4����\ moY.��}3�n��Rfi��;n�wT���GO-�{�r�/��u�:+"���$����n�wj�U��X��ϊ�.�ݽ��\�¶t�SR�ZgfB�	�|H��վ�5A�h����P��>Қ��tE�ͪ"�VM��b�₰U�0mf��/�����p��٨�Fs�&���2(�i�������#-�eN�̋vuȳ��*��qIn��6�rF� 8 +���S�]��Ҟr][ݹݛRr�\�����S����j���λ�Q�i^ئ�V��5qs�l��uh�����\:
݈6��a����s���/E�`'�y}�G�ql�U�"�C���*��{&�n�9��� yG�����F�.�M��|�'Q�g�Z��	`a�Bi*�9@�� ��%.u�Y��l�v�tt`9+AWu�7F�x5��g��3.�b|�s*ec&S�[9��ⲝ'kY	��d�tT#�4Ɯ��Ǭ��b�n5�5�oq��`����K/��t��:�~�4��R�)��֋�X�tĝ�ll�j
�cC�6��Ӽ�qG2āG ��r�+�[幗Ʃ�V�Mj�_'M�,]��w�mS19��:��h���p;�ӃB����}ڱ^�򔘆@HmAI4~�/Ne���A�ev� #��u�V�1���	ޢF�۷*+�9�{��`�7�%�;����˥�TN��n���At�E���n�� �i�2�d؂Yo���i���xs��`Ww݅e�}C��l��y[�z#�"�`�YBSW!F�V��p*���0q}w�L�KB��ᏺp�TX:v[:��A�_7l�p*4c�,l���=��r���2��
`](΋U[|C�p�w�J��WN�7qˤ�����.�����Tj����Y��W	R�Y��2sff�;8�d�����]����m�� �M�H��e��R��3s˝��Gm��S����s��c8қ��ŗZz�i8R�Ϝ�Ι��8�p�B�ٮ�p�H�Ɏ@�O�֛O]�b��ܾ���k#%7��n�a�5���M�lͱ�:葑�+ܐN�s�o.�ׯf��6��.�T
��d�p�IŝGGuy�!�mE�<��\Y:�Q�J�^g{��(�Gϱ0+r���y>)X��F��uTTX /��^�p������cu(Jgz�]�����op1��i�����5�v�
֖�:Ȭ�]νq<Ѐ��U���YR1��4�Z��R�V��]q{����c�?t�pÃ5��b5���;8�r�����j�Ov�W"lfZ&qGZ:4c�2^���}�]��7۽�y��栋oo�	{� 0M]�d:��+"^�ʍ�$�l��nQC�;-w���$�١���u@�d����̺���(V�"���(�s	 Xt+%���OYj�e}ƦॼU	���<2������Z���0�i��pO\����]Ԛ�R^��8������|T�Yg�[^s�!報IZ˷�`/P��6|�{x�Y1p�ʾXLG�J+�[x7���CUx@w��~w7DX�v�S'D���;f��;9�����*������Iľ������3	�|Ԫ�bn���X7x�����`��۬�����Ԑe�r�*3�ɼ�ol���f9��mӁ�r�yw���M���	��|SY���9fD%�+���8�+gq��sZz�e��v��ob*@��L�8��aeG^A\�TnJ��B�ݻ���2���@U�[ l�U�E���vC�P�Y�wEܷ�+����{���LI�8�;��񨫾��!�39n�J�lP�/�"��v�v��U���e�u���`���.�d�k-9������}Ҳ� Ԥ�>�2���J��0/�\�O����%����Fl��}ٜ�M>6�nY6���e\�й�;TN�/��OG�&��p�Ͳ�7}�v�2��R��lo��㗦��q<ct$2=ڷ溼�^W)�)OC/\��N��B����n=���X�{�S<��Y��(�G]Fj@�@?�N��oϢ��Θn
�t�Y��`�I
͒<8�K���5[
!6u�8���;��5��0�1v�:��� ��rk�moǻ�pf��؝x͈iM�<�i�����`�Aq�'�t=[J�M꘷w:n]^��� �������J��w��κ�i�8���Ƿ��!/t#�E�Ayc�ĉ��-���-��2&�q��� ���yw'ucy�����@"�xd�R��&��{��כ�[ԅ��f��G���̐J�o$������&����Ƿ8<��Ͻ�!
|7�E*��ۦ�\�V���#ٙ��0�{D$���-޳tm��AGv�C:[��k����u�I�Mɽ@M��=����sԇ:�=@�ߐ��=�{�q���x� �̩v�ߩ�˸��2�X��T�LjY�!;��V�h����J��3K��.�s�y��b��2�=�6ƺ�3!��T�]�4�:��j$�6nv.@3�ӏ��,�s����w>�лO�����z��{��yI�EHĆ6y -�#�T�j�mf�m����ј��ˮ��c_>��RƶeIر�Y�N9���\��n�4N����5W�~�֮Kζ�|Nr|	�IvE�<u�=� ��+F��ɸ�f�yGN��`��k��ɥ���F�^Xzg5�e����!���/���W��ZE�
��e�$L�k�[��v*i�Q�B�Zf)���fͮS���Ү�Q���ͨ�+�[�����%
]Ӷ���l.�{��:c���H�7(�_I�_*3���+��sE�,xS�4��u�
��*�l:8�3p�:�K�B��L/ۜ����������*�r�P���mN۸���,��D�y&ҽ��9��DyW �n��3Y��X�[�_*��6��xN�.}��}�Wj�����/��϶�=�=1���e�P�z�F�'K�ޑ+:�';wP�m|���,c�� ����$��0�S#��50�^N�Pm��I9Z �d�9�� j�32gE�X .y�V����w�Qj*�r�rPk*[��dS���%i�`�&�f��ގZ���P2�>��fv���������s���2�������ЗG_\rS�ֳS���q��k�)���[G�X̛���ڑ����
���aM$;ӌ��ք�.J���W���Y�z�]Gn���Cu��մ,uu����,F�
�q��X�,<9��;Zn�2���;Ր��{v���d�\z��.9�|��s@�f$1^�QE3+y�y��7��ͣUju+�+Աr �^�/�{���B* ���:�����y�_��������ޝt�wxjpOɃ@T�fs\�?u�ۊ-�'�'J1��Q�=݈�銓8�tB�Ẕĺ������WF ��u�k)��u�T�F�Q�79wm�ʎ���hGyQ!��ս�V�¬v2��%���Ѩm#�V9W*HD�P���o��gV�wYY�-�������CZ㼺�w&�]�u�l���}�-�0Zw�]�c�?�H�H䉈j�&�gyh9�#* �ZFe�73w3B�����z;�� u�u8uGHi�� �nwc��l�u2�,y��8�Qqs��-��m���Na�K�9n����`p���/�+q�Ǟ`���L3��O�˻(���B�������dT�YA9�DW����� �1P���h4��Q?v<Nn����3�-�\ں�jb��i��)���3]{�Y�r!�-��6��t("g�s�M����G{u��c�=;���z�˽3�격�׾��wn֛R�t�Y-ݳ�kq`|�ق���:D\���0ޝ�|Y� ��)��S���UBg|އ��J��k]4c^P�ǡ�Wܔ�Cuq52�޻�5;hǜU�7&!�H�:�Y��y��}�z��=̓S����2�*E�K�g1U���s���rfL(���Q��wh��h��v��G}��g;��GO� �K�w�-#�_N���×iK��mǫ(^X�f+z��mT2�4����b"#��6u�h��nYD>���pR��OU�A�tؔNV\{�����`^�Eн��䤡R��L^H�<��`є�I�C���h�k[��0��^5��������Ί{�c��UmKM2\��t�i6��j�a��c�K�엷�B�j��l�C���\vg���}4�F�D���˔��ʫ���ך��V�������]X��zhR�1�s)��Gt��Wʠ	mѝ�kA��R��8�C����׷.k+iBJ��>����{W�'8߅�iR�YR�O��oompq�fe;�R�]�3uuH�o��$��ޢhy̮YrU�6�I��c���X�]��53��U��)_,ӛD��ޖU����b�޺՛�=%�+Y9*Xۧ�>���VU/�9D��k�	7�B�
���G`+��wn�c�U��f^1k�*�ƪ�.o;���{+���A���rR��Y��V��f�=�0X�-���C�8J���A�6]�Cc����M��k�}�jf>����(�q������.O4�"��c���d��r�ͪ��Œtۦ^��v��u`s
`[;~�z�E󝻹�2�Ix�;[]ޛ�J9�^VvN/�F��qy��\��Q�:�K��X�����F_^ώ�3�oj'�n����ƞ0麺�����]@����Õ��qY�z�2\϶�7R����^��JᦘZZmn��}�=w	fY��L���ݔ7B7�H@lt����.<�p�@p�zo!=��oHV��ɥ7wW� �Zk���B_(Eq5b�x�_7�������r�3����rkj5s�f��÷����J�ES㠡���n*����8p�ɘo�o���%�\6��.�QCJ���v�7�sS;�����C�l�ՂL���O;�&M�Iux�Zau�c^�Q̱V`�{O�4N8��EB5=�7c!�;���q�t"G�9��/yn��ك�wݜ��(]č�}����&c�H��Ʊ8�GN�j`��Ϋ DT�I�9�7y�OT���;��vu�8]��!��V�tNMT@U�}�@�3r��T�7F��PY��]Y����sR�� @;�>K̾�Y5`e��bЭn!o����Kt�Sf�<�-�ӥ��h�[i����(di
P�l�ou��L�e��4*���2���
�iRF�wiS�&^����*İ�/2W��]l�+Uh-�.�K����'gt�W��z�]���:�Q�ys�����q�T�_L*�����b���[OQ�Ep6��4� �@'/	U�6&�8��p�r ��̀�KxpJh������î�	r��D\x�3�ﴷZkf$NP�Rw%z�6�� 
�Sy�7P���{5mg;'7Ue�PjR���h�]�L�pqQk�K,�H�윮��Y��}4f��>����&�G�u�v�:Ʌ��l�^�^�Me`H$��/�K��X��p[x�'E��+bk_�w�)�\#��������ec���#5rBE�t"�J;	�����6�ۏ�Lz5���$�o��\F�o����!�w]9V;����n���.(�-�7�%�+�q�Ѽ'�v`>���r�
4rƟ�M[���V(z�n}�,;��v�R��<w��eԫw'u�؈�u�;M�G^I.L���GG��ޠ���v[3L�;f��ga҅�j;t(�#�����`�yj�u�9:C��[`�Rw��V���x�j�`�\�؁�<ݟ`���*��[�9�o"B˫�Mj/V�ת����"�tE!�t��޻:��.�(w#�RY�v�6�����g[y�cVz��E�e�ɉ��B����C�O'jQrP����^\�RE�X������
;��>i�v��ь��|��n�����V��6��털b{�xe��(0H��u���"5e��Z6ַ�w���3hNNM[7&�P�o�h��ϫP����qvPԉ���y-�v�����WV�4y��X�t���Y�⧹��I��L$u��wf�L �u�������>�g��U�kHһ�X@uӶ�������!!8�Yj�٫8���8��M-e��S��sڰ�Y8 �����s����\���YոUҨ˔^��#�e,�ٰ�{Ǔ����ϗ`��M���$�m�����1���%�g'
���������S�=���Y�l"��R���x�ɮYkk6�ٮ�g�4�,,q3]�v(�M<,9����+���G�<�""n�w��	Oz�8�&���˼�9���ˎ�X��$b�v���{�t��9Y�o���>7(�����ۯND4-�جo��v�3	z�k{5� �5�}s't��w`�}�4"��4uWG
����bZtj�o(,�ښ	�|~�P�8^�ڹgs{�W�v�$/�g%�Q��w@.����|�&�1�8��E���c�Q��.��fv�������޼8ң�뮝���u�9�m�̉=�vO�>��nG!r��%ԡ����{-�Vf<bJS�����j���M����f\�0�W�����[��������d��8!���Kvgi7Ag����-��o��<�g���QR�)Ј�lm�>���9��8�G�H>���`�dG��s�K��D�}iBJ��`��C'3�]ci�+6.�	jX7�=��ɜ��m_D����B���D8q0�פ�L+�y�j7i�;P�ARp��y}��ub��s�i�;��.[�$���s�y�*�)��6Ӏ+9�z;,�!�f��&�췖tW���/-z=�'����!�j��p���V�ps:�x�T����H��6��x
���.�.�7���s�C�~�*P��m,��r���i����S!i��}�����ܑV%	#w
�Gg�7�f�s�sSηnu��u�/��Ѡ��
�^�/8�0o%�x�3<|u�i��D�Q���'n�@�w8��%�{�쇭%�8�v3�k�<qm��bg���J�c��wY�U]��[q�o(ޚA:�ֆ۳�-H�\礶���[:�Ʃd�����r�0OIٝ)��
�&��am�8a�S�@ fqN�aK�̗�R��n���=��v��(����ٓrۋ��Y�
��N�D��N���]O���'c̒Tڙ(�3z��.�-�7re�����[`3��R��=i ����)<��+t�*J�m�5�N-Ɩ7��#kX�8�͑A��ѕ'%�3�pγp�gF�h�.+��m�sڰNZ����<8�F��8����B��IV�{kf�iڜtB�k�!�it�����1{(L������T�*�Mo:Cr�Z&,�g:��̠��LE�^�'����d�#W����e�ɼ��L��Jؾ�=˦�&3���62�������n"'@���iOd�-`���c��^}A���nѨ i���r��I(�j�K����惏��M���ve.�.�髧��:^:p-Ql,�\�wpW��Rf=1�ŏ��8k:A�H쵏(-�ݰ�uE݇��A���D I(.�b�4h��R���>��y�7M��{}�9��{�87{!�Ӹ���p�r+�5�w��9�}%�z]�h�(�gj�E��(bhlÙ6�B��],̂��=�	����u��v:�ު"<f0�d��	&��N��q��U�g�D��8@��Fa�qGBb�4�X�X��ͧ%�JO�b�O��f��۾͂���+,�k	٩K��\&��q�]�38��hs���{������Jق��زW
z(EӲ�寣��7+MՕ�Jo��^��q��B5��F�fu�6��z���)��S��ZV�_`�"3u�u5:,PYd�z{��:�2�.���Ti�S��5R�O��|*�Eٽ#���v��V���
���`�\����:�,��h�O[e��g���JR�v������4{�K4з�k�o���b��nG&l��uH����Θ�vd�t$�d���X�|�L�+0�7E�v�[ZŔa�P�_m���7n�X�j��kenΥ*j����K:.ڣ�⻴�kJ:���r���
J�@ u�w�bX�mvp��[�;�K�-Vmgj�wl6��Z�9�N��xE��]�A4{�����8�}��n�[5��l�X�<܀�ݸ�+��,r
�#�y������C<�i��u��]��W-�b	Z��\�W¯"sN����rC[�*��j��r��y&1k`ŷb�̾���׵�Ks���n+l��h��f��G���������v�ͻ�̌�qV��k�����-������.��K=4Ҷp)�m�i`	���5��5�q�[�u=x�F=5�J���A�N�%շ�1��I0��`]����!���*u/�nY�iY�m�(1��#�j�G�|L�X�5����z�6Eˬ�'��Aް
3O���i��8=a��;�E��v�^X�F�z��C�B@�ǹ	��#��,�'ݛ��9洡��W�F4s�7�v��}eNhfebo�onki�+nå�Q���j5׼^���y
S3m) ��AF�lT{"��{c�\�{tFVJ��n��=��6��2�"#v7�����t9ˬuw�5j��6� x��s7-��1�vsU�Q���}i�K9�����w� �ȩ	ʸ��H)娭r���Uv��ܴ����	��3P�g�u�*���m�asp�zm/��O��8^e��jw����8%7�R�p��ӑۖf�Ͻ�3�z���R�V�[�%�7�1
"ԩ6h���Gs�3�f�uN�<(l
Y��Du7[D��w�WF8՛@u������{ጷ}��>�u;4�e�0��aV��phP��s�1�vF��I�W�L�9�zҲ�i��O����*ƶu:�U��;C�jM��普l��"wh�h��5^x'��z"s'��/1�-�.��"^��Y���`]<T�(H���CI��'M��y��/S8�8��Mm�@S{�%�{M��+�̄�j���7M�a��;h�%�1 ��K�(�[�-f�MX�om�~{�(�gtF��7ø�o��4���Z�OE^S/��wr���|�/K���`�(��F��N��KP�Pc�iT�yz�з�c�å�v_%]i]4�m7T�>Y:�c� �J�����oAT�'g�N0�81�=CvP��8��Ҩ^Emp��C���Vx��r�h�ֈ�q�o�gܫ��<.�D6����htu:�Z=SX�j� А�=z��yw�-&b�ؗ����7��+Oj"�0�/Sy�� xYks����:����۴N�wS�V��e��?����v�^�k�x7m�i��|��p!�z����!G^<*��v��ǽrs�;N�ż3�T�jwB��'a�H�Q���\����&�V ^�����x����l����3e��_AH�]��1��y�Z�r�iy[�lIebBh��-���oi��u�Wk�qHe�{�$�Iq�5����Vd7���OX\{`{E�wҋ'*i7���;+p}z4�4��� �5��`��-c%�b-�n����ډҤU����Rۖ�<J�cE��:���I��ۭM�J��Zl�+y3�c��W�R{yƻGk@��1b^_d��ood�3%���,�R}�����ٴŒ�xc���D���)y�I��}JK���{�tWP'�����p�x��Uyuff *�`����0�VDԳ6����pmj}���Y��zھ��osjJ�+ �D[����c�I�F����36��{�\��X�E �d<�����'j�`Օ2!��TC`��7�xMҋ�KP�$ݭ�wƙj�BWok��ݾ�@o%wgr}Vxf3H��.SW��c��vт�{�^�CB�3�]�r6�O�`����S���{���l�(}�WLW\�+�ڵ1⮃i<��Ԥ5�%i#'fpĭ��w�&s�^��]Z��|���{�^���<H�)��������E�K��,�(Ձ̍fP���#uȫ\�D"��J�7	F��k�����,�_�_W�}_U}���ؽl�r���="�W]ޅ@.G��739:��Z�/_Bh�[(q;��
pP^���}qa�jԆ�c�dH$&]a;��u���I�Цb G��w��b�[����\�*���K6��Y��c���� 7���Q�1�Y��8���<�'���0F�`��V�!�g�3��gو��v���#�<�z�[�kn ����	���^<�0��pE�deW��;���X(�s;�"��'Zj���۹���޳4%޺߻+xȚ�Ad���g�Z�jfp'�l�������OsqG��Z�������z���u��Z�gާ6i�T���iܝ!�R���HM̭�K�W}��w�5�/�E�K�W+�1���6f�l=oN��D�F��V�nͤ�����TS%N����1%�p9��E!p���ʹW�z��	��|�^�[z�H���w��~���U��G�&��-�	z��a���B�����4dn��]`�J��} �m��>�Փ_hxs^S�{={ϐ��5Z-:�0V��w���N��Nb�R M���gNҡG-���A~��˙qt��r,-J'��fʄC�X�J��:�5yW3p �e����#ٴ�61sܶ0Ag������e��e���V�&�n�?��;�Nn�P!�M�ۼ1ѝkM�u6�}��Y:q{�3�.n�7�>������K���R4YR�%��.f"R� �V@49(P4+@d�@Rd�R-��
ģFBd�4B�PS��d+BdP�Bd�Bd�!B%(d�9!�+�@9*d�BR�JU��"d#H���J�	��	�VBP�)�!NC���!TUCET�(^�y�����T�f�����T���0s�8�;t2��bQ}���z�pr��ê����d���&&ծ#y�6���G���ݥ���GV��+�T:��?3²�8*+;;�8���_��zh��{�/:�w��m�Eç��,�`��C_xe��n����ɏ��3�${�x;"�d�<.�;�T#/.���u,����!���抑�F_�_l�J��x��g��^J�T'b����V+8����f21�]e�+�뢺��9��W�.���u7W��4�sOGm�sa��Д^�5�c�+v�ˉG5x�K:����t���sY1yw�s'@~�����bלj#���3a�fĮ������LL�a�ޅ��sG9u�����=�����D���4��f���➲|w.�U���{��c���*+׍�r����}���v��_1�y�O�V.���Sǿ�>ެ~��_&3��T�4��	���s�9zf�U��^oypG7\�&�<)�������`OŠ�v\G3�8���h�Tۏ)��{<6Ljy�ZM��t��ֿI�o�#�9�)��Eu"T��k4ރ��q�\;ֶ�P�+3K!u���>(�����fK�"��x��*�o���u֒�'��]������ui���HU���X����;��Ú�#cr�S��N9��m�w��(,��(�E�}.�M�v���w�Ş*>���f��[����uCv(л �==�f�WP��:3).�6ϻ��*V��^쮽�Oz��J5��c!6W�Yλ��Al/>���l��}�ߠ�}[�ҝC|���yY�}I�-��1K�0�ʼ���D,f��mjs�x��c��1[�	��t��E�6�iҜ	Э�c���E�ͽP�lK��"a[<*욉[1l)�����/����
�1>�S���f�XC׻Nnx+[={��J鋬V��Z�D�{mC������K���r7b�8�n��#d:�#������EV'/�lL���\����ً1� ��ܜl6��1	��[�#n�W^0���m���m�d �p)u�B9pS}%L���Yv1�b�������f�����'Sl&'ʺj��y[l͟dJ�#3�"�9�K�٪Zg#o7�eY�92�u�V��;��%���.m����ʐ�����Ն�'vs
)�ٙ��oۈ��fIzum�D��΢�]E���_&����d�5	`��r�DƧ��]�V�'��u��\�Sw�*+-�.q�͎���r<�p�ӱP�8�QѸ�e>�+pھ�i؛�Z��Qx�tg)�ή����r˚�	b.^��h�9��c){����~S0���7��_�Z���LVr�+[��rʪfq��+'u�}������:VeBx�o6v��>�����0�j55�������庎�q���G'm�Y�����V*�#h�§k��k�3:WV�wUK��Sˋ}�&/Z�K�[�~	�z��z���A@kk��toR�ؤ��p���U��N:��.��6��%����)�Zc�k��SA��e�\�w����n������Ux����n��+ޚ���΃nP�w��{�G{��7�콸2r�K��hT�V��~[W�Y����8#B��ۿSn�3�*D����`.^��]�,�o�����ΪD3O�
y>8֖˧;�y���L}w���7�#�^�n/T3����"}xC���]�R��J�uՀ o�]�m���ət�Lmۛ���׼�ӑ;�c�"����C�5'NqD缾�f���Ty�GW���� ��"VͰ�"�f�ҰNf���|���]����ζi�nv9��j@VƶxW���������;Hְ�;8��*M���V����[	�����#d:�#�l�h������(����Vq5�K�uح-��q��X*9�JwN2,��Z�'\o��S����v�B���7}�E-����|�Sv�9��+����i�d]校������W�Q�9Z�܈�uH��gT����-%U�Qi�usFkCܷ��f�^q[zg��Pn�SeF�񨠻ڀ�-��:F�^����J��;����Rͤ��^��,�U+�6,T�ӌL7Q��t�v;���b���5k[k��}��r[]�1�O�ˮ��-�� ԩ�ܺ���q���/��O-V9<�{�T��U�ט5��`9�27EOq;vz������6̥��ڤv�ȌϪ���2����pf���tz��o�>��iuf� ��,[��2]Yn����b׾�W���h�:�OM��ҥl���g^�k����'Q����5n�S�u�>�+Y�ڂw���Rb}|��ZS	>w��+zu�=��cDK�eֿJ���^A:�\�A\&�Y~ħ��e��ъ�	2�Us��{�s'oI�UD2�Ex>�1�k������\TTK�ie\�l5ǝn���T��7�Uy�V�ym�֫��.n5\j����ۊ��b���������S�'p�����^���^�	�r[��z{�o�������6�ҳ�w�ۮ��Oi�¤��]�C�p�3��VrT��gVMzV�^4�N,/��B2��!;���c�u*�G~a��E��P�y���;����:�[���^����)�'�����y��=q�(����g��k
2��b��̧x����m^�=���C����Pn�7K8���ך����ڊ���9�ǺYʮ��G%/6)6g��wH S��������w&}Ɨ�B�u�+����ٓ����<��p��(�I�[H�)�i}�ON=�#`���Ɠ�V*60��$���o��֦�}�R���/k�B�']�_[��m[R�w�"�ܘ�>����)��3���N��W��U)�xgz��x�<����OYn��3#|_�s��=����F�)���jW:��sb��/r}���󙞬�Ǳ�!y��+�xOD�;�].+׍�Dg!�j����i��y��. �ہ���;��kq�<S�;^=�}NN�|���><�\iO�*u]k1�X]��:�\�f-����Y��)�ȃ���uץA��b��!V��58P�2ᙋI����>�����7��z�,�ʂyT��+��]][�zi��f%�[݋u�~�N��Oy��o�uy���˯	���P�z'�mE�4t�O�"�h�{��wg3��lO�ߵ��{F%6T\�]�7K�ձ[�Z^[��pc#�]t׷���=/[��S�N�By�Ɛ���]��2:�q�ǀ�0�pS�{;��Y��mͱd�Tu���l�c�[��cΫ��I�ν�1<��3XЅ!ߌ^���'���;���.K��v�Qy�*�_U�!���hWl��X�
u��4ڼ1��Z��b��Q���'����,��>~-lf�����ث�=C����ڷ�Y��݆$6�2/�����f�s�>��i|�/�R�[Ƈx���w77e���q�v)'��7��'[=���J鋬VƜ�9�� �m9	��Z�=�D���[2�8Y	ŵR�#��6?�d���Yԛ���oc���[Jӎy׈��c���6�qx�Ѧ�c��6�ы����ڲ�[��9۟V7Qw*��	�p&�1Pݭ�1֛9�+*�$����ܘ���2�Fm@Yx]dVSW�**2���Q�ا��F=.����������q{�ɍ�Q<��-ޔ_�ܩ��K�S��M�9��[��\TJ�糹iW�1�j��f���򙇭��r�P�~�һ�/U��'���A�c��eu;��\Bi��o���O��l��iGE˷YO�u����z�����{�����U�O�{ɽ���U�+n������1Ju��+�y	tj\��5�4��%(��^Hi]�#�[�nҺ-VR�Ӱ�ϡJ���HF�Þ;0<�%�A���K>}Z���K+mF��.Rv���!;\\��gK��<a.w4�<y�/m�"�`�+���-���"��l��dq�[|�8�'�H���n 噏{�L��\�}��V�^Q��j�)V��@O���yυ�'e��r�k��/��G����^�FW����.Z���:y.�\\��rw�t�XW)8�Z\�D'�Tc�e�\V�Av�������n
�=�a��N����3�J���ub�l���Pc�pYZ���M��NlY�ʷз[Y��/�u�_;�Ȧ陎N�w[<*
욕�¾���'��z����r�[V-��qߜ��%�����9�t��:��E�N��7b�5)fJcg����G��s�����Ϫ!p��O��v���ݘ�ZvS�
�5��9:�ܒ�]b�^c���l�wS��`�s��Vg��!�,ě��Y#z��[VY��߇�G��9��ߎe;Ǣc5@�����r��a�Pi�2C-�v��5k����':�ג���{PK�K����O��u[�x�j.�a�e�y�<��\1´����c��f���qe*�R�2	�f
��h|1K`��^����iĵ�L�iV�K�5�ד�u+nˀb&�q)�gFk꾩����;7x�ݩ\�;r�pvJ\N�;Z=W,���%����Q8s%^ZWR�g��tS�IS�}%���yٮ�{O�����-��6s�,���Y$��Ó�9;Z��C]=��w�\ثi��Rͤ����VG.�X4�Mw!��̻|�Y�_#{n#��^6;9�Uk[��5�M�ܬ�O:ts�V�٪f7;}]
+����l���Zgu�Fs�<�\O.!�-YM��t��� �nW<KRH������s|N�q���䅤����/^�+�#V���k[V%c�z�^:EnQ<�\�A\&�Yq�+�����[��֕�)�{���˗���yE0�F�}�9W�/�j�@�-}��w���_+�ܥ����u����*�щ�+G����9��L3QxJ��$�Gcs;z��ve�n7^o���[}�}T�¨{�&:��:�t��9E�<�n�]R��!�Z3�ޕ��͆�l\:Z�C�7�6L�4N�Q]�a(֚�6x�FBD�����B�_ɆOd���^���cQ���dY��[�J���a�/���	�H֦8�$uy��y�а=�o�ɖ��]����Om9@�I���;�'R�f9΀��V�l0e{K����P���+.`�ĩ%�a7@>��{x;"��Ņ�s�F^\$'}��)k��{2�T��^���k��Dz<��E_�� 2������z���`r������̎�iFKwN±o���+�.%:�Y��r?>Y����mEb���).��w@�\�Sv�_8��tj����^�ג�JuyH�1b�(��=YS���7Ɋn֋绮�ڳs��k��9������3�v��w��QOd��cΊ��+�fsazݽ܆����vg�Y�{�@N������ޔylέ+ޭ�QLUw��ƚ��ˊ�y8C���m��_�nףVt��1�°e(�j2��{T��N�3�z�*�mI�*�K���Ӕ�o��䶫�v2�=����cLU�C��$���y5KM��ul�gr~��zu��ܼt�,��'�D���(�"ђsH�d�D�@x�Δ5�S,
���N��kR�;l�]9�%��1���:&l[�VKj 0\�rR�:R�8ԗ����\��P�p�v�<���Z%�=�M�{y�˩�vrfpV���r{μ�#��������[�w�ֺ��Ts�n�WZ�Iլ�S3Z�#�vΕh7{�O%ϞI2�U͖�k2t�Gqn>X������S�8�+	P�����QhL����ŏ��ҫ��/rL�JXr	�DBsڡ��Ы#���,�J(Wo�uJ���@�R1\`t(��p� k	��7
l��ÒO���Tu�^�x�2����Bi�iCH�������s�[.��$r���5�i�ݡ���vX#3:n݃��_2�;9���5�Y[�>�k�Q�rGxO`�"��^'���;F�s����|�W[H�4'+a�ҺC'��<�w�Z���|/�{���P�?vMn��$(�g\tk�ݻܜ�]�&c��d9�w)!)�u�]�kY��E�z�j}�X:E��\F�+^��Ȩ�,���Ym=��t�/������n'�ţ����K@�{8=�TK���b`���!�2�![Vj3Q:��c� �����Y�+
�.��5�(�B�]4�0SyttCzempLx�$^��3�62zy�!G�����{��ձ�v�n0�,���"�,�,�X�\X;wh�l=���6�h�D<�9K-�G�r�0����ΛG�^QHt���V�;�lk&B�h?\�t��EE�m>���,̌�7�7;\��f	��i���^�zUw|��.�&�|:�5�׼g�9��M������Z�����v��b/�����
<ͨ}��#ni�9�G�M|5�5_e�����Ú�D�37j�5�MT5鸸e�S�ض`�r�C�Z�� :p��.PU���s)?l��)�9{|.�����Z_Lvb�zBX���t��&M��q��gk5: '��8wZY�`��p+��`���[�cJ�VoG^Y��&��n(ӥW4]�����/�:�������D!rfa�*��\G2�#y"���H�H[}�;˅�B�k]lԩa��`�%oH��k�"AQm��Nslo��l�d��"�+����
m/��J4�l�tP����M,�w]pӇ��ᵗ���E�����˃+��!`�<�0v�yŋ
��N[6Фi�5}0`l�3]��k��=�<x+p�/�K�IW{VW����GEi�`���gw�T�o��K\@�����f��\6�g��i�SY�:���T=�P^!�3�������$���`��ݝ\z�`B�Cs���ˮ��v�]�F�+-��vۇ��ڎ�Q��P�6e��Q\7�K�4`�Xi��r/Vլ�ݝ{��k��'�5@	IM(RE%J�+!H�%-�E�NLC��YR4���MPP�f+�P� PSNK��HҔP�B�M%P�R�D!B%@4B՘d�E%"�H�ER4dT�KIJЅ QE#BR%#IH%R�&K��!T�Hҙ d!B�f	BQ�LH�fPҥ44)KT�dJP�`�4TW�~��fuuv�S����1�+�ޑ�+1bT��թ㪭���̕��qM�d{�Dh�w�,jN>{��^���ٙ5jU�6�Yx�·�P��o�g\C���������f{���� ]lr]}��T�AN�>wq�JU�M*{�i�ף���p���v�\����a㝣��ʃ��]z�����S�o��K���/����<zW��'+�2�Y�<%�B��	�W[�	�iW�ze��������9����{{L�$��g�]s�+f-�1\2qf8iLջ�j�ګw6y<C��imvX�����Rok�n@V?xDhz<�ΙGWb�̮�[��I]|-��g�R�e�'a8�n��6G��hs+�ՙ^e[6s����\eoT^c�g b�@���Es���y�ΚإV�'��Mᭊm�Ce��ˈ�sX�Eܺ��s�	���y�Z9Ř��7ka�Pq]��S�V�d���NJ����J������sc}TN��6Eǋ
���v����q4��"x7OS�Gd(:WZ!���M���+�/�p]�j_��y��_�t����.���GRp�a������{�#E�ј��W-;ni:��#Vz����9O����.1�1$��G����B>|�r~��'���l�N�*��KSY*/���~���e�8�y����f��������\�͖�ޫȌ�3�CA�1֤*S���w�k���
t�kyp�kr)�ۈ��P�9�͝�/��Tbvt������{kz����E�b��Y�9ۇ�f�&�oұR6��-���L�B���ԯ�8�%B��|&���Ħ�w>V�<�|3� [�i��Kiòr����0m�߹m;s�7�����]Ҹ��Y�pu�w2�"kǵa����?v�K�10��אc���UA}tm�tH�{H�Xg&��ΎK+%�������k��)V���5�T�r���m��B{�K�s��g�)�����OeB\��/��Ks�棫�቎�xT�7�����ow�."�@�;�ݯ}��{��Y�K͆�t[�����6D�[<.�[&���Ӷ�z"�A���������Е�bA}��f����x��.`ä��hZ�]e�u��s
�N��^agvG^5n�1��ؗw�QpzGfG�����N��`J�d��7Ɇ���6_Lۭ��	8�^���L�}N�Y0�@���F���'���e�����.|�q�Hv�G'�]�w��F��Dfk��7����1pߙœ�uv�X�؀�l�wS��p�NlY�V��i��<�R��p������w��Q��1MW�2��=���{�����Xkt:�Fsa���|�&1ޚk;�E�>�ȕu���d�Z��pk%⫫x����IFTf�-h�'�����zG�϶��&���:���'$>���Blz<9���g�ESg��л7�=� y��nA^}��$�z��y+���y'%7�:7/%����{�?����#�C��������t��ވ��C�>�g$�677�՗�Dh�{G�8�ԟH�����@{%�dh�ԛ���tn<��}��K�؏��r�]_C��t���?���H�!��|Ћ����+Yw�}k��=��G�A�b�~���>c�A���&�{���y��&�ܻ���GRrNεѻ�����tn^}����q�{�<�5�
h�.�fv�?r�E}�`���ֽ��s7�i��]����?Op���W����7#��17'$;�P�]�G����ܝ�}�/���;;���wf������>����u���R�X����\��w	�}t���pRxf	�?C��u�J�ǝ�r;���X��S������1�ƥ}��^e��t2'��|pYz�RǸ�c���3�}Zѓ��b���1>�6��zp��l[�	����L�W�[�U���X�@v��E-N���#Qq��O;{[R^�~�np���!�%��U;��ֺ��৲�����M�u�|w%��ܒ��/�9^���u�ֿqN�>����5nG�y�9�����A�ܼ�B�y�}/RjS����AI��9��0���c�"�����ۅ��j3"���s��_��s0=��u{�؆�7{������~t~���#�|�A��_^k�cԎ���z���߽��u'�`�R�wk~~����^zo;����~Ϸ�WR{<���;�R��S�09.���'�Z��rs�V�@z�΍I��]I�|yΑ����@��";����D�}���e[7����}���z�S���ܾ��Gr���07d�#�1?C�ҝ�c�C��Ou�HnC�5��?�<�:^G���g�1b#�zbs#!m����#{�\|;x�ps����ۿz�=C��r˩}������}���Iߘ�/�;>�rA�rOZ�B��s1C��z4DE<����9ϝ�_ћ�z�}��7/�S����~�î{�����^��FB�~�\��w�!��%Կ����j;�����C�%?F=��"$z5fD�LN�Fޡ;=��5��n$z�{�G�����1(7/�S�`�>˳����^I�����^z�:\�^���>^��x�8"��E�b=�G��쬏�}���sr��{&���A�g%rr�~���Gf�ѹy!�`y��rƹД?K��=��G�y�z\����gK��~�d���#�4x��\�\�Ck��:%|�u��Hy�����C��]�^B�������G~�r�2���wӐ~5ΐ�/�s޵���q�=�M�lI#i��H]���E?x�ݩ
O���>��������y'!��/�;�pWоA�7�y��>�Ò�2���y/��?�I=�=�]3��mx�|t����Tf�q���Z�j��Go���Q٨�"�ͻp��kY��75ɴg{�㋆)�O�e A�m�`ԃ@��Iŝ;Q�*�pk��nN��.S�oσY�AÞN/��^\;Bؙ�)-�81����Ư�w�y2^��U��VD�WpڷHʻ�g���>��?Hq��ݎ��{�w���nC�f>J{���w��wߙ�;�pR��/�r^A^?`:�pwֺwJ�>��G%��G����������0�u�К߳�.�0{�=�F=�Z�Dh��G�c}ؿ�<?s��Wp?�߷�䚏%�z����NG~`n
W��t�pR�{��w'#���<��?�=�~���|y��:�޾�����H�'�F����F��?���1y����B�!����s��=~�?Gr����W��;���G�����k�wyu��~�|��~��k��?��9��}.����^IoC��s����R�o�/$?A���!?o��s��O��"${�#dď{�D1����}�7Ϻ�}��>��kݧ��_�u��_ђ��K�p?'ئ�ܝ���������:�#�5t���Լ�&J{�G9�k���}t��pR~��s9ߝ<�?g}}����~כCpy.��aԏ��<;��w+�ΰ9.�e<3r�^{���)�w&��֡{�}��~�@�m�:CC��`��;�A���_t��?KU�ﶝ-o�Z��}��(}�N��]�I�`�P�>.��y&���A�^^Jh�˨}�A��M�rM�Z�G�C޸��8D|=���Ow���s0�!�k<��κ�\מp^��x}�{
WPy��v=A@�kޝ�Ժ���� �:���:1����MY���O��})�nC��~�]`���~�}�o^�����������o�xy#�ߺ�俤���� �_7߽�+�<�>�z���׽��u/�`�R��w��_��{��$w�j���ug��ߛ߷^�}��}ν���7�I��}/%>�\��^C��|�2��>o�)�?K����)CoΗ#!}?s�IԺ����^K�w��x�����߷���:����$�8j�ڝ�E���Gk�m�Y�M�x��ۜ�����.%g:�ɹ��yeM�����z���5&�.�sq�@7ݲ�_׽
m[#%���,ט�b�
�.W"�ୱy}��Wɤ�}"�o�0�����D3y)�����Z�ֶ��ps���/ҝ���>���N�~�ܜ�׻Ξ��'���Pn_�S��Д?C�y��/!��^��D�����x�y�D�?E�v\�����=��_������7=���}�=��=�J~�9+��u���˷��C�(Os��7/��<�:��{���$z���޵��to�k�ϱ�f��N��b=�DlϼDyr}CP�}��;��;<�������{��x���������)\��uѹy)��tɹFIg�g�����}��_}��t}�(}����x�R�~�ݮ_H��K��~��09!�>�G�����;<���^C�~��K�/p_ �7��AH�z���Z�{��o�U��O�W4g��h�=���b0z>���?k}!�u/����^����v?��{�o��~�Hy��	�GQԜ�r?y���;���_�仂��g��ԽGO�A���SϽ���O�z�}��z�Ի����������o�>��?�M��b����z]����K�~�Hx�>J����(]���_����S�f/V�(����"�X�">G� ܼ���P����w'ɟ�9//�}7η�w~���t���?���B�!�}�r;��>��~���c����[U���[��z=b �}�G(^���?K��=�Ԝ�q�����w�ܟ�uѹy}#��!�}��[�K�����v�>�9�W��{U�h�X{��.�qD�y���Lz��_��Xu�ϝ�r
GW�n]FH|���9.���Sr���O?b����G!ո^~�C��u��z�w;:�?vl�\ѫ�Bw'��^t�I�N���;����7��<:éC�����.��7.�$;=�ܺ���z}�n]������^᾿o���v�8C�N:nT���?Av�k�,��粭��U��$�Za.ݹ$�)�^��׀�'I���'�
�$;6n�b3�����B�yQ���=f���U� )u֋v�n�j�������#��}���෹'�(�)���������:��+�т=CD{߹	�B:���:JWQ�>��
�s�pd:����9��<��u��Or;��K��O����{�y����t]9��陮��#�z>�<�z��t�����y�H�|���>�2GP}��\���׽<��u/�X�ԿG�F+�y����w=������~���>����߻��z�y/��9����� ���$>��{�W u�wΝA��]C���:�y/�����ݯPP=����.�%�rj_��TЫh}���\yiq�1�`��'��w�r�S���C��~��]�!>�[��^I���y>C�)�x �_����>&����rG��ߏ;���}��ߚֻ�5R����X?�ܿ]ǝ�;��v{���.��C������y����׎�y	���d���x �_?o��g�ϧǟ��v��~����}9Q�#����t�.�`<�w���üSR��p<������ }���i�ޞI���k��y	�:翼��μ��g��o�X���]�z �cޱD}�}��{���Wp�f��s�W��Η%���X���>�GR���>�ː;���O��<��{�rG�s��r�)��.�W�{�1{�G޷1���'����;��d��	I���s��J�/��ݮ}����]C��C��䆡��:��'��{��7����x��]�;n�l���>�C�B ��/�rN��F�~������=��u/ђo|������>�R�K��}�����<u·!��!�brC�?O��ϭ�:J�e
����bR~�EG�F4E{ R�� �C�+���7&��#�_g��t�NJy�:7/%���7�@~��|��H����?v:���;�/�x�i�?�*�I$D���;gKY�2�#xwuZ��iUr����i�Ñ�o{qlY.�K�dű/��A_J[�1ݯ|ʸ{sY�Re:��9x�R�}ĥ�"!�w���L�����D�O.�u�"x}/��‷�p��Vݳ�;�u�׳���@�Y��!}���bjM��k��^AK��n^FF��GRnN��F��_g���K�؏���ܼ�w�~<�O��B=��n��V-��&k7{/yg~��9�>�ww�~Š���|�H��$�/���9/ �<�P�]�G�؎�����ߥw%��=��=x�g�#�TUmR��+�=��ߥ�<�K�C�����w	�7�i��]����O��?�γ�_���&�uw�&���g���r�2<=����}ȩ���Sb�(N�l�����!r���?tn[�����C��}�]�~�s��>�By��M�K�)<�p~����WPn<{��w+�α�!�=xՓ	�<�n����=����5�~���ލ_�{��{��:�#�5�Hj���rS�{�z�R�9�F��u'�`��R�tc�!�c��}<�zpv��;�ؾ��"D!���X����S��ܼ���{�!��ۿz?Z��_7�G�\��7�CPn<�c�~�z��s���PP>o����@�:ݷ���X�![U��n�����{�Q���~�sߘ�WQߘ���ا���u��3X��9�΍[����:5'#�u'���:GS�>o쨀=�1���>����<�f�dtk�/PP>����u9:�5��<�Gr�� 咻��1?C�ҝ�c�C��Mu�nC�5�y���}>��,{�" ���� et��Җ��U�yלP}����u��ݯQ�������%�:�亗뻩�~��p>�GRv`r����w!�#��Jb#��~{5��q������z����]I�߱2��
xo}�?K��=��W�zo�{^�!{s�CԻ���K�]��;��w���;��1#�|=�p��0z�߳@�5�]�����q~�$�^�mм{WnXS}��X2ì��F�͛o�g�b��v����o��!eY�����騦#i_Cc����v�Hv �魒�I��۪��<k����ѣfC�]���LU��Y�[�����svF���6Y���E�'������k.�<{���:���O���<��<��<��R�IA�AO��Д?K�s��y+�=3~��{+�CY����w.��`���=���g���l�����)��|�������^A��\���p��F���K�)s����r]s�(~����g�=K���������#>��=����1��N)#��u�����������!�vy�ӨC��!�w.�a|��{�9+���7/# y�t���9��LG{���d��1��;*l}���ν�_[���=]�����}���bnC�5����Gx}=��9���r�
���7{�O#�_���tr^F@��Οa俿`��|�����w�o�k��!�~�����Hz����Wr=Ǽ��}�!Or�A�u?���;���K�)~q~���
��Џ1Q*|�X������U8����v��w�~׾��_�H�?o�r�]����!����{���_���c������rMG��=�e~���07+��K�)|=��;�����w���ߺ��~�����5=���q���(����-a�]^��xj]���{�.�?C����b�!���n{���ا��_��Xu+�G�x���<��ϼ��Nw�������߿��߮�}����C��G�✗�vs}��=3}<�w�<�b�����.�>�q����p7�A��w'�{�!�;����s7��7�\��~�����~�ԯp{I�:��p:�Լ����P�]�����ܚ7�G/�=�����[��CP�~�\�I��A��<�rBu������]��_]gY�9���s��y����{�%�
JC�?K�p��C���Qܮ��r��S��ܺ���{�)�w'f����^��~tr֠|��CRn<�����~�=8Z<�h�hh颉���W��p���wִ!=�E>n�\��w#��q�'V�޴=���m<u+2.Ue��
�t�ç�M�^����e$�O]f��[��N +�nu�E��ޭ���e>"�w̽���������(�L*�ވ��i�6�cD���y�j��H������K�)<����ǣ�;�$�u#���������˨}�A��M�rM�Z�ܿ{�=��1�U韧�ͽ���,��DF�!�z����_9�{
WPy��v=A@��zyR�2_�è~��Gr�;15d.��O��})�a�C���u��x�^�`�ߒ��==�G}f:G��9��|��<���<����aJ�7ϻ^�${5�G$�]FK�X�Կw��x������$w}o�����&r�7������G+�F�=۸�W�3_m�1;��sp�+u��e��^�o+]��9��Y��CJ�\��l��	�O�qI��N/�hQ�{;�n;=��ݍ���gv��)��U����5j��qM����2݇�;5涧'3�mx;����H�=�Z�߹ԋΪzª�p&�0�f��g��{�n���a�8�ν5�d׹��yVUme5q�**2�pf���bZ�="R��wG;}¡�܈O����y�5�mxUᨉjb�T�ۻ��yD��Rt�l�T���{I��*-�ۑK7o��ּ����P+�Gu{�W��BΙ^�S�jR���<[��az4*#����giН1@���3%�6(4�o&��B�͓.�c�j��Vgx���AT�l��5��N:��V�˂���q����ht-���%S��D<Ⴄ��4��3Un�3��,rDAU'��vn��t�;&����b��gRzDV�d�e�=�Om�;@=�0v�k��j��ɨ��{��4b q[эŃR�!\��
�A���}j0�œ9��N���ݦT���w���S�v�/o�D�|Ü_(�i����Y���]�x�1({-�8Q}޺��f7y��Cv_@��V��H�~���ٻ��3�f�"�_<� �vrr�"���/c��¯ b��liص@>D��ۖ����oD��ӤoDs7�ў�5��Bu����|2{a�D-�̫�����9Pͬ�0Zj�G��>�t"�@X�8���7l]�Q+CZ�s��쮽�%�yO�j(<M�׻�>KO���b����o�v��A��]R]nb#����9;�2	+Z������[�׵��rꂃ+�ŐxʳM���t�vo>W;�-d��&ƅ��UfVś�����B��Ý�`��C����G4���<��*��-��S��s/��WA]�ĞŲ�
NMVC��?u�{��l���l�]�7)`M3:����;"wu�4���2SO�I����4{�q*��s�D�I)��U*�Ҿ�o��$�oh�*b�+��\��{P=�f��*<���lۄ�a�0p���N�:m�7���d���j�{cv5u��)�.��e���d�&3�6�^0��K[u�A����y��,��=YA����:�A��v�����4꽤)�ʜy��{zcX�i&`�-]�}�t����L��{{��Q^�7��#!�I5�UA�\N:�����C�� Q�,��t�D��0o��B�<�����1>�!��k'$H��/��n�֊�<(�tsS`R�|���$9X�M}4���k^�Ch�X��@�U����Ue�y�΅c��8Ýz��n�Q�6�L�*���\�ӡ���j����#׭��󗷅��������oa� �k) ���u���T����{!�+]L�xi����E`���m'}�fs!����s�9�D�5�E�Eл��]Z*���Jf�圁��-gǹu�#�15��+��4���3Yx`���v:Sm�ϱ�*����u��<+c��M>G��w��H�+̘[����0bw�5��L���ֹ�]��2�����)��Ӻ�p��f.�%AHFD@��(��a�U�B��y�����C�`��=e���/oL]�n�N�b�-s-� �k�2���5�Ǣ��{R�yuq�,�ع�Rۊ���Df�͔�Ξ�J:7)U�w�X!��OE���N�'\9�v�������zw�^��ގ��k]*���iZz�rJL���
������E�i*��)
����"Z���)�
��h(2 �q��0�230������*�p�rc1)"��Z")
ZJ
�J�����"���j�%�i��h)J*j��� ���0��"2
2l�r��0�����##"�J�C!ȧ3"����a���ij��"�i� ��*����b(�
B���a**Jd� ����J(L��h�����
H�����&�
��(�*��'3 �"J�*j"�����3�%���r�WG��g�����N��i闏�ۏ���8iJ�;`*�=��u,M�ݚN��V�����U�y5W����sc�k슈�lTg1�Tkv��kr)��U�P����j8�R/l>��h�c�+�D�b� ���嫂w�zjo2�l6j�ǋy�|�!WZ*���j	�R�)p�j�1%o_x'�Շ���*qeo.�+��*�nˤPQAvW��Q.x.��/�B�[Q�u=��c��r\�>��.��0�LChtP}�9g��զ�lu"`��^��[��,�����Z�����uz1P���g�A]�9��y�sEO�5i�պ�:-̨�o�e%Ϝ�n[��N�du��,�p�%�à3f�d^���^�S�W�o6��_���ۮ�t������ӍL�r�Yx��G����E�MD���������\��q^Hv�����b�|r>�zE~���:���K��sY��b�^c�����
��K�����۫�b�U�s�,Qҫe@�X�ʩ��Q���o/@��/���ݎ��(6��u	�͚��6Y��\�$-�F����1;fj&ά����+�w�R�c�3��hXY&R��SuH��k;0N�&{;�F��K]�z�-�{�>��ꠟ�)މ���+��s��Ӆb����+�
����_�$2'6�}0�̝�w$㼒�\����;3Աx���V�xY{~��.��/Z�6�u=��+����:������Jw��y[�=ڍyƼ�4�G1���y�yU��2����ONJ��j*2Ԯu�ͅ��z<�w�~���'����]j���+�s��QQx��ZyU�-ookL��ܥ�2�ꊧ����~��MgN�F���}J�qW�
�s���dD�B�Y��9a�Ԫ�.Y�)�ە���+F��u��I��3�bޖ9S���=�6���a�W��>X�K�P�
*ܯʥ�U^�iT�nm�X�=��N�S�V+ŗ�LB�٨I�>�����a��}�v�^m���'�B`�dQ����)�;E;���cR�zT���]�>Ҫч�wFME�Z��P�ʝX��G֬��q�V�����-�e׍6�g\T�aՈ%*�\lD����n��8���lgff�$Wf�2�oXBg4�������P4i�yߺ�v�����+E����vqˆצ�]oMHei���F꯫��G��<4��j�����j�+^PP���zs>��zb���5nOWK���q/��ba[<(�ʃf)�>�)��93Py���z��9״׋���r�
��︛� ˸���Q^E�j1 �*��Yy���=
����ry��4(��l��A}�Q+��X�7F6�E�.O��;�]��\L��i*p�,��0�Ӹ��[��:�
�ͣ�b@�Y��I��O��<J����]����(��Sv�\s��wE��̮�Ӣ:r��Z_S�o����/EN��E��ONs�7Ɋ��h�s��b��Վn���̋�Z��k��ߔg8b�z1�+-.sẅ́FOX��ƴ+mH[�R�Y�ٮ:�*#l�E��^xk���J���qY�1ҽ��Ņ��i���5���ZL�w��N�����.���
��8��/����(��߸kL�T1�7��,TwHn�pې�t�����-�t�m��0��5�U�vo�If�t�o�߯�����:��s�G�~nEp�#1�OaX6�o�c�qo����1�u�V��A�Iw��pn�(�F�ӝ�	3XR��W:�(�wu�#������;�[�C8}���^��4�TS}�]�BX�oٳ�N���2�5ʃ�wu�s����y��/[i���Me�г�z˷������l�}�ѝy����N:�*��|��bR���4�\>�q�s2Z���#nM���֞v�OJ
*��< ������iwqsv�͵�2��ǩj�QWW��&i�Ъщ��QC�h�� �w��Y�ގ�Q�b~��7�W;��N�gMڮ�̊UP�K��h��l��isT�����0����r�هoXO[su��T)�t��� ��g>s}�j!�1��x@�w�w=\�ef�+�J�B^l&'b�{P���V�z�b�-�k�p�#���ώ��l�;[�e�Bp�*��n��Q�Tʛ��}���˄YWo}T<�ηWiIױ�b�@��⡰�}*�Kb���F1������1/�S�wh#j�����κ71�FFjKM�u��j�턴m�]����,�{��:�W�׽P�]���	��۞�(�D��i���3�i�l=�D��h�3�ғ�3�G��L[�W�-��-�_������G���̇�c1��^�V-��E��ʺƶ�]���bQ��&2� F�p��y	�ݶ�r��Xz��^�3j�˕sYM\Fl��0
����c)-Y�.����ou-�Ru�W���zM�yB�׉?���Y/s��Tpo�_t�f�=�����>i�s�έsb�-��̜������◕�;Y���+�?wO#3l9�QW���g)�ʕ�o/ɦ�)�f�R~	=P���߻}�b���nZ��΂�.�t�H�R�7(@�x�{1��Kޘ�'�^'T3���2�1K['
�4���\�:EVy/Pѓ����6�o&41ߺ���w>�N�ǚ��Ohq�J�-1/:�C
P� "�����G<N�)A���G)ڬ��:J^���˗��;~�N	�Ȭ�@!^{f����48W��I�
q"MՎ������斢��/F�b�r��X��:��-����
���KDoN��y0!�o1�������|�'��-�j��[�ސ�yA���j�猻r��!g��Ӡ�]���s�>U�T�[Q�.1��� �wu�n����,�f����2;�u>°>7����>i�;X&�$��LA�y�Ke};���W�W��|����}_|;�1\#��1�;�%͓���t:<�b�S�f��⣭=���p�k�R�lb3�-_��q���yxc�M�Փ 9�O�� �g���Ѝ��9;��X���[��3p���hc�2;H��o��e/.�~�L<,PÕS�$�Su#4�|���+��xn�>u��ౣK��)�*�=��;S(1����i��S��O(T^�W)�u��ܥfC�46pV�΀�.�!���r-�x�����êE?>���9��vM-�|�4��QPk���tP�΀���\��8#�d���,vl��u�(oH�)U<�"��x��'흢�_����qQ���V�zm�'��+^u�]��iEr�G��sm����i�8�S�kf�ӡ�/g�j�FgK`�/w�@ϱ����E��}B�#�)��*4-lJQ�a����E��P/ٲ�:P})݌�}P���W����YtҡU���m��."԰�)�F��s�t`3T���P"uˁ�Δ��3���u��ֵ�%��x�Lv�K�3	���M�m�ti�b=}�^fi�Q�q7�U�q��\ǒ;N��\�۩W����s� ΀��3ٹOe�xf�]�qX�ʯ,��0���is���匕��vٷ�n�(��-=iE���Gh�?��}�W�U�h�F���F��WT`�Bޥ�S�;TS܆.�6��Z��Uh��kn�J�k%f����ϟj�[�O/�C�KS�G<�O��Z�E=�rY ��n&eC��k���YF����y<#�wA�eٰ�K]	�F�	��[�1�*��r�����R5���|w�`�e���&c��x����ۊJ�͌r�|H��J�_U.M��G�k�v::��y��p.
�4�A�\�]E���;3:���N,��%-���-��MY>/7�ܳй��!F׉��;Lq5�sNxY�0߳����R�)���t�^M�9��@ǫ�y�ʮw �=d
U��h3�}�U�r����GKX�إøk�[׏��|P�q�=9		��p�ډwv�B�4D6aYؒ�mM��P���{�K��u���R�\�Ҏ��)����������r�N��ǣ^��͟^�E@�f�ҵ�o�s�C]�۾#�[��If�icg:߀Vk��^J���Csh�9�r4�k˹�[����t�,Ӗ���1bI3�Q�S[i	�0֜ޫ��:̥��4���=D�5�{�B�{�)on��'tu�L>|�C���һhDS��`��-�m]=����3Ό�.s��9��o�Q�U���X�+:m�9���ܮ�̮����ĩ��"=�G������M`!���i�C��WY�[�B�&����t،T�P���j�>%���5x����s��4��cl�V�f�.pp������پ٠��g���8��1={NM�?p��fj��J-�©���|�\���ޥ��A�O'��
_S������G�༽�T�!i�oGSޑ�]+83�;��q�S���C���O>�Q|���r��l����{�[ͪ��8�Zm����tT{�7>�f"y]��������n��ܬ�������\dI2�4?P����y��8��&�xVx4�2�ø	�ӏ����gC�u#5up �=h�S��e�'��.zhi��ꂸ�h�X��_o/EZ}���^�"xȭ1����I�.)5V!�K%@iΉ3�O��xE��G�
yk�?��ha��k0T/����E���n����߽	ʺ�X��|r�&9T]ud2���g�d���n�	���U�C����B➻�k˃�( ����{~h �W�iWxb���ޙ&��p�V�n��	���=�����%�gV$���ذJ�-cȲ�{�C�1�k2�ٖ2������q�v9ƶ���eD��m�ˢ?V�x痣�+��x���*u����p�-�]��j�u��]n�\瓣Zv%c{�~�����<�m�-��&�����ǐ�а9��F�b=s���?	���B�g��e%­ΏO�PFi��*q�L!��¡��;5��9�N�SQ�2d�$��:Ȧ�I���{�ܩ���k>�b�I��TE�;1�����X�F�����	�g�Ý1�$=�{(�՝���P��'����x^o�������rl�v~𻏚��|�c�]�_�5��( �HP�*�m-��B"{ĹC7=T�
��B�Iy�����{�i��ȭs� �gsZ�@!��.����@R���HJ��)Ϸ��<2^R~n�&�ϒSn'I��ڻ��l�Ct:�I�F�p0Tg:d��Cw�%�9�n4�ޚ���4�������0;$�#�jk��>���D(�ɎD��R�&ږ7M,�\�I�u�e�17��U����<��@�)�����+�x*�Up���,G#�]�\:�����}���t�vj�~�.��A�f������k�2F"�*2P�<��gOf8C�s�CD�s�Į���+��hQ8wZ�4fR��P�[�J�/� ����y�~K묫P�7	}>���{�ڋ]�62Q�̅:��de.g:�QR�h��3Of�3��H�kYw@�gG�5��-m��
d�\�o �YV�ύ�jQZsaʶfo꯾���c�κ��M,���1�~���_��70B��&c]�S�¢-J&���e��,Ȼ����6���a��hc�/T�RF��Vb��J E�#��S��s� �xu(�>5�h��q�6�\�֌�\�y��_��o�by��@ ���=��������ں�%Aw=O�ݥ��a�ӳv@�v�ڥ����z�S7�:�����]J&��-�rZ��+�e�=gVZ��\L:h�W,�;6r'���·G��X�]�WK#z��{,�MM[kT�~�u!�r���;}� *<NA�O{�X�B���0���TʋC;m�چt�a�<��ɢ�t�z���&�gx�&/.�~�,,u�*��=��W�3y�m���
a�;]���������Q�1Ő������G�����~�
����~dV]�:�˜�@{x�f�hP*�ZM�s�6��4�0���ɹ(vl�0ul�v��E�î��@J�2��T��%�j��Q����E<�
5�\�,E��ɳ�����!�ۛn�*S)�z���'p����P�h���m���^�"����}�������i�n�g7�?[�|%�n��T��[�涍���-U�2�6���YZu�g�3�F>�A^L�|��P��cpVwM)��\!�mM�&��w!{Ht��ha�ϴZ`8͝����/mۇVkD�L�^����]٨���� ɣ���V�=T�CGos,�����˄��Ƥ��SMà�٬��:nɽ�Nɾ�&�`qkp%���Obr�k"wv��/�t�F�Nz�:�,�6����,#وǤV$�h�bP��w'���<�*�˰up�,���(���ζ��
���,ʽ����2��;WO4�S3�g�����G���n��X��v�n�ZU�g�g5>�c#�x�>�{7���])���bsf��/�;Z��ܐ��	�\����Q�A[�=���r�r��}C��σ��]ueo	O��ӌE��g�8����xVn�Yh^����,��[1�ah;�v�c�v����K��Qi�䶶v C2쬄��NrU��'�n��C��4\�`�qu�8�p�M2�NuL�	),KrTKO,�r�iO#zgd Wfflŗ�.<Um5�}}��NC�2S~��}�:v���Ny�Сu����a��������1&ǆ\�ŭ�a�a��E�kH"��9Y�AQ����C�o3o�`	7�&�����w���m<�h�ݒ@���Ț��|� z�UvK��gU̒*;����ǳq�ySa�:�F�4v� �*����@��N�%n�ߎ�x���6�	�ݪ�T��7�ۊ����}��1���kҙ̣�-�G}7�y)���:��2l��<2QW��S�d�W�4��	<�AJ<s"�f�Y!8)�\ޥC8=�(p�Fo]�e�w�w#�>�l��7��Ƨx&3�]�+c�@�Cr������Nw\�hj��[j`y�Ak�\���o'�����G"��-��-��9Ao<�p��y-ʺ�'@��&�%�9�uơ]xK�Kuz��90�!�ef8dB���*��l�Xt	YD�(n�z{�ۊ�eљ��h1�7���=��1ҕ�*]��5�j�N콖��gEMBC�:��vZ�����6�k7���������Q@�ݷm��Fk�<ý����4\�{A\J;�J�m�j��z���r���[S{��b�	����˶\UҔ���C�C�}0�0�)��� �vAًi��{C��E�ºf��qf�)��>8�>�Ժ���nP�����P�ʂh0���j�;� .�����{�YbC�w:/�@�����!�r���OH&(��Q e��TPԫ�����"�8��c�|<��F�J&4��}cⷖok�E՜��b�ɛǎ>����ݓb_L�Մ�S~Ɋ��j�Pb�k�K�����2 �bY�j����L��ރ�˖pE_��*D ��ID$��$�EKS�A$�QQD�AQUTEP�TIERQQU4U���E-�4UT�T�%U�dU$Q#ACU)UB�CUE@UEL�UP@�Q	EAM-SEDEEPA5CCES%6FS!IQU5TEDC��e@E3KAA1M�QUIE�UAT̳U5T�MD�AD�@UUQK1Y���QUQUQAE4TT$UDE1D3�IT�Y�MRDTQTE%$Q�RNNAPT&XE4E3X�EUTM��33U%5DFf4�LILE�KCT�FfE2U  �y��b�#�O{~������{Ru+�/�h�y��ͯ��u�E��w���4���gZ���ړ֋���z"<�˺�S�x�����z����L+���[HҜ|�<^�0`�kι 8Bڞ�Y�$�Q5��3��v�����ty^�k�<O���d\F�MU�Φ��i�i쳳u�-�[��$��!�0�ӏf��:uށB0�FSf��h(��L���Jwa{�+]�r� ��j�vڝ<R�y�O�vܰ�)�F��g:gF�1�*c�DuӁ�PG�U�{+t�CŰr��c �Q����i[�t�짹_��6�l�Q�3 �1ԞSi���r��6�z��iF����b�u���>ηֆ�����.�"�;H\���Y����[��1�Ȏ���`�2���,]t.g���xz�������5JzR8�)���|��`�^����_?�6:%[3�}j��~�yt�������c|n)S�y���\5R�T=Wˉ���R��:�E@8�9�T��s���,>��<�3/0���sk59�Ĵet�.�0��A��'I�I�6h��E�|Ձ��lq��P�I��%g��'��ae�V��:"8H-.�%�*��̺R�8	mʹ�H�I[tԼ�oB��c�ǫ�����!�)�ch�M�B�]E�gvb��#��d��d��7t��ҢUm�{�س���lƛ5þ�ev��;��'_�#���Ucdb�Mn���G̱Zn�p�,,< D�u���'FMz�;Mc�@��i��}"���ɽ���_/�q���j���bhtZ�ck�.���6h���v�,vԮ�H�TaHї=��aԡp���W�.j1Ll̮,BS.NB=���;�`+��=\��fFH�q�+H�h�9%�w�2ܱ�䓚�`�0�&�&�|��|�E(
�S��x����<2�÷d��M\�Y,p�̚g����j1S A���隵vWs��-�[�~�,:�R��Ȱ�(u���X�D���7�bcj}�Ǣ���W�Ң��m�)F��$/�}!W��c��Sϗ��c���s�3W�):�I��/����ۼץ�ӭ���h�>�R���̱^���̥X7Ny>��z����R�g�Y*��f�k185����w3�\�@���5�d�Up�l�zrE��,z�]X�s�t8d�e����싖�1^f'*��"�v�	��� ��� p1���
�r��<�J�@l�=Cj'����Lt�P���t��Z�8���ͤ٭sm�ޥJ2�[G52n��b���K�t�h�����̭|�Y����K���n��,Pɑ�z�4�˺+�:ksz�ֶO8!u�ա��Nt���"Ox�W�� Ymc��t]��g	�9.hmę஝B����S�yc�f)���M":zUaE�w=��d�HLksB�S t
'��Go�]/��
�r�^��+E�F�zηr�k�]p����h�}U0#|��Q:,�����{<�C�ߎ7���L��B����k�Hz��WB^�b���nlG�d�c� y���b�ʠ#7��۫��23�s��c;<��Й�ܻ9y疅�U�L_��bc���82��	+���f�˵�B�p�hTLQӓ^���9
�F�f�4ZsCb�:����E0��5��kH�H�JF�����MD�Ph`�,���.hk,r.f�Y�Y.o΄^X���}i��h����C��t��D�u`r����»<*#�f"����b�U������� 8������U�Y&�>DJ�|xKK���/�l���=�����H3�EN�N[��%X�U.�4k��2y���{q"�ѷ�Nt���ɦ#/��F�mz�R�&�C��*0:���w!�}�c^w�ø�]�}�t7�e��
G;w��=K{SU�I���lxG�x�+�{�G�:�{Ym�1����}�|�5gzg�5�rD�����N�ue�����L��c�}P���=;�g興�{�SX��6�#��B���F������2m�R���o�س�n���f ���Nz{���T�S½{T�\a�
*2aΪ/!K�jX�=��C�cz�+y���Yy�q/_�ڈ��,����s�OW�E��x*�Uqp��Ӑ�&V��'J�⨳Y[c��)$"��j�{z,+>�V�����1�(����ԕ��Z�:7����jYGiL?k��~f�t��S��h�d�L�;��EE��Pa�-��=�ֹ��^ɾ�~���z9����B��z
ΗLjs`�Bz "�".f4�lu��Ľ�	��n3�.N��L1^x�Ey���<�>�8,�0�D��"�5����{"�����l�11�ٸ%�Xr5K眭������a���UgFhm��/^ű����k���/İ��#+�ãY�@R�|�h����z-���ߓ�S�&����ܤ�팊~ŷ0+�HDϗ�'�r*�5�خ������}<5���5X��ӑ���&��uMn��1\�SEO����3Nm�I�浺/Um���YS5��28+Q;!S[7:jj�E�;%��������
����j�O�T���i�-��gw�����V@�E�WdWSuLZl�s��W��}Y�����m���n�s����rʒb�[4��r�9M�k������U9Z>�=����kŢ��;2�sKbE8�5�.9��"����^\��x-�*��8�S|<�~ܶ��`�f�v	i5ս٪���L1�xȸ�A���V�� mf��Y�0E����Exd����n9���=�q�ɳ���^�ΥGw}=B|=3��@0<��<�=֮'�r���e{�R&O@ї��F.����$�
#N�q1\�����<K0fb������BK[���|]����!;#�Y�kB��&���{8S"/#:��VF��JB4J��S���1�~�v_��f���`H�7-���e��NdV≠�]~��27Eb\�������cT��b��m��-��F��F �2qҁq{j=4x6`��ʵ���a�J��΢ŧԴ���at��kx���̚!���.�3s�ëXw_G�
&b�2��pB�},����y;CQ���.J'z$�ʅ��\���K]m���iq�=l�g//��08�L��\!"�	�&�c1��+O��%6U���A�9��$��e'{ӹ�.����4x������*��윶E�o��×�X��-ͥot��ŗ+�5��J���:��G���N�Q���]Zēa}��e�4!��Q{�Dv>�<����z&7]�}�u<���o3cnf��:��rPu9�Ғ���徵t>���˧�{|����ME�s�{��8����Mz�J�m��q;B\2*\=eE��tyl9uZ�|�~��!z�ڿ7�/՛�ާ�E-3�����*�!�`n��T�y�^'��ՃI�Q#�o�t���;�iu��^�q�\3��4t2�i�r��s���/�y��]7[��������e����B�/���:w���wJ֍SӜ���F�ꡄ����7��8�ZYT�B���}�UK�
}u�����1�2���S�p��z�0hwRĸ�ʁY�)ki�Q}W�c�2E0ǆCr���Rd�P��x_��IUy�)L8��%eE=m�!��/{��Y�eȅt&h$X���p����)f�����#����z��L�u!��� �����6/�:^��E��:��t|�S��
�D}�Vbckټ�]�U��n����wZ� ��8���绲��p���i�%+��u*�
���X�ƶ�'��'� 3*h+����+[X�����'i���Kl�����N��D<đ���.b�Ub�W^ٚ����>8aS��oV� �2����]�T)
�r)�DG�Z��[�)����+�Rqiym6{�SϗƟ��Z~�3�R�Ux���
,H3pg'~{��ˣ�on�.0�{=J��mS�}����6Y�}���	��ם>8��Cԗ,�0��&&�a@�,3^�j3��.��:\��=ua���J:M]*�պ�uо�'����q#�ط@W �<�>Ei�c�=/�C8��\[C��1�2����H`�.U��R�{zzhi��S�U-+��q�\�]�p|f�����Z�}�T�e{�з5]{���x:����7X5#�)yp�蔽IK�-ų=	v��}օv�dg��������`S��º��'j�f��і�k���`׭EMVqq'B�}Lz������𒼠�������p�a�Z_RY�>��F�%�-�7����4Ƅ�`؆����[�,)��7�������-���gwZ�;�� qr|�8�*&(�ɨ��뜅N�SQ�3#!'P���㔼`��u��}ѳ�ti�Fuf�öU��e,���1�[x1َ��x��s0�a�
>�5v�e7���������}�Ή����R��cfU�M����}���}��c��δ��qǲ�e��o�MG#;�W[��.̩߽�z7`6�hc�'���O�8�'�|h`ꈹgf+1��܍S�k��V�Ȉ��3�W��.}h������,�#�$�p�]d�輤�R�\<%��ꯑ;g�D�tE�Wd���i^)�Ό�&% +���	�\5�l��B"V�(f�U1���GN�޵9�i&����O���~,`3��+���[6�~�@D�;ۉ֍��rs���n���}4��I�Q:"ߵ���C����x823�2}�pͣ�x�#/�#b��T���*zʺ���k���~�(T^�8�D(��BW;��R�&�ڦ;�ŭ�:����%���=�5ݬ^5�CO7:k��-��:�ʮ-s��^�g�w�(#ך�;���'s���c��tɂUC���Cl���T[AS���[%l�L��"���k���ďR�p̥��^��0�m�)f!�50QA��o�`sW��yh뇢��Ot�����[��~�Ъ��Ŕ����^��51��`!�P�|J��ADۋD�%ɀ*�sa���J��$�8��ܙ�7V��&΂;�Bn��V�T�ݔ��X>Q�u�:��+�v���C��h��
�|�t�.JeԣG��qY���R���@�U|�'���Y,�[������g$1�S?�=��v������N֓X���L1^x�E71�S����y��D�)31�f����w�Pf`a�T�'��:�������P�GY�oEp}����;�ç�>�BB��q��q���2���5���&�Z�,Z��t:<�b�/��B���s\�\�~�qQ�m�
X�B$��lL��0&��p���^J^�fV�ON�?L�:�ef�}1�z��"��Ts��c5�����cK�a������讝a��v/�=w����q�u34�$i1��x:�u�a#���o��^=����X�u6e{(v���;��}�P�O3#��b�Zo���f�T�0��`�1�}���V%�rz����gg�B
�v�ûs� ������4�;EF����S�\l,V��W�4T�Q�(p�k)��ߧ���c>�+���qQ^�T�l�:J��������^N�Y��䶆e���q�o�և�Y�:"���ס��ώ�:gV;��56Ū�'������߄��+H~��V��Ze�KG���Gut�yF�����W�E_T�0 2%�TʘC��/GP��cy�N՜��ˀr�F�w�8պK2n#��;	��u'S�t�����O|�ɭ��l���2^Y�v�;�{��{��a-�j�^�bu�r�i�lf{����)|�!P���\��@�-��9]p��fb���Bǀ�q��f���-���~�1�m�F��g:gC�V����$��Ȱ�~p����U��)A���D�a��b�{=��������sHk���α�	�����s��T�θ�'bb`hd��x�epb�},YN�z�6�5�{L$i�m7z,J-�y[�}���� h�."fXwS"8���c�׬��}t!3Ȩ|'����)�"s	Q{��h0��]�7�.�Qq �����UA\D�u����SU��`���;̭t_���o�C�+�}$D�ʩ�^jQ=ʔ4�A�����OYӣ���}�Ϣ�+9���:���u���*���*{P`D���H�2�T�y���Y3E-�]^�Þy�U͇g������i��Zmܡ����|=d
U��h1��SE�S�Ԝ�6�zT�P�}%�O`c~}��B�w#T��F�)�6���
l��� �=�����F�]�M�y�iJ�}�3IcRs�Z��ަ�qfDLTvOB+��[ ���Y�U�PE�<U�k���t4R�1���n�Y�k����!����RN��a�ם�d+��������O��n���Po�F�Y}�Mr�E�ra7�bz�G���ަQ�	��]�[�Ω�r�5^��m��V��g�d6�:�D$�'s�:�z�z�,�4����j�'��bkGU��b^���J#*R��g��x�-%f���
o;�"���P�����������v]�ׅJ	`�B�;��C�Z�%.���f�P���m�S�k5�D^{s5�{1�����-���&`:[���F��d��Q�<15�޾��
A�;�z���_sGǹnb�
7�6�UG��x��n�!-n.J����J�u�pR�:��8rԧUq|�K����QC����I�ӟm&�X�Q���H�
��p�4�&�tY�[�'N�d�ߛ��\E�u��s6�%����M�g[�d&�ïv���L���MR+�(ٌ%J�������םZ�U ܄Y�1�˧��jo+qM
d�r�Əw�8�a��e�زg�n^�DC+i�%�����i�d��;%����-���� +�8M���oF��<���(�;īF�������S;q����Nr!!1�Z/{u��q�f�f�9z����LL��:8���ӛ}���[}rbVq�ɠ;�����ӑ^j�[�z�y��A�;��5�4 aW��3�/gO��`��ǡ4*���O#'L�{��/6uQ@#LY�v���_U��{O�ɽ���'�h�W[z�B���	dkAf��,�V{/�
u{���W�`�ҹp%�s��r����Э���;8-�*��M�1��F�S+����֐��)�s:*��]��vT���|�\; |jar�CS+AΦeg�+9�o�����)�L�"��h��h`ҳ T%Ƙ�짩��y��c'$�rL9F��( ���:��Nv��|P:��!�]�=w-��A1%��1<\כ�\n�R���h�^������Q�#s9����yy.�=�_�@��׼�F���;�Jޢf7���u����U2�
c�zd+�s�@��7 x��-;�|�˩6%����E�V5&mY&roYwG2�6B��"`��K����g�K�Wqa=���Jw^jOE,��\�ȱ��)��/o_^h<��2��QT�@2M�ͨ�o}�}�9�>���ǵ��b�0p:��3��~0m�X ����^^C�h+�Q�D&��8���b�����Sٝ}��E�p���^L
bú!\���n�������e�}P�zv�B����MK��i"��m�����&�PZN����k
�dʓF)m�U�dT#^' z��" �$L�TTQ��UQ1$AUD�$QI2��S4T2LMPUU$EUPTPQ$U1QE0UALQS�1��*�H*i��H��j(��"�&�*�����������	������*"���
*��rĦ(���%�����()�f&b*"�i"��h�"j*���H�"ji*���(�&���"�I*	b�b&(!�j��*`��*&)�*�������
�"�$�*J�h�J�*Jd����(`�h)��*��*���j(i����h��*�*��bh*�������j�((��(�)����&��
*&a�!���׽zw��7vu����q�>��v!����+������e�M����n�a�;��d��ۖi�����Y�n�F%qR�o�G��b�dI�w�AO@�mn+E<:�CT��٫�NfjK�ˁ���z.�4Cݬ��a�#�����|�l�������r���Rd��7~^�D�y�t]w:�3c4���R}��}HY/��-Fп�Y6}4�0:<�p�n߆��x�y�9�u1jMM��ʻ��2�u ]��Ts�Z{��y�i�ΚB�*M���0���*T���}�7�����aV:��S1�9�#�ym6w��3ϗ���5���(��x(V�έ#g���_r{PW�)AЩ���'GT�;80s,[R�_z)VӞO���=Sq�,��ٵ�
�<�l���la.-D��tÁQPf�ډު��t��h���b=6���������]��Vn��z��g�xW��
�-���`
�� n0�(�0�*zr/r&T����Fl�Q��+aip9�*a'��qjc%"�z?:�}Č��]fU��L^�ML���h�gi�oxu\=0����^���%ن+�d�D�� �����<"���inkM�Ze��k >��=b�9��x�y7FQ]��w-���do@�ImVn�*�A�d\��/�G����gnY��]L��j~`�X�rS��g'���;9Ÿ8T�i_V��J�h���zM6�3�jɐ���m�fI�� b�UXu���}�F�ן���|���k��*^;��{Dsꩁ��W��u�LLoeC�0->>V��,��U����.
�:����y�WB��*\�\��p�[����R 1slV:���w��1g�s���*�>�W���,gd)�4Zs*!9vq����)�+A�X��+ӽ;����Y5�k��h�EЮ�x:L�cG��ʝF��7q�3#"I�[�J ��wM��J���{���ȭ�MG�(�<"ICsƆ�E�;1Q����X�:�S;`>H��⇘�wc;Y�t����o.��9RK
D�%���B&(�f����5�޾�署yyHŌ�#q x��nʸ�5�p��D�%�/6��iM,{�[�w����v[�WQA�(h�sث�Y��\3ai7��w�-�qq�Nt�h.�5�1��\��2�,����k�ez���2T\ų\\ʙ7r��ƍ�A
�c����:xv�U��-�v�P���&�����/w�f�w]HWZ��iqa��mS�m�	82b����c��ݭ~�r��[���a��E��P�7102�mBĖ�����u� \�4Uп"Z(n�g�a�TF��S��%������w_f�M��raˑ�X���9�9���ЋqvZz���R��a���#��շɱ��]q��{xP��K���ާ��|��Y�:͋�&~��4�s�ף]D�Kda�����O*���v*�s:rˌ����fv"��+NE�\;!^ދ���Y�8T�9�T�{Ƨ���$noV�d��Ȱ^U�Ɔ��Υp�Of2Kޖ!�ΊY�E��n4`�0��@А�:�VEN���]	�t���4K�
�Xu�hb�ֆ>�KF1'Xa%@�%���\��AS��l��a�UG\�2j#��=��H��7��'�MI/=�P�j�h�ѯ�n�s�ŵAb�-j��#�$.2������ʡ�+�/��b��6��܃��7fE)7���8���:�oİ�ߦ
\uѬ��Md�-�{|�kO1��\��w���&�9-kNv<+���홷��N�W{"�����e/.��ɬ'lɣG��.��'75�ڡk�=|;�@�;�"��⢹�I1Q��@����3�,w׊^�Ny����{���\F��p��SL�$'��<<1�6+�W(C��lϑ�8۲@�p_�T��m<�2����j'ie���g��Hw�8]�+�@j���G@�\wrN�7j���f2l'v+o�,8@作r�6vcף���k����^���8(�1��'�Z�<w߶��yY�l^�F���R�n��W�@`���G���lg'	"��}Lf�o��	�̎�J�|��.�!�!��]m��Y��<�5�j�8vI���[U��@)}N����	�����7�U����.#霻l�W*�Q�'��m�B�ӿO^,g�%i���|�����0f7�5�^�s�'�n��9g��y���C~��U<&�i�㡲4�sGc���� O��[�.���$cs�z!��,_�c,N�T*��S@��Ńw�E�Jjm�����Xu)݌jaᅍS];�;m�������#jb��
�1ƨ���oj��Ldtq�k ^l�����*�b�:�	��<���)�z��9�;�Au�UI�iCY��OM�~�1�A���&��㱕��	��~�� �VlBv��=�o�U��]�{��w�)�(�A,v���A�";"&WP!�#H�l^�l�����r/W%�Ӈ"�5=�T<�D�T5w(�C�D(��,v�<<�sc�U��㾋ګ���!�?�Y6V-�})ӧ0�XV�� ;p�o��GG:�˨���oh���k�=�=ؼ�E,�`��X �);l�Y�,��5:�+�ɥ�a^����.���yn�6�)I0=��=Œ�m�l�k�|�P���م
{��Aݢ����Z�͊���Sc<�sp�H�yU0(���T���A�\����pv��Z'/�x�k�ґ�U�[�G����n���wFL8>����#�VK��Ř1�G��k�ZQ��$��N�ޟ^�M1���bp�;�5M�hx@��[�����Fe�|�Rx���AK���F!(U�:k\��#��xw��
a���wTz6�58��z�'�(��vtl�e��^��r�\I�UM�Y-i��bI�j�n���F��x�E��UȿP��xw/
J�]�7�����(�a����&JCw��y�I��EN5����qI-{Q9��M�)j˹��$h�>���\"����*�?��7���kl`�<��3k͝]�~�T�Q�b9�s���\M�{s���4׋�PJ�hK�6��ɝ��[ы6'Nal�q^�a�f0VsvE�Tn�Ntw<W�{�qI�Ƃ�<s^��S]]wo�ϝ�J�^N�R�̨�ʊ�N��OS��<9�*-�b3)VӐ�W��ɸ���*��k�AF��CG\&�W���A1<��� ��Kݝ����I�J�����j���Ǻ7�g-�:s�h�-��#��z����L��o$��Nhs��su�Y0�Җ�{��Dy]K�,�c5�g	��w��ي\���|��$�z��պNj�`�OR��WPp����3�w�6]=9��c��f�	�@S��lEU�c����WC�6xW�}n��,��� ps=%i��.�.�\�ۤt_Z�u����%�G 6tmҨA��8�1��ҟ���_*�%��.
�4�|�l�KNg�ݳ���8�L'�^��BcU˳TB�D��;rg��䡚���͆�GX�m�ݻ�z��,*��|(*|� rSq�h��C빁��W���1J�\oS�K[�8nu�5��}ϙ�)j���}��ǩ�+�/]1J�!v��+ݐ�7����{���Ŏ���@|!�ʃ�D_	�^���˔3�!M1��U.��:B���%T�P��\1�BŒV�x���b2MCg��B���;5P{ӊ�F�*�V0k�:��'��Y��g#��]Gi�Y����Mq�#I>:)Z\1�,k��qU����SܭT<'V^ﻳ��e��*��l
N^�������T��+˞S(U�.���c�,�O�X��|�/Z�'��Dg)Eb-A�·76�3�`�Ʒ�>�
�g,�rc;X��9���)8��!����^�6�5㈂3]�L��7���&'z���e������Hp٬4���`�6��=i[�VC�?W�s����/D�+�\�7�|&�
d�@dI�\<�hᆀ*�D�C5q��o6Eڊ�q� �dU��1��tX*�_P"��`k6�|��[Q#"ѷLM����1��ݻ�ZԤiK%�e����0\�1��ip0g)d�ܤ8祍'H�/jnN���I��]�V`!�+�����D�f���ߨJ�8+��>8����e�K*�Iv����IVp�/ֶ�XYӢ�5�t�Y#��A�,lZ�d\d�`
��[�8�@�f�UF�:8�����7o�Di���M΍�{z.��X%Y�r.z=Bꞯx�a��*7����s�G��q��IOnq��R�N�N�DW�3U��]�\;���I���q7�*�]ӎtꪝ�\_lOY��7L:n��S�A�/:_5:�0��+��΁����,���uT��l˙�\�6��TC��Bۘ�oτ�+�̺�ks_mS��5����5a��DP,p�1��&;%�aqv{\��P�}\"vh�u��k��)��Z���s:�șB��'6�mx��9`gX�O�L0���ɴCfEYD��s֟g/�kmJ���4
ᵂ:q�i�ﰣP3��q�_v�ԡ��!������O$(A������u/8�٪��S;���tX	���	����s|��{�w���v�B��J"�"}\&דPJ�'�g�bTN�'�k/kY�&=�nڨg~�]:���"���&|��d�K�\T&��
�L���L�1n�&m�O�`]�����"�aa���r�S���q	��1Q��"n%�S���g^|ّĊ$���::�,���=}0�W��8p�(1��1p�Ȩ���-=���Ǒ`��rJ&S0�����n���^�L�{(�e�d_'���:j�A��ˁ+�U�Үe+J�s��b��/�%��Hp�ԙ<%�Ȫ}~TI_K�t]n�z��e"ڞL���7qwm<S�`j"r��+�~���z�x��u������N�f��6�me62�����_��l�����x@n���9f�=:j�X�i�As�w*P���e��Y�K�;�sNjކ�/���T#.3��1q���瑿y��^�Q���#KGnоv2s.7�\����9�diA�ꅸj��Ʃ�����ݍ�G�z���uw�/=��fR��؆��_]fVWzH���*u'�+�ko��e��u��S���:M;��6� u��H�����c^�j��v�4����B�k��[��5�\$�voE�؟�(P�p���k���L��묁�چ,�KI�:�']��
��9u�s����ʕt>����)���R��:]F��==����#G:��Yy��e���9��a8�{�Uh����j,��ȣq���K:Zq�d��u����j����1���R�ǫy���>9t���)%�Ѥ+Z]���=`��6�z�Z����\>합��Ć ��'���|&:�;�f�Ҩ�I%��UA\�u��<�zԵ���<n���$t�m�8wK����+�Ĉ�{w0*�J�~����A�R_ ���E�'�ˇ�3q����Q�<��l�1#����/mҳa�T�����Z; 8:��ڬ7���>b�Z�g �b���S���3�c��,V��yHZ��؀���n0�gr�%��\�l΂BG*f��K���t`�X��2�sC�c5����c#z�q��s=N�͚"����J�2���]>���_�bI�j�\[���s��ꇋ���l�}�#p�P(;�B��"}4�*8d7��Rd��k3����q:�z��C��kj�z��c#A\�2����`4l<ꙶ� ����q�J`nj[Տu�ϲ�'�������\N�&j�L��}c3d*��(�X؎!���'�M�fh�:�Љe�W�"4�d@�W�3����yO����S,��\v�;��4?Q{N�k����aQ�nS�]ag�i"�>�q0��KL�w��Zu��k{³u�����s�׵; �b� ��n�h<����e.��e���/>V,s���CV���Œ��$Q�)8�����/�8x� `��nȼyQ�sМ��z�$_��M�+�����<d]�7�Yz�5��I֊���p. F2��'���vpde�QmS���a�SMY]t��չ��9���^����TyNcI�'L(
=gd��؞Whir�ь��2'Y�쪧wϒ�83����Yx/������r��t�t��	ч���yv��]s�[èŰ��NB�(j9��n)T �D�%�g�� -��D��.�6b�l"on.��Ǻ���zt'���0�L[�/zr<И�r���Q*�+��I�Lw�Bw�����v%�;�L`n)b2����,��B�[呌��N��;�]��e�P"�pc��n��;�mժ)�Lk��tP�r��P��]lz��+�t����f�D1<�vz3�Y�d`��n-��+�vv:;���u�IכV֘�� yK�/Q:v�k'j��7j��՝M:�n�t�`��̜¯2�U��룼 F����t=~��|5��D5gM!��ԎG��3��]״��w��dq�Ջǹv���i��Ae�C|�gS��I'Ճސe���Vd��A|����6t[���XBީ��L�Q=�n�p� b�^<�+7�3�Uڇ_��w]׃��-�v�Ȅ�Biy_!j�71m8��+��wX3�"�tѹ�_i�,�L)�{�v'�1U��I=u%�okU��i*���JS8j�]!�붅�{��VG$��T�91eu��P�>�w;E%K�|Xg��Y��jX� k�k��'eZ/��yx�ic�L�*��C���nw�+������>7� V}΄�.t��/fR��i>�&�Å-ė=�G�
�Ml���cJ�u`]�&��4!h36��L��/��n��s	����S��v'Fo�Ҵs�z��t�l�Տ�ӞavGX���=Q�Nb��!�x%���L��N�BVټY���}��^�ʹ���H�b���Ѹ:%UĐ�r9�n�혡ݷ�Gq�E�=�j
e�c���6�>u=���GZ��-��-����jaU��)*Y�K�v-��.��e��	�1���h|ȇ)t�h�l�H:���L��[L�8�����=�d��q�~��ː,��p�d���ѻukd�.��dʚ�V���ynL�iC����so����Ws�%ݥY|�h�6����a̅4�=�F�3 �`z=�y�-\��`̣lۜ���{=d�]Q��mw`�}A��f�W�Q3a1�}�!��m���V���p9>��6滕���Y�->�B���n����O���J�G�垐��v�`�Q\v<�r�1n�C�2'����`pѢ�H)��7VO���4R��:,"��ŀE�&7|�������G�M�x%�������nT5Xk`meޔ���4;B�1�A�7uyBu��8pҝ�+��d�
��=٪E��ׯ���$��e,��5j]B�긥'�f�0�w�+�օZ�|��M�J;�؉y�T��f�{c�٥����g�]���8�+2Էs��Q�7�B7Y]��E��n�+������Ȼ��|�5��C-�Q�o#������0z�ѵҚDT�*W�ܘ�Y�	��3��=���j��.Y�T�e��I4B�k�vr�����o�٘_i�"�i�I��n�zG��n[p���.)a�q��I�����:E[�A��۝�0�j'z-�
�!�8cvb��hzZ�G��*k�\�Ƚ�r�ʃ^�/7W:��:�߫A�0�<x�ҡٱ�x�KOUŷ�fA�t�<v,��R�F��պ[	��E��I�w�1%A�g�k���������	7څ��)��J�j�	(�*������H�*(fi"	�)*����R�(�(������"�H����$����$������&�����"*"�H���)�&��������h��h*�&J��f�(�*��&�"���(�������&���
�����JbY���B	������(�(������(bj"����Jb���J���H��$(��j�**&(�����bb����(�"*��"�"��*"(b)���*�� �()*��)"h� ������*���"`�(*��("	 ����a��m��c�r��㏞dv�����xf>B����$���ڏo��J��<���'�>s���B\��b�{v������VQ;(��#Q|&z������4Ƌ��T�����^Rc�Y���"%���[�W���g��b\*�
�����i٭(=��*u���C��o{�N�ʻ��ݫ]�9��K�k�����G��4x����I�\1�,k�/U�ey�>ZƷ�Bؾ���\��~~�j��rl�ò��B9RK�J�q.xmL��qò%�T��Rr��!Y��1I�S�<)�*��@�O*���8a���s��La��qk�^�c��)8����n��,`3ԠY��PXN�����EV�����]v0%=ᢶ5�9�d��L�YUta�*/&1���`��L�{��W��[Жc���:��ǫ9`!�{yr����>���������8+��j��o���08�O�{�Z�D����@{���;��C���l��8�q�A���a�O�J����s��i�už�:��^�q����\fCj���	�����݊�8*Ǫ��9=��,��VZ��y��x��Ã��%IR=s��݉�P	���ʎ^^ح``�gl��W���[�cX;�;W�)������3����9�p,��-7�*��o;�N�2T�rRtP��d����j���k���%'��̧S��0�jp�e�k���e�Eߜ���u�	��p)�ʟ)�nJ��
�72<!�{�*~p׎??b�a�뫗�g��R�9,>n��>��	z�!�c��V/���Tִ�=��z��g.Jġ^$CF��TqS��,<qL1P�uж�9|'�N�{����[�#6���D �Y�. O�pUzLuz%�a���9���W@�]R$��U����cw���n��^�z:��45Ԙ玥pM�"�Xc^Hp��Cԫ5:S���٥ֺ�����έ���y1c"����O"�>ʘ!ğ��xk��斠��.�����'7ߝK�����G�\;�"���B�OnI���iq.P�k�N��22q�K䎓��GO�xE�b���:a��f������e6��a"b��w:��*���K���XWaq%q����c�$VNVu[��(O����K�������0eʼ�kC�~���]ۇ'��^�%23Pk����M��M�r�7�&b�EA��v� ��zF�~?AFÍ�ߓek��s:p��(⫝`u��!
��ce!�ȝ*��V�n�=|�'s�h�\$Z������ŝ�h�-��B�޾AQʟ0ې�)1j�ZP��U�Dr-b�G\h�v�6�As��өTn�O,�౸{��o��d{�n��9r!�
�٥r����7鞖=u��Y��t�/l��BO�˞�%:>� =�^\���Y��1����Əb��μ����{�3��5c+��.}�r/H}8s"/3��b�����k���~{4m�׎�ol���Iyd������3m�6v��)��.3e�.6Pu��̈j�鋌j���s����
f;o�6on&ߝƑS�^����S�U8҃7H:�N�\Ŏ�j��طL.u6�a���}w��4���~�\�q�MX�t�=Y����9(1��b�t�̘[&�f%�/X5��X�,q�Ƴ/%�r賹2�i�L�^u2�C�
7�X����El��}��uؑ��j-|'����pu�<�f������fet���D�u��;��j��n={���nK�K�슸WO�؆9T���Dsک���%@��?eg_�^4v�l�2i��+���.��GU0�!�#*���/b�+2�����ѡJ�qzMa�m�b�hpʚV�#&�'��u�-��ݡcCt��{i8݋k�QC��k_�9��Qk�1q]q��7�}�aZ������G���}�ቋ/;��{3�Jf����M���jS�!a=p�5��F�;�P���:�yK�S0��8�3
�/l��q:���LK
���_N��׷�Hgd#Lp�2�i��yH]�VX^:�Ġ���V������X@���R�#��L���ıQjN�gE�'����7U�	����Ix�S��8�n4c���.٢*f;Ė#�::��,��xL^�1��=u$��;!;r�vR�Z�;���n��Æ���^�[D�iDT���Z<�L�Ɩ7�Wy!d�}��[�p�=����I�ؘ-uB�Pܔt��#MByw"��߸���O�.&��ri�re`w�Z�
��;&��b��[�Db� �n�h9�F�w���Κ��2�Uh����Ҕ��]O;7��t]�)�͚
/g�́��9�"�Tn���Gs�q"�8�0�3�a>mQ-lw\�S���F3g}5D�eR��eGFO^��gs,�mS��=ױ*c$���+��P�/ܺ�_-SqX��S84�����Et^���q>�O*�Kq{�ж��p�UmV�>�H�=����5����̬�����<+�eN@��` ��N� f�d7s/g��tf�-���҇����C���l9�難&^���]k�,;�#��SH`kU�{�'�+�l��:/�����]���V�k:*�/���5яw>��M7��O3g&�����`��\s�RR���>��r�V�ݱY�p>k����;Sӑ��P�s�:6�T!P��IZvT����t�#����xr�j�*�3d��e�aa�,}�����1oD��Ȇ�ƫ�va��2�P,��d�S�t�7�"��>�:1�*UN��y(%�\(t+|�2���k�7�9W����GNg���.7��v�U��r�bcz礱��+��C�[�����t�(�H[Q����p<�o�!���!`?����mѥ[��hU����r�vB�cE��82TX��d]T�'u�i�=-�gǏY�^�[�| -�kI�%­��x:�U�X8<�,�g�8�49�!�^o4��;��ƋN]��wP����7��x0G�/%���P�W)�S�[�!�9����9Գ�WZ��eK��#T�\' F����鸗wp�ʒX�"V����.���ES��nQ��iB�ab���x�������O*���p��65)e��@�5z���i�B�����(X�0�^NYxX�se@#3��J񃰙�`S����=ŝ0�0
ٯ<ɻ�Kz���)��Ĝ�2"��f�3���[J���k��.�4{L�ܖp��ѓt�t�*�F�s�=pDv3{�`]�\:��l$�i�*�p�_K�xS�x2wi�y��Q��=���lS�XU;z��!����%:i�z�M�_��QW
a�=|���#/j����[;�.
�g*d�3wK���4��Vk3x�l�׫i%=Y�A��ys��3��ᛪ�^�U��V�2�^�Ty$�0��`u*�|��'�5mS�b����E��3P��5���2��"��Nub��x���H��,:���3˝�9a2��\;=
��\y�#E�A��v�ɤ�W��=
<��e_��2�:[&�e�<��dq��c*|�b�1�~YhE)�n4TD�-�՚װ�2�o�U����Ļ��?��Ϋ����Ô�7�҇+y]�k:�4�^r�ػP}9] "�Ĉ�j�T+���j1KvXaz.���#yKy��PS�Q�ܷUq�D!Ol��/-Jj�6H�Ӭ��=e�zX{OXZ�ĀT#�k�^���U�����7\z%������pI��*�y]���Női%��k��5�=��	t�����t[��%���	�T+}�0)c�����v ����l���{�`FBx���k�b�(_%��X� �F����+kj-*kX��J=��GF�ϵ{��2�XGK��
9f��o�m���Z����t�D��z|8^34���bݶ�om0��&��0�Ŷi`���2s�`�q��Joo]�9����/ڰ�`���,gr.�vAa���X�j&B{rLWc4�9Gb��qn'�l�Řl*���'I�^xf1�I|a��f���3�qA��uB�x�E[��ճm�d��T��J�g�mq����c𗈊_T��3Q�m�Hp58��T3wGӁ�_t��x�d��١�"(���'�HC�'Y��Rd��O$�K�tz��s�3�v�	����f����	X+��^
�_�g�q<U��o����x�z�`n����S+R�禘��I%�I���o��3��#�F�ꑾ��GMX�����U��Y�a��X�u�G�t�٤�q��2/�8y��y��1q���s��9�E�k��4.1	�
XV{�F�p�T�Oz%�y�ց�/�lFl�E��S������w��GOy�v�Y�6��_�ȸ����!�!�SzcDuҁ�PeF��%S��t�������2	�+N����i�����Kr4[z��v����1�*=*&&�ɫ<�9(1	�7-Vr�`�8KNA��AތU��n�[Z���·�+�nr���&�=в�yς]�[Kh��yϝ��J�`���b3|�ֳ�Eн_na��j}�s���$������'��f�Ћ�J J��R�ק7����ɭ��r��)*r�%Y�h�׭�cYȧ��×E�%�ñ3(;�������V<I�D��7���/7x�ʴ����l�/��9�i��7
]��ai$���v�;:J��]aZv��z�4���mX�]3n���������+}��ܲT.P�W�U�YA
����|��0���r��̡(��;�(6w�HqO[��n��u��0 �N�ù�ڧ��6�7�QZO�qȩh��sVa�.}{q4�v#Lpa��N�
�M��]<&a�����a'��O~���L��l+�£\��ıc�!�Ƭl�V'Z��Ӓk�g[Y�֎B�X�́�ܡd:���jU3�_���_�Y�c�ٙe��&�����c䖪o�j��!�N��PԱp�*C�#I5K�2�����Q�k��=ٮNx������{ I�m��U�CrQ�y��|�]Ȱ��/�#l��⹲4�R�ǻ\�"y.�`�q��1y�L�)�u: �b� ����i�y�
}�Ȱ�����T&��C��w�k�����rG��;��)�P��`�_�;e���D
�mЬ��H�Nnp��Ik��\�J��"ûw�Vɏ9]K�p1彖�w�<4s�y��͉�1��T���,��77ޯe4b۷Y��ɯ��s�Ӣ���Pc(�sL�l5�́�����*7NBs��c Sk�-x�(}�E�-J���������4Rxk*���P. F2��'����ge�qc�h�wB���[y��N�K��٪�
��l�U<�i��� m�ϫ++fWU�����p��n��T֣�G"��j�{�*��h����ۉYx-=wC��=�Qn���� �����9�b��m.{�dn����C�
9K��	CQ��Ѳ��)�RV���48�����V3ڑk��/�r޻^��@-A\F�AW�>�y>SAy���Q.�0�D��sKwv��� �9f�
�8�8Ժ,Q;�ˈ�A,��C��Y˥{^����l:.�u�z6��^�º��}��*U�q�<%R��6\�ً��S�WB���F��9�ԗf��F]�������b�����6��D!�Pbc���S�e���4÷�������jN���5��sb������S�<l��<֓�V��2ꏯk���{+
�u��X�I� 7.�%�ֵG��Z>�'�;��Hpںb�һ]���b�xT;t�]&���ʐ��Z�c!�7��e\�
�`Q�.벣@���k������+�Yv#!)\�n�m�G�K��fv[�/3��v����2m�C�j��c����F�f�4Zr��c����dS�k�q5.xD�L����W�nƳ�!q���MM!A#�&t쩸���#T�\' F�l�;�ww�%�R%ap!Z���m�g��sj_o�U�Q����,b$��v��t�2`��2�ʸ|��PZ5,�g���jΜF�[�"V�(f�U1���y9e�cA��P��n�b��FȦ����|����e�3on$j��oeA,,܉�#(�k��GR|�z�_k��n�;P(�wz��ᛨ�u�%�W�~�b�rq�>�3����f�L�eLo�,`��t,�%��+3_P�i�沛>�i�/��҆�qkk�;����ɞ�YC�nt�t��Pw�����i���C�,0a�yU�b�o�i��Ӗ�p�Y��W��t��J���W]{�y[�CsA�܋<�6=2U�������4�s��w�R�N�N�DW�3��]B͞,��Q{ݙv��*81'H1��N
�,��,3yL:n��>��/Tעp�{�/T"�$0R�z-�Z-ǣ�,�U�x%��g����e��9�[��8��ݡ�Y�rsʎ�"��S�d0��K_H���)����0�-���#3a��nj'r;���Ư�����sހ؅��	BxxM�Cv�����:�C7͘�
w�%��X9'q⪾�WՓd�����tCG\v��Q����PԝٌNV��ΎF�G �3u8�ޭd(G�3R��y#F�V�E�wJ`�Õ��K�^Z��ml�!�[6niy��ZfǓ��]d��XX|ꛄ���N��W�1�_w:PN�}��ۊ�S���$P�>��c�_��Ǜ ۣ:�o]��-����"��7��R��ϲK��Qr�m�1��oo�i�Q �����=ׁ_]��gb��ޕ�!(#�OP�ҭce���"�ն<~����gX#C�gD�A{9�����e�W�6���V��!�EJ�v���h��xf=yw[k�u�9����W�mR��S,8NQ������ų	xwX���y����2�M�l�]��2j��qV�D���Tb�nnq6���A��xS��Ɔ������]�{�Κ6H���A��ްym�"���)G
���C�mM���k������ܯ��nn����vښ�dVf�ѵbnl����A]������eƮЪ���P_]3j2={�+�r��X��֖ŷ15�n��s�K�w��=l��A`�73w-竆L��0Ͼ���/τ�ZV`*q��&w���b;L��͛��J��8����$ε�����Sf��Z��O�b�-�c�Q9�N�)܁�1QMJ���u��U8��á���F����&��GFO�V�����u���[��G�iկ�'}t�[׽}g6��F_p���$ܖW�G���O�.Pr�X8*Y},�X�P�[P��C@�2j�oN{��N;�1{�ڰ�ia�S6��/78o�}n{���1�}s֞��we7)�'(�jɓw��C��s|���,�ZE�,���O�{c���dn�i�0& hX���r����CO��m�y2f9�A�ъ)DD�0�VZ�%�j�$m��'�j��,�LT�+� �6��L;�M�wn�D�:~q��F%݇�G�����c���
��.q��e�B,E��|�tg,ZM�>�}GF{��nz��<6�{� "ѐE3����n�t?��*O����t)���恹���:V%gwRVs�N��͎mp��nv7��V��yǆ�g�hx�2�"�K���v`mE
�+Fu��b�l�����a�ײ�[(\��:iRمw���"�c	�}�d��Ahq����j�Q*j���c�2�I���e6������7�ߖ��Wvr��Jj\�]�;s�Ϡ����rj�V;��b���L
�k
�ŗW\�N�T����"Z��*��|�(Z��*����(��"�P�)�i�������"�" ���
�������V�2r)�*�������!�)**bY��
�����bJ) �

B�iJ����������*bJ�hJih���(�%��)�����&�jk11����R��`�(Z��hH��&�$(��f))"!ȪB���(i����)�����hi(��H���X�)�
ih���)�$fbd���������(h"Ji�"�J�C$��b
T���"�6,�m:����Gv�)��6&�;�%�.	;/`Ǐ'nd��JQj��+fgfv������'1۽��U�D��3�}�%�௼�
P,�#*	��:��\MF)a�m0�y��&����P�)b#��8���s����EcTB��1�@c@�=&8��8J��T)t:�U3�\��w��<+3j��}\"����#_
B���������}��
F��b�dmbxU%1X��c1Nz\���:-��ɋNzͧ�P�϶�B�R7�Õ.�Tk���w��u�Ct�G����T���E��,:=��Nn*�=�&�ۀ��-Syy+�L<�*��.+�І\�����V`a��9%ߺa��Fi���~(1��X9ܶ�pV,z��l��]giq�)��c𗈊�l%u�=��ǨzH��)Q�`��#��X�}���΀��d a�=�q%͜�g���d�s"�~TI�}a�uw�%�r��55�������. ;(i�s���',�+�~5�q<UZ:��~*�y����6e�K����I��~�8"s�T��V�l�:OD#�EF��+�����𿏕���';�,뚙X���Ppك!ؘ,��j���-b�4r��N�iqrK�^�ᙉIō��=45V�)�Em׽�Hy��x�E��J^��O����Ӵ�/�{FĘ�Vc%���d4�� 1xUp
K0�G���0��|l��V��9��;�bRj���/�E���ȋȌ�n�^^2�d�k����ɣn��q��'�������+��i��_�S�3e�/eS��T=1~Ʃ���s��ob{-owy�֨����~�6�+Ǧ0�p"�uҁy҃7���J�e��u!M�p˪��Ɯ͖�)���ڏ;T���.07�jƓ�u�L��Q105M�E�� ���La�}�s=tWj[êl8���N.���f^K��gre��s2��DvD��]-��˙��EWk�X�7gFq~x��XL�7�����pu�<�fԺ!ł��IA�c��cy�Bbכ������DU���h����WO���r�|H��{w0+��%@�ý�!�w�p��T�'���]O��OYޙA�9�bEz���e����ƅs���C)r���$�x-�pB�[��^D���9��{9���׷�Hg!,h�X�5Ĉt�ў�1c���=�c�6��y�#�qʨ\q��"p��Ѣ�e���s���(?v��Ѹ���+Yf�/�]�->J����4�b��g{V<�,��K���=��D���ĩeҮg*U�
gX����|h)���,�yҮ���+����,�i���qw|�G�1��xI�uye+�e��p�/�G0b�ٻs�77U*˞�����F͉w`0E�x�و�n5᮪�J�V�uf?9������v2�<[ݐ�f�B5�5N�!�jWy���=���'Ҵ�*P�9qS���W=�U4��(-�W^�5/T��rI�f��5	T8����F����)�����$Ya8�C��B���W.�^�c:�A��(�c�����S ECwKA�r4�kθ��2�N�<�^�����4hF@�/�N�,]�-͚
/g�3ќݑq�*7H����C��l�F�#Lt�/���MK~��n�����9�g5C^(�p��[*+'���vp�k�v���ѕwaއ'�! [�t�U����6Y���kJ�;��+K��T�ꮠ���JJ����M;�U��՞6OmR�-9��c�"ݱ�Yx.!=wC��=.P5n��4٪�	e�6N���
��i���r�ʞ���P�rgF�*�)MҒ��J�^�q��J{�y�C�P
��2EF)���

���C�a�z%�N4&5F���������W��i�梱q�<�AA�=ާ�DoS���]ZL��S�	2�\�r&ݮ�ͮ6��(�Ho�5��Oz�����Ҳ$[�d�U�Wo'�Hh��md���m=Ժ��5-�^�U{Öj�\9�ӳ���_�����G��k�K*�ڻ�XR'���<Ժ(\K�Mc�#0��m�q
�,��@�jjG=������JӐm$����w0"�X�����]E�K���C�[���������}U���fW範�P��d,��W�F�o��y]�Fo�4=�j%x�����3���f��Tp�}O�:b�����l�6y-'�V��\1T�u�<JK%jȟ�kR=��������v~�K�ѐ��sq,iyD�ĖtD�$�9��wj�M��8`��8��;1Q�vT��,u�5N��#`Rr�ܼ����T��85[�0i�o��l��e����*��K���W�U� ���Zix���(Q�˥8˄�jmmv������5��|��^[~H����si@#9� �u�������ӵiZଗ΀�ν��ihۆ�7�x���*�7\2ͳ�*�_�֎@�(���9��wt-�q/nP�X��k�;��Õ�g5B|3u&|��
���H����eX�����1�#W�̸y����8;��(zf�q}��G�'"�	]�}�z�sF���M�ӹ�*՞z_�	��>x����i�9Û:���O��W9��槪1PeLU������:6zXAԒ��Nn.]�R#��LZ5��nl�ɶ��ӳ��^�<�Q]hi�,ۉ�=�ƾ�pc0���j�=�Š��w)O*����o��L��p�YX6��4MZ�u����7u���Č��Uh5=}ҙ�Kd�l���-��)��C�O��Y�;Z�G1�OeM��3ij�?t��LLv���{X2�5��r�-K&�1K�S��qO����eẊ�싗��VK�9�V�)B��P��Dj5N�:�*���R����J+�����c�_�̥9{Ct�������=�L\�� 1�<(T��M���({�o#K��<ߛ�CQ�.J�и�}\"��
ʍ|)�멁^x�Q�XZn`�l�c-�iW<j��ap�T;�DeܲPy�x�׋�:.�<��,�O"�[�KHD�Xx�b��/����8��uv��8��:b�I�Py�}R���ox���w,EC����3���]�mN�Bɒa�n#H��(nL�ۓ��V`a�mi��⟍��V]E��ZS<��/���>�N�.�/s5Y���LY���98���
��Y�mZz����ݠ��V�lTv3۹�9�F��m�lޜ�P��kR��:�/m��Ul�����������|������e��;ږ��/k}��Yi��lp�����*��t��3KI��8]d�xH�jpL׻m�"|���6�+�g�I�����_���`J�`c��X�B��(�H��ć_�Ϭ���|+mי-�_z����ܠ�⚊�^iہa�CM�4V���ň��8ɳ� �ٳ�P��rᙉ�Iu�Q-ӅYWZ1������QPj�[&��x��#�F�ꑫ����,y0wi�o��W ]��z�r�"ے��E��Yl7�P��gS`��<w�[����V{=s=^Ay�t��X�n���bM��P���������N�cS[�]���t�b7��ۉ��\�z�dp�9�:0���sk�
�J�J�F��*����6j�K��0e�O/*88֩��L.ȧ��5cz&z�\I��A���Y69b�[NqإV�U��_h�b3�P~��-8�O��;cY�S�b���gs�,V����Ȏ3���<KK/yOo^�GiXn0�j>���S�<4C�lw'�,ڗD8���^�ɸ���4�����K��o7=��C0S�xb�i�MFYq��65S�	S��-:J�P̗�fn�+�������c*�AC�a"����e��8�[��1��P\	�IOF�N�ʹl�N�ܞ��e�N��ӹ� �۰�L^En�k�}P9��.��u�ovͼ�͍�W���s�'" ����T�ޛw/�%y��e�x���zt�I���s@U~�ˆ:;*.gҒ�P:��a���zW�p�������ɣ�ﶃ��Q�w�9\5ѥ鮍
]�i$vϕ.u�����׷�Hgb4���������L���t+4�r�]�����ng��+���.;�K���:4U�s��J�d;�gsR�1�7]�C���ڇW`0�#f;�c��B��Gk��N�W{�u�2�g(�R�q�q�c�f��P��F��L�v:�4W���.�I/�"(`Cl�z [1}�v;�+�8�o�����Z�D�� /���1л�K���"p����u�l��9�
�tW.t����z}ys\�Re�gc�:� w0T7t�darWw&��rJǘ�v*ݘ�̇�&��X���g�e�c�Tl�ty�0Tg7dlU��el����W��~~躓����VY���X{���W���.�b�ǩխ��d�!E�.���Tע$�v�ĭ���P�9�^Vȓ�v���rn���z�i�EA��+ז��+���=�`~�<� ���d=�� N=|�ƆO8�$��ص������O5�VKm�$�C�������U�(��͢y
��Kgp�a���[T�nE*��r����WF:<�2g�ndWL(̨܍Q:cw��:u���<\��1)ݡ������c��1��J��i��K�{:�]�JowB��{�1��aQ��Y��7��!i���=9���o��:��|�a�ZW�����v��C��o���g� -�h�Q����@0�L=��4&5]`��������<��Em��bU�=O�Z:S^g�^\K���Uϭp�דC��)�Y�|�����/z�Nws�i��#�Ϯ�0�(�9q11�礡���̣��n����Wu�!\�9r�Bk*��Z���C�p��h
��@T+�أ[�sB�s_��*�ʘkU2��w�U�^�!��U/�����lXsQ(o��$�3����k���Z���s�j^�uS{�,��Q�t��гe�u����i˳��a��Y�=t}����ս$�l������b��2�0v\�ي�s���ac��p-�"6y9zn^]ø|d؉��٥՚�N�כ�.m�,����������Y�"J��,c��vE�%�˱R�may;X%��Wy��Ӏr'��s���H ���sT�v�5���un.��-$�&��u:�]|zr�x��&�ǖd��=���0�K�Q��v��.�+��/9��cK�0��R	ă��<�O��% 8��8��阍��#s{��1��J˪�ٯp�����/2E\%�϶l�>���d>��q�tuo19���a�7ʀ��;ۉhۇ�ɽP����*�7\2ͳ��V����s�wI��:�Zs8	^kz�UY��<�����9�g5B|3u]8�!��s*_���x�1����T��o�b٨���7"6XdյLw�[\.Ν�s&jP��,�"q��QO�֬v����`�՝��w]���=�+N[uñ^ނ�-Ƿ]Sh����~}��O/`�n���Pzɲ��P&+��"�+�(D��ۅ�e=��ʟ)��Z���3S�� Τ�TX���
�����b�uH��Jo�hNL�E�{)�M�paYw�l�eɋ���jS�=��!+T�5,sʬ1JP���# ��S���J�&�KUv@ۅ�u�/i'5}������y]��9|'�MI/=�L_�O@��@�q<��|��t�:�,��St�A2����'�^������Ԋmt�g�t�~�::ܨ�xraBɇ�>Y��xUf��#Ӈ�Ӓ��\8U�t� �˖��^��v�-���Ҟ5��A��Dʷc:�S�.{4"�GqI�m�J�A������E)�Ow��V��b��+�n��E\'\}Ɛ��S�J"�M�[��-#kv�ϾS��W�!1�;��,vl����S����ɋ�ߓȨO��~��Y.`��H�,���vT�%˖6�bX김'l�uJ�����G�ώz�Ǔl#����&_��:U����0��D�y�7/�T�VN��G���8�$��9,؞a��T�udv-��U�Ր�Xѵ.�B
l��l��C㴢��W1�^+'+	t����+�#�ˉ�|��Vd8�C`7a�t׋�A���c���!������cWf-���M�~	9:,�y^�� Քw+p,;(i�s�4Tk˹�g`w�2l킇f��+H�X�ZW�u��A�^�;E��8"}���E�Kf�`N��?(r�G���#�w��X����ݶ�Oz{N�xO�f�x��24�{U��lX��q��IF69�qҮY�m��y��{J��BtzE���SF��P76["�e^���d5P��UV����'���[4��i�ғ��c��W��z�R��1�Z����l�|�j�N]����!`a\��ݧS:ɑW� 1P�
�ʍJ�fF�
�:�5W)��aZ����qr��Nwm��|Xt�XaS�.��Y
n���[�vt��:�����F򑢱��F��}�j�� }�X{�����;铰սwG	7��44���)ِ�d2�n[%�-�pmB�,	W���=��g
ˡv�=��e����
J��Aܭ&u�u�,���3���tGȨXH�8��\�|Hѭ�]rNޚ7�[���Â�]/�J�
��[�p2��,Q�m��u(L�rN)��8ms`�nv]	zLN�.�G"����6��,��=6�u�����fU����;���Cv����g��Cpaɠ�zw�5�!돁y�n�]$��9����i�m<P�tT�&�+�	��0Eu{�@�ti ��ޛ�`�����YK.�l�+�g��$�>�s�n����H7Ocẘ���0�lhժ�+���.�����?f�m]�N꩙���)��# #��+U���x�����l�#ZS3L�}����'��TC�Ɋ��v�:�,������*�ӹ���A����"
y�fV�/����G%c1w.2�r��Ln�W��;D݉,�f`t�%:^pG��wՓ�5t7x��ω�w�nPi����m�}�^ ��oN�C�OFn5��N롺��'�͠���w\��N�g=:s��ZR{gk>�����GЍ���+��s.<��~��F�֝2��镄��{|,��@"��#*��ֺ������0#n�,=��
gro��̄s�-V�,Zv�����uk҆v�H����Ug�vwEe�|�9簯p:�Wb�-osf���YK&D�3K��yݽC@;th�����}�p��`\z:^V�0����j�5t��Y��DYvC�j}a�Y6�����pٴ:��7R���Y�G(�f��ըs����1�&��P�:nm�N,�͹�ZKN|����W�r�ٹe�s,
�-���`�:*�u�wC�,�����2�KΩ�Վ�:xa�'���FT��45��0:Cv�Rƛ��y�s{D���9��������2�a�骋W,��nʹ9��뚞Żwj��j윍����sGM8��x(n��Ϛ��+^���j6|}>�V����p5��c�i�Z<����e�(�W>u4��H�D��Q�)K�97Vc����55n�Q�lU����N�;m�aqqS��-~�g�GA�1���m,h�y�H��2��u�xW`G	��e��Y	���iu8ԥD���˫�'�8�[����������#7��wu���ˇh�7��:�Q1�DI=��]�`�mc87y�L̲�����w���k�_���)T��1
R�-!Q$JP�)M(SSPP��PPPD�$D@�!I)J��cED�K24�PTCQ-D�P� �SJ%RPECHR�HPR%U4�4H4	J4�Y��Vf �44(QBD�(�SBR4*�P��B�b�	H�J4�R%P�"�A@�ҙ&M��KJ�Y��	HSIT�!�Te��Z�b��K{� ���Y��A�n/��c����d��y�#sb� ���`��-mu�.�޼LZ!9@wM��N�z>́[��Y��рl�bɅ�8�ʍ�]EV��ی�wJ{[Vw��T`��==��L.�{����7��g���L�����x��T�-����eO>���������KS���>��N��r)�1n]0<�̈��^Q���}�[�^�ߛ�^O�;���V�)����&y��xh���pu��,�B�D8��]~E�j���u߽y��|����������<�s�R�{"���62�m�����1�Q�5
l��r�tv)��e��_��4�A�ʢ��0��;��ז��{ׂ\�"�u�\#�_��w��P�t�Z꽎�
[8�$��yJ��r�b��.}{�P�q7��.���U٧S������)�St)l�Z�G��7]���/S������:B����x�q6e����㉉��~smC����Q1�nO�=ã�t��̥���>�M�v�����3.!t�~F����#�i�!�^bD�kJ"�(��[��a����d�&_a��}z��j4�m�ypg�tϵ���Xb[G��]F���և,��I2�t��#�v>8��*o�޻�.�VJ���c���Ng��,UC��&���H{�!e�.�a-X=Mc��|k~�����M1u]G�0�N����6���q�m�D9���1�⠥0�lCrQ�o��)�T�m�O��G3ZmgV�F�#p�J�^B��;2i��s�֧`�*`�2Z熧1Nv@�WΣP��{:R���&��bĤxAV���^&i��2)uJ�J��2�]3n�OxM�ᚸYg)!���O.5�>~sm�tw���fɘB&�T��eE8��i8�6ga��Lu-��]+8#��U�^�j��[c��ܞ}���h��f+`P�� 35Q��ҡ��tT_n}���C6]=9��c�"ݱ�Yx.�t"y/`� �f�6f���yo�ۭ� X��=y��Z9SӐ�J�@l�ۥP�eLo]gu1����+˵EJ��~�SC�L�R�E�B�S,}��C�0��.Nո=1��\lV�`��q*�1Je�\x��H<���B�.Q5�r�f��179w+��uz�]�jr�vq���{Du�빁��W�\r�&9W����a����Q"���q+�vEqAWQJ�5��|:<�c![��\;����蠙��˞�.���oZv�ݡm�e����S�+5ݜ�@ͨ�]���e�R���r��z��=����'rD�K2w=���؁������ok�MY���H=}wwOf�fa�;Μ�t�[�<볮����b�J��#�-�@Vߚ 1\6٥[��]=e�OtPm�T�dѾ.Όyi���G�]��S��'K�x� /�g��b\*��:�)������1]k�^�ߎ@�ܿ.�.c9���ЙtvL<*n%�a��˝����J�&��h#I�,\)4�ڃC���n)�sp;�ˁ���)9zX�+n�l��N��д�(N#�R'D� ��^Z1��R�]��v|_!c*�����v92E��ч���( �T����@[G4Vz\����cE��y9e�4be�$^}��g6�r�C��`Z6�~�@D㽸�qhۇ��Λ�,,�,E�E�5׷��]�����[�������K��9K'��)%�7���n�_:;�pK�-�+��	�"��5�糚����ꭁq�D(��D.wq�Xd��Ct�d�{8��t�����ډD��R���D��lzM�<3��,a�0p[<��1s��#L&V���TҾ��R���Ck%ǧ����3���W<m-}/[����o%��դ*Ko	�@�ޫ:j[��D �E�����䯔�������#	D���(Ys�xr͆�K|$��ސ��O�].T��u0^M˹��R>�!TY��_><%��<�1rr��FҚC�9:��y�QN�Z��^����Pz�&�5r�Mt�@�['�Q�8�{1�k|ګ��3q��x���Ks�z�ḺN�r�2�]P�G"�=��ɬR�9,:��qV�0i\P����X���a�N�ȇ�^��5,sȪ�C�
P.	B0�S���J�'��#�ؑn̸��{1j�ј㫂U��9��y����)�b�D�*ࢺ��m�Y�h��=���_ӵ�o�J��:�
r��xEw��y�B�]L
x�Q�rf�[A0�����H��y4J�9��Aߋ�:/��LX�s�o��T+��@�>������Z�з��u!�r�0X틘MN��� �f��]�܂ã� ��D{P���1<Y�W�2�����yÀ�ߊ�v�yp�)�uk	��o����������)����q�.��:C��Q.�C�6EEkf�����U�0�{/i��DV'r�ue���n�v�[�(L�w��bC���J�/��]�E|	ے��^���)�&�\P/�{���ھ�3���b�F���P��ET���
���	����8Z�N���g���������I�:��8�7�4	n�樗s��jx=Wݻ�t��qΖ�W�u否�=;���V^��8��]D����(�YJvc�2r�p{Ǎ����+��EuT��n�;(i��`h�k˹����d�ռn�őү7=��f�[ׁZ�G�^����i��*�OCs��(`����L�m�smLv��)�0},�3���?_-�J�c��{�n���X���� D�h%�o�z$�=q�b��7V��nNѠ��N��B�MU4k��A@�f�diA�Jwc��*�Y;ɼ
2�>癑�a�R��v���{n�J�z�	dcT�*��u
Y��/:Pf�aބ,��x��Ƽ�zv��������������ol�Q�1�
�M����,wK��6N����0�@O����<�O��!;cY�{L\9tYܙb��ܽ9ke'xY�p.Q�ne�߫2z��]O@��������#q������	��1�Ҹ��Wa�k�[������д�����īa�G����+�.��Nt~�Pd9\Ã�A`�JE�HGI�j���d�\��1(;*K�L��T���uR��1!Þ2�:��3��F�R���p����Aa'����lb犬ٽ��<�@��,��t�On	�@7I U�|����&�s����b	=��7��䶏�x�Z�S_'ea���J���l��dW����Ư�ti�]���Q�t�'x�8ܶx����mf%�ݪvn ;�
��֌��t�g_��p�A�g���Wb#�*r�v�N{�{rz���,�z��5�$��p	C�@��KA�{N8�v���Ks[�z�TV��UY���w#�|p���E��0v#t��&&�C0�9���$�����S�,3%�0
z�{í��([�뇅��1�3^],G!2�l'!�N��^�X�)ʒXc���"�0'�����"��ʦ�s�2B���825�'5��Ī
�rQ�y��!T���cfLɞ{�Ԧ_���A���b��\�\#���*�?W倿��.������3q����\3Ǜ�e�#Mjθ�ol�
��.p`�����-͚
.6p5�va�$r1%:���\K�iwq�-�"��f	Ύ�sՔ��f�N}�g5j�e'\)|�N�,��'�ֽ=$��W�z����!Z���&�ڦ#eM�ñ���_�ꛊ�c�;�V����V3;��y��O'��;�΋��2Y�Y��33��.^��c�"ݱ����	�y�Y���lϭ_���!ǥpݥ�C�E��9ʲb�~�h/$o���AyYD�Cث�S����Z<|�ڛ#w��Ҝ�M�&���j�$'�75.]���tz�^!u������vp��;���0PTOi������鷎7OE�(��n(xS�K�cr�).����=��Z�&�X�x$�a�k�V�V9SӐ�J�x6th��Yn�=����\�*r���G,�y1�����E�$:�P�߰���d8�O�ށ vEV�g���T�\$&5ߥن*�%@�%q����*].%�&���PA�'8GNyVB�R��{o���2%:�H�S,B�D�9s�먡r�a�+-J��]_p}��=�˱��K��t�[�wH]�xHඌ����B�EeOG��h�Jq�K�ݺ^���6zX��4ƋmTp�����Ӧ((�W������x���+�c \Qwk\�yT!I��Шꋞ;5X{ӞT�5g���	˳ю��u�LJ0G.�&�JM�(�pp#�r�ML��h`ꈹgf*1N˘�,r.D���6֥��ۤi�d�]����r�7ʒXDge���B'�k
3�/�;v*]T�E����[��Lgf�@
J@��j�[G4Vz\��2ō���:���>p��(#��v��FfU�^��#O�sY�ܖYG9��H=���7iG�s���L�t��T�P01o�<;D�:�L�[)ok���gGgeC�Jn�U>�#;����_=�G_=	K]ҸNV�XN�ͪ��6/e&˙�خ{�wlsF뫠XҰ-�I��@D��ċkF�<FNt���ɦ#$W%�h�8��ud#OiB������1�״�+9S&��!ı��5�1^�
�s��)���1C{R���=�q�}��ެΫ�a�
+&-\��t��QmS�cֶ�\�:"k�5�"�.3]<ɾ�S/΋������Y���NO�KX< ugB������v��0�Zv)�N��[4��������X5���aa�2�����j�@�WKd�R�7��[P�^Ů�f��;a�jYGiL8֩�v߫��PzUAb�"�=)����^%�|�<J��u^�kM Q�d����ۚ�V�pA���|ΔԱ�=U��)J�Y(FQ"5s1�"g��n�bb��XHP���z��ǵ�we8;�p�еWc+�BX(\�4�
�ͭ�cqo��th��Dd�Sf�����XO9]	�E9]磬߷K�+��V`r�~1�H�5�=^ǧ�������e��1�&��;6rzPw_)���Nx�����hX�Q�:�f�i�KWG���]�"QPտU�M�Ckv$���T�|��q)��V:ui`C��G��j 5�!nt�[�lv�ʎ_gWW�[�N��'PbĎf&�Ʀࡏ*_aҶN�:�f���ӆu��C^��ni�n��j���*�UuWxS�@�}�P��C�ڥ��%R�ᮢ�95�دl�(gw�w�y�OVY��N��;������Q0���&+��D��v��UU�|�#���S7}�p���Ċqf����1˪ũ�*+[4��Ih�\U0�F^�1��5�P�wK���ovk��!Ʃ�3^���ȸF��^��V�|�����b|yk�	س�xm����Hiɟ(�v�����8<��0��A��~S(�EtT�N@vP�q��F3�0;j=���
�H}U*+�:D��2�]2�U�y;E��ӂ'5�A�T��Cs��8����T��.Z�Y׉��c���4�f��qͩBb+f�x��24�{U��u6��������p��#q��ګx�r�F��:/^�Q�x��,d�SF��h(��l��A�����j��Q�+�oG>uL^5Mt��ݞo�8_������&��JոɅ*�L*���w�\m0�%S��t������-����o\�"`b�;�|&5M�2cyC�Q�U��fxs�ͤS#����ug5��4��b�S�P���q��p��r��6g`��t�뮨�7�N���
:h��4�75�
��N�*���B0<��jg.���af��V	u�j�ѓ�`(8�tV�Z;�:���r����d��:�7���KS��	�u�;cY�S�bܺ,��uq6{�b��7=�����о$�	�ȄK�}̫6;�X��XL�7������9cP�yN�����x���4\l�!E�,-2�\=*�68��hq�E¸r�t�����x��ו�8�o;	54�[��`?7,� 2�lĠ�.UO��9����.�!o}Ϡ��i�K���+�k�'e�� ߍ
���u�<�nbPvQ,o��t�y��U)�Ԝ]����$+���͖�Ᾱf�=zƚ�|$�w �Y��<ւGi��v�j�CM��d���33�y�4z��.��F���Cd#t��&&�E��1�j�`+F�l�a�6�fMlؔ�ݹv����}�UK�,:�^�+��zq�ٙ���u�5N�!��ԱU��z␤HJ�O<�����Dߴ�*<2GG�eB���s�Y$�k��P�C��(�8�V^x�=��LY���HY��9u�^�7˟^B�+)�/2i��:F�@��V�OQd���3�CtU���/��1H���'|��%���}���SHA�3�e}�X�s:�@��i��t��5ӻ���Ps�J�5�o/#�Q_b�ۻ4���٨m����fQ�ΐkoD��"�D�b�b��-J�1�[	;w�eҐZ�f�fr�3E֔��4�η��@���[���k�����\v��c;�]��'���y7k-�)ͣ5�`�F�1��}�pݞ�kZ��/�{�l�w�7�Q8�8��ݜr�b���K��*���/���̩�Y��M�gp��J�R�S8����50�f=9��;��W=��C�̓�'�)K-ˆ�eiZ��.���p��-5���0,�6 z"���nnfî]Z)�}r���G�D��z�њ�@\���1`��� � ��՘re�I�.�v�N��>�;��\�H#�oU7\D��r؅aj���㨛�fR�+1C��H�m(skLX����ηc�>�[i��"�1���x��xMW
�zL��AY��f��-��]V��$�����w@}r�&
i����w���*�cX�F��ֳ;:��qv-��@]��L�ߎveJ}9`���lI�+Z�y�^��ܳ��`B2S�.�G��j�C@���+�D�K��ol��$4�z@:�D��Rqig �i;���h��f$n�..ޠ.�he��{X~�X��°79${W����L6�x0連$��}y��L�b�05fD]��ʝu3�v���THh���>�WE;u��<]|/kA\�q��Y��1�X��M=+sb����ؽ��D�����+�+��v��ge�H�+	��v��|lf���6�T���!�V8�,����Ep�1m]+���P{����Ր2(BB���2�c�v������L��扙�(���1\ۢ��7]��o�0�◶���h�2����q��F��_]=�1���nk�ދ�wsF�,�f����m��0����b�ڻNJ'�CJ�5Ӌ�mY�ᓺ.u7oI�v�Pْf�-[��/+��p����-j�9P����j�L.����Ϋ^V����Z�ON��}�a�A�3�{-�r�c����H@���2�+� �Z�<nN��(gЀdR�<^gN�ʡ���w�$��B��ZY�:0�8���MP���Z�]�E5�}�u��k���^>v�D	��V��:*H�0#��lJ��eg�׷JV�]|���PP���G�'d67x�zx�����!u�CY
SAPnj5Ʊ9��*�D�.㶉y��{J�>9�cH��w}�t��T{&�a¦h�mhk�H���;5 �d^o�c�J�-��!��M
�>']�kUt�5
��c�|�TW�q<�ᙹ�uW5�H{�x<@7 8:�C2��z�<��Uu��Jc�m�� 2f|�E�'�V^:�H�M-H��m�=�L��!5��m�|�����F 
V�b�
��
����F���

� �)��bZ@�B�(�(�))���
F�J
��I��(
F���*�*�F��J����"
J
R�j����(���R���"����J"22�����*%���)��P�hZrD2�2��)J�*nű4=y���H6��,Q�1+Δ^L]2��ο��S|�N�,_33��,$�A����'�5��2�rYMu�N:񫻯ѝ󰾝���X��f�.�x/���9:�"��������Xr[v��0�1p�����v�T�E�^[M��{�U<�V[򙵳�Fl��^K��P�,�k� 	;��]���Ϸ��@~�x3���QņME�LF�*��sПW�n*�S�EMvy�o!�N�G'#-Z�++6euY�e��r3<����t��E�ܷl{oҮX�V� �J_?1=~{�8*P5n��,C�@��\���T��C�(j9o<5e�3v�}�g�C�μ(�Ô�1��Z=*����EF)���

�>�tWm�tј-���ǚ��d��h;�-�1��.�1Je�\��ɞ
K���\�j1���M��K�$#|�y�%��G�5���ݾY˥F��:�]��e�P+Į�eNߎ�kH������:\ny����8���f{iL+޺襪ج�BO�����B�{~h �pۭӕ�6G{���z{z�����Bcj"�=7���4Ƌ�j��ľ���b-�.\R�v��q3�T�~O�J�4��cyq߹􋯎���p��j�ƙ�՘a�j�F �A}���;@�e'�k�0嫹<i���i��ϯj�G��ј���Cv�<�W}��Vk�{����F���KHW�|�ޠ�=�]�.�$�$��K���|u�]�O�c� ��O���=s�f�P{ӊ�F��7q�ӗg���ñ�;:����3��kǣ�r'Rn@��yB��THr˂��g��t�{U�=p���[5�M�D��%��o:_�s�:�D\G0�uQ�.d���]f/-�|)B��B��:�D�S���]u�綫55����ي�&% +�����=�[G<�D�7.P�ȭ���r�ڭ��r���P$߽a��m(Vrv��I�s�"q��H���m�@���%���(�z,gfí�'D^*�A��..2c���`��Tɞ�|4����疂��a��3Fi;~W�w$3�cfx��է:����YA�Q�)���76XdյLw�[\�]8������k��̜\4��\�\e��t0{Sʮ3!s���lx]�M�D�g-��N�E�\�o�o2�ߐ�Nʠ�3Y�,�kfy�1�[(D�uכ>����;��x��Q���c*|�b�1�~���_��7=��1̨+�&��n��@BX1�yZO��Cz��<O��mO��,;�r������M���]���T5#�둨�g�6�	YːT�Ǚ}/r��Ox���P�yo:b��4����z8A�Y��T���{,0�����n9
�u�ZɈK����9�%�}����c�X�uv-�sF�ա71�����K�9K�*��AHҁd� �D�W
����q&K��[M���;ZMF9a�m0�C��BṎE�<�&��)�b�D��6���l��nN�k�W�Pf`u��éu�n	\^e�9]]<"�:���4�<ʉ�ӊ�q���O�u:
:�`?n��D�(Ep0�Ƽ�%͓���:w1b�s�r/����M��{s4\bȨ��슃��48�KˆEK�\T/��l:~Ojy�������|�~���ڵ�`?;�"��T$��fx����;}���V`a��$�[��9��x�9I��c���p$�PcK��B�"�[2��Ih�]Su峝���Jr�;��G^�����$W�r�����(O��p+�ĭ#���ѐ�Y�q�Od�잹[L�YE�othT�F��B�eL<s��QPk����n9�5�T�L�~�`��&�P;�{�0�X��kh�~O�U�a]'���> �8�%��8V�gY}}if�B�!QQ���b�;��i�E��ֆ�UԷ���/u����]�yh�`~��6��^�}W��c�DT\x��+kg^�
��D�A�^�9��Y��5��ݞ���G)���,]����k8-\��]��ʆ�9X]����������NZ�8��2=i��=��:��yL��Ƚ�������T���Sf�C��U�1{j�K�s��#�t_�}�Yb_��bM�qu51�%���@U0�fw��^8�]x�S�F�B�ꅦ1�}��ntw7�;�s�t`3�++��L;��n�l�|L�s�\������N�.��5OOm�avV��vk�~®:̚#\�j�6[;dj��5��n��͸�ӱ103K&��2�� �@O��)�Ӟ��}�p����=�??5�>�)o��ؑ�"@%���a�L���L��#�Xo
Ec��3���<4A�#`�Wm'�E�LF�!5�e�R�I%�������T��/���8��G�m�i�Ubcė
݋�su��a��m����`cr�P(f�&%eI{<"�x��:N9]fF)%M��+���r�Y�1!�=o4]9TTpaTCڃ&:Ѯ$����%�uUT�`4������d��v}n��؍1��+M;�)M�(��y�R=��4ţ�������u��j�:X�{�*Hmř��]ȫi�I�˻���w%�>4�iD������:݅��JV�n#V:Or���"���RM�q5"%Z��m�V����M�_v�}L�a
����۠��<0^P1��hI-��{�M�H�ú
֤騍S�E�L�����<���0��:��+�;�����=GSSà��Ձ�{����7�Y��d��X�6fit�p�S�p��z�0DV�e�t�G���o�=;���l�I9+J"�ƴyԙ+���+U�D��qPj�p7I�r�;I��{G=Ұ�u�)�����$Yc����++)�/љ4�� 	��S6��*�[Z� ]��Ts�ZDs����\K���Rk�^�էrtE��.'J���>A<ĝn>[�U��
p:�)�0TFsvE�Tn���G\sՑ#^t�Rx���ou!���G˻6Q��-�������
�����ņM[T�5[ڭ���M�jy��Ƈ�s�ư��敖�/xF���V��Օ�2�W�F"��#����t�����d&&eeCu�V����H�Sw��y/a(�i�讖 �<��$-0���8gU��z����.���%>u��(�Ô�1���:��Hu|�a�()� u4�덣1E)�7eF�-�tφ`�%�E�wu`�m�_6��.�K��ۙ�/Y|�V��6p����D!���ǹ�_C����YRL\�x���6X�.u!5��*��˥�ٶ���N]�vu��CK��&j�1�bD�M�&7;:D����e�����V�i�7�xudd��Y��	�Eц5L�T �3�]K��˔IκV@WԱֶ��5ωwE�s��{~���^�9l�{Du�빁��Q+�\LLr; [����r���o/: w�ɍ��_F��{�BV�b�;�,;$p�[f���u ��I,�oPnu床���#W�c�/��.P��4Ƌ��G�����b���� лnc7p��5�nk��a <�R����j!�lT*��;5�҃ޕ.c�n�E��vz6��j�[T���.�۟��oaq��Y�}rI�?�K^Z)4�c�ōqx�|�y���eo���-��D����~s ���xK��jʒX�"V�<6���Y�(FYa�`N�	�+GWS�;���Z~�D
lJ Ts�2�<���hᇞDJ�r�܈�c+�f�1��2\3$�#ƍ�v"<��[��'�@����6��@��{q"�hۇ��2�{���T��v+�{6]-��p��a�*.2c�.�,��<4��yh#���k͖��Z�����r�e ���b�0[�1<���O�Zut|�Ua }��E�,ޮ�*-�۹x*䬬�2��<<���!�	v��4B���A���C�oo��{ffIc:Z����T5mX+Q����=R����B��HT��8�
�}����R�׬��ё��[��O�I���p/�tB����kй���l�ɶ��Ǟ�c1fтy 6Op��_���e�Z�u^�4�b�]g���FZ���	}�;M ����/��׽<�nT0�Zrۮ�KoE�xxF����ە\z�@������i�'�]��7z���.�5wr!�Ԯ3)��C�O��Y�;e]�V)���'7�f5�R��e�
h^!���k7��/�ӡ�e0麎_�}hg�	z��ƷU��+�#J��*����ԑ!�z}4ry�}�E|��u�S&�Kr#i�)��m�r/��yCTB��1׏d�eZڧT�J�a�ʠ�y�(Q�V�n��m������U�ތy��O��l*��8U���%��\����8޺�玥pM��B&+�£�j	C�g=҃��t\��h��K�z7֞�=��~�ٜA�����*`lB�R7���c�.`5��W�__�Ż�)-�7Lňi.�{�-�AkV6�����7
�<��u����Kˆ8߆��xnf���q;��5ժ�op���E�"�[�+�\�v�p�<�i�U`����6,�Q�}f_]�gB9P�7!�8��^��gʄdl�ekd������pj�ٜ:�Nd�˫Tc�&�1C�d�(�݅��d�O�9�w�^��P���{��=��'UYo?{)�f���	�"�PcK��4D�6g��-��,ES�i���hbJ
E���i"6�pL׻m3!	p{^��BǄ<�5视ᗾ�e1h:�ōNԑ�/%��
�w���ݹ��0��*7|�	�/3�7�,F�L^嚷���������z�ث+J0��,vl�2�Շѳ�\�8"}���Q�|q�5��t���=]ˤ������U��cH�����P<n�i����2/g�v�V�k��H�����w`��=�Ìx��y��m�g��,_b��Zm����������ΧK,�&���è�N�f5P���T�M3�w��dp�9�:.0����SV�(C�9��]vljc#�C����y��7�J�e�.b�y5OOl[�dS܇g�~®'����vҿ�+ܒS�i<��`���LH�Y69{�H1Q>�,�KND>���g���S��Y��9�ػ�N�Gs�,V�JjdGW�WB9���j>�<�DEhjw�k^ee�zq]H��ם*^]Px�9p��t��[	�v��=K�%��J�˕��Y���eJ�C3��s�u��8��y�LX��{�:�QTu�(�Ә2��ܲ��Q\f-v��t"�,�n�M�()>[S�T`��D4�K�mv=^�WC��m�R<G��5�\>3���@�vI.�����<�r ��W�;m��#'������lV�����_#���
�咠Yr�EK���s>�h�(=��ξZB\����t�u��U�<�H���f��t��p�?c�B��8�$��x�p�����j���Yq�/��~鍃BgŚ���c��,V��yH]����x@��u<>Z��ȩ5_ngE�r�h������-�u΍2��F��L�0��{I���܁p�ut6�P9=\ 6���XHc��C�{p�ђ�Mc�ٙ\X��#T�Zr�0�ES.�>�k���,x\j��m�PWf#����!a�sc��I3�����gs��"v�c�w����d���%#MByw"�G��`���ϊ׫V���઩IJ�Y.<w0�>��X�2����gs{`�r]g^�S��4�Hˣ���:)f'+K���ʅ��͊Әu
0�L� `�n�ys�y9���\H���S�w��^�7A��n �v+Jx��k,���9���G�r�R������\��Vv�,7�����2g(<��^AOevF833�i{u��;�vi�m�5�nx6]+�vX�(�Y��y:�{�1wr�t���s�����*Z�C�Q�a�k���l������v��G���wYZ�z��/�%�ɮ��5mS����O��a��,{���������]��+��a.z�*}0�TE�E��Gby]������&�K-B7�����g91V=�%eඵ]�l�7�V�	�� �� {�y��+L(=y\2��T�V:�Z�ݴ\G1,j8:6T��7JJӱ*hu�L�w^`s��Hwʺ�ǚ�iI���9{r�[�K!�����/zr�]�aB��I:��O���3�xw��K��u�l�ަ��!
��g���3/l֧�#!�9t�k�#�ULa��
	\r���O)�IJ��Q����p�Q�Qvw���,{��]��جwH]�xH�^[f���A�}�Fa��jq��� 1,�11��_	�}/��C9cCj��}.��[�,=	�kF^�X���n�pܭc�l�O5�ĸU��p�૮-;5��8��jb�0dh�`��J{;��<i��S���M�U{Uo��- mA�	,��%�40u�vcb1Nˑ��n捅��<��.s��#Z]�+��ʛ�rq��'�ٵ�Zv��xp�U';�|������M@u*8�2�_kY0�2��{ݱ�W�f���6C��we�2��jkǨb5�E@NZ�S��hT����PC��I�텓l�<ҭ�(�}en��9�n����;Z��rjZb2[�Q	5�2
��>=a���Th(�-� vRb�>�E��n��jON��-ΨZI�zŒ��RU������_��o"[[�����u<zw�Wv�,<��\5�e%�(ʙt�x�>:#p��7�|dA%5��V�q�j.�2`�;;ü:xhT*PYAY.�|;Z�sZ�|d!s}�K)�w��ó���B�Je��ɝ�w(3x��,�\�ԫؿ��2bu�m}�P����'�7f�Ǐ�j�5�={u) �Gb$���V��yք��v�E����ۓ,��i����ܦ��<8�Gt�*�Xք@�kHe2m��'�opt����)$D�Vr�����]����,�W����@M�5fK�=muZ'{���h���5Ї;����x5���� ;�U�3�v��]i�.�8iM|ӫT���0�.]�&�	�s����XF�j�ۢ�y���b�9�A��kÜ={���Q��c��|a��L�Sƹٚ8�65N�F�F���;y�3�Z�'u푧�:�XN	X#�gW8�B����{�Q�²5u���PG�o	y#��j؃yV���yCq��g�^1�8�oB�-�@8v�����-�����	ךьwPY�{���r�#]l��K_�q����c��s³�5���!۷Ɵ|���Mg�2��ft!.;�3q�5�Wlq�V.@�;��>hɤ$ �[��c�r6*Ғ��\(\���E:�wo��zl���Q~VE| ��'zٟU��ɻ���#����(7T��jQnd�"�<u<	�8,�E�����b����e�r��B��	wC6ღuID0Y@\גX��f�Z�J�g�B��^N�x��^̾��̑�vy���BӔ1#�G�
P��|��]�&�FK+�!�w�7�Bշ��#Y�λ�o��u�Y(B/�fֹym��9�{f�x���I���s���ҭA)��oY7\�fjYJ�vZ�Ŕ~�	vBl��&F��G�;3�]����d@�p�C#9&w����԰q{�t�ޞ����qBnCr�0���A犾��)�5�}�b���i��*^�D��[Ջ�f��a��+7jrU���04e�
p�g�Gř.T�վ�k�����ZMI������ގuJ��i��&\Wb���-j5�f�%��칦�ac�e�h�-|<w�D��Ϝ���6�S��i�H�Ԛ+�H�w]��
�ݏ.#��M��wq�d���ǋS�ЍS;}�}�ϲo_�P;{q�B8�mHIm�S��b�1Ǻ�N˹݁�߱�3)�@�$� '�$#A@��B��PR5T+�VfP�H P-H��Q(Ҵ!H4�d&H� �4Д!HR	B���J�	�R��)TPR)�d�%4��J4%+@U-R9�4��)JRSUK@�B���B�@-��eBJR�P��4�FT�Ӓ�4*d�AKM-�5IUFf%4�Hd�P4!HP%
R1PR)T PU�����dzr9��;}�G��Y�+IA�ò��EB�C{q��]�r|���!Kh�V�ݝ 4�V&S��̕�Co���\��4.��@�!9"6'/M��+�"D�mr��^Z1ϩ���S���4�-��"�W~��0�e��d
�ĠG9)<���m0���g��:������c�}ս��BdU�Եp��р��P!���	��n#��n$_�ѷ�{�ُnƛyve.T��.	Af禐�����0\�b��.
��L�{��� 	�w�ސ[��EשX�Fn^Ɂ<��&g�劋ڧ��D(��D.wq���&�x	�]*0ثW��Ye��)�ڥ��mp�:t_��t���8�(�9�t�Z�d\d�`A��ر�,ï�l=��ZY���v��L�4���YXxtV	WG��.z���*��� tG�'�D�^��]÷u-�wx��,@Oj���a�]�c��f!Z���'j$�k�u�U�ǳS��s5k�`~������a�u	� �	z��ƷU��(�i@�U�'&4��V�w\��Ĉ�e���u�ױKsi�)��َE>Ȧ��à����p �z��#n{s���T	�8�S�P�����=�eax�� �7g��%t��u�~1��g1KF�<��*�-6^���'l܋{ nHG--�PhWA��ج]��գ[�/z���}l��s�]B�쉼lΩL�%\��:��vu�����#��H��D���ֺ^{d��v���ׯz1+�^�r;�-��jו�K"�S��������`S�R�����0P��
�c|�@��ɝ~B�S�L��Q^��h�ǫ"ݵP[���Ӯ��T3��&R�ᒩR��ʚ�ly�p�rv}9��ﻯ`]��jxod"�d�n�~R�t�dD���|L^\1ϛ��F�*zI.mK��N�ރ7@���V�-���a�f���		�"�
mD�����E�?xg!^^��.In�ҌG�$���n�s��Egӕ��nOx�8���J�/�����b��_OK����z���z+|������/�Ж}g�9K����I��W�:�1��Ε��K�|,���J]��(��,+�~0`!�����ֶ��W����Y��f��3~1������d�>luw#5�K�L^�۽~P��q�#��c~��J�L��ȥ
�png�U�Q�ofe���l�W�����d��`V�~Ǭ�*�,!�o�l��a�x��X��0R��ۻ�)W�nʼ�YG7��-�+��O|ދ�Y�6�<��"fu>:t�Z�y�Kj��{|N�F�zxm	C�Z�6�g
�!<����I���s{vN��ݝ�0��δ��sN�WE�
�Ut����~yr��Ҝ1E[ϞJ�Ա,վ���l�T/�zc��4����#��VF5QNl�}Y�P�F_{������U� ��(�,3q��*]8���Vg��誷�S�1����y�!p��<�-�|3�%��Uh���*T3��T;������KS��	�t'��\Ω(Ov�d	ID�'^`�.��]w&X�73(;�������Vv0�j=�_�ĸZ
�����;���*ϫ4O���YfԺ!��,-72��|��kY���}k����t8Ob[��P�D�~��ȫwK�؆9T�$F���	O@p\��
b�Qb���y'�jXռ��,G�s�V:�ÞF$TS�z�<���8^pGW�����'i��l�:`�F��]��Lr��'EZ��eO�x���bpּ�-M�hx@��J�,��]o�|�l΂�Kgn���~��9/<�`��xXۮ1�)�#c��1�K����~Gx��v�;t�pQ5��7P���[�]�U�N��]�·�^�^�z�-5ȶXB�@;��<���ê�X�rCԴb�s����{Ju] 2��ܬ�aޮ�����rtoGFt��v�0����=<�/#p.�1�뛛�y��7b�-Jr�������4����8"a�k�1��/�q�MTE[��4��N�x�{l�2��``cѮ��O��E@����g�g:�~���{��(�&g����m^�+wb��Z+�b�F}�Oh��l�����;7͵���c9y��,���(ɍn֎q{���X2k�͇�u� o���_v��4�G/zq}�?E{-L.q��بykw<�uDs�5繦^��r6�<��e�VU�=��	��	�Ȭ��E�Py��jlW����K7Qa�cu<LwC̴��s7��)���b�K��j*�1^�RyR���TvS��̫.N�v�5���+�mĬʈO���׋�1J'S|���|��ڨ�M�ٮ��ֵ�awe�:�7�r�R6��*v��R�)p"�6t�k�Зc���Qۼ�p���[���ɵ�#�\:�����p��)g4�p�QW�p�3�'֛�K��MJ{���.�׃�щ�m�� Ŏ\�{څ�6v2�ސ�g,�gC�r��Fh}�^oqjq%���ʲ�������m��Y��1}�{3Kn&�I�B{3H�$^5ǯu #�q�v�b��
���Z��Ƌ�݊�%g��̈́���Z��v�������=G��;�;[˗n��&cӞ��Av��&�zJ����Sv:Ga��Z'B27_sv�Va�Z(TA��1�k��א��b:VW���/��eV\
�4὘��[Y}�#f��ϰ��u��.�ȕ�l)�p�N�c��7S6fZG
(�0�k-�uｾ{^�^ھ7x��
�}�Q+g�Y�ll�+�c0;��w���k\3.*b��ڂ��6o���k7����Z:�������ӎy��@�L�K����^��K��[��#���sx{LWJ��з���n����X�lf�|�Sv�_8��zcl���`+Ŭ�oxh��+��ˉw>���3%EF[������ykB�� �j�K����^�Ɉ��=���?Voj
2/��K�ݘs�'Nٽ�nurGu_��ѭ������ʧm�^�Ut����6D�U0;�r3vԶkJ���CE�9	\�Y&kR��\:�������T�Qf�]]S���s���T:�oWI��lMC�]E_6`�,�O_:Bu��頯�Zxf]���[R�X�vV}�ͺ���/=D�>�.Cr��8VӺz,8�껇ܶ�1��)�Үӽ��dl�Q�
��u�S���U7;<殚6W�u
��'���_��ՑM��J�AZ��^9�^�<�X=3��\�V:��׆{�bҔ�;�O���z-E�}j�Bk��CM�V���kX&x��T:^QMe�J�gR|��䃕Jv����mmE�؍	�j��c����+������cR�z[jn�8�qVe娽No'��r��}�S�1>V�E�Pc��W5�!ul �>u�Xc�K).�Q��[��۸��;��}T��{f2:��Q�*'����ձ���e��i�ﹴ���E��n�-��sp�<"c��_,
�җ{�X�Nb}R_�z��:?5�˄��Tr{P]ӿ#dh�M]FF\��yN��Uo��W~tyg|�8�'c�X5Qb�$���FHW﷙:W	�-
�:����ir�t�F�N|��p���x�:�GZ$<7�)�
��=\]^�.ݫ��o&���b������x��y�<.�_{�n�߭V��l�!��[n�F�r�dX,�1s>�5r�p�j�.۾��'��l�ã�C��WiK|iz�|WU�I�Q��S)��W�8��}ǧ�D�I~K;�"���«=X�^d��q���O���x	������h��kE�=�~Pj�o�֞ߔg����R�\*��N�ԯ6�.�5����N�9�N�c����v޽����&�	�^��r�֞-�H�[�S�W��g)�Uk���Z��ɳ�o_��z�O&��gx�1�
��V
�N�|���0yR�Ҟ_�O{"��ʐu;�B����R���*��o:op��A;��pbu1Q�
������pY�w������c���&�sV)c����PYpT�x�U.z�p�����뚞h�p�l�՞WMjR���������:���aE�PO*����klO'ƣ�5�Og���>-G���T��Oz�>����Kl(��}�c�u�(V�r���˿�D��M%��|��"����Bx,*���7Áޡ�]��a�Z7s��*^#�+�
�>�1����Z����K��ŗV�¤]�]�#gV]θw^����Ӹ�r�
8(�Z6��'����7\���t9q���~��f�w�!�SR����ԝByf6�Ѹ�8ͻ�F-Wq]V�9ޜuU��T�ene@n����^�n����R��|��ܮ���"hF�[�i@�XC�E
�ݓR�m�>�8�����4����]���V#�S����j���Z�lz ��v�n'K�Tw����}�&M�x/���H���F�v�%-�;�l�^�:��V�\��җ���9IJ/s4��!�5o{�����0�(����\�%;�M`�|F�\���e��ay
zNy���Ցs�b��e�a�X7�f:Ӑ���c6���Ox�<�R���\�v�+);��Q��s����C�[��uG<�&Y���fKY�S:����dcv]f�'{Vum��N��ή�6*-��D++8E7.��mI�Y�#�\rݭY�5����1J'Z���b���T��1;c�F����q緦������x���!ä��C�6[b�NU����@j�w��ևJ眻2�ĸ��A�q���p[�����C�L���E+��]Gxj/w���޷�oi9�:fK�K�ҕGp�y������ScM2\�Nվ�]ӊFz������5��������K���޵Tgu������ğ��:���ԝ�4�ޅ�i�ە�
E'��{@?mg�fzf2�V��OR1�q���}ڲ�o_@O������vZ�����Vi�ף�=���Λbl�z���U☷���{�S���.�x9옜��fq��mOqX�<{T2��],>����{�Q+S�="�
 Ji�#T�M��"^��+G�x���s\k��}{~�YIs��ⲕ���Ʃ9kZ~�ҹo�dݯf�����K��f��aO��VY�`��y�ƞo$��ݿ6��=�7��5��`�ɨ�L�2J�];��~�zc2A�U�4�S�]hˊ�alRok��;�F�u�u�Mfjk|h�s��D��)�p�7Ե��K��g��5�N)��W��LBwN��o}��7��)e�,w.�2{��԰����a�Ż3B�h,:0�lGȕC��dX��HZ�ԣ՚�-�}�o�w�5Y%m�;E}%Mץ�tD]T�8�G��c�h+��v�;���,0�r\9�܀��bG��V��g��zi;:�z�e㸞^e<x/�_7��h��q�KuY|�cc'L��gC��ǫ���޺��>�㕫}�,��G�I���޲��R�m���;�	��1C~|ۆ�4�mOZ{W�)>N�T�um��7���;�(�(N�5��v�?kHT[O�)f�y�~׽2�9t@��� �0n�^:�*��<|�x���N�kyo�c�7�q+1;�͈��z:ZA�<��Ի��O5Z_�s���ny��Uo����|{9�{��/V�so�,�z�ֲmTOGLRbb�!il$��|�����櫒볜]bK�U�tH�T
�m_���K���Wvq�)'�=��Q}8�['���{�f�f�y%c(w�X�]���/���w�_�vw���V[�p�x�w�p�R��O9��4&��Elt��;��Z�f�_����ꯗ��TA_�TA_�QpED��* ��Q�ED��* ������"�
����+�DTA]������
�+�"�
�AW�����ED��* ��Q���+���+��(+$�k>�e0�AM0
 ��d��Ho��ϖ���l)I��R����-�J�
� �I JJ���EUMj*��UFڥ(i��&����4j-���c-��L���Fm6�ZJj������5X1�޳���l�w������&f�*�լ��ڵ�f��RR�L�[-��4��YeQN�;CPe�klҳ[,�[[2kl������j�V��kLU3kmJ��������-mi[iVcVlZT�SElEjգR�ȳm�̶��VfmmE�٪��ɦ�e�� j��Q��r��� 	�5r��
5��9
�tc��ҀH�5ڶ�IM7%�@PUv�e\�-�`Q�Zv��B�J�[���m��V6�2���֭� ��AI6��F�Y]�89
d]�uB�E�Xj�)��f�5���bX
hh�kp�SY�� +M#�
(P����m�Jѭd6T̆�{� l(P�@B��y��P�B�
-��(R�
B��L:  P�B��
  P�î�  B� 7z��G��^��*]�#n��ʔ -�pi]cR�n�vR�Ւ��J�Ci�� G���cmk4Z�������֨,��UH(��4� 'nl�@:�S;����N�In�5�T���]�:��T�η�����Q���(���U[4f�� u�R٦�AQ�ն�j�Ά��Ք4ւ�:Fc�m�J.�*�*��� ��nR���r�:Kb�Ӷ�Sc#FҮ�4�s�ʹZ���P�cS� k����Snծ 4)U�@J�Jm*�*j�F�QJ����J]c�p:���j�Ӛ��5���[4k���hPi��%f1XřMaK6U+4�  6{ˡ��T7vn��k�tt7\�hU-��� �� �A;� cK\� �f���t#P ��ڤ��5�VV���i&�^   �� 4�0"(X��
;� q��  6n�Pk�;p U\& k!� A�]����u�lZ���n��km�KEcm�  ⊡U�pCn�� ;��*��w*��79��N� �NΠ�$8��	� ni�6�kl5 �2�[W�  ��th��  k0ȃ�nN�J��
�⊥:6v���` �:��T���ᡡ*��M�S@��n�ҁN�S�*H� h�"�0IIT ���@`�4��~%Q@  T����J��z� &�"l�RM '�/�������4��?�����ޡ��ny�[�p�[��a���]@������x{��{޻���B�R�HH���$�B����$�@$$?�������K��"�!?����v��B9�`>����J����W:�ni��4�!�ʳV�H�e���ۡXe��r���t�AQ�iQ�-&�]��!��!!�4�n&��{�S��f���I飌X�P�M܋h�2���\�U8�_R�ZUh^~�>]�$M����3ѺFL����$$��"j,;�w.�u�P�xp�؜u
�r�����t�+�彼d<�W�b���nm���hZh#n�z���B���@�Iz��RʼB�>�1kD[�[�kF�XIU�t|QW�e�%/Z��Ð+��ɃD�!S����+7p��<˒w2�8�ma�k6Z��z����ଉ�[.\+ �Yn:�Z��!l�`h�%B'u	*��F݉t�c0�1LmF��1n9Y�M�"1��yKd!�U̬�-����	�p�]6�[��
�pV��Q(��2����GSX/�ܻ���XTgi�<9L[OSX�݃(�oM��s$��)��i��iB�ͳ�c�Tp��MW��!�����/d��.�l�e�yfe\����� k(	��Fs�e��gĬO��{i��p2˕h��z�f��ER���^ɦF
ܬԃ��R�1����,f�(�(�Nݳ���!Bຊ3b�}�)ҩ[hLJm����fjel�U��ijٖ���Dl�.�ã5�@��R�QMF�A`��|Q=�D�W[���[Gb�7l7WaBeT�E�j8�g[��ǹj�X���6(JC}�v'�7Cx38l{c�5�f,"��t�)�'4l��Nl��3(�hإ N�ܽeXm����(c7(F.i�R�Hu!e�5uP!j�H�抌�7T�V�t��ŊC���M�t�wR2)�Bٱ�w�m�mi5y���X�ňk-��d�8I���H䄜��f����� �����p��8=球麪�.�-�+LDnM�7)ػn�X�kڑk[t��*�K{�f�̄�zj6u�l����'�M���[� T6�� �ҧu6�]�݆�䰨�7@ae?�-f�ܲY�kUFbz-˃Hb5kNZm[YdRf��m�Ѩ��2��-��^d�2�w��X/i��C,J���f�:��ͶK�@���N��j�#l�>eBB�Lf*$nS��ڷ�B�,��*��$����J�I�CUI-?[3ب�yK0e)t�̠�B��DEŵ��H�>��[�F�faf8|����/#�x`�J�,!�>)k�D���X�4�����qe�K:��1^Z��+�VA��.�Qi�Y-��d��sr��n8a2�	Bh9l;Pb�n�E���0�CRm٭�E�2j�b�U�K�3TWOh*g���!�Ȗi���v��0^�%K��@�{�x�o]X���Պ��tZV��w"U%�&��7tk���R�4B� ^F���j=b��rJ!�ZhѼ&L�^�	�Hch��uH�)���jv�֕N�Ot��j�q���K/����#c����W�C�;����44�Dw����b�m�ݰO���!� ���<iVb�J��%]6��0��j�X�u��VԽzAA�f�[��
�M�Ox6�O�����Zh
j�-�w+f�^ܭ����$���b��J�j�wr�֎3�!w��T۲]��i�b�S���S5Q���E)�F�A GM�e�e��ݬ%�Y��.0�`e��4X"�A��VM��OoTz��]�JU+R�oj��b�[ɛhX0�	l������Cd"�l�vM`LK��f�&��x%�{&�[����@˥Y(�ǥ�h���ĖωyV.�Bc�.]:Uv5yH��1�a��a��dj��zMڬ�j�*�y���B��"5/ /wpP(ވ���[v�љ/Gn�|:�+�<Ĝ6��j�{D��3�w���fG�:lRyV����.m�E�X�Ղѭ�e�P.��.���],z��n��'{��w�=�N��3E�`��(�K��0��$5a��T�n�B�1�q��$�Wz�W�*�!<:(�+e]�R;��#�M����r��8p�v�ǂ��n�V����<�j�v��6��e#���E��K-��p�
k�Jg�J�V�0ٜq�D���|��f欜GA�g>�Z���9Y$J�
���[I�c.��J*���(s�YWt �|fͩ���\ <��	���en]���X+Jf�1q4qf���c�M�b�v+��a+�r|g��1LmyBd��t����c��t����K[H�Y[Q�W�j��R��bW��6`E�7�*����E�i�*�[Ch"�����P�B�5"�Jyn4H���̄
Յ��ޱ�����W?�ɵ���^��6�j�2�as�\��A�6�P9�`Ȋ�SR�e3+XlXqK�⣻
ٽ���ߞ��c��m�ζ�� �,��f��ڼ,q�8�5MV|Q��m��ܧx�� �,�۱*L�F� -+y����Y-�̽����r)��Q�DY/JĬ敗[����4�3%�������Dn 6��R�N�\x�,D�,l�VYW��ZЬ��c��]��F5�!d����"
F+��Fn���켏u]˔�5D�M�&$�T�J^��Kn��HQMem��*#5��a�m�5�nc�N������jI�f�w�Zr}�`p�3&5��J,X)1���oVᣒ����@�*�(n�,˘�HJ;�^�O1���8JֻC&S����V�*�a����:r�[ˀ�2U��,GN`	T�%X��	�&�r�e�fO	{h�r�Fըխ�$P�B�V�Đù!�Ź��p��Ym�/��:*X�Yˣ�*\��"V�Q��k���QKR����2�¾�2潭�
�f�)\t7Y�Nl��O%I�	�(Q��n�wh!LU�IѲ�ج��Q�y��4J�"Rӑ�yӃJ���$�wQ�eS�'��3h5s�PY.#t
�U�h��FУ	�yG�X�m�,n�tFۍ�BGN��Q�M��/�Cwq��[�|q�ku�2���ܺ�s<���ق�9dF�@f8�-�yn-��sh�tn���t\WF�S	R`*j��A(b8r�lܗ[$;�\}wOP����d���Y�N�X�/D�4��(Օg^!f]Kp���kv&v��ƨ!i�#P��j���kUqb�`"�Y2�K>B1�b�̺��˫gL�#mSP�#ƕn�%mh�GX�E�rK�����4��+A�W�nMq'#V��Xq�\ۻ��HaUv7E,*�ɀA��$�ܴ*�$�W���st&lC��a�,�q�fm�8"d�Y(�m��R-��MhJ���%Ey�0fC�o,9�� �+U�Z56i�V�N�浛�%$����(�x��q�2���gN����f��(J2��Z����鎯K�$���/1����nZ�tv]��Mk�/�Y�{I�4Y�D��M��*�bk �t��~�tw2Q׳�Lğ�P�m�!�S.�ح[x�AU�f*�z��Wa�W���#�B�Ø��J����i�zE�&�rM$F�b�N�Z���C[
�
C���j�w��X�Mnse�Y��>�4�W�մm���c Op�
�ĶQǘ��y���J��2=�x31�r��ۑͭ{�ճX�ݼui�z*�C&��"��2�I&S/��e�5+&������X��$=3o0�\N͔ 0��w��D��B�� �P��@Oh0 9x�|[5w�GF��R8���f�b���f`��Jҳy�1I
o3Vn��g�2`Oq[/f;�(,��2΄��Y"�M�sI�v������qhp7&JH]�F� �:���kh�Yj hL �kY�4Q#�]aٙa������"cM�>Y��K�t.�n0��.��tݽϩ�1^�&e]YwF��C�S�$���McQ��B�����p(���H4)�i֩�����EB� T�:HE�w��(�ye���Ĩt�[m�V�aC���1j�j�v�c4Ӽ�z�fKDV�u�:K%��Cf������GB{re�Ȇܲu3>�� ]AM��0cv�!s7e�(�|k�7������L��hV�O=�a�[1��`��E������p�,��h
���(!�.�[����6�b
�Qͭt�cWui��t
Ki�KFl��uONmn�l�ᅇ�d��(RL��+�M
��n�V�v��PYle0!���S'u*p�F�xޓ.�k�4��b���w[���9k@i�ś�E���o�6 x*�hЭ@�p�'�Vw�`8)����V�%���R���3����e�i�Ѝὔ�e�h�P�Ь$�.�A�($V��>Lթ����V0�f,9��Vwi����2]�tШm'�P:�/Z�]�CM�h��8��%�l�J�v"�XH�n%��ce`�P�[���V���7N7t��&%.Jh�OP�PD�ܡf�Y���/�l���y��y�M��#�K�4曬�-^-����a�&&�I�r�8]^������֛+b�K.,Y�R�3e���,EN��8%�Ȗ{zX!����[�*�3R�����c���&<��:�!S0U��w-�I��wS.^=�a�"�Y)Tyf�]K3/P�Vm]�z�s�[h�ݽ�Y�n�+�®�O����f����:Ckp@�b+E�a1�V;���:U^���yAռt��zH�%OR
��N��j�LD��黰���-��p\�FnP�����8�]b�t�U��R)=��6���$�z���;MHvʔ�wP�������"2�{"�6X�*��T��b�w��ҫ"���%�Տ4͆Fԕ���1+kn�SA8Q����ɡk:G�u����׍��4aE�`�ß[E=��V-K�vŖ�BV} 6N�D�!P��׻�֩�k�ۑLY����P�Mr��
	���wX����ś6*Ս�a��q�X���;�D$��V>݈]�Y/	�ޝz1 kJ��{Z�&�K�m@�7-b�M�64�D�D�ڈ�V�t����7R�D��Q\�m�z
+���˼D֑AGYJ�ȩ�(,�hT��(�����-��ۚ��B��q����աl� Cr�0��x�;ٕ.�cI�*�x4�/2eZ[�[N�N�@�n�3G&���P�.��;0�Z]�+7T�l�Q=0��zx�]�`e�P��&9��NI�em6ÄA�2�G`MRr�-�t��Q��ا�;��M����)^��'�Y���f'zIVK��H�H�QVP�(�Jе�~[zn�fLX(]9�ѓ S��n��-�U�0����Q�sG�U3�^�pأ]bSD:�T�f��q7��fV^�V���ƥ��"4�EA�`���v�S��T"�r�m�[Sa�K��ZYИ�v��vY��h]�lN���ƈ��Y.��f��/p{��jͦ7"��[+���&j�{l�SC�C��,���Zn��2D�l�Y�K@+w,�
ו�����)�c)K���(ʬ��tJ�zpXȇ֭�4�L���F�f9&n��%�#]�����^�
�Ti�8���f�]��n�nJ�([���"U�O�JԱR�a��U�a{u�3�������m���"�1�Q_Ċr٧p;nq�Ϭɔ�7��4�`p��J
�ʲ��n�y��z����#�%�W{m�-fv�$fQ�S��AE)1��3��gaȱ�"]�p�{���(kڇ�x�v��c@�0��Ϙ����'1!YmE�6��]ԙ��͍�t�݀�9l\�7h����G<&�ޭZ�rL�q��"ϰ�J�:�N�>{r���B6��VVl���Vhj4��Q@`(��ac�m](N�nZ��2�]^����!�0]�A�Z
0���teB�I��f����K���fT��PN�H^�P^`�B�e�iZkU�*e#a�8���&F|X�LR�B.��Sa�����1޾OqJ�εE ��mQ�[�yZok�;�ҽ2�Kf0�`\�2K��ZF�j�k�V�K��T�(�.f�9�m�4��0]�[Kll��%B��CG,[b�D`��#^%K�J�aa��GU0�Z��t�+�Zܧ$�CN�Z�˩tl]���/v��T)�&����pV�5f'tu��N�{��|*�%+V��h��1c�sM�۫.�Nl[S%Z�Pb�:���v�ׂ�,K�n�5n�҉�4m`F�ٳF`P�6���$򢴵а��\҉XN
�3᭽t�-�X �+Iov�7��-v~/�g�L��k9xLhx�c��ڵIB�G ��K`S*�(��E��0�����-tu(%Ht`��ɛ%M-P�fE,E]���ŶĦ`8����<��1�8�ED4�f�o7]�E���q��GV�P��C\���X�e
�(���W-�t��k".�{&�2f�t���AekȫFV$�x�0ˎ,Tݵ�ceF����.��7�t���Nxb��P��l�Rљ$�f�a@����05%H��4q�m�Ku��N�L�]��쉚:u�*ګ5k^�:��dF�;��U�)�M����Ar�l��z��I��]�ޥZ�Ne,�F�E[B�^K��wP���ڦ�a��4��Ȇ�jR5-2���oL�e@��ܑmV��GyI�f�A�0Q�Gǧ�g�ǐɈ1�i�n��6��V���KsU�,c�n�Ӗģ#d�����X���*��c̙���������ާih��=��������*�(���wj��y������+o�u뺲;'ky��l<1���Y�s{4�c:��`q�b���>����zT��37�G�&�q�"�MM�������˅�۳�3��^�P~���%�O�\�i�����n�:���.��k7�w�;��T��>���;۷	��W�J��V��ۜ'�oN�aBrC�1�N"�^��w%��F���o��b	���۽+�W*�{	[ݶ@m�{�� �":�G�9��oBd\Xg[8	O��4���K�͙��C���e��;s�����ty��Qk:&L��v8���!�����k���&�2-�`��__,g��i��R��:r��6�,gx N�o�ݵ�J9��»$.{���K#�է���e�*S�}�y�%\f&8�w�E�����fHe�uv�nb۸&�t�R��7�^5���g���nܦ���,��ү�qiW�^=b$w�7�
��3;uồ +,�L+6o\��9cv��V����Ǘk�5�wgoW�s!�ۉ��L�]�#:�ɇv"Yst���uɭ4���@\�y�����Hgq*u^Ws����T�86�������L@p��x��N���0X�@�6���pr�6���a�A�V�u%�sxL�����OF��
�3aם:�[�K�n�4�ؕ%Md�θ��6��BS���c���]��]Jv�A�o�q�,ٴ)ҷ/��v�7����G�Mr'wZ���G+ ͒���X[ˬ�Y@^PH�΅pc���Q'˩h���re��X�8;�W
އf��r��{���R�43B��*o��o86yfS; �HD9`�ì<��ü<E��ز�z̼�3����"���K�7�
P�d�Ig]�뽮˥�K9ô�1M�/���v��b&�,��k��\���
Т�-b����5r |�u_I���m2�ƥ*��������ԩ.	�hn��gh{+�.���G|��>��Ai����=��3����Yx�������E�;�8��x�(C����r�sr�����>���V��.���"^���C�c�VN�A	^�!&�zp�\��ݕ�m"�,��3y�z�E��M�%l�E��1�^���i�>�Vi+|w�/���uA���ޖA�`��M�	��]��yZ]��o��s�i }QoN6�o�iէs6���˦A��P1�t��n���8Fǫ�;n���,g<�������i+��٢�&=k��w��^�'y�/���YV�Œ'��ON�GS�¥e\������#a�#����)ۯ9�k:�g6��:��� �gT�k�H˺�irALVՐ�ծ���^�I-(�䢔z��64�ʻ:�w�g�#�f���,y9��BC��sJћ��L�@�U�> h���q��~!*29w���ob]RF�ڜ�M��ۤtiwv|�ݐ�YO�+��H�O������`�/` �[�є��2v;����R�@�s�c�N�9`���-�V�5�u��������N�ِ�|�C^l��:��U0:^}����9Qiڨ
��GƸoݖ��Ǻ>!GJ�W$ޗwH�Q���D*�`���Y�H��mc�e�����D=��[}�dU'y�����6^�G���⋱�.������y�� �6��p���������ʽg ���qӪ���b�FO!��.�=bP��E�Ȓ�]g�}q�)/��hu��/W��WT�;��VI̾��B]˫��d�sG'è=��}2�G���	���\�q:\�l�]�e�:� �Ǎ�򗺛��j��p��	�.n,6�k[h���"\�PN������܉>���[��Ƹ��ػ�e�����,�nm���:uhL�y�T"f��w����5s�s�κṶ̆Y�6>��:..�����N+��5�"puK��p�ۏ�@��&2o��CDbcˁ+����9{�	��wS���+���óǽ5��Ń�6���_���l_䲺+ݽe�nt��T��zk�WAHj����0��N�*�ݾ��`��ڵ�jmXd觼�_m���v!D	�k��ı*%L��wڼ�V������4P��Y��<��O&�͏k���.�]�������;\�N���j������d'V��c�E�s�Oz�!���}�Y�g�E�s��X�E��Eډ�#v��b�l��ν�<P[��iue]N��%��\̡0[�'ZK
Ɩ�έ� �[���s��^ɻ3��"e���sjb� ���]2,I�^�b��	��k�l�0"R��
�S!Vl�z�vb&J�*�m�J��	�u&U�w2`l�5�x1^�Ȇ�NqN�O�wR�D�q�,Q�C��X ��7�/�1��n�i_k�.��
�T.c,Z`�A��4�/��n�ms��Ui�� �a��c������VP�SY^�֗.���W�,K����w>:gV������EG(�˛�i˸���k�j�eP|9�n$���%����fLpL�hA�}��w���6�R��0��+<���8�7�ԺU$��3��n�f_��-�wC�/���֙��I�.�opsx�d�z�B��A6���&a�N����U�$1hOG:��a�`����6��\k���W�)����{YC1e��͆�#�'Y7%��%̣�ͩ+�mRVu�h�� 뾛�qb�7Q�.�)\���=�j�,N����D�)}P�)�(��%N�/�.�ٮΪ9��n�=��;i�-E�i�œ�9o]`���o,[D;��/Hو��$Q`��Y�|�}I��@�f�v��f��vu��n���Z�Έ���]/�][ޱ�5%_M�j�ˆ�mؽ��TG���V�tV�M2������;�PD.ܻ���[��&�'<���;BQP�ݫSz���V	y�h�0�;�|�]��౓��vS��*2\ԃ�[����U�����	l�U������]l�������[�� ��ф��{'%����h�!��W�,���d��뮘�
��g%�쳽�gn%�nS�2���}�x�!�6�����1���W�̵<��vJ��u�=��&k��#}O�7۳���U��#o��[R��\���V.|�Vd�b{w ��ʈI�kL��K���Q]�����Ω�-��rm�q��#�v�ۋv���n�*�qޢ���Ѿg��M�8�-����<O�.��2��?d�̖�<����3Ns�{��� �����V������,��-��!�Vh2z��w�&����B��nnSݢ���h%�GJ}1u�1��`������
H%�;��9�B
��=�nÞ����gO4B��͌�b��N�hֺ���Rq���+//J�'��cS�s��bC��v��n[�Cr\�
��:���(��L��wa����������<[ �MM��Z6j��xn�Wz�ݪݩ?7}�nGK���<�v��{��uu�;ҡe^����+���c���!hB0G������@�k���7wi�W&�,))�ZWY7`��37H��z��҆�4FCf��J�pP9�b�N{獖��s���Z����A�h�n:�+�c�#�U�t�m��w��y�=�L�����Ӳ�fu�mҖ��'������)�m^��zJ����32e
h� @^<w�W;��n��38jh�ua��E���}�ڝL]��T�1#Nɨ;�df\�������8w�JQ��:^Q�%#�J���kH	����+x޽�w��wf^��!�A�D���1N��q/��I��O>*þ�^.9�;1�Ίk|-ed"�B�9�wh׻��rv��n3�%֒.]Iuݐ�k���	Z�ĩI��Z�>���vYj�S�9�уX��ݑ�SN�%p��&l��f��؟=OoD�9w�-8�i����v>��Hbv��J�G��JpF��G�o�T���o�
�(�G����V�ۋ��_J�"(�L9��ɠo��}حGn'�3��2�2�,����9��;�ct���ALn+�Y��VL�<�=���Vo��$��L��	�TI��T��|�Ҍ�U�B��^�4,++wfax� ����`N����c������՗��o2�ʝC�#;s{�Aߣ�]�x�ˏ�kdP�f_4d�d��v��5]4M��-��X�5[�8�b��X���9m2���s�/{�ҏ�'�����-ҳ{��@k �\ǚ>��l��)��gKJ*_o0k�i��C^�KO�^�)�{]��L����k��^fi�w�	�7�!�]]�FJR�s�"x�eenS�[-Ŝ�1�t��,��Ԁ�F�$DөH<�POm�3n���G8�AB�$#Y��s3��y�%�8���X[]�z�b�bbӁ��e-���m�N�t�X2�7�q�ګ\��|6Y���5ҕoDR���	^���l����%JV���-ձ�{ϯ�m.�
N��@���rI�G��iݮ�hގ����KmZ���ι�������8پܐ=F�Vb,3M̮�ӝ�����Y�_$Ŕ�l�`��`�ie���g%}����ꏻm}B�B�y�(ߋP��}������w �y��-ft�Bk���[7oq�鄅a{�"�G�]uip$R�N�tnmXY�8+p�]��ue�2I��eMy�v��N�j!�<�\@Vdmwf��J&��7�Z��:)N� �{/~�o�c���iF�����l�v�^N	,�����,��r	T�Wp�f1�bZy�H�I��q����z�'bf��kQ���2�}@ef�A�W��-�Gp�tn1C��]lL񖶖M�Åm�kg5I��l���ںJ=%.�T��9�a74�q"4�K�F���J�>�h�e�4�d�l��)�9*U�{PܵK5�t\�y�u�<-��6���m�P�ސMZD��+M��%^��ߡ��fɞ�ˁ��`L�@IY����.�	@K�u,W�SW�W��&�U��i��t0&0L�9�o��׷�|�1&I�� 7}�ٿ�r��hd��i�7[J����|d;�4-�ska����1؂�we���V�A�W�!��xӕx�����
�k���(1V<�PJf���������À\Z��h����Q��z�{�惼:x"rl*�^�Y��l$�m��,h�ٻ��d��'P������ :�K�n�W\U��f��$�(� Sd�����	�)wY�9<J	s�3��!|z���@6��Z��o3v23P�v��x��/�h�j�&{�h�Ӊ�۠�sɼ�
^0!6���%�]b��nڮǃ����s\���Ō�cM�x[�b9$�<&*z�r��ƺ��i`+���n��7��"];6��ғ���I���������:�oL�S�w�Xm�m*���i�����w8g[ڒՓ�g���RH��:�P�7�,wi���5ٖ~�%��Xv�ô��`u�VM`�(��v,8��P�^�M5��UY�3;���7�jt��8�>s�Jb����@��0^&5.��5/%6o(h0l�Tn�S\�Ά���+Bcx�/+RC�B�\1c�Y߱Xw�2z��3fm�gx��ê�q�^�-̑�"��l�r��/Ueu��9��ѹ(�Ŋ�����m���޶tS*Kc�R��5�U7���K�;Ɗ�=������t�n�]���Y��Q]7u������Ugr
^��&B>e��	l�e���9�Z$ax��͎�m�=�p`��Cr�c �Z��$0�&�;�G���$|z��J �gf�R�^)'m���Qmڧ^(�b�+�Q�9W�������/�}p��x�ȠCL��o�o&`�Y�/��vYx53ȫҷ73%� ]"���-GD�a׺;1�����9aD����4�ܵ[�S6(���\r[����ĸ*��ቴ�b��W6F������7h�P�������;
�ВXUo9�er�ǵ��rok����Q�~�kO�:ά]�9�6g!����Ƿ�|+��r�f>�:9�y��x�Qu��`u��rG��r�@@�-s6�5ج<)ǌ�3x�~�æ-W�ޓ�.n﫛)��aT����S8�Fԝ�u] �"�.��q���p@��t���V��%g�f%H*I�P�g#���ӫ��:�m6�rk����[f��=n����gz[2v?l[�(�kԘ��	<<��Lh�Ռ��0��n�u��^��y���6����0V�e\�	d��f�	X3]���Ԥ/{�F-���Z=0��@��]����w+�اK�m���K��E>���ל�&U_^�WnH�K�rCjq6��*ү���(d}�w�7�m�m�<)`<g	�����!�\;w
��{�7W���b�s��`*��d4:�U����2��G���0qS[ q�����|j�������[�ۜ�w��{��\�A�V�s��~��װb�e�E�'�P��@}<A>�kew[L�9�}��1�wnP�>�g)t{o������.���#l�m�:ή�oe�_v�Զ�nfn�
ާV����Z0��ou����z���ܽ}h�����P��IO��j^�c���w'��n�.�^��W�[I�Ż��^|�����[s���m��m��m��m��m�z��N�_W$�@xs'ɗ�gi�ȧZf�&��%=�q��P��:r�t�[JV��*�:����E[��]�v�>}Wu ��'z눟��]���Ȅ �$�	&��V����>�L�]�L�.Һ�HJ�w{�Or�Pܫh�8�)�:3B��Y��꠨@x�y7b[`�v��j+�k�x���>�n�Uf�R�z6���r[��G/�9k�bg�#Nd��xnݸ7۶�;�W�Y�8���t8�4V�GR���SN��AV�DG��ߨ��&��������L]LQ�9𤠸�׆ �e�v�*�鴪R�O�$�̵�:�h���ԳPq�|`Z�6/L^���9Y�j�R��P�7�8�s���EQ���}W�wnƭ�]aH���3�����{Zk7�������5�=�t�TJ�c�3|Ͻk����*�ay�:k��`�C�=�P��^�j2ƲXmݲ;K���7������u�ڈaqn����ՇJ�)��r�cfλϧ@�������T����[��B�x����S#X�/l�	��<6f��l�Й�y(�Ü�8��H��B�z�.0�X�"���}N;z	2�,��Vz��
�߃�ݛQ*���� �voNU�ޥ�V��lNoo!���:�N��d��~�9���9jL=/,�ҞN���h��J*���6w��-).@޷(a���f�gw�q�
���P��Q^��TWx�~I��nm$���	`'�������Q]_#}�q��;Q�, �l��X�l�m�Ŵ*��z�ؽ]��z@�+u�����5@�gA���m�>ƨ�\�� �s2rz)Q \�^LB�^����u�Cǻȅ��,���=�-a�G�>&#���z^�Bp2�kUe��0����������w��"o`��6��(���Գr$8*־�M�Ӹ���6]��x��sz⮾�3�#��9�mu^�͜��ǽv��:q�{̮Z�=�f]i��z
����_	v'�vRa�I�)��ML�����p[����i;�\�J2�ktֺ�M���R�e��Cv���i�n�78D)�-�����fz�=��
�L"����̜̕�Q�u�������F�emg�bN ݬ����ff����_	A�Nuu�]�?�؏oxY|zRk�͙�`!އ��S�VHh�����V�M���t����
��^�Ѷs�f�k��d��Lh鸫w��a����pͨ��k���SQ6��ZpC����5(>!Ġg]�]5Xi�xc�n��L
�Xb��WM�iV���ل4�
�o�!�d,�6p!}җ	���Z�"�Z�5tH�rGϷ4@�<O{��r=n��k�/��]b�r���S:qw:�S\!�k���I�mD
6o����@}�J�Y�I��������N��dSt<{����J���,��]�X�	�D_]����e>�yTt�!�5Chm�<a�,4�XE�-Y\���� ��D).�܉��8�ֆP���Ը�s0^,�ye�I�$�C�G�����&	�cZ�*�k8�>��re� c� �=��8�T�U��M�ϊ�M�be.S/�5WCB�:�4e
�՝ZS1���	��<qC�t���y�Ė(�
4n�A�SL�eͱZ���j��	X�c1������j�I�"Y�����oU�8Wf+:A��>�[Vq�h�̉���AsF=o�yo�փ6d����w��܌=�	,���,����MK�U�"�y��B�e\�V	�����h�yd�b�rt��J��(&Ȇ�m��(�L6�v*�׊�-e��c�J�-�i�au����9���<b���U�F��M!f�����$���[���0�:�lDz<�!1��3+��E:���t��E���2�ަ{��,+���R�c,sc7E[�-*��܀��>:R�wk@{��h���(�m�%�s{x
׃ތޗ������Y=��c�'��c]ge��-�����B�����|vV�8�#��@�ui�����f�N�� }��P�x,��y�NՍm�X�e8&R�[͈���`S��X�W!6@��0�-+� XgJN�FU������Eڼ��e�fAL2����3��W`w�lN�`>&�M[Z*���؅�1��M�w����v�+����� ��qd��Q4�	�)p�뤜��X��0�k���[�t�̏��D,μ��.������\��n$���G�坡���z]���#�x�{����J�1�;2�Q�';w	�cMv�՟�F��'�emJ���=fv�A��Ce�L73�:=�f��
߰т�Y|���w�V��`MM�6�2v�֪ayI�d�w���IZlh���+i��4e�A٦�����Z�)Y#�|�ڠ��Ua���	 �i�*��f,���� ;\cUCh&�hDo}m��pCO�h�������GE�%���3��{4�b��$�s6]�1f#1^�).��,N���'�����8�,�6�� b[W7X8"fan�eᖫ!r��C%��N���&=$��bYr��h�nRL�Ǯ�]Y�5�Ȉ��m�jj�e��A}�ݵ��D+H�vgZ�˄bQjTC�{Ϫ憴��T��K�0��O��)W
�'͇<E�A��z��������6��P1&]�N:V�BѼ�
�"���X�����u/8��ȍY�EW%ɫEf����@)�]���2Q���U��X�ѽ\�17k��*�HЊ�]�����Z�p�܃�B�v<0�S���x�׭���V$TErQJ�������^������
��"��]L���}{0-Ԡ�.�~O�`��y�4p����İ��\�_Sd��X�KgI��dE��2�]��v5�㋠��M�<q��7���w(��� ���,r{g������>��AuҎ�;�Ћ��Wx�يG�b���:yo��c��.q�^p�h�n)^Цyc�h�F�S
߷N��,�x,����׼d:%�D��YY}3�s�>�Wp�{�7'Q�;�%�g)[�L[�*"3gn ����b���j��uw�h��f�׳�G\gv#���9Ϲpt'5��{T/w�"�Fo%
���ms�p����Ip����ф��
�U.�`�F͂?9�<�v|�d�R{F������b��T:f�[�¦3LiQ�=��wj����Ȑ,���48�BA�A>=�z�
{Ԋ�|�qs-��<�E6x��Z�8w ��9e�l^�m*+���	14�8#��f��Kl������:N/Fа�A�:Ŷ{J�Z'��̻�K�@k����0g;��&���˦u��n9��� +�Uۧ���7)�
ġ{�/7%t�ӑ��`+�f65vf#���b|s�T��w����� otѺ�v�F^��U�����ۙ(���h�K�-�W\��D<n��n����f�ƣ�������t�*]��0������nU�Q�7z�	��J1֚���]o�a�Y���	�t�T�W�暑t��6�Zy��A�'���I�an��"-"��H�WP�R����5�*��J���'�&��Ы4<|��ٽ��W�A1u>Ɔ�c���Z��%x����#V3h,�ب�N�^s���h�_%�o�c��k�?w*�������.�b�vm�ſ����jT��<�Ve�x�T4�X�C�.�A-�lv��/�su��ӝ����h� X=C�6�.�)[w�z��6�a[r�S+CtY�ѕ������]W�|]����).`�7ZP�6��@��7h�G����c���^�8I?[�n����1T���LU�����+�T\��uԮQś�JG"VX�8�{81zSS�a��ȣ!Y�`��-�Q�^-��3��oojka�zP1�����ǫ�u�4h��\LB����ѫ6ˎ�G�|��֡��[/Hup-�V�Ze������֍�B	7!JBy�3�u��哇��3˽l�o��-�'�4-��sF[�����0uH��5Q�y�	��v)0m�%�G�u���ݫS�=�an+��h��K�.b�;{z��kf4���c����@V���|�9�̙�5:֌�.bҡ������j�����@XXc#Y@���;QtV��m޹j|�Y�2<V��L՛�-�#�Z�	��7f{K�}��J8��]����F�Z�y�H3���2(&���[h�U`n���2c%��r�+ֳ0�}�ct��_R���䔕�\t�Xm<y#�K.�⧎D� �jH�9\.�t��[VY�e�[�Fo�0��w�iM�mv�zZ�*����P�ɐ̂�Z�w�x�|��4��X���k:H��}�d6�հMYD��Qr��/��-6آ̬�������:Q�R��f�N��F���HUՊ��$z�'5��!��FYz�&q�ۃ��x\�K��&�����bL-��#m�kk��𡒃�V/J{o궹��BJ9��T��a�)�6�/�(˶d:���C�z	1s���_ۭ�rVp�t�7�`/��칣��_62������7�7N���K���$��w:`3R�/ڄ�5rv� ���q�;����iB|m�����ɜso����X��77d�%mNyN�2�r�y8��2���̽Z��.v��ӝ��ɻ2���`}��{~��������.R�'^�[�5,Z�L�.�MAz�rɋ��j��m27t��$��6v���x��������5���2�SC�
oO�L��NfC�����W ��	��m`έ�]��T��o$�I�t�J�:�ʲ�,��ö�{E��d��b��Z�-�٤U�L�I�0�93V-��+�p�[G����A�n��z����V:�$
�j�,���of��U����x���6�R��P� �凎�+k�%�1����|�4�93)+��Ru���gd��Se�<*z�V�r�Ha��&�էD�^��/��0�C�y
�z��}�tu(x��)�br���'(���l^�ݲ4vu�<IN�!�w/h��R}0���W���eٗk�)3���&���U��6rf����B����W�m�|�@�����fһ�{��hJ��J�;�[���\'hdÙt�ov�q�P�ys�X{Ь���p�鷥ɛ��\14|"}�M��8�f�T�~=�%�ƅ���v��$/���Ծ��ꖂ�8O+|���%	B��{@W��W�f���{Mu^��$�%uM=ʳ#i
YY!�6uЇ��6Q�2�`j?�^Yv�ZF���he�}��36��%���qx�]b��Ѫ�v��9��+�����Zxgd���9@ZtUͮ�]��s�o;��[��NQ�U� �Ӳ��V��J����B������7�|�S����s�m D��YJ��<-Z�������Q���g��]���c�����k�<�F�P�����p;5}�*�c��ȥ
�YY<��ᦦKg+���e{|��n�5I3ɮ����m��)��0��q��3�ۤ�jɶ�P���8x�zp��W`(p:�c�K�Y�V����ۅշ�֗_��^�T�$��	��V��tI�1_'�ٕ������ng�y��+ar��w@����3���;�p�p�v�q��)C@B�t��q��B�&�%Fڐ3f�Ov�K�܎�10T}8r{އ)���f�CS|��ut�<��+UsB+����`NuD����ԁ�έ�GM��ۂ���1������[OO7� ���>��/+�Ѳ0>�I��Y.96V��i�+��]�'�{¶��7�d|,��x��N�8�pK��4G#w>ը����VGB��Q�σ7�����W����[�T�Y�a�QR�Һ�N�l�)��_\�:]�n"��Y�]����!��D������*�+��Ŏ��vY
���P�92���y5����o��u�o�[�cR�<NؾKs9�Ky�Ǔ����Yl�Z^�q[�b��Ƀ}����0��9�]s6f1����{ͦ����|V�ۦ�=u�_+�o_[�S(	��Q�#'�<a�� �
�[ɇ8�2e�Fyz��<���E�c�#�o�m���B�s��kq�+:��{�S��#aU�H���:�X�$�xjPR s��.W����(�*�Ӽg�:���˒�m��%[F:�͚�a���Шb�pļ^3)�c��ƹ�(��8n���v�E��ۤ� �W����l�Vl��t�`]3�zZEL-��KR�-�Wn�\�}�_QX�]]�:���A91������d{����aa��ޮ<�|y������$ag���]�:g�}I�����Z��Ƶe���x��<�Z�){�Y�«4��`i�u�;�z륑�Pzv:��Z�h���:|��s�T��:f�xG��g���XN�-�Ex���l��v�uyR^�a/
������i��of�pǔ���7YDP4�p���KwHb̎�Ë��֌�E����Jt�e��tƥ)r뇶L��{ԥ08vm�]��jVߨ��홸��Sњ�32Z�u,f�Kpl �â=q�rp���}X\�P9E}�
hP��u�.����/	���l�w^���
n�+jue�8��N�譋13��9��P!w-6W���\�򈬭w��4�J��<0!�.D5XNN�Yd[.�B�Х�'`O���L���&2#�^��=�}��-���M�;kD���4jr�yh��1�(3�i���J��$�t	�-���݈;W�V�1/w�
wJ�3�̚�J��%��$�������x�r�է[S^G�����=�z�%T�݇RKO�p�LQ�-4��8�՛�͑������3H���Ǌ�5�H^�Z�47�h�t�;���}|��ͮ,-�b ploE�A�^���YD��G�Q_R}�
�X�J<���V����sd�}����WZ��JQ���Ƴ�3�7q����[v嗀�ۦ;NZӕ�U��m�WVosP��xpYʸm!0:��^rn�m���T������t.�]ݤ�z����
G��{f�}3"��=��Q���	'��T(�d��5f��:{l�ġXʙ����[���]����ne(BU��7��4XkY�gv��}B�:F�6To�l��p��֢G��D�N٧(�p���V'`����}��Bt��g�]�Vi�BBNgY�����l-{	����ɯM�wI��g��QϜVy��������y&j۪[���WP�ѫ��S�Q���f&n|3�Ī��XỦwM�G6�!���M������L8��N�K���|l���*�M�����y���;q*�Ø8`4�j���l����<
tEr�h$g��7v{v��̚�3lWN��Ԁ!�DU��u�H���Q/cW�a��TҎMjv�	�|K:�d�S����\�=ydd�������Zoٞ�9�j��/����;6��m�o)޿n��3����i�
ʑdZ��R��m,eem�ֈ�0��-�(���i�9�+"��jJ�(x������BB�TI
�Q�J� T���\a+��!�fZ���*)�fH�M�aG�X+����UPLd�(J���T"Ȱ1�eaMXX�F(���`(V�r�E�+,��c
�"�%jA`�1��
�d�
((�EhB)`m bLCH!��\j,�-eed1$�)���%dR� �U���&5��f3c��`��}����u{:ZF���}��2'�Ƽ3��`e�*�4�-�D9c#�T4�CfX(kY��TFwخ�G\�K���ga���o)�����V��uU����P�8;�vܶ�%(Gl��q��Y�{�,����ۼegPZU{��m�iU�>| �����r��g�����A�OV�'(�~TH"�8 �Nd����1ӐjEt�V".�:
'!�g�B��[�L��u![id�oռ�����FC��h�J$6C�U8���SW��yT^
D0���X�kn�5U�jz"챂z�W�eC�p�lF4Έ��p,�xO�;v8l��{�W�U�9���"6_$EZ��0u:��x����b<��5.���Q�j�ۭB��rK%��Fér���EEA��E�>ީ�����5�FK�/����GH�6}�f{���:,[/ѿ�I��G��؟Qu��x}+���ѩ�E��79�*z�kR�]���٢ӱ�#�zl=jH9 ��C��^�]Ss����o�ͱ��N�ګo��A��&���;�L��Ѵ���f�h����/v���T6db�X"�䗞��~�qDO�9� �<��4�Pul�ʃ���a�w��fhz]N���/��~��\���ޢ%�Y"�m�y���b��%ޫ��@�W�3ǾS��~����(�$�������������[i���ݶ
� =�� ��V�ذ��њ�m��[�_����r�e-N�/\��n*WFM��5ylH���C�νO��2�l`M`}~��\�P�Wt�N�.�4;R�Af��:8&���qq�(2�d�RΰE�N�x�9ӊrUtVϗ���m[o�ɭ��������+;昺t���P�x��S��< ~��AX�����V�9��]�<��$tζqt'�
��buE�2�l+5�ɚ���s�Y}p����/�"c^#�UmӋ���(^��B�B5[�U�x���r�MU��䠚22�G,�~�ٕ~�j��Лn�I��J`l�X����&�`�Mc�\�e�p���\UΩ1�+�*��۟kd�M�NLP%l�8צ�P%���͆qv�b��%��4/��؅\�XѴ`�r����[�����lO�_N�]�0�3d�:ާp�(<,�4�A��x���A���m|�g"���Ϻ�y,�2	}��$��]3�&��Z-��Qv8�F%��q�/�qiၼ镑tn��S{��;o[�_�v�:�c��]�`����V����6Oi����ye�_]u�����˛�%�*�gR��Ȱ���L��n�g��Mr!@b���܇��rt�ձ5�fE_�u��wV��z�x�]���%������|\�פ�B"����&�d�<dN�F�,6�k�cX��1��&��0jHhEG�E:%Y�7LإRs�^�t�&`�N+��%Z��)�1y/^��
DC���A���	~�/�H��#�`�H��SjV����/{gTf�����^���A���P�Q�QD4}���CJ41bv���a߷��q�g`�l�.C/ �P����v��2�6C��+�ñ<lV�l��yj����&��MT�[[r��*�H�"��e �X�=�=�:ν�p1OFeC#o��5�RFM�y@eŝ��b�f�EE��=���6�8W��λQ�m�v�u���R��'g�@���>�|G��b�����Eu��1��C�q=u��p1
nx0�Gs�z�W@�~�{H�v�:�������ؔ�qW�@C�`Ս��pDu�WRz��e�s��^4��͛R
讎�Ẽ��-L7Xe�$h*��]�
�S��WY/�]z�����u+�	�'Cqd��.Ş9�N��j����-9{*;��}[����͓��ͮZ]\L	
���̻[c�����8'�U#���@��X0����o_}�<G$�D��
F?<�^�n.}j�n������7nЭ::��Ce��(�h�"���d䷞ns�*-�]J��a�q6�ҏzѭ�/`��6��K�#��֜3'���;�Ƴ�{��t�Ih�x�c�DYpU��˴k�0�ي}@wz��7)X5'�)G����c����ҹdΊ��=�'-�����[��#t�hE���H�D�dڪ��'k�0}�p����w�.�w[S&��A��75�i�4�������^@�t��Kz��l�o`���=���h*i�Q{7
Bv���B���2���@���Ë����W�s
�R�2�f�U�lㄮ����@B�G	Nloi�C�c<"`�]�V��T�p�c2��vN��o9�OC�e-���F���le:�nPB(gU�c�f�����Հ5�u7-E���G�ƆKG��z�=R2�NC>�.6/
m�m8���A�L���;u��9X��#6�v�sq�I_O@;5<�s'͋u���d�X�NK���Dz��.���&�_�Gگ=�������c�>��T���K�)}f܉zVM�=��^�����T&s���s<�̅l�_��l��fh@�sқ��kw�.Y�e<�o�a�l�Ԥ7�Z�PO����y{�Y�mmVj��冞�=��w1��(���wF����|v�/��_B�g�9�3EE{��1X��S,���l�;*gX2V���"��sup9�\[����$x�}J%M�#�&:|@��bu���]�̹Fm��EE��Յhu5>���B�o��p�2Tc��C"���j&�R�	LZ���(��/M*7�Ϙ������霄#�B���s�6�_Pq2;�d[���A|�f��R��Hl����`r3��Dh�ڭ�R�Q�TX���y��{�������s��Q�F��>u��.[tz�����*&/W�p�!T3�ʋ�;
�e@��/%�V�q�}�ܥv�s�E��p<�$T�H��������&:r��Eb"���(�l�`�cj$�f��j܌2�H�=t����q�7�E�%�ǈ�J$�=f:m΃0���cFϣ��oYh���gx�
�́�)I�.�W�@��ŀ�m7�,xR��xH��V_=���=��2�:X�����q����3�L�����#��F!���*�1���Dy՗�&@�����]�^]W]��f"Z���ߐ²�x��R�{{h�pf�2-���2��+t�%�\��8�U±�oc��}�r��C�� wJ��hN��f}���Ő6圥mD�dѾ�0�"�dn޴��"�R89�y�.T/��gS��Dp�5��j�^eM�)�^5�����_�}��s&n�0���N�F�I7;�i�.=S]� ��llc��r����<+��r��������fD^�[�Y�gl�okobڣ�E�.e�P�/e<E�b�EV<��uQ/x�s�M�O!⹜q����I�j��/!�qW�:�&��͓�92|��:����
���[������)_T���^��QÂ#�*C�pW�t���j�7��E?[�_pv6{���^w��$�g3�é"b�k���T!C�νM�jC���V�-{�>��9<� Z2/�>���b�V�����*Q#G���
T,�JY��'n<\�N)y]���9^��B��
,k��>#�-��M1tN��xl5�=+�� �u��]9��:��UlX�u�yG\��ht��aBx@�	�� ����Ǭ���6�����YB7�Y�Z��}G�z[اaS��>�{*��qu!@�1z�BtB�ȇ=�J�XĊ�̢�1Zؖ��&��9���7w�,��h�6c�����Mc���`ݷ�V�na��m4���]�&�)�����:���������n��[�֔���'�+�ľ��T�
�88��<�{��.�L��4xV7֡H\W>ˊ�پ��;\j�%R�2�͹/�ka<���L�ʿK���>��ЛӉ��X@ٸS0�:��ң9;�Pzv7q|���O���ђr[�; �*��gr}m��7	Ɋ�D�6��aVD�}9W�^��>�q����yo�J���X���:�S���:��c&sZ;�ļEnC\�:*$5C�M
Ѷ�jA��;J*/׌���x�����	�P	s)0��[Y�;���9��8"�q[R|دE(F�"��uW�P;EI��rĘ, �w�Ed�Ԇh���ʦ4����dՆ���>hEC`�	Vg��6*NPz�ͭ��NN�Ѵ�;3]d>����(��D7�]<��̖����¦	�&�vn��ی��������_8L��Ѱ-�)N�xEB@e�p�*�}�qK(�;�QZ>����Ӽ7��u�˹��m켣�a#��=J,���p79�n���W~]B�����\o%Ë�<��f�:��ַs�l�=��U{i4Ng��Ҫ˭[�0� �^��8 �^�$DmAP&ֶ�&�"^Q1TH=O��hO>̽ԁ�b�yw�x�!�<,>�ת�:��ͷV����y�w��ThK�[c��k��{ް��l����#"�X��������w6�:y��Q��p\Rѳ�'-�+�U�4�i�<_N��ek朗�Ks�5M׾���E���ߩ���z��)Bz7���e`�Gï>�Zx��4�\�JK���j��7��X��-'¸V�˃�<�����s]��]U�ݼ�(��{ϐ:��Ɂ�ơ^x�P�%l��J�������/��sX��35�Cs|���}��f�1��sNuN�rD�wj,�uW�q�}�4}�nfͽ
�E]:���؀5��*q&�nE��zEd���P@�[2��������E)���~7<sZ�<�3�bcb(~ߎ4������Ճ�?-��wL�ʳ�{ڮ�mւ�O��;O/�ipnz��qB�>���N
���@��"ʌ�^�ƗD��tsa�U��|]=���}�j=g���F Z��B/�30.���"��M��_C��g�8��%8���(�\];W1�-�pURk`�:*l�N$�@�ٸ���nzxɨ�pM���:�^��rk%As��*�� �6P�q#�d��4�..��Â�R�@������E=^��1�ifЫv��@�X�gx�$�5;vt���ä���7�\z�3:�ꕲ�Ί�Y�'�9��:EjD8G�s/��"Ѝv�X��+�l���@�s}���IѸO�c8�5��vN�	l��8�x���h]�*��9,Β3+�G�p+*���n��X�� 7�6�Ø�j-���v�����B�fTd����U7َ��S�V�#:K�4$zX��Y!�����;v�MvV�i�X�d�z#ap���R2
�r����@�����2��+��+[�V)e�s|_z����<as%�sP�A�A��k�T�
�صU��l�^B6iͪ$\V9�w'ft��������l�ؿ7��:��ңc�h��al:��b3�S��uv�����^rМv�t��w<ntF���_6r�N;ΨvN���+<���&�>�Z�7K��e�y��G+�*�u��7�h��*ĩ���'a�uJ-�z]�ٽ8t8�E^��ӛ�=���=AV�EVǪga��p�EҦ�M�W��+s#��\���W�����w5��:���+��K��莙�eG�ǙQc�g����=����O�2z`�O�|�����NO��ba)��1.&����>��+_�τ�,W��;o�bg���
�h��+j7�,��Ťe�.\^xw�ü�>��V-���I�=r����f����U�.ա��H���("�幔�o�aW3�
;��$�W��B�����B��~#�ya����u�֞�gz]o|Ei�u���ZR*+g>�\u�ہ��$T�H��2q��!�q�T��"�v����'u{�C��W&��\�VQкll���
Q�ȧ���7�FC��h�J$��wU8�9b�C�� �ؾ�<�ce��x��]7�)I�	p]�r��w.-�8"��<"�����������'�WoT��U�;�M7�'1��t�-瓹��1�="��^e!�9���3���g=}\�@/oT��FR5��j_��l�NV'�O��EuDC�����}a�2�a�,v4+8mC���U�4ߺ�x:���SX��r1�p{�h�1��X��f[���h^�|�c���^��f�hߛ��&8G��S�_�ا�U�'?��VG2�[#E�]v�5�zu�*0�n]!:�c]e_����s�}�nQ�P�p7�Q̐�9�0q�I�gt��`٤ �A��Q	y�����r2��<;BPs:{t/׏}Dw���a�ޝ2��D:���$n*��ኡ˿s>.��?^���������vD�d4��~@�d�E�5����ՑJ[�w�g�z���f�=�`��*K��tnჼ�ܵ���7:��z�'�3{q7q��ydc�3z�!\Γ׼a���E��5U��:���a��n��qM��{�~}��4�۾D��z�S��"&��/u����ônh��U�쓰��r�T�G�{ai	�W�^�.���Gݝ�6��]�W��_<�vzC��
̇�+zӵ��{�1�}��=��^$��ޠ.�u4�:$a�N,��w3���f���.��5�����7:ŕp����g�_���e�0*��ng�(���6Pf��M�nx`�oZ�X4�n������h/g���e�t��%\G3�����b�g�``��Y2��h�ұ��οv�I�E~''�z��/v\R��ɻ;R�*U�6�@PBd��U����>�f�J�9|2�N��\�L��
ō<+|���z݄���_[�Z��.V]�"����u����d�u�#g]�}n���}�O_Dp%fޞ(Nۂ��J�,r�a�p�)ps�ت) 8S��2�"�R�=�#�p����&�E��C���}0�=-�.��$v��}GfE��H�¼�l����yE�v����T����;�=��Z'mĤE_Fs�}x���Z��,�{7�y0B��"�R��N�[�S{u��#,+!�f��(vP���s���a�"����<�?�ͳ�_=���3��hC�=� T/P)P�j����ĵ�8X9��]*;KV�[>ET�Jm�����p�� ���E���ـ�.�(�_K'en
�Ӟ
�t�;�:3�P\:�dԌ΁e{�n��׵�i�'eǐ��C*)�͇К+��j[�3�5�ƟK�� ��
���wA���u��q��s��A�ćX��y4��9͛�������Gu8f��p��ː�ul�V�ժ�
V�a�E�s4sgY�}�h��*63i ���,ww)5�q[�ofs"s�]C�ץ���$����C��>���7"ν3Y���`�=��k�J���X������q�k����@�8q�ƅ�$t��g�QS,o��W��ů�P��QLl��g�Ci���r����-�-Lw��O%R����-���"�h�rp�<|7|���e��ݛu�q��q��8fn���� TN�)L��τ���؅I�j��V��-�=�r��[�tPw���binaeM�(�ٷ�EjQ,��i"�\�Љllü�+�]�3�r�-
��:��7`��߯��4ʒ�5Z�Q_=M�(�򻋮��[R��nT�/g���Ws�ݫ�޽�p���;Sr�%���� �Ū��hP��^�(�6V8�Zzo����F�C��ӻ;�8�1�4�3 ���A�t�ew��}����}m�M����_�o�������(Ad���*��Rb �*ŊE�,�	UT����dX�T��+$��1�"ȫ (KhAa��C)VAH)
�d��VdY�P\E"��F"�r�*�ʚ�"�)"�̥ *�
E�
���,$�)��hAdURAIŕ"�H#VTP��A�V*�d������T����2�9HV��-��"��F�X���@ukb�%f�0r�V,E
��U[lIPY1�$RVYY(ł�B�� �+"��2J���
�Q@U��B��VAB���E��h�m��y��}u�{|�'{�����w�M�:�N5��*�foU�$�va�Su�7u��2���j�F�E0�I�G�ٝ&6������:'uG��R���������TE)dk[�������8����m$S��:)g����^���;"��Ka�*�ڵ<��3�d�w���w#R��_�l�ۼ�~���M�!����	�� ���A�v�^%ˌ��w��L��\���yl���\Lm�۪a�qu"�1zBBpB�U�x�2�^ �}���7�,߂�z}�nB���m[�q	��V%�\�i�6�8��ஷ��*�ιW���Zظ�f�Eq��yԃ��ue����8)���G���?J���e�aU��
�͘��ٵ]�G@eg�GMz�]�u�E�F8�;�7I�U�.Գ-y-�+��z��O�5��_�vӼ�5��z����A��y�������6����rǰ�A�!�7�OM)��S�HVFՈ֢�"��+�^�#\����\dn}@��ӭ��3t7w�cPVd���O*�e�#��M_�F`Ԗ�P$6@35�ns�r��J~�=&�>0MYt�Z����]ը��K�~��g����AÇD�����i�̓��Mf���(w���~0U<Q��H�8��p���U�|d_��}V��^A�o��92
����;��+�	Ldѥog�іF���ǔ���A;tNp@̮�uD���[�2��6簾`�%DC��zu�����
�-
�_�n=מ��|��ɞ[{��Fqp�u�b
�5\:�U�1�|� �����������q�,y��u'VD�	�騝�.�2+m�a�@�2�E쨇j�ǈL�͛d�qp�;O�rձ�:�Sˉ>H�O��5$V�ܼ�5�U��}n��RUS��,��[3��,�LT���=���:���+�j��<ޥ0ϑ�'�z�e`u:��I.D��ʝj����Z>ˌ�1W����z���[����-%��\+].l���>��̽��E����[��9�;fT'K:�A�y��Z�����D��NKAw��_/��v��M'p�g�uw%���L7���^�F���j�iq��$xPe�݅)]P��GYU܄爼��1����J�M�7#�2����dt?s��Q�U��OY�3Ɲk7���p�os
�TN5'�H����ド�g�Ãt5`�*�y��;�	O�k�r=e�"�Fn�P�o0��\{��.��L��1�T�B�Y�2k<Ϭ_+�+�[='�e;�"WP�}��3�e(�׀m�Ȳ��P�fgq ��;�����;��]�[�Cu�Mgi��h��)�Y 	}CS�����CM�9�3%%�>�d!#�¶�4MԱ�����\/!1�J�D���!�8'�*�S̙5,TWP\�vŽւWn��u���#T�hE���)����V	��D�
Y�fEÊ\mQYm#[���Q\q\¹k����+����WH������|��b��ig �ڂ퍏z���}�Δ4��+����*L�Su��H�5��.,8oN�ɫ��ƭV�5
1��GN)�g6s'�J��]��7ὦ� >�3�&
|cMc��o-ܽ��C�#`5t�����,��j�?��V	o��f�F{:��	VÅ�̸UD�g�,��y����͚�%�c$�3荊�;��q_�C���B�{���.�'j�H{�z�B�,}6[��<�L�3lym\��la~u�3U��j�����z^QD����؉�}�F)�s�:2���{�+�Z9�RT�����hP��L�+"��0*dfGo�Ҍ�m}U2a��^;(Gh�q	Վl���ê����#�Vk�_�W�it���~�S1��4��UA�E+͡9��u4v
�e�#�,i0�m^3a��вVy�/A��/57�ۤ�r=rڌċ�¡�����(���<�U�Rf`���ǝ�̩�ns�6fʸ���w�����U	���JPNQ���zWt�Ր��]Dr�'���*4��ځ�;�Qnz]��T�3&z͛�x�����;�[E�VǨL� D�P��E�ΛR�������f�g]���}��Y5¶_�q�<����Qt'DtΈs*=�<ʋ���fO��_��Nv��~E��^0�WE\r���d5��(�>
K�����	�����t��zgC�A5�[+����x��w���r.�]tw�p<@�j�	|�2]_�^���`�:X��t��RDqc"�o%+3�E�t��ll���GC�O/#�&oD�.6=*THlV�R�Y�6)��8���cT)9,�)�U�2S�Ɉ�8��r�%C�qa�8"�L�[�!ưf��N�w{��8W�!g�Ñ�jׯ�}zn<p:
��L����n��;�Q+9-���<�ױB�V����k���������Q}�\�7�` �-w�t7�W��%�v����GK��F6j�G�i���-
4F��:�d��F;.u��y��B��7A5g]o'G4����R���`a�]���wM$Sr�9��rܼ�2��&��wE�׃u�u|vkğ�f��Fb�8�(n��EvĜ9At鰍���D��X��c�^Xʚ��4��Z��<۸�V��2�D��0(��9tdE����V~��V��ݹ~���Ŀy�)Ͻ�VK��>^�X��b�EV<G��ԲU��H�W'힨���Ku�kh�ܺb&z5�W5��l�-U̴.�����7* �rF+��M4V����٦ ��>��Q	y�6:3]����H��;-��5���
�b{�����]#b��
�t|:��S_{��n�r!ޑ�ΰ��S[:r���|��3��Z���G��R�==���ʅ�)K#X"ݚ�o�������Q���s�+[=�G�D�ʩ���Ul!��E�NP�Ĳ���#�)ݥ���T�<�."���pG[n��q�!XSC�[
�u	��3���Q��F���"[ٍ�م]p��8u>[:�WGZ�F3�Ua�qu!@����!A/�!yw��]f#eүES�ɵ!E�������L�ʰ%�\�s��F}�/����K�y'�s4�R���l�;4\�l�
z��r[���_���t����'*i�Tɼ7��=b8���y[%1<�<���'i����;,N��O���gt����)j�
e�{�s�w���h�vrQ���s�����p�Jr\�������$�r �R��1�m��&f���j��i�f�����P2�zS�:`���y��l�P�v$;�C�#�r���yJ.�:�"��h�98�;�DC���{�|���X�[�]@�N��Vy�ؐ�8��C
�� �:TT^2��	�h�u��"��y��0�f/%��H�9ӂ,5�'͊�T���.�t�(,:������^u�����G�F��Ij��t��Bu*�m�}�dմfIhE[�DNIs[Ճ/Y�d�m�\(B��,]zwf��vPY��lZn�Q�=��[�dεu$��Y�p�,�#�sV\^�s�;�����
�#8�tUĻ��PC�*����5�%]�c�*)27v�jMQZ�yo����_\5�g� ��c^�ڨc�����!�P����]����1�n����'\M���^R��
H��n����Q�>���xk`��#�܁w(9H��t.���=��Ѿ��[yZ�׽�^����Oc>������W�b�T[����YX<���=Ӝ9Y��h��=�,�~����v�烶\\Nub��]�`[u�%�P8�Jd��`�<����i�7-ZĪX XH.הT�VZ��+�h�9ַˏ#
�:�ӡ�.ڽ�ʕ�vn��И�a��ݞ}Z@.��ȼ��s�����7vm���X����+떣�<%8�c���t>��ײ�Z�~�����D9��&�s�@J��w�{=��/;�5z�´:��w�_��A�y�EB^���$te*S=���E�c��^;�N�-���9\�/p���؃N�A���\J�S�ٷ#P���j.d��-N	l��bä����>�����>��;�
hR�E�p�;̗-�B�9�̅�4P3/5�gt$]r�V��ˣ�j_*'�).&@�/�_j��plj����g0�X���r��ܭ��{+n��1�B2��dcU�T߱Q�4}ߥ�t�����μR��Z�(#g��Q,�oG\�F�>��ܝT���U�= �f2m_��Z<���)��*��Kd�[�s��e��R��k`��S`�N$��=R�����uN^�%gY��z�S�t��S��σ��C޴�`�����Ezy�ONev���y����H�G�E���M���A@�Ks{�a
�t<"`��5g5t�.!� �9˱����1��*`W�U..��e�di�# �g�}���._��8��*�S�B�/.l����|o:Q�ý��ݽ�o!��NnD/u����kq��/�鷽��ڮ�Gl��'j�ϟ'j���ln�t�8!�;,���=�6�Z���C��b���S�,����v�+9��r_��"�z��$I�R���:��O�a��)+��Z�J�Or��Yy�{(�2��Ud=�aQ�c#US��d��]9�^���?[��6s�2��g#��;55B�Hlan�fk§ �'�&�뮜���Z�m��4���m8P}���S9��+�Z3�LX��������-�Řl�n���]��3�Xj:�}JP�ѕ��7^�L��#nr9�q�A�Q4�t����=��'"a#>"v����{sB�Uz���w�n���8.���Ξ�p�'.��՜�*^+q&�
����c�&v>�
ee��Sڡ�(�i�}V\�l?t��ǆ��M2�(h_��:xEG(k�,"�G��*/�g��q<:�\�D���~a�[ځ=s�>!�=�-������] ��_*�7CI�=gυ�nٙ���Ԫ����`H��.힎��Xw�;$j�	ܹ�����cf�To�t��ID/+�$�������Q7�^�K';b�z�t2<�����.6<}Ip5ۍy���\�N��|�hGxZ�ε@�;zN��NvE|�ˉS�i>�S�[�ןf��Dp?lݕx�BH��R+չl�N�T�_j5��[A^H�m�ʋ���=�_uƹd�,���E�w�
���L�����ξ�>�3�����v�n��`T���>�M�D@�:2\c���*ˋ�� ��rs7g.m���w�/4P�0�]Rv�z�⦪+�v�>v:��x��j9ʦs	���ٝ]���cg#QYD$-�>��r�Lfe�A�E��RS�����(�&���004����ь�������'�{ ����9J䢫:yH�SW}m�\N�}E��!G��T�{<r/|پ���28G��jf2$]t�ۼn�K�c�Y\�d?s��uK�pm��Nu���Y5��$�֎L��
蚜K*���Nr	��+ļ5�|���v�M.�N�����ռذ����C*k���,�ᡷ|��6���/XV��c)�ز����sCL�B��+F��"�SuQ�X|k��2s���o��|뢺�{~����Tx"��ʤtx?������$R��q��)msiѵ�[�e�X�_G���N)�*�u���c��P���1tN�����>SsiT4!���*��hմ�oy�(\SIï�f�f����s��*ƫ�l��!g���̊�۶{'N�R+1Z'������G�3w;,ra�������a�5S����[��F2jS���:���X��*O5J�r]����n�Q&e�Ӊ�sTL�ֹ�����j��(��;�ͳ�8C��
����D�	��"qUM�L�D�dV�w��|껺!��qc$l-�=�J+��S��>�{&ۧR��b����
�����3��=���P(�62m�Qfr������\%�\�H�M�u�lk�p�m8+C�˯w�����UH)�� ��<a{O7@�����H,�/�i�TR<�6ì�:�C�L�d�Y���`x�Ru9�i���� ���âhFF�Y����G�@�@�:^��1��]QCf�����c����+:�Sv�E���bq4�T>�'�{�\�+x^�D�
�S~�'��u*,7�'��q��&��|%����}���CW� xG�S;�j��� ���rM��IRy;�4�'�T�P�9��B�c-��,��a�uI�Y<�q��A@QN�d߹��I�*y퓮�HL�r�j�c7r*�:=ݿ(��<l{�2v{ܚf2W�O���ֈ)�
&�Vm ����C��=T*���L�ef!�;�E��H)]�?!�1&�P��z�g�
�鏒���O�4&:�'��؏C���
(t��N�P1&�'�i�d�;�<>�,+
�2w)�s �1��Y��&�R
u���M'�,��a��7tB��4���H,�{;܊m L��Y���l���yG9n#�la�����{7`g�JŚ�y��H)6K�f�d�ߗi�N�������^QOL���*f��ɷ�f�w�H
/�������� �
��p���?�v熷��	΋<�B��w����!�̟�~q'�Qg��&'��q��3:�H>�<�4ý�Ă�-�����SϲE����S�P�OP��O�w.��'���
�'��~'=�q��x|���V�<
D�?x��1o���.�h�[N�3j��aʣ�A�B5[�ٲ0�5`��'���Jm����z�q�ǡ	���=}	�y���@��_u�i{�\�{��(}̚zBқ�j�䄣v�]�up�!|2֝�u����(l��ٵ3~6-�q�V��Z wrBh�ǒ������qj�)u}�4����J��nv�jv8
,CҲ��餕,�7P��M�bj|��Y���;n���Ŗ0s!�)�o*A6���Z�q�3"f������ ռ~c���P�zEG;3x���oN�7ʘ���gn�
��OP�dPޡ���ރ:$�\ǡU��է=O��\��xy�ع�5���3��
l�Q;
Z��{oB�\gQ�QEA��+!x�M���	e��C(Jޛ�W�o���\rZ+���,g<����_�tQ�ֺ��&u7;���!躼x\�Ī<Z�����.#��a�F-	�85M�ڧ�o��p޻)�\K�O���^y�ڵ�x֨��t����Ѧ�qn�:��ci���,�Us�t�>�4P���H�#%1��t}���8�hN>�r�N�7iv�.x�jm�6�]f�q��v��r�Yh|'n1�����������gM��`�����h>�rT�^����s���4ɡ�>bub[f����bͲ�o	�ɵ�X��t�e��96�p�=f��m��RB��FՒ�,�XV����6_$�A���m��l#�� ��+hF�����;0v?|ΰV��n�|�<tFSJ�s��fb����6{������%�5�|��1H���7�7-���-���J�kT|l��7ʯDF.7��bx�t���̱��雃�?wf!w��Ŕ��&�!1v��;M��jȓ��\�<�Q4�NX ��wPCk^e'D�E�MIz�c+�q�K�8Ц�Ⱥ�p=vpQ6��evXi��6�)�92��R��[�|'<D������g���7V&���F-�:��������}.fʮ���{_5k��;�Fr��
������I����"��,��l�;������~�T!0�wCu���i(�M��D�8I7���p�6���W������dmO�(wUC˘��^]MB��p���*����:{��'k��.�X�s��Wj��H�T�W���|�ޱ5��Y���ׂ�q�Ρ��U'��<8��j��|�Y˸m�Un�:4L�4��mݥ$]�E�E5 j7A=J5�mu^��!�M�ԭ�àɕץGWXX2��(�r�ke��^n�s2e�F����)���ͽr���r.�e�th�`K/_�}z��r%�X&������ �O��oE,�U@b��*�M#�9i�F�4��tfx�����E޾'7/��:�5�3��͕
wWjՇ�UE+K��ZInַ���_/߷��^~�h�,	�%H��,��T���i�YYa*)
ŕ++��3*X�YU�Q�E�+�*QB�&0,�+�A`���X&!
�*,AT�Jŋ
�RT�aPDb�EY ����"�i$@�j ���B��
�l�b�PX�����P�ȑH-J�AB4��	l�d+
��`c "MZ�P"$�	R,+%I
¡+ 1�bP��XE�"Œ-B�����b��I��H*5��6����*`(+l�0QK����<��Ϸ��|���9%�Z�׵�Z�s{���@D�yG+��}�u�� c[6+W:{WRp���;�I������|+���hI�mu��H��f?�=�h
)Xk��i�'�9����9�B��V~a��'��<Ն3�J��g�ޅ ��aI�eH>Y�N�Ê�I��`q����4��|H=�.29s�vs�8�R��L����=C~�����"�?yCI
Ü�jm�S�`�ӷH��O�i��<�d�f0�³L����Ag̕<�&*�������U�L͏�����"=qQ�����|�+��Va���;��x��*)=wI���6�'uE �d�_��aS�H(nw�(i��ɉ1*,1�M�����~B��	R��ߏ��j���E|#~ (���;��&�0+8���4��񓩿��G*OP�S����7�B��\�P�T��P<�0�>I�6�;��|Ɏ3}��T��&湅M���`k~ß��"�X�t�$� c�"�>5d�Y:ʜM�3	��!Y7�2j��N�È|�AH}i�*Ɉ
)�vs�|N T�}�&ӌ���!�p�|¾�i1���&��%q�9��������Ͼ���W��E �w��|���X�a�Y��&0:�Vjo�g�*,�Ϙbu!�����Xu�"����$?3~�&ަ2b�s��>I_ bwZ﷯��{���{�zy�C�>f�7����VaY�h����d�5�IUR
|�E=Ag\a���R�3���m�XT���a�m�TY�옛a�b�}�|@��ޘ��#o�5��X'�����bAzw�C�g��b��a�3��i'P�1�ܶ�a�5�)1����lՆ�_�5�§*M����'�^R��q��� LF���+�䦗ɛ컞[���xͤۉ?%���I:����P��<?w�񇺰Ğ{� m+1Xo�͠(�VT�w�
M$�1e�~d�VM3
C�ߺ>q�L "@��?�|�I8f��*���f}�6�i��ꡉ�'������W�O<7p��̕�o\�w�)>C���'�ʁ��k���ҡ_� i�Z���Cl��E&̠��� 8����)�����;�wff���yk��˽%wS��e�M}�SL�u���{�h���f>jM��NiK ���<����|5�I>���z"����u�CWrmw.��+Q�,�B7�g�����%ۺǠ�
a�Z�����p]e���%{�{�c�a�<����Q�P?<��
�Pѿ��x�2c'����J�����Y�M�p�}�l8³���C��Y�������N�GP6��Y�����]�+o����t\�9���o�����N0�
�R�z��Ш�Ձ�Xu���N!���&�ŚN0��n$�������T�l�l6��4���M�a�\0>I_X���ۿ��_RW�Wv0�>�� "���D��*O�~�ݓ�/ԅq0�T�!Y���I�7�b)1�]�`�B�_4�a�Xb���%g��S�@�����8�Ś�:�o��?'Ȥ�1
�?}����?2oVs�H,�ϲ:�*��Z+'�'P+<5g�4��?9�wa����M�}�i��W��;�)4�ɂ<�#��=���0EP����;�/Xt��a과�m �8�e����g�*(s���g�16��Ӽ��A��+
�Sÿ�Ri��d�ʊ$��0�vm'�Vu�s�w͐����1�{A�J�O�U�bW�y�Ms��)���O�UT�����
� ��>Ϲ���!P�}��O~aR{?fͰ�������4�S��M��=Ci�;��m1�2c��&<\�ܾ��%�y11?|6����@Qa��N�����O�V{���E�����I^�.�{��&�^'5a��z�R~�~�s�'̼�~��m��9��B�_rg���� ��`�
�d�_M�{�V�b��B�:��i1������4��|����ɮY��RT����Y'̶βwT�������βT��hS�'�'��>��6���9��"^����9w�ɺ��;>��C�+�;3�
T�Ϙs��Y>�)�/�	<VT6ZG�!ܰ����A`h�3L��ϘTS�
�Ϙbu�~�(m �a����,�
�r#`I*f��I�K�S\�p=1p:=�gL�CH��J�����i8�f0��;��8¾X,�e ���I������T��S�,�;��^R�<��q6ì*~��m�Ɉ|��7���D�?]��Z:lq�W$�JYM�s��W+�<�|N\r�j{@u�T�� ��D�I�eA-.r��gf�#�� M��I�_Q3��|�Fю�����w�QbSަy��Ia�ɤ�a���7�����Λ���Y2T�
��{���s�k!��z x)�O��3�?&!��y��6Ş'Xc3�$�
�r��ٓi�a��z/�I�+1�
����i�+�M����J�]M��u6�@��/#:hA��K�������0d���#�(i��>�O���si�I�%�!�1 �ɹ�r|`��d�{�]�x��]��t�P*T�{�U&�Qf'���>v�L���:Ɂ<��z�n��7y���xT c���@�d�� ���������~fϹ���q����'����O�J�4s��0�QU��S��[�g3cX,C�Vz�3�L�ALgbt5�P�A�����iq�@�*��S���!P�%t�Ϭ�'�+:��w�=����i�m�ܤ�s�T��V �M�޻�F���>)db�z�( L
A�~�]����`y���&0��Mꁌ�>LCF��i ��n�&��uHy�9%b�'bo�$���<>�CĂ�l�s
��:����L��;}KRx��� 	�}�0�$��y3x�d��a��~LN W�Xmwd���=�&�V�M�`i �k~��u
�S~�N�`�B��ԙ�&0�i�^������}��o����vq �x�9��~T� �f�T���üʆ�=e�i���,:¤y������Փ�ON!�1&Щ�'����HVa[�^�@�1��ݾb��{�J-��O;=�M& Q'�M󙴃i�7w'��p8핞���r�$�1���4T1H;�gy��h��+�RW����i�2�V�V}��|z�wC�� >I����I���+�~��m��`o�3L���Y*�C��L@���a�|����ӽɶ3��Cýͤx�e�%H)�h�0Y�?!�*=헗�sT��J�{{vR�)����g����B�{�I����5��s�I�=?SL6��E�?{���ԕ�{��g̕&�����OSL���'�{�M�� �XfPϻ��]�֌'ە~8h���U&ǭ�����Ghf��]u����joX̆Wr|��+OD�wO��\=tw���[��;C��4��^���|:�qv����*��}o��Eh�<	�ka��@��U�+V�x�9D\@<J���,�a�$
ّ��J�ﾪ��}ٞ����8k_�C��!���'䨤-�����z�OMP3��n�$�g%@S�d�*q������
��-�������
�������ޘ��b�p��L�{s��]��>}�>E4ɧI߻��N�S���]�HV!�w���x��Sy~d��'�EIS�
$���ɤ���ܙ�!�B�זN:egP�q<����D�q����ޑ�g)���o~LL�)�?!�󚇬6�=aYӝ�4��+���w��
(T9�4�h�����d���C�_�i�d�)<�g̕:���f)? T��0u�0�����{߹�����Ϳ_M����~3�Xxͦ0��}f�6����y����;��3�8�0��Ϭ��4����p� ��W]��&�Y����I��$���i��_h�l���*I\���r���~�޾�/�����g�J�C���N�'~f$��'���e��a��{�CI�'��_~J�'��*|���xs5��Lf��Xm �ٖ)���*����~���s���~߽9�JɦT���j��4��[f��9�T�OhbC���7��E:���|�T$�
�'��C��B��7=�M�2z����3���ɬ��d $G�vnI�"~�m�w�s���N��Շ�B�4fdZ��!��Xb)+<��Өq@�.�:�gW����+��;�mE������I�y��ϙ<�C�a���u3a�����SYːE���l��}��>d��6~�*�8��� ��<ayM c3���H,��b�QH}<�6ì�:�C��ɟ���6�u�HD}��|㟺�v؟�+�n��&��۲b����a��TC��Èc�����CL8¡�=�sm`Vu���E�ɴ��{�M$�}�O=�9HVa�։� ����}`Dxm�nۓx�5�������E0]�w�6�{@�3�_j��Ă�9܆�l�RT�w�iO̩����`���m�Qd��0�bJ�ݳ��(
)�O��m8�Ri
��������"xuX�"��R�ډ���`�yC�j�UӾ$u�n�����Yɶz�ё�:u!N�.Iʘ�j�oܐ�t�{ՙ-_��0��,(����Ft2椥�s<���΅��`Lv��Ʃ��I��<��o������`��W��X����� x|;�JWɜ��&߹HT?�ڰǬ�Ld���4�d�;���u�
q����H=���d?n��B�y�a�河����"�R�3�,*~C�bLA&|6<*G�U������n�YJ>~wԂ��~�̘���M�	�o�I��c>d�w ~ʰ�+1��N��c%N�p�rmU �Xn^��|��\a�w��!Xm�Lf������r#�7/����^Shj��@?!Q@�����x�C0/�JŞ��0�������l����\a�;�>~�!�����3�J°�u���~`Vi&�����@��VP0`b���No�t� 8'�k,;��,�R��g9��'�T��2~I�Ğ�E��Sl�q����B�h�xm�{a���1+8�+4y�CH�u�:�}�I���2�1�Rs�{sU�>C���z��\B���@�C-��@QJÿ��L@�=C�w�謟f�B�3�2m1�0��d��w�H)��RqYR�{퓻��R{�w�y�}M�gνy���=�~��ޅ`x�Vx�>�3�
�Av�m�a�z��1���a��"�=���
���m��& (���&��@�7S�g�O3�'��L?0��&���Ag̕=翾~���>��}5�z�{�~����I�T����l4��Y�|�ߩ��
�l�gy�Ă�w܇ɴ=B���;����bO����~�V/7E6�I�
f��bO5LE��T�O��]ﶟ��]z_v��s3�$���/)߳ ��*�}���g��f�^2u6~�8�Rz�r��̇Y�����u�I���a�|��m*>�i>d����*A���O=繡��߾�d���4�9wҗ�`Tx>�
���Y⤮�Y1N2�ɿ3	�����}f[8��Xq]$�֟�VL@QN�ӝ���q���Y��'�v���!�
�ɤ�_���Z5}���˭sg���+q���G�1PÝznD@��	&�5�$�YR.�`~݇��f�Y1�Ʋ�S}��>aQ`nyq4Ϙbu!�����,:�M���$?3g�ɷ�������_���W��a|��ڕ{L��Nw�L5l��;�K�R7����>D׀G�*�-�y�|;����3�5�A�O(�T�'�}���ٮ��<q�[o�iN����p�59�A�j���,�n�ىL�$��҈O�m݌����v������=�弛7o9��_� P=1q� ��:!�|ɼ�C�3!X|³��:�q���aRUT��:�"����0ֹ��)
��>�l:¤~Sl>M��
�4�SL:�C���y���z�7����}��|}�����%N���~La���2!�y�&!�hb,4¦�a�s&�u
����P+0���)1����lՆ�_�5�§*M����'�^R�_ڿg��}�������{��7�0״�!Rvn�3�>q'�u�1 ��N����P��<�����x{� m+1Xl�3h
,��5ޘ)4��T6rřl���8�M٤��Ϸ�~����8w{��{�w����v|�PS��I����j�'��9�Ɍ>a_�6����?2W��s!�(��';��'�ʁ�)��=�*��d0+Y]�
g�*)-��_�����^h�}�{�=��t<JϘbmY�I�~a����� ��~�4�:Ɍ�Z���+����	P��&�y�0��
��k!�H,���4��UT��a�'�,ӌ���ys�ߚ~���:w~~�������R�=�0Sl?0��c4���<B���a�b�:����y��6�a��q'P��,���%E��T�l��x��X.����D &<>�O^?�Vݞ�V^����y���]�C�J�Y߸�@Qqs�m8�Rx�MsvO̽�+�a��=B��Y1�$�ě�i��ɭ�6�x�H:��ɴ�� R=P 0&<�#�gjݳ���n����7��~���"�����ͧ���1
�������~dެ;[
�Y=;�GVc%@S��+'�'P+1����'�v��݆�z¿�=��H,񒾞w=�D@��-_,B*f����e�������VT��������s6�Xj��3�4Ͱ����p�M��M���w�<H>�b��E��H)��Rc�4Ɍ<Y���J��7f�z�gY<��;][������=�~��˾��<aY�w�~� ��<��i>IUP4����
�Ag\}>�Xo��C����x��
����L=LCHW��f�
x����O�A�C�bŚLa���N��<σ<��x�����O�����2t���n�YK%�`w#���u<�<rD�.�i~�_�u�%I'K 3ۨ�9g'��]ç9QX<76��5�6N���YGeTs�Ou�����ܞ�Yz�-����ŝUU{Ԏ���� <1��Ƴ�����J����O���(��
���h���a�3�P+Y�bI^�/	��O�6���<��O�I�����?2�@���l=a̤������� �~��I���g�=��)<C��"���`l��@�c9a�� i+8���iE�F��I�RT���(}^�9�{�Gs��5��B;���`7oC���K�l�}�|2�b��4��*�>�ʅR|���`d�K�(Oi�4rlm����h�;�ޠv�i0<><����8�ÄC�)��X��@�p�AQq���̃�LFb��k��+��{@9��G7@��|�]�|/�ƞQ����Ip���8p7:��*�ę�Wp�T��թԨ%(G9�cDLhn��<RDF/O�p����4.M!��7���#c�`;T� -��Fƹv-����X{#�F�T�H��9���7O���~��	���*E)��'!��l����t2)��vy3{#�����&qEb[\o.R�l!��,�۴�x���F�N�͏/x˘�JNK��UA���������м��R�=��<*�!������hx�������U�'���O�!��-�Qщc֑��5,�r��.��=�fwK=��Va(�W]�2�.�Z��Ģ*�ne	�lw�u��N�WP	#����K��8�74t����ݷ�S��aH�5������(��<S�	�fl�1��AFn��Gfd<:�{����v�E�ƹ��nr��,G�lX�j+"(���ga��r��Ì���8IȼuxY�)^f�k�
��!�U0>�D9)�Amɫ��h�Ȧ�"��l��s�"�&Qu>�g��W���R}��z�U0���ؼ�f�i��NP�!1*��p�JՂ��~]7�yf��|��R�������w�aChmV]�=��,��W�`�ӣ�q�����fufK'ݔ��hh�%��#l��F��A�N�D;
�lB����p�)�F5��gQx�6:SO+bw�v6{���նj|���
�t|:�*�����e�_vN�yg��o��^����zA��cc���ѣ��\�[B�Ŋ���tx8~������ή�zs3=�n	S�Y�.=�s���͚α}���Y�P����6���`%캎�g�B_��+�{k㣀�{�֑�C��
�������$��eN4J��p���b��N�dl.�מ�J+��S��8�dߛ�R�Dzg���:���0�t+%7p̜sA��Su��f�����#\�������Yw�p�����w4�foxz�W��#%ctZ6�S;���YG0�]Θ�l��:P�t�i���6��4��E��<�S�Va�8Kְ�H����X�v'�� ���n���Jw����z�>+DT�D)>��E-M��nB����>���̩��qf���jk�1'�Db({��q]����_W/�
�Ji�>4�Ղ�/��7P���j�\Js48�ڳֺ��X�Gr}a�r��91@�ρ��C쇑d��A墖��T��ɽJ�,�'�E�����l�e��2���L�܌�
C���z7
 m`E�*0{����7���B�����x��0��N��@���Ո֫b&Kb���9���g
r���v+s�="�P�Gt��ғ�)ܮ�.R��� 2:�W���Իc�,�3w)s8S�v5�}9�9��R�q0��eAzTD7��];��^HD���ƣ�k���T��u'�T�! z�wg X��'�*%��B��1bRu���ʞ��b��w���8q9tc�1��ך>��c_Tt�h�mm��C.�}t��:�����3B��-�.h�b8� 5n<|�W�;�q{"�xDSf.||�Q�8q�Ϛ�Ҋ���(�e�9�H{���{��	Y�Cb�{vkʔ�Z'���;˱0������S30����K�-C��X��T9V�ĺ�nC�{�X�'�eK�iu�ݶ��Ĩ�1w����[L�o��,daS�MОы�)@����*�Uu� {��Z)\'����gP}��K���jpz��q��^����R�d6&�j _H�n����M����	paXɭ�r�w����F9�l��W�wI�m�L��',��4��4{i8�1J��L*C�E�l��t���y����%l���uܤ�N�P���
B��_��8������V�jTAu�0\�KE�W�%C'9���Q���꼖y�(4vd1��/�%3�^L�D�Q uW^*�.���N=x*�,��oY�˜Z�gu����u� �|n���1Jܗ B�#!p^�p��w������q��oy.������<'ϕc�	�@W��*o��z#~�Dm�}6���w��/*�����st��T1�qK�����S>�#Z��B,����1>����U��Ǭ�tn@����"йp(�܁�+F�e��T]�8����%U��#U][�����:Em�i�d�0T��?y�]�!�)�G@�n�ww�vj��үK=V;!��4Qy��0�1@��yqwrGe�Y���|�f��%@oW���)��5��[v���_~��1�v��ǿ^N��>0mvFT�6�I�飠�[�4�/�q���C� BK+�E7-Iz .���X�hK֋#�%�^��5܄uۧ3.�F䎤��}V���h"2�;��;���4FX��=|nf��mq����)�w�����o�X���*p!ܖ�aٚ����:ۄv#�K�'B�K����bA�&zl]��a"�qH�XT�J�Gvժ�A��%C���Zw;O����ۆ�",���'N\+���:^���rPB���)�^T���rI�I�q�p�2U���U�JB��0w�������Js�{�����?x�و�oa��ڮ#9m���fi�fu-{P�����8G�{�Y�=�H���c3���r���{�φ�:�ν����%�ҁ��ݺ����ւ�vP�)M+i3"�n0([۫H���i����׽�mB�yItE��Uvlb��K���d<�т�V:��T�$r���o:0��x,�g.��-l<$M�]�H�WHO{��h$�l�����!#�r�xt�S9C��J��@r���ꢰ��;׵%:'Y���V�Fh[���N7�o�oj�F%�\ �+Z@�8�޼# 6���ډ=E5���y�
��gaw�g����S}V�08U���彸+^cf�Ȓ��vI���ǘc2�N�wxK�2�fh�&�d�۹��ʻTy�:P����ΏoTeFK]�r{ɰ�z�rbλR�rZ�F�a�J�[��D' �2Օ��m�*����[�NV�m�q��4h�J�{]7X5vq�����awh�X��('��tU__9t+�Xl��W�s~�m�q�Q��6�̨��n+�]3M�����ܚZ�A��lں-������u��%=���k{B�D��� TRV�1(v����Q�lJk:�:t(V�=P�6��D|rx��9�u�5�٢��C��YW�`�&e^
R�� {rx��U�ۼ�z�M.s�.��"��跻sQ��8>vt+4E��n�Yt��K�8%;���;���tyR�itl+:\{�a7�+��A hꮵ>�Z����}�0��A��Lw������t�A�W��5U�7��c�B��������8U:u�,��e�t�]W1X@��)�:��g���=�d��{�ɰ��^��w�\�W&�-��ѳC}�M�K0�<��OuE�wg�=����$g��c�\�+	5���m��5����}��A��+n+g\�UۼT�aui�[p�D��gi��W��3�r^\���z�jE)��P1ۮ�6n��'�u��Ϛ���d=wQЦ{v��෵���e��t�H	�������uޖT��f�����⾖��E���k�P���>#Q@
�)Z�ւ�m!m
�Ԩ��bC��ys*
!e�eQ i+La1
ȡ1H���VL�*0*E�Xe�@�2�"�ԅH���!��d�Ph�	RcKVfP�)&2$�Tť�,+��L�t�
��d@X,��Y++$�XT����[��
�VAE� ���Y��-��$2��)(TL`�$�ELf0Eƒ��+U
�-%nP�F��P+�ɤ���֢�,
 V�%H��F�E1�1,"�R,X+iX��\��M+$�@U}L|�W˲t]704�3*oF��V�;�l����7�}]���t����Mx�l�-���P����6�7'��ۛS�-~���5�3�b�ŷ�2�A�x/���~.���|��<��Ӡ�
ʦ塴�)���������Фc��	�F�1|&`5�s��^��T5[��vz���Q5wԯ�L�V��Pb(b��C H�g��Nk$�X�,� =�6*E�W���<�s��0�+T+��a2�b����.=fL �L��s�{6A٨-P�����N�ި�y�z�:��u;��1`�c*P��m8pF�+E�ņ�_B�g�彑�k��;\��i��5��S,[��>dSnl�F�^�t�nOD7Hsg�L��D,-&�dԖ��F�#7���7�D��k���� ��@p_Ӑ��Xf�]:l��s�O��kC,HV��a��;*��u��@�]> U���L|��Ä8�Â�8w#y4�'P�'��}�f��ٕ�d[����I�Sf��P��N��%.J9�
z�g��*����==������=a�!)���q���噦��&�E/�qU	Y{yuƏ���%��4��{ƣ����}�Z��N�D�ç h*�d�NE7��s�\a�C�"��n��:�(r!�=D ۛ
��1���wiӱG;�:�$�ur\dx87ӓ�{���e������w��en�M��������CcA�ꭈd	��`��aA!��r�[<6W{D�LU���	�.U�U��&���=�2��8(Lt�R+��l��AAk!��둰U��t2)��w+�A���7Od��mY¸�J���0{��z|��|Pn�/���2�����{{�g����[�)�:�O�ˌ��jn�J�y�"<)|y<%'n�!��3��U=2k�I@+ŉQ�#Ԣ�ظ`c�3��b�b<�`�j&�+�B�LR6L2��̴���N��<Ӊo�~���ߩB�Ox�
sfr"��8�h�MB�L�bdWy�k�MɭGe��|^���6��^�,�_���7��_:ظ�S0��ױm�ٮ�R��]n�������jL��ޥ�6)��T
O?�>���P~�����A��Ad֊���28�ն�a��e���;%��AV������5�#nO���"�! �%�}���&̆�TyS�tǝ�Ir��{c�3�Z+z�����"T�j�jU#b�Yt|:���gv?m��7����}�S �{+�M*˫�[.u{�A[��M��+��r΋���<��ɪ��Юw}rCݻ��OC��ۂY�����Nh|;zn��W�N¨�锊>�a�<�Y��w
&�ɼ�M�_]��  <��x=�Ϙ�qs�j><�7#��X��'g��>�E+1s��5���q�*v����b��̳I��܂��o��T,)Kֈ��wn<D<��0��V�w�0^|B�]�� <�⫕l�a�cDʅ��A�	ʽ�S�*"�1�a`e���;$+
ht����ܺL����W160�t'D
��B����Nڬ��i�дl��Fߖ�^���ecb�1�x���:Hc�8ސ�!Z#�V�9�>����߲mHQU9��w�,��c:�\���y�{�y����Zf�V:������0���4�bK�{�~�Efz%m��q���Q�tר�q��d���r�'54��Hl�=�󦆙g���y�L��$�Uɹ�T��6T᳻!�(���I��g���J�*�i�*� *]Y8JTj]��Lqw����r9���<UX�a��t-�Μa�z"����7{ꕦ�����v�B�/�V��d��U�B�W�QRl�r��B"���b�� C�4�"f��\�����P9��wB�42�V���!*���U�jN���������͑�o��"w`��6��7z��V�ʇ�.l��Wgh���IA�{��v�+�h����;!���Ft��oB�z֋y����[�Ի$���u�~�諭��d����ZaI����E�
�3[6�ٱK�9��x>4������h�@؞Q��;
�l��LV*�������qWE��H������#�pT�e�<*�^�q�*���)��}��e���v4x���GH'�������Ɣ,Yj�6�}� SZ���D3}�5��W�Pa�^l���nY�,QU��{�����8q���G�<y�H~��٩�MI͍|Վ� ]]0�^�Qjr�'��k��=���+�7$tB0`.�m�1��o].�T[�N��c+b�i�����]��8��Y��*JL
UT(-��e=�՛�v2��l4�혱1t%#^�Z�=ˮ�1Z��^e7n[0TIVЮy��f�&���~�2���R� [��S���bm(�t�o�iKs�T���0�vo(��}{����z-�zd���x�ɘ蕱�)��;��h
T�o��N.����n�]�|��p�ӽ�N9���XƎT�tS�%ğK��Q�w�[�.<��/Q���-���}W�N%]���8�|���1gh%ײ��B�y��"����5������S;^�^p4l#�:ݸF�׋�fP&�c.���U��Q��X{��A;����Ў�����!v�������sc�R�a���p�R���?��������ibNV����l(���)1�.)�ݞSp9���*q*1C�l�"�?S�ڝi������}���+��<�:\z������q˿utu��\��/�|#Z��B)��M�SsX-��wu�=�0Δ�*�3k�3���GC2�r*.��w!��W��Pu��hUf4��Ԏ���(��@�;9�L9�dQ�'�*n:Cya1���ν����J��gD;��CQ^�hb�;,Q�j/gqצ�t��u�}�&`�l�j.��qD�h~T��0�Ta�sP)���ˉ�̗Ʋ4��4�:�<�R�/&u��ё�k���8Ft�,jFa��Ր��'Z��|Ϣ*(=�!g�g��*���k�\v0NC>�.6,aN�`�1�up���&TX�n��{d^�AP��t��Y��عeJ+u0��oμfj��-a>����4�m�i��#s����b��}����&CR�<T�F,�$ˇe}���Ҩ.�b3�YC���S��*��)��i�.�����bd,�/����7�=�$�:��R��f���+ޑ=���~�UF��y��Rf��g^��ٔ�&3[1�Y��O,ۀ>�L�5�+g������+y�eq5�H��ynF���Ok��8E��F��ȼ*�m�u|<��1�n��&&WtB��9�FV�DŃ#s���*�³ǜ+�r<)�,ｳ2��r��@�έB�.u�_[v�F)�*��u��D���QqC���F=@���:8.5����ѿa�ټ�.Z��ԫ@qڙm�nn_��)>����#�0����6��P�Cw���bgc������W������w�L&������Lf�48�Z�tK���9����tC5Y̲�`��(7!쫑��]�g��>���\���:�$��x+���"�WL�zT!�q¤WL�@�u�k!��\����t0�5�ppG<��V�>��K:���T�A�`�;�Tt�aM��0�\�Yw[ؖyi����w?W(m�Q������x�(]}���D,xR<�;v:�+��hة�5"�o��tz�Cc�J|�`S,G�l�Ȋ~�4k�F���]���q���9�ˊ�nՃci܍�o"!�	�\_��5r��4W �g�)�(n.�\n=����[
��[V彵o����С�L�]2�R2��s<��n%t�.a�ҵ�pE�[Bڄk_Px�W!��
�Y�����Ry�"{s��������
�YQ6�p��������]S'`b ��<9@elP��蛶=��x�q}o)7:���TtZ�O�*��F���n���b��L������fn�=2���	��Ǳ��6�j>�t>Kv�"E�^�Px/���{�,mB�0�0�l1u��k���e�K����렌��9�`�W2Љ����^�̐�c*pCs�l��\!cΨh����]z�⍈�9y�Y5��+ְ�ce{��S��a�Hخp��{��K�N��������ڷee�~�1�܈y�djvzc��W���ؿ6-���;��;�3ӗ����5�Ac�t"�`�JYՌx��x�yՊrUt
��D�>�ug2,P���'\5�z�����c̴��ny����Ȃ��V ˽�bvHF�L�Ot����vvd�3���Z'��	yFWR�����	my�����
�Lsη2\���;ѯI��쉭x�\��F���(b�|�h��؇9J�x�62mHQd�CmG�W��k#�]:|������}�����y/�����+zZ�:��Eb&0,�|���%�+�I1q�G^e��-�s�q5���K��~�¥��(�D�r��8��n�7���V��c����mܮ��� L�=,wr�:n]{R�vxf��Ӎʉ9�Xi�W��M�b��<�ޥNT�����P�}s��^��  |R_�h�MD�\�Ɏ�[����a3�>�d�M�rb� ��Hl�G����c�q��b�����:뚅k/�RѴ���!�(���Ry}��~�lH*��.󩎲��Z#1�=1�5�+�+l�H>�����\_�OV5TùNB���N�<q�	^�=���	7g\~�+z�Ġ�҄c����Q9�����S�W�")�nf+|��ƺ���٧E��]�nup3L&fI�A�r�t���lR�9�ǃ�N��ʹ�V��+1�������<�}��tD'�qC�����D}�H^�Y�Ԏ��R��`�W�KrcU���O1Z5�e����n�Ƌ	�~���X�dTQh�)�3�CJKNWL��<o��7�l�&���y��������f\C�V���^l��(���Kf2|�MT뢯%���`,��g95]VzS�E����̔��������oU�������}�r2bQR�Q�����P��cv��)Bt��1����{����?�Ӆ�ߧ����^�$Y�����Ca�~�;��}��r�"�>Xf�7:��
8���m�/�c��'�7L�G��<6��ɪߏY(e)V�����lA3�����W���b�yz��0,{���^tmT����%;�I/%�4�ׯfhѧ��YO0����]ɼ��g}�  ���5n{�2`}����R.l�(J�5���q����+C�y�S��P�m��}�Y�k.-��Of�0�핞�[V*Q&�q
��k��b��υ?�\}��ʙGn#�.M2in%�V�ȴ&�qS �J-�Kg�������:¿UD�$`s^�J$=�TS�䡚�^��̝�`�!7���:�!B�[3�x�ʛN��j)�Èr�&�[ϼ
)�k�������gc�p�C�h�=�✎��'Y_���M�7,Ϣ/��V��f���{�qB�۰Иܥ`сS���C�PpN<��pv�ʗ�G�k�)U���z�ma9�S�O�Eq��|f!!J��ͻ �`��6��(}au�<����	�\��f�"�I5ɝ�B�T�c&� G$�]G���{�"�آ��<��*}$`�M�7���7	�c����zq�1���WJev"Gd�5�hS�������7L�~_��[F�1Ue�$�q��^��0���e� '�4ӈ������ˉ�̖vv���2���������}"���ә*�|�	׍��Id��Y�V�RWl+�8�g&��iʢƶ�g 6���4Q������Ė3��$Y��r�5䎶��W"/��;8�7�+B������&��ajd|��We����2Wot�@VzrI�䢏}�x m1���)��߀�l^+>�전gIrƤfF�V@���M�c$�}QEnuK�Xc�T[;V�f��}�5����v�X��F���2��9ɕ�8g ���$�R�89�.�X����l�F���3@U�E����l�X�HF�1����E����a���ܮn�h�K6��e��֙�$��ٔ�}���# ��ۛ9F�רHGd���\�o=�=�nt���c3r�08��K��;��(��>|�*�����A��B�6P�ޅ�9�$�����f���[������S��lWXn�Ix
�"�e`я`��y2r�f;u�I�K���,���)u ^2�Gpl�s��R}0�����qcd�V%/��z#\�T��S*/߭��W����!)������&t�i�ûdt\����N�7�#�g�/��P��`xr�E�88A^��21�*�7��W9�qЯD�}���1r̢6�>u�$A�T�H��PP���>��-�9AA��np\����{�b�����Fds�����"���eڰe�y֚�P*]ID-��J����=��P\E>D���ٳ6���ڙ�ypk�a��D�j�v[�g�>�l��P:����9�j8RXج`L��q؏v�ەl�7�F���ײf�^��#7�nw,:��ӱ,��2�ڸxh��$�]�Ǘ{[X-;]�,��f�|]��j�8�/��M�v��Yؘ�*X�]R��W���h�F�f���5"|�]�b��Zm:�˩�ח�<��L��?Qm�Z����s�Q�3Ҭx5M���%M�������y�����X�kE'NQ��]�*"K�vqWU�$B�o2�j�e�Ӯ��vu�&uB+F�C���W�G��i��|3o�]Mn-o��s&[Й���j�v>�(.ƛ�Qz37��s<D�����F�j�ngY��$0���q�X�������J�yɓ�N��@�I2��ţ{��
-t��%/�Ve��Bᝃo��/#�pZ7/�$�s"&`O������(y�ٍ�Xm9)@�0H������+ň�.mV���?�8�6����wU���`�0IoX�#�R@�u�1m.\ҹ�!����W�jT��`�7y۳��ٻ��¤<7�����9A������/@��*�a�|E��"�}�U��3�͠�.
���\�Qj��j9ע�e䈩��n*��p�������p[��ۂ��Xi�#��҉�	1(rۜ�<`�U�Flr�޽{�J�t-�kqM�wd�d	��i[�&���;\��Y����<�0"�9���z����;��՝ǰAK�����8��1B�t�!���`%�W]̞����=��ANV�a����&�1-!�Q��6.d��}�%�x~=��٤f���_��8<�g�������x�G���n�_�;;�^�j5�7��J�؏��U��g	}I(��y���J=�{�آ�#��H����Уw�$���FU�Ym+W|x�Àw����62�|�n��%�������=dlٰ�Y&���iח�x��	N�S;���Gk��X͍�D��[B����s�Z("�CtVv� �l�,[]�K�Q��%s���6�(ڕ�yF��QWr�oR}�������3X
�]��
�iz��.��{�_3�UK�Gw�0S��ܜ�{>8���f��u��0�ǉuC�aoB�/�f-![y6n�����d��*���m(m��N
��X;�y�w���L1�sh��ź��z��Y�Z�^m�`��g_ی�ǪRCy�l�
@0da�_)\"��i]��Ȗ-��4��ŏ�/	J�]nj�ٔS�v�ve�ӎ)��i1�Fb�t�P���kQ�.(����,"p[�j[�fWU����wx�V��k���.g�iڶ�1	�nί����5����Fu_h4A��.�왢q��=�c���eMu�]U���j��7�yX/ݴv�������N��E���H����,Qd�WDUPb"�-���#j�F
J�ۦ��aU�*�0U��@UL� �b��(�#UD`��WHV1Z"*"��h���
�,
����"�FZPQ-*Ѣ�Z ���)"Ȣ�Q`#�e����"�IP��uC2�ZY
�%DQF*�����D��E�QPL�b�E���� �Y++t�Mb ��*�b�)�c*J�J�EPX�,"ʕ*A�Pƫ2��*M3E�V��Ŋ"�����T��I���{���CPc/�u���t�Ӆ;CCY�\�3���QA�γw�|p>��f�b�݇9E�n�� ��\J�?�����>[*���1�:/�,����顐��+�^�-Ԇ��)��}1|����x8�i��%�E[]�A��u/�ձo=j��3�┡��=D<*��xO��c�ơ�^sa�i��N]��;���g��S�G��mgT�o�b�b<�`�u�
�^�~V<��h�Gb+�!yC�.�ø-����(7�9B�ـ���%4�ь��Q�����s$Gu��"�@�c � O�*��b_���'�)�X �}܈���遬�qMvq�˰֝3O����1�=U�ړS�
�a�*�f[�ɨ�ssa0<�{�}�ә�c������+�,�򻝒��k��4Pf�Z6ˆ� �4��+#q�v]��R�np{�Z��
#[��	�5�ښ <:x(7܃J�j�jR6+���7��룓����3hc��p������שw��"^u��	��=����R�;�ŝ�=Ca)�'��n�z�2�����aR��E)gZ���q�!�V)�U�+�7}����������5��h����}f+H+��[2��.8��0�_k�Jͪ�l^�:l99R.6R���-���6Q9Jf���W�#��r��h�ի1�ή�=��^1S$����_8�x�Cy�`ic��z�/��$��_ob@��ׯ�b���y�*�9&���� <��n��L��P���4c��nleR�.Br�mZ��*"�1�ac.�R���8ׄ��q TUH�6h9��p�EО"2�Ԣ��Q��������F�A��4��	ڳ,೭k��[i���J�dXR:b�W>��5����/�z��,�5�-�x�Zuah�(nOW���x<�9�W5H�*��NςS$��=&�u��`,��^�"����\P��� W2�a�g�}cY9R���D�*!C�V��R��:����X̷MmF��"�Jr;�6�6wd;�2�����	~U��� j�W�9E�����oO tQ�~�"� 98\Txˎԫ�Tù��(Р�9ӂ�*ޘy�ά��;�"���z*tF��RrB���Ϫ攔2����pn�(�X�N��Ek����<0#kMX�fIH2.�L�fkf��3�(]�P}
�FMCs8hi��ӧ-L����b��Ƈ�Q���"��>ɖ�MNy�Z��;���T<*�xVw'3��=q���]����{�2��]���a*C��Jʄ�=ؽ�_��O�Z�z�[Vէ�³Di�<�.����sz�{�9޽yi�w'���.۩���xv��fS3���ۯ8�>��|��)�-M]d�6���6ig�<<5�Du+G�5�vL~*�R:ԎÿK�YF1�H,�?���L�~�4�p��7�&��4t��ƛ������U�2�ob��Q�q�����/dQxn$��>����kK�9�wx7[���N��a��m�
/�h#)*���"�P��_E*~�0K��5Ӓ�k���:D%)��������C�''EH��d�W�[l�+^L�]��8��n�vRWs���V�i���F������.��Jٔ�1t�`�ڜ��v�+A3z����#�nOs�ԅ�^��mBuK%�YHr�n+ݡW�@Gզ�+iD-��"����ث��r8���!�b�m�.d'*�n��bf:%lq}UW�`r�I�v	*��E���i*���`[:�Xl�
�s��v9֓�_��2�ʘ^�_�C�����˱�g�F�P�����yО��	`�2y�����n��V+���-��n(+�%����#��Y6��};m��SLR6�U{�7��U�F�W�ʗ�G��s`-��U�m�]c����t�[��3iV�/6�`^=����]7Bf�o�V�����k���$n���s^���Sª�!��"{edTlH����!n����Y19���e��gZ�%�(5ݿ�ûIU��{ө}��	�Q���$���:ye�_����o)�i�i�B?t�hE���Al"6K�DtйP`��no��GC2�"���1g�v�{��[ьUe�v:h�4�R2�R�-u=�xlQ�g�-��4��MQ���7��QBn.�ÁQ�Ӹ��!�;& ��hS���É��X��{w���N��vh��[�WTK�b�YU�wz(��@6����ԯ��E/r|��G���gE��fN�Y��cb���d�#3�ܰ�L8^�Ր��%�.u�Dok���b��U�"a��eL�Ȯ�r���Sdo�˓9�L����鞘i�.��z�����g8uMC]�>�F�����QX�m��~��-����{�����y�s�^f�ɷ,ӛ=�
�n��}�_I2�3^J+�C�FA6���w,��@��9����\jVX�����1i������..]���EXDع|9���,G��C����Qt���V{޻e_�����w�_{X"ݧa�u���Pخ�ݨ���(�"�e ��z<^���M�1��y��`7M�΍�Y;ڜ��6�4�WL���`�;�vd]~�ryM���#��h����%
g��Ս��ǯͰ��x��a����6�&Vm�OM��R"��n�,���w��FI��H�;3U�T�Em��1��n���Ǿ. J�
�Z��+�
{�����d[�������x���\�8z�ѧ�5{}FhÃԨ�uIgO�:Q����̟��7%6#��q��¯Z��oc+����t
�!:!L�C�%�aE�{+�#c\��z;�®��2��&��bN�¡� ڧD7Nd��((Lt�R+���"�GPP@�Y�{�Ȏ��0��_V��ƅ�X�=�����_)� ��6��R@M,h.���C�]��T�'6L��[���1�Ḫ�eVʇr���,4΢!c�0𔝻cqM��T�c���y��t(�ty����L��PUy���p0�^�h��g��.϶Խ��꾤0y�|�9pCu�N��S9Jh-ɩ�h�c!p�O�_1��Au��'ݠ���=*���s��r�?yJ�,};�a�����ڊ���K����Wq{�vi�]I�p�U�ړS�
�P�qWh��uM��ф"�g�ʨ���7D�;��}�a���T[Z�=d�ְm����29��s��e�싔�!d������B��zu��� ��z�Mu����UȺ�<�nup��L�HN^��"���^�֨��cE=��L>��v�(�u���<<�#��y�f�]�|3�u�Y5x�l�6�ɒЊg�t
��5�R6��{��a3��e�uׄmy�&�����##c�.�	��V"���/���{��QӬ׌��ʞ9@�I��\�w?��`?�ha��# �uU��h��/:��f����R�.�zl����Dv	�W?{\�N�[�ڌ�7>دP�E)z��ݸ�X��
��(+v���\�wP�>|B�]��ьUl762�A!9[%Op��ƕ�l����8ϝV�U���\�a��
H�:gS�z.���S9���Os�V�`��/����VLoH�T�\���|���ĭ��>�{C�dw���@b�P��;�=J�x�uCZ�����jG����f�{��F�y;�#�ٕb\+��-#t��`����
�F��PZ��޹#�F�w}K/�A
v�)�.�`e^ð��_���2�x���O��R������i{��}S�E�4�j�-�R��xS�a�3��_F'gD^:6R�sZ�~}�b�x��Yb|a����ˆ��ɀ!B^�ur�l�'u�Y��<0C���;+�h`�����C��ʎ�6�[�Di�uY�ʛۙ�}J�{���b<[�[�tľJ.�,͚��-Ԩq�M��2�{�??2�8e��:��6���J����O ��i�,
&#�2�.���2�**�qc��Uz�a�ߓ��CB���u���q�8�E��"ԏDT���B5�'$+�# 7>����+��E7[zx��		�8����9Lždc��M5SS�E��0z���x�6*NHW��[ZFL�;zfM����1y/^��%DC{�"��\�5u$>0K@�=Ӱ/�7�tV�c�yS��K��C��[�w�����A���p�Uэ�;"���Fy�3C�5b��z�ַW،���Ou3;2�x.�0���̨�����|U�Έq{"�Q�.�O�e����`ϛ�F�����`5�M�aE�3%+��z-H��47����T��ᜯv�ٴ��m8���Ĝ���*���6وV6���j1�M������wϘ�]��^�l�	�R`[��@�lŉ��ExvT+C����wV�4���1�z�d��^�Up6-	�0ӷ}��@֋X�o.x/�+��B��r���d"���T+ӯ��^w���]�햩�;�����a�g!�ٴ&_C9�X����̝v��p�o1����g\[�&.��=��w��X�g�����j}�o�*��Y��Jp["�M���=�F�E��mE��+�D��Υi]v~���%�0޷P���2iKs�ٵ �P�x������>��| �r���[�K����Q�u�˥J$�E)��@��:���Py���^4r�Ӡb��Iq(5�� �^�_��Q�(`�V� <���%c�aE��yN\�K�.�tߓ�u���V�A��}X�w"�0�u|ϏWQk�LP�������}]j���t3:I��M������9'v>�M_I���l�u=�S�L��z7CL�F׼j����}xS,"��W�ְ�"�Kˋ�fC�9� ��Sa\S�4��6*N�@��sGY��F����eA�ѭKBT��T&و�l��Gd���4ċ���+T�Aq�o���qg�7Û����*��D(p���ފ0����"`�>1��9��
�'o�67�2��R���2ܧ�����ד�6�l^;>�2�^Ϋr��Âmud�{C�	��!�R�3�5�����p�EE�[R}R2���aQ�~�ݎ��/�GM�{'{e�a���$�n����G,��h�H�{v'k�`aT�#�t�u�`�e�b)��`��#Տ�qνڞ�/�EK^���\z��,���'�0��O,o2d}�LB����{g� ��9@5�gcP��m�h���=/lvVP(Ʋb}��j�K�_ A��{_��ڼd�Q�n�̗������+	�E��4�m�71	��t�%F+����Cqo�������v���e�26f�Q^���ЬFx�(vU���/Ju�p�z�s7������膪�͛�a�\X�C�v0&�2��Q$M���r1s��D8E�y��\�%���Г)���7�
\�R���8.��b��Cb�۵C�T(�����9�Q/�[Q�-��1茄,OB��-OAR���,���������+x�_��ߏb�N��N?��F2\H��*�LL���eG�롡uOXnJG}>�q�Jw*���J�Xn��@�N�tM��};a͊����gʺ���IX�uP���a�kx�<	Sɹ�ld��-l	�]=�]w1��[�}��֩@��̟c�(!	���*Et�tGPQ׍=�o[Ț;ͨ��H}`zxh����u�s�}��D��=꣧�B�WX}�P�T)�)�u��
����
R@̧����*ˋ��g�b�&
�6TH���d����ѱ,��;	�۴�/�0�yo�P����9�i��D�M����^ˇ^X���(�'M�����;�	ɰ
�^��w���sbݮ����؊��w��qG��K����<�b�Q�a�,�;�,H������}_U{��8�.�}�3�P��2*��{F����T�ov��S,G���CQYJɂ*�̘�I;�՜��ՏH�è�w|�u6t�+i܃��DC�ЧOc�Κ�p���	ϯ޾P�`ex���	�;�׃�!bz7��';���xW��|�A�VSt_M��
E�:�Y}�=e��M�R�#�^h�"� `P�qB��nw�e�yջ[p3I�Q�N;�,E��ن���!\����l�6��/�AV��4Pf�Z6�U�W'�%=b��2�՝[���k(S�<6��8<�
�lXN����t6��V��`�u�b��숣LVr���gJz�R��E�"T!UU���7#��X���KW���Ю���^�p@��4ؕ!gb�]G`T"��A�$R�}�X��qX�8��C��J�%�j�;�
SP(���L�#�Wd�4��8=㖗�5�=+㣀��=g�� ���ԋ~�n0i{���}qewZN}��JTv�*&�Pt�p��Dj��˸���yoX-lX�O�*�a�gd��ΰ�7:�r��4[�.��h���񶒳�{&|�0�GF-T'U#���m���;i���(��^,�p{���i>[�B��=ޭ��&<�r�c�B���g[ظ��/�4_3ņ��h��
��x����[8�5S�|�T��{|�+�n=�ѱ�@���0]� B�r#�,V:9���ٔrotb��t:(�mN�� ,	�YM޳#�}u�Ζ�Nԅv� ܋;te/5������YB�9�N�tN�Y�sILIc�&�q�o����5\}#&�[}1	��-BVF-��>�CoUE��ލ�	ő����ZsE�yf��B"��8�+����RkH<h�ϻ�%]��`P�8��uս�hd�����Sw�nѻaU2�=)�U���-hjܮ���ѣ�͡�_QQ�[.�N�)Gu����ސl�t���~y��1�Gw���m����d�j�f��$��p�v��m]՘$:6�;[����d���)��ª;{�`��+��^J��}\�ٚ�T�0��c�{��^�0'��޽��vo��y=. �7�R�ŭ���<����ފ�,�y��8mhhU��^�o��bh�|��s葫������˴x����v�(bb�q�Wr(�t&k�!*c(s;r��M�!��������Sq+��rc�ҽ�VrK�&��������eє�p�GG���w��ⷨ��r�*��8���%,��S�G
�����製^2f{8K!D��iT�]f����d��
�N��]1Y���m�ohH��+3�r~�r̺/��h�Dmjk�K���iv��5���M�K�>�<y�)�V�M��c���zGW$����Μ����1?�����o,�l,V������+�����kK� ���m �溍'@�p���ƶE@��q��ќ<;R���^�ʼ��%^�x�*f��8x�t�����*7B�+��+w�����'�X[S%�1��(�p3*>ӫq������4��Zx�	u�,�X�;��Y}i.b]�p&47�>�"�s�^�v�K��%�$�i'biiIP���)�S�I�+��Hm�NuBՎ#�b˭��p�%�w"#�m�����}iŝmk⻈��#F�/gҢ�ܖ�.&
ӵ}rsP����Э���h7�s�e����gb�;D��Ѧ�[y��|��f	}Z]r���U%���b����S���CЂ݌�����{^[&	��/� �[��T�s�HD��y�;��>�4!�&�M˜�<-ڡ�K$���x��웕�tش
��`R�{Qdz/m�1"�W����܅|�K��R�Ft:9LKW�����P��{;Ƭ�h:�\����~�Vʕ��ֻms}��
�nޓق��|���2ڰKC��9h�Uł�PDU��Y��.&!��c��ȃ���F%-2�DTQS���DC�J(�eĢ*��#,���4UXċ
5�CGq(����Ⱥ�D�(����)G*E�iT+�Q�ETQ�q�`��U-)�J �W�RV�V�Af��(�\J�X*�Kk��VbJ�[h&Z� �QUq
�խ��-XŊ,X(��+#b�1��b"(� �-�b(��e��PF(bTF1�Hc�TF*�b��DU�Rڢ
�������k0�Ve����PTm�(5��Ʊ��,R*�Ŋ
�Km���+I�E �4K_*���9K7�`�I�{�
���	�y��aj�Ď�y�{'^�&��8��9E�z�9�=��ط���=p��WB��=���^o�yϘ���Y�Js1�c=��K�dXR:b�@B�G
��riW�j��`�F�U��P�2�m�q~&�����;2��3PR�]KΩğmx*
�l�'^<o�V�RE����Erޙ[@���S�z�
}L��~�%χx��r�jTuz�S�3���S�ŉ��G��H�Sy*C�R,h�p�ݐ�:��<��]�]h���Z��~�����T�w��
�BEÀ��EA�e��U�UL;�N���[�����`�eV�}:��sgN�g�*i��`�#\����FFxCs�JNe;�VN��Ⱥhaͬ�ln���Oܪ`���C�5muyS>�����x��͊���\7����"�8�N�F��}5f��M��Q��q@l�&O����
�%�y��t�CV�$Z�`�	��h�����a�����Ft�%Y���c4*+Z>���f5���h��8s�K:�w�jP�(�r���ή��u
�l�.�D;�ǈ�U�Έq}"��}mC�\B���L�Z@Z�c�a��e��ݩ��]�/e+gy,re)��B�{��Q�xCCF����y� �-d����=���tSU��;x���**�;�T�kgP��]�ŅI�6o}�Å����w:���o��	���7�c����y�O�ͿSxo?rb�ݴR6�d=t��+��U/�]^<i�,�V�m~�\�sՏx���:����ϺyX��~lU��	��"v4l�+k���
r���'�y���](�({W��T���L��(iA�٨���\�F�\�=xЉ��\����j��+̦��uK%�:2���(�n�O�@[��bB�wt�ɋ�|���C�@"攷;H�Q��Ē�As���.":'V�XQ�K]9\
�NVl�ʾr� l
X�N$�-H«�p2\�������G{9Sm�1-I���G�K��^f��3�b\�<6���K�T|87�Ճ�?-���E�C�m:�S�'Zo9��rō�U���7�Dn?S��ܥ~4`T�(�ʌ�_utu�W��;��ʵf3/v!�t[�,�+��֩�ЊJ�z���F��+�x0����֕�����oi��츣��P}qt��a��(=T�Cq5 `i�6�8�B�N����Q�}~xy�&�M� i�Oc�P����m�(6����[96�\���Q ��N�"**�Cv�fI@�5�q�������z� ��¹��D���#U�fo;�*|Gv&>��'fb���'	���&@�:��VMXHnE��˔��Nޜ��ʨ����X��j5���_e�@�*��&��`�HC�kl����{��IK���k#�@�[ܨ�{��:�� �t���׎��Q�[�ފ0��@:�"`��4Շ1�
}�{κy��9��0j�%����g��F�f+;>���fu[�0$f]Y�(Ĩ
���=-��[��I�E�}QKEmI�d`���J27v; �1�˫���>��p��uu�`����b��7M2}^ڷY+��I���o�?y����3���z�����$3��f!�|}�˽�򾅼�)&g�����{iՏ���n���n�[���Ӂ��ô/s��Dk�R�N��7�,��t;'cEO�D��r4�1s��:B�B��8�`,����@NQ���s
T�RްE��vXz1N�R�}����BʋM�Ù0p�U�C�ƌz�3��8P�l����+�
{���n�re?E�Y�#f]�m��-`���х.,P��:�3�J=^�P����{׵&-�& )J�Q�~ܘmM�5�K��̦m`���k���P5r�}���	�/Fn����3�}��~5��G{�hEA\�G�$&bC��gha�؛���vnT��n�v�S4�ۡؔ��z�	b��3b�GzFܘ0���k�T�y).����N��N��	���[�&
U��)=�>Σ�9�`xr�EÃ���bY@�u��_N���Kb�El�\s}5�:�T�H��2F?R���ND����ȵ �c��Mԝ�JROo��*C�֎�ˑ�T��r��jLޚ2\�J$�z=>Hi�7���1j~�줞��{�c�x��]6L@�'2�[�W�
�^M�w�"6��3�]{ⵕ�u]�|�r�*v���y�P毙E�q�h(9�&[�������b���o�[��yg{:���^��#X4:F��5ߗ�6t����}�����P�CM7�q�;�z&+8nÞ�,�x|�~�U��}a�Pe[����uC+	
�f^�\�н&.=�f5��ױm�ٮ�pEԟG�S@�I�N@*�\8��@�}���A��z��q�ޚ�#.��	��r�h�sd���L�Њg�t
��d��g_�30�U�+���f�K��4��A��Qռ�Lи��#*k�ñ$6Gu��u\;}�N�M�=����Sy�X��HMެ]��V@�ݬ�ވp0h)�I�����y�[aȬ8������M�"���u����]0����n���w�*�괪_[���uZdole	������+�{�ލq�vq��w��oD���hwr��l�l*��J�]N@d\��P�\`�P�_i�V�>�;_w�v �]����9.�R�WS���qa!gb�uu�ʃ\�b�
�P%K��[n�Ƕ.F��˾��ݷ�+�o5UV���T�WXn�&������_�1t�������5�=+���hr[.��R��L^�B���#�.�*P��5ӊ�%��=Q���A�\��h[#;h<�)�oS�Po���_D�t'3��X%Ӎ2-H�1z�!
�3�^������Z����mʭ�C�,�&܅�k!�ߑ�veY��Ps������x���^|<�c�����\@��,�r}\Ȼ�] ���\�vV<U�;L�ϯY9S~���t�]�4F����{6�bV���b=�)�CJ��H<��ea�9��:�b�e�iz�H#!+ԥ:�ę�;�C�CbGHQ1�CmE�.�p�� ^7�+h��+9�D��q��Y�\�.���c�:��N�ӭ����y�~yk�S�����,�^f����QB�i�>�u��߱�8��R���f�޺�Us
�CFJIv�����0�*�w+������;�c�Kªwk �(��
]/�h<��:BۙG���`
s�W�;j	�nޮ�[�\�ߑ��QW]igr���R��_�廒}Q��X�R̜�m��V�L��<.k3��~�@>���s��@�F���x�;�QO�~�v&R���ѽ�ጕ���Ql�&Z�58
�$��(=�q���gv��ι�������F{:��/�#���t)e�v}%���u�WG�K�|��(���]�4��b��۷����U���HTC�V��e^l��-U�Yv�%�9��"���2;�d��I�mm��[�[v^�RU���jx:ӝ&kX5a,K�R;ugc�R����/�V��,�F��>n��
��w076o��<4�Tl�(-�@�x��:p;e���9]˸�^ä�x�
ָ=�>X�����(j�{K��j�b�|F������ǫ�3�Z�����D�����H<��}�+�M�JB_DW��L��Kh<�>�\}�xgyԘ�|�H)ҋs�[<e�c�i;�/6�[�:oW/+��=ƃ�7s �b�My���@�%μ�
�[3эU�ٍ�U���j�6���.���%����K����1"�q��Z\����7z�s8��!���.9!C���+ ↃVJ�d�?):�:ˀ:/��X�œ��n��=����H�d�s���<fI!.�.n���]eVen�gv��u�~���O[�5�-�Q9��=}=!B1*��%Dul(��yI��p�]��>�Oj\[��Y��Iʁ�ݷyS�ъ>���q�	��U5���0�T�Z�&��������Z�v��QƖ_��L�mS١�LF�
�}36��$GMT<���Enݸ{a)����ܜ}C��GwȨ��w!ۚ03��¸��S�$,0R���ei���j�lOhKl�H�"���NtG@�n�w0Kev"Gd���4�..p�MWm�/Z'��mk�S��n�V�������P:C�Da-͍�XT��B&O�Ɩg�OΔ���;w�8��V����u���K?k���j�).4���G�>[HEgU�cFaƜtp���1���X����Q�&�v2Hg��[S02)g��g0���l��u�g!��i�jᘡfB��B�,�Op�5S�ŌO(��>P��#\��s�u�k	�An�-�vv�U���wv{��g���@yz|�Ȼذ�+�[��f�#fi(�i|Xb���=xڰ��k.b�0�������8.����E�<�ѕi���q�6�>��Pغe�/f�����h{�vP����{�X}�s�7��nz���)��!��]ǀ�Su��r*�fٰN�G ԙ�\�����%����ѩR��f�R�=�'�����꬜����G���q���7�,��#a��լ�h>2���,�^O٤�^(��ά�>r�X� c�E�lZ�r�v�)w�n�v�F)�T6+�)m���RA��<����u��vfĵ��(�;(+�4c��3���
e���[ S��#s�=;�rZG��1��k�l�)����Ey�
\]	�}U�`�(�����|%�|t�Ȟ�߀�|�]\��s��ʸ\����\-�v."c[�sMEtLb�����t�������٢c�iw:�/SPdQ�ć�]�>���\�j�	[�2F?R����>"�{rHz ѻ;��==��������!����*�(�g���9:8hp�pcƕ(�[��\��r8���Kڞ�c)7/�aMZ��U�ld�
Rs)ż�ĉP�\_��-�z���70w��T8m��¸P#�.r����5j�F��������T�m2��L� q'���OmC��2�_^�M��`ݵ8����F\��0����"�Ճ�̍ީ��"=�h�c���zN�X����h+"^NBNm�hpE<4��A�:���.`�a�.=����f�6��ǝY��o�寀;���W����볲�9�gAat�X�?X&�H'b���^Pw�C㥾�/vE]3��.on&M�v�1��<��?�zs艞���t������dՉQ�j�d�X��M�aI�ī�|�-+�E�]b��W)ȓt���.=iT�{<r/[7�Ox:���>K�Ot��}>U��)�Y�Y���)힨���u�j���b�C�c L���ɬuy&�rd��P�'�tLj�{�&g��������T�#��f��FK� �����o6w��n�����-w�;tUN���������-��.���`T�|.hi\!ت���.���:�Ǣ�`��mv^dg^��rWq��;�;�3���;]GT(��s킃��"���j��j�]u��b<�"� �����Þ�)�u�+�7}<���+�3���ʎ!9Y�Ղ�k�MB�mG:K�Fy�qvO�����{��d�aM�>N��3��]J!b��q��Τ��wW�16ra��aW\=4=�.��;�cX�{d�q�E�����;���LX�B��Ⱦ��b6X��^(�62mHQ`Y盿.u�+��P��s���/�=�`���n�Pw��sݲ���z~wu�0� Y� �jj ��,畸%v�0�s���f�Wc,nC#��i#b��P�[����u�Ӹ˨	kE�g���>�a�'��[�7���3FӚ$��9dTz��'�das����r��?{�3^��*�7�u@ٸv&�"��%ι˝�U#��&{g׬��Ё'99�t	�/�5�#�QA���'��=�<顥K\$[ƥeb�0ף�[����@�~�z��H�����5U���lH>TLD��FP�p�g
����\p��\�x��)\�Wp��_y���٘��9Pp�v�N��=S`+�R�k�RrB�����o��pf�,����5�q~�]ϵP��{Ȇ� ��k�I����h:E0z���r�n��*���^��z`1���PT�2j��t��t1��I�d�j*�O��SlA`�Jޮ��C{��ゥ#,��E[���GP�k�պ��,��Ȩ��D\m���Ig{N�K%���=,c;�:j4V�۪����>ː��1� �.�D;�+q��''!VH�bS9ܣ2�^�PvE7��O�1���I���Xk`�d(�4���;����t��t��RG�����<������y�t
�g!�''}R*-�'�±�[���in�V��l�y.9G��y�ۼ��NP�Z,d��ܲ�l�z��7�*���8=hE�ӐكY��Y:�rCn�_�ol�F������S��+��2�1�u���7�_U��/�E+�2�p�N�"��-N|@�'<��}�+�k�[qwM���RM�`U��H�mZ.���4uFA��'��b;�8�:d�Yu�#�=�f��.�
�jEo83��{�u;�a
B��`� �v�l�9�k(��F��麌+��������W-�RPv�V��Z�)���n}o���/�����+i'NX�'a�JwQt��ֿm<�w�������c�Pݼ�8��/I��ZVh�}�[�E����VGQ����ѵ�z�Ǚ����D��۶K�"��t՛�4j�ɸ1��h²��t��T�h#۵���M��f����b6�U��z�ԥ-e�p�1�Z���#,;�u�MLn�[�;��#�.l�eut���[�w�M����=�[Yp�J���Ɋ�ѷR�gP���T+uo���TF��1S���C��9=��2l�ɃO%+��#�*���c,`�b�����W��}�oE�ph7iv���<1��4� ��j��:���qlJV҉f���w�����v �[ݴ6GU���Md��a�������p��b�,0jhxuwɈ7q-/��M={�wZ��������w��U˒�Ζ>ΊO��w<ī �7U��j���vrov-��L��Ku�Yf���s���D`���tD���A�PЂά�˷j,�2l����t�5��Eu�O϶�]Pú65�fA��",�S�r�2��o�\�=&c<z�3蚡�b��V�DӤ��k�O��6�uq�B�q�͹w��͹�t�MM�=,wsN� fG�}+n�������+�Rn� \v3��v�0�����j	��
���*��|*��WZ�X��X-֢4p�hC�m@̕�ݫ�ՙ�$�[GY�gN�>:����J@*�7yRoJ͹�[C78\�Ӯھ�E�꼽8+P��T��8�8c��҆d��`�D���N&���3||�B�HQuq3��BI�b)�v�[��il�35�|���gM���=���B������d���Y���CE��00��pB|�c��7Q�w�X.� *�/���O��=ڳ3MƎ�Si�a川�fC]���uXp�V:�6�u��^�ٴڀ��Ot̷7]���&���փSkget#yh�8t��y[�N�{��� �p��H�5�@����q�:&SRK�]Dw�����-�+u����p����!ױ�����K���2ve�E=]-�o��`��J��6��E*�kN����dW��y�Ư����z����Z���{S4uz���'0f}��"0An4DE"(	�.Y�dp�QE\�8���E����b�Ql����D�D��9B�A-*
h�-lc��;lDU�(2"�"��Dt� �UIZ�ADU-��UTX�`�
��EEU�V�DTDDQV(A�U�cV*������+mP�QEUQ"��U1�X�"""��b�Z��
��b��T��������cP�����P������UQX�U�b0U��XƴF
��1*,2ш�Tb��F#QI�R�� �$F(���#��*Զ�X�UA�TcYjR�¥H�j[�V��Р�V�EX�E�ww�������c�'rW9)�Do�=��[{r*��\Ok��5��f��fC)#���wf=A��c蟧��Y��Bd�z����_���YQnYt��7���w.��J�-%��
�T�=�p�(Cwq���S��yF�^oDj��o������:�y���<�[/=%�zgo^^�;�p![�LN�� N��c��@���b��o��q*[���g	���Ê�(�0�i�{bܱF��N��;ݫSHotlK�(�� ��
j�(�|Z�~�G�TS�|���ζg��0��}v�y�I�����4}���/���(p]X��~�|87CV���}��9:���EE�{��O.�5HFX�@v5��M�H�P�6}���u��*Q���C�x�Fp�K�1���7�}�j%��-뇴]K��#�'B�/&� R3@l �36�i�^���������j顁�l�@u�C2�Qv*��n&��tT����{��%�I
6f�u���}gY��,�*�R��.
���P��;�'͔!�H옂�W��g�i�;/��pw��̡���qtx�sd�u�t���߷��!~T��B&2kdwb�S�����x-�޺�`����
M�4�Hg�12YogZ��m�+�?}�g�D���\��ހ�^�
h�!�O!���	$���W$U,cW�eWV	 �Ӟ�u�J��c%��z#���z�=����X�w�c7���W·����M�3{Z���t�T
�m")w!��RŘ}tՌ��V2����Z��S��:=�
�`��!!����8{�jՊ����t�>_ G����JFAV	�y��"�6Ed<��3�l�[�q���Wl�eE����86E��{�2}�_�Ȓ�R���Y�'=�b�;�ƫX��������� ��>Vw�~򾅼�)&lFF��J+�_2�F�Ʒ��~S�5�:����h��}�R�*!�^����2ˋ�C�v3ɡ�;�z�`�lZGD7���������0T��F.|ghX�\�.k`�UT��)z��'a���b��T(�f�Wy+�TQz�Ĭ	p�P�W�'P�ZF�5cJ��]�}�EtPJ�9�q�������}p�)_��6�:1��T5��<T!�;syչ8�L�
[ڵǾ{��=����.�t���^CB��(Ɂ����+�0k�.�յʥU?aM�u;/����>�6��ۍ���]�N�£Y�f�5E첄�J��U�6�}X�OgdWY�wE�s�܎�_.HN]�Z'��S��m$��\��+����]�^]Y�F�2g5 򝙐mlz;����Bwб��ب+���؆hǺ8oR�ta���z�h@�Ӌq���������9ܦ�68�Г8q;t�+�������fA�% �O'���W9���ᗧ����!�82��e���Q$.�IO^�q{���GjGV˝��[��T�8�Ѵ�����ьU�W�p��3mN�B��Y�`��H8�(k>��WW��m�x�U��>��u�i�=��;yؼ!���dC�rZ���B*�Ț�w꼡s���C�V��5�N�+&^o�׋ڽ�ڰ��>�u�d����EPhlק0�덍�(�+��;�5�s�7Im�!C.��F&�������>��:Q�~V���m�p��=��~ջ���DcC/Pj�?&Vnk��¼��OL����n���xC�f7i��1�е�4F���:���լKI���m���6�����B �l���WR \����s��Vb7��0�aə�����,��ĺ1�#tF�+��w�YD�]�V�A�^vv�>�0�b�
�bW��s��$��֕Zm�浩fP��D���$rt��|Ck���$�vn��9���0�>�\��Lǵ��v>X�S�[be]tgV!��p |�Q]�Z��՟#��v,�����P��v+��S���2����{be�}�7��_j�J�t�ߡ�R������4E���/�z3�anOn�^�y�;�W�/�]�jq����S����//A|�U������ѣ\�u<�l�+U�q�m"=�F5rE�e^�ʙ��{j�psCYv�y��k�9��h��Daz��t��Z�OqgLѤdػ�y��ͩ|ѐk�Poΐ�G�:N"a�����<H�?S�A� ��~���>�G���i�)8%P0�����n��Êy���Qv2�խE�*2�����!��M �(k3Yj��/�y����	�Ţ@��
����m����p�FM42��ͭ���k�nҝ���e������D�J�;�P�c��d� �}M�&d��Fz0�s���brwMq�츝S;N��[X`:�l̭�L1r��s��NO6)�CQ�rža2^�V�$s���=*1OS�=^i�NFT,]�����~�q��x���-{�Im),i�,k/@�S�KZ�kS�ݽ)fD��=��E�ơ���lc"wq_����t���{:���R�2��@��{�JK��v�����6���S�U�:o.P�hY(<";_0�]@1���m�@��5���v������2�c�'�k����ۮ���'�o��Pz��(��a����[ٮ���GyX�lU���w��Q��#SY��\cUAՎU�w�;}�jݲی�Ļk���PvQ��F
�S6�|u��x?Jl��E���iv�O|�j�,w���(�˾{�&{%O7:�3��ãH�:���Mޕڅm�ϊ�mZW��D&��,��1uV0��ls�#GP���G��ej�	z�ͥ�*�]qZK�b�E�a��2�K���A
�����p�SV�Ò��k(����b�)�{k���H�>m�?<^�DUtb�Q��l�<��|��� :�X�#�I�0J�2;N 8ю�u��[��)�n�A
�v��׊���Y��/�d�7�/{	ѫ�Y5i �MFŵI���1�y�����D��-��aT�c��v��.\*���}�J�$ꑯ�r㻥Y\ȗ�֙�}i�)(��}#m���[�cb�F+�//�_h߻�#�n�p}L���)۰���'ȹf�,NGEHdD�e^��/�dN�3�l�G�#�ݧM���k�Vj��ͳo'{F&_!��to&���U�nh*�M�����At�U��s;�wΘ����Y�f�� r��\"��gӻ���*��{Bެ���UK�y���ׇ8��p&v��qO�U�f��~�uv�DX=5SkP�cA{r������+�w�X嵉���j��������IC�%����fW�q3��?OF(�R^cr�+E�z�{��j�lhJ/l����6""8���8Ԏ�Z�.�ج�}s�1փx��e��f�Mu-*q9��u���C�C�! p�ڰgZ���A�~�L���C�DUv���Sw;��jU�� Ԙ�ufy������r��E�Y��U�FQ�w���b��O��l���#�q�ʍby��:V��	S?s{G&e��ۗˣ��ΰq�#Yn��|�k��Wz>�
N���BP�#µ~�.�l�m��(���k����T;�Ub5�x���]7�%�����YO.�|�hE�%��ջ��J�C�xH��-��T5�i���$�#yz���h������w��\��2�кk� ��@Nb�l��8�]N�9������DYz�u�_r{
ޙV��|ۊ���x8d��n�+���l_���sȘZ�Í��*��D��n�Ju"{5D(�ܲ��a�9k�O'@o�W�#����F����\L�m�@0>�.��y�'����Iu�fmd��U�5��|��ֹ�w(Q�����ی3��/����9+r�3Ӷ!`h8�(k�²�*ۚ:U:��-L��[�ı(7wj'�A�h2!�>j*i��߽��3Q�ғ|���t�|	t�5�̶3OQ���}��7�Ձ��>j��A���Ϊ�B_1q��Ouڠb�ȡGz�Iz�ג����b5�U�#�<��e�����ge`;<o��5��x�+�+�i�K��|ہ�oy��-��c0fS�A�ܤOL��$����T(�V�E;x�N��)��k��rk0�T��w�v�cV��n���y�Z�]�7I퍤(�l_-��ճ�\���}w�F;�Np{��"�cf��b�����>ƅe��z�+�UԦ��vu��.�ы���n+�����.�)��ZF ��R�#cVOm]�8]���'��R�����N���G �^��8};V�m��(>���mE�@-���P���B�׋����εл���)�\U�2E�u�����H�Z���[w˞��ځdcI[��>�\�����P��p��s�o./OI	;����P$n��_.�����\!��aOB�s�Ku��].bs��h���P�Y��m.��a�\�3{�^T�*��a_T�F���{Tg\�Lv���[��z2�����z/5�#�s�·7*���2%(���ҳ�8����m�|��!��!l��/��˰�����Փ~ԕ����Dypir�F8f��j|Q�l�2tn`;��M����ޠZ��NB�86��*�
�wNpu�뇒*�����5Yہ![XUI� s5w����.�\Ei���WϛP[�o�՚J����-=�E'�FFZ"�8���^�e_X��8�5�p��(E����s�OD�H8�CY�v�ޅwa��\P+��~����5Ք�>ފm��mC�CQ�Mk]�B�>
!��o��:���}JZ�J�h�9M���A����o�r���.<���i�\�������%����U?]7G�Hg��%�����"�YsT��%��-�S�O�M	�*�c�v���Ƅ��sHj�P��3���b�>��ef�爵�ؽ >jwJ�ʠ[�7����2�ߎ��_�{m2�y�S���������R�xC`�l�]w��&�qU�\�r�����:��25�w�[.s�R[\�އauUBDF��5�k\r�)B�%Ճ�Ʈ;A�ciq�!6ՇK}u�m��»J����ib�$p�
��ٗOdr6�AZ��ugJm�&���@i ���w�@T�Ǉ]<w�y��e\�J�զ�9�=�۩�+�ͦ���#�kyˠ�Z/�;�ZFV�vgg]e���{p;�I��s
�d�UU�{�ΞPw���5F���F�~�B�H��7z:>�n�w�i^`m� �|t�Sދvk�[Ѱ���D��<��ej�K�C�o����EB��U�76�i��m�v$gCl˵.+�4*�R�1څI9
m�1[a��v[mD��k������g$�i��װ��Wn.��۔�pܼf_&��,COs��H�����g��>�
ls�AQ�p����<�y\p�(t��&120e"0:dr�D�mđ���Xq'��1yy�a�y���r�i��_]ùp�V�E7i�Sh:�k��S�n�L�xe��붃�4H�5��Ro=m��Q�SdoE!ӗ9�6���k��HqV!�|2���|"��gӻ����k��T�������>S�C�t_��Ok��L�Q\>6�lק0��x�ލ����i�V��6'j���g��ܥl�����Ҁ�6YC��˛Iڌ*諀�N`�W���	�e�����dj)6ܝl.�.��\G(���惎r� �}�Or/�j§Jĕ�Vƀ��M���
[Z��$�KGF�Ǐ^���&���Ć	�ܡ�f!�E�֤��|�
(���}����s���7Ha�T��B���Zs��s�`3��$��KӴ2�������6�3���i���o ƹnp�2t��k#tK��P��K6�E2J�Eؾ��H��(db����[5W^n��1R	m^�΍l�k�HU�s���/疲��4���UΕ6��Vn�ރ�婷׷���W"�o�*=�ƥ^����r��(e-�>�XtFGi����(q��AR��{zɈp
o8C[R>i��B��aU��gYȎ�ntڜ専��7Zx!�:�Ū��(����C�����f��L���O��<��1Q����~����d����pvg��칽Z���ؠ��cãu:�uV�A�E�e+���q�4�v���o����h��7è��:	�M�|�ZrM�F��i�e�D��	���k���@U8�r�FU�s������#�|A�Z��5�*"��u�����=x�V��j��҆$���p孧�1x�K��RAQ�1�u1%�O6(�
�mM|n�bs�]��=�o�hvF�G���窺��!ܯj�f�rƳ�j��I�;M	Jb�h�[��ڞ�k�oN��D�i�����μ��q������{)l�(�2����:�.����Vŕ�j�!�Z/YL}���;����E]����wT,�����*>���3�\ӕ��U��z�L�m�����G��7��ooc�ɷCw����PYŮ�*+f�X�i��V���g{�Pr��Z<�s��YZ�m���%��-} �1s8�|)����P"3p�1]om�~����Hy�P\x��c³#�9Eli�eW���R�t����Gq�Z1�j��y�Vhe֊D�AU��^��p��y�$'��}۷��R�Ҿu� ��Dܰ�,.!�
JгF~��p����C���C��"�a���`�R㮃p�(��f�!�ٛ���R��'�e���T�[�5�lK���[��ud��dk�@�.V��i�݊���*��/x�
Yu\���uF��Q��^�M�9���a��B�m#Nr��� ������@�>̾;��5%�MLe4*��F|��\��0v�<�w8p���%�J�V�Y'P��}9˟v�ɪ`d�'y��Ð�{͓�
1�W�V5GWX��yI��DUô�q��ږŜ~P����jgsN7��wZ��&+��A�c�''���Opɫ�x1�)��ʇ���,e�g�k��:H2w�y.'s��\�ҷ�~���ǺjE����QbZ�X�KiH��"��K��\A��QDDFA�J��V5��E����]%UQVV�c#iTq�"+m��(��T��X���fZ���+b*F��(�V1�R�b�E#�*�QTX���X,R1���X��īDDV2ZUT�,��Z("�#QEDUT�,
*,c"��AUX�
�b1T��A`騊�V *�,D�����
ر ��d�
E���R�**���DEb"�ES�R,�(�"���X�2+`�V��H��QA`�TX+�U@D�aZ ��m1�5�*P\eV0ST�115l��#VU��,+J	RJ��EEUF*�`�)mUQ7�ǹ�>��e��~�gOm�&�M�t�8�4b��,��p��K�}Ҥ�Y�I1|[���L�G����oV'n���U}�8��^�=Q����~{+~D��js���x�����¤�X������8�Emr��ծ�#2�%O��Z�j�Ͷ�n59��o�roCS���i�t��d���}s�ZF �֋�[q�xaL��Y�Q����k�m��~�ͨ)�U��X�k@����'�S}{%��ԡMw;�pʸ���Ok
^�������GZګ�X/�MlCݐ��.3��Y��P�zЬ`g8�ڷbe+
z+��������g`���'$�e����Ƒ�E��}d�)Gq�}����$6̰�wؼ�!�vԙS�Y�8o;��l�����'t�p;�������&�2mű�F��o���;�瘫�>�ۙw-�ڴa���`�f^__�9<"�ұ6�j�پ�}�*ڐ�-��6�:N"D=x2V�2�5s�u��C��_�� �:�Ի�����rw��6���e�*��J�Z�\\:Eu���"9u��<k3 -"30�Z�F��nOZv�_Yj6��1(DźMw*GD���k>��2ú��0�i]��#{�KHT�b���%��]hh�)-��䤋�)��4�~�>��߱Fk-X������Ѵ�mr��`9���^�s���|����;`�&�A�J�p��ʶ�&��'1���kr8U�cl�O��5E!�4�7���QSM�hk>��{j�9Uѣ�TH�
�p�־K�U����4%��c}��T�z�1�W�q��Y�+'��Wg�t����y��h�z��.�-+��ܹ���R�T����[�m_��V�J������ ��]!�cB���;��+��:-X�=�-����;ڢlPl^����.�)\n��1�������d[�(ߗ�.+����&��^��/|�^�6ڷb���΍;�ć��v"J��b�Ry���n��fv,�.���}�.*�b�Uc����ugD�u�������P<��+�
z1��:X���)_d���}%�� �4�:c�L���+����^�}+���M����[yD�L�T�WC!sI��4��ć@O����tɡ�W{i���ˮ��"���ص��y$��-���I5!n��p�btF�{�v̄��Nlg%Ou� s�`�!�'� 	:��p��! �M]-W�����N8�}j��<gq��2���+�=�qݐ��ᣳ�p*���<���U���y�#/�_l�Db~�jc�E��Q��#��omN�.(c�^��� #�/]�ҸL�Sb��nwc"���۵��jE�����i�RQ@7�Hm�C�D��{�de��%�wf��J,]�ܤ��G�;�L�>��A�
�5#-H{]��9A����yi�Z�t��=���igC.�F|�lz$�A�J�jȞ��f�mY��x�OGU�C��*��#z)�n*�h2�Z��\�cۚ]lA�n��
����:�W�npU���P�A���/V�7\vM������?��z��f�%^�S��׍iZO"�u���lMl2]�P0ԋ�YZ������kp����+������u���xE���ۡ��4���v�2��D 'ú�̾�حn�n��Xވz/y���F�k�;]��[���om2�L���x�� ��[*�ó�)6V��R��u~Uu���m�I��c!����5�ޞ�26���BY9N�3t�������+��|��!�G�ݱ�=ᬬ��}T^\6�|mcc���g_��7,OlI��G��&�;o_��a��^�a�7�{Y��z(��n���곁���q<�:D\���3�j݆[>s���.�oz"9T�J�O=����/i�����3�`ζ}s��m.�)�m�*��((Q�R��Zq�:��tyw�~}vԮ�(�E�n�w�q��|Qh�̼9qK^�U�w�u�Oi�S�Alr���N��4��#=������0��̥��;�>h���cW'ͳ.���?,CB�ίKF�*b֕��N����ULaM��h���W��i�V?:�i4�K�zj�����vk��&d`�Ϸt�s2��:����A��;����|��$���6P��H�r�dcv.Wy�kg�=>�R���6؅�܍�i<^���W[:��рY{y��u�G�82����7�t�"�uj�-nrљ�Pc:����]�ǝ�ުMYG����Ӡx#�Z�@ʬ�OhM�ԞD9�h(jm8���{z��;[C�ȳB�18�DBx��]��[���������Oט\��:�������:�،5Z���|5����.h$ J��ڰ*򭹠t�>�n��ME���&걨ŭ�ؼ�6КO�QEM>Tȝ�wW�.�i�#3FӼ<Ѯ����b�B҇A�v	��!��|"��ٌ�ZcXڜ;���)1��}�5�-���HV]�����V3�ZW��"�A��g$���o1Y[7,�r��6+�z��􀞭�g*��[F%��M^��5��[����^
�F�h�8��h�e�y/j(Rc�suӵS���Tmc��Oz8;��8D�X"u�띯V6�{���B�61M��r��j����Z�gZ����Q@;���دª�N�E���ܺ�d�9q7W����R�5�ƣ�E���J����a2$h��*�*���ߘ��S��WV�"e3�J��,-q���NI�b��i��]��v��hU���8��X�ܝ��ޤ�]�P\�q
�澛ЄD0�E�.쑳���v�pjٶ�{��l�Qz��F:�+JU��=NaB8N\0%H��D呬Ȥ����W��x��;�����㏮Hm�v!t�/(�5f��A<��8��h�Nt8�V�e����|��8���FD�������%�wc������\�Lv���wJ�τ���Ki'��=]T�>2�:�Y�ڝ]R'T�hm�`�!��H���U���r7��-�w��P���e����
.aYY���k��j��;o�t�MF����]�~⵶����s���^h8�7ׄs�(�{ӫ2A�j9�Eox���1zr�S��� �&� C�rCQSM��C]�W{�'�tUҾ�ŝrN�w�o��2�:��a(t������͖���*��u���a���	��c&�0���o�{ci
˶Ŏ[X����Ar��]�L�Q���B��w��P���tק0������HaЬ���=Z�C���zp�X���d��H�o�ԫ׻��9�n÷�ͻ��մ��S�y���V64b�A�^���'���^텝���x~��VPo:��ԩA�W�侉�zcKo���1$�{&װ�l�h3%�Ă�����^��0��_�C��gaN��>�=G*��������]�R����Cf������M�hn�Ek���ی��	��[ފ�zث�Nջ�y����3<M�_T%�R��w���L�V��<�Avַ���.*�b�0�漵�za���˝�QI�һP���W�K��aOGES�)l�S1K'�@�bj��"��`���YOZ������х���#6E��z�2����������44vzp:�ol�V8ݶ������f�,�څ�kv��fU�ˊ�?*^�S�U�j8^���\_i�ś�˸�zس[������rM�dJQ��:i�B�_w�`ZG�u�罻�|�w7t��\L�|�X�OdRp+�P��g��N��l�3ܩ�s�'@��9��MT>��4�I���q�˔C�"�7�Ya�t�4�ј��Q��m���֕�Ю���1`9�7�����%���������7��}�V1=����=��nK7�	X>�h'�m�K�-�oR�U�6���(�R�̠�X?h��:n'6��*ٳ{F[HrUk�&�����OBx#+�Q���[n���
S^8Uc���M�n*�A�<3z{��V^�7�*��91�z'�W��4*��oz��lO��P�5}��}�P��s$���\"�C\f[�U�z�e�ur����F"���yl^��c���Vtgj�1����æ3)`�u뷎��\��'�}�qblCȶ������e�c���ef��}T�� r�Z�:S5�s-Q\��q²�Rw_��ܡx1�C/R�^�ޭ��}]~{�|�KU{p>�����^���򞔱3s�
c�$�����s���%Իޮ̮���H���Կ}Μ��m�X���+�-�S�;��w� �^���Ȣ������b9�m�Ҋ.)�دN�E�}t���w7%1�qx�b�3G�c�j��{N�[��S�ОT5���ᙃxmms�:�M0\1���C�g��8���\�d���@Du��B��;S��m�)�%E�2�6�����<�UOI��v��B�U;3��c��nI- �]�ܝ�6rnڥ0��e��2��KZ�'��uu�!p)�r���IS���wX�����4����1��l�P�q�!�d�B�ӷ�N�no9\zi�z���Y�n��Omc���d�V?=�w#D9��s��ݝ�/�e�:̑Q1���Y\̼���-=�qM�:�>��\�m�別���0�oh��O�"Dcd`�X���)ۋs8�Q�:�RĜ�;A�Z$�*aY5��:�<@��gD��}��s�Ǯ��w1�	�d��CQsMaq8W
��m� t������ڇ}�t��iE�ݨ���y4&�|2���|"���'w���8��/M��A���D��LM�R���(og��	��h�y����l؈�Yf�JGfM�9t�:\sc���]'���YA�帚��1��5q2,uf������w�E��M�wYT
|n��1�C/R���սC�uVd���v{q���,�<�2s,(�o[�Y�870�`�]Ҧ#���j:��l�&:.���I��˚�q��l�TO+����lWry�I�6x�S̊ˎ<���;�k5h�;9�5��Z�n��oA
�~~{��c�����{�̍Y�����U���8�#ρ�'j݊�D\� ZqδX�ט����N;��hL�a���	�������9�v�N�nv�A�[֭��Q�4.�.�*α�!��gZ�]��P�.ШvR|P�V�8��o/��h�e��Z\��\u��m[�����l'�4v�<�;����x���o0RG���}���硫>�!�e�.���$����G��瘶�6#}�0'8KP{Q����������U��21*ǗX�8���#�!���X�Ѫ���WV�fT���3]���P�������z0�� �P+͇^CmH��[Y�����t�]��q�{�PVl�َe뚰Z{ �5(j3Yj�3�]���1Y�U;��d�uG:�F��U�آ���2�dy��-F	��q@J��Z��򘫎���>~�¥��[{��� ��N���`M�m5x�U�G���rՆsA���j&�>�z��kY�N%��v�\� 8���f�g�����/-r��&[P�]F���s�C��.]�:�V45��v�;z�B��Uǃk�ʄ"���4Xi��d����9�|�c�,,g*�*q��z&�1g@!���7�GV�)�MShk���/(����+Zu9��3E���ƶo=�O7�l���``渹�rm ��۝	i����!t<ޥ����|�����{-CV_!^��|��b���ڤg��g���/hn��>s�1�*�_lo35�vu�A�C�IÆK���86��Wvr�ds����c�X�V��"�0j�b_ƷbZ�P�e,��x	�	2���`�aS��S8xu�-������[��z�+�'uj�*E�Mh��S��*�CZf�SM��T�Y�0ke��EЬ�A`�VԬ�ڐ�\t���8�t3(V��7�����\���Z;9pW��v�w׉mpʷ��z9C�c8Sݣ�_�'��Mhi,�`)\x�q}6
�7n����J0�)iSM�-[$�N�@m�}ˎ�xμ4���5Ɩ�!8^�>9^�`�pQ��
bâd�a���������
�p^�!.y��wذ:��Q�C�)� �v�T*��j¢N��Y[B�;�u��������%�I�/�e����Ȫ9�A�����f��R�ux�b��j�yYB���|O)��Fny|9�f�>�*�F�wp�݋�K0J���i�;3����gaR�+{Nщ��Ե�81�ӷ	��1wj���R�)��r��F�O�� ��Mb܉�ܮcKӠU��#Y��X�W߅6놪�����䦭�=G[���}AEżfu}Jz�=���u�����U�g	[�����œv��#�"���-���]vhsh+��� ��;�������6�;���V�p�L���#;��X)�
�@ҷV���rYڮ��7hAҟd���T��l����7�n�")k�o�:0gN�b�!���S��l�)�Xv�4��w���yU���;*���H.�͂u����f�N��{�7�iA�1�7����F�L�_Ír�&�W]Ko�)q+P4�r���$|�$6���3��+s���y��1��!��a�6����[���m�<���4�+u�V-��.�*+��9t��[/0��@*<V�e���ْ)�/>x��AE�[�A�텁�a@��ׁ�^*<(m�g�S�4�Z��ؖ�A�O]�k�k}��1�g�SH�hqM�!�x=3��[WM���c$����&f��Sz�����Y�yh���e�������g��ִl/�V���&ݨ������ޥ1����C��BQ����԰�"Жwݑ4N]�'�\{�o�t�*w���c��;���"��3 �����F#Q�(�YU������- �*�b�eQYAAE�T��H�*+lA",U�ŅJ�Q�b$
�������EER(���X,��kX/��1A,DH�X
"EU�i�X�`�cE��(��)���b)cb��P��k��cib"����d�b(�b��fe2Ҩ�-�(,�bX�(#�"$��rؖ��((� ���(��X�c+�b��)Z"���3,PPY(#(E�%@Rۻ(,�V"
�UH��F0PQ`(�*QX
E"��Pm1��QdSI���5\��Y*� ���k"���"����PU Y�a�d11ci]%AQE�X,*Da�d�UA�,D]y�xoݏ���~�1զ�[�b��q"����d�|s��@�u�!+��x����r�}Y��>�#׷]�U�N��9[b�\���M�V*z�R�C����rZ���B�X\�R���)s�C9�k�_��XmG)���Ok����V��eU��=28�����:���DK�f3)�{v��ݤ(�lX峰�kͤ�MmE��ۊ��1�Q���ڢ��y�����¬
ʢ��0�^�Ag��E�qs�~��R��6>���k��/6q�3BwK���:�6��`�k��o0��{�~�N����qm�u��k��Eb����;Vל;���v���I�����B�=h�e�!�b����}�.����#s9s':;�� �fHbq"���q�#=�������t^)p��`�;�$�k�ٱ��#G9�'��H��j�/�]
}�e��N.�kx���gD���]aOEb򠆎��<���Um���d����A����`=����Q�/@�v50� >�eޱ4�
�
��
��Nkv�V��j��β���{h��sMg�R<E^�4Qfz�!���n>��݆V��f�ە7!�Hܻ�M)Z�ɧ��Y0#��Z�ۅ�u��Ȱ��>ƮM�e8q����`��j�;WOJ��F+�z�	�J&h��`�=���rM�dJ(7�^CmחM�jlF�g��P�g!�|0g3��ߊ�	�N�y!�N!�2�zM\g��Bw�����lP�<�&|4m,�t��bZ��4�O��^��3�X�b�%����d�«5_]-�e*�eoE6�N���;+A��#t���֊c�d�
�҆�魷uyWjkŕG)���(�G+Dld>2��e�������A�d�/�O45Ƴ�����9�k���~�f�"9�$;w�--o�Y�gj�W��5��w��_�nN�����^�lꈓ���K�e��>>�Vn��\��w:P�6`�u>�B�S�erH��OՕ@��t�b@�Ԭ"���[ٮ���� ������]N��<�#h资t�`������&C
c��\9��}�{��J����;�S�ȯ) �T�M���d�2�5Y�<����2��Yw{#� �km�ݼ=v)������<'a�ۻ���^���LBw��ٱ5�d�rI��^B��99�[/O�Jfի��q���\ߵ�w�[!�vn����S9l�.i���rI�h�J�6�4N�nx���څ7AM��Ѻ�9qx�=��nu�]���E�qT8#��:�� ]&�c�urol�f�����^gw1H�����㏓V�C{N��-�Z$h���t'�0z9��5�oi{����j�Qc
n�+]��kg�ƮO�f]�K�~Y�4-�vS�Fa�Y����%i0�#
�gu�/�=���M�R5��,Ⱦ�*1���B��ײ��T�ӈ�z�l��W⹙y|�X�i8mP"�yo3}s��#�!�K`Wp�D��ht�����d�3ˈ�a����z���<�W*�;�a�?��㦉|�n��s@�D�]w�F`bioE��\�ؼ,{�UsA�}��2�t�g�kO����cx�]�\�
�����߯�V�Y�RP6 �у�M�{)�S$�e�z2�����uOlمv��#��!��W6(1g�z����ݫ9�y�n�����ji�Tzq%��5�[���c�'��u�O�X7sE���{��t�u��8~���Ļr4W_f�5�kec��� �4&��CQS^|"��wq���v��aHX	��#Z��a�U��{:��:{]��e��*�h��ҧ���=��+��:U�*ﰋ������A��O���^�/vN� ]�\a%OMo�ڿ}ʊ��^R�YTo�P��6+�/R�^��N���.�w��GcP����zx����yE���;V�VR7;E��b�Yh��ܦA�f�m�:��{��U�Q5�{�����9�v�F��:��l���9uަ�$�.��i�>:�e6�gZ�]��Q^v*��1..���c��5V-mo.��z�g��q�v!�RQѡ��]�ӑ�w���h�f��8h�=:�KtS_S��'�>J;��}<q��m�t���b���v��RW�Z^u�C�8JP{V�/Un��}��)Wպ�Ǯ�g.��v�L�����^:�#ל�^��ϬO,�����K��rs0��l�{��HT���&s��ݽ��d�}�&���O��r�jYm�w0ڮM0ޞ��~�rqGp)z�7֫+GD .R��"����w��]��i,��Gj_.2
N(c��/����^���g�lc���߸��N��|�.,J�V9$ZfD�*Gh8���ج�F�+����Ԣ��?^�v
�D�mĐ��	0���j<kk��na6��-}�2�/V�L�:)��t�v�F	�4P�5�0(��jfYK���lU��1�}��	C��a�3���������ݗ3I�j#�K���e��˷��ʣ�ϵaa(|���VOeM�;#+����y��l�{�O�¬U�k���HP˶��/�9D�n��xuf�t�i�U�W�G�\P}V��*f�$8֭�Gz��ý�WDH��eTNO
[����!��9��	����S�������f��cՔ�	�B���Z4Hz��~�����T���-�9ٸ����A�l��g�"�o�%��Q0�תpĭ��p'��IVt�p�]x���D��gR�ϯ����[7��'yLQ�N���{,c���+��|z�����^��'��d��\��"�d�W��>n���.E�ϡ���b΋o{���ݩ��O�|O)s�\���25�o}��Qr��g�,�������W��F.�����N�nz�Mm.�j��%`:X�mQ�Gc��k�[�ą*���9���ة�(��V���twB��&�L��+V�kb�0��'���z(b�4uN	Es|��)��G^Ljsr���`��a�Ds�DcW6�J�.1�����{>��p�^�r���n{}�rR�k;�_�֞��k9&�2%�6���W���X����=�+#��i���ߊ�e;����{ ��������M��E�Oc�,��2��>8�8����Ft2�4H��.v��^�&��Gw)+��%w!�hK�Dh��&������Dc(��ۉ4�GB�s1�f^�v40�ǳ�(ɠ�d���ۺ����������^�u�GQ�aXFQ6�>'��:�;Ӵ8��ˤR�^
}���P�ܹ�'d��}����T�p̓�U{:�r�֒��N|�g�Ź�-69A+��V���)�CY�:�x��.稵psYE�g��`�i:�n�bw��=L�|�`v��6x�ɜ\7b�xC�c�}�Z�4�ESCY������^]�@����OD]]������A�B�Z��Xoڢ��y����tק0���
���Ȟ+;�.NjS��&����ƌ�A�{���k��xa�s�u���ML��$��η��/��ʠZ�t�b�^�h�>oV�{]�v��:����q��5��[������w��D\���=h�e��#e��MI�ԕMZ6��u+z���Q�$\�D\��J�����ˣ^Th,�_u#\\Rz����}���Ex�\�pZ��)�uw2؞1�R�vu.`�z_k�����p�ӵ=c��:�8����]�6*N��Z�Uv�z���%�m$���\�f]�.+���/^-�uSɇ�*1F�~���/U�w[���{�]\�����O VG^�DT�bW��Q$p&Ne=�J�/[Lm�WpZ}�x㦣�}�ޫ�]���֋�K稷�:�㖔3B�(���MH;�N��$�Y� ��JT��dEA̼�8��c"�䮮.�	m�/H�	ߌik����:*�]p�۫q�)SR1ǳ�w�E<�3K&�a����m�WP�D��}���M��t��	������qa�%M���Ν����k�
�c��hq�V#82�9mT�z6"J���rz�.�5u�YLtՂz$�\ԡ�'
�Aρ�')n����O\O^�֢�ݼqZ�����=��4�d�CY��WW�%����l��*�ޜ��+��U&��E0}�:M	�7�$��T�6�9�u޽�t隡�yHJ�<LC���>T�qlo��A�v�l�����7o�"�˽*�,k��,&2jsN2]�o�2��4Mec�����@C�^S��&��(��C6���V���;ԗ�N�}�6*^��c�*��ُ	�ةV�>����������"v�������꼼�UZ��W�W|Őu�\z�-�μ��R�������"v�N��j������R/;\q��.�H��+7y�CQ�%����H�˟fcBV�)�O̐�r��2<�:��O"뻍�"�����iie���g���0��u�����ꖂ[�%�F��9��,[�	|��a�I5��ɍ����N ^�ݻ#�r]x���,��Dn<��l��S~M��;B�mG;���U�Mž�;uTZ��	W�lQ]^)5+w؁gغ94X{k{�:u:��bBz�����2��F����O*�?���JQ�C硫>���|�;�ԭ<&#��OW9��W=43��!�T�t%(��|,�U��/�:�����t�yKWfJ��$�k�ݹ>�̃��c�^¸Ut7W��+��8&;:���[���e.2�����i�RP)���m�C�*��0���Sˌ�vL�ݾj��|q3��ղ��j�i�Ю�Χ�5��:H��}�h32yV��&�.#F�Ήo�h�-@s�j0M{��=���,UOiu���MM�鳇��EoD��J'�}E��!���c9[i�12����8^
��.�eQ�l��䡹x��=ʔ'66/ �g��4�[�hA:"��o�D��d��([Ր����+��H��unB��WU����`l�6-줼�m[ri����ŃW���f�[;)�}�1m�Y��jDxw��;�<My�
��h����̞����0q�ZN�u;����-��]��O�vO��4���@NaV[�v��7�6����k랼+�!;xS�c6���=��,��;ڢ�}���f��V��޹�SVr0G47�G�/Pz�1�����^����w�G�6(6/H|��<!aU%D�m�Y�����;�C�;�U��s�q;��z(���)p���ʝ��=qg�pZ�o���݊�d\���3�[��d9�łmu
�+�.��ͮ�Z���J�u��=�P�S$F��=E&�i\}�F4��6�:f��j��kj溱�	�u����*i��+ťr�w��Y��cԷi������0�ilq���yN�����8JQG��ոhQ�1�˹�uvSmA�)�{z�H���ƌ�e[����p��1��ɦ�u���i�Q^�;�YZ�{�]\�dRQM�Ǽ��}B"�:_a���,@��΂�g�����D~�;�F䛹7)A�F���B|}�9tk��q�3��I�{^ �g�*.�Y�˷����#ux�鞸��a�ƾzS���]��8c鋱�	�� D۸DV3�y*����<݋V�<u�U�6��&g�¼�iqm�rІ�����
�PU�5���ڽ7Agr�&qa�q&�fl�S���.�M��_^2��5�^`'�G���Q25{0�{��-+�����6�)ݻ�&��,����mh��{F�؇�� �K�&)=��)V)�y������0H��hc��w��am&�R�ǧ*�ʳ���KZ����q����C��y��hS�_�h���.�v�n�p������#��[~�X��Xޙ�D��CƭEX�T�*N�Sgvv����7;"ihir�=�wS���h������Ы��I*n�RX��y�i +z_	���O�n:K�H]�j�Κ�f�Q��I���'*�;Wo[�����V��N�N
��Ҍ����Ԥu�#䯻 -��+Nv�L�5�N�іm�"ɷV�[u7i�)����]��(�p��5��J;�9��t5-����`���{.,O����,o�k���aɹ�J����xF ��"����G��1�i���x�PgR3_g��#����-���d�#J�\�~�Z���J� �tR�s�hRЎ��+qlkz�:q�*=�FT2YeÂuCM�|X�$�,�;��i��E�1j��4�� �����K��N����Z6�JWŌ�ܫ펃�BI�!K��9���ӂ]�QF]�ٛa�����Y���p��b4��M�
?n�:}u��U�3g�v�];Ɯ�l��K�_�N�oj{� ��#G�ȉ�T�k�X0�YP����ۺ=�<�=�a4��ۣ�N/7Iw�v�1J\���,Qɱ�N`n��(gL����`vjB�k�x.�+����;/O���Ղ�g����9D%uv H��d`���R�pOЇ�mΙR<���I�Y�Tw�^.�*̗n9Lg|�C��e��h�P�8G۸��Nzbe<Ī��*v�%r�O�Α
�B���%�,u4�.�,�J��%�����N�0���d��ǴvM�"N��C��U��dm�a��������e%�(�(��񾧳��-�l�y��Ue�I Q�T����ݨ��`�V�w���l�Nԥe��T����������8w�`��Wf9"�9W��F�M2%�y�����4F��.��؆Gi��{}{ڈ�PU|@t��X��/��٤4m���B��P��'2ke�8��Fլ�c< =�ٝ;���h+��M�ΰ=�G;T:;�.��[Ӧ9.p��s�ӻ��$�՞�{�����[h�"�b�H�(�T(
�"��i�2

"�,4ʌb"�b�,F����Q@PY>jdY1� �Q&Z$,��
�T�Y\j9eC)H吩U�����ؙj�B���26��:ʐ�J��CK��*,̡�����V\�2�U�",����(���*��2�IPF(����1!U
��Qj!TT�¤m�J�ɴ***�L�LT�R��m��X��AeIR(�ъ�.a� VA�h�)�2cHQZ�֥j,ib�%b�R-aXVV�Jљ���ְ�V��Z����m����@�(���(*�J��(�
mC.PZ��S0����a�2�%n�3Vh`:��1��Ę�h���H����Y��eE�b��0����"��̲��n��s(�DY�`��*�q�>@>���5{n�fj��k�䲑MJr����pQ�ܴ�Փ�9���i�;��=��;�L�c9��ݶ�&�k��n^���8:�=��Oi�0cdn�v
�D�}a3�����Dw7�Ak78��Ġ1(f�|}A��4q��igC��S�{���2TO�ۂ�Ĕ_��5-}\T��'
�C$�4X�n�S}�n���A
n6�ݜ�\�(��#���&�A��C|?Z�'�ʶ�:g�k��,ҍ�\�]~ǇG ���E�$����a����98bs�?R�{��ȱٽZ�m��m\�)��U��v���)��|&Wo��:�&ǝ�̲,GӇA�W����8С�h;�k+7=�������h�m-�YSO2��x1�Q~z��b��|e�Aײ�+E��[ʪ��YqO�E�T��.�/��W�������[��G�:[��֋���A���܎�Jz��y����^��k�X{�A�\U�'j�kZ.z�A�S�i��ˣ�-��u��V��M۬s����L�ǩc�6�6�{\)��0�f�H���sZL�U�-� Ys6V�.�6qA>��dNW�y�����/o���T���g%�fB�k�{EF�����f>�/x����7Ϫv��j)�M����ubgo�c6���bem�J(�\U���K�U��iFn��X�*r{y�*ǔ���q��t�N94_�;S�Alr24r�W��X��	Auby��+U����kg�5rCl˿C�դ�����:����N{t`Oӎ�%�Dv����;��}�=�`k9'u�Vi)���M%��.a���:���5]S��Q���n�T���w^�9Q���%؅^ձ�p[Y#@��Sc����u��'э�I�0�DwX���vf�A
�c[&y۷5`���>E�!�&���r�%@űe�n�ur�F���n(����PmC��Z���A�%fkmIyi���(���{������ފ@�A����Z��|"�O&:%q�ܾ�*�W5:�s��b�W�.�E�Hgƥ���6�٨��x.�L-�٬
���p��}�J�htP���f�F�%�\P��U�0�� ��]���Vw
��j��ר�`�l,fZq�f���B�CW���Z`|w�K����4�d �/���1k)�-��h�n��x�q�f����ɩz��$�'�u�	�wE�>���\��jJy�������@���2��4�_``!{�懪�3�t�1�{T�����S�h�@�Ǝ� ���6WQ�7]Nv�jz'��5�o��9��{����wY~���M[����	N���G�Y�Y�9'�����נml�\�f�k�X{�N���F�Q�&��1R-"�Mە�Ԕ���Bk��dk�ۋ�����mEat�D�'\1W�Kq�)��V(N!@�P&��Wj��G6�؇�I��e�GL:׹j����D�3�+��������zx����z~�6�r�A�p��o�Sۣ�/ܸ�X�hb�4*��(�{U���u��!A��ru�t��H���>� ZFA�n+�/m�*���}���:EDZ�2VQ��J&I,���f^__�96�H�� �t��4:/�o���޵y�U_٭'b��"1h����KK���.qg�F'u.�[Rn�9`�t�2oGV�ժǒ,��@{�Y;�:�D.=��p��gя�'�i�*���}�T�jL��%\^�S�`G�u�L����;G|̡pFޙ�6�4���D��0���Ǔ��5Y+sv
�e;v�����ؐB��Mm\ދ=}�_���g����{���x���<U^��.S��p��������"%��tw��= ��	�^��B1��d��Uq�D'>�v��yN��P��$�S����V�:-����9�L�w����Koī3�*��ȱ
�rj�YF��.T���miچ�^�s�!0�A���2R����T�>h�"�vn�s�*Y-��u0뱙[���3ܷ(�0D1n�F�H�P�Q��<"���C�S�|c�o1��;�4���&❳�3�܌-�G����.=��y��\ñ-�\�
5<��q�Q�J����g5�]VzS�^I��e �^��9�-�!�u�	���}�_�r+�2�(���g��'��C�HU�ߪEE��=D�h�)���|5ڌs��p#:�4|b�@�\���K�e��:O�)
P{%`� ԇ��A��N�V�+C��_z%\G4�/��RIkr�/L܈���5^� �S�#�Wx���j�Y!G�|߱f���6�N�xXc���S��\�,v��Pf!�ml��M+����[q�@����"�shhO�4.i�.H�{��4Z�V���	��F�}GBy�w�hԘ�}KMCC�^����u�1��g�}��Z�+��_������\�9A���O.��9�/%�w��xu�{�)���Uo\��8����A�:�9�l闂f:&�/��D�09�*&Ű�Ȕq(���Q{��-&C�E��'%<�vs�'���;F������8w�@q�h����J3"�=�Tl
�8��yɎ�1JF9i�@V����bf�*�G;0���{^Z�N�qb�۰ܥ4k�·��]��գg��CZIߺ�#*N��v��oR6�r�%P��2�[OE:�E����<N�bV�\ùx..�4СU7����X���@ވ�Md w��S~(S�4����b�"ʪ~���Y�|N����P��˂��ֆ��;�b��(C���5�hS����q~x�sg3>�/����]M���V�|b���)�k�Y/V��1Pp����9�0+υL�6\h���aU���.���9�f�uiaG�r�Y�nXJ�(�U���Yo>�J���)v�A=��k��=������j��_i�;gi�\t����YBom��9�ж*�`�8�oU��nX�����8�zTL|���0zI�)`�A]j�s��Z�7����	\��-�=�4�	$�/��CfMt����"N�@l���=�0e�=�$��5�����̺W��+�3F��@��m8���A�L���ݹ�e�b9,zv��N�{������v�*�?"}�łr_?y�[]C&.��q�]�(���/�[!㾘t��{=��f	��s3G^����6���1�c�Y_?P�k��d!7�[�՛GR�-����*-���đ�+�b��Lt��� ��*�zm�0*DE��b$���;�s��i�^�E�	�p�������I�QqC��@����}4�����)ڌ��ԉ&,9q��l���M�W��1[�m�no���/�E-3Ң�nF��=״�*���Dk���8�ʋT�+��:�!�~���ƈ����ӗѴ8�ھ������"a��z��b���A���2C�W����G_�����b��#��_kw/Z̢6�?s��"��2}���1ӐjEt��Eߡ�P}�r��Xh�:<������n�Vp�<�/!s��Gd����D��ت��s`�7���ne�v�9�v�qW;x�i�f"^AN�1;{����l�����&�}->�`���G�%�i�K��ۜٚ�"����bubzK��a�%�0�7ăF��Y훐ѓʅ�XPL���gc]�qT���]m�n���]i�v$�z��`�����' ���D�w.,:'[L���0�W����Rv�u�<}}�
H߮�haܽי\�P���MǏ�*Ω2��`������Q�B�\]H�p�iX��]����O��{��㢵���ס}n�����r"����Q�P��>��n_N�D��-t!9Q2)�p66/�슻G#���BO�VC�X	T�{<r/�p��ZaU�[ө��t�/��d��=T��$T���C��G�2��MBۘP��V�TP�\�;x�:���ܚ�G6LH��has��L�\�k�8=B�ZX���kB�E�c'`>��ذ��њ�m���]���r�b��ԤlWA��Y�哣s;a��1�G��0���|]��}/:��j� �������v!��֩k�%5��^�&��R<< ��T���R���iۏ9ӊsҫ�W_�v�`����{���V�NsB$b�T+�{�j��r��Ny�S��Q\��Aa�yUUK�V�[{cwwS#�&܏o�Mq)Y�Ā܄�q���5�C�E�=i���!w� �Ğݜ��f��l��V�# ��'%�K"y�}*�>�9gB�}Y����9�B�)jJ�c��[}�?����  ��s0�Q�u�@� �.���CyFWZ��q��#�ځPjE��d��.$G�3��]A_;Q`}t:���'�Etu���e���9H�O˷�NDŰ��UXJ�����X�A+D)��s��������W_])o��%��P��15�;J>���̫�sPE�n��.'�ׂSd��G���"��e������;x�O�R����zWI��K�U�;����d�HNj(iED�1�m�̻W��^Q�M�.x��>�V$��J��`d����7�O-�:'[t6$*ɧ�^�����w�y���^�ԃ
 L.*/8��x��j���Ӡ�-�:pFň��j�5�Ǔ��""}�K�2�i�]��x���|\�^���T�/��v�*Va�6��q��7�8��s\�b�t$"�!��S%Y�6͊Rs�>�;({��8�ҫ��j��w�u�!{K#T":���/��'+�G�D�u�G0�Q���V�ZϷu�@E�=��z�e��B�#�aCYF/QMW��{V�o��=�d�VI��<��PxR���ֹ�+"Pi�\J�wz"f�4S�7��Ѷ\}��I��;����6(�`{mtxz��|�X�X՚�13�r�4�?"7oR�T��S����fv;hT�y�"��s����LQUfMTo�Y@i��z!�����va��U�2�lc,A��Q���y:F�׃�K~����Y�&���̬����X�[���S�S5�]��:�@a�Aʽ��jpAn�u�{99'E��!�Ğ��5��(���CBNN�T��vOA�y5�m
p�my25ڌr˧n2���-D�.��sJ��Qَ��0mi.�ƸV�a���.�F�<���RC��tl�ў�%�mb��w�u�z��[j2V�ȑє��WD�����{�5�V6o]�>u�׳e��G�;Ӂ�3},lې_Etv�s#��]�=-�2�	��^��ʢ ��w����P�N<ڛZԪ��-��2��d䷍�Q�veE���X��~r\L8�
�����/s�ൡ~���W�xOC��(ݶyɎ�1���Ӭ��]�T�&n(bێ�=t��W;�ɵ��a�����ܥ`�@�r� �Tn	�.�WG[�#��gݕCX�3���y��c�u�E�;eP�S�dԴU�,Δ�8)�77���,�0̹��.����Ĝ�	��G��}�mh%��X4��m|q��Pز)^&M��ዻ*�飽��K��9U��9\�OiRxu����lJ�Vm���}�(����=t����i]�ǹE�y�����ShKсmf��q���J7P�\uq�Ӻ���K;(`����_ރN�|.��2�xlTDYO�t��S��u���kX�7�bQSqw,C�Q��w1A�uBFP����{��H���O&K��y�*�/->��{r8�fz]���u��i�aH�h���ګ��
�Ll��*+��U�Kㅮ�{�d�M�c1�ؿag�r�C:��=�U��WF�{C�W���0�aS,�5��w7x!W�1[RjFA��3���b����f�s��*/��ޞ5t}��mx�F<�����G�T���?P��;����fvv
�}Q@�z2�Ѵ�8!g+y�n��M�;.���B��5�}G3�J�����TW��B��2\��0��5���x�y�������s�`�'j�j�0�.,:��;��+�O�ʪ:}��,A��V���E��-̛��T|l��]����]y���[���	�(�=�t2+o���-�P��P�!g�S[��`�A�л�yL�4�������YЀ�]�H�|��f�����B�� IO��IO�$ I,	!I���$����$�xB���$ I?�H@��	!I��$�	'��$ I9H@�XB����$��$�	'��$ I?�	!I��IO�H@��B��$�	'��PVI��Fv��7��@���y�d������`�p��L�t vuB�p�ED��  ɠ    ��!JT� 	�0  `20110�L�L���I�@Ѡ 44 Q!53H=ҙ3H=C�Ѡѡ�I&A	�A4ɂe���&�2� !Dg|�*�;�*���P+D����w1�|h���~�6	�\T%?U�,�$� e1��c��^�d���x�z|�U ӡs,��[�i�G�	���Mg���v��Pӄ(	���^�w��ieh1SS/����UE	��p XmCɼ�n�c�$b�~'v#d*4�ˬe�.&*�v
6:٪�1$��.F�l�lOy6���WJ�՛N�`�7qVfa؜ʘH�ܘ6��"�S�e�|��^z�#�HV�ugM�$�ꁱ����i0Ω7㛉Σ�y�Q���[Ot�l�
�uU�M�S���%�E�ݙ�£sUVf+���xv����mws�[��� <�{����s�����-��L��q鬕��3�����Y��z��b��w@����]^��V]��4�Q�3��8�c������c�.�� [rC��A�l�=Hk��%G�L�:O:�æUJ*���`��'6���p�8� <d���!"&�4 �
#�� J�j[B!>9�4&D4��̨m���2�F����Q�T$O��d���]�T4BR�U����gTcx�y��2> FRHBHD�O��z"7�/���F=�<:�Xmy4�M ���1��ǋ6�:�`
��쪶`�K�.�F�(�W��ݜК���0�@2L��8e���T�V��[4*����C!�d6�ΠlVm�\�U:[�R-%hA��f�4�A��%G
i�0ع D��_1;��N��8�=ލ̗�w�w�������ug�6�����J~�Sֺz��Vjj^T�y�t� ��Q"�k<�jډ5ʔ���,a��4�>R�I^Z�"�Y
�]���p�:le�"@�(���2�;�<��X�'k����9���U8��i>�ׅF東����Q�P
t�\��y�An�H��#=��&&v$h�"��%C���"��g�[+#"��\��-s���#t�鱗M^�)�ТG)��^$@CZL��&ڱX�}u,��2̌�b���g2v�sg'5��
�:t�MX��>Ƴ�g�'gةb潙�<�{�cA4㙭�!�Xظ��] ���{j��57htR���pu0�v ������\`�.f��d�HM
�Vj
':�:�v���LL�&�`�T��	0�NAvI�N�7Ir��w��-��~,r/mA�7�xp�:����aZ��h���)��*&0����x���m|v�ldj�G�����1�%~�T78�@~����L	��i�ڍ�w(��ff�����D�8L�n99�D�ts��ښ��F�°nb��GU�F(mIᷴuG<�ߏ@�&:��^[l�>&��;�
�璉���LtҌ��vNRE��M��5�Z��c�M^$�s7Z1Ww5�2�0��u�7��5*�n�3��ݧls��Yy�d�OU�R�H��lPܼ�nn.��Zȥ}B&�G8![K��(���(j,
	Fe��HJiޞ�����&���nfiJ��-/&l��U���ҺP��$u��L1�~y������y�F�
��U<K� V1��1��m���V�23�gN�L����Kt*�`�I)��k͒�\[����1�\2�24��Mg{�!e����s�k޿I�Fy���&�P�K�N�/z7���q^H�K(��Q'sws!�x˄.�\�]�ݍ�=6�VS�h�������6������L�U�J�֡�ֈ�"�K�ɷIe���娓J��? n�L�;�ы}�$����F�W{��{�7���{!��Ȯ�T����:�8(�����k=�O/-��b��]�������'`!3b��8O��dfV�vT�D�Dy�=���R*�;J��clW���**���QF��׎`jsq�&ø�F�jeTU��W�71כ}7؛�D|'wq�W�Oq�p�	�-���r;�<{I!ʊ�$�I�%*�ZQ��U ��B�UP�T�V$#��(�,�k�l�y��LW�s��e��k
�?��ek�[;��b0�IL���fpJ�Bhz�i��,58P���K[�?Zq���$8g@�9��Ѯ9��>Hn��f�_�D!lˇ,�y	dS����c�,�qcF�:\��,�K�w��3�AچM��Jq^����q+x"�@�@��!%hiN�U�KI ����T7VI�m�(g�������uP觭},􇸉A�u,�ĂYD��؂a��F?)�6P�T>��I�UPL�)b�ןA� �So>y,`����A��)T�)ى}mV/OL�Br �2��2E՗�Dp4ؠ�o(�-X,�>�,'9u�3#q�U �lR����A``�^�AU��9��J�#>]��`� t<���d���F�Ԭ�;9i���9-�a�
�V� �:T�,/C�%�!��B �l�ˤ��T���I:��,����V�-jv:\�����q��3���w
�sY3N^}C?�z�7t����u��.
���z��h���%϶)�(���,9jz����ن�N��
�`0B��f��B���L�)"ܡ��D�9㗶���`b�* �	���+�4�!�*�����ѳ&v�\V��r=灲'B��@"���H>,"�gy3��n:����qh�����r0�ҩ�8����Ŕ4�0��N�s&u*��jc
��� �5�W��.U"9Й%Wm�cH�
�J�,��6��7.�7����^̉��8�xx���l���ȰB����8o�����`3;�؏���ɿ��Y3M���ׅ�@1��'!0�{�>\�X8WfFB��^�l=18��Q�^+�B�d��.�۸8� "����Ά��=�c��I���y��09��u���ن�ш_;|,�}�spI@���R'v���8����)����0