BZh91AY&SY�Ql~_�py����߰����  aT]��%  �@�RG�TPk@
��D 
  �   {�                     m� 
)@ꀠm��HZ�2��!�Ȩ*�� �    =��
	�-n@��n�$�B��0z�����,�m��֌HH`�����)W1_]HJ����{iS�Rp�Ԇ��R�M:�\���yH
����Ӑk��֘J�
�� %�|�� {.��rr	gs�9P�A1�w@�{2@���d�4�P�P�A����@u�<�GCfP� �4�'0
�A��r�(x ����xv-� d4>�:�<C�����^����Ijy��Q'����� p�ܡE7ñ � i�N �8�v�*� $t�I�   ;p � �rC#��:h�qp�Mk��á�vf9؀�Q]��� 3���.c#�3�v]S��i�l�{���s0u��LC�����% � @@w;��Gfd���ɻv�GFƣ�v�!�g�s��W �Q�PSrE��N�e��.���R�YY�;�� � w1�p                             *�7��UTɆ�P24�M4�2djx"$�R4�dbh�` �01��R��J�h2h��� �� !���� ��@� @��H�I�M&���'�G�Ɠ1�b�����*�` 	�  ��O������h��p�q�QUt�I[TH���g������}�>絗������l�yn�<�=�?�����xla���a�Y���G�6��ls�^��������o��Ժ?����>VJ��ٛ�ݣ���<s���\��ݛl͇u��ѷ��6�UUU�p�Ն��~o����~_���?
��~;<:�������w�{����.��{$�i�Iy%�p����^DF=Q�DG�Qu��"7�v#M��UDDG�LWԈ��DDm>��5Q�DeW�\�^I�$���$�����߸ĳ{'��I-w���xK�'xI$�jܗ�8I,Βܰ��":�&�L�"J�R"'k��4�U�Dec�"j�$��.�{����xY��F�Q�Q*�""+�DL�F�5^aD�F���y�Ds莢#�j��F���e>�#�y�8�}�aHTDqR#_qG�j
Dm��#���m��?DGy�0�#XDDu��2�Ȉ�Dy�f#H�"4�}��N)�":�DF�FT�")N�e��:�݄yYy�8ޕ��ڑ�"2Ñ��6��Sq�m��eO�4��ǘ�)�i����G�"#,�s�h�:�㌶x�DFQ��:�#�#�H�#1F���5H�?DDF�O��X�^�a%�׸I%�1%���KKrZI/d��Q�O�Ȏ5���#l}ʈ�:��DDF=QO2�#ݨ�̣i�DDy�Te�F��""%���$�X�K�,fI%�P�*�8������(�#1H�"=+�0�"3ʈ�#��QE#�y�Q�����FQ���#1FN���aYu�#(��Du�"5�u��"a��$���I%���w�]���Z�}$��8I{仞�V$���DD�5y���#�D%�a$��ė�^�jIF�k�DDFݎ#(�1��w���I%�֤��Mc�F��DDz<�#Dw��FQ�q��"6�"�Q�Dm�ܗ�$��cWrK�KX��Y��I}�^K�jZK�r����Ϊ#��1��e��xFwQG���#q�B6�=��0�Gv�z��v��k���������DZy�S��EI/<=j:��z��FR�"#�F��Iy1��K�1ܳ$��j�K�-w�$�:�X��$�[�:Ԓ��M�w%�S�$��0���#q�F�F]�DDG�\y7��$��^c�I�Iki��VQq��Q��<�"n����}�"z��4���<�i%y�Gq*�6��K�$�	}{J{��%���e�j�"#���0������"&kH�M5ꝯ��M1���U&���r��v�8Ī{�Q�DvV�2�}��)��Q�G\��Y�N�4�*0�8�V�e�U�OV�vs���$|<>����sOc�򲎹U�D�DD�GYL�D{�����g	#��$�OTq0������cU����8�aL=J:��0�#�i����*#����F#�2��фa�a%q��l&덣L�IUG1Q�y�mG;ZF��VֱQ9\a\8�f�8�V�u>�DDgզ�O��&j"'k���+H�)9Q�\0�MTDOW���}�NTDjV�DLTG�z��/f�6���"5�8�L�Dq;Q�1�&��1��=�K]��V��[�δ��S��}�Ta�UTm��=�I,jKrK��/$������"2�r��c�L�DF��":�j�H����DDr"2��TDDF�Q��j#$�X��K�טI$��I$�a�E"#]�O-�Z��V��jU6�m�����#i+�%�3�$�X��IJo��La$��I$�	$��$����y,��I�%�8H���}D{���q3[DG�����'�I$�>�I�$��I$c�Op�N�ZcI>��䓼$�m$���8DDDvTaDMVXDDG��G�DOVQDLW�G�yכ�yL�;�G�GQU�""3��"#ި�h�Tm�JDDgU��DE#=���;�����v�D{u0��\a�G�^a�מw��G�R��f�'*!>�e��#qS�U�������2���h�}��m5Q�i;Q�y=T�#�qk���j����R0�2�QG5b���TDa%S���a��N�i��u�Xu��uH�'��TDi�Ds��}�oU�j�xI%�����u�$�Yc��ʈ�'\aڭ9��G�\�9���u�r=��0����qYyۨ��ң:EF��#�|�=�����jg차Fc,��m�m�#.�g�m�|��2�q�D�����O�#I����!�DD�R#�I���4�Q�j�٭��m;_OW���]q���ӕ�2����{�ym�8�H�ѕ'�S�
���"8���:�f��kΩG%i�Uʦ��>��7ʅ#	+m2��H�����k�T����M&�"2���i���i�MVQ=Q�]���WXDgF=]F]f�<�Q�i�DӬ}�y5]eǕڌ��7��"'�h�ʾ��5ZE"&k��L���ʍ�7*���*)=Q�D�DcH�\��ȧ%u�Qڨ���ݨ�e�̪Dc(��m�u�Vj""#���$��K�s�.�}�Im�j2���0�4�F5Q�"<�"1ꍲ�0�����"N���K6T���K�$�iL)���#2���"#q�S�O�������8�Q犈��#DDDmQ�F�F����F�z)�Ta�!:�Dy�D�2���㈈�mFQ�)s�DFZLTDGF5XDDo�%e�Qi��F�9�c��NW�%��K�$��$�_X�
^K�%�Z�Z��$�u�w�ĒI|����%���Y�,"2���"8�E:��4�y�GLq�G;T�Dq�8�"0���ۨm��,�F�n"";G�g��yDR5��&��VY�:��$DH���NE7)��De]m������uF��(ʑ�q��ѕ2�������w��e��E}�4�m9��V�m��#}D����c,"��(�[�S��9��Q�����?0¾�F��,��c{n)�ն�b#mF�j8�GZ�;�G^�6�^�GQ��Zx�q�J���z�a>�""f�yDz)�j�D�Dm���4�1wu�G��<��vTaǼ㭺Λ#-�"#�G�H���l��Gv��>y^a¢4���Q�e%Sh�b�ͷD7+N2�b��Ʉ�}��4��J�u�O���z�<�ҩ�#9�e��DiI\q�]��YDohD�GO�1�N�Q�VXuDG��F�Xe7Q�G�D{U�[D�FQ��Dg�z�4�ң��:�""j��<�_G��9Q�J�D�Dc�DLW��5���DerV�Gj�4�I�j#.3UUDDD󎲈�9�����쯩F�"5��ǻ�X�9�}������\����/��9e����[����Lm��J�!�ɕXA\����s����i���˛BH��ȇ�xI�I0��Vy�e*�����'���vqK�������]��Ab5�/��'��)�j���ru��}u�y��^�e�b֩�K��Z����͞q����μx���׮���~!��O��s�r l���	
�F�^��o]�3�s@<�t�U��*�n���B[s`���aV�2>���싰!`�Wl>Őb�,��sssM�D`�I��!��}����v3����=ߝ}��5��)脦ig��{���`�)�gm�uFr������u>q��`�t���K{�̇��N,�ug!�K8��$���> x������vӕv�UyK���DX>�}
&��l�����l̝���^8wݯ=�FxNFݥ�m��1u\��*P��2}�4�w[̾ېj�m�q�a����:���k~��?ϛ�J?D�?��4t����Ӻ��8��a�I!�7~h`���Х�q��1V:D�o�t�C|N{X�b�e�7L��,���n��AV{������Ȁ���^�?,�D���>���c*G�,�I�����^�g�A|E?'���->BҏU��Y�"A�������?���`? �s�ߏ|*r����j�1p����>ZSoǹ�M���n�Y܏�jT�	#�>��ss�x���V�T�{�I��W&5���Y�����fQ�w��@gO��=��Ě�L5�ދ����daw��n���/��t*��i�t���2�����^��pw:�zU��b�]={LVЎ�ߞ�]yk���sN�sc]+_�P�B.����|ք���0I3��>�ex�>���)=r�����ϝ���,m8ɖ=]`S�NfnNBAh�W��]i�^��hέ�iy�=��$ySu����k+�R�+$)^y�H}y.�|�ӕef<�0&o�;�ۢRv6$*,T��#�zW�}k����ۢ��n����&]�5j�|��#�ba�^���z���5�Ӳ?1��zϬ��]������2)�Ǜ�f]�4��ui�i�:�S�?�5�~q�Vd��φU�g�g\�`-�ެ����4m��0	�޽��]zw*l��ӹ9�&Y�GW�	���4,]�u�)�9��$�Y���6�IE�[$�y����M=/aE���3���I<]D�<�2�m��0
^��fm�q'�w�F�,�Q:x��]>�*Eg�d�:ô�͸��8������O���R���aN�I����*w�M3޶�0�3)�-�%�����9�r�4��j�cz��ׯ�Ȯ�s	��Q/��f��;�m����/e�=<����Ř.*W��~|�YXI6�t��K��s"������W/x�'[��}���r��Zd�5ܤ�e;J��':FU�nzK�3\|-��ۧ	6Ý�9���w�͹����nj�|��'J5��u�{�9��M�NҰ��������rRZ�+��xԖ�Y^��g�^ΰ*���9�2n���)�k'�#MY�(!�WPw��'nvw&b٘�e���0���˳.<`���__[�>��X�����
:z�2�W3�g�,Ӆ�p����]�=��(���Q�d����sc�T��ynt�� B�Ҁ���<u�I'����}޲@R�����N1��"�
_�[���1^763���4� {b��C#L����|�Cb!�:VF<I��^����W�]f7/2�]w+��2�ӽ�"&np��ε�擻L~J�=�#I#�s��Nlo=����]�c�A�O�:x��6e3��p���$N�t2�5��ט������\��/�_����G��@!�v�Hiw��f�k}z�d��t���,�z�}U�)�Ϯ�f������>����;���v���D\���w_:�ݽ�r����,��pb�ޣ�੟7��W��_�s�
��iO��Ϩ�Fw"�Gu����u�^\4�S����n@|��3Ŗ;ti�)=��	]����c����QON%���������/5'�&NZ}z��ҳM��Y7���n�͸�9�nvu��=ߡ��iߴ_w��7������y�:p���ϊ�rf�V�.�s�a"w;�ɷ0|yӄ��z|W���+>33�Z��Q�Hz*���FI�[��=��[}����TcӒ��3��Ї�<iO�x�A����oO�0̈́�����Z~�1>7�~M�bbn�[8����5���r��t���Ouo�L&V�R�x�S�d�+��OHp�K�]/p��^p<,_f�3Oڳ-����������.���t�3���k�렍�Cβ_��o��'�"�������-:���9\�̀�û�6�{����}{��/o�;��؃���t��;��//����]�l����w�I�J�w�����)�&��o�����@��HA'r���Ѻ"e��w')N()���g{Ԟ�1�'v�=#�.�aj�y�{�ODGL��(�ɚ����@������AwJ�KјPb�0:VE��.CB�Je־���}�7	���{�v��!��q_9.���ޛb�aX�m��a�Ow_{��HD�l�7�V�^�)�{��I�ޗ�Q�4��>�m{x+X���F�����>��eo���z_f��\��D1�ڏM,�������|~���W���p.��H�6��K>�h��uM=݅����|ߏr$����W��
Xd�g�m�������K�i�	�ޓ��׃F��?w�㭢�d�s!��{�<1F�Ϗ��Qʞ��ϻ��fF7�G`ԎZz^��������}��'�M$��0ǃatx�Q���r����v�;Q���x|V69�N[����Ϥ^]��Tm�4�џjOݳ�a>�����
?`�o��xq�%������Ӌ�w����y�>�C��z�}9�i���0P��5G�1�s(����Ov^�b��}�}x��Ϻ�7��aD��8|rMPp�Nc�z��Y8QǏ�}���vc����9«fp�V���ԍ1��>�w�+��������	w^3A��*�D�F���R�&���}���r�&��!��J,�I��8��n��>�#+�J����r�Y�6cˌ���>�\�3U}<����{D.d�s3�w5k��[z@ڡ�gD��`�� Ax���Ǜv�⪪=�.t�Aol2�İ���ɱ��zn�����݆
��b��uu���c�Ҥ�:C�y������i�S���Z{���ʸJ��p���^c����U�K-:azt<�����Wߞ�_�Ýs�Ցw��~=h����g������U�U�i	;�����3���6�K>��&����v|�������<�ss�l�z�μ�e9cå�<�WW��^^6C���6a����Or�s5����fk��ۍ��g���e#�Z"����-c�a����E�����~>X��Ү����Y�qJ��y:��v'���n�-�gS	ݾ���3����u횱��3	�%BI�t�Lqj[�1�/��Ù;�1�-��s����g�j��8	ʉ~ע�kvv݃'2��]ѩ�c�<k�ᝏ�?�|&NwaZ]��i0���9�LG&�{�Jq���s>���S���w��N^�	�a�j/���?H�ju�Oe�z�Q����a;�籼��H@L��ϿgN��=����=_�h���?gٯ�n|Wk$���k�%��C�3�N��?��g�����z5�뷜��Ɨ�sݻzf��ҫW�#0]�{.R[|�h�b���­����u��i�֏�c������'Y*͚��l������;���ݿh�]����Jgu������n���{�w>��嫩8��*W���ŏ�2�x�u�h/����+K������=�հzt��L|ތ[c�e^ӻ�Q�Z�i�ξ���}�P�������,]�o��w^��=Q�7شڼ���~g׻�����\��#����x�����|^��,�c�x�n������3����L�f�?g�&
��_����n�j��U��lϮNۻO]y]i�������ܢ��c�B����fǷ�o�|�7��#�nBaS�5�q[R�����ƧanJ���7��� � �=���s���I7�w9�Yۅ�5�O�.Tc�"n;%�����̺�껶�gp�^��=m����y������ۻ|z�����D�p��m7x���n������m�����out�u���:�cs�o?ݓ�������S�v l��2sn^C+�ވ�v���q�q�c�X�ְb�]�4u�ߥ��F$��"2F���rB��ꐮ�<��cee���,�vS�����g���������b�����99*� �^[Ŷ�h��ktr���n���K46��y��¬m�t˲������h��iޖp��#�5�*�:�b���̓��腵T:��t��1�.0�Q8����x�c}��g9�m�5�M�#+�R�!�][�1>����]�����Onj�6��;qMwY94Yk�����ǹ�~'�NB#G"�q�vqvq�uk���n=��e\$b��hBC��(��Q$em���X.][�3ݎ�;v#-8�."<@̸V#S<J[I8�v,�gj�����j#�i':{X�=���t�{{�Gm�Ҟ���n͵���u��sy�3��d;j���n7y��]����v�w�i��^�+�nxh��M�i.6�ɱ�<;<�cs���F;sl�Y綽���]���@À����d9$d�A8��Y�N�v��I�wǞ���ڷڬs@uڏl�m滶;A%����� �0�<���`�kՎ9��o�>1����[��k�ւ3d�\�g��v��%���>��2�[aܶ�}����P�EqI��j�V ��V0�I!M�.S���}����A�<o��9ӭ�mԊQEJaiݦA��Qe����F۞>�c=�h٬�b-���w>|�����j�eN��g*6�)(y`qsqLH��L&e(�D(�l�!��
f	^n�cؚ4Y$�H�A��%k�p��`5��w�����7�E6���"|�.�!k��q�⌽�a}��w�������9�Ols�3=-<T![@�$hSI��f�b�0R�B�� ��
�Z�$)A`��!���A���6p�I	�W4㵤I-��`��� �Αp�6{|��V9��쵸շb��V:�����"v��)�C����wn�^w\t�=���Ii,��ʲ
��Rɍ��������6�\!�"�R��dp��C���+(&�.��KlF�\ȸ-F�l��9��#mO�n;>�;|ʿ��w9<�]��L�.�)N��.[ܷw�l��t�Q��Ucj5MS(m��/(��dv�:�ϐ�?���7�������R��\�]w����c�����S��ߛ�3l�>��yu�>]�f���>�s�m�����������K���ۜ��M[�p��Y������f��-�5WV1�u^y�X�?ߋ�ٴ�٣ס�� ��hxC� ���C� 6�=G}� � ���9Ͼ� 6��`� ��������מfSɳz[:�um�[(�@Vb�ef�1� ���&̦��1�e6����M�fH\����װ4; � >;!�x>O@l  @ ���@M}��|`f 6�s��v� @�NI3$�nI�ٯ���1C諭��S�ɴ�v�Φ�ۓ+7Q��]]cw�<d��d��l��v��������2C���`��������Ͼ��{!�G`>@ ]u[�]1�x��V�(^�6V�51[j�6u3�-ūy�5Sv�l�7%mJ�RG=p�C��-[�9�mɳ���V����M�56�����LQ����E���ij�_9�|�w��`ٛ����������?�37���ȿ�w�]ߊ�/ͱ~$��I%�(eDya"#,�":��(�Diu�\q�#�.�[�$��I/e�fKRY�$��JKR[�$��nԖ$�I$�$����#��<�8�#!!Ē_K�%�IfI/b"2�,�:��6���""4�H�l"#0�R��l��Dq�a��F��")�qM""#H���)ꑴDDya�y�q�"0I/$��K�,K^�j\mmN#�8�L�BFX��K�$�$����%$�A|�f�� ����m����=�w9w�/�{=�}<r$��
��\U�s4��V@����㋲wN_gu��cSq��i����ӻ7S��sS�����d��{' �p痆Wu�qq#��3�N���4=�Y�v��/��n;?]����6����"RO�vǤ�G��;�羸�,�vy�����T!G%��:0��6�wC�WP�����}���5t�`��۶N�x����hF��Èїp����N;ROm��ΰv�Wa��nݶ��N��ll�"na��x���7;}�~Ll�;��?�V���n�;ki�9�:��ɶ7�9������W4�U7�y�rR��vv �չ6=pݵ$vc���y�t�ȯ�m�Z��e!%v����Q��Ä��$G]�0��C��4`��o.��q�YR��s����[�N���L��9#��M�A���zDE���Ux��힖�5��;�a:�m�g��K�C��vnzK��T�:�b'�\�9����\�.�����]��F���2N�a�G7n��s�<#pUc�3�n�t��O��V��Tr�n�\ObG\�l7��G0Z�*s��s��n������r\B���5$�V��n0)����{���v;;�N�>���8l#���Kgs�ϓ��m�c���q���	#,6�M��l1�5ۊ�q�=�<�^�n��t����b"�L�2��q]�]j���{j6N����#nj�[�q3Ɏn��
�i�����¥�ۯF��J�粽rwOn��M^n;zr/
�馪r
�]�ݳ��g,u��|۸ ���p�,z<�k��R�u�����?Z��m�|Fuk,�����֞s��Y90𝶢���ˑ#�n��x�AE�%�:��<u���w0�s�>�]׵s��;�"O(u�6fdڶ9�n���>�C��s��đP�F���n�de��N`�C=���.������yluW+�ٝ��۴�`������z��v&@7`�J�1�y;&�mT
`���홠�=�@ηe7:W;N��D����;�q<O%�s�um���K���X+��z���um��|���Z�����r��<mv��YC���`�^����u<��$�����o{�������c����g��<뮺��s��9�s�o����������[�[h󮸏-H���#Ȉ����L�҇�=��H#�DPB2$�Q��A(�0&<�Ib�,<�p��"�(��n{dr��	����9f��!s�u]s��Ən�vzn�>����V��n6�=ڳ���㹦i{l�S֔��91�GaK��=H%��a��H홌7��@�fn-���uA���4n��>H�=c��g�����tG���f����Ϯ����D{5�'�sn�|T[���\,)��wg��y�϶��w���7y> �;!	OY�!KQ-1�t�rR,oT�(��ܻ5�1�r6I�u^�Ta�ʊ_��!�p,cI�t{r|j���R��?���l��d4��ios��il]<�{��ĶC�a�8JUu&aA�]VC�\�s��ŉm��G�����O��ե<?��T���B2�Lc"cN�+4ãcxCKL ��8�	�Y6��M�Iu�Gj�^�-hB��먮Be�����!A0Q�Q��E�L)���s�U7#���M�12����:��u��)yDy�q��i�Zg�b�P����SlL�C�*1�i4�>rܪv�ٟQE.,:����F�x�FS�r�\��3�F��(p�3qF�M���� c׊4�f����7׎�mʫ^�֍" �B!f�0����Afr�s��U:p"�ճ������-���n��(˦4Λ0)@��l86A��s\�t�Bʫ�Zz!фC9�h�Ts�^Lꩃ��xZ�ӄ0��S�6�"#���"���G�G)��e�>�_}��yҫ4Í1��%6�8s��a�!G���FBx���4R�c���Rp礑qa�t�R+5�3���b~)t��A�y��K)�U�.��ɛ��m�<�	����!�xX�F�+��d!���A��7����#���ɜ�>g�~��N6�H�l*<�f�U�<��C�N�䪭�T`�)�0�e�����X�I�,��B��t�, ���)�����G]qE#�#��"":�0Sm2�_s��Ռ׫9�)�T�c(֛m��(��uUT�Cƍ�-"�5(p�`1�o[̔۟�rz{i��Wb���q个�n����45�'ya�h��{uM��NaY�dUe�V��7�5��iuaf�pTu�)�ͮ�oƃ(-��X�����:A��XQ���j�`�Y�!7UM�Únͭ��ƖaB����l٣�6l��E#�#��"":�0Sm2����8Z��w��xK��1A�x)��^f+��"D]a��f�n;��Ct��c�r�A����eG,�G[ ��v�h(6]�8B�D�HA�!�~/}�W n6���JH�a6!�I�J��@��8o�(ˏ�7�d�d0�t9ǚ3E��:Ib���,��!�qTE��Z2��p,��2��GP��� � l�GrK���-Zb��e�q���(�n�{q�-tb�,��Va����z��ޛ��.K=�29UW$ᡮ����.�bn,8X2��J�N�f B�(Y���13�lѡ`hzE��m�͞�8;5㨴�--8QFei�Q�<m7ͺ�׽r���xi�eSq��d�r��,Ұzod6b(5!l��Z�f1X�6�>�}[i�qDu��R<�8��"#��6�,��ǫm�1Cڢu�LugQ�=����7V�n�Sulμ���m��jͮX�QE	@�5�>2���@c��a�r��4f�85O��<���e6�O�9U,�����af&CDG�9h<զZ�ѯW\*G�l1ôA��A���1���u�w����==x;��{S\�*6R��9�aM�~�0�״ݚ<gG�CƑ��f�y�QNJ�u$gM��E�T<��E����bޭ�ya�BO|,�O�Q���S6�<��눈�y�q�x��gM��Qe�H��F�1VF�a�m��&B��"ٝUR�e�4����H�]Ʉ;E�UUXX��{�u�������y�4���v�h�kg$e��=�#m�{v����s��߰������߶�M��aQ�l=���s�@��W�I8�[΢�NQ��E�L�66͔���I3~�%Xy�ѲӴ�_|�xvl��{n�Lc��.�j���������,�:i(Hh'�>e��yo<��눈�y�q�y�q��i�Zo�3U��8ҹ��ag���m�tQ��Ql!���#�>��� "�aVf�&�I�G�t�P��-���2��ҹ����f�ن�P`Ս���T�98�!������K�`4+(��x3�/� 66,%E%��N"��d�T�BȒF�=�њa������	x��ag
ǡ��5�o4�0̲_N�6����P�4-�+�Ҵ��犩R�g�X;�ᢓ

�(�����K�~ΙW~uHȶ����-n���O<�"<�<�ͰSM2�H�x����m���$�f&���$m�I�3�c����-r�d��o��@������\�s�6X�u*ݖ㖛q��#6�|V^k�ׇx�����<jq׶����Gۏ�`�g�_l��Zkc=�ѩG���q�hӨB<�Q�sm�H���A��W!��2�	#$���G��T�F:+�TYYx�}C����q!"��/C���o�ə�o��f��<�ҧk�=�KFB�+Z--&X{�oP�)�sF�ɮ"�v߂+F.�,�
�F`�ª::���tgm�k����(f�7��Q�<!�[E&OP9�r�t�y�UUNqaгE�X@�!$@�
!ҕ�Z��9*�EG����k�Ź[kN�|&�HƃAF�i|��xL9�쀒�x�6pj��n���d8@��H�ҫ��q��㌺�"�uŢ"�yDyyǛ`��e����o.KI$��
PN!�� �y�`��@e��
�h�Q A�����QG�0���
8۳�I��t	y��:q�7I��CpkI������1����l��SqӦ�lڄg�J*�oު�w<�W���g�V�<H\c㢹�[�,� 8�ܷa�6���4�}pB�m�lX	�	���I�xs��a��{��Q��.�l�`�0�+�D@5���d�ѧ��2���+4G� ��V�u���Y��??3���?b�1����b�ǖ��e�ulڢ�g�1e�<[[l�V�<�-�4�laV�[U��y�+�1�X���Zٵ�Kb�Ū�kb�[6��l�ص��X�Z��-lZضQ��̱�����?*+�y��EE�kbUVco1��3�⭋Zٌ1kbՕ��V�[6>!��6?��?����2������?7�t��;���pv�ص�j���Vͭ�-�R2�Vƕkb�Ŗ��mV���ŭ�m��L<M�<OB�G�����g���2�E��x|<����k���Q0~pl~6H?Ç��٣�1�z<O���<x����z<eL�ص�����[�Xa�kb�kb<��0��ůkf�-�[?$<Hx������~��83M�����ƶ<l�����1��0����x�<��&�C�����C�lw����jU|C��h������a,JU��:A�V{4e��(,@�	Ӑ�́���٩=Թ�(��Iz�gm��a�x1�i��|�a��$	�ׅ+����B�{3��g*�P]	F�v-�c�f��a��+T���45�mAXd���;��:t��asN,�LP��� ���� �?����!-��g�����{��~���֦�)�{�׼��s�����9�y��u�s����ns����9�y����n-խkGQ�V��E��yyǖ�R�m�Ym��Z���;��A���g��gC&bfAbdi21/���HA�v��;��vx�y�\'K&�b1�|-�v���7y�H{��
������G�ɡSK����U�q�i�6@)�Ɍ��-�;8->ul��\n�<�x��
�I}��^K����'7w���4pub	�%"��e�Q)��\���y4���f�	c�I��p����hd�*!l>�o��-`A��p7ĢJ�70�i����wO�~�:y�w�2t�(�Z�^�pń��/����R��h�A�A���n��5�yM��l��s|�3o�O��uuWm�?�H�cVۻ�gkl��ӺwM�w�y��Q��a�Sm����[󮣨��"#�8��mfT�m�[gC��~`�J�#6wYFْ����b�oÒ�6u�hи3��L��NJF@_}�����a��>�"��/���J� g��/�gϰ(iH�aHD��F����7�I�¯$�X�=����dbȠ�����wO>��m�E�,Hi������8S�ϼ�V�4#��g���-�y�F�<��u���M�[�u�vL���R,J�z�k�I[� �4h�e�!�S ��,Hik�����$m �b�!��r�i�c ֻ7�)��eKe���"C��~�I�׺�N�
ot�:�4���l��p��n�v�<���Al�h�[ �`P�P��ݎ���[o}'���wM�TH����n��dXD�gJ0�F�ZߝuZִa���4t`���P�m���'(�a�	�bĮc�$-�N� ��b��(U�L�B5�3�"M[t�dw���uYm��f�r�T��}໋v:�6��my�7k,mۺc*��� ��ʍ�x6�`��fF�D���>���F�˱^���0��"Rӱ�P60_k�e�� x�oVa2g�ɔ��D�.��S	)�f�N�:08�06�޴��u�͞tݓyO��;bD��jD*bd��BGc��16�ϥ��D;����\O(��tnPAhcL��e@lI��0i��	*�ӛT-A[-����#�|wLђ������C��m��8����yGd�_aߎi�#%IU�<>2��؇�����]�<XS=��w��:����q��xN��ѤHi0q�ф�;!�i�m�m�t臏On=��`�D9�� �ᤠ����6�P�6|�o=�S2>�l84��{}�}�o�`p~(ᣭ%DŃH�T600���08�S믾�H�����> ��0��כ���*G6Z�9JS�n��Dykuտ:����E����^q���&m��om5���e���C>�	|�ic�1-��lb�@@�`G���D<M������<����Վ�C��u�w-��{+�;������0��m���_����x-�km��K;��C$(`Ьbߛ�Bl������"p�f���Msm9�I��Q��í�6�OE��O_�c�`��r��m��4�2Ɓ�g���頀f�����c˒	�"01�*�Y
�*S�U����zD�!d~�����L80���%�͖/st���:�`�M��l��C�6r��mۿ�����\�H�#����ɐb�-�cQTIr'�5�T�&��S��H�`�aU�Yi��� �9�E-16��>��Ｗ��ߝuխkZ0�ukyn��ͭ�L6�-����f~ˌU'Cllm�B�����K�4���_0���Z�u�EW_��B�(��F��Ɣ�	�&�3 3C҂�(a�`�I�����m��x�DΝc8qm�{��k���7���
�(ǰKm$�V��� 0- #J#c[�fm!�|��mB����Ixf~:h����*R��\wwlb@���B�.q��2�P��j`�<ʼ#z<��CF�����p�il��Y�H���7�rQcAcH��cw���>P�o$;k9�ӭ��DBss�����YN�Xhc(�42�F^sy!�o��&��Woe��g��:�u��>�,�q��tY�x<7��I4�2�*a��|�e��E���͎�W�Ӈ6֙�m܇+��P�piO����M"�1�_}�1�������-��u��E�h�-խ��<�̩L6�-�۱�F��k�ز۽m���h[<��,S5�.J�P�����<��v��vY�ӄ)�h����䖊�����d>�R`��:|m���R�ᕐc���͉�`!��T��b"��,'7�h-p����MΚ@��.�f��_�p��!��8�3�f�m�m�V��+����h �M�A��#7�%s+��Z[��G�"��^5�� i5S
V5}�q��%`�i���16}�vt��G�Ko.׷N�:X���s��KͻT`�!�oaH^L��M���޸��7dy���Sr��;�[in�8�{&I�P��<�e�I���F*HK�	|��=�{'I䇆�����<�;h0���҃
m l�iCCH�ER4�΢ߝu��Zֈ��Z�n<�ͭ�)L6�M���u��Yo�A&��޶�8��ӆ66��T��S)~��൲	�V�Kd&���{$G dĤT1>o��?),wb����{&CL�c��v���I���p�7n�E�ں��Llm�s�q��zX��9�.�锈��]%��ӹ�|�w��ʽݯ�B�sw��E���a%�
pe����f�K�.����ߑ5����Ke7U[4x�:[zC��d����<,t��K4Bپ<��q+�yG��td�҅Ѥ1���D��aL�{8�S��X��臭m����;9��6���|,�S;�����ii��2��v��KjH:���J�C7K(�kE����64����MI�n�����!Gcn(׆V�j��:��)�[EB���D"PbY��>+>+E��"6D���CA��7�J�)���vM0�b mp�`���������$|k;#��t��8��b�6C��+�wr6���-���)Rԕ�~{���n���Kp�U����Vx�X [@D����0\ �4aê�y3�)�~�IK��O A�zn k�}�v�B�+T��L}�ַ~eO2�ߟ�����"ֈ��Z�n<�ͭ�)�0��0��Llg!V��ˤ�TFې��.��lm�4�-*r8���9Ct[M�h/M��E�j���S���ԕ%�r�1Κ(|E韞:���g�۷^�G�Q��E��f�C��}>nT�R�����ƛշgz���f���s5|�
����ϵɹW*�퍚FL�� �f$��� � �iĳDG��Q��=c�i���Dh�Ç�i�� o��)#t��=Il�t2�ݜ��F���߼Fl�ލD�X��`��CKJ�5����G�-���iY�7��ʥVbGE��Fk�I(�['����v�s>:���g����� �LTy���r9��7�(j84���pePk���S�*�i���E�??:�ȏ�D[n�h��q��ʔ��Y���n]U0�qF66��h��9d-��Ce!1��޻�*��>��\�2ic��J�ph\���(it=ѤΡ��f�D��,i+iv>�$X�5��m#�2$3x�S�ܶ$�sq��&��\���l4��/)�A�0`R�V�W-�/8-Ȣ򰶞�q�I���v���V��l �4�Gl���0�_�J^��R�`b��I��8+��4��8�B��6ꈯ�{����_W�q�FjmѤ�kP/M��K��RX1���>q�\01�PЩ��V�A�M�2�wf�R����Ķ1m{���ݣ���D��^�;8�:��[:��CKZn��&��g�>>>6l���E����a�ml�L6Q��a�M�R�)�e6�om���Bh�
/�E����*���s��)%-ә�:XZ�*JʳY��Vŭ*�d�R�+Z�����[;;n��un�t��u^9�d�&t���.�cyƷ��IWd�*2��Uc���u$�6��@`�����:G���қ���L��0��#g�o����1��͌ �GƗe�)-�`�1�Y�r��Ѷ�I�j�ΘH?�i0��C0�0��ƞ�ֱ�wD�+|i���MV�b6o��uEv9��#`��$4��5���1�Q��"�g��魞�:�oV�a�OK	�~��N��#��tGZQ�i�3�L|e� ����j��i�<�-lmg�mK[[�-l[������p�ǟ�~F?6�^Y�e��0�ٵ�jykg��ضf�Ÿ�mV�y�+�꺶-l[Kf��mlZ��-V�[[�-���VϏ����?'����x~�<S�Z�W�lűkb8�=[��<O'���x��!�����¼>��0~G���mC�g����OÇ���~4N��p�,�6<oǊ��p�<M�<W�g���~,�Y,�-lZ�Vŭ�ml���ط�l�a�EC���Q(t?>>#>'�'����,�?��	�|<m�c��c^���
����&�x�CĊӌYV�ulڭQo3�eV�-��-�U��il�1�1U�i��Db?1�f?0��kb�ū�S�2�-X[�����S�a�ql<�� x����Fd'��3�g��'��<L<O��Åx������&a�8x���g�����L�j����Աb��� �}��W1�=]����ٔ�CU�ꍓ<������z\9S�"����Ic�]"�%>ΒGT�k$$+F��b1�V&O*VV�ꊟvEz5ӈ0Ť��\p�l��\���TY�{,��CHHwm���2"~���<u-�/o���Fشڐ%̎	� ��1Zsf"�:c��S��շV#�$W�
G�_��{9F@�Jdb,̘�$��)
iꬑ�ሇ�3'{�.z��
^�
o��$`�1�#j$b5@� r"���R [�t�^u9��DP�r�=�-�N�[d�I��m�䌬���qET��}��˪F�z��l�d�Ѧ�����YC�]Aڥ�2-v�NB咜u"+EDimBR����JXxM����5(�j������t�2�'*�m�8�lm`�(Ӏ�.�����	�b�=����n��0�t�zϮ�s���u������yG�����7W]���Qe���Q��v��۝�xrn0�� �v����Gv��[A���aj�Mc��2'�o��݋�wlw�F�h�ۧ���K�W~�[�{�'k�x,g�u��C����7��]N2;aj�g=�X���>�}���9�{��ֵ�z��s��9��{��ֵ�zƹ�s<�9�87�9�k=u{j���$u�V��-�ֈ�#�6���Q_��('Q�q�"A�\,Ec��>���8I�iכa�_m����V�*E�����^���.�n2�V����֚�|h�9��[��Hҡ�ɃvW�z���v�s�<b��w�(5�8��<h:Ch�Zf�]�v���{l֎烷=Nヶ���c����K�#��/nS�ۍ�[���ݲ�.����Ů�λ=�6��l����{~]����nOU�loT�e˅"P�S�0.�]Q+�PY�+��ܷ>-�����>'�椐h����ۖ���\>RE��[�/u���)�����o����x`�)��Z<����їݤ�c�JJlp�lp���1\/��o���p�ᤰg��x��16�cD`xi3�Ii�H����]G*Kq�4Q7��G�ˎ�͎'H{wyA�\G;�n��
��1���c:2l����9�%���{KC���f��r����"<1pghh(�gT\�c<a ��5��v�uUP�piyQ�4�I�Hٲ4.C����c ���1��b�`�[�
����"4`FN@�F�\I� ��~�ne��`c����|3C�pf��j�
,j��8w�|���*�T��:2趜Dy��먈�-�֋Yy�eJa�[i��ף5�g��0`�2&`�5��gHDn�@e����kg�m��zn%XB� 0b�p�d Y�ŝ�7V���=[�n��B���=�([ZaAE��C1_�������*��͕�>Fem_(���?\c���}_?��]mJ)_8��P�^�r2s�Wr�2�w���".��wF�+�v96;�p�v	tg>�s��е�B�Ҁ�ȍ�ja��͹N����B���,��A��d,���L�L�궧��og���ˎ�l����}�+>}��m���]DDy�խ�8��*S��B�n��֟Dݵ�r��@ ��ѻ5�7�и�Px� ��7�1��!)�q�@�&2��l�m��G��^�,4�7};�y��6�0�FG%� ��xa!�&E�Ir7����cZP1W(��n�)h*�־�Y$x�]�N��ƞ9����<A���(m���(}4Y��Ѣ#�J]�9�TS�d�hra��J�T*L�K��z9�7���{���U�t��T���2�`�F��,UwJ�ο}N����b�3c_��0{ncꆎ�a�g��u�DG�G�V�Z��6�&2ae�a��u�m���	Se�66&>�ѣ�[*��:u��.�9a@�6�Ƹ�_(��h�A�}Z=W����*��I�X4�I�R	Ϣ����C�_�D'��h�$�-��������ao�c�_��e�^���yR���4�@�aZ�
F�$�lt8O��c�0a�P�ٸ{�������y7�q�gA�O��4QK�4s|nh��ޚ]>Q����~o�Li�LJ-F_*���<x�]0�����f�U����{u�[E�"�u�DG�G�V�Z��6�*S��M��/4�HBB��b�a�B	R#1���A%�r7+(����n���/(#�Ra�Xˀ��fbMH��N�t }o�����V�397a�u����������3�ǌ�"2�i�ۡ��Gy�t(_R���I��hϚ��oK,�ʂB.:�������%֝���5�zv�oo6�A����i�ߩ��M���u��E�tFۇ�LTB�1k!�J�z>8t(SC���CG�(��4Rl�6үvI�~;>�Jt����I�3Ə�Ѵ1�}:e��0�i�p�h,2�����m�ghgP����M��7"��%�mF��t�d��4~�"#Z'A�
���6Y��j�/��*�����\Z:�DG�G�h���m�T���m���R�9Ũ�D�ۖ�:�4@��|l�Z4V֌[C0a��7}>rF��f#�ۓa�lo�cVx,Q�v���m>���W8�*������)������c��m�2_�A��	P�8��4�d�F�+e�����xl4!� �|YGZJ��r�k����4�u-����ꓢP��;�u*�_�K>����}�s�q.���X0�c\G��s�7*���aj-htP��X�]�tР0a�\{hVo�|�$,�٭q2e�֝G_�uբ#�#��ȵ��m�T���m�����Jb`��C<C��U(VX�6Z!Z�%���	�]�$+X��!>7�GA���dC<�YH醎�KA�ý�$�U:q�:�T��FK���\�����|Q��P1�6��2�B"��ͺXX\\�
��>(4ogB��1p�e��ϭZ��d:4�t��f־��Es�A`�K�&���l,�C���C����/VԦjl�U{ܶ�F=��Yo:��-oκ���yDZ-duq�a��m���R��V>�?S7MӦT)&3ccb`��jo�R�M�WjV��uZ�gN6\,P|��8認��{�Tn���g���;n��� ?m�t�t�gu %����w��Z�g�#�h46C~7�_Y���Dr����}�
�/[��5@���8F:�ǲ�O�7,á�y�Bژp����b���(z 8a|oA�`�C�E��d1Y�>��QG�˿~{����͔�y~G�]ukDy�GQ�dqp0�QB|!�h�!�
��啭'eq�j�")�<��=w.저l��m��[m���V�#�kqlG.��q��ν^zۯ��(�ݝ��ǭ�q��Oj}�[��[k.��666&/խ6Q�s^���׶y�]�w�xt��XѬ��4�)rv2[��h�us2���^�0^���lUn����g)���n����,X���>�|qmo{|�uUGgrR�gJ)~[L���}_GQ�:�&Jg�m�r�7��R��k�^7��t0D<��x����ܪn�0�P�0g�Um�i�g|�+�>��6���%�+]~>�ٺ>0��{]�p(��6��e�#A���G:����"A�6�� ��3d8�P׼�l�l|�b�o���eB�ϓ��>>4|t�����Z�y�y�8�6�0�a=�3l�?]pllL�х�k��,d8��G$�*͜�G�%	��(��o˻�f������Ųݸ8�Y�@`�MW����Ε
h�ֆeh<�SĎaЮY��ތ��r���'YQ�씌y����)�UJ�:�Tn�n�����_t|�z��#gK> ���Q��L�y1ʯ3��7j�W�Þo,�C�7�P2�������mճg:��������Q�Z�c.���:�W��ͭ�q�^*�Zص�kb��-�m���~c������~~1���űj���Zakc[8[�ٵ�ט��u�[[[�ٵ�n�kb�Ÿ�V�-�-�2����kcǉ��~$~<W��(�n��o�V�u�Zf�Ɯ[6�-��⭋p�����������:OP�>��{<F?c�?Ɗ+���?7O���t��x��O'���<x�^!<x��,�,�����<y�[�[�ٲ��m�6�)l,�(t:<F?�!�����Z0�|O�|V���m�`ǡ�|x��c8������8ݓC<����x~O7n�ᱞ�!^<O-�U����F�0���~~Y�|O�Ǌ��x�����?O����pg���Fx���&�h�(x�c^ ������<O7�
��z7���<���T�<6<<O�ǻ���OuW�[-�\槶|�z�k8RƄ$!���:���rl��賷X�91/���H���@�F�NÌ�F2��#mo���t�y#�3�cs��N�<�7ӯ��!ة�P��("��,A`���'a�+������dz]z+nBs�P�I9��Ժ�-\���JA\�p��1LUk�o���?�?$�%����d�\�ھkZ�y�s�z��ֵ���s������<�5�g�kW/._\�%�w�.Im�GQ�Z��8�,0�m�ڴ�6&�dV0�*?�Ң'=9^���K�qsFVf.���u�l�`τ���X��GD*a%3-���������fe0�ɘk�tJ�GE2�QԐ����֜Tɗ�����l��4��@�ί/��Z�JE^����e6A�f��K�9Ќ���aH��;ç[�٠c�U��mh�|o�Ş]6`�c�E7]6a�}�Gv}R5�[��1�����t�_���գ�2��~[��:��#Ȏ�ȵ��q�Xa��a�k����+Y�J�\���1�f�f+8s��;�s�U^+��(c�Ɠ����a�i�EF�1��Q�q��;�ܨӶ:��~�'�?�ɭV����gJ,�r��1�f�
>F^�J�C4f�1�g��]1k�QC����(ln�Z(��$�� �3vW���N3B��Ɠ��q�1�`�JTI]Tac- ���Ɨͻ;M��>}�9u]��R���i�ږ����FT�<��a���?>�����e�G���ukDG���ml0�QBg�S�^,�D%���k�8j�LP{�#Q R��	C

�I���-q��f�*U�I�bx떲��'#t�C7p�R��J�O�Ο���֍ɣ��3���-�*꬙;s��$ͧ{b���
jK!D�*�P�|66`����Vͬ����~	��C�����-��~+ۨ��ֆr:�o}3#wm��Q���Д�2��l7x��>��GU]�p��c6�QF����>o�(c�S�
/�)�
⥟,5�81�c>�6��
m�g�;����[jR��&j�X��ڟ��
:1�c��n��G4Y���V&7��ע.-ѣ�u7J���������H�����oL�:�VPㄌvT��l�(�&`rV��~�@�=`~g��@#�&�m^��2�1��
�XW�C��-�mn���<��#Ȉ�ȋR0�
!a�0ⷺr^����KD7�}�<p��@��T�!}�U���#%����I���E~�����a�~��iy�?d��pa��0iu_��D����|Yj˴�,�Ό5CHN�����
6����6jQe2�BG	E]6��F�Y`�_��#���"�MX�TAԪf��v�C�0`轲�'�c?i�W����:��a�O0�v���o�uZ�u�/δ��o�<�ֈ�"#�"-H�8�,0�!��o҇�3�c`��/� ��e�ogL_���5~rv7�3I�(�mqmY��JY�3�f�W��0���P����:Y�������c·߂�):��7"��Nʎ�PRZ�?��R�T$�g�P��-�Y�7�CX���\�U�8l�9�����I�G�tc	�ڳgK>[P�	�ы,��,^(,�Ƶ����4TLe�a����YT��FϏ>?���1�0����.���&�H��
:qX�ϋ0Z#����[�<��h�"<��3�0Ba7�r�6SM�fhll��Cv7�^s��T�����[��)G���wl�~���a��~��"�q�j��Uk!:��.��+�4a*��yzxݞG�Lg�e��7�dr�3lm��cx{��#�ha�tx��uMh�|]�0��8O���ëƓ��Tݚ����n�S*��AXQ�Y��t�U��(�3\6p���a���7߾�*��C��>,��QL;��Z[�yh�:����Z֏"#Ȉ�#h�l����eM��Rᄧ�]����۶9.@yn��m�tэVF�r�V�P��n�맍���}ð��H�i��b��2l޲�
*s���ۍ�sz��m�gr�V. �'�4��-!�A @J�>o�����Dt�`�U�6f���]X�ݥ�+u��,;�=Q�mhf��_#��j�y��"�c\�g�G��!��E��W��������|��A�k�+F�������>E���C0���m���T0�(�rI�p# ̶��Hl�C~o���a����=�{=��0�)��.0li���t{�V7�L�B�1��}6>T*�.��W*[#��T�[^��D&�g��p�сp�b��0��g�C�qK��}E�0f���~~~G�ZִyDE�F�e�m�_iT�&uY�Xk]4\���b�-&`iC����a��>��$>���.4!�ó'����cnήB��&�}�:t�Y�[i�:7�xi&0�:ۤQ�y�=�Gw��q[0�є0�C��9�����P�;_eJ�%s���rF\L�cD&}��F�)	&���(�:0o��բ0�,۠���[�p�}N5�f��g�ZY��F�����@�p�\�8C��i�_�hêu�~y�h��Z�o"#Ȉ�-�m�Xa��a�2kCf7P����Yc0���5�E{�y.���ts�Žp�
61����Or6˯90��e0�p�γ�)ʓ��
4�ΐ����tæƴ�1��s�S�Wp��v�1�n��箠Իk�tU®��'aG�6���g���`�Z�d��&/��V⌖l���(|p�����5�9�6ܕe���W��eOaC���yuE��QѾu����wr��p�h�0��2���U}�i��N8�����#�-kE�"<��R�F�e�a�0�޶c#�i�}��Mxll�-�r���l�����)��2��ZZ��#�:�mGX�������i׃�^�qպ���UT�����, �d@���QN��41�,�Z��l�M�ų�V�̓j5�K��ٲ5�"�f�4�æ�������z�n���a�����!e|�Q7�6��bƈt�0��R��L�E#IXx��:x�˒��K�$��I)jIF��Zֲ�Z��ԷDR"#(�#N��8���"2��$��Z�^InX��J6���"#.��4�<�4�qi�Dm���6�먈�h�����GI-�R�I$�KIyb��Dm��a�"#0�")ƙeqQ-k[L����en��IjIn�ԥ/$���I[���6��-h�kZ"":��DaG�m�qmm�!
DR#$e�DG�DS�!�#���;��*w�ǫ�OE�����$��
$Lh8v�!m�A�-2� \����"�y(�B���yU���W��4U|�3�&h%(+�K�&õ:edY�<{u��)"�M�&��a~�ë؈�̬��B�H_'+�y��rs�ĺ��X*젧�F;��0G!\.V�7$޵�T�L�$�E��K�3֙�3�,3�T ���E��,B��XԳ,X,RB�j�`��}�_C�����B�t�����H5Ǖ	**dQ�٪p�4��In�:C�D�n1���z�������-�I�.I�Ja��������Q�L�)&i�g��)R94&Z���{!&�C�1	���&�Z��Qf
����
4$�O"���@�{��}a��x����-!�,@��l��w��*Ck�St�JZa�+p�^T1 �>n��;Mpu��&A�:�a
wB�(�<�`���V��;\)�p����&�IQ$]r9���sWn�u�&���}��F���󭮺�TMc{��S�zŵ�v�V;��S�U;i�u�s��G��xN��g�5�naz8�2Um[/}wn�q�c8�����v�k�/<�u��v�E�kQ��X}0�Ůk���P^���7\q��]�ؐ�"Q@�$�	�Tp���û���z��ֵ�\����8do|;�Zֹ�s�����kY��b����-ykZ-�DZ��6ڈBa8o�8�Tʡ�uR˭.�.�Ş��+7g���j��
pOA�D�I�u�.��w;�j�vܗ��k��x^����x�3k�m�����:m������	�nK<x�k�x���m[�y��=����E�x_iq�y�ɋ|G a�9�^�@��6�����;���n�7i��4��cr\��onz:�n6;Svע7��@�n��q�N�\\�.۶-��*�`����s'n�רn�\v�ʶ���U;)��66&h>m�6"f�􌥙h��	w�]�.�H�ȸ��K;ZGR�v�k�0�W'��"���f1E���uӾ�Z��|��eA�!p����O�~����.(�J9�5Y������^�d������be&p��l�E�0�h4[<C�å�(�na����$�������|�p��r�ǜ�e�R��V��kJ������G/N6Q�~	��=��0@s_�<�;(�-��`�lt��v{�9q�K/����m)d3�1?�)�UVm���^�x���a`�#�x��c��U]+�)���^~G�Z֋Z"<����m�Xa��!�[l�G��<�5���tllâƴR��[H_h��3G��CbŢ�m���!�1�)L����8i(��9��C�d>��F���>(�(A�y�B68�}E�F��cD�J�!��A�{~*L�nꋒ��%�r�[%]6��WF��s8�֍����z9����(��*��`Ҿ�q�^Y�4g�b h�a0��R�X�������l�K�6֛W�S�6�DZ-�G�Z���<����m�Xa��a���r��i�6Wn����c�{P���|mR�p�J�]6`�\8ۻ�ӳ\(����t��ٰ�r����A���>�`�����HX\H���B Dl7UV�Tu��ʽj�K��CJ���,d{���|q�C�S4hf(��>7���1�ܓƗ��6�m��p�AчA�>$�3ƈ��&�՛%T�Jψ�4:v�����C�Qf�+X������8{@ԏ-ku[�-h�Z֏"-kmm�a��mO���u�W�1_��{��;½[	:&h���oF>W��`ǡ����Z� ���� ��8j@�n�\?)l"�K�4��7Ӛo�N�XE��G��1��u�"�<b������!hc�eC��Y{��<3-|p�����,a�ڒ�ak�-�\�=T�Y��C*)��ʸý�}>�bUs�0�6y`�'|��)�-�p ����������jn��aiל[�ȏ?-kZ��DZ�F�0�QB`ߤm�3-Ca��0@�Æ����km0)�W8�p�v�aÇ㱧�;�L%�QQ%�[�4i�� �̓d��2���e�[��u溶�z�f���e���v^]/j�l퇮3]l��Cս��۵��j�^5��x���A @�̲�"#���,���R'��_�T�8�ڮp��4$�|�^�3�������u�m^���
�n�'+p4���@��s�-hb:���4X���r�0k�J\�dR�:=C�2��P�.�kM�o����NN$a�h�aK�}'��Dވ65'Ŭx�E�⣦1�pуt�K�)�6Ht�F�|3cu�Q|�ґ�8H1�+<z}W(��n�p�
A��!Ob
9���� �����Q[e`���������b��j��a�\G��#�Z"ֵ�Ȉ�����0�l6�V�6�������Ϊ���4qEe*(��KB��F��o|������]!T��li�}���!��Ō1|�eP�kkYf�o
}��O��KN���>4��1�0�S,���m���ս�PGd��vԼ)˸NCv^�??��}��|̘�9p��:�k���H�ٱ� �p���E���]�wuEIQ͞0��t[�N7gv>�ٳ_7�_zO�4r��0���qן����kZ��DY��YD!0����Hm&67;T��l�q�J$^������`il���:n:�m襢P��(��(8�`�^X۳G'���UMxt�����6QC���s�4H@�� ����Z<}�4D(���8ȋ����������ڥ�7ﶸ0���-湶�X��q�����۩Uu�������ڝ�0��~�i�}���Y�C���ݖY�닅�5GHQ5c����a��~e�UQ��]2�,+�����:󨷞G��E�k[Ȉ�����0�l6�)���mT�0a��ŜӦ�w	4nF�ea�V�k��ã�{90���7���ɜ<�ڀ��3��	9���XLr��z(�6Dp���&1�7�����D3�CD>4Y�{ZF��ʊPo�"����h�E%��TO�S�7��O�v�L����n�'"��n-�6A������ٯg�^�������Q����b���v�S�Z�m}�"��Σ����y�DZ�kDDZ�F�e�a�0��9ˍ��gZ ԹM��udF[ ��C[a7eAp�(ʄ��
M�V3L#AM[��YU��b�	��'�JK�xن�@�$���&��0U!*�$��b>��p[��I^E{C<lu]�.��9y��nv�(��~݇����˒6������2�0�{㈕�P���!M�=���}Xl�Uv�S���H�"��$B�o�鹴en�(�v�tzzO��x ��bi��a��?eJ[̷�$���%\��{�����V��14ё��aq�Ңo��䯌=��zJ�(��Q&�\n�n|�&�t�k�B�c�e��P�1bϲ��T�o8��4�F�Q���\��K��w�~a��;9�GP�����Wq��[dr�SqQNH�_3G'��ϗ���l��B�M�!9��>�|޼��k8�W��:�?:�"�h�Z-h��[h�L��a S�6ؓ;�#wpcaI�m���M��N�YT�$�,ڇV��\��K�{{��3���]ԕ�C�(qvB6p��CǡC
F �������A�E<��xo�]W�èӧT��g�sM���f�(a�}�Gi�(�Ѿ@�>tse���,(a�n�=�nt�)f����t�ʔ�7N��(���	$J)�{誻��w2� ���x>b#��/*U�>!0bd[T�p�0�ˊ6�R-�QJ1a�[��DY��<�:_��RD��9�W�_��w�u����#JI/��IbԒ^ؒ�<������ah�Z�m�]u�DDDm�F�%�%�%�RZ�^I(��#N��4�<�"#HR"�B"#/#h�����-X��%�$��I%�ay��2����"#H���6�mB"0�B"�a��Q��ֵ��-juki�ZDR#ȏ2�)�"4�""8��G�m�Z�[�Rֈ���>��"0����6�8���6���aDeGQ���,��"�U�|��U��?{_f�-����k�jQC!~���,&�)��R �����dͰ��&K (y�J!��NX�e�j�pc%p�BÍ�ɋ��M����F��!@à�t�Z�"���s
\ӹYW�9�T��3C7��n��q�h�Cnu���c-�$m��(�ʦ7O�d����f�n�"�{j6��.s.��q��0d�m��q����d6�>����rL����O�;��:_r����{��7�k\�9� h���9�kY�9�s�s�7��oZ�}�r���v��\�+E�-h��"-m�m2�6�oʴ66a�i�{4܆�����k_j4���g�8��f�k���eE}��L���	Qy��#G�(�a���4i2�9&��� ��q7��HʪUS�B���F�R�ձʎ���D�,�uTQz,p�z)k���0��$j�:g��ʔ�3�c����#*5�[$e��`�c
��H�q�C�c���@�<�0=�F�84� ��6�wY�2N�paBh��E��ky�$0���i�[Z<��ȴZ"֋Z":x�L,��CS��(���qFq�G�A�WZ0�+֍z�6W-��%�<@��d�FcV�xP 1���2֘�	��F8aDC�~��G-��Z��a�ga��0��h�Nm���z��� ��7��gs�cZB���vG$���JG��0��`���j�|sQ��g�y����[5Ce�(0a�E�^�I�(�۪���\0vE��S��V4�߷��\Fa�_�[���DZ�Z��Ѷ�`�P��!�$�R���D��
�~�u�������^�A�:��[i��?}�·��&8;#Un�d#�\�ɜq�v������Yڡ�i�%:R����Y866aE6c�砤����o͞�ʯ�ې��ͣB�ޘ����RE�<P��!��:�E�_p��ｏȍ8u�;S`��e-h�D1}����(a��3��ߚ�_?�\N���v����ah�(��
7f��W�9X`��i�l���s��[j�A�c��>��}P��K�svLcч����Y�����d��r�n���g|�t굣�r7C(�oŪ,�(a�v}꡽��Aӎ�ݷuM��N���k�$����_n?;�6������߆�4X�)m_i�g>�{��g��<��u��u�]Z-�����"-m�m2�6�qSNE�
���5���]�TDc>+��xai��~�<�UPYe||t��1���{��D:��#!4�0�ע��۠��F}�_�r[�ZnQ;����f�|f�qh��ϹNU5����0�ӛa������]���MCϔ�f��rF�b��鋘S40��B���p��r7���|,����m[��a����_7�t���m�����C��-ƍ�y��>��Ɗ0���]Zߖ�E��kGh�!0�2*RG$m�li��z0���J!�:l���%aӆ�(h���xkj�;�u���aG��'#r�a��a�Ǖ�C�ϓ(a���g&�wd��"���/smv	\�j�?�i��6\�eՎmt��J�(Q�������eq|`����$a�ã"�(m$��Q�aþ�̟I%]��h�����۲�-�Pta�����;���~�5����iD��6���#a�;�ҽ�O�m�~[�����kykZ"-h�m0�6�l���SQ��pll�H�߽ں����%�Ç� X¶��4��i,߆��p�DUc9$���� A���Z�d2^���9�DT��0@��c/4?����'�6T��`�6Yfsc�ȳcv���U��E+-Q�0�x��a�D����>,��rp����"�Ep��֋��N�hgF�P��}2C���7tl�O��12�f�iJR���_�GV��Z-h�[�Zֈ�����0�m�����(�YM���r�B��T펫W���irQ�{B�V݂H�$\����)J�����D��e �g8�7��U�PBcnz��jW�:�"9���N]ҏ.w+���~~�n�SI�{ذY��vߘ�W[,��%�s �]�$�U&h�	��� ��[�m�s)�;Պ ��-��h�>7 �69
�A�x��h�5�B A�(B�y�����~�ffe�kk�V�G~�2���Q�c�d�e=�G#o�G:aZF��Ų�71�a�to\;��k,l�%:t7���F42ơ�T�l�՞=��e�޵$��*�V���}�d(6k2�F�-
�/���X1����~!��:�@=����I4^�t��ѭ�Vx"�l����4���ra���D�R��P�Y�������4γ��i��~e���~uխh�[�ZִZ���a�m�
4-��:8:��F���:��6ϴy3E�t1��N��h��;o�͹u�)\����<�O���6���f�!
��G�UL��L+:�ì��?j�8��s&TɧG�3}��UU��̇�o6ݛfh�����W�����ꨨ]�S�`�k�'�����m�y�����]y�:P���ޑ�D\:C�
f-yY����!N��G���>��V���5K�7F;������ٱ�5��C#�6�T`�>8Q���u�h�DZ�Zֵ�֎6��0�
;n��a.�Ccbc<p�!cZ0�ᠭ׌6&=���f��4�4C�/�Tl�QJ��P���2g��x��ϟ6����GD�n�T-�r���Dh�cq3�>C:C�Q��,6CM��ge�!F���9%V�6��<=}�p�
�H_�Ѿ�P������Kc[(ϛ������&Y�#��"+)a�+�$�6Q���Jm�ň�x�1���e���uבh�[�ZִZ���a�m��_�ʿgU�a�FD�-����e����]7E��Y!�����0f���j�+6ycoQBh��8�l�9~լ8+D���,�qP�XmƳIbuws�M��ɵAA�4E���Z�s�ل0���-x���n�GNp��l�+�Q�>4��QE�,|���g��G�x��&����d1�!=�ߩ�L��tf�몕_cr�	1=|h�ء�#D<E�>4iy�?{�bц���4��DB#�.�I/�$��$�גG�GQ�#�[+[�Z��T��u�^DyDGDF�KrĒRInX�I%�4�<�O"<�(����#�E"<����:�mRR��$�Z�rK2K�nK�.�$�����I$�"#(�8㍴�)�aDS��""2�2�R"4�škS�[O4�ֶ�GYG���DDmDF���#�8��[�-l-h���DF���G�yy����a��#��4�"2�#�2�)�<<<:�,�vw1�˝���:)�ℜ�F��v�"眓��yD�%B�e��T����%˰�M72W���9��{���!x�'R��̜��nu��K�Tu�G�[$�.�(>�E����6Vs�u�D��"Z�6����C�Z���W�
��XFbŻ&nM���"Y�(JQ��Bu��d�k�yF�����P,$�(	d����ua�x3J�]Q��
L�ow(�Q����3a�Wt�E9�(iJaF�9����?oc��/cv���(X^06�v��ő�XOB$�u�/X��M̓��*�E��E�<�#�n��3M-l%4��FAtj�@��]�u�5 V�����:r8�]K4�A���n�m �W`.�6���%"�=�v�
j�[^��m�5$�A,,�'(@�L��C �QG�PZ�i�J��C
4�5[dr�a&�1��u�	 � ���C�_b�!�9ӻ�e��]��nJ�{D�%Y�3��j2#����W?OGu�a����$Y��]Z�+qC�W;����K��֨�׎9�u���W'��o\�x�/t ��ع�vv������c{��A4K�`�;�����8��qp��ӺZ3l�Im�m�O9{V]�����&�gm���c4n\q��� ��-�����3g��=%��ggp��n�z�8�n7�i> �u�6{�q�&X�T����N[a��w@crr�/cv[I��BFJ�PMy���}�ph��˟g9�9�9���|���<�9�`���\�s��ܹr��vﯮ\�-kykZ֋Z8�L0�����F��Hb-�1!8�ocr�a}�-�Ɉ���m`d��5�v���uq�����n]��/�ur;'1c�lU�x�H����m�t�g��hZ��[&����W�mk������O���W\v@�}�������ƽ#�;XGxyO2�m�0ѷ��,�&w�,g�A���X����8{����Y��\�ŭϳ���mh�WPۇ��¼7#�����8	��EX��t4�!��ea���C�D���3I)%r��L���
�2ȶ3-��ɫ�����ʖ��w�eUA�6��h������=1�83�Q��D�Zm�6, C�V۴Pδp�c
1*GZ[���V�G�=�E CGjWV��A���|ē\mc4h��Cz�	����wC��X��h�XaJ�~5f���],4|�yH��Qͯsn�u\��/���#��<[cj|��P"u��|,|4`��}����Ţ͚
g�R�i?�z5$�͔t�����u������kE�m�a��m��윯���lX�M�dJ��C��D�lm�t�¼��)1*<3}|rK����Z�a$�p�����o��JKࣧF����Q�����Of �W��a���x=�{��t��J9^�&�xgOn�4�.�a�L�d^�λ�N�
��}�B��ڶ\�v��3�Iݽ�>ֽ��u��i�8L�7���(�n�ڦΚ0��ap����?������̊���Sbz5�o�]cI�U~m����]u�h�ȋ[�ZִZ���a�m��gt����kc��lmؙ��g�O�7��m�
81�)4l��L堇<�۝6adϬ��0���1���B�2p�˶ҭ	�j!�F�ťȘ)�::>!��h 44b,ٳ�f(��?!�>+��.��,"�i��������U�ա�>����%��ݚ/�$��e��C�~�kG�F��:}��˫S?"�u�Q�~G]Du������Z8�L0��aK�	$��\�����m'�cchf;����D�8�NF+]�0�j�7�+#��C�T����� ����Q�gz<'k��۫N�7�k�q�@no�4��xg��}n�y�-u3@�h�pa裏�^��~��a~�1��eo4�?S)lL٧�j���y�6��gU[�a�g��!`�pv��6a8���J�����/��*"v2�u֑����<�Z�Z֋Y��MYBa�\6�s�^w�T|��g�a��m�T�X䄔)�K*�6ւ�"âP��c�	�v���n�����ǭp���G���N޸�\��M����'�D����۶�n������>����=l�����8 s�=X(gN���Y���5
�⧮GT��QJ�����.{��zk�ّW+n�'p�dn2�B�I�cH6�/+��u�.5�aOw�~t~L������?4��a��6���������W���f�VaA�xc|���|x;��<{�����0��[�ߛ����_G�tD\Ug�pc���\�n���Ӊ�D˸�.?T�c^ Y>���r�l��Ai�5�& 鎴*Q���9jF�Zɦx�ь�t7�������������g��>{���}���i�~u��uy��h���q��B�(ȭ�#D�cchf+>C0�ǆ��_S5���^��ཟ7�DpHZ<�E�$h��cF��"cp0ٱ��s��>m�Q]�RgO��J����Ç#q�QA��cY�*8K�q�*�=�<���.��\�:WNB�Pݳf��@�-(PR(g�P��M�b{�	��i�_��_����3pҋ�4��A��o챨�J����uKu�G�uh�<�"�Z֋[�Gi�a��e5l�4W.�q�^��3ǆ����tp���x���o��፹6�Ϻa��P� 3�����e�񄡶4š�T_K�ӥ�<m�~��ݪ�%d�z�v�Y�K���c�[xC�>��9�x��B�$AG�(��ݞ��.����v6�-}���`�ڍ�%�É	>����\���xi-�ţ��3�t:Z1olcOt8����[&��ѹ�?:�ߑ�V��ZִZ�[��,�!0S]kCM��U ���p*A���H�!��֛ؓm�Z!�_9�S�)�ލh�g��N�p� ���!�Ր��iݍ�UYy7��z�B
�GEnUUm-TY�E� �*4Q9��9*�(t�;:l�\iuFZat��S��Ƙ��U*����-��c��{�(� �耜������0(� �Żn�[?��S�3����B�|lgM�փ�<�-��ߙE���ukqyխkE�Ŷ���0�l6����,5����!���1�Bd-��N���\����a��P�s���ђfB��R���<A�b�J�����>zz��LqJ>��Ã��'�I���>��2��u��o;m�5N�=:��#��C�$laE|�2��3���R�|�QGS<Auf\K^,@-!��F�I5��,t��y�>��aE�e���8�b��8R�<��\�t٢�>�g�B�Ɨ�	-�F�s��N�6�h6q5�n㡲8�>�9f,"\oj�A�'�^���684��b8����r��h4h�J��
�4����%�\�r)R���S g�E��"�B���nϞTMC$pZ&���yMS���QS?`��b1�r�I����y�T�uD���T:�F��3�6h�G�"8�<���ִZ�[h�L��a&��V�TS�7��`�Q5���Eߩ�Ϻ?.�|f&�aa�Ͱ��F�g#����E*���+�Ey��W���v��h�ﱵ}�|n͖V�6Z���7��SM7�68�kp�=��F
ܓ,��I%���D'b���'�/��w�(�������b�՞4���95m��3b@��:�����(ↈf�޻%S�ގ%IR�It�u�\u�����)Da�Du�FP�����"6���FфDD[�:���,-/��������I-�DDa���":�8��<���Da��#HGuu�eHB��Ԓ^ْK��$��,Iyww)$�I$�^�Ѷ�eH�XauL#,0���4�qH���)�"��[o2�ֶ���Q�!�Q�q����#�<���֥�kDDGP�DF�Dq�uyǛG�mq�!�0��#N�#/":�(B"8ƱF�S�u�D�u?)U��ʃ㲌�-{ ��Q�$X�;�3PdLyn�t#ԏ12w}���^�4�V��_�1�P;���}h�DF�^6�T�D%$���{N�Aݻ�Jk�|)Y8��M{t���,E@�u�ہL����B�U02I4�A#.���rU�i�DLM�6��t��!DM�����Z�h�w�{]H��#�"_��/���O}�������˚�s�s�� >o{��g9�9�� I��z���{ikZ�m�ukqyխkE�Ŷ���0�l6�H7�m��<��:�l���7�-[^����Ӓu����?��w��tx�P���#vv��ے���wQ
��)������[�p�߷1��~�-18��0�H���C0�[�
ЍJqk�+| ��C��2�+���m����4�<otQF4K(����c��$b�J�iuxcTR1����e]��C�����?S��'2���q���뮿#��Ȏ��֋[kmi�a��`km1��bU=�2�+n���m�<A���q��L]4ZaF�{GHlF�*o��ڬV�:�Q/ک���~5s��w��E�UwE[���uJ�<z�������G��S��z6Ot:z���:�w�Cf�AJ�8�gѺ7�$�>(�L�tP|����e�&�pݼ+ꄓ�v���f�tx��7���|��i|�Ԧ��}$����lՕ�J��q��[y�u��my�Z֋[kmi�a��m����)�!F;[D5\i����q��v����k���M�#�'�-�:R��B��+��.���qz\^ls�E�t�@v-��z����ݷ�� g5\�m�d�W������q�ݜ.K%f	�9�M�J���Ҧ2�=�&D8J`���ăa��};�\=5��܍m�Ʀۄ�w����p��U�,+�R��-�Ey�s垇N*4Ec;�RGa͛n��{U-�)�J��?9U_)�x�9�0�����_O��d���c@��-||���t�E+�E=7��qڕN[g���;����t����	b=y���(iZ!��Q��yl����u�^F��E�h���ѶYa�m��_|�~Ǫ�t��^b����&\�Ư�m�:%m&���Ht�B.���l��ׯq�>]���p��M��x���Q��I��[D\V�ᲃf��D�;Y�T�W�����4�O�l]�t���x��ƕ�ݜ2��&�c%m�:n�z�A��<m��sw%�\��i�l���a
[��x�۲*TQ�YҸ:6��Y�tsa�a��_r4���6���uז�<�#��Z-km�m�Xa��C
)��I©�f6�E�ȷߚJ͐���#�,L��G���J!Q[N�T?h�>]+�$�͸2=�'�6�}�~w��_�w澍�S}�c�\.�`�N����x	�7)Si���9�����г��ç���p��gi�Lie
P�^�
mZ��a��Sv�{�8�46YСoe��h��R _m�h�v�饖�bI4[��x/?�E� |�Ee�~o�H��Z8뮭m��":���ֶ�F�e�m�	ڽ5��T�6�Yv:,�ǝcfK�`C�,���%V�Y��8}oG�N����l����3�ސ�"�R��e��ט���Y��F�aAE�>�Ԫm�S��|]�I��Q�D���H�nIa�И�i#0ל$8tٲХn��.�"��ho�U%QP�Q�٥�w��]��6(~:n�۹$�wu�#�t�}˲}��#�?<��㮺����DE�ֶ�F�e�m���KBM4��q��
V!j6��c���"k��e���)H�1``�e ��M:��FQ5��2I{�v���uVӨ8��@��v�4�,gg�; �����_mQ�k8�yۍ#�\M��'3̒HH>��q�t�8���vÁMi\�e���GΙO\{m�c)��Iw�)�Q��J�n_�Up|��6?�D6�aI��ou*���t�h���7&��ߍ��5m�f��I���yt�h�5��奱�w\G�E�m�ԣ?y[
l���#��R�N��qW[�Y=�L����%ˍԐ��4",�H�����d�m��h՘�_̶�B>������*c5�}Jc���u��]uh�<�#���Z��h�,�������m�=ﾱ���g7�t�4\N�bjkZ$���ͫ-O�[}>(�'���p���Ў0��ɘ2.&��o��h(k_7��Mk�(�g;:b���p6=�+!�㼆�]f����~%U�mhD"��l15l�ݻ�Qiݑ����B�;J���VC�8����A������F�<a=J}�T�S�٥��{ce�������?":�㮺����":��#���h�,���ßsj�2�:�8�r]�kG8�lՂ}��)�����\�skCGNxv���l,�Ԥoi$YQ�&��-�hb��<Z�&�Y�i���θ�WT����6��!��0d)j�1t�<��%QD,f���@�nז��m��Bt�ѵ���n:f��#%w9��"��4m�Ǉ�Q��E���
��6>XB���ש��F�a>ˋu�G]uխ�y�GQ�Z��h�,��a��m��n o?
m�����4¥��(�BHM���1�<|��^��y�G�O
�`��j��v�v��up��.�;N��v&���~-�||yp,>k��Y�>nA�:�����AdG h�P��>�A��k$Q8x�5j4<�L\_@ �E�#�m��<Ԣ����jk8�vWӬ}��SJ�"�'G"���A�F���7c8-��}M�Z��'��Pn-P�q��q���-���"�DI%�%��o%$�y$�(�:�)F�\q��]�.Z��r�˗-W.[�$�I,I$�[���^I%�qǞa�q�����0�����#����"<ێ0� ��$�Ԓ^�%�DqCM4�"#�""#h���H�m���FX`�"#�,""6�2�:�GZu�!H�4�-""��ַ�Yu��"8�"4��y�Q�^Z�Z��Ե�"8�R"4��4�ȧ�y�u���a����"4�"0�����<<���cǉ#Mn�$V�J�����
$	,��+AG
�đ$UZIQ98�"���?�ZXx���T�&$�R�mD2j��i�h��Z�D$y*}v���r��rV)Ϭ�0��~a�j���li ��L�ORa)�N�/Ui��r�!P�d����M`u��ZA�t���s�S	}i����Z/'��c�b��#�B�DS{�%�:�uE�p��]�*�)�`��ޥ���&J�L�4[�,P�a�B��4Yf�d.�u�X�
��M?(��-/��x��E1~"R���.�o);L��m��0w��e�1�B)�:h!����%���We��q���p��zw�.Dg���!s>��pBA4�]�ϒ�� ����΢�}�&x�zhD8X<�ƨ��lᘄ�-���\�%;Y�3]�{[9�֫-.P��a�l]�;q��,���� ��a�^,���K!JPQAO��MFag�xü�y��AE@E"�l�؃��3D�k�.:,�q�h���s��$r��*�v�$�����=���ع]%=�s�n]a/���7�m�|8�ɶ��6m�-�tdU�m���P�\+�z�;=��:Ml�ݶ�a�4��k��z:M��lm=����|�vqǋ!a��'<�ҍ��@dc��Xi�n��������
��u���ץ�t �:Mµ۵H�3�rcD��ջ-�Yw3�8h�%0Đ&\H� �~/"��,�h,G����C�8��gw������w���s9�y�s���|�3���9��{�u��ekZ�u�]ukiy�Dy���6�,0�m�����C߮p!���0��\�=r^y�!���(l����r*Ko��Rn�p�������g��q̸T���3�ڸ�9����[����m�t�>{��4���/d3����e�t�P��C��xs���N��ۮ�z�h�v��K��
�Q5e�	�.��6۴����uтܻn�d���ۮӷ��ױ��{�~~Y^;&���0�ya!>BH!��h�i#Jt"̏%��d��r���w����w�U�'��U$1��,�'��	��}Ժ=<{�OP��-6dB��o�LY=��a��I�*��f�J�����!�xbf���F|R�ß}�bSA�%��#i������q�0G�Ty��Q��N����(�M2%�Yݧ���^+�Uf2�nb��rҞ��B��עs���C������΄���,6
6�( �J& S��Al3�:�R[urYL�S1Cֺ3Z|4nF3����g��<g\�tsz}xT�QzZ���um8��u�Qm#�":��"ֶF�e�m���1@�Cr"�D�6��芰aÆ�y�$�p~#�"�J�Kd>gN���B-���W��]U�X�<�g(�Y�A0��3����Տ|�;��ݹ,d���4Q����M��|��$�N�(��GL�[�msɝnq�N�D�v˾�xx�^-*3ck�u�R�l�3�m�2������nΌ1*��t�MR�m��xb��9�ц�&�Sal6�,���yku�]Z�G�DuE�l6�4�4�ܪ��_=Z��`�U��00�&k��{U�ѳv�?q�R��7��}���Je�2���Q��P�!kEW��i���Ȭ(����>�8�l��*!�8��1�#���v~�e	��4xl�j�T_u7�,��=nUFtgѦ=����Zx�4�|��<uGW��*0��JJ��D,���Й�i��b�E��n,}9UY������G]u�F��DG�k[�M0�M0�μ�Xh�m�����m�0�E�<Q �f�����A�(mQ�E�X�a��H%CEu=�EI&�JHFHC��`]%E�{��?g�1�s�Y�F�>|3avvm��a�v��TW�Q��:i��|oEZ,���3.I!��j�6y����&�ڇ!�u>-+]4D/3H�Y��	�k�aZ�՞&ۦ~��l����?m��)��U���Ue�4��}��������0�Z<뮺�4�<��"<�Z�mJi��,g�����E�ʍ�������@�@ECHSn܎�h�$Mp�!2�����~m�>��yy5ݵ$�aj�d,�v:�@m���{	�-&L�]�`�٧Cv;
�����q\5�.���U)�t��`�5	�o[�>�$�Y6�F˩'�4<c�ޝwi�k��!1j��Q1�a�m���	��֭�M]]����ʂ������gf�;^�22�.�"�?�h�Lڄ>+�s�V��i�E��gp�f������4��ߣ��\իj�3ᥭ7F��iԄ�KkcyyQ�gَ��[�f����<I��,�3��TT�#�m�uuW$r7	N�t\�D�0���"��KF��q�]�o�a_��4m�~�~yϯ��a�F�E����뮺��G�DuG孆Ԧ�i����{�V+x�l42�3�}��}��Y�cC/�T�:��j�8��m���s���U���k���P�1�)t!��lѮ�-�,��Ie�	���$q侀ʍ��QE�F�N�6o&]�r�]9=!u<��;%n�f:��8�cx�R�������{����B���R!�6�����-b)�紞��D!�W����f
ENZ�Z9ҏ8��-�\uז�<�8���,��1�B�,j��#�� �^hm�S6�DbR੤��m����a���4�Q�ڷ'�GJ���qxa��pg�TQ<>��Sr���a���G����F�Gs�i>T�&��r@X�GH0�E�+��ѐbTJ�,@ta���z��(q���{�e8T��0�Ŕ�d�c�����P�bef���R�)?6QDh����P �ᱯ����Nl�ڍ}���զ���uխq�V���#���"ֶR�a�ZS��l�սM��TO���ws��l��[�BHр�����ᅯ.� ���}�;v�QIԛ���N�Cv7;�q���vݵUQ��F��:0�F����y*1n�ʧ^{��WwF��՛[Xx�mY��oAg�A����q���XiPQ�F�1Y��:W������1��!�u���V`2��/4UT�8R�hҡ�;��}Κ�}�~��#��ӯ�θ먌��#���#���jSL4�Jl��gt\m7���A;
U+n���7&�p�pBJ/�)��k"f��=��ٰ� FI	M�(��R��c��m����Aֻ�p��g;�8�ٮo�����s=�7w\�N=��;G~�}-i!!��{Ē@"2)_��q�3���&����X�
�T�^u"��	*�v����FD3N䅻��9�(����^ml��ᭆ�ֆ��Rn�����.()(��|l�7�������d����:���ZgM2+-�q|E��2U���DZsy�gdZ>4�P����og�i����E��PZ>9��T��p��$�)WCd$��FZ ��D����"�`C�y�.�OD��ra��6�x��kҙy�u�]DeyDDy��ڔ�2қ穏P�6�p7����G6��x����C�$��GUc��Å@����A��6h�ܜ��ET�СqM>��iM�@���$���u����>�G
Kk����nb:h��(�GW�${������%��r"x�-5l�u$���
-�<5�7꽚4��;]m�2���[�NTm�-y3eZ����Lv�}�J�Gk��F~�2כ��X�	A[�����Qg���ӤS�"<���ڑE6���0��Q�Du�qH�"4����8���"4��$���.\�r��˗.\���K2[�%�%�rI[�nԖ$�InK�%ܽ�d���^Du�qJR�E""#RI{$��I%�$�����"#m""#jDDF�im�G�aR�"#0�Dy�q��0�4�jB"�GT�""�Z��-ju��u[�<�Σ�-m-k[+�rI,�bX��KR�Ծ��au��ZS$!�DiH�����گ�������c��R������s#��L��)����*��4�}t��{U$�94��Q �`r�Z�)��)�kY?��5˅4n���.4�rj̢6��=����!�<��L���o��*R?0>!��<α~�:﷭Q{��ޓ�T؂�|Ćx(�"t����B7�1�r�Xx=Q�B!����]���msZ�N4�Dz)�UBQ*��c��ޟU~���1�.���I'��]����9 7���s���9 7���x�������]u�V�Q��GN�:t��1�YE2�F�`��m�ps�p�C4�^H�2�wd��[��a�"��V�m0�U���l����6ތ\[?<|�a�d:|Bm3e�6��ۅUB����q�c�,�m�
�mC�Z���xN�������nʥm3��{ح�t��}Ih�� �H`׋��1��Q�K�Q������8�A�o�����.��{L�Dk�u��E�:뎿#���"""?-M�M��-+��u��m���څ#۝(c$%C�V�wm��c��sc� �}w$�o�z@@�~��&�	7���B0Ѣ��}5-��j�ڳ�G�*��a��@�+,�ڹuTV���p6��ѳ�|� ���e.��r��S�YN�����ѐ�o�ClyÅ��'G�F���Q�f6�Cix�f.����(���X>7�n_wʿN���6��sUkQ��a�Y&Zu���:뎢0�<�""""��0��,c���U��[�-��\�"�������5��<R�l��厔�n��EԉAڢZlL�g���j ��R	�ݠ��"s]�����a^���;�]vM�ܘ��m��ƭ
ګ�: ���KǃM�瑵C��H�n�hc#S�Q���^[Ǩ����	dƈ�lu��)��S����lb�
P`b#E$NM�:Mx�J�d
��c���,�£}^���m�N4��EL6qaE��DsI��.������:QG�-h��Ѧ=��7����&g�����Ɍj��w����g����*9�$���=�(g��n�,��Q���p�xD2G"qF�iC���%��hM�<6�g����Hw��>e����.t��Y���?6��u�Z0�<�"""#ǌ 3(��^Ε��P�XǛ�m�`p�E�h�����zK>S��7cуفK5����i���?����6ޖ�0�f��[ª���������*����>E��N�~s�%��i�n��c:q3��(L��X�����,l�v];��h䬹R�a��q�����K�	ݤp�0��}�~���t�)lh�u{|$f\p^�UU	�Q�[�}U6m�^m�^G]qխ�y�q��)��e�;�~Ϫ)R�Q��l+��t6�ugOYf��E�������1���a��_�(�C��'4Pt�ǰ�`�2��\�Ì�u��l�r�uR��1�"*%��he	���1`�n��+(��a�g����6�Შ�����r�Q��Z�|�l����TY>J��2�_o�H��صS^��9�41kMغyQȧNy$�����۰��cvb�͗�ފ<��?"�u�V�#�#��"!�Ǎ��Qc+���ag�P��N��C$en�m��ߪUr�u�ϫ�Xb���ם~O��v�s�D�F����cf/ЊbqW%I��N&ۑ�����h�d��'7���_7�ƬѲ��|���H3f��x�A(��x�k�N`���&�p�������B��s.IP��^�a�����Ƴ�U��X�
p>Q��j��j���_��Z���(���!�1�ClÆ��M�<xۮ����<�8��""��(��  �{�I�%-����1��DJC�G���iF�"Ȉ�l�&���@o��>]��F����#������v�E�'`ڌ� u���B/OqoYS���\[M���T�+�c�����$����}�V����Hd-��Q�aˀ���������(p�ѹ��홌�w��ܕL0"gguǗ��u���&)�U�,��g�S~P<5t<����e����ݔ�U1�,���)Du�gf(��VknHJ[���)ӻnI����=j�*1������`h��/Rf�h��S~6�������9�=��Q��Z~/Ϳ�����!�<3zX���I�󰌯�H��Dh�ʁ�c<�������AY����ѣ ���C������/��Y[��,�ޜ%J;��8�~�N#ȵ�뎢�G�GDDZ�`��e�����g����p#!d��l=eh���9�v�G+dXQ���HݑCg-���g� t��a�:�9�&b���/S��Z�Y���ȶ��QI�g0���3�>[Z�yp���6��F��|aTx�8l��3�
��Bۧ*S��eX��F�6��j����p7���-H��%)	Xh�G�Y���G#s��Pq3��cq��X6�#�>b�_�K��Q��Ϗ��:�ayDykq��ݝ:vN�EU��QJ-)����d��Rm����i���ԗ�<5�fHIfs����ǜÚ41���Ǒ�.4��t��^Ԓ0`i��VG9e�i����Fx�F6m�wM��#E5�m�òd��e�wyAL˘��ƭ���
��nU2�+�V�	C�o�����/(�8Pg=�O��9!�7���"Ȍ�ճ�ѷ�� -���٥�GKT�z��΄|�A�������g�E�s�@pm�/,�<G��q�n����#�#��""?-�
m�YiO}�7�Qө�d��SR��Zm��"7i�޷�GM�5g���h�E��VQ������L�ҕwN�]U�%�HS�*E���߁́�E/R_|O(�x�(�Ș_X����G���GN���:!��(d>Z,W��8Wxq|������sM��u�7���H���ru�)��"��h��tQFϾ\4(V�������f�����o�1~R�Yac4�pt}kM���8�O����ҖW�UUUf�l͇V������sӳ�"����v����,l�ݦȝ۽�}�u�ӷ�[�����Kl!翮�;"",DE���-�-�E�"-�"�M�p�����DDB-�"�"&�kmdDM"E�Mm��mDE�4Y���"�"&�h�-�h�����4MDD�"mm��h��!�4[[hE�DB-�"�!��"�B-D��X�m�di,��"-���""h�mDE���!�"""hM�""-�4[Bh���D"Ț"$[D""��M�d[DDD��"""�&��h����DH�"&��4Ym���DȈ�������DM,D��BC�3�DP���&�kmh����DE�mm�&��"h����	�E�YE��Ț"$[E�B-�h�mb""-�dD[D��E�DX�4X���-��D[D�m"kmdDYDE�4[D��h�&�"�"-�""θ:�:h����h�&��"-���"-�""Ȉ���[D�dDMD�mm�,DE�����-�DH��im"D�mf�$Ki�4��d��D��M"�d�m"X�I���ki$K$K$I���$��$KH�Ki9fsim"D�D�[H��4�D�d�4���qk$I��%��Y��I��H�I���4Ki4�m"Id�h�H�&I"D�E�%��ĉ4��,�M"X�"BD�d�4K$��4�M"[Y�D��"[I��d�pultK$�%��K$�Ii"�%�%��,�KMXZ$�Id��-��E���,�Ii�K$I��5�4��Ki4�"[Y�-��m&�,HKi5��4�m&��i	m&�[H�Ki4�&�I���Y�i	2M-��Kimf�m"B[$��	m"�	m"[I���M,HY�&�-�K$�$�Y�&��,�-���$"�%�i,�$�Y$Yf�i%��B��4��H�E��[Y�I%�i4�d�[�%�HI-"�ZH�-$ZK5�ȴIi$KY��H��KI��$�Y"ZM-"ZD��5�%�K&��KI$�։m�$�ZM,�K$�BZM,�I-&�Z�	i%��M"[H��g�$�$��4��4�D��$��Y"�m-�K$K$K$Kk4�,�,�-�KH�X�,�"[H�H�Y��Ki%��%��Y�����D��"Yf�d�id�d�d�5��ZH��f�D��D��Ki�f�4��,H�-���3kg��sd6�[f�Lkdm��m��ƶF��u�.�qs%���cX��l��m��lke�kdͭ��-�ml�Ɔ�4-�m���6Иж�-���,�[:Z�M�� ����b�ZBB��HY	BAd�HZB��D-6�BBА[AhI��i��k#I��Bi����&���!߮����К�D�5����i���I���Zi5�YFz�&�Z5�H֚#,��4�d�i�-4�Y5��kMM5�Mi�4Mi���Bi5�De�D�Md�Mdi�5��5��4Mm4Mbh��i�X�&�i��h�#-����&��ɭ�����:�uÈȚɢki�kMX�&��M	��&��i�k&��FD�ki�k&�h��h��Ț��5�M4Mm4�&�2M	�����&�i��h��i�D�M&�kDe�M5�M5�Ŵ�&�2&���D�&����h��dM4�&����h���4і�M5�DК�kD�&�v�éF[M4�5��4Mbi��[FM4Mi�i��Y5���#&���Mm4&������B2&��&�4M4�&�ki�2&�4�[MM5��5�h��k&��M4�Ml�i�����hMm4�BhM4�M4dMm4M4֚i�i5�M4��4Y���m&,�4M""�&�dDMc��b�"&�"h�DDE�Dő"�-�DE�4Y14Z$M,���&,��DDE�!d�D�D��"DE��E�M-�[k"h��!F�Ym���DH�$H�Kmh�"Ȑ�"شH�H�d$Z7�]���-		�!km�dDZ,�m�kDE�B�l�h�-%��5���[i,��	�E�[BE�"��hH[B�H��Z�	DE��B�"Ȑ�$Y�gZ$B5�Ő�Z&�"h�Mm���Ț"-�dM�[D�"E�"E�-�D�D�DBh�Ő�hHY�M�E�4DZ!����4Z$M�dKmۙ�"h�&��[kD���&�"h���hufq�DȈ�"-�"E�������"$X�m���Ȉ�$[E�"��M,�E�DYE��"�H��&�"h�"�L�""Ȉ����ֈ��DE�D[D�e��dH�$,����D[D���",�Y�dE��-�h�E�MDǾ�����q����������3Ì���o�������fkM�%����͗��>o��z������>�����o����;������������o���]{�]~mt���8�>�o��q���|�vx|�7�|�uؾM�>;}��gg��?�����g|�9�?����������������������?�>6�������nE�kp��K>f�k����>﹏����ߵ�l���3��-������~O��'���>�������6����^?��ʏg���n��x�g��aؿ�ovk�gߞv���g3��9��v���n}�<y��<��}��?^}o�z���߭��i��&��?���|��u��lٛo��c��k1��Cp��@�i�7�Y����6�!��1������8q��?.z�ι�������|������7v�=ٰr�(HP���盌35	�e	3l���~���}�f��[{oO>��o������}��O�����C���?�����׉���~���2i�3a����]m��Տ�����������Oͽ#�>o����oGl|wsٛ��~o�O�^�~�vo��ȟF�G����o��}�-��_����3a��K}�}������s���~G��������>f�,6͇e��8ٛ����~��o���?��c�>/���n����s��'��8��o��f�w۟]IK�ӛ��[��m�l9�h��^Su��ߟ������5����m�x����5�}���S���o��|�g�oL�����sc���z�}���ٯ��<}�fl>��w�X����ϧvl�Oo��f>�����||��/g�~��u��6z�O��_{~���g�ݿ/��k���ɳ�q?/7���o�7���;lٛ��|�����m���ߏ�6f�ɾ���}?g�?������F|Ϝ�F�&v�7��ߧ��O�޲�y�-����7wq�w��n�|��n��G��dߗ�{��0{�z폟ۻ:~>3��nۮ���{{�Ǉ��6=����/��s���g������t�[�<�Kz7��|=oY�׬��tS�|;7}�������՞�>o�}3� ��~��0����~��������o9�����`��v۞��_�������7�3�}ۿ�������g8�Yl��g�����ܑN$<�[ 