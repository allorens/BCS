BZh91AY&SYF8��ۺ߀`q���#� ����bE��@        >�ᵒ�����6�f��SjXe��bɫfEa%	�D����[3Hm�cj�2ٚ2j�klȴ���`���j6ML���֕35m�����a6���R�ͫ)�3bQ��֫)6*�Z��e[2�Q̒�"�ѴѶF���V�VͶh�5JJ�e-�(Ģ�3, G6��h�6�f�z ��l�3Z�ln<���YT[[e6�*̭a��B"�k-�F��Ҷښѳ%��Qk6��T�ɰ�b�[kcY��0�����R��lZl<  gu��-��1mWc��Ժ[K�4wuډQN�ݎ��i�P��v)E�`鮔���'M�v�:�2�Y��cM`���m�Eo  g�A� 3]p4
�`��
 
���@( #6� J�껀��  wN �R�N��  �/wB@ ��Ř�ɲ�k�ZMc��� ;� �;�  1��  .�pt����
C�ݞ� ��>� >���
�҉�>��s��  ��MYe���Z�Y���l6�  �� t�ӻ�{�  sc� ���x t��Y��4�9�p2 ��sm�נ�u7@��v�����5�J4��MSkii�S4�cm�V�   �;� z]�C� v�\�ݝ5M�[��i��s��: 7�ۀ]t`B����@ ]\v�@��p � ��m&e�+[Zj,�i��   ���  ��� �y�� s��  vrq�t:,���� +�ӝ���T�	�8( �D�8P �\UL�i�6�f�fʒ[,   o �C0@  �( uox�U�S �Ƙ t�l� �����q�A�ҴUV���[Mj
���   ���1�  f��h��NP��� Wp ���D��
(P�j�� X� :9Ի3j��Z��5V*YX��  �����w  6�h ��:A̹� u�� �� 6u� �s\
(u�mp ���S[Z��ɣI
��m� ׀�s�����t
�� F�  �@uW4��.:�77�iZ��π     @�
O@RU(d � A�"��Ĕ��ɍM0 �L�#LE?&!)UM d� M  �))J�4� L�� �db0��i�TȦ�)�zdOI�zG�1�OMA	H�z����l��M  ��M���N}(t��3���5���`W:�i�+&�1l��ϗ}��ETW�<���� *�
����� ��χ����������%g����u2��DUEh�iJR����
�+�`��B��Q?��o��G��S��&e3	�I�S0���e3	�L�f2��̙�a3)�L�f2���&e3	�2	��f29�̦e3)��f&09�̦e3)�L��0�#�L��09��as#�s�fS2��̎e3#���Bc29�̦e3)�L�fS2���Le3)�L�f29�̦d�s�L�fS0�9�̎`sL�e3�L��0��3d&2���`s���0L���.es	���G0�fS2���a3	��f0���0��̦e3)�L�f2���e3e�L�fS0���&a3)�L�f4�f0��̦a3	�L�fS2�as	�L��2���&a3,�a3	�L�f09�̦e3!�`3)�L�f2���&e�̆a3�a3	��fC0���&a3	�I�!�L�f09�̎e3	��f�L�`s#�L�f0��̦i�̎`s+�L�f2��̓.e3�\��09��a�s�\�� ́�\��s29�̎`s�\��f29�̮es#��͙L��S0���ds+�I���W0���`s#��)��fG2��̦ds�&G09�̦e33�L���2���&`s#���G2�e3)�L�f09�̦e33��f0���.ds&`&@̎as#�2$�#�DsdÄ9�2���.aQ̀d@3
�d̨��2����P3*̪��0���#�s.d�(��0��T�� s dQ� 9�0����Ps`��I�2�fD��3"e� 9�G2 �EL��s(�"&aE�*9�2�ȋ�As*�`E̠9��s�aA�"9�0*�U\ʋ�s"�eQ�(�"fʋ�@ʋ���G29��`&L��S29�3 f2ds�̤��0���ds#���2��d3���2���as)6as�L��S09��e3L�`s)�	���S2���e3�L��L�09��`s)��fS2��̆fds	��fL�?�M?���7�=��v����\�'������x�\���j=�Pn|M(�G�ɺ	��Ɔ���
�"q��R�EN��Bn�i�q�#.W�ML�]-}څeǘM5�@j�`�nj�ţ0d����DI`\��/���ͼ�IT�s�O �允�e�m�t�Ȕ���IA�w���Ė\��9�)'�����Tq#��鵙KE"�E+�S-R���{�H�I��,�T�M�T�L �n�d��;�V���V��%�9�넜���s\� Щf�sh�]46�8Hǚ·eA[B�BL���B��{�
�4/�&4Iۻ��4��T*A�D��u+�&R���)&����3cB�`�J��Y661y(�D�K��ʅ�9b�le�2 &8RK�K�4�J�낥h��"{@�:�)d��Ū��8X���zU��T5Dsl1�q-�A��z�6h�7Xi�H�rV�ˣ,TX�!5@�\1Z T���ĝ�iʀP�r�97�b�@jF�������$Y+F�ݸ��t丂�5�,h(�1� �0]ALͽ���;,�%<�y*酚b�-�P'�%E o����i�:��p]�,I��Ԟ�M�S�ǰf�pn�go%����SU�7.K��ᩔcu)^[�2����2��-?\����im9��H2��������Yc-��SX�©��#4˒�)�
����+{whғJ���$�e��A�����LҫI��Pم�b��q�4]]�(��ر��Z�EY<��K1P{�+&M[���(ș�z����#n�0�,'?l��36ے8�]E@���r���͙���m2fSp�x��eE���lyfk@���bp1Q2
��c.F�>��U��
�
�YǕ��sZ�3a%]5��2��ҡIVh��=��c���m�
�;����em)W���i9&;�ҵp9��a��\���o��c��i�`F �/�R����BM,�-�Y2頻i�ue��2nAW�ƹ3@3Y���sM�%d$��m ��6XX,E�Tx����W4���o3����a1�T���9�e=@��VsB�4ѫ�8�Zn�ʴ��&:{iا��ql�"(ݫ�)3&�&��R{5Xy,��N�2Z�ERd��i�U<�n�4�YR�0���p+W�nDT�
$	Q!.�k-���l��7R���	�oB֎\:�VV�	�����7��L��bQPQ��n]+/�^R�T����z�wZ��^@�K*�`�K��I}�z^"�"D�r;a]�p��-ww��I 5=Lb���mJf�lYʱ.��"&��F�ǔf���Q&a�gqM�[n5���h	����[[��-����`딎�M�ķM6��eN�[u���/(ZW*&ۙz�#d��@��׊��O"���*᭩���׆`^�4E��"k.��@�Ӻ
����=aˬ¶��,�j��]c�����&̩�	�X�i����1�"��a� r�@��n��7`6tR�6�Ҍ|�a�#E�/.uMJbj��\��G�3PA�3v���m]���dBL��ą:���:S��iӜ������ݹJ�*5��ؒ̈́���n&�il�{!�|��#��ۀT�[�e�R�#D#8���)RqR%��$si)u��h1�uzS�3*h��ѱ�-bS7CO�͏sy�V�e�A��rՋ,ͣ[N�������EY5�ۦݬ0���ݰ��j8%m��*|�n �`.�ʛJ��KH.�ԥq��u�7��ޖir�����#3Rܙ�3D`DK��V��ej��)͵7�^Y�4�{�52�v��O[zKzr������ifd�*�6����cN�qӲ"�f-d���8��+&��$���M�Nƴq��ʨ3 ݺ�- �v�ķ��&	�%]�Z�#�"��Y�֠��5����Ye�ekIܒܣ�������.�;yBI[�]*4�U6&�2��N@C��.�'vVk�f�)�T�qڣ39Xi!G��؛*ܼs�2R`��]���d�|�p��"�81�ân8uJׯ��֖��͵Z�e�ZsJD��.�����"4Ր��HӢ0Q�[�Bz�̏j��H��D�f��sp������tk�i�٪�B4.����'�9,ٛO
�΄ 8�	�tq�hzijp9��02�P���iS0է�f8�r��F�<LD,;˃PJ���%�*���e��V�Kb�أ��4�Y�nh[
r�i7��ӊn���3L�``9]fml%(썁�c060|��Y�,M�U��  Xd�{�
�ڨΘ�2&!���cE,h���-��,�&�#Q"�sM�Vt�d��٣d�5�_mnc��\_O���8�f��""@&(H/U�2�����B�&���Wu�ƪK�K�&���1�t�]
W�)�N#�A���i���%*��Cw+% �"���MCq_�n��`$�d�X��� =�Sń��[ǋI���E嬶�h�2"ݛE��h�J�&�Z�L���1�&�*���aN��`ZF㵨Eiz���9�SfSw�֩[�H�)	L=�	Y�l�SQD�r���f���4h	���Bw3BVm�*m*��S^��h�5 VbtI��(�C.���Iwr&i����3�,Ȕ�^�0]-Q�����A���L���Ct�e�-�������]C@��k��6݆T�"J��z,��,T�o 	:n4Y&:�)b�B�埖zK�˨�y�Y��Yk�F���aߖ-n����z΅���<"K�tܧ[̼���s4	@�Y�>�^'S^:qŢ�o�3q�0���#���t�]���T��LR�R��{�I�R*���
��D�U��ca]�s)�Y��K=�<fBi�����a�F��Jw�Z7�GM'�f,e��h����p ���i��������56P���t]Iq;��,�[Qx1�K*Q:���٪:�r�m�d�e�G&���`��^ێ-�l!Q0;�YE���mk�j�Tv��;U���2(i(*hǬ� �J(��*�#`��E��i��ֳ�ZU��F��P,�,��g4⛪Sɹ1�۠�7��6���wh�5n�J��1�e��p�.=ܡ����M:�E�1k/k$v�Vi<DR�k 4�(\��֋���n�1o���l�X&����H$�"�V��7Fأ�\�@��0�K]��K��$ҩv��f7(*m÷
-`��)��٬b�����Ѥ�ږ�T�ti^l�z�㣨�Y��Q�Y*�j�YІ�ooh9B����t�oM�B�]�L���6�I�X���C�[;b��tnE�'��gD�u��V���k����C=��d�B�u�Ԑ�����)��7`VK�J�b��Q�ͣ>�m��	֛�@���U�N�J�"p��&9��3@Y[
�6��`�OnTMKh���g�/q��A�U�5�v����o^�WX!b-bX�&PE�͵O�I�1lc˸cX�*t�O�T,�������Cm@��kr�ehޙ�R���#=)�ɣ��������Z�Fh�`B�U�>{�kZ�WI�3�I�R��k���ʰ�oJ�iY)XK�m7+Y�
�a�Mo3
��j`rF��u��t`Ǯd�]�4�n�&L�
�D�
n��c��[�u���~o���f���&:�4Z�X�Y���R��舱X�hR�jg���Gf��8ȓ\�
-�q�I�Պ-̂��-i��DV��*8Ѣi�¨�4�B��a�4p��˂k�$�4�+u�F�j� �K Fm�nbYQ�Ƌ�M�^��
P=a*t���6Ƭ�Ƶ��n,R�R��("�f`�m�Cduq�/T³q�"��"��.�1l��N���(��5�f`Ƿ�{N�يleU���� J)jZ�Ml]��X*�V�I�0�0���\�p�����E:7�%H��c˭�7t�]��e酝q��m��P��������dAb��b�x9�:/n�2�L�8�A|+L�;7�8��יq�X�� �a���+�����L��D1�or�P�M9�`Z�4���Q���%h��� ��3b���Q�+v��^�lHދRMvV�n�4r%�1J;CA.e��Y�~�ki'��7��x�͏�@���A��hѬ8�'4c*�k$�Y1�I&A&�ֲ�E��@��j	���x�e��^�'��gY�1�ט�*e4i��B��fw0�YkhmY+����imk�")f��X$�ƨ�zk4kʴi*r�m�a�/orR�����j��k431�
��5F�(ډ�L�э+k0Ƙ:��v�1��6����a�g];T��N��V�flʁnӕl^�`Tke:Jݳ�f�N:���@�z�T۲�YEY�b�e^�nH��QǙ��-�6LjàTUclJ�4GP "l�����V�,�{x���R��ER`%�oi�Q`�=�n$�Zh7��VH�-���fGN����d��t�B��ڎe�e�A�2���%�L�t�/V����W��j��k��^����f%���@#7u�ͦ�<p|Ƒ��u+&j�&j����5KV0�Cj욎b�#�����ՙnT�7<Z��&^��BI�z�����ʱ$��z� ˁ9�)h���0c)f�kq�+�*ͭy�q�*<(��aR{X�u�fYCx��҈�yCp��Y��������m�!r�ݘM�z��EdM[vD�s,�=F԰�Z+nmJRiIJ۫.�OR�L�g��r�42�I��M[�x�w5��뽍MUSs+.�:TYz�4�30�!7��Y�:��\ϯ7-aʆG��D��=gN����$*揮j�ǋ�YN9�n��mn��:��u�2� �m�Bi�|��FV'4v&
��ݨ��`ظv}�n8��Q@�oj�&�z�ݠ���2��v����Wr�v�k*���ɀ�"&���2�j
1�4]mi�{����r�Ƴl�˰Ti�Ԧ�7��#��Un���t�3:��Lz�W�e���+����d1-ɔm�B�0c��%2��֩U���u�X(�qjWy2M��+`Ŕ6=���Cz3^��V��]����V��=�
n�3�j�Æy��h3�i��Ju���{s6�1"��D
Pc܄,N���p��O� ��n�+uc��h�4 ���f�͓UǤ�
�ىF�ě#I�5z�5):�g]K"z�Yx�E��[g0kE�:���w*I��䷃e �Bb'�V&q�v�@�ǘeE%R��/P�.<s	�[�椰)����8ud�#���
W�����^�*��Et׋h��V�l��w�U� 7M۩#X"%�9��jA�y���a���2Bq�(ܒ9�����t�nDij�f9)Sp�tIA�D���2�Ҭ��8�B)�,R�9���G��IW���c�f�����ݡssh�"����)H��7���찝3%鎐����n�[�'FlBi4��`N�؂�+jLkPx���ܬ�y�cU��Bp �"�m�)v��g2\��&�L��T5��NV��q�Y�QJ�MmжZ�=Фm8f]lA]�5��n	��Ɂ`�X	x�G3f]�A�X���@;ji �y��Y����ˑ��m�i5�lĨ�޴�	������e�{�L\ �g�{����f��թփH���F7Q�6^���z��kn�Z6]D��[���D�E�׵�r��H�U��*B�qG6�M��ƲլQ+�lL�ʖ䬥��ڽ���7	sSNkF�Ia�aH�Щm�%y�ZMAd�[5�0h���yx��������"Q��K�
ŔШ�ˎ���L�XƳ�i��t6�5*)f�P(Hהݨ�4Rq[����4kL�V�G.䣒�clLl#�x�� ^�E3Me��$���u��A�2���34FhM��F���4,�d�%�T{Q"�&�������lyZ� ���9����[&V=M�����lx���:^�lǶ�UOOۖ ���
Z��!,�e�2ɏe�X"<,��V7�-�L �;1Q͏i��,j�0ը���V6�e����������^*[�ȡx�|��lwY�פ�y +C�e9 lӲI�3*�^J�ע�-JIB���f�zD0����!WZ+I�k�����ҿ�s8��,�y���e=HvBp�"z"�ԧ� ����V�Tz���`����1�L�ˣ�썽�Ǧޭ��y�����
�jq��gۦ�v3�K\9�\��\&��sz��u��4ӌ^��/V+Յ�
�����!�ʐ�0�%���'��9#��(�鍷e�dʸE]��@�`tVP4l�����sMcH�q&����u��x�b��[�j]�锫l������5� ׻��<�����)��5sw4�pflp
�"�����#���GEA2XZ^��X]�\%mt��)�y���7a7^$E���eȈ�zx9���Z&�G�~�y6�{�oW.u�Vf*9u�hv�P��p[1:帜�.8��u��@Y�Xoh��W����T�k�"h��{Bķ{<��հ�6r�4����%m�W��b\1Ro9.6�0^�v������r�ҹ�"�>I�T/&�E&�B��(����UOdR^���mf{)���/1iH��m�:�Q�(Y:H�c/^B��od%�ԩhH����ֱgDq�N �]�EaG�\�C��V��Z��Zz�C�2���+e����i�	���/21�Ξ���X3K�yF��nJ��E��f��*g�8�Ѵ�#�<@3�١�?�E��g�����^�����B���m�_\m��I$�I$�wwwwwoo9�ܙof�P(�Ćٹ��]ud�y��jݒ��w�U_m0�?�+�* �FSW\�����շ#�]�K��%��� X�t�udv-U�.K+y��C��ȯ��g����$�觋r�^!�wk�1ƌg �nv��w:� Ei�dʘ]�M�Ǹ�����g�S0r��Lp)��X������ ��VT�w�i�}��<��e�Jul�nf[�Q��������X�a�\��E�z�(0�Sv����ڤ�f�ko;�	aW,F�o���
5��p��ol:�4�+�t�-Z�:���J�o%�$ҡ�Q;���V�"k�%�Gy�j�[��\�j�s+�m����#z��&�*�XeN�$WZ�u�E����f'�5޾Z_R�in)�8�+���7Hٺ��#�i8P5���̵�P��pn��v�88+k4�JG�d��D���֙Ƹ�����bT�zf�2�%m;�1�N��+���$v��}`]��:��:�7��c�X��-b�C+��h�)��1uI�\/�N�+�;�7�us���WB��)�̡�F���ns�:+Z�$���/��t�������N�(iP�	Cr�X���py�HfI��~�#�#��+�j�%�W;(R^�Ɋ�P��ĭ�|-NV9��K� ��+�Yx��{5���'5NН�̈V���Ķ,3 fN��tV�y	`1[�.���v�4;�Hr�<��#{���[T����:q�y��C:h���sE��Yd�d"�T�8UcDv�NN�z�����uX�P�9��򃀙�.v:}t�`�T�U�,V�0�7�����k�.{�'p����#�������$�/�S���d��KF�V��fv#Y�mZ+:��-�$,�(���,DR��v�;1ю��}��6�<@d#�  ��:Jfh�#>�Z�}�@�FM�0%�:����X �\��@�(}%0��Ȧ>���6Xx]\i.d�i6���n��=Ӭ'8w6m��
��4�� �6�S��ͬ�e"�hq��
+T�E/�a��M8�޾�x4u���N&
;^	���S��'J�W��ws��|���Vږ�9�3/VjAl�,dn��x���m�R�!|��"D��_,�>�.���9K�������qt�A�7�B��'Jǋ�s4oQ�PFr;��n�>��8Y1�Q��wv�_ƺ������n}k.��l�x��^ܤ:��G�r��B���ʾZ�"�."��.�|�Zrly[@��Ι��8e��:���ֈ�	�����h��I8Tw�Ei��su��!�NE���h���s����$��{���U���d�4+�q{ۗ�8��V[7�P�`D��/�̾UNb��ҚiJ�:��������(�%f��c��^�|oR��X�2R� ��$�4��6wgx��Z��`�!�=��[Q���AM-��^�K���i�0�^q9Y�i9eg7�s�����n�Nʅ^�Q��)��4t���-�cRf,ۮ8�ʜܚ���yAJ�v��ĵ�"$N�9����˓'��3�Ttc"5���C�T��6�f��u;
����ghPCWZ��!b��fU����d9Ӏ=�O^�z�I�������K�b�*���R[S
8/���;߅cum��Eg�ޱ����a��My� y��lq]�����HVfт�Sy�U1:J��&�<��lE�ϙg�a�z�&<�ś�/4'Cr���L��t�1����i����-�}������{��ܹ�XGm�5x���@+�Q�"�S2�O�����k^�Vq���>�,᝭�59�?t�ɸV!�<;Z�j��s;j��ho��VU��Β�sHH�j�:J��/,�hI�㍨V�����32-��J��ܙ|�Ύ���1��/B2�(��@��ǲ��w�]Ů��oe��f]�Ҁ��Q���:+��).uMi6u���u�D� �C��e�1t�ޒ;[ˉ��[���Ny���6�]����>ȎC[o9}���i,�ý1�)T�4��*+6#[��ҧ=:�����c�D�-�u������i�W=�4r����8MJ�
bC�wݠ��+T����.�Z�{o("z��<��7aGƥNUʻ3
�ee3A��7��
p�@��:���VE�&�̮/�p}�	��}���WD+��ܐ�׆��cf�ƦpLys��־�T���\Q��i���e�ױN�)��MQCi*�Vi	[�u�D{�;̇�N�W�������^��o(_�����9p��a��1�o*+w/)��3�Z�VUs6wص��@E�=���MRǽ'5��U�q�r<8�;0q��"��2��DNX����r�>�>�+���Kj�'x�q�wάWY&�S����Y���k;� 9�V���Fҧ���a��;�DMc��������j2�N����o�VO
��V��z)��Ң�Q�_oF�n��8��y
*��ؾ�]V���qL��mo��K��֊��R=w� W� �K�q�����[��H�5���raA���������D�Z^���o�ۂ��Z; �Ѭ:���uz����[C �������S\-�|��>՝�Tۚ�*��K�z��盻���p��X�Eo@	ұLgj�7�t����eϳ�9��QOw'B{��()*Y[��2Sz���"q��^R�8طР���w{��!n�1�U�ȶf|yp}�l�l��C��x���2��D�nh��_
;�l����od�k���onC��&l�w�@�=i%��֏�2��
�@��.�v�iܸ/�m^�&�x蝎SF�Q�"ǜ�I`5�h���J��գ�9��-o��\`���=�h�\77bP��*��,�{�1�ou�����GW����r���bF�E �A�#�웅�����mi�3o72��]\r��ꜚ��g��ى:��!��#P��oC].<�*�E�Jr�]�6*�o�޽�P��j�۔$쭥B��;w����b�n�r���ﳣ����By'�[/��b���khR�t�{����T�r3��쐁�T�R��WKE9+��
KYB�`!7B��+XgV�ށ���tŶ�ʍ�!��8��y6�[u36f7rJ䖍�`��C}��gh�٥�}�����{��q�AW�{.�v�@p�}��c$.��6�|P*�{F�t&��>�iv��M[�о�Vy)ێ��ô���X���jT��5ח�CV�ݥu���ǝ�!����;J.����f�V����S'uY�Qȴ��r��dG�� ���E�C�ׂ��� #�4ĺ�)��P�7;��:}V����.�<4�(ӫiOAC��tm>��U�D�Boʘ��:��r�\���j�X�h!�n-v�gu%�25���.� ��qp5�T/Z]�n��p��
�r�7�l�%0�f6��G�#�4�Vo���2V�v��9�;؃z;%%���2�ns�D��oPd�	�u[:��-*�v�8�wk1m���#�o ��=��^�Cp���-I�X�����X���ỹO&`�[��!I��Ss��(�u������D�S^;�b�β�Yy���L_䘩�7��B�L��ZKr��wݴmQՃ(�$�p=w܍.�̅H��df�+���g�Ꝺu1.r�9;��d[8�R�)��P���!�G.��2���.]��j���9��nE��+��уͱ�;V����������l��o{�*�Ŧi�v��#�L��]^f'+F��l�ݛ��Π�$Ԏnѕ���=חP�;��)4��h����8���q�rQ3/#���ʻ��sh��Z�S/���g�y���qR��в'b\�M���.�=7��F�S�E];��6�)m]�9��W5:�i#;y�m�TEY7�!�:Wo �M����#��
��^t������
�^�5|�ܓ�C�n�y�\���ս]�4��(Ε���O3^W4m]���Tw�]>Wx-�*EP{ڀ�0��qWh	�e��J�{|Z��Áͣ�ئI�Yi*��DEu�� MBѥ�m��l�0��_s��:U�)e�i�*�{0k����N�N6tTG;�5��gT�{���ݺ��\e�s#�7p�o��`$���j<�otw�k-Nw��M�]�X������V���*�.LE
v������ͫ�C�j^>�a]6��W6�.7�R��8apoa�mS�m5>�Q�:�b�9V�	�KQ�Z�ϳL:��e �q`�v��}�-��<e��L�«��@õfG��ٸŏ)����H0�t`���g��1�C9'��t`���ˎP�#u�:�e��=6m����+���g>ܚ6˚��|��l-8�}�t�;�lF�]�����`���Z��28��v*�A�wR��D�:g�����^鞚�|j�!��o�`��6Y���K��.�'%nQ���Ax�X�c�i���c�P�k��/�LY#0V��<:O��B7�%{*uJY��u3���ӹ/{
ǀk�@�{�hEszn;kS�F8��\Ѹ��s�N��hA�
۩ӆeG\��)e�_%t/vJ���2��V�L��讳w)W!���]��#�=wt���TC�Z���ms	qN���q�}@լ�J��k�7;�N��:����a�ܮ�R���*��ɹ�:�H���V�F��ȵ�aێR���L�ڢ�b�κ�t'TB�'�7��|׼��tr�8om�=̐]�A�L�.5��#����q۪�fb��;��[P!�)����(��r/v��\ws4+�4ѩ���h(��,��v�ONG���U�ׇ�5lv��-�����INܬ$Qw�T���.�$8�z`�����B!���,]��}ַHUo�A�2r]1�^��������dD�Y�{EL! Nyb�-�N8ʫ�ҹ0�2�j�r)�707�M�{���h�V���h.���0���Vw�ʃPn[R��G,>m�ow1�_r@�\5�p�t��ì�?����]�ћ&q�fm��j�P'��/�cw2�Z4E�=�i��.x�D���v�v;ܨ��h�x�!�)���c_&�lS۾�W*��$�5�-:��"�b�<���V�(����H�XJ]�9n�nn)!:;*��y[���0D����+����ۊ~>ӕӄ��RՈ	���46<��gS��ƕ���@L):�(��	y�X��=��;�btGZRJ]j�x=][�w0�J���ӂ�ܙ-���2��ڿ�x���H-u�����*-"Y�c��y�͗���6�$&λ�p�D�?��-������3D�=�f�G�w;�Kmu��y�=����J=L$�ܕk�*�v�S��̝y���[���\-�X�i��l��ToN@"�G]��y�,�$.���dT�v҉s��{0�͂����{\��O���Փ/X���ޫ��=��D��K��N's<+5��!������z����$�l4��w����bC��m_N�t&��q� �yqu�K���٦�n�� 5�Y�+�y67g9���l�L!�.������mא�޺u��av��ag�m����(+���`��r)�/�5�eess�åΎ�Ę��nc�$34yV��{�Efk�:*�������]��X'S�=lǰ5;;�o��DT����7v�5��ɻ�[�c��8�hb�v��zm�yl�Z�m�
��j�4�qvӃN�;sI�}��Z�z�8��
�Ι�leí��*��,ym��*Ej�>󕅘k���zᬷF�ٴ1Q�Q�-���W`����h�,�]�Mup%P<��|�I2��D���9y	Y��VF�n�
uh'3C�G�օ��7P�I,�����f��K�Z�P��1o����n��f��6�2T��tY��Ck�����J꾩K]%%޾��V�)J�ٍ����dHâ�H�.�9�	�ӝ���7�� 
٥敷�Oeu�Ƀ�{�������΃E�p��Q!��1��g����n�I�	��D��jM9�s��ݞ����º�]^Rh�uQ�W[0�zi:�G�kv�t�W#��Cdcjv+��Lgo�S ���b鼂��N�]7U����-v�[���:�P����}w�|tw\vd�����OzJ(M���ʛa>�$�sww��h� �d�Hت�UE� 5Q�b)��
}(��T�%���H,�m7�ܢӧV�`4��T�~,�%[�Y�K��t�l����M�:��T���$?K��L2����en�B�L�$u��0%\-�K1�v��
t��SeP4g8�R�H��7�
un]<*�or���A'�8h�(�o2�Pv,0B'B�U(�&���E3B�]2h( ��ŵPMDPUh�$�V5F~�`4@���$�dPL�PL�`*4@���R	G!���N@��5�D�*�Q6�Eр()B�g;s%e%�Ptx�R�{ b
�NӤ�AQ�i:`ւeTlT_8���(����4}�h:G�
DD�?W��0|%��OJb
1����-�&ɰa�J�v�@�j�-FT
*6J$ڢLb�@��Zd:TR�Q
��E�B�P�66U'
��:� �`��kT��c�
���>Gå�C�hS�8�~!����Z?�����`��ӭ�~ʱ�E�q��7����n���������oF�س�汛��M�^*�]�
���K�᚟M��'#����;Yg�3��i���]�1��}	Y���2�InqPˈ�"���nF�%;5�([t���W5n�PfέV[Zb}V$���\�]v��M�#����I�)�-hP��,>��u�Si�{��s��9o�JSK�[BQu_b���tsgJf����@��r�֧WCB�
ҽN�v&�1�N�$w���S�B�	Þ9��ӗ��N�_`�W��]��4�SH7������j��� ց�1����V�rJǽ�����#o8[Ȍ�����Cb�9�Ӈ�6��%��j�}�_U�WmB���&	Kj�5�%,dʄnc[E�U
n���W��`��h�R(�<��s�[�hy%R�T�/c�?U@U��hI�2�:���T�PY��n��Ӗ-'�����[~ 窕*�.K}�� (��$�{,�k�;Zj�7aФ�J���9H���Db�Ըv֬R�q�9>��z�K��J�v$����,T!�Y �),�]�yP�j����xl�T�Qw�L*���R���|lD�9�+���_�|��i�XGn�L��4Nta���Y���"�ͼ�+j�cv����d��[YAfc5���J�Y��O��U0Yo�e�u�أ��V��ş���������ׯǯY�ׯ^�z����=z�1�c�c�1�c1�cׯ�ׯ^=z���ǯ^�z���ׯ^��z���ׯ^�z���ׯ�^�z���ׯ^���^�z���ׯ^�=z��ׯ�^�z���ׯ�z�������ׯ^�z��z�^�z���ׯ_^�z��ׯ^�z�=�z�9���=z��ׯ^�z�z��ׯ^�z��׮z��ׯ^��^�sׯ^�z��z���z��ׯ_�^�ׯ^��ׯ_�^����ׯ^�[͆��]�MTVs.MPz�}��aF�_G�϶�����hL&�oC�u)V����ifu卮���M_]�Ύ̏VSޭ�ByȞ��;�z��x;�����_[\�+���"�d��T��p��\l* ����F�,�!��U���s���K�wh��ԃ";j��Ʌ];���ɩ�'X��7�y��W	Od��$�`�Dތ�uü��Rf�ﮱp��-kM|�H�7�;Ň�I{���_��͕��J�=�:����w����+��M%�̘��/]����>�[�=S�/���$��8���M���z����J���c�}����%���X��8�r�nٷ���C��Ti��̶��LiUӓ��;��Z��î������y������>̼5���{�7�W D�RcJ�+S�Ѩ�+:إ�0��m��
=�ċ �z}ݷ,Q}PB����1�sݮͫ�l�:�J\�1�&gM�䤪Ω,a��֯`ˣ��`9����r-�!�I$̖����s��ks�K!9��:����:��*�4��OtQ5{���m�4�7(=U& �.�s����[�����w��pIm��n ��rBE+ţDS�ow��Ͳ���[WK�@���#
� �-�|
�q�s���e����o{�x򃗑��=Vw������zߏ^�z��ׯ^��^�x��ׯ^��z���ׯ^�|z��ׯ�^�=z����������z��ׯ^�~=�z��ׯX�c�1�c1�c�1��1�c��c�1�`ǯ^�z��z��ǯ^�x��ׯ^��^�ׯ^�z�z��=z��ׯ^��^��ׯ^<x��ׯ^�x��ׯ^��^�z���ׯ^�=z��ׯ_ǯ^�z��ׯ^�^�sׯ^�z����랽z���V1��1�p�1��1z��J�j���n��J��*PH�:uJ�:v�W+�)m>��������%�h�D,�i۹W�]n�3LNȝ/v�*�y���jA���n�LK��Ʀ���X?�Ԛ����R�1ڕ0�����twW�f�	�'S��v�#�R9���Vt�ؐfd�Sr��d�'�T�ϩ���������a_����n�0Ά[9����μ׆說���C�ci�*�U�2ȓ�r��dl��֚޲�����fNMaO������w��6l�5*�"�[P�:ܹ�y�BY�{���'Ǔ��Fh�6��ގ��@�q�s��w���N�˴�0���v���©��(�=����Ď��"����5z�g���%m-oo<����WsV�EX��o��)B�����mR��vB�+C5������"��qu�kӕI��nՕwo���ζ�(�(�q�)p��7b�E���5��R���_6e���-W*����x[XT���)\r��p�\�ʰ�ct�5�	I�Y[��!��v�M��y�����8�gV"Hr��Q���S�z�R$��a����s��v��حj�l���H$� a�S*b�({sT},�ԫ�4��+���%@�wʑ�0p��2����8H�\x����P��M�N��%�n���곶%�9�b�=+_-�˝N��.���*h9I���K�;�̙D�Ul>�	j�\�x)�ǻ�s�w�V�{S�f4_Xf��׵��h[I5ٸ+��ΛTX�:����$�Vo;9܌��5m���^���vP3���=�����珯�Ϻs4�7�N^&��pMߑ��Q�nۮ�R,V����'@\��WN�S�ӈ}ٝ�>x�:�BV�=� N����:���m�XrTа��u���$ܩ`��WWu�X�͉��C֘'K+"]�+h�b"� ������������o��F��㕝�f���Ո��b�yG�I\�mL|CNl��;�:�m�_L�+�p�勦��[�q��V���B�� �n$\w��N7Y�u���Q
y�����ٓ�`���V��L*�:�tH|Z�t�J��2�����]���*�eH�t�b�VS�t��F��k2�M�����Y��#(39�N��cNǀ�Npy����V� ;f��f�)C���a�κjzkW�d���+2�@3�Z1�O�ـ 2�\�8wu<]�G�x#��YI���9���]��wݨ�Bu7�t��q۾u�I��IOB��سT�5$,z�8�:.3����&��۫=�U�{��6�r�2j�O���	Fn�ܷr�k<��=�T�Λ�y��͈�֙�B� ��e_T&]���&��˟ս��ǐ��T�ꯀ��jd�{Z�J�����J�'/�p�Z�!Z,��38��SX�=�vCC��!����_S��yWU�\���g1�fcB�m�г���|�Ԋ5x/vV��_l�V͕Y[�]
�w¤�!EkfNCs���C
��ѐˋ�2�#��3:5��6��"T	7���cy�+��'A����6�5��ҷ�� �%E��vhP "i"�(Ņ0k��I/{ 5��q]6��}Qd�j�w�9��9�M�F��*�T����m��rE��K��'W*���]�T[	鷙@�j�՘C��x9Q�S�̴����ڝ[���5�)�
ڠ7�4� �J��p�U��ɠ��Ǒ�m!�(&]3E᭹P;�Wb�D�����h�����T")̽J��ѧ}&�f���P����A�p�)Gt*d1��&�e�pM��N;V��Ji}�7�ri�5��tDB�����������f#oS�$̸���J�w])@�A5ԇ���F@B���[�"�ܾ\����@��שl��k��v�o.����e<�v_u��YcZM�;t���_l��oVE%��Ol0�Weq�J�
\���*�M[���3#�z���_F�Uշ�r!b���`C��InP�ޝu˩�v����x�.l�*����v�R�92�9�5�lKW)�]�6�󍋤cIH��$��z0��z�W�Om.���k��ɋz�L6{� Lqu�z"&؝m^Q�Lwp���gGHkov�Q�q\4�`R���	W+4؝3���xz�a����䭘�ݭ�i��J��YEVQ�94���w�ޥ9Y	��TH����A����ӚUZ��M7��H{�*�ef�L$��z�J�D������t�)��#��mvA4�S�f���j<
nZ�V1�7 w��t���:C;f�.3[Ti�дЫU�;)��@�u���V�ɭe%�(�^���X��P�#�`e&":]v2�J��4I�g�x��,�%r#9`�38�҅`���̫NP�^wM����	�z�mp��]u���*ٗD�\��d�&���-�Ep>H�˲�6N��QuZ�;�p	��ju�������M'ҵry��j��'�bW��'��S%�l�Q\E龲��:ʼ)���&�����`���j��:V^��u.��p�(Y�lR�l��Sp�e� �vRV���	�M�g;Ό���ъ�J�x�-�#EуvJا=�D�Y��س⅋[G����&$�Ժʦ��7$�o��(JΩ��\��;���o;�^��6�A�Ў!�&I�v��d`_e� �P��
}v1��۝ip��5(��h�r��v	*g�qC:�*8�Q^r�V����0���:S�����䮙�Һ�H�V�F¬c��-��J�W"�Zq>�GUԦ�Xtå�5}�tE�+p>��:�WK�8�b��L58�M���D�e��7 ��*��x�&����������ɒ�]q�!e�L4l��P�r��v��ܧe�GT�ڥN���fj�:weGZ����Ư�eB�;��,��PW����Ӿ�ܑqӲ!ڌ谹��� �-�ר�Ҏ����&>�;�ܡX���ډW[�Q�	��s}f�f�!G[x,/�����iX��.�`6������2��e��Ze-
-��1X�\�V�/>g �G>�6�ѕܘ1�&fZ��~���iu�%��x�[����7���K�:+,=�W����Mꂍ���0�Y(��Iү���|[�SpJ� e$���	�WQ�D��8YS0#ܓU��X2��xj�R�w���y���N;A]r�+�>�@Ӡ�k\.���=`��R��z;#�*ĕ{�G�f��;6X(�ɪ�>R�%�V�XwRb�׎��u��R�v���jH�xH��97A"H�!���pX�۴���`-��D[�GG�{j����&s���*��L��iЫ�B��`Me#�f-غ�'���0�r녓5��ǰ�ܬ���h1cUZ-��.=5�sq�rp�I�Pl�|:�r�f�:�dO{�=�q�؊�z�_i��nQ����x��oqc�Z���̝�u�����U}�&��W�[P�4��V`\�v��u�0���_H�᫨��".��e�e+��D��N��t�*;�U��(��h�n!�zncɒ�ì�+���R�S9�Q������Z("ye&��E;Gs�x@��d�kn����ո6�͚·[@p��2�p�l� ������m�A��xاAL�����r����Z���Fj�z�|U[�uo+E�7��?�JP�=}H��Z����&�f�m���K���=�obB��I]�Z� T.�Ѩ%��R33
���MK�5oIwբ�v�����䡰UT�8���R�^��/q�G"I�V�y��\8yV�m
�v0��K�ݹt�5�5���#��AN5�oe��v����B�S�C%�XL�u���[}�>��g��\��[Q�b�:���!�����aP(&��t���T���Ӽv��	蔆�	�f��j㖢u�~X_<ރC�b�(�=R����9��:�t��#�$κ��IY�=�U���X���ʚ{�j&�9�#�-���Q�1��v��ѝ�)�ֈ�\�G��z�Qy�x�Hz�L�|T�v1�����%{]y��Cy�3���ٛM	�Vy�G[��[�2��Yѩ��Z�d�=NƁ�rme�8��!Q�/2�Z���%�.X���u)Q�WY)�������H�
T��ݭ�S�oj}��� ��+S\�f�r��HZ2\����Nv�ו\4buN��c�L��Ï���̠�PcR�Z)�UFo7��֬�� b�@)"�&����5*͵���z�aZ��\�b5>�ϭ�7&��d�$�y>���̦������Ǆ{֘�t��]�{g���Ż.�.�"��H�54�*�ʅ���m.��g$��V
��S�ޛ��;�@'�*_`'W^.��zkt�CN���/\\Q,�L�VuZ ��μ�R��Z�J�������`9,*j���cL�o�샍c����aV�#Yz�`]o����h7�C|�5�4+6ZS1c��؆k�!�AՓ��Cj�c9������	Ե;k�j2�K��,>�A����	O�Wt���r�5)��^����n݄��ia����+��^)�/K[h��YMc�w�V��'O��lC�V���!��[��[���k�^���I1������9����'��~z����[��^�+oE�!�Hf]�3��i{���:�e���R�Kɘ-�U+�ac���Ҝ��!]X����!��lj����DԳSA�������7��P ���)w�����t���=9�H�UkZg1Qub�3Z�ΩBP�� Y��|�֥x$|��%��� �:����)�|��]f��R%�Fl�Ǻsy��{�T�w:����CC�.���)0r�1��v	H���:.��ͤ���&><:^j�X\w�C&�u����ZA��P�F�q	Yk�j�j� �r���fu-\(������'�.���m�Ta8b���V�t��)K�hk�����<�$���b���_=�����xP��]p\�Ɩ\��k�Sw�D:8L�޵��Ɖ>��n����~�oioWu�V�(��c�w(p��c����rn�ᗉ��3`���@s��%�L1+8��6�u]bu�!��b��Te�6��r��4�U���ψ��7h;�.өs�9ي�]���x8S����ݼ-�X�2F�C,U�ݽH����뮙Lڲ[[�\�ƶ�k����Q^�P<�:{�{}<�w��5�y���-Jգb��j�֥igO�W�E�$���
������� L$�n���Fb������WSy0���E,*岺Y[�__qbj{�^��7�1rrH�p��iV���J�CG����)�T���BЩ�!��K4Dr�밸�[sUB�F�ea����W^���������X���\S\�gSbkŕ��p�B��n�qP�5LO��.�6����嬭��r^�:mla"��ΞӇc���i�-N��ls�^�;�=�0ր��wf���"�o��wE>|��fȋ9��b���`#�Cہ��ѩJ�����%�Z�>�A���$S>r���?N�Å�Pu���c�y%*�V)�ʎn�t9d �۽��i(��xf��hom��[����Yݓv�5���6J%W �yu��C]1��i<�mN��uRoX.�w�a�q:f�:�6�(���{���%,�l����e����j�a�'vh煜����҄(lyy���%�-AM�c�>��&�R}�*>�;μ���޽h�/�Tx����kqM:I��Ui���m�ݜ�g��oU�Ҍٱ<������U�{�6�^e�0��)��54v'Y��4M9 �Y.Ii�_d�����R�o�}2�ۓ�[��s������'f�w!��^.����P��,���i4� ��M0�	���2�HSt� "�4�$�h���d�a�	� Q`��F����lU;�2��@_��@x���R��:�2mO���_^��^��z��������ׯ_�=�/�@�O'��� r_J�q�T��>�����=z����ׯ^�}}}}}}z��� |��~G "����UUN�O�: ��t�^Z.�����(4&�Yw1���@r� �6Ԛ�E��5y�t-!�6ыF��i�EM����b�0h*��\�i���et�((���\�-4���U�Ə%���y<���h�����F�`�Zaт`�L�3�j�|ëV��I:��o6�w�p(��'mG�y�ȼ�գ7'�THUW0`�`q��
���S�2ܱM��ם���-%�c�V7)��;J���^Bu�� v���;m�0^�ޏ.�����r'ˇOp㋌i�j��]���,Z�+�T<=<��ݩItv(�������WRt��O�٩�6�����V�V��1ӕ㚻'��^K�k�Y�i�W�}�ם�hc�]0%=	�!;���x �U�t3����P�-��߻�~G��|�����ݔ�o�4����x�#%G^�1ک��~��υ���@;�i�uL{ݣ�_����k�����\�G�kIA<�k��[��
UU 䪄_gK�mT�5��f���u��������;yξ*�}��{����g-9]�oE��3���nÙ�f�����r�4��x��Nھ�M��*M������7��j�=�D��z
k�g������];	Z.�{���(�������ﱟ�����Q�NUvX�yy����X�hk�f����^�ݛk��y߳ޓ�|=>�KQ-�G�/}#�3�&�G���;7;��~�%ڇ[���^��[���	�Ux׮W���"~d����u��u+�w��6�
��z�u���7��v�_��՚2O��)�t�[���[�ɧ�e��/�C7���{ϖ^r��I�d�K��gV��h�ɞ=��Vn#�׵�����||a����z�FF/�d�>a���~������{C�����74���k�c�OK u^�r��+gmU+�ƅ1W�!��5����t�U�r���s�/�f���P�Mན��㽕\�"p���__�VuO���''����#�Wx�������S�Q�����ڰ��t<�~i����,��Vq�7𦧬d��M�F��n�Oh�b�S����ק��e��5o�{�G$��W�G57����xQ�|���1����{�'y(�v�~�{����L�J~|ǜ���Xd{��_�Wy���{�t�'tW���$���O �z(s�խ��/ٟzy��(���v!���g��ݏ���s�{ͩ�̵0y�3��c[2�=�����g��K�ً�`_�����y��'c�a�U��ڥ�Ɛ�x|^�,s��]ˬV#O6�K�������s���vw�$��V#��F���}36�eFd��խ�=�[�n��.h� 4�w������f����ǅ��l�1i䈮��Nj�(8��"���4���H�jDiӮ�x��ܻ��m��/����o/5�|����eΌ�c�����<{c5��^P�����|P<�ܺ�|�2I'l����C�G�h���v}���y_���y�%p�	ٛ�{��Hή3}TU�`>��tEP�Gϒ�����w[����駼D]���l*M��5v�t*���@nͯ=z3�#�5���}�0���x�t�����$�;8�u[L{wm�'��f��n��W��o��U�I.�Ц����5�v�g+��Jq�WW�=�wN����|�����{��k��kz~^f	�*<dͪ��q������'���x�}�s�b��{`'�F���HU}��}�j�����;���ח�����jj���+���6��?Z�'��vzV�f��{�6���_R�}龼�\���-�?G�d?X|(k����]�V�kgφ�����4g�:γ��Z����_E�ҽ*H�P�w�^���\ 2�Ď�>�V�۫8x�
�o�Y�����lTgK�H�{MY��wT���5�V�w9*���֋�0��X��u曼�!y���\���nS�g����N�w	�J��������mx}H��9|]w�U�^��@���wM|�W��[�Y��o���<��^D�jڒ|9����E�ՙ�t����v��+���|�S�5���q�.����|����5�̪^@���P�۝'���v��&rg�w��莿]iƌ���c��m/k��M�=}��p���Y����sY �'x~��_W��w����K��\�������sA
��ҙ�k��ӖG����2�AeT�2�z*=Rb>;�g����ʻ��J&���K���Ë���#��Wd3�-�
e�}��3V)�uo=�r+���*����9�������t��}���p!�f�������	S��v���Vp�/{v�t�d.�/���{��x��J��i��ϋ���8�}�ywns�}��,&w�3�P}$�)�+k�곊ߧh��1tN�j��M�M��:6����L;����\Ƶ]�fsϐeڮ����58^��a{.��M+�+s��$�n��h�����ƍ ᬅ��i�Y����y�:C�AQ.c���h�zhջbt�������Ǻ�޻\e�۹��W߶|Y���D� �H2�$��xx�C�������FH��;g<~�eV�vQ�1���܋>��c=;��&��_��Cd�\��ը}Cڥ��ªg}阃���������)����~Uӕ��~5}���t~��*�9U�{β�Hja�M��~��k�S9ٿ}9zn��uEG�����h�T6���k�]�L�۞��R�.�M�}e�x���ܲxz���/⟕�<�^�7B%��ڂA��ܹ�]nI��t��|�W����s��>�{���2�b_O 2Ь�z<���ni��2�K�P]^�����^�y<�Wk�r��9��>��ȩ�Ǳ#!����g�Gc[sm�V����W^��tUH=�j�:�a�^Z�9M�/�oO�����c�-/A7�WzKT�^�s���l��}`��fs�i�p���_U�����>UNW��}�J<�ϻp���z�^���q�PtF����۩ʋ���2��[�K�1G��Ax�q����>岔�uؗ��]��}j����G2� 9���l�,Έ"k��쳡+���bE�)�y�L��W̡�v�p�7/+��E�W�����uM�*m�xxy�yۜ^�2���󶷻'�+�;ݛ>�y\j�:�砠�W������2uv�^��˰|��#*w����w����/w�s��fE<�L����[�exe��s)^[�%��u��<��h}��(���:�|���yow�Ǖ�g��f�S�W�uӑ3�K!Lϛ�z'Ar�c_������혴��ۋ٢u�(V�^/ت��A��j.�Y�A�.��yg�]����Kn�����Ԕ���$�|��u��տQ��kWW�pY� ^K�_w�3<�c���OP�}��\��'����UV��1k����q�}���u�ڲ�Zݽ�����)R�+����
�s�k��Î�o�۾��z��<����]��	���#��Y���g��bv�_���[Ӏ8�'({����9�N_��j���ʭMû3�'W�Oz�s�-F�"�yHJY~�!�<R����k½N&��uޗN@�C���� R�L�z�&�g؃�&9��ot��(�E�*!��C�\'˪n`xF�6>�fM���[�e��q�ٚ��;�,��,..�=�+�5���"�?�����R��)�=}�zk'l?J2Wy3U{� ���>>Ky�i;���kn�����.Y���c���b�����π����X&wʫ�n��c	�^���]E�od3��������Z��	i��g);��Y��ә�{���=\'�e�O���p$/o���.�����{%{��ҳ�S����}آ
c�n�U{��b,3ӧ��_��?_�'dz���V�g��/�ӗ�����پ�(<�j�R���@��?k����yn\��؁U������W�]&�{1}~Ub>A�:��뮘߾�������߯Y�re����t�2�������b�M�ݠ�B������w�kF�>����p�����o4�k�wgtJi�Z�����~�M�����y
�w��o��wN���2��//��Gu��o����β}�I���o�9�R��Y^\W��ޔy�
מGUu�̙Lq]����8U�x�����V�oV�2'�� �M�V��.��"xuv��Sn��<V��N��ga�~$U�)ڵ���|�Zs���9��Q�)�2M��K-l�ή�'��S���q�29�w;Oq�f��s$z��\o�����A�k3k�|�<*��y���&p�<ܣ\��q\��r}��wG�\w���$�؞']�?s��7x.w�1V�|=������e ��}��[JPJ�b	\�w�t�}�խ0�Q9��߼�??n0%V|�¯^]T�7G�:m���.�d���Gݓ�"�>;K=N��۬�g˺��Ej�QB��2���JN7P{��ܛ��t�R5
�L��������ow�]g\N�=�/s되�u>�x59��R��Z��d>D��#'
��0�y?^�{�f�<߶������;k����
����es��LUR\t��Pyg�{�W��{GاxV����X�F���ׂ?{���2��ǠY=b�z�ϝ�*�5�zr�'��񙛚�Gs��sݎ���^m��[�⳦�+D��|�`8m6ѷ.1���s¸�z���=ڶ�H�tł������\���;�٥٧-�Jx���g��Ԡ��bIﮧM]�<��x�'O3�Ѻ.z��߅��υD�n>���_�|���4%d��͑<����ڳ����K�GH��ó�̼T�ٸ����?�-�5q��%^��;� �i��5�����9ō?U��vyyU���W{�]�������ϻ]mn�]g�"�3��ܩ�³��2+vgc� ����F+}�(�%���z�Z��yǾ��q������}��=ﱯ���ޝ�O;���O�ٵ�.n7�����{skUz�hj�$Ձ�\�'����&�'z?��eyO}qמ�ebb��z�����cd�>s�z�A=ua���5PN{�s��j�8%�X��]���qn�	�Oן[�����]���V����ju� c������/ �֜���oN�֐݌_0�g�|	�@����3mnLs�Uޏ�x�錻둍�H��Ǻ�@�i~�7�ծ@�]����S28T�����֤�O_�]��\�z��W|��@/��u����m����ywe��p{UY���s�WW����a��1�:���:��^Mӕ����`f�Q�"*1jl#l��P�~�_d�6�B�KY9�FB}
4^��`�y?���v���N�����2�}PW�]�bulpwq�|�o��lu����[�fSTQ�͜�fv��f�	z��s����uu��ݾ8��xxxaٛ]��ޤI�!,7bs���O��/�OWb|����><��wxg�b7��#uX����P�6���?�纳|��Z��w��K�����:���������9�ޒ����Y�{_QW��/�{���������ׁ>���9�{��9��=�j�Q�[�-�7Y���x��m�i�\[�sLޘ��A���5��s3�}�ݝ��S��_�W����tܻ�^�3���a����]�;����߫�J�}oX�v��#µ����������>�tj��#�sp�����9�m{ٓ�n�Xx�	z�^�l�+�z��MT��E�c���嚮��3)�uW�6q�B�ޠ���SN积�� �]�ю��C>�o����ӌNe���yΌ��R�p�H���*���|�|��}��C�����-�lV��_�<���������}w�%�%����-���O	J&�n���m�U�P����JR���j�Uͫ���m�W�����N�bB2��u59Z����b��s9���]>�uTٻ�E�b�]�sے��@�PY���E�F���>��NvG��]��n
�.�͙��u�l�^��L+ib���)J�޾L9�y-��W�\�b��Ce
��lt��{�Ae+S^	�T�	9Z�N�2�sE��F��T�&m���(��M�)�o-Ns�s cUJΗ3�Y�:�R�,�m6��!������9�����3.����I�C
�.�ҔQ�^��ң35�h �Q��_*֧i@ܳOW{�hє�S�Ʀ^�1�\i�P>�ӝß��Qٯ��@����NjN�
%2l��W����s4F-:���5�n��ʮjn�MW_WAx��X�:�!E&$�s2�<v���kL�$��EGJ\Gf-H��2[�n�(��>9{Qe��Q�V ����$*�Vl]C��k0�Ҧ��Ņם�{�9F������۵�nf��N2�iih2'���*���e]�	����X�_^i�L:�\�"EXc�(t�*ܮY�qشL<E�7W�9Qs���#��՜3P�N=4xE뷝��=�z�+n��gU���rn�ĵ3׸{��R����/{����<�wR�i����+���hx�h���pJ�5��&��&���Ղ�ζ�h;���DMZ`Z��ȉ��E���iﶒ�W>\:N[.������/gZ#�����3)>���ݡ���6t^? ���e:�_kT�0�4�|&d�J�;��!6oMth�!X���õ���kV�����`4ډ��GY'\�w][B�V��s��)�ڵ�&S�n�nw@&^�ӌ���\�d�,�9�Y7BJbpUv��]c�ȭ�\�)����p��/>�¶�]��`q0����V�T�ʝMI'ܪ}K�-�-�s�e'9����wR%͠$q8��)��]3F*c+�xފ�z����a�oE�9���Q��8ũW�����XΞ-kC���y�˒:�e��e���3z|i0�ˬ?[�c�^U&.s@Z(T�.�5}zB�5�*.'�U��+_ 7.��]�83r�u�a�zx�#�K�G*<��q���Ž{ ���W�o0�i:4+T/�Z�Y������s.j�c��]�:��̎���@��Ms�6��+������VYš��mA>b������罳�pc��]�.�1��36�:ܻ�ALn�1Ob�W_h�kz-�}Y�a
�n:
�>ݧ�5�������;{`�EǕڸ�ۉ�G�l��`1n�I��'2�� \�+2�f�wn*bv �p�F�? =�<L$~E����W��%QT�'	S	6͔�S3-EL3Z1݈ �5�\���9���z���~=�z�������ׯ�������SP��$��+�clE���|m-�.�m������\|��ˁT�8��ZNǰpj������}������~�_�^�>>>>=z������� ��yɤ윎�⠴��LZ9r���foKZ<�\�#AE��ŧl�fnO�� �9Q����#I��I��h.41Q�\�{R��M�<���`4�0�����C���D��sc�t�h������{94&��*��My'�Y��#�s!�!��U�rSpϐ(��'�? "��J���5�!�����9K��*��j��Z(�y��-F��4SE7��~}����(Tݍf�![��ݦF
��q���-�v����%*W:�zJCry˙a�3��i���＼|||��^nQy��G�h���ד�O�$�-��4��i��9�8��}戰@r5��qbk�wA;Rz�hwWs��K=�\���,Ȇ��[}w�ι��,8�o r���0逶q{Z�6]��fl�2��P`o�l���߇�?hte���q"H�K>�����A�m��3:.]�߷ql��y.,�t�1��l�g��ĘO���6e䍿�= M���6b��^���QҶ�7Z���N�>�{r�'YK=4��%���ߞ��^�K0�.ׅW�r�rЂ�u�5Q���d�W���䬵�6Nɤ<�ٌ���E-�(���o'���Q��bh���7�ϝ�Zq�4[p�y�/��Ȇ8�ۏ�5���Z,m�)7X�H+b�۵��v*g�ǭ7[|�:�y���d���h{�E��!�H;Y����3��1�I�p0��
V2M)�ټ�=B��Y�ӣ:��������ٽ�[�ѭ��,Di��0= �7P��k_K�J`�:Ü{zs�<�̿%#����O�L3��W+[:և��ɑ��pƧ�����Y��9��� x��sf ��c�G����^�c��F,�T3���x�w��:]bu���̝�ܝJGOS�x3���Y��
U�d��MȪ\Ŗ��`gn�`�<=R�6��:�d���4�@�wU���b�������18���J�����"��Q�h�q��띩VQ�TL�5���q�����|>c57{�{7��}�׏��n����k��d2�0Ϻ�	�ޡ1�3�>�P$��ʬ[��([DU�[hC�3g2ԡ�����t�[?����$]�|g���CsN�����&[wJ+$!Q7�կ�U�O�ݻ�B�:X���d��[�}8}��j�Py�%U�!���N�R��#Zy��cR��|�C�;u��0߹�[I�0������n.�F*`�E	W�2�����b���3��Mef>u�}N}�[-���"> B�f�]���|����޺|ϔ�N��>�+�8��Pc���LU�%��.���]5��qd�J��(Pz��t���C_�m��A8@���|�oo3WcV���H���M��h{�w'�pe��i��z.�G43gH�8�hk�|�6|��u6\��L�+�˝���S۝��H{���x|��8�j�^Ɏ���@��kyǛ��0�*��ߋE�*��k���W�ۋ/5}���߾z/����7���Ɵ��Bv�焗U_�vJ�8~�K�<�(`�^^E�;�j算�>>�6�Q/�Wz4���D	���	�7��4�<���Q/TY@�N��m.ݻ���-���@���҅V�6V���e>I͜Ź>��B.�ڈ�7�p�����z=�c��N�r�uc;m�4�X��	�̽x�Űf�n�|�q��HtŻ�k�#]e�\9�����x�_2���Y�hQ]t����;�#TZ�r��ɉAH*i&����������T�N�ݾ���c�����e��u��i�t�>5{���{gò6�8ᡬ��E'oJ|�}�+))�e��_��[�1^��{��w!^;7d�|�:����"�7��dN7�1��{�5p��TU41����4�\>�V(��C�r��3/w]�U��Q�^f��!�]��OF<����\
�ȴ���B��}�Z�e�F�&�~�<��ցO'q��'phyZ��WC��ӗ~V�
�����
=�{�s�K�"9���b-|��s�]ѧ��� w��:�\�4�P������*2*\5���!��#HI������n^%��h ���`#�+��_OC	�u)���y�4���ڛ����@fH~��{T���˜O��({m�zl>�H��7T�����(n��a�}��:i
�}�N��z=���s�W_^�r{��1��488�\ ˚�stˁ%5�V�C-(�HW@�ҹ�z!3�ɰ������Yu0��ӏE���q`��y�ϯ�!�2"���Ȩ��H�c_c��3���i��suy�v3�����O���?��NR�=>4�Ox�7G�t����Y�d���t�����b[cٚt�!tpV �=��T�gyR�v��ɜ�!K��n�!o���\%�edɗRgb{�J���*�5ǪuqZ;�BXV���X�\�fЉ�(�w*�WMl�YۃK:�3QW�'�h
&����u�'����������y��]�����\�)6�����D��3�G+a����t��!�?Ro��Ƌ]af؊v�^��g'��eś�8��@@�����j��~$o� r� ƨ����>:���0-���5�N�������Aڕ���}��VC��c������m[�@�@���K0e���x��^Ӟ{����79{��\����,j-l��C3��2h��t^'�#��}d�6�ծ��f�+�j�U�*϶�G��NDذ�~#Б\��'���q��&�9�ͻ�:�"YJ��y���{%�PZ���c�P��Mlؚ]��4�(������K v�I�}-��l��e��ܗ�����H �|!v�#yk�	+��Gf�͑<��U�)l�5�Ψ�l�Z�8	L�C�kGT�ʸ�<L�k�	�n�����xL�����SD�L �>�=�]1�bj 5;$N�ſ�rͬ؍���v6P��f�"ޮ�S�*�vz7��Bm+w'�,m6��9�@<��8�bfmg4����	�[ԍ�b`�9�Nq���
�Gm�<���S�̱�Μn�_]��&Ȝǩ}��P<yYf�1�u�)E��
��Qܭ���j�,��6������
f�$v��W�*�^�%k����}u1v�w!|�1��X�J��^j����fL$t�
��Δ�4�f������G����P������ia����+�o�:~�>�ѕ�K�޺���Q�H�����c'u�y��L&.�����d=��w�ן��{��xd�s`3ώ� 0M\�\4k#0�p��ĝ$w�q��s�%�<����@k)D�Q�a��1����?��ù�.zA�\��u���Ӭ�c}=WVr�������Y�u������ t��G��P]�<��u���)��1y5����6e��u4sn�O� ����n>�`�s��qr�m�}���0��zM)l��l��@��Ȁ�d��º1W^4
�����^�F���~.E$��b@��t���y^�q���QG�C;�Έ���Lr�on�̀��aߚK�7��4o@g��`Bpi�{=v�ӑUsy�ՍP0ǯ�bk-���EWc����$
���m�E��F�����d����ĕ��=��}�-���ʯߓ�C���d
�ge�Ys��C���(	ƕ��v*���ZI��&�2����ߝ\�)�Eݗ�&�V%GA�q�>X��V�C�L;Kd�m������>����9d�����c�N�%���>Z���S��{�c�,]�-P�t7��_u~���]B ���6�/����+�u�.n�W���t��4e��dl�<�Lޝ��c��.s� ��f: 4�EnT�ٸYC�\��{7�����,��F�}3s��Y�:�)�/��Lef_�����y���y������ �"�gY��DL��N���	9!(�j�r�97�����A�|�-U��6�cp��#�귣F_�1���|>�O��Y��M)�o�N*Sg�
PF��x.b6��:�\�cN����go!�E=;-���-dg��`3̟)�����bQ�F���x�s�2�z�]ў���onM�ƾ�|C�,�
]�!Tuˑ�
��{#�Yֱr��b�����r�^�v,�U�T��ܬ�Lu[6�j���.��ϻ�W�Ph:��v�0��8��p/Ǿ���\�t�;��V��N����2�
Z�CH���pn����vz@ҷ`O�+/Fg٘�6,��:}�ۚX_��פ���G�YKM���q��8��},���y�4��Ia�xW�(q���I�� ;S�Y�b��`����@SaCz�c��:N��&������䎙�i�����dǦe�s�����@��� ��O'E�T�}n=}���P����\�����[A4��%�����Q����kL�,��hi�z���!yj�9딵~~Z��ۻ����9���0v�$�Kog~I��3��Vh��m%x�'7R��t6�z���̲7Ì4�]/s�y9���[�}Y��8:�0�w��*G�ٸ�+]׷���cM�9=��2]j�]l��¦��3����G�|j�/��^:�yNo�`Ц
&�T)3�ח����y����-���Yw|೺{k�o���0T#��@�{<�j�3�ֆ��'fO�����Xn�Ia]�۷'�ia���:�G<I*���o
�D��x<��K��)�H����_�8�����x���ݹ��2�lp�>��{)����7L��k��2F�78�ٚ�g; 3[s0���:����Cl�c�9�7iT�Aޕ8��4
i>s�j�@�O<�U�D��x��Y�q��4�Ε�Ә����i:�YSCk�����*γ�d	�tV�xZyM�j�Vd?j��Ak�c��{�3�\=P�,--�ar#�n�l��E�G�����c0�n%�*,񑏱��ׅ�����cc��%R͕Wh{a�y(-�X�[w#(od�4�`1�H4�o�Y����V���z���n�v�����YԤ�!�pC��\�e<����>� �S��tt]�ϵ��4�Y�Z����T�c�n�����y�7�l,��=b������y<F�q�m�	2�} l�P���u���V1f�wru�ծ��{��˚�(q�sYt�P�EoG����S�R��⸶��[��gٮX�z�b��g�[Q��T�L[�8�,�4���d��'X���s���h��mϗ���C5J��7�W�}���O�g��i<_^�i�;��bJ�����ed�|�}�V2�w;y��jl�+C��Ӣ��M\{,S��bK�F��Q�a�<�潚��^�~?��7[.Z�s�'�.�O��}n2!za��7�g:D���os0��L��W%�W�m�K���խ��z��[o!��h��A.�9�������g�yG��	N��}V����E��^�3vw�����鑆k�s� .��e��]�-�?�_Hc�p���G�B�/:7���Y�v���:�V[�\p�=���b|5��^����s���Ns@��?�t�FB�'�,e��&2$�i�ù7D�np�%�a
p�0��e�)���ɏ ��U#C��-�2�l��������E�]�&�֏#r|À�Q��|%�`�v/���[]��ox8�ޮL&�3���ُ��_n�)B4Տ� ���nwf�� }^0sB�^vծ$D�ո�l3�p	7O��_S r� Eϻ�^��ZV[�n�է{6gP�C�����;$����k0@�j�L�QGRw4n����z��o%>6j^ˎL{�:�ؗMv�=m.3[�%�Ԟ�ȑ�u���'�l#�=t(b��mR�b�x��QGb��#�1���C�������a6}��2�,�gl���~�	�.$E��{��~U�j��R!<à�e>D9�R�&�[��l6�7�¸�0�;1�^Ǳl��ӬX{�����2��Y<a�U��t<}�y=K�^`B�7� R�]%�-��4J�j0�d�Y�9]��Y�se��BT��
�oU���U�~�����M��:���K{H���s�(tf�)����r�,�]����m��� Q���˸�qB�!=Pr��N�!�!�� ��.+��C@΅�:�ȅ�0�oy@v'����G­�����O|�>����aa³*�A�ٷ@q]�~/9�>\���1͡���i��_��yE[a�~�׬�疋j�v�P��
ٹ�b,���ɰ��q�@����<}|��`���SS'��>.�Nu��yv2X3p�W���d3�dq�6��8� �d��TÑD��Fv�X�d��都+���Ϣ)���mT�[�C��8���I��ǿ:~+���� ���;�&�l�5��CAì0Ѿg��2]"�_�t��xý6�&���ڸ��wF�5{������f{���ܔ�4��Yݢ!I'�nc/:qf������{-�u�?��e��@��,�dkx����NVM�3"��Ur�.��i�ݬݙ����A�����6�ɶ��R4k8s]��i�v�� ��pZk��;� 9��,��Ce+��Z���S3���m�̈W@�/�ͱ7��_2�|2��z~(�R��j���ǾP�[�j��'+_3�Ѵnu�|��YRd�s��0=��뗙�ރ�r$&(�L��P�]�vov�sF�ɜ�!3�[;&:żl�h��B2���8�["�;uv��֖N{�|9��HU{���?~>��y����k�u :i�͆<����ԙz	�_���ţ2�����"n/wą%��N�4���M�������$q]�c��r�~�~2ͳ��F45���b�sH/�E�f�``�#�8�Ve��Ti�x�C�$7��3��:	B'yVzh�O��Y���jq����t{F�����:����?=�j/�r��]ӽ�y��g�/W�>�u5{�=<�QT�������'V(�g1L
׏3Q�ʛ-Z���>u)Ǿ�=��9 �µ�6&�$�u�{u�2Mx�)2�1�1'�i�ЧK0��c[����*v��f!�4_Qq�P4�����.�2�A�O���ݬ#�^:V2M�ԟzqO�l�ٍ�h��:���ZP�d0x"�r2q�R���/�~r�&�Iz��,f�� K0��J��J;�fxUdj��mD!�v�m��s���F��YA�3\5G�=l:��i��t���1:��3�4��̵U�c\��~�;�ܼXz�_���YC�4fp�a<� t�>�H����A53�(�Qn�ul��xy�h`'c����W�_������u�{���,/G$]�31�b���������;�E*�
�.�喵�lZEb���0a`Ki��5-�} 1�0ʲ��].#�s\$��a��Y����ĭs1,�Yn)�f��7.J�v&�y	o��L��n�;6��6X��ǣS�N�Z�ٛ�~��C��z���y��LUa�+_H���I��o��m�8�И\ܡ��r���J�&od��Z�d��"�8��{��[Ð�\��ӯW��EB'ѕN*��M�,Ń{qr�T���"��f�T�-�̊�X�W5�8&�T��].e!���Ӧ�*�5m�7Kќ���f�Q�!f�uhOI�'��`�����LV/�e3���3+uȡ��y�v\���;�(�r,��Y�Qz3����F�QE���vuss�£��~���D�Q:��iW��8��$:� Ne�����ڱ����|m,���g3:p��iK��23���M�f]�]@T+[x
˼�;.dur�|�%��Ư����2��o{U9s꺘S�єɚf���3����^Ň�T�p�{;���U>��c�a�<�]5qf_N��Q@=�ө�X����o�
�^q�Vp֐��c5��$N�1���S��|!� l]��s���%]��J�WB�ĝ]�n�vd�n�K�R�tk��:�Vu��&�*�D�W'��"���=`<�ѡPǫ�љpd��]��t��:y�$���ZxT��f�of���YԻ�􏀨x�������v�F,�te��<�4j+F�5C qǦ��e�ZHrc���|M]Y���/c�W3p����\�B��n����ݙ*�:ᐅ�,><��f��2�x�@G��v��+ ��_%9�s
�
�:�M L�m<qX��J��tj�j��|b)��ǁ�9;�sl��*����_�m�����]q(
�n��[ܖ8��5��ö3Df���NVmRYv�1�
�7C���ѽM5��p��h\�ܿ�ΰ�������D���y���>����k*�@i,�	VC|�^S��iD���6�t�u�3�V!����
�vz�Q;�����JO>��ŶK���\7�dq�W;��s���Q��:A����7Vga|OE���^��+��Z�TsTtԘkU+�q������u��ZȺ�w|�O�=T�R�9����wc��{Z���*P�W�٫��p��>��]�m���'ð���V�S+]�"����3n�Xԯ��v�d]���u�tx�.Y�+#����|�\ãs)[ŏXT��D��~��8a�or���Ą��@f�՚�ۗ\cA�7���㷒5�2����ì��7n��
�4*�1�� FNՅ�n����n�q6V���)�'cU:_2ڮK'%�U���-ڍ�r�r*�ͥ����8��1�/qk���'��I�[5����õ.f�!7�6W<M�h)@�mv�d�1Ԯ�d�:ʲq��4s0��5>ił���6�"�RME"$����z�4�4�:`���T>B�� Z"�`�`��]8e#��0�!*M-�I���+J:��
�SNT,��y���y�{�o����!j$���6)h�U��9��}~?^�_����������������~��"�b*��*�����b�9��'UAZ*�9�_^�z��z���z�~��������������|ƎZ)c%%���Z
.gQ'�j�&yJJ"J�.c���\�:]44���M�#�4�FH�UM1-���4AK24EQE@W1�
 ���)��������)��y��1;��5��"$�`�8AA�����cRӭDQUE-���/v)j���h*/j�vq13IT�q1#y���>~m���.ci�j).Ұ.���1��HLJ��U.bHVT.�r8�	XCbf��i+��:����!����f'u+I��4��H&�nN���W��~����q�"&�-�����x���@wo�CF�[P���x�guO��Ή 2ex�y�����%���`1���7yWz�lT�H '��Ta`sY/6	`��}m'�a�d޻�L7<)t�9gə��t�m.�ȁ����]���m�r�����1��1IƸv�NAL�>'6�*�r��֠aƼ��7=��M�c��.vz�=��\=l�E����CoTx��hf�!�g�1�yͽ�b[ģ�ny����jΫ����^�dw	�=m�G'��jW�`�*�29ދ�oN��gHg�c���o�i��&�[���3���י����5���c�;��ù�6�#��M��z��n�S����}������)��� ��N���2/)v7C(i�@�`����`A�l�=@'@�G@
�{�N^בx0���-W�̤��J`�3r���J*��d;��ȇN�b�`RuL��M��"�b�m�p#'T�a��9d+���n��^f� ���e����od��>�͔�^�O��Lϓ�ɚ=O�c�΍��֫O)���m��g��M�5��z�UOl������U���E����E� �@~E��q.eF8��b�Cm�Ry�Ӧ:�_���M��{X���og)J
�Z�Ty:ۧE���%�2���0;�*�Cޗ��;��>[���[�^��uW0��m>�Ynq�U��ٷPkP�}ϗpi�r�����/f47���q�1�;�St2s�?��y�������򺬼�R�7K�|���&�ޱ��Ƶ�2�FW�����l>b$�S��,��m��k�E���zb�u���k]!���J���i��Ʀ�	�Q�n�%����*:.��[L��O���2+X��1���Uu�U�C�X>������WB"���y�aXe�Ǔ+o�,#K�|z��r�1ө����=F2�n�=��@��g�c4�p��=�8�-k�U_Gi��U��-.�+�7F�X�M�Oe�.�B�5ۓ��l�����[Y�!ߛL���z���Y��3����;x�[柭���Noυ�톗�v�}�QU��-�%��������<��m ��'�i��
��}ow��l�Fgf��-����w*:��v]���C�����ü�D4sq ��v�h8��{�M�z�J�I4������+T�V�!�\���i�)'O�F�Ƒ1�G<�s�<t��1��0�i�JW�H�����0�WS8���Q�Hy�vrA�ȻS���ϙ����k��- w8�c�O�.�)�ׂׄ?P������H �ru�i��n�񈗫aB���l3k�_-�	Tq�O��v�Tx`��(������F���(K�k����+`���#�l6�Z�xH��e�l�RPQ��i}�L�F�b��Q������L�}�KJB�;C;�r�Z`��ڃt!�R�����(S�W ow���'+�Vͅ�[o��)�Qq��[{�d���8]�͝�h�ʯ?��y������� y�+�|\���=lͭ��~��W��}|�H�{�{���-ė��OI��do��u�=�Қ��մ!�{%��2*\��v7���&���3��(J�-�S7��ɬu�Xc+VSC��Z��C��$�l��m�5y�rj�a`�1g|�q
�|s�å�E�ۘ��R٭y�7)�����a^\�[$
y�����}��z�PY���Ml��L�m�hö�R�l�\
�ΌC�\�C^�Y�@�[���|sU0�+c��w⪹L����j�͑-�-��y��S1��gm>�k���Ot�z9�>�a%kYC|���]�GkH�Ȁ(!�L#��M�o��1�G��#Yf�ާE)�ݩ���$�h���6�A��[�{�m�> <�B��y�7<��Ak���[Y#���yU��atM�k޵PC�-��aza���ف�$7� X�a�b}�`S�������/�3��z�yfd:B7*�p�kA������rm��Ӻ�t�6�;��Gپn�9/�<;��Bbǫc��j�zƜ��W�P�<Z�Hݮ9���Տ~t�c�E��pN�3�`.�2 ��`��& u���̧j�k�hjg��][.8n�%�v�. Tw���CA{�/�NS��FLyy���xd�4	�${773���2t����u,�sTs�ސٙӐ�s�L 1��}�,�h�]�4�*}��{��c��11W��q7Zi���x
�{�8��?�� ���ef�����P� Q�:�Lv�G�q�v�k:7��Cs{������I�p�]�R���0���:���ݭZ�c���[Jh��f1�55߻־�3�tqy�����4?Q}�㕅,]����c�S����(���M#o�@ڜH>�k�o�kd��i�l��sW���d�y�1��a#bS�Z[�{��!z���&ϊn.r�"�>�����m���q�5a�E�܏�Q9͑y�=�<`.��`�.*_[H<F���o����,a�p��Apzu�9�	�����z�&|НF�u0�>g�UK�Ӿ�}Z8�hf�%Ǟ������*�n�nɷ�õ������$zs�}�D���D��Y,|"�ӻϻ��l�-!��'�x�q���Q�Ys��͍��.:Z*\t{YE�@�Es�F�rʣ�E��Z�vs�S���U	5�[ӏ
���]��{N��FK�&��m�;F���Z�'��V�I�(�`+5nޛ��Iv �l壛sL�39�e��c� ���F](�{-���C�~�5�criLn6��μ���0cd�"�� ���^�~�\F�Ⱥ"��@P��C�0�h )vWs�W%늯t}�.����V֋��/I���.p(%�DwS�>h|�٠gT�RMu���Qn�مɄӌ���X���z�ޖ�;����ɢFuY�{o3ː�����n�<]ڂq�AQT��I�4i�=�UWy������?���'��JK��C͖���_N���=��?�[����r1���l�}&��ƫ��/<f6*mI�V)���nCČ�s��'�z�iB�䍟Bho��l�GM;�i��E�;]�4M�k3K��p����l�C���_��څ̯�?�s��8s=A'�\����a�� t�g�i�5l�;����zgc0<`���7M�xE2���(ׯ^m�e�t��t��nQ�
�z�$k��x?~� O��_�u��3sk'���@<�cH��e�BZu���dn��2��K&�+����N��v��Uls��;�լ��;}�����J6�tx�����iL��2��쥾p\�c��uͺZ[SeaޅMqW|zZ�l������Dy��Hb��f ��p[u�������d����/}��U^O�A�������S}��վTG����S @}z�@dyW��$��Z(x���V�7��l�:C�B}`�/��g�� oA6{�G����vl���Q6TQowvl[T��y�f<����Tg(}��8�/����}f@�d�_'pE9iS����d�1��4�b���e�eNNgm�;�F��~�N�1�CJ�?]d�|��x������]�)��^����������-5|�6<�1TE(���8�4�Bt�
��<C�lH$)l��a��u6+�vH)/S�"�k�����*���x<x��>�>.�����9�M����5O��z��6���ת;���_�@�ڞ]��՛���K�q��oj���Y������[>!��]	}��z�M��	:�������l��Ȝ�a/Q��Sʙ�ݵ�۶)L3�e,�w�8=�p�n0��]3�i1	���C��&p�1(��������W/
{�Wl^Z�k���#z �aUk%ȁV�qH�W��6���N��R����˨gL���Jd�^K�!���{:!ce��[�j�*�|Ԙ]ЭYFل��<��B+(q��S�J&�'��ޭ�j�<O���8%�>cH��
�y+m(�Į{��#���F�����g �'$S7f1��d�����w��$�C�����P��{�Dۣi8kބDلw�����9��-j�u�ӫ���>�?w(u��Ѱ~�;�[�p�s[E4%��}�:z[U)�+�tq]m����[��Y-�feM��:�g0P��,��z��)����ߓm	c��;�zMvC&�s��je����ڰ�����R��";1�3�;���� �-�!���3̱����w�_�U�e����6Z6������#-ʶ��ё�Mdŷ��������`��sN�p���Y)wl�
��1w7gQ5w�/��e�\ɏNWI����bz�bw�+Ɵ�ǅR���߲Q���آMG'�=��ww���$��5�4ƼDWG�f͛(�D�_l�$���.E��=?�nc��0��z/�#������ � �tC��a���>'��y����h���4d��d7lq��g��p�|czD9������u�2��T����'���������%
��$X6n�(��]�sK	��;�Y1ʧ�4���g-m���إ�E������C�}H�@^���L'я��؟Y���[�6�xލ��'��SSr)E֋y���;6
�i/,� vƀ���Ɵ��n��b^������Ʊ��5��ZHm��9�1��r�u�du���p�Ȧ`�7j\����qg7��<�[�>k�L@���:�S�S�_u{U��zZ��.�����W+�8ջ�j��\Y0*&��f�k��ü��;���:�g��j�i���������Fsy��k�
�	M�d򻡾�� 3��ؕ�_�T���m��A�k��U'���Uz��۴!�7ɫ��g3� v�qYa)���Zy9!+�"BG�w&�����v� �j�������K�EcH��ic����:�ȊJa�	M�J,�%5|�
�1���ɸ�W~3����QWg>=ӛ5o�_>6��w�8Ha�'�Ӄ�LG3]��F���}@�(ؤ	F{������]ݦ��s+���n���j"d�{��^<U.�Fo_��c�Fbk�rž/残5��������6l�E-��mvۅ�}��kz����do4�J��Ã�#[�qB�͚��Sa10̳a�k���^�WU��y�C�mF���dhG8b��q8{�;��8��8�)��	�:}#W@z=0
=OyµK]���kTR_��|����{8�h��p�����8��0�}"��w8�2��upkw�ވ�C��ŕ���=��<�ϧV=�p�Ë��`g��@�:}�h7�i�7q'q������4�E=�F������_��"v-_|#!��v3@��Ps1���Q{m����Դٖ�&���&M�
�뽟+���Wr�K?&�슛k�����p�u�f8�ۈ�nI��O|�mg�Z��u�%s�7v�͙�m��e��V3�����e���Vw߽����LI֐9_�w��_�K@�&��/�X�ۑ��Ӛ��]�{���!�vp v�s	�tӭ�Y/���7��{���k������c�[ʚ��v�5J�-�jmtN�,�䭤4��˻�ڀ�Y��Y��S&��:]I�}�O���.jnF��:��+��}��٫�����;��T���z�����ʼ�|yT�R�0�IZ���o;�x: 
V�6�H�?`��;���q.ޅ�k瘦|�ڸ��z�X� ��LeX��J賷����S�9�:�%b���Xyy�眦�75�x^y���J�x���>�?��<=�x �xy�guU�ZM��r����o���|�����'�N��I���CW�����p�>��k��H�m�!��e�T�SU���:�S�	5>��EK��Sw�2(�^����s��&Nr���a�z^�MM4,��82x�L�r�h�a:���6F��i��֫O)���Gt�7,!�5��"�ݘ液����
�b�|_�3�M��A�J{"��a>ׅ+ i�̆��p�BX���~�ֿhs�>?>pV�ň��L���Ǡ?9M��3�޸&9,,�ca,�q�:�;J�p���ݱI��K���5r|����K�	�4���|����ιK��v�^�c���[�3&����]�ͯ��u��\�bl�2��kn�驉V&����G�P�WO�&�N ����i��U�F�]W[t8Ō(�k�5�;�a��$��1u�CT�k�6�B{zM CD{]sX�����;z��a��[@
�=S���;���ʝ���[Ss9o!a�6G��8.[��ת\b�8CBf�y��؎L2���ۢ;���A�.r��KL/�zb˓x��[�͔#Y���w`O4F���S��|%���S��5�;o�����z�P�_C�~T�h�޵s�s���5_��q�ܻ��a�vlR� �dmb�7��	���:����8�oMt�71�k7QW.�͛6{�{����S�Rf/=��st�16Am�cj�����3-[ƭ�u7�.ӽy<4�Ǐm=.L#��Q�%=~i�18����;'Zڏ�� "���Al�B�\{[g1�v�D�z��v�FV��f�w@�cÕB3�w��Z��4��'+bp���ӕ��O������v.FT�x�m��������k��y�ڠ]T�\���1&�MW:�s�EPװ�����9:'ڠA��%��f�ol��&���C/��]��õ6�z����^w����%���%
����Ί���L͊�b|�4���vm�R]фAV��:]�Ͳf��ކ׃2��E\��,������f8-�MA��iRs��I���#ܢ��Z��#-����|�%��v�,!7 M�ۜ��ˏ�v���&�|7�;��J<��T+E+�����1�c�Nת,�6�Wا
����b��vä>�ε���G�^J���Q�]t2�gNd� ���W�ѭ&1t����8h��(~칀�؞)jR�)�uDR�'"x�]�;����q��t������cU�m�i��\Ү`l��e7g�B�K�M ��cs-VJg&q�V������=�"�Jm��5	r�Id��:�d�����ӱ}mN�����$�1�v����l!wɆoh��z��9@��Zǃ�\85CS��oc�wQ㘎�B����-�fnY��Cn*ZӜ(W���¨��vB{=�wd��QR�C��IT��\�&T�E1���G8��+횠R��[��͓Z��m�;4�w���X����57p9��P�Z/��A�aokS��5*o��Zy��+�Ԣ��8*����S���(�sݦ��*ܬ`�mܧԎ�I`��JY�uW=��:jGf�;�<�eX�'Y���6��`��\�Y��t����J�^��BI�-�����
�e�1�$+����\��E���
�ܫu����7�&������.#e�O��a�^[��"&��f:0�/yX35������b�+9vg&+��M���W0�> �kvSj�x��yP��+2\O\�4�qS�N;:�t�k�u*̥�7u����SS��wP�N��QtXe'%,�f�L��;(�X��an������!�۬U���Gsf]N�qL}D[[����M�����D�qǤ4��\�N�ԃ1�ł��t��ȥ� 5ItZ�21,�S�M�����7�IP��~/�~Z�y.{�GW{�Ĺ��d�����9�kTZ u�v�B@Z�����Jh9�d\��4�E�����M��J�C��h��bsQ��J�͠��'rk��A�eV#4�;�5��Ov�����L�D��׶Pa��n���8K�,�QӃ`�u�(9����&�Y��[u-'��_Q�Z�w��V�R+��v�a�u-��oWw)8�㫻#,n�]\��k��V�W7���o'1ly�b��|[�/��ü)���`B��/��S�L)HQB��U��|��i����e��.���ۼ�❌���˒g)Z�����δ5,tW���(#��j�-�Ȼ��t�Ky�e.lD�WlcEs�+4�荻�ġ���1IN����c�1>vJO��׎�M����K�G����!hN/�s�e��Ŵ�F��*��]�����õ"����Ï�YQF�\������uN�x�n 7x��㬸[�ޜ�Y�;1
Y���wMΩO���=Fdr�{��T:.M��E78$9T�6VKy.�6�'�J�Z���t��;�O�e{�;F��H-�)c$�Y1ܢ���;޳��F&�P�1{xʖ�Fjqc͈�3Ç/9�???�=���f��������vח8f
g0ED�A��������~�_ǯ^��ׯ���}}}~�_��֤�/��RUkP�LS��)���EW/����ׯ^��z�^��_��������:�E4W��@b�"�6�s�TEU4�D�D�T�P��+�ֱV�*���9�Urű�e�("�"18/�1A��(�(��=�UT{8�-�[V�l�*-�QDLUQUlb
���ESh5DZ5UA夂+����(��������"���X������+��EVƩ�

o�嘂�����٨" ��!�lU\�s4$QDD�5E3s��#AAOK71����j""��y~{��S�W]�|�&!�v(�J��I�WK�Z�{�#�ۊ�r�n���*Ur?���Ft����6M]L�s"��~����x��x��)߿?�������<{G��j3�9�Rl����} ���DN���j�t�9@^�3�@1�
acdL�
.flε�����!�Yb��=ޚֿ3�LZMT8��-�4E.���,6�	-�N��=5mF�3;.1�ս3�]oG��ك=0$��{;�;���B_��H���,&��ZX6�7I�m����͜»�HKF����8�崂H	���C�'�i+��ϣ��DC�̡���e%�Ϳ�+�J�%��ܭ�Ot67���O17�9�8���"^�*t��5T��HM���(�œY�|��;�H�/�����s��	�hv��9��7��˪ź3{svorm��,�l0W�`�X4�����U|w\Y05T�z��u��Oّ�Ob��kr��7>9!��9�E?&�[��$Yl�����z��v���:��$�3݉���{K�%�Ŀ��S"-۹*�+�X+��X�������=F�]˔���5;�M��R݊fީr/�s���AddǞ�#"i����tKw�"�x�.'_���-{���0��V�xL݇\gU��8���U���3{՗�mmo��n�=�� ���(֔�0 
BK꼡7�$���^�*����ˊʛ����v������s��{#X��%kꋫ�Mu��U�տG�x�x�∡���Ͽ����9�?�^������T�v��m#�S�:�+f�ݬ�5L*=�@EX[���V <�R4���nt�1�`y��+5���+�
�Jl�'��
��,�ĭhf�gN%og�n:�;gq��X�|���T7sT�\"��O�����؄V%S{_�i��UE�{�pU��Z�i�"���2/���4x�u@��ƛm�d������ȍ&ݴ��N�؞�f��U4����M�8��%�fᰉ1@��D����V��p��P��n`��@���8�k���}/5�ӭ%���c9�	��q�>�>�ɰ��m���zS����7�C �Z.v��9�;���6��f7&��9���\x���3<i̎lc9kg���o��z��Lg9Õ��0dm��O)>�����ya�:���vY��=��ٱqx����΀��d\���=��7w(�G8kɵ*��f=���׸/�����A>�����(���w��YB�?����m1���4��3����/�~�����:��N�M�(����u2-�ǩĭf�_�$a�6閲���vrW�7��P��j����e%~M�5Ƹ$G��X*�o��Ճu�
�*��!*���i�U"��Kn]R����Y�w[>�3x>�jI;gtdۨ�Ẻc���r�'���FN�AU�{�s�/G�uy�mn��VU�4M�#��弭���PO��x(���<��M0������Ē0�a�9�}���1:�ˢ#�����>Q|Ս���qH�:�כMs�r!�4ק���Ze5��r�����J3�w�\���,M�<ዺ���.O����O�#�Hn0ԔmS�嵙�_)��]��vxr���{����$s�:iֆl0�~�h �k9�	ч���Mᅅ�)�ƩT�[C�}@���2�Z��D�2�����*0=���N�8�Ɵ58�|��u���mNQ��n�Q�y"�W<z�k��l	<[N+�>�[�p�4�M~!q#+�:�sc���?���J^P_�&\v1�q G(V��d���9^K$K@8�MB7��GU����ݜ�`v�|�nLT�!԰�\"���k¶���ƑI�6j�ǛsSԮ��ݩ��B� ;b��ҍǑ f=��a�&�?(c�A��Ez��eb��-�Xb��Mn�2���C� Rzn�	D�T/m�9����v?�j!�g^RY��O��CP�J/9��� `�oӭzP���>�q���s���@�r��c�@s{��C��~���H�S��ݭ��г�"�I��#�i���d���V��C�M!�WVJL�X�*Mƈ'F��,%��������O�ϒ����}�j�L�+�������]K��	͝�NG��w=�j�c���S�k-���������=~?��W�<����ռ+���O����Ǐ��`V(7f�o%��>�K�|�ٱ�ȳUwM�a.{ge��4�-۹ڄ!C>kL7�p#Z'�iۘ�i��E	tq]m�>"��9M����y����FV�ě��D��_�sH��W�"�T�B��4�i�x�>�Yv͝1��y6L�ٶ>Xv����xhcl��z&<m�r�ͅ��k������3#y�5����w���6��4d�Zg�n|Y�
fΦ�m7�A���ۂ���=�H��4�"��)i]ɩ5䃘�Z�� �}�B�Q��ͤg;ǅ/�Ua�|~"��P�hY,�?[6H�hǟecg3C��'�����1r��|���8�;�tӭ���q��+P�,��Vc����x��D<=MV�,K�a"���ix=��`���0��V���ci�6�������f���,_~1�f�J���"�X��y��@��@�w3��N�7��'������1Y��p�ȟ�����R��m��-$8��
�=�p)ڲZź���X�f��t��:u�!����p*�1����W�L�v�gc�����2Z�r��6�S9�7�����f��Z(��6�V`r�j��-v-T��ù�x���w`�F��Y�X����\�����3�pDyJ�#f��*�^���V����7��yǼ ?�� ��jj�y'W�
�uuH��碘��Y�m/��~>~+�H���p�v��ᒢ[f��N�=���֫��^�r2yE�y��Ų�G��s�pW�U��Ug�w��y�Z�׏M�Y9��JbqtiF>��w�ׂy7��o^*�YU�\=��kfM0=��a�en��h}��2���r��	�W��gv����V������e軇Vo���8���r隰!_�3&l.5�r��l��/Gt�4�B#x���mn�Gh-�6�[(��f�Q7�m=*�f�β�j��`!���(�_�"���xǂ���.�����a�*4���-�;͉�vsTi��}>�Zz�t"#ݯG�cp�(�,Zi�%����r�}*OЫ����Yk):t;��l��C���y>���q��`;�m!����4�>&W�1�X��!ma=�݆[�O����s㸟��[{��~n$�g]��5������&�~�TG8j+'�x�҆03S	�����������s��6M�V�؆�d�n��11�T�z���3�I,�E�e�=ӟ���R54ޅwv:L�� oޭo�$�2oϭf7[�y*ë��a@e{V������B�k���+q��5�U�L����xNַn��h�BXz#55WuЛy&��|�ܫ{Tn"p�������}�� ���������UF:o�]@����a�5��Q�����M�����٬(��S��K�[�"�A����{��k2.�S9je!���(����rl�6���Ø�7&�<�튰��[��y��R������b4?S��
��aq��E��#�ߗ��k&+�O*�J����&�H�kf+�kF(�6K.N��Z \b�f�R�@�p�KO�M������F�瓃EL��U�9ì��D�E��#x�mX���z�v���g0%�ې���.ߢ�Nl���7*�sk�P���cE�4���A(���U"mfK;Ty��i�Ct��R���z�ͻ��Yl�5�0��s2��k�Gz��Q�J �n�L"�қ�"��\K��?n�Ne%���=G�+���UǘqcE�����O�Ӯ�̈Jǉq��JX�O���2�v�S�2�l_y��j<D��QG(b >�G&�"���P���/t���Lw�i(�x}8�� ���j�N�(X�kМ1~��g�a�	{\.�~\��-u�	��EsS�g�Ӈw:����[��o��Vz�)mΤ���� ;��vT-c~�V/9���]]�B�jx�R�߰R�B�J��hL;�9}�to��4�/���Uk����v�F����*��S���V�`��,�k0�oR��wf���w@���tC'T�RR��=�x�~?���ǏU8y~�9������o���I$���ߵ,���Ju5y��k,��#u���6�5�� ���%�H2��El���uU�p5-��rz=J[�F��'O)>�X�h��f�L�xX`5z*q�I5;0�Nc�� ��L�4.#=`��O{gي��4���|�d�K�޽�{��k� ��#��!���*��9�ÙKX��|�m)��	�\^���*骢aOλ���d�h����U�/*U����3�bm�O�C��8�	�͞V\^�l8M���ۘMW�T����uݶ���W4��A5ݎqbp��'[i���r{$�շ�oa0�����M��;�Q}#`�@�8@�(�	��k����h��3 7��̟��QB�ѽ�&�32-(-,T��iz�b�}��u:'z	`r�ţUK��N,g��ݩ���=��+/��p}NXCKCv��qƦ��P�q>��<���d�D��b�b jzwz��v��/�
:�ݛ�,�l�v��	H5"��8��*\!̥���k�
6�DŚ�ؗ\B�A��a7����ܩ�����BJ�y��Pl�A-7ʲ�U�Z�},g�@�&�+4�K@Ӑ����{���^t-Z]x
�z�3!�9�/�d`�S/����X�ڌ�cdD�ޜ/2���N����>T������s���W����}����Ǽ �[WS�}屈����ܧ��n��t�fx	�}���F@����i�����"�c�r:���o�n��d�����fK����s���6����h��'E6��*,�uۥ����7A�%���&���.x�X�̎oR+$R�#�z�����j!�9��)��;�6��.1f��]��'bxb��L��A�9k�s��-)bW\��G\���K�*��l�M��1��o����Q�g<e����������붭�?��c��(��y��3�XƬx�,��'���W �z�����Z>�U�F�
�L澻?�ӯ�AwG����'�#�Қ&.�w�687�Ri�� J�!wYU�ox(~bh�)Om%�����>L]흜��M~Uٻ]�b�Z���쭷j-�,�f��$�8,[�ir-s�ф��C�@�9�z����&���!�Ye0�ށG�=��ü�_���'�����5�����߃�j'S������թ��/�ù��/ݏ����'��!��qط@���0s~�/~��Ŏ`ZC淺Q9�rF�s���*4\V���w��p3����ƾ��]�F��qY���^N���ܺG� /Ʋ� {Y*�b�
��r��Ce�5���<���gz�oV��r\,3z�p���l��?~y��;�|�=󟿿����*x�� ?"o0�,�W������e4�ɺO��賕�g�f��U��4�|�]4�C6p���5��uĭ�}�BI�p�τ/<=�V;��&r�x��țl��ךy,��g.���f~�.��mݽygL͔�5��|yf�	���4�]��5N6)C�tT4�t$t�Ȉ� �Z[2�g:�e���/���m�5s�V������H���>Q2��V�i�H{˥E���P���i`�v��&��R$�D��6]�Q��g�o@փ0��-Ȭ�pdRml�E�n�V�އ����m+E��m�W#4�L&}֘eAx�kdx�>Kѵ9�6��+6�7n�u�ܰ@s"g�Λ�P#6���O�+�H�h�Y"u\\4�[4��3��w�Nb������{Q�C�+d\�s�\Z~Ƒ�����V�&�tB�g�L�U�L�������ѯ"��i�ʢ`C������6ȿ��G����i���7L-j�Zky�@�J�3�D�aQ��
̠�3MW�gT�|A��W�g����x�aK�G��:�+��}A\���_>�L?f���]��������c��Y�ji(W����n��;��o��i(st�ɜc/jL���';iVv�m�P�ls��� �1�.sgv>����e�����of6�5�=��ؖ�#���g���?���xI�� ǉY�
�t.5q%��u��D,z8t�$I!5ۘ�a.�ɺ�zc� ���ױ���p��օ/u�WK
�|M!'�at�q�Q�F�+H�x�I��g�97"GT|­���sp�7�K���Y�V2���>B#���ʆ_�Q�o#��4�@�cy�4�sc��;z3��Ƽ�[Y�-x�l!ƕ<7qц[S	�!�ԁ�^�}0#zD9���줸e�U��Sp'9�v7^x�<��3����/��_g��fk3�Ӡ�����n�G[:��{�eF;,('�.מg/����	8y�|�j��~L[���𗞻��ۜ7�uM��7����A�=�d cz(�nvlk�lSi�q*<%�M�|�8H�߽�~�����m��uz��?}�t�ڢ��r�r(d;��n�e>ba��7$+�S�ɮQٵ7���C^M��Ah:/���EҨ�m�ˎ���i{�~J�$z̪J�}����9�̽��U��ac���)D���z1x��H�ؒ��� � r��T�r�x'�G�8���{kR�ϭ�n�8R4���u7�.��:(����׺u�s����n+�[�bɖ{St(���&vKڵ�rM�f��fU��9u;+		�!�� ��F&.坙����7fC7*��4{�(�d绁�h�gLYȒ��uΗΕ8��5 d�xΈ黆��KsS��p��]sjL�k�+�u�b�/ }�b�(>����q'��1r�yVqu��F�Q;���U(N�w���ɇ5eue�k�B��s��������vЛ�f�r�B��#/@�_t�0U��Vf��̧D�jcE��S�9�ݑ��5��P���tW"|���W�A9����c�ץ�#<>�j~���o�����G �Z�J|N�#�T�x�J;:�Z:��c�2�?�(Y�����;��6o[.���2ʠʑ���n�C�Kqf,-z.;O���v���n�=�0S�Jw���̈tU���ٱ��9��fX0.7&�!3�@՘r�����V��[�Ϻ �,Y�+��7�]Y��R3.�Z9%��WqQ��ي�8wj���;��+f�y6�Y������5Su��U�gp�$�\Ġ��f�pռ5ChQ�⮴뺸�
��$�J-,4*�[�,#��ʱ��)����meҸk��L�!�2�ƆӔ��tLEo�v�֧�ݰ�U�3䲉����5:�j�ާ�ΚY�B��U�
�bdl��U�\t�� jڧI��WK���d�R9x�(d9�e��A�%W����p�CU�R;�*�Zj�`��Q�1�ti0=f;���� �TE�
�ݙ�[ɉ�w}�f�QtN�gi=���{��{C��+�=S�U�M����榷��=�M��n�L��Zk�8������t���¡�̵B4R���M �\ �2ZT�}�a.��\�Zֲ��f�O,�^��b��m�訩`T�bk*q�\��[�z!aۍ��]��ظ<`�yg�I�q�o�͐�-ܻ�W�ce �j�x��Tx�W˵��
��5YCQ�c"����&;-f>4�`
�a��GP�G����sO�qު.�3 �|���:.B��M�\RVe=�Z$>��i��H��X��%�^Z���o�}��)v��{�kS��[�� �'(Ƹ3�z��u�'���\9�x�a�r��/xQ��58*ҥ�t�l�pB�7%�}O�Tl>:�Tᙃg�VM�yY,Uɥt7\�.�op��v����T6��s���3K�y�]B�i��^�ܣ�0����+"�r9ˍb����w��y��E��� ��q����0E]��g�f���W�����Ɔe�ڝ,���� �8zq�	֎LȖ�\o6�[�r)��wx��oU��'��7�n��,ޒ����qM�����@ּ,�~B���7L��%�͝���p�\0y/2Y�D�I�����p�h�e�(�RB���A� F���(��A� Hx�ˤ��"�b@�F�4�-Pb9J]� ��L0�/�{{�J� ��BMl����[j�uV�3DQ�s������������=z�������������4ߣ���Q�ETET�1QEUSATQ-G6&"���)��������ׯ_^�z��ׯ��������~�;�o�ATQ4CUQETE��>aē5Em�����)�*�b�����`����"*)��t	����R[��`�4EP��:�����h��*���*����Ѩ**��(|٩9�U�PU)1DLP�i�SDD�Q�D��4UO��;f� ���*bJ�	���KUTUEUs<�%D�SE�SUDID�3EUIQkE[��*�`���Q�c�("g�ꪊ�Nl�乊��*�����������$��&`����b�&&����
"
(�Z�������h"��b�����
+�ƨ �@�B����U�0���M%C��w�U�̚v�iB�B\�ռ�P���a��1�&���hIb)˳*R-��cn��|^>��%�	6�X���Vl�v*Ql�f���ީ���q<x�R!R����Ͽ�^�z_��3�L�~fMۍR�qy��sǬ������*��P�y8�}���'�mlVP�n�ǻ�l�\�{%�"�����ک��v����̈k�p.�k*7osy��޲a�At���g;z,ܶ;,&ǚc�1��S�_ջ���Z]Rm]����ѲYn�<۬�s�k4;�=������� ���''ş���a�F������+뛽�[l�Ə.R��U��&^J54����P`f4��t�W܉+����?�?r��;�K?ǃ�%���z:3'F�!w¶� �� ��[0gm�t��N�{t�ՙ�r1�7��ڭ[t�1-��}��B�W��O��!�2/~h8[5���r���s:�7>c;υ�@ƹS���G)�}�a�&(b��PLPu�M�@����Y������Q�٦��rI�BH2����Mù1�B�1#����͆t1�vbm�>���8�=�M���j;��?r�V�<�͍��]	6y�����!�+�y�Ar#�!�D���C7x����0�O���[	�-R��,Â��c�?+kG�U�v���f����QNG�/h�C��4�&_Z	/�����ٱ���� *`0f84i�I�[Dɚ�-qR;��/"!ŗ��SpG�pwp�X�g���,�w��j�x�VoX������l�9���Wz���U//?�� ���:�n�2&��j|�v��C4�G7�����o�t\:i�43i%��Zg/�������Xْ��)(<<�T.<���ؾ_t��j�#�6�Ao��\�5����ff���W�Ww�ӹ}F3����Lqy��}��~�?^mz��9(�u�Q��������5�4$+Lk�ww�ӌ��E���&C�	5>���Ï$�n�Ž\�Q��$d\*�Ȼ�;�:r�)�i�� ^Ż8\h{�T���gL��R'����?��lk:�7����wn���סf�Ky��$󭶜A��lަ�f*�ج��v >�dd=Cw�yc ��0e��?���K0b#���ڎv���I��o)�0Ϋ������-F<o�n,c͙����OL�u�WoM��(�R�&1��Xǃ�3��W9��y���c�_d�u@��F㎑���<m���[�������g:)���kS�ݘZ�`%�Y�4�$���P���έcn�'4̝�y�0�v�ƕRι����v�I����i���?c �gK
&݉����f/"�������������o�VDf��ל�+����.����Õz]mnX�0�S�3�y){j#�U`gώ�mkJ�^�y����r�a��p��j�t��7O�:3����t�`ɟq��o���d:�"��A��&�.��w���U@///*�����3��c��{h��9�%٬��d٭�CBe�M��"�ۚ�Hؘ���&Z]���ja�f��C&��k �G�'ӞV�E��`&����Ǐ����48��^�Su�U�S[銢��tCF�|C+_���rn�e����Y��և�zظ_��(h4H��!Q�ʦ�1{ֹ�~˾n�G%����od�����Z@�}#9�y����>��bs��-���P�g����z��5}�ȉ$���.S8+|ǪA��9��Ob����<�V}�s׾%Y?~:u��H����w�j�~�$��Z?�I��
(���>e�h/q�RdM��n$q��0�rO����^v��|v�~dM�-o�߭�oK�+ʕ^_��.��QV���F7�C�V�$�:=,�o7��܂�At7!ְ�viދv6�ۥ�lu@��ϕ!��0U��~I�W����&��:�7��s o�ס|����H��b�"M�I�[@ط@���G���?��?+���Oc�-p���(�i�օ����Qv¨Z��"Fc�Q�g�ϯ���*��:� 6�	���*bDe�}�rh��S���;�����Qǯ�ӼDo3s%X���<)1A5� *F�2)K���Vm�I�ʕ҃��bv��{�aQ���e�N�$b�R�1$�����չ;�U�Z�Z(J�վ~>^��������H�v�gT.�2(j��|!����D��Y�p�\^lBM��/�|�V>՚��6ڎ=_ �2.�<��U��5�/�ߝ���y=�v��l8��kL����璱��P=�s�0�m�b�M�n����W�YT6~5ῒ���櫙�ڏ{h+[E2/[�5�7f8�6��'5S���UJ[{ZԴ��\�N�� ���lk��;��,�T8G5�[G4R�	��3�b�U��~���N�@�u��T���ˡy�����BƓ�ƶ1g�0�Bgh�������V�v�y�5-yT�v�/R������[K���K&�Ⱦ��f�O�@Xj+�լLl�3�`V:���=�𼒰l�J���'��̄4q��3*i�t[�	���,�ib	�эl� �cS�\��͖QU\{��?���-�~��~W��:����fˍ|�L(v�i�����k<É�yq��M�l�����Y�s��|��c�Rq/������A_/�ۄҷ�]avgr�;��
����n�[ �ʜ<��ڱ���f��=�!E�	o���`�<��o��DP��0af�}S�ï�P�b[�"�𵸍���T��QHQ؛#�T�R4��\���t���h\�OH�^�1Q���qR��
�::�cv*�Nȟf)�h����ﮜ���{�tv�v<�)� u"��nu��ju�5�m6ڝ̾e9O���о������6���K=��<x�	"�.��wg�EUY,�V�Q�;���;  �J�墂�~P^��ΔM�T%��8����Up�]����K�a�9��{Բ�C�S�s {=� T�4��CUˑ�ǵ��(�٪r�Gtga/��u�n�Y���F�^���)؈"=6�"���]
�۷���F��QzZ��{h�����3Wnc�4R���ᙉgka�6z�=�tQ�x��Ms�G�^J,�$r����i�:(�f�w_"�ყ���M�f�bD��7�q��%�8�ﷻw֧{2��et+�ݢ��ݽlS;��Ti�6E����jݺ\�9���@F1�K Eb��-�9�I�y�v]��6���t���rk�ʝ���A�;MQ�dߧb�[`:�I�_�1��m>�ʆ�8���ɍW����~����h$�v}�6�L�k�� ��<}�����v�r�C^s��m��d�-g* ��>��%"7�\�j�J��2ۓQ������ύ���E�"w���3�3.'�P�D326���9�� �Kf��KBz򷳝�o�yY����߫+�#g��w��b��54m�6��#O7c������Q�Q=�Җ�g.�Ӵ��U�Y���Ы�dt����ˉr��^�=W�-^4C���s�<�U���c�v�n=�x����7��Ua�|u�`IL��N�{��㝻q�-��q�<����R��~��x;���p>'s�p��6z>g���������CA�ׯ�1*~��j|�}.ܵM���>3U��3X�(,3c�g�;�.6AN��Ci�i�S5c�5���֥kw4@�m��h���!FK�i^]p�'��ڂͦE�r�౷)�v��$	�m�������B}�渕-c8ێ6q�u��'��\�� ���o���۔�*}7�m��b�u��a4à��I��W^���d�u�q����(�c�#���N�˳��Y��2.��l��Y�w3s��^��`<=V�㞪v9z���N�>>���,�䭤4��dɌ�8�A�&�D�.h�ܕ����x��&������Y�P9��^�(+]}������8�x7��M��c��Wz>	m����i'�4Q�3���ks��MH���#Y�E8t�Q�v��k�n���KD)۵�r�͙�k˲oƨ:�vs�On�j<z��X���	�4�ƺ:��r렲�$��: ���s����C�ڵ=L�Ԛ �j��0��f+s����s������V�al��Sp����o�qޙ����ЧC��I{Y�krJJ�²ј�q�g$z(�ھk.����
�.�^��L���5VNe�X��`���Hun�x��p��Eu�Ӽ%�2+�� ����\�q�*�ogN��_����~?� �J�V�f�����/�u����)X�9:;�-H��Jl�3���p����Y�Z�+�Kv�GL\k>��X�Z��/|�3\����(�mu�#(u�����3�/k&�#��l����:o��P'vǫݘ�.w��?���N��B���+/1Nl�7�f;qa���H�~֟C#�"�F��� Z�Gk�������9�tD�S=��s'snZ���wb7-�����L�a�S5i$���S��l�+�3���uP�qY�'/p��/5׻uv�VE!�niW���C�4��v���M�X~�a0u�s���0��,��:�O+��)�S,��>���]%�(����y��7|E
� `�V�#y:<>K��TWm^E�)>�	�Zm�S�vũ`k�e
�s�4����y�9�C�i'90w�98ﺫ0�<��W�>sO��_���nM�����鳠�7y��h:���vfۭɈ��s���br��Z�˶D�lPj`�M;�ߌ���n��{���|��$��w�ԯ����V��1��\z�\��JMͺ� �'�]caS���X�>�6J*��c�Typ̳\iT���u���E�뽵.�q�]�u)!�&`��*���hI�ӈU���q���-+49�J%��>��%w���|��o7����H	��f����Br~� �v�o�tf�T���J��񰡦'�]j��TG�@��kV����TTvCP`�N'��x�����c�|���V�+����QZ�yp6�̜��
������|��l;ms���H�>��p�2-b�+�����P����Ct��3$���'��s�h:3�FFc���/�SmZ�#�]�����@�v8��Q}T˶�r��s3:O��z,V�x�OGy���f�*�|ģʽ�6��iUQ��X�Q�^�qW����fc�O@��2��u�@�`Neb������BO%km����1���I���\/JU���G�cH�l�5��EcH��V��d\UwHi��-�\�';Q�5�n��9�0��2*���O�c�u��NK�4�a��^v�`��g���)�nj4_�)�L��Ag�7���Y>=��{Pn�"ǣ�N4���4� �48v}����0af!t�P��M�K���*������d��Ϙ��?�F�Ŷ@"��!T�+b:-�_/���x�H9�ƣ�g������l��6�.������͈��S�n�oV��Ͳ�YZ&=��t�|4y":@�h,$��I����h��1ǜ�5�Kv'�>�_U����9ڑ�g3�0ιM�+�ﯮ��ݲ���p��fSU��=LP��K���W���%��q��$�@�1�˳���!4/�h�2��ͫ��|��,|<�2�*����+�����Iv�;��N��������e�S,�7qq�����"Y���(ې��(�;����F���s��04��)���jv�C�����kF438C�>5�9)�����`�ټwo�3mϳ�6r�Qd�œ��_���6�/JE�~�C�x���Jۓp�6�R�yj�Y���R�b�IJ/)�ֻ�����l�#��&��lc��6�`�N%�3�6W��UR��[`�{�Z�*�1�dy�k m���)�`�5T���o�9�Tr�á��/U�0θXuye��i���]Do�"����v@J�M��0"����Z��H��V�"�u�*f�L�([��>s	����iL�M΃�\�UbSg٘4q$���H����gV��`D3x�I�(ZT}���LOkC5SC4�0퉏�Tec��5���wE^k[�o�/}x��z�.�)i�dA��������j��4)�#E���)JNX�t��R�g����#�/�p��~Sv�ZO'w^�9���
�bPvfC�L��9��Pڦ\�=W]�g5�{*��t���R�g2�_�8��^R	�|	x]l΂eKf��2�gvZD�
�-�]�9M*��0�s 3�^�}�ٻ9{i�Ln4��}>@7��=� �@#�/��Y���xM�P���Q'e9��߻b��H�f<Z��؊���٭\�sW�6NJEy���Fa-�5��1��PI��'�,w;	���?�nz$�ۀ�!gE]�h��.�½�5*�cO�ի�<�)�j{����#90�<�g:͎�R�l�(EԿb��1l�Z-Y�㠷n��;���c�v��ж�I��ǰ�'g7yF���4�7�����J����8�]�@nm��!�Y.p��/f�btoo�K#�J�<Ŀ֦����ݻ��q��|�f����P��*�������3�>3�qj����"e�S]w�����m>k��b���,��~���^�W�?v�	���F�H��d�D;Z� '�k��hu�,��w���mQ�:�K޸���da�w�i��!�+���pbA�,k�R�N�8����˸��9�f���p�?+�{$��w#�y�#Ao�p�Ó�0�s�:�=if��Z�dh�>Ȝ�Rog1�E�3�^H�"^^�uz�ѭķ�����N��Nk�	�%�7��m1�ݎũ�=6��w�s�DrXt)y��Q��dK��9ܹl��b5�ē�gb�K�]F#�5��]�k.`����v���fP"�Y�E���ͻwr=}�;L_���o7݀P��d�p\� ��<�|�d������R~/`�P�ҲSz������EKeAb��R�7�ٮ���;޺=���S4E_d��SA����Y�.��׌��y�{�=���[�v���yc*���z�qJ�6d�־OҘ3`�{'lRWb4r,g�U�o)Zn�R49KS�S跭�����6�b����#]��1&7��J�Pv��b���7�#S�`�߅�r���@�9ս[��[��Z�C�9ź����@A��+S���:��F�{�2d�涖��. ��2���m�|mG��_1�Q��=Wv�<�.t��5�����ga{Z>lgdq:.�L�A渾�:a�3\ 5ρ����[�2��Q]%�㜌���<�U�Sv��+���4[0s���p���^�ݤ�R�hu)ך5Sv�ƿ�<��MA�vpn��� {D���R�7G�+dn�F��o�Q1�s��Xyx7o/9@�c9-6I��.l&.��r��\�*��"���E]�7֋��۬�B��G�f��y�<�Xt�m�0vP��}f�m�
ZM���(��P.Z��n���9jٵ���>��ѓ2�s�6p�TZ�K0��dd�AV����u�X��縌7%��K�*Ʒ��ޕB�9c�܈y�I�U��3�GK�;�������O>���^{�),�s쩖J쉫�t|3�c���r^nN����
���v��&b�aZ�e�ϊ�y6�K��Wv��[V�}:ᙂ��n������W,��`��.��Xr�m�*�5�Į�uqL�0Ռa���7�EI�ӡ���K	�Cu �����B�_qyoX�wT��S3���GT��XT�m�t6�@a��Z��+w�����.d�H�*�e������A��v��@�]�J�b��[��Q�W=�.��έ���.6zwiڛ�һ">�Rwk�C������{IdWw����zT��;Zoq�.�C���u:H(�_��X�Nend섻�H>�D��ڳ��R���;�w%V���גt}A�l�[��|غy��t����;��/+����^kPa�����<��w2qJ�zĩ�	:�Z/d���CVC`�ᾐ�ѡ+l:����9ٖ�J��6����+d�6����,�lui����)ӯ����->��C��t�,��[hb��^���Ů��&f�ڸ��{�����W����gK��RƓY���oq�X�`tv�r�s���&=�gmp̍q�'��MX��l�ˢ�W
�r�Ӭ�v�s��cn:@]�ƾ�Mp�
X���Y�b"j�*����(�6$�"�JH�)bJ���������������ׯ�}}}~���_�ףڈ�)��J"�����f����
/6�&*ifN�QQ)ST�y+��%F>�ϯ���^��=z��ǯ____�������֪�i
Ӊ�"������J��
 ��"���CAILkQ�ib�f��� �hZ(�����"��"(��*`��f"!��ZJ�j��b^lST�14��D@Q0RP�,@QT�rqHU�h�*���T��@QM����U/��T�;f%����������e��Bj&�**hb���QL0AZ��T�%�DQD�RL���RUDMPR��CP�bh���Jh/�^��
jf�s�*jr΅�Z)"R	(f�"�J����y�M%͢ ��&��
*���"*�f������?7�~�~~|��>�=�sm٪#��nmr��T�8/2TΣq��ޛ/z��S���_�׈?�������3؂�Z��ߛ�LM�*��F�@�X��|w�v�n�o���{9�3�tO4l[|�[�-l���7[�V�����ݯ��g���Gߕ3.�rg5)qI�66 ��"ʊ���-xw�rQ'N*w7ʠG �7�!��"V� Q�=P!�a��p���'RzQh=JXלf�LZ�[m�w?��<��N �w)�k�'^�u�x�od��ܞMqj��ƻ��Tӏ	���z#�^�w�Sl����,V8XHgP��$��R+$R�#�Փ����jP��Ç}ΗʫK��)a2Lz���ou��~��Kť8hrj��	�hJF�]4D�ͻ�m��E���eR��9^�VH/d?��kL7�3�bwa�Mj� l:��<�Y�{������[��[.�wB/�.�V�(I|ffSY\-ƃ����t��F4Rq+_a�8�F\И����{�q��ws�:�AYy78���٬�Ȁ��Z}˚���ŋ�v#������C��:x����ɥ^G�{�L�j-��6��+��=���)��f(�/��B�Z�r�_���;��xeӣ��u����erH��d>�t��Gu��3{�[����('U�YXE�-v�2�h�ɘ9j*���m�N";4�c��^9X�	t6���ڥ6�c4N�,bM�I�^�[Tw�&�~?�����j�~�;�{��y��<���Z�p�{�c��ZL;�cM�j��qy4���A���rsm6�,�1b٫확��SU@�8n�S�p�:�Ez��pk�m
ϔ�;�H����BY�u1�Ƭ�WLi�b�/��	�K�gX�`�jL��o�\f R�fV���{�i�`ˇj���K�'���2#���'�����q��p�
,�xz:���̻�u��⻮�Cfq�yR�;���,&�/d��H;�.���q<;F1�ϋ[$�4�o�tõm��r]4re�&v~���:�jn� v�8sq�QL���#��ۤ���M;�S��n.YWt̻�ܧ�[,���^�q�M"��)�k���D�b�"L�W ;�{C�Ü��kAu�ɲ�^)f�����=�"MV>s@21���FFc����	��@��s]����7���x�۽Y�"�����؋
���R�<df�H���5�Q�ԉ��1z��tD7�D�.͋��tˋ��l��T�(�En\�*g������y&��*��`�j6Q���χ>!1��Ӣľ옄ڼ���R��}�{����2���z�����ztXG�t��&@ U��9��[!ЇX�(�X;���D�
1�7`�1��s(�3"4�h�J.���P����ߓ=�D�u+>��Ϝ���y�lk�k����>���p���v�w:{���N� �=��W)T<�w����+�xU��9�L�KG��i��n��{����m��]Zs����]��k�8�-�;<�c	P�X�b�2&س�؆�e�#��8�f-;�Z�˶b�Kv�&�Z�u�t5�����+�:8��F���ᑬp3�
%�Oo��%+�շo5HȽ�*�$���I�z_��Dϼ6�WK
�|M)>�I��G��s��1;לn`�m�3�O6���"�Ť�\5:�w���n�T=ƟG�*a.���ұ�t�FS6��S���:�<7 ��Ɉ7�8���@8�p�kE<n�F����?���[ok"���M��gf���*/�UH�6�C��pN&�r��������X���2"�ٙOen\�*�6�xʨ��P�h&��^�K�L�z��ŋ[u��ۄG�'��
/�L[�lޗ<a�43��-fhܜi�vݝ��$�X'�sQ^�[;M�������QD�t�6��;\�}-������k<X��SZ�ר�෩��N�-��\�Q5L{O[jd�� b�f��P�_�&��̋�W���^s���G��s�	k}�ead
�����/G@hj�O�9�;�~�s�w�i����;�<����̺.�n �+��@�$������/qy�4��]�N���U��Λ�[W�u����wL�:���t�i��Ӽ�su{Y_����>>5^�Q���kwG1�Q������a�t�\�.m�	G,O@G5L�	76d�݌�݇n(�m\;��Z�;�q�̧!���X�1<�z��_�Ц���4O<|&��P7W���moGV�e2�|D��t*�d�<4�j<�Ԝ��.��)�/�S�:��tL����&;.锼^٬�N��S'��S��
◘Jw^��x�t�������"���/Y�k>ژlRwo-;�hG�Ύ֑��l��%0�m�4vk���N��0�yދ�"�ED�S=M�%S�O���]�Ri{\#]���kW�lto55���^I�߷�,n=����V�L�E�oK�+ʦ����b��� 5�ZLŹM�zS��֮��;�׵=�y'�i�FcO'�����V\LuL�M��,��:q��qηQ ���p̌��A��e-�5�y�$��k�{É1R���bU����:�8�� ����,,��y�h�FD41�٣C1B9�fy�6�c�uh܆�X[y�K���p�0�k��g����{�����*�矬K\�ԡoU���RM_��v��1����+���S��-LA�P��8�0�D��n\�[�2^͇�|�R
�t^�T�,�:��f�)���[l�'�� 5��1uv��@�qD3f�ɭVգ���Z��i;ݣYݙ����W�\����Ã�ϰ�m����g��^�zsf����bI��)��ֹ�t�=�=�?F`���j��o~1r�������4�6w]Ɯ��o�|N՛���~�`�s��Y��m�����s��,�81i���0�O6��G��ٝp3��9#�B��!DW0�z�Lfjt��y��Y�5���i@0��+�O��ϩ�X���۸c�`���@��A"�S䥒_��i�C�_<N�t�C7�%�dܺi�o���t���_~.���r�_��7�u��-�w�b�̵�F���檽�VL�	<[H�D�w��,��>v�ုr�T�I0���K8�g��h9���rN�+2�5����d�{�ʓ?<EUƇ�[�pfP�:'�����Z{�Փ/�4MƢPc��P:qmC�ΎkZhM��A��(�j���&��z^%���Nr��zׅ��a֝<��<�"���.���f��#�֤V-�.�]�^~E`��]o�C�6��w֋��Ց�d�6ȧ�\
���q�j���)�))O�v��̻ۘ{^uk�-r����י�	��<�Қ7��$_yĨB��6�.8�c�3m-k��#^ӊ�����չ|�jc�P8 �\�hX�8���v�����Y7�_8����H��V�|Aӏ��o�@,��c���\�(���<5l�p���|��� � ���E7>����sϜVϋ��B����-��v7Z�@ݘZ݋tPv�\;&���[&mq܉�u��t����vP���;Ya����3�g(�����=j���SC�*�)	z�|ws��j�I4�~�{�Z8o��{[�??�Yy7>����1��vO}��y��_1]����acZ�}���d�v�((RP'o:x��ˌ6�zz��Ѧ=��M�/�;�.u�]��<����u:��3��ݶ���<�JhzΑ n�&A-�l����S6`o=;q���o{,nֺ1(���*�5��
���v��hD&�?{���ܜi}�V��τd���;z��gwf,{���;��Q=�!�Ƃ���g,L��T�z={���ӧ�K=�4 �m��.i+�9�S�W�K�l�������k2��+�GSX^�L�mS��A~����r�o)�n�`�O��jD����w��]����xv�hj��ߓ9�k4SP�K^t3lܚ�w`OW�U��s[�P�|���Ì��j�fh�tS���0��m�^H�����{�p~����]5�_sC�<5��	�V5�$�ӹ�dn�o|��n	�Ϝ�5#��G�'��۴R`�ࠎ��*�+9#ۙi�C�S���@��4� �5Da��k.h9�ٝ�,YV�'Cг�iH��4�nq���\ �E�"f\�QGٳ�o+�CûAy|jx��2��!�����߽�>>>�y�1[��o�=�"܂]�>ۇ1�����~D[мy����\�ԥR&�b�"M�wv���h�v4�ڪ�j���-~��F�eM��Ϲ�h�q���ъ�g��)�6ի���.�T����W��2r�M��b*َX���!����Vzc�mqC6!&���y�k�Ħ[3�/©��>;�z����0smN^�Yb�ܸ�;x�{O����qeE�SM�u�s ���mI��+��?=T=�XT�4eK�X�AZ�L�v�-���!]����5 +c��Ӛɺa��O��c���,S�)S�Je�γP���~�ϵ��β�h�]6�:N�)�)J��(�
��r
8%i�H�Ob\[��_{���"��P�J���w~Mu/�z�-��=4�M�E�XV���x�4�x6�����-m�*��A, ��|jN�C��	<٭Q�����h*.2x�|3PR-~<t�
�n�W<LZǯ���y)hi@,z.����;0�0�o@a������o��L����ǵ��=���a����$~��;6�#+E8���#<�:!�.iW;-�Ӟ�B���o�H��/���Ru����Ad��^����|�Tc��.����Ll�V�v�]fo�#Ȗ�0�V�ݰ�d�z��m��[����ãu+j��������y������ђ�>]_�W��H3�����y��j�׾g%5�b�Q]�;�&�O��9n�>1`\W2��q�ژ��gE�v�g-�r�x��!F[���c���i�TѻZ�ʡ���0z�b��~L�ƭw����{�AAw��/��(���[:�5�@g�	ڶ�<5m=�.�|\���jt
��E���(�`�5T���܃�33��5٩����i� ``������-v�ǒ�"&���/����H�b%P[6�#��l=���I�����L 0�>�P�M@�zG��N�L�������v��	�J�Ή��xo��1��כڿ~�Rq�"|���0��Pj��p[�ϊ1�[�m�l;�]Ee�9+]��X]2W5z���	\���'��Q��n�@�w�o�̓ؔ�*q�l�]5�t&�dW�G�ƴ&DO�L#�a)��)E���n�v�<Aj68OW'�f�x��u
5�S��~9&�p�
��}#�sn|��6�Rl6i�N���N�5��zBTO겉���?bٚ�������5����V[�~�u�|��
�7�i��4����2�ם+ֳU[�>�Y(y W�5�k��0��Vt]f�Z�QWc^�+�3+jA����W��*KP�J[LDc��>��ѱ���^0��{��ڻ�X�Z�D����;�a�!9ƁL�D�N�j���;m�J���y����Qx9���KV�df�2P��g�.v0R!��K�2��P���P�I���`��	���9ڣ��O'�����Ȏ���Sߣ�&l���p`����a�.p�{ؓW�����-������W�l�$�y�H��1�͌0q�c� ���Ypٰs.k�o�j�/ H�a�eVn�<�`��$�t��$��Ѽ������#��b=Y��y���r���8A���P��h�己�*�kuuc�ݬ���Z����,�k����t@�~��w�\����gjg憮����om]��V�"iN��iƽ,!'�M���+ͻU#4��x7�.�f��^�=���Yl���<��]����h��l����JՎ�x��]�7;�<�cS�ww�\jV���t�s��s�mn�?��?U<�Q]��\@�*�t��iM��D��%䌏.�[pƫe�ڎƋG��}�ɶ\���r�F��w�if�jvcL��3N$�C��׾[!��4וW~4�k,X	��!-��҆d�]��)��}9�Ǜ˵�����A!������u+5X�U\]XmM�0��l�s���.�֑����9�t�k�ż��-��Bm�9��t&R�[Gk:m�ˊ9��h+|��_U�~������l�|+��є�2�F���Y�v.�������9��rh՞�9`o�:"�,���B�@Fl��,���u�Z�-tRn�o�EkRK��c�>OA�V�v�?dܝ��lq4ͤ�[��f��2���<&�+�q��xR��.�y^@��J�#��.���-�3�w�[�٦Q�� ����1��1M��N
DzA1�����W?�OV�N݁��no�c�3����;�|$��r�*��ˑu���;�閿�C7��cu�P$��D^曲5��4��N�f�r)�˝����(O��fp�dY�2�喵�dw���MZ��-����"+^�����A�l�3���fQ����+�1�
�ɼkfbMt������fWL#��)Ku��F��vV�|�[����;�E�>L�����}8:ݩ�x��l;�.�	֍��5��-Fٹ̘�@��{*X)Of9��h�~L+֓�������g�m���u�U���;��Tȃ'���-z�`2�7Sl�O���Z��ӱ}"Gsܴ���F`���[mV�M��t��x�3�[q[��s��/�H�:��[SW56c�
NfĚ�m���軌4���\l���2Y:�vr评è8о�z�ɦ>��/i�:�yt���>wG�f�u�^}�S��Mv��ϐ�;8V��li�rb׫�[�;4��zu�,�7x<��ohmbOR��bۭ�9��f��sJ�Ƀ��wf�}��8����Hk�'�dNΓ�)��Bn%�:d�\�#�]t@���\��=�v�[K�RT�cv�T�A�z�R���lQywRg&!�.�֦{��ݲ��&�͎�.
�]�}9��Җ�0�cBs�WP�c�yM���oi���Y-�m�bu�7�d!�Ԯ�!���XN魮ZQT�t������*J�r���1Y�i�Į���HIٸ�\�y�hCw5;Z)���P���IMFv�k#���Д�qL���  ;c�oܩ�zt��o'��B̽y�6��݆%�2g(j��"�5��
�g8�o97fb�,a��&���=�2�8���yH�7zP��V����U�f,q��V����ܨ�VY� [��gYzL�-Uw��HؙcKU5��%�m��`^>��æ@3�TY-w�wY�� �&u(y _9���8�Fe�ÁM#��<i���/F�F◭��Y�.�$�\;���.PO�:��/�X�!�o����z{L��
D={�:��^V��o|N2��fSc�1F�wL	�H�gL���n�j�oz`���{�1�H���ݗ�f��m�E�T��r�VS�,��K���ȡ��yj�O��X���.�7S,���v�騫f�.���M�1CpL�A�5w7���]��h��D;�pZ2��Jg��&��e�q�!���}����r����x�Řjf�6�Ԝy�3^�}���3z�d4��}p�����:�v����;��!\m�:z胘�Զ������1i�2��@�,_�ʇ��޴�  }�I;�����v�.����-W&sQ��}�Q�!�Lt���t:�@v��{c��w^��z�tE]l�98��Y�=t���Z�S�� o{�H�Ng��[�dmC˦4P�ָ�c�=}O���m�QF��bc��y݀$�=o��x�u�(��}��L�|�#�8�p��sWG�ӊQc��|dԟs}r�)�V�#����Z�t���:����˞ݽ�;B�9�=��O0��{�������K��k�'�}7w�Jm|U���=���yk�� V�^㫚��-�}��ޮ��ٔV�Gj(�@!�hS��i�ڗ���A6�۩p�S��}V �����Sc�Ua�8es�����7�N�[��%�!��-X��\ґ-ʙN�b��ތ8�f���;�u�i�pU���l�C��������!�Ov%��F�B�֕ۖn�!���V[~'��qV���f�%/t��.�TiҦ�
�d7H4��@�b̻�>��'��9���������7燞)���(�������)(���((;�LTREA@�I�g>?__ׯǯ�^�z��������}~�_�N��EM4����TQL�QQ,T�JU�h���(��f�"~��>?_^�z���ׯ^�=}}}}~��_���Jk��b)�����b��h
����U�QD�34D�AZ]v5QS@�DSR�MF�sT�>F�
")(��"�J�Z
(�)(i(� �Hb(��(�f��C��$��*X�j&&��֢�Z9#�AE�QG�kF(�h"�&"��(�J�j�� 
����飒bh�
yg�TQEP�Ƙ�N���

�("J}�4ҕA4���AFƤ�b��((��I�&���"%(���N`��TPDIT��PKAAEP�@�BSS153͂���a�}�dP��P�|әH���\�����f���5z����9t����G��2l׽ľ-T���aja�[��J���
�@�"�I&ʢI*���^���y����Eg`������>���g�']��Z`2*94v������Z�aU��n{f�q��ڎ<�%�ivk��ɮp�!E�GSP�ދ�����=�f�J ���N�q��Q7ʤ�ez�8����
[6L��"�<��V�I�0����
A��`v`"�v��������5E;�z���e��=�rz�����;nc��J�H��h��� s*i��S�z�[ЎҸQ��� ֫�vw�;�G���{I^��l�Pu��Ycz mx3#�MsdF�f:=�W�)��@���աF�����ژ�;�,1{VKV�V�����d���	��*l��\`�P�rnzǹ׽5�ܓ����7��*P.K)���͏=zݜ��z�́����n�8v�5��3���)�n2:4y]̼����AV�BS����Y�軇�&�5�"AZݏnV�����*9�^.�����p����龝"v��0��[NXI���
#a���CcӴ8�W_�c��^��҈��1/�c0T@��/4� �C�K2�;P=�0&vZo���ٖsa�B���`SEa�TK&7]�����-Ü�<2��4�����k~����t������p�;.'It'#��j�U�i��B���z5T&�fi��5��c>�_�7�����1b��G!oI�a���[Bh��?C��)�(%���S�#'�f��n<��ڭf,g��0�iѹ�X��`��o����_�dn��a>��d�9g�Y��J8��3j�UH������źJ�&�+"C	���hv����:}��H�G�3�ao�E�4��f~S��Y�������U�j������q��<״.(�ɬ�j����)}��|�� ����z4��#�oH�;:����q�'9�:9�MD�-�;���Ka�5����Fل�� 5�_0���@~��?\BϾu]h,�����=����*��4������`�c�i��=S�>{���k_a��#���|'��zmvlka8ݥ���)=���LeOdG��k�/J���l
�_���~<����yf�������b��Ιd�!P�k���0e���}4�	y;	D M��]z��D�B�#G��n����g��%�컻W����4h׃oEvf<�oS�Jd�X<G����Br���h�=��rwq�<������sf]�dwb(�U��N�s61���pw���ʜ���_V3�k"�eӸs�
�0�JWq�z�x�Z��3�f�ZKU�Z@�S��w�j��}�
}^o�y������{�e�O.�M��O�2��X�Ɗ8V��U4i4c� ���t�"`���fji����)���8�f�����U���W6D���É�vT��a�.�5c*�b���<7O/,���Vs�i��1&'�r��(�X\��^��wy�����f�\Ig����E��˖"C��v�a�݀؝kΣy�d�f�};#�,m7��Š[�0�Y�&n��P"L{C���<_���Ўs��TJ�W��ںC��S��6�X6Ӫ�U5��j����T2�{:du����=��j�͟C�N��kb�u=Ls�wwf��;{���z
����ά��9���pݼ͉X�Ɲ�9	qY��S�g0��v����-��Ji����̍�[�ۜ�9rsu1�eU����S&H`����Y�UGvR���g>Pސ�zA~"����4����v��^��W:�TRW:��>���/(wO�߻l�w�hA�c�.fm�	�>�xn�J�^�0��Y�g@�9S�2���w�z�0�v�#�'�������P�]u�1c�χ�(\8=�k[�K���%k���ُqz{;{����[:8�.�K��:<�ʮ�������9ݝ���������ӱ�B �po��FM�]��Ã���Nĺ������}�zO[E���7)�<�>�Tv�T�o{��jǊvLH���s;��eq�SXR4WT���d�l`��t� �T=.���gt"?J�a4d�Y�}`�!u�¯y�ԕ�Y�!�	kF���<l�P���tIgA���Z�-2�m�!�vhWQ=
��u�JW*�ݣ֩<�xQ�j]cc�SY�x����.y��*kq,���V�u^��l�P���o����S�e��͚p)��m]�Y*�)&ZEs�n*n�5�ĸ5Y���L��V�/��Ә����U��M��mܻZ[fa�6�,�Z�q;�[�x����'��	'@ېY��~>���;��m�Ƴ&f�9�w�#�h�.��ĺ���_�qq�����[Q��)����0l^�$VN�V-8���]喙�߳oxqp�-�T+,�Y:��ۺ��Έգ1�7\w�7RQo&���K��8��X-����]�F:���vbǈ�������F��\�[ʝª9w��Y��X4φcVН�}�#�����)�@7k�X9�xy�|p�������Ͽ�{��}D�\�����s����ݾ���Ve�x,W�V�U����/�y�n�p��Ox���}��밥�Y�>�;�>q�#۟�������N{ٺp��%�a)%o���U�Ϫ֛΋�\�˽���8�]VA��1H�8���rP/3N���c�A�U������b�T%�`7V�N�ؤ��Z�*�:�W+�mf�Hl3em�p���}�Vw�oF�k�u:�8�k�U����*�V�H��л�HWZP�W�t�`�j�CҖQ�Gy����o��|�@zɢ�u��7��x�U*�qj��ą\���~wg�h<myʵ�X�fT�g@�����ɆQ�<>J�P_�ʻ��S����Lw�Y��"�[W'id�0��[�2��F�N��`]r��[q-t(r���K���Tn���S
���9gW��v������oJ���u=�[׊�vs1�?h�5V��jP�db�'Ct���d�MӇ�����I���ȏw��Lr��w<�[ҷE�8�ۙN�M\A}_��y��7�����;<-TMKDr�����
�� �8ɣ�Rᐯ�����tçm~������wL{+1or���J�]�{F�5�d�+�o,ԩ/;U�͍Z=�ϫ��^w-�J��癊ڇ�9I���Ss�D�ZK�y�������C	�oy�L@��j{xs���3WR��K��r�wg��:�Y��ۆ')��ӌ�no�+�k��abЗr�n�`�q�9ۃ�����֡��{̰9���C������)tm���Uڏwe�-.}���ia��i��;^' ���ì�G�az[\�����Do�&.s۾��\�Z�����m�[ +ˣ�i�z�����3ߩ�{:���E�N/�}p��^�kwxǎ�U9'�:K���M�ָ~��#�+����[��+��C!ーQ�2��~�����2�Yp�Wv���q�3��z7���CʏK�H�({5��2���G?p���^�alKz����޻�� '��7qb"�7&���3��}�1��:���ld���7����*��ԫZ��{'�;oF�s���XY����m�>�7 �}�y�>�3zw.[��X�|��>>>5꤆��N�_ْ���}�'F�{4�h�ڥ����b0�=�]5�cm��uU�J@?G�8鞫�&NVw>�/4M����us*�+O��u;�+Å�+�f˸,�ƜV��EJ_<V��Qu1[b�s/S�ޚ�I\\�n�w�o38�3����0�y�5����Z�RP�Xw�o2�����߽}���=ԲG+���Yą�e�L��5��yCf��T�s�/٤��2��@�^�����Qp;�������{��/���k(mU����-��������+��S>wWE_O���z�L�"�&���{��މ�ÞT���K�,�9� ��y�[��%�{7¥A-ڵ�������Wwk�Q�z��ϝ9 �xe�w���y�ìؠ5sG����l���Sn���Rv��;n/N����P����	��ӷ�0���@�g툯U�9x�f�U�s�MT�+06Uo#��#�|O�����ݞ����㼩b�����ػ���Z�"眛#��kN����G�7hhؤ�=�)k���RŐ��U��^�>��g؎_KnG�sv��8ȃh�Ǌ[����7�o7�x���ڶ��O�0�^�R�+Wr�YKx4M#���@d2��H��-�j����A[Dx3������Rg�gk��]?;U����飲��~{����s���KV��4@��2�7���x��[��=�Y���gm6��X�	�kj�����k{�>7��G��`��U%wB�l�೅-��ʉJ�s��Զw�7 ���Zm{(b�y�v�"7�N��S{/�}u���]=��j�I��y�zE �Y]���j�6�\��fQ���-G�2�ꊩN��"tDl�����<7�x���7��T��h�Z��v`i���ȦY����u�2�Up����my���Tڲ�j�g��G�XQ&$�X�ǘ;uw]=��mD��&3�O�]��ΪU#��J��@y/O���n֮���Cg�tG$�Wf��U�d�Gd��9>�w-�ߥ��0���� 2��&�r�\�|K)!(��׊P����un�g��z`�T�q��z_�K>c�z�C�#�|��4�;4F�MRj��H��k ���L�s�WJ7 ���"���x���%���X,7uX�������k�s�;���A�2+��*4���EQ�ϻ��������d7+�� ĴS	�Ol�h٨ȿ�By��Z׮��%�͍7���̙���ۛ��v�S��v6L�@���[���"�	��V�&os���m�mnN�Í[�;�ӗ�k]5!�o���gJ���UyL�*�96n�5�x�kw�66�bKx6�G�K��`h)r푐j�����5��J��c�;/3�]�i�i��>����ηs��.�[A�:�71��~<�m�U.�����͙t�&ٶ<���V(�lZ��<˂����~�7O)�g3\>�++k5�K䷱��7�{{ݵ -���᳷1*�ݪ�^���ݭ��Cf��~�%�x���H*��Ӿ��0S���g���/P�9�f�	`8����,
��>������/�t_k`V����p��]6�F\b����3�vJȎ��H�H�[GT��t�l��5iU�FΔ�I\C�l�ٮ��[^��܆v�{cZ���{)Wg,RS��@�gk"��(�>�D�Y�q��=��ۻ�Ղ��a��[��%�S*t�ǡ�,p�t�[f�wF�u�kM�ʅX�m�r���ra�w���y��ﮏcoD;��`�&K]j��.xPq�C��e���)���w����$�Ϊ��Ͳ�u��E��v�R���3 .~�$.=�������kCʋ���ɞʶ��ƃ��e��h�R��CC��t�@zC�I�ě���8���{n#�;�x�S�K����9�	m ���}���bvw}��U۱�����ҹײ+U^��b��R]��pڪ;�J���5Bh��=9����kmW{�R�y�5L�M�W��̖];<s+��ѳu;�ZLhaۈ�f_��)�yC�lJ����5j.�;OߟO>��z��'�>?��+������_�IF�����f@�֥F�Z�F�aD�����-��8uǝvl��<�ھ��V�[�Pn���.���T�}�U��T��c5p�,2����a�Ϥ�����qj�n�p#�� ��e���3f:�T�J�ְsd��_� �#��s##wOP��M`O%fe��T�"z�J�[@\�P��U�,�i��ރ�aH�*h}7z����l�k3{]+�1���Tt������ﭛ�b&!��w�����:�v���a������
ɓ��ԙϜ�l��c"�ҝz��D�=k:�C:�giwج��$jc\(6�J�����o4�p^�95c��G�3#���勳 נ��y��cV-��E�R�dJޅ��]Z��R�%qe!9V�̬�c{��p�Ú�m6v�+@5����x�捧��i%����̛�:���x�(��w�ה�*zu	��ņG��yu���T���u�S�kV�%��,���+��=��cs7{)�k�p��op�o�x��'=^W�;�~�{'���ݻ�̡0P|��!)��}�vui������+�%���׆�c���;����;�i떌����-���!E�n�������߷��JUз��R���A�m���eh�Z6�v3��%�Iշ�NE�tiy/���"���od4+P��_],�[nh##f}� Ňk���=�x�V7iTA�7;v�.�v�w��g�*�*qsI�;�-�@MH�}C���i������'mq[n��)ֵ������1[(%"���q��� UQ���9�(.��f�6��2���1�h�B��ޫ��d����T2m=+ES�F����?�{mR�7%��O�&��rņ�H��?r��K�4� �c�y�3��q�i
�&J��u�}���&_W
�x��8�U�n��D���8X����H�;:�U���
0�o6s���LQ���G���n����4�GX`��&���ޖn�1ٳ)Qiv�]ܵ�.I@����ӻ�z�V�{H�0�S_�T����hhWW[��V��+���;r��`�q
���S�s;z0��'��aՎܚ!���J�%���s��ͩ�\��V<�>��N�3{!j9O�:{��}ϗN�5�)J�q�m֐�n�!�N\���S{y]QvZc�;�n��ؔ�U4�4Nu�HQ�z���Y�΢���b�w�Z�J�x��N�sF�'<�k�l�s=��
�C#L�Eӧ"]��EK�Qiqze7w������b��<���c��鲹���m$�.I+-�E	�N�f#�f\p��]I���<+4���nft'v���a�M�hel���Q�HQ�y*ǅ:�%t;���;�p���N��|�@,z�^;)����pS�f���KXF����B��{��^��k�Q2�/-��F�[�쮮Z�`��!�ة�\��]�wk��N)��X��̸�ɊWl��mu΋��U�Q�wz{)"#a�V,���-ѭ���-���h����<�6������yQTRU�^�������I"�b"�����4QG�觘�u�������~�^=z��ׯ�������������DE�#KE)Q`�IT4r4�1%U5K�?cE�珯�ׯ�׮z��ׯ_______�����I(��*J*�J
B���� ��������h�� �QT�RRU$HRPRD�4}�!Z&(h��JJ)j(�� �
�SM44ԔKE:t�4LM��(�-�N�*(	������j���&��(QHUQH�T�MICA���QT��΢H���f*�a�NN�����&)��("SlRD�T�@U����MSA�4SIL���*J��(�� �CATQU��i����9�q@45C�F��*��vtPDla�C���*�lQR�S�E1-!A$<�AH{8�m-!EB�&�K�uM�8����q��󿟻��߇�K�f��:�������%�R�E	����dZ\}N�����2^��%M����*i�c�����0�s�-�iaF�'�׿{��F�^;Xc�\���P����Y}�CiØ���Sq��;zҶ�n�f�~�����<����ei�l��UHÛSj�wc6u�_�	os��4���%���O^�R#8�@a��t]MI�ƚkj�V_m1��A�	P�
�q��o3�*:��?cB]�~�jSꉩ�?d���ֱ��������?��0�;lP�ؠn��F�\�A�5J5v��H�]��u�3\1�-[�L��k�uLQ�v\^w<Hw��Ƌ���w�c�n���c�'��_� ����������]��]1]��������k�v�՘�".*/��N����UQ>�"�.���jT�Bm���E��	�U+�d�,�׊���٥m(Zy��+r$����_momf���>�Y9"��k�HJMtZ�̪�Բ�{��Xp;��f�A2K�@��i�::�WS	��	�~�Ƿ�&�4z���j���T�f�{:�k{�=x���#��}�L[;�	'o&�����.N�c�G#嵒�j�7}�Ԩ�E�Ih�{�H�V����X���E��MN�>^o7�ެ~�����"�!��7��c�-vImJB]�@kג��6������ɮ��y�.���`g�1�}
���/���ѽ�T��P,�Z�{U|�r��!���˺���^�,�������ן�J�5��mε�
�]9�6��GS�Y�� �v��+����k�*��k2��C��vU��>��U������y�̵-�u�O�
�գ���07��䛧��"�n���o�Y��w��#Q�nj�]5��Q��ټ@s#}V��:��1l>U�fn<�[ Tk���1�U׻�����l�ڸ���5YY�;r�����6:��p��}"�Z�[ƾ_/e�b�ˮz���;5����ڻ��@��a�Bg����ȱ����U?���s=4β�~�ή��7k)x)��v�q�XƖ3ۚ�d��uMtn񱚥��8�Sj�r��y��mަ(�Ч��[RI$�7O�,rYՋ�sUޫը�f�l�-m]7AX;(���F�ܩ
��Kxz"����xRRHK��';HV<ʖ�h-J]��ǩ,�7��ubπ̳)�:(�+�����.�qYjUōM�1E��s.���\�P�	�Y(I�e�h�T�N�{��o0f�7lm���P��ǫ3�k��ʉ}R��O��ng��T#��Km��Rص�q�)�ɻ��]bڐ����U3>��3��@Uoӓ(v䊚^��S�0�%&�	�:��)�YQr;�{+�W&�Z���{�<=�6�tZћs�1����6뫟bW�ݴ��fuj�qǊo������ ^A��Gr<S{zjy�
��kv }xJ�ҙ�![�{Y�UQQ��Ւ*�oO=�dǍ0�J��n����Nq���O�-8��)΃����b�z�W���_i>�A����%��?��W{N��,����*�y���4��{2;6�ԵQ�ĺ���@�����؎Z�5{Q)��5��,�\��Mѩ�*�bG���gq�K�x*Q��~����\�+���;ĥ�#X	��B�{}�*̜\�ܰ��ў���hP�J����u��e*)on�a�}tE�ch�X��u�#��J駌γ�]k������Q��$Qh�t~A�O�GC.��ۅ%Ԭ�0M9�z���m��`���xL
I����{�4�'�k��O����֭���y���9[ݝu�r�"/ǵ�A�J<�����ٜ�;�[{�O'�;�5�E6��ݡ��\�h�bv��-�nutZ��Dq�k���0�%��Z���E�W�7)��螞i��9�o���l8�e���c8��?vk9��+)fH�v��=ʝk�l`k��=��ym��zorr��x�V��&_����pwsU��A�u��eDlv?s���)���ݠg�� �ey�TϪ���%t�B�9E�y6I�ū��P�������S��$�P~h�G�[�S�L>��d$���[�]�^���旣�Vϗ���6�d�u��^n;@ȖqXok됼f���[g��^�*/kK\f6�=�Ǳ�n&��٬�-%���`b��ꢴU��j�dӶ�.#m��]�{�ۣ��+C�,l�{y�*��޴^J��2�/M��^6��F?V���z&�f��A8'i�{5�Y��Қ�uv#K��S���J�ɹˆ����wK\����(i��W[���5��'�,�ʕ�#�	�m�O���#ms��/]X�%g��$*�Ê�}������i+����>>o}sw�z���k�,��ӿ��}�F3�W�v�ͮŰ%u�q��V��6>1�x��WUd�V,ӯ^��
Oy/��+�Ov6ny&�[�St����5/,hw��|S$�q�ӵ�p�u�nf��O�\��׏f�ėv,GyD�������h���S����f1��k�].��\�5S���Y�i��x�OcoN���ג���d�����1� Jc�a�8w�'B�CóN�b�zbb/q���!��es.z�����=����lc�\�P�ƹ���9��C����V�K�LO�w%���Tp�����[��PpFn���]������>MW� .�&�S�iG.&�]��+�3S2`3)��ҩ���� 9��Ωީ��>k��yӌ֗V��-�
ڪ6�2��>��u*��g8�o�A��G�-�����V�~�x���5��o]gzǨl�_���[����`��(�V=̊}Ȉ��eZ8rv��C[� ww�w�I
N+a���Ӻ��ZbJ�Hч�0Wކ�aMދ�Gu���P�m��;F8Q]oXM��ռ���l_ft�%��n$v��y{�����gox���B_2I͆T0��ql�[)4��� L�[mC��x��˴v�h�{������g)uy�_ԥ���d��s�c�Q&9���|�$Ѵ���kX`v �n��b	ǄOB�5]̬��P9Fe��l�ln�������]�����}��:�ZN�ҋ�W���f��¢�U�|��e���$�ٞ��E��ϩRU�G٩NT�Yz��%���u�e�������m�������q8��K�]�g�:w'1�D,�}��5�[U��;%z˛��Z�
�(>�Kt,���S8�4%��5��۵W���3f�>��n��\��ǵ+��,�nU�l��͖���ƚ ؝���[��o�t8ʽؑIZ��J.�v,4�Q����@l{v团��e�˞�˞���SM�z���oT�Қ+��^��D�:�f�b��`[H���3�E��5-B�h�PU�bx7.Y��u�5鞖)��+��snk��d"mvΗ���Б;�R�H��6�͠E)����zI3*۔vr�y��٪M�o���v록u���j������uC���V͛��wc$���$$(A#H��3U�������绝�3ݨ�{t�[�\=q|�Yݳ��Ë�
<�^�҄�Yx�w�}��Fz|��E0�C����߯�����Y�H��)�\L��������M/���`$W�ʘχ3S��ܦ���;����ew͌�'&���2k���*���Xڰ�ns8~j"bk�w�9�z�+^]��6�����/q�4*B����#��^hUc����V��1�]�{QNu�y�ȭ�꼞*`L���ގh��_sU�TTr�g���Bki�3�-��kz;�۷Ǣ 6©�v=C{�L
�7��`J�Ӕ9dG68aIV�n������ۀ%��4�(�r����S]�����v�q���z�L��� �(c�'�ѽ_*�c=Y���z��!�Q\(J��y�luP$�p���.k2�^���ݻ3]7 OR�UO}�00��G�,� ��oDF����nԂ��N�z���gwZҨ7$�Q���ź�����a�Հa���Ow"�U�cY���!�(SQ�t�����3�t$�^�J�`�Af��Qg>�����rq^=���}��N���<�ꔷ�^m��yy��o^M��sk_�Kj��^R�xɦ��(��N��]՝yr"�y���"��6��0+���f��Kx6b['�x�\_Zk���%6�gi�՘���Ӎ��ٓ� en��,��)]˝���Db��ڽ߫���X�^�������5��B]wW���y�:�\�K
����q��
��&Q���2,9|y�A+=���b7�<����V�ƺ?~|@�ƞj!x�$��Ӽ���#�R� o�����/�i�`�gRT��M�(�jt^4+�kk`h!�{����{�p�����/��)3��� ���p��z�F�ȣ�c��8�jaw՟E��+��T�5��a����w�?�@_H��ګ���/V��*���4FvxH̺3V�3�to
9H|�eOM��6=��s��כu���g���M����v�	�4G3��<bB�f����,��4�\Ыi]�߷���LQ,��#��XD��l�&Ku�D��e��&�f�u��IM����*�{h��9�k���,���PO�U�\�}�k���Z辒��w��k[J�9�`�6�W�
u����`�������?=�w{��Z�]%ǩ�YV9A�����V��,��1V�T7=�ogk��Lwt��̵7��{��h3�V>�;4���YY��tQ7<;ݾ�B�og��j���#�`���2���;��&�0p>�y7];������x�ޑ���y%�jrT�T�G�QvƗ��\ˑ$����Y�Qy@/���vEpa3��]��g�=�+6�Z�Uϟ��'2������w�57�\��u;s���Za3|`X��	O�����3�w64���ʐ_bww7kbȃN���T�uǟ{6E�8����_]R9�6:^:&�]_d�ؽz͓x��=�����m[ �
�ö8ܺDnR�r��[��׬^�oU��g��w�����p��G�^�i�Vt|L퐩��_[;�[T7N�GS�?����%�*��n��~��D0$������!�����&��e�;}�:�>���;u�5v��9у0_�m�Ө�͡�G�ܕײ�U�3Ք�Y��3z�
Y\zL%��-�Нk��X\N�7�RI#@�(�;n����!�B�n�����׶,5E]���y�����B�M��mG�����;mY����ֶ瑝�<q��y��*�Nf'Ͳ!0ᦺm(ԺⱲ_�>�}��� j�)l	l������s�������e`�t�h����t��p:��}��b��eϳ���`Z'�,ȋ}�B�[/6��a�2��m�s���>'v��(x��$
�&`!�'v.������:���ג���BmA�5��:��w�r1�(C�<���DֳYBuB��~��g�_}�4�o,�\�r�ݸ�,ϑ>f�ty����tM�ǫ�����M���Mk�e1X�D�B��R��JnM`�i��ث��\&&��5ݧr�8=e�����1����K� -�����A?J���х{9�娐O)~� S�ܦ\�E�OXֻ0����f�OZ�%��>m�f�c��]D����MZ��,۩3�B��O[���8m-L�%厾��~ڻ�3ڦr��HtM9[rM��shy|׺Ģ́��0y.ٴ�zh��N:��-	��'���s{� �nc؊ߍ�V��"ٗ��B 	vV���,m��4M��l���V�f�*��Rioa趗�%�ת�j'���Q-��LB$y�p�B��@���4���N��t��fW	p�k�*#רN�f��9�Y#��rZyjj֮�tN��*eD�]��p諬Y�2ϻ+ ��ȆZ��9�ov��U��q`�F��G���X�.U���!�v�ѳ�vw�3H��W)�R��.S���+38v�T�:�����q'�Vb�w�.s���;1��	����];|�4\��\�2�LL�Q����������������R�Y[7��Y�HOq_���췊l3T��0����F�e��:��|�,�ӭ�����cz �5����4��Jc�t�1m|Ʋ�^r<B�YQ�s\̚!�_Vꮄ�sOp�f��]S�JR����a
�+���R2������d�h���"���O j��1y�ХQ���2�mI�[X�^�3l&�lŎV�@"q�i_Gv�9ٝ�
]-�dv�N�r�3�����]|<�,c��K\pYSz�
�5�=�5��bq[��0ݡ*P,��H7e<,��NV$�FB��hfާq�ZP͖�7��(�i-��\����B�K�擒���T�l�}e�2��Ẁw"����ơ�nVWs��˶�f��/C�������ϥ0b<ѓdT��#���`g�Nv����J��.��	J�Z�Zp';s̘6h�j�`��yC�p�U�y�JV��R���&�鋜���Z-<��ޥ xT�ȭk^��juy҃�+"ާ��I�������b���ޔD�bي�v&Z|��VAm]��i�
�Y�[J�;�L"�o&e�VT���n���$������pe9�Ҩw�p���WV2�����8he��V�h����P 䶳dYx����gp���J�2I����X2wE��Ɖ�8L���y!�+��Cz���N�T/�q�ޔn��,�.jp�ynX֊rȒ!(^�֔����k�R�JSm�w�2�ثO�L�%`c+�욟VT�{��a�Jw�u��P���R�QT��Z����Op���f�$���w��]C�����a�ɀ7SB�t���5�7����	��q�����&�Dv�Q����φ�29|���HC3���4D0�M������]tܫ�+."�ם�.��gY�����Tk�ν�}\����=}���M	m3Q����ϻ�����&��;V���5]Rά�Ch�Y��c-���:�"KD��tJl2�g,v��:���䫔�r��s���-�Pd)��8ɩJ��aR4�O΁��@ �P�|X�)�|�K0 �U%F��F&�f���P�����%B_6"���UP�D�4�RrMd!4sd(��(�H��<|�����^�z����������~�^��肎�)���*��)*��&"G�i��b-h�����9�����z�z�^�z��������������d�����^΁�R�h���������W��T��h4h�� ��iB������"JS�gH����PP�1�����ǐr�$i�MQ@�Mr5KK�t�IM!MUBDHSCM%%	�J���4Q�(i(

C�fZJՇ@��IHW�y��yih���)NN���hR��
@�JZ�
�&���|K��1"R�%!T�UE y{!ȣ�����  xPᘂ�F�����ϵL�`{��;���>�^�ʜG.gD[���σ��,D㽣8�T�1<����9�ɱL0>ѵ�@H(8�P��R�2�eQ�K�&�G�~�����ob�hg� �=�������K�y*���c+Ɵ� 3,�ю%�c�>`Nٝ,�6�s_Ԫ�SBե^�˫�W�+��p�c�zY�K��H_z��Yo��y������ �מw��u�t�B[��̛ʌTF��� ��F��[����f9�jr�P�����3��ՕI��/�x��شKՆ����ױ���_�׍��<��u:���8��wl�V[�cT���fn3/M�d��k��Fz���G�u�
�zV��|�ݭ���<�j��_5g���<��!�>ޗ>�^a����>�}Z����hrg�QU���;�E������'xU�@�]�Y@�6�3��ֳ�H�����.'�c6"w��X�w�l�:+��d6 �
�y0�:�����[0$3���7��p\Z֎��L�V���s>�p�FvԕP����Vz��n��VJ������\^��G���2\홻�kG{.V.j���I�B��n�．u-ޯ �ٯ�̴M�yy�ό˄��ɆLr�oť9s&ʋqozu�ו�Km��Jg����S��H-��>-�>��|~?v-�;z������*&�_�������e)K��|y�c� xk���fckU��_vS3�f�pS�.s�+����2�f�hNR55�w �}����^d]�{�ܪg�z�duow,�3��B�CB��C�e�w�R��Z�=��w#��dWM�J�UOݙ0i�|�pY�98��Td�;=M)�1��{p<�ݔ�Ir8��j�V���r�,�]�u��s�AC�4.�ʙ��x�5�z��zsK�uf:���je۲�����������L&�ı~X�vǝ��p�.So�6�+u�a$��m6��a���ʰ������ےţ��aM�E�ⷨF0��Ž�}�sQ��W��Q5���m�^�%��b�=xl@8]�M� g��86�6��\kV�M���u��~�m���w�g��/a0�ӽh��.�5���Mu=��� X���wD�?�MIV����w[��'Xo0���;q��n�*���ۻ����Y����j7oT��E���;��z�1wGp��O�������k�i��E�W��9a��),.]5�ۛj��|�||�UU��ݧ�ש�1��{n#w;'��4��/���I�Ȳ�/�W�59��
Ϸ�*P֯Ƥ�͗�}�Tj���b���5����ظv��}u�"�gX�闔f�<V�Y��5�r3���k�����Q5s��Z67��9bVc�l�36�J7��Z���'j���=qoT�<xbY�s��%���\u�4��Y��2ZYd���ӤT5����jـ����I\�D�ް����;4�-���z;ў���@�lϰq�=U ���tM*�6�]�ݼ�z;1���]	M*��U3�eEY[
�#*�8��U7W8���Gv��C�m�;6u��w�_��Rޱ��dm׮�L�zh�Fl�8|_Ml&��^�ʺ�5;����+CN�����=���v¼�ܶWVbR���z(u�d��]o=l�ghz�Lq�R���[�Oqqz��v��VC]6�]�=��0������C:�u�ǽ$}�����L���b|�8>�W�ϝپ�cQ�y*��=�3�9
����^��u��	n�j���L;P`G ݮ۪`O ��쥹y's�D�|-]��qq�n!�r���V�wh_��������]���c!���3]��͟[�����m�h�T����}۱:���K�v�2�n�����8{p�*��4����~��~+s���	?I���+����~��������t�:�8vx��h��s
��eO�VD������;������r֨�0�n��7��}��v�c��X�r{����8,�bz��:��b��K�:�Tk�S�[^���۞�n�9�Z��45�8��3[�i��L0��,�a®�5��Z��eh�;�К����픧��i��C?�<�o��X�!gCݨ�5�2g{g�~_���]���k�Mw����ʹO�(��܆c�gr<�&z��؂*��ӕ�76��7�-o	f&�=�L�`�-rv�:�̙�6(�/��'t�,�6{�ڈ�A�#7����XͲ�qV��ķ@�14T>�U1	������P�h�Mq;�m�)Ku0�u7M8�-�oN�Uw�A�5srr39v� �Xs�������D!LU� Hw���Ǫe��i��]�r�8��='tv�d���8���rjNJ�[��̡�S�R�����\ow`�\l��U��B�R��n��臒����>^>>�2����Ki��b���}�淊��bΪGoZ�]D+�إD>���W�T�vtk\�c+�S��*�joB��!��l�zlt�lҋۚ�����ޣ��]�br���e�ϥz��=�>�qie�+^�{�]�R��ή^r'o�]d�=\O��ٽٗѪ*<��ȸ�\N'�K��۫}9م��2j�����n̓���V�^��[.k�r������Y�m�\ψMٹ�-�-� �U�͝�PY]�;wy^��^���=Eyմ��j��ѹ:�m �]�U:�r��6O�[�U�aQ���l��`�̾�
ݧ3v.���\��b#l�#1+�m¹�0�}5o�1QQU7�$L�K5�r����,	˛g�T'}xsUgv�(9z��mu����W����	�d7@�[L{��C�|����P~Z�B�m��y��z�є�5(������jb�o��6K}��;�%٧Ѭ�+e\�x61�u{���We�B��c��':����ˬ+z��#��Q��1q�9WpȄpo
4vf5��9�hʋ�0.̑�z{S=��K��sr�f�����KwK�_~��d�h��k�n��k����,N�}\�;n��/q��[sX;L���\c%��R�sw�ԁ�r�3ح`���0Ԧ��wh��g��K �-��[�5!q��oB,���F.���snb�6�m^l�lw������2�:�z��sHHS�S�Z��h�ǧ�S|-.y����A��5���ר1��5�ܗIE���+�Xh:P��Y�t=ꨱy��%�}Sޛ�O���p=��k�ݸ*\5�S�Y�z���m��T��t������q�]f=�z�NH�g����p���MSr/:8�3};͙��yZ;��kK;z9����'��	�Y5��dv�/k[j���i8H6ӊKt���~�C�����+z���WQ�W�^z��}��7v��5`b'(�NL⦮Ρz�t���oh�^���^u?�!f��K���2=��Cù#���nC0��J��-ܼ�r�og�<��z�EL�R,T�d�-�<���u/&�^�i����F�|���h��JK2�=hr[؀�v�k_-G�_k;��F��v����j��q뜮���]����9V��H�q�����>:�"�g\�;Z�Lyx��;+��w���e9��0ˠ:���uD�݉aP��%x���u�����ᷓ�O��fr0_�9��f�$�O0X�wUc����u�̍YXs�v�o%�o�Y �� �ˠy��M�]���2U�1�V�w���7�\��@�^8��پ�"����(�SF,uj���50�D�{�(�E�U��n�^�Wqp�Cl�{r�:"�m����nm^�ɋR��j�E
箧�g^Nk���5GXr�1�W�S�䮑����ں��麳��mo��C��E�z���w�� �_+�y֝;��4k�s������E�2

yK��H�X�Ū{�;�<ܛVk1g���#�j^���%�K?���֤2�T�j���x���N3g��-�:�r�;|u�:��溔!jٜlxieå}\���,�\�C�/ԩ�ϟZ˓(�����(���ϲ�����Զjsɾ=!�Q�FE���9ć����]��( ��R�UHA^i�[�;(G��5L�Ev�2��E�P�ПV�.O�.ۛ����9P��N���&b�;���1���멉쎍�m�������9�Y�ba���� b���������`����f�#�7x6ҏB6��6�c�}�n��ȕU��D���ݧs{,�sNv�׭a&�`�Jk�p��4�;[����]e�v���+ζ%�n��^^CW:�x��82�uݍ�l��Oqq�Ԡn�og6VL�EW]���gv�vR�B/�˘�6����սq�S�	���sm0h�1fܗ�|jf�l��R�w.�ۮ�nh��9[�1�a�9n[n��䬞g�x���}�e
�)�`��T�Ͳn�ya��{ma��2:\�t�.�1�]��P�o����k{1rĹ�|�Í�f�~�w�ٶ��ݙU{�r��x/�9�S+`�3)W��+�q���7��=зՇ6����|���s����H�G�c Rpٞ��]E
ץy���g�n�	\���uձ�eC�����9�d*��غ@��.�ݎ�n�R�g"d�c�\�v��^��Tb:�Z����f��T�6��f�j%����U���kMuf��>�iV��FG0�:�n�_�Pd�i]�mgQ�{ /��m]�Yգ�����Z�s�.���/��m:��������~8�3��=ܛJ�`���z.���R��o/�+��u}�z�k��7Kc�!F`ڳ�6ִCMGk����|ݢF�#���@�8�G����:��Jt��S��s�x�7|w6D�'�k O}�ǎw	�Rk��������*��L8�2��NNq��u� KA���L�Ӽ�Cmz����f]���׿_.u����/�{������0�&-s�5�)��:�_s[P��'lA��˙5o{���ص�����hRa7�X���t�yF*��9��w�N�𝋄оK�^��0�;�q�y,�y^O�D��]�^h�ɧ���٩��筳�z@@K���F8�����q=0�Y��\�KKX�,����3�[dVآ!�y������m��wfoun?q�_����V;iz5���?v��FEGss��(�֮m[�r����{^��Z�U��D��O���`Vǵ+S�ܢ&j��m��B���T[��ngf��4V@�V���Sd}�/�@%�n���z�!��Uڵٚ-�]j(�b�էJסjO3�]���qoQ�434.�ܬ������f\]O�j�/꽾��yy,��C���|N���{#52ЖgY��Tb�kͪ�ǋ��۽5ۅt�b7�^�x�f���o�q��׆�N:T�՝��Lbmb����ʶ|�%��i���K�>WEBxgf���Ӫ�N�3W,B˭���ҷ������}l��e���`,��O�%E�kl݉������_����ƾ��n9���c���t����jeb��vUq�yU0�eV�{'���(���9����y�1C�����;���'\sG[�,���G�5z�H\f�q�TN�d/�-�}z�Ǒ���f�U����A�z��%�f�CN9�6�i�ݞ��F5�A���ʺ��b��0�x�7Fd�D��|�{�J`U!���zy�5j�i]��3Y1׳��Ȟ��Ue�~[�*�ʗ�mz��_�À�҄d,ż��M5�b�'���a��nռ-�gTӻ������h�ЇA|8l݊�����"�U�9���]�;�dv�z�f�f4NB_�ݍ9� �[�Sr��׵����}&���"��K��n�n�,=p�]{h0GkWɮ~_L����z�,���*��Œg]��+㤔�Cl#J�\NԶk���ۭ��hk��b,5S7@7��\kt�\yFj�9���3��+u4��w��>ĕV@ �3�w �N�2�kQG���*� HK�������K� ��(��%[����sr1*�*s��.u�����3T�N�]��d����F:%3�<���T��Q��;R޺ͩ)zuN}k��;��'gs�3�a�.��۟gaU�&���zPO3���.�ê�X�������\�m�[l�'LT� [ס�$�9]2[�:sY;�T�Q�}�=��@0���)�o �fV����P�u64��4ا��,��f���#d��%`��W�uҫ���ݑ6]ӗ��AO����օ�f�eK��Khluc#��9�Qӊp%5�f�9F�b��u�t�L����)��tm���]o�)�B�&[��Qa�f#��#�G.��c��ҫ3��e��o�v����ۏ��}���bM�n��M�es�T�T)`���8����L�fCH7E��!�#j$�-)��J��2�_;wgҐG������������ ��H���M�'(懊�C�~��A�,�%��.\Q���!�}�[OTӵ�i�S��*�
�:'�j��u�<gen���5[E.H��{�`��x�����9en��m���������ao'���)X[��u�;�m�7Ԏ�p��w`�2*L�犢�f��;c�q�pAY��R�rb�+��c�p�iw����b��m�s(=:;�&k��ɭ�ѡ�>��4���"�ƫz��5+�`{Ҳ	dWs)����(*$K�R�u�,7\ș}V�r\�mvg[�g�����k!�N�F��n<s��]��Uί��]j����#�4I�����Rǳ���h�O3�Cb�gb���;��P���
�8h�E L��d1Q¢����z���oaU���3��lNh���gxY��P�%s�Xv�)G-t˭X��
B�Ȅu�n��.VԹS���xt7�no.��#l����EϤ��\��Ar3k�l��J��7;20�K]���7�Tǖ�k��;�)Q�or�5h������� 2�pU7XE<I���JonZ�����j�c��|P������m����ǡ�oqP�71v�V�ǔ½�	����4��YA78�'���{{5L� W�(
����-BP�LCI^�:R�
������?<_��ׯǬ��ׯ^�������z����&���(��4?���B�(� ���x�����ףׯ^�z��������������i"6��RC@htc1UJUT!B��gCT��He��HR�ABy�(�<M��j�Z+�4QA�@�+l�4���9䇐5��R%� �Tk@� āT����%<����о,&��S�i�h�Z�a)���!�NH��%o̾@���Jb(M�D���1�hov������\�LPbNT��}>�5bZ$�E䱵�:��Qk��B����>]-����ȵs ���1��la�r�(�K�s����l�=�T�U�}�ٓ@n�mZ��ʶdr�q4V@�^�m�~Fe撘�e�{��[Ċ����v5�*�rY�+��OR���=ّ �cl]K#��v{6cc�:�PܟH�+D_+�l�ÝU�n�i>�y*�}\��fZ�׉wyF�뱸b�N�N�z�Q��d�.Tۘ�D��6����g#H�	�w��O���Tx�Ƕ���Uz2%W�	7�4����s"�<�3;f�jF�k͓�h�/e�ƃx����Ӳ��~��
I�t��� ��wL���T���c�2�����Y���� �`yq�>����\�]J���ͬ����3v�_V���q㢽�7��7�����<���/|^�sm;|$�׵�7{(mÁ�}��]�=�_ ��mqե��H$��[OOgkmm0OL����!�+��͗Ւ3]���AƩ����n����u�-������>�J�ᇖ��(Uʶ�!��v�w�d�S�z�6z��L���~�R���j��<yo�<v�y��hE�+�j�m����q�
� �wҼ4)��ō��	w;���KvN˓�������	��ޯn�;����67�&y�8�=j�X����I�{�Ԃ�g�D!�w�s..��"�n$[6�8ܖ������h�yڹ*��?�)�ɻ�?������wg���wH65Dc<c�6/����b�!���'4���9��>k�����9|跩m��|��9�7)��.��Q�m7��L68�5TZ�sx�}Yk/-Q,�{�=O�}���_Bɮ����ql�2�ɝ�h�&��M���3R�����cCO_G�`c%R;��V�՗�J�ӡ����&���j���5��p�* ���r���V�W����3h�|o�X�m�Y�=[�Ϝ�Qm
R�#ϛor`�F�t��&�oR�R��S�ώ����M��w������֠(��6k�+���d[�V%6#7(����F�f;÷�HK�m2ݏ,��4%탄/_�`�ϫ�~x�Ǒ2k�2yT@PLbw��׮�^U�5��=���
��%)�:f���]y�c��qї]X��N�Ng[��ҏ(p3�y����p���M��k��.	�N0w<Ǒ3��s�U�Ӂ��w%�,�i�����g!Q9L�$ckr��nb�	s�h\e��-�Tsx�.�C�@
lPd��I,8������1��{�6��|K;zڵ�ݪ��
��=eG��{M���_h�6���1�������V�Cm��j��S6�V���+�sT*0������W��m�	�B�����7�|�i���q}���G;*qmk��vOv��!M���o\�=+V2:�����u�N߅uy���®�[t��k����ƅ��-�r�Ҽ�ɺ}�� 5`q��d4c]�4����ʅ>�h��cSP�C.%L��E�°$cgf���B�<��eLr�s�pl�塲�\��,�k۩�mhb�2�L]%ϩ��(j	��e�o�/^J�I��/�RN�7�+��<3�~�[�t�+�k�咕W�{5��fq5B�'��#p��=��(� a}��ey��{9	�zN�mǣ�wt��z*B��L���
�{n�L3�_Yg���d)�lUW�R��k��J�:�f�+���ܗ��i�0No:�$�P��Fu��b$�:`�tۃv^n�f<F<���]}����@���9Mw69������c��ٔ�懝�m�ŭ��B8y���N���3OC�����:�V��S�N�x/lnU�oU��w��[>U7�kǪ�# _D�jYz/�V���D\A]���󱟭TJ�pm6�Jv�^��׷��B�D"�^پ�,�3�ѫ�M��{�͒�D�{{L�wg��l��Ԓ���^�u�\Gu=���m1m�uLnb��|ѱH��-ѕ�Y���G-PW�>m���Y��y�ѡ��=q˳���"��\;j�u�0�ҝ�S��!��R�WB]0�7f���(�~���šR7��������f]��fq*���lϜ6�v�k���ӕ}�n^�H!�&��񃾛�6ۃ�\�}��0������W�S8�_n�z�<�v������v^g��}��-���=������Ect��u��Fn�v.l��1��W�5�xxﳄ����=�슪觨�13t��g��/U�M��W}-p��4���������hl^�����+-ْ���'X��qHF]=��WJ�GN{�ӊ�`\ eQ���E�/ޞk�pw��wj��@��h頹�0�LU�*R�yd�7��J .Y*�������\���u1�fm`铆�|q���ژK��~�����tbg.2���|}�7wݷպL�bٯd3�d�#�5��r1ЅFg7�Y"���E��b�;\4��xc�|(T�c��Җ��13�	[�$ȶ��jԴ�;��qy����#�좠gQgږe�7�S�����p&%0�I�����l�ٶջ��-!�2�\�\G�K3�G<�_a�TCs���2]�Kgu�U��fMLF3�Ï�{��zu%�-W�V?�t�Ws#�ם�U�IO0�5b� �9xy�dS,]j̼��:y����Qz�K%V��v�wj�d�Wo�1嗮�y!���i��9}WS�!�AMh�����]G�^%yh���3sT�!�t�MoV��T���D�J�5��s�]Nq��|�Y�ybMQ�+Ǎ1�#m��|���nvba�s�/`;v��oe����D0,y��}���F<%���b�����
����w6כS�fnY,kʲT���$��aaB�j0�l\ĳ �F��xt7� S��u��d'&8�����������V�Ӭ������c�,�6��g;���n����	X���=�w�#���e:���y��d�)��;{xU�_R5�wm�9YM�Y�έż�c�s����|>�Ӯ��Dg�Ĳ��ңʳ*{��Y���ㆰ��o˸k2lhm�[[�&fL!��.q����v��Գ�aE8�-Ѿ�E�b3}����i�SK��dŘ`�g��fP�@����}m��s��x�]�i�,!ɞ_?Ă2t�gG(����4�^�4�[���D능�����u���[ξ%{�~�{��0���O�T7=�I�:�h���̘�͹�]�o\�*ܶ�\&_H��`���ܓ�o�����8jI�v*��ʠ�L�L���<.o�8Mo\H���Qӊ���g�P��Z�S��\N�^v��&Z߲��j�^|�Ys"��ȵs�}��a��3<�B��ZquTW^u�ƣ�
�;I�E�V3�ms�*k�UL��ʋ�s=��r6�[�}��`���T�\�����
�6�Ϙ�]w%�B��m�,)�Kg֐�@�(b�͝�ko�vT��c�eVyʭ$w���
��'�t�ˏ��1�3-����]��u,P�T���2>�TX�J;���h��2��HV�*c����V*3WV@���N�]�֔�>f4�z�GcH����ssG�/wp]!���v}�2�3)�F��C���%��O����	z/ћ�}X�¡��ʧ�*���2YdpqO�Ů��3꾟�J�^���˖:�'�߹?{4����/OQ�ny�-�B{��3�-��F,�ۼ~`Nr=����J�����.�*4�l.k�+�>'ܾ	U\���f-�m�b��s[�l�t‖�*+v�p0�x���<`�WU��ɽ,�����Q��k�o%��$�Z�EG�s�ڰ�@d���r0����t���*�W��ڝ�=;��c;��-4����R��#(�v�wh�*�z�� �\J<�+b�Sྒྷ�-�4�q� ?i��鏧=�Ս���`�̠{�\X�t
��m�V�/5�(y�>On�*`a\Z�k���;���!��ƺ<�o�2���S�nO��ڸ����ּ�	����>�*�F�CT�:���fzr�F׷-̈́�2m�9Lt:׍��Wg�z�dם�����9�+U����>�8��Y��!r�(�"����)�͆��N����a�ҽ�g�kE���n�����qٽ��n-�p�dAA�	��X�Qj@�5���q.�W4dۛ}mPR3j{kd����׀^kR�s[�}�ᔽ����|������g��\fM���mHdo
�<��,����C���geRi-��0�!�m/(e���|���4�*oE�Zd�:�|��u�;���݋��Xx,��Ȋw���%���Mj*%�Y`I<:Es�>�oK;��zo<��^kC;�]��ߤ��7E�PG�o'���oe�������^R�i+�[㰊��OF��Eǻ���Wo�*c�ߌ�Բ/F�z�����yT�OW���{s�5�`xro%+6�*٨j����0[�y/5� m�'ˎ��v�t5n�H'đ���C9j��]oI휵`-�Jk��ܞa���Zn+:��kN��a�'��o�ȍ��rM;���]��oܫ#/��6e���i��m��E �n\�}��nQ�;�\��J#Ҳ�Nje)nҦ���]�4�f�_l����m�6��Dn��m�r�}W"2�2����"�M�]�٧���=����gl^�9�+�7Q�l�3�a�'$m8���{��\�����V7�^|�~]}���k��׏�^��*�����=�rǊȑp���á��=w�7�.=�NL�ֳ���]��r��|}1��;��K�8��L.�Q��}V�v�����{��Mه�SҦ"�&���){�Gc�Y}���c��|���M�/k��Y|�6-<����=�$;ڍd|)^��=�}~�;���hkHn��o����ޓ+'�6v�29��hD�-�6/��v����m��a��zo�\W��C��O{�ؚ��Lw$m�$��s�K<�+��@e��VhUn��h��5�_.��b{�[�X�#!�(���x����B誽�桜�O�&y��dN�sU^�Y���̢��Qms]M,'��N���0��G��V�4?	���iWB��Uʮ�*fq���d�=.u��u/l�ϛ�c�b�4E��B}C�8��9\OD���N��w2[U�y�,�܅SS�7�7���!�S7��	��jGn�d��ս}輘�{���(e;�;X!���P����^l��q��2�,F�zgגə�̺�#��.����]".w&B�W��J��n��y@����ޱ�G�^�ت�-�Q�^Ի#bB�^�7 �Җ�7���݈�3C/R�1��RgN�}�S�7��~��Zr������,����U�g`ŝ���gD�V��~�Ýg���?s���s9�Z����^������tʘ?��:q/�gU�ڝO-��"�O|�Uv�o{}'���_H�,7)���ڷ}#S�|�ܳ��*=�.��w��K��ϻ���W��������/=ѹ�̟v�mKem��1�״�w�ݘ�2)�t	�����9�z;���U�<fE���GY���=���H�b�;9q�_sC��^]�u�����_s���yZ�k����������;u�Wu�c||	4<fk�9�,C��R\ջ��)% f0�ީ��ic�Y�.�S��Ds�y��x�\w��r&=�.a�;��p�2 H�p%w�۽��Նx՜6�*7|{.���gM�ʟdk�\���h�g�}�Ƈ��6�-dL� 8r'7!�CDǞEbj�QZ�6ֺ������1�i�
k��V�Е�p��gMo����t�Q�(���� QQ����D�(�'�� "���1�����PS2�L*��°�2�� C*��0�@�0� C ʰ°�2�+�*�(ʰʰ°�0��C ʰ0�C �2�0� C �2� C*��0��++ C
�ʰ�2�0� C*� �2�0� °2�0�2� C�0 �0��C*��2�0� 2�2�2�0�+�C
� C �0� C �2�2�2����>x�C
�*�(ʰʰʰ�0!�*�*��2�2�0,2�C*�¾Xa �Q�U�!�a�eXeX@� !�a�aVV@�@!�``@�!�d08aVV@��a�` ��U� !�a���"��0�0Ș�������"� � ��"� � ��(��3��9 @ @P@P��< � �aa@`P	��@!�@&�Di�@&�Aa2� �0L�4ʨL �2�(�10���L*�0"M0��0�9����
�2�LL*$0�2�3L�C*�¤2�4ʻ	�!�d�W�+ C(°ʾy�x C*�ʰʰʰ�0� C*�U� !�aV �U�@!�e�W��`���O�UQ�TdE��|���������fx�p~?3������!���2|�s�J��~]��a�<AQ^��<�������e�"�+B�~~���D$�����ԇ�"�+��x���Y(��1�MC���'� ���!���+���i fD �P �Pd�ID\� 0 � BȀ�(  @� �  H2� H�" H 
� B  B�*B�H��*��� J���) @�ʰB �(���,?������D�Z ��H��@�P (8��w�g.!J��.���qETV��P�ۡq����O=�P/��C۔���􈪊��C�����?�?dTW�Q_:��8�Qo�;G�UE~����?����~�|n
��+��s�ܭ����DUEi�}G4>���"�+�;H��T��g|���о`v������y�DUEa����~�ETW�03�e(�^��c��e>ꇙ����ɜ����DUE}O�_��� ��ߴ�c+�T�� *��7h�.
�֟͛����S�����)���^�����0(���1!-�'��D)$� 0&��J�$	R�%R��SL�Em��6h� �"P�CmJm@���
H�B�b%UJ$��띌�Uj���s����q�ضݎE��ZegN�skmk27mWBm���6h#f���Pٽ9���j6�f'Nꕫ���-[Mk���̶��S������m6�mmL�髦��VkJ�n�v]�ګ�v�m�]��c!�l��]]U3��ӝ�u�:�묻V�-K���m�����KJ�[m���ԧe�fZiY��<  '��E���j�� ����V���l�j�[�o<�k�m=ѵ\�m�B�ٝ����`�7=��Ҭ�n�Hj�h�+M˽�t�7]�-i���\T�k���  �nB��DHQ!{ﾯ��BE	�k$/�7$(턎��P�Y��잮�[+lz��OM�m�ys�U[l�����ziVղgSA�ج=����2�s��mM[T��5��k����\��J����  ��P�jZ﻽[j�i�7���ͦ���P���^�%r��6��S*�q� U)�R���TҕD�s���m6ڢek`K)��
*��n�KUW[�Y��  �R�e-tqҭ��ɀP�}�v���W<\��t`)"�i��@
�aU=��󠦕VO84 ��ze�i�z��w]ǰ��6f�   ;}�ـkY�q���N��U��֨�	ńQW'��GM*�(�۳@(��p
]�A)�L��M���!W2��us�؏�  6�$5�����(���;5Puo{�W����X��QWk^�UD��f��PUPlz⊪���Pq�9�n�[I��mej�l���;��  ��eB�:��:
]z� u{�  �w��  CL( s�@{K� [��t ���  �י�w�V���m���v>  ��  7��� ���( .'p Cv�`  n;8@ݭ� �Kܻ� �w4�@���  mڻ;��e�i�֙�T�m��4� o{�  /;��  7[� V�]�  �x�� j0� �[p  ��� ���� ���  ��ѳ��c���u��3Lm�]�|  F�  ���  ok�  ��  :�x  twu� �����  ��N�*�0 [��  |"��JR�@@��a%%J&@ �{L���Q�@  �~%)S@  � ʕ)�#@��H����@��K��Oӿ/����ӿE�Mfٔt���喭b �62v��-J�����諭�����ϝ���mZ���m�����jֶ���խm��[V��mV�mm}�����|O��	��!�Wj��L�P^�'��*�X�&r�*�f�z![%`��V��4�9��b)[PY��5��+)]�M�X�Y(�l5�����zrM���_G�w{F!����&�v*f<����ռ:ӽm���c���u�43�����FV4V��yMU�Z��� u��^۰��i�/��B���6�kF�ѠZTe�	�z%�e�SP��7B��@]L�:���2���������?��rdP���OAGTCFE��M�Ii��!$�������eԺ[f�X~'��ɸ�7�˸��5,�@�B\���ܡ�v�U�U�������Q�T6�s2Z�(wN)�++u�ٷF,�3t�7��k�~�6�ӵ1�1S�D�j�e�&�up8_�d�
�>\����Y��Q�z��ED��t�j�lE2C����\�wf��!̚�f�Yb�V�]�(�Kw��V-�0���X+T��ݔ����\^����n�3��Tuu�gB�0�*TňR�1��b�3�R�*cY^�a�e��l����٬��M"��P^�-R�3WX0jVR!Y��!�&B�
@[�>��cN㭂ŷ�X���E@e����5[�j��ҥ��l�N���4t�WX���D1lќ�dz���H�c�:g<J#Q;*-'n�m#u�j��MP в�b��@�RbAf�
�L���ˑ��P��z�ؕ)��S�L�ׁ��![��o]���K���������0Cei����W��2���W�{j"�U��91Z3 �coj�Z)�����^e�6�f㶕�,��ű��*��{*ҠM�טΈi�7�X	�YKN�Ԓ'f�Q6C7nmCX
/c���mb��׮,���(`WQ�AUӭh[���Rܽ��kU��8m�j?����nf���jb�@����|�C�AW�-���TA��*�$nC�7���U�V���G+v�ZRV����� yE��N7aͬG6��$�ڶ¨�Lɘ3ES���l��[n��7de�S)k�V=twpEl�@�7�cHHF@�A�����A��Jm��wp�*�1��5l�k�cØ��W֣XV[���f��C[ucm](��0��Ǘ����m'`��B����Օ ��������1JĀ���t�켻X ��t��\�m%dW3
�YB���z�K���L�t�T�:앹�V!n$p�Э���[��!��E�]:Po�ڼ���k.�-DQ�[�p-�DiS
�Z"�K��їY0� ܭ�F��� qP ͸{�}�tcQ�.39�a]�C�����rX��6�kyFf�N7W1Q����>�홒L�'@��`qB��y �X��6�`ei3t;�&Q�I��ɛn��!ѩKi)��ʛf�҉��Ӄ��	�iP��o��<�x�x��&�V�i-��J*4�e�b�����TPF��D�f&w~@LQ������2Э�[n�G.��Yx��5R�*-��Ĳee�f����Af����aB6���[���]��l���U�PZ�U�����È�����R�Aw���1�f@�fi���#z]�Й��i��!ے�3�h�olV8mРh�x�=�pT�k��۲�=��̓%'ʆP:�����QjZ�f:�hU�ynX�hnSbFQg�D6�q�j�*��b܁��.�
��=D���B"ek���]*©[�n�w��7aIh4#��j�2毂*� ��&%��)��;�1�m �R*��^*TSw%@�e�9�S��EcīM��(�[K�A���*U��14�k�Baz� -�#��DssJ�۫t��à��V��lJ��Дբ2K����ʃdZ�Z[Yq�jڋ!s��W)} ���buJ�)\c�NݺAvZ�SU�V�Ӱm��ݩ2'&�A5�pm�HZ8�,�Ouv%�^Z��&�6� ���l<Į��XQA�!o#Fҽv�jQJ�יK[�j�.�ol�t�����v�D׀1Pۻ	f��2��^݂�9Cvj�t>��k�ۭ�*�j�75X�Z(mr���LY�hm:��g#�,��T	�,:aݫ{$���������"�-������%�:�ə@�ݱqBqմڋ��κ�7-�M`ֵDF0��Dل��ylb���Ģ����6��K[�yZ1�%�*���|R�6"��.�(���٣�̂�.a���&�ӆG,4�H3��Z&�`ʺ)�w��ȣ���c\;0�U�J,F�̥��4�U�Yxjӡa|)�sa��=�N�Jw
-b�v��t��ƙW�Ac��5i��E�e�yl��}�FE����=	�I.ۥ�jC�Rl=Ru)�J�	���s	�7�鉑��ĥ�3C*D�,̺Af]O�AX��y�ᵔjȿ�&�ˊɭT�.���$Y�Ŕ��IJ��AUd:�uj��V7j��D*��:n�6(ћ"����cp]A �v��p�Nж�疑�ʑ\��Ly,@�@%�{[(^�ElIVҕ�n�rSVi�l-7%$*����vHY	Zd��u$f[T��Z���p�m�e�e�2�S's]�b�:(�Zc4��BLU��gţPa	�����ʴ�%W�J��=b�䄲��s�P)���,�C;Vp�5�q����qjG�7F�dR�m%,�
;J��C]*�]�G+If�9��Hf�u'V䴨�Ȓ�q���K�2�S�n�c�ϬZOkm
cT�7Pƞ#L rV`�O!+��Kr��jm=�����(���a�1()�X������ӷh�
�צ=��T�L��*�F�u7q ER����w�hQꖝ�v�(
x�pVB��ۺşC�-�oX�/t3EG�Y��@w2�3oq�I9D��!d�*lR�h\���m|�������j��]����ʀ!n�� u��X�nf�������n�kL=Tެ�&<�X�<��"��z2c����� �cɆ�	H�,�K ��-�YRֆ��$�鳭���s
��Yv2ܨ޼�Ec�V�$�ńIuy���j<@+���;oK�6��AA2X�X�+\�]"���Y�w{�M��z�ӆ֘����,�TC�r:/V�j��E���B�z���/���cl�LT�j�S&2��M�#��^g̍��9�+�܍�;h��#S�2�fI��Y �4���Ę6��X�
���?@��&V� ��6v��)#�L��\�Z������ca����-���]\vt�j����#C�!pLܠAh�����O�˂���V�j�e�9@�L|t'���w�X����QN`�u!ޜL����ݏ��f���b<��䬆l(��@W��*nk�쎌-l�m;�!�Uy��F�ЦCjV��cmі�:ʎ����w��I#�����ݗa<�̈����@;��ջ���^c4��g3Iy4C���ՙwx
�"Q� 3B!�%�m�X�����i�xj��]:�dqȯLZ�^(����'^f��I��	��JN�Ve�&�/���53&�/�2�1�N��:�^��ATͫU	,0�v��[,��L�j�`Tհ��إ�l�2�"^eM�����K�Zu^"T5��y��Á]��D��h����-����r�r�=b�Ȕ�R��T���f�6V�5�SK��>lлŬ���QC4�mńPh๐'�V��/�� n�Y�Ed�խ�&ѶJ��պ6�K�Z2��m�j���ZQWB��껰×M1�x�h��w7aQGG��4'YvZ���ww�� &�]�Gd�D��9� �{@&-�Wz*[;j���2��V��(�0��K�v9v]:��RqI�-	5�][� 1��yNA�N���^J͘�]7"��I�h�B��n�v�,e���-M�a׍����V&���⦜������"[�jj���kv4�#i�ٰM��lR��8��u����I6)�;�H]J�ʤ.Z��VJ�X�g�
���^�9��B%����BQ#-�E��\�4��a�S�ݦl)���H֒j:b�B���� �.�^Ayl!�H�j��G���X��ct[�y�Jx؆�n��h(r�/Y��
��$�f�x�Q��N�X��4�R=��
:�3j�
SdL�jv�eԠ
'eYV����<��P��7`�k�����SU-m��`�����Jۦ��0e"NH�cۣȐ�h�V�Ƿ�� ��崭��0SYNb(������/*�`�Z�e	��TiV*]ù�,za嚂dقP!�X�)����YA�G3Tst����1��2Q�_����ɊE��vB�p!գ���� ���/dS�����Z ��&"�ICf I
�[w�Yө�r*��j=ț�ϓ�8���2�{[��4�]�c�wL�S�4iۺu	G�ܹ1?��kt��@<[���+���PJ�K3pd&eL�R�l���3P"�����(�d��G���ԳsGG#���,���-#�-`����̦,֠�����Y��ecЁ�u4��/L-9m�d���$�sM�/wG�*&h`�ȱ�x�[y0]�J�ɷ���Pʸ�j��R�73E�#�� ![�ܦ�76C���kaۻ�J+V8쪼��.��ò��Y4�M��\���x�r8ր�6j��xjhU�j��v�-\�	N�]H��(�ͧp����|ڷH=����Y�V�l�{�]ӖVc�nn�J���)"+���n-�t�j�IH��h{��k�=`lHZو��إh���u�)�bzV ��m+Z敮4�t���!Kg�E|�轇�@�zX���(�k0�ֲa�bS�s]m �k��x˩)1�`7��fj4�4���TV��w	Wl}6��)	�meR!=ۆ�i�M��mF��@��5=LС���X[լРi*��ص�(���R� �HtV3�2]�[ڬ[p�M�pJ�/eae^�6¶@�ʈP/F��sC�`=A2-<gw"�K7�Vb�<Q|E'KPd�];a.S�3q'sXUoj�M�xݽ���i]�Æ%5:ܢKͤ��*ޠ�;��Ub�V���-�+mÖ�M�S��l��Gk"n������B��;u"����54l��ݖF=s�M���W��`�+\y�I6+�� �l9��*�����{��/ `���b�Rʫn"��[�$p�q<Y��ѩRn[�n^6֓bІ⦝� � �e��IWL��ge
������M�x�����h��h�o3)��sm�M��A����R
q�zFFb�i�K)�����mD�-*�t���ж�@f�/kF%e&ߴQP*+TX�����3m�/[I���\�B��Cʊ�\��j�T�Hҍ�^�fl���rܲ�S�T6o�ա��ZjC��t��{Jn��w+5������M&��:e�pFi�5ٻ =�����ȥ�Jk�	w�S
_bb�Ȩ�]��ז)Ռ���E�'V6!��e�� ��,�?l�%:4�V;}-����yucɥE�Б-|Q.в�������vX���Օ,��m���R�i�Y��i�Vn�4�T�d��杠��邠���*�^AxTOl�cIʴ%A3�yfT���ˈ�7j���J�z��]m�(�c�:�{���e�l2�*ݫ���`
��-c)dm,캳\pV���ٻ�_�]2,�$�oiq˄��ƶ�P�c�wf��8C�E+�yGѷo2� �2Z!E�֩��.	j�Ԫ�$]+t���l^Ȓpӽ�A�������3(Y2ᩌ���rF5jj���I��i����6�Ћ�^Pz0+F�,�"���3t<r�I�f��L Ѡ�5��`:
�T̸C���b�I�m�{����/7Zø������)��N ��v��	r(���-�0�$�'5�X�Q�d;۫��ݍ���)��J�o0V
�2O*
Wt2]t�llʆ+�S�I�;��;Ztx�׋&�H��4�����V��W��8��hVF4�hACi�Zڰ˭$�(`5pS�DV(h.��
�o*��n ZFII�7Zbu�k4��MT�r,��t��Yq�Y�����K��8�U�÷��]B���
Z^��z�ts�r��IRb����XslZ��n�ԏa�,�XW�AjR��3(�5��4�MR��Սf7f�@R�5��P�B�Cp+\PT��YPĝ
Y�X �h����z��ohQy��ߔ��lQi:�N��4���ۉ� _kn��:����Ea����
�Z��w&�-�Zfd�l�?Lsv�VC���W �r;20�7�X�ԉk�����M�iud�9�)e&�4*�M`otWx�l�,veX�(f5@��6b���T�����w���)���Z։,|���e;`��f�v1���2��S�j��*���׬%��$�&=4]*�ݺ��虗oi �'�$�7$k1KҎ�V~����H�^�J�aԭ=Bm�u�6��X��ъ`�j5< �G"y�w��ڭ�5��D5`�an,ek0��嫱��	n�^�4�������M���G�~J]�d��/#Um�Dhmڻh�Ö���֠2����hI�2�1�Ze�4-R�-�t�m�V���J��yfi�v[GI]�e� �ԴjH��2����²��=lc�e&���;&�VdE��)�驥=t�&,�PEi -�^�R�xI�(+r�ռW�M��� �c�M�GI�З�T%]$�	m�� .�d��t�;��\%~t:��>����)R#��jrW�������QBg���J[��{��pzZȗX�3��Bs�H1O�s&@��g���P��e��+�ŷ�iH�	�h/%O�)UNj))e5�k���7;e�fK�J�g-qn��u�4�"�<��yw��q��Ӄ��X��;,�sHU�W$�U�y������-S���78�n�:�o����!_I�s��{�6IH�;�;�;�O]�S���,}��w5��~�.�*�U,2�z_KYcm���vu1'YoJ��Z�T��z�(*����X��UUj(2�%�sc�~nLz�o��_Jgf`ŏ��\�.U��=�ۥ������w
���̫�u�p�+�Xڻ1�R� Z�ݾ�\Z��f�L�-�MdZ�ff���M�/�-��i�:�r�b���l=��7���o	ܞ�7�)�č��OG<��}N�%�봡wu��<�5��m�\hJ��^L��hG�9�,�W^�/eo��Z�y�ʟ+Η@�O3ٻ�-I������Ek�^�o�`��\���G��`���\�tGv�;��^}�Y�e�<�Ю�_��8*R���.�h����^����������r^vP�l�����D�E�.��aW ���]6d�p��/��t�0F+X�V��s���-�31�h�MJ�v��J�a�����v�	4;��CY��u�����w�#wqN�����I.�l��/�[?L�X�[��ZF��SGZ�+O��޺O,wT9|��LMG��[
�����V�2�d�:�`0�{����4})WpaN�Vf�3r��!�����%{�]��E�`��euʓ'-��5�0������-��v���9;��^��[�N����)�gfu�q@�
vV^J���r��Z�@�^����i��7qȮ�1�%>�7,`��B1l�L�M��ס��u%6
[@�ạ� ��5)�|�ј��.�X�iȰ�a�/B݁��儁�r)���8]�;�&^��7ċ�A��Jo�C�ؽ��CfG(d�E���fʨx���8�tWz�ua�w>[��4�W��K���d��En݀����b�
k!�{��k� #�b�ˎ�c#9�UB��I٢��*��#��r�ر�;���mX{-=J��t����+f�Ћm���Pf�Ϙ�k]i��L���1$�g
�[@�\���8٭|by'v}ݳ��Q}m��j��OtR����m��!I��:��Ѓ�b����Pb�d����XX�{�|F;�,�鴗xd���NL���i}��f��Jx�,�y���f]*7�G�c�3M5���T�x7!�m��k(�ܦ�i�3&�����0��j[!��B�-X|�ix)Ve�t�Nmѭ��R��Ё��}�2��晳�y�% /��-߄�mha;�u�ޭp�Vulk,1�z��5���ζGsL��f�S�J��Ւ�ۺ���)h`�5�s`lJ��F�{x���!,M�8�5|uݽLlѲ.w��<w)�a�ڲ���Ұ���ѧ{���]ԣ�Ш���#/�[Z�:�17KKᆉþh�O0y���v��GLQ�V��8`���S���;q�Wi,���r��L��o�^��e��S�b��,�Kޚo��aV�;G����ު����V�ӳG���ᯖ�V���;���@+��5{5��
������A�x��iQ��T�.��,J"���9KDsH���6���'*#�:Z�M#6k�F��6�3st�+w8���kK�R˱�E���(�\�ҏr��^>��%���U�)�XH�t��1
�
����]�M�\i-�H���#���7��a��e'�n�E;^v�(Q���\������_�����4	��ߛu7���@cCA�d�q��p��5��[�o���;��UVF[�۰���WrY��vOs�b��5
�wOpG�s��V��Y/��V������<7w1�7���	�acE�N䵗���سVړ�Eo�w�^.�E3VYk#﷐{�Z��Z�ti��?��o��kR"M�@��f�H�T��H;����%n�a8Z�2Z,+����n+�Y�/I�{�0*���.��ݲz�NK�r�Nz񢵽~7�'5����DR�8�X�R\��wPެ3���s}�W{E8v��}ձ�X6c�t.�7�G��oٯ���}�|HV�i�o�;c,*�A��3s����d���ɳ�����#iW/�� ��j�m���W�_� p!}��l����Q�ֲ��Ktv�8�����x���4��UnJ�R����;j���ݺܰ�+U���+��:F�,ܲ�	�*�s�㫗�Н�6av�Z�G�����@�V^��PZ�1������ՠ3�ؾ�]���Ȩo��M��B�er��[-ZI�aw<���(]-��daq��4��Uh�&��S��B����).��-���x.�:]؛�8�I���'���ȸU�Z��9hD;q&�ޜn��F��.��F�E�;}�%_`J���u���������m����7�{/ryݱ�y�,m]��]vx9Ԁt|�N��fMZ����P���Ӛհgn���k�7���Y�s3,9���A�s�s��{xZ�o"ݎq�Fo�y��TT9\ò��Zd�wU�	֠$��+���*�����B�uv;�j�b=˔�>ٌ���������i|F��A�hbP���.�ѹY7Uk�6/f���	Z����7U��ڠ��O������U�6}�4ۗ�/<�-ۺ<Y�oq�(9ou���`Ƚ��B���^vU ��[�Ӊ�/>N��vr��Y�K�7`��R��ü��[�5����t�v��/| Kղ�"_Z�x����SX�n�q50��p�5:ck�h̅�mCc�F"WY0h�5�]v��� ��_`��6�Lŏ��X[ �[�ȡ��u��]:Cjw#B����r�L��/�y�p�m%�{^1ܯ2���k������>p<uP��P��e�;��c ^d��e��1�qő��i؋�H)��:�3�{�l���V�OJb�z�nS�eѲۚB�kuM	�3�jݑ�8n�*tp�ݵ׌�ҁ���>��vVH:>3,�Y{���a��xw\-a��d��[���Ɠm\Kk����MW��('qb�o^��NQt� ���3H��ҿ�u�y1-X����cX�;���y��V�]���/R��Ӝ��0E5wQ#��\t؟U�ܘ�B�"�[��*�� ��0:��9���o��Ά;�S�G�9����ԹɎ��4)�8�x֙�{�un�+�Z�wqPLCD~玾�w�{��F3fGVv�[y�V\OS����M{���`�0��kM�I&��z��O�i0��\B��ٯ|��	V��fi�9�{֜�Cb��bay`���x��3��;�.{�>��i:S0µ��@�>�A����^�o�7=��ʓ);\N�
�5��]�%L֣Q\�.�T;ۗc+��ŕl���m룡w����2ǌPo��`�I�A'�{��N��������P5�	�ە���Jw@�np�t��KvbZCz��jXW\+�v l�ʤ�-e[{��˩���dkC$Q���鳝��������z�:q^ 
, S��X�1f�{MA$nI�q ݫ|�y63�X���G��|_1J���aG�՘���.��8�1R�^ކ�T�m�WZ�w����R�˳@YX�m��/\��2�m:4�QgK`	Ƭ@k�/�c�C�I_w!�����wt���۟YX�Zz�3Y�,��]��w.���\�=*�|�f�E@Pt���)iY:p�Y����=�h���P.Qz�S(��^d�3��Ú��}j���Jm���W��/U$0��SkU��gL�3NJ�"�Pɗs�7�~�f�����w���W���Kܤ�l�r��K�&�Wc0�,�ַ������E�--�L��jt���m:��N��fW�)��9+��A�x�J¦q�l
Z��-k�VZnY�o\�'\/C�D��9V�Z̭�<o;1��v�� �Q:l�R�je���f�n��_�o�t%��ԳgfF+��N��J���K��_���2B��a7i�k��V�-���%oJt�0�:���C++����n�����b��2,�pu��'c�d��P,hxY�Рu�v��r��9�)|MMG (q����`�nԺ�H�E,�6������b�aw]m�a,ȵuj ���
�2�)�F���Y�+B"���w�rS�Z��W]�<i��h�c���IW�v�y�N�T��Ҧ�i����4�u�YW�Sܷoq-W��vÕ��Z����Js�U��ba��ҹw��hG ;4K���A:�gc0��[�,��I1{�z�ܥ�㵨9�m5{�1^,iZ帥�jeD\�}[�ى�P/�Y6�K&�M\���x"�{���	ME;y���F��F�a�od'i��bQ�����"�MK���VqO%�S2bW����v��N7�w	����\.E�:����'���'�}����y՞�8�V0�0����Z���;�η���Ykc�ې�ٙ�bK����6l,��.U�mX�{ʹ����^Ҙ����B>4�Nz�#{}�J�v�]��拮k�=���K�}�Lw:
����fy�BO98�{)Ǹ1z�שּׂ9G"��%+���x��
gJ��sΏp�ɝ������ݦ�N�14˵�VL�K�f��7`��Uep�.>���EUa�0�PI�:Z�a�8c@�d��9(n_E˥A��0-�Kֻc҅4��wj�[�NI�.���#fݜ����O\|z�!�T�ͫy��E;��NwX����`��O�m8)�pޭ�6���#5�e&�w�h{Jj�jW��E����:�u�mK�l[]|5�A*�r��*���/�-wTؠv�4Y��]D-�<����w&��G�ͤ�=�������ᖔ�5d�7�.R���I01�bQ�e�n�¨��3�j�tw ё0���,z��yT٦�܄?+W�o!�؀Y{��0yl2n�o�-�v�����	^�b��h���I��5 �aWهP�:_�o	���D8��RN�A��vm)�wF�J1�b�3��E��H��Lg�Zb�8z��·���%ܝ��A�G_]������hR�j�K��(愋���N+6���E7I-ܽ7,�c���9�W{�5`�$�S&��~���W�Z�К#�@ۡ��p�[��R��o!��62�����B��W}����s<n_f@8rɣ�������/�l�����@�؂@�6�L�����hW>P�j�w����^�]���q�"�D��Ň6���Y!H�`]؏�Y]e��.a��GYW��1u�Yeu��":H���/K����^�����c<����'dDS��6�Uݯ�bn]�PQ���mg�]G���a�ǻ}�k�]�W�{�A����3BԺ�;|ݷ
�NG�n_�x���5�=�:�V�����\��ss�(��!���xFG2h�l5\�X���/CڵV�X� 뼃�r���g��T�b��V��u�,��PG���7"��G����c8�3	�}8	��ٳ&�aE��#$Z�ݝf�*�?02L�V �a3�0=K�$��EC��17���2r�_���� �MG.���(�i�L��W���'��iq���m�(������2�ܸ������,hso/J���[`]��gG��Wl�>�=�oqTC���<n<�����ۮ���X�
=KP=w����h�wǝB.Q��5[+ݤ4�3����f��N��n(}�םVh�9���3r��wx��D��L���x�]��4��i�{��uVrIVs�P��^. I⫬(��ൕUȔ�z˴��^�+�C4Rч��#�k�q� �4�x�x��ǝ�m[L�kx���R}���E�֠��8\&X�Փ:ù�B.�p�R���C㽔�ON��<�}Z�Ct�	Ƚ�]M��r�Nx-�;7q��W� �qt�:��b���E�C�7P��y��+?ey�
��J0��jᚴ�ﱦ�U��%F�me6z��Iצ��ny�����S�x֗����9�u��{�!���繙�駘J^Q<m��Igq��V0VB�'�꘸iY��jC� k�Ub���Ğe�7Af波C���Z4ƷƧ븏E�⦮`��h4�K�ɻJ�ё�|k Rތ=.�wՕ�'�w��YnU���W:ˤ���Ѡ-k:�ĸ����j�D&ٞf��q|��g.���Õ����`}�5da��;b�B�ߩ���#,X׀�F<Y�Ʊ�b�v)��I1Z5�ꡮ#��c.��,r521,�.���Lы{�L�l���Y��.�fus�1����u潔�OEV]��\��8�6J�qQFt��_�������op6���3Z�����8"�+�;m�ں�&$f��
�Jn��`]��o�(��o��Sm�^�4v�"�ʉ���8�r���C�J��\�fͪF�N���jA4�V�D� J�[�uN�tu���:�h���	�Wgot����)IP�	�Xgh�"_AG���v�Yϛ�z���x{]�1{G��Y�}8�;��J7&Y�҂���6�b��N�W��L_N���j]�Dch):���'  ���uG}ȕ����qٴ�V�\J�
���9K�3���u�M	ǀ����u��/��xS8ĳ의�)�$�.�p�Ĥ��I�2{�K�%@�v1[�����U{������ڭ�����֭km�����}�?����wW�����8Gr�Z@�K{�3F ��x�bij�ܒ¤�(�6q_I� 3F�O���N[�{�3��"`*���m<|�M{V�n#�%�p���`H�_�ݛ��}�m�-ob��5��l�yDx"�˭O���.�����LO�H����^�y��P�������n�xυ�5�&�pd����:��NQ
�bECD�)'l�����{(��U\����xUK�l*n�^v�p�Y�T%�T����MD��ILz��+�2{ ʴ%8g]�k��� �Μ2��eV��h�bMU��ڔ�uFu�ì:';t���F�(j [�z3v���T�7zұxb���7��i�w	STk�@OŒs�\�R�9J�>Õ�;	��L���O��{��v%�k9巯x3���9t3�A`�R�e��6�caՍ�Q�ɼV��v�/�����z��A*�"�]D�a�f$��K�N�D��:L�Y���6dC��1�-�gLK�Hգu��tOX|�93��]��m���8_hֶ���0 p� [cc�.�n�{8��h�}{B[�t��Z��3X�<��L~��'sۛ�E�ݾɊ�	�{M�a�V���KH,�vѫ�|�T�%�BBۻ��Y-Iǳ5{F�ڰlF��޶���i�m�p�3)CJ�_l�Ϻ�$F92?,��J�8W9�A�t����:=��U]��i�:Yp�b�GrA\Ox4����wx��-�ix�6�(Je�W�rR_ �A�<TՔ�s�,̵ʥ%v"�̗6���2u��Rl�h�|���<F×���u�|�k(Y�K�w%���˩7�n��M=�.�'o;y��o��!1:�3��t�se�_-�b��J�g
B�r��C�.���*ӻUy&%g;ә���s�� НDU�=Vn�P�����(�臷Wڬ�Aݵ/C�QU:�Q�0`��ek�aK �AR�g��Q���*l�]��ס�J8��˪�{lm����Bs��vb����셋��Vf�}�}{�D[.��d<$�>�'@��b�a`n�N�b!u̗�1�y���.��N��V�w�]�+���Yyd�Y��(�/i.h�X�D��t�t��I�/\��+ɈcTv�F�*$����\wEVg���P�k�"���SX:�&F�|���u�O0J���{�+G��js���<�O�j�J{ޚc� �%7˲��e��T�x��/K�e,�ev�.���Z�т�\�ie=���_NË5)�"���}�l]���{X��fK(X!r"���g�d�<�c��צto^ �sk��9�H�.��!�1�G3�7�*1�����z�(���3x���1+-^�+%��]{z��*���s��'#�F��A.�D�m�(p�}&����˹����C\�Bhx��U��N��d��+E�+�n�s-I�+ٳ�Sʊ5"�nQnp��k ���`˧�����J��=0)IM�%�W��_C��&���Y5�_>%�&�X�n����F�E�WU+�B�٘�E8n+���\�;�o!�`��zjQ�-e�t�fw�[ý���ܙ�Q�پ��v=���Ў���1���A�� s[k-���uxS�m1`ʾA#(ۛw����7q٥N4�^m��u����Z�6Lw�^y�^Լ�h���mM1�
���JN����w
p QW��m�еB�<�����Ze���r�N��fG�H�\���Ak�wWnb��i`� QZ��]�-&Os��J,�V{x'�v�JP��y�QqZܵΔ���pk���<l4���7&QŔ�_B��1���!�.��V����>��6�����.opC�i�����_c$ �{�`ZSg�H�:s�ޜ�zifݓK��e]�m�#����v��6�5�e��-@�f�%)�;��#ZD�\*�܍�#�q��S�S� �-2���n�ɴ��읔��|N�9� �Bld��B�teYs��K�s}'�t}�R7y�t$yu=��ԇ>wk��ȷ���,5�W�akt�8G�ԴH�vh�
��γp�i% ��K��iMՂ��
}B�Ш�T��2��]!]�vS*�K̮U��0��C�xr%NW��!�,l��x-��#��>O-��,{s��'i��,�7����iC���1���x����ծ��f��q����>h�㥦���v��k�8���V2���%�i|ظ(j��^<�T�(]r��摆^�33"UA�O�,0��rG��w�Et6im��a����þ:8��)i��f�gd�v��ჾ�ѝ��w%qv\>�_g�y'���ҌH�X�C��&ѮH�x�7J5�۰�����u����s�B���V�`�38�?�m^,V�^��@V=�uv�Vɴn�Y�T��Z6�w�h�N���X��PG�\R*���3P6������l���M���v��]N�]1l�͢�|�Q}(���4@1�%fe�ѣqPt��ӊF�Ea2��fK� 쌚���!�*��Խx�y	�	���/J(��V��?'2Q�����fuBTv��+��u�-��*<9��E�6�t��M�Ĩn�o��S���(��xKQZg]���~ف���F����r̀R��Z��yP�\�m�'^��|{�E��e`�eӼk%��y��k@s*X��v�j�����;��BoQ��qۮ����s��v�ȴz�V3���椏+�af�o*&]��hT��[B��zvs��ٺ���nv��q��h4
8F�r�t�v����6�w�Y�p33�Ol�(�Jl��}Z�YgX���л:v�.� y��w����yx��{zc~��d�l��7q�)ժF�a�o�_�#q�N��\�G��)���C�}z�3e/�Ja�:w'��k��Wx8���f���ZL�R#����2�%)�!��f�(���Ԗd���w�7�*�2�B�2CJu:V��|��i������ۮ�~�R�����g��3��w:�͡��#)�bB덍צu�E�
��X�:�wۥ�Nd��̤:��{4>tӹ�Q�@	`�X����+��kRV芹�bOAR`�XdT�ˉ���B�E�G�i[��9���3�����k&��#���Cz�u5i�c�Ac�/���;���G�T�KYh�l (�tt�"�qZ����5zI����(k�B�α��dѷ+���T�V�B_��,��� ��N.#9�*㙇�w��r���'���i<�������e)�̮�w�F�NDq�tA��&M��Wⶍ��s��ʷ���&�E������O��sKh�Q��m�e�Q?I'�K�)��³��O^j�gj�S��ud:�����m������V�f�W�:���̬�g}3'.�n��Q?C]�I:�f˺�+��1�G�|�Z^�@n���'���A��;�s����-�w/i@Rzۜ���Q���Frin�`~��g�rzQ�I������%=Ԛi�����-�� 9dҬ��ve��շt����hva�
r�����A��3:�[��+w��r�=�����P��uk��&�ׁ��p���I�,)n����˳��r�[�5�&x���,2+J��"�z�F�[4kLJWu�d]�Luv��j|��7��k�]'tfÂ]*ʇ���oh���K��ދ�>�#8P�ȶ��Z�p�����j�uػ
�d��\��
Q�t��3E������).{o7+X����v��	%b�(��S�+~�u-L�]4d�h�l�!��*���4�^t�[0_��-��8~A�p�k�YLP\-�Ǫ`���9��H��J�����5���O6
�>��gIQ�η��WZL	�fE9�"��<��)��W�GpM��Y� ��h����;���Zہd'�u
ѫ0{2��J����2��q�%���#�ե��p��=���C)��"eԂ����}�q���[˨�ƈ-+�������bu�A�gV���2�VH3�U'�p(�xYVv�؋#m�գ+v�%����X�nf]���[�6�F�+FF.�C}�ٷ��|])�/w68Z��6`�x�&��tw-O��JZ��fu�����Ŷn�/������;��8^�wӤ�׎iO�b��-��)ڽ-�HN]ְ�aL{���i%�)WVc?z�(	�Y[�G_̡�E��n)2S����طUAB")�9ʸ��w#*=*,��.��0�B���q����ƟΞ;�<��m��d��IQ��t��Wm�3��u,ƅ�Y�����uP-�:
�ݮS�ծ����K"��cz�Ni3��X��k&�H��U��F�D
W��v��ec�R��:X�y����Ƌ��"��y� [:�;y�.�昩�)�dr��Y4�[C�ay��΍��vͧk�P��I�5�N���<$���H���ǫ�:�u`NO+"�_`R:��+�%SSJ�=����Ӓ�ﷻ(,��Z�oq��m�_�nL�II�^���kTt�6��y<4gw?).���=*���7
'��U�ح���-�W�^�:��Ij�t�<[W���v�p�v]wܩ0���Nw��(�s������4sv���j�Pݱr\�+%����aD�R���~�3��+{N�yK:�w�w�W]a�S4^���k%�f���i��A�����V���Ĵ���ؠ\=�GM��a��v4<�.D,�U��x����e�s�ĜZub32�W�J�"�-�Vp�xIXCQ�ͩ�<PK6�k]��L�=��J��֧n;Z(:P���C��WF�N�3P��.�۱� ���S�]�;�Luf�"��F�������v�K_ܮ���t�����U�	�	گ�����&�}2���f����)W�f�7u�H��gy�����+�o��'E�
�a�Ki�x���x_.̜{I��b�HsWzmVc=/'��h}����ɓt����m#�'�V�w�fD#�5�b9u!\���Z]���#��@Y<LLW�ud5�m'�T7ÊԣGz����Qm��;��f+X����rS�����C��Xbv.ot8.�zk�ətZҤ�����g�~��)V��!�c��yr� p��/��ma��!�\�ӆ�S��n���*�ց�`���:����w1�ܝ�@��B4��z��lؒ<a�nP����n��Ŏ
� ��X��ȶ�x�F�5o2�w�{ �r��{|;�z�Җ���x�扵}��ūmu �T�4�Գ�/�˔D�U�Ky��%��O2a�('k����TN0XK)>1�@��V�L�V+�D{k��z�ݷs{�>����x(d�R�Z�ʋo�F�,YA��c%P��� 5k39�z*2�����.�v�l�L�,:we��h!�nB�8�+f��2�1�����'��zq�Ǒ�5�
�r�a�|����C\:���m=M��K�SU|��b:=y��{j�8N�Уn
��7:�ywy��bpw*����i��Z:��y�\%u���4ѝ&TH8�4) �*��m3b�5']*4�r���y.ZSn�Bô�#�X�J�h�w[A96όR���r��jL7[���֞1)��J�M�h��%h���ǇG)��x� yf�,ɔG|��K���}�z�S�9l�эl��x�<������ /���8P�,q�=�q��ñ�N�bMY0;!����j�x�u�H����J�+MCƔ�k&ۥ�9�x��ں��<B�G@�.�����u�����+I{M_%�hD�|"��l�}R��2�r�N@�uu���O3�+yF��j	2˨�GD;�R�:νW�mTf��+�ܷn؍�i�!Q� ���r踘�w	��jrYy���fA]��,Ήvr`m�A8����x���B�ר6s�a�)��s��%t�#jp��^WRb���evqV�::S{b>�xP6U�A���53�D��E�\j
ډo�oUv�������i���є�U��:�D̊�9�f�2�7.>�.����oq�0���嚳Z؜�j�f՘~��J�:���*�[+7�R|ޥڥ��D� ��F�8�0��R���
E�J�v�8�/1�n�1�΁�x$�i�qt(����[v'��F��D�+�Y�Ĝ/
ތ�_�әْ��)Z�{���8�-�þ�X�} J�����ڍ�%�A2`�zh���WX3c6�pS<��( @E�f36�����Qu\��s� 7�vt�Cd˨�7���+��wB� ܤ�Z��d�̬E�\�M=]E�1^������vz�;�`�2*�t0	����4��@�k-M�*MU�::�;i��s���=�|əU�>>�X*f�3����V��z�{���X�eT<d�#�h��CC�hƎ�軝0�w��ۢ%��2��Z����n�&��p�j�5��`r (Ž�C�����X�X�;�n�!\�� ���A�uw�(������;[�U	ҏA$Gh�9�y%δjڡ�k�J4�N2�����\q��B���J���$�wv���m2r����dVM�C���̮���Մn"����|�q�2"�*N[�u�<
��+{�N���t����[��H�+�|�w�GM���gg13�X+R,�i5�Oi�~��ǉ�k\d΄�m����jQp�Q���w�_�r�_y�5����~�-M�{WE34x���t��h��תZw����u2�4�=k�*����������w��O|��涽��rwW�A�2�$T�G�^�zӫؚj�|����=or��df�^��cj���U�Í������a�w���8�`e���-�)�e�w3@a�����O'����,Y}C���}���Ly+�<�S�R��*���Y��֚�Ra���޿@���h�odc�JzL%~�v�a��=����Q�Ʋ��h)b��ά���;g0�����B�^�8���l\	�o�}ݝK���:J�a5H��{��Z��C!�*��|��Z5��.�:�����G�l`�E��7rS���[;$�}RvA��>�ӛ���܅�b�Q�CN�Kj=����o�uXu��/�88��C��B�=ݥ����>2��x��m�2��:P�	i�&�Sm�J��nM͏��{Kk�A�B�76�+����|G��?gc��7r��+y����W}�=+6�n���l ���lBs��v<�}x1�ŏ��4���C�dy���8���1wEӒ@omf����k�k"���ً=�����˺JS�1�<�Y5�6�����W]�ť*f[�;�Ogo`���=�B<��Ǵ��~d����ʓk)���u.ښu��6�?v�����웨����{VvĔ��KI3�΄0�Ջr�]�Q�,�"�7�26�LϫĒƮr�������ssW(1\7+��\��x��\�wv�Es�QnwwwM��r����%DK�zj�"7��t��t��j�,QHn���.]m��l��d��w:��\��ccE�Σ�D/:�1nd�(ܮX�3�s�pd;���n���s��V6����.�Pc�@4�םG����W.ʍr��L�x�G��x���ӝ;����#r☋����.��wwu��fDm;��,h�4;��wv�r�H(r�Ph78R3[����O1 QQ3H�4���#�I#��WH<wQ븯���*����/;��/:�w��s�xub����At65�b�����ֶ�^�%����R�C�jUs��N�� �;���G��kv̆x{s'��t.��C~�Y-�'kj]G�)�)B�� Ff�/���S=Z��Y��U��� 'n�{�"0�����![����ito�`� BIY3Ţ���C�ܦr�iE�������� &#���e�c�A�o�o�q_���
F�P΋��w�]7.�����s/��f*3�pW4���h����얌T|rX�1�TsV���=��޽J�2x��߀[���.��%T��X���mY����KZ/5]�Z)�\���WT`vq�#���u(	<)+��{�@�낽U�
���oB�4V	댎s��C9�o==o �,�'���ͫ�G���@UR��T�<��\�;��*p�ͨ�÷|6��4; �����}v��JŜHh�U��:����>���C)s�����Y#w�]�ռԖJ1�g���;���GN���Q,p9�׮�\d�?W�a��J�k��iKS�r�%�zD��а�7)��ۘ�Q�W��`���:"�<@�%�T���(�a�E��w�}�[��n��)fb&�q���eR���v�uuh�M2]Z�.���<iL����ۧ�|�e��+�͐2���]�c��^���C�i���$���B��]"<�+����%�}q`��~@�7q��/�X;/����P9�/�O�rLuתfK��y<�x�ls#�i�N_��}pz������o��ۊz��Ee�n�^e�yK�C�&E� tZr�e��n�P������� ���1�{\�ͼ��N�n� �4��
K�zɒ8dKT��vT.YQ�F*u�T=�xHcm�T���=����#%j�����ni(�خgL�����%#��~c�uD�ʪ2n�T��)�*��ݼ�.���=����fT��
H�tYB.2��J�Ð9�����&��A%Lm-�u��!|�6��U��&�Л�\ā�?.:jP���$1�笕����ۮ)��xOu�p��nbӟ��St=*��}��K5��G]m�j�p�������\h���d�c	��,=�PФ9�MP&+����V+�p'��ތ
y�'$�k����SJ�Oq�쨹�1�0����A�� 23��.#�q�p�;I�P!	�h��]���.�ڕ;�,�ĺv�v�a�}_UKUa՞��1�B���7μ���~�q/.�F��;�Nئb}�(.Vg)V�1�8��Uk�>8Ʈ5�͞�	Y�%Cu��݉�{�?[c�6(���{���ν�#9��,�؟ ���Ҕͽ'r�gEsVy�����w.8�u3����0�ҋvC	��YÚ�oפէSԶ�*����y��u�z�ӎI�V�p�w�W������ 8o�k��y+e�tX*-���fYDfr�*��N�k�7O�ҩ5@8�����_!:�n&��)���#�%R<.g��K<�ٺ�g��d��֗oF��>�i<`�:L�4"��x��׵<l!�7s`���f=�ټS��R���u����=�fH<��VZ��M��9�h�9�Ƨ��-��g������V��7��	�&v��Q�k��=U�Qz@�SW�3��̡ıc��Xj}�^�z-*��i�)�2���hi-��'�]��LGeDO�� _��̪�W�����@s�,fC��h����9�g1Үqa�x����;%�p�*���@�]�?v��Hlal�����R�r��j�qt&�/��"9�
��Όw��;E�;���o>j�G���a���Y g��85N�\�V;��M��tm��+�.�
ϝ�a<�B���+ׂ�tڛ �{PҤ�bo��Gq�02�p���.c�_�U9� ��%>�UZ��\���� O���v�J�*�~�<�1;0��̹)�K�T��I׹=G.OnDr�E��踑	,8t*�)E�keA�O!���3#�����k:y�"37%�kZ�՚�Nmwa�Wqr��e��C��u���a��@�듷.v^!rp]PcZ��;������}QY4�k��xf]��j�+�ĝ�!�g��]��(dM���Z�+o;-t6��o�x�^���a��,F�
s�L`ޡ(lq�T&��_c����p*V��(ـpu��8`	��O���;A���n�+��|o�h�1�	�K2�f�B�5�cS��K[�t�:8F�	�A��x׽�P��ͅ���Q�����C�3-,��pO�Z}�F�3{`�u�!9�D��OӘ~N�l�9�=CE�V�\��m{�r>�����f�ڞ�K�-9�f��@c�Q�Ӟa:�M��Y�AR�]�7��]Ԕފ�]�2�M��5��o&�����@�{R�u� ZR��E9����Ȏ}r��mf�����;���g�B8��,u*.g�ɖ!i".;&\71�.� ��5��G���8��|�/- �ʏ�����U�e��RQ�g�px�\��rʈ�]�(d�,��2�i��
�SeZ1����r��
ڑ��+��qFxO�R�}������φW����nϣ�kBQ��IM9��m�^ �-^:�����a�3e�ˍ�Ҧ.
њo�C��@�Gu����q�W�F���\��z+�g<�<�M�f�����uNё��+���,�Z�c�X��r�L/��F�ӽ;� a����=,����p�!t>��4��ldڔV@�"�= v\UHeJ&�,�d�]�jQ�+0����D��Æ����]��<�E:%#p`����'��SX���R�T�N��8za��tBο��Sľ��;;�X���"j���Sq�'�Ji����w��x��v�Ǚ ���|����^�A��!��hB<�`�u.�yW�w8 =K
����ܬ�;�&&�VѸ�n�	�"w��/������c��d��ܖ���쫓�sٌ uCy`,�T l�1�pg�2�HZ}��c�'�R����>'���M	�=�6m��q�q� ��=��°A������W����𲰍�Ւ����i����w8�0���:n���ڛ7~�Թhŝ�Z���=I��y���E��y/n�_���nm�+�+��U>����z���o��Oi�5�	J'5�IJ*��?!*��s�,+.�^��]�w�<(]W������c�u�ĥ�qbI���C�U�v���wG�+ɘ����J6)K�:�f��۸0�&��׸x�5,�95U�zU=�<�ы)����w)\}.]�Yvu�;C���k�m�M�&CU=�?3�n;o�r"ȱ�,��}� �g+t�ʙa�Y�|`���c��t�C������/�^B�u���*��s�y�5�	�X���.����R�z4�rH9�A��u���/4/�t��e�V,�CG������3V\F�!��Pԯ`�/g/m�\�^�j�gi}�-ϥ��5�R����5�o��C !���)���O�ʺ�p�4����7�_�*�WYzXL�4�cC��Lh�ju����_N���9uw4�͑?oU罽E�=�8����a�u�C���!�Ǵ�r��*���+��][�^i�7 򨗮�=۳=��h$D��V 9�z��U��E�ɼ�>���9e<ǐ�f܌�zx�ua��գ�
�r��c�&h���CC[��l���-�k��V�9yn�O�E
9�0���H�q�`I{�^y�J���:[֛��=��@H�t	��]�
ȼĪ���s�	��u�m���SRD���tE��2�Q�¯����93�s*C�R۫�<�c���iE�������b��"��s������n�
�}�l�®��	W"�C㲡�B�7�!XLF���_{ ԕ?5��2�C���f�[E+ǑF��P#J���۷+��!�^Ǎx?*pt5=}a���a]�,Lu^�T0��Զ�G��\),�z��p4N���Z���N9\��kR�h��d�u?���kN����]� �^ǳ!����q��Y�큠�b�3�L<�*f�.���]u�|�����g�*���fj�
���>+ԫ�^�V9��&�`"b0��z��,)b�T	��s�� ��s�y�خޖ�>��R�d�x�E�~D"+���O��f�� ���c"�dT9�%b8jD�ʪY3��so��}�(�Fݙ��qS�2g8�X�ߵ}��X��6���B��dX�M.kC��(5��x�ndT&���������|��g�����j�{�wT|�"}L^��yu	�eEW=U TnK�V��D�]q7��dnu��X����s�xC7�.>�Ө�t�b�����s����c4�x���u���0��^��=OC����S�ն�����J�ʴ�Oi�;F/x�pڦ���r���1��K? m���d>YͲeo	�EMEWGQ"���1/c:�B�e��K����uގm5�<,�=�WbZd��1�E܁ןD��J��<ʥ��	V����\����Y�lU������C�2��芷J����'��xa��htd_iy��z�m��*dْ�oo��(̽�\�F����M��ϸ�J�����D;-yH�ٽ&�?���nSw��M�s��͊�Ӻ�8��)�눢��\��O�j��ܳ-����]6��/�4[���#[s
�1DT��K��XG� ����_T$j�E��d�w��ϭ�Ԃ�T~q����dh��8+��A�����BF���v�$O�K�n�9SD�|%��ܵo|���!N�i\M��-��s1�8Zrt���r+�J�	��^��p0�\C�׮%u��]��. ���\�k�aK�Nr�L�1)���BɧD	]͖���r]�V�>@�3�?�ń�}��u~^�xL���w����=���؅���"��&&���AD���4�����r"r���n���s�j0�vX���)�SB��l�q=[}���-9U�M�P�1� ��x�e�͏��zsratf���4AܘL�+g�'%lJiF�:yHW�7fJ!�F�N���<oމ�2���qc��*8��҃'O�~�Y"~�.,����L,�p��gY���<n5���	�n�GI�Q9H`���8nD���U�y�=қ�>y/PPZ�H:�ڥ[%۝~N�������LTs�7Mg8�S���̡��ҋ:P�+�\C5���klXy�t]f�`��s#�����a𙗹h�!���Ω��r�nC%'C`I_f�(��Q�y "�s@�N�3����'.�ˊ�*�L¬�jkŕ�kUwQ_v��-�V�^����Q;<%ZU�� /�4=����/�*8&�8=�C�.J�j�8�a��Z���0�Ę�_L�f�QB���F�2e�W�"2�]�r5��6�\'T-����uUnh�p�2H�Ne���5óX�F��Jn&��:��9%bT��c�����Iw��	0&=NM�c�]1�纐����B9UA�zn�iTD�|�,��]�lً��]��r�#��[�p�'M����7��B*�l^D�U��"@�Ȫ���"�Bp�e͑u�>�2���D,w��e�q���I�F2
�,p����rP��R=��j�[��%�Ѧ��a�XE_�ID���*�׆���'ʱ�	��R�I��嘃��.��Bv����&-���<̢c(�xl��2�A��i7�4"����.�RP
	�S��d���N3w"E|;(�Et�%$au<*}����3%|p�Y�S5Lv�4�VT���ryQ�Jˍ��#�� v��X-���~C�G?�y�.��2�ղ���/+)Fc��{�`���� }�;k-V�j�(-I��{�'Z	����j1Yl\@uA�{��7[�ոe�_����.�7��j�W�1�(�3Ώ��V��2�p�wg�=��M+��]N��M��e�,�.o-�q�r����Wt_lvJ�i���U�݌C�U��9igV*I
��@��I����Pꩈ�p̹+7�t�h�a�������ǀ4�j�Ou=C=K���_:��>�S��Ƣ����62f����Q.Z1ٙn(��<��o{
�ގ4-��ª��(��@Lw[�c����/����ͼ߻�q��r����dGs���������ڷZ��`�_ +�(	<);�S9��Ϣ���{w]O�����3O��fl?��5�r\�9�M�+���C /��O9 |P�{�N�SV�7�m��Nwϫ�T@�F[�^s~�KG���։~]���v,��b��N�n��ӕ��N��^k�aza����M5(h׆xo}��a�,h9)�L���h�<-�R��"��TgI���1t��悸�۔�G~�1¾
�cLw�H� E�|��ig|�S���j��\E�e�茙A޼y�@�l(gQ�9�/M*�X�1�4���Gm�t=�u���]�*�ː̐�f��ˣi����A����p� ��������R܃B����u������ܝi�ѽݾ�#O6/LX�C��]��U�W�!ӷ����=w;�cg5���v���(R�\v¡��N�Y,�7ZXM��B�I�szb��\4�x&pGcf�8r�����S]4�N�n@�om֦E�$�Z����*.�xH/!����֯����^ʕ��`T��-�J�./I�\3l0��Y�{r���y���}�hO�zav��\;�:z,�d#u��I�䵶��]N9&$z��=qt6y����v��v������ n�v՛(/4��G�HX}�b�E��޲�}�����58�#��ڊe9)j�ojK���l�CI�l��u�M�s��͗#i��r���n��K��n+��k����}t��b��w�M�Y�V�wpA�FE���Oi��wq�=z�m��3�THf�\���d"u\��X����_Y��.ZC�{3��: 7�%S�B��̫��C�o]B��D���E����	T�R���+��h�Rږ���d�.�<����H]��@-}g7.��E�㙗B ����Ex��DөQk���卖�9�;�7s�����(K����2qtZsXɫ���H��TՋ���s=�^/��B��ܔ���:5g��x�i|�Ѳ�ȵ�G�����M�z�:4?��}�Y{T��r�fB��t�1�ɋ.��"�.�P��j�f됨��|�7ά@�7M=,�g]]�E$��\7��
Ӟ��WaƟ�eJ�j �fެiVV<{�c��ܫl�'J����6&L�/ ���n�`�+n>��/�	%��D	}�| ��<�4�;~7�w��i��wc����їׄ�6�s��w ���K�$iŽ\]�÷��
��{��-�qr���$n��p�w�6��
��sx�=�����I��0��8L؉Km9�8�3�E�)'8���:k�)�]B�Q��.�����[�jiuK�j;\��[����Eq|~Ӯ+'!jv[λÓ���gڰ����<�^�W��C��;�Q��9�6kwy��z��ef(kF-Z�9�7���BWKȪsR)�)yǙ�S7׏hAXs��v(L���:�����ՂN��0�;]�۹�
��;���c��p�Ci��I1]���5��g�������A��֘!�m��Jzf*Ş��U�'$x��dIR�ݹ�mL[�{�]�W�X����WGC�n��2i}����w����ks��	��Mz��ٳ��袄ۻ�v��Ю�7g0D}#�._2LA�O��2�!xz���&Б��j�R��ʳ�7y�FQ;D?����=�����Ŏ���T�.��_8��<Wuj:��ea�kX��,B'fi�T�A�w-�j.��u;Z����^1[��n��f�9vu����l�!��RP)�a�M0�
��l^���l�w�j�
B��x��|�L�ߥ��F[371n`�X�(���P�;���	/��񹢉#�&�:��ڹr1�c`������(��r�2h�\��
+�"5wD���b#RHd�y�d!�h�)*dc;�F77dco;�7�u�wX ;�ĒPPQI���h��D;�6�����FQY�$�����\R
&d�Wa�&4��v�w9��oO-�@Np�%)�^K���I.�ݮQ����;ƮTwQ�6���]Ӻ�lX�����]���;�/�d<�n ��#r�ܵ͹s���I�'�ĵݻ�rA���DPWwZK\�A� �v��� +�9m�h��]KJA½�T*��\p��ˢ���A��X���ܹ��n|	��mݝnV�.ɮ�x���6�We�d�@��IN�)�.j��!;2UN����U����o_=[�������n����-�ί�G+��_�������=޺�o���+�^+��_�r���^��;_�|�?|��nU�r�|������c�Dd���d�c��)]S�"�J�x-���1o�s~��{�_������}��ק�Ѿ'����_[�W�������zzW�^=5s~o;���_[�x�+��7��_����h ��>#r�7�1��ګ�Y�#��{��{Zz�����ڍ�����+�?W������o���?�W76������kzW5�|�׭s��⹽�}�{W���|m�ݍ�o���ܿ��������}#G�9�r����Z�|�ň�G	��=��!p��5?zLE��{���^���j�_=|������W���}���nno����ս������7��[����z�|_��u�z����� }msfxZ��u���Z��E�Kn[�����m��jz�|��^��}W�����x��s�^���{�Z7ƽ�����[��zZ?/�}zԖ��o��6��Tr���矾�ڮ\�����m����1b"DR�J��^��c��]�`��\�����W�������{{�nU�^��ו�n���/wu|W+�n�^��׋|W>����z����WŎ'_X���@g���"#�� ��?TE�>���B/���N�7���d�޿t>*��Y��H��$}G����c���������+�x���޿�W�����~w�~��x�|~����m�����r��^��ž+�����^�UG�FG9���b|~��C�}$�/�1�K�^j����j���G�!���m���-����ｼocQ���b�y��[��^}���k��߫�z�y{Z7ſ^??{_��������-��[��W��}W��=+��گ��sr�����HU"4�5�{ܣ���H���"#���M�7չn~�>���/��{y_V�W����Ͼ�����m�~|��z^6�<{����nW?/~���n~/��h�1�>�>C�1�1��D���2ӧy������<�D�H��~���Q���������\����<�9��_�{oߟ|�Z
�k������+�h���>��׃�����y������/�o>��ߪ��ջ�����x��s~��ߧ����m]o�|�t%+�NWv�(�ƭ��m������)��}����kx�*�a�xjҘ���-K6k���9]MOs��G��/X̯l�ұ�]#�\�Pk_m	�Eq �WK]=z�y��ܸٝ���_Tt]�M*J��@ʨ3rɎg]��W�w�1�bf�追����j�_����?�����6��_������h�����/��s�_�{ҿ��x���/w��^�����_�~��_U��m����zW��^5{���D@0�}"�G�F�l*�V�ea�}_mʽ�����ڿZ�����[|W��kſ>uo������_��Ʒ�~��ŷ����W����߷��m|k��������}d5�;2��z�wWwzvדzo�x�~�n^-�W+��c�o��/K�zU�sno��כ��[Ź\��v���|[��~w�zZ?��]�������oz]�����\߭����y�^���!">�V׮
G��-r�<����8G�"C��z�\j1��>#}=_}~1B>�����o�M���ux���?���ţ⣗���/����+����zo���>u��ݽ��k�_?=_U�W���oʦo�3����I-S'({�M�nk������_V���5�����o��-��Ͽ��{[깿/?�}m���-x����<�s_�r��m˕��������y���x��\�w�U���G��6���̞���Nb�Y.����� �DE��Fa�B"�} D{�~�o�����m�����\�>-�����^��W/=|m���sr��}�^׊�o����/Mx�>|�^?7��x���4U�?S�}���3��=G�ۻ��{}j��?}��Dz	>�x������ڼW־�W�~|���/ţzW瞼�����ƯϾ�����o�r��>�W�}����ۏ�ULQ}>�G�xA_!_���DC�T��W
q�R�wG����|V
���Z+���i�B�B���B6�s~6�����~�o��|W?��������W7տ~����oϽzZ?k��^��o>u��7�~�]oo�Ͽ<��} P����i٪g�c���E-���z����r���ߛs�7�x��ǵzZ5��;z���^-={�⿚�7��������_V����ݯK|W+�j������"��������D��=R�}c�>�(G��L��;��Sʦ�ܕ���������r�{o}���h�|���_���k��x�z�zW�/�/�]������~����������ޕ�^��^��k�ƹG��������DS���|��@zx�u*����$�V~u;��{[�R�V{��(��CU'�^>��Ge�r�����{i��Ud��K��d��y���%��������
�t��K��(�v�c���]�"�Ѓ�q�R�cCX���ov�R;Aŏ����#��1>�>�;��o_=��W��_�}^?o?|��76�z���������^-�]��~����O֮Wֿ����zZ7��~���������� ��G�"S�U�4^]zv�,���M�� ��h����8h�?}\����M�ϫx�.�u;����}�oj��}_;��x�+�n[�.F��7���}���+��o׏�מh�#�"�������"�7�4�T[�yY�ݾ��=���b��FG�}����zoK������������|�ǥ~���W.�_~z���7�_����U��������^ץ~��_��|�wk�x+�n��E��[�������C��/L�=V��oG{�D�=��{�j-��ߝ�6�}�������o]��^��u�o��r������Z
���z}k�}^��k�?�z�J�+��Z��A_P1U���U!Z*���~o��{;�Nb�����VW���|DEb#��z�y���r�����v���[�z�����m��U�����C�ow�o���5�ߝ������Kr�������?r76�Ϟk�����}�x�⎟��hd���Ǚ|�܋��{�>�"!����V��1#�3㳢>"D|و��+�k�����ŧΫ���u=�⯋���צ�7���5��^6��7�����r�������[~������
$�\ίr����>�����.�ѯ����w���o��������Ƣ�"���8}DB�uX����P��]�o�����~^���jKҿϭ�h����W�W���~y׍_�ϼ"'���󮦧��.�"4G� ���/ּ_��W�~������x7�_/�"#��������1DFľ��{��/�}W��{<�J�[�����羫��ۗ/k�z�>3vo���Nd_{����C�EB(}~5�Ϗ=�r�+��~{��}o���o����ޕ�|W��;��W��[��_�y���^��(�=����_-����z^?�x���߾^���>*�;_�}-?��ux����mrg�P�|DD�r���_����#r������]���׃���[���ߟ<���������x`���"D}cξ">b�|�b$F����߫�����h���w��W�}X�$DCjp�(���Li>.7*�Κ�I�a��mP���~;j�P�{�u���^^�^.���L�wwޔ��ɂ�q=�F��<-r���-�8�w^�L����#�+jn̻�?Cq>�+�qe���|<�&�^<�-���A��Ȉ���
���6/I]��W��}��7��o��^6�n�{�uz[ҹW�:��|m�����9���6����[ž����������5�ߕ�ׇ�o��Ʈ_�z����o>u����߭�o���1 ��[�~q�����WT��R��G� |rۏ���� ���lx���k��������{�������ߞW��_U���s⿟D�>��Hg��G�#Ԫ�{�)�E-�M<�:�Y��8ݽ���H��ϕS�H��$���R����w�p�{�\"^c��\�Z9���;�c��p]}�W �u��A�U��%�/E��}��n)���0���2��0/L`n<�N͛�� ��UZ"��2��t�h�a�c�E_N�����ja'Y���мzs��[�_d�i���J��f}F���V�Qg�CuZ&ڣf��GY��71ȶ^�zig��f��5�UE�
X�9(��yg��n"�JɆ����jy�=���-��D�
�'An�?h��\>��|,+.�^tpp
�> =�d���h�<۝����+T��F����ɗj�^F��;�n�nY���� �cCt����j�]-���X�*]F�
��,n�Es���?A�r88'������������Ԛ��l7��}��p]����yKftBN��� ����O�>�O0�8�T�:�/c�t��
:���P�?h�������Y��O"KΝυ�^Á-
��Cl����k����{)��м��#� ߈�6�jqV�]Iv�����J�I+����fcݏ���e�4eBR��b�,E�\x`u�ƴ��s!�TKF����:����R���A��q�<~��{T�Pvu�L�v��
�+錸]PQ�rD�U7Z����"�'�V���6��[�b��A�/&Pw����-ԔWe鯕'm�H<3v��<��|��5�q�	�����u�C�䫀	��޺�O<-���|'��ymK�:�3W��ҺՂ N��!�/T��0BF�'�,���p��K��FT.��\p�����ݛ��*w�ʲr�m����:����@��O��Q��'Nn��}��+������l�Iƍ�;���{�s�7�~����g���؝�)�T�P�"y�e��<>�ū"�X}���u��u��^�����c��"���=�\ā�����ݠlV�A���]��y$*0��8���2�����W���u\ԡ��*s|����{�������ftZ���׾õ���V챲t!���(:����B�)b�T	���Q�sd|��[�~~
�k�Y�,�����r��V�˫O��~��esUw��e*䊢�����c�B�����R�	ͽ�]�a�)2�<���EiR=�B_Oj7��gc���T�Y6_*�'Y7%	ԮRz�T+\}̕�����b&���}L# ���Oa��-Ȟ�����0��ú�A���@���Ѳ�}��W�u��waޜ��K\�{�*B��Y<�#�J^ہ��{\���iX�~C�c|���d�Օ����]�(6 qf��P��@\>�:aә�����N��Vr'%����^K/v�]��e���'�z
��.Wњ�
��1�����θ��45و+X�^<���I�ҡ�-��Oc�"��3��:�.5HF+O�;`�:L���Lo������ �]�gM� �=!��s��Q�R��M�
��J��I�X�E	�ݦ����u��/i����9���N-�ü2v�����Va��SY�<���Vz|m�'��W(��M����A��U䱷���g��S'E܁ב?(�J����eVm}�̌�0krk�ס=ɼ�qjጃ�Lv�΀�)�\!�rO)��@#'�%#���q}y���b�W����3V{�ȹ�=�rDr7D௞Z�	�D�c$�������~�(�<~��2(M����@k��v��z��k�e0V�19v��zta���[w��xy`Ŭ�m!Ws�����o1a#��o+����SZ�F8���/�Sm7:��{�:��z����!�n�"/��G���:�������ܵōH�g�s��sF�O��Lդ�&��l�:���;�dC�"a<�v@�ɥy��D�Zsm�����,80cr���f��,��1
�}θ72�� p�3p�b;&.��2#���	dLU�I¡-ț���Y1K�$f)cv6P΃!	�'V�Ή���V
6si��W#lWK�f���<�����I�i�u���X��(C���0a��0�=���)��V(M���&�ئ�k8c�I���z�T1_�Met�=���T뒬�"������_;��cAw0�����!�)�ȯ��'U�G*x�ba&�YϤ��6$.���o�����.�!��9�ö����w��d�N��Ɯ��w3aT�X���/c���;Sy}�AҠ�����ʴ�d>
��C<�i�1�\D��<s���Zڸ���t3�U���9��vH�>^@U�\"�'g����+��d���h@iS�6n�(<��B�c�C���z���2➇8Q�vq��Mw��g���_V��v*[
���ܚG��������%�uv�V��ۜ�WD�]���ٸ
���ɶF���W�(3�'-�)��&d����k�֦UvGZ�P�u�!3[i_^�X�NZ
s�զ�͕룯��\}1I	�����o.��r�kU(��&)��җ��WԜ���`Na�a��Z-o23�u��>���o9��R0w)I�F�y�BF����z�G�^om4�7B��,��e���<�t�cJΜ%�.dV:�2B���7)����gA9�����o�*�wJ��|z!s뇐�,`�7�r�WKǖ3�٤n���M��җ�On�tRC�&-�����U��\b��g���#�,P�&#�T;��/>����]a�+P7F�<%2d���:�0���1�{_N}����5*��L��Fpt�{se���A!?�ш�\�퀄�D7�"Y��a=��P<<��ɤ��5���{@q�p�F�m�}��y�뒐�&!2V�aQlLLR��qa���y��D�;7��qzv��Qn������^��X_z�	��!A�����]�!
��"����J9��Y%����q�,N�L:���Ñ� ��"�Oݲ�.zw"n��D���b�@)U��t{{\*���qg��a(�<<�zO����T&���N�C�v�3U��n��ܶ�f�W3������͛�M#b�*�0B�N��/� ؞`7��SjnS�n�J[�	��s�<�f���yn�м��$��'\�l�ܪ���%(��[2;����m��O���f�:��nU�S�8�k�t_j��$���Vc�A=kf��"#�O6�ir�+���-��Ţ�S0p�|�
q�h
�7��1�f"~ki�ʙ�8����d�:��H	왻�fϾ�A^V%������!�YzxX�8j0�J p�E�;=[�ˮ�����hkT�SW���]����v����/�p����`���/��N���X�P�hU������c���J���*zh��b������ﷷI����ȩPc#t��Ӱ7c)s��co�X�ҙC}�ƴʫ�x�%�91FŲ��c��{���k��9��ZC��:3�U�ce��z�K(>1����c+�N�Yu��)�1Q/���1Ϋ�vpz�u�]���T\�(Fү�0�6#�i����0�"��nl\o������ˣ�ռA,v�UC���@
�.��Њ�:"����837�8c�y=N¼SdG[U m|��C��E�4O@캩r�����ʅ؉��tJ7�ۍ�em	�}������01(�P�9�Y��#���# ��nh��1�wL2���W�2�ݸ/ΰp<7U�}��d��b'��)�uj˖�Ci���a��_G�y���{�$L.'	��=q<��Xj��˩[���6o1���i�P��p�('>��d6�ж����'��KÓ���`����
"+;(%�>����c��'��$k�O�'SK"rf5�V���w"���R)9��RB(��5S{ Ѥ�Uv�1/�������s��'_S}L[��\�u�\B{qQ2�@ꥊ�
Y�G\��/j��>�4�G���B���yw�]�_�5�]}�َ�~zT��g0����ʯ5�&yP�z���Qj�\Q׮U����1��N��(hR�$�e��Q��z��yn]ש��C��X��꼈���;t�ј�u�j��������nT�2/Sfulws<yHV08�ڢ��0�ͯ*B���/������iȱ�Y���
Ѯ�x=�
�-��K9�9.6�?Y�c�L0:T4��I�+�rX��컈Y֢�a�0O���)mE����F�g�y��}e�gS���'���-�{S�r�}&Շ�kC�|W{��"�vrZYʥg )fL1���7�̽9���)��˙zhT
��Ox�nf3��ѹ��vf\�T\�#y2���:bD��[?[j�:� P�6��Ϭ�sYFɌ�h:}h���ܝ�-���F[�-����w'�z��\���Lڽ�K�e�S�u�7Ss
UȲz����+1Q��X���^pN`��Y�	P�Ϸ�P��E;�KY��q#�'�sc|rݒ�z����4���כ֕����Fk6��4;��R�2+j��:]�N|̦��W�@��X��رt���#��wU_j�G.l��(�Kv�ˏ�HZ��`�1�����s5R����zn���0]��*��ՌV΢K�+�3�k\wK���k ���e�g�]u�S�;�K����[92�!u�w�
R����>wo)�Xz�o�!ͨ��Vқ�9���O$���4У���V����V���(�<���k-�̼4�[Z?�k7�Q���#�B��� )�A�˓g8݇���:X���j�[��ݣX��X���[��q�ک;�)h"���:�������.�QBޣ�ɶ���b�9�ae�#b���,�\�T�>xB�r�r�qn@ ��e�й�s�PhJ��Mr��kio�a�Q7rS{���Ͷ�?��#8H,�:�o;LaD����7!�l��B�I���<��%����k1] ��%hS8Rx�l�#]DMv%X�/h9���9Vh����M+�c2������"��g �Lݼ��y��6�*rn*,c6S�V������ô{�z�(Dp��y��s�I�_�Êk}�r�;�h,$]+r� 
t&t��
#�cx"��6�+�蠫�@v������	fvm�,ԣO��s8�J7�o��f2'�Veh�����-���Qv�\Ŗ�HS�f��V6U���F]ކ]F����GB\jC�����J���6Ѱx�m]��R�v�G�J�}�۽V���0��e���	 s�l���({D�mfIΙ���Պފf�8�g��X�{�>��4��!�����{ٹ�9E��=�P��]J�on�i5�n0�]i%���i�W��Wk���⮺땺=X�L>5�*8eu�dΕ��X��Xj�%@�쬙6���91���tvb1raD���8	�@��;%�D�G�*ZW�AJ��=��=�H֙���8�7$����P[y�;1�˺uh��H 9�d����#�fi$&������}j^�r\K�4P�==��D��Ȯ��u��^`�aٚ�k�V҃�ڻa�uq6x��;E��uo�f���6R�8�Rۂ�a сy3Н8��Ҧ�>������\�"�[�\����/��@3wL����u�
�P�8��u)<���Lr����F�j�s	lXV�ң:U��D*�f����^XtaP�]*�K+c1�8)�"�_����2>t���H�8t�t��j=�+&Z4�m�[���񿮮�d��rV�(YV�En^0��w�r�.�e3mτ|A��U@U2 ō��p޻��λw:��wCP5�E�ۥ7wc��q�����7#�t�m�Şww;�4�I�E0 ���#;��i1��݋�ݍh(��\��ı��0��$�.r�aD��s�77�v�3������a�dgu����j��0l3b�	0
:��]+��F��f+���r]ۥ�m�n�Ix���!�k��#�&���r�P4"X�K��#	F��&�;��&��ٓ����wt�d.�3��0"����1���s	14���9ۻ�w`��B@��wk��1˴��w\×Qawp�y�+�BaK�q9���\���O
D&��l^w4A���IP$�@>
�> t�>e;�tz=3���f{�xFu�M�h�>��֘e�=�� ��k�k�d0%�/bp��^:��V�r�9�������購L�	i�|��W+�{":��G�+��ju����0����̡uM�f���Ѻ�I��U�C���Ų���]����Y�E&�#���?R�`:�[��f���S��tU����M >��s6�`N�����C�	����QP %;�'�~wj��6�.�c�'*�[j����܍�h���|�;H������X̧�����X.p����ip�����q1@ �[���@8*�o����{�����|�ƈ��8WCܹ'3/�a
�w�s���ٔa�T0��Y�1c ���8>�D>s���nY1����jƮi��
��9���SѝD@��Ծ�|M.�He���j/�W�!u�����àk��W����H<��\�r��y}S}<��t����n�%[��~V���yc�	�)J��]����ึP�)�����m :�*��o���1���Ӂ���^O���/PV"����f�ۺ��UlB�a:�W�qʖo��a���T`J��l�H`��~�C�t��NdZY�0up��p���Y��`�#����Xݿf�qhl����mٽ�
����q�=�)cٰð���4\��gz����ΉU��{��U5�n��U�N轒�BH�5�5;���\GK������+K�}�U}�o�>{|VR��U�x��C�5G���^���x���MgOғˬ-��-��bV8ַ��Mp�<-ҷQ�l<7���4�&�DLwK�:�u��L��9����1���|�g��u�݂���wI�ʗ!VjO*� Nʬh{%��@yf�kcҜ�;K���V+��uh�om�Txӡ4�b��[��c:!7��v�v��V�̻ʬJz�XO�m#���!�Oα����]�/F�"�r0quE}G�u�:{}ժ��Q��t�� s?LF�vn!9�c��tƎ��㡽���	@�ӻ}��*�9����r~�Ы�1M���#��]�y鋁��6��Ӧ7�=�(�����|v���ܓ@��&H��e�UH��]1�a�<4s:'u'���ʐ���,o<2ڕ�:vav>�u���6�ǩ�b���.����>
�ez�YO!g��W�t���D�+�����=h�iR�}$uA�1ʓ�<�ER���g����<�����R�J�x�m�V�h�Ƹ�v�˜�q���G��ٴv�j����i����̇)m����'#Ғ*��Փ]��{fs�C\On�_e௣N;OV�1v�{�z޹�^�3�-gs�
�lEu�C9ǀ'iK�ػ�;��'@q��z��φ`�w� �H���:�u�eQ�F��q�Bc�T<Y*Ɉ�گ>���.���O���2����$����X�L`�I�bᾫg"���X]w� ��F(O��-����T<����~��9���lgX���ԅu��� ��y�����o��� :�\�OW�u�u�4gt�f�n��}�~Zs���CL�F�yT��)�I����:����፴���r�V3$<? �ԩ\b���r���_3�:�^?��
�g����}��cןy���|�r��u��L/{�����V��F��{��V|+αpg(+b\֨�׽�����U�n��2#�Ż���flg���k�Yȗ�*f
�<�Z�o�{v��.c�5��p)�F����@P�L���o��e��y��k�h��b��K�6��/V�Ou�ǩ�g�!i��1����!����e�M��p"��H���,�v��X<�	��	dEz��:hu���7)�,Ōy1�����K"%�(�ݙ��[�4H(a�3L�2��[�NE\8j���ݳWM����4&�J�z�?�y�@ws�ܖE�ĉin�e��!��J;��l�s������hd�v%�Q�r��D� ���j�u�q�N�J��V�X��Nѿ�}Gћ-��Qu�HPl�۬��R:*�%�&�HuQ{O
��צ5+3b�jK=�3����=���d��XPEƼ�����j)Y���;n*��T� P�һe��n�}Y���+Qc]�>��¡5 ��0�9�2S�����b
�,���)�<�>+G����YP'�^���n�����A˔��xx?Z�,:� ���u� �Sq:x���|�$]�{a��h
�4�w��l���.뉿�T6Y��{�;�O2�R2��K(@��RI굛[���c���(}<{M�����'_Tkj�.q��j��w6�y>�%���R^�۞׸k���8߫��sȄ+!�M^�ˠx`�BT�ŧ?>;����\�gM޵�3�f�����E�ѓ�uϭՎqxb,T�g��S'�~�W�7�w%��ԧhP�ݮ��n~ɥ�A�Xuqȗھ��t�U�/9`(2߽��|�im�U�#�����uEnc���t�=����#�E�4��c��~?p+ٯ�7n�J�*j)�5�*~�͓Z,����F1�j1��v��h���;{m�r��m�P��\�{�ԥ���'�N��c��ڞiSG4���P����C/	����K�n�R����P�6��2'Y,:%�i��:#��t���̟�����_n��|Ϗ�E\h�w����0@�bc��0-�A��Ԅ�
!�&�7�5�z���YX�o�=]
���{�^+=�P�>Q�@ʌް*,�l�D'_p�כq!ٍxn��WSw�ܶt������	H�GQ;>��yT�9J�ޏNu�7˼{Y�D����]6�P���H���}{ii�PVa�(�9)��Ã��񖗠�����=��]l�%-������N1c��x�O��j�{":��V�B�N��5�4�pu��yY~t�̲��yIj���G��Ӂ����q��zk�J�!�A8T���ѣPLF�}?u�X��G���z���[�����j'1���n>��I�C{*QX� FIhiF�9���O����mX?X�6��V�mBF�,��a']�2Dj*�Z.2�E&�$-.�Z&a��nΘ��,��A���e��(�K|	Oy��&0`a'1�8Zrt�Bl���d_t9gQ
d�JLT6&����}<N}Ja�Nو��;��xꕹ�U�L��m*O1�m�4����Ƴw�ǽU�l�W�YBe'�Pڙj]���w���ZR��Y�����-�����.9�/��&�-�'e�;�2��d+�d�O5�����r�R����'�˥a��H�3�'�M{��7��fW-�]�=}�G��7��L�ʹ8t�vMV�z�'U֟�P=�7侴׉��!_b�7pL_\F�M�e��喐�X(P��z��D70E �:�'�v��2�0r�u-w��,�b⏨h�\F�J{#��lEK��c7b���Rj�}�j����su(Ś�;r�z~n�&y8���<KW���_R�wo`�b��̘l�f�� ��Pl�0�T�=��0�wA]ԟmuf�U�G`��Ęc*/+\d�l�ia���N�3���u0���Wb�zٓ�Av����	���*')���*6&�}�k�‛Wq�/�;�3	XKz�����w���8�ux͚{Ȍ�)~@U�U�(�����W���4=��}ٜ֚nU���&h� ?�.��l��yZ5s���]��b5c�*�5�%~+���&����cO	���F_k��~����g�*��?<y�S/;˂<߫�W��5G΃��u&ov�Y4�;�}s<9S?tE��3��K�f��օl���|q�ۮS�x���avn.]�����E{2O{+6�
�t8g��n�:k��9]��	)����+��j��ũ�(i�ul)��Vu�����=�y�pT�Y%�A�+��仞M�ʷ���PY��7'v��*y�\{�lyyS��Μ���}DD5���%3�@ڟDQ�&�DM�+HL�>}p����}0��2�O�]�@5%3�wXn�1�Y�a��p�舠8�וRD�B���
PS:%�IP�T���{6Ѱs�E�in��Єղ�8w.�\W�H�3 gQҦ�(r���ު��Y�"�����G}�h�ߺg�\F"T�ta`��4%�J�T��.�
0b\|I6)�Fu�ݫ�z��b��멈bƃ�	ހ�绑 TF"xv'�w�7�/+)/�J���q�[Z���ɍ��چ#�,l7�l�9�b�*� &*@Ů�@�2oJ����9=���jW|�z��|f<K���1bcz@���GSTE�H�B6 �=�î�|��n��I���1,A��Ky�^Z�'�����<i'�E��cT�k�q����͂�p�-��%� �gd�1G%���W�s����΃5���pƚ�;کU7��ؖ�ruW�/,Sݎ+}�a����ğ�eD�B^�#��b� �܆�Bn�o�+��?c��DLklω*��"�n2}+V�׻���_�[�ٶ~"	]�R��Ž�끚��9y�y�_kRi��p��24�O��1�M]�� ΊƊU���і4��ǻ�'�Q��b����_I���z��Lp�j�7��UD}}���p[��ƅa�[�B e=��P��s�]�>�#���e�>jT���[�V1��z{�����]ڛ��z��,��Z!�<�/�����mV{]�0KM	��aWc��z��Uq���1����1���%�7::���l���T��.ivsN��vo�7�&$ ������TΕ�N��>Sj�
��7)�ƙ��X�9S"�.m�e��9L �<z����-.5�C��xT��z}���qe3��FV7��q�
�b�Vқ#J��e��}q�0�m�� vL�:�� ����ӵzS��TK����j:��E�������-�2���a����@�-�<�|N�V�X��Z�μ(���Rj��<��!K��<88{$`��i	ӛ��d�r���5eR�Y��������g/��bi�h���ν�<��z����4�5��M���;�s�?>��{�4te�:�`/���VI����T1m+��|���
cc� �P�rj��ʵ�@¦����$L!I�ol|挧pÝ6=��}:�#`v��xX�<�zӬ��-%]j]5G�Q	I�jöi�U��x4��꽤u��
���1�>�q2��z\k��vm@�,fQ�ۥj���~��#舎�m�ۂuP[ ^L=~�9qt�U�"B���vy�W�]	�+�v��W�+ϛi�Ef;�~�f����O����0o��<M�j�d�G]r�X�Qxb.�< ��oD�jT'��L�$�c$9�MPf/�3��T�+�	�%���D�}�r�'����s��oݭ+��~�z�l1q�8ȿ��r{\Ć����n������+����fl^7��.��]�oH�>�٪�:��8�> (_�����k�h;s"�NH�Q�$�Ĕ�`57hy�XvT�W����H�g��?-f��ٽ1�}�@��0�/��u��vE:�b+;�=�3�=<�X��A
�꩝��i�j���vz}ig�J��b����K��gxF(����V#X�+a"��6��յ<n��4hȧ���1��J�ʴ����R]����2�D�Q��+��j�_�wq���h����o�����p�t�o�Mg�	ja
*wu1ӳV���֔gB�փ2�{���}NX땗�Y #��Sq&#��~P;nډ��=�7��t�GwZK_=o�-.ݩM�lu��錔��ȋ�ۋ�jV�͠���j���	�������]آ�mob̋�p�ű�����;�
� ��ސ������pwJap�ޤ,G�;:r��!������_U'�}"��>�޻�����U�
9�C�s9��r9������z���}��g�Җ��5�˞�&@f��?A�t��=��:�.���$s��Dr6�N���*�}
��_+��z���$&o�����$L��,B��K�B�Uq;O��1�q'6N�|��w^��Χ���q��"�-�vX؃!+U��R�c�=�. �.���;xN|vh�ohrڌG�|!ë��oH�{�?2�aw�K�g�ԧ��U|�30�����=��7�Z�C^N��Tkj�{*��mP�\|6X5Y���[\���{�csn���J�ܭ��K��y��Z�)�D��� ��g� Lsu�*�z��w�գ��6|��}�݊V��=I��~O{���,��ߜH���E�����*�,��^����|�f~����9H=$B�yX����zP񙯴���wMk cN�����^|#'��M8��R~}�S��	��V�]�
��+���򕧀S�����C�8��~S�䶒}ͼݫ���ͼ��6�E��1B��v�,��I�XK�m�X\�G�p���_{���;,�[��ޛ��(��n�d���X�Uqb�"��ч7�>=r�v�Ft��+�f���6̙�ۍS`��� �GB�Ft�N�O)iL{_#H�.�0�ōc;�v-��x�����sZ�U��2���ii�t��XNe6\Q�����*u3�حV��'�ܼ�n��'��U[�.V�B�c�̹;��P[/�����e�^�W�ȧ�q�)��ϽVFD��P�Gk(C�1,�6�d}�c.��YA���;z+��:���keZ��QӮ� ��&�e�̌�7p-O;U�!:6:�s�l���e%խq�ڣ)[����\V��[O�[7n��^v��ǑX���Ƞ���o��ŷ�P�AX���^��B%��2k�g�A�y�n\s&J��õ���{�*}���G����#�Xeb/�E%�A�����V<v��I$��T���T���*�LV�ͮ��[��htc-6�K��yu�W�ݚ�a�qWT<j�y�]�B�\$��cw;���t�rH_:�h�O�i�nv��X�f^�������.@��7wY�+�M�I�F�e#M2����k4��)�s�2),0`�K�t��̬9��ue�en���"H��*R��f��`n(��\���$�ö��Ǖ�ƻ�9�����	�̼���j�1��X頻�\:fj�U��IN|)��ɨ&�gjG5�FMV6�j�zNw�R���<��CQ���Ƭ��lz��n�%`zPś� �����,׶W-�oNԀ�bZ*]��;;Pу�Uc=�Et'c��#��fƀ!����s�V�y\���eM{�+!:O,�*&u�3d��Qu������tL���X�Dr����kU(D���Z૓�%�#y&��޲�=����v�.��~s���[��>�9�X�Ykd�f�ޗDϔ#4����[XS�'rNF�ꖴ)��̘l��@'����%KՀ��,�F�R��剬�%�����:=�eTO��T̘q�R\��s!(w3�7&�\�.j��Ks���X����n�U�`�&�U�
�hh�u�x�im��pP@����\3��5���N�F���!3��놉.�̘o��l���.S�ц��||8�C�#�l4/�{����ii�.˦S����6fV�ޢTtޠ�i�����=O��'*�V�̦��~�u���=1�&����W`~Ju��2��](j��*
�i1�#��y�#ܹH��N���EX�y���or�e'dz��M:��K|�A�ܠ&�ҭ�*^�5a�n�#ED2���;���	��s�\P�{�׵)2����R$�nWsq2�\H�DDQwm���uܺq�ӕt�˼볻�8\�$�O;y�����P�Zs]�;�����"Y�H hdd0�K�ҧw�pH���I3I$QH�ـ&K�����4le�pGws�j9p��#AF&Yw]<n4`Q$L�&	H<v�R$�]����I�%(fE7A(�k�Բ	�L�<s��$҄)�����dnv7;�fS��Lb�wvM��	�9��w�d�I�!�r�Y,�bHf�C;�Q�ĝۈK�"��\���L&�R$Jd�H)@�7u���wu��)�%9��RF�^w������lݔk�^�.9�2!ܱ@N�,���yw=&n�[M�B��o���I���WG�=�V|ǹݜʛW��������K96�*yҁ��<�\OA��i��/ *�R�}��}~Të�$Ԭ��o���v8J���ќ�]� ]�o��|��vs�b�f�ܘ�X���|]g�R=h�o�;�&Wܾr-����J@�[2"�Zg"5��7"�������ߐ�nS���p�!�_���<��1A��Hh�\��r���R���L�eKT����̈ٻS�N-|�&�p�"���ٸ���������+"HL�>}p�'ON@�v��ȶ��\�����z's����d<?Wk"�@mϛCΗ>E��jU�:']'�ˉڡ���ȫ��׃/Vc+U+K�1���!�T�(�G�m$�9��*����ܵF�XSy)I��3��ɌE�����}'��1	�&X/����ER�N�eNe�˗��۞i7�i�aKp����X�nph+���r���"b�r̻��֨3���n�)G�ى,LZ��.	��a�ϻ��/�����;LA�1��O,��U�[�d��]���J�j���r��G���:��L2L㕕���'��kȖ���S��u��>�Zq��!��&�R:�YU)5�8e,�ǧ��ݧ,����\�nغ�l�H�<U�ʣ�SLw\cB������:��,��g#W��p-7mwVm��q�����>�>��舾[��9@s�h���TGT_Vɨ��� E�ޠ!_'f��5 6X� B�P�_tO���u��o0&�'qz�Ep�1�[��T^¬��r�j0�!Ȁ�YQw���}��wUhY�I5~��K���/b]��ǅeg���k����:�$�͞<�+Q��e��L��榆�'�\j�-�G�%�u��>��U
ʞL�zɦ�2g#r{������%����m��6�_�T'��_=5�r\�;q�~6V�Ue�Y�ܹ�?r�s|E ��`��T@�O%�u���A�p��n�"��ԃ԰άݥN��E��G�em�Vc8���C��%�7
�\'(h������}�Ͷ��sC�7jCM�ۉp~�j���_E�˹L�kyM�����_7�<���y�$�y�Nt:�Vu
�+};��'�������T���y��Kh�P�����ɽF�oì�����|:;
��J'�|�-��hOƗ{>���j�B�\߸�Q���[W�TJm^�+;�eї���9�A6�͊`�����k������L�����գ
���G��g]࢜ؾl�Z���U�Qckj[k�oڔ�{ ��L+r�=�ѓ��+��w�sT_c�#�k�U}�}�ɯ{�.�戟}����ɷ���ތ����(�W�%����	��t�$��;P���ˌ}0��Q}ܘ�WFL;�4��WGF�(���;��.m-�������޸}u���Ի�:�G9�꧖w1="zi�R�Ȧ�KR;&!Ϭ����Z�]�W=ϛ=/���mp���l�nV�ԜkH�h
��
��+��[_X��Wy��UNm�(��v��)�Z��Q�����u��l;��� ^�k��U��F,sDs(�'X���W��c�3���mT&���p�1�8t[����HaUS��4�w�����'uĻ�N��'Ɵe��σ����~���z�Y]l��r�P���L�'Ϩj��U;��2�>,�xr�z,I�{"	�ǭ�R˺�S�q�8��OQ��<gVl��]�%}J�
���t��
g��j�����P�m�PΚ��0���Zq8����q�gsY��;v��,�
E��s
�c4,EY�&uKWdl���J�P�uX�Nbgp1��(�Z]N�ZfGb5v� �ݵ�����������34��T}��i�;��_l���UD/m.���u�땕�8�����*ĎX�갖�����ecõ��	
��>��UgE�ˈ���\�Iי+5�"q?�9n4�E7�U�\'����%Wƻ��Գ�+�F���G��/9k�������#�.n�;���k�[]��);�a�˨�Ҏ�s�������Y����˟5�OC�臫j �n�v�Zؽg��[|�z�B�Bʉ*K\*2}7�nFX����a�x]k�v�љ�k��K-�vVԸ3�]����ǎ�}v;�}K���f�D�f�=�j9�^���0�T���
��V����ˀ��L����:ɣ�W<�s�L����8¶�K7s���r��Y4���i#Y�r��4\�W�=۴�����C}M�yNGT'�?+�<.��J켝I ���t���U�{y�ku�x7�n����O4R�v7��R����B�ՙ���#�v��K�_�zJ��[��i|��w{!��pJ7�*��K���{u�����{��)��[�yR��t�Lo��DS4%�����&阮|I��ﾯ���m�}A�K,W�p�f�כ�}���MCYg&�p�*�T_n6:�e�g:�ޔY���'�TK����ʧ	��-��������r���IQJ�q�G{,��o���{y9���j����Nz�w��k�1o�=(�N�Z�y��'�O譭��.:|�~��.��O��EI=�ϳ��}��p�1cᐖ��㱍<CN���k8������ހvf�<��rO�h)ym�U�;o�zz�Y�m�����ᘂ�j�[����+0-w�ΣM���#ke�o�b�x{{�cj�b� K9��[�Q49��i꯬���<������>o�
�͵U��sf.�V;M��Z6�o	��ןJ�;�O����ϝ�9�����ɍ����OB�s��n��x^�Ъ::�K	p�h�.��b�@������Pu�K��r�K:bQhk��S;H�DVb��������|Gm�x�T��V:�߳� T��v��|�٤�7�x�p�9RB�������O���#�&ѿ����[id\r]�"��\d�|gl��ZA�U�:���]$ ����W��}���R�\]	��Gv��φ�9n�w9V0%P:TI�z��u����vbT.��Ś�z��I��F�}ԞhWF��1��*��F���|ᛌ����ѫ�IV!��#2���)wM)�����{
�a��\����k�iKC!������ͷ+���VNve��,+��Bks}���j*����,ߵ|B߸�x��ɠ������a�vŏo�zB�I�MC���ڎ�p���{��B��V��Y]�##z;�*�]�1�.V1w��o�#{�9�s0b�e�Sќ�׽��<�\�E:FȜp�o��:���[�נ�gNMC}9�UnuR�?�k�7!E|��O(�sÕ����[�3�Q���zg��ϩ/1�>�[7մ���6Wm|���><�������74��gvサ���z�KT	�;�dݬq�\^Eꉊ�x����j1��Q��el�4���eu�C6qXW<!�;P�he,T^��e��8G�˭P�RW.KMm��A�W�®�o����)��G�ҰC�2�T���rT]0ƺ�YN��s�xh[v�zJ��Qn�]�9R���b��kfܘ�`�&�����C�d[[��}��W�!�1���1;�o�w0+����Vq�(�]������}I����z	u�ܕ|���$�,�q���6�T�Z��~��\F�U���X�ʙЦ,� j�.{(�[�E����=�t G���!���b�жt�mk���;��Z�Wjo%M����:�����T��C̷\�M݆�-J�?��a[�pJއ�oF'-��	Wád�.��u��s�y�]6�ps0T^���a_t���e'��r��(�t���h���e������j�b���s���uէջ/�:���h��"��rv���7�ԝD#/Q�����W���ח�e�YQϝ|�i�ˆ2�+�Ww6]\��.9�¿�<ʄY�+c�����ͥ�l������6���Gݫ)�:�PO3i���7�q1��𱞌��h���u{^�����q�T�yM���{�Cs��j��DYG���R�郰�jzF���`��9xQf�����h+�[�-wiԛ�ܒ%����<�ԵV30C�����m����R��DD}�MN�Ors����я)�a�>���;G���V׿|�"�I��(7٪Y��3owq�k�f#����⾇��ByM5�k���8�pjlo��7�B����jiX���0��l��Sn\�F����"'zC��9Y��͎�7�u~Z=Qo�q!GGؗQ��0��މ�TU���W��fp�n�4����A�=EAڎ.6��R�~$[b�)u~{�ni)�<�om�g5���W��\��^��w���!v��6����O,��q�:���i��o� �쫈LwV!(N��Qt�䝖��T·F�n�Q�V�ES�q}Qg^r]�{.��ϩ�������[i�D��FM���n��5���spb%lLE.J��]�5H�I��w���јy��GCU�j����488v��U������>�>t�э\ۧ`u\�'�q��r�W$mVV���ҩ�<B	�K�yݹ��o:�*37*���]�r!��7(�hܛ�m��|�����z��Ԧ#ÕY�9�g�r�4+��e�z¹:��b������c���K�Yo��J/*aٲ.Φ�3F���ĭ^���ﾈ����iM��R�Uָv�p��@�YS�09�����ǫ�٠�S���K��Zs3|��X��[���[��ݙ��zU�j��W��.���.O��7&1���aP\�8���z��r{
�a�V�O�!vY��ž��Y�W1�W$�!55���+�a�M\�cP�5a�*�:k+�@
��9�睞��f����}U0r}e_�����>��T&����w�}
���9x[�+8
cUO�Y�q�T^b��s���{\G�@����J~,�_�f2�5n��ye�y��w�W���r�x��;����5�)��ۉ�Z���Ӄ�\�oy��m_����m��cw'�%C.c�*���An���"]N�����{�a���{��"�"���8�)F�U��*����-k����^��^�y͞Q��'#|�m�[C8?c^Pҭ����Ӭָ��PfwK��1J�	���rW[}J23�0���]�Fќ
�V	@��[͒��U�süqP&Ꮽ�UƧL��o�����T�����g"xɆ���"���g�)L��5�
�klb��Nժ���ﾈ/5-�n.�	�E�ڈ����r�����Ӹ�e�}�����{<�N�j%`��4�5�g*����7����J�,����US�m5�M�k��ŨN^�P��@$��;���eJ�;�?o�qS{Ƨ�����{�Ƚ2�]%e)�5k���k��hY��Qג\�K�E�Yb�Z��<%I��J�61
�9y���ûm��彈�U�0%P:T�5�D}J���\_pk��8���sĦ�|�.�MB�N�jbjNMط�U�|���[����]��s̸�]�Ju�g4u��§�fʘu ��FvASt�ճt� vP������n�B��a���@��*8n�7Κ<��V�۴���������=ב�W�}~؂������so��׫�8�#�s_W-OW�䍉�7���l��Ɵm�YQy��ޙ�X�&�#]>���N�.�n���YRN��ݧ����i�Tz�������"+Us�)��*)������)�%nd��O�e�����x�w`Sy^e�u1^��AL|Z���d\��J��٠��U|m��[�� ؍`�-�R��5i'd��Woc]��e����ۛ��lEVw5�X���, ���h�[=�ر�:�3l������^.E��B������<�:V%���S:H�v�u�U%�VE&{��R����ǒ���Hҍ��0l�\j�v�q�����g)�gp�JS
���Y������+���7z��eř1h�Ϋձ���Vւä]��,8\'v	�s���b�ڏ�7�����2;r*ś�Ȼ�ٸ��R�PS~�1a7aQ��ܖ�\:q�8Q�t>�����Q3��z��U�Y6m�%��f��e�t݂��ݘ
f��I�im�W;=�Қ����:[/���3^��ت/���~��j�Q�^�Gǻb]M�^�^8�����nK\�2+:Kޡ�SSDj�3[��_3��}��6��SqZ�s���ɝD�C��K[��$��]�x���ޮ���6d"�ePF���؃RD>��c-�z����xNi���Z�^AH���2&F+j�^(ٍa�Pu�F��5�7�"��坅bj��q�
������nʓ�]�m]8-]Ǧ$(dS�=P��oG�/7�.��U��X\����'o�)�%u!9)Zy���nU��tڢ9�yyY"n�������O��9Q,	w�*W
����(��J��<�e+��jORrp�z�u��6�:��(���7�gO}<|�6�H`�kM1�0]t(���"o��ّv�I����}B� l~����L��/%�ʀaO?7\�<r�2ŀ{���+����Q��^��/��i	*o���h��܅��S�=,)���^���N�N�U��� 5�1��I�p����ع�O*u����&��u��+��+������/
�ksټ���r�[����T>ٯi�}�����;q���2�E�W	�G)��ϲ��x�ӫ�DS�j����¹@[0b)O�9|�y/�*J��6�"�cD8n�WAl��^�S�Cvpv�ӰZ�ݭ��%��w$��$'����jI�;�A�@9 ^�g҅�j��,U��*�TM�P����p��5��f��P�@|t�3�TxWv]F�JОq���Q��p�~o�G5I΃'�5��<mܣ��E�ڠ� #�g�`�wOY�+�):�K(���<9=��Ү�t!A��l�G�{9!At��.��"�Q�~�4�CY����Ϯ�왽y�����JX��g`W+z� T�B�}jĉs�2�p�`�fU�]$#�+{0
ݮ�\��Z)n�)�TG���[ݺ�/8jC��d�jԻ]�נC��9���߭�����Y�)3M˞�#�݆)#"H�1�Y ��1��	(���D��B�&d�)2K��L4���΅���@I`QH(!6k���J�ɔBe��vJ�m�y�k��! ɓ�ݖh�dJ$N�t���!hNq#
P���d� %�(�0n먈d�M'.�A6�A�@�L�n�\�×	�	˦s� 5��1��Q"W� ɡ�%$�ljC�⒉$H��%$D�370��(����Lwtv�ܹJ��h�d���\ܺ���f��.\�$&%
T�Τ+�'w(]��H*QIH���Ax�x�!�0Ȯ\�ws���$L1  wWD�_� �TP�A��ՙ�aN'v� �z[��(�P���3�{�r�.���m�M���gnTt�Q
6�k�P��EB��T:Q�����S<����L�B����ځ��6��'�p:�|����K���C�o�f�k�{=''�Y��T��=Gj!<�\�������Zi��K�(t��=��i0}Kэ}Cf�9��s�o#���<CH��tb������(g�y�����Q��e�W۪'ꧮ�]\�s��w ց�.N�B���=�n�J���_Y�Q�9V����_<O���ުך6����E+�^b��^��e!T3�%A�֬b��-R�S�O�Y��=3}Rkw����'?Z�=/��F��J��O�0u1s.zL�k�P�1[��W�o-����7��)��m7� mm�]K��.�J��֢C�^���݊������o]�-,��5��v�r�u�֮u���*����g9H;�g�P�E�yq���M)}֘�OE�S6�+�{���V�T7�2e�k$�~�W�=�Kw�7�i�>�ھ�w��[{VF[
�5j/X)��!5:����G��y?Y��0���{�/�w��EN�u�wr���|�Nz��-\2'}�J���+4��=���=?	��)�7H%6�hߣﾈ��e�1ڲ��Br��ڎۥ������P��;M����<'�n�����Ř��Vk�V�g?*�%��=<�6��@b-G�����{����O��1]+�ͬ�2%vMb{���{W��V.֦���|�M>����N�spxg��T[Qy�2z9�~��Q[��#cY�U9���-�ɨ})�v�1�]Ao�¼�}B�]�v�+����6����t���O�}�踶���NrpkN�z��/+yj]�
9�'���[AC��m�~]�5����Jq�ƸՑ׵T�;��wwq�����h/z��=QZ�G>.���Wǔ.�F9��\���V�]���6���@��m⚌�͹�W�*��Y�X�v�>c�D�ꨩ}ܜ5Y{Z�9
�i��SͨO;u��Y�+7cjS��V�E�K|�^9;�ԍh�X�Z�*5�EjKw� ����F���/\�������$��~j��~y]��;��2���iFY���Q�|�9A��q����!�iGP��r�z6���t�M��b�xu�V�7�,>�m�\,��ᄤ�������yq�w��E�8�W��9����kF��8�ܖ�\{����8����beJ��܎Z.f;-TY�_g5Q�<����)�
�h�+`�nA�/��:�:K7�+;�/�eOA��i�W���s�q&�����3t�;3n]��Av�Y�4o1�(���,%W}��]��&��=��S�:�u.xr��]�-�����ʿ��r���sЛ����n�}tl>=8N��M��s|���O(�ЮT�0�@�k��g?$��v"�o%v�n۾�I]5��o�۞�p�!��.��e\�����l���*��n^Q�Gm6D۝[�"�ܼ�ݸ�y�M�6=�V·pUk�Ml���FVy\]����2ܱ��YQ��F�ڏ��*�P���
gղbHOC�[��$+��!�������f�U�+�mX=��o]��T� ��(�����%l)&b�峿�j'st�\`�k��;�j��}JNW���;���,>���R�"�2 @R��R0+N��I�ʰ�<�95I�N�)�(�f�ŋ�}w�����WC��m���%�&���yҵ�Ï�rҽ%�f`�G�}�\��n9��z7'��=_�	a�y��ߊ^ұj��3��D����"�!��uH�x��qz�Wя(�f��2�V�7�{9�<4۔���^c16���z.�l�q]����u�c��6hz�����_��������w���Sz�ΌZ��-m�܈m�r�x��+�<�Eg_�xl��o�˻�
�o&�:�8��r�7=�;ƚ܊y�Z���,Օ8��HK�������m}*խW�yU���J���ɵ��#�\K������J�O<ϥ�ڶ'��쨉Pbw��%ђ�>|�6.�|VG#�uB�5;��z���ﶥB����+Wysqv�GoY��E&���n�M�ҷ�3��9�<�X�S2W�]��Ȼ���Z��Z�Y�o]�.�}�J_u����T�Br�_�W��9�!��}]0W��GV֘Ԅ����'���ع	� ���0Ȏi������yo��q����[\�4����C���l钭t��ک\R�S�4�.&��`��n�ci*C�Y�;K}���z�^��><S��Ꮕ�Ǣ��r��՟�}��L�5;��� V�rc;���	��wN�����p�'f�އ;b�ʔ���U�T�0�|!��+.�'�p�Gs��w�8���s���M-�ҕn�
�ȗw���2�4yf���lC)r�5W�>so����
�}5�i��m��k�O}�T3�N��P�w��.ڣ�2�+�`{i��Ψǅ�-DL�J�էo��.t�*�b�P!x����h]���^ǧDM�}v
�[���D�y�渟���C�z��׶o��nzǪ,�b�R����8׌�J�n/���r�=5�WR��y���Όv���\���M{���7X��
�ڃ�u9�����c���3�۴�6a,庐�in�L��Iy�v�z{����qg�q�F(�Q��Bl^��["�EO�9����&oQ��^�.e����J��ڕ���=Pp�l^v�!�^8����i��uRT
S�/�k2�$.Y�.��^j� �
h�L���]�M+�����#9�FI�$;x�,�Ґ*kM,�k�X� #����R�oe��[3DZ�]X���v<
�G�W���Oy�ŷX�nb4�_t�	���T��p���ŷBP���v�R.��z�����}0WvZz_\=�Tk�nur��1�s�2뼟T}S:h~�iO-�[�	��S|�Y[i�T:;	Ιم�'NGo6��U��W�?SMb�V��i'���5�j��%܁#���~��]�R��`yC�,��Gݴ\�ޒw��5�k}���	���ლ��a�"�`j��*'����/��M)���>����n��[�RsGz�^�8�T�}�5�W��,>̅W ѳYKM��z��vgH[�r֟��_�W��W.b��v�W����!��2��Y��Q����&lVݸ���t���ث�����>�v=�zkc�sm�P���6�K�^ou�ӎ�p6���9��k5Q�=��4��SԥU��}��h������.�v�>�⾇��w/��97J�l������愻��i�.L&')��9��K�t<joJ9����F'�����Ǜ�\��\�cH������ZE#d�mIv9��ܗ$�!�n ��U�z>�d�����!��]l{a�m�x�����6Y������{�d �*��J�h.;G˷�m.�O�Eu7jU�)�*����~������[*'l���M><�fQp��+��L�F(�Z�(�+�b�0�#]���+�W��c[����{����*����X���� Fܾ�������prw;Z�[��Yy�|�z��TzƔ�ܲ���nWJԞ�mt	�_U���Ʀ��ۑM�q�1!]y�r~��u�>>���"�Q���kK�r��TE�V5�ќ�@�OsRo��*�Q���̇6�鼽�!k4pz;*TJ)�]+�>w�OC���NfMN��������s��U������*�%��.���]K���3.p�UM5�������N7/\�P�]�#���J�����s��رYSvrj��uc�T�wY�����P�j��bU���a��B�����Wn{YW�[
�x��8��c �s���C�8��YZ�7jn_=��Xs��l�m��n�&/�	U�چ{a59�LE��7TxYB��L��i�yU�o���.����!�TF��#����H�y���Us��A��'û�����I��Wc]L�5�<7s.4�K�����q�������Y��y��g�2m>|�7��^�9�8�f�s�æ���*�S{��!�
�E���w�y�Y���2�ٷ�x�<3��j;���B����1D������55v���B�0V\�F�T^b��g1��U#�����[=w]��V:�U�(s�p6��hQ��z˃�=�߯1���b�6�D�}��."D�u�IN�FC���i�b�hl�[�5�'�+�p7*�ʃ�����S9) ��K���(�׽ծ+�E�s��>k{]q߱�ʎxwl���Ɍ�j��	�C��M�����kZ��R���;n(�����L.������jw��@��[��ugE��_i���i�cMnSͻ��ы(u=yg��d��J� ���F�mJ��TY�V_;�T����Z�Kxwv�p^�8�s;N�bO�k{,u��}�����-�/���x�ׂX�1�W8q}}7����g�:,�B���o:c��ή���Z���1�eڧss�-ʽ�N��lr��.�@ެE�+�1s1�'�S⭗�f���ڭ	S�3�E�n4�/iM�徭]]/�vj�bP���Q;�/�Y)�e�.8֣��Ia��i+n{K�UsYO����z:���V�д*���R\�K�8l��t����$��=\���V�i���ۜ�br��;���(�W�iA3{1-GQ���N�a�e�N�J��5��phW�Sq�T�ͼ�<�zӐ��^��X�p���[X���葪�s�t�)�����{q��b�*2�v<A!3%#Za�A��&+��[��!VGs�j����z�Uu_>��Vd��,���}�T�)f���l9��8��m
sƊ��I�]�r���z*����)�t��6{6>�6��/1U�7��9�s#�
;K��m�_���5O���n�Nj8���Q���;��$�<��~�=$+��I�?;������j���;I����p6�#�h]	9��1��s����r�C1���i��鯠���-6��|���p�z)2�g��Fݣ�d��������cx}����buX��7:�:�r�U������	�ݬ_F: �J�PN� 31ӎĒ�����Tβ1�y�s��������P��{}��Ь_���-͢�m/y�����s��qt�^��64E����seR��V�����D�ڣ�K�{~~��E�f���Gw�h��v��!�+j�"X���=��6G��s�Q����T��;�'.(%�z^:�C�͜Ӝ|�om�P�ޓ~�rڥ<�F��m��C�~�!p����D��u%�y���F�{�6��o{⯲��L>��Ī�[ƢT9�+�O��[Z�f��7k��G����c���w��w��}�N04-����F�&^\ս����]�D]8�������W���}4����FOН?k��mR�s��=��=CGy����IrR�Qk�^.K��/��ա���U���f�f>j�Nj 'u�˗K�WO�j�f_z}5K��W0�P �M�\=.���ÄJ��8+����Y�W*c�kD+Q\�ya�c��T6s/�c���m�GפS�:&&^�]�굷����0�ڰI�jÃv9 ����a���ȅLmaB9h��x��Z��lp��Թ@<�|S�`�ijh�Uԫd��v4�̸8֍�OV�YEBzP�[�*�,5}ș� �HX�:�e��fZϔzh�8�ݎ�G�.�fM��G6����yIL��73�$��ض�w}�����Ch���i3'�]n����-J� e�+sh�oVe���mt۾�[���VB��荬�7�`MZ�cI�y'nod�K�t�^�X��+�2�\2c7ź�X�N�^m[Zb���/��DD��i���fw`ݪlg/Vu4�_���)���%,%HЗG6.D%҆R���Z���"�z�D/2N5��������F�x}�P���Ζ���zY�2:�ۥ�ڽ��Qƨn�b$!�nE2˺��o�W]�ZUjb���Rk��J,�X友r��]Gz��P{wm�@jP?o�r��G�����8�4��M )����q����9�N����u���oC�ya�&���X������5�˳;��)5}����1�J�n��:���.E���+�rP�P��IZ5h�Q�+�%\���h ��ʲp;X��@ua���_`}��3�U�ܓ8�J`�ݼf���*��P�2�w������q�f�M/�J9C��/��">Rǻڽ�O��88��j������g�5iX�qz��;b����*4#�d��o�ekPV
U�VS*iF�f�Y:�C`XƼ5�C=u�bE����WdRj1���| ����Fˇ���ʽFE37F��̔s:+����1 Gc�\���y۹O�k���3]Ž7�w�pnn�:ʲw�}u��8�8�p���,�2��OJ�U�˭�ˮ�8uJ�L�ޖ3n�tb֐�J�啩oN�ʣ�0������Y�Y����4'��uR��c�s�V\Cx�qW3�\6旙n�d��!V��c˳�w���f6T�(L�X�^��u�Sa�-}g�>~�#��rQ�ԧ�5z�'>A�z�-=��`�FrQk����=�gY���d����BN�l��9]��v�e���*���[�J,ʝ$&+�*��6M�&��]��+����Fq�G���t6�q��S �/��NN��u�b�r�R��؞'�m��۵c;��=��b& �Q�W\�n\�?u�� N�fIf�w��ݮ�TPۥn;c�d�m%y/e�#7�͚y�iX�x;Qf�[Wa�
i�p-��Xq��m������c�V�ų\n��C�w;^x�o"��w���R>��u�����R QW���{WP�D^�u����RV7��J<���1kK��Vqz�e=]-c���o[�r��v8��3���H�UۊʽX�;��l��o1�Qץ,�/-�
�3%A�+Rhe6*L��qo�hzU$����ue�Z��ڤ�DN@�y�Z�%���ɉ�`�SH�(b�H��P�JH���D���Da��`�L�d��i)1�����) ��)�	LdL�wY�$M�dD�(؊@�'��F�E%*D"B6T%!!I#B(a�n,�bJhf"`d�\ܔ�I�)!- �L�9у"P(y�$F��d��J4i�,lQ�D@�h�����d�#�#31!��L"0^v��"e&L`�fhT\�A��(�/�d1�,�S��LB�%�$)&"T��1�Jh���+� U���s�)֞X5�Y6���*tE�ٔ��ϒ��7�RM�
��$Xb�)EY�)��dN�˽�N�����cA���>�U�����,����+y�4�GT'�%[1?t��6��Cf�Y��{�;Z�y.�n����
�t���=����k>�>�f�g�R_Q[�?fV.�>c�7�-nW)�\cy{6���>�!զ���&�|��u�EZ��uI��fB�c7�_^c�y����9�+�q�C�����ˇ�w\��:�ܐo�4���u��GeA�u��Uv��}�/:���79sE)���v{��\��P�������2�9�ܨ.;*TqM�>Ŵ���*{'�����rNP^&V�~�+7�������ߗ�{<�dz�:�%\��gZ�����w6��.\�~��SX�ߋ�=ލUo���19�� ʗ��p�;�mkν��G������]�hjos�i��Rs�U��==�8Y*���.����}	�](T�5���Ԫ�*�,��j5;׼�e7��8w�G�Z�.WE��(�
����������˧i���{v�q:�+�lG���dr	���jI�x%��Qa�8:N��_�(��A;��r�����gr�6띾|w�@`�>�h�����ɯ!u��R`�����B�o��=k�㷝�%�)����y�����N���O��u��ؕGc���J)�]���>w�<ҧ�R{\��ٗ.�[e��5c�ڃ���)_�*�%��.i��]
,-��Wl�Ju�E��v�w+z2]�V9WT#�W��#�^�igc/���kw�bP�s��U���Z��y�dCc�}f���U�� G]�3�f�JR�{dnVzU8�~�}�'�9�lZ��*��U�1�7�4<ɶ2�os�mU>@�f;&��nM}���W1�˴�M5�u���\�M�])����DO*Pv��A]�i��[�<3��ڲ~ޠ�51[�UL��s.��{�֜��<�gFG6VY��)�D^b��f~ŀ�&]]�ʌwW����B�{[A�6��9M˿��,��o�ʼ�_^Nt�|s��b6km�ܷw��\^A�M_˧[�v�����z\vU�&�I�>�$T^w���C��e�x�h&�vT�4���ldtr�d(
�En�_f��ZU�t��� 9h�],ӻ!�_h[���	ydU޲�Z#yqGioP����3Z4�N����}�ѝV������f9�G��N�7Jb<��`X,����]ۖ�����dVuB�L�
�Fs��T�~���w�5���ͿF��gF:�Pb��w;z:%���M}�.y�=�zaaSŵ�lm<�T�9�ÊoǞ��\���{�Ǐ�^��!�YuѭC��\!��[�v�NXG��n����b��DE�v�oNV��-��'�eRޱU=��Z�}�!W}��{�f�����_��c���cC��='�t�3o[�s���G���~^��*-���(�v�Y\|�,���i�i��y\"�܍��&���n����k�����-���䭵�{f\�3���B���^>������V�wm������q�}��m���{��V�����0Fc�6*σ�w��_t��_w'�7�.�N���TƇٙ[�`f̈�g�h����+��zf�w�]�a4��m��:�m	�WG;i�W&Y;�	�a��s�]fMp1�2�y��0�ٳ{}���.�P��{�&��%e��E�񕓜������P��0ا��j�,��3A���GPlxCv:,/�dj�lb�6�3��������wzG�ǈٽ�牲��^������{y��3-rZ�����e67���ؓ���*�s���V·��\��џ�[G���b����2:��/HKuE:ޭv�&��N8O*�7�NC���OxBF�3�<����>��������!���./4Ց�AV��P1��W�U��Y�{s	���:'kn��Ozv��ǗiQ�ϝ��rC�*�C��Z�Q�f�\}�5Uj�\r�7���?|r�5}�b]��lޭs��he���v3�G6���v->���[^����+h.:qM�麺����e^�i%+3���3n��U=y��z��6�G���ڜ�g���8�\o�D:�SkUv.}W������s觻I��ק���ݍ���ֶ@�o7���'��o_J�\����֚�CZw��|T<������i��H�ʲoo����d?�lLV��2y��V�	�|�-�ڝ�uM�������
��X�h�&
ɳ��L��{2T��u'��&0m��1sj]���4������|�6��B����K-��Jl�;:�f+}��6����IBGq�U�J��:y���jS�����M>����J�p���E�(\&�j���!*�m�
��Dߠ(YQ=�n'��jo�]�R/�B�o�dQ�����l�lq�h,��L�����Ga�2:�dn������IP-{�<C�Ko��8-I�h�r�2�	}����	���w�'u�f<�K�6�̿�ֵ��9�\8ja�����iY��\J׆���R�2F���IwD�c�e�$��9�w�f��rvU1�!v٥�\�c�k*`�-���\�Wsy���ޠ�r힇����c��<&af�=�6gQ˖gt�{���c��_�S�}����>D�B��L�#�s��-QJ�� ;�)vٵ�y����j�sS�WN�Hq�*�fj�Q�.�>s;[Ѹ�bt��>U��1\:=Qm�O�
��c_WˡuL�Z�Tf��⠯��HoB�Ck��ڞ�k~��.:qM�>�>�n�������;mƬ��K��M�_$0�w0feVΫ�v�F��6�v��,�E��ܱ�u��	[��,��]�C��{%�]' ��Af&@�_���A�A�mw��̙�Z=o2�G[���FEs)IpIj����jz��7�m.�eI���(����Lo&�����������f�϶����ߧy䊨"��/�%�5����w��?S�t�����4���HU��r�jwٺ��,��J��O�se�=��M=�w���eoTY�a��qjoo��_nD7�we���C���(g.����o�d�z����VyW�W;�j5;؇��kuF��;�kyr�ؤ���x]Za�[p��Pz;+�P~��b�%FJ��s�~��k{��u�%�o�7}���춄��̧L�`�;�;���*pʓ��"y~���ѧ��������z1ܥ[�� `K�W�Үqג�{�z�����ӄ�Lސmv?C�r���O����zj&K�m������:���a�e��$�r�i����y�or�Q��=��ɾqG�W��o�Q���.�N�=ۀ�w�u�;�T>W�;r����̝���rc�@�J:�.v*���$Y��'��N�=�&�]ޜ�-�u]^ٲݡ窛]H�]ȬȮ�$%��^�	�vi���f�L��7ە_V�_��v=�ۃo��.���0�����|ݠ��0������[p������^�����䀝��1E�����sNc�W�rӯ{��"�~<�a]����6��/�xg�X�f�PGV��C�56���wtjy�_"�"E�����}ȣ̯�r����6��56�E]ڸ]!�5i9ƅ����K,��n ﲢ�ݥ!L�$���n��XҊ���\F8=ԝ��V��<�m��|+#\�.J�Y�6�;�O7�}[�َ/[������T�����k7�Y�iysz<M9u����駵l�/˻8��{X����yq������m�Ҕ��/.�����f)0v�eOR7�b���/�U�u���ZVT.o -����(�C6��i]��=�x�b*q��7���1	BxiQ�V�_Y�Qe��4`G �U���p��Y��z�5�)0�����bz���P~�ދ����*�N�-�y�8�8��\���\=��7�U�p;
�ZWã��ɢ8�#O��B��ޏ�\��1f�b�}jׅӷW�Ǔz�a����޸���7P�%d�hIQ��.ƥ+r+��`,]��(մ.�L�fK��q���'���[�{�6���@����0�X��cb�\2[�?n&��p]y x���f��������L���M��@ث�K���ҭ��P�)vk�r�D��v�š��f�����G*]�'Һ����(ܨ��Z�5}<WI\d�����ƫ��ɤw�5�u���=H�Z�-���|0%B5e}=2���/��.�:�%j�m(��}��5�u'4s�>�ws)c�iuP�,�e��i�$~�?M�Tܛ��5�[��U�/%!|��p�D»s��tf��}~�؂3���n{���]�'j����=v�bg�MCv�!�7;�d�=�7��Z�1���S/�NW�ﻴ�c�s�zBZ�:�M@����B��p:�4'��#o*_1�D��S�Nc������w���P{���t\43a5D*��'3�k�z�{���\_@wE�-��O�
��c_PٽNx�߭Z\U�zjp.���o���� �� ����.;���5Խ��J�C��j��XԷ�R�{��޽|	Ί��n���E�p�F�Vŋwa]�uT�n���Sv��d�zk�۫����y�7 |���r�W�u��]B2Fx�Ww�i��;��rl��%�#p��&�~� d}�#o���om�~��|�x��@�ӡ���o�B�V�'��.�f��Wq�ioGGSùI6*'ۛ��Ǔ����y�T	���W�Yz�kV�]h=;��
���s�R�kym��"��<�nC�}p�%O5$&]iu�f>r�/�蔢{�_d�;ˍ짎���نz
�Vx�0jkԑ�ʽ��6����P�쯥��R����*x�ҷ������j�����Y��m��6�u��;-w�QЯ$��
\��T+�P��v���{+5�ʊ��I��;V8��SIʗqT#�0�W@]�˯�},A�p�M��x�Ku�}�5ӭ�3�:��Y��Z1<�[qO�\��������J�0�2þ�ϾN������]�|1T����%�	݌�9��ħ_�jW)�V8�W�پ.e����aC�nf��4�UTLɓ32�TX�f��T�y�w#Io6��3q�L�u�K3,��b�s�S�E��e�8�_u��D5�zE���4���=�ш���9P;��A}�ٔ�¯r+8�oR�b��^�p���x>ppx�����M��ڭ̥gL4ۃ,_c���1lx�b�"�;9t�:n�}[�����jܙW4=e=�����uoL�,s_n=���4�uNF̉ڞ�2,��N&�(}^^��:;џ���)v��>vq4�����a)��e�omO,R(tV#��hY��\�.;*+�����bzRv��
�h��dUub�qC�Z�1�ٸx.c�vͬ�8��s��@:��	f����M(��ѝ�/>�Q\��O5F��X��;;�\^s����T��C�;�q8��o뗶1Z�X�w؋��o�%<�����e=Gv7���o-/�DJS}J��+�#��c�i��S|�BE��R�q�{%e�9*�\c��[ƾ�u����z�P����Jc�c��1*�sԐ/iM�実�y��hZ�=�Ge}�R��|���2)���j����G���J�s��~������)t	T�ʒ�
\7q,\�c۱Δq�#�eGV;�=;�jژ�Y���v5�&�MV1c���kkr��LC�qo˭F1��g,V"=\ؽ�sx��;����[�����1��2k 7"�t�}έLE��9Bb�8j��͑�u�U�&��OI���^�,���ǿ3��K#�b���|'�u~��U{w��(��WM���#¹�7�n�����ܺ�F���AƜ��o�����f+��C���6�,qv�P7v�K�#�ݖ�ҵ.�������2�;s��v�U��hK�z)b����L��X,]�P�ܸ�KCyY4:�����RA��QJ���E�����]�����jh��=����[���aP5Ǳ(��y���G;�'v� ߖd�>�����t���W��y��@�3AUWa4���ӵC��ݚZ�g��"�B����Q44�H�w�a��b0(�s�љK�h˾a{���(���
V��,�8��=�i�=}N�vr��l�9��Vv�i�E���.�e��yJ��s�����x

�(ك�v�yF6�gǷ�ڭc��oS��9�w��:��d y�S�t�y���ŗ��a�-���ǅ�뜽ӊ�s��\�+�����S�f:$�y)�	�	�-�V#�V����6H�0�]��=���\4��D�c���P�B����~��<���4f��S'0�R�f���Z�c��G;��;�n�/*M~i�2��(ssP,�,�Ջ��4�V
u�C�]@{IO.�GӍ�N�X
x��F��3ܭ�����s@��_*;O!N*as{0�8W܁�S� ֖T���4l�{=��`-)]&�oe�-�"��"ʥ�(���#b�����ghY{�7�`�`��rZ�M^������4mB^�Ӝ�f=� �P��6훢��퐖��h���,��|5�bpYV���}������c��dm4E�51=�*Y�dh�ϩӽKo�ڌ�v�c>���3�p������i�5.1G��<=_E�%�oc�<�bp�[b�e4���Ӝ�8^-��;U�4;��j��hh���uX��{R� �Q�.v=�vSH�μ��S�S�u9o�Ȇ�����5�'=�����%�fm��E�F�&:��,���OW;�VvWj
A�f�:��eܾ���hr�ζ&/z^$j�(R��@v�!2~U�2$2�2�
6��e��*��[�]�Mp��9�j�c�i��mV��s ����҃o��m6� asw U&$���F�\�K]/I�8t�D��]Y�yw�(���ŕ�ν�ՄR�קn�.�5�R�@�CX[�]��+�4%[��{<��ޜ������R����Cힰ���t�(%�ޓ[W�"���ו�T��P*a��e��sU�ыnI]V��u՗OwK����ᒀ�Iu��ٵhv��j �Y�z\	K��a-��rۆ�e2R��ahy����9�խ���VŌ�@
���
l�ci%"� ��w(
I �1	����60�]4Q$hMIAh�@B�IB�"�0�Lȑ�DD�6 �� �v��Q(�`���Lh�(B�/)��HƂ�6\�hę˖� c�1���0,i$�L4󫉣E �$cP�&�d��R�&)32k�L1���,I&I4�)��&H2D�)
��,V#PF#x��lX����E�,@Y"�.��M%��&6�F(�DTb�ěH( (��>:���ʽ�$��/������ժ7��`��aO�����1e�Hv9�宝HCt�^�ƺ���� ����r��;�z�%K�.S\��4��Ԟ�؇t�n�JDjK<��S�l����G�{m�{�IVڻ���.�P�_\'��Ѫ�Y�W*{��y���מ�S9(�� l�\��bV������'?%��ʦ�ZP��N,�7��";1FZ֔�b�L8�#�+Ȋ`�+rkݰ�w�u�5�7�m�Op���y⩾����K43ѐy|�|�R���������&-{5YW��9Q�b���.-5Oa"y�������R�7ou6_{4��,g���//A�\E������1������+���&}s�>Xx�YN�V����ozr�Ɓ����\m��8�3��ww��n ����3Z��uK�NwE��b�^���>�3�Ou�N����+3�h�V�#�=��Gn�?|Zf���k8�]��v�R�~(��ߏ6.{�ݨ��A��T�Ư���h����QԲ�fe�r"�+�C��U�R�Sz�5~Z�^���V�b�[�;D�D���ʕ�v�;��n:�i=b��ꏑzɢ �>�̃��˜U�7Y�=o�x䂾<1�9��3�+9r��CB���[[���!j_�3u�$�%|�&�����B��NW�K��4�9t�Z�Q3��&�*������W�s/F:]F�{���*�M�o�`��K�����W�S�m5�M�|U�U�.����vWҡ�ϗ$���6�3Z�P�{z�[��>v:Z���K^�����Ǟ�R����ģ�z��#�F����I�+P���t�+{5�4�|;s���N�B:��u�m��_ :��@��@�YRz~<��.wq�U������A��k��85,H�gr���w��r�UTK*'�B�w�]�	�%�1�n�.0�4��'tnD�zs����C�2�T�su����V��wy�p��͎m>���T����֚��i3I�B����t������`�:j�p��֤����P�iz�Ϝ���wz�a5��z������٧��S.*�wh�͔b�f�\p�r�L��o��Gӭ.2�_U��m���v�����Q�Me�>���ۡ.�K� ^
@����j�I,�)���a�u����F�샏���/3�_�o]Or��T�s��m<�;�OI����c)s���
�5Pw�:�z��I�V1f��զ���a�y��{g{*/1�^=�z��M�F�+�褕�GgOT������;����ޫgG�-���V-]�6�V������"�%����V:�����fo���vG>���SO��R�^ �:���i��<��O�2�7�y��9��^A�!�C�\9�.��cn��nT���>Q}������vB��d�iW��%���/u�sNٹS����T/k�3��W�뗧��Σy2�yΨ;�t��FG����߫�ܼW��>1�糂�=�׽��}�\�]�G����.n*�<���L�ڨ^���1��?g��Ǳ��;c7���X�H�y�i(�*>�C�;ޓꞂx���8܁�jW��چ�C�uǡ�[,��;������af)�=���u�����g�mK/�no�Pf⌏TD�h-b�j>Q֓��"c �/ˢ(��]����s	De�D {�Mɗ�OLl0�تvMq���W��.n�oM�c:�}n
M����Cp�1��665NQ����<�K��P&5�PܿvP憧iW��"�{ވ&z�t-Բ&	��2�7��H�#��T�>���[m���K/Ǵ��e��p�U�/ l�ٿ���*��7�͎7֪3+j(�_��]�ez�>Ī+�u��#�;ģ��'����r)�S��>g�LL=���ڪ���v�r�{�H������zV���{	z��z�_�3Ӵ�3�w\���m<��:���
��u�����7蛨��e2bb)*�;���i��]W%��������S�6E/rO�Bf̬�O��&l�	>��`�MSGr'*=���a秤�iz}]>7��b��r��G��[8_�6�$�ex�GMP�qΚ"��J9q��]�p{M�n�;ͯq���ﶡ��%�#������SEW�z9�O�҆3�?m�{ڜ7�z$���i���3=8FN��W�����[T�_��F�ϙ�'�V�<ٜ�Gy�F�۷o�s���n}���1�#�ܻ����?fv���=�sO	���#}7X��@�ίg��O����}�<a{���F3ڠ�w�-��`�B�(��Uh�ɭ,\FL�7�@��G�~ζ��y��m�^��\�q����A��h�W�c��b�ZB��l��(��g���Z7�;q�q��~l\�WCr��D����g�	�~�N?N��a]�<��;�Z�Jt;8\�jv����Gr��fؤj_tE��Y���v�̱�8�^�/^�M\:�į�cҼ���~5��ɝf�ɟ�ю�~�q��;�+�x����ޙ��3O��Vma�
�֍����
�n$�jnjި{�S7�L��r9�C�B�o�.:���������k�O����W�[��B����¶��ϡ���pe �n(�&��s�坊/{<���ws��|��M�Ci<�ȉ^��G��Zo�o��}���J�����@Jd�!�8zr��,�V3��N��B�9͟_[W�n!�[f2<��ϸ�=�p���E���n��Br��~^�r�s��y��1�;�YF�h�8}+�3g�S�hU�^,lA��.s�x��N\P���;�=�;"��7���Fx1+��̢c"�W�����ǫ�n�>�W���W0��?l�j�/-�����Ȑ�T��B�=�2�Q~����~=�&��^�Qp����>3���*7B|��<���G�� �#΀�~�7\NDσ�3a���h�~���������3�	����W[�����>��7�6n��s�UZ=��)z}%��Z{����ͭk�^��Y��
��mYW�/3��K����V�ݥ���d�n�%\'��sηo���p9�o)�GdX��D�0��0�!R��)�k�p����g�3��W���*���=O2�&�$��z��dV�43���Y��u�]���e���f������Y��Q��wqr�o�u~�3��pfkY/ƫ�4�9�L^��G����o��aϿ�YzO���w���� 5�������xe��w�g���.�'Ei��Kk��	_�<����J���M	O*p��JQ�h����5����3��Yܫ�A��e���k�����͚Ӭ��莦�+�@ϗ����N���t�a��ƽ����bG���5����i�9�T�;790�#=]gYuH���v�R��ډ�����`�V'=櫂��8dw��rK;�3�M�CՊ����n#�&^*�עG�dfn㞯o`�`^Z���ީ�}���Q�����q�F�"����늦�����e�S�M��P�z�}/5G��ǾS:�����:���z_�Go��n^+�Ϛ�V}�"�(��=�N����hle^���ɡ� �>�*.w��mK�����G��Q���'Jy�\@]R�u��{����ڐ���R۪��g̢o�+���a��Zg�鋏p����#NUDz�^A���/)SҺ2.�Z��fa��|������B+԰��������4/�^�����������Mm'�m?�T5�z�s�2Hӏ��� ?f$��O�u�)ӗ�\֍��U�s�UD%�}EZ�0���X�n��;%#-�7��N�N�׽V�\A��2�m�z��q_ �<�KJ����9���p(uZ��{Zu7�aȭd��q�Y��`���dp�����j'�o�@Of�M
�����g@�~3{z�����!����j������9�U����{v�<�tF���D��ڵDS=�+���"yIʚ�[���ļ-�Ly��-���Is�~��̯QG �CG�')���N��_�z��3s����鑌��1�X�y\�CȎu�Ɍ��@��ǘ�B�W��;�<3��?drVe����~�r���O_�,t��s��}�ǫ�Y,\s��~tM����]���d�۾y�����=�g@�a�r���z���V�q�^�}��f��`���$�ψ?|�nN���&U]渽�F�����n�25Ĝ!���NT,7����i����l�gO���5�Ⱦ��M�
��3Uo�:����(r�{����Y�n��Ǟ�~Z�*���`UG!��\��@mϣjxm���[��T��"����q{o�ȇ�Gi�)�T�w��P&K���wˡ���r�㌏m�^�{i��;~��?k�����(�9%�.���JY��1�hN�sv���ц��pl��Q5�HUdj^~���ƈmZ:W.��Ƌ���f���T��~l�s=}�tԈ,8o5�Ɏ�6�x]��/���y>�/�t�3���H��r-�u���-�l��[�#��nc��ߛ�_��KKY�ɟ"�9�	O�to�����/ƾ���_�R�ξ�4��d���ܿCl�����B��M����`Q�@���)���P�:_t�^�p/N�Y�F�z�s�s2��X=!z#k/G���Q�½f��ۉ�p&��*-J�u�Pѧ��x��Zf��o��{}2r��3䐯���B�z�,�˦^��8�h��}-�G�Pj���顄ϷR�����h���w:��s��(�s�p��t��KCd�ȁ���*�F�����9fO�����^��<;Ng����J�o�]~�����(��>q��E�9�$
^�Y�=���F�b���.�w��z/�l�El�tV�c*��쏽T����霏T�o�t�u��?*�����S���(����~�@�e	�ɺ���W������q�|;� K]������s���o���:Y���� /�r�
}�3h�e��u�2�L;�=]&�K�꾯�S
�QU�&e����x�
�Gݾ�Ϝ��g���%��x.ǰ�f�C������V�~��T̜����3�1S��6�ѧ��&f�J�$�l���5y"z��f=�6�`�Q�����ٕ�D����*����k �%�K\A'S�u�B�����X�=(h��!"�����jw:����w^t.�3/z���W�Gڤ��g�ne�g��]�##���P�����:k�z$���i���c/=Z�^׽�u����3,4�le �G��8�]3||ūyl�x��Ί;�ʉ؇��p��N���Jv�����.&v��A+�{�f�}y(V������'�*"�{=<�S����k6��9S��Oɷ�}z��"�t��d֖0���� k�#�}M�-)��86ǯ�f�Au���W�����D�^���r�_�tSg>��OL����t��L�7�>	�u:1��?_����j�紏�/v�>�r�xw�=�8o���L�Q&�SMCb����n2e��@~�W�p+zk1�Bzlָ�eu�9��e�_�Å�J�~mK=��DS�2�[7XM�z���^Fr7Co�b�%�nW��y\{ /Sg=�|W�K�O���mK.4��PT�����FAC��|�M������&�x&w6XU�b����ӽ|���3�w {i��}1tu\��5��˫U"�"�ɝ��|�Ð\����T�Zp����\�H�8g��7���;��۝�ee�6\I�-4&h�����R��ŋ�y8��|2�1;�ib\���yX�k�M��F�t�&���EIvz/9k=:dT1�[����RեY��=9�xn�&�S�ZP�V����*�1f��;z�$@r���U�ˉ�ϒm��u����zǄ�D&Q1/g�\���,z�n�>�:�<���a~�mm��o�[�wY�z4� �#����u���s�2�~2�Vѽ/ǻ�«aܽ����cݿ!��Hlfl�,���sZ W�`T<�]"r"j�a�m�m�ӲEc�ک�����8�{�=\n��ϸߕ��_�նo��� ���Wg�֒ǉv*|7����V]fw�������T���_�g�*�5��f����Ww�����8��ߪ�y������!���r�����z�׼��h�O���6���*�tV��}>j6��Y���Nw��������^
q~�	����ʯ5��U��cpk�r$�;s�ˌ�qb�f�޹}q���4�	{oȗT��K5oޘ�;�Y�O���{GE~c߻rؑ{�5��=5�rHêf��ڇy��7�@�}R<6:�g���9�����*�'Ϻ��.�������mܒ���=7EWخ��L�lq;P���{���:=�Dt���~ӛ�~/��������Uƺ"��Ph:����6? ��꾎)�C݂��h��)��@=�)s�4�ɴ��Z���My�&8&��	r̕:�Ұ�f����ǈ\��lŗC�M��g��xKv5����跽lU[t�w@�	�2Rt��`���Hp����\�ބ��Ӎ��ޱm�V�%A�+0��4ճY^w�qH��-�M�r�����������,�>�W�4)M�!��w��0�p>UܷSFe�&��2���X��P�u��_
ŋr�-�c-�|��J��jO��oW����\W�w���x��V�j��i����[4��i�ғl�(���n^��86�'+)�5)��W�{G]�j�@3���ջ0�.��Ǔ�E�'���a1�����>d�VT1�2���7�8��/Vf�W1�Ps��FȤ�F�R=nP+:JγV�W��9�P�j���<���B��٩�U��A��,���4P�D��Kij�c{r���-0]�j���F�$lU���� ��yM^L���u��q��t�"n��&ڄ_k�5�T���H���^_*E�k~X�{^6���z���\��2�fy�zx�w���JZ��ޤ_s�ix���wq-���99+��ElJJ�1
��F��E�v+��żәޕ? w\�𛝒�g��I����Uw�@�����n�n܆L�$�^�O��>��]dV��Z$-��&�ī���
ʲr=�CE8�p�ݳ�ۙw"�"K�V%���:� ��gP�p�� b��{�Sm�.��1��w�|ã��b%�Y���5���[-��Ef��t��5��,��pT�b���=ĆEr�v��O�){���K��ξr�0ě�Q�D�&�@�@� ��ﳔP���*����,�ו�mCr���j藤�u�]��V���j��y�3�u�=�@5��@J`T��	�?�{�<�6=��verN�ޕؕe�Y���G++�E�(LK:ۮ�W��v�a�I�#�2jJ�n;/N��5ί2�-��-v���p+%�y��Wl�3Jr������%IqX�f��'��]`���a��i8P��ū���AX�&n����U���QW7�D����r�b'Wg��a�*9��{Y��=�Ӈu��JǗ�L�U�S,�ՙG��48�p��u����_"Uθ�f����=��eh�H�P����E�t52GE��uq�6`}HJ#��e�������V�S�I��s&O>��2��Vu\��͔��Vuw��� .�HgM)��&���>K��r��)&�dQ���P�� �(-����=7�W���~E�ؕ �j)�d��?+�u�J(�K3J��F������q��twp��c�5 ����іitM�s �Tt�VQ����](q�اLt��iێ'q�����?��{��߯�ȋb7��j"� �F����ɥ*dh����\(т��.F�݃Q%�ʊB���^7(ѱ�۝ 4h�Y"ƒ�5wuD�Rh�z��h�4DI��W6wr�m)�+�r��ٛzj梞u�i"I(��#FH�)�Oe��r��1�6��%Ő�2%݋�#���W-�b���$��]�F�.m�
ɒ���;�ҝ�sL�Q2�UˆL!%b�)빼p69�Lld��h���b�.����wU�6��"ذV9��r޻�(���\�5ȃPQS������{���"z��t��_`G(^�F�aa��쇭���8,�F�S���C:!}o������Y�4۵c�'�:@��ɑ,�]��o%����锦/&R��2��}��W��QF���j�*�=DR+�n�z�hǎ����Z��o@�~�� ��#"���ږ=q��CЏ�������>�r��/s6��2��m�p���\zl��r�7�Rۊ����&��+��F�
��b3��L\{���w�=)����w9��!���� ^z�[4O@nd�
��(���#j�yi��G�1E�TO�� /фO��GwR����t/����<'�@<��4*��9��/.�9*��WW��wU�x}�޸���Z���?W�{v�
��䊈^����L��D=�oƽn�=���;J+��Pi�Na���$�G��U��:Ϥ��t?m�O2�JNMT4{G��&N���c�X�$����h�_\�27�>�\�\;�����/�~v<�d�T2����l�M[��:��7G�7<�dD�G��oC��|:M}�t��=Qʬ�.9��������%�z�#�=ǯ1y	��;V`{B�iېE?@���'��{>����en�w�m{��zx��`	����䋏p���֔(�V�5Bk.Q��s{��.'������\��fٍ��������_&�#	�Lv�׌�[>��t�)T��������Vi�~��]C�K^J����ů싢{a���7D�o���:
��GgB$����wN+��/�v�{��<���h�&Q���շbG��Z/�x����;N�<7�ꇛ3�~��zyyArb�i��{ky�܊� =s�~�e��<k��u͟ߘ�f��܂,��i�X�֊�k�D�F}�3�6������\�O�4�鿸�Yް*-:��~��o��W�ʞ)�Ν'�Z
���0)N*ѯ;W�(��������'\�Dk���#ٰ��<�����_�T>��\�>�w�f����k�uIe���f�~�@M�2���dϑyΨ8���:�=���9#�~A�W��b�+������F�L�I�*fX<�~��϶��K��~�?x1��^��[�����ǹ�[,o�Re�>����l�ۚ�b��*-J�u�P��tGy����˩�G-gU�F�oRg=�|d{������2 ��e��d�  Nё��bl��U�}����<J<ٷ���y�Ts��T?UOg���_�Fze����"g;���Y
�������P�P�;�0=�4�ƟuD�]~��L��?I��ۗ"�yT�/���w���V��Nw��+�BG�#{)�:��c�h���4/2KZ����������.�;_m���u�*B�g���,]_�G�<�:5��F�]���Ϸ�h�P�V-����i-ε2�ww)W�P�q�Ѹ��Ȗu��ά�ǌG��k��KiH�*H�=�<NS�gFJӹ�/
��c�=T�/�_�n#����I��������f�T�/���=���t�ǻc+���U�o\�w`�2�U���ߪ�j��@ �#nw��G��F�JvN �� /_��&g�uNT=���L;�WI���>��r��y��g��q-���S��`��>9��� ����_�&�גQ˟W��b���{^4���ߗ�K]���qg���픛���&}�Tyz��uG�_��bx��Tz�ʔn#�Q��a؉�c~g7��z˿c�o9���r��q��t��ū�G�3� /��y��n+�M�^�=�띣~zT���򷔞�a�P���2kO^O�i�Fzz8�6��j���~~�F�ڮ&���X�Q�7����§,/N��Fv����Hë"����������޹X���l����u�`S> ���}-mw��0�;��v��Zf27�nJ�z�*���+�0�g�ɟ�H�r��͎u�����QT�}ܫ��߫�\K�CF|�ƐY�ӛ�a)����w�yX���YQU?!����*�ˋw-_줽f��Skz��f;�4q�;��Xf�@T�,�$n�'$G_��M�B�p��i�O'���o��E|�h׹��0P%ػ�\��àAݖfֳ1.��'%e��&�W�_G�Zks����f�yI�D���nH��X��RQ����,�w9z��~�+��z�<��[�����E;�<ٸ���0���߮{R.�j;�r�^��J��G�}�~�����W�_�g��,�e�������������띥�/f���UHʉuȜ>g�,*����~��g��.ߎ��5�����'/*Qz�Ξ���X����xق�۪�x�;��̍�O�W��Pȇ�\�G�����{*3�����H����,O���(���� >���,z����l�\�Qjz}K.�o�uw��;Hd/{�ܸ�_<�M��TZ�ȉ���1������_�pύ�����4�FW��Q�>8��}�����Fp��P���>����m�m� �vͥ^�v�}r}�g��q���b���s��/�@��G��v�^>�;�Mׂ�g�
��=�r�����t{ݻ�����~?,~�<�á�m���i̟L8����V�c;Sd�`���UߪD�,����Z�?W�f�8S;�z��ͭ���Zo\�k��~��ƫ}�3ʜ�z�~�8�����' �ξ�3ß4=|}�Ѻ�`vz���r�G�e�O@��D5 ��Zo,.�Z�����2��'.�C]WR�=�f�F�MO�9��j53C�7��N+��#6';7TR�G�M:��nu��`�EL�q�~.9b����FV��ٕ8c��	�'�#��/+�X�͚�q�@�_�L	�W���4����'=��9��[��'���O��/i��|E�]UN�=��u��#\��-�č�ƨb��8�Y{у��X���{գ�/m�ý�P_=�,�D�=7Eb�����#^�w�Z�C����>��k��9��~>]~��m�]�dr�����������ԉp)ܚ�Ǘ��{ �Sێ�|�:#'Լy�u�9��/ţ���%ڨ�k�YIy�ef
ູ�$L��,���r۪@MO2*��ͩc����1y
����2����#��O���_8Ev,+}^�w�;>q.�A�+���l�Q{�<�i���y����O#��N�x��UD{���#�pǊ�M���[�%@{uR��z�>��jX|�^���\�,���G���4=޾�x�l�[�P��{,d9f��$�� 7����D��3�b�}���ލ��ϗG�6�&7�}�W:���zv����~ݹ*�k�|Z&�H��{j�k���r�����aض�xw>�t�(�����Y�Y��ǽ,��D�1c���˵:f�佾_63]���(Z��rwkO.͠_ǻjka���4���ü��9��W�NZ� ;�x�k���0G%�V�*��J}'v��5"������ςC=
Gt��:��G�#�W~9�g�v#մ�:~�{2ꈾ��߲;%�K �nߙ�z��#���z1Q
�V����^����m׍�\?:S�:���f��vv�����G�Tr��}�NO��ܴ{'*=��V�w>&�΃;�Ǒ�Xq·�*�����g�{�|�#*}���~go��'���OT{n2�L;ͯq�����m0z7LO��ִW@�A��\�R�G������}NO?eP�uߘ�f���9�o�5�k�_�׊{�{�9�uNa������|_k[��Q��F� &"�g�Ns�_���Y��ȷ�5�׽�H����nvXĨ�)L:Q�����kc7ў�NΆz{��mg;�:��~��n�\M���{R;��>}�K�^�ݰ
b(��^��Q5�^L��Br�ώ�^�k�s���=Ɵ������h��=�욼��zQ�f��h�NN��Sb.{ŋ�ɝf�gȼ�T�����yϑ�|�5w�s9|��^n�Rn3 9D��F{��ao��*M��e�'��ҙ���������b�c�/0:�����7F��ӫۑ�lu"�Es£}�����ȫ�`1�@^�/����
��Y} q)[��D�>>��׫�Qk
�����Ƞ/W���Ö����f���&��82:g�fH»�I��<��^ ���M��7Yғh#�}��K�����E^��.���qu��G�  lMC�M��Z���|Tu�Z�>����=g�z�C=���>������/%Qe������f��#֟8�P����Z9--�"�"6��մ�&�u�H�C��S9���N�lC�W����Ce���.�;5���+{Dx��V�
�;<�d��Dl��X�Ȝt��o�ģo�t������צ��il�{�v}�� y�0�&)�x�Ϗ�i�^��C��W���_)xi��{��4}���Ov���f�Rz��@����Qײ[�M'�x̪�O���r�,E9��� e%>�i��n����z�ٸ����z�4�艪�<na��a�ў�����	��#$����z��䇬h�fد���7��<����t��Qˉ�x.ǰ�dÞ�� ��x
*�ײw;���i�L�mBf�o2�9���҆��樣_w�Os���>�>�겋��J�V�'����ҙ�7Ł6��ϛ��9�s�٬5����Ҳs�ŕ�]_��#�_���}|�f�Ϧ���)�x��v1���b��)Bf+z�1b^��Q�2��4^�`P���F����v���[�ذ�e[|76rE��/FY���=Q`��Ԛ�[W[""7���^�U��h������qH;����F�b�t���a��gw$�����,�r'�nv�ˌ�ү�+Mƹ鸎�`n�p;�_����319��LJ"m��7��}���/�u�1���O���U1�gK�;�z�w�#۝M�;%wO��?A][�r�v���z��uǽ��g{�Q�{��9���6���+�.2gY���O1�O*�S=Y�]y,��]m��:�=�rǋ�����tiI����`LWz����z�������Q�x�L�h�{*��^��+�s��~\�V�|VԳ��DS�(��t.~��w)8ք�N����6�W�;�/L�����=�B�6o��Gţ�>����/�+.�qR���&�GGv��H)]��^ >�!dO�ț��<���,+j�O7�l�}ARg�HϾ���Tk�U��3���!b�������gi�b�:%
0t,���0N���T�7�,+�ᴪ��	�I�^���ӻ�[�s�z_���Bz*��f�\	�"&Q1����	h���%�vd�엢�=^��\�X�Qcgf�g%�~��{w"EC����U��&@zj/�iS��e,��O�Ɯ�يZ����3��,f�q/���]�����b�Fh�O� �Y��ȭ�ǟ�Y��1�QE����`�8M6T��bt�Wkm�=يxZ:������S��Xb�S3wPyq��=a)��JuL�2���lr]���Ln׍x(�)� {��h[��ۆ��3���c�F��o~����/9�]�$|-~�Mx6��z�����b��?Y�p��"�g���������=�{�]gg�>��}�=l����c�O=lfk�6rF����Ϧ3�$�~�c��w�&�}^m'q�F7�̓����t�/Ig������o't��tV��\�j6���#�>j��Nc��T�V�����9;`{�ϳv�M���j~�����|y^-o�=e<��X�t���Τv�۷�}��>�����|O�v����*3�kE�i��O�a�3��mC�OQ���c2���y(lY�6�Hў�����ߎ�}��{m�2�{�Y��g����!��Ğ ���םЕ����/����e���~ӟo���ؿ\o�|���l�+>�DS�骏S������e��`�EV�?_���L�1y3��ĝX���w�9/��i�X�6n��FBG|$�vfw��-9����F�T���SȊ��-���c���C������k�I}Qy�r�C�d�#�r����i:{g�M��׋����������wc ���8�r��T�-�-�r�9�l��@�n!�ѵ.��R�sC�`\�3r�>Ѯ9¢����y)7�]���	,�����d�e޺G��R>�{����éŃҏ�q\{���;>|)���j�z�e�Y�)y��
�w�&)��o�e�j��U]�=Ӕ����%����;�yD���A*۪��J�, 4}mY}Sx�,�=}�>�^���(\C�RG��/#�dp�����n�@�>spH�n)M��ّ�G����ڭA�n��wrǼjJ⭻Y�9�H�x� �Q���G�ȩ������+��B��ｃ��El�;��x���K£��+��L�>��$��`\o{6(O��mS��!z�e�����w�9Lm稏YZdc9��,m��7�϶����.��_d������B������+�*J�sr����{y[��FO�I�tݦ=Q��b������w��^��u�W��P�F�v|���c;r�@*���Q=Q���0�6�Ǽx�[
����u��SjKu�=�C���������ݘ(<���T�ܙ�t�ó��p����	�1~�R�*]�}K�W����#���*t�^����A�Y��ȷ�5�׶��d���3�F�C}uE���5t���gLβ9f_����ԇd�_c����c[��;��^桹��iO�eW̑���S��ZS�Y�	�����0V+ujq�vG�e'`��E
��ߗj����S�p�7 ��P�P��;��Үm��r�K�C����*iWE�z�5�[x.��X�V��Ys�z`<�?r�Y���s����GX�HH��`�����4�]'�S���<�v��Ҝ�YG�n�q7�l��[���H� vKi=2e�����ʄ�&������f���i-�ģ�Պ��fl����!z�S+�Y��&8
(_ܰ1�J���g	|M8Շ��v���P�El�{��^�S��[k{��w=��To1����x.���t���/+T�
Z��DY����w���38�ˢvv��)vJ*�^SX��ۋ�oD���D���dұF{�9�O��D�pt鞌tu�����M�|M(�l�d^+�+R���x�]piP[xmM@�=�� ��g ���]���dtٻ�8�5s�Y���oq,�n%(r�D��6��N����e+�P���b,�S���4k���j�)TΣlP�������X��}�/���
���J�x&'eQb gǕ�U�A�����,k"���u��4�{t�3��u���!9Py��Jک�X�50�ނ�;c��CLZ��ZN��~�$�Y����X�y>}�5jTy��񗦖mH���fnj{��-��0�[�T U��K��$T�{��m�I��!�u�2)�P��2�b��XQ̭K��f)36�#/_�w�f�wt)0��'����+ट6:E�k��ds9ϡ�L���4�4���[�����a�$�P�+OC`!�tȆ�:C�$���n�cwfն����)��,u�c����*�I+s'���ڍ�m��(j�K3E;���h}�P�W#p��q�Mu�+ �ݗ{]���-A{BA����������X02�	�ˁ�����fMW�_U{�N�Qn���[
a�\�s#�3��Bz5�A9+$�Q��*�n��Fn=�B�o�#[W��(K���눤���b��;����_fj��MJ�:؍�x�,q��o����wg!�{��y]ޥPJ.���۲�
ɫTl�s����t7�&е�ѓv��:�R'6E�p��}�Z�1����V�9��G��^��w�X���w���ES��wE�L���/_Y�)顎���6dը��6/�k{x����ۧ;)�V���y�E��"<C�h|��y�nЅv'���,�����:�KASq�#lT�GXA6�g�����kq��օ��8�xjhbY�;�6ossF%����KsXZaJw�Qw'�V�B���s��s��+�@�r�-t�������^wbɢ6���-�й�[��\�s\��Wwmnm��-wh�B�#�ѫ���s�-;΋E:�sm��n&�*D�W��6��r#i,E%���ۜە;�;��cT���̒���X�s��6�\5%��<�Ex��A��jw[�s�-�w+�ͥ���m�y�srMu޼��v�ܓQdJ7-�h���[�;�4��s�znx��ntwb�4.]s��v�W5�ۜ�5��$w]��sE�\܍����"�>�@�> 6U�ģ����	�Z8�{*�tp2+�	L��c�ˣUu�>#R
��g�*Mٱ>_fKx�Y2_t�9؂Q��ٕһG~�����Ǯ2Z�������6���[����9��G^�vR,��p��svV���W��%�}:�A�EW�Td֟^L�/�r��#�m{<Ƕ�����*�E� ���J����uk�K��������D��=2���,,��o&|�Ϲ�c��:)�7Bzҩ�������B_3������w�'�9g�R7m�3,����ҙ��������LvK�����Y��Οk<����ýX=�����J�yH1���v?Q���(�a�Ȧ�B�Gr�K�0�ģ�(�yT$i=�ȼ~�����.Ͻ�F�����dA��L����<r6[���zٚ��W�%WYX=#e`>��^��Pѫi\M��֑��(�s�'E{-�~�����"$��������dft竪�-�XZs#e��J�{�����9ģC���b��e9��rR���R@���Dw�*D�E9�Ҵ�@,e%�C��~��i��_1z-�[}�T%u���Ny\Ͼڝ\{ۑ4�k�@RGzn���x����h޹���,b� O�E������s"�Y�*]������tJ�y!�*��P��@�v���|�F��E㬡;�W#��-ܼ�|��6�^����H�pY8��N�ַ-�rP�(�]�H�~�!or3)�x�t��T��6�dhu���e付+��{M�żsir��P:X�7(���}�J.��D�n��/i,{=�l������N�p/g��9�MW�순�{y[�zzN҆�EO���2��w�PPl<�u��G�b��uG��~t�|�o�D9�D/A(����]�p{Onr��=�}�ba\ע��*������~5�_�9��{���q��q�s���蒎H��^���	���z���X��O��.3�B����ٞ���Lv/\{���ޣ��۷s]w�nU7�<פb�c�<}�A>�s�6�i���kJ���7�o���7����zx��ML��|/��l�,a�}ۮ�n7�s�.�]���8�*��ɭ,a;㌁��H��{��m$ꛝ}�\��J�����N��l\�t������F��ʓ�O_�UƱ]1q�:����n�k�>��r�<���o�T�ڇ޷��^g����^Zg���#]rES�5z.}-%=ۧ}������U~�~�e����Tsʇp:����'�u���J�,��e�?Q�.rn{.r�kw����Q�&)����i�϶h4Z��M��t���^���17��"�����H�dn蚵��2��̀;�4y�c��tb��2�6Ǖ�����V>(u^Ҽ;5��c�S� ���f-�q��Y;oI6��[�i�d�Gr��]�G��������`��;�EZ��O��czn7)�+�4��ML
-]�ɘ5��+7�)!�� -���z�%�D��,y���ø��h,~��_��_#�7F>Fϫ�WfꪧZ�x3�v�=�:}%�8%� 0�d��{Ǚ��x���*���ʅ�aw�u�Z�����=L������9߷2$S�sp�����̢c)�{N����]F�M'��+����%>c=�,�c}N���`��z�m�_���nsf@|o�î����e�[Z�{G�_��L{}Ɋ�yU���L� �P�z��UຯA�=�%鮫�����CcB�m��l���>�|^�T&s��>n@:}�9�<�r��н��T�����]�}$���n���rP�����'|gKfwK�wp��uG����+{���Q>Qu��d/>�I������;Sg��?���g}��m�d�_�:+N����`JW�犜�Opx};��|�k�z']�zq�j�yI�����c��5KA�?Ry�����S8��׾�ݎy]�.����o�m�y�g�z������ߘ���h>[��6����J���{�k:���Q'9+轾��U�}��#��Zf�*��і��J���X�k���J/�.�(r���c�/s^�ُ�gw	�ӡ��͍���n�u�|�m�=���[5.u�N�u��Ԗ��ޥ�PD���2t�?���5Y���	F�W���E{-���<2�{T��:�]�R��K��j�����3P�g]�^L�e}�,m�����~+\_�7��:���Eyv�	׶�q9����5�./�]C�~�*�Ρ�ѓ)�\dϗ����״����9�~.�-@ڡk����KW�_���]L��⩁5<����-��ږ=q���쀧��;��������6�SR
����#[������z��mK1��S�eHfH�L�@�=�m0��+��]�hנ�v��'�({_+�ϟ���ޞ�P�~���+}7>%��%@{UHB�%z���ٮ��d��Y���eǛ8�P߲�49ש#��H�4w���~�MC_��6H	�9�y*�o�����}�;�a���D�C��x�zv��7�@dF�hy2�tz5X���}�7I <Q�>�(mD_Q�ì}�x���x�z��^,�����[@&xǪ9�<;���`O�6��Q�H�}9^q��=_\�2*5����Tr�p���G�G�3���"�l�	:U0��VE���]I������]�Zɧ*.���Y�Τ+�N���j��n�)W���3��~V9�ZY ��3��x��׼<�{a˜�boJ�b�6��I�'�.2&{`�#�M�G�z��X�V.P���:b����{U�"���Ħ��k��%��_��g�uN�~ d/ez���7>G�"r��N�}���j#\�3�ǐ��#�r��g�L�M�v��(�]3������{�z���)�צ��ڐEGz�'���OT{o�����T�[Tq�+��x�5�<��?K����w�c9�~�rz߶�H�^�Z;�O>��L;55��y1��j���}��Dr�ӣ���GS ^+v¯Vx�z`���_{�kE�mO�1��Z�}R���k9�^l�p_��ۅy>W7���o�>��΀ش�<z���^�Q>�^��Nm�j��z�¬���^��z}��eSY5��L�/\����#�p׳�ߵ[�h�{�~Y3o�k�Y����rz�͟o��9QF�ܩ-����*�s�,^L�7�>E�}Ψ:���՛���)�W���M�_�-����v�3a��|af�U3rm3,	<�_�3����V�G�GNy%����C�A汉��^�@h⇾����b���w�g�z���3 �J����׮:.���Ƶ�xG)|Uf�y�� �M�p>��#����g�VԲ� l���b�N���*�{F�ݥI��[c�;�JMc!�˨���.[| ]�$;���x'�.�׏Ѭo�۹��0��n�g��/��{�M��{[L��J���R�k�nf�Հ�����<�G�,�R�G�Z��	1n�ɲ�b쫎̜�E��]ۥ�;'�deD�l>Gٓ�.�q������"��A�1��{,IKG����[�~�/P�d��rC�9�R��#zNdF�񨶕��:���zgx�f����yV���[��Y�Y�~(�,��/����0a�C�L�S���<V���Kև���FFe��L魽�T=N�N�S>�}:��;�0��sD�P[=su�2�LM5[GY��ڼ�c�u��<��J�co&����g��t<�N���ˁ&�^�	��9�NT=��0�n�X�ͪOtw_r��|�}�}����Hh�BX�������s���>9�C�xډ�x.�i�y�y鬋�f�wֶ&�_��z<���n�+ͧ���f�ڇ�Q�_�s�>"��u1<m��=3�(֏G@��wᚺ�6lT3%z'(��e�u��d�l��X�L�`�^������tY�v����ψ�5��������Ζ�&Jҧ%��i���&��>�u��Olby⁦;�L{��i��WnA����r7�W�ʞ0��wK�Hë"��������;�z�m��̩Y��bL��Y�e�]�*)�٧�w��p� 6��]��6XW�k�hw
�9}��
W�VJ�F����	����F���j��L-�Gn�Jta�����Q��@�A-��w�a6���u��Օצ�{=To�%��S����h��u��XỶ�������3�~��ב�N��~v�g{�Q���)�E�=3�F+��6^�9e��EDƽ����T���s���^g����藖��~�H-be�l%:�񬌩C_����y'�ע��R델�-�ɖ�G<�w��^��+�u/Y=1pWT�Ժ�4�+�L�}���7�%gp>"��`=�����'-j�����q��zR>�|wO>�qsnL*B;�{4�j�WZc�~�G���l�ٳ�ْ=��p��qF�
�-��-��1*�y��S;9��̛WDch�I�_{-�8�O��0�0P{qU"I�g>.W�dl�)�yc�'&��<�N�Y�b��\��J.n=�t���q"��S���	�6`����D�>�a:��R�Wxy�K�<Ѿ�	����|==5����0VC�����D����
�4{>��o�7"=��)�3Y�Q�^L�G��[F��{�L{r����W�ޠ�ʐT{�`TC���&)k�fG�ii'��-�}W��_����蹧��V�i��/MG+�9�͛~t�s3���t�����Dc����s�u`�Ual�t���$?e��=f��y8��u��R��Da�q�����W�Y��k���dԦ.���x����ǅ>�]�-���n��m�*h{0���]��@9����=i���k���V^�P��V3�{��R}���'%�����'|f�e�35��=_r��y�ݟLnq|�����q�~���F�lz��j��7Tl�G��zO���T�~�p��'Ei�s��`Mח����T�RY�����B�F�oV� cT���mX�~۝1}��n}!��j\FW��q�5��Q)���K�+o%式x��׈�W�>^�z����	�7�RʨxMR;��V]7�z3�#;ћ���5����΀�7�o�\���3��B�{�Y�X��ՄX	}��c�N��"ʟQ�����q3�n0�f�e�az��w�������?k�r�O�ږFtLm�����h����d�^�6=u^b���&S���&|�<̆�s�i�����L����ɇ��{��NY�oH<����$�5��9���L�@Y�U0'�DW�>E��RǮ;޴=w\ �Yk˱������z���$]�w�>�K�G���f8�Dq��H�L�@���)��W[�D'�y���Ms��+ѻ��~vǐ+����F�?_�=g"W�C���nn ����!�DV�Vhu\�s쌪�"�3�J��wuǞR%G�� w��y��g���i���FZ�Z��7k�I�髺y�6��X�v}f�Ru0m��Jj��|T��j��_����?JW�g��ճclb�4cUcs�YzpUĪV.��(v���}ϱn=`�eq��S�B�o;O_�]p��RG���ԑ�~�@�~XB��h��Qd�L���l�<���GkӸ�Uy�<Jg��Xr	�̃�~�޸���_�|rx�����r:�vy41#�����u��G��g��L6��DM9�;��%�Լ.=��U�q��������i�{����x��Q�uD\)��\M�y�#�+L�g|w�2��������zGx-����`������3���N�� b�W��&��ޜ�{en�y>&�\�3���[r�p�ewRZ�zB��%F�a�y�rz���C;r��@���'���=�;�����@�W��s�+OY�wJk� �^Ψ���u9=o�v$\/i��z$�ˉ�w�o��=�۳�����]�F?T;�ڭ7_�OK lE�v�/V����:n=~���hDz���⮙��y��q�k?&x�p�Z�ꢷ[kN���j�&�V3)�f�޼�+(S�]}�X�U� ��9�S��{R;��']T��Miw3���Br���m���.|��Uqٗ���|�^�0̸�ݕL�%���,�K�ո��C��r�����Z[(�{Q�[�-�H^L�yR���yz�t$�ԏ�Ӛ��ee_[���}��T�����,1E��g��U�jzn��".��+�ͺ��c�UۆR/Ju����������y���n#��DNN�,��.2gY���.��k�/�Y�ͮ),�oEz1Rg���8��^�r�\n}�uό-�eI�T�U0&*y-��&z��{m�ǖj���򙆮יc#���d{��=����� ���v|�+�@@,��l����7;���.2���h
���>�چ�������;��ݿ:ǽ~�2mJ>�K�xwk�=�t��<o'İ7fA|��%���چ�D[J�o�^���(�>�pR���[��h{L��B�PJ��F�<�A���Ҫ�s�s>��3e�մ�&۵����OF��$1^?�V�(Ks*��ģ��/?]?;�t@��>�x���ta��;��U��J�w%���5G�:����Uu����?L�z�`+�~ۉ��Mz��KG�麇���b~�j��]k%M@���:t�{=)pKxO�^B�3��o�^7�����P=w W�|i�q5^Ed}9P������7j���%�8�wN��iZ}W^+��b�Q�~r�9���MK�%߾�u�(��a�#��h���]�A�N���N�6�L}�S֥-���V�X�+�g֎�r�2��"�*��t�ju�ua����u�{��z�W��6x�qw��Vga1�0'�
LEe�اf�����ր�F���@�Vk7���j�+D������]2�V���5���g���c�2�Ҭ9���ϭ(��k��V���*��w �Β�l(h}�:�p3%by��F8"����WcM���n�֊��T4Z��n�s�u�c����)�(K̖��C���֘)\2�{��dF>j(3���z�r�*a�w|�+:A
��:�R�^��Bm�#1�WA���RDms�H����N����[1f��h/P�KN^m��\m�� jc��[�Ar���آa�;L˷��(j�&���h�PT�ۥN�+�����y,��]���Q�q똯g-OIs&_:6*Z`L��7kYq97v�6�ks��L��ަ�l9��W�
ۧ�	�VݒS�A��q�.�)���tc�J98-)T�2�;1��$4IN��J3s�JB���Z/9Z���edt���+9H3=7�B�vݪ�T�z�X��$��E+���G���j�$��(�1r�X�уJ]7u�T��d"����`W���w{].kf[�n��-<vIV��h�Y����[�;��s�qձz��:����e�Ͷ�^M�W|w.��v��#S�Mm`��֌�쎌0�]x�̻ɇ���n�no��w5��~/S�Tnf�-ʷt��d�k,�Wj��1�����_����^����F������Ё�k�Ĝ���#�����|�兺@�S�Q������r�d��U�,�0Ō�k�P|�=����Oh*x�~����ʧ<��i�U�Y�`�ͷA�֬z\����#9��S͹A��%o��`�Yh�<�2�U��#k:@8-)�'������Ѣ�]�o�؂k��v�1tz��I�X�):�6�nщʍ���p^O����5[��!.�[c	�]�r����۸쌫���yg{�#�
 [�qm2ws+�f5z�N������jU�v�Zp�۱Ȯ�f���}(X��3%��[��]��-2�[ɹ-1���3�ko������!�2N ��tU�u�rm�>WNs�V0��_���Afy�9�6U��\�r�[l^FX5�V�uu=���ۻt��P�^��.�,U;婖r�+%]s�K:�X�4�;$�������{�+��Ƭޮ(h�@�`mLR�hshͥ�=|6��!_�y�eu�c�˛n�K�G.o;�]�پ���P��)��ǘ�2l9��Ig�o]�o7�MW��Q���:�QU8��]���S���"���
Yx�t�M��^�+��܂���9'Ʀ"��f����Y0a�Ã��07@B���o���� _MDMn��ס�}
GhR�W!->+���˸����w�5cr"����� �����ԇ���˚�wps�����r�D�q�r�N��p����Wy�s;����nW+�Q��;�t��9s��i��오�\�.j�Rk�عF*��ޕ�δB[�����r-A�D\k��Z��+��S��݂�U͢9���\��ۛ����(�ũ6*6�ޛ��W175�Ϊ�dѯ*1;���]ڽ/�zj�cTZ.�k�r�Y+��\���
��5����ד��s�r�EF�nZnƣ��*-r���\Ѯ;�w"J"��y/p���j�4�C3/7��Y���LC�i�΅�M���hژ{A+����Åb��X�W�cT��n�V�(wf�J��N�]2Wk�;J�v��;s�_�\_����ݨ��\o��f�j�E����uS�.6P�_�U�/I ���]ꔻXE��z#S>;�L�ZN�/b=8����,{�n#�~�~��|����6��ڕ���(����j*���ϻwn&����Jd�>�Cn'i��:WFO�i�r7������_k��ݨ�1��~\�W�[�X��{�����F����H�|�Oi��)g�LeDd֖0��I/xnLq�P���o��C|߶�v�2B����zpo?m����b���DI�'����_���_�/�G�.�^�莙�72��GT��ާ�|���ſY
߶��BPW��)��A�&|鍝�~�{.j�P�&c �W���L�,/��Ý{NG�W�U���^+b˱�;�Y�&�l�z�`~��J��l��X�@Ϣ����٠�M��[^������>C�m�L
����.K�kҏ��}�2}�~/~��9]T�TK����<��l��-��>ǽ�b=ܪsv����S�R�1��3���n��mz�D�n�T��{Ǚ��x�������b��9�nl(�Iaۣb�E����e���I�C�F�$��Q�6�&L�6z�}��{��[>��X�T�_M�Ŷ��"��h�2�ծ���ͻ����"LM�ݙ*1K
V�:1}��0�̔<c����dÒ�:@ֹʳ��I�C��hU�L��(�{d�;��D����(�>d@��U"a��5�	��PG�g�'a�`�O������$|3�R�����0VC���۹)�zn����d�@�c��/7[�w��>�bbb�Vѿ��{���Q�+���W㾗@y83�P��}�r�H�yM�;���ۋ$��Y32���ṲG���l��������	���h�~t�G�3���!����d]^/%
�p��;@?%���*r|6�����3k�ke�3:�+����5β9��[3|�O��u\��zʘ�Go���nNٿߤ2��������6���>���Zn5��gaX���q��X�IJ�D�@���u��W����V&��۝1ހ{D�B:va��W���\x�Mgu{�}{��ڧ�+��x��莯6���K�~D�y�q��BE��Mh�^�]�>�Hên�@�aߴ��^��]��a��^�w��� c���ڦ�{����;�|��q�&�/L���ٛ^�+�Y�6Q6,����+�����o�&n:e���~Ӿ/�mz�4��{�s�r��(
%*�|bz�R!l�+Wb�y��.7����I"�j���eͮ�D��*m��ցi'�އ2�!����=b�VY��G+���
�>׳K�K9)r��kQm&�<��٬0}|�Uз_��(	���ZK�?;jV��dV�ޠ%�<�T����Q��6=qL	����S��ɟ/N}�h;�w;�j��y82���N�6�����7�F��,��"�(��j�SȊ��ȶvK��@�u�n��V��}��>�<���pT��iP�=q�*Y�|%�@�_UH�-�.�Q�^�ꞅ���(�F����z�C>��1~�5�y�@�{/�a�j=p0Kf���ح�yå~R*Wz�ͫ�c��[� ��y�mCO)#C�ש#��H��#�G��и~�MÉ���@�f���ժ�Z!���@�ٺ�K��KGv?M+�p�_���s��~���[{Oӱ.��]���z'T�@�%n��He鹃��TD�9�;���8K�P��G��W~3�U5��ʘ�S%�UO^�z-����|�ܟB��ǽ�<���a�����}��=W+L�{>��Eq���j��ٯg�q䧖�������s����Á����O��7s�+"r��m`}���n�k��+�s{��zs8p3�^�Y,_��z���Ҽdg�ېGzVO���ُg��f�O�|�G���1T�}F�c�ݥ9��(�����G���nl]�{ũɏe׶�\���j�rSщ�,oƤ����6�3p�c��]k�FiH����$gk)�[�0P{N+l���	��.��'�{���;��^�Il/�Q�J��b����:�i�%+��ds�>"��ܕ��݊М�?EO�G��DpeR���ksSw*v=4x��gѝ�
�6�N���L?Z�`_ܽ[�2<�����s�w���_y����>�{�,�}@f���ܭ�W>W7������@��@Rs~.��og�<�Z>Vۄ�Й9���V���<t_�V��X͈ɭ/	�Ltk���#����G���6���Ϭ�&h�2S=���)��{S�юvKg>���*�s�,_�3��EO8}������.R6�����꠬%^��s�w/��K�Q��?Y�{�T�ě�������XQ}^��6W]/�l��ޕ��&c��v�,gK���p�ǲ�î^Z��o|�G�>�x��w�IVx��念�Mr�*ԯY��� �M��'�vΌ��,��ϥ��k2'r�n<��@w�x)/��{7FG�%�@�d�}��iTO|�֑��(�^���Jw#ϯ�Uk+T��=y}t=�Qq�����㈥T>F�0�ڍ��QҸ�4�^��^sJ&�YSz���غ�q'��:��t���N�www�(���,e{_���[�6�1t���K�L�@��LQ�Z�����X�(��m�촞.dEz���ޱ�K���
lcd����5
���J�<�:K+D�T��4�gs���n�>�' ÄO��GL�%����(�#n�W�*�-xO�!�:D�=�`�V�<�ÏF��w[�#M���G3���ngީ��\Lk���*	h�}7P��L/z7}QK"L
��������J�h�:7}PʎUd�ߦ�WޗC�q���2!{=6�3>G|3�3T����{q���s�z5\�^�U�kO�����EGb�lg��2���P��:h��0C���Y���w�e��/Ӕ���f�G�6�ǃ�g�ڇ���xls�>"�=���=�`:��9{��W�]��W��\�)�<o����b�Ӂ�ו\n4�,	���;�\Jۇ��gmF�V�]�2�+��2���:�c��
^�Oi��Jq;Le�֕��p�k������?/e���O3`�w��m���E��9�v����j���}�<b�{Mw�,�b��6��nke�?>����3Ϗ�J@��G�c:�$^4�̧s��{�h{9QF!-�.��L枯{J��@�����V�{q�A��Y���6�zߎDo�y��O�u���4��V��3o3�����Lj[r�Eeȹ���:!T��.k��T�s�� ؞�X�M ���]���_L=u a��Wr����+X��s�u��龁��eRq��9\����z"��r�',w�o-�2РGj�e�S`8�U^���Ir38���"�)3��ÿ��p��sʊ�U�>�^/�"����9W�E���#�Ts���/P�|�Z+= K@Jd0:�����/>٠Ѹk����^���y�M(�F���9�R#)M�/��]>�q���a[R��$6l�m�H�D�h���X�;�,(6�u��#�v��LT��<�g�cT����3��{#�6\����Ȁ�ɒ4���|����zk*����j<�(^vW��U�hS���R.s�t���w5�9�Y�|͘(=\��Sd�v��x���c�g��H	����n�>�W�w����' j#���~�3p+zܙ�)��qr����J����P�6��k�?k�n4�ǻ L<5�¼.#�U~9���L� D�^�aٛ�؜/��^����}7��JKï(�?���9��.���ev��j�î~�f�`{TR
-�k�w�u瀾>�ww��x�Pϊ�j|9������>�����ɭ,y�ٚ"K���̅��*���2TǷ�(�~���gjl�G��zr'�����z����댝�k����l��� �IqУ0���e^EN��I� ��-Vf�6�r{=����_gx^�I�[޶�m�x͂��p��ا����_50C��̓f�v��������q���Xۡ0ͮR%��37*�̬�3�Y�EF�ц�T2Yp5G�����*�'�k=�����/������j����s�;�V�q;0�ԢHY��;>´r���xz9Mi�@�wSb�[ Z^��'cθ.��;}��_��k��G|w���.��>���F��U��+j:�WY�@ǲG�(�vb���/�Z:��� �ǖ�uή�����)����h��D�=7EV+�w�;�>���X���_��o�����T�S6��ov#ޱ]����n���Ef�4]��@��0/�P�&S����/�9�qT�k��7��ܴ��
�q�wJ�h��=R��Um+�Vo��f�%Hn*��O"+�"٩b+��<��/�<�i����[\�#����Wqϟ��ng�=Y�TY������l�|�uL��U�jw�J3�y�Bë�^
�z�P���BR=��#j��V�n��ׯڎ̇�o5:�׷��nό�ET�-S������j�=��u�l�G�(�0k�WCcd�3ޖ33�kު��>�U���}��M� '�t��|_W��-�0�zJ�\�{�zv��������6�Ƌ��Y{]I~���.��]-�}�u��b֨[$M�{�T�hRg���<&C!��q{���QϜj��|F{� �N�����r`�S�w�7Z��1o7�Z��|i�����4���^7�N��R�q��c�X�8C��B�1 ����0�ћ�"�Uz������Ϧ��Z�&�����sʄ��������|j$YK<�J���xF��2}�����,
��^�-�CG���cn3�G�"�i�Q�wǽQ���f{�L��w��v%>�>ͱQ�׍�[��.N@� J�������:na��auCwT(��~9G�*���j=C$�3'������9U���v=���t9NG�46Z���	Xn}>G�"E�LKN��q�#�����K[Ɠ�@g�Xͧ��%+��g�ꏈ�u9=o�v$\/i��`l�z0���O�kiu��ǌ�蜠��,u�e�]zU�xea��}�� ��	KӞ"��W�ہ����w��>�+=c�o_Y<s��#s��\em¼�+:������#�W ���o�� �1��n4�����G��#p���o}�<m=��=[Z
ʦ6�kK����L\k���@�Gc&}k�9{Tn҆��=�{�� }T�_�΢��w_.�����T��=2�Ϯ{Ł�*rf�Ե�J���q��^Gz�;����:�=^�q.���\��]g�ߌ���y|��OGh���Q�J�>�o3d��D���3����\���\!4�h���醎��K��*6�B��>�sM��m^�<�X$P���ݚ���>�ں���4�@�2V/Cq�u`�؝�m_Vˢ�������+}=��R�>Z�G$eڊ���;���G�EK�_O����wv����z;�K����xuĺA����c�'�u^��w�ސ�x��²}K���(�PjW��چ�<�\{ ?Sg#�'�v{���gQ惻�Wx8�!o�Y�:W�%��x�tdz���d�}��7�%Q��i�a`�
`W�{3s׎��l�����g�}%�=��ۊUB���9�����������<��I.�>��ѵ��|Nq(��<]�r�T<�t@�^�l���YN{�E\2�x�{=ΗK�w�_>~�=�2���O�9�\C��M|��sD��ƦUTG[���3��M��뷖O��ǳ�}���=��ʬ�.�_����' ��<r�
^_��������DB���y0V-����a^:�:=���^*9X�7�Q�� {Q�	�ѽp��՗q��YIw�TR���{6$��˦a��ݨw�^�q��3Q�ƛ̿�T|E�Q-�u�S���}�7�����	grf;��(�z$���ó��x�{9]7�i~=&�����}��f���Z̈́�z*�j2�B��6�@
���0E��:}����gX[�o�nʊ���2`�6��!�{!�O�6N��I2�W�bE��]��yK�zO(�G��4��Le0([za�g������@���^֙�ܙ9<td�R�_D�t�_gRr[
e����3]��ӹ�̨�~W:mzA=��
���\FUhW��ZCÀ/*��qh�r[�w�\�O�����<��;�\���\M��nxůi��|E�S,]��%�ܛ����ǽ�ǵ�3�n5�뎩ی�l�q�ב��h��_����\�\C�����a\�����l�3��J���n2g�<�WB:���r5ϼw>�W�\��4[�������w<�гl"�?F�4���6��j<�w���P�r���yP�:��q^+�h(��gW���!M������m�a�Գ���N�2�[7XM�>NZ�٠�t��=�dJՓ�uoWw�L�US�}ߎ�aa�[�=�(���*@[uR=Q.�&�%�3�xl��1�=2s�w|��.>"��n�	�o�ٌ��*L�N��[�w�}^���ٳ�ْ�|g=��D�f1x��n��w��c��Zp���ca�S>�ٝ��wO���,��>��}�_z3�O.C��<k��&&����-��L9�������f��	� ��$~��菣����#�>�m�鶵k[o��jֶ�[V�����Z���յk[o�kjֶ��Z��[V����km�Jڵ����jֶ�+jֶ�[V����Z����kjֶ��[V����mZ���յk[o���Z��kV����խm��1AY&SY`��Ǖـ`P��3'� b=y��x�K�!U�Q+X��d�lP�)F�Uv�a�UQ"m��A*A�UR��)٢m��F��Ɣ@�Th�MV�I)�����:����n�Y�qQ�9;�vU�ٵ�K�wۻ6��nj����շvM͚��;\�Q�\���gm;����j���j�������s;���G]��U�֗7k�]f���6��HUƬj�;�];Z���]mt��i��vt���Mm�fL�ETIY��7v��Ֆ�kb&�%֖�˝���3Z\���b���U��7;l����.v�u���� 	��ھ�:�7V������;�S�Wqw��i���v�C�o<������\ �޷�F�����҉�C�]h+^��k��N�z�Ll�9�խ]kl| �|(u���j�n�y�u�:r
�����QE{�G�(QEs��>�(��)s�}�EQE���ｾ(�QEE�=��E�(�u}��QE4Q�џJ�Z��WU���s��r�`  o=���>�wg۷�{������.�t=S��.�N�ki{��������z[׫���3�w+]�׳�h��o;hZ�=��յuwk+��q�\����I>  ��
�(K��8��ͮ�hS]u��Yn��om�L(n]ov��Y-;��x{7�:u�m���.�������]ޞ�����hڎ����GZ�y�v�wwmŷ7wv�v��gQmn�   {��_+[Pd���]�NٶF�wg�-�ͻ�n⻭�f�5ۛ����uݻ��;��:�ŹZzV�@k=a��捆wv�p����:��궠6�ڷR�kZf�ӻ�Y�n�#�  �=�����wu��^�:s�c��z�]뜭M�w����:�V�qԦ���٭�7����-�.H�{ޡ�Ys���w���T���n�n�(�������m[/{w*�n[��wcv��ka� >  �ύU}wV�m��^)�z���W{�sӭer��{�{�((6�{�����ۏo=5��n���s�iM����^=�oa�n�Ʃkj�n��;��{[ݶGy�Tmo]���V�c��k;�l g{�v�����u��-ݦڇW��s=�@�ލ��r���q�L����;���*���H��o=zP�w{��w�[:;�����B��<GzV�\��uz�Z��w[�����˺��� w�[2�쵶����yN�6컍�i]���Z�g�t��jhivx�w��u����:�=[��=o^�r�Mv�ݻyT޲뻻i�z���hr����f�w`#���q�6�.k6�wk���֭� 6����fSNw{��޳��ˏ*���Җf�n�m�����ӵw���k[��۶�]�S�5�i��^�Խ�jmҵ���������.�޺�xS�)Gw&�U�n�;|��*��db41��$�T�@h2d0�==2eT�C�F�O��DA� S�h5*R�  �M�I!2�⟿��߱����f;���wWC$_�7�iح},��g8���R������}����>��t� (��AQ�ED��* �����Ԃ�
�����Z���&U��'�rN�����Y4:P�M��ݚ�Z�Z�����u�bV��de�agp�{1����Ҳ'V�:���n,��xY�lj�V��zHXd80݉���>�,�hl�U���Ә���Yz��- ��`e���1���mʏCe��N��D(�
�\{L�kf���(7�1��R�
�[�`[I�"��',�.-�U\�1d�1�6.�y�����q#Z1��(J:�Q���*G��;j0�e#jY����M�zR��kB�V7c��P�Ph�`S1Z�Ht�*���@Z�JK�F�F�Ӽe=�o�j`�Ȭ��B�EOK6�JՃ70���t�
��tˣ�ˣ�Jؖ��`y�h�����d9-����(o\f��ݶ�� S.�J����Y�dܬ۸%<�W�VX�~D�r;�n���oQX�)����^��\l��.���h�vv��r�6��1�-��2ŵ	VA4�ǚ�!7���G�Yf*��B�M�W[�����"T�CP��Mw��q��Z��&֭C\L[��KQ�%k��Y����9&��SK��5���n��O(m�?jHv;Fv79����l�$G��N5�5�-��Ӗhy�=YO%n]1BW�Ѹhͤ�4�K���V*\�Lx�ڼ&���kE�	�k��,6��6;,�*�$6L�v�n囧$k�Z0�a������Ʋnn[ke�EBr ������r;�I��TtN"[��#J���2L+'j�F��l-2��`ZBQ�n�CkUh�ta`:�/r�`��Xp�sp�KbúOv��+cc����o��N$:r+�5��x,s�0�S"��`E�m뎍B�ʫ��&�{ۭjhF�"Y�����,�֣z�Id�Z��W+5�M�I���p1/~��Ѡ ;�hvȲ�̦�x��P�I=9��"�)�`�H�T��TmP7�+.�[*̛��ۈ^*�HJ-e��Ok-�d�]���%��oP���/�s�d��H�KN/V5��3'����R��q�:q@n���Y�KD�:�WMQ�6VF�n
�YwL��A�p�$n�]�娞�T��l�hc�g252�ha�n��f��	�b�.̷j�٤�������K Or��T{�l	u����佬!��l���sw&]O��-ӵ�F���:��SN�G�7I���]�TǺdȴ¾ٗ�9#ImDȷ��@ۀa��@��2�����#Y��`qhJ��Y40��:�9���2"�v&��&<Gqadf4�d��Rц;��E9P�M�aN첤y�j�e��J鈥G1�����*@��:���*�z�ӗ� �fN���{���yV���B!��Ս��Z�W��he����4|qS56��c�QW��4n�Q� �V�\���[��ƵD�Of�l�5��c�Z����X��7���{�\dF�a�6�l�$�n�*�V,�l�d���)�q�y�9��G'�T�s��j��W�dn��L�Q��3vE��gV����{���f�l��-��^��-�Gv!��J���iI�S[hk���J�]dPeщ�b��i�[N�Uȶ˕��# ����1;�6�%��sJ��w��� �f�(^4��T�K�01 E0�ån4��([y��uj�&e�J��)m���:�Z�Wi��M��`4m�o34͕E��>���(��OR�׭+�0S�Gki�փV��{a���G2[0�t���F�V�GI��ג�HUWD
�in���ǗCQy�m0��$8(Wv���ٳ0��Y�^}�Z�����5a�-AS��� ��*��������:�q���T"%��-,�(�М0k��"���Ųc/I���tT�M��L�d;"����cFf��Y���0�w*H�R"H*�`��LZ�e�E7I�&�*�.��ը��;�1^�NI�K%-��u-���8# #`5��~��Q%���<Mq�>'�qobO�9e����3m��Q��ΕJ��o��J�2����Y��V�^a1��IN�!@�˭���d5$�͙e�EB���aG/u��Y�c�h�ˇJ�h��lgƯ�\�C*CqMғԝ�&S׵{`�#K�����,ͻ�Ǳ�ߎ��v��v�ï\L7�:�Œ��i�x �Hek��eZOV��H�j�ܺP�3Q�lV)�	ڥC"�`�lĀ�0V�l)��CF`!��*_V��]z��׿X�[v�U�*�"e,,�%�kqK�J"9j��|�Ffa?f�2yy��5%�+
�i����f��n$�O�&֪��v�-��VuYTdY�AhR�;��B����7�����Q�	U�E�F$�7��^Ӹ�������#+3w$t�6�Qj�S�U���*�M��d��z�H��5ukR�%];p�Haez�V8Ĩ�/L�/bQ+nۄݧ����1��4#W@�+��r����$�[���Cd8�mQ���*Y;nlOE�X+��z�	�A����V[�(�r�Cl�I�.2"�vR��HG���LU�@�h�B�r��LJ)���⫺��L	(Ix�7�4dHcy�8-�v�3���0�1��[Xf|^(k	j�k���ȶ �-`��D��ڰFQ�%(�.�W�eD���]Z��.��%F��bAY�p�ո��d]����i$�@���w4�̭-	�xN� \:���*��lr��z�aM��Y�����m$����	�c�7��cr�)��ב'��2�	B�J	�4I�5s^�˽��k[N�l�冰	Y�w.7�V��m�+������6V$�Вsl�tM,�n�2&@ʺE�4��u�&ZgdL'M�!��0���[�V4��~x�Z'(n^͑�����q�hЦ	V�Pz�(U7P�ZXj���X���En�Y��ǒ�����n�)�C{V����.��<��V&r���-�7f]*�'I(@��L^�\�$��S6��M�f��R�wm,j�j+g�1�8��_m���d�*T�I��n�yk4�F�nd�y�h��q9>F¢k�B^��`+�֛�$�bL�e�9!�fT.��M��&I8�
i��f5���#2���A���޳���aOv��w{�l�L�������F����^���D�Xt�ɪd���m�ͷ�ε3j����F�ӆ��u&�@c˒�����v�-+MKF��^pO]]<�"���kb9{��r�ȳ'5�{q�JX5p)YoI1�+v�^�Nc�˥y0S+Xի^��75��#/�nS��n�\iB�+�.�N-��7��ou�f��Y�f���"ٗ/mۀK%�"b���+�i�违P�.^R�{�f=�ԏbPZ�9�A*,��K�X~�[㻋(�Iä-%�W*Dn*͡������ۓ+
L�X�z1@jJ��<��M��2���j��/��hCZ���8qq^�����1�-[���Mt�)���N��m @���Z{ J抒<��+hQ+u�J�+bC
�Jrl��c�-�QXm+�Ąm�)L	��+0�T��4c�X�W6&tfT�D+���hV�h�)�(ޠ��lշ�贉&;��Ujkr�}��ۉ�gb�Yl|�*;q�$X�.����U��S4��#���E�͢�˶%�5�WK0C�A��ee�2�1�R��D�)eBV��]F��v>��9Q��Xˀ�5�{g-�$͇a������Ӎ&��׌n�#�$���h4�T�m��4���(JY�S�j�i�/6���bi�W��
 �4�)�nUŘ^6�Hf��r��]�.}4K���(53U��a��*i6�i�&jKn�����PE��+Z�E���]1A��+2n���sh�˱m��M�y&ɆVk9c��*�E�j��d9`�@[TgQO
W�m�	Y��+Y�9&V�7
*�\Ke�\�%�qV�"",9���3<K6S4V�$),Mfҷ��&5lݚ��e�РU>�m�Ҿ�J�qyҴ�D���]���#T��N��J2��n]�q���31k1R�m�v��7-��E%�R���n��υh�V.B��z�9	B�1�)K�v���mF� "&�v���b��m��CPR:��d�\��b��{LTP0����a3f���dn�.�e:+Mi�w�0���/3C�(��h��+0Ы��i�� Fݚҙ��aAp��Z�g@��ȅ��F��:�|�&�M:�B=6R�a+9v�3V��8���=R򠚙+n�4#�{$4�-�ɰ��Qܳq�Ű�Ղ���5m6���mM�I�lm
�%YWv�^��h�V݂��dؐ$�bͣf����L��"���:N�x�˷�^b� uz��:�BhX�k�[�]�U��jL7�jrX���j/^:T~.�IWcF1Y���z���-�^�&1�	O;�;�����v����x[�Z�!K�ljU{E��*�I�.�,;gn�S��K�14�<��� �@��la�5�;ym\;�b�I]��l�q�}�G�B���]3��`��>4�b�j�Y���32e����h�+.��#��A*�X�;1^K � �@[-+�,ݫ�Ӎ��!�����Yr`�2\��7z]{ſl�^dn5���	�S�f-!-ͤtF-����dP:�U�B�`�NM����^C�i{���MeaH�b$���G3 GsG����0׎��RUN�1�)��I���QA,�, �YR;��!���X�{�rˆINm���d7[{���U��eK͙�v�|	ǎwH�Ê��E&�~�+'��L�L�Xn�f�� �EZ�oX��r݃���H����͎��9��Kz�ZFF(���']�8-5�p�R����JZ��X���m���sX�p Q�jT�D�h+�jh:	:5��N9	!����>ʘ��&č��,f	g�6�?H�wx�n;��S4�l�M�φ�Ӹ!C����47`7�Qn\x���F.=��"Ū�q�]�����!!�z�"��,&f��Swp��@@I�9��BAY��#M��l�L㚍�� �{�9\���l���%���d�<��f�n����D��ق��ਂf��j����İ��JݪCYP���F�#7� V�����MJګ�r�������wۦh���9f��X�zv�p�[ ϔ�������2����Z��DD�¡�q�3�w!<�{ٝ�ﮠ2�]^�4�)�v�Y9�YGs^F���`Z,*yi)���5�z,nZ��f�d�Z��i�
7k0	���G>����m5��N��7��S��ȃq�� ll��Z���i�y��V�&/4|b�ç�{;! �f���N䙥�,R�l[�K�T��������Ahߛ���bֆ�Mʐ�����;5D�Y�F޺�7�,�Sn�[����sX�N�R��m�g2ۈt�cGB�`_�z���1St���Cc
�@�W��o
8�4n��aH˻a+�Qi��&���+��	�5�������TM��R��0iyje�d�*Q*��.LG2	#͆U�{�t�x�qav���ۡ)���6rM�K)3���`R����+L�wBk_��E�	K`���f؋F�l��TU㽫��h]2j7�0ڕ�(��5���k��L">�q�[�)����홂bJ3+2k�ѯs�y�qf��7h2P6��Nf^�[�S��k�U�sX���3�7@�*�V�Sp�Oe�[����֤�N�ю3����-���ʄ��0�\�I$5b��+V�ͬ���e�:��G�Ī�AR��0z3hA��!�Ւ�ySm�W��Н���1�Ol�n1�nQ9x��2)/X���E?��,ȅ㭩�� MH��������D��Z�ӗI���vA�ށ�h$<�Ն �-"sX0vk0-Cu�-��p����e����û�	��2Nm�9����q��I���y��J�5�+ge��jf��(�8�-Q$%7M޷W�&�CC�� �B`ʓc:���b�k^��
��N��{�d�ŧ2]#PTf�TqI��j��t��Hm�9[��������lD�mĝ�ix2�Mқ+�"�{!��Z��{.�.h�Q�B׹����6܉��>�R���0�j�	�n�	{����c���n�x�&�ۀn�A��q͖�Zl))�f�YY�`��^�7IL�{�^X,ڡ������e�n�Y
6�m 5%�;1K*݅���A5ՓMA,S$�C �ߋ�9�%9�c������M;0�aҸݑ�(��]��R;��k�I�l�1ƪ�{�h�
�n�k�Ne�j��j9�t�%]�p�]�+��ƴ�"b��37�#c �3Z�G2�]H�9
��t���xP��+�q��!��DFӼ7��w���NH]+�&�թ�$1�r�孴��Tl�5�
:�ңN��4�4�4SWsnA�֠+!;�a�2�1�F�Ɣ,,�:6=�G
)��{��Mћ��xsz�U�n�#)��I�%�H�afm̖1���`�7�m�X�U�a)i��p2˕w2�#���֕P�uV�c��%�5]ic�O((4��&Sp�H� ����a��([:�"�0��<c>����#8��D��y����^�&H�MYyk�BU��D�I�09��lq��)��5�0f���\�z�b�6�&�d��=Os�r����8t��Q<�<�Z�8-m�����޵���sj�ew;u��I�e7y��2f���1���3��q%��t�l�m^�
S��g��(M(�6�����y�u��g �j ���=tHt�\����u��n�^��YǞׇ��!�%1^�g��Ll�]�=��iSe��Y[Zn��;��%���|2=���W:���P�*�vSW�!z���V,�����zd�����{䯅�u��޺xҪj��Q2ZVYep�d�p��E�<lr&F'M	���m�el��qǄw[�u��t��p���1�v��e-�@��V�!6�m�N�˲Ƃw��|�f�V��X���Nc���y�{�:��Xb��M���Q}����䮭u�d�4�P��=�Y�v���������G�œpw_#�@�ѡCU��71NFy���M^�if�u9ڍ��S55�T���,��ulZop�lJ$' ˡ��z�C[[�i&u���}��}�B���n������p'˞%��I�r4s���]hY-�c�PtԷf�]��Ȗ�'R�����y�θu�є�Z�Q��6T��w��ᙍo�6D�\1>����<��Y����v�q�/���m>�s/a��z*���a� W)
n�w�jk�2j�9`��ff�k�(%ּ��o��m��'6A�z_�9,v��˱{z;���4pwh�x7S���`��͹L��E��'�U�85h3#=�:#
Dmp�l�] �\���.< �2�������b�յ�MN�&c�/��R�u�u콐�T���������B'�����o���؋>����L�<��ك� ���l�4�(��� ��%�T����џ+Ru$C8���fAC�/NR�J����*�YR?K�z=���+�.j5RU]{��+ƨ�BtI�M���]��Kl;L=�6�lP۟v��FP4���OʸjfL��3��q��3�i�cv��4}����o� ��!�FM�f�ܘix�^r�9q��V{�0�+����l�������p��{�dQ������FU���-ko�����+n�Ǚ�l���/]���7;��xo��TY�IQr���&�?7����ˎ
��v���!���)]=�����d8��H��aۆ,=J�棬���o��'�\���]��8Չ1��y�3�n�k������;���8`}3���c&�����ӑ�J�Ӌ�Q�G��%�՜X�I����!?��e_n���
@Lg� �p�r� �^��[�{vbv����P�R�Ur���b8�@!b��+9��𼷗PL&Pa�|x�D�߱��M�K�f�VŅ�������= ��'���/+q��f;w
᪲V�˯9j;`��t�W�A�vʸ�*ظ�[\�b}�ׄ�Q����]R����͆���ؤw/BA����Q���ys� �rY��iѠ�ņ$H��l/0��E�!Λ�|�ۘ�Ⱥ��ܳ��.v�Fos���Yc��n��v&=.�|t=#�<�*�.��y����[Z)�:ӇY(ؖjj����mps7#z�@�㕳Z���o+�HaA+��ٟ��lf�K�k6�W2w2M|����6w��#!5z��N��.P�"�k^�����9J�qy0�{�/�U�t�p������Z� H=6=T�&���u0��U�����\�V�*���iK���P��9N����4a������s��ĺ�cu� g�|a�r+��ŀ���x��P�0�ԇ�m�`�+}�.��}�;��7)}����k�y���%�`�i+��n���D��<�����e�F��4���.:}���{�a�C�kNL��$�ة�?(e����y��C^���'Rw���#܁V�cQ�� OD�XL|���(fn�ћ�p���R��9��XNQ��͕�.^���ە�ۉK�(����
8��0�;o<�Eܤ
6��`�Gis,�Ý�<m�d�ȶZF��y�fa�'��"m�ّA4�^H�/�m����V�عx]�f��՛�x�[�m���7�򋕑q�4G��]0HQX�����-�Եi�u���H�)��W��<�@�ڴF���F����r�}T�Fv��.�{��C��gZ��bX��9��%�۫��X��;r�~e\��p���yGuH��柫�bE8�v:�0�ۦ����/Df��X<�ҏI��X�ʝ�Kqfn(;�9N���Y>3o��{m�� �}ɋ����QJ�r�b�2�FI�p���j�4��3'��;�����&���
�U���:]�q�
���/P��>]ww#ۂ��o9>_k�ak7&]�������i���Wۛ:c�!���S���`ݾ�_@����wJ!��Zc ��C��5&gg���*nz4�h�br��q�೯�X���L����?b��C�E��[�ٸ�f�b���B�H�xvva�*�x汒���Cq��u����+����3Ľ�W\�۵W�zݗ&�-�\�κ���v��AC4�R&]LJ�˱�N�/o��z$�Xp�׸�Z�ZA�H��7����̛{���W	�{@F��Y�<�R��.
қ�G:�ͥ������u��r;�">.3��ug�7��LM�dpkU{7m�����G��s�2S�g7��ד�����n��fVC��.�יz��EG������R#�[�Π�o���)s�R������_3����`�j���9*KѠ�mL�іA���)�rN��řG��^ۯ#6����K��=K$켳��f[�<�FuK6\� e	��B�)�)�Y�ˬX��.��i*���#J��Ӵv̨���[[,DZ���ϼ=��k�T�����Z�;��s������a[�wur�ܺ�+�l��Sw%K��DB$���o�^�V-��[N��������b�Mv�9��)]gk9R8lr��y��n=Zږ���<���i7q�d2؅��jc�>ͳ�	�{+��ͱ�7	yN`���N�čڈ<R����5���
-���̄#o�]c��>0�ٛ\���^�0��A���Haث��~�ԡV�LÝ�N��E��>S{Z4��r��U�!j��]�)�b�ۼ�}V�Y�ccc��,�S�-p �Η*N�^<�f��v�I�^l��(�ѽ`�\P�����\"ѥS�
�uT
K��Wł�J�9ë����<������3Fz{�ƘY���R&��/���$!BW�X�÷�.���Q�F�L�u�����V�Ǚ0�(r�.z�x�Bۉg�O�7t����j��4�M����u�OQ�g��h�MツI�F��7ڭ��64��(�*��7��^͚�/d�ځ�A��ȅ��o\��Y��cg>�'
|*�4ny�ۃn��](�fG�T��p���-y޽�����>��xGI�V��i<�r���3�����p��q�n\���b�M������D��g��zM�t��_'ᜬ�r�eHn�:{�F_)-qa�w�c�N�63��2�_Do&�뽶3D���F1�	�@Gq����b��������ˏZ�3EmJ�SKy��|��Q��_>.�jՖkok`R�!�i곋:�4(�q5��J-�ջgE��Έ�J9y���]���5Io��ɺg�p��֌��.r5/#.2wP��v9��>�;froX�ó	5P�y-Ϸ7��<(��Տ
k�%@(�� 㳥ѼH8�Z�.�}�\�]�f^�|;`۝��4qf�Z�q��Z1 ��>��;r�v�^%;�ם���xt��ɐU��0mmM6��i�1�m�sh���6��Ųr[C���=�Ϝ�a[�6�\���6�ک��Uv�0���
m֘�h���o����u�PhJ��%�j�CӬ!�Q�6�[s#ɔ��}7k���{��3��HD��r��xۨ=
��i0�E�z��uJs:\��Z$76e��&P�����ڤ��e.3{9�e�����T#z���L`���)ӓ��K{\���pHt��`ɖ�V�%��|�1�2P�����͐������]yc�jv󢸤�l5���w���9	������sy�L��
���^+
��i��Fv�Q�W���[HoN�3$]��@�6�m��[��!�r	8��8F�Zn���%"�&?��A2��p^�";ܶ��3�-K�`k�����e�(�ǹہ󻮱�N���`X�D[�'4�ST�,Ѓ�	�W,yiӫY\m��:4u�x��Җ��l���b�	f��,�9i=�,��#ŧ�����Y&�7@�����0 n�w.��m�BM��c֏������꘳Ot7�etyM�g�Ɵq�o{(y*{���I�i7��/v_��4:�S�9J�M��f���A�)�gD�V�|]V"�ff[K��S��Yi�9F����@�>YO��y8xb�ZF����]b�D��D9o7���pæ�$�-�4�u��;��Ջ�
�80�qî�!�©���R�K�t�}�%�^�h��OF�+;f�4 U�	�tE���
,�h�azs�-�:N����̣�}nF�아E>�����w�3厷�.5p��c����ğlg,��y"�Ƭ�&0��&/�0;P�7l�_'��~��+ywf`=ڗo�g��{\*���, �,�Sj,���5�4�4��1�;m:��l���{{g",����"N :}�"�ݹ��[��yj����Q)��=��{_�o=�Zg1�cO f�n�2�q
�ZD>go�����+˴�}|n�7��N\�rp<�vU�Z�����ϙ!l-`��K��J#S�+*��1qhL�0��C۔u�ۍM��{�2�K*�^�c�7w�dP[�ef�v!���w3�3
�0j�YZ��"�_��+G� ϕ�)MQ��-��rې�f�N�q�4��0��uwu�n���K�i�$��,�@���
އD�w}��
{�(mp��.t�b#R��]��Qk�<I�>��C�����\���(�#m����\ce�%����uua�:H��6�b7	�2r��yT�N(n�C7b�v�{�G�[�|��q����
l�����'@�r������Y�$�r����Td�b<���hF�Đ���Z��P�|�B<ʖ���hV˳�gp�:͈�v3
<u��ǌa�ݱ0Y��겿.��
^�?`�{C���;���铤�ka�� P��k���ğS;sT̲����>��v�!{�9`a|a���Ә<�<o���m�S�W�nW\�L��&x���}�'ER��<��ܢ��=;�MT��E��r�#狖
�,8�d�x{�_x��k�ךJ� ��.s*��sZ��_c�ŖtGf�Лu�#6W&�>�Wx�T��89@-ч*˺�7�ݵ��A�G�V�ͱ�`x,����ݔ���ᛸ7#��2�f����b�Z�e�W+�rtIG�{zqD��|�R���47t�l���cZ|v�,�$���K�ʕw�k��ʼi�r�<(N9K�g&�#a
;��.��Y����%6��z�w�"�ᙎ�X1�8��Txg+2��R��K�dV=�a���լ�K͡x-Y����J(9�:�$_;P0�8ݷk�C
&�x���z��*��w�Zۉ����Ih�{�#__�P>�-�Ǌ�E��d�8���#��>��ɬVr���]��T]�+��M���C6S:�+=vء��ڨ��|>�gx�IS>��w��ȡV0�����"�>�{�
%u�ظ�1s��7j�{�)>��v����X��X���5�1{В��+�8d�e�.� �������D���T�s2��$>�\��8w��X��"~�%��+�B2N.�B��NH:��Џ����\k�<2��X����]��\ל\n�6�7i�;��wM!�v�W=<�Pv�ǻ|u1a�e�PJޗ��>�N�;s9ЅU�Pu��8��7g�������>_Z��7��fWk����zq��B��<�}�Z��>d
���c�ח��"F���y�R��2�&9�X��8]���e�\.������'��A�����i|����_��w��f���༷2\��h�cM[�-���/�r�/��@�2	�mr��ƞs�]a|�r'.�#�)�iV�(���w,�w\��9e���U�y�;e��e�9�ͻ*0�Q��^�w��{�"�z͂�T�+��|�%�:-l��;�q�e�wH.� �W1�i�b'8�Gr� �"}�j����˓!k�>����l]��\E_Q�9,�UM�W�V؃��t1��h�Y32x��WL\���i�F��Ŏ�9ʧ}̟y�B��T�\�*.�η<.tK�,mM��+��E.(�*Ul��0��5��g8�6�����!��2�!bshuVg=�5.�Kv��H�@\� ���eQ�W���jk��F;��Չ:���֡��C	����映������PH�v����u�2���k����7�Z>�c��t�@���Lh�hc��ʅ��.\)�]���퓻N`�F��JZ�f�eB�U��2�p�&^v��9=��R1C�0�h�+���C1�VPC�����A�n�k zlL��S���q�/�Gc0Ŏ��
eb��d��5}�|/I^I��bu��N����B��8&eo6C�L���Q�Qܭ��T�5/��l��?���Ȃ�� ���Њ�+���k�������l,3ԏ;� r'��ӵ9�f��V0��jȉfӏ��fvAV+k�67H����c_PQQ9��x�Uxd�T5n�a�K��x�~2ʗ����;�.�Q��S[���t��������v�����F*p���	OT!ug��q4&a}euq�ܺg8FϘ۷��|�Dٷ)�w�#�m�En���d�P���N�e/��yeea�8e�0��+E���m1PӐ[��Q����񝥧�K���*98x�|:����)�7	;���L�U5������Qrq�;��K�;�|0h�f�9Q�Q�:�Vˠ�*��l����c��B�gqD�� nN�b�i�b9�s��Yt�e�h�;��樕k� �5V2���]�Ӛ�t2Ƒ|La����2)�1��n���'c@p�r/)_1�%�;�΀����U����<�5*O�q���l��ڳ�U�iM����u�_q��k �m�ͅ�f)b����nSU},�U����H�Ȭ�g��(��W[1�8��@�z�qYw�:�����|����.����9g{���r6M�����4��Oɜu$7;kˎ�����T���K� ��J
��,k�KM8;M�b�>Ƶc=w/��')֫L}�����$�zĕ8� �lJ"��E��ܧ8]��{`%��׆8U�k��3΂U0��Kƛ�\��gg
�ݜ:��5iu�W�R6����M�\�D�8�i독R�(ɏk��t�����Z��7j� �В�BJ�L�R,Ӄ�Z��2�e�t#Xqs�y�e�쮸��F>�9v��ec�I*��ɻQb�5v�BʣT\c��� y����4gr,:ǒ�|�M��<�������C��m��R'wLk�{9p�ϔ���(��v1�7l�q��8�s��j�
1�=V��u��R�˫'E�6K�n/��8�j�yr�=nCB���;�3�1G��b�{"�����/Ͼ��t���ט��h�H9:������Ta���^�j3��!��zi�fkd4�e����X�nV^�ކw+��_�v��$*�m�<��B}ǽ�m���~Xz�d��u�>T�&@xA�ύ����Y��Q����LDWG���Txq:��7F�s�L�wE��-n��شav��eqh6���x�S�+�m�����aV���ED�*d�\6N岐��ht�1�6���;��"��->u��#zD���;V^���7��j��1G�����G���ڼy&Z��W���,��L�I�9�?�����hۜ����x���·;ވ)̛���ط.�ol�ܙQ��l'�Y��4�%0k�|�|aM`R\�$B�+�^KP���$�N�ڵ���\J�9EJ!k=��K�O�-R%�`>B�_��o�AF5�u&�7���e���%��1�`�(F1L�K��-bHnn$:3/�(ƪ��rf͵�-�,-��-�n���F�"��~������s�9��'>+�^�i�y(^��*��|��7P��_C���f���V�s��9+.�z��x�ޗgi.�s9"MZ��YOiG(��ue���%�}�!�;�r�R�Ըa��l�c4�k�m�i얥�v�s�Kx�K��}4٢q�ĳ���ԃ��Ý|�`��_rtR�\����k�iٜ�^�v��v`�@^�X��*�5��cy�G8����ՠ�{�<S�:'6�j�󈽮�b�b���Ԧ��=��Ky0�]�.��4x��!��j3�'v����5�*�B��w�_� �|4�-��(�RU���F� �ȴ-N��ϫ*x�a�֞�l��X� a��}g�.��;;��sv�m��{xb`��rd����:�H	��]�e��s�n�(����#��Keb7��N�\am ^	/��ܾO\s��벶�s,�E[@�/Dy"�z/��A�,m�3�/e�Ͱ�]ӫ�G�o�*�0�v���x��q���]0ɓ����	���."Eź�mo*[t�Pk3pRt���o���l8.��	}�<A#�� *9Le�<�e	��V���ww
�18^3��ϙh�#�X�[��e���=5�����˛O�"�c���8o���z��Y�ӆ@�6�Na��^�Y�*�#ta(��29��iW�(]�ض�=��[�}wAP��f^c�ecjÈ^��ٍ�bl7������;���B����iO�S�Ӆ�*���{�;0��.#ؑ.�t4}��Û�b�ޛ{)�+J䥡������繇�;�{��d1�����r�3K�[�9��2�{�_Y�*�of);aݔȘ(�F�.=s������+��i�7��wU����2��`��ty�LLłf��4��;�Žj�:L��&l��+1;!d���k�F�	�v�ntn�%D ���V՚.�8�{D)U��l಄��K�ǂ� ����<n����l���Kcu=ӯ�T��l����ɢ���6tG���W�m��e���i����}	�)��lc&wT�.��7�9���.�f<v���j�ˣ�J�&�.�޼��KNM]�^��vg������[���>+n+�[4_Sk!B� �����v����Lc����K4�$����$�7'�ͧSsJ{�<Q����_h}7lɢ�޾��f$㙭�c�c�Y������s��M��@'c�Ǚ{BU����	��s��*ǣ��S��G:�|m�7ʓ�m�����Cc4��4G�Tsv.�u1����n.��Ԡ�P�8��1�ϡ���Ʌ�Xu�����]�պ���5�]�b���t�6}��Tq�^�ӵWÖ�l�����f$N$���;�����^EՕ�	�Ȣt���	�T'��Ƿ�W1��Bu�7�������24�\�q�1#�WI�{#ys�&�WdN�(��D|�ӊ�۾,?7��d�Րġ���YYN�<��,�vwp�)kS�ٛ�y��M�,�Ax��&�$땯��kbq�*fKѰn�t�2rf����Y$�G3��p.NM��t���]�Ա��sL�uh��-8���M��w0�6r��������Ww���qw���*W<3g������o�C]�D���^EBm�h�rɛ�����bZh]���]q|�d.u�<[ߒ�yj*՛�v�-��zkN�~I&��\�H��{�NS.8Ε�+7L���顶u��T�#��}t�P8���j.K��&������f�H3<�w7�<qR��	g*��;�g{�$��n:,L��ﭏCl��0^�=��������Q�2�R�sLs<|�{\�K/(�n���E5�r��6݇\�vKN�Q� E����z�kS�����3{oK�w��{����εȭ6�9�̊��:7������[}ǘ,�Mvm0�G���ø�K�<^�)�M�ha8
9v۸ۑ�{A�z�j㝻�+���P[�7�v�"�ſ8����l�3�gK�f'�������y�;���C�nݭ�4�&�$X��5���eN��7GE��qb���"�sB߸�VSJ���ӂ�+�"���I�l��Y������-��;̍�R��'$j��I��]t�^osB3���]	si�J��D��@ã$�7'���Ľܝ��YN��W[�ؕ�8����hv'��Gi8v��֟,,	��d�)��jI�*�O�%�i[;��.!�j�׹�P�W�V̵�q��}M��c���hf5K$�VVV��K��m�tb�ø(豵��6CJ�@�5
;�Rǳ%┷�)�ǎ=#P5��94Q(�J-L�P�"�h��w(��6��bE�.��A�����I�U+�o���rcY`�d�T{�����BS՛�os9�X�	�rV�%�04�c�۸��k�.��#�����wX�V;��9xK%�;gJ5-+��������+9O��ۨ�}�H����Nم�� �IUf��z�D��|6�S�at�֋���˖�[�-������2P���ODq�E����j�P����fU�w%�1���AӆNd���f�ڭ��E�7g[�{�V-��扖Q$��.���ؒ���c�0�N��������0�x�0��E�E�w`���R�|klK��a��Sɡ�.��f����&�a��ѽ�n0]��i�#j�e?�B�WW��mRT�;b��V�6;{6���tb\I�-m�[�P�����)wsc-�t\�34ң;���S{�(��,W�ݴ6d��*��nl�7�gl��*���N�$'-��֛:$���Yȳh;hm���P�L�,0paq����w�qPz�7U?It�������yǯ�UVB���W	s�*�O�R��XwFs,xfkǍ|�<O����.g�:�-�����u荾��l��$Cs]}����l4-�D�S�V����d���:F��;�X.��ڱt�
KZ<����Gp�'m���Ť$��yGd�^��Qg��ž��������y��y H�S@�h_t��O��g��87�-�Q5�f|�\47%M��;�
����L<�4�»,=8c�V"�މѬ`�zx�1��Q�-ȸ�bU��;z�WՉd��H�h���:3`�)M���.7�ٔ��o:��kb�8W����wMy���َ;xƫ��mc�x;Z!�`�(Ȧ}�Xx6��w��B��<kFm�czsl�2�ՙ����.{.su]��vӳd[2�<׳	�#������V��7�{AFʍ��{cӢKVz�$}xbcVbLU���(�[3�嫈��Q�I�n����e^i*��Ctv;^���"9�Աa����[p���sZ����fh�����|��N���hO��-QӔor��Sc
����B|���ͺE����
L�l�(�<�$�zK�q;��]�dy&1kd��]	۸��pd���w1]�F����{��78\J)�PD-Κ�je�'BN���d!�ޮH���.,���*&&�D�m9�����D5�s����](`s�=�D�rw�]Y�2't5��Oe�5y��L���/3���e.��
g+��K��7���|��*u/����#쐊q��B�Up��j��A�dy��+Z:�x����;E�<`����h��BV�G�͇�;.-"�fJ=�[!�CW8fmN�b9ֵ10vq[f�؜��nP�;���ҵT�n����$��l���W���XI9���O���2��/���^�*K����<��qo��s���z��1�s�1#��U	Y��l��Lِ��v-�Sj*��7#��향^�6�fP-�Zh覽��T=;`���(�,;x�@��(;U��rXvwu�%�/f�L�'�ˁ�&�ή�4�F�Ǒҍ6 ��"Uۗ;�j�8޹*�\[o$��]!��a�ܺ��KS����C��>O�7��L0R�e����M &f���+Φ��k�&�t=������fEp���y�$ٻ�Oh'v�p�KJ�)�Wƴ�E[�l�j�ͥl;jعe*�L#��1�L�&�Ն�u�Q���d[[.�����%n���!��o�F����vV�È��)��F��ZVR�1X�d�5��Q"������d:G/�7�i�OSSw~�U ��wLT�t��By���(�%Ey���ް�)S�ڑw�Pf��T4����s����º�W�p��an˜��sW۰�)b.�b�yN)fģ�S9�a���zm��f�}���V�^l���^�dd�7�V��w�66=n!�|)W�p:Ë����g]
s��ۋ�Ô�h�}�x��C�g5==QS��L��W��){t�J�nN��+��o�`F'm-��i�7/ "��Se�2��f�Mo�j�#��w6A�Xٙ�	�0|~�'�Y���6LC �T�/t�o�f:�`�F�ᇻn����ŪE��Zl+��-�r�Ԅ8*��,9���%�:ʍ`�+M�y��)���3�rݑ���ښ$��@T�xh!�1L2]��}�;��'r����!����\�`Sg�*iٽK�Cb���"2������R���MV�b���aޝq����״�0��̼�\W=kMH�K��Y8��F9�4��י]V��4�yU��%�0�om�}]�cR/]]fpfH�IS8rr\{�=��)m�'��[��%�,�%\ah1vJ*l�;���V�.oa�� ;�!�>��HHr�����z4�4��4]�$W�r�ض�.�%�o^-Cnp���C�J��t�����x n�e�Ҥ6ֵ5��be�B<���Z'8�Q�4T�Ó����_���ձ9�������3��;u��%d���NJi�n����J�uAK�X��mU�b�����NG&�$�o��r N��޾�N���CwΚ t�]�MJ�X����%}xu���b��
y �A�ݨ�F�a���u&rkچ.K���4]�h�s����s��Y��;���� �aM9.ĵZ��n���B�L/� ^K�0}a����n�5�����Y7�
�^-]��L���3P��w�ݥC�xw.3L�ij�L��X�R�����Cq���1%�Nm7fi|����z{�0pr5=�p�\�Ld�A3j��$�+y7�ܽ7{�9v-�z=3�"�*蝼�T���KKD*�g2c�4�*[}{i �lY0̀��]�G1��;\�2$��"z����Gw��������ާʆ�%(�%��޳GP�����7+�yx'X��hв	0Z�ٕB��Z\������/9�����A<�A���\F�2c�XbGB�zs-.����T�r-�̲/�.��k�W�L6X���׾�x�~���d.-�Q��$������}Ǝ����4����2v�	�9n��(�s|o=���c,���`�'n�=���ݚ�}�v�
��)��y^��ݱBO�hj��
a�#i��j�r������Ѫ]�f��j9��0X����+9�����c�9��n k���m]�j���q��DV4�>&�#3<�Ǫ��,$��l\���wH�������Y�a�yNB�Ē��3����+�u�]=�8I;��aݗOS���ڰ�	̃cH��?r��ipy��Hò��1+�[�`5�=�
����9�1[(�a�]��҂��q9�zOC+ـz�c�=��@����*q�s"��g*�$V�Ib��e�VU���v��Wu]p(w
�t��%�������{l���>n�1X6��sA"R}ا���[MH6�"��n�\��ӧuy�9y�V��U��"�7C�yy�ic�-j&��Uٶ��v\��i�l��a��"� ��kf,��%l^D�{F����g*�L�:e�\�֛�>��_�c}4`+������]fѧ�.u9���Ci���RCÆ\��t��w�8��ˇ�������/��E��Umy�W-ݤ,�}��u������ ԍ)K�	��JP�e@�@�#C@&J9�H䩒!Y
P�BP��J�&@Y��H�d�KIH�%�*���d�9 eB4Td(d��Hdf`�
.HS��&J�	NJ��B�%���+FB4��VH&C��"d�dوP9	�	NA�Dd� ULIEP�	B�4}��;:��_{���,�s� ����Fx�9w|�a<�n�{&�E�2�i~eEkwٵR&i[�4���}J�|��R��#���t͵�JB����P���.�$���|��YMJ��=|�=�VQ�e��ΛT-Uzo=)�7�#�B�1�(1S�$k'*m�F�lP���<����d�:Cq(��f�7q֯��C��7�C`Zx+EBCi�`_2��->ݓ� �ֻ2���;R�9�.��Ȩm�B��V+8�W��{}gV�|�Z�ݩ��E��S�U!ʸSG'�2�*�pr<��<���Y�da��9�"uY�ʉ(�d�����B���
5�������*{F���>�N�#�	<����mQ�����N��[�w�	㎵�j�qz�z�ti>�\�2�5�-����s������#��>^�@�o���K�­α�D���Ic�\���u�%�[�zr��A�m�efw��I�3���5�X�?{]E���ԁT���=�֯���=�9��CKj�	�nwR�8�xH9�a��OA�w%3T�q�P[��Lv��\���dƧ����9����P�i��y�ƛȔS,͛���x4ۡV��B�J�A��p�^�NX��&��ǎ�ȍ�]@ZL̠�Nr�������r�����~j��SQ��j:���h)�7dn�Gy8�sՓy��g�{���ą�[V�Ppk�u��o&6�͇��r�3���)��=�	wRmJ�a�AC�#Q`�c�
ᦰ]X���]�'i9�|V�<+v��f�ŁwK�jy�l�E�J�r��h>���%�в5l�U=�D�x��.^m��U*�ǆ/,�c���E�����9qz�Rx��lS~�g�;��j���W��i�SN�L&��X��cV���=-��uٌ{��:�S���.��:�;�5�ۭ��{z0���ƚ�z��*��B��v�)v6=ʚ�s��V�хt'n�/Ttn�����震ቮ~+PZ�ީ��E��W��Wҭm-W�S.1M��gR[�O�h�ᱷ�����.���go*'��ʶ�=������KHn]����-7Fy`��{1{]׌�*:D�Z���>U��B^�T����n諚�r����iC4j��ww�-Y�'_q����]|���u�h���uYDY��wǽ�+��A̧}%����\s��q��1���f�B%'�%�ȩ���֍Iq�8����v��wpp����tn�ʸ�Nv$�A=��o͋�g�jRp����
��"uv�\e��)qZ2�K�t�.[��q[Ц1:)��q�5�|M�T1�t�\�{}�zKA,��[��}��,���>n��z�f�Rvj�9�^�C(N^>��n�"`�֚���Vy��/ueR���n_,��UR���JUij[S��oZ�ݔ���d�ӹɚQ��^&/M]��i�����V3�g�w�^��\���۵q\3kɊ���w=3�Q�5T�y�y�q��0Qэp1Y���ⱻ��ԛ��au;5���wN�sK]�|�tUNq��܌q���c�X�7��s��D��=�G1�!l�&|+��t� 9�QT�k�y��/�'PX���y���z�5Ys�zu�v��dųp6;:��<7�=Hyf�X��>��U�G�z �g͊��7MH�>�/�pX2������Ҹ��}Udaї/ݢ��'�mf�����m����3�|���#�^S5x��/�]z�
ӷ$�q��QIq����k5�w��w��@c�m��t�>΅װ�>~i�l����	g(βy`���מ�1sܳ���i&%xL�㚤�v;�+����LC�X4L�^+j�����;H�b�޾��VNM���79
��TJ�ɚw�C�N��Z/'_��23 I雷���'�#!��>
S�2xED�%H���&��=�mM���YՀ�3�&%�>��X�Td��Ĝ:�=��R���XRɥ����#w:���N+]���8��]��o�h�ҹ�{mi˻)�(�mfn��e���;.���&�:�{�*+�m�!��3t�s���9z��sٻ�����b��N���eE�vqŇ����3��t'�����jܭuQoo-��r��"��!T{�j+��W�0Lf7��\[�z�\���x�Q*�5�oZ��ǖ���ॿpW�t1���Y�ow�N��z�qm��u���|��|�f)�_[�#4�욫mPZ�k�1n˭���+��^��G�-���z8�N�#,���P��B\�M��:
<o���m>w�mζt�B�I��	�ԏf���^����2
|;��S%ݳw)�>����_!9�W�g+��kɮ���k����������uZ���љ%N�ה�Ħ6����;w�^-?%c։2�8�������)��rX}�P�n*��=S+�9��Ê�c��\�>���G>�}�0(�=�%^,w���<w��Y(t�j����bO&����okݬ��S�	��p8��sm���W�Oiѻ�Ć��]��ڪ��c��;5m_�[wQp�/��v�G8q�v�N�ĥga���Mn:�{}+�3nu����zR��۽���ufj�'3# �.{*�.��2���s#S�Ḽ�X�қr{<.��W��{R0}U�\��p���m��r�# �\����1PX8r���[M����]F4ĩc��Vr����K�ܧ���$��Ĉwʇd-��1^S���^-�9�ٳ']Ū5 y5B�M]����K�NNv�S�q�l�#�%��#��:�/�>}wN���o��!�[F�.�.u�i�Zq��Q�f��w��N]��^�Y�M�Ӵo�Po�L�.�^+����`�?,�S����qd>'�=���M�����
;�m���V�U��aw�����]�9�h�u9��+&c�ͷ0x���/3Ձ�;�W�Y�;�ϫ>���Vl��e�^K�3�����+,8�w瓷k�T޹�ɟRs�.&[Q{�L���<�^��7�̛��|�MG�ا&�[k}��t��������W�<h^N/�{��w_izwN*}���ڷ	�W�r��ox�ŵmo�������ܻ���`�7qz��KSyG�u{�n�uF�sl�׏ʈ=7^S��\O.ځ�=Y��{}YΝ��-���R�|��B6�ȫ���7K�շ���ӻ�͜q�4������pW�ܖ�_����uZa���[�������P�P��5���G���<���<n�ҙ��ѣ~<\��vu�%}p�k�k�a��Y�Ƅ(��b𗃲Nc(�Y���)*d�'_]4/I���%]�h�9c9����:f��K�G3b-�/�ӕ#]�̊�Hoa�ʚ�~��$ل9�\S.t�Om�PR��wB��љ�)����25`Y��]S*�[���4�h����M�� ��fԢ��.��r�m�OD�B�Wv�=G����aˣ�����GRt�e�uj)X���^�u��oI����0�i��[T��[��ۜ��W m��]9M=�yr���q��]ӑ��ƪeU�Q���J�5��\�^{8v<�u����s���\�L)p�ȯ6�Bc!H�Q�W+��=�V�RX�o@i9�ҽ�e�;�*}�Rp��Q�0����3����D��Nrx˭{DL躷&�"�[��QQ��ֻ�O�W8˘��OT�9E�Vk��dڭ�$�r3���˷���0��]7݋S�Sg�������f�v��W��/.�7�\�0sͱ�-�D�(�cQ6��P���E)z�Y�)%��j��o_TE�٤��1G�+��{��u��YK�u�/�W!j/x8�HW����{p��Ʒ+��&&�����%`�4'Q�s��5�4��U``^�<�um��{��XG�t��MJ���H�⽿nK.�H2���~0��F�SoF�E���u�ԏ�DB��,j��[���;���!��}�kfM�qd7��D��2��oGj2�_�����*5Ҩ�|��:�m%Y�,v��Oŏn���w��ǃT�Ð��(y�huF56�;�Өs��{�Y�#3��өO7Xw9�s��8.�+�V#ڢ����:�ۣ�u�e���92`�۵�.�<��/�#w8��ٯt"�w��~'�q�w�')�O�	o�S�b��VX�'�#e�w*j*�p����ж�xw�ʞ?,y-�Y�ӻy���ݝ�qcT�ߜ���N¹11���f(�J͢��l���MJY����]җ|őv����ͬꎕ�	��R�`��s���ᗕB�+n���عxt􄀽W�M�+���c��-�'+a;#|���N���2&������ѓ٘��U��\Qs�	��:�g���qٮ;�oX��u��q��Hq]�zp�{���WQ)�:U�n�TgC]ht��2���G�u=��Xj� ��WM^�� ���苣��!�y@�haxsl.v�;���M2�[�.��tc�Fvʬ���&wfB�ԙ�$U9n������Z�u�#K��_/���j��㎻M����f�l��[w��QC���I)�ẫR���
�>cf���e׸��&�:�{�+؜���<��wm��i.:�^����:5	�n�*�\���/-�ͻX,#}��^e��ĳ6R��є�Ա�.uV����n�7ӷrV����m2T�m����B�pT��9!^�[���ڌk^�K�^W�$�+�ϕ�ߦ�14�"*\Aټ�'ӱ��7c9��iO!��wl��6�lfι��&�ϮW����e����iA�)����۸i�	Է�[��,��]�ۓ��/���(tMb����q�~|��	|M�
ѯ̶���t���P�3�c�:&<�S���;3�C�{�Q�UOw���{Bu9�j�f;�Z�r麦���� �6ʏ�ǹ��D�V3o��۾�~s�]z�x���:k���A��/i��\���<�Zk8��	�}}��������뗘��ᓸ�[�j.��zD�N�7�
�@��>̀�0ɵ!yz�'L
�_2*���/�Y��)�Z�xo��,��Y�����n�VƷ�/�����c��SfRCm`tn+�˭�4�{I�Y��KgtfD�w#��v 6s�n,�;۾�E۬��e¦7��x���Bl(�h̔¢�L�������3υyK��-%�;�̓�vZ|�m_LvfK�fT�UE���	��g�5Gܼ�]ܺ
��L֭+K;�a��vB��D��,�蜌,�b��X�V(�<�f��+��OfU_k��ѝq)�
�q�K@x_����g�9ŲS��
5ݧ��W`����YWJ�΅9΋Mh�,�1���$�cHOM�I��K4��we�͞��n��Q�ѫ}�|�n��ɕ=����M-�}�.�p��bf��NMs��i�Y��_�ܴ�+�\c!��JN)Z;{���Q7��{t�2ꂛ�wY����.)v��T�^�gu�嘱�����/�qۇ5��/ڶ����1� �m.O@��@ʻ�pc���R�Ӿ���˒����ۚ�ʕ�t�[;�h�ӌ����*����F9��5G:ة##r�/�ז𞹥�OX��wP�fM�f�W�V�b�1�=�I`K֮�՗{�ۄ�_����Ĵ@~��fr�T@�*�r�.(�ܞb��Q�2����KC�D��u�\����巷C���y��j�AH@x�
9���&��x���E��:r	�� �N֪�.�k�������҆�?+�!��D�]4H���kT2ӥ�Cj!y�b���	1�^`��p_,��,,^�`!��<+�����)�B�soX�T���^T��8�?3��v�/�כ͎��\45؇�y��������S���!�|�M,�����-SHMr�"����wU�NG	.�1��2�绔������f[޻38!�ǯ6���u��^Q����O���(���S4Il��u�|x��"s�9Q���YO(�/c����ꇳ��ED���&
z5!(ػ�N6��{Q:��3�d�s��8��XU�w�~�M3�I۴+�NC;]��<�����{���Iݻ��� �N�uM�����K���(hG�|\x�A��{�~(v���m͇�4���M�N���iM���PIy�)o��=�v��* �?��N߭ݬ��t����=U�.� z�r"�Y��=��7�z�N�=7�tr`��J=$�ȣ,p4��|��w�7����I����e�tW��uL��-�ĝn�x�$$��s� K{���V��.�R��`�ݢ�Ws�h���̵�\��Ё�3L�p�~f���pQl���eꝷ/q(m1��pu�ϔr&�s�v7i���fcR�-9i�D���Sʉ�U�yN{�,w.ͬ���z�o5�w���#�og���W1��æծIᱱ�y�*ߠ���u����&���zN��,�;g5;���P�Wg��<<���b���Tp���¾��l1R%�ZQ�;���D^PΓ׀Z��LnZR�����,'j⚕�OV"������ޮ8��`�f���R:���L�����繻4��E{�����U<�k�zW����:MB:Ф+������z�ڭ�p���Of�;��)3�]d
)�v��B�&|�<R��a
L6~J[�bb��zg.�k��C�stIe�38�;��Ȧh�K3��p:��W����Fp22^:�&���BVkY���QtiF�B�M]���]��;.��^v��j�e�8�%bj�R��Z4�02��
�+"W[�I�;�J��V�iʇ�ƊsP^LR�C�YEEu�L9i� ��LʻB�(�wp�f���"�V~��"9o�2��	"ӄ�/'�}����!*�hJ
��
!ʒ�����)���j�(rL�L�r¥(s0��(B3ʐ(�����$j�����2�H�(�J��JZ)(��)B����(Z
�j�Ȥ�j�H�i�)�%(�p� �()Z
)
 ��F��i(�i*�b� ���* �
�(������B��!������))L�
��((h(B��P��i
Zl��(F�(
 �0��~����]����l�J�U;��y��k�,V���';�i
����1�<���c�Ou�u\��Ջ��ڱ��|'�p�?K��˔*tC�t_wL9q�)���������#�z��cΎ{h�{<ݫM��/J�y�=;u�_��]0T]Χ6��N
bݺ���<��|���*;������K�s�n>"y�Fsj�ڝ�R�s�_*�gS�K&��yī�ϙc�Y�e_�拷��y��2�'~��ꉖZ��N�u����57�����
je�#�!+4�����j�]��Rs�3����VN�[���%�8��n.G'3')���) |�s�	+M�Jڨ�趞��!ft��ǡ�T5e�B��Z'�U�s�M��R�)���G�̭9���������Y���^F��CS�o�B����Lw�E�_Ќ]�e�	-6��<��g��5�L^*W�v�IØg�W���w��u�0//�QZ��Í8��ᷔ�Uܷ�TloC�LJ}��8�!�9¥*,ݼ��Ҏ&�9�O���qh�%J�BD1�4)�Й�xFk�^������=��G^�x^�����^�F��C�՝�-|�=�Bc̄u�w7L�f�b$�ާ��ɝ�
�x�s,���|�P��zV�~!�b��T��W��K|�f�����w��B���P����rc��䃨��7�^��Gհy�̩=�W��K���#�T�!TsEiS�h��#vw���3�Y'a���q��>j�ƮɯR
b��G=��`;���5B�knx^ORU.���F4&3]�Wʠ�t�wU��jX]8��/���v(�ΰo��f;�t�;ë���1+m5w��[��*XR*Wa������;,^$������z���){}��.�Y"@Ǐ<��OK��zk�O�_B�n:&�9M
��],~w������މn�`ɑ?U�m���ɨjL�5S�!��B�Q�62��g�u\Ԗ9�l��%w�^lN?KmR�~n�뜭�rc�)�i`�?{�薵^<|2�}Z�靭���n��t�݊^(���H>��7fvt����G8+�3l��u���g�ʍ�f��aN�fJ{���0���)��Ȗq�L���H���3}�W����f��
����}$�W	��ۗx�̎�ܗXzrJ��/��S����Tl����o���Pc��w�5���m����ܞ���HOR�t�|����^J���E��{"��샊F��D�s��������&H.3Ec�>�Fb��Dc�^��9�Iú�:𛒮��wwJ�约c��E��U�=F���ע���4�ƕ�1���W=t�or���%�*9F��s���Vj��[q�]�;s-w�3��R��Jnz?^��{R�~�n�a���ۢƚ��
��gd�%C� �?Y�3-�^k.uV���V�zsX��3a�"�s��FfE�e�l��p�����^�q7��f�+�*�C�dr��w*d���\��7�b�M��j�L�˃MF�0o��J�cׅ����CX���/�<���� {>.n*��Pe1�}�b/��Q�q�d2�-+e��<w��{�=X���6uM�&:W��݋ZΊRÔ�9(-φ͝��xFw]s�Q��U�<�a	\�#��,َ��/�S�Ә���H{'���UX�>~��ɘ�Ѭ^�]��0.�qN������\mõ3�v��ڝ��ڴ.������t4�o�$K	���V����<��I��v�_X�̫�])��W�Ö�c�����3�c�Y���@�f;��>K٬���7�>����mw<���{�D}��,1�G�b��Hv{�}��{~��䚑��z?O%�z���4���z�����2�R�A��ђ����Y�o������߹�w��@j^����x��O_����wb����!�����W��7P������}��<��/�w/QO{��:��^xp罗_{gy��{���5�|���9!��m!�`�:�@{/���`�C��vg4.�:�i}�ܞ��;�����ӹ��x�A����ﾨ��z>_FF'3��߂�پ� �u{��Z�_����=E<���9'G�}Ѯ�^I���d���{&G�z:��_`;�u�tҝ���^�ܞ�pz"Dt%?{�z��Ͼs�����|��q;��:����_b��x<��z�}`��ԟ�Fu��N�oM'��^x�C���� ~��y�䛔���z���}1�;�쏳I�V�+W�z~�P}/qϷ��B���i9R���kG�E!�0(%�`zszS��o�#�~�rMG�;�ZC�<�e�a{�x:j~���mN�7�����ϣ�":é7/��W�2]�sߴ-�{��H��:��0�pK�����K�����/%��h�Jn=��`��:�_w|g���Dh�菩ϡG����h{�p=���K��q|���+��-����s�WS�b}�J~��S�<�����!Hd���{�~��w��r��f�����S�y
�+Fu�x�8/������z�&��M�zde��M>�t��6C;R&�u'���p`NnM��N c�]�Z��
���=�tS2�c"��O]����]{��tXtd��e+}�\���[����/[��R���8�>��?���I�P�����r�I��Z^O {�?Aԇ�K���y'�x��w�α]O���~���������}t�//{�%��.8z"�y��x�Ov��FK������>���z�:�}��z{惒�Gz��z��%�R�{���9�voH�/'ӿ�>a\-���6�~ۥ�.��(z=���/�?I�~���<��g�>�/��{�9P���{/��<z�=��z{��)_���]������:������� k@�
oݮ>�h���
�}��莞k�!A�c�e?s�)�g�<;�:5'��d����b~��K���>����u�s|�?xk��u�}~�ٯ���:����瘻���<��N���ozS��f��ې<��ޓp}?K�o�䁩3�d�W�zk�9/�����#�=��RϦ]��f�Z����Og�>�J�ֻ�K��~��rwn���n�G��iq�y��r�������]N����A�:>�">����fT�_�߱��{����=�f<��|�N��nr�w�]+���_�w>A�Q�����������׷� |>އr}/S������aE}�_�ݮ�z:����D��~h���sz2_���1e�1z�?@}/A��G��oC��]ǝw��_��a�C���'�jG���s�����ϲ�o�B�"#�~}��%�7���\�FE+�:ߺ2]�#Ѭ7�,���I�u����~�{��5/ �K�gg��R�5y]�[��}�zG�"Ǿ�t�\�+���u/���~i9r�������:w�+�w�~��Y��j�^��܇�{��iS�{�ϯ��٭k�f�^*���5�V�+y%E���ʹ�|�����Hm�#s/�,�0�yxyk��W�+:|$�މ���
���#"��hC֗;6m��&�l(�*�.���C_�pʜo{�gnf�b�Ōl�'e���)D2J}�=��
����,z!E����ѣ�{�"���뒽A�ټA�.���{�O���?��)��2Pnl�w'�7���.��}&G����^Yþ󾵭���9_����q|��z�?`?�4w�O��!܅;��>�rW�;�ZE+˷��}/�Hv��)��N�oB|" �������ިQ�\���r�>d�e�`��������g�>���h�T�rS�jz��/�rS��<�������Pj^GO�hZ^G_����J����s���
�udo��ε�?;����> ���}%�~3��$|�@�;5�~���^��I��wΗ�܏�w&���e���^��hy5�G����3��
o��}4�E/��~���)Ͻ�P��ԝ����r_��Z�<~期g����zu��{!מiܯ�y�^A�Ǹ��u�Q��<���R�<�Ϲ9V;���@~�}��x.���{�7/Ҟo�=����sHR�G�ѐ9�b�?��\��N���y+��֕�=���/���N��ۇ�)�6�h��/$y.�'7�~��sx���O��4C�������z���K즠���h�|�R��'�lD1��=���T+{��.""G���h~������1�pI���r:9�����xo����?}����p�h=�5�h�z��<���g}U�o�/��+���ߢ,z,{�=���z������]�C�_�eܻ�C�����s��)��oA��Ca�?O�{��ޕ�z����o�R��ϧ�ǕZ��#�=�1�F���CR�Ru��y/]�E#������W��t��r`nrw�r}�c�\}R�����=�Y�E�屻��0C�w'�R�I�H �I����j�W"�[x�Û��kR�3����y@[Jn��t/��o�t�A���9[�>�MI��g{
��}'�a��.��<�Z��[n�/�+N��*k���H��akse�	<�t����y؝���%M~�D�`�P�~ޟG�2N��}ѩܮ��XR����_�z�w!��r�_��b��G�����rC�q7!��Fgy��ߏ:��[��>�q��w���/�n3�^I����`�A�~~ѐ��1��(L�p�������������?O��p�yO�~+���,�Xn��}p?@j܇7�JrӸ���{&�z9��w=@v�rw/S�Ú�<�$��h����o�9�^���~��'޲b!��z,g"O�է�������b�!ֿhr�*}=O��8}ޞJ�<�oI����>�K��~w�j\����Ծo�2)��s�>�}fo�P�C��=��Z��+;���H�����}��N���C��h2}����y>�����+웎��I��W�|�Aܿ���}�9�z�5����ءŹ�T�?�B�����4}�h�}�>����ݝi���z�w!�^��J})��4{!ܛ��1���?\��F������޴���(O���}Ϻ&��Y�vUq]9��V�ހ#�=�&#�>O`2~�Fu���ђwH��ZC�9{/GX�HrO~��&�=���;���B�Br:��rG!��uw��m�}S��Z���#����y���}#����he�btsz�F�׶�y/kFC���1g��]g4���y.�r?y��u/ ��g����|e}��h������!�`�Oj=��=k�H�;�?Hy������]I�>�@jPto<���}�����|� x>߫#�|�_�n6V��K�:���5���G�a�K�){p!�/"���@��w�α]O��i>��b���H{�rx�搥�t�NJd��挃��_$�~�y�{���z���v�|��繌Ȧ<��~�7JS�O.�F�E)nL���{kEzLRn���ʷ��A�PA��Wyeѵؽ?
t1V��Y9���|�A�s�Lrɬ��-�q����f]��!�isy�s���8�ШSui�9��_S������a��ӗ�q���=�׳����"����_���]ø���;���������������'�w�voG����O�K�SP{~syή�GU�A�k.�t��Ԥ���`�H�����O�vu�y'R��~��z��P����Bs�O��y�}oH������r�����{�Js_]���k��[����=#�z����==�h�����	�~�R��ޱOd�^�ީ_����.���������v��NLC&*ϽG�������M������_������܏�����S���_5��\ђ~��{>�FK��	ޱ?AԾE'z�?C�z�z(_��w�/3�^�y�y��n���tA�p�M���!�joc��hHn;�4�������^��|�$w'Pk�d��3v!�|�����|�N�`���������D/��Nyf���Y�Z�x����=��_.{��<��;׺�n.O��)NF�sG��_d�>����/S��Ϲ�;��;cN�yF��%� ���#�G�@��{�������*οoϾֺ�C�u�}��\�wnq�X����~�rs��;��jG�9���/���������3�"��DEk� ��"W��z2w���w��w���׾��{����^���~�ܽ=��H�?bu��~:��'�u�r�O����w'R?��;��z��ߚ]�ܽE;�����^u�\�����}�����u�N�����/��tϠ=��b���C�g�r��:�e7'oX<���_#����G������b,Dh����qv�VOM�Ò���}�>�����I�^��)����2^��Fu��N�7����=��}&��{�r���9�w)�h2}��!�F{Lz4{��X���7�o�}V�=�N�z�fPO%��{=לm��S��͛6�)��!�q�y_3^�G�Bʳ屺;���j)��W������7�'�>���cWc��:P��}v�ӷ�ŎrTo:1a�dLҵ��ZӛFd��mcrDUu��GW��qdNjW[�����_��{<�9��R�ɑ�>���}��޴K�R�����)�7ބ���>�Fu��'g8h/м�֐���P��콟{���{���W�e��ߦW`���=��{���끗����C�5/ѿ��/�df�9R��sZ��)߹��=�Y����NK�u��gX�%��ZH�X��<��G���v��hΕ��w�k�~��'r�?>�Cܜ�����}/s�|?bjCq^����7�NT�#y��_3���M�^���^�#о:$G�������eM���B~�g}}��ٯw��$�:��2C�;�%�x�H�'�h{��=���K��>~���/p�+���w{�';�u=�揤?Y)��4���u}��ϵ��}�מ�[����
C$����P:���2g�����X���y�%|��δ��@�~�R�)>�C�y۽����s��Ͻ��\3�_G��~����2b�+�K��GC"=�G�cG�8G�����!K�}���/�{!ѭ�}���=O�`>�Rw�t��Ob�tw�){=��r�0�}��ϺI��:������G�{�<�F��{����'��=�d?A�{�|��W�߹Ӑ�&�:��=���X��u/G{�J����iw.r���7�:�{�������B�D�#��B"��'{�JnC�ٯ�����I�<��<���O��=����<���9Py	�X���_'�xu�}/P����_��f�|�t��u���=�P����>��� /��1��%�7w��܆�^���C똛���^��3p��K������Y���������'Y�y{|s�������8�R��	�>C�����G|����ײ�N��~�r������Sp���s_N��'%�9�>���w_`�A�<�3}���~�K�̶���A�q@�-�aS+���C����M�e����w�����Cٮ���R�"�W�`�)���M	qv�|�R�3Uc73����G:}/g���a�h;��l(��&�W8�w)3��6Й��*�6������y���uӼ�A#�c߶�H{P=9����Ȥ�X����uҿK���1��z��'��7!�<���L��ߚ���&���|�}�_asY�3m)K�`�X��{G�&�d���R�����%�R�f;���f/f`C����w!�k��wb�'q�C��hܧ �;�ߺr���3'��p�\�ތ��}�^���;���z]�ܺ��g4%�s���Wpu�td���Xn�>Yy��$�w�#����r�o�j�g*c�]�gB���}����=���;��w;���W����{=�y��NCܽE=��t�%�;�R<�~a����f�>�W���.�?C��[yIEܽc����u���z=�=z���r�NA���K�v}޷+�;� ���'r��O7ޓ�����}`��P�X�]�ϰ��1^e�5�n�&:�,��{� ������Y��jy�\��; �}��9g��&��:s\������E+�g1>�ؤ:��NC�f'o[М��:��&~�������Fw��3����=�"(y�5�?I��:����S�~�|�r������ܞ�JK��=�\��r:w�"��w�h>���:ֹ����f�}�[\�}�K>�"$G�����$���z5#���kFC��q�C�O���M��z�/S��{�����>���7G�t�#�u���(�-�������(��*�7���/��<����ԝ�>�!�}��ԏ%�zӓ������z�|�e���;���:��@����u.�ϭ�4v��h�V��_rA��#�=� |�H��v��I��]A��4}!�1NϹ��Od�;���4�!�yt���s��rr?=b���^�<��_j��U?���n����\FRr�?��[�)w#��%R�r,贻� I`�͝�V�t��Jc%�Ю�F����xuf_ ��]Yn�s��O%ۍ
6��2+�l�����!� =5��t��Lck�Q)��-�U���X5!iB��*��Ћo����Z�j^Ui&��|�dκ1��{ThK�ޥ��������s׫����3��V��Ʉc�y��_O^�G�c)X�"�%]��A;s�ڡz����ʲ�s������j�$$hs�^��JZ��X�*�(�6Ɯ(��T�&��z5�M�ߐ"S��*ʲ��];^ه�_-���y�J;�_��hǢ���#!Ӳ�ҡ���C�|�	�S>3�����=A���Gm�����־�z�D�����;\BfZ��6�͙���{Qm-����h�v(��{ѯ���׼k��RzA��.8��{�:歑a��Q���=���&�{����sc=&�{wb&��n,��L63���/+����)�\������>B�ܼ��E���fӽnp�\��Γ|�y#̝���`Ni�&����=�;�� �M�WN�M�ҷ����ܹ�Ƞ]ˈX�O^���A�-4ܹ��^v�w@�̆���P+N;uY�)�n�zq�Jb�+��F]�sq��h���o��K��-TX�M��3V�f[�֘��^�f[̦	�U�{{dYEV��K��tH ���F��wǲЫ��<R^�OIs�����U���{�!���%o|�9��[oy���q���=�
��s$�n����_K<tܲ+^+�e�֭�Eǒ�`����8����\ˌ�Bb�����au�/اl���<Y|���ƷS���i�&l�Efv�6���C5*���l�������� �P�ɇG��k�J�Lg#��R[�-�V���&���lid�/{/��2�r����"���!֝�(�}1f�m
��k3�C)Ut�h-�1��F�!�tiuvB��7E�g��t\� �p�?1�p��r��|��tU���`갔�U��Ƴ5e�;`S8���1��}3b���1I��Kr�O6�Z�������mo�Y�+9K�A�m�ZrQY	�ӫ�TG�3g6Sׁ���gDUD��x ����KJ�lP� a��aL��J8��R�C�U˘-,��7�S��K��em�8,\?a�� �x1�6X�����fe��*�k�w�R��Fg���kc	yY�P׆�S����%���mpwP��V�ɁJ2u���	���p���{����];'.���)u�[�R��]�R:��{Ce��h!�6�g�+�#ġ����&G]��v���"\��CsA;Z�ڢ�F�8M<sȞ'.�0����l���FD��a�.B,��S�(
&f
�F
�
��Z�jEvЉ���:�ϔi(����((�$��L��0*�'#��$)��(Zh����*�
��h"2$��*��*)��0����\�231�%2)*�(j�1�rc0)"!h����)*�"�%��)[2�jj�$ȡ��a�%*�h�����*�� �Z#$��3%,�0������22,Ī�2L�l�"��&� �h(�!���Ģ���02
�j��r���


J�"���I"
f�""��,�j�)i�*)���()��"� �����(��2h�!��I��A��tJ��*<�1ҽ�9Y�w}Ә�I!1J6���R��!�y�e�n!���4H7���pxq�� Y�]���|=��ү�g���L���{���_����t�����7�=�5�|��7�?8��1�7EL�6S=�KY��Z��v�\��l^$�t��kU�Wl�g25�k�=	��n�r<��XC^1K����b�ޭu}�^zt���/����2�0�+;.�k�}r6�E0vv(똊*:�1֐�E��m�,Ha��F�4rUް�N.��,.�S(6�[�g�q��/�c�$
^vs��ʅ}N�x�cA�z4ghJ�c�~��FP��ʼ8����/���o��F�l�5��T�����2�U�ne���?%�c -���B�/`���޾Jm�jb�6z��p��y뭫V��[`��Is7�����Ώe��u�;t!�>�3�6d��#�,c��ҝ�=����B���b������r��8�`ubz�}�W/j�t�1��!��s����N1q�`bM�Lx=<DAf��
�u��A�Y��EH�c�w����<ȇ٩�ߓވǞ�t:�ي��d�Ÿ��^'2�Kp�8M������f#Қ0����,�ۡX��9���=O�S˂�7���iԵ��q%3�ވ����A�[\�GRK�c�n��b8��и�
S�*1�,W���YL��г�������cq�KlJ�.���Vv�1[JY���]Yy/9�M_k���1��N�'�9ő�|�od�tf��V���}�d���JT*��ݫ�����)�Iܾ���+\�VM�-��}�S��b�b�+6��ݻ˖�ٲ��-0���eE�͸�tD���Xa���Z�e�N:����Ei=����F_�S;�]�u�׭�=Tgq�T��ZW�h��Y�5�Aek��;6��Q��v�&3ZA��sw�����Z��{����+2;�cj�}A������n��Bl����oc8?U�gg�s]���p�n�&LAC�#Q~:�S�sGNN����{��w#��e0���J��9o�8}���>L'^,t?Dp��`�[�[��>	�,r�06����vS;{��͜"����0�T1v����Wn���d|��!�]+�v��>`��E�V�Y��k,{�)\R�^�J<Ѣ�{p�(�2���]Ma�༥�I�[Vt��Q�$�X[���{�lb�	�\���;�E��kg_��k�z��u*;�X�zn�s.�g-.��22��9ϫ�T���׼S��:��π��'z��w�ŕ����F��bǇ�NX%/% {{έd�Ⱥ���E�v�X^�8s��~��:�nL��%[�q��JڨO��Rp��묋˼����s�;�㫴Tt�v�`}�m�	F��^���S�a�d[��Ȟ6��]�q{��
Uf	u˄���ۊi�ȨL"�'��ǚtGN��5Mjah�s�ĺU�n���Rp��Q�0��@�1WS}cB�5[�7=�ݝ��sՄ,�r[�O[���M���
�ͧ�71Q���c��yn�V�VԷҔ�uʣ�*����<⡬ySՃ^ظ��3��>�f��k��k6�
�c���sq93�o,��Ơt�G"{�Tm�3�j��b�̺�K;�pN�A�l�d��<�-m���=�!w����Ėj�AhF�����r��y���ŕ;w=��cϸ�F䬖"���X�a�Jcǻ�P�Q
��8�0��\�ǡak-k�Һ���Cr�Q�zz,o9������Qގ){��| ��"vz?Vk��f};��9�9sw��sX��;��ӓ4�dpFU��R����i�U�,ufW�~��O�����vˌk��Ԇjbo ��3U�u��"���V�Ǯ6k��ƅ르�QX��m�y�K����\G\�:�ݤ�7Vr�e�7R���|;c%ڴ��<L.X�>���0$��{�>^J9��tweK�WAm�SNx.s�ױ,�\(K�72�*Wn�2�U�J���(����<*!y&6�P���>{�c��)�ڇ�d�ŏ76�V�Ծ��6f�R�hhG;btN��i�bZ"f\�x�ļ�,�_j��K��׮r����HL)f(��7�(W�긲�����<�γ��sk���)��s�P���*faȕ��^<{5g�������B�g�ҭm\)�k|*�lu�G7�;�ڋ��c�ߎ�� i���CM��<+D�S��W�+t��#�}b���C�𤜚�-�x�ꝡMz����G���Щ@���l>VJ�d�7��J���c�Rwݗ)��DC+jw�/�N�I;8(�9�[��W��Q�Gc��}��G���N9�s�5�>����3��VZ��v�0��$�ӷ�A�T��{��������8��~;yShӕ�r��nJ��Z:Ԭ�<��j�v�-Q�ݝb��Q�5�1�ˤFn���ɻY^�o*��{x�������c�4���˽g<����^ث�<�y;���1Ҏ�7-evm)P�	���9Ee�+�c�N��g_�f�Zzr��1*�m���Q�,����BZ�\�LVrB�f;|����z�f'�J[x�T�����U}A�%&o ���b�m7����v�_ ���G�o���n:WKѵ�)���,.�;*���T�:�=!��Xũ��Ov
m#��ϔ�gN)�<��x\M�_�L���ݎ��_?-g�w�$��P����G�iN�W\b�-���xL-��E6��*m��=�`�NCr�q�OӯU�~��M`�VNd!��ˮ1�P-zh{Y��qdz�f]���s�>�U��X���{�4|�YNzs���t��Sb2�+��n1BV�����)��g���R�O�w�{f�\���x۾��>�o@j�~�'����W�Q�$�:V}Nզ�[�3��[�T�`ſ)XQq�Y[�v1*�#����w�d|7���5���z����f��[J��lCl$�����m��h��̙޲9�������dzr[��7/���u�}�2n��y����faO&T��C��2V��1Le,�w�τ�RyB��;[��i"��q���$l*eW1X�����3Yj���n��J���u��MoLu5��'���8�c���^�Tv�-��y}fƞ���-}ER1'u�z�n����b7B��	�'�9ő��x_x��:���9�U���y�o֩�\����z�'F�k��˚�p AWy&��Mv�K����7md��E����u�\��'�w�;�f��:o>��1��N�{���g��������{e��Ϣ�R��uy���i�j��X��7�T�WCT�@B*Z�㻃6��/*#�Nۻa[&Znʡ�eX��Ffvo.�J��;:�\U���z�}v��Jv�ybͩ#XN�d{c:9���U�}9�GvNTXz�Z����2�m�m;�+��9�)��,���n���DG������w�e�uW�'���ݛ�෣<_0���YN�A�2x�=^'��75�o���˩���v%�����i��%���R�y>���̓5v�����̱�ߢ�J�|�x�����j�{��f,sɶ�s����9��2�\q�����j����oz���eX�)�ԝٕ����2�$��j�Pû���q�.�\OSį�����զ�\�H�ͤ��T�ū9M�k>�߽��X�OW:K�lū���W�����/1�Z�0��OY��*��T��]z3��ʜ�.���Kb�z0�=R.~�o}
��W�;��r��1RƼ�����ĭ��� v�e��N�=�{S��i��!UD'�T�w�Ey�1P�*D��Qi��w�ٜ��c\�5r<jˊ�Ց��2
�|4���\TG8�'�1=b�7����l-�pg2�_	[�ALm�e��Y��C�(W:���T,�vj&�����Z;؀�9K{u\�1Q���Ξ�.�[��Fև[��G�ey�6��[N�x#n*����c�`�c�R�u�vLݘ&�ǰ�+�u�;	-ѥ�q���kmԙ��+�G-�}����7o�L���f	�y6�)]N�� �|V��YO��ș_�����x��l���c����q�4Vv�9����<βw��Dk%��񊹌_�yu�^�x1�%btSkgx��W*�;R����ԯ,:۫�6������JZ��ҏޟV�z�ON��Ĺ��6�NԮN��=�%��2�T����sg�j�<YO�Z�����r��]m����!�[�ht����@�y�e�g\-�ٴ�+X�'r�ǧ&'ѡ����}�-]Bb\RQ79�^�%RtwV�4�,��5�Am&+!�W !C�n9�}o�o�)�n91��v�_*+���7�1�.���f��"���.�����B�83��b�t����iĭ�N|^�(=Y���9L�����p�����ʙ邸,�v��w�-Y.�r�햧�N#�Qyo���8�ܟJ�x�6��>�}]0u1o´ۖ�c�o.�
�쭢���e�ZK��&3�2:v�qn��97g����5j�/�*bk/�N�^>�(��4r���	B���G"Ī�Imzc�-n�ߢ"=������M+�\ެ�U�M��jJ؀џ=�
��A��c>�{���$�=ZBжJ�;'�#-��:�yw���Cw�\�*s0�!1	�k��C5�{�Nff����N�>�Ꭳ/+ehޕ�ɚش�_Y}1�$5Ch���w��	ƶ4uO+M����Oe����"��3�d�c;�vJ*��;S�wv=i�b�B1v�a]\��j��-������m�}8��;J�\�:9*u*�<"�,l�h��Z��Q�Vv��9�Te�{Ura�dnB�m�ܛ���9��}��]Ny��Df��5sk4�LpJ4՟fr���/&u8���V^���Z���}��]ִ�R�ni��&�,�<�6�>�����6�w���]�ז�*�=9m������*Ŝ����t���!�Wq�iS���^�/��Ht*�O���W������&
��d�luc0g*Ҳ�e�Fs�G}��Z��	����`G�;I~�eV��G���jwF�2�rrju���8p�'Kԫ	0��Zx*�ֈۧ���*L�En�֏���p���(���<�c�9����U�=�i���\mW)���D{��S��'ת��Oޭ�����m\�]T������^��9�
�>���^�J�����ߦS�<�aw��uK�;�e.�7�RՋ��}Fc-E6-M.A�K���w��&���LW��%�a���q�,K6,ݰs[X��PЬ���]�mr���S������É���d�����R��b.�]�_}=_R��d5�m깴�K�gc�T]�VZ�VX����*��h�~첤O����\�����=�*�u�9u8<����$O2�>\DP�ߟ���/��e�5�LNG�����EW�s��1k�3�93v6�-]uCU�1S�LBb]Z��x\�گ�^u��2�����}����L����+m���W��+�g�i��|xq\n���(��gtn�w-�=��܁���:g�9Ő���h;K�|�B�Q�7yei�lŝg�Yg/�@Z2�ئS��:hb��)*�^�&��{�;^U%��;���h8\S�����bv��4;�9k#S��Lt�Z��-�����"C�$:�����X��v$�� 7�������t�y��iN}X��s��͹���Fa<�`���z�W�����a��,���sHHK�Ъ��79+��Wv�4������C`���iݫ��ĩ瞙��vt��Q6~�l���\#u��㖨#j�ۗP?�d+�t�yp,^��y����&+w��I����*�hr�1��q��aYpt%�.)�)v������؜Ʉr*k�X=X�
�w:��y�9i;��;���R.w���
,�6-�L� ��Ჶ1���	!��:�k.��/g	V-_N~#��G�'0�0;��y&,ѻZ��
�Aq}� HΩ��A��8��+`�����xz�|�]6���:��&��H��z�����idډi嘮@��)�oL�
���j��Ҏ��o)|����+˹~� �ӱ�����Y�*!�����]3����nT@�M�b]���8zA����4��xY���Ť�M�3o��n�%��y�	�̺��$�H�֢���7���b ���-ww@� 8~��V����}k���!).�����+&]S�ꋝ��8���"�L^�[�[}�����u�L�fN��R��+�6����G�3}�rJ�z� �˞�б>t�[��Ykc�2ygQr�,��ss�t�k�52��+��1�	�ǖl�SQđ]�v1���^>of�v�+�t�;{���e�uq�'갫5�Ev`�Nv���6X=��˫e�;v�]�%�,�/)�`�|�k`=��Z��r*ڧ;���kt;K��"���v����m�#�/��B\�ͯ����>��2{��1ES�z=��R%���`�W�kIm�H���&�&��p֞�w���'f�o��Nv���f��HɆI�oE����GhY��	f���j��.%ȩ2���|�f۷"�z�Z�f��_�d�Tf�F:�Y��.m`7r�5��#A�?���J��y���bJ��V�\�m;o1�`�}�Ʉ^�ݖG�Q`�s5�a|!ԕ�8V��;��hB[LVx��'��;�X�Τ���R����Z��-�)�u%w����)�)���m]���4��0�D��1��c1t�Q#C�S^c��v/�]Gś�S��aɔ����HA�QȠ5���ִ�T���iRy�Z�F��-g�Y,X��ح?��J�E�B��D��Z+R��iF��a�?ZV�6�M��\gEu��.��dܬ"bQ�.�EOQ��W���@Pf��Z����Z�̩��� ��j*(���h*!�"�
����������(�1Ȫ**i(�j�
*�d�*�*��"�H�R��"
�""�h
(�������(��*�H�"B�i����������*����(���l����������'# ʀ�f%���������*���b����	f�j����(�"������(*������̓"��*����)���������!�&(b�*�"����b���(�)"��� $�����2���)�(���q�
��*(�&�3#"bf�B�����&�$����b
���*�30"�*���?��vv}�~כ�c�y��p,w+-�-o��"��ku�M�e/���|��[^]��w�"��Yӗ���r��ff������곁v�	�g���=u����p&kE¼"_ c��K�kn�)��h07�g18�H�L��m���N��Ee���S�Ѥ�G:��S���7�-�L�uK�ǂ׳hH��f�ɶ�T��U��6TW�11p���S
7`��Y�<\��NO?-^��ŋ��^o�˶�*�ޙ[*&��H-��z�M���{�ZV�'�q�__���\%�Z�]x�۹ɘ�MG<:�D�4�ͪ|�桎;���½՜��w�E�m��)�V]��/�J48�~[�;�����FļaO��N��������jj%��P�k�˫�6��Z�sUp�ۚR����v�1*w����^��n�65���XP;�9-V;d�p!���a�u��>����������=��vQo]�*^Ozs!c��׳;���)LtH{b�r�+�W={]*�h1�@���f�8��.�F�0ݜ���]�T��آ*
՛e	Bc�1J6w��h�d:u=����z
�1Ȳ�f21�9�X�M���fjƺ�4���s93��mwZ���F^�]�t�귀��zs�n�fB4����{<��׷ �9�_Y�/:��{[6'J���J�&K���oT���G���<Y�w6���I�=ە_{�;��lx!J����+�:����-�׬9w�+N���;V$ٚ�mVՏ_�R�O���_9[5�h��c�1�����6���1��*w���K�.�㣛يN��PSQZ�5M�*��盛e��Q�97��*.z�<�nBp�ڎ�D�lHsp����j�<����EӄEfߎ�T�g+�9{Ft4�7�{\�t�\���ζ��R�$8�@�ĝm,�G%�S�Ҟ����^/S�6�i��n��j	�4�c�ĹOqqۢZ���p5d���o&�eE�y�C��1b�W-��=~��J���톽1�Y�� .���{e�X�~<;�1�CY�J���j{�����5�@�9��W	���毑��E�+W����c|�W�z^�������8]���ʁQ��t$���N�����g��Yp��_�����4���y��ZWB��_���/MM���`x��R�6���Ot��b�}�c��� 5�]Uw�V�ڶp����VuoN2������G��� V�_DG�=�	���/7u�"&Oҵ�ŎS,_
��W���|�}��a�pU�Yl,��"��S�i���dż{ZU��d�/�a�0B�p*N�n��D�q�q���b�҃|�LV��T\憣�s9�k ���t��� !Ҩ�C�,Gύ�\�/eg��
w9��F�Q�ҭ�T)�vλ"+�z��褡@��D��*t !5�-u�Y�Q����x��ť]g���k0�dCY�b����,�2� :bE=��������f�I�	<X'n����"(<�J
��l�����r����7a�}J���1<EC�B���m��{�eU��tK���8n��w�a�+)�F�����`��k(s>�]4�>��˟�K�{�����q����N�}�OI�O���~Z��;#�#U{�p5�UN��`ʎQp+=O:�zp��\^J�-�qI�	�\�es[V�e��W��/o:���eWe�C�t��l��d�m�X8|�x���K>U�W�+hxJ����7���Ny���{4�9q��£�\�r���[0y�HdLTн��]hY��"���Onl��[J*c���iU�֐�`��*J����ޡ��Jt���j&1ì��WN>ԥ��'.�.��A�#=5;����|�T� �ڲqY7��:�#*�z,ߣ��{��{�=����L~���V�6����Z�'>��Ad����B���#��JЉ2��g�@o#�k�;\9"�\�Q�4�ߴ�o1�l�1]�z_%6m��
G6#Ҽ�r5g���ĴX�]��>��
��aƛ�Nz�����X�����Y�U�Zܿ>Wql�QPwiͥb�!�FRqi�W\�İp���������&B ��w޾a䚴���zj�~/��K�kc��.i�`#h??��ʉo/�Ƕxlf���t��39�nws��W�Q1��1_&�1�ؕLW=%��4GR���1�{cl�&'s��+�T#���1P�����i�ʐ�N�(
��\���sݓ����Ă��M�WB�߼a[��)㑪&x�S��r�K�7q�mGJ�Q*g+
��{mD���Ys�(�&xhD���C������1c�������F����+`JLvV�ΊI�is�*~�Pc��}p"v�_�������ÃW(7yA��s�g�/������m�ie��YV5��j;�M6�T�=�0Kޓ���>Ef=��*��>у��+i`���>u9��2��n��`j��Ԧ�oPm���{�@9�D�c�Td�c����kL(�^g(�;i�_�>��1��v4��۲���ҫ�| �|6�l���nYl�5���4���C�K��0��%��|oK�4��u���ݴN������n2����u�C`[�Z*/ԩ"yH�a��ӑP��"���g��9�'�#홋���)p
�R>���g�!�V��E�i]�4��/��<M�C��Y�m�S��U�W&�����hq�[9$�r�$�q0�*����&��J�4�dB��[ӻj��4�r+`a�8~�u�ٖ^���5H)8�)�`;�i�Z���YY])Uo6����"P�K�k4�x�{���j������ᒰ�}TB�<�J�[/�A�:9����mo+�����h'6�E>�Ul�l�P/rPd�a�D�y�i_�=��]=��3ƱLX���X��S���ҍ��9�
�ä�T'�T��*:׾��ܼ0.ލ�쑨�������9��V�s�o|Ӵ; �p��z�����1���P.:�i��(��+���,һ���s��\m����vp�H�xȸʙyY�ۮ���.1��������{s�<:p�G]��ۤ�-�+��s{�a�B��\�-��xZ]Q��8��3t,gط�L�rX;���OT�۲A���Xu����C���T�}X��S�Iٗ]��Y�WlEK+���y�C7t?MDz�bx�j7�y�P7|̦{h1A���}n^�]�� >�}NJ׉=fr��:>��@GYh���9�0�"q�� K���F8EzPu�yB�+.�v�X���T2��d\8�AS(lK�J�ًV)V^F�ל�8=Ƒ���q���9���;ÚQ����i�<��_Қ���]��^N/s�b)k�	��l#X3��s&{k�Xq�,]��3�0��Is������JZ����W���G�!�{�r�/RFc�w�V�b��<ub���^�.i�E|a�(�|�b�~̇d<���k��Zg�^9���$(f��Cn�l��V*.�C�Kj'I(�'�Ղ����m� ���J��Ih��[�{6u��n��؇��V@�s�ơT�#]
�%Ý��;��k�
��.RX�B�R���� ����t��� ۘ���jbS��aNǥI�k�ļ1򻣠�^KM��(*�Z7e�f���@0����1��i�}���� W��V��<�׺��}^9K�j��1�Pq1����|p���x��wY�Ż�)lSG�ZE%3�M� wN�b�OԂ�1��-!Ov��([No��w1����e�=�y��2���ü��j��̮A���Vpr���T���K��O}��}_R哩�f�U&z�c��)����'u�v�]@�y�Uo\A��c�>Ϛ�.���'�����;�j�tnն-�@P3K�a��ّx����E��s���bH�[�YldT]+��<��r��r<�EEf�(�Yf�J��C.��}[��g��S��q�eyq�b�L'ި����2.�W
n'�E�p3K U�	���V���r��Ʀ7nw���_d�ݽ�V�;ԁ�B�M��*�������ص,�q��&��,+��V�romq��Wx%�]Y�ӧ�<�Y~g�ɧ9K(P�@�KAb��;���<1�3��@����fs����Twuj�ktw�Ϗ��k֦ z�����l�A����(?ST|�.�\oӷw�����1���"}7��
n"p��d�OAJ�KK���jý��~)��6�ZBϛ�,nSac{!��0�	����2���5����.�~�X����e����<�v0�<"�g�xm�Oa�λCY��b���3�Lk�D����j���C��sg����*��C��ԭd��Nd�XX&�^U�x�s�(��@�����ڽ��o�<�2sU��I�\C���"KӼ%)�l��Ɣ�����&����=�k�_V�[��R�z_T��ej�J3��?π�����{����
�&
$�b��2�Al��t ���`��Ї�㣓T�X��!�Fgp�Y=�M�$P6l�k4Ǭ	�x�r�*��X/\,b:�V0/^�c�˾��q�����]X��t�"�:��ZIu+�1�=�'�'U�k�y��<i�*|Pg&�W�^��ԕs� q��;ă].z����K�ޔ*�Dx=A�im����W��%��'�(����|k�%�Lk+�i̠��F�<0�pl]g�YC�b����/LS[�θ�z��2���yr�ϭW�äxh�c��ׁ��$�,:�VB��$��~�^��/{��"��,������Jc��A3���0F��N�75��9=�m�.��3����ٝ�۹blZ,Q���u\��7�i��ʕ����'���l��qZ
or�NP��ޖ6#����bX��9��٘`��
gS���\I��ޞ�3�)��;s}՜�o���ĺ�-����E_��C�"P�4Ua`��PpP���&f;!����D߇vfmY�<KC�9t�ǐu�3'C%�n�^@�����g�l��=/r#c�NMf!�)ʽ[BlV�f�\�˝��8��͎9������8]Ď�mzi�dK�#S��3��滻�S�_�{�sKƞ����T���=�Z5��{!9M�p~uu���[ֆ=��7l[��^�%@����wS�zOd5�״r�$��Q"�����k
�uA���!"S�5MB�ԃ6ޛH�׽=y��pvxa�:��T�8-��.��zVDK[�.*�0Ó(S�1í���%q�׈��̒�yb*�8��%O$"�lIT��8+��iC^v!u�`4���{(�|]�5�[�W�P����s�i��d�<�J��ʚ����R�#Y~������5w�irn�'��5��RE�iΉ�R��ĈU'I�'OL�'��
>�ֽ�k>�S%�ྒྷ��5# .���9���$ו�^UF���ߦx�ެu�yNpW�Q���Ô�.c�cGS��R�w�I>N*�� \"�h�J�"aVa�<�fr;у$�g���4��>mb��o&�y�E87pD�N*y>�&���$�q�L�=�R�kst�s�!�D��9�f)����2n�_�>`o�!C]�u*��K�*����xm7�P��qfU�U��Z��6�y8����%͈Eკ�X�veMR�^�[����X�D�A�Y����|/I��8��m� �`_[��۠H�-^���\����ڡ�V�z�+�6ڰcF��ϗ]�en�_�}�}T���z��Jglh��c{jw�و��YȊ:"}fь�L�k6h(�(3�g�ש{Jzf,�|s�}���}��u����d�CeT��-�gC��"h�KNt�5���G��.П�zPF�^~(s:5���s�%\7��0*u5����/�WZfn�y�̱���7�t+��]���{!҂Fژ��R��E�BoM
J5�w�Ģ
�5�o�y_\�]y,N����m����9�����R�ڂل#.��̨�����l�s�U޶1��r�*�L�b���O/F�E�R_c�C����+CxqR����Z��7��	d�8C��)������-L�����(Y��.Vzx=p�\ά�=�EH��6C,T�xN�W�#�D�;`�gR�}r����M�8l�'��}�"���{�ud��He�jhTs��%�
�aJ���xzD�Qv��u^"� �Y��/o����3�����ۻ�*�Ш�t�f,g�D�3�|D^�}&`1 I��:��ԛ��)�{<�K�sY��V+��LN�ye��
��w>�W݆�͜VO��4yٔ�+�Z`�&�-MS�Ǎ���泌��N�Y�����{���р��V����]H���� �e[���Y���L:<͸�'7i�2�)�{stp�(��J��Ns�fv���>�Svm��.y���2%�J��3i\�&orz��t��D>c��Kb���U%���*4hB��/��*J��]I䝇^N�_/�^�����s1��ͥr�E_T1��'obQS�f�v`������e�O;1nl��ʊo��oل��|�2�F�p�9�X�j���8�ol)O3�G��L�]sk�"'�������u2Y�QGӨ�#�����Ѡ�F��	��r�˙j� �eP���Y�'A/����s^q�*�&��6��ҎB+ۦ���	1�	�¡BJQ:q�r���Tנ��h�w���b���F�y�1�{G�T�y��t������ϒv͡�xj"�ˬ+�s��q&m!l�����=�h"�iƑ4M�|{ob�{"Ü�� c�J�j*_K=���Ekq:gy�M�o1�]Y���x���s&�G�;-K6�3�B�k�b���	�(�4������u.u������u�3#�!�N|()-]�sC��V�qA��#�[�Y �[�.az��(�\^N/z�5�ï"�b~���#�$c�3��
���rΟ[�}ݏqch�wf��ROTN��WE��qZvsm^:w�:�Ƚ�"`͞;�ˆ�5#N����(Ш�<�ԘY1oe�1$*���=�6���d�IY%%_`�C/)�����i���M�;�Vw�-��5�w|eF��O��&�f���5۸�s;�Y�ǣ�l9�����;bh�o�;��nK�$�z���B^�-;Nb��͢�x���mk������|������j�9=��u/z]�����\�`��X�m��r�W"}��U��Uzʥ����+��W�dk��z��F�N]Y=d��o�L!���l��F�j��5�b�*����V�ٻ@�5�9�׉�гaK��k��X�&'�ԩ����Q�C~�#(���|.��{t��7گ#�P�-Tq�g6��YO��i�V�����d��*%�Kh�ə��t���*�NĂ���ǳt�ôx��/{ۺF\�(�9�R�TtSz��iiz�e=ʹj��.�P�|D��
f���b������ԮNs��fM涯~u�(	��5��#�Aw�Pjmf�IV�0�G!W�y�D}�_b+׼<�^vPr�S�)��ι%9��pT��,(+ܔ�˭����fIe3� 8�)#{>z�+�1�@[�.��47���f>�`�	��y�nZʵ"�Y)�
i"jb*�)�bh�J����"���*"��(��bj�	��h�Y�jj���*���	���*���f��&�����"d�*(���.�&����*i��j*�����jb���������h������J���J&���*��"*���`"���)��(���������
�*"b*"�i"���)��"�f��*)�(j���������"���B�B�b
b&)��������b$�*)�
��*b�$��(�J���d�jH���(�(�&�(�*
����*�i
(*��������)�b(�������(�)�i*��(�()��(�)�����*(�����b�X����y�~�=��nb���y���3=X�$���M�$�044���uG ڰ�O�A����i>]����.�=��~�}�1,�8[�`�cd���Hu���#gY�V�6�ֈ6�{��5
��N��kئ��V�O�Y��u��WpW�=&�&.2hu�$	F�g�)�C�f�hCah*%cnT����ӳ�
̜@���� ���S�-�|�Qx�f	�Y����I#U1��}����kc�Bt�� ���VW��7S����(�^��(�βZ��՘ϼC$��F:r���feg4$p�|��oS�=�	u��P'�`�q�c�>GQi{)�Ow9Pߵ�)l�V]p�oft�1�\\)��5S�"��oo'E��q@�ϗ��u9�G6����:��J~��a�\�� z:�i�xP��)�EFlÁ^á1t�1���}[�mp�Ȗ4Fq�m��q6
���1y%�nt_g��P�Z��^�.{6X��H�{H<�wp��N�e���,՛M�.�ە�:/T�;+�~VH�s�ަE��N>'��x���Pt����3]�i���d�2�'[	uv���*�2�ɯS
��҅F
�
M��:͸<7�jQ(^��[�l ��zŖs�����n���U%m&9+�T�3��&��(�����~����$渆��q�b��.v\n4�R
�7^az�u�l9�tΊ��f��x
� ��֫-�]�ss�������kX� ��@��Ⱥ��T�;nu.�����b�Kݘ�f�}ؐ������x:2���ϥ��ged�MJq����������r�����'�������Ց�׈�n���8S�2�D�4�$׺푌e?:Ǘ-{||ٳ��p/OJ���T����d�=uF�)�xi��~�3$S��͑�����R��Z2�r��P�=(W��a�U��҆2����=WqA�tj >��F�|ԫ������Ľ�aMrO�Ʊ[�q�D8�,,�Lmǥ_��鍸�e���{�ǻ�Z^����UQ��*����0�Q<K���dl�1da�o ���4�����}~�)5�X:v���`��	*(W�f������W-��9��f�{l���@��R�cʫ���{9�|�)�Vq�'D��P�Lw��+-�۸��҇�	��mz�my{�e�5��^r���Z���`�=)�"��p���*���D�va�"xC��,�y�2i�c)�"j�q3c+r��c���S�V5ay�2��;��R��8��8z����Y�Ѻ��v;Tժς8�!j���������&��1�Pw�� �hڠ�d^�&��|#M�����i3Ѿ(��gIX1����x�f�f��{:�#��U�\i/rÆ�7�=Q�嫯c�A}2c�wM/�fN���J�:�)���ވ���'Neέ�#2đ/o�U�Ef:�~��P++i�p0�(;��W���Fg��%��F����L�;#�}ō�N<���|֊��V�����P�f���ޖ��s�MT��%ԥ���z��q���T������T��͇ <Aֶ<n�4 #q��3Ԋ~~�Y�*u��a���N$1�_�!�n�u�1p�V�kN�\�C�UP<f��I�X�?pȭ�!���.��5a�a�:dױJ�%��u������HT�(�~�%@Z�Z���V�_;EnR���tmY�!���at�0��Ӟ�QP�#l�X�}ƣ�Ѽ]�����ݯ���q9���R��C��7�cGJka��^���ȃ����Yy�c|�^�����>
���t,1�����w�B�]��M�,]�,1o�"Z�Z_8������\���$.�^J��O���({H��5�/�"w��׏��e�|�)��o�I{kF�8�������2�����>�+�O1�ףZm?��!b_8�8�~��LV���v�T��yC��r��t�lmtt�u۹gt=�ϣ�aN�X�Hm�g{�.��RnG-�G���i��E�·�K�p���Ů��;;����I�Aǁ�3-����Uv*S	s8u>,�p�:U��3����z�V�gf���U���DU{�Ge�a��̸$Ҧª4P�ń�仪������8�Ce�`�W��vs|��׍��E���D��L6ʬ�~�q:$Ԡ��e���m�U���CY���C��]z������sD?��by���]�*/emg����[�}S�/����xzҩe�6��4�f�����
'��:˻��)"G����^��OX=e���P�[':�Ex��Lu��25�3���������bU�!�'o��kwcGUOd�w�b�ޚñGhՖ#��1eQ;3�d���
��a��W��9��`�Ǖ�e�=>�3��������-��Wf#�/^s�/ّ0��;c%�}�����!q=��g�n[:�\�E;<t���;��;�绳�Q��WS8,UCŋ��U�:�J�7nl0��X��*RSu;o�:B3��[{Kz��saT+������ԯ����<�	Kˉ銠ሪ/�] �#��tNTN�����;�
b��p�;�j�;4��<��{c�x�Y���U�F�,ʺ���ܮ$�3j`��.�|`q͉X�"9�݅�'Z��ύ��\��q�}&}�Z��f�����>���q����a'k.@(
yK{T��P;�d�����s�6.���4�x�N��Bı] ���3ԅ�L�Q.m'�q�J�v��Ƚ�l՞�^�{��\])`�4�����8_ym����p�ݥ[�7����9�t�8˗1}��I����.�Ш�s;SP@�����9J�M![ۈ9�Y�q���A��^l�B�p��Uza�����
��t��9�%���8j�ttJ�5�OU��ʛyEԹQh�>��U<
��Ŝd|�$�u�qU��T��ul݌����ϧxZ�OV����VPv{�h"���j�t',�x��h6x�����A���p�n���B�*F�H5�,�T*�H���i�\�@=w�l��+B�á�]>�UT4b��%��#< ��(���� ��P�\X�=���^�{J�8�#�z�F��m����X�#�����FF��I�sb�_M��� ��{g��3Lǋ՜��p��M~,�������nb�/�P�����пc��9��b��@6j1�#%��$�+K[�n°Pɾ�P�N�X���(�\]�s�eM	�0����[[����t��+[NmLt�S��P(�]�%��Y(1�=G�M[���5K����Q�]C)\�Eegf6��E������__��5x��%JS���.��ӟ����.&&�a@�<T�c6�V�ռs˶�u�J�ӹ�i��%�&DfA��*V���˸+���^5x���	�x{Wo��9J�w����N�x�����^���~:�X^!�b��~X��b�,U��/%B�����:�K/r�mEJ�;h_މk����QL���p���P���D�`�K|��W�%XzV����(�%��ֹx6����A��Aܾ��h�:xMB���*���,�#�:u3�ߩ�[X;ߔY�P��*�<.6�c,1iy���z�M�lJqЀ�y �89u�TT��K�w'���w� ���G�k�TK��YꞾ����ՑfɊz�.�����i�@jGIݳ�����!�
%˞o�X��
��,;���;�ݘ�3�+L<uQCk5�����z���u�w����^�����+(�hXD(>5�XB�3�V�텇�=@m��;w�t]����+��^"�q׍?�4ı�%�a�X�~�4�\,b:�CMR6�_�D��)�硯K�%jX�s�"{F�Zi���zC�	��h?���Y��ZHW����t�[�I/ۛ����U<g3~x�+>��_5��:�<:f%&���,Dm�물ǡ��c�+S�S�}�O^�&=��o���S���ٝ��S�sTZ۸�7�d��ҧng�@���E��������{5��Ŕ�W��B^OYJy�a�}��^5�Iu��5
a�b��a7�'D�u����E�0�df�s*��o�|�\V�ۗNP�sL��UC.J����F�Ce'U���� �ް���-y�~]<��$�֏T��_]�YQg.X�p2 `���uq7Ư��Z��Z֡�W��$*/�bH��E�	���:K�Ƭ�����z����%8��O@�f�e��է�mOds���X�=�^����LG\E�`��y�d
�PuI�q�����Ԯ����\UX����5�C�K�g�����K��lx�԰�t��q�3���jˡ�C�R���CE�Aܺ�-��npT�5Ü�GA�=o:]s��K�WwU���u�!����Q6�ܾ(1~��LYs�j�+B��P�ud���6���������T\�ȹ�^���0��h�AWOj��)�C,D�Em�f����չzr�T���f���������Z�M�}ZСC�������Ըȳ=���*��ovX��Sx�2�iq��KЧl�B�/�!O_�%�������ld��:�|�,�gK�3��{p#Q�Q=z��������\�;ʜȞ�'��un>v�����'�����Q*x��
R�AET��Y�.��zy�����QZ�s�(��vYb�@irs��1��W@�AS�	�,]�>��Wm�����uո��+��[+g�9�͍ڪ��,�.�߃D�0꫐�Mg��;G���/�9������&v��/��Ąi~�z=<ܳ+�tx,46T*��#�aC�r����<��$����i��6�)�lmZ: ����zX�sU�-4"��<�l��#T���/�3=�&�k�9��9^�2£{r�FC�g@&2-s�$ߓ��L�d�s��%t�#ݻ�^`ƭ}N;n�<BxW�DІ#��u
4[��U��D��$P�����=�oX*�w���9���U���WbQ/x"�l�U�+���U,��N6�w�u
N�T�G�H7s������R��pu���}�'�2*�l��v�0�u�Zv2c�7��-	���vJܡ���F�3�H1��4uT�Aog��c/�j�aٺ�I=�c��L�D��ӫ#n�2�ͬq�+�є8>\F%�����%gN݆B��dC��mF���Aa��O({��C{��p,h4ޑϿK��s�h=����Oח��$�x�<�u�+a��"MhRۣ& �.�|��zՂx]�R&k�\׫����+躥+�sJ�q��eR!��Q۽��;��*Cn9ѳ�Y|$N�;�ȫ�h�ŔN�ei�8%��Tp�Yp#����Q�W|=δt�F񺍡�m	��5�C>Ş�x�0{����1u).W���rud�D<s���^,b3��.B��
��ݝ�oǒ�b%*�k��3�ɋ��3�pR��vV]h�)u��d�D]�B,O�����FP�<�)�4�*L0�=�b�x�� _�zP�UH\��\qܖ�E�'�o��d魵��BDe���uȥ�V(Z(T��3�֦"���@���t'����V#|��M���x]9�6��gd7y&��c,�<ub���0^ɀ�D-%b�L1��s�[̬�A��)��׶�E�8�� ��a�l�m��sBb��3��X��N��4�&:s5��'�EjN�Aau��[巆o�<��K��J�u�Kɼ��}�:=�p�V{�T�m1���[���U���`��T�l�A{�A�����<�;6�t�&����lsU�P�ծ'� r�H��q�J`nj[Տu�ϳ���5��,��������������������',�Q4,n�WLo�9
�_J�(��#v���7uxz��RFl�9]���Z�y����`ۉ엗��k��&?�z2u��ߣ�O�8��-�q�t��4ǂ�Y�����y��{��s�Y�6<%a����t��+��rAh�s����3��D�ͫy�5
}͡,��$�������յ��4|�d����TlrԘ�P'�o�	�["��|1�^е�[�M8����4��e/�w_�]k��Cj�^.-�F�q����ռrâ�2�p̚[܋޾�s�}�_pG�'�U��Z�0nS���
�aИ�Ql�2���֙��W�«c�D����]ɵ�g�*�hq�łrX�Դ5<�BV  �Q;�(<�u����}[�i.��c������v+��l��N���ZP��<-J�l��0�LP)�M�]�%e������r��x�U��X�5�G\�Q��)7 �g"�Oi��+D�������k2��p<�X�C,P�<��WZa���V���鐠�1p��V-䋬������2�2�]2P�S��,bPՑ7���!O��<�Sļ�EO4��Ԕ(=�ק��5�fp���
�-�¹�=+�t&�]�)k�va�6�.o6�����j�HVQ ٵ�b�+��x:�7 t�6�����ny�`\��^�آ�<u�K�E�ճ�&�M���R�t'��xڙ��u3r���0[�ݛ�q��De:34��9�����y%	f탈�<W[��4]��C�.=�w���*��D�Ԗ]��WG9��f�;)L�)t�@s�������n+#�qW�Z���N��ջ�8��Yg����#���F�x�@���o.N��_-<孖%d�31ͧs4L��g�*q�cHP��i�� ����t&�s�gE�{2��I��6>)n$���=�U�kd;��J��ݤl���fMkCţ1�׸�nZL��u�L����*Rb��3o(��0}�J�<ѷ"���� x}��C���z�\�;�8���L��84��9m��%l(p͛Ř{;�i�M���F�#�^�.<�!�{�j`�zr��C��v�k�-��e>��|�[N�
�/�R�V7��ƭ"5Vޔo;���h�J�{���&yIPoRV�@f�%˧bW[�Ɍ0�+�G���5;�=Ҥ������|ie�:8�O[�X!z�ɇs���CKl�p<��=RԂ��d�.��L=��T��X��έ�ݸ�˛o߸]
�l��q�m�s��r�Y�yv�h�(�c����Hd={�>L$��НP�T���2<vj!yt�Lmf:�vO9���^�'�ҧ�^���nZ�xUi���G�0ؗ������NF/�˙�(`�i�fb�B�:�U��!W<���V����Z����|{��_C�z����<;),W뻦���AG}A��W�o����Ӱ����Z�x�u)��͠�G%��bIW[�ϲ�x��j�(�-7AJ�+�\0Q��4�d֍���l��;oUb(�� �CW[ �<�;ie_j���#�X�p��7G��p�1qm$�7C��ؘ�&�W1ӭ��|�u�9z�95�÷��i�5����!.0wo$��S$��i�c8Q�n�ǁw;cL�;F�Qg{O.��������H2c��g�Y%wF��rbיLZAtr��1�t6�d��/1����4�W��`T�j �����������9�7׻�F�W��q.���'3f�U0l΃6�H�ݲ�Ld��fA�c�gej��X�	�+o^�%�E�h�Jd�>U+�԰��ћ�L|9X>�e��ߛpǮ�.s[|��f��P���]\���Z�f���&J2�9�C������jT�|�+]��I�60T�ܗ�[�󞑶���d\�<]�;4�(�_9��m4�� 1�A���#*�
�u�dדiupJC���w6��|�R\˝���V�u����̿}s�o��n��<���S[�ۥV.�48�*!o��DQJ�E]rD�e���fٚ�41eY���_ZE��uz0`�o����j�
	%����*Z�*�����B����I���)h����Jh�*�(�������&"a��*	�!������������((�����%���&*"��(��"�(����h��
j�"	*
���i�*�����"�(��������)*�������Jb���h� �
�*�� ���(&i���(����"�((j���&����*�%���)��"��)"�����)�"Z*����*h*��H��jI���)�"������$�

J�h"�&��*���j"�*�&*J������>��*����K/���Z^���KB?!���+�~��A4z�[��pyщc)����T�HM6l+��5��������EjK���E��hϼT� Adq�B�]���WU�a�^w���㨺7Jz̺9׻=cwR��GEn`!��5�R�(D���B�<>߲�-)�������D��o���7sַ����Ž"޶ֵ�<�F���b���K<&�E9�v&a��l��c�u��>��\L�S]�����ݜ3���^W,D��R�Ӧj���X�R��E9�7��8��B�v���V��G���:X�Tˀ���6t Q�7�'^�����ӊ�ҲyC䳕v�����/֫8���S;䪌�dS�+�qd�^uD�ʐ�Oh���t�ͽ�0�9��
�'hs��÷��;����P�ѫ���^Og�E�.8�s���W:!�
2�)��� ���
�!o�����o�����>�O�ef,�u1��v*B��#�K]l��L�r��>���a鈑��ȯG=���K�M���,f׏��a�'�כ��2�d�b&�-&7z�IpM7W��KT�F�ѷ��2�Gy��*�O�z%[]Cؽ4_������|�7M�}ݻ��.�o!Pm��Ѓ��VF&k�п����t;Y]�!���Y�E���z�pbYa1G�+雔� G`������;�P>*�KL�A}��^�J������&���'p�ګ�.Q�7����5�c�T����pq>}~6�sD_�K�U��.5NH��َ�lxإ�J�k��'��{U+�p<^t�kT��-��ֈ��U�{[��qL.)s<p�^㋱����U���u�9�N��W�`�V*D�)CDK1P��cOa�Z��Ev��8��[�s���Y��b��2�U�p{+n�p�	\&��5�(+�����S��I̸��Q=�q޸�B���C&�O8}A@t/WVC��7�g��]e�<+m�D�lg0�e��H.��z�y�7�3V�ю����L�ߦ-�T<0���
X�����=DW1T�C���Y�Pi�~ScB޻�y)aY��=�P�҃����q��3lT��x��ZB����(�~Ӛn�θ;�Uxm�(l�v�EE�'lM�")<=���]�Y�zޅ�$7�3-��^z)N� (����U��|'�M�	\|0"��x*a󩐭hz������z�r��(��hb	՗�,�k�B��晽"LOs�$׹8�w�Ud
����;�/n�����i�8��E-%��V�:doVѣ�K�q:U�+j�B�ǳxF���x8�Kɹ�{�n֞�a}�ڻ�H�(({³�(��a�C}��"�����yQO.��]�Y9�
�(o�U	t3�M��QT{[6m"���k���i�Y��wx�z%�a]{�x�^�wf��v�����v��IN���Ch!]�k!�x��ڨW��b����Y��#L*o�UrGz�$V�ĸ�����I�>�^6O���뤪Ybq�<_�}Yi�Q��f�1�j�_+APACN�Z�o��	�����o�Vz�A�x�9GD]���soeBNET�7��<�#Q~�Uc�g��f�PA�.�f�1��.��B���Y+}��ٲ�W�xV�}R���Eu���'K��:��+�pͨb�����{�M��/�n=��	�;�W	;2s<�o�Ӄ�V�1n:��:-x�d~I��Wt-�N=Ǹ�b-څ�����{{w\r�z������.�Z<�Դ9�m����r9�bzF��R�̽�J��Ot���e�57��Aa�vġ]�|�1u�����O'�V*����t\�V7���۞6�� u�ay�q�LR� w���LZ�T,\n�n]Ccn���'6�кҤ�B��]�Nh�5�+9.��ʸ�6|�/��նPO��e�ѿ12�m�4ov��җ]�\A��v-�R�DE�%s<����b�k�p���~������|��c���
����.sj�����5�O�°[�,�=4�Aro.��[Y.ҵ��������4��f�5y&��Le��sBb��3�`p
�1(o��m֖Z�պ���.A�
�Ä����c]psfNO�8�P�&l��n��B�V*1�M^VW�{�^�S�ix�|+Ru���Zi��v��ݠͧ0��C��B�rZ�z�ui��FZ�ځ۲4�8R��A�	C�N>�h"�娱c��F��V��gv�\�M�^ESA�W�I�Yݲh�g����҉�)�W�b2ߍ�(�������]�y�_�K�T}�W輣�������4$\(2W�u��8}� "���ۙ�L5ɭ�2J͐�TÖrZ����UѪO%��������
{N�}J�N���*D�P��Y��YSZi�"v��Y�3�3q���n���:P���~á9j�ƅ�w��}t�)�9ͻ�>�Ͼ��X��*������������-a�6X�+��Xkl=���ɭ'/y���{�ɑU>y���b�krjvt[Ȫ�B�ˀ�e�0hK<�~oJw���b��Ŝ�o}n��4A�rhoW�fcb�譳r�h�c��X�c����l,@���}��VG�ʴD�#��Z�Ϊ�)<�Vw\F�B6��\��YS#���Za���л�Xع�&���:�� �8ul&�^�Z,���>c0����WF�\�U`_zS���{%g�e�W����<O�Zճ��B��,�
��%˩����(7É�5���;��x9H�8�I��cb�cJV��@��K�{c���Un����A�[�Jͳ��,XzPj_Zd��V@<:M{�
J�J5r��ӗ�� %�����p�P�T��.x�67��N�cV����!��M�4����Q�Y�ef�\�m��8z�A|u`����k�^�+��٪�{fL�A�|ŴK�Ӟ��6��9\�,�<�M0EF�L8N˞o�P��x!Q�,;����ΩCc|z���ɳ��l��jۯ}�� ��u��{�}�Ik�B�)�h�)�W	���ꊪ;nOٜ�zQ]o�`�q�}���{�e	]�*���LTı�%�nR�^\j��X�C�s�.�����^�q7!g"0�U�82�4���ŀ�K&��T;�d��w�^���Cм`ͽ9=�;���ڮN��1�bQ�"K��da�c\�a7��~c�?��Q �6;j���GkX^��K׫
����z�̒�v�96�����/)���T�5��E���o^:D�j�C�P�N^c���(m���ar�w�7۪�ᚎe(�8�p.���v���˳U�������R��Y���g{�:�>5�1�m�#�zo`���r�뤶�Jv���<k"U�͝���c=�N(��3�	�ϒ��69Ox�w����d����Y��=>Ϫ���7���mx��T�R�YS��FYu�~�<�����p��ؗ����F��~�FTjD�c�*�a�W�g�k>���o[�gT��ŀ:��cӍ��^�p�~�"�^>�+o���&>���j�J���q���oK����$��w҂&�zPf���EC�;#],(>s�i[�n�Xb�f<o�W�N���j�ٞ�T�C����M�|��8v�Z���؋�1��D��҃N�I5���|��T�j8v�R����]�E>8�<P��Gc%C�%��C�V�D=��c��2Ls��l}��z�\n��z��K��Dq�*qb|�i�>V2
T��AVh��U�a���9�W5��T�Rȁ1Ĭ(g�/Pg�E�Ap��X�ѭ���G$�n��[���e�{���{�[�yG 0������0�h��PT��B,T"����;D��x����B�j�(_%��X� �%��-c�+kj-*kX���}��3�WN�I�ź�{	�R�{�

�l���qY/&05�r�W1c�IQ�k�/M��T:[����}&1̺��]��d�=��\;���)��;B[��{���<G�5t�R����ʏ�������l�23�S��UP�s�l�z�\5��G8�vP�f��ʧ��W��e!uó�=��-�(:��,n��c�B����_X�xR'�9��9W�j�2����
��H�,H�o1X���l>���ݭ��$�S�&��Wci�cj�� D�{��q�)V���S�)0If���B���3������[�oLXcҒ�u�y�'�0�kwʉ7[ާ^������O �}~�y��nЊ�}KG��v_��A1]d6�k�
������/#�	pH��ݳb�C.�U.�r�#v�`����G4�4В�|/���뤪Y	�ÞS�k��SZ<TT����\��{����팟066B~��(X�cݺχz�[�N�8�|Uab�pI�[P����	.��=&Ls2�!@�nK�J.�f�F{�7�r�o<�([�}��X���k�y��fU�tz�Yb:����ˁy��*�ï5�.5��ns^q��<�-�x�R���u���hCo׈�e�ؿ8����2��do�Q�0��=6=�괙�|�b��d!��c�k��j��9	q��Z�\������H�fr��h�un�Ab��ɨ~:��u�#VNthj[gA7�(l�9��g|-8��rnzY:��[���K}|��yN�g�=�����\��cn\W�@��\�aA�2�S�h�|��V�˳�}+o��R���f8W/:ظ=�&.�Z8O%����y�����^^�퇘tD�sLO�Ny��H�R���X���p6zP6���e�7:�p鸳f�~��E����R���#�N��c!)�*��:�a#`Ga��w8��]A5ȫ�S@�%#Vꐹ�X�S�n:���w�i�2�<ub��`߷;vk��M����wQ008�Hcl�Pwc����&�;6��A�4b�W}f���n�'7�$7,�O6|�¨TYҵ�>�*$�J�C�0�/��z�g��]=+�A�7Ӛ^�h�^q�7ủ���{�91rߍ<�~��&J��I���J6��QK�^^ٺ���Y�@ǘ�`����/}�uԗ����tK9O�,Y��;�)���=��Y�}B�l+z�A�3< ���5$�禡�#&�X���P��s�V�to�ɭ�v:ʍ;Ft���.��{q��L�e� z�Va*ͷB�']\͒����ˤ��\w�n��7�a��Ƴ!�ލV2:�;�־.��O����41�����#c����J2K����,��܇Q��Lm���k�e,+Qۙ]1�Օ��T��h!�t�����23Æ�>�&� w�	��p�T5i&or��ɫ�:�HqХZ�|�"y�clcc�<��7�,��(a�t�i���1�!�[ZQ�����������|
�}�l���9��b/R+5���ɇ,O/0���o��j�x��:毑�:2�%�#*5��5;:-�葱j'�E�p*3e�1���q<;���T^�_��W;�g�iW�u��ᎴxR��G�7����:���"Ӵ�y��K̊�ĎŢW�_���EO^���Ȁ�"����3�Ϫ8�%+_1�-ݱ�ꭻ�mV���R���=��Pe� �/�����{�@C�r�P����O;۽�#A�C(>�:�ϒ���8��5ajȊ{�h砷\)*����){�����e-}z�xD*����Q< ������XՐ��5�^<"��G�c<���M�ϟ/B����k��OD�5�s��B((g�����Ck�;�d��-͚���h+œ�t�+rKD[٬X��C�#Hk�c���;8����]&$��\5I�G�,z��C��CՙKan�H������5�b�G�J��$��V5��2�ƩJ�gy��}�]���>��[�1��O��V��y�O�xTU���Kp�Ix���[�^j�q��x���W%��B���(�3%��fVx�@W�ՉOg��
%���o�^���7��P.:�*
bz
�c��y�ھm���)���w{�_�dH�r� �\X�v!U8��p0��b	�x��K=�Z����|��k6����?L�٪sj���1(�nɢ����)�V�	#ip5�.ao$��d�b��.hh����7���N��񩗙^L�=R]��V�-�f[܈�|Sz�r��W��ۃb��<�"�X�%H����7��:r��Yc�6i��8!�^�.�򤞧��1�}Ҙܑ�P�fڟo�#�"<o� ޝ,fy�eJ��fmZ29�̗-ho��8���:��r����r��;��e�Y����+<iN>�Aǅ����ޮp\evY��p��$�mx�X�xG�T�.�e����r-	Ѷ�
�B{�+�~RV��nkx�7p�Q5�,c�v��u�04�pQ�֊�U7���o)e����N�6Q[��:AQ���u=��+�M.s��V�Pe^�1ٜir�1s���'^���\�ٖ]䷶i�%/��g�b;`e0el�Y��ǻ�}5kҨ�4moa�ը�����=���܈���*��U�Giwz���X�bS�i��,�[��>~*N8h�7�a�Mz�kٳN�3�Α�;8��c������}Ή�.�V�ә˻3`�"R���a��4��$���Uk�G�,v�r=(e�c��6:�2�H��+`��֭)w��:)�#�O�.oT�dÛ�ܶm4V8�ӑ�V�<�{1I�k&c���.,��V�4���c���]�Hv�{>�I��|1�XkD<���G}���ӑ����e��t�]j�~�⃬� �?%����i�^Ӕs�%C%6�2����,�Xp��%c{ެ� �"����>��}E7@npH���`���!b#���;uN��;��w�������v����f�N�K(�e7��r���Z�d��a��j�;��wW�ķ+�؅�9+`�@m��p����n�S[�+��/@��i�yw�AΟe������.>�y	��a�4��s-�꩗*[T��h�|���Z���jl��Ch9�1-wԺ���)=�ظl��q�P�Pf�ͫG�4�=��MQ��	8�oe����#�'&��u�P%�Z�Ug�-"���yK/��w�P�ϪR�7եv�Rhم�=�gR�H��w,v!��״[9��O�O.�	�������ʠ�%\
GG#ìgym�x]]M�kk�Q����b�P�{]XҼ�љ��D�����m;7_���bxnf�-�}ܧ��[z �#�c<�������ٕ�*�<�et�^�QݞB
�Ģ�g��<`GZ�dx��](ۀ1�սu+���K�6�]�e��zrn�*����x�żh�H�o|�'�}�#�<�؄��r��$���T��|k��Z�֟�T�3.�`�*���V�D:��	��s��&E�P��Y{�
��;�U�d�"䓒�"m��}�p���sAW��+��K�Bѥ��VA��ѥ�Hc����#y�ܐR;���iB����ChW4�R
U�Zƴus��!u���F����Ά+Gb³l,,Tjem
[e8O��QZb�dm]��tQ̤�
XP�򬫚�T�:�������[��:Ba����-&3We�ϲ�Is)�v�	��*�oMyP��l�SZ�w��͐5%<�Y�f7Xt�Bd�;��1�Ɠv���Ln����T���n�:�b�������pH����%)���K9��� � �ː}qѕ�jm��Vӌ�L�3pl;�Y�jH갰ͥM�"�́��#�J��%%A�B�4T��h*X�� I:U�7������"Z��
��"s)�H�(�&*hb���)h*���*����"b(&�!�
F������*f�"ei�'&�����((i����iJ�� &����������h��bJ
��R����((��"J�"
�R�ZF�bhJ��
�����((")�
�q�"�$)�i���
i��
B"*�)"�
(	�)"\�Ȫ���
Z
h��&�)JhJ)���� ������
)()h���(�%&"I�J����V�"h)("JJJ��K1$����(i �� ���B� «]N��]�lv�����s�<Jl��K7�i^C�����o���Yx=�xxO��0pI:��v+lù�IoŅDK�|qu��,f;��ˠ@�v+�e�gei�"2�u�\�p�w�cc~��x��"}N&8PL��V��Ew, �yW+a3q�uP�+�]]�Ku��h�农.�&��G���x\d�d��+����x���_�y��8�%�y��w��ޑ��&c!ܛ��b%߇Tt�Zy�c�T�WV�C�	U���z����˶�P�<��4-/a�>���>1��n����|������C�XRX�snn*��o�N�us�7���+	�pj�ib�}��a�]o�t`a���&ye%{]�7���R�F-���$"��=�:φ��ݩ��� �b�X�����祋��
��N��9���������E����W	�kWV��u��w�Q"���-�ޖ1�V�.�Ff�_[}���"O�MR(�,{R�m��E�L��ds�ţKwΉ=b*J�K�%�7n��Alt'�={<�tI�J*���&+��m����=֟���Mnɻ|e�,��^���'�/ID��&}zO20�;В&�X���VL��	��ߋ�Wh�r����8 �]�)m�n�4.R/7�1�&fG]8Q�n���`Y�tE^#�{�\��G�j��M���0�yi��F��\,b��������r�nnqs�aX�U��:��v�L�8���[M�=J����؃��������u&c^��٦K�׆j9�Wf,"kUfBf��4ܔ�C���������+p�G:�/B�λ�wG�~�6=k��+�/z��2�Fe���A�١��tcSb�Q�*��Nhc�[z�u��uR/�K��4��U��:��ּ�f:�������v0+~����/
<r鯺v����o>uW��А5�g�����=KD��-wy�a\��Ϊ6F��1�N��s��լiR���ѭ�p�.p�ɋ�Ih�<��P-Ӧ�~�&�kM{|�a���5���^ƪ3�Y}�q�r
�&Bı\�)��N}̉�}s_S˙%Z�>n7�/)��x1S�C�����{f�\%�1��H�{��ř/���αN�x�H�*k|"�<|.��t�'1�m�Iz���X��#^݈��7a�b#���~��0��@�6��Xwc����$;ٴ�� ɛ0b֤�d����x\X�lQ������P���MlMP�/sSS�����c�6�7���驌ʃ]*�^�7�������̇3�)�ʴ{â���YU�vQ᳴儺�W|�a�Grt��d�״�u��� פ��&�&���4K�qd���f�#ܾ��v���e��<V�Q��p-ID|��i?(h�[jdl�7����n�p"���Y��o]UD�b�c�5W�zj:�+΅S�^�JKA��-E�-�o^^�`�&E�cۊ����g��*qp���� �Rɯ*f�Ez]�g�i����e(�?JqE*"��}Z`�@��N`�E��s��s���� �=7L6�W^v����o;a���E�^�ߝd�LS5��p`�ⷨ�]��U=WZ-�r����^O\ommbU��P���>���,e>"<��8�������۵2���S�@%��;��ߦ�H���=�<��k=U:�:qxY4=5�'���/���?͡c���{��5�_��ѱބ�\C��Y��Rc�}��_���f�ϭ��!��hs�����c�pY���'�/�
#2ts(���p��+����,���9��N��~XS"flBD�{=���\�
��R�w��&�:b¸W\�V�H����j)�Q�	�/q�Z��Jη���*!8x+B�їڸ�ͅѩL9�Q�HG�L���+���
�%kH�5d	;ޱ摔/\��=��
sQf�^�s�ͨ{�i��.\��O��G~�wΌ����um�$��q�7����N�hnL���ۖ�;ϳ)ɼyN�h�H}S�(�+�7�P����. ����ç���aI�-괶�%�1M�[u�(�g�
�E|���D>~T9J䡟��޹cV5dD�޼ELe��k����k�4��t 1P� #�'��$B���>\��;��+k�˭ ���ڢyr&�Í�E&S��x8z'�,�P��
��Xz�1S����8[oA�+:�E�{1O]�P�W.�E��B%1�z'�,�2�
�{2��!�i�Tm凢4�h��~6 �5ե>r��>��W����("�UlK���,8=�0#Anw7Zt�S�&�-��4�9���c�S.`���X�DJ�NZn��t�pV����E�_ ki:r]9�5{x�\nLR7D��� ��zl�=�W]�Z�'�����Nw�����v ������q;��S��C�ucP_��/$k�U��!�x^��\r4��_A�t��#�;0�)ZD͌��CFK�2̸>+�$��,�t{3Eb�b͓D��5���+��D{�����L%�Ϳ���GE�]-+���مuF#�Cw�Q�6J��
���'s��>������� �s�z5f)M��&Qh�-��ܲ�7}�=�Oei\��n����nF�}VUٍ�z܇�]"���LkvÆ���YO�:F
L��a��a�]Þ��Z��vrUfJ�é8���w������:����t��ܜU<"�p��V_J�f��P�;����ݺb�*T
�f��ޖ�w�)�S���,o9Zj�ئ7(��YS~<�Z�uL��tD�Cխ�7J4�<�q�7j�7ŋwn�eN���%h,�=c2m�5K/��iou�B�V�aܪ)i����WK�p!��(s�#�1��Ǒ�H�ng_`���R�;=wZ=��R�-ǪC(TK�Qr�x�`�8Щŉa_Q�f9�3:���~�N;̯%/oVE�)P���KD���Q*<0�	A��T����[���x�u�'�ef=�#Bu.˷0�Қʑя���ã.M�0���T��es���ŝ��P�f#'��hG�WZ�c\x{#vtȫߦ8m�g��z"a��g�� *���m�Y5k�"^V~.X�X��:X�9���pnf��X��9�P9�bH,��9׻3І��6M�Ga�w4Z�!�v��M�P����Z�4c��nT�w,�6��q��x�V��`ޙgAmSeK����׶��	�ϙW��y2���H���}�59�vZy�_w��\���pX��?p�ݔn�RW�
�Vh�w��C��YT|z�e4�U��h��uw�i�`��2�m���Kx^>�ѽ5��j:퉨��<%0z%�ۦ�j.e������|Dõy�9�J�%�n�R�����PIp�EC�"� Zq:$Ԡ��Xi�%QBku
4��+j�b�Y�_LZ�v�]�E87�$�`�u��stx�eWZ#���z��=uIT�U���+���a�8�¡8t;sh���Q��5H�5�5���y[�9�@3�܊�
\�ս/�VH��	x�	��\Q�fٌ%�xd(��7�4;�twƄ�Z{�{�h�K�Ž�)��3!��m805ٲ�Cϡ�F��P�\
͔�R��
΀���U�+8�\��E�����.��Oaҁ����Z��C���)��(�}����F�^ڽ���%��B9u�~��F�mTc����}�
a�-L]O����hs��q���|ek/�%�Y��ӞFu�x���]6�f�Ø�+�ܩ���Wo�5�bLM�F��*쫭��j�ʼg7�5�q���|R�1�����<K�s=؝\�ļȧ|�v*84�]�R�|	EӸ@�L�|t9���#Ӕ�A��V|���7/[B���19S�_��Vۺ�1��v�o�7ځ�΂�$�c���BZ=�u-�l�=W/������q�.���uxXq*w��%�!��%
p1l�����AQ�'%��T�Ĺ���:��d����hL�ج�P�S����)l��t�����SŊT*˝�@�w��H\OM��R��z��j�VL�t�Y�(�yl�,�$U��/Z6�c�lC\�0��h���QJyW!���3�^t�+wT9����X7��7��b�wh��뾳�X���L�0$�0�KjPF��G����1'�8��ZW�;:�Ou�[��u��&��ֈ6�2��j�bEC�4X�(7���"�Y爵�쮅u��@Vڣ�-Jh>�Z��J������"�K�ev�%��:���>�`̿ l�|��{��S�V���t��ulذ�3�Q��@0����� ��s�D���uwg	~��鞚��rt�/P��x5[����&1k�Y����dǱ����Z�%9;�)-���j�!.:�v�A[��,��W��xU�]Cp�./�cI�PHQ���[G�+�هi��9u�[���-���g&�ɚ׭��wsF��rw+g��b�"���Y@*>ި/o�s�U��`O�em�[��ZϏe�<�ʴ��:���k��_`��z<d�:��±wiz&г'�c�l�Ο99�qÃ��+��w
��t�g�#�k�=��~~:r�(nm	ьoD��
㺉�K����Fq�.�K�+��&+_��6�U�c|����h7�ո��l�gӰ���yC� *=�G0m\���q�a_M�5Q�s���\,>�3�;GY����y!����ؾ[�M��Ȯ"Wd�ɨ�S���'i�p�=e�2OS
��:�1���j����voJ(Q�#ԬdX/�q��(�5�g��X�~{(;�փ_WQ�p����Ɯ{9(�/�`p�l�@�6�)����(xE~Lg��6��|��5k��/x�<����֩7���r���\Dk�
�@�T���8Bk��l��6X����MͿz�R�@&�6p��i�ɊZ�.�ùVic4��X�C�<Ig���P��9h�{|/.6�9�O?0z��3]���f�z���m�5�'S,S�,����8f4R� ���ƏN�a��p!L���O<k�P���3��A�K��u�'\P;��;�̡(d����m�f.8Dx��FW F��KQg��w[�XGf��U��u���ٍ��b�c2d XN���OY�y��������Kp&O<aU���&M��)��Z�k����Y JnD��k��g�ѽ��cw.2�c2GXY�H�Q������^�۵Vv7&�.nJ�%}��9�3���,�7��-K���-�4 I�/X�w��G)��~��rD�>tn��iFb���?*��fZ�� '�W��(À��_�*�}���->���\V�,�u�J�[C�V�����Gk���x�Q0���*6���5e�vgWp��#�-����,a�`{�hz��굃�(-�%[��/�uV�ӎ�η�{S��}�,#��y�>��yث�cW��60e�q$e{P�&��z��/���^V�+{��g���b�<��
���� �`	��z�\n{[��v#����e9Z��s��]uM��oIy���:����9x3j#�Xey�����Lvz5�C�K�K� �m�o�/7qͧ���B��f�.n��=F�و�N��D����E���cgeb��'2b�S�S�V��[��ޞ�7����F�Cu��+��p�u{"k���]F����9��w_>D`����Oi�\�
�%�:%���\
��i"�=�H�Z�D��k=M�a+[�.�Vt��)i�\;�	���اGGr���ɥiE�m�պJ~S�f^g�����Ҳ#.伀�w!��>�4���,�x?.�w;~<C�-ĺ뵮d��x.R�����1Qe��/0�a)���z�f�A�V�w��d��0a�i�6Z�Ί�pyf˖"]�uGI���c&
�1Ύ7%���������E�ҋ"ơ�R쫅0�ұ������ã_�K�^�鄴O@Q}�����xE�>���ۑD�zx]��P�����3�����T�sY�]|2���<+��`3p����ӥ��%��~Lc&���ɕ��O���k8|/�{:`����2`d�`���t��l�
��Att!^Nc�#�+g�����y�*�����0���{���}H��_�U���ރ��p��#�Tm51AN�rP�*�)�e�.�NP'L�Lyc�s���^�t��=Y^���T.xV�L
���~6Q�D��XܠF�]īNdMK��5���H8̚��@.j�"|���Q	�h<��$�RA�X��9��w0^؜0-���,+Dm
��p�#^͚/g/�Xڗb��qN��7�����5���w}�d������Bgx���n�֯���i��n���B�vj�FC��DQUTjUѨ��p�v��A�\��((h�m�(�3o��wģ�J�,�u���p�n���cc̝/���VgP��Q�Ur���@]sAؔ8��S0�R_�y�v{�e�R�v�RDo>H�_��s+��R*PJ�u�!ӈ��	�9�q�Y/�5b�����c/2�ԕe�X�jR�w
"��/�#	����^P���V����m���;t�Ǝ�m���ɝ�9�w�F���
WQU�
Ιe����N��h /��S�MbN�w͑3;h���� �n�nT�yG�>�EF�lJ�:
����s��A�s� ��Z��֑�������)�y��ʕ%04I��66���-c���Z�$������<��s=4���*Q��ṎXgלK�l�ԬT��VtM �$Uݛ[[�@��5M�w�����
��޸�9���5:�������Eև�q���#�h�9T�ܺ��%3m>�K6f��w����5�t5��a �V���K{6Щ7����Qݺúص�*d��s���n��ӹeC��g�!�۽�X)}ͷ�-<su���uAˠ��=È�}����7�57wK�����4��r�J�`��Ǒ���n�-�P6I 2h+$�a����b���;�N�=}CH�d%�q-��W����}���]W����Z�������)_-5*�{ ���Q���Y�n՚A��qJfX֔��ѯVZ#��ke^+�]�(�;-�iohFg�lf22�:�M�'[˻���S��M7O���/�&�Z%��ۚ�itg��9��mGw��NK4Ѫ��eՠT*�+�k(��+��v�Q^�c5�c�\W�i��z�25�<����5	�\�E����,F��3�U��X��j��l�(�9:Y�����U��%�z�٘�u�g�Oz>&�6�v��x�.}���,����U���}ǵ�+�����)�A�c@Әw���{ī�JAJ�tcӨ���4qG��wM��>�S�M��|�ݢ�����<�����{�O)F��J�t�u0����yN�:��_���d���cY6TĎ<���>:��VDv��͢�P/}.dBͧ۸�M �P�WC-�'S1�T��WH�_wI�>D��ATt�:�+/��yH�kc�4#�����-� �Y�i��r�b�X{�ȯ]�i!�p�o}c�q� ׳A��V�a�n���ED��&�H4�W�E��t�)�L�8���`���{R��e���<�)�i�����3	ǒ��p�f�˼�f��k.� � ��dWVĂcq-w��H����sZ�ݞ5���TK�x.G��ן��,�p�H��L�g*6��㥂�С�Ovd!f,���;w_T���D3
�B�i��U)S��b�!-��H��th��ò�(ǁ�*�`ʸI5��]X�  �r�}���>���(

JZ
F�
�hF�����$"R��J�$��i))i)()"*�JH���*�
R�%hP��ꬢF�"���@�
JJ)*$*!���D�
)P�JbbhJ��Z(V�()ihZ���J�J��(���h
�i�"P�ZiJV����V�(3 �V�%�h)�)B�j��)(�&� (Z�h,�)rB���!()����Dr�|t��hE����>�x&�q(��칫u&���hV�[���˗�����nx���&܌��d�w9��y��Oy[67�s5����9�0���9�����7�޻t�\�:�i%C,�o��R�[���7��b-Nϭ��=N�:��V��w�=�:�X}+�M��n���Y4�E���p�J�|04R8��WE;8t\$&��2.	��z�ONxm2�ˆ�;h0"׮�x��ۛ�aQ+0����b����6�xS�q��F>�~FA[j�����9���m��R��=+A£�/#] ����s�i��I���,V���ʹ1)��q���'ȪeR�6\�.O
�,=�R�y���g���a=]pk�gG�n{�N��q��W�����E/T���_7�Z����4�?:���G���퇦�Z�3�.�ۚ!�0^ɀ�-HGl�P��⹈ls����Ľ��a�E-���v���)�>Z�P�Ѿj�y�b�~p�<�Mx�RQzЇZk�½��yO6�o�8��23`�S93����;�5Y���P�X��L����%��iOxt���9F;�[�Y�3z̈�tϵ���Xb[��tQ��Mff�]59!ɉ�G�w�^ݝQ�:�����G�yȱ�<NV�^�5[Ń�_{DT	��{�f�d�����&7��t.6�q����MᏠ�epq7s��[d-)�m�%Bӏd��c�^�æ�X����@>��j8�m��������J�2�O�=�6��>�3,�C4�S�5�L�%��2ToP��3< ���	s���B����=���Ap���hɮ������m�����{�~;��Vf��֨^.�	�k!`[�7��H2{c��p��*��U���A���ϲ��.�βү��P;�q���[��l��z�2wN��L�6����cF�=`+�����eN��tƌ�ڀ8�؎nj��S����x$.��m����x�ݸ�k�^��Y>�NK	� k|�=
�+\�j�{`K��� b3ǉ�W(2��o9�}7�Gu�E��pX�DRG̽���4x�mӛ�������hU���%aa���1aZ��uv0�$z�2K�����|mV�*M�Uo!s	�
��j��u�pxlEҤJ�m��9b���/k��qg5m������3��i�D��F��,��Fi�G_�W��T�:��o�dHઅ�c{v�{r���-aڕ�)G�ݨ�Xd��O���a��	��sR�<�v����!�Gjm'�E�E�U���nml ]�T�sJ����|�~�h찻�$u����,q'���e�j��㐺޿eifM��q���]�O"���ڝ9]{)�\�u��;�i�7�]�h`>��$��ƺ��Ӿ�[�[sOA<�SO*!;���b+�ٲb��T]w*�,f�#_��{�.xa�(E�W
6�u�
���͛u�R��uS�:ɇ��(*.�C�P�^8x'I�ݪ7/���-���W^� ��5������c�ne�`��x+�*Q����������{�p��͜MA���P�r�&�\i޸X����x����0#~�+�Va��n�1[v��+�X֭�<�6�}�LU��ŏ��t�K��\]���ٮ�0J
08-tH���yZs�i$P�{-Y/���_�u�K��<'ը7��-���o�s�x��-��K+�1O,F�^�+�Y]f������C,��q82���D�;0�B����leGe!�#i���*�YCU㭤���q��j@�3�8=�juq8�%Q�tq�"����n��v���W�gbͽk���jp?eJ��Xq�8���:�܍�s�T�lE��Ŋ+W��Υ��r�3!�����b^�%#�!��J3���H�ݒ��@�ޫ:j[��D �E��7� 	38�sM��n�-��u${	����9B/����v�,�9�n59Cx��5PW�%C��%������v������L�e�{\f3�>P��n�f�仱7rs������Tj�FeP�E|�^�mz��\<M���%q��7���0(��.��u������]�F�j㞭�aq���b�4������x�ʉ=���?8}�e=��96ݵ���´zw�x*��c�>~�����>�����T�P��u{"kl���)�.�F�mr�n���R�As��+B�"��e��*>Z6�Z<�$+FKd�@yg��k�v�����;S^�,+����N2b��᮵�`��/���d��EV��7�N}��H��b���\&I-��?R�a�솶�TF6�m���&���ױ�c��vmR�v�y��C	Xu�þ����l8%k�co�_t��e!u2ы%V�[9�'��#�E�uW*��[���P���D�<�MG���C�Z=�y�f�X�o;���%�k�K˖�e��ǇT*�^4G��ץ5����+
ϧ�9�x@���[J����g'�m���w��8ݪcD�WlJ�2P�ō�&��z/r��+[�{�9�^*`��NOEěPq�S�@����!]�\�a3t��:�/�!��{{�;t]�!l'���`z����d�-sj��<��n1o�w\YS��Iۚ^הX��!�rm\�}�6R(��G�ڙDM=u{H�9A�R��ʜ�n�ۉs�ی�"LM�;�M�q0����tI�Jd�'��]"hB��g�w��GJ��0�F�{�kG��Ai�^�K��H0�������F�&�D����g��} %ۜ���"���÷6��rh(��8��@:����K��cc���ݮ�=&7�c�j>�<= ��$,	i����'�\�����(u�l��B��]N��3i��رUb���{�;��=�cGT���6_�Շ֝��n�/�mC߄�<l�V��.��,����Mވ�ܝ���;ޤ՝����il_�l�D����TB�f�"���0Bi�Ϫm�b�{�����u��g�HM锵1u��O;w����Loy��ԁ
�)QS8�3:��¥%7��Әb3�(Wq��h��WcȎ(=nٵ��3������On�X�S���� 9s�������9J��w�!�/��Z��{��lM�pOi�]P��¼�^��#"����ѩ����0��wme�ZOkb��[$����'�˻���m�ϡʘ������{�v-�����$�ݤ�S�%wg�ٚ/e���gIp�K��K�׽�z�":d٨M�3��ppdnp��ԃD�PH�����;��\�-)�^��!RǞ>0�r��(��픅6*N�2��F�p���@gt�y�|i�l�(ޕ.}z������<�����k����F�:�Qp�3��X�h�F��P������n����ڠ���&�ze�	��9�;y}j�s5�-�w�r:�Q.X,�%��p�*PF�Bi_r�f�]�{�kX;)�([3���~U8!&j��/M-��F[���ޯ:���ҶS�/=���A�Qj.�xhU(�;- �jg��N.�1�+���Z,�5���Wl�l����z=�X�f+�;Y�񘭫Fņ)���4\t�u⃀�� �ǶD�y�m�s}Q�'�W���6
��+�^�6Z�~u��S�a��тC���ob��u��IN�=UZ���6*B�r�`�S� o��lX����NiÎ�6&a��^�(e�ed��|��-�CgOC[Q��:]���{�4N��zg��u9�Ge�����`��l�/�i�l6ה��y+.�z�]JH�<7;ix��-3>��	�������qK	���U򖌠!ǥxn��!ݢ�U��Y1j����7�p{ ���N��T[�p^�Yg^Ql�r
��/v�%c���bzlݰ�qT�!g��y��$3:��g��6�\1�VT"���<15��mN�>���7{�&yi�1!~��/:�K"b�{m�v������y.�z��N��t�_���,�H�\���+��c�}7�Gu�z�ڎ��wE��|�HHh�>z�s�h�>'��^%���]pW�[l8e#�kp�2Nv��G��FR�v|ǬW0�D�`�[���D�(�.u�3��A���-N4 �q���R�9�k�4�����@�F9J#���Lu�|�;�z�o)�j/�L�,��l�Sb��=+7��
o����C��3�N�(�
���C�^���V���=�9��K�6'\�ծ�x�*�B��4�`���a�:Ie:j��1�wpu�T>�f�A88�
�{6s#���r���z���\�5J�I��0�"�;)6�>yUk�FI��ϗ����+*�Al���A�n�C' u"`n�����ۤj^�YS���iz�.�N�մ�����52p�
�_t|�9�P��q����^��>Rs�1�=H��r�O �z�J3q:mc�^Nd������� *�����9�A^#�������2uS��@��0�{�n�U����G�I��|"��=��z&c�ri����+2t�B�pnY�#���Z�]��R5���/K7��/�_Q��TT���ԬN�L�Øs�J��i�YB!�l�fG��,?l���K�2	�q�T-䡬�V�7��8:�c��r]�o$���T�T����J�Xu�^��m!,�m�V�,��b�홣��ɠ��Wd�l`c%x1���ox4X��1�������ׇ��O��.�=i컺����{�<�Lm�pv#Nq[��uq8�i2�փJ���>Gon�d�Nfe���s���DU'*���ٞzlc��͖^mh`�l:�SQ��]mg��E+�d#֍1t�Gu:�o�em�D{�Z-j�Q���}�[]A����g٩�n!�}����i�Y5ǹi��p�KN��R�Y�~q5���t��Tڇ.
�(���ct��KSS ��%�pG9�N[lq<+G�t����o���*5����]."�8�<P�U[��T�v�%��w|3��=���+�\},X��o>.�j.7P����Zg�b}6Ug{w5QgƠC�sQ�#|uA��>U��,At6�d�i��Pª�z�k�N;�=�I2�hQ�������lEOYw
a��c[rXR1uz��ͧA�˾�.
i0YUx�<�W���J�n�ǃ�{��g̙�ec�V�;X0Tx���14���Q��]�s��3QY�d䷵��E2��)��؛K�k����s�䋸iz�s���>T�Jt0��D����r�MPWDޓ�}��o T�f���K��}ܾI�e�8�z�NX^��!}�EZ����<H�ŏ/�e�f�;�S{`�ͳ,��Y�rk����"��j�h��(�bD:�CA�F��t��V>�xc�<>�b_�l��R�5�<S���o����p� \y4I�o0���"J�����y��\��<zN��CEs=�K�S7�sLߴ�11ܪ	5��CaM��N'D����
p��&�,���Z���Ԗ���2�=���:ǖ�a�]�.F��qq,���r0�4�I �����^��o�u"���w��Y���sl߷&����8��@:�uBy:��5�A�t���U�ӭ^��R�p�@3Y�b��<n��JNup���pu����`�L�MB�3�Gpbz֩�Zi��2N٫�HN߹��"��^5�kO�^#��痁GO[�2�T��ړ=�/C>��Bm'��z*W���.����ܼG�X��]0=%�6��z���K�SZ���4T�˝c;LZo�vJ�,*N$��wM��
�D�)O����,ɽ�rzG�v3���xl��������SEU��l�4���+���G�x�Z��&��p�gv��3i�"ۑJ�N���E�+e�c�7�i<�zv���E��B��qcx�~���Ok�04R7����=T!���
q��1u��M���2I�3:�OY���2���-anP�	ļX�))��l�Q,:�#�KYJήr�f��m�1>����K�9�.Q+LPB�T^)�|��{�"�x�W�&����۳Y�
�E�����r�n�pߕ��P�..��'4jXx�{�� ��{k9�[�����4zWܫ�{>��>Zʰ�Dr~^�8�<�݊�1z��u��+-E�@�f=w�i�4�Y�nhLT9���08T{�tOJ�\3�V��t�ݜ�N�w����A���=+D�$�Ԇ��Y�X��E�:`� ����J�"�b�5�bS�{M���,]�zpTE�;g�6u��n�n�;�j��t91�:�o�o=���Hи�>�Oo=ٛ�
7�Ib�j�B#�W�C�8�N.�����[J� o3��K�Lw��}[�2A�}*�����Vգb���
+z�u�X7k��)�����c�=��6Z������Fc����_�����{8��l��� �R��Of66r/��2��8/$�:�9KL"�n�+���.�+-q�`@�D��j��<Xh��V�F�\�ُ:��ѯ���>�|$�V�t�9�v���>�M�'L���[��[os��9��;sZ���ٻ�l���̉_q�ʥ_(.�t����l�S,M��� :�o�B���Z�׵mf��A���r��
���&��Bk$?FC��w�������_���l:�բ�W�*9�/�ڱ��֖��W<�=�s(�ag�@LL���0�˂��]d�0,�ͥo p�!�N�)��Qvu�X���N��
瓍��ie���.,�nG�)M��ؗ�F�q}ΰ'�db��4�b},��޸��ݙ��C0�a��O3�U�t�z�'p$� �2`��qݎ<y�n��'Z�.7��/���fh��g�H�a6��8�ʔ�r�a�,ؓF��Ec[���NI���)b劸hw�Y�ѓ�~�z�"�����.A��0M�a	�x���ג%�R���'9ㆵ�et�w8F�>$U��A��Ԧ~�O:���Vn�f��s5�d.Κ�AtCz�졿P�t���%.�!�'�Z�/v�p�p`_i�ޥD��������tS�X���2��5s����vɑ�7�p��p�Lk{�M��^o�M�m5x�U�A��sƭ.����J��J*f��e�aw|�J��	J�qԙ�m!�Vw���Z���Nw<�"�.�9��o&�a�ɔ�8����^��#H�N��b�46J�۵tv�0�<�C�`�*S7��+�4��Kgd�����,���sNu閏>�di�[�#��z�$���*&gs����p�b�.L�\��qv*�b�N��>�V>u��7v�O�3�x�C��yJ�dz�텐ym�fb�p��y��5���fe��0��Iܷ3���-c|���̕���W5@�ur�*m̧T�O�:"K|�7��
��hJ�}��]Vgkf���M^.�^��u�R��W>�k�2�0zՎ���
�]�D�ʲ���+�P�Z�'�*ʡ9t�5�L�!��z��lǡc��k2�s��o��J|vjpZ/a��E�˱e͸V�i�>�pi�^���Y۵U���I�{q�s�r� ��0�>)[����S%����eX�k	n����M
0�^�a�֛h,Ծ�F��0�D���8��Ĩ5�]�*�"»R�ʱ���Bb|��0�Yv.��K�xk�����S�4�o��Pn����nRGt�C~*�֕��(E�wh�d�Y�D%)l��Ȯ������5y����V}e�]�� �!@	M#��*�#J�-(P�� �%% QT$QE#�4 R�4�IJP�)@%4�	J�!CKCBR1#H�E P��4�Q!@�@P@��Ȉ�� ɡ(�W2���)��1R��%
 (���%2D�
 %��rr 2ɬ��
�W��}�}�����s�y����*L���ԙĊ�Ž՜�n�����\�5�z=� ,:��HV����ک�Jw�ݕs�ۃr��u2V�Q�[,dIY�'FlA�F}g(�p`�㛸�g�����Nt�gTns�Ou�v�%��*�?����� ��b�}�sMf:����!�}�+�����YUZ�H�PGg����]�^(1�g��>��9c��S�-�n��_?i�	m&��ǲ�����;]q��)���ޜ�p�W��cG���"�T���S#��}�޹̡#��B�-��r�f� �� z��s��r��F5Q�s>mU�9��g]�}{!X'��:^j���2��\X+����<L�4�>�GE�<<.W��@\��L�<�2I�:�3p�Gχ:�Y���-�w�\X�Q(lo�<n5�2��{s�4�>��}<(ۭ0�/s��4Ģa�<aJ�����.zO���R0�{�z�퇣zQs��վt�;ͼ㾂�!O!�jǨ��G��4�BKK���_]��ݐ�a�7��4LPq=j�s�*�o�QcVy��1P��]�r��Ȇi�+��>�.��a���i��݈ǔo`������,;���UԔ٨^��F �к�7X32�4�q[6�Om`��{����WJ<oҵ�Eu���W�
[Y1�8���#��l#1���;zk.?>^/��L{\��ٺ��U�5���y{&f�_C�Z7�-ݷMa�w�'d*�ނ�Γ���P�l�#z�y�S��E��L:��a�{�z:�g�ڋ�uQ"�˳Q=1��j�������x<N�a!�8�|��-1�� 5�SЬp�-�'<G���٭����=��l�H%��wC�Ƹ�DLf�{BjQ<K
��5Nx^���]w��G�2_�gm,���������H�@_F�� �R��c�^(�U�Ii���'S%���T��U����N��YM�-�p���]0�0���2�԰"��
\���*��q;���ƙ��"��h��X�8ԉU�'oO�K��)��������1�$;0�)Z�`����F*壬�r�t���ܧ�V�B�ѳ��Z�l'x�Aa�~�!W%{����rNG���#�4RGyf0�R��>��X|Isc���Sc<��	�s�=�¹��E��p���Ł�Z3+�VӖ]%<"�،�1R��!@ؽ�:��w����k���T�u;Ė�m�p�,(g�:]S�lN��9��zv�#��P#iׁ�D���_�9	C+*tKxb%S�T��:Br��������>\�_*8��p���_���I�|��[TgA2��K�ox��4|Ќt��x��̤�5�EJ�tlVR��t��:��������Χ��V�|;m���>����z]����M�]O�0Vu��>D�!:?U���??��Y:&-��fԡ�%�u���1�itp��ה7^5>\lx�1�`���fMw3s�8�*"[�;SQ�}:��P_)�E9b)��%,HH��e����wVr��V:�8���j�$p[Se����r+;�0Ó'�c�^�WOE�]xWc�C��$���ê��Z,�G�������
��[	����ŀ����g�;O�������_���S�N�t�<eW	�,Ml�φ�I�;^�r˞Y����̇}��~ٽ5�
պ�QqN�!�!娭&�79�(u��B$���N)ʎt3m��p)�#gi@
>�OmC����3�j��4IULJ�SE�"���-'Rضױ��}&ha"o��L+��L>�PI��\�U�)8�j%V��a��{���ȹ= خ�ZUT�D�e�y4�ΐ%��RJN*y>�&���$���ڼy�гHPf귢�-�n��w@��j,&�7J������oj���p�i�+�@����^n����v����5����*ͤn�w/ue���`>�'�74�v��b�Ff^����v�,�;��Tc��a�u�?f8���=X���	����iAd~���:Ŧy]����(f�O�Kpu_�Ǉ��0<�9�G���B)'��'��2i<����:�]K�)��Yh?�ƅ�6�
Rs��P�����P�k����V�K7"t����af��<�)6ycGW����:l?��j�cd�b7���n��w%Rľ���s��p>��X�5�Cc}c��}�g-����R������>�����O=������v�483�@G1�Цk(һ����;ၢ��F7^ڸ�g�
x�oJ�s6���M����gD�ݱ��xh��x0oD\�{
�<g0N�[0�.Q\�Bͽd̫�Z���KG	�b��zV*��F)V^{] �ହ��q�������CJZ�Y�,�0���8�� \��Q�UHrQ|P��R������E_cX�����e�a�sR��h����G(/V�D�O���WM��9��O,�=��˽B��sj�{7y&��c,�:�P�0^I������l���O��P�O=4ed˃8�I]���Ċ����3R]�x���l�bbQ�^+ńe칪��9n٭�j��I�[霾�0׳=e�Fʷ"�%>I�O/l��p��]��G���u���{v{�4����MlM����}y��Cg���O�E29B�1b���~��zs<�Bf�Ŷ���y�.���x��ix���^��=a�)�_B�ԡga�%��F����;e�u��n�n�6&n{��5
��:g_���Ts���,䟠�z�J�ڵ��_.Z�8*�i���\]U�x�_8�u�\1'�����u���.jP>��h�ԗ �>ϒ�xe5��q����X�'�	�O��́l�y+%o�G��XIN�SґT;ڬ;�d�K'�f��n�v0��]Z����u�v��BG����J�8i3�q1bj1�[{�$(��\��F�봻��o�h��yv�
g�Tz��qq
c�T�ȼ}[������ a_�!V�=��s��JW���q�mr�8_�%�*&63f
�:�-��]���;��h�������ب�z����w�m� ՟}n�־�cZ��h�쭦 �� i\��r��c�h1�07�Y�5�;6n=]z�����e�8��z��GFN^'�b��.�UA�֎��qV��2��
1��"�tؼ��<r�!n��E�}k��T:^{�^���ѷ�ֹ����;�gFǝ�G���U�=�x.�~�u�IǓ�k{�@�
��D��1���nA�o������wZf#չjn57�6�}ܡ��JuL]44�P �s�w����ǰ�z�s���|��Mc]����'���#\$̪���l��b�P�Z׾J�����w�/¸�R�B��2�� `�!�NX��|����yLzx�N|׸�+��a�B��J������=yQ�n��O���s-�dcH��vO��XĚ�<�z�-��@���c|��	��@�H�咚*��۲�`�
v��O^���a��+6�[s%�Tk��@���K���n�����y�R��Z2�r��P�҅�ø��;���5�u�]�P�+�f��z�-�Y�Э�F�Gc�݊2ϾHU��%�\�����t2�i��kmV�qԯC��e��i7�=�#_��:Җ�8��?G`Q*D�v��+�����ߖ�1pϬ�����<lH��洢0��qg���X�D��_0�zUi
a���Ӊ�U��K��-�Q���/{sw�5�sj3��]`o����<��sĬt�|ZC�d���;�r����os�Hz^o��%��׮;�,n6<lX�;�^LjqD1�����C� ��1̎�]����+��o0k5�d1�}��LjxċN�����$�:H������E��w/\����PY'���:=�	v��.�#�6�G7�7F�K��bnU��ziw)}�����3)Z�6�F��D#3z�B�V@������W��#��ޱ�gýLm���Jl�V���j����N!�3�Z���Uf0�f:�q�*ia�l�`
�Jp;���sv�z�Oy��L����[m������.�-�P�E?y�;��J���Q�,2�����ީ��w���5i,öz��ꖡ�폹<ӷ�%����R�m??�>�.T��}{Ʊ��:���Y�h2�DX؆��3��<x.���-N�ϑ�Qޫ����X]�vU'xj �6:�vɴP�~�a*W+bK��5�R.J<
�YH�g�]Wl����|^�)��$Bh��������_)�C,D�ٍ�YbO�T�J��]x�:}�JCԴ,��<�Y�9�4t��D�ì��]l�����TU��<�A�Җ?w��n���c����	0փ�)\,�Es�R�x*�����Â}����?x֬&;n��2_j	�z�q�cͼ�o>��������bcZPb�<JԮ/	���e���[Ps��j-��x��KQ��>�\^�k�T<F�v��91�|!̾�d��c�WG��G}{�|zߏ]yp�Q]�R}f6�tTл�Ί��/�\�-���2�%�J%��7}x��a��6�v��P�h�"ĩ��D��v�c��G�)-�P�Z61j��y�U�ۚ�[��K!�0rp��:����R�^�������齛��\���M=,33�c��ؚ�Th�a�=�0�=<�۵����v�ϫ}���a�3q�I��u���ߛ�{<�tI�� *��w�+8,�׋��Lz��d�Y��N�н����=�H���a0'�iO�z�ڵ'emm��;�;[�aO��M���j
�����дp[4��M8q|��5Օ�[���no�ƻ� ��a��n�ʮ8
�����B�O0VT���C�8���L�����>�Ӡv���t�����\�:����7���|%��u�X֘�GG~,�6��=]�e�{$�~�@�����+��
��z*}汳����"�P˗��A��c���{���^�Z'èV���~�Q�+���DO:����{j❜:Z&��1^���K$�oӈ��Y���&P�j� GTb�MF9bk��cT���#U1ntF�j��c#(��dCgʶ�V:&ޙ)IMY`�꾽�ʥ���a�uyH>�T��38Zo�U��D����*�;�-U���[�hf*�+>��"��g>аp ^:�v]���pg:Xh~�v��o!۹3��#"W#�z����i�۳,7��|�z9.ވ�<�e�Q����;� k�.��5^�����ʖ��c&M�g�uEXԃ%s��v�퇳B�ޠ}���a�!�K�*	Zr�Jj����\�(@�wyGiO�׽��V͒��Zf�\].�U�=��׈�E|�[e8���8,���\�Ԝ��6���IE�s���$��He�y,X��,z�0�4�"�;ed��s^���x�e�)�Ñ�8;w��QyӘ��!p�k\6��ʷ4*:"�0j��č9�n�jY��v��i,�D��D�sX%:�N�Y���n�v<�%����\�/�{`�9K��os�n�!�L�C�^�s<��I�l\��@(��P��8s�u��B��+6����t�Ȩ#�h��K�a� �>�KEᏗŖ3�񎍎��ͺT�n�Wf�m8T��E"�^T���^X9��6�KU��=4�'%�O�[�*zJ�^��oo���$Ni�ւ'`w�g������P��� �ʑ#���-DT�r������p��/fs|�Z��8�^��^^ډl`���l�gir��do��D����o���X����ȊK�s��,�̤إ�Px��S��1�ɎI+�&`��g@�+���R�&ц��ǹ���:�j1���N\��ib<]��.���os_A�.��U��Q��je�0��T�ȿ-j�0P�� 5�I�Q�GE<�¬SV�?|�Kw����0�m�b�<j:�^>�����	��I��:��ȝ>�2��{n
�5*tZ�Uh�V�xU�p+6X�'B@�QA�Jאޜ
Vcg;0ʒ��X���%�2������fx�=L?�R��r�=1xx�z�¡�*8����>�!���r�B�%;�����e��^�G\�Q�Ț�q'Y�[��QjQ(B�Ӯlpp���z������w��3��\�G�U�s�\�1#�R���b��ͭ-y��E��ȱp�)d��m���CVCVG����:[�)�#H��`1P�m�r�޵Ʈ*����̙� -�Rc�D�녕=}7Q����1��
��+��J�R���PoS��|�o�����Թ��%�G�:Oa۾�CY��f���Z(�5$v�2ݤ�kP�i�t:��^/�k�b�\kyq`�y�2мL�6�Ҁɒ���4��5�U����a��6ʹ7,+�V�55��1�"�'-T��k^}��	�u��x���g.
�f�SZ�w�s�ר\����(�S���:W&�L�f�y����R��k�T�xW0b���㵭����f�9W@xsN����C�9t[���W�?|P$E�Vw�.4��ǥ$�wT���Gy`��ܸ$�ν[A�"{/o3)�|:�X��Ո/���䛧��ϯ�7���"�<df�YC���9�����7��cU�c]��M))� �v������4`�B�<a�ݮx�Jȕ��Q�UoK���ܴ����F����_Y;�g��Ǿp=�0��@�F#�1Y�x+RC<�Bw�;o|��$Sp#�ܘm-�i����ܦ�*<8�Gt�*�Xք@���9wN��f<�g+�,�cޖN�Ԓ�1j�Cn�j�B��Q�m��e��)�s=�����.Gܱo59�����B�OK�������h5�-��gu�(k\�S4�*$|��2��$H9K���Pi��ʴގ�*l�)�9m>;0E�B﷪8`��;��P���v;��ˍ����_b;���B�Ò�jۣ}O.V<t%�ۋڊ�J9���ӷ����{�I��y����
���(�u��)v�B���u"��<]�P-c>��}�[�й�qu=��U�K�5nT�,�SnyU��=�S`�lk�%��;�F�^���/���:4��J��l!Ң�_cs�Z���`�vmɚmt��[O,�� ظp���TZJ�B�a��Lu�"^X���`�F����J.>�si�.[����%��(�,��j��2�E,T˾�3��/A=cc��3X2��k^"���]_#T���]E�(2:9����VSЩ�R�O����T�ap���w�3n���\��;R������}�&Z���47�S�E���t^V����P�H^��qD!����smDV�e�&��9k8d�B:�ֻd��<�^N��y���O�e����,��)1����缃��7�V���)�ʇ[(�m�
�:�ۉ��Պ/�������U�����9eH�S�=�z5�̘��ܷ� ��eȆUT�;�nX���x��q=�(�H��m���We�u"����om����"��E(T)K��W �Ȅ~Y°'[ƫX�__@�R��ݛ�m$X��RF���@�𻛇.�)V�x����ǹ4]Ⱶ'%�2j����q�=���cN���F�2�=�xp�������h�\فEK������7�do]e�D�:��ͷ�s{�W0M���7]*̴���$�V��;';n�ݵdEJ���t���u�K��tx�`GV}���z�B;"�W��������y�僤��V�O��|���:�|n������ӛ������cd���~>��4#@4��%U#@Ĵ�^a�H�.@�BQ4@��*QI��+JR�A���(R-	@��QMRR�#�&AC@ґ�C�ѐ�4Q@��@R�R5B�`��4%	KD�P)�9#��B�d�)@ҙ&T���%	���ANN@&@d��KC�d�%U��BNE	J��H��� PRJ4A��}��y޼��~oǝ�[Gu��\�3o(g�`��{��Y�����8J�џs��H+��a+{�ʳwE���a���;/�Ѝ�9�򈉁H�eP��mE"X�|��O�BT��١���o#Ι�����Ν����ze�z���� t�x�'^�ZQ����k>|��j�j��&aT�7�=8�#l��J�z���n4�.�9Y��)�V|�tI��L$�+�"�B�꧶�k��ħkg��p��S�5���A��/)���9=V��L � �;b�
�t��龓�#H2�	���81�K=��Y��~ӂV�F~���o�&�2�dZ�``�x�N���R���!Q~[FTjFȯf�wU�Fc��˥���'� $l2,jy�0�׮*zյ�mh±lk�+:o��r�7�U��S�.M��_�>6:���mC仚���ZP�^%N�[JE��t���aC[��r�^��Q/[T<pR��48{A��nY�B��!cyR/`h~��H�S�v��U�0[M�cy�	�%��(��G�2nA���R�2_-)��sEz���(4uF:DױJ�%��|���v��\�
�%�$
��@��k�U���x?���-b�#Os�X^>j�!����]7x���)I��	;f)4eG���*y��˧�-��]!1�P<��eLz��u3�#�[���(���;tu�ځ<��2�����z��qf�Izn��XS��Ki3kf$�U�b��.`8.pdX�a�"8LK�P���a_OyA�0^��9J,^y��YV�֓"���^W^��N�2�Z�P\���%*�R&�~��.�0���ۑ�����9�58��Wu�c��Y�rk��= #���*X��������[�֌��_�._<���B���nύ���;�c��V|a���R��-|<�.ۦ�I��G1ۗ��,�zx��b7p�_�k���~V�EE�� j!�z��70�x;�%��	܍Ď��\��WB����q�SOK�����^WlM*�����_;3��{���ܞ�E��NUK
M���+�D��s���ߙ����i��u�:A|ֹ�{����d�#�o�Ѥ+�F�5���=M2���pTq������&��=��w���kvU��_�u4M��"Q�Xz��=i},���a�)�+-1�>�c�Օ3tk������t�n�Q���5��7������XU������n�֣c�4�	M㕊km��������O<r����kvʎ��%�y9X�� E��.{8bW5b�R�W�z�n�$�`��:jrb�C�淴2���Q�۳L{��I�֯����m�Fo �ew0D-V֋��n`Kcm�/qY�vyf{u��ڱZ 䔃%|"y��1�����>��=�����R7��fozp{s�>�q��q���L�č�-����� ��q2�D�ҠVt��Ҽ!���j�Cۜ�Z�pۈ�GJ����c��Mm_�g��d�W���/��/�^sS�?���6H�!��[U�ڒ˙�8.����O���
<=[�L2�&.�Z<�-&�~)anw����� �����D�t)�Z�t�F�o-�g��Xs��=�&.�%�����J^\OLU
�R���W[j�Yw��.��������Y�wDL1��* ��8�\'%�)yN>��-Z}h�����>��*B���u���7��B�K��l��׈�E��*�]�w��U�[QOyفz�`q=6��9��S�g7W'��2˷4*:�C�X$W�ۋrK���;E.Sδ*��'�E�9��D��kT6��ʷ4*:)ׁ��:{��0��z	k_AB��0��T����5�t|�M����g��n��؆���`������=��������u�d�^�a�ʚ٪����.����3*��]Mw9ђ����ss/�$ۜՈf��B|���y��r�jbL�e�î��rh�Vza��07ת����
Cq�\́P���2&ӱ�6Ɏ��v�N������˯dxz�g�u��-R\�6P�Q�=q�$�^��n@Ӂy)������F��Aaxu�ޢn�bJdҡT� ֖N���J|kf���gpS���#�rrud:�RX���=�`3�NH-s�p�5��D�͙�1�tՋ�5�nJ8��|pVYH���Ll~�F�3ҹ+(Y�����Yr$W�������cr�혜}��-�����ܙ�#c6��-�ņ�U;66��8UW�h�� �=�D�58D��7ޚ|�c�� �Ss8�-�޸p�xP���Zg� ��'�桱���(K3�\����w�2]�:���o���_�։�o�u-���;�����V%�>�-T�+U?>�Y��.Iծ��l�/���WS�:�|)�h�3�ަ]OD��yկ�}�enkSĎ\�Ƙ��_Z"v�w���q�6L�*��B�"R�X�ɋ�(U��÷&V�̰���7�rŇ�����/s�}ʸ�%1<`)B�f}��K;�4����oF�6�JT��?go�s�3ݖs�oe|q��ib�G9�A��������3�z�${v���p����3s6|�d�э���C���2�0j�o7��Ĳ<ׁ�Q*g|V�����y�;k�SU�鼆�l�;s���g�mե��xo�g��,od%dy��x�g���5����n������&���X>
U�X	C]HB���&>w�lC�'ޙ�����Q����	Z{hћ����ߨ����W��k�c����2�ꂆ�aߪ���CP��*x̓�a�>��*^�;��ZcèD�O^,{�-yhVeS��'���Ьt�P[.#<h�pv�������Z�=Bq�J�׈�X�^)��1,z�x��R�ߖ����Zf���~���Sg��4�}Y
�v���x\�X�D�@�k�:�}Wp���k%�ڏa���<F^
p���i�gt�+9�aL83�d���N���9Rܜ����o��t�',��e!5�ً��c�Ƭj�`�?�����+KxV�v�&��yp���7�FA:�H��о�e1������âV�F���4�էsٸ�u�>��>�0XX\�F���t<)3�Y�1�{՗�*3e����q2;)�h֕28�2�E�Y�%qՎqa�W4����hLt'�;�tQ(>��K�I��,�-�(�-I{H�}ҹQ��|�N��9c_wWR��1�fu!��5@O��Ξ��y�ce�����r==p�W�ǥ.�zI�gQ��1����$�&ӫ�����::�nD,�t�\C�����ύ���;�^7+y%X�x:�M����S�"��S��aC#[�����hۇ V�ڨ`�G{�����N-�뚹�K���ޔMoK�Z�ֈ�~i+Cy��.���I��k��0�7�yN����z(B'��#�1�;����T�ܝ������z�pm4�Ou��ŽfΏ|�/Ptuh��h�
��N,B<�h���0�ҳ�tuwe�v��р�����j����z�B�i�f��b��<e.k�x�/���+�4��{�<���#�o��v�k�|І�T���P�Mp:�L��/	(r�sT��CztY^���Iн=6R�w��e!u�
�(y�kJT�XR���X��v�{F�����=7�Qc^��u���¡9"���NtLJ�AbD*��=>Wu[�ś�z�z�5����d�y誴6�� A��wmM=,d9���XЋ�<��Cg|��9|t�b�#�M���{v7X�;��=��7^ ��eB[�S���Պ^�_�k����'���
��l����ł�kto{���l"���dMq]��ˎ�p�#����N���홗��Dq�.4ok�ΙakW�������6�Vl��/��4��g���6%�ۦ�52�	U���ef"�?s��kܜT;�Ud �2a����������>נ�Z�	U�&+ҍd6��EeO�ɦ^t�.�l�[�vu�L�N��FAx�t��i�k�	"Q�|��_�},�g+������S���ӯ1H̞@�S�;����b�{�$;�Y�Pt�&�axX�ڿ,h��1f��m�P��ܵ��ZY�F��M�{����0:�]N�c���c�V��U=�[��(��󚰰�lX*ϧ���Ƥ�vX�fB��r�Vl��Ҽ���0*�z+>��l���x��pn��ix��~����x�YlfV�ʃ*ׁ�G�o�L	w��Ww��|}
EօD.��C Iۥ��j�ʯ*qY�	�
a�SS�x?��hs�
��eR@߂fٿ32�4z᡻V�_j���]]W��t���,B>�F��a��R����7�R��zb�8��H�y⩘��*��W8q�tB�<]��yu(�#�
�|	MX�+�
�Z�@�Q`q��(�{��S���_�e�o)��\�ag� *`�oeqV�ܭ����B�����0�Eƥ_�Y2Vf`���[ѭ�ǹ$�G0�8�.3����26�<T6�u��Η,�f��V�іR�7�+�NŞ|;f�����׋�W��JqRň����R��c�	��d�*��!�>Q�W�1��o�u���4U&T͗2�f�bxޞ�N���\�z錳�X��9���rw��ƙK�UO�t��.0��5���1���s���Y��z7z�}�7�X�٣+�1�A�{EAy���l�	��>�賢m%-TF�5�˅�Y^,f�[�D�:��t�#f���Υ�2�;X>uw&.[���~6�ޯ_�\��.Z�8*�m���\]%+uܔ�S-s�ytR+8�*�{]ה�mW-��ľa�	�)�֖�¸�n�=�ȭ���J��G0h����+�A�z��+�NH4Ԑg���p���c"Of�e٩��!��A{�⡶�@՝�}�&1[S��G��2f��Tt�N�}��Õ��U�q<��x�.�>j���s1m+�w(e�#�5��Cq~S�ףU;2/V����g3DW)w��jd�mS�S�x��`�'V���֖����?3P��ش��_��aC%��]~"���vt�&�ǅ�w���\���pP��Fe�c��JA��	�q/�2S�ڑ.l����۝��{/ar�#�Zj��r����R6����ۓ��d±��P�I���(m١����1���u��ŶS�c���g�׾�i/�o}u�K9%$#ʞ�(fL���� �����ԫ�9nٿczYb������' ��B�=���ټ{��y�r���������/�y��W8c��|)�#~7OSu-���wV�E#�8���j�Q.�bþ��V� 9H�9��e�1��B��5�'Y�#s�=k�ɵ�{��d�J�N�,d3l�9bŽ��>�mﰬ%֐8o$6�J�O����{tb�8�&��;�\J�q��,jƬ�K���vt�4%�R N����.�O���hj#B�e� ��W�I�*]��ʺ���!�>͓O�Σ-�3�(oj7�o�|�a����,S�,��<0�B$a�B��a��پ�C��)�1[��]�����rf��LO��u::�_xR�~����Ct��	�A�+����k;I�hy\���ވ��_fu�7δPn� _��0*[`]EW?�����-�hZ��>�Ms��>��f�qf4��Ab����S���-�4^�,��U�ɽ�W�c�n'k/3���(ɼ����+�_Y���p�2c+.�,Rޛ�*��)�ֶ�+��X^�;��g�n_f�ec�=�0�V�OTT&#(az�v
]ڧsK�tL�n�Xkc��O5�P�l_u:�U�R{����[��:�i�1�hQN�&���u)�~��e�Q<F��o��C�Q`{�	ϧ�г�^��3	~e-s$	u=�z+2��
*t"z��`���[1p���X�7�>Ll�h�.8��U�Β�w(Jj�󶮖FHT��GY�3�FV�`���v8t������!dxvsg�o3T�V�淲�kX�V�NeĿ7\8��m����Y"�xRg}v��/c
J�xXqjA�׊d%��N�>�#@��6Of�~�L����X�����'��`e*~����8�6��ͮW����PD�oR�Їe��u�xdw'=�eTV-���Mcu�y�Lv��a��Xؙ|X���@�q�Q5��7t�Q.�F���[�t�!��ޗ�Sw'=ݝҭ4υm<
�q�P�'����5�Pǒ����*b˘�5ee����j�z۾{K:�h��r�����x:��\&�Js
�|sڢa��{���=R�b�Eh��Z��x���3�m'��,T5��([�5���٬����Z��}�W�h* ��TW��* � ����ED�* ���TA_�"�
��D��
�+��W� ���AQqD�AQ�
�+�PTA_
��W������ED�ED���
�2��t�U�)�Z�������>��������"��T%"���D�UU�@*J�)EBJ���R�*$UJ��HT���I �*�"��TIo��R�� IAJP�W��V�FJR5�HH�R�T��U)R(�
��J�CT��($�EIB�hJ�h!B�QJ�T�*�UBJR��Q�B
�URE+�D��UHUBJ�R�IAJ��"�QH�խR��� l\���,L*���P�kf�E�l�[J ,@5R�����+Ej hҰ-
U D�f����"��2�HT� ��hVX�$� 
ҩE�[X�a�J�QcP5B6���� ���mV�F�cU��B��`PQEJiC6�T"UIU�ܰ
�
���B�  �B�:w
� �E
:n(P �
�.(QB�
s��(P�B�(��(n�����UCU�Zkh��m�Q�JJ�R"N wmQT�5akV�,�b[@��hUE,��@PYl��HCX֔����aQUPJ�kAT)%J�N �Ҫ��X hJʦ�Ulժ�[V �����i�RCV4m�0FT6kl��6���JTmTJU%U*�%(T� ��4 ��Z5�1��eRְc@(S1keP����ɪb���X�j�YJ�(6A�i��Ac�-��a�Ґ�J�� ��
�5�U%@C3A�cKV�CSF��
6 R��,�+��Vkj�Ҵ�VB��D��P$�T%*8   ��P�@+l��SZ���aT�2�5�TB��� h�0UU%�
Ed�JT�R��**�H���   l�ѭl����h�UQM����P�`(Y,P&
6��m �Z %���Z�$
P"QP��  ��
�f��ICS+R�E0�V��T`PFR�Z���il�Xi���)Ybi��n�B��   ��RTTLC	��4M1��$�*Q������hb#i��&�&	��0`��E?�SF Ld`h`#A��4�`���d�=)�FOS##F�MO5 �IfUJ���&L L�	� 7�ݻ�i˗��/���B������[ֹB�/-�U1�Ԭ���EEG����?*d�:�*<�E���C�!'ȡ
�**6D��c������2C�0����%�� (|h��뀕H��A	 0��������僚X~�}���,�����B�oZ�~A��p;�k���Ԑ�����B�J�g����V����/T:u�Sw(�qmm���_���4��C*V#�&��(^EI]]��J�r�cf v��0�)�Nc[�NB�i�&����R���U��Șj�R�3r����6���KK8��p���mM`��Q�zcqj�a��QhAHA.��{!��Fv����&F�L�[ad��l��+X�e�����G	0�{���D�iPWGwn��I�O	�b�غ�V�J<�V��ifXb;�ef�`�f�kڑk[t��(�24��	z��l��O)i�N�-����0@�m� #Q�N0�m��
�fe�aQ�n�4�$,4����쩔Y��X.h1-եt���m�&j �n��-��Qv�k��f�قژ1&�v�i�`ZT�K7mǔ�*4P�0�ו2��bڡV�����	1������v,[Z//VDEHM3a��%i��!����S�t����S4�:4h�.��+VHw`�V���H�>�ȷ�� cI��w���7Oj�(zlRn�Z	��ed�U��YIR0�mKO���dA��T���ի ��A(�٬��w�CI��[r70�N����1�f�1 i͸5��n�a�j�ٙ�y�R�`�Ff����T�1j�wq�܏D������"�H����Ѷך�b8�a�:��������购<f�D�K3fn����2�)4uV��	�Xj<{EU�{R�����`�{KaL[�$1�r9��ےܽ�FR&'i�aT�Zy�V*u���t�Yk�3;z7�Io���C�Ԍ��W �TGq
pi���Y����`�峧sT�J�W����0`��[>@��2���zh�j^<�&ַ,��aG��^�������B}os�g��[��D�ٴ�VL�yR��f�[�$�fEQH�����7�^e�+�SX�7L^Jz�B��Ү�D][�Q��n��2��w��Y��H�FLz��z\z��g*K�{�ŭ̽���2��	�T�ި��FC������f�E[%��=��t��l9��v��l�j�X�$;Ld�4�&����ъ��ma{M�vhy���� eҍ,�fc�ôi���Kg��Ƶ���ӣEe]]醬M��d9�]�����#U//�]b�Ֆ���U��@��Y����Guc�t[��,�-������S�s'�� ��r� ^�!j�]���qL��GM��43c�x��;��{��m�Y��n1Z]��]��Ut���p��);��f����m2Յa�ۗt���ҹb"[jBH�{�ҩ���c��1I*���7�U(BxtQ�!������j#:��G^�weʊ��M���u�@]l�3�E�y�Հ��`mU��GI�pP��Z�k��B4��u��h'r�ovJ� �� �#4�&�O�A�yxm�Q�����N�$�U���fVRm^��΍tҊ�fۥ��VU�m�p�5j�֡e�m��
a�^�	[�V��&��¶d�On&�C+��'�e<tR���c�g��pGi�ں�N�nk*���,ñ��͠��ŊX*��ڳ���̔j�l�	R��	^^�i�	IԖ��R쉊���/a;J��*:ۦ�Q�LU��>jE,�Ÿ�;W��;��w��x�v6�Gs�nQͭ�M�P�,V�li�U޴�b�]Cn�i�h��u��M!�y6��Ň��*;��M�ڡ,���LV::�݀,�n���B�r�q1�iǴB�Ԏ���)��-[�k�5�ᅙ�v%I�(�D��o0�Z��2B��[ޜ(ܣ�tKV�HU�x+sK�e�������Dn 6��R�N�\x�,D�,l�VYW��ZЬ��c��]��F5�!d����"
@�[w��q��+7��b<�w.R�/V̵�'�]�z���q�
m� ��w)�Y[��抽r�d�x0l�86)wz\ē��:ݻZr|Mp��@ХCjQz4�c�ͷ��dS#�շ�KM僗W![��Y�
BQ�X�`6�Q�k�œV[.��&��KeKW������B*�sKpJ��#�Ԫ%^�� VY�Q�Z�@�Z�ذ#���3qdj�he��ki%n\Ih8$:M��i�N��[z�Ơ�ȝhcfB*|��h�r�{H/n3��;A�j�j��Y�#&E.�Fc>4Z3eG/(ӓ(]b;W�����I�4#�3�Km+��S`�%©mӤn`-70m�,խY�f@�����{IʧPO)�f�j����\�)�ج^�r�T�l��P�����dXݲ荷H���[2�v��0��� ��-�g��F���Ŧ����!�:��1��b�W�i͹E�v�[�`�) ܔ2������L7&�tj*A�MP����d�0�ը襻�l����V�]:#>M����"t��+B
�M5���h���n��+cz*C��.�PB�U�2[����}˫�+fi٭lB�!��v�������1H�e�h�-Y׹� �2T���&Qz\����{omd0�,�J�r�\IňպxVE,�6��o(RU]��K
��`j�I37-
�� �v.,L֩����B� "��l=(f#���qKH;��-�h	f-����5�*
�T�'Id�+C�7�n�!eb���F�L8��)�\Ɔe�I*h�fJ+Gii�C[u�d���٦96����r���F�#^fH4'�@im�j�I��v�
kM���݅+2���o �p�Q��FټXͺڼ�)ϛ��Bl<�f$�&0چs9֞�Y/&�h���T$Vľ���F�FBN��	��,R�b�md*P�6������Zܣt/�з��Q�h+v�#WF�W�	kC�z�5�բ����#�d��1��c Op�*y���N��K`J��+��d{� on[Zޖ܎ec̶���V6�B�N��-�Y����6+Y�{���㑏�ɢ�Uؐ(�,v/%c�g���16>sPC,<�&^֭w�V"JQ�5
o$�ST�	�� �U>-�JJ��ܬt��{Rֺ�����Dq����`b�ǗC㬙��V���+SwhK��e2pö���l�d#3[{y��8��%$.�u fn�㵴sF,���& X5��՚(�q!t/^<�F-$6���oЉ�7�|�KtQ.����Z�+5F��v�|-����ʺJ4��Ƿu�>��@�AL
��5)�(�8.,G���*U��Y�re�b��cn�V�F4+k2�6���r�w�Zy-�J�[{�h��3� w�L�e�AVĐ����7��d�Ea;�Z��4�^-֫x�^MD���!�@Ӷ��"����� *�
l��wV���ȕ�Џ�O5��ݙC(G�b�́�u�t�l�E��������342��-͏@m��J7.��s�PC0]b�-\�B��U���.4̬t�F��ө�U�̕�%����j�*KF"�I%�V�L��l��k�&����.�������/ҙ9�S�Q�8�xL�ɎD��D��wL
[z;��ր�W�76��%!4�Tl@�Po.S�n3��:\Vpj�T����lYQfb��nؙ���z����kR96������d�x�I��I�ۦָ
Ԋ�P&j����P�����ҳ����ɺ*
L��u�]�B��m9z���J��m��.�J�BTK��Ez����<�m���.c���V���7N7t��&%.Jh�OP�PD�ܥf�̨YƐ�/�l�V�W�aF�(��˛R�����t/e�%)���V�$	��)=�&�KT�cH���7K�
���*���ře/�C6YK^���T�mÂ]��`7����x��r��5(Pk��&;���c�	���3^}r5����Ҩ�F^ޣ�u��%]n1Z&���/6��B=P9�6�R�9��ڇڽcњ�*$d�F����:Ckp@�":��a1����J �QI��K���M<���(�`�Z�8I��T�	x���R��56[��์��1�v���2�8�	�pЫ��R��af� K�����;MHvʕ�m�[�f���3v�[v�5�X��,�P1�b�4����2����fC#jJ%��VV]���6qV4���q�*���jV.�^]@х~	��}m��V���+CvE���i�sI�&�[3[�,H�b�m1��.D11d
ViQTE34��y�᳈��wA�[�ɑV �׭|C�່���m��N�+n�.𬗄��&����YZn����+3�M�����op����j-7�V-8]��
��s�®h��c��J�z��"kH����@�TԔc�*n`5
ooi���ֆ��nS��!̬h*]Z�N��)�p�c����̩t�H41P��4� ƶ],����@�V�&��]�F`H�ג�j�ՓGc��kK�%90�]�͗VÃ!��e���`\�Alf�e6��R��H�f�Yt�v�5'*�7Ih���z#�E^хX�7q��Xj(�[����w��d�@R"$u��
�R�t�m�3�AAR��e����L�n���eXF�WHn9�
��.\Z5?����
�l�ں	L�rK5�Q."bUŮ��z�'vj^�#I4T�2mL������Z��X�k,�ʘ�U.��2��N�����R4.�6'LKT�Y�w!�U\Yg����ԓLr�� �ό5l�z&�t����mM+/�]c;P:`��r	��$Qdm,�+0Y�
�(G������J]ddT I�:�ñ����鸷`��
@�	Զ���.i̎��@J�b�mi�j*5WE�3v�4��dj�"k[n�G	W�0��K)���)�cb���6��X�-�7�$P�5j+��CB�4�m�.;���2���=����W��1+�4&l\ߕl�
�	ߝ�φ%�ұ�D�I��nTt57D-QJOA1k�81�
�4�t��)c�Ǯ���L�4hR�����9�*���a��m��]ԃ1�26�ӷw��"��n�s�5h�*`�pF�b�ے�����iT�Vi�<�I��/E�Zc8�f��N�a6��I�%���>�Ҁ��yV婻�֑AGu�`��A�x�ɩ�z���j-ѕ��&n鐱�c1n衷�rmA[E���Tm7u�Rem3"��%AH޺$%f�|����ض��{�%6�����;l�Y׈���u�){j����]@�1w{�@�+� P�ُwmln�;���J�h�U_
��\wb�����Psn!w�]h�Y��
��X��B����F&�J�ҕd�ñ���dX��+*��3eF�wj騶�]���b���X�UrM��MU�+1͠n��;���v���C���jм�*a�����V��NdYPJXE��Э���ʵl�x)R�$�v��V�(�SF�l�4f��o[�"O*+K]-���(��pUБ��m�im���9�2�%`	ڬɨ|�1JYB�2�M�`�L�u�t^�,[��b#�n��+!�.�8qԖ�N�
�ȝJ:��R�,�rf�SKT.��*�`ĝ�	�-�f��]��Y��8����N�ݖ��b�����>��0V��֊��Y���r�R�t���Z�W-��{v�F�<��^�J[Z��X�U�($�a��e�Tݵ��%F�n��Ҩ$�[Y˴S�^���32��4T���̺
6q�B���MUa*���swk{)%�*�M���-�쉚:u�*ڤ)dٗw�c�J`t܌;��U�ڔҦ�O�i-�GK��flxv��������%X�N
B��p��V�L��:u	�񸍪m&�1�J�܈jv� CR�)�����6T�A-�oҲ�L�u���1Ӭ4�!#�Hk�[�J�Y�j�i͚cL�t�So~�I<�-+wFj����n'5Y����	3�V����%y"����a�O^`yWXi�a���7E�u�t�̺�t�G���1��f�2Rj��Ll�deB��j؉9q �hƾ����ѯE��0c��D�*+�"TT�A�E]�B9���l��׬O�w��R=�NXݱt���fi��ި�?[��~�y��O?��=:���o���7��4�G�9��P��<�/�C�w��#�HhnU�=����ɯs���r�U���Ne���2C{���{S�ݮ��º�LZz
}G7*X*��3��J>�O'C}��9J]���Vj�v�$_r��8�z]L,t@&�쩆�ܠƼQ��W(�bn{o`#���D�����J��Ý\�4�e����vP�ht����G���5}�y��4a�Q@m�5���p�U���R����WؤF��a̩����X�vТkd{մ1c��e��U�q�a$�Ǎ��� \�%���6�:���iwKP�����^>���j=]C`�G��sEM�:� ���X���N�lgp�ň�P��a��=�*��盷�Z�w��Ϙ۫�lԬ3�U�̀�u�Ϲ�����IB�ѝ8U����b]ǝ\���W�el;��d6��Ȟ	$��G/3��!rr�Sc�l5�L�f
�b�e7ج�g���,F	/c{j���R��,u��͝]���膟n�	�;��V[�e��e-���k+�8�l���C:��Ǭئ�����'V����Sb��Ew���R8��0��&�e�prH|�����8��uH� �"s��D�а���-�*C�+��3�N����Qi��舷�
V�T��6�Ƣ�)����Z�>�jQv�FwQd����e�Lډ��ݔ��,����o:�/�%�NSP�qt�ev�ǐ�u�zN��"x�Y��Vf�YӍ���:ʤ��)��͖�,�l�u�1�z���H*�b�5�����f�����ܫ��^�J�7�n����f�=�\�N;��PΦ����1R=�/����xw�j;l�u�Y����
��>v\�Mw'![V���gGwBWH�Hp���u-4b�U��v~��CI��J{X��+j�sN���+r$^����^S"�Vo�-��}��=��Y��':��w&Aю;��ၮ6Lw�V�6�մ�Pr�*�aeQu�1�qJz�ma2Q��U�a�l����ui8��f�P*B��<�Od&�'�ay�Y2�����3����؊��NY�{Q(��i.������=&�@pQKzuȶ���Ю�EoR+X9|ԕ|� �g7�w�\�*��꾇_n�L;�)��Z:P}�Ԯ�Z1���}p�u�
�5s�����
�v�7 �Y��/8<��-���B��4F��*SZ���Vہo�C���G�q�*'���[�t;2s�:��E�b�"ݽ�/�틧����M������g�R�KN�$�Z�������KF<w�R�b8�����6�;Mՠ�����hwW<++�v�(�.�ݝ�#]yZ\������_�/q;�������
ء���!�9���Ͳ�̔0c��"�Zޘ�R�mwj=V�R�Ȋ��L��I��./�9���Ҳ�G�M��1�^.Wq�˹Cz�kP�)����w`H-3�lK�ډ��䮛��n�U��8��: 3lj��S��96���k�r��#m��� �1r�ؖ%D��$��挖1Q';����K��w7�;@�y6�a���@> �RB�]��n�ܜ��Lsr�5sa*+�+ޡ�r�ow��lIK�H)��/�O�'�r�O ���q
�ݝ�SSy<U��n�z�G^�P�g[���`i�V���tc���oU�,@V�YzF�ۈe��l=���s"�6���-Ь����tJ��y�#w��oBW�h����66}4Vb��C��^�to(Ne�{rG�5����r��c��$i��{ݥ�m9�pYL;h�@�Lٞ� ���0i�Dbꪸ��$&s0D&A.��i��@�[W�X�M�|*���a��c���'}��b뺱�t��,m�{��7�Q���.�(�݀�q��+���h*�H�3+m�Z�i8���kuخh�z�;�j&�c�D�|4r��H	�q�nf�-a��KM�3Z�Q�-udu����+����cޠ��;�u�����;pV�E��u�CZ���/�[���'��e[ȕ"kN+�{ņ5��Lt|4��vEu'j�W�ycbQ����m ���c�D�c=�qIVv*��`UN��YÓvz:Z��\��}���*̸�i�P�����N�ݾ�6���r��9����5�٣�2�}oh�ȧ�9��S��@V�V��d�Ɂ:n���B���N��Ba�>��I6!t5 ����X�֭�ݱWh�C׷yC�c�e��]n�&�Nˬ�H;���Y�m����wd�Ȁ(�]`^#ֳ��x����h��f�M�E7�h^�$�@����j��g���mX�W�E]S�Q�s�-�*9���;�[>h�k��]l������V�����݂*&
Η�Ħȝv��pN�93���`��a��\���z��P䝛���s�A��π��:��1�T;�be�m���XZ��qW��-C��m�P��,J�S��}�:d�م_)���0[�m���]NZ���Nnq� ���2n�@��o�����-�Q��{�}k��Ŝy:�S9݂�tm���DrJ5�`��e��<�\���2pHK�լ^]8�J�Ն��uu��YJ�۶�}�V���������sv��,�/���,���jc�THh�����7.���1��R�d�Z�r��:��,�L]{�c�8�B�)9rgw�i������!IQ���P󢖊��2�K���Q�;6��լ�����N'�P���^Z���^7]y����JIW1��]�lʊ֧�;
u����ݾa�;2�Z΍ޞ������NX���og�i�R��]k줋�3��=5��޴��Q�ۼ�؊ة��^��њ�vPń�5�Z7x�O�st�p�-G
L�L ŹSE�[��r�IX^>���[����5�8���b�9M�-��SX1V<�Xµ4��@��
{����L��8Z6־�ĥ|]d���]����S��ʑ�g'�����+ç�n�:�0�Oh(Z35�P�s��(�3�������H�µ�zg�u6V�ˡZ� ׎�
�z:�n�NS3����7V���/�xw@� .���ʜ��Ѳi��n�-u��v��+���'��aޗ'Ksd�x��X��A*�16��D���F2ǡ��x(j�3�>�Uӝq4�q8���e1�W���ap},o�B�8V쵎�
��W�%�e�ek��M�M̷5��Z�3�
�㘆�td
�Rn�ǥ�X 4�ge��m'o��y�����2���c����J��t�Y�B���<���+�ۘ�p_�;�g��r���J��A��w���F]%�t)R�$�@������{0,��X���s*e2��� �(��W]��q�^f��\�y[ق�Wn�L2����:7�-��D�B�G��vrC:ˢZKT��{|u��.�:�;]��X֔f��:�mM�/4b��j�Bnku
��8�;9��v�����sM�4�l
�*tio]\�˹'�k;:�(0gWM5�!��Q� D%f��{��Y����V�q;��c�����we^J��z��;��Ru�2�[�Y�������t\�\����+^�"���K
1�.��ZP ��Yܖ���VL]�or��]+8���y��b�qOm��2k�wV�o�V���aG�ұ����J6	U8�K��t��B�o�Fh��{Vӡ�0�y��m�,���GZ!�t�bB5���3շ���-v��!������e4���m�5�Œ�Y�KYC�!G��'3��w"x�p�t��f�:�o:��2�Ƌw��i����x@�#��Ӷ������M�>�M�ɥ�X�T�ݹd��a�|�4��o}���ꅍ9F&ժk���+���p�8I��Es�^�JJ�zs��֚F] ���b��Ǔ3�k5�H�=F2$Y�C�'��-�6d��ngWk�κ��	Ys�!8���O��M:�2�3�w6Y�~ܭxޡ����e-=�����f�6�T�L�ǅ3Φє�*�C/���)�J�ٰ�qf�3k�g�(���H>珗P�Ko	@:&5K�k�ϸ��~Aݾ���y��Υ�S��=�|�+��U�E��i���f�Z��À'��ƪƎ\[ȑ��3)up����=Z�Is�+���Q�B���l�x�R�tp���s�����=�i	����C���6��b��Ed.��U�v��*d��Db��5�Cwm6)�#.�b��d���5f�D���C2c�S�5��KUu�ո-R&�5[6rBК�(�;��eue �[0��..��_��D�T�H�*����go Y�^+�_� <]]Q��i�Eح����{82�_�e_K8��V~]�vsw2(ʽ�[7船w����|y=�$�7�-�wݎ�k�W;�v�A]�]IF���������9̬��.P���ۉ�
//��eFN������Dl�L)���:x�p�4*m
+R����oW����v�L@��d�>.|�Y���ST�T{Dx��G[�1ŗ�.�o����;u��(�uooSD��q�՝�v�`N���a���ޕ���Y��6t6`͛�=	���a.�s�d7�6gNNY�y�v����Ve���mg��;�ķ|�W�f��T#u�.ge���mXT�rR����W ���c9Z�����u:Ӵ8h�VL��pn��$�9��]]�j�m]+�:�q����6���\5p�r+[���&jC7y�J�2�r�{�̤d��@[�q��.�++a�=6��3�kK8$�����KW���K����6�8L�c��C�W� 7ƞ������R�(�T��ĖR�켒�h^������/�t�������3��1s�����>7�:ŀ�i�u������溸���S\�Ά�ܗY��Ǌ )_�#�3C��s��]����j!��	4bT�Y*:��]��[DV6tܭ�jc�E��\��spJ+f�AQ@t�8dCTɺR�[K{��n�"hN/%����G�*o}h������y��!�e�	:坯��Idޭ}�L���^<�7&��̱����s*vX�U��?��N��ĕ4�Ԩt��m\-l�i��]]�'f�\�5�L@�t�F��\%�N��_R�ٷ�[}��"�Yv���
&Up5�ϣ��ǃk�?��ρ
_7�wYBMK�]��S;�$y��Ƃ��Y��B����0��F�U®�T�f�<C�
UceK������9�
;�wJ��i�ȋ�E�3���80��'F4�NF��Ur�p��cAy��$*��D�罜).�t�B�Ͱ�pyp컥�5-��\�7����2�w+ig(�+3l"�����nQ�0ٗS�=A�Ee�nT{�/�s�m�i��n�s3i��v̥}lj�������:m�m�e,�2�����\�2�<�S��*Y��g�c#�I��|{ogf;n����и�V
����Et���u$ʾ�;iU�7�R�.��z� յ��s�c�@0���(uV�q��>YƑ�����f9W���YaRv��z�R�x_+�Bk�v��qgº�I�"�(��M�ל+MJ�{d	|U��Iv�ԸU�X;�ٶn��d�o� �5ǂjL'nLᲆ�w}v�=��z�:�ZƘAàq�d.���f;����`��,��ե����;J��90�U|�z��$�W�O�N��OUaV�m����,��c�t��6�0R}���s6����u���t,��R�.9��l�Ӌ�z��`u�U{��`AI�՛�=3�h�����n�E%F3�XĠ�}���Y9��,]�	�r�Cٱ̮^�W�xh���"����2t��z�AII �v���V�;6"'fd_rJ$���Rl�TY�<��q���M]��76]J���C��#���'�TV��޼[�3{�@��o?L�4֔g�V/R��A�G;������v�W.�����<�
ԡ�6l*�ˇP�zL�z2�}�g]ʝy-�ܸ�w_�m�nq�d��=�$�I;���I'uI$1���+npY���ur��塷�,1F���BTJ��-
i������k���uJW�e���Ym��4�ʋ��!Fr�ASk�-�n�٧	Y�O>�b'f�.x���q�G[u���Q�{e���Ր�\j^�̷i�ge�;�H>�OR4-ۦ��_�h
�<@�P�������hc!�*�L��J���t*�1�N�)�t�v�3|��^\7I��!	�V�x�i{dW)���;�˗�i��h_f#Ox
(��ZB֮�
��;/�����i$��
��(��QFɍ1ʹ�µݍ�`�6�+�Wו �,����N仝�����x�S�tf�V��ֱL�9פrnHQ3���2Wr�[j�R��	�Y��$a�Ւ��#{�K#�-j�V��]��n�񩮘��b�ۥXr� Հj�v��N��AV�De�{K��+ޅ��Cz��W]ӳ8�M��d�i	)�Ze�Yα�𭮠�e�a�:Z]=���
?e�9�g]�0��+\&ʒ��Z�|�������.��[.��H��-Wֆ�R�7h*r�#�4�r��SN�}�i�cX�5����y���-�)+����S�,�����8�ь�k%�I�΍[���Y��*"����"���&~FG�3�<��$8e�Ut�BV},��2�nf�$&2�S���;F�.U�-��"�=&�L30�l���s�DF��1�.��4a%H`������c���$;w.p�H��iw ��Kds#W���EuL�x�5�f vp$�v]��K�����6�u�Ra��ydv��2�r�:u���<ũ-�޶j�����Q�"%�:M�x`=.�lh���M�4�w��Kv����I7X��#:�c��^v�.CB	t�:�%��jV��t��ȍ�gy[S[`�4��:~1��I��z�3~���i���z�fd��F��{^ܬ��S7��F<8�ڴ�͙H�m�"<�U�0E��/\�YE0���������������w�ء{?�YY��D��f��}ySs��T�;nd���o+}�u�(ч5u;veu�Ol9�%�Z�7�l��u����U�T�n��!|��V�e$n�ϖ˒j�W�W��At
G�[�͢�M(�DC��4�Ӛ'�`\�B�<l��Y[ȴ͋�I�p�6�q6�l�N����+��;��e�bŤ��j�ucD��;Y���1J2��3SJ���gW]Kՙ��2�v�t#Y pT(��ʦ1Y;�������٫�dЦH��u�'�\A�]������TV9�� АÝ-K���h���)��l:�g^+wn�\�R۽��P	�I뼔�Y������]�� lB�7a]6��P,* ��Ѫ�Xw��F��h:�:��Ө����W+T)�����o[�J�+�&�ڻk	��Xx�>�z�S�w9澣��*߱r�ԏ8����^[�l�?f�sx����E@W;J�M���n�Zy�9��<��ޭ��у]9�X9�U���л���S��Q�<������AXXF]���<F��h ���"�v^�[]3SC��oR�4��:���V�����M���R`�Q5�B��Zvq���T�\D���r���;ѳ32�)0����Z�L���CBC���"��>�Ԧ=r-M���9����]G8��*Ԧ2��Ž�1Jq�oj����*ր�j�ݗ0�uo@#PH{R��ޫ��.�T键�����/��˻d�e������x����*��䷑"�K08n�+M�g[��]eE�d�1��m���{�/�`��AI���yM��v�ːN_�X�*w^R��Y&Z�%E�(b��-�7��عL�e�����=L�
���٩6捈V��������Z9l��tʎ�Cw[H�B�xp��v�9��X��ө��^��Ϭ=h��%�Q�[���K��M�O2����ͨ�;.��poR����nv�'B��u�$�
����8t��5��2�>WN�K�vR7��A�9N�\fÆ�t}ۋ���F��*����o@ �nT��[�ed/5�.���{wB��Y{�rZ�W!6|KL�o%�b�^�I|�@��bo��kt�1�(_g���Jx��Gr�E��*�`W��NI��m��b��غ�Z˭����Bn�N���M$�j.v:�'-��*�OY�q�e��9p�v��']y��(��Q�ߕ=u�wH�N��j�ƈ��2�+�Lm��mc��x�
�b¤a�.���\ݒ����?P��i���-�Ҏٝ��8(ni�S ���ِ�2��;� R.�@�kw;%$��^��m��Ȩ'/8�G������t�	�� VRm�Ev0]9]�:}�e�4����V
���$�.�[b�\V2��k$�ᢩJ��뗂��q�>��0��YR��:~���z.������W�l��[3(��t �h�n'��r�q����72�+y)l�w/� *�U\܉T1�)�xz� ������uv�_&�T�t5�؀;0rF� ��E��XL#SU/-�/��*���[{g��/r%%V8����r��"�Wv��W�bmo}��*�2}���Bg���k�U�p�5��_+�n\�f_V�5��J	�@��AR-�I�r��gQ�.�ܔ�mXe����8�3��T���vr�%�*�xX�ѽ\�cԫ��<:�����:<��tV�c�����<1M�A���Wz��j���Z$U\GyW�:*�T�e�۰J�M=���:BV�%�^��%��_`��A.��������k0M� =o��G��S;J��BG�60͎��C�^�a�<�B���w �Y|8���Ѭ8&��*Ϋ	d:��SV�|���<&���F^�^v��+���g����mEVp�U'L[踩܍��G8v�k3u�����k��9�'��ev��������S�"^]�T��-�!���+���o>�	`�V�f؀Ȍɻ�'kwq����u��qH֎�];����:�*p�h��ͫ�>k-�Ѻz�'���pC7��d�F΀W�+�KIp"��ls�b�s��֩���W��z:���J�nwD�%�ì�U��ǒ�d�mKβ�o5���i�5F��+�eXn�5�����c(eb���ΤE�Ƀ��ڡ�ᣰ�bЧùK�r�x�:����aV�h��0���4��6��A!�V橭S
��e��f����R�3���Yae�f/�52�m�1���:��esr�T�S��%���M���7�l��
�u]ǘ&��o%�G;�Kx�ylk���@f@[ݪL�Ҽ�XiU��w-��:�%+�:'\��L����� U�H֌��F����ڧL֓C%.׊�b��N��n`���6
2�,��w_:�i$��\�깃:��XMuq"U�tM�1� �+���$�Q��7�T���X��u�\���;�sN;ͼ�{P��sTz���V��N�[6���M��9�B�sl,��0�/�)��.���F�O�q�YײnN�b��yӠ�D�(��j��(ٶ��[�&��fú�	���[3'E�=bռ�(+����aɠf�m���n�U�T��N�Z�S+���2#j����̎��5�Y˝H�헪���).`�7@��V��p-Wcu�t�[`��J����w.�(bSi�%��y:ܡz�uө�s���e��z���"��Ap��g����.7n�c���0*<�:+�,6��� �d��S�n��������&��q�]>��ۿ�Ф.;
>����:Bք����LO+Mʇ��z9�� �[�`��k�s�X�/���N�d�t����9A%).������0a�燴���S�)��{�o`��WE�B�=�c�0K7fl��5V�2�k�o{;:��+-�T{��R=�� V����#�}���;oz�K4n<gq��*nfVd O��G-tG)}�u�J�(gc'^r��d��mLt{�Ҕ�����S�s�4	i��$�Ɖ�ެe�9#�pwm�ʧ�1�]A��� C��1ũ�/+�e��^��+���U���ܒ��+����� dp	eڼTR��2��,e3:�g��]��&^ř�wCS&b�)������*��;���wVۚD�۲�8]��㸴��b=�N���P�|�p�N�kQm]��z�������:YQ:m�jn���{��/�蔅;7��e��r�ÄT(*��5n�����,�L�*�y}�d����7E��{WcsD���P�W{&@�7N�s
_c�X�}�e�͒�1AArרvnU��*�"�bFk���׺n��rfg��ù���wZ:�K�&�b����qز���t���%A\��aM,�Ǵ��ǐ�eZR�1@��]�>D��ݒ��ڮ-��N!�ۻ�J��306�敕˩ۆVNV�'4Ν�/A�/7����E��8�(�sVގ3�mҐ��U�9�5Z+����ŏw��j-u����sbLC/^h{:�%Nc���;�//u�sΩ������ʮ�ȶ2� k��;kks��G�ȵu9��XmBf��8��
ʙ�s�-sJI-Wul�F�6�8�ܳ�Y}�mʻ����c�x[]2:W����J�8� ��o7�����Ԯ��5m�bVZ/Uc�,�	F&U�5��2i��[�S^�9]CA�a�cV�����ebDxGcyH~@c���*�J���J�-8q��륪}�;2vP���,DI4�7�bj�Jkk5ʎF�C�ʉ˾���
�+��cb�v푢����wDuR�r�N��W�m�[��m�.ތk����P�'jsӛ�n�L�q	5���kC�ܜ�`��u�W���;ܷ��m�����-V��H.�,��
�
]ln'�8h�k^NK�t{jYM��a�hN��㼫�U�|&�	�YG\<�@A�g6OJW\je�}�۪+�baČ;���Y�����\HE휅;�%ռ!���fdE	]QJ�nU�9���le���B�3�:K)�ͭ`�GX�e��
!w�Yo�0V��]J�G�+��� �v���9;\�6w�^�XOy�.�n�E���G�kV¡�f*B�M	�ZX]��s嶮�n����%"�}7Lԏ��vŉ�H�ޑ����>l(4��v�Wv�oNٕ՚�lv��Iv�[ڜ&�u�c���RG�wJ��>��E+jE��[�T;X:X�#���[ֹ��$(���nj�p�ˈ���X�e�Cd�K^sVWbٮ�Y�����{��*��ZL�����#�1w&+�WZ����$F�p#;)N��^,��UqW�vz��ͭ>U�cT�м3���:���K��>�3��H��/e��d	��V����/u4��@��N�7*㻬_�i���&0!�h���o2�W4"�i�J`NuD�K�9�Ԍ���ϯ-u�2�3]*{6��r�9�iNb��^s���l���y22��+�������ibFVe�\�=�GD�����j�s��]>����M��0c���[WE-ν
8�O��+��m��%�Rqvi\R(�}��_\�d�����9��F)�{u�vW��Dj܇tk�ڞ���y]�z0�[��>8*��U���)[�Nzݳqu�Ȫ�#ܪ�|���댞�Wj�}n���cFCA����K����b�EȞ;`����z��e	*`g*��%L�d6�e�S�=u�_+���Tɑ,�.pE� ^�x@7B���q�d��hu���J�:e5��[j!�Z�$���I4�����]9��^-�����v$�Kfgbo���u�4=�'km���h|�탢�bt.Jq�QUH�U�3^Ί�ko+.WJ��ـin���yozE�9�������t��6ƫ��W5���#׍�к+�4�]�j�(�QE)pv.1��(1Ҵl�Wp�Sotc����7HX�YH�Y�ʻ�	F�{�S�}�!�;��� $�]J�&�c�VZ�À��q��=�vL�K�}�t�x�<&�^u�[x]�/7��TTt�rs��X]s��,<;�IY���M��[n^�	�/�$��Hu������-X7�<�Ibd��vo:�[���u�0�C���f��l����KM��ѣ�]�;
驫��U��.�������`�c�W���I��᳖ p{O)-ZU���m�>�v��yE5����Q���Q.b��G2;�Z|4��ͦ�nI��X\㎡�+��Ye�;]����څ�eb�2M�|u���N2`ێ������V���7�,I��t{/�s�.�sO��+�
T(�K��W9]I�g�̜��G��h�4�����j|�TԜ7���o+o6���CZ%�mV���5<�����f��.�l�Dr�L��N[Lefb]�I���Kg ��wb`����R��muM����+>=��k(<���/����������<�����_�?� B ����&@����J02����2?)��vO�ʱ^�U�r��;&����<2[��g&��� ޼��q/U�n%c�x��y���x��K�@��n��������I�oo���5�o��yP�7s�xF���:hA���*Us����n����f�	})�yk��ܕ7�j�"z���y���K3H�3t�z�(���x씱F ����ѹ����uvJ�s
��q�����y]�����3��4\tFX[��0�0^�QݓD=wrU��p�涴S�~�=]�-�[����W7 �+��@������3e9W*��vNUp�L;yLKM!}�k3��V�h��6;1S���
��S�cGd���G+(���B��HA�F�;����Y�J��%m�+�M�yӊ�N���۱&t���#�{.⃷�N����Wc����4:H�{J�r���W��dE
)gˎu1bu�:��<�O�!��f-(�/��V�Y�[YE}��}q[ࢵ��SӢ�W��W.�@�o+,-���h>�ig��\�Ѹ� �_r���ˮ~�a�#�M�p�w�%��Vu��罨�W�
t��X��/����[x�7����*ہ��8/N���{�X.��{X����3�\�u�x*N��#��p����";T:=�n�5o���q�{ڏv�m�mw)ܳ4l� a�қ9!�DL�T�t��(�O�{�7���Yﺪ(�(��PYJQm����k`,���VcF�l�,mV�Dq�fJ�b�jJ�U�!Q�UHF�R�Bb �b4�M$�P
��HV*5Qd��q����=J�kY�XVM���UF��LeA2�u���
��d*����$PLaMP���(���[�Q�XAaTY$+R�)�c%`�QIPd*AHi���10d�֢�E�YR �R��*E-�`
EX$�$� U��X,
z�[�d^���Cwrm�K���@靭�j�ZGN�멃��l�/^p=Qţ9�%�����m�[�L��a >+��)Χw+{���A|1��o��x�՝X��vX���5-� .Ү������ �u�4p�;=��|�ce��-g^�����Q�Z&J�
v�1���M�Ujv����w� �����������N��'c�݃�kx��Uz�^Δ�Q��S��;����ml��n##���a {ƫ4����䦘�ja�����u 9��}H+��~�݌<F�1]�������Ő�U*�����6�O��ێ����q�s��^�rNA���"��Nti�)�<=���Pȉ���#��S���0����2Yg��7���6!���Qf��� g*���(�t�Gd�8��Eu�3}��ҽ^$z�&����U�H��=��_C��@�>�Xd��!��vR�Έ�["k��`gb2��{����i}�}e�0���,����Գ5�0��չ[]���-�&��Cb�[�14z���h��@�Fnӽ?�a��]��������G���c )N�0�+.^���ʵ�szm]��Wc��`\W;��Mo-�f�J����
M�w颞l�{	l*��QNKp�!]�ګ�A]y櫝b�Ⱥ��E��.�>X2}⎜8�2���$�'�o=E�fo�U�5/�������ӥ���'F��5a׶C�æ!�����#P�s����Jo�XE�*ܮ��4z��J����lŸDY��±#wo'8=�$����KKmJ64/yWXk|]ic�wW6e�Ck��H�V�Ҝx��f�yP�CM`W�&�I�A���V��?q��}��y��oݮ�d�{��}�w�dc�
h)�0Q�Ϥ���2�����PQ�;�Y��ҹ�� Yo��}�X�a����,�"�e(�X�����������1r�J���1<�m��l�p�aF���6<���. ���:�R�ôԣ��4�.D�f�d��XΞ6n�7A;��zr���*��|����r,��N���,A7�!�jQ�c��@�fb�^�9qh���?���
�ȼ91N�%���R!"����|�K�\8%]%q�!]��������wt�z�7���,A�|�\�����;��,n��(ܽM�7�#4��E�q]�l����\���Y�	q�Ԡ�y�O�	E��,wQ�
�wo����4�T2�L��LP�{U^�Mc��S�28�?���:�4r��S����,.��p�P#i�Y;�9�g�� JsS}��Q���b�#c�2�")WE���u����=&��^%�<[;�O�
_/���?���S0`�*�xm�Qc%�Q���o�K}�'֘��h:|sȅ��
�u@��t�W��V&�Y~��N1��r�v�uJ�M��u-�*��@�T���Rܨ�j. =�@�����7|W�=/bG�}|�bG�17,����ݍ�8hl#������K��F�W@��7s&7X�'d�Bpp�+[f3Ls��k�*�¯<���t��>��p�3��b���Ӗ��Lh!�Ʒ�ſ����A�?>8,n��g��C�d��o��m�?^��)T�7�V��<sce��#o�"��kdv\��GqA��.^��؜���qnF��N�Ó�`�"���J���S�X�_�įGݳ�N�����|4���h�{��xv�5���3g'��[�pU֦P�����ţ��1wch�S+"��W��i�yrf����*^��p�E�+e�C6�Tr�*�N�k�
 ���`oV��2��s�`����6/ִ�ʦ�|*qxz}�η������PԪvo�b69l�}=y�]$��
,�u>�H�����qB(�#�k��[unf��|M�!d���y�_!��AA���%�Ж�"D^�>��8S�Î9����ck�����DԷ�̓����,��5�S���*Ea�j��R<03��3�iWXj�[��̣R����(��|!>hw�.j���゠P��:�/G��y��P�Yݫ�r�f�p(��3���V�2E�}�1���e�n��3�rnI�\�]Nq)ۜ�&�N��?d{�m<�y?�t8;��;��)����>.E�+\��Z/���qA� 5U��C��k�*�,�Ч����Ր'��%�[�)� ��n(#�i�9E���j*�~b���U��X���Ť�Ԇ���#؈���On-����d��+�l��2����>�I͜,](��YWRZ�N�S��>�f�=uD2��J_F�"^��p�orW��0���uK!���+�wd2��qr����N1�vpX��Ȅ�s�4�Q%Nv�עM�-�I���f�WӽM���!�+U_NY�b�ǖv�.r�W#3��ER���H�����&�ݼE�󰖩�-	*��_h�|�*4�Vc�2,O[�o2��纽X1�5Cw4q���H��j:*��{9�,X�T�WP�1X/�uz�����8�F߄AfB�p�f%�)yu�{C�=�~�@Zy��<L�.^�4��0��ͦOJ�'�Y����߂�qIO�Gp3��M����n��\��! ����iB11`��.��G�i�6:�t,���_C������ࣅ�H�\q�w��d�Z5�����c�i|��P���ME��P��SǊ����ͨm��7�#"K�ƴ�'Y)@�5�Eh�vc\#b�EtX�"���"��
�,o]}�_/*��י�q��'q�1VDA9d
�2�]Mnr��U4Ňcǽ�ٕZ��#wɆ��^F��.���������g ,�aR�*�HdW�ۆv" �N�Ξ�m~ڨΊ)���U��O�%�*4Ҕ힇���ӘB�D-SB��{f�t��q2���.���g3-WN���aYo�<�#��pt�C�������n��OL���̜m��͋"q�ʴ�B�j�F��b�����X�f�}JCsTj�"�|t�t����kkj�W_W,5����X4�Μ[R�5
Rtd��w��:P�������]�Q�v6�c���^x���t].-)u�3�egH�sj�WÈƕ�u��V;�J��H_����w >�}�f	��Ϳ9RV��=\P9�->���k)��S��:�ʫ��Iu�b�C�������}�P�KU�y���֊cg�#]d��@�c�jY���2�$N�\�w5�?Wv��ѭ�-�d_o�r�3Е�'�:r%�0��ؚ�/�AZp�#č��l��x��d��$�>�3\��9Kx��ݯ�
�gw��Ř�Y{�w�7Һ7�U�
��#�n����i�D��<�v[�!Kt�
oo�+"�]!�ҋ#��	ñ�eRT������\��ԩ�ؗ�A'7(&:���l��5���l�R�����*x�W�v���r�XY�bFd
�ެܱ^���_�n룷�5FR���h:�t�1O��u�5j��Ԛ�;C��=ܩN�ީ�Qu��
�I(���I�(����܁���.��O;�ܜxS6\}�3j�N��(�o�i\�w(^@Uv2d�G�ػ[��qD�ۖE+j'3q�F�����M�v�N��eH��n�G�nm⓾�X�@X�7���X�C�P�ΫK����0R6Q�F�!��괦�#u�b&�)=��|�4T�]B5�\%�le�I�lz�\L[r$��h�*GS��b��$ib`[�"J��k!����<p���'~G^��{^T��r#u�X����X@��5�u��q2c���|�4���mw��[�.-:]�Z'��8G�7�>^��F���25b�5�����S#ƹ�����������S�;��ә�3��� *����|��;Ҕ���:DY�W�XѻÚ蚻��Z��s`2$�Y�iY�����R�VV
��؎{5Q�NT����Qp5�0�|ً�xlP���S�&'Ցu�鸚�=g8����>�^��>7}��&� ���R�XZ�*�1N{cMU�""��/!��q��ڍ3��dן���N��<�s8~����������ì ��Ua�A�}�'zp�i�w�el�}n�y;��!+�(�]�3�v��sfTͣ�#����xu]�ڶ݌�)��ΐo-q��g^bsGj�����}��zҹ��}1_T�%�Ղ���n+~O&�f������S��O�W�����;�Iy̧����^������N������u�L��os�*P��Z'��wNg�����J8]�S�׺�-W�����c��0���ָP8|�TN�]3<V;�P�2���^���٣暯(r�3yW7���q�
'���ȰD�<���dE!M�^��ui�\r�JqŸe���ӳ����]#vzI[ѻ�uv��9pn�N�g�ۛس;�BnE�\G�]��u�:a�0�6�ޔ:�[��e;WQ�{I��4/Ӳ�WS�[�n�.�n���P�5�S�q�s�s�/3�g�j�r��
���aā+D�S��]�����)۾���;P�j��.�7����O0Fr<x���@� ',�o�.���p�1���&�v�3H[槍�w>��8�9���q��c�X��Ϛ�<��0�H8+>��wQRqV���Z�22(s��]��
*�8f��li֙"��T��3b��<3��,|��K�3X��^*Sѫ� ��M�	�c��ǜ�Ei77�eX���WekrL���:�ʕ���ΠL\�ho�׷S�cU�=N��f�Օ|���B8�Ѩ�T�\eEEgMu�Q��&�c�U[=��Mv6�n�늢}kR���]�+ ��C^s�����6��"Ga]�r�5�r���'�1���s��Qt9'��N�Uzݢ�w8(��'A��O��[�I!(L#yQ�=�w�֙;P��0=�`�"Gr�0��nv�M��Z����`DH�fG#
��P0�ʫ/a�a��D�l�`�;3S�,ozL���39�6ǫ�&��#�C�'X�E���Y>��Ӭ:X0�t��q��#3�L�-ş���͊�6fyi�Ѱ�b��|i�#a�����@���+v�fI�b�Gk~��,nCQZ���x`߽��_�gÞ���W�,X���i��[�lQѝ�/f�gI:o!�D3
4$�]�NƝ��lw�1T]i����+�[�e�k(��=�R�" �炋qIO����8�FDr;�[E@�����lY5�V?GW���t	��t��>�Zt����Y����.�+G�wzpd��:�"�7�b��3�S(�S�h��>��l�2��8x�D3�;�}�4MG>�#�Q� ڝ2�h�\8G`�p��ˣ�Mȸ���3V>��N��5e{�U�.��D� *u�n, �[$����.���zP�	Gt�IK��bg1'�rQ���3����0i@�5�(��(����zg�ʛ~A�q��͡�&�;/{��X�<y`���@(��`��'�\A=�*���\7"�{�ɽ^.��6��K�� ��_7���Y�]f|�xzP�k=`=��g$�RU��Ȋ��	�y��qfA���eVSX*㍑;����J�I�%��>��Yf����wJ7�i�u����)lI��Q��:��-U��h�|������:�(��Ɲ�&gO!"��~��Ϯh�:�MVPF���)��4���'�=�%Al�	���d�榀�|���^��h�Ʀ����yk����gŨ+��2V@
2��^�=w����̊~!�ek�'�R2!≳5�Q�OH�:l���1:�p��-5Q�3��٢�C��-�*c|�+�0�u���,׆�w����'��o��^���El98BM����@�Q r�;[<���{2g�{�?�DA���x�+���XkΜ��^�+��z�� u�:#��
���)o[8�;w�h�w���M��۟>��P˾D���:�;"�#��N�ѶJ�YyS1��,m�+�X���ޥ��&���i�ӧG�N���jK���˥]��cg�i�C�/nQ�lCg�w�SH�Gj�x���v�����lW%yw$Ou�|bX��)��P�P�Y����d}�I��캍��A
�G�k�g���jE��tx��W�p<�Y����)*�٘�hK2r�ז�V�������]F�>p��n�i3� m.�}#S�wm껥CD4�7}J,��+���B��8	2q�o��p���n�Ԡ
���h�&K�B޵K���f�.�f�d32E�&�����K�vAr��32�]�	��o8p�Zk��nP�%����'�շo_7ٛ����B6q�'�^���ϥ�*|���Jͼ<V�˛]M�`^�	�|�˾y��:�v��X,�5�q$�����}uv�Z0���]/l���@k�*�;}�*��U�r�P��6c5�-��6:)f�y����Q��(^Ed;{,h����н�z
�]�]���雾�y>V�mt�z��@���5��%nFC�6.�7W� *�����ۊ��	:.%𝎲��,N�����_�޶��І8��ِUd�v0$�ED�Ż�?����p<jj�{{�辈Dʹ;r
Xge�5NI^�����{���V�`r�;L.ѵ�wb	�;��ܮ���lո��l�F!<_f*���6F�&)�
厡�Igl��7��:-�e�4�:ݪ^�rv�C���X��,RR��g�����a���^ۏ9�w�U͹���Q8�Y���2�9|��ͣ��U����f����Aze�#Upe�2C6�_Y��Ʌ־�iΡe#[��h�2.����;����a�O;��<
�К�ݱ���o~�����,�4B!O7���7Ϣ6�iA���i����>�~�� u�r.�`�N��a�N�����ݧ��d�H�CMn��G#��9S/^E�Ö�HN��%�]v�u���'��l�/6�������f}tB�e�|����y��ۼ��R.�;[��r���ǻX�`��7�t�N��jֱ�wO~!��5Zc�j��.��T�AuE��D��o:�H�:2�#f��\r�.���u�i9v��z����-vq�Ty�6��R��/E���h�Xl�_޸@z� *���
��*ȤRbVI��(�Y"�0�PH*�
E�)H�AADd+*�d� ,��,"�(j�a���T�Aq
�YbT���""�P%Aa�dY �X�EXA`�E XH,ST-��EUa$Y"�`#
���iQTc$PQT&�*H�%B��)�T��PPQE��(�V�F)���°X�UY1+��TL@����)b��CU�X�(�EF)"����
¡Y
��)���9}=7����>_}[Z��9��0�ei��ƥk���XG�u�1=~����n�TO8�]���ò�7ߪVi�99mHƏ;۠���t5k�V�eZ�J�SWi˪�eP�fRt��2/{O�>�9�G��(�s{~1�zQ����8߂�/諡��J1ٹ�mmi�����u���񍏳��݆�bٓ`���}[#�wU��U
f�5{��~��S��9�R=���G�/���
�3���p�	����V(rg{2���bԽs�7��[����C�PƩl,�G���I����ܢF'��<�Z��&�>�	ʄ`���X��\E��N	u�P=�W{CS����V�Ha�A�5��I��D3'}�O�i��ڑc:x�]:[����<�jY�=�d���N#��-�0�9��0�B��u�*�>gTi�F�q}��=��ü�Y�jg��n�N.M�۽���8��DX�MF�ό���E���,)�:���������3_	�lLp��j����������JS�dA9	�� ����zEλf�vUJ�Z`Ծc�{�]����J���}Ѷ���T �7����@_A�\^� ��_�^�ps��
����\@��v�5���?���I����آ3v�1��v��i&��b��'C{��ҷd�������x�߮�����i\Qtx�w����Th�d�ɯ{���\�UV/�lᢂ�yNi�A��UnYHVa�J��n�J�8<O+��-(裏� 'q�|׆�L��a�
+u
*��P_cU������9���:uf�|[r��P
~�Gx���mzV|=s귂tƅ�Y �OZ�o��v�ʼ�O^�UW��e�)�c�S�s�����]f|�1�yZB���CT�6�N�ǻ:9�\��}κ�ٱϝ��eoT�����
�8��؁/&�z��s���\��Ow��/�ğ�豱��՟HIW�)j��)������P�_ܴV4�Ь���dթC����Gk|HP�53
�t��JI�IJp�7�`��t͋��+r&lp��uvQ�:]�%�0Sr7íW�v#PN��E�K��T�v��:���u&���&�*��i�ɀx��d)�u��#v wB4ܷӁB(���4̘�]�d�IfS�g��_�3A3Yx#i�io8��3v�����Xk�r��N숕�)�me��b�D�;u���}]Gx>��F-*M�o��-�K+bUH��!�t�2Y1$_ml��f�Y�HJ�Y�uEy����͛;3S�[g����c"������\�uϰ(<���'Tz��"4�Nz[��"��*B�+��U����j�E�i�:�P �r��]~g�3'c	�
8Z�]p� H9\�ͷ����e��˗�Ž�A����Q�rx�;}.���:�%�N���S��p�=�!Tn����QE8e�P)y:�$P�g�Bci�GVP�)dM�aͤ�2&a~��lm�6F�z�ħ6��D�<�P(�L�=!+1*[�uv,v;�`lV��n,U�󨞑��I��dh!��`��E_fC]L�w�l���}����(W_���/b������>�6)	[ Na'^臎e6ߨ�={�GUNM/w����꼰�W>5�Տ�o�֝aUp�k���U'7q�x�Xli��_tcފ�[�akG�F� �L�DY�r�ZtD������ڙl�؟"��#�(sʳa����bb��mA��9����x4������K/���;U�I^l��];���H�C�>�cj��y�B�A+wB�X�U�q͚����Y��\ȁ�''��d�䂑ξ���._\R��
�i�W��uЍ�����Lhߤ�KkMżŬ0J��(�����(�u��:��
��Ӆ�D'����v��Ӱ�aنF�b잍d�[u��"��8��;`1= O�,�7H�fJnmE����Jx����|\�n�nA��k@�?{E�]�,�)��h�1p�oϼ�c;���(?~o�x��g��ʼ���|�j��[}aE�;�:aSv͚��!��6B얢�� r�peT�V7���͕L`��N�)(ޭ�=��4�q�L�Ah\#�<��#����Y"61����#��'��
����iH���S����"	���;�#�9C��ĺ��Rp�U���5��ջ-Ŝ!TNC)��_��덆t��T�J�3�w(�j�=�F	A�W�y�l���c��8��-��Ti�t�2^̓荸�P��;�4��P��#��tIʏ[�#�FQ9#%8�y͞����!�v��Z��ԧ2���lE���ئll�؊�>�h��IZ������Cj���X0o����G����6�|jWC�:��VZ���養nV5p�[���SW@WڨnN�܎�3^f����:�^v<��K���^l��n���@�.n_s��J���.;�s�M�qT'�i䔭NQ���O6Lq��:��>�r8ׄr��Xzh�,������^��PW]�<�t�(=��}�r?>p/#�2�*܎�FֺR�qT()���W�`�j�]{���]d�8�vl��}��Um^�4P"F�@϶(��*cBܡM5 �w:uYy��w-����q���ᔭX��5W(>��S�ӥ���%�˘��=朾�u1؇1k��RFǬ�����}'E����4Uj��Ӷ���gLf���̈́G�V�m����;��uΔkݎ�>N0B�Y5Yt'�Z�k�{,��u3f��t7֘4�1�`�8�5Ԏ�	�k�����x���Ѩ9�ܔ��ET=��N|��J��om��K���-p�:+P�'�nX�ΰ���I*7a�O��Sq}�#k����^��R�[�u�َ�Ph�E��*n�a��=�}O���(�=WVzۡV��gл;�|tW:ӏD��8~���?��0��b�� U=?�B�Nu9��nN���t�u���ۜ;mҸuEAKU+i�<���.r�`�0���'!&��q��%��1���XVeY1��˅(��,^��FF�[���yU�ҘZ��C(���<sk.k����v2zz�D�S<��@G��4��	�����'i���R/����imyב�5)IyY���f��s ����B�A���6"Ψ�C\�C�y�	�����4"Sթ�l�s�A��8v1�B�BQ�5������\���;��&z�z��y��E%��x�Q��;�xҎ�< ���y�[*��F�w�(�آ��݌����4M���\�Q!�ʓA)�dIn+�@s�iYtx�(sG�L����*�B�,%��-���N)`�ˁ@\��z2%���nP4
;f����W���wyU�%�S��޼j珷��>Xq�SX7Lqg�]b���Wث�QV��ƫ_����G�+�'� fo'����Ob��-���Y��L���J������Z[4ګ�OϰV�ju+OX�M�^�Ve־z��>u���"�J�Y��1ޟ[�\� ��j�\h���K�/���>\��O�	��j�g���1�������A�({9�F7u��ûw�K�lL�w$�]�GAε�\yU�V��vҋ{+"��X��q�m�>����P|b�����ų�
�ݗ�0k6`�ۓu�K����r�R�BOJ�yR�i�f�����P2�zS�:e.�K��N�o/Uz�0���8]�՟HIW�9Y�r�*m��1�x���0���e8Ռ<�������l�3JGP���r��p�<wڭ]8a܋IT�ћb���<W.���
GrJ��,��1"�r2��)Ed-.Gpn�8GtH��x��n��MҶ���.yL7R	ΰ��܈��a����>�H���n���P�7,�We���ڝ���,F%�|k�a�y7���@��Q���p��&#Tz��(�8r���-gwW/#�9��KQ`6���NؤS�P,t�
��^�����qhlr��ʥ����<\)[�*�F�]S��m��/ ��*�tf��F+�:ԇ}�D"���ݴ�xP8*�0W���k5�J�F�0˸��U�,�9�RsfHۆ}ڥ�7ko�S�^����:>�S숌g�0�{,���E\��J�L:����A˾���^w�bb��>�JG �+��Y8S��ON*�'j�0<n�=�½�4A��m��n>���B�ɸ���p��k��z��t�K�}�.�9�2�6��&B�v�V��Fն鿸u�cߦ_�۵.�=��~\vQ�W{�l�i�
l,��)[���"�0�e9؇��o9Z�E`+�XGj�s����0i���*�yn����ڷ=�%qb�����c��k+O���\"$W_�PgH��1��:����(J|��AG�XeU���U�o��tȷ��S�S�9Ɏ6 ������_t.�χ\��%���<z�5�W_p1#�Yf��ϖ�Tw��i�
��y0��K��-]-�\*K�췕t)��Rmc�����~,��ȟa@Ռ���h�rC�&�L��WGV�S��-��':�13G�3�4��A�>��E���T.��NƝ��OIZ(�.�%�x��O{9h�z�+��<��gAQkURf~^��PC������O�V¬�wW7����M����t(��G&0���ePGԜ�]r����b���
�h���?)�6�~�])B� v=���Y�>����5g4EmE��q������\x��.Q��6�cuf�@�B9�Q��p���]���fNf�!����3B�t�S�+��k��S����Y�C�"��v�\!8x�r9;|�T����i$�dW�츕1�V��%?U��c���AQ���L�V5�l���ݮ�����M���Θω����Gj��[|l��k��d�/��2׽�\[�����v��:B��[,���A��z�]*�Twx4�H�x5�ή�k,�P��vC��e����c�[�أ�������ًgn���;����	����F��:eޔ'�����3�ur�q�n�a�,�Q���Y��9I���K�aNvhi�6)����؊q��Fq�ݺ�Q���UXN���+�,����BV�6b���:�jJ�zX;�@�||u|qc�����*�y�KnlFW�ڴ����>�S�*��`��T��*�}����Q���u���˴�/������X���͆��E'` dmHQ��Lj��LSR	��*�B�
'U�胶i�
6#\Y�ٲ��a
�̚p���QcT��n��}�'������;��չKiԙ��s�z�H��Y���N"}kE/����x�4T�j��U[�]s{ZR�������;ʝ�8���U����w+�!q�p8ٱ��y���`|zr���1��i8u���l������s�7�X�t͙9�,�;%i;u�HN3�x�7e ��v����W�V���>�\Ŕ����.y��,�Ϻ�\�ɶr�r�E�p5��m\z��+$Zz9bjS5��9�e$����1�{y�sV����2
�����'�|�x�c3��&7�κ��fv4�1�V���}�O��iZ9-����H�ʩ4Y�8��o;��<\��P���h���(c��r��m%H͎u�jWBA�isg�U�J�<�Z����� R-º����
�υ:���㢹֜z%��#���Q1�5�� FR�j����Ti��d
=3����mH����0��t��k)�8m���:sȴ�/�{^T^Y>B�K!�Q� aU�9�Y�t����n��F�ڼ��'�l��6�;�>V�J�;^5�o���d�x�1U"
������FGy����g�+^��C��Ϋgܘ��e�#P�t���ynק͸���s�w�0�}��={�&���"
qAG)�lqd1��ѾR�����f�w��=�D��˩od�Q�g<p�u�Ȕ��@׈�&M{�VĨ����0���Ҧ�Z�4j��Ol�=�H��N�3�����6ի�	F�#x����$o[Y��oҫp����Qs�b�75hm!��qg$5ظ!ô;sd��őp�W].����܅���s��S��Py�l���D�)%��գE�a���%�ifL�(E�p�Eh���@�7� �]���뎯,�%��V���x�Qi��[�
�hQ���+�Z���Ԡ�|�^�ɼ��/Sk-<[:���V��:����8��e7s����8fX�`��6��T+�Uʩt^9��es�ܣ��t-��=*(�\����ٔ�t�K[ܢ2�S4��j3zk�]�ۭ'[CrKEbT8�8�m���1��y˯��t �ˈ�mء���3K�y��WN��fJ�
R��'\w��!�F,��Ԥxt���L���i�����+�r�a^����8ǲ��
��qf7�4�ڑ��"�2�=�#z5#�$!��_Ď����
�jK�V"����ہ���ݙ�Vr}��V�{�R�+[w���7�&?�H�c;75��N�U�,�촍ʉm��8:P�wr�Ʀsw����n�	�3����k�4ɡ���z��S[z��F��fM���lg��q���rm����de��]�Y�zr���
��H��e�J	��w�2�M������n2���,<H�V�����6sH���}C@����*���hݒ�;����2vA6���wo+kV-ɜ�Zk>G�}ZP7ڦ��G*��h�C*aVQ�ٚ�y0��]u1�i����׹3�@p�$���@&YI(�qm��^A���f���𬩹�l�H��8
Ǻ0�5����w:��	���t妅r�Kt.;����8��:����Iw��$S�i'w)1�f��=������q��8"�x��0fvX�V���q�`1���\C�+���6�u���7�dpE���q�kP���@�LYl]5v��7K�A�2q�˽n�
��WO	��26�a+BWm�Z3��ing�N�-������a��I��0ۘ[r�%7��0[���
V^���;�̘��A�k��Ϟ0�u���p �,��n�3x���y�+��w�V����mve^:���S�^E�IY[3��5���&�na
�i�I@��WyJ�
n���s�ky(�!	۳);���;쩺�c��^U�kxܬ��&c��^cSi˖��r���l��n�jv[�A"�J�u�%���:�w�}��)u�@�yQ�
�n��EZ�λ(�2��q�)�j�6ÈmyK\~ �W�@A�Xp'���G *����uܛx�[;;��z๛�L�R� D��C*�w>��S뜱HnV��}��9�rՓ �4�����*���i.���u��>�ߝ�������?"�*�D�"Ȥ��p&�J�eB���b�B�ʘ�P��"�J��"��R�TY$� VAb�X,���+��a�� �Y!X�aR
J�L*�2Aa!RE	���$�* ,��V(
�R�&��� �X�Yf�V�l�d+
��H�2P+$�$+ X�%CV@�"�$�P�	���i��T��h�VP(�-H>�DG�/�g�OW嵐��ne��b�Ss�՜o��7_%Gw�/�z��.m*Lb��仛���̴�[||�]��r��=���*�u���\I΍��\����i�=I^{`b|n�iXq�l=a���Y������H,�Or�bԂ�x~�i�Z�^ٷI�0����h�������v���eE ���a�m����s�����/ʹ+�Y?'-�g�L@QN�C�g<�bn���N��/R~߹6����q��bg��=IQVʟ���쉾��}�;�}�$z�Q���Q�Xc�>ԜO_:_�ԟ�d�QI���g�1Ě��w
�_P*��h/�4���nj���8��bM%EIY����I� �~��r��,f�'�� ��>@���>GҌ�٤u�\��n~d�?!S�;��6�Xxw�چө>v���
ϙ+���]�4CL��^'�̞&�H/�<�AՇS�4��痻�Ѿ�ϿW_����������,�N�1�ϝM����OP��2�ϙ1:�P�ڐS�4��Ó���&$��>�M��s���~ޡ�a󟯶&}�|���F�B9O`��k�������2�?0�b(xũ��@�=Ak57I뤂ϙ��u6Ì��>k1�|�~9`c�N����0��ɿy�7<f�d��;q'�vǽ$}4�q�'(�ߔo�X?dI�9��톘|°�t���T
βoZ�U����LI�+�/,+�a���k�N�]$��x���8�Y�,�ͤ�Ĝ�����|��uK�w��A���E$�0~'���8�a�xsxE�g��}l�N!X�q��J��7��J�d�8�1E�0�ӻ���'�y�8��c�g���d��I>��}u޿5��3�Gk�h���}Gރgޏ�>��|�]��5
�E �3ü���&���rκHyl�
y�� (��r��$�I_�>C��m�@�T��f�d��������k�W/�g:rm��I�&0�!P�J��O<�0��C�s��h���J������Ag���E
Ũ��z��:����`v�Y��C��̨�٪�0�1���������ʉ��·�O�7˰��*�k��Q��:ڍt
P��4A{R��1�RmՂsJX�]�h���v��G�[l=�|��3�|g���"#x�]Ĥ/{,u]r�(��&�u]En�k&Ez�s��u'l��Xn��%W��u1X�w��gY����9��$�m���W��ơ���i�vɌ�{q��Y��O4Rz�I�+�s}�@x�����~�z����=�(
�A�����'�6�t�}E�|	?Y�	��Ą�쭇�t;�N'��4���̡��f�x����"�X|�`~�q�Y����%g��u$���,�lRVa�� |�Q��]����Ϯ��w�"W�� ���!���%I��t�~d���t�§̝��?2VVJ�a���h�c%zé�����a�q�C�R�q~̚@Q`ro�v:��{��������|�ǋ6�
�hT��`|a�1=g��j`x�O5��T�Y1M���¾'1�7g�4���h~��l+
��j~�w�!Y�J��a�QH,�d���-I�޼���s�v]��}��z�a�����4� �=��0�?3L*()VLa����ɤ��'��t���@��=-����La�TR~B��P��ͤ��I�7=�u�i�f�ٷ��w�����7�?{��8T<~J�Y�|� (�'N�Y*N!]OsRq<�!P�s���d�m�OwL�ɬ���fb�Y���M���Ci�5���8��0?5�Y��~��]}�~Vߎ����}�i�@Q@��;��=a����8½b���z}M08�u��ٶJ���{̓��l�'y���ɧ�w����XT�&�t���%~f�f6�O����:湻�t>�jfg�����LE�٫���r�I��OZ�ճ��Vb�'�Vu�&���� �0�M�̟�m��Xw��}d����,?0�&�3a�tOP,�Dz( ������ϕ���g���P�s���}�+>a���
�ZAkX~d�(q�P�I_�
��Ff`z��.3�La�*)�
�a����6�_y��S�Y�
����]��y�ӝ�ٯ���>ڏzO���RT+3�>�!��!Ri=9M>>�c�W�P�;J�Y�}�iEXm
�*O���q1��^���N�M!ĕ�d�Y�y���}����+\�>ء��E������6����}�a?�/-vk���詃n� ��`Ѳ�9>�f��y�;�[9�*��Ҭ��D�ws՜�>��ʷ���9���s��&���U��j޹�˵WNA
r0F]�$f{7��zEE�i����I�O�ͤ�(bA}{�&��?0���v��Y�~O��M������|�q
�d��RV��k:Ç�ᱜd��N2wVq���l�D�\�ҳ����Y���q����1��T�'���^$|�_';�I�x�Y����+�&"ɾk&��,9����Hn���eAf�0��*O��i �a�xg/�~�����ַ罛�4�|���Nn�ğ��O�=@��I�G����XO���M�~`k���1f�s |�k�G� ���OK���3z���3�>=La�e �z���Y��H/�x��mq�@���OYY��7�AI�
Ͼd�I�'%�t��|�ܦ�x�8���u�iY�y��MM��٬��ǉ�z���x��c�7��
�������Y�Nejϙ��͡����';C~���?���vO] u+:��ڇ�}�6��2bN�{��n�o�׳���ﶗ-�
�)+;�x�H%g�y>����n�g��e�d��`���'�3�i4��:��T��Ăϒyn?2x��S~�̚zé$�<|Tx2.�3��|s�WI��`|ԇ�w��~AeH,�l��T�����B���oy���>a�5�v'�̘��"èz�8����T*�n9��0��w�|î�R���HO��wk�g���c���G����TP�7�k[H/<��O]�8�g�3�La�y�5�����I�=x�$I������!�4����ި�G��W;��t�履~ּ����?p�M$���!���a����6�\Jɾ}�f2T��f@Y�%CY�Co��Lx���&�m��'���f�6�̧��C�m �z�8��`	>����8�U_(5k�%�=}@��N���Ĭ���bAa�i18��~Oi����J����k5�{�63L�&��L��Ԝ�m
�d�ǯƳ ��!o�<�<s��ȳQ^Ua��W�b9Z3c�u��yo���z2��{2ub͖X\�#bǶm	��d���,�M.�i���Y[ҡ^ͫZsr.��A=�Shf�us%��zG,р*IB�1�aZ���]�,��yjl�E#W</��xW���'���1H,����~d�R�5���%zÉ����?�vr�f����i�gYP��8�
��6���5���T�4�<�i ��L���F2��j���73���~� � q�?=�a4��T>O;�s�z��WHzÎ~�*y��&��
��?$�񒢇S$���Y �����@Y�&0���4�Aea~�5TN�ן;|D�Ï� I�Ͻ��@�aY��a=vɦVk�<����OS����dĞ�_o!P���!��a�8�I�(c=d����`,�%MO(|��2|��ύ~��s�|�[9�wd��l8�IvвǬ�a���z:H,�'O�����E ���u�O��{�ì+�V�>��m��P8�������
,�,4�gS�I����Axņ�.�z°8�>����^��]���k�3�0gY*��Y�Ne���bM�S���s6�Xx£���8� ��}��6��r��}�M3�J�S�������0�>g�5��V՟�YP/O�����<;�?�����g�tR<b�z>C�5>��6�g�1'��<t�S�<������w�8��N!P��	������oY=C:`o�o[g+1�M�u��J�<���]]R��7p�=��R�'uf�m���k,���:�E ���,�m�����I�b���O�L�2��r�RmE'Ǽ��9�ɉ8���6�d? 	(}��c�Sr[����er����(t=�L���l��*�Y�&����Y8��mi����w���2s,�5��M��Ĝ�g���>�*����L��*�O�{��!�����?F�(�H��(
/O��<M��������6�^�K~��aX��z�Fq��$���N�e"�hT��'��0+��{�:��뤂���1�����Vg�?}�g�}�:|0���R������T���k>d�Y��'<�"�Y���a��B���bx�0�4�jAO3�4��ès*��dĞ�S/�y��z��_��������V�WN���֌΄��a� p�P�S;�E۬��7�`����Z̤tm�猍w�v�v�4��'6:�=w�*��M�G*�ӕ�>��r���;������9�Z{&���ބ�_Z�~�� ^�r��������?�����������3�J�T�wZ ��J����~VT��?w!�����Af�q3Y���"�Y}�4���1 �I�b
�'�{,y�j7z��C�|>�A�}�ɤ:Zq
�ydĞ�*N!^�2|釬+����Z�����ɤU���7?}�O~f�@�y�Y�a��<7�<O4��;�ܾT�韐�A��D}�=�� �:j�ʓ�q:�?��Y�S��m�����LgS�@_e������
�^�S�kD�0��\î3�J3�<�f�YY>�u�f�����{��q����27�!Xi<ݚO�9��C�޵<d����*Ag����k8�H.2k�5�'Y������+6[��.��� ��vK�G{jk뭌����bi�0Ƿ0��S�Ϳa4��§���&$�σwHz½}`bi�a�zÎ~������l=��;i���QC�ʐ\O?Y4È��ϫ:��{*���M�_z>�(�gw9�a�*)�>���z�&����y���&3^�ЬZ��{��3>�b�o(~CL�LC��?!��B�}a�~��+�q��b���F�5J<��5�}�������A%���~��O��;�i�Xc����N������jɦ������<I�!�m/i����U�!��C�Ɍ�~a�7�b(J�#��K����K�� A�{���L<aP��SL�%��H
,�&�wz�2T�!S�}��N?�0+N���~I����
ϙ+���]���?2W��s'��R�w^M;���J�?�����1�$q���4����RW���H,����Hm'�T��O���?!�۶�H)�׌�@Qa�滨m�zɉ=~�Cԗ�;���T1��{gqΞ�]zyu�G��������|�Y���ɤ�z�ɭ`���Z�]{`c�Z����Ag���p6ì��7��i�|�,|I�b9����Y6s|����& /����~�cs!�[73�nE�
��3]���D��mg�׷'��&�=yV�Al��[�܍�z��3�9�GQyEHz�E�|o�Y�uX��2n��6�R��g.U��'�;ن���۹�m�V;k��S!�,��]�'9��<�M�R�l���u��鮬����hC��w�Fv��Xc��=�x��c�B'Gk����I?!Y欘�������_�Y���m�V"�8�����k QV���I��B�C̳�^0+f�)�Y:�t�_�l�Փ�E�rɌ��$y�[�u��u�^�b��'/���P��;�I�m��&!̡��T��8�߲m'��\}b����M�Y?:gXTY����@Qg�6�՜d�6��>q�����~~�h񶳧�y�>G{z(�}���q��d�>�R=d�����*m���;�&���i�I��y��Ć[4�<9t���S9}b��q
��Rc����8���6��T�}��{�+f>Ί��h�O���@�G���>�1����P�%{�&�M���C�s�y�gY+7�~�*}i�3��06��P9�c�a������8�Z��~eE%���}���~��
�zkg{�v>��Y|,���H>Y8�M�����V5����:Ɍ���)=B��Y<�)=B�����m��+{ߴ�%@��Ǻ�@QV���&�i
�<׷�{�����-���Q����O�	q�i�f錬��'�E����O�!����A$�����7:��O�1<�Rb(J�&��wp�N�A����d�|6u�'k*���8��������]v�f�TY��5%@Qg-�����&��i?2~q������'yt�=�c+%}a����T���7n=a��R���u�@G��#¢=�k�9u�of����/�>�.�=@Q`w��6�
��T��>&�1=c�2`m���̊z��ِ�+��&$�uǨ}=��
¡��:�HVi������ x���f!nVW
U�U��{�ᷲz�1jN��5�Xx����[@�T����8���QC�icz��fd�Av���Az z��������ݘ�O�Vs��m'�*N����9�uo����]^i�Xi�g�Sh|�*f���@QVLi���'P��sA�n��xs���d�m�Nv�3�Me��fb�Y���N��$(cS�͐$�ѕ��M��,�Um��r�訫� �6ݡ��\�!HK���#7��y���䉇n�D��-W:� �����]ƒ����i��ξrhJ��h�J}�U���x �g��{�?/��"����(�i*f��I���+�@�1�&08�u��\�2Tk��Rw�6�Rw�04��i����wG�=aSL����lg̕�������}�Y�߽�Z^�*Ag��i��S`l����É�4��d���:���� (�k���1B���H/�>C߾槬<`~k�l18��$�L�|��$Q���(��1�7T�?zt�	�CL8���6Ì*'�̞;������T�6§�H.�O̚E1jZE���>}\`z��\g�8�Ì����f�y�a���nj�����]����w�M+�1[��ڨ�M
r�tJN0������x�2Sr��k�t�������>�[HÁ�\hmT��Ӫ&�Ɍoe~��L�e�C����w�?e�ab�\;�-��u���,��g�bf���D{�`�V3R��K�
�7�E�7C:�*��X�qƆ4kO8f�B�e�5o�kIo���CH�zX�{ب��ȭj�t����U({,���B�j�9
T<p?^������a�eÙ�u9�iD���Ve'��c���ߴ[�Z�l�L�'�Š�uĂ�s�2�24��f��{6]	j���~���Ҽ����i�=i�9��>�H�X�{������?5�t�=3��m����ÅY��b��*dR��%�Zޙs8�o�#x�s����N�nC}R��D��uu��}��B2ك�N�T7�lG�����p+;w���-���Z��4��+��y\����>y��J����3��.�x�@���x��.�|�����:�Xq�s�ru�r��C����|4�#�(k�+�}�i����������V؇2��#;t�܀��^��'_�Sz��Ѯz����c�Nu-M� �(uE������^�`ϸB2�Г^JFD4b��7;Zc�ʵ=ke� ͚jP�j��[���U�zl�@������u�x��K��O��\`��"���P�Pð�ECp0�&4��9�x��Y�\쪎�u�[�-I�H��0g�ލ~=���`c��j�ԙ���2��F��z̦�� `�g�*(;$���?��h���R�H�|=�s�4Q\�p�q��R�����S#cV�"��Kz��I�y�!(�:l��"��8`���,�5AE��Փ�B+/Xۮ�6�j�L�.c��X�u�H���}��gV�Kt�:`b��v�}wl�R��tN����'��r�n���H�����cI�}�\�JlC˯�M��u��
C��}�*���"|�Z;�f�};�2ħƀ$7X�Y����Lz
̢�����x����I�w�;ZvR]���  �vw�EDB#���&X=]!��b��\���n+��އ^cTڄ��ۤ!�K�y	��T��z��f�PH���V.h�9���U�8N2�K�'�� �/���Ҕ�%Am{�鱑��B�r�"
+`��9�"O[�M<����&͍}~���� ��X��ݷ~Gy����yǐfԢU��,���|r"Eڶ{#tl�=����x劝,Д�q��<rAΊ���������!}8�v+��xq�&�Y�Wu�\n����F(�RP���_�����֕��5>���T�~�dP�.��A"-e
�/ )�i�-(�A:B4�n�F�ʔVtVo�|i_�r�[8�)Mm��,X�)Z%ה��&��� +�Kf�J�2���:?D��C8z�����	�^�{����4z�w#�pȎ��{S�C,��o�_x�?d�����ʋ�9^�H�^(���b�c���c� ���d�x���\"M�H<�Eǃ,�ZH~ےV��YT���&������#���j����@`r��ib��\�j�mݩ�������G�Vd�,E��Ϸ6*b�@�sz�2��^4��)�MQË�v6s����ﾪ�4�ܟ��q�垭U�x>N��S$c�	[(y�
~�I�9�O�<�㊤�%-zŞ���=cbp�D^{g�#�Y�m5h�WY1�i�Ĩ¯:�Ց&i5��z3���1^L�<��t���C#T.s�	*�=���qS�Uo-��K9�ta�DU8�#ng���j'(���`QnD�Y#�'�f-�ks����1�8vb�5tzܣ@`�W��`�����i�ע��2x�tf��X�^�
�t@�YJb���e�6��! '����ؽpܖ���x�j8�E�7x��#MN�����ͪ�P��`�0q�^2\I.�Mрz���-N��"Ě��d%�ҝN�<V�qdk�@�>NY`�L�W�#�	��)�m����D����DW��q�aW�F�]
{|m��/6~��y���9���2����z��&;���M�B��^�\�C�i�9�N��*v�OVE��ӓ,I�&tY�Ƨ��R0��ga�ٚc�T��t�	,��hmܵ%� ��n�b�/Zb�@��^;���;] m�/$�IY���L��j$Vk�*��E�4��̹6�o3�.�Au兒�q�:�����6��=�a9�U�����҈*v��J���[m�Ϋڈ�烕gXYs�}�d��x̼P� ���E*�9JJ��jhP�"��Kq=IªY��0i�.d�c�l�0�W�	ӗ
�,�"l���yt\�P��"�K����$�	+�+95�X������$<��S�GUlN�l�U���u�z[�z2A�V��R����Rt{��]�㣑�I�ilΥ�ų%�yы���SՍ���X<���m�������ݸ������oGi�d�v�S]oF����dv5���[�lR�V�fD'Z�`P��V�[kF�e;���{څ���O|(���6�YV�7�9�c'G��W�Gn�9Iz�鷂NҼF��Vo�#��e7�t;M#Y]!<a��a��Ѳ���\������	L��E+�� U˲��۪��0jH�^Ԕ`��gCӈ�4,��=�]�-(�%v�cq���+�vԬii�q�s���Al:�oUoW���-�<&�oU�R6,]ro�ڧ��W��=�;�04�D�c����G[�m�'�`�I���[�����N�woB�Fu\v3�h�h)���t>���T�(Œ�c1�G~HTW�2�_�f)Om���s¶%�q[S3�
��j�������jꖊn���wo�(�����۸ӧt�@��g%�oI�8��z� M`�y��KZ�PtԴ夨���\����:��-�,k�+���[�t��Rܚ��˘���L�T��(��WZ堺���,�]����	�p'>�v����7���(�lY��f��]�d���P�)c6ށK%"k%��h���j�֚ے󅍊n#��,A�F����w��2�c��9g���YkvO*Ղm��P�[x�P�����v�}����f��8���k���V�X�;0`���e�2�A.�����XTZ��K%�*�ٜr6�)/D��Ցv�4�YR����=�����V&ܬ�P�)���Y@쪸������1޾�˓^�pC{j���t�ε��|ɤ��b�b�[ �jZ���o��jmpRb���������ڑV3��4�٫�YC�Ui���G�m�F�Qѐ�늠��Pu�]o�W���t�l�#�q�@3�Twufj�so�Yͧ��{�3�퐴�N}-W(t�.f�d�[�m�:uUnm3��I;V�@�e��R��AgF(O̯�qR
F�Kil�\a
�$��B�J��
��b"��YIQIK�C�f ��
�+4��咤-�:�%I�-�*
AI��LH)�����3��ӌ*�%@X)$����b)����,.U�J�d+	YYd��q��I�qRB�&["�
ɉ���j�3"�IRV
��ċR#��Xɤ�1�֢�(@��J�d
�)�I
¥@"˔4���) ��#ީ��?[ߤB�3urQ�9BK����X�
���	]R5���ca7A�<3J\Vfَ�g]Z��,3�1������˝���l'Ԅ�Zt#����t��
5vtO�i���S����j[Q��:�Ѵ�|Á@��1�Z�5@�F�h�����2p��c6p�ލ���������׻�ԑ���JFEu8�ϰ����X��F�-&��+R�����5�r����Y}щ�tx���������:�,�Z��ҋ�\\/��g���� ��ڄ��U�V�>Y{щ]��7�����2�r��ȬL'$Du�b��p*c58���}>�����ܶŀ�;=C� ����9`��OգLL.S&P����X6%��5j���ll$T��tW�蜋(˞�}w��P�^&������i��V�Tn�<��Y����,󆣎�gL��1�!ڹ]u�p��QN+�}U�HÁ��������]�K_f�߱�tfK\;9lf������.�������F��V��ꀢ8ŦhI�F����!̜]��7%��򡸞{�xꥀj�ؓ��,VS�ug\a1�޵�~8���_���n�g2����U�s#��p{C^���9uv«-���
@v	5����������30Z�K)4$�̃�Q����������qͧ<3t�R.��C#J4::�ʸ�V"q��V��,邏�{!+�Tj�3R���	��P'b��B�c���)��W�1^[\h�s&����ӭ͖[�!@��y�V������Lg�D�?%W��2��
�2�~� ���ݬz=��q��}0��@2��2'�eB4(F�+ٲ�nxƖG:��R��Vj��Iwr��P����{6��Do
�΁b`_@�ܢq+m�
y����ɮ}��۔d��E�0�4:4�BT�EE	�r�\��,�����;/�O�8��yq�r0/r��Ŕ�g�It��o@�~��y0��}�E
P�f���/:�Ng(��`�yz!N�:�!偔8�Y�=��A��h��:A�]ʬ�t��S)��+Ou"������H�.�Ɯ6j�iؠd�D��3��7�̩}y7�F>�5|	~�@.��c�t�F�8'%�F���(���U�E��v��:z7V�s)�G&�.u{�A[��M��n�:T�h����C����&*��B���d͜�on&q��B�{LM����+:�̒q;�v���S�,����u3����f����Q��}_UUW�^D��w���W�}��k<e�A�<�:ǟ��Q���덩ڲ�4��K`��؅B$g!��W������Y~��Xn���3�EqJ�.r}�&]ǧ(|{������#p�P�v�q���6��T�\6P2�*�A��#�KIS�s��g#r��	��f����Oh+r�R�j��8�G�g���`�c�I{6m���)L�նb�(l�o�y!8����_�-�E+��u�{h>=�vS9���!�s�$��tkS�l_��AU�(�e�J�V:B���2�8�j!�ûI^��:��1q�j�L9s�Q��0�o�BƜ\-���Q<��lu�o�b�_F/�[����"Ō�w �q�$8�B�rs��G��Q4`K1K-&�S.�F�8����,Д�q���!߱�B��Nv�VοLk���hq�;�CD[M�OӔ0�9���W`e厮6`��B�:��Vg��g)Z*Y9�.�f��j�2��1b�]�Y=��a�;l?������o��2Gm�Q�N�H��2�����D�g&`5's����X	�{����4��Rs��Z%��9D���3V�2WwuVUp�7y�Y�Y�+,ez��,��+�ddsxrV�ɯ�uk[ۄ�����!_���z7�����Hk�#�Da�d
2s�W��j
C�wAc�ˇ]X9��\[7� �*���k�n���5�Z,X�d*�_��r0l��3a:ZU�Q�����7�9�nL�x>�^��uE���/��l�̋/}�ȍ Fm A5�GT����f��{OP�V�
�ʭ*"�P̑QqF��Ű�<$�Q�����_����a�q���|���:��B��BV��i��8��vm��L>m�=�=�u�����}����vr�6m��r��cp�؊7&{Dc�Z�a�+�d4�i�,uP���V,gͯ:�U�R���n�i�uNȕ'k5�ǯ�6nX�h��񁧨�l@�E���"��;B4�0�����r����j!�j �p��BUGo�#`�Q3e`B(��q�ث��
��+��+�*5��]���y��Jb����	>�T��s�Wۼtt����ԫ=����S��w�zu�g�����Bk!V<�Z[W�J���{�w���ez�y�Ѱ��n�#Q���j�ҔŪ�])����xӶ;5��UŚ�Z� < ��Ȫ�͑�h���8�ܽ�<x�da�f}���ʘ%��
#�0.-���E�9
]�(z+2-;�Yޏ_��#`:S�u�M{�R=���#AN`�w�*$�¬�Q�b-p�h�IA2�ȡ1*�t-Eza;��_���#K.�=�7��l1t��t+�<��e
�/ѡ��?>�����^��m�\V�/"�7�R��S:�F�Tq~sՀ�)dA)Ϻ�2�͊���t!�VA97,��n=�S϶õ��w?Δd�Mz��@��1�R�2k8�>%5{V𰗔���Gy�)�����{��O�ė{�^�喇�	;�N��}�^�X�+Y�*�� '.�Z�k�4�0��l��4:�	��(�4F�Y��u�#>�(��O�O�g�p�t	��߷� <���U��xt��Į��.��b�
����ތN�x���s�.*��>���hʆ#��b:`��|j���#��v�uj��޷@�t\U�����W$���\'H�6z=wVOi3��ӿ[�5��Kw�\����pqu���?E��{�A<r\�N��s��v�\��2Z}���xu5�i������Gk��mhٚ�H�r��ZnN�)��������4nX���`�eK8)�G�S���P�|&���u�65ą!�t}��}�s����d(kU�Jƛ����	��s���L:.�
��T~F��TlH�>�v�����kՖl�'W�R����x{�e�IZL��P���+�����[*&��b���7" Q|�]q��=г������"��p�,���Ŏ,Q�ɑ�N�No�����c<�(�T\�n(��ΫUǊ��cU�������1��ݜhY(��F� �q�j�[R*܄W�0�~J��)mq���wl��bu�?F�lS�X`�I��\9�����������^�u��C����݂U��v��i�9��sڌ�C��w�Z��̐ȣ��;��(���<*ˋ�q���[�"�QD?k��$闣m=ٰ|�pt2#����\���>G��Zw!i�id�n��g���.N�J�)Ӯ�d���DgM�+�=n���+*ܷ���������k��Ԍ��<�j������`�ݦ��]R�����Wx)�Q)F�S�p�ByV��R�1�+�	��|@9X�$u��[`{�u���n*���C�V��6�D����������$[ �4��U Y��8��I���mv]��g�qZ9��P����S�wֻx�.�>�/?�X��WK�^�8��.�sA��ks� M�b1r�q�-ӌmz�dE�fTt����3�zfh��);d�D����s�:��؈�f�5�(�v�&׹��pfx��%%�Jׇ��b��Usf�H��%z�z���^5Ξ�x=4�O"53����Q��+]f|�A�9|g?)d����NA�!�b�;uɎ���N����/j0��E�J�5�Y^��,ؐn$b}��
zd��y:D��k`s��9��*F̓���)æ��1�N���kȹyY��:u[�H$q��V/�3`И�>���5 o%^g�:G����=�VvU^�S����0�u�s<E�#�Ё��������E�g���|;�� cc���h<�Խ7�sO/�(��%W�%
 ��]��{ZfK��>���s9�vͬU
Fh�������蝿wJ�=�W.YL��}�]�%�V�h��VBƇ�ŏ���+��bY]�Du.��5�p����R�d!��*&ގ�qd��c�	�w/b���i��Bz9bjo� �.���R����zDw���-:��[WJb�:�ŁQ��HF�d�p��G�ي(]o�U�U-m��(݀���f�0�a;�5�zr�⺀kÚ�NYdR�ڽ�;ut��)i�b}6�ל�z4ף]3c�x݊���8u��C��tTt��b�����oge��;~/�M�I.��S�aҮ2�2���ق�9�RR��&ᡛ�7�Y��j��8Êf�Tp�D�8�DYC+���)�%���ocs5��m�Q�W�p/^3zM���+�j�az���b��ێq��K�U���6�����U�H \���*0>�Q����%��W��.;�s?S�7���4E����t�qB>������kБV�Q��������ҡ�D����o�X{�i�<p׶ 9]�U��س�s$W���O_���BC xul�L��|��]��Lv],4]dN���#+g�>�Vl�i�G<�V�*��5�1�:��e�%U@W�1���S���&Lk����ʣ��C��w��нɪϏ��+E)V���0[����[a�RCĮط���{v%mr�d� ���J���8v�N��+Sy8�0K�K	v��ɓ��t���UU�7�oq*a(���!��]{o�%dɒ��\{��p��{΀���8����k/�[w������'ʸ��>�`�`i�Q<Fؙ�����B�9DO�'��:Q7�\�ܚqq�ʹ߮�,�J���b3}��'σ�G/�������"�]l�'�囹�q5�V��7��ʅ���,r-��*���H':ˤl��2T�[�����Ɣ�r�/��,�:13^��up���(Pe�n"�v��O=Υ���e�Q����yE�:S�ӧyu#}�ΐ�dh1�R��d��s��S#���G�"�'#�z�[�(�ݔ��@Ҳ�_
{|zu>HV��/�Wm�\��y�@T�Jgen:&OFB���C,�i�_x����rao�;�*7LB��Nr��K"�S�t�3�9���A���#�K�r���Iȹ�}1��W�=��Wˍ]�J,C�}�Mg�(��)�z�� �������˩�����:�U|�,���k2���J�t�o&��h��SX�m�� l#���P��ٮr��6�
�ϱ�NZ�.��ᎆ��eM��j�`�Vp��)��Hiy/1��֭`T��+��&..pFRvz���_{� H�W�tL_l�l�6�` x��zk�;�\�~<f#��u�t���Q\��O� ��~�m_�����'����F�����FY����sO��;��}\�D�	�ƈ>Ɇ���26�!�uQ�§=����k��c�U������R����wA6���aitn�D����J�����!��hK5�Mn��q���z]�ZdrA��ؿ)�F�v,g��F��X4�Uҵ]A�c_đf��zh��{���9C�5"�ß�`�{��#>�b�"g���M��] f��)����{�ʎ�nB,-�������	��+���)��e�m�����	��H��'<s�s�?:����h?��F��u@�3�1+�}A��frp��&���B|Joj�P��i�S�O�M���:��Pͫ]�=�ȅfp�k~(�&�tO��f{U<�:�ꡱޜ���_QCybg�x䄼�c��+f�A�Z��V�	K������[s	u��V�ȓ}�h:�0={&kE���5y&u�la*#z�|�U};8��͐�I�����VP�N�wm��.�y%���,��9���CWV�3�E�U�|�_`�̠F���� u�犮#)V�43PTcX�/�w]6��F�XW��*N�Tr�IL,���w"���R�W����+�ʤ���0�.Em�+�H�=�9�|���uyNQ��]\�엢)�vB�Ы�f�Bm�Ztm�WV]�ϕ����Dv�-��ˑ�����ȥ]������0,o�� �������mT�}�3]A:��]*�%l˽����qЧZ����v7	!��\y�&!�.����ײ�O9�ӯ{�L䖍�o�F��B�.�:������օüZ��,G3Ov���$����5>�[S�9S�C��@�47{)�H�ҜN���^h0�s&K.�!۽��|-���N򻪎�76��� �-��$c��M�+��oA���s
����s�]^Y�R��0�oVjZ�9\�n�k�k+O|��^J��(��誝��EO�a��<ʵ0�f�]̭T.mj(M�5��饪�Ts��X�RdblYA�]��c c��.�٭�ב�WGt�sk<qds�"zQ9A&%[{���6��j����<y�MJ�sVhv9&^f�o��EJ�u��o|�E�ؤ�Ǩ]����W�7��V _��Jy�r������5׹����4.�[�Kp���fv�G1u@r�QCi�,��e�4�jM�+�i&h���NƇ%s1+�ԁ�u�U;�]��Ռ1�9��YW����w;��u�4\�����Q��ogoU��=�˂���6^u22�6w(^GZ�=c=���M'�0�5�N�"]�&4d���B�bu�(6.c�/��ի�5�&�k\�H�N�j�;�ǝ>���DM��p�$�'\ 'J["��Mۆ��I�v�:=�q|��ge���A hꮹ���ķ�]1Ԩ]��jl�[q�iփ���Sz�um�k��j�2/h�|�V[��#֞�J�^I�<�j�x3;(��j@m���!�<��]p��Q�ـ�ݞ��N]��Ψ�Q�om�*j:�lvW���) ��*�[GӷH^4�7ev�l��*3ػ:�``.�ڝI�˼`�%�V%��.���rڬ�+�+H�8��2�?�����5�h�Zu Y)���Qt֨.t�CT�����K����jڜ�.SI������)iYt�m[��i%�y��w�����ςQ��%C�`�z�LAb��\�YaU(b,1���]01T��V
�L� �	�c�`,4�cIF
J�c )
+����m��Z 1� Y�,b�L���D��+%t� 听RVTA`(J0\��dS�,+a�HJ���i�(,4��`9LCR-�
"�,P���QB�F1 ��0@Ri��ɫADb��5	'ď~}�OO�U��v��f�"\rFp�U��lӛ{�d�4r�EZ�>g+�Y���/�#�,��!�rw^b������wA�{yح�����̅x�"n@��@�Bʚ:��+���׮ܧp���q����B"z�4������d:�+T0p�z�r�f��l,{x�k��\�ǩ�9�p���n��4���O�^��l
�x��u�BU��A��J²9�*���Jc'�8��
,��!Е4�6(P�VN�+��5��D�~��� Ɨ�P� �O}>��T��/c��JI�{zGʪJ�#�f�E�=⅚�1O���|��_��YA��xWC�G�]�6��eŬ�%���Y��]�.�I|�dG�m"��㮲RX,����I΄�%/����Wt�Gj���~A����G��	��*�*���x�6M�vrYf�F��t^=�<�m	y�x���D����:�F��T���$п"��[�F�	J�Y����/-6D�Ϭ�o\�U�����ϰ}���@��=��# }*Ұ����8������Y��a_�ٵ��qŝ���#�:��O3.�N�ިxj�F��c�����'4X��4�+�V�0��w���Ε)��-����u��yec�7����u�����'7� ��G(�,&�4I�5n*�bQ\�*��<w5���&��}0�(WM���H�#�lQ��ʠ�#f��j����N��tQ�W��{��%a�lF�W�_X���`���Y#h'MB>��W��Ҵ\38�VY<I�;.�v�lw�	�E1>N��F�9�(�#��5�������}�#[��j�����Ob����u�|�l-O-��4UtJ(��Yj�V:�;�L��A������Cج��j�!Zu���R�r��x�P��<r���J���)S��"	6�͚��}{:Q�Q��	ߑצ�h�th=�?�x�WC�N9p*r�U�y��LIx��~��>s\i�)�tq����jtf��tA��YE�R_P�-xQ Ȋ��x�ɾ��,���q�*c�^t�a�o� �u���Ԑ&�s���V_63�躵$G�@�S������(��ձ>v�߻�z����9�6vb�w���
h����kl��� �UNG.��zqj�{��@+|j�(v��Qz�-ꖢ�C�s�3k����,�Э�J�[Vզ�v%Jjj�g�-2��̧�a�<�2�a2e[׫�ū�7k�u�!��P�ci���i�՜'՘�)ϳ���%���7�o#4�nT�׍Po	´�|iZI_&L�os�NwsS���_ʯ��v��wj���? �X4@q�5&��/J�@V�W���_�^FG�����<�=�S[F�)'5nS�B�ˌ":C�`��qB>��e�E��d@v`d����G�oT�#�Si���u��6t�d�a������g;{{δc�
u�Q���fp8�V�ܫ�z�) ��PxЇ��iS�X�e`uXxU������͛5h�Q��n�ۮA<��]�0�>x3��/5�a��2�P��`�ug8t�Uky{a_K����=`h'�xI���>�ݍNTG=�0i�O#F��<��B��+�`U�WX����F�p��=\�)�91Ϧn5	t���V�<�e0Ud�T�-蔌e>�~�&�w W�*�8ʅ�a����;�.�5��>|Pѯx�����=YKrc��s��	���^�7`@}�ܽ�x��#Mbf��unf©%�S)��7R��&���S
�������)�Zt׹u#{#�'E��S�V(�b��+V�G��~Vڱ�<;��7V�]7[Jo�V��P��i嚠�wn���e�k�M��&dr��ƻpZL�'r$������W66w����M�G�'��tx鑌Z��6{r:�.��J�xϴ���/�MGb���]��E�,&�J͑�	�C��>�Z#M�0�=�W��C��u�nj)tck���Ot7��Nq�`��t �ۖ}1�ưT�G�h�'v䱺T�8���L�ث���lB�;^L��a�����'Ȍ�L���)W� j�SmC�yOr�-�)��Q.Eea�Mϴ���J����Yr}�"9v����XsmVM�Վ�PB!��$Y��v5�.҆�றU`Cy}���5llr�:��l��9J�m��ߪ��߼�:�IWB�ã���;"�	ꮼ�o��f��)�Gck���6��帋�(���h��#E[�lq�,/y|*�3����2Y�+��(�7V����OC�(P�!�[���*,��zˮ=c�`��%��5j��7<7x�K�n�]���Qlm�!�Q��]�v4�s��{ c����F�����W�����M�c'�zK'#�S���w=��Q��]���^{hmv���u����3ۯ��G�n4h��KX�H۴-]���;�|�C�Vz�t�`�k���n��SV�f��]е���YZ:� �<-�X"�4r��d�/�{���bө�:l���O8F̞q�TwG��Y�s���]�n�_Ǿ�y@�\4�q�T/����A���B?zjlT�W!|��w�WB�"��7�x��ӄe�g��oVF�[鑖��I7�6�P��D�G�8���h�#�q�o���W��YƼ(wM��@�Q�n����@��GA�8ب�B�P��#B�
dz��d%E�`o�7��_��S.�v$xm��T��z��즘���c��P�~�*L���'v�DvE��Z}^���a�.���PL�di�n�Q��o�d*.b1e�# �\�O�%8�4�;������^���z~K4�!</�z�ט5B�g���	ˎq�����2̎�!��mu��5��10f�!�})wa���C�^4��ykՔ�'V�Z�3<�g,<��Z�m�� ܓ�˦��6ѕ��x��L�ھn�?Y��]w�̕��R�U�l�@�\�������C���}�&�Pmjd���Z����y���G:��8�k8E�t���]v1��޼�8��Q�r�)��2�L�t$�	1����7o���z󂝚㘝v�J͕��"�wg,�f�ϋ�R�K�����@d�l���O�ف��ȃ9�XO����E1��]dK���R��}�t휇���>ݝԂ�YZk(j5�xr;�b��ʅ�DV���9>8,�C,��H��k$U��U�y�h�y.��@���a�1�P�n �iu��;3�P9z"��Ow�%�{{/��4���Y��tc�(�#��G����@g�����if�KW�s�-jH2$���}) �faci�X)T�Za��,vw>@�ʯ}ԍ�,�?���_���	~�G6#���6p7��ܵ��^U�`���`��閲�]k\ՊնX�T�;}v#�q����㠎����]�i�=^�V,�� �a{3�s��@��ឯl:��-��님�erH��ÅV�c�{bc|V�d�\&����1�Sq`������K֝Fǯ�])�t��QGHE��6����&0�*+�b@�Y8Y�Tam7����kF�o��[���S׌\Ֆ'�7\5�&L
�뫔�&����v,���!�Ee���40M��`�!���In�j��޸"�p����@@'�˓������[I�/ Uq�\$���Q��Ɗ{�|�|9i8��[���%�~���Ӎo�~�P�_)�Q�u��"��^����t�ɍ,�S��4q!ᷳ��#;�r�"�/��F�Fώ�n,TW�FN}�:T9C��5�Ι{�ѡEε�xJ,hp����;#���ExN
�(*��$Z����;Z(����I���lE^ni�BՑ�UY��F�3u=�Bb�ld�Hc<��T��m��ȼ"�Y!�p:@q�5'�D��`�Q#�j�1x5[���	�c�{�\{�z���,��"/�!"}���b1B>��.j,�"`�E�����%ΠY��U��ˬx#��cP����.����*ּˡ[��gAK7���q':c) �D�P�6�QNr���`XxV�����Sf�	�������F|,`#C;��_f^�:�v\N#T.뎞����m�o�{@�S�W[��s�+�9`�����&E�$��h��V6%^g�Y��=�vR�얩�9����o^���b�O�т��H]�U�R9����S[�+�:*����t���.��<V�<�������D�����wpK�t������v�qC�]�6V����c�_��FhQ]{ݳ�wLR����ɰ�BI�7VG�c!(���P�dJ���g����9����\zIUۆ��.3p[)�j��~64Qo�<z�T�/Ǧ:��u�5=�!Fi�/g�τ���� �d�gw��x�&,��9�H�����f�0xV������y�%�mřlF�J�iZ�$�� �Ō��	d���{�:t�S�N�r�Dd=��Ui�}[}�-s�i�*�A{�H�rh�����E8���7e��4��:��L*x�ft�^q�^�g��U�ǖ�>��_|��^8��t��b������z+N��Y�H���gr,8QN�9X
��APϺ���7��A{�etγ���6"p��Ԩi6�N�]�a���E������L���)o�>(E=O^6�t������u��
fa�jUT�`���X��� r���n��*|4"w�9w��_�.����)������Ex�*�]at7i5�k�:�Tp��/���^�ţj��'�GL4`H漻��Z�ɯUKu��J:��e�ӡn�ebѱ�$x���יS�2�<�k���T�Yë��X�w^st�)w�u�y�FsB]�tUwU�7�2;������\����qp�A�;@��}Ӂ��m��gtK77��UW�����s��;�%��>�7���?fq�Ueרȴ���k�#�F�ΉMV�0�v����{#�Z/|�X{��e4U���:F�>�;*U�y�%��f�k�h4���yB�rŽ��&([�sǙ�=�:p���n7�2���z�z�6'��GNq�\�}"��cKqg&5�b=��������f��S�l�*@ˌ/Ds�h�N4�F��P�G��t6"�ܓ�]�2"��f�7_(�I�ާ�4���nvB�}�:G�BC������?}s��c�B�V���J�ˋֹl!�T�f3�(�D�X�@���%���+�;|{e�����HT|=��gJS�dFD��}Z{����@׺e��H��8Ш�mH�r�j�ռ�k�)|�:o[�3����u9���fΔ܁������\Ǐ�tv�U~J��x��\���oit^F��,
�]'���FC8��eZ���$2(�������M�.�p�7a�C��c~vU�f�����Y�Ք���v�^��b�ӡ�{$邴�z#��#=Tt��Բ�P�y��!B(��:�������8�j��{)=؟	�|h��Ԋ1��}8#�)E;��}TW�Ol���#��~�.g�`8��7%�Q���O��^�D�j ��������qt�y�ŒNfJq��t��f��<C���� ��u�v$FM�G73\� ō�
'6#��PN�	��צ0�sG�VE��p2^�'����ٚ+�UcU<4�[W0É1��
�A������`�Ҫ�x*����;2E׋vvσO]kĽXt��jĔE\-ҠXz�Ll��Y�`�=Ʈ͇ؑJi��� �M]�v�t�Hq��h21��U����|	^�@_�83=��rCp���9q	���|����ʫ���� �q:���6�@�n0�PZEA^Mv׋g}L�oq`qf-^�)�eU�������r�����������D���8B6C��O���'�S�6���}l�,mC��yV���;a͕IR6g�Ƶ�]U-�u���׍܄ƪ��q�6g|��ň��hL{��Y#[t�>ި�\�0�EQ�-ԍ�������\#���t�2�j�Ƴv��)��� �u���=R�CO��{S/EtlgD�kݻO��Z*���ڻzN�w|c�B���6Qw,vy��t:/� �U:ջ�q2q��a��`:��Sɗe�(�h: �������1r=���Q]�mv��[��F���y&j=e�g#wVi��=���Hu��S�/{"nF��k�X�Z���v(�$��Nޖ_U�b��w�[�s�{��!њ2���͚a�	���͝7�e
"�@U���-��nAc�X�O���ɤ�q�7uhD��V�}��WKYLTB�� [�B��ׅ;zU^�,��qע��C���iK�ٛK@3���53��_HZ�Μ�����1��=t���yG��{v��l����d���Nw����q�Y�C��h�����I]pҐ�I�*;{�`��+��^K����(��w��*��e�|��`v(w���f�-���V���mS���b�V�ihX�����b�׳��Ί�c�M��p��Ыy�%ת�Į0X�%�K��qFH�:�6��]RƘfP��1�Q۾����Y�9]ȣ�Й��������}˦���p�B��n���3�Cde�^�(l���a,�����O�����v�
�U6;��\K1m=�5��u�<V �>�M� �˪귽�4W8�P�k�JA��9^�8�`B�"ial��W�-`RT-Gb"�ހRz�-g(>{{���b��ڼ)��ћ딮n�5�s �ձ����勭�I0��N�=?u֛{׮r�)W9�}IUb�k^�8��B��V�rUy���ׂ��m=��x�[J���5�u�۰��m�"��lm�i/�gN9�U��`K]A&�RA�z1�Mkz3R�R��h��fۥdoj=��
��o ��E-�,� 8�k̗l1��k�-Y�M�9�I�Ғ����t�
�oo3N���-R��3{S\�<�Cq��n�o|CJ�lB�쵝0��sYW�Ժ6p�tq.��Z��\r�����{�1H�6�L� 1>'�m���C�z��i����*ݱhZ��i���,�7�}�}v+��S��&���Ot�WE`�bsN	;9٥�����u�ǒ�۫��xt��7�a7h&5޲���9�W�M�ޖ+;�䖢ʅ�-�l�+��9�k@�Z]��[���W�o���K�w��-�V���=��t�䧀4�ik�`��ƣն�jo_&�`c��Qa�r߮�(ԷH�]J�}tV�k0�G�PJ�[������WE�/�10ൟ!%�5uջ�+�]ޤy˫s��3�g&������\�.O�G�Mzy��]�q�sK��]`Z&��_ w3*��L����=�矏ڲ�ڬ�11���Zŋ ��iV��\LC.�9j�1��R�)DX�%W*(`��E)q
�ˑ�bLh��1��6ʆ2�ˉD@c&j�.�4�AUkm�4T+UW��b1a��b*�\�Q����R�jز.Z��X)mFMZ��
e�(1*��Q�b�
iV��1e�m
��b��ŋ�����B�E��&3IQb�((�m`�X��MfCC̫dZȴDƣYR*�EJ�l�*
Q�	$�TQ�$��O��S�����i�����f�Wf֒{u��f�\r��O��X	��7��n�O��u�tJ�JÇeX�����������pFW`z�[=|���܊�.��N�-��q�E^������9�Q�%�n;b���ʸ�F�9�(�#�	���!8�~*�"��9�x։�����U����lA�l:-B�=5�e�N�T,����r�K�ȳ*�Q�*�=c]ǚ����.��IF V�l�Q����.Χ�$ib`[���U��6_@�Y8Y�Q��N���7CF+�����Β���wS�b��b-C>�s�q�5)�tq�:Y�N���m���Q� �f���q��G?t�2�Уg�<ro�Ip�2�@i��wawѪ7e-���I�i��1�	p]V�����F�:�LT)=�uB�E�*r�X�S�N��k7y�36"N8z���O���s�ο�.��)�|k,����ݬ��|��@���
s��L	��+�O<�V5�>��)�]�q$]>���$&�.c�4�oP�-G
�̋S�X�E���@�b1B>��e�E����#����9S�[�bM��ʚ.��J��H9�+�|�	�y�GZ��g/��Y��Rf�Y#��!� )�Wv�/T�\��� �Cc{o�`}��Ye@���T�k���x� (~�˃�!h:���복�� �OCq^�-9z毫=��}�s�nL��Ss��4��$Eʲ�!��x �¬eP�Q}��TE��d��.�J8{W�90�0x�)­ě���Y���g�>���К=52�oy��c3d��,�]��0� �ь��z�O��㧁�푏WP��i/p�;���\%ӎ
���1g&9�C.��?��[:��LVU�!�o��<�W(�ܧg��ފp��C���*W�����Y���lH�y��B	�8� x�D,
}�-�7~��������#Mbuw6&���κL�9ٷM�O^L�RJ��'�	�P�z��'Tz}�y@ӥ5u�Os͇��ҵW�I]���#�c�A�&����q$A���E8ba#vS�{r09�{/%_A\����8�9��Z<�p���,;叁���#M��q�į6ǃN��{�"����|���z&�;3���(
$��߂"���7m�2j�Ю��Ab�^���Us��4ϖ�:~�:�Q��gsW��rul���`@��y>����e)�ȸ���KI�[��LF��'C������o.������2�8�(��s`��:"�>sV�Х���Q!�Vyv����~pK��#(��a9ފ.�$�uتP�	�����O�D��{��w�q�$%��o"�W8S΢z}����Y@�A*F�רw,�#�B�[z��W��Fi0'[�}��� �*�]+�[�=y�<�]�q��	�ޖ����jћ�"�Q�����%]�+�A�i�nP20��X�q~�&�)�I�'�:(�q�6�l�_:´��a#E[���Vy`C�^�`{u7�K2�W��5�rEs��t��
.{j��/�`��-ۮ9�&�fQA<Ӽ��,3�E���f:;��a:i���	�
t�d����ӎ�k�v`�jå��WEc��e�����S:�>�S��,(
@m��x�wT ��?����>L�����q��>t����_�Q�>t8��������<��%��ͬ�`�O�֙@Д'٭,ٳ�^��3-�d��ž
���G;�kbVEɔC�		���OX���7�lY��Hl��t��);���;fm�ɶV>��u-i�=0�A�"���^�3gfcj>��g�چsc�6x��p)��LВpG�@�l�y-@܎(׺:�'v��+G�]𙴓�A���8�S���0Z�� ht�4��i6�΢�C	�����{3͎���68��;���R;<Bw2ug+��r�Uˎ��:���rvS�d��SH��k�L\17>�]\����,��e�}~of.�]��HZHd.1�Y��l9�����ز��`V�]#d�Ȭ�n�i�b��A���ܐm���c���
L""X��^��@��*D�9g�蓜a�hwO��F�r����-�ysl��C�^����W�Z���HG&0� a�WRt;�x-��T��*��/Y>����a��1��)E��
�l;��F�$3�d u�7�R�z���̊أ��CڬIDU�ѥ@�����㮲%�äX������n��'6��%Qǝ�(�`��@`�T���T���j6Ј�;a��F�6텪&ǞK�Y�o)��/hefXVp��󻸽�f�nJmN9}`ܻ�I���GV��9H<ݰ�n����M�"�@���=S ����9���ޝ��^Fy'��;#,�m��r�N�5<;� �RyE�܍*D�+R�����.�+[fi<~�U��dH��WS�������)aB���
�^.�y۝o�߰��s'��QӢR��2�(:�N�"��d�]�J,�\�������3���n�/q)V�1��".�s�����fSX�ڳ��ϕh�Y�49��v�=�gO<es4DfH��lE?��t3ƴ7�l�R�#��N�c�:j+cn袸ΏRH�/_�_W�[�)�lk�<bG*�
Þ"��GH�@�	��v�rOy�*�I�2�X9�@8��F�Caש5Kak���,�D]�AU��h��ˌП�t��b��D�׳hU[�"��(N3�8�^B����:��`:u��Q,h�gz-&7S�G�8V Q靤n�_@��,��ݧ~F��E��@�3�e$�=�#&|��8�!i�8���)^r b�4.񕺴\��x<���hc�zWZO�N'ΤEXG�X#_k��]��kƼro�Ip���E�^�t����L��W��8�-����Ψ�V�U��:�Sv�.�|�v<i���F���\xgc��t�h��ŕ2�|�$ӳ�^����הMu�Z�ܙ7�����v9@�wgp���-`�1�+[��r����{�]��t�z�����t������U[��[�_63���[����Uj��Wɝ�L5��4S�\����r��{����+����|��1��/�=����=V�^*��gMIL[�FD�#b<�)�`Ͻ�+fQȀ�/��Z���nl�� �9�k�t�q`�J��Qb��EZ�j7Ǉ���qh%50̉m����F��O�t���t�p�x#��xXxj���h�Y��Z���1�ը����a�%�U�u�'+MX� V3��j��V�rӱ(h�}~)��^�B&1�w�_o�� ���E����p�ơNa�׶ s�2P2*=�`�雔�̮�a��Y�z����!t�z^����S��<r�=\V�ȕJ�[HK���F7k��	6�Ov��=	F(��*z���j��+}���y�C�9Φ��Z]�hkDτ���ܧ�����~=>��[+���k�.E���㾄K��s�e��􋻴�$����N,�@e��'�{{�޻��7@s���I+���HS�Z�-����%�g��w�E{�N�vnX����4TȺu���c5n3"[3��و�O��(�+���o9Mr�i�9�t�_WĒw���(��LW�Zj�cA���=�-�7b�F�ܽ�#���pu����5��G}Oܪ�ʘ%`�8&1�U>�.�Tz�J4)�w�/nʙx�{ �z�3{�`b�A��tȍ�*EY�]}OH��j��jce�����;z�{.F�]W>�q�Pw�=�Z<q�0�@�b�1�{݌�5�M�8�S����{\j�q��C�+G:=��ϭ���:"�>sFބڅj��K�9'r���2Ta�{d�.Q@�q�bS�]r��-�`�b"�7/��T&�0��Z�K�0>$+�тx�qX�^�5Uۢ�xVO������3~72՘ŵ�^|�%�ҕ�[�L�1	X��]aEQ�/`�.�M����'iȜ��sõlJ��}�'��F%W�#/��'�>ZUyud�3ʻ�I����o����9*�w�Ʋ��j��A��h:뷈��v�|�B˥���n{���⭇��6E�%1z.�5l��ˡOD6����c�B83���_ulVf���Lˏ�!M�έ_-��ܱ^�Y?b�nZh�k�.�K)숦$=�]�f�� "'4C�30ѩ�+���؅p�D�2�ܢ��^��K��.'���$aόy^H��yB�r��bb�L��n��s�hœ�Ĭ�gg���+˕eP�T"��q�z+��v[���;�ods�\�JA�f<-��S���{�N:.�VԵU*�`�G�<8Dy�Q���_@�E��w-���<^�V}Y�ܡ����N#�ٺ
�*�h�Α��+�g�M����ܧ�<A�ŕ]���m��(�ʴ�-F�<��bf���=�!�6G:M@���6f�D��t�������H��q�F5Zy���!]2��D���l#c37��e���Hw>��z�v{J��k���FGb�0t',���.����qu��7|}t�H}�/X�o���VpWC=���ʎ�pq ʵAs�b�W�57��,z��%@U_�C�w[PUt�K"��-���4�;���}q3���N�5dB ��#]d�t[�>F��r}��q�6tY�=�ժ�ov�Y`[Z�\�vX2�������Ea�~��S��ޫ��.`�a���i�35XT�-<�� ��~o-|�/�ޮ|���D8������w,Kn
�z�`�mܲ�r,�{*cN���V6��Y��Fp���f��H���%6$���2$��*q����'lذHݫ�s�Z�W?�i��"����U��E	��GZ���:�L�rcv��\�J���Gz�QcE��$������W��y4{��.����U<��WB�3��Br�]}N�$�^G��[a͞���BMJ�� d��L�xM�k1ڿg�����z9��+ꌧFȜ6�0�P��Q��2}�#�l��(-�LjA8ɍ:j\�r�^ӻ8���}I`��o��ꅊ�������5G�����������~��w�&���Zwy�[��;<Pz�
ʇ���r�Ɏt|)U��WT�5�3ߍ	p}��s��E�s���ϡK�c�ѵ��V����ؖ�������7쳯:��~+�����C�yh8e#Z���e'AИ�"�F�v%]�7�-U��oT�9���P�<ӟ2���-d��D�1<��n�㠎�@�L��f��@Ų�s��v��"����#`(ҫ������w]͘肸�4�Lېi��g;�V\��O����z6 �I�M�r*4�1X6We3
�;v�I�́�[W��S�\8wUT
0DoV����nl�:mĘQJ.CGN���̱d��z�
���t*�x���	�(����;��c�[/����"��֨�0��(?D3��3S�+(���7������anӿ#n�hS�]ب�$����]HI8qU0�9���C"�mT�y�Q��c�{���� �n�QWe�֬�OK�m��C�����jiyc�1ji@x�CPeN�������Փ7C;1=~'�s0������ˀ�U���l�!�j�t��*`�Nl�uR���^�w*��;$HJ{ X"Kq��Y�i0h�C�}������F��	[ʹ^�l��"��R��ʧ�����b=C��x�Zy�T�ͧG�P�mh�=�V},8��f4��
�ә^��ߠ��%#`t�1B>�*�M5i��oٹ��i�� *{���??��[���x�K>s`'��{�}E@��}+R#�,+�ʔ3e�*qvVχ�`����Bf|�1ޕo0����;w7,&��w��F��q�%��Z �p:�w{��:P�@�eW��p�5}B�#LGXh�{՝�{�uˬ�N�5�R���k�)'̝�\�����ѵ��Z�4uFA��'��b;�8�:d�Yu�#�=�f��.�!�܊�pgE=��u;��B��Fȷ]oѐ�L��$@�ʭ+�N�]3�׊UX�=b��m���)(;i�}�i������fގ���C�+)k�ӐB'z�R��]&#������>��s�Uv�b��Ivލ!u�nb�r#�K[&�C2[Z�9�;�gh���r�Y��&7.8m�)[{�l�D
-^�ڳ|��O�pb%�H��e������y*=3���#h0�)�W��Y�-��~��̩JZt�TK�+[�\��v�����V�o�p��m­� �U����6�҄�[�\"��s��Bip�J�����r{S]u.�um�A�9X��"�vZƫ��S5''P��j�!ϫ���	|����g�RR
�AU�,f�s������^�%��v�k�nS��m�K�	^�6�mӡ;�;�`W��ĥm(�j�]7{��x�pG`���Cd�c�v�W]�P��r��i�Y�#牌�p�nV��+���ڙ݅;vuN	]�<��0�zY�5{�9g+7Fi��ڤ���1*�(M�`4ھ}��5r��:(���]�5:��u֧s4���;I�i�8�9F�L$�It��ͻ���u�:�r�*ys!�nG���m(m]gd�"�mM�"q���Ν�$,���z��H^F��n�\�Vň��]+v]&�vrΝޮtoj�,�C��)�
�*�G4DU��3��oj�|�ێ�^T�*�,"�[w7W3[��F���â"43*>ө����e�f��ᮂ��tW�;�����7�WwN�s�d3Y9,[�i1V�6B�W�recW݋��2u(��/&v@E�Y�2�����;��>
�cC�0\V�偗 V���l�}��Ek��۳k&WI�Ȭ3�����3��AW��>���W%�W�������YH���x�D�N믹S��.�6�/�ba��Q�w`}�Op�Ng=VEɏo7O4p��SmS��@���(��(�[Xh29�w�&��t0%j�id�R��O�Be�<
�j�Q���=���^V�jH��u�c ��^���b�*�vZb�)�R��K��P��[[l�z�)�C,��E�VC�����Ž��V��S֢�$X)[����(4�f������DjQPL�UE��b��eE�1F&!X�R�[EQkX墾�DF"�(�T��FEY+UU[b�*��,`�V1U`���E�Qa�4�)1�YJ���Z�X6�4�X��EbŌE�(����E5J+Qb�֊*E+
����J�Q�*0��X*+"[� ,���1Qƪ1QY2ш�T��1b��FF(�SNJEm�(�(������Z��Q@��J�ږ��h2ƥj"[ahR*�EAADAu�.��}��tz����.s(py��'�������腹r��%B�`��SY��ЏW8�`q�X[�Zo��;��0�{�o�|�����)����p鎁B�S�?�U%C֨����ۜW�|�f����N�p�.��IW�K����U�M�}h��4�1�e�/U	�7٦ah��֯�?8����L�1��#N8�)��N��N�T��w.7cC���(�bH��TG�x��.ԣr�
]\Gp�l:`'C����wpcu.Oe7<�u ��Q4�\h<fa��{�y�v��aϴ���rL|� ��PE��Ъ�&�"�{+�a:�saL��{�@���7*��w:��r������ә���y9��\Yk��g�R)�(�#��l� �CU"�8���hoN��[Z��u���Di�~���T���o�K���*���F8�dg<���3�ˬ�o\�
��t1;�4*3a�q}��Bp�yX
MQ��}�˝�Zo��3��-p]Mm�"F�g$\�2����';�.��k�
VӲҭ�N�b%cj�Ps=�|B�Ѱ�0�������u��Eh����Ú�@��%K�����h^��d�u��(y���})ؚ���ޞ�:N�������@#Զ�R�v̗k*u̻Q���+��Ļ�Vev��������S�zF	�)�c�z��6�~^�����[7�\�1���fm�ʓ���J��J��
�>������\�<;=P�ǲG^=�^_g/h�A:g��]	�tx����~D���&���5��
��P�lq=P��]so�ץ�T�3NG[f�C*���.o���-(��eL�Rt�ҳPǒS�)yYŒȓ�q>���@�5e
�rŽ��hz�[^Z7�w�nD�E�����w �'��IZ�����H�P�>�Zw�Ej�x8�qgv<:C�s#�Vs��C���|7�xtoԚ��Z��3���l�N(tR��}J��!�Y��t\�%N�̬Z	8w`&:�lE7$�_��W��;4'�xT�>�Ӥz�t �HYqk�r1UD���6�q��դij6 p
8�,qb��>�D w`sܦ�h�R�PprHB�������0�`5h�7�klv7Z`ҁ� z!��"b1����Ba%Mت�l�����vEu�gt]w>f�cpF:������z]J��=��nK��#�W��1��8
��/�Ȯ�z�:���^�Z��]siQ]�oD�PȸnJ��{wp�5f�Lfkuj�'Sq���>���S���(n�d	���5q�;
��R��6S���SqS�@�t"���Ŷu�9�'}�<s���|],_7U~}�,ல�-k��Ȼ�B��p��m'���P@��de�5B7!�Qw=BxF�F�7EF�WI�Øe8��Uj��/Fn�� ��#��d�t_D��mVQ9 d�lG]�v�m){|�ْ�syz��k��	���J��,��_"3�&��H��JUVӭ���B,����N�@&R���2�K4߁c�� >�5�U�u�L�qt�ϼ��],��3�t�2�;MK�zxm1�7�˚�.b��m����vR�o4t�s|&�pOx��.�Z�r"��sl�da���b���2&l"�;�g�"Z�N8^�(��$ir���{�P����G�Ъ9h,�#U���k��lM����e�%�g����؇QL.!g�2��3�~΂�[��yG����/U���K��/�4�hF���g\����O���]�PQ����]���ї���P[�NcX��0^^'3^Ī.��q�q�YWPop�˶<��ͮ5���ȴc8���ʛ8�j��<z��DB���3�����y3��j*��my;Q�1�E?�r��K�z�Ǵ̾���?v�ٽ����[I58���Y�^o��}T�n/+B�{Qs�q�T���6�}���NSI_�[�ו��W���=�o��!�93ѵ�������֩�{@&��u�)Ob���E}j��`��hr2Kj�tNk���M;��Ui�m�����k�r�)؆�����d�����9�=�M�;���OU��6�e�Ư�P�O�9^�DO$�P9j7�#V�M3��O���Zk�ywG.bS�����\C�9��!⡙�4�Zv��}4��Dds9��t;�ϹU�;Dug�����r�jX���wK����ȗ�zor�Vф�D�p����0>��TG�-��Z����*]�mw�hȍ��:w�Gj�hi��&ۛIu�gM�[���p�y�O*����{o,T �K�<f9.���/��n��3n�}ٸ�*޳Gs���oe;���c���j��:r�����W�Ư�r�rIAG�� OxҨ(�[��y՟J�\ѵ8�WG=ݕ�Ðь���h��k�6k{�����:��S|OM{p��WFk�}�3��#^�k����߉��23+��vK��s��;uCx8W3\#4�'tPk�x>�ȫu����ppZ�t��6�.:�g
��P`;c5?V�v,p�ܮ�����9���Nǋ[N���f��|��X~y�-��$����� ֞����޽V�8�b�Sa�s1��;��t&��y�T�"�]��F=aNr��`�.5؜jB��V�Ux!��йH�p6yCT�ݿ1�Ǌ�Ӛm$����=ؔR�9֢Q�T��mU�]t���Fh�퍁��L�~<��}��b^t�@C=�݃�1�b�/U=���P=�Lu+�6F��T�����-��7r6�%`��H�Ywu�h��e�u���EB�3��r�unW3Ȗ�O�epJ���w7�����n0�l4E�G<ˤ����v���e��ޫ����4��ܕ�?�Q��7Gc��7��f~Rs��彣���DO�lq�6+�эfj�%#E�7Q�e���m�b�Z�z^�x7���E+U�����Q�-'�S���w�D���{�Uַu�J�7E�~	�X�VT�Y�͕]z9��F��دNZ�D�����u�����)���M��*��u�#{�B�Qq�㋢�]W��P���Fݚ�����;s*b0	Q�9�7�u��{�����'�ƺ�(MZ��V5��D�LŤ�tWt;��ּn�(��SIVEu����`�WU�����J��
w�q�mmv���}���Ҧ�s�Y��t8=�Fà�$�Qk�:��&g�Q)�z�����m��X�6֚�(fד�2?v�TRf��W�=Y~[���u����9�檔��J�8��~�]V�{{q���P����.�l�����fwZ|��e؋�~g��\}y�w�@Vv{1�O���57���f�c��ۦ^��'��b�a� ��ۼ0X=ī�WuѮ��^�o�jR>��v.~��C���9׉���F���C�:�E_E1��ݥ_$�R3��d��<��c*�ڮ�ް"lI�Tq���ٹdeu<�4�p�^���%^��7��K�4�co� ���9�ی̩����t�l����ۛA�ԒP���[�ێS�

|�cEùiJxg9s�e)�w;�o����U(ޯbg;���FVe�Wݔ�6;����'h�'2�F��X��{�%��y=�|�sMo]X�t{��(+��ⱇ/m�MM[�ʵ1�ul�=��-3kC�g���{��^�&�{cm�B�
��H���캳;��;����K�)=��u_|�u�uu�c�<5��_��5}�up/;���[|���F�5���s�
7��*��5qZ�sŬ��7$�߳[r�E��w��G��ùꕬ#�<���t2��w`~���l�3��@����v;M:��PJ�����p�~�oV1�Ŝ.�L�
�j�@v�O�Μo����O[�g���K]��m;C�y<���5�ܵW�	_ky�ǎT,�D ֭�g7�����D�~��̛T�*L#�W�>�q7I���ԥ7
�*%#=��U�re�W���'��ezk�Kr�{>y�3�Է!}Ó��1�Jٺ6����q�.�8=�S���Zj!�N���ٻ�jn�VS��oq�|kwO�o*�[�*�RyAq�����gn'}4B>��(��k��|��R3��٥5�ګ��(�� �R��X�`N�u�f�1��5J}ܪ��r3���]�n��4ml�"��l����ɵ\�PT�It6�\��������$�s��n������k���K�M-Xk����Q�M�\�Ea����%�{)��gU�N��\vpg�9fA�u�p>�='|�S`�ӷ�#�-�S<��������Vg4]_\���̃O��K�8��8������l劮q���<�5��y���ڥy��uV�y�l앩���i�瘤�QG���r�q��VU��;%6�Y=�n��w|� �L��.O�:�W��TD�i
�v�=��n+����tt�]�(��jմ��n��x�
�Hy'�W`�����m�n�/kC��ֆeH�ýێ���*�[�uМu��̦��Zn�ᖄ=PJE�/�2*�P	�є�h�<�W�T*�ۙ�}���j��9-���4TSZ,;���l���0
/ ��Oqat��Q��].�=��^К˫�6�O���^*����w�?sV�k��"k��5���-]Lg�%�|���H���w�dnq~�շv{[���&��D�=�pnA�Qr�>���R^x�3n�r�?W{m�-U����]o�!��bfsf�ȀN����;�O�bg���e�|��P��
_n��8<��J&�봂��7.��<8�Yy�wf
Ŷ��:Sl�4�GJI $�ߋ���2�6<8������7F?f���Om^�*wD�X2ىL�<�ú�ƫ;p$+k
�0Df��vr�[۸At!����>�UU�UiM��˜g��Ͻ@��sk��<ժk��.k-[<*��K�{��uTe��`�H�3S�-#>�N�v����h8x��/(&���2���ՄԷڵŕ��Nu�UG}�Ґ��ڪ��jt��B퇥W,ASA�*qs�H:{AHBv;�q���q]/�'Y�;�*��df����1[ؙ��Ȑ�b���n�ntl�i�x���
{�vѭ�����o����Kޠ���~�J�i�W[�^Z�UY��قWUȀ�U���u��wu�oK�
f��$y�E����s��qǨLgE	�p���w��C�d�t,u�\>:�~�4���W�\�a��a=^���F=m=����5wm�^�1���Uʭ_�I�b"y�{�5k,f0?����xT�|&�ɧRj���ش�"���*d+�[�)6��"���S� k�#*���	�V�t���ɫ����Z2.oLۏ�Iל���p��567��4�G�j���/�\*��S)1g|��ټ@�~1�H��In����S����ڽB�r���T�ZOg:���%k�{����v7̝ r���v��t��>�,<�-ޝ��L:�Nz�g�P��iI��N�j���{0b�ڽK��+8
�@����������4��fs�L����I+�-v�tޖ-L����GʻV�5�wi��m�b�V�9C��?�2��^,:##���r�C��:
�f��ЎL@k�SyO�jG� 3�S�^��[R���G;[�2�9oV��,�/`��-�`	��H����:)��d�y�J,���q����I��(��{P���C1�nNvwz���k�~�3��&o6�s���1-��<�L�����C1>����wg+���7"w� e9X�cn�R�#�&�ovvV0Vo/�e9���=cYt�,{u�	���F�Fp�tr��sX�������ëO%�F��F�آ=X��[�ߥ2"V.96�l�]��̼�3BۣuK:�ȣ���1���ָS|�Q����kxF�M�Q�t���S��Le��;/$�Ѹi�Un�6�h�ke(��hض/sëqb�uw��{�:r-��b[t/^P�o��|�N��j«�h�۝�Յ⧓K��7�֭���_2g4Y���e�Wf��T^�:��ݰy%� I2�:.����jIG��CVi����ֳD��)j-�V��1ۃ1�{i��B�oS�Q{�*ӵ�@�Wƒ�)�Z��9�+�$d�[1��غ]�f�%�*.%��z�A�Ŭq$F�Gp��1g9k��k]@�Px�,tn�8�Լ�us��^�"7H��5���5=n�<ơ�����U��][�y
̭S�i�A��Wo!A�N��d��
�֥�yZ4�a(��V��-�6M����N(�g)-+[#{����	˶w`��+)��&�\��>OM�3q�Au��h
y�WZIz�����X�RQ��卐v�]*U���kIW����S�h�SM&7.'����E���nC]����ִ��+%<[�+mwa�v���S�V6Ѓp��&搥����K[���A��V��8�,F��Vp�c2򷜝���WFK,pS����������[�wjl��1�[d�jJ��<������z��ޮF��R�[����9Aj�RV����h�}�I)��h��[�{��50R/{��@ܩ�M�گS�L�YF�I���Zs�g��t�YS���$�Yڹl�c��;��|vڷ�r�xp������ݩ�B�_Kl�
�uUdm��Ct*�[b����K��Q��QE���E�j�(���jł�2�X��fZ0Ab�VX��Z"E�(#2Ջb�������F(Ԣ1U�b,QQf5X���b1���UJ�Q�-*�1TDb��-`���(�dF�QU�*��(�`�EDF,u�0D`���(��1�+W)T����R��������#iH�
-eX��cbS-QAH���PH�ib*(�X��UDb��`�5U�!Dĥ�2�EamQ���K�2j�DA��Zʨ��J��VV(PjB��j�UQDU���f4EATOG���_s��EV�C*#�\w�+9˭r��w6���9��so����+HM&�l/Tp�::?诫ꫯin�%Y�����@g>n�:�����Cg�?&�x1iv���²�d��/s_���M@�Gs���ȧ7����L���t�x龼�l ��硵���Z�QU�-����e#�E
@B�Է�>��u�x>��4/�Y՚�U�#���=C#�pe{Z���k,3=���N&7�;����LU����ОS��1wL���W3}������J縫6(62轪譄a��Iz�Z},�m{+�,�w}����5��5���Ϸ!�S�03�6!�	B����;+�T3.��7��p]ʹKV��mJ8�C�"�(��5B[����SD�]�0����Z}��(ެL�X�g)V)�k:o2�1Ij�i��R&vb��cN�U�6��U5ݎ�z�+�s�G5�X��ܘ܊�~��z�	�t�L#h����="�6�d�<�Q����]��߷��aG��~N=.�׼�:���;J`��:�}�g��7;P��	C�F��%�Uv���ÆS���i�oٳ�1����
l��Ď�ӝ�V�V�y�3@�R7�1��Z�m5����^ӛ��G��Ak~�N	�ꌾ0-��OSi�o��;{�y����g��{J$dm��5䧠ꌜ�Bq<Tk���8���4���dH]٢pQ�=G�³�y�q�:;'�+9Y쬾��Wj򔻩M����%5�!_EF�2Jq��R�F���vLf�M7��R�#a�/�U�5(����aö��7���~7��.-����Kx�UuZ�*��v"��5�H<�4єXy��vYN��j�u�D�蕿:���YwQخE.�3�ɞ�ό�t^ҙ��o�)q7���p�ܼ�����X�i��,^b�孷I%8��9f�y�;���l|4.ew��W0-��^�<k��g���5�;>��i!�ꘪ�l.q;���WX��	�.m���Cj��[5jD)t+�.�[t
�T�<�,y��e���n|������0�I�{Զ�^�4�-��u�͂QM���=q�;�#EX�߇&�ܹR��K������mWB��1z0�'��z�\5)��7]� �j��|���k�MjN��O
{z=���ZޑNy��s�o�B��Q3̠'����ܰ���
�j7N���y�e��1�n��r̊�Wc���z��7��y�t.���2����vt���Nǻs*�#�B��9}��r�dt��l�7g�� ��+��,��^?v�Мj�>ol>�?G���L��Lv<u��3�C8(�=���5C�oq���VzVϹޱ8�|w��N�.�m;���D�٨�������2�V���ys�,��iȵ�j��g��>�jQ'"�p�_�5Dh��Z,8�� e'���|3�yt�4��]��M=:!�Hz�0�}^7�=���G몝��n�:x�Z��x~�ne�&�ktcu�g:��C�^��Z��
�-g��̾ZK����<�[�Gj�V��9��Ga��Ǉ�[��3ZI���u�&ɮy8-l�_wb��##"V�av��7Sgv��fܐ�G,-��4|҇���h����8>U�5�\k'1�ۡ���5��4�:;:��fmm�v��5����t�U�S���'�Dv�ob�c کr��̗��U��:�E�.�=#�e�~��xo��+�]�u�4A(� ��%S�і�
#oKʙ�57�㙩v�����߹0�*�z�&Ȑ�}����7�&��]	�V�5j����A���2�.;q!�.qm尚���P;�
�N�;��i��W�0b�#�x��hw���{b)�ӧ:��P�ْҸ��FD��L����b��'�9�.���@���ʦ&ES(/{�sAe��zI�~������S�[��z�3���Лb����9B&�$���\���yx�s6�Iy�u=�Wµ���M�;�?"��ӗf=�z=F�� ��֌�;���ˬ�((�<�������a�K�Q��M�s��r	*l`<�h�,�%���K4�
��ʁ7h��ߛQ�6��6�	����M�(�c]�u�95�
ή.�un/��	�K��\����d��[�Ԃrc��d�6�J�C{GUP�Չo*�H���sn�7��~����S�P��1���H{ X���4��	ͤbMv
KNӷ'�9fh�O�ķ��⃣�t5��E�"s����[��.��(8��έY�<�DL���a��Dӿfv]�|��mq��g�����k�6��	���2o���Ȕ���x��|T/�:j����O����;��|��b��ӊ��z:U�i~ܭ��qlߡ��TW��\���[$^s�����[���^�ؖ9�-�q�Q�(Le!c:Dz�nXs�	�6QF��(��P����jGM<�ڙ���;��s*�53�ßPr���wL�ʊ�ثMN���dsY�����ثcu��¥*9Ұ4=C�W��2���F�,���S�ڜ������#K�#wN׷�����]� ��;���R�+*B|8\g�:�r����UU��.+I9�ת�Cٗ��j�ә���T���R���v��O�X�U�٠��e��ǋ��u�Y.��p�p��p����K��m�u֩r]oTV�٪uc��n>]7����������T��v)ৎ+$Nݪ����L��!{���Z�]OU�w*���jǏiO f����w�q&	5|����Uo�^'An�w����Ƶ�v�L�mu���

�N�+���=�f�w�o����:u�^T�����WB->h�^s�*җ륱e57徶�Oj���ۺgѮwF��'�N�&��H7�
�*��q����x[�"1T�����׼���K=��^�PQB@]ghb��E]s���l=a~���՞�w�gWz�C)q�jǲ;�&\�8�s.o�2t]�zfD�n�h_fڛ�ח��$�%���y���)9����#q)��!8�-m���'�s*�NC��*�h���m,�3*m9��8�d�=sI.ݨ��L�M�޶$<��j遷a�������V�9�	��ƙ��{�{`s ��Ayu����I#�ꎩ�_��o!	����E��L���䋏ta�'?B��ms�߼.-��({�,�U��)�2���U���~�b���篪�t<���󃛐U`�s�Y�R��!U_Pp*�䗫wqcr�9�Mm��6_lP\��o.%���x���㉢&�$�V�=�JRUJZ���7�n�}\T��ű�-]�yz��3�,��oj�m4�m�pu�ۃ@�LҢ��]�������J�S,W�9�o�ާ��K��ݸ�7s��R�7{�P�]��j�
x��B�-1�+��7��T�5�z�mL�Y�I���ڈbi��o�n��QNYb�9P�R&y����I9���ɭ���F$�_��$Ӿ��PFsHW�5^-F��o�� \����jA�U��]�u8�'��k�*=#�K\{.-�H���p�F�ޣ8%�����t�1��w���Gg&v2�ga������}�g�eeOxf�l^�}�e���W�2趺�tP
$D:��9/�z�����oFRALfr�1$;r���&���n���@Nu����QK�o;j;���}�g�x���Ԉ�!X�Vp�y��peve]�I�
�bar�k]� ]��m�)���������;Z�d��$�W�`(��:�2��潎=k#%�( .E�:�����K�/�Lg�q�������y�~c�}�𣀭ԇ��A�yȩ�ߍ�|�yґ�D��bhs��Nc��Q|B�p]-���%��9$#ڏ�2���I�B�H޳>S���&��GW�����`ݬ}@Ä)�}ƓȯM/E�$�ˆ���i���,�T��Tv�� ��A���S�3N'�]K����/_-%�7��0E��Nv�e�1��
ޥgb���WC}��j¦��kb�.ek֕O!5������w����L!��ZF~����գ`-u?U��J �>���z�y!����o��ںHV�<A�;����		5g�|R�	��=ٻ�K����ƃջ���<yI��n^�զ��R�%�Ps��s��o5���Y2gf�io%V�y=2�(OG,uf�P��\{��2�V�6Rm�x��ӧ�:;!���:���U{���L>ޡt��w�����T��%@�ގ��\�J��٢4;���)-�l��~�^��wR޴�wb�$&�����f���;j��	��$�`�:�Mߦ���7S��Y:�	{��w�8\�"랃����{'�����S�U����B9�=̴��Fm0z��	��P�T�t�W'F����߫�-���}�J-�v�����9G0�^�
�YЗo�F��6-P�N�gp���c��SKv���r�fX�zz�\.��Lvyƺ�yc���H|�ve�VU��oٳM�1�H�ዩ�ֻ��_Oh~?��)��zGr��"��@w�#�"����YƳ�U���vK)y��A�&R4��8�m^�N��3�Fݖ�5�*D�7ʎ�Ed#�,�rl����W�~6�ގ�=���8!@�ݱT��q�GwE�� ��ĵ��Ht�e��]�\�n����{.���+p��)�|���k9t�Y��!�і5��=�b�����"�B�5r�ޫ�O�kIv�K��}N3y;�����^AgR�╴gF����6r��"�-�G�f��T:y�w��4��+����Gx]V�`2KMyk�ތ����������N���Ԏߞ���0ՎЂ��*����nDU֝�\�r�~������w%�*K\|1Z/��/f36w��ݯ7�W�?,�鶯�oSԻ���-N�T�͞Xs���X�'���&�tf�m�]N����v��J{����8G ���9;�����&�t%@��I�t�N�n�UcȤu8�Vg��5짯�=6�9�iO�w�m)�s֍��z_�hJ�]���G��u0�y~��p�Я��8T&3� �ܯ.P�p�{[�[.�e�q����S��٩��a�*v�n=Z��M����9f�<��ä"���4Xi��d����9���B�����U5p�3Y����dt݆�,)�Y�Y�O�j�l�F���\�L��	,*�IE��,�s:�5؇'�ʶR@N�.�l9�;h�2��#�8�El�m�FJ�V�u�+���r�G���9]j�����]k��3,����Y;��T꿂b��S�S�vM�6i��Mrq�'/\Ǘ!hsή��U�� ��8�{�M<�S.U��0j�b_ƷbZ�P�e,뻶����&V�-�T��3�-7~PW���[��z�n���G��J�}�-2)��c5�3(���J��2�n6X���(���P�UmJ*L�	��HRn잘r�4�e�p-�^[hu�}�_
������|�.n�.�s41_D�yC5ʶB�y�W|9Ѻ�]5���5��!q�x��.�@R`�г�y�6kuj^�Q���8)S��E������D�+,+��̚��ǁ�8����+�UЩ��hׇO�+WC��L�#Tx����}z��uv�<w�v���_#�u�x%9�b���c���K�bZ�&�[����s�+��ڃ;mN�;��.��g���/a�k�o74\s�2�)}�}����zښvvuJt�-�d�����p�:�Yg�-ٝ�u�:�[Ogn�V�/m�>@C�&��Wz�;oJŧ2�;K��v�� !B��B���&�zgrd����It��{�!ÛV,���خۤ
���7&|�1]�mr���hJu����]`Ҷ�Y�LS�p���0e[��G@����#B尦�Y�����*jٟjj�,���H���˒��P1i
��M�\2��:��j�������-:����7�ظ�P�0�`�I4�=yѸ�#��7�
Ŝ9��
��b�vn�<w�RA���=�\5�hּ�P��V�X4�����+(�X�,P�h� K�q�-�`�yX�0���2a��c��t+6�\���d�Q(�����]c����<�msU��	�XY��w��G+�p��ط�WU�7�sd��P|HtɖBx�Z�{�U{�5Xi�ܦ��J|���m����^�#���,Tr�5̭:��G[¸Tٮ���8�����b�q,�z��snLS&�+��
S��CXPڄ��h������3��>�t��H�� �4c�ny����eh��]����Ց����7X�+d�L-f��ʀ�źِ�p䲵;ͷZ�o3��W��weg=:K�ӯ�I�i8�1eFdS[��hަ~@��V��߅���W���N:?�X�gԱE���{J#2؊�S-��+
�Kj�\�V��JţX�K"�Zʕ�X堂�eتZU�1�b(�ִ�(*(�$FJV���"�.XVDAq�>k,EA-
��
U�
��DEk]8��R���Ե��EUJZ ,�PZ1�Ds0�PYr�TU2�3,Z�@�sF�r�*��JQE��B�4j �UE�˖�L�d��QbȦ%���c[#ZJ���cR�V(�+	ib��j�dĮ5Ơ����`iֲ[b��Eb�Vk
�Ҷ�b�""
�(��Q�"�b
(�*�R(Ҭ��m�5���2�\B�X��J��fU(����e2�q���m�PYR�ڵ#l1��a*"�T)hY*J̶�LC�l����Щl�E�"$R�ڪ�2�G�j~��7�R��|�߶�k뷻 ��YV�{ǰt�C>k5��;�RYB�v.�iV貮�L�yX��ww2�"�Z�Ȁ(���AUty���zT�P��v�J3BuT�r�d':�M�mu{@�'Ͱ�����{;���4��%{��[��\3+�e���V���8���ڂ���VUJ����2�9����&�/O|Z��B눞�(є,����̩����!yX��ѵ�84k�e��x�k�ݥ:�9~��x�m�3�닠sZ[�� qǦ1޾�~��;T��2;���q:���A�͡׆K��V�#��؇I�p'ȩWm�I��kl7y�q�D�\+�
��v�W��S�Ol��5���ls��������f�7�sEd^iG�^d�i�̓�|�U�oi������J^y4��o��u�f�ʩ@[���4�:��R�d���眊sw�fh%��c-񂎾���{u0�偫�`�sz�"��^���X%��VՇ��9���Y׉�K,u�:����!U��Y�@�'T�X�}�����B,X�vK��9D�gQ�|�s�r<yu�^-;;�1�/@�<��z��<W�L�Q�qX�qƖ���s}��8�lm��v������˘i��Z�r�ХhY�h�漮-�Ql�TUwo23Sv@�Ʈ���|������ ᡔ�W�6s�W&����ʱ3oi�omn�;v���7���G���S��jzw:�ư�+�*�+�O*��-]{��5��7�4m��������2e��A�~��^����"�O���2�{���S���婪�M8�7���.7����:v�[Y���]䧲���J&ȂU������v���Or�Vxj��f����Y���o���Y�bw�tw��?,�*���[�s�Ol=}�lս��P�N{�6yz�����vj���o+���^zFl�m��m�QT����T�u�:�]+K#�Ǥ�(3���\ Jˍ�o��s\yg8�ls���;���[�,q�	ʯ��xJ������k;�3�����,bs+�E>9h�S��V$��ј����dQ��0,���C�]�J+�aK�D�;w ���9����{Lr�߇��{K��/.�މ���؜�G&ֵ�a\BW�q��f���2�Փ��*�y���\�c�r�ߜ�ᱜ�5�9C �{��9��Nn*���R���f�s�k�R�s���ދn�ԏ-����ZG2��ѝ#�y�c�'ϻ��S��5�|5�Jo]��M�9��
���C��Y�~#%���e���)����;籹�s\��7e� ���R�k�sZ0R�������:��[�:q���<�_s��7�/����c�\
6Mӡ3��Ϣ�V�ي�V�R��m[��
��M�j�w/F^�{�G0�J5��UҟB{@�*}��g�Ҩ������Ց�c�W'��Po�g/�	f���x�Wrڧ��/g2�l�)�bj��x��'�8=�FeL�������N�"��Q=�fDg#�T��H�*#׌��H=Y7v�w�)���q��9��ͬl0��	� ��u&2�l�8����1�7�hjf��en
�y�Fj�t)�R�Q�Z5��׮�-���@� 6Cϻq�059ԏ$�U�����΁�{;>���6�n{\:o�>V���-qj�l�YB���u�~�1۫lB}�F��r�W��e_��:�ie�M漫L:ƊDN�I�g��e=የ:�wgv*{C�7�[n�]�%m������C-z������s S{��g�G�ʝ�Sx\	,W��렑]��=��m�7ѫ}�Y*n*m����`�3�3Y7��"'Uޏj�3~��J�n���qoQ
2�;Mt��|�O1m'�˷��T��l������ז��@r���Y���t"wSkә������C��=ś�a����ݻ.��PC8Z9���:�^M.�����C�}>��^m����M)��S��w}o���A4���6�T�'%M���^�zg�թذ{9d��x��		ܼupG�m΍���d�f��)U�o�:�A�H���(|��;4P@gq��:h9W{ܖ�<2���`�*w#��)9�7�Uru�rf�;%+(�L0�p�B�[�ʝ��-�x���VE��ѱ9�Z��j�5���kG�vd6�▝�����#g5�gd�0��l�p����nC[�ӏ�QM����7��t�FY��U�37��v��y~��P۬	y�@T�P�ίF_Di��b�n�4\z��a��tl�I��t%J��.��#�lB��J.^Sy������y���Y�k6����ls�G}��'�5����ez�h��o�z�j��x&�e�p-dO���HH��9�:�W:�k�p�vC��g:|J�^9n����Ե;׋���D�݁�غRGNb�x��5=o����.k9����R"�v=�J$h�;�y5�b�$F=��v�a������{o�"h<���Nn�+�XD�0r=m�Q��Skv��<�r�����룤6��9��3��s瘕��7�q�H��n^�:�b��sUՒ�ڡ��k���ɵ܀=ӆ#���9*v��aB��Z��U���)N^E�ou��e,s����5�@;w՗^IG�B�ivە!9��kw��^�J➙��]vL�a7�õ;LU�S��X�/.F�&��˶+d��R�L.|��&����Tlڱ�jQ�.o�Ӝ���&f��4kN�r�r���O�+�C顣��N��sKé��{��:��}�g'�L\.���Ձ��V�%��F4�;<-�QL*�h亍�|�5�7��r�tm�Q���+�HZ�g5��\j"3)��"-��v���cu��V�9z��i	��т��ҾUr����ⵉ��e9�k� �t;v�q����{���vyX��rR�[����l/����튷�TUm�M��U�WC��5�M�Pz�:��­�Q4'fb�$�Z��OAO��;Yj:��
�2��1�>�d���N��~.�J�b���:��4(��mԾn�Nۗ�]2%J�$�xuz囬%5đ�y��c�V`���G�(g+���uW]B��1�'��4E��f�(k��-�\�я�C"��#�X����q���kSs��+�<���?{�-dTT�Eu�]r���E)�ړ�p	)��ZLJ���9�$�nS�&��̿<�=6���������"�{����c+�����wg9'�l�d�:�����m�Ln;݊�n Fs����*s��CW��:��:�8S�}	�Y/�z���rA�aA�ê��m�i��R�v��{�gi�ާ�9[�����O!�+3��%�BW�q�3R�k��'����*��Ǽ������a==A�����+�������z#0�A��í's׶��j�Kw<��6+�)�}�QB=�����mj��b݋��҅����_jm���4N��Q�������T���[ZkU?>R*�P��a�bg9�q�B��{bjfcx��2�]�^%�֫�����8��_m7��Wo:wFu��R��/lt;njP���h�5 �m:f���:��6WJ�+�7���JWe���
��M�a�R�u�Z��Wz�<�9"�6��t�ڗ٩ٗ:�;��a���/z�_*��b�g�rצb��K�~@��;�������)[���L�WTΫ��n��Z�WP�D�"�����N�E�]z�?@T�S�F��;}�J|!=��1F�'c/�~���(M��{�`{
�(9ў����,[��GT�.�^�QT��ddk;2��>�*�PU��v�P��Q�rҁ��9%]���':��BO��N�ǭ��!�_��Gr�W��eX{(5I��8���aZ�[�N[�bG��Y�˨Sۏ�*�]
�ȏ��B��(�n��ʋ��wG��kQ���V���c6����޼k��K޼��՝�mlPc����7`d)hT�������:�7��+�A��\�N��@��q�Q�*r��^s�������V&-���r�2��,'�&�F�\�3��NZx�d���@N��W�����mwpZ��ܶ�ǐncWq�oϝaOR�ϩG���rű��+���M�F^�xv@N|cKA���]p�� ��ԩ���ͳ�4��x�w!���wNV�9�-m��7��5�?,!������_�?}�t(|�OsU��{vdl�{ΰ뫕������عg�9���^�6��JG1}�j��UԹ_��q����w%ꗱۻLbsb��^r����ē�i�3 ����5>��^OU��]��D��w%�t���^�+�R�9B�S��S����^&*a=��1<�/(P�)���*:lWBCig�uЉ;�
䬛!�L%պ�kw��u����O{[܇c*Ҡ�\VZ��;�l�МBj�� Ӌ�;ʆ�y;+F�tPT~������:��bLL���d�$j�Z��A\�eh�*��>]GK
�brks&8�i�<����]��n�̹��oO1����2Uc����Y�H�S��ՏI2n�k^4�+;=��	,8�"�uչ����W/��ea���<���Iy	�m�a�=�B���Jxs��F��n<;�aK�e��_^�Qu�����/v��Y�[V�zn�t���B��fc�-�KVC;�a�������(	ה�,�1���9M��*�/y��^R��GsL5tHǹ��Q��D���k2�'=Sq�l�y��l)�X���[Ch�N���4�K�X^���6�h�w�v=E�<��.�\�p���U�|��}y��^e8�軣�-�6�G{��h��.z��j-��r�9�ɭ��6l=�39]�H��l��m���gy
${��+���W��;�ht�.F�&���ӈ�s+���e�05��euW�WQ�8_�6C����S�hVc;Rݖ';�i��V�q���u�yq�e�P;�B�9��7�U5u"j�^*�s�|�Y��};ikQ��S�WBZ8�I
��N1�dU,|���gU�n�r���L޵J9�,P�R�?�`���Q���X;�3~xni�ko�Lk�8/�X;e���1�tŶB�``X�
y�b������Ͱ[;w�\��}�w�t�# w@�sQQe�r���JN�j�z��Ÿ�syW��P�Y$^��k/jt�9m��K��QUa��	��Qǡ:w�L�^�:^���J�k(�n���Gwn�I�t������YJ7٧;7)E���tԵ��O`�)<��J�sU�TP�� ����s�R�7̗M��o�,��zr��|�:�p� ;��2��xA���V�Wr�9u�@m�WZ��"��{�[V�Z�ܺz�GS{���T��aVGy�����j*�HIT\=j�N�zs-�����H�������Jf���Ӡ��VK[W�ISv%$T�|�X�XN굁JL;oGZ���)\(;��k�2�`7�`���U�v�η����F�^;�N�N�}�iFMc|L�RnDk�#䯸9��7��ɢ��.�a�f>��'C2=��Pˡ�Z�[�f��8�������U�rĘ�Jm��9��r�}�Z^��xwP	}��A��&m�}ց܏v��}(G$Nf+B�}YEpW��X�g��V	ʭ_"��Y�"��9�,��\�xE����,;m�R�p;�؝(�kӉ����`�tR�s�hRЎ��+qlkz�����/X��R�k�p�c-wM��dAt
�
T�d��y9��s�W�4Q&dyq�ȷ:ŗ���_���䔮A���Q�;�CM���eu�����Pw.	�����L��^��i���vE�m�f1�2Q9�����M

c4�ݺ'�;�).�]Ɔ�;u(�/P�_1q9|�]J[yV�3Z�p`Y2��]n���^����5���p�
Pʺ�N�����Z3�(�,	b�pې!�5��A���r����c1�l[��fm��j
R�K�^�*J�֍"���ܥ��]F�r��4��7�U�a�%�������&sVؘ�T��0ћaM�w�( ���#{KEf�X���)F�}g@f�C�h#�LP��˱Ve:Q�%�V�=D���B�$��Xcf�����îG�㹣�"Yomt��G��2"k`Km��r�є�9n_�KE׆�������{��������4���v�ٰ�:�#X9;<��u(���pٌht��wg[�lֱ*Fo�΢����o	�y���sp���wc�'Zt�x̵$r��S��Q�a���[MVU���mAdPm�"¥d���+Dm��3������#[aZ�+YQ�DR�b�,F���E"�T�)�YbV%eAaR�0�E�V 6��U��J5�ƣ���a�+
�T��clX6���-(TD��VfU�h·)X�VT��Jԋ1r����̢ਢ�*��1��EX���-��J�&10j�e�4P�#R��VT*J�V��EB�eB�hU��j�4Ԃ�Uf"�++
�Y[m�m�Q��)R6�Eib��iZ\�d��l��WC�H�m��-jV�Ɩ(�V[eX�֠�-�m�%ml��Aj-k
�6�ŭQKj�VX�ʊ���KAb�*Fб
6�2��
�E�3 mm�[b��(c0`9eq
�@�1��jc"��%d��*	�QLq����IYQk*���e��:u���2�Qb`��*TH�����<���(K��gy�������غn�:�|�����fY��ղ�>�:�� nۍ"�v���h�J3�q{���IKT���;U�x�M�dVg;�n��*���dPi�KȩK�i�����K�^�s���]�q��K��v%,ʊF:����jȏ0)��tg9nŢs%=���7Z;h���C`�U=Oy\ˡ�����Bvg�u�{�-^7Y�-��u�(O_-U�W/v����[�*z66�*�:�gnbo��9�T�٭o�V����Ү�>�'��>�2hq���:��*��]��^���>��]B�wf�ϋ~�������˰��F��� 9�;q��\�q� w9O�Y��מ���ɫ��̼�ݚo_nXC�=/йW��
���� WiRN��W����#&-^��]�qC}����^��Y�Zb!e'��j)�|�!G�M۬s����L�t�*�y��v���]ڬGy�h@S�D;��dҮqf)5�%fن�V	�%��Wj��YN_w1��
"ӈK"۝�͗�9}؄�.��v�4/o�)������Ls#Y���y�0�2E�R{���P{���J+��Õ�M5�z��stb�7����T�q������E�h�nY��^\�$U�M]]H�q����cs���������5ͼ�}
�F��wU�d�m2�>�4�?7�[War�y�nꭇ�����q8���Rx���*��K�0�����}���v�v�?N��xַ9�9(�j���Z�'T������:�&Y���je�T�u���jT�.��Ò�n���bV����*P��5�f����#[��Iי�� �z���<��m���St^XVQ4�W�3����H{n�U.U�D��E��N�\�R���Ǭ�(]Q�ޜ1�^��T]�g�k���:6EU��A�8+ޙ��Y�<���윽���Գ��R_�0�B���<�2�]�Ђ��A��eY����՝ �Z�����lX,[��x�p7�P��:SY�s�3������k�@W^P��Uj��h	L���yي�Qth��=�h�b�J�A f-�8̷��IR�������:Ӷf�n��Yk[<N�jW,au�iHȓ��%r�LQa�"7�&��c���w<1u
{q�'CJ�Qo��	��<��.&;��qT5]뺑V�ؔ2uuQ��c�gG	OL�j^I�����5v�����%�w���7'=�N�D)Ꮵ�of�h�7�rRkq����=4!�ӌӎ���b�����(�\�P&߲��S�9�P�7y	昺�[��H����\�3pvQ�������)�8D�H�ҝ{�O���t�{�J��ü���|UǾ2X/�,�.���*y��V�����ɵ�@[�b�mb�j�u�ȥ/�,�_�L�0���:j.[/W.�r2��]y1v�&��d�}�~O�#�M:���a�vSX�������^�@NhN��W/m��SS�]�w�Ym��	P;j�u���F����f�����㳉�� �_W1���~�o5QU�n%`kH.��wKy�Y#V�1"�3u�ܾ�2����P&�]p��1��;�M*f��R�^��b�(su��u7����7!=�oN;�>V���)uI�v�w{WKx��;�1�1��n'���	��N�Lɇ�!�LGM���X`��B���n�i�x�e�vӅ *���֑BLu��gcw��m�*�E�z1;v�$cy�e�R�(�쑰�U9kju V�;�tf�����ǔ&��=���)9���'�;Y�%E;����g�d������OZ.��"Z��Ⳳ]7))\�k9"+�؆�F-��]pk������f��8ZB;62g�}�ת��y[Y9�s�ņ�����4�^�����.�jx�t��w�$�0#Uק+k�8�о]���X�]�H�-���o��+����=��Ui���d�N�
�Og�ܶå!%I��be/7.�jr;r��[V/^���}Y��WaU��jвuK��˸�O�����>�\�`��!��'Y�j�޲m����S���YȻ�ޏ�V�w&��;����I�]o��>+{U��Ð
������66��(&�d��mL[ڊ�����^�ޖѫ����ͱ��J���}�;��p�� �T�XV��W1M>�Cow�3�\qX/�������h���R�8c�o����7٩Ės�{A5�cu��qIh�#��M]���,��s4ҫ���Zr�������F"I����t�}����o��AN����ՙ����Z�֞ۢ�Թ�]���&����׹< �:��:�s�մu>ݭ�֮_���s��R��.~���W�Q���G/�C�Y�.ӊ�[E�gc�!�M�t�}��tz���\�:��A���$$�`�Yr�hn�򼱷������9oP�U~��� ���=pi��~�b7�'5���A#�5����\�'!�)�����3tsg���M��!mS���&o-��Xv3���z����ؠ�Cf�]s�{zOw�D�,�f�z���\p*���=�
�� �0�K�e=	��;�E�b\�F�S��4�\ov�bi����*%�SWoC����E:�s����ܐW:���k�r��+Q__Q�ӗܝvt����n��rN�/�uk��ޭ���H��}��S�̽N�E�7��֔M�m-a��š�4	��T{`;�O&Qugv��f����9e)k�c��XX�[�e׷4$민��W��]I̹͂�T�%F�lNc{Mz2�P����n�K�����k>U��2^A���"n�rq�r�_S������*͊u�jǠޝ�-��Cg����)׉,�vӑ���:���}���j��Nvvt:
�7	����&��6D.�]mM.J��{�z��{C�諞��g(�rΉ啳�H�n�#���ϻ=Ӊ���S~�ʽ{��n�4�<����d���g;#�bGGH7[S8��T�5n�ϑ�j�Wc8(�]�L�
�p�j��U��H�J@�B�����w���>8z���Q��ڳ�6f(�Y]��2І�:�a�ikkkN^��������V�'8�;'f-ܓ�G�ǦV�	�剩�J��9}�O}��8���x��Bg�v�}r�� �;���wo9�o[##�l���m*���µ�s��+���̮	�>ޜFZO˽���A:��ҷL']�����:�܇�<�#��Ǿk����(b�:�[7V��P��@�ܪ���(���;���W�Nk��
4uY"n�^c�Zx.�R�B�w�N�]ދe�s�v��s�+_��f�5�є��z��kx
T��oy{�S�=sAm�M5gh�A��8fJur��h�@މ��t���D���/_`�m5����%�Gp/v�f�c�V��ٸ�\7� ;��K���j�5���i��������4�T�h N]���(_&��4:T��/��U�%mE`����vj�2^ɦ�';��oJ暈zh��?\���.��8�bA�e��"�[�-�U�Vvc9��k�#{yD�J�^�|��vl���a�����=C�R1޽<��h��˸U5�Ap���7ev��Z�"w����q�ީ�ѓO����}G�ޟ4�������j���l읏�uv��A���k�x��d�ل7y�[K�K��ޔ�s���Z&^���<+~�5�m�
x��F��u��}X�n
�}�k��t]=�l�͹��}ݓ�?.��c��ڡ3�/j��0,�EOS��"-��R�t/ue�s������x�V�}��7�i3�ݻ�`���=1e�q�3����[J�9^�Xh+� �^߃�`�ֵ��ک�=�x���ݴ�T�Z�.:3�'������Aڣ����-TN'Y��D�v��6o��N�S���,�`[�9E����gT���*�幫�^�����I����ދ�ZY�Y�b�X�����bzѳ�f�����,s��#_*<�.�=0X7�:��
f�X�n�n��&��v��ot��]�~��D����τB^��J��h&�$�����[IT�y]5�ؓ�urlӦ�=-�p�|�e�`��%�"5uho!kgL�yܰur���W�Є1lFNϷ��a�6ף1��D��Z�+�eZ��W���,�Y*�E��3��0�=���^֔�i°�ձ��'$����r�^t���.�T�sͬ��P��8��v����%.���0R�8�9�ӵ¯`R�������v�=\���ή����_f�}:���b��p�͐�S6�t����Y��S�ܱԥsH��8Zgܸ��C�;=r�mK�r.:5U�F6���cw6���֩�z�X�⎎��KGN̢/c�� ������Ϩ��q���$�ش�kT�����܌��1��M1�ȌMX�#T���v+��-�# ���yI7������!A]>.�CzT�,��C)�[��u�ݸƟ��82�H��b=ͳ��<3m��i�����С�dR�"G��38b�ʲ�i��<V�c��u�:s�\��í�ԉ�S�'5�h�r1�q䢐f�8;�5�0���7V�	å��Oh���&*7Ϭ��!�^cjs�tユ����Q�o��Vd]��W��X����ij�^����P*�P�g]	�Z8���zTYw)*��7�WEE���Q�i�u��\%�)p7{^P��cTF���N��ۮbR��2������\)�U'!���~�2q��ϊ�σ����������{y���>���[�2��.��&���A�U#�^��J�DA��lW�������E���)��|���{��o.�߫5o�:�f?u9��W�g��`͒|��B�������K������׀��_�w��ĺ����bTu������2��O�/w�j#T�֖�y����(��6 evg�bs-��Ck���4'v��Ơo������|���������O섟�����
V���a�HJ
*5�:}������
�EG[�͉��JZ5�z�ƚ!a��� �F���M�k�pO�LL?�s�5��@� �$BHm��P(�/���#GF8]��A��M(�rm�����M��S�n��-���5���d��2�![��x	�Q��C�^�Ȇ7
�Щ�JO'�[�O�����4�T~g���
�:�U=�0\U�(��B*
��� I�S�8ɇA4(���nzv(|t�e�C��z6yǚ����(��U>�}j��$!]��b�	U�[R	w�����B�MH{J+)��R��n�m�y�0܆4�ǝ^밻F�2�b���2?��9o�m1��2j@$$���?��}��>�aCa���p0-��Q7]���`k= ����u.BI����wm����$=�JT'�����u��`��;L�����y�j�=�׾�S҆�c*
*6�,s*���\�C���_Z�0
�u�P������aN�������Y7-��ǫ <C`WEz7�����sPTz��3.>���z�,�6r
��� ϼ9d�҂a�Q�*�9�
*? ��P�a.{��%	('��g��6`.^�
 �E���seD���X@� A�jԛh,���d�Q�E�A��D�q��n���/ZJA����Ъ��G�5�J	��X�ɫ&5�� ����wg��&�8(
*3 �G`?6"���uŉ�~��4����:�r9����?�%I��Ѭ;������	�L?�&A���PTx���n��I<P�
*���D�'�@QQ���/�̚�@�_05��秳4�CGpM�w�c����j�=}0*BT��s6m��W��� \1:)�Q��&��y�S�f�l�vY@QQ�.B��`cÂJ��u�]2!߈P�PjvnS1�i
�7�XL�{ȝ��lR �*?�0_&����e N���6�q:���*=c��M��h\�7mf]��1c_MP�Zظ�F"�XC�(��Y����/�rE8P����