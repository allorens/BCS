BZh91AY&SY��� ��ߔRyc����߰����  `^��|�     �@�$�(
YAH�_��|>K2
" D��n��(��B�uJ` 4Jc�� th��$� H3q�QM6�.ۡ$Y@V��Aٛj:�@@Pv�4�0��݊���U��hxP     O�B���Dʅ)H5<�L�UU1i����10 5<&�ISS � ��4   �!!��#T�S��䁲����@�D=	 USBb�`L �&A�$!R���1@i�@ TQeD��5?%?T�OPi���i����b��6��(8H�s	&�HI�C"i�5��1�i� �V$��G)�|�a��������&~֎�e���pyJ%Z�R��H$)¦�7w�k�1�m��pn�! H44��4��`q��E$cm��bG�]e1#�0`����Z�u�Ϟ#��7o�����:�{Q��[��6��^��]�.�c����z<{d5����*r1��i��o���Nǃ�$�<掭�8[��k1��5wG;o��Ŷ�xm��-����"5���8.��(�î
%��b<�7��k9����Z�G"��@�9��k:�WX�b1��sqȱU��9��9勣kN1o�º�Uӥi�p�
໴���k�b���0v��t�ma�/7�Y�G�*]�"ذ��b,s�<M�UQ%��F�Lm�M�*�u��Pݡ^ӂ�chZ6�G��}�bps�;�Ҙ�ts���b�ݷ]�-���w;�xkZ�4-��գ��m�g<��o��n���(GG\"1x���c�k��$5����ݓ:�߳�<�\�#�GC|��P�:��%�BlF����s��I�}��@�o4��&y�\5���nsm�i�ᎍsH�5�L����}$�IIIyRv1����o��.IZ�X;�H [���<�Cct���=%c���y�F#�G����6�Y��q�o٭��LT�B�[B�^����&&+�^�9�&-�n�F����VףO�'mX�D�$&Йo��q�o��Zl�(5J8���b�gSB��>Ǩ^lC���2��=�{2;�w��cc�����pC�`�j���a�AP�5աwH�\g���w��c�籪Y���Y�T�#]��E9���Z-Nju�b�w!n�ƺ�}P}�F��}�A'G�Ic�>�D<CZ5�j�,�)����ػ��b��[��s�օ��V9j��1@s���w��bclGX�1b��s4p�4s9O���G"����'�W��y"�]��,~���������mo��
m>RCv�c�}��o�!���>�8!��d������:�V��[δ�zCYn�c���پ�l��I�l�����
�\��ō��8kLf44��?6��qؘ�uÂ�4-�mb�3��-����B�V�G&4�պF������I�y��y�Y��h���f3�i�C��W�ee���~�Y�'���+t�C�#"&��f�y�m��tR C%���"d'�-�~ާ������Ty��{��zT�+�ú*$%�0��~���:�I�Ȧ���F3;sղI�х�0z&SJ�[��u�iE��+2j���n�r�GՓ�3N��57�0?`Z_S�)(��lv"�^=!a�c+eeH$)��v{rN��~:s}lмw%b��ͻ��Y��f���i$��5$�wu�ƻ��T`�����zWz��a�Ib,θd4���Vcy\�Ǎ�)�b-׹kxWw��W[u���m�^S�b�r|u���+s�7zTE��ڋ�g�����I���¤t��Vݝ��k��H�8V��=�fJ_ry�Gl�v�0):������Ζf�/t�wK����ɗq��s�����w���f�)�(�-+ۻ���L8"�"�����o�'e�ۇ˸rW�&�}Ǟ+		{���<�AB�c��fJ���EUǺ�){ݞu���dm�`đx�e�K�kѴnܛ
)�,�@F��6�L$�n�l��i�u��u��M�	����.�Ԇ�Ӧ�_z��gpa�C�5\��{��/4{ԋ���J=��(�Q$R/��b��[��M�(��9�0�͛�J��el� ���2�:_�3F )O����9 �)HQ��9���N�g	(��;ŤD�c4
A����z]R@1ۺF����s�L��/\$��L4Ǟj�P9L�xI҅Zt�m����N�On��z[����ޟu�P�%�_����D�ۙ�F�SbR�R�D�h-���Rw^�	x�N� l�j��f� e ���*���I&=0��ܘ1���������ۙOF.�F("�L��
ǐ[�����6d���rnǗ]�o{z�y`��1��H�DzPy�'����Q%(P=x1xn�fAI����
A���
ӭ��C%3�1ǹ�<�E�_n雱��eK}� �e���1@����9�9����U�=�%s{��u�v�F%��Y'p����R8iA�a�]tv��;�!
]���/Q���ĳ���/���W��"t��ܓ˯!��Și[XX�q���!��ǎrz	���(E���e��o�"��.�u�����8�*�i�rZA�Ekrҧ�N**+;9�8J',���zT=]�w��#��)�H؜����m�'��(�#P��AUl��siM6�b�f:�W"ם��'H|����o��S���m0�jOc0+_.^�8�c$�u8�U�V�����޵R�L�,@�%fUd��G ������ ��kuTĤNe���PkNm�����T6��Ie���ES���b���V��n���v����^��i$B�A�(B"��A�.��:�jb,����f�n)�����wP���$���U�SA����Q=,��pI(��"P$D2$�0�	��f:}v��&k��s��\'[8�Q�2;�3�F���7���6���evκ�B�P�8� �SXN�bϝM|��!H�뎧sn����$��~ɽ�B� �2���+
+���t?F�4
�\�$��m����+�� ,�I `   F  �W"�8�Q5M(�Jk����!� ��:� �    'ȉ6Җ� ��`��D�	����� � � ( < {�����a@�%��ڕS�$]�M��GM&Țq�`�����4 � �� : X  Q��M4�I�¢�����U>4�|Q���p0�@< D*� X@�@v��aK�jL�b���ΖTJW@��  �!L @` >q$I����M󋊪.r�'9�` � �0� �  � ���|K�\I����s�P� � t �!U �  0  \o����T�9c[��"խ�%t�y'�OH�Bʔ��m�i��O_����4;Ӈ��y��y޶���r��ñóUv;�c�
��U!�T�j+V�Z�y	yZ��B�����Э
!D(t�H3�F3��Ph��G��Fs��mqXJ��v���K_��8�-uȈ��`�-+���iS�J�-���|vP�TnX��Ə[��D���WZr��@������2R.�a�D��H>��@tp��� 7��P����@HR'&��V�k����"�ۭ�*�(�����*,q����1!Ny3y҈�g�wG����9�����b@��{���$��{���B[����i�{���	����`�����
o��'�!߶J���
)m�\۫=����lFX��E�`�/����E��Di��/�D���㌒G@����^�N�f��q��v#�⯛i��Ň����Chu��$jn9��7��lĎ)�Q �kf�(4A���gC���d�U孭�\.8�`�`67�jy�31����t4iEkHl��{]8a�Ä�7�9J�.���߻˵R*1Y�h�����<�ί/
$��B+F��Z���vS����D���r��-ZX���h�la���6l�(��j�T1��خ.�Gj.��{ʷ�ޘ�#pT�l�-m5���뛫��M��*3���,@l�G���gy�M/mt�zS�g�����!PRT��V���鍌:���I���h��Y�B�m6sJ�F1mT�9MF��Pg`ڌ��7!&+6ֹK�4�����p�h,�wܞ�f�.��:��]�Z{[P�����U&o�J��H�b-P{Xh͛],�d,,���~�^��m�K	Hg&>=�D b�R��;͕ɨT��]�R�-N�d�Ҁ���8 x����8�Z�v�����"�J�	
�t=�b�b���QG����Mt�A�m�&8��M�H�A�K��<��5lf*��7+�l�o�q�l�&�V������s�3��d�apՌ�ī�v^�1٣:c�Nc<'�#<Fx�$~<U�"����G���~����t�M&ǯ���g��	��t���<3ǉ���,ٲ��4?Cͺ���(�~z��>K?tľ��O=�굏ӭ��B��9����N(��}��קN����}��i�g�|4�E�k�b��_uã@�f�Ϛ8���� �[l�m�s��m���[l�[l��X�a�(B ��	�I�|�KHk�@�i�Xh��?^b�i^�q���*�t��h�R�Km��i1��0hk�m[�4�^i|�kPٳD,�����G���H��T��KI��5߆�M�ZM+�")����y5ƅW���b�W��f�0î!�\`��y�,�D^-B��P��"��d�����l.؛Z����I�*R;lTB�ˎ8�E2��A�m4
����Ziu	��.�G�[h6�%�2�+<�b�%��S8�X�'ϕTD�m���G���M"Ɩ�0�g�x,���E1��"G�F�J�,+M!q��܅b�L��fWI����F��*��!��4���0�xa�Abf���4��1ڣ�ƩD|��a��6!U(��q��)�|#�0�@�`Y���4��&�6�[�Q1��A��J"0&�gKcl�q�b>�#���7�l]Mc�鳳���k[�$�lҥG�X<(��܌������1M@ �W�,1��V�j5 ���&�K�� ���H��4����:t���ݯ��\*����+��T.���΄�xǈG�ц	L����шh<v�D��$�LFƊC4ma�n���m4Ah6�h�j�����c����zt�\p�ʑ��ҡ�T��j�"_��I�������i���V)�qiuZ,0�c)!����>"Ѹ��D5a�+,JR��.P>��G�q1��33�Q%D�'�+�/��R���:���l���y6S-�N�FҠ澥�t��A�/�5�nא�{�yR�����`rqQ�!@ΩI���E��1�Kk�M���fԪ�v�cH0�G'j�%��/U��:1�����J��%�i����*�D�t/�`yh�Z��֟���l�aE�[�eLz���:Y��<;��?���G��ϓ���>_)Wi�^�S����6�����vlƭ����a�����)��|3��xg���G8l�<L(�+�"�3��=Q6�P/S�`χϋ~x�1�H\!'�[G��fkH��-�DƫcR�,��yU��D<Fdx�C�����.I$�KW�L^_/Z�P:�$�10��H#�n=�o��U�춪�A�BY��cq��:`��0APB��t��&����$ j�e�EeV�Q�QG�P
�4�㄂��4Y+��HP�T8d�'��r�l�B,���@�U$,���~���k��r��m��[l�s��-\��j�!E`0w�=pȄ��T��
5mmV�Il2���Ꚗ�F��*�b��(4���V�(>^������͔KDK�P:��6����<i�\8S9�!��`ak�keAĔB}���G݉Pi`��!�\{{t�Ӵ|�����Ѳ���Z+j��=աY����0�����V���l�).�9�ç]�R��u��l9񊍰�0��w���,�a@񋔠ύ�F��߸��5�y�+j�N�UWwWΛ����x�u���6,��Q�1��P�>E�B��3h��:a��(�a���C����%c
�[e�Ǫ��i�i5v�5I��(܎�$MR�Q���-#�1�^6�M"���,���QEX�(Z�Ҳ�fc���mh6�����<h��(�ad\�� �KG(�@v�g�b�!���V,,g͌�\6���\V>1��[4/&����TۣK)V���
6v5�8���i&y& <�@ ��qy�a���T�]Xb4��f��(1l�(;x9��c,"�D���~6C��(�a>��&8��鵠�F���7#�v�BIe�%�|�!�6�5��}��F�ë�!�Jx�&�Q��k�_aQx��D:�E�����xw�k�>����KAW$NF�}˥a�P��Kq��+ՙXѺ�b ڍ̱��+�%�����XgW����(1�j�z,�L<5���<�+H������UUZ���D�!4vLQŮbn2�\j �|8B¶�qkV���6��*G�EXe$`}��;*:��m��J������E���ctBϏ_qEu�����xz?e�+���¼?%�ɻ<S4x�x�$~0�6E�>4L>'����3Q�='M�|p����|x���߇�7����d�x�?K����Qꉴz�z���:}�{�Ϲg�]0����ȵ=���[�Jt���E�n�|�����1����� -��<�۔�m�M�ܤ[m�m��m��B�c��\b[��"�P�B���?���V�����c`�H�j��ťbz A�������T,�3G�YD4f�Ʉ�
DGÇ��"�٠�m����,�b_+l�ZK�V�԰�cxaaŮ���7�6��-��:U\*���KW���׿5���-��Bj����[��J�lv�v��*l�Q�$NR�TV@dQ���|�ȕ�M;\�e�b2Spr�Y�B�~E��i^yg	)�:Ll~�͆�-b�����n�WFC�J!��ti����7k��-`}�҃�"�H��}�m�&�^�8�8T�����,ļ�w��og�0���p0m������"]���|�)�G۠���gJW��(��!��/�ae+���V��iWQ��ύ�,�gEm�f���\�A�?9m�m*:�mZ�m�e�f�t|2��F��Ɩg 客$x�F�,��{��}c�:m]ymr),i�����T��3%bKƐ���1�f��:z�=�x�pm��F�>E���نU �D͝c���ePJ<a͟&te��͜,��8��ȝ�t�F���IhѬ��$�Q�uU�
�Z�0���9uTʧOV�rʺv]5�D2�cgrƏ��+�
41���DR,	`x�H���F"�FY�Y��ލ�l��3^IuX�^"�(�Q*F�I���(��`a̓c��*󄈓��@�N�A2t�U9[zF-��V}Fp}�#Q�1�+�k]4ltYK}�~Xu^^�Z����"�kݚ!Ѭ1Z8��!��m�=)��4}zm7g���Y�^�+ǣ�,�C��)�<W��*͐���x���!��=�d��l�t�V��ӳ�r�J�z^��Lr�/K�t�H�5�z�
�QQ�����(���0������t+�l*�i�Ӱ=�n=��תklCP��z�&�iC�#�ej�_L��1Ĥpa�{V�8vM]p�T��o@-'(i��.����f0�������-H������A�"cMK�U�d��J2�P�;uU�r�q�r��c�D�Tإ`6�L,i�5^	�ƭ�KP2Kґ]��Nm�M�hF�Z�㋱�.�Ow�v�m��r�[m��m���h��h��xF@F�=�d��$Q"�mIe0�H��qI(�-e��ƅ�R=X���6<��9�mC8����0�_�٥IT�F�(�#g�H���)���QhNܐB�@��@����".�m֑c:x酌��~���#����5B�Z/G���l�㊕�(��>P���se�����_��Y����:qԶ�c�G-�4V�Ep���imZ�a(�le���|��!%:�#�F��%G�2�i�������G)Y��Å�i�>Ib�l��4k���#l��͘��(t��"��M�5��8��ZM��:�6���t�qE�gƍ&�Qt����6�rhH$j	�ID����wG�F�c�Q�؋��GU"�� b<�H��n�+G�4�R�>L�_4P�V���G�uER6q\�<���f(�t0�ӱk��ڳ�[\>��Q��m�Ρ��zG��|1�����:Σ)��P:�XbƏ���B�e�����(�h0�6��IN��9�Kh�Gˋ
�!��$�EV:��:�����r �� K��f��x�E&R"�(��R�l���%6�,J&x鲌+�x"kGǓ��u߆�P��Y�F��Q㣳��4�1�:�wpdH��z��KFmt�|�"k�8Q�,����/O��i���T�L�Vժ�R5S�:�r�`EUMX�;X�ɺ��}���ϸω�)�Q�lm�h��ݪR��Řt�����---�� 	L^f�b�Q:^��^(�����\11p�lO�48�D�B4�qi*C��f�K�ih�Β�[)�R|���s��s����r8b��b1bŸ���<�4d:pLc�ppl�0������x�¼x��	����p�<YeY���%�!�輮��zn���ݎ��X��eӳ��Lt�/K���WwN�[�MN/�SQz�G���D�Q4��z�����}�揓�����;��@D]z��.{2g7�m97�����=�g��_�[m��m��m��m��m��m�ۄ!MX`a�W�!�C�m�Z��f}�p���GW��j�O�5$�K��h�tţ�ŀ2���ʈ�o62�h4o���w3#N3�'���Z+��L]����-�;���`������:MQ-4���i4qD����f��V��T��Rb�W�.%ĵK����N�Vmک�Mj��ʝ���th��&�{j��
\�Z�K'KZ:�I!Z;v�F�bkU�E��f.|�c�
J�E�o# �h���aҍ���b�0��"�0��f&�"���V|Zj[C�H��m4�g�=�l��00,î=uѡ�0n�t��{�<W(�7��v�������^����AD:�-i@�>���f�ҏ�c*_R:�lÇK��u��7�1��~,��ߗT�ڵ�k�j�^7g�&~��m���k4�~-e���F�Ak�ǧ喙y��۹h,X���r�au��4֮5Iz,����^,Z���b�d^!ӊ#�G�Y�lr�uZ!�fժV��g��FiG�$o��n=�H�������L�h��k�GȳE(���h�
-�Z��<�$�.o�4E��QV�P�ma��5�FF7Z�x"�E|����';$���K|T_�|nGJ#hŵ���G�՛X��0]F��z����,�N�1�}Ě���T�<i�H&�5%Q�i��4��1��|w��4�#`ހ:����R)l�MR]>�Ms���G�i��im#K��ϊ�t����=O����htx'��g��ǩ��R�a�����?QP�B�D�q�˦7]����7t˧f:^U˦:^����<>>��lgŐ���<;(��dO؆#�!��3�p�#��wP�,)��N�3/[h�����~���9��"ؚ�6����[M���la�:X���ֹ�K%�m�뭪����i*�#�9Ca���B8K��?^s������M�I�3e�`�球޾�}�H=+!�$�f;��P3�elPB2��26ԤN�
�ơ�ty��[[nHFh�V��+��J�$g&Z��Dǁ7$�D�6.+�4�O�C��i��g��m�M�ۖ�m��m��m��m��QE ���e-��mPq��$$���"��94�t��K�)Q����b�����nġ��֏i9��<���#�*�%��24ƣ���$�eX���p٣��agr4�z�k��e�FEVD|u�~\������*�|�F��Tm���(����X�p����ϋ�C(��akJ��j�qDM�ː͵8Fqi��y�ZF�DH;O���3�o���ÇǍB��Q���&(�����/Sla(;�qu�Tuf���ix���@k捖�$�y�^6r��� ���M~�H:����w�$����9���;���C�����؈��0����1��b�4�yY�K�k���F_�h��x��
�m��_N�G�Z��pi�f0�5p��ssF�.�ԆiQ�����v|��G�����77�8`��`j��y���*�_$�8`l,߭
�Y#��|F��æ�c�].�6�g�o��4�#���6mqk�H:8lå,8h��JȆ�(qyp�>^(��Ը���o���Z6mH�y��m�L��7����0p{荂4D�
Jj�VD�"��6��0p�qZ���>�[u��$�G�<�&/�=Y����)ﹶ����/t��2�,^�G�����t�"��-	�W$�z4h��1���,(��D1�G�Cv�r飃Qt������w�?Q�m^��M�x�IWދ�{�f6�,U�t
�s2b��/Rޱ=yh�����#��tu�	��?�+����htx'���!�ģǊ�F�vx�0��<��Q6=�&���l�Kì^3ռ���W�Lt�/.��x6O��c��/�!��d��g��A�$�|����?.�;i��5:�ڎ8�B��v�w:�����>z�m��m��l�[m�m��m��k"�(���?�X�z�[�K�k?��k��*���<�����ld=u���.���_��0������3H�\\_t��8p8o����Vt�llzD�'#l����8�M���_8��b�O�uu��N�$�M(`������\�_aKӚ7�vݪ�h֫R��P���c_gQ�~�/�
�h�k��E�0>�`iq��ܔ�۷n�H����Ce���|>�y}�p�Uk`ژ�)�b<��mE��1�m�6�9���ȇF�lk{�O��G�l�DO�cv�#K�GRVt�ï���ވ���)u�*^M<N׼qE�1�#��8AhçC��S�?�ZF�>�>�>��,�ID�Ԥ{�a�im}�jыKH�mpKV��L]�T_ �����-Z�\KR�w�^ՐN�\��U]Mբ�9Y9�80$ ,��Up�H��+)ͺ���66���%�ٲ��䬚Qm�/t��;������u��\r8�D���1�(��c��ߕ+0����P������9h�^+��T��m3�F��K�-qoI^A��h�Å�8Q�ꓦ��E�^��t�z_#�jvG.�c�U]D��>>l�m+K�Ttk��N�Gt�Z��E��COM��b�1�1ҵ�)u{R�9K��[N�ѣ��:�|7��|��6m}��T�oȣ�.�]�ԩ�CDc��>(���G���<?G�:����<Fx�<J���`��<a<a<E���0gƏ��|t���y^�˖�N��yt�+Æ:�@�D�Ȉ^�O�E��*qD�^����㮯S~����*�����w��9�p�SrBZ�V�Yp�������KD���U�ӗ1���s����f�`�(1��՛��	NOQ��o�:��I�vk����{�M9C!S9"��@��U��JV�����d��&�X]-nU�_ѧmX#hȯU�s��:W&i��"�A�:�9�=��#�m�&Φ�\���4��ZZ�dX2�dq\�E��V�lL2��r8 a��;�^���m��m��m��m��m��m��
0���d���sf��v�)�]V*�M�f�[HЩl���
H�#������6G!>K�qq���64om����/-.��T�p�\>�χUR�u���x�������I��I��F4WWXyiCK����zj��E?��]F*-pccED|���06�t���Q�t�"K��B�W�$�ҡI��TCip�p�6�ŕK[�#�D!��aGƪ�Z����!N���T/=ŋ�`߳�P"�X<��|qpf:`p(����i�iَ�k\�mJREC-q�ʜ&n�[��!n�q� �CW�j�.-�e�֫hg�gȵ�nB+�-v���T��A�y^g�aȯ��)�`�t�f���H��)�l��R�K����[�u@�<qx���=�bmWE����F��Y[z����[fܬ�QP�q,�ё��m��ul��mCE��lÆ�晹�9F��(�k��@��ې��{ךl�>>�T��Ά��g�c�kK��r�1 ��BQ���}�[����E\�bk��M�WQ6֬�J�lq��f�Dq.���R;X��qF�^5����8bw�@�p�H�	E^�(6A���S�D�c ��D�Q1L{�M��L:�}^[ڳ��~ڳ���JKL���uv�
)%��^b�fL\�;�л�=�}M�'N\��ӧ-��;0�٪�$$!4!R!.�BP���իV�量<l�㧎�:t��ǎ�6h�x��t�H3�Fp�������0gvO����\�y��|xUO�̹�Әw=��G6f_-��z��$��	$�V��I\��LkL����U�P�Ƒ�<<SV�{3< ���������^W�宕wH�L������X+���hYի�倊f��(u�Pɧ�t�<����T�����j�� 1�����^����xp�Z��m�{7(}�"U9\0}~�,=�b�u��/b�ۺ�9���z3T�<�u=�3�ztz���|���m��m��m��m��m��m��X"� F��BOG��OR�о���&W A�u�g����6R8��+�c�7EgS��4��1!�H3!H�F���#GH��&�m�,�F�#i�j��Y�m��_/*�z|��JϏ ʽz�ث�D��R�8�:); J�U�h� K �I�%@�lpt�"���z������#���Q�1W���ҵ���p���{��P�#-ql��>O���l�Ҏ���P�>d,zF)[4C��|-PѥT��*5���Sg&�$ص��jǘ4�>o��|��aE�z�f�J)� O�-^󯘁Q�*��a�t�yqiD��wVu����l鲃����-Q�-�h��ӡ��m�h�:��IJ��S�g1:<ZGx�4��5�6V�(Y���зޯi)�٪ ����c-�}E�-A�*A
�dDlcN��MQ4�2���@}FȂ7:έ-F���˞m��Qx����[IS���|���GG�BD0�;v��l��-,�cl��
�lڣ|h�r1��:Ck��Ǜ>E&�[k|Z����A��'<�n�I�|B�;�^��hM�x/gN'  �(����Z���m5GV��T�Qe��2��2Kp�CT��4Q+��c,H�V���g�G.T��R��g�Ů�1��M�/��:���N�]���[�e�5?/���"�źZ���-ŵj[m����1$2�}��=����4�c�J�ww�e[a��ff���"BhK%���v�LY���H#6 ؁�!�-Ke���&aK*`�JRRȥ
RR�����i1$�IK
T)d)R)H���"�JaI��X�X)d)b)D�IJ�R�LRb
T�T�Y%,��"�JX�R)`�)1,�)�)QJ�J%,E,�JE1I�b`�)d��K(R�JE*E,E3I�)R)dR�)H����J���&��%*R�FJK)�FQT��,�U?�*�),Sjk��*��--���l��e)1,��l�Ģ�e%�,�S|���J��QV1RbQT�J��U0��*�K(����3�*ZU(�-*�*LJX��h�K3�4�Qe"ŉ��%%�U,��Vpf�1B�K(�T��Z���1)TX��YJ�
LE%�,��aI���B�$�B�%����*�RX�YER�*�*UIb��(��T�T�R�K�YP�����U�>7Wk�[Se&%)VUT�V���*X����,T���X��K(T�)eK*T��)�)eZE�h���-E��)e,�Z����T,�W8�EU�)e*��UB�K)b�T,T�������R�e,�X�eK(X��,Rʲ��YR�,�*J[m�T��JJ%%��RX))%%�))�X`�
--%BŒR�Rȥ��%))d�E))��L�XR��
T)bR�L�0Y%L�cL�J�,E,E*IK$�
RR�*IƽF]�
0?S�� d?K����H����(��?���EeDBI���$Ɛ�����4"%������k�Y^z���xQK���zJ��"��{���T1�I��:p~��rT���OH�uy]y5!���XlFp������:R�JY�f�	@�m�o@�&�Ǉ���DT�z$�T��Ӈ�!!���~���/�ė����)?Z�$�8G����U! Y��T��i����ԟ�u{~H�V���+r=0��#|*.1�K
�πJB$e:�>;�!�&��)x��0�s���7��?VX�O&��Ԫ����49��Q�D��z�P�'��K-���S2��F~N!�_[D"$L�M�
RhS�s��D�W�c��=Ǫ<Ìy��Xҵ�f�V[�\_�s��q!T 1�9�!$L��}SI	I!l���!"$'�$�$�4���&$�i1$�M$�1�F�IF����(j�ƒ)R Sc��6F2bd�}os�j��'R���M�J:,�@�HF)THZU!-*���RDLRB-�b�P�/3���cG�<�_��;Ѫ:9y�yI���~�62�f~���l��X����Z��	�'��<>
�����g���g�Tu����{d�+va�L>	>��\7��F�?7�n>}<���ß!z6'~﹞�$�{>z{�%qi�_�5l�T����^ҍh^��"W�s��B�Ya�3H���A!�w����H��It�	����JW�yX�����wd��>��0�EW��O&�"D�V�DH$?�^)���O&�\.s#œTt��d�]�B�苤[C
4 �ďтD���<٪[��em��>Vu��GS$�HP�G�����9i!q���(MpL0U�DA�h� ��	������^�H娴��CTe��AlKH���c}�����'h�H`2OC)]*�̽�k��zRi��	8���U��X��T`��IsK�Sk�v�������`_��¸��	�H$$�H�N�I�>���t��N��Oy���(4{w�h�9��dp�`%��cB@$�#6y�����%VmX��ğ_��Gb���H`=�M��^�a��Ǌ=�����M|ǚx#�n;C��E�J�"���F�/bm�UJY��� ���`.u0�@�$��D1���#ã�Z����<���;�٫���#T�F��<���w�nx�D�C�jH�"����hΉb`h!) ����Ğt�l��ߺ�w99�����9��O������lzyj�0�p^0�y(��J�t��Z�I�*L�=�A��
���5H_]����s�y]�H��~W��I�N�PA��$�>*�u�%�X��tT���K�LڈIC��\�	��]��B@�+�