BZh91AY&SY�b|�_�pyg����ߺ����`�~=V        w�@�P   U9ƀ   4퀭 h-�HZX@  9   ��큐 �0�          �� �jz�on�n�-�+�&����������y������{{�����]�M]�������k��w�ֽ�vs�����w=��{w�n�eo{ޖ�f��7��X ��v�z���m�ǯ{y��[��:���VG�������n��i�n��Q�]�h�=�Gyv�Nn���o�g{7�[y��n�]յ\ۀ8�` ��7T����{���z�p������޲=��u9�4om;You�g�C��(���=��yx����ݺm��']�w�Op;�\�u�3�n��xx��  h��3�mݺfݷp�v��v����}��۹��y<#���ι�.vVsuswm�W���s��m�����׼� � �x��g����˸z�koN�n���w7 W-m;xO#y�o��sϾ\�a��hN��U��n�u���                P@           �~����JR����@�h24�A)�����&�� 	�CC F �Rj��L�2a4h�&#LL����*j�&F��CL�h     $ �@!�a2hI���m�zS�'�@�j�J�F�0 	�b`L��g�����@}a��xq�� ���A� 
!�A����/㲪��H���'��/����������������O�lT���6�f�ͻ���P
��'���UU�)��gմ��ڪ����ޭ���A9�G��s�g����{�_ؿ����U��'�?Q]9{'��88L4�f�&��w�^��>/��i3i9��w?<���9�q;I:�H;�3��_%|�.�!�5'*�ލ�I��A7�17ӯdv&w�N���Y�9 �d�Hq�q$2�3Bf�0�xɜ/��úd����|o�h�d�&�Z	��(k$����h��i���C�Z��lѯ�&���BkI��~���)�$G�"��u!ߓ:��d��1�2D��&Ӧ����N��):�w�|�a8s�u�J�I���hJ1�p���O	����I�l�d�ˉ;��������]���P�����8�$(���Nm"hr:N��e�'��DI�"k�e�D�'	�+I)�Q��6�L(~�-,N�
/���:'�ȑ!��"t������|�Y�K���1"$�L:&=&q�>Ft�h�$D�H�JL4k���И��K(~�	z5����%�|3�M��H�ԟ'bK4;��0H��&�'�tH�3I�I��gѲ}h',RQY�ټH��9b2��k�3d4��I�'D��a%��7�H�ٳE�}���&m"u:)�Np�3I:g��U �p�Qr#ܨ�ؘ&&����<����L����o�5:V|�)��w�"pnpM�F5:^�ܳhfǱ![���9���DzH�d8?Y�M���M�|��/�}�<���}�ک������ԭ���i2�N'(�9�+z9iX��+�d�ߨ�R"^�Mpg
�D�D��h�����.�GS�z`���^�~ʖi�=��i�=�3�ڗq/�j��N����d�5ek�j&cQ5r8D�ESR���\�\�*��9&:�DG�b>L5���""Ŀ��}s��TL6�X�ʈ�8Y�}eTDwuChIʟ#�����DdL58A��"�a��G;Q����R�u�&�#*�#̨���B'*l�����YfT؎�Q0�j|�$�c�DG	������"/*'~�kR��K �|�i�J�Q�j"oMJ ��#�TD^T�ڈ�ϣR�9>DeT�c����*"qʖCZ�"9���ѝ���jP��K �|����R�u���Dޚ�A��GZ����B3�3mK ���Y�M�f�5"7��DV�s"a��1�8Գ}�Ϲ�����]w(�9>N�Q�vPS>���O��FP�e�;�9D3�&�"76#̨��`�,��gK��:��G$fT�u���2"sMN١��O��v�B�$�I�$%�>y9"Bt����'Є%Ғ����e)��V�����9����p��(~���ӵ0F�Q�+���t�Y�J��J�ΝgM���rC_&�J%�}�,��,�Y�C���TIQߚzp��7��u�:Ùa�����Xev�v�wR�'yl�m�3�2�C,�LE�j�{��T��*;ʋ�lӪ����G�ӑ���c_lk�F��k�}���Wu��{$w���n��TyjWp�$FG�9ƣ�ԃر�T��*jeNI[L�'D��p��-ʍ�N�oSf"]��V�u>rt{o�S�s���C�:�Nrg���}�MeTԓf�H�w��2<���̓⋩R#Q��=�D�u����u�fgY�L����ew�mc�i��淪��UG#�QɚjJ2�γ��!�K�Xnw��ɾ��rkdvI��G��eGs4�ʝ2��S%�ޣ���Y�\�}a�Cd��Ragsl�,����N��|�L���d�#:V�O���>��r	�;��vJ��3��R(�^�W6L-��BtI��:qɻ�i%���a�:j���bpG{��ev%�'F�'�����ؗR��*�7	]�NT�8��벾~�*��&2DG�M�~5C�k+��,u�_#ؔi�P���2W�ߑ5����Nr"�W���+biܤLw)w+��JD�2�h��Dy�VAYD~�K֥"<�C�O��R�4�R&?DEԮ�:�_?<���jU��%"me&�a)��|�R&�JDβ�h���c�J��eY�O��JD�]4:�}ߚ���r�1�".�t�5�_?<���jU��%"me&�+��ܤM<���ep�����hy>{:�֥h�g�$��";�K{U��2�~�jR�W{/�;�T�t��9%���Q��ȘlIؘs��7��7&Ʀ�H�B�ȎL5؛gM�H ��_?,�(�j��rN�ɱ6�WE��ea�Έ��gMv_'Rvf�l֤����b?p�,jX��$뺮�p���MI�ڔ�d�-�~����"59��$E�&��U�U8�<�B�:<����D~��CL�&vA���<�s��������9�D�g��_��pL�\�t�:j�q��F7�s7+m���]��-���Y�*��Sr���wq�yw��I,�p���T�'nV���CJŕ�2�k�T���nV�*s��Y|�&�Ԇ����q쥘Z��̭J�!;�͹+i���ǵ]fƫX�V��$�Θ���vf5��#Ѿ��Lp����=T�.t�;�Y�o��&CEꉨh�)T�Y"q:�/I9�xIu&tⓩ�o;&�5�H��3GN;&h��Ζ���}�XK;�V�P�>���Z���Q�B���T����YO���cE԰|
X��fJ��B��A��������U��IY��7�SH�a��4ӓ����Q�`��k�$�樚J�������99�v��{��'�K�5Lx�y�$�8V�	U7�V^�\��d�I$�l�ԗ���u��i�7�K1/#�aT�)�r�9VcI$�<rާv��J���(�Z��==z��}�w�D/%��zjK�� ��q:�[~�]-_E�9�ӵtua�̱l�U��d�>��i���|�%��y�?$��y9�qq�W��Ɠ�+��$�L�t�}I��u.!Ǖ.�&�ۻ��P|b�M�kI�r�G�yy��Ȼ�_#�J�7Wb��D�L˭["NȔڭC@����V;�FJ�߯>�)�,K�"�U�y����ȯ�}���V����#=�گ�7�C����������G5`�h�����K�ի3���CH)�Y��]��b�Jv�r�Ӝ7�O!��]��}���Uz]�b�i�q%��H�[��e�����)9US�!����"�H��d(N��T�jr7�T�����W�if*�i®��?N@Q쳫}x���E�򣱪��i%ݳV�J��b_.s�m�yN?w�4�lVV+���{�/&�K��K&�U>���pz��|���l��I.��x�bIE��6��R�I$�JQԒ���ʒ��W�ҋ���-M%��ݚ�%u.��n��U�VcU5TQ$��z�*�{��s��o��xqr&��'��|�,�/&�I$�K5T[>s���.ؒK���Z]汽I$�|�����ID�K�ъ�;~��$�Uu��&��|���3�*oӪ$�J�Ə i$��߹|��&-G��I$�J��R�RI-Z�^_.ow"I��H�j�#;9�#��3E�ih5�_��2Rn/��Ց�1����9�CzL:�!�>�w�3�{u
�`�u�,�RS����3��B����!�g9��4��E�hv7�G&�L��JB|�v�'�ۤ϶p��ّ� CFj���a��0��H�zL"1ɐ��<,�.�G���	f{FUݤ�[3̐a�SA�&��J2�Q�r�"X�E�F�*Z,�%�0�%�#��}H|���G���ţ�2�=��ތ7X,�[D�#+{.�1zY���3~X��5��L�y�fyfO�3���ц׊9ך��VHWt�H]��Z�	��jҰ��9^$Z��$r1��.!!,x�ȉ�*�̐��CY� �$}�AY�f�=���m�9ׇ4m���9�8�#���ƚ'P�č���"m�1!O3��7�RjĈ��x����hӇ�sh��Y�%ՑbX�%�����-��^$[I���/�3�<�ά�,h��C�\H�<H演m�����VyxYr�l��cQs�W�B��b�j�G̨\y$>��N��.�K<�°��H߾'��.${�Y���2�H�0��y�,՞�h�M�$Ch��4Z����{��z��Ӽ��NQ7�G�[�k;ûL���k���J��'V4]X��R��~�� �ϡ1��	��rtu�v,�*X������O������<���5���Vh��wش�gV%�g�$e�3�C�"ı,\��Ļ�='�^n$�h�J�RZ���,��eIR
��UE����s�21��/e�q��,K��6�h�g�>#|��:�u�YQk6t�w
&�bk$����5��eTȲ��S*dnU�YRT�SBʒ��*Jԧ��d����KE�J�X6��o�����Y�`�y��+��Zĩ*J�0�Ưc�����ܭʛ���*p]�!�-yV?"Z�sH�&6��kY�sn��:6�,Z6�w��"Ʊ,�Ʊ��bGF�DAלX%�5���Ց���7�ۤ7�F�49�C[��M]n�p��CyMi5��o��/P5U��;���Y�:_�d3�mP>#/KeISF��M��H�sNe}��J��\��)���2���e���22TȒ��fL��d���\-aՕdG:�T_3�Y�Y�\�ǌf�	�]yŊ#m �:�����t��5�M��{g�a��S��b�6�`�=��oVj���(��!�h�<�]qa�9�w�fӊb�H?�$[��#%`�H�B���#��C�8���V-C����O�B���$���Z�oB�̅���G�����:l�_f��^d-�TH�,H�I�=�h���p�أʈ!ZMEl^x��Þa6����,~4f��E�Ȱ�Ȩ�^q1׋I�U��K.9;��ȡ��G5���O�DF��^��ucE��Q��G8��oY���bL�	�
���>�5��#���"X�Dh�
�$w��~"F���Ď�Bh7�"ʍ׋�![�˷ �sll����D����W߯�]i��՚�|��%��N�΍\'J❍�j6b_,q4��N}�>��c�-_O�����H��V?��?���O��#W1�O���|�}��!��O�)���?Oӛ�lH���b�ͭy��֬�s���tԩ�fV���V��u�Ccy��w�=�jq�vso|�\�g�U�z�+��QVD{�$jC�^�{N����C�	��nj8�#QQ�w����B~��y��M�5W�o�X(íY�2V�v���x�
���Vݜ|�#QQ�3��Ҿ�����U��ww�/�.cF[�7�9�?{}�T]}�Ë�x�w�cA_(&ǣ]$m���}�ը�]�����Y���ĵ ��6��|�����߹ā �Ȇ��0Չ`w�5��7�}e�O<�ѝ�8�	_z^ww<P���������u��wI�O�x�M6�j�{ǔ�Z�,9����p�o����k��wX�؃x��1�i�C������J��U�,�px����{k�X�ؗM�9ol�u��Mf�G��&�]�D�Xv�]e���̺�q6��J�;��u& k%a�*��o�1����#l5�84(�x�#bbn�,�,�r�aR�C�"9$�k"6��sbPRR��!"V�emT��Eyj���^��s���QÎ6Yn9X�*$n���1!�T��Y�vXAY��Elۉ�Z$�[������x�,I
R<����_n��J$dA(�*��U_��q��xē_'<�H�/M�E�fZ�%ZY�=�D��&��Xy,J��8�,q��HrTc�J�>oSך��,(�,�)�3�|�7����ĖFZHs¦��Fab�a��2��E|���`�	.h��)��|����h�b[��+5$\w!(ˊ�V!DK�@"*ԒO*t�Ȯj�*%X�\D�LJH��B��X�B+��<�r��5n;��!B�A�A4"�B$HD�sK�nR�*@�+�̅��p58�em�#�x�#-P�����r`���X���1<��{^c[�y5<� ��ufM�טel9�3<�V���f|����@�֮���_��J��-7j��fր6���m\KI 9USQS����I���qg��2>�|/������1�rXgk����2�9�!��"�jT	�p��qY������,�Y�[Y�cEF2v j�X��;�%�A���%A��]A,@A�w�k9�P/�L�Ϋ19x�$KKGR���yjL�nj����ܡ���~�b��U@ ��;	Ο*���������-c�������}���_�/��2��YUib���ׯ�����s�X�Ux������X��+�U�]���iU\WJ�j�U[Uڮ�W�V֑UU�U�t��Uŋ��EUUEUUV�U⮕W�Ux�*��iUy�W�B����'� |g,r�m�����[d�*Ȋ�%EFE��T�*��ڮ�]����U�iU^R*��UU�Ҫ�����*��iUW�J��Uv�ڴ��UW�t����i֩U�Ux��U�U�]����Uګj�j�U[W��r|�|v}�!��V��˫l�0��[C)J�
f�9��ګťUq]*���Uګj�U\EUUE�Ҫ������������ZUWҮ�W*��Ux����{v����Uq]*��b���Ux���ťU^=>;��Ͼ��'Ą��|HI�}�V�������*��b���U�t����]*�*�UqWJ��Ҫ�T�Ux�UW�������UҪ��U^�����U^-*��*��*��*��*��s��9�d1�A�$ 	Y��96
3j3QM��0�\ƣ|[[o�wn�(�I �"���|ϟ�?j���0_��6��ү���V��i�>��>��(��4}�	�N��:'舉ӆ	d�M���(�H%��:"c"X�blК  �DK:& ��"%���N�d�F�؛blК���6!H`��lK�١4C��(DDL�,��B"X���'D�bY���hAA�u�Ye�Zu�\�5��U��|��Xe.�sꬬ���d��Q?�h��ܪZ��iRF��!\#���)X��+�R%q9ju�����d�=՚-Q���mRԫ��*�ƓlE�Qڄ줊�b�U�[L�I�%�
�J�W����	#�Q�3wZZV�労�N���#��S�)M���6��ob��do&�1�ptUH�:��b��cXڄb#�C�D�E]�<YU�Rc���ZY�	+V���ҭsQ��H��YQcB�J��!'�V�uX�$�V0U����kdO$D�N�\b@�i��bZ�z҅������)%r6��MT�*j��TƘ��u�'YG0c�ƠH���Ċ/ƹ�[!e�HE��6��֊�4ӄ�0NQ!epMҖ��h�%��4네UdHtCjV���u�`�N(�n����S�ԍf���1���M�i��OThX�Kl��(�v�!��Z�HR ��6�8���X���l-n)�s��j�Ǣ+j7��TQ�AK2O�!�\dU�X�%���A��
RDB���6Q�CHI�pyISX�"�e("��0c�$"�
��!�A<,<PX��Ȅ�CՅBex)�`�Q1�֐�1����Dlz�L$L����J�,c��`�G��DId�o!q
NQ���&�ǣC����Bttk&D*F+[��$)(��4)GGc�A�q��6�o��%F�qGDR8ZR�xԥ��1Oc���i��	�$JL�K�6d*)4LC).!:6�JH�B
��t��"��	�<9�-"J�e�.Ad+-ɐf7r��ii���!4mƠ�$$WK�W���B��W$Ǆ1��Y��(�B���#�]2�"�;��C��E,Ce�tlx�pd.Qb�Dc�k�,g����q�t�5��ˑf��ǔ��8�.,eD��	DD\���yL�CT�-2�,)q���D��l�HA��q��Cv��	?p�PҐe���!�Cr�L�$��B�h�]
���J�Sa�GA;-,�x�\��mJ^��)h*�t��,8;����[�hQI�n6�PcQ�$uR����fi�o���]�*�Q�Օ���$�!�e��]M�km6���R�St��+IY(�����mI�V<i����剷A�q�W#M�R��bqE"l�IkPn�m�v�0��0��U�V�H�*��"�R'�aYk�Q��H���li4$'�4m�۩��$�%D�VZF�RR*�n�u�X�6�i����!9�YR�(�'q�S������ D2�	D��F�X���	ds�clUҺ�1�EJ��UUdj=�[�گmI*�2�F�ث"�*
�VI
ۗ#M��n5Èm.8�D ��]��5��JRƥB�AD�AB:(�;#M�\j���8&D��4D5K*)S���{D�%S6���7Ts!X�j�U�*�+,b#r�ؚqH��@��T%Li�+EeCr��b�K"-,����H��+b�,j8�UUu"H�si���S��-H���\�v4��YR�&���$�k[�ijDk�ٺ�k��rQѨ�CM�Qjq�O��^���'!��bv1d+R*�u���jES��!#U�\��Kev[`���hh���n�G"�c+���m�6$��kV��˺֧��W�{�(��wwk��<{����yEU���_��������{�*������>�ǽ�{���U[�����T��U�o[m��V��뎶�ӄ?����B5��G\��2WD������*UX�����V�A�UD�*���ux�C�i��V&6Z�ꊎWbj(�B*J1�r9&Q���h�D�8�9c��l�*n�j�R��J"��21
�e����$R���x�b�,�V��DB�B�0VTQb��K(�+#�������RB���TtE.�YX�X�#J��c#�9r"!e,b�!4�q(эTG��T�'$��6���l�A�Ri6�$���I�9*dD�֢���q�9�����W��i�e����i;F���-k���Wh��F
�S�����l��9br1��QG<�IL�C���������o��g.؃�u������
��{|Fp|���7N�C���3S�yݪs����%l sѩ�_w�/b�;n��5F2F�V�+T�HR�>]6������Ur�HF�%,��kr�6�홿���:~��M��ɡ�K��H�nF�CL;�������uN]kq��gh��h�5�ۭ���Ē�p?�������㧄âx��t:t�4i$�UbI%���a�)��n�s�r?#׈]�â��Ƀ�M��I�!�����g'�1�AI	M�g���&�'j	�B�,��H*N��Ѩ8h���;0�7���L��L�qIN8ۍ���:�:ۮ٢˯��$���$����"cI�����߅�8f�ݽ���:e��l.G�n6C�����B`�H�3�s�Q�s8Vٺ�+^�v��8d�3���q�bq�"іñ��I�#r�GN�Ĝp<��I#�p��v`ij�p�+���a�����z뎸뎶�F��ԏ,Q�#K$�I%�r��Gy�p�G��d�J9#�.�1�+��I�ѱ�v�\o�-U�M���^�4�L�E�l�2��\:U�b��9$B�L�JQ��ȯ�pӧ���i�i�+U�f�m�x�޴�]"tN��::C�'ڝ+W����8���^j�h�)3��n�B׮]��Z5�q�7:��7bt�V��JkrjI%�}Q��n��w7����z}���9柷���|k�|{o�yiN�s��%ҳ�g���ίw����o�5(I�w�w���y�9I9f�J��+����4�p��I��t4J5��;;t�􎃔�m�N�v��Sv���còR[���I4�Q� �g�x��3���s�c�69i�GN��NZ36BL��i�V���뎸�n�q�m�'j�X������v���Ε�}׽p�������ۻ�RI,��|L�vWUE��͆&�pl�EƝ����\r�����bY0�K���J����v�.LO�3�A��
$,K��0��G%3�v�(���`0�4��Zf��N��]q�q��px���!3��ˤ�$�X��rh�B�P���r�gLTK�p�I��S&���	N2< ������47;�O���1O����y�H��.R�g�t6:d�w#gy$d�ݸ.ع�d���61���QvFBJi�gf�W1R�:�J�5���n����[���n�q�m�,�DI�$HʼV_�\!��3��q�z����4̰mãm�Hu����	�ᢜ ��t������w��)$��3M�WD��l�i�4]>��s=�5~1Z���H��F�f�z�^���u�[uÎ#oYg5�na�.f^�5����4ՑN}�k9;Έ҈�(
�U�u5WP�>(�l��	Ҹ�JY�}ԒI��_~����������<����rRv󸧄"�k�np���7�*�o_gy�H�A]o��O_�<��{�rOWW>l>>�~uUSf��[j	uҰt��%p��3]0l���E�<V@>�tށ�)�L�U9��X�IZs��s�X�.����nvK�G!��GN�(�R�BG-�ej���Eu�dJN+
ҽ��zۋu�޶�:㭺��ӄ�I$��<˞1��C��L>..��=�Λ�BF�ŝ*[�MJ�m�0�I������w.��0�$����T�6�t�cØ,G��z�D��-�c�cM�E�>3Ｄd �p9av�d�0��tq���jq�*�$D�co��YE�0Zm8��Éi]J�󬭦Yr�u���Z�u:��[�[Gkx����b�Žb�i����->q��|����|�KKK����u�O	�6|x��9'��8J�0K�ÂRO�X�;�1ձim�i�[�[�0�KK[[���K^$�Z\�L9rc�,ǉh�-�o��4�4�L��`�\e�ZT[�I$�DZD\�al��Z-*���z�Ҷ�oXa<M/i+	Ә�b�b���^gͧ�հ��Kb-�Ke�^%��ش��%��in��1'�c�x���E�TZE�z�Դ�VE�K��h�+	h��-�+Kb�%����+���y~�q��3[������f�t�ӌ��x6����9�LPؒ�/��.������?�-���r����lI�39��/	��[��_/���x�ʬ�+����n�����vS��O>]�{ڵ�ޞ�����������|�Oz��w}����Zֻ�ڗr�����w.��ֵ����6���m�ַq��p�N��f�	��ą�ޱj��%�^��ȄA��;��`�4GqftFq޸�#<ke�8�����	�"ѐ�`r@�$aD�������I��L�,���a�h����J,6 ��(�P�уuIV \�J�(�W�)��Hr��,7%l�`�A�'�Ű�d�����I0�GLF,�L �/���60t`�.<�f���J�1Ȋ���'�m�]|��͸ۏ\x<"C��9�����y�/���	:���Q��*P�� u܌��S�B�e��/٤܊,&3b���$S8c: 87&�ƄICw�o�6�v�9���o��=�Y7�>P¢�C���iPߺ��eF������ù�����dXܿ�oZV���wg�x��ܳ�bS��(\,A�Ґ4���
�MaŁ��7 B�SJ��*�̯[q�|�k?��8'C�$:hᲜ'!?/[�豟��vE�M�a����M�E�_
F�yX��α��g�I�;Ub���qyx޵vs���!���4�fT�~�o2���>;��!�}��,�G��.QN�:��4i8�( ��1�V��;��'�z��㗄����>��.����4kid�%�P	
t���;�(�"�C�4�yR�"�b��e�Q۲�S0h���������G��:�sgz�4=�n!�Ɔ����%x�t1c�����|3E�g���������:�\���䈘������)D���j	gw�Vۘ��cSN$a��w��h�v�|��v9ٶU���D1�$�l:�8���-g,#�:�'��'��C�޽|�ׯ�>q�m�������s�ܓ�D��S��/i�2���@D(���S�yGsSo�Uۦ���=��k�8p��Y�4�t��;���;�sNd�-6�l�qô7P؎F NH�l@����1�v���-$�&�&H����3�	��K���	��Fe�Y枫]��e��R��H��H+�ll$ Q$0Z`gġr�����Np���ϟU�t;��M�;i�Zw�*�T+h�q�]|��>|㮺�ӁÇ�p�fd��Kpd����q��֧ǫ�toS�Y�>��4�۴w��G��s,�姄S���N#�ռ���������t����Y��u��M�y7��KNO�8��u�j��f�����d���Jߥ[��C ��� �E��� w�x|{�)��)��j��sIg����)�W1�א���n�η�����EHǥ��%�4�0li�#��r���bו��5*�C�%s^���d�#RE�i�d�
b�4��AD�Tl�h6�"�`TR�w�ɓGO�d���l���ǃǏ�:R���?�}���w��kt]_�s�}����d����r_2�_5�G7���ڪ��WHQ��D3Id1S�xk6��7����Lv�I�����s�)aB�k��
��3�j۷"�[)�	H�$�� >�v&a����� �r�18�p웴o����魽<�>]lb-<,�t0�ł��"�g�m�,(,x�qR���U�S�,e���Ɣ:�^d8�n��e����C[�ov����Q��=d|i�Gz|�oH�X��ZUa�ECuf+m���z��8뮶�[6�Kk�_$1��C������y�gA^Eר�����z�ITi%-�����m��c<��Vw�Ʉ��1���v���J�4����|n|5�t���;<��׆����Ea��7y��=��6w��}q�+�w��w���{}ا����!.�m�L����?���@茂(C� :z�h��!��o�Dv�^IF� l�8b,��Hi����6"{{%e�0 �Xi2¾7�$�b�Vg%vʕW(� Q�3���^~�^ �j�)�A��Mq�ԣ�9��;�w���G����o���noɌ�:V���S�gDt��ӤLŬ���C*��Y�d�� :j�d(v��;{8����r#�X�����f���
��[jӌ��Ϟ�u��n�qŰ�m4ν�<���J������HI0�T�h�$��UUEC%\ho@�%�K.F�2e�kp�2K;.��� ��F鯊if`ix��5 %B�U�֞4�1b8b�q��F!ƊxEͪ���� �K�!�) s������ˊ�����)����Mǥ�'�C��ԅ�`u�x%��C1a�c��?e�XP����u^V+j���q�=qo�u�[><<#��7���&Hv4��m���t Nͤ�W�*T�~�����P���W�VG�:�>-C�W�jF�����3q����4A<`��.�,όA���ߔݻ���s��2��q��a�Zu�x*�+�41.��G%��y#UM��$�l9Lפ��BK�%� a�G��p�NT�D9PB�ƽ�}�T=j��1�$�y��Dk�ɠ�B@����Vf{�}n�Ɖ&|i�G��i�^䤨ʏ�4��έ�-�]u�N��̙��sfp����l�)��3R�z� `�bтX��)6�	笠X�<�b��5{��<�c��d>�'У�B��F�G�&`�A,�L�b�eP8���`�qb����q���h�ϖ4@���ƫEm�"I=ʏQ�v���80���X �0�$[�,_��-����0Am��<լ�X�(��fJj�9c���6m��x�����a�~	Ԯ?���an�i��Zu--'Rӫbӫc���ilD���Vͥ�b��h��[la"ش�ZVVť�11ih�ش�N��SձV��kg�0�x��&	�0~"Y<HxOř<c��<N>ckc�oX�,��-2�--��-:����ql=[%��2b��,~2%�	�,��,�0"��ĺU^Է�'�����o��i��M��m�*��x�KF��Wq-�Kb׉lqn�i���fa�H�����-�OVť��-:���m��lz�)i�WRK�"�&���%�KH��a-*�H���-��x��>�|܉��u&;�y�gF�pۧ���!r�m�f'��"h/;ͻPq:�_��̍���5^u=*���ϑ���5�>�Վ�������)��=��QMLo�ƅ��%���`��/}:��!T<��S��7�21p��~F�v3�7��*)���JN���6�o�s�g����I�d�k�Gv�u�h���g6�"/⼋n��a��L5n�y��v��ϼ�����&5�����9؏uBa�ݞ�u���gկc$�kRH�A�$J�蘛Ʋ�	$��A���5-mH����Y$��7ak�ӳ�=TuJ�b���F:����VH�X�JE�U:M>��_&s�OӨ��c~��o������ֵ���U�������_{.�~����z��{��*�.���w��{����,U�]����Ő�8p���q�]m�8������3$����IJ<��A����,��!�t�*�bN�6����I�܉�"�{�F�k$��#��X�G+��L��
<#��+(P��<� �)
TU����6Q�!6��%���� U(ʥK�x�r�#$b�DXEr1��%�.LB@�.H"�*�GEr�d��eM�RP��1���A	AFBeC���EG��,JX���`�v.�4ԒR26	8�(�vѺ�Wj��V
�[S��)X����Q2��յ;�(Ablk!	���N�ESO�6�u��X�y$��T�Z�1Y\)ѯ6�lR���cq�y��əV��7�sO�����С�;{���E!Ž����r�������W���;;��y͞��w����f����Ԯy���}�>܂�-�z������,�~2g
��bu)��Sbȍ�)Q��P�&6�,=���&�!Lr@��+̅48�~�BB�����K�����!"��S�%�;�Î�)��کq<6i!�h8�N��0:�.j�#��+ eՄ<S°!{�zy�x܆�|��1��Ư3������e,>06���C�Ƈ���%ƛ6z@�z���o�[��[���F�l���Gs$<�������ˉj�UU+�F'����$><]M�D\��#�g,�Ǥ�����FpA��ʹ�e��1��-3:#�Y7�M�N��C�tY��#�E+A�VsbUfW��Z�G�͔��j60�F�WqІ�7_�zS���f�<@ff���� �] ����*��
��qP�U4��գǕO�,�S��V�­R�J��z�ź��|��u�\8�6��jq���c9sUUR�X���^!MJ�{�w����(3�2�d-���4`�����]�%���Һ�7rx�������(Lp�!1̔�R6Rf��7C�<O��d����:L����D#Ƅ�w���)���fhU��w\����s�gbY�CT0l<nd��"���˷L�9����!
C#k���0<��ݻ��p��$���M���۶$��:I8�{���L	h2��RaX�ǭ>[�[Z�:�]mӁÄ6|l��Ѥ�a�ʪ������.Y���5Fq� Rr���i��?(>
G�T����)"��!��CNͧc���&�Hp�J��$����ʺz!���ur��1-���L�Dd9�C��d��YCH�T=;$��e\Wնñ���]ɑ��kna+.��Dht%Í4@���%�d�%��̓'��F�ٱAe��!��W&U�[O�uŭ�>un�ۮxGO�J[�3ʊX�䜕�G�E���d1�H���2fHG�̺�r���$D���޻=��m��C�1u��z���k�oO�����iQw��Ǻi���!��]�G4��gR�]8OOS˽qw�}�/w����G9��>�~'����脆���|kak�āAcb��u���&�Xt@�E�e��:#C,E�2��zˑ�d���7#T�]�a�aq0�8%l��0��7�^�T.S�cd�<`n��NH`u��g��-Ƣ�b�f�IC������f�E��B�7������G�1G���ʸ�b��d�����[����<\�ӆ��>uku�\8�6��{����wY����Ν��q��^�WӔ���]��M���Ͻ}��/y��ģ\�֊G�m��lɲ�������k��g�w7�ֳ�3J���:g6v���'c��������U�?s�I�}�����y�$��w�"R��K�'�UT�}[��RU�}H��"�ג�5p�d,�,�=~r�X���]o�[u��C���Pa��Lh`��(/��g�f�Ι�̚c���P�<B2��?�LΈ'�/|	�E�����Btnp�^��B�q�ӊ�2\00N�����Ɂ�� d tl�շ$%�l�C��e��QQ^�]V�Ȭ=F�2����V�խm�����������MNc:�ݪ�� �	%v�ԽRY��z�tl6rP`�h�e�d.</��.@��hzpp�::����"�5�\��Ɂ�C�@��h����f�V��ZTu�47ie������8d*�$�W����`�S�������ǸB�2  ���w9�y�8!foS8և�x�����dHe�'�1e�v<caÒ�M�>z��]|�ֶ��������`�G���*��@9�M���.���z���d�Qu����ɲ��|c�kA�Y��m��u��KD�����nh]�hp��ѱ��Ȅ&���F��h}�����X���A�2p�Y�e�HX6!Aq�N�.�A��\��G<f:��c��a�	P��# 4y���3�|r�Wk�e��m��]m�_:�������:p����j*�/�B"��<�>0��ْ�1)��g�8��Ѝo!1�-�'dWl��6�m���w�Lo��&o&���	����Fy�0�40ð�a]��<!����T�٭T��w|�o,s��M�]�]��{�M�f�V����3�Ř0�X�g9��WZ5WV���W��)��2`���<m�������*Ҍ/""�ܰkH���?��L�/رb�gCmZ��nW�Ր�u�6;I^IR<�+a��J�1�����$�Fs��߼{�\�\�@�H�'5j?�:g��-�/�]�+/�u�Ž|ۮ�խm�Î#oYg��&+rg0́�b�����]*�?׎�T��W^f�!|�sO�:�1��kY��9]-Q�)Okv�c�$�����f�7�[̧V3��gLX�D6g��e��ڄ�NM�lC�=EsϦl�Y�Ř���^>+Gٮ��2:�q�y�-�C!�\ I��\���y2�\����S��5Z�I�Ѥ�KN�q�#��-��H���E�V�Qi�aձiպ�i���kc+b�ޱiiiiԽ�--0��KxŢ�Դ�[�u.Iհ�Դ�G�aox�OĶ�#	ix��4����[�L�u-�K-�E�V�����3�|��'���+��>4'�A���G[Kg-2�l��-:�[)$���*�L%��iV�m��6�J���S�Xz������u����|��[����%�g	i�f׉��h�z�--�KĝKKu��0�-=F�)u%�d\�"�"ȴ��-���F��Zi*�<�ោh�/{���~S�������޴���ֽ�~���-��j����N�]6{~��zxE��w{���b�:���Y�/F=���cߵ�P�浛/�4a��i�\{X�S�*��N����s�	�n���~�W�:����+J��]߽�{ΕW�o�w~���:U\V��e������UqZV��w�{�C�p�g<x�����Ä6h�I�X�*��ʄ�P�
�㚢K2:4�̘�
ap������Aɡѓ�Xd�5���&�紅�1f
�_�u�[�֊b�����P�j�y!n��=V��{�{�x�Xp�|#LA2A��k�ct��-|6*e<p1C��'���>��t��#�>u�筺��V���8��,ߗW~�r�UUH�<x��z��x�^,��U�L�;��C�4�X�K��U�덽YϹ��n��/U<g�{Z�Z�_q[#e�g�U�ɏL����*B?Q�J&�Ox��H@�q���$&]Th��{Vޫ�k���̰ۮ:��n:�խm�Î#oYosŽ��ī���G]cۻ�5���l�ʢ��'!��&�|}��>�}͕	'�����8�NpK�H�}>�UT��Cz��G��9ػJi�8S��B�y�?�խ%`��ޠ�i�<��ݾ�ؒ����vNq�6f�[�*�o�0�����+ǧ��,6��%��&�!`�"B�4K4��ESիHQ�ۣOz٢��2�+-*+&����SO+:�U�q�,�Dc��d���vX�Pxx>��/tGe��h�cG���n�n-k[�t���Y���m������������o*�����л����.X/��L�U�L։E�(ȇ��or{�l�v�D��@�=A���f�>������S�Q� ;��Fÿ���Z:�]3��L������0X66(��n�,66i��iX�Q<V[a�V��[uո��:xA0�{�W��E�ѭ�ڪUT�*�P Hx1W]�e��Zt1��W27G���!q�\���\� �՜�J�U�=^���"��b�;-��&i���\�h�4r��2�}�|�1�I}��O;�e�׆j��m9$i]4�o|I���n�����o�Y�33I	o����"FZ-�����[źۮ��Ǐ:xA0щw';����y;��*�og-��v]��.�9�7�i	_c#���u�1���UU %]h�`�k?E��Z4B��=�1XD9ϩ�l��ܸK��e5�)����d���o�/�t��1�5nj͇[��|�h�UXh{okH���a��Z�iO�z�+���zmQ)�;Yq���<u��q�έk[�t���SX��1*��R�e77��P;��n�758��Mj�Ϳ�I3�޶��#m+Ti����9ߕUT���ts�;��gN�.�9�f�}?M/t9Z���k�����7�+�!�5��l����O{ǋ���>�����m��٧��W��Q(_߯���#9��Q�|W
�I_����j�Q1�m�=a��
8i��ن�q���D%w]#�������Ⱥ2B\�*�E5RN�BIs�c������Ϗ��ĸe<!?�YR,2f�gL��ƍ��߉<0vz�6�dhy��VO�4C����&ym�Uc߮I���jo6�$�
�AH1j�{\��SW����]u�[u�έk[�t���Z�x��Ĭbg�U��M��	tY����Ȑ��J��j��x���&11���o��R=D|B^�O/c$-C��=�`����oX�w>�w�ٯ}��9��*��b�����g��2]F�Y�����YX�W�Z*ΗbBz�Y��Mh�&�V͑ WJ�LrcC���!��5ǯ���L�a�^�㍸���V��t�,����UU���w�I���n|f�^�t�gNfh���i2e����.B>�S.}����:~ҝ�}�8h�����2�eY�J�M3^���&�F��:�&�(���,lt=(l\��g#�^8��㮑d��f��x��BB�r�68v]s�����8��m��m�����Z�p���V�fI���\,��I�HHX���J�d�y���lp`����؏ĕ�DF}[��p%`HBJ7��Qq��!�C��\z�N��ş0�0^T���Y]̙������������k��8h����u�9yͺ9�~3�Hb1��-��� [�d���Q����m��!$8se�x�I�t�p���:�u���.�i�Zulu��KKu�q�z�O��شf����K[�OR�"�l1ii�����-�u�R�ձ�z�Od�[���-�+	il-�M-�KE��-��:��-�Ę���$����&-.N�h�ط�d�<[�O�+{�4����[8�������-�L&$���*�GϘ�|���m:��q>C�<CB&Hd����c�!��<_�>/����N1����^e�o���י�z�V�In��i�d�=J�e,�"Ⱥ�U�E�i�'RҰ��.M1rx����x���w�����9�zNw�s���y��_�������zz3ݾYű��Ȫ�שlS�f�y��9K��%��K/�;��`�M�����N��x������َ��zή��gQ�|�n�!�l篸"����n������W:*���p��iF��L��ð�S��VOq��f����7M��E妚iH}�u�|��9�6y�s�ۏl��T�{G�>�7}S�t-f���^$�9�F�3F%)-m]��������PM5�,�#��,e�J��M�Lh�W�$ �ZuԭC�7��%�Rl��EkU�T��v�|��ʸֵ�үz���ޛy��n�w~���yګjҷ~��{����U�]-߲�����;UmWKw����p��8p����ֵ������Vf�1��*Vs�JG[��1�����j�X�P���eyvd+#�������&�%�q:1:��J��ę)A7(D�0���Ҏb7
��x'��$F:I��	
D�)K���l�EH�TF;!mc#!FRя2���n���e�S���pM��1��[�$T�B���4�Y2��L�XǗ-�HH$d&�%��"C��+d�P17E$c�c�Z�I���T7q9#Y[�te��F��D�ԜnI�eT���&&�&�����d��lkm�myh�V�'h�eJ����Kc"��˥��L[B�H)����U�QT���7����7N�������_q�=���bj�x�Û>��~������ߏRU���sZ9�~:R<t�<�B#W9��sM=�v�4�st�oC�\ҩy�P��������B��4�t���3M"1�U�]y�Z�a���T7�BxIi(�����z�`�(�"��ʮSH1|_"~LoOp��!d�g�3J!�x�<c�R��I��x�����C2�'%ID�q��8�]m�V����ÁÄ6d��\٢�j��$0�֞������£H"�Z|h�V�U�B�*"2+|ѢgIL8����5���}��4�"<q��/�P�y�J�X�Yzj�_6����#�ב!��8g�џ�pY��!����^^��l������r%.7.y�[24BÒ<���ѳ�q�n6��έn-�8��f����1ɽ�tn˄��-��޺���Cgd�HMn�����X��[��-g��u��t����ω�!b�������ک^ؗ�א|(��%v�4��J�B�T�ś/���hM]�W6;s�e�h��ޝ+�j��|�y�iUh������?uiV`�U��84T0�b���[o�|ۯ�:���!�%��x��H�1�UV�W}$�M��ô�U��8�Z��9^����^=6n�����{4�I)�Ź#�$��J"���?��r7<0��D���t6ptn82B7ex��VB�)� пX�f7�ɐr�b��!$�q�°n�_�LT�kN+�e&K�+Ƽ�F���$���u���E�s���Ŷ��uk[�8q�l�fk�BFQ�3V����2B���8��A�,��f��)���Wk��6��m��1�k��?�_������v^N��N��1{_���c�>2@��e)�Å�(F���h��Gt�'g{�+��ުk��m�����*�K�!g��� ������ 䏺G�B���Q��.e��M!����D�$���`F�̠����6��Ι��c*��*����a�B��vb�i�[!m'�=�!
�'GfL�W+L�h�n�)�L��DgU�xt�M7]�_���xۢ�n5Y�s�+!��x�*	꘬�F���^7�>|�m�m�ϝZ��qz��j�_v󞕙�d�4:�޿9�/���y�?u�N׮������s�����6�m�d2;�m���dс��4Q5*|��"���I0j�=	9_h�l�CNm�e·���Cc��$����X��{4B��>3DC��=?bk8g�wrB�֢Yc���-!bFI-j,_G�|6:y�$,:#g�:fHt/��(�׳��y�z0{�@�,�0C��>l:pb��:x��ζ��:���8�6������%L����p�:�r�z⪫I�u��Y�c� �i�n��~��\��%�K_��D<�:�q���~�����}q"��)Ӻe:B�6��*$��>�CGH�#1�q�������f�T��VHC��	"�%J��MӓuW{�f�[6��W��o]m����n-�|t�ÁÄ6h��u�j��$3�*ʳ��!�[~�"Vρ):C���3�)�3������F��/���&�me�BQ��m_���?��0c1���G�����k{zgL��E�1$!$��W�!�@�(r��i��bG:�:!ر!&SR�N�B3��fO�(����
Cp9"�G��/L�sٟ�n�Y���[���m��n�n��F�!���#��^�鷣�i�{CM��a�s���3N�6�\9י�5a;���,���L�)DC���~m��$&%��̙���=��7�<ӘpM�̷�ٙ�Zo}�뿠�7�8QD��f���t����r������ӿ
M]�:ʋ�c����_^5���cg�����b�{�P��W]�1���j4K�bˌ�2D|gO¼���+-#*����� �zH�r��^��P�^+�j�2�n�T��-����G*!�}\T�U��i@,3�SJc�I���ݻ[w����thV�nݫ�ǃ��#�\f.��?jc�r��u�޶믝Z�m�!�6h�5H�W�^s�*����q5cÖ���FBW�����?��2, � �G���}ҽ���`d����e��/�%Uexbf���m��ۭ��/Rx|v��)V��Ӎvv�����M���M�!��Gό���Q��u�xi_+�Q�SL�*iZ�]kV��N�u��mn:�:tN��tDâ'D�� ��"pЂ$4"l�:lE����BlM�D ��8"pЛ �Dق&��c%��6&�ن�,�4%Q>HC�� �"P��8�n�ۯ��[H���Z���ǎ<��0D�"'M�,K4P� � �%�BlM��?/s3��%�_3ۺ��=�/%^���j�y�5�O/C�3���MvoKӾ�������.�u����{����NvS��+w��V]�v���r����۾u���"Wcr����Z�y��O���_{��8M����9������f�<��q%��`�>��v����������Z ?MϞN�|�O/&�\ۜ����Y{�W�����9�{׽��+������������͜P�ʏo�}�PW��w����W���v�y��J5��޴w3[�U����Ƹ�m|]�q�pi�xA~�-��M;ƼV(�%�J�"�'ݟV���k�v��������	���=��p\���}��Oo������l�Y߷�������j�[�~M���Z��F�H�?~��O")}��?�Ĺ'�9�|D��%ʕ�Ev|������i^֗kQ�^>�|��Y�d>s���U�{��o}����3䘮ֺ��keeiֈ+y|y����^�9�ܝ��y|{�w����L��	(x]�-̹ե�ݞ�g��/�U��a�'�g��u�������Ћأ".�H�uY����[����\}]�f�O(-CR�*� �3~����S������\�=w��{���������U��߮��{����ڮ���w�{���ڮ�t�w�{�����v��������o^�m���kuku�qf�?V$�g;UUi!���Ķ�V�>i آ$O����>Gà�Ft7�!�K��ơN�Cկ����KN��y�v���ٗ�<4pp`��cR$���E�v�ؤ�K6(�F�r�f���d	 �\��BC#r��S#�⾮y+:I��ã枾|����n���<xG�t���D-l��ZW�UV���5��J���i���ٴ�h��=:N��澼����u"{�ξi�j���y����\i�a��"<�&��&��"Kq[vI�$!���eT���d6�ѲQ�DX�G�g'6��!̶,�m-n-��]u�[�\q�q��!�	�bMV1FTDeYm��sH.�[�,b(�q����jӉH�īm�N8UZ�U"�UU���5z�m����~90[�F{�я��<�o�=�v���:�l��7��0��Fx��΍s�%N슕p]�5o~ϓJN�^"W�T#�2FK}��E���`�3���|i�W!�O8B�8<8l�����-I��h�����F��v�kd!4hZ5��N#ecAP��'+�����I�|�}$��l~4��~�Bƚ�Z�H�.#;�kq��^׺pc�-dz�uӇ�4��[�V�^����e�2�Og!p�Lc�f1�UV�l��d���ʸ�,�+LS��ODqW�#OiLx2�U��g�U��8m��h�8\���5D�ѯ7��� ��5K[H�����6p�S���6�%]g+TG+���a��-BGT١��C����a�$9�$�w�>��i�[[�\[�uku��8C�y/�$�s�hЖi���2B2	�=��yϕUZH(��I7�c�OLg�,�!�G��m�2ʛ�4ǜA�g��<CD5����.`��a��#D�,��P�Q
��,�RZ�|WRpۆ�!
���ܑ�� �h3U^,���v�IQ[:]YMY�|J1Yb�V���_-��]|�<%�:t�J8a�h���r��n�����fHȚ�yk�s�l��{ǖ����ޥ��o'&���4o_*������:�s�T���^6\���A�0�ۼ!x�~0k8,̼�|O2�bJ�>�b���D7�BB�0BeZ$æ!�>
p����Q�Qi	)4W�Z"B����#�q߇��F�!��-˴_m����Meˑ�Q��i.B8���=mŽq�V���\qa����V}�m:�B4�d&��V�J*�+�HҶę-�d��?�m��1��ݟ�9y˨^9�G͟��]Ӟ枟��;����'����������C�>����~8+
O��4�W��^��U_�;���&��=C�	���N��Yg���u�(��d!��z�	X44\��zu��!G5Ag��)�}z�3�{��đ\e�$���Wk��e���	�eu�����Z2A����ioXF�I4i_u�Q��7S�����,B���1�����衔�3�E��&g��m���t�eպ�k|�V�\x���e���=_o:SZ/��cY[5�*��D(M�|��-�H�te�᥄���?NF��Hf���!gGd.p�x�`�Ĩ'cQ�]��Q°V+@`���ɨ�)��#4wQn�2��ʶ�Ʃ���b�#�Dn���k��*4���>z�]>:||tᓇpM�,~�ŉ�$Y�&pg3�d0g;UUi ��IQ�(���K���ې�lp<\!��C%�\��*v�ָ�Tp��9��ʡ�A���d��mGf�Ŝ���X��ꖊO�(�}u�$��������+�$�V����IS�8<�C��ĺ(�$s񌻆ö���pl=���x�r:x�޺�պ����Gm�,�0��Q*��$>+]C�X+U+�I`��L�4{G��J3;���0K���C�'hl;X`���l
)dv:�N�0(�cq�&Ŝ��Otp>�Q���vj�gzm��HMޖ�:6tf��m�Ͷ�km�ۮ�뎶��: ��8'(D�"lD��%�D�&�M���D�b&�Лf��d����'"CD�b&���%��6&�١8l�6%Q>C
 � �"P�6?p��6pش���:qŭ��n��q��x��6x�"tD���XK� � �"%"lЖX�"x�Qˬ��~�5���3EL/w�G/��8���n��WT�H�I�����*�)Y[Hc�bŹ糯e��<�n/s|��ž��S|���������l>��W�J7&!kfw���L���]!���(�K>vcB�d8ij����7�������,�U�e5\K��K%�����(EkI��*[q���l���s��K�^W"���.����uoW��E��%�ONs�9ƕ���������Ƿ����v�70�j�_)�qsbIkU�J�Ե)��v�ڱ
4uˣJ)�$I�eX���VQJ��kV�4؛�&�+bjv��!#`�������V�Ǯ�]�w��{����Uګ�����{����ҫ�����{����ҫ���~��g,��x���x�4��ӄ?�#�^(�����qK-v��%(��$�Xө���n�5K�R��T�����!`��UMN�H�4�B���AI-�Y$uBY�Kh�Y��*�,V�܈�X� ���St�P�L�@�rex4J�rDG[m
9�X��c	�Cs�Ԃ=�D�*�!
�+dC�B�,�S
$��d6bA�)��$�*8$�[)V$ǅ%�7t��&h���h����W)IHZ�K(����֛��RR��Q
R��H�⨲H�	j���C����ʺ�w��#d�Im�*�������5�IF�EmF�$�bYb�飪������Y0k#MVU ۮ�"���YcV5S�',(ܗ)#��Ͷ�n����^�$s�kU������޽ �A���n��o����;�"��މ2);����oO��ޘ�%G��ƪS���f�O�e��3�DĕD�����0���X��:;63a�Ab��Zϼ��5�\{co�9||�2J�>2Vʰ�%���+�+�����[%J�JK���V˗�L�(�EF���`8� �p,�4՘=fH��d�%|h�㇎ܜ:p������4Y��$*��%Z=��ۄ4��N��.J(!�T�R�����h�Nۧ�go�>4���_�Y�t>:�h��\ӓH�.PY�Q���_��<�8~jR���`���ł�����!,�p{0����x��e��d��)���2tѵ��ַ[i��z˸�X�Dc�ƕUZ?I�2Yb���7c�d��m�E�s d(�M�iᐧO�=�-����oL6i���z��/>���j�,�I�M6�3�ÿ�>(C~��l�gmՙq=�c���
w*|V�8��}�n��<��)^�����4`.B�wG!	`�r�h��I���+��u뮴�[q�θ���.8�0�־�R��Yg�9��⪫Bx�چ̕�TU�d�.��B�,�ع��ٜ��ZB-D�|����$��s��2׳����ɪ�ܾ_�{_x�h�\Ҳd����g�F���S&�C<g�Ѕ=�g�F@ɱ�*29i���nH��ij�|W[|�_6��u�x���!�6h�o��.-[��u�!���9�G��t4�[h���"D˜6�m��O��'c4_��%�N���k�+-f��s������[���ruGӇ��<|G�ļ'�9 ��<�:k8��v��Z/z�j��ϯ��x�����݃�߲|��vCBC��?gxg��hh�<�x�ޗ��L�ˣ���Y�S����<������1

F6�hf^g����6'��[���~�:���Y�j_o[ܻ�/rNΔ�1���S�O��/����ޝٝ��&�����/ik���Wu�a�|�x|�Yֱ��������ku�O���,��f����V^��^03�^m�z���ebs��sx���u�mȋ�]���w>UUhO���VRR���j�+�`����d����,xw�-�19z�0yu$(���@�w�<dˋ?��6�r5�=��J4R����KϏ�����@�%w����J�c#k;nG�N�|�u�Z�m�Glт��v+�UV�J���2�dYGܓ`�����jI�erU<<���f�?Y���{\6*}���
�<�B2a���j��i[Vڣ�/�<<9�ƍ=���1y��)����ˬ%IR�;a���M<=#�Ul�q�����뎭n�ˎ#�4sz�/-��%$�����НO�2�1�����
2���vi&�̷&/�Q#8W�h��&C�z)�B���� X��m��S��j�/<$�su¼V�!cdOZŻ�+�g��A���(|{!劙OqBJ;�p:���g��8�.l��_8��\uku�\qa���&&~�&��(�rQB�(�!d5tt{k#r�&6;b��y��m�ʷ�:}<��t��ry���4׿_���F�̻��d��g+��Q�_t�/��E��>7�M$��4����e�$s�>J���e�Ϲ����}�:{_�����*���}~Oc}��CMۦ�_�����F�4h:�ٶ÷D�8Ք���ueՊ��V�Yx��C}�JMސ�Ň�a���B��:h�_s��c�HW�CG����ҭ�R�m��?m	��Ʉd!!�k�����
=O
n�c�h�/�u�u�_-��q�pΜ?h
�om�[��m��;����p�ǅdO���E�� p�v9��0|��̰]2�}�!�;�zp�7���CѸPb2�l��������e�tDp���	$��,�G0q���l�m�I�h6І��N������3���FN��6x��tDN��:'D舉ӂpᆄHlD؈����D�4"X��:lL�؛0١4A���'"A6 ��'D�&	blM��6hM	�F	�e��,(O�A(M��6�L��׍-��uZ�Z��:��uu֖����׏:aE�f�AA�L��,؜/[˱�t�������{_�u����<�_w�Z]h��ݳ���%>�&��w{�����D�{��*)��՟x�9�N��j��od���w��ְ溺*�D���$v�w�{[���^����9��U[���{����{خ�V������{����sޥU����������<ZU[�����g0���>:p����e�8C��h�f�����mRR,+1�7Ӓ��R.��0�9���:<N�+�!��[I_!wp,�P£*�:b�G_<s��]�S ���ٳf�̚�f���^�������+4�\�֖�孷�6�:�g�Hx�����D��FQE+ȗ'��Mj枪��o$�'׀��X��!w����\m���s5ÕJ�ݕQ�xz:C�ܘ��g���������t�(B`�j""�+�T�ߪ=VVBՂS
˫�D���}���VU��W����|�o][n����~>:CǄx}��G��R�(��`V�:����"q�+����\�3����w��9�l��tټ�7	yÙɤ4l� ӛ���d(��5%&������8S��L�y�c;�8�U�)�ٳu½���U�8�t}D�0�����J�Cq�h�w@��G����`Ԓ�k�F�v�쉦NEEx�j�䇇���+���!��dsclŒɾb���BI#�RWJ/�']z뺩Ҳz˭-��m�\uku�\qci���^�]着��`�2�U��Q]'�B2q���������á�w��9``.��=�!�f�P�Pp���A�~�=�!��0|����vH;�)�?�7������po��+ ��b`����vU��rt�t�iV�Ɯ[�]m�\uku�\q;&�[�g-ۥUV����we�F��"F+j�õ�q�Jr�_���:d��'td<hnom����}{�\8h�$��c�4<���s�dv��h8�M���W��N�rj$B�ȓ�}���V%�ҙLܧ�O����ͺ�ku�][����M�guw��Pg3�9l�1l�'qY"�o����w����-���_s�Gc���>��B���z���ĝ�i�Ֆ/++�Yz��%�z���w�����é6}����rV��C�Ƶ�w��������p��ԣ��˚j�}�JD��]?RQ�<�����ؘx>筚�����a�#��σ����g��~�_۔��'*׋X���<�pp:3�,g4G��P��j�aƝ|�_:ۮ��?��<>��<�i�~��WY���h���"�Xj���"e�����uآM�j��G����z��ч�m�I�s��I1������}��g�J��B��!9�<u��7Ǐ_^�u�����ê�}4�Ə}w~櫵�y<|fʓ����g�$BHL�0htL�x>��4�<n'ӽ�Y>�Z{��˒�@��VW6K|���Ex��(�����p�Pd��Ĥ5�\%Ak�Ϣ�H"�F�J���d_ȁ�	���_V��/�[km�\u��8�8vM�'$V8ڪ�CZ*��V������ϻ�{�O_Vx�����U2Q0�p5�U+��wF2ѣY���*W�R�����u�^=���
�[�/�1h��{�$�n��tᤅ9,�|`4���.��>F[i�;q�θ�-�q�q���p�e+�UV�j�Iʫ+�% �&9��jġ��Uc���a�t8�ˀ�:t�Yd�7|~UR|T��+�ݼ�}�u����x�I��^:���rM�C��$�
��HQ>�s>���O��'N��<tG���.�$��bBH�+8�UZ9P�]+���F�ɺ�Q��'}�i'���Ⱥ{��G7�kD�p�����Nnt��o�%��F��%�7u��d�p�s\�'d��$ppn�0�Ia�w�`�a�M��5^�r�ZVtiŸ�m6N�D���tN��:""t��,�(�&�DD�(A4%��	��`�b%�٢� ��Ȉ��0�H"&�D�6'D�0�6&��(M	BP�h�lM�(A(L6"`��,؛<Q�D�O<Y��'D ��m�Zֶޭ��x�,�ΝAD�4hDؚ��z�Ԕl��i��Ȟ���_z�dI	'�QT���Uj6<��Z��&$_�\;���vͪ�u7�E}�Q{��T�M�����_B�%G�Lߖ�".R�����i���?��O*�q�F��C�?iޟ0��6g�-61x~I��W��;ٛ�zrX���̜&�5���]\0�Qtx8�_8�1���t��Z�'w�����>K�?=��v	�-�Y��MJ�5�5�����;=~�4���&�71
�vj-Y��f݄L�pB�bl�̞�m����9�oޤw����`���Bmi�qTQ��&5n6P����J��wW�=�OL�����^^��U[�������{������wwo��{����U[�������{���*�������=z�����㮸�����z�3}�j�����Y��%"�&DB��$$��2�"�eM:WG+���$���*yP��a&��D�Ȣ�:Љ����E4��q�؄Ah2D����qD���8QU#%(�+tX��ҥV"\�̢$.A1�B�"����!��eYJH�H��%�p��A��
������,hUer�y�� ��E(�D�o�Q�e*(�Y2����,�$w&P��#ݘ��m�Zґ6崰S-jeJ(�Q֝�"RKnRIm��l��LMT+^��H� �eR�\%��Q���.;Gm�[I%X�RʣD��D���:"�V�3�c+Ԣi�P��(2\�dn�ڢW��Q�'To�p���UU��y��z�ӫ1w�yn�#��7�L��Y�8#M:��D�Q4}��C�����K�gW�g;��v��ϼ���v�J?!zjﾯ�Δ9�>���o8�=bB)���FgMB��Ia�������gB���a!�ǥ�!��C�t�!�Hh9}�l=�;���s��l�GN����hp�B;�"�!8�C�Zh���;����d��`U��Z���[u�uŶ�8�6Y�o�q��ID+elK�R|@���LV��l��D�&�&A;y����C!�F grFp��^�,��+mh3~~c����Q���mu�I�Sj�Lו"<x`�r��T�W��s�&���[�"'N��<p�N���F���E���3rI%u'j�la�EF�C+ޗ�$. ll�n�L�礐�$���ᦌ�
8I!T+ߎÐ��S���2k�ٴ,�d<7z���Ct�^��Gm��ídt�.�7�X.[0��͌xۏ��n�㮸�����{]�>�I��$$�>Md�$�Xt�C���jV���+ �1��˹k��!�a����]�.6��!CwY'<�43G�H���4�����V�	�xMouu��5G�ڕ��S/^<x�V�ku�]qm�Ǆx��&���4T�g�R��4K��S�U�ޞ�唶%��k�Z�m�m_�I,>g�'d\�s�9�oy��˛���w��W9�O�	�E�YS�ÆV���7�M�r�fN��_m��]����-W|��v?���p��sK�8bi�s�Ұ�t�I�T�K2���i�IOI.6c�4݁�kK`�I9�B1<$�ēl][�8v��n���p��Q����v�|6W���C��(��ɉo��pp�t�i�;�'��J#�\a�6�u�uŶ�8�6���IW��x�uv�Ӌ��_���v�[�t{ó�ډn����O����\���^��z�7l��$�ǃb�98g4����Ē�љ?V7�.���s�nrK�g��L^+��\�"K4��<|`�+�5t�$`ۯ{*�M�leq�"%��
p��A���w$!$�>=�&Gsm��G�Ӎ�m�qn6�:돛G!�e�&��I(�vƖ
�kV����z�a.�=iu�{��7X����L��=��Ev�9��?��7nQR�Y%
c2i�?2g埂�1㇃Ι�!q����Ͱ�_āM�@���b�4�m>,4WĆø��d��DFH�-����n�㮸�����z�~��MT_��F�Rb�$�IN**a���b��w�&{O?KR�T�P�!$����!�O��A�,���ABq���)��u����t0K���6�+{�J�N�
Ƈ�dKn�4T<R}��U���bL��
2��$�c(g��z�Wkn��j�{G>[O���o�q�\[h��l�LW��̴�s5�<P�U	n��TK�*��jV))+u�nG�9y�I%��Y��_>BÞ9N�{$;�pK�${�����"ь>������.��E��:x�����g�?��>�y,u�q�s�����խ��k��}�!�5�7v�'���[0Z�F�{Q�&�ʽf�����f��>ʒ!즁�ѾD��-n�Wdt�����Ð�A��Hpr:��B1�oPl���8��ϊ�N$�"Li`�"X��~K0f�g�1����e��덺뎺����:C�ħ`C�ӎ%�I%��;���(n���p��ĒH�6۩�H�J����e�����L1��S'h��Fo�&�7�ۚÝ�3�֒�V��Gm��$��+U��O��<h9�0x5tY^<q�J�{��z��y&�|��u�\t��tN���8'(DJ�؈��ӄD�&:"'�6&�٦O�AH""X���0�F�DnDG�'D��0�blM��6hM	D(�lBX����܉�t�.��t㈵�o���(A(DK8"tD�,O=[֌,��,��]G]e�YdM��,��_[�en���r[�J��.��U3����:{o���5���٭������6zo�u�#[Ǿ�ŭ��k�Z��>�I��.}~�;�_yx���(ͽ�<q{׬U[�������{����U���_{����{�b���ݯ�=�{����U[����fYf�:"q��8�6��y*JO=�I)�<�2�-i*���0;x�0l�e��P�kǅ2D�d�Ń��=6޲hٲ�$>|l\[���CW.�vBM�0�]9=��q�c��u�Y	/����	���p�g�$�GF����ފ�l���<|�o�q�\z��#����'�I%!�=q#�{4�@�R��4�ψ$�Qcl��}$&�.�ʧs�ӣ�s��ޝ�;����4?�|<g�L�x�J�hOX���n��`i��&��^ֵ̲��u�ͭ�;fٝI��u����No��o9�GP�t1��R�`�܆��r�í>i��u��:㮸�g#�HO���^���kǛ�)�T�d'Dv�>��v��N*��{�\K96�u�Z^8歺�\�vU�o�S��}������C�}�5�,%�6���m��9�8����6�!���{��r���3�����99����������M��эsy&�H̼-rLp��\ܛ~({<f�L�d2Ra�f�4�66�d	��I$��MΆ�؆{ѭ`cw���
�\>,�&�B�W�;�N��4�))<!�M��uj�%��z�S�sn�5e2��x��$�)+�ɧ����^��o�q�\z��#������,�f{���ƸMׇźvϖ�Z��]�1�L���J��K�S>�1����̆��B�(�'��HCI4|�d���):�WUj��<����75]Ym��f�<Rr�����5X���\��L��^V�Zu���[����ǎ�Ǆx���܄�?wwS�I$��ؒB��I2}���R�ΓR��L�
�&B�a�P?��|<�2��?�������'����Y+%�����%n����y�x��W�;TplBÐ�q���ctJ88og��
��Q��8p��m��y����-�i��n6�:�Vq�<t��~�w���]����K�ߞ��͝��\K���c}�:o�4~Υ��t�?$�F\����΄Ca�t���6�3�ȥ��=~i���=�ny2q��a�͛!!�F0=�K*�r���\�4�����{���m8S�"�������.b�S&�+,+a]a�޺��q��������8C��'VHЭ���|��/2m-X�' ���Jq�,��$t�4�����z�������_K��Ȭcuci$T�%G�K=�?z������y�����.��
����ר�Û�.f���v�.q�*�83�rxy���IU���L��ݜ�w�5ʝ.�>�.}տVu��k;�5ߋf��}R3��yO^s�j�JrY"��I�s�v�\t�ɾHB�rsRQ��!'6p�X+"g�I$�(���Ѹ9-�q�g���,?aM4���/ÿߚs��YP���CsNF��.x��La\�L�C����:�箺��q��|q�m�.V�-kfI$9t����Rlp�ht�V����=wl�i��������Q�Xi#���,f�ܽ�F���N�H�����"Er�'�L�b3�nR���\Fig�!����X���.i�/[|��[�:۫8�6��4�!��$S�$�S�IX��7!�f]=5��U����``ܡ�a�L�k'zW�MSXvw�ԗ�>��\%U�����k����Ս�vy�5��N�*d���h\bCs�፷�Ҷ��n��S�m���oV뼓���<:C�0�Q+��v��$����ǯv;��HI(z�4k�6zS��[�����L�M�f�?~������U�<�hhƛ]�)�೑�=<І��kg��\�cY,�ы4h��IT��·�L4�߂�i��S{n��t����6���~��iK+�j�R��6�q:~����������4~��]mbn�h���x 	�<����Y�*5�k:Q^�H2��>=t۽Mh�I4�h��I-2$�iE��ѭMdMF�ZM&�Ѧ�K$�h�mid�-DL�M�h��d�h�)dM2�"h�$�:��M$�"4ȉ"h��4I&��h�$�-�h�#M��"&����&���Ӝ8Iid�ZdK%��id�Y&�F�%��I-&�KKH�&�Z:덺ȚD�Y&�ZY2h�id���#M$���$�kH�-�$��I&��$��M,�4�M-"$����MMh��ɢKKKid�Ii���Ť��4�&�e��I--&I$��AĚD�D�I$�&M"M"M$�K"M"RI!$��&�I	$$�HKL�i$$��Y$�,�BI	%�KI2�d��$$�H�L��I$��I��ɒHI$���4ȓH�I!$��Gn	d�ZI%�K&Ih�M"BI	&Z-!$�Y$�Ѧ�&�&�Ih�H�H�K%�D�$�Ih�RI��4Ii$��h�&�ZIi"i%��i%�I4��d�"��ۉ4��$HI���I-,�ZI�I�Rȱ,�4�idM�d�E���E��4Iiid�"�d��Z$�"�$�H��D�Ѥ�Ii$D��d�d�II���M��I"M-$�I��H�-$�Ii�H�ZI4IidȖ�ZIE��KD��M$ɢKI�"&�"DDD�""&�4D�D���-KKKH#��m��B6��B���F�b̅��l�[bl�؅�!lhA��p�a��6hLhChF�!���n��jʢΦ�b�!0��؅�!l!	��4q�2�M�-�1	���Bm	�f��p�&h[4&hX!fж!m�X!m�fB6��bЂ��[���Y��B�!	�LAfBbd,�CBbhY��І�2�hLBhM�psB�Z��-��BК�Y4H�hB�#Z$L�"h�4H�Kn[r4�dM�5�Dj��hɢE�"D"D#YDE�D�D�"F�-��X���F��H�H��4DkDD�"""D#H�"&���D�"F�D�D�\$H�$MD�"h�"&����4"D�D�DD�4h��"h��",DDѤY!D��""""#B$B&�D�D"D#H�H�H�DMF��"&���"h��4D"ȄH�H�H�i�H��H���!D�E�""k97#H�H�$M-E��D�"�"hMFZ-	��h�h�"h�h�DY"��E�4HM��h��-���A4H�YBh�&�h�E�4Y"A4H�$Z,��E���"E�Z5:�u�Bh�HZ4�F�E�E��h�h�&�"h�Yh�&�!4YD��h��h�"$Z5��h�D,���--��!4i	�ȴZ"$-h���Z"$-�!4kB����\�g4i��eК4�Mh�Bhɢ�4i�4H�F�F�$i�4i�L�К4К2hMhM�hM	�M�hM	�M	�����q�FMF�-mF�-hZ�h�E�hքі�Dдi��H�kBі�"hDi��M�4"2hD&�DEcMD��M&�!4h��D&F��4"	�Z-F�i��I��ѭM4Z&�h�-4ѭ--�i4��-2�4Z&�Ѧ���&�}�S��)�b�\=hS-!������v�Vf�e����k{�@�}�_�3������g�Os�����?��?K�w���q����䲈����t1��7����Zs�3��&��ܗr|
��Ą���w�no�ܟ����� ��>%����?�/~ʣ�AU��|��������ʃ���H� ��8�0� ��Z @	@���B|�������>�C�W�h�J]�~7@�q��b�O�������!���~Q���ꊠ3����>���Qr��CBXP��l��
]bB��7�?��D���t���"�H�ۜ�]C�S����6>W����,����/��?'��n���f���:ٷvf�:��c3V`�f7��3�Ͷ-0m���ƛ������5?Z����j����軰�'�(��L�>C�����`l��`ƴZ66�H��Q#cmA�K}o�~T��}lZ�S��k� }�Ң"����~���O�<!�W ����1���'Т"��~���1y�?h|�A U@l�{@n�`>o��g_�o�_���������K���/�� ~D�[��R�����O���������|����g�?�QT�l��/�}�#����i���t��~l����   ݟc��*��O���� E~���S��������r�1�u����C�v�u?b��D.��0������#�R��������d�9>������6i*�4����)�>�B�Ҩ���M�G��ѴK�?����(N�稔'�����A��Ȝ��?W��_Y�|��TU�����К~����������><��_e��0}W��]-@A��>�T���'�i~����џ�đS�}$�������wQQT��n/Ũ�?@C���/�_�
jj����)���j�e
ڲ�2�
ڲ�ee
Օ���+++V����YYYZ���j���+VV��YZ����+j�j�VVիjյ+Vի+ej��VV���+jյjڔյjڵmYEjڲ����+Vի+)���++�YEe��յjS+��b�X�V+jmX�V+�ڶ+�V(eb�MYX�V)�+V+�j��b�X�Vح�j�m���X�V+�m[)�j�X��
e52�YL�R�Ք�����j��j�Z�V�V�V�[j�B����mYYMAY[S++e
��L�Y���2���jիV�Z�QE5j�+VQB�Q[R��V�ՊԢ��5�Ԣ��52���յ�V+jڂ�MA[j+(����MAX�Vjj�b��X������mX��+��b�X��P��X�V+��b�X�Eb�X�V+�V+�jj�b�X�V+��l��J(յ
j+(�QX�[V�YB�jՕ�V��Z��[V�V��5ej++)�����ڊe52�ڊe�MX�Jj�R��5j+j+P�E
+jj(QB���)�SSQZ�ڲ��(QB��(��B�5���������eeeb�����YYY[VVV����������(�YYL���YYYB���2���QE5V�Օ�VSjjef��V�ڶP�j̭��j�+
��P�EmB�mB�e
+)��B������VP�LVSjmZ�SQF�VQJڍYEe5j�5a[(���mE+jVSj(+�
�b�+�
��AM�+��b��X�V+j
�b�X�V+��mYX�V+��b�X�V+���X�V+��b�[jQJ5mL���Q�+e+(R��V���VԦR�+P�
�ڊ��+j�+jVV��)�Q�J2���P����+(�R�(R�
V�����j+j�ڔ+(R�+(Ք����������eeemYYYYMYYYYYYYJ����ڲ����++VVV�P�J�B��eeej�Օ�V�VՕ�ej�Օ�VSVV��Vղ��
+j(�j+VըP������c�~n���S�"�TD\|�Ч��}�&��>�:��3����NE�H���*����������(��۔���ͫ�A����ê~��+�0�.%?�	��ݷ�d-��4eQT'?�~߭~k�7�*�i�����?1�2����������?��x�> ���@j$�~���V@lz��
���J�/�����A"'�X��[�D��6A���~��S�|��	�O�J������u�����]���g��w�d?bU(``1S��'?�rE8P��b