BZh91AY&SY�d����_�py����߰����  a2���   ��_@        Y���   㻩��$� H�*AQU ��IEP�
T P �^�Q����p�Z�(4� ��   @ �       a� @/k]�={�{�l�����_<��w��o{�U�uuG��W�Ffٓ��#w�= ݷZv۽ЮA�w��]����\�b�7��U����z��.å��nf`Z���Og�� Zrz�n���e�7}pziO�}�2�$������[2���v�[��	��w��M6��
Fs�Jtn�Ҫ���������x�f�n�n�ͳ��ݯ3���MyՎ��b�m6��h��x>B7p  |�yl��9�mvM�6f�[�Y���z�M��[=���I�e�� J�K�C���g�Gq�����,��˶	wy��y����Ή�l�ټ.�4�  �:0�o>��5�Yn��}�K{6�S�ۭ�.�s��{ʋ< ���w�Z=�G��q����%��n����yJ��%������/ x a�  �Cޚ�
ަv��ڃ}�;ݞ���{�t�������3t�m����W}��u�����9��v�q�9J�k>ܥ����     �  P	Q �    
� (  J��4g��*Q��@�4��##&M�j~�D��! ��4`  �0F���D�*�`  F� L ~� �%�����LL@��a L���=OHʟ�Sҍ�̚�M�(
�!�*QF�PcPh� ���� 	���?!����4�R����ؔ�E@i�-_W�6��I �� ��R�C�q�JA ?y�B��������BG����7��W����j����A" E��І*��IAQ?�����)�>�.I$�H	���Q�C��g��!�g�?�����ƍA��L�g�+��+�]�A#D���	�Fd�x��,�	8$l���f!�Sp�p���$����p�:�L�I�7��8C>�߯�	19�P����<��$�I��x�ȝD�5(M7g�q���=�L<p�"{�WNɂ-�iҶ%�&�DL})��X�7r��D�WvV	�:&>��<�_?c+��̑�%�
�G��+�~���%|��N_DѨ���_%��9�JD}�se|�ڕbq�H�nR"ܯ*�s�%"wYXp��"9��At�?DKy)Ȕ>�}�5)��D[�y����^:<�������䮉o�"Z�O�W��r�8�Ok+�4��%|����8�:�R&�+N>�o�JD�r�<�����ҾM�����J��R&�֥'��+���H�rR'���~�wӃ��be2�K9�}�'Jd��G]��gYT?h�U;��g�&$�T��t���E���x{��&cU���+�d0��t�ږs��9�3����D���U|�ϻ�eW�����<w�)h���r�#�+OQ�ɩ6z���>���N��Iѩ�O>��5�W��Rpt��&�UVh�L=��u�jt�����v&����*���H"�4r��L�#�m�?'�A�|��ܦӖ�6�{w�z��vl��T�L�K�v�*	���$�BeW�ʕEr'��j������g���U{ݪ��Ur�q�U�U�j�;��J&�@��������[�y�bϠ���!9L�}3#�������N��y�N�vW���Љ�C�?�k�ѻ�>�y��1��	Hv��T�7r�A2�I���m��v7:HwS�kߥ�v��ڲe�{�NT8N}BH����M�M�t��jOh���<t�:'^��͓�:�9h��$t��Y�_>�\*$��ľ��u&�|NY�9�:�/O8G�����!��Һ���M�G�!7�3�I�~6�q��I��9�W��OC�bDL���8_9'8Sr	7'�8G$��Y&��t��} ��3�Hc$��d�=�Op�=�p��|o6��Xp���t�Q�"P׉ҍ���p8��hyI�Ie%2N2pNq"jx��#����B�~�"o�h��ߓR�JDԱ2�(~O"Q��7�4�dR}�?`�d�~ϓM;Γ0N�������8A<�tH䉂s/N��搿�t�M��i"&�D�����ƶO�2��N���K�H���G~xO��2�$8>�M&�ç['��DNa��"{�&%�!0�Ğ�ӥ�=i�R��N���҇!�i���P��N�D�O�6QA<�I4��&��y�x鍓�f��
�DJ�DՒ��
����Dt:P��,DNq"`��rH?%��S��$M<�&ĝ87	�'�O|���t���"'��7xl�!>��}��)��%��4�a���#���� ��"#��i�='D�
.&�%%��ϊ�'Q;}"jh��}#�=�>��`��r����$��9v�؞��<wӖx�9�'����N�#SǙe2Æ|�G�Q0y0K�54�&���v#�'*Q�Y�#Q$Md0~��Nϸ$��K=�Cp���x�9v`��:�K8�U���Y�:�Hbbe�=¯�u*��#iXg���~�
�}ڈ��#�I0O��xm�N�p}����v�����ީq��޺��?�=��G�Oz'}�:s�Ǽ��dr|�ۑ�L��XWD�eM5�션J�!#S��y����}3�8a�x��*"9,Ly'
g�x�"#�DE�ӌ�g�#�Q<[!���ba�O��*�#}��"�'fT�UDGݨ�Ȟ�x���ȋʉ��">ډ�OyR�y$O�W��TD}ꈖ�(Hz��A��dƦ	�q0�5>�����d����N�Ȉ��*&��(Oy��ϓ�T�&�=S�<ڈ�ƥd��*P��R�cSD��:A���SN���#�����t�1��>�/ܨ��Q4��B{�N�v}Bx��(Fv�&�j"_�A��N�����R�f�D��:A����8N:rD{̩]숭N���[S�w�8^��?��к ܢ�A���mẂ�O���I��#��P��2�{��$��X�z��Q0]�:&�J�ީ��ϧ���6�D~D�ښg"x�Z�M�6]O���x��w�P���7f�J��a�=$:p��O�{>C6|�Y��3�C�B>����xG�0M��釤F����y´N�SL�N�֦	����Z�/�8vJ)9��9S���'�g{,�lC�_1kS,a�VQ�J��wr�|���|r���ɧ$9ճ���߈ϗ�Vg����1��3�Y��d_>�ͨ�Q4��irar<��G�S��G=Q}R�ԭ�=R�H��r>��Qݨ��52�����ljU���Qb��T��;R�U��+�a�j97�_L��N��r�W�#����v;�r�[�N��s����)}{��X���,��yc>��>��1k4<��/+�{����u�v��gO�C�V�'�]}�x:�T�S�����϶�6��[�G�g�<�~gY���|�����m�/�꽥9v��ͪ�f��Ź�}���j���5�|��0��I�ߘ��^��G��y��	�9�V{c>^��^����y���X0k��
��U���JrR'L���Rh�e|����DL�"pvId�G��+�~���%|�ģ��4j"t}>G��(�rU��"9��~ʕbYoe"cr�E�^8U�H�N�+?"w�͕�ϺQ��JDv%��o�JD�r�<?"#ɧ���JD�^�W�����YI���|ܤNDO�h���_?,��8�:�R&�+N>��o�JD�r�<�����Ҿ~rR'3��%���k)<__W��D㒑5�a�G�;�c�8P�&S+��>쓥2DnA:�W�3���j�vV��؛sT��t���E���D�ؘn5^0��<vNN���s��=��6%���}��C��Tʡ�Z�������#�b[��f���$�ˈ��;��5&�Q; �G�rD�������O})4��U��T�GIGj�4vI���8�T�SǤF��ț��5U檌<�;��i���G��}�2��vC�#�}7�vsr+)ٜ����������N�=�t�;O~Qڍ�gG�[������=�ֺ��{Һ�{����F�k��[�V�H��v��^�o��~��.��]���]�闲��Ӝ{�t�q����k"�jp�����<�ŏ/����w�y��r{�ل�{�E��O���Qa��O����6��!�!�!W;$��;EIi�	��55:gJһ���=�S!�<�߭:���O�iϤ�}�՞�v����Q���P��2��O{�w���K	&�~$4�����E�c?�9�d��0�3�a
�pi�[u���|��w�y��8�֘k�`�hxly���}�&L0���x���i5�џ�A���_8t���Lr3�)�0�g�:��/<����^i�\hc|�q.�0��M�ͽ�c����5<�/��>s�0<t[[)���t��<�m������N�|�1����чʅ�1�����qS��d�4�v}�����N��� �q�ܘil8�7��ϖ�1So�-��i�󍻻�O�e���n�9֪Z���Ҽqn��ۊ�xe��i��0ȭ/��FXly�.֨m�X��a�]xy���m6�<��C�y��m���N�����6���}u�,�G^~M��
80��~el��+��-m���>_ʓͭ�n�^ml����STL�SOl� ;Z^���6�:|a�N|x��;��x<��4�m��u���p��:�m�ו��3ۅ�:-m8�� �m:����i�G|ۏ��f����d��ä9�歷�c!O�tç�@��Ҍ��dq{]KiŴ:�#Cm�;��#8���̹�k[O:�,�`sM>��xe0!Hqt�I��:B���K#�Ӹ��C�����S������?_�g�K�@Ҍw��ݵ�8�J���:�O��_,[�זqC
3ْ�@�Ҝ]���'�>m�Zaj�q��i���1���ʴ�a�Xa����F���,��qhc��Fi��|�]3S�@�Ha�<����:~}�|tgFi����|A�������R�I��5٤�d>�ҋq���!��O���9Fa���&�|t�����t�����]����B�e�T�G�{:�n�Q�}`A�4�vt����oyYm�l�T�o|��<�N�2��cܼm�֮��NK�6�j�n��L��J��~�',��O�xæ���i�S� �}8�������	�+}�4�
�w8��kw��u^�?zx�L)��2��:q{d�y�4���j�ױ�UkiS�$tP�1w$����fM��E��=Z_�|]>!'�O�ӊ���	'���D�����̐�"]>>:x�@�����<�Y=���������>��)���T��<s�~��?�Oro�D���!Ν=���ç�����{'�g(iD��g{���X*C��9{�|%;��./�źHq~��i��@�N-���y���sM�O,�R�b��e)�Ӊi�N�E���?�)��*���B�͖YϏ�!�ސ�s�NaZrzqX\��8��T���qR�X��`Ҧ��a�Nik�+����S��{�U8ӫT��w��;���*m�_<���=�⦝q�\`��^�>�8�m�8����v{�! gZ����!����Ϥ�Ϩ��_�<~8�4�/N��ZUG�zqS�M8��	�_�������L-%��l>y[i�k]��m�:�e��:�̭�[W�B����4�)E�t�_>4��li�)Og���ӯd:|x�:O�!7`|w,�7��9ྌ��6�̎:��u���q�l��K�Ǐ�K#^s�P�0�g�w����wd0�O��)Oqkym-m��n��ͪqn{X�i���[�4�Ͷ�,�8��y�t�c��a��ύ!���␄>4��HS:a�;��F}�q��/#�y�^q�Ze�g�1����9��w���HC��)JA���'`Q�Fi�%Q�>�p�Γ;=�&�
?M��kH��;�Ҥ��u�e�mm�����J1�c!������h�����ky���u�e�qn��,� g��f})����|X�Z< L��Ӊ@0�a�0c}���S�����ز�����|`�oge(�@�f�7gn�<c��a�Ze��:���Һ:�4���Ə�Ό�����);޽>�AAO�;��t�x����}��{4���┧�n�.h�~<t����1�x��������?���JtL�/��am�`���?�t��e�Ǐ��~�?Ze�a��]4�]�k��M7{)�<t����8_' ܜJ&�Be��
C��x$��Ɂ�臘�0�xD���f="���&<2����2�l:0Ъ��n��*�Btf�{ӧL!�d��B�:s����}���D��>;G~�>�=)JC5?�ў9�>�f��:iO�Q�>�a�����
B��-��?-��ت�8�������'HS@æ��T�!��3�ó�?��BS��Ҟ)~���ƽ�������ƀ�;��hߧƟ$�v%D��a�����l�H|4���Ŀ��JCǆP�Ν��>!�͔�Q{�:xyc4���L=;�ftf�~��tJ	C��'��aO�'Ĺ:a��|$����SW[<�ӿ�a�> ���RP��R�'O�c���q�q������cH^�3�!Jh�Oǎ��m焺�m-�[,O^Zm�^a���ӊ���_6|9�>æ�i�c<iE�����}�Ѯ�a=Ozdޱ�e5u��cҚw�X���I��=�l��>0��؟�a�>>��0��I�w������կ��h��MN�����e1�3�)��o�:�%q8x���̘`���S�57l�^�k�L�����3���x�c��Q%����tA�O2�)�f�{��~��%���Y��>�������*�0P��0۬��q���8�3���;�c�*��N�3?��'��͏�K�ӧ���7��o��Ҙfvz���T��6a��fz}rC��<��y0ï�.|`x���;$><xo��&�� �@�M>>:n>>��2�O]©İ�@�G{4f�fҘ|SǃݜK��}��쌃rt�鞸h�s�RO���{�T�|�x��v:�{%��?�ݟA��Xi��њ~�'�����a�:Cg�=��ݚx}�`��Q�]&e(�K?<��Hiџ�Y�ɝ��9ӟ��ҝ0�di�\�qka��I���r���4����t�0��y݌\�w������A�i��0��q/�x��Fa���;�!�����l0�PgO0<5_ǆ(�0e'{8�4 f�e�Z�k<�����wW�[J�[ ����M���m�w�Ǖ�C��#�|�������L;�*|zd���M>)���4���}+��ZL�}vZ��<A���:sO:�K�����O�q�1�y2�tZ���~e�C37l��l�m��Iz�4ێ2��	�1S,<�<�O0'SL2�Ӎ\��m���̯�~h����
��/��~?��|$?a����e���W�!����?O��V��"�VT�@���\Br���mBE0_���I�"��������q�N@Gps�R�r H�b��&"."& ����Uv,�r7cV3MXZOjQ�My���p5D�ips>��P3���5M�k�Gc
es�O �U�\��{ �s1&�QJ�CX(�*����*۱�D�-���+QY�l�R��ꄗ����.�pZ����J�@b���ky5B#A%S�U���U*4\�-]b@5SR�
[��L�r�U3r��ZR�ZV����"cT���f�Q����.��B�L�Z�̔y�kG����v��%/�sNj�8�h��q���k�8)U�G�r���*S�\p`��X�����8���Gu.P{Vs.�7����Jδst�5�1��p� �5`:�*���~�VS���E�p;��Ng&�AZ�<j���o)���W�3�tQ�3%2�5�,sX��Y35���Ϩ�ND1!����kS
���!pѺ2C{Ūn�p�9�F�B���k?P%��q4Aj����E�3���تv�f����*-��z@�J���"@�q/����q3Uv��ȩ�����'ܤ�/T�"E9* j.�T���*��r��yT�4��YWpn!���B��#�W��wwύK����~ƿ2��� ��{��a	�g@#�������2�����O���{��4AJ��@?2(HbB~Q)�?��9�������*�UmW��yU�W��U_"���UUU�������U_+�V�^��U|�UUb���^*��x����j�U[Uz��U򴪮"��-*���U|���n�qZUWU�UUťU\ZUUŧ��9�k���j)j"�C��-��Bb��@ņ)X�؅�)ajI-b�*�-#ň��Yd����>�����U\ZUUťU|�W���.�\EUUU��ZUWUU�*��x��U�^*��UU�*��*���U_+�U\ZU^�ګj�V*��*��*���V�;ޯUU�UUTUUTUUTUUTUUu�d��@����[$HKm��RU�"�$E�D1@�
���b�$Z�ղ�aI-[V{e[�]X������������J�U_*�U|��U�+��^�J���UU������U�iU\EUUX����������Ҹ��UmW���iU\V�U�Un���UUUUb���UU�iU\V�U����}!�G�>*H%�lZ1X�KV�T/񄘮�W	��'�����߿uW��努��*��UuU�UW��UU�*��x�ګ�^*��UUTUUťV�^��U|�ګ�iU\V�UŊ��������W�UW��U�W�ҽ�ݪ*�����*���U�W���[UmU��}�>	>��
�Dj$�� H�" ȣP
��2(��Ejk�f"��� �$@�B����VI�Q-DZ�R�-��Ғ
T������@@�A�?�?�@T �	!H������������_�?����o���l����2�8�<"&���D艂&��&�� � �!�HpN	Â%��8'DL�LD�O%	�`�""i���D�4N�tDDN�A	B'��Bh��0N�bX�pN	DH""t���B�B"tD�h�&	�,�Ĳ	bp��(�Y>A�#$H"X�G�'��8Q��4�L4L4N� ��"'DL4D�0�,��� �:@�HtN���}g��r���r۷�L�+d-���v� �H
�Q�H�C���Z*���DA"iђIeHQ�2�T�� )x�%mR��tM�&�UV��P(��*��U%�ʘ7j�j;GdH��\���ZBDլD"��d�i��Im�v�Y"!�AF�""�&�PCRƣ�����t��(��n"�,` |qF�	P��k��ԥ�Y!�"���bj�MAUe��F���d��"	,�*�-vId�$�Ԉcbj���"��땧�(A���-NE� ��G�u���QFY��ࣤ8H��8���ݶ����:�N�jF���銡Q:���7�VG u4�`�Tq��+l'�v��>ZXKY	j��)k�� �-��8D����A��yJ� A��
IX��ζ�M0�P�4�%�RI]d�"[�9SMG'(�q�3�N}�Y ƫ+rXݎԨY��5Dܪ�+���c��d��P��W�&����"�'Q��d-�LL9)I\v���Ɗ�2�
DrZ'l���P�I-���ȣ�H�(��*�U���,�V/\�����Em��|trҡ^Q��뵁X�U)]v"VҐ�HVH�mh�+c�a��WV�n�ꡊ��l�8������G
�X����PdF�u�
[�ZA�� o���NM�DՍ�\N�}f<�,+���ҷk������ٰbh�q�kTrE��.��b�8ȉp�#��:8����c��b�����5"�V0�r��v7Uu�F�����jU4�R�QT���9,��Uh@&5uK`ӕR��*��0j�S���@��G��3*Mh�j8R!U*���	�U����D2*���hU:�Tc�N(!�U
'Elh��d� tl����P���:ԎFAWe�![n�P���И6���N[(��"lV�Z����GBp��PT ʅF�s�GKƕ��L����RUcQ��V�,P�TphMDXH���)��,dPhd�7kT�~��(ख jZ#��X*��
��,�X�+i�m�N�0�qZ�J4�|��p�m���Ƭ"bc�[t�����i��J�r#P�H1����r@U�eVט��]$��]���`�Za�vf_"�U\n7�-��v9��d�9��U�mX0HC@��WZe(�jnA�Sr�RzAJ��#�	�B�9�u��em:8B�,����ڬ�nr(��+(��B�BH�e)F"���YEUl�oř��[@*�v�K+mF�N[�9[h���ԍ�k�uKm-L!#� � 걹vV��|��#@@J*�J�p"mț��";`� �NIj�����,�B�,b-�V9mN���J�����܃���r�[�n8�ڡH�A�Ƙ�Q�K��"P�D�m����("�l���*R�G�DID�V�N�mN�����9�1�6�u�&Z�]R��qZ����R�R��8����Xf2V+o%|+�I������UmrZ�UTV����	c؝1�|�5i��q�O�K�pE�bh�n1i(Ih)b��P�KStv��DܖA����q�5d�	���R��u�b�B�F��IBJ۶��B2�Qʧ,��7M���P)FZ�M2*"���*�8Չ�;jj���9SqUk�%T��"ăq�Y-K�"�x��dF�	-�����juKtNYeac+��Y#�hNY��	��GS䪫d�
Q�u�0r��
9IF�*��%	KilpC�UFNѶ27I�KSVکmj�l��XԱ�HX�bh��GY)K+
��T��Ch�v u�+M�&� �F7
�;������MU*�%��S��R�HH�Mһ�R��6�jh��XX���iԜ�7ʣ,��(&�F���(�*�$�"$��"7Z�`ӥ�U �(
���H�V�l�T�0i�	�8H8�E-�2�Z�I��VX�n�Z@�VXԖ[,V&��;Y��Q*�uV��9jRV�;"�:V�	l�H�ԣV�6�i��]t�����AZ떏����Y� �Lu�V�L�K![��UV�tL�R�6�v�����F�뜴;I1K)�F�n!W�'etR�*ESHrNIU�*)e��v��
�1���7h�T��2�䔰�U���������RU��:9b�Yc�,d��UJF(�q���B��D@	�J�XWv�Rv�x�00N��c� Y!]���9�aʙ��X0�˶�`��*��L�I�U�^�Z���E����ki�NGVc�V8����r(�EU"m�UZ��A�cu�8�h�6ԄQ�؀M*�#�r2�P��H	�$��9d��$8�%
�����T9F�:WSj2Z�r&Fs��7�R;gJ���8�)c���(��������b��pI�뒃�d��9T�b����k��V�*��I�j��B�HL� �N�N�rÄ�5Un���Vڒ;��"dp�H�v�S��Wyb%q�*��8Q�8�#��6��l�D�;+!!��Rq�[	)Z�r���MLl�m�*�	�H�E�X�728̼au����3�Dw��~�UUTUn�����}�J���UUTUn����}��/W�,UU�Un����}�/W�,UU�Un����}����>���~+���.�u�8㍸��q���T_��~͓��o�e�Z�v6qµ ,E�Tr�C���i�ix�:H�v��Lc�	#+�9#"���
�-��*�+%a`�UZ�Q�7U�(�l�ʋ�Rګu���#rIX�Z::ܩ�ƓP*j�I`ێGj��I]���B�m;Ec*�-�9Ec&XV��Si�E�k��y����"o�[�Q�J��X��8��*���A�X��PTCn������W�Ю�bU:�"��;s�Lf^b\���n)1��#b�e�2I��P	�$,�j�ҊDے�1أN�I�*�!D5[LjYVI+rB��L�]�	��-r.X�L��/N9ʆ+X��q��7\��UjA:�D�l�P�%*�I��GhD���$m :���V��q*�2��d�ae��Il,����
41#��q)�n9��m�*"��U|��c圍����H�v'+b������'P �s����[{���+_�����N�Q��p��nx�;�/o��y�?w��9���=�����s�������m�o�H�6��qH����^�O�ԧ�,�ꩍ����]Ro��=r��oS&b�s5xa��K�+�7R���:�0�brK0y����Lm��Q�r!V'�o��w���P��sx�;������7�:�z��ߏ�Q�l{o�6�@�UѣřZ�~�n�܍�jkBs��4�!�˴�ḯ���������-��������m�޸ӓ��971.���%��������%L��&��Iwr�����'�`ܒ���I�A��fI4u#�ͮJL	̦O��6Lp��㢝C�=K�h�����k�{�8��~���7�v�z�o[�.�	2ZZsOi�pG�9,>�l��]!T=��!�=E�}m{w��w�-+��z˯uׄD�4O%i<p������N��.�����9`�N,UX K}L�̔ˉ��{*������+i���M:zS�VJ&���ô_��%ej�Q�0�@��co->̐d�V[P�r'��6.>>dc��a�i��U�۸|��i�#�Ѽɘp�a(��bZ�k�I�B�g�2���G�S�SML��8af~<"&��x�(�Ha�]^yd��猰M�x q�}$�I��0��Kb�产��qݎ��f��$���������]�'�-��f d�ӷF�F�&KN;0L��B.��9TUS!R�0�s�o)����|̪�=6Sie>+��շ8JQ㱿�������8~,O�xDMD�Q����(<� ��[1a�u�&Jږ�@�3^� �뜌͞ϻ�w��/(�VmV5�J���Ge���}��"�yn}���{{�fo�}f_F�=���Z�Hc���l���s�1���̇�U�n銼��'O_\�b�<a��ڈx��W�uνs�vvv]ʨ�/LTK��n�+5�dy$�E�"|�Q�Vs�詹�Or\f��2�Ö��v�κL�0b�	��v��I�$���'�p�r��o	� p^Q|��巘����g#9��7�V�3��jFs��WV ��Q�H!���4w��Yg%U-$�So��V_2�.<i�_8㍸h�0J4�x἞�{[,�9'*YH@F��eJF�� #������-Ӑ��q#�~�!3���+�b�������4ഷI�'G%0�$��i��Cn�9�$%&~Nt����Y�N�fI*[vQ�+2U�wDtR}�Sn"�&��AI��%�ғP��'>���.�bj��bLmݲr�XY��$,�fN,DO��h�`��Ha�
�Ih�o��������`�f  ����d��V)}Ƶ��H�O���f^I}�B��J��J�S��Q�pJ%I�&D�iY�1g���f'[0v�:���S� ]X����[nf����H�h��u6��rc��]%LUyNL���HϜ�L�l����2���ܴ�q�cA�F�Е<.2�a���.OX2ڲ�.2���'�D�4L0Hi�0��	����8��*�x 4$%:U�STJ��au��e�&�'��_�ܼ��^�=�7U_s�繛�-S�w�RQ^��M�؈��ӴJj|`ַE�Z�*����ݐ]+n��F�5� M��:��n�I�`_���*��7���/H94A��L%%��>!g!��p��OǄD�4LCM!��}&�I�Ga��cG^T4��ׅ��6�z0 �;��9ޯzorY=������>��ʮ��]�,U}��g~_G3z8��u�W��n�w���^�Ι�9%��M���&䠯c�E�ͱg�ؖN�t���}S�V?�O���̋,[���.[f˿>3"Ő�����w��n��7%s��5>ڤ�{7w\����̑�j�(�5�䡇Td�r���_a��d�y�h㔣'l�9�$n�]���_� J�H�))6���%�Fw	f\�8�t`�4#G���.�ᄯ���!�4r���%Ċ>�����̸�71%�s-������a����R��fڸ�Y~�L��2���m��4M��Ha���~��YUH�;y [��⋼]�ET_qm��3	.7%���M�/��(��-cy%j��{���z|�E��;֊p�Jp�>J4�}�&���
i�&���[���3�ѵ�PR$��/�$٣�(�ㆈX�4ofU�$���`���'���k��>����o�����M���g��~_\ŘA'���������G�h�~'��ò2xa��<X��'����p�'�t�'��㌛<;!�'�eC�GjHG����CĄ=#���d<L��<C$�<[�h��n'���Y��^+j���0�W�î1W��ux�^:�W����|O�'���Ǉ��<>8>!�x��x��O���a<OD���O��><5��Ä�+��\�%$�S��;r=<>'����<O6)<�����x����3�����O����g�L�e�>������bˏ��H�9.�K��՝Z�V���Xbu]\����N��Vm�/W�}c������|p���<;xHx|O><����̞'I�x�׎2l�솉ru��,��^�j���.׫U�ez����Yb?0���*��д�=��e?��f���e�����������{o{74Z�w�p3�ӳ���gj�Qfj>}�x��i���|���o��b��'�~���ض6y�W��qSb�{&Ⓧ&�o��;���G�{�<�����&29�Q���<�;Ml�z�w�J�pW/%v����&w����s{s����{���K�^��	�����I��w{ڋlyf.������Ŀ�9����~����{��~�{���}r����8����}���~��*���9�?���>ݽ���߷�����ʺ���8����7ww���������߿:���8��|�{���y~��߿~��?
��s���)�ն�m��6믜q�Μ:|t�x��,��d�J**-%6dey!!K�l��'�,���X�$_��Xy6���~�Q��F�1�H�KKKIc:�Df��d��G�/H�R�E�uLM$6�pY�I�BS�ͨ�_�����5an�,�jV�f�h��zGT�!��
u�����i�v��r!��&�8����-�]ŧ%�X��wK(��r�䋒�%��$*/H�>x� |�j��d�R��8��Mt�j�$�����s(�J��EtM)��R"��AdM�b�IJ`
,��K4Y�|�m6�o�p�+l����-�`�i��reۆ��**+BB�Ѧ��D("�lŎ�
0Ģl)J��՚W|�ۈ�)���|���s�kE%ب��J�-����Wk�I�n��N��9qYOe��A�D8`h�)��R��&���Fb���Yapj,���LI�aP�b���L�������T4���@�B�t̖��컼C�n+H���C�8�����Pj��]��B����'ZW=��ǆP�	1$+D���Q/Ƒ��n#�	ԁ���l<�MT�+��p=s	�-+�	�,����h�&����K6@�5�y�,��.K�Q�4���3�LK�>�j�����:���А;Ňvg����r�/y��S�E�^'�Ϩ��}�Va'�޵���߽�[���{�sϮ{6|�Un}.�i��_jϪ������~�îa�|���m7�.������������{��Ou��,9b������OvI�9R�=��^Ul�G�A�v�s3{�svL�}קRw<n_���z�>���Ϭ��ֹnOn���N��>j���6p����;��^ံ1'��8�z�&��0,̐�T�\��8@��B�S�)"�p�5	$�堙�F��+�H�@�"&��ʫ_�qS��!��kC*�T|n�.�S�ZClWFW�qM�G�k�r��(���E&B쁧q����� ";1�����_�����Ŗ |;�}� �"�H��Hi*��1�.�R44�'��I"��/���[�fL�-'/0�_3�=��?EL)bȱ^+�C����<A�C�i)C&�ѦV��J/���a!�ӂpK?���xDMD�44�"p�f��r�c25"���Q� �/����`:b8"�b�bj}(D�dZ!x(�r�����+��cf�˭�U�r��%���	��) Y���Ғ! `0Q9�Eh�9
�P�,B�D�p犬�h�Hb!D��M�y���)���U�'z�n�ٟ�3x��1��N;z�����
8�6DK � Q- ��JL��=��U������6"n�B�.`�X0<b3�m���X�Nd�A
zQD8�ӗ%�X�!��bO%b�O�We�\~z���p�0M4�Q�q��eC�T&[pn�ޢ���$(�I܋wp�6`J��ʤ���B�,�֝���������G��,0}�im8h*.�H�48 ��UJ��q20�h��&�pf�S<vP�z�!*vm��Va��?2}�Jҳ���*��s�>:��&NZf:��ȳ�&��q# y�Q~a�6D }�!!
��*8\$�IL���\Vx�ʛ��I���a="�X� PQ�����$-wt}�-�H|�ed�v�P�]�ƍ'"�T�Hf$0Q��4��ۗ[��U���&�`�rI(۔�Yy���@��(�4��ܞ��z�/̺��?��8�n8�N88xNV\�J�J�@f�/dɬm-���Y�H��"���$(�/��),HY"۶��'$��!)pCI�(��ڕ������hTl�^k�}��}�yo�n�.�x������luV+8^3!+�C[(�MM� B�!��G�#��š�u��*|PY;�%+��1�!hq(�3����@��k�k�7�%iZ�n,�*R�g�̘X�,UjK�b�G�oQF]�b4PX@�>(�4�6[�a)x��e��!撎�2U�"Z쌛�$��rR�@�Aϻ%��b�K\�L"e�a�zW��l��O�_��8���H~4�Ӹ���8@�uŃ�k��%�F��.Sz���Os�Sz�o�� |߾3��t���7,���I�ڴ��>�����q��	�sI�}��_�3�l�J�/�����|���{�w��g�s��{���u�{E��l��/��f�}�zxܭ}����=�z�4UK�p��n�����ޯB}�s$��uw!q��Y��8\V���x�J�~&#
s�1n+YG(�'��ܠ�U��J^��'Hx��`d��)�Q�&�<�v��h�K�F�����c�i�VH�e-�LDj5�����n.� ��$�m2��M.�4m�a�YM�\l�E����A�����d��@�؆]�b�E�}�Z��$��ψ�aM�Q��"C��8^1t�ӦBa$7��*� w��n��:��Vs/7��Y,�sl�Y�ś����>��C�%���7(�d��Œl�����Ñ��L�i_�e����tO��4DLCM!��
+����BHL/��QQZm'�9m�i�B�iT0� J)��g�R���w�oR.�J
"Z��+՛��>�w2�Y��y�G��Ǉ)��I�Rʦ���Z O4��e8ta��h
H �Lp�M�Po��֛mh��n�ɜ�M�>N���'ŦvS�%(��}�����?��e�]�L�,p�v�nH��7�>��|��fd�QD:�R���i��VzkA�E�6Ra�[`|my6���^2qGb�=�j�E��s����J��/����)�q�߆'��������u�_�����m�i�Ͷ�:ҟ}�G��L�2�BC.� kE�e����$�;�̼���s[��x�8e�f�a�6��4y3�pSiޜm�����y)3i�z���'�%J-1���i�(��5�ۂ�l��x�c�7�l��3��(�
�K߷��j}���-���e�MÙ����f��8���ӄq䉴�|���O��2Rp���¡Yx�@[F2��Cdpb��(�K*I�BI���4J
�A���G�g昜��ǙR��,�^e2j�l��OX�Gev@3��	���Æ�r���p`��|[�]~|�6�4�f�V�ic^��-��J�n�6��c�0(��,���	�Km>�~�l��<L)D�Z�MY�[�2�����U	\��nq7���=r�aU�U�M<�IlxC��L�	nl����Hm��~$��GgV�Nަ���-��Sʑ�	L��O���2r�N���-k�]��?m�b�^�UFJ@��r�$V�J0�+e��`]HR@בo�+*Ϋ�e�Zx3+K2Ը�����G�#�7b6��Ɩ��d�q&-���l�]�7�Y��MC	��B��➝(��kD�~!�N2�?���<O=s����:x��,��g�x|M��W�bޯ���i�α�\�V��v[�;-��Vt��^�,�m��\��x�W��u^�U�:��4��ת۬N/���\~a��'�X~q�����u\^�c��X��<u���W���W�������<M�I�x�>!g��=4Ǥ��+�<HN�+$�(�O��:VI<CD�4L'������x�W��۬u�Yur��/K�X����x�����!�h�<'�����>65���x�0�Ä�l�g�.�H�}}.#�D�>�"xO�՝\����gWO1oVm�<^�ɢt�'G�Y����<��\Gć�uz˹�����:�s�x�^�í0��>Y��z�zWe���:�]+�\c�W�ܫ
�VVVql~a��,��<�����]����y����������ܕ���'{و���=�}�2���g/3�U�=[}ڬ�{��R���)7���Oni�?9��~��f�C�3�h�p���혷�T����o7����6���4�s#��vv�`_���^5���T�������g�W��>oƖ�^�^�7��+��,��#�`o��lY��w�z�&��۞=l������ܬ��ok���:o����o�{>�<>�K��4'��s�}n�0��۷K�u�q�������~x>�d��qt��:���mZ�tV�:����c��؋�z޵���u���%~��o�w߷���}�{��{ݻ���������ҫ�����~����~v�{���yZUW?~�?~�|�?{gۻ���ߺ�*��/{�����Ī�����l���]|"&���hi�0�a�z�˹Q����d��P��Q�AƠ8Օڝm�8�\��D��QW+��R9d��h���bmT�Qh������C����]q�&�l��"��XN0r�D	��q�C��B���VԬ(�c�q�T��eC�K%��6�`�q�T�ݕ��Wd���FY %�*��-"�^Ie�*`�\�)UH�u�%�"pv�+k���\��d��Q�[pRW,cm�D�m��)������m�d�Z�P|���-��4�lm:�*�c��!mE,��8Y+Q�K#!��X2�[���jQX襎�
�Ԉ�����#��PlQ��@㰰B('�����,�G$���Bi´P����[(���nP�����r��(���Z�
ܒG,BKZv�rYl�R[\co�W+M֠�[��`���*���,��*V
M�7]B�D�n�+U���ȣJ:�L��8"��Q�m��M;d����B�ؤ��'��b� ��8*��V���T�&�rV^+�N�G%d��9kcb$M8�n�f��F1�c }��ޟk�1���_��?f�s�~ǹ�����˺C���WY����=�Õ>��x�g'6�x���g����������[���J̪�DX��,w�Uu�Ok[�n�s|�;���x�A��)�-�L���f�س�G�o~��-C���F�Qd$[��qN��"i�[ �.��l�vh�����d���i��ĳ	�n��Y�q���Y

�����V��F���ͦJ6@��jA��⩅k	��$�$�烢��"YF(�"P��$Hh�Q�Z�Y�af���aO�SL���g�au��Rt�f%P�C�ϣ���ҥQ������(_��#Ta��ٞ,��]�n����F���'�qb�E�j|��Y>}̽s:n�I���g����Y�"��}$�`1,�Q��~V�2��n=u��8ێ	�hi�0�a>0ٕ[�|��n���nT։f�s#�1��%J���Eb,mYY-w�?c��)�2�!�.KWeU��ZB��"6@0�R=��܅�R}�!Ѝj������J7�wU.��Dm �١�	LSiE�F��.�x�N�/όXܰ�I�����<��,�8��l~�#U�O���ܭǬI����q6��mH��>�D!�'���fX̸C(�v7���$���S�/�p�|�h���Xq���m.-�
�\8h@��$aA�I�׌*3ot��PQ��P�lS�f|�M��I��0��e&Ԡ�(��/̿6���θ�n8�N6m�iֈ5jA$R@a"�� �h�J�1u��Zֵ�%đ��*G��Pք�C�5]�n���^���f�SP6@� j#�IA�jRH��E}N�(� d�F$!�	I�M�ܻ0f�~+�h�@�$�M4�u�I�p����8�KC$�\�����s\.�t��ij���4Z~�=�P�Q��Tl�(��*�7*��y�RdB�&���&r�j&
�����d�j$2��v{�Ǘp�z�<h%)���r�tl�Fm��mZYtL�p�D׷���γ{w7�^��ɞ��O4�n��h=gő���D��IA�=v�&MK%��HB����2Q�Ş,�����<~4DLCM!���۟���r,�x/��>)j�ŕ]���1��$"D���T�Q��i b�7�캌0�M3>��5>�T*�4@��vl%�_�{W3���㚛�L՟o-�y4$�O��Q�m��[K>h�YK���񬇘d�2����'ǉ�ɝ� S�~�1��%'�0�9<����J�U��&'�U)��弶�;c�biW�k|�Ef�򞩯�U��Ŭ�Q��I���&�%q!��j�8@k-�L'���Q#I�i��y*�*.׊�K�0;w�� ;�	QqmS���
K�R�$1����%.zSJìu�I%���#�-�4�,4�㬶�����&���hi�0�������W	+����b������;��1��,W�b��,����1�I�,���C��{�����E����E��"Ż.���M���e�^rr��擗%��y;͛�]��+�+��ۥ��7����/^潾N7ܗ��{0�^�7�b�w�n}�U�}�9����0�|�����:Ȫ+&aY��׼l���4�6����,�';�Ά{,�I�Ի��Ry.�|����F�i��a������*�=cW�h0�d ��-!�m=m(�8��w�n8�DɁ����
�^�LL݅�K�Q�t����e���a�����55()_*KQE��������h��6��sG�j$�R��aLB��5K©>̓F0�"Lx��IADX��D�Ƥ�Ya���Iۅ�,��Aʗ�G��&K��Y������#���ZjbVHPQ�-�J/�EV�8eVMn��P����Wk3p�k��y3����a�4ˮ=~~|�6�4�f�V�:��F�^&�C*L�JK&U�
.��&�}�1��D?SD*DN�����#E{���4lxRZB㸗�S_x�F$��8@���ջ���/+)_K9��a��50�[2��NH�mhimd�t�
=�$r�h��y�Hv�D���M�&�B 2ꬠ���1���d�/O4��:�D��Wѕ��{�`�h��I�So��C)ģd���h�[<�X::Y{J�Fފ@�'1�h�����q��Ѵ��9 q�ލbIxѤ4�|D���q�㬺��_�:델�8ٶ���P�O��Q3��1�`$��	K�(>.�r�oIE�M�+�B`L�*be,�o4�����UHTK(�\��'�2��-��c��<S�9������t��a��b&N���"�HY/��� ��`�U�#�l�S&�R��*$߽R�J�SD2q��WK���.'늌��i��
\�s-ݕlC��x���E�CD]B�)H7���\�Se�N�]$1l�U(�h��T�]+v�p0��a�W҇�ڷj�c�7,0��C�R6J)�b%�RQ��T�x��u������]q�q�8C��eV��̨�1��*�1�7�7�q�c�Hh�h��/��{�8%��!��U�~HS��-2�"F�h�;�<��"�P������ݭ�s?�[��*�[�/M��7'�NQ���єH\(�"i��kv�5,+X4��b�c0�-B�I]̚����GI��-�8�>K(q��fX��B��@/)N���\XŐ M�	!�%�0��	�I���p�L%�w���40B��٤�1����
�D�`Q�Kba3�,2�Xq0�H���L�$��l���Sȧ[`��1'�&#œ1LE�b�x�<u�q���?��0M4��\(�>�\h3�4���׫2�Y^�Z7����1�4%�Y�2O�	N�I��z�����e����s߭����k;+���w���.�g�w纣�r��d��u)��w�Ǜ�3��w~���1�)@�UϢf��`<��d���靭,��{q���z�y�|<���P����ߒ�?|�(@uD �qx��bUQ�2��k#4P8vYn Q�>�� �+Arq�˽�34�t�
�(@H�I#Fs�c[:HԌ=�
n,fʝ��g�v3�v�}CEnP$w��R�
9���̕2f��G!ÈV�2�<�P�ZK5DH������X�;M9��[��.j��Z�Vqd"�ߤ����%�с2@�D�4@�G)փ12a�R��ua�Q�Q*� �=�'_z��p�~������q�VtUV����b�$w�D��Pq�O9-f�!A���^?<u��ϝu��qƜlp��]���RS�=5mjTӋZJȅ���ֵ�i.$�x���:�ч����C�!5F��m�}�E�UP��a���H�MQ�z.��r�aޘ�l�ե�Ѫ/f��(��ruݘ�:�L�,��m2mÔ�D�iI�!D>8�`�II�%���@��,��d�O�Zm8�@�R�wꜧ����C2����{�ˇ)�'�!dk�WrTo�i����;�kt'4�`��:���I�^�.ҚL02@�O���I�:�\�.�脃G�t���]8&��h�OĬxa�|O���<O�|Og��ć�Ǚg��<O��Y�N�������ϥ�&��Z��1B+��G�'�_������2�]a՞�Vy�ê��g[ck�q�Y��]q�\a�긮�c���0WM�<W���K��&	�x�x|O����<pu�$'������c����^��������&����O	�bh���h�1�I�y��<L0�~'��x���O��/V��W��X����z�^�m�<>:���d�|:��։���E%��	���r�D��$���$O��B'��.>��L�Q�+�����D�òa:[:v�D�8p|Og��ć�Ǚg�Y6x|C�Y�N����=�ò!d�����^�jέWJ����uRN�	�BY%��%�Ř���e������1}��zB�wP�ܪv���fVL�w�Þ�f{Ӟ��}u՝�;�q5�v�g۸u�ud�o6��^ǜ�x���<��E��m�}�&���k�Yʬj���r�fwk9TW&�
�P��*/�ϵl�����D���}1m��ws�vo<���{g����cri����k)ݪ�o��<n��-痟��d%g����*�E{�ḴKO�'[��?���Ux��X������������U��Z_�����������U��Z_��������w��U��Z[�ۿ׳�i,��,�N��|�6�4�f�V�8/�ˋ��6�������@�u$?
I����7�-�ki��0�����hBC�h�'�R��vD�Qm��6D��x��ì̓�O���!-���!��Գ�̱R~�p�����o� ��>WSN�!D&�6%�2�a�A������5��g�Y_Q�!�`	�p��U'4������/я%���.w�}R��K�	v]�zi�V�$0�!ւȼ:��x�7g0���|�<z񷎸���κ�n8�N6m�i�m�����.�[�5���\�a�����RQSMgC�h1��z��pC n��>ݦ��E'sn��-�D�/��͊8_}��4���Dc��S&J&�x�;��ȝ#����2�HX�$]��Ět�L�(���W�,	:)a�|�9��0�+r�ӭVBl�����fi�.�sH�8N��GX���n��7�����o�$����,�RC�I:Y�Sۜ+�F�*u�Y�'�Kn��ч	�!�ř<xۏ�~|뮶�4�f�V�9��߄#O_Y�K5�ӻ�av^�Fc����%�L˙\墢��$�uίb�����v36w���ϲvG�����Y����vg=��3����^��9�f�o�w\�׳��m�_`��3�OG���޻�!���z��3$��9�Y{2w�w���X�M��W{^^�oW}�ǎZb���7VO3�wm�g~�_z�y�YяF��n[���7uh�&~�"�o�2���>!q:���HS���5$*�Ra�-��gj��W��
l�Rl�'\p��!)�leź���$;\�<n6�oUd!_4f�ԩW^�&#�шx��5��yQ�gҐ��>K3�t���D9���HL��|C���K�10��f k)�Q!�|�G�|�M�o&`f�Y*f�8�&�JN5$�-��Ii�oe�2�0ĉ�	��a��U��m��?>~~i�]m�i�Ͷ�:�O.j��3�`��r��UEUT�E�ӭ���+�-!��B��<�ŵ�tl>���8�BQ	�v����o-�]ݒ�m2|Ӥ�����못/e���rY�c?K�J�~a2���08Jxi4�2CI�4`��#��	�$�5CO���nh��75�c&��޲ke�jI�҆�z�j�$1-4]�}��B�L��
!�:���b�YaB&}�Vv�8���B=z�?2�/_��8�Ӯ�ۮ8Ӎ�!��<n���.�&c�D5����А���B<�WT��cYY���oΜ�H�o�OI#Y�3���-�e���o���ǯl~���s�ʜ7Nh	E��H���zG/���z�fMGX�/!�9]��a��m�r����UZe�Y�C�M���rDd�̫�A�� ����6!o������*���E�e6^��L���XCV+tae�e�e�i���~|���Zu�\u�t�p���{uOٙ7��! �{�QQZ�V��kgy���R��!~��9#��K���sꯏ��n��Q�{��v�ܐ�XWi�sw�rj*�X�gN��U���!d,��������o����.&z������N0,���6d�r0�@}�T��zG�e�ܒ\n���x��Rn.�ӪM:�������>�5D�mt�S
�{>Vf2j5>�==q�|��[|����u�qƜl�j|x��M]�Z|7��ia�a�du�0�c���ÏQQZ�v�7���y����ۅ�ٻRi�^���sR��s�t�_n�^�SΝ/o7�����L��^�۷�}��{>�����9�j�#}Ggw}��w��ߝ&{~��ӑ�X������{5�{lϻ߾�Z�,�e��g��yz��>�n�k�L0�+��އ�����Jt9!���ZsA$�A�KH��0d=԰�
��Жp�2�a�{��J㉙�)���ֿBC�(���aY�Ԣ��Z�sdl�(���f�>-�`�T�f�Dp�6b`��J>��>_	|����O��dx��1nD�q(��!
�#xɇީ��@��&_2�ǯe��ϝ~i�]q�i�Ͷ�:涡�Z����[�V�2^��.�3~�**+BB�X~Ǳ�ߧ��g��]U����C��=�04C��oӮc.29�t^3f��BM���.OrN� i6m�`��e��4��q���[��C���ǃD9����nv�Zϯ{��K����f�`:��uE'i4��������5>>U;2柤��z�Q��m��0ЉӲ��<�*a��ҩ�a㲮����ϋ�>e����_�u�\u�q�m�N�� )���������$BC�;-I.�Uփ����|!`'c���J"z�I�%�J�u�l��̐�ф���|��_�L�8��ZM�N?9`h���Q��˘d�vi.c�RItC��G�2����%	�$��T�L���BM�r��gz�,��S���6�R�꒢Ԓ��&3�#��D��˪d+/_2��Ui�Ǌx�>���r��'��a�^6��>�]u�]q��4��u�o+W���Y��s����I���>�1��Y+�rrm*�(��Ɇ�8��Jv��l�tH�l�t�T���ɹ�6�L��#/"X��vV�u_���4�z�t��٦�ưaVx_��[W�O�~�(��S�����ce�C$1���sVfMئ���+Ʉ���qjӜ����}l=��<<̄���벳�ӴB��!!F��>�$#���i��L�C);��a�n�d��F�!��&�"N����~������������<'�x|h|O�ǮC����<y��D��ܟ�Z%��t��v[]Z�/K:�{l����Y`�L:���Xu^�Vu������:Ë�Xq^/u�u�\c��u\u�����|�^�����|^�����W^����t����
O�#��0�'��x��x���!���a��c��G��:L��8x�m���G��0x�'��?���xЧ�̍���|x}��:>!���t�I�ك�xO�ÒY��,i�f\�xI@�\D�^�O��\}��z�/U��gWK�O��u^�1�a<_�>/��8pd�0��x��<>4>'����'���^<Ώ��[���+�����t��k�Uժ����u]U~b��Y\)�b9�������z���a���]~S�o}��ş�����E�ӱ���WݞXw�p�������r�Ϟ͞�t�~�>^�~ÿY>ՂfD���#*s�j��&.���>�N��m���w'xU�znΝ3-��+��o�z��ݱ���+�{4��B�UΞ2�����;C�{|�3�7�,h����}곙x7,;E��|�L��w�&~w�{3������d��n(��U�ƣ��X�VՊ�s`(�,+`����&{����3�j�U_+K�w��ww{�������W���o�����n��j���U����{�������[Uz����o�65�Xm����m>u֝u�uƚ>>!�Ƌ��Kl�E�mL�1��QF�
��j�mjr)!
��Z�*��T�8"R"��N�-���@+V֘ب�r��a
���I%PM�$�KE���!�%�o���P�tn��\��$�	#����(Ӎ+iD�[�Aȋh�\N�b�
�
�#	+O�F�-��)��Zq��$�
�v�Q�I�bmU ��q�����qI"�,�n�]���QT�Z'X�t�QZ�1NJ*N7#�:Q�kRKcmZ���ll����mDWU�dt�#M����@�mE%�EP�#J���W��h��9Pʪ�WbrX��(F�*�*P��	aX-�Ik���*+�;JYbb���Q�7�� *2�+-�إ��F[a-�8D7,Bq2� ��m���ډ�F�T-d��Yy#iDB&;�8Y�bT��X�UL�t$t ��mUʬE�T�#r�lB�H.0rȫy	�`G`��>8�V��dEL䩜t)6X�w��+�*n��
2 TU�ҍDYA�ǝ�6�m6���ۿ�����F�/rw1���v��S�[�w��S�c���]6�˽��>�[�>�-���f���^w��W3�w��3?f��E��U�gW�]��R�_-��깥z�W������]gsMՒ��U��4�:��I	P�<��=2��	+6C86�2ਕ2C�&$���Q������F�)U��_OĜ���Q�HOÜߤ��s��y�s8��G�Of��l�����OrO'���F�"5��Uq�M�C���]|�r8!�V~tQ���a��!�w��C����r̼n�&"�"Cu�?I�_=���ٜ=����f�pq!�f#G����<i���_�u�\x����������8��k�~���k2�fK��i�(ن�|����$:V�/�s����xUY���s�W��5�C�w���UE�4kć�.��3F�Nd!N�Ya�ݖ�]���2y�찢��l����t�1o=�K��C�^�^~������[5���kXe:��e͞�d<��OvCʥ��,ma�?q\Y�����X���T!��^:4j1	���]�m[۫;y��O_��0ʸ񧎼q�ϟ�i�]q�\i�M+�\��ڻ��Dn�^���!|�J���1�[�����4|`3*zRu��m-�;	��t{L+�{1��5&c+<F+}r�������7Mɳ.db �MLǵ.����Vk�*��4x��y�o����Jݫq7�W�b>�esOF�����f�KKӖ�>���Zg�u��s3V���u��L���q�˺�������W/cz{4�z�|a�z���玶���:�<x���||Cg�Zd�1�m�$$�(d�Hci��TTV���
�p�J&���"Xl�U���p߈�*���v&�
mMڞLXeX���o8e��8���o���t�46���fYS
�)��{F�/�����jv}�w\杜U��uR�'��c��	h������:�U+�ɝ���6�Zda
�����V]\�,�Ќ����[L��瑆��<��Z<~W��>xۏ�?:Ӯ�㮸�F�Wξ�L�6���I�׫L�E���웉�I�1㡩%��s��TTV���s�oZ��rf�z�뻡�����ϩ��+��g�3s]q�/�j�s;�}����Qy_�f�ǟ�a;?]{-Y�c���qTB4�qI��e��_�Z�K\��7fA���w5�ߌ;�Y��_��׋��.fa3̄Q��6��2��2mEr0�q����^3�6�k���]��'�S����R��O��7�;��|{U�uum�4O��W,,���)vX�����Z����ڜl�Z�b2�ήW�$�;�?2݊F�O�|��l��H�F@�A��aH�TEd]&S}N$��<�0<C��8��Ϝ~i�]q�\i�M+�X�ȉ��$���3:m��e�`l˫,4B�$�	���Q��N����I뺲���d��ʹ��q6C��]�F����e���eIY�n�'J��L�&�Q[	g��u0!�ƨJ�fk3Ψ�gZ��6*��
��n @�\��+ȹm�֟�<`�ƂZa!��o�;4a����*����Hc�>MG���/L4�<z�׎?=~i��_��~?�00���!\.�l�8��"fB��w�"���$=�����V�EIx�
��:����?&0{		5�2��Y,��G}p���4Cx�^O��3���T��� ����331�f\��hj������᳀&��_qw���c[���
˷`��2gp�w�h�4C���G�%��s�H�L�p��+��!�xYfU��{�M�m��=M��}<�g�?[V\Rն\_e��ͷ��U�fW�<|���t�Ӯ�㮸�F�W�.O1��A�ˑ�\�̴TTV����Oa��6����烢,9�$0!z�/o�d��15��j��|��v�����͏��X�Fb2���x�u޳�S�7��V<�����X]�������!�Eￇl[�?k�Bɂ�5KD4Y{Ƀ,B�2I!�}����mO5&�4㑶�����̿+�2���:�O��u�D�~0��������$�9�0��j�#$�\&�_��**+BC�������l�qa1�����/�/~���ִ>��F�9E߹ɞ�=�M����Zї\�5���B��ݬ̪�5s����ǣ}��N{Ow�Υ�X���"�1_d�DI�o\�sn��\�ӥIX%һ��Zc��-M�Cw�S&�P�,����<����Rs$��$!�K0����0�Y
|��1����G�&6O���;Bo;?��K,�'.qz�z�s��K�/��k?Y�'X�!�RBt�����y)�pk�|Io�dy1�.zʜ�Y�'�HB���k;��"�������C���9�	���)8��*s�ב�2���Q�0�b��z��~a�l�q�?4�֝u�u����>gM�7�P^%7(�� �i������lXk[�EEEhH`M�Č�zJ!��=p�|�n���.��v��oƨ6_w����f/7�ۜg+:�Ƙ���X�4�K��y�\b�T���~��Q��<]��Q)5V�sC�'r�V�(p��j�x 6ԍ�#�r�ҝ�! �M���	8Ru>bgi

���
W=�q�m�̛�b9�_6��ƞ6�YSA�"&�pHA�b"xD���!Ӆ �!b"%t�"pN�<'��Hh�&��h�&��h�&�i�M8"'�"&�P&�E	��D�dӇDN���pÄ!�%���"pA�'DD�0�4O2i�:p��q%	�(��#'�'8~p���.��u�m�^��l�ۮ8ۮ�˧]W\q���4DD��� �	Çq�VS�:����y�������a��<tS��2�|����ea�%Tͮ�$u鳜��飒�1���L��?w.�a؟����w���7���;d.�z=�}�>�o�)�e�Ӯ��gI������7��w�.y�_�=�ܝ^s[��@��~�}���{�$׻��ׯ5�g_�r�0N���r��92M�N���Hy�[�����}11��{����xbܼ]���;3��d���I�ow�5�~�~�|��ew�W���j�Ux���������~�j�Ux���������~��V�[����[���������[Un��w�l�6���l�m�m���Zu�\u�>>!�:<��%�h���	�wg���s,s2g�>9^C�eT�V�I�I׉O4�!�V^�ƒm�$�M�č�5�Ϋ\��p�8!���u�xƮ�.�sX�F\I1�L�:�~C�}�2'��m��LF�vV8y.��U�xލܑ�[ �&=�����h���$�M�Hl�*�N
2B�m�/[x��>~i�]q�\i���M�7�J�a|�2�_J�\��/|�**+BC�e��v� ¡���?bI8g��y�&�$=�	��I	9f���q,0B�#^�&��VL�t�_z����ׇrD=I~��Ht��$�L�8�Zu�f]d�a�1i��nF�dpC<7���<��;B@���e�[Z?�}G���'6`4CN9K��-8��!$&�.(8C����C�m,!�0���Ӿ���<6�4Qp�fO8x�O�i�]q�\i���8��ܾ���z���"̈́��tiطs8��ˑmD��Qr�����i��i��в�o���߲���=vY��5g���y!���=o{�F<�:�^����c��{��9�����z��ƪ��˿O�ݾ��|�JX{�{�i�^�>�[�l]��͍4g�w˹�s���7�������1�}��ә}��K�Ә%��.5.�k�??(�h�V�PY�YKpZww�x�I�CbC䅦��!!��n�D]��Vy$$ܚba�OeQ���!�|�o{-��␽�g�~KT�*�!&G\2:>s�S��l�����i0[�b�Q%J2y�Ya�a��˫�4�G�8�b�L%nTk��FY�$�~�#�ӑ�,�rY�L��4�ZW�6�/_<~~u��u�\u�i�i�g�pNK^H���Q/S�TT�����v
�"��:qp�3ZB'.HˆfP����i��bx���Ҍ�:�O�m:x�Q�>M�넖`��&O��-�	��n9�zo�0>8�f�	!W��U�K��M���L�f�4�Ԏi����ݚ�?vK�D�~;ų�r�p�wܒ]�a)�ಚK.��6�d"���aK\��&w���U�����i��<q�֝i�]u�]q��V�}�}�g>��1}��M�!�S��f�QQZ���E?y4��F�!ԣfNl�O~G�;y�p92�(!�0a�y6�(�U�@�e�~�%��g����mgDɼd��bII�NrTϰ�4�4��f2�/��[eLry�>@��tCϏ3xC'�:j�������v�O�r��4�+��j�G��u��M���x�׬�|�i֚u�\u�6l��4l�A	��j/n�n28!~�QQZTktl�]���Cv�t��j[�V�x�e��Ry4�����L�*_���|�^a���˙�s�&Si�$4����>�f��9u�*�t<�4�:d���:)�˼����~y�&�=�'�ʅU�2�N�0hِ��-2Y���R�z�F�|��Ofv�F�����<n2xʸ�O�z�����N�t����f͐�F���K��Z�8�����g J���qgݍ5��}���&����ִ��O����;�mTi�竧w����[��{�={W|�����VrJ�7�n�K��b�{��9j�U}��[�uQ��k��m��ީ~6d7�Λߢ<���;��H���Bl9�3���gl�c)M�_z�_Z�9W�}�Q�z\r�+����[XZ���ԏ ��z��a(�����Oq�M��:��|�{�!��<u�e�DzƘ�i������m�a��ݹ�����̐��Q��8j�0���,}Z�XX5u��H��F�M/I��LC!�J`�f�a�C��u��yz������;F����`h�!Z�������Î��玸�OϚu�\u�i�i����3���yX��Ȩ��	*Q��U&UQ��|BY���ܒ;��s1$�m=����»&���M%�~Ļ�����4�N�l���z���]�6�O$qE_dVr��T�_�����Y�2���6�Cź-S��8���(�YÆR$f�^�J�76� h���zndd
>ˣa���ר�we:L�h��x�p��x�o�u���i��N�x���O���|&Ƶ����IzVp���EEEhL�:f��'�.�p�4wD��7�xNq6ノ4<v'��f��$��	FS���,�%�C]Es��r��{;Da�����|u�Yn���P�5�'Sg�ITW1�C|M�-9R��S���|GUH:��J>m��zl�,_���Ia%�j�>g**�>�?HE"��ǩjk9�� Z��%ը^Xi�_>x��:��]u�]q��WSZ�_��`^���r9�%�l�z􊊊�׋����U��z��G"�x3�0���X>K.,?	 o��LZ�Y�M��ݯx`Z�f�u|������&�����8||(�~<��t1���cRi���s�ۺ��Lvx��+��A[���ك������F�U��"��S*L:���i7��HL�
2�ї!��Ǔ�ѳ)�ّ��q�k��:�����?<x�*����4L(A�b"xA4DD��:'N � ��8pD��:"xO	�`��&�&��`�""p��!�%�"&�pO�D����b"`���DK:N��<p���4D�L8!��bxO���xN��!g��Q�8FO�A4p�\u׎���]|��[a���M4델�u�u�^:믝~4DD��>�8P� �t:x!�O��r��5��t���om������/}��3}wvh�����{���Z���3���jĠ��/ۺdS�ȝ��[��޵��Vt�擓2���vk���>�,���+�y ���F4����زM�|����ŝ��_������{wwW~���y�}�b��̭���M�d�w�)��iʼ��n���߈��z^�%Ư�N��Ͻ�o�����콮osqV}��o]^O�y��f��҇V�{��{��b����tm���ܧ�����g덯���]�x�\j7_�e���i2mX��s�3/�QTmo;�o}�W���[Un��w�n�����Ԫ�U�V���V����~�J��^*�ww�������ߩU_+�V���~���4�M8i��4�i��:�:�4Ҵ��c]�����[���c�[+��H��9C%�����䶤���K$���$�q�+R8q����KKx)G+q6�5#��[l��l$�Ȭ��]h$���A��Z��C�������lCN�m��E%b�A	�Wk+9 Q��p��;�U�9*�q΋j������v��-d����\m�-��q�۩�8�TD�]U���Z��brY!�	d-h�u��n��Dƛn�j�����RÖT:�Tr�Y-"cTA
��\-nNZ���8�:�
�IJ7++D��I�A�\�����"��(B���$ڣ���j+e�&��IcpC���K]��%�Dm(��y$���C�4�7c�(�����FUDR�v&�,9T��,qF�d\q�ؚUZd�:�2��y*
&���ܮnI!*�,R�ƣ�����ʥ�4ڒA�q�lq�8ՔN��Uu�cv�c�\d.]"Y��3H�
�l��R�\aqIj��B*�PR�Q�ePW��WF�VQL��/ �:��5��9.��~�������8���(��mSTs{��~���^]�1�;4���h�~i�~�|�J��<�	Ozay�}rcϓ�s3��X������׸��9������s՞���j�S��ҭ��k����������������e���5CU��t]�|�9���RO��lh�=Iﾊ�����M�:~�nI�z7���'(k(٫���$�,n��FpvG�U����ÜB���a�Cl"b�v��̶m�e,;�K�w;����E�{\�*)kˑ��ۋ]��dM�v�mf�����p��!���K.����[��F��}�/U�4���?8ӯ�ݽu�]q�M+L>q�ۆ����1v�ܬ&�j�XE#�e��<���0���f��Q*��D���ӹ2w����C������Y��f�������-[��PupHת�P�OZorω.��87�M��0!�Ĝ��f��N<�v��̥ѽ�������\���o��oN&u�����Rݘ��h2ps�\_�;%ԓ�Q��z�C��r��>9�,����HGnS���(��0d���i�Z~u��u�]q��V�|�ԶnW�^��\�\̻1�x���2�'�_/��'�'�8sX�
(��ɗA
Ą������ـ)�����dN:�`�g�9.L]�u��Fn^�m��%��<x�+GL���OɃ!�L���8m�/��}&��v�&L�C	�&��C��Ʈ�KYkn�߬��6v�⬰��a�ñcZ���x�֙i��8�OζӮ��4�J��f����[
�uQQQZܩI(���oK<�J`p���N��4K���Ie�o�[&4�'m7-����NQ%i;�NNU!Q$d+�j�#G�����	�h��2`����6��l�3q-)�`�XS�Mk5W��bn�Y��)?h,�w�j#
������ƙ��`ڡ��Ν����1!1�%#�l���82S�:�pq/ ��`���A��`�e�_4ۍ?:�N�㮸�m+I�_n�_|�]Y��r����Js)����ja/���EEEhO���nY�ߏ�_}�:�����0�ɳ�6�ۘg�_�0����,���xx�����,�ݚ�ߚ����|g_~߼Y��or�ҝ�X�7���VE���^L�s�H̗����}.�����~�ד|���0Ӊ�^��3���9�;������=�o�r�}�_�{}ݲu�����u~���.��r�0�����v�{�':��4e�V[.$�����v��V9_rN�Av�2�p�A�F�f�%>�H�1����'Xِ�`:����|Wط*i��̌>�ݿ~�z���~�4���;�f��àsromj�6�Ϩ�>��I$������drjaߖ�4ч��:��_?8�N�ۭ�㮸�m�L>c���GDB)#|J[9G�綴�������A�x�!>z��_���>�*��|�w��aG>��w~���x��~�'�>4A�fM��V���)�]7�����⏈w�Q�cC�%�����|�2�%�9�����3.�Nh�Lŭ׫�N?fGf�$M�#��^ԑ���)���L�xi4=�v��[�5>��\��r7&�=WXi�_2�M�Ӯ��N��4�j��M�S� �.��TTV��_r��E(������RU`,��i��(2aG��Kԁ0c��x��Oa0kē�����&,��J�Q�6@�Hg�<WЂ�%n��Q���YP���ŎF�����<SlE�}���{df��ɕ��,2�l��-�A�X�ѻ�a�����'߲{2F��٭V�4i:���N)��-h����i��e�]i��u�Zu�]q���.��n�DR ���Q"�T���EEhOU�����������6eoq�/����&��P��s1�.Gq�*
,S��uy!n�6,�䐄;.v2�P�Zd8e4q�2v��cR��%�>v��&]+5�i��.%��p͟V����e;YR[�2GI��ND�s�<�4�<�����k���fC%�FM|Y柝i�[u�\u�m�i��k�w),]���EQ J���ݖ[@$�Qdh���Y���k�h���l�.�'�s��1���}��_vu�L��MÄ�s��Q�]N��㝹ǅ��7���ggw�ݟNIݹ&�U�$�2H�n\ʻ}��z����|��j�����Ǿ����fl[�	�{�֓%��fCFRu%�1�&݅&'�G5�϶64h4Pː��1$�,�i�i5�zn��|0�H���&�8H:��t<є�CK����c��x	�ny<��rً,�iU����w�W�(ü����D��'#�3۸J�+M�<W�<q��~i�~u�]m�ǎ�8C�l�����u�r(��L�+%µ+0YZ����**+Ba�׏cOY>c'\_|��6�qxj���Yup�ߛo.cvL�*�O��ڸU���Y+ݥ���F0�i�-Z�O������5o�vy���5:�=}˓N�^�?n�FA�H��1����$���2�ZZzT>
<�Ō`�e2�(,쐓���Kv�6Ƀ��#ܹ4�E�a�x�K,��h�DKD ��"'�M�a�<'Nx� � �i�p�Â'����xL4MD�4MD�L<t�,���"a��!�8"tDL4O	bX�tN�� ��"";"aB�D�:'���k'���:!g9�(J�%���A�q�����]i׎��i�M4놉�"A,DO	��'����m�]a��Ç8p�t����'M�5gd=5���2�(�iz�����>a�;?1o����uy�>�Ns�:��D�������}���e�{��[̋�5���W�kK�gqzw��{�3���}bY��~�E��}������oߗ[W��>�F\���P^?���m���ƽ�;�3�0�׫�}�7��6P�W}?fm�����*���_������/誯��ww�M������*��x������wwww��������������������-*�wv�64���l��m6�N�ۮ�㮸�m�blw\֑QQZ9��v�����4a�Nm->t���zp�#�)��$~�&(��냉��iӺ&SS�����*ϫ^��4є||���ۍ��m���!� �0���C	��i0�4���`�I'��?<//�[�p��=�B�u�y4�a�_:U[wk$$�	ߎ�~����ڮQ깿cؾ��>��M��-�ۭ?:p��㧏>8p�rf�}7$)�� ���r�M� �������П�I(����А<\�d"O.��϶����uYr]8^����6�ŜRʄ��Yɐ;��i�}�Fͤ2jz�Y_\���D���+)	��O�ఁ��`�Era۠�WxUUQUU^��)=�Ķ�Ͼ"dr���V�4����$�i�i�Z�d���2����o�?:ۮ�㮸�m���F����G��ξ;t|�7u�j**+C�Lt#����~�����R����4������ܹ�O�o�헷��7Ҿ����w�Y�]�Də��ҭߢ��ݳ;}���X0��Vt�Eq����ӯ�V��Xu����ƚ�Y�d�{��6���\��z�1����X�B|m��{g�o4Qi�Y��U$$�d6��"C΍�$ˠ�|zP�z�N�J}��=v�ݹī����Fc&��X���V�#���FQ�I�.]�d��̓G!'MWRx�*���~�ʒ]By�뎯#z�5��9�*P	�fGA��g�uu&��D�$f2����!�Z���p����m�Zq�\i�ն>��j��cSѫ�h�cD�y�**+C�$���a��ra��L�-���u)���2\��̙�B�R^_�0t�·�fL9{��'����+�gd��IG�I�˕�*x�]�L�\�{�3'#���m��e{��ջ���1C�*����/Ԛ<�1d�zk����5�{��T��y�g����̫�[�[e��~i�N<|t�����I�����̂�G��**+G9��"���lô�SrH�`���&�c�~L4ٟ\��r<�=��c��Ϲ�`�.���U�2�&S㾒�O�>u��|LL��T��FSi��<Ѧ:��t���n��fU�����2�Wn���!�Yi�Y�ĒIz'������2����̿2Ӎ����N<x��Ä8;���}��UKkW3=��QQZ;r�Q(�{�FT�u�2�Ot2����餴�,;��R�_޾\��>ꏲv�N��t���N�۪��,�U���J�3Hi���fSaC��"Ț��y��}Ne��F���m�&1��Y$���N:gKG�[��~;�<��nܦ�MXa��GM%�Է�������d:W��f�<m�柝m�Zq�\i�ն>��Z�L�mx��n���9��Z�*J�m3W�Tur��ol��������]=��;.�����M��s'��9o{����W&�.�+s+��}st���B�[rva�M��w��N�3�o5���i�wF��������&�-�5F{Ӱ���<�j��1ϳ�s�3b�w��n��͔e��9{��<�߲���w���a���~%lwp��RAc�~�|����V�z°Y�$ۃ�=%Q�8��R���֌8C���%r6�5���w��)U�v�V��Z��*W�?|�+���`�t-0���E�,)�_hj�yHwRl)<-� Pj�>���I�q��Ҹ�2�s���B8��A�wd�&Z�������>,�-6ۍ:�n�ӎ��M�����t<�-���\�z���(�ai�'^�u��Ð5�UUt���?=&�V'��f��Q�?a�ʤ�T9�5��'qe�i8�n��̆H�M��O�j+	��~����/���o��Hݶkl��j������GM�&���>�U��n��}�~�tvd��e��%	a��4�˾�6a�c�~e�]~qƟ�m�\i��������U��&��ɦe�fe8��z�;��EEEhtQ�ueK.�d�I�&��F��|��-�fS�C"p�r9�R�%h8��9��x�/�p���/�[2;cݺ]�̊���o9�@�?�>J��&B������v� e�a��� �M�����Ǝ�`jW���JJ?��K���e�g�zL�owWng3��W����PZ�)�<M��Z&�:a��i�[u�u�m�m���:�Kt\���%�˒��"���~0e8�7���&g#O�'���s:��R�U��F`Wq;����?G�w'rI�H:L���������;Ni0��I$�q�n.&����7���7�Ĳ!��I}&j뵠44h6Q�'$Q�%|l3r2I���_L�|>5�N^�����'�����O�d?�� ���D�B�DK0M<tM<'�(�A� �	�(��,�'DO	�0LH&�"h�&��h���	�J|D�K:"""aB�G(�b"xD�DD�<%�bX�x�,����dDD�<P�$�A<"h�'��%��p���(��FO�A<"P�	�����8P�i�L?��"A,DD�4DE֟:��̰��:t�Ç�����m>�$ZW�������{�����d����x��������o�~�'���wz�|�w��˒{T�욇�����|�c�g6��m�?kta����Ɖ;�O�mlǇ��w���u���{>�<�^���C���ߋ�ߦ';zw_�[��v����nj3�i�Ω�ȳ�3V_�ߵn���Gޛ7x���.����N|�6���ū��������.bm(m���}���.�gG$�w���gC16�󳹾9���۹w�X��Y���0)�Q�uD�V!�*��غ��ý������������𪫋J��ݿ�n��������������������UqiU���񻻻���*���V����ψi4�,�O�Ӯ��4�4�j��_�����s�.�<2�Uee��Rt��v��c�5��dS�!�EQ-n�+�8�"u�\�vRH5'�am�Wkh��*�N�2��A�24�Q7KQ	��2i�Ɏ���VZ�d�[H�*W%��$eH�"��m�nN*J�h��(
��E A�8Y#p�:�bd$�,��Z��a%���*��*���s�䰶�ER�l(�i��d�RGr**�d�^>Y��nJ�F&�\v�'"p��T�`pNQV�KF�[�aqJZ�PT�!\��#��"L��Z��"q��[�8�m��'���T�U-Etv�v2D�A�@R�x�pV�e,����H;c��S�5X��ISj�;-N'#C���Em^T脭�*��:ܲP�<�\nX�T���X�X
�[,���akL
7Ʋ�U�%JVQ�J��V�v78�b8��p�P�(
8�r��V�@a(�`�v�V����Q>TՂY\��T�˘���dK��"���X��l����g�n��n�r'婻;۰ɽ7'{^���WƎw����+��3�����o�[��ug���f�V?g~�=��6Y������]��]k���M��j2��}�;��"y��n��U{�{�ɯ�'Z��N��b˳J�GyR�w���h��׉ׯ6N%h�Zb�.L�ߧ�Y��mǇ��[m�9��]Uag��7E<�nHm�n\��<tѝ���$u��������6tɧy�Ok���s�.d���%?qt��2���..L'Jgd���~�E+o�q�6��?:ۮ�Ӯ��k�^Z���9͍���8��ŕ�f9�YL��sSR�!"m-��~�����l4Ւ�p�^�ў��~��|�U��T��<���#�x_-��kK��Ʈ���e�P|'b����~�ENN�J�xs0fb��p���f�d��$~u����G�r=Ŵ�}^-�ح��[��V�n������I�cCG,5\�@�CO�q�^?8����[u�i�m�8|Y���� ��0����a!!%�����̵��s��~�<xng3�Ua��QԎ�0!�i�*�U�ОN<�$`u��fv�g���$��W�.�����Պ���|�����dR���%|�S�Ce,�4`m������bn����Y�uX�jS�E�M/v&�lNY>~Lr� �h¾x�L����_?:�n�㯝q���b2�i�c�LƵz,�ie�9�HHH���ɣ/�(>�$�������8�OA�e�O��^���ܖf��k0���3eU�g�
�u�&�'OrY���h<3Ed->^�j�~�ӏ0�ץo�w���UeߓO���R��|CwEդ:�`5$��
c�ƒ���f�C�ۄ�xm��2c��I�ն�m��6���]u�]q���a�����U<�e����^�ܞ�\�*��!N�� @��;�����ו��$�rn���u޻�>�=7������a�C*��vg��=�o�}�Ίʌ�A}s^��;�óL5L�s��]�]���Nu�Y$����}{�}&����ŉ⭖�7񙑆����Θ���H�&���[�w>�ufzK!9Wx�10I��_y,�e�ө����=Uy��Ԫ�u/F�ZXD�C�'�ɔ�zb@량�U(�7|��9��i
8e�UUT������i��1�j�ǳ��̗��\ŝh�<�:�'
�?W(�00���������uJL�
溦��� ���ޥ��np�m����i��Z����z¾u��_<m��κ�n�㯝&i0�ў!���9;ڹuT1��Z�ln0�)j6�OWՇ�~�t>�?X����@g�;��T�Sɜ�r����9�hw���a>'�����?}����>�vÓ={�v<0�2d�4vN���ꡬkEq�h��I	����v��I�?p�B9�:�g�	�!��uwu�ZN������h���Əu�]q�θ�m�m2��q{c�<�hVҦVV�/_��!S{��$��fOh��u(��&�.��a��1�F3$�&�/}ۗUww&$�K&���N$��蒃Y�5Y>��G-ptl���4�&,f)��]WKN�v��j�i��˗�R�;�FL�Xh4������çdή��{�S��.�fQ�?l:�Y��p��&8�0d��,�o�8㏝u��u�_:�M����{���%�K�z�!SU��3S5u��p��LӠ��	�����'q��~Ǚٵ�/{��3��i�WVw�|_���x9��J��VlrtT����9$��>̘+Bh-��M{�Ҫ�28�{ia�ɩ��.�u.b��<vHH��m�i$�j���T'��PF�6A�5).I��c���!�U֋=x�^2�.<u�_:뭺뎾u��p���k"&L%\�1�ӱ�Yb�1���9� ��𻽭��NH׮�wM�0W�꽞�b��I��j�����u��aυ]l��d7/eY���O�[]��y��sٰ�g׳��ݧ�/[揤�L�s֯����~������#���Sۧ��Z�]�b����z����>3�2gZ���y�K�0`�����̦L�vu:��ܯ2_�	�s�Q��v,���l��;/k��1��"�5�ڕY&��k�!�7�<;M:½�Kh�/�B=�77�I��Hh��+@��R��E��F���7(}��ϴ%��V'���+�Yu�?8���]m�\<l���p���7��&�%�X�����jձ�1.*�N���-W���*����ǌ��-�s$0�@���d+�	��6�9�rŶ�%�.�epq�D˴�ܞx��#!��!���lbĴ�X�q���+f�����7F�e�6|h�Ŝ�� ���D�B�B"tD�DM��Ŝ8 �� �$:'����B'DL̘i�h�pMD�&��"&�&(D����4�"A���J4DL�X�%�d��@�"'DDM�"5"#�GdM�Ĳ9	BpJ �FO�A<"P���A��8'�M4񦟏Ɖ��D艂-��n4�Ǯ=u�.�t�ӧN���x�<'��9��Y/���7���{������f��{���K��k��è�������.�W(���}��U�ﻂ��\��s>خߵ���5y�W�_]����{�	]��Y��Oۉ�͛��+ۆU��.�ٜ2_�̲j�Y��;�OD��t���_}~�4�31�jeM�M鞫n���뫽���}ۼ:�}\+}����TV�K�~oYqJ�?�ﾝ��B�se��fu>���.n_�ۦ;���)çoW�������v_Yn��o���^�ٚ����Un���n���������U����www~�*���V����l����߿
�����ݿ�4�i�NY���:㭺뎽uƛm[i�X��Z������[!�D�ټ��l>����n�{��e�h�;��W(\���:m����~�?g�N{z�w���M|\S	�Q�7���'y��q{���L4���t����ܵ������E���>�l̐�M'�:�u0p8�Md�M~��1Z��t�I2�t��5�D���=އ!g�6Y�Ǐ<㭺뎽uƛm[i�Z��+�t�]Ck�TT���^���=Y���t�Ĺ�;�$��$��o+��e�h�Y2�Š��
�ϗݞ6�O�Nc�W�=��d�;��px�v>N�6���C5:UGn��Hn��(�k�g=u��tt>:l�Z���N����8B�ˋ���q��a���y�V^2�-<i�:㭺뎽uƛm[i�s>��y�gT�0��ϥ0F���=�� �?�'���֑��]��a����\���=�{�p��K�9�^�n���C�,��o��7ӽ���1�����s���÷�v֪�mM`�f<���k֎�Z��dS�xn�!�n�m��4���fd<��}�u��o{+��~��dɆY��d��l�I�ko��7浪4�#�-�M>�N��V`�-����y��f�<��r�rIur]�P���c��BBy�
J4�4�=��˗W���Po0�Of�9a��ҫ}�߱�Ũ������w:�5�����u���w|`�Y�0��.��|��2aZm�̸���:㭺뎺�O�!��˟P��{��^��4e�:���}� %��8�|�m	�Z;_���Ǻ������}�(h����x~�i����~'��Bb���>m��.����*�`�ٸ�BCI��h��'��W��}ո{�v��V)#��y9��#W��`۔�M&�9zi8�}'�F�i~�|ND�}�1�=�ҥN�AK���㛱����_2���~|�8�:�Zm�m�_OUY�3Zն�W�d����-���5�[vQ�R���l�7Dx�&������,�I���WV��x���{�&阍��W�K�k{�x�}��i���MzHJ(��M��ew�o�N|h��*y��T�Hߤ�۫��,�<q�$�M7�Jʺ���|��\|�8�:�Zm�m�Y[���gח�YbiY�f\w "���T�{įT�r� 	�/sx�]G�Y��mL��+�$��*�qw���N�P����$M�O�W74MOL�Ě��j �V����I$��h
|�q&�*Rx���ۻ�(��d�^��:�:|��*Iƃ��[����,�Ӓd�
��Q�`�a��2�IE�WX@�-6�r=d��x��l�x�󏟜i�q~^�yu�T^]A��$@���H&��X-��k5���=� )3��?-���Ͷ�=գ��#o��=g	^��~�t�t�wk�#�.�Tr/��"�����	��﻽^�<��uy!Y�~<���>/��VM�N��3�~��w��9��ї���{	帰X��o٤�S�/�ޯٱ9l9���X�Y�fd���D��(D�O�M%�L�L�69*ț���U�ӣ\Z ��$�*�g~��q������O-p�Lbp�z�2�&��KQ�N��6a�c�8�,YŢ�s�&�����*�O��Ss���z�rh{Ϥ�nB!���Ou�θӎ:㭺񶕧�(��p�L��j � n4?L;m>6醓:�Ux>L��;�UUJ�Q9xԕXtF:��>>~Kvl�����9�,ވI	�ᬦ�;M��9���iƴt?T6!�UTv>/�k�'6�����;}W��|�i���d���J�a�Hȧ��&ׅ+��~eǎ6���Ɯq�m׍��ժ,���[����d�T4L]{����qAC�fvj�� {�~Ydcww�we��D�T��W(�Z[1Jao�={N?un�M�ͫ!6�H�0������K��sb8��3Z�fc��>L}$ۂ�=tgF|��%z����e�;�Z�W�BUg�Zm�����!6��Bw)=Ǧ	����G�ɓ	�0CG��e׍���\sv��m׍��5D4�'8��@|0 �k��4�q�\�>�M�*�jQ�G�>��W����̎M^�Y�0WZ8�zx�/��S8/�O�Yz��#�)L����d�I�H�ͦN%���Q=�ԅ]܄�~zb�8�/�u�q0�}�s[L�2��/ãg����*~��d�կ�O�T%!�  @
(������_�8`��	?������Q� @v�29���o2���s�DaP�DUB����1)e,�������*��&,��eYUVJ�����K
��K*�QUV��R��YRUYUVR�UYUVT�K�b�UU�U%�YUVURʪ�Bʪ�UVU�b���b����*��R�T���UYUV*��B�,���K*YR�X�*�UU��YU*�UUIb��U*ʪ�UUJ�RT�d�*�Ub��UT�J���T�UUb���T�*���UVU*�IUUd��Ub�UV*JU�UUEUUYUVKQ0��*��b���U*KJ�UU��YV*�T�,UU����Ud�U��Ib��U*�UV*�b�RTU*�VJ��UU��V*JU����Ud�%R�U*KJ�T�*�T�J�RR�U*�VJ��U*�VJ����J�UER�U*K%UY*�T�UeUX�*&"�U�b��UU����V*�b�����BʖR��*�����U�����U���X�U���UVUU��ʪ�����*��UIeR�R�R���%UIb�V*�b�VU*�VT��UeR�UUJ���T�����9�FUeU,�*�eIUeUYUVU*�R�T��J��KJ�URYUVUR�,��(UYUVUU�eR�P�T��J��K%U��T��)UeUIeUYJ�*��UIeU(�eKBʖ(�db�bRʲ�(YR�K�P�Ke,R�*�UX��UX�b������(QR�X�b�b�)b�)U%�X����)b���R�,R�,���*0�,��,�YH�������#0lP���YUV)e���R�R�X��YK,�����R�,���P�JU����9���IR)*�
J%%��RP��������H���H����D����"��g4��RTJO��#�RX��%�RRJK��(�gL����*��5#E%�)()*IIa),�RXE%�RP���i��DRTE%�RT%%���$RTJJ�),
0�bAIAIa)*%%AIE%���%%I),IF�RXJJ%%��RX��Ĕ�$��)*
IR)(��$��RY
K��IIdJK	II)%�)*
K ������HRX�II�E%$RJ������K")(JK$�K	),���P`,T`1@��`J�%�RX�%�)*"��)%!aP���XE�E�(�
,B�QR(�IE�E���E��$QP��T�,%�+Z%�(�T(�%(�J,EB��EH�*X*X��
�B���a(�H1��T� �1RD� �H0R$�
�IR�J�E0�*UK)R��ĕ"�,�J�*UK%J�U,T�H��T��U,�*�T�T��T�T�R�Y*UJ�b�T�R�E��T��T�J�eJT�R�ET�T��T��Ib�A�!!b���a�X�Tb���J�R�R�U�0H0�X)0�1 Ń1`�X)0 ăH1`��H1jET�T�T�K)R�JT�R�H�RĩJ�*R�� Ń�(b�HA�,�b���b���R�b���`A�,bAHbA�,�a,A�AH0a0a$A��b���U,�J�*R���R�K&Tb�X�����IeH��T��T�K*��*��"�K)R¥��K)T��H��K)T��K)T��H�J��U,R�*�JU,��Qb���R�)T���Y)e)J)T����U�K(��YI-*�R�e*�QJU"�,R�eK)JX�
0�R�JR�)JX�)b���ER�U,��,�R�U"�*�R�eK)JE�K�,�Qd�X��X�)e*�YH�YJ���,Qe*�e*���RZIe%�K)%����(�)e(�E�7�(�E�K�X�X��E�X���),Qe$�E�KX�X��)T��(�D�Ib���,Q,RX��RKQIb�)%��Qe%���K(���I,����(YJ��%��R��I,��K),�))T�Ie*�)%�YIe�TX�Qe,��U"�K(���I�&��RYD�U)Ie%�.p�bRYE�YD��K),��,��YE��P�YJ���(�)e,�*ʖ(YK)e,��(fa0YK)Ue*T�eK*E����eV���;�l���k�b��JP�(O���~S�1EE�@QPX�VHE3RW����5�'7�w����I���K���(?I�?q�����%����>{��a�,�)C��ᑡ&�����i�_�������������G{�������
d?"���}���U� ��%���?��A�����Q@Q�@�������A�VP?�_���������D?��?�X�)�Z�l���x?3���������!��6���?P��?�G���@�W�B���??� ������$-���k��D��������@��ַ�F�~�?����,��)�fB!������F�S ��2�BL�#�@�X8p�H���  � �ш��HB��$��KD�
^�?֡Zf�\�U�����`�d?��������tYDDZ*��KETH%��A�1EX�H��B*�K���M�0~������M~O���{����;���l ���������������?���* R~ր�����[�5�������"w�3���6C�+�?�?����4���?�L����!����?����������?�?H�*���������Y�����O�>�����N����U@��@T �/����_�?�����iE���:{�e�C����$�AJ4��ʑQ˕��$!��x,���Ԁ��))������1��(`sa062���JhOפJМ\���������R�1�^	�#�P��?�����������(����@���"��֟��1�X������߿ �e��場�b�����O�?Ο������'�tg������G�����~Bu0�(
�����R��h"��������fC������}�	���~'���?B� c�3��a>#Đa�IC�s�G �I	&

?�v���Ki��/D����|������k�\7�p7�`hҀ��I���?��a*�O؟������2��1� ~V?����>8�<�8�O�B��YT�s�Ht�����O��O�DP��?���?5�?H�����>8���ИJ���Z]�Z�)?Q������W�!��T!i����������)�c%�