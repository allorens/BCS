BZh91AY&SYt���߀`p���"� ����bK�|      ��@U�e$4�@гDV�A-h PU�`"% �Ƥ�"H(h�F�
Ե���CJ
[���Im�Gv��YfZ5Y6���Z��e`������A�lQj�F�-��L�ګ,�k-�U(�Pi�i3mm�(*h4%*�1�V@@iU�w��[3f"@ѤQkV�؋m����[kZ�f�	4Rl����i�6�%1��-�j�dQm����ْl�6�b�Fڤ[4��m�;�jͭ�ډFx   �z��n�M����������=(2��nn��]��c����ۢ��^�v�u{җ{�����^���h��T�w���z�=_l؛-�Ƭ��w[TU
��  9����B{�޼�Th����=V�S�\�7+�	PU����Um�V�s��*���ٶ���Ǵ�
�j�=�*H{[U'z��:�)���n���a>�*���i�Rk4��T(���k>�  ��|;l�Ol��/]�� '�Y��U��U(�
�o�K�}����>魚4��;��� Rk��=�mU��(o}�>=�T��UO���Mlւ�����믮>���<{�m�+V���V5��i��  �w|�t��[us���}*����|�ǩҴSA�麝b�W[�׳������K�g:�z=.��y��j���v{�㠪z�-��7��{SA�;�z�YkN��zDFբFZ*+FC[mHg� ����i�m���v�QGmA�g��{z����y��y�V��S=�򻴺W����R�T��B�ʕW�=�w�����Z�z�禤)�/oݲ�ܒ;�Ѧ�3Z*���QV�� ϕ��*Yj�Ѵv�֚4���w�+-jm��{m�AC�w=�z*�i���5�{iT�v�Kp�hR������.{9R�mf�7����J��Oz�(��VCc3Y�l�  =�e4ҷ}{<z�T쭶wS�jڕMjq������ݞu%zԲf���[�g��n n^�4��(/y{< =i��w� kV���U$�6��fY�&���   n|�P
��� =-���n����
���{������^ iC����B������^�� kvS��=<��dZ�ͬF�k�J���   ھ
���^�z�� n��T�rw�^�k�w���]����`+n�� k:��� X�3=R����m���XŴ�QB�  �|J�����{������9���9��;� ��ޔ��W������@�h�^�xk�h���V�]>     �  S eJUF 0   !�C�*�  �  1���OUC	�M222` T�U5Tb4�10LM4�2 ����ф�d`#M=CA�!%$�ꩡ=	���##��S'߸���������_�!>R���yל͝�[���FS�+���� � ���?� �fidAT�Ȣ��(�
�����O����~?⨀*��檫���*�X?�����+������?� ���|e�0��?с3	�����eX���}`�T�eYFoY���}`YS���}eOYS�T��}`_X9�}eY���}dYS���/��`OYS���=aOXS���}`O���=aOXS�@��E��}`YS���#� ��>��0z�>�����ʾ�/��`_YFa��XD��}`_X���}eO����"�"����/�+� �/���#�`XG�A��|dYG���}`_X���}dYO�@��s��>�/�� �ʞ���!�e��=dYS���}dXG���}d~��A��=eOX� ��>���z�����~�A��}a_���}dXG�A�����}dXG�������#��}d_� ��>����� �� >�G�E��̯����ʾ�/���(��>�/���>����"��>�/���e=aXG�A�=aYS�T��}`Y>�C�Q��}`Y�*z�>�����xʞ�/���
z�>���dOY� �'�)�zȞ�'���"z��� �ȓzʞ�/���(��/�zʾ�l!����Y�E��}`C��aYA��}`_YG�����/�)̾�����"����/���
�XG���Y��}`_YO�"zȾ����
��U�\�����+�*���+��Y��}a^aC���}`C�P}c�  |`~0��U_� !�
+� +�(+� �a=a}aT}e}`Q}d}`P}eD}d~�YYY���(z�
�Ȩ�"��(�������� ��>���C���}d_YG�U�`C�=e_XeYG�Q��}aXW�E��,��(���/0'���"�`ɑ�"��i�JD͏>L>9O�ȳ������ڶ����ӔY_>�.���x������\q��H��6��R	�ш�w�8�uXx9���AYӚ(�Zh��*A�I6�̻u�����E�k<��9ݷ`�m��5Ju^∽� �����"Nᡱ����k���'�}fg	e7����C�Z��½/بޢr+�).	k7��9Iٷ�K�p�eKӖ��v=�~�7h��9���D��i����[c6j�
���a7�]uP�r9��a��>At{����;܄ۍNvt�i�,�㗐}��U�K���WpI���pʅ�g*�wk-<)d	X��ӹBa�M�ڃ �t�ld[$
>1f����t��=�UI�[lحۊH*Zn��'��H��q�VS�X���CF1[�ਣ:���,+k�lUnɪ�RY+i�K	�kn�؆�.�������1[�Xn�9�S�*J[�8U�������,N��!S�Ӓ7�v�ޚ,`&��m�ZΔ�h05���3��"�k4��ćW�U��X��%��s�.n�uni;�<�7�l��#Ɏ��gi�;�԰7/p�r��3'S]�I���L�r)��������<4��V����<®Kpb��h���2e�yHv��7�e�^߶�1�82��������P����OT�V�+y݃V��K[ܖ�v��B�����p�#.��ۻ9�'�Qx�̓J�g���JI7i���ni3�md���s��@//@���q��ч������:QA�wNV��J/��Y���wFu5���`=����2\r����-�Gc�Y���ִ����c�{��:��v\�����!"F��\jZV�dJF2�#w��e�ُA�sl&l�S��Z�om+� �C�;���e�� {4�@I}U�ŔK2L6tJ#Y����J�5o\좞�4����Y��4��ݙٗVA�!�"���P�wn��{%��� u�ZV��[U��z#M�0BV��n��x��e:�o%V��W����d��ړE�N�Y��L���<�b>��9a�S�P���j��<Q��v|VoJ�ϞwI������-�ÌMYP�q��i�������S5��妯����(���qAT�*
�@�s��i�A���kSȬRZ���bb�1?�j����]l�G`Ꮡ����.��:�{�%� �L׏1ToKݗ�L�&v�b��ؐ�vP�ˀ�/e��p*�Y������� {6(�S�T��V ���=^��5"|����I�W	�h͘"��y�hb�����anK���a(mrvi�B[��~"M������u�1.��,-��U�`/��e[4�P�� e�ZwWSN���Ѯ�h辤���T2�A�Mc��x���Of�8����>O������EOܬ��-ˏz��ɷz�i���rκi����� ���y&��k$�Do�Mk�^�c�&ꃰ�e-��3/lG��m�26*��Ն����;غ�^{;V�{��f�v���q-*�� t-�ß�5�PJ�З�e�Eͼ��c�_l
�y��흢ʜi�By'mqa�`CK�e�M�͛�nlN��������K��:r����iW�Lx�@�Sv��u�֝�c����/&3�����x��`߻k	�f�!Mn��;:]�T�^���X*�[9�7,9�{+!.�J"��#��N;Nȍ9�3s0��i\S��V,3��v3�x�8��RD�v����}�������6L�v���:kqg��K���Ņ���l�jf�)��tѽ���#d!E߰]���5f�4NAs ��`�U�g hƎ虻�耑Q{�-���ۤ�0�6uOe���/һ$��&�fu�����l ���p��jج�qS��pgN�ݰ�����4-2\l '}2�:7i1٣B!GA�����c����>�i-�m`T|-%s�X�Fq��!.�^*�B'\�nll;�	�%�7���NKs�t�C����Y,L"��e����kA�\����pA�cӋ�Nĝ��&niC��U�]�(���ɛ�N��jIi{uj���i�ҾW>1�T%�'�1MӸ�YN�P*Ax�Wl{��Ź�O g���3M�����ga�/ ���U̙i�eV�����Y�ƴv[�6��l�+���U�^ť�[f?��ˌ�f��v��yry�"�ڟ�2��I�B�F��Kn��5���v]!4��SM�]��P��f�b��`��u`<$̌*U��n��%�l����ʯfڦߝ&��7O�a�h��	�B]yN�2֜osod�gI�X.uW�bZK�3a��m�Z��T����Y��r���L�b���U�����g(�5&L&�o6�u�L��nӡ�Z�99S�\HՃ![��̵:�5=F��,H*cy[�;[�\g�Nܹ�e\�*I�^���#p�̨iGn	9�5��:{�P�9-]��B�_�c"E�[Z
����42��*�'l3f󖝣I��xp����,b���^Rz�w9��LՔ�@c������.���L�1>��t��Bc����,���S�H�jf�ZKno-���as��^>�#��: �d�����; ���vc��H:(���W��ckh�566�N]I�1уh\�m=x�ثKP�[�eJf5���4$�� }1l8�b�.��շsU���=����D�:�^�`��͚�٣��o5)�l�]���
9FAf1 Umx5���6-�m.����v�G��f�cٝ`�4(�l[.���yh�c�9�)������g�����n�b��$n��E�N�L�G0�V�6-,��f��n���/q�����Y�h�#��+)m��f�
���CJù�D��zJQ��+�sb�ch���q�%.��UDP���<ҵ�ձu����C�)���\�є�5�r����e��\(:&Ovp�9
DQ���X�+��M���͹0cOD��[.ɛ�&FC��l�f\_n�ۧ�g{������q��i�uo2+�4bӃkpL�j4���9B#Y����A�WWعuv��*���&�Z4C�N�!�$.sݸc�anB�-];n^�5]7LV���M�C8pМE��k��䋞���FkٷT�&m�7v�7�@4f�Ŵ�:Eq��f�f�>�iɦm:��
�x��=P�H�x����{�M�mu¨01e�3�b|�������Z��a��Z��z��-wY���RН�u���'1%.�*��e,QwR��f��4�æ"e��:ſ����|�,�N�	��Y|��1gm�NoV[�5z��5�S3n%3GXz��R�x����{��{ #^�^�6Ɵ�w��('NGF�+e�v\�)�6��t_=pq�Yⴒ��s�f��:CV�'�5�K�qi��y��*iLO.u+�@��߸����M��B��I��""R�7�Edv&��ݛ���=���%^��(���6$:�j��x�v$1Y�'R�Q��Hm�7�U��;v}�t0;2�$�o�k�`��8E�AN��[n��M����F#b��įD�S]60!_Y���8�iG"
�n�qTuyNB�yf9�&��t ����K���%kvY�RQpL�̢��( ���nSa;m��0_���f4F�zl���t�΋P[�#��nr�ŧ�.G`ӐūVZ7j
8�M�*Sdm�l*x0�˪�{��PoK����wHYǙ�i3%��1�̦b������=�J�!���z\���\"Uehj{s���ǘ�Λ85������y� �x��]�Z�,�Qb���Y�է�~v�h,����������(嗇r��O�U�2-\���ɗ�:Q{0E�=�M�ʩuX��W�B;6��R�K�3n��V��G}˶���݋�od4���.lۆ���0a!��n��W)�V�م[z��򰹤�u9�%ǒm;3#ŷ� �
x3\r9Ou^@�Vr��阒����DsN�]V� ��wd�F��5�����oZmڅfKܟ�f���6��f�&�Ӕ�
)��[��m��I=U)3�D�A�I�\ٕ�z/��:�	<�@�{`�ITtY�]gXo�dں��YG)�-{q�|r�B�s��Ɓ۰�M��m��2ι�F/`�0�y��F����e��ݳ��S%�2��{��՜�Q3��-	��Va/t���;�R哲:Nӂ`_P�㯋��9 ��7p*�`e��J+��a�\=v����r�փl�����+��<Xױv�s�vE�Jr^R���s�$�g��=(��Ni�L��D�c8P��&���T��mɯ9�ݍ��x����M�]�s��v�o"���9ۛT�JY�!8�F�j�u�v=CgaЪ�SJ��U�y�vH�WX;���X�ЈYmQۻ�RV�;�O�C8�w2�g
��hq�@Pw�m�0�wα,����"�8&m4�b[W���؍tp��f�'(
l�u:�� �4�VZ���,�r߅'e�kN��\�.b(�,)Ʈ')Q���j�q߁3��ހ)��C��U �-;�sb�gn]<�������pa����89�:�Ylb��5�5�8]���9[6��4���zTuZT̩X��"W��9on��]����=p�s@�(�;Q8B)gl�t����P�����G+&&����N�%iٚ]KXm=T�$6�	X��
����Cv^f��zMؤ�U �V�@����[`=$m�����k7���@��V2�K�������ۛ��Yc�	M��jY��Z5{�� ˂�����NF��(̲��4�sVe���=�{�����8
b�H����t1�)�;�F�w7 �,����]9©�D*�H<�eΛ�e��ق��ܻa�PK��7E|v��!�vl�4������tm� \8wh�0;�dc����w.�\e���3������ӆ	w�F��U�T)qhh%Ԙ(�J��W��Fhݔ�0�(k䰼go����*�Ҭ�YC�uj]�;�a\���ZH�K���cKA٭�ne]����S%�j=N��_�FIS��	������f�R�:�i����K���tҳH�iQMS%F+�j)v��SP�M�*;n�H��n� Ļ#װ@˶���%�Ƶ,��tشRm��L�4��yn �X�]��7�!���d�.��s������f!MU�a)S8�ϙ����c�bTe�{1[��X��2�8����n�BK�\���Y�]��oIwK�f��ӀN�%ɵR� ǎ��9@�"�!T(�a�Ĉ �aUqVe�kG5��ܽ��pmP�31�Vdl���jJ��T�ݵ5lR��KPN�\xġ[��P:�5��Ԗf,��h�Q��u� ��=�-�[�7��Š
C���KR��һi,�TGÛ	���\��\��t�����HA���8�C��霳X֭���7�-�T�Ե�GRh����}��!agq=��+ �b��p;��$�6��w^O&V�t�%R$�kT���c�sF˗����6n����� ���o)�8\�&s2��f��z�`���p^�6�d�t9ӣ���a��I����&\�w���NK�Z�6�І��σC�i2UŰհA�tի~��5v��dg33�o��Na�/����P2�{�;s��5�R����s&N�[��N�J�+N|�а�H��"�����&�g�{�nhۅ���p����l�r��%u6i�śY�Y�슧+¡s�@�i��s��)L8��˫��?SQ�>�y����ˋL2�G�4Nk�`���3�Yϱ��霯*��.l�a	li��^C��lvU6�N�\�,;��(g�WN�kF��|���V�]7h��C�^N��i9E�WlFF�֍{��ЩR��r��{�ͼ�Tu�C���;�q/���olr.��0J8k8:���3�ߞ�M��)��hJ�1��� �t�G�5K�v���>��X����S�Ȫ��2~�v�~�,�'��ةO2
���Vt�����7�$��8�5�sx^���b��b(W*cr}�852�\>ӔE��9��m6�m��ƣw gq�ڂ2^�q�����-����W
h�ư�$�_!�p����Λ��,=N��
%�7I7$S�����f��Ja��X�������¥\��N�㚢�sVn�ށFƵ+U0�#�r�e4\�f�cP,����oaG-9�~�n�G=tx���as9�ͬ��Q�5�oFX���^���J��*Va���4�=�w��r��(e_!���20����A��s��P't����Os<i�����Ӿ���K�:�9������f�M)e���&-
��4%�L^h��Y(gz���������j׷��FG�Z�䊟Ma��TmK�2�)Y��r.�G4Q�	�6E�,���v<����y�z�#կ:�kU���|����Xפ9��̧;b�	{�&�т#�Z��u�,��=PoL������!��Hv��ǒ�q��=�x.Ɖ��ݔ��1�}�0���j`$�$wo�z	�;f�\:���9y��ݔb�=�0s����⮐�Z�Z5�c&��'�f�ɵdtI�x#�uSPb���V����*��77w:zS�g�����,��{A�g���n޿�T[�F>@Kn����ፈx��yĠl��󬀝]	��ۭ�0�j���~��������?�����O]5������I$�Iue����eڐ\e�0�
����nw���w�uku����m�2�[�ݥ%�.+��Ga蚒���T3�oj�3���:����.��eM�o�W��Y�$;��<�"vEǗa7xx�řS�m�|2�i��/�	�'��_��X�z��A���
h��v�ӹ7�y�V4��j;@�I������Ai4� ��հ�^��zSޤ��feW��Vv<��S/5*�Y�t��$x\Y�EEkp����`:8�����ڲ1|���r4�{���d���jwn	��QgN\��̇�X��{LKBK�;�,Ȁ�A�$eu�%�H(�z��or3��U�^߽������f�T�B	S���*³��U�,Ss��d���y݌!�A.��:��k�������W�ǺQ'n���2)���OE�og�n=�ء����s/UP�R�|N�~>�&ӝm�ۢL3:�_i\������J�W�U�C}3�vXVM��ؽ|u]��-<���H���m�x^I U+���x�s,����J�U~�ϣ�����Ys��Ճ���=d���;u�}���^��PzX�U�9}+L�a��v*s�Q�}qfuU�Uз���N�U(�d*Mo�t���{�q^��'��rm���t+`���sAX��۶:f���cq�ё���s}M+�ç��5�K�J-�:w�fM���JD�����.��O��3�$�7�g��k��Ю̴�D)(5���/1x3�R�����#=������Й��c�Kh�`gQ��[��9�.�{��k�,��B����=�_�y�ݝ��J��Y�N3h��d}��%��(d�E�x��-YN���fw0�v֭�;�\
�&Cn
����1y�&�蘶�+u����{�2�p��xܛh�n�l؝��U��Đ�klGT��FN��A���G�A��0�M�ε[�~��.n�ۯJ�XԫHZy��l��z�@>$&�dl�NgFӷ��W��^^�R��-�mb��E��s&K[�S�E��~����p3�n`�#.���g0��}�M�̚�-�{t����&�#Ʉ�}��;�Ç�к�`l#�Õ��{]%	���mmK5gX� �j���wv;BQ��Y��S}W��l�t��C�V�p6���(MG�P�cSӗ��q*2��2%�!��A���lRW6�U%O*�i�lw���w��-u�@�5
]��&�n�G����<��>u��r�Y��1)�[`CN�Y���KΌR�e�k���k2���w��]��v6��à�f�˒�)�24%��u�Af���I�غF~�6%8aβ�_���OFWzҙ�DlQ��١CN�p�Z����Õ�]fK�aB�*4�ns��wl�|�4˅�H�Q4ie�ubi�xC�d�͙:�����5]�^7�΂�G�i��:�gC��Rr�Xc_��}Bk�Q���qpu%&��5��(��,�'k�K���˸��+�c��"���:P�x�{7׆{8���[��ݍ���p.s�4"�
�3NHw����������'b)F��wLߗ?]�T;x�����p�)���4��8q�=����$�sn5G���;*TT���郺��v�YIc}
j�9��OCͪ��w��!b'WXO��:�ʿh����v�x��V(l�i�Jz��r�L�ܣYy��;y�&��L��Ck��]j�l��������]z_.�q��aw.;w	����0�jn��d�t;�V ���Y�k<�X��ޖv6��%��c�R��e���/l��X��S��:}�KE�t�-��mw|^�.�^�1S�2��W&�f�M�p��	̰;��Z�����mn;G;���� ;�3w�y�$�s�]aZ/r{���{>q���C�r4�^�`w;�ǡ�<�f,.Wkʡ��أ��>W��u�ѥ� �^�AU��8��,�n�=�k��\���en��I��;��T޴BC%q��xp�;�MB.z�ˉ�n��E+��C�[/�+��[��M��,�lR��C\ݚ�Gr�7�O+U�
������o[�[��Qov�)��(,���{W�w� �&{���tYg)����V���ן*^��� �^nl�"p���ܽ:��I7t2�gn�6昼3��˵@|	}�2�=�<�g�U�W�Ur1'��88ٝ#���pۃup �;	��6�s��{A��Xr
�&M�I�dw�a
�=��NpΨ�>�8��%�z^���to����\:r�"�.\�:�V�n�����Ԏb�����:E����K�M����ABv_l�^8ks�<��˾������}�f��e��)vnn�1�٥\k:��8����_�ƴb�朹�)�8T�v�=�C�Z�}y�ž��y���}:�z����yG\��J}�4E���]�<�R?'1�l�f=2�7�����Э�	QMӡ+aX dT���n���,ܘ�nٛ����sq�ݻ&�A;b�;���~nq�xa,�Ԕ;=��+�WV����,覰��eK[�L.�{z�I�"�	b�f(��+;�H������!o���Q���,�Jj��m�C� Fx��H�;fx#BO���r-��:�ƣ���L�y(�Y�����Ѻ;�42R��6�@�$�:�v-���UEG�3tL��8,����@^@Ļ�yz���El�����Ec�E�S����J�{"�!��7/E;�3��C�f�/~�u�rNN�R25���&���[6�7҈"��B�8_��$��./��;\Q�]�,O�+:�Wl��Í1ȹ�إ�i������>������Y|�>�A�L���e�K�`u�|\�6M�x��}ԃB<j��C#�b�\�
�^�7٦���z��*��Lr��-�R�n�4(�ĉݛ׆{A�����w��74��:��N-���+��2��� -��>����Ɵ%������q~`.��U�(��]5�6���Kr�=wD6N� �ؼ]>���� �sٶ1]����=e��lf8e�k%�R]\��Wj��ZS[��\8݋g�@��S��u}��W�K��НE��ٗL��8b��6��4YQ��	J�� �x�?���³�AS�Ҿ�;�}�*�������y�]B�-���Q���"�@L�wݪkӒV���IA],�%�j�s�5�W)^.�xl۞,�x~�.ͺQz����Z٫�û�%Mu=+����ʢz�ȑ�?x��Ⱦ"l�=�3^����")ۂ�S��&�ڄ��u5{�i*�=�s����d|:�z��ˉ�G��������ː�K�����/d�+�����Z���\��9�F�ܹ��5�Y�m��Tu!崏�Bh
KD4���Ծ��샅���Jb�[me��;E16�9�E�VA�����Mr�ŏ/�~W�x��3��\�&qo;ιS�i���5s.��ཾ�e��,��ڤ��rxn�j��6!5�\x�Y����д�r1������I��^lH}�wU�W��J��n-�2]�bEm���dQ[�U���� bxo�_�`�5�3�oMj`�1�z৷�u�V`��e�6C�H�p��I��*l��x��a�G$)�������ܪ+.��ݹ��ON3����Y��l�s�� �ʍ�5k�1��U���<�����ń;Ǐ��;<7��e�>�
L�shv7���J�p�Qܣ��
��[Z�N�}��ֲ��p~N�s�^*��E�xf�;��b�������y������W3E��sRy�g�w���7����5�⫐�5���J-����*iz���Pw���p��mX�s%r�{����q���`aΙ��2�h�/I�!J#j-�ӹ,<�b߀�_o/]�{7�S҅��Z�E:Ӕ2:i�Ü�5E�|�f6 #z���pt+&vc�Hu��y���NV���&����g�cc/.yv�y����n9���#zS�0l�;��������YY+8��SZ�����.r�t���b���3ƭ��ή�Κ-�\�Cb@�����R��xe,�Cu����i���Qܛ�x*{��h]���X5Qr�R쏔�+j�!��oMNsﯬ�7}���+G�}��&�+᝚C���`؆�qѣWҌ�5%��)��h�W�6��r��#_,��z��Xw������O��=C>��d�!�b����t*{<���0�	�dYMn��]	���HћH
V���۫���NH�a#L���o�F��m-����VȪ)sD�P�m�X���nF�g���z����-W"X�99�$�3oWM
s|c�ή���.�c�q�GwA��/{/���4�m���-9I7B�b'g�5���|p�y�{��C�=ϓ�����u"�EYį{Rv9���{�<b���r/�QB{gp���u�Z޼���R��i�,��/"!�snѾ�d�:tw��t17�ԩ-)����x�WyJW[u����M���aN�-�,:�4��	����=�e�Ӌ�����c���=��z���)�1 �ޣ;$�=H|��&떱5ig�T"�Ӧ_+��vk��*Y���[���N8X2��CeͨaU��o����^]Uv]����&�Y~����;��	P�u�p#b癮���{��<+�j�K���;�=F;.9��6Ɛ̹���$��w�c�^�$jާI����;�|r�쳌��J�*l����N���.��^�˫�v�!y��!�V�ډ����ۢonuj�O���0���v)	x��	|��G�>��^�	{��Fò�����#L�ur�6:�d#hN����lh%�+!;�]"���h_Z���6�0ro9]��;-u��Dh䫙��g���Z E%��遏�p�]��4i�2�W�m_m#�G32頛z3YJPUE����d9$������[���]�R�o��iC�(�'ƈ��f�s�n�����.��G��":��(��]Հ�ÄEz)�q�un�ˮ�y�ۖ�c9�������oA�v]�����[ط�:��xSP:��+p�TT�E�cR��(�����K��Wq+]%��z����<<��]���qw�^��ѻ�Q/{(����$�u�ƶW����E�C�]��x����ǻ�;E��*�2
�M�t�W���>�Nh��i|o4)�J�.�\�墺�kN�T9�e�!��/�&��$o��-w�L��^�6(���q��]L��{�o�{�\���ޓ�5��/t�=�������_�X���5Υ��A��=��"Pޓ|�*�<��	Tq�H�x�U��ݧQ�&�G:�2���C�S��zn۹�������~���헗^I�l`C���m��eTڀ�S)�6��B�7�N$��/&�Bl'�f�|��ɃgCwXȂ����dP\�"�;̜:�N��E�f����֫��9 r�"�����v,9��<��Nm[�+2���' �9֜�Y�v`B�.�ʋ&i1��w�3p�d��Ɲv) �m@O�M̦KC���R���ji��Wgs����x�]��|��U�W��z������ޝ�Sh���k�*�2����csj3+@�5��F�i��n+�K2��}G�!��r�L�O{f:�v&��,Qrɽ�7��EZ�PA��'���f��d�r�Yx���\�{�EMCƞm^��v�Xݢq�86���+���c9���:����Qˊ9�nL�_/u��_���'���n�k-����s�-�eU��K�L��*������d��-�����+|�tANE�������vŞ�;(�'	�h<����w]9pR';I��a�w`[�Һ6.�#�t�E�wݴgw����t��d�݁�Ǫ�pR�z�/��߰�*&  ���7}5��ō�o^���3V:�-�����5�RN-�sM]�CFqMəڥ��WA�n���7*,��l�5�V܌�.�X��t�ky�PkN(]��f-�(��W�n��k�j��.�����S(9&]�Y����,��n3;|��.��&��ȫs�Yb$az{B҅ �ivm��H]��}YU,/�3	�J�\&���$���Z���oxi^�!��Οm�Q��ٲʼ��N������r��PU�w�����.���z�L��v�X
T�=�i��"xz�8�,z�p�%'ӊ��f���b�s�g��z�ːZ��zx�c\T�\��R�2��Ta&�.b�oE=���no"�8/1\�>�{;>۾�8 �-�0g��ԧ;i�ېa˝=��8:zx=�`�:Ok���WJ����υ;�nB9�=/��ׇ;ř�җ
�����F(|9w*�(��Ծ�a�hh\�3R`��nFa�Ԯvd�r�8Cɳl�NI$�I$��T�Q�!��)f�<٩�ΐ���G{���n��+L|'v����q�	��u��yܤ�E�wSJ*���}ˌW�FV>Id��u=GM�Bfl��Q�q�UX��$��$�I�I���Iܜ��m٬���d�DJ��@�dQ<n���Տ�5M\L&�0�j	���K��Q@ڌ�J�wK���k��D�)��K��C�#7"�R.ź�QtbM���r�"7����TQ����[q�H�b���6$B�5�̤E�[��#E��E~)*`���j }e��TAĪ�=J���hK�q�6�b2��P�V-R@��	H2)jE�ʻ�@�NQ]�|��0� �&0�p�?8�"Be�e4�"d�QM��~�
����/j	Ɋ�����d%H"\�� ���yF	�F돞w�PA������
�����ߧ����40�o�,��~��~���T|�?d�O�'Y����Ͼc7�}լ3`����L^�o$�tyvtd]��}�%�%FS���Y�ݮ�%2�	�u&v��݁�<�B�K��.��x�5�gzn]-u>�����Wض��{��G!�Vk/�]���G���r ��B�wW����R��	E�{Gm ��Y;�;�O�+$+@5;5N�M�P<�6.�]��Иc��U���Q'��W#7ú�_o<�c����ad{�`7#��s�
8��[977�q�ɔ��>˱�6�K0���iX��|����!o�N��$�i㤍w�L�p�b�8�;]Ś�<���Sjr��OpZ`8*n#r_�wti�1�]�/��Nq�v��@�N%�ϜݚoNʷXvaC�����8��� ��r�ϲE�&�V舦��]d@�}�	�A�Wܳ5���v�`���LжJ���ve�O�N+=P�۝H�M��/M����t���vo�pP��Tt"8E����x:�g��	v��������4 ��7�����7�SX�8U.��(�(r�[&�t�ǣ�[��|��I3^ih�a�w�z��l�d�vI�Ny�ߣ��xb�������|O��x�z��<-͹�f�rU��.��`K��F2{�
�ۘ;�[�%n�wR�c�p��3����]�~yo_Y���|;ѓF�2��_���p�5\���^^����4H��=��C�~�1sU�8y��U߶�a�g���i`�S����(CV��u��:����&�L^��Z�3��*ا���R�e�RR�4R.^CSwB��;n`gڏ���h��)0S5�e,��#�ׇ.�/<Fx�6x.g��=G	�'��ؼW��,�K�AW�3}�z��l�ڶ���֣o
������qS)f+!�=����2���OK19��%�N��s�C���Kt �O}��ɽ�mHfRP\�R���EԃͲ�1��Mf�Ai���̒W&v��<v��6���&��`p�I�}eN����/�2~�H���H��{r��Ζo� uh�᭒��Z\�]�Qz�7v_T-�N��Ƀl�O:6;J����[A��)�TF�֋�U�9ö�������q���9�p���P���ҙC��x�{��H��Z6���Q������^����8.P鵏�.��nR[y��]8��[��7˕�s_q�K�)I�ɦ��C�U���j�C�i�t�^��0��v�
\����qЮH5�%�:���!h���7��S|t�2�F�搫�%��x����Փ_ ����h�3O�Mbޝ�mI}�I,�v����ⷛ:��7�/Z�Pa�Yu��7�:}�J�d�q��L�4r���w9)j����L�2�9�6�����&�b�?mU�%�'��05��Xt�:� ���wR�z��@�K�����m�
X���ɼ�"�tW���jډ4t��zH�G���
�:
���([+r�^$��p�R�r�w]X�����b�dJ0�'K��ٲ��5�w���ԫ�z��k�P%͇F�Ϧ{�8.ݏo4�m��v�5��Ʊ�R�;�����׫+�UM��}�4�v3��H̺����Ӹ��$n\P�c�3}��)��d]�-�t�GX1����ɺ�=�tGp<�lG�������$����1�ey�hPŸ�𷶸]�*��[���fn�6Ί�c�3LNPe�Y�xw�˹_E���A�G�|̎�o>7%�7',�h�nGL��^�W�`�d��^sS�J�SZ��캒r��v��w�i^i�F��K$��*
��������{}��;lY׺�<��12s��!�WJ���N��Y)U�Z�K�Ψ��
N&��M�;Mu��Af:DCi�ɻ��6tb�c��4 G%Z���3j�搗<^����s�0x��V�	K�!�=�N��{�\���L�{z�t͔��-#���q��0r�b�ށ�;p��V
Fr�� ��O��v̎���Х)p���|��uj\h�pz:,�ON��اv��/{��q�h��SV� @�#�-ޖ�V�v�
���7���*]��7��n[��^+�3��p�~8;}�h?��+Z��?^!s�>����GQ�s|�M͜W�d�Y(��<���5+S���­׺��i�}7}2{;���H��'��y76q�?��s��*C��/��b.�:]���tX��mf�\��ULGM(s�N����26�ʈ�sZ�2hG>7zY�1A��ҳ�fY�vR'���#�5I/�]BR/r�������������M�����ƾ���b�pm_3y��F��A	�y7Cd�fWٍ���ژ�kj�-��u|	c v��B�{d۴��@�z�z������ʇh��G�F�k�����=��u۾\�i���8���BJ��i�n��b%��9����<J���.���"sǥ:甞8ô�e�<ُf��od�k�G���2��N�2�)r>�ʫݾ{��Yʥt�r�{7��.��˨��=��,�[F�AR[�
��k8)�� ʑ��u�{>+^�"�:y'rd=�_+�r�u0]��]����:h՚���9��ӂ�񆫍��9�S�!2�)��� �W��3�9�ț�0ӭӔs)�*wؘ����JőS��}N�w-�9\�sd��� �=�������k�5w�T�@�Qv��Q��љ���R%�x]� �ﮆ��(�cc]�'G5�H]֝AE��*mn\V�-N��p%��BLM��%vN��0�m~{�f!.�£fiVK��`�s�gU�2�R˪ۚf�,���D:�bF�i���:�,��,'�u���-01�Z5��z�*G��'v��]�bC�3;(F	���N��#ۀ+!�;�[i!��Η��$(�ҜZs���L�'M�@feI�kKd����V�S*,�Tx�ȝ����W��7����Ì���nnF{�˱p����=��ў�}w���3����p��5}~�eZ&�zk5-=J�+����D���I��n����\����8dYY���\�7�^p��ʻ��1�i7����@oCpM���]n��Fr�����l�9�+���ͱ3�qXp���L��K]*�����֎�u����O�8&�X2�G9�l��w�  k��`���$ ?g�=�[P�[����u����"�Vi����{=���*.{ٌbV�<��6�Z�YY�8�
F��xU�5�>��a��UkD��K�a �&� �m�����[�3��ͭ����b�M��T�v�Q`8�	�"��v���:i�Ńӻˮn^�*�î�C��Bˤ؍m4{��V)��k�ZƱ2��P#b��Ս	��O;.��`��{y>өA�)

��3������ۭF��&��
1<����e�5�-���4�XaU$p���|xA7vu��V�e)fz�W�pgnu��w/��4���E�׍���	e*�}����Ό���p�1�C��f��Y�*����m��x.�n�H3�l[���:W���O�0����M���0	��9���;� �Y��G>�j��r7�B��LE���QT���8{f�c�=ÅwVť��{��Vn�yR��qZ|�{{��ϊp�!@�LEG��yw<!�q�7uV^�rm���1���l��Cvq��x;'?�Kܶ.��(uF�gJ络�5Y��sF����e�l6��t�6;7�a�=Z)��\�L��w���h���x1�*��p=��L�40��ԧ����Dtl]���~�(2$y��=@���P:��X���gc��0�i��v��v^U���Ɲ�8jw�g/MJ�+vAө�� �����v���;s����r���VXk*M��l��1^o�.U��8I�_��T=�ZɊC�}�g�����l��wF�{�r�Fby����:]u�NQAi%�N.ˌsA����n�j��6ˀ��r�v�v�\��u�,�%�t$M2fm3��܆n���g�K2�T�����|�ByjRR��ŗJ���+_)7�x5c�!�~�8z(�t��:�i����ydEշYy!*K�:gdx��h�d���=cw����k\V��T�m-+T��z�n�7��pd�χon���Q�Xɕw�=k�;�oQ����Ud����u���L+�+d�㞹�����'�*� ��E�_��x}�z�+�;��hi���Z������j��):�s;u�����Ȓ�ٍ�2�= �whI��ܫR�Z3Q����<^�;G]��	�T�oF:�q7�&^��{����m�Z��Z&!����v�g!��q�֋�)n'�}<��\h>H��3����/��O�Q�+G�����V&���q�4{��{B�����N�# �Wj�$w����6�ȰX��6~�g{�g��|�,z.C��"b��R�4KˣX��.�$��� ���S����eIkEj�6O�ۡ@��)d���]�ۛ�v��8��9��͍&�a�*�%���u__D����������:�l��V/�v&^a���w�n��o^���to����&<�`}��y��q��b���U�=��+��o�Z%�1��k��H�G�c�i'�\r�cn�����fJ��"�ff��|
3	��}�$�53E>G� 6�Ș�#�YO����'D����>����.��y��g`z����\7^[;�=��A�G�>\�L��A���W��ͧy�B�[M((���V�J�uƏ)������W��������6w��(��Wn9��.w÷h�
������uW�l�㾠���'�zy�r���尬Mƴ3��`�N��Z�.����6���oc�fǶ'(y���$P]h����������9�J_M}�l��V��I�[n7�/q��Z��)�%#l�p֙��Sw/[( 7b6Ck>cS�t�f��87�V%[�@���l�=�t1��ӌ��s%�Z�U�Okr�]V�{��t��v�s8�n��eJ���^�*�`����=�݂L�x�կ������e��P�d5g��nX7d�_�,�H<}qu��ށ�hzWѮ���^(j��B�m��Ǝ��~ɛl�j�k%�u�LuK5�d\��	�$���Ԭ�Cj񋽻���Eu�B���vt��3
�&���e5,�9j��}IT�un�]7�1S��g���=����C�d�y��J�]ds��)��Ȫ�R��+�r2�A�\�bP(�Ÿ.h) ��'~�F�7&�:L��wyv�dq�g��:� ��c�>y^ZЪ���'�k�w�sB�"N�X4y}p��#��J��ǋX�u�@��UISf,���v6J��腌^�D ߶�_g�M��]R�a;��{y
�;��l��}:xd�V�a���>� �$
/��V&��5Eָ[���`ɦ
���v-\�v���>Y�x�c�3�{$)l����Y�4��FUFE�n�Wp-�=�1�+����)ޒ`"8(���rzz�po.P���+B̻�
otG]M��q�`��/�v����eˏZ��k��x�|W]8ʆJ�#Kvz��"�M1��xo�.iYaՑ�6�#�}�s~Z��!�H�HL�5^=os,;�FZu��ˬ�d��o�ьpRG�vYEt���V��|(�uh�p&�;��b��ʉR:`z����',��II5��nn�T��ep�j��M9�V�vgW�*~9���Q5y��}����*�`O.�"�g�k�:�Ԋ� ϭ���(��Y6���;f@앍N۬��ܡY����#A�ů�+���I�^��m�M�b^��"��i���V��*,M����	��C�j��5Y&yhe�
�ыt�!b�x`�8�Ou�z��_����Gw��މD}g[j�����צ;S���~�}tC�#�ջ�r�}���L�u���[���E�La��ϲ��x��KW�Wp8�qY~ȟ�-�4<�ϸ}�eǈ�w캬d�۸�B���TA��z��P�W�ɿy,�]1���SЏN�R&�s�,�ߤ�������Ж�.?L��7�����~����ڲ���9�(5�c���N���L59��@��y�A��}�F^�u��S�-�,�.��h^ͽ�}��s���&��kCbs��܌	o�{��=3F��\<�g�x��A��9�lۦ�
�ݥ$�^	��u�ߡ���v�Dk��U.��Iog�����B�0�<'�/���5z ��o�4Ϻ�P]g��3�Ow7+B>Z+//7���}�����˩lL����>���t��,s� �O�!R?��j»��4!u���!cd=�<T������Xb��Ĵ_����#	��*��H��]
��x�ǆ9�z�t��V��fR��$fɽ���YS��&{Nֈ8B5<|֪�8=���zE���-}��C��-���y@��j��P$�C4�{�@��hr�����"_>�v��ŵO�ҢC#�T7ċ��	��_ s���NR;}�fo�<���~ѵ	�s��jj�AE�[Fԕd٭P/��ͫ4/�۞ՍAo��x^*�b���N�xe����6U9���~�2/!kp��[�	4�W�oZ#Th$�&q=�W���tj��2�U�rnٽh:��Ώ(T���c6�g:m�AP�����(��k��������Hw�<)C��58`Ӭ&����������� 
����~�������W�s����/�߫������kkkkkkkkchmmmmmhhhhhmo����e/8\�RC��"$��y���_�$}�|=����<WKë/Wh!$����3Ĥ]7�;���#�lY�Ù"�w�C�H9�wC��6�ؼc��`�����I�}��t+&)Z�Ϗ�7�cy]KO.��"Fi�:z�3����0L���<.7Y,���E����j=�]M�@��_=��È�����l���3�n�<1,���	��KV������n�vkVU�EJ�K# ].�����QV�}S�ci�+o�X��۾���\�����7;�����^�U[�"�Żg�x����L�Ύ��^��E�הN��^(�ɻ�&˦����MuM��־�]{u,�F�'ȳ�k]��/^^�==�p��X����3]F�f��5���l劳,C%����8��\�β�mN��#/^(/j���~I���3��w'םs��ѥxZ^GQ]����kl�B��M���z�#a`��n8��=ro?o�bJz�������bH�P��ϰ���xnL���o+0,�l�p�6�]¤,5ou53���v�[Y�VR��9>���%�L��R)A�j��yoV��݄�y��mC��}��S��g�`ޞ=�H�(̠՜ݓ�Q�6��r���JT���aM�^�bA�%jG9A5&�P)�ign�M���u(�%u�
%Ta����'�N2Åi�e�!
J!-���(�_�_���ׅ�c�QE娊��E�KQ���J���qAU��[`�c�"'Z*�6ɉ�+Y�-�DT�ն���C�?=�ADD�SSDN�TCU&�1��I]�D�F�U�MV�D-4h5���"h�!�h*�ձZkF�� �b
h)��������*�**)� ���:��;`�����SEZ���i�PEEQE�U�úpSE3li"�����(�DAU�h*"&�*&��Ń4lb��i��*X
gcMUU��"�1$T�F��t�UEQ4�h�;b��Eբbh���(�$�Ӫ*�(���;h�(������*%�&��	�lQ%}�D]��V�kmV�����"&�����z6�S�Mm�����V*(�"b�kj�1���v�ضt�Ղ	��ћ刨��1��ڠ�"+XjB��&�&;=USm�-����"B���SL��
���������A1�Ɲ�j�)�{���:@��)u�4��o&��ʞx�W\�e������O���9�|��.���4Y�ʣE���L�k/�q�@�+>��PӺ\f�h� =E�����o�������Q�WzD	�{3]�=٪/��9��s����^�j���UNSlوԓ�&�K'�>L����s��Ɉ�]��r��?6}���{�~���]��ٷ�F��	��6E��c�1w �;�f;G8�:�b��~�ޏIoT����h�즺F����~���>wA��/:�����B����q!�
w,�p��S=3s��?do���^��Zgqʛ��i�=i������`�<���'�~|c���8���?m�#�>b�����4��E���X�H%��]��6�߻\��}4��̂z�"�B2�O>�{w��������Ɠ�l��*�6���@�Duܞﰣ]ޛމ�C��~�=<�-q�7]�xݮ�]xHOog\�)x
�y����7���dH�o*�{�+�T���m��D.�0O��&w3�IbY�;�5��}C�\��Mn�-��WHˡw5٫2����9�V+S[@<�'��j齇�@���ײƼ{�6�A��HwW�6۹�(�|�R���,���������{ ���،����mw3x�G��%�
�l�\d�q'3P�o�zW[�����.���}vz�n������od>����ƷT����>)�?e>S�H�/��N4o�Y/|&�k*f�یc[���m�8Gqŷʹ�03��y�dkF���H��_z�=-�<�yG�u�r<����Z���S}{��췕���k��\��-	�����S�� #�W�'�A�6����5]�r�~�����Uj�]��	���d][���+���5V���2�=ʝ�������5�nL�b�ݸ�����wvml "����$�l:�w�6����͛�G�{��AWj�3���o��Pջ�8�}'-ڤ|�Y~��wu5u+��|�/��|Wa�2
y��{��� l�`���&������3���9�./n29J��0��j@��zx8b̻u"����9{^oU��۶�&�8S���Pa�9뫟Uc�re)����c��5���KW'ٖs�K��8�uU�rc����Ѽ��O��b��G���	x!z���'�cj�y;��i��90�W�X�Ν�GL�P�"�v];=���9��^����n��,~��w.��uf>�\1OB�����n�0]W����7=*zz�gw��$՜كO\^��p���Q����&�_�������y���4���������JyMs,��#�8L�~���x�{�����tWMߜ!-�4���>�x3{m�w��X��:jX���l�pe���U\dy����K�_5���}䏮����$�Q��Y�H&W�o��}+/i�r?���5+��O6��B���|��ǚa_�)�<��ޛ��L+$�>oZw�l{�Zm�;���h��v{棗57�����UͫyPڙJt��C_�foE�\��5���e�p����1�Mη�/joT�{�{�3a���q��\�x�Y@�|���A��"�;U�C6� �w�&�1���D��/n��:s.�Mho��@�ك������U%���kW�a�^ܮC���.�p3JvS֎����[\ ���������<�eG"��e��׹�}�9��V��^���{	YR�n���/��>�T�u��s3
��'��h�el>��%��:	���hw9���u�RG�h=3��Ius[�ԉgd[�����'s��=d��%��`��U�of��;�5���)���\���=Y��]{��޷[Ih�}�ݿ�� Mz��yH����K��yE�z>��I&��7=\S�>��ۤ�2v�d���Q�ڶ�:�5A�R���~����@h�T_��q�	��'���H�w�2F�<����'Q54{dwݧ�'xj����2��V�B�
��}�=�v��!�u��D��ެ��o�gu�)TʄU w��fp�5��6�3�|.Mƹ���;�s%x��[�;�Ƚ��������Rh~��Fku�o�a���x�=���m���g�w��`�2�[,�h z�@�͖,`�;��g~�ى��ƀ�ov\��1�GNe;wn7a���׎�$"1�շ����9�j�������YTO����\`�3z�w?�z��v�cS&�I�kվ;J���M�|���g��@��F���{{=� cU=��yl��;rO������h�}G(8r�[�ֱ#ӝ�.#��>�]e��ص#;�lǜ��8�6�yuJ��Go�;��C�M�ڶ�^HG�S"�9��Ż�;�9��I�ƩD[i am@R3�����H+����J�B��ܓ�h�'��*���ڧR��q��3��C�'uʮ@~+�Y��,Z�w��?NR�:�}o`Z���;�����[#���&��<l�e�@O���R��������G�B���)��7V
�)��8΅š��	��B:{lʬ��/ێ���;5z�#Ir�"�o{�g:��K��N�P�Ӛ��	M��-���?d>t"A}��ŵ�W�V�,���O���/h}���;��[>��i��.[{����á�����Q�0�g׺Aγ'NU��Ͳ5��3�j�l��3����� �\+z���ҝo��Lx����pt(�±��~�x�d=����ƺE�ĵ������C:�k�'d\���r� �OY�7\.�~W/^Hh����c��2wl���ٴu�H�c=���� �Z�:2�e��w1k�A�|��{X~Z��c7qL�Q*ҷ&\E9{����.���7�%��w&	�X44�����e�/)��\}�M�O�����1�J\j�����o2m�;�����xeL.��hO^�N�wӢ�qB�k���E��t�U7,Ҟ�����d{��Oy=���"��J#��yDs��t��\ovr���[Rw_�_��i}!y�_���o>�>y�N�Cx��u6�O:��9�8xs��C\��{��۽xV�rͥ�j)����;�����Y�Jk*�P�;?\s(���y����W���?`��}�a��jW�~ǉ�_���Y��4���.�_�]9i�z+���Z3����Z��/>�s
���-���)��Ӎ{�m�Pe ��T�<�9}�*R>'�G^i�9�C@ם�vA{G���f�ț0ca�di���٤2_���8�W��s��A�� �u{�וL���Q�{�;�����מ�����R(E�i]�o8k�I:9Λ��\�vE��XjV��d��j��Z�<d@8⻢&�r��[�Oq:vν��/qFJ�w�Y.�x�7��Zx�&uWs�=�f�l;?V���V�aa	ڊ+���傡r8UƱBö����=�r�0(Bu
��oOn��3)��V���[�\;��L4gԛXQ��٧��Ո�qgG�~s��䥭&�]�ȕQ05��-o���|�<�/
��շ�}�LR����宇]\�RXŰP�"�h�f;�l����>�W5'[4�1�\d��w�3V�<�ϸ�W�Ϯ�L��6�>�c�ӱ{1H�6��w@�jٞ]�����y}����jn�r���ofׇc�nM��tj]��'9�9����[t�w�9�Ot�����"I���/I�˜���]�j�L�<��lV�cw�I'����C�޸�V�7�w��]��/���z�#1�ƁBvg�6~&��K47�.�bnfn^�YMo�Z��w�}'�^�7�:�n��c��nl0w��a�q+�h<��]�t�ԟg�����zw�:���W�5Ҷ����u|���'k��Q��fyxI��8��Ыyd�ν�Ӫ��"�d��+)���}���
]ߧH�����.�v5�go뭜^�ܠ�Jp�k��N{ej[���Ԥ�S�s�,)�^+��Z�B;��r�ö��m}�����G�˗�X~ۜ�E:X�c��9F���_n9�3l�ӥ�N����l�Agj��G��`��!�Z��^�ϝ��r}ۑ�ve\ڸ;ޣ�FDk�g#{)i��BP6R��7z
ܻ��њgM��M�Q�^;�������`-?�|��Y#럗�0�߮v�B��\X��=
�	׻�PM�C��{Fy���iy@�ގ\��͉�w%	X�]�#T��G���[��F�Oǳ��%�'�5��� ;�殛��0$������F�<m˩ʔ��Ϸ���i�����3~O�ߺ�- ��}ʪ�N��_7��L���dp�S>����^8�w��K9y�
v���o:��t��&Y���\q��(Jm#�dS�f~�q�5��u���Qa۴��L��=��e5sW\�YzPj�5 >�ȭ
t!w۔�����b� ���wt]�]��^��ǝ�_q���:���e7�ݲZ��㑏P�QՕG�j�	m
�Q	sB�[�ly[�}f��J<t|�{õS��xW{z�V�
ʝ�é}��l���+�eG�<p���Κ���_����Zͼ���R�m.��]9`�3������.���648n��	�3l�hJ�ѶI0@�U�ټ�:o�9����=מ�z*?禡<,լ��(�����]>}����c��ח�po���{zE7<�m�U�|�VS�B������ �9���ͧs{�M��[��~?M覜·�#o@�̩ݯ�d�lkǬ�n�e�j;9������c�P���� ^x�����vW��ɘ�&	�����<��u���o����qs|�Z��������+����%E�+'D.��3���{���Zcڜ=��#[Z�^k{��eܱ˕_	�^��=T�n�ލ���PK�%��jw�i�==��®��A��'��qV��=fI)˕���5^��~��f׬*��[�qb�i�߆��Pjfπ��ƻk;�$A�s>^�q~�2��������ݚH����!���s�V�r�ǆ������G�|57����i���e��9�V:ra!�-d�N�-�y9��e�9M�py�ZB8=S}�XR�sÝ�?��-j��<�������@X��v�+�q�̾�x��cQ�*	wǘ�n������g��Pb��W^o�$ݧ����6��:b��B�D����W���H� =�����5���5'�WW��Mސr�SQ~���x�1�_/_8f��K%�%J3;!�S�s�H��������eH�z�8�s�k�EM���q�N��=|��k�ߪk:�΄x�g�8�M{h�ͮ�!Ι�&�t��kh���s�}\�V���7��Tn�����?��O�m�a%渴����xtm�;�'�OK��������ĺ����'�M��e?eq{'>�0mO?W��b7��͗;הp���\jrYʺl��k0��¥��@pr�!�-�ut{bv�W�U�%����λ�f=[r)V�m�v��N���뫫+�K���^�tnXչ5���y'���7�/^�zV�U>p��rͯAO������j���Ay�ӱO}��ӽ�����ɘbг�Ÿ(��n (�4�3��66�7����o۟��>�����������~�y矶��3 ��ɗ)���=7�,2�bw����d'�A���ޙ��Tk��wRWʅ�d�*6q_o�R����f/g�d��q�x'r����_��f��MbFl�$uT�*M$���M�\�����p�j�68�^�%FZ��Fo1��k�[Z�A&\�Fq�6s�!�c��]]�����}�S
��������֯e��������;��˩�D���w;j[��M�u��B�e�OYƘE�{��8�I҄�@5��β�n��魋�����.o_G$��n�\��W��-�e�|ҀKݬ �b�F�nQ��fmdt\��q��RM�#Z�x�,����a41NPJ�W���-�k��<4c�͑��zP�̉dN]��N���Ԋbt�i�rr�i�����AG)�}�yj���I#[١-P`)k�/b��r�|��l@�>�p���L�o6!�¸�mާ��G�:\�ڥ[e
vg�n�lw��-3��ei �:M�g�3#�o��wx�92oWA+�Vv���;��E1�q�����̓��r��d1�;��[�V�#�jN]گ�p̓�ܙ�trnL�^c�[Eq�ƕ�
���\�-y�ԻB,���w�{CF�v�����"WV95@+�P�.��r�U����i[���ƀ��3r͆��ٸ�o�� �${o�R��=�c�����j�&w��@�]8Po:a;�I1�;{�����Z�i��j��e����1�l��{fNV�8���^�=B�mx�#ca�vZ��K�\�Y/�^b��9fn՛I�GIz/7�]֞ƣع�mib��}����$.�V��I&�����O0p��DM��w{�h.&;wm����æ�=3mN�e���^�YÏ,��f�W]�޾�}�����L̺���hr�w�W�%�vwޮa���/��q<�:�J�+-����0��-���#�$�A�����^�NP�[��vb�l���T���5�-����=��<��;X���PeۻSxc�XyR��VϜ�q�:�b�#��>�f��ޓ�uh�\,kw�u�wHP�-���ΆQ[š�W�=[�y@:p�/���I�����F���X���3[�b�V�!Ÿ�]��3vl�rv&h�	�����4�8�j�F�Q�[�B�r)ڌF*@e�Sc�Իh`O���}N���cM^��q��v#�YL�+/)�.19����"9���BQ���, �H�z4��p�,�9�bf�V���A�@]�A�ŷaf�v�:�%*�NCvb�*�з��Юv���e�ն��o�²
�L��5�{WSʂ�
3s+�e��+_P�:𲜺����dJ��N�ϯ��u�F�S�@Ʃ�9Y�ά���z�D@�/mt�|��v|zEAt���&�{WG��S�~*/��o�����I�������s'2h�?qK �ĘA�D�ւ���S�ɫcmlkZCKT[ij&�j���}��(:>�jt�h�)�Z��b��N�N�j(�*������� ���b�sl��M�ն�mUli������~,�A��j�>�����P��U@D[.��Q�����e�-�؈��4̴�����5{ۚ'l�Vڠ�!�c(�v�1i3lJ�b��lD�{4��qGZm�M#QE�����N���T�0U4�K`4��F�b4[SCILDE4�kZ��b�I��!Z�`�!�((�N���"���l{h<��d4T��M\ꈖ�R'ݪ�"���1���ܸ6�Tk445�7�OF�h��ζ���t�6�<� ���h�w8��Z�Ӡ�<�S��s��~~������}]g5�}�:.F�0�׳ O�c��M�u����r�zI�e'�̸vp(@Ξia2bF�����q~�ڼ���̍nk#�=#���9z��'&�N�	�G>��⯯,�׹������~?B���5��9��n�v%l�w�mq0JSi��3U	�Ws*�lV�I�S���陾�0�����)��h�иm7w�f�����x6׹K0��b#Ϋm7n��9�r�_�ܥ,��6�g�|�%�j�H����Y�|��ema��4}�^����@q��}$��i��\""�zw���IG)uv��}�<5�"��Ɩ�Q04��*��2e�G8�n������y}�?�����J]�l\�aW%�uN��M�e�.��,nE�w�H�h�{#L��)uٙھ������}�O���o]�I�����ڔU�`N�����;H��g�Dl_$��WJ���۹�_�%����Ro��*��D,�O8��4��(���[��cbn.\�yC�qb2r[.�.0����aw�} B��и�h���=ڕ�X.Q^����J�.ݐ�|x�q��fc#:��3Vn|�w�4}r��@�	Za��O���1@'>3���^�`��G�{����"���'t�w4ƣ�S���ӽErF��B��sk�χ���'l��(_Fi7_o\XJ!Y� ��[;N�G��¾��j���o����!�!����Y��M�j]����u,f��Κ���]���z�E1�_(k�S�}�8����׫r>���l��:YAԓ�!�2��GKB}�0��Mԉ��"��뉭ͥ�m��F��vWJ�ڮ��{�8�p'�Yq+�1�1�2�	��G�ب��h��3O�^�/3�j�۲O��񤽎#�c����e_zr�{�H;QM��[n�d$1iE���萮����vM׫����ң�K�]1�����*����㑏
b%[��*�Us����Z�>�X
��}��0�hez�vu���c?���`/Z-��5���9������^6���0�f��_a\vi�KW�M�O�>Z�P��Bp@��|�gS�A��\g�s%�����mN�w8��zܭ���"���S�������i|쯕yD�Ԙ�HQ�o�zE���P� 8m��� .Ã�e�9>rB�`�k3���Ζ�U}\P�3��qP�=��L"��.������F(U�*Z.;�aIk"�
����`��s{_z����"���+<Υ��A�|T�e�-��ܦ��]��Dz�P%�TQ��{����M��r���^��y*m�჏l�,uf(�ߗ�D�"�m�ai�=�^=:��1;�翛�����nG��Q�ڠڰ�S�pP�A�CY?*FY3�P�	D�7�;��j��t�Bo��6|�,惩LY��,��%��hF�>����Ws	�1���K�
�<��r��#R��VŲ��n������Aq�5R��.� ��G�w��s�[�-�����3����������2���\֢����z��8���1���c��˵s�«���H����&���u�"�����l�g��6[!s�Q�<��;�����׹z�T��|����/k��3F��5���̃��|�/���{�[N&��9t'%6�5��#Y�V7����m�s���Vr�Г7��f��e�:�N�}�@��yj+��b�ә����w���~&K�L���L\_a�k�z=�H>�J��t������^�㡰���j�j�!�|�K��H�q@�\��2Y,��'�a��w�1`�J���W�W�i�hZ?!�����9Cr��_�9��|�*=�zhUw*2�l�T'�Gs��%%�֨}pvu��E����wO�zI��MZS�is���>Aa��J�	dsT&ʍ��Q�z�Oz�b�/u�3��	Ы@Kz�7��Sȃ�(R�z���- �U�?P�M3�Oj��O���
ѭ5ĭ:]�5��γ�Ϻ�Q�z�e��9�,��c7�a,"���A���Q!N�קbO�$����̎Y�.��B^��P�W���Uǈz�:���[u����2��,����D� n*۔�kh��Mi�Zy37{��et�L�֋��V!1vÔomQO��V�ع���k.hEl�����M���a���f���
�l�8��Yǜ^���,��L�=.R�kPV.��}���0K���������Ws*��(d�D��i�l$��f ���#�)�<��GK��
�D����1���]4=���n[C�oE�,9�'=�1��ݪhj�X��P�o!,F���r��d��3weG:,e	�[۝S�c|���1]ʌ�[��N!)�b}�n�gU�kg!	�E)ƒ��p2���Qm���N�mݱ�ʈ~iwƿ;�[e�8b��T��P
��&��U�c�K7�szw�,B�25��D�����m�����C��Mz��I���]]��E�g=�{�(Z8�0�vM���7q]F38�0�͘�5L���ۭT��{�q"�ש�+9��݈wc���@y�cT:n��U�%�Wn��P��uk����%�J�7rSM�V�Qw�1p��\[L�����(]Y�X�����ӳ������&5�Y0��*pM))��Q~k]�C
��[%G��4�K+gy�1/:�E�r7�#���S�F�Ӣj�x�E;s�Ȗٵ%�>��%O'.��G����l�>����`qa���Dl)FVc7ۖemE��-�"��v�����6�ȴh�C��Y8�$��=�1�f�1q٠:b�c���[�냬���M[�Ï!��y��
����@��˫A�E2�l�h3&ө@V���"�q-7��yS:��?y��S���� ���Q�O�%z���-�~wp\g�k��^9��"oX�L���TZ���j�@�P*�pL�\�ܥn��~�'�[�n��?���݆���	�(`2�|��aNG�ɖt�y҈��P?59z������*�˽;��ZqG��	�ƢFK�H� ��e�A��)%�m/���|j���ٻ��=D�PO���'�.�*V@��PսP]i�����|�@�v�@e--�}e,9T�����AA#֭Ǡs���6��!�[�5���W��4P����V�숾_xe��X�¦��Ρ�i�hh��./|�����;v�1�p��rvnFp�c��ͧޙ����1�O����i���%ĔnAU��{��Vc)���N]S�w��?���vAGC�#	o�Y�Zn�m�e
�Cȣ�2位�w���U�$z~�xM�B���k��Ch��ӓ��}����S���Rʶ��l�3�M�������f(����j�\�ccB�2Zs�v5N9�l붤*%k�(A���b�`v+�lҲ��Ʃ�w0�n��U������~���3S�L�9j�%; 8�7oL�����x��qS�2���[l�9ƕ������p���55#v�Io^:�To�����a�rٚ2�X�����N��+�/f܄nM\"6�D"����c���6��`��׸
|6Q������d��6vh�ұ=,x5��WR
��33@ � �3&��J��ՙH�Üx��:_^d?���uσTRr�ǟ��"ʍm���N��{ŷlM2��jGsb��ϐYY3ЎH��*���e���)lt�'���T/�M�������g�2�,fFzv�w��$%U���v���Ȏ�.ř>K�5lt��R�d`&�Oa�R}���Sx��Kd�Ҽ�o��ν˶��\dg��|�o��܀�=��x�-6M5�.ۜ�Z�a�7h��0��+;�+�*�j�׳s��Ԡ�I�XE��q�`��\���9b������f.�eë�yB�JL� �䴧����q��YP��c�H�3��&�� ?�y}i�)��ڍެ~�n���@i�S�Eݑ�^��/�-��g��ӝ���+H�`<��we!s*�����O$�<��g<�	p�Ec�y�F�t�;���Y�#4UZ�L`g.]�oj��ۜ*���q�O�Dギ�'���=K�7y���@?S�&!�J��x1�����Byfѝ;�X��^sb_3�b اS�����H�x����	��6�[w��Z�;���8�T�!�PT"�#�B�,�f@�F�2�'�ۻ��ӭq��}u��m�;(���Ѿ��[R��� ؔ�[R
�p�M4_&�7sn��)e�s�3��ef��f)�gw��_`U�"���,v�q��� y6k�����l���	����0d3o3���1���yn	I��K�܃L�S*ݑ�@X�W��(K4������<�ia <=nǛ	�Sc���S�v`E�Fw�3 �Ns8�����C�6{�T����ӈ����?4�z��@\�����I�j͊���m�2� f�z��a�A��)�CT��K9sCeծ���Z�F���Q��\�4Қ�]rt���-߶�Z
�Ocײb�Hzik��2���ε,�[c�kxSW�d�?��n�:�#n5�&Y�{�n���7u&��	O�yS�;��=��>՞҈/>[~���/؊�� ��~�VƉ�Yi#|;�.D
�G�,^�>uE�{���P����䖾�[�!�:���-ϱ4ﰺ�-m^�kU�׫��c��B�3���H����z�a��ȸ,�f�c��<�3��,l��w�Q6��l���]c(�\��)�ie��sx�.M�G��Y��@d,}Ћw����GWn��ہ�5�R�t�y4��}����A�I.�7G7QR�ך�!�ٛTZ��gKo]=nyL�LA�����h���z�5��y.�L�V�	0�A�U�(t�O{}!z�J�9�М�md�)����Z��o���rsW��p�����%Ȳ:�r��@�,E�8nUYc�*�ߠ��u߽xqTC#z=�^�aUzr���1"�w#fD-[�
v��q�p�)�m��
���߮����jڪ˻�}y�H��7��NĂ���r�S��Q'���,� ���	`Z�<���{=Hp�~o)�=���f�QP=�W����|+6�=x��a)-��,�o2��W��cY���yB�"����L����B!�?X���6K{������:7�$�K֡ʟċ��ʝ��x*{��o��d�<��+� �����8N?��18ke��4ɍ�*m��·��N�~(���y޵Qp�1�n��F>��Ij1ba�8f����p�����a,,"�N�|��/�<��~{���y�_-����R7�8�c�S�z\�뽉)�N;�:�A��U9C��ꗕWz$�љʱA�̈�����7�v�xA�}���KB~�|tޑ�%F[���1zk8�>�_tB>��2S���,5ջP�z����rGw�2&p���AX�u�&♙kOU�]�T��0���Y1M�J��>�Mi�i�����d�/�G���������<[�j]]s��?=�_�e�VT;���J��0����������|Z}�*���JT?5��w7�0N�=ɩ�<�U�u��oiUt+-��+Kڧ���rl��*�8�b����%�6���+eA���ѓ=%�wP�[b���j�Ū������  ��_�W�>���P�'`�y�yDOl̙'v��;��(wp�p��c6�����sК�sZ�a����;-��M*�vj35b���s.����[�wt�t�Q��>dEN�ef�Fp ,|@f(�����)D�_^��&�]}M�w�by�x��˰%Tʌr�cys�$ _L
��W��4ܻc{��ֽ�6�����F��U�_��.Q�?D�L,��1:�����8`ON��y��)��<��j�r'�0���ro;yc!����!7h��Y2w�"��������`O��T�p5�j@�hw0��80����҅C�E��^g������6�W�%��1Qoa9"4gɹ=�PK�M�Ֆ�c��4t8}je�ݗ1���&��qy��gL�#��8������8鷲�[mAil�԰g�2}��8���1hl\!���-�Z��k��;�1�x���~}�QN_� b�Y2�`Ea�{74���YG�U�VۛѼ��,���n�Y�����64���(���Yt�O��Iv���b����'���|��H��5ߥV7t6Z[��>OLKF�Au�y�CB����ϣŏJA&��/Nr����^��9��̍�V�05��� K� OP�BM!5ʙs�(�:l��ܥ2��G������҉�j˟G�<f��ȴM��HGz̳����@���7�ʁ�\�f%6"M�����.�z���b���An��ڐM��Ӗ�i�E�Y��-�g��se��]�8Uv	7�=^�nj���0����B�c�^��C���U��R��`���Z<�w�y]��:DР'a��OZn��ʻǈ��ƻ��
~��R
P*P ��2zǽ}^�=�e+�D����a��9
��0	��	O��VW�0f4]n�`!��U�P׺<,�Z��6a�Y�����+mR�zS��m�*�x�1.�2*(��Р�"�����oH��ۣ����J(�"I��lO�p8�Yެi��#�(�k�ӻ�j�����P*E�d�kof�<�������TWow3�!�Ε@2��v>xs��&�Q,�ӟ�u������ϑA�W�yL&ә��[��ں�Vv�,���s��v��<]{ׇ�e����������Ӭ[e)��`ʭm� �ڥ�kk��[��Li���S�Ě4�Ѝ;��k��^~�$�`�W�I�=q��B����c��O]k-ֽ�}<&V��Ed�vǲ���'�O�A�K&�Iy��4�Q�|��$=��e̔g=�s�Yq&��rhg�t�*�Z[C��}� �Q�
�:�:!?�0�0��j�` sT�˖�FC^���6����wʙ*�][?��W�^1�<	[`�7;�+�K{�hO��yo&ǲu=���ƓY:�u�5șrT	i�\��{�ш�zo{��z���y79pI�r��?D[֦�����|���������������ŵ������������TKڊF��rl�=�a�kdWl��o7�k��o3��'�w;@�I��nH�u�|0�h�6Y_�y��:|4��\�f۫+�Ӳ��3L׉���+. �J�ל�b�w#���#��'{9�,������
dɂ�TG�h��}y��H�+��h��\.\øH��$)��\����e�K�Fv�)l�]7���@ܻ����bm��ďv'�5`'Q����qoZ��Z�j��)<��[Ԑ���û[Eb�|U8��ʞ�M$��2>z{P��H�34�wT��:�����+'��u{S�N�;R@Z�j�T�A�а9��q]z�;M�5&/"���˔�nI�^��_%���Er]l��1����FWwW}PɡiU�S��ê���mm���<���S����������>�-��p��5܈�gT4�U~�2���͔F��Vfc�0��1e����i�w�\�9����us��z�x�羷��rb�Ӟ�<��6�����3tg@ef�A���:����V���sp���_����oԟ��&�����-�:!�儍��&{��g|�w=���n���Op�����$�k�r�Aώ�q2$Y���v�#�'���F�!#(���;�H�:���vq�U����)����^��Q���R��K/�6W��ޏ�Dܙ���C4�*#�s������0.ƣ��Y�������������35^w	��$#Ǫ�)@�O�c����20��P��k��w����5�d6��9�,WI�#~�������n���s*�R0T��U�TV��k�G1�w�唬
}���(���=����~�O�q�$�aAe3�GyGo�S��e��픩[œp�i�b]D��GsRK�n�:p%X>w�{)�J�<�\�p	���K��{8��8{ɒ��I\�����h�=޾��XNc��}"����|{��}�訢v�P�%����Ϩ�5��2H{���Ct��d��ɂO�UΨ���<�l6DL�i��A��L��%����sx�w�v<b�ԃ��'X�Kt_�4vv�]�k�v>̘�ԣ4�Ud	����%�p�v�l��{w�xvX|.��ɓ���Ԍ3ۻ�kƞ�nwv���~�N�ǯ��I�m]�%B��'����.����Pخ^�E0]��`��ޯ6b�i^��-�KN�.�����d:,�M���)�8��ON�Tr~��a2��7�Q�B��3��tw���ٞ��'px�R+������곒8�}�9�<a�]�&s��ASM��s^[6(ϕo9e�˻{�/aTk~�L��)��:�.*ӛRm��d��:��N��\9Ifҍs��1I��a�t���;;��R�d� �[��z��x�������zu|�u��R]���I����89z��u����Y�A[ϯt<��ŻY�&ڧu�}z����U����=��ݽ���jҘJ��b�E)jrR�Oɑ	��H�d�Ī���̀�M�ۼ�ۿc���vRPi��،�?��m����70i�n�v��|��Ƈ���fcq��X�ZzG�(ηm�$�k��6�;���	�Q�J�187q�O�X-���4�7[��1&�0���M��F���u�c[�C%�)AP- �wv)3�w ��4F����ְmh*����u���3�.#���l�rl���[:�8w�`�5�-j.��jw����UF�3h�l�b-��G@F<��k|˪1�&����nγ���5I�ضu�f��Pf3�N �����X�b5Z�b���X�lpCN���n �1�3e�6��Ōk�<]4Z;��n�wT���cWgmؘ�U]�óX��1��W�g�7��TTDX�F����kD�i��k1Ӯ�l�f�ٸ�v�X�h�F�	���ح��=�}��4UM5�'�ǝ���h�b��W���j�:�[RV�F3���:N/6O��؀�`�
h��b)�$֍8�*�^X���:5T�5�b��huli�"A)2$�ĻcMy%����Oyͺ��Z�ݼ��c[�(s����#E�0gIƌ�,�[���9����P�����vvX;j���+�x|5�������-��E@����
ҀR-
��
�9��l�� {r��B�_Z��<�>z�r��vy�=yf���]}e��t=��@�폭䲲8q��f#WE����&�,��S�P�P����SƇW�Ã\�u#"�/`F Uk��'{��_�g.m������|<�8XX�L|�����4/Z��}�����]yCKX�|�P��4��7u�.���֧jE�@��!@[�0S�X�8�Mw���'��|���!8};v���Y���q��j����nb����L6�pU�jsΗ��@LMP,�����g�@v���-N�]J�;��z�b�oP��`�����6���Z>y�V���u��c������p)�ڦ/�En�uv�8�K�?��]��͉��nt������õ�w~�i �{HC����c�=j�*8p���F���w�Ɂ2кitzbC��2��gB��qM�:�z*��2���8^��3,�ƽ�L$�ۋS.�ˣ��fତ�˞ϟ��e� lj���;�2籊)?7��C*�\��v�vd�����s�lܗ"U� v�E����Y�!w�-I3���Dl�ش���o~7����Qt{�v���u޳��P���&���R��܉�\�c��w]��u�󷅙�%�|]\��ث�f���>N �9&��&y�5^�畍��]�E��;ԮE@��̶�_^~���%��w=2�uB�r��&�V�=�U����� bY�� 3B
�KBBB4P��B@�*3�����tOY�~���&�X�z��Co��
E�HI4���gzU)��kf�p \�'���v�k���A�r*�:�I���S}A)�R7^��9���͖��cL:e������8�lg���=���t�S͕!�_L($�];�T�G�
��N#�Z����_M���'4L�dc��Cj��l��X���<���O89Jy�8��K<�y��z}`%a��-P;b�c�/'z�Ӵz8�h�5�LBt�&zS��E�
�Re�m!q����_�˟�;���q�z�0�昛�eկj 硓���q�-���]��|���6���X��{�
�H/�T�;��cA%���[zߋ�3'�ta\�r �BpKau��!�����}o���ɟ�u��o�kw�p��+��y�l~��#�\��5���b��Y���;�_�:��@�需Y7U瘱$Ij*��U�G���u�{���ngV�G�o3S#��,��S�YuAK�5�\Ј���&e]m\�3ƳEή�"#`�aq�Tюq0���1��j�؎i��X�=�0�D�����dٷ�x�����8������d�Q���Ղ�%*��«v�o����oIX)����*��*d�L��}��n>ߘ=�jBlj�3/:I�\�����w,�g��;��7*-�S7R��(]�Q��Z1[�ؚʬp��\��V��G����cj9��� ~��ċB4-)2	J� ��@��J)JH*4 D�H�!HD �)2��@��h��.��_�d�E6Ϛ�H�£Jg����vs"�y�Z^�x�q�9���̬�;C�Bc^�[�κ{עo� �7�.F:F�5�Pn[ʌ����K�jW� �UM��:l��x�����*���������/�Dڦ��=�]�$��R�Y�&͗UqF]�R9�Rm`5f�J/'+9p���d����ŝ��i.v��>-�=�B��Z^�)]�d�цu��&��g���0�H�%{3{�U��Bnr�u��عH���}�
�c�p.�n�-]c�.n ��+:��7�[�ST7��hqGܤc���_l�}Ry�?D�L-*������:�)�\
��6�m�7a�!ۓ>0$�v�7h�	�Y2F�\1�%;'�}dG77�)ֽ�N/�s5��|My�p�<.��R�l8
M���Zy�_��X�����bDo�U����|e���Wes��_+,ڦ�J�.z=��P�'c�,A^�:^#H�%��6�bCR������@nQ�Pً^�j.�n�x���c� 8��#��9�����>����@�-���C���Ѿ.�n>v��Y5(�t,�혙�nYV�X2�\�L��א�+�ꊅ����y�*�}���"��&�'gk�)�7gZR�bHzk���j�{��틛O<�}���3�qH o�����'dWD���ܥv���^I�a�~��bQ�F� @�hF�I�)���hJ�P)hE�� (I�B$`A�� 0bX Z�7/�\�ΫWq����MD�I�����.�W����E˷Ks� �䵎���-� ��D�n<e�fkqn��R�K�r�tz�^c�kH��%�	��c����Tק�\�?5�\��d���!�{�t�GgV���EIA�1M��Ll3y'_�;c�O��:K���������>S4����I����{�0�v�=���tt��;�n��2}�ƀ�g�t7Y;�ݠ�w�#�ɂ�ޝ��xM �W/Tz6��a�� ��_��#圢Zg��U�e���qY���K),TI�O߳����CjE ��XN>�hC����2�1�j����WJ���!/�Z{� j��/�O�w��>�R���ZE�{�S\�U���1x�)��%sM��ha>��"y���Ї�yʑm���ܚ���37iȅ��mSϮjA����:d�-D�m�R�۳�'Z�b�1-"�7( �`|M���˽ٸu�	~�uLSnHU�.�t`�O �烎wE'\��)9�Ȧ�Joٮ�Oȡd��OJ���]f�y�]�,]��<�kT��ɷA�o��a� ��2��*q9����>-}ɘ�W>J��/��tp��j��T|o���Z�y��KZ5 �~����_5����#��±DN�r�m��^Mh������&�&o���]�S�j6)ݛ�1�j�|e�Cݣ��kd�d�|Oj�M��;�!;(�W�>E���D���x��.DIF
r��� >bİf$%��Q�hU� �V	�Q�X (�	�
�h@�iZiB`
U"P�`Dv����]����gEc����|R/�d�����, ���]�cK��jWf![�.����5^o=!�P��)?j29���X��!��}^h�퀮� �z�74��&)O.M��������N˒��ZYI>���c�[g��Z����EaZFx㭡>�q�H.s�'f骍�뷨&_�
�)�ٝ"�����䴧H�e��g�4Se�o"���� F^nL���ke��}�ow̅����_��S�<��4.�r�a�vy�=,��]%��$a���=�W2��u²6����G�'J	�6�P�����y�I�L���I�hFE4���R���E�i��<-z�����d]��X��A��&݊�H�+@tqƐ���v̍���3�y,4�Gu)ڍ���Ĭ�<L{�+1�1UY(؇^Q����s��h�Z��9 T.,EoM�^��X�p����Z� �QE�	�z��U��iKo��;�es�^S��.�%<��R��pO�J���*c���2H�b�vf_[ZR�b/���ӏ�P���6�t=��V��׮��<RY9�Xy|�������&f�h�$>�_���n�ɦd���ӚfN�(Ⱥ���fWj[���� #�k����1�[��!�������?A�eo�@�o"&�6r���7�%e�}�]7R�	�K	��h*v�"_`��w�ɠ�0��`K0�
P��iX�i�&@�B�)�)P��� $0 �0iy��Q��a	ٽz��c�jp>�����ױ��=������JY�} [� u�:0l��h����==���ʈ��`���K�>\�0Z�c�gJ��Z�/���NS�X�dgNf�R�1�l5��[S~�����s�~�CP��R�����JlkИ��{=�����v��D�uf�ڲ�'�,N�9�+}�jH��l�TZ��,�u� R�]��� ��i���S��-Irp�M�N�I~J<���b��Ӌ����^���SH���	C-YWsrnfj�M*�7Xٗݭ�"z���̴�`�:�QL��S�n������|�G4��uy���m�ǘ
�R�6��%��4h�4�RU<�;)�˛c[yA�У�yc�-����l23d.��B�gؗ��p���[�<�2(�Q��aa#%�c� �6��5���ȇGٹۥybq䅒��g��<k�P���Pnc���צ�w)2�8�T'��k!03%���z�-� 
�n�P�H�Ä́��^|�"!�˨K����X�m�I��@����ZMgsi�AjF��@�K���1���.�0V�&�.�M��ɋ�;�6D��ZaK2�c����l�O�ڱ��0���,��v9Z݈��?Z�\���Q��#u֎b����'�1��+&�Z:��K��S06�qB�u�E|�0�fd�ZE�T�@��EbE�)J��	T�b(
� g��~o�Ǿ����w˭"�=�}�G4]x�SkP�cAr���N#��O"6<D�Zo�la������RjZZUҠ9��&�=8�U�Ƽ�Fz��w�������������K�>����~���q �Xke��5���k��0��"��-l����^
�ţ�l�9Q���Q��⍪��u�J�9(��MG��=��m{�T1�FF�Z�%��0�8G�`}�A����u>fs5n��<�V�])�/����������T�~�c��8/`���T |��x�a�\���
�UѼ�Y3��(3|;�i�R�Fã~��@W�Vi22z�#�����F�;�7���v�=��-Z���n�cޭ0U�)� �Ia&͛]��
#�_�¿P)��p�Ǹ.�¢�2s*���^�\U+ֵ>R���uE26�����勿b�mAk��%��Tl��#ó��ǢZ�;n�`�3�A�x-�#��)��UL���M��m�Fd��g��UU9i��-��A�V���eS ��r,��;�ϯ�%�	T���%V�~�I�������㇆<��G*���K��ˎ4��g����F�����|R�/���N>5Q��H�g� 7�+�_���k=��^�`�DCn�eǺ"�e�����A�6[��Vm��:-��u|5tzu�����Ob�0+&K��{s��b���[9�̗V�b:���@�(� �hT�Y&�B%���JAhJB	R�
�D�)R �H�l߳�;��kU(�!fA����[F廆"��&��>#N�P��))��Q~`'�+s�����V�g�B�A���\_PZ����;rI7�[k���λ�ק�orp��$tz���d�V�3��/�Z�q��k��d�I�n-oc�ü����q!�^��B}, DBm멖��Hn�YZ�Ԗ{�΋nq����-l����=,�0��1��c=
HXj���N4]�}����@��ڷ�i}�;O,42eSʭ��$���ҪT�3�|7�*�n�@��� 1u�J�*�9K�
��0��ؽz���9-㐤Z�P�0����mO^�}�S^�����+[y���÷^�j�p���um�м[<����E�k�=�3�9���{$���܊q���OAQن��b�vנ��S.���dB`$ǭ��B�ykD�@����d���u���®;�lT�ŚP�(a0j�NԿ���,�Q�b�S��G���{=T�>�p5�錶`��Q�|���-3/W����ƃ��z	a�޵!H�g��R=��:�,!�J-G�ű��O��ҿ��j_�������~>A7��hԂ9�:��Xfi�����{^�zV��y+�/g�hU��uq�9��@�S���a�I��@Xl�
2��\�p�Vv<��#�N<P�p�g_F�:�z�<�8���O�tq�L��՘/��;��1��IK��)/�h,_��~�D� �!B�(D�RHB,�(D P�%�!��(9�wdo��b�H�I쏎w�Zô��e�/Bf�Ԯi�ƭ�}�7�T��&�;���Z��a��T��WXO�W�0)��!0;����g�\ȕ���2c�Q,�������ֻ�;;Q4�=v��!qY9�ѱ~m��Q��^FS�;��PE��hGD�p/�):���)9���~���-bY9Ǟ����e�]�Pn����*]��84Q�� >�<���|�͈�h��n�=�;��^Nu�?6��y[��{R(�R���r���jg�>Y =L5l���;bd�4Y��ꊽ6��T[�OݡLy�z�r�ܝ�ؖ�P/�48�kـ���ߪ�_���:�x�ᘢo�k��K x˴�t�Wu�.�%4��zZ��������XE�^v�;��ؼ�6�dL,Y9��U�ǆ�rfs�,�����}�e�iOi,��{B��Ͷ�F��s�󼶫�������{�� C �XH����}./��dU^r�O��lsrz:}IW5.�P»)�#�\���/剑m�{%����b���D!�b�='}07�Jq��?���h�=��Ŵ)罙��Y0*4葎��/([
5O�W�ݯ�2��^�`�9�h���N�r�_�2�+�nt�KSa>�Xπ��P{:	��5�4-�&%�5J)��j�j��Ҕ��]�
�[�\xd�Yӊ� �o��7Kx��ڂ_������y���
~��� �*R�*R ��@�� R�K 	 3Y���?mWb��<]V���5t���{yH�F2�"p����q�z�H�k�����+���*�|.aQ7��o/lG[�`�0�36\1�_��}�'�8Eb�Ux��}����B����j\�w������k�^ݸ9=�R;��z��eL�{*T�ˬ�@15��;}���u��M�Ke�
!5�yzl;e�49���^(P��4�x}&9U;?(�u�����X6�ӆ�֛���A�I�e�Fh�K�8��pN�ԻȽ�a�!��)��}S�7������t�m�O�����/�Ϛc�:|O�8�>��3�p2�Q��"�y��J��΃(p)<󡭛b��y{���e+l3;�Z�/3����d_\;�.��+7eu&�s�!]���ʚ@�Wƍ]�Ǖ�v#KS\<Z֭t7L�s�p��qY*X[I��k�L�i Y��P�@q>��^��g7��7_�
KPu2���S�M����լ�c�������
wzp�}�V�]�UL��P���;�.� ��:B��l�<���s�^[��l�u��#:s%�ҥc0,�L�MM-����CkkkkkCkkkkkKkkk&�ֆ�߳���*�QX�`�0?L���/6䱕5uٿ��c���mPȊ�������x&�u'���7�VEth���C�
��>A�'JSyCՏ9Q��Gr�c��\����5o6%�VɱW5������pBTn�Ur�c:�����ʧ{�eP	�w��ڽ�}��nJ@�]5���A��g����/�R֝[yr�+�v����`v��צ�מ�PN��� �:��WpY��QhJH��旳�U����t�Ü�ݶT��c:!{�Ou䖪D�Yp5m��c��:[ō8�p����.\�x�����]eL���l�bF���	C�xY�լ�b�	w�%nVu�t1�ّu�ݐWf�	�&�{P�5υ��9�.=����z�3�{�y��d����&��Y�>�-�d�_��inG�����zÐg�])�wn�d7�r�ε(�T�m�eG`��ϒ"�!1�j��Obk��Ὕ�3)��i5*���^��A�\���x0��n�Xd�ȷ��ճK�0�^��cO�)b���h쇘�ݹ힠����#��h;�򮰕�^q�G)�#��-��k��y�z��F�7/GF1�l�ϵ����]gJ�񗋎�ޓ��kr�z�5�
����'H���r���`Ѽprq�S��)Φ^�o6��25O�[�9��O\z\��-��>�TWҜ;&��/q��# �o1�B��OM:��a!˽��F*�n0MS49')s���T�J>�+�<�C�g�ܼ|F�1�\T�bd�������S~cu\j�ul�Un(.�:����zE�ʛ1 l���N�/�l�0����Am��q�^���lԻ�9�9H���T���l����9W/������xr�*�讨!"o �E�S���F���W�F=���-Ee���^*n�$-]t���Z���ܥ�����LQF��|�r���Ԅ,ŋ��һ.�4>�ɫ�K���)s���95�zu�\ �I�7Pr�j�O����we��j�M(��F�͡K8n�t�����ғ]�ps���˩]�ȳ�ٍ΀���ʺl*�T��z��<����I�}��h�}2,R>{6�$�4�k�	V�0���6�/�!)��7�_m���Y�o�roo�hW�+'M����^g>��@� �5�*)Ip<"Y�����cJ�>͜Ugp8�/�78��oj!w�{�G�7Ls�z�I5OsKٳA]���ÏI;�g3�a�9�t�Rmq�dw�����f�	\�7�u��uå@�,^WK��1�̹t��`MզjCb���ný�Y�4p�K2�$�
�8'��a�D���~{�{ ��3ݢ�;���h~����R*����
�);N��ѓ��Q�K���5�;vT�����(�q,2'�Z(A ���|��:��TR�CAEDt�ѻ>GO�3v$��k�I��^A���4|�(�cV��EU4iLT���_S�������?1MR�h5^N��͢����)4�e��H����I1^ڢ&��y���Y��D~'MW�8��N��X��'W��pS�11%��鵊����Y��/0�Z������PTRl��5�DDm��j�;Pto0o-�*B�CF�("j*�6�bk�b�$�i��~�)"�TR�P��qTE3����)���%QM?!�c��$�%���(bڟ.�]$I����d�g~1��$F,E4�|�*��ʴ4]�}o�H|٤�/��rSQQU堻���6�%v5iLI��DS5ELCK1Oy�yH�K��Z�ez�/]oV<��g,�:��{�=����"�o��;�ܥ2y��x�1�,�5X8t�C�T�:�(�J<��F�3X�~ �?%( �+H!@@!0b`�`;�
o�=P���՛�/�b��d<�a����b��T�]�����k���~��e�M�%kj���џEʥ�X{���q�yM��hȮ�2i�Jy�%��&F��Y�t?�/*�3t(��<3Ωa��:A=�IM��l��LD?����c�gH��@\<vdvKHaf��grw�QN��w��O�l�5ȋ���1+�%���m�̼��|3;V�HL�Caʃ�]�\��M�\��n$j1�dsE��mb^�˒�C�!d���`�/]I�)(ICŞ������E#4ɶ�'�ZGGD�q�������[���ʃ��s�w�e���م~��6J�Q_d�!�G�c�b�G��(*=��Í��mN��24	���U�jsr��Jn<�CQ�#��fV��^��o�ݪ rW���4]�z�-� Q���ϼ.�>�s�k��S/S[qww��VJ��)��zS���3���6�|�Jw�`^,=/u~�-��rQ~�C��\'d��ٻU���"e�� �ﮙth�g,�k�Ɏ�U(q�aO&�1jdے#і*��8ޜ��J�b9�Fp�5Q&��m6T�ol����:��������&���P�.�V>v*��p���D�骨��V��ou�����ڽ{���R��.��Sɾ:y���̖zx��T;���y=��U�hWL�N3�;�~�� `F�P�� ��G��ƘZ���7�"'�-)�1gS-άiC?�f$_ߌ'C�h��}��硫�ҟwVH��"�{�}�6Yx��i:i���'��4�.����U勰0&O6�^���	M�S��N]t��\Nz��\���[ �����@,+�e2�	U2.p.�n�Sl3�Fd�F�J�p|�*���S/�����B7"q�M��v@Q�%2�/|�]0��Sw`J��7r�kU�L�m�f�k�n���E��:�Q�b��F�#�c�&��	�Y2��.84��1C5���hj�sX��Ψ~Sn2�Ҙ؛N�渿��Z���W�Xl��@NgWV8�1Iov��d��{"��;�*ώ8�5���%��l*�AtcsQ~vx�,@+؇H��D3�s��}o��φͱ��G1�\�����SR��,q�J4���y���9c]�9�q�@^�􍤽7M7{���u��R�]5K�sH�3&tnoT�v~;i����>��¥�[���X��^��U�!Nϕ9�N�K�㯭��Ҍ��->Y0��,}����jz���Ć�L�$�h7����@Y4�>�t���읯��[�g�z�}���<#Bxz?!�����# [2��;�r^W��߾�������f��Dެ�sze��T�ь�9Q�{.�~�ċ1f�ń�N�Yf��\¡[YP\��Y����r>�����i+i�>�pvEY�[	�r��8�Bp�DXS���v$'.��~f`	�ff`  �>Ȝ����L�B&�]a�O澻� c���d %��y_,�q��r�l1���]�w�jc�z�'���=��L�7EHek�(�I�d�۱0Z}3�Z��'!�v�����m籸��Q]��*b׫�ې݉	���{<�_�M�d�*��J8�g������Jcj6��J�ɝ�֬[h{���pM3R~�2�O�[H~U0�=�N��&&���)�/o���j'_i�{w��Bj=��6�tntת�2|��K6��&�z���ǃ�i��v��X�3�S�&��}���-�W
�(��EЍ�au0<������\��2c�Q,�,Y@SjW8�KA�0,�P�PcL�5��_��sd��J�Aʁr�R5,<��ћ ϣ�h��Bu�F(��vi�46��ưX46B׊��a�~C�潵�g�+M��������+�4w ���="�O?��M�bd)
����X��癦�ۡ�-9:��ᓌ5�s=Qc�t1�zJi���O�.9��F��!�kf�q��k�`���M~�.Qn����Tx���`4�B[@�،pd0p*f���:)vlD<\tU��|��zL��~�3��:M��}���S� Ūb��z�]�5��mlb��٣��j#/(�Yc�>>xV��t�0C.��=c��h�Q��7F��e��詬Gz��.Kyp�3-y����͘�$)URJ3��R�3f�wI^wM��8(���ɫ�;`8MKP&�A?�tGF���vP�
���Y������]I�Jn�Rm����a�K�vD�*`G>�P%��:_{.SJ{I�d��s>G�4�aU. �����~�n����)��=�В4ݟX �������oz��"�w*$e���S��g�aȍ��19$�L�g�+�y�6����NtK�~*
�[L�	!0}Nԥ�E�������*��	lsN��ʭ��w��፸��UX��	i�D.�n
�Hly��p�k�[��(��q	���Wd�!�ǘ�?NP��m�MϤdtD���-S��#��N������{��}��%e?�Z'r�I��$��0̆v��Y���CwA47z��5 ��)mP�qA����H��z��j���'U��
L�l���0?�\����	�>�k|ޘEk�m��Xl��m߷����	�=��"��,����B�B��8ػ�UB�Š�ln�x4��KfN5\�ȇ�[o�x�V,wt;�m36�Ŵ������w��js�wT�{Ѓ(p����W���r�����a�6=%E�.}i�t�{����)R��K�W/u�nfaA�y0��V��9�+��Ӟ��N�d�H ���ڇx�7È1�!�o�,�;�����(����\y����{�����lg���ūV��C�W����MFʰ^�jNf�|��O�]={�_��|�����	kU}��ub#�z��AU���n�g��d8GV�M?Er��/�zick+PYs����P��Nf�����ӑ#5��H��Ϟ�����88�cQU��-W.�~��ҁ�Ť����$���S�M�z�k2��ﶞ��!�A�-���_����M���m/�je42A`3n���
ua�S.~������R9CnL�Lq���a�C �9�ݍ5�R��t�����c�F<��0�¼MJb�������j�Ӕv��i�Ϲ���<.�B�,��T���+ǲ1��,/�Y�����I��U�8�U6�`E����W��&۳���!���a�X�p��]����C�-539�P=�^���Q�Z*�`�
�m�gYz����OAdw8�	Ia!i�XYi#�w� �庝�yw�SOa���G:�뼽��\�I��{Ȭ�����3�`��TW,nD����^�����a%0�RJ��ܙ�#à��i��\I~X�ҝ���BGs٩΍/�Dq��<�!���W 5���O$c�N�UxN���n���6�{�@�D�???X�yX�e׭�\�P#4�\i�����+*�<�����S�Һ�n�,�/O	αu@�i�nPМ��،�;�fѰyr����i֚���{N�oc�9��D�>�q�����Q���������d��N�R05����iS��Ɂ⮋v�(�C;١W1�F6�v7��Jx���}Q2�D{[͝*T�q^��?�1lQZ��ڦ'��k���
>'c;6�f�̮���� �˦�4��h�Ζ��u�<~!���1R��������V��-�t�R�_'w�/o�w>�Q|1B��z�����u'�0�x���=��6�%�5&��i����^�ő�q[bEU65�BKEZ�[i+�
�Սx0�{��"E��G� ᠅���T3$�G�[�/�0����ԋ��4���Ʊܥ����~����U勼[Q�G�5>�.��S}Ϸz�o).����C�v�2h���k�:$��wL�[�J��s�joo��b���E�u��룂�;Dmvp����u?�kz`��G C��V�C�t�F�<��K���Jn�{��z!�����*l@j���$�C�q^��`Oz�eL&�����p�L�q�	��\=��v�O�����|W����~k�n��k���P<����ۡ�9v���qm
x<Z�Y6��|�������n^ퟚ~��کBy�E��8��삤��v�R�^8i7�ÆfFm���P��ɶ.���aW�wM��1�����n�[����d�V"�ی9/���#*?�&vu�:곆���t	�q��Z~���Wgw�}ԋ���[:�o#�q��(!�	ဒP������ܹrOX�a_[z��tГ�{_�:�\q���{O�� �;�6@�!�b,!>�/1�vxZ��#��U|����M4�S,����vR�@�Q^J9�屯��oa�G'\�	�G
��N�;*9��/�wg/����U�)��"��q�MCt�Oˠ�YYC��Lk`$\��{��'fE���Hݺ`�Т4��ܐ��ϔ�:���򻌁��� '��eqΑ����	�jXc�p�M��mCC��hGC�8�y��u��${�6���J�c�̎`ѝ��zbo%D��n:��K�쑃���+�ADbH��d�??`�d�dg�{����^�a���gpb��VڎX�2�m�v3�`2x�C{�^AH�)�,0�4,��@Nb<W�\�ܻ��yGkI��x�X�o�l���ٙ�3I�i���2�1�j�����q�o�V��?W�DW+�D��ͻ$��V���'�GE�*�i�O�*1z	\�e��v�."6;<p��=jӽ5f��]�ۧ+=C.fE5И�njGj~��~�0>z��5�+*�ϭ��y�O.�Ν=c('��a�է�	�D�Ȼ˰z��'�}|��F�j{;�<��<,��mJ#�PYwx��m��wSm�����`#������<���E��ٰ;ju�<&3�2L�fh�������J#�wo��� WB�_+����}��"x��[uSw�x`>��e�&#��eݫzg��g6�;���p$�
��h�ܛ���彍�JE6֢�V�͋5(����tl�}	����K�����S!wZGm�[��z�Z��ZruH��Z�a�D��������`SW��a�ހt���k��U07�.�{c\�2���:�C	���u�u)��Khu�ʆz����E�#ge�n�>7=5}���:i�K�{���	�7+�`j3�F0C�l�We��<��6�//#�	u��9���Լ"��y/�`G?E��8�A��Ҝ��7G�K�W�v-n[�uŌ[շ���� ߛω#�F�ya���S
5{�
z盝4.��Ra�k:s�ǜS;
_����٥+^g�g�c�)�m�)d[�V>�'�\\��}��='/oǶVږ]��;��b׽����ea7H�����s�+��D.&ܬԌ+�q���9�L�C�<��WV�0b���/�}kѾ��X-��[ے8/N��a���a�D�~B)�yI�FG1�Q���5��V���LW�0�ޣ�*t���MT��S;X� �[aXU&n�����w�����Β�Y�p&����ɽ��CۃrH�w����]!������b�t�YL�F���u�+v`*N�|:���	�'���d��������G�LA�2�I�V�S�5�` �x�~������N|��pM�Cvd���F�O|�s�@���<iy�_.--����R� ��^zA�]Y�[��
.�ё%J`���^�z;r��,H�ya4������+lkC���ͩwƾ��j/լ��ϒ�1Q+��*��G���إkE%I{t����y̽�7D����n��a���a7�5��|Ix7�)Ә�uk������H��TFE�ej�������~�=�\�m�A5�t�d��g�@�u�!�(W\����'����"?�Ѯ��x�?��8qDo[u̵���u�|�MScjt�\�P|޴�6����)�qU�=�,)��t��Lw�4Y���}�����7�,���ř
��֭����T��ڕ$�m
ǚW�6�ml�6��	X�����ln����m��4�Z�6]/D۠�Ӓh`3@�Ry��钝7��M�.S�zW]������3M�w!��nU+���ֲ�Æ�|�����E�{�S�g�AVM� ���_��ή*����L�bF���uvB�A�o�q	��;��PN�va?�q㼦�j�^�#o��ж4�j��}�D���]���+�S��N�]�A��Ql`ØuT�m��j��\B\w�A�[�)�Q-���#c&b�fx�R�+�ǻ�wr���/!hɣ�����XW����?������ s5t����tn9<F�cۋ�Ğ��ؠ����i��ǩ�}�}���GK���34��,���}�]Dc�Xdj�S�����gf�i��~���ӷc���}]���{�'��!ho%j\vxoO'��������}��b��Ä́��H%ן5s��O%����P��]�M�f0�Ho�Rt�����X;BR�"��sE��`0�s�\�r �-�y��Q�J������ձ�Zi���s�L.h�������B]���<^��Igמ�� r��v�A�u��\PQ�u�t��C�<?l	�T">ZD������_m�����F�`k7j�X�X'��ٛ}���{��uAK�^
�Hwlv7��3�A�߼�q�!�Z�>do%��.�{�0LL9�8���V��^�X�ތM4|�tkW��`8�D��?���k��bƮ��6T����;Q��γ��[<�*Gs�9�pć�l�i�#]#|S��g)�2�蕤��Z^�Sflՠ�Q�k��n�4�M)Ƽ�Ь{��py&f�lH�2t_���ȿG����rr�n�S�M$�wY�Z���
�іS�5��:�W�r��
3�[#�M�*�����s13�455�56��3������6������������474�73�)Ļ��~���*�a-�K�`�{�n����V}�����sF�iÃ���	�{���%�XN*��g������lݞ�5�I��w�ʛ��&�x��^��-��#]R��;�K����j���Ю�����w`�DS�}9�}��aن�G�����Q�y���ݻ��gHp�&S-ht/��k9�3����vj�Rw3���O�O.\ޢλDv���؇c�m����LU1Y6ct3t��2�^�z-6��/E�p�2_?x!�_\O+�����x��-�O\��W��da�`�R�g��L����4����\�!��vb<��`o��;wV;W7K ��Q!�R��sjV�)�J�v�]왖��Ι�`��(�r�]=������S1��u��=�MZ,�_�{�^v��J���-��u�mcj`�Ȓ�lI�������/�>�.,W�t���\q�46�K�6�d�
�Z�@�
�{�M�~�<�/�p�j^�-ɹ�=��Fy�),Rhg7�r��ϡ�d���F)���>W������h|��sxc���s��7��
�z��0D쥳q�t�ܖN�3�%^ a5�(�T��y�v�L7��{Ue���!��sY�~S����<Ҟ���z|��p��:���k�)J�WIP=C����.�^)z���!`oj���s��^��������u�p��Q�$�ՠ�bܻ���4e�^��bhZ���X�X>g-9����(�'=�{	��*�l���)h���m�[��MM�h�A�����DN;ϱ>n�X4���r�0+!Z�Q�;lc��n5���^}s�p���L\��s�4R�O�J���W�5O��#�<k�j36]=쩒,�f���Ã��G�p��b�����b>:�<�� 79=��󜙿_Q*1gP�M����|���p�(�MK�k(���;�P�y�:C�fCך��j���d��Ǎ��2�_%��MMr���W�Q{{�ìS5Js,���y5���e��5��m�hً\pgD�'��H�/��]���B�B;k�����Q'0��+��c�^�y&n���<-���sX��{�R�Y��Eb#wOʅ���R�j
˻:RH�L�>A:��]��>y2i*� y���8��!������YG7BME�yٗ�%.�G?Lx���,�"�Fg���U��&�n��o�.�U��-�@�t��(���(T�/.��L���k�}/|�n��JE��[�XƤFof�9��1ӕ��J<nh�j_�IY�d{��N:OL9��U�<};���&��MBF=׹	)Pǈ=$��K��u
���yqQ������z���=m����Xv§���o/l���u!6rS��L�s3�w��3���y���vX��]>a#ٷ�k���e��I3�9&壎I-d�u�t[��n�tѝ�D��&"]��57�݊j�MS.�2��h$)��D,Ddl�d.PB�k�EAF3?�S���F�)C"RB���;U~;ϫ���2q��Ό����wqϐ�3�)~�w��uO�?$:��%����4y����m���h����ꖼڂ���:K���F���c�1�vꞻ��F!���6k�S4|�t�n��y�P�%Q�n΍&�F���Ƽڣ盠�&���v��w�������ǘ�|�a��@bT%���8�?<�#kI���&�;jJh��}A�i>�8���q���5#�A��h�R1���#mTPUF�;Q5M����<��;��I����y᮷n��)j���1ME�#���O��y��1W��xO���n�]y8���%5F��4RybJ*>��� ���<��7���(��Ӂ��|�?����3��;vY�)���^�L�v3xX2IDe��@Zj"�)�R�	ާu&�\��*�A����,@v�ͩB*��r&� ��L!]�R��i_�� �vJMg[��� ��w׾e��	fSjĪ�8����]�@�֪y����UB�{��Kƈz����я�T���;!��j�=��>���Tb��rr��Z�2ﰭ��ʢ߬ߤ��zhֶ�؄&h��8hN�Ռ|X�z���`��B�}�/=dㆍ�_��(G3���{�����b��%冄k�1��Nۮk�Z�4���z'�KJ]%��(-�3b/�O'�Q������э�@�:E���C¯ڷ�J)����N���wu�`�#)�m�����MKP9aBOǾ�������i��ω	s����,`�*���}��~�E@CWbr���B��gM5n�)�Ih�Y^v�&�Y���;�O���տ��e�a��y�x���_���r�cU�j|�>8�1��<��t6��<-΀��&�%U�T�w�߶���Z��'�'X??[�a���4
{����ގ������x
7��Oc��R�푂XtEr�\�
";�{0�B7�_���~0!
�8�ɍ'��{jr�u��y\�iI�#�8#ɢFvc�M\'�
�+
&M��6F-��31Z�Kp;|����]��e�z-�p����A�#3�z@d5Y�}���1����R^DUv���/ ���h�.[����ާA��wh�(��^�m���^&���z�28�n��[hq;�(�-Ø���5BXIF劭N^���͞�k�>lE�ѷSQ͹y>֌̗i�S��RCo�Ӫ�C�+�O^�y��WHNg�ăl�s/zY.���cc��zj<j�m�;�b���<�w��꠼D�7#=r��6a��n!d��e:u�dD!�N�^�>cϟT��"��LL�3.GRxV�}2j�K&�6`�9�Gd@y+_�-��ӽ�����ei��3���;\QD�qb�Hqw�Hא�b��9j~�J=nc���欼�;��h�L��|�^*)9��)����+6=����>�b췞Mބrm���P�3$�ZՅ��N��B�4�+^�'���P��6�X����]4c	)��1k����F�F>�v5�:m�ï(L�,�g�=wV�\"��QI�RTx��ʠSX; �6f�^.�K����=�B�>�Qx-3� ��s�ch���:�2�r0��٥�]<�>;E�̪��ҝ���S
d7�B�x\�/%��H�{N!�m���{��4���GZ�ndɗMy>Υwa�яU/NN���\ZF�ez�Ń<�^��%O�.�J��L[Rn��C�ffT������a�7՗�Z+�85-�� 3ej��O�974����7yT�cy@��l�μ���%����A3�l�eCAum�b��hTH�J$E��s
p�0`�k��J�з�߇抯>��ivo�Dhh#c��M���[�*u,�B�}\F��g�r^�>������Z׎�.�E�ΞĤ������ג��. ؄6�)�i��۲�?���М_������e�O��N�����K:Dm2�Z�1��*D'+yF�|�Pϑ��{�<t#�p�� t�m {�ks�C����CޜF������Q-�@��o���}��oeF^���F�kԇL��)�ϤnC>�E���#5.Ph�2=�0$������r��]c�o �&�_vD ��Dq��+�Ӵ��5�����^|�P�̹��vr��7czs]gN�Eo<����5�:�P��)�M�ycSKָƠ#.Gf�m�1ע�Ѻ�s����'�c�3���Xk�֊.+aފ�i�=�_V~���%��^
~�mB&+w:"0,V��m�����Z�/�=�9[��$ߩ�Ս�G�%��Ԛ��>#v�eև�f�1��n����ߜ�!&����%�la���n���[r·cMl�7��㠑IN�Z�����Ķ�֝��پ�N�>aIYT+�R�d)�)j��ӳ��:t�Ao�s���!mM��	q� T�7�)���s���!|raU)�7��ǧ��{�Z��"�K�ص�v�r�e�v2*��n[�aT<9fM#l#[��0f�鮝�ޜ�;�(��>jZK�F1ju?������~�%>D�V/_����c�ї��i����b�s�ʄ���>��P�	1�x~`�ߟ�7D�QL��S�2���z,��n�������7�/�_�<���Ǣ���˞|�7sͼ��_6M&	�LS�����*>�m��n�M����PJV�_.,�z��6��D�=Q��yW�S���&Y���'��80;��*ї�,1.�>��4��uK��Q"Ɂ�^���_���1	�z%��s�g�f/AG�סy-�T��.6�;�	�dw>5����r���w�<�t@WK������>~�%�{��ݝX��	���/-�%�=�U�ĢL[ז�0�3&̷s�Z��{.�C��Xטe>�8�7:;!吂�!�Z�s@2N�TkGGI�I�l�Ϯf`Ǟ��b �2a��f��R�ל
W���u�8�����F�l�Єm�����f�y�}��9X��7TGuQ�	dN�s>O��6emA-�5�],������E����5��)���2n�J���v
�ȿVG~���
�v۫rW$,_�ۺ�	��ke��mI�h��nOx��;=x�Kr�qm��śX�^X�ٿ=��+s�sZ�v��Ɋ\<�{�{xV�x����^z�4^���63�=�bѰ��{�#ք͢ı9(��F2�l/�����o8
ݝ�&���JĴ�o=�D���Uѭ_Pn��??H��1r�F���픳)Er�|��=-�Í+���\����*����X�G+�a#�G�k��ʏ"��������w�~�qX���Z��ٻ�-m��Jh�Rj��fM=���H��0� �L0ֿ����,Ь������oA��oF��:���&Gl԰�~�6�ܥ���[�k�U]	�c^�l>G޿|�^w\ص-0�P���I���9I�i/Dq����"y2[m���.�7qE9��=l+�~|���z2l��\G�n/����"�Y���r�]ц�z̩mz[���k����Q�l�3�ɜl�,)��=�������Y1�v˓ọKv�ʽ��:vC��N,:�E>:�O�k����J��J�a�:mx�	������N�m1뙎}��MA�SLZ%�3���0��	>W~3�PK���Gs�]t� 5$1�|1�����y�>#c)D��Ѷ�j�l$DBb��~�m�2Z��_�`�!���>�{~~0=��,�2���:��J-�(��n�Ѻ��p�^��4�c�n��v=����W�������5��d��?�*k��~�z�dŞ�����Cg�`�bu��C�4�=����t��6h�M2����hyЅ1���,��?��{�r����F|��7
���?�8�\,RC}G��9�`��֘Κj�ԭ1��[����C�m��2��)d�'r���A��
�rG �>��0�-� ����<�ʿb���`�}��7w�x?Y��fp�wDZ�[�;"4�O��4?6�;;����>�^��ױ�*G(��UT���C5Y�1���"�ހ��4P3/ʿ/; ��Τ�����0O�x�W�`�1	�:���Wn!Y1��qx�nj���;�	�G#D��N���OYΒfP�}�=vE�K�5y��Y;�ό�ŗ�5�,d��fK����ڤ�!��fөc�z7.���H����LZº�0`ر�Jx�!�
ipSĿ����v%�2�⊔ͯ^J�,�ŧ�T�2�t`vN��W�S�C�\Dg�nNByR)ZN���Ÿ�P#�%*&�N�U�^t ɫf���6\_t�Սmh�̜�T]2���Nl��{��1چ DO;5�PG�l���H���NؽT�:�EZ�t(����lsal�9�<Ҟ�ٸUiM�gԌ��F�&�_.�O(����d(ѻb�s���w�����e��dŽ�@-��.G�-��j�u��]��X^:
����<=k���{3��g'��<<�n��-�x�۸��ނ�%��0���&�Y����\��r�ו��o�ܜm�r�=ӫ�����<�|=����k�_L �=�,�4�����q8�a�޷{X=��!Y�Y��ҺWD�2�e�^����ne����y�Ft�;H�)�E��T_�E'��T	z���_�H����wh�����L�C��(K�)�2��ɫ��ªY�t��Q�F�i��R&4\{rVP��Ù�<����#_lP�!�ʄS�ޱPNR�b6�t�{��4��꽃rzX�o��2l��AfǬ�y;&�.�B�X�9N�'τC���^�M*uC>t	�w�#�b)�R���n���*�sG:6}@h�1�IN�P���=G_��/���c�c9Z3l江$�{�}�א�S@߃)�_���Α�F�u���D.&ܬԊ�=���,�����%���%[ $>����)��1s{C��m����2GDW!+�B���/tۘ�XWWLev��!����v�P��C��,�N{e�;+w��U�CT�䜕Px����s���l������ E���c>
e�b�/G|��w(�^>�B[��M�!��s�tvĉQ�8-X̓��7���m7)�M�Ca���_1�Wq����Jy��șN���AK��K廀g�$J{"^UPz��Is41̘��pe����c�U�>D�&��SΫN�IR=Z��w9n��*���_yndEl��U��S��LϾ\�.����`}��ީE@�N�S�ː�ܻh:*/cXˁْj����%ʦW���8�4��|��Cڧ���u�:�������͹�^�~��� ��5ߴ���4���y��F~l�t3�P����a,�[�q���������xp]��L�M߼$�j�)�q��O�5>��1�r��;�2��6��ש��ȱʷ\]�[P�E�;j��vSz�\aOW�ceSx��-P�nY�������锟���#w����j�F�������r����B�\��i	ޗǩrud�,�f����=���(U��<�K��{�)��g^t4�j坸>�,|x�Y�7��~�ρ�V_˃�z��?�1�^�o5�i��vw��ZZٮ���dY����p�)v��5�^#�B���yH��o�ў��W���Yʇ=�0���zH7j���d�X��խ49j)�0�~xy���1(��n�hYk�,�9T�*�(��b�ɗg!y@�|�.��m���BŸ�+pdS&M�����8|��>K�ԯMN�x��s�d�0�KF-�����x����{|�uy_��"������v�m7��p]�iɧ�*L��D�7�^�����7���:���i��O�<I��Ż�&ɋ7���S�E�P��n��<o�t//�;���\o���1�!	*>`�5�w���{\�q��5�fsu�1�X?�}��X�	I^�����UM�@��r�(�ʒ]Y�!'���U/�4�	�I�� P�����4ōD�)��3�=I��cZ��`2_���pԭN]wF��Q�F,L6���3.V],��#�r|������NHv.��_DNMD.}}��V���jBi�{9œ<Z��Bꂗ���]!ݱ��A�KO�9	���S�G��y�Xiʑ�f�oL���S���~Q6׉0HIV0j+|�!�]tD�,`Лتr[�F�ݐ��l ��W��6߷^e��_�ß6�"�Uc�y�YpL;a�<Kf&���Sj�%M�[֨���I���%Ƶ_�\�V��4�MZ�[h��cޭi��!�(�ᬧ9����]x���z"[Q��mL:�є�J�.'ŧǥV5�� 2~�b�e�������&a��q��ܹ���6
*���[���o�G)d����G|����^�/�EwL�Z�rZk��F��������6c�1Gbz����{�qVTyc�9��ۡ��[ml��Ɛ坭�\dC��s͕O���^����=���q���X,���:����8��X)y�.(�nI��孨r:�ݽpmʕ� ��rU���@��o>G܃�5w!L��'>+ޢ����ɾjƌX�O}x2C�-7�z���xVM�Nu$���؄��a���O;mvA"�����~���<��R���^���&u�^�O�lk�|h�]��OM˥���~��W����D�,�V�?���g�g;K����G7��*�nq;a�<n6L��F�m^�b�}�;O��9�c��%��LJ�OJ�����G=��P�z���"Κ���u8q��8ڔ&�nW�a�(������s+�[o�z�H����߽t��q���~J%�lg�#�f�E�E)A;��Ž�݅���S�w!�����P)Ѽ��/�!{ؓ-���-�=��2g;z/�;ko��Ƀ����ؼ틔�x\G�� ��Oy�5}���~^ſ�,yN��Kl�}�c���mL?m��DZ�3��k׮�tĴ�P]i�����LXL>�BB�/vM*�hĸ�p�!m>u����&G"�u�1w��'�`��ˑe �1$kJ&��1�pm�+f/���װ��Q�>hC3瑘��ә!�/�m�vy���$EM�b��C�kF���A�#WY��5��sg�xh�>��{>��h�wH2�rm���;��v@�E��Q��2nkhmijmjo7�������-�������������>7�v��"����:b�x,�V��]���h�'bP�A���^�%~ۂ��O=����H������3��:a�g��^�O����C��-pnu��Z#����=ܶp$ |Y�ٙ�E�)박�+�}|76���=�{�@���?t��s���.&��L�Ʀp�WY�j¼��u��wh;z_+Jнv����鼲N��<fz)>��?-9�l9\IY +%�c�5���r� ��]��r��[�r��Ӥ���A^OzLo��i˝�r�'g��+�[?�jao�g����5���ـ��.X�hvn�#��_[�w~�\F���G�ӛ�7��"�	,˝2�K��v�y:����.����&sN՛�Y��!2`��[�+��U�d0c���:�A��E�>��cdƯq��t���N]���B�=�ڵsw60@7=��z٫%�{^�n�`��B`꼛��bօ�U8U�n����'Z�(���SN�f��J��x_���T�pSj�{7�ĨY~~nv�J�*�>�?,����恀k�3Z@����tݙO&W;fDc#��ǂ5���{���6�WE���)GNή(�� �9v���vy��n���m��Y��q��l�a���mΘ�����{sw�;�`�ْ���䊘����1��x����ȓB����u� �hsa�v�ãe���k���M�+e���NT7FϤu�Ю�%'0��4��W;�~�������R@ZU��~��f�����f��=�%�PVn�-�=�#ua�ϧ�6_�l������5z#똭�{b�՘^��8@vp`��I��MUU4����6�Õ�q���:Y0��Gvp���"��|M�q��6���Cvxf�(�2��΢�f���DmvcI�]�ݛˈ���Y#��x�y�SF 3��]1WY�Z(��JӐn�8�v]���6�q�k�Y��ShWAu���bZm>�����d,RW̠�j������>�x����{N��c= �;��#.���G��-���۸��*vf�Rx��J�ӧء�y�eдz���V�>�O�l�龙Weκ����B�˾գ%� x�vp��{�<��f�l����Eo巚�lv�ͻDAa���Y�4���[��3W���:��v��;���%�*�ֆ��"��5��;�Ыz	�I�8�%Xf�HMS�۫}�QD�)W.�*-�AN�oι�^ơ�^��g�x�z91�f�Jw����js�X�~�S"j]�V���Ҵ��|:�@3��{�l��:�d�K	l��u�2�km��ݷ��KKc��k�m��s�8�7C'gg(ǀ�zc����iv��&����ģ���9��*�����j�h�f���#�L�M	JS���OMyytWT�0���;Z�����<���In��xkN�h�o%�IL��q�V��6`��PD�ZS��.���16��DV؍��Ol��Kӧ�)46���,��PkO�u��1�X���qh���4�1MSo/<|����t�m���=��`Š����͢�4�7s����8����|���klhm�h��;ik�뭶�K��h�1殗v6�7g�讷gon��$����y=~a>]���i�lkE:<�Q�覩-c@m�h�xc�WZK��u�����7�F�6�:�uV�ZF�����9������|���W�u&V>:����;��'�gC]��ؓiv�Ѻ���5{��\�T�?��TK2�O���J��PLMQcf.>/��s��#*�ivO
��];{2�ȗ�5\��8����� VӰ�3����I_ʃY���*�AF�1�S쫠o�<�c��0�d5i��ZE;got�#UFz$���v�n{�<k�1�ɗ�����J���葫1�ۊ��we��t�sV����
�<u�x���>QÍ^�b}�M���Ƕ{IM�d��&�l���>�!7|ʣ��s�G[���v��*��
{R�żI�(���j�}B�cjA����{JM�"��d�9L��{�k}$xzl�C�Z�WK��qDp�,]�*)='�iP%���PG� �1�'�y����I��s��qX�:�?�L.LRs��Z	�˽�I��r�����ړ��wl]�\�B����|Rعv���;�ʹ`��"�Ø�~�S�P��z�T�k���3o�EV}�|VLIr��+�b�kM���Z�=�cE6V�;�k��+τC�����H��^�ƕ4�fȸE�U�~�8��KUĝ�Bׇ%F��TF�����g�Ӧ;QMB6������d��?���'�{@�==D�ȓݶ�?�vާv-̰и#}P�j�M6�j�d����óz�__��E�� 	���,��b�3_�W��w���{w����n�B���}X����t�:NVjU����S�>�O@S�rWT�k_P�A���6��m[���g�/���,O�cZy���F�.��jFE��a��ꕦ�瀯*D,$NUO�)����/����ݐ~�����*����;��6�9�8��;�3�4�Qq�sb\��J6��4����H�� �~g���.<�� /t��l�7fK@m��c�璱�Bo�Jvg}pI�ğ�>}�L�V���E��3�yw�Ou��*t�9w��&׻�F���R;ٍ�s��Ǒ�f�3m�f�C�q�H���������?�>q��+�Bd��B*�)�]�'��^���cMu�k�mؼ���/5��u���8��� ���褖����P��G��"�"����M������:s��~1L�G[ׯ��P�j*B��%�+o��"�g�]?v�䞬~��Y�T�eͬ�w9[Ԩ���D�P1���1���	���L��R~��(^�J��f{�]���ۘ�xz���aH���t�փG�=��̇[�6�K��Y� ^L�I��	?ZS�M�-�z�E:]5�:�j�a�5"z:7%�r^��;�i{�4��Կsu�̯�Cv��P[��ހK&�]�9�uxQ)C�XN�2r=��=����Υ^�k�af�t�K,�g�����"S�+h��I8�؇j��ֳ�#���{���G2�V�S0v�q�� �\w���J�����^G�������E��0=�1�I�.j3!7� Ä@?�"��uUu�� �ߴ�6���m�V�P�޷�=V۳�����~�_�/���w�'i��8=��ku�[�_UY�
�InO�jSu��n��k���`�����|<&509���q�\O,����]�f]"dJ�&\Jy�x$d�X�y��vt����H�a�;���Ur�%|2�[��Djuu7�ʅ_r�.̀5=%�2Ғ�kSF�vm�[��?��_����|8x�A'�V$}�QC�O7�QU�f�F=
X�Br�����{1���.�ʏe:��kă�u'G
^��Cl�D��2��!=����Y>���tfިkE�]�;lG�~�	ߔ}��S�j����="۫T�8WP�e�FMy4�սئ1=�W�nB�v�L񐺠�99V��G�2������.9�*P!�ۚ܅y���t%��4w��>�<�%��%���ފ<�H�@�X�'7��T��O����4R�=���W��b%�.���l���kk�L��t9G:N������}�������g��@�m��
Eu���[�u!#�zS5�u���%���X*麃ם�1xw�ۺ����T]�ϬS%�O���CY��3z�S�+��I�<�Q�ڂ�v)e�[F:sc��� i���m�w�iF�&,H����r%}�>^v�럴���2Vk�r8�	ybk˶��%4�R9�����q9,�f>�������SG�\_����*4M���t �7�o�T6�l�Ϫ��J%�C�"��]0WKfu+;sN������-[�R3�E�Z�����;‛���GD��zPf�吭�fj���q��]�[9TȽ�i��s�'Xo���ZY/�3��C����փ��/��a���Tû[ok�	Ҟ/`:�N�XJ�7rSM�-ukq{k��05�b-���X͔�uZqf<R~�,�%4z��y��H�b��T ��ZҟO7_�@v��6�k��<�ƃ�x�o��B���w��DS�TQ�ѥ�s�P� �\��G2���S�O���Nw�¤��vl�T����Ǉ�
�L r���bԉik�Z� (Q^J9���"2-v�fUl�ro���A��Ghs��&4t?>���e���Κj�R�y�ժ�O��+�I=Ч}�,���lY��� �ą6�W�Y�|��)�ŝ�<�A��mw�٧���F�s�,�̶�]��7��ڈb�٘�H6��̲�%Yz��j���
l�H&A�:�m�/	*�P�Ģ���΍]�T�>�s�u�����qc=����8�t9�#G�g\� �N�RPwuF�LgcM���(a���s���d�?,��y�������hC�O����e�+�6b[6\����$��Q�&��-�r��jkb�o�D}�r���nr�pֻ�%,;�Fs�q���F$��rn��|��v_�r{2�U�{��#����Z�sȴM�72��d��98-��D�T�p^��Q�RW�`ۻ�fGe?�)>I��Yi����Tw��Mfd�n�,�PC�fͻ͌��(�躼�̟^�T�r��/�P��Ñ9П�	�0��-[�f8�����9������9$�j*;s�Z�h��N�ͪ�����[���=;�j�����/A��q�L2a{��W&�M	�R~�����Z�t2�ů��iW2�|VP�Qp��9�8�����K�F�ؾ��l���K�šF�֊�v�����,��R^��FȦ�*o��a��C���-�v�z~�|� ��~�,{���%Y�U���%WK��R��tǈ�^ժ��9d�-h<�C2�%%�=g��ͼ��8�Z}>�_m�l��n�\�莐e0R����T���7����*6�R8q���:�w�8GD>�u����G�;f�c���a���pD�N!Ul�<ܑ�Ȏ�}���!�qv�O���e]�87�!.�j㓳^���롫Sp�lܝ�- n�*�܎vE~��|ek^o�B��S�@g��˹Q��sᐮD7þ�}A�1���R�ܺI�f��vQ����j�+}ez�gU�%b�ʪ�^��i�3��r{�(K8�ea`_d_�r�ǽC"3����_8\�;j�pl[}1V�^�G72K���k�����sr���$�'�ȧ��������Z!��Z�C���C �d�,4�srz6}t	�i9l��4#k!��s�Z���+4XK�55v}}>�ze.5lPǮy�Κ��S��]C�@{�DZ��{K���@������Ht]:J��x�wjFD���<Of�v��=�t�[Ӭ7�)���N�����ۿ#���C���	������R��\3[t�s�����.�{`Y�F,z��7��W�~�W�������9��>�Bh=���~Ww](e��Q.�wk�qug�W_��͎H{f�U�i�)�u]mQ"u���S��[\K�Gf�<s�:�Q��ZUT=PX��+�(1Nf��;���S�E��[��3�\��N��>�9-��Ɉ顋����O8vF���Z����^�v���ܩƯ�b��R��dd�o:~�!5����n�>ǹ�˝6����LT��;�1������
F��~�1��T��L������;�,북����A��d(A�������o����$�ϔ��B�#qS^�����J�Vj�a-j�!�uC��r���r�45댈�G����b���:EWA/#&H�M�cėԚ����nP�M�s�&h�UGb}��fxf�=�^�\�E��(8��2J*0��}��wL��<o��2���b�V6�2�K�V.���H�{R)ZB*yc��/t���k�'3�؎��7 e<�Sx��n��QLy�
i�H�r�ؓ9��.�	�1���P�~嶾?1�sW��X�)H�ay2�\Ӱ�9�:��S�o.TXڅ�&sC><���Cs�#�ɷ�^�Wuu�ӷo[_b�.�yO"�L�a�.	�<Õ#E�׎a"��r)�����KP�g���}����c�|��	�D���z"ub���
�;�qG6a?y(%�b��kT>�i��F8-a�I�}�Nu3
J�>+��_>�3^]�W7���M����@��ȣ���O:��.잫=5�X��>:D�>�,ށ@u�AD���>0�v��|�[;&R#m,�J���W.U�Fus�n��L<�r�v�J�2���G8?'t<SԞh��~�D�X._s�Y�c!�׽�����>��A�1���i砾��M?�:ke��_��{l~@S��������PMk��V^������+܏�I{�pC�f��nG^s����C_������X��o�G|�����=y�@D~XD������؇k��w�ڹ�1��aP3�i>n3muE"�Y;�MV�ȉ�8\��cK�\�b��Cٻ*��.���v�n�N��bmq0����Bz��fv��uNK�S�ڔn���n�d�!͘/j��-�ݻhk�<��T9	�)�=�WP²^p<i�xЎ�}M�t����<KXnijq����b����h�^�	��R5�*�6��Ԛ�PǳWWlG%s�5����F�Q��p���z.�[L���FF�O�{j"vjo;ʟc���i=q�-�y�W�qe�Gu]
�\;��K�yѨT�Fv��0��Ǟ�U�'JN'�vh*T���kX,S%��U��E�.�n���#�,��dd[$^��6����]1mc"z����3w�TNʀ���ޚ�{�<�L
�M��*��8�@��|5�,�U���_)��'U}Y���΋~vE�M�.4
��^�(��*x��������%I�ֱ)H��;�4��I[|��3��^��Q�����Z�s� �)�J_J
���|�z]��;�:�M܃�m���\"�&��7T|쬍��ܛ���\խ�R�v�-�WQC,T���!��U�\��ސ��A�L\��@�]���WT�/|
�%��J�׏H��R.Msz���DH�����2�����75�����}���r�I|��@�ڇ�O���"O�t�mصB��t�78N��;L����Ͻx�|�v�����j#��"�oH��c��?b����΀Q�⽝�E�`���f+��69����RN���Aø��ށ@i��@E�<���&�PȪ�ٛ����V��0jF�B����ܫ;���Y�v^Z7j
Ze��r����.#��ܡ�WKRy+�ן{e0����C2;K����˾�%����I~Z��D����;��M���7uyUx��u�{�æv	Ϟ� �B�y�M�nHLow�Q�nN0���b )V;�3&`�<�ܳof����ys�&;�zGS�o..��������FEoi�k*g�6\vVs\uڗ�ڮ��(���}fg��t�|���И���o�К����'uJk�m��8�ew�����O3k��׃VS���."'ڥ*�!���@��jg ����������%�%�����z��f�rW�
j�|��=��v����N��|����m�T*���r��0Z��4<TZ[@��R���t���}Ŵ������+���.�=O���$�8T�F�o����#����债���l��r����Ak[{�,}	��E�����'#N�W���Jױ�d��Q,�o�-�n�H�QP�����������7�|�T�J�o��w��	�����hGD�{�.{�Si��-���<e)�v�y���d��.��ʻy׏C�έ�S�RH�7���|e����a[
w��0<ʮ��09\�KȬ�R�a�Ǹ-V��4V���ͮ�m�r�ٮ� �#0�x�'G��S�."��L�JKW���b�zo&݉<��1�6ۻV���d�{���=�'��/��� ��g���Ӆ�����H���
z�q�9wD۝���Q�F.:5��;b�:�eaO��`��ʢ�����-��i�6f�r�C���ldJ�T�2��2=�=����e�ܰǴ�t�d�軭?��U�������~oI��H�4e:�:h�EW����;=�<О�6}}ϧ���	����d�zC�>=.�g=�=�s�Y�C3�>�k�	(�zO#'U�I�����s�F�5U�@��w����9��T�Wl�H�p�]�a{�@��~��=��s�ܑ�&2��%��d476�55���[�6�������6���������4444771*[\.\BwU��a�m�]�7��'��=yz�����Nf`]�^�b�o��ӫ6��<X�g���y^���v_�*b/P����v}��ҍ�t�,�F{��p���E�t
����Y�`�Ҧ�/wi��T��s-SF>���^�ʴ��y>w5��d�Z�ӷK2]o;m��I��N������b���SB�N��5�oj�a�|����j����B��]�QL��M����S�U��Y�b0μ�͋�6��w��f5)��"Y�pN����X����7 ne,�ǒ(�d����#(�x�d�FB�`{N����y�(�x�=k�R(��xq����[���髗���f�~�8\}i錐0�E�V�W��`�1��bxԙ09�>�ۨ���w_a�c���Y��A���;'L���:�N�o�zťԻ��ZV��Α��I�<�a��.��5c��i^������v�9����)zڑ]�8�������v����u���M�n�d�ق�(͸�^*�Xɕ"�tJ�dm<�]���@[5Acܺ妞��ML�Z����Y8d�-������Y�*��B���`���R�����#���ĩ�uu���X��g�Ҡ�>�a�a�\�X%г����1��nN��Ka6tNQ�Q����Ύ�ku}$��:�r��F^��<P���!XK�Ɏuc|DQ�T��9�-g$�L�[k� �����^�4/+���]-��7�J��4P�����+;*D�S���Ձ8ƢدF8̄����X�ڠ'+��gG���h�~�8�b`�|3bfi,�z��@��{����Cxx[!t8:�[콦[d,p]��*��o��{��(+�K�]`�sor�l�@���R���U9�-=+:s�VI���ޛ�v�Ap�u����bD�sP������څ�$�c�� ]��+�u�
�E��������r6-u[w����ʖJ�}���������*l�x�j�|2"'Zr�5�ɝIp:�YE��.��伞��f�/�������dɽ�@�ft�	ι�C��~�쌋�Tk�Q���l�R�6�쭮���Jނii�T�R�<맔P�|;��2��5�F`�(�A�\���y;��jYwvS��k�}7;��G��l�q�#E<��9-�����	��cx�n}ud+O��,̵.�;K{�[�w/M��⧂�D��՜�۞�_����,�����}��d��c&	����@J��[ث	J�;FD�gso�=R��n���XE<ɷݏ����<��zzRGDS���"���M��$]u����c�"ˎ T��.�k���]�zʨ��N�㙏�W[�� 4������^s�\���s���mD+/��}o�Ğ���(�8�?�,��H��#&�+�	���$4�.[aFE�5iT�
Ќ���T@�a4Q�6����ݵm��e��C�Ƌ��4R�KO��ד���:�l�Dy�*�����5F����5����k��7�B�͔����q��������h4Ūmi����A]��5�.�t��ա6ˎ�wuV;6�8���:4Q�yt�m��x�PZ�F�mc��WgX�[���ES��G͒��X�GcQ1W�]U��A���(b*��U��h��cy:<��㠪6ߋMѢ��>GX�2k�<�v�����ǛmPbu@Zƺ��'Y�Ͷh�-�pm�c�:�;kl�tU��*��7cy���j<��)���Al��E�-�����>�>I���W�lG��k��DM�Jw`A`X��L���L��
�=�ʁ�k:��gn\ܾ}q��.c�Z��.���3�j�v�rUV)^
��SU�U�` ���!��p�^CU�WX���L��~�֯�"{�0u0�aoZ����&�ȿCV�F;-z�N��)(���~�T+���}c��zZ�}� ���T��ǝ%�I�,,�O��Q�*`Y�aW��:^��5*��u��'�M�<���mKo�c�Ro��{S����)W�5�F�y\@���F}Zʶ4r�՜��S/���˻&Y����d:�!��"%�Tc���7$t��07��Ǝgv0v�FF��[s���됥�"�b��}j��S�7_د������Ǭ�	���!�w�m�T��}ݵ7X���Rԃ:n��o�-T���Q�0;F<&���Mɂ�����r��u����F�={u��\!��D�G�)-�i��Y��9f��XŮ2z�:�ʭ��T�lOuwۛH7/]Z�^�_^Pn77'Ѣ-�ȟ�7�E�*q��dߘ&��%���SK+-�F�>�;������OK�QL��%>��Xۓ9���{��Y�|~�Qp?r��${w��Wkc��}���P�2F�6Xt�9��T�{]�-�>H�!L��wB�K��ɩ�,�������?%_���s7�j��YY�CI9�L�8n�Ʉ;��]��r��M��<���w�Ȝ�9����2��w���m�z}�o�C�^qŕ)�2�o�����[">�6��m��=��ު8Vi�;ݹh��=m�f�zߌ��{���M��Ld�9�_���mW0�2Y&5<Â{mi��g�л�OH�GcG<��l�@� ��vY�
h�BY���UR�]�'w�б���j;�e�%�[K����anj�������N�,��$�����Ps���UJ:.6�h朢s.��������dL�k�^\H;؟��zC�t�����\�&�Q�n��m����ͽ2v�LV+�j�k�g�5��H���r|�T�����G���2��s�1��M�Yȩ}�<��Nvs���/�����;�9-��i[�Q8��<ꂔ0��Z�wkv>����A.BN�~5�?�r�������AŞ_Ghne;PݎN��zd�X7#�6��ܦ��L>������D祭���Ƴk#�՟|i����{�8�)�!:ʅ7_���P�i�}�m�=6U�xf��9�۠ox����GzY<�
����0��r�P���eo����PJ�E>����Q-���&��qt��^�D?ޮ�t��FocM�����视����͌����ߗ���z���h�c-P���O��f�iՃg,������Z,ů��-�Е"8.�t�dYeW�o�ʮw���Fm�/��>�zQ��U�rR�ZVD�szv�ݫI�b�M��Ѫӊ�U���)�M�F=�X}���-o��*����,^���ϭ���J�BRh��Tם1��ǼyaЉ5��^m��Q��lC�O0.占�S��6�	]cxQQ�1~k��⃸q��6�Z�<�*^W���yk��Q|��G�vD�ޓ�~~�ML2�Jn�[q:i�*<�y	�Y5K��fv�E�Q����=Ր�^�[S�..�d)Ћ�W�Ȥ��?6�[eW�x����fn���2(E�#���S����֯I�ו�-Jy�;���P%W'�QͫW'�U��r�WU�n�m	�ҞΞ'Q�q8��v!�ПH(��͇s��R%�s]3N�!�)����j��V��^T��N���?�>�J9C\��`,������Λ%嵴f뢮ぃ��U��Pm�%��K\W Ү����	l�3�ѸE3\�:z64��?���yf�z��ec��v[��S����5����Ot5[�vbZ7j
ZgB8�&���^C��Q�ׯ9{ќ�����$'�R"��o�nˠY�M����vű���mH(��vM�=������K���7��J��s�� |��B��á��o��U���'����߭�_���2`���;��.�9f!�NK#��ju��{�vM�-űQx���.�����`o�^���E�M��A�ETv�zm]��Ձt����������Sǿ�� L�0���s�@D=��N{Gmz���7�x@�hmӭ�u3qZ݌�rz����i9�k��3G?�3��r���4��	�q�eڧe���]�.v�Ƭ��çh0�p�6)R�>ldV<����W9+�>�eN(�=?�LK�@�n��@+d"]	M��VCO���?V���ڟtq8�w��+(lܢ!��N��+/B�<�H���Mz��"�+V�c&'�]Q}�9�i�U@]�{u�d�)D�l��*�m,�Tw��yk��(�u����X`�/m�r���wR��@�_l��蕏}Йs�yO��P��
/��Ɔ��ħOb&�ݳ�Rӝ=R��m1q�\_=2�p�5-���1S�c���Z/��17�T/F3�յs0g냚�g���ѓ2����Y9/B;g�9��g�fO���޽���W5��(r����p�hY�����I��c�/T9���~�`��s�,B���ʀ����?��dC����L�6���7z��r���1��2�$a����Wma���CjNncRР㼚Y�4]��N3�D-���xH��Ih�`=�V%��}�����BX�yK�t]��A��>'*�����U�ªGף�/vZF��׼}z�G���:�{&��⼭RM��m����5�M#�xj�p�􇗍^Ʊ	Wm�E�6ħG'=��R�R����L�;������K�p �������zr1�@�O�<���}=/�PY2]�P��eA��6�t��d)�W\Mi���Zݕg%���9h�EW�r��lvF�����>����������f����z����ć^)\��򍷤�g�F�IN7 Jk�>ϕUc�{�#^�^�^E]�r[�ak>��.�6�{�W� 8^��.��3�4�A;q�cq��	-��a.��~�ކ�Xoޒ���g"w�ZC�����(2�f��C���7&�e�Y�:c)q�Oz��@�c�Q�W=���(Y�fDO�N0�Dŷ'pM<Q��j>��U}���c�͵ޔt�0o=7#ʷ��1~�|�����s��b5�����k�e��E�o���^��qm^���36j�a2��|�hw�C�7�(;�m	Ѭ^N/�Pq$<f���/b@�I���~�),����]��][����|�У�q��!M���O��h�:�U�'8](��H߁Tj
� �a������u�Y�_sǍn���T��--,���x¹��n����5���.��^[&υb��|m��	�_O>�֟��w�z�������wT΋�̋-uw��1��& �7��Ob��7jf�ɯ��.>Ois�iYSq�����ͷ�s>Y|�Tۨ)�NXu�����\���G�U��J&]W�o�*n%O���4��x[%*�Ь���рo���g�g֩=��(����o�:��w�~?OO*��^P�q�Q [㸦kq����}8Fc�މ�3��wNw:;�w�l��Ҽ����Joo
G6����L3�za���:��Vb����~�������=x�RM.6�V����qP���A[T���iv�+����.��	#Y��#~�=3�j��Œ�=�޻�SwL)ݝL���-�̴G�5O��7�ݴfo��K�W��~QWlT���wg����� �����d�X�ua�.ֹl|�K�vj+v��r(2�v�.�Oqއ�SZ_-�o�t�1�X��0o�B�n�%xf����n�,]��gV*G.C����
�<9Ps>�ژm27��:��3�h9�ɁW��{pC��6�� ���nܡcz�H.'���Z|44�otOGs?���V�,� SY���I����&}�4�j����缅���1i���]K��=4c�*f%�\h�N�~}n_`��8���*��L�|;�{[�<X���h�PY�S�1/S�B�ւ�6�	��A�9�nJ�Z+]���s8{��������,�ؿ�s�#�7�#{��r�ܩ���Y����on�_��Pg�v�)���u|���y�LQHl���W��ܪ�d���8�m��o02�,�pSwZD�p�����L4����3W���@�>�>~s3qD�ۿ���3��_�J���������f���ߗ�Y������#��Y�c������]�i�)VF�ݠf��8���W�)�,w�P[��<�Z񌢳���>"�nE���8�x�y�5wAY�J�''C��׋k��(�5����Mm�����u�65�+�C#� V8i=����l�a�Ld�7��Y�9c�SUK��e��l�9ڐ9t���ܑ���9���]����p�-vN����7n��p�*�����pا0���>�R�J�ԥ�n��zcM���[{�}�@�W��ř�n,7�}�[Ѯ_O��O����%���h��5�0�;7����>�:=�]?C���R�hVk��MqP��BL����+�}��|��������9��#�%m�;�:�ńq_g7G���ḝ�jm�c6*M_gTj���`&.�'�d-�%��Y S&v�T�M���p��fb�a?4"V�ʸy�w6��e�狾�s[���%<�N2TY����NC%]��bg�����T�Q$�"[�[��!��>�/k�������3�vbN�sb����	��o_$��ݩb�F�Wu�2��}��B�>�7�)��h�>����bY�o����t��6X��̙���?B���ޯ�(RO 9��J�c�#��w���N�T$��ؕd'�sF��jk�O�5�z x�e�z��\���7u���l��~�v�=�.��cGϏ�
�h�*u>ኑb�m��{�y��]9��V�q���f��^�2�_�HbOV1[BnV����Z튒�VȖ�z����~��|�oVj��e�H�nE>�U�d��@����w���^�P����N�r�%�u���D��9���W]�m2v�qV�*�&ض�l��xC��dM*���Z��1���N��0������`��f���ʅ�1S�p�s>s7\�[I�t?M�~����j����1Ej�����������(�?�Fy���:z#�k�|3@�%$��rv�<�7Ǹ��;�Yd�����J��(M�%#�X1��6��O���&�����^�c�!���{y���ޫ��4
�¯�v�#�v�=�c��H�678�noV�4�6������C��5�T�/28;C�ܺ�HְՓZۓ��\\����Wwbׅ�uا��{d���n�{�Tv���n�V�t�.;�޶�Q�_�v̀Q��f��7,��C�<�b?��+����f�޶���,�Sz��wW7-�Ƭ��~4���Oo��>hD�p����".���ٞ{D�̟ʳ/;�} �[eeE�p���=][m�t����D-&�T>�#�ږʊ��j~���C�i������蛧�n�7�A���M����]\�������Jss���# ���9~��UH"��Q����ht������<�2N�}~��P�sE�r3�f�����y����#����y[�:9��޿ Z5.�ص˫ ��&��[��H����<D':�ܬ�3���S�emVc���c/r��G�#W�b8)ɻ��F����|X�{�ǳ��z�H���휋8u��e��
�̩�͉+����ںwrU��3�}qn�y��]������d��w)��.f�Çʪ��%��"1���OA��.�M��N�V�|�"/n�F�s8��u��^�ٛ8���FN�9�ٰr�i��RT_P�Owf:t�]�k&�.r�flGLLN�Զ�q	�&xI�έv�h�nc3�F��NjӛT�r�x����1]!�i���]V�KY�w��Lv7q�3O(ݒs�G?���� w ]�2�Vڤ=�����|1�����ɫ��ʶV-N�nL�_c�o�JIf�G����wle���96:Ym=p�����i��ӽq�f�$m4�<9��ҷI[�R9� ��K�=e<��jع��'���[8��Q Yz%�7�yX&���d�g�+v�r8�B玡��wm��<�X��k�?{(��Y)�zz�W%\S;��tĪ͚��G��]������m��`:�K��=�-Gr1&���������<���ky�kkkkkkkk[kk&����ֆ����߽�%�c�>��]�Ԓ��e��̶�I'���ǵ�3V�R�*��/>6������
�<�[��A�I�M�!�_=�4��@��+�#W�{�o�7m�ˊ���0�<j�Q��V�����sBƦ��.\�ܲ{����gp���R����f����6b��@A�V�YF�V�؄��-�^���F�zTd�#=��WD��g��ứ�H�����ͷD��`MQ��~[	G�O�a��9��7��<�k��qi���Y�{�w9I����D��'L:�&�"Z��|�}�&�'��];	r� ��%�j%=g�Hz��P�d/7�V:ZZ�f�C��Pn�ī��{�,J�O{m��*��+��M���7S�bpރz���mގ��,���y@nc�z����<u��aS�޷٫[B['_�<Я�nEۘ�t�zkf�Jm��3����eu�n�e��}���"��n���˂�1غ�7�8Q�*}˶\^��xx�_��SJW��5���Y�wd�x��z�Y����5�s�c$Y���G����T�}��;.�D	�xI|�B���wg���)����#u?d�Iݨ��e��Nr�b�'.Z�a6�.��ܡW���K�=݆6����^������|�9;-"�3�ݵk+86ڕ�@�zN�60�~����<m�<9���^A�@�K|��:�Z��8���L�u���eZ"��V�^�^����ᦉAQʩ��U��=K�;[t��_Z'
�X?z&�ϹALi���c���p�ܔ�R0�xsnĎ]��칣.�P��ɀ8z��o��ܵ\�5r��k�K�9�Լ�x��&'W>��Ź����O*j�s�+\1�"��;p��C��1mtdXy��Br��7�T��%⽏H���2J��?��{����~o��]��0 {��m�Ү��N���I�.�J�=p����Z{+�fB�R�t������[}L��w	wz�m����ܭ���6�G��'C��{�9@��J��v����Y6ȵ6���\��ʰ���(�ﮡ��|���s��;�O�����x�{�w}�	�����pu��s�0Y02��d��U���/b�Ϋ� x�Fa�#����kq�BV+�V�G;�=�
s�����l�l��	�,kr�^�Iޤy�\�W��G�ˣ�8w�M(����>���fM��d�*=�Y����Ŵ�&3	Z鳹��GSs�bC->˵X�&�7)�nLi���,��AZ�;kI!��|K�]���dڗ
l��P�ɲ�j���z��9�%���g�]&凛��I�����d����a�u��N˛�p�L�_>�s�I�B�EG1vv�۰��J�y?'��8l^%æk����}���a��U���GU|^�]r����M�1{��?e�b��6���=�h��B�=ԜwzR3��{���7�)���wT�;��0��%�H"Ȓ���:鋭u��h)�mcS%1����ض�񢫶5��+m;kc˪.�ŬDth��Z��*��mS[��v4kN�PQ1:�Tv�SL��Em�*6փ�m�54�D4���G�|��{q�m�I%A�F�ܔ�c3U}ڏ<�:�]b`�֘4굊"�U����1Q��Atw�j���w8�h��cV#�Uu�i���Z����P\b��٪&
�c�h'�kF�]�ઢ+c[�&
/�n�أ�ꉪ*��"6�A[b��v�E�Ul9�4ED�t��ALME�i�q���Q�S�1QEъ(��DCF,�[�PQSM���h����[��i"��(��4GF�lITZ-mh3ES����,D��(��5M:�DZ�UM^۶��\�;���(�7t=רR��u'�m���齓��+>����f�׺��&��7K�y�]���>$\+GF��s���|���V~}��H.��<3a����z#W��u7&��u���.8f�vH��rhÍؽ�R�l�c6Yq�z8۱�L��Cl�R\�^�Asя�U��$�A��i��#Kia����яU��J�5sD@³0�ں�9��_v��Ԭ�	��Ѣ�^ή�ʹ�����S���x4'oD3���f�@���[oH��SA|�w�Tr(����߈�n�{�ժ@���ٺ��@�ݧ�&8��a]�2��|�=��F��l��[�T"Z��A�c�f�?tߕٟj�����"�UA���Ƈ3\fsD��+������ʡ�&�����S�=�H\MA!�m��ܡ���6N�df��Kɼ��H)/���i{���z��=�	�Lvj�u[鹿L�e�}ݖ�׽��O���%+k�''�ժ���`J�1gd�C�;J��&'k:�o0o��|qk2�U����Δ��q3�x��3�ܨ�xc:}ˆI������l��Kc'͛��������!�Е��h�X�@�wel��mK�Ƕ��\��ZZ�eP����у�.{Q�{������_I2����L���>�Y�� ly�����%KM�[ 
W��]���	ƭ��'���+�o�I��˭P/���֑�2�Z3�ԭ`���C�4�6z`=N�0Ѝ�u<8��@��1�+�G�9C�U<���퇨{M+tM�Yc�k��v�VG1�gl�؇�w[�& �q:���lmf�c"v��9v�i=�h¤��2�m-x�7_|�HC�of3洷d>��{��u AA��2����\���"Z�א���Y�e[b���~q��j��lX��,��z���:�	���~}�ل��_#�f��E�8�kRA/E�o�f;�?a��/����7s5��˜��{;2��9��-r,R��h�V/6�;�ycm�6���*Z��g.�����	u�/N������9�Q������ɷ����s7ۑ��ߥ�2��[��=���?�+�8��B j���/.�qEv�oTa�86�+�z��@�[����K��$a���z�U�ژ��*��ރ�`ބl���%l�pi<��>�Շ������u�OP�uj�7J�o2��vF�R|`�/JIR�����ջ�{��7τ���|�.���f������Yq�T��`5��Qu��k("7I��Z:�J�W>cdV�/#��P�ӕ�yO��������� �<�F��ͷ�n�Fg9�M!5��H��@�jV׊��)eP�j46�7;��\�c�w��g�Qn��l4�8���e�Y&�I�/ߵ��K�c4��_x4���^��'�q4w!��t�hc�/:�l5��e����^�xK��&G���sx��[���x�Fڐ��
k�!l����s>��o�*�<�o��f�@r�AF�%�W^SGZ�3�\�w-�
��Wp�7P�w鬋��3����O����
9&�!�u��95y��nb�o6�nη^ػ�ۻ��O�:+�Ϸ3�h\���Ԗ5f�5�V�"����_4�wW=g���PV��2��%����\��J�l��CKs&�3���ź����g��^�d�q��Ҿ)�.��VCM���:�k*R��=v��kA��V�m-W{���n�C�?��ym���{H�B���pe�k�;73���P�o���˶��h8�p������&N#�Θ�y�����誶?��	�^�l��imL����|�;�z��J��9��=�U���s�ڞ��5Q��ކ�|=3�3m���0���q�C�W>�FGj�7vG�1��9f�����bul�4KH~>����e�Q���uۭ|{�LqQ�㇭��� �9Q��n��N��~7��{�3\R�u'O�\�j��5��F���dDd��I`����3�/�8��5��u�[�{�/�7h���nc��w%�Y7#���NW�c1s6��/xe����Ou��z��6�j����ہ�SOj���6�Y�m�!e.��&t;G�r_�7��nx��~�_���uO4f�=����Tt�W~�}�q�S��=af��=3��i��śCʮdQ�R-�����=�q���(��{�׭��oZ�Wkf��8�;~%"mmlҫ�Wq/V�$f!�&�c&~촷���ʖ�s1jf�㛗��2a���z�6L��}.O%�E����Ѳ�=�zq��x.�d.�i����T����A�>b+n��Z|�*������{Gz��K<@��Lb��\�p�O���hf Ρ�:�Z^��[�`��f��;xU�e_��h��ed���*���`��#��&n9�\���w�"�T�s�}�E���z|,�~|�K�U�[);An�Gt��0�7�'�~��3+��vX������2�1�g��MԵ_�"J��閌Z�N�랣Ӵ�^�RP��h���c��_`;�ϻmC��w�����Q���TQ7�=yˢr!�"���{U���Z�I�C��Н��o>�	�p�֫Z�t�E�Y���Ho-��Gt_r�����ů͉r���z�f ���f=�O�L۹ʉ�$Ϣ���h?qi�`n8�P�4�ҾZ�u¶�d��֨`�ql��m{�����2��1�˧]�@�ξ.�Xr�/KT1�K��z�utm�Oި<J���S�m��~�u�[�����o�Chk�N�]"	O��z��@���z!���\L�6��^	�U�#�|V��w�X��KR�n�Zs�C|���~��|��e�9�F���=J���Q;>Z�����+�\ji`q���V��\Z���/�[�b�Y�$�+�嵝
�J��K�w=NE��=��������U�c�vO�!p�6��l�x!��zFc�g��ɚG��,oz��ֵ�Ɏެ=g��#z
�5���-S�l�w�T��4i�G�n�Oozz�tE�;3� �Ģ���w�Wo8��*�X���Sx�!֒׽�ǲ��;��.�������::�	JT�rI�TVd�U*��4��¦�v]Cnj�j�BGs�z��b;A�9+J�u�Z�v�A�綡�nzK�4w��w��UJkG��kTfw4�U���~q+���VS2�[o6o�/��kHq]),��y�s�V��:َ S���ƴڶ�s5b�nژ��t,�_�ЉeO~Sk��U�j�����X���dۨ�,�����գ��'؂�v��\�f��p˭��k�M��7[7�v/;�m�ueIUL��Ϊ�9m��i�|��"�:�6w�����(F�'�(������_Ki�{]DF=��xc�U~�oϾ~���d���M`���4*^�<u��3�N���7��Q��>p�_��P� }���U���
�V�����ǎ�:���꺘�3v��]�5�cg.�)S�LiG�nܡ�;��]H"
A����3z����L��o��1Ϻ�>���]k�n�#SA'����|��퍻�M�9�5�Z���N�����H�&`,3� m�~���������T��(�����^pd0>��+�Yt�&���}�U�c�*�zC��M���V�u�@/�'�Z�[ө�lL�M|�!(�"�o]n�d4黙�͇��X��	$I\/x+­�9Uz��=��@���)@�/���a{22zT;�g�x�x��P�(���^*e�����k*����kkQ��G_T��R�
�I�X�ju+ʽ@�P�|U�QW76��۹��k�]�3φw��m�������3z<�
��ڗX^��:2Ѽ���Ю<V�q��U�[(�`@Ǌ�;>c���nSCW���v��:�FFٸx��lMvf���Y��Q��9fB��s}�ۼ����G3[&vL�����������V��1�����Z�����$��Nc��:N䕗����BהV�˒��3��n��[s|�}���n�fV���6O���+�m����^���4ބ�GkM�}��]�!���jo^���%M[-�[18)�����Y��vθZN�~IR�Q͝��#hĭ��3�:Z�nkd?oz&���;���p�
 �Md����II}Һ����\�<ד����c��Nbh�/����S���3�qEL��G\��Wq8����T���x�T��9��}�8H�Ʊ:+AF���/��U,���|ovм܅t+S�W�B��`��ʅz=�!�ٽ�á��d��G!c��+2(�m���.����w�����#m�������a>~��)8.�JE-�M3.�(n�����3���=>��ghܴn�4ٟ��xa��d�F�O����j��]¾Ȇܰ}�e�<�3�%�V�!��@9ԺZ��������~F�1�s�Z.}�&N�c����M�9g��	P�j�����0��!^͝ɘ�^O�鴈��3]uw���a/#��E�����P���K�t�3d���U\j��ONӂ�KE�m>�r���n����8����\컯�`���.�eqhC�g��?#��χ_�e�^���� ���A�+��&}rۀt��A�q�ת���I��T^����SB�{�}11t���[���Ef<��k�UTa�P�缶n��������_Xނ�ƺ`>����r�O��~!<�nCef���3gl�铆�ӕ���|���oy��F�:�T\pѭZ�d@�y��e½��xz��K���,�*jo�qԋ�]-wWŬ�b��,�����}�פ��G�{3���+�(�[["�\򷺶0*=&N�;]�E��!��;vz�,
~m>@N� b4��Vx��*�s���&\�J��Ndو�yvٸ�kS��dag�u�kЁ��D��Z	���;Kw^��u3S����Ѝ�|<_{Y�R����e^w9"5oW� �Y��ұuWq�K6*���.��B��7ednP�!7�\ ���k�ܶ�{1g��ˬ��`?��6�^�9L���e�akSo���o0[������E5V�^���]nN���$�������
Ϸ}k���e�0h��,�5M��W��'��K�O
�����`�_yK�0w�E��K�5�i��Y.t���{���0��u1��ś��‾b����Ι�s"�2m����{=�FOv �Z������,g�(t�ҙ��Υ�:���$�A.�觊�e77AtX�ͷ/� xC����0o!}H�������v�|�f@����-�k��a�eu�ȳQ��wv�q��v��6,�������֦��ڱ�嶘�������h�l���͔^�B��QS�J�7=s�%�`l� !/���I��u��P�F�M#�ߤt6��j�tVz&��󋻗!��<5Ҵϝyƻ�muB��d�q�Tͦ]^�o���Ǔ��W��&��PwI0��,�#�,�d�d�L�L]ٸt���+zs Z�x-E�t���rϵ���0S��[j��(��#zP�Ae�9���g�lC �����R�3�Q;�b��4��ם,�K�$���C�q�;�-��R7쌀MrcOE`�VI�eÓ��wOp��s�ԸG�����p�mU���%]�K��:S��g.�V]��z�ެ�����M��O��T�.۾�@nfM���������hmmmmmmmmmlmb������������;��_��"�-�)�l<�GB�o񄊻ɷg)�5ĝ����Y��hv_s��7)��F���亮�bw(+�9G���j��f�8��q��U�T=�B�*g6f��S��ė�;8S�`�l~�ߎo������/�a�m���5�>JJ�x6�U�9��}N��P��N�7b��ǘy�!*ԽWk�֑3��i�2�����A'-�p\��b"�';4�~�vm���ҫ=�:'��T��D9�HS�U�8j��众-�j�������D��S��)45s*�VBW{/r�wp�hd0���ZF�#D�A$[Lb��G�V1[��{܏+�G�0�t���V[Z#���V��[�i�Y2���.���i��׵%��L,g<a:�tS�g8��v�<f��`7��]B�%7o.��D�w�w1x:�n.Q�w9v�jv-�E.R��e�v�Ѕ��5��&t�D�VB��E�F�/_U��s�Xy]�&�0��\��o쬔D"�/���;�P}[)X@���R��[���4q�i�8�@1"���7/)���8�x̓����k��䋟vt݈ts�n���}v��ޛ@k�-��yM1��-Vx��۳�V<o��$@�wǞ��gNce�8�t�=���9�۔��$�%���F�+��c����HUȷ��,�>���׮K��ͣ}�e�Y��Ȋ<��-^��kv����d�󖚒�h�&	��`9������� �,	EeK�L��|�Y�3�M�}�W��L������9s�����m���	u	� q��:![i��Xp�պ&[[y�AT��iEf����qٷD���L�r�,ܴ#w^f<V��y�P�rV,�P���].��h�����l.�o(l"��F��շ���nN ��acbƳph����)�����⼽��M���)�%
�C��m]<.v��������}Yx�ώ���#�&h�ЩEćǥm9�-d�o1�[�=]}Kw(A����Pk}"+V�+��N�Xer*qE�|����q��;�Z��L$ɰ��^�ۜւ�o!��j����͘O����QA�����=}(ǋ�3��W�T/�ȿ���7���J�_5	C%Y�ô��M5u��Hp�:����#��%��3Ǯܹrq:x����]\L��T�}3�SLй*������ks���`�w�ʯ[���m���e� ��DӷT9�'������/qz��m��=7g�l�Ņp���$��ǰ�F����e��S	�͕I�A�k��58�k���j)YN�_z�!�V�.�����Z�����+��@ �P	e���2�0YH��$Eck׽���o���k���S{<k]:_q�ԥ��:�唀��0>���O'��r}\"�/��=hg����2�
��+NR��g9��mMp�ܒ�f��������LGcHF�	���ʒ �*፣
ǕTa�N�[t	�A$�E���*T1�"j9	�y�kwWSݷ����3�clX���E�0͵j$��uSSD�ST���mT:�Ql[SLES%V��e�E"�lD_W_~i.��v�C��kC���"�jk�E3QQE�3�m`�����ƫT�TEIi���0Q�b�<3���1Z3k�� ���������#�٫cAQT6�Q�h�tF�cf-f-�4��Q��ƍ�5U4Mt�S#5�u�]V6hֱ`�5�`��$_��f	��UbM�q�h$�c$Uv�Ѩ��D�7cvu3PKA%QIMAQ;j��gU5m�l�i0U1�DT���ITy�CVƢ��ֶ�$y�Eu�"�"��4I;&����F�TIM��
�ƀ�c��ETV�LLT4_YqUE"`�#cM;&�cVڂklMT��*�4�5������I��1ؚ-��뵢��Ӣ`킂�:[���i(�UX�������E�Y��E$=�w�l�ǩDn�^�Y$3�t��%
�F�;R�m���MwJ�Ӳ��Z"��o
�n*�	�
��ͱ*��V8l�-����6}����F	ܶ��f�o���w>G��z��I��g�>�\�m�Oh0`�D�YѽBg#r��5����=k��Yƃ�g}���͹�ȇ�:Ԝ<A&��=kv��l��^�1�؁����*	w,��C�0���:C�9�F{��� ���ǜ��U�����ܝ*��x�}֔�Vo6�!.�������y�j؋r\x7k��Y{�����9`A./ݖv�$I�"�lfC2 �~:��3t��e{]��ws�9��a��cݑ�zr�*z[-�[*DmY��Gw���-]6v(�n��D�	|�qY�t̮��Ȫ��zjz��.�@�2R^1�~����_�q J�^�g��lR2��	(k�WN����;;�*�H+sw[Ib\:F�XU3X�N�p��m\�i�U�;}WZ�Zk��}"&�]�kx��P�O���H�n���z2�;��/��m���0d���V����M�%ێH|�ӦvP�3x�Y�s��'����%\��D�/搟�7ͳ���=�}��l�X�+��d>*�oR�Ʊ�`Z{�ʞ��M�˕��.�S�&�Vy�����(�!0�����!��Ӥ�SV�>�L��5�y+���\��X0vp�i���;�Ć��32������n���	�Pl����L��*�� �
�rDF@駖��h�W�Y�C�U�V�bs&���fS�:f�:A���?�]�7���	�S�gUOf���^$飕�F��i�=��v��6�/Ơ?b�Ye@�ⱋ�-�]����9]�a�J���m-�+�:�gS�YQ%X5#chp���^�,�?o�1b���o4{o���WP
|��N�r�f+D�s�jʧ��uՕ��K�͛�WL��1��X������H���C�~=<��f�OFi�p�h�p�8��.�B�1��F���t��y�7J_m�m�s�x�αr����wٰ��d�c��J>����=��W4�_;:����YX��� ��}G kg:��<};�lX��Ӥ}���s�)Y�DE�l�)츉ݴ�Z�7eM[�Z�Z7�(���h���E��V�?��ɬ �C��bop��0t�"���4�q;�#~"�����}���/Mc�ُ^
���c8@Q݃�y��\lg4�!;��J�{��h-w�������ܒ�u�@�KL�i�3fK�s<0��+`?|����s��m䫧s2�Ϫ�(`P�/���[l��Ô��N��ze�_�W
]}�����8�W>�9zh`ɋ���ʹ;�F�BT[i��	�(K�cp�{Z%�)�O�6 k0����������1��z��k�8�^�'���݀��F�
�c��:Թ��[a���E������4���뽐R5��X�_��mt�XqUb�x��U]��H�l���ZY��m�S�o�{Oq���Im�K���|U]P���3λ�3��3���ȱ�|3��0N�[S$������	m�R'��wqʶ&���T5f"Φ�#.w7b��=k��qپ.�5����W�J�r\-�h�tR��L��^�����u�S���~�_���R2obZ	�U�y;ޏ7��C�8�Rbons1�<�u7v�J�Y鎥{}����VS��m�,�{!�m�
r*���u}w ͤF��~���Mi���e��u�{�ص���\��+\�n���6�ڒ�D���K1���-o���#\���u7o� ��_��d�І�k���ǴH[L�����>�w�'�坥gR�y��{{��.J��2�����9a��tkZ^��v�&XY�g���UM-�}��uŐ4�:�̂wVXH�im��6�p������5��q��S��͘1�Jҕ���M��t��rޣ�0b��VT�]������3k;:���R +��W���2-��׉~�
�Vn�o+ٮ�Hz~��?5�qNu���",_N��;#�m�Z*E+sWK��o��_��i���IO*��{>u��h"V���#gu	�q��[����_*��k4��NI<t�Q��(&�P4˶�>�j�t�{&��\w]�����z�y[OW���f�����Ey�"�1?��K�-�|�!��z�d?;��{h���A�a���CU��hQ�jW����\<��uV���zU�����!�13����ה�fv�6���k&�F��"�g�7�rY�uG{=g��3��KkU���dR�B�����0�#�4��\ٗn�?l����uo���i��-��-Nɛj�
���f��ݗ�ug�p���e��Y�.r��N�[g��ߚ�C�4��[�z��qI	���}�������G�̣��ݕӪP�ARsy����5����*�t)����e�5�w�b�QcPU��F���úR�JWRɔˆ�,S2�V�������.}���c���<V��b;M��J�+���և��k�މ�.��{���휲N㜦���n.�ڤd�>��=oF��4N�ή���,k����N������E�����e���)'
dU�0�i��ʍ����z�򐰘y%r�����2x��w�&]�é[�od�ע�;z7{j�!�S� e�|�R]�*hjщ�]�+�'փ�ov��A7q��V�v6�'
�����j��dl*)�<N	N�vŏ��cjKk����
!0��l/�$�#��g�)��0��,����f
��\�J�J����C�l����E }� >#0���Z}�oX�u�]Ú&�%]�x|���[����ڏ��s��{��^�ag^�<=�X�I�9�V��c*����{����ƾ��p��P�f����&��` :&��'|N9ɮ�D�����#\����.��ܥa��Q�?�着�d����`��W7�9з��˕'n�Zsz��Wr�_�tMx��
�!�2���b���j�[�ֆf��L��階	�z��f4f��
�r7�©��P����=F��꺝��G�����e��O���7��.�R}�]��GH�l��$��\�����%�ؽ�r%��Hzp�fCҫ�:�*_WW�jv�4����Ӄ��,�z3���s���?��j���s�b=�zof�+���Q��JKfwt���N�;׫=M��ʢ�!�[-�.4��r�+��qn�
��^�~�:��������L�-���r����r̉;�-n�jڊ=֕�ogGN�����C�������b��K7үݏQ�ئ�:[��f<:�۸J��g���^K̻������ƽ�]и������G/����ٖz�};��a���FG@{s{s���*DXq��d�����]q�
Q*�影�W�[�s��=�++��=��Q�=�2u��W�f �*M`y���S��2oQ=&0�l����.��)�z'��+B�gGe������7C��u�짧(c�P۽8M��7�k���S�D M��Q�}�޹JB[�����D�ve��v�|;�$���E�4�l������rh�U���;�����޺��tEc�y]v�Y�p#-D�<Z������؛~�&Y�7l�r�:o�HӛtN��u��oDdwQ�m�"�:C!(����5���׾���t~�[��0�7�'��n��M�ꖾ�:b�i{���C<�i�ፌ�]�Q�{��n8/�T ��F{��A�X���O��Y�%���UT�#�Ƕߚt�;f<A��|sLt��������/�}8��]�[Y�C�u����2�7����,��p(���w���/5��m����6(4C�ޝ0�2$��oNP����RcY�E�g�T��z>lG5���s�m���8)Ns��t�o�G����7�~��lv�+�v�&X�D����-ɴ9�۔��w�4]Q���9��-���F6߰:e���[���BPTQ��P"�~D��*�H܅Re��юJ��e��4E�������r�z,���G�v:���ote-�C�4��u�EF�2�+YJê#g��E�}���ިdu������#��,�*jhۭ�Y{���Ⳇ���.���W]�U��|�N]���v륄����Ά*���ܮ�"v#��eCM�۩���b�M�}�gc�C��v���R2wlQM��6KF��ۭ��0k��)����k�]ٔ⦏oTM"�q#r6�u�u~�{��#Z�^��~ߨ��@���}[�2R =3���]o�6��l�p�l�w��s�yQZ�%,�+$o3	�_�vC�x;��6���zN\fߺ%�n0����>R�+�$�tNe%�-jm��g`|y��}�V^X�w��W��j����-�m���t��/s�m'�Ml����Eи2�j(KC�uyO�NCk�7�����OX\g"rtq�&"�N�A��^��[��857b4%!et���F�M�-�m��:���Xۮ��%��(�ju���F�p�E��2g��m�{�+q��
� ,��-V!*]9�c;y :��R�Uk�OR�D�%�Kxq��Ⱥ*�hs��|����]ќ��rڰ��R[�l�Zs��Z��(Xxv��XoP�0!'�ZD<a����#�oV�S���Ր�$�k2���b^+2"ʛѻ����=�zy��ͥ�ѭ�ׄw�k�:�9�`b!�����9���y��_Ӈ�I��7�M�L=�e��e�o"b�Cg��Ľn�9[��e��x���v^����=՝����o=��OE,��:}���w�-F�vpW�Y���먢z�Φ�!���Mi訾��P�AM(9\mmyY�+�tU�G%�����`;���[w5ZJ/^�	ex)l�ɆF������0�ڊzӦ�G��E�&CG�a���Kk8<�Ў��D򾖨�p��OD��-�]�c ��c�zs&��"
i��}z�z:�1~J�,Z�y������fY܀�ٴf�wx��^V�U��d���9�^��G�m��a��G�V�0��V>�I+:�g��7���k#�ۄ̷�i��c�Eތpn��[&������ZHL��_}��M���=iS���2�������S�+N�59��;r�a�]X����gd�,��R�]ZRCy�ʯ�Z�����F��Sw2�ǽ-��T4%y �î�`;����C���ʄ�Ǩ�zZ����u!-Ռp+ik�q��a��ͬ�m�T'�fˢ�#R�L�gEn�Yc��J�E�>�Ij�{Q�۬ٓk��I� �W��Bg	���y�X�vG?jɕ�*�M�sU��ۚ�z|�؋�m��؈��˺Db2�nҾہCV�x�gݩ����n|��篥�όx~�{��f�ςfpw
�Z�ZJ�z�=��]��%�dv�m�rv�H�*���Z�<�B����yvz��U�N5d�}�@��vgpb9��3�i+���$l�ʝdI�п.���]�_�</����Ov��)��ϵ/I�����dC���0���9�����n��6t��fe��NTLbK*��K'�5"V�1Q�o�ӹV����}�YmPSj���y���\���85��mhnjo77�[��kkkkkkkkkkhmmmmmhhhhhmj5/��r6�L��g�C�2�Zz��3�^nl�Zuq�����5��;:���[l�-4S/_x��׾�,l{�^o�	�fRqZ�\���A�xP��Ds|��-yGnr�lA�!߫Ȅ<���l,�wV���z��1�^||��׭5	X�a�7��c�@��E�^;,r|���i]���8y��>�F�ՍZ�@R�|q������d�䆦ޭ�EF�޾x�]T:7�)��mc�����������5�V)��"��M�]6t��=�
��b��!#��h{�nŁo.TH�	�nK�a%I��"�r��W����+)x7���ڞ��1P�C5,:|�N0[Τ�s/SΧ���#��(+ff�N�Q�D@���XkjL]o��|�<��:�ΘY!]�	v6	��}�wB�.-u�=\m7r
y9�S�K!𑢥�qV�S77�V��%l�xB�ަ�T�"�
'k�R�5�j%��O9�sj'�^�8,��{_P@�.��!���W��^�L���7!1؞�����z�贫V��˅,]>1 WU:\DM"�K����zzY�D�3[gPB�����㗶qk�ܖ4���}u�I��+L8(�ql���0|�,A�`�zOb^脞�����W�p��E^AO�P'�]���,���Tw��6ŀo��qY\7ک �2��ǽw�ₗ��5��歝���^ǞWs���F�T��{�B�`�Gh�QJ�	�1޾���;�M�A�?�T��]I8�G�7����Jr#w7eFB��Yj������3���^���Ym"�\&fVC��t0�P�5w��+���"Zr�Q.T�uf��U��2��T�7�UbƜ.�Yɯ��?KM]������a�����-{��p
=��M�p���W}0;����f�>"V���e�5���N\�*Cx����7�bZ6`�P8֎Q��Yy�������Ma��Yy"���Sx��z�4)ogn�v��e���@�6��[���y�RӲ:�$,u�(Bz��
u��Lh(��e�Em�;+�����c��F��X��;1~F��
"��;+j=���4��6��<Vyٱ{����,��3��p+<`����Zv9�1�[iT;��y� �h�u�.�U�y|F=��+��k���b�:ukt�Z�J��oHz6ڸ½xg
���etl]���4ZC�^������9��D���3|�(�\}�ks�$J`9��Ǧ.�5εt!#u���4�J�_����E�|f��Sa]�i�y�X���3����7��4�¹qMHv^��xy����������ߍ2�ܑ�(4^����]���A)9�njlcb�h9�������gWJ�����Gݴ��`8�ֶႬB�^�t�&u�C�wss�b�fE��_����r�:�����)~�����a�ݽ�ݽ��IE`E��!1!Z�km[m�;b�c{A=��uPGX��(� ��!���8��"kX����'m���w��ui�;8�e���k���SM�·F��E���Z��]�D��pmtsU����]h�Y�*��s;j>��ͼƩ���m�;g4U<C����U�����*7���ƫ����#b����֪�븶�(�"i��6N��Q�ł��!��]m�F$�ՍZ�UZ3U%wmAU"��D�X�q����k��������m�b�3�J��DEOckUUQDkh�Q���b6�	B��؈�Z���&J������cͺ"���y������uc4Pt�:[b�N"��`�Q���T�P�EN�h�P�]ے.�U�QUh�{�z֨���+F���gV�MFآ�*)��Ly�cA4G�����)���D[�� �m`��v�D�3TTQkDl���3_zHG�{�b�Upc�S]3�令 ���Z>ǅ�OVI��]+ ��9�e!9
�sy��q2`�N⭭x����C�5~x;к�z�h���$����'g��8AW�@�xk��!Øj��	�K⺌���}T�[�i�K(Ot�AYe.����2�G,|��2ח���B�㻷y�7�Wm�s%H�]��n6���J�K4J���u���p�>α���r6�
����.F��r���;3T������X۵/���w���py뎾�׉��
%�ͅ� �="��v���ڋ�~mr4��<��O�~��ͻ`�!ʀ��$�gk޺��Djy���(��3q�,��@�3Z��=e(1W������^�&��ѿ~�k��"x��ò����hÝ}՚��z��Ĩ|��V�sN.U]�O\z-DIλ���̘��B�������ɩ�~qm��d��>�(A�{ȮɆ�o78�О!-��P�ww���cC�*�����	tRx�.��rj��c�ث��٣<}eټ��>��Z��]���,]�.��e8osE4����$�f�i��l����/�Cש̑�����u�mZ�>�;ĺ�?C��$��T��%����o��؊>Zv��E)����:NwoC�͎����jJ�D�*��/3Fo6�"+�]/g��P.?����ޛE�>��~�Y��/���'=b���<�I�~�	%���N�cN X��U�3���yR)�ҟ��@s����i�3�O-���������ض�E,�t�{��ڌ�����[�t���nQ̰�QMSm14�&��{m�Ϻ�]�m�VJ��(M���Ħ���-��9�g#9��˼��c�] �7v;�,7�s�5��%.W�U�)]�n&2�W;իZ�沩kě���!�qhݴz��;�W���.6����������ݑ���q�1P��흶�w�k&8.�uŠf�F��F���5���/};�����N�{��kfW<���g�wY1�z��8�=-Xtdd��h��:N��'U �(ߗ�c�Yp�6Dx^�S&�\�b����ۥ�u��*}덥����?_cs:w���b&o^��|	7�ł�E��Q�م��'_�����Z7we�����৶��5��K�T�����<����g���3ҡu{{_lf�|C�n<}�
	Wa-w	�}�[���u�ɆC#�ٽ�;��h���,�O�S�� �2�� �t+��`�}�$�d�ף��2x�7���Չ�-��k`�=�=us5Qu�u9V�`�r8��"^�2a��$�pb�,i������/]6ت�׀Ϻ�4�9�!H�Ѿ���ٸ⮀����'jI솰�P��S�W{���{]�T&��yC�9��>٘
͋��[<��ò�.�y>��{�M��L�VxA�Rƃk����B�&Xc)�s�6krƚ�Ku��qj�{�z�c��y�����iW���n���<���[�!��?�qjW"1~�]{�Χ9����=��w���H��.�!��l6��W(���ԙ���n�V���}� BڑT|gT����X�E�5cE�w\wn�h4�=_�=&�N���]�1�Mq4y@����+o܂>�	Y�����Z�N��ꞻ����P#X5UUs���!\a�>��K/��i0��;��-� 3�nz)�t�,�q�����Y��Fg��j��$�]����cF���gZ�Й��8mwg�y8�l�̶�)]�_��wd���@�hѼ�=�gH��Zsj�#S�16��F��}�Z�c��9&�,���_��R�P0=_�17KiWU��[F��*}}58Ҥ̆(3��d��W^T*|_�n̹:7*YVwY�ܑϸ���JsE+��.'�n���4 �B^��-��kp�ɮ��h�5��Ƙ����(���E�1aմ�gV�/��S)�}˸��<��)�X7� V�����^
��~̟qY�31,$�vZ�zT":+y�U9� �c]�o���^o���\m��ZD��[�|3y�#�o.gkh>�ݲ|�\�J�t�rt�z9lO^:��ngt��{BR��O���f��,�w��Kvz|��<�P��/�v�@|9�e.~�Ks�9����Θ����0�k^{�n}�a���x[�]�#�a,�8(�E��a�����y��{�Q���-$љ2��; �k:�"�|C�쩽���>�U�ʶiGۿTb�j��x�k�<0��ez�/x���#��1]�;0t���v3N,�7�	Cfꈻ�����8�q���>�|�	s��e��3�Q���O3w���m�+��hS!�+$�F2ˤ����!۔ڋ�E�^�M*��Μ��:�bP+2�]�L9{�Ӡ�����8������o�I�{������^c��@����'/{y4��a$lڄ��OSY̻�hNv��{��E�x�Jj-aaBk.n�ՙ��l��3%�>ee�����^I���{��I�mB^� �zL�&�[z<�a��]臺ꛚd:{j۟{n[��*wcĬ���)K��DUs�7CJ�&Άbb*/��N�wS�j���|�u���4YU�
�n���x��Q#�SY̰��1e��Fd��>$8��9�^Ж�H�C��W�-�Y� ��I�I=��`o���Κ��o/�t�8�\0���JAB�Զ6��C�g�	͆�k�ܜ��=�x�n^ʈp�0�i�z���<��Ҹ���Q�r����)�)��"�;�c�a6�� �W^n��P�\��>���/��6��Dfxɸ��׍��B����奼[�U�Y(Vy�i�wF�Ci��Oh�씜��_m��?�x��$�(Z��G�`K��R�W)�)#.h�|*Wr_J�GN��:ޕ=��]���h��>�N���!��L�v���:�z_Qۨ�]+�6�dt;j��Z�z�]ݷ
��X]%����+��3��a��^6�^=������u*�oIp{ύM��Ն�罹�i?�O;��N�9v���1]���X��9�A��&ۻ�p8�\aIS��-�������άW���āx�y�8�mW{�>��ڮJm�:a�vKHs�K v�ږ���3�n'K�5�����+�͙���zA~-'�\��3 \�Y�;�8�=��%j��v�l^kO��M�o`���4^o6����ff&9�^�s��v�o���CL9�ؙ��ZҸ��&��T�y�g���-��a�c�ݯ]���T�ՌÔ�xt5����0*�潖��nB��Z�㷇VwCt,'mxg�iv1W�7�[��;ly���\�лY�͜�z������m�Җ-JT^>*���q�b����=W�7��x�ϻV�#sǼ�sNs\�
Xu߷],>�M��G�)�q�Q�Ͽ:�muݱI�KH�q�q��l�����A۾:}#�L��C�H��+��9��y=Ɠ�7GY�N,���yp�X��&�[9+�k�J����F��#gvΛJ�{
f����9a�agSnX)a2 H״y.*-;`��p<*nɖ[��2$
�a0^[����Ý&MDC5��d~U��	k�o�o�"�O�9�&�LB����W8����ަn��>Һh���^ɠW�'���or8.�j�,�o�Ͻ�V�ZM��u���Q*�I�n��8�й��NMX��?�pC?z��L��a��{���f�g;��GUK� ��m��C�X�Y۬Ycܬ�͋�S��;��ٯ��1WʨE�[�۫,$V����n����Z�����Np,顴ۿ ���j*��K��>z�#:��z��*Y�X^!4���{ӄ�:��}��!�h��L��\�zM���x�#|�ϓ'./��k��o�13�ϻ9�����e���		~�Kƪ(�)�����v�r�"ã
HD���x�W�^X��t�p�+Mׁ�x�+bmZ_e��vo[�w[Ő�H��/�#xX��&�9S�ΖT���)��GQ�d=t�VА�jn�	��#�H=y`��]=���4�'�'z�R�{�ݺ^V��7���͇q/wSR�5ֽ8�%Nx8�1T̤����&Kխ��&;��=����#���U�N5���}�5�Gq�f��0�LdCݺ�珖�������C���f|�P)�B�3F�u#e������L�DBy�'��csD����uщ�tQ�'�(��r����/�ѱyW�v�^w�ݥ͐o�/I��eڢ]��2�}|�eڂ�JY3���f�KFF��ɑW�^���D�:*�7U��k�'�Xe�8웭��6��C����!��u~�~d�̜pKz�W�L/E�*��,|�`������WR��2i��j��;�ܺ��*�T��%}Wyձ<n��n�/~��%)�㔔�x��Ç7I�c���dM�^n\h6:��=�R��!�z��K,��v�,=���~3�����蓽#s�9;��R���qU�7�<t��O1B^�2�'=&%�j��W1zl]��[�|�pK���&f�+����=�iil���H}�}0k�k��L�͙�K��-�ٙ�h�<��c�����zs�!]�@<֨=� �=�	$"���j���Oگ��k?�2�yꝢ��Rxmf��I��N�p�{����da9�Co3�j�kj�V�Cwcqҋ_ud��ұ�ʊ)�.��V5r0��.�J�����h��y��Tm=����u��}�on8DSGz��o5(�u��C����^�:g/k��ea�Z���qu�=����=�p�}aw>����$��8�눘��ߌ{D>�ó��oX/����1]!����s�+z/��>���R��ŗ�|M��"J7c�wN6���FR�4�(�V&����<vl�{={�j)f>u��'��ۯ5G�+�z�Ff4f�$�����[��yv�]Ͽ)�n�S�&:N�B�R�|^.j*�B1�V���1���J�V�ٚ�D���\�F�V�-~�R>�}V&���9p"�r(��}���^m��5!j�Km,���f����˧��ᇍs�/z�gF5����v(�<�ុҲE&��[^+2���V�As�����رE��7ͿV�~�\�i��V+����&�P�[��C���1Z9<�HO%bǓ�u\~�ik2s4Q�&q~g�X�d���ޘ��7��K�T��Wat͎��H�:6]3�h��E��FP�D�}�oa�v����Y����9%�J)�6I�9��AY�M`��	��q�hN7LaT-�!ͣ��*�������'�9���v��*�jX0�����Ա񦧻��������gw`�Fm�6�}��6W�-�#L�-�������]�n�k���"y������A:���e�����e|Q���s���Ϯ6�>�n��u3���D��(��s?v7��~�'�_��Ʈ��uW��=�2U۳��Q��X+nnQ���#Xs<�ܴ�#�Y�^���'q�l�{|��.9a���V��7aق!b�����D�f�VU��3; �n����3�� ����G{\wx��a&��Ȥ��������4�/c���bqSA��k\җ�<g�U}�N0����8�ԑ �l�#�<[�Qe9���]����'�;���U��U�{�^�Ù�@����,9�P���b<�A|MT��1(��Ȑ��(_���c[����>���������/��W���*��
�����?�H��P?� A?݃}��� �%�fE�`Y�f�`eV`Y�fE�e�fE�eYdY�fU�FaY�fQ�`Xb`e�f�3̃02�ȳ �@�*̫2,��̣0���(��� ̫2,��"�0,��,�3"̫0��3̣2,12,�3̋0,�� �2,���2�ȳ�0,ȳ(̋2,�0�0,�3�0,³
�0,Ȱ��OdY�f�F`Y�f�aY�a�&�`Y�f�`Y�f@&�A&Q�2.aY�f�`Y�	�f�U&�e�f�`Y�fQ�VT�dY�f�Ve�f�dXeeY�fE�e�fE�eY�a�I�f�`Y�fA�dY�fQ�A& &E�Fd�fE�F`Y�f�Q�eUa�!���"�"��*�a�P!�!�P!�P!�P!�!�A�T8{�8p �(��UV UXe eUa� !�U� �UV.  �VUXaUa� !�U�UVUXeUa�U�Cª�( C*�*�2���!���� �����0ȰȰ�0�����`X`XeX`X`Xa`X`X`Xt8dY�f�``Y�f�����?c���Y�DP�E I����?���������_�� /�������c�%������_����* 
������?� �+�?,��*���H��i�C�?�ꨀ*���������7����O�7����?>����+~� ���#*���D������"B(��� �*�@���J��(�
�H��
�J�,
�,�! 
H��E��!��?ޟ�
�Р�@�P �%���?��������������ߠ
 ����?���?���O��O��~����O?{�_�}������~����� U�ʈ�������aAW�P_� 3��T�����0�7��'�=�}|�<T@o����O��ب�*�/�i@~?�� ��O���~���z��C���G �
�_�?��U_����C���_��� �}'������ߕ?������~L�����*������2`� �����/��O�W�"���|`��|�D������|�����I���
�2��
�H�z:� ���9�>�3��oU%P��$�(QD� 	"�*���RD�H���jPUJ����*R"UU$URU**�H�D�Q
J��՚�HUJ�)E�Z�H[V�m��B�$�����$��*
�T�R�"�J�%d�(�*Um���E@�R�Ts�*�b(�tvD�"" �HP�+cU%!6�-�()#l�#LT	@�PR�EQm�%Kl�HM�ˡ�@:5Q}�E;iOY]h�   ;�״[*ҹ�]�v�:�n�]M��a��Mܙu�[+�dv���*��P�ev9����۷n띳r��t�T�����l5�m�:��q�j&�	UQB�
�mJ��   ��ж ��@��Ӏt=��B���B���(P�h 49���
f��׮���N��ҭ��m���h��u4����iʷj�:�������A��;Guε�wf���aR�֫�ԨBD�   ���J�wm]�����m����ݻ�*wj�\�N�U[s��n���ӭی�����;��8U�Mr6�;��إ�.��몕�U݃���vu����]d�U ���!x  ���3KRV���v)ΧtT
t4�]���;�n��k��U�5l��Mٕ]P�WR�ʳ]p�Pj�I�mvշ2�TTm��B���DH��  6���ѵ]�p���;I�ɬ�6�\���vm��rG5�V�ͳ���Jn�m�SQwT���V��Nr�V��'8Z��:����E%Vإi���  f{֎�)ٝ�F�ꎕ��&tv��9�#R�5WC\���X�j���s��Bj�IwP#�v����n�(�P�UAӻ*���  l�U:@rn�j����]4��Y�J�i�k�T*���r� C� ��s@ �&  1�  qR�ET��UUD�R�T��  	�  W�  k5w� 6��  R   mU`�3  ��\t m�.v  Z�  N�@��R�II*��  ��  F+��^�  1�� �, h�ˆ�ZW]\( @( ;p ���h 2t҂IR�Md��R"&�  i�  ^�v����X  s@ �` V��  � i@� Ak�� �%��(�S�)J� dh��$�� S�=55L�M@ �JR�  Sh))P  $ʑeT� ��[�Dw�5dc��w��"L��J� ��-Xz����K��T����'ؾ���UUco�痟��1����cc�� �6���1��C cd0m�����2h��`\Q���4s@����ai���)dwrλT��V>�\�� �!�t�ۘ��	Ҥ��X�Բ�x�]d��I�a�ӲF�x���=�~�T����-�3oa�SYY5�ڦ%��#������im-[t�Z��������@�yi&��S�¥n��	Tnڣ6�;����!�?c4K�eά�ʑ2�sF]A���
U��ynV��-fE�H�i=ϊ�1��Fc��hȥt!w�8�e�b��\�5F�8j�	E 1�ظ�"�Q˻�-�C�@WGc��eRR�P��,C�y�u��.d����R��f �a�<- �Q�B�&�U�h�5��v�}b'	l�������ʻ� 9�F�w6e��KC$MB��f*�巳)�����면�Ҕ��hMtr���B�}�:�� /I	*d�òz��,�Ӕ!0g�4.m�:��KpƄZ� ��� 5fe(���.���U��O�������T9��'�vk�Ǯ�Uv��2nY\Nձ2j7`�l��njݬ׵������:a��K�M �[ttf<�{��Є�A\-�Yi!!�f���M�n���]ϬfG�1��C���.�H�.��Z�t	a��[hG�MV0��S�s6)�ܖ)�Te�Uk)r�mM�i�%I�Z��k2�ӱ��mm�c/n���,�A�g;u�ڽ%;��DR�@bԭTw��̺��w���lf���2��������w��G\QƎ*X��n�0BƧ_�;X)�ʁ�MǓ���]+�2ܥCnY��],�nSusvZ�FL�e�Q���Ԇw{-Q��ΈUqV�B�ʺWcmB�l���%�RM�������ҵ-�*i��]n�E6��� ���f�t�U%�zJ6�X�jEB��U&�^�6��.��։a7PU櫈^<&m[�Bm��c�yLi-$�U�A����
7n1Zd�	��j���#���6f���B��y$Ln�nj\�1�*�l �7[Yyy�\�4,�֋l�E<��^%�a��J�◎�#�[�Tf�*�7��Xr�	*ĉg`qH��-���a�#6s(ǅл5���%���F%���oNX۲.�]��V�v)�ذ�Őbj+5�Ɲ	����e�QEhj�@�#)&2�������u�=N�8��wA-$j���̨Z�/q��|_>��2�;�m�Q�{07��L�d�e�j'���*u���d$���4�u��Ɗt~M�ݤ�E�);��eVQ8gVEi������[��D{�dpաZhSZ�Ŧ�V��$�x�p^�������ϝ��u N�_�Gn�m��M�,0&��UX������gsN��]0%�q-�I��{ Į��5�t��6���l:�u"�;��GL�2�\y�:I4��z.�����M�9��q��F�S���l��"9���[�ehVe��3uX��pS���Ԣw�����1����$�b��#Yi-�5D�έ8��n�E̀V�7Q�
�k�Ƭ�QT.��,W�c(Y2Cz�AYaP��/B9�nJ�h�L��MVd�{B��[�!���޺�b�2�]Kj��J�Ȑ8�:�NhU�t�t����5P���\�q-�DVM6d+e@��������υ�vp�ĻY�X�qȦ��E#4�ӌڸ7^��+%��2�n5EU��A�B��cR�8�*�R��w ν[lS�Q���Gx�W�R��M�n�XŨU޽�$�*�hR�uzLS��k��ZQ:��[�� 2�XX7P���1D�ȃy���7&��)Pغ��B�yu�e�n�Z]�\;e�X��Xh۴ь'���n����;���Ed̀)Gz�n�1�	EK�f2S�"��1bYue�XH�5B^�%n*-Ďm6�ɖYO �MI�6��'���M���U�u�[�zTXTO% �*FK#���n��u�J�­d�`���g��$1l �(S�x�hZ�w�5+l���\�X����<j��-�I��kR��^"֫6U�ߞ�gVS��N<BP�U��PX�] 2jt^�RX�ZjVG7���Ȁה3N��MFt�q8�jV��چؖ]d!���V�u*Tӱ��\�f���t���@�b:�Mk5�֧��g ��4���v��tX��ua�j��Woh��ROV��������i�n�M&˧业۬K��+��V�*�*ʽq��M�9�L�unS�X�� ����,ckV�A�KF�/,��`��Ej�4�4kT#�i,��[t�QǀIV�i�l�+-��˧��AOub�],T��G�rZQ�@iwFF2nM^)j���(�0�nŹ�vDױ�7�ݫ�-�q��a`��`ڥ�EM��&�5h��Ң��O0k�д�l��jk.�V�mg��-IeZ�R! �`��͘ �V'��wSt^���B�'h�j�^��@C��T���̠T	
qkJ!��M���:��n��v��&n�ݒ�k1�m��qTQ�78.�1x)V�����]��b�y2&ZX�9.c������وǲ��Vn}h�GU���V�&�6Y�Ny��[�^��g� :E���Ѽ6U{4,�y��ߍi�CtZ��U4'�KȀ��������t4��̓n�� ު��v^��%Ӵ���봞_�'��"(^��i�V���+mjJ�*(����ӏ-��l��(��7Oi뙉V�W�ef��&�Z��!@�M�I7��L��RQu���a��MZ��ѓ.j�W�T$5�fk��õ��[e�w4�V4�8�`-%J�ڸC�IAP��A%6(µ�n�t�;9yYQ4p�b�Sl��pT�5��F,-�n��ӃR�'�������r��ђ�R�iW��eU�u�m�ۓ#����n}jڍ���;{�V$-��7jH[vM٤���7a7�K��d'3,�)A-L�m̂�G�7je�q�ʴѦ��gv1 �X��R�I��F�˱v���Kfn�,T4��ݦR�RM	OK��i˶jU��6���ti��-g"71+ù{H�U�@��^H�� mݹ2���X׵�H8�kܗjf�`��L�=t4��A,:�.����1Yz��Q�r�Q<��MV\zՆ`�r��D�K�0���6�-j�+���l��P�r�'{pҩ{�pb֫V���3V�j�*ʳJa.�X�}kE �^��8+E�F�r�j��TIKQ��r=�	N�]ƆC�2�Hq�f޸5t4�"+gm`8�Io1*��Ա#T�Xe@�Ҧ4�B=9�h)=��ǉj�.�M��-��h���Żj���h�ujǢ�t��eE��Ͱa
�[gyR�p��Q�vS�M`�O1���GK3tVC�@�T�J������f����A��Ld!��Sa��k����Z�B	��9[+tۙ򣰡� ��e�vFD�� ��Zrڬ	#��r����b�`2���cv��ō�0B��`�,�2�nP�ĭ�j�Y�z.�\0$joUj���7��7_�@�+cj�j���ь���M:��j%`fZ�mm������:�|�ս��QF��mڱ"�q^�<���B"kUm5��JY��	7h��5l�ܛ4���0�Y��Xi*�"�`ň8(")VF,B|crV�W�۰,�]��Q����%�-/��9�k�R]h��#[t� �m�	;�P֕:�N��jбy�<�	];O.^�M�ʹ5�l�t��q�6jKT�雁]-���M�bS]7S^���$�r]ܗ��te��.��J¦|��ʆغmC�%D.�Ŭ����Q����).��[�YQ�x��s
<
��]�)Q�'%�"�������^�M)����$�(���)E�a�|�4�,S
 �FO>���n�Ѩ���^�{�pǮ��.��3p�����eH-��݅�Sr9kl�c0�t&SS!�T�@�{yF޴��p9s5ެ��û�Z��J����J՘RO��m-�����eMN�>$3ko*�z��m�v��(Me�j�n䴣�m��C@O�3�swD��}�Kݢ�I�N�����`V\�غ�&HNC"�d$]=1�H��;uN�B�U���5�J�[u��[u��=�^+��B㫎b~3n!@e���)Kq9�G��$��6MwD�ME�<�6X���!r�)�+w/'r��x��v�B��Y���f��)Z������F�i�HeD�b�1�37Y�����*���o:��y�ewP4���r�Y%�Q����r�a� �j�cK�e�#������W���ڶA����if�d����[�t�V��L�n�V;R#*]]@���X�ڕ)H��`�����Цr�G\�0���v�*�*C�fH�l��eT�f��V�r�=pd+v�Z�x����X��ؐ(їN�:Y�uV�W�L�κ�M�;��ͤٲ��1��p� ;$�+�t0�z�^���rV�ٲ�a
$2QFw�%�wRi�M�mR�Vde�Z5[u����V�`�ҙZ���Fl�LZl8��R���CP�#�]F��(��\�70�/d����7M àb��=��-fe *�5��0��n�-�TAc���R@im��Mû�͔oE�i�%f��d�!Ƒ�E�d���6lm�F��v豚k\y1@��tU� d܀��Z�MPT��6�����4vcְ��M��j����Z!�z(��tQ��ښ�1�L���F�V�!jSI�z�;���1�L�5��������@�&+uհ��V����:U���kq���5���2���j3b�)݂�ͺ5fT���'.j21�j�x*��If&�h�E�4PaW��v�#���)Vn=3Cg&DaC�5�^:Z�"@&6�)3�Έ�1l��f�@�X ��`��X؈��VU�-1e��Z���c�Nť��V;#+r�ك5�6E[l�Ĕ�a���T���&H�)�t��$4΁iVRU�/��E����(�l���"�rܩ�Iz��07F�qMc(�����PGLLݢ0�n��ҷ[� ����b�f,��
�X��&7	��)�1�M�u�m�N,,O���Z��cĪ�V�R6l;�S�"'.fEWx����ʻ�+5Pf��T.S/J��f���K���6�m���F����iHwv���:DJ7t��)RAl'1	ɔ��n�`�Be������Lw����qƍab�a*i�X*:��և �9�{.T�R6[Yn�@1-U�Z4!��	ɹNbʼ?`���[��uwWӫܩ���*�U��13-�j�՜��ř���a�tf���R��4sU��Q��z����ˆ���͋�mn靛�e+ұ4"�Nܪc"�XH@*b��c�U2�~��}4��kC.�,�k�"�TyD�Hi���ɑ��Ӭ�f�l��Z�v���6��J�����Em�hf��`˰��B�`��u!�yOj-�m8ʻz���jj~+�l���m�uyOm�fb��SѹU�BME����ks2�IJEH�Y�H�jEnU��49j�P�Z��Exm��a�N�O^��]�{4��5F�x��]��)�[�8�[YGlnU��30+�P��H����uwV�&�Ԛ���q�[��8$��Fn�fU�dfVk ��ePL�e��X�{N������D֙+V��r��Qr4p�,��J!��n�哚�81��%�Hb߶�Sp�y��
�U�R�k:�t�̶�pU�U�Ŏ��� IW �b�Kn�!:�J�{�V�J3V�	����n�-��2��W��5�I/з�7C�R��3B�f�'�NT����b6i���a�n��	w)FC3P܅Uե� ��ۡy&lYWN�kxC-[W`Ja�#ÿ>����w�_�7+fʃ\6����+I�]�ͩ2\X��v�"�V���־�`��3b�^��ݠS�Z(C[r`54%#�9v����v�n�Ơ�-��٧B�
��kg�Lx��4�M�T��bF�c$Bm���^0����q3��3kj�Է5����ا������½.�c���Q�L	̲r���F*+[
�]�P�[ E���yF`�7�)ۦ"D��E&�TN�a�wT5)w��3��f���v
�'
�z�ƣ۵����M(%Y��(h][�%ͩ�"�"�9��P�Z�k����
�K���jRԘ�u^(��� �)n��3��/R[��76�֠´��Sс]c��v��(�Ѹ��ʃ%�ae[X��,8�Yv��a���i���ط#�R��i;"�&�VR�1 �g4}�v �/�-�:6�髰`1i([&m�R���Cjc�ː�AU�:U�v=�"���a&����ȓ�����mn�!��J�[��c����8�Y�b(��b�JS��j��JEȭ�e���w"NV���tȐhD�����{��j��[�p�P��Z4f��=ŀ�.���ʃ+%M����Ffػ��=�h�jPTU{��]Y���a��iB*%H��GM���+lO�̓f��#�Iǭ�v�b�e]p�,��t�V3���N`46�s���S��=Y��v0����q�Ȟӥ��9���&��od���;�3=�c.��}mL|�R����v�f_�j�Z�Vq6�D�c@�v�fТe�O\���`�P;�Z�f�r�.(^�t�Vm�&8�Np��U���2-*EZ��{�^��7e���Sr T�jC��F;ĐS0�Y �������xlٳ/lZ#4�R�� �@IC��WN�^bD"`jTuk3�Z&���G��ڱ�]�w��;W'R��λ��3x�r�qe�Z�q�:ƪ6�k�(i5��nK��j('�s�]�	���[q4�O�1W)/���Q�܏"H���K�6�<��m�l���YS/m�:Z���7��A_q"���#4���C5����!�}�e� �t��-]�k�qZ�8-�.�k�ޞ@ڗ\�LguZճ�� k"�;�$w��r�֋�#5���ڨ�T̇E�ϛ��d�7�0���\��nҬ��n+�U���H��Ί/e��t����պ�eu��Z�vZ��Y�bf֝�����X]�ȴ��T' z<ˁ�ڜ��#,T�7
�?YtV�N5)���5^-ʪe×9LY=T�w��Ҫ�rM�&EF̖{���#Iful9YK���i����o%�M�N���i��cԓ�%1�+����F�=8/ZX��4z���F���y[2�f˸K;��̓����c�{<��C}:��WFw��N3>f61�L��5��k#T�cy�pul���]�����Z����Jf�2�|O�g�c���x����eŇ1���^+�%o=u���{-1sx {[���j�9Tz��-P��Xo��ʐ���[�r�F�⣛דx(�N���m���Q���r�e�T��K��V5�N^+j�2�`�rd25��c�r�վ�_+�vFM��[g]��:�#�
9���T+]�('����{,!K���\�r��f��kɴ��Y$W�t#�K�d
���]����v���4xН�7iP��[W�q�g==�����7��۟mJk9�ͅj���}�0���˸Z"Gx��E��	��C^��t���iN���XG�J�k�@ҝ��>��L7S��i���ʭ��ۻN�a<�������%f�^���mi�O!�Z�`Re��V3�e�m(9�����}.��LѓoM�ǺÆ�>�����X�W��Qs��]��'9���`1��{6=�4S�a���n�V���=]z��1c1c	]j˨��d�]���à5>��u-h�6宥���ۙ;�4t� gcW}�rɷ|�����ʍ���S�F����وQ[)�f�� ڻ�mذ6Fk\��]�e�+v�-��|�S"��iw���݂
�0����Ld�}nv:��_�y����J!#���:=|��fŃl����eH�F�*�T�ɇه6�gu�e����k��0�K+�6��;n��$��w۔�*�;L�Z��qR�'d�l������C&ܙ&�3]l
r�P;�	1��(N���;�e��C�>��n#R���{U��@y ������
� m9�d'X��ܹ�+�xn�`Eu�g�]ԁ�ܦ�Z��x�n�Cz�y6�Zh��n�$��}��a��nńY����ծp�@MĞf�a�(7R�2s����|�Zo,gYr�v�p��y��5�����n��'j��Xlr�����V�_,֩��8٦̦��Z:�V�3Ɛ|�n>f�c�4�U)N�k��[��B%�f;W�W���;*��0�Ik�O[=��p������Ʊ�lt՗qu�������*�w�mM�\�բh�����1�.��s:`��F��Lܳ9$��f�Dn;y7mR���AЁ�h�w=�y�HHs�!
�ͣ���'l%��sh�t�����,�XfMmk\G.Mٳ;���H�]�ɇuw����*EE]�d�}:�^�ԁP�g�՞�`�o��g&t�J�|�X+����O�8������ad��C��$��N��/�a:1�ws��n�:���w�a.ٻ����D-k*�/e�F+b>Hed�Z�U�x}�w�	���qp�R�WFu�|>ݎZ����t�PJMIof�����)kTiTWV�{F��.w��&mG������@�וe��Aٖee�[1�rhA�����4ᴮ(��u�b'�=r�.e v�x=l-t��1Y��g Ѕ���g��rM.t�����4e�=�nm'��^ʙ�]�F�m=ʴ�Nz1b�=�%kO�n�g�;��(��w��:���־��鬡��R}�cַOX�Q�`��|��[��p�^=�|�ђ�*����w�-\v��7	=Y�p��W�кgF�:�h���)\w����ڎ̤��d���(+�nT�8E���J4d�UI
dK[�Sw��5a078A�8X�ʴݺ=���U�C%s��rQa(��Z9��mY�ʢ�T�.p ��y�]q5��S��8t�����FS�I�\D�N��CB6�Sኤ7b�ee�P��Z�5���ho���JkB��H��Lf8w���`_L�r�D�A�k�������I̺�f�^�e_i{�Z:�C䃮b�j򮆬o�(u�o%�(�V�7+�>u�CIP��x§^���sɐJ�Y�q����JU��T^o�:�lH<4��7�x��m��'����k#��Dw��2 1��6��ɩ!�����upfP��'<F�q�$di����ɶ��L�V1�\�u��A*�����(>��̾yiλs�� v�"�
=�@�v&&vfv�sn�����Ja���4f��Ib��S˒j��I�):������˫*�s%fb��`�oN!����!��V�)ŐJ!�nX�<� ���묾���0%&�V̔a�6�����U�F���"p���X��|5���՝BC����*�'YF���KZ�A�d^��N�z��S��#١�}�^�'ئ\�q�MN��Y�(�J�Vt�BD�e1�__j�c�t]ώ��]�<� V������[����x�}�on�DRܴ�ĉ劝�
���b/���W5�$�դ�ԳNJ5����v�\���n>]`���S?>�U�5^-� ��OvNbv;绫�d�LE͖@�,��!�!��r������g�V��mhHwvX�.`��e���OX-�N��]C��s�6R�̈�zԉ�x�����p���<j򾮍�������66�l��}��b(�q�#�֭t�Pn��|��+�;���4Ѿ��ʹ�4�m���U�@���C}�ky)�W�u���;#U�wh��k4b�ړmr}���j�`�V�LJ7u�si�9��Q���a��Wc=b����,�*���	'e���N(�N��[�Q
�*쥣Bµ�f܅A��%����;��.}��tv�ͨ�3�Ӹ88�>|lU���4��[��^eJ�t�t�nYnF�V*gu�˦+�'��r=�g��LJI6y�#�En�#-���g��.��u+r�4�3۔���_S����� ��[��71#z�moP�ڛu�R	�.(���k\�F�a9�4���.���#��o�N����8�U���u
�5Z�y�����Z,3L���r�f<�������U��a��(�s�2�^?���ٙ}.1B���,�B7��f���\�4��˕��֎RV�;�s�9P�я�T�K�����8��k5��2�gӷ؛���ĀWd�g5�MA��V�q�ă��`  ͂Q�Xޑ���x��Է��]% �(�e ��U��*ݗ���s��g��5��!]%u��7ͬ!g&w˰Q��t
Ti �	�O��بoh���IW*��n�Yq�ܒع����^�0�5s�m�\5���#��%T�����c%�Yܥ�k/uMA�iX�9A�c�4Շ!�h<�K������T�[���Ț$[��x���f�Z���]jd^�f���o
7]Yf��{���wc��B
qvJ��`��54�2oV���g.
��%��,�ݣ�Բy��䄾HI��A���n�u�б1��j�I2�5�a�5
�(���XBjxz��T��}q��!��7]�/dH�'4�=+J�+L�H�}�3_��;@�E��m�T��EMi
Jo,fZ��2f)��42��z#�0�6��Q�ò�|/�r����M٭Eނb�;�0��v��U�ҙ�W��t6�V�Ø�b�4e�=.��[��H>���+꼜�@r�˫x��ʁ]� |T��O��|p7Lp���������/��,�۽y7í��Bh�Zcr�F.��,�b�v8����!(ˆ�$��S��o�u���7g����;n�اi#���n��Z�U�j�'4��ұ ��&U�+�Ӧ�;Z�/ZH���q�k(.t�]*/m��`�1;�A_vn�|h0֝4DX�T�
�e�v�o���.<�f�e��s[��^�r�D������P�hT�{܆!��2\[]}Ƭ���ޓI��LV�ӳ[]tD�or��5gdE�-�Y�Nk�Xy|0�sL��0��X�NӉ��4�W���xg7�3�U�ԙ�{#��ƚ����Q�{{������2�m[��Y�-�A�)��ך~5�'R��1l�S�6�Z&;�;xm[��eVR�AB�E�K;E�%���Z��4��fw��<L>y�S=u�q_�ݽE��]���\����u��9 ��Ƨw��Uq�
lkk̈́�{7n {'W[*w;��b��֝Z�c3���4 `�js澝3B>��a���bpFF�U�#eqՍ���q��B�g0�v:�u�����B:
k����quZ:��̗4�5�T2]��h�4��6�3�oܮ�<��E_[xs��rs��hRu:
غR�<U�#��YM�k��J��fc���+����(N;��&�k�N֊ˍ-a'@�L�xX!�Rd�P���DR�9��a�Ɋ��,��%�z�-f������%r��N�[��%G�c�=x�K���/�(	F�7˗NU���\��*!VݪsgnT�{J�âQ�h��epAh�i>�=͋�4a[���&r������&���u��Z�%��R��/�P,]4��z�u��:�f3�7��C[�܃���xӮ�O�Y�J�ص���`��Gw���-kHHy>���QM�K����^�#ZR�h��M�㜆�=��8y�����ږ(;-$�>�E��h���~��Emf'M���8�EJ�[/��`}��^T\sS饒�K����G*.�+�i6�\���a�C^b�}��<��)����a�4�><�U���ϏL��}��A��@c���޵!e�G�d�8]�^M�M����v�X� ���4����$���������{��T"�e�!Rwn� �*h�_a׬_I�@��嵘�k{U� ����YҮQ�6�}[Q4�e����\�B��SB��4i���%��Y��I�o���C����E������u�K���\��MD�1ְ����tc�'����,�ʙ�5XX2����̓��(.<���,o�S�|�@�U��C�A�w�U�� qe��'}�_����$X5�J4Yo	���,T�����9��W>��U�Pfm�c4�8����'&Ӭ�p^�)�&˅�A*`'����r�/P[�Td8��X�=��E;V�v��Kuub#Tq��3�JO���œL��KIM��V�6�\I*Ƴ�G	i ��[I�X&�;��Z+��� �7�#}f-���`��{w���cPp�sEh�(El�L�ћ�D|�
�����$��S٭`�`���l �DV��������-'�͓�[���Pꙮ��ٯm[m�tQ[��!#���z�|4��+FU�o�8)��q���GU�yt�	�pU��v�����N�ˁz�ū�f1(%R�RF�?�^�to)���so�l��p�|�(�ʺ޺��F7���v�v�1>�k�#1��O��N붪��+V$Ӝ�ٲ��&�t�u�����j޵ū8���:��z"w����9�݇0�,�̗���.���ə�Y�śQ���4Fh��s�A�ͽ���w;2�(m�����vY!�f<�[(�ծ-�G�������-��1c7M��f,�u��fr��k�t�s�i�G	���ެ ̤��ܚ�P�f]�Cf�qX<n��q��`�
ވ�ed�զ+�VГ���y���>���Ya4'��ƚ��o�6�O-Q�+o���
�5���TQ[�	҄�q]�VK���K)�@�ޮ��lTm��=B��r���;'�-�Ҹ鼗��;=��O�� �Վ�-z6��4u�:�5��S\���pb�d�y{���8�R�}�M+�j����I[�Fa��R�w�8�J�*���)�/�j&,��֙��#Dv�v�9X�I�g	�T�(F�T��=�sOI2���%�L"��I#eZ5�	FV����o��Mz.�ǁH�Dx����w��ۣ��j<R�)eط�cͷwմ��QĶlƾu� ���
U�^����J]���e�i��g.Nv��<��<��@KA�)�;���f����(x�EP�0]j�-q������\���;�ؚtk95ch�L^��Cu��3�W��ĺ�}�o:��I�r��D�;�ܢ�q��s��X�+]b�n�w8�;����91��dZ���]%IK�����壇
��UB@�2�.%�wNYktn⋬sZz���tq
�"GG�=�O9}�M �}��|�z�i=D��P�s!�Rަ���v���}{ljX�l_U����fZ�.6.�nĥ��+_p�k��v_>�I��1���|�(n�,&cU{M�ڛ䗩���
�7��[<�H�`3��ם��e�;9���h�<����ՙx>�WD{�@�)���mG��'+;�	�"�L�s��ݬw�ʷ'L�0��s�1j\�K�ۜ	 XPD �PH�S���˗zou�8ӳ����2�f�A
a�-���P�1����A�[[�LĤ91%�j}�~ {����?���}_}���kG]�>^y%8��'�$f4��p@���nkv(�ܮ�p�nM���]�-�	c�T��sm��ܠ�[I�̃S�s�]�7��R�G<�V����=�A'0�U��0��\;�5��x�|�J��l��M���|��!}!ꛊ��Tm�׭�A7ۖ��5m�d*����<X����WgN�Њg9"9i�Á��Vo�"���9{&�Ӑ�����NHy��	���u�hM�^����=�����&�˹���ڋ��o /8�l�t@���v���', �&>�ծ�v���\8�#X��2�f�reu��u�1�b�:8�h�Y�yPWrm;ܷ����M��	�����Mf ��t*�d��U�M��$Q���__�Qc��3���qieK�­�`ai�9�
������Ha���[��ts0�/)�X�;p�(U���aW|NC3ozК"o�!�H�(6��&(�1J�)yjX��!��h}܁mެ���[sr^���YuW��mx"�E����aJ+6Е�wl08b���U�9"�.;+\��#��
%�u	�r3�V}@�;��r,��K5���N*#�R�}>Z�E��!v�V;�B��}˩c�ͺ&(���	�ӥXOq��j5b� ���@^�����|	�,e��h�`Ā�y]E���������1"t\���B� �t�2t��ƈXF�@�$��Uz�x�`T�T�KyZ�KF�#�bWj+��BQ00����cv�À��J��mS69��:	�r��\�ب�7)��*���vuE�,�q�{�d��=���F��Hm�J���?q��"�6 �93���V vU���0�ZQ�갱qlCc�#��w[�/�p�g%W� �K�]0�T����utxFq��Ɵe��n�qf�z�2��X�XٻXT{��p�g�EQ.��N���k1wGw�7mN�&Y��r�N[���A�evZ�e�e�이㵕���X쓬g:�r��Nٝ�)E�+�.��"�8�!+��dK���6Ʈ����gbΚGͱ|�� udt-ҵ��T��y)�*�%.3��={����������13T'����Kf��v��fͦ/:_*��cld8�L�uִ�1 �o�A{����:^w9�	���7&��Tk"�z^�J�m�弴?;�~o�B�F�_G�5`�]4����m�aLmp��*�6�4�x���I}��L݋�z�r람���\���u�x�� .=��ژ�e�L�
>����˭dc|�=1'];@�[����c���W$������Oc��)�����ݠ��inZ�Q���Ǩ���+�[ETi D�_פ�)�����r�L-�Y�%�����B��yVw�[ͷ�Jt���륗MIf=i�U��f1��kyzl�uh�� ~ӻ����]�X�����$R�'t�H";s�`��Mo7��f����ٕ�">u�#;n�Jܬ�%R'	E\�2i����s�'|r�;S���D�T]�QI����VW^
�=�핳&u(v�N|��]\W1.oU��R�Xa��q"����ܾ�P���)WF7���Z���.��2��o���ń��[m���Mr�W]J�P�N�M�Bx����e�+ �i<��Ȗ�r�C��.H������c�Y�B<2ֽ���}���Jm��'z,;���U1���6Ը�+�r�Z���F��[����ڊ���"&P���^.��'P��e3ډ���L���り��D�[��<n�actb��SQ9��'Bl��wtm��Dӆ�j�E�V�mӥ��vM��m�T��'��|�
9t�]��ͼp�oqh�ͳ�DgU�M�XHds�
(n@'[m�Ѹ��.��놝�WۣG	�X���*�A��6��:�]�kZ(b���.�ġۂ��n�����m�Yx˔�����n5�qu����1����I�S=��0��P�M]٥S�LRc�2Q=�	�3+���p
��z�!�s$����/���R�la�v�j��$sg	�m��C��kJ��8Ҏ����o��o=�*��9(.�������,���N��G �ݗC�L�-i��i�؋я���#��RX�O�\КT���2��t��۬�J!u��zu��KImڸv� .7A1,�5�o{��GY%��f/���ݻ��;C��
�Z�3�G��n����R�n���푧��l��ǪB,���m�ءL)N�GjʍdYVo؍����F�onX�� �!���,�X��ۚ+�Lʎ�I��2^��N[N�h(�9G�x�3� Sޢ����Y��O��EK&շY�BC,V2�J����K(:�O�چ��@�WfU�)K�b� �Vf � �9���cв�����`$���qd�0���T�U��d%�6�vR��^�#�杚"�hue���Mtt�:�)sv����a#��S�Ȟ��k[��qd��D��o�nvj}� ��ov�!ր_f�t�36e�)��w�Ja�b��U��u�!e��!p��2��4;�aἺ�r�f�N�p ���J	�����[��wض=�d��AzF(kii��l�®q��`�ܶ�"�W*����������&���n2d�oX�d}sT#ŝ�yõ�.�b���q��s����Lϣ���B�N6:���*l�Q���y�;S�rz�=��o��Dݙ*�wz��p��Jo\HSOC޷���1����[2'�U}Y	�;9O�Mv�_Ov{�뗳�,���J����c��W��@�ݽ���*6��gV��F_\tC��jP�R�WN\)v��]j(r��f����$��E�k�y �q���9�Y�N�x�
K��k��kԫQӥ���E��oq<7��7������E��.��+w�u�{h�� �ʡO~����油���;��	8G9���d���͂��f�q�ד�5�K���=g%�׬�W�.qҖhV��T��0�d�{;�2c��۸�;^����+��7	�L��DݻOR��7�~7K����6��E�vWJ�h�(�Ť��YmТ�+#U��{���dv�K�v��'�3�,��2))z6�}\;ǻ'��H��/���
ھnR�K�G��u}���a�p�NQ)���Ԍۥ.]���&|������Ѡ�6EFbfg�hTV��gL��6������l]\���Kl����<ʹ�"��l�痙�ĝzj�I
ڹ�Vv��Ty:��veh�!�3���u����}}u2�ӹ\��x�H .R���t�!��]�_gd!qQ��^�V��w�,���+9Q�ݢ�,Ll�]�H��x����M�Z.���sz5��&����
A��x�F��!���1�WR����	�y�Yt{���	�4���E�]5�V��[W��]œ�v�s��m��Ђ�e������z7�ZOm���0I����w��l��/�O�f�r5.if��U�w��q���LB�d�c2L"��W����2��e!���.��S6�r�|����D��&�E����aoi�L/�7����U�h�j��Λ����z�N�U���ݠ���KzJ��*��H(豴���]�{�mwV,��,����B��
X���t�]n�_f���&�J�r�F�l�LFXǖщ�]��U��!S�7R�@r償Z�#�"4�5Uؐ5�(�;�̬�Y����v"+y�9�i�8���R�[���.�}�k��n���nK<�oC��e`C��w���Q�QJd�bpv;pi2�mtW]L��2�'�]�,Q�!���b���bJ9�if��I���1=snY�g�4�`w�7�����2�*8���L�8�O:�ʂ�����j�;��e=γMɷ��D�o+7Y|���rm�9S����e��e�,M���A�-$:ˡ�ota�@b;Z�=g�E"b��&�0�a$�E�Z��Mц��VR�����B"�[qKa�ki�3-�AkV'�L�|��;���HǮE]����v����d���І5Zd�S�,X�+������[b����1>���Jr�(��� �V�v��W*��~�I�qfV��r����bzq��sc���4y�5�앝)Ws�95��I��7������5kP��h��k��F.�jp�B�m��oL���W6��8wN0��o2�}�%$��;q��N�^.��V�X����eS�����v�`�X���Ю�r�*���8U��ܢ��'k(�b��[Ķ��P��`'���<)j-�+�k5p�ȣ��ܤ���,!�5�66�)����Y��;d�����I�����L�^J�t�k�hk����+�Kk��X�e'��:�U�-7��=Wø#Y��u-K�\�s�V�8YZ "���hy�r��7VC8V :y�qѶ�VЁ���w\iR/�uk����@mې�u� Uٕ���J��]u�h�đ�/���J*��AET�&�Cm� ��gݔ$�r���yY��݀r�1�Xʑ��J��q�yZȥuջ�T"�>�-�Wu�����G9YfP���!v��Ĳ��ۆ:j�%�����u_n��ܲ�C�[�¶�[��N�ui��t�r�[�����{ɝN*�}}rh�+�;�su�o�q]���L�p?��r���b|v\��4.Н���(+�wk��Z)�P�}\���8�� �]&jY9wT��`Q�:2���Ս�75�l2���4��[B���2��������ά�LV�\��ĤW{e���3T�V�Hf��}/,J�k<smgDl���cAt�f����v�ÖX���&�̗��J2�L!�6;����,��]Am<2���f%.�2��f�i��7T2�J\,�Y�UX��cG`�o�vNU�\�x�(n�ɫ��{͞�H�QmNW�U���ܜ�u���c����k1%W��I���QL�+�������⧰=�Ҕ�!8�
Bu,�U.j(��W}zv�ë�Ws;�Q��ġ��ZĖ���.d�lf�F�RҘ:|X��%gur���D���Q��j�+�CL�e��r෇]5V������Kz�*�WrU{���
C|&��S8�������:�<�vS[$����tq��q��xǓ�`�`�V{>#{�uN��F]s��m�u*�B�{!��jY��:�Nō�xs�b��)����%V�i�����I�^�-#�.�*S�zc���r�;&�kp�EG�w��������򭑫4Ú�U�[Ec��\-J8�b<�%&�V��=I���*]�*\��,�W^�CnTUl���Fc����m�.௢�\�'����C('YS�:�lj�f�u�}6�i��Vޔ��nQ�I�p�j�|�Ҩ��T�=�z�� ��M�ԯP���Σ�Ź�1�/��Y�ںƇo ��+�[�U��@�v8$6#;.4>�۳.mX�@i���7��{�QF�6P��_t��)HP��ѻ�ʛp(�P��A25�M�C0�1��Y@Ӓ�'|$����m�o(��)F����4��/Z�X��H{@-�^S̏�ī�.QDp�D��]!�s��m|j�l�lghU,:I�"���|��Su�vf�;����]CQ��A5�����4�=�wl�.+8���ݛ�fu����8��Y��X���;Vd�ɼ<2ƧE���n^(��g��7/:e�X���a�<*�,���@=*�u�Kj�Wx�j�u�+WV�W�,ۡ�	q\�Q��pl�����j�yY+�IWsT�Lc�q��VE<��u�K3SR�+י����̇yQ��Mg蜰v�� �{�
��u&[��y�p�}�lٱ�@o�|cM�eYH5��7v'nT$t��vm�j� ����	�a�̱w
,7�.u�ڻN]���Y��K$�[1�1۱�3�����x��ız�*�*r˸���<p�h.�I�� �n�odŌ�w��%
/+��%�j�.�*Y��j91��kk�Ru�,�P���9;O-��DAw��.2��*�ҫY0��:��j�kڍ���y]�WK8U��RY���\������2>֨T5��0؈�tIf��,��]�2��͹$�W�"���N䠁�H��@����G!$�	�Ct��[���吂��)|6In���Y�O& ��u��7(ZԵ����.�ĊS�*�:Ս�3H��S���&武��$��6�ʻ�:�oxu>�Ŗ����}&�c�̧8�m�ڽ�Oi��ٕ4��"�1��=���w\�b���h:Xu�vf�Y�N�<&2��:U��F�c��H%�d��x�]��Wf�fw�q��F(�ٜ�m�Xc�B7H#)�媶����u �'A��5K
T�����(�Ø��\S�ڝX�G�t�ق�y�) �b��:�Z�D�R�n�kY�#,N����`�S�`;�f��x*�MP)��RƮ�F���ka����:.-�9����_s'�X����|�o��]�Y���@���u��{)�01iئ�I0�p���!�U��7o	��KJ7�Cz2�Ŷ�N�w[kQ�[mZ}LS��NbX�%�a�Ş�̃��lɝ�px��B���K���R:�ӇS�3�uX31�8���6И#��ۄi��H��y�A� =���x�r+n��s�wyE�+z�[�;�\.U���8���,unf���қ \��_��J�,���Q*��6e&벌���Q�3+&T��3�\fC����<��h���J*�n���%�ZZ������uu_����1���?9�Wע{�<?O���ϟ���Q�����9蚩
%�MrQN��4��1���oo�-m����R�q���8���vV�'�s�C�f)��Y���x���R�,Ƅ}1E9r�Ywҏ��M�*uܛ�1l��j�P3���GAƍhCxI.�^S���lF+:�|7�*��I66t5�,j�zd�ɽ4S�qV~ы��S���o0�Y�ł�in��9܋�N@j��a]�k�GMC>w5�\�F,k��H_u�%B�خ���}��fˆtX`M���p�S��W�4�@A��&�>����ژ�mu�K����W7�ik㕲�c]�+�3ʄ��N�l������}�1��{����{�,'D�fRh�P��f�а5E�c5�y��Lt9��U}��gZ�[���ω�[e����|�9��T�f�2�'4wU����N�Nf�5Mp����Zhp��S�r��eb��7y��J�����э��L�%2u5w٦�i�>��� �\F����Սf�y��e^���ۃ�9@,&�c�1A�"�rc���z���/m��"f�{,8����6�o�1!-���!��*t�bi�-�������NN�ajޭ�S�'K{ȗ���(�N�Y�'�j���(�/=���g���03���:�ue)֟<��ɻ	Wa�sx��>|�V.[|���՚�'��e`4M4>5b��E�N�����"��,�f�f�"�Ej�D���U�'*WY�4�r�)�nB*��,���:�"�\����Y$r*�Z�ˤ�����H�\r	5�F�6H�"�Nr��FT�ثuJ�HIUXL*�$���S��(���8\HUBQ\���&Aj	�W"鲮t�L�����I�]�(\�bBI�4s��fI�2�1�QG��ĒC*���jh��A �,ʩ�Q��RU��raq&��ۈq+J5���9^:� UpN
�I�H.�N]$�n$ȓ�ӤHn�U�NP��H��	L=ZyR��iE�8U\U���$T�S.�ӤD������(슩6BG9es3����!"��DYR�6D�F�T ��az�N!P4���u�!P��gNZ��Q�"ꉑs��IK,�r;(*�����x�ETD�C�F�(�2�B�G�� A��@p^l��*�w|9٢�`�m�NƠ��۲g�G�'lu���M�����nޝ��:�v�xʚ�X��G�sT�k�nL�R�ޗYd��^�[�ٿ���
�VV'��1}wv ńW��p{�1��$P�^��ю[#]O<F��.��1��/��v�OP)h.K֫��p�f��1	�[�f��0ԲV��X���^O�b���CL�!�2� �˩�=	[���[��70��63�k^E��gG����A�A�#0�R{N,3))�]�Ri�TnTt�h��xg�璴U��쉇w�,1m=��Lp͒FT��Y��}Os3��(����l�)D^��
D*���\oW�)��z���ײ�n���rϑ�;�o�Cb��<� _?�]#9�%@b������u���J�i��V��[��Zk�y�Q�lY�أ��b����3W���Z�OHtd��v���Y�����6ܱ�����S��KF�3Һ��^������+����Y;��bɫ���ۖ�F��:j�����_����
�x	Mb12�暡Gφ�+h� ��I��0-�Rܼx�BЗBk�����Nh�w^�����3��x����X�F��s,�:h�KAMn"D�*t��ʨ�6�q!��(N��{gJ#���mr���O�:o�y�$�WT}�v)i�w7�2�x�Y�#ic!��Y+)�3�-\(CS,m�����:Z8.!�Ǵ�r����~p��<�Q�nzs�����*�Z��-�3q5����}��O��h�p�W��{N3 ZN�C{\�Ӵ�B�7�㺁v=��������C67�i�u<8	
:�{(5O,(������)����YHN��c3��NӽoiQ��6��/<@l�)����1���	w\U����*��m̼���_��q����q���W��!I҇��.:�Q��s�s ���a�̻L����FBo[`wo>�)�RϞ���X���`<��A��J�ܐ��a�;ќ�C���WDl��sOY| ���0��na3���J��Щ�s楒�礅@MPjN���C�<�G��٭�N��
{,)5�C	���߹U���r�&�c[<�S�����q�紵%˻�^m^��;�v3�����Q]��0���f�.���/�S7�\ ĤLL!�����^���am�歛�q&s:~ǵ���~Ҳ������]��b(7�#c��^l�h*V�F�%����9�m<=Aꩁ��[���:F3�gZ=N�3J�A�d=����@m�ˋt'���ˑ�VI���&-�f��g`��χG�M̝ (��v�j��bݐӷ�]Kj҅�0jUK����6/G#�2��1e<�4�K�CGb0��iV��/�nuu�#��Au �_<ތu�CL��j"��[8j�,�k��y+e�tX*��Vr��FUYB���uBfosI�i�ޟ8^�lU�{د����6�X!���8���sʋ�<��"�v���a����6���[=�/�����Y�kL�V+�����q�/�4�HwCVWh�j���Z7�:;fbGE�l�Ḗ�gŇƧ��ʖ|��$8A� �<�Z8�';�Y����5� :��å�[�X�i�tux`�z'���r��B��^b����$��r�ÇL;\�gd_ꎹ�H*|�2�q7y����ۏ�|�p���^1�H�PB�s9;t]��$v����� �ȯOO��*��n�$Tq�h֫���m�0h��{�Ds/A��-]��B����F؂��v��V��Sj��z%�|�)���VҒ�f4G
��+#ѐt|�h�j�o�zJ�V�>4�����urW�CC9=�-�ct��:�}>�/�T􀫺��z�%	-��G}�f�k3k�f�>�v� 1z�南8��A
4�\�N�2���`�/s]Ku�gWu-��8�唦R���th��/��n�;�9��A�/�䘪Wg<6�4D=�n�_1:�41ZYj6,0�"���Ue���R��<{����d����X��4��B��1'V�yy��|+���@}zVKܬX\���>��|����n���Ug�9��Ƅ��Ȅ*T�X���7�|sF�P'La(n_�lr7����#eH����y�ѩ�w1;w�N�v�s��8c�T8
;��V����0�\L�,7&�>��ٿ��W���u6��i>��Z��?W�7QD�r�������$��p�r��ɨ
vX�#��<Tt��5��L����7��N!g��>��E��wV�s�V�PT�v������K��K;1�R�:L����h�r-U#7:��z{������F\U=p�N(M͌xϏu��Kh��=�"�*��Tz*�qɖ!\l�B6��o��seӤ̃L���E>]j~T{�!u
Sqn���3�A��e߲�.65~�#Yxf�:.$��!�Zs6��!*��8��4E׳��{��̇Ҋ�7g�UN�@�)� �D�K��x�Ő�%�g�&��1�kt8U�ɦ��'sQJ��l꧌7{����í{ ���b����ܠ�k����9�G&�Ԕ]�ۨ��\s���>#Vnt�dI�-�hA�2����jc*���I�&�˃�����5:�2����8rs���*L�|a��>҄Ii��ڔV�p@ɭ����B�oº_T��^���y�"�sk�Q�XU
xh��'i�h*L��D`�r�+��2�:+�%�>[��T��r�����ω�^*C��d�'��:����\������	�rB�e�t�T!������؛�|$H�WH�4v���	M8�j�p_>�P��7XȒ��t�lH��GmLSY��h�;�8	�r�&b��&&)um�0��	�#���}V�.NË7�S��sS^X�FL`UV����
׆ۢ��[#\��^��ew*�~����+S����~y �y�͛��f��U�/��L�r�Z�`Pc����Y�d��y��ɚ� �祮�(̸nt+��3��0���:o���@yG�Y���1G%>���j��S�]S��L�ۭS:�n+��o!��]m�l�=�Cʜ0�p��W���f��8�R������g����,+/��y�1��|@}��P���J��yA��"ܯ0\���������U��9��\a��#�`e]�N�vkn�|�:�v���R�jwg���C��K���YWq����4a]1rᚮ��-���M</�Bs$jE8u�{u��y�nq+�<\˵�5Y��bU���}a�z��%��X�ǉ�E���V�dpǱI���@���s��ϰ�:V�<)��d��P�{���.&q�v�U;�M_l�w�8��a���ô)ș��f��u�)>p����P�0.j��Txx���-�EN��ss؋����ξ�5�R����cZv뵀���4��鞕���L=.#\�;EwvjY1�yR�;���e�����p�#-��^F��N�Ġ:��$�&�0W_J�\�ސ���Ṵ�w�-;�2�����~��8x�;7[��u��n�u9������Shy�U�Ip�ˬ|)}��i����=�q��1I��c#	q��]�����y�q��p�=3�xCwT�� ��� (�^�<��c|�#�>T���
��M��cU���$ ��"�S�Dq�̊SQ@��Þ%����t��ɔ�O{��2�)���u�J���S��_5$L#!I(!`����S�rg0��S���Ɏrfc���yZV,�K��_S]PŹ�E��[@l�޸~�Diu�U�n|��N�y�`���rV��RΔ���&5A�.��"A�ޏ��lz�5M����ׯ���:��8E�������9P�c�%.Y��V����T%��c7t,<n�ڑ>��ׇ��DGz��[���o[g�}󖎞j%�*rR�S&��r��)gi9�4���܀�/�?��ؐj�Ƈr�9�	�lQ>�)Ϡ�(m�IS71i�ύ�ҭ��;�&��^B��z�.�R���^�����eoE'Q���ɠ�&;eqʬ�,9
b�T	����v�Ԃ#�o�c��g���{��6ǿx�Eq�'��A���@	���2QXU�:̡��=Ty'x�D��kԺ$�.k� j����e+�;��{�w>CxX1OJ]�����8�������/�@��������'�Y��p�o%C��q��KôK!1_O�ǋ�w��=�F2����95b���ݢ2�U+Vh�󨝞�j�p]#^�uP7\�oT�i��eW�p���#Uf������J�ÆÖ���- ���q��jp��Qs9��&v�v�By�/>u����,߄Z#(>W<|��p�]\�|&jrlM�3�����M�SY�	Ƹv��}+:h�8�c^�|b�9cF��{���q�9.�r�Tm�F�ꎹ�@YB|�Kt���q{�k�)����8�ulȪE�A��<y�dM�>�u{�v�n#;c�o��E��V�T��iW\�Ŏ��s�fr�2����n8�v-�۷J��p�y[u���(�]��Zڏk2�3J�v7��t�N���9��ƨ�7lυ�����]F���{s��1mN��(HЬG\k�4TsyqQ~Y4�� �s^%D2*z}>�ʃB�۲4T̩�iz��][�w�V^O���q�!�_C�8*_]����� �JĀ��pu=q?L���C�M��Qc$�=���+��:[7f4Gnm�+ȋ�[����
��
��,�m#��/���f�eOa��b\��0��3r�g~f#���4�i�D�Qo/s/�X�3fv�^�w�yG�:�	�T�]!Q�X���Hj2>��:�r�N}&0a����&u��ݼ���_h�R[�'�:�[�??��"�
��,RVi����>qˑaa���k�d�}���A��x#����˅A�2�1¼�|o�h�5�	���{���PK_������iʨ�.#f��]�����~�M���>F�#��8��0;�Mh��c�9�'�E�ˉn�*Ҹy�3��sˤB5�X�Ϯs�t��^��Vu�U�Ncuظ�k�L7�}�]8嗊F��t�:�U�_[�GAϓ��5�����t�D�����"��Jo����6���#����Z�f���rDT9��N����\x^�e+��+����f���p�8n�s �з�_>7�wH9gu�|M��ˁ���\�5sc%��vt`lx+t��)Fs8��VR�F �}K2��@��j�xz��/��e����N��-ʶ"��|.k�ԋky���nH�S!�B����8O@hl�Dm��o�F�P�����a�qcf�6:C����������m�m7�#r��EgPw�a2�eP\mSW��-������zۄ�6��㓢�v}��@�J[ۡ�
 ͞���0�P�VD�Χ�p��}�U���\X�.3y�<��6r�C���B(�v��OQE^��; v[hYU��y��R#�@;W2{��AÝ�/�XW���I�F1��3��}=�=%� �bԙշs���G��z�΋0	��^'t�9��:.�OB����S��x�Z�qw�b"�l0'_Տ�'��*�/� �;r$.�]2D����Į1��q��ݶX�SB+�P�w�D����.�A��l�{=wD1��X�-�L�=5}$
j���H�ݴv��jw�]��>�u۝Ҽˏʑ�Í��#�L`��>X�D
0�e��+E��x1�{Fg^�G����cƙ0�re�}d��0dʷݳp*NS�Bv揅��M�9����J����pq�����4{��9�Ɯ֭]s3,k��Ц�p�Znr�E�jKQ�*��BP�x��˖�+��)7c�}L ���o6��Pq|�Lw�DPʺ���t�5//�Q�ʋ�~��3+6{����T�\#d�-K%nA�#E|(1�y_*�����ݽ���n�)�9��-Jf_By��3�j(���D�p�Ä�H\b���2��R�����N�g>�����j�^�.ׄ�8�J�F.���g�뢍�Za:�lXh� <�����������EA=J�p�p���|��gظt> :ݷ�v0.?I罓k}�|�1����/���s��1+ �n�o(�!U��6B��^s�J�q-qy�U�����w�	W�)]�Ѱ��%&Ŝ�����"�c6F�G[f� U�)=���.iH|��sHq�c�݅׹p�3�^�����cA��|�^���,E*Y==�7��1��˴摁�ƣiU�����'-��ۘ�P�jAgVu�lJ������UdA'u�_]����l��dU�"��x;v�|�l�Ȁ�����N�2�h���MK���bL��ׇXkzE����uD�p��+��N�}[�|��9D�wH�����Z�ݮ���3��̎T��o�̱/�t�������Q�+�S�`1C�z�JF�)�j�!ɳMv�li�,���u�5{8�X�I8��X���ie���!�'lw�S�b��r����c�ҝ�RJ�o�/YN����1a�3Q��;���Ǝ��n�J|���6�p��<��Y��4�u΄�1T����2�+:���,_9MV�#�ڹ;�gCi��|���fpjvq�4����3���Vi4y��l�0�c(&8��\�igGQ�p���.U
��]�+��$�S�(�b�uJ�m�heֽ�[��.l�N����|:��޼�k�7�\3�i�q�m;!��)��J�	�|x�433���jA�R����ʜj|U�+; �����MV�Ų�����2����K����yIڼ����ҵɚG�-���U�:��S�zn}׎9әūL�եJ���\7�t�FZ�d�{��I�N #�l��\��67iv��3l殈]
�n\.3��K{���=5��ս�l�vx7�����}4v1�j�0vLo�Är��ݙz�����<ŝIƺ�T�vQ�*W»�Еrb�s@Rּ�z��68���P��%,��S6�������Рށ����u�x�3N�n���z�ֈ�JO%wH�}� �ݔ�׹���u�VPws�UA��"S�>5��\�����^�[�:��r���q)8���ق���q�F�S1q/[�&Z,��ۧ�{���M&��n�;��hD���(֠�jU��}f5���j����ea��P��$��.�>���G���Y}�ˣW�i���ڷC;�(�:"H���T����R�V;C.mp�a)�m��RF�vɗMn�a�OBE�}Zz�Y�V�:ȴ#wfgӠ���Z�=<Y"Ԫ�����f���+��h05*��it]u9��
���W�m���,������:�m��E�8Nѕ�Q����:os�D���Ҵ&3k:R���1�a�������̕���J��S��Rj [϶��;F��(Ў�]<l3+x+C�s�1J���(�Vź"�d���H�9�ո`�\A���Dc�v�Yz��3'u�enϟt�3V�+n�*є)�Ս���(*D�PƼb'a�q2�g^�6�5k�T�[��ƕ�;Sc�gG]�����fYN��g^>� ��3�e�`������ظz����aBr{����=� ���9i�ǉ:��"�N�-=��Vvv%eJ�莣"cE����aڊ���������\�l��k:���:K�7:��18m�A�2�M줪u�5�J��u.��]4͍�֛���@̫}�;p�aQ������]u�|��Vߕ*���k����k��M27��ܭ�t��}�V�cn8��/8�k�SUw�e}�:������f�N8�xSZ��V�ڇS�0�81���J7IdS6�d�eǉZ�(ܖ�
=�=��4S�j���;�ȝFoD�t aɂ��E�ʢ1B��T&�g9\"��(ÖEʉ�&s4:��l̹QVg��[.G!#C B�)$�Ў*+XgNvU*V�%�3����i��E-;��"E�±b�*$+9aE�S	*L+�+$LP�����$.PT��꺈�x$-Z�ˎ��
" ��*T�T�I\�+Z*'B�!(:"�J
I8^D(�R'(����r����Q�PaJ�(�NQ�T�QRfuӋ
��aTQ�%9)Ur�!f��b�UQ&��UEB`�h�����*9�r ����4$�,ۦTEPx���Av�"
��#�U2��Qʩ%�B�M9G"
��+6jQ�Q8�(.U�\������������
�(�1*qӹp�"���L�ZQh�иr#�Qʪ�"��"(�%i˝2 �QUF��r��\�i�$�*"��Ȯ��Qx�(!R�H5)�R�\	\��"* �x��K"��H4hP�L �V��dz!���=D��1t�r���N%EJ�p�1F��9���喟sQV�k��dy�sJ�YO\V�3ȋ�ݥ1����:��#������~�ߞ;�©�["o�� ��d<O�qۿ8�8�^�G�z�i�P�iP��OP�����0�c��}��w��I'�y��݆!����ɜ�_zchV��N�BP}Hx����sI��;���}~pvvy�}cק�aw���Đ��T���!W���8���t�������ۏ]�8���8���C�?��	�@ G�(D�D����?f�}�UM�h�l�{ (@�� *"��(P=�o9|N�}BN?ɽ}��ߐ�;J��{�;M�'�s��>u`��?[�;H�]��!{o���%p.:|C���]�㷝�]�$��/�ߞu��߾�����><M�~N>�κ�;������7���®=O��oP��y�]���8�oN8���m�;v�;���>tn�HN݇���+���7�ˤ������>_�@�$]�޾��G�λ�+��:����ϟu������;I�}9e<v����7�?\~C��}?s�t������8�]��~yÿcq����޺���;��u�6������9���8�q�߾s�z�!���8�u������:~��=�W)z��DBAb=F,A�a!�}wJ���p<M?�ӷ�����!�����7�O��9��t�������q���aw��ۤ��w7~{��a�\
n��}����;�W���,�k�ݽ��|B�w�4��8���>Q���?;�'ο��M�v|�C�}C����}��{�m�?��8��	8���e7�N'A��]>�I�BO���ݿT��*����@�doz��d�l���q I>;{���л�i7H]�}�n;�p.����r��~8�C��&���p�0���^?\{��
���>�I��&��|q�C�����ĝ�I��.y�痝��]���?}�|M���������&�F��y�7���<v�c��7>��y�]m�;��Ǵ8�v��]��&�	���8�탈x�~'�}���;��7�t�T�GP���ɖ���9���~�N��p"o�q�?{�>�,����z<C�q����9�|w�8��;���
��ĝ��΃��9�ޱ�w�iۿ<���&���v�޸o�t���);�[q7�'z������|���}�U�%rݭ�ɗ!qU��we�њ�j��@��7C��S��;!��jl�s��In3�u}t*�[ŵn���3
p�Х�����Ap�j��S����)]3�xQ�!�w(XnS1`�I޸;L�8�DU���-/xvq�Y������_���G]@z���_����v�w��[�:L)�����ۏ\O?}�hx����7����:��!��C�����0�~��~C���_H.��7�ݝ�߽��~y�ߟ=�:�u���~����~@�4�O��
������v8��n�\M����>��o�~G�oɷ���1��;뾝�͏���
=�dA���f�W���61<����zwN����e:M�	2���8���};�h��;�[�����$��X��!�k�7۴;L/�����p��<M��x~��oY�]�v{��DECQ7!��N�>�j����U�NWp=�����X�#���7��[w�t�]���
t�׷q4��D����Ԧ���G����'��7�ޡ�#?��aq���ߝ��#�©,��:v'"���NQ�.w����wi��֓�&�����?p���H&�Ǟ���i�Bw�~�����q�A�N<|z@�w�i$<w�uc�:L(uG��q����1�!>��3C}��1zD������~~�ߩ�ݡӸ��߸��0��whx�!�o=���>&��{��t��w�ߝx��7hN����c����Rq8�<�q��)���O�Z?E�|D}P����6�MG�7�y~�������8=
S~B�m��~}�q\x�ǟxx�'�����θ<M�q��޹��I�!'��q���������8���z���=��i�ỳ�
����*���2������{�L/��?�u�M�N�p�o�]��c�:O��^;����M���g�p�>>8'~M���v�����0�K�]��yקt�H
)�?���[�`	vm����2��r�+�穪��";N�㾸�q=:��w�8��Ǵ:L.?���u�n!�����t��4���1�v����~O��o���~u��1&�	�<����pq�Oz�>��G�#����^���sa�-��;I!�����SHI�������v���F�P��q��:�'i��!��7�����
v|��C�:C�;>�����!ߟ�|@�$�� �1bG�P��"�Ƕ�;1���]Jȯ��I�kZ�|�d�}5F���F��8Lh��;��{n����8�J9x����g��Osx��X��w77vaջ�<y�B)d�����.�o��/��/�@�qp��h�KZռ��HY��.�Q�#�^�۾��D�!�@�����Aۉ���m�yÈt�@�'��|ۤ];Hu���C�[;��BM����}9t�pH~q���������aw��������ߝ+��G�"y��n�|���ͱ�y�6��7ޘ_�?��zy���돈$��Ӻw���M'�!v�һ�k�~tn��0����1'H|M&��S��~g|q��oP��Ǐ+��'�|�����AFo�"]���q[����D���:pz\w�k�o�N�>p���t|�÷�|L/����ç�?��8�q9�{ю�;�8���:�:L*�~{��v�!� |=�\��8�}M"< ��#�0E�Y�G�;����T�3y�׻~M������wN7�>];�������<v��}zC���7N��I����t|Tޡ*���7��8������>��qǿ�s~N��@�U�� L Ls�7�q׳�c{?�~���?|��I�H'�w�[s�i�_�XP<I7���N���M���8�_P'w��!Ӊ����������?�������EӴ�|������+��|�M����{�����~~~>?:�j�[`�w=��!�A}�U�>�
|���i�o<��8�Wn�M���L>@z��0~{q�w{�t�}|M�>�!ӷ���!�����C����y��g��}���w|y��^�����u}��~~�^aO�\x�����&�������W����zۉ��������F흻�:v�v�yǤ��aW'�P>�������d?'�q��h�� ��"%=��͈u=Q֖����]|���{�^����G�8�!�&������8��{ z�ɧ�^}����7�H^}�q:W����ރ�q�������N�~���pw��I�q�Tޡ*o//�������������=�������}N8�ǧ?�v������w�7����E=w�<C��p���S���ތt�Ă�~|��� z�o�?�'��M�|��ӧi_'�X��N'��u���y��
&{�ܬW�s߇� P<`{�I
G��.�v~�M���ǎ8�����B�g�s~t�8$:w{�8z�M�x�L?}�&��7����p	]�����<C������Hz��$s�zs�ޮ����R�HV�hR��d��.��&J��R7}[�M���N�
���0�_T)3M��'���� W�rur�*��7и�]��)�� t��:$hl��5���X�ӬT1�붅�[b7���`ָЬU��2D^�1(ԥ���l��[����u�ߟ?{����&���(q��w��:���ݡ�	'��۟�����-�N�v����}��oP���y��{��;�<��v�8�����7���:qg���|t��*�O�JdO��O����?{�®�?���;����e����㾧�YN��;��>Gi�C����Ğ��:v�����A�C���;|O���'����Gׄ�� ��<�w��F�s��;��x���k����s|C�4�ǏϾ���aw�~s��W~v��X�o�q��|:�L�����g�c�I�aw]������N������S�
f,G�A v���TL�<��G�߯���7��w���޷�|O���L��8�q+�����7�I O����{��	4�� �:x�"��e7�_��'g.�����>'��r1 p�>����L{�w>��no:�p���{������㾦��n�����ю���'w��C���q�����O�>{�H�9���D[6	>GĬ�,F��A�Œ�ћ1K�d����mj���	�nӄfm��>��X�"8���N����U׹�.�h�6�$�ɚ&�y��~��d�F�3���
X�'#��CV�P3˦����j�/��M�vM�4�7c�T�Ce�B�e�����<�S�tZ(?>����P�7Kv�-.-�}�Ks��+#|��b>��m����O<��;+�1�^��Ԣ�v��~�G\᭠=r��
����}���u�l�ˤ�Y�>gG�+��F3P#��3ٴ�4�F[�}�5b$cf���l���ַ$4̂h��u��e�u5��E}'5˱@�L}WYn��^'RК�z�����j��x���kS2n�wJ^&�L]N��,�F.�A�Vm˾���xy�:3'fm^:�����Bۧ���g�Q��2������Y"��e�YQ��]Le�2վ;��l��J.#^����
���U 3Mll������=�Ύ櫲-F���m*���Pxo�岑�
w/��G���/h��"v��4�t��,��=�`G9�j^�gCD�Jw�KGD��XXOr��n��6{(�Ϋ�:V�3֚I��}�b�̀T�nF��p�\;�ً�mt������O�	�:ދm�וNj��w��9P{��`+zo�#͙'D7~�TE���5��[�޷ZVq�(�܎Oy���lT���9u E�}R8AF�'Nn �f��ٟ
SQ@��p[;��E��U8�6�����<�5na3_9��{!��U��0�P��>;J�8��2R�5��{��kh�Q�9��&+�����3��9������*[��ʤ���
�-R���N��ݺ�C�rC�~�YLo�w�*��J\��3�f�M�wn����nzX���w������3���R�۷V9�ሺ,?v�)�,t!LRj�18v%���ᾚ������<P�3+���F;ʝ>��}�K��7aỻ�ޖ��W�"1k����wO^��֡��a$W%h�@���;#�\�|�^�6/��z� ����R����������=�]�f���M�Eeig{��hQ9����x{�kx�n)�v��c��~�|�1iȱ���Wf�Z�ay倪��@	�����7��e*SU�7�0;#�x����B���}�2%�rP����r�W�'"��;3��1R����3hVp�f��q��C�s�X�(w�m{��5	�e+\.[�[�=�9�H�Ŝ�v��M&�U�r�h����X�g�v_�W��X����Ύ�k+ӯ(��f�w똗�2ד�گZ�g�2gzb��!��_e��l�6W3Jv��{SŎ3CV�+t�,>��+0�E���QV�M��K϶���^:l��hڹa�B{��f���̾{6����T���NPu��gנ��@�:��%5�@O*�֕o��>���:�]���{ǵ��%����dn��Z��l��1�(�T��2�"o�W��(���=�����H�¦����p�ܔ7�by�GnOM�DP��H�ʃB�ԣ��y��|���"�;��xk9P�E�>�9�H�&��bp<�T5:���#F
	=�����p����+�]L̡����8U�[��_d�(j#���۽�N�.c@�i�@�{��'q�Z�cR�,�w�c��W"�M���r����y����Q���5$C�4�:��D֌��P���:2�ȯ��#�5��Q댗^���=v��<�';���ru�p,7y=Ƽ�`Ξ�|ꂇ�=u^���F��*g]Ԉ׵�lap��ƽݮ�CE�F.��dR��"�J�e��ê������͉�z�x�f����B�c� �!����VG�!�b�7szm�"��N����gf训��ݝކ��R������Bbx���Q�m����v�
��~CGoهT��u�A�fΠ��"8SJ����Ǆ��f�U��D�˅A�2�6�f��8�L���m}�q�7��Z��n����q�s%�Q�!
o.���ٕ^�Z#��6̤k�I���WS�_��l��{J~>�m��=LK阠�g��<��N�r�{?'s6q�$�^�oO��VU��n�'�w%�g�W�K�y4!��6s�s�Pڮ���Xʃ���Mؠ^�y����S�.�
0�܁�nK�q0��E�aC	�3������J�|(S���o1��f���0���7x����K/�bj��{��juIWx���2�/
�5���W�k̳<���ko�t�cU$=��ً�ɖ���`%znя/-ۭ�N�'yj3c2����yLVoXU5�������u��k@�͘��XE����wHv6�<�*�gm�e�RO�[�R�d�ݔD��4���nm�e�����eU뻂�����{�w=�3YV��unRvGZ��'����a��ܧ��Eg�t���y:��G��u�K�)f_A��_TE�zy�����u��"*�̇Ҋ�7��+6.(^��wv��HlH��D���>�y���i���qv���v�"��2 $�w4%�;���@�ݒ�C�V�i�T�;: T9a�P�T�	�N�1�㥳c`�}P�y��j+{�]H+�k��̣�0#`.�U�W���v2zy�K#x�}��e�����k	��#�s�U�>�麬�=$+#��E�$M��d�F_���JO	�}d���n���T���n�n��CO�H_[̂"˘b4��nd�������:7J�=�j5�S��iK�;���dTĈq�´\5�l��]+�X}����4(:5��+���l�:�Jfi<������\���uG<��L�j}�N�;�xD���I2�eN�����T�p^�'bwJ�g>�0����B����&M��_�fg�ˤC"���=�T8uɳ�Nt��i̛�w�+q��(+G:���m��m�U��I���uM�c���-*�i��gi������JY��Q�6�)��	5�٠�!UV�́�����j�մ��8F(�)X'⥵��Vq�y�Պ��<C'�p�ʂ���191��\O~��S���FU5� 
D�������B+�R����B��B5�:vy9��_>��������|�c�"��{��0.��T��P�
�a��@W�� ·��8q��n��97xyǕW� 8��l���k�a��w�X<��[��++���gÀ���h��-0�2���o��Y7�q��8#�Y|���Z����h<5�_���חF/�G^d��H|�c���K�J����;|u�c�|����Cƽ����Q�$p;ynJQ<bQ�r
�{�N����
�&Q�0G3�m*���Pxm'E���9�* w�M\K/�.�aViYۮ�W*j�
��V��%�/��!ŃEBt{=�O��GC#�i�N_��N��y���))��z��e�#qĺ#��T�S0�Vy���hE��ƴ��-�j{6�̓���P��܏7� m�wq�k�h�%�neI⺞�!G]���Dq8��-1S,nu�N󜡑1��T��o�-쑢��d'.j@!�ڃ�zP�Q�~��[R~�򢱾�NԬ��RN��4��-�]m��1�	9}���ܴ��j`��y뭭�\ns�d*�UF���W ���D�9����4"�k��I�g� ;4�*����j�zK#W����NIJ�4󫫰 uo$ڐ��oz��dZ���ꪯ����������4����
ɑ�k�<n�ޚ �Sѐ��"V��E?�.;1§�q�!m�Zzk�K]�=ے���a�C�P��7�Ź�E�ȉ[@u�y`W�.�GoK�Em^u�M�8����x.m
�}�ؼ�9��Te}�[90��J��!��#9��UJ:㯞��̓޵:JӂHQ�&�5yQ�T\��k��&#�PiMIc���f�k&9����>����+�ߙ��#��H�7��uٮ���s�Y�� m�e�+�&�'�n��(ghA�*��_�E�\A���׫�I�d�8rG>^���X�Z��l*��1]�s|;�ò�0ŚD
���1�#����i�������:b�%��s��'�Gm��K(]��ԯ�X7�u�v �ts�s��(�߽�;��3k|r������̍�����g3�b�����}�i�_
ߤ�����,�aY���u��Qh�r��
�R��rf�K�`�*���P���U���D�������0�l�X�u�����g4խ��z������:v��u>c-��L4Epq6�s��?�U�l,hV����2'O�ѣ����4�jJy������g3��ѭR��H>��.���X��%tO�𒻝�n��i�T2���/B�G!�#��!�ZF�$���`�x��a>в���;��!��6&�n��gj����	��Dd��������y%e��WL�&��ΈV���m��Bf�q���S�VEbn�H!�ɻQbpL]*���1���}ڪ6e�B��[�fl�W6V�������':
�;-qw�^�FJ�-T���L���ݥP�t�
*��d̵o:q�J�P�ᛜB���l�B�����*'5}�`�n�֩n���	�h�ޫ�d�7U
�tB�n�4���I�+�ʶ��%E(
�;��ɕ�Yh�8�]��L�D�!�*���<.��¬Rﻍ#�{t�{N��-���J �!;ā�ѠaƏQ��F�2,,��IT|]�k/f����Ӕ{:�5�E����=ťyǲm��܋��Z�{��!x�f3R[ך�ڛ��Tet}��k�K��@3�+Z��{��ZyU��s�Y׬�̰]��������(\�Դ��U�X3�;x�ܓk���z�r�8�B$�&S,�I��t^��صt|(Z��ww�7YO��X�g熮�l�����Ƥ���ة �\��G���52��������ˢ�����E�
m����	�u��|����[��S59ܰ5$�џN�}�y�e� iG���%�j����	��m^_ٰLVC��j�U����,+��Ý�N���Ұ��oTڎIu�Af���^ɕ���0���
Pn��St��*��Z�y!SWrF� ؋8�@k� &1p/j��u���J���<.;�,�tkE=�	��V��5֮��FVQ�ՈN�x��а�u-�V����6�'�U�����9��ʮ�aZ�c��f���-=���^��E��Ҿ��[-������d��q�vY\����m�௕tt�e��]:\��n���t�n��:N�#�E@�f��yG�������Y#n����0f����P�Q���������`����5w$�ۓ�:;��n<<�5�@.���n*���X��l)�u�l�4�=���mY�G��v�+��0\C1s�s'P}�V�i�j!6B�m�zj��((殾�n�֝��ѵ���ЈR�U�[Ĵ�i��
�m.����:v�V��u|���3��D��3u
p��A�P��'�;2��N���ʄ#o3��YQ��ƫU�a�=�h�� 󂲥�*ۻ��"�*T��5_w����j����5ɱZ���΃]���՝d�q�����=X���[��d��m��p���Nފ���h��"a��\�O�++x�MZ�<�7��Q�Ҳoaak�������Q��Cd�N���Y����˳�v��AP  �jh��DZ!2��A�_��!]��y�WDEU�]p��r���(�EJ�
畐�9TQ��d��r�r��*�W��XH\�i+TD�S*�B
"
�����YPZ�t顉$��L�
�E�I�&�,+�US�y�8�֗"�`a%GU���V�����qBN<^\xrYP�x�L�5�&a�:zQTWD����q�Y�������8�����*%hT�^��<K:�Ȃ��(�sȆJ�8
��"���q�ȎȻ*�t������s�c��9QUV��DS.UȏV��^��r�EU̠��"9ʥ4"� �h�AI�%�"�u�Ar�r.U\(�A'U3��7QPB��Y�QȊ��AP9U˄�g�u@��Uz��Ea���ˮ�{���u�z Ζv�Z�NJ�:|������
xű��oJB������r���CWҲ���H����x{�7h�O\ot��LV��{s���5�hSө.5�@sʻ���}1>҃�kTnX���c�)iL�^3�{�6|-���W���Q5[n��@����~Bxs�����!6��]���٩\<��B��(v��#E'uU�QEߠ�s@��d>Y�ib���.�^,isB̂���q��_t�JS��d��\���F�uQ#�>D�\�{f�%%2�8s��n��"bK�d\����)���\U���dƈ��z��\N1X�K�=���{�gE���ӵ��D��Q��#�"��XBD8��0�t�s亙��/��S@p����Z�=����+�2�q�J?���i��A.�0厵+���[�����d� &7���fwY}*�S�&0A���LWO��(�[�??�yb.�
�V�
��慛9u��ّT>��r��ٱ {�4�'�\���y������_M)�cE�h�sY��i
�YA���1��@�"�Cn�@YG�!d�l>�Ӏ�);�=5
����;��g�Mǳ����"�Ǒ�x՗�d���=,�%�7�^�Jr���GVГT���bhq|̴�>��oD��jwL����<�ǉ.�euca��|,`�ӎ�м�ˑ�be>o��R9c��xcX�Jrr�K���{�B΄�+�R�m,z��1���ћ�^^>��d�E��� �mΞ�w)��$�i��G<:��k�-������������鱊\B���@�}6�����*����!���Z�լW � ��þ��/e*��;<'֕x<�`gj#׷���Ǟ0��n �w/vOn�	K�\�X��vۇ�:,�nf䋁����*.��b�Vg�����\�[��+X��g�q��q��S��[���t�\J���ziBjb\�&�3�w�<O���1Z0g;!:/��dTݮ��ޛ���y^y��e:c��KVX�o��v9UD�7�/�eh}��j����ļ��J��-���'�>	�g�C��=� :tƞڔR�E�/�]�ue��e0����$ɒ7>�H@��Ph�;���5�<l��<�`�	�V��ծ��6��{J�m3��P�#_:!�l�ea��t]�'�Px��NF�Q�S/����d�6�qt8���Zb5�ʸC�rB� �vĉ�Y"cc��KDe�e�H.���-���G[�i�aU�g/^+)��[�U�s���[u����y�]�v�{�j�<[��l�ԼyP�(7]�F�� ��M��x�YI���t�׏�f��W����lN������; !lcn���S�˝}M6�ub�p�.�o� �����y�=�Գ�Ǯ
�{V�� �=�D:yV�:s.�������b�֛|P�Z�5�%���.Y+��b&b������.���S ��Ŗ����>�}U�ֹ�_V���ǩc)�mc�5�"U �
�F ^{]TW�U��R��T���q:���m�����o���S�ѿ^۾+>l��u����I���/�F/�cq'��p��PΆr����mK����f��E�ó�Y�"21Kjp &;��1��n8Bs21�M�5��r7��Ø��1T0����nE����++D�n�:��xU�� +Φ>#T3�)g{���j�WMi)�����2#��{���eؕ���I��[�Pخ�Xɱ�;\�7��E��h�[�Jz�.�E�5L�b����T5u�FF�5�|�(��6C�U�_�����8-���w9�s#��,Bf��A��̨�B��O(h��yS����/ �u�r���uB��Qps�T�'����Y�B�^�ua@A��N[<%����f0 ��!��r�3y��v�.����ܵ�n(�*}�uL��Z��E����O��=�`�eK-����C�16�dW,C.��T�nm�㜩�E�)�����E��%m�uI����GXy��p
8����v�#R��Ks��n�򧿼< �o8`���`᷒bt���#	`]N�r���T���w��q��ڛ��[v�ګ��̿k�,��m��±�S�G6����C����N�l�
�h��y˖eַy�v�{�yn�q� �N�C{\߬G�2	��R�!t�:HQ�:�A���]��3y*�O��!	�$q�@�g���p��T����Bi׏U�q�)����'��T>�&�E5U�nt�n�n��
H�S����������R3�N	�|q�%Oa�	�xi���\�tc��jM� uC/,�����*r�\���e#Q����1��F;ӎs�瑗e��u��_�O�ze���WYP3�kWװ+�K�(����4MPk$\:=%.4�CK�������A�*���6�%186a�%bL_��^�����D�6$�v�k�B�0�~̯1�O��d��aU�!P�)��̦.( �g�j��,��ڈn����_ν�2|����c��/���D[<�Օ�:���Տ[GD���fW8�F�NwCMD�x�דF�A�l%}�����������Ž��wMJ�5���m,����|3�[&�r�a(U�x �נG1���˵�}j\;Qs�-�o��렱aga}
��gI�'*����������s�h�Ʈ}�~��pso�Qa'Q�uN�zds80u� B�������Y��Q��=ۘ�s��j]�d�scHƵ�����E��������Պ�y
w��g^Ӥ�G���y1��ry�<�X!����U��V�yT�94�y�v�;`���* X�{/��s+�(�]�qJ��-ڔm�	��n*�s!�1p+3�rɵ���{��)�\$�l���]bfu���l؉�#eO!�$8�i�m�
�� O��*�;���h�JpO�����߾%�>�7�R��:P�6\���	a�b[�O^ե��Y��l�1Yڹ����8�M���	�!p�J���#E'u��Wz74J�dL��i��L�4�R�Ğ�h�)��ٯE�>g�"�}$V���|�w��:q�{�̧eh���t6�#4�Eة
���@C����f�����Ɍ�[��N8%=�	�Rp���B��c�q��w�P
2�"But��r:2,��"�!�S}n6��O*�����c�.�[5�mpt{��K�Vᩍ*��փ����� �7�?ާMw3�X�0�߫�W3YؚZ�#y?�1��c�Z�V^MW��yr�����y�k�ue��,������]L�A�\u<��#Q�b��+4ʼ�3CWX�s2B����=t����|[;�&��o����O��$w����M'�������i��[�,���VKb����6,E�5%���@<��昮�\���孏��K��ȵ�ՁJ��"U`{̩�-�Ѣ��f����T&��UP�`Q�2x�m��f�⧟�fN����r��m:�:�6f+*6���6�2-�1*��
����L1�Cˎ�.E�o�>Ӌ�`�/;:^��X��=~��
�f�ו{ٯ���C���S���/g��]��ȷ���֬�$���,��!B�"�vF)�Bb�b*�V3���n�730�݇�*l̶}���͓�=�a�G¯e*�N�	iW��@_L�Ƕ�_]΀���eOQ�{�G&
շ��j��F��<�\�.3 �o�E����|jQB�g���mY1ݜҝ��1b;#�[�j�c.���+��'G.�*H��v&��S�ո7Y�{.\0��с�n��a��*�eKU��a��H�dS�8\Jδɑ���˪ś�!���'=��v�-k��-�.��Vt�n��g�{��{�=�5]���!��}A��38R�][�Z������`ǒ���v��KT�J�QO�.���5�
N�3��r��ZB��/�=Ko�㛜$iZr�mdKp�7�Q&6H��� =��S�<��l��F)����
YL�:�a���s홄;N2�Iwo�ϻ8��Rל���d��*�*�U!�Ph��aC��<4MBN�1�I�=l�`a�K̦�p����;)�C�T^�Th��a���xz��I�ؾ���j�M��*'�Z.t��.�5 :.H�gnD��.�"E�@��R��egN�=Z�эx$�����(VoW*��@�u�.Ǚ
6�P(�˙�zo������������.�i^UQ|c���ٸb-1:*!��e F�*� +�n����@�0�vbyS`ED�����No�}�^�}�nɨ�+K�p�Ɗ���Z��6��9K��gh��՗{�}�3:��$K���0ǆ����7��):�\'��1�(��ETeʞu.�Xޑky嬸��N���jK�����«�"��f���wO7�� ��������I�K���kM��E����g�֋+u�a�,+.�.�֙��c`/r����ɕ��d������S������kwP�Օ��:�7*h�,�����w��5����mlU�uh�� 2��dV)��5�e�CW7|+]�0��{����Y�Q�v��t�e<�F��Tɵf��66v�֜��k#۔����u4�FN10��0$�:��(�� <=�S���K�ٹ�=Eq�r�B����O�u~��Ov�mYκo�Cb���{��Yr(����͸G��ݧ��h!��p�wq;�T�����Գ���f+A��k�����7�s�V��n�B��4,�	�\ȼk���7�t=�LF�E��x��ȝOM>�ނ���42h`.�������0�:`3Z���Pxm9L�v��U-���z�Xյ2��nd8��Oc�lJ����.*w���|P��ɔ�w�����ͱ��/ut��4�O>�q��´�r�ؗ9�����T�-�1������\*�
fA�g�`�y��X�
�+����r�0��ڸck���|��tCwT���]O JdD��#��Ψ&b�5��dNs�΃�
&)�RG<��-쑢��dRt��`!����$w�����P���O���t�v�B=@w���L,\n*�T6Y��WC� �u$_�f����e��5���j6��͘ðΏ�ON������I����'�J��]��8~{����0dܞ���ҕ���yk:��xw˥7�ۀ��|.�Ǟ�l[��}����X����t��SM�A»�XX��0���p���c��gN��;�"�7)V�y�b��t`ج�N�J�C�{۽���Oy���q�3�\�1�@!a��:�+DE��}9 ��WbdCv����wz�:����p%�=�L��<KӒB��&�5�.�sѲj`"{e�l�+����/�A��*�JH銆�b������H!����l	��U�a�Giif�WSs�L�x���K��� Wϥ-L�g�d�ƺ��y3��g�g� =�_����O˞�o���킍��|'�wr��@��B�s�u�G�ޙ�����:Gt��=9�'�T��n)ˋ쭱ג���Hƽ�xF�Һ���l��uyĆ�vE�9`^����]�J����pNNA�Tu����k�di�����q�g��k��e�M�[C0��_O�f�Zg�j�wJ(%�3^6$�Y������*�O��\��-Dc���~i�M�0�=���e3���>�;=T���� [0�k1E��|r��<��)eLe7*�cK.��0�c:e�TH�l7A܁ב?(��M��voY���D�Fݺ���A[�s������^@iJ���ul�"tLu-�o�.�:�,�!˽��fm��;�.ov��p�0�,8�vh�Y*RO�;:��~�}��	+���C{�p=¯���ZYi����x�\{ �E�3��D�����<=��3��is�tO�_���B��>	�p�z%�܎j�����=%`��z̍/p��mj�/��븍#���ct�4.y����ZS�sԑ��`&{`�h��U�T4o;$����"�W��F���5�S&
��,B��%3����nr�Ժ䮷qW�)n��"�Z߽���זb�ʮ�a�i.�D�9�XB������L�"n�7V��Q���\���I����ԥR�U�ޒ��O̢L6uzn��sĉ�	��wq{Ə�� VfN3˹�>�N׾��+�Ҽd"��L P�1\���J:��۪�c��m�;����.8���}hh���Ȅ*T삪�x� ��t�'�^?��b^}��]m���ئu��6�6 �e��Y��BuE�g�����p�M�+�
�:��ݣN���b��D��rc���`w���4����].��g�y��Kc[�V6jH�I���Z�~p�*p�9$�
�Z���U�+]E��ʾC<�O�YҼ*}T�2��'��zm�ez��n�pCV-�*D��M�l���,�qp7�H�6�u��x�Z�Li��ٓR��,��[�:5��f�;�z�re	�YM�XF�K%�MBypс�F���հc��εvW#�*���R�@$�in�Zl��A����T����������S�e���DW;�ZBe=��&�?�dś���U�qӚ�E� 8�>=�[�;�V'=i���M�f�'/x���$U��652+flԠ�rRj�-�W�5�9���Z�H�˄��syNk<H���&����Y��91+b�9թ!�!���ܾ;K;B�	�Q����s�t��ɫ�¸��V��P9x�J�s�j�9í�V�`fE�p�f�u��\N���1^Gy-	.j;@l�0�j#6�R�М�Z�-��}�#2V�+�;.�^r���9�Ⱁ�J���
�z����wٶ�����4��0�(wVp��{iN�z�)p�ph������w��`�ԅ 
l��u�-�������(�����b��*�ξ{Q���Nt���6nK�ϴe�W@���=��d�뾮���
��;0�J��O�)���sk���[vu $�!�̛��ZѼy�J��L����1��0#��2P���_�H'��zK����w��w�ND�nI;lc՜k�Lf�d��K�$�%xr�=��6)���)�*�Z���@�P����ځ�IJW��a�wu�V�ƴt���]p�i��N�LdV��z���P�pC[|=Z��7`�W�kj �R�I��G;�"RAy�P�r�1ft̕���}��\+y�t�&��Q�d�׺����qG�����#�X�`	�r-F�c5o`լZY{�@([-@y�:,��W�9��A�.�J'.�0*81�b�7����:�u3@4�3rR5��q��p��ދ�%�u�R�[�M�lV�9�c(��-aC][�M���!b��׿t˔h�w*����<���x�s��E,���L��Hfvu����ָ=��}�p�2[�գc���1)r(��_Y'�mo1�yb*\�H1�ȑI��;ғ�=t�Щ��nQ}Ρ�Ǯ���L�&�뜪A��8�C��B5LީGf�e�[�]��늯mm�X��zݙ�wC�l��jGs�IDPMA�%�A.�l3JMRԶ2��<���T�J���fYB]���]<��S�AS\�в��YW�.Ω�=)�j�%sm�S�}�5gJ�j��W��^;E�ZM�Sp��f��H-6t�X�`=�VK�ʅtT������/q�:�o���(��j�j�0���q�1}���ڊ3+��ʈ�Mm�<51}6R��!`Wu;�d�=�*(��بʊ�-��9j�|��s\uvJ-��Z���mi4(((
�B*#�QTD�4��0�H�8\��\�Y!S �"�E�Ȣ��c�i�A��(*�qZs�˗9�+10�9/T�^�jE��g"T�)���Q�G����dd�e+TJ��P���UW"� ՑP�
z��A\*��*�"��Qa
��I;�(�s�(� ����UTQd���J* �!�1ݮhUHDAt˅T\�1a�QD������$���ʫ9�K�"����2�"�� ��9�.��Q2�rr$kB��"�C��q��q∊��t9�l�p�ʪ�"��uH�Tp9DDW(��U�#�
�s�
"�Dr(�Ç�Q-4�*Q����(�W*(��(U�\�*��N�U�,�������TD�"?>�s�u����}�_ݿ~}?}9`�Ge�5N����0!{[��%5m��y�_]$]N�G�J{�i�9݁����ڪ����U}U�S���t}�īҁ�9���)jȬ����7�>zk���vxO�*� N6�[��8�������Mޮ��@:�˼juʍ��-B�.W,���-���p6����(v��M^v�zd��k�R��P7RFs]|��HQ�WWB�K��E���P��T́&�]�ɫ��2]��}�<8;tDr-���M_���i���x��\<<z�B��r�k�;���n���Fg��7g@T��;ǥ���r}p�'M��n�{(DȎx۳ȍ�z]�L�k�x'����
�,��"=Թ�����Գ�_-�1��'T
�6��=Y��f��T�g�
��C���:먨�
f�*�&U9���)d�����^((X�]3�MN]ϧ�*8�\���=c&�	w.H^��h�!u]2D�Q��/$�/hggn)>kQ�	��a�RP��B+�gН���`��f�%q�iʕ8��F��Sg��7f_^��±ңcH�|j���ho��eH�L`���\�b�>�Z,uf{7a#W)/m�����c�x�+"��8LDt���W^�8��tK�+1����xJ�V4���7yb�Y8z�2:Quxp-����Ҳ^N���[������gl6⤗�]�"�
z���-1/�_p
%ׯ7���E���حjŜ�򩵯Y�s��	��Ek߇�=�{�3So��{6}~���^Q
��U�t=.���ʀ���;6nH��.�e��'8Z�4��d��m!��%n�*"**��g8��%ƙ�	K��fg�.��O��Q62�{���X,�[�Cxq���(���i�\<*��`B���N�0vcr�L�0�γ7x�(b�6�e���������ĭ2��պ���XVM�b�F�.�~������.�Ab��{h@�o�nO�u~��{�-�G��K�=uv��AHb6��t,nuwZ]�1��gC b�E_:d��sb��	�!�7��5Ǵpq�A�9+�+8�|���"^�=G!�λ���;g�&As"�5���ޘanC��M|ԡ���®����36�v��1�(Q48�`V���ɔa��1��R���2�\uʣ��l&kQ{*�_J���X�n'Aqy�,Н���eGx�����ɔƷ>z^T\�o"N-<���A��7��J�qp��K����iW%þ=�y\���}B{R�v��R.������f����ck�є4V���%Ɨ�]{�'�x��������)���N�|8&��7������"]���^u*����_kY��t�;s�0���.Rǁ�cmM��b��y��tڴW�興����]���T$E�O	���`[)����_`�%q�!lω�تTD�&�vT�Zq��G_���f dmvP�O,(���#�|��/�LlW��2):sp��kU��Vl+�x�u�p�g�騠�xs��;������UP�jr��p'覨��B�<'gU:��Z�C$������9����Y�I����c��"��"�QR�v�ș]�;Z���<�TĎ �ӆ�V�_�?N)�w�C8�3]�.���yI��Pv<��ڸ���S��]ֈ�F��9��䐣jj���*0*�卓_0����jt�Tv��Жn�ͻtmpֺ�J+�9�����4~��#�ٵ��+�\.3����:�O���1���Qp��3s ϻ�9̔GAa��E	5���|$��e��޳�BD�|��j�J.#[��/&0`l��f� Wl� rsiٌ��a��9#��m�9�/^�;��N�Щܞ0�{�Y@��h�-f����K�i�z��<|B������܇����QU���s����^��J�;6����iN�ɍ.�+�ɎN����t���iχb�R��X�{��t{rC��]'���[�A�'��AY�.�vl��ڭ7����N���C���=v��46� M�VT=ECѭ��Ä> �/X5˝����0�'�F�6l�x:5�߲gzF��힯e��gA�b�n׻9�c�o�M����l�G������w�k�V+��Q@q.���.fz�8{��
�\�쏆���9��H�6����bo�2���埮=����Sө.|�i }Tz��p�T�r��P�dc)iQ`�q�`-���[ȅZX���'���ɪȓ��v�A��ت�{zSY�T<�
�/�{?p��8	� �79������. �ԣ��kŕ�Omm���עb�04�r�Cg�����mBF�ħ��ED24h���]
[��Z�Y{U*�URݨ!� 6h��U�LH�*_�v���D,J�Ζ̓lo�f�޿���"{ò�\!��́:�hƩV�u����=f7�!�,1��[w3�
����Z-�t�V��u3��G0��2����?���iS�t�,�z�i��������w4��V�:3�H�>Iճ��Pjr"L`��醘���6n�u\[��{طՎ��Y���D�b�&�d�a�`��b�7���$$PS�NR5�PZ�!��]�G�W,��F�����c�-�}��*�n+��@����1��=9S��C�k�Hmq�J�s��՜�����q�5戩A�l���F�S��TN��m�w����<=�{��Y��vou"�������
���cxȆ�@>P�u ��AL�.�"y�=��ฬm�=I�c6�6��FH|i��������hn꡽t�s2h<��zBOZ<�`g�0�³�c���a�N�΄=�=��TEGK�v���D�'4gv��%z���X�Z;�~�k+t�:L`��eAŕQ^��V���gVl���
w�c�B9�`{��~p�~�ފb��ܭ���������G��yd�~�
g�K[q����Zb�}��'}��D�䯸�m��r��ox�㔢]�d�=Nj���^ʭ�\��6��{�_e��JV�,�Ӽa��1;#��u�ԋ�W���g�P���J��z�5�sPֱܤ��c.m�����Y�&r��%P��`�[�Ԩ\��˘���l5�S�t;�7Ԧ�{�3�=��T�G�R!���z|[QB�<�i���a���~o��v�Y��7��â퇢�`I������#�1��.��W���*�@E���,[��(�.��qEPc?)�2��wY �GIi]i�M��讒N��`�?�o��|�곕��uS������icx\��H(��n����/�ۄ��t�]|�K�w#�[�)�o��	S"+�u��r?n���T2nvJm�o�Y���{��{١^8�V�D´{�׆9�p��@'��g��{R�Tj���W%yZ�ve�-�ͤ�t��q±ݡ�T:=!y5�ME��+���y[M(���'�'>�9n�W���ۣ�w'6w`��^I�Qҵ��{;�E�M}�o�z62���E��'';mk�]Wɨ|�9W�����[��ݬl��W��Pi�E�*�fc=��%��<��O1��6�FwcC�Rr�mwg����z���'Wk�'+�L���;���y�=w#�i+�9�,o�˩N�U���\v��,��>�cmx��M�ޅ�����Wo8��>�i;9]�m��]���/�Z����?=�}O�*�2\b�t�^�6)��i�5�/�nM�7�^7s�� ��m/������y�O!WY�>ņv��,��fߑM{];�yZ��n����SQ���z=��-��׽�@�|q��xB�c̛qXW�r���f�D�:�9[Zz��֚Dݤb�N���qRv�B���o�0i|�<����1��1u�7p�N����s��h%N�]�xߑ�}�o-��"�CW��g=��6�vϊQ�,+yՔ��u�R�щ�!2�G�9�*�`d��_boվ飌\�����F���:��m侣f@��T^V��3O�y-�|�7}]��0-�vYBOH-��X��"Ź၊׭.����i�o�v���%:n�c�p�#Cq������w��ש55�1��!'v1�v�ל�I�����:Y��Җ�8�y_D&��m��e���s�3�Z������C��9��ûC�t1���Oo�+G"����^�Ь�}����̸	�^����K{L�����9���+���l!kp�;�И\�%��F�>�:؆.^r��!,�tj\ՊOIL݊x����>�S���&=޸�Gy��O�K�;3�e��kυ�n%o+-;��k��$+�����}'%;�*KM��SoMLmh�v���m6- �l���Fʌ�����+��ّA��g�E��@�9�,�;nݪ̙��ٝ�	�f�z��ѓ&vQխ�'7fi?�x �XA{й�$7����l�)��{�@ۣە��l�9�w�D���r����N�*q�mF�kOu7|�(Ɔl7�-X�|ة�C��.�ݏc�����z���{;����b���5��<-�F��{F���k��xW�V�\HQ��ݥԽ��MOz��� !vzxi�yy���I�>��D׹[g�M���x�ʈ^�]S��a5�4���<�3[q�6�������EPy��UF�4V�Y��&�ƴM��K�b�[Ŵ�&�/��/���ܫ��ʷ�˴�5�ץ�kb���1�Q��{j�yWG�X��˶V��[�ݩ�F�V�a�TZ11�g6�8I���'B�	`����ƥ[�W�<��k(vnS���n�)Զ�0�V�f���>���	&خk��5.Җy$BOn��KƉ��Aޱ�a�FNʳj��k3�80 ubjZ��L�%,��u�{�bc�X`�S����vҢ�6��P(�n����yPht�}ƻ�L1�d.[� �J�-ibA��m^u���9�a7�Q *<�Ņ��RZ�ۨo�N���M���x <.���^�S����M��؀���R�>U��^>OqJ��sZ
8%N5T1	��ɳ��sc��r+�%\��[D.�PD��嘎F�prn�]p�^V-	n\����s��L�AyM؉V� �Ĭ�aZ!\��ݛ�����k�W3���C�:���(v�j����Zc�A}���\V�gM�3nm-�_�UkL�Κv�'���P��
�hQ!�[\�sZ7u�k��5�Jg3+�M^Z�Ǻ���j��n+9����c��)Ym)Kr�m�[x*���~-eA�u�uy9Q��oTo���ѳi�ך����%؏u��:V��� ��u�W�P\v����]K�l��Yj5�t�m��Oᜡ�V6���j����[dx�s��Y[�H(yPa�-��w��/�ǜض��;�N�^A�䯸�	�;����'�xj�ԻX2w*�=$���r��WN�j�(_,����b�w�Qh)�gH��s8���<Ɠ����xU�DYǔ�d|wڻ���_J��ac�j�13U�����
t�.# �n�l�s�G�	]
�\��G����Ӻ��#�C,/�xz�=��=��7�v�՜ۄ�9��<L5���vjxyv	z�1��]�o����V#S�ΧVSw��6^���{���Wr�".	�9g5X�v��Nv��=��%ƅy,	lO�R�{I_r��o$�3�W騄(�)���Zֳ����0��;�)p��m_l��a��U�J����E�q%�I�(I���r���L@n@��ԩ��ֹ�p�D*Im��W$^����i)	�sgyP}���5��Ā�\�5� ��C��|~㞘���H9=%�)��W;3�|�]p��8�Z{
���r�4C�Z��)\��ڞo6��k��2�&����WɌo���C�R���;Y\	ꩅp�^�-��ñ�,�{����3�k�''���{��}�ɯ�'�<�L���6CL+��j>���W��,ks�����<(���dם2�4�V�wr��|}nhw��c�l�>�be���b�
�\�v�nvfe�����4��Ӭz-P@�B�z\�r9�(֊Y$�,�W̞�
��>�U��8Ҷ��$���,:'n�l���9,X8(��������6�o�,wGV6M�B��譩��@�N�����lV��	 F<���1��F�wʸu:�9��k^m���VP���7w-6W9�+}�D�jm�q1�����_w+�6�gjݻ�)u3�ն���0�\V�+F�Z���Q�n��r�WҶ��j�����x�ղ�l��\�n�X�{��Vm�d,��wPش�� ��GD7�M��rہ8�Z��r$��f�f�{4�%s�q�f;�l���V�c�[���U�o0�6���:��>z���]�Q�C$��2�S["��N���q��2�3%�e^��Ϳ���F+$��XU�N�/1����	��W�Ok,X�}�nf�]�v�����8� +�<�n9�cv�_9���#��r�c�Ү�v�5�=�/���୴!F�Ʋ2�d*��Z����@��m�q�N�u#dD����D�5�R�[�#�n}��[ׇ&�)�NHd�6�p�Tu�·��"� ��m���U�Lѷ�*F��Ur�y�w��He\�xk�ϝ^��{b���2r�L4]�<���"��̋E���ʏ6G]��IP�l���6��ZWo�ݏWEKhhjShnK�zp.B�S�vq�N���=Hl��F�ŏ����Ũ��d�S郘��Ӳu�= ��}K�r�,r��[{�@h������2S/
�a�]�Ѣ��1��q�u>]�7{���N�K� �N�TU+�
��>XU���ktz���E�;��[l��������,T��tK3�Rp��^�8��QQv�((
�3,jv>�r=Jb��f�l����[]�QL�G�|/a���֓sm'�KU�wY:�Ն����D1^i	Q��#�o4�VP`1��ͫ���������|��;��i�]5@k8���d��<�X8�J��W�Z�&�Io]l!�8Tp�*b<��z�Q��]����>�h��ق�;|@XF>���r��kk�념M�o����M%e��s�:r��N�Y۷su8Cc����ʾ2F��Q��i��yvi���@��R�M���D��Qa���(�w�����@�ۧ��sf�f�ǁ��/1�Kޮ��N��	,\͗�[LS���Rpl�Vx��w�n���q�5�چ1o�AU��^s�G��ʫ��Gq�m��[�kM��؆��%����_E��b�mɀoH�Ӿ:w���P�n��]zb
;�Nb�x���ɵ��
�s��*R՝i�s�n��<t�'k����h���aQOԏ9n�g:̭�	��;9�����𩙆�bcM[̖�B�k;r��(��n�I.
���ݳ"Qv���{N��΂k�ͼ���	� Ukઊ2�9P�]$�"eY!�B�$��e�;
�.�*+����
".2T�RA
��UQE�JE:T��dG#�A3�ap�PG �/|.AL�i� �Y,��"���vʂ*��VIUU�EDQJ��^��T\���Er��9Q��Q��Z�ETEr��U�V\!�*��%r.�d£�*�\���W��p����2�Ԉ���H(��A��E���^���Ўj9��O\�H�8QL�B�ՈDr���E$���u�	$�0�u�$�ɚĊ�oA3<t�7HG,���P�2hz�8�s�TQt�.DTEETDJ4���
M"�"��~뾮�]���R��S���m�w^õ/���=Ok:��Fj�\�NY���[�7�qKr/r�����Sf�!�J˛����e�W�"�v/��B���-����au�N�Ҽ���FVcLr{�A-�2�GmAn���8��\l�˩��*�GE���ż���	So����7�ns�����1M�5�c��_��+�n�9l�3�7����S�{�ev�˳�=kj��tUۉwE]���P�kd�:�����	����=G��4	��b�R��uz�'���wm�w=�ap�@�[&��.�x��Yi�K���XV�D�c���B�t,�d�O}q���Hk�f�N�vq=M���J�`�����(�s���6	�ዞ���v\g$�sYp�wm�ok⭺��mb�Un��ToHҁ��g+� 1�w�Y�q�e�����MSK	m��v��N{(V����Ѿ1%Y�������ȍ�v#�]�j]�4�J��T;�llúS	�̕9G�]Ȟz��m�t��H�`ݶ>�H����m���b�hQ�N�!�ڕ.��e�{k9l�Vuc��gf8��5m��p�Y������s򾓹ғ����Ly�y:�x��f'�a��j�,�軴V�=sW�t�N͟Z{��M��x1��S�g�h؇�wfX�����{���$o�;�5�df�]���	�!\0��(���@}���{�]�/)���u(P,�훛�o^�n7��i��edu7p�\�һh�ڶ�a�X�-U��!<�6�K�ݛ�Y���͚���Cu�5�q��-�j�y���q�i�܍Ӻئ�r]d���g�T%E�s��P1��I�m��T;G'���Q�{������}2�^��V�X�;�����Q&�4o!7�p��βٻ��s6�&*�5�)87�G�_j��'+�Qz�E�a�����T�k��=K�-��)���=��<��C��ڨ��}O�p��tH��c�f�˺{|�tMb�
~������wu�A6�'��.߈^ߗG*�a��2��;cw����s��&�ZK�U��v��^�Ya.7cj%A�i�^�u�Y��sW	��ɩP6�Юl)�[ffp�=.��f�wsH�t��tTi/p�x�O�-�y![r���]by��iW�zU�j!�[\4�.u�]K5!�k���H��q}m�t�ܤȇe�����gK*tz�Zy��UKٱ[gc����;+�n*�ȮH�U���Ϟ竹W��{�.��4	"����k�gk+s-�\�r�$R��d�����k��Km�myͧ~�e�����}Z��S�������^�O4*"����t�z��)���9��]޽�J,d�-��9[z��Ct!������Ɓ�vX�5>v�ל�\����vO%9z7	��[�Sϧ����	S"���C��w��4ɚ<�19i����y=���s�P�vk�}q>w.E ��]���ך��Ѓ���V	6�%�6�����S�g6^GSv'�r�]�VM�Y��^���i	5}�x�/��vj��{�eBN�
��+a��i�P�6*���p���x��OO1���zy�����W7����f},]�rmk��(��m��wr��Uy���j�ko�����5�|��ռ�9S�w���G�%����	�Q�u�a��@�oK��9adF��b�G��n*��XblYd+]u��	V�;wuk�9�Iy���Y��m
vZ�� Gl�v��z�	��XیR}S9ʰ��u�5��*�wP���7:�%��>������p�Ù�ݹ[aغ��%��*>8����'1{�z��
�X
��V���S�7��}����Z��� �� 7��ns���ʣ���T�n�Kr��T6xrᵍ��:Yͦ�Mxv����uī�m+��ͧ��u�$�r�"��p����K�,c�����mga��c�	�{:���.;>�4�M�ɨY�qn���:���N-ocml�֯��nf���:�D�d��kY��bUJ$s�:��Tv��F>�s�c�a��������;��u�;C���*;*T�boh��w����Z��)�)&�t��n�p�x����a�YRz|[Q|�QL�Tn�mw`t����y����ۖ��}��<�g���$`�)]��TC��$��k;�m�~��Jݔ_$j�c8l����r�[c�E�]7���c�����LB����G'r���n�}������!���+�/Mc~�G" ���|C���fIwx=�w�A�}،��yit�39��Fdh�[��;���ea��Ҙ��/���+����-Q�s�k>}E��+c_�T�Z�=��������.2�]�f\qN�I�����
���Mc���r�VX��n\�HC����>�@�Kܠ1�e��}]ʺ�����8㙛Sb���pα>�*,��L*xr/��|�%z_e�7��m+[w��TU�q|�%�t��4�`}�kg���,��1զ̺U�6��5���z��e��V��o�#:];ePS4������n�3��Z����:Gc�˂����P�g�o.l'���6a������7�^�JOM��w��X�2����$�h���of�<8ݻܵ�4�k"��oryi�"�a�3O=�R�����H�b�uۖޭ�U���¥ne�\�^���^}��*�sҺ}r�Q��lj��Չ�HU�O"^�����L��W��n�)<ѥR��o:\�8���)��g��4����u"��k�	u9��N�6��#��c�pv�i쭏;��S��w9�J�8F�G��)l�ЌK����5m-�Oxs�1���M��2G �/��*g�֨�hҴ9�ee���4#M�4s��G�E)zwV���s]~�_�0շ�6�O1Я^vБnur��X+D���`*TkS��;�ǔ��S�^w#4���v�6��a�X1�۵z��^���;ՙiZ+guhq�ˌ]1I�CM+zok��-��=��������/xE��vf;�k�ַ[��y�O���Þa��nG�sw��Y~罹^�K�@JF��X!��}>m)��{�n�C��2ɜ��k���L!k���W�\s��WGu��d^F������\����Tf����͂R�˧��i��AwM�ºs����"؝�\oaC����\v��$�]Npw9�^7�A���=�i�؀���+aɥ��"��Um=ެ�\e��ޤ�]��qZn:�=>F�K؅m�B�I;Ag�M+���w��s�ŵ�A��?wS|�Qo�(o(�#���3gw��t��y� ��4'l�X�OX߷ns&��^j=����ķ�0��]�#Te�YI���2��z,����ޛ�R��o%=�Dɒ��B\�[�/g&���',��ōy�[D��i��Wse#p.;�\X��#�w[�a9Ƶ
�`+� 㺶��n���z'���z�+���˃hv�7:��NA`�VZ.j2���_;�����S�z����~i�^X\po����\���3��~��A���y���~��c�S f
ջۃ��"Z������ڏ��^�9��x���F����U�i~�N:E,��;�o�{�������Z�|���W����N�U�_��t{�;�b����C�(g�V��Er/]�I��k94j�A쌸��+�$��\�t%%.���t-��yBi\=�����ZC�l�Z�+�*��B����
I F�Er��ԻE�"�u����n�l� �S���)��q��Dܯ��N����"5*��{7��nRW�p&�d*ɶ7m��%�otӝI������;ge��C���|"n˩�wO�{��K�,�]��I[r���:�<Z��<h��CZ�l�tgP˙����e���9�sdk� aݼSBv�b������K�������иm�\5��5��j�ܻh��S1'�9���ӄU�{�t��b6hIs�e��f�����mR����T:v���S簭���wN�Y-�N���$}6ys��/^F�)͘���������"F���'S'5֮uM�����I^6�*eo y{I�L�}������{�$U��U�ˆ����k�s�����w���F,{�J�׫�y��G71�>jblc��\������Yg�`�������b�Jlˌ�\ڹ��1M��Yt��p���\��@pF"���nT�Pr��y����xx�jz�F=�K�e���z��LKt�,.O���!��i��tyo�{H]xPg�򭴻o9��6�p�h�o�wE�h���=�5�'�N5�k/|K`��>Y�5�*��[7���8�X]��ʅ���4��E=����:���h�4Wr�R���z%׍lH,'9\j��ղ�F>��}�������y�	o Q|��^�Ϻ��U�O ;tl�i�pѱT�	t���d�ɳ:`�Ğw8v�{w5Y��C2��[]|i�v�#�q�_c����-��%��zA����{�d�J���{�fԧИ����JÁ�A
ځyr���*�3�����j[ߔ�v��}���X�+ӛ�s�7nob�p�*v�ys��L��m_�6߱%\�y�����X]a��P����X���j�ZV=�	�y�x�	�{��O�o<0�%a�b���@eڹ=/X�Q��?#���x��8�LDX��҈4+p�K�:�Qu���upݎ}[]q�]p#\֙Z�5w�6����hwB{��h7tj�]����b�k6�G!2�����[�i�pW0��j̾gtOE(Y�r{��w�Ӏ��e��N^�ꮝ��Y ������,u��kWѹ��{�5��S�lUCJ\�	"�;,�����]��a�gi���[�	ԘԸH.9�wS�k����u��lU�m�UnQ�g�c1�xg)c�:�;�ji_cpf����|�X���sT���u
���cp��]i�t|{�~a�Ӻ�A�ڇ!0�J���+32��P�Rހ�o��S��X�F���`��@�r��܂��k|U>��g�Kz$ۮ�h�[Q�_ ��_u�e����uYՅ�[�tV,:�|$ߧ;o�*���V?}�/{}��Ԣ�D����o�Eb\|�/��J7�ƆrOkf��.�c�A�=�r�p�*򠪚��{U��S��l[���� ��z��R��)pݾ�Vv�<���w@J�.��U���6z�wH�FXL�[5�����r�.5�ɸk0>�\ޭ�)��(��o<��.c3�5d����[]-ʧ剷�[�������)z�8�V]x�^��=��e�+j�a�I_�ԫV������:93�-��k�u5��������9)�yBۈ�gw��Wы��֚I�]��19l�k9�~0��{.z'�z��-WM�3�[]x��O����y��u��54P��^����KG�� $���A�}!��A}�L-����{}9�8��cB��C�rk4�N�����O��ek���)BI�7��������tՎ�v^���H]}3	��*ы�q�cfn}��f�8�Q]�Ԇ���#��-sJ�������WG!ve4�7[x�y��2U����̉���G�7�Y��E��d7��U�ڭ�4u��Eؾ���i��Ƿ�5����U�\9\ʷ���T��Gm�,$��^�G��!����䢐�`7Vt��h�`cY9�n^��q�]���V�kL�9_GC����^h���[�&�[�Sv�:*�-�
�Ƅ��˦��:����E\�(p��-�Y�NB�lt[#��h��2�1�k���n�We�x�0��tr�u��6OJ�lA|{��.�ڒ��8ІB3���Z��<��x��o������gf����Aklu��)ʝ}3�*2��+��Uڬ��D�3��N��t�@eoU�9��=}-&��(�\��]Yɸv�[����Ȫ;Y��2I]X�k���a��5���dQ�!��y���|���s��KU��Hv$8uX�&�èn�����: p
�F�pT�r�%��6/�;�p�놻����m��b�xc�|�� ꘅ��DbD�)mڽ�n
�e���w(֘�!�	;*^G+�{��n7kz��9kTs���3s5s��۹tL�}�֠��@dU���y��R����캎����K�/s��^�lTn�6�Y��R�!��
䱔l��A�Ru���p)�)�7�»���/U�¦݊c���{z�
�x6�1�h�c��W�8�����5m[�Lkf'���{Q9�H<׮��l![5<��+@X㕵��ӷ�,�y������ށX�ԛ�C^˜6&�j��r˵�\�V+� l1��*nt58'N�c:e���΄OZ��W���Zgi#�{ �lm�l�M��t��L��{Jk�J�o1{U\��y+R�_v!u���ޘ��8��3��v������Rt�f��il�4��JK�HYt.B�t�M����[A7�X�$	�҆&_�ƚ�N��Ú>s�����	��ޔ*=�$�ݳ��b�tQ\w�wt0�+�C6�m�ܧB���|F�'.f ]:��v��xe�|�RQ�u��b��qΙ;�u�pc�j��շ�*�H�T�Q����f,��3M8��DLa:\����H�2�ĝ��q���!�7�}+�ˆR=`h9x�i�*���^>Ȃ��b�[2Lj�pKo,e�9Ic�Yo��ll���T�.p��n���SfT}|M��+�F���C3	�J��v��C]�������D����*�� �s0�ͳlsU);��>�R�z���ZRf��S;S���M�Z�:��jknq�x���u���^Φ,�y�މ���W�	��O�ƵP������[��N�ֵ��k\��{�{ZЪ���-ͭ�f�,;��۴�$�%�/{9��*�r�rq���lϷ޹~��("����hAQ~W�PE��PQ��\��dUx� 9&Eg�QQ�"+�#�U�*��p*��ʢ�2(���u�Qp�K�r;O.
�U�q!z��c���\AK��㨲�r*()PUӖ]�QG;(*��Ep��x�D�i�ӊ��dz�1��qN�n�wX\Oq��H�'(�XQEzzC���Dp�W
#��þs�G��N����Q����G^<�<d�)�zu��\��L�yÜ��'qn����=E�w��I��j4�T���N8��"L�D�.V��+M%d˦s��(+*�M-OW9���Ux�#��(.\�NR�2�E��Y(���	��[t��P!V泣��ŷ�"�fȒ���6�glO��e0<���8>D�r�	��n-�YiՋ�Z���;z��Yܫ�"�O�������c����{�J�L������m�X���ټ���Bu�3hWrR��v�s�8���ʄ�Rj_�r@v�Lu��)^=ա�'d��p]v����H;�R�0�E��N���9�I��e��Ns/��������j�[���f;���T���FZ�*«ǧ.�>w�F+�o���m�7��r�s���ͥ5���A��Y����~�$x���\�UN
Bk�^e�nP<��;��E����[ܤ��A����4&mu�>��mw���ξ���B�~\��r�����'��n��.S�s�i�iRq��[�8gM��u��W��V��bW!�M���ܐ��o�Y�wI-�B�m6D���뻛�i�qI�Z�Û����;.c�Et�.���b5:�T�M��][/X�ּ;R���S�=�j��bj.����{���=�
v��,o�ƃAi��W�Q㚒ꆇ;�v�+��2�{��&���de�r藟j��M �r5o��c���:��۽���?D��y팯R
�I�u��
,w%�^�Ym�(j+�c�;���v��>&����K�����w��\�Ì���F�z����]���O]�-,oD�}�ח�]gJ��ܟr}B��	�hQ7pT>o1r�(̻�p���x�ho�>�p��OE�U	�p!)�0�tgK��-Ns�ͻɾ�6�q{�	<б8�bk����1ͽ�Zږe=u�����{���,��u�����s���*���b�s¶��Zb�������D����5�F�i{͘'=l�:5���/ ��daњ���ʰ(��z���W�Dj�4��x���o:k�=��L,��)e��;7���q���&vsm�"~j:��)�^b��x��Ų�P��}�Q=:y��7k�(gj}J��m�h�e�ˏ��VA�ꈿc����:6�=���r�RB�pډ��;�8�1pS�u5��r�9DnP����g���֞�U�N�����a������LQp�l��/��0򷵽��o"��ǃtm��N��Y��ܨ���/d#�� ���yn�Y�6�9�AT����Z�r�wWڴ�̹��-����$)X�C�k����3�_h�B`{7����6� C&b��oZ( %pn��~��J������v���Υ��z�C���r�*�{��X��,� ՜���3�[��r�.ߌ{���./79�Qn��'�Q��p�k�o�}����=�gHx=���P&��Og�S�9����y*w�����}�p�Ct��aFvz�y.�y���)[��o��(�X"��)��%u�N_(������$�p����7��
�T]��֖�gD�A^	`��+R*��f��T���ۭ�I]T��I�)����ۄ��m��P���:�P�ӈ��p��uiJrC$6�����{54�!��ۇ�&��c��SY���j;y�Ӷ��]lc�'�Dn����xԻJY��P�sf����c�X��r��޻�����]3k��,&�t�n��@v������|&N�=��QO	w.c�f�a{6^sE_y#-����VzOb<���Y9�c�a6�W��E���:׃:����-Η�B�Z��w�̗�&Z6��WP}ɸ��U+N�w����N��v#��孻�����T��Cn�PJVNM�'�Z~����M]�O�����2����|�θ�k��%�5�ߏ��[���5���^<��5���Nn��%�/srM����n�p�#DKLv�%m]��xν����&�oR�!���*�5k沝��������_=���	��ֶ�Z��x�^-���f��J��t�O9�M>Ax��֧Q�[��E=�K�j�{�����k]^NW�>�B����b��j��V�h�хd���y��O��r��7lqZg�w�Լ�Ԍ~����/��y3N�J꧳7��o%Q˳�԰n����ʢ�p߯�{���OQ��>���_s�m��m��+ͨ��m�����	Y�Q*kF�Rɵ�5*��)���pԝ�����e�֛�c��v�>�o�4Eνxzmƭ�۾��K�
�O�rxWax��}�;a-}؁v���UO|�� ����.���7�n�)mC"�(�fe�u�X�j�aK���f��D�U���k-�JV��{A� �	�:6C3s� �j�kǴ9$ݱ�v�٣Vc,w܌	�E9�6�8���v!jM*��9kO.0���ȁ)Z�9���. \J{����<��z�_xFʝy��\��1�V�U���ÃYO8j��&�!+ɢŷ+�:���S���Cr2�����Qk�\b�V����RJ�&���%Ӹ�f�;�Q���'.U�J`BR�d'�av]�y�
�tfOU����]��\��K�t��gx;��h��"��T]"�{�N(�;�c�l3'�RJ�y�򡶹����.6{��w=*/ŭ�{��5Y�GOfk�J;1��x�A��:�A���vʆ����� ~i�9�Y���*��p�p�q�T^fխ8�ήz��̎I�|b�=���v���ִ�������/1T^=�Zާʩ�#�d�j}�*�h����8}��Fb���+��X�[oE��bzoT-�lk��B{q�w�>�(8u�|�1۔��y���T4��Pq]��f�D˗tND��������m��F��[uɱ/��d��{�������-V.].PPC2A;�ye�i}\.=�i��2�1�r�)t9���grW���r=���]p/�Z�k�rT�K�[��[���{��~�'tc��9ԫgb�vImO����Z댟͸����TCx�36� ����?o��❮G�^O�����P�gu�s��������}kw���ӊT;Nf����sͪ�gP�7�n�������S��������Pһ�R8b���z�N�����p�@�F��3��hd������~�m�X��[Gq�ַ*���D��Ae,K}�w-PO�:y�c�U��Nc�;��f�@�{���)Rb��c���B���H����ypd�ؑ'���&������t�\ʨ�	H�J�*j�7�{ \v��Rn2hnm[�Җw�}������s�{��<*.��f8)p��W<��-�����tk��^���_\U4��U6�'.�Cr�úNf�=�@�N.^�ױ��{�����pʇғVk�fF���4m�;_Th����l�l�oD��ܸ]2�]�2����3�5em(��D�����a<�\�C��IxgA�,��4g ���?,m�!m�l��P���r��D�+�g>�i;c��Q7b�>N��+�khme��K5��զ8{�闬4󆺖�_~���i���b��þ<��-���O���r�J�XzOes�*�v^S�.y�
�׻�u�!��}�i�}��ߣ$�������Ӻ}��*�λV9�:�P6���p��W���?T^cި7�+�ϩb�)w��|!�����N�����!<�OE�C�3+�)c�ۉ�=撓�s���P)u/o��e�]����E3j� �>R�y�a�5-lWW<ٍ�/�]Ϯqоڬc���sb��Oo��덐�k�]�]��Z|�v2㲎�mJ�R��uz�'@l�˅��oղi�5�o�dL���6��{c{JV�K�J6����B�}y+���[�ݦv�gm��w5���I-t�Awz��5}h,,�,N������9u4vlS��wT�R��|���e�v�[~}�E�u����U,�Vzd#o�Ĉ�N��ex��A- ދνY[ �r����z]8�]Z���R:���wkA|����g[ۯ]�#7����FO.�B�[�X��C2�˘�AК&\���%K
M����/��U��~�
˔�7�6mdrm-��o;��*a�w[(���
o�e�-mn����-���U����W��d>�e��s�����F���B)�]���"�u;2#�]�N�#L+�_w'�і^Iz�����.����70�9��S"�ߣ�E����=���e���y�ށ(�{&[Q}����yA�D��PJ���̰�gs�#l�vMP����V�����N��8�ߋ��wXw=*7ŭ�{VÚ�$)����s&� _��u<��|�f�%5�p�4D�Lvٿ]���UM��-�?���Wr�kFq`3��\�:�!&�f��S����o TOOeKt������[�����=���*���� V1!*�]P���sS;w�J�0V�׾ y���9��z���Z����7��Mz����b�}�F�=����F=f�;�̃�r����o�qߎ(}3q���h6iO�ЕSe�Ѷe��Gj��5�u>]w]_LV^p�������ر�"�b�=�7ȕ��>�Ox����	�!A�e�ux�8��;8	W%�*Ug���L}���+�
�e�Z�f�l��W��X�r����oz�y%��Y��፩����}�e�Q�c[�Q_:��z��f؃��Or��n�;�[s��:"�}������iO.F�6���4����������.����j�������e���ܨ)x�;7�����^��e.��3{Z{�t�Ms�d�JZ�/���,�����]��
��j&�yt{
��2�C��.[QV�偍H�>ް!�v;a�ڇ�����Udtٶ;sApެa���47S�Q��f4���How�_Z�Kz���ہ���VêS_s�.�%�K�����ƻBڮ��-ba6��}�_9�����j��؉�Z1и�OJ�ox�Q�ž q��o�\�M�W��gf0�R|��V_be|�!>
��;�O^W���q�n>.l>��T�c��M}��ބ�2��W_�9[�B:\t.��x�x�vj�2�C�H;4K�[1@�}�[�s15[��O#@_:6r$�Ř�.��P���b��[����GЮ�Ἲ�Ub\h��ⱊ5�M<�t���ձ�ٖ{u��:˺Rc[����}��t�'W�ؓ��=ݬ���s4mn��+}\o���ж:)�Y�l+�Wbs�}W�wd�h��d^��KF��)���\��zzXn�W��A.�U�݋v_�*p�}�ݲH�`��e�����R��;UX��w|�����v��%z�c	t����r��S|]A}�d[�_^NV'��T�*���t{*{t��+��q�>ڧ��:]
Ϛ2�YQ��u�!�	g�D'�|�v_�n�i�p���~�~�1����Lx��Tg���<T�v���Y��/j�m}�1֩ʋԅ�q<��mg=��Fx�2�-�d���i�Xu=�}N�-�/��U����[�ܴ��[���;�t%5=ɫr��j��q:�Kw�YM��QկX�քM����Xm���ν�<��6׃�@����%����ѫp�eORw���yl��f�8zm�լ�{��b��H�џ}3/l�fH+a��5���)h��e�fT���	l��Ѿμ=}���K��mp�0M��>T�K閺�fe
i@uc{�kv�n+X�DfܡM+�:ٔkMqo������t+��tQ�9�n���1\p�[�[}��2��!1���2�`���\��`6��a�d;9�lp�ѩW��Y����w�m�
G�ŭ�k�V��s)�YWl�N��Ql��8v����B�mڂ���j(��
z��u\b���źt��:�
�}��8�sךzhH��W�yN���\[v�|�9�;����1�
5�&�i#���Lە����c�>��e���ZjgM-\�&���,�u9�y�H��]\F2��9L�f*�)[Uw*t��&a�4un�g$����G����,�45,����]�6����v�����[{�S����qjkYC����2̎k7]�-�']�ߢ=}��#�;sx�@��
U�vf��}�f�A��]�n��/O7��2�W��3���T�Wk���i��d6�S�Qr��N��u�sn��:��]����pn���՘�3�G�B��Փ1Q6�`k�dV���h���b�h+'���T���YJ<:4&s�du��@�����}�ж�/&U�do&�u�(ݛƷF�s&J�#tNhHL��T�}�)4%�rK`�5�\kNP��ͬs6R�y)M��jG�d��n������4�U��6_ڰ�}�2/�_`��0�C���aYr-�"���ؕf�)�j�����"�G��唆J�:Wm�bƫ�],���Z7��,�M���w�V�����Y��S�k��F��rǽy3�+4}�"T	˳��b��I�٭�z���6�%�,�7��j�m6�	4i�&'��x��ջ/�;�f��7�6H�(q��L��j�Ls��. �����%]�G�y2�nB�s�Ӱ�s���s؂���:Ԥ��[�/7���E��v�-�l�\�7tmKw�B:_8��-Ŗ�؇N"�4+*NŘ��v��hܵY�)⼕��Պ��jܵ]N;o��:��2�6�%VW>:��+w7���i�+JtDٹ�r̵��8'E=���\���a��ݼ)�il�� a��C����a��V0���m^��M`�V��W1�=�6slu��U28l�s*5(>�}�e�@%sGf��:�Dg�;2YJ7����c'��T�7�n1��3Fv�z 0�+sS�v^�pc��/���[ǌ���~��T<�`t��t7�^�܏�]N���Kӷ�ibR��7���ͨ'5�0�:�B=�ڻ�)�DF;b��+�y�jgf^GZ:�pGL��L�Md��Z!����A�:Qs�2�<��A�x��s�S�W��(�֊��O��g���*Xh>���.PS>|��j��ծ�&��A;$\U�y7�k�M��h����z�3k��ݾ�.oR������I�	X�ߨ9)df<C�(D�t�QHt�H�!G\�%ʢ-H��*+�$�X�N�\y*�y?tp(t�U����bk�W:z�L���P�Bp%�$�C�����5=\N;���(�yǇ��*hn���"��ǏyˇT��-r	�-�+�(M9�J�"]۸���ĉ�fq��W���N���퓨^�qN��\��	�B��p[s�擏��'r':�1!0�5�%X`�T!E�Q$���R1I5u�9ӕI7I��&�Ij[Z�D���﮳�$�1��<	RL�sL�tʧ�+Ot;��b@��2Bn*UPv��:+u-PMME!�H�"q��Ah�a���N9�"�Z������?~O�.�eZg�T��Vяf�apw����أ��A��˻�ǣ�:�d�}�K��}z�Z��R�D�����/��'?����M��u���OE�;��<r�%���oD:޵\"��w-�yM&��F�w�I�rNҚs��=�j���VT�Nm�z Y��1Y�Trb���rlZ����;�놩[��Snw5�7�ܺU�w֓��?��@>��f)�+rkݸⳓ��=ܖET<�����;�7������˰O��Q@�ȗ�/!Mvǝ4�ܧqr�b��Tj�aq\1tUz�< �t��-0���O�-o׌�oh�;n�J7�9ՑT��T�H�.)���Ʃ��M�;�+O�	e���8��V/N��u���C�����gN^3�����YQ�M�6�k�\�.]]�-]Of��ﱛ9b���:��^][�_^NW��A�Q��mqr��G������I�1��칫w�/V١⡬�]��v�R��j���O��XM�s/ "���95���2�?X![HV1N�i��7t����01�y�Vk]��r!��;�G(�̭��bA�sC�+-��؆�Z<x9y����mD:�
R޿��j[�u�CNV���I���=~���g�9j�CJƫX�~g���7[�ؿ���:?u����?f�16��� �{Y=���B��}S��v����:Le[��j�su>���[�j�_���`=�ҍ�,�ue>Zy]�T3�������7*��3�\&��o��쫅�uc��vWҠ)�)͙�X�w���%{.U��U�o��:Z̆�[q��AO���3�,M��R�re�}'��uEZo,i�l�>n�9B[`v�H}]�v3ٕ)���-���w���}�J����C]v�^�Gi�T�f����
tr�	������'	�=P9�!��)�Cް�ށ�6��GeΣ�L�KV��\zΦ��{λ~>W ;�"�[^!�҃�{�bf-�S�GDV�n�5�:��Q�y�MQ��L��^B�uS:2
YF�հ܈3yw7m�������[��Bu�D��9X+!�#DL4�e�}�9ҳ1��B�Zc��k޸��c�ˈ\w�^���㳞�!Z���q�,\���@�i.n�-h��Mï�F�> �{�jon�b���c�F�Rwh'x���ȷ�R�D-��b�p�J8��gor72�r�CoU}��1���Sю\g����=��r��\�ɸ�{	�H���S�JZ��Q���E&wr�8����W�k^�?V(���n㜅�1ans��m�h���\�"뵾��h\t���VeOM�]J(=�Z��&�x?�X�o8��pݲ�*˜���UDb�a�;f�<�vqfuv�;���9!j�3_��lƼ���V٠M����8���NE\�Mn�Xg��U��ʂT�p.�o�W�w�5<�F�����ַ6������¡�ʡ��BzC��d�j׻o�S}PU�\'��	*³v��cu�{���й��xX���V9Y[Ӹ��c�;}��nFk��l�{��Ni:��s�����Uа�b[QB�<�jE>޸|�T�ʺ��<����F���3��l,-����zzCj)���t��jyۭ��J��;f�&�c�7ru����#�y���uӨ�䳊w[{
��V�T۴���	}o0��3:�GF"�ֈ�G�Pى����}g�__I��-'k��̅��L���oIe�:��\�cW�����+�b"庫8[�V7�x[α��ju��d�6Rvt7�7rz��>������mǢ��ȭ������$�v�J�m�ҘW�4��轄�����\�A��B eU>ogi��|�u��v\@]�q��$�[��l�f��+u��\�}�b��:��+o��W����pk6���ݓ��o�K�j�>=����9�tê鈠®=�ju(��Y����Y^5�W��oL��5���Qu�B́R�7E�3/��Ě�N��|S�c�FV�{r�s��U�kV�1X�!t�����j�mZuU����!EFv*o)�b�տ�_WQo�x2��j��ij�<�R�M��Ük���f���T�)g��9�d:�ޝڞl7!�H��2��[�f�}1�Qc���ecü����&<��ý�ֽFy������{TB��u.�ش����Ѯ)���23�^�d��,c7�P������p�I"�9�M���m^c'���W���i�<���,־xc�]�i,��@�Q\jf�@8��ړ_rݗ������H�p��x��t'\�6B� 蜾�n��t+(Ҙ�#��K�F��h�����<��ɛ|���V��m����3{H]�g��ϱ������u��w%{��G���Jj5�^�BOZ4jX>��B�n�J��z�9yT���;�y��M&�dS}P��߄+/l>�t
+����(Zn��wF���L�T��Y7�ڪ�oy�����]�o+龙�-W�'"0j�3I8�әs�:����42B��c�W�5	4���^úJ��*�BOX�=����2�f�h-���̍޻��c�}Ӱ����=��T����y��F�����F��^!����ˆ�-��ڿC��3�s��H�m��6.W`y��W뎲�F���dWA�&�%��Sa�wu�2�6n�sZ�u�Ȼ�q�T%��C��:㱀y^4��!Wa��:Z��	<JB�v�M�Ƚ��2�!T���T�l���Yp_h��y�qLۜ�E�^ΤXHH�T6���f>����Ã�F�2F�q���|+��]y퇰�]2 ��Z�ݜ��
i���g�/'>S��Cy��ڵ�\귩mZ[,Wum��of���7�C�Їrun
}bc�C��m�6��5T�I���ƫ�Ek�\Փ���3�z��|�������3{���Յ4#1_��|�%yt�V���^m^Nb@�V1!*q���)�mԾ�� ������� ����`\���:��ċÞ�ڇ��R����5�����`tGj�dw+I��օ�U�U�Sy�r�M
��c]����@���*ݯ!���x��1�@�p�����W������'3[��w=~�'׮{�u�Zyhp�i��v�=�3�M�=Q�����o�>���5�ti��>�����s\�����s�~���~�F�6�{L��P�̈́_�L	���^��;s{V#�/��xފ������RѾ�V|5״�?O�Z5��%�Tck�YY�"���R�~Llj�YyoMg�s�X���X���Qs����R��=�Z�
|Ό��.9��x��Tz�.�f9p�f�Z<�Y^��]���胒��UH�>e�W����}�����1~�=ǲQC��a����m;��o��:Ͼ��G��G��;���Q���K|KGٳ'���p�ԑ?}�z<�2r3$�eW�<$��Y�����v���imo�+^�ٴ�嫺��]sZ��˛tT�`���K��N�U%0�֡-����\�Ɏ�����/�}���"Zn���-�6Mɧ%��`1ʺ퉪��!b� h�u�@�=Z%��+����n4��ֺ��`;�;�G
����p�^�� y��L�٨�4����Z;�&�GFz9�5�+�/^�T<�2�w����9�U������L�!;J�,z�Q�i�{�� +Խq�]���E��x}��G[�o�3�}'%� �#����ר��f=q7Lv�?�x��ӳ(��^�ӷ���x�¸��oN���2Ʀ��os�vLd{ޠzn!�=Q�I5�>%靑[�q��ϗ��_(Z����Bw��{'�΃+��rud�\/Pw΁��ڱ�1R�VM��}�Sgk^�)^�G�����t�ǝ�a�y>��=��ge�6�_�rwg��}~��e�w0f{B���m�,1�B6Y=��]f_��D�X,zޗ�wq�����)�����d�6���^�eN�#Q�κ���y�9�g�L=e�f����q)�(��:������oJ]�j}������������{�g%�܅�G>y$v�mR1o��z��sٗ]��}����.7�s>s��^��5��7��x�.�i~�Q���(�=�%�'r��h�7�bx)7�b]�~���yS�aؕj���&NvQ啙����i��PΑ�)N��5NŽ�"�MD\�Xn��,[����]S�����$j�<��]Ht��R� {xV�^���N�TK�O-��+p����'u�N)j�-�.}��t���߬��(�<,�g��3�\m+����M���{Ƕ���D�b���%P!�����`�ag$�8E��*��$ߊ��*��O"E�S/>ڨ^��|X��ף=�R<]z2�^+�=�쭷)�]>s���Yh0�To}�Ez��(�5�7H��
�{�����X+ޝ��T���oQ���<��M�a��8z}>�YRʀ��x���M
-��%�텣�j��m���;^���Rw{�+����G>~��g�]:��zK�gL|�P�B�zr�S+�>���w��m���ә�^g�ވu������(矨#��M��2�P��V	~�Mg}w�"�C0�}S9�s�[�~�^&b��:0�Zu�tC~�Dz�_�3Ӵ�3���
��+���&�᪟T(����v��z��>��=q7Q��d��U�u�ބi����	��g�zUz{>q���ʉ�ۄ�v����z��"��� n&|���C�����t=>���*3�&\f[<�ա+]j�W%18�DbTX]P�f���BO��C��c7j���7��2�	)�	�����ؒK�f��mm�Wp���jf B����v��Ƶ�5����8d��ߠ�#+Dl�x'�I7��5޶�T�Z6��v9V�n1����j@��;5%�܎���Gn}+eV�(`���K��H���۴��g�%U�F;EMr�W�ιА�T���_��F�S�;Nu�pt��#���ƽ�w��V�!%���Zo蝖2�ա�I���v��t�,�x����9C�l���/�\?}�ֲ�^#���vu�\?mΛ����r�ff�*�ϯ3�b�p~�&�z��B��k�����ލO<�g��}���{D�c�1�*<5G�������<�C���Hf��3�=�@־U#*/��E��4{~yZ:�����:��u�b���S������/ۢ�9'0���㸮��u��ɟ�����d5���~W<��'n�v�w
�R9NP��{z�Y�S�(%;P���C�S-��P�N�4�5�n2h����ܽ���^OWa��-��~��W�̳��DS���̆�^U'�zL^k���t�y��FC��?+�B��_��,�9����^mK/�Pz@��Rs/c�������wg�3ґ6���܍�>Ո^'���gǷ��ߙg�]���t|3l��yl��6�|�]�>0p'qU�j	��Ð\�͟P�Zn��Pϟ��s�������
���S���\��!����`�y�3�=wb}An��*e����'�+��[��"����݉Ԁ�jj��oz@�Zț.�Ǆ�=���|$|t>68�Tl,�8�4�:�冷W@�cs��ak������Ѣ����|�<�b�b.�Y�L,�$��{�k|�v�{�W�0?B�5��s~��N���>�i͙h�Ac���=�󼒺������/�V�w��~�ՠ;�<���צ���[<H�߄����7_�r�����>�n�Ewi+��z��z��K�<��5�~����(��g�m��vl���[$���$*�#z�9娃�⹥�T}ޤ�Cvj6�z���^��(�:�����m���χ"h�+�n�&<����[>��v��_��LN�4������y�ϗ�����8����`yG��Yxel�z�ަ%Vw�U]כ�1����O�C���댝��}>oi���{c�a��؁�<�|���S�H���}�{�g��5���z��n$�v�v��y^����i�r��X���o)q9 z���_�+������A~���(_ڴ֋�=�rO�:�aٹɇў��z�mT�u��ݴ�3�i��C����^u���?_����w���%���ᇦB�Wp��ɝ�����ty�T�E/=E��@T}�]����w��+\G��x�ۭ�Gz�*�P�͎������cv��9n�;v���9͙�{0� _���b�
+w�n�l���N��%`R�-E�&w3�]v�4�n.�fR���g��k��T��Zn6�ߟ%����!X*T/���]P,}l�}J�H��ކ��BV�S�ޅ�G5g欯/a�]l�[�.�5����Wh�2J!�Z8IIr��њ���%Vȝ؛�[��#xz���
ĝ̗\�_}�eX�9ǝ�F�TN��jǧ���3��(N�<ۀR3hn�}�d�{�I�_u� Lbe�xc!�[%Clي�Wڡ+���Ƹ�� �o���٢k�zM�NҨ�U���2^�CΝ�Wѥ��&���5�٧ul���^�c`,c�OH�2���r!��&�N���k^�'�[�N�i�(��[��[�zE���L=o�/�>�f!��4֭���t�d�o��'�a%&�a} [ˑ���I�Z� Dtz4���u|�R�P��e����e���J�B=TU�M\F��a�⏮�+-I]]\��U���S��V�EѺ$�z��Oeij�m�՘�y�W��@L2�:�J��&"]��%C�
�3S��6̬	bwq�-X����:�<&6�`�G.�����U�����M�!':���u�Ξ���KT5�+�(�e�����Jgr=��(2��P�ʋ��1�کݷP�Ra�z�t��.��74H�Τ2.�Yu�����u�ˆ�i���%3��m�'���$.����}�g)riusI0��ܚ�{mI���{/�vp��1l0A�Ր����(�ۜ�%J|mp�t��,���+��`#��v��1m8ܷ����|�$��勐gE�ov]�yd}�:�����ga&��OV��E�#�$;8���t<,l.��t�j���8]pY{h���7K�;jR'֪ő@���:��]O'�i�8����fn T{Kh�X 6�9z��R2u�%�ǌٙ�r:�>��Y����fюE���A�6��.t����Z�x(��J��3uWP���� �b�v��daws}La�:Ų�C۲���к�W��e�,H�\o;]���.6�v��E٧Í���5��*�s-�0��& ��GW1�r�/�����S�[u �� ��9I�t���}�l�2O�蹦wQ�η�(vYl�F��Xʭ�D������X���\�x�Pln�(Xm�ȋ;]�[�wT��"�@��m�k-m�ኖ9�rTj���J<����*�n�u�F��"#D��cLC�0����.����`bt!���wÍ�5�1H�ѫ��\-�>�+7��Q��g�������A��7u���W�j���vΊPv`v��FMO�.��T.oy�|i;Gn����@)*�O���v�U��uf���SމK��oV��\Ka�wV�VE���=aL��
y��.M�Q@ŭOYg���f�D ~<1mE�2��dW��xa�C�,�z��mW@��o͒�{6$��]����~�TEP
%J�]� GC�[L�Ed铂Mi*Њ�F,Si�*SjlY&(Qj��l�4Yel��(U��e��G|8�Xh*��!�*t��hYr�:c�!9df�W �I�E˅$Ta��2� �U�|������wiUW�T�N���-+����qhJg.K%-e',;KV&M�ՕTYTpCL�͓)"���Zj���I�s�'E��
�;��<bVG��(�&�g���$8�k��B:�0��CF�U5"�*&We�E�%�IȮ˦Ad�*��I�o}K��\�J��+��#*�NkN�RI�A�t��4�D�.q;)�P$bTFF �qY���dQIRBI:gV'!P���ұ8�J������5(1���U��2H��&KAmݫ���3M�v��B�������an�;�H���۔ft�%jL`7�*Cu��Xs%�D��
�W�c	7K�/���25]y�1ϰ���瞩F�{�㚒�,�H��h�*��si��Sޕ��1L�$�#�<<��J��ZȀ���Ͻ�R��>�K�\z5�׊fEͨ'�\�����^�1���7Hn�C���&�¼^찹篅?:c�x�;�B[O7o�گq7+�>�˄<V�n}d���T��A^��>%��ن��-#B��cAM=�j=�֮驷��O�ϣ�R��#���Hߟ��p�9ޙ�V��|_W����שNNz�tei���wֶ�'7����k����S�x �{l�Q)�������Ǫ"�X�}�F���D
��5�����h��Gt�}������W~>'����W�e�P��Ԥ�L�G�w�<yZ��.���w_�����Q��#O��,c��\m�u�s��ǜ��v��z��6�1B1����]~D�$n��M�5fއy>&���7�ǩ:�|/�\\C�zf%���|�]��3A����yB�A�=g�'�v�v�z�+tøͯq���3Q{lI_��j��B�9Lu�Cu~L�x%ښ.�M�]K��h3�*�
:���Z�" �cr�)��j��H��jK�F��c޺:�<׋l�G�1�̎���u�>W�\v����@�Abͬ�R��Y5���C�#}/��\��2,��It]��."��2ns������PY�s�mh��x�̴v�v���T;�ڭ7_�O\禷�o��i���u��fg���`\y΢�Gz���ݷ�����=E����y�Ek0��u+^������{�c޹�"�ޞ�p7�����N#ݱ�\r>v�+��m����98G���E��%�#��:�뷋7�{G#,퓛1��H^���U�ϙ^����x�;g�~�p��R���{"k���EUw^�y��Q=�ӓ��g�˞G�	�l�	Fһ l�t?z|�����n�W�G���ڪԺ�9UOw>�>�~}g��g�M�SuL
<��L�����O���4n�pF	����7���ȑ�g����H1eaw>��z��@-���p'�n�7�x�ن�ɂ�L5�7>���=��E�*L�K��dh�����mK/ ���77�zhT��~��̼���8���/f��F��3ڌ����Is�<��
�~��\�@��A�����wnl׬{ׅw>�X��vS9�����Į*��_�r=3�J9��#������ߙ �߻�wt��B�y�1]%�΅ǣ�l�u�+1=6��K��+!/�Y%�΂����k��gf�.�:i����cE��T�*5V�l���a^��z��W��so x��*���3)'WQj�=�s��C�3�[�9l[�t�R��.CC[�:�(>��sXv�ޫ���Q��H]B�4�3�>>��qzm���{����Ǒ~�s��o����.�]��)n{�^�y[%r|���G����11MV��|7ycn!:�t[~���va� ���m���h�xk�D��c�d^~���#�u���
���k�/O�ڿK<])J�Uo�
�Ǜ}F�tqVl��n�����@J�u#���v��7�(�;�}y��/�>�Ǥ*�`���{&��M��R�&[��}�f_�/UE���<o�۸�@yG��$��>M�챕��L�g\RJs7��y��N�M����g��_�=��o�'Uϑ���\M�Q�^rI�:�1��Lm�o��n�Y�/�fz��O�F^Mi����i�Fz{:Xjy�o��c<G�[���,Ws�uV\�~��B
�:f���������9'�ueSQ�ZX��g|n#\���;��-�*ڤ�m8�칧�T������{O�^���߼��1��[$+'�a���t��L�7�L�'��f8Ǉ����j���.�~��o=���y���x+����~�H'�%ʉ6��jި{e2��d��>W?a>����핷3$4A��~�yFP9�DO
���QX�Y�4�y�N��ݕ=�G�jk�^�_5E �.�fA��*>8osy�&$rK�P.��6��e>�f��Yr�k�1`��8{+je��R�=J��ǽw��w64�MB�d|��mDz���$��_�[/��lx\:�lV}*�=p�DS���f�3ۙF'�c�o�|���ZٶD�C}@��*�&����?+�`^��G�K+�G�_�g�� ��e� 6FT2#"}��Nl��9�<��>��D���n#���w"6XU���[f=�]/G�Q�p��O&�e@9�����]��|jҪ@�YE����g�<T�s���QrwtD�F3tϻa�*���U��{2�K����Q�����&2"�W��ĵ�����z[<;�L??q���r��O�q����� }�߱�۸�_<�M�r&Z=s >5~�>��z_�w���z���}�Z�����W�Mx����k@
��l
��Q73��͆:�h��N+�<�=�95�uN�+{��L�G�Tn<���Tm���/�@��{!��&��9�s�>���ϼk�wڮ����o�?Gz�;��Fk�i2it��Owc���Q����'Y�{n���yG�';��uM�Q�������R:vٵ���N�Ӭ�z����#�zq���#�o���P\xt_�q�=�{ъ�F����zK4D���bmk�"Vn�	�-� �<j�t�ڊ�mͭ����r;&�qJn�d�8��{%���Q�p'SVrϊ�0��Վ�:��z���,��Wm�6�g=7�Y���yo���JҲ�����K���s�^�M�ʱ{Ey���^{MĖ���C��+�X�3�~� o���`b�@�v�xe��Z�>D��Ԃ��Hh���kG�	�='�ud}UemC��u�� k��U3_{��D��7�[^��o�`~���7����ߟ���^�C�G{�!p�h��سӴP�F+�g��n�~�~s�S�N���p���s�~� �qΪ6�k��;ޗ����Fߵ߇"Q�h
@�`�^��V.��,վ�y���=Z��FL�K�+���Xy]{N?O�Z;~�#r�\nC]rʙ*KڮO`�zva.��}; v�UpSȋ<=�eJ��{���ʫ��Ͻ
V�~�q��j���mx)�mk]��^����z'�h쀕�T�W�-�M�^/r6�T�����l\�!%�8�e7y�h��g��o���;�G�������'�72��^�d���چ��6��ϫǨ��N���������~#�(�@xW�~��1��H��SB����̥K���[�M��^�4�&)�Q]���zv��Z w�̪#�r��1Q���X��J#!�R#翨�6p�w����S^�}p��W�&���z8�M�y��7���Tgu�]�t5���e�y�:"�0gdz"V{^z4�۹��jW��n��
\��O����/���&��R�1�Bn��8,f��R��ٕ�L�����vs#�vKgsL�{����T{�U^+�uW3�;���y��}G����k���.�*�r7�ލF�7H;΢��F�|{��:�׍�_�·����+w�%ǼI���3m�s�^�}��䔏\�G��n�y>'Y�gb�c�4O�B�qE�m{��ݎ���;������s��]x��p"�`���K����V釛>����f�m���r���+���pg�;|Ǔ�,��@mG�]��֋j�@�g�0�C_�׍R{�o�_�ܧFnZх�o����/]���8�9�z�3^��?i��x�>�ge�^Rޘ�}���_m�辯.��j�f���5�3�ѫ��n3ӈ�{��G�+������#��C}��[�ux�!�ޠw�XFMi댙�1z�'7�걭z���>+��;�����u�53a�m�W府����<�DNN�^b�X�ɝg	�i]���·�O��2/z*��ye{�uJ�v�����W��ό,�tU2E"�j�<�~���mL/_M>,tϳޙ�ށ���Ĉ��@�
���%)�u+�n86��e��y�L��+o���r��K���&�	�g�����iq�Y�,�0<ޗw��L|���A�Ӯ����O	�U�u��
�h��:��w���R�A��xҸ�;[m��X�[��[2s&��!טhf�N��xKG�{�#�� ŕ��w�#�* ���j	�n�7�x��g+�{���u笼��uGsw��H�A���}dh�����YRYk�CsD���zh>�u�~:&=]3*x�䐿P>s�+sj<�<J�!׭#��%�G�N��e��?Uz�ρ��|�:ꌝ���P�[C��P��̀|���~5�z�EdKW�7���Q���iw��![�������V'��6ZW��DGAh����v�������>��P,gC~�G���c=;O�7���r�$�)��[����̃Q�TQ9%�ƦnW���j���q�FX�M^Iࢀ����%�ܽ���^�>���;6�����	>�n���n�W���Q���ox�|��"�olͫB��+4���o��@yauC��͚#���eۈ3ax�ٻP۹�"�R��wU��%�ܺ�L�����l���_�rwg�g*c��jM��!%'�aʞ0�w�P���]u�.}^����ד�����oK}����zkYD����g\U�mΕ��_��u�9U�bw6�Ҭ�/����R�}B���l]�U)��ӭd����,����R����"��ev&�J{�X������y�9Y��Snis/�����c��l-�@wt�K+�IqS�˦'�&U�����{���h�]���v�С(b�G�`��s�t�Jo.uh�1�;�f�ͷۢw7���~��F�k~Y���秾��`v$���d�,�{��e ����]�v�we�K�V�p�	m�1���n$�
Y�SY5���ɝ��@Ǯ�b�������0�[Z)�R�T���U�3�g�����Z��F/�)��' ꍨ~8�X�q���g�;�$Ϫ��3q��JKo��v�?q~�q�9�;�<_����p����)��M�����w�%��O�މw���a[����<���������r=��k~�_�mS\�:����fPdl��c��g6�2�w����t��O���d�h�~Wϡz�7��h���ĿW�W2ʸ�~����d�d
|;�\��>9 k����9X�;�,*x��[~��dyI��I��b|��ʄ��ň��D��0��}��=dP��9تTh����r�߂��h���k<'�!�DND�dg�ם��7/�� ��n�E�嚅p �U��(�ϩ�{NA-�F����s��X���F]?i)�i���Uh�i��=�����!��iK㤀���	��մ[�ۨ�7+G��lTo(I���u��t9՚tz4u�Q�88���.������o �v���9k8�P{�Z��ꍫ1�9Z�&��Һ�tس��c&�l׽|�+����t��.PմӚ�WxK.#D�i��Y����{O{��G�׍ǥP�9� +�{l��D��>n�c���~/I�b3;q~y��3]�"�����=�Q����To?Q���q�K����ʒk�|Kݾ��]��KŹ��N��z|D����Y���'Y���4��.��'�q�^�.c�	���wq���[y���]��D{���"Kgnv�ד�}�D�؍s���`%^���^�x���m�r��k*�Ӽ�^�]$�/�GnU�}�8ca�'��Ih��;P�'�XY�Zu�3ݝl�7�T~34o��q�ޞj���R�r#�^��m!#W��g��w���>̯��kƗ�yz�j�ȬMUy_�9jY�:��G������f�wz��������{M!p�h��3�M�=s�r�{ޜ:���w\�s��E�~7��L�S��ƽ~�����e���p؏l�)�.6-Ƙ>�|�o&��f�n:�Zz�~ꅹ2�>R�m+w���N����/Mx�'��0ǅ�����s�Ѱ_Gb���Ӟ�Q��*@[u^~��E\�H��R��{և�3�G�*\ftsvhj��<��5kF�(����½u�ц�쁋���}��;�O�+o���ⷙی���Rڣ�Q&:�YɽEY�
Y�<�t�Y�������m�	9]W��O��d_^t�h[�V�xnmr�Ѫ'L���.��x�0��˸vd�e�ﹴ�ns�����ӹ�>j|c��qN��R۪��[(�¼�se�P�X�0C"����k�U�Ǣ
��=�����C��ǲ���Rc �R�G������U�͆���_��йb/�S������Y*"�n����p󝸙�V����^��_���r��j��=||JGvy����*��Y�>{(�z� �ʈ�uN���o����k�4Z�
ޙOW:����ޢ&����S;���m�Tu��+��L�>�^H����^�����|fvr}���t].�^�8}c�z���${�.V��wǳ�SLv|՛��s��y��S�ї�(�U�e�Ew��NＯ�{M�l�>�r}�_�u\FV�x|:OF��f�u��N����؍�ldL��n���S�}�3��i�X�|�T�+�	Xn$�;s���V�y��=����A�3���#��--��L_�ｫ1�L���q繂�,��t���gn'j�3�P��=�;��Ȯ���v:g��=9Ԁ���V���\k�vu�~�87�h����7Q1�uI��rEve��8�M3�i�7��!�l,�xoX�LfNH�A1J�]����[�)\F4�"i(0D�7��驑��4�q���3����O��0�`;K34�����'Ҳ�}1M
`�3o!�.��n�v8��{S+1�jS��N�Y9��aմ�d�;�7/z=�گV\��Îmh�bS{��Op�0�G��yi�5ѩ��I�:V@�#���g7'Cm9j��`��W�6wb���U�P_7�5e^�W���TVi�j ˲�A���qX�Rw�����22�C�b��뎱\��0m�cT����d|�F���ȷ)��6������tj�AZ���X�h�׉�]CR&e�rW��#x��-ng(b��������r�p�����i�\ywl�y[b�iаt^�b�k��E����1O�'Xz��r���E@нA��@VM}.%�c.��ұ����1뻲,7��15^T88<�ķ;/Q�]F�5��F@��;\���.ܕ�K��=5�I��Y��VF!��;�{����w3�qt��������Û�.�Eڡ�������t��kM�{.[P���n��u(:�V$/�E���v���ׅ%��B���!u"�`�KLO����u�B\fު��=��u�MIe��s��O.`5�MQ�Zs�k�鹖6�;P_%8U�2����L��;���>����c8�h�H�J�����{[z�G��7y���n7{o�1��wv)�_�iu������[�ۼ�4K�7���=h���&�nlE*ړe����d�K�������z�V�.����֧�e���qb�̎�GK6�
sF�dՍAԸ`f����Ż��`������#+��:;+�
E���CT�í�V�h����R�a"#�}.��e��j��bi��*V���I;�\�	(��@2��t4�}]x�՗γ�%-��z'�48�D�c7���-!.���$�D����js[4���J��cU�ai7z8���W��:԰�tV�yi��XW�1�W��aHb�W�Z��ܜ�nALwhTy�!�T�j�f[�[ϴp̒��$K����;f�cW�[K�\v�3D�4��q��p�E�и�>t��HE����5a�U���c�8Ǧѥc}�ipo�iq�f��GSiWJ��M�D����k�j�y�]7����������*�>B;�G`]^|�ѷ3�#c��
U�錶K��#c8v��ι;r)�C�W9�Qj��QD�zP��z���.�&X0��`�e���h7R���w1w��U&�#;&�5�)�s-c.���:�m���f燨@�wy�fZt��j�=�W��k:�Yj�W.�lsS~�y���Bz�j�v�����@��Q9Er(���R(����(ĉ�~�Ey)*yȥ[-L�I��L.Y\#��*hsU�r�$�8����rH�k��r��<�%K;�Y$�px(���"�QL�;I	:��U��E�L�S:+h�)ĸ٠����.�ER'5�H�z������i*-J.kq����L�v�.'Nit��K2��눕���I8�S��qK[L扒��BJ9H�L�!:��0�zw۪Rjkv�'	EP��p�dr�#q�EE�t�B���I%�J/U���UJ�T�Z��8�D�\څejḭ$�z�q�D��(�UQ�Yh�VD&dm�B9�I\N�B�뎙��G:p�sA1*-3�URd��D�,�i㸋�ȫS�V�r��)ݮ)"���քP��PR��އt$�sb�Q��+���/%�urD�g�s�q�����;��j M��=DwKƛ�����]�l$oѻ��u��̅{��<�1o%?�5.�}����p7���\j����^�e.�z�MLg|�ݒ��\N���
��������R֟�Oz��Y5���L�.5�Nz}43Z����W�Wy;�=�8B�>���x�׶�T���������rrp�`g�=����:��mT�q��+-�a�]mƪ}>��i�W3�g���\����{ʏ�+��R7&�SqL	��@��_mT//uya��Z��ez��|�Tlx�W�#�%#���*e ���v{�=sd���8M�%&�v)�I�OTt8����,5�a�腏�"���>�XZ��dh~�W�Y2��'�nk/ދg�\N���oE�t��*��A�H)�0����\UïZG�����	�^�wB����\��:'}��-��^Y�;��{��hނ�ә/ƾx��[V��;����H�k.T��q�"t�w_���=ޭ�C��v�&���3�S��чҴ����l,�R�LV$��R�Q�ʷ��8Z�lϢvtqِi�ר�rKG�n��O���j����Ѝ1�9jwB���<�d��$�x3|�[�������"���1ؼ�O<�����]2ƺ�B[HI|j�i�Ւ�֠�%vGQ���ƴ�u�V�1AK�:֚x$������d2�\%���]6x�[�x8@MT���R��V*�r�9�n��a9���c�:f�]���S�7��B\��3�~@�O�i�u;rF�VA��� I�9�D�C댭�
���OW��ob>��y>�w�p�P�f�.9�� {�T<-͚"��x�(vi��>��G�+�]�f���E��u�<5��m�_���dg����ݙ߅����o�m��:&��}+m~����;P~��-5������̘�����g��,���#�{��+��}>x.��V�5Q
���Np�$���r��Ӵ�\d֕��p��Ζ^���Ռ�7ݱ��}t�b���VZG�ݞ��gdZj~��H����n�<>���������I��&����}];��9~�$z5:l���t������y�R/�9���?�t��L�"�C��3V�H���E��`W��]����߸��י��x"��:�%o�S��M�SsP���U޵\�;={Ѱ�O놞Oh�������ڨL�S뇃�ߴ�y�n{>�W��xs,��"W���{ђr��ʖ�s+=`c�Q`MwZ�S.�&�F�?+�g�z�9����|n}��	W��P����H �a*�>��n���ڝ�CVG>6�2v��9��F&=b1|� I;���i���|�L�v��� �
E��.�2^�x;9�z¬�DE&�5+]����oe�V��[ˣN�q.R����]�MV�����k���*�Bw:7Ur�3�˳W��� y�[R'�q6�3���w��X�M���<z�|��7��PB�h\ve�u��>ݽ�Q���"	8�Tj	^++�4�%�^�r��紵��r��+զǣ�R>��} s��d�\�.�Ah��10�Qt����W��-���(isݹ:�h�P�{��>sRTG��T{Հ>��&��s-�$�b�&��F���`d�E�})+�UD#��g��Q�6��p�yU���L� {�`W�=R����Z�����bg_m_W_w����
�rO��>��zz�Q������ �d��?N����j������nU^mIT�2M?Ѭ�Mς��������cL�|�X��y�^�.aDo�Q�_s�绳�5�Zq��ίf-�w�{(���/NI����x~��wO�2tV�:��3{L	J���?y��!��s�3y�@��(߽�bn=�p�}��9��2}Ņ�5�Y=I*�����'�ۙ��#^`{:�.<���ޭp��/^��q碻�D�a՟UCÓ��<ǣ��ף��R����֣���#��X���N�oL��Ã���ۏmT2��f�۫��^��K�@�Ù4a�����O�e�O��b��jWU�s.&��.^�.���$ߟ�rǒ���ر �a�J��z"ժ�ǻ.[�VCR��o/W���N3����������U�fKBgqG�ʿc�5)�ir�ɱ)�Z�w��w��O}�@L�u;�ֽ^���O�_l{.7�����Tt��8Kae)��}1<�ۙ�&����Jo@�οBS��ԯ��Vw:����L�Gw��7F9���T�<��O�_�����tE3s�۪`Q�F\�H�FT�������)�:�;�E�,��O��l�C=67�wO�ܼ�ǰ-�f;#\S�pT���G�l�v0����,Q����oh��P���W��3M��=���Q��o���!��zwT��|W�a=6{Ν��^��%ؿ4�k=
�Ρ�h_��ԑ�~�@��u�¯��E��^����$�]QQ9-��Ԫ �Y��V���:��r	H��	�x�i\U�:����O�������yT�IK���£�#7��>K�:Ϧ
�H�S�w����2����G�����x�NJ�Uo�;���w�i�W��̥���t�A�#�7^q��=Qr���w�P,c�;m׍�$� hdm������NV�ܐ>+Fun����W	�Ԣ�O�� ����j�*�6>���
�����F�ݓWs�7�W�{o�����2�5S��v���y�t�a]�CE��]C�r0&������&{���b{�>�gم�x�iT��(�5-���]�KT�u�>y����N~���Ɏ��k�|Jӑ'����CY;����8�/��ǳ�wf���z+�ª�GI�a,v���b�}�c��9R� %a�/���B�N��f׸���E&mg{n	����`3�z���w��E���3���֋��'�\�Gnv��8���Nǽ���V�w�y��7���ζ ��v<z��;�Tj#WV��{Mh��<v=h��8�W6�����ߴZ>�}:2����JW7X��>�׫��o���=���#~x�*�n潩n�{�)�K�1��27M�V���UZx}>���� |��C�z��o���fc	��}g����}����)(��K%������Sn{ŋ���o��6��Q��VOt�<#D�c&ϻb��F��X�~�3�~�"]���~�Yn$�*n��1<�~�ˠ�	JW����x��6�JY^��?W���u?^������xr�e�4o�;�ǼG�x�+����kkO��gc������/��ڏ#Qo�q����p��d{������3ⶥ�����|)ľG��\�N�:�2ڠ�TwXL'�l��m�bZ�6�"�[_ Gd� f��q  !j��ã�^�[���$f���=3���'9��4Mv�o�Dƣ��&��K��Y(�U���vʛE�}pQ�-�u�oZ�v�Г֪J�7�Z�s���ҁ���>�چ�CĮ*�/cgO�L��W��ck���f�Ƹ^�m�^�; ��

�ʨQs�r�F��x��\:���/َ�j��ܫMQ��K���
s,a��{,��eS���w�&��L�9���\{Ac*���~�6=��6�y~��']m��x~w]�z��%�Ʀlex��j���������!�t���ݛ��+�3�ʬ������K��%��=vA~���#�u��[ى�ch�K6�u��~�f�sJ��<��1П
^�(�/z����wc����d"WZ:nR\7'b8����A�����w�����&��\o�����~=�_�/UF�X:{�۸�;�f_Tr��9���=��4_�pn����U��N���c�3���{��ߣ�q�Ox�M�� t��2:�u5{���s�x�{K�6���3�]��Zo\���t�;S�Af�-S^�㯍�uwM����P
bc�w.5��g ���;����wַ&��y3�7�r�.%���8����mk�b.U�}W�F��)\�3j�T�3T�6q�m�9/@�:�@G���4�3��6�̗������,<��̹�Y!'�n]���y¬�}����_nV8<���v��̾!�K��9Q��7*<+�0��]d�es�ԭ���ke�������h�ÝP����u�1otSg>��O\ET?�WL/:�Y��@���;�v5g�e,�=N�v5���#��^
�塣��S~$1ܪ�J���\���Y^w?n�g��θ�ᖋ٘^*:�\<�s�i�t�Zמ�_�0L���'~gW8�������o����;fG�^w�n#%2�#Xl�?+�dJF�=�|{�C��^G�V �iP���|'�^�ԫ�/�=G��f���+��0T�&����wK	<W®��c�w�������N7�k:<����Rtײ�����2�|`�n��Tj	^++�3g�9�}4��s�
�ʺ��j��r�����c"=�E�����\g����e9�YG�鉅�LdS����S�S��GUǺI�|�s�����M�2=J���%��G�|��ِEC������� >=�z�#>�f���i�쵼=�t��iH�b5ҹ�W���z}@Nڤ U�`T<�K'��RrT�?.[��?v�#������#_��x}��n���;��h�)�}�yz0G��WޯS��p�av���>z�)���6N]��'Lv��S�P]��$r���6]\#I�d
��!\':��	�4�QB�m���	���Zu��е9Ǚ&�-��Q�`܋`�2�w=�|p�"��{v̏��\x��Aq���fև�|gvX�2��N����ݟLK�z=r[�=��D�{Y�����g~��,�9|��ӵ�����>����\�j��(8��(]g���V��|3��Ǣ�x���#_G�*�[����{MĖ���C���/�f��F�5��Kκd��G�_������@�O"o[�DJ�CF{��Z����[��?O�ʔ�m~�!�[���k�Ѿj�g|@������^��7�~��u�G��i�-��g��O*�L�t���b���,�Ȱ����q�;�>����wq��������>꘿�?k�
�U�3Ր��O��x���r�~�@R���`�πϯ�p�2e9�ͩ^7������_��W���;�98$2���ӑ�W�W�z�Kڏ���q��ϊ�IʉRۊ��Sȋ<=�(?{ԇ�g�y��mvs�_�~���v#�>�q/�����n��H����e�������>�N�ov㲯��7=i_�O���/�{�������QO��Yȕ�P���;���F6"��x���)��W��T�#�,��ff��	�CN�R��6]�6�ڈ�	��N�����tƂ�#�AQ��̳�w��x�gdڼ��%�/�.x�*����3�P�N��#��;���2�l�A5�|��/3;k�V�K�i\{��g��Vd.�󿲒<-ש#�?u ^G��B��_� yJ@]�g�+��۽䲇���������	��z��!�_�r#ӵ����� ��D��V^�>��R���/m���\n&��TD�9�;���2��s~#ʫ��ų�>M��ъ����í���|�=�=�*�<f<jX��Q��V�����FX�N����f���ﶣUw�S�:�W�����S�.v���&����I�<ja����'ä�F��gml��뼌�ܼ�Or��h����<��9���X�C9R��V�Ʌ啺a��.|⦦$�.��P�vz��)@�}�����^�,����ڏ<�/�zkE�BO%��|$z�	P�~��_;��h�9:��3�cO�zn3��+�V���Z�:��_L���kC��i��]��ʻ��k6Y�l�*�]+XEn:�+�j7e ���2j��;��F�7U+�/q{l^�z��^}�,���Dw���P������Lk!9]^��ׯ�ϑ����B5TI��hl��R��?K�>��O���X��C�F���Ļ�_��ᚭ�O�Y�ɋ��.̬B

Vs����z�켒��#S}��睳��8P�������|�Yh�3�߄�<�Y�A�����]?p~�%aXi i>yR�����yֻ�	�Z_���%�w��Β�Ȝ��X=���βifK�y��ʾgi,�=�����o������3��z}+���>0��2���yF����������9'��dJ�]�vya�C���:i�c?^���%#��^p�-2
��;މ�JowK�*���X���RZ�y/R&�����G-����{�nJ����W���2���S4f�_��
�g�k�3��N ��}�@�FKG۳��>������ȏp�����9�;;�>�z�үP�ut�p���IU
������P�+�r��NO`j �JÊ����s��g��4��$o���㠶z�baz��1�t�,c��G�`���{I�7~�~��V�2=;O�9>����;�k�Q9%��u�|Lm5[G4x<@t�\��_�Wz������:-�kŹ�	��:�=w����,��(���$��߲)�^�l��j:if��f/�ާ'B���xhJ��{������,.�x\C�4G�'���D�'��� ���d~qoQ��+kk�6J��
��e�b�u�#�E�V	C	�L�����t��N�Z�7�K. n�mK�iiuҮ��n��CN;��sڍ��X��Z�m�9*|�ۛ>�o�+��;�t<�\b�3�H���Cc 0޻�M��M�
�"��)&���gk۽�:�!*��i��φܡц.��F�ǳF֥���*�kR�����	�|k&��m�'�rn_H,���^آ�����F>�ZB��wQ��&�������L��h\&*�n�Y1qN����qom����j��˦�{����><���U�%��.�����v������qJ�t���ĥ�ʘ�^ok��n[;�Ql��:j���h��gZ��ʐ�R�{ 9�[@om����[����noS2��f�޽��fs��Bky]Yo��L�*p���)t�+ޜ�Tozk���`��<�}hQ��,O{@��2�0����`8�������i8,.�'s�]Xu�к ��y{�]�񜤐Y����pܣ#nc�zn�){�N�<�\�꾵}��\;�EG�VZV,��Z���՜�oM��Z��u�m��=�3���\+����'*�qa�+H{1�S}\b��K�Jn��&΄a
���K1�έ�(�1+aB���+S��X)�9wPYh��]��jE#+�2��2�������Q:�_'.R��]��3s�Q��1g}i��|��b;��	 BM�,�@�x�i���]���TʑԶ�mR\��������*^;,���*�{Oa�.�Y�[9��Zi���n�N`����9B�;�܅�e�Z#KJ�+�st�y"EP�B�1L��ݵ�sb�!�p�c+��©��V�
ʙp�ř���(��w��˩��x��+�;�C�V�sP�S�:9�R}�񙳞d#H;��':҆W}�� >㝈^�[|C�l�de.�-	�& �>����Y�ݚ25b��n��ABd��5N1.v��e]a�ǋ�r�Y�˖m:�0�@�:�	��R�Y��]
�u��t�չ���k5>D2�����N�&,��k/�:�O�N��QZ�C^������2'��s�Ў]�.-��>�坴Ѐ�z<�W�@=W3�A��o�2'�Q��GQw%,�|�;\���x��o�n��\K�E8g�,{�],�a�<+yG�a�-�c{��=���*�;�4d3ծS�V��J}�]vՇYq��vN��t�����n.�(��L��/V�B��ݛ7����U�ƷVs9YVj�=�R�t�{�vv��F�i�5&�7CvT��NX�S����0�힧0N�}'d���̥�*Z�QmZ���.���@�b�)w���M��O�Ա�vv)@�����)�|����N;�&�u�r�&��ە��!�R�f�rD��ф˼�ъ�����M��-�TUkU\�z��Q+���Q��ɼ�RN�K��.���^��D�L�T�6Y®^AdC��
dDt�EB�B8������H��.R��W���
�O9��W	�D!Qp��!�UB$F�����irЙª��.I�)2L�.e�����Ih��hY���dEV���uFT@��jE9h8���p����H��Ü���'e$\L�2S�rn�t�E�(���@�"r����&Fl��,�;��|�A���Dt6\�JH�D��(�5gC:�R,0�W8Ie�Y���I�Fwo �[
�,�jETHZE���s��ﮎKeD�*�V)P�i���AVd�;�$�Дs8��C�	;g�*wpE8:�*	������N�l�"�ɬ�\=���Z�L�B�2�$��(#.�E�Lt�-��g�.�+��� �-V�����s������������%�f�Tz��� �;�L��V���j��v�ACv\�j�Z N�%u]̚�c��,�Cӏ�N���_;n���5I�0z��{���m~�T|E��ͯ{�"���/=�Mq��_��(�	g%�zǾ�$�����Nφ\zp:���,{�o:X�������L�S۹�I�^o��wK���_TSYS��N�D�P۝�3�]>���#}7����b*�ʅ@W���7��|��Y@�NqQ�To��r�'�{I��}T�a�,Y9�k�'p��hіD�;QKo�mz=롷��$^7MߞV��~�C���\����"�ڨ~+�y-V91.�9Ϻ-�*��*�X��=�,SQ���\5���#��@w��m�BPV��)����ū��ڷ�b��6����蚄׺�\a���j�x�S뇐9״�G�[-l_��u��S��w���P�hy���}�=�E+2�[7G�Su�w%2�&�F�?<��^��������yN����"hw��:Ҿw��^��������@�UH��q7�<���
�+�Q����]jm��R�>��=��n��x�{���S�}�^�����0x7U*4J�XC+����c��6:�;�B7W7[3q����x�G�#Ԗ��ke����o��jw]����kK��i��,����[��D�Yه.qR	xF<(�2",N[���|���2fk�i�E���<L[�%c�;��p	U{tˌ�Z���X{ʗX2-U	�{�n-_%�+�sV�_��e��J.o���y�`"+ݜh;�y��"C���"�@C&%g�Ny��ݫ�q<���H�>^�6P��*��
^��=wk���"&Z=�����Wϻ�~Q�z)���Ɣ�v#P��'�\/�U~9�`y����y�~��s����Ot��]Z|�?���
�Fϯ�"��^������'b����f���<���1�+6��o�l�n�-�~c}9RJ�d��3��Mς��6�<�𞍖4��B�c��'��� �|�/��1�=;��'vV~A�+>�S������7��Ie�ȓ�v�k���N������޹�Ϳ*�����K2��~�=���N�`�z��eX����L_�@Oi��-���yq��,9��y�eG�'`\5�ހ�F��},��Vu :1U�������G_�e�B��碻�D�a��]��"��[~��z�1���Ͼ�z�oﳫ��o���WCó�+��r;Ӟ+�ա�ye�c>�i�B�8M�"�&<Vt���KY���}80���߱]ǯ&wӃ�+����^�q�������4�D/η��>�����G,�Iq��0`-���~+�A��Ι��yWPz��Y��D	ً��#��橙ЉY��U:��`�췛�-u����ʎ�Yj�ԫ��*���半���ů���6����R�|�q�=��8��a�v�˳�˗Z�1�}�,�}@S��*��_z��L�>R�z\�q�״�k�ԞW���iYֻ���qh�}-��2᭹e����J ,ڦ�O"*�F�ʔ�슠�y��^��������� t�tg�*\_���y�d�,�dk�vo��U#�2�D�@�7��.3n1�8Ȭ����r�az#;և�y��5�{b��W��Ǿ��\�ǝy�atX�Ҧ��g/���;�����R/6a�-#B�z�8�ԁy����Q~�r-��78fڭ�2����m�����p�x_M�&@�j�hW�WSÐKGv?���Ȭ���o�xa�� ��fM7�:�׭I�m�|�@���"�σ�`xz���N{N���Ӑ�^���*:���߉���egRӗ~hvxWMwj��B��y��'r@I��^�'&a���M�y�#�V��kó�e�{������=H����ra������ӗD�3�^�>�L5��z�7��Q������%��z��}�^��4O�B�p�����jǱ��TG������;P�����W?�cQ-@e~�VW���ib�dC���ss�1�C3��y��Y�ꋞ{4��������/�����5���k�bf*�]=��Gg��O��ٚ�U�69jaɟb�K�ϋ��[��c�6�%,&�FH;v�0��n	��C#B�i��kv�|E�J��<끝� �J�~�O�[�du��݉��hIӜ';�զ�GVV��s
��_�{)��I������?~�[ Tb�`_����W���:�\��}\�����p�8.r�ܯ�h�F=���xv'e��څ�>W7X鸞u��>%_�8��jR��c�<T�{�[��n�O�=�X��"�8:'��=��Z^���G9uz�n�綁�2K�=h�D�Uh����[M����=��;�ϻ�r���%��98\U0,���:���B|z�~���>j|�{��ǳ��I���>gr�O�����o��¿tU3ro����=�U�2����`k|��[^�@�l�^G�U	�Ł�Ճ��)�~��u��Vq���C�>֡m-�P[�N�@Jo9�s7�צ�@��R&�0�^��4jߺ������5��N��~�:C�*3�x���vj��^��5�<������KGۑPѧ�\S�RE?IE3��;1�53�����wS�<�meP�U^��"!��Qϑ���4��+�Wz�M3ZO�:��~輟+|��m`vﱪ,������@��c�b�L��[�-n����V
G+�V�@�o�7L�3��Y�V-!�|�R3���ˆe�|*��Z���W=:b�/�-�v���yF�S��l���]�Y��C��z ¦��N-kxb={����K>o��m�
yT�jG�baz��N{�FDJӯ��]+FS�w�'1nN�<��U�Gr��O����}>�\{ِb�W��o�-����ו�bs�Cٶf/
��}�Ҽ�Q�<7}�Lm��Y:�׊��S��@�z��<�'�S>G^�N:KO�j�j����%�1ތU�j4�>�����x��ȏz�|o�@�������2�x���<��T�Im�,��3c��f�G�g�t=&k*�Wtǡz��7����<;u&EW���^�f,�g��8mxIG.e���'e����Ɩ=�9Ł�b��ǌ�l��mD�%ήέ�D߷�'�IGWLc�T�^rI�7>�6�i���Ү2|+M��F�|w��ߍ#��8�v�#n�~��x��r=��7X�*������]ďY��Le}�ZX���̎u�T���x%w�|���t,�T����2E�jV�]n�+����r��W���}'0�]~�D';��B�y������;,���fu����#��~㑾u�{b�^
�^Z2��	��^��P�f�XA��-���e�N��kB���p��l�>B�j*P�W��O>�&;w�X�[\t�j<t��x�e��5b�n�cw�yЇ��i��m�Z�7\e�n�I�]x�=��6�j�V���s:%��2.yB�Z	{՘Ng�{��9ի����;��lj����T;2��U��J�ȼ��~ӟG�e�F���=��� ˙��gFwT�.W�]
��[+>�H��	M��w�p�Z�&�F�?+�`^��p��.�����RK3aڪ�/���>�O���L��.
��T���r=,y�͖��9�Є���6w�|�'�+��?�+��w�a���=������A��w�+�_�V�ё� o���^X�Ⱦ|��m��Xu��hU�:��A�e9��F{2y.j-�����šh��7s6}ϼ��Gj��6e.��|=^�$|3Ԫ�|�i��Ӡ/y�0�7���h��Y�0=Vof�g���{xߦ@�j�LR��8=㺡���?
�{ʯ�#��,sZ P�몘�2��垾�|����T�o�ٛq�B��Vɭ/O��ؕ4r!И���6M\g+��Q�f���<F��$|�]�Z�Wl���|9�n|�mhw;�5/I�_.�<t�Ɗ?,g$�R��gocf�G;}������n(�{n���yG���^����t��~��_d�#xFG�^���C�
��F�{٩|:�D$1��w-Y� �egx����:��*VK����:/'*܀@��j��a"���E=�n�r��fmeuv�w�=Z�����\���q}v����5X������Ӽ��Sy޶oPru*3�Œw�.���˄sV%~�g�������xo��9ޠ�{��S�T���	�7�����Cɦ<%c��n�#��)������Κ�z�Y���Ul�m�.%�����Pǆp?=�W<�=��e�=֒�S뢲f:ϲ��b��Ѯ@�m]���/�^��K�աW��8)���R�f�<�΃���!o$��}3�M�EWخ���3�����uQ��~㑾�x��U��B�*3|iJ;�Vu{����,wỌ̈�^�����vS~T�ҽ*��/��^7��ö(p�<�����9��p�r�3���-���Eژ͆��+>�Q�� ;'�߀Mo��Gq�Xk�����l�v޺K2��G����lw�z��|�>�]����Qf:�������R=)���{�Gpea͎�I�4O���nFׂ���.<�������DmC��#�
�M�ȀCs�p�4�h��������CW��\~��Q���RÄ�fF�4��f���l����]�l��UA�|��)a ��9�ڽW>���$��jhT��8KGv?m+��]~��N����5�K�V�^����0Л��a����z�5a����{�'�o�k�'�6����O����m)٦�)�n����zr��A��T��	n+{��Y��]�_|-:F����P6oq�-V�|�Q��{V��Ċ֕�u�O-��r4/��S�OjT����d{&}Dj���`��DLE9�;��S/M�k��ocS�eIݚ�j�W��k�5����5&��G��C˯Qg �4z�n���Q��ZdV�����K���83J~Ŧ��E{��P��ҍLz�)�s�<�L��s�V��>G�麆�w��˭�L	!�̪��Hw�{���n�3u0�:�|/����:��f�t5D>@J�r_�Qɯ�{~κV�9t�)�6���m.7�9�f��~J�~�TY��6���P�zkE��eC{鷞�l�u5�<l�D�iӳ����l��eAζ ���㈲��{ �}����Tg��5w��%�|2=�x�̱��,]�T.�=J�Ɩ�n9Ϡu�������n\�0�f�y������*��������r��ƴ���@}��+��_��f����L^�	˯{��c_�9���郎[+O��5	�^G�mjK%������0&.{ŋ�d��͢����{s�ϡL�u�+��l�����=���%ڨ�~�YH�T�F2�b�K����l?l>�����T�ե����a@;��w���=)[�.h�y=Ae<�8A��"ڝȺ�G6���"�.*`s��YM�P�q(d�Ek:p�;LV^����L!}--d<���b�P+AF}�2�J�t��������Mwm��Z�w�D)�*��9ͩ���Ō�����4i����Oz^�dy���k$�sU�V����Ѿ��t��Y���H��+��mCF�-��=����{���=�F�����\�Ճ׻�S�Z���QG���:s>22 �H�h�qu�f�*�s�H�\n���k��:{�w�p��߯�}�Iw���ASUB�.|�d�ә��C�v,=����.�MzbP�㙵"���O���R��G�w�G�#KQ��!�ˢ�-��&�-Y�9��O��P�>�����]^�/��>y{���&Uzb�ҩ�g>�N���{2<��NIh��7P��iI�7�P��P�Wjr缉�}����Ǳcm:�t\C~�����S�.tX��y�J�1��!Ϊ���Y�ƽu�#+tø�]'G����Å�vk��w��9� y_�����1^�Z-��zҔ|oe���Y�㱷���������f�w��̿^�,����j�ߐ�p�m�Y�˶�;>�8n<��r�&|���2�8������zM�t�'�EH�);��Go���ō����˭�u�܈|1NV(娜���)���նC�U�4��"���Sө�"o����+����d\k��蕦�Lꙶ`��Q]'u�X�ȱW�͞	ڷ'�7�oq��do=�goG�Q�枑}�2)]�r���p_g�z9Mh�O(�{:�j�Ο2I�=>�6�i����B���
�y�9��6:�}U2s�T��<:��>j3�<���r#ޭ�q��^������V�>_n��E_�?�<����us^\l"Z>�H��wCn3��E�t�퇕���~�C��mr1otSf�.%GGz�3�3�|�����UF#_g������2g�<J�ᅩz��"5��ܿW�\J�CF�s��/-8��y@ͅ�������)�6���?Wz��(.�B��}P�@�^Ӟ�l��T����״��������{���O�dC�N�2�[7E�4����L�2=I�dz6ߐg��9��?-Q:ǌ9�w�"점�^��~>?�ڔ}�d��T���D�T�&�,y���I3��I�];ލ�m_�O���W�z�1�ARg�N�[�v=>��P`�n�[^�U�^��>����k�M24��ς��Ы�N׋�}9g���pD����|��E���c��ʒ�Mu��b}L���m-9�wq�ܤv��`t�8+;�DP��?�x{ӌccm�� co� �6���1���m�ɀ1������ ����������� �6��01��S co0�m� co��1����� co�01��S co�`cm�� co� �6��1AY&SY�Z��PY�`P��3'� bI~��%u�TT�J��RB�
�� *��B�T��DQ@B	PPE�$)EB *���AUUJ
�*�Q�z`+m��UR��AT�A*K��J�� �+A�����J$ QAla ��o\��*�H�Q٪���E";lw)T��:"�J��$��*�
�$� ��U_mQBREJP�I��;5HP��*J�IR���"(�]�|   d��[k����ݧn�r����n�un�:[�ӧΝ*nj;���{�ʪ7
��M�6L�V�m���`6�:8�Z���*��
� �S�K�   :�PSCƲ��gv��r��n�롧m}�� ��N����h
:8����ѣwp   t��GGEQ�:3]�x� ��4 �q�F�QEQ�)H�D��(
D�  ��ޯ��Z�:��j@vmq\�
ΎQ��Yn�t�j;a�7}��ݭkcm��jӮֳmtp
t]�uR)TAm�����  =��zb���*Ӽ�큘��tp��R[�nm�iww^����:���^P;�vɯ4��W���C�:U
Ѯ��km�9��n@�B�ʨ�B�G�  6��Է��=n�2��jة]���٣WURJ�u�n�m�oV�@iI�oP嶎�+�ި��q�oNx����:��m�Q��u����/PΝݻ�v�ݲTJ����i�"�D�D��  ��{����[��p��nއW��n��cGv��y��;���G: 
ݝ�9���sf��KWOou{��u������v���������a������&T�JQJm�@!B���  1޴У�����ѥ��k[nҘ9�m��rp�om=��;6:5R�����M]�&r,�Gvw�ޚ�e�v�ҳ�ԫ�Js�hV�uu��RIR�D��J���  �=W����p�v��n�tm	mW���/;��M��0�]�z�=n�Gu�^����Eڮ��:4�wm�D��wr�x;��^���]oR3�u�� �N�**@�J�Q	*]�  ��oMnht6�����P�pu����WUӸ��;=�l�{��*�{�g��뻻�9N��
��VB�ۧWJ��n����b��{��Uv��:*�P�T��@�J�%_   �u�f�v�������;���/M#�7�[�:�U�J�=2��Imu��J��{Oe���î���nպ�Δ��[N֋��F�W| �=��2�)P  E=�	)*B �OC!��   O��T� 57���SOP  $�D��Q h�������|�>n��o��}���݌�
�F�_x~w�����~s��$ I=���$ I2B		�H@��	!I��IFB		��?:�?�����7����f��{��q��>�Uۡo�u�.�;ӻ-�1��f�'n1�H�L^фe���{x,$T�i{Yr�g]J �K���ֵH�J�/J5�b:Q�3)��)}��Y4��n[����^�����0ʵ����^2.o�n\!�ػ�ƱL�50b��M�%ҹ��S))or��A��Ct�ͧ X���/k�n�B���%[7�4�yNTn�R�	��i �n��ZNk����M�x�f�y7�'c�����X�R��[����)<���Z�m=���%�Ǌ-�5XH���Kff>f]��\���9�KR�I�wo)�bt���**N�WR�o6��k @�5:^�S(�tC�+ύ�l�WC1�C��T4��v��2��̠ƻCa	M�Vb3h]�u
�mBڢ���ٚ��6��@��-�L�)mi�\i[�e���Q(�	H�1�7��n�k&��wN�+Kq���M�O���xq�^��#�JY4=ʂ*�x�N�b�Nڔ�SwF��|U\Wc���>FZ�,���,��q2@c�I ��F��-��V��l�E&1pIoQ	�څb;b+���a��e��S��0֙����s.��j�0��͎C�c±�RV�
�\"ȫ������
F�k�"D��#�h�t���iMsKVpd�1y�e���N���H�.����Z�+�dU���ǿZ��q��K#	�tS-dF3A�oM)��"f����=W��W�k�C���08ǹQ�:R.STFH�,�.-�Zk�H!�6)R�(bO ͺƍ��mڗ6�L�~BC��z��L�KP�@R��R�bƨ]_Ȇ5��$RS��I�����5�ͽc.��5�TV;�f)�a���=Tem2�&�v�m��P�tJ)�l�K�&��++>�Ov�gm@�����R��S{ᛡꁻ�vY&)�V�;u�^�VF�̠7&弰�D.��+a���Jb�-Kj�q�[f<+흌�\��t)ҽo�	�>�c��Ď������~�u+Je2H
��ͫb��zej�C^���$d:l	�Qf������m�Ke���q뢬̕�<�N<��P�������4B����iz�M���
��k�c~���й��;�1�Q�>�Gs0�lg5�WP��$��m�'%<���f������맄l�+>�2���)��5x-�A�d������Vj}��SxvYI0r�����㣚��)�S�=�3����@���.��S��
��F��t���lR�X(�[��i�V�F�Fk���+%�ҔP��%OQ��HV�:�����Se��nm��
u����"ymTZl�L���dQR�ʹ�6�(Tj��@-ހk�wn4�2�=@6�օm��-�FVS5��Ū-�̢m;8��]�L�50�C�D��ke�"�?��́*�ْ�Z�5�SA*�>��v(���M��(���][n����7Z�
�����u��mֻ�sjR����XvS�f��n�[��l(ۖ���57X��ML�l���j�K	d��U�kX�tv��I�}+Uo�LU���-�7.�8cxMˤ��S-nKt.S�z�f�5�f^Y��=h��p㥓m�+dNK&X�JLQ�D���
��˽݀Z��a5dk�.)c3q�jTW�b�a`�@d�M��)�Ԋ�,áW�t/d)�ж���E#a�@���Dj2"ډM[�������Z+!�ɭ��[0��VM&P����̡޴��'9�r����m�����c/i.�1s�O]aY���VݹRG���Y�S�D�����*�j'�2nbG*�f�ÖU'�`�D2v�4Vwl�c.J6��kZv����A
GvK��T��<)�W!ʶ�-�!�+0�J��!%��f^?�e��Q*�P���mLA�hT	m
m����[j��˂Ip���ccG���w[�4)ٟf��h �S,���A����pP!n"wCvk&��[[�!MG1:4U�؝���ǘ*���A�Iϲ��P�-�O-
���Yc ��53N�KN{�&��ɋ	��U����*ׯ.�E1��7�������i�a�H�EhhƤ)@)�I������Zd�l`��n��[�w�jմQ��j܄ 3 ^��L�D��j�ݛ9��+	��Y�mPϴq�O4�7D�bY�J���Vt�FM�c���M̨�h�
�+R�a���X�����sa'lT�[��E���ٚ�)J�+��&�Г�X֩r��MU����5
��e1-e�c�H�@�T0U�Bj{�Y��Y{�X��MA�H�T�حk-u�JN�X���w�E�ڙ��1L)�t�Jf�X��Y6�� ��%���O h�� R伥f:˕��j���+-Ǳl�Y�AV�*�U�V�.�14�iK���e�4k�xr)������˷�R�h;���ۄU�z6)��(ĩ�r�:��n�OVd
�m�-O��!�J�5�N�U�����rlɢ�W��@�I�՚�u5TV�(�-��F�6�!��;��T�QT������Vm
�[/f�6�<�W�Tke�̗�Z����Gq����C��`A]Jʷ�iب�5��Uj��"��E�V�����r�N����/1�MLr��t��@'�3j�aYYf���٢ݷ���Jm4r!�LA�^㚥]ҽ��̹I*�j^mf� �l�H;��^����S���yw�f\ܻwr`��95�Yh�K,1�zAڒn��՗�������!L���M \���F�Ff#�d�DsJ;P;�	t�%=õ7*�t�����v�44!������yOu��e�}X��]]1Ւ�k�*�����o4��t�h��p��4�U#�+DQ�(�R�r� o)����-�
4��
�t%E�o^�N��d�A��Tp���B_^��o\�|3on�%6����ڗ+5�l#K݊;N�]��Mݓ�X+b��Ȁ6���bv���يl�v��y��(H|\���kYRR�q+
�Ȧ5V1@�n�0x��� ��ku���vܖ�F|1�x[_*˼�&�S$ؕF�Rڻ��B�[C�j!k գ@��ҩ2Ҷ���H�������k	����/��M�+YwG%:�L��AM<��Z;ca�ncMe�uv�`ܽQ<Z
���rK�zrk�ňX�b���tN��UܹF$�)e�Y�T�Y{���Rz��z$�V�	�$ܵ�ks�C�ʔ��h�f\z.�c��NWm��R��֩|B�-��*��Z~f��U�#�v%m���V���OIUi*X2��+@�jml�;o���"ɘX�GaG�ui 4��	�u��-8�!GiCyn���1�6�V��%:�R�݁i�a��aR�u��f^�^�1�`Ƀ(:�n�	E�R�!
����eгH�x0�	UW��)nP�ow�XB��5
�%�P�Ƭm1�k�y��ޝ��n?�d��v�Y�큲�'FGV@f��+kEݖ�)L������Q���cZ/fPĲ���GE��άW��k�2��)�R��G�˹I��K`b�f��kE�d����v�Rʙv��Cd7���Z�Z˘*6��X��`T�Y�P]�LR
��ժ���$�3�z�Wq��+C�jA�6�H*4�y��Z�V�Ne��.T�Sܭ��fe���yR�q�q3�������7Yߜ��X�,�9��c�<�j8��l�� D�]\N��m͗b�vɂa�f��%71�[�2ԩ�,����Ze*+5]хZ�C-��څ��=n�JKFT>WݢF���6�3su��f	t��Y��%���cG5R�O,K�
�hR*�)eY����j�lQ�0�haTC�kL�h�׀�ؙ�A�RX���ДE\Xf�-&�oSo�`�8R@3��1SF��V6���ǂ%�懖�ɛ[Mk��^�O^��Z�P*lr+%cҩ�`��q0uf�������D�%�zc�r ��]�"\ll��]�P2��/N1�IS��t
�2Q�����6N�D�2	A��x���IV+	�P�W�VD�Y�(�O4^�)!Q@Wʲ�ǆKm�c�D 6�-
L��Tܫ�:��!�F@;�[Zl�v`�Y5����V�Kt��MHf��Ub�2'E�Y�VQZ��ʓNH/d�Y�ӷ
sVA��\�i���ZWNc�͔uU���Pl�+��XӴ�*J����m�l�-��:*̲�ghṋf��>@0���%ʆٺF��X6ՊԞP[M��2��t�����f�#��\7S@NF�5.���k�Jf���d�^�DR�݇�`��w����.\w��d�ؓ��k	��V���Z��h��]Ԋ�I}nH��/ln���A^�5ԽU��*�+���J��nf�;��Y�uKd[�䂲��f"�����&�F��Z�-�	�9Vի��֝�ɼ#&���1��v+�h͇Qǻ>y
�P�d��ZwA��˷N3���grevK����қX�آ��I�p�����7-ۣ�eY��d�����i��?�Q
A�xiˬ`��2x6�٘������y��Y�a�ű)g%��f��қ�F�z퓨H�sP�v`���R���.E���C�=_&h��(�s�Z˅�tn�dǃcQ汙�d�>�'���-���K*2�2�@����0Rn:�[�'[��eۥ�j�<�߬JT����@����Ҕ��#/�F\Ane!t���6�X�ݴ���h�MA[�a1�A�n�j�4e��Ju�]GVl��fn�.7KXvҧ�j�fC1$bF7�To p�m�����a4�A��EA��BwX��,JS�-�ͣZUnU�n�j��!,��u�m�vp�V���x��$��Æ�Ve���6��B�ꦰmV����A"�i�) ���Ķ��pwH�7
�b�(0�5x���m�`��00v�+5�l`�ӫ��$مǅ���A� ��� ���4k���b*��l�d�dd���wR�ܖjJ�֩`��6Ƚ�/����%��m�,#*�nn��n���B�F,��4L�4SjR�Mʘ��y�t�"[����@�U�L���}*=��H
�.��m'9��.P��8��n�@�S��¡�Tƒs]](%�0^UȔ��`����F��V���ܽp��лݩ�cʲw�BN�
5�d��H��Gd��SlfݙO5Yu�e��	�U&�/����ŕ�N�EeA�YiPa�$2,��'�Sc��.��RV�ɑ\j�����td���$Ř�VU�	F���5�os.�"��x%��; \2m�beejAH*-uJmXm��V�#������[(��
a?Bkݭz���:�A��H��p�fn�$N�(@�WRl�r����3�4��LAW��ܠN�@XE�V���k�w+-д3Nk
�^����4�7�n˳����W�-"�|��K������.��Jق�<C�q�D��/$��NnE)B���w-��wQ�&�4KݽR��8W�����mf=p�a$ҕgl��d���!��b��vݢ��jtn�-� ٔfmӢ���3E,��5HT�[{�Z�M����me�]^XSSۈfԷ{h�0�J��
�o+2eb3Ne�ċ!�{.�.G��OW�6����a��BĔD!�6��mm
h4�������v���Z��}*�)x��R�%R���@��7oq�F(�[r+q�הƽr�ڔ�K�D-pغvk)�ݖK�(%Y!MKr�E����n���v-�K��nec�uJ�
���*=�oZR]14�����m���C0��&�#���J;�b�j��7C�+HQ2����{��Z��Xb���cĵ��V��p���[Đ�r�wX�ؖ������H���h��M�5����'n��f��CW��m^�y��3e��	5���Sb�P�u2��U:B��t=cn,�V@��V��f�H��:A�j��u�JUaPX�nib����Ul�2��2�<Ne	��x���;W4Ŕ����h�*4a6T�ݪ{.P^;�v�*Y�nf;x�'�4�43RаP6�{n���KҪ��UL�fx�-����u`�2Ъ�rº0e���y����͐4A�!�+�R[�n�wM����n�P�@��R�k)A��jUҩrH)���C*�ފ�������RB����`֜��Z�.�褊� �Y.��!��Η/U��в�A2���cFj���Hޭ	�`�sOn������2�-���Bl�ebִӻ�&��t�'��)�B��ٍ����t�r�Y��%co.F�]{��B0v��v�c9��`d\:4M�n*�5�s]������-�9af�3Z�����h]�õrB$9m�Ƹ��/4*M��k��哊λ�>K^��)-ͻW�#R�P+c���]�o�Z75j����l�2��A����V�DHս��;&뿊�f�,n��J�5�35��M F��2�(t]�$������rE${��cmL���W��ѶE;����6�݁"������v�:�b�q��v��Ԣ�p�wc�ӇP`+�w+ EFE��=JLZ��10�۽Պjy�[�ڭ�x�Vl�S�5ҥ8�"vy׳��C�2�o!�T��銘"3���O��#r-���\�SOR����L�K�N]S%�����c���[(rt�Ѩ����n�%6"{]G;����YY�hG�M�%��$R�<�����Et���_A�9)���]Kt�!*���g�ڕ�����2sv����M�Y|
ٶmFper(��/Jw��\��S������cVgN��u��]n����|�aL�vB��s�gv�a��ԡNJ$�Uj�6{t�1hr\�n�x��[����0��O���d�d�5]n@������0�
��r����i���kc#I�;��*S�ӷm�uj��x��!lĸk���ol���e��P�,�t��U�y*,�x����g�̨�p�5,��]o6^7���pT�خ�v�Љ�HՊ4Ȫ����u�wF�baj�m��5�fA�hpٕ�]��S27�賐\f
J�1A��yBay5�u��OI��A��Yzw�i���N��Fg���z<�{4B"�mҵ�(տ)ڍ;��^�ڒ!On�ac8�j�
�$<�%*��T��w6�m���HJ��3��5?s�fpnc�!h�ˎ��Z�j��I�(0iɽ������>��[��Yc��6�t���ΙO�Z�����WuǷ�:K<��f���׈d���im��A��W�,$#Ҵ��t�=�����wnm*B+�9Z��ۋ����2Eێ��vU�)���X��#4��$-Ƒ����u���z�G���|Q8����M÷,�I�¸�	WF�FFq�&��t�
�|3�vnSj�:D	�R̎�|���C����sN�%�e%s��ʆj���Hێ�7�9�ٻ��W5���J��]Y��.j�Σ�pX����K�k�-ƶ�監@��Dn]����%=�Ef���u]���e�\x��.a��]�"����`<�xm�!���kom,$�����T�L4���߻fHB��fJ-�wGɉ�۶��m'�;�WL���\<�WQ���:�R�gW^mD0+�[���R4���c�twtl��ohW�~{n�<^LeAKëM�:�Y؄E�$�9�ng$�>$_'��V�tQw2m�Ea�:�7)m���XY/ruÛ����]	�͍�l]�PN��RI�<�J����&�Tj�o�Ks�\���%w-J��o��]x��]m)&�n1�IZȘ�6D�-װu�G6TX�	c��rVE�t-�-����t��6P�@�%�yt�U�I��*�X��DL3V]=I�Z7��D擽�e�7�\�G}ݦ�h�Kr��(/O,;ݍwaU�kQ��fj�z4m[�\��)�^����XȨWG:ά�eE��O�R:��
y���P�f��uw(a��ewWNt��P��W�6<��]��(f�z����TR_�m�q&+xɒ]w:Y��R��f�A�<.�iAͲiY����v��^`��u�a%O�DEw���6�����/�.wC-R����c�W�Xy���۠e���h���e-J�փJù*rF;Uʭb���޶�EֻK��1�I����aG�Ӣ8�`�\iWv�����{@R���w��T��fA�VK���]J�{{3��v�Z�9�Z�,���śZSm
�����B��� m�X���h�}ǰVr�󒵱����Ol�>\zE<I7tUuj�|Zٶ7�$�P�y��'Vs��q�Õ(���D����������Fp|FVP�!o���]^u:t:���W��SB��J�1����R5���siԞU��Z��9�����ަ��PVp+Y���ۉt�f9�%�o1������֪�oKζ�u���sl��]n�vc����-R�2,�pu�<�Qg,��Z�u)��sO�U�i�ɑ��n�p���ӺU��fvn6���^���f��W:�؄Z�����5���w8���M��
��ԡ���M塤L��X�ZQx���wm�v�]��Qt��d����35Dh�k��O~w3s2�f��֒�2M�fJA�Ǥ������]AK���ML��7w���pa뢦� ).�p��\X6�N���7c���!�Z���~[H���a������pŵ��Xcr&������(�w��Աy+��J|�����5�{e�9����ۃh�r�f�m��w6�}�]<a݇J��,*�3<B��dλ-��<��m<��.��\~�.]�l� �6ݾR���p4�Wo
рe:{CMTB���y��v!�:���vyrvF ����t͏��Qk�;�^�5���;n�M�䠴5���:m�W|.��ӯcE�W�O_cE&{uꥭ��uo�ڀ�^ufh�w�l�����N���}��4�X^X{����&�|�RQ�ٝ(x�d��f�i�W���ً�FE�fF�[�{�J�]�ּ8��{��ȷ�71$���|6��u��t<�Wy-�������(�B�p�[Ѿ��8���P*w�5`��5�C�AVҽf��D���f �ܗ*�Ř��6��	J�4�Gn�X޾�CE�Bm�[Y�J�J�]WEly����%��2�r��R�ϲ�c*�)������u�Er���}Cu̥P�l�bJ�Վ��������85�tyr�zsf��BWs�y `Y�wv[�[,��˴w�s�ft�J:Ow:��{��T����N��}F�w6۶��Ȼ�iJ�|��6.�<*�P������=�]�ԫ':P�|k;�]A���!����$�q��MPJ���{��o��k3C���[72���>�EЦ2���#�O�ŬB^b.� NP��d=�|���tm�Y3�}n6l�wH��Z���b1o)���X�v�r�F�j�;ݥ�v��z�K���:�6/#�#���K9Xy��EPn�J�q��홁�N�AA���W���	0��]���%F36w1Ώ�>5�lҰ�����5kT���=|2��7(����C@��ĳ�U�:��ci�k�%!['n껝@r��n�J4��N:4�	�>����EAuՃvƔ�̅����c2'J��ũ׻�3W0�]��d`�;Y>��-��79����F��s����}����o�ގc���<�ڰ�إ��Ұru�9m�{x�#th���3)���ʟ>�x-ĥ{��iTw��&n���ݚ��t�d�r�G��k
鼮��V����Co+��vo5t�w9��dE�+�Ci]f�"�T$c7j9wà}c�2�[�p㱛�L��y�
b�	ѡq�Զ�C�����u5],���_fO�.�u��3Fk�9�7��I��؜���a�673�L852���0���'�Ԇ::N��=��v8[Ĳ���Ue�O���}�4��8���Q��!��1%���b_?�Cw�*���k�VҭwN��MUӜW�3��d#4��ɒo��cg5�v��[l#��][�qk2��g�J7����n�;ͼ��|v���Ѫ��˵����8μ�2��06R/p8P��ώR8��n�ӷ�#��-��z��0N�@�sU�qVg���T�[�N�j�\� 82+��8]Ύ�X���Uj�]�����K��n�)��G��wt�p���.��I��Ve.�mq��n4���woC�ҥiLR����q�pu�3���P�2Sz�IhQOP��L��/8��;L�{�V&��c'�c�Af�֨��N��>B�/��z�XTQ��yrw`����ռGR� �9��FX�8i�X'�������N�8�Z1^d:��a}(�Nh.�79w���� �ɔ;��D&#�|�[Z��v\�.BAÆ>�l�Y������ol��Yٳi���뼧���AwبJ?tr�5+sx�p���]; �B���٤�9��c�p��0\�B�9���&��z띗K��G��ʝ�Ou/���xm���C�⎺���
���w�]X�o N����W�F�i�֭snAAt���JC�=k�oZ���(�S��tL�599*����al�ʌ�i;-rμ�e4nsZ7_��l:�ewJR���5�17fW�܋!y��e���w[If�|��ʻ�;k��*[������{�~YS�Y�-�6�>v�qW�ʊ)�z�5��\���@:�+1�����G�h-mu/5=�3�+y �Amה�DG���zOr�K����b<ⳚY�VA��.q�;V&���k�W�+pq�Z���C��-b�r�|H%b�q���S#pͨT}I]�g%�k~���͡˳��[��4A\�c��⛹���U6��/ P����Q[� Q�X �V��c��p�6nrY�.��Eu�6�V��A��f�5/�5�d�s\D�C8�St�͂g�I��0����
P]��B(�"ŧKA�z��L&���8:XP��]��i���p������zr��kޣ�O��uWs�L[�����(�[Fn�l���!��<j�%۔G�Z[�&J���
��eǎ��nG����]g�\�=�&>Èo0��D�\�lN4���k"�b���*c{�vJV��5�F�@�u��u���D�5�o"ݨ9�M������u��'���t0X�KZn���.vv�O�mef5}>��k�vJ���������bҐ)u����W
d��V.��1*�wp˗���>�].�4��:�Jkb�1q�3U�
�󷄌BQ�[cp�����;:,��Ƨx�h����x���g28�x�1�]�n0r\�4b�b�R�m�A��oF1�q���WX8�C�w=h7�yqrV���M����=y\�|=GS��c�e�Rk�Zʽ��ת,��O��f	��J{�)�a_^��uc���)�7��ymSr��sތʹ]�oq��A�(��g�_<RK,"���+�9��7�e��-���F�=�Wb��� I�+�8�]ݰA�����s�o�Z����B�����,���`�1�鈤F�K9�㺻��Ϋ}�RQ��,Mb���Z��o�)�4��,u݃��=C�T,V� �p��u{��`�<G
�2�<�"�#s��=5ˊ��P��H%� �N)d�2�o<;{��ȍ��������T��-�,�����͢k(�L�dsySp3\�Y�u=����H>8YZu�/T�c,>��2h$�`}����C'tپ:�]-U�4k	�E�i흔�"��R0"L�7s^�G�X0�=J��w
� `���R�C�P�6�M&�[21yP�Q�K�|a�d.����a&�Q��tUg� ����YbR�J	�l¸xܛ��k#�`��qp0sQ.t�z#R�/C8+iM|,��辅���'$r�����θ�Dj�;�����`�BY��,4U���H�	��]�ս��}�땮��њ	�a�,�r�s%ƱJL�9��/��i��O�o��|5c�|�SQ�q�����N-hR�x+*�κŮ�d��2���o§2)��{N�Q��N�*��@COT��^o1@<��U����h�0;PHgM޵ �H�c��^�����+�q�6v�z���"��V�ߋ�(��B���^,��=���ޅh��,h�Yf�"k"�J�ճ�q`�cE��ʓwb��"%ڥW���a�-���v�t��&�9<�������)]p(ʻ���w�i��I���lי����"= zh^UG��:�]5��3n��Ha�7��H�s����ⅺQ�{e�`F�����JS7�a���!F�&�݁��gl�#�6�%�<����|IgŁ�t�]�o3���ޗ1>����<����Z��c+��J�c RL�pZ��������	�Ĭ�wԗ0.�"#�u�����fI{:�A����J4鵹��mPQ��V�!�����8���VYә�kGN��v�xx��0�ד��r���+0�V��gn9®27ڽ�|�P�n����)H�w��J�CQ�sQ��{c����}��uǋ"������ɒ�ľ�ca2�.��tU+��v�R��>���f�����Wm���}��D���ldPZ�V�Z)��2;���A�+toy9P9�l5{����7B�sۋ�=z�9s��n|7;�d�Eͪ2��s����ý+T�CV���h�픽�Թμ,<������u�$�.m;��̼gWU�	�F����Y�-��n(�/�X�/v3��v�#KMͱ�ݷ�g:�.	#�t��͊B� 4��nr\�QT=��$��[����P���³����uJpśp�;��+��@5R�K+2_M��4�5Y���L�M�9G��ޥ"��#�����%s�l�.��{;5�����W���cy�
�Kk#��%<�3��� Xz�Öu�Q3�e�N�������-��;�[ 1_Åk�5��1����V/s��ԤzD�
��;��T�繻݈f��8�"Vf���2!,�c����9�u
���^,���i�Ke�Ε��F>}�-�˘fe�\Vv'�;N��xsUu� ���Iz���Y����jCm�5x��\p���X�Δw�Kޱ���}�k��UgR�e*֋M�8�EN��G�.������"���a��y�1��'��Z��Z�\��9d��Ş��w�����%]X{������	�sۜ���o��ݶ�oi�a6���o�ջn�ګ�v�x߼_��8�~���Z�b|����=O���8<��-�i�S����X��n�=�w���������K��m�ƶ��b��{[�����HH$�	'�i��;�|x��{��h��ј��xV�Ojm�N옭�>��=a6*K�zْU�w�l��wó7+��)��q��o�9����+���N���o!<Rm�S)(�p�8�*`,	c���8��w��X�."�NNَ�{�}�J͸�e�����u��d�e�e�ʺ�n�pZ�bp�NA�*Z��^>zk�uk�wK��Q�X��Pc:�a�Ňy}���]���1V�m�g�sA�����NBL�

/�].�r�5�)����C4j늁�^s�� E�d�c�h]v'�ko�`��u�1]���]Z��̾rA��i۱J�f�*�[�zT��z7nܰQ\�__.ǫ%agx��zlZ�*<l��7�^Qvj�\�:�i�/�|׳wt����� ��(����䋗�����o���`"��ȸqت����x� �����ȡ��kӿ���Q�8,P}	�@�<]�Ee�2=ŉ�c:>�&���iR�6�ަ� �;����Nu*�]��.s�t�Y�E�T�O,�U�_UkX�(��Y��'}��l���=���{]i�sh̒3�s}��v��]�yeQx���y���Rj��5b��~Q�����υ�t�o1-�e`��g�w���싳�(v� .gw+O.�𰍾�ty��ʱ�Wv��\�R�K�h˿����}>��7�Vƺ�*�E3�vY�c��M�Q�����xuuG���Qh4�"h�X����m� ����]�N������o 7��-��ɪ�Vݞ�wu���Q�������6W+�Z��q�:4���Ś~��7�C��Ge��ӯ����ҞS�Om���M�Pu3&��g�O���v�I�P���n��f�9�W`�
�	������]l	6�ѝK�tĬ�N�X��Z�SQ�5����}ۖ�(R}�q�uy|�\(p ���|1T���R��NV��E�I��T�tL5es�U�ļ��⾧r�0�;ڒ�Ɵe��t$TdKY�����>DC�M7.�]��"{�����iE�0A�v7�]�ds��v{�JfS,)�5m��l>�+șo�kݽt�,hȷDC��m�y�
�ɣ�5^*�t�7v�>��2��+z�w�[�r���]�.�Sݔ)u���V�XgPg^^4�ef�b� t��#����Ouk�e_hB-�G�o<�͋���s���,��\���!De��"Жv��Z�77�/�ɉ�j5Zh�uɵ���P��*���۪Wj��j����U�Զ��A�1T�3qQʷ�'Ʒ�M�%FEl[J�<{m�s͛B�X-Mn�8�ǖ�הe[Pk�W�[9>���re�]\��5�]/��;���ls73��ԅ���2h櫮�m`֎�E�KОlHn!|�v=HL��k2�~�CjIC�Z�LR��6�����v�r��VҰ'J�r��-r �,�̔s�/���0>8��O��έ��[=8=9�b�������5J��9�T�Z<�����ܭ�,����&��#]���(��2�V��gi�3)j�f>��٣�(�$�ǒ��X�>���G*��0K�8��J%�WX��]���s>�x6�b�}e|�}��}�,m�o�҆���gemk9��i���F.S���Y���M�h�XŊ�A�ܐ[�]�E����Cv�,y��bؚ�ut�}գ��[����CA��uG"�R��mp�i�ǝ-��)�����+w�������l�(�l?v�b�ܺAq"�9�_U�'n�s���]gKi8��q�8vP�4�������Y����C�w����)�vI����A����Q��ur�`7����O��wY�h����r�dw}��*�w:�rZf�5qH��֏���t��-�}�L���ײ ���}́[;2s�ؖn�r�QŎ���ި﷟<��b#oVt*��j"w;��Y�em�	��4 �-�q	R�N.�7Nt`±�Z�������^�\c��W����p�<���A��$[ӵZ}�:n��z��`K�s9ʤ�S�B*���ǐ3qJ��K��)�}����
�J����DT������؋��1��ڥ�w����o��]݇O|k:�]�VWY� I�z�Mn=ڜg-�ˢЗn��7:.��N�`b��h���e�)�*��)h�٘�n�F��b�� ���iC��N�,bgE8!�בX�մ{]ڝ@5Q�I�t»쩷�tM܎.�#�m@7F�z�s�w���!�F�X*�v3�"I���ϧT}���<oj�-p=Ѹ�>KM����v�\�APܼE�E�6�(^l��w!b্̭`�V��'�Ét�u��w�]�,f:�ص.�v�f���7R�7��^��w8�H�e�73�>�	��O�����_t���s��8�;r�W��Ur�f�#��)�\�!ٳJ{�X5��B=�BM�[<�+�>I���GR��+۰2���9v�F��;��J���6͝���S,���ã���S��m3�0��2��>�n��E�c�I�v	�yH(�!ם�r�-yW�Z�mΓp�.�]K�y�|�#w�	Pg��B�"(�y��c�G���I��sM� 0Rhg#]m_R��e�]ݼ�_v��):� s�J��X�m���4O��m@�]���Nd�
��p�P�l�@��s]k�
J�4N�ە�x�й�B0+\f��=���MbԻT���^��-²��і .��\ytF^(��pf��j8;�˕)m`}riN�32R�g�����.Թ�.��:h
�<��$�X���Q�{׆�x�n5Z�X�}f���@�f������1=��\5�v*�����5��2�춷t7k��0wǂ�"�����v�Q��Ʋ�&	q1���'Hv�Uۊ����v�;�h.��ǝ0
yd>�;���q�;}V^][[��,iffa+S��6(K�n�浱��6�#o:u�β]�����	�g^C�P��k�38J�C� ��9mh�u�L��'�#���v�A3����8��n�!��fʓ��pY�T��k
u;0��Y�T7N� �IH�!{���Vë��p̣�V��;��gv�
ɿ�N�E�̤�n>�N�Ep/���λ���R���n��^�7+��Gʺzh��Tf7���J;�e�c$�Gj����DH��b���hEB�����|0��X�R�Ó~��b���-��{{�w�Br�ˋ���=0��/��,ckO"l�aD�.��e̙oP�-(Fi\U���yWݺĳS�pH&)�����nmѫ���5�>5��AƇ�.�
�1�v��;F�R�����}�����Kl���#�垩�8QT�j:C8�hR�F��$-ۥ�6=#p�cm2�"#j�J�Z��˧��l�jWN�^* ��B8�2�Dw*����gW0�v�cg9��ӽ��ӹ�����˫����AkE�1�nl|�w�R�N!:�q�l�;A���dY:뉫j]��9a���|��j����%�\)��L�u����ǁ]9&�]L������uDʕ�������q��oi�(E/�-��m_2���ki�&�q�l��t��p���=[`�#F�ZuZG��v�A�v.��p�\��}���W�V_Z��z����$�[04V�.!vKj�H��ܸ1v����T�h�<5� ʲT*	M}u�j�f+�70�i[���Q=X9���M ooN�UH��j��\�=���������jéL�\�Bv��2�����t�FŸ��f���%���*@ C :h�,<�]vuZD�n�c&;*�*yM�E��$pđU���V�Ɩ䭱}(J�r��ȇlo_os�oY��aԒ�綍��np��ba�h'�/X;n�R**�)F�?7�ud�6���2�M�����j�Iɸ�fK1�}x7"�u��+L7�w�+5�U�\)�@+'Y�7�!\��s$s��
��C��
ً�[�Y�b�����/�,j}�+q�d��Lֹ]w���&���Ŧ	:�n�mNv�Źh��hV�
�.6a1$'d�n�Е����B�7ݷ��v�Q�e]e�h�����e��Ip�^��+d�@���f�Ks���؝�k�ɌųE_ر��c�z��I�6�>tj�jzy��|V����nRyHrox����b����0Z�f��ґ�CU�žU|}J�LR��qܰ��.�������UBU�ѭ�m+�����W��$�t�͗iMֱ�t$��3��}��u����5��
�RM]_#��Z�d���C�b(��Uo8����;vL�1aڙSMϸs��nu�yO2���(�|���*W5��+��7�o9����7!�l<���p��ٵ�zf궷b����j�2�TG%��!�d�J��ʈ+n�8D�C�KR�eW��=��j�V�Z����l��ɹ���z�tgpR���vwN:o�
И��1 l����z�}�1Z�f���y���U�\^����Q-TzX;	݃*|9����϶��1��h\�����ke�ἬxXС��s{�v��9��� F�.�-������n�@]���Z"���Q�kV��oQ�S���u��9j]���Qߙ��6q���:����%�7*�Cj>k�7�*Xu�Xu��\u���L�g,�wL�m�/.a�up{{Jv�$�^���M�
2�mϚ5��VGt�Ue5���80K&�R���qf��[}|��o�P���k��Ȍ4o�ËöN9i�-�s�r�a뒸b�e��u�5bfgb7-�Z���D�t�VUomUf��
���F����|�\�RS�WE�WJ�V���Z���grզ�[u9ʹ4Z��	۬j�k9=���ݙ��=| o��(p6��*�5Mkǅ�j�啺1���TJŘ:��ep�;��l�t'�}��P�U';E� �!6fQ��l���!w�<V�G͊؊�-��(��������U:�������Uh�>s\��L����h���ctұ]s�ViK��Dt�!��LU���R��NV�I�F��uR���wGmVs#�ڱV3�m�-�qtX��4��i�����k�u�T�:�W[e��hn��m��oͮخ�e
���r��䦦X�;FV����*��e���"���3]g)����E�X�W&[����q�U��X��ݰ��ʻ4^⩼���(Q��3��1p�'>���룂�k��:j��%d4X���������]Sǻ�yq�_�i�D�ݖ��J�KVk�B���l��(0u\I�7�J]Ѹ�$�Vs�[��T�7�&�?�@���{�f �v��ٖ����-3�⛘by��SI�dT�rԚ��G�O�D������:ڇk���{ۧ�7�����1�^�!�yP[�]�v�Z69�(���0,KreI�P_U�,�w�X��|S�>쮆�@/��tui�z#S_*�� p�>[ʠ��f�8�<�=�X_E���̠^[גƊ���1�e��:�or�;0�z�^�W�i�	�I�X���:�W(0^�$XA,_gu*���®nZ�yD�EF
q��PJ�آ�|�ví��)�%��-4B܊�=����%T9�	�F"�aыy�ZZ��sn��'��v��t�+�70�6	��	��ؤ��a��6	/v^V��h>��\�#��Zou���5j��}�7�m�B4Է:�xs�M�##��y��ܠ�%qt4�a��I����u�>{��]�"Ln�8�h 	*���n�� \����̨64K;���+O.`=�o)Y|1������+�|�Vn�����VX�q.*�TY�����&�c��̍k�>�.��`��n��a�r�]Ϩ0
��jޠ���+�Cb�\���1��g!V=���o;qʎ���-]�ڃ�!µwYJ��cg${G]��Jqܡ@�V�p��Z7�ʘ�=�ܑ�{��T�N8�i����3�BWt��W��>�]���-����w.�a
����W��x�%�����m%Y�N�݌=mp�r2d<\<TǨl��#��-�H݉Ymn}2wL�ٌ9	�-����w���s��WHŔ�td
��b�Wvڤ��*���˝GGr�Q�]v��]����k�×ʢ��1����C�'O�!�Y�,���c�v������M�BN������+^,�jn)6��Z9���w5��{�\.�M_	�q1+V�'O�Lu+�ꕛ���k�ګɬ� �OYHeҫ�-�٠a�Z���Vݙ�c����e
�aěns1����Tj���.<��V�O ���E�I���d�ۃ�$	V�.�b��Ԋz%�M��1�+�U�=���s(�͋���iQ(�I���VS�(K�9WLy#��"�[���;���S+R(t���{hFkNZ�!Gt��V�r��GAѕutf�@�|�H��ٜ�nM�n�cƖn�y%t
Fq��{N���v��y�#�Hwp��PA�)�w{�lm�9�-�4�b=��u�l�����ea��e�t��j�����utOq���q)r�gA)���YyGG�vX�V��w}�i]N?��L��Z�2ud���d�Y|�V4l��,-H'���H�4�>8���;��V�^f��ݖ��BM
"	����U�U�%#�Z}�� �Ϋ�o��r��^p5��U�$�CQP���쩡^,F�TB�V;�G�$����(���5�*�#��Y��W"RݪV~�D{ޏD{�>�m�)K�����hj�Z滤H*�e�UdZ�l��s�z޹��©�`���g$�V�$cͧ�L�:��D��0��o��_T�y�]����󧸀��`���I.�jִ�^�C��Υ�s���u�᠙$|�g�Bӯ:�AO��N
�󲺦{,JͰ��c5��"��<(�F�Ǜ�Ø�7g�s)suZ/f�qhBk�i��׼7w��&Nɑ*� &���eؕ��qU�j�V���u��H�OWV�g�s�s�s�QJ8�c�a�ᆳz���6�aQ�:�\��Vh�wbK2�;�o��}�y՜�I|��4ž�:C����l��wIVޞ2�'�nQw�0JfQ�^�c�}=2�f�yJ|����yݍ+��o�W Ę��j�1]�<��@���ެ�����++�!�E�9���<.�5س&�[Y>�oL�-37�a�'�1�]޽싶fV�ө�դ��|�WY�OY�[�ň�jTs�r�V��x7[����X�;'Sҥ4K��Jok�Y��-���f��2݄�����<K]��®� o*wWG�pIZ���_��R�`���$/�qs����uq�n��n����k�9�s�ǧHk�Დ���3U���ك��V Q^�G�Vӽ�s@��km���M�m��Z��jشǓu��b�o�
�F=��vm�mkڎ	 ��6��/Y�����s$���@K�òea�����JD�[r�sH�+g;��є3���W��r�Or1u���v�	�  �Z���Eb+R��ETU*Q-(�;�*�(�������X�""�TEUD1�kX� [V#Yb�Qb��\�eX"�Kh��EE"�jT�Qc�AEm
 �1EQ�UZ�J�kڋ6������Ң*�(��Ұm��*�,��W��T1�DC)`�Yl�j�(��YJ��X�AAb��7lb�`�UQq��h�"��ՋY*�R��K-KJ�wj��i�*ETP`��`�F���F����"F6�F�jV �%I`�҂�Z#e�Zʬ�U
����D��FV�1F�T��kQ�ر�V"mE
���ifYc���Z
�SV��Eb,Kh�T����ƍ�b�Pwh�+2�QUm���(��(�mQ�*����mq�*�-�����[U��*������,E�h���QjQDb�WiV9J�Q���Q�V�QUKj*Ŋ�l�mPiV*m�Q��Z4E��)6ܴb�*,[j�+(��EjX�)UAD��Mfb��`�J� E|� ����9�w����;E��.���s;HT�9���<6�Wtӳ�Wk�x�ޥnp
�{��,NAۚ֕��з��#�[�/X�l���׌�
�k��};�X�e
�� �g��	i�l��������5�!8�g�L[�0�b�vrmx��4D�6��;��.ޮ'�x��w����J5mgB�g���@u��v�&8�Y$���ע��$76m��P}��nX���Emֳ�;)��ͽ��.�q]��jtZg>��A!�(������*V��u2������ջ[����g�
b�:K	�x�1-C��(��'\a	�lŗ\k��=g���Ԏ@p�R;L!r��M��#��R�U�V�m�g��(>���Ss޾���o��9�:�ח����^�[�������EYj���zP�Eˡos%�kP��s�����sURu�􋶈�#պ�׹W��q�3��w���Z&�/peq]���,��A��G/��][Q8�x�}�2�I���xF��Dhֆ�ؾ,�Ǌ�ڭ���&h�˹w$h���4'.��åq8uӠ��B�aaj�z���ѐ={ՊCtɮAw0�Ui!z�q�w�֙IԼ�
5"��7���p�������l�`�:�+bC�K�J�u�H>Oy	R��,�����S/x��Y���,��3�Q�h>���@n�f&��k}�l�W=��
��wGL�򔲶�7���Z���ab� ��(3��>d�`��y�7�Avv�NP�y��:��z��t�*��������<�� =m�@y�T�����U��{�ێ���E{4z�-§�
�O�uζW:{�.L]J����pt����^����y����>|z���YҶ!<.�_'������H�'�Bh�-T��^��{�� �m�IS�W��%j����A�-����?NO�W�B���|J����ElU~P7�3��喢ek�o�������e�N��C*�� �c5�s<I�끹%�"��%�Û�����IW��[�v�μ� hP �8,����'O�sN`\�uS6��%�l�I>��f Y46��d�ma���*Qp><>��*�*#]ጳ���a\=es<;��74ʯ+n�u��s��E���C3Q��ċ�|�I�f�N�_�5q��\U�8�x� ]Gs�fr�m�Ug�㵴P�`��{���]K�W��R���f]�{N]����j�b���S��(����3�yh�#��Y��7;Uw<�D#�Ι'9��	v���$�}ٮ���Kx��j]X�׸)��Yv{�^�z�̸F�w�1�Q�
k�z�͠3 �g^�ueZL��o���ǻ8���J��'D��O^f�-ދ��U�L.�q��62�^T�}y&�α6$|��.[��l��ՁߝG@w��@��F}��[�.�+�z�:4mj�qE��{\YڷL�����)Y���Ѩ����V����UA<]�ٵ����rU��^���e�/���	;�UP�b˾�aN\(����F�\�|�&�i\,���Z�8��J��W��h+2��`6q�cX����R�������\Lc����sT9����9�Y��;\��s}�+����8�����Yt�,� ��%�4z"��=�3�q�[4�0���5>��}��X��V�%y|쑈�+J:��j|�� ��h�8�t�ۼ�|N�J{c)���*`�q������TfY�;��Տ��C��x�ZȈe9Z5�{�^�3w|g1n�;d��r�`�YY����C�=��CW�j^	�!�᎛�XS�3&�%>�(W�e��ڭ��d��/�9^q,.1��^/4�8�ފj�#�\�vz->��:���|��4*y�Cy=\Ϟ�Z������U�z�L{\��$�^ur��l��-������Vo:<�ws҅��u�n�J���o]��Kë��r���nf��9m�B�y���Z:4������[�(w0�%u�(&���2T���n,}0�\�lG�3��>e��}Հ���2�6}V�����Fx�J���ە����*S:/^|�"��>�z����*�d�S���)vg ���E�3p۵��
ܫ��m}����ڄ��N�ج�:S@E�=�/&��s��	ޡ�y��^��l�q�ֆ��;�-��s��q�����T��U�y��W�*�bc^���Yn� �Y/�vW���L�e��E�@������~�rh������)��o�<GO�udr��N4�W�u�wг�PO+4ڹ�KSqk�te!5����x��[�ѫ.�j�Ta���l���'Q�~5�r��6�n�X�IX�mW\^Y��P�o��Xc��OCȹ�[|}��8�r�g>�+Vv�k�PV0iw�ߵ�i{��[�[�<��X���:���)���=�J����G�������x7�������m��p���p,�iО1���]�Y����d$	[�Ձ�u��W��$k/��JE�k09v��Tw)=o@,-�>�5�@N��\0��W1���KzF�	�9�Xe]:��]왚%=��2�u��OE�4=��g��ׄo%�1��%wM���7��w����+`�ux���������r�,�k���/�x���h}N�z��G]�|���r�a߇��/�x	Ό�E3�"%����Z�U�w3YDm�1���uG�yeZ,O1�m�If.�ǹ˨�i��禋n坖+����"}���t�QfaR��V�g�z��㖝l�ty�k׉Ʉ`��ϣ��a�I#K��rή�/�JtC����3���/�L1d��m��u�/^x���]�ʽ��l�׼@4:�{\^�W��}������̂7��8�"#ȹ��m�lv��������+W:8<�����ί���Yq�ys,��(\�<z��HY�;��@�y}�[�T�s�&�kU=&=r�3P��gE`#V��46��k�~#�GhV���s:[�}����4���0��5�����Ocٺ��%�%̥�j#�N��#X�xp�M�微������K),��n�h㋆������#����z�� {A.k�;�=����7�|���O5.�gQD�*˭b�Ё�O{��יmO��{ ;����7�g�$���%q���*���5y������������um-�+ا5q����+B7�U�U�׷�ݾ�r��װ_����,�u�t�N99��Yx"�CB�76��-NI�Lo����L�Lo�c�r�Ϥ�n!� E�H<ǚ��y��r�.��:q"�����vX�1�����TwjϞ��/m�&!;LqEO�wz��>���i42;<�v����>����ky�)Ϸ�טjz��������c�3�8O�=�6%�M�آ��yy{X�}���W.]�/��{�W1o6�R��:*�)�LJ,	m¯'��+:R�au�ی��v�ʱ�v^�?^1�9�M?Ng%�R��}��6>��``�e�}�F��-�R�E��8D�fysuΨ����ر'�Qط~�V���(J�5;g5��\��v���ͤ�W��c9pV���V���ɯ��У�1V�v� %}yݣXn��_>����.��ꛯ=�mSۆ���S��L�����ڵ�wl�>��GJ�"���ݹ�5��V:��>�nx]Kyv��p�u��"�_�pmY�:�v6=Ρ��V��z���{�+d�v����ׁ�
ܫ�k���8�ɴ�=�q6|+FU>q^����4[C�U�B��_9���L�.h�y?�	�V�h̝�`ا��n�[k�b	ʼ#�5}��I^�Ѽ)��<�]�e��s�zõW� 2��ӣ�ٌ�;z^l��|	ʽ�����^�Bw�g,d��+\ޢZ�M��踅e�;���Pt7M�\��ZNs�rŚRWN;�5	����}��Rg��az1c��]���9K��%~��=��I�1��o�7�ަ�Ҵe��J�}X������Z������$���O�q;�ܑ��_�������5NW�מ|�/|�<�j��8�FXx�зx����<!�Xz�m����N����QK�S�l�yo�-'ȌzT�\��g�c�h���ո�&oU�V�t���ٔ7�ޫ�À��x�m�(�AO�=�h��>�E�;���r8e��u�����{hdGn�E��;����}\���]l�>v�y4�rx��U-ų'�ǽ���<y��,h�]�n�R掗�Jh]\�����ə�K�V�Z�o��̓S�Z}>e �lx*'�������z�w(�����L�L��;�{�:Ɔ��F��x�����0O����WD�s[rC�������屿b�|�ϝ��Iyi8�B�U�������{|w`�e۾�Q�˄��]�y;J�������_2Ix4[�!r���p�:�7�k��w�x��>�N�]d���q}�.��R.���a�j%g.Z5MN�sy��4';^��o(�c��k�V�T쭦���t��t�]�п|J]�zP~cK<<�h{.Lژ��M�:���j���L�.Nz$)/q�u�r3Bq�suX_(�5Ѕ�ӕagr\e���θ��1�9���f�����/wNEԼ�{��sӱ(&m]�U.�KCwr����u�4�þh}��w|�8/i���*�*5hU�����D��JI3	hoJ�A��|��u�W<G�
Oh�'���轚a��.S�����q�S�s�ss|���$�נ�p�W/RtK[IbqPs.�%�Z�?hC�$��)�nM�n��rLYA*�~�Y���1t�+�ĝay)�k��M�­��q���4�l�T^Q�Z����b޿/��l�xP�[�l)/��X����1�%��to��3��>Qs��C�Ղ�XS���^3�]c�ZPώ�Lu��������A��n�z#	�wOc�v�����~}���u�����j_S�{�^�xz�WL͘��7���܌���?����#A���\�rz��5Y�a��h%���9�գ���ߗy��[w<�����}|��j�Kg�`�fi�O�2wS�۹��.]0_f�3y���/]�dh��x!��t�3h͙�W3���X����"�����)S��Y��)��.�R�ʼ�Fv��+VY�����ݼ��:���Uw�<[t[�Ք�L�-���g�a3E�<�:�jn05�ɺوV9c��d���*��z��%�-�gk�	'n\����E�ޥoteVs��ۃ�k�nm��c��x`��Y��4z���7K�u%S��ci��u�sR�2����գ�}8��R=Fy�$�["������ڗn�/cφK~�2T	�t�(*~u���ږ�n��u���7ԥ��g����^_rb�K��1ʬ޺�s�|��6U���0|��Q��~�S�{e&�j����yɭJ܎v������k��y[q�w�ٖ��\@מoA����)N��8���gCp{m�Zr������{p7��{2l��=��ݵ��2�"��W�Ԫ�n��_�9�����y�=}7
{��|�e?jޟ>���cr����>>	�����\��l34Y���n�Ŧ���:n�u�n};��4��o1y㷁��k�7�Q�N��zp�sR��A�.�Tr���R��c޺Ӛ������Hڻ`T��apLu˅Ս幻��֥ֈ�"` ����9�0�){K~��ڏ��{�O�>&�;kn��J�C3fhK���`n<�%�.�e�=��fs�TS��_d��' ^wW������[K/��,�ws�-p�YY�i�=��th41���Up6��M���t���S�7z�X�VED��1����B��&"t�l�{1
��B�WE�Dr��2��!��nL��O�{Jna�H	XEZ���)���P] cڠ���)/�m�b�!.67�r�=�v�V9���
aȪ�]��dDQ7�0�T"���拌K[4�LPM��pخ�����X$
*�]`�\6X=ӆf+�6\��г>r��i޾h��i�&�����{�ũ;���2�':�@Ugu�N�T8��u����JI�d��wW��ǱWD��2��[٭rj͋�^�V>�1��H��'>�%�\�/kX���CX4�zv[���ݹ�5tBj�卓A��(�Іʐp�獮^\���z�^��Ҝ�ˍNj�LB
cm�(�S��:�F��%9Y{yz�����9f��OA4�,'PMh�'c���l=�W�.���Yu�*Q�L���ϡd�Hv������H7ٶ�x�9E_8�m�Gr7Cy��DZ/&)��-���*	_A,��Ը[Χ �Uճ5��:���X/�;1�,�o��v��w��ҹ�i�:znnt���	*�Ս�]�����ՠ����ϕ�o ��������t�K�q�����*Xp���b
�Z5����a�*�LO�Cj�pYeC�&�2�fc��b������ӂʪ����O�eIf����l�m�S�A���b�w�n7�b��V�B�)J&}�^ o2&����Y ���lT�X��}d�PRL�@�f_LL��ӽsq������*�j?�j*�

T�.����F�amj����`�ҧQ%����a�ɼ����h�VBGB�P�u�.�̭,��¶��+��I�J���n���o<vM�ܢxd�-'�56f�6��X�g���:^D]����,H4_
�k0��Y'Ҳ�]�!��װ��f����
��{0�$�N�V�R��%��@�n+��2�T�]�G���;4��P��r�k���;�)�Lý]ԓ�3YQS;�/:4�;�o1�J�J����VE�`��{�>����kj1r P�(K={R�Ӓ���vK��ɬ�W����Ϛ{���,|;.�v��	��Q;O��I�*V�ch����!�;�yM��KF*Ҭ��h�����ޜ�Q�o�
I��t˼6�6եD����7.vr����o�#���T��U,���W���C&\�WsBR[�cUi�V�+����X�����都����4���.ٚ�r�.��1��ϭ	�wksZ|>>���޿>�����}��E*UPD���DJ�V�b�A`����TV(�
:�Q�2�h�Ė֥V5��q��(*��l����b�UF�Q\����,c�Ҷʪ�FV�+QQEA�2�X����6ն�TFڊ+j�Tb ��M7A��5Jň�DEUU
V�Q���A�,�k��RV��b���Xŕ�ȱB��(*��`�R���TEdPUF,LJ*�rؕ���,D�1V*�b�Yb�X�b��QE��%�����Jʪ���+XV1R����QD��J1M\�10b��	c-�e�T*��%��mJ�e��b�.`(�Y0Dm�+PV�UQF�%`�`�j1DE��D������
�*&-b�"8�\j5��"�Qb�ZV"��Nd��bQdQ��.�b����F
��cmU\�r��2(�mE��j(�ƴEJ�جX���Db ���U�"iUE�+i��"*,DU#b��1j��X�����|����g9sgwB��)6�Na*�Ǯ&��&P�ӽ�,����qɵ���X��B�qq림�F>��{]�h\�Ov�ٔ�A�D�\��̎��!�k�����ԗkTm��x�U�h��������Iǀ}��Ш��c���s�ݓKnd��/3sos9*�2��p�6ل�}��{�S�z�HR�|h�vLdŶ
��Ag��m%�:'�ZfS�n�O0��r��s���GR�2pl���7�j'3������[_�1�����rN��Z�s��(�Z�����:�3e_���T����ko�E�%{����"�uXdɠ��W�����n��⎑	� H. â��ޤ*40���ٓ|�|�m��6���b��f
���F/�ژ�S�-���,[���I��ns�������ϩ��j��_WP�UJ��2���C��z��׶���݂�x��g���X��"�1.�e/�V�a�PЇ���n{�JA�{�o�O����?#&�z�n�M�jNڿ��/�X�Uu�m���nS����H|m\�뫖�Z/қa���;����t.�Xz뤕i�0_:��(���k��禩�43���ۃ(����x=(�Κk���;0r�B��E��db�����r�p6�C�&�F.ת�Q}��ݞO�3��>�Ō[ ��g�
8W)ζ�����/�w�����Ŧ��v�_w�{����Ό�[�)��痛�w�Tڝ�ϜL�y�{Ֆ���*�c�V�>�B�j�]��zE|פ�:�x��>��Lq�{��ψ���¨<=2��+��4���loWo��؞���w�n�G
�>���[�UD^�\�[v}���ű��f�z�tqj:��ף�r\d
��d�;���ѕ��j3kj2(>1~���d���M���޼���|�ݑ9�)�"���}��_!=��2�}�N��7�:9��W��\!ZW�h/9k�M޼��:�)t�h&�x!uz|�0��K��U��u�{�o���U��o�u���,�H�x���zO�Xy-=��Ca�����e}ֵ��<�7k�`k�.&�x(W���]b���N�!�,�s�״5����f)ܶ�.%��N���C�)���O+��ս(�`͊��g��u^�K7T����|ied��m���>���{etf�W�2��]%<�/O��(k��^9UZ�_�Y��-A�jb���v�Ub��aB��,�}�Ŭ0[�w�W����B�ޝT��SpG0�M�Շ�o�>:���^̸��W��`J�M�e���*`�����8w��<�w���L��������Jg����V^�6�~FMژ;-J�0{-�NuR���;���bV�ρ5x�Lk2�f3EQ<�\����4lþ�M�s��3ۯ'^�ى�;��zN5�iCޙW���%_�œ�@�Jkٞ��|�/�7��
��qū<ƴ�m.y�fa��+��sy��Їz)��wdZz�1��q�Y�{�.�_e�g��^�\>k�}�8��p�j�t+� ���w��ߦS���M�(�n4�	�=�5[r�nk0�Z�oy�+ı݅4&TpS>���Z�z�'+��ucy�2�bCk,O.G��#A�yla�YZ�YF�S�n���e��� B�x	{����n��^ŸE:�^����i)oVRET�;Ԃ�Ϣc��Am�l��f�k^�J���v&-��}���ɂ��AcUl�Y҃ҩ|�2$
�#=�3�_U-�hd�?͙����{��_im��{]LxS��f�&���nPh_Ľ��(�[�G�����S&���8yp�8܁uN�T�&.��LFF�m�1���ͤ\�]=O>��j��%�zeI�c�٢�6��M���XW��6AZ��M~Y�\�L�z��܈@I*���w����X��}-����[q�l��匽g:����)���N��R3�M'��'O�u/hi�N��d�0�x�[}��3d��t��.��ԇ�p���>P�}�J���r�8ü�I�XN�5�=aS�Mj����mo�	�!�!�xɤ>a�,8��h���I�
�֮�|�W�7����~��C�|�i;�2x�^���O�1�l�0�P+�9d�a��,6�I9����Y4jÉ%f��i�9AgY4�$��}����]�t�g�����~���׾w�����x��:}�>a1%Ms!�d�M��0<E����xɖ���Hu�k���0�d�}b�I�	͓2�x�̛��C���~���ͼvo��}�v���}(@}�	�=_���Τ�;`~CL�E�>�J���w!�I1��;��'���� xɖ���@Y+&}���I�M�E��'�8�3�b���]�+�;��ԛ}�1����/���+�����Bt�g�i���o��'�N��/�s	�Mw܇۲M3g{��'�d6w�~`~a�4��� Va���P~��?2j����4?��Vө�5��4Wf��o����$�hQ��(Y�Úi�?q����.>���jڗ.բeU[�r^�͇t5ȫ2��d��i�O��f��6�vw�v�	h&汎�ay2�7X��P�뷳���UW��)O'^?9�o,&0?��'Y�M���'�>d�<�'Y'�<�I�u	���4��,�?~�@~Iĝj~9Bz���j�4����X~}By�����k�߼盽9��O�����@�$���+&�c�e'���l�<5B~CL����$�y����5��'Y:�'�Rz��ZsV�N�ݜͫ?p�o��z�xϥm|>��~/���'�������=f�}�,?2O=��QI�?$6eXi��uY�i�F�I�M���XO�Rq������w��'ز�;d�����o��_��Om;�|ԇg�,��$���'�>g�4�þ�ROY�7�|а��|�p�4��e��i��Xl��N�����=I�w���{��n��}od��'�Y?$��<�A`u�����Hq��o�����<�dY���oO���|�=NsYO��!���4��,6=�~����,���DOO�g��_S�����$� oZ�R}l���N��Ć����M�O��	���Y�'�8�����&3��s	=B��{��XN�.���Oܥ���sey7�U}�>���q�h�� zɩ���'̛�a6��q���N�=?s`q��<=�C�+	�o����N�	�d�u���=�3����oy�w�zI�+yEI��OQd2ӌ��9l��d�ِ�`_Ԛz�|���O���'Y�)�I��&�w!�
�=s�?^����L�+��?%�ݾ�O����:P�����<d�S���VL�wI�5�,���?$��6['a��~�N04o�&��N!�!�~d�{źln�)�?���>��i�c���V�V{��x�6{�u�~f�<7̇Rm�f�s$8�P�h��u'���a�����Ld�Ԛ�������%[Y�y���0�DnQ�h,S�Y׫��=���V�&�l��m\��Wݥ'�q
��I���զJ�����b��j�{ȩ���[c:&�<e�7�O��2U[��(��븪f��3ˆa.=//b�����:�gY�r��T������N�l�r>����R�WÐ��2i?�_��&!Y����	�r�!�O!��!ԟ�1o��bCA��N0���0�ve���">�v�%�T0��[G���X��ӶO�:�x���10񀲰8����$�
͆s��N���z��,�y�Y<d�a����b�(�_~}�ŋ��]���Y��ߒʅ�yW���ΊO�$��d��:�f��u�c5�rM��!�~��:�hu���a
��8���E�����M&�O�[!���x���?w]�>߹�w��Ϸ��X�O7��zɲ{E&�P�Mɖl��,8�x��k��O��&�c'Yԛ���|�l�G�sRJ����eWY�����=�������S����o�l6�g�d��g��Bb�<g�M0�{�	���<��I��k$�Bl�}I�N*�Y6���

v�M���n��~\���j?���UW����wI4�ϻ�䞿2O�i4��y�+������a����?$�g���i�[�N�O�o�d�K���S�����&���Ԏl��O����Y1'8���ڰ��q;��9�	��C�?��s�=`z���w�,=d�����l1����Rm��P���'�Ǿyn~�����{��I>d���~E$ח�OY;l���`q��Y0:��?'�'��p8���'���nI�<5b��Oɨw�,�ġ�֌��>Y��r���	���W��ﺾ���H|�L���,�ԛ���I>}?Y8��`h��4O�:�׬�vC������I��z�1���5$�1<��������6�K������Ns��+����?$6e�$�'��s)R|ɩ�ట o�O��}哩6�����4�O9d>`q���>d�{�<��쥘��w�$:�����o@f,���� ̸���{M^�Y�s�$����s�@c�E�n,����R�ƃ��3���g�?��	z9��x��эѭ\�(Vo��@�v�i޴	�,�
�ڈ+Yk�j��{i��n�:RE���/){�����K_�>|۔������2y�+�C�6�ͻ�}��a�{�8�8�O�B~���=d�RT�q��y�RO�6r����g�$����2�?3���u������o�~��·�*I����2m�Rr�:��LC���$�a���(��CG,Rz�%�䟙;l�-�$ѿ�L'3���'���<m>���ą<����'k��% z�����_}��Ώ=�C��ל揘3Ho�'m��ù�:����(�N3������/?2}l���:�n�<�N����>�7��?ߞ��t��s��1���D����I�kܟ2N3���r3�$�=��m��@�ré4Ɋ��	�+'{E�>;E��a7�_����W����o�9�}�Jɉ1���R|�����B|��������C��!����3�ԓ�=�C��w���'��3�I�&"�5̐�%a�zr��r�{�����ߟ}�ޏ,�ĝK��wSYԕ��Z�q���o��8�~A}`c!�,�Ri�^�O���9��)'Sr�!�OHn�g��s×����4��޾^����>d�C��C�B�RN�l����'7�ԕ�ɩ��%fk̓l>Hu�C��g{����M��:�T�;��9�q��{������������^�h�M=��8�Ʋ����xɖ�G��@�4�~q$�'Ȥ��'ܡ6�5}�P�$�l�L�	��~CL�C�;��.����=޼�����������2~W�~�J��v{C�XO��{���d6w��Ğ:a�{�T�!���+	�N"������ڡ<C�My�ē�z�����w���k���o��~�W�q�a:~��i��,���?$�'Q��	����w�n�4����|���<`x��L?w�Y*O5���'�1�Rx�̚a���gx^��]Ȯ \�(<���j��awۻN���ɷQ��畭R��W���zmW�촃�i�T�n�3�;�\�.#0��s�T ���#�H#�k(i�<律�m2���4��8cęP�w'�r���� �H\��^+�+����Z������� �����?o�!����(x�<C7���)'��I�,�μ�=I�N�x}̄����;�_O����<Ŏ�~ÌRx�{dw��+��%��d��,�U���}'����;����l������dѿrq��&�5�q�^~���`l����d姓��O�O�g�OX}߰8��4}�3�s���cӂ�w������}�	�<�'ϼ�ɦx��=C6�Y���i�F��$�&�ܓ���;5�$�'-�ğ0�ާ��$>Hu�6g����x�������o���6�e|?�����u�d���d��ɮ�$��k����ٖ��Oa����:ɣ|�a>d�,��I���'9lg��;j������7_d��:�ҥ�~�	�Sgu���O�:����|�Y1�y�a8��I�{3�@�"�d�&�aᔇ�8ɭ�Z�|��s�9�<�~}�}�;�?�ҍ|>t??}���q������O����P��~g��0�'�$�Y1�O�ڄ��!�X���h�,��Be��$�RW՟����A?��D��s�� u�����O�5�d6��u1�Ԛz��~�N����<������u�2x� w�N��LC����J�w"���}���ܺ���2��0�8�~Q�_�M"��o�2v�l-�Rm~��H~߹�XN&0�&��'S�s'Y'�|�g;���'��ɦ���̓�m�gy�m��޻�}�����i*�̕�5�,��I_�?2}l�N�=I��s�$�s�g�a�C�C�=d�l��8�|é���m'����9��z��,��~�w��uw�W�gǬ��b,ϨN!Y;�9d�aÖ)=k	�MdXT��Z��ԛv_��C[���M!�
d���|��C�<����f��ՍS�j<A�7!�v�l�hZ�N�`�k�l�g�]��%qT1���3�Q��9�xLό��Ϥ���h9�8��]2���=:c��[���Q�L�}N�Я��';�r!�޶��"m<��z���J]�q�w��w]O�!1��#�S"��F������������x����m�2�|+oSy{Q�sA�OȰ8��6�����ayG,��4��sٙԕ�&0�IY��2M��!��N�N�y���y�o��cb���y�PR�+�����6�U'Ss�����܇�u6�2x�gy�P<d�C_w$:Ɍ4g3�XN�|ņ'�'=��=C�~dy���~;�y�5�7��}�C&3���6��&��<a�N����*i��]��$�:��rT����Oք�;�<dա���������N�o��y�}�}��w�י�O~����衦i'�<N���3���̇O�6y�hq	��x��8�&�}����:����ĝN�a���L�w�|����yO0�4��?w���ߥs��t��3�o}> ���~̹W@}u�h�I�?2m�_5B~C�My�N�O�6y����s��&�8�'�P6��:��(O�N��!��&��������wn��R?�,A��pNR�?}N��~���S�R���<t�����$��}E�L6��Rx�̛g�Oɦ��ta>I�Y8��7�	�N���T� q���s�s;��M���<��~��~�o��2|Ξ�ǌ'�7�ra�z�x�X��4�ϻ���I�g~�Rm�
��1�l��x�2~�0Y'�5��E����h�~������\UQkk�k��	��|�+︑�fHq��s,��$����C�q�$�;�u$���s��a�	�l���C�Cya�d���N�͚�}�}�=�~~���~��}�I�N��ԟ��|���N�|�Y:ɴ�~��!�Y�������?���2b;����1�s�ೌ���5�d���i��=�{���f�x�ۮ��>���Rc'��锇�:�[�i$��'��>2u��$<��Ěz�r�XN����2xÌ����&?J�ݏ�t�����[-�r��[�-`����M�K�P�v�\є�umr����FP�)�L����.��oN����Gu�Eghf��
��Ъ<�"<5�,���q�"�I�ފ���޾j��F=�Z�3δ��9�uqfB�ѪT�X!kM���;;�������_��A�?{�
a8��y� z�Mϒz��,72��2kkRO�6gp�~a8�Փ�N�8���g����u�a�����T �5���i���ߵ�_���m�����m$��y�Y'��,�E��ӌ��;l���q�����N073�&ޤ�O&��!�=I����}���K����A�j	�������Oa�
�t�����O���I�6Ɉ���	�J���E�qܢ��8��'�I���8��'�'�|��Ҁ���g3��c|������6��vk�jq��>g��6�&����C�4�����M�b,�k�ԇY*���IԚ9E��I+��c�'���_�>�O�?�x�򹮏��ۯ��*���,�L?!�,�Y�M���u�|�e������CL�*C}�C�?2b,��0�RT�3�Y'|�M?����^�,������oB�O���C��VN0:�3Y��'�8�x!�=I�8�g�a��M��d�!Y�>惨�Lz��M���w���L�v��th��-U��T��d�7[��}P�>L�=(x�v���~I��2d��oܓl8�o�<N�6�Xy��B��N#���$Y:��"�:�hzɻd��0	��w�����a�� m��O<����h���>��O�N�a4�<�̇O�o��gM�����:Τ�r��`u}�J�������."�\���/����ʀ��h���Cha�L?{܀�+�s<q	����~d�'���3��<�''�7<�I�:���}I�N*���{��f{�<�����ﲇޯ����>� 4�>�st�Hnw��~}d<�0�!�Hw�`T6���VO�bd�i3c&�gY'�v}�w�5�P��!&�]���l�b��k�*7�v�L�p�ob�t�:���ˁr#J��1f�k��y�wI����4∘^}�Wn�BpjB��+^�y�"3n�Vr]�C������u*ʥ�C�ի�e�(D�)��}�ZJV�<�A AA�b��嫌�o�⭗)�&:p�6��34��Ђ�vdʕcX����Yd8s%�%_�9�֞Lcb�Ƿ�icO���R��-:79�d(ܩ��7�nj�B0Pq8���a�t]�Æ=�2�����ب����'駚���K��&�31�@��۟dPc���S��$x�����c�oW1Jp��������ɱ��^��X;v*��}�2g�f�.��9u*��k��{���x�L�8�UΨcI���Ⱦ��\fn�e��՛��R�y���\��ݜrs܄�᫹s��]=�_uoeC�����'*[��Zp}��2^����,��1�)�U��%������`R\�&��/���ݒ�4	������%0�Ck)[�A䈫�G�"�BAٻ�^�[{.� ���:*J9F;�"�U�%og3CɌ�B*V]N�HuD���+�x�㙷�+2��YF��+�@)36$�:�z�l�� &�]-�T"��s��-�7��4�ӡ��j�XW��pv����>��6�<��R�u yce:�Efk�W+����r&����u��n�D��`uC*�aR�}h$��yۏ1�t��kxv7X/u�`�G,a�&a�[���L�u�;�`V��Q@�1�+b��U7�,�"��0d2�+1��U�(��kf=4�ݫ�c�Fi$
��k�F��: j������s'���vȘ��J_�a�Y��2(Z"�{IN3��t�`��T�0���m�-]�U�6��ZZ��a����5u֒��Ա�Ĕ��B���=��j�F����d�LRt����;`��B4�^��ٺ�\bf
��b�I�,LYP8�_�}Xu���������)ئ�,ͫ	���h�R +W�F��t�ێ+�5Z��#3�L��*}�ۀ�yЋ�
X�`\�[w���9���Y��%ˑr ^-[��]}����%�\30w<���:��Nv,��f�WX3�%�V��C�Q��Jc� :�(F��"ổ��t�BZ͙(�m9OY�7]#Ə+�t��}ۗ���R
�~B����"���V��vɲ17P&7]�ժ\�a�\�n��E��s�2�+��(U����䡮�>��T'���%I����_ !�ͷ{B��*TMQ����+�%qN�J��G��l��+���釟Sư�qF��8�s�1y���1&�Q�����Z��I���AIf�X_]`����l0]L�ɺ{�.O }�A��v�v�.�k�[���C��Ͻ~30�EKk���*~j�F1��Fm�T�*��AQ\@�%�M�T�ED�+�(�PADb����PW)b"��5��-,QE���PH��łTQ����ň��U\�TDX�UV%�H��dUTF���Z��nZDF-J��2UUM%U��0��UDUF#��`��(�
�ŌDD���""�Y��A\h2�U��DV( Ȣ,AQ�jʂ#�"6�+*�EVF"1Em�e��QUYZ1X�Qt�jB�EPDT��,�GT�����-J��U�**�QF"����t�\J���c�X��,X(ZQAV�JEb�(��U�E�*���Ԣ�@eJ�VKh�J*J#�b̶-lTbF*�ŶU�Ԙ�(�{����������}羱y��|pvt��=���+u�Ƨ1ҷn�Iw�C�4�&�o-̍F�d���3��5�������u}s^�߿~���������'�OQd���4OY:��OƬ'�Nv��XN0�������}���z�!�X~d�{;�&�c����4�Y�3�������a���=��w繯;��4�������߸O�I<$�'m����'�IƧ��Hq���9����'�<�p8���'����~~B�z/���_}���2�Ј`���~؟_*�o����E�l���~a��g����&��$�&���:ԓ�a�Ì[G��|�������`u;X*����u��6/��ӕ�ޯ� �R]���ǽ���/z;��WdO�{�o���Pڹ���ة)2�>y�?S��=W |���=B��R�|_SCݓW�A�,.(�EV�9��mn�[�OSn����4]�HW5��##QHU�t��g}�V�9۵=�e.kq�M��a�O�]-�:�=�T�7M�];�ϖ	�.\�^H^�1�����RR!�O����kp�1b��{G�3�J�X]^�7�R��U��)�2a�$��i��ŵo�=O��
c������+���C�]�N�pL�\yV3&}�w.���J�c�>Ě����ͫ�;n@�8���#��I<�Uy�]�عWI�"���u�kS��3���|E^76���]��u>�t�L'A�L��;��	�=A,�뛫	��f^���.c�o��ڎ�lq����������Z���V�{��<�G�}EWQ��i�3��ZZ�~|b3E9�7@5�^Vc�z��J2�nT�F��������VX�f�Nz�36wfmVn�|SN}�T���ޥ�`���p'Y�б=�)�������Z�9>�׷0^v�9�s�e���w%E��pْ6j�mDÔ�2�Q�N��u\A�S踤y������+}ٻ��Qv���K5�[�v��,�^�ϯ֤�lVy����4�N{c�/����<R���>��+z�z=�Ro�Z�;ɗ�&6�RC�Տ>�����̵��a��v����};���X�n�y����i��(��ڏ��xߝ�S&����\��?3�S�!���ߛ@��`��.:�����}���o��R��a��1�y=e�yǪ��:�5g2�V�E�ҙ�چ�q��Ľ����^A1�մ;ֻ(0�J�ჹƭ�J����f���pvv�����}gѬ�$�^{܂W�}�t�:Y�z��
���=AVY�#�}iʳ����1��%������w�l�uu�+5�z1��\�����gMz��9v���^����\�\�sݛs)|�+RDf}�ө�W����tI��~���0OK����N����v9�Z��}�3�sݟE���τ<�:M�,iu)��|z+�2���N�<��5��Ac����pa��^��|�m�n�ყ�-�H-��4���[ԅ{���_{�!��,V��=o#^��&��_�&T��5�[�e�|/�Aڅ�5�7�z�p�ݧ�<Z��\Y�I�si�&��
8}t��ʋE���-Xjxn.�߷���v�6(��&������PGXk`���6�U��g��T}}�T�����O��'���w�E�-�r�x�z;�w�͌>�Ks�Nj=�NR<��͜�V�^�x����gV���`�`�u�]��x�u�ݺz��a�[��;�>G1������Uz��5�Q����.N�ŝ`���B��t{�X�e�P3X�PUF	��{�q��CR�n���㝕�TU53}$�5t�W�	H0�p��RY��&,�j�kZ=����v*�uk�Z�Df�S�"�qհ�)l��
��廹}[�9��xy\�Tfn�#&�!������w����}N�Wj���G0��Q�5:���j�9E�UQ}ZV�6�㊂�d��KsM�^WBp����n��p�ݵ�l�,-����o�fWz]8�T�1��G֟�k��}X�&Gb_�Ϝ�ӑ�Ӷp$-vy����Nкׂ������1��;� :����/�D5<*�>y5SS���u��S��eO�����]|�\�_)�wr����ʝ���H�nS�3J�\�D^.���d<>�U��qv���6:ɼ�Vߛ�b�.s�'�٪��xr!	%_ޟ;chR�����xM�L�Bh�)g��f{#�g���E͝�k$��nY}m��.&6�z{Q�Щ���iΌm��YTݣ����C��(P����V㭊!.��[Y��}�z����L����^�/zu"��������l������q�Oh.n���IA��2�����:򺹩R\]A*�S}Ӏ�دbU��G%�뤞�]v�����!+nDƋD(���k'oW��u����P�����_P!��)��I��`:�=�p[;�bM�ǀ\�լC�u���A{;�U}���ө��E���܁��ͅ��,�;b@��{�r	{Uy2Or��n>���BE�Vj����J�ׄ���2&���ϵ�}b�s�o��'�|�ds����HGY���\��O/%����Hy/�V���:��X�C�O6��ņ;���@�6TIWƕzi��W(��o�2V��<��c��Z�`k�|�[�{ہ���H7Ӆ���lz�L�o���n����G����^l*���������5&��l^�����k�٢�`���밠��v�7X�d؆yۥό�WKQ�º+�\,ݛ�A�v;Ȼ�[<`���"v1��3�L�陌�P�9y�9=Io��B9Z��NN���ǝ�}O���#����}��Ǩ��[��/4�/%�٥���FD�LX�؜`��t;�j���g�L47�y[��k;K��g��U�TvE�sY����fW��iL@4��'�JJ_eh�K�TCF��-��˥^{�V�*��N���y��*���Śk;4�Z��3�Ӷ-PںGje[	XxmL��?i`�cD�8�#��t������f��"��m�S�f�����y�c�W�I0�
�~���_��Xޖ&Z�1d���s��»�B���~�k���|�/H�y�N"����=��}��e,�}��}���!z�=ھ��;}�_l�qI/>9��.T9=ѱ-m����X`���ڗV��=����g=��"C$�L�k���2b��oO_5�.!�y����o/�D���b�9^�ֻ����o�=}Ub9��V#�5}!g�{��Ee���;�<4\�حxo.��\+_�m@����(07R��ĝ�B:̴6
#�������ݹ;w���'����p�t\-M���7�T��n란q����FŴ�t��׽Xi���d�)dc��)|9�����8�-��-�-��<{և���6�|���I�e�󔼵��נ�[ޠ���������+ �1X�VE�����9$�8��t�֖��Ek�*w��+Jgu�zgX�����r2���!U�H���]�t5%3�=CD�m��glgWz�_N�A����Z:���3��,�J�8;-���}_UU2fZ��:^Ξ�y~���{yat�����/��jA�n��G0�+�s�{^�������6iQ��c������a1�
���,{P[�~�Vo�t��������c�ӭ��f��S��sK�]��(
8�v�*�b.2Xۍ��	��]Sao�9��\9�`����bKO���9=�~�%k�������\��E�=ٯ*�9�rK3y;^����i�w���]@��c��+�ԫ�_W;+Lyٱs۝3���y}�.����c��;
��H���GT8�3�E��|�xxr���fl�[<����:�}��s�!m���:0:�=�|��ivaH�9s\���W\����;��nW�9^,[\4v����ڻ�w[��{�&�A�F4��U��q�&��:�W�����>lZOs��Wg�>��ݭ[�A]�5�� v��E��;�W����=��ʹ#m?�nb9���b.���(���Bj�b�5��yOj��d��W+NgZXܩ�F#�.�s�r�@k]U��>������DP=ygp�jpR$��эv�Ϋ�0K!�:��q��/kg1�\:��D��C��?�|��">����Z�]��̀�>ۖ1Sy�z6hv�7�[�d�I.���=3p����Ǐ[tS��
�'��dQe�����%�7���PMߤ�	�B{ꏣR�bKIv)x��
�5X��M7�=��Q�C-wr���{�������s[T�z,��B�zOS���X�Ү��;�'+h@ӎ��w�ON�+ͷ���Z���� JR�5y��T�`���c֣�)k�T���{q�#��7�\��K\L$N��]�l���㭳���p�λG���&L��q���񮥘rd����ZǮ������A̭�K�]�J��Ӂ��l :��H� #�u�F}�.��9ߛC~��q� ����^�Q�sG���Y!�X"��]4J�{Ӳ���z��?��4OҐ�k�*}ާ~y�1������+ٛ{L����]V�Q����){M�WGs!Q�k�N��G^�e�=�����)��u��+{(��X�]��ٍfũ�cP�Wf���վݾ�J�)�)6�gԿW�U_}^�T��2��r+�_?v;�JNV�m�u���ch��No<��,�b*5k�v�0�%Q�'���QX��|Z�%��q[� ��L.X5�rTW}���fu.�c9S������H2`f/s�r���zvt{4�	����k�'���u�|mzD<�o�y�FD�a��y��@
�;��OS]\j�`����s��7��ײ//:�����!��~`[I��%���[MM�8�^k�B���j]��g
'#��T�{��XyC�\;q� <�6���X{�ԝ����[xM�;<�^L'��@|瑥i>⟵��vyin���޺��c䮱�W���$����j{ب��𗔙�����M���9X�6`��	����ݼ�7�z���<�ݧr���fV,�t�{�(�aVw�n:�p��9���됪�V\�1dS�wD#-�7��STXv��~��n���U?~T	�iZ�#��`���[ƷG��s�(s�4$�%���o�$�̣ٓ�0��v��YK�v��X�)s'�vH�r :|��N`���p�|��z����|>f�~孚���a~b�^L�ap�9��1����${BV[��U�'���nߠ��6�M	���/�B�����]+��j�=�_EXh?S��yG��psr9!瓾���}V��v8]=�O>�{���X�վy1os����}�W�od�˚g����`�]�F��\�τY�N���ft�����f}o�c�mR��|l����E��W�ϸ���-�JW,�W��	Y<�R����������=W�v��Ѝ9��uc��m�u;�і��Tϡ�w/�Ԫ;k�nm���\������ku���x������1�k��ؽ�c�{b��^/~��:~ ���\7[�7*� �:�;x���sԖR�����h?R�_b�Ն���e�h�9�;�:.|ܪq���b���zT��*�Щ�]�sM`+ �r�Yv���f,�s΢9qM��8#DU�&��6�m��GO�{9v[e>�7�j���]�4�#�~{{,��N��<+?)�����ł��tѵZX�u�_1K���ڌ�:�Ko���|�4)Pf���ʱ+�h�83A/+l�Lvĸ�h=;jY�a�35d���b��R'�R�5���⌧k��''��fN8:Z�!|Y�V��m��1v��#����4̮��t���z�t+�e�-���*�S���Z������l��
��2�onX���շ�Edf��Et�i�y���RϏw`�B���F ���\*�=�Ej���U5���k��q��;���z�ȱY6�2Mm�̈���eG���r�9Q����$J�:n�N�C/A5�{/h�\2k���d�c%9'�:۽µ����f�[��;}�T�q7����7�&����b�gl�0�s;��r��}wh�*�[zV���Gk��I��jp�$��w]��YP��\;l3\	"�G�+�9|�r�OU���cGv*�V��h��%඄��%��A\$��x�[��Bܑr�=̪����r�'d)�x=X��tۼ.����s�� f���rUh�Gycǋ1�wU;C����Sՙ�v���˙*��_j�\�f�*�U:4o���t��ױm.Į!]������-5t��ۢe5�7��sWU�m-����\��v�{�3��"&	�+U�E\��d�S7>B�e����;�@�;9�M@[؎�/�"�r�ZL���V&Ŷ&U��;XN��/��	�*eL������������W��N�b����K*×����}*��0�j�ᕕ�dA��Y$�D�y�i,HC]@��"�yY��B����j�����Y]�k/��vwj�yѥ#@Ŋ����ڑ/Xbn��j���h�I�Ñ�T����6��2�W�-v��cĮq�lӭ��/��B��}$�WE�O�GF�ʊ��	��!�	rȤ;�V�Pfͮ���1��Cavk��YK ����	��ud��Ӛ�՚���.ۈ@uN͊�\��Ȥ��$ÛI-�+7���2g	��i���EE��o-���rv�2j���윯!]�]+`I%`w}�X9�珑=&��2��z�v4��Т�:�Q���ͧAVM�T�<]o]����i�M0��3�!�K���1��e��_+Q#o].����׀ᠩ��v�[�WC��5�'r�W��y��3w}�%���iP����m���8��:�]���˦���z�e��7P�R�����4�Zr�}����ަ��\֔��^�G2��B+'1�XVĩՂ�ؒ2K����ܩ�˰́E�l_WQ����Y���� ���%K���1QZ�-�h�����F0D�V��iEUKj���TP�(���Q��H��b*(�`�X*��kJ�1�6���(�mPD!iQT4у���P����X�#EUZ�DUb��uj"�Ҩ*"�+("��W�6�#G2�A0dUq,E4��Db��Q�m����m�.�E6E#[B��vf(��b(*���**��q���U�i��$E�2�TQkDV1"��"��X*���Dt阭�X$Q�V1rՈ�QL���s�J,S�Ҡ�*
��TQDAQAX�̶*nԕ�������ȫRUA����e�*���"�EUTk%Vڂ*�`�Fq,DTTf�&�TAJ�b�V1
���˼�Ɡz���Yn�ե|��y�xu6>��z�r!S)�Wy̠t�}2�U%5��P�nvX�<*uP�y�z#��va��By=S?Dc����ږ:p6�{Y��;`0�'^��t�o��89[��eQ'+_v�9ԡn3�,����$������t�v8Ȩ�/��,�>���ҕꪓ����~�(�aru6�]�>24�\�ob�=��s�sB6z�ÊMY|,��[�=��{��A7ٍ���d�}��N,�L61��եC^���o��|q_s�U�_(�j�z�c�s�Pwu͞3P��z�ފ������)�=�uj��o��s�؂ej�^4L�8���:�;e���н�Z�L=��q^��˫}�����}�L��+�V�qs�s�z%��st�'�7:=9��<'���c\{��y��C�*��˾l��t�LĶ(�S9i� �}����]�H
��-Q�[:��7���Ez��]��x��7�vzX�-�u<�R����7X����GZ���#z�393�ޝ������: �����{�F�y[�p���4�.i1ž���F5O��y��i��&�5l�[6wY�P�m��NC�\w;S�:en��n�zN�*��O8o��d��u�G7A96+��N�S��v���W�}�}�:y�m1��Z뱿<��F�30a�-�lh�Ӕ:_����J�Rݿ�r|����Y#y;�Fcv�{ڭ�SY��o]S6��^�h�ڛ�����1݁9�"�L�x#�K���|��Lf��Ӳ�����>5�Dٷ�����k�İ*{��!��ͽ��A���$�o�p3������|�^'&oU�����r�qd�8s��7t'z�L	�b�{腬�y�&<�y� ��A�U�ږBb�X���Ls���,�y����V=��o/�x��4�V*���k��L~���Y�sփ�Ow�?y^�����9@���{Ъ�ȶ��^}<�<��2���0���N=��{�}�<��t3ד��h[�ijº�vR=K!7S;[�ns����'�����c<�|�������*�Z6k�ZP�kӠ��S�Ә�S;�,mL�c\S?�{|<���~
��s���4��s3�p���&��
��K7[�\��$Z�gk�z��M&%�;;�}�� �޽:٭��ux��m��m�+�����s��G,��վ"�=�mw���7�{�P��Fz�;,)��vD�\��<�}��c'K�{6׻`^��� ��߻�aް��S���U,�}u����Ts7{0u�v�@�x����;h5�����n�����N��8繣�:]���;����\��~�;��C���]�~��2ʝO:M5��Xp���=v�:B�x�v�H�݊���U�v���n߸z��\�*�a6�8���@��Ixs�{�+��3��\�T�M��(-O���\c���X4��z4<6�	7�U�\������g^�o���}��4�(�X��๡��Y��[��&c4S�P6xA�(.�yۓpp�Lv�~|��5�j6+:��a�s��$��N�Jv�Yi��3h�d��f;�����h��d���x����Nۍ�ƌ�[�ui�#�l�s׃i�;ik�]�H˼<�:1��Iȯ�g��Ţ�]Y��ɻO)�)e���a>�+��j�-���T���˰�;_���꯫�OGvW�za���:���|�ʓ�J:̵�Q���eK�Y�����d
h�U�rٵ�Y��
f\��"5㷽uqf[�= �.6�U��V���o?_j�N+�>��|��'~�l��+~����&ߨn��:tߒ�\]h��X�>�x6VQ�`�o:|����v�4����9������SC.Ax��t���e�������i'�NW�Cj�畻�zu���Nӂ8e���Qq)��eE�f�H�m�֭�Z���רtq;��+�xk� |�����h�^�,�6��44�vx�'�z�y�|��a��~�i��qA�X�}��<^إ��͛��ڟv&Mu�[�|߻��)���y��R>������v�~�q�]7�������iQ�+�����q����I�4����ɻţ�ExF��P�3��[:{ԝﳎ)���\���2�&���P�d<�[.k/rh'���Bv�)�Tr.��K���˝���^��[q�V�9j莺D��_/��]gl2��{Btܮ��)�yX�糝�k�R��_uZ�����������N�~2X���}B[D�@�Hs�g����k+���ksV����4)����I��Am������{`/F���d֚�v�m2�Wں�wvŕ�;��<1~|Ԏ�#�TM����3걝�2K7�{v�l�j��	��ʫq���hkT�M��+�M�v&�q�غ�T����wc2�
M�c[��QN'��A�/�	m�ύ�@M"y��\��^�3.@���-c6o"n��1��v
��An��3C�*�q�P�]���o~�:_:)���W���n`�}Y��-fx����9�����3�U�r��Jy�ps%�&��u��3���U�ݏ,��y���b��c6��j�����',�����k�-�΋J�=�)|�N��9���1�w�ː������V.�P!��*�ϝK͓����vX�����J�fLN�cZ���;�����Wd�ڰ��f��5DV�\��_�w�j�
��l ��=b�蠟W6�8h��+sج�>�����,S{"���vj.l�Z�n�ķ����]y�X�t��WoBL���ç�}Ε�z��+��N�w��qՁf4�U�+t=�ww_M�'q.�t�}�v�ζ.���%nv�%�
J���#x0�<Zw� >}���ݮ�n�W���b�+UP�3�׎��/@�øL��93�iΈ���LU�!�VU�v���]~:�JK�C����ˉuf�����}y�9�7ʸc� �I>��i��v[�^���b��49H�������5����ӱ���'^���=�sh�[��߽�=�ݨz��Ns˛I�aN��A�L��N����:�����W��ݳ\֐P��<��������ϳԇ�N�d�@a�j�d #|4q3���pSg�z����5���9�M,0>��j(1W0��'�w���0��:,t�WmAa�p���B&l���O��������I�N��&
�`���	�F����^J��oft���Tr����d.��1��҇2�XnA�y,`�ɥtS����^��wA7�jΛ�W��`�e%���Zr�FT�z���5��I���w��xT�������{�2��s,��5v��p�b��W4�4�&i�eܭ:0!p���!VA��ʎ˝@�z�{4���ӐY�<�z:.�����
��e�2�1�$uH��{%�J�t��k�/@*�u����>@X�ϺS:`N���6��[Pql�џ����紼i����������%o�&}Ƙ*���z⫤�{��+��,g������G��wy�Q`���A,:����f��>�`��h3�~�6q�ư7{��{ȇ�̺�����84���6�3���R����>0l8*3�����\|��0/�4,�o�չj����ep��v�V���K��1���Uk9m7GQu%�`�8���<eg���ߦޘ;��X7׆Yh�=Z2�X��nT%�c*7\E<<MP�0K���������s^�m��X!KZe�Za��D�cJ�It�/���-�S�w.�yʴ���P��y��p6�\c�R�󭽩��\$8$2�4�J�S�u��y��c�?hɜ�1ᝯ��v�|�`l[�~0U�Jͻ�O�p��@a���S(S86������l��޹ҵ�dƇv�c��2�z��B{
g-@H�@l��!�|Uf�.	٢��fN�m�;�>�XP�xzSP\�&������V�FŻ�P��v�#�Un�ZY�p�id4w
U���
�ᕜ�،S����t�ܒmu�WÁ#y��W�ꝨR[�<� 9,5�A�5c���о5��X��_T3�\�뒄k��ֶb��F��9ҵ]n��j��� \���Z�=6���W�> 9�Y�^�]�xvW�M�n���։�����Y��u�Z]�bxҔ\@�iR��szs�Y�ك!7zJa|������pt���'1�daaѡ��О�i��F���$� �_��W�ЕƠo��'��N�>�&*�wQ^���xԳK�����LH�KS�����8}f���*UN�'���VK������j�D����bh;�.���徶��F�"w��#6��Nj����oυ �� H�g�`�S�)٬����{zy����apV�ڌ>�V=CV�pw�03ϙQj3o��@ܗ��" 	�Z�rR咬���f�Dz�W�����w��]8)�0�0�� �v�;�����;����pQ���ύ�5��jT)�ORr�G��綉��G�n�7�T2f|�#��Te�
�z�[3v�o<�]t9e��
��B��u�u�p����՚���J~�"nY�+��s7M�;\4Xe�����W;���R�)�t�Ο�T��G/�R�
�9�lb�~!`���]S��A`UR��n��_G����}���^%I*���XX�uޫ��y�{�d�/B'<�-P�]�y�n�d�R;��t^I+�H�[K����n>�����J<h�1�Ӿ_1��<pvwƊ��*VpG� >�ݢ���K.���W��u��aԫo`�����j\"�L(��PD��ȭ�l���eC7�=	��^� �2Z���r�J����.�X�;���^�p{��l_�w��Tst�CƲC������Ʊ��(2!�|��ԝ'�!1��~���{����N�VJ���(E���x<<��I���&��{ܧx��T�5A\C�`9B�N�hҪ]�D\�H<�MGxJ�xfx{���o�s��S;%,����W��[�TtUxV9{VM
�b�sć��ze�:�f��e�>����\�������J���X8}VPy�	�a�t)4�'�;�f���zw]K�z,�z��V�֙�vQ���E�!��[�T�u�"��M���v��d]J=��1y��AB#�T����Vo�C=��d����,_���I��7^�u�slW��Fo����{�gj ����^��K.�*~^�i��5*T�I9*Ν[^�V�eͧ�j�p��^%�7}��񨡴5��}w��^��ji��9�F��o:�]��-�/�ل���������E>f�ʵ�f�K@�jo@�W��&� 0>��;�W���|o��Le�� <Gc������-wU�������ɞޖ�#r��-��������nIR\���	�b���T�@8U�s(.���S���}�1V��U�g|B��}��^.���a�B��8>Ea�5K���^V��uZT�{�E��2�<jS>��mL�9����	�0��kpH���^3��������+��d�b]�������@�3�M�6�V&t�OHS���V�@{��Wmd֢�5��r�{�+C+Ԗ�	�j�P��Dߖ�:A��Ys�U�4�t2`�׈��n��x���A�U3�U�Z8:�o�����4���������!�k7����˼\R���N�0�K����	�X/��N��r�eҡ��ߏiگh5�`�̥�Zα�!��T�A����`%޸۟(3���U�Ll�^�r��Q��ō�F���k���!^{<i�����l��Q�p*g�ey
kh�Dh�ts%��s��fOW�|��~�=��
w�U�<$��^�8��`
)EUfRZ���E�1m�+�i�dV`?M(��V���Ӕ7�_s�x���U)diA⮱Z�������Lf��$�K��k�0"��]�}3���P��C�F#�t�;�D�2Kb����Gq�`�	��Ź��t���gf�&�	�W`T��y�X�(P��!��x/	E.��$����Μ&;P"oh��׹V��vr���tk:�i�;��KK= �R�Q<bvi7V�:崰R�y��eKĜ�� ��E��`��HX���f@� ^�钺�nL]��T�hFIq�+Eq2䊱h{�o�Z��ڹv�\o"E�d��ww�Џai�rŻW�j',��hs
������]J�,@�b��t����'���3�b���.����,1WN�{Ҁ�"������.TT��z6��ܝ��\�a�Ѧ�Q쭾¥�W!p]#V7�t��$������R��@s��pnx��Dni�\���J�MMR��tX;+� ��Vs2�*)d���gT��ɔ�xV���6�Qynv�d�q䫻���B>C�bޙX�2������X�Y��l;����A�¦�oL�A.�[�7;D�,��;7Nr/j�<��#v�ҩ�i���G-�d֥���Ј���l��'dӡ�sl�7L�s����d�}���m��W0'A��\oxݖ�����ī�u�._b�k }�,�X��n��s5o[Z�ʏC�]u��Jr�%��R貞�ˈ�=[����ܢ��qD�x�h�t��CG5-�vd�!�D�ǩ]��w�h�cH�x7���X�5����(:V&].��B�s)�T�z�ֻ��궲�9�r���ͽ"����]�ub�Gj�o��{X�%��4�κe�u��{Ԓ���m����Y2��i��l&7�#F`�ibX!G��PB�x�TkZN�Ca���]�N䅗�J�C]r6�[c�)=����d�z�Oܠu�{O	�v��*�f˝#�]�ͦ05�L��ʹ��ŭ���P$ޓ��^>8�AH~<KO��uC�C��.볅�(�<��̮��ܖ�4����7��fV;��V�3�Vi�s��;%cV.e6낉V�c�5+��+x���['k���i��Gc��nRH�ἂ�aV��y:��������zD��Jv�6E�Ю��n�w�u�97��L��0oB������lu�k�,E��WL����7Q�br�瑪�5��Y����)>���ø��,*�z2�uh3���]�T�s�sU���Ǣ�g��p,�@
iN���l��}���[�IǑEO��|#}����*���]_���jY�c~c��cp�x;��b.����}ϵ!��+�Gvk�����@˗�]c!J8%^e�o�!�ppno-ᯬ�9��oWn�p"{7{L[Df���}4�*�X�����K��f&�.��ʚXEp�ݹ$�����1ݚ���T�Wd;0Ŭ_O�w~>���j�Eb*��1V(�Q�EX���ڂ�[DR�$��,EEAEE�[��dQ��PKk�j��AV6�Fm�,U7K1*��HS)U���,����b��h�DV��Q2�8±UU����,UQQc"��V
��*�+7B��Q�,"�T+�*i�1���m�ff�UX���Ȋ
*V�*13.*��"*QAQEG,��QT�,b���EUA�v�AEb�1"*�EY��a`�-TTUTS(�QT�)��s
�Ub"�#mDIE�QJ�Tr�QQb�w�1˴��*�(��T�11��*E��X�ň�E��r��PQEE��PX(�U��R���T��U*�+T�ĭUEb-V�hL]��[ټڝ�����i���ղ���q�m���ӗ��e��70�WC$�����gZ3��ڷ�b+�:�� >�o{qs�)>"�?��$�����f\���8-���,�7�v�Şɔv.@��%:��+�ߩ�:pc�9`�<kG�s�l��8���)��*X�X�Ikާ�Vh����6f��bd�9>��j"�i��ȋ�YV���m�a�58�K�P̶��oFF
�,��ge���j��M8&u�x�A4G��ПKTL�1#�GIo�߹.����zv���Fٯ	l��N:V�4(^��<��%�8��f������=9n���Ѓ�-�U��}Q��*�yo%�uz�Ȥld�WJ�B9��{^u�}įJY!��[���{Cb�ϫ�0�Õڛמ/v��p��������6L���*���w���حӀ� #���J��|�o�,nM(����iR����9�=�G�f]d���#����x:���}3֩�3i�����5�(A= ����vN:�k`m�Y�N���rz��6�[�ϲY��u��^})RzVcՃ ���d3���ST�IegYف����~� h�,d�;0X���g��"�ٽ�/�`�Ŏ�D�4�Wd�[�҃��a]��=}��%�R�̧������MU�i89��{��H<��
���kç�9�l��F�����*/Ɠ�����:����A�w�]�w�f7�P
�aؽ+�B�
]jZv�'7�>���:=�'��O\�y����8���yeo�E�s����+D�X'�URW3�1�ŋ.86�no��d:B�;��8��,$A��8�OrčO��Y�}$�5G-d�;{ծbe�P��tq�_ �8��|:Hȹ*���q�fb�&(t��+NE"����|��J��<0����&��{V��������Y�e���A�.��8C�G)��͞=��=���}@�@DՒ�b������G�/-pڄYbP��#n��Ӓ�<�z�^nQ*�K�P2�:��*PUU��V��hNi��J"�j�F�+��������l��<'6YFf�U�S)���u~�*�|F�tة����(:���ݕ�Fzw��}��Y�"GV������0��s�紦uĐmc H�g܄o1εĨ��n;�ot�[ײ���w	^�[�0i���o46�Nkɽ�YO�Ո�@I���gl9�4�gbpsQ�7�2���<���@Ѕ7�gt�2s�J�nن	4�|q�3�]%ո���R�p5�/�5j����eF��L�����јI��,%0���X]<�S�;�)�;�[�0�7Sf�=VV��z� ����K����������d��E��v���%S��Kk�;x�=V�J��z���X:��>�-
�U7g��z�]�iш�\j?���$`���Z(/i��!�P���CN�=Uޗ�R�|�|/|��oFoW��]��]�=ACFҮb86�b��?��1���gUr��O0��u+^�N���}�٨�\���N]֞�,������������0�=6�cɅ?��{�V��-�ODJ��	].�M뾣�EP���(�@�d���4�������K�P��mX�y-;��87��3K�>�^}��\��*����[�us�7�h<*�.��૕)cH/�����Cᣄ��u}�"{��I�hӔ�Qw��~F��W�Y�w¹�Vhpq#����������<��������N\�!���T��C<+��xR��]R�z%.Z$^I�^��osѲ�$��̅��߳���x1t%w�O�΂�ʐ�u�X5���C�õ�r/��l�~h�#ր�����wSxZ�����q.����)���	���jR�6�56���u+8:��Y>����#vAZ�c�<�ס�ͱ�t�����k�m,[������m-7;s�<7�׭��k�"���/2�I�	y;C���3�n'k��G�1����㮝o�H����ާ��<��ߧm@�R�a|�+)�>�(������u"S�6���v���C7.g*lM@�S���&�m�	+�B`�׫'����u�@��y"[��r8Ǯ��t<�%���x�f�)S�sA@plhe��w>S�84MX��7�V����n�va�l��bj�p(�Ksw�c�&a�uCyi��i�<��jzTZ�a͡sܞ�ޭ�~;4ll��h�3��g)9��]�c�w���X��<)E7�j��n+Hd�������6�2��.;��M��|�,�K,�P��������P�w�ٗ�j�X������^�p2�7�A{ք<��/z���͎Z��(4+�첌�ɪ_�k��~8�J�P�-�Z�-.�S�x�M��c�Ul���MB����&J����N����/�W�2��cՐ��'�����ħS���áݾ7� �:���罫o;�m��*����U���ɋ��Z89��O��ұT-tWk���B���{��ң���!Nz߹���X�����䕕�i �r�F)�*��{�b�+���P��vx4��5�k��l�w�Uc�i�s14�j�WH-pw�M�ܧ���{����݀���R"���;����[ �������T������E�e�~y�q���fK�K��B� Oq�����u��[������g���-ļ���Y6�
���*�ϸ�QC_�4�E����P�I��ݶ�o���-u$�����Do��@ߙ���x���#�eXό�F��E:A�T�����C�	�<�����-�Ӈ�긃��C��r�A�;�<G�%�s�qeXϓN�UY��|.Y�`�Y
�~K�ka>���T+FXt*�F3��k9�&���5�;B�}o�Ǵn�,3N��u�;ιo�9+�R�%+ `�>KA������[�Ձ��>	�!$�4��(�-����U�c}��O�V]7�YB�JVi��f��@�x� �~34&:��w<M�~Vm��{���"{�Ut1�C��+�	f�|��d��>�AVG���:�;�+Uw��g�OVn���fv�A�ԛz�U�	~���
V�o\A���ҿC�>����{�mm������6��]����{�0;���6ͼ�P�%{���kB��b�8V��s�vQ9V��}����l�n�0��hCGH��@�c����ט�sm�ș�`���.ћ�)Ns۸$������f:�	K�VM�%�R߷���E�w٢j��ά�.��UR\V��;�dԟ3�ǔ�[ ����Y�یEy՘��`�Z���[��4G+}�i���%��[^�ౚCＯ��v�z�-�����l��7z��W5篔�RuG��/:N˥�԰!�ԴOP�| �����u0E�Ú��te�=Ws:��g9�L�����'L�-�j�������0�u�C��/��*y9T�X�Y��<|�8�T�����~���DfYhK�,e:�
5������l�I��dQs�N�j�5������_�b�}-��c�*{f@ͺ+�:�ҮS!
�C����u漉���]�4��\ZK���0T�ll�T/���f\X)�\%:N%�* �b�\Ѧ.���k�ʪ�=Md:B�vg�\c�P��a#$���F�¥y�\~���F\o�}�����7n���(]zv�X˖�!�p�9��Al��ovTۼ�z�J��e� [�!8�S���q��Q��Z�뎡U�Ϝ�G�E�I�ܰԊ'k��{:��;K������W�Š��.�]f��Sp�#�o���k��n�W\��"
��G �ڕ�";��=���r��&�ڼ�M��o;4>�����<��PL�M.�p(y�4�EJ�v����ﵻ�@=�+{Q�v�{+]p�{	u������x����.�l���;=;��]tL>μpG�����w��ή^L#��ґ���a�1�*�K���UR\�_[�κͰ���R!{ٙw��}�r<���a
����醊��b� ��r:�*n�b+�Ԯ�8:���4`��Y����y�9��9���`��nc1]�6��=�hT�ҧ�8���fU�q�C�#cԵ	C/2���o".�����$f%l`>V��v�gJ��n82��֚���Ō��e�͎ }\\�>��y��T��7c��w�U��/L�;���U���K�,��Ëy���7��C���W�6ǐ�YB��L�=fug�V�/m����-;��1��5��gf�86_�����''����m^L���K�!z����"����k/ZLZ����7�8�	�}~����N�	��|��F��ܨz�EJ�<�^wm-�D���ftlҺ�[�T�<�&0?n����nEpO�'6���U�4}�ǅl9ᔨ��lf�t^���M�HT ���˹\�]��B�R>2���uO:�ʱ+x�d����U��o(B���[�V� ڧ��%^�����q�wtM���V�j ���BV���Ǯ����(�f޻�^�����L_T�+g��]�@9y!�A�5]	���ϲ�j��;�;ꝥ��s�[�[���+z����oy�����z_w;���h���^2��Ԥ��4��S��6x0��FF
tH!�>�
ӝx[�cEUd�X��w���>&tk�hC��J�&�+��oǦn�w5p.�x>�Sn=q-~{�^*�w�tY�{�i�X8!���,D�$X����]�`rƩ�Sᱱ��^(V�c�=0��T4� ��qg�}Q�^�U�XN�A���p5�Ma�g����{��|���}K�Fxm�sMP��-O^ ļ+8}VPy��[T���Lzh5���<���Z�:���L_R�F��LCp���B���1b*��+ ���f��֓�o�^��UF��W���
��r>�QJ��V�F��3Ú4�8#�B�q�/�7("gxίT�<��@�tڼ��oX�Z����愱b�OPT�@=(]�i�3C��T`a��#��/i�^z�Ժ�@7w2�ϝ���[������%9VO��g]K�>���.Os.���%6^�g�VÕ�CjN���5V�~�aZ#][�5Xn�W�x����������"淞���뫮���l�Kz����7F,q��ᆘ�!5�L�a::#��y�w�e�!�޻n��e���hڬWW;����x%�T5y��=�rJ��O,d�XR�V ���8�_Ȝ5itX�j���R𫮗�/K=�_%=���.�4�(��+Vۦq�:�%�g�Nv�ve%6cz/���ħ,��xP�į`�}Z:Xw�x7S�և�V�[�P�]93Jƹ�W����2lA�b�W3Dn�~�d;�+�Y��V�\V��tj��9t�Ӧ8>v�?��;����ʾ�G�][�op�T{�%��p[�^W}N�K�FOn�������U3�h��p'���7T>G��s����%}t"¨vI��k���G���1|�v�c�f�8��b3"p�?e���dX#��:V�E��lx��A�\Ći��SRy=��ڬ-�NK�,�5��j�<�(zD�ȩ-U��(ɨ�t�5C���yot��V�R����(H:���gsqø}�3��X�����9�����ŻbFn���X�*4���POF���*�Y�u��-�]z�=­�ZNR�tnP����䘮���H�64��ٱ�ѥp%+4�}F��w�UzK���ȣ+��Wmׇ/{���O}�[����f�ڢ��ܪ7[c�s�Y����J�����Y��λ髴�'_��wċ��ǹԜ��͂z���WvP��I`���3x��:�����v{g|g0�V��m��Mt�����fssZ9���3����=��CjV���9��[g0���JW
L����p"��j�r��(Mv)G8�QRFw��/H�n��2��wLt�h-�Bu��䘘�^����zX����܆cs�c[���8����*�9�����'�:0��
�O=Є뭑a�����O>d������g��l~�4�e~�ʢ���'.��mu�6�K!a�YѴ�
m	��<���١�f�
���9J��<�A}��/+�r�C�J�v������,u��s��i��.�����˛�;��V�U��*��J���T�)��UU�W�Y>�St�G�T�wc����������ʹ���y�[>���uH�3�iC'R��r�=>���K"��p���b^�3��v�Q�[*T3S�(�m�Q�e	���z��I�q8�ˊС���m�9)#v�3�;��d���z@e*Y-�w���c��j>��G�8f�:�4�<S��v�}�Fzj�~��2fS�d���.w���Z��Ӑ�ފ|+�ﱱC�+�:�D��	�3v�������h��kZS/]�Y톬MSk�O.�T��n��q����P����V�<�}Y}W�:=ȝ<"�X�j`kY6�o:qU�w�v��0��y�܂frjK���Öl>&uo�fv�ɭ^�}�B �Z'	Y��Up�ة��Y�;4K�メ���D��+��Lo���ع�YM<[bo݁B{�����ӨNK��/Qc
�7:H���m&�jWKd뾴
b��f�kt��MӘ����@��9��!
�yZ:J����6��[��\�r�{�[H��ŁVf�x�̏i.0��-��o�tJ!L���
�{:�Er�MQ�Tﳟ8��q���gBR� Zټ�N�����p��2��>��uK�Z�+�w��fۑ��@t�`��/������J0�#^��!�G���3��t�3�V8Yo��͛���3�@��dȪ����wLp��J�WOvʷ[�v*��k�J��H���j��ҫU�aܩ�u�z䭮�Uk#(�r��s���w��Щe2(h�����y�.c\���櫕Sa����p���,�Z����@�K�B.x���S����7�xjw���U>�䞇�us_uEsp�`���V��X�so2�!|p�*B*�]YV,[-�r���tBNxE���=��/�ݴ�<�!��p,,m�x��34�(�
�6����`�2}�t�؏%5���+��Z�r���{.�m�ѭؙWKn�*��y:��V]]��+�+�]#��3���Zbd��V��̅�f��g}�鵏E
�ԩt��YBj��V�	�MF�.Ջ�/44��*{�݈��!�ͱds�ݴnb�������u;#����o�E.��鼩.�u\H��O��<�^c�]���pu�-��B��� $�6���x67|7��w��֜`���7����bT�=I�6����Z�T��a��ą��=\澵��ȋu%|	�w'u���ss�2���t�w�p��
��.����#���*�oz�����{CM8���C���,k�V p����W��i��́�9��݂Q}�U �a�������,��GZ�ka1�.ھԘ�جI@��Ǐ�P���A,��&�b���^j'+���ַ>���>��i����D���%�oo-�.����WKZJ�L��ԟ��F6��v����S�gu�F7Z���a�p��W���k�ޢ��PoV�Ë���Sf*��WZ!���F��GJ�J�f� �����kШc�[���!x�hl��U���� �Q��\�&Wv��f��ќ9Թ1ٗF�^(���	�l4Z�۵��W':e�t1SlJ�;��i�`�٧�aס���qhrIu�x�2GVG.\����>Ң
M�\�����;=;�2��S[�;�gx;ťc��k�=�2�WS�A�95���yK�5+�gI�O��#�֋�L;[�9ގK�V&�ޥU�۪c[��xy�H�X�m�1<j �	�e��r�Ab�j�5EQ ��V���*:f�:AZ��(-���(�`!�,L��&!��Q���aR�F����TFbi�U
�U)T�i`"m�jܶZ���E����D��YT`�2նUZ����V�[Uh�m̈�[*QF�Q��aZ���Dm�ˑkKd�FZQ-�Z�	J�Q�ih�e�Z�1-�e��V��6���$��!c�\mb֬D`�b���kjZ��!������w�D�e�Z����Sm*�+��U(�%L�cQj��+KK��m��TAX�YAV���i�����R�m�`����Ak(�J0��UE)j�e��Q[ZJڕV�mQZ���Ue����AH��������@���7�I*�T�QѪv��c,�B�9ڶ�p�g�'����?d�����bu+.��=���InUҐ��6<�0N�`�����N78n*����R�N�q�)\���q�.R����y"g��6Ю�Nt���y:�v��!���u&.\8��.�:�8r�>��>��Ü�%L�!�e��r²����&��W��؋�d��w��#���Ϥ�9�akVK�H�oF��qx��U�+D�ޚ��ؤN�J�|��R�Q0�/It�]f��Y�:�`��8<�ݜ�����z?tyT�����z��ڂ�T��
�|, ��N�Ru�Z��\N�T��2l�g̢��|���?i�L���<�ϵ�4P2��K���'��겾�R��򺕒���]��륈��.�mg��Y�S��W�cY��BV��,y�+��+�����+]��\���(�ӕ���	_L`��B��k�He��0*t��*�s:�C���ͳ�O"��*C�\O\�ɬ�Sk����1q"�AS|b.�b�w��+���Xu)�W뻧
��^�L���7��)} z�����ӯ����TG��Y5��h��=�����-�J z�Pk]`�B�y
��^�ZS7D�)%W֑�ҟ��ݨ�[���N�u�Mr�v�`!	�.i#�V��ÎC!�b�.��ގ 9�,�)A/4���O�zr����X+w���n��(��`��j�vRI���Z������E+]�zXq��E�FN���pS?vÕ�h���O����]��F�B�HJ�,�*��0�Yb^��tq�z� ��N��넭.�zLN���V��ϧE�bS��v��{�U����ޣ�Χ|	���9Dr��t��tW�;�\<;�L֮㢍�zR�n�k����ΰ�O����.�]JKG8��{B��>������^��70���ܧ�c7AQ��0y�N���V]�B�Z1���]O��)Ԭ�vb0]Z��ч�%.Q�b��Sv<�>����%UBtd��_1lU�y`�a�� ���j���4/,��R1�m����Fzd�~�X8�Y�.�p_�D�,BPٴ,D��"�����z�øOJ��iæ�-ue���y���i[�uL���Fn�V�Ռ
L�phK�h��w2�.��N���f�(�JO��\[��r�G���@�T.��<,�S�V���JU������Ĉ~ޫ���̓������9�k���'X��ϵ�D7,\�bׂ����pcL\�*�򤴩���5u�_ekو�:D�:�[.�����__�5��^�m)\]:̞^u�U+w�Zz�BL�F(�d�u��A���.P���Xm�8#ػ���]�:�X���lw�-��gCH��s���1�>�9��"��(f�E׵�TXܰ.�m,�9e�L��t�umu���싥S|<�]Gj��Q��5�p����}r�]Z�N��0kE+>n��-�|��V��z�4�=S9X��p�@����EX�S��!&�)�O<�-f�}S2�Ŕ�-}�n3[f�z�v�4�*���I���z#�F��h��M���o����p�!�o
U�qf��V;��R:���# /Y��u�~{|f�>�4/vR3f_0���襖\��qrxr� �v+��:��Ւ�P��w�<���_��'.�zt=�"X���ul�R�ʌm�Y�%g��ߩ�ݬ=P_Z��{I}��C9}�+��C�u)��u�B��Y�t�������[�hہ*�Ծ�/<n����qZ,�6�w	�.��9P��lu���Vko��H��K�����Ϻ�q��(:ñ��Av���]�:_e�N�K_m��[�͜���g����y�%�f~��6�~���wо���h�g&u��޽��q@��{X�I��+���[��k�izr~*�*B����^wι��(Q<���Ƿ�5]�ǭU�E�s��y�3q<�Y+&Һ���ݧ���@��کs�`k ��,�w�Uȕ���k�M�0�gR��6\65�ظi���F����w�qb�S�����}I�u<�x�������e{�}�,f�XK�簧^G���PbS˘	�30&+_L
��D�qrm��$n�1~��s���9���Y񖰉"^G�8��Vp��r��TO��y���4UUD��^&��+QF[��/G��s�2U�7^��sf,��k�Lލ��)*��#��;�j��`fg�}F�۾������A��T���H-�>�̛�M��|��VJ�ʥ�DD���u7�=@���d��_]�O
��GՆ� ��1�lHۭ���p�.1����wSb��j�gӪ��"5oj����C�}�4��R��j� ���ch�è�|�Ҩ9�T�|���=ZJ�pUy�[�Bż��w�[�)5�R��0�a�qpJe'�-��Ow�փ�q�Q���fl,��\��F���ї2.�y�̂sPXaY��Ō��q��v�h�0}1�*���i1�H}x��_�͵�/%��OK�7�����o�N"�b�=t��ZO/Pw��V��W֎O-����D3͋�Gz%�<���H��ADඅ�������>�<)�U�+�>#|�X�{���F��;ͣK�!�(�r9� 
qJ��kR��)����R������ӏ��!���Q�C1�W\�gd��U���,TEM��q����,��禲��r���|d3�k]�Y灡�%��U�G!�7I����\iU���I!T^�L�,���S.5�����[�u%��'e��6���g+;4�
=mǫ|wc���zF�N���k9��eg���"�zeB�l���B�J��Y�mT|ϋ�����v���#��%��z���zB�=��;-���ӫc:��}~9���Y�]S�����U L���!ы�z�u�}�(k谑��!�f��]#��.݀�����*Q�6}r���6.^�9V�*D�:Z�T�y�����<�X�f��׷�D7��=�@7RH.��ŻL�Pb��[8��fQ�u_��6N����ԯ-�8�H��k��BԻ�b+x��b>�'r����P�-���.���/+��:R�Y2�'�Nw�Z5��;�A<�C�<�]��'�ؚ>�Y�ׁݑu�1z��&I��a]�g�~B�E���XL���f�fDߥ���{FeG�
B��b.<���A�j�,����Џ���k�{���^.���$i|*.�@�+�k@��_Uu�\8Cz3+Ѧty0�_t����RuN��
&�1�,-�\��-]L��V��-3��eK��g^u޳��05&uESu،��j��}N��M��޷t��������'V�E���$%{z���T�үi�lݧ���cxz-����{!�
�$8��a��U�-]!����|���eg+Ꝯ�ySߤسj�/�4�h����*�9�\A�����)��H�T�]��Ĥ�S�*
�N#oD0�����u���q���Q�Z6ڿ��5VJ�N�G>0U����'0�]P+��,y�s�.�6e��S'k��+L��z�f-1�Z��eT0c�L0���M�Ch�%K�V�����k\;�$���v̧�u^!n���.�ݺf��Gf�i�z��
�e���
�����d��-ק��[��(u[�]�pg��I`jUI����z�1��*=C�����?�B�:��t�(zr�G�_x:"V9��Ykf�]�5/� �%(�V8�c��WʏPG�Ap�u9��cGJ������֓Ʈۋz�v2�l�1�#"�7�FP�D��p�O�z����'k�A��=�*H��0�����iiǕ3=i�Jt�p9ʻn��s��a���T����z&(ѡ�H���dNw;�ռ���b�B�$͠c̊��ybkȡΝv�S�u��MD��Y�5����v���E���k���cl����y���͂.|��+E��=��:�oR�|��H�>;��6�Q������O�b!��{����icS�J���BO����o��*v�ӄ�:E�:�Gjrc����w�C�k<pTeW�\�걡4��	��oa���qy㛹Z����<]�]vej�S�V�ĥc2w��J�Q�=c�t=&��(T�\�ސR�S+��̽�˝T)���|��ϒ�u�5��[2��'�>�E��Pq�&�˚��;��evͻ�CסXE���U���E��k!�R��n'X7֡��4�3r���J!2�{#��Eת%[Y�����^Ҩp���kPsV"�[.�h�4�M%�2C��(�Տ6�����q[��!�P!�UD�*�qv�#պ��٣q�I�R�K�s�('{T��$���+��c����¯���A���6}5V�'giL�g9V�%�7�����{A]Y���n����V���AA
�0R�{q�:��!,oY9�P�޶6��>w�u��?\�:Jf߾R���f��^�C C�,P�=nQ_S����2x0z���rq�ع�-Qșz Y8G]�,�S�ݎ��z.ku�B��VkMSK��Շz$�z'Z��I������+mN_�zw�sc|ܫ�%-��$F\}��̼irΖ�ޏ3s�Q��mѺ��[���My�BX��_�Nm<?>Jؖ�����6��r��T���[tW�꧝���b�Cv��oӟ��XUw�}3в{M��r��,;��rݪ�'�֌�:˖�y�!��Om�ɗ����.�@�_a�����^Stf�e��J��E\)^� �mp<�g6��4�U����v�Xb�d.��8�9��/g��M�Խ�4�(S��N]1����&T���^р��cI���ex'~�0[�{�s*f�w�\�ݑPe�$�Fnj�p��j�o���(M�޴3#ͭV���W �9j��5�0A�2��<�D݌1|���u�>�����T5LH�&X<$�vj(�t��^[�0��52��'z��aO��e�ϫR�Y�sM�w(т�S���a=F���	�i{={J���B� �=���ӻx״����ŉ����vk.����=D�_Q�}�xe3ƛ�v�b�/��Q���s��~!nN1VoP���K�GW�E�螚lM�f?
�iV���A�5,���k�k�U�Vzg�����s�;(s�Y�v���z��q�,(���Ʊz` ��%����e�<#q#ݗ���+lmn�Z3���sm:Z�:�֌J����/E�whV�n�݈d����U1�
�M��;Fc���S�\���ǭ�~���y�Y2�*���N<�*�h�U{���� �e�)��7�3t��|im���Ĕy��^�AVyz���'P�]�k.�F��
:��=�3w�10�9�N5��{�ܷ~��X#j�W+����W�������A��gY�`p��7�¥�R	���Ī��f�ޜ��`�u�s�b�M�VV��éԴOP���d�i
�� d»5�ڸ��-�a�w��T���sZg���;������>�R���w];_u�E�C�CѿV�=-�g�<��k�C��e�b糪x3}]g�̳� �r4�_PvpU#�ΰ]�p���OĥÉ�^����q��8� �n���Z%��g��E|`�]v+8��hэ�
��@�v0R��l.�;�ĺ���}�\�~sP_M匹u���3ڮ&EH�n�����N
�����|� ��\<�Ws[1z�z��†���}�����lF�{�
f|�s�k�ϮR����g(.ã��b>Ơ���q̂?�p�b�O�u�(0n��@Uv�S�YkX߄��Ÿ�5_�B�3_ey��-�͇�7�P;�+ڒ,�.�,'s�(a�pfvvѰ2���8�{���V��m}�ԏ��o��wJ�\�o��s�*��v�o	�\��=�7��d>;�9�RT����Mg0]`f#a ����[������l�R��(�W\ϰ(��6�:~�n{A�;_h�v���\�Qϭ��d2��ϓ�@�_[�E[��8Oz���5��,�ě�|�i0/dBR5�q��#���
��� /���諆�X�Q��V�������ּ�Vp�@.�Z�Y����}�����h�e1R�3����U��f��W���ӧ=4L�Bǲ��蔯!�N�dYφ�!+>޽�Ǜ@�ˀ��{Օ���n>���V��Ԋ�*:,���Mĥ|0(�L-���� ���T`�9���y��a�󙴏�����/������o�z�!�E��,S�+hǠ�����p2Sg���0�M����>{�cS���{V���z�պ�ӈ�G>3�V�z{ݒV^b1���a��)~�x�w/�w�T�|f�\��O�G��ض� �_��0R�=Y�[�f!��h�l�P<��\���e��=R�&'QĶ����#�:.��>C_�U��	ֈo&�\#��W}{������jYW�W^@�9��)[5!��uȤ�P���bǅS��6�لW.����Wj�M��0��ۛ�<�X\�u��k\4�D�dv�t�*c~���;J�JP���JN�uU�����$��e��Jm����L�\���ɱ᳥�j�k���1��ܣ\��cv]�2�l�:'V�rݮǗ�����鮢���̥��KY)ޤ�K�W1�7��O�k���ǒ�𚶗*
�a��!��y�h��v�ëq�Q����&ܓ;o���2��1(����DD��b��
���n�t!͌��˧q��)��u`'wi�Зc�e�*�=u"���9^Tw� �Қ[WS.�Pv;4�	�)<�T6ƈ�BcJ�;�R�$wΦb83-r\���{͘�i��c��*=r��h���y�,kV�;��bn�>$��Wq��U���0-t�g>��o�rvI9��Pnv� ��B��˷eq�	)_v=q.��p��Qە�=V'!�-<�d`Ya�by2C��z�,[�V#���,���{/��#�ݹD��Er��-j��u�>T��n]d�t��[���c���oU��[d|2��r�>T��xN��o�>��=��|'e�������� ���~�/u��$WJɭ���V�\Vh�b�޾�Kj�2=����-�z�V�[���}�M�jn{q���1k[������}V�ƃ���x��U�Ğ����V����B��)H��{"қf`�N�w�3ҡ��GwC}<�%��Cæ�ܩyp0�'�F�*�ym8��(�)b(Ig�hp�xp���P���%�!*�Ib)�f�F��S/�XPH�H�oa8�RFAQwH��V��U����e��Ҵ೐��E�Y2<����T J��64�Yjj9E;�#�/s :P�i�)˽�$�n�+q�� I�pfL��Nn3�!��ͮ.�R^d�T���d'fӖ�̸���Kh���mA��
���^����|�v[	���U�n|���>�����IJ�gԕn3R�WX$O"qov.80�Hv�[�Vh��u
cv��xb�Ɩ�]��2�-���V��oJ�t:-��nr�n��+2�^���_u<�'N�����"�R�9��M���Ej�s;oR�U5
��;����a�A@"$v�r�ڭz��C6Jw���]Ƥ�|�Ҥ�X�|�wm������,�g�n$��Zc�"��t���yA���F�vf��x��wЖ���+P	z��T>%�g>�����{za�u'4yU��҃�ҷiT�k������H\t�_rU�:n�w9lJ�jk���E��
5��ئe�+��)lL�]��I�0c /i�:�^͡��vU��_�:�ǯ�i�����nC�MSve�zz� ]��|i
�+�k��p��.��M`W��<G��Z�d��_��|����#4�TG�b�Y��s
�[J��iX%���-�L�䵡kPk
5��YR���Z6[m�+YV4e-iT�G.c_��������R�hһ���Z�)���6�h�E+mcXҕn����[D��ŬE������]e:�L���[t��rS-�un7L���\���U��f#��fU����V��am�e��Z�����-�w�d*�TB�m�5K�J�[miZ�m�7L���E���S-kZZU�V�ҍ�5��A�`�ض�4�#,��Kc)l�Q�QT-��JҨ��SN"��Z�L�)aZ�mPj��mT�R��9���pR�1�ҭV�R֭S)R8:��؛f(�[-�(�X�Dc��Bۘb�Z���-JZ�.��,���h��+X���Bƴ�`�X(�ik�T[j4KU���e�Pm�Ю&��\�(  �G�@� �;��v�82���]����5���jӡս��3�C�8��ֈT7@ښn�F�i�ƺ*��LQ�Z��C���BEWڕ]�%Z%�$�w� ш��\��{��~P>��<�a�����n�gf��=B�:�9Dr�x����u)�4%���eR�i8�FWtӌ�b���V4.
F_W�w��wC��� �^=�T�.�����*{�;/r
AS�����!<g���P3rey�N���V��pmԬ�ݺVUu=Y��It,��qw)�h���f�TzUʈs+�8>��:+�L�����8��Ke��w ��̪]�;��i��Ծ�f��:�"P�6���m�Éݝ\�Y�6�>��&��1]|4^L1�+$�E�DӒ���U�X�jŻt}����]MW&e{�s�:�d��W��|��̭R�jj��D8�-O^1/
�Ҽj���h�v�n��d���t)ש�w���5a{��<��u���]b��Fd�W����֧��]j�/�x����s5����� �F���3N��ݙ�ݞ7#]~��j�SH�\�uBx�vM���(p���:҃�1b�QE4�L��-�N��Uy��� >;�����
Lu(Lں�T���+X6#�_S]C���m!̃�հ�����<�W�x���K1>�I�5��fd�r�C�S$�Y��=�]��Gp>�����3�*Z�O�_��u��w�W{[R�g*p��R.�#���^�Γcg�h��9
�>������Ky>��֮���U�+V[�y��'[Eo�P�mcz��G{^>%t.ݎ�lW�1�z�7P\k4�G*P�������S�|����Ŀ9��w���J�w7ڻ�'�`|�:�;�}G������X)�c-�+�t� ���f�({��f��y�	�������ǔ6����]���x�C�g)jb�%���R��yZ�����N존빻N���gi�3����!����^�R���hD;��n�{뾧HdI���q�������p3�KI�|i���]�ﳘ{���N6πwl�!�B �R������� �b�V[���Os1�w|����n����{\F����U%�1��7�*��5#/gj��.v����B��Ҏ�P�JV��ex,h�����S7	��W(�dW��"�_U݄�le����H����8y֪����0>��a���T�Q������t�d�����<n��1�Yv�Y�b����nv��A���w�b��$��5>��뫞��uְ,:���M5�U�e�_kmC$�T3��M��v4${uux:�oGj�n�^fgB����i2fr ��_$�]ů.J�1�}�H���rY=]�?Q���`
�J(K�2�`�7n��_Q����������Uxt��jv���ͷ5��y&9CW��`����Q�p%+4�z�[������P�{�ָ���]�+�{�A�]6#J�tLa	�,`��vk.�.YB�JV|��<~��i�� Z�ڇ_v�t!�B��v���7��1�sUQ8�hK�^]�K�7�N��Oe���Sg/4v�w��ݼ0}
�C|Eã�����Ps��ӓ«>��I��Uq�QNG ��]���L�Y<hP�U�Z�]7	;�UP�e,'�+���Lu�zo��k�j�+��g���W+k\����au~h5k!�q��^
����*�����&e/6�V��5 �[���s\�l�����
����E�łz�?�R�����"�fk�b�"�VV��6���NE�Q��%Jkֻg?g�!�9K�qVr�W�c1'y}ڛ8:�ׂ�,혼t�%�u	��2���\�u<!�����2��LƂ��u�W��k�9>�ۑB�R���2ل��S\�5tժ� �ǎ�>/���"�T{憤����w��M���wX���W���b� ;ۧ),��l{���Z_P;��2��������R�N��H�O����W����f�-�tNV��vu.��h���
=���s��i:+�����e���~�X.�v�N�����/�Yn��}����R����K0�Q�ӓ�AU�
���p����5�rq�1����^m���4f����ܟU�R�eЩPV����<��C��=��]s\���.�
U׈�0�Q��{�D�m@+�[G_`Ξ�5���D�����|*�U�ׅj2�,�^������!eɯ��++�oc���h����و���d����(b��[8����@���j[��w"��Ƈ�R�j% 2�ztNW2��kE"}�2kpW�TB�F�ʚ##��}k�l��|XN�Z�:Cƴ�|)���u��:Рr� \u�m�ӹv�����_ph)��2�ݹb�����	��Q��f�,T�3]���~�y�aݫ��XD�@���b�1TB�W�s��9��zm0�w���W��^�xp]���S7�H+1��"�30�B�R�HZ���b�cӉea��mUZ�pt�ޞ'ulw8[��=t�q޼�܁����N��0�JԉIP������z�wi��;;_=ЅF���;TL 7���-l��wWyGd�X1��D���ymLs9)�ʏa�j�����UX6y�K�n2Mү��Lqo�Qj3o&oúPW%�
�ĊT��A�� ���
�ɾXVV�c�G�@��=��UV����hoNOz�'\��_��[�Zpo���O�1.�ǇMJ%3_:���*�<���3|�2pF���o��ᑮ��f/���pFy��~m�.W}���CՖb*�P��Eu`Z�$uJS���;���ߺ7����G��zo�յ#'g�=��)��Hq��R��*�}J�?�x�^i��ź��J=���Z�4I�g;��k�6�ݽ7�N�ү��J!|*����8|M���:u��v�p̈>���x�iI���f���uW�G!�|�[�+Eqw�U���4�=Ք
���t�TL�{��	�#<g�nq�X�,E�""Vu�%�����^ ��震��	�#���{Ow$��;ᢄ<�V�NT_;��i�@�V�Ϗ_Q'ЇB�б���9�xV?vxE�5}v�L.z����}i���8.kVU��ס���R`76
�HT6J�B�S���e0,+��[��-��l:9����';���S�R�[ke�i�������ݸ@��`�i��q�Nmg��W�?%]��<�w��:gH�>�R�RJ�}[MN��0я��XI��B:�I�k��{����ڮ۝���ԤŢ�������������r�G��B i^��2�0V���!���x�v�Y쏖�:��KQ����W�շk(z�U�u�.a�S9�XLA[�W��'X���vQ���w�T/h��t
`������h$�,l���IW��J4���Ph�|�����4td�ś�b(�v-��G=�Y�;B�aR.�1˿O?Y� ={R�b�
�7��fe�6���m���=��ڟt�ӟo�TFS�5�T�rT-"�#����;4og�4nTW�N�!F*F:5�sU�他"�;P��������'P�u��h�&�����o��[�Z�Tm�QB�xc��י=c�)��sM��2��Z�}B���}A��N���3j`�9���=�?:�����R�]����d�1	KS�릱��5�E�C��F����{r�w^7�{��G&�wfu^X��q�\0p�k�dq!N�L��0��1p\V��.��ͦ�7�w���팾Ȥ�n�0M���T�Q}��K�lK��A������L]O���W�]���0�K��J�7�������Q]ȱ��-�ǃz0�`�TT����T���9K����J��F�i��ocor��5�1|���Av�P9c��v���_wJ�[]�����m]je�b�:xU��I�Z�WU�vxi#������Uނ�w+�hƼ�c�~{�o�k�r3���o��SM��	��ЇB&���V;�t�/ws�o��b��,iJ0�g|��PC�[��)�=9?^�
�:�Q�1%�X2լ�z�]5��@~�@�]�h���P�I�}}y�'~�6�C��ٙ���W$���EZ��[M.`g��P��^����WQ�����x�]a�r�!U�W'0:�~�.��F�U��X�-ه���ʃ�Ȩ6퉸�K��[�k��e�_`7Nϔjo]H����˚���w�`O�q&K��,����Q�ܦ��3>��4=g����b)��P��W��+�A�]�֝0]�)�tj" ^r�I<&��6�|^W�伹矵����q�#��,g>��JޫT�;��%�*-���F�޺v�����s�!#ǅ����o^��!Ul+�S��(Sq[��V��^�б����}����9�4)\]�W�Kn�WDr��|�b��J!���Ԙ��_����:?z%��p��NO���6�ݰ7C%�Cy�1oS��`��%���2��w���><�{R��=��7Pq/�� �ȭ��r�eb�ۜ *2n:2��`l����Y�Bo>�Μ����E�ȲB��2k{5-eG$��US*5��_���&?}��rժ�`���Z�������y�`�[�:w�1D6Jv�zMɸ��^����]�� ���g�k�t�.o��t_�i����*�w�z��X�r�̦��_U�u5q���O@p�`���*8�]�(���5��x9����vu���ҽ��x���f�r��z��p'N�/�r�(��=G�^����RCr�o��\hc٤Fɘ�׶;�F�r�h�FP�T���;��]t��t��qLa:��;��,g�u�K����NU���+����[\�*�B2�
���)hu�\K���o�՞��Wu�tvؓD�`���q�Y�/��26�U����OV�R'��z�tb��}�s�Y ^�w�ê�-����9u�єo�{h�?'o�W(�}�딠<M����}V�*S�j	�Yfhi�[}9,'�nG�,C�!}���'�c�ɿ���(&��ڶ] ��v1�VLќ�۝��*�Rs��&���k�@ǜ�hN�(�(�ش�4��Y�<`wg*�̂�FF�8�/>]�VF���K�y�4�Ce:u�J̩n����Ⱥ�R�wB76�h�m��-�m��	AK�t�,�ޣ0\dڙ�{Q��^S�Y���O���a�\-nf�Z�f��}��}�o*'�ﾯ/vj����z��������S�U�B,�pxI�.话�QR��+>�W���L�+�"kǻ�;س��E[u�a��|vґC5d#p�gF��f��S(\wm�M��D���m�ya3�Z<)W+hxM��t���[k���=D�Y�QcO�:�;Br�L�]��iч�6��Y.�Ԭ[����0��*̖��J�!�ݱz��v��i��_���u�13۽��[�S���CjNv�齜NO���s�:�ז�@��Mr�A���L��C˝v��ckvqwW�d�yz+����0����G�����yP2<��WΑ�7�V=��;��̛ݽ���g�S&�P9P����j���:���n�;GsV�����1�;�U��^![Hu`�ȡPP�.
��v����^�bu�/P��NV���o0��_���3K��Ns_�)��.���^�P�b�R�,T���o˫:ך�Wx�s��1t\����yN�)��7�[�W�LU�`�Zb�u��_D�hk�:�5O-����V�7ò���\y��Ah�[���}���:.��VR��v��d�n�@n��aʺns��8A�Z|s�zۮg�.Z�-Vk���̶����d�r�X3UYK����_Nؘ]�Y}����%5yO_R�UO�Tf�c����4�(�l>�nK�`��u�='DW
��{P�n�[5�|���0�l�u���纩��*�4�3u+��1��yDDJ�a.�{����WK&	�)U�{<�8dp��>U��.�Vg�.Rה]��|�i�G+^³J�v�X(B%�{ȍ3窖en���GYӺ�
}��"�����z�2��>"T�ү�ڜ��9Rj�5��89���.z�9L{`R�_jR��B'u�DJ���|sm�G��r�;��l�ǙFg�T�#8����/z4��7t �a����s����ޓ����:b����J�}ٓ�.�m��N��G���L𬒯�e|Дj��R�p*�����)Wf?/�	'���1�v�Qf�����P١a�����Gg���j�3c�*PLW\�o��'km��1�lU������8ɂq��@{2 ��pL|���p�HϒV�F'\$�|�: ��>Gh^dC�ԅ}�LV��P�hmD''�M���vd�k	��`;|���⎬)\�8����YbЛ}�z��x��j1Q��}����ܕk��*��\�¡�P��v���}W�4J��\ f�sA����sTX݊�/ؚ�s�����2�y�H�7{h��ʆ���7s��m��X�;���������ՍVvK}b:幰78�'Gs�� ;MN��.Y�N�^i��Gz�:iǽ���\С��r �N�s�����sOVCr��Rk
Z��*�Õz�֯k�0�ʂ��K(ԑ�f�}��p�dw��޻��mÆ���1ff����=�����
Ijx��z�͛��rݍ�i*F��t���v��[���n��h���+Y�T�{W�^��b���a�:��ϚG�z��&h�S	�M�� �_�8�wZ�z.ٸg;�`�N��u��`�%���K�d�;�m}Ö���Eg��Ҋ��N��ebd�Ѕ"i���X,���pUܜ᳔T���yu�^�l�.��**1ᨭ�e�glʳ�*$��v/��K�է*	c��$����v�Z&�,��m�`�N+X�M&�t�-�C�6����J� ��*�٧:���,e�2�Pv��b��oo{�����p��!�]��.��=�ʊ�`�l;�鮇1��k��dֳ�t��t��ne���w��;�
����.�*왇5�Wop
���]G�tU�h�!:S�<^i�w��:a�����Ʃ�Xvul�r:��w�*�q�M�i޻sq���5۔�5��݌p���ӵv->xOX�̍Ӏ���V��(&3�[��c�FV�a��wh���J J��f0`�Y R�IJ�,P������M�jYd��a2�6�%�#�� ���23v�r��B���A�ʉmIytj��e��k2�a�vl�V̒�5c㔔,!���
PJ�L����t��צ�X�è^�.���e;:��F���m��C�R�>�����6p7%��}�6P�ye�u��*�^LMK��	�������{�(����h��U�m���� ��9�+r��u�jW�T�,�b�b���54���t!���M5]YZˆ능�jw(�]�Z�r��N���#�Wus��T�l�ڮ+&�Xx+�$Je���CYwf�^�w�f(���A�ɠ�ۣm�0B��W�T�G����-�s�9�gq�?��5�sRt��q���#�jY�s�_pzx�i_]m,�	��i�yYڬu5��KrRS)������5�Hv�9�ƍ^6._vu���S�ԇDO�0�g$漒X���{r�V�v�*���4e�� x���;tTt�{E�g�]w	�5>�'=�X/����d�iV�c�C�NW�:��j�z�N�8y��l.�g[���x�YY%u.{9s��6	���Md��\c9��[�)�X�v�b;�w0X�uuuu~��mƑ-Z[h#m�\1�i[j�Zکm-�P[l�ʖ�-���T\���q��GZTWI�M�\�-Q�YU[ZQ�����\��T�\�m
ƊV�ժ4kn�a�����Qո�+l��uj��km�m��(ܰ�p��Ụ����%��l�q�!mE��ֶ�T(��
���Z2�ʲ�Qeq��YX4��3+E*(��G31�l�m+R�e�)Z�#F��lR���V�V�UkD�f\n6ҨҢ[cj�XV���������[aZ���Aj]�pU�DeB�������0R�l�R�VХ��V���U[i[KV,�1��W-f!e*ыwIr�`�T�++Q-�F6�kKH��D�Z��J�R��]�(��UX`%�(V%jFlAFūm�
���X�-e
��wc�� ɐ�Ll̷�[5�)�����R�]vM;X�IX6<	pR�����fp/�X��ӗ��cŽ�����'���>����abf���se�S��������#�S~(/K���N��y�S�ܩ;r���<i���z,���uĆ�ul�}�C�R����k��Z2����w���7
�/iENY�˪㹺���~�xp읮�_AG��O�&�vjua`A�iz�C\V�V]f�㴕�e��.��CT�^
�� ן��8�f�eB�A��9��Uᦚ��uA�ʵ��=s��^�D�Y/���t����l�������6ϝ�%B�v����W��u�:��B�%��Te�2]W>
���>�?ߜF�&�z�xSeYӑ�ȓ�Z��1I<=��YU�r��yQ��Q<��x���JZ����W��s�Z�̩��-�hY�j��k�$m�A�dTKU08l =�����H���u����r)zu��ܛCs�����l�(A¬��k�W'ǝ�P}}|&�,2�`�7n��@�Z�[�hz��G<�A�;g`mWM��19���/(L��
��i��5(�R��i�w�hk�d7��(w���07�[{����eV���U�ޗS334��k��Ѻu����C��a��%\�p��Q�D���إs�mԝ�rs[��������y-u�[˷�[]�lK���&ݪ�V�'�)v/m��u*�����E�:� � <ͧr�(���mg �U�^Tu�z��fS���0GR�
�}YtW�.YB�JS�{
"��y�z0wJwn�e-X�U*�ѽV��檝è��:�\>hI���4��7���\�;��x��^�~
�&6���*��B�[��۴C��u ��\�Y֣�3'�x�}���i^��ekF��Xg�]'7��B��"�e�@(�r�&�q��&�m��h��1���X�[��M��܈0���փ�*�=S�������QI��q���oY'c�l!S��u��P�r4��M�o�^�}��
��N�X�O[x����T5{�y�;��YR_��Ֆ%ݪ[|�%��1?�2�m���������gf�ɞW\�����o+<�	ڥ�_R�p��mʄ����O1:�������.`���7���w%�����{�0l�z���pRw��/�s<9.m8�+��aޞ�c/01NJ�Y��v�y�3����M�()�&�p!|]��s7��-�%ֳ�������7B�U�tz�t�lR��;7���]�m�j�tV��WV�v�p8�B�����}]�q��]�U�-Q#4'��עW}@��KH��qrho��}��(��ʝ(s&�L<|GMnVL/���3��e�:�Dֺp�t��n�#�UNG��04�V�|�h�8I�Ns����xW	��@b�K�QՀ 4r�ژ�tΘ��@�U�@k�o����|�2�����@���G�goЩF���ʂ�����
�AV��%�j駰�֫48����E������I�.�'s��I��O��'fj�s���@�IK9��B���jR�:��3<�j){�]qz�ʊDƿ2s�|�944��֞��l�׼�O�[&R]e��������ZS8<�]Q�mAS*_W�&p`j�"����C;cP�� f�
���j6���;w%��合0�eu�foL4k5fz��o��m[tJ}
E���L��$T�SGJ�(غ��*�Z��[�s�CdS���
�q��]VV����W�ND YBs
�N8O��yg�2�ИD�Ա��[���[���mOC�g�!C��@��4}�@���`�����2c� �L=!_�8\H�S\Җf�n����#O/����pp��s�����ӭ�m����W�Piw���sϒ�Ai^e�WEp�j�!��S��2�l�r�=v����������������q�����#yff(��t닍t�xe�kT��
p̚���n����q��Ճ���q���̊�]t�d[� T��P�뵳���:�.S�)���WKk�i]t����Bť�9�"������t������b��z�Y�A���@��r,R��HJ�g�T�������3�:M4x9�2$�����E����3��Ӣ�1)˺��`_Z�8,�|�#��ʱ�y�L^~�U�nors7_d^���޸`��ɬ޾ϑX^Tz�>Z6�%��$+G]y�^��%����u��{�;�y��R
g!��P3��u�1�녃¬{P�;��7gvO�����]����;0���՞oDm�Ҏ��xxXɝp�U�r{Q�BY���}>#��r���3CK�=�.�|mp�3��D�����v%�現N-��0�����I;t���-��Di�Ϊ�:O�*	P!���=���]h$:`��L0��7�X�vTߴ����;\�)� �U��R��Ta�*�Fi�~W����/}Z�#�ڇj��/Q���"ӆ�OyŚ�����~���	C�l"�}<	��t)���|·F���N��Ĺ}��S�;��W7�[R�TnTÃ��w'-�iV���:�����^�u��ƀOp�+��7)g{( M�&����S�T��o���=vo9k�c<^u$��;Z�V���o:��n�ʓ螊մ�*��������v����\e���mw&�Z�v�5�t���8��8 ��²:�U�P B����b���o���N�}���y�~k���������P�vl�LGf��B��.�8#��d��Y���LlO�����չǎmlf�4��N6�h��Uc��B8>ް�Ĉ����\mn�^�aU�&*<�����n���FPrr��*d�S=
�v�-X��ju�hmE9<)Q��^x�=��t�+ɪw/ԛֆ���[3��	��?��+�2�/�&(*�0R�jt��U5G��[�Iw���7}]�w�㙴=�~�Y�'[�>����򽤲:�(v��0,���d���4E�ɧ��>��옎'��x�^sö`�wE��?oR�N�%ZZ<������ָ��{
�X�bpgH�k�C��C�;\�wo��E(J,;�Ao�����>��ΥҜku]h�w�+ܤ.[',P���}����m�����⼵�B�|G{4��J]�g�NaPs�Ah��=��u��z�G���E�tW)՜������v��`��ɺ��:�������zt�x�i�h�v�V8��7[���T�X��M9la��!���b�R��D�:����
y� �ft�)p5�˚�G��a�Ʈ�-=s�wM6�\⯅��kKhS��{a�[+w���g6����=�4<�����?h�Aw�F��ܾ��8�>�+�S��uz�:wgi]E�vd�[&n�V#�"ʱ�ӣbj"� �����H��,��ܢ0�Sn����<���t�b���9x:���aD��c�*�|R�2�̤:M�n��_�Q�ǽ�n���ę����Lr����B�N`�r���33<+�3<l ��ia'X 9�e��r�]r}���
}�B|-ܲ�v�K��/>�҅ԧD�H*X�HGf��:\���/Z��5o���S^�������K,=��3�ʔ���j�a��BXb����Ud��xE/Vv;̓R=\t�ǩ
a�咺V�F=�PU�\���4�D�!��檢���z��u2�{7��]�bƋ'������ �[A�����$�z*������ĝ}�sw�����n3
�]�������^s�ϝХ'#kҬ3�8+<]������ǆ�%$�<��:������n0�.&1���<�͕۷�mא��{"�,ڗ�,����uv#�|�DrT�7+v�vj��s��P#��07�2�_sGr+/S��5p{�*CZ�X�b���W.Ɔۗ����:�S��Mdw�T��+���?J���R}m��$����,��9*�+r��ΟP��g#&U�PnnfG�X��K��5�	��Q����S ����	o6�	�Y��y	oj�<h����������AAo�R�8_R.�mʄ�F��xLN�\����0#���A�h��b��|�Y�����rz�d�Y�������3�b2ݧ*!ıbˮ	@K�+UG6��N��`�O�
u���E��K�N�R�춸�Y�����W�2��|W�{Ÿ�d���]�������p;u|6*)}�V]�UUu? {u�1_n]qw�������<D�O���.R����`d�e�]}�ܬR�k���l��:��r��2+m5#'1I���vu���z���x-N�>�<G�H]jw0طa��}r���9j��i���ij��O�.�>Z$�k��7��#ը��u�����*ٔ��1�mR;��oX�S�]��&/It�Ye|��Z���Y�3�R_���j
h����]%{Ǹ���P��@9\�X��/X}w�m|�B�j�F���oYFݦ�罗�9���#��[i�ӂ���1y��ݮ�9�5c�<���v:P;��k���ul繃T��<}>���PI�r�j�1���j��r_Bt�(v�u����xE2��w5���A]��dؗ���s�M1yG�-����7��C�ޟc���g�֯-a�]~��is�pڧ]��Ć��i͏�P� �,~��t�o�XE�
U\��ᴎڢ�j�][��0�`�zn=�v�RF|���+�8�>��x�	��/�Vd�H`>��$�^��=�]��u�Z���w]�0sCjd�,^q"O_���ݶk�] j�bUy̪�� �� m�xe��JT�=�XK��)�#��8��\qy��{Z5]�sW�aHV�gs���T�q.�E�H��Z/�Z2�����p�33��}б�S��Z[�Z}Mfw��}<ָ���m,���O ��݉^�"��F�pWR�JK�^��G���h��z�:�$k��/{t���X)�S��D������pY��b�Pr�� �"�����M�:��qL���C�������z}+�Yu{�B�ΗPtN8;^f��	��-��+zP�:8���^��3�}�R
m�>�A2���Z����p�xW�����tW[���
�ꜷ*�K�H1g��>����֙g���4�^ԍ[�{��.i�~
�`�*p�Q�B����Ox,��[����(R�o����4)���?vsYkU��)OG׫cY���}�&�q3�r叟MOU��^�q�w9-+��t��}h;Rb��v��AYSF�юn�2[���kg=��ЂK��ʧ��Y*�c��{=d�g�L�#�U����u���(\'�rm�x�-Sw*UB�k4:�߬/��!��ɗ27�,D[�.ޮ'w՘*\��gH��J`�����Aݫeė��A�[cmU�]Ռ	�EKB3[DM
�����#��/�2�ʹ���#���u���`�q��W���YAIꢀ���:��|��Gj�ۭ��+��=�O�x����l��dA�!d�A�֠�!S~�$WZ�`�M���Zg+�8D��������;}yWV����`֍(d���A��_z�d��^�N5�Zb'%�asٛ� �)��B�����Z�0m�T�9�T�%BБv���̉����75��+���]^.t��s��ohP�	Z�h{ԅ�YLW��u���+����MK�OB"c}�IƝ�\��ݮ�>��>�j�|�Pe@bLPP��Q*vӍ�esg�3;Q(d�q;O�g��C&��+��������3P�y���k��n�'�kR��8-$�{״�T�š��Ṕ;\�R�V��+;�)���{�ņ����U�wQ_m�-À�]R4G+��_	`rK��|gN63F�B	����xXt�'X�h�b5�e��Q�gRSƩ����Y�5y,�
�.����i^�$�:���.��z燂��J_5���!t����a*ô��/ϯ�W�&���{6��j�aމ��S�~Ί�pv���O����H1����B��6����4:*�"��RJ�f�sJ��Ri:P��K�C�s|'�ˉ銠��t>�^ .�pu��+�}�E��x�t����y,�u�+%^�2��j����J�|�*����v�r4��Ǣ����eOe��v���a�d9����ζZd#^���'"5��0�z��(+��$_3{[7�����ϳĩ��^FCuc�2��EuAUCE:�Q@�S2�W=.Ff��1�Y|�|��K�6e�y�2�� �:�kr%�{YV3�����)�b݃]�+��!�ל\�y�V��
��.R�|�x�+�N`d�yB`��
�Y�̣P�)[�/�����L�9�y����T�Q�Y�#�������Y%@c��E=��uA�~�u Й�Nj��,+oӥ�|gfV*�v~t�΄]aj�B�W���sUQKT����Pa�Z�Pⴞ�ߘ�F��]2	�K���w��I�4�%��
K�AN��`H��SHЦ.�W`b�*=�9����Uw���+��6iu�t�#������
ڬ������ HH3�"fʓ��9PX�mL�|���.�k��@�j���z��e�vg5���1��:�枍�n�a�j����!��Jh7F�FD�䱫,w]�s�[h��H4yQE՜'����ab����E������"�d�U���V��ۺv:]��b�:��K����t�ӕܪv��o�	ي�7b�Ϙ�6���o�qeaGv��u���Ԛ�U֍�3��+�ؾS%�����2�sJ����;�k3T]̓lhɕ���Y�r5���CBy���:�Z���
�˵"�]p��P�WC��s�5mM.Ѵl�D>ʼ�Æ�O쬾r�y����E�u�G+��^�ReeZ��Wq�O��1u�Ix���8���a����7`=:���O3k�ܬ�����v�a2���G��CX_ʙ��]��g/ ;n5DP��x��z�.�v̗�����-���+��!�8iVw��<�o�k{���Ȯ��o�Ğĳo�H6�fE�k���7i���tF��5���7D窛��ݛB��]:�⼸���$yI��b[�*`<�`�b�K9Z�Y����Q}��2�<�|QNf�+���am�k��^P��u\��C!\� v�Q<���W�f5w{W�Qt�+�M�T���Y�5��HK���uǶX�*��9V]�B�Jғ�-e�M�!�E��aF�@A�0n��&<�a��w]���6���:�tj�5��Q^����/3+^҇
�B8�=Z����+v��̱f<ldf`Pc ]Z�S��r�^;4Fm�d�\�6�"2�lĩ��w��U�(sVI��^��;Gm5��d��R��o�X�����vw[��C1!��t����M��h�Dj,;�eo1�2�"v�R�T�����謟gSS:F�.Dh˳�(2�������Y��)�Y�������VD9u-����T:�Ý��v��q�n���f:��Fq�ۉ�v���R�X��f�R!M��^�������p��-WS�4��b���oe:��Ļ�:k�me���h`�]�
�@21:ꂍ�9���2N��ᬻ�+���%T�Ruέ�)vF��d��N��w��-II�d|�R��SV9�����C�llҩ��(-8N���p��5�熻R���iX�i�v�s@��I�D��W"���b؍y9e�G��?D��>��(�h�k9����u��ٷ�b��е�Fn`5c�ɥ=\����ähc��W�in���cw���S�
�Y�-�Q*�։V�Jh���֤F1�����Q4%,��+X�e*V��TE��������������c[a�.4�������W�2��Ҷ�+DQ�KV��R�"�Z6�"�Q�������
��"*�kJ#ik[jT)mQ3mݮ��U��Uh�Y)m�TEUUVڠ�%�b�]f*��JJ�勖��2�Pe,��Ե�ikD�F�ڭ)B���U\-��"1]�D��D��Z�F�V��1*QkDkc-C+t�9h�E��UJ ��aV��5*[A����KT����"�����j*Ц�F#���50Qe��TQ%�*-���V���*+m��ֵb*ֈ���R�kP-(��(���"��̲�J�[lQ[b����J���V*��U��R���6�m�U���mB�Fm�4��.U���:L�jm��DL���!�a���f��N��5i�;�u�Ŗ��;g]���2I�n��Z��W5�澆��n��]���5VP{V"��-����J�����f�!�������S'JeL�ׅN{��z/D�~��C�PK`o����]���A��������ߝe�^U��1��ٻ����GWmWU�zid�z���=��׎O�ȃ�h8�e5���^�
��{��xXZ�X��㸸x(M?�{qܧ11ϱ�����/JMZ�>�����++7�1F3�����Eh���S \+��Tq����@�sJ���'��w�s��;��X7׆-���!�_V3	}��	����G��vN�F���4f�ǹ����g�v�C����PvpR���/���.�e��.VQ���ӷyJ*��d輫���L���3�ۢ���riW��)GSP���tw�;w�[�H���>��=C��[��׶��
{s�t	mu\�^:�hT���n��=L#c����dw3=�oH�3�%�����P׃�x���C,�v���*Q�6}r��%�{va���WS�,
-2��[�ր��j�DYu���-F�J�k*�J��7�ˢ"��J�+B�	 �t�9�1ʌ������V���E΢�B5��Ճ���xEʞ�56Y�n���]7Pa͂�8{�&B߈�v �!pp�/�W�xv�]�V��Wp$��/�k;����,�±���È�M�t���S�²+�l~��u��2��ˢ>�<9ʇtT�����S&�&�Vg6��Jz`����vTG�T�`Zgϖ�(�z���5ck��8-��`�R�4�~s���� 0��{�Ƙ���//�U�h<��.�]g����'1�m3�՟7�A��J��n��\IO┠42�(ŀ6�����.�l<|v�R!k5d#��e獃������955���p���t�JFr�9�u~�(\�B��]J�giϳ��z��͏x�g�Z��1��+r�:�{b�4;�.�M8Ot���6�����.:fK���˞w���׊Z٫t������.R�o�@u�P�����긽�y�fH�(+�EHHfـ�ݪ
�c��+h1!�C鼪C.��WN���h0��^��z�4������Pḫ����	����)g'Feӡ�5VO�����O�
�Y����z��e����R���3hB�Jf�`j�n	������A�O�}�-F r�AW�]�O�<��������K�ŧo��1�v7٧=���5��͉���ȶ�N�8�un`����;q8)
��4��Z�x�)�*ipQG����t��N�^�Z�ᱠh���M׳��}�/��i����x��M�#C�<��-ȶ��������:#C�s�x�E1lqw��ڵ@\�U�YR߯��q��;3x��Uf)$J��S��*Rs�*�7�kx��LU��[���1�L���e��y�*���&y�v�S2�^�I{]b'z<��_��Ay����JxU�&�N��gw&<8d�m��:k�'�t<qp�p��s|",h��l>���Ƙ�FE�|U�s�}V�Vu�@�-w<����L�}a�xW���N�Ve.*�'Q�18��������=�-����KK�)l�4��I�5E��ïk���>�`K��4q�.mVU�=!(�^��=V�<�&�~�*n���`N-��tP�.�A��D�����-m�N%�\�k�����ᚫu�K��T.��x8ӹ�UK�����O%��x|��ϒ�|�i��fͻ�m�C��d��l��(��!d���`��
^�V|���������:�xL��L��P��b�j�t�qJϷ֡���ȟv��{S��v�C�)��d:Ʋ�#�K���%��zw��z�|H���t�����;9/l���"ZX}~h˭���T�[�*�I���Q�@58�H�%]�"r�Ս#��o[��t�kkvj�1:�7:�o[]�X[��<��,��i����N�2���:��g��O��{9tO"pI�e~��;�A1^9�T�=(\E�¬��0���`;�B���m��9���B��,Os��Q��{-��@/��GA.U��Al�u��C�qV;jj�}n�W�b�:�;E�;赑�=�n�{��5{�[���-�&� ���C��]�<G�s���1�c��U��A��%3�z��7���N�b�{wf�yԴ_�xg�S�린8(�/::�1�i�
\���F�k�tU:�a�3J��<�����0M�m�d�8�Q�F���P�3GPްѼ����hecC;K��[p7|��w�[�|�B��6ĹA�ǆ�gp{���{��t/�P�W}N�D�b��zV*����]���ð���]:��Oy�3�ٽ3��t" ���P�Z�?�7�S~k��+/�u�hB&��v��x//�=�ڐ�N�M��s��>1
�ж<z�&ҹ�A�N;�]��2���TG��$���ٯ�=� ���s*f���
�AnȨ19����h�����bB	d̵n�9�Վ�m �� ~���̪��
�m`e���]Y��W�d���{%��x�wtו�+Ljf�pJլ�E�]~��j���k��]6�����܎�:�j��smh��m7��{h� ��s�,L"]��:��]�,u�Tx[lԸcu|��~��Y��{+�|=��d�3Q�9K*�2��*��LM1����vɋ�d���5��Q��t�#3�[�19���/(L�Q��c�jT�q�²M#���\&��͎�dI�r��E/�-E���^��}ڼ>b��R�
�[݋m�	�s�v��S]���uU�9�9�4Q؝��!��c�H Ź>�c�����;wSt6��at�K��f�Vt^�4(�u�@[�2��>=q�
�*��:�!*&��mn��mܢ�֕���ofj��8ް5��f�`3/DŊ�'`Mz#B�ƪ�=��4����ej��K1��E�OEH�v^[
��E/�/a���j)��U��o6W���A��&n!1�B�J��hR�hW��-֗byg�k%�X0B����W��9\�Tj��G�9��e߸B��
]�#s� \61������2��é��:�^��W����g��^�u���]w�ru�ZU����[��S��imH>�`z�A��,_R�p��r�(F��{�Թi�e�?!����~�W|R�+��S���g0��z��pb"���PC���y���%�傌dXe`>����M�/9F�d��-��ni�鏐8�92��\v�P�9��q˿�+	��]��Է+M���!�L1��u�J�CJp�gze���*��
U'd�l���w/�d޺)���s��Z��/y�כ[>�n��}Z��8�;:�d�Z,�+ ��1�%���iX���"��l]��n4����������vdf���s�z(w���HP�j������ia�Y���kӌ�M�-��)����ӎ�覇_Cb�R��S;U]�WG�N�Nkp�2��C����͹��(kι�$g�XVRv���ЧF�|es����5�_am��'<�) ��P�_PT�딾�FTȺ!�<9��wqC=���]=��ӫ��\�[Ҡ̿�a�ٕ��ڶqK��C������QK��8-�VN�9�j��5����7��Z��T��J�C�:K��u�n��j��x֔�)Lm	�'��#�����9x���^�
��V
��UR\�,�/4��|v�R!hf��X��þ��}8W��m[�w#�{��5)���r�9�p��rĠ�]ԭz���J�x:a��v���L��Oib�[�-��1͠aS�WHT��W����*�Z*a�_pI�����²O��au�3RJ&˥��!�g��z�kG�4ϼdq ���z��.���wls���zmU��y�Cmԩ5��&.��>�Lܧmrc��Q�2���6ź��5�LN�(	�����	���������m-��L\-�q&3�8;�cC[�p��:��kC��u�ri�nZ�~*i���4_���U�@�,�e��;��v���XX���(���s=N-mX��V���.��O��M�y���X4���f�P�Ko��<o�����^<��ѫ8����8&��1hpp+;v%�<1Cl�]�~̮�v	�Z@m�����3/��Tr<�w�6��y����u^	�Jx"T���x��/U�~�U��j5�OM���P����������&DJA�x%xLK�ߛN�	����upU��]����̕��o����˺��ԃ�&;^wT��\����}.�X�;2����D�5���Ә[�>�xU3��®T����cGF�D�xX���!N��f�E{�:���U<mzoO8-#�>^J�?�l����$�r���yה�ð�8���q����U����f�\v���J��-�`��(_�hX��u�Ax��<�J��ʩ���9(G�v�.fU����.�^=���!���(�Y[4I�׊��xEҋ;���k�u�; o��(j�a�J)\�,t�\;�u��`�+��/Z��gTUg�κ��w�j�&����z�bj�YԟD����Y�[a�}����zs�Um�ظ����^>P��;�r!z��2��>8$�^n_�ƄӢ�����" �D̾���OI�}�0�~o���V�����^�C�����K²�>�('�M�u����u��h��Ҟ"�g:=�D�^Q���� ���5�D/��,��GR/
�겚�P��%�^C^{���jr��B4B�5���8o��K���Ҁ�vh_�0��m�9�$uF�oSԶb�[(��慈��*o���q�rcX�1�0������<Z������e�и=����'2��������#����vJ(77*�@�Y�4�W�.ǉ,-<���ݮ0X�v��VMCյ�5o���5��O^��	��:��i��	�*���8�gt�y+�{���p�|N	��3՟	�z�	��J��81�x;�}H_Z�<���R���Ù����3�`�:�˒��Nf�:���]YWq��h;Լ��<��N�f��}�W4���.�^өhu<��wωw�N�c��k�9Ϊ���j��S
f{-5xUu�s���7y�$�q��o�.|��K*������N[�Љ{h�u�+�Y%APb����J������x̮��K:T#q�*��ib�;��8���j���B�+�7��+�B��|�b��C�q�KiR�p�����x1e���2v�����6뮽�ڛP�6�0<.���K���Q2_�
�^1o��U��9�[UΡ/D�V�N7�U����6��V;�G�w:|MA�RiO���|���j.��UX
�\X�e�f�s��_	�������� ��)��t̬�3ۮ��&r{�̍�s��g��E��9c݁��+��r��rEC�'���D���h�<U����Ȼ>}O:FU¥��ϡ�>㘜�����I����,��� ���:E�½���y����|t7C[�֥(�6i��{�1S:�p��jj/VU�Լ�0戕Ѩ0]�b����бr�ʯC)���5p��tUǂ�O���v�̸n?D����,z��`Y����h�1�U�q��?Y�1յ��=�v:\��Ylgs��D�T��UQ�	�s����Ԟ�e�Up�Ҫo& ������0�<=W�6�Fs���'�:0��
�N���m/V29V��pl�-��v�[�/_���/��kM����_e�bg@8|R�y@U�E`�i�>��ș��wA��6�\��9��B'��VtD��њ�)+�v>�Pٗ΂��]��f%�$p��Ԟ��䂖Q���E���s�i�b�E@�,\K���K<ZF$����{)��W^�L�U��T�E9<*�Ny����T��G
Ң�zN*5���+�6�19׽�i�RXӭ��=��Y�r��6�U�5��M�5��랃�Wz����b��)�Z�m���=KD������谋�/{Ǚ��K�4��s���m^���~̈́Gh��⅝G!�˭R�/�}��/>ە	Cѡ�}�TyR��#��7����QS�/�~�����9Q�f �v��|�B��A}K�v�u`���'�^��\���l�0����؝O_'�+�K��_�6诎�]<��X��)}C���~j��z[��$�y*��L��Nq��]����JgD���z�ukb�R����_�V��%�����UU>'j"�J�vg�\c�P׃�x��Y�Z6�(�jjٍ�]+$f�4��ѯ7ՠ�S.+���\����5�ʔ�-�����a=&`�F%��ր�B.��c'�Ml�;Wf�7������l�?�l-gQ���W�XX=��k�ΎEj�$�]j�&��Z`��ƻT�/ӳ�� ��H�GK�wZ�u�f�K.��޹R��[M)n)Pi&u�(�ŏ(*L�:ͼ�"�����;�}��]#�	�u�rPi��nl$Xf�Ul�
Է�I5��-�X�����9j�U�"W�����g8���/'^�\T����i��yk�-�P��d�/踪��Lbv+)��s��d|Xͻ�nw^^
�^�b��,�B�]���=�'Y�ܥ
����퀂.�tsP���8N���nr�ZT��e��m�F�9b�������Yڌ=���E�+�%�C�#��'k��x\�;w�r��*���0P��ڋM�6�r��(�Wf�%�RA����ê]���`ă�.@ ����2T��!�X/4[��*�w�K�7Q��Nt�9y�jI�6��,寭�A�G�@�p�A<���/��+B.�`�����Sf���u�B�B���!R�wt3���enGٲ$s6�ZAa�k���Z�D<���B� �H���q�������9%@�AB����ՊW0b��q��ES]j5�ޮ\����{4�`t��\�-0��r���
:i.��*S��j���0��cK 6��Wgf%8��pc�#��.��2���Y�\o%i��P�������`}A�{��Le(���L���^c�>e��cj7G���e�gܜ:����iV�=�H̗C%Mx�u[6B�� ��j�r�ʕ+��F�a�Nq�H,?v�X�d̸��K����ç�Ot
�R�ڢƹ5���@<�Y+'R&9/NV�˙���ٔ�E����_�1`m�޽{�WܸR��yœ�EOqM��T�bܬ���f��>z�l���xц��ǩwΎR�aW��ĵ(�ok�x������ս����_r�{MNã�.$���o�L���2��bviN)*ܝ����]p�(_���Ya����.&�W(��P�+��@ZS��F����B����<`�|�%p��ѫݧ�&��̣��X���V�J��sM�&��a�:�3��	w�:>�v]�/�֮ �ɶ���G�_] �
$Of^v�#��+&�e������єN:7�Y�9�OZDN@� :��e�40������.��ӈ'c���K[�hhy�uy�5ؖ�H7�`W������U����:{)��K�-�ox��:n�>9��6�*(���#E�M���˳L�e6���^��ˊ�S��Gt�5Q��]1Jܫ�;��t�S�iB���o������ }_J�,�o�H��̲D���wkqK]*bޙ&. ,��'K&����a:�:�q�n7�I���ӭ�9���V�#��O��#�qdf�{q.a�-;
��%�����S�u����Ԕ��xr+�����}�p�j�E�栂"���(")1�,E�J�U���V6ʃ*W��m�Ŋ��Z%����`���1��J���m�EX��ň��mj�(���-�AeJ1b�EF�DTQZւ(�"*�T�iV ��-ULJ�̪�Q�Y�!iX�,UU�b"#-(1Q
ܲ��q�e�����V#-���KV��b*�+-*+ib�eĪ�Um�*6ب���ֈ�QU�*t��U�[��"�-�Ҋ"��DQT��"�jX�DE2���"6¨-Ԣ�X�*����U��Ҷ��FʣZF(�EEU����Ꙓ��DQ�k���jւ�q*�"(�6�F ������KE��m�G����DX�X�������f��b+m��J(�Ɣ��V�DQb(�,R[`���E�
��*��Z��"*��($Qb�����r�؋Z�l���U&���B�+iej���ߏ�dz�%+��۷����gT�*�k>��Κ3��7���.�m��gqhoF8M����f��xV�-�3�F-��vs4X����̊4�|
�u']�p�%��u�W�_U��!�ZS#,��Y�;r���Or�L�t�օ Ö, ���u'^���])-8��E{|�����'ƺ��t���p:�K� �����H��0ѩLT�3���_�� ���X/ײ���L�lg��/s§u�z-�ε^Ԅ�z���(8eL޸��d	�[!=���s8.��".�3�;��yJ�����|���hA�sCjgӚ�����S��v��{���^.oG���@�����ZN�F��a����7��8p�WU+ͳ�N�ˌ�������6�w���2h�g���8(zͩV+b���&GNoU��x�Ξ����K3h 9�uӭ��cd[J!yOA���B�!+�ES4����;t����I���X��w�p~��s$h�Y���c��F͵�9�u���1��a���Q7�*%,P��P�O���M�g6�ש�eKے�M^�WVu���o\1��rh�q�G��s��j���-Y�e���do��Y9hzo>���i��V���}\���[jXDJ���m#eu��¸�괯:�f��R��а��2�×(��pq�f�x8��N.!JQt=��;:u��	`}O�rj�8�F��A�b�Ov��r9�(f�.��z�	z��%�/9�Q��O5D��'C�W���c��t�#�]�X��G��'`XU������cɜ�;M�ׂY�:�!`�2�C�n�!�'X,��x��0�a�7"�r���Xu��O;s���VA�V.�kN;�Ew�lyj|L�׶Ї���?	���u��m��vo`��)��z�4�C=I\8'���9�����M�D`��_�I�]�fR�1��zj����y/t�h�FW�4�涜���
�
ςqmX�Ӣ��.�_;��%��'j��d,U�Yo/���i�)�L"U<imL���J�R6:�j�t�x�Es�=���Kz9^��Z�O|-����u]\��ĮQ�^�������!s�Y.1bp�ׅd�~�8|�����_I�ޭ��^p4jbemf��5���(�]f�u��P��Y�gh[�!u��2��k�1jH���|�Ǘv��D.6O���xk�U,���<���Lt�A��y�+k�!f�n�jz.�/<�Z�m�=[���7��.�g�r8"���Fh7.[���F�@�>b��P�C<�-ԋEƌ�r8ӡi9�|����:��5�
LEW��-���RwR�۳��
�B��n\K��4�E�u����֠��St�z�zElX&�_3z�dk)Ȳ�S��L����x�o�i�+E�=N-s������>��z�r�t̶�T����MCյ��[�sw��G)_�d>GQ
���}�݅��<���W�c�j����>�mHG3��s^��un��^׷�s�ޗ*&_���W �wp�Eas�r����
���!�C3J�&9�Z:zB��X���ב�Y|��l�����p�(�갠��G.+D�@F�Op����Q����&9���I�x4��'ʾ��\!��v��s�v����[�'Y��d�c]�\��"�T��^t^�i��0�������	d�!Ј���/O�`��HcIх3;z)���X��6v�G��btΔّp��B��Գ�Z&/}a#֙׮bC4��S5���	����0��/3C�trt(�Kfs�Z��2���۫Y�*�� ��;OB�4޻+�y���Q�w�j(������&���6f-�N\��Ȩ1�\�Z���@��g�����ɰ-�5��Q@�t�z�<��s�8.^P�*%��L����4�	ҽݱt�:����S�޳ڤ�'���X	����h6���f[>[ӕ�ht����^_c��{:Ɉ�]yqd�䈵�����
�����7�ҝ����5����G�ȉAH�j��W_[��'ww�c�Z��Sj�k}�jt/��V���6 ^[F����`時�п��YV}�u�o"��fS�2M�M̤aE�22�yT��J�hM��<�0+6��[��Z�o�u�ҩ-�n�,geJP��P���V���s��W�mU6C4
��T��.����tӐ�P��T�7��c�Kt�c�4��&�E�v"�4�G��M�Pg5U�rxP�^��Ί�O<�+�� �md==���>��8���S���>YK�-��u�'��i9p�x`ok�ld<�͔�� �)�5ڱ���YXRS5����3~��9���U[�:ux��:�+R�T�n�o-�M"�u��f�ݷ��F�_`��)�_�։�o�R�_d�)}�UHy^���-ԧ<"�ѧ��K���`�j�g\eI�
��yx�gQ�|Z������%��r�8.d��6P$s'0���j8kz�r�>�7��r�2�g���!W�;:)Y�V8�[���T	��:Q�ީΙ������r����Lv=2�w�dۢ�0S���ѧ��R�7���}�m`�Zv��a�n���q�=�B�ˋ���RƲ,�w^�i�9�#H���AD����L��GX���Ú����4���u���"�!ꚦT���ޥ\�*�2��/Ju1RZU�؅�r� ��r���ڳL��u`���q)h|�PjNZΊ��)�v�p>K��oxs�T1�y�Y��s+�U�6*�ϰFEAY�f�p�k�3��"R��v}k�it=��1�
�	��o���L''��;�������yF������#;r1���pst���5:p�XCt���}��]��r��.��G���>2���/j�ϔ���
����2��l&*n�i�dl��i�ͬ�.�J�,Z�1}LA��r�ش��Au�P
_U�{]x�5��&w�Uj�޷V�����]$���_;��/�°C+�T������:�&*薜N}��ڽ�)d��g�f�KP�����j��s��ȗ��O�
B��"���b�Q��G�GEln�k�<U�]�4'��X�B0o��z���"su�	��P�)r���rwYZ��w]��v��C�/�
�%��C.!+c+v���q7	�P�>��ϧ5�HGf�/�{���ykI��bٕ�����R��M�b�'x
��)���(%������v�Zc��ĨPwwR��y$�2a�H��:�SwU�U+��.�ע��Hݵ�"��c��&)�R�F�:��T������}Ϙz�g�]F��-��6�ᫍ�X*f
��IS���u*{O��)Xi�V*�Q,8��F�;�Y�^�����z�q��pq��W�S��+�;A3�P��
EՃ��ON0v������zb]�;�p���`�;�JP�ӓ���r~=^�Ҋ����,n�'��+ -�J��պ�׳)���m9���'1:����΍�#�9�͊��%\]I=�|�tU`�f�H��Mm��(�_y�J�'[7��X�{�w�o6<us�	Ng��H1�)�'^�>;ټ!��V�tyh��%��HV���=Lv���_��b�;��N�{]�^�x�)�S���Tr�R��~Tv��������>1���l>�]J�wn���x���od�$�q�Ʊ���d��>���_
����Nr�>�r�����!��<�wr�Ô�5�F?Ob�d�����I�0�<0�P�1Q]��&z��i����2�ڷ��n�1��~+�q!׫4������>�(���9{Vi�R��v�`�kP�,�H�6��U&�h�b�:�֡�<j��郎|Z�2�J�J�a�xbR��x� ��Y+q��,v	4�}zs�Y�i�5�h#G^��S���n�c�;V����R(�H��\�{*��B�]l��	�`D'a]N�}`�I��2�����l�oR:�S��^����v�n��v���/�BV�7VM�:�=��1�����8����u�^;k��KP�]�G,i.1buF�+K�F��0ٛM�&���1z�Xk�J�Ph7�
)WK7��Z�{�(�Y�vEm(o�<WWA"���9��C+)z���'ٮPᜁ��JlMV-�u43N�^�P�ڦ'�"�-ݺ�j/9�I�ہVW�o*��hcz�H�=[��#���x;�7�x�8*NU�Qv�{���3���3���;4�*�r��`wo�Slez��[����t�ڲ4 �U��Yy����N����@���7;�<�_�N|��9෨��ko����o�}��]�U�6C�)�7dJ�ּv����u!������)�C	��V �<��к|GT4�a"��Z��`�S��)���!ߪua`A�hl�ˠ#UWp���乆85����Aw&�.��m�[S���t:����ONv���S��'FK�
�/>�S|Vٸ�����w���.�U���_�78�>wl��!ЈD
D�7@��9�S%Ձ�[���ö�X�7^J����[1 ��:�C�vӫoa��5�v����W���r���'f�(��v�ם��O�LZ�|h������D�w�˒Ѻ4��Y�l;!Yl2Q|�X۽�_Q�ݵ0ݳ��So8 �smU��N!�=���^b���5���Plݘ�u�����?xP�zQ�Kw�r���z�A�9j���tYL����#ȇ�ń��בRZ�eJ7�S�{�=��"�W>y�{2��c��xl�5	K;7]-+~\�ug�E�"K�E9j�9L:J��r����3b\�*X�4X;㡱�5�IߣZT��T��ϣx� <6�ڍe^Ϋ�T3�G�)*�����i|.�1KL�w�hz�W����s�/<
$����G�����}��d!.�A�.]}ҁ�7��M�C~���>�Ih�2��E�|u�_�b�1��)V�s���o�gm߶��* *_UP���>�uF�M8#5}r�p��}�82]�v)TS|K���kY煎�/L��d>��TF��h���d��U@���_o\A��($�:��4�k�qx%2�̮����U��>�����ly��, ���*�H��Iw�����ݒg5�=�%or�D��4�V�(C�a����+��
�V
P-t�t����X�(G���dL�糤�SHΞ��j�B]�Ї�h�uqKΦ�[%��W{r�@�#\��6	!Z���X��g(�H�t�n^��3����]6����(_p�Mh�s�*�,�����q��+�D���u^7��K�W'���&˚��������łz�8���Pɋ�mh�����E�ݶ�X��!ʕ)�B5c_�tƘ�r�:�S�a\c��6�38����u-�����p�'w��3��c�7��S���sZ6��̳v9ر��%
vvٙ�7�Lg���7�3�cqZ�&tp�;	�0A]L<����W{f`�|JJ�U���	���\�W�3˴�(mK	�-�%�����k�0Uɽ�f{W֊��cy�/j��]i�n�{� hp���ՀO�3��箻)Ƿ��
���x����XB%Y��7��q�Q�=>�J	��^�9V�*G�ҭFT��W�Z�8y��tj\;��3�LNJ<֫��7w0]_��	��R}r���r���E԰�D.��0��O"�5�9<n��~���<���HC�	ܠE&��+����.�u�R��gn�"J�G
/]�}�ٝg��Uq^�e$y����L��xT�YUZ��([		�u�a��(wA��qq��Ch���+��^��ݛ�i�;%#t�Ně�f�����):[�g��00�3V��{DtM�k�T��	���g��qc���\�����{�P�k�y�1�R�vձ�=;i��#;:�.P�wP��I�ѻ5ؼ�t�=��p��rq4Znv��i�3O
ۡ�)�G�9�,�ʂ����*:�U�.T���C65������f�P���놚��	�V��䄭��X��'0����Ļc_B�+z�	9�{����g��y�	�a��B��j�J� i�x����!��\pfcB��i췗�钔[��:OCf����v7c����R����p������e5�y<�ń 졮#��Ư=�*֍WJɅqi�Z8)���(tmh�?I�J��r��9Nt�L��Ks�hEy���^�зy��莸��br�{�����G:\�d�j�K�p#�����e�V��^���Khm`��r>�Uf-�*�њ	pU�J-m�Ojq�H��/mxR���c�
�����d��-ק���Ԭ�	X%��X�d�V�@0ާ��k��|�7Z���yC�.Q}Qa�����zD�~f��<5��6�n��Vƻ�M6��^q���ͷ���aъ�P_UΎ��zމT�6Mg��v��$��	!I����$��	!I`IO���$�$�	'���$��	!I��B���IO�@�$����$�	!I`IOB����$��	!I��IO�H@�P$�	'��$ I?@�$��1AY&SY� Π�Y�pP��3'� bJ���"GX����5��@�U**Q�����dkTk$[2��H	V�DU5�m��[dCf���V�l�RR�R�%Z��$�fQ�J�i��im&��_X]���՟wB��j�1UE��fյd�Ɓ���&�k*�R[SH�ٶ�mV�M��F[klm��{�^�qK�Y��mV��j��)XjF�Um*�֖hؑ�U���Uhٕ��[h�h>�u���b�m������Z��v�-�bٲ�e�id�f�kVi�Ѿ�]k-�S#clπ  wW�(��n�U .Wnѡ��C��>���-�A^�\�m[mQ���[m�[ON�+l)�6նŰ5���m���N�H��ҋm�#j�QC�  ����Z3����K������ҟs����uzĴ�:�v����Asyr(�5�#�w��BT�=K�V�B�-֧-
h;��4�l=e[�եjD�M�J��(��mn���  �W�\444@7}^�(z=
 ׏x�CCB� ��W��B�
  P�xP�@  ��^�� P�B����y���hP�B�h{;����������US(�
Z���a��֍j֘jڶ������  ������}�5Ώn�Z�V�j�p��W��a�^ロ����oR�T�[ziN��J�ԅe����T��c�֮:R�����PQ��֦mj�X(u�l�V��  ���*[2`*hT��ݠ
���j�o���lV��:�u��z9�MS�t�f��旜�P���{ޔ����ݻSA�ܫ�c��f#-Vm��L��_   ��\�:�_sv��Р%]�uz8�C��.:zu�]Sn�ׂ���hN��Wn��m�EU!�w#l��h��$E���H��wU�S$;�J�ј���  w<t�m���wR&�+[wvv6S�R5Gmr��հ�=��oS����Wv�s�5�{�g:/ev�=��-�L�ͺ��کQ�6�VlhQY^Νd�ճj��   }����4j�wnδ��T�  ڕ�(kwlq��z3��Vc�P��w8�QC� ;]�׬��icjJ�M�i��M�   	� ���� wu k��:�;��-S i���θ� �v� �u�ʡCL��҅�����Uk/�  wo�:ʻ��6��:(,cJ 7v�P��:� ۺ�� Z��]\ �4j
 ���eIT�FF�Oh�JR�  �~��j��F�O��SS@ ���T �� �I6UI  O���#��}���9�B���'=��?{�Ҳ�G/s䯌�����V�{��$�	'=�~����$ I>��BC�`IO�$ I?�	!H�B!!����k��F�F�̻��EMx807�5��2���j�1RBn�
�ʀ�Y�;�Fe����y�謳 ����D���q����u���n�w���z�e�\�4hCQb��El�U�O�nb��w���t��nU])��H��u�XkP�W��ܐ^�[�bH��,J��Ռ��YM8�B�%��P$#e�u(�Vh.��MTu(=n�4b�����W ��*&��|�<yf�ٻët]'�ƑL�����+t�A=�b�ӸǙYMV DB)#�935?xHGG7b~`�h�ZL�V#Eg�Jc0�B�F\�c�3/FKF=@`��+��UJf��V��W��5��n�]�=m�����w@��@5鰐ܨc[��@MIZ�Џ���ZMJAt�(NAz �;�a|I �D9���8�����dL�g��7[u�5C�1&�aZ��Ŕ&ڙ��4�Y���e�1�"�����2�WDh������p�Fe3t3��v��z�DM9Y>�k5-�1x[۱	�#��R�j��|�mj��[cZ���E=a�`Jʐ�ּ�O�-fAI-�³U���b�b�UZ�H��� �d��ҽ��⭝��H�)�2)71e�[Z����V����n$�����!
�[�6Fށ�����;��;��6�"6�nT���m<6���(|��1DF�
+P��YU� ��{�;c/vV���#��I����HAq&�\R��*U��M��M��J�M&�IPsoуD�!{tvA�ٴw*�hcAV,R&�1!���;�,lrZ��lN)n��H"��%ժߕ�=���E��;�E`�Z����sE��m�Q"Ff���9A�{W��rT�v7j]��h�v�Nɪ��Cg�l�Gh��DkJ��C�@�^��&�$1}�LW�saE���p
MV�T�Q��fb"�ӎ���I#�B1mcۊ�[��̉�3`���d;ܥ�Mf�]�� d95D��ܭB���խ��tٍ"����<��L���'R�X)f�Iaf�c�0�P�I*�ٹ1�M4�m�O7��&��R�-˥I��W{�ɵA����#n�4�P��2=rm�s۬N6�3"����D��W��J�-��q�ғ���^���{�]��5xF�%ݺ����:����Ol��X��b�I���@U�$he�X����0M��%��RSe@oݫ٠���r�7&�^}��X�v�ZU6���^Ҽ�l��J5��Chlx(ɯ���$��ǒͥ�д��7���b��kK�a�Tk1֭��nBK�]��7,�f�H%�
��7S���d(���Ow/A�� �!���H[��,Հ��ݕ�p7Ԛ~ �uk��OF��N��x�U��
5m��<&�y�WI%��֝��nɽE���
jc�DL%(A��㸩�9��[�L�8ff���xj	��S�ј�%�d��w�c�-S��Z6"�f���S�^"��kl�/)�v���r8�jǢ�4���p��	І Al��u�v�j�
XTn�`
ܛVVQ�Ct϶�]b�T&�Mf�D� M�U��K��i�!^����xӬj�en4�Q��SwMf�z�F���t��� �D9���a���ws(6����b�g;-�!Em��Q*�đ�˱�en�=��� n���[�+��iw�#Z%=QC�b�@��4�h����ެ׈tV�
<�+Hc��u�B���V݇�Um��"c�񡲦�(�W�S"����	45/3�����HJ�dJusd$��YZ��k�ǲ�T9F�)���qRF�ݿ�*l~U������ҿ�ai�L�9yn1��ˬ�ô�]m��Pn��rZ�Θ4G���q��l��U9&�1ؒ9[�aZLY��+��f�t�d2����C�!hAY�����6���7f*R��H�̐���h��B91C��M���Wz���"�+e4�H�p���%�uy�R��n��O4%.�J��4�6s%�2�n�i=qf[&T�b���VX�v08,*��$�J�b��.{#ۧj�]��r�d��bK�ѩ��a�Bg�����G��<�P���>�y�. �&���t�C#���@�fE���Y��'��`X)��,��[[���T4�QY8qG�_����L���Pf�l���x��qX$��h����	��2��6��h�4�{�d��Q �Z�n��б4��ى��g�q��xEk���+�U1ȶ��T���	��ҡ.Ӛ���YS[57l���m��j�e:�Bm�T��X��
����q������m�$+f+ˋu!��-�u ����G�Dv�C�vo-/5�P����G'�r���b�dFA
�O^�V��Ņ9��2�;�=�kc�i���%C$�쀸@iKk@e�u�F��$�l�o��]��j��'�|`ZΌ��U�2��
6VVJj<�v��ͽ��� s4f}�h	�^8�
��0^�iɲd�aƶ�Dʃ#��iBe��*�t�56B��{!�n+ٽ���D����G�A9B��r`�L;������dȅkw�٧��u�|�sy�ޘ�E�K�)1(��Ցk+Qj*�bí��i�J��Z�|�JX�ܼ�T#�ķQebId]h�{�����բ0aˬ�p�A���V�S���sKE��6H7{��wuZ서A�
��*,������[H�xBL�/2�+��6/m���EZŚ&Q�(�՗(m?���ei^�Brm��L�vz8�;��r@�wZ�̴�V
xN�����ƷW
�dդ!Cv"U��%Y �`��@��8�X�G��hw�[�-� MU�0Gm/�#P;USm�I��
��(��֊{W����{���4�a��d���H�k �)c�Լjf�-����h���t�V̀�NԬ����9*ҋ0V�d�'K�P��W��<E��n㽕����C{���:<sy�7p��R�\ҕn�r�/S����:�Ԅ��z�1���\x$#NhVN��ݓEa��:��^f�L���ׄ���� ]�)��V�ʑ�wL|M��8�R��uCNR-l�ڳ�u�N�ZXP��$N�ݜ�u ��S{����2����2��{6���i۲	"f���e�tT�3U	�/i�Z{!U(k�jQ�	�v��hKP�
l�Z6iZ��� Q�a�+�h�I���a���ݩC/S�Ѭ�$�*��ཕ�a%�!W1a�h�w*
*�$��h��ؒ<�����ͪ!�ɘTe��T�j�Bf:ڳt5�ۈT�HφE^����M$L$e�&�H�k0<	�$"휢�B�7%�[�]m�^���Al����w��z�3��mɷ��S7j�9[����2]9�H�a���+�I4#�dA1k��L��wl��� ��;U����!�#͸�vor���2�
sC�Y������yi�$4��q&@FQ2��ȍMF�Ɉ2"-����t��f��yi-�V��<�f��f*����v^�]��ް�����@��H5,���U�r������lh �U!X#ŉb�#l��7�*�T��q�N*�2�T2�s�S�ݒ���YK�8~1ʛ����a��De�ja%�2�݄ò�$ԯ�af{	��H�<��g"p�a���j���%��H��{{J�{u��XR��E-��;B�h՗I`��#34ٻn�ѹA��e)N��\�7&�͐�@2�5�5A-fQ���A:�n1���Q�%�s)���t@���UЕ�d LpԨ(`͋2��ne-���Q����sE�KjAy�����-� ����(j��k*\T,�4�
(K��;w���w�b�H/�m��U�V��H�㌶���T�Y�
�֐yH=7y)^-�Y6�ݑ�z�١Q����R"hX���(���J�Y.��Orn�gT
�]M�.2c�2���f��p�gv�?f�j���j�V�9�l�����щT0�]*n�=����{}�v���&.�9l�@�n���$�#B�Xy$���X��sU*j��\��&� �[4n�x�;Cs#���5��N�m�Z�Q��p� F��X�kVcEb�ܡ�c��l��&"��C2;��0hؑL�5�����WC��4[�^��MՊ2���[�R��a��&'yL��"t*�@֔+�`�ͻ�M��������K�%�&1Na�wϗ`��M᚛$T7m�G�𢯫\����j�'	*�p�u���r�������i��SiV-"��%ԘӁ�Z��5͒gy!��Gc�D1�#!hd�ti�K�K}f-��S#qk�{v�[6��B�`ؖ���AKH�+]�lSz";"5g^h�1f�z���H�7Z�Z�;�tn��p70֫gb���,������mKT�#���g@e`��k&�۹Sܬ�9��\��<F���B�qG�l��n*U�{6��V-�.�����5�0ʘv�Aj�<��-Y�����{���La���Eb.�J��׋\�s9B��v�K{v�j�4n��t3G2�Ԡ�n�vm(�϶D(�E��|m�.;w)4]�y�Fb���{�;�pC-��M��f����cMLWF^�D�Q{��H�L[,�F=˭b\���ǋ�q4Oѻ3E3
�+tL�b�n�i����,(��Ȟ�ߴ`���(�}�����@�{be�*��^�Ow2�{,j��ٺ�R��9Q@`?f	��Խ��D�jԗ�S�"R����l�`6uՊ��x���fn��;aᑐ .:�6ٳb���3bۙ1��#b7����EW�ܷehNZ9-��!�`
�ܱj��Ss^)a�A��x6����7L��g/"���!pu��,�iس�Ş*xl$�-�uTh�0	��{xiۼ܏)P�E�\�8�>���N�w�a�ݽb�P?V����f�t�YYI�V^Z{� ���d'-��I��E�56f�`W+5�Z��0XB����EF6h���C��gfb��"��)'0�8JY��4����K!��!������=Lc�����e-עe��#t^�x&��/o�5C#��9[qF����J��A�U��[Qd�jIx��ZNcT�r]�2�nf��i�Ks�4���j��P{m鉺$�!S�b��f�͔ͤ�����4�:P-kfQ.o F{�)3�r~,�\�:|���bDk]ҭR�Aw�i[�4�x��i��=��!o��������مD3��y�@�fXd۠�UBo��g��tŰbX8-��2	f8͙�=U�蛍[�d�T�ڰv�.�Z8\��a��x������5-(H�^ř�t>�%=��Lər�"���C�Z�@Q���kg3$v���eZ���ܶ�Tj޳uTؘ�(R��B�i��6�[G�:��J��/�.:`��ڎ�'[�cF�ٰE@J��tؠ���)�Ǧ�(�X7u#��q���旇Dݴ�ٵ�Mϱ�)V�Ұ�ײ �eV��/0�ΕJ��4
ƔgFmXf��#&�E���"[:ԎQ���"˱�{�*�ܸ� ��	8��*�'uU�  ��5�U],��j�����+2JB �G4��[Ykl�h����	�Fj���6�t4�e��ӳ�Z�H^�GA5[���!jEu�*F�i6�vVг�J�5e�]Y�%M��j�.�4�Ĳf:�j'eT0�˸�C��话�L�ͺ�QhhR���:'n��T��BJ4GY�)�X�݆��ҽ�ɱ�<���� v ݺD[�D�Q7gUn�qeLWtL@ۙ�0h��{Q*��̹I�ӒY�V���-�iBu�*+!6�@��j�%�5�T�A�-�`^�go�!}�ATȶoEdZhǪ��es5��(��^)��5҄���Z���9�6����`-՘庈U���r�۰�kEKQÑͼF�cB�42��H�cf����c&��!eGw]{H�)�����vvkʹK	�ú���X�������jy��7B�EՀ���DdM-\֫�n�V,�������W����(dj��fnɎfP	8�;Vjn��aҎ�.e`D�/�X�񻱬�J�Hh^�U���N���������S1�M/��U3q�����i�{f��l������6!vm %��⅕�Am ���Ln�V��M�Z�{��J���
�4>��b"i����{Zȉc�W�3cقmA�6��e��(��R�v���j��09G��r�k���kr㕹��e���>I�BJV��m�Z�K7lٸ
S�z��)����N�t��n�d�QǙ��eY48�\Y�3�S"-v�٩�d���&!��	HϢ�٢��R@M���q=7Y*�5)\����h��fK�}��r���0+��に�#%V�E-�m,0S�V	�=Z�,��Ob��xd�1TY�L	ad���p]�R�1J�]
d#mܡ2�^�a�ZA��h���ˆ��c`j+˫ɪ%�j�õۆ�<lC�Yl��2\Ux���ϯ&j-n���p�7cA��)*wZ(�)c+#��ä�aem��"��Qh��dޭDb��7j���@V[f�k#n3��6�!��:ú�Y��J�kq�u/h��jG�kDx��ɏ^��eU��%�fQ��V	Y�᭰�A�D�+&m������-p�Fŏ��T��������hHY־����/^b�Ð�[�-.�਼�,�\>y�fM�*�z����KТ����d�(�V�a��6�а�N�:7��u���S1����̕c��{ysn���'^rٜօ4�ӝ�����'%�c
ZT�`"k�n'WY[�]��QGbgm+�Dq��TZ]]S�F-��^�ت�n�d;/w;�9�.�E%My�/���7�f�����o|cޤ�CչnVzB1�Iܫ�sI>�}�qu>���5wCk��祪J����Ő*Wh��x�G�����)F�}���́{]i�Ł85r촩�>J�ݹ[��b�țQ����)tU��;7,�1���v����ܴEЮ��o��Rw�S����S�S��Jz�΄s���ػ���.�A��4��	|��|�t����Eܫ������7/���o6�
9��qp�%�~��9��9pyx���_G��r%�[��r�-<Yk�����6��zM�轧�\�Y��h5{7K�s��7�os
�(��Գ��\^��0�w24enY���{tk[m�0��wkJ�/n��n���� »h�5�b��.g	�_�����ܔ�1���tiC��<9u4�s��gf<��<����V[�A	��]�Y,Gq���S_mWk���5mW"�?��뻛Kr��#���4v�}||Z�k��k�Y{3�d=_Y*��fɕ�{qI1V龣�AԵ��j��gQ�΃�Xq�}�I�cq��8D�u����:P�\x��e\Lܣ���]2��8 �=�̌������ ð(�U��s�֡�u��^+ݼ�T��"��o8Ӷ�u&Y�s$'�����\9v�n��M븓�7��[Y�3�ӗ@�~�ºC@ƫ�c���0 }8d���w�y��k��V�ӌ�wE܇
5/,k�j��籑P��L4������H�������YӫM`�A���"��]��L�Wp����y�����q(�vDu�����W*�!�jۦ�]F�Y�A\��%�s�:�w�1�����2Ŏ��Ild��%��%\Z��7O3��t�4l�ߧ\��W�d�\*�[7)��Y����e�FO�e��۷w5�5�AN���9CL���T�K��$��z��:E
8�sj�7<l��f w=�si�&RU\|�fG�� 9Y{[��X�h>y�*�م��Fi��죑л�&��l��Ԯa�%����tA�8KW�
,@vz�j�A�}�z���:�w�
��Ӝ_qv���\PZ}�>��:+���5�`�{������Y��uo�0Hb�*]7�Vr9w���=���)�z�
��o��"��8b�m�=90f��/�U!�,�=��(0�z���A��ǥ1�n�}�Mo0>��N���2����
Z��#1�r	M��	EC�>�]�;5-��mӷ�ק��n��Gg��3�*QQب2�n9s��]}F�"q�)����(��#���tw	�`g�ڡ��ԟ��L�3=���}B�go��p���u��G\zn+Э��[Ė(u_u9��f��C�b,-���7�6Bph�C��݉x�]��9��F��3�7��w��e�^�*%�cIk�bڵ2�n>y�eE�ݫZ�����'�;���khE������~=���-VN�(s�1i�1qCxgf�,���*�V�M=g��>�kIѻ|�7�q!u�uv�=绠�pdDAܐ�xu!`�u5Nپ�/zH3,#˒(.VPG�WT�7.��5G�R�:��M�d)�3@KT����^]�W�Mp�`]e�;<~���i5���oش��q_G���q;�2��p�2���g��sc�V/;��Y�3P��P��/i��=4�,`�-���u�'y�����+#ݙQ�Jȏk�l�9��LM`^6}�"t����9�_zh=�H�C�Ntf[i��3*,g�}v�pI*�8v�TC�nm��ȵ���m�2[��J���3,��&.&b�u>��̃4�$�X�ԫ��I�I���<S���Wlڼ��0`����W�3��P�k��X7�����eCW =W��K
.�$�W��kR<5a)���$&�Bb�n��
j�K�²=Y�؁�렝�R��R��������ꯗf�?����{��z���2V�Tust9��]{Ƅ˚�ud�$�3@�����������͗�Ohv�gTT����"�{
��=&�p�Nlt5��+t�()����5���io���<ܴܥ�T�Q��W����/bX �M�sb|������v��-i�շy�̎άW��Uփس�K�XS��b��;B���˽� C�{�(����2jVf�wv�t#e{�{��c�wM��q����kZ���u}�(K=y'[�W����2F��c>϶��]�q�f�Ď���-�Y׵kٚ��y�}{�e;��w�����b/;a�����O[�$��Ǻ��+A�o�;�xqj�MQ�q�9Ԇ_0S��.����P��q��+H�p�\^�k�M��Z�\��w������6�B}ǆ�>v��%��@$��:w'�$�'��W>?>�z�p����{=��+��G�{Y lf���"�V��Wmn�X�÷|�k���!��b����Um
k���r�#\\���A�sڈm���u?{���LV�V���1�O��ƴ�Nݛj�q����f齎�:��hf�Nٽ�;r�������i�$�*!<E�7ǜ�he�Ϧu�8��� z���L$�O����Ol��Y��i}���X���]�Li�=H7�4�]+F�	b�Tz-V�m�	�Y��Yf�48�R�O)tNZ��	;�2/`���wU4����h���9�3/Yh��9Rt�K���)��'e�e�q�0�y�o2��:PT��0�{�*E7�̷�(�#��&Ʒ.�e־�t��ֹ�Äޮ�)px"��zE���y��!]�Nw�Z[v�ك���G.�|��3���R0����tų�K3�|��:E*�5O�]�0�离�Y�6���x�8�*��Ѻ�$�ߺu�E�!76=
>|���*qw5� ]$CQ1q\�a�Ҟ���b�����xs�p#6NNh)P��.s�NgWҐ�E�ÜYޚ�q�6��3����,�f7'���Ԁ��y%� w:�q@��x�.�I�']�! ⒵M6OL{������d�.5�R}���#z0_g@�qe�z�� �4��W��ӝ4�������1Ҙ��%�1ne�]j�NŸWW���b�a�ڠd)F����Z(��b���z������1$he�'����X��c�������Y� �(\R��ƞ�ziԊ�.hT�ֵ�����G�r����Ml�;�o+<+i����;Y�a��~�¦�q>k6�w*�*c�v.g��Iqnqk7��8Uaz5з�LhB�vH�Yܑ�6�Eg�ޕ����P��sՀ��/e�7l�ݺڱejy�I�\$�Έ��'�;��^%M�l����E�h�[�>�U�����]{�����O�l��]f���u6[�b�;���{��HyQ�w�o���F��V���y�r��5u��������r>���0-����0�YFwe�{Z8e��|Wt�m���H��sr�h�Wۺ�W#���uմ�Y���5:�o5��3G�x��Q�g-��^]�瘭�0���8�`H�QS4x:^�KŦ>�~-�#���f*��Սn:���V2q��F���鏲ΨU���WF�=u�@��	�=W�:;����֐��D��Q�Q��J�o�$e;3��.��ضEl�D]�3u�装�@�Y�m�Z��澙�������]�m�ݷ��-g&d�-� -�r���<�M��V%��:�cP�+=^��Q�i��b��^�W�gL�6U!�p�
͆��zzС��=�ҳ���*�V!�u� .m�����VOi���|k%�/�x��.�BŘ�D�j
A0.�N���j�%��J�!˞���.�-CW���y?!:Գ'4�o�B��iul'VX��QW^t沇5��_�9[ΐv;僥���o�ZRyd���G~)�����j�oj����2��*�UK�L&�$q������-G�v���<r]믍�uw�q�'D]�]Ƴ�D����tSőf�xq�ҕ�Gی�Z��˒+�b�-�h�	�n��#>��C�n��^�{V��]�*�4�+��R���΅�A���fj؅=7�i��fC|eJ��j}�6�'�'l櫍eҽd�1�-ͬ��R�K��5�`be��"X��N�-���:�'�`��{;tW:��hM�U�H1Wy��6�*��+x�v�yN�T�#�[b>j�K�|����*A�|	
��S���]
%#i]��6{ޫ��.��X���\�o���ﱳ�RWS���#"J���v�^͏�v��z]�b��[D�)%����]q�����us��R����1Mۢ��t�
����z��Ӱ�I����*�[�k��C����[��>��?��%��k#���������h��.M���Y���� ��m�@!�ӵ�K䵼�N,u���aW/ �sK(�z ����b�Q�3l�|�h-t��h:���;�G+���z?d� <׈�%���[w�/N�شi|_n,�^,5��P;��-޹��"����"
�7ςr��5yj�O�{_�9[,Ī��2p�o�WVNy)=ݾc�|,��S�SaY&\ޙ���F�VmD����R�3�Y�J�)���kR����1��T���}u]%���v�ٺCg
i��3��z��#ı��t��/�Ӫ{���E�Ff�oV�`I�+��{93���N�A�q��:X�*c��̺�aX���z�hx^Ď���Gws�P� `��uw!�% +�#�M�y��6J����_�iW�Ɛ�8=�+���g )�^���T��oZ�.@oE�������v�]�Rخ�ɛ�)���RV� ��߬�Uw��ψ��x>ɑ�g��O.�o��'_$�ޗ]�DW�0�<;Q%jA]��yU@��w䴵|Fbg�h6��d���imi��^+Ⱦ�Au6��M0��y�-vg��eE��yx��-��܎��uÉ����e��:�ǎ�ޤws�n!�y���aT^��h���VWu��]�`��1oD+T4�ݳ�yA�o�|+�vd݆��_
���T�S��c�)�����<�W��	q�چ�o�6��HL\���4��;35�� ���ΎV���#�6[�Xu�`c4]�Sa4���w6��]��#6�y�$�L��t8q���Z�63��d�+&�C��3~���ilX��
V�8j�M3���+7wZ���'W8��X���cx�䓯v�=�vWv[���Z�Y%���ȃ%�U�8���Tʫh�S��܋�.�{_I���3µnuz@��oa�&���;���]u�H�V�x�Y��y�nf�d7�,Y&9[9EQC�.m�[���x��=��T��5M��T�͹�VuN�d�|L,!\D.#1+���H	�5c�_���7������u�򼳙 ��ֲ{�֞w>�o���m��l@��G����{��5N��A%ӣ�#3��8s;3��zo���+�7uf�{�:u�P�6��cu.~w��+y�Q%�Qȵ���t�;�,�}y���/[��`�\����B�#*+ٯ�{3ٵ\8�aɪ3��vn�k(%�ww�)L���0ԧe΂��f\%Ձ���+�k�b-$RD䮛v�n�َ��N��l��ZЋT�X�cC�ˑ��������o�t~���*��g�S�j#��d�Z��fy�x�v�9��1����.P�s2UzN���,-�tVܨ�γjB9]�뇒d�D�)כ���0�\��5g��I���ϊܾ03�vV��R����7RK�-�XB��-����o]%�S諭���ۂ##�cS�,D<F__��~�mw��Ȥ��q����:Z�s�B��OIQ9���@(]6�¦�{�5��Z����a�k���h��ZmERrܤr��N�M��/_<��+�E��j���7�¯��7o;���Q�]{��������FD����oD�ϕf��uPj�ףh-n��qnK�)g�N�P��.�b��V?���b�6||����a�p��?$7\VզS�k�T�bH�Hs�TrRzw~ 5ێ�>�{O�anVaB��}/������6�ry[� �s}Y�Uڍ���bI����7�˰f�k ys��v����\�ٿT"Cp���HB	���+gK�ښ�	���ǻN�	��֒b��<��:'��W��M �ӭi���F�t�klE��Vc<�nT��:h�E����Ә�Zxv�(ÙEVUŏ�ܛR�/�m��g3�X�/ 8%��Ԑ���yI�z����%}�ko�s�m�)�
�2�g6$#�ns���
仐���PG�+���/N��s&�VlJ��ܫ�,7]:`���
��t��A������{�{(aO.���#O��7h�M}��;���]�@�}K���Rk�es%:����,�o�Ι��l�v�
݀�����N��I�v&U����U-͘9v^Fd(v�{�XNց��/B�BS(gW
X�GlP"�[�F��&n��S�^���݈�a�uڬ9���u3��w��y�[��~�޾Є �	!I�y>�?d�6�m��Ef��/#3�Qt���#�N�l/ȱ8��*��L4KB�S�3���p����[ԏ����,:��E�$	Ӱ+4�6�^�4�#�ٔ{_?��C*]�3�؆B��Ne�LZ�z�����g�[,ojt$k�s�+�o:��:X]Ɋ緋]BoG/�]�F��N�|�%N]xP3�a�n��ḳˆL>G�����ڝ�Mm����,'�,A���/�Y9&i�w}���'�A�$��r6Ρ3/�	�n����2��Ov5�AN�$l9��+vz��K��QU�^�������m�vOm��8��P��/(�鹴no@�Bop���^x�F�����_����p�ܟx�]
+��#cŕo�-[}���S[�f^T	�JI*�|�`�r�x�Rϝ4�3h�7!F�^�/:��8�]��&SQ8��R�[H`��h�;(�s.��j�;H��4ޥ�(��ӎ)t۬湜�B���.�9|,�������f"貱3fs4k��-�w�&�����AL>ʔ�Of> Y*��rW�o�8�b�!G�@;Vzv��gն��Ǐt��mYy�ݡ�tj�{�p���p�67/g���Vn�M�k6H�ۻ�z���v���k�`���O������D{�����xw\y���zA�s7�a�h޽���19L����<��;�_�����u�2� ��7�-Д�t�Y{R��[[X�����\��Q��t
Xꛮp{
v�:�C��G��{@�Ev�	����g׏x��{}��Hӹ֙Ѕ���D�uH��F*�6h���92V"�tmӓ�p���
�΄ᩩ�|�N�졸�e3�cP�����*����,����`y�,y)L�<�1fg��X���z�����;PќvB�U֘���(����Xt�3��mF��7h��V ��Q�E�M�YR���w8tc�"�D[x�Y|���fZn�OݧT�A��$���i|'�eN6W���mEUq�	���۽�2O��i�gZX�*�6nS��(�8�=��w@�݋�roc|�=S��$ٝ�V�/h]劚DĊY{/�M�,�x0tw9征u���r��Բ���w�V���X�f�96��a���~6D��&>�b�����]xƏ���土���.'�O��b�bx]�F'y���HҺ��G���z^��-�8y��:lT>tgd��쵔�G|��+Oj�gZ�.fi�wY��Ǔ�Uo��/=�k^^B@�	�po�4�W��r��U�y@��V�c��
N���[���/g#a|���~�o�<�D��B�;ݧ&�OU�6�k�d���fU�ת�{e{V��	"�Qά]�f�f%%u��A��b�\6�1�ۗ.T-�3��K��t���7aAL#�.�-��V�#x�m�bz\o��i�{��%��5vάp!ڕ��j$�Mt����Ԣ�G��8ɛ�.@S�Rc��א�ߑ��|��nEJ����(=W�enu�/*���;�>җ�ٯ��Յ�[�Ù�#fM��I�cB�H[�I�.�=dVv�U�n.+\81�S?e�ᵈ4�& w�ݩ�Kr�ѣ��%Kz^K[Sh;����0v���=x/lg����"Iov+f�G�N��=uy&P�e��|��օ�(Ř_v�*�.�V�����I�Z&�։%	88Uh i:��K��މi�kAǶ�R�VR����K��m�ț��{��U���"Xɘ3��VU��x��b_m-u�"�&+FK*˰��t�ocuy�jT`�����J��ui��5��KƦB��AJ���6;��g�z3�%Zg75�=Dz�m��vn�T��s(�����د���_.����������]Cn�-�_��>���A�r9`��7V�}�!(����ϩ�hޱS��8*b�ӫ�)f�(���4����t��x�pP��F��7ٺ�/(SX�1Eu�V�[��2�po�4s�heX4���]+�1�mWJV�lՊ5J3k-�<�����M��C�+Q����ꜯb�^G9��®� m[[���9;�0�[�n�	���.��|��g�3"L�,ѷI��["0���x�&S���u�a��=/�މQ��=��)��nH1��E������>ie �Q*��X6���E�k��JiG��ojnwQ/��k[���(��t���,�T��X��!BC��6i7`$�d�o�9AM�-�ɐ62������a�8��nK��F{HFb5�����;�y���I[:�Ro7/�7T��.�}��s^]^���u擃(ˌ!�6o�1�P�+4�`ѽ�z�}f9`�|�ơ����ŚM-[6D�'�)E>xm�n�/4U�7��Hޔ��j�,��|
U%!َ�&����r�fV
�YQt<�����j=���dI�Baב�5B�A\]���k (sgD�W�q�)Zb��a⡏	�jm� ��u^�E���V��(V�Ο@�To/��u��ܡ ��.ͩsM-�OA��_��֝��a�����sa�P&�eK����='/�ɥh���X?'Ѝ�zW/tql�S�R.��bx�-v.�Of���,J�����f]�~9_	*�����dj��a_P�,M��[���|n[�"��v	�,C��ޭg��]oH��:{,�����Vs� 9˝8�nP���*�XV�Z[�RBV�B}�a�T�͖�{S;�+Ә�)7�d�Xm�V�{,�1Q��cHSCn�b��yΉ�b�
Voaׁ:Ӻk�8�z&\}��=�݃o@�v!�=[t����] �	��|L��fh*J�xw��2!���JMى�yČ�bև�U���nP��;J�@0Vσ��pm��8��֣Kw����ӄxzk�8mL>z;��4&�D�wYmw
����̤��k�O���+V�3�Z*�+d�1=�of�W���/��W�6j�X�6V���{a>�/�1��UF.<��(���.�fޞX�>�ٱ�(��Sn�����E{�U�:�r�r�v�Sj22d��C}��:��ͼ��y�+��t��GD\Ǳր7~������4F��F�~c����;J��̛�k�|%���C��۵�րSM "̫�k�-2�+N���=\�a�8eMn!};9'h�����eV ��ʁ��Ua;�bVp/S�F<y b�f��s5�����R;�d�����fD�����M	p�����yp'�+q`ЮY�J�NfD*��=��cF�^���Ö�F[f2_7�tX%���Lҵ
�o׉ͤ�e�M�-lʱ�]	��M��u�a��.q[I]����G�4�p�u�/uP��@(M "�EhO4V�&���\Q�[E0��;Vt廰Z�QӬJ�\���f,U�Ӓ��h|,.�on�ғ�1_C��|�c�:�3Z�+C��z[�0:Wm�iv�ͱK��m�}Ϲc��6�X�Z�q��k��	�1׺v�֓:6[���5E�m�`���^�.;�ewM�K� ��·"ݍB[qE��y}ְ���ݳ��r��I"f�?n��/Ua�ޔ.�ޅ�/:dh��D�Vw0��&�eJT�a�[�^��ڕ��_V��^w�^�O,�̻�TQc�ܕ(�n�Y�	�8�&�3s��ٹ��u�r@����C4�rm�)�a��[���b/I�+k�R1a�6-4]龒x;��=@�=�t��E��V%v�̥��0�G����I�k��\�vJ������|(m�iq�u9چ��h:�3���^��<���1-���B<�sA�3�W@��r�����uw���@$� 95�m��1i��쇯�D`��k.�٣���T�Zx.gE/1�g;�8ֶ����y��M�ug�=���i�x�H�g �R�Ħ��JQ�]�kL�܄<W
��c�dQ�CiXL���8��KZ��S�M�,@��|3�-��%�'��l����7�}��(�+��^1�����b���'�����T�vn�z�1*�|st�|H�&D%��V/zU�z�z�3ALi�*���&�L�s��<.���E��a�g!��6(���0�
/�	ܔ'5rY2C#�E����9;�	}�=�
��U̔m�&L�y��oSYP�2���s5X�:U���!�M��Ԟ>�%��8��^�]����C]��$Sq:3*��d+�S�={�.�'s!t�u�A��R�+R�jY,��Qߧ��9�Ha}Im>�mh�9N�(5,��3�V �]?\�'ޛ0J�o�u�}^�zzʥ�xz}�,���t�k�9�3 ��-j�~wtUr�G��-�XtW Ƿ�F1�"��b���hV����#Um0�=��o"�n��sk'��9��2@8	j�n�\�{*;%p��P*@�mnl�f�tg.�g+As2�it��'L�`�I��1�v��X�Xq�G���Esn��v��.���_H;����r�5WuΊ���#�fP�)�>7݂*0]><���$���.�<N�*;
�ז�T�\vH���ׇ��w�4�ﱛok�b�AV��W��z�Ш��s5��g_"��y��XgU����z�A��+k���1	g��ES[2�r#��g7,�ҧ��j�)����__:@_ʹS&��闪�������]fXW:V;!f�%����7����`�ɚAØ�^��cx��0X�C�;}��A5)ZWgf�����a�_̘��x��S����mZ���Ds	�S�s��}17nys���:M[sW��w٦�,��j�ׅ�h�ܷ}�l1p5��U{îoL�*l�Y2�C"#Y�n��r�Y]B��@���q��Ħ�b�cz[�\T�n)�AW_+mF%K{�ј��gw�b��j���A�n(etCD�$�d�N�|ynT�(�����8��˭o4�ʂm��˵� 5��5�V�V>��{q.����ein�QP�����Սy�i�@v9'N�i����n,��y��*}GjS9<|�4�i�fM�,cS��[X��M�A�m3U�#���0w}��<Z7C���k=D/��>C�|��o�Q�@��ol;6�d��g>U�fM��M�7ucL0�a��'p�2�E�'7E&/4���%��W^�{7�Z���8��2����l�o6FBG`��������e?f�:��ZC����ev�����E�u�@�D0��%sG���{3�=��d�m���y �����x~����
c��w;e�����9cY���{N!��0�n�j�ژ��Zd�dEu���tz3�M���Vn�-��#����� �|�6���#f�]�k����Q�Y��hpj�	�`,���}�9+$�� +��z�U�+	/@�8g戨cC���yLk��7X�:��We��W�|IV{��Fv	]�u�n�/��WxI���~���e{<Ґ�%��-K�^���\�k�(F|�t��ֱT�%eٹY]���b���[�T���ȵ��/E�;ǄQ���o�b��W�v�p.��g��♋2������taY�V�W1f�ހ����������vw��٥Q@�B�zn�y��ɨ��k}�F���u��-�.�'RUU�����q���IVn�s�Hl�SP�W1���,���B��Z�!d��q���0c�[�g�j셼�Z)�C��Nf�GIˁ#Z��@;��vn�K5�6eTX3]�Y�q\z�%lL��(^k��ffU�bjX;P�%��"�U]gk��D��Qm��YGsO%���`6kI��<Ԇ�YcG�by��:��6���ƌQ%{�q�`
��U��6��seq�;TU�n����1]uk��hˑپ��m&!U3E �f�ٺ3\X����i���|��
���;][�շ�COݧ�p�a�Ӛ�h�Z�F���F^᥍ʋr�H+r]h$<뙑'H����l�����6��iv�خV�_#,�G+��Gn��r�����YbԌb���sY7�&}Ό�]�nf]�R�Yvf\ɹ�Vݰє��9.�y��B�늎��g�#�o!�@f8��<��:����S�H�]�:�oN�zy����إq�xwa�*Dz�7{@;YW���R��n^t3OmKL�M1�g9�mK� A������z�f2eurɑk_N��gRHM�KE�-�o��ߥ�c_h,F&nfu(�rq_Lp�H�sq�4���s��a{�a�3�c4�������X�ƴ(�o���6�:y��X�'��x���9n�R�u�B]C��tp�E����������)���nM�"\M�b�c2V*��9WΤ��%��^
�E�#�~h,�����v�5���Ӕ�����&�
�X
q�9+�0l�c#�d��;| I��� �#�X�x$�*�J<��L�%gԯ���uDm/����:���� ZmŤ�eŮi9:$��kg���p�(U��U��轂��<���IXcX�ۗ:mV���q��]q���`!�k��d�N����9�G״b����;A��ݗ/���芺�iؐ��r�q��g%ĹH�D֏V���3FZ�Ho7-y]v�t�O��{���È�k�{
�����ȱ��\v���a$��]Y��wp�u]�z;��Ļu�{��	�i�s�t士��U�ʺ<A������f����vŁ��z��n��^�s2�C�Z��^^��l�-������+�O��������^�UV��dڅ�7&`��RH����#��p_�*_NA�+��w�_yU������Snb�/M��K��6�Pe�&Y;A���H�"�F�&x_f��|U,ʄ�q������ZF �� ;���k4�r��\�F^�h�P��c�t��ŜR�B�Q=��������7;s��K��5#v�$�!p�>&��W���:�
�ȃ���	=1��@s�z��V�u���� ���S惆�r�� �e��i���+�9�Ū�`��J2ۻz2��/�������#�wc�N]��>��WӶ�,9 ���ܵ*0s��B�Jp��[������l%w:���k<���:�	o�"�rmy��kIjZ���R\�!�o���:�;��N��ȭ������p����A��Iɜ�����#=��;�d�>仁�K����p@A}�W�L�J���w{��XC��=mS�M��8�%b�LeoH^b�]��,@̬.S�7�WJ=�5���X�,>�%�����=�nⅭݩn_?<߷�`�,z�c�*��W�"���&{���hS�N�z{��%P�n$��tD)`��4 ��[*;��MުP8��7�,\�Ԃc'X�-U^�k�}o.��Ny���A�]�lҮ	�hx)�w�F6�����l�d-̞)sP0c1]�ջ3G͞��,��v�����]�� ��k8n\͜��d�t�@ʺ@��0�"�]�zolEKG�AҕFIf40��73��u��a�}g��2�̂8�����߾֔DQ(��*�"(�}KEE*��X(�"*�������UF(�"*���b���PF*
�YF*(��D��
 �+��*��TF"�,b�ER"�EUX���ATX*�b+mEUQbƴZUE"�(��UUEEQQUdQ�DETU�dc��X"�TX(�E`()���V1EcR�b

���h�V*�DQ
�TDb"��TPX�X�� �������UU�������(�UDQ,AEEJ �#�
��"�*�EADT�1"(��R��"
0UQDEcE���h����X��F
1����Tb,Tb0b1X��"EX�*0b"�1EDE���Ŋ�X�V�(�QETb�(�EE��"���� QW�E:�{��p�j����D���,�|�b������4�q���[�r�9�9q�.+���Z���GB�go��m��7���:dZ4Ӓ=�^M�ƺ���!s��7��/�ւ��rL;�~ՃGm����9�;���� �M_$x�W���Sh��{Y)�lh��L��u�s?w�uz�6�tE���4��"��>��i���z*�N)�~n�.��܈�(�F�~�Q1�Q����l�7ՒN*���l,��J�r�oQ׳�~İ@m��A={h��5ƾ��P|��{.�3̮p��&E4�\�
��΀�Lr��8��ؤ��sѬr���X�sO֕D�ys�妬�|]�6e��r6�b��6
ܴ�D{ǅ�ROeE7�T�[����O���T&�<��f8P�p�Rrc}���	&��Z�L�B=X��8����=1<T��0�'YEi�_ZՑ^�7��yKW4�ǉ���J��w��DVb��u�EiP�Ƨ�1��&9���)	m�Q�'פ�#��
�/p�Vb����V��l;�'o}eE���;�ީ�|]B��o-�ڬ����C���ܹ{nwd����o�����0X�w�=Q:����':���t��w����򧾪�<�id��+���;D=��y�B�I���Nm��;z������òӅ�K0��[ύ�؍��Q[�W�Z�6���2#������T�Q���H�7ڌF�p��e������0��_'�gX�-qy=�38��}y%���:�l�k�G7�@��wq����]>S�^g�<����x�wZ>�ɘ�(��
���S���ˢ-�*�a����Et-�;w\>y��Jvo��v+�)�X8��B��d^
����O^�G�.��~a'q�q�}9͖:t�1��Do�����Վ3�j��a��e��t3�p�;}���N�!�F��a����&'m�1ýp��kk���.�;�ڌ�ۥ�tE=���K�~FT�o�.��U���������q��c��/��8����V>fY�X'��wu=T��f�X�m�����ٶ�r�ʇ%��x�[K��&�Fw<�V�ʊ1�m�5�ŘƲ����AOY�9ּñ���� �Ic���.d�q�5tp���k�P\`ީ���G]�gpQ�x;Ӵ����pY�n4 釧�}W@������i�����F���뽸��O!���C��p��"͕��QJ2�B1<�a�<gX��G�q��3�
��ZC�jv�%�*�6sK�ʎX-�X�%Շ~��w��X�)��j3׺곴ˮD��w�Ӳ�NQ^KI��������WK�#��Io�tQ��f���ˊ}$ޖ��<�<��D+qZ�I�ݔ^�
hξ��ծY�D�(��i��4u'ffXΰ�K�:�3
8n�Z�����a��q���D��t��s�Z	��7��F+J�сaЋ|�^w���9����s8�N���%z��)�������NO(l�4�
Oeqf�	����r���Җ"��-�EoU��n9�ؓ�b�W�+֔�c.Y��B��Y�W>�H��U0؂���U��8)R�1`�yj"�~|$�=)����<��}4�:jA�w�$�ma�[��kɝB�ٚn����HX?m7�V�ӌ<7�𸯾\@��'�3�~��ǻ�\1���:�'+��T�wb������ZәN���^m<��B�����b�E�$�b%(��������F'sR�)l䖩ȰҨ���ØH=����f�8^c�TL�p�<����u7ѺՄ�����هf���sv!pRb��X�9r�Ssn��;Of�{E�&�y��t-�笂�J�
}.v��������*}p�@ĭ5�j�]�9�į������(�il1`^g*�3����K�TN��.�_��b����q�-�*vpm69�w��+|���,`м�&	C���>��U\S^dt�k�tg(���NȲ���Zz'\S.�2��wox����QX:'�C���Aҏ��3��WAt��
������?��g�g;�6>�Q�&�b7JjoU[}�WS!�ف]Im�'��X݃���؉sV)���6E7Fc}1�C����a
{����6o��u���j�jp�1Os�D��j��51���G`�@�[�_����AU�cx�Q��*�ղ�iT�w���W�g$M��60����a���ǥ�ۭti�Xyb��r�����RԼ�U�O�C�TV]ˑ��˼Y#f�+��
0�1��X�޺�<�^��S�E�Σ���5-��\�Ɛ:�*l��z`f��X�:۰�'���h�z~]ח��-���a��R饜d����w��ξ�LK]��X�>�urK��9���B���V֍��[2�t�}4}��Uv[�]�@�->Z6}@؍5X�	ɤ�*��tHS�c��� .|�8�+HY�uW����o'���,b2��͗*�<,Ɔ<*�Z����$P_yu-H̼/���*"_^���A��,9�N���i�]�k#��ʲ{���u��VljMKK̜�R;�+�W��H07Bb��Ar�cSg��)z#r��w�wH�-5G;U	ۜ��j_�_s�X�'�	j.�O�֙sq�A�{�W+�
�M����+bF�v��ǃ�C'K���f2�0�Y��M;�9isK!�*Z��Lcg�bbr�t�r�����k'Zg ��9q&qBR�S�e����:^r��<�;4X�Ӷy4+�;�r���n��⧽/AFMj�}'�Gɳ#�N\�,�=��H�kt���oo,eq�{;#��r�J�``��[��<|�WD��LJ�!:P5¯��.Kȁ	*j>��z�A�-�U�1��A��=���	��J�3Ϋ"j`�t@W 1�$5�]zz���4T�Y����>ic��ݿ%�	!X<�q��ϋ�v%Utwb�&��Y�cU9�@�F�hud��n��1���*��x�p���,�F�rpIh;��14%w �pq�>��K:���X� ��>6����k�ђ��J�+̽�8P�
�(}ñհ-Z�8$�OB\�t'Bh�˝��X�S�W��6֥��?-��i:x���c����HXc�r��;��D>e�����7�|Z'Z{(��75-;8B�(�s� �B�m{)���(Ŝ�0�{h(�N���2�kK��B�TK�05�LT�ns�eO(/��J�Y���J��d�H�X��>�l�Sד�Չd9r�T���k��
�����P$=�k�jǘg1�WX1e[��r5z�/k�Kg�%7.T��NUƢ�Z�Ls�?I^�L�^C+/�Ns�*9W���"��~�Շ��A�x|,��t��T�lcLܻ����ώ϶�W�'�D��V76y�}��ΙLV�� ���j�%\0��+�~b�UBa�
�W��xX<��l�R�Ώެ�L�p�'<V����0�),:�M:G(�r�L���L��Ugܴ��΋��M�R��l�m���1U]"T�@t�AG�?���.�� �o�����������j"1��On琢��ژ�$�g��|�HZ� f���]���kɰF�39��kMMm+�-�,��H}r� ux���0r��@t��]��:�c�v'�[�)�[����]ty���-�H�k�N����p�7��h�¤�U(�RtGK�\z^pg�1���ٹt/�\}=�MЈ2�@�h$VE0��3ܸj��ɦ��^*S��S��T�>#G�+5\ه	��d�ʫw�[��К*F�ѿ}������M<}�Hw�8GKۂ��&��k��[�-q���q��/S�j/=<�/D��cF+خ���s�FR������P����FeK�g�E���y���8�LP�m��g�t�̬?%T������_m�.z����O%N%m�c-��[*vÃVP?��^/���7Γ��:�]��_3��9a���������,L�M�e�n�~�&v$�L��cM�8������t�'F����6V�f�M=']�';��$Kj��y���c͝�A������<vfU�\+/��8�_HG�9�ow#<M:���~X�♹�Շe.����Y�S�f�o�e�|�`�p�(��F�V�=fsqQ���x���C,��*�	Ұ���֜�z�D�o{ U\��U֫:u��zw�83o�viF{�
��u�hui�a����+AŽ�H�2��.QWd�+�@�̩O��Ͷ�ec����^���X� V�O��}���)���<���`_U��*�%���nC�dSX�6;�<Tn��r#|H3���{�B�U�ī����.��޿m;�/Ɉ����DP}t�B���Z.:��
����A����-���˶��q�z �W�d�w���t0h!�G��{�RtQ�p��].<Xv�3&�6�n.Q���c1�w���߮qZ3>��j���V-��hK�pV����=SX��;��E���j���FzT�9�VÎ
T��l@b�Q��=,�������43V�����4���b&�)�Pc�;SBA�pF:���Ч<^E�5*����R������G@�B����TM�`�s
�{j�sv!pR}kӬ��˛�t����O_��8v5\�#�N:�J����(��t5�nb�C�q��D���]��t9���y���"�7�=;��l�~𖮺U_���èJ��J3ᴬS���}*�Űh)�#i1�b�1R��ʼ���{V���6�3N����x":Td!p2��#uU�����U����j�cWx��;��1�$F��W/��t��xx�AvWz@�A������5vx2*�ݹ\)�dͽ��W	��!���dhޜ= �#Ҷ1[���̾,LM�g����Sxu��_�x�+�\�l�^�O�$=�C)=1.A9X"W���mh���U52�:u�h��T%h�b텡m�÷υ<iK^e��ov#��;�ew֥��h�.el�^�&5PQ�N��
+7(��T�ͭ��H�9������j��'p�J�/��*�b��+��m���*11Y0�\Պb㫍����trl')@O���\X[R
�	}�3c���_�d^�k���ь�'{�7.��w<@��ɍ������7�4��W�c|_�Վ���b�Q��h�㙈I�țj��WN�L��Üa�H��Oy�{؀�BϘ�����bǄ��!ά�ؘk�9g��BtCr�Q�.y��5]w����ɪUa�OD���V!ri:٭�o�NO$��r��Q<�{mϥ�ϋ�m�0`������f���J(��Q��S���J��zU�ݎ���6�QA�d'V��N��덝��w�\1��ۿK=7]�fV��{�z�{�)qEb���T��l)��ƒ5�[6|�ӗ�7��6�Z[��9Kp�Wjuz(Os�ω��%���V�����S�˞wM�A�{��R>��}ڔ��o��s��m��||/Ʒ�p73c�N�҂�R�F��p�.n0t�>�P�v.�}p�jeo,��`�YL�=ꓻU��흺s'-+�蜋շS�OM�G��yK��n�;�cb�k;a�+)je]��7S*sS2��'{��)����=8i��u��2�������6��ɜ�������l�(C�GqSq[
q�L�>�5GK�T���
 ���6���}4�m�2��.ie��H)����Hl�p��}��U�H�8rm1��ye=�O6O��4B��2���9]is�⮼��lr0,R�sNK=p��'<n�hP�9�p�t(y��S�ڭ��>�������肱������U��l0.&�5�y�\i�a��{�ob���R|G�����a�ʌ§f[�=ޕW.m:�:9.C=�i[�0��N��k��, �
����뉭b*�WMX���Cj������B�����!��u��;ӥ��ޭ򰃯tvΦ��u0&ZK��Kx�0�]��&\Լ�i���1i�Iv�5W��wa� �}�*Ls��o���$�}Q�d�rЎۇ[n�Ĥ�8;��d������T��ű�q�}壑�E�F��* �x2�9`k�2�f��6�Fi��#��UhE�a��q!Nj.%���X/8��W�#!��&��/"���z�k 3����*��ܱ[_/f�����lZ���uq�xݻy|�٫%�����	�>U�:�nf�2f�Wȍ�HI��u�I�,o}�Cl��fJ>5�U8s�ZԶ�p�c�Iݤ�p<̫�[&Rh���ɼ�+yc�z���t�Y���$�3�ˮ�l�1ՏF�0�Wf�q�wt㱚���/��'�.�dl��'vѬ��`�G
�+� 0m��x�,�p�ԂÄ́�e�\ͳ;�jB**2���@�q�r�zu\~A��M	��R�m�]g�~�����Cu(έ�j1oj0M��Q�H;}�v���H�CH�҈�Z*�$�@]�s��V�B�<T��5�U�������j��zwc��[i\��t]>�b8�d�Xk+�vYW�X�}�#]�tm���V굘�)��5S�p��o�b���ͷ�S�iF��A�5��dWz�7��$ݹ�]V"P�}E�0Y�W����b��3Ie��!�Hh�t� ����껖3'�.(���t%���ȩŻN��H���V����z}��a𬮞C��������5�!�>�n�z�W��B7���fux �C�kOQ⴫�ػ.w�CKؤ^<��L�cƳ���:L�rM²��3�/��q��Z���g�P�ե�i�e�a<��ǆ5D�ڀl/|F�LW�����7��Is���7=��&�p�
q��)KF��^Pf�����P�O1�� �Z�g�a��yܷ�("���� N�6�j�2��f��!�v�5g�ϲrKV��CH
N��&���7->|�$
��ll���X�%p��^��	�Y�ė�~����Q[K��wRQ��X�pv&��9�Jz��֨�gUN�pu�����ZY}hH���T4V��͜�Mk�1oFn�T7�J�M�L(WQ�ٱb����aŜ0��ݵ}�Y�Q�͗��/���}�v	�,an���cHjfL0I�S����h��j�4y�o%eڬ�X	��ȫ�b+U������XWqYi�[B�hB鉓E�1��W��]�\Yb�M�.�m�G��4��:5���CD�髼�.�{Ĺ� ���R����3N�"�)�"���XFf��ɨ}�۝�"ۼ�f�8섊{��}an��Z%�X�����5Q}�Ѝ��Վ���i���*�lYkH^[ӹ�v�N�s������Z��p��4��p�A�l�;�,<:xk/��[DQ�vfԭ# ��sk�97ɴ��Ղ�hY���(��ꗁa��ͬWQ�c�Z�x�-m�e��[N��KZ�x��Y�������\Ӗ�A��:�>.;�&�:9)*ˑ�/���ُ�\���1"PQE��V1��E ����V"����E�"��Ec��E�1U��AX�b�AP`�`��B�J1H�0Q��A1U`+R�XʔTEX� "���Z����PE�0�UQ���\kPLePb��TUU� �pˊ(�X�Ujb`0UaZ��)*�Up��AER
[L�r�����ҎZ��G)��VҊ���PY`�TQ�R1��rʬF(���&5�Ub*����EF)m��H��0�PU��#+
�,Q1ڂ�aPUb�**-J��U�%�-�b���>�A�+o�q#��,�#{+��N��E�r��ܤ#����;�����ҥ3�=�����m�hIm������P�4qr�mg��}���.
e
���c��I�Z��ڴ&�Ʌ*v:�ln�f��nj.�����
!ì,Y9f�����gg��>>J%��
��&;9�	�a�r����3C9X��%YiM���=1��g@��)-�t��ے8_�TJ���0m# ���-���s��7ˬ�>���~�Ǧ�n���aD�"XsS��JW`��#m_]�;5k��E�q�ϗ<�L\+/���w���c���B��\�"}R�M�����i��4�����Q���b=0}j��1�n�a�T�F>#G�˹��{+�k	1���HܝP������k��Q�5R��Jŝ�V4h�b��N	�M7�.X����Ι��1^��K�3&'��f;���1Q>Ÿb�8�����ʊ�AN�,�6=��X�}W���9�,;�%\BfbQ�p�X~J���)��]d;��C��65v��N�7�*&�9��P-�=h���[���o�'O
t���7�^��~��m�TJ� �$`]�����U�m�A�CzrE7�}�L���{-�
���Ky��!
ǁ;xM��9Ѝ�� w�U�����] ��Zڰ�7b�87�S`��Gew�N^]ד/yg�����ufME�e�|�:V���⻔K%��yܢ��=ã��g���}��ނx�[h�}=ú����5*'�������d�z��4�i��t�!}����z�/`.�z1���c��䗍Z�h��%_{��;���{\^`��T\Eb0{K��f󻸠�}X؝8�pl>q{�]b�Z�xq�	~T�jYp.����{ytAs�����T䳙M��-�'�'e��x�*������zmm2w����v����!������˹'��l��(~�yU0^q��31R�l��x/�A��OD-�Y<�9�Y`b̴�Y+����z\���{�^5�4����5���.�-=��'���j����Z[j����ܹ@i�͛�(x���vZ�UY;\ݩ4	b��_fu_�o
��1���8a�f��-��:���ݪ��.`�(r
��֪eJj���S���':�e�
���q`^�:��Up�V��,)r�>���!	|��P�)P^D 	�DnW2�%��Y��=|��,B���G���C[���o�'N\�B0���KۋW���MЉŒ\�V_��Dq�(��Y�N]펃d?t7C̳����TqIl�g��}�:f��>X��P��u�Ķ�X�:���3p���<G��T�vQ�8�5s%�{׍��Y�t_:B��sf@鍬��DDE;��YB����|譡~a�qq*��LN�B�:�71P������������׋�뺳��v�[�j���Pm�sӳs���J1)J��-��Z`�)7֩������8�J�m��{��ڱ�B���M���p��D=�T���U�(�R�8+�G^����'�gE�������b�cn{���}A�!��.VDҸ����ßq�NӚȮ�Ȯ��W{|���!���\���Αs^�L{c�'M�U~��x*P�P�U�4uz�swt�o#�6�N�ha���q+DU��pn�^罦e�b��:i�Q��*$�bv�_�*Ѥ"il�Ѱ���x�=B��q�w�*@�79��0Dd��96o
b��TS���f ���=V��Sv��6�'�ܕp������؋�MS�H�~�#�߶�X��1��5�l��>���(�����6������;~8�r��.jR�Ѵ,Ve%|h���C)��I͸.��HZH`X8F��)�����`�ŷ���F��;A�P�2����VԬ'R۽�T��ЯFPK����Es�g�=�b�����1v��GEK�W��D�����ưd�Æ`{�r �M�͑x^6oό��u{"a<�"]ȹ_@�;f��)ԓ���{�xj�Ԑ.&�vW����<�����/ܬ��5�3�3,��L���(��ղ�	Hp��L!r�*��N8�w��d1;��	=3�f���A�������+�FE�R��MĊ�bD�ב�:�LF�i��aX�7��lvJQ�?y�D��K>&$lI�pC�F+:�^@�>)�:����
�_.Obc�U��k5����S���=v�mt�u.���M�cڡ(A�諘>�L$j+��V�B�kA�v�#]����L��Z�*��8��7?3�c1k�E�N���<�a�Ս���������i���2T�T��ﶶi���HO����^#�J阃�%�#l,��c�,�ة	nuť(�8�lU�>��Lr0��\\՗��к��wN��Gh�]Vܼz���P,�ޮƈ�7^��KʾC����w�CV�&;$6 �]7V[�cVD���x)Jm��5걸���C{���/t�br�p��e-7����Ur��:�������O�G�e�ʙW88h�˟y|��xҷn�4Տz�V:4-��L��tJ��cq�yow'��M���u��ޓ�]BSZ:of&��q��55�-�m>]���`A�w͵�Af��T�F��Rtv�ߗ�P����>���/Օ�8_B_b٦��	FC���|���b�Z��h�ܼ�.�nKT�w�Ǖ�{�S�^��z#��ݮZ�m�F4���>�']5&zU#�̈́'���Ib�Ԛ)oz뿩A�+��W����I��s�`'�'�p��I�i���<�2��3�Z=t�8�k�i`�^����-��X��2��rÞFY��F�iN��[=��RaeAbӥ��G(c�����:�#k�r����4�ߒ����A�Y��~��j.%�4ý���l^��2��� �#e�.�aƲ�/*x�����M�	
�P��eL�I��[���~�E�qz�Lv�sY9������Q7/W��W�K�k��]�ϝ�.��;���M�L&NFa���B޵�ooofߛ�s���k$N�t3Л�[��a3���q��a�҄�1h��K���(7V}�<���ߵ��d�ܪK��-p�*B�T�J'�<���@����q:�\Ό!�^��IJ���P�)w�����΀��#�BL�5]I�@�G�;y�T����0'l;�f��3�)����&:a�8��c�4z�Y�ַ��\T��ErqoL�&�wJ���Dt�\�;�6�䥋u)�������z�*�{=&*ۆ��'/z��C�K�%9I7�&����Of`+wt�(�яܪ{<Q̯����|�i���E��8i1��w9Uo�̄L�����ڙ�'�U�xG���E�69�+�:�J�ب���xY��0š�w�J��E���x���A	y����W�T
�|�8+ȱZ��hTO�tF:���5�t�������P���6�5gc���<>>���p٘�}a�\��`�	�'h
w�T6��h�HD����n��Mιt�v7ns��S��=s�T�9�"w�y��t�����s��x�}�wK��]��p�MOb��:"b��LT%��ġz|5|4���՞
�7mL�}eML?�Ρ�Ѡfz��+h���>�S�E�7�D�Ly�Ց�н����=��l�����n鵍��F����	�x�w��ذGW���<�w��m�0�><�X�h`ȸ����o�� �wEl���g7=�D�}늒�a��)V*Y �Z��c�x��\Gq�:ɼ2v�r�����T��Y�[嬄��X����Z�(Rg�k��mA&��DA%�adŸ�|���2_el�7����GP��z���:c�`|�t��Dvܠ�ꐎ7��w��E>���@m1*�%v��0��{K w �}:�#7t�%���8ۉ�����S=���+�μ(�7Ƕa�xq������Y���_�K����b����t��Y]�\��<�ˡd�V�oz(l�s��U}��\%9�]��9��� �TXoS��<N�~u�'3���Ӯat�8�v��b� ]���������eĹq5��u�1�
ya�JT�7n�Dc7<����t���	󱟧������\ZC<�VT(y�Ѡ�2���a�/1(Ƅcn1�)�{F�!�T1�g
<C�j&Y�\��1'��0�{�-�$F��7�]:Ȅ�˘��
�#��R����S�>m�m���B{νLr��i���.��
_�}�t�m�-M����9��xU�٬vz{�������6�bx�JTK����>[8�*rF�
i��T����{;"T���\BU9~
z\�/�����`����uQh4/ܱ��/|��ˏH�:��W?��&,�X8~��Y�㒆����$�d�OI`��lPV����aϻ��)�ۊ��[f��������\`l{.'h�Y	�1����sr�Yi�T�;$��a�E��;u��雘�ٖ!(�޼`z�`B�"𧚺���58�W7��#��$fٍ���6K��a�������:#6ۍ�3_>�#��l4u�yށ���(PH\;����|%�*UkL�*����_*�It���I��m��ִV�d9�'9�Ğ�),�gI������v�&�����J�N^u�f��$�f�:�I�\I���ox�f��%�Lw��G�W���^�˓���dW�<x*}^4y�*�ѮT�@�),��M�RƬd��k:���n����b�C����=�ga+;F�����M@zb�T°c���>3��b&��}�\�rUXS
'��˹sp�l����=��/k�\�-�H�Ʒ�n#�)<��e�R�WN&�C8)�U\�VxO(ʵ^�S��Q�y=���6�Q�C��o��!L��I��q'�K>{A��,9�Õ-:��v�gZ���T�T���]��5w�R���TZ<���V��)�U9P_Z���C�������ۣ-ʔhp������f4�'vz�rk��Q�q2�#	�>)�Tj��(���9In�A�6���^=�ٳmΘ�����\��U���<kkh�J������߸���Z
\��Nv���UϕQ��Bu<�)S�;��Vnd���o�~��=�t��D搳1�66�f{����1R��p�\)�8ջ�IO����`��p@Byy�h�@�ro�%-�1��]�G<U�5#]C�]b�V���0#Ʊl�+6�9:`$�C�uw��7��ﰁ�urڬu��3v,n���B�u�Yv��o,�-)��|�UC�t����W�m<��?}�>lw��]00Y\\����o�M1��;�w���Qw�ܭ,\��WT�(U��7����\��0w��#!�'.�/o';�U���P�ˮt��N=͸��~n�Y:¾(!W���1�X������[t91���i��R�o�z����l�2���r��!H� ۯuH�"���n+�
�l�lR��fX�y�eG'����H��_'f}�\�Bg���G
3\����@�LY0��dpٺ�w�Z��p�LԵ��iJ7�W%K K쨩��Q�s����"���_�ޯhZ��6��'�GG���;w�A��.����`�;�ہp�����	�[٪��P\@��k�f�Ҝ���,�bS�	Vk���a���@�]V�>0�9�,��,�[�n]���c����-=54��ϴ���I�	�jМt�:0B��j.���f�4B�ِ�]71!���={>�px�cf2��M�>"��g���I�:�"�(r� ����<�Y���`�C�sy{��t<-Պ�ڻ&�*uk6e�5�]s��=O"x��y��U!{kz��q�K�9H�&ֵ��f�e�`��ns	��|NZ\������,�CˇS��7^�lP#�����i镶�:�%U�7�z=��.�ZN1WY+"�|��>m[�����ƣY"u���c�5�p�k�]�9� ��̠$#�yc���U�Ҹ kܹ�&1��Ch��j1
>J�B�!�s}[~��d��X�ԉ�޼�1$��A�*�z�r��9�nO*�c����t pM�o7+�z�zo(����/��;)�wTV�*b�l�;��L;�8��|v����"��2���jTa���C�L[��g��Hb�[�%Z�yT�:4X\k�VE��!�s�v>���:�������ĥb����bh�7�d�^uu"j0sfC��Z���>��L�=�X�!I����%7S�"�0���X���Wo�.��]r��w��y��6�r���?NMJ2����v�8dAa��3���g�/�������,-�E�Z����Op7c�ze�޼�G�$��~N������W���tg�,��P,v�������kнMor��0d����QtS�E�](�)�S�8E�W�<>���a�|s���r{�.�f��)tw�<yIٞSw籅����u)wA��1Kڨ���v���lN]a)k #u�1}*�u��q�ү��V�:���;��<���Q�@�RL��؄Ah�YՖ�rnH���Ѳ�B����|�,�x��d�L�'г�¯k;��E�K45Nc�޵�Iě�~�c�����2'պZ���B���vU��oV�/E&��$����L`�����ɹ�7;��y�&��MggN_!ÖJ**{,��>d�l��-�I[v��ķ]G�97��X����G%���4d7��B�&$)�B����+o�t�>{�3��f�]��Y���f��p��œ��R�u&q�\�Z��nV�Paf�e-���a�KǲM�ٮ��d"��׆�����ej�HiT\��d(Pj�F�l��2&n���}آ�z�ݤ��w>Ê�u�Ȭ)u�ci�1#a���x��$��w��!{a9����EaWݏ�A\�pov2�)E����ڟM��poSe貪L+�
U��w����H�;����(h�Al���7sEj��E˶T�P��u����B�!R�l9{���g��J#�`͔�cV�7�$��8��D�3��[�Ċ����6#������ C��LԭL���ܬ�K�~�����_F�/k��V�����a�Qe��K�f0n��	�Pȟ�3,��CT:�9��M�*
����T�
��evGP)|�>�Q����ڋ��*!��CJ>����m�3�Kb�k�'Hz�1�.�(�`f�e�C�ob޵Znsw~�J� r+�z䬦C�pr�Xn���yL��k�+,>y���$���"�vl:hū��d�����,ӈa�v���c]�J�����܃"�Rѡmt�`M��� :�B�S�vSy��z����^W�Q�0�5���u.�!
�|�f���>�ß5�.��j��m�,�Pp������ЪjRo�����C�Ĵv��ه|jR���)�P�*����9����pS٨Mnn����r.��L�c�\�G�VS��;��2���<��}�X:��秖�,O�/rt�/ss�}E�v�ދR<Csմ���Dl��ʝ;��<��`n����u��q�zU��{(��uՆ����sH<}�w\I�i���}��+Yvo�*r�B�v�+[���[�v����a� ����7���CK��xd��e�`��'n�����f.*�u6u%`�ޘdDaC��w��s�)W�Sc
�`�w��Pi��������$&�ӐoF����CWPC̹�H�����ӼS�{��RՄQ@��j�J�A���2�t������t<��������sp��'��r�]�0�F���"I#�s&n��k���=�D3�ʹ�э<e�z��f^^�m�^�ۗ -q��_i`�,<N�wv��@oRE�EG��������B���DDU�E��+ADTX�+DQ�DDd�h���1��"��Ŋ
�,���T��DRVX���(���ơQh,DEdYP���aT��ZƩT��("���V�b�EU�c�*-���AX"��*(�5UT+AEV
��*��"�V)AF��e(�L�X"6�F�TQB� ��1U�P�(�
�l���(��+G01�Dr�1ER�mT�("8�\eb¥Q�Q�Q�W(�Ԫ����iX����b)kj%�Y��Ĵ��A2�V*���ʰ���>ER�(�#lY׭lx����Vl\�,������5n`��kk:�2�^�w9��nj�k��u^ �0&�z�*�V8M����z6�6����[|����A�����؍(3�|��9u�fϣ)�TF�(�'��ޘ�Wn��ImSsHW�i/oEl���s��2���l<:vmdPc$����U�JoJ�Mo>}���Neʹ��Dߓ{��7U0� sj���kV�̪f������h���D˟���&������'���%b9�l�%��� (���;�{���S����Ϳ0+��Ciԟ;t��_�V|�\d�R�aH/f&"�]��(:��u�j����=cyy�����[�gS?�����ezv�a�R
矴q�id��Vq���9���R
s�gY6�����P�����>�M���9�!��!�a��,��Y���I��7�u��ͦ�vs~hu�{�(�LǢf=���%{/�Xq�ז|ϝ�c7?S��eE���%a��1�X�'Y�s��0����������L@^�'�Vm��z��v�;|���������_�*�����xU/��~aXm:Z|�+'�3��� ���J�O,��HW�_�+���{<���u8� �sZ=d�Y:�Y�J���;���A���@��7�>��|�����o���:���`zצ��z�gl1�"�R��~��~a�1��1I]��LՒ�βQ�d�
,�Æ���
M�D�����fЌ�A��}��3~N'y�v��f��#��}���ǽ3�J��{����R�;�P��R���0���L��g]$q:^f����P�i�C�t���1:�&٤�H{��猘�����w�o�������������
å�8�!ԕ�,��sG�>aP�9�agY+8~�u��AI�(bJŨ|����O�Z�wY��Ă�|�>M0����j�]�����ޞ�mb���m'du��{ǵ�T�Ƿ�o�������>����o
���]�s�u����=UvU��֡���c��c�0����9�:���G��\T;y��u�SF�j�]#�~�;6�.�E!ycwv���8��M���Pe}�~��| s�<��_^~w�����6�O�J�°8�+8�g{d�OO��"��+=d�8�>B��ӳ}�@x������A��+&�gXzg�*��ĺ����J�q7x�~`V���������\ƚ�Q�̬Ϣ)yL)3Dn����P��E��X�|�yCi��������HJΧ���M"��V/y��O�:�2{2�}b����;�x�i���'5��{��������to�IPY��� ����4�2x���n������?2VVJ�a�߾�����5��"�_��jÉ�i���P�i���9�jm��Q`|ko���wk>ϭ�oS�6�~���9������l4�'��sP�Ʋyd�^�b����
���֬�!�J���i�aP�{x��!Y�J�M�z~�$�N1jK�ݟs�+�y�Eר4��ϲ���o�{U���Ofi'��Ă��0���aQC��@�+�]��4�]��^0�%OKa�+9�&0���Rz�g�o�4��*N���g�c0������U��[���?G3V��7T����yx����U���H)*�N~��<�!P��3��d�m�O���=d̡�����S�(w��(y3Y
�8��2m=q�Y����_�\?)U���fxu������(�����x�0�3 �b��CL��x���%��sS�%@Qf���)'oI�&�v��ﻣ��T�&�t��Y�%~gֆ{J�R\���\��VZ���?K,9�c�R>���5q�����OKLa�Ă�;��f�2TY7��4��Vu�!�sf�.�uO;�O�6��;�N?�1���а��q�w�tO�mI]}M��<��޻�yӻ�ٝ��=aP��-�u�B��MSL�
���ܰ1'�����8�B����`~ˌ��0�*)Ý�4�Ԭ7/y�����������~aX����w{���i��_���i���d�t�rE%B��~�!��!Rb~�o�a��q!�IY:�=�2M (�S�����Sۧ��L~`W���g�N�M!��a4�;�Fk���=����ח��wP�mn]'�r�'�VM�Π�j-�H��-3)��M���s2���Y��B~���f\�u�IM�I��F��t�}^�]\:uJ/f��Z��}E�oYx��o\f�,�AM���.W7�=��G>\�-�����ߣވ���w����gg�	�DϢ?}�d���$�Ӟd�VT��w�8����?�6�P6�.d?0��|�3L��q����06�u�����%H.��'uH,��}������s��}�yϿoy��'��9�N��0�
�2s���x�Y�%|��u'�� ����a��Y?}��0.X}�������<�ؠ�L��
��Vq�e����>�J��{��9ߖ{`˵�i$�����[�ğ���|��'<���G����_�'��rɶOX>�����?0��|Ad���"���9{+k#�ڪ��]7��g�>La�ް��ĩ�,��6�_���8�gT=�:d����d����
O���;���N!Ry/~�c����x{�6��1Ĭ�q�wXu�i� ϻ�yAAc�E-��P��?UxUH)/H�ǌ�L y���c���뤂�2w(~՟3I�S�z�';C}�k�
�1�Mr���f����x�P;��i<@��u�Q6����A��ۂ�X[!^��+�'+�Xc���=a��g�0g�J���Y9����P��������L<aS�l�8�� ��Kq���Ă�?}����LEN�c�,z6an򝝡�����񘋟G�I��jz���2Vl�rM!RVq6fgPă��&�M'��`i��`bz��dXu�$��xI�T<a�ϯX��
�u�]yHV~[�O��f��_�w3�r��O�}��|�����l�u���
��S��OP]��u�sY3l4�É���II�,?=C���H/V��d��"�Rz�_����f�������o]���b�9g�i��0��sa�8�VM���߬�%H/m�Щy�6�ߙ6��'�fM0��'��L���Ͳs)�X~f�b2Lǟ�"�����������F��+*�_8}���|@���;��Z�Ĭ|��i �bT�z����a�Az�%w��c���$��2T��wL�������!SL��z�4�������Q`��h����r ����z�G�e�^Lw;��C��C�d����~�_�h���e"u�̍�q������ �&aY�ݩ�uI�D��3LR�&���8��h%_oԝ�X�K�ƨi�o���0��%9i]��:e�h|��z�aȦQ�������j6�F_�z""=^���x�o�z6���C��̗�T�ZAx���Sh����;�Y����� ���*s��
N�Y����6�\a���'��@�w�4�S�L�Mn�i��p�ྚKs�x�L�*b��vgp�I�����~�1��<���u�i
���4�T���&$�tyLt��W�����AjN3�'�h4é�4wϵ6�A@�����q7g>�ؑ9���O�g�"�=�����gg��~vɦVk�</p6����n��%I�޼�(i��a��a�8�I�Y�L���.���8�H)���CoY:��g���=�W<���b�C�@�E$v7��ϣg�0I���t�Y�'�w����QH)�s���~�a�v��Xc�l��l�@�+��z�h
,�11�XW�=��i����c��j��}��y�F+�~���t��b>�Ơ�,�'�xw�jm'�T�'yt��Xm�N]~�|�;H,���o!��%�VN��H-a�bzw ��vn�i�6�0��0����a���>���_4�����?~>���낐Rm
�8Ρ���u�CI�|�~�Y<v�S�9n�Xu�~���@�O��w��i��~Me�!�Θ9��l�%f0��N�T��z��;��>;��}�מ�����o��~bԟ���tݚa�Y��S���a��~��f�H,5�M0����)��:�Az¼�N&�8���>����E'����=d�>g����q
��/�����w~w�w���{���y�0��˔;��u�8�Y<��U�iR�&!^�|��<<�i��_�5�t}H,���d�QHk��<jL�gg��5��U�^߰�>�r&":����"���	�U.�7�zi��0���I�m�0���a�6�^�K~�ơ���и�̔g*h�&"�̝���I�*~a���a�{�:�Y�I<�)O�%O�0@�B)t&#���ʭr��:��Ă�'{�4)��vs���*~g���q���&3�+8�-1����;�i���1 ��a�'��CL���?C�@Qa�5�U_`�"����])�ҤE�[���;�x����8����q$}�MEq�j��;Vb��K���07�2[ ���b����nd6�J�'c�Jb[���Xn���c��(�[U3�I[�P��pr>灙��(�%\�ӹ��\�e��+��ʓ2p��ޏG���^&��%~������ELG�Xi�러��k"ϙ+<aSa��{ ���p<Vm&!^!��raPZ�0��3��1�<̇�i��g�4�׈bAt����y�}>���'�]�u;ݢ�eU���"}�	�y�ɤ;i�+6�Rz��ɤ�B�z��;�0�
��>q=�kRx�:�Xy3�4��T��~�M$�6����:��6��g���Si�Nzx�����N$�{��&���i�z�L(����z����jVw�u��4ԛ��M3��� +�وJì+��r$�s����:�>��i���O%�4�����PG�,m.���}�⳧14�#�\�	��~�:딅a�ٻ4��}ۤ��7�O+���J�R�?oY�*Aq���Xq:�!�6����L�+w!�����������׾��9�ң��o��=�����L<CL�{s ۉ>x�3�h�@Qa������<f�]!�
���<a�:Î~��?Xi��+<a��a�H)~�Z'�'P��Ϲ�m�PZ��g��w��o��ϻ�������Af0�g�V���]�$��LCHb�0�}I����f`~k'�ܷ߬�������m������W�X|o�O~aXz�uLd����������u���������>�ߛΓh�'�X}�I�+�'N��?0+a{��OS��Ac�y'��i����`V��i73�m ��Uw<���0?5�=Lg��IQ@�VC���u�r��=�߮�������I� �����OP���(m4βQ���w�@QgY;�7�
M�S����׌
��|�i?$�����³�J�%��bAx��4�E �0�3�x�����;���繝>׾��4�3Hcﹴ��*J��|�H�4~���!��C=�����g�y��Z�Ss��]d�E���چ�X'�ܳHz���a����T��fd���6^U�����������k}��L��N�f'֐P530Rq�R~B��`c ��3�|� ����m�YQ`o���X|�|k i�'Y�xs��V����So��L@]x~����������s�q(��s���jy�o4C��=D����(��/�Y����Ps��MKǡ��Y�9|-�k6�����Z�vK<���e=��z!�9f�9A7|JlM[V�t��x��՜6�$���eB�Eݰ��Z���a�����tv�mM�n�N̫84�)�߮�����42y�������q�M'`m�VTW}I��d����I����Cl8°��Ĭ�q�d�oX��q+4Y1&��Pٖ|���Xc5<���u8� �}�h���d�QgY+��{�7ۗ3���w}��|H.�;���a����]v��i������(+#���Èc��)+�0��vM�gXTY��[�mE�0�wT��Hh2~q��X�LU�Ӯr�g�V�Wge���ѳɯ�I:���J�������R��j6�A3��	�,8�f���֧_4�<��8¢�SFP����qC��c����8��f�<`Lz��W������������b�=a��
÷��C�J�O<��=a�
�Xi�N�D4βVl���>���~sI+��7�x��8�׹a�:� ����i����z���j�1hB�f���QDZ�4���� �d�16{�4��`i�m�����ɿ��E'�Vx��p�!Ru
�������+'{����T4�3�/�Td�_��D�1�1T��ߒ.�~��~Twl/�0��
����|�t���Y;�O�E�큌Z��)���A$��a��1����R���O�w	�P<J�e�9�i��P�OC,��@���*?��Sܱc�\���y?}T�\�
�;��RTu7l?j�Rbbbx���
�d�n��%ed��9�5�*A`h����LE �z��'Y�9��1�Ag�����1ѐ��E|��缨�9y϶}bg�v�Rx�f3�bo��4�4ɉ�<���`x�Ob���b��2�}`Vx���:��<��L+
�P���ߴ�f�+��<a��P���&:�?���x�%ܩ~��d���=�Ӧa��u����LH/��0��0�*(}-"��V���ɤ��'��Ax z�6[YY��1��f"��+<C�bM�Ru'ߏ��>7�߻�n����
���m�J���<9��U�p�p�AIP�����<�!P�w����i6�'����&e��� �=jze�����5a�a��1����G~�F��y�wv3�y[�;�{-g��niXܽ���X���������U|;�>��2�.��ͫ)�;Wo���z�͝�3��i���%	PT�*���DG��J5qQOg��j�Y�� (�bT�7gXi���Oِ^*x������Ƴ����=d�
,��sR{� ����i<a�c�O�}�0�¦�5��öDT�O�%O���|،�_O�㫏qG��R����a��X���݇��i=���$q�{f3L�
�'�Y�:�gY���.�uM��������a�=2b�kB���!��M�5�ϳp��&���T�c�v���I�aP�x[6��B��&��m�NZAvj�Ĝb�5w�X�\I�>q����L��0�*)�;�i�Xn^�]CIrcɵ𝎵v�9�s8m�옉��@�Dc�k$����d�t��"��Y�n��Ci>B���1��~a]��㴬�q�o�&�T��M$�����a��
�\����׉�)��/�}{^dtvv}�~�l������|���X;�su&{C��rɥa��a�P�J�S��^����r�C�
��c4�^1I^!�߲`m��=��q��(���߲2�g����;��ʫ�}}�b=>�|fN�|�i+0��N~��5�Ag̕���<E ���W�LE�k&�������0�3�PY��
��'P��8��������-��I�������1���\�}^gXcƳ�l��xɌ<嘋��̜�4��*$�+�@��T<��u�!Y���w�Y��,�\H)8ũ�����0*��q���nޑ?8�\��Ҳ6>s2�<��5>��f3l>Lg�5i�Sl��$hz�f�_�TO>����Vk�Mꀢ��+>�jM��
����1��a�<��m��c�Y8��x��w�n����2|���ϳ�R
K��>�m1�j�0��>N:O�f�;�4k�"�Y=O\I��ć����U�>!����� u+4���?��U@UQ���3Y���d/�o�\������8������� ��J�4o�h�1+4�0g*�E��w)֬1?2x��=I�6§P�j�z��Y�O�~a�b)� ��� �pz2��,�/Ő��p���?~ʳ�^o/V죄k*��	�h��
�����r��M�uM�}Y;����֎9B5
���2�s�x�����ԛ�lS[}Ȇtu���YT]��U�r,蛻� d&��V/�w0t|\I�
�9����"%���J�,+G�\� p��ѿ�<Cl8�Cú֧�,��*,�{�i%B���3:�$��6Zi=gcMw7`bz��lXu�0כ��LB���}z���W�ڿ����C=�G��͕�_�3������^�4�T��;�1 ���f�m
��S�ܞ�C;��2��nO�r�
�Y^����4��IpC�F�=�u�����*�;"D$�N�|SGf-�]��(�s� �B�וAy��s�wWiU���k:�I�:����������q&`	}�9�2��W5��Ŕ7{ם����Dܧ)ۍ$MϹ�"��fpl쨗'в��k�]����"n;-��u��Pf�k9,䢨<�ƨr��i��Y�����}f�T+�^�q+���"�dى��*׹>9�1��HNĂݡ��:�Qw�X��Z)E�S
{7�ӭc�Z�����	��c��g�g��e �d�WD#��`>>N]�0��=S�rTP7}����aޑ-���ꡱq��Kj��^�ԌnB��$�u�϶k"N����]<�l-f�E.y�]�p-���U�Ց����ǥ�OF��B��="T����jЄ7!�\7�K�9'����\&�'e�����F�9���4 ���X'�FCu����wӒSa�h�ɇj��qe������X. ��Pf3��4�u}*�Z�<Y���9���}�7GN{-��%
wϔe�G���v jMyG�ѹ�']տDG�����EÌ�ۂ>P*]��`��{-W!~�X�9�H�y�o��.*%՛
7�T�k@d?���#�QӲ�c��IW��*|���{�.���v&_��dD��E;u������	\�0��� Ɗ1Y�R�z%�w�'��W��ʽ��7����#�ٱ�&v_���a��I�|�w�bQ�X�'#X����TLb���Ѷ�KQ���{_������l])�4���pD��fbQ��B�6�QF���c_W���cI�}O�������L�U���ý}��zn�P�C��
�Y�&�&{#Ov=�5�r[6���V�U%�{�loV@���h_���|41��{�V�㤡��7��5`�*���gS貺��x8����)�η�A�ţ^��ڴ�ȳ+5u
���flq���x�Y�ٻ�!�W��ȐDk�A��,؊��|g�/_,Z��<��I�S�����R��𫨔���U���V���ɯ 0f�?:6�(�;ج>�V:��T��i����J���;4p�6���-�c�wt�)�1�ݯF�	-"fV���A�W1A;�u̞^�|����1�
	��Aۋp�N�������+z��7�u�QB6(/]��ud�Q53Z'u�]p�l͗������T��o�\-~��Dz<(����y��*W;?z|�*�pzW��MJ���uce�)��%l�f6`ņ���uS�Rx�^��e�z6x�d��z)�V\�>�5��rSZzX�9[Nc�d�
�U�z8�!gK�H����v��]�	�
'�����h4��(���:�����˩�<:-�S�w~/��"���V�*�J��
&��0��0}�)C!U[�9Sǳ:��h�Os5]�Gj�:u��*|�ǵ��1�C�檸)���>���F������g(��$W�T^g�23�S�Wy״�^���5@_A��H�	�#�U{�ғy���~{^7Հ���W#F&�����uct���1ӏ�LwCf�P�A�qq���]��8�\�79jf�a��3=c�ø9\:i�zz���	��Vʾb�xP�վ�m�A�&6����)s��sSe׾��&���@�5&4&r��~�=.h���p�f�y}A�W]j�����n��:3Ӟ,��a�d[����KvT*Grk�Q���a�������T��Cp�"K�
�^4,��؝d�6����Ҕͩ�ѿ���[�c�r���Q�:��0�y&��!�r��sE�QfVӨ���׹�T�	P^Li�B���b&�X���rSz�`�>V���C�t�*3�tTQ:���nY����7SkuL\���f���j��3�+ʜsh���'�z���C��jfm@{�%���%:�8�cEͩen�Ć�"a��<g���/p(,�h����o�α/�fWG��0h~�7.+�d��Jc`�w�o�v�� �5.Nܫy�W���a������L�Ո0�='L��7.�ܸ�΅�;�<�<v�*^�(����1�GM����ĳ�n5�~��gTS�Y�<��6'i�22"U�ϲJ;�G�Ka�p ˫��a�]�� ���W�_f/�Z�
S��w�=��:���e�1��e��iT�� ���5�%�vF�o�!��k��3)i�y������*���`�2���.Iw��������v "ux��r� �X.�9Ae�!���;7��[3��Ű�I��B�oT�o^����4������7�� � �p::�R\�R<'x*9�<�ݼ���9oAW���dB+i��ˆ���	s�����W3��l�:��<F�\��b�@�m��j��Mw�75�"�x���I���vFπh^mH�(+Ӭ]j��"����<ox��gs��4��i�ږs�e(H�E�ٮ�@q��E�t�m0h/�1!F�{�i�Z�`��(nF�NŻ�Q]�1�(����
�5�t1���F���8�¶�\n��M(]4�s�A��ᡢH�apB�:��碓a^ݛ/ݘ�H˒�`G5zvA�f�&��,�b6n`|��iyqA<�)�r�秱�57�?c��֭�>rkR���)��DZ�y3�BL�h��v����;��T���~��,>3��;���,���}��j
fc(L!R��{k���39�4�P2�Xխ���V��e�x��S��2�Ԓ����4�o�������3Zd����2qLM[V�2��ݠ2ݱl	i�)q�Ǣ��l_^�5��*@�(E���=���I�hNIu%a��/��P���GK`�P[l2Aؚ��;����O7э�)OdȕJ��Cj��7n�7ii�l:�����+��hT�#`���n�ŧ�|��Tr���ڲ� 2�۪���FS��T	��ݱ7�C@�$?^����LS�Y"_;���E��2X:��^iSYm@�7t��� �%�"���|`^��dd�o(����M ��}m�7k��
��]	\x�3��i�F]�)�u�,ޅM���]�T�I�/Uڢ��Ӆ����,/3��Ǣ�M�tm��)�wB�2BHPZɩ�hP� ӆ��k�<����F"����--`�h)?-&eQQ��+��!�r���F�S8�b
�D����.s0�Q�`����ՠ��
�JF�RWq*�[��T�J"���"Ŵ��aXҕ�V6�kTYX[KA*Ъ�*��ؑ�mD�[bP�����+J����
Z��J�V��A��ڋkDF�ڪԢ��Emee,���VR��QV��(��`��T�%���[e�(�1b�V�Q����[JYR��J�1���PkD�UUQ��ն�UDF�VԱ������*�b*%���mb��mJPE���Q��,KJX�%h�AF���R���
���*�U������,���0F(�ڲ�g�����xA> rߋ��E�[j�T��6���CJ[��6i�M^��F_���A������F�O��6_
�;�,��ꩍ�G����	�6T�He��͠��kc:�G��.	�5vxGG��0���X�bׇ�m�+���^����6�m�ً�sq!�F�_�f�J�4�Ħ�w��__<v!���e�K�.��Y�dKi�����>�L�T��S%zOXU��;�
����qL�ε��M%9�i¥�fX7��T�Ȃ��1=��jw��������^��[���^鞭�G(���aD��c��N�8�[�w.n���Y���;@�a�ɟ��X"���&u�UVh�C$�Y��`�1�8����^%ٳ�l�ݕ.S�&Evz��s;�ȰQ�B�=>X�P�V���僮q�B�s	�a֚�;���x�(cʾ�/�����s;#��ꉐL�����>C���T�-�����qb�E��cMr��z�.�ʚ���붎�c]6�]�P�t�/$�E��g�\L�uY����Y��H|��|�q���K- ?|ジS}�ٍ����U�1dK���g�;�><f�r2����ƫwֽ����=�ܝc�:"�ޡ�`�0�1�����Q�t%�����A��W���pp�;W��rN�.��N���ǎl�*@h�U��m.��K1�d>�;��=[��Ò���!6��44�ϫ���꯾�6��'x������E���N�IB�l*\�=�N�7Qr'��Q"��8�����	~���z�R�P\xe3KK�Υ�B���=4���)�ԧ���O8+0;nU�2���]��q�H�9�R"p�B���t1���)��U��\[Ɓ�]yASu��Y�J��pHa�ƅ_=]R�p�*�x:tv�J�Py�q�W/n��"T��G3�wG틘ɲ�R
MV��A�q90[��F b��*I�O��ʙ�<��Z�W)��w75ų��/۵r������:S��ܹ��b�Q���OlN�b(�*�wĎ��}\�fҐ{'������5'=�")	0���&.\ۢl��$T�<�
I�G�f��D��W8��y�����#�Y0�*�}/G�#v�`^q�Q0�-f*y��
O+����zjOӄ=�=��Ucd@�1�4��&-;.'eD�>YP�SX`c�5��c��_is�{<�`�4w��"����1۫��>
μ>��:C=i��_@s[U��N�=g(fҭ�����z3q�'���V�b���Xt���n�����ɱ=��>��fTu5,,�ayl��䉡�v�^ֻڥ��;���)�FQtZ��7I�4�Ұ��bo9����c�p����Z����u�sC���	��>�����^�Yl����}�/Ȱ�w��hNC��ŚȘ��d�Ƅw6���Ssn\'e��Q��1:���z�|ٳ�l10,�򾚛�������Kd�M�����)������ha*�&:����z�	ɺث%tzM?���<+C�tY��ܨ�����ڕG1b�"u�+�&�#U45�[���T�eöF!]Pǃ�ۻ�~F@���'� �c���2��TS���j�؅-�*^G߭�{��b�Rit7�[k�O4ߵ`��ZO�����f���Dƺ�zT�� Vg���rÅ��w�^=ž�b,�j���974��g-�]z���5<6���u�z�ٚ���:��(�6�ɲ�eէ~S�lc��ה9��ho�b�ʬ!p;{��C�u�,�S����|�Jc��Mɧ�:m��%�c3�Xfk�)v�Y�`N7op�jefp��Oӄ��>j�Q;*�F�/;�ۜ�U�7���(�ni:���>�!s��# gX��W�ۼ��D���622�	2��5����9V��<�*�F��3x�xz�Z�&��ҡ�R�SY�Hx�Q�s�g�˞M������^֫LEk]�9�V�wI�/7^^���\3��"u��E>]���M�ͮ��շ��_R{A��Y�l>0�=�"5��y�*u�Q�����I9����G�����m��ۓ��?���X*�}�Y��s@�<~��)��э�x\�t�a]\���}M�v�D��zx?�ʍk�k�>f%�<�?��^�ef���x4&��]��}����8E�w�{U�����%���������Q�ŷ�/G6Ԙ*p�E�^tX;|4d֒DNK�����Q�V�����@W:�E�`��[�k��`���L�v�H���i����I�/�"w�=쌉�ʩ�������mP��W�nx�7�P���bI�Ftr���q�*z���ڜw�MS��a⽜���Z��K/x���N��{]˰J��&����[J��':S���"+]x�<�Bຨ��ay>i׺o^λL���^�]�Wl����Gdi�P5��[K�x4tuܨ������ ��ҧ���覰��V�/�G��_�ב���]Ѝ~\��!��W
��2�)R*.�u��9�b���o��u�i]0؃�j�N��SpZ,��j��u�$`zq��])��>�V;ޓp{p���\�/}gq���dj/��y[��,2GZ�YT�V����=ڐ�\.*�,��v�t���3끬W�2i&�ݝ� ���n,����/�1��9B\ݜ���DG�s��y[����� ��Ӯ�=;1��I�[f�P�A�qq��l��$g[��M�TC��ݛ���=q�����4��裡&�ʎUӳ=��(�N\M�"�Z]][�Ƿ��Q�PǑ��P�b�"���Y�`�S�9���#�r�������M{����um���k�fe�KUO���kA�O��q�[e�uK�� 5���r�bu#&�Ugcv^cyݩե��%t����
uS��t1pM�����==��.�|��-�Ǽ>k�ߨ��"�qz�{/��ה���6f�'EL\K��8��2��)vk��[֓
U>��E�)�W(�b���U͞�q�F�s\+�J�a&jr�::D&p��� cQ�F,�Ss���Ǡ�di��Z�t��I1s����.;֠�7��T%�̉���jM{��n�,�bzW�
�f��[����#ۧ�J�,p۟\�@��l��Uv]˛N�||��2��(�;�ܴ�;�{i%�g��.�Zשyp��Z��01��%:�Mp�}����N%�S-i��I���������Q�ݫ-��!G�U���G9=�v�Wy֙0,�-�}���<���e��]�ӹO^Z��(�.+�����Z:g��Q��{y��=�{�r'�����\�v����<�:�^6mPZ��o:�-����.|}\ŏ���O��������	N��6�,����cPS7C�<�&�=V2$ǅ:V���X:ֹB�sᑎ��tF�Yl/!�E�3�;�����j�c����>N��ƨ�U����-���W=R�$Χ�ؿ&Ϯ�t�����VN��:��գ�����r�w�y���n�s��Y[�o�!O�H��vR~�����p��}�ٍ�9*L*���%�b��O1'�'K���H�AهC�u�ˋwI&�r���<`�R�P��}'g���|�ل0g]�!o��0��ʿ{�����/Ǆf����u%_�puS����Zy�5p���2��Ot����.�r�}8�f�1���\�*�tU�@�q��m6�فb����dXs_pH�Y�O�����d�9DĪ!:�
T/ǂ��z��Ә���W�B�gcz0�+��3bD�����dJn���a@����@b��*[5|X��;؂ͤgxF��z���49�h��\��uү��ܹ�qA��Th+�+��5��N�_#�T�$N993�����Zyy�D�7B���=�Oa��պ��c^�q�VN��)�z��S�F��P�H���Yr��D�س�����>T���880aJR�G�N����i}<o��֦��2�sT��颋r�<}��*eqO��Vo�TƷ�����z#���a�v�g��'7芈��f�⧣�D$���Нd��c7xC����M���&��Q=Z�Z�/�Q�L�^�nǃ��w�x�W�{��	�}�*l-�V��B��*�o��p,-;�E1�ڪ��)1�5}�t���xu���lX�9b��X�'�SV�P:����1����83���%�lO�(<%����Jɍ�|�7�p��մ=~��~�>?Y��苈b�EM���<��Hx6n"��;V�� �u����<�q,:�!I�Yl=��˱��]�={>��/H�1Z(�CzhAY�p�����{�%�Խ�7xW �
e.O*�&:�ήZy������e�ܰX~��p�m�`gx�k�x�N ôa��!Ե(uy^Q5��csV:>�Ё�����V۞�R�7�e�\�X�����t�N�L�
%#`�qW���!�[�:EK�����}-}�w\��;��޿a����P�4."�WG�5�C�y�=���.�13s����2�1���ll}u�7JX�w�������g&@y]aQh5Y��he�:6O:Mm���N�N�s�chr�"�N��u�����r�np�%���]��Lf�kЅ��ȋ�p6=�wc��_0r�aɻB^�.kk"[���{�6�f�۞��y�Ҧ�ln��{ވ�f�*m-�W]��~aKr�akZ��g���V�O��|�����\#�x��Ƙt�ƽKv�,�[�z�t]N?:�U���&ʭ�V��I׳���S��Q���Z�;V�8�T4�uuJq�.7��|�G1�F���)�ضa�M�Tt��B_{��}a�`�tX�@[]�+�ۥ��*���(C8H��ǲvU����r�"�9�<EXsaצS�%�#/uf��55k���s�H�~��:O�X)"!�d
?N������!�)Q��z�Ժ˖��.��]�8�g|R��/���&;(b�H� ��Yd':|Y]�l�����WZ��]��ryv�(�݉�8����'+J�GE���V;<�u�'���#R^7Ӓ<9R��-��LCon��>1��jΨn�{{L�a�Tl����4��r&����q�Y����>��������Ԛ|��*2�&�dM���2'�*�Cʰ+���l©���3��t�b<5����X`���w!p\����||�C��������&��cy��)鉠�(+2�Ⱥ3tìG�]]]�}���jh�\�UƖD���G�M7ܝ���4d�KQ\z;�������Hta@s���Ar�hĵw�W��!emHi�;�1�n3Z`��e1��;^��4�;�é�l����U��?�#�����^��#�aK1&���
�ю��p�������s��>u�D��qɳosx��M����T��8o~�6
�z���BN�G�»M$5��ηn�Y���(Z��Ѥ?7NT�(��f�v�%Bw8T�B��jjc���c2����X�W%`��S�3+	�n��'���1�����-�7�d\#Q3��'�@NĞM9��ly�~P'B��>]��q�./f��:r��鎓�O��6M��? ����uus�K5ʏ�@���!꼏<hᘠ1��\�Į4�"���M7ʺ��*�����8O���^;��g���2�����Q�U� ���x�G����3{�pYj�xb�=��}�+/���D�ηK��zM�1
h*�r��5���R��\M`	�fD�(l ���Ձ:54;}�Y�[��:2C��.VE�� B��ەC髳�S��r����!�jٹ����o�zA��C�\+��4�;��>�=1�F��3s�)�v�8��ô��ǋ/zV�"�L<.r�\&�޼=Q�Wd볼Y�/z�]�h3J�tU��Q��6H���X(9�eߑ��(qo���ΐG���w�D9��]\���`�[�5�I�>�^m��O^�1v{�nl��������(�J~�ﾽfv����Z"k�]9(�1���LBL���::D&p���p�]���Y���Id{�ǞN��s��{E;0��q��[�fX7�E$�H���w=�n��N��Nh�au�TS���"�؃�EZ#uT�U�Ս2��/�^�o���m˝�u����2cr*k-�s�q�$�7��%�qѺ-V�񤍇�Tt�o�b�Ơ�^���`\3���D��ء�yp{��4�Z��bW�`[=V0�.c=YJ$��l��% �Tl��sK��Չ8��W�6a��a1~E�l�6�j2�ڨ����]�:�<eW��+}�k3�/]�e냝�:Ct�Sr(6� X�&Ϯ�t���`��]N�^���8e�<*:vpve��n�ؓʪS�ź�ȍ�=�o�G'���U��s�AU]#5KLRVB�-b�z�3�wa�|�J
t��oGr��^���rmC�x�R�� �I��.:�.�;�V闅Z�ngq�uȕ1��X�%M�lB��SSF��1x����MŻ�K�y��uA�+m�y�슂���U�Z��Zp�g�Ϋ�QJ�;$�U�:��o]�#A��g�����CխMm���^bv�"����A��.:=a�A��ʶ�7zd��$�ڧr��X�ٌ�R�w��M�}��`��j�\K �4�V��w�WBA�n�2�9�a�h�q>9�l��	ov���_q�f%�;u�����옌bYrWE��A�%��gm��<���Z!]��+NWc����սɄT���4d�]n�ƕ�.�>�"Km h��C�溊�F�J9�	�XY$�6�b��St<^��d�E,m�nY9Lp�,k���k%F�t{�֌GRv]�TQ�����8��.�q�3�u�/������o�h�<t4H�t1D۾��`,M�SC�K��N]N�ލ��ԩ�`>IovM[��<�����!oa}P��܋���f�P�>�;�'o>�Zא�9Ҍ[��9n1o\��-�l74M���{':Z�	��}���4h�٦�E�Y���a������Pƥ�mo3ڢ5��:�t~���SA�Aym�b �C=뽃�Л��}0�츷1�uԚK�6�WS�ѵ[S:����嵎D�
 "+(�Vr��3��s��w�],�&���_͔���&��5�-p���{�puϸ���#W;����0Sf���A5 S�ms�\��&����|�����s��.L5b�b�������lo-�j�ӄ�Y��g�f����]9�]k�T$K#.��ҹn�B]�vsq�"\�/+e�SG��T7�%���X�%6y �t�B�1J���a�^�.貲��v��P(Q��f�M�)�,��B�`�������P':z�ɘ;:��Q��;�6�6� ��������<��o��	uWPE�N�Z��*��fv\�1鼴܊�7��V��R�+m<�)�%1�Q�q8Qw[£�ϕ7C0pgk*�BZvT��IC���ٜ�:�*��r�ܖ@ճ�˭T��TZCX�I�`9���)��t�m8��2'��8Q�N	J~PxFtn:`�����np�Xe'j��8�;��F{X񆠧�b�����
�qh�082;�EX���e�1��k)`^a	���4r6��ORY�7<M�KvN����ތ�F-�Yy�`j��\xT��3o!��1t�8��'�U݌�H�bЍ�hf��Ҳ�Vh�D��ۨ�����I�=�st�T0.D
����.*�!l�B2E�sU[��6��AB�y$�,Ț�����^����0g���6�ˌA���D�Y��/*�=��T6n��p��M0����^��ޝ޷zx4��r���;���P��+�Vx�EF>),�Xՙ�__������-���Em��[
�"��m�Z1[d�Z��+R��UE��-�����1-i�R�h�U��Z�Y@m-��%Q����J�YiT��Z
(�ekjU��TKiTml**4�ն�"��Ԩ�YQ��,l��Z�
6�V,���l+X(���ZP-�[eeb�6�
��-��+V�Q"��PT�V�l�"�Db�Z��h��b����
RЪ�l�֍R�
#Q��J6��DX�*R�m��E��*T��+m�[Q�VڡX���P�Ջ`��iDJ�Q�*��0D֑E���,���kl�UmJ(,��H��*
�*�(��VT*UEQKV[T��J�J�(%�h�Q�)e�+ak[`�����Jȱ�E
��ؠ�D�(�h
���3��SW��k��S�sw�0�;�B:sX�c8E�z�E�vzb4\^iSs�)�u�����0�\Vu�-w��~�'^ux������;�_YB^�(u����/�lD���T�u�-Y��~�LR��aqβ�/�F���[4���{B�c��C��GX5�<;g�b���{]�ɜ��;��e�7��gn9��3-)���M��}��
�$�s� �����N3���M[�����g3���;���z��oNQͿ]v����->^N�H��)��ٰ0��N�r����o�b��M/=ua�͍����m�x;�"
�5>��%ͺ7fZ"b����:�cg��]�vܻ	�*Z}���J>b���Yxr\��Z=� 紩�S�r�V�d�wh���ͭU]�vb��Q�zx�_Ȧ6����xp��｡�W�~��N5��o���=�1�yb�1/���򮜠q��P<�뼪;&�ᦫPɿ��7�%&�Wf���P�q�"7��dh^r���.>�gO��9����H:��!lc�pJV�gW�V��/Dwo:��KL����0��=N���7.�1:��g�g���.�c� ��}j�ݞO\O��2=4xjJ��'�t�2R�~~� ���H��?f)'=�C���EX����@0d�]�-��(��PïU������+��7��ڵ!���n�Tk�\T�8]�2t=T�C��{۹�g��V�1�M�=A��U}W���>���^�"�B��O��P��T&79��oU�ի������j�
�9{"��݅�by�9�$���K1��iT�Z+>U�G�j1�#��e�3W���%f޼]�m�W%���>Z�Ɣ��v�S����|��4��9�z9.�h��(Ov���p�|V����H�s�P��Tߨx��h+�3�1���X�0.��k�Tw�ђfu|+�CL����I�Ǩz��Eæa���bF�)>��A�j��g�OmwJ�Ő��r�yT�:4X��`�ޟpuY��x��9?�x����`Jfⴰ7lOnu�d����l����$SD)3�ҸS�"�]�3��/e_Rt6�P�>�n5Wj�Q��T-Z�'�,90[�thDm�S�����p�T>���;lǹl�����������T��`�H�{��s����+�R���0y��Zb�)�#v�	e��'GX�70�$z�ٹY�扭����ʧ?���A�m�)�떡���"@���e;.Ȣ}j�#a׀�LN���Y1�K��t���9�^[��[��1z٨S]:�`�ɫ:�ђ���@�J��ӘIغ�;��-b����#.U�57�{ا�j�?n�o�^8�g;vh��2,�A�Gx����i�eC���t��29a���/`���Kn,X7����1wi6�u���B��:&y���¼n�f�zR+�|e��Gx�s����[��zE�n���晧�t��Q*N��q&{p/�;�O�ӗD\KC �q#gb_U1/A��T���f�o-A�Kͭ��4�7��4|��KȆ�H��������<����L�Y� ҹܼ��n��*ÖÓ��.�2�z�D#���������97)����׎�S}B���^��YƜD��r`r;5~5�	Ю�Q;����QA��zX�7��Vrz�z=�wո�%}�_t�8�Y�sɔ�|T��#��1�*T4uRwJ2��(N���+�ֹ-�A�BA ts
z\2���d��䉳����+h�{WT�1�QV�Wb��Տ'�jjBʡ����1��c�wB�a��F�g��(	ؓ���uQ7�^s���*��v��`��?Z*n�d�
o�t���.o�t�I�}'�pٷT.<�0�Z8$���#7RZ�^<�Ο8
(�pMJ	e���cP�\:iݻ����s~�=���tr���b[b��)���نjݷ֖C��h}d��e�Z`���;f�˒�/}�r��$����q�S��}��SΣ�Ҡ6g�~�˫�}�Յ�8�a�*L��/W����1���Ҝ"$~t�Ę�\���d��Z1e��;&�b�0��*:\���tOͪ��f%/�;��[sA��B��DJ��@缣#�
[B��*���G��Q:���{�I�/f'd�¶Ǩz�5䮂�_w�S�����髳�P��ݥ��u�ZUY/����Po�q"�y\�-�y'�q��d��==TQ���Vx�|�⪏�m�yp��Z;��P��z����j��|й�O�N�����P�DWf�z'z���-�El���L���>"2V\a�F6�
�h�����I��/���{��鬨��[���s�Zw�w��k-
X���VMk5�H�Cgy�3�(z�9\��}�W��:��#$@�^��S�f7d��o�)��WT���FLa�2��Cu�4mMDs���s?b�b�`��YћwT+{y�G,�r��o:�����k�ҏ��dI�
6z��,�W��e��%W2@R0�%��A�z�gq���v�+�?+|���Z��fm�,��v�r�Ͼ��\����W$��,������S@ ��Cؓ3�E�Uo��o��AزVu>��a�J�ʎO#�����
��VLM���c����X�Ȃ|�`��i�T��KB�3Ky6�2tqlJ-1�[Ra�D�oEu����fA]5������t��b"��!�q"�7Y
�ظM�]î��7"���58u�V�ᣢR���<����Q�9X]�c�U�����j���W�W?}��×�ˀ琁��*�5X��`�7rGAd��.Z�X��g|(�J�0%D����e;S���B��@�R�:NM�6�1X�\���:f۫�+�F���h|%eŲ�xO����L�R_�ps��^|z�3�-�mX�{^�s�3�V�;u+;x��rUK�84ñ�)�:v|8��r��5���P�a��7��.j�__�zr���b&�I��k�5�k�FQ�l��Q}��ju��iN�Q�%֫�~������dAt����3��&�6������U� oo��_�^�K���|ԩS!3o)��<�绑�sp4����qA�]��:��wy7{���M|������V�E�͏u�/�ȉ��s(|e&j}��d�
ܸcn-vњ����ڭ.`���;�$]���[Ĳ%�jZ�K�+G��bNj�q+fґ�z�u�R�òwP����Ro���K��i䥦�bWBu-!GO�W'����)�E��6�֩Ԙ2����W7�;<۳-W���ǯ���*�mϖ��|�V�������2�d}N�`I_=�E�����jx��^/6�Ed=�s����f�I�/+�� �*�֊ckڪ��@�=Ƨ�Չ+�#�H��mKT0�U������Q&ۖ'��tǢ�;Z������ѓZ��e������v�_40-8إ9p����D�uz[���	��y�&���i��l���p%R��fi����=@��IL��s�!��~4{(�l.�>�E�U^.��sݞ�h�B�$����� ޓ��]J��$:��B�U	���r]�V�'=]�ƬP����s��J+o�߃��_��˩f+k�"��gѕ�Qi5�¥��J���Ǔo�*��w�n!�ٲ�_Ҫ�'�h#��у(1����J�2�� ��U���Y���=v�v]f؅-�*_J�[�����B���;�I�3�T�=�U�g�Sй�����N{��gH
5Ǟ�1l�$˘���I�|G\b��a�q3<�ؑ�
v��ˇ���ྦྷԡ�� ˪�ns .�J�����>��=��琡Ρ_uEs'��q�ŴD� �Ց�oVc+���N1P�r��<�ɤUE3�3�smx$֑֕vV+�v��u�ljto5uY��=����-
=,#-�"�={�n���>�_N���{z؜�HYb8��r���}M��V^�Y��N�8�M�=ݽQ����Y7o(�ŸU�����y�μ#P�06���m�)�>����Y.��.S,�Qgޫ�Rк���<y��
�bFT�MDZg��9�`���eM��8a\���N�ŭ��e�R��J�q�x��T�� x)�g�2��S�B�}f�D��XƤ��ٖ�tNє�\=C+��?M,���>i�����ށ�%���u7k.��.��0*6�ͭEDߥϋ�ZF%W��ȐG���M��.�+�
�k.s��#��odS���74����*%ɾeĘm�������T!�	�fr���Н�S��-d����b콽����Z��4������+u}�>����A��^5!B��+�}���l�u4&J�������a�x6LVS�~� �vp��,��V\��||Ϟ+�ɇ\(IY��Ճ�T�Ex׆@7���־4�ɽU��y��I��(>^{.��
�:���c��md��z��{Ð��zzF�q"8:*�.��Ǝ���Ί'ٽ=Y���kx{�g2&�#}�������m�Z�wA�{�l�����W�M�}�%:	��ۥqo%ŝè1j*�'�����s�HsSb�=X/�]�SM�����{�*.{��[s�v{eM�(�{}���v�xpm���j�ٗ���|x����EU�3HCP�uV��*n#ϝ��ג���r#/~|$HC«��+�'���
�Y6��tۨ�x��g���ߴq���=
r{f����W<J;S�Lg,Q���������L;5�j����J�Km�Z×&8l��75�n�������V!b9[������yq��ӟN��0��	dQ�iO�:�/ҸtӸ�}=B�4\��QP�����q^����3�5E�D�w38�a�ە�[�c���R���N�yS��kGep�JV*�p�٦p옄��G�GWy��\=�>dq�V���5H�Y͊��G�R�+O���4��q�e���
���������{PE�Kv�l�}{��{� ��q�	lp�듚�)�{1�l�C��3�A�Y�v���ÀR���Fa� g�����CWPu����x�_�;�3"�ׇ*i5VQG�}��zg'u}�Ňd��U�G�<�����x����@�{s#�@S	k�]�a˭e\�������b��  _�|Z刯e��f٤T�CƬ�T���s�x�X��B����)�(nC�
'cN�zS�c}ֻ κf�fOIa����尝�g�o�o����j=5�RVL�6%����B�U��62{$İ������cm5j)�����y<�A%��%��.�s��nyvȣ�y��+�����m�;"�^o���J>Z6P6*�V���)�h�^�Nc/N\�M�������j�4�'q�������7��ꌑA�ae�Z5��ȓl�F�;u�FUv���Ya�n52&��T� K�]Qa�)sL(i��\c'7͝��~}Q2/j���^ �V;>��7Y�W�o�ZUD]��9�'�(&�:��M׋=�1yY��Bs"i+�>C��WV��T���7^N�0C���L�ʅ>�L���+��G®~�87��>z}�Ւp�EH5�t�_F(Ţk�7U�1�S��Pq)\a��M;���`�<�==.�wS�՜h��,���)�)l�N�8V�3�Rϔ���٥�Ծu%U��XW*�N������{���M����=Ja�U`�z%�b� ��
�N�FJ�T��J��^j�+��������S� �9�/�Ž# c!���eP��!LT�0��Ր��������7���;��Q�8��_�.|���0R��H�d�y`�m~�k����hu�5�O��\�:���� ��\�m�&s���AVh�X9@��Й÷K�����=(��s�V�{�����5f-�A�Zz	��jy�r�؝#ڲ�Ht�~/��ê����f�
Z&�M�9�t�-��=���m�Q��}��]o�m�ϖw��B3���Ur��&\�P�.e�Pb'L__"U��y8��qٔkoT��
�zS���"��M�N�#eX3��OGg�ABJN�|�7��i�n�9S��2n��b��+�Fg�~J�G�1�*t�v<�?*�I�]⍷.�"���U�lR��~c �}�)�!�³�E1����D�@EKB3Iue��=�ۥ1�;���ڨ���q*j�8�ou�*N<>��@��;f��xo��/+OA�s=+ͼ�{%wI�d�)Nn҉\N�`��>�ڼ��T�=������X�sitY91ʪ��W)�h���:X.ձ7���L)���Wm��FY΢�w���w��'6#k��ft�o/b�:����(�?� �����}9�!�pV�Bcs��Kz���u��u�w\o_��k��b�u=��������x�Dz%�FW�ME�`��M«>�>�q<�$��A�)V�>��oXZl�λ��x��Ij��'��Im�/�H|��b����uZg�ŵ����
����̾�U�r���q���v��]=��g�N�g�w�Wv>���u.M�uOx��>��$nV,��w�cv��÷*j�W��T�������O%�j��r�;�0����d��$�BH�0j���U�]�J�M��*���um���hX�]�h�N.�0�A�P������ɸ�;�=Ǣ;�s�9�Y���E�/���]�s9�2���w��V��ћʶM\�1�l 6��P�X6��3Ɖ�7WQ�S��M$P������3S]P+�ת���f�ͩ����o�v��9;�5��r�����- �Km1�t1�f|8�5r�M��N�H�c u���L���"�c'e�0�,�iK���_I��F� ��(��Sz�kV�����g�/z�*�Y]Sf��CM<�J��M��w�{�ד�sh �y;;��ӏ7I�t��T��x�uf���6�fB�#�F�{ܞ���]:�5�@2�m�P�!��c"��T�V���Nl�B��@qŵӒ���5�f�V�B��9+�u��GϰśOnF;t֦�q����.٨����e�=�z@��6�d����ӄc���\��K�-䬣8��W���Fv��w<;Rs{�,����;,�%�ݒ\{i$d�vc�i���,���+^־Q�N�������Y��mD���x��n��J����/�΃���fbF�s��i��v.i���.�N��%8+�Í��w��&tzpgg�9�-�λ��fɟ!��?�S�A<�,>S��{s486�.v��9��.�䤫ܾa�\��yk11�)%�Æf����)�g:��Y��Y�D�Y�@�s��紉��SI�ټ*�-O^�ӻ���{l�=̹:��Z������9����&-�2��������P"k=y�^�*ڸQ/,�T\U�/Sq����]�;�S�X�n�x��+ue�-���8��S�~JpIŴ�Vl�鱂���@˼ܜz�����,wa赧����:�V�+�4�h��h�L�ݫ��2����|���t�a9�:?��7��$��7=�����Yh�p��-������}�v!Kϸ��'l��jݬ���O4!�����x�s]�_B��;2C}&���M��As�p���=�$��~�Pĸ�ٺK�ɴm�ǰ�V�dY�G���Wcos4��tK��$�����|Y/XR���D�5�)i.�<s>!fg[ڠ��V"n�t.<�z�Ê�x �E��W�+mg�4�ʖ"��#K�J�٘)$��af�����T<�:�o����:�]�;�(��Az�8	l8]�7_{H�b>���ų�m:��KZ�/s���!�A!͕�ace�Iշ�_SΘ�Ms�=n�I�5Ir(n��t�CGg� �\s���MK����cٛ��3�<U0e�����j6��̗���A|G� AG�
X�-��E�J�E� ����m���(�%��V(��R�ִ���b�Q�B�UZ�+`Ҕ��J1eQU�+XU��m�J�X�
���im"��*R��jV-���*��T��"�[am����
"�#[R�R��[Uk"��mUIR���������k*ZԴj4����imP�)h�e��V���R�����B�QmB��P�jEjT
�+*X��eB�J�KF�V,��R�[�ж���J��j�B�e�X��T�"�ImDKE�F�m�*�V�Ume)`���-���Z�eb�؂ԔTQh6*,D�B�֍KJ�bU�Uka*QV
ʔh��¶�-��kJԵ�[k"�1�����ڪ"�ek+RVX�kYU�E�E��i����T)F��P�-T-�bVTh�JAB6U��UX����Dm��P  �G��n�ϳi�i���=�9gf�Q�=�p+F��W�Q�^��ᔙ�¦��`[j�K�4nG�3ܚ��Qfn�Y9�[�;��ٯkyK� �dW�д��!ˢ--;ܶwAxp�Z�9� ��*sy��ˬN�ٮ��\}����V�C~�5�*��*t:�4=��k�������@�@�.�R.�y�c�!�*_J�v>8��d��Ai<F+�P��F�������d�y�]RŅ��l�/�
NS1�N�ÿ'J���n�\b��a�q~y ������}	�`.�鋗#p;��.����@mT\����W	߸<���B�%��G�+#�{��S=��z ^��b��#�Πl��#i1|�Lv�B��O�tル3tT�	mew�����n�%���'G�,Z2�%.���o�i��*���-��OG��ۍڥ����EXSn��QL�ҿ`.@�7Γ��:)=�ju�
'��;7�M��k��K����.L�����c"L�Z8�hn�U�Ӛ>5��փn�ժ���P��L���$K܍���𨌣����}X����TG�=}>�&r��۲r��7����q]��L~��o?Pu�{%wM����LϽ�ɯx��J�'.����'UFFhL(AM��[�H�x��w}�He	㳏_&w�Z�%�l����[�;2�lμ��B��k�C/{r�q���X7פ�Zk�����x,�Ւ�����c}no�����r��}"TC{��w��x7++;"���w2�a�V;�f6`�K��k)`� �wN�Y�EpQA�k��6��=��xs�-�Û7.}jr!�;Z��A:<�t�Y���Mꮠ��_>��2-��pg��rQ�J�c1�y>/�\4U��[)>*E�u�'�6c Q.r'�D��]] ����yk�=��J�0�IA���a:r��e�mX�f�27,y𒆡y�Ylu�,�ue����-�`ĩr*.�u���� �w�c�0�)Ȃ��!LT��ݝ�j�N��Y��\��yc�:
&تai�u[*napSְ���A˗7�:q�	������f�K�n�����\��F0�N@�::�D�zuT{]r�tӻw��!��-��4�5[���s�
ޫ�9׹?B}��E�PS����~$p��]�}IPC}�cn<��������˞�0Z�S��·�f!I	6mp.����
ʲ���u��N9���5�t\�x�T�ޓ��s)R�Fi��ꋬОk�eK�����	�[|9�E�4혭�|�X���U�9�]��a�ؕ�{�*Rc�&x5��|�dD�x�qd�43c��-� ds��۰t@wEX`�{5��NP�}2����|�h0hz�tҸ܂ۥC��J�Ө�����i(N�j`�s�^u愇^�J#�nςd��F�ґ���+LfD��1��S��Fs6�*W�q�&k�'e^�����xi�z���k�����n�ydq���vjN�1�!D�LԫN��	�٘��Q�=�s��v*�6�L
��Up�����U��;x��|����:����++'�=�{s��8ǽ��5/�x��|��b����t,xN�Y�Mzӓ�z!Īp3d�N��]Ny�:fa
�!q��~ѳ��Y���;@�	j83�o䯏�X]�k�zI}ޖ]�H3��Os�S��n�zn��Qu��Bھz�V1�ǅ^��.�%��:�8}'��\7].�	huQa�btX�����'5��p�� í�\֞p-tUv�y��K_P7���x��F]��.AI�A7Y.g�o%��e4���n��y�M�����D�7G���X��Q*���yP����Tߺ��
������t}=]��Yk2�U*ӳBtT~�*�
�^(��c����8����%(f�hm_��m�˛���SjX�'e�Ư��t��_uW���N��4��^!_��'�V���o#��wp��^��1��m�3�1�e� &���������|��Y�Ǹ�������bȗnb���Pq)\F<}��sy�ҧ&���O�`��۝�=����@:q�V7�P�֎����R�e6�����^:�\8��Q��t��a�(�A�	���D[�t��Tߢ_eT��W�<�l�\�g*M�(O}ж��nb{a��΃y�Fɽ�a�]x�$[�1Z3ǩ��A}~>oH�ȗ3�����b��c������2�yW�<�ߚ1�=&b�#�7T���y�\)��P�'�D����~���Ku�ʊ;
�j��p�ulU~~%�a.ze�g��r�a%�܉���T�N<� ��lW��MkD�&)��U�ҝq	^��eK��X/Ğ��ٞ�f�^Էj�?'Y=67C�O�	��lx�Lo	�N�Rԩ�ӭ��Xc�;{kZ��9uY�	�c:��7fd�y᪎�ŝ�����~����5-�|le��.������2\4�f�F��ЇQϲ�[�E�~��E����(i��yJ�������n��2[�͒ٶԖ*l�/��v��ax��`��bx+�S�My`����y+�a�@5���-���YD�S\���I��;�*��\�+��V�盋F�my�uwG���81t�H�HT�r�Q.R���c���*�����^�~�¶,d������q)٦:q��6�4F@ux"����to�\��9��6t�{�ĆÛ�����;����S�uYlv�ܼ����OO��c�׻�/`��\MU�V{V��0����k+�`w��£C��=�/i�T�j��_��1_vb����qاg�k���vtr�`�b:I����AD���QiQhs��2� ;�q��7ˬ�>��>��H*^Ө��[��<j-��k�wLt�o�s���L�뾴����'Ӄ�m�1qR*_J�v>+B�,�/�\tp*n|g�(g�-�O��/pmZ�Q���(�wq�����S	ҘwqSxҺ���K@�������U2�--]"�a��'�:]H+�3��Ҧ�6��Q�:nx��t�����nr����2r��iq�v�d������D�1pG�a��l����rE1�P��mS�s30�/�XԼJ0��m�2:{:*�:|g��P�|c#ƹՠ��|����ɒ���]�I|�{wM��7G��6���"�=ڳ�"��[���TwKt=c:=���_�*3�!�z�;��g��y{���uhr�ݐ�۲e��3�-�3�����0�)$Iv]ZPY�R�	xlJ�S��T�Dl4-'{���:�1�����]z{��\m%�EK��=7�`��W����-�\��f(�ӳ�Ll��Ys��Pڷr�K���E�I�ŷ`��u��dI�q�ӣf��m9$־�̛��b6�{�N;�R7'$˄&R���*��&&j���/�W����)�9�y��Ɲm�T5�薌��!B�nu�ͤ��Ґf�P�5�{��.�iD��T�w�=��.|������ڼN�$w��g'�m0=Q�X>9N^�c�:c^8'۫�	�[�ӽ�A�6��p5ּ%�Nv^�,L�ͯf�:��j���L(�Zmqa�sWN;��ؖ���]���M��|�߶r�f�Lz=Ռ���c���(��]SLy�3����ND��oCT���Ψ�ݾn�|a�>>U�y/y]���ʝ�hld���J��g;��V�T��.Yr���{rb\f3�sä���B�)ӕ.�<��d�����pAZ���+cM�UZ*iC�x�I���<v��pkG��=
p�,���p`������#��>��=N��h��*ۑ�1\�E.���4�bR��u�
U�ܬ8���^���Rw�Uⷃ�'J>�w��d�\��I�ռmO�2{�Sò�`^�3w56y�v����SC�T���Ju��M��D�>퓡2+��s]�=ƨ��ZZ9B!T���[�'.
m]:�R�J���'�6�eGl�ְk.���M��f�U��? ���E
���Y���u�z��)�����)�5�y��:۵���_�N��P���xz���}(��b�ԊÈ�6()�/))_;���&��ew;V9R-������l�;1
v��GJ�@缣#�
o�ny;��S�8�8��
�j�Hr�_�����_���WAt��
�����%N^9ʦv�R�{iPQk9J
j{z����ʹ�1ۉ�)�BsQ���ɋ�N1�!��p}�Ůnt�v%]�T�[0�Wa�H�)�� 3~��Hb>�/_Tߡ:i��!RΎE{��Atk%�=�Z���<lW
$���T�|xX�`����ܧ���.M�s1��9tMKҽ#՝��ޏR���%V
��2�X��*�0��Zd`I��o����G^]E��r&r\5ǧ���~����v�)yh���I_t���]my��uX2�>�m.��IDmؽVr��=��}��:�Ց*�*`���)���V�z�L����C��.G�l�$���/S���FGS�N���_b���f����u^8��]��8��}��K�ck�*�oҙ�܇j�:Y���	Y�)K]��jL���+��1MS�Iש�y�y-����$P0�e�F�`��"v��Ҟ���^�C�aѢ��u5`�D���'��W\�l&"�%q���g�[ꉑgF�0����K��ls�&S�xt�e��"�j�A����PM�ª�.g�n�s�=��L�2P3p�jq��|&;�w��P��P�S[���ʪo���겸-�U��}9y�d�
���u�ЯT�ll��;1����P�8�]��}�C=��D "��e����\��.?��&a^+��u��_{�8K^�o��#E`�;��YJq����P����PnskcR8�ka�w��ls\aͮ��e�l��7�q�(\K�U[&u���2:���u\��4������[ԫ���L\b��+�.j����#�9�3�DJ�5I��]yoWj޹Gw��~�Z6I��=52ڨ�#�{��5���E��'����㹲��!����1*gsCK��p����'��-Z���m�������MZ���啮xZ�DN���lY� ��ؽ;���8��IF G/9�١����v��ZR��s��ۘe��OfS�YL�"���|Y�*�r��(�0M�/#�:!w%*#�Ǒ��༾ʲ�T���nÓO���&η�*ܘdT���.[F��bu�%��5��%ͥΒn�<�W�n��1���w�`oSQSsO
�s_ �[������9*XȬB�Q�����<i:v냤Տz�U`4�\C����sWs�Y=x�����u��UQ�%�۩���<�G�ZS}uD�|e_U}�(A]Gc�*7�'�[�}}s���h�`,ͻ-��ϼ��ݖ�z�SXz�b������u��� or�<��Ɖ o���0=dB0�i
�@�t�.�N�Q.mq5�e��t�(c����b��[�u��*�b��WP���<�V�T��\�=��Ĥ3ӲXy�����rlELQӇK��r�ծ5�{ٵ4\3�^��6Fc`�Z~�z`�S�uYlv�������r�l��Mbԯ3�^d��7yzF10,�;*l>"�0,��n!�S�Ba���ʙ��٭�:�É*f�4˳��}j�N[JWv/a��.]� ��4K��R�T�y%7����us���Vy��'9�8]{��m�U�S���G	G�Ee6�蔻z�[�':�Oj��Vta�M^;Hg��!��:���>>��hZY�nG ����`@:aVGcjs���e�i'�=BUZ�r�,�EM;����0���k�^�O8h�`�<��]~�Ԧ��6�Y]��s�[A>X��a��mݫ�z�s�=syZ�b�J�y]�� ����'�Gv�U,����9���5w��6��S	�0�v�^4��{=����D�{�N�uI�Ӗ/T(`K@0�Lj`A��Ҧ��M���`H)��6|�w��r��RXLu�}p �S�M�ܸ�S�X�(>b����\Q��+�W�+8ؔo��}˼m�!�n��l���K��6m��%�=WQ �0P�^����/�K�L��}9�]]J
TҪm���5�$X�.���\��j˖����ު���7Γ���D=�R���Y�x�	}�'~����[�h���)��vm�GX�*na��zx�n�o=��X�ꝍΞ�@)e��T���0L��x`���z7�D�D�=e���U�X~x>~����%��F.g'>���X�2�Y�.�`�_����Z}��}�f�Ov#a�mS�ޚ����S�b�F� ��ok��MAX')��ӳkh1����4b�3"�rk$ո��7�'�f�0:�bჁl��X)����k��f��Kov�G�'O�X�W7����{ME�rur,��+h�ו ���t�`�C�C��xZ��@SaJX�r�v藛}CV�DBm�X��Q�r�ԝ���	����1�A��-�v)b�8�y`���s�t�����&oOi�YL8��X_Γ��gp�0\�mp{Ns{J�W3c��u{��6xS�2��9�lg�ֲ]�U&�Ko+��7�m`5�A[y�ٸ�ەݣ3D~�/�o���� �-���F!�
�9\:!� ��wnn���>����;x��;��u*�*�ZO!)��86u]s(c��F^�A�ྜ�+]/^]�F�#����Q}��qA{���ysE�8��0Ȼ����Vi��7}�P��MԸ��K_,���qs����f}44%�ո�J��zc�]�W�Y������Ch��]A�*2�SOo_
�S��	C�n9��������Ld���\@�*x*x8v��ܭ��.4���ӵ�9��
\���t��*,�v�����tYz�1u\��I�Q ot��	Fɓr*\_�" ����ۃfj3��o/u��cY��"� �=��Io"�ij�k�'ٙg�;�`�w�;3B��\w�����.�;�Eߓ���R%+O��7|�ޤ w�O_n=�ş��G�D6��O�,��	�ֶ�Nw�b�s��qJ����i��Y�ڹy��t�{+;����A��ϒ5���}y�/�r�NLv�������Y9�9G����IF�SQ������	H��	�/{�.�U�z�@���cM�vNCV���,ki�	��C�g_m3�0�A�X��çn먁�*��k8=7�ʚ�"h[������ø)�����x�Ӽv
�5W�V�CFM$.��Fң��m���ڈ{�֠bą�o~����k.$�4s�"Ga�}u�oA���ͼ�Ĭ4h�y4h&\���-_p2��B��m%��&�L��i'+HP6�#T�dH���V,��� ��q���ƍ5�5B�F�T�L.�{�ݷ �L��Ǵ]��n�	��i9��� 0zҍ�����TՊ�J��j��G���A���I'Y�5j�0>�3�5!�P=gK�2>@�#�1�s#��'��ߐ8��A-[)+ւHJ���a���Ρ��a�WL
P�%��:�Fo5,��I�����������m�
;�>{ܜ��C���|ǌxdc1$A38��W{�ۅ�q�+�v�@KK�Q@��K�VoU����93���fJ�ԼNPՕ�-n]�LA�M�k��#L�&V�[�Q�"3�d����-�B��q�սu�>s�)Z`�v5�x�����i9���r�p4�f���o߄EQ�E����-�E"ʅ`��J�J���-�)kJR�D�dVҲ�DUJԱ6�jU��)UJ����R�Kj�Q�J���Pm���E��հPR����,�J�T��X�,��QDm�YYX1X(���kPDQ�� �l�T���AT[m��ږҲ�F��*,J[EQ[E�QK(�m,�Tڂ�cX�+Ѷ�Q�
�,U�(�+UPEQ"���+*�(�E�Z��m%�F�J�6�+Km,E�)Um���ڕ+U�[DZ���J"�,���mKh���5eQ�*0ZՊ"�

,Z!c"*+iKj���DTUj
PE-R�-�Z�KZ�j1�e*QDU�)TAh�U�ʔb���R"��,U�Q��(V�����T+j�(�m����j����6زڵ�U���Z"�Z��J��YTj�E�V(#E_� Q]9܁�H�/j	�&j㳃�|�Eb˗���r�-���l�{���Y3a�S�x������3'�f+�vgu�A�����[�s�����^T�''#��S�a�5�;="��%\��H�N��!D���E@l�v��t��y�jw���;�W�9V�R�#��Zd.��C�'��	���}�37�L��.&�3 Ʋ��9�����u�؎�5��/ܑ�C�̓I�"w����ߤ�7Ð��檴*K��EE�n�����hY;Q���Ufc�كs�,q{�)�жq`��8f�gĆB�'��NaY�m[*n�.
LZ��"�.F-���c#'o�blg)�ٌ�����tB�a��J�>>P��t�.�b�֡�c��w;a�i�ٜ���������˘���0;WP�.۫��=B}�}(���S���}#��h�M�ay�6��+�c������.��6xh�[O�4A�n0���UpMs#������Qșgr�ݘo(<��%�s�\RA�~�P1Z�lh��D�d4�.A����&nj`�s��-�F�q�x,h������a�U�U�Z�V��۞��d'5���91!��r{�����˹*E��&��Y�2��ׯz2n��ݵh>�*�G���7Af������G��*�.���v�{3]�ڢu,�,�¦��h��14	�OO=�}��k]��F��-肃@T���t��o��1�&Lʡ�#�pW��]<[]��0������{��u�]g�$l_�����o�1�
��^��L	=h�%�����kq�s�
ٻ�f�ޙ�^4��J%S�p�Ŏ�l�M��e�K�FI��e�I�;���S��'][�����'�홸J�ѫN��	F�̗^�VMs3�cîU��nh��"�u+
�g^p[�}�^������Gҽ��u=o{�Z��h�T��U�y߬�2�=q7N39ॲR�WN%L:��m�d����`�-��N�x_��R/|���]��Y��7�h��#Yk�J���u��L_WK�)�,9��tX�a1l�����{�t��l���VzΝ���@j�=��8%'�q��R�U��ALH	�RX~M�^gt�,lXU��m�+��x�-³�������PQ+��Y��S�L�*�G�yt]��-�6���!�߸��z�c8441t�P˘�諘1JW嵳V���N���6��{;�fm�h�#gy���.N=5��\vCf�IB:TK;��YJq������MS��*k=����{l<�Z�
���1͚���3X�ٳZ����LX���;�ޅ���v=3t]�^���\�1�
��lPv_s쾾��\�᫯:a��Wcdm�9�wO�MUc4x�� c�\��P���Q��%w�W�fy�.�ɗ{ڢ��m�����aM�WM5n����qSuC�M��P���ʩ���}�C��m��Q�}C�2��ێf��y3�ߞ���b��,�.j�ZY�{W�1��bQH���Os�i誃�'�H���a�D��ѵr�yzjc=���]�����F��Vu=8�v�D�n�%�ьMB4�Nդ3���5'z���L�+lrc���0@�����Fdo���Ζ^_It�ܩͧ�a���[���Vx�&(�Jy���ԁ�KC�V��r���z2���3�9�:$�N�|S��7��y�< �B�ׅY���
��P�Z�v�w���\�T7��� �0�z"S�&����-T`���M�nk��=[4�(z�CsN���ǣG�0`�f�s6`������%wbat[�s ��a�)���M�뎤�Y��TOJ��1�Uo�Mʜ���^�Nz�K�HdD��>�ڼ�3`���s���a��η[�"���M;��D<#�Z
ь��L)���n����r��/�jW��l�m�\3)�(�lT$>[(
k^M�Ȯ�}���VJI�A�˛���V�f&��j�
Z����:���;�1bD�'�B�R/C�R������޹ʙ�tQ��R�ۈ�t��o*Z��:��:u���v�T�Ift3-f���o`T��x>u����E��]��K�
�]Y-��7�)4�NlMy��I'�����g%\=V�'=5�LnB��$�7]"v����0�u+_z���^��g{3��׆���p�V}�>rc+B�ޞ�N��n��p�|�:A���#����]K3$��oN�
ks]�t���z_��
K�:���]{���Щ�K!D� ���B�@|##��j��x�>���¸=m�9�L�W����Mx��W��.|}2��8�,>t�c$6�L� 3�2aH���OuiSwM�QC�u�_hw��nN�vEE�g��\�O�[}9jr5�ī���k.'k�0#%��P5�i0y���kc�\9�Z�j�\��?]C��������Pϗ&�޳�3�V��?��ޝ߮�[߻E��,��+��r���=}�~k���8a�.X��5�#r'�'��0t���^�r݈��Ox��s�g�aZG��EL���<i�4!�2��u����u_,��Ri�(��w~����j��YΑ��4�
*��:Z��p�IWp�P��7B�z&.���h�W{,����,Y^B�����7��v�3����=�7+���J��ޗ�T/���_N�x^FIolN�e�M�=h���мw�6p`�,�����}i����tJc�_q����c���r�E����"5��?o��r���)Ŝs�a��Ң\�'|�ˁ;��o��dw�N�Qp�r���Oj9���^?0c�~uV��e�C�_Z��}�x����k�KoZ
�P�L���ݳA�{ٷ@k�
��vVʡ�X)����k��Hw�Vk�
�i��U��U�O{s��.��Vv\�g����d���Z���Mm��V:����O�z�I�m:V�ܧ
5º0bz}�
\4
������߭�Ѽ�@��|T��#��Wen�<�=�>F�L'U�*L�����˘<"��3ʪؿ&�ʖ���t�4.��7N'��Z��Gt�M�OT�vj!Mz���)7Py�1��g�8��=n��ٹ<s3�f޼U�lz����^j����<e�4�n�¸5�JL��Z��FV֙�S��޸�ۚ�r[1�q�/�!�{W�%�5���iL�gmJ�h��OeW �z�|hPt�\���M��.�"̗"@ݵT�i�<�M��[�pn�p�x��A��E��Q��9�@�,r�Ŭj���� ��s�m;N��I�m#���O��t�O�����Q�o\oݠۍH-�L��wƕ;�--[��}Qi_W<4�9U�s�up����ʾb�?���o�CiX��OrA�l��@��2�A��t���~ɢ{ې#�9ƨ�1�g��1�5��k�k�S/0wu}�'��`8ʣba��\�����:���q�o.�ag��qX�>O7�y)��N|��ɣ�Y��T�tNN�fa��lp�듚�)�ɋ�is�Ƌ�Y[���z�:����PT��4�F��+�8��*٩Ͷ}�=J%	k5��ob��oo�yڵ��q�� �v��_�E�dVEW�֮����J�E_�P��
���W� >��z����f!�U"q��c�զ����~VY�W(�B�X�Y�k�,��s�B��\��T������,��)��l4Ve�C���9����G�FбR�4p�SR�����~���0�DB�X:��_U���*m��y���c�m��'Q�.Td��5���r�y,��-�/�H�aH���]l��HoU�'E�)�.�����דb��x�jV��e��dS�$I�~L%��
����`�����$�'�,:�uǳ��:=솮S ��N1��#tN�]Ù���Ξqci ��k5��c$�O��U���JǎB,eS��9���ړ�/v��TRv�F�ܦtY�0�w���z]_1�Y�51���׃e���'�X�"2-V���S�(&�!c��r���x�(��{�ǝ)z#r��wj�^L�a�>�߉�����2L�uP�h$mL���-rv��	�~r�pW
o�ٍ�@s�BUJEf�ۘ= �_���J���癩/���H��'�j�����!�4�[�&T��>�����H��t��;����������|��T-�;��E l�q�B�YY4ݻ�K�8���X��p	B�阊&v.�a.k%��\p�Yk$l��5��):ȋ����Lw�t��pW5q�����%�����6jCso(�c&bW�Us�j�/�M<��v}�t��X>VZ�5,0#��=�Wl����%MU8��D���ó册b��:dz���^�έj��x�|�j�H���-n.s�+��TR�eJ�>�;q���^ʇ��g�x���<i+U��VȊ��
���J��<��f�S��R�en����&D�1��]Q��G
3\�j�8�+�x�tr7�⵽�5fM��_ �y�0�g�Z�jw~�an�"�U	���k�����E8:��ا��볹W��Ovu�����u������񩺆�R�o�����i���|�{��nr6-�aN���.'��=�g��qv�#��'�5
Q�e�Ӓç�,â��o0���b:7jң7-2�4�whn�E��F��7�n*�L,�4��z�I�N@���1RЋ�b��D<�=�GKg��(�{���d�Z��V����d�l��NʉrVT8�a`���P{u�@��c�e����8�[.�!�ۊ�c&��\��a����p���D����YgΏ����G=�S�bb��P��W�g���/E��Tub�'�v��$���]�d�.��#�;���͹����E,��zú�LޔvTȩy1��6���ړL����ܸA+�1����F�0%�a��L仅����Mv#��NȖ�H��.c���`�uSuu�Y�.���'�0��*��Y���Z��Q|;|
UG�t�Sa�J��I�}׍vZ���
Gz'd�؜OL*��Z<�%X�T���K����4V����E$��rj��m@!Uq�{jP�1ܵ�'�����5T��IW�E9�a^7]�½�W�N�s���Ev�"��X��ڧqT+x�p#Y����>}���V4K�/�C�{hRX�W�4<c2S�am5�]Ez�^���anZ!�k�:A<��C�����*��\Λ}���SF�,6X�^�ww���ķyvN�W�uҟz���A��َ��j]ٳ��)�Ǔ��X����yA�+X�~���:?_:�u^���&���	���g����e���Sri��(K臤D���B�lW���
�b-�26�н��'�eQɑ*��:Q����v�8dA�9�=r�&n���L?\��q�e�V!�;W��-��7-�Q���(��N>�Lhc�ewBcS�w����s���4rq�<�Y\���^	��;T�B�T\(��)ћޥ})�Y}G��.�g_w�Gj���q�V) ׹X�21��5c�c�8��,��1�+W�L��Vy����d��[%P�
��sB�� �3;;�J��S���Q�L)b�8��8���yu~ɧ��֑������D��T����p�l���Ȭ���*S�Eh�59D>A�h:؜YC�5�OE�e�vD1��ᣳs~O��~�y�X���Ǖ�����e_�;a��´��3�]N�Q7�^Q+��U��'�>cj�b�#ҩ�R4b��`�{��-�l`�����Zv{ @��u��S��^F�=YC�M�i	<�}�F39�6��36K�����j�]�)�Jf_�G����)���J<^Jܫn㵘9���M3��c�}2�-�+}�1����e(�Ggnc��9F�X�Y2���>���*�Iuh�
w:/<�+E;�k��-6fT�CU�Dn��0wv2����x:ǎ61W�̍ˡ��A�CѪ�J�
T�7������9���N�Eݾ���
]��B�fՎSv3r/B��J�i*�P���X�	��
�k�Sτ��
g��1˰ޢuX;�]]ӗ7t�N4��P轫�Y���F�*kC]�7t�����Bۛ�Κ_Sae�����7�R�f�{B}Jvrnc^#1(�N\M�w�
��M	x��������"^�|H�,���*�d�p����M���x5��*����*LS}j�ia������P(r�y�@k������):���M0]V���Kn�8�Zg;c��Ű!^�����Zj������dDc91�!���)�y9��U��̵M�wv��yQ�k&K��0*�L�Fc�wƒ6/���~>������d^��r��ĥ���S�9����Zzjq5GlV���S�4�� im�U�ác�]3V:���V�yzb��J7r�q>�)���9��4��ş�3t����{��Ge(W�S+�
�nh��t)nqt��⮬^�-3�Cɕ�P�\��D�����l6��ÐVSݢ�Z`�Q�B�f�qk���YM3�j��T��t�=�
IԺ��o��n{Ip4� ��C];�e��N�z+9MU�,oD��v�:�	��l�z��&�Y�e� ��w�`���On�%H�a�>#x�w�U,��OXW+q]���P��Y�Q��T��z��Q��ټ&S���|��W))`�HeM�;�e��#H�7�6�u��wn#���1�	j�S���/\�/x��$p2#���8��t0!}זJ7N�U��η�h_5
]��7��^L�>�Gq[=OB�r�8if�N04t�/������M�-1�ؠ��~��B�w�{e,�H�v�,�P6�nž�nA�R@h�z�y,d�5_u��8�nlɎ�p��^j�K�]}�kT�2r��a.���`٫:����"�w��S�(\��"�8��!+�e�,�M��["��u0�c����tn�k�-!c��q�ZW��"��}Z9aq��ۥ�Tι�1�=ҙ�8v�:���pJ:x����-�ل(���߷�	YSn��֤ype�-�Bk�5�e@k���G]���
SU,ͭ9 �ڏ��t�)κHB*�cp���6�˷�w�-�jv��KɁ��l�L�\��"�Ã6Lz�����mwf�o f��į�.ýŵ��������+����Y��
���_(�Z�SC��謴<�G����31�ؠ�b�<�|�g��Cb��Zr��̶�~EH�sq\�WnH��Wg�����#cvO 52�+��?v%
�pR�?	N�$-�p��风؛1Z�v����e6�<o��P3�F-�Ɯ��3�=c�^��D���CW��$i� �/��"s��˽��a�>�Z�r�����-ڕ/��[��{6�΅�~����I���Ks!�fû�V������NI���*c=L��vS��GBm�%YX��̧�`Y';�����D��m�wlk7�>^.\G2%0.4�nS�a�AӦ�O�BԏH�Sv��2E�}��o_��w(��v�Q�cȑy�l[�]~ڤ����Ct,���ٸ7`�\3i��Jp�%{P+J����9i�W�t4oS�Ņ��
�	.Ǯ��Ϻz�#1�|zy���=�{���n�D���Z��v��ԫIO+)�hf�W�F��`�@������Y�Otf���qmqΣ�[�C��yɫ˿�*��.|���]}9I�d�٧;)�kEG�_oFMP���ڶ�8h���jĢ��-���d�Yt��W~�t���:}~�:����� ���6�����9=���.�{	�C��q���-G޺}v'�7),
�e��,��qV�,��ݻ��(���ZC��㹑�8r�[zʮ9D�Თ�P{�s���¾܃j|��#N�{/�]��6�5�S�-Ӆ=��c�a�Z�.�>mD_�+b��D���e�����5,J6�+�����,U�¢"0[J��Z�`����[kJXQ���6)F
�k1bZU��X�+b##P����TX"�Ŋ�D�V+[�FZ�DQ")mQTF("�QU��T�(1���meE����F+��B����DZ����X���
���-��Z��[iX*�h�
�"ֲV�+m%A@D���e1
��kV�UYm�������aT"
����E��b�*�`Rب���VTj�5�Db�ch*(�[A"���"��T-�U�
"�m �Z�kVҶ�E��6�QjUTQF�D��R�����AT`�������ť���+�F�ZTF�b"��ZQ�2�(�QTDb#�(���4��R"���5����E��F�(F,�%�����Je��ҕ���mA���Z*�DKh�� �	 �Ird�}���hR�����R..�s�ˉ�t>˚��ls;��wIW&��{/o�`sŰ�1̢���(���U�d݇.�C���7�QN����0��U���̌J�G���b�,�؆�^��Eq�IQt;�\�e�>3Q|��~�%QYw.n��>����d�]��-C�F��+
�҈���+Nr<1E���BE���f`�0qT8�΢��y�y-��}Q�($�%�[ʛ��F�﬎*�O�kD�)���僥;��ԟ��_y6.LE�рq5צsY��N�8e�X���F/k�
u�h+8
�<W���A�����A7T�H���n�FE��o�{���|�e!��h�D���y�a��5�Jğ�m]�L;�Eʖ�.�#W5�[�/��A����.>�����[�h7��>����}C���
�c���=�)��#�oxW]�z�C�x�R�� �)��ó��!*$�w(��9��$�9��jJEdY]]Р���4�]G��w^U�S�x,���8����`�U`J�!�yy\�oNr���!��M�"u:�����ݤ�F*遂�
����j���7����le�����0b����N���NL�4�z�	g�t�/<����sZLWn-���-�N�*p5h��Ex����GR;�����O. Y'��\3���c_ˢ8������z+
�)�h����:��Q-��e6���)nY[9����L�G2:\)
�
����k�+`Ŷ~�v�c�ᔱЭ���o[火9]7O��k��;/wC�����:��U��[��R��#Q�׆b��������^N��W=7ҝ�tn\��C�6Acö"kX�')1F�S2z�lWkt����c��}�����S�HL��'].n&�>�S\�
�®j���7�>�$��r����Z��-�r{�M&�j�s5�(�������]�n0�Բ,����r�R��eV+��f���7T:0��Bx�_X�6�j	"e��w�m���;��������3]S��Ԭ�(�t�ھC�g�g�ɳP�v����&}
�N�ګ�g��g+
�o��$�t�Ӷ��WmT�gV-��Q�����[ί3|�����+hgz�'R��'��,@a}1w��a�p��qo�Ⱥv�ڦ�r!�c�ї({[��qg�� yA�~87�j�S�n#ss\��!K�?m��=w��K��A�� ��۝�&u9ռ�PO�%���޽�V|�'B�5�;��/Y�hncE�("%&��[V���xG;|����b����q u�w���3�dTjd	]]pq7��)�u��jsX��ː,�%n���V�+�-�x���V)�n���,�%�q��:���k��+i�t�r��ڕ��9.�]��R[�77���e��Ѱx�����\����M'�Յ U��Z�u�!��o}9׎�A���=�kӥUkW�@�N���ڤ�-��v޾���a��t�Cm�q�x��x����rb-�me5�K}��h\�Xm�n/�(͛��*��]�8�`��qn�Yy1�C���׉t�ώ׻�@�9�N�3���c�)��N��>��W��{-5[� а�[Im�a�"���Fr�¬o��ȚL���u��]X{���q.���.�V��*���+հ�����e'Y���0l];%����u<k���l��8l�X��k�qa���Q�W�V��P��D�{2��;yY����q�ˑ�4X�j��<|=�7��cl�3�Qv���f;��v/����ŵѼkk�ErB\F�O�{r����h{:V<�=�	FU�\�5pX��]*��+��:u+�[�"�V¨�M��F��ڻ$���^�39I��nW�����c��P�ݶ�v�y�������8���{N��2���t����E�i����m����6��ъ�s�&+9G$���=�P���T޽��7ّo����ұ��T��CZ9�ȋӇkv�p+�s�6�ܥ\)5�N������w#��Óu=j��� �{����p�/�ZS��1,@��j+�cb�<�\�č�U�F[������&v=}Lť5oSy�i�Z���P殶��;g�����)��)�
�q\�)خ�RҿZ9Z����[$�En���3E�wÛI�!�}��u�������bAF"�[��I-j�F�y3�җM�a1�>�I�=ڟ.׳�x�����z�:�hX�8ӝ�-��/U�j'S1��e�����@v�a3,�ӥw/��{z�:�K�ͷAe�5��!�/�W��\.p�}��v�;�:Q�D<�r�%�0�9J�0 �;	;��,4�B�kD�Fؼ�엙u%��|�q4�6�b����!E����MZ�'�ܸMl5j��=����W���L�QF�0r�V?}���߲��Z��܉�v9��I�]O��5k��ܮ�Uk,��T9Ņ<bu
��}P�d`*�Yzg�<m��fųK��ǩF�S�{:��/o������J:�w���<U�TVb{�kT ���0��u/�}0q>:nf;�5߀�3�V&+�0j%bz/7S���S�hp��#�7�1+]�4pQ�c]�X}/r��dao��y�������6iXgYT߫��y�yl��Q�y�N�n�ө����N�ƌ����[�3le%��U��'��.�ǻ��:]�<$8$�=��9���[Hc��C2�LM^HN�x��.:)��&\�v�K�k�VtpƆ_�w#��{�(���
�r���Q�$��|�s�ŝ�/�Y6q? x��ݾ[�����d�-t�m���T��w����\��y2���7	������ ���c���tf՞HẐ�u-�@?������^��C�tԨ��{Y^u��9w�s�ퟧ�{���9G�N�q?bb��e��-2�Bb��j����f�rr7��A"l#�j�n�/��t��f��N�:�C�n�}p3��ؑ�b��İ�K��5�������؜�]<���\�ܞ߼�Z��~��Gq��۹O!�k`��qem�g�rU�xYȫC\[D��bվx�N����Ǿ{�:���g���k�(��E�겭e�����u^�b����e�;�9}���1}g%c��\�}f9��pb_)1�T�zON*��N�p����'�U�K�����kWs�p���V�q��1�dEGb>�.�>��jF�[��P6�k7${�I^R�t���f%7�늭x�U�>%#CF��ˠ��/�l�<��軮q�w�֘���q,�
qS�:�f+M�/5f뢳U5�6ԃzZ�"�b��Ԡ�N����q�[as����*����
�ֶ��y����*��F���JsF58�Ne��cGYd���veV��
F01�����^����F8�y�n�J�%*�ʉLK(�(����p�ovfzhe��'1R����=g��@g�����$��wI�'vp�� ]�L_��)8*�vTPָwF-��f�ZQ=266�V��U�7�e��G���`n��}�b�X[��U�K̈p�e������˛�ǏN����_��dq�{�^i�����/V��nO��ڮ�jnE�Be�}MC���vm��kh�Z�&�
Nf��&x�oRq��Ѕ�-$��qO�5ӻT�ꫜ�o��W�&�Ҹ՛�V���p��q�]P/�JG�S�r�>��[��]ZH�����eWgEs9�R9�[�S��<�Jj�#��y�7M��.�\�4Ę�1�Q���Uo�k���:W�R��<j�Vk��8�p8ͧs;b��b�<B��_Fv>���hK��{�T��UZՓ�Q��j�v�񸧢�.�M[mekɴ�;s��!(��߭�����.�9+�]c�@�U�.�8��q7q���}`7��ķ^�Z���B�P�(�X��yZw�]P/V��tς�:6����JbZl ��8���5y��ђGgW�|q;��s��r���d�q���7�Qi�7ݏ%��V��Ɏ]��Y��0�������q���۬fzt4R
��[�ҩ�(���ptccq�R�8ȳ7��Vv�s�vi���mi�꽸�o�R��|}1Vq�.E `2{�u5xǱ{*;��fq�ƌFF�1��|S~u7P�s�Q9���Wz�˼R�j��Ն�h!6(3"�ӬUk�4qe���)���P��].i�G5n�c� ���ew�c���B�(-B�ھ��U]���Y�ru�/��a-��s5i�=Ƈ3��y�ѝs9�/�q�o/"1�}���b�Gn��r�b�]t�&�L4�n���sНp��^V�,3F�͊�mYj��x�0,:�}��0�m�K7�M���X*�o��S܌Z��]��1μ�F>ܝY��y�]���{"o285�P�H�{���CkCogr����(b�E�9֗H\��N�Q2�m�
U�xz;U���s��V���n������B�_S1iMZo����w]8���c͏Ϛ�	��w�Κ���s8xfهj�p1��79�)���]�Պ뒒�v�ۯm�r�ʕuL5�oa��U��0)�o�#(��ٸo!�}QNd_|�eh�vޢZ=�V�I�`V���� �t�2p��֊G/��K��+�l��������])�;h:ٴ2��D/]o��[�qyy#0��8n���6펴�v�q�}9͖$��Vԝ���g��"�j�ف��fu����F-w~)�-�y=׋ʘn���٫�ֈ���ZEm�f4��wF]F���ϵw�����{�'#2�!�*���\�95�N�;Ô�:�o���h�&����۶4��Z���:�8�����XsѨef!^�!���������ӈm��䤊v��1�~Nr��w�w�
e3��TEdb0q3��M茕)B�mn޶l����U�q)Ey&,�YW��8�ƀ�>�Ń��z�"rEX�>�$�nt���ܻ)v�ҡ��p"bk�^Qh��k����ꗁ��qT�m8ՈM�S��p1u�Mέ�
���Y:��1��:��w���5}z
�fС9iV�t�dn�r��.�v�:��B��iur�YcS�z�M� ��o{X�pƜ���@�I����1udԹ�/��A/sǱ��0PQ.�.�[fP|Va�ǆ��G>BՙP�w"�	^p��6!�4�v�T�9w�;>�)�j������Ɨ~��M)�j���1Y��g"sg.��w��͑��vj��Rf"�E���
m�W}�s�Rj�{�4o"�;��c�w�7s��zE�}�/$(cT/E���p)�=2ʼ�-�y�i4ۛ�>Ŷ��6�r��d��P��_r"��d��\��o7���U�ӛ�ltR�~�~��a5��v!ӊ廜��H�+�v�=���;���5�];J����o�D0����5:�!��s8��Sպ��V�ۻ�-�إ�O���^��[�o�A��f!��X�gf�������kk���D�p��"�pc�)>��EN�k%�ͤ����9zh8�uɻ��Êy�=��x���H�⚜hGb���픚RT���;���w �M��Sx/�Υ�J>o�^!��*���q��@{nI�$�u���:�tUy���e$ٮ��lquŚ��"�.om@գt��t�[C�V0k�0�����"�`�[#��7yn��y���QwY�U#������7yDjT`X"*��V���\�/P���*�_g)yf�� ����;�Ƙ��nN�7���C>tx�zS�\��)\cr|�n�����sV+�A�'�kwe�{Z����ͩ��׊?��'�1�{�*�vO�ͣG�`�07���wF�MW�I�]��1��@�/���j��˺?/U19��wGL��^���ɜC���8-NmuŜ�`u;�d�N	2b���F�%���*e�@��w�^�JP���r¬�m��}�z��Pû�/-V�P���䙎�%�yҺU�K�qj��v��'Ode��Ј�Oo��-L��ٰ9�&2Ks]\Y]�t'3+����甆j<�!��R�97�f�1���TAʸ��հ[ʴ[��i��i�1�g�X�Z~�����Y�
��i��ޛ�״��p� ���Mq_ù.j���]�AW�'l���	FF������Xz�[W�\�R���G����h��q�I����^��U-��T��*Z��7���r�\ʎ���}����x83֎��"'QF�:h��w4�M �́�yq�q��F}�˺�U6�3�s��*����5��Z��-��[0��6 �pa�9a\vehh��t����Qv��=x`Mx���u
�MR�v�8�?X��*+���t�~���)��
���y:�YE�v�D�m�0�b�n�O�dN���%ui����W`��	���^>��f���V/�t�s"V ��m
��ܙU�2�S�<D� ��SСiU���ym'nn���ƛ$>55I]u��x${��"�p1^�
��t-��H��W�E!t�#�DJZu���7��u�Z[������pG:��£�s;�\̴��uw�d!^V�u�sXu��]3�X)�[�qt�9=0�|3{���{kƣbF*C\[B��uf��W��G*u��l�Ne����(ogX�'�[4��He� "��M�f�WjY�S�a�1S�����5���j�ѽ��J���pFI)�8�W�7F�.�b��$�P\��E��fZJ��H�y7�����\F��v1�܄o< ��k"`*b��F�tĮ���`�Gt���Jܕō 81
!4�F��aN�N�uë��X�v=�^`�����O;.yf�>
�D�eඩn�4�X*��*��s1H�{h�e��,L��j��YAH��ch�F��y�$�#�>�zI��(�C,�"�wv>hb��8�7�mC-ư�LC(2� ��T��r�$�+F�H���TgBU�]�����,ڼ'��pil��ϑ����\�Rx��?/�	�r�Ib������+�33~{��5���}�LY�ث(�բ��h��2("(�X���#�[�m�Z
�"�6�آʶ��Tb%e�(�U��ZQU�J�KeX*���b�b��Uj	iZ�Q�U(��D���A#*�m
���c+EF)U��j�mE��YF�)��*�R�iUej�PTQQ�T`��"5+QUH�1UQUb�E����m[h֨���XF �kX"�����Z��EJ֫U���(�+cl(Ȉ*ȣ ���,Y�,J+��E��UJؑE�ň��5*�#[#V���5
#Z�QjUEX�1�E�lAEdH�#Q�[DTb* ��e���E�ŋUQ��ZZ"��FP�E"�@R��Q�bب�U��ZYDU@Eb�b��E����1TPF��PT��[A�R�֋^�����蝕s���犟gu���3�y�5�����``�Ne����f\�[�[��q�h܄%JQ�����ukd^~���_qF���5��8f%�G
qS�:���kz1*'kqG^�lh�v*#͸�*
Lbj��H�} s��3�����^�E�+U�>��/ُ/l�jq���>ܤV5}r�M�ur���ւ�r�]���F+�����3Zy���,p�(��6@ǹ��I�8vZ}�uvh��g5�@�_a���1T`wӘ(E��u�쓤�ns�5��Oo��]�P�'s;��y�C����V;`7oz�(�����W]�x}�a�wn�6�ͫ���R� �,ה�<��򮷠�����t���kRF8R{���M���;�������j��,��vT�z$]!7�A���f��|��"5>:r�@����t���H��f��(1�u������J1N��ͮ[���a&h���
�c��sʸ+/%e��%�.���2�q_�[������5k�.��܁�t��L��lG���&��MmO��+�^�=�էV5�^���#��D�RvT���H~Q5�
�_w��5e��2�E�5Cy]nmjR�T�n�|��S�Ч��il��B�R�`��\Jzlj�K�]�glk�i;C���ӝ��<�pxr��mN���ӐdX�s$o\n���k�e-a=���u�����5Ɉ����s����eOtk�����sS������ĳ&:��=	5]ϫf-���W���v��d�J�0*;����꽎n���N��1�X�4򅊂D������o�p����*���L�d`�X+��m�s�6$�v+_�dT�iս��fӉua[8���b�^����#��wQ�:�I<��=S�֜��iUw�3�ʇ�	�Qh�}45���eEbf�,�f�nx�y¯�YrG>��EB�{7��eyk��o����m����,�3+7�y�E=���x^a���mB��s{%��~�ׂ���b^�w)��O���Ab��)gv��Ǵ7:�y|N�@7{l�ڶGW6��{!g�!�l8���鬝�f-����5�哜�A���=�a^�f������TQM�T�"��9�Ї���+J�z\-�����4��+1���%e2�s!q�E�-��������x�-~?FW3�[����	���g7Yٞ�G9�j��k�k/�z��L���\�(�/Y����>�];N��<������Efp�yn�zr����Mn��PR�m/p��Ӵ���e���Ѱ�cӺ[z�	�:��If�ľ&v�
���Jr�U�[ʁx�bޒ�*�4\'k�Cuj���P�֥ۮUӊ8-��Ʃ���gL���,#&q�ћ���Ih3����:���1}lri6�q�ӝmܳʝGr���9�bR�]�J�	uQ:�������Mv�u��3��N�څ"o*U�c{vf��d��1U��	uZ��u˸e��`�=�.��5õ;g_f�/�b���x�(�Ӑ������}�*{Kvy�c���u>X��,9�<*�VE&-m�\��b]���M�T�H���3��g�;:���%m�<��J]m���Z˔qۀ����#��t�xihL�jh���`���u�|��M���6B�{�i���|��e�\K���
)bp�-�i�Jc���ə�$��u7.����
�v�ի}�e*W&$o(�5�rp���/#C챱0BnX~Ï���	
7ٝug��	s�j]�����;\7)0^z]ĳ��F�����|q9��������Ʌ����Whq�ym�y�$Ŕ�(�9O8P��]��
�g������{���Vk0�Ciå��Ne�mg�8(�5�-w5��#��.�"�o�4�����P�י����G�>Ml��Vtwh/^�T7X�j��+�X{Fe@�f��q��0;8�>�=/+�U�'�j6��.���}m��У6G��f���b��z�)��q�N.�'V��+Vg1�Q��ݺ�������7F�6���Q��j����Yy������O�C�SO��w~h����p�6�r���;=Tvy�6rU��V2[��ئ�;Nw�zؿR�c�~w������x����#T��9ҹq����PY����[�-[�$�8.>��:1p�j09ܓ��3���;-��,�_@tXv뺅5י��rծZc�sL�=(͵܆���KcD��b�Q̦�W�]���}S��y�ӪL�UT:@���]r��s�Cz��d��|� �T^�m�1|� �:����Q�{��o!��oٽ�f9����L�5��q�4�y���>	{�Ͻ�O�Z���#Ym�{���w���@b���eE�T���y�<)qf�Dl���q]�ₛ�~��R�%7���Y�.o��KJ�Â$>�u�SQ��(C�oU/LD�&�΀軉w�p��]ˁ������巯��O2�l�="�Vg+������۞*b����]��Y�W�7ceE�VH���g��g�qe�c�Ţ�����ܜȐ_��-4S�z�UWlݚJ�r�����f_�v��=��{�E*��ɧČ\�⽶,C��$���}�*��w n�}�+I�bys�x�^�y�܃�Gj���l�7�n^
/6G��e��E���wJQ�7k�q������X
�/qX�YUVh,�����&r��?�-� I叹3��:��o�%1V��q�j�yg�Cqr	q��m�.�~�(WȬ�b�Z"壇���7������F���]���U�T�⽃heȲ�*������Ր3����PjU��4c�jw-dF��g��3λ6���ۗ�"���\��6���̫��O��8����#)=��l�nn��ݿB=�[��(al6A�c�ޡ�ý��q�bkY
_8������Z�8o�zwl7x���K]�OMy�<�t�خ�P���Q|��#��sѹu��Y�g��ͅ�ol����hj�<x�J���F��TҸ5��l�m%;}�r3F���|�������r1��u�(Ia�>��N��:ԭ������髾3�s�Ә��XJM��]�)k��׳����)C�r�ImC��`u-sԔ������S�:'S�zࣆ"�qn�Yy1�J�_U��X[s�N'�r�9dX$7�*����?6���O7����S�s�a�^ju՛��I�Z���tэUQY��F&c#Z�����m	Ï���sIO�,�8GǺ�l�Ψ-g���k_[����
=|}�@�-%�H%2u��A�;�i9w� 8�2,|7��gI�}ӫ9���܋���m�-��::L�+��d�m�|����h��e\9q��v���u�6l�޶;�+�	��,2�'X�V�1GeK�B˥|��C�k��|�x���fS��)�,�>��	���w W��&3��]jT����gjr�i��N+��|{ì�hξ����&���8�㈍7<�y��Ά���H�5��J�1��if���V��s$̩©^]b�L��d򄓁�ׁ��֣�[�|Y�Ŷ�͇��n���XTq�=۽M��2���0)3\���җN�z�˦F�Pt��ݝ+�����țQ�x��۹|O������|�we�uo���;u`�qm4�'���m����
_S�=:��W����ܸ�����*�ou6� ��B��W��F��k���d8�]���v�����k�AV��I��;�c�ζ��&�FV\F�X�C3��]D^}̒���^M���e�� �F���Iz��n}o�ɱ�5���Y�w.k~�iQ����j$ˈ��>��L�֭�O����죡"����.ԏ�c��Ըs��,ܠ�s\��˧ãm�.�(u��HNR�"-�Hv�O�]�erQ[��ՙ��u��|�wOt4�wۙ�3wE�ԃBbk�V����}�uB��s���[�]Zg5;��ܲ���3`
�5�v.���8o����
��(�✙o"��9A=3��lv�FAu��n�ڪD�݀����dR�u�Ň<bu
��b��1�e%{�Vk͙�<�j7��gy�aW��pSܻ�g�1)��ck1@�^��.D�J&�.r�:	ۭ�޷��kF��yE$ŘN��3��3��w]Tf$�p�_
�^�Iq�8�-lc�ZT:��+u.��]Ub��p�a���k.�&#藸Fu�Ƴ*�'9Q��Q��,�5��u-��J� 䵥f��vy,�#^��-'^�M��^eVcՅ��U�������3�/���
�����߹����ey�8�J�15x`Rcd�DEʙ��x�;u䶘�'������y�3�VZ��y��
�f�>���<Oլ�Ҡ�c�:���ۙ��*�>�Zrb�wn���1K����"WF�c�iٛx԰�����X#���^1�~C���L�v���ܧ:���e���r:'{s���6��+)(���TC��L6Y���î�܏7�=�e�a�P�zh-�QM��b��uP��JIo
M��>D�V��qz:�۸c�](�%wH�phҹ[�G1Iq]Wԍ�5�M�iV|~gGq�6��Ȋx�tL�ő��[zҗU���pJO���(K|8x�M�����a'һ�7����WM�̪�ܫ�`�O��ꈽF�.�����j�����Enwb�p�'	e�nS�=U�w�1\�0�p}Ô��G�Z�ў�)��֚r���1��\"��E>i�����؇oܠ�+&T�5U��B{�cH�U�et��oz9����R���`�߸˞ȉ�Dp��^�\Y�/�Û�ہ���y�-�{һm\�s��
9�&�s�O�_��� ������,�|T$�&-�Q珽j7�Z��\غ��;~35��y����,:N{S����L���J�̰�E�������2K4E�]�ܢ����&] N����ݜ�G6d=��,ďS�#9�&�?.M�l�1��tS�R@)��6��㪰���L%�3�j`�aWޙ;dD�لuY��d�^X{ۚ�#��OF���nqx��+��}h�;Y�gV]j�	�F����#��-aS�Y�d�B�Ԃ��#�܄O*���0�����
6�M;�ݩ}�+5�;�z���E��^���yJ�~��ފ�{�m��a���/t��2Ȫ��[:�+����"�oqH�>گүU6�ϋ/�uٷ��6��;�[toQ�n�N��vwT
�&�EE�����p���x�k�޳�yzzpˋ�d�MV���Ξ���`8u|�)������b.nR>R���[hfv��1���8�%�D��*�Ӵ�/�&��!G'��Ҿ�]t���N��O�wFsCVD<v�h�t7y�����tkt��z�<��+�&S�};�c���_<���&c��77��	r�o�r�;hz(<�\Of4U<{Hn	ae�w�JUgFX�"�a�X��>�k(s�h�;�0@ˮY�w8r�o9�#�	�T��b󵌢a�G��F�V��$��M�ɻ�����8�v/ ޼zM8gi���Ǘ�a��!U�{��y\�Z�`4 �]b(�e>�,q��	ʸQ���
�l�ެ�[Gm��a\�6wg7���.<���<�!�L�M��*�"���͛�HA�ѩl�q`6Q͕T�������{o��D������J�l_c�!��"���*��KħXX��;j;v�buw)�KrJ-4�+�b�٬Ӄ�Y��w(ee�������D䣣�U��"%�3U^K��JYW�XE�Qm6�&�"+;*v,է�����39 �:����/�cv�Wu�x�Qf��|t p^4��2�=@�7�f�8S0�.���P�h�{���{ō㜵XN������s�#ɵ��2n���\B�I�ߺ�=p��u��.M�弹κ���ޫ�dѶ���co��cpm�_d�M�#�<�0]���=��#O����X`�y���.aB�A-�J�T��-����
�y��;�02XO��M�I�Lꕹnff}�7c�[���R�B����ɇ���k-��3��y�[Y���e�]чR!5C��5�eD
�FV�x�hP��[:=�U�vN�FCJ��
XB��0�M�ľ�']=���.^}"czR�*<���P��*^,�i��%�z�9�<6��#fV}ӽ�����Tm"��_�nuf{���JI_Cr//A�y�U�#����X�k,�z����	g�FX'��rd!o-^1ɎP3E<IKIM�^9j��j�)�Y0�r�Ap�n��l�VZ�a��X������)�U�h�²]I��LH_�V�g��HO�`�T,E��s2u2�f���$P��H�{���ux����8�NҼ�(�q�Ԟb�S;�Ӵ�#�Sg�r����p���\����
�Vi�%7W��&U33};�[
gI��E+��;U�_r��� 1dC�>5z��(�OG�=u���`"VB��kz��3)�����Ay��r�\�\�M��o�\�r�=�I�o��SW��Z�0V��յ���3j����V���Ug-Qk�Qa)���$0T-���2��q[��CN���5�Y�Y��7[�陬{����N�ںX/U�;zmk��=9f��#P�������![!���l��,\�1	D(�n 2��^8&�Žɭ�R6F6�� #!+a@݄���B��e�F7wXp�n:�1�&��M %yg��F��C���qS��lE%���7����`�V�e��
�9�~�P

�`��1F*6�TTE`�aEQU���DQm�"���lE�#����Z"�UQb(��� �1ƴDX� ��X�Q�,�e�	Z��AT`�H�*�*EXT�+"
,`�����X�mUH��
����E��*�*��UDDV1D�TUX�EDV*2��V
�b,`��F*�QEF*��b"���*(�b
������ ��UX� ����b""$Q�����*"*���c�25
���*�AE����U`�VұTc-j"����m,���X�EAUc��DH�(��*Ŋ�����UQE�U�*����Tb1X��TPH��UTDdUQ�*�b��E(�Ŷ�1��b���Q� ���Q���*V�ET_�$�I ��<	vq���=��n��;k��S�r�s�^��ko�Y���T����(���~Dٝg�Ҷ�.\}�5{��a߶Q^o�)�d��eweM�]d�-f-w��'���㸌jbk�(K�]D�v�7��%_���t5i�L�r�{�Sx.����@t��Ԯ���=�睂c�.3g'3�T<Z��Uw�U�(�[�������8�)�N�0y��Ԩ�e6.�F#r�эx�Gފ������x���Y��k��UZK���	��"E۾8���N�^�z}G_��xv޴Bk/[8_Op�'���&C��0���hk�����؛�hVR���N)��xz���
�*N)'�a�ekシ����4_m���+<����W�#��l1X�.3
8n��*u��I��6�^
�N֕>]w���u`\eL�#���������vr�>�Ւ�U7��f-�OҧcN0�n��p_CW�W���Q��SW�Rc�Sǲ�G
OO�̜��K=m�=ю��OP�(�1v���D�W���{����^��K�Rg�<Up�4��-��g3B�7���W�7[9��R��#�G��������v�	��GNJ����+,g|�(�]�<�]����x2��(�{�* X%�j�S`����}^~�uS���r�/����)C�������c3�/5�H��	��Z��O�8t����h��zc��:�+��hd�RW���.sm�e�SZ��I�iSA�!ӊ�z�T��6-����H�Fۊ��f�z�k�x�coܒww}9�ݱ&����s9�����-�7Ř���>��Ů���S��Eɳ�U1eqJw�T�r��xs�;h�n*�:��9��B��)�ۓ��9��vJn�����uXqO8���لeJ�S�+��QpHw�-�~F�4{�-�r���(̀9k��ڰSr`$ڰ��C8�w�W����W���*����wL��qi�y.�Y�p��ҙ�b�9��z�����wGw�L�u�F�犃	1������u�rQ�F�f\��;��z��%����'����'`ܯbܖ+�RW�q5���3�8,L�����=�؝����ԔZv���<x�zt��W���ii�t��F��{����:�B�6�c�E�L��Y�2^�X�!���g[���nzbE�w�@���B#�b=[7�bV`�Á��t�5	�+�7�ڊ��vⳑ�8��c��P�Ƨ	c�׸(wn���*��}M���SN�W�+J�01Y�k/0Ѳ��8]Q
���4����1��)[��h��i�Q�+ʣ���/t�ۜ>�u��r���`� ��s&����zh�[����~l��s(���Q��LM^��P���̮�j��N+������}���;�w�O7[Ly;�_�߯
Uo=�ϩ
H���i�;�:�EE��l�$��Ro,��ۮ[��V�[Y���^��lQ���}iM��8�>UU�uCk~؜��y�s���+�3�^�k���Z���8HesB�����y$�k4�0�E�Zw���;�����w,�5;�@�(�4� �T^�b�*;ٵ���ıyz餷0��~/�9i�޼��s�����vъ�n��un�YG�-K4&�Gi-f�Ǌ�.w�*��	]/B$[W+�SK�'����|h��M�l7�bw��#�0�9kͩ�8����F��r�ol��qUGQxѭǐ���x�-�µE�k
��{7/��R�eN��{2�F�N�Pq�5EƂ�Uὧӥ�o2V糮�Uø��{�}v����sqm��=�1\�h��{k^vM&��N�ܻ�yR�P���,���(u���5��Nu��dc'>�F@�y:����%��L3VO����DK�e��鮯N -<�����1`�F���ph�Q���:�n��8y2=�6�$p;��pq������=t{0��Ȱ�y�<Jk�NH-7
����/�(��a��w+A}�1_��(9J�cz�����W��)야U�q�a�P�m7��+�^�<+^l�1/tɨ6mU��e7:�I�j�V_k�sڋo!�g���:��n�hXj�*��j�N�S���穇��l��5\��N{ZG�)=�v�<N�-��ݾ�����՚A����[8��rz�o��\��HTmNU�*������voM���xg�a7�tW���у>c3�n�o��d�aqʈf�{���恃%C�zc�]j��`H�z�r�ow.E�G��KJ-�=�wu/M>��NNX���[�y�a��ˈc��;�(u�*"Қ�����+���F$[�u�I�t-�ZwK�zպOw!�@�WN+�����%���5��Ga�绢���A8�C2����;|��8.1��)o&�qPg��iA�WD�D�y��k}���H���L����^+����l��9a�w�G�Js�@��>�Ƽb���U��]��c�f�c����� ^LZt��s9�c����x���*y�L�f9w=���wd;xWMҫ^���Ƕ�ރyL')FqMD�#��m::V���(;�ai�f�+T��a~�.1	���<b4K���E��]������"~����,���:�I{Q�lV�1G�.�����EĿC\Gy�I��]bG�k�+��v>\#Sf{W����>˅T�E։�˄'���Ȑ���f�w��I[V������e��L'���`�ꖂθ��s(ν����"�U�s��l������2s��Ȣ
F��SD�=]�v��3I�M&��%5�����x����-�Ɨ^�AI�V��{r�ﵝ>����^��эN)'�a�ekゝ^5[,�Jk!�C�ʧ�%<03l�cy~�+%�n�Ta-�p��y�[��K�	��A(o�)�;�)�`3�L���r&���5U����!�n$���k�r�)�å�kz���m�^�>X�^HOb�EAz��u�*��<����6��w��;E�sv�7oܗzol>&kp�R�k�a�cF���E"����+;ԸժBռ0�j�'����Jw. }G`�k��U����}ս�d��ئ�3�Nj-�y�O<��q����$��]8���F��=�/���ES�~5��h������Zi;��`��M�NΫ�2Eʶm�q9ZokP���p}/��h�=8���6�������+j�u��ޚ�o���Ƭ@��Wa�����M�Q�����1�/�n����	\ב%��S�4*O�:�T�1.Tێ�Ҡ�݉��za�F�΍�&�;čv9��.>C;��g�n��w���;'��t�}�t�tkq��|'�*�.�`[h�I�H��`�F�3���C[X��\z���ò���YG���b�Iuc�/����� ;�`�c�]��:��o��5`EN�3���K|o�����r���j����1pu(�r:5UVb.3v��`�Ӂ���̦���<^ߧ�;I�sO"^ľ�;g�D�nj�n^s{{X{���4s�靨��Q�=���La�'YF!3���xi2���]�έqa+$rp#��Y��՘�-�=�C��$��׻Rx����Gm�:H��dvb;��%���`V{�b�X�e��e9���^�l
�v,;���x���Ň	p��k(�;ʣ���/t�^d�#�I�����!�k�)ʮM˼��[� rV $[�n[��<��kz��৸;�V�����n�ؾM
�.�Q	k�K�Sz�n�����zA2��6D�Qԥ�"h������)�W80�G��:+��@��wp��#�#�N�R���ef�qwX�(�9qʼ�
w�jH���i�Я5Y;u���#k<�P߽۪�5ũ�'�0�m��(�/3K�D�"L��5ޅ7��s���o5�Z-��#Cj=��_f��3c���MG��{\��<�t[��:88�Q5װ�&\s�b;��n�w��,t��i��>~�W,��_�q��W6%M�����nb�6��v[�����W���)�G+�.���.U����r���!���OgЖ���S��c�ζ�
�T�*��Vkj=z�q+ž��>��j4f��&�T���w����Fa0���LN�1U��^���Z��qMٜ�P}7j�XL,M�wnY\���|��K�~UB�f�1��A᫼8���P��XZ�1i=[�p���cQ���� �`�>q�ĭ�qҙm<�
����a�g�z��0[zbu��޴�����\�,��i8�k
���1)�A��k��
8��V;�����H���tR�Xv�-<\j��x����ɕk�=ᇋKع��s+zTt����skQ۬ɧ��)�u%����@�s#�"^���f�Y3'4��0zC�d,��wWj�վ��o�(3��Z-��:ȁ���h�4=�*���ⵑ�J^��#��湋l�*�26(��m�83[��2a"I�F�h�e�������7w��m�t�m,6sB{M�RZ���rl���^1ʚ�`���n����i��*�p�9���(�=�a��v2�}��[���{ř��ǟ���̤p,>�p��if!�l�l�܆s(�͑�ڤZ�9�n�mm�gK'��ف�f��6���|c�=��yy���������j�\
��V{r�l�9�X#�9��k�Z[���;uyڪ�m�ti�p�؆��]�_�f��L���ׯ�U�:�ף8PՔ1�I��t�>�R���F.J�7��gC�^Q���[t�Wt��߷HX�Ԅ�yz����T�z�n�y$�㏖��x��*jr��z:�S�Kf��	ᆕ��[�]ĳJ�i�\���v�n�.�ӽ~�hI���\㎕�˭��ǽ����q*ѪI
��:5�b�p��Z���k�zF��T^eotL�ͪ[���s�	�{R��۪��}��ZgS1˹�x�c}����UR��E��=e��'�������
����Jd�z@�X9��G6�k#s�e6V<h����>�!:�c�E�j��;Cy�����x�;-S˩k�ݱ��+�[��	�d�r�#�=ҹ!wL��wQ����g��m��˺�/��V�aT��SS��EC�b20�u�Ž���܅=/\�S��ُvwj7�\���b�#�L�c�<����uR{­m`����9E��l�L[�ua��e\N�U�r���N�Y$�2Q��v9_`��L�r�����0���hk�]�VoLX�;xC(�e2��\���9�FD�{
�G��d�mf�=CU%i�����C�i?N��}���cyq�Q���u£�ۿ5���m����'v�Ls��P�ٻ�~���`q��e�V}X[��%ej-�*'^dJ��%�w�*���6ɩ�p�z���j�1�V�nN��k���;RG#`�}��(j�\��,�ݲ�}�����r�_5�!C�G@�]M��r��[$^\��ԅ�\�B{�t*廈���%;w���=�G�=�߂H@��H@��	!I�r��$@�$����$�(B���$ I?���$��B���IO�H@�r��$�$�	'�	!I��IO�H@�8B��@�$����$��$�	'�$�	'�����)���5���,�0(���1%l���@Ԋ�TUER����$U
R!�
-�6�T(SJ��emmKc*"�6��[h�ڔk�*��j��)R�LڦfR5�X�v��ݻ����e�l�6��,)��Ɖl��U����Y���b����孶m"ke��:E6�cme���WRe���V�fm�a��5�UjdciT����֔�ٶ4��m�[�[km�����Bƭ-*jmZ���q���a��l�m�Z[m��kZֆj�nmN#e��#Z��  ��=](i�6�����P�Ju\�
�(fs��
�v[���Ue5u��Z͓�vګj&E;��kYm-+`P�T�mnk��ee4)Fl<  ۞5��Q�w) ڲ��Z,��eUSF�ecVճk-�s�Uf)-mv��頳�pt-�m�v��f��S7Zٵi�)Ʀ�md��bf���  n�x$��ZXm-�@�ڭ\��$]X��à)r�n�u�J ڤ���iT�m;j%�*�j[]�^hP�@��v��(hhP�B��ݬ�А�B�
(=�L�&��i�l hV�  ;��B@(P�AB����
(P�BB��aB�	B��{Ǉ�!@P�B�=�{h *�c�:
u����T�fgN��J�&�AJSE��,
6p��d�V͕a���k'� �������R� �\8:�*-� .����V�X�DuZ�WCP ��s����F��n	����q��Z6�7n�4m�  ]o`j�����.T�]ˎ( F�Zj������  �N[��(�p ���C@�ݻ�l[m��٭M��lSm[�  ��Ղ�Gup�N�nQT5VN�	R���U:iQ*검	9�J�����Q�R���wv�p(Ӗ��5�����V(���YZ�   ���Ԥ��P�Ғw8hSKY���U-iJTܺ�Z5snZ�c.�PvĴ�ەE.)�m��ГL�jʶ�h�n��6͛Vͭ��F���   ]^{�@j�����SKp�u�SM
��;�h�ikb�������d�
7.�BJց��Mf�h���4Z�Ci�Y�4!���T�l��
����    �z��m�ɼMN� V��qr�C&�e�M��S�� W]ź��Mmm6���h�lX+j�J5[a�չTւ�J�*��@� 5= ʒ� 2 S�0����  O�x�UH���aS�A)TC�����a4��M0	4�&eR��0F#'�~߻���??�����Ϡ�΍������z��k �H	�z�#F^T�w��7���ٙ$ I3Z���@�$���� �$��	!I���$�@$�}���g��hܟ�lF�=DMf̚���u��X0���qV}#ʛ �h�t�Ѧ�:
�"��eE���V�{�7W�Cr�5��.�}J�V��p+nk��l�5�8��f������L�x�T��4]Э����*(�5�G~�I��~�,��R��4���͇�aV�hkԲ�D�0�%m���.�"�yZI�;U��y��MT�`ߔ� UhawXs[��5qi��qh�:5b�`Վ��T�6�I�E!�V�:&-s7J��b�)�5�B6�`+���p�(�Yr���fԨZ�p�p*����2���k�I�2�a�5d��(�A`M%)��2Rגhy@m\yI+��@�f\2�\�����f:()#��0�+A^G�Ĵ��|�H�ݛ�����u1ʀ �p�"���62�jew5��3[G��+m��ͣ0�
�c@ұ�-�f�E\�դ�:���R�-��R+CѤ���wP�ܹG@�Ѳ��²P Uͭ�E�Xu ���n��GM!S0e�Ǵ�+Cde<��VqC$��Q���D�5�\�4s(��Lge�YN�u{���+1چ��t��B�6�n�4�A=��@h��GX�jı�Mɓ2ƀ�&��EXE� هVG
Wu�^�F�X�V��i%��]^(�[A`�t�v*쒠��0��>�ʙ�V��8*FS���.jdX�1+\n�n^J�"�- 4)hi�����ӿ+gQ�,�����Bf�Ğ�X�;g
�Z�L��i���"2H�e��>k�y���c��@���¨[�E�QdŹ��������oT�Q�����En�l�/5�@�R���hWR��(�U[c�D8�HX9�%
"U�HOA� �*ۥs��5�Y%��0��L�gr��f���B�wY7Ke1�VXF���k%H%� 73&���Ⅺ 3�͐�4.��孕#���J���3�EŶ�#�M��Q��EF����K3UlŎX��ڙ��n�b�k�;åEFf=��\ӎ�0���)D�e;_To:�ju�ۦ��{��jS��J[B�Kr�lt�v�bB�t��&��ne#������k�]L��-�7Kp�T����U�B��j��y�,e����Hûow%:�&������%(sRy��݉��V	3rd֫d6)�\�{St�	��e[̷*܁˒���x�D=%�m��y�����N�ل��ն����K2�a��MA��\�J�v�9�+E��"ƅ��S��@co)ɦ��F�r�g"��n�E�^�&�#�O�
��+0��Y�`ͧ���ksj�ȅө�m��.֚t�F�I:�&��]$n��"�e4�nR��EJ,�r�Щ��gN[�ySP�M�l^L��ƭ1�D��z,�Pe���Q��w��o~Ӱ`�H��%��n�i�FH���bu��/q��1�R65��s6�e�XT[k4B�˥�nR�v������	�ʱX+e&��;GY�l䗷�`�Y[� r�BfwX���Jl�������/!����1���q�_+�LۗS,�Z�+ib:sq"�A
v(ԩǍ�`=�Ep�tʑM٪�IL�wy�ndLY��i��\'YWK�� f��w�Jԫon�[�z�x�Ț�t�"��`b��b������
�L���&�I�c�P��nĸ3]f=:�1�$��bjť$�ցcr���"�>Z�d�݋�j-Ǌ��e±<�1��C�H^��-�m)a7$(�-#hJ%�v��{�+����Ub�^Cf��1G�02�%a��u����y��n��[�yzV�z%$�ĩ�țX�6���^c9&bں�I�Ht��X�,1Zs2��`����1�e�ڨ�$E�Fe���*8ԁ�2h�Gn3cp-���+J�I&��ˤ�X�Pô��kD�i�Vb��v���JX �ba=p]�\Kt��f�Ӵ�t��.�^Z��)�C*cZp���º�zp��`@|I�[@�![�-��&�M�J��2�oP�KP���:�a��rU���mR�$��]#L��9uZ�bZ�j�h��<��Y�f��f���yf\0n��_6rݠ©d�V��#L�Z�)M���S/m��\����ͮ<���l���i��{6T�d�7`��a�jl���oŦ<��Wj 9h�4��G��$����l�LA�/E�SU�8���i��e O��i�{6��u����S&ys7�CRY���)��x�)xn��.eA7E�C'l-�Q;���8��T��2�W��ۥ�L���N9�Gel��4ɵ�L6�L*����V�헂��PF�� ̣f))8�87d��d�����b�býql��:.�cp��L0��,��_G�.�K!J�12m���n�Vb)0.��X��>�s�n���S'�sFk3��1b{�
E�u]K�x��W��S�>�۬�
��mc:%M#0�u�4hf�D�y	z�oz7Mf���V����RX�q�x�k/4�e�A�2��V����.⥱%��E�uy�T��M��aseXӺ2��$�� �0��d�T@�z���l� ��6S �LٛW.�WWFU�I�Y	U����E� ���P�]�յ�0VY�Ɖ���N�K(j�u6"�!�4�]4FFi���ָ�`d��e���GQ�m���r�b��Wn	�q��VM�ć?�M-�X ����lgm�NP��'^�g%躣o�0֛G(xU�-1Zm��O@��cJ���!nB�L��X���{�`͹xê�4�n�p!�#��Ov8^hRe�*��VG��],6m�*m��r�4���E˝2isn���j��t,�֛ݥ�bŜ��6K̓j�d���4�y[{j�Ѣ�m�n�ݜIY�.hH\q�25�����-���J�:�f�΋˩2�k�6�:��v�vMLQ+ײ�R�8�;gdY�Œ�G�����-ޘÒ�Swz�#.C�Rdږ�J��X������Wx�S�.�
X�{sH�����0����v�Yâ�\�ZD�ONb��b&k��eh��mGt�Z�i!�t5i�D��?�������d�)��Lېޝ�י�M�-�Y�6&4�;O^;9��:�6E	Ҫ�/�ph��I�z7Y0����b	�q$��7E'�Ar��
�S���ɛ*ͪ1���Y�MV0��n&��֨�Yg�CiR����^T-���BŘ��:F�^1���aVL��B4�+����V
�F!b���JhѧlhP b��'1�z
4Mb�����J�%�c:��E�Q�FpJx��o)���f#���*�V�寉tF��3*�����r�B0Gy�L����96¼�V\hA5�+Z�9�e:�p7ː`X[�.Ordh�^�V9
c giܫŨ��k^�L��M'�gE荺Kf�v�`c�q唊��>�L�@�O��{0�11�8��F�J�b器I�."r��!��N	hT�5�B*f��<EwajU�(���q+������4���d��)�LR�m��,�>Č������v�8�؅&�8v,���s^�\Tv���݆	t]7Z'��oXP�Z���Q�eV]MX��rK�IP��<�N+E��B��e������9xj�#�#�p�����3A��I����.�IL[�#v�`�^�w>��ĥ�W�X,աrM��^e�1u� ��a�bŷj4(�u�v��w�m�J�7��Lukp�.SF"dp���&�ˇ5i��C%f���$�Z�*�j�y&	��zBЈ�t yt�ͳX[���d�
r��u�]8�v�J�IdN�h���KA୕GwkC �M�E���a;f ͠�-�Pa�A��q��6"���]4�ذ,¨ ����q�CU�����Ǘ�oM���w�a�I!/q'{n�b�Ts-4�rKTÙ6�;GA4�i�-��ܷ��p�vХ�L�.��:�ô�IA4]m�:�m�C,��p�yB��Ń�Yܓ���`7�H�jjE ����X���R�V+Vem�����;Y��B�b����B[bѭr�kY Y�2�BM��T������Ld͠��/��`�i�rr�n��V̥l�A�o��-S�nU�`��q����p��]�z�OC1���	�YR�*,i�l�(�fޓP���{��a��a爦�Y�M}<ΝQU�n�N�,�ŔVN�M�{D|C�]�z]3w�)��B'�9 ֪�׭�71���x�fU� i	��4�k1TX)�Y�)S�[aޥ�-�.U�
�U�3.�(�{��4F�P����UKM���'No`ǰ�`='�Sx��h���ʯL������6bV-=f�㦑CP�C7�ciЕͦRĪP��1.+�nU��Jj�P�\&k�X9FC�O)�%ZM ��n�^F�2�Vv^�,�$Dc�M�O2�[� �L7f�շOn0�iA�RЫ�]��mm����XR�̹� P���1��nGH�2<	�iȕnՑ�Jw)`:+oV��7.�-��#1J �s4t��ДnU9i�>��yr��,3.��RĤwC��4�1�m6�U��/+%i8-R�F��Vh
�(E��0&'���{cP��$k����)��/K�r�Ѓ�0H�q陻o�
�4��i]Cqb�3)ȃ��4�����`�����kXZ�Q�l|2�|�ޭN(%d4��A��sBӂ1�ɫ&��%����C$a*m+�pY"�Ґ� ��Ŋ��]��L�Z���<n�VS�kgr&<�|���^��NQ�!��O"c(G����Z���6@�5�᐀A��W&'�f��qn���fC�	�0���`��jw08�<8݀l�Y��LУٖ���4�A\f޲�����뿍'3v֞hJ� �O��A-��v�ɂ���g):Xnֵ�P�xe�8rhje�Z�Vn���H4����XܹV--�u%�E�w�y0/2�xd��%J�
r��	.U�{o.���X�CJ�Ȳ�)%`�w�o*h<XV!n�e���JR�ę)m�3�0}2BBx�(�b��Q̼�k[�R���E��E��d�M�v:o)��!S�v"�U�HR��E���ejDk�Y�X(m<z�!�ٲ�Zz��)	OMZS6�j�;�t��/�9o�Ǎ�д�];¤X�^�������eM�X�4mj{m&F]�CEal��/+$ݡ�W��3+���[J(pL��Ő F�R$*�V��Y�7m��]��35V`hィsR&��m�( Ϋ�^IW���f/��Γ:�;s��hXFR�A���	��rس{��.GJ��T�WM^R@I�k[[���R�����
�6�U�lE�k�<hb�XT��c�vXfB��jR��_F��&��򲀉����7M����$��[v
y��E�2�މ�6
�@VP
:�ve��]�wS�; �Na�9�b۪�z��*�LW=4%֝[E���V
T�ה)�:U��l��l1fD�-����^Ǻ�K�/o�Ո�cj��� ���.3��l�1%�7�Ԓ�ڲ�5*)�U�w��Qcp��U&� ��V(^ۏ�u�t��-B�S�
�jOY�^�����(�� �N��B�)��klҼ�M���Y70e�I�F�5�mm�^�h��j�[X)�si G�VU��N����64���A�ܨ�F�i`lv@4���ج}tVqy��)t�|i�&+�)Re�w��[�"�!B�J�d�n�C�ǉ��5�Ӧ������*n�ҩ��|�*�F�62]n;ƃʒVR5�-�kB��hY]ѫ$D>��������A�P�v�|���UC+u��ڙx�5�X"��n]7D��ԫkl,W�5W���+dG�.�Y����t��!���S&���G7av���p#4vWV��f���bD�])�d/�{X�[�#V,@�\�Z�n��%� *V/�;����92`�uc ���G��B�E�h��nr9�N��yy�	��,<!�TN&`Nk�����5c2��U:i1�ƫ4���*��]flYkhRl˹�e�ۦ�A��Kb^���KQ�i�a�������KV%vg�^� ,��Eձ� e�E(div�5��j6���ݛd��Nc�n��+����oR�{��j����Q�nݵWu����V�5�$�2їo�3!x3�����X+i���!F��q�G#B"�(m<�7V��I�<��>ô�bD&��{Aj�Տ|=����${���ý�D:���V�j�?���;����S���x(��v⭙{���$�5�lߡ'/U�O3Lxޣ%Iޗ���NU�m eֵ�#�6�L�6�o!��qA�&�i��z/C�=�:�'����`��Eô]�*��sM��b|@/ ��P�{WA����J[4��I:ID�y(�IʻNKppF�\��Z�4eՅ���l��>�m9��Q&M�v�C7$U{n��a�C;y4,�5wK^�Y/.*�*���5+Q��m[PVV��j�:4�r��`��
T`϶|����u)Q;QǒH�z��7@���e�1h(��=�-�źk-U1w�=Gr�J5�[r�ZKk1�H�|����f��<�dɑ�-{s�mʚ6h0�KY1JS�r5�����+�9q��؜�c����7�nib̢�z֮q���a�@yoa��[\C�(����)hV[r��i�M:�/�oM�}+q{�t�b$���i�� Fj�U����SZ;��H�h �N뮇�g9�*�4��/[=�HQ+�t�;�7bW��pLژ؊9m+۝�2]��rZ��!.;�ؠ����E��P��w%�(b��N�M�CN�l���Ȏ&��VbS���C�:�+V<�"����w�A��jn�=�ՓX�T����d���9W��-�T{��Wy�\o�e�f��ٔ$/���g遡�w@v�Ϯ���Gt�Ь��jĝ�t}��^�F
�O�A���s���B�IQ�\�cW˱M��%�r2V��˽T�,zL����(z=�8sTD&��cε-J[�c��^���烨\����x%��~�[����.n]��b9{��'a'Q�n�{���%q��E��l;=�6�y��5t�L�_���v���ȇ�`�57�����8�j�3F;'5oL�7�;�J:`��k�t���g-�|��LPoX�5�.���i�1b�X6n:n�:�W��Ʋ��L���`+��\��J�w_���'�ݾ�������B��b���L��2ٿ����n�g��m���:���ky��c�k���5�Z�4
Y�������g��nGE�����ɫ!�$y�;��T�oed���{b+���w������&F:����Ј� e[D�ț)�[�fmvv�!�8�<��t�d��W�()��vN�xޱ�s
OZ��R�1�5����Y}g�@��d}�
��6M8�7��̻�XN
����Wu��&3�j�sT8�onI�ڵ͠�e��*�.�t��y���ћ��J��_j��e��:��-�{�=
B��E�m���o{����cc��I:�+oX{bA���|jھf�;A��>���޲�K���Y;zb�����)����X�R���p4M6ի0�[X�)V;i�/]�J������[�ü�gp�Q��;�F_7R��X��7U���+��u��rsur��q�)��;�ظ���k�$g
v/4xH��3Ӽ3��=]Y���x:���W�]	h������Ɩ7��A=��g�BÏ;,��i��U�I<2�����t��xa��.Q<�NV.NꝆ���!�L�&t����ʲ񣖨@�f	���<���OԔ��)-�e�n�lx�7j����rsE�=�s��
��o��b�	���k�=����~�!(�3�ҝ����U�5��~K�Jñ�ޞJ� 5 ,���@�E�o��U(2�bAR���/��t�vd��Y<G"o+�`I�Aم+��\�W����tz��Sc� �"��*��y�ܡ<N���-nd���K�Wm��D3e>�d�+�E��:7��Q�H2�i�t�I�C�C(��%ng��wv����T���8i�9��^ywz'i����G��8�����c3��O���Y�H�DPZ;�U��)i-�ԴKNS:-8:2�V�L���7|S�V�R�k�wCrPm2�d&�c���unRKa���U�Vݽ��&�T�v�52V��AR
���.��m�O�:�"0.�΁��cT�R7��};%�}����sW�x�1D9�B�h�$�>����>�SXqP�]� ��z�ǻ�i��Mُ�ҍ�Ougv�@'R7��'��"��/"�hnyTɧ�������D�2K���{��vOXB*�9��4��Ws,o\��`4��"Ƈc��V�@�U1ہM��a�����7�U������5<Vs��te�+'YPu��X��v
B���5�����huL�K@�͙;I�u&z�}�ޞ���j�AU��+`�GN25�b9p����{� 1�z"�X�2P*�%�)$A)��'T��o�9k8[�{<�'1���b�� :�ާڏh���&�}l_@3KZ�{ӻ}�gU9|�)z0S�OTN|ok������بv;���L�����~Tv򱤙�������{�ʑr3=�,i�~˚9I��o���[�yP0��E��]v�Ns�Q
7�zf��%M�^yK12������Gֽ�~������r��*� ��@�S�IiMe��|����r���a���;MC�-�mL�'k�7�(��嗨Y �8L�۞�b��T{!��y�GU�;s�d7�w��T��2̒7�X�.��5�Hރxw���5�48ㄜW�8i����ჭ�z���w���u���뮨�	/+�q��#X7.��n��]'ċ���J��qй�30���W�(����x��k�;er��	�+������[��Oy޶�P�fC��B|���: ��j�	�׻�t�+*Vf�b��ӭ��ɔ�\x�E,)ǙQ��.ǜ�Tb�w��cܸ|�'5!V%,�jKx�V�`��e�h�����4ÛUOM�W��С�7�!^��>�*�ug��J�[-�ORų�c;	��� ��]�m�xC���P}ONܧ�mj�:έhe�����a�=�[t��5���Qok�iQ�f��Kkt�Ө�����Z��x$��T�!���-a�IK�#4g�U�:������b��,��S���{�bZ�>E哄|1�!%ͣ��H�p���� �l㖨sep���9�QD�[���M��b�;�ԔM��ϟ����4x�jy�-"��K}�1=}�A^�%����<���!��C0r�c�����/yo��es;�����T��bs�xYܷ�.Æ��[�9/k�u��TZ˭lVZ̺�Rde���[�5�c��{��M��K��YE�������(�ީ���F�NX�XE�V�#Y-�ȃuS7���=�TFn�H>���>��]�Y��҂����D#V�o���|
cz���Ig�N�!��;�R���%k76�M\Y2J�ĭ�}n�)���̀p�c�%ۅ^�$��MQJ��mo�-̡�.m���()ˬ����+�Q���S܇y�D$-���75j�dtP�^�}�_B�/�چD4�ꈕ��#r�U�֏�j>v��*�F{B;���k`�u㛎�Z�#���>�,�{�M]�.�]Go��8��%܆�$˃-��w��H����;\w[��%�qY6��8DO���^�"c�+��28��|��,��|C����T�Xo�TdDI5�m�+� ��U�X�F�	�0q.Ss�!`�ghX���'��0���:v��!�u��;˺�Z��~��!����$(�yO:����x��G����������t���Vi�/o;#�h�����}��X4*�=��C9�#Ψ�� �5޾���%�[��=9�h���z�$3U5�^ȶ){��}#Bݗ��>�����)����;[�~�c>l�v6:�u=��7:�k@ھ��7;S;݅�j�����qW-l��u�KCw�8��F�52�!;i��wK���n�C�=��QH�TAthh�d�_^P�_E����Gf����I��,/����Y:�ö;
nK��\xě�ҏ>(̗���ΰ����][{5��;|�Җ]9&�m3٬�������1J��A�ܾN0�Qy�Q�zG�8q-^��O]��x��ܕ6L��32cѠgc�>�xˏe�ѯ�k�^;�� �`�zc���)BT���#;si��C�su��O�3X�y��:����m$�b���Ā�wm1w2�٥�Ewc��$�r�i�k;`��x�*6��1
�)XmfP���CKlY9Q|�MwO楇Á�r�˨ᖓ�w�P���C�dM�c�y��~���#C�z-|�}�q�^�T&�h�{"����1{k���FZG)�R"WG�[{�C��t�)�$��h<�s��O���M�C��>�Ҏ�a�	b���5���i͚s�4��{B0yWX�ۺ߷Z����P�M����!�f�yi�R�)��Y���Vp�I�)�0�) �����"c0Վ'HS�ٖ�]��.j���g��L�.tW�$s(��Ƹ�c샷9��K/��1ө"=)��8��(]7cktS��Phs0[����k:U�\Gf�)���v ��iJ��Ы����X��+��a%a�q��-Ѿ7^̗�zpp��:p��*��`2���d�wu��ez�F�D���s`��K�GEeE'-���LCN�D��=� ]Mg,��D�3/��r	Mctz?'=�|
�|���ؾ�E5�"7����y��6�=�F�M� f�6��@-�vkWְT�������z��R]���վn5+WS�U�c�Wx�@�ӫ���zv��WK�)�m�<�Q�Te����ic�Z�v���T��vq�T3��ݶy��[�&��}mK/0��5[M+z�:�6$�}G�\�FUs��S�Pn=	Q��[�� ��L=[�V\Z"�1�#���6m�X�����65�d�4��.��)P���@�V���{d�:5��碕-��*�|��}TAUtp�f]MxVK�f�#Ed�6�QX�<02��3���kR��Y*C*��P�ʕ���TK���h��Y��ݮ��L`�+�9
&:��u��f�o�u��:�Tp�����
�	�Z\�
%���]%��)/9|�Kœ�I�''��<�HB���Y.��ẏ�}��Y/����S����K5��b 5Q҈X�L=�P�*��g7%��«���W^�����F�Ȯ7�Y�@��d�� 	�/h]��v���t��n,U���s�b�v����ݍ��g-�l���'1�j����uk�ư���"�kс��e�7� �Z<���M�H�LZ���f"��_
ũ<G�BQ�u�w"�*:!�ŅX[�[�	��P�i�i����2,J���êR_���"d��P��y)7��Z�)�.���ԭ�@�{1��;!8�G_b�WȈvj���3�K9B�oF%WkL�\�l�o^�"�]��v�D�B�X��"��u�mh���E�Y�qf���LN�u�V���N m>W��-�S)�Ҡ�V�s�K�LJe����it��*���ѵ��C��J��I��u2`
a���C�)���y���8�7Z�3=�* w������4�&1���r&��pC&ܵ�d,��c�p˵I�3��"�ȇP\r�;'Q�n�
x&WαŢeu�0@�,(p���vS��i3�mr)���K���c�A�����U�';�o1F55��Ȫ�B#YN����*�ma��
��x����&��wO�.ڠ�5�+_�ϮV�F'[��
�光�L���Q*7�j��n\��S���E�3��8,�=f�J#q��v6��G:�Z�Ol�ŕ��I�l[���Q�YӉ�P���8Z�V���w��&����&"���ҽw:5�s+��嘳+���R�<
��7Ab=@ݔ��U�@���F�Y!] yNK�7���
������r�`�z�.��cGeה�0p|��s�T&�'�J�N��,�=�:�p�f�^�n�}�����n��1�۾�]�U�.*O�f�D�h�zMD�9} ����˧a�n	S�;Vn��F������;ұ| }���/��'i�N[�'w�^O/3�����`,��%\���{��c/�8�Q�}�X����r���Y�O4�������X8G�Ē�e9IF��^�XE�F�NPjT7�1�ۺ��"��(0*���R�ї���@Y���Ȑ�mg�#�u�F逫l��J�g��i޲�-W��@^𚎹 snkB�p������w�U�4�C�Ɇ�����`�]�V�v��&�x.xBs�Z9v����c��L �d9�\%�i���*���y`������.�nS4>��׋�1]��=����X����q#k�*����P{0(�9Q�H�D���T���/6/m����CXs����J͢��n�5�V�M��f*�� \�Ѳr��wbA}�<J�sU��{F*�ש��5������tϫ��������l)%!��ؚ���,V�gg�p�(� }fq0m8������n�m�"%�>��o)�1]\���3FFi>bhS�A�Y�*�#m�n�g�wr�J�y�a�|U
7�:�<�ħ*���;;lq�B�Y�q ��b�ݎvp�d�Ux����Z�n�.��\!��}�q�)���G(���!�F	AWlJ�҄ pk��Z4.�*T��L���jU���4V9������$���5�_QOa��)�AiRp\��Ū=]f�K< �1� �glm��N�y��r�1�Ipb+8ۧ2s:��0�52�)͙�}��k��w��6``�{�
�Z��֝Vz�au��ZRT5']9���[�rG��EZ����JR���v^�+��R3D�$�-7�7V��(N�?��jة
�8��o��؝ڬ���[���+��-�����u�n�KgIHUm�vs�H�;S6���I����f�J@��Y#�g���3����E��*��LR�������oE�]�]rT�I:8=�=W�����h��v>r�o��U_��)W�ڣ���A�V�����P{ð�s_e,s9�����Z#л���x��)쒌�[u��S��Y��ǫ�30F�X�;w��]T�ɶ$��M����������/wf�����I��N��w��ڻ���*�t)?�u�y��Wd��Yf�א+��s�5w-�r.co��Tšzoo�a����w�����Z���߇3�~������O�����$>���Y뮏�9��'�-���ǉ4�����m��oF���r�k>\C����$1X�^�r�N�|�1�*�j"�"�h���}�r��t[���ˀ�7u[]��e+�l{��)�لg^a����4�5b˴60e�ʎk�_rJr][2ct�qB�=P-��ԯhep�07sM��a.����s��u�v�jC��滽�z^�;N�f.k[�4r�GWwENX�v�M1�W٢U�%�'C�9m��!�6#�7�k7ӝ����	9ܷã�L�ܥs�`ή��J�s�H��Ү6�f��B-�F>�f�8Cפ*R�^7&�����xz[-;-^CH��j�| ��Mʵ>�U�؃�ltY�YW�{ӄ��ܛFm���1$�/�QѝL�ݶ>:�Α�¦-B��7(�Emvk!�C��V(�s+S�S*8��7���$6���X�7�F{@Ub���g�B��g=Ȅ}���pZ��1=�p>��XyV>�ݪ��<s��B��0��DO^��!t�[���ݱ��[�8^���ԣe������+��9n���4�㺑tK���y:��{��F^vg�ZK9^��|׽�*�p�㴎�����7�M�_=\��EJB��ܱ�c�F���״�9tXN�E+�a\�����U�`��;#Yg�եfո��F��Bۓ/���ƭ�[��>5|��Ӡ�b���w�h��=�A����@�fU�s�Ʒ]밨�VF}/%�f:}y�����g��V.Y�Z�%c���,�ˇ�8�ժ ��B�����*�0���Z�"�U|�;]M{w|S�f+r�����8�]�DVS����3N0"�;��J�3����N�� 井�`=&)G[��B��cף	i�tp^����-�0g�޶�.[�u�	U�~�\�n"��*���+��=�h����&�x���>�]��к����ډ�Br�fo>u�dϲV!���#�;bJ���qn���y�yE��ȥB���Y`�+�pnv�Jz!�R~Ĺ�k���<a����ћ��R����|����q�6�f���溓L�@1"X� ,'\����a��C�ŧ��� �����Ukv�O��jq��<I�k��7��ێ�k�I˓���s�&�{WJ-�&.+I�{G}ժ��T���>��l�bm�-5���Cn�����)�]
�d���$���V��ܒ�Wwc��H�ڮ�
GG�q�*�'�\��t�Ѻ[��&��P*�v^��]�Q։��N�����
���ŹR��~���z�M�V����A���J���l\�e똩�u4�?����'D-��ו�Iu��=b��W��TH}s�{5���frݮ�����]�o��@�n�j{�hF�$:۝��72 ���#�z^��wu���wa���*�ζ�đ��,�c#9����]�(4�
�.��8�a�Eꋺ��ɽ�#L5S�:��Y�*�Z\�;8����M�'Xc�o| �&�{%Jh��.怜���q͙�;�x��E��LwP�!��:�;��MS[��Ga6�����r%��zl��9�1�_cDe�Oo�P�lI-jD��]j���%bd��t�|E:x]+�x��qi�ĥ�gg��B��I&���X9b�l��5����>zG���2�|�8;s� 3�i��=¡��c�-�JGӼ@��/w��T��gU��MX"r��m̠*�fm�}z),.��dH�Go���tX�����.�C����;Y&Ҭt�ќa����m���-4�����)L�ۢ\��_}uz(�`��7��6��V�٩�uJ巎��'jGPmI�����-���oL.��gc4Q��4p+���A��c*Yה���\�ۮ�/D��H���������������Ԧ�P��^J���u<B쾺�|�(��䫜�K^�._	W@*ZǓHZm�ܢ[������ʻ ܭa�2����:o2T{�`Xh/��H�G4#�}>y@�dZp��s�¦̢�����/4Á�G�(=�y�� ��d���1��n(e���s�H,۳uܜ�� �1����=���Sq\z0��Y�J(�ۡz���a�,Y�B/!��@&��C�Ӕ�u�W��⧒��m�KmYO)"(�ӄ �E��0���1�z����e`	�n<�AV(5ˢ9�W��-�r�`��V]MW�廅��w�d����#:��_:�����q�&��>�Է��] t��}�8��U���`fK�mU��j)�숤�W
��n��Mc��
������u܈��y��oF�1��TXs�����7tp�V�0���y���6|{�d�>��^�|����5�gu�p�]Iu�ٝ'R��L����-|�J���9.q�ӈ`cEx1B�#��[N�/����u�Z��r̬�C>����;סx�=��}� U���,�t4ghEh�]W�HJZ�c�Sjvl|��ˎ�<�T^MS���a|�ڻ\�߱`�㹩�v����(��;F�Y.�_�U��.����T�4j���!�K��{ϲ�μ���1=�K�����ݽ��٭��]WŨFY�o�g���Q~�B�mk��q�>d�)���3�u)�,��\tZ�!7��u����óOm��0SБ�WD�zB�g�4Z����-'��WJ�Bu)*� �a����mP��7�d����및n&�J/ 1��&+�`#��A����F����Nl�WT�+��Uɪ��1�LC���7�0z�.U[4GL5۞��kr�s��Φ�#�EXÉ��</��j��������ʞhO6%��	�8��0�e3g"|�Q�\.njy����E�Uw�"�){r�R`yyM\��:�̫���[�T���C����he5F�_io+)um�J�*H�rRv�S�mp��(O.�˖M2���=;��_�bj��mdPv-�뾏V�'��_Ky�۽����F%wڈ�pb�b�v�{1zLg���Z�U��e)��_!n%���v1��H���/ a.+t�0�Ei�9�2Cf?5�!����@����|5�$�0QWS��{�����[�Dm����ה7]p	�c�AD}�Z�z�Dh��������z	>9*�h�����f�A��h�������3n��$�ؚ�#zU³]�N1x#6F�ov���t�Ҁ��v7�d�8�q�p��eU�M'G#�	�{�fa��%��]��<�F��t��s^�p�i���;�۝�	�k/��z���˹=O����_g=3 a�Y{@�8侮���I�(�d�I<����_\ ���V�j�SlV�}���<3��I�*����8�
0S���˓#�3�4j7�kC�2����7�/JD��c��3�sf���d��G �Lz6z�.�F�o{7)���� -F)�^N+�����w{�����|m>���n�U>�ܵ�f���3l��`������c
۳xU��>u�A��eD��}��	O�q�r��k�_?�j潥��|{�Y�]�����b�7]evL��=Vl�y�ԡ[%v�l�Xܙ̭g!�yeku9��\�»>c�WjL�R
�_��WQ�;`�Ɋ'r�+lYU�7��J�}ܲ:�k챙''j���13|z"�1/8��DH�Չ��o�:�n6�7D'ӷ�36��7�n5t�j\*�A����km��бi��͹a�0D�`�:h������`��LV���w�Vپ�T�_p�lPz������E��Ŝ�>�]|��T��P1ҨT���\��-īN��Y��bX�sڼG<M����U�c���k�)1�o�]st�� �#��N��?<ɉ�p�Y�-(�mh�5ئ^�#�d��[���@V�T��Ж���T��1�2r=H��ŕ�V*{��&��Y%#a�;�ۀ�l�hK딑�����⟖s��ZZ˱>g&9h�<����P��B�u�{� N�h�y��L*�En�8 �v[�3��sv��2��՝dX��q:����;	�j�+��Ś�TP�5%jó��c\vWeb{8�y�T��W3�MR;4j��0��T�P��ٸ��X��i,��х�Q*T ���z��<��V�*+�Xh���]��>{@^�n���sN�8h�:��
{^�|٥u
�0n��8���kt�6!R�ͱ���pKt{{�/Y�8� ��@z�'��2��4+�@����{r�$�X��#�ץ0��AӞ�-�W��Tf��ZR-%�־&���%� ��}�"�5O�ZnsA�����s�Ɣ�a��r��,Ө�'�aj��p���lGݡ��V�R�t��p�,,�
aP��: -���;r%ۇP.%���N���.es���}���og]��;��-�u^�i9�t����L���3kܺǸ&��cS���]�����9��aP쨲Fл�N���n �^X����M��L�Z!�¶�$N���z&{;؋���_�S�b�ܬ``:�,E�wR^p��R�6�����S�`��g.NT���s"{4���!�:�l��Jh�؂.����*^[�-�o7��GI��T2QJ�Gj�g7[��]��϶s��48��n4�\%�Ӏ���1S@�l��绖��H����j�S�Tg�S�Ć��A�3���C��`h�q��wwF1Z�Y�m�{��̲zi]@o��_�0�������ا@�K�{r���/{A��ʨ�׶P��Ub��	�%qW*{�6eI�21!��w�.x�W��uã��C~��0�s~����fK��t�rɇue�(^��u3ԫOd"�Q: �gf��Y�:<�ۊ��89<��AUS��o�v���b��6�7��궶��E�i��3VWR�U���h���ç�EKk{�Z�]������ֹbz!|_]�6�3U�Xj�ܝ�Vɯc'e���$mu��*��(��[��8��܁�/a;�>�ר�.���j�'`��I�jm��:�Q�önx^k.&�
��C��\�f�
N��R��y7�r{�sS�6wk�黧�RңB]��J��I�*;z�,+EY�����6���9�Q_a(����	�Vn�nuPɝ�8}wٹy�,����f���V
ϐ�q5��ee�T;�7��:17ٳ��]��l�vvd7K$��s ��M��GN��e��6.��O�����#�	N���v�n_L.�8�j�wF��7�*wr�W��@x�}m�&���}Q�o{�n�ٻ�mh����W������
�^oWe7�+�5j�P�ا�o�nW� �Ṱnx�r��(��l��{F7��O�Gv��A��o;�twNX���%�=��;f1΢5x��H��P|Wq�/;VN�����-�h�h�}٢(��PL�G-9��u{hHj�똊Ȁ}{�j� �� m��? }��-p�ً:��/�5��DsL{�(�U���s�Vb��.�1���l*Tl��O''�d���R��!9��1S��{�ޔ�̚��}��G@I�bP�9�[w��|p�9�ڨ%�bIr�d�!9j���o�Ԋ���E-�(���AF��]��	�+��*nG6Ո|�2�qh�W��:��;>�먲kJ�!d���3�p��]+�#V�c�]�Ђ�c�����M!�y�=f�s\�2�V[	�	���'(k|����4�C
\�\d�BOM���k�UϜ�kܱ�(�ғ�#�tmQ�C����%_�Vom��X�r�"��A��jTQ�đ�f,L49�Λ�j�2���ڹ�.�6n �nYgb���}��"�
ԌL���Y�w���a��/��@�9��iv�i�
�������V�I�	_T���͆2^���P���(� z�)�z>�$��P�]����RU��{�؋�mѮlM��餓hD�8�i��7Js�j�J9y�f$��^{a���	ý�72v�i����e � �u{�9B�����N �y
���#��R�S��vU���Ұ�{%������G���-{�I�ыn�뗽Sd��v̺��l:���Ԃ�)�;�T�{����Q噱	��0nSS@�2]f�F����Z:�c��M��J>k[\�Et˻u�/L�k7�ӱd�2*{34���D�rnUw'G�u�U�Pe�g�>쾺���[�-H"oGŁ!˒�����)��=���'f�VP'��x���ٕ��Nb����:���W�3%��]/��%u��ά^ݳqny	h�-����)7�
NM���P՚�e

Q6��(*r�V���M�XfgGO1_c!�.)v�N�fq��ή��*:�r�y��<P�>��J	\�ؼm��yj�A]��b��\h����Ә��U1A�5��V;-0�lK�&��VK��odI�ĺ�ș�;��6ͻ�(��n#��#���M:�S�\ꈸ� �/�e;���,c��[�⮦[�)D�ߦL���Ӷj���ڏ�s���/�;�zܡ��SF����r�	65�z�V-��İ���B۴/T�f��k&Y"�Q�'8�����:��7�\b.�H�I��6zApڶzw�[/�w\je���5�^b�b[��)������|o��1�����)v��&1��Բk��Cr�R�Mȷ}a�f��+��� �b�8iL��s�b��� =��{@i��d�y{�seE��h/،Q����j�����*=J`u�;{I�P���rC�r�>c�q�C����m�+�\�Ն��9(3Y�ce�a��d�S>�ϫ]p<J+����0�l�թy#8K�IC ��݊Z��:lR��4k��5V���U����U��!\D��D������b�V�Զ!s(T��y����n��s,^�v	�dXB�RN8MjZ>�!ۨT�f���~���ɤbg}���[����$���:�������Xcm����H�x�:A)�`e�T���"�Q�yl�<C<Q�X����H�"d6%`'�WwQ�*K�;�9�a����j�Ȅ/u����)��cV:𡌻���*I�q�\1Q'`���Et�5r^����r���Z�e�b�
�@�4u�8�Z7x�m��ٖo_XH�K��zG�\�w,Ym���ԃ�Na�C�-U��rjP�;�{���4m@�D�X��%GBr�O7��WISpun�F DB�7wr}m�Us�b�J����){�(�W���A;éS���;��Ne$�֌[�̨���iS�%�M����yj�%8��m�<*�@�x4%�����'^ߴ\xM0��8Z�"9q������6''[���C
�����q��$;��w�,��]�n 5<�@Թm���$�do�e�ĸs�:�v���}q�;�yS�q[�:��*��R�ٔ��o����O4����%`�6s0Ʀ���]��c*D��M7BI�wj�n�r4�k22Vi��2.s��'Ǻ���|)�*�PQZ�b����q��YiUem���J��֐�**
�m
 ���EDDA1(�Qb �Aa�4�V*�����F)m�b�TB1QLr
�*���U�2�DDX�6��1q,C)Q�X�ZT���
�Z�(�+�����Q��j6�W)X��Z����b���
��-��
�R"��P��+m��-�m�1V"�+b6�QUDD�Z��R�B��D��j�h�\���D�+UX��E�؃��YDD�Tأ[�����U"��KJ����*�e[X4���E�PEE�Qڕ�TQQDDDY"�J�F���1�b�
�E"�+UaU�DR��R�Q��# �(�DTF��b�����QQQVKj���,b��6�bDc�PTF"6�Z�(�-�"�Q�
�j��=���{����o3l;���>e[�eO�݇�ny��R���k���o��ފ�k]���ʜ�*�|o$7�ۋ<�����}l�98]�u��ҝ��Ӱ0^��Lݢ%u�:^�y��;�Q��� <�3�,�a˫$�S�i`P��h�����D)�u�3/�ά:9����?���������9�Oh��&u���ZՃ�Tŀ*��9�з�.,^�G@� kUd9�̑��xhh�z�b��.�cl���Q���S��'I�\t}��o��ƣ�J���0c��E�INw�Ng�m��u���>�u�=AN,ۀ�6���r���Ds���q��%S�5�x��{ѡp8�j9E���p;PU�X�%��ײCun&��f�B��V�mV�}��M��Ϣ��EԆ]t	��sy�p1F����Pz���1�b�:^�q�_{�����c��p�(��*2�K�F�́9��j�pv��O�K�W_7BO�_M�B��FŸ�<�J��3�ܟ��>��&>�����X��j�s�rj��i�{ue���Sl�Z�L�`f��+��4��K��$���C�"�&V�D�QF��,��4P��T��s�~U6
w ��Y.D)�.�3^�ڮ�Gs.J�W���K������n��W�1��N\��1w���i[Q1�.Wݧ��jG3V���&�>��Ȟ�wk����i�]���Թ`T@G*��!d3���L@�l3($�l��ۀT�&�W����獗r�Q�w=<��:p��ˁ(׆՞����x��*�+����X�ֽ�?}�}�ڭ{P�4z�O���	���K��Δr��#AÆ@�N"�pt�$v�cvU�sS��Ѕ����Q%7�\`5���'�Fe
����.]F��Y��uN˒�q�r���0�܃>��k��4�.v&��z@nnc2!����k�nk!4�pw����W���h�Fp���9}l��[~���-�E��@`����7�#��Գ}B�y�|֍��Ė�u�(�S/����+RD�n|�K���8�u��	�Lq�y;�o���Ǣ%�2�z���ˢ����E^��V�J7Ũ��	�򖣎S�v�_�N�LDr���(4�bB -"��g���;�$3X�
�z��D+3nM�]�[�wlD�����§݂��QJ)P.�%\�<iB&�x���=э����=�[%��5_$C��5�c��/�|6���Y�V�� #�-��X�z� @~�d�⟫���#p�����T���r�=s�y؃Y�Gg��ߺ�v+��"�J�l"�	�v��V*�y��gx��e��]sWu�Ӧ΢�Ge�wwo6��+�n-�*����]yڰ��w���Y��P�L���3��
Ac�ׂ���|V=0�l��;Zz�Cq�ϸ�����bk�;ǐ7Df,Εn��t�]ϳN�%�;�Zu��A��E��|�C�v�.������	�*��Lk��Г1��wl��[;k�GQ�F���O�x�)W[��g�ը�2��d��_��k{;"��9��c�>⵰=^�XP��υ���<U�����1�|mE9�x��~��S�¦+��z�@F֐�Q�*�/�1X��݉OW�\����4
,]SUy7�t��YE�4�uXlsB�d��^�A�^ɐ��ȡQe�u��@��z��oe)�7ԯo��<�*��v�(����{��dX��Ɉ��Q1wA�}6��-�s�!kyj�#}��P(K|\=w�/��y�Z�۾�?MW�جZ�������pKWd���s0�����F��n)dRN���vW!vk;)y�w��>��e�/Q�x�尽0�"�7�p�x�˘i^>�%ۮ��b��9"�u���C�{�zת�>y��cVϨ�mL6okb�|�+���ش�@䧉1wz��vlE��>���@S]u��y�;��+Wa�b�� ,��(�{!�����s�s�xVor�ܰ��'�����:+�Ј�:e[��Y���L"-Ȗ��lMaR���!ʺՕda~�����`�q"�:	h��9�]
�{5O��w�h���w�W���K���a�nː�#�hf��+������HEO��q�	���j��^�}|ŉ�7	�f�[55�z`�C�lױ�L�F��Q�� B�
����.F�t}��"Y��<j�.���O�zl��9�#T��9�K�-�}��ת��WY �������{��Z��6+�ꚐC�&T���P�V�.�U�*g�-���t����>��m����}*�&��"���$�_F��+�>�؀�u3�Q�8d��(�KP��r��۞Ȣ���}�!��L5.��l���o0HD?
���&�W]�$��rc�:G�� ��gcpe��4I����6'n���5�ŸXfnW
4�sJy��2��/���1�ű���(:����&@n��X�ȯ�
�2���!Vv��wx��q|�3o(�А��Xv��m^%ӯo[�R��/i ���#�*�M�=�;˘X=��t;�o���z,T>�kGu�	��ݭ�9v>1F�@�sm�z�����^��-�^w�n���&�מ[���߅�����ir�ʣ������m"�*�"Gl�prr7��/�Lm@j�Dذ_F�f�v�-~����v��]}��VPR�8f��"���:���ʘ�ONe;��k䅻�o���o�������4��	w���F�w���u_�<�<����q���n�j8��o�Pg�9� ]b��QX��י��7�A>��HU��坎��w5�ٰUCdi���\	ѻ^�j��"��7�ɝ#j�QcGTp��wh�m������ͽ�n�7>���b�t�d{�42����K�K�a�8Ϙ^ٽ���Gc�gGlAZ!����p�o���^*�F�	=���Sӽ☁����7;lf�oݍ.����@��_�c*}�^��B�<^F',������
#�v�	���
]�R��B� ��~�z.��!�Y�G��nj
��B��o���o�P���������<X�O�E�Q0nA2#;����t]P
G'}иފ�F���.Dt���yB���.��Z��#1O]CJ���J���ZW��"�"���Ef���'_s�e���-���@�;:�2������[�IM%�|v�<*sfo�{�z�˝A�6��n��}�5Y��:c����$v弉I���`�!�(��)�	G�l��W�d����V���^X��a�/sf��Rt����`[�0k�$���0Z� 0>����+;�;&;y��k����uC��u�T)ҍ�Se�XI;�q쌠�hI5�	J��G"m��f��v���
�`���P�(�h�eT%ʝ�9}�-L�4�X49�:�v�5��o��m��䯪�#��_��<�./�<�hl#��Q|6�tK7�3�\�Ѭ^T��MGv�F4mD�K��p��j�٩UO�x?��%:��x��	���/b9&;�yNC��{����~��;~�|�E{~H�;:Q�s�o����2���pҬ~�)�IƟ��N�X����U#[��0�Q^�n⢍�<dB[[U�<�Ts��}�b����
gqtN���0��@b��&u�2#��띠E`T�})O������|D8qV����e0n�:͍�)�00A��c��O��/b\�N�H^׵=Q��[}�)O,[�:����$7��(������m��3ڭ�չy|C92Lsf����ӃJ˗�9�e�P�8�!o���Yʜ�Ƿ����9U��G��s}=�^т��]�A9�8�2����5�ʎ��Ši�x��ڲ6Āu����[��J�QN��]N}3Q1 �ɽ}��+U��!�t��2φ��*��s�v��n�N8u<nw/�#3,hO��o9%*�I��H�Ƌ6P����Ď5�,��{~���\iy�#y���9U�/S����gS��-��(ӌ0�53�Ҩ@F�(��je�N#��^��0�ͭmպҌ'�E���VO�Ɏ����K�g�D�D�r�<��������Bz��Fv>�J�'��0+eC�����0�w1qI�Xx{BJ��`�T�諪\��u˥1��J#j�3�z(�S���L�㭺�m��E�Bk�;�p7Dhd�JV������z'�c�N��0�i�y=;�Qӥ��S��6 -P�R�p� �@���Y�^t�wa�]_�sBsb��n`J���'�!e!����8�%����9���j��u=�	[� �bc];~!�hݞ�5����f�+�t�Ľ�[���ļ}������w�Ν@�5��9�a���"��V���>��1��,`���tY��z�h����ũ��p���UIW9��i���ci�.݃�J$����%���!�ڽN\1C'ҍ�[�`���[t�b�oj��(�&�<KyxRM㣼�o���g]�[� vܣ}�B�p�2���h�:�3g>W'GFvwU�An�]�u�ʀ�a���=4(�H�tō�!�2p�a��B·%q�zɘ�-��r�=�:v"X�6]~�P,.�u�Ȃ4Ror�C�U~���� ^�<�LN�|�9������ᬌ(��L�>��ъ��׵f{�p��^���p���gq�e5
��g�-@R+�	C[|�	�m���͜.�
>YO���YX��e�x�H\�)U��ɍ-�\j��=p�!=09���U��Z�!����s��K6HU즪r�	�7RQx�*���B�#vZ�!���q#w����KGΑ��P\]^��@�:s(�B����9��Bp�*���V]o�!N{��j�Ht�T	fT��m*6�R?^�������v�*�Yé�:C9�ݩ�b�)�۩���L��v�K7�ʕ�.Mq�k�2w ߪ}�͜!q�=�WGBƨ�쐝2�ӓ�؀���[�S9o�u��J����9q�I���D:�Au�����rx;s��SEӭ�y$���	�=�K��~YѾyPGy�Ʉ�`�oc)�C��\�M�p��-[���@vV�"��Rk� -�N����Ua,W�,�Re�mǄ���؇
�v�Yź�������Q�����]u��ۥ����:�V@7��㍕f�d�Ib�sck�A;��$Ԯ�=���/�N�tC'1I󽔳�L y�`X$̭��eJy���G�g5��Mp1�t^��M����Ҷ�:ѵ8�}�`�s����Ƀ�b6�3�_A+�Y	��؀�.�A3t0�gb��y�z�PJ�b�cu����(ߍLExs�p�D;u&g�����!�Ŋ��o��v�Wj���{�U��q���d��o,_��l�'������.�ƃ���]=��{${���ß��)��'(�ˈz��<��#{��`���S�Ӂd��:���p�C7���P�X�9�NՏ#��Π��!��N���9a1�)�=�Yk�ܗJ7�s�c������7DC���p��Pr6i�6��HԕQ�Dl	��e�ܿC���u�A�}�Ax\K��v둯
�0(\=�E�=�W�*�u�9>o��ʌ��Q��CWTW�Ve�k"�߇3<v����.0��R�(�����l1Fؕ�z�k��'��)�KQf�@ù<�\	�l��T���J����un��Z)�N!*ZO�ա���֢r<M�X�h92�n��+���~��ʽX��|�X�����7�_ ��W�qR�{�t�{�)���'S��{��p�wū�#D�MRt���
GW>�[��+/�V�aO9��ِ/�g��r��;�^�<�qS�xz�NR�j-�D���fOT"�Zr�q�n����2���q����M͠�����xz7l={��^�fm�=�'��3�w�W��%8À�R�-�ze+�^F�e�gq|5���dm��-{pWӝ-��5���"|ym�F��@�?h�p�C���K;�W�Oӑ��{V��g�>�:��s�����Au� ���ʽT��gr���;Y>�Q��s���"S�u�%���QBvI�"��H=��;#�b�+^�;K{v�ǳ$l9�nob;v#b�n�A�y[�G������G�f{<����{��i��ԫ�cAp���눯B�(؅6\Bq`��`�1��J�0��k�ރ�j��v����?)�}}�۔��.����b��6Kw@�YX�Ds�WS����M�Wy� ���'jB�2y9ˋ ���l#�:j H�fRN�e���a-�w�7�#�ܱ6IoW��*����b�Ե]�\k�d��x�C@���e���t�/D!��Z�=��E�)��͵lV�
a��LP�F�����\��h=�E�\��is�W�8 �=�K8�sW�wu*of����Ad�iǢw{`�E��|�;���K�Ʀ��\Oh��R��=�T�'�6��MWol��W��Q}��G�\���O�����O��M��v�=S{�V�{/�7-�6�8o�:�vB=�"�]�fП���l�l�}���\���hL	<���}�"tE�^����f�|�d�92�v�/sLo1T�^��#!�M���ob#���o�rd(���c��N��R'[g�o5�x9�n�
���0�;΄W@�k\%W�/?X3U���z�t��C�N���,�l5�,t���i����˃&p#�h(Kf���B�9|'R*nD��*T�Qھ�}���cg:��\��Hv��S�f3Mg]ef�05����v�|֐g��wQ5��MJ��nj��\�7HɌQ���f��Jd�.�_j��wsN5xn�#�k1(�`����9i�y��l���&9K�a���xz(�b�I��V;xE4�$�M�FJ9�c\�� B��������C�	}u="ڦ%���;Pg��[��;mK]D*�n����w*�.s'K����ެ�&��i�}���\�˾$�ө��0��ӹ��a���9If�u+ܰsfc�m�C~��]�3��#��e��$h�:0��#<y ��PuZt�1��ʔ>�HQP<��D�6�m!�b���tx�&{�&Y��Z)70@��hI�O�-�B��a��DX%7q�
�3�ڙF"j��_ڶc�Ę�!Zi����x�a1+2$h,6ڡc�-��]
O�ҹ��C&+f+U����h��?Z2���SLk�����/.�9���u�
m� ��Ǎ�����^\X�V����*
O�Y��Do�!vn�L�F:B�Jqܧ��c0�0S�*WtYU(ݛ��2�=7�C5�i��S�2�'�ۤn�j���q��DYب�b8FF�y�mڠ�D�
�Ck&.�Dm!o��ǵ̛��h�+��$q��j'��e?�溌�l��a�2��%<�-�N�hKm�8	E;��#�C,����4(��:�t^@��p2!���������@��hĺS��ay��4��9�M��h�O"�Š9��#c��5��7mf֚�U ����n4�P[Q�N���
��iԜwjm͂���V��F�⦝Ѵ��p��0ɴ>F8P�(�Q�tСQZ�5ͩ�k-�X�Q,����7j���Y���F�*�b25mE�*"ŊU*�Z�*+
*��*+TR�� ��UZTcʍj�JEb*
���(�,YX�
1U#iQcl���"���X��PDQm��j��E�AB�eQjX1b�QT�(""�����d�,F-�QT�E�b�-�
�*4XV*�jQb��jB�Q�"()mUUTAm(���%k$A��R@[KR�Eb�+(���(,
,PK[*Ȣ��Q���(�,UUQ,Q��RTDTTJ�2�F%���QX)-�VUTV[`�Kh,��A�PDV���#-������#VKJ,��UAb��T������*��PU���YѬ�*%B�lR��X���0g��_+_2ʖG���
�o�vl�{Fs8���-e�g3�Z���܁Ql��h[�}�-!�LKr	m>Q��>��S��{�nN��n����;y Y�|�ϻ�q>��Lt]ˡ�cJ6���8x\L:��D�7��E���4]2�dA^N�(��LF���C��IO<�1G�q�x.�����t[��6+a�A������#�8�{���=��z��������\�D��_�&�X��n��:l���D�����I]���f@Ϻ������K<��q��!7p`9rD�j�uE��yXTD�T�s��>��n����0�7�F�o.+z�#�b7c�[���E�8&'�q#��g�^߸�J�͑w�5�tO�����3C�V����{oMJ�d��rD���U�!
�3���+�a��s���Ɨ(����תܕ�����b^Pf�z�ҁe..�%\�<k��Ȫǰ�X�5�I��"-�j��S[vb��mY}�HޞO��!����</hIX`���*z�=C!�-t�D���J��q�k���2����Q{m�P��9�P4 �R�ݤ�(t���:u#к���g4�M��>�P��k�eN�[B�����#��b����x�]m*�S�]2�-uK��]+o�D.��9e'8p��h����	��%�e�u���o,s�s��� r� ��YSr/6���+���N�����R�m�~ŵw.���]~�"�v(GN�� �U��=�����ў��ڥ�@PK��><��VX���A�fQ����f�����	�3���}��%��o���e:d

h�Q���e&6Z���_�xW��2*�<�U`�1;��=����Y�+Z�_)uW$��!�H�,����9���+�3HO+"!�U�c�V�>F�f݇c�qE�X>�&��B�,�;+��q�ȭe�k��תy.6��!����ݡ�ˈ� @�tlʁ�]T���DRo.�w���9p�by�Vb�B'�oQ95�V+)��0��xd3���2���z���$��[W�Y���:"9\�;�����j;�異=�-@R�+ʓn۩=* O5��kg�����z'T���ӧ�sm���X��]�z�>v��ƣ\ٗ�c#�x�f����p;.2�R͛iB�V6az�7�٢,;��GJK�T�Z>#<k����=<��j�/O�<�\��彖���np�:�ӥ��Yn�QQ�P��GF��=����P�D4��ŧ���-�a]Y�D,�n� k�M�}jgT��}<�6�	V�b	j�P&U���-+����1���nS����v� �ܓ��iq����G�bJ�/���RV�����E������{'�lns�+�ک0��X��tو�(_7B�e�sx��p�����	��:���p��B	�"���
������h�8��;z��<[��F�qs����� #�2Y�JGB��g�����zko/֟�����N�-k�]̐�"'\X�(^�L�5����!Y��sǓݾSqW�.�51�b�:nc���ӵP0�b�B&��|��:
W]�S[��fzx3�E�Y�/C��x��4�ڂ��w�����YcG�Ϋ|��Ah��F����f�f�&Y���#FEzԇ�j�t)�,9I�ݻ�:�q��ί�^fg6����J+uWKn���e*��{<w���=s�HR7��X�J�4�M�g�Ը��C!�(a�e��u�i����ui=+b���p��J.@UPD���P���&2�X��B������u�棷��C�����\��T,�E�19!�4��2F�l�1�UHٺSƖ�lK7yu��5�\˱��.R�H�^e �+��j��I�w�>�r��`�Z�F%\�z�shѡ�&���`����7�ч3�ڽj³����]D��X�0Le�]Xc�	�Gzἂ�2�dHV�L\���Ju�Q�����z�����h�Q�k���cR�R�4q]u��FlQ�6��3�f3(+��^�3qB�8�<N����恲|6t���{�����_��j�莌�tJ�vt����~�1 �����v凾�녟{_T/�*͛��ʋ�#Mb�p&Ƿ[[De�ˇCGv���w�-���6�E]�Y���37a�a;DY��!�v��b������0TǂY�jؼ�Ŋ?=��8y몢8�!t*ɒ�ЋQi�q�P�CM��e��A��kw/	��Iv�Sou����OTR��Yƥ>]���݊��!)�/��D3�Bw���c_�IkGj�i��%�1GO�'h]zbGhK�qb�G-���hvFX;�[����a<�OW)[��Ϗ��|=hD5��Ԓs$k���Rt-�]��T�&dMurŅrk�VH�����Q��0�'����%�ܣD�mΙꋤ��#�DWQ��9��Ql)�8��
̆��#�;�V��Q%"�|��p/���ꇖ�����Hny����ۯ�J���	oo��}q���0�ٓZ�YoWq*��0�yb�ˣw����0!WSs�cڢ�+9�m�\+���MwfЫW�VD������y}�Ki�݊�f�	�<���ʈ�*�s�k��9/S����"�1&�뵨\{��w��ˮu�Q�
l��Np����00�\��~F[���:Ym��f��C�	������Er��$\�������}�<���e]r
�Ռ٭3���bY�3�qm.��y��=[����ց�W]S�T�'�m�:σ�<-֦M*��|)<�\��خ���f|vJ�wq����}�i�Qj�5*�Y�JuK��4]�bros��x���g�����m~����>��Q^�g�a���;A�ҍ����(,�1v�T�����s��*�c���B<������'"f�	���]��q) �M��	����:G�zyT�o�u�UM�WB8�sz���~�K�
̑f|����t�����>�o�oz`�1!��vr��������L|�o��K���yl��'�It^�ʄ��P�����+�b�2��u�V����7�IJ���������S�ںuъ �G9��c��np�ѩ��"�t�B<z��R2�ƺ�¡>ۍ
�Gԥt�+�eXc��I�c�!#9�w�X�u�s�9�u�v��D���]��)���c�Y�h儨�B�^i�F�T���V���W��KX���0�JY�ڏ��].�.^%�sV�/R���Y�������u��]�ZqM���{�;g�����.muE�J�/���H�rʹ�΍,�m4OJ\깜�#5Е�����5yL�$�u
�pT0��3���/��6#��E�N��s�� �=ˤ�^R{w��"�r�n���>T�_��;���%���ѧn'�;v {jH��I�h8�#��ũ+���w�]�Yw��T� �g�X�G����!�u���Q�<����>���U�y+NAm�L�e�^��J���X�$�i��Z�>��0���=D���?YO��nv{Fr
Tn��\���T�z�7#f��n`U-�����FP�C m�nH�/1������r�W9J!l�n����`O���`�c�
�!߬�)�j�ۉ���[p�Y���}FF�>�E�$��)�$��ob`�:Ez*Y��
�c������ʾ�J�װ�Z�v=W'BIl�~��U��a�g�U����+M{�V�1�M�#��:��t��l�r랚w�8�5[�\����ʧC�v�J�~]T��$O��J���zMcY�a����q���$��f���]�qh!�Q��K6�J�+��͓���Fr���ǫ�"�I��ɱиu���.GKg�xTp9�殝�*��gLC�N�*�+���/r�S�*�w����{������N��B�������l����SQݹ�O��v룷�^�XveU��;5p	MN�u��Iw�Q�rWtVj�o�*��a��=�Df���B��(����y�1�I������wf.K�A���s}Q�]�+ޘ�N[/'���K�6O�EG��nrB���6!)�\*����g;���6^����U(�|�`�I��T���_cC�誱l%��=��Ѳ����*�W��{�ؔ�}:`���^!�⛞p7*��gX������L+�
)��X�m=���ü�{��"������E�%�;�����C;��28G-բ�fTz��l�R6���_���m�F��6�$���ڽVk�h���x��p�!�
�F�H��J��9[g<����92��(^�,Q�MA�����*��P�=Ў<��X��{w+D�wÕ��u��S�p3�)�E�V!P$�{���8�	՝��"��"��	m㾥϶�' dnV��C{(��N�w.�x��W����F��[m�_�} +�x��W��X�fd�yc���2n>�b,��I^���fu*����ّ	W�0���OF$�TTK�+&�u��3Yt���w��o*�7��.އ}�pC�f��V�;]V��a��,U>�92���u�\��+lt�@uyL�`k$U��t1��V`R�V9�Aٳ��>~���h���߳e˗x��J{gr�����s��z3��W�}_T*�Į[J+ q��C"u�bVݨ�S�_��$�m�ɵuN��k���̘��63b҅�ޕֹUI~�;�W��q��=}�{��NR����d���
�j�M.�U!��G毫�Y�n݊-\1�~X<���ؓ�I�{<�h��n��_C���-(�bS�^D8}"��d�D���Ѫp���E�M�3k���Am�o!鑳���mtt����������(剟qF��#^��(�V]Y�8x	���,�!x��u(fyתo�g"\A�}���cUW�o��=������FؗD����tg���u��k(��
�#a�x�N0s�o�7�nH�,O���Μ
�k጗4�ƫB�����vo��Ӳ�cn<Kᷫ�uu��z$n�x;�?3��c�׳#����o@&��NI����ס�I^��V��E(n3<�{E�h���<�CD��C/wܺ�}����+_�3Q$���Dr�3�w���BqgK�}R�'��磦jQ]�9���.��y&(�����Mow4�-
}�`w�k�rk9����(��8����b�qB����2�k_  ����n�Jc��G�:D�p�(sqP� W	�BbB$ԹJ.��q�{P�F�vmd�Ǎ���X&�1=���!���9��F�%Q*�h�M� ���f�9�v�C��y�9+���UGP��(�F���}/�̇QK����};&�y���h�wf�ͺ�͎�J��lS0�+��8ק4�V�>��lB}@�~,�q@�����e]/��)�硞��QkgH�S�����Ntx��^��jv�el�n6]م�tb��$�GT0!�@��-�"��^��r��q�oŐF��ܕ���f��v֓��`�U��28�n������z�`�:�b�&	;{���I�5��s�x����; o����m�#�
�j��|����J,Ot�/�n�^vuM�w�0�E5��z7�﬙N`�|�O���qw?S=`��gv0�!��Âz��(�j9u/cN�׫@ȗ!�ĄuuS5����	ȅ�LF���3������D�����%d�$���f�:��G���^�����j���z��y�x�O�Qc��� ��lk��n^@z���'ݻ���'�:���g�������FN��j�A�ؤ�|����I�����2��RZ��׫5K��<< �ՙ�c5�KD^�5èɎ��1�l"g�X5�����ͺvP���K(�rB<@x݁�Iƣǝ�_`�G����1ts�/��y4��Y�ǘ�^��QPSL����-�<�q\��O��\V����kL�p�]�/+���1�Q8�nI�c�H�S�ϯv��݋�s<��鬌b�wE��:��B:҈G��=B���ˉ�C<�Hz�fە��cmuN�!�BGt_4�#���*���8S��=>\�`�%%�(��v�$뭙�w�����,�g��C�Y�b��w<����3�;*T^�Rd��(��g[�y�ʕ&cs��{-��زhT�9x6p�Nt�ܥk�F�_6�z3��0��2�b0�!S������U�p����s�L��B<���c���	��5��W���ϧ	�h�˅�V�Gj��0�iTH��X1 h�� v��Z�E�G�U���\�KOm����q���}�e�&Ԉ�Ρ��F�/f�Kha%8/�Y\��}]4��U%L�$ǆ=�8�Wʭ�1���a��J���?9i[�*F�0ń��8���,^C���~�m�A�t�i�Y�=�;��\X6r��FkU��f��_p�3�g�na�Ghrv@���I��<�������K�SEwi9�]�C�.��i��j�C�X�9F��� �Nl�*O��k�6k뒜$�J�+]g=�Wu�6f�e�����e��ଋҕ�v�Uҩk ̢7�D�d��u{�޸��]�SA{^ξbe[����1��Zh4�-�R��)�+j�q���Z���6���o5�noȵ�J\���d����gU�;um�+��1�|�k��ڒ�^y�z��v�Kxz�;,}/�z&F�@�������ʰ�o��"�J�C�G�^PT�����e�4**1՚ܧW��J�\�Z�t!�|�=�/pL�� �݁�te�0H��R��)k��Um��yo=� ��!��f���<9��BO��HbQ�3���mK�pnN7�s�2�x����o��B����=�|��ޙk��fy��B�0ve~4�"��G4�j�ķ�:�����n>�Z��U���әJ$�!��v�c�.J�B�X�ɶq�8��htz�{����������^���,*�~:QN#k�9W���^�hO|/�`����K��g-T��nP張��q��~뚧U�g�!��&�x9�7L>X�Mm#>�x��C�xۿ8z�	Y�If����|�7���MJe�]w!�U���sK��H�n�AS�˟݄�f�_8\��h�q	����a��-�N�uF<j��an���q��l��S�d�A(˃���P|;}&3�5�7����"2xK��%�dՙb�V�'����D�.��iOq����+$O�el��8nƌB�*��U�A5�E;���#N[�ts�����\��Y�\ϔ͋s��DS�,��w�͟w�Q}{!]܆�՛u����k�)��۠�D2���u�A��aL����"Nz�(����h�Ĉ��VA�̩�Q�[y�c��tx.��b��g/�\���k#�T`k���I�x�5Hҁ�1��+��/���j��-[�ͅ��jӋ{K(e
0��I�ͤ���M]Ouy&*,Op�<8\�{�H��ޝiN�л-eh�MC(�\W�k�׈����h��`	��~3��xU�-tN��u3�2��(���'��ٹe�����a��6�Y�}�>�o��lă��*"������r*�I���溽�|�=���<z47����&�^U��)��I�]U�`��&��ܠY�w�^�2d�kC�ʹA��[��hՖ��c�_��*saz�Yx�f�� e�{�9YĵY�姼cc^3#����؅B��N�QZYW���ZK=N0�pkۨyTye�t�Wu�6��%��M�x��{��3����^<��)�<u���ku'��յ��ӳ&'c�環����Yׁ�K��֖+8d�ѷ��r蕋Q-v��7����`���g�j+2�z��ڔ�/z��Fk�Wh:�I�DHb/�N��b,X�YZ�j�EAjV�DX��D����*����XdPm�EPc�����H���Uc��b�b�@UT-��X��(�b�EmT�,�Ȣ��b*
,DQT����EX���(�
�ł0��Ŋ�
#E����(�H���E�"���Tc�Ab�E"Ȋ�Ȫ*�((("�DD"�H�Qb��)X�"@D��UH�+�1��-��QF(�
�-d��A�
,X:lU"DQ�(��QH�\�T��9ePr�@Q��`*�(�EƖ�UT�b��)D
��-e(#"*E�E"��Vb�J�Ur���*���ww��xs�g��B�B�WcQVM����k�zv���o�{e�0!��󨯙[w����b%�ot'}�L�'M�d��}U�W�-�!w
j��sЙ�F7F��k1p�$@7���|��R<whj����B�\4���V�r�WB��h�Ny'D��5���b����vԋ,�e-���^֪!����*�_�J��D��4t�E8!uH��6��Y$vY�J%��[Z�+G5�Hn��3Brs"�i}��A��*��ν>�mr�]��꿼i
2��e,��1{{��ɟW�jC<A*�B��
�NȼR�M��L�������j\33��Jq;�[�����Ɏ����$X{�Fa��
B��7�[u<اJ����R�AQ�Ա9��K+���q\���R�)}�������ذK�����t+Epf*���#6 �E�j*��M��]�mOe�����oʥ������9�KfOr�r��+��Z!��e��HB��l/��Fs��&�/}B�t���s���4C)�7<�nR��,JΕ��hV�s@�}Ǒ=]{�0e�I�D��t;ެ45L��݄�Um�®!M��l�=�&l֢��,�i��E]f�6
݊�]��[�q߽{)�M�ѥ[{�	�L挩-��{����)��_T1s��	c^Gy8�J�%	.���Kk�Ӵ�ޠ03�u���]��9��g���HBJF�G�   �['�'�K;-��C�h�}����I�&�k��)Uf�����-(F���dU]2񾦺İ����7.E�"R��9`��@"�qQk�zW�v��Ws�)#Ĝ�0=����:���(6'�4[�G_���]{6U�'�F�$�uFD.����W�M��;%����v=椨}�بS#����0�t컻f��3}A9�
P�F�m�-�_!t����ù�S�u�NW��Ƞ�C�Yv��[��d�m�ɿ+��`�v��$OY/T�+�6+R�W�j�̸{�(�����I!Hާjr�_Fyӡ�ߍ�Az{e�{U���%
�uAS!��98D(g*-F8�:Y��wV������r��lS�\��f��ۜNdw-�:������lE��d��VC"�)�U��R�5���֒�*Y����vq��a
�<�F�>��-�;��+�g#
p!��,���V�ĽC�rIk5f��y)�>���/����jz�@���^gO�M���m���y�W\�D��;��A��5���v�5b<��藩.��#�:v f�r��yn������Sˈ`5(�ۿ^JJ�U�p���y�[��tt�;�Y�8�.��h�zb<W���m��՜7:�tIT�;_W�B��:� нJ�� � �Sݯ)����$X7�m�2L��N(oUo�6=�!b{voxN�8�E�y6��}����,V�2,
��({!��l�/�U����8��%x��}s���"�!K���U�J:��8��}Esଡ��)ƫ�U�4{a(ꄣNp�CI'ۚ�3�r��+\�]֨��O.G����H��Y���Qc&}�ƫ�Jq��T7F�UQb�u�R|��tNƱ}O���ݔF(��hꔵu:��*� ז�kDG�T�]C�ld��Ț��K9@k63^ѳ�P�%��Pg\�8gDvE#`��P\"Q� ��"��q&z��rk����CU�!P��(�F��4�#~�~����>���J�����Y�pI�������T����wR�Y]�'*��|�~�GK��P��Gf��x�S}�fۻ�xu��h2>��_�\qCD'OB�F�)��<��&�L,�x"�2h)���m���M	&��ؒ�/�ϔ����0�P�n�G:C�,g�w������7B]�41��1u���Ԩ�p��Hیt6�rcP��^u��7*P��n�G3�C�M7;�[ϱ��o+I�Kn�\����7���t�NjnL��l�dɹsC�Oz��쾯�H*ܗ;u8��8v\e�n�g|<�=��W�ն9lb�OG�4y��3r�F����HX+(A�N����f�F�F�������Ջmv��눲���5�%�S>��P{��|]����b���K�y��y�v�|�{X˥/��>آ�کP��I3�?���}��Gt\},���5���x�QX��;���N��mֺP�r{)�8ᬇ�Bp��.C��٠���gn0����Q�F��2z�B��^��tK*/�M��/������H�3Ԩ�/����x�ؑ�UO���)dzW�ܳw-T��|������3SsY �g�,j�t׶<�3m�el=���xv\-ڪ{X�IP[<��S;�(xX���ٕEk���1�$����v�ܺGֱ��5/�OS"�gG������>�p��������!�9��2�ƺ�\4\����tl>��w�s���5TD�bCqa4�#���%m��4��b�J��(����<�s��{r]�Jmi|��p3�.�h�o��H�7�%�� ݇�>��u�(�ǆ�9;�Ş'Ѝ�gݙ��x�R� �W�/k��d��=���K��jsM�^d�w�)�ذz����g5؅��=��+��O������P���n.���X��L["C:�>]**y��9�ݗ/I�7���Gq ��FOa�Z�u�O�b��<<<=�����j5�Q�I9���dq4J�]��]9�+���5�#v,m\�`����"���N[�Q>]г�����Cx�:�����d��H�B<�%Y�/��A7�ߝ��|n+�9�F��2:�1Kl_
iu�����%T�Ќ3�X�L��}�2�y#�v�@5xv��-F�Yq
�n������Ob�����Q�E/��#M�:�	��Ͳ�3D�����6�-X�Č#N�j�c�C.jd�2�}^SN��Q���:}O�z���=�sҰ����姕��F1�G\P�2N'D���h�pL���LT�,�aۅJ��4Ҫ�����7�����)}{>�FB.�Q��wMK�#�0B8"(��:�������u���;���H�b:�pv;99�b��}=L�D���t��J�auS�����bm�.�z�*D�]��[Rb��F�
�YL�u8k"��,��R%D�1���4�;8䉅'�أ��^��M�O��r�,V�k<��1y�ٮM(k_�!�|��Z��3�	r����ͷ����5�q��n1W��oWM�x�$f�����>�F������M?g0[G��j]�Ee�ݶ�ɷD FM7o�?:�>m�H��f���M���W1
T5U��:#0�I���H��yŹ� �|WV����j�v�Mr͇d'�k��Ť!�jG܈��;�o��_,��}�ɼ�BXz1XU>��z�)���O�}�}_s��c;(���JUl`Y� ~��9�/��.�f^~g.Y��0����F�\�m4����=W28�fJ:��*c����ݴ��u��P�F��D�q�R�jk9'$sܽ�˒�>�W]5�+���9�NN�t��gX��}rF��y�2�ʷ�'}ڻ������m7(-:�������AS;��#���(�n`��/+^�v�hs����������]�Jk��)Vk��>�ԻN����M������ig �z�_G8`��Qj�U���>^�C�]�	E�!�rA=Gj���ÓJ3�Į��~�8yBb8�^}pv�P���05a��Ө���k��q�<�^R]Y��Z��7 -b�v�]l��i�������������#��-�]�z�#�Nf�͕������QM<���}b����C!�
��q��2yro��f��0'0|{�g��Th?�������E�#z���
X/���Dv�Go#S�4�	��P����{0F�s�z�0�Jf�����{��
,��=ѹ�OlW���a��-7���&�/����2���&�.��	���ꇅ:sws�xc2�`��1��!�������y�֭Έ�ٸ��%=Xoe��Ȱ�����ȩr�,DY�s"�T��F(�YH��.򛾲�ݬy�ڵt,w$�z�r9>�62o��0f�P�TkA�v�5^�]�e�~���iEob��;X��Q�i26i�69bJxJ���/�����3Ղ=�|�㿁�l沷<Ф^_m��v�₟���j�@�q\�I��͸jda��JǱ~N�N⅀�Ef�UYy9�zMVs�נ��\��T�������
>+/U�`uPgry�n4�B���;�1]��]L�G�����O�UqY�<EdЮ4�TSq��8㺉[$���/��[��Tg>��:�����d�W�Tt���OK��ERa��<%D�����g?�a���^���+�zl:��Ÿ}NY���ݔFx�DO��h�WP��t�� 5�NDx�E4{w'f��o%f�ъ{'Xx��.�r�uv�9�H��䢽Q(���^�L�������}+�Y1`���摐��Ns:8@B]�w��I���Ô��L��U�qƂ/���,��.����9�(�.p��tQ������>��o�^}�&z���tK�w)Rn���p���t�I�!�1XJ�	W�W��f9��x����I���#Հ�g~�u�T0���P��Q���,ʄv6��3��IC'�e�֍�z�����>�}T� ���]��>����b���z�]�q��2T�O�>�w���'c�;�A~d�0���Q���I��a+N�������)r�>��
�Βb�4�J���$��	PĊ�vg�'�AH��q�l��~��4�ĩ�Y���$��7�&ߘ6g04��^5��s4}�ޏ�ޒ��:	��^���~�����|���>~`6�O�Ï�� �I��i�
i
������ri��f���&&$�h�
z�!����=a��T��d:N�W����i�P��_D�${����*���qO-}�룗3l�����d�E����w����=d�Ru�� ���}a��i ����AC�X_l�i ��~7�&�Pĩ/u�C�mbȬ�aO�0y}��W��q1Y5��u�]o���z�� x��2T�l���W���+��1��2u��+�a̡�)6���:� �+��r~C���f;fn�I:�2��ό�0*�����H)���?z��߮�t��׾$�I��cya����c�z�H/>L��;aXk7��f٧�1����?��J��!��6�HT�������&���Y�O����x�@@3��ײ�n��A���+y��~�0*O�W�d���X�xL!P��M���K�&:w���^0M�޳I���H)�*�{�v��Y�z�~��I����p�1!��s�߷�����wG�����_|�cP��ʅ�L`V�ĕ�~��&�>J���p�����9��>�5��� �X������3��*|��;H-I�}��a�:�H{Ԙ����*�Q5�?~d��|\���O��ϟ���>�i:g�~f ��*�w�<~I�1�3�B����3Y�i"��Rg�14�Ɉ��0�
������CIP+�~�b
E��|����eIs/�݋��3Z��%w�\���]Q�;�25��G}q��se;2e�k���y��6R�KZ�F�s=��U|Nw]wi�b�����Ӻ�B��91��dc�eL�X�[���ǎ��WNZ��	r��*�!�;�Lh&�KNor��K�����R�������H@dNǽ�1��@ğ'Ɉh��8Ϳ0*<��z�!�bA�g�*��~LOMw ����c3Y�H/<��6��`q�ޤ�6�^��~u1���>dt�{�O����]�
#ȁ@�'��j��{�0;gR|�=}<�h%O�w)�^0*O������%~`T��bE�J�>�sP�~d��oW��A|`l7��u>C����o��V�l?��{[����ҷ��,�Hda�PӦ��|���1*A}?|`i��C�c<�rM<C�1��?s���x��P�%v�2b�^[?$�x��9�p�t�̼I��H))9���~����H���QIߩV괧�S�Ԃ�̕;�a=}|H-CL1�����Myf;`T8��!�I�p��i���jN��?'ӽ�Ă���c滇�iZ�&}��"�>���N����!�^�SD	>��'��m'�+
�����P�vt�YP�1�����8�ݿ�'����:�>�*���u�N3�2{�1�%T���g��D4�'�I�k �{V���]�4yU���#�|a��4��@�|�钲��c乒q1���f��i*&�0��'ڠ�U�Y�N��O��&�8�>Owa�L
���X�d�1�������1�bk>�kEgo�<M�z6N�� �1���;�'��';L�'Pă�}�@] ���y���5�g����J��)���C�>a���E�ơ���r�3�G՚�]����՟ ��ޒ ��\͡�K��'�����2��9�&�R,P��0���Af�<���?~��$��c��SL7��q�PP�9��x��H;�N'�6������φ�ѳ�=�M)Ͻ�2G���}(i �a�7�,�R,���������d���
��ְ*O��*�{�{l"���a��l
ʞ��m�N&}d�d��
_z��1�r������=9~����Y����'�i��a��
�'�)�����P�P�Ax�ϲLAv¤��2u�%eO^��@�+%e}�'�1%B����i?G�U �}�>߷k�}�q}�/����r�I0��VԬ�'�
J���Y�h��j���'�O�K�gNȩj����'��
RCb�w�����c�!=�{)lY�`��-�(��04WA-v��H��!Z����J��ju�[�"�ovu:t����}U�{������o~��4���m'�3�J��T��'�O�a��1����i?��i"�d�7G�!���3a��4�^!���kt�z�@���sf=@Z��@�� 	2|�>��?u��]�;sϷ�}�������%I���Z�`�P���si�0�ɞ��E�P�k�C�~d���M!�K���봝B��L˧��6��b�C;t���}dY���D[�(��C�ە6���:|�&v]�h�R4���,���z�gg3$]0*
h;�<M��q�{��Sb
%w/rjO��h����Ax��ε"����I<B��Y1<��8�a���|�I�x�o��O=G����	 �=���q��0*~~Ͳm!�Ϭ?{������
�I�Oڲ~e0/���Ԟ���k�&�RUI����bAxɹ�0���Ă���!�6��-f*h<�wz~��[؇W��%eO�����Y*j}��x�Τĕ
��P��u���>ϐ�����>d�O=��zɧ�<9���2z���v�H)�O��|`�|Ͻ��>u���*�O�k>w�����O�����K��}f$��~H���S�c��_����:��*�&<B�S�;��4$��Ow<2�X�<��y��3������ q��nj�'�����#km�^�&Ь���Ͱ*
E��a;ˉ�O&X)�=x�s�c�z���i�������P�VgS{;�sa�1�P��Ă�'��F�����J>���7C�YZ}�5���I�4ԋ'O~Φ�i
���ɝ͠~JÌ+�5@�M�X~ְ4��
���2(u��<`_1��&v�hq�0+��P��e}d�'�A ���>�%�m�S9���=�Ͼ�`~g�*����<O��Az�����i����}�����W�8�YY�F�a6��VL�1�8�V~��E�,j�O�ċ�gɹ�����}��~�]@���-��X�[��~�T�6ɷ��{�(i��������_�����a���ɧ�����`9I��b��&��-AM�{��kY��8�!�*xM�1���K	=�wW�����;YS78�j�|w�ҫ�z
�����v�o�����'˗�)�#V7Bs>~�Sۄ��T�x<S&is�������eX�� G���![�v����}Z��].7��`j*�L���t{\�{�= c$1�&R;���P�fN����mQ�[�q��O�IX<��c��v$�@�ts���7����1|��@L
b�
�2lqb<�U^���e��8�G�;b�M��qq��ֱ՘sj'q֋דn��t�\їf��q$|&H���k��Y����4��lC�H���}yt�7�����%�f��X-9S/�������MfS�h��oC�fg,xi��軓�G�p��8=���Ȳre�7�`+R$|-���n�q�u{%M��1M�-;��	X�R���ؗ�W��;G]n�Zw-�u�J=cd�j��Y���e��ff����NE�%��;;��/L�tR?&w p��`>1��pV4�[�n`���i��\�m^ҷQ6u���Y�š��t��Vk��G. lsZ1�[�:gN �ǌ��Z�Zub�'�r��ˇr��XI����g�@�qr�6���Kif�u:�^����;,�A�xLm>I1��H�o�/�k{d�j�<hη4h1��t{)�X����}Z����M�$�I[1��n�ָX�Qj��p�*=����^��}ۗ�ΰ��d��=���;�_aԫ����Ǜ��(��]�	��uz��YQ2�.-(�����2���Z_3���WYt��Ʃ�#Y"A�������qqXhJG�/%��C�$r��n�e���GwVq\I#����I/Eh�V])���|P�i�x]Y8-cuxnd����CL�G
�F� �"T
�,#c�i�eՃc2�2���p,d�1�Y0�*;����6E�"*���lf|ѡ�EW0L1�Xk-�@YQ:�l�ۣ��J�Z�՛�f�8j8�eb�HF^\��nڈSa�I�H���
L�㰜>Hj<���HH��c��q��XN��-ѡ����R$KaO&J4PK��l��]Z"�}K�S�C]l�X�=n��2�w��-1SІ�g�C�xJ7'���6{�~����HJly�P�D'n��l����TE�TE�0'w��Q�Zm�CZ��7LjG`�����&��HVV��'�T,9k���4V��/Z�a�'t�V��נ'@U���M�
����Y������RE�đ�ͽ�Uh`Xl0B�x' 1�J22��2�]�L2a-�
,�EX	�G1���)[j.v���)�^�@�ʈ���F��cÙ�pVJ���S���r�(��:ډY��ݻc,��@ʔإQ()��$��c������ƂF�a!l?n�i_F��o����ȤPFDg�*-O1UX�,Q�"��FEq�0�j�AQ��T@F*�"0Q@X-E�Q�#��`�¥UdP�AV�J�ģ�EĪ��Tij,��T�(*�QAk(�hc1DA��q�A@Y���X�D�j�ET�*"k�.\pLR�"���b�(�kE�*�QD`�b�H� .&3(#X* �dQAb�Ƞ�"�bE"����aA�E#i(���`�#QeB�Ȉ6�X�����"�mV%a��TXEU#hJŅkXV
�a0g3���J_	{�ޜ�w{�˽׌3����ۍf��j"W���$�ڷ3��rb�gAp�NTE�����g_Z���< �Tڣ5ə�qj��<�M�
�$���3O�T��Fu��J���by;�"�C���?w쇉1
�Xl�7�0*
G|wW6s�i*N<t���N0+�����dx�Az���x/�K7�]Z��Ĭ:��ᔘ��u��g�~M$�:�Cwhz����湁�3�H���C�z�L~C������M�w7_��hV
�:�|(�'��%�y9w?UF����ᳵ٠��|�1'�}� qȟ�u{�}f�
͛��>�$��?Z������Ă�$���R���|���?!�8g04�d�b�xwX�<k%eN���&�4���g�f��]��|�m�������z�ͤĕ��d���#߷�R,����	�i��q>�ֿ�=��I8�z��1������h��MjAg�߰7�'����.h�|����3�}�m�RYqM}Ͼ�����݁���t�<B�+Y5<�;���1�C+�Ă�
�L��1 �C^�i�ʑd��q�I_Sl��������x}d�N�_q�q'�A �:��ë��}�<i]����zx�&���Y�%J����9�Lt���;�L=OP6wX��R���;�r��>f!�<M$�7��T?'�1���4��1�jE�3z�D�".�D�3G��&>kv��[���?v�m+6�Ol���$���u�۫`,�w��E�ӏ�s�f�*������L��
�}܂�Փ����u�(,+Rx�H,��u$���I��W9S�kf���X~����~���i+��:}I���� ��=�L5���ORbR�����o��La�����C�E����<�"��]s��I�����ϻ�R�����3�4��^2s?W������g���}�s+�ᆏ��#��]>��*Agϛ���g��MZ�i<z��H/��S�Vj=̇Z��1�üͦ��������1 �|�ܞ���*E��o>�wﳟmJ� Q�����@D4�w3�]`m'��ə}`T�n�{q�Vq��a��4�l��f�|���~H-a����
J���]<	�8�Hr��9P���1�^N�y�Q�����ξ���r�Dޢ�����������sv��8�|�:*K��V�0�6WX�9����;�kbaoҦ��!RayM��iu;��.���.ӵ)��؟sİhm�'Qn��Z�ՠ4�ޘ9_"�-�/��U  ؚ�H��]�?���#��}������|�2l<�M?0��5'�wZ���?!S��g̛@�V�����$�~<��i�~��ʑN�|���=�+4�P�l�>M���c����~���\��\�>���̏2�{���O��?2��g��<C���j�a�cs�f�2i1�<C9@��N& ��k!��ɹ�4�^��%�d�c�8����!���u>��~�7{���]�|3y.�߼*�G� }��L�������rO���8�����I�+�s���Aa��}��H/�8ɞ�1�i�M?0I�I���!�H�+S�ذg+��IU�?�XcJ3{Om�S�{��8�!�=f&$�T���N��1 ����a��*E���1�����wy�P��xo��$��L�̙��c�Ԉ��.$�;���}�"�1�l��}�������z�w��Ak��2��� ��]�4��!Xq<N:H,�3{��T�����hq8�0���5���T;�1��I�ӷ�d�%g�;���g�d${���Z��1�ە7{���|���y�0�+��

E�z��_��Y*�p:���c����8�2���ۧ�Ag̩����i�|�2T�O�>�w���'c�>�@�%{��+ѷ���R���{�$|�ֹ��9�]<H�1�9i����L@�޸i���ge�	PĊ���rO2��I�Y�L�'\g���8�>d���ޙI8�z��O�
@$P�
:}�,���[�(!��B�:vv�Hb��5��#�Fǽ'�>`}dR���ï�� �I��i����a`V���Os�蘛H/P�,�!����=C����!ԕ���L@�T<GyS���ͬ�/��$�#��M�|}�G�A��M$X������z�R�����Aj5�m'Si��ﷀm%a}�i���!�o�M�bT��XϾ#�@�,�'ʝ�ٝ�DnN}_,���~�vE�8�;e{?Xb������i㌘�į��XW�f�9��m�a^�9� �P�Ϻf��
��]�ܟ��y�'���k�&�u�{�%O���@'�օ`�]u*���fw>]c0&��������3N��oU�]Hw>�h��K���ʮ�@���	ޮ��V5�Z<�PPv+|5n��{b6�.	L�;�|�.W�2�J��Ŷ�:)��.���{yZe�8�^i�OA�dPF{;�Ӎ����շRK�]������.k�I�G���#�����'��1��Xc�����)�'S>�]0�5����i�z�|Φ2VW���9�<I�"����tzɿ()|���'�3�{��{�ܟ����ʿ��
Kz����4���i����~䞦�X�xL2W�Y7��g/l�����AxȥMKCOY��>��v?�S�T\q�ֳ�z�xp&$���ߥ��ڬ�0�IGU?x�$
 I����0Ǭ�l3�i�Z��+����M�q*��������<�m��y��AH�I�n'���J�5��|H-Iyez���i!��k߿c��>@��O�	*_Y�@$D����>|H,�xg0��@��g?s�<~g�1�3Ф+��c53��E�Ƥ޼��m��9��4ì7��|�Èi�a_m�=���O��h�v��{�[5~�:p�>�=��͐8��J�yI���� <�`3l��Af�;���i=LHx^9?$����bgh���c٬�������]��7��4�L��Lb����D3gӖ6�v���ѕF~ǰ�6�Y_߬I�T�~�1�>d�)�� �u'�3��;���S��2W�
��=��6�ɤ��O?s$\d����g��VOƯɴ����{Ns����{��۶bA&�WS�+yCN�:�ϙ���6������L�C��rM<C�1��?M�L�=d���m}N2b�_Y���0*;��4ə�P�i��p��i����K����@$����{��Y�J�ְ�Ǐ��y�i����O?Y������봂�xP�4��V<�CMI�b���>�$�>C!����B|���c쾈*+~�w����J���D���{iĬ1�~t�нͤ��a^xkF�()0ܻ݇H,�4�C�>L퓉�����e4ì�����$��8�����*J�{��%��+�?����:�7:�ߋ�:Cd�����!�Az���o�>O�/�*��+
�<I��d��2VW�ٮa6��R[A~N�}�P8���'�����T�9�|�G�Af<=���b��\�r���џc��v��4w]�e2���ϻ3���ɨ�mt���f���&ƾ-;!y(#������֧�����A�Y�Ǫg�;��ˁ����..�Y���[2�=��s{�;��܇V�]ӵI����g��]ķ��2�z%a��gv���|�٥�4�3y�@Q3{r��-�陎�A��� �k���p��b3w:����`�������L���1H?}���'����e �!Yĩ��`f2_�6w�?'��ý�[��bA�ﺨ��B�rg�%t����3�@�P?~�x�`�P���Y	:|Wà�s���_�����߾t�Ʀ���'�L@��k��>Iyz����!Y�&e���i��h��Af�<9���N;t�Z�>�����u<M0��@%�>@�$xྫྷ#Z��}qj���É��1/�D
>� � ��zJ#�f!�<�P�Az��l�q��:��Xz��o1B���=M��
��x�J���ͽ��Ss��l3�Ă�O'7���>�XI��{�^woK��2�v�#23mA���}�Q���ޡ�MCT�0�$ѯ2@�8�v�M3G�4�I�k�2i���d����<�Y��i�_��^zb���ߟ�|�_L��d��ɦ���4�̕����O�
�OY�H�v��l�A!P��?ag̗�n}CmM��n}�C[���b��?0G��r'J�`�M���u����~���� ���gg�~CH*M��V
z���3�����c�� u*5�	��~d�O7x�Cԗ�����N�_X�O�hH,SA~�#��|@qu~�e�*�g7��g���m&��H>}�`i���P�9l��I߻���C� y=�eC�%^��>f!�?a���<�ぶu��8ԟ���������i�X �Dw�T0�9�U}o�}y=/P�߄�M!R���wl!�;��?8�S�{��&��L������x���4��]�f2i���~���Ğ����rM2�������O���l�? I�%c'�Rq_U�om����_{�O|¡�X~t�YY��<hm�Y*k�}׏��LIP��T1��d��Nw	�ϐ�����>d�O{�?2i��O�f�c��}C�v|,�t��#W���`����Z����/G�I������y�I���|�$��z��'_�����]��8Ρ�J�5I�����4$�=C�w<0+֧��Rm�|Ɍ<��B~[=�MA-i��.���_�g���Uz�/rw	#�������@a�W��s֠�����j��L�R�,�0�t^��N�������{� y������%׊(���$̳���w�EĖ��� dS��p��"L���'s1���/�RJ6�l&]rEmR�(8v��$�|G���P�>�������g��76�'��ǝ@�ꃺ(��DAJJY�PZ{jTZr���:V(K��T���S�5�GX!��&C��J��`���<5	}�n��X�C�ڕ���
�E�$�r�/'-��p�U�})q[�D�H�bh�
������j.�W��0)a�\l��3����y]�iW��y�p%�g6(Dj��d��w`.��]Ƙ�N��z99o��n8�3"�U�2���'�ԡF�T�j#�d��g�`���{A��%�q�6�D�#�#{�/|mr8��J���_In��A0|�A}~f6�NU*����#װHV�v�l㮾�-�"�D�˼V��k,�j���Y&@�or�# 2 �
�+k�R������x����z�g9�;s���|�F���ٮ�M/&�J|OdT�{Hf�|l]�:υx���#��yg
o��/��}B� N#�Uص���}���Ckw):�2�ϣ�B��0o	�1h�Y�'�t���=E��%�n�w�D1����7�2=~���y���j�N���i��J����`�K�ݔ;kR�29��va���I�u�܎��{���j�F﹑-VoE�����s��z�]U$W��s~N�������~������2d���Sý�^GxF�j0�F�#}���tӆlr��9�y���m��޿V�{�ukfd�%��ozx�`�}GmK��!���7l B$��gX�T4�)�n0�'j�?�=��·}�q�+r$:�|��^�L�ɝ"���d"s��"��`���9j�q%k�<6+v��c�/-��#�}��|sa�(�1����z�`2G�+2P3%���������ƪ�(���]q��5���1��޵)��k>)0ҥ�</�w�՞zN�x�^���n�[o�1)���Ӕu��D_�(���qu
s��T���t��,��������g5t~:�q ��c&C8[��b
���%PY��(����>v��V>�<f��]Rs�%����������X6jC=~rP��{y�Q���a���N)B;P���	��9�jF�n�Gw� ��Wư]�H��U�m�tB��ՈM�9v+�Ĭ�\�3�d��k�R��m%�K��\Yu{�[�`�ӷ3�=r�@�eY�r��ZǽzrSo6����#�V=��*f���k����t�l�31�3%p�[���$�s��4t�,ȅ~Q�#7��V�oscX]Ʒl|�2I���$�gʄmǦT��ati�3D���<C��݋��Yy��_\�4X��=
p7:<{b��Вz+�a����$��W�g��k�3 ��w�r4�﫱�6{a���#���q'��;�od�k��A]eAFi��r�3mꉬ�w_-<���0Gdi���gU�3e���$�o�g�^�+	<�#]5ME��k6�j�����v�嘈bzw X���˸��'Ehv�K����N�����'U�JK'v��drj7�M�F�)��,ߩmi����j��cF����x�U�������yC?+J�;�Vf�D��V�G� N��C7o��k�z�,g*��������";540o��ƺ?6_t�f�N�I~�����#'91���9��/�D���^��@`���Ъ�|�7h��U=��[i�J0Tq�gb�A]g���UvS��p���LoFa*ڮ���)]9�l���]�7>u��1��q�s��u�o��h�]�kG��z��� N\�'�}M\�6��5������-�,|���뱨��l)�gP�#1�}����L�sz�������0(eE�J��p�X�^N�SgX��D	���jj᭬�kږW�{�W:w��U���޴f�g��:=뚨�A���U�����ʥ�ǥ�v��!�݁�q,��e.RD��$7	�{!S�v畍Q�F��WiV���JZ���L}�j��E:��*�D��g:2u�w��fXN�踑�n^5+k����x8x�W��9?�� :RUE�ǀtwKV2����H�n��7���.���[o�r:I��錊n݇��vY�JE��k�
�����+����\6���/|F�Q�wt�ZJ�'t�#:'5�YgNHwkX	�*�oH��F�v�D�iY8T�Vo	�2�oL�;�abĞ����±*���؎N@T��?+�U ��8�0#"������۹�V��~�]c�����F)�q'S�ߡ�!N��d�(2t��.\��f�t߾�Ջ�h��Y�$+����9��I:%�5�����&\q�};�Tb
�*A�GF��0��ϗ����*����a�=�׊��ȋҩw;P��F����L��~n�߇����{U���~Z#ʯp3.�E�7���?\�]���V�3��k�R9��P������c�<ù�WEV*<
��uy;�N�G��%ÇwF�O���x�M��p��*�q����{Ks{�V +c&�-Q�ٸ;��Y�6�,w<����\�O| *w9-�Z�{!y�|�v���i
[��Y�	���E䅀e�d+�rL�f\,J�s�=ٜ�\���'�O�oK�g\˘կ�B�V��o�zo�b��]����yg^���݌^�]����qA6�i�=��	����jGǧ�3�rc�ccrp�ʖ�R�r6�۰"*���C۷��c�^79#n�kz.�L�q'D�U(�x����ӓ���Ry����i3�ZC7��V	:>��Mt�G9a��N�=��q`7)Ƒqq.�_`��c{&�����c�����de{�u�=��y��֛��$�|��r���֦��<�&3yn�{��<�^�j�*�?F���XnY�W�xڕ	ØxB�O�S���Ck��)�gs��v-��sF`FgX���=�K���i�k{l��"�H���J,C���'4�����V쬌V{�s>��;��.�Zԡ}A��!PR�tZfx����鹄}�9��)KƯq��7�xڮz� ��@�ɞ*��_Fd�Un�W+��e��C�"���Cnn���{�)�(q2��wvV�K�x˱l
o.���f����,�F{�3p#�����qkD)~9�iݻ���d��Z'�ͱ�sx
���U�?-t��������9N��{��N�1oc4\x$�\G�z-N�v%�}�S�'L��> �u�r��O�v�/�|n`�W2pR�gpr�HDO�����{�ݸ���ʠ�
��}yX�#�(Z4��m�<�� �f��ϼ"��\wϫ#�	j���L�����E&�xO`7�<}ׂ�S̓���KNxvu[མ���
���̉���W7n�?�/f��t'"9�W�q�h�#68�;5���ѱ���EK��j�#dkJm��	��Vxs\��ب��gM{2�W躆h.���s����V�Y��G/�>�K�;���R݃�mv#1�2��;R���p��U�0s��i���e���<��~c�Vpa���=�`��'��@���M��J�"�@���23�hi�s�P��5"G{v��с>h����v�k*N�tN�(�f�H�5Ŕ�� ��Հ�3�����~;����g?KRV[>��6(7�6��sa�&:Y�VO\,2x�!�,�j�z�M��l�o�+k��	�(�X�C�W@�n��N�tU�RO�q���%�<�C�i���(����U�o��Y��F�Mxs�bn���;Z����z���O^ю����Dt��p�*}ƥ�ՅȞBh�e�K����5	�$�����c�<cљB񋵚��`�Y�p� 7�e���RU+��׆wL��Aèf>7�C�iw��s�ܦ�*HWfjLK�C���i	��{j.�i��,8@b.�2�^�K�FꞞ��q�v�)�I�,�G�����u�[v;Y�R�7���bv�Z�Y��5i�3�V�ۨ����R��Y��G^�gb����'0�:��)"��P�\�ѕ&g#sD�ո�|_}��3%�j�h73&Vpb^����{�'8�M�R�hH\C�=���⣁lj��K�>�ϲ��4���:��{/;5M�T��؄v0����æ`����n���У�-�G1�S���x����n:�#�H�Q�YO5*c(�S��X�g�$�\�ʌ����2!�5ī��x��-W{�AM�i�(b�b��Y�J�����ٛ>U���\[���f�o)5�T/���J�mU��f5�|+`[�-���q��8?&��^Gzj(�6��|�iv���Uֺ�D��t1@��� m�6�{*ܱ�Bun|a���S�I�FQ�*�woMb�� ���${�7�x�<3K�����`������(�w^w��3Z�fÍ�zx����S�����
���l�#����;��'�xc�����;�I�����\�������n����ټl�UM��@�;�w*�0��'�0�* .b  j�e<%G�s(ѻ�%]�,L*u����mT�p^P� ���1[�k�U5��ٺi��ܳ#^#g�ǡ��C��)�d����BQ�ѣY�T���b�)ѠT����H�*��M�8�4�&M۪��^kA�Q,�����1���h(ڶگ�N謘�֜�6e����2�ʐ�c!,RX9MP&��v��7���v�C*�V�h˻ʻ�a�	��%��%���@gW1P���E���R!�j���nY�3��ȷ^j:����Ij��Q5*Z9+`FM;E�P���?H�5�@JW��ihT�F�Od��]\���r�SY��Y�QF�P�D�K]���)�.:��^0�lpy�q��O��/�b��X���|�5�4�I��V�c#%xh�R��dXd��'\�BN�s`�C	wgI�Mjض<���m�r�8.������Á�x�v�9L� E�J&&fF ��)l7��Y�����s_�~��AbȰ,������XQ$Qch,X �kBԫ
V�AIKV
�+*T�mFTR���Q��T[j�eVT�ed�"�5"5��%B�QDb�dR�(-J�j\LI+*(��ŒT���Z�QXJ�+Q�Y �[h�E%`��V��-�X
��E�R(Q%`�1Y�ذ����m(�AA�������ill��1�֩R�)����[J�2
��4e��-�.PZ0�YR��b Ṭ��eV1��l���.f"LQ�F�-`���%���q�aUU��8e��j��aJՕ��¤�iU
�E��`����-*UmV(�"Cbbm(����-+Re��[P���&x`��L o�3����e&��ۭœ�	v�Ĵ��w�4]VَaA�A��Z�T̠��62�S���( �>;��ױ�*����9ka3�SČK&�Y�]��;���9�|��S{P����T�\IH(�w��)t؈�v*_:��nF ��{�j:�7'��gA�9
��]��j�Ȭ~:�Ѝ�6,J}^xWn-����k�ޜ<M�m�5�eg������~=�^�{�L*Afzes���7��5��v�il����v���m�2,�CB�[q"V���0&�#����]��O�]fY�N�H�vv�iT��WQe��`ŵ[0����S���i��Jp�zϵ�>崂a�)����[OM} �ʈ�GÃ��5"6.�~��h�Ս�P�b��+��ձ����,`nܩt��M�0|y��G[�yLr՝Q�ֿU��	��=��Y�O�Wه^��5�l����~�e}��Đ*��3�W�\�f)�.��
����{����d�nrCx=��X6�k͸:f�|&nȨ�#Y��s��e�d�#�%8B��&�_)t-�7j+�z����[$ɒg�x̍�;ID�%� ��ݫ9m�
��ٙ�4*(S#wQVOsY��b�결�S,��|9�1��g��I)]�VgH�:�{�xx�en7M�J)U�}�(X5��P�I�T&ޫ�d�N!��a��P�k�G�]���]䣁&����	�n�1rVqh�����x��̉Nr1un��c�J1�oX�������:���N��߬N��e��׼�db�۵r{�9����y�>�Y�_f<�v�����Í�ն���`��x�i��E����7i�ݔޕ��h��<2��ᩝ��ⓦo6�����*n#����g9�[��c�\�g�h��P�F�Ou>�C����N��tt(�Z
�}I��
]"]��6��hc�n��f�J
{���s4�ݷ�$'M���)퐦�(�g��N�뎽S3f'AMd�uC]���-�G�R��K�#�����H��MBX��g{R�����P�Ecz
�=a���
��e����8����>93Jh�&n{�#s' k�3E
[�;�����Y�Z�q�&z��,h`NN�����b�xe�E'�O%n��TƔ���u��g�+ |+h��v,�ݑ7��
�u8���菕Tn�׽ݽ�t�b�fW8�5����c�4�}h����4�C,�8�^����9�u��̕&.Q��{aa<¢_�6�K�����_:\�r�{�͞��MǛ��g���Y{��۶�َٯ�%,���`W:˞[J�Qmń�𷁜M�Nҳ�P��CRy�iP�q"_d�ŏB��
��*�I�ǌnT�9����Y�{�=�2��=7�m,�Q̠ܬXJ����C�ʭtcܝ��n��9�j��<,	�ʆ�n���+޼"?m���hW����O�Oz�b�K
�ח,<�࡮��k}p�X&ި:dsp����-py���B7�la+ɱ8������q�1�E'��;�̻g9�v6�s������X�=C�CX���^x����[@����z�yK{�Q7���r�
�ve��㓯gJ�S�A�}��>b\����ŏz_M/� �T|�q�o�h���}��� ��z�|��S֣�z�''K�c>���!����q�P{c�+�MO�7�K�@C��)|��6P��VṞ�>��O�9\L�K*!Sf']_���[�m�x���d�W$�k�éPb[��X3�h�rĈ�o4p����v�/��zӮ|q&�L�W��u�n�yޅ|��BMC� ���ȩ�c+���vT���X�VJV��C�P]؃��$7M���a.�|ء&җ�P���f�ik��y�?���-S��7�n��xq�L_W�������T��:�����m^���p�^�p�U�vH�N7V��`zz�8Nh�J/���_M�2�P�]
�Ǒ͈Z�졁\�k�^��1�2���SU��Z�[ݕP#�Q^U0�%u��v�d�R{*���ڥ��+{oe�ޭ�OVV�h=�6$&,O;r+�/��3'�S���
u���#�n����8UK�`��a�L>�N�f������z0TD�K5���k�}��&'�v��H�N�\��aW��ڰ�mc"�k�H��E�꫋If+0�ޡl��ݛ�Z}�t7|��y�H��j��y�� ��gG�β5�"ӷ�aջ��D�a?v�	�e�`�7���e�w�y�������i��$YE�a�H*Qe�ݩ���6o�ucsN%�i�a�N�b��tX����3^�o�ݢ{4�m�wX3c�)�B[{�����<ngw�>�ɿ�:��E�S��CB��\��ݝ��i���ٲ�$U+�f��,���7K��*�����}aX]Ww
+i3{�S��l�� ��y�yE\[���?16/zf�W=��oW��+{M���\���F.o1�E�����=��G��ݔ�c8�����h�4-�uSA�9���{�����uJ
�1S}�a�h�u�ݮ�3%�#8P�Y[���b�� �o�5~��Ut�>̳��,�{˥]E���a��F�5�ץ>���;���u{��g)v��:#PI(����Ci���N�x������z7�/�MγF�WM7�a�Z�|��]|�M�^�Xo��@W��j�p�Q�%k� ���t��lli��Iҭ�t�f�&�V[=!4Ӝ�r+�%u˟-��d#�:b�fE"8�8��v,���.��(��WM;���9ﳋ�/rP�*��Dt��k�OSޱ��C^�X)�r�<���jZ����ňq[�
�b98�UQ������v�������Mu�Ah�Uڄ~ۑ�ָ�x��b�\M�+�k�A��fd�3�!砂k���/=�i��SbSx)m=�/��[Q��ah�gyf�������3qs��s0�c�䫤���iGm�����x'3(J�4��	�m.؇�~���hш�C߫0=$��op�o%B�h���{u�f-���L����-@��$t�[�A����?yY���V��WR\7˦�[��^�m�)��g8����g�S+r�׾>o�?g�O����[A<����*�ŧCjؑ�/Oe+�"���3�ʓ�;~����{�l��ʊ�Do���xߤ��+��^Kr��q�>�hr�l)�\��yj��g7�$[#3�ȣ��ﻌ��ս~��QyQ{��e�ۯuFN�9mCJ��C���}�)��Pm2��\�>�B�tIH-�1�TRoU��:'kӤҾ-�D��d�欹d��u.���Y8��k�rcJ��ƙ�{V�v{qT���gȩʺ���>��-=%��o�O#yl6a�um�f.���f���W<��4��r����u���eKK������u�O$���.6����i��_.�QO�}U����H��'���r:�t(��T#DI=�u.�K��F���}���O���a�(�c�^�����r����`*6�Jɠw����k���}��Ӻ�Пu��7=;p�@N\ׇa�8y��J��M����.��j�6ά�x�[�X�U�����U*}ϩ���Z[c�ln�2�vZ��=��J�h��v�׋yC��岑���=�[�4�Qbgokw9峰�Eu��`pW`=J1�K�ͥ��T�TZ:x�Y+��o	���֤9J�ZÛ�9�>��}@�̗Iw�΂�_{�[�����l��;g5�a�Ln�#7��{��9�����f8뼕�TY��8�#Ji�74a>���/v�����"�kl���^�ٽ��U�gl,�ZاܹUS�����꿢�Ϝ��}�xW��Ak��t�O7��M�hG�ǚ
�7�uoΗ��:d�[J�ؖP�����(a�OCE��<�����0{V���ь�LU{���͍E�v9����|FT��H�ٷY����M�]���7���x�zѷ�HV0r�qTz�wu�z��'E��S�L�_}���u\����[�����c���ޡ�+�W&�We�<^&Ԣ�a���؝�mE0�!����TZڍx�.ܗ^\ą<��7=���by��/g��T��U�[5�c��BV!fP0:��Z��=rҰ6t���OM:1iխv�R�3ͦ�pS|Rx���jW��+&�#xC���}�W���VZg_1�{-�m�l��ڻ��ڎ�v�I�q@��Fԉۈע�f���z�J�r���1�+$���]�Oa�{P]�1�oNKtݝ��V��f0����R���O���T-���S��s��� :�"Vs���kUו%4�U�K�"9��ʽ �}70�/��{^.���]�[Q�!��u����R�Vu8u`�9�r��}z0+��].�k@l�<���N]8��ٛ�e��{]�*�ȭ��x��s�%vN'���$�-~��#żF�T�y��[�L���*qo�S1��Ԗ��o,u+Zn�Y|Xr�v8��(�-OV�*�UYFw����U�3���]rã�wz(�a˚�Iin�`�&�j���X�B�l���:���}n8+I�rs��z]�S�Cjz���Ճ�gN=������}���L=��Ą��nE{��ۣڒ�oN5�վ�:y��Þ�<�޾���a�I�����l�.�����H���Y���Km^�Ӕ^�#Z'��1i��{�l��	���ELn�G��v�e��7T��G/��`Bf<��L�B:[�S�\8͸��+�ML�j��E=y�b���~�;��Nr�!����A+��N�УR�Ӽ�TOf����V��W�{���dz�Z�\�w�u.x�hm.�ۜ}{Q��.H�oK�
�I����F������O"��qq�&imҝ�b�S��%+���ѝ��#7��>���X��	�mxZPUz�2o[��}������iW�IEO��U�O/�}�)���W�����b*�\�z�SO�+�2o��[/�����؂�A�ߛ�wp��{��{�H���u�;Y�ڜ��e��}�����a���$[�M��V�s�}�v!*�h�7'6e���v�6j	�|�_]�J���Đ�Z��k��F�c!|Wn02;��$؉tCf�=ٜ����n�*j��V���r��E�0��l��}O3�}OEu^m����KKaP�i!^�MX�]��&�gB�b;��sm[oy��'q�9>�+/!�XBT�U#��M��s4�Q�6L5$bñ��ifGFڬq��;�t���-�{S�s��+����Zlz�
~0����[��9%���zSBC��J�ȡ�WQe�E,}�$uV�0Q�X�K�\��ɡ��ߩ�2�ҰS�E�7���r!L��[���7e����HY�1!�9f��9��'���Z���wp��6�c"eܷ-�ۢZ�R��S�;n�3!c�ń����\��ouD�/}�^*/�v��l~���1�U����CF��]W;X�K�t6C힡F�fn���L����S�;S�ujF�s(C
A�QoWVb7��>Ob��?s&p<gTޭ����v�c���ȬyA<���a�Q�^ҍ���B]:���mT=��kd�/�3!���n)כ=�B1ntWo��,�n!��=xP4<b��i�'��F5�g���W�K��r�~�t����,?3���ި�2k]��&����7�"_�چ����@�{���˅��L�'V,*��l��+�C�ޮ��S�u$��W]��.�k�#먩԰I���Y.sSn�j���,̒���7����('��x �<���o��˖�O��\;f<���F��2�Źe�!� 7
�E�fmm��ޓ��"�&��:��%gӜ��_���%v��z�C7}��V�%h�����=/��}�����/�N��K��g�C�Ѭ�����yh�ꇪ:<=d8��I�[qDլ�5��mp�����Ҿ[��9�7$�y��קh��	b�K�+��&&T�VDdh7~ېQ�t����l�u�oK��uqC:b�ǠAuFޝ���Z�,���{y;.�C05Y,@���u�w����4�/EgA	N<�8�0�<���OC��r(��V�}n(��l��"/����9b�I�yϓ�T�Q�`gvs�zH��:c����dէDJ.�<(�<3���;��+����r�����7����=j�gW��T�q�y��"YCݪHb�lfu&��7퇳)��׆F�1Y3��nqL������U�ݬ)S5�+��U�l�W>\�L|� �n�����D�hэ`z�}�&���-��s�;\���9<:��3��ep�D*Pa/�,R ��s;�=ڃ,�w��u]w�N�F.w���|�>8��S�sMN�#��&;��y����Ւ?�ߚA�<�D/j���K}�L��T�m6)�E�2tԟ"ĭ��}˶��`�;�*1��̢
$���2��9vJ��AǴC���5��ݽ��`�l2�gE��l�f�a�V���Jt/�Ib�2��;���᲌��8��͌T�Qd��O��\���0[�U�k�E�
�r6�Ҷ���y+|���@��se�`�xsJ6�yJЄͶ����a�#d���(Vֆ;~k.K����[{��PC�R����+LEQ�Ik��f�TJ�2/�����ٟ5�B/خ�n̖��XX�hq�%�nF-� �(��F�\�Nᳯ{�цwV&�f;\�v�n1V�'���l��opjv^�1n�(K\����Yd��V5*[ΥTl�!3jC��N��ʖ��#����9��o�sK���1 5���uz�<��K���ט;=:0�Xe��m�ۨ_P����b-g��
w���9lR���c��ˡX��6�n���j��_m#��Pƙ��"�/��خ��p��� =�S{%G�ݛ���H��;�����V����t���W�P��}����~���u�F��ꑀ6&����̜����Ԟ��1����AZ�Ua�t��2p��L�꾫Yݙ�Pw�����J[L�"�g^�<���ɌtŃ3,��=�iƥ�.W���ߙ?`LE ��G-V��j[Z#lV5!m(���Z��`��U"�UYPY�Z��aXcD���d�Pʢ��T��A¢[`�Z�#j���eJ�+F**�RԩV�4J�R(2�V�����TJ��UP0�Uk-h�Qk-����P�C�*��m�*jԊKh�-�ڔ�j���meT��3PYk�d���Ȉ��+n4V�[Z
(����J֥���TJ�X6�akeU��kFڈURҤm��d*TV�EŶT*6ܳW(��ԩE*""Ҷ(6�-�B�-YTEmZ�T�F*�73�B��VQ�X�Z��h���d��DeETTm����0Tm+(���Z��b�QV�Ih���Ƶ.c�>�N G�}=�R�*�P>�vB�]ӵN�&w�rJ������J%����]�e���e�R,��@$n��;�lINht$v��n.�}xj(��j|�2m�QSY������&l}V:}�%�ƫ�*�M@����=qdg^������']��fܽ�ѱ<�^�[�~̣)�ߞ��S9y�ܞQ���\�Jg�g�Wzꁼjs�L睱�J�\�`w�5������jQ������&ڥu�8<],1�^�|�c��ʆE������	i)���|Vۤ���_i��~kaP�}R@�و�/��O����3$9ΜΩo�n�[��ΰ�����nz�6;!u�P~�i!S���Õ���5�'���.�Sޝz�n�Ӓ�7g��,!*�
����qc2��;���Fz���٧=Um�I�N�	�7|Rzs^;t-�d4�Jl�f���m_U�(=OѾ�]���	�4�Z�u��������_nU��DU
δkr_V��"�)��R�)��΄h�[��
���>��4�Z%�3`tk�z�W$�T�w�OJy��:�E��{]tU�wfO���67�E�F�:"��C�j�:7ST��ȉ�*���t�2ΣC
5���-��aR$��7aҮ��\�����kNs]�rs���a������:ŉ۞�/����e=�
�OgVZv��32�ӻ��ݙ}''��9�#7��+�#X=��P�r'3�FF4v��><���Y����}�}�+t�������D��K��f���K;|�1��wY9YM�Zv!�����E'��b\��A�j�Gt�P�B�#�����v�R�A�B=��t+y:�p�'A5���4r�47���
C�����C�m�ۇ����v�X�0��BV�p���*�j�Ӷ��i�L�16�!�G%�&з�uV�4ztn��k�U�����kz �}^��E��;L4�l��
�ke�@B��51�Q��-�^d��^W��}z�}�('���&��|��B��8����W1+�V��[�축?Dm���t�w>�;����޷M��0ʚ��|u��[��f�n�a�=]h��L	�������tY���X�������8��=��z8���u�0�Jb��'t�y��}��oe�R?Q/H%*]+���yM(��/z�@�n_��m����t���R1_w���cNY=���[Ԙ��Y���VR�O�P��V����t���^���Ó�\�m�$����Wp�ͭƑټ��T��ylh�i��+��
u��7���ޢ�74*v����8��M�PU0�s-Q�U�R%k�/��N2���J�����/��ee�+l�N,6�E��
�ȡ�R��݉ۉ��q����.��ӂ��Wθ�Z8ZL=��b[$s�"�_W���o<v8�����в:�zt1��+-YL_nPŎk^OIS�0�cyD�kgG�g��~����__��ImcQ���.�}7}�Dw��~o~�gtvs��=��ƒ��1,-�cp�*o�ee�=��C���>񃳽�Ɩ/��:�M̸mde�ٙ۾�sznw���!���F7u��bY;�b��M�؅����(��߻�6G��֧n\t?vM�&nh�|D�S��Qj������ +�q�9��)pK��z��Sל�ʼ7�n��4#���7,����1�7�F�l��	򽸍=��$u���֗,�l�u0*�/";jvh�2�:鼶�N����u5m�y\�m���>��R�Pa��m<�y�����&��;��|����VMV��+�1��ڹ=��s���7��i�穽)<{�����a���޵0�o����D��Ts�p��j�A;�����)C��7w�yb���v�j��;s�9���АU*A�d	|���78��A��t�@��ծ���Sj:Ӱ�m,S����HT�j�2�W�qP,F\����^�W�����/�<7��s����%@��Q���ҹ�*��ge�yi5Ks���mz���qV��t悙S^ΧՃ�Df�nw6K���^�N�-�Ԫse�v��[KO,e��Z�U0˂��|0nhWӋq�i%�뉔�k+��+�s.ym+�L=�6%7���� ���T����Y�m(W}#��~:)Vȩ���⽂�G��w�Ӊ��㪼s\R+���ه}R�4ZQ/��:���ld˦ZJ*rl��=1пw��������`��OѬ�S�{۱#�����RN��''�j,�J�m+h��
���5�f�"��Hl��nB�]O�9�r��ܹܮ�b�i�J����b���d�Ӓ=Su��5�T�S���q�y+��]��3��E[��$}���<�o�R�����s~��������2@��Y�4p�����k�N��MMGUz���1�'��8c�4��yY�P�O�b�6�^�FV%��w�ю���B�۠�=�S�CW�[�A���{��ó��_v$�i�NKw4��1jr��:V7��zM�Q�~bOn�"e�G�^Ie���W�k*�����NN�Ar*usx��~l�9j��	k���c���K�}��-A]�V��Tk}Qʦ���Mp���WH̙Y��9"G��K�c~���T<{d.��P�P�¥�M|�V>K<g^`�rӞ�1�k��+�z>s��n|{!Wb�Z�r.e����Y�U��9�Ե�rR�:�VS�~m*�1���%�n�c�J�����F�P�m�}o��ܾT�7�c�#��ZMV��~ ��"��D��*Ma�f�3���f�Y�f3�Y���r;�6�6D��h=Z��ٖ^f&�o �˙����wU����/������y�ݙ�K�y�{��K�7JT��M��ښ_^����XS��G�r*��wUB}��󊷧$kǎ����5��̑�QztYZ�.�����U��;�V�����Fv�v�ӓqVDMb�i#�W,y̩���j6�D�ܛO'����ܶ�9������;���A.ͻ����R�`���/��&�cШ��ǈj5��v�8�>���B3c��p�s�*L�Ӷ�s2�)���G�6/�m�g?A8e�n<�
=��5�vSX�|���YO��߂��K��8\n�t�4q�.T��ݿk�1e�؅�l����5s��_F�(4���K-�X��Jkz�0u����d�Ob�jF��z��߱�A����6��Oܽ�v<ü�^��fk��hf��������W��s�CP��B�Jǲ���8��i[X⇷yt���/��;p��UZ=T�Ǻv佤���^w{�VW@�u�X��[wy�R�Z,<1�h��sڲ��9myZ�����fhl�뫛Y ����0�KW%A��ܩ��a�Z��v��t��ޙ�F�j�@E�x��½c�(�0�z�^R��2VdO]ަr>o67��Y.a�a��y�P�0��]�̿14�г+�:��N�`��7��b�孶�Cl��F<a;m=�M�Uׁ=�W��J�HƎ
)�\��gNb�ܡ����w��O-�)ihvWjq��(��g��zX�zq[-��jb3�L.K)t˹�w^ �o�NHn�R��Y��[��Q��J��c��d:5�Е����'uP���=���D=���3o9C��k�Cr���G*���l�^�)׷V�ή�qR���>|믵T����y��M�W�J�^�TU.$-v\LO�m]�dbu1I-�b�qm��ї5xVJ`�n,9�/[�]��+��q��T
pc��a�ɘR���
粡P�(&h�-��w�/���3�I���:�/k~/Mj|�������-�V���'�%H��L>��u������7=����8������|�WfX��h9E�p�V����*q�l�ȳ�$�X1�O���W���n��?��	�ƽc��r��f���	8#��qǻ��n��ٵ���|�ֶ�_;��i�����Az�o*�U���c���O+sI��fܶz��m��!�;�������Gۑ-�^g���.�k~u��]P�c>K����ֻ��9�}�"���B�1E�Z+'#�C�[��g�󭉞7��F>s��Щ�Ҷlb܊O#+��ܯF�df)s�~�9C�TM����y��f�J�Z���Wݴ�E�^O#v�1rr���)p��eeZc|g��wi��^/;K�eL�犸��lK�8y��6w��/�K����8�����z\=������D�s���8���i����$���uM^n^ �^�k�DԈ��u��5z���j�T�7�˙q��lw;oZ;W��{#�6���T#jA����Q��؂�ў=��]����s�T�utw�����[v�m+	p��Ԑ�<������m�۽�Z��*������9+[�۩Kx���ylo����k����q���pRb��כ���g�����{6_{�k�O�ν)�n�����[�Z����eE�C�#�04i5i��z4����HoV,� l��}|;i	1S�Ra��p�Э�#9�/�^���I�������ۈ��@fv���1=��Q����e�J����mӏ9,���h��@��<�=D��t�k���s}Z-c��Rev�'����}�p�(��l}3��Gk�O8���۹��T׳��u`Vw��N�c{�֫��gVV�][H*g�%/E��>U.D7�J����5��4�[<���c�-������sB�O 崬��Sc3������D���Z躚�[�+w(�l�H�%���e`��hb�45d����pS;��d o*t���7C3��[S^�z:�NfB�;�Xc�;Q|��5�e5غ��R7�w�F���_�߁�?>GuМ���R
����㞻�}��R1��N�l���o��w
�׽y�у�K�@e-�w��aO���U:��8b�BJ7�^��[W�#+��n�J�������U����H�ک�͹�օ-�C��7�c�����v��ڏRⓚs�.��9+����d=��(���]c�l)����{r�]�Mv��E�i)bBz}�{6�-w����;�Y�b���A��^y���	q!�*���o%JbT��t&�|�-j�/7�t���"���=������T+TuTƵu	E��3c�ұf��66�m^.���	�\��������aP����U*N�/����PI�,���8N��۲�ܖ��b��97�ҷ]�Z�(�¨�KM�T\�r|s�F�$2�d�m�01�ݵ�'��c���%���7(n��x9�KJ�LF�'5Ny󑘺�uT'�a�/�����{&gN��u���;�.��X�(�1AZ�.�	��G�'S�\�ڀrIUw7ۨ� ��`m�M:�#�hYր���J��S˥z�FI��IDWgv^bt��T�1�|zÌxS���ܺ���ӛ�K���u��ع��r3��af	�:N���T�LJ�w��T��v���[=�bI&��du9=u��\��3r�f���Q*}�0�&#k��s$k����x50�Z���Z�+ǘ����Rܮ����r����isRR����,L�r�̓�Q3�����P�}b�V��y/g�}�˅����@�K����3e1�nI��*)��0v\��J����9�h�T���rN�	a_b+�0�}Z�f.�c�>�e�sC��{��H,/s��g�AE൬�<�~����X�N5��圜��Jѩ���{��w�����tZO6����T���&�[y��%�4�{�օ����9Y\����'>y��k]�|��Р�����ofX��os��:V��N��Ơm���.�Ho.ISY��b�YavV[7��Z��(e���K��ȇ'�}fh[�ݙ�J�hL��M$��c]yg��F6���F����Cw����y���M�ʈ�I
X��a>��|�o�ˇq�Sj�2�x�.�B�2Q��L5Gv�m��U,dGq�M�Ϭ*v�\���:^|��S]vdGɏ�z�y:w��8jV�w@/��P��C��"�s���p�Ϧ�}�{�W�{ �x�����*[�t-�׏���}�yA�`C���Y�Y�2�<��I:�1���C�B����B��T̾��MJJ��p��;@��ڃY�j�u8"+�9�g_�V�|��2��`:.�w����ҐI׬ؾ图���o�eiV����1�%Y�[�oo@vN��Oԭ��؃>��I#ݠ���N�s`f�h܋�lBR���W��;9����V�<�Ns�XP���KR�*���qK�R�f��KECM2�ݻ���v(fZEq��RӭL7V��,/r����		��`քg�,*2$|�D1{t&�����,�I����u=�j,�h�����ّVr��f�����
F@�J%e�%CJL@���T�Jvu8q�HJ[�l���?j���!V�����2��ӹ�#Y4R�(p7o �vq�J�c��;��̢�e�C�R�<1V FHu��"��'"ɾ>�^�H'�ZŠz�Za�l}z��4Z�kXK��V<R��@J]���6�r��`�a^C!�7"�Ѥ��$��#4�u��X�1�1�0<�X�,�U��V��梲�A����(�&@bO�M+2�2�U�@��*�_�t�"�1�:x���4�����SW���Z_h��zmۋ�w�D>�5�c'"�j-9L\�x�j��ãڂR1<R0�<�wj:�t315I��:P�V�Ffe�XR�Jey3j���Y�RRͦ�i�ʖ^Jkdz�0ɬl���7v�� m���X�-�M��%DBT�e\bV�-E�%�`�X���[h�PV�XT���E��6�+P�Z�ilX�mF�*(�m-)R��E��E�[Z����F �mZ[����1kU�#)B�+EKJ�linf��R��Q�-�UX�QJ[DT�V�EF�
���V�Z��eK[AA��J6�ƪ��U�U�E�[J�m�ڍ��Z��Ң�(�Z6֡r�ţ+K����-�V�X�l��,E�(�@l�F�U*��Q�c�1b�-��`�ƨ��b�m�m��FcP\��,�X�++mZ���Fڪ�*QU"�V��QJ��r�b"����A����ZS-�ۊ⠢�[A��""£mh֢*���h"�1b �Z�X���т����j"��m��5iQb(�Xʵq*e�ZL�ZkcrQ�2�]�T2�-���9�=�����}a;ܴιn�{�K�M�o*�뽻���Z_{y���G)�o�5,�VѬ�d�Xbq�o�!,�8���S����ʄFv��z�'3�o���d�bghB�������q��5���=�9H}��{�6G��Z\r�3(�?k�_T|3b)�qy��k����������$�`K��qMmE�bv��ƴ?j�m��6�%���4��ޗ�����a>�#��BE]�uP�|�)�i��u���[������R1��i��7�+�O!���J��[���_Z}9���[�i*qb��;��!�'�K���=�ѝ�\C�S��q����W&c��d\0u;7��OsS�w<���:���u���+�@f����SV�z�wN�J������Hs!��I
��]�wQO���H�׷��vQ}Z9+��oU�����4A��o�vf&f�ح�7|3�Z�,�l����g:3Tp��3��̹��g[��1N�-,r�"�e`8�@�)$�wHNa�o{�:��sh|ŋ�E��vh]�s��W[R��f���Gu����	Xƀ�ta�����7]߄�o�w���2���wv�^�:��'G�m�}��W�94�R9��<�4\-t��rr*����)%z^�s�Y[+J��Û�ȡ�ݙ�=�9���:������ֹT0%nMb[�V��{��1�B�b�������*�=�o��������3�j���y#���l�I����(�R]�����n[Q�D�ه5���۟NfW�c��ČNGU:����&b��ɽ�b��2�+�6���`��������X��]�R���B���'�铳==������Ck��ߧ�ܠ!�����q�B��E���3��5�P��"�[(bw����t����	}���4�{�<����vVp�^��W�H�\�q^� ���ױ�-d%�<�c;Tۃն���f/�]N��"��ع��i���ס_c�Ng���^A�J�Y�^�Ю�}�Sr��K�����
�1s����[U�+N�l���b�F��L�76]Ĳ�X�,g� egu
G5`�;If�O'�����0�`��|��q��ռy��0A�[�(�*�n���X��seYnwa��/y�����w��G*�\�V�j	�;��N�W*T�S�v���`��@&���[R"0Ҹ�}�o���1�5i'оFO>n>U�}�{vǞ��vݞ�U��H-�g�!~�M6&���*�TU����}��v������Esѷ�%e����p�F�*x�nǲ.�)�N�zs�m͢���V=������ҩ�@s!����s]V{}~�a�N�<�e��h��S�K��_e`O�^��V
�zҗ�ݴ,J�Y*V_jJC'�x�kj.V�ױ=��\����T
a�9Yj©麠m�gkgZQۢ�l(�!���Ҭ��#�v���Z�C�J�ߎ�� TIM��+���v�ް�n����.��OGS�+�t����$lk���/۝�M��ĞUec���l����Y�����P;�7s��E���ݲ�i,]qN��.�m����9�Nޜ�s�+#��+&\��&Z��.6���ƔjK� ժ�s���#v�<�%��8��+��-`'�������¼�ۋ�y�S��������B�{�^�#׽h=�����X�㩬$�VT�G_K��d�m�9�'��|ݬR���x���c#�	�-���p���TN��sv���-�`NcwY9C؆:��(N��{�>�2�m�̣�&A�٧OkCs��B�
��`�t&���UN ��8��(l�{8�m�F-�ښ��w<�҉]*2{�؛G��F��6gO�?mT�|��œ�c���n�r�B��;�ѷ3yA�֨U1�I���\^���x��.�;�nc���2OO77��q��a[PWH*�>=�<�J�-���ƹN�O�_k��e�/v�oj�~;մ�p�Jq-��{�[��i3���N�V�M&2�P��G6�ٔ��I��s�`�Ųa����V���*�������as�3T�����ˉ��-��7J��զ�٬��ҥ��CQ��X�]z�v�Z��,�Tp�U�V6�^^���z��!�;k�֝2��Fy�wk�"�e͂xs~��gf�w[܏4l������XNۺ�9\)��O�5:M�k�H����@|��ŧ��y����D�����m��D�gw;͖���>d�7Lra��#�vv�˻\��:��9jT�q��A\���y�Gx����BnqO[W�=����g\��qaM�Mࠦ܊e��~���'3�e����Ĭ 6"��s�	�1+=o�W]܋����J��^I�˥���zlE>�ڲ���݁>�ἥ3����W}�W/����ճC�g1cX;|�h2�V�i7ݝj���f0Su죙^�ǆ1e��y籟����t�4�|�$��Ӹ8VMͪp�O��U鷪�'+؞�B�!\�@��jʬI$�9gba.���h{�+��#�s괻p↫7�Q�&�]D�ԧ��sS��j����[8>}�ߔK�=��zf�D��N>u����|	�T����ʧ$�=�'ݏ)�uoc��ͱޓ�S�O!�G%�bnd��μU+�i�\�v��-��\��-��M��7��W�i�:���-j3j���&�=�הt�j����Ws�]n/9s"YSH�Z���S7�"�`�YS�2��.%38[����9"�Y0f`��r�1�j����é��W�v��L͑���N��t��ܶ\=���ǧ�P)�M����h��۔��f+Ft}4��r�P*��l1���Ve�^�0&�hP��B�ߵ\�O,=/v�s����q���-�+� ��� �bOq�}U��~��W��dBoɑ�ܞ���J�1j��]ï,!*-^��z���Ѻ��sT�!�5��yկ*��S6��r�kmZ���|���)��`��jey�����f�nv��m9�ҹ�S�ReH�N()�"�����B6�-V<��L�(���jWu��r}����P���U��6$�EV�`صº�rl�{��O�ث�bLJ��o&���
������LN�1�Cv� ���������ku�
�5)�;j�3!=��X��A]�ɇ^��罷�s*4'=�y���K���d�@�?EJ������bHr�t�X��ɻ��y���܆��+j�&�`���V��9���+����O�8c�dtUL�:�,W�<��~���O�ݰ�Kޫe���=اo�u�-�5J�����1;�G�/Gu^(���*�z.�L�*�_`|]��j�wt�	4�`�>ᦆ�ٷu�滅]�l��N�.�Y6�E~��:��vU�ѯy
�X�u%�����Ǖ����K�����E'���`�W����qP��mI�]32�����%U-�T��;mj�X,��$�/�ޙ��߇��*>F%*�\�Z�u�$�)�K�/��[Gfjw���c5O�CRQ���e�t���BV�Sـ����;T��������x��U[�?zx6tSc�٬�w��B��y����q%Or��u��++�W>�ʭ��y@BH��V�][��\��u��oK�X�rj
�H*��	
���g�����^Tn�wcLmVk{�\%��?�������j���>�3�}�}�_!(�eKb����x�O�f�61��k��*�&��ؒsѶ!)/��ˁ�ʦ��wV4t@�bA��l�W���0���qOM�v�h*�7A����}Y�M�u�4��.;Ua]�0'#�UOx�����T��r������*����7['Q��0��HQ�V�����uϳ:��ذ��'�� ��q�ڗ�Y�g�0��j���f]̵�]twҏX� w���QG�on�mu�3ct^���U1�"'#'3B�=�4�m`X�d0U��ɥm�c�G<�7�����B�Mv9�]Oz�Hr����bNmJ�}M߽��F.����-9�D-���L�K�F�w�U���mr
��䮯ː�O�nMb{CB��c����ٚ�j�����j�kSa7cg�֡�]t�ʤ���Oc���D������}�kh��ՑU�֦o�����mJ�i<�ݵ������;�۔�V�1��=Y;T�{��a�?W��T�z�mW�랭
U�dUe*��h��\�T�[�l�0}��v�+��c��N��궯m�æh�X�:�u��yxA"����L�j�����1�p�x�Gr��>����Y��r<B�܇��}jp#�}T1U{.��'�$�5y���w�#I����]ݼ�����b��̠`r�����z�J�
���QZ����j��j����v��<}��IA�����w��:1����b�0�_w1�z��L�x{�M�z:�d.����UOdG:=��t���]ī�S!��4?h�s�)_;�ԡ��[��zv ��*k �w�0�[�0�Yj+�^���t���hk"ȓ��>m��}9u��׾�;��p�b����SxU4�:�V{�C��7�z�g��P��[-���g
�,��%�m+�ݕ�N�ڶ��������F��U�N���ぃmt�\�غ3纝���/�D�*��*��|�ͱ|l)��v祇Ҧ�V�t9h�Ⱡ��'��=�FO&K�ck8�Z�l��/E�x��Yn�uq"V��pQB3F�=�{=�EK<��羮�xE6�qM��WQ�m�TT�#��y��%�e#9/{6�uϺJ�q9�}~Sc9��j�MD��!CE)�x���m����ە<�qٌ��QZi�LF�9��0a�!UNf��	5��?G'@��Q�X�|1�� ��{�aR�s���b8�y��5��p�a�}�
��~9����9���:��Y�ER�nBǚ�lǂ�C���ʷ�Ӽ&�S@�c.�BsΕ^O|!'ʵ�h��^�%����hac�f�!�Ja$�/�����X����97�w*y��7��u�{a��WG�j�I��L���y]ה��]��dԂw,�z=˧ݳFC9��9����[G��
~A��j��k(k7П����A`}�	��t^���X��LC���6yA�K�=��do�ڡ;>Ë���N&'���:z���&��gÆo5/��7�:F�b��X�ԲUȷѵk!+��u'	�sw��o�ܞ�n�,*-���}�)��W�a=�y ڭ7b#�O72�=�� ����H�:��W*	�U�	���[��ۺ0�Oz:{��w5�rԎ���c#���0�6�!!B{��=7�{�ut�%-W
���o{/Y<c��p����7~=p�a	Qh3�IHhZ�S[�p�+槮�4�*������=���SX�۬���΢��O�L��§zv�]p�(�T�_P��;�u:{�*i���R9���\+V���\�<�7U�WzV�X���^3�<�V˷%��J�ȏ �&���h��3�
�=��EQn5ׇ9p�Z��WNu�c�6`ťq�϶�|�0�k"H���uPa���O/m�z�d�O5��I���JVr�edY[����<��,��u��cB}EE8�݂�nq�w�a	{M�0W��r�l=Q�.\F��r��_,����*M�֚ZA��tY��^`�G>���哵lm�n
j�ok��ESi�����z�d|a�+,��7��Yz]J�xo�h�-�ٴt��$�V�m#J�!��lvr�8\n���"X�Z�t�w�P=�\�T�9,AySa����ⶦA[��L�Ă�ܬ�*��dR��"ԣ��a�:�l����8>��糜`W�\�G�q�q�����5�f����E��� �X��Gw9ޗh��|4֙�d��8=��Ww�#�.�Y˾⣭wz�V
tȭy�֘�����C�C@ ���k�ȾF 3θ���=!Y�]^h��tY>��tyjL[ع`��X7=�����ݽ��|�*LT�3L�c�<2"_'�n�6�yW����ݤ#W
��e�}tN�u��:�/��:�3^���9��Q�lS�,Oޙ/���7��5��,�!ƢJS*������z絴8?��$��`�y�nA���Q�WZ�J�(F�w
aKV���^�z���ݬ/���oֈ^f���{A����!�b���a�w��6�s�V��FVE˗�aA��5�
��ɺ��Msz�Uy��袪(|w��V��gi�����G	ҕ]�3:mÞ�]��y���o�����-,(��G  M�ݧ<�	�c�;>�}}��enm&�1j)�7gu�l�(]�E�kt�sNRnz,�N��j9�FK@��!}i�1 fO/i��1[�2�|�#��պZ�j�5��#�Q�G����C��	�dU�-�77Nw���g��Jc~��^��f�����.ic���F���6��y���iY��bn�Sf�_g
���.<�P�Y�k䑄�K�m-��YK�7���U�J�=�=��k%�V����+�m\}�rR眯�Qc������,�y�3t��Q_dp�z�!8L>Y�#�ь���u*�O�K0���Hv�;��3)��$��N<Ud9u&�.��Y�B�P��W{��t����vV�!�r�T�{�h��گk��M��}r#]�˨��|�o�X���M�������NIE�ߌ���o�k7�
�$�XZ=��a��BG�)��\o�ȋ�$l�|"� �s��0�:���/�2Ljs�=�I�h�F��s�׸"cD�Ȅ�͍�P��ۘ���|ʬgo�g-gQ��b�,e���EL��k��.�����|B��N��U,����x��4mZ*�f�h�͗Z��3��G"���\��M��1]�f�}:���[�Ws{�1�;� ����������Q�?b���@���L�nu��3�����\��=ٯ��	�-�v^�Fj��Hp2��Od��ø7��0ݜ�̌��m���[ ���=E��MYb͡�J��9����_'/{Њ<7z��VG�0 F�
�[Q�"�Kj)�k*��b���EF�1����kS,�3)*��[h��V�DF5���m"""V���*2�������lPcl[m,m��Q�մ��ZѢ��e[J������)��cmm��6TF[EJZ
����B҂����,*)e,�"�*���D��1QF�iF,�\eX��m���-YVֶ���!r�EV6������X�UFj#iZ#��-J�
���
�Db�kT[V�ȕj����2�Z ���JV6�Em�U�kZ�DA����Z��DaZ��IdR�E��b�*�0�,AZ���((�6��������F�ՋQ�LqW�Q���̮2Q�Ԫ�1F*&fdKIXڶQ*�(�j�1YR�[�������QG,��\�EDX�RҪ5,m�գm��EV �J1����"�J#J��>��ƾ�סoJ׌^{�M�sv�� �����#
'6��]�f�Qk�zl`e}$C�T�(\w}���?[׼XO�ܴ:*M�TOJכ�����9"�^�uںJ��J�Δ��z��#���V���}^;n�3*S١��k�J}�0���B�=�_j��S�+_��ך$s�u:>���<��.�ٝ`�{����a�Pɉ�/L�s�И�\�ǖ���sX�L��k�X�����Ot���lu�:�� nSw�(�A���=ȯ7���e��JK�b���hqx�˱��b�r�3T���|5j��'�.�(�ы\v����73�ފ:�u�uc�`�g=���߰��ͥԻX�2��c�~��l �j���Us�s��6��u�����qq�ET�_*�B�I��i���s�k���Tz���ᚷ�X|Ե��A��~|w�>�~�v���O�\k��G�tT;��V����箹I�^�R}S��|��a]A�f�� ��"�$+��W�n��;L��m�v8;�b�B�{�.%yv��5m6����ܗ���v�]8׏�SX ���5놣��}#�q�f^jc̻;���i��7�D���&A&r���a@5�;�N[@-7$�j�\vr�vd�*9�A�.���w�ϟ:�m��Aa	Qkʽ���:�ba�&��{��r�@����Սv��q�ꏏ���>ǎ��|�����7�U�w��Tި=N7ך����4�_Sy�=6�����{.�9�jWOAk�J��c�	׎GEB�]�+s��U�[H�\w!��9�\�����Wsu�f)�N�����ː�ℭ�'2���Bȯ]z�L�;�lS��齰L�y.�9���ϛ�@����6:�p袷յ���eP�^��:L�7k����t���"fQ��!�
4Ӣ_`STp�xb8T��m�3cg4+v��;��$U�̀���u\}	%���=pʮ�����R�����G�|�F�$;���Q�:VR#p�ΆXs�����x�q*|j�_�zn7������u����z5�>m��v��Z����ނjK:K���P��d)�3������*h�z�:5�5
n�iվ�r��i���2��EԳ���g��ƕ�W��e��6���@7Z���ȱ,,γ�D�z�~Պé���]�ʤql;s�1 ��ݫ;�w�«<��Q�o�`R��g4s&&+����Z�.u:�]���q��gvLӸvGb���{��/ )�\�n�u�SΘw��W��O�o3���H�4]M��b�;6�������o�`�:�o�aFß^����!�6���Q���:X3k��8�z�����v7l5xF��m҅�aP�P�/��WD[)gr��Ui�y4�8�g1)K
$�t�̑�8e8.B�b{:��k�H�mT�V!R$��\�E�a��bq�\�{��_�fϨL�"P�j�5�AR;�4�wb���(V�< �Ԡﮡ��4<XOl����lX�7�
$��L��Pn������g�t�"9ɕ��=s��c5�Nkd��5^�R�/q��P�q �ž:͓½B��]`N��,�Ƶp���
�6�^�Vv�1����"��'0�R�%��Ӭ�ҵ��p{L'�Ӻ5���Pz/�/}:MC��u���5;<�ݟY�H�O����Do����]��q	�����ۖҌ!z$2$���J,B�p"��I��Y6�)�/��޸O��@|G��[LdW�㷴�bA��gU�;x���F>Y�Zc
԰����� �a�bl��<���;�B�����Q�ݳ];
�u��X��)�:A;b?74��nU�=��v<����C��*ݖ�-O�Nx!��u$�O�����\�T�9��l��7���$-�sS�%,q�g�RΒd����ƪ㎊������]Պ��k[�b��Wf_,<|=�SsvS�-eo���J�y�V�e�tڎ�6!�>%�T�}�3�!(�>�x�q�o�X������> ��n�%��U�umZ9��)1�.�8���؟U�%��7n�5^�]>6��G1pѽ��xS����<膝ߣP��MEa�{S��%�9GgO��u�am�5����97�E��U�bF�jY&��M�Ӯ/`J�䊪޶�`~vū��1�L^jtםyy�VF.]�VCla�y���`���^݊
��Gh�ފ��K\���8;`c���ǓzrL`��[�4��๓�U�}
�d���]�I�=��q�U�0tT�rk�n�R�J�P�}Y�ȝ2����T�tN�!�O�x˙�;�~��Jq�0^F+�O:{;E�QS���[�$y�ܽ"���qd,�1ЗP�ʝ��� 5��z��ph��#(�I��4��NF��)o<2��z����G#�c�6L�e�6a��|yF+ڳ>)����`3��D��l]�Q��g1+/���j����il���2^����+�y���������?t�����s�5����^C��k��E�B��������DD�eY�n�C9�H�8|�T9D��md��jȧ~�[r��C'\��S~ݥu�{���<tOb"ǂ����3�āDQ���I˧+���S��{�����8��� e�������^�=�O��V�_?(|P:K�����Mٌ��w|d?*Z���>gl�z)�S��6[��S��m퉫Q��b��
�1ۺ��1�%
���(F��Q��dv){����T�.<�*��[1<�
�yu�IGm��,NP-N��t*�ƀ��
�e"��[Qd,�hf�;q7�^�ڔ'�9;���10�iQ#���똬$�熧��]5#���Wƽ��BU�59r՝���[����G��TXq%��N�����?B�{n�0�����S\�{�GY����Q˨�}wf��2r��`(��ymS5���H�n�dWC��\�w1kfh��5���kƖ��~��p�Tf��r3��$�s~�4F��-v&�<�����z�=��U&��	Xz�t�U�g�T��BP�P"�e9��w���ݺ�9����|xY�m�m����z�x'u�t���p	����ǡ;�3;*�OP��ZWs�\ނk#4�
���N�ь������5�}oP�]�YjК�V2�絩�u)!���P�9:�k�(VN�%æq+�bs�7��5]m~��t���55Gx����Ӵ7hh.�=������*��Q<>������u��,�:��7e��]�| t�l~�^�wJ�ڕ
8BQ~�9�c�=�e
(ة�Q~˪g�4Z�n|tʍ+k��wS�oK2M�k�c�`7-w�`�e�ۜ��� �u«������}rý�Δ���0W�����{'	j�/���z'(�n�!\�P�"��3��[�rI"j���v5�si)�a~�X��4ɇ���E�^Pf��ʕ�IJ��IM�sR������u�t�x1{6MT����)B�t��'IFk�F���c"�kע�l�3}4Ku�܋�z�6�U�t��$�;$��B<�2G
��ҕ����Q�s��f��)Q2�M�w\�;Uv)��U��tl-;E��W��������Y����Y��#�N���<�x�>W�Ժn��9O˨	�*�c̩����9�%t���[BMd'cD��AFF�Y%#\��D�c��
�kT�0�@���0%W6|vPtx� �g��Ы�f�"�>��ѡ�+˝j���q�ָ�E�#�=�OA�OL���B���m�DWяx���Xˮ��Lܪ�e}:���+ܹV�;���rS�ó�]�W.B��0�8k��_(�6C�9T��Ĺ���j�#����Q!�oa}��r3����� �B/��,�j\���]5��������<34�&"�K�����!�@E�Nd<:klm"�&�h	�!����%T�H���[oZ�����Ui�ÞmGU)�a�����'�@�AX�d)�3����wԉ����z^C97�on'-j��h$�n�s�J���k��4X��_��
Ct�?�n�u�<��~]�k�ܿ} [Q�<�\��n�jVl��/�7$XjQ����9لP��
6ĺ�Q�!��ꐬƸ����[�]n�7܆��6_�I�Z�[�ג�U�i�U�K�f���L�2�7�y��-A�8��n��J�yR���,�;���Aݚ1��>蓄qn5���^Ҿ]�+{��[��4!k6S�뭍V]�{@��4&g����2JP�Ua�����݋9dW�[��X�z���C�v�*�>��Sp��\��B9�%X�&"�E�T��M���T3��b;cG�6�iT�-�p H����nI�5�m���a�����{�-�8��QWv\ĵ]W5(�RN��!�
����N!�w���'�Y�Z�uT�������k֦i�u9ͧe9r�w���:�t��К�[�/N�U��گ=q������O-z���!�X�C�\��D�ٔEF�3��Q�D"z��]B3y��y�,�۞K�/ϸ�'^^��`��E��tu��9s��%��0yX�	�t���]ꁗ�d�!Ӊ�����ى
������4�XN����A��!O9�
�Lqs�Rx!��D��Ն�|�bU;�_�9C�D�����=	��"�3����a���_�9m5/�'d5����uL�UԶ,�n;Dz��B�T���R�j1���9��+����t
:���r����s���ʗB���ئ�xc2���b���sdV���[^"�������ü�d��|�R��0���v]3�|*R�;J�������s�^�g8�x���w;��)���8�C[mWa��l+68S�y���+J�Oz_��z�����_��j����=S�)�M�9�OGg��-�X>t��[�C{ù1r��왗���Ζ�soh#�!�g�q��'c�s�lcے9\���Zt���𡹋SkM�0���Ɍ��Y[ҫfZ�&wG.�9kN]f'CDp����T!���|}��53�#[{���]���BW�1�ԇ#��9�о|o:AU2�(��rz��ٮouE�Kq�]���m�7q�ͽ�v\�֝~��b��˽
�Z3,��(��VC%)� �\�UAx�۱	�do���9oN�/��%p�qӇ	�4pTθx.d��қ��qn/��8�n�����w����7m7�6�d&��(sˑ<g˕�J�4��v�_o�8~]C���� �u�^�<J��}.R�uȘP�T�!\�7c�qdg�k��B�X�B��&:9��A�6E�0)�(���{�N���3�����qߏ��G �3zQ彡R���L�n��SsϡV`�Ll��#Y��}с��m���N)D��]F��$�gܣ]JwA�7�P�嚑'��0c�m���3^�A\��Û؎��<цD�F��uӟ9�)1�c��k�7����C�Z�����2�����E#��'��S<Nw\/n��TsM�S��Fv�D�SBI� ��^�g,<.�ˣ��u�0�{G^$z��vtIɲ�C���l5S`�Lm��x�E �����
�(a�N���!�,�v��;j�p�+���ۻ[�Q*�/�_!ν���;�P=*�t��z䛪��.R2ɝ�W�9w��)�'�r�U�[�5G���wv'f���D�p'Q�CFV��$�;8�֒���N�W��	BOO�;>j��"���b�<=�<�c�gaǇd�#��ߪŖ+Z�Y�3�b�����El�j,GNAm�B��+�0G��23��wk�Ԯ�D�O�F�,���fq:���dW�=��3h��1`�t���VQ"�'���o9�+���
������8�:�	\ڲ�3�!�ذ_d���FE����ը�3�{x7����i���Ʈ4�N7�ʁ�D�no��o��w�z�o_�~�2N�Em�@o O�ׁ�Y��$3�Vr���L�T�>�}��,�VP�/j�,h%��\}L�S��2����3��ve���c�iv�r?�DU�W����R!�h�S%�l�JWj��0����rΡ3g�Zu�o�(�(�HȑVc\wv���0�T��ՙiLdW��+��r���ʰ�G�D�����V%P�n,W���m�\��@�S���$�1��Ђ��dC���>�����Q|@��sk,5YEۚoi��g��)���n��ea]]:E{���5�!�>x�#ƹ�۾l���N�9X'���9����,.�v���'K�'.NL�nI^���faO�ƛ5��}�NZ�Y�!`=
/�\y���5�0��:�>�k��ͫ{A�!����11�$=B�c�G�TE��R1���Tפ��]5T�H�T�񬭵y�e�����1���2;ė>�]�D�Y�#:�yM��_d݂!����, R7��̧��������#U(�G� # �HX��+��[Y�)����7p#�觕pT�ˠ���fmo6_>8.�	\6*r>���8��s�E�qXvn�����y|h�K�U��d{��b�0�H��\�w3qBܘ��H�ga����h�ϲ�����N���h�gC�g_l�WF�"�iW�|�6�ɼ��&��`�y�gl��+y��'_)��U�����T�.ud�x��5ε���Z4����Uu1�o=7��uj�*�%�4�6	��Ҙ�Ř͔b��s�|�罛~�[������f$'mI�,U�����IrL�h�zPLg"�
��e0��'{�h8����a��|p�M9ԭ${�L;tcU�3w���.�.jϳmӏNQ�hvx.{����wu��¨j���;_�g�HԔ%c6F��x`7�w�s!e�L�_--r�*u��9尊X�f`|1��c�Ie�g=S�SP�w�U�`A��šy����rIi�q���ю����	8�]�I�������6b+��9�CEh�m�����ϳ��2�܇F�!��I�գG�.�`0�R7Vy�V���YPc�J3-���]���*�&St��:C��
�$fTid��,e]�l�v0&��NS��.�����eػ e�T.�U#�*��E*u��,��ue]c���N90�u���Z
� X�2]�&�N������X�I)Z*C���Mx���ւZ�@C�E��Y RO�e4pF�8U��TQ�+>X��Kx�$��jF��dn����
��V\v&f#DIi�k�VKK	�	RLhS%�,��F��Qtq�1U���X�-ʙ��s������o�l�hZW����Ȳ,�D���?@�#9��J����M���&Ӟ����s����h�<1q`�%H(��P:�).!a�]4U�ڡ�Ll��N�C�G@���h�'!T�_���f����#FI6�5Јmfj���Ơ���8'|�[֍>&��4�%�u���ޠ^S�����発�����"���n�(�^�"�����U��ˁ�F�x��39,�w&���#�bû5�U8-!$
D��:�V:��[V�h��V�.����N��)CoS�J��j*�0|.��.��X3D ˕mT. �~|.��2X��͢.�[V�Bo쐅�ܻ�V�8)^��B�!F�� 12�2�TiFժ�V����Z5�E��ʵK
��kaiAJDZն��Qh�2UT�PkF(�m�,�T��kU�h%��"*[Qc�em�1�KiZ��KiDTUAR��eeF�EQ�#iX��Q�im*���KB�PQ#X�F%j�b
.5Q�-�k+m �����"�-a��h��*��iEY��Q1�,E�+Z1F+jQb�5
(��P��"����1)�d�bԪ�*"�
#EE,b�h�K�+QUEU�ԌUb�T��Ej*�������B�L�m-�-���
[UEF�%aEX�ګ
�(�[Q
������UQUUkT��[-�����"�e��1����D�FJ�Pbc�Zյj�RҢ�+�V*��ьFйj*�a��R��X�ʕB�k,��b�(��6�UU"��5)j�Zƥ�J
5(�+R�X��V6��EF"��OƉ����C�Ztw3��X�κDZ�����Lq���6v 2��M[�֍%��L;�T�{��4�m��nCm�v�Ri=����Ж��D��g�A< 'J�$؈t��8��g������'D{�+m�Xvi�j�+aYR4�O�oh��Ю��>X��<+�e;M�\<�Va��lO��v�����%}��,��4v#�n�v�g��:�o��S��d���R�i�{��f�����9v�v�F�-n��kڷ�ҝ]��%��D��wʪp袴V֙7��	�A�jj������FNLY�2Xͱ�PF�i'D�Q2l�.	�H~��y��lT��9�z��\�j<_�N��U��a�##������j\���6���ʂ�7,}�˭������H�q��6C4��C��<��x��Q�-�W���[�k~z��*����	�ɗ���A��ذ��?��ҍۮ�p?
�F²� 3��։�����&5;��������tLcG��4�Z�-uSJtsU�mu>�<p�܊�'��*��n��)'��-k�'���6��M�7�IX��w��Ұs뒍�a�r��@�����k�=��P5Θ�N'��4{��\�̺S�JΫ~y���`Ż�=�Ú�cGngg:-����/�_�=w� �F�� ����	bV�xku�qWL���7�t�_d8�ZpqG��g���~
��h=b��q;��]�˪}"V	��QB=6��Mv���^���`�БM�N�Ƽ�Gn;��m^���OE��(���Ui�lU�7�+/�S#�ܕa��6�Nj��<`�[�ܧ�.ǂ�`���uI�"$v��>�j-h=K\䖏�#�xJq%'8���
���݋nY����}86���p��6���g�����S�h�cd�p��s�����5�gbg<�&q�%���]��#���"�FK�K����(^��g�.y�T`�Y�<��В�S�n���]V"�NQ~	�q����]B>����Sѳ��8P&A���莙�.��E�D�����]r�MlW����.�Lu�;�i�=�:iԲ���c���i�^$p��)���GQM<�j��`q�$2$k2w%�p��d�)��qVS�=ܟ��hd�i�c��,�M��0p�;�j�
�����A��.R�o*t��G��v9�TA/�n�C��M�ȭ�
�2�
�3���p��Ee�<hjT���G1V���{�4��E۶�뱂��0gϨt��!�wB���ٽ۞��$g.XT\���#������a7�%<�b>�o��$ST��U{Ʌ�v��8��a^�}��x���،J��:���q��t��E-[Hg�ۆ�m�K�BJ)^��f.%����)�����2�]?��U�v�.$�kA���?�3���{w.���k�o�#bV���q/�Y��װ���V�H���>�Q�-ڻC8]��Z�9�z6�3�]�83&�>��ޗD�x�����s���9���l��S���{���=��i��%l���r�^���1I����}�1���"r��X*��#z$�O)�����~UAn}��F����(��U���+;��)�������֬��0��s'���B؂�1n3�v�;�`�7p�ode��QV�L2�+�P���%�@�5��n��|���Pی�r��t�|�{V
��-�+cm�g�]"4�������H������d���{�Cu���}��w�4�;�î"�r�Y��Nn��v;"�|�p�(�q�	�X,�ݩ�#�f%l^�J��*F��h>��-����q��`�fTI�'QL�0J9��6,LVt5������z��v��a�@ƲS�x'yu#Dv���u��{h[�A>Z��ԙ���u�ז+rh/;t$f�s�,�H�/'�[������/��p�J��t�u��nE���u���FK���b��z��˚���TW�V�C�����&��`t�o;���r�w��t�ڙ�'άR��7&C]!��Oh��Q�/�**����7�b����UX����ݠ�Hn:��v	஌2l��d�"�ܼGwv��Z#�̎�݇$z@�:�g�;�!�v��((ҍB�-��Y'�J����RP��3�؛'HZ��=�ױ��*�i�N���L�W�j!p�m^R��o�}��*������tkA�P��@~�a���ꎯ[���OT���0��mE�C3g��f��5�{au�8d�x)�uxlAn��El�j,��*rs F!bs�VM����ӥ�Ѵ���{���5�کQaD�go��W1�^��ٹ�J����aZt{��Rft�2���=dI�g �El��2�:�)�̓�R�躁���FA2�]���7Hdb��� ����~
�ûQs9:�a���ج�.ܷF�&TԮݷ�x��"��D�F�-E�nF�:3�T�vz�$3�Vr���L� cF��޵�G�i��P�|�7�oy��l8]+���ve��>v��Y�U��'u����/��nV�lvf���]�o�iCM�f�ge��X\��=tC���_�ಆ_5J:�/G�	3tF_���I�s�;Rt�q��p|���>��,꙳�/����c�(׊6R�(]}l;�놪��4�=��]eX
gv{i�
�$<�q�4�NY���΄s�.�ˌQ�
��@wH
]��K��Փ�k���kI�x��W����S����Ӑ�i�����;L^�^��kb8]دX '�-��L���DЎP�M���ӤP��(�rH��d?oT�tR��I�T�ze�w�c�{V"3>'G:��Mo�T�\7��������k<uF6g��o1GZw��	n�w��`�D�o,U�����(�0-qDn��^������<�]�i�79v����,/}��fB,����>v��_��:�o�U	I�2Fapӧ���
�f����3m{����OD��!���ڵ�N�}��Γ~�@�8�٘p��e
�% �Eis�݃�v����������;�]�R���p(�N�֌ɳ���ds��H���N��5 �;��Oq��U�W�Y�����v=f��]�W�5.,�~i��WĆ�dΨk���1�u�Ҭ�f�V�:�&g�P��-�bS�]d���]��44�)�V������O�Ȳ炷x�p�<g.�C�/)k������,���E��V���vK��(�X����J}9��Q�L��n��X����o3��AI����8h̔��t7���q�f�Kl'�����E���v�s8�>%<UG-�W��U�%�s���wed�C	]J���4XU�])��IXp��@�<|���H�I�.�Uwy���)�Gܢ�4�3[�=���V���ч�Ŋ"��:Ӻ�r>�ۭ��2I�c��M�v���ݓ�	�*J�5#�x��W�s��E�0�lK�e��Lol].Vy�)�����=�>���
9�u�����!9g��^&�5�*��������,s��-�c=;Iדzv*��(>#�k�F��p��S��NŸ�ܧ���R�����#�1�B��s5.��rC�u&8�D���f�dq&B7�(w��M����ݍ����p����-�J��b2Շ��.-l���5D����p��4�r=B��u���t�j�-�j�yŅ=�NJ���,k�;i�H���1�O�R�3�ĺ�:8�Tb�f��^�%��+`[ʦF��Yn(�a��UQ���0-Oz6`�@�J"b�9ۢ!�J%�(��Ua�wP\����s9�;�]���/��Kpx��Ax�˗Ig>�&�U�
'��J�P��i���qbȻ�k&�)U��JtvH�k(U��A-�ͷ���\��|Vc�3�ż�uϫ��@�|��Bt�q�q�Z=VجT+ݿ{�v��ϝFԝ�5��(��Cb�{�ex���'��G��$��r$�*Ӡ�o@�!��y�n�i��B�$���e�[<��V�m�}�B�ި/�'������v�L��5�����랒Bޗ58��Z�̥��ʇ5J��tv�Ŕ,S v�����^�"�n݊k��3/��>u͑V�g�٘"
���}����H��]�r��>n����#���E	r�.#Hus"��Y�qf%�h��ۗ�\����0<U�<����Ʒ2rtsܓ��1��g�rHX =���ꚠ�C��4��:���9����"��&zi�;�q�s��m���'�W�/������y���Zi��X��⯢A��b�w\�?N�#�����{���۴�6
8�*�v��s�N<�#�l�Dr*��j���ӤÔtV
�"��n)O��z���8�׷`��M�Z��9	�WU�	�۞���TYh�=Zn�u��s'��B�6d��n*�5�����kW��O��Y<�'�:�}oT��XT��ْu�|w.��2��eT��Nn��OԜ�K06�R�Ѹ���:�.���o%��y���0Tu�1��}y-��a�HQ�y8��1o�
�v��̦���$|����r�w���t�!�D��N���N���<��}K��Ra�K4�����D{���̮����=+��*����sc$����zĬ�E����ג����ҵT �4>��oˣ�vy�ug<|�&�~���0j
���%��I�'��.=�(�8}�*�Y.�Z��� k;�������U��;V�G��]�4�>��v19�l=�8_���7�x�Q�(�'Kͻ���@ ���ik) �j�.�rb�^1Wg˶��h{.��o�b�Q��w��Y��C���֪soH�O\��Aj,F����~K�x���fQ�osЊ|pp&#��غޝ�����2�,�퉰�I�A+��>�*E�H2Wd��3��QKq�f���&wfy�sY��}��r��Z��kɌ�k����@$q�͠�V��+ҝmD��3�ݕ�m��U���QE��r�j!���ʈ��b��@7�����Q�GNq�+�߻$�\����
�\��]#v/�Kȉ�	Ď�,��ʍQ%��N���1�^��Lt_��,
���}Q��pz8J���2�t�f1VU�q�L�W�;���qTV�KU���0�@9�F���w.LzU7�YÈ�:���$�M)�}�fB�+�C�s�3|�;�Y����\�v���rfa��u���t��[ҫz����µ,]��30]N}3wRSX���&
YF�ip���^���pSA���e�n\�=4�7�����V�R���.��pOw,謪��hf�U/�]�ʹC/��6oc��Չ��*#�{�blB�S��܈���U��
�̟�r����b֥�����w+�]��q���Gh�C
��Dn��PBQb\ᬞ���Lp�,��35�����u��@^uss���ft�DQ�y��f8��"
!)lUC������]Wb��A��;�X��<�z�v�!�^9�pS�v�Vt#���L2�D*S����{DN�i&�?\׾��*����M��Ӳ!$i��ЯbT8��wN;�Bșj�#��5��~+_]�5��J���~�$�t�IW�
�"$�(iM���+g�jt�T��t�e}���o���5�B}�F4 �G���c�7N" X�Mgb�>G1�ù,��yJ��ܜ�_���b�qG�=Ts��J�@�dHf����=X6�uא?�&뀥�#ƙ	X�K�;��n���R}9��F��9+��l[��b���O-E�ò��R�	���N 嶆����.V���*��e3:8X�y6�F������M��2�n#�͡�b����d�� ��3�.���'*AQ4�s�CJz�a���T�{}���c�M�&�����'�9Ϳ5BV�{�;�:���������:��6�=Q�L����lm�T�C3��j�d'D��4Nco	)Ȏ�����x�(O�4ZC�]�&ƺ�$��Ɋ�D9���I��ȓ�:%�yMQ�`��N-�a���84Ɍ
rC�5ceV4L�a�����u�J麚���B�c)gj�)YR>���}ê��jn/a8�',Hj$�О����e���|��^��YJzr)�s���"\�@s�~B��;�s����Xt<�F��GoºSnĳu����y��KzԬCofI`\��۝�G�~�پ�J�`��Ȍ����QN@N�%��U�[�x���iRSc�$��ڒ����6Hǲ2��ETq���K( :٬�����Z�;a��=^�Ɩ�_�eH۸��~��D�sÖ�{
ᑸ���U��u�OB�/U��ؠkE�u�-u�J�$�8�eё,��؃�,�|��E�[�nS���=��U�(:>U�ri�L�@��8�4��gĮQ��Z��g�r��}�[���30?�!�o'(�C*�bb���+Ab�]c����1H��_�κB����[��M��M�$�(m���<*��.�۽m0��ev�.�oj!�N�zR]&ɼ�{�x)k]A6�G�J}Վĥ9O��\�.[KQ��]O*����JTsn�೚8�ܫ���c�Q\�6z��N��Er��w%��3�O�)3QQ��81�6J�ʊ�ަ�^7!��F
��:��)
^&�V��]����r��+)v�c��:�z�O���Cqf���j9�ũX2��Ik��n�5Kg&FO�]�OOh��<�9�:�]�j�m��_�E��Ѱ�H�1��<�,�������]۫�����],�g#O�rSȟJ��=���@~SMK��Ce,B��j��\=�ܰS��ŷ�lvu���{�A��0g�ޚ�{k�Yչ .���[���-�kȶ�'r�B<8�S}��6&�8In��J��t��yyZ�Y��ږ�Έ���t�^V������j�i\5��:����R���[E���z:��q��*�|��ܼ��n���ͭ�Y�����.���[�w�:`*�
)���)e=V���ι{��W���ȅ,@s��³8[���4�܋�tM�e��Uݩ¡K�[,��F�8�kXe��[�%���jb���Թ3ܱ�M��|�
��
`�,&�u���D��A��U��L/�ʌ驔��(ᎲU�XT*�dvʳE�j��Qxyn�ʬ�(U���eYg+�c�a�Ki�)Jё��lXd�V��X��B���,��k)����eIv,�80شZ6.�m]����
���<Մ=@2�"#�b�-Tf�8D�t\&f]S�i����L��4�M, 7�SRĊZ��"�r«���n�C�e�6����`QR���˥�� (�k �-I�)�W�h#7M#Ld7� �ō��	��{��.����[��6>4��
���4�b ^X��#&c#+;��67WV����h��g �Xzjd̚%���`J�F�f�o�*�Sb��,�`B�j�q�N�4 9t �	�O!*�ʁ`yt�)��UZ8�&��5�]=�а����/�/Vx�}��x���"��͔��гr�c6�̢��fmM�L��ۻܬ�l�� ���?s�6��J�b&��m��t�3�im:�J�DK�QK�*�j�ͧ�
���M�h�J���j�iH��-e��	��f[�D�
wy�  X �p����TE�J��ZUTH����Tdm
��Z�(�(�QF"+�A�PTU\�b�V��ȥ�Z1E�֌
���
��EPT�*��U���-J�hQ��Ų�*�)J��2رX�DU1�6��.Sq��#iY(��`�0��k��"+iD��h%��m��
���-�b�h�(�Y.%�R�X��jUTP�U��ƴX(���Q�X��#R��V�b�����m��PUD�"2*���Q0�Ke�`"�P��X�mc[l��-h��,V%���TQkU-���X�R̵EU%�U�Ȗ��**5��Eq�����UX�(�V%�(�mb ��iZT�V���lQ���TA�*QUKlQ���+
�EE�ZT`�E�[J�EE�Q��PX��T����E+*�V��31�A-*Lj��(��[UmZV��lbER-�XT�Qe,��J�Ш5(���E�ETDQ�
�EU�TT�V���Z
",F5,Qh
�|>�s�̠[���<���֞_1����mc0�8�w����!�1�-�Hz�<s
�Z�t����\�l���^O��r�;2$�r��ڴR��h���m#�<o�
P�ۊ��
Q�g%Ƶ{��D��߳W�:==+�7�;#D3�`tX�RL��{��!�6.g��hky��2m�V�#�Į����'L�`��ytBQY3����P�uC�M�#�ts�})�[�D�H��8����?\q�O.
���>�7.`P���l��eC�8U�Q�iԳWI�yTΨ�o�v���e�i����/%�Q��G�E��1�x�y�)v�>��c���Ҵ���̇\��F�Q�dQ'm�8�ԭ��Q��e.���;U}�V�ȔP����ϼ"��o�p�</�k6��n���nF��!���W`��۫��9R����YI�S.6�EPdW��5έX��z����="ȮL��Df�,�<ܥ�<�ީJ�hI�W��3�}��������w���踍!�6.˦zυi��iX�ƽ�
�נ/����Yث���61M��lJ�Q�9c�>�s$%�^I*$Ҟ�yoO<�ܢ�`��1��k�P��D��F��X�T�V�dk��.�Ϻ�9�[@٧���L'��0�|K��僶���ٯ��U%;u�8�o�g��6^���r&�Zu�lo,�F��58Fee���ހG#{�Z�w=ݴ��X�Q��p��67׽'N�tV��b�2<:iA;�q�{�W�q���o�Kh8���f}3S��1{�d�t�_���b��͂8�h0w!x�)�L	`c��&��zFd�;1�ʜO&���+ݶ��Y���|V��>mVx��SDAs�I�6PGr�cs��h�5j�<C�/-�Α�5m�E��v�,�YZ�F�x��HV�P״��HpIQ��i�1��R��ʽ�x�.f9�÷�Z%=Uy��s�Ȟ1r�5(�ä�i?-�^O<X���6���ɜu���ǵ�ħp('�6�n�땖��8Q	��3�ʠc�Yj2�^Uz�/e�X�b�5������AW~�%���9:��ù2�>J*Y-�*�����Ih�����\�N�T	��V���[��j��']�~�#�D�b"ï�̶�cݞ�(H��k0J(>��	�i��a(����s��������>����Kܧ�R+�l1}6`�sE�0�y`����<n��غ&y`�S��3a��+��{�̧=��T�����4���fmj9=:�Ü�V
�ǭ�Y�f>TZO��U�H8*��N��8�jԈ]�Ƶ`q	�ɮ�ף��E�Y�ФΩ��3��w��L���~�re�9l��Ov�v�a��I�Χ�7�mQ�kF0�ufl��L�(+��{3��c��y�L�xE����g�]�����1�&��,�%�B,|agx�Z�i/N��=ۉ"^5y۝�6-��f� ����3����.�D�������a�H���0�Y�.}ʳs�ɽ7���[J&��|�����&�xlG9�R���A�6�*�e"Ϻ+����<�u�2�vX�_�$Ê�I�4pT�Wyى�[>�pɘ:�/���z��#.�Y1�Gd��gKȉ�HN$�,���,��wG��dW���wNv9.�ʆ���1ьOQ,h�(�ΑB�F��B.6B8�Mm�S5�;w������Λss�fQ쏸�3/�U{�&ã�F��VVߢ�9��x�b�s�G��]�5�<9M�;	� i���݌\�����]���DqC��SO�������*Z��s\�=K�e٩��="��N�HGZ��W���1�����rU׳B�.vxD��W�%+�s��L�K:���<��z����t�\͞9a�َ61L����c�Vðg2�R��ƒ��g���"�GǾ�e,�CP��/����*����
2���V�9cf U�C֨hwH�wG�$������3;�F�u�����+����� N����xRH�#.�e�y����A�ӹ�2����4�6=F���r�vD����T8�Z���w	 �xb&����"�b����ټ�����H��L��"k�<����)E�i9:�Qy�m����s:I��]1�^yj��^ԑAa�R�2L[$�9�#�3!�}���,���}�ۦձ�Xޤ��OY�^�0�{�-�U�T5TJ��dHf�#�W;Y1%�'�����������m�=>����]�T���)��۩��%`���Gd��v��{kP��l�429F��D�C3�j�b�Ga�A�dco	Ĺ�W2�<ƶr��������ѳu���ǁ�Fǅy`�"��2��B�8%�5G�G���8��0�E���jZQ�F ��B�"��`�c�f+�|��_��,+<<�I]�.-�P��wgR�VRQ�F���U�=��~��#U���z�dć#�C/%�ו]�Y��Z%6�N?<�z��U�FxL%r�L	���rb�,���!g�)��Tᬉ�F�}N�9����^y�5g��Xy��Z�uN���)׫z�:,�K�k�켡�_
�[Ǚ�±I]��8ʿ+==�k8r�'�ks|;M���^����6z+t�;(c�����mi�(��Jнc����..�n{f��Q\�;�q&�9�-��p<gM=ևxK�1��[���2�9j�͍�0p�sv.a�u��W�+�)�������/�Gڠ[��F�I8�`���	�R1�nt���]r��������܂ݬ}EV�����S�����t�~��ʛa�~�`�B����˸@<�Gj����g���E1�*���1�Ԙv"E�@Ȟ>�_@T G)��-)�tI�2�����W�y�CB���]��;��`+��m��3�4¨UĞ�*��GX�iH�d��V�s��{;�33}��j��J�\�� #�ܲR��dʅ岦Ԓ�ӴLܙJǹ���Jgi{8�U9��)^f�:l��9�P�s�;i�Jt�w�ӎ�Z���3�#ђJ�Ugs�.�T�N��|�GT]C�F�����Ui
�{����Fzx��T#��s
 ��jc9ꠘ�X_�����5�2[�ug�WE���.};�+��`��1��%伊91V�ЧV]Ì��E�=���8x���灮ɳT����`���fC��n�d)�hފXju�����D�#�y��(���\Y�a���f�f�z��*ʁ*Θ1��(���5�X+����/�V:. ���t�|��XR����3�?hZg7+(�r�c6Q۲�)awG���K�Y)r�E�.wd�\l��[������d��}F������Ε{���r�����PL$יS�RhS���ػ�m�+��O��D+L͛�zX�(�3��P,�<�GVA���뫁ا��,�倫7��>}���WM��Tkf`��r#�SN���9k������`;�hV��;u㍩SgF�ˏ+��!���^��dnոgL�`9������c�3�.g�Ru���Vn��� ��9�K۔�+�"�+"�[��٥�s�8s��m�m|/{�j��n�����x9��:%�H�rA����;E*� ^׶�FܢMto)�
�H�'WIk�k�k�<̆�]�+�$.�|�`����m���(Q`�r5s�{��Ύ�W��gl��jJ�g�O~l{î���r�`�󰄥�������N���*���n�Xi2��WVI�����j�Γ�{Dv9lWH�N�8�n\�(�g�)0���"<+�,Z;o5Jcg�|+^z��'m�/co�3�+-q����S��
P+l�
y5u��/{�*͍ a����^w�d��z�Z�^�9̄�����^Y�M�:�hҺu+Լaê�]�1E��Z���u�������Ǿ�':��R���ŀ�~J�Nx�����p
�nk��
�1ɪȷl��~�b��#���J��i������Q�}b���c���A r
x��%�n9�os\ak3�Wjg�e���tP��0�څ�	Ӓ	b-�`i{�t]P�;��q�Ti��`�ס=�3��5v�g$ve�;�}�� 8?����X�U��.����!�wh+�A�Tw��]QJ3���?Wr����4���~�{�20���>ETz�N���{b���]n	����Nk)���u�8C�8t߆�w��Λ��N;�M ��P�,<�M3뮁];��J�]��})6��pDZȣ��5��;�ps�j�ɠ���9�:�l.�knB}u;ȸ�|��ZWbJ�!��B�gK7�t�B5�&P'D���{&,���Ƨ���������Ǡn>�ǎǂY�)b�7Fz���2������ƈ���*�$�;m�\&�P���1��ba��I;��(�#EE�5��ٺ��SA�02��NIo[cT�+5����Y����J|��.��i�ۋ����鎻\'v��l�z�Q7��]����(�'W����{w�>�^�h��w)fK���)��w��M��ٮ�h�f,����zF�{�����Ƿ�p0�Ҹ����fB�Y}Z8s��+�h�d������ G�e.�9p�j�Wz������}�d9�\YX�;�As7{6�h�8�О��4�s����p��	��Fx�~!`����jJ�	�϶v��7�jEh�;����T�=�i���:)��	:��h�L�Nac�H�^���~���
��_M�'ا��:H��Ҷ�4��N�c��G=}Ƒ�|����8�2�Tȅ�SA���Wu	"��8�S�v��YЈ�ܮ���z��+>��>��D줼*��*aU%�(�k���D���7B��*l-�q��j��-�ˤ�4K+eL�r�g
�p���I���D�s>�u<����)E�wZzϢq�X�lw�"?e�?^xPyj�$I�%(�`*�E ���߮��Zӄ��.��;�O	Ů]��l�����׸�ofW��Ӣ��5�����tq���S׮�n�S���p7I �D}��X?vK�=e�rr�yb�uR�E�����	z�8�wb2�^�n��5�s�RV(ߏ(�$,�!�̎{V�C�^�% �2N��f�j�#�����>�ң}ޭ�����/TW��Α��i�K���(EEY�Mh
Rݙ����0*1��_`Z^a1n-��׬��u��$H�Ƹ�S��O������hU�t�]�a�n{K{�_U�lB��������sʏ�Gx�N�}{�0=�>cT�`C>g��vxW���Y&;��YA�/�LcTV���ø�F�f��m����Z��H�EK=X`�ǘ�J|�ŬU\=��%u6��(�[3	]�N秺jjǁ�L��_j�� ���~��f�6n�dXL|D��*� ��6�� r��rj��/�:@����j��a��]:`��j�E���_�����b�]u ��\d<���w�h��>�oK�g=���[�^��V��Ȍ�)yS�1�f����u=l��bKF���.�2Fc�s�jK���ߥHǲ�;�I���;�|o��v�����Qq��fѾ����,{bJ5z����F廰���U9�n�uF4�\�����"�ݩ�j��렖��C<k�Q;��v���d-����\BY��r�r�ٝP5����/:��)��FyF�U�UĞ�*�����Ў�(gR��Y1�Br�wmr��T_��;�7��R�,�;��Ӿ�����0����oiu�y�M(�Y��Y���u�������V,�W����ŝI�������w q�r���i�Ĳ1�r�_s���Ϋю��O���5b7V�u�ۊ��=@\JX\�X�	��J5�;�j���S;ȩ��ǲ��/v	/uF�&�wLP;y�{y\wZ�B�5||,��IB89�]t��'L�`��wH�P �
�s,�!i.Q��5i�������l������t�{�����(�Br�ggmk=y��04�����7�&'a�k�m��'i���V$'s�����UƘ��	؈��/������j<zP�h/���ӧ7�9@`���`<��C���RI��6�;���6�C
E�e4��8�8�˳ū�6'n��9튿l��/���@"`=�T�Po��Z.�TĎ�(���i@�O:�Qձt���v+��B}M�0���y'ە�6op��9���vȇ�N���9����toS"�X,����)��N��\�r�iD����8brY8=�NIeݑ�<�N(��w�l`��n���������z˄�)����Y
p#!�*	�N��s��m���쳧��M���n��c����(�/�X�LYV��p*rBr8���(����	'� �$�� �$��H@�XB��$ I?�B��`IO�H@��	!I�P$�	'��$ I?�B��IKH@�>BH>d$� ��H@��$�	'�H@�p$�	'�H@�yH@�z��$���
�2�ϔ�nH��������>��������;ω
Mj�YH���H�TEJ�i�6j�EV�IT��� j�����+Va�T֔�4��i �/�=^0�Ke��[V�-X-Z�%�Z*� �	���Vfm��l�Z�UT�S�lM�1�[mZ���M�L�j�eZ��kv/=ތ ЉUH���&��F�h�Vͩ���m6Y2�i�mV��Z6�`کJ[Z��kjգj���YYj)ah����V���m�����ѱg� �y�M����V��� n;�*�Fô�s�Em��Ӆ��c@ꃺ��.�Aj��h��àj����-�Y��ʵ�3[u� �h5��ܴ P�:��X!ѥݸ����P�&� -�u ��ptE�&��5�ML`�R��<  x���V�`UF�قA����g@u��f�0
�wt�ۣ�h\e��P�8:T�9�f�emi�iU�Ym-�� o^�52c Ŷ4u�V���T;��(��(��7{k�Q@QEQE��x��(��QE�n(�QE{��(
QE�W�QEQE�ǥ��Xe��mX��� {�
@:w�r]:Wgt]m�ӧ;l�mlQ�ܸu�l����Ku�n�Վ�CMS\u��WX-��t�۪tk�Q���J�]�n�U��+��M&ƛgx  Y{z�t�m��;�-ig.v�0�waUn�uT;�8���Ӯ��v3��j�ֻ&�qZ�u@v�i]v��Guͬ5�5n[Z�;���[��5�6Z��kZ����x  d���S����wu:k���u�k�[u�n�խ���c�F���wJ�ͺ'u��5Kmuڮ��;b��j��4�9�����-��Z1m��L��j�aL�  �=;��Uh1�m�ҩs��%��n��5��S��V9P���`:��;;k�u�.�c:t�k���͹v�:��hwu��R���Z�Hf�CZ��ք�h2�� ����Ӯ����wuƆZ�����T�t+���ڷ]v�ʶ�wsmW-�tP��4�m���::�ƶ�C������FB���T��w� {�;m+MZ���T���ɷ6Ύ�E�vnZ�k��V�E:���ٔ�\���.�mgqWqWm:.ͮ�vn�ӭl��ӻ$��>�  S��I��@�h  �~A�TT�      S�2��� 4     ��%R��# � �����	� ��Dhȧ�mL��OQ�jy��H���U 	�0 Lp�â��8یeH�^�<o�3�1h2�+V��)�3,dg��Ri�u�1l�S<������R�h
 /����Њ
�O� 
 -����>L|��O�P�}a� ����H��?��$�N���R������u�ΛX��]}���"�G�4���j�&�:��ye�H"9���4sղ/7��\�����bq�燰���הU|Z���)�,��d���2��3L^e\3"b��,e�c�82�Vi%+�JC+2��l�: +�ɭP���km鲬��WgF�D��<���`��\v�N�&d���R"�n,{YJ�[k�nVhlm�+�7,Ru#y�\)��!ET��
˄d�[���Ϟ-�k	;�n�le�"�Im�];Z��<�n��]���&��M�����6�K�n(�݁{�+���Si�ŧ���V��S\�9fY�ܳ�i:ǯ^f冣+0�|�T��]d�M1t�T��F�1<��tٺ��;6��g���Ĭ�aS�^r0)V�����[Ia����XcDڄ$�K�iV�'uV�O5��P���rd�1&:ɢ��n0��Z���dϮQ�x[k
�2Z͔Pȵ�;{eL���cr,�K���ghQ�x�:�̬�Vq������D��Z[+CBV["�ʸQ���AܺOVjoasc)�j��4>�R�қ���r?�"_�yP����T������V�6BVI[|�R�N�#]Z�^M/V���bW6�5�K�˭&�U&`�xm�QQ �׎嗙�C���S,��r�a9b�5X�uYl
���b{k��́��F]�oU��li7���Sp�o2�E3�(Յ�ͦv�B)�1��:y���7X2$�GtlJ�fݼ
R��`"�h�Ɩ�
ͬq/�����f0��-pĵh �m��ԅ.��V�F�e��u��WgJ˽��ؒ^j��$KдؑFV����i�8θejb����fmn v�9VƚY�i���]����%U�e�n]E�d��xPr޽G�O#ؚ�ꐌ��`�L����oۺ#";e�//	��,bEj�y���Q�fL�L��qTQ�kkk6k�n�&�s0�rJ$d�ɂm���=�N�00��iж���1�#[���l���$�w+6�#p���H�t]�B�c,��l��h�w�*�=D|�u�̩����[�P�w5��w�N�ʳ����"�U]�oҀ��6�	�͌#7&��S1F�m[%��Ň-�}�>tml���`�B��(V�M��Ȧaϙ��4�@�fB%�Y ,�Z����՚(�4�����t�̅Ba��c�{������n�^]sP�E�*TBJ���8��3~0���V[�8�r<�dv��I֐��Zo)kv�Ѕ'�:RhU�*6�=@L���/m3��p�Z/6�e��Y
���b�j��9f�L��\
�P�Y1�^9��*Y�S��Ӕ��*R�e�ܹI��+	0�ͽn�ZN;d+5���.��2��o@[@�q,��o+1�Ғ�3����qA�͢��*h݊� )�l����$�d"`e*����aQ�"I�f�+t̡j<�V�j5z�8SX&��Ū���n�B�v4���q�&��#yz���6�B�	��§�76��"̰�k+h�t�<���y1Q��<w�DLٲ�Bk�
�[�ԦF��Dh U�[J�6/�#U��V���X5��3Wf�5�-�29oV�t�6G�4�q�D����5SPb���MZ�FҸK���hE��������I|�øNQc���鼻����ۧ��ӣqT���3�y�3A����џ�m˘�]�r�J�b�cfnQ����Qh�-��4K������˲�4ad����:A����Iwnl[u�%�ڑ��j�mԄ��7
�6��1ۙB�-׷ycq��f���؈�i�Wj��VŊ��@:F�+�f��pm�V𜈨^<��.�B���,1�Vl�>&�^ӥ{f�Cyb=��i��N��n�RU�����i(N��x�+���쇗�F(7�[�õ7c$�pէ��7�+����@m;��i]e:ےQ G�e[$f��ԀZ�[�%8���3l�Jj�5�n�Ƅ���ã�ni���T.�:;�7Q�[yw��_ʀ�*" �U�Ua���E�&Rk^N�$��`��|����;��cPn5�۵��Fn��ȸ�����@Ӭ��ˬܗJ&�J�a������ca����}m�4��V7]����<�h̰��JJ�9P"�.9[���5����9-�Ota[˕^�
+(�x�w�#�`�@!�R�b|��7LD��a �9@l$7��uR���CS���ѧ�X�	E�u/,9f��]�-��7A��ź]b�x��"��n�?,nw?������ޚ������F5L���٣j��w[P]]���S����or]��	2�Б��RY�F�z��"]�@Ό��0�-�ݖ��1�zu�A�E�R\��_}d�_D�0��VI��ɺ*ä��];1�y���TDmڇiSZ�LƦd�k>6��0�q0k*�CBw�	m�ڼ���SecE��޻�N����!a�zP9��21����2�q��b	�l�[�j���l�7i7m�+D8�ŕ��K7(�����@��[�n�<��r��U	EAo6@m!�rj�A�wɖYN�ڶ,T�o)�!�ۖ+v�U��:��&iڙt[��G�U��K[�\��3]-)��N�?j֫Q)8��f�� F�C1�YGt��u�v&�[���
���fZ;H�����#�4+:��qMK[*�y2n� �R�RC:u�{*��"YR�re�Kqb�7�SE�
�,x�r�H2��,+t�z#x��{>ǧ	�!P	yv�8�l'�-*�{o*��L�ǡ*[%�W,ڴ BB�W��+j�$�(�Dc��6n���b��/�9����!�	L�:I�S��`2d[�G�̶h	�Z��)a ��*�x����l�ID͈	�m�	`���҆��.�)iQB�8��B���Aq��-�fnia�nJ�V��b���e4�#k2�[F�	9j�5�fT1Է�Q�d.��)h�5hu�L�N���2�<�˧M��V�(%)��Pw�"��CM�8��p;���b�A���]]66���� V@o�WsU��^�W���9V�\���ږr�п�v��m��mW�_$RM:i�7 ���.�Šmn}v��[j|⩘�l^ۦ�W$;wY�!�b�E�̩���W�R����Q��md;btb$�u���S
�U*���Q�t�#x�B-���⼭� m+I��:���(i��zC	dך�[�t�!�n6��TEu$��֜|���'�0�{��Ҭ+m
bҁRd`�_�if:4��7.h�S2j JF��7v����"Q:֤]������.Q��ZQ�f�f@Լ��k/ �2]n����<a�ݼڰ�����R�KɏbP�&�n�ܒ����`�jVIx%�+/h*��d��t��d��7e�Ř��V�ũ�Z#�&����7i�<!���a�F���Vn]2��FQ�,ٽE�Ò�S&C�c7N��9��;��*)sjf�-h��I��J �.e3Z�ڼ�ॉM�k�T��m!W�ʁ�5�2�+�M3Ź-�n�B]2,T��'H1��<��$Y,�Ygv���t,6�S� Ajy�'f�)��SL�Kc,]�w72��	����F��ҵ�"h��Sv�A/Y�"��fdcMcT�ɛF�w�D�$
�^ȴ�Ŕ����!��X��m�hlC��Q�q�{x\�۫����C�(�×J�f#V���Z��C76驲��5I)���G�Z����,a�y2
L�z�~c^b��ͫn�Vڔ2V)�HRZ�S-Qj���{�2�/XH�v�AcI$�y���7�oR`�ؑq*���:��i\��NT4([���Mls$x�\�F]�W)��`�)Ys7)�~�ª:ə��hۙ"�
�#�9fu\�y�|�k)��A�ǵ�e��������"�D\��au�1N�e�@QM�Ϡ��i���6M)�B�-}��Y�-�k%��@%�,!z�h��{����6�I�.��
mR�*V��2�+4*E<�c͊�:)9�w�n� �_eAZ)�L!II�v���b���Tۚ�L���Qkk �Z�u�f��T�:LƦ��2��k���
;WU��*�Ʈ��P�f�k2�Z�.���N�AS��r��3 oH�Ȗ+�Y`b_e��:ɥJ�(��6j�T�̼��!��]�*�@	�� �֖�ɕ
x�7�H9�*7Ou�%�Gmb�=�-9���r^ȖVn]BFN�쭑e��r��g�*l�W
Uɺ�T�VrJ�m&Ui�)�V���X��R���NP�5��ԾE�t�ʋB��(�E,�s$�U�ͻBޝ �4v1���MVHBBʓnE��2[z�Z��yREE�z4�t�M b�,�hx�3�Zl*L:�U��ĺQY�j�:bVBڤ���ہ��мwcƯEiR�i����N�^�7�i�Q�&������6�XY�vT���)cYmXD���d f�j��^	Wf*�R5���nJ�ӣ�!7&EYd&t�Kj�c8 ͚f�(�32�"�&���w3M�Ys�7���w�w4��d�GWQ#��̈́`���5���SDk)V�w�{���!MQ{`c{Y���Y�Z�;IG�ѸL%��ZIf����x $�PҒ��h�t�,+#"�Ze��Ǎ\WkN֔ɑt6�\�;˒u��Y��p�Y��T�j��q\���M�����j�x��-�d"��d�������qR
!�m\��V!�8�-,M��mb`֘ڭ���OF��շ��(|�}�T`n�,��(�J�-&���+h�\"�Lb�P	�L9u�hi�w(Z�}�)!AJ��9
v�JGbD�B�yu�y�5z��V��i(��!Sh��%͌\"���z~4+F��@�bN��ֆ���Z�Ue��+�����[��L[�T)���'��w@͍���5�e�k�|@�+l��y�!Cu�ÙI�,��.0��75'�8^P��Ʒ��
�wB�L��6���[.�Gu�(�l�՚�Gq�z!gC��Ǭ�+G��3/.�TH ����;)�wR6(DӚ����uuv�Y�()�Mk�����(�9�$��m�ڎ�]��kp�tz��r�KrL�oFk{x��V�f,��wSr���ϥ@M�٪r��d�$�ue!���m�=���b�0��N�F�iGihw!ob�x��۱�îg�:I���A�G�b����, M)E�o4G��Ի� ��[dh:X��X_-QT��ԇ�H�N��6�^���qy��-���[�[��EOF̏�(m����D0e=oPx�%�����;ۢ���VUk��`�/1�.���!�Cy&VZr��z5`���#ux��'M�pB�?DAK��]�j���7����=zr��GF#o�)�v���h�`���օ��u)9��	κ�f_5t{�����i������V���$���91��^�U5Қs	Yw�-�a�N��[���ְ<��h8i|�X�i
t��yI5��T�h��4&Э4체�[U�J�6CQ�[��,��[�kz0L�F�\
]n6F`�獢8�sr��:��T��
%��M?�n芌F!>��;�2�y�P0��K�&`z$FfA���� *�]T��qj� �_¶O�#Z�h��S�E��H��ؤ��|T��[[ʂ�%6G��DeG���T`���1I�����*d$�7L2�2�˳/%Zb���^�)kd�D��ƭV|�M�AVR�JE(�մ�K�	���Z��m6q[v�SJ��#7F���v�݁Q�^Sl��#cŖ-(6õuusj2�]G �F�^�jD�����T���VŴ��*&]�׷%��t��q'[�b��Y���n��07�n 	�l�
T*��n��+
�PR�X�Ilɮ�����X�����L��.�<�70F�xmk�k�L�ݘ"����M���sh>�X3c5�*v0=��f�h���)�R�2�I�	�(�,�T)�19(P�2ɤ]\$l��
D(u��o~�K�v�hW��`.l����������4o�rĂm�ōAVg�-P�N��j��2�ys/X�M��u�Ѹ+��L��I�����@ᗓ�+`�+�y�Ϊ9��Jա���؁N7NFڋ.�4[&�6�fg�'��d���f���+�=�{�x|D�Py��F,\��M���6�AR��Q5_����ߺI$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I)$�I$�I$�K�ܝ�*Hv�6�JϬ�e�BM�K�����[����q�<�X����+f�)�xD]�;�������]����hԍJ��]���P.���H_t�2�N�<gxk��{F��˼%F�7ښW5�Ick�g/sVγ3�F�d\j����Y��y��olI����wk:�ؖ���-D����r��i�b��C�ڴ�����j�̀�wH��2Lr�m<6f�|~��ൺ\�A���L���N�k��y�Jj-�}9n֋in.�i� ��®�W�sbڄ��hM�4���^m��=y`��[��C7J��&.����oMü)4R9��2�u�}G�L�\3e!������[��B̏1I��0�T��b�d�1f�ԛU(u���T˷�u�*MVR\�.S;%�ۓ~z:�dX����t�忂�f�Q;�O�;��m�6�)q}hs'S�
�쾺�fdMp�PLT�����8�	3r).˺�<��l��J�̢�T�t����.i����%5|�W��'Mf�D��֛�[��ʗ&%4���7x7^W���i�ƒM�l�0�699M��U�aJ�(�Q�bs*+���ym��}'n�G;���n�_)�/^�Dy�EE+8빸�{s8v;a*��L��zU`Y�I)�st�����b����'��٧s&�<�(PZ��:�L!ύ��c��5z�DDL��6�o̴��Ga���aV+3����JS�.%�sY�(q4wdSr��ۻ��B��د�="��G
��������e=Ȱ���1[��cZ���n�H�X4�T1z�[�b�]�X�U���b�<撊��(�ޭǓ�I�)��m��^2��41����A��2ۮ{����w�`�]�]���A�W�w�I��U�s�9z{�3f�;��ZM�8�m='j4�_Β�^Ǧk��^k՚���i��6LHwq�R�3��=}>(�l.�	�J��X+Y��_1��=�V���V�*�.��
��'��<�:ܤ^��:!��o2U�6���֜w�-v_e��I`X�.����oQ�����
W ~������Z}����)��;Y��;a��U�&UJ3��`4�Ո�(�tɖ�5�����Am�9���^�zU�-b�A��z��V�[�a)ۚX��kq'��{�z�hw�Cv�&���VB�y���NcQ��A�:��ܕ��;f�y�N6��`�̖���h��J���ؤY��¢�ʾ+�n0�دr�'DU�|0�3t�(��f��*�+ZU�&�hX�V�g�E=���y�n� �������n��r�+b;Ģ���5JU���Z�@���|��V7v�)�V�Z�th��P� ��Hj�ϧ���p��W���õYZ*֫1.�/Q�����)[�Z̫�[U��;�󫒡Je��Q��0�>4����WS��V����)��yrR
��R��[k�ˮ��@�a칒�l��6_9g��,��qK�
2��mɖ��=Ev��Mm�'�K���ڮ�rJ��l^	���j퇵�犛��&�<�iX��L/�W%$Vm���2!��Seb�1��rs���Yz����E�/hȅ���
�ά�B��1�l��N,1��"���2�*As38��	�_	���c�F�z�:�J�k�y�)�_KZ��/W�^^-�Ĭ#2��q�7_o]������5W���"���W����hQ��&�W�T���]�dEi���l�eu��o+�魋s��ۍ"�8� �Nt�Pb����\&"��ƶ¤Vq�=[���/�1�օ���D�;(7J���C�v3~h�%˭k�Zǃ{�@�!G��Ė6���ӕ �vV\�n���
���?�[}����G!�V���B�ޗ|��*@y]!��mc+d��'�\��U�i�b�o��iv���<+��O�$d��8�|���Fhcc����)�|�[�X��L�1r�6�݆u;hU��$Ty�{Xgn���U���b��V_^��Ms��%�ɜ��Zᘷ��|2�U荃@TG�hh�n�
�Y6�v�n=�;EC��-I:=jPҺΑ�]	�����ڛVd��y��[�*}%vAy�8� +{�sS���h�.�Cf��L۲k�;4,ϋ}�x��A��*s"y{��ʺ�����щ�u�ys���`�|Mq]�N�	gRos~�Tk:��"��kP���e�4a[̮0<����<�����5�;X��)iz��77�RpXf�q"��ʥ��!��� ֤��]��TIw:�lɓ���_\���T�s��Z�뷖ǣ@���_ mVrV���w$\���DFPmš<������Y��ݫ�u;s�d�H�TC�����{sz�59�2���s�]FζQ��yל$ ^Sc��¥�U��/�S�Y�D.����^2�iH1���ױ��X��Cv�X��b�VX���ޕ�ݠ�Ut��O��7s�
]EK�3cX����ύ�U�z�se15ky����x��,�������Ԥ�rQ7���GsG��S��o3^�V&�zT���f���*�c��خb(8���v.�Ig����c���iضV�̠0A�S~�B���s�VC��Hnɶ@�.�/�;�R���舺X�*�{R �ٱZU���X��>-���7��a�.�	�2?�A*�c�\ܒ��&;��R"z�,�N�V����S�a\.�~�-���+^�z����K����ս��z)�hAh'���n�`��5��gvJ�vn�c3M���c�3eN���u;Wb͗Q��HWH)�������S�͘ f��Ve:�vX�ZL���Q��t�rk�VK*�G�v ����=yhS���x�kGe���j�M��`�ܷ[�Tɭ����
+�äE�"��zE&�0�����,"H{F��^��԰����ϓ�*�H����\V�wcK8e��b��˔��=�h��d�3TҭZ����Yƴ��S�P���(ژ����; Ʋќ���)�nm�"�B�jm:��J�<��1gg�Ceqq���+ɥ����U㤯���;vf��\y88E����n��b�{OY\��ҙ�q�աJC���4$�k]�yN�*��N	�Q-�$�!�ZgE+B��%]����B��15��F��9m͡g���-����}3�M6�m�y,ñ�Q��a���m<���oW��k�=]�Q�D4�@�cY1������&Y@�e�e @�rݥ�*Ǵ䡸�����LZ��-��9^ۛ
�:�E�D��_jB�tڧ�d�l��G#�Ն�"�Zʲ� �`�«y]M�jU��k��� �����sl����'R��n����|Jg(���Õ��8��U�1�Is����L빚C*���*=�OP�tH%vȕ�[��\jH'3jt��Q�e��3�)���ܪfM�݋˒�p]L��ޠ���zhT4�O��[��l��ɹ�u�Nb���K{��;ĜLlΕ�L������%3���G:!�Z�,jj�w2B�v7HYg�m�s���^��[{J�z��n��x���r����ٔ�����W�k���Z-�R�l�}�F�۴;���Sk���e��	5c�ub�T1ڵz�ɺ���\ٜOt�e
��Ap<�Pf�q��ܨ�5Bs��4V@�c�2w!gdbP�2,�pB�Wk�� >�=|��};�L��wg;2���ʐ���J
*�2$ڼ�/Vt综��!]�&�yE؊��!y�K�`�]�T�ɵ��;�X�͠��xh�Y��T��V���}w��!���J�9$;ӢȘ60��]��89��Z�ި�쇤�N�H�	L�#�t��䀩��o�7��!��j�L���k ����)p��Ѕ�=���Y�t[��i��w5�2�Օ���t���d<4	���3���M��`�j���[Ɣ��N˸:�튗q�b�ңjK��*{��t�OH"��F�¾�/`���׹�I����eG#&-]�WW
�"{[�Vj�w΋=���CqW_T��q����oBv�=���w����.� �
���\�yƖNV@4k���������{vm̾����Z�̨�en�]1*d%�ސa�AR�g9˯����5�gu�=��"�ܡ��.4��L@�r�TQ���T�����d���[�9�����*F~2j�7ƙ���r2���ef1A�R���@�1�SdȪ�=�^������&D�s�u2���f���撂��e3�,t}�&ol�~k��i�]�+�`��|��t�ڳӲ�d$t�s�T�*7�Q�iְ����T�uܳ�����c&�)]�^�F���`]���"=�Z����V��hwi�ن`��bݺ�]\��+��YV��<���EYzsr�qtږ��IN��Mtq3��{qsk)���2���ԋw�q�"A+�	g��٩���ũU�D�����ҁD�w9��J��=Ԯ��7�ƹC�'����O!�½ib�v�V�BSy�]���d�P�q�%M7�&���YڛKO�z7{�-f�8k E�2 /f2�B��ItN�.��Y��1�9��%t�k"�X� �͌@�]m��mw�f�wa/��b�IV��_�(>�ԺqcnK���h�0���謼�x�=-�5yR�Zy,h.�9-<��ɤ����*<Y�	#Jjnu+���XPZu�0�a�O=
�	{DXT�l�m��}R��ߤD���4��`�n����� �^�g/��U��,I�[�Q�Ěo+�-�7.��F67*.�Ⱦp�����Qs;���%�n��Yƚ5������"b�Z�tީ*1�e9KOذ�I��1-981ֲ7]�7����K7BORe*�;�9���+r�8�-�ۂ���w@��Η0��^tJ�͕��8�v�C�݌ts6�"�����;+�޾w�fd�Y)7�,��Bi���_N�N��rKթ�{F��][��Y ��c�Ӗ��J�Nr���C�
�v�F2�nMh�ug���ܜu�2�Z��vm(�vl����q�.�ڄ��*ɺ�Ų��Z9Q���t�d���·��=�G���ꚬi�=j*x��+�j��ˬ<�v�I����X������vC�2H��jq�|�ިAXt;�QE�VRj�δ�F]t�q�;4��M��;�=�1V�z���Jʖs3�n+u52�,�����eL����A�kh}�_9�	9�Fw�1P)���o�5ed�/�FQ��fG܁� �v��̇��⹇�J�o����X5�k}���R�aY*��ҵ��5����mS�h��1��ik��OGm3n�8�K*���m�y�O^��8� 헺��-���҃�2�����Rѱ
��5o��Z���.2B7�t��7�Llʅd��9f��̂�0���TSF�����Z+]��>W�%T�K]!���G6�G���3)�O�o6�&��MD7��w�6Pt&2���"�;CV��i��s�]�}��]��a)���^�u�a�Ǽ�Q���EO��3���e�
��9��6%x�G����,��h�-���)��^��֖�E�=�\��3�պ�ml�cɷ:Yg��C֖<��J�33�m�๩:��D�J��P@zc�F�*��9��Q��\�%ggF��z�����,ݾ#)��� =�r�����{���d����7O.�+rӌ�mr��D�7�ۛ3�H�(Du��N��EcmG��d�}7ޞ+̓���xC�H��Y���M�ٯo�h���9pO��W��[Ǝ���F���ҳk�&vǛX��uI��β�EG�y�mN�wesf���:�>�{���n�{�µ�cҪ�4Y�s�S��ܗQ��
��R� �7j���NZT�ehX&T��3�-�功4�ܣ%҅ͨ��G#�5)V�HwdNwLɜ�N\� �I9�m��jf^Α\3麭^jn	�TsLS��K�ݠs/D[&�>���g$�V
�VG9ʗ9��NI*Q��K�f޹�ԟ�E!1:���A葽_S8��%�s"r���yt�S!F�v:���ݩ#�X|{X[�5���e�V�ITmCNݮ{C��@%G/v}�*��n-��M�w�L]��z��T��xVL퍥��CC*��l^��r�㦩Ȧ�]����p�u3t�U�TԯJqG����2\�0FN�n����3y)6jw>�9�ԑ9�I.�9K�LN�ܒI$�I$�����?���������v/�QD@]�
V�X�|Q:3Qz�3Ӯ#ev^k^��M���ª���D6T�Q=9�q��:�C�n)JQ4p�}��g��gfޙqH�U�\H�ˉ�l�Ǚ���9�sw��,m��wi��7%��]�|����wYT�X2�^r)�W
��jEX-0.p�ז
��1�U�J#&>�pI��T\�6/B�eKj���0�ù�-�WCyqŜ��kK,Q�p0�:�4A�4m��r��%�渭1�/p]c�N6����=|B��ijT]u.��R�ku�xܴwB��.�]̡k�W��z;(� ���qA���S���g<yP����Q�W�4v;��R.�9�d��M.N��_��$�s*���=8(E�O_�|^�vu��p=�&Wf_,F�h��xK��	1�)tcn^�c���W=]�;_��{�U���y,���ڙ/2�U��Un����]q��.5�K���k��h�P�4R{-@QIEFj�I��$/%d���DG���P��+��R�Q;]��1b��+'w2*�.��E�b�.�Y�K+����N�ū�X����.٣AX�\l�n�}�r{|��TP;�ʔV�Ea��d)P��eì;�O��ܒ����4﷦��%VP��~���e���Ǩ�%��>�,ܳ�x܌�6����zO]�yfuPf#M�
��[�YzWd���ԻZ�4�c[̆�=����l�A2>
����%F���d� �%glV#kc�ځ M�j2�P$���^�F��k�j�+�GY�����T���>�l��t�j���3S�|��-��y+�$�^kg�\z�d'eV����h��;p��άʶ�~��%N�@s;o�ӹI0nM�Vu�w�:���ӱJJM�p�mн��ʰ�*��%R	��r�te[���M��1`XH�L�R��qk��]p��5�"�Ӆ��hջ�|�w=������k)5nr����O����f/��׳N�'���;_B6�t�ɕtz�����k]�t��#��^�u:;n��<;�3d}��y���1ªs�����3��j���bcU�n�ڙ�D汙N�|��om
׳�W1P�si�J�:�;6�+�m��Fɮ�â��<�����HӐҦ�m��]EY֯�4<ˎVlʶ�K��P��Y�pΖh=ڔ	� 9o(�ge�wE�q�.�/AM�X~�9o*j<{{0;����Hsg��ZS	��v��S�S@#���PHb�S"2n\�i���n�|��S�M�y;&wom	B�&�������֕vP�Rv6e�9C|f2���tҔF��;݂�/3m���s]ö�Z��&�X��Mr9]�r�tΥ�J�1V�Ѭ|렳���t���v9R��q������4��i5�(�R`'%]橑-���/���7��d
�V�%E\fs�VT}}O6�X�*٨T��ӳ�q��h����ܥf�X�S����	���Em,T1��s�	��u솴�J[ �C�����:"��%5\6�������I��V����T��gn��t�̣�%�w���j%�2Yq�u���|�j���M±���-�K(tR�i��c8|̈́�7���օغv�󥯠Y�6�����:��bJ}j����ڎ�k��|*K�Y�k��pMv)�ں�Y����M�;{ ��u㩙ըR2t�j�9EX|�L่b�'f���w|�:;��%[)��0+����%�\��|'I�ۏ6�����J��QYe��=xx��U8�VVr�������ê����[��۹9g:�qⰏS��ۑ��S*�N��E�a2��e�\�v�.�F]�@L��ڼݩ��I�w:<���������Z$���R��Bmƛ���J֫y��������iv��<Y�tZQ�R=�wwbܾ�?f�(nG���ohz��K�}�]�dB�˚0�{,)�Z㕸$I�WC�5H�(�w�'2ɰD�9��V��E��6��qJ�0_KI�qRQ �_7*Fh��8W-X��*w6G/�(.��b;�(���Sx|=b��KJ�=�\桊��o�7s�|��KqPX:q'��p�&ёVgnNjȡ��1�1p�����9,����gr�K+<W\����l=���J�ɪ#)�����9�XTT^c�b��lT,�V:��X:Ӳ��	�!8�J��J��ݏ&ԏ��!�����4Xܩ����w��`yiԅ��r�����
+.�2��j��=· eWy�!E�Y9ެ��)#/��)�i�u[Oc9����������
�rZY�]>G_ ��4WT�_�v���RtF7��.b9��{R�(���m��%�˦�'U��ִL��Lu5��KkB�]�jƹ\9�d��M�XaG�9+-={@�R�9�ggb�F�=p�k��CND)컍p�9�K�A�}w\�bJ�v�L��X$%��s��H�C��vm��򳍡H�]�ң�]�Q������ΓQ̽ڽ��vE��H�D�[2�ݎ��2�t	Ґ��o<<����uҕGy/J[i�#��9��S�ŅQ+�.w�t���2��3��s$0�S�V�j�E��k\�ꔉy���J���@�rMK�	+,�֥#	��--�l�y�-��BE�"w����#�"��U�)w[f����r��$ӱ}�$�>��r4�z�V�c#�wbǥj��Z��J����OZ啕0���b�����pHc�[4S�%����h2�e�7�����pX<%��tRzffLWJ�T*,���O]��wud̊�㫏�=9�/b��۔S��% :�j��oLW��������_����nGw�9Jh���_E(>T��
���y���<΋�[wB63h��Z$��V�;U����'k5�l7/�x��Օx�I��Ya�u�O\J�Hi�U�n�:G�1]C\^IFƥ�6��nd��F����*���ݲ+qW*U������nrQJ%��y���k�z�*�5��!�u�ʳ%�X���Pu8�*���v]*z9��\6�z^����oPoz�K�u����u���5G5-��b�Np:�-;x�[h.��g'+��PI��ի�)�KC���u�n��8ԩ�[�2l�������-GOt=;]�������(�ܣj΄=ʳ��E���˘`��<��K^Ӝ;5��|�Ȇw[[���%����Ag%���޽����8�fݩF�Y9P_�t��)]�`啫wb�5#Ɠ�+�ޙWg�n�bY�WV񜨫�-�l.R�@�S	��jé�iJ6�c�Ng)��9
�õ%.n������;��YX�t�ν+ n�2��СBw�ѳ���.�X}uG�NrGH�̥�,���yPX��<7��i�v�Zn뱳zV]a��M���G����uE�$�71����=µhâ�� q|T��n��˨�A-����7[�h��ѩ��/a
o%-gF�X�g8Ê�uE�4�(����5���I+��`k�k6��iށ\��ڶ�k�������ã#RZ|Ѻ�mi�ؖ��I�N���j�Iu��t��>��:�W�֝d���v�歡��.�t�`��� p��u*��F�Z�;X�aR��\��fi="V��X�6i
-��̩e+aa��KW�9PI�(
�|0f�Z��rp���(�e�o�V;�w��3\����;e5+�
��GXx^�[`Pr"{�&��e*�Ȯ�+���ĳ�KN�}�Y-����k��ݡ���#\з.Y8\A������v��Mɠe
,��� ��ΖE�p�+���՗��%��٩4�K<U�����'N��I�S��wu�IB#Z�m�C./�����Xޭ�V�.���j䔶���,j���6�݄�i;Z.p�2���OD>y˓Px�q\�����ɯ�d�K�ڧc|hЬ�P1,�,_B���B���EL��W9���8�OTWm��'j��| wWC6�t�GiO��@o�Y�K#y����P@E���Ͳ��q��H�G
���t.�*�v�qN���,���ۣ��yt��ZU *ϪB��t�Ƕ��U����6�8H�4%��Y2@8�1m�����˨�Mi>��e�[TVJ�8_L�l�si1`�|��oy�Nc��i}+��2��]m�`���Lٱ�9tDCv�B�h�y-��I�:�y�(<F��w�t7#��b��f������#B��/C(V1�؇5h�x��ʀQks�7�8f�W`ʼ�]-t;sv;I]�S*�j��X� 1�f�8�|Hr_)��&tUY��x���5l�M6����6!U��sX-�����[����]Y��U�`t&Dɹ k��e�bꕴʫO-��+{p�yZ]u�j�#a��g�{j�.Nˉ�t��u�����SC* U�略t�lAb� /K�k!LY����@%���9�����͘��;���9�|^it�Za�H��+O!��$�@F:�@$]_-Z���.
���γE�j��
��KћL�B��ng=SyZ��F����lu��*�b�y��RR��Yei���Zb:��@�n����ңKlP�����Tf(�aA1Sfwa�W]���.V"�c�9���Wp�h+�଼u��7)���똛c��-�i�s��BI���e
{Cd5�m)$0�1h��mk�v�&�8i�{�Y���NQ��@�lV`;F&��ި�Ⱦ8�3�N�;m�}+6n �y T��s@�Tu9��w.��]r*�gq����� p��A��mWX�:P&����8j�ٕ��z�Y���rpQ����óo�=����v�<�:����=ґQ��k:jjݾx�n�� #h�6���9�p�ܴ�o.�wy)�� �NJ����l�]!W͑"��Z+Ov��F�Vؕ��ýZ�>c*$Im�`��U���w�W7j�֖�N�[���5��w�U��w�0��7�C���4om�Yo�=!�I:e��a�'2�zN��ԩl��Gay[�OQz�q���'L��k;yyIMLc��vo]��;��:4@��J���e��)��v&0rv�Y�5R�!U.B~/��U�ӾǶ����urli`��.���=Q�$�e���P��m��µ�y݁��}Ϛ�����
9�46x賙�ɽ�\��@CB��]HF?b�̆�qھrn�����T���m؆��ǜj�B{j��Hs��r-�9OU.�*����O�� ���P�Pj,�9@L[ó8�3t>��6�[�]:.�t5­�ը��D"[ǻ���;��	�$R������$N�l�����ʝYn�e�����\Y�U�{U	�jbuN���1�T2���˺��@-�&�i�Ek�q-���є�Ѳ�k�2�s8�ٜ:�^������J|	�y�#N��B�q�P�������A.vb�}KFW.k����y��Q�wQ����BggK+��S׷��#Q���rl���H�Szf��k���2��%D�v�-�n�a�:ڌ�+@�G�V�� ���+sV�ƣ����bs�fW}�k(���Q�J�)}��(�^)m���I���)��>�Jw]bT��k�Ҋ������Jt��8���!j��&]�v�[�1�0�K\H��L;�kt�3#7�q�rZ�=���H��P�O�s2�yZY�)0oP.�^ѧ�f�2qw:iwHKKTul��cOg7k �`��y��YgA��t��z�#wk��1WX���@&u�+4�r)����<,n���'ub1�ozS�m
Bf�wZL�yF��q�w/M���2'9��J���bB��\wA�3���ء+�Z,��w�,m�XX:�Pzج�٭�֬NU��!���Z��)i��U�;���6���k�{�{���I��se.��+8���Q�v���\Ų��"����%:�ojD�i)h����4h���͖hϹG�����F��v��җ#�L���Z�u�Ơ�*T��j�,ݫ'lG��`H�읥�,uBrq7zqpté�**��.��}Z���'X��^����ΕA���j�N�U�k$}�v�J��̝ƹ,iVP��|;r]��p���'���������u�Gp]��%l7�sJz���D�S��;�T̗X�T�t2;"9��+��J�x������$If�X���F�@��g]��:���VV\=a��;��nT&�R�31�{w(Z���9G;L<�*x/��:֧_b�������\D���2���ᴭj颟*�qv�88z�:W]m�W2VL�[O]��r���o�~L|%M9�kE�W���nIZ�Ρ�"�A��.��E�xw��<:>�K߻7��I$�n�T;0���elɱ�9�i� F+2�':�1Nո��p�m	v�v�&c���B�tqE���(���!�]F��rG�Sӵ��R����EB�w�n�dJɚ�WL�hD�z�1���2tR��"Q�%qQ�0ѮS��8��(�R���^R�w����y��~㦼��5~��a�W����eg�H��F�,r���ۊ�5���3�Dn-�B�!�1�'���Z��Kq���9�坹��bz�/��ɳ5)5Z���R��Q��{g�E�6zĕ3�3��/�d�2W`�×�-՜[pX�J����յD�aN��%�s��Y;*+$��͗Ύ���)���}؆N�Mi���ˤ�>�Fꛕ�a��.��wR�[���o>��R�$�;tfϤC�
�������<"�r̰2>�������仚(��^X7�BTf�Ǚ�;��f�1b3�@�y[fLv�;�ȉɡ��Y�z��j�7S��Ҳ�H�L��.t�Y{����������g�a���6�m٭Ф�|�|3�,�N���Asw&ů�`��ݓ�L�ZIC�tˆ�궞JT��r��oR��&�Ùֻ����f�[kC�L�ڒt(Ul���d5.����(.�̬KWs�^M������}����$ڠ�E,
)Rc<�12�"�>�c�T��(����EX�%MZ��(*�dYıU"��ƅU�J�
,\k�y�6��L�v�R�d���(�
T����	"�*Ŋ�I���A��(Ȳ,"�(,dXJʬR5���	�*�P�*�*���H�E�Ƣ��3Ԭ�Z:�P�:|͠b"�r��!�g�j���T��?Z
�ДB-IDQ�=f��>Sl��#�Vى���4�d�&�̬PX�(�VL|J�0� �q��+hT��������V`��dG�M'��Qa�M3�I*O6镀hq�±a�b��m"����U�ji c
�Xi��L�?�n�qUZ���j��5�W<6dg��#ӓ�p�BfZ�F�Z�&�R��ṙ33ui��c���6�UnɳQ{)1�?���;�-��b꤫"�zꍶ��td�dT/ܯJbR[��]W}��؝���U���]CHu��^�8yC��+̊o+V>�0�b�-�}�kЅ���c���Hj0k��Ex�hEdg����J#��u�N }��D�9���|*Ծ9�v=�I�^�魆G�D����YT��링����cԔ��\bÐ�͇���`+�>�#��u�p0�@�ʩ}r���cjGsL�w�����!צ�"��^���3�ݪ䪖�:�GD@�B8���r!�b�ʚA�;)���C�(ݧH�[U��^�p��2���7��)r�����uk��=Ƿ{�
:\F�r�~�(��Q�ka���=KAu�ȯ�5/l��=�![���	㔢}ވU�,	S���<��2�_L����̢��iZr�dۤ�\��p2a�D^��:n8G(X�(��Lؘ{70������Yd͋�uk[,��	w������N!���)�56����Y�L*G(>�ݣq��C�>�;ŽD� �N��	[F�㎤�r��uG��clw]FG����M��;ՃȑV8��N�9��v�Wˣe����V������Yq�nE9PqYXcb*T�ΐ�����*�����!B�+��<�oc�X��+�i��JY���S4���%7�.X�i�uz$�L�����vtR(Q~����:���=�ɯ%L옷r��
�׹�V��zvk���
Ol�y�a��y�t0T`�n���#��Fp�Rv�ԭ�,�wv�$�cmI��� ������ײˊ�n '!"'0d��E�PhψW�)�����=;՚� �����԰�yv�k�g��2���8<Ϩ|w���;�|�j/���0hѡ2A��A��>Pm�\4?��
sUp�X���s��R�%x]�O��4��<$�g��g��a�k}A��U�?����n�߲��jm�[�+�Υr}�O�Vw(�ª{^ݙ��隇�0<�u�(�]���=E�v�.̕9�DPԥ��."�ޟO)�q��>� ��o�K���t��ʋ;Ȁ�\<��v���[7���^i��m\����;=��MSM���B�\֩��+��/���D�)5�o�R�΢�0�����Lܷw�j�FN�r5���%uX˝l�|bT�<�v����uh���	���;&��&�J��Dn�O��D�*"�3l)�)Q��Yр6��y�^4��޴91q��ẒȾ�CI� qɥ4:��������U��l�Q���Ocr�y�����H��7P��3�돉F�@�0�x�k�>Y��U�l�Z��yݵB���6�q8���^��f�\q��eW@G�qo����\�b�ձ�e��a��Z�kjp�a)f)��Xgb(:�ѱt��q�,Ż��O`"�q�8��J�%�8{��6)K"	�,�f$4�q�ƨA��w���<szT6��]k��Y����T�dn���p�,�t���f^(��tFJf�Yy�/.Ȩ��FB62U)�ʟdH���c2�b.۠	`�\]0q��W8�d]�ViZ�C��7fa�,h�$����'��y�3~��jv�|��mu�wNVQ4&j�O#ob�:�l�,�q��D��!�z;�
t9*�~\/���i�e��]��������/����]������c*R�M�-T[��1*���R�'��(Q�R���4����P5��}h�MU���W@�iAC�E��|���)�-ΥM[�fn���%�2-�	�Wz��ev79��{�V��|S� �T�hM��
>��}cXnMFlP�8F�c�BQ�+ZYh$mt6��6p�]��D��{�=�J 6��[�0�V
OX�o�rH�2\���l���t o�ҍy:�<B#7�e#�0F�=�]����Ƽ�yf�qН� O�o����8!6jR0��7#TP�T��s�i�۠�˭���Bܝ�})�eⱯ���wy���h�F
O�(�`O��#2<��af��v �<��Ҝ�wh��F8�&�H��P�}�+��Ģxfժ�>P����Vy3 i��{݊e���������i����z���b"PuQ/C�����}���N�����4Ez�[�A68f�5ok��(Y�#Lo�z���B����!�u�_Mƍ���7��0��S6%M�^���c��#J*Գ[N�ٛ�S�F!���.'/)��w�j9Y���].#��&���]m׮����b����/z���nza�_4�8�(����d�3���y�{� n]֌�zZ/�{���b�r;�Myu ����dyq�kP�d�R��.�=�4�[ҷŮd1egl�5�ܲE+�U�)�$F�v7G%�C�Տ0WS���<�5�K��o��i���Fj�{��'e),��a�P�/%d�jEqŎ�a�nv�wB��]����Kk/�:����`V��?�B�k���^����/�>��i�o>����0b=�I����k(�Ӷ%dH�P�㭽ͣv��A�܎}���c0��rX|S:9Squ/��p����Q�2��Ix��8�W�\���29�؉I�Ѫ���j��xkz������㳛�y2��Ĭ���]45����V���2tw#���L������IH�8O���]��yr��z
�Z�su�ی��فVvj�ʩ���%��}��_n�1)�k=R�����(�z�D�ՠ��o��-+��kS}�^�ߕ�'ј�rt	�RM��*w1�NgE���:,��]$�K��������8w��hK�n#�X�o0�t�WY�o�G�T؊����:��",�ή��F���9v���Ե�l���G+�EJ�}�v}7�v�"{�e��j[nu�T�5�����T�������0̣b�P؄���z�\�D���6':�'#�U�k'Jw)�Y�5i]s\��:ƴ���'�8N�������t��)���El���;W�J��O=�j9��4����4���z�&�JҤ���.��t�u���W٪�j^��D�V�s\q���]��y23�����+&�)�����Ō��iT���4by۷L7��t��RL�!�æjV���ӉP�;m{ث�5��g���>��b�=�J�HL/_A�U�i�t^T��FjvBM���X2���Cc���K{�雩b�|�5+���]#��Ƈ���J�m�ȑX�="-����F�&�M;[�agG>��X�Շ�1�w\�/B�rv��(����En��lDE!>>;�G�>�v0�/P?'��9!��k)�R�� s/%�<�*�N7��p�� 1�U�6�a����WJ�3J�zn$dy�;mp�&�����¦�Ԓ�ނ��:I4�;�>qr˼�ڽ+%��߮ �I�r<vecwt�� �R�	�E%Y.5�bJS��,��O$܃�������'�����"y����d,���Pv-��8p��*xH����G������[{O��R�'`�j�]�{�nGX�������yKo-=a#��>���n���U���:؝}X��T�� ��ƢMݬW|�wCL)�bo�5�甭T�CoU�{�n�)�j�Bu4_Ff.|N:]l��X��)�I����5�yoC�����8m#�dD^�,v���Ɇ�!�3!�%��ǠUs��Y��_��f�*���k347�MN&v;�8�e�G���>�WG��0���{����̼#n�FB]���y�y�ܘ���6�+�ƙ��!3�GC�!^z�P4���#������N�T�޾�j��!ZsBrX��ZCŇL���9
&���l�,�nE*�r�J�-�t��Ru�2����J����9���R����بq���Z��V4gN��u�Q<h��5Z�M�da����h�������u��Z1�$=�Ԙ/�!p5ڵ2͹@�.�4\�$�f�rދx�M��X� �lYF�w�a��P�is]-s�f�v�j1̝�\=^N�EW]����u�{>0�p�y�������sQr��ɛ����p�6�dMb�uX;�o(S�ӕ��Se)Ҭ4�A��(0����edH�St�ڃ�Ku��U�e�h�E3M�)��he�.����	�[w����+-������Z|������n�y�{�+|&X�p��^�|�I�ew��l�����Y�\�F%[�`7�s|�Ǳ#�^��k����{M�ZyK���Yp��+�~9>^�eN��%y�/tP5xm�l�H���|�62g٦���3^�S�Uk��Hј�y��W6�_ ���Y�ü�&�([�ٱ=3Hl�L��F��ܽ�T�gD%�l'{�i�\��u��fݩ)B�ph���H���&k�9�·}Vū�1�bAa7[Ϯz0�{�uXq$y;��x�S�zuI8E�p����vG㷛/��.�W��M�	}�]�YB����Tռ0�2���1�Щ��,E[jƬjgX�ƞD�T�	eC{������ْoö�g��#�K��W̦�r8�w����q�;X�����G/�l,ٚ��ͪ�WK�2�#��$fڵx�W�U<�ࣝcfל�xC77�3����MMj���ܟ
�e�ӝ��f�i��ڊ�A�vc$ӻ����6�j�1�/��d��V�v��Yu�mZ�Q	]���rSX��d�q{/WY��=R
���)���%e�WT1�ס�q&�j&�9���~f����L\��:q>ReW3�5�p��y�oy�s*S{�{�l�K�c���'t�(���:q>Re�3�[�ە����ɸʼ��bT�q��r�D{��C�4r��B��]P��^���V���'���.�U_��>�u)�̙�1����-����5p�bT��N�8C3{?8<�א�=R��B��s�\�Līl����'Q�v'���o^_+���d���;/p�j�ʼ����K�0����X�@�(�Di��'N|%�U���/���������r�V�޾*pa㋟sQu�I�h�4}}jc�ͨr^M��5��F-�z<�#��w��&1lG#�_y T�>�he,�����r��D�j|��e��X�����=�����@��������ùb��'z��ϺV�.�}K4-V��ݛ�U��.{o�/�"��e�O9[�\��GC�����JyS�oz�fõ �-�V�{De(/��e��P�a�3��#BҺ�r�H������gf��gk��W����굑q]����B�i��bUB�O=�`(�`T(�ñ���5bswW1�� �g�G:a��)��>ǔc�ozvr�7��E]�>���%�t���TP�8�������d�s��z��� �-�)^�|��ߪ��ut��W�fC��:dT���jW[IIs{yn��-�15���ﻩ������f,:g�/�&| ~�=�>�I-����_�i�/�ʵ�&�yՏ D�źr�}%b���b�W�f:;� �S8�O�뜇k��yt����Knf+Z8�ki��y�Lu%�&p�%3u���������M���%b���'e�X���cb��r�,R[�]f�N��0%#;����å�ǌ�(�A*Uy�:������Q����b�e���1cǲ2��˗Z���G�6�i����
qJ�3Ƿ3Q��C����2�kua�ʴ�l��o�87����-�(ܝ�����}��z��;+]�uܦ9c-dN��fj���-��;w�S��P�u_<MSAÕ���]�<�-Z'7�Xe̳J�+�G�uꍂW1�dAv�[G0��VN��#�kc�^T�.�����V�ڇV�H��
�Žщ=j�d�7B��eG�w��t2[F!��ڨ�!c�D��2\��rY0��ۋ��J�N��� .�'+nD�r/0ѴJ�-_9J��MM.b��_o�	�F���]�C��0l��z����%IN��Ǹ�-�*{�T;�攒�.�r*���y��t��BB���}��y)���
U�в"%t=�n��ܝ�S��K���b��ܱ)�BS�&GFʭ�Х������5:��"�u�]�4;0�I��vt�&�F��u���)Z���V��-W��k�?���I$�IA���XUDΌ��r�D��Y�w��M���Qt]����W\͘.��H�հ+I��9foS�iY���f��l5w�k�*/����s������Ģ/���5�O��-��UˏGV���C�$�<&�y���`IG^�x"��.��p���G�ڻE7�r�Ǜ5X`�ِKI^�y6;�F�k�>}�$ף�7�
f_`�C��qT*Y�i��EN�h�'n=T����M��v��V䡸m�,���c{���r��G����s�s�l�b�*����\��3em���]�6�;��bM�\����+4�*�j�Z�.��X��v�g$�QM�u���mAw��Zgfn�-�'�`ި)���,�󬛻w�5Ig0�y��7���{,��ա���^Nrr�Ѯ�B�/�3]�Z�
|�E(�����.:�L��X��,<�i��w;piy�i6�V=��)��%��pY��K*�Q|��g�CB����o�wp(e��r�d��T3�Ǌ��[� �~~iHW��FmL����,��~lY��I�w\��T�Sq5��g3#��O�|�%��
y��;�����L�ާ��x�Z[qa̅�H�.ԭU�nU��{W5&���(����ȧ�A��6��
H,����T%g���%`c1 ��(�H���!��,��R
I�+Xa�Q"ŀ�i
�X��n�N!PX��q�(
�!Xo��ɪ2�~|d�&�x�1��2:�)�4��(��] .�V�[i��%Irȡ�d��T*�J��P"��|aXm!�|M��Ȍ��`�X
���E��bcY�\�6�F++
�XO̞3N�6��x�Ev¸�L`i���7O-�3I�1����C�B� �ۊ�#�����ȡa�+4�d�,�Ð�?���{��~��F������*#-f�䥔n� �p�A��#�M{. Nؗ[p�;>��R(��Yõ,Qi0����nb�g��"�ϰ}��H0�k����:p��[�ĩ����|������+�����X"-�����4~�P���Q���������3'��R���?�8\'��zޯm����Ϙ���]��Q���k�ߕ����6<�����]yr���uJMl�3vwiU^�[v����1>��5�fM���+��g6�{��&���U7f��u����>�����V��)�ߑ�W�y�{�*�=����.W���yy�9�_8I�^$(�<�����Z��I^�"���1��	R8�z�N3������I	��g5��+U<���a�ݑ�*:�m�]m�=�w����g�|�(,u��vH�6�� �Hд��O,�+b���Q��z�Oݪ���>���;:�����Z�%OÍ��B��;w-��`Wǩ������y�%ň|�WoLt4�M4����e��R�f/�59z�ڊ�;��1I�FL���PM�4m��Y]5#�^�����vǿ#��(�	3�k���R�f�fJ|�h-�}�w�]��F�c���T!��(u�:��'���'<�97�jO}�5�^*	uEbg;�B#ah�z�ɴeU�C�j�k�;�G�~���;R��}/j$̅�9�,�V��j�����gϺ���C���Ϯ~�+C}���S����f���WV�r�B�h���F���O�>��㊆f:�L7�!�o���+�S̝R��T��]�ˡ�����r�+[:����4ܘ��q=O9$�|0�L&n�/�HRe�A��[���&�H�m�j�JV�QJ���z���xn��\~���)��<���]�R�6^NMC��������⃍�}S�y�>h~�Ą�47sA�0(����'���ɣ��9�������T���X�e�#X�Z1*�;����e�mv�sQՐ�*���p�˅�|���0�ҵW7�L�Q�$=���	��B�ܻb�:�X|@q�<U.�Z������?�����1�K�ǟv��*i�7q��1�XL������6�@9k�;�P��2з�5�üE��L|�{:�6�k諭��ۺۃ�ݱ	���8�U���������X�����^�ltu��9�N����3�Ci�����G)Wd�c.�dƻ�[��s��q�˩0��̀�&��qߣ�t�O�Wϼ���g�q���#A������i�m-��O����Xm�ͻR
P�×Z^Lv��c&z��s���ͻ)6����Ԏ[��~�8�l9 �G
�UvB��������ę>��axvǾߺN��/=��ϱ�3k�n��Y���3�YՋ�'�z��<6{'ԥ�:�vӵ���:%�F�1�w�����ܢ�!%���=l�YC�z�����B���HĶ-��ac����N�굔�O�&q2�:dT�����]{�D��&��9}�cɧ�-�3�3iwS�@�N$)2���"��e��g5	�'���nm׮�%Y�s�%�v+~ɖ����Et�T�H+6�"0u;"�$��q��Í^:�)aڽuw�?h���~+qp^��${ADc�z���C���!�)�Z� �V��� #"�E��%��VdӃ^:�'r>���q�v�mw>��qz����⫐^p���E�B~{ˤ�<���\ˬY�y7�z��������L�G �Mĩ�yju:��摹�]h�^���`���;q4��Kw�3�@ƶ"Rl�F�E(ވ�I��[�k��%�ӼNn�{�.VH�n�\�@e�X����^T�6{шT��\��Y8���2y�b؉�mx��ד�$n4+-{2��Enof�rK
��0���mD����+̜�z��B��N�&TE6������Y~�IE^;[aj�`={�j��x>�����Z*��:o�u��ؐ-�k5��H�O,kz����j|
P���(Of�k9�b��U�\�M��%K���y_�<�Ҋ���V����������p���/��"��z��j�%YZ��'�n�AViY���اi����i�L�|��Bb��yOO�͈��^/�ꑞ9WHT�qQ�_V�j��>�Z*�nY�cs�#+&dh��'J�E�̗R^�k��1>P�̦��{�uc�e�̝+��O]8�YQ��Oa�U�~}�P\����ճ��hN�X��c�ozu��tfkE{S�����gS�MTcw��:%��6
��S[L�uf]7|�b숼p�뵫R�}Oj���5�NT��`�{9];�s�E�OX1�woo-��wK�@J�Jaz��y�Z=0_��c ����U��G���<�n��,RO`�p�GB;��gm���8��.5��t�y�/T0Dn'%��`�r���ǯgl�E�v0�Wy�86\'�.�q��b�[��.�<!nlP��:o���Q��hCO�L�`�X]��U䬚n{.U�?w!�2�]%i�M�?GI��fd��`b���m���`�N'��]��E'��_N����a[������؝}>�sg�O�v>3/o�VO�K��R�z-w�J�M�E9r�k݇>���e�9��o��2[4���_��� %�[�-������2�9J�� ���$_=��Gq��$q����S��v����1�]ͯ�F�Κ��ۙ`=Q��"l���o�{�j�Su��ߖ�v�wf�k`E%�I������h��cR��s�4��C�f�\�Z���\f9��./t�2:��[���cΜ��Hm&r�#i֎j���tWvS�ܜ櫸��v4څ�NA���֋��q��\d_;X��*��	�KĞOe^Ob]��r�X�h�����U�{8�#7��K�~3x����ą<�ژ�cL���S<'���Z�`m`���ؽ�%�����3۔԰�9�/jy&d-!�zŋ��Չ����i��Xsy��Y4���r�j�ﻩ��u �,�ڡ��o3�nyIm�Xtȩ]
�Pj}��2����K��S�1;�[����������B�
�����������Vέ��'N>a9*�k�����˞��qF��p�[�����Ow�����N�~��M�7����Td�mF���N�����q���:�L)ۋE�a�nGi��K+�F-$���rgwzR��jJJ�ns��~�U('�{ÈU��\�����=雔��]�K{m��
s+�G'���c��n����h�A�&<��t-�tg��)�=�]��s�1��;S�.3�1�L�M��T�����GD��7*m;��m��ս����V�X���ݲ��:��F;i�ۚ�_٣j��yܔ�T#��1����|����/���_���u+�y/og"�o���m�H���o�(FL�4Л��W(s:����g$��w�n������q��ڰ��ͅy!5V��c�=Hl��[�I�M��/$��R)ȡ�&�G*n�Cΰ�ݗKJP�Ü#�K�ۊ+>aJ��摴�o�%T-���.���-���8)�Y��d�����:��➠�rkg���[��e{5H�^����C��.n�2]�tu�l�h��学�}a���)֧��@�2*s/.�d�Oą�f)U޷�t& ��>R���M��6b�u��+)˔���͘ks�,1��X��/ ������U���r�I���v�悹s��d}0�d��v!%,��:�1�߄��s!�T.��byC5J����Tezp�+w[�ofj��9�x2��d��)�݉����E������ݺm�uKS})��d9�æ�l^zVO�55�$���O�S��O-.�8��a:�LByC��&UgL��і%dO�'\˭Ü֝�,.=���,ailjO`ӧ�ˮ�Y3{�Hy���g�����W�lJȟV)��X#��,>)����w3'��T���i���Ã*���.�E%"�[�ɑ�lE��$ޞ�]�����<��]+�~�eR��U����r�{-�g"d��I3��|a���	�d�|L[ s9���(kɩB}��y#`l�n:sJ}�����G���o�%�=�U/2v6Q��y���9��e>�f �w3�s�&��^x��Y@S��U� IU�F&il���w�I���]ǰ��̉[�4��Ҙ+G^�=k����K���Rn;�X(��73��wC\�3{�Β���� �s�t���]d���
�u�]�.</V����9M�;Z�SB��������w�+�+]e�B�<nnzN��t�!>�H�k����oSי<���f�뵚�^����D,nv�_�d������ZWC���y"�tvQ��s�m��̘~u���]�_��i���j�*��2Z.*���|Ħ�S�u�i���g����l����C�+����{}[p��7r���ظ�~\�{���QC�8����d���yr%������z*X����o�\��S����fC��:f�n7��k��Pf�uɘ�p�H�q�,��Kr;���O`W�8���j/Ƽɩ�Tŧ7^'9��lJɡ�}H���H0�k�O �Vs�WT�2ٺY�ܙ�Zok��N��$V)��j�E���f��1ܫ܃��:�:u��뇅1{b޴r0��ϓ��]@�4B�0�d���h�2JU;M�o�,;��U՗o�*k�n�z�5�Â�ή����j��r'��\���e�זЭ�eғ9���L��T_�� �I>�@�\��s�	Nc��AIFX]t����y��7R���/����ȭ�8�<Y��� jL�F���5���9�u^J��Ar�U�8�6��u6�{l������f>I��ݯh���|&W��l�#l�I�.�74%Q˱�][�Z�su�V��=ۛ�'_Dk2u�m������RҔ�2��B�x�r�����Z��{������=�H���BB���fr�����υ4&�3��r���:{��ә^|��|��m��Ux����Z,Gd�CdRfE�F��h�ɭO9
�k�:����v��Xm�r�Ǻ;/�֍����1-#�N]�/<]��9���檅� r�Vn;�8ςe��xOC�Z���t�OU�:��z�*T!�W�ef��]��(cdb����~ZSv%[i����D��h.�z���U��8f�N^��]����wu$����˥x�q��k&+��4uL���D$�[�Gd��n���x�v��Az�J�rb(�����z����[���JZ�Y�E���2�<OM5�f��\ۻ�v�>�pT��A�3��
ّ�E!]�#�A�F�nV�K����5S9��)�	�Tާ�l�ͤ���toZv��A��愎����]KW����o/z���9u���gb[F��d���:�_:5Q����L�����"�H�\X(��-H	�3qV�ԣ�[Ht�\�K��]Yf����X�ڽ��7�B����T:j�czm�5�y��-t�N�����D`���J���}lYߘ��<7Ӯ�b}z�����߆ܗl��X!�g�@�\�n��L���ݑؗ!��(E�qv�ӔV�>|���h1Ӑɕ��n����\�	�
KL �]��3PjQ�r�,fh���h:Z*S	l�a7Kݼ6�v4��o���7T�1-�xAGEs��pob�B���I�,u�͊i ��ySwf>�D ��X�Pņ`�*�`,��uIҘ����m3w��F^I�[	����F��NϺ���2�:�]Z�t�<�O,/hT�+�4#LrV�ކ��:��,�A�BG]r�j��6.��8-�Q:��u�uJ���H�e�P\f��1 vu-���~]y�$���I$�B�,�;+�-U�Sk�t�=��R�g:�OV.C�ʕ=Y�����h�N�zڐ��P5�­��T�3g
�4 wH�wQ6��5mי7Zuk�b/&�++��!S39^��7-��K;yJ��%]WyΞ��K+k�w@@D(��|#��Y`�k��^��e����۫��|���tӐ̫�u�r��q̨��I&��P��E)��=���gY���;Ztn����p= �]1_ ��)���U����)�Ϭ�D9����I(q޵��u�����]��$B�%�@�3ܠ.�Υ(R�c&��q�=���N�v�tǯ[���椟6�;/�\��Xk����4U-��G9_|�l+��`��m��+=xl ]��(�k�P�0䣘�^�{��!WKGCW����!K��yKz;�<8�pw���de�s:��ŵ72��k�ˠ�b�d�7�5��%�6��2�ՙJp�շX+fdh��c���
&��Z�ޕ�]�/R�+V��f"��o`-�E�+�r��5i��aZtS��
��w��2a�*�\S-��j@84��Z���*�Ν$�Rkh�܅�r�++U��wo)���t̕�#l+'R�����۲�F��5u�8f��9V�J=��O\\�(���5�P���O��H�܆3bŐY^�b�H+���H�|a6��M�$�J�L�0ƙk�b5�lĀ�@1+�$�m�cAB�Ш��Y�ĚB�����(`�@�Ib)'�]��AH�06����hCh��Z��
�<CdZ過3i6�bi 6�2�)�mY��f�6��7�(�	���°��T*c1���5J��q1@�6�m-����=ȱC-1�&:a�l�YLr�V6̻�e]"�����+Q�p�Ŷ�fZi��J�1�S2�B�)X�ۃ[n*�۔�&�a4�j��J�n��(��1%T_��ʋ(���<vɤ���g��WI���P��*�`,�.�2bi�\�ˎ5x����%B����2��&��Ĭ�VUaX�+QCi�I�*bQ�J�@+[u�J��Hc=��ꯩ�ټ[ů�ܘ���zy��N�W���338���*n@.�U��vWS*�ˤj���g6�����e�P�75�z����uJ��׷	�����?�>遍�Q9�# �fdI��slZ�!qӰ���X+k˽�Z��#�yu�W�{2?.���h��)aӵ+�,Jɠ���⡙���U)P���۷|��{o͉B�{ˌX���V�3��Η[ࡗ�La�~Z�ov�y��a	��)��d&�T�u�Y@�7%dD!Wu7ۘZ�1S��Dyp1m�|S-��&y��g�� *��u���Խ��^�ds53�f�ѻ��ᮐ������Іf�H�0
��W�T�]��S��\�hīx�.��|�յδ�4v���_��ű�l茙�P(M纮�r�'�ռrM3t�q���͎�k�����'���2�tP�#٦�����v4#�����J��w��3<xt�i����N�V�#-�<��O������_�;����Z�YRU�fK���53;��;듩�ƶ�td�J�]�t�yv6��ǳ6�e�mlݏ}g���\��wr~�UWt�N��Jձ� ս�6�Xz�f�W����o�f�=2)��K=��ڞ���}�KK��JySv:u���۴�x���u)vw�t^�S�z�Ú�d_+X����yXP�k[$ɫ�`��V6�m��x�dB8-�r*[���ˤ�R�ܜ�i7����)��r���Xk�q��m�+&�Uu����g(���?�h�4��I2GV��yQZ�3��aӎ_a
�)���^��U��Ӻ�����i)
�:�j�P�̦C���R�2��\�o�BӔ������A��mߩ��"���þ�}	tq��;�L흗�=ʦ�Dj����y b|��($��
:�b���;	ֹ��:�-���{"}X���"72X��3M���/H��!]}G�H0U@�e��zI���e>�D���m�jM\)239�:��*����:Hw�WG؝��-�U��"�o8�1f\Vűp��K��iwc{�n��6S�N1B��	�vwIUbj�#wp�++�{�*��  ���s�3;�>s���gh����'���2dr5�-���'jy�ָ]8�����'����m������\��ǵ�R]�E�ɜ{=5��O�@�p)��� y�no]��tV�気�v�K�{<��j�¾����-ݹ��č}6���&�*���u�,FT�l7%#ܡ
��|�9��lQL���W�7��;ܡ�V�5���!fuK�5�p
hH�H���ܩ��[�~z�g�ϖK�:�_5�����j\)�B5O����J뚞[�L�J���	���&�P���擊���+��X��q�!q�iڼJ�i�q���r�TS��f������!4o��JP�`�؜Q��%�|��E���V�dD��졚�{��S�q���@XtO�>�ebP)�=n���6*7+w_�
�{@*��w9"�	ҕ��ƶLuh�/-�YG(t@0��;�-;�
��7o+�`�Y�tҒw;I��Įwf+���{��#��*��˗��
0,ʶ���m��l�0�,v�,Vp�K6+�������V�h1�;�����w]�@V�Խ�䙐�>Xt�Z�kcY�Zq����s$
��y�!l�绩����*q#L�����:y��o�<6��0��5=ѐ�=C:E3��8ǀ�zİ�mL8�5{==��/E����*�׼X~Սt*�8<���ŻWuS�n&��gZ&S��2q"]v�o�r^D��MԷ<n:�z��J1Q��;,s�����F����@t�+�/ұL�Q�/#��m*c���pP���޶a&Ά�2ly�zi6�9[�XAOl�a���\�G0�&��v�ᖤk��h��[�|�nw��k�8���w��ߢO��� Nƛ���$^6(f��7Z�m���B���׭.^��y����ӭ�Y��;L��x�ɤ74/�:3\�f%�Ub	�#�:�S�����>�wr�3�bf��un9R�ޚ�T79���NݧC@MZ��w����t@a�خ���Ŧ߀�3&;���.�F�bS�N�E����3��3�\�C�㠺�����NR;�cm_�ﻺ�#Ǽ���-�T��� ���ۜ޻�ϓZ��ݛ�RG����ǒ���� ˗'}ـ�n+���5�S6E���%������Hf\^{VfS�69�k"紴���__���nyo+
7�c��Z��t>�7&�}rm'�Eܽ3I�yh����9�.g*�]��+�8�����!u�]���z�m���}<#�T}ލ���݄�R��Lł����)��.Q���ȇ/��}��ɡ�Emb�w�d��7[&�>λ�MR]V����)�}g�lZVM��-�Ǘo&�Xq���[ν�`�m�X����ą&Uf��Fؙ��΃�{7���ҵ����Q"�-qlSg �n%I�C��Qo�t$��Q�77���v��b�#�3���/�f�90oÞC�8�w��M�_Jc���>��p��s_Vò�~���a^�q�ii˩���w�z�A,{=�媕�o,�u�S�Y�jr� �%	4vܮ�N��.�@�4Yq���=�m�^XM\w����u���j�����K��x{�+:����*���O�% uKw�3���	6k����K���D�i>�-L/ [��oJɩn��(P�z�kF*xբ�S|����OW����=���1_�%Sޖ�R������`�s�`=t-�w��5%�6�z�N��J�����M�9�뾔�=)�x�W�Y��!�ߤ�l:<��.g����V��ʫ�Q�o�f����T��$]8���PH�~m�������T��<��ov] �u���%�Ջz��ʫ�����}��Aϫ�2/��~Ī��[˔<�X�k��Ȓ��&{p6��pL��X��)����x�W�T���8��f�;���<��f�z�Z��	��d�J.{!um����#�$M�tUމ��'+3��Pz�}��/��x(r��o$V���Sw+o�\l,��� �K�Yb�7������ے���*��<�5�+_��v+~m,�f���86�gRwrm�טn5�_`������'j\	Qw8�d�K�(܂��L۔�O9��[q5Xr���"9/���xm.���^.�Y��m�=
�:�MT
��S!�3R�2���[�ێ����H^�xv����ͨ{>0�{���O ht�|���t욲�}�z ���:MW�t���`S>���,b�ؠ��4��gQë����[��wݨ�8��0��P=�;�b�k�9���ć�2w:)N7�̩ƽ�z-B���0�!e���.e_���n�d��� ��*֧���?'��L��{X0՗Jm _^B��Kuֺ����^@�#���x{�=%Z���V٠�fM�&1lG3���Pז�]�ɀ�N3+s�1��v�2�uMִug��$��y��M�������h�g���iwt4�U�x���#��c���[��vl+�k��������6�+)n�6�lܹ�SM���w�r�x�uTKsrLwQC^�h���]�{+��FmT;^WG�V�t<*f(%���`ᥫ��{=nw~���Q�,�K��G��Nn4l�]��<����}��.��:�jc�&MF��n�#�5�c��<�v����o{]������ ��k��Ҙ������Ԕ�c���Hu&k�*Ҿi]�c)v�������+���v;֔W�9=�ºh��~;hO��������.��Se�-s�5�����4ϖu�����+���xۅ�nKno�o!j�QO��YY�|�uՀڨ�8�/5�Fy��3�K��}בk�a�V:�QY� ��S�]{b��k�+T�^��~����3{��C3p��y��[��6
�	Λ]�6�!l�܁����{ �*�0���h�ǉ����[0�3�3R�2࡝4�,<��(jB��tMn�4R�
��}�kΔJ�*�����Nܬ��R�j����Ɣ�������O:���j)��!7�X]�;E���y��ڷz�uu�������RT��3��:���@tк���5�B�-�y@�F�?c�R8�B��F�57.��2��=�/�w,j��ql\����N��TGj]��3kkk��7�'wkP�7/S��v��+�b�"2���|��hW،�Wq6�x5A��N�VŮ������^`�/P��(�����W>���s�3���#jxP�S�`���$�ֳ2l>&+��3N$Ft�����cA��~��.{;e
�Z�zщV���ng4Bs.L��/��)������U��~y�*�5O)���[ �ܴ���e��h������vm���3NN�L�Cf�Ʌ�ށ\|īΉ�^�Ԗ���k����f�w����}Z/��4�ϩ2^���2��-�\��O�)ȡ��$�1ͯ�smBt�tu�]h���F������=wY��ȫp���ZR��<��;o���S-T#�#��
�R�Kv6���=@�V�T*�����E<�m���4�eV��w��ilmj�0�Bva
�UFӯB�ۄ�h
Ӝ��a����[J�����L���,:e��7��hr�}_��w�qV.i�yU�Y���^4T<�^[��-\$Ȍq��Ԑ�$<�3�����P��o�z��U�va*<���A�tG{�L;� ]����|yx��w6Ji�fZ:��d)��q*� ��+�]b��J욝�?hx{���rLZw۷_��uX��	L�fZç}R�2����Mq�C2`,�ʫ�5+;1�b]fq��>�rO`9p����������M:�"��s}��7L����6/�P0ąŰٸ)�^
L��H��-*W�SL)���s�䞪O"k�'X"9m��f�9B`�9�y*���/�9c3�#�1���w�RR:��̞`���JM��Tb�9��[���k����Vc��������=R�v�OX�'��۰��]V�M�Gw���O��{�6&=�b$r9�r1��&�<0{]`�~-�/ό�n�+��:w�$���6�ɺ��dq�\���0�7��W_Z�aq�z��k�+]<�ݫ�ת�o\�=��x�Aݹ�����܍��Lt�# _$o]h�ܩ�:��ݛv��� �ll��g�3krz���B��p�4�H�哶�Z�<�ҕ8U��:6o�9dYz�lj�eu���yR�Rk��R��W���I_����貛DZ뫉�vwmɟp��Y oiΠ�:����u�K�����v�7A��Es�s[��m�4&��=��Fz��^m<y�ߗ�v��X�f�C�۠�f��� �NK�QI������z�֟+3���T�I%5����'a�����]�<Ն�Ś-<�PmU�m+}mGaFnU�޸�m��C��1�a��Xy{��b��W>t�ԯ{�rOAXog4�U�̩gh]\*��j�JJ�芫Hw+��j�c��v�K�B��8к�:�J'X�{���cN����
�8�[g5�P
T�Y��ۆU��ۑ]�䅉rT�*�qM����Pd�߹��s����ŢC]�o$/{M=�2�i�,%Z���Gl�����SkF�;�����Wp������:y��{H���6��c��"�!�yN�%�L����ky9\��Z�sϜKu^&;v�fښ�$�T�f�ނ�;���#g)(���F�Z1K�7����|�]���v����]H�N�����vfNx�����R��R	�',���
����խ3K���Ìv��q
��tӝ�Wl�n�֥��'Le\�vn��sg$1L�h�ܕ�����}��(�̙�Ϋ��;�kg Q��>����siI$�H!�l�w����ܳ d��)���F33/1�
Z7�5�*���W))��а��v�Z�9�[v�Zd���Z�Rv+��_t8�m��ٜ���G���B�K:&wub��}2��\6�q�P��ŀfBv�Nf�Ҹ4!� ���F���uK\��/'���z{�*��Q\�ҫCo+r��-�����s�Iv��3^[C@�e�V�1�낙�'m�r�"�v�$��5!Jg,s\Ū���������u,(T[s/�[��n��;T��o���iʫ�BTԠ��PRa����Q�PwR}ܭ}̕xլ
�4lu3x](.��'��FGh�4vg��@o"
R�1�]8���Y��Her��r�]�9����۱�+VQl�6i3��x*:]���]Acw#�l[D�+k�l�s�yJ#p����B�ڏ/l���S�s�򅳈Z
�]G1x�c�r���a̭�<SR͚�t�9=�އ"�����qp���!�Ѱ3uZ�m�����LN��s���os���(7ڕ꫉���C{SK��Fs�L]ˈ�4�th+�kGy�4k^��t!��\�P�G-��܇I��a٦;�d�*�n��>�gTw���V�4Mn�l�|��k*kww�-Z�9w%�|3��{ďY�a��X
6�R	�c�fRVC�7�����b`�L��V
��2�`��L��V ۍ*,X�T�*[d�bc�j�I+3�vX:)�i"�a�L�o �=Ab��PR�Y}IUd�J�YXM E1�YS�Kf��:@���&>[��&%Bi��P�P-H�E�}�4�el�B��+1���"��F)ID�IuC�.Y�d�����&	uLsT1�&����I7��M��.��Is0*c1�Y5LE�VL�AE���.�Xm��i0I��̪�=³�)�10�T��AI�,Z�lEQAC"�LsY�Er�(;i4X� P!4$&WdY�_4y�`�7]��17����V2Ѝ������g,�BvH[�.�������^�oZɵߠ=� ����K"(S����w��~ɲ\�}-���C�x��M�ŊWֹ;Hlu�,>>:��4Bɧ=B���`bYY�ʨ�r�b�C�bSS���u�i�Z�L�·�B��0���δ���U�w=�;�#ǓK���{P�fןY��m�
��)��<�r�f<��F5n�T�ec��Z���S���zS)��,:f�lb��fw!zbj	][����p�54�:�,���û��O o�8�&Q�C{��8������(�}�����S�GU`p1�,PH{Օ'�#^�����ml��Y9-����Ӷ���St�{G�7�����9# .뙼O��	Ng��-$Wܡ���,�Վ�/����H��Jy�v�4�x�(��ԙh�Nk��"e����K>�/�H���q�P�=Wд&�]\0g=��,�	�fK!\�C�����_��õ�JRGZ�ظ�&���ϽOΔFm�(�Yc�R�E��Q|��\[�ɵ�Z�ܗ�h����
Ն�c�!٬_[�#/)\�:R�������Og��4}��7��f1[f��fM�1lD���luaqQd�2�N�A*<�py�²ָ�^�gӽ���$����^d�j��M���[�0�L����_mʿ���}�X�7��o��v���+JWF��HҬ��9��-�Yʶc�!�M���F�3]�䧕<�c���
�V�����]�=\�R���h��Hu&r�#V���Q��E�(����w-0�sE�c���ს��ה�B��\��j���K"+���s�yZ�u�i�,<�C<8���+�8�Jͫ�A�ǭ¤Z���Vj�{��6�+��Y���.o/.Ve�ʹ�j����vW]{p���r�S�{0g�2ug8��뺨�������m3ꗸl��	Mi�X�hB��o�/U���弦 f|�k(����y�MjWq��;ѕ7��]�f��z"�ȓ(����,ciwX�]㧣��2�X��y�K�0f*K�:;N�ry�A�� ��ne\�r�k��x�Ū�YZ�q�e�`���z��"����.��xx��R����p>��D���Xt�=��r/P�*{E.Bn��\�Y��3BT�_[lJ��4�ą&Uy�j��W8�N��yͧm���*���r'�(OqlSG �n$B��t��͇q"�`X�5i=�<�F۩̼\6"�;�-������H��:zTT��lN�	�������3�n��v��~��JM���q�7�0Ay�$���n��&@�>�|�]e����B�Z��oZ1��<�^�q�q��������b}��'֎l����Bxج�#����C��榦�{��9���ɫv�wf�؟k���ճ~���υ4/�%Pי@Ƭؙ�ι�l��Z�Jj�koU��vm�HIFU���)X���V��y? ����o�����1�=}�m��:r�·8FC�)���G�T�Q�c]=c�o�@&��\Ax���b�E=k�(!�Ub=X&�Sr�g,UdvOU%�cꙙde�i��IҾ}ڳ���[�ҺN��c�6gvf㚴X�[K5������z0F�#�V���UO���;Rι���=� .�p�/��?r�G3"�Z�J�����Vn;�L�R�Dָݙ�q��8�z���7��E)�\WK���"�k�ڨ�&౻�6ES�z�;�����.<$t>�~+&�Q�x!u�N� V0�����;^r��k�W;)�>.��.>�e9��*���E�
�D�Z�T���9���wS���JfS2�a�>�]~���PiĒ5�x��]�;zMe�;d�}�Ԟ��NW��׮B^�eb<�fk�|�,�3g���U��o(bB�ئ�A���ɋ��䕭��B~7�E�R�[���Λ~�V����$>)���u�x�'�nF�^��fw��ch�;@��\��jz���dϹ���7J*�9����ʎ+�i.�g�f�y��p�
�䬚�ꦮ���������˥c�17,���y���d�ߺ-���b�b�_5���&���w4��L�L�;B����dsؠ��"��6]9���R]����ɔ��3f2�[[F��G��4��u�m$�fd�ٙƑ���^f�9j�L%�� {�M�x�-��	���9̓�d��}�I��Hxw���x�<>�X2�ɈLd����z��;�I=CL5�:�Y'�~�}�A>����u]��d��|�]�o��vq&2|��? |��ْM�w�rN5���9�I��Xs���?3I�;�?2��O��LI��rO��!������G��/�������r�|9IK�Y'�;�u���<���>jM��? q�G�֡8����<z�~O'{�u'�w�N�?!��Oy�=a5��P�<4�ˌ��A���,����Q��Rߤ��6�����M!���Y'�5�u���jyO�8��I��'Rm�������'P��2N��>`y���xq��(��&��]���uG�S�!�\b�$�/{�c'����u&�?"��>I�7ga>a��'֒zy~@�2x{d��6�<�q��(~!<�K�\_7W�5�����D
>��U�q
��
I4_��1��X�fC�>d��<�Hq�5�;�$��N2|��9�>a�u'��8��>�����i���/����k�=���3��t�a���Ւ~B�|���:��VO�`j}�N���֠�8�����XN2T�M?$����_�N��Iނ~����V�d}�$�Q�=�@�H|�����	�CS�a�Hi&v����1=��	ԕ5�0Y'SG=������P��<j�d8��/�=O�Qy��SZ��>��|{�~B|�����'�Hz����!�'�y�m���O7ܓ�6Ɉ�\ԓ�*js�
�	�k��VO��{W>�*��i�ie�K�wN/W�" G�O�;���57W�IԚ��=Bu7��=g�JβO�{s$�B}��!�N���d�I������(�_�Q}�i�矝�t�Ev_
��L^õܯ�ۚ�\�^�¥�4����"��ن�
�J�p~5!���g�G�]��j��vE���d,�x'�7 ��%Ӷ��nۏ*�Г�l��6��}A\��e��}��W���'�>�t�������gߟ9������'�c������O,����}B(u���:�=CE̓�=��{��|A>��Z�#�'�O�zk��xxɍN�����15>�B��|�fI��&�0��!�����'�P��8��B(I������G�,ᖯ�@��Z��׍r��?o��)'g;�'̝���%@�&55��'Y14sX��u��°������x�P���f���!Ć���d�:���}����w���^g��~����>d���,���s쓈����ԝd�7�a*�<t�ݲ����I:��fB��~Bn�$>C��@�P<Ͻ�"���
��3��}J��d����x��?"�紇�?2k��,'����v�&js�I�N�����I��� �+0=�~f!1&���AO���}]��̋�7)�*_b�	�6ó��'���L�E	��������{HxÌ����I<@��䜶�7{��O^�9����6�?��È��ޮ�xO�ڷ�Ѵ��>�����|É{���4�S�q0�3~Y��E	�,�';l�=�~@�M}��$���m�	�9퓌6������s>�:b����*������@��#��aR��>Ld<d���'�6���|�	�M0ѺqI��7gY:�!�)�'9l�=�~@�Ϲ��`zk�3ڐ�?V��N�]�='H������2'X�gYP��O�|�8�5y�2qP<�u�|��?"�e	�OXh�8�	�MMӌ��A�>d�'��	�;!%�gf�K�臨����>Gß��9C�>Bq��'P��0<�ܜa8�&�w�u�?}���"���u'�OQO��|����]$�$�����r���Y��X5���
�/!�Ȓ��F�G����2�C6t���m8�{ujj����}�G��i)N�P$$`��_.��l骥e���S���;�*t�è��4�c?N}����F��lJ_�����U=�gZ�9~>���{��&�̞2|��&��B|��>��|��́��6{�Y'�*h�
��'[�
��R[����3���Έ;���u��u{�{�HH�]2O�l�|�oXM��!��d��Y!�>���C\����:�m����0�&'��	�J����(�N��ݸ����$mV\��}ӫ����������O�<�Ť>@�n�O�St��o�l�d��?2Vd:�����XNs�8��:��y7�!��I�YE)�r^�4�qJvRcޢ=��*,'��=�VO��o(q��'�C�[�P��S�'6����	���<g�>�I����a/����f�9��_��:K��}� �{�_H$�Ɉ���$�f��
�$�7�r���7�:��&>��!�辡>@��:�g�N&�������(�+�ϊ��:����� �{@��$����w��:��&Znwy	�MsX�$�o��*O̆��H|�O���C�1�x����t���zwN~W.)v���(�A}���x�'�͏q�Ğ{������ԝd�,���	Y=d�Ms�	�Mg2zԓ�7�`T�>��}����q�W6z����m�=���}�~잲�=;N�>Hh��hi��3�"�d��क&��E��_}�q����w�J��&5����J�}�I������u��s�[�^������}
��q�췬��<g�y������C��id�,6��N�{�pY%a���u�&:9̓�����4�#�h����oׂ��;�I~�ǻ��BVN�����&$��`T=g�Cao�'���Ԝd���M2u�>g䘓���=�<I�O�̒m�;�f�龣����"f��;ڪ�퐁]��p��6if��C��%�Rf5f�A�]@����v�2F�v���&W�ui��m6զăi��Xv��{*J���-̾���ަ�|��^H��|m;\�X�I>���F����[�o\*������~��C�3��=d1?~�3��^s��?2k	�C��γ�'�o�i���5垤�'QCs��'�A-F?��fmo;�ۇ�{����
$����쓉<z��w�C���L�,YO��p����~�$��~CN$���{7gI?!��'Bw�o��F.�:2���5�>D'�ȁ�<>�d�9�a8���d<N�����uY�;�'Y�~f��w�!�G9�C�l�'�m��,���!{�����8�}��=޻������J�$���:�ְ��^�q��ɹ�'I���I�ܤ���~�ل���{gXN0�����G�1��<d�{����k{����������kϺM$�&�eBq'�;7O�d�a���>k	��>d�O2y�'a��Нd?}���	�<��'��H���#�G��|�7���߾w���+8�i/(VO�`v~�'|��)Y2x��t�VI�
ΰ��Iy`|�OY<d���'�П2�i�Z��9�0n�1�Koe�
!�&'N��d�B���QI:��
������̞�!�O{�|��M�g�N���d��<�x|@��W���E����KFw�ݷ�ćN�'�>Hi&v����1��a'RT���E�u����Y�N�|��:�����q�F����3�v�x�ީ�ʮ���׋��P�=d�Xq�����u	����d�a��0��LE��0��*k��]Y'Y�l*O�d?�>I��y��@u�]
��������o�jL���V|���������&�P�I��l�gP�}T���Y>�0��Ɉ��'Y19�,�����+<@�O���B��_xΌ�&rzP��f"��75����Y��ov�n~!�9��2��"<�U��n\�(p��+m�xOE����e�j-�Q���8��6��
b�o�W6���r�D3��]e݉�"��P�a�d�{�ry~xxxzh� �����|�8@�=`z�kxz����8�g�P�{d1����$�nd�E$�����E�}��zɖ���&3�O���8����9�.�4|<��| �Y>d6_������MY:�z�ky=BqG�C���l��2a�0Y%I�l�E$�ְ�'Z��s�kY�o.�~י��^�����d�N�ܐX�>�'�$�!���T�2���x�Xy�'OS[��$5>��d�g�bO�E�T������������B߯n��3v���G��)ǽ�y� ��d��$��o�d�HT�s'�BbM}܅C�~d7oR��=a�8�x���2u�H|��1��������sy^l�s�?����$���}��xɮ}�r�&:y�u��R�X�ۤ�}��*g���b>�
������)'�h�W�����#��2;�r��R���	t��E�����:��,=@���'﹭I<d���'�~N{d����������p��C_����&$�ϧ�DG����>4�,�����Y�i���I>Cw��,��jn�2uC�=a�N�'�h�8��3!8����'�RO���:�o��H~C�4��<0�z��;X�5���m����G���d�vk!8�Hh�8�$�����N�	�)�q�<`~d�M�r�|�����Bu��:����N�0��UQ"r�Z�ro�G�"��|�8�j�2q��y�d:�l��g�P�$�����0Ѻq��I<~@��d�퓌$۰�I�;��LkX~�/o�]|�2�����8�����>B����ԓ�~ϐ�O�`n}�����,��C���ݝՒ|�fS��5�ל�0�:���l��g�M���M(DM�m���*��%�<��e��dԸ�o[�ݱ��_Z�"�G�4˝��י��K�W��Ҳe��8�M��9�ju|�#�Qc�N�ӝK�<.�1Q�[d��5�*��u":�b�Q[����]0��  .�)��7/����4��9�:�k|�����3�f��7=�,����
,��;aY>E��ل��=jKHq�4nϵa8��(�V�5dܟ�~�쯾;��-_	#�h�{�?d�m�'��u!�=f���8�h�q�RI�]���&&���*j�E�u59�d�l����|�i�|5�N��_�cVb���Nw���>W�';�>a��N����<g�M�ać�<M��Hu	��0��u�I���q&�1�椝ISS��TO��>����)�]nlc�8�π��8�x}�`x��}a�0=a���IԚ7g�T�	�߶P���7�u�~A�N��'��|��:�'���u'�L ��֕��"㉻��~s>�� 	#���VI�>�
����:���I�j���1�z���,����v{B(u�'�u�z��̓������f��,����"���G����}�� L?2cS}��'2���>�
�o�M����4�Cɪ����'�P��8͞Њ��k�}���ó:b�C����_���G�u#�AI?rԜd�?C��TRcS���d��P���>>̅a��������P8��h7�Y$�~~�\�r���s}?k���|$��}��@d���IR{�'Qa3��';l�m&3����S���RN����x��?^d��x�P�^s������s?<L��_xxa�������2|��6������a?s$�L��jN�u���C��=M'��rx� �F��=|`ι}�kV��7��¡�8�v��'�z�g�d����L�I5��Ru����!�d�?w4�x���rNZ�y��O�<�w<8�#�h� }o�j���]����JV�ٝ��\��sL���K��6���K��x�M��4G^�\�Ԝ�M��]/Y�1��PS�r�J8Ut��<�)�[k8�\�*�)T�����AU�U�P8�˨�1��q��=�m�mr����;�fP�&}���C.ʴ�]Jus�=+���&��+����@�]�40���k:�3��:�s�]){��J츾yq䃊ڃc�s����J��@�P�W��(�CP垃
�Q��p�4�+�3��Z5�@|��E��/J���wB�T��z@�sPɳ4�N��n�v�>��O{xY�bR�<���zb���J�,�x���G��uuR�4+�����^ass\�)_NiBF��Z�f��M�Z�s�H]t��Ϝ�3d���^ɕ|�wSr72؜���	9�$EQ����-,����3,�����4Mnuc����K��]b�\W[���W��P9%d+���a��g�Z�vmn���o�$�KaA���tX�k�?E+���-�V�;���9��N���mwP�a�t�� ����\w"m�ξ5��v��b�7W+q5בl�\4�R��ap��%��!�7������F>��=%�x���7B�]^�O�oU�h�M���sE��MN�VTu��n��/o+f5�I�8�h��d�#��!�<9
H
���0�\�
M�**�%)I>�~ܬ^���w}-�C�]h�}|+`���ݜےI$�I5uv���LU��.���\�V�{���kl<�]KV����C]NL��]mGI]��M�P-5�V�0R@:�wa88��5[w}Q��t*�Bk)�R��;X&�h��Z��[Ƹ�BE�L�cG�u�{t�� :k�Gz�ȓ�3f��@�y2l�0C��B�eMG`Vg�.�-O��[ŶoY��=u��.��[*h�;�SH�)YB���tP�" �K�ݮ�t�c8b3_.�96� ��JXۤrS�˝7^^�l9R��&�}i�9Oy��}	j��Y��h��\���M	ĺ\<H�G�6i�	��\�+-^Y4�]	�W'c)۬g/���{J�<�,y����R��gt-)�-"��˿z�#���5�/dB�2���%h�S���]����� ��l>�W���@��r���dB�aV�&�Z���ʴ�gs�̘�P�Vt��:�6��n�w�+0����<��RK�k�N�z�]a'�\-*u�k���'/94�fc+��7&S��g��+�����]�L��K�гy��l�*J��YȬ��A�N�Ü,�8�����Yyt��R��t,��'q��Vw&��!�kwke6#�˘��jJcRF��$�J�W��)�V.�U�*�|�&+�d*E�E����aX����b�Ż�J��c��5l(�]ZE�-��-����P�P�E��Lf%A�&Z�
�XV.�PƪʅJ2 (x�(,Ģ(֠�DC�oUKj���&��g�B�'ΘO�X���6��"��DE�����Lk�� i�d�/�kv�Y����*���:£T��<��1�A<�
²x�Rj�q.ys�T�3v��w.��U��ۻ5�XZSW�3-*���@m*|��{�����PR*#�,(���e���Q2��*8U��̦AX�MZ��<˅�S[�L��뉈{w��0���>�   �DaL8�jP�&4�%;�5û���jR�cX�+CF�JT�8�I�7x��\�Y{[iNĖǔ�"mN�-�U��<��W��c#��<2`�3���gY��Ma������LH)�C���:ͤ>�y�CI�RT���Θu�E�~�d��Ì+���@�'��y��Owx��|�}��y�ǭ���Y�^Z���� q��;����P���:s���Lf�|��m�g�ɤ>a�?3n{�!�J��f�
~f��:�a�YP7�>Փ��w)1��@��"Ś���/�≯}%�E_o�-������y�A��
O�1��z}��N��S�YԘ��=q6�w�&�'9̚t�QO=��>ev�����b$��l�E�A@�s,��1 ��ه����5۷��%�V|8��h�q��>�G��G�f���@�}�4������k$�m=g�1g{���C����7�P�J�џ}��L��B����fز~�A��}�Di��F�P�,:�R�!Ȭ�R00�S���L�
7��g����p���0w���3z�5
�+�7z�Qῠl��ܩ돳d,�����(�r�&�1@������}�58CkW�K�h8�X2��ºQ�tӈQ���E�X]!Z�E!�ZY5e���//g�܈~}<aq�ȍu>e�}hfѨ.�_	���L(8��u�gFN^5�Ӯݵe��(�ӤDR��Lć�O1�ӀT#�a�4.��W�]��'�=�=��TA.�y����ᢝy����\�8`������>!֕B�گy��g̸���;�F;syu�FE���t�3s4�>���M{n��b��jS�|�T�J���`�WfÂL�U��'(6��fn�@�Y�I�j\u8���(�3��B�������e��r��hr��V��rY�Io�{���gc9[����bo�
H\]0m�:f*YdH�$�]&k!Z�/1ʹ�5+��لr]֑7R�v2I��(A���yC�j"��`%=�	��Đ����{��M���(ף�M�TΚ�(�W4^E���3��ISfh���&�m�y]$WL��%�Rp�3`�o��uMŎ领Ŗw�Y
d<��0�w���޻�%z��i�yh�.r�����3��t+H��P��\c�<ɼK�b��겗3.}g��|bV���B�N�$H����3��mZ���3�r\Wdh�ƹ��C�R<��í�F����]���1F�̘���ۦ���Ӓx�F_JF0�\�qާH��Ft6�G:�D�a����O����}��lmD�2��E��eg�\Ōr'ܷ�$a�
��=�,$�7I�2�R'�Ý��D��K�����Hք�h~��t3R��y��7=�qp�3_�qM��E7��Sh�wx�?��щV����6��.h�[^|��C��1ֆ3��lغ�8:ȇ����X���ɫ2�m!q�*�Q�"5����R�n���u#���P�ko�6�}T������s�z{$������'LP����B()�9J�ʸ���0`����$�G/]����62;O(��f��3��C!i�^T�(��{"����)�GY�v��BNw�����1[V<�^��W���p�g̴挍�L�g��Xgb(]*ٍ�҅���;�#5��W�tB!�G(;�[�����\����ҩ��~	�͖x~�>�Q\!���k���a�V������F����%�Hg	�$X\e��v��'�zH��K�,]��z+(�;s,��he�*��L��I,F��Q����O�c��+1� �ar��Bkץ���������u�����%��"��u^����r�Ak�ѪQq3�~j�Ć��ҀsdP�=�!@�({� c\��q9#���XF��Cp���:��J~������Ǟ�AU�-<1�J#j��k�N��S�q�搁Gp�κ�z�DiX��ŁNX���Zϐ0��:�	���X��(i��f���E�j�;:��3�7��=,��¶Zm�졾��3>q�o&���B�!܆uF1���JΎR�kzԽ�ڕ����j�d��[Ⱥ�μ���v�b���9X��>6���,̤� x
[�R�n�f��e��x�D����_�ҧ�ױҡ��+s~z��"f�ij5q6ﵦXɾ�!#]��u�7��@���_\\8���0pFy]3�l7��,�)�ά����ΟǸ�Ӟi���J���(_/�_�f˃|^9���֨�c����K��`��.{s���>d�L���gU4<�e3-�77)Z�7d��:�<�xq+8��׫��-����R�]g0]xC#�3���(�h��YF08��X[�;OX'�d?K�js���Y���̚nz�n,��Y�yi��0V��؜�;�ނ}AA��A�q�H�ق����
�۸�[�0(%A��'}��Nfs�B�h���E]:�X��
�zgJ�l���r�k��؇
j�5؏x�O=ܻ˥�<�ctF�J�W 4���U�X?����|�SXt�s=�ϓSkW��ɠ�3�b��3J�Юs�Hg�'iO��Q�E{�&���iO1�!YY�_Tz�}A�S�+kQF�,��I�̛�p��K߲7�̉��3��E#i:I��3M؇�����=�ѧ�S�Ep����ӷA���a��@�mmdI���'ق\�n�tRٮ�xn��'Yb�r&����=)}���]��9�����vԞ�@�H�>�ќ3��5�[r]����b�Gn^��׳U����mM��_U�xS�7��ETnǉh@��|��E�PhϢ}�����'�����wnۡ����Z�3����T��T�k�i��.�� j��y��^0A� ��J��;��}����9���<v�Ҏ���{`"w&��,�-
�ۓ�&�
��)Vdk^Gx�V������a�}�KA�ZJ���|��p�B�ͻ�Si��W�9���:�p��2"��8b���a��z�j0
�2)	@[�gJ.#;�v���^Ho�OZ��o"��qb㽅�t�î7b�����#3�6c�W�VU�V]�I��[�I�dת��H��,‎��x�}.���,ˊ,�wU��� +�:��܈yܫ��n�#Q��������AF�#je��$lP�p�����ya$�;�Vb��P/�\�*Ƀ�FK��t�K>�Uj���݊-¨���2vo�3Try�K!c��T���m��ö�k,�ļ���w,]u�;��!�����8�Woݣ<7�3�XkM�8�d��9��v�Nv������	ٕ��e9S�be�����+��K$�O�&����+{T�*�]��K�I��� ��פ7��r��0�\>p����r�w)J/"�HQ+cne���T�U�"�N������Xgb(:�ѱ!Κ pT�`�^I�lN$Ԙ���v��kQL(x6p{rg�3��g���![Wk�g��u����*�W�j[�7��w@�4R�L�����B�g�eW6Y��l�1y�2�
F�0�b^,�n���9��C��v�
 �`�\]0l6gL�K,��$�Ee����{s�ru�a�P�[��(���u,�c$��B�ءG�8�jc"b��3=��Nh]�'ҷ��K�p�hYՁļ �����qA[��
����y�Ǜj�ծVNr�E��r�oBк0�Q�.�*�/x����p��N�U�i�Nf��o�,%=:��O��l��/������3���	��u̠T��S���u=��sY��co������k����<r�G!y�p'�PJ��oE&���^��%ň�1Rt�e�xM�u����ֹ�3!ׯM�Uk��qN\/�Fܐ��U��/��t��b�w)�4;9&����F�yسvp�X�wb��-p�JM��F�!7�9܌n�]b�
��mՍ�+8O%��� �O=a:)F��-�3��+���ʩ�8F�m�6�֝����A7Rt�^U��gB�YKl�2ȟWI:h�`H���X�땄hr�l��ۑ��y�I{�ʛ�������|�١�0r������Q��B*��9�z�˻	�2S�]�N��u@m	"��t+��x�ѣ&Q�B�R6&�<m�"�3���Ҝ��S���ǒ�Eő��1��=��g���J&���7�ו��Db��IZ]�2p�F�q��LԹ�FTB��$�YQ�N��ȁ�3��6�/pM�K��O�]_��v�a�G.H��@�Qv�Y�`R�b�3�ea�JKz�z^����OǔrY�VZ>�<D�W��d��^�#k�e��,(���M���V\����DqT�p,�o����@�<X����(R�-�1�֘�w;:ޅSҬ�1���%��	���	�¶�dkÞ �;ڛp'�J��V��y��,�%Й1<i 뽋g��޳�e��:ݠz�"���6yj͓��q�i4���luV�6[ˇI&�os��e��y�E��0я��R�))H0ԅ��i��u<�0�-� �դ��q���R���fOϾ���s����`�T�N`옠��Q�񈜝�>��\�Cb���}6���f#$k�]�<x��&�%>�J�q��֪KxȾ4&*:�Eʧ��F��M���Ʃ�D�B0p2/b��'8q�y^f��V�}pbF��2i3��..w-U�t��;�ky#,9r�i�p�C!�7Wu�|L�X*v�Я�� �>Y�?t7M��[�2[}L�F��GO�I��Lő�O)�W�ڱ��![���&�ji���o�T�::��������4��:�u}JW��qţ�k�=�ޓ۲�1�9��/9Z�<w`_��:=����Lm]%S���^%�/�.��7=ܸ�[�����bC=�yD`��tzyp.���TdjQ����s�p�:���X47�Q2�R�*bݞ8F(G�e�9ބp��'LW�Q,�8��.�d�X���Ft�W����re�4+�JEʞ�85ϲ�m#K%�4��Ĕ1����� �ث⑆��v������>Z��r���J�����,\[V��W�u1z��'*lX�Vg'OQ�bJ�=�/�����$>�22d9������[F��cJ��p7s7�s�2>�t�Dk��[�)�p��%��m�u��tTN�+�u�r	;1gO����Q�r�yXW�����gNP'�4/���ճ�����]���4`=�`��3�K�-E�6=-\����-�/��4#��3�^���g��3���̴*o�n��Z!�r�HuB&j���JO�*�r��`�S�8{H�<d�Q��U���?<��/��3��IW��o�Z�O�a:O#z����U��|S��E�&�q��=>3���;V��B&3�ن$e�SFp�Rv�ҭ�-�,*>�����y��3^�<�H�����2.*�z0�09�#0d�E����~���V�/��A��/GJ.�F��*Q�D�l���R��	;q�p�U���unon�W]����5�G��"�f��u��k�B&��eV���4`z;��";0�����n�v[sǲ�<�n���j4��deF7<nay�24�2��d��,^���hzN�U&�o�YI]����6�2���$Ȥ$m[��A:�������ya�&��q��l:�ޗ�e�Z��?+��8žp�=��U[�﯌@����>�1���cN���X����1�-٨���R��f%������Ȅ.+k���8��_b-=�΢7N,ᝲ�9Ĺ?~���]ұ��;d�F�{���CTۍ���3�:�v*�P���#,9kD_��lw^w>�d{ݯ9*����C	��ن1K8�#��<Q���:r̿EOt����-�w|�;��M��K��Ml�V&_2������l�Q��R�.z�a�@�U&+F�߷+����OD��W8*���F���/��Y�+�ܲ�U;�k�
F���K�{{;Y��P&F/Hu��p4a��`�������(�=�6jt{"0&-������m�qb�i�iK1^��}����z'��tk�z�v�A�6�rs6���-��L�?J�4#e� HX����Q���{����Ԧ֘�F��u����k[ӶQ�Ɨ��K#Cqz��`ߔ3�W�K3J�*�l��=c�s�ܯt��gZ�m��yc�b2��f-���'ˋ��gM���W���b"���ܵy���0=^A8l�晿5�֊ʶ�+�X�J�
g�ءG�8������p��w]���9���jpAO��Ok�R��-�Q�t���<����|��ԤD���m�\�,uD������ǖze�
K��m�.��;��X!�͕���7�7�AWZ�8�s�t&h,�RdC�Xc�s�K���n��/f��C/{/�%��Wv����p`�s��GYv�ܺ��8��'�@�[���C����qW �z�;
!{*[]ݢ	���a�R�����"}&�!��nv�f�r�r>2T��5X�J�͙A*�������ׅU��\�ʖrR��P�y�M���y+�M�L�X���p=ǹ��\�������\�+[�(N�>�S��*U�zoVS5&�U���ݻ�荮�GVӣ���]��6I�.�0�)�r�{$��B��Gq̱mn3-��,�e����z닄�!9���I�sE��S0+m�3uR���9
Tx��c���p��:�2����1�H�q[J�D���s�Yy[��+)�Nq�:��Kdw���,��Ǽp��������zH��MY�����@�O7r7,,��
ێ��}��ƕQVP
	��!T�;�a;���5-t�lj�P��`��k�.�]R3�������%<h�ڝ�J[�o1��-�r�Y�IpS'xǴ����dȚ��Cљ#A�Xf+'lb �W]xu�����"�vM\�Y�!b�LWw���(�I$�@*]Yzm��f���(�:�RqL��J��rN��+����\��VD��)��� ���uӕ�^o�\2qμ���@\�l'3R���̊�VJҪvSP���u����ٮ��\UM�\�]>qYd�L�=�̥�7:wVRo2��ݑ��CS�M*Bf�ȝ��"��o��ճMjLLDμ��L͸5K��W[;GaF Mw%���-˧�L���wp�}H�*�jź��V�ݬK����ɐ�B.}S��:t���ofe@�k�&Z���v�]$�:PSA䣠�Ֆ�Rʕ0����ŒwRب���ŵ/�}LK�n f�+o��r#v�3����y�ױ5���ڝ�w��a-b�� ݝ��B��.L���IvJ�[}�i�Rc����6�[}�M�P�
�Lb]Ηٰ�����5I�n�:�OW�r�����'3E<RM���L��/e�U�Dt��|��A�Ή9�ɪ]�:��*���	�E�j�;���*_E�����Vĝ�
BNV�ʡ���GcYs5�v6��L�Yҹ\��ns١,�Qܼ�uٔ�T<b�'�,�܈u;��9+���at�_K�:�d����!�r�(��H�L�yҌ֜�n[�r�ܘ+����݃�I��o� ��ym��J��jI%�!�j�]2bu�d�+1+���iiKZ����TAfҊ�Ve���vmQ�,Y����B�Lh(���wj�1&��.R�K�{|�#��a*W�P�����0�2��AMU�.3"1Ty}ʬAUT�h%�c�m�QLB��AJ������ц`J.d��M5�f:t��[�@�Ze�(#���"�iɻ
0R"�3�+F��1[��"����U��c��n���˫A��*"�+3,ո�+QTHŊ*��iv-�U�hͲ����X�<�b*��Q�W���
����UY�7�b�*��J�EG��ԬQ��-����QF-�DQV�=��,bDTSM�Z��7J#5�	����$�����V���}[B����Urá���E�֢�l���FvC�oWj�YKQɘ�w��n�m��]�xxm�v����\L~�]�A�5� �3�E�7�C�����L{�� ����O�s~�ù��*ܵ��J�ڈ+z��
�l�SS�F��W��	N��}&u�hf��\C���~�g˥DJ�y�ӷ���Ǳbhr�����Dg��5��7P���zL}{���8yG����͜����:G!y�y��PJ���I鱗�&/EZ�����]��X�R*y�1K���Q\���F��o]i��,�#un�B��s>Ry��#.�8X�U����	�j�]�
�*sjs}���NMM=;^�NV%��dvf�a�"8���N��ɔv�}�E)� �w
�QW�7R�/*��x �Y�rĦ�4&�V�� tBc�z�
P���K��~o��P+�����w�����[~��Y�Ñl��س��@�Ȭbt�/Hz�B()�9~�\u��&�1뷆�wU#�b��|x��(�Ҋ�,֊u���RL���^^]n8_euC��<"/o�2وo��Ok���y���Q�3ņc竨���Bz56�=����'<Tۧ�J����%��㴑)�wnn�%�j�j剑�W-8�W� ]�+���U�Y�Z�6�vJΗ
K��P���&��@�
B��R���!@��Y�:a�m�Vd]*f*�3��X<"�C�X�5XuD7Y[1�R�б,��9AX�{���e��T��^čC�����潝��&�M�(�ႰY�М���b/��poЁ�QW�"X�]��7��V�E)�*�0�1��\�~�AX��0a<,)����-xu��d蚎�c
�q<�h]M�fVA~Q��xq" s����	�h%b�|y}y
"%�!�oN:��+j��=��]1��i�\���s�JYq��MTo,�Ƅ�W���i�i/� ���fWz����QC�u�	A�����԰9�ħ�x?��x1�2ޖ�ϦO+�*��mc���{�X�ug�y(��Ҋ���u��	A��B�%�_�i�u��5�'U���{�Z;ς�KC�� ����#J�r��v�kW�3]үo�SV;r_�u�wxE��s�X*�ѷԴ[��=\8����:zw��Ŗ�鄃)��VQ����R��v���QxqmX&॒GX3�%b�*���^�m�s�|�	0r�*ޅb�؎m%y�Lǹ�.-g$�E,���XL+}},����Y��A�,�8V��yy��ڵ�	|<�ɽ��wl��n��Y�@�j�J%dk����GdU�<hZ�,�j�k����6�-Y��/��w�+c�FG�q�r;mm�ڗ��T��t��|�˝s;��8%�l�Wz��]�\�3�41��1Q.�28�;�i2�N�Q�ܞr���:1�U	��N�-~S<��Y,ɯ7=q7amK*����6�sy�<5��2_�3��g�@�n�qF���;Y*a�!��V�����
I'{f���&v*�t
{����Uo��f��y^�2�BmR�"ɤ# l�t��z9W�z,�����_K="�؂���v"f�q�,	S���ƜFB[T�RY+�cs�v"t���^2�w�J��1~w,�yQ��s�Hg�'EK�԰Q>	l�|a���^��F=B��"��Os�5�,#,��Fp�Rv��Yc�8X}��e]F���-k�ʓw2X�g&�q�3	ǉ��H��L<Qd���X�F-#�ଡx�Vz�}�.G� C�SqD�I:�ݝc{yY�4KUƎC��^�4ޖ�u��`_O�!d��2\yE�.���;-G�^gZjmƙ��.�c9���Q<��;e̴�u�wJl�u�x��n��-���߀{����fon�q�9*�.�mH�,�hu�!ᑅІ�5K�I;qw&v�ԥ��ʹ�WU�<X�$��A�x)�x�Z�`h�M�\�Lu�k�D��4�I'7����x`r��/��ʜ�z@��Rk֧LT�ʊ�7\.����|+~��{�2�R�ݖ;���ٛ-�R<t�����7�s�(C�XyK:�2��ԫ~��6�fq�sq�k��h,r�D^��yJ45M��n�C5�9��c��HU�@��Z�=&׊vawb��o]�~LP��Q�J��R�XR�r�(�9���n���,�y�_�����ȹ(����o�94�D.04d;Sy��vȥЍ��Y��D��3�'�JE�]Y�=dA�lWQ0K�Z��^w���k>�\�鎸��M+���R[W\(�s���bA;��fv��T�^�0_��[9��;8k���z7����nD�Z�E]:�r!(f8>"�����S�}\a�.�p(L)��JC�*U.��v�v$v��4�������泆;��k��w�8�w������ ��ȵB��A�����va�R�M�X�!�.\0Yq�s�����T1��ˮ0�Q�h�Q�eۀ�dӃf:�&����{o��V�oEI��M�P�:kǗ��!c��	s�=�Uv�Y�գS�T��3ռ<���������d�2L�q�D�yC:ER���8dEnԙݦ�=�s�^iFz���eHȬ��c2�b,[t(�`���f0�9Bj���(l�s}lmw!Òp8�xn���5�N��Vׅz� �܅8ؐS�k/L�u����Z�)��WyQ����ׅ֠�Y��Wh�r�+�.�p�.3՘,:ޤ�J�6.����S'��n�睐nN&�#6(C�f�Hʺ��0�i��Ŏf/{9H��+�5ao��c��e7\{"�x��X�SN������$��ni��ǜ���9�z�:8ҏy+p���g�WH�/;��(��J�5�\������E/U%��Ь�)1K��dj��T��s�i��#`=u�i�:`�<��=U���M��m������&x���4
f��H��y]ps���u�(�R,/�F�M�����%���x�2R)�Æ�̃���W���9m4с�[�]#W["��l^��Yɷ��v��c٭9�:�
8�}(ɫw'A��V�X���U���i���_u^;6�nΕ�-M�kmLj��5.�Z��p���J�PUH�Td.i���+>K���_@��pA�<�����M]���g.M�f�����S�{X��.�G�z!�`�2��r�Z��p\��uK�L���ݰ�/ #��f���6,��1X�A�0�o�qȊ�W�"�\��Z1�c���bzl�玛��,�Ɣdj���\lͩ��	xTi�v�S�k���ބ�e����
�|�:��|�'���iH�r������24R�b��͆_�^*9n���sG�JO���<1т�Ӧ�u���
��fQ7e�͡]9=<J�=�]��q����Q��
�Z6��f7�Quz�y�u�,U�B�N��AZ��k�b��9쫧r���A/����o�� �S��4�}xѬ�ef9,a]ԵC\�{n	�����4��/x�"��TWܰ���^����><TU�}�pO��L;}[�����7skM�Д��5�9�VU$7��Pl�<�{ ���q�˓������wz9�ל�@��ӿZ�X�+�oA!�q�t�ܧ}yxjf��:�w��j���l�S�G�fca��Tml�]���y\��]�vn�
��&{F�v�gpt� ��ۼ�7�5�&m��39�Rr�s�益p=�rx�Nl��B$��0P6iƍbp׹K��+�כ�Õ�����c���u�֜��2Xl�#b#NV�G*搁@p���`����^�K�^�(�S�ERnZ�Ů�w�e�2hj�5�W��w��C �.�.�`�[��xbY�^{�q�Js{.1`9
��z��6+��S��X�K:�wԠ_�ʮ.*f2�����p�\�[S�\�T3��WLߵ��8�3�õB�(������#�(Zǻ/:we�(C�+kVR7�\��[�o��F�J%�q�9�1A����G���7G��;�tVMTzb�nV�d�
��W��8E�oa�3P,�g��VG�����엽7��=�!Xs���<s}jhP�U�.T������,�d�Q5�nU����u;��98�H0�TAf����3�"�e���tLu�ؘE���2:#U]�,�m<UΒ�YpŹ��PqYXcb2�W��pȠ��3�l<����L@��N��ܩ���c�"��f�x��\�/M�������X�H1�%�u<�ve<�5�+�S\��@�<�憏f�<��9�z�˙�nK~{c:��t8�H��]�u�S����Ӕ<���-.?m�j�`�"�H�f����]0�����MC��o`q�:F���b%C;#�؂��<�����\h��8h<N��*�cw�{���9�Ot�LS$�25N���i��JY�1��u���x��Qcw2 #�3�*����6Yxȸ3�n��ږ ��}^h���S�%��=�	1�����l�-���5\#7g�0Q�Dc��(���=Y�1�4�u۽�]� >�p�.�pY��w)��MxW���4�_�0��5K���V(����rL�ߗ�����x���B
�"߅��>Pm�\4:���Up�u���4������X]1MK�~��a�*�?OaH_%R����C���뫋�K{�j�X�\��8�IUa�k�G�F�ϟ��1'�X�i�.yk9fY@T���N��
��T*��ॅ�P��0k��,oO�r�kTۍn^�,�اr0$�Hʲ�q�Ra�U��q��B�P�&��"\(�Z���,��HFyO_ڽsL��~n�������L1�[K}]3��a�]����8���_N�lҗݜ�x�؜n�|ڣM�gƴݜ�j�*����-<˫lW:����Z�g�K��|�po*QZ&D���3��oe��v��)�U��{�Skm�����,�9N��JhtB�FC�8QU�c�E	�3��^b|.�m�=�|b�g�����<|Pȼ�8X�Lz�K���jh�� ��<�4럹��Z=�Gb������$k�	��hq�"��}"�Q���{���,�Pm��j�ڱvF�ƿL���B�,��8jDpJY�|E�6!�=��.0˂�!���1-�����(Q蠗F��-r�ꏗ�=aK"	�T�&bB׵`oD2���z�.��9(����xvӶi���>Y ̷5����(gH�R���9������<a�8���L\qc%R���HȟVXG�����x�\\�E����s��Z�]�|�4R䈁��t{�i��V�SG½1 �ө�x����iMC��Ǘ-����}���6g�2��׃��-�-����s(y����2��ڱ�k�1<��+�7`q�Bh��U3��HK���.ƞz�)���v};%p�7q�J�6����X-�Zz��E�D{��%gM�YR��B�JA
Wvz�(}#R�3ga\߷X!�K&ݭ�iԬ�;i?�o]mvͫ�GJ�<��vZ�Z���T��	����ٮ���䟟}B���Me����䦊�����vyu{����y��0�V*G��q��ԝ�kxtC	�
�̰j�:)�Ofp�j:����rOcW�M�
ޗ+p/)n�!���s8j� F�JBb�Y���T��s�im�=���x�#��דgi��4��:p��"E)'M�	ґ���r��c����8��bNsU�e�Ù����W
fB术?;��k���	�����#Ad�3�;�lvĳ��T��ް�(��,k:"�L�g��т!=n��]N�)\�J�v�]�����͔k���ߔ,��'Lb�w��.�(0��,�!?u-ݿ9�7��S(�Sdt��,�Ҍ�T�]:���^�]���`hA�'�vd�;Q����=�p��N��?�m�xc5zZ�5�9�:��]�Vd)a�z�m`�������)��}bX8KQb9�k��xT�����*��C�kY'������R�/��"n\�Li��1����Tf0[����y��i^�c�����Ҙ92'���Iut.��5Q �cG�g"ܺo엔^]�Ɗy���<�qB[J�|%C��)]�ʰ�Տ��iˬ�}�����V�pwb_$�������R�"��ժ��G<��t	���1C�W��2�T=wd�l��a��R��Ӷ�+y��]�t�IA:�s\�ջv�n�8�igfrZ�\C��(�.�:��4��o|XV���
����iܩC�G��#q7����p���@X�+�;��J�R�۝΁�.��V�� �6�����v��CP�ƒf��*�բ�Ҭ�6�̘�q&��Fk
�+D�MԚx����S9�Y(ȏ!Q,��ƚ�\�}utL��=�XF	��S&�}��d.ӚR�ְ�
�����>*,�.��&p��i�n�����h@��E�|g���{vIYb"y�U#���Պ�oJ��usIl���I\���1�K���]_
z��.�ӻxLXk���2����W�#��d�3E��1�w����ͬ'�ʋyJ!�;{մ�5K8c ��R��ڒ����ܻY���脊y��b���� �"��Ѭ"v+5��¹v��ʵ˶&�A��m,��ct9ܕ������k`ѻ�vȅn��oU�}���[si�Av]m��8H�p�n��5^�U�
��rI$�I Cg�g�AT�η����U�rq�W��=k��2�W��i�y���ȋ�N�X��e=͆���O��榪 6�[V�Ⱦ�y�s�f��Բ%۪c�B`��m^��6W�c^��|�2��o+al\n��d��b���n�{[;��Y=�9I�'od�͈�̂�35W:����o2�'լ`U�_9��n�M��լ�Ty!f�'�p����C(.���ϓ�S֯%dmY�Nԙ	p�j;ax��:w�q�nЖ��B��%#���[o%]�M:����ie�m�9ث*):���k���:p)4* ��+:�3o���v�6�ԕ�WWv5�\����������\�Z��VF�ɨ���dU���죓hb�v��A]-̭/�`3�������m�FT:k
���jl��'vWB��i4�y=���E��fWp������q�X�MP'ܩѷ�2��,�� K�
XՒ�=�ɬ���)���čs�2�g�]�����NI�Z�.
Mc�`V��(ghT��W{Yzc�Iphϻ@�o����;�|Cܵu�}z����t��-���Y���-��k�ϵc鋐�0�S;��5̛�Y;�}�AD�l�R*�kP�7��\�IiI$���|�0Tԧ�e�c�Ɋ�m�Q�҂�X�GL�g��+0f�n���Tg��Z�����բ��5%CYf ��Q��V"0"���[�֪�2�A�"Ȣm�%�v��V0QX��LEQ@U"��ۦUJ�Q"��IEƊ#�`�T�*DT?%E�b�#D���*�"
�E��Q �"(�h����U���#[QS-DA4��l�wh�J*��EUH�"� ��E������cP*��1��J����eOi�1D������*�EDQv�q*J�����DWID��"��H�0AEUY*U�UM�
�
���1�2��Db�X{��,TPQ �<��(���X�����J�Ъ��!���t�H��.9|���n�}������_HWs�^eή����s�ר�}�����f8TBŌ�t�+
Lmϓe���S���[=����"��U����.H��(xV�ל3��j.�@��@���J��1�M�}�Jە6[μ�����B��)���LE:󈐨��=A1��tBx0����ϣ���Ί^�7�HH�> /@��߹��9Bkץ��/�-M�W����hʝXC�SƲ.�{6�ѯs}�}�\E���E[Uʃ�+ULE7�/��j�������u�FÅ�%�F�8k���y>g[�Õ��KEeg+����ɎR<�ޞ�#
�d��[!��.i�P�Fu��t�8�n:��+;YؑU7פ0�֙�7Zd=�-�ς��7��Y��]�~��k� v��y&�/{RZWޯOWN�Pd��׶l+�"�fpз=q����Ceo��|�"��������.�Z�jNCH��(�ʥ�\�S��gpׯ��"��k�����nk�N�:X�D�mJ��GmJ7�Q�8u��{LSˁ~_x##R���9��Eݭ+�5���z<d��[G)������=��j2�N��k��1���u����*Z���\N�
OM>�k�^�3���c���fp�����U�v�?op�o�Ĝ������;z���L�I��C��/i���s���߫ﳛ�����%EX�6+j��u���"�"�e♂P,�gz���;~�%<^��w�X�x�8T z�s��]\N�>qS\��L��\��u�x zzv��o�{������ʬ�q��:�,�L�\xh��>t�p{k�)x�<=<9�y�M���u=	���v�!,�ۆ-��8�pAea��˥^ˀ��^�B����6�p�.�l�Y�<U�5��lFR�zE��S5A�'b4M:�DB�*z]7QY�e,vo-;��at�Gl�a�f�|d2h%L옰�3^Tf�8��ʰwff1�-�i�;7/ԧ�Y(�#�3pf'��46����}��1I�3nbb�b�rނ�����gLHN���3V3��n�*��g�=T(�NU��_�X�`�,������;y��>�o�}[�5�]KU,�W�֯��`���
��X����m�O��[w�_�V��f�rL�,�~�������ܿ�@=S�j�ܒ��tA��FQ�r]mnS��za�֡�V�5�[s+\��I=u{V�7n�cz0K�``��)q`�,
.��Os���q^��SZ�Z�H�{����GvpІpn�꛻Ϟ�*7f��t�#�����_%2&����t�_�{ىY�a����<9M#�5��zyM�Ѳ����i��h�F�P3l�ݻ��3���,���ǔ͝w(�*��{Cvf�Θ�}c��ڎ�-ܓ6ə�����y��0hgJ."���9J5�m�盧��q�o([�r�����u��RF0�i�bL���O\�OC�]At���d:W���ǻ��q�v͹Նfs!��|Ђ��Z�jT��Bz[����B*��!��d-�ר%�MNB/�W��R�3���)%U�tO	�}kF�Zϖ�'+�E7ںar�{�׃��(�nU��	�^��ɚ�k�qȰ�|�\Vn,uK��Vw��CGӳ��e��~]!Z�Eh�ZnD_��b��VU��h�Y�<L����~Z_!m����V��B,R�.�#{i�!�#�$��*dA5*��L�d�{�Hv�sΞ�N�׽j���u�hC�pF������E�"��=���y]-�X��]گ~L�f����WFό��
�x�1�ݷ%p޽��E���i̰f���#�϶�Ŋ�}�f����D�w��f�ΝmQw����Z����G�H�nN*
������v7�g&�_I���g[3��3�����X��n�W�Ϊ*1t��.��`�+,#X̄hd�ۯ�=0���7Wv���S�f�ft�P�8WG��PW��È����
h�W�&!e�5�����
T�,� �.�T�w���E��a�Z���22�}p=ڎ�~�<��ǢV�򷷷'X��'�zI� jf��J�1ev��D�vA�����U�N����lvf^��-��F��Ω���4P�l�a���a6�g���h-9�Wy��k��9X�m6)oB�%�:bF�W2���2�������
u��.7���y�����kޫ3&ǁ�s����̡J��(�}��NqP�w~��'e�=4���对5}�[n��c��I���!��� 41����
�81��+�Θ���A9�-ڂ<y&�t"��DTwEv�:ug�	�v�ϸ��l�����mx��w6�����w�,b�#����<���$tE&]
�q��z���O��v���S�y،��48�zHDK
���Z�-�C�9od|km⿥Z}G0|��P�O�V��)�ڝ��M�N7H�N�V3�\��N\�1�Z���m��'�f��O]s��ZT3�vO�-V�&�_g^뻸dBRv�N	+8O%���U�S֌���i�`#>�(ڀ���(ս�6�qdV1:b�������+�d�i9S�f�����2Ͼ�o���XyA��(�V���<h��HdQ�n]��Ԛ�B�&XTq���a��>����xK4�4���Ej>�K�����i�k_S����������ņv"�t�f7J;b��.�{���ɬ�-��+7m��g\��m� l^Ċ陮l���xV�ל2�ᨻ����4�>>�wh����&ցޥu��7
�[a��@:�F��&l���ٔ�0�F�:�s*c�-��؀A}�D(| _{B��܈������k�j�9S����<��e��dOGP��;�B`�9�JTǉu�
Cn��A���Y���nM�=RggAn�"�OdT����PP5�n5����."^O�}�Nn�Nrt��;[���=����,uO�i(vR��U�!��Њ�FF��s���-�p��vU�؛��fԹ�FT��
��˗�*�Y�����\Ȣ�lz� v�K�Ǿ9��'7~�Q'n�ߤ�f���Z/�˷�ؓ�AICx-�N��r�3d��-��ɜ���mȵfno���5|=�2�{y�������![^K��{����U�d�hb>/\"M�&b!)ࠎ�{X�B}��Mz�Z���)�lڻ�(&gz����Y�`͕lI<T�[|��2(d�ܳѓ��<P�t�뗪p����_i�(e,�n,��kp{�~{I��0���8��>F��F��!di�^��9F(9�6�}�Ȭ�ؓ�W��뵑��0�Y|#&0�:�Ч�4R�
ڮ�j�1��0Pg�-w\��^��E�m��Ȟ��02ރ�L+]�?��r��?\����v���Iz�/Os���:�*%�,ČTAf��W���]�[����w��׊
^�S�P�;��J�grN�H��v�)Ę�^pAea���t��b8f��m*܎�u7�e���wu�[�T�`d��X�J�́��lFR�zE��32+s��
۞�@��Du���e��b��;p�	E�\�1ߟ�J��1aܳ4���h�~�*��[9Gend��q2�ݎ���t�'"6
��N!���iSnܭ5��=�@�L�����T�	��4u�b^>d0g4��>�"�'5|&MD�l���c{�L�Q�Jn��;"UmNc)I��;�pV�̘��l';�����x�D�����MxE��_��
�ྫ!��������}A�8f&���&nS�Ռm��/y�B_Y��<�jC��U�Yl�ў"r"}��2c��=9���o��w�i.��I��8���Xƙs��5,�k�P5�e�Vn^�H)��t�J���؁5�[��8Ç�rLF��������hvׂ����.MjK{+_J�Ŀt���CF�r���cX=������ZJ���+����J6vn[H7%#��L X��VF�k�Vw(�F�p�=��3|�L�,��r��k�ٙ݇�vw�����'���	t��t�;�yIs��H�"%�ʼ���4�9��/`q�h�)R����B}��2��\'8Y�%�o��d�v�C�s��J���,���j�� +C��u����>O�xs;*wغ;��j���j3�S,�O�a� A�Z�;>4�}��삺>��֩Z�1�q�P��CY` �c��wxi���Sf_�*WW*}��s�OO`�u���2 a�4i�@�}Qe5k&���զD�U��;��;2Ɨq���*���9����(¢��w��ߞ�����G8�'�η��$�.�SQ�t��Ͱ�z��e�UlH&��	��Aq���|����G'��eM�ո5P�xn��Ñ/Ck�O��dUӭ7"-)f)�$,3�Y<%q�е�-��U��gMxX��laz 3{�LÖGlI{J�M	T�t���3$M��gf��-q�ۨFx]OFM��r�a�5�r��C#/�e���M���+C�*vV�5/'��kBq��\�p��ˑ��aT��x�P�W�޺�3˫FM���os�u��P#��@��阩e�� �}&k �=���]i.����CV���)���$�� ��(Q�"�jc!�� ��5�5�����\ ܓ��Ւ��[�ʺ��c
��o'�>�`ζhM �6`"*�_D���^,��^�d:�0_b��tqV5u�[��nD�V�S|����O�����/���p���G�{;�e�ᔽ^��4��X���N����P�����x.�d샼v��my`{n�ڐ�6���c�%_��m�׭�h��Vs��#YV����hȲ*�:�.lr�[r�Q�9����"��1���#�ScÊg7z��31�3��p�*�`p��t��چ�cټC�x���a��*��{��z�{��▅���Zd��(R��F�����ʧ3 �a[�8�{oyb�9���F��l=u�k��A7Rt���Gb8��$��f@t\�XS��~Z嵒�������L�S#:r!�����\���T{Nh��J"']T�:��H�D2ʸ��K*��Ȟ[�(��/�Ď��ˠx�Pʉz�~�7��]�ݗ�Eٱ ��'U��3jx�����Gm�q��qdP�'LP���E��9v�r��-�����>��S,蟦ȨS�M��Y��jY�s���s���ȕ�q����%�ʍ0:\�1�(t��;nYʁ{�X�,ֈz-dl�<��n���*��2%K0Y�(,3�t�f7J;V%�5�(+�K�	+��u*�Zk!O<�܁��39�-uS�/bC�fT�L#ő�ϖ���F�-�g�&���?9}���L�w��8L1"��-��7:b��`Tj���6E [�;#mF��ڲ$����M�o�Vzl$VN���z޷#�N����{g:t��{�Z(�;c9�s)�Y(ө��s}�k/N�S�t��v�ծXm����vDh�C�J�K��������J�r;|��8N���b�K�
�ϓje�+�&yN�����9�#!�e��Xi��*+�&��e�j�[��8&?wP���~vk`������0�R!}�$%L��h�dV(�J��W��4��������T43Ue�ϗ*�Ex�P���R�x��%4��~[),�B>�S����m���9�X���cF4��f�\�(�hF^95w5;����Ia��J��؅E����!c��;�N���D��mB�At�ޙ����k'28�)�P�j�␭���j��������WB�G��oς��Xn}6�2���gܮ���^��8��t��{"ڞ�2�S<OjN�J�n�q��2E��vܸ���թF�s�k�lqV�^�����;�~땳���p�����xIG���}/ÅoK�>�pe?Zf�\Un�>�ofb�z%���28�>.��WD��E�S��\z���>|�v]��K�� �㧧�4L�Ai�눭��S��w��nEZ3�]�r���ȹ�YR��A����I�8�!���ݾ7R��r��j)mH	�a�6BڌEv������[� ��
F.1�Ʈn��t1bTttH�H�6F�
�)�r+���{R�-*�8]u�U��r���eѬ�vS�{�k=���!;{��ۚ�Y�Է>:��etλ�X�veE��m.���XW��*D5�S5�{�596�S\�oDO^=;��Z ��Kz��u;����Y3wKwʕq��|�N%$��\�Vm�b�����W�Qd�P����Μ)��;ƧSl�5���6�!�4:m��m����� �����nܙkv��X�-;ю��Rf@�6��S˰����W��Z6���8Z<_t�e>��V�a �G�	!Ϻ��l�A⺎�SG���:K���Ɲ���|b[�Om�R�G��ܣ��N�c�f�ܠ��N�%�$��R�%h�����5�,��J��@�us"8)��;te�3kZʻ׻u,��9��kӁT�<��ǹd��ܭ���=2kc�$���v_�"�h賓#��Yoy�Z5ʶh9�D�I�W6o������X�<c�Pj�bd���]�\���h�	W�i��s����9����m�h�@�v�^�/�ZYᑥdV���:���XT<�xa׾e�ْt3yv����A�ȗc�e�Ԥ�I$�J̳�[��ϲ1Ԫ�2�������$�le<���h���}���{� �b�tJ�����}�Dq�r�Ѭ���2����񁲗��O%���wN�I,ѻA�ƞgnմ��;�Y��ԙs���n��
Ы$-N
��C�%�)T�U�����|N�BuEZ&k�{�(
�6>�n�yLlV_%�mP���*ʼ8��r�u�Qqe���Ay��r�K��[K�OV����`�S�l޹��m����/IT\��R�6��&�v��j�mجW����7V���N�s�[μ�Fmn.C��6dW]�L)�I!ա�4��7nE��\�����:�ɏ�m�C�Ňg2J/Es�i�V9|:�Mϭ(oD�Z�Y�V0���澧MA�Nw5*Yk�49���-o,��j�z��C�3���3��h\�_�Q�5܁� �z�P�5c��RQ(����=�����]�)E�nW<[���>��i�����E����WH�HC�'Q0���g;S֑u&*����� R�ծw[�Eʛ��dtv�m���Fuf�K3�f*Ϣ��h�#$&.�(ݲ)�u�ֻ�~K�ous�����Ŝ��Epr�:�ə��L�p�* B8�Ens�oJكbmwF$���I�s*��Ċ�������b��H��QV(�kT`��R((ꕑb�J�R����B�őq��j�`V)m�,m10��M!�`���Դ�*D@�2�(���U"�MY<d\Q�ƥ��LE�B,<J�+��(cj�T�UW� �n$���U��Q��(
Ͱp����	�a���!�[q�T����1��*Eq�X�%Lb�un�Eq��UUE�PY�PEE���E�V]6**ChT.�c,]��1Z�A�)D�Q������qӃ
0�D`���.f"�!Q`�"���W��#��;�E�eb#R�V�I_�BV�/���RyL��H�eGʂ�:��حJ�S;�Sm�<���{��ɫ�a&}��>W(��JV�����>�����1��v�Y�y��'�uD�18���-3�p��Q�����4A]r�q���gN�M�F��[u�J��~f?+0)*!�8�;r��B6z�5|��G�X�\�탲XH�*�V�_�F��!���"T3�P����ԓ��V��jk���Cރ��C:<8!t�2��Y�s��e�|d2h%L옷r̈�MY���Xqq���RH�ӓ��>��G�>�3�n��ږ$e��	����=kއ�D%�}��綇>(��ϖ�RτWN낪f���|(�9	�TG�]�q�Z����-��w���� �s�|.!����;��c>����Q%�˩���'�{�A#�s�B�QRt��f��$��b3y��G���!�Y6�f_�G;�H-t�'"�f����F�v�i۩E�}/3�3e�o���`/׷}�H�d��������`�l�0�GyUa��)(L>�YI]�?ZB���!}<е�MRƼ�l����:��������n�R��!3ͭ��hD�[u����'���$p�Oo����,Ժ݊��v���2.XC��X�47fZ�/2oB�1*�J�'U�/5q���H����MNGNQY�Ÿ�ޱrd�1�og^��@=+3y��-�~�r�6�D��$m[�t"�8oO�B85M����3���4���Z�Ry�L<���"�5Z/(����t��x���|K��#�\0�<C*"r�o>S���
*6mC7L+�ǀ�!E�ZѨ1?'R�.�Ӈϗw�h,��|7-f�q�,�/����Ѝ�2�bF�s�P͉�x�x��e�ECD�qա'��<c�; u��ս�͆�\M�b�21zC��p ��qw��n��,��tӊ�0|�r�4�u���/"�H�+Tȩs��=����S�{�ة��ܒ�|K�u9��
t���¶7�R�MC�GtIz)S"	J,ks1r���jy[��N��J�jV�uu��١��d20D7�R��'!o9�e-��2��`�O�pO�l���قb��b"�+,#C��d��=�]�D���9�yY�'j*�7��阡,�%L�bV>�f��S����5�=�/f�
�e*FeQ�};�y�ál���L�[˚��{�WM9�T	��{R��n��.��:g,�S�3
T��:��)�n έ����΄�V�kL"c��y4���Y�Oʯ�Ꮪ��X�z�d��ä���(A�LP�����e]���k����<�8�^-��iS�p�mJ5�d���7����c�D]��}0bR�re�]��\��� WxϚ��hS��eօn]�R6%E|<2�����o*vycuǲ*���yWW��Z�-�&�Tl	4Ɍ�#̠h\c��zQN�G3P&�=�fr�j������&^�7���/�Z�)_�������P�y~�k+����*��M\�V��Jw�W�����|��^�Ô���S'��cZ)}|��t;����Hc�/���)ljk��ޞ0����r�l�
dgCnDw�R �D�F�ӫ<0	�wfȾX���GR�8>��.PL1WJ*����Aw�K����&]
�z��R�g��fI{�c;^�a�^R708ڎ4�HEdW�e��ځőX��塎^Elgf��ckW�JS#	���Q=�On�:^LU����#:8*����Ƕ�y�f��o��΢A>{(�W�:�SN�wVX�0��c�+2��gk��9�'�b�ڔ��0m����f�����By��T0�a_+�%��t�H�o�=�.�u�\�&c�{�Tup>������u�带5w�  S{����ٺ6g��i;L���eF�:Z`�r:B�\�g@���#�o3��3d(Kj�v���Qbګ2.�3!�3!a�NV��eY����Zu>7�E���g,���*����2��E�Hn߂u͖x]
�ϔ
��О�'�RN�/b�A!� /uׇ�~����7:b)לD�5L��3d9��[f���c������:,�,'jVZ���&L�0g����f7�L����s�QC������ufI���J�i��Dtq�S	=�4k܄��s�BRˈ�C[��+{�:��(�p�{�}S�ɯ(6Es��[�0P6iƍbp���'7km$��e�DKN��w6n�=d��.��/C�pL5��5}F�A�#K�3*.��X����dg;��߂�Ql-u�_��i�	֙4���X�#1g6Y���􌉻���aq�K:_�F����j�炐�͇���`+�4��`��3M�k4����v��v�a��I��6�\��ƭ��^�.����傀\�DIt�ͱ�a��A��,3˺�I��V�r�ck=�zV�{��Ӿ=X̩P�

�k��a��	]y6H�Rvs9���N�HJY��GHJ�}\zp�K6����)�n�ݖd��ģV��}(�����Q�WL��/T���v�hso��V�<ހ�DM�2͎�U]�㲋e����22?db8oȱ�#����9ݼ��|��^I���ƺ�c�Q��La�]�2�;���K�+U���Jkl�^�Ħ��!B0�[PYdq'=���(���hP�D(�s��L�����PfnZ]/62/��(��Y�M�\M�@���,��>��9��,Oz�a�%��Ҽ�C8�z��dxMUO)��U;�q&�8�pAfB�;B�W��_t�q��7M(�B�89F�hΗcelu̍%�f�����R�HuB
fd<�[�ƥ��x���TC_V�"�N
4�2���4"e��%K��� �l9c�<mrlz�ŋ~tf�-���C=9:9�VJ>eby��CjX3x�ml���H�]���^(Jp�>i��1A+Fk�Vܗj&*8ߡ�f�
�rnB9늨n3��2����w3[��S�m�p��-��Ip�wu�K��{&c��nJX�5����Ō� v�+Y���7c�6+���e�:^Q<_\�t��h�[ְܫ��9�,�42f�Q�t�o���Z����n�wLB)g$��f�-Md�΄��Ԇ�]0����kM��Y�4G�J�<QqџD�]��f�I��b���R2@�d3k5��J���m�Έc�P�@�. M$��[�8p��$��b�fsb�9�n�)8���a�<���Q��Md�U�ha�x�9��S��{_D���V\���������2�s����W�<:89���ZGxF�p�=��36�J�;ﳘhd_(��Ơ����3�(+�U�˨d��Ħ~p�)K�^_��]�ͯT��0��-F�U��!%RF[�ƴE�c�P�(H��
�T�/���k
vB�Cu������6�Ό�L͈���<s�.��p8�sC�L�0
��v�t����%��ǺWc�ބx)�q�;���<���b![weBYS&�
魼A���ī�a¨]�Vm�j��f�r�'�M�@i3\�������{�`g�A���iD��-x�³��Cn�����ߘks�=�\sV�aG��]9�3�^�^,B�5�!�3/�B������q�z\0o��W@#�h�m�ޏQ��%�s{�OX��2I,2�
�;�߄��]3	��YEQ�Ӝ�h��=ss��v1twm��]�����}�m�PQ��{���ס�p�hvk�z�u��-r��>^!C؊�T0{ט���-��z�
 yk�]H���`4���ć�a�4.�F�C!���1f5t�3Y��i�ݭW���E�a�:C�fp*����Yѱz�����\u�꧂��9�Ѹ�y�ҷ�d�^d�`�D�L�`GW��*����(��i��C��4R�˞��o��r"�)��K����bF�CQ��Ay��3��u�&&��\�R��t�1TΚ�(�W4]����7��ISf/�w3O�=���M�I�s{
���H�C�v߼o�W����*�.%>��> ��iK�F��Zo�#�԰�aO�-�|�6�d���W2��.1����uXHT��n�����XÌ'H�>��K�-�@E+�pR��6z�k>�5������3s��s%8��G�y�A�#��#o]i������Nh���W���3�qP^7��+.�HF�(+��:7�5t��1HĹ�i�F��+C���yÙ�x�����{�i��>�����wdrq�q���FU�,j�&93{\�?a��ڇ��Q��dl��������u�X�n�{V7Ow-�K� �7��c����-1��u��49[�qL��mȇ3�/GtWl`~v%ZO��̻WN�����������l(�x��`d��1��[AX藐,BC�L�.��7��U��/,0�ne�ʕIh�t���П-��\:��X���ő��!�w�94���hdv
�5�)�#|�x�E�,��v\�]/ô��]��+�g����˪�t�M��t�D�BIt��L.V�Q]m�_�c��i���}�E,^�7�zj�͓Sg#Z�ת;A�v}�'����g����6�DfU���R�Rsc�U�^y��B.��ntb��^��E�Ha�34����ӵ.��h�m�z_n9�5ۆf7�!|gM�U�F΁�
�HE%8b)W�D��E8�{�|zy���'%�1^��,h��he�+`�8�3��2�)�����1W�(Fo�&�� �6�43;�C�&��������^)yp����ؠC�"߯�^n��l�Qk/�ܩd����]h���*fͅr��!���`ᬪ.��t���nm�i�Yu]�(�d���pj�VsnWM2	�pqV8^&�z�WT=;�׽5\�t�����C�jvV-$;Eғ6R�ٻѼ��F����6��=p�sȏ�3�i�o*y@9���%H���Pu�|Q�/�D�6�$~��l]��zK�S�x?{y�d��C*��\�:r��g.%�b,;��y�j�]}(�Q�,_��V�\%Q{��b�؅���-�\KC���ק���__5��JJ]�(���������X�X�S���׶l+�"�fp�1Y����Vg=x=;��SK��!紴?�=\8����YE�t��\�R�g2�j	��ꙍGNW�k�C����V��>.���x������p��|+���k%���R*goS�6w/�0����>d�L��xn�!��O,'�r�����A��(gJ�K7Gkyݕ6X��ބA�g�����G�� E�0'����QV�r:�]��#�V�dT�Kޟfl��%�-�TN�@�1Q���>��9��o��*d�T�gn��v�`Pd����1׳�{���qN$��%A�W�
�D�y㭦<CҪ����N�`��a�㦠 ��uu8�s��zbipx�O4%6cܛA��f�lIC+s��e��n�k�cK���L6��-��-t������x������|�"g�#4�
q�R=��Z�V�lp{L�l'9v9��Vv�N{�To�"͟��j�Η{/c�L�3C5��lFxR�zE��5�*�9����:�~� !*��*�,���p��Y�z&Y��C&�Ֆe[�o�ۮ���Qo@�����9�^j��S��F�ebG7RE)�c�S�mr����L�>Lř�	�3^U�%��0])�������V[>�[�\۰�J/i5�8�3��n�&�q��']��f�N����R06G@�ݿsW�9,y)�E!�m⣵ǎ�p"=�\@�'n"Ì8p��$��IO����̥��<hz�{%�tp��)Ӧ����6V��d4`*�juF���^Ƿ"z���n������%�,�U���p]c]A�
a���o� }E	�͏{�ZTx�|���ݭI{�r�]��<�,�8�
��*�~}B��(��z} r�k��B��ʻ\�N�]��g)�X:�v*�P���#-��Z��ꯩ���i�\M�Ti�U��o��C{�͔Z�����]���կV�Q���+X�Y�/cFe6��M���b�ʮ��E�}،\����֎;�Ż���j2��]�$���{V{]jQ�O,����Ba8Q�:��I���<�s2�N�����-���l��6���P�|���_�)����˭�o��� �zA����E(�p������s��j��ŏ���[u��ۖ%��Zi����� �MfI+�����͆�,�zDL=XbvkM��Ճ�����k��]Kb�������a��kz��+��A�|) +j��oT��6�F��{��fs�r5Y�Ĺ9�bN�WR�$�нRe;�:�!ղ��CC�X15[�x&�1ۄ��`�%���Z�(�`��̝��
g�Ź{�t�P�`m�l5�N����W�����c��黍�!ek��h����>���\�<����k�^MH�kqkø�����i��Ю�.V(��Β�EBM��b�;R����I��/)�YS@���*�t�;��O�����U�5�;JJ��!	�ԷKݵB�%��N;�N�w�K:0}M���:�`�ⶑESI^r��.I���W�grF0_=�أD��@(�ƴe�W�a�!V�d��}𫘣��N7��疸���vT&��r�Q[n�	2�i�;���2���gu1��VE]
�	@E��-�r�A�z6��`��3�8�	:�G$�I$��30�/6�-���֣�j�\W�K�R���vC�e5�1��;���c(k�m8��-���I��i���L�	$�����MkMj"��ȳ�jZ�u �%���I�K:��M]��5�r���f� �y�u!��O>ëw;1�������`����-<�&��`�[i�pٍ��P�7 �ڜ�=�%C�j��]��I�Nb�ӫ�O��O��+9[����8�9�>Aܛ�	"=��䛮Z��%+���������:1�8Ï�O]$:�C�V:�k�Dý�z�+\�WwWU˙����j��M��IV�qm�e;W���G�T1���
r��A��tA�0��$��jƥPK�
n�#B���рk��V �k���I��?�L�K���-��GY1v�VΥy��)�jp���k���omfiQ�7w�F�I�2�[��uZ۫�*4�&�aL�tO71g7�f�X�bۭ:��]K��d��<�ft����.�]���Ht�F4���6�P6"��L�}Y��s���H�1.�;*Ver���Z�!H.��:�V�0	\o�uC��0�"�>x���d�#16s��Z�̤��A�옪�n�0A>��q7|nj����[щ,�X����`xi�$��	>��QAV)�(E�AbɲՕ�R\�b#1�dr����dQ@�X�0`��b��@R��>C�EX��1b�OPTQ��c�������(�c����Xk�U� b"
Da�����qdXm�_-b���Y�%E$�b�EP��"����X�P���GM?2֘¡�3(jЋ""�A`��
"�f!Y6�X��J�E��]����T��_V[Ad�yj���X�(Kl��P<O����(�I���;�9�몇'n+{\��B�T�a�G�R܂��^���/K�m��;x��5���-�}�ϑ{}S_,锿 ��Ju�s�UXk�H�!)�+�W��଱���!� T�Uj�5���!�2Rl�k��w���o{�zQ�28s�P�x������)t�b�vȤ]{"�k��v��Q� u�Pⅽ�ͷ*�o�L��R�Y�^��&V�� �F�F�}J~4t��BT�F�(��]"U�dU��i���6�1�gg]�oq�;)*0�f����/̢G��j�|&���L(�9g�:37m�n��G%N�a�f�����
Sѓu����r���d�RE�����;�^A[���ap�,Pΐ��
�*�uo%�Fe5XU<��X�i��r�6oE1V^A���`�D����f4K,�S$x8�xl��i��M�$6�1߷�sΌ3-�"@��#�d�<Ĉ66(W�(q�Ș��!�s�E�Múk��v�=�P�'�~��\Տ?��O9&�f��Tًw3#��9l�׭�++Fg�:�o��.}T^3a7�z�rڣo3���u\��)��],.�]<��}#�������e͝ʗ�%����{L�#���Kau�&�������JV��}$�J����U�v�}q*mU���ޭ�oe��gL=����1��pc��4���:E��c�o�7R&:��`�pՅ[�Ĭ[���(m>yȪ�����q��>01�X��g!
��yU��2��=C4��Ԙ�\z��9��?jKO �!�}�w�}���8�"����N�z�j���h�h�1?�7��$S��|��*L�o��[r�z�N�,�4��:p�&x�5w92�/UWj
XH�Q~-��#2��#\��8�Ft6�GO�3!sK��ӌ�w�O����+���,�\��9� �w!Qn�ag�K�5�nj��NV�L������t��ѓ,�n�#�Z�6�B+"�e���`���\��JKU��jƊ�E�����(�X�@�V���
��a�ڻ[�j��^ǲWH�Z46���Ӯ6fԆD�bK��`Pt�h U�S������{[�j������u�Y�l��tè�挅�T�P���a6��xOa�*�Y��PK�)��J��-���bW�G>���1ΫJ����n�]=Ϳ)�����]֢6�0d��Kd�5Y���6��tq�u'X������|v5zݪT�T�;�9��ݸ�w ��%g	�b��{՜��<;b �Ӳ6�rއ#h̷���6
/bEt�צa��
C��5�ܝc�םO@��B�PD}O��v���劼 iS�ޢ�借/�L�������w'}��z�2`΁\�
�:6�K�ux�c>+������0g��±`��YG'��W�b��>��,&��������p����v}闂��oR!�°���gs���^��니���EXj�ķ�sdl9�
�In8�@�o����es��섔?$'5."h<�3M�`���2�����p��Ux`J�K��UeS;��BK�x�U�o�o�
�Łwy�A�h:���iyk3���&���Sw|�t����I�^Jf,4��)�c�CN[�^ٰ��,Z�ww�.��K�wKN�J:�)��hж'�[�H��Td�w(r�f���9a���Ȼ�j�c��2�ךch��_Q���7�8`{�	eģd��$����Tn�<b�j�O7�usz��'�Ff����
��Wr��_]q�ވ^ΆQd��V��ޚ���5�k�j�K���tr�F�ï�g
�hM�RP��d�&7I���P���P�ܮ�7]Z4��Mm�si��k�������m��WSW�q=��r�S��Q��F�^Q�G~n��	�>e2��2"�ëu-sS�����a�L��>�(Qa��Lt�����k�X��'����N�k�T�T����z��^ͤid�&�s�p�f'Y��Ϥ8g�DT��=��־��+9 ��z���:�4xzj�
�|ߙ�nh�JC��Y�� �me�	-Eu4�L�ì�e�G�AK5zgJ����24�9׻�����1��R��+��<�l�-�T2������\d����4+�0���x��R���&�t22ҝ�R�Y-:�bùFh*2�x��
�Պ>_T��
���Gj��%�WUpnRμ�R[��k��}@>.���kC��`�>S5c>���V��n�^s3v��B�ⲑ�Th��T�����H�DĵY����6!J��Y���6_v���eN�ܢ��5�0�[�`���qi'n"�aÆ��0��15��{�[w;^��'��VG����~��0��6�l$׭Ho��ە{Kbq:&���mI��7�\��}��yC̃*�t�s����<$�:������#&�슑��(ԛ�^��X�M$R�W���:��ե�/�K8]˘��l';�$�����r➭hs�l#�)gM�f��!^6Uk�CF���ps�=�=g��:m�γ��6;,���x�Š��y<�ƺ��^�����a[��X��~�mo�H%ޅ�=�:�J뼴}`��3���R�u��C9�'S��,9�}�)9����I\"ڛ����3��ث(JJ���*�yD�>�����4ݜ�����K�B��j͉؇�Q�
B<��;�Y�ߗ��Qc�Q����Z��8��rp��r�����"�c)2���^Q�ڙf����C0I�b��#�8�{�?-��k�D}�9^��j]�Q�dk6�4-�[�Q=�P&����*�sť!���%�i@q�"�e��.����)�I��=�����8W%���˽�W�j��Q���x��P�����3į����Pb<"5ᨘP�jkŃJz�rv���ݾ�]��?>a3j8��]OFM�#����C�׼r��� J���� �E�œ���R|�l�{�֧\\\�̚�d�X��*wQ�U6Q�]���b-�b��pS�Պ[��ó��F�Y����e�ׄ�)��ܡ�N�t{��:7��0:t����<��{:t㢯3����nq1��w�k�������2A�N/xM
,�a�AUEBo�á���v}j����(���M�gϐ�X��G�����f&�У�%qt���阩e�>S0Y��f�;�.��I����ԯ7c]K;5u�H��C��g��8�MLdLRvL��X�q�9=��1�ݐ8�&Q���y���6�Q%���s�`ަhM%M��eT��9J53���1�z^�W�{܈;�Z�p��ϕX�5ym��B�T�VPՉX߄�߳6)Ot�o�OcG�ւӎ�_�=�~�Q�$�#&'��
�̠j� dk�.��龞w	vZ�7�Y</�t�B��N(��PR԰1�+a�ff�~�K݊/T|U������UNU#�,�;��#o]i����דu'M�!�	��+	=c����#czz�c<y/�#2�T��ݳ�dgCnh���q2����V�5=���''z�lmD�2�k�
���g�\9�Sʖ�k��W�Ս>�m�����Wn3�:[��-v5#��6^'�j"ӯ	�)=�t}"�t��w3���@���f)�dP����^�R�r��6w.����ᩴ_T��tj�u{D������%��1e�&[�P ����UWJ��};ڧqTb&��&6:�	����x��2�4`�GMz�R;f��X�/���r�\8�̯u����ʒ����Y1��1z���BC��	��K��&*�<�`\s�
��;cs+������,�R�m:�fo�C#�^,��˕�4D��-{n�MEJ��A�j�M�ْ+!ˑ>�,��Q�2�Ʌ[O��t|>�]�i.�=G|Dj��C����7��E��,p�E#�䭁P�m��wL�B/"B�F_�TT#��Yࢷa��b6�E�=Zg2���^�41�Y����
��-�n0�lQ4�Bk��6�{b��<A��x����	��>�xv��D(Y$��s=����p��f	������@tD�l؅>���(�]�zV^���$ҫB����N�Ւ��}5R.!�qZ�1-�����!�d�#*$��i�ힴ��k{=��t5���5�R�&�W����c��]rd�gk�:mdzç$:зj3�^�z�\���V���=泽�-?\���҆nt��ڶ�4E�Drv��n��[���S��sE����H�ˡc��[ij�@-6�U,�)�v$U����w��g:���_TM�98O%���T����Ȏ8�x@���Y����J#�����[��m:�ay��:�F��g��;\9&/�(�t�ƅ�$ȼ��_�ҹD���ՍP9O]{g��K:���]�hHd_n߂��.��)�_R���}p���{ "��d�+�U�"R�}�)�ά�w`Z�B�(��������슴'�V��=�d0gI����zϊЕ�J�n�r�VG~Q/c�s�b����wT��O�TH���fS2�3m�^�^���Tn9'����lf��~)�(#᲏��YI�t��1����*���:c����H�r�N����i��fKq���1�H,�Zg�z��ޚ�;�S��A>���WJr��F^��x<��
�S��sFy* (���ⷹ⛭��ص�-�=r�׀@g�Sj��W�Y4���o7�imt�	ٲ�]�Q�j��#�븁��~�2E�T�p�s
�Ig\i^ĭ�9�&נgŪ�(�tK��b�����Ѐ��wguι�н1�{�������JI��F��o*=�Jn�󳜱�LDS+���"�T���I!ō���:d�K���tu}�b����X��rl�KW�K�=���~�'�;�iŬY\�ɠ�3�bùfh*�9�f͈��N̨�M�:e�`�Pq�K��3��~����f��ݩ4T�i"�>�pP#}��v2<��gC����l|P�gk˘"��Sų�s�D�H�r����E�4cњ蘟5Y����,��F]�щ7*�%�0-��k�i���.��5C����aÆƹ&�m���\��������#��p�l�������!^ɲ�\��`�GT6�a��w%áOg)�O���}RG�0�<�`$�F{�G�t��WP��u�U�A�!Q�Z�#IgjS��q�u�W�{Cve��%�=�s�Q&
BFպ@�t��7��99՘�SE�R�?>�i����}�:�v)܄����5���䫩�W{5TC^.���j�,1�����R��d�[�k�J�s"���!��ԡ��9��g�y�܄U߱�"�oB7�2�c4�3��,��/6��
�t.������T���s��<�4�^�5n�DM��K�k�8CyM-O^��Z���9m/��;�I�6Ì�_T�ړ��F-L������κ�QZVt��S�
e��tgRwa�;�ʂ�G����w�d���==˱��V���˦A<o )�5�W\nT���l����oh3mʸ��T�s\��W�93p�@%w�&��C(8�������azR�����FQ�m�K#�cq�-�]Wh�`S�����_��J�i/�5�t�>Z]���G�t=V�ɽȩ�kQLx�А������]w�u��`4�Gm�;+k�R�Z���C���%7�w��4l�"�BQ�D��t�u,�T�8f�a��\���(F���zk̊"���i��X"���Y�B42ċn�x�`����gL�2���`��!ח�"nڳ��=f�C��lv����֑"�Y�I3>�(A�Č<��PjbyZ�JB����'�9��uI��YA�A`�:�9*�����u�="���$��LМ7��p5�n�6����Xa��.�yD��rh�3b�E��e]Sq�P�,�AA!�q^7�u։��Si�W���^r�g��WS��}��и��~�����V�����9�����S���f]���vt�v�3�*#m��#8�.�f�]�U��:�ލJE:���@ܩ�w+T�����z����3Hr�Lv!5|�"Շ"�9u�R���^�t6�٬�bc�T����<�S�gp�z��t:���bU7��ȁѽ�e�}rxg���J!o�vm���+���5�sV�T�!ז��R��66����r�Y���V�6�Lm��	K�ح���� n1R0�Ʈ����%3M3#�[Q�yYܫ{U{�e���kj<���H��w|�����'��$K�ʔk�+tp=#���R2�s���nV�&gn95�k;�Y��H��n_�M}(ͼ��r���T2n޺<�ɪ.��f�wZ�`6%��@��Y��RU+�/w<`7���xQaM]):�-�[�'P��q.�z��x���p&R<J�,:�
�R��9����%�=���8��8��>�Z���\�,$��#�/ K)�v9��^�\�%F����%���f�m����%^Dh,�) ����3Ut�\�7md�r������pkR�m������-��kZ�cJ��3�x��:����^+��~S����-�*sA� ����)�N��-`�8����P�����!��_ع��1cwZ��C�w֭d�8�rU��9��P�l������8��I$�J$����pvr��^VЩ|%ַ������R�a��]�zfdi��V �,j�f_D{�̾��m�rL#sb�v�5/��3T���旅M�_�>޿\���=y��P3SR�[0l����Ef�f��ܫ�O^I���:�/5�;�L���%+��W9�/����a��b$�۽�3]�V�Fc���ې�=G����Vrs[����w�SfY��P�M+b���o	�AG%Zt[���e-���%&M�u���E�Ir-��:�V[}w
[xn`�y��U�īd�C�L��\
�f�7u�	7��}58I�yo\w���=*Q���G�\�7+L]C����H��%�eӵG-���jQ�,.�w��0 �/i�48�����/�����o�:Q�[�����:=���)*s��S݄`�8�k�N�t.���v���h�Mbv��wx�ݎ�rnާŰf�t�Xe�ɡW\U
����{)"�&3��ںu;w��-p��M��z�d&�豳y�x��̎�,�ފ�!�Ԍ�k�:5�+	#�ә��RP0Y�Dt�"n.�7�MnN�鷇���J�P�����gw9���aΦf�I:9jZ�����@`�ANs�q��Qn�������%%��._� Ϥ�<�������
E�q$X�4�a
)�X��3Y ��V�	XTCL��,�b��L�g����X(,X���� ���(�V"*1S�2x�J��$X��UJ�E
(�
"�CI
Ȋ�����"�'��hJ�j(�`��;j���@U��ێ�P_�+D@IX�ȱb�v�@X��
HV"�Ȱ��Y*mnj�PX�~J!�X��+uhE�c�PY1!㌀��L1�e���ȰQHi]$���`"�����CHV,r��E��(i��*�_َ�+"�b�}qDX��&5,E�*T%��VbUm�����	�Ym�im�Z��cO�.�ꙭEX���m���@v�RV�t]�;2���tE�=ס��}yaݕ0GOa?f�5��+c�K��c|���}�<�8ך�i��6:;K)q�wWtRs�v4��t�Bg(
z�\oK��ܔ�#[��
��uG)�:���,=u�i]a�&�N�"p������ݑhc=w�W��C(zS})��׹XG�:g���΋mІw,e��,�����(D�{!�:���;q�8)OD.�h�E\_�9-�
w��Ҷ��S��m�WT���9W�
Pq/C��p����F��0?m]A8������8��60�����}|Z�őC�1X�A�0�o����D,.�|��zzeB�o�\��ֲb��ivD�����\iF|�S5t덙��D�BIk&4�����"c ��;H�V���~��/W)qA���t�R\�]�E�ufE�J���|��#8ptײׂ��p~�TrY�<;�S�W��d��^�#h̷��T��Q{(t�؂i2�1��W�WJË�TY��P3
�ᨻ�x6��劼0�K(.2؊4z��R���^��컽�o_D���C��oz�9�R^��_^�y����Ɉ[H6��]����ɭ��q���,.�:(�XrC�����V'vJY�0L%�"���Z����6n��KֲF�v!|ַ�j���5n)�]��7nSqNz�����P��������mp�^�w�1��i���x����p>��"1u�TUr�״�C��(�.>��H� 0l�u-mI�
��$H~�䩗m̊��A���(��#D9|kj��b����ߊ�bSfz��8�CxN��������>�E�,J��[F�ڻ.�=��)@�o�4�
8y��]����֑kv��s�O�/�NV�aF�h݉�~�C2���V� �3����S^�J�o��nK�ֲ�2�4�1�//�\݊�w���q������OW.^C\8U���F^L��)��xyGb�B9�v�T%�1���bdvEzО5j\F(�*�Ħ��a��o�P��粫t�]H�[U��8�9F+�}���J7�2�����3k�f�K���l�↊�X�V���3υ��,���� i����7��1Y'\��˨̓�\�������/)�v�����m�hצ�Su�4�r�={@��N<�1p�v1[���rGJ���3���7�U�eG�kV/�}�z��}C��癶nH�]s�#̣�\�taJj}\,�ږ(�_�Ф�:MU�\��	�z\�Q��k�ef�4K2i��U���Vs<..�k����k�yg���{�4B��.�-��~�u�%z:�"|�]���4`n�W���]�R���TCA
��J����Q�
��Ƚ��.���5��]��GsT�I�[Y�DJ�;!�v �fC�$�EK�2F	S�a�."�v�,��8�����W�_-�׹|~�L�\ |N�L�u��a:�%�ߨ���U�_O0�%:��I���{�gj�@1�"�N�(mK�2ϩ�8f);fhJۂш���f/"�K�#��,��%ם��޺нqUў"s"@�L<QqџD�tLO���ew�B5���V�/�������n
��*Q��B/�]`����4��~'k� �t���l�-0�G=������E�6/��텮�A��>�U�\Lvx�b|=�����l��������{�	�g��~[�Z�h/�#*+�7�(�l�+#J6�;�����}�%�h��5��gz�ͺ�T0^��(!���%n�3���ŊQ�46a9.؎m����0�@�=���ޕ��5�\��%�y� �FF����ʾ��VjD�����ۍ��D%90�)Inw.��6;2~�Oޞ�)�Ii�?jN�QBi���u���/(���<��g)�Q�����l�Z}B�����՝�r!�S����ܽ�F(̊W!��H�G�1�4�A��s%ub�e����n\@��Dp�,��]@�b}z���/�G��o,0fr�v#x'IM5<(���+f��|`o����U��l�
7�S,ױ��ڞ)�~�ݾ-ENA��0��YP�q�WD�����|���,�+Uv?�n�f�exu�.�t�wy�qj��o�b�3��&k���2��WJ4�q�(�=����c�ˤ��6�k�{����4�XJY���(,1��R�6 �â�f�p���v�ݾ�S4�s�k�9ѥ��5��]ҦDR�����ֳ�V�8��q�Y̾�G�mG�}��탔_��Ʋ8�FY�n5����(c_�x.H���Y�~��V\�@g]olo+���HȑYcMb2��f&ۡFO���m��1R� ��J���V^
�=t,%O1]ήT�+p�J�cŨ��]{�{ FLb�uiJ�k_n�y���d��|C0�2�o�.����nH�ǔս�B�8��B�ƪ����\����I^����\�4uyj���ڍ���o�����w����<!�� �7FG4�|15���ׅ{*u:"{Ԫ��m�m�e^S�=�7�E�Q�`�0����-���ÙE��"y�0{���;u�2w}��s7mӮf,�.�i����Ԑȼ��P�ʲ���Ș�.�����ktOL/D,t2�TDזS�x�q�Q��,Mr��h����ޡ���T���x�Gx�p���F���}�R8�v���y��PJ���K޸6�VuJb��U�k�x��0B�T�1C�܍QC�R69���(����b�Ӽ���+���Yϟ���I�8��"iI:h�	ґ��V�V�S#:8M�_TK�$��������uH��q]���Q.���/�(K�A�=b��n����=2y���9O���*��	����
C�q��e�h�G�u�Ld,g�E���;QF������\9Gt"�mqDqdp�'LV/Pt�BAL�����q��Zw��m_����r�wd����VVt����s�gP���a)@q���z�;�o��I�u����vڮ�N�u�Î��D����Q'��j���ː�z�j�2'�&w�]��Gcïj1Y����ؠW*z⍪�I,ؔ���CyS��"��6x���V���u��ڐȜBIt��L.V�u}9�i+�B\�����@�t��,��
�r�t�uiՙ��,��r� t��=�G%{������+f7*Y���dH�(,��4C��f[�}�L�E�H�85�L:����95ِ/W�,��i�8e7�TU��fx�%�Hg	�'�Ee�E���Fͬ�ȥ:eX���s���S6:L�WC�:1��n_	gá �/���3hΠ�I��땼��3 =��]�o܈��*+�^���q�ٮ*\�1Jʜ2�{|�9r����]1���MB �G%L��h�dSS47�C���N���A����ا�A淧q%ti��٥�Y��\D���4�V�������2Q�[��i�-i�G���*����1��E��J����B��X��AU�\���������m8�5��3�v���"�S1�1�N�ͤF�6ߑN.c6�2],[���	
�*;�|B.G/�e�Om
�*.�������g1��c�ƶ��ëv�4���D2�� ���*һ�\ZJ@:��X��sR�v�t���>@�|V�$�����Y�S�
�6�nIX��އ�T��~�.�aL�����^ٿ;�"�fpչ덬��A�R��~_+����a�t��ʽ۫�v�w��Qa��<�����v���C*RU0��P:�^%�6�o�_�S�)��������>���<�^_x*25(�D�$���{9�F7�u�^]��+٭���8r�1B}�Q�,b�h^�<�za��N���ס�Ę���)zћo4'i�g,���]\N��b�/�|~�Y���^]{�YL�&�q�r߮[��=��YKhϧ��9e�X�(о�f�:�?����n�)Us��ϷRW+�/�r�޷���<J����>�"��,&��{.8dPr��:U콎�L�)>�&g��Z�����?��b0W��HuB&�]rITߜU�X'�p��~9 �}ssg�Ov�f|R��U�s��׭x'�'Ny�dׄZ�G�≾�BY����V�iTYpϮ��w:���3�3�a:fuVܗb8X�q���(��V��Xɨ��>�ֶJ��`�bC��:O�n��>��P̩��0�.�X7_��A��0"��6JE�%j�з���pӆk�J�Z_p'M�`��j|�G\R��/)ӹ����Bie�L�Z/���X�3�5'-�?j��ROzʓWu�����
�g�~'R����C���F}�&m���@�4�7[j��݈�Ò���\fԌ�e��B/#�`��. M$��;%e`-��X��۾*+ �� �Y��pY�ϔqp�ꮥ�퐉�d�U�sC	Zo�S��7y3�.����3˼tm����д��ZU,�yh�k�\��VR��a-���s����H�F�p�=��3~jt!�j���q��(/��*�����5Y��*�ek]	�^9g�7���Q��m��n�C8u��S�U'3�'z��c菋��ɭ/ѽ�~���f]Z�Bz�##��F���:1�L��z|��o-�m9x�|�u�ȹ(����Hf���\������U�;dPQ��S,ۥ�=}�yc��ں��^��dA�z*�
�tJ^w��ZϦ*�u1�
^��F�R*Y�5*Jjxq�Q6��^/Ht5�׌8�!et�^:i�	S�V�|����9IV���gU�;��\	����e���V���u֌OA��`5	�Ŋs[���^�]5�NJ�;��S�r�{�j���ʸ��$.U�o�h�����}��hEL@]��PY��i��J���Mk�����7ɫ�O65Iޏ��>
�3V*p�iK'�U�}8Z'>�_�D�Z�j ���8a�3������f�B�Ap�y`�ɚ�(���Ԫf)34������d�`���nU��i��U�t)X�!��C3����_�������R�Ҫ��ip����q:�lK�Ў���[�Jc��#"Ee�k���f-��,�\]0l6gL��Xxl٨�[�rw�� �^�D`D�g|昏�)oEZ>d7��=�0���3���ۓ�^2^ä�N�>�4*q�A�1`r]���xg5cΪ()#�C\�#�R�r㕖��X�.	��i�5��1~(�����	a�!�y������nb��͜i�;�َvyH��+�5c\(�������=�X���	�ʣ`I�D-��Ӕ�ȼ�͕ςty�Ù@�e�L��{3��P,���w�j�8�3]<`��֩�HڹT�}v��͞2�(�+Q�S9x����s|.��
�۔W��ӵ�ѓKs���<.�E�c6�5�n�6nS�f�aLn��hE9��mΒ���+�Z�gR�k^guΘB����Ă�ݙ`��]�Nk�K�=[\ֲ� Q��kyy)�FƷz��[�,�N�3�i���f��i�Y��}�)n�d�M��mT�62��&x��)'M��7ґ���r��*t�>��wݭ�
k8M�iP�
�B:4�y1�).�}|�/������nk���7hv�ܴY���:!��h�q��L��&Q�@[�F�g�Bq�z���	��vEɬbC=�Y��=�4,��'Lc�P�d�c�i���Eo���:��]=����1�D8s�N8f�4�!Z�j�:�fl)��],����{_��s�we��v�`���Z�Ѭ|�%�xo�ʖyx\5�/��U�����eK�so4S��mM�k�����E�[1��R�б(�����C��!��T��ݨ����F���.��W�{C����oBF�<+�hG�B��b=z�y�u�*��p��9��{ֱ^�N�gZ��L�b�1��"U�o�&l��n8�̣�[���5�ʾN��"���7����7�Gi�������@�ʊ���Ρ���*Ze���b�p;�ǰ������(" -"Nt�������0KY<����&Xf�����%o[*yT���Aq ~�j�ʵbD@X
�Hj��C�ꆶ�DlegD��wR@D@_I�2��6��[]��~��7�çC�4�Z�*E+.*�}o|^ua���_��������w�׿@$�44{��W�����D���
 /��IZF���$8�_������?}T��@��9�x�{P"N^ " .>�yOڏGT1:l4��[�B�c%����I�=�ڐ,���&z�t!���8��1:��G���v�?��r�" ,gh�\�;jz�r�鋀 �=P��͋DD)��Jms�,ҝ�v2�^��T�w�������I�_�nm��WS�=��$=ݒ�*��D�f����|^g�2x�]�����!��l�%�.��Mw䟩˰6}�\���6_t�в���|{K�u���&�����zu�R����'#i�"�x��8xt�C�����g"�h�w���"�ي=�" /����_d'd���5�(.��i,>���EE�se""`|���!3�2UQ`��#c"�p���Y�ѡ"��K���s��yO�1����{5�������@��v���8 ���_��Fǳ`!<φ����7�������'oV��Yc�t�B7��OS٦!=I��R�����������tnA��I�U��{�	�" ,����la���O3=�O����&�������hK�2!��I=\�P ���9On�xo~����2G�#��������[_[��" /W�`Ϩ2��"��K�;�	 ٛ�p�6��.7��,C֖�Hm�!D�X�`ڃ�<^�c�:�D@^#��R�]W����epBʜ��Җ.��"�>$�٧R:w9?�]��BCl��D