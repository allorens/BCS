BZh91AY&SYR�=׏߀`q���#� ����bC^�     =��P�I@ (�H PP@TU(
�P� �)A@@
AB�(@� )RJ vj�H T��"�%J�**��J*�@�D�!�IP@��(J��T%!**I%)(��B��*$����T�%D�T�� )B)PT��IHJ��JH�H�� ��T�J�Q���*�R�	JDUR��B�;:UP��j^�
(J�  Q�j� d�١Y+%���*���UPj�PU�5*��I*J���%D)� 1�Eh i�( j0��l   @ k@ڌ  
�KP  +5�  mF i��f���;���)D��ID` � ilC;� �m� X������i@ �� �4L� A:��@�88  ��4  7!!����@T�,  3���PO8 �G8k��  \���u@ �/p�T5V �@Q�+AA5h 0* 
0�P@� ��!Q�   ��  &V  XA@A� -+� �� ��M *a` (#( c (�� �EII� C�  U�T��X  T�P  `@�fV�P fV ��#C ��0
 � �J6�c�(�P��!R(��  � Z����0  6I`  �L  	�  #V +0� jD�)` �JE��*$T���   8 l(�� �� j@�&�  ��D���UB�@h��%Q�IB��UE%� n ��� U� ����@"��Rh�
�0(���PZ �:D%*TQ*QN ��e` j�i[eQ� P@T j0 (mR�b� 6�$�e �    �A@50T�T`F  &��� ����2 ��  Ѡ� 	�	� L �'�
J��      IMS
lSI�M4�� )!3RH&�4��F�� !�㦺��j�Z��Ӭ���iy�&��]�/(�����|G^�9��=y� |~�TW PT��P_����* 
�q��#��a����Gj��� *���UW��D U���I��C���
*�����9@�2'�`O�"}�)�Y�
~�D����2&�l��
m�6��aM��l)����l���6��`���l#��l)�T� �yeM��Sl���"r��Sl)�T� �:eM���yd�ۖ� �v��A�
m�}0�l�d]���l	��
m�62&�eM�&�l��D�*m�6țaM�&�Sl�6�l	�D�m�6�;dM���Sl	�Y��m�6ʛaM���l	�D�(m�6�2;e���Cl	�D�(m�6�;`����� �vʛdM��l#�T�*m�l!0��Gl����v����� �xa���Wl#�G�l�� �v»aL�A�c �6ț`��l)�av�a�*c
m�v�;aM���Sl����+�T�"�v»e���D���A�� � �*��QGl���ANWl��P�*;dAv����� ��"��Al�������Pl��@� <�;eU6���� #�AGtH
����E� #��Wl(��E� �ev� aUvʀaP�l� 4ʻe���Gl�� �v��*m�vʚ`���l��T� �6ʛd;ev`2��l��T�*m�6dOL�6d���L�:��1��}������1|Ƨ��aGA��J�w�Q��i�n��%Pq%yٵ�,P�L�9����O0�(����*�o5E���l�Z�_�Y�7J����
�v�ˢrm��onȬ؎��%KͫsG�n/<�e4�
����� �ǀ #�+FE�y����P"R�T��wB^En�Ehf�T�]���Ц�H[C3H�QĎ�Ӧ�e-��m+(ӵ��/h�9�ֻ���7�kH:�!K�V�aKQY���uE&�.PJ�ha�rXÞ>�I�{��5�P
� �l�6���Ciӄ�y�+voMJ#M��4����{��MF��f��'n�x�:�YP���!�4���J�j̤�M��=fƄ��n�ۧ�s�1�-T�����!��5�34��pYn�xM����v�F��:m)����K%��-T�Q��<Ih���/�9����4�b\M�f��
X�d*�&լ�P�)h5���7��Vm� ��ˎY��HG.�
�)P����MX'�5��-�d���M�\H�
�r\A[��4V��؂�2�T7�h����ǚ�s6�\��@�M�v�NÖ�D�v ���66����#�1���bęhI��d8��kG��v�[�JZ��5Ycq�.��$f�(ܕt�)j򈫖��u�������-�04)U�1:���h�`��r]e����n�\Z7Cu�A҆[Yb򭉩&i�Ҧ�1����[1ڤ��	T�*��L��]&)�w5u��HYڵ��Zi�y�����X�#�O^˚q��w��x��{�4�H�X�ֶ�7����6��37u-6r<Un���-ʏ�y�VPQ�o)��u�gi���S׬yfk@���;�8kmYz�V!�V�
*,��X�+��7."/��+"浚f00�&J�k@e�B���c�k(�+u�*`�;�!��� n��h[�d��{3[�M�4i�zv�]ZOpӢV4���Oz�L��p-��_X�픬pm萓K!�z�GL�h�J�ފ*nk��Г���Q8�ʳ/�JE����ڷ��՝��v�x�8�wv6!s�Y���W5a;VpF��.��Yy�9�<�R�'漼�CY�N�7Q I��f+:�Zv)��\G�0�7j�j�L���{2�RoU�M�=s0�kt����*�$��28Iu1,���e[�6MZ��j�QK�]�Yd�um�WYm�>�b=Cq*���F�-hⳲ�ehvNXr�t7W�j����tTE�8���/�^R�T����z�wZ�^@�K*�`��]�A;X��;���`5���-�wM�5�pc��{WP�j�#�Pwh�Y,�Y����n��IkRތs�ǶK����R=��
2G�T"�$�tΫRU�{��eT�*�RCB����i�U��{]yƲ�qC(�z�] ��X�|e\5�0V������ 戳q�MeӔHwAW���P��5u�si�S	��Hm�OVB1�4�ٕ2�7K"ҭ5�����S�M� �$K��� X�1 f���{�������̦f+:����u���4��f���f���I�`�Z�����&������T*� �%��է��4��<WU[u�d��i���D��]_��,�r9v��=B���h�.ڗa!��fbw����5γ����K��s�z�<1��2�.���L���n��v���We�k���b�`bm�oe��0�ѭ�SE�g4˙,^2)YeJ�'�f����b��jf@k}�c+t�V��VZJ���x�����C�2���f�8�CVvۤ]�k���']�"%�X�GV��\y��ڛ��ů,�M=��E;h�����%�9J���x��4�2byw{FH�^
�+;bb�K-�+��۵�R���p�C�rdq�K�2�����)J������Sn�&��ˤ�[4���ư[��,�*��óHX�l+�w�wFm&������Z�ã�+0˥F�V���Bf��&Vi�f�ø�-Ee5��JM�2V ���{�f��q��I�>guV��V�㛶Y��7�e�*XD�z�F0�94��«2�i&9���ñYۡ��)�N�b'�PȰ`��y;w�ǔR4�wV���LY��X�);ȔlїnbnRמuxc�N�a�-U&��*ѵD�ۼ��t �V5z���)�i1��S��w�s``��6�U�b����W;�L�M0�n`��iU�F����%JV��D�i2�H*Dr�;јiI��b�n��nj�ѫ�$�4ӎ�a�7�� 0�J�6��n�#lB��G���o҄.�˃H!8�����{]鎮q���F�-��or����aT�vD���͈+��9��AR	{f��w�Q��Wgs��T�'��L뼙�h��v���IkL��b�&�Z�%V͉q�9�5vq��[�Eq��ĘGv�¶�^�X��#A��d�˦[.QU�N;*���X��yC$Ĭ M��c�e�2c�jJW.hX�.��t1{k��:�b�Y��X�8�-�vɺ.z�$�Q��4�.S� �3�')�<m����\�Χ������F\��Z,���W�$f�&�:j �*r���s4vQ�@M(�Oj���oAP��iPԮ����G4�.ʶ�)$q�˓h��kh�*����]�j=�s�Ùhݷu�Fۡ�ٙ;ia�g]\6����yv�0̭f�cA1Z��=��2��q^è��N�2V�f�k\�d���pnZ�l�/r�m[����p/c/bZ	�	�c�ܸ^m�H�6e3V��;�AIP�Kyb9��~��U���fmeM�l=уRn�U�������^̕.[�N��7�^�G�:g5��)�HҮw\Ad�gz���
�ͱ���մ�z�V�#H��
��l+�c��a-�]�ʣ���N�7c�A��5a�*�J�32ЇUՙ{s]��1&�34��2\ -n��h�5u0�Q'���-���e]�qY6-=�U��)��w�p������w�q�Z�`��{�Z
pP�4lx�b7Ia�Eˬ8�WS�y=�7�T�^����.�i(*hǬ� �J(��*�#`��E��i��ֳ�ZU��F�%��>:�ξ��ioH�Z+kt��Z	�l���,[�F	�v:W@�LPZ8D�sw(m\w%��-�^Baħ���[AU�j�*d��cE�[Z�p�Y��f-�[�]M���`:ݛq6��^
�Z��sK����{o�[��ui2�Cr]RK:�`������R+�a���y��W|+d$��kr��k�Z�=��H�u��e�׌á�qM[B]
�,"ynY�BM4}�ˠ�=n�zq��w�@�kbI�G7����CV��[��C�RR�]�b�����{/V���_c{�pm�J��vH�v�y&�	cԬV9�S���ۭ���:�v(v�9���҉Q�J!�.�\^n��UH>��^aI?�0� K.�	Yie�F�bdhYf�z�+��
�\M�Ws\�6�*�d�&'��̼��7m�SZ�dc��bVn<�Ja��j:]�0ٶ �`&�ݙ��Cm@��kr�ehޙ�R��zw�j][�z�j�ת;s��-�Z���Wo�W���|9�@���� Q�_lɛcs3J[@���]ӕd[�h7���]l4�k �W�fa`��&�$in�P�JA�@�z�HE�w�7Z����,V&N0�vs%7AJ��,�/A�[��Q�#x�.\�p�G�\Z��$�WZ��Go�-�HL�ۺJ��HWD�"Ms (�,����i
2^ج�f=#q���ܢ�
�q�J���U��ؚ�Y���0�A�M11�;1�ݥ���̱hA,���dڛu[��Tw�1��i�e�cJ�%N��#���ՓXַ��ŊZjTy��/U��}r��e��7�/Z�\F�� hy�p>���	��uB�c�wi��#3=���v��Sc*�T$�QKu�kb�
�W��XNe�Ø�u��5;Z�7.��!��B:x�F�H�X3q�˫b-I;֯MA2�@m����/�a�JBa@Ƿ�f�7��� �,��"yXU񨴼�SUf2��811����:�m-&�Wy��8H�;��^��V��������ذ���������ܒ�n�i Rf�L@K���F�/|6$D"�_X�c�eS�~x�����%��Hj�yr��R�in<8��Y� ��'B�h�8�A�Nh�-c�R�X���]��) ve�Ƿ7��kb��ڗ�2Ian㙁���4�M�3EL���2AUVL� n�1��K����)���E]�u�M�j�-G��@���F��-��FV�nX�::��]ۆ��N���U�^�G�DӐ^ݫ����A\����R�1rE.��%���:�u�����t�e�m���|�V67��.�U����/:@��Ct�O*�,ǧ����24�G!�.B���ܻPֻ�9/6�8��`m��ׇ@�t��u��3P "���Z��jY���iJW�I��
C	��@E�t�-���L6+�n�ŝ���e�";Q7�f]�ڹz���X���՚ŭ���צ�9w��M��h�V���,�bYkjT"3w^l�l�/i��eE����sw\�̢e�O.��`!����5ņF7k)M��2ܩn
x�=�0L��6B��v�GFit�)��=6e�×�t�PIӘ���a5���X�fּ�C��RvD��=�vJ��3,�!�XP��Ee�.�ˬ�.����^�����8F��7*-�{a�770�0�F�[)��2�^���n��=JM3ɟ3q�n��ʑ$V�yyc!�8�5�4ܮU��ۣh7���͗Q���.�[j�.U�)^yf�!P��TAlzG�i���Vi{Ca��e7�������jřrLt��u��iڳ���p�D���˵��6�:�b��z
j��n4v�4��WH�+1	Cu �+%⒍���+k�,`�j��j��}�D�V�,Ls& N@���(,˱�^��ڊ�T���4��ѳr�[����w5���I�hgst��K�7`�����K��On.e�������e�t�]PY�WkKƱ��a@*^�=jl;��H8�	Yy2M��+`Ŕ6��Lj��KA�ڗ�J�D#jn����d���ڰ0�ec��l*ҝee���͐1�{H�(1�B'A@���	�'� UA�pZ��l���F��wX��{���n�CG=%�*���(<��*�uivk�F�k��_0ͥOr�-��e�;�	��Y�VM�Y�y��e����
�<�*)*�az��q�NR�G5%�M���&�ó,�ݣ7�)^f@.�;1z�X�
f��^-�/	Z���jV57Y��U"�wr�[&r�e��wkp�t)��V�j��������N&l:a���F���g(⫖sfK�e����gE��.ۗJ��N�d-��B�i̲��T}�n]Y%^���7�7Kv��͠Tr4��U�i[CIᆯI�k+H6�+<6�>%�n�[�'FlBi4��`N�؂�'j���07+0�i�g�P�^�l�X�L��ZJV[ҩXO+,mfH<>�ؒ�TҺ�ڙA�7S��J�MmжZ�=Фm8f]M�`f�ų ӭec�m���<J�f�%n�2����@:�����3e[Y����ˑ��m�i5�lĨ�޻���D����%���yB��D��[�ϗjL2����A'1oċ
�5uT��'j��6k*&6t@��`�y=��sV��$e�8�MV�Djy�j�fC6�&@��ӀH���ձL'.�=���m�,T[b�k�/qÆ���)cZ��l�\��k�776D\���d�0n�-;�`ee�E5J6��F� �rA�4+!�L�-T{Gt[J�㚖T7m��t4��� 
b��O];�U�c2�qat^k���*�S{H�.��7-������Э��c�(��M��&ŷ7n]hi�G1��SJ"���)DPP�B9X��s)VX�fV�тfJW�CCjKo1a�w�ͺm��j����!c�^���%���6//P�t�,�b�U�FfR�V#�%�Y�Re�Ҙ+�̼��D����66��f��`�|�/O�3��Z9ڠ��ͦ�;z͝:��0�e����w�Z�4�O�{(�oQ�4t�j�U��E��䬥��ڽ���7	sSNkF���;D��J����r�3/HKQ8He��T�7M�ŋx��w�!�'u���˼Żx�^:��-����E����3j��ɣ(�C�t���b�ٔ%���M�-�jV��
�U�(Y�L�[�n���j ���P�.<�&��.@��Y�t�u������ɔq
5���в1�ԗ�Q�D�d��CHkc�s���jx�Z)���p޶&L�z��I"1+֞D���q	c]Vk8��z0Iw�~�Y�rJF����b[���;�0��0ن�$�
n^J;xͫ[�pVΓ���x(���'�j��AuIu҅�A�� �����r�Wd�������ٗ�v�U
0#Nݟ�
��i:�o�78��g;�v.�P�����S�e�
b��#76Jw�b�,E�g+:U�
�6Gfs ��M�l�6p��N��2]�X�ԕ%F\�.��]�w����x��s����iP�瑯��">�)d���l�NG���+)��1�j]c�
�*<�iF��7�
�w,<kt���{u��v��U���b[A�������B�V�[I�Y���SH���$0�Ô�cy9}2�Íb��:M���ƓZ�|��GnF�mܫg�at��RY�w�1�T��28�5˷y.D��P��ެ�w��C�zQ7j[٤y�wa7��������LM�_�y_��W��~ ��F0��d>lJ��9�,1�DDDDDD�I$�I$�9�97��� ���[���G�5ǑmQ�J�/.�]ѻ)Vt��A�C��"��)i��I󃩵X�rIË��]��{xe�O]qH�
�c���܃�z�g#�&orm�!�i��u��8�3��8�mޜ�9�r�7t����C�U���d�oWw�Ϟ�`�[Z��S�Ա-&��J F5WC����;#�
v��wB޼9Ov�62����d��b���ܓ6]��ïB��Mٜ�E[����ڤ�f�ko;�	aW,F�o�!'
�c�y��_p�V�ͯ�훢��r�vBD��ѫ�eh�4W[۷���zʺ/���`�(�r��VxM)�;:���I_1,���򙔟��W��z�Et4��:�T�*��W[96���ɞUP8m����]�r���,"��]��*��8n�ے��%��V�˸j3���F�o�u�wo��Y��M+���;,������GG
pQ"쥦���1r�3u5�D�W�j
��zz���sm��%�]R�Uu�HEe޽��C���A�kJ}���g-{2vuEFa?7�A4Eϳ��C�OVe�>2�7:4��g�K�.�/[ѩ�j�u�������{yQ�Vj�vm�xw+��q�{5�4_����h	]�Ua'���B�U�v/k�	g�Sr�"{�3��ɢ�l]D�T�S�W6�p��$'	�������2ح�nb��xo!$���\������5��Ҁ�ç���l8;J�:y�gs)b$�|�v9��#�Qy�GW9�C�����Z�sT�,ܠ��]ݣ�*�oMv����%WZJ�����>�{�cѾ#oʏ��]�N��F��ɥ�5�ֳ�:��k�f�̷�ʜC̒�u����ʬT�׭m[W��C��Z�
�m���ѯ�Kl���Jdf.�=�GT�qN ��V��fQ��C<�ƾ�wu��S��b9��'Nā��F�ߧ�Ɖ�,�9w�J��H�CK���ל نh�co�4j6n���WYz�ƹ�}e9r%�n�f�RGcη��`�PB�!]�4�Y尜�f���0���Z�Ӷ��&�s�f���ЙW�9�J����X�L]n�]�ރN|��>�9[J�k�I,[kb��@�\�&�|%`,T���ͫ����{���S�^���N�Ρ��_�S�����Y܋!r�Jq����b�ˊ��K��h�k"����0Iݏ}���\��b��Ά��L��]fF�q9���,<$9���%��j!Jw�3�]����9�e�Z+{�h�u��;��M��G-�Ki���e���n��[0��Fi�����T8R������l�K�olymfC�q���f�\gQ�.�v���X����y�t�w>��u��Ds���T�Ձ"��Қ{��
����oU� ��V���Q̙�u^�/����c�2%^2�bD�9��M���iλ�ՠ��b5�`2���J殙��"�,\��i�ZȻ�^�RZj�T^(.�C|
u�:��ⷉn��%��hxk��!s³zMӷ�rU&5�N�	�v��(q�,5KE��b/q�@]Ť���y�q��&Om��o{d�g5�c}�l���[�����Ix�1e�7��i��LWT�p�j�Hu	��lr��TW)��r���1�����ؙ��7���m��W�5�����yr8F���oX�x)ȉ�^�.b�a�R!�9d��uv�R�*��{5�cz��X��
��
T�����!�
M+�96��gvl7�K[�r�wA��G/��Tܼ6���N�B7�]�����
�m��9D���h/t�6慧34k��u�zR��F.�n�£%Y�d/v�+c�ﳦԤx.���﮳S)�j��^�H�]HN�h�K�YĆ����t�|�E��Q�ѥK�&ҁ�B�p�5567�Po2�i�]�֟;��֛�u�����M4��q����5�Yd��ĉ�-�I��k���H�e�3C7YMܻI���=�q���1�}�Aq��r���.�qCM�)F�fk˒���R�z��rU�m*� ̰�w��ԛ�E�V--����S����j�N8���Î>�[��w�;�L���PZ55�6�b.��:��o��v�H�%��E�Ww�p�#����,s/���Z���[���˝L���뮕Έ�2���g���c�����x�&:���VN���AH�����M�A��uj*�a��K��/���!�2eNY�v霰��e�u�M`�[k2��>7W�Ug:#cm4���o��><�2�Ɏf�.�!d��]�N����dl���L���5�Vi2�� ����M�(�:+ҷ.��t�n�S��Ϝ�f�	��s�$��w�� �W�k�9H�U�J���W�v�8��/	d���+*�7y��{ Z�"�M�#�vؔK�&*I�)����E�7n`��ج+��O��)��o1-	�(�cʄ˯�ZR���W\(�uەb �ˆ�_:��F��z�s[����P�����+�хmT��U�{���i�f��U�C`��dRf����:���6"�Co��o��kqgj�è�O���fp�n�t�Y��V�V��+��ռn)�.tں��76��՚w�.�#�P��Vl��̔a�Ā�Ϧ�9�s�ڹ��&:��.������)i�Rc)�d��][�����5��AwM�(�8ʨ�A)	���Λ�7k���<�t���΂[·�����괸�^�F���/�J{M��t���.�����q����tm�����.�&ůIIM�K�{F�kB&�P�)�hp�)�{�״��6-�(*k�;�M�ڼRµې�Ƿ�zu�S�.p��,� ��o���S��yyT[�����Ɠ���l�!;{�v z��;��l��;�ؖiM���T>��hmK�՜�WA8;y+8��w��Y61�x��p�C�;�z��SZ��zNP�[��s����g���b���T�;e�}�n\z���x[�KZ��	7��t6�s{"�+6�I|{�lV�!H��W�r��2L�#k�u�5wa(�ϸG����I�c��3Ep8Q��t�A�d���x/Z���c9�L�d�l�r��K9�u��|�+�4�W�c�{T��k5U�qbh���gb0Y=�i4�m�u�V�|���X��j/@)�b����7�T�(8�f��wGK7�ڗX*PGZەPbS�Xg	��p�-��avm��x�6;��ыD^}��1צ��Z�2�Ic��ɶZ۩��0�����z.��p����������Fnc�)2���N�M��fU���t�|��[ݠ���|��pD+#�Bn`��>�Uν��ٝ"�Aq�����֬f�+�_̫FP�}����h7���;�d�3[�s��I�8�h�X��~����]���S�c����;�;mӵuw.�{	6�ͺ��o����r%�4%Ї��WnsS^B豭hW�s]�,�4�Z�If��E�h$2���4; �ӌ�y��
�m쮥f)�1u�\�p��ww�rgJ�u'�]۝�jO��@Huu�@�]ӂ���S+@D��U��8�i��p���s29Dos8��V#��ɓ��!�uJ=Ɣ���t�Oi�����v�}]�����a/k������&��bt9���Twl�T���Ъ�h�kd0"%\�%S:8l�ۢ��,j�Yɏ�]M�9�Q)0��ːЁ>x/*�Z�EuHlQ˾�JJ���@�b͞�V��p�f��/OrDT���T� R�hp�ݭ�=[���6�"l��bal.htM�*���cYd;9]�+�.�t��񨫎ҽ��M��M��w*��fX�ޭĜy�^[���8�4���v�*�5�x����)�5�ٛw�X6M{e�6ѵ.´oV�8�a�D	��9���/�����"\[���Ѵ�,ׄ(�w$��j[�+�.�c��ۖ��ZM���v�:[Mj9�v>E���9��헓�_i� X�pf����8r3F������*og�ٴ���ѫ��te�<�K_^9���t��d:��%n��a�aT���h��� �ҟ/m�q�k,v����IJ��ps�WWK���H��a�t�x�h�&�b�S�v�Z�[Qk���}��_�f�*wNՈ-�}��Ư%����SCn��d����Zm�	0���u
��Y���n���$��[y)o�˖͌6�6���'$��� �wu�[�捇s��j�92��l�t}P���n�#�v��3(%]�J����Y�p����iGy�Χ���[1���tj<���YA!
�=�U�+;,o��,����g�h�%����j�͘�{�+��To��ۗ{����Q�
��\X	+�ň�u�f�nV��Z�&t�!l�w��CL��f�s�ڻ���w^��(�&��*'/{�
֮�n��:m45�3��*�P�U�JaV9���}7 ڢ1v�����pX(DUԠ������7UUg��s
V�<�*]ɲ�Ǹ{����@�[hb�7.���l�z&�͛7K�����0�B�17���7B�b���S���U:>��N�R���ԮZ���^9���-�NQ�ote_>;C�݉\��0�N�toweZp�7,��k}�+ �B2k��sbHu�39��]���٤ou�IK�����L��V4�ou�1ݎE��P���Z{��]R��J\�j�!�^>�+.Z�0����9ѻǷ��,4�Q�f��v�m���fs�>Ø�h�|�X3B�{�	*T���&��.�7g�$-�&�T�W=�IN�4�C0��h��rg�k����i֫F4�T�Ucz���`ub劫 
��֘�C����\�5o`�S�'�e��������*���a�l�<pV'Y�<U��KR�]$��������MW<=4d�SĶWjnS`!��3��.���-��U 47�n��l�b��/����iM�Fpܩh�M�g]�:���	R��R��լ6�k��tY�A����[��FYV�v�ny�c��y��J�(Pue	��OV��:͞���S%-���n_ �,�b���ۋ
R��!n��0%\TF8"/(k�}V�^b�n����5: Hܜgx`;K�wA��ie�c[wۘ���T����C\�ܳ9�`ۀʀMR�Yf�kx o�u� �/�k��x�rd5x�P#Y��{。����E����	Zs>1��+NJ�7qZݡmXY-lńv�9�4<s���9gZﾬ|s�h�(�m_��:�����N�
Pu�y��&c\�t/��'\Ega��݉�5��/7D�o�\�κYA^n�v1,㩳snՍ۸{d�R�C�s��a;	����r��tu5'n�d�=z
nƠF���d�D��ݽx�C#-1�is6�]��\4]5��Ў�z��xG��Wq�a��rKr��wt-7�Q�݆�թ˷Υ-d�Fo����O�{����mm��P+I�6X���}P���C���]���Ί��ö�;�d3�	���#�x�P[�"��1h��WJt\��V1Y:�&0n�N�ʽ����e���+�Ci�4S\Vu�Q]��e��w�8�NXXFt��\y���3�;s:��e���c�Ǜ�(�|3{�6�і���}E�#�ۯO�i씈ƢQ�����Raj�h�9��q�%�w/��1�a��^�i��ƭdZ2j[�gA��P{�N�lhRBmt�J�s(���Y����6���pm�֖M��8����p�C��[��0m-�R�S	1�%LM`]7·k�������N�S�A����J�j�<�p�.����u�;G6C�ݑ�G:��.l�v�i���V�]�_��fȈ�~O{J�K�Z��4��ۤ%ͼ��WV���u�{7lp�j�۔�,?����وF-&�fd���nj��#.`;��A�g<P�Z43�)�1���� ��:�������*���'>.C5�9-N�:]ۉ�6��y��_`�5�!�^t��U�ӐVw��_N���m�b^	�3�1�{�fɌ��<�4a��t��35�^O 	�ͤ�'NF���a�cV̫��#�e�ʫ��(�Zn(-�f�i���� u��/U��A5ǹj@	��p�p�\��r`���lb�bԡdD`Y����c������xL탪��-ͅk��N_- �`�6ƞ��i�6��~X��J�z���hѬEḱ�o������iC_vΜ,�P�v1�1��X��5d@��8ئ�n�-q���}��j�4�Xge���3kv���ԕ-�V\�����,]�Zr"�Cuwh�����%�>���{\����&�t�{�����>	�nΐom��,N�6�]�j��՝R�����ܜ�HX`��\1��QdW�$Q�'dv��7�	�ӝ��Y�M� �iy�m�:�+�	��ۓ��,�;D9x�8﮺K݈2oa����U�bC��fP�FԆ�G[y�e���\*�ُmv��ckD=�]t^s�^Td;]l��4�KO �U>��m�nm%9q.W[\���w;����{C�͹����<�˷/�U����sGi�!`�![�RUg\����eI,�.C$�t\���l�c��I"�u{�����ڦ�B 9р� jT��L�h&�4Q��N�*%�Z�Q�˫D�$ L�c���G ,��mP��$~��Ĝ��T�S���SeӔФ@5N��Q(�r�F\�dщ"�h��Jo%��4R�	�*f�@��t�Q��[�r��$|M��|� "��D4��a�҆<~.R	�*�T�F�B�!�1!%#D@����,�Yo8:�+�:+Yf�]~� E�~��?7�*�y�/���Ч�~�EDEI����q,��YmY�|�iiY��
H�ݙ�F�/��kZ� �o6,Yk/�����j��u|3\���l������������sv�Cq�3��Ro>v��Y��e�X�m��j��Lm�TC�f�En���d��غ����w�\����/&m�5�Q�zu5̽�+fbLQk 
���,>�Ve=t8�A�R幔ٜaz���c3���w]#OCV�U5�7���8�����ȷ�����(���8)���ܨ��Lݙ�1Wb��t�e��V^ބ��|��<뀸�-T�����ّ��5��e��Ğ�}���t�.e���ז�o	:6�1n��CvމE�p�a!����2�o]H,�� �B.��*u��a0�RN�����n���L}A��.��8^g��1l��|�ڭf�w2	��lW۸a�@�e[��C��qj,S� \o���dk3F��,o9b�^�+�EUذq��9TAD� ��囼x�kMP��:�wZ���3�c�y�5m���� s��dɹ�aҔ?V��uee��:A����}�j��sX�u]jBXi�:7�w�e]�Y�@�wAhi�x�嶕\[׈fkI��H�w��cbT���&�΍�L���̾��Tx�G6�5��cv����ܲ�U��bv�ݦ,�*��}q�9>/��V��j��<C��R�2�3�Ļe�=�E4�Gg
:��ܪB����(����>T��c\���W9��Y�8�R����ҧGu��m��)k�p�{v�KK�����N�4��]S�uCԥ�g��]�]���u�Ь��r�fe�ފ1���ibQ|!�Z0�D����%��;�՘�@�9��EV.��"�Cٸ�1Y�g1�:��/4�֜S�WM�K{yq�W[�:�6�@����7q���u��n��Ұ#�a)!���e�k������1�d�1lԨ_@0��;kҸ�$�z�v�n�ŗ����y�;=���U��O>�-��8�t�3/Gf�
�G��ӌ�;8h��Nؠ�]�gU����vd�3�#3F�#xl;xq	.������&]{2�b��d��p���]�rC���x$.09��B�ʻ�m�K�ۆ����sT�� V�w���q�;4+x�;ܐ����aaZ��]�&9.{�ۢ����4)r��L��1]6ߒ��%�;X}b�^J�CAs���[��HI
}��Cs��wZ�N�}sINY�f���z!�Uڐls��fGx5��ï��B�:+���uh�(+S4{U�kη$x�����AKϣ4#��B����7�fXu����+�/Iۨ�"r����4El�"����<6�7h�/�]�.ё�+r�h��vIP>8EN�hܕg��9�=�F��Ғ��b�עS��5b�Y��t���q��ØB�TuԈ����D����Z��;[�ucl� ��%���DN���YD�]�3=؍C*�R5{b���h�N�uo������7��j.��a�Vআ*��\�
�Y�P�1s�������o.�\�F�=y�&�+��)`���mw.��ҍR(�ǘ����iS�c���v�^T��R�-e5���N�ۯ�ΰ���b�J�q�n���HQ�z`�{�$|�Yd��(�ұ���o5��2.�Ʀ�e�VQG�u���i����u���h��vV��JX��3w�4,�ҭRa`�Y�*	T+E<�Q��O�U�5d�'ݤ���c�1i���Úr|:�Φ7I�)�dJ�<6����>{p���G0��k��i�����ޑ�gU"�%������X���,e�����C������qa^I(��Wy���5yQ��3>��9X)�Z@Z޸-��g)+tiRc����%d�Y|�]������
�JႵ҂]XB��-m�RMe��r�C�P�kJ!��4p͙�Fi�b��TU[wuGf��x^�IC�g[��1,tG��Mb���;� ���+_`�%Ƭbl2A��u�W�$�*,Ʀ��hs}ιf�A�(�l�k��&���J&��Jcf�����v�2��@�v�ں�`��N�ڰ
�z;`�{���C�y׆QF��QΚ4��6tY���9ʶ4�`������M�8('RQ랑G\<����M�s^j�Nc���ui7����\�����q����s*t�:��a��r��QR$�Zo�7��e�?�� �Vf4���bh�r��cɦ
�+tj-R���8�+	\��S�ys"�vwze7��vPb����.��k�n�{Ɋ���J'����t+Bә"5{��cxT�bb=�A�[[��oc�2�s!9.�s�4�IVec<�y��H�Q4�):W[j�C�ѹE�bmi���A�� :��.���(�\�EB����9�e�#�=���j��ёkp&�g���S�c0�;Ȳbp�mfǢ���gK��Nf���LN.� 2���D���HZ�+Y���5(�lֱ�z������v-��2������*=��:aPe1֣ ����.��r��7˫#3_j�Ou�\⑷IV.�e\�t���Pj]W�^�uXH�b>!𨃬h���B�xVB,��4J�K7�X�֫�������ߴs4�Ὦ��[C��MOe��H�v�d�me��
+�uڻP���-3�݌�����8����%�����>�qU����Y[D�9�'#U���}سT�5$,
G.΋��d�|I�;h��V�|�ɪ�����k	@��#��_Ga�����1�M�J�G�J9��y�0���6y!�BX���V�Z��IWd�Y}E[�䉯_veMǭ�,�n���x�P�����Fv7��F���x�t��!�"M��U�ۣe�=�`J�����Vm�;�F�g�n��Р��9���I��'V[�[�S��)-�ٶB'N�ۮ�;��^H�"����u��+�_
S�.�Y.j�&п2[���r :q�3,`�pVd�}q���ج�]��Z�H��7Qؕ�[��2�J�IxMD�k#OR'Ƿv��8)%d�V��ux5�M�o`5 :�n�Lչ�y���2�
}�;2�h�M
�Hm����\�����W�{��Ǯ�vN�+%tWqLhUU�cU�J�ۄf��+��o��:���"lu�,(�A��h؂=u|2�8�jqM�0o6�-��Ɩ�^����Z��E��2%���Y�1����L�8U̽J�#������r�i^��b�[�]���`�V0=x�P��Ea�W���Ǻ�6�F�כ��/M@!��H�����*�)�T!QVv��8�c*k�.�1\\�u������rV�k���=R�K��r�Т�c��z2�2��5����}�Wy�Is.�X$��c��T��:j���շ�Jʰ�tWU�KŘ.wa����Q��;��sY��TBv�
�ɑ
8m�����Γ���=�$�k\�ނ��y f�b�j�"���6P�޾�՝S�}�8�H�/:�,5ƮKRn�H`�(��A��]����jktͻ|�b� ��r"0�4/�ta�1;�m��;����+���5�9��˛=&��|�e�3]�B��%_Ҫ��-`4GQW}�y��x�Ӵę�.
�{*�{�w�S��݀�;d��՛���X��G�9ӻW����|�W'�U� 9�3X@;�UD���r�[u�v�ҩ��)^��:A
��
��Y���$+޸�Q=������y*MH�>�d��oN���u���U�ͬcm�CQUlM^��R+)ѫ���Ɠ.�W����h�q)	�t'H���d��Fp�_j�7�Vum�Sd
�G!�-0x�Η]l��u/(�6�6Y�X����m�e�덵ͩ9=�
��-"�ۡ��u�t&Nk==���<��,�]Mb�m��0�ډ�e��P�sq8sn��0h�JR�)��]Ԋ�V��,��m1e�f�w�w�c���yf�U�W��kH7�V��=b��烒���t��t�Yxr��B��<{rm�«��oJD&yU�	���d.���h'�36�5�,4O'F�n�1E���Mk��uu�X��:Y�'���j����$�鏸DګZTc��C�XE�Mc|H����$䉪y����l���Z0�T������Jc��׆»�fcɛ��.�!8XG݊i)T3��^���Ȏ�U3W£R���7i�n�T�f쬣�lUEU��भl<�i���x�̊��֣g&5o��v�-@�B�U�N4.����lJ�j@�.8k�1n1RiTJ�_���c�upF�mh�{y`RD_����v���>����3l���q^�1�M�r3G^U��igs���63M�zuvf�}��tX�r�*?Kj�P��m[[ݛh�
�<�V%&�"�nS���JKʮ�ڽW�d�*t�y(��Em�3_�v���C��L�P���5ݑ��ʏ�Խ���Q�[ïQͥ2V�X�c��*��!��CvΎ�;jh�B�9�KeCX572hV3:��xb�u�z)7�ͥ�蛭���MԮ�|ai�X�(�.����c��ی��9�q8W��Sz2���e&fZ�\s�ݽ��t�{]���q��g8�5�r	�S�G�k���Zi	 ƋJ���*�4�jVY��RTD��͸+oU�t����Ԣ����)�.�bo]H�u3@�� n�#ܶWM��H���3Zk�һw�g4p�[�1�V]��&U�ۼ!�=�fo��
:�_7s�1���Wk+_B��2X�s�����J��ځ��0��5�lhAodW�k��j�&��#�NW.�A-I 2��a���)Ǝ��9�F���Z�d�լ���ύu�a��Ȳ�"��͕�p�q]Z�Q��y|���iwv\�퐂�*�7��R�ء.V[Q��p���J��ʜ.>5�nH�_]އ@F��9�1~��R�Y�=�E�L���+�4�)-���]U[��ֽ3A���jYΑa�'��c�Ǌ�Ibv�(��dT��`�Ӂ�Ŝ"����|!��$]�Ŧ���/5'6�:������5z�F�y���u&d����F�]��m-�1M��2e��Xu���uZb�F�B��(�Bm��\�U��'�Rh��DS�jl,�!ޓ�����q�#Wr=[�j=ٮ�.���2�\�9�f�m���u�n��}���r�(ǫx��$=Ck��f�Wl9�{��rv�Kb�u푵.��œSd7���n�q�v�h��5N�N��b�.����aY�BDب����u��5�С:
)U����S{l��>�q,ɴh��։��nw%f� ��,cw�f�p���Z�E"�����Jظ�����$Q���K;B��ﮋ��,ؓ����3n���R��� f�b>8���Җv�`�߬ض(+��P&ۜ���Ҩ۝�8��0�5�U=�c�֑[:m���ؤ0�.�P�}j�h���:S�'9N�S���d��I��ˈ���ӌ˭��R�-ő3�Y��+�u�V�����R:�#���0F��Z������@��NJ����;����]��;ڗfGvzK<�b]e�X�v�_Lܲ��ୌ��-J=�rl��� �k���s���n��S�R������Dםy;��ͫ=+���Y�w+1��85/F0�0�Vj�a�����T��.փ��Stp�P�k�Š���:�vmӠ)	�ϴ4w�W��ݑ��}��x�[c��Qݎ\k�6Su\t!'��ݲ�4��mV7K����RL�+�V䢄�nV-�݇z�:����Y8V�=�n��,�f̣4<�)V�r\����+'8��R�����<Џ�L+��k��A������j!�,�z��e��O~heS�U,:�E����Z����u�"AZܙɻ�J<=oGEf�X����T/ea �sDi��l�m�SxS�[��$�tŵ��K�CFn���P0@jt�xp�Y�-�d��&��+�4׵Kx0�y��&���J���o溳��!r<^��R7�U�8����$r�����gJ2��%uFٵݲ������{���Jf"��8�ٹԖPmVV�FP��u}
�s:4Ma1��)rh�j�w�p��.�=w�:r��ɘ�a�"���w�륢t�"���H�;޼Ӗ+ ��U��-���q�5�ή��.9;��AL"��
Pt�Rm� ��[��3v�*Z^�PY����GEh.��q���k3[́��]	���"Ԇe�p�l��a�pdh�Z⒀�xjJ�(8�ѯ&�!k�d<5!�qsx�:��y3����jY,�[;aN�M^k,�����2I�p)����]0�T�����G���f���7���
��������1��ywS��9ܲ��Cµ֌�/���J��,N�8��F^���a�fXk*�)�WvoI2�3�ùٶ��a6=F��c���|R`�c�ݰ�����pz�W�%��W�Q�j��7�O	A����*ͻ�\A��X�#A�C
�.����\�����蕪�n�iu��ĕަ���#���jT��El�N��U�Q�_V� ��7�3I�Z�V(���tv�1�����)�dWJ0ѻ���eJ^V"��=d������.�ئ�8�U��.����w�j�\�^�Ç���y�c֫��1��A����r�%v�E��K����d�Y�wO1m�XJ�7��+�*���u���/�kU޼L>�ok��İ'U�����P��++���z�kS#K�#�<[w���H�/Y;��x��R�\��m[��4 ����z����K$d.Eƴ[.�pP�@�B��Ǘ��������>�����E{���u�����'��JS�����ok���Im���t��]kT���xZ=<T�;X�9��']�ۖu\Y);�S��g2�s�����i�֯L(�^q���ZV]0sT�5�;�]�+Y�ñ���5k���S����呑h�I�r�����v,Z�S�w*�,���g*�Ǥ6q��ݎc�	A�;4�Rq�B@�K�v��+���׷�֝�J\��fɽ��;�
ڱw)���;1�Kp��Ӈ���p.�m%�Y@`8�{�S���Υ]�tKikh
<�1pد%��$PX0��i�R�n\�˓+�w0�`뺏YM�ŗ����TG�e�.b���=ʘ�hQPC	�1��/��1��Ny;ʰh͌p�_���]�P5�V7���"��Â��1	Pm�/���'�����ҍ��ܶ�gXf�r&y/͉c�+wQ�n��o��u�l#r����^a��tEr�`��w5|j�Y����!�\v5u�w0j�e��pյ�f)��T���́[Y�j�<�J=���&5�a�"pc94I,^Ջ4��[u��,�N����]���;T�[��;���n��T^V3�&�g��p�S�]j;t\Lk��5H�I�o����]͊�wʫ�`���E:��<�{8+K	�8��=5� �F���e0\n�s���]n����·��촨P7�@4Z�<ʢңN� )�M�~m�q�fgs�z�-uZ��I�P^F@�R�BUw>��P�P�.��5Rj�H�L�� ��²B�(R���H��Te��)@deT�A��4��d	Z��(B��*����X d�Bd�fFFY��NUM&AAf4RY��!�+&�!�
)h2�����Z����\���)2�����ԘNF�QE)E����5�jhr2S ʊZ�PDS�w�
�?WUΆ��y�;�����%��΂������(v�9�Q�������scb�xp��f\�X��-xuԁ���^e�� p�}&�x�����qo���'�I��6�L�!:wV��+AYq�Hr�tdq����Dvޚ���A��&h��a�-;��mʏ�	�)��rF��r.�D{o�zE��O��v�k�8�<h�5�"�v�mTM��&��0ѷ��ǁ"�"�z8�n6�7`�m�I͙��~�N<�{�q��ew�L��gv��h	w� ��� y��b����j�\���UMAo$����x<����I;�PWClw���c�FzZck����FVf���u�3�Y/3�gbEsQ�K���T�e�.����;�&M��݄g�6�Y�O���$M�pq�n�<������=��P��&п����3.�*{|�/�6��O�{��d����4��6�Ӕ}'o}^�w
�yz��=�I��/�}Lz��0X^�p"��;���[��I���.�oو<�����]ye�=���j�bYU���ʴ׺�k���Z�2�5�P���˳�g���nX�����޲�B�����wsoon,V�n�r��{���O$Ev��sP�B��{ׇG$�fu�w��q@�P@�)��l�W��!��ᄴ���k�E?�{��S bV!�^#8��R�o��GtVz��EQ��{�{�YHW�����D;X|�l3�9�_@x5���j��-�R9�������O���� �%`��m���P��>�D(;׻�B8�WO)�s�M^y�-��#�����*��y���]D/�E}gy�"?�u���[������q�^��H�� �2=m"�����^�+g��E�t���{j�p&�h��Br7x� ȣ�fc�s�]��s���>�M�������1�R�~hS���7l�U�1�>�y����g�A&�Ϸs��=4� u�1��=��}Ck�B��%S�9�N�jw�'��`�;&I&���Z���8�LH���\�[�v�6���ڊ��R�9Fۿ��EM��y�<��!�Y��w�� �v��c+rb�I��U5�Co,i����o��tp�@�c/�k�����ЎgY�V��^���̛��Hz	�}Ng�\֗�8�r�^�V�.wt�!qأ�Rgi�-&�8h�xa�
�;d;�i�~JϽ�9�֗V�u,oWyb���=6�艪�E�r]�HO�~�z��#33ՀC�'y����<�oҲ����=�/rsnD\*�z�YB<��Z�>{_5��zd�^͞l�����/�'�ˬ����,ʶ�@S{c�7�p��nC����g��^�D��xQ)��a�,_P���q�}�?j{�>���~z<)5�z��y��eta�Tw���ޏ5��q�ё���zԃ��JThN����2I��C�����=�{��N�� �D�����P;�)K�=���Ӟkֽ#�
z�j~�"2�M�@�LJ�lw�$i3�}v�ԍ��u���߈;>x4_k'�6�<���<h���$�K��7W��!��|s��[W�2a��DLn[�D��jK�w�ۘf�����v<�I�f�<�5�^���j�p�{��}" �q��u�}���\��zWSnU��Ջy�}�۸�I<����,��\IZ8��p��L�����
��W�uj�(qK�`KAW��`7&x� �*J�ݫ�%��K*s��;��+͙���o[�1}RE[.�P��$��g;9G�c�7r~|�/�N^��4�{.~����?��v��!��-ӭ�C��6��6xL������t�^��\����٨[O�uh��i�[	{����o�q}:����Cb�=���I���c^'��j�}�ۧ;���u��s3�����e�$XC�/�����ϣ�6�t74d�=ݞyj�5Ҥ^�="�{z>��W��3a�Py��z�H�9X��oIޞ���S�F͍�N²7���<���g��sCz�
t�P�<�끽��׳g}��͚a���H�X��&{���ޒ?*��h��@�<��ޗ�=��9U��1K]�?%�ؖ��g˻�OM-���Y;�_>�k��>y��P�}�Ȼə!�w�����w���������;��=	����x���e:���:�u焟��X���hG�'��� �%��fw��,�
����y����#q��8�C���<o��M�a�c�Jo�g��ѕtm/#�^i<&d�k&��ee�'+�ɉպ�خ����I��9t�Yo8��Q�Fȵηl��G��N$-��:$oQ;vXi�Y̌�uݪS���cDfaJ����ج�#+*�E(��]�fatH=8�_��w�����Dd�r�&D��Oy?���#������3>���.�W�����yN�D~�?��s
�0}+��<�>����hs�9��D���Y>��=��76��h{Q&e��y��^�q�!��YFF�9��{�	vͫ���'eü�$��v�q�'ټv��|�}�}�/&�b�_j	/zKV�H�O;~��b�߾�C3֭�px���z��^��?F�R������^-���6�ǭ�u� ��$@��wH=^n�I�M�} ����;���DZH��\Z�Ԇ�������3�{�*=�qm���g����X0R.¦}^�=�:|�Wu�$~�ϯ�w���à+ݝb�+�wk��7y�&�2xa�I�}��f�A]��<Xc�����n
�b�ˇ�>&c�3)�S�+1��e�ܷr�,b�ю8���q��_}���݆T���ذ(͵�M�Gk�hˮ�Ґ�xM���6�5ŇG퀴��b�}e��vQ`t�Z4�!e!��x�ho�)bP�%n�t[AIn-�q�V���V��Iu;���;�_q�G����O�����%�|a����F�[�=N��Sd��yA�"O|���I��w	=3Ź�Խ��m2�S�u|'����6W}c�-�B;�>��5��k�NI탎OuM[���O9����gf���Ϩ[�s��	xp#���}sޜ=oI��|��+���6�����Ț�E�����L�FpZ<�$,��;�oӏH�e8�Lա� jK�l`>1����p9��$��N�;��V�(�]-����7����H����!��u�xL����ۧg��j�k����������-�"����f��}�N���K��o�<DOd1�5���qS����|A�F�=MY�{xvE�"��^���L�����o��K�%����4H�d�dF�u�A>��{]�x�r���Փ3�W�w���¾�W��^;�R�3VlX�5��`�d
}u �+_��L�� O���1]o@��U	\k'gny�~���&�>���[�:���׳fԀ�<�V����80�FLgu��R�,�}�/J��6]ˆ������	NM�M�5mw�'�o�q�#;ɂ�yA��k!WD��Lk������A�Ü�9�h��B�۹L`M3�&c��/Ƿ��2������A��.N-�I�$�I���ο��8ULV���y�}޾�)��̘����L�����x�����=��G'E�YYVz���i����׽1j;|*�U������2=��k�ţ��H�gK��t�/��򄆻��ܾI���n��S��P�.���zv�Ӵ�����7�/���~cd[�}ž��zU�|��<��o�7�X�1��M٢�<��;�SWw��R�5I��v��]UW�N������9���t\p����v�<�~p�Mpwr]'���K^=#�t?f���S��|upzD�w����d��Թ�f���u���S�ޓ�\ݐE�Lz#k�V}�/o��Hs&SWD�}���й��F��Qc���.wj7ט��>^'���"�����w�~TsBڻ�Z*�z���6��*�M�
ٲ��1>o'˞�uT���v�I��3ov��Ð�]-��N�ޡ��c��ũ<�$��0s!�|EV�p�!-${û�>���È�_I�l�`J��C�m�+J�h�H,E��M��a���'���_2�z��'���Z@�˝^�gw�r@�N���t��h:��ڿ��g��Q>������iɃ�e�����'������6��ҏ�Dk�&Հz�z��Y;�3��B���G���צ��1F��A<(��=m=�r.i��E덈�`��ݒ�͞�(xy>��ӝ�}�8<�쇬���fA۹يa��lk�9,��W'kz2S��[C�0|��~���Og����P�������x:�4foyN����|φH8�˩�N��珞n<F��&�"g,��0h��ɋ�M<-�m��؂���ѐ6oǜ�gg��<��U!���(�6����y�-!������p7��z͕���3��7�h��c�w��-^�����n��}�����_�H����AnÝ}�Y�7࡞8zs�B'�q��e,}���������!����-��|��'5 ����U�#��J�H1��{�aS�崬��΂jMW|zV趂ʐ�8e���/6�E���o�TZ��<�G���{�i�,�.<�~ay��=6(]t��x�''J�/�_���=8_��= -������}_A�':��X�Ʊ[7s��bj��;
�#d��s��'�Ŷ>�>�z�5wԸ2)�Ù>I�ٵ�O9�9��D���Be
6o�<��MF���[��A����na��Ԯ�u�ƣ��۸Ί~*��xR�p{ލ��Df�&A�)׼���e�/z������N���k���	�e玁k��ln���������/!==���Op�H���`��/ׁ�c��vH��K)׾�e��꘡��O����=��]�{~/j�;�J�y��}�KΝF5�J����ۧg|w:Fv��hԚ'��f�TK�Di����sj�~����A���0}�ŏ|���w>��j�����s1�\�Nda�UK��� �W;�p'{dj6DY�:ϫ_��T챖�Nj���B��u�)O�b������B�SaWV���C���MtK��"�Ĭ+D�j��g�{��Y����]��YK��J���&L̾'h�%k�TkS&k��w�Ī��Kq{��7��E�]�m��;����p����h�Jy�T�q������BF���_�$\���/o�f};�x��-yWe���ݧ�`��&A$�m���sc2b[�١�:U^e�tO��Zԭ���Ճ�I���l9�{���4� ���Cc��}��ۆ�<�8{<r����ڋ0Q����(=$^�7�5KW���pW���1o��9��c�����u��M3L��I�-9����c;=G�����a��`��3XK�a��`]�f�dᡳ�i���oA=�0�NdTV>9�cR5c)�i�5�{�>yT��9�,ی���4���٣qN�x>��fD�߅�7�طd��&��<E{Ä�a̼Fw�G��/�yV��*�s������WC��^���ވ��iA�ś<�u�h|�<�<�'ӷ���|v;v��w�����������L�F��Ǵ7/��u�����2�z.T�j��j�����]uY��,]-��\ڼ�(��{�z�۸9[T�f$#)[�SS���q�Km�C_fe�G��җO�rޢq��Pغ���ʂ������4W�Nl�hދ���f�G���
���z*Li���E�2�X�쬂�[�h���z���Oj��·`�柦#|Ň�u\w:].f�p�CsK�E�K$�k}Wx�}0,�ڌ�aR���k�{C�g'M�)�o-N-1��j�Y��{<'N#%�Y��m;�C$V�K2���Jh��uu�e`�箤�:��-B�a|�F˵4�yW�d4���u� 'Tq�ʵ��P�,����^nG�,Y}l�Y:�w-�8AW��*w������l��o�{(�)������āT+��<鉸w���jn�Z�d�]H^ȕ5]}]��9��YB�6���H%ӕk`��7���j�r����;�E=�K��[� .dL���՝�p��h\CK�̾�w"WA����Y}jt�fVΕ�\;���L�]� �s5w*q��KKA�<̾yP7՗�(uQو���E+aZ�A����ơݱq��I�w��9��KW$�o���9V�up�-��7uJOh=�݃%�ҕKg��H3�Q��Kƭ3��˫��=�#��2*걥G���D�]���yN��J������_�;u�bn�ĵ3׸dW�8eC�.M�X�m��K��4�[B����P1[�m�n?�1�iX�Uf��tַP��=���%..��-BZ��Fc���/��,N����p���Ӯy������$P��٘�>;���֣��Z#����|b.d��o�d�1<�]~6�[�C�R�C.ҽ�\j���M)�^�L[s4�7B��òًbSD��c�gj�-�A���t8�:�t���;ti���A�.{�xo"�F���ho�;ֳ)� nT��s�W����L=t`f�Ύm-ѕ����Ӽ���	G���p�˒��u��V�2��V�}�oM��I9�ގjǼ��Ӹ-�zf�V7:]D��˻��+u�Ʒ 8���o��#7�!�Oq=�r�$��j��)l�'�tжwAʧn-k����8w5UR*��跸��+d�6�(�"7sUP\�k��ˢ3&=��=3��b1��+n��k5���xE`jd\���9]������G�����d;���AV�u6s�#4C��垾8Ӷ[x(�[h�w�Y�;��d㮆��8M��R�r�4��H�0�W+��.<{�/l�%3J��;+����*͐�^1G�!�S`!jm�.���)�}�!���c)⼫��]�_--[�:5�P�!���P��k��y�3Ew��ⷃ�r�^J�v[���9��]�m�\��1&o]�Re	����iIiˋ7w9�p��<���|��fk=�[S��|��JiV��ɠ�(2*)��A�F�*�i2�&�&���5+��
rF��2,�X!��rL,���#����N�uQ��a@VM�BDP�R�D��CUR�4�&@QN�tZ����!ɣ,��r �Q�KX�cFAH�aE)Z�p�Չ�É�jZ��3Xq:�g1Ď�11*[,�̣�uZ$�ʉ2J£$���"��L���bDa�f]��-$�	��1L�U�e�fffd�5h,�,̬����1�ba&�%�!�-a��fa�����j�20��(׉�~^^΢��}��շg,���7jxj[K`A�YL/S�.v��X��)�os���K+
-��� �G�_y��)O�_�w��_�Q��&[����0v�;���H�G$/g�hy�=J"�{���3��+��;˪��m,��Ƒm��:����O�q������,t��K�{ؤ�c�뾅�ZZVn��ޭ����s�<`X}\�Y�&�-������n��߿@7 ʔS���s�L�]>Xy��x���_`q��4u�,�E��f�!M�K�'b�>;����~�j������O&�-�w���\|�ˢK߾�k^��ޭ�^����@�.��Ly�V�8��S/�D�]M$�15��I��嬼�89D�/a#4�ĥI��;��F4'�p1�$>Q<���N�[?c?^J�Ӽҵ�CB�� nI�nx.��bS��S �%I���9�y�.W��3V��y������l�=�f�}���1o����0���a�ِ��z�$�^S��M�-.����c��)n�OTJ��ѽ���U���@�D@�`��6&(6�G4��*]��&�z�1i�g�H%���l���iq�Z#N`+f���o}��~���_��{��.�q"����n�ګ��M��@����O�ݴ�z��z��Z���kq�҄G	9�$(0s�m�Y���7J
�Ջ3	Q��5�8^wVZ���v�s+\���Y�uvMn.�N�C�r�鏷pN�,�2���f˦r\ŦY7H!�T�3�hds�:��4,���J|�6�o5�u�K�]{�o	�z�9�_�θ�g�I#�U*W��\����})������7�n��ť��c�M�_N�5����a��Z���y�s��fƖy 0�?�yݛ\����uٖ�����u���Λ_+�Eje0�Ϭ���=:��p�u��:$wUr�\��u��y��a��ݽ�?X��^�=���'��p6�U�;_'ә��a��`$�Q��_�9j/a���i�J�ULA�v��ռ;>*Y��B-��9`.&>�W�#[�}��@;��P&h�Q2�Z}�����W-+e�&�ꉷ�����*���x����*^�!�nG4��_9�=8�nu��]Ѧh�.���Uf�qmuY�pᆟ���>��� ��?5���x4=�)�0?�ol��U�>��y����T5�y���b{_�<�����1j���3���8ʆ@�t��N�`��$��������e�((���{�����.��Ư����xa��/K���c= u�5eEÚ������[{����EZ�5cWI�߀�|Nz���M�jl�cPɏ����2ײb����*��zlרs>>����XW�|�m'��U�J/��Ӳ�7/o�R�ȳl[��@+$�R� ��.�zKT�1Uڭ�f��J��.k��˭����]�v-����k����u%���y7Nk�}H&(�*�l)4`��z6C�q�kSǹ�F��x)���3i9S��V�:�mBƿ;�q�H>�;�k��X��3�r�@k��훒��Gd���	�p,9��(XT/nU$���!����S���t�f9�
�[F׺q�B�>�(8�C)�n8�n�P�Ԩ� c1O�魧�P��˄�Z{md<�c���.4��/A�-�n���i�>�^�7����K(�4�
�M3���Fg�!�/H%6ĺ��1�F�pFh�~�4lU/���-�x��/����7,'m��ܥ��P��RaTJ�X�BO\�Ƈ-�a 'x��7!����l�����X$���wy���ٳzAl�WQ\�����s'\]��E��<Ư��[�K֮݇�E�y� Χ&��j�k������	ۓ���G1����gR��Zx�o�s�K})>6uAa�B5�P]�"7!���2�˃!�xF#��4tsH��\�Ԁ̷�Kc��䟦��ӯ�t���.�/a�S�m�,l��5Cs/^��~j� 2%�<8?���y�6߬eK2N�wK7Iܢ��a�֓Nd]�c��ogu�#.ݯ@��iD[�s�g/��0'C�whOl*-��G�ӅO��z�)^��
�������1�cn�ָܳW�^�f���'X[�Q��<b���e��7�p�����$��
P�o���l��_S�ێ�p>��vp;哞U7�B���E��H��n<b;����{�"�¶��.��׸vn��n���旧��u�U����cL�|���r3"����c�ӕ r�T��W���.��l;G�5���ɻ��\�]���,��5,������^�U�B�F��q�����go2��:��&ن֪m�޼�� �渑sM�k˷�J�Zڽ�H\�@tR�p������xe]ڕъ�U�eFoN.��z�'�Ô�
g�8Bli�0�}#���g+��nj~"Se�!2�-��bm���J�/���7r-�����E=��	��鄐���	��֠f�!77���9�5p�m���n^+s�q�a,`��n��з�x"<-� �{ɀBy�c@!�8�0ӛ6!y3s����O8n���{j�:�ؙt�Kvzm���S�_8k����A�l��.p;l3�p�8�՗��*y�@lCKH�}%�}�]0�jQu�n�`�˷�~b�^��p&����Ӗ�v�53��,��ѢuL��dIӴ��*�*�s�I��~nCT�~jN%À�2=����y̼]�{׬C�?�c�h-0�kv�Ip��`[	���F]c�9���s���~W�w��ʇ7���~�իPFɼT�j7�&g�_m`�1�x1*)���5&5����m����yn�5+�2]�&v��ִͷt���Hn��z��.��p����L|O]�k��]�����spqޑtok�͗����K�Ô�F/,���.D2ק`8�p�o,:<�������j���Ҝ`��J�)c(��S�жpŻ{�Y'�]�/�������0]��GH`�8t�#�ȇmtӓۏ[�6ɽ����v�:������P���6XF}:�L��{%���Phc�0�����LW>��-�t�sX�ke�qb�rHf��%�'�I���v�J+���;�vv2b]�L hͫ���\�R޻n�c�
�.NJ/aTf�&������	���"�Ӵ��o����{jVv�3��k�n�o^fqw���sK ���7'�uE���wP֟n���4ׯ��%T�7ܤ�����&]a���8v��l-��avPzX*��}_/��Yͯ.9�3m�)f��M�~���՜�x��y����P5�9���R�o^~SG]�@��Eޟ�åV4�P�P�fe=��h�-Y���[k���j�  ŪњOr��
=�^��x/B�� �d�e�	�1̐p�z��U���^�oRt��A8�Ƚ���+�&���\�ΞE=�ă���\��M*�K�@fف)F:R��]H�W��݊�I������.�v.��=kU[1pҩ����*R��_q�j���̷X��f���>4�rK���<�*1�T�.�k���Eº8��f!�]�C��\�HR�7��AR�>"�g5,>u�d����#E�����d����&�jBa0R��p��\�69��u/�9�N��)�y%I����<������.ѹsT����a^#!�ZE�4�lLXc=����K��);��F����o`Ke1��;��ɖZ�~3]��f�SN����{a��9�O�QA�F��Q{¥�A�M���`OI�6�T�M���}�7e���y�B��Z��&i������X(�g`�s���u��D��j�kob��g<�5��Y�s��^&G6��-�@2�q�����ga !�;�������xW:ot�[�%D��l}�-���3,P�5�w�ғ����L�z�s�5R͔6-ݛu�5�����mU�h0ʯ�j5b9��V����T7sG����L:�ƲǰA��q��b�aǸ��#��}�MN����bѦ.�g����6'�w���4��$��H�v�LW5 _�9`3;;uU;9-8�V.sJC�@��^$Y�8M10���j|5���A���B(���L3񚤞�p%�o�oe"���!�_zo#��g��^]���i���\��m���>�fY�h�?�� �UU^�X���ۼ-��A:�wqn*�w�U�k�2�R��F|yj�:shEQk��x��p�6�T��':��a�.�b��i`Yx�ua,��Gc���qn��ΝN�wuH�+T�Y�C~S*ܗ3v�I�j�r�����l��������u~�ߡ���*J�v���CPH˵���h1X��"�[_�\+��Hڱ��t忑$Y�=�_�O,��X�M7����\­B�Oid�j	�z�l�*�Ο�]�a�p5V�����ͽ��w]�oX/L�62������݆OB�	eE�z:�����\x3�Stj�
�;Bm��}�ͻ��.2�T�k]�3lZ�as�~�k�1I���J� ����`6}x��佛{��=������|g^��
�]L$�#r]�Od����2O~bS�Hд�ٛ�a6����#w{��e�)�F�0�;"�{���H"1���?��Ð�}�.�E�K矺����:|2�;&Եξa�T�Z�7j�)�\I�lA�/N�e�0�qh!�!�O�0�; K&�υ�`�é���E�#v=�I�I�қd]c�^/B4���Msם���\=� �k�9���:�[Y]�o	��y��!�3����*�ki0�����.Rz�%%�[N�Bxwf��������%A�	�2Uݫ�FU͊ k"�/)΃YB���q{�Uk
Y��iT�������{p����=�yV�i��m?����Z5:��P�D�ٻ�+�V�(y52�.�F��L�5�W�j�1p��,~�^���y2����`'���1���Enٰ�)�V�-XH����6��[�K���P[[}��s,l�LI����II@OEU?�ϛ���K�6x�����X��
9�tm�2)!�S�o'qɺ:O���yTp������ݽձQ!N����zC��fpF�0=���2��Ø�R		�k\x@ƚ�:�+g��k�ƥ��w@��`Pg8g��2�h����߲a�'DwL;�{n���q���m4w\ݨ=�;�[�1<���91݁��g/:��@������!�8�9(�0�-�s4۝����Kw*)ŻǴ@<�� ��F]�l��&�׶3�0%�|0V���h]R�����yd�y��zl��>̄C�_8*���k�"�m�t=C��A;n��;�s���5�7�W8]��<C�q>����X��j�ʩkmJײ�1V��W�y*:���_6fF(�ƛ�����=u�0��*ytS>��7���C��i�N+Y,��b��	��`&M��:����Q��uD7ivݛC�פ�P����p+��o"���-�'C�	�����#�O0���ӂ�oS�!7·�-��ŵ2N$�MjR�o�V�ϸ���$8��HP�z��Bz�x�v��6*amkb��˶��F/����5�+���iz��g�T�c�uk�˳ܩ|���(���F�ig���/�}P������r6���woR�7&W)�1�\�,r͐�v���Gf����[}Zy����K/�K�vXj�<]*N��̶�=��S�q�!R47��aS�c�:��ʒT�P~���s	��ր]����"�吻R��Y��z�z���2�q�I�}I�{"���J.���PZj���,�\�5!�+2��ܺr2�)dE�1i�!1��[���dQ��������`r-?5�$�X��P��m��1}Xb�/��l��A��s�S�`嵤��@mM'V�Ɩ-�슲UzY~�6�@��[A�1u��3^�#{2<9���En*4�R�\�_������-Lo�Z�XR�[�V.k�|V��++�sM;�N�Tq{��+�i7rʹE�~�4P�%���C,
w���TՁ0e^x��T�SC5DM��7Y��#&V�:�	�F>���j=��K�A�� `3p.tB.�V���)`�S��M�7UZr��r�P��}}$�Yx���nzb� �b�:�;�p/k0��t1����ʈ����f@���A�HBj|�)�^�a&�@;����	^������ܵ��1Ƿ���:����P~�+H��u0��D��}hj2H��I�/�{��������7����B����G�$p�Ϫnc+&�c�(g-ѵit	�����h��ъ��W�޵Y���8쭝�5�i�5o�r^�@��ɴ��öd���}���������:zI4Ⱥ"���k��G0�
����ȹ�h��x�=���?�U
���*���/fVQ<Segf�w�\�z�o>זxk`К	!Bi�de9����׷&m�%,0zn"ю��������ǟo��w���E,���8|���.�H�x���ρ�|���I*�������8jf�Y�vk#BUOq�������SZ�MV��{��
=�V�o���A@����cZ��d����w�U�����~�ţ��E�0�q^&%�{H��ĥI��"�],����W`{{�Y���v��jk�UN�C�
%;6C�9�cO�;$�ן�S���%:�H�I)MM�;'�ņ?;6�� ���;|�Sh����3c<�3n�pe��p��K���4��yNRn�
O�U�9����Nf&�3qjX[�����=0 ��9�jc�l�O5�*]�������S�T��m�S5��L�W*��^c!��<����	=�|)o��Ҽ+��Ѻ�N��C�����=��tAe��(n��V�ny�x܌c/\c��3��b]�F3��y��?sȇd�_ݡ=�S�w]9W|ٗ�_q���@B�ƻ��I��-2m����;�+�'z�2���Qc�<�zg���O�������zyyyxv��ٿ5���2,�oGs���g�Ɨ�(�R�Z�teڹ���hÃ�����t��[)�s��v+�4J�:q���M�M���x�&^�c��}�؁U���gFw#�oa�]#���R'Aqf� ��j`���Y[3o�P�:�?�D,�o�����V�Н�8�4�1\��g]��+��4+��n�`�����(��5Րh������[:nf+�Ur[��0C{���ˏƐ�p���XBy�j���;�o�i�HU)��V,j�_y��̊������6b�Eb�ж2�Θau�PX4n�wΔ�t�׀��me��:�p�]�2q�Cn��EU�z���ӡf�N=ɲ�T��}Μ�&f����:�B��]y�4�����F-R=���Z��������m�����;4�2ʅX�n�4����j����%����|m,���g3:p��iK��23���M�o�y�U�{��hD��xa4��Ǜ��F�N�d����ok�j�u�9=(�BoM���A>�8Z��^ĮU�P䪏Z�&����V���Ͷ��a�<�]5qf_N��J���^k3ϰG]���_
W��w'*�3dޢE�K��K5yW��$߅�bă2�8d�j�$f����S%
�����u�� ����(`�g[γoQt��e�ɢxQV+����Zk{��S��I޼U0�yx���ú��˄�k"�J2r��z�R�����[��K^@r��ܛfr@������m�ʶ��-�G��N'��U�
�e��|<�[�Պn���fV���T��ʑ10��=�om�ۏ�)a�@���c��K�����93�~������k��i9��1�����B@�c�ǝ���ݥU�-�<f�ܧ���_bZ\�U�{}Gi:2A%�ԑ��Q]Y�������I�a�̡82���JJ���TP��߻����u��d"rk������7�fl+%j˾x��#n���y��$�Q���3�73oȻ]Da.�+2�#T���-ҽ}#i��\�t;������>�l�`H22��s��.�%�������s��賥�u�E�|(��)q����Ns\J`�9Ʌ)
(\����f�b��P���GK���_�	��#�i��W7�.Z�톛�c�6v����Vwz����k;��n�`,dc�8����7��]��1&�i�mB�Ġ�xM�*#NX��*��Jj�����Vv���6�f�yn�3u��MM���X_m=�[�g-�*Q���Xu��E�9ڇ*	�D��k䑴��&o��IR}]�O6�,43��l�a�T�����{j��j���ݻ�ʗukm�ܼp����S��Oj�������G�Z�s�R,��e�5\�s:��X����b�g7a�R݁�|`�[H����T�::.�y�:��E��f�֥��=T��vSj��k�h�YCrȔ�G�X���t��6µn|mm���SM�1l�8ָ-54���Λ�΋����̀"
��# h��O"L�8à�C�Q�����n�-X`���b� P���f�&	c2 �!˫"�,0�5a�LI���LT�`f�faR�eXYVdc�Q�j�5Q�fف�kC���k21�0�Ec��ZѪ��e��R�hkD�%X�FFNIf�N�'�S"�
�Ƶ�D�Y�Q�$dfa����#Pde�kT�&�����M��hŬ��,��
�j���mRS�N�%�!r���(���!�XdZ�J*s2����(�(��� 0�h���i��5kFU:�+	�"$�b�T�QY�R��2ը����2l0)��0������fUUa��L��U�¦&c �M�����ȴj���!�ohb�����D�@��Z����X4�������%)aˣ���K�k�\�'$�ĚYe[�wY����T�� &D�}���+�T<��3R]3u>�r����zꆿ(�ƅ�}����/�,rz=;Ƣ��u��Hwno9��s�ѹ��i��p��8E����y�K�bz�z�]�ͷ�h9�5�$��Nf�vi1\�Jҙ㗾f���G�z{.U	~d5�;�l���\!0��K�scjF�]����4"�L�voqǛv�V�i4��H��L���n���5��y��["]� �E�5��I��N6ۜ�<�s���H>��X7���N�&hZes�%6� ��˴��Z��<����N���F0��ȸo}����f���d_k���T�
ֱ� H8�t7��H2F1���P��^G=;Ǭ�s�m(+b�kgLrm6M�p[Ρ�=7�E�ŹQVϩ� �[��A=}YQF���ɿTB8��_Z�鞧Dys�W�b?�k{���ȅ ��q���m1���as�~�~gZ�LR}��Хr�0�\�Jo%���I܆'Z)m�����9��*tu�����O5��ی�����p��	�{s�0�}����������`��QӒ����'��F4� �a�e;r���z�������:�W�����_���2�i����dt�{9JPV��£���:-��/�.y��.y���V���^k�1	��3m˒w۝qTC7 ��K˪gN��.��u���q�t=�Յ�\�Hn�K��X澹xLԤ���,�P�I��������%S;羽��7��~�w�6��y�n$&+T����D�7�8^���N�!�9	��9c���H��Wļ����)b�i9R�Ղf�Y�09��K��=5�^w�~y󇶄-p�˱|��9�g�^�ޢ���	y.��:�aTJ疯x��OW䤱��5<;�F�>82�U;I;WQ9�uh�t�`N�r��2"n�(���s`�P�nd닰	u~��V���������}`��P�;e���sPe�����hbڃ,ZD	�*4u�T/�ԭq֟�k�PK���β������E�_�܈�W{�ø
|:��3���i��f[���jR�[�qXV�vF?`�͗��Tv���1�Fj�u��h���<���_90!�
��D&��~�2��'M�qI�Hx�D��pD�jf(ZT�W(K��]��f]�p�ld{�[9y�]�dh�.>�Lu��o}Y1Zy��br����n���{2-����h=x�4�2�'D[ �tM�o����VGSS-51}�r���HAv�	����*�5�v1�fC�D�� �x���W~�x;[g��yxx�u�5����j��C�轨��Ŋ�D�#ܖ�G�a#��Ĥ����w3~4�Ҳ�l�\ʣ!���ܥ���1\�e��gK<2łEP<��n{�Ǹ��E�2s��U��Y��)GjV�x�J3�v�ڠ#����/r��Y�K
�T���k�̑��=�� ��[p�b�K��L}�,��KsƟ��|i��s�r,leT����M�kaV�D���nmc���͊Y۪�áy8�nb����3�r��0Lv��1N2W;R�s7��_'�;�_����n����)C�[��}�Y�՘L�B��X}G�����̩<c>Oa����y��y�G4�x1�.l�R�3�J�؍�ǭ}Ǆ�o��!Ŵ'H>7�=��l�'�;�]��l����`���:�hF�Ot�N��K$�<�ʒT�S�_8�=��z��d���\�44N-��3W�93syC����������E�xX�\]"�X�6W����0i� Bc��#@g���{ӽ�C�GCg��yn�0p�hQ����P8����O�a(,[й�_9�yښ):S�̈́�NM)� �0�����x0r��#[��SEՍ7Z����>k�ATe����$&(�^e�G��[��ks,)z9�KӇ��}>s�lc���	��L��M�g�}4ͭU|u�C_Or��^��W<����{����`v�
1�:ur����R#O�~>V��~�+Wt�/�i����Q3��hnUV�l3�2�_d6�3z��tv2�s=�oV�����߯[;�E��\��ű
�Ѳ���f��&/�uض�yc$�PQ��ⷵ6�P�\�:ư�-�۱3�,S!�Ŏ	˝�t�I��<���\z�h��^y����� �*�*=s߽�{׼���~n��|����%I������>�rb9��f4g�<1��`�v���6�>l������!��α�mC'���ͳ}(�X��C�"m7�H:"���Ž��<�GK�K]h�ʹ�ռ;�R�{��ĈJ{/cj3]"d1̛`�{����- �M;!�&��cw=U�c��X�?���j�᝽�C�KJ��'s�av}�כS����P�}��EAN|�5s�{���$XZg��Ƚ���)�����������1b�~myq�J
�&VK�fm!=�eB���#{�6��PcMi���ZGh=����O ��[Xd]��֭���u��wv���M0:�EN�%62b-��(�0�ј�בx�OB��N|�ޙ-�Υ�8����m�R�C��½�����N4Ƚ�f�X��5ߢ;��t�(��W)>Ȼ]�׭ɲ��ߐ)&%;6ÖnA;d���Jt�<ħVH�TJ�lW�j�L�6s0:����3]�򥗝E���83[L,ϭ���;%�)���'��i'b�����V���e�x0��_�Ś]Z�{b�Q��gd�DR5�f(2�.#�y�S��ٻh�D)��Ȯ����2A�_��$���X'�Ѥ�{��և>�UUn�yk L��y-��K�"���׼��ɞ�\���r�cWb�o�����v/���'U J�f�c�k8�qq�*���P��4�"!:�7�=��׬���7�U�R1��>G�d0�aA� �Bm��`��`.��v�o���R5p��k��Xˤ�ˁ�(����bXa�ӎ���8Q� C�_��\�;��VK��c�Y�i��m+c�gZ�[(����^�4�� K�o��X�������`�x&�%���ww;S���}�n3X'/�"y�{�}B�ߠ�cY�I����*c����f�����=(P=F�Vkr����.\x��vV�!�?��ϵ�k�ՇR�u�e�`��WY��j/�{�����4�����5��s�e��<p�ŝ����;�{L��i' �%��D��E����~�`q�]����;�k�[�����3��"9��\����;05�ݐ�����l��$.�7�j{;��r�ni&���e����.�0v���}	:�ON6ۖ��A�V�>��%T�����53�٫�e�����.�Sl�W�v�[�Z~h���%��q�cx+�Ʊ�uN�5�BӍn�Z�5��݊֡�,�����A��E���l� [:y��5ßo�ڨ᝶]O;�B<��B6⦵]O��0����B�5��_g��yi��:�6*#��Dv�u5��뛕fs��H��1��"�kP��M����`Ŋɓi`�n�sG6�^��jҺ��s�c���׸}H]����v܂L�Ĭu��h�2����<ֻ�;�9��Ϟ���%
�B�J!JBA - ���(-*�(�=�I��y�(�78|�����f3r
�eE[jr�w��	�8�[�ű��[��I�=h�k^��<s��'�Þe:����)�P��v�{L�&�2as�� �-{&):��Ф�́QӴ�(ֳL歵�ssw�,�rs<�=�k!�׈�L'�*T�UL$�4��.�$�����	�p"̬ʁ�ω7^򹈬Y��hY�*�qw8�Gd[B�:q��H F4�t��;�j�0����x�{/*�+3+�==�'e�T�1�t�Bb�1�V�D�7p�6S����@��'����TҥI��w���1�؄u����N�eIOVL�"��敥�m�\��z����W�]Y9�C��� �1��L�x8h`�	ok!��z���t�&@�yj.RzJ�%��������Ȯ��K
��S�z���x�o��;��_�TW/C�K��� �E�ygO1�WZ�s�Y�n����Kw��������T��*���(���O�(LhOH���4-[�Z�?J�:Z��'OU�����vx��5��-��\�Xw��0��gt�@}N��R�w��+��^>�U׋�J����/�О���Ѵ��l`EսYnU������B匱�n�v�3j��N�^r��
b�>�ז��R�tt޲�LnE�A<� ��H���OD]��!�]|r޸zѐ�e^3ϐ�Sc��Ln91��p%CET֒��nYa����}��Ԁ$�!"D
Ҁ�SJ�J!�$H+H�> y����oUq��]C_Wv~�SZ��3N׉�nj�az�3�2%�ހѢw�~ot�oF�袶	���LǟQR�d%�i�����c��̻H:"��g/�^]� `Ky�+��5�Q��������y	��LTkwp�`�u�4㇜= �z@A���c������-��)��,��r�o3�bˇ@�U!)8�F��=�E��^�cf9!᫜�r
�r25��p�z�������Nvw
Y/��@��TS<{&,:O,�w4^e�eT���k�B<�9��gT�ɐ��,����e�8��[ӌ.aּ��魻�i�9�F)�J��*`�P�c'��Su[�\���p���jd��+�4)=�8�Ӻ�1��E=�� b�S�!�7̐l�O��3���Րx��{�^!�:�Z�'Sc��JKԥ*������¿NS�V*��>,a73�f�M׹���&�`�k8#A�^��%:��%�u��)��&&t�8�̘NN]ˑX��^j���0��m���%�n�h�����EL-�F��T�����=Z�(��lY����!�6k���_/�L��U���v�b�s�~�B�	O��q�_o�/5G3]��D}�vk75���Q�z���&L��b��Pڡ���&sSE�{Z��U��'�PV}�6Ir�}�=z�W=k�]|(?B�H�� �$H�D���P�( 4�%�0��� ӵY���]�b�[��]�Ty�h0͌�prٓ7vNJ�֧e�9���|P�Ԫ+ɤ��vm,h��-�T�9j�q.l�?��M�1�5����u`����-��R[Y����C�	�'9r_y����K sH/N��k����6%�?�ˡQ|n��q֎w�S���2Mk
�=+��PK�=��cu��L�t����<Dqp���N�1s�gw;;z��s� .a�S��Sl�
����S��N�1O�mW��E]{}���<�NC�E ��]�W愄e<䰊/��]���d3l�J.X/���x�zA�ŀx)����fS^k7xe�@.؁�w�X@!�8�f���f�X	��[v���s��8����N|U:-�ٛ�w�s3V6^��v� ς���0�����҆Ai��I���{=��ln�i�����j�*���b�-sC���@�.���m=sͼ4�ש�}b9��N���_�UO��
�:B1��q�o]]���KU�*d5.�m�R�*�6�5�Pz͜OX�o
�H�x����E����o�*V{�5��Y��l����̓D����Y\�{�.�]�m�lq`�ٚ�9]�3(�0r��wV�$>�X�:9�{u��%��{*��@�u;���7G:	�B�_��q��v�s˳b�f����}4�������N���Yz�^�=�ͻ�2ERY���y�\ae���Yƾ�e��R!
 U�P�Ti�F�Jh���B�)��V���J
UX��@"V�ߦ���燞�~uz��:ۜߚMK�ǟ}��&��	�5gD���}ꀽ1���o�|w���z);��b�<�Kn��)!��� v��;2�*��?B	�$�M3����(JSWDr�ƵTe۪���9�uUmɆzt_�H�>1<��S��ƐD��<��S���%:��)�l`j�ļ�P�5��k�*� �@F��P|��4G�@0�m"�m��,�d�"�K��wQ��N����M#/�T�u�h�UϺg���a�D���}�l#�!��Bm���x7v�4��l姝��7VZô�͝�]��	��y(�����^�'��5#4�����c,sH�9Ƙ�����N�e�:�&%���Z�[(�������Gs�,g Ļ�>3��69�M]M,����9/uAv:�mu ���Rsf�SMc]�Җz9�.3v�j��awL�c�ٹ�C���[gSdvy8n���;G�q{����i�j�Ja�Ʋǿz}]`�澷��ܰ�g�;���(̇�B��a�8���Ŧ[ƻ���4��$��s4��N��v��Z��^�?[��μ�7g 7pR�Vc�6����j�M�ܛH���y4!AT�2��0��y]���w�_xa�PU2����ء��GIV�q�V�v���:	I�'��7�קy��y�q���=���
��j�V��a�Uf;Y׬�*�( ��B A�h �Z ZP�	`�
Q	��)A(h�<��xoz#i�J��A��j������ �O�'�v�
<:��ڑ��8T�rTVǈ�=P���X��渿Xf�}h�qNɩt'q!p�O^�o
��%�q�ߙ��Iы=���4\��gW��wn��*b_�S�2�3E�]��M�^��O���=y���%���4�]��4OCve+|[�}�0N���ߦ�}]{�Z�1BAŗA�pJ��$g/����lgOYa���t�mI��H��R��$B�v�yar%��F�����O�� ��j��-�Ƃ&�6��p�\�+4�]�ڨ{d�\9���à\��Jq�1<�#T�&�d���A����X�J���i�f�*�t�k��q��%��''�Eê�D�s�s	;N�p��M;�k:��+�
ukn�k�Z�t���~Hе~�I8���Ы��$�!�&�Y5�۷ߚ~��L�?; ƌ;|
�I�1����E'��4�3���-ᄁ�<��2C2+�3W
ޭ$K��@�5��N��RSՏ6Ⱥ�1��+K����z�w�~~�O�>��o��oO���>>><�zyy�����y.�1��ך�#���2�v\�[�s�t��KR��"�i9nc���z�m�pG��ҷ.�Vt��z�f����*�sp�2�����B��&�w�����.�Xs��Z`��M�]ϭ�g^a�Բ�ۦu�Yy��oP�(v�Q�靦7+tIVTN'�u��h^��\��mCy��,p������k�p��O�]��a�G�c:�^@R��%��G���VE�T��8P�#G]�QU��(��S�^�8��,�e���!�4��V�aW��sˉ��MN|]�K���fl٭pl�4�a������h��%]��^�/G��Xfq���{c�ʻz�I��ә�͈/����8*����	Nr��주�i��
�4��IS
�N��$�ƌ`��Ro���W�fC�E^���ꪉ1X����UKf�2�C�5��"7*���!�.�m@�֡c0ث�k�9vC�Wjč���
�ܷX�����5�V�)p,�}�[�1�vGeM�-[z'X+C�y;燷��@̉<�L�{��%�X�a*��Y�4#[�R5ndTUI�z��A��6�f�1J�{�'�K��zK�8�V0zҡ
�:��8�݊��a���z���i��:�Aa�5g=9��b���K+Z�A��	N������Z�8W�k���ӎ�oM���6��
b�FVZ[�4��Nv��JL�}D�ʺ����':zٙ��a��!Z��C}Io�@���`_��sO�)l���.����w�3�{�A�e�p��|1��^+�{e"+��Pb��[�Q^;�����G`��7[}c��%S���95�Dw;��,�2�/2*p�����X�p����mER�JF�#��<r�.�
���5rzHk�v����y���%H��~���[N�rP�
W�q�R�Wc�0Vꨎއ/ �++��Tp���sQ ^�فqJ�̳kM��4��Xe�|s���{R�ǭ��&�ާXy��&'�ܽ�;ч�k�;�#p9K+��n�c���� �$:i�,�ә]��6�K{3p&%#KYc��K��c���N;w*�v)ZK%!5��X�l�oOQ(U���;�`��w� њZ�F�1�W��������1����̣W)>:�kU��n�ǯW^��č7S��;
�۵_��l��I{=��*�������IP��k*=��]�ޤ���uI�g0�G4�|6�̏*�8*᫔�t�n��OĊ7}�d���/NcWu���c�(����r�� ��,^q�;�����Y����7���ta�������^8�G('�o	�)��n�
��g/w49������b�v�J9�u���˰�!,��s�e�C����aw�vM���4l�p��2��i���>�Y}��������4Kų��=�d��Po�H��B��6fI�����A�MTMIJY�E%L�VfP�LS��DM��EY`MQQTVc�JaL�T�EQ%DPUSMMAESJMMAY�E��Y�ETAMAVXQdb�%TQ��^f1A�����������$����r�
��3b��ʢ������`�l�(��,�j� �#*�����($��Ȋ
��&&����2ʈ�*�`�	����)��"���*`�`���L��(��*���"	��J*�����'&�� ����"*�f&���#$����1)���j"&��L���7��f�]o|�fo��:�+g$neة���'}á���U<_����.��a�S9G��!�/&�i����@� ��$�&hRd�JF��b
TJT�RaZS����)��m`�[���]�E�^K�ul�¨�yj ��OVRcC�Ӱ��4�2E�����h�M\ve������K�Ɉ����uf���0q�i*�
Y���7͕x����w���[�d�ɮP�S݇�5��Ƹ`��[�0}ni��1���C�д�/ɜug6�YÝR��h����?�zc/�맠zW+�y�G�x�O	J�~?M�2�Z�m�N@�S���7Y��V0�V���tN>�&Y�I�nm��^�{���z��(ME���̹OUosuM�4�������f�;�XW��.�8˱�b_��lk�[9y�y�m�˛7!�]cB�F���7�$�f	BH{�v�{`�m�19�L�1��6x�C�Pi��I��t�D��۳��ow5�Y�xlC� u�Z�N�?k1��o�+�uB�u`�rC�W9䫐��y9�ޚLբ��6������L\?s�>L6ä�b�h���Oh�aꖶ�JBנ�FDut���4�?d��.�jD��G\={zq��	��8:)�����	�t��v�a��:@w�����Bu��j������2���7�\�-�T��,�<�[;1��g�S�|��a��������K���(�6lm�s�K�`ɂ")�Kw;j������E��6��"]P7)���o%R��{3���/ �^��g<�k�:�]s�|��y��@���P
@iF�TiA�
V (JAbI�iP"I��^l
�{�ͬǄs_�)	�F�+�Q�g�u����v���d��(ͦל�c$M���]�O�϶��^�<CH�3�O�Jc`1�NR��1R��ټz��xOV��J"��v���d�^�q{��ӌ��P~�L�c@B}�k��锝����/7E�IJa��|��	�E�{ ���}ꭃ�s����"!0<�.Ct��y����c�t�B5(���^�eL���y��01�[��:���C�������8zhfƑ!g���&��"N��(q\u£O#(,h�v�b{�釭5Ϭ��%С��'��dy�{�ɵ���^ښ.�Ű-�|��&a�����fmE�g��~6���?Z��Ӈ��#�F��`�>`�_�Y�cQ��XS|:��m�3�M�J�aA��iA/t�����,�[��GH`�à8"��"P�S���S@�:��d;2���/�Kr	���ϧ^�L�5�,Ľv5&"�
۶7Y���\C2LA�{���^����n�f�����e��^�;h1^>?�V�;.,?���A���\��ͺnl
��W���i�7q����7pN�?c��|[k�!����/:@�y�j��Vٯ�*BJ*C	7j.��o:d��ŉ��r��P�]O�	�wwi�2�F�\�B�]v�w�,ƶ6�bb�!�+�r
��b�������UO�T(B�B�
T"i	U�@�G��}z����`h )��}b!��w�a�����boʰ�UFt(�M3�X��D�A�[���=E�*�ڧKk�TF2��>��o�b*c�=�"KSR���>�*ϗ�pt��K��k&���~�Sa�~}��Lд�a�䮂�K�y�i�l����U��ï��~b�~��	m�Z�J�>�U���9�5x����fڇ$��o���S�9A�ٳ����t	w�`qm�0�\�15m���7��t!G��N0��v+�;���d�����(�0�,:r�����`�F��/�2w��W�^B)�͕00����2UsW���1,��Fi��R��b1�I~ů*�k�_^�}eol��[��y�P2LIvl�&#��=�y�?D�I�9�N�kss���3�N��6]�[P��[\vO	TqZ?J��J�@Xk���k�~}��S��.���Ȫp��L�id�Z�
����:�NV7H��Kn&0���솋a!���K�צ86�k��s��7!�rw��F^��-R�>Y	�^�1i� �+���bXa��-��}j�/o3��[ߖ}����#������Q!|M�B�-�:�;�v	�	��t��c��7*F��,%����W��*?��)�YR�B��y��^b�3�-p���ńh����(�K�/:�B�a�2��U�Ezp��^ϑ�볾9�՝�yߣ�>$hD��F�J((Qh@d�J\��Vn��"�;;i��i��i�k�vQyYYK�T�8Z�8�;���v}v��*����^�9��ӵ���=���WU
�6H>�z�k�R~kL�z�s�5R͓N�A�@x�n�v���77
]٣��!����v�E�OC��v��Ԧ@��u��x�>6=z�߶�K����3�N�.ik��#�B��?�?3�-�����c�������%��W�e\Ce���t�7{��+�D�1\Ÿ[����s�<�� `PZbac�R5��)o=�ͭO�*�5͵Wj]HЊ�4]�,Ÿ�w�,�sͼ"]�CF��k����K�e��L�tm�ggi�wO�e %�kǤ�jM�\��M����y��^��os��S�-2r*���^Ф!!��[o=�\�V��H� $P�1j ��#Ͼ͜dwZ*q�b��q{;��q2E2����4d���1�3r	���j�����0�	��	d��F��l��y����;u}����Ã��Z���UwE|k3�>v��u�P��G���eN��?����q��-��f�9��@��fĂyF�Nȕ�J���i�@�fu\٫n��]3�cttZp�ݤ�ؿ[��{�T��_,/PU��!"�ݙ�[)�5V)���t������p��'Hqk�,;[G]��>�(�O��L�P�"/H��x���Jݱ@����$
�  �P5�|�3~�۽�,/�vD��U&ˮ-��.P� ����]4����r]�ChP�����;f��:�˞�D�W�W*�qv#�O�"��o@cH�H8+y��f����w��;r�ը���/L�wI�˅9q!1X�"��L�`���yA��������4��w������9��`��@�W��0�u="f�X������f��ʒ7����*#��É�˧� hq���7s��?U��7�`p���;�[�\��a),f1چ2MWbٱo���u-��ʨN�kû4ip"1�8|c!��t��^���\��ȣ�̖���T�����$�O��z�2W���ԍ�a>/v���n�`�}n���>�a1��ͻ�hM�lx쎐�b0<Nvk%]ԍ�+��V�����Q�P�l��z��fpF�4�|NVp�ζ&"Zb��ꆾ�,�x�0�AjU>ci�nܗf��j[���\�s�D���`>G\w����Wܣ��E��x�/�Tú.��Y�Aܢ¼LIv��]��1���+���>�?�kE_L��J�-�cMOe������qg�$輺k�H��J].�w/b� �q�h���ꙝ�%qn�g'��V�n�����m��J�@m-y�Ǳ�?}v�����G;�������s�]	��;� �*��Oc����N[lhuY{�x�Z���o,�JE"!���Y��d�$b�BI�B ������l�P��8T	�!s�<��#nq��a�2,�P= ��8A���b�cFn�	�(Erp��W�sM��Pز&�(lg��&P�.2}Qx��7cZ}����fxz�t��ʽ|c�_쾽�w�P�$f��;\e�5{�.W�)����ӪWn|o�U,��F,g/�hF��+�[�v>������C� ƭ]
V�z3��:���?M�;��F�?(�MKh�lҬ����{�4Ǘ�T��HJl&dE�B�ܣ�k�zv�i�S�;@@Ŵ�Ȼ���U۪������������<��������RX&�)P���������,���*q�9�!Q���Y���!Ŵt��8����ð׏���n�xd�.v��2�����/b� ��{��~����֙�_�5�����r�v4�T/���dQt��]D��ٻ�-i��X�5��!�j��A�,�^�=4y��#�&�6{�v�v҇8n]�*J�"�p��|��(����ƗJ��'��g��{���֑#[�bK��z=�v��K{���gV��뻭]�T��_u�^��s����/g��G�vw/�����37�$�����T]������9��p�ͣU���]�M�
LᖱZ5�_��q�OeK�n�Q�Z}��>ޫ���s�s�}����f�
�3��8og'm�i5�z�����0�}�|�����3���5m��Q��,��5j�w:��Ӈ�p⼄k�ty�cS��#^T����wUXF�ק&�U���[+
Uk
��(%�S����f��E�~��
���f"�eu�n�۰�>��t!�w��ra�q�7:���
����:j2=�}:��siܖcu&o���ެ�2�9�2�� �~i�Cξ����۲����/��	;i��/.r�]+(�"�?���gR���SDͻ��~���Se�^����F�cf�]OeJ�ؼ��˚���s��B$Ӵ��o���T?c�=� ���{d����_�~����6{����O�hȶ�?o�](T�f�.��׹�}�-R��#�=OH(M{�� ��i�Ef����}^��Jzܙ��⩛p����	�$r��l�|i���"����E.�1p��3����oxN3�t9��yq�Ꝭ`U��K�!62b-���Fq�ј��{!F�&��!�6�w^\�o׋�pP0[0j�4�& "G-�FB�f�A8DĲ.��d�^�Vk��gd��vr2a��q�>�ʽ4U�R��]��!X�ɸ��\��9�9�he�߯2�5��ueVn�V:�?|����0�}V+A�!���i�Ȳ�L�򈪭m�����yNģ{�R	�$^��u�����Vf�c�ڴ)��_Gi�{�v�Z?��y����9��yS�����G��ש���$(����a0R;A��<��S��,��e_Bf�1��5��uX������
T���y�ϑp�= �5��ۢc�)��[��z���[��6���.ר�E�+T�d��R�-�Ø����}��a �O�<�M��'k恫y�/e_tL��6!�Uy�>%�rt�/I�R	z����0�0\��C��J{:�]rH��^�C��Bq0��_g�[�ݪ���vQy��5���zp��?h5�Hxn����?�X����:���S��#=�y�C�~4U
�V,�ln	�k�L����6�j��cc$5�n�^�^��ȡS)���̧a�?��ݛ]��~}��Bպ�ë��Yc�G<<2��ی亳o�ѓ{&���q����H�uZ��x��ŝ���{j>��47��Q���T���*��q��%����[��b���4G3�`PZ}�\!s_23m���r�QT��q��$�W���L��]����y��CdK� i������??��b�0-!��[�J'4n@H��w�`@��F����.�Ѱڭ�cE��m_)q�F*�8�f�<9������@3���}1� ��eoF4ln3�:�}Z�%vE��R˒���T�5RJW�::�����������L�Z$E$:�� > ^uosg�|~v��O�&q��wG�2�3Ey�I.�
�d�v���i�q���ŷ��
]�x<�!.�5�pr�y�-�=�_z�o�8֝ ��nd
�A�#9T
�f&�O�'߷��}�~C!�:��x�`d���a��T��&򢭫�T����	Զ��2'��L������vP��8�c=��YQp��fp��v�ɉ�i�Y5z2;Ph}�+�����Oܞ��d4;�C^�D3��<�(b4)B��[|�'�T\:����z��Y���.����->��^����Ʈ�.�*R�Y��I�9�N�2)%RN.�8�{"�t�?�A�m���Ġk������&C�:�÷��.��J�,`&*��"��D�7p�;�0�F#�c��^���ɬ�! E�֑�sB`�>�,�_v��RS����E�.9�-/#[ͭ�s'��zuU��=<�g�yߙ��8{n����z���]F���ũ0���\���)=^��]L�kV	g�Ӵ';���v�)�qD���cm�t�>�
|�^�\W:�YB���N�����<�3�=a��W��w�q�������&����7����y�j� �ONV�i�E�<�l�s|��BP���mr"�ح&i�9��=��:ju*:#�SMx���o��ٶ�r�����+7����co�ڊm���lӗ� ��-���e���.����tuY��dNwŇ�t�5`+�a%��[��[�B�)T�-ԭ���^�%22ղ�gM�7��Э��%W�%k���+^���֪9��z��P����?�1��|ݒ$�J9u�vtuU�3��������sW��@߂~�ױ�a�t����z����ȗv�n3���v�"��z+s,ZC�w�ss��Wt�t��,+�K���`q�kׯ2�'D[
݂�U=D�hGI�6����/������F�v����s�Ǹ	foE���	�z�Pl$0���6�q,j�ʹ�4�����f`P&Beā��ؚ�Ƕ�|k�$<5�4����������Q6xk���h�M4�m�n��u����9aV'�z���]��L�T�į�v���t�f��r����T�D�J��}�.b�μ��BcN	��!dND�;�]�30���vDK�gLl�sk��,i.(&{Fg���uȢzw^��V��Ol�1�+#�C�37t^�<��!S$�K�z`w	��/��V�!I�Q:��JHW�R��ټt<��O������yz���w����z�^>�W�����s���W4��G����7��0�7�cZ�҉�n�X�5���ݜ�͇(p�M]��bɖ{St(���&wtJ�}w����	��٧�����3��s�`Kx�����6��y]�#z�:dT���Q���=쑜���m���	���Q	��Ȧ����y�4n���D�5>�8 )���6�ʀ��}�\�Z�Z�NgMvQ��^���k"K�ʳ��-�6R��_<�����w`�n��͖멃l�9d���YB���-<H�u}��5�/E�U�KQݝׄ`�ܲѽ�ˆ�/[�ڀX�|C����f�dE`;�d�`v'��ٺ+�?�����V28��g�k~>闦c��@����9u�7k �Z�J|N�#�T�x�J;3[�A�F����&��	��:!<�;����nP!3PHtZ�86�sh�x�
/N9-�P۽�Ǫ�d�6�d�����&�"��N���G�Ё��:�o�f�H$�S�`��ܚ0��=Va�N�#�[��+\����4EpVL����V�����!G5�k�U�0�Y=5-<�-�y%�݇uN�YY��Z��Ɏ\M=�wt�6���$��MfS"����{j���sx虨H&x[M��g�Z6(SqY�~�2�IC���wj��lBF��_R�:��L.&�������M���+M:��f5k�7y�X���x�(bi�ouLn?R�PJ�ն��B�}v�*��-'+�R5��Q.��mء��7hǌ���b���*38=�􌰞N)�5��8�>�î<�Ժ�zv�m�N��,;6H�\݉��2vF�"��=�;e)ai�����b9����;ǈ=�MQ�y�5ZNV:k2VbS"�����ԭ����;[J͎�Q��+J�^FH����7gm	m�mfՍh�u�#�G���ԬB�������o��☬��,�����Y}SxW�dꛮf.�rC��g&-%ʶE[���2��:?wVVp�5kt�" 乴:�ځ-�xQ�Hք`5fY��D��F���Y�1��V�\��ج(����:9�Z�+S7�ZE\ܘT�r��8:�5}�R���dtn��P�u��&��%W�֥=���i�9=,�on�֛��X���mV�H�;ΎUก�,���f�Té�t�*�"�h��p�� ��Fj�D��ڳ�� ��d������P��)��\Z�v�ϕU�l�ڼ�s���k4Ga?�����񆳇Sǣ�U�e����30����/��zr����C������ݲ7Ln���wR51����y�na�xާ��/o9��3��b�������T�O����|o�F	z��X��2	�(7�WQRZzi4��f�u�=F��902qbԱ��bL]�1ogp�1�Pܮ!�`�r<�ݰ�����&��4�$�ByHѹ�e�O1�拜��̾+��3e� Tp�!J9ƻh��a�Y�˹���M`�,�*�m�@��� F�$%�"T�U!�I�Xo�.yʸ�3�.����*H5a��`EA�e��f9LADՑ��K4Q5QXD�T���j2*2�*�*��b�*���(�)�"��Z(�&&����s"(*����
!���*�(���\$��*��Ɉ�&��)�
��*j��("�jr0(��e�"*)��RI����"��� �h"����"�f"�(������������#(*j��(b��r�*%�(*�b���(b�p*��" ��#,
& �h&�*���3	��"��"�)�b��!������*���(�����)* ���,�
�����
`�����"���*�����i�
�3(�h�0ʩ)"g�2��*"�VI!1UMUUTUSTATQQ5�%A3c�1I5Ya�QMTMDQMW2dLU1IDUDT�EQT�Q�����{�ͣ�YD��t��3�V�2�5�q�[=/���k�m�,C�;Y6K-�����hN=�z�⎨h��u��Nl�/��+��� �_�����><�����ٔ)E<[�[����*`�{�k�;�R~��x�I��O�Iz���vꮬ���L�"��]Ds�c@�f�r�k�r���J�W���y�.�>���,v�Wv�nt�V��}A�Su�����-���5g��Pͭ1Buz`&��a�G��$�uM��.k/M9��Ê�2e�Y���Q>.l.��C�Ļ���>a�6��#[����V����2N���6��M�-Cyk��	Te��#��X
�w=�9�������x����ü�~��3/�5xy��hj����e�:�����V���J�%��ڸ�w,�C��?T���,s#��g^fV�l�A�/���C�~l�f�}��d`�Ll'��c��mɈ����MM��z�f!3rb�;�
ֈE�q𽍨d�^ݐͳ�(�Yx��7�'*����$�5-��)�nc�B�
1^oO���殱�GD��A��*l��Fk���{6g���x�coK/�Ө�v�~��qhO��v��-�;P�^ȖxBK!�[=�N}�v��?�,}��5��M�ݓx���~Ue��h.Z��_ ��EҼ��4JI�y�c�kڔl��M�$^����SݖԪ��m֗b_=Ż8MX��t(�a�]�������/y�ӥ������{��(M��{�Ejk�k���K�m�w���a�����Ŀ��=�����P֑���n���t��K��EgN'�^mṡ�Ö����@gW�/umwp�̄(�|�U>�z��͵jJ����[�:��6�r��l�z�n)�����z22���S�D;�`��^!ּ�G���0K�b����)6�1�O��(�0T��wb��{*��m�䩷��x�^��x���0D���@D<�[ ��U�OЂpK�"���ٗ�y��s6����$���Gc�W=�����2Eg�%;6T�0]� ��y۩�C)�TSm��s-|/L��t��S���%)�����.s��f�t��pLpd{(�T��J��$��NL�npa���wT�'�9�NP��-�Ú��/^|�>�E�A�{m[�}�F�SF���4ݳ�6����Ƨ���P��!7K�����N^ƕ ג�a+�?���LObƜn��\`�mhRýO̡�.$C�v�mt�wj�j㲋� �F���)Ē��Y����ߍsb�o�S
]������'�:�v/ǦD��S�k�wJO̴��������DݧS���n?�v�p�H�.�ݫם2�Y1�Mp����]1X��3����X�}�Z�jt!LWڷ�yH�����K�`><9���k���J�%
�ٚ�Pq�3j����ݎ)�y���u�;�H-�=���R�fKw�"J-��+��ح
���u�wM�5�}WR���wfS����?0!����랧��������<�m�l͈*:��E��Ө�ݰ��}W���������'�~a�ۥ�6{C���|D&->����6�����n�C�v�u5{�	u�H9�<\��i� �	���Z�{���h�gh���43�"���M��di����u��M��3Eڀ&Y�qr�3�DYz�o`"b�2;�o���??�rW�>o�-��!����4\S{_�� �@̳L�@�]���A���i�ֺ���URg��1T���Ŭ��L�	wC44	���ؗ�5s����#$U�A�P�4�[-1M�1uk�]����t3'���+E�:��e/ߋ�9�
�ݺ&�ʊ���O�"�^��m	�G�����bᮇ(�C��g���C*.��ft�b$��x�k�:ɤ���O`Q,�R��]x@�tAq�r�N�b4)_�RaL��ۥ�w�1��-�
�^�V�}T��J����xm��e}.�N��nr�;���W�T���8�Gd[B�����Ԅ�į%:�.��X)��G�:m�1s�ܮ�� ���:;O���\�z�M;�ncq��e��ܮo3�_Z�N�iLs>�C�ȹV�o7e{�u�:옛54�Q�ݕ��S%�Qk�ʡí���®�:11Y���/]���xx�ӴOLU��|!�É��A�v����v��T�g��@1V�"�j-#���/-�٨)����SK��oQ}�e����c���pG?[�eZe�nc��Ͳ.�1�̬����F���Z�f���w	��m�s�韞\=�����%�?WQ�D���yb�5��p�� գ�w��Wk�e2��4��͸�~p��%�&5:�������p>�����]Z|
��o��0ݝHۋC
�Θ�9�
�X�}l���p��mn���������e��[j⪵�R�b:���C[W�4,�0�Sk��'�Z��[�maLs	�N�q�'���N��.C�_�߈{��'?n�ɡ��I|CjY��m��@�~�װ	�i�Է5�w��_��g�{�dT�·O�����o�D;�*ǐ��<�~��ٵ,�:��n��(��LIv>��c�LC�n���⶛G��x�q�˛
X��l���yw��Eh�/"S�
���G�Y�fE��= ��S4UK#��^���9(Xe�e۴=7gD��-p�c�2�Yq"3%'�zǦnF5
��=Ѩ\଒��wՆj�����-W>����𵸍���T��Q*���"�������i��6d��s�U��+v��&�J���W��Z{��u����>k;�3%%���ƒ�$�Hi�gd7R'QR���'�u����]M5�	��S��9d=�> x G�^ Eɮ�<ǻ�ѿ�0�=�w̅�F��덷M]1p�)�0Aaä�D]�{�vF�:��gs%v�^j�:�T���B���2>�t(�J�ߠE����d�1�t61��g,�Z�x�I����ȳ�}v^]8ܮv�����Jl�^BeѡI��Gc1�cռ4Z��zٹD_�ҙy��_�Z�r�V����ݕ�E�<�����ħ ߒ��5yJT-y���	�B��̬�ٝ�u8�]�^V������\� ��l!�3;�od� �1b0>�9込f������_C[
�[W-�~���s���A�l�"�|�v4�U}Eݟ����/�؅m���ϦK�R�Xm�cG:��4噃k�ik���kW��&4&cFݷ<U\�t��]v�P[I�U��^�E�气5�ҡ��w����CM����{��s���vn����T��}�:��:rEh%Q���;�R�έƱ/N�7���gFp!5,nN-|Q��;L*<���\�KoX����Ju���J׿#��ڸ��f��y����5U!�~e�a�/:
�dލSM����OMK��o/f�������D�(l2�	�0�[��B���wU��j?�d��8<��+_e��Ӭ��Q���d�9�&$|Fޔ��:��gv��C8n�kS��̷����8�2��ݱ�aF:����-5�P�'Q����yz4������@`�
����k��d�6���M��Rc`'���gӯ	]��r%w���/-s!��ʹ:,3�����D"�!�_�� ��v6��_��:/2:_�XW]N�:�kۮ�� n��o���)��u�v2:%�r�=��"T�{ڌ�J���i�^SSK�M�Ojh�`��@qhO��v-��ױ��g� ����sŎt�]f�mTڋV�m�S�wH�Ệ���}%��U�B��K�y�i�m�k�;˝ٜ�=A,�w�����
�!��"22��cП ܙ��.�3l�2�*���	�$r��͜N��^8�
I�zd�w�۝�6���(3Gy"���k�ߢ���*��V'b�=�Jl�eM^�f�����2�4`�¦�7u�0�{�Bޭ�^��;�'�"X] U3CC��dGgH"�UsP~���z�spU��¶�F���c~;ܽ)R�=ߦ:����৷x��vl�0�.ƀD��� ���w���ʴi�qtD�\�����H^�x�$��.�c�0�g�x�*�a��?04�<��qZ�+�b��T�ktO^8��|��Ysɝ�y�zˏ:�׆IF^�s��v���M[���VS��(�bm-\nN��@��P&�q�|S��\�b�cY������L0E�ۺ�
��o:<=�Fݞ�7!YA����Pl�=\H��N���$Og�>�.���w;��O��Rr���m�Laz2}A�@ży�r�<��[d������bb7H���^0�v8�_I�O�(�Ҥuf�v����L�Yݗ�x�9��A��gd9��k��M7_�Us]��^id�e/@��{�Hf���R�����^9V3�y�u�,�]����#ϡ�?T+�G��)��6��	>��T�ՕF��Vn\�7n1t=#s�U d�d��E	���~�O24��ʧ����i�jRnC��}��]�L5wR,
�c�=>qL7��i�~�����63�~g�!1i[ӦʸA���+P������?W��N��i�D����nX��� s�<h�gm���!1~���{q}챈���O��S����7<��hEx���@,Ÿ�w����O�Cl7e�����D;�`켂�i&:��m�=�>��f����*a�m=�+0vB�2�k�is�װ���)����++�7�԰R6�~��.y��v��:A�A�����z�]�r7����y ��Ur�/��r��Q��D��e�� �'�^1�:���TἯn�y�گQa��������ݴU֬���&I�/�$�%�}��Lw$D�)O��B�vG6�j�
�:�W'�9�x����B/��<����7�W��x��x;@�	W_*ǔ�~$f*�3r	���n��}�:��8U��{��E2��8��8>�](�3��{l*.ۆkA@��\e	��a�D#{$3�y�7wo��{�������Z�V��):��Фޱ*�j�q��.P��y[���ϥ�Y�<1榭(���ҙ�L$�!d�p��)��?Bd�Ø���4-X�I8���a#�-�c����:*�oC�fo GF3�A÷YP���6���&X�b�@��wO�E����Z릻i�K�����F4Ð��`���e�i�%=X&m�u�y{'����ew.ۘ��1��y�'�������p��r��^S��B���e5�T�cs��ln��B-���\�z�����������8Y��X��q5�w�=�ή����m�9y�����2P��Q�<��ƷR
�XHso�|�����9������.^b��6{��j��'$k*�T-2��;���k�J	{e/�4��֡�aߤt���rV�ʷX�gu'��Ǽ�]�@oP��|j�f���ǽ�f�/3lB�>N �ฬ؈��� +wv5�_`�T-�/At��s诺�1@���N��r��R��N0lХ
{�S��˳6�+r�(TcG5�╶6��(���28�Njh�f�խ�E�o
�u�π��+��Gb�����;Om��=�f���E�1Ԥ����i�f��.�1dE�kg�t�R� dKϢp�XHy���ʖd�wC7�����\e���e4�b�d�߿8i��u�_Q���{�.�0&tFv����n{��(�aّe�FN����cWv4^���;C�P84�e�A�ʺ&�֟Hv��`Je���O�EE��&)"Mޭ���e��C�U� �U�y�\m�j鋇\�ρ�':Z_Z��a5e��UQ�J2a����|�1B�У~	O�ѕ��S��?MP����侾��b�6�"Y�>;!�8�\�KsP~"Se��	�hФ�%�vzw^���,.`I�+�u�T�O�Ƴ��1l�A|�	���G6��%1�9䤰M��ffۆ/�n���-��FNc�>��z��x�������O���;{�!'\���Jk�h�5uM�ʍ4V,n��E7P*L��^ˍ���c��փL��$D&����"Tx�|���!��O����d/�[�w��c)Ӣ���DWe���^�n#�B����Bl��_d���q��Ė�S"���{��,è�v��lS\��c��3dx
��mv���E�Өg,]���7�o�0p�e`����ݶlޠ?�z�[���~�����-E'L,�Qu���i��?o�{j���-�A;6�!1���<D_�O3�j|���T)N)�ěS��oE��J];�1�8�x=�C���a�
��nmvq!����^��GD�;��KW���v	Te��dw:�WC������-.�R��}�n�7��uOW2�������	�޾�-l�Еk
��{	A/t��7Co'��m��ή���Ȩ��(d[S����@r�߄;k��vm��ΛepU&6�S�$����Z���{�،M����iz��5�.����Lg��t�ӟ؇�۪�߿hq��{|��u��z9��5j:����rC���+�C���!��D�ǐr�4>"T�z�6�[y1X6��'�/��T��ci�C��D�&��`�-���.�ĳ����ĢJ%�;C�V���m�h�Yz�c�zǥ���5�p�4WAa�t�R]�ϯf��,s�<4�<��g���FX�:�Ob�tDwy�S�Q���~��O=nL�W�%L�c���R�d��;��ӷ�Ǘoo��>><���yyw����С������銎�� �1�aХ�V�G�#]��<���85U��+�sL�b���_$�8�Tά�C�5u�X1B3(R<����p���D����a����u��s&�ϖn�L��JP��t�/~>R:��w�;��{���;���6��|_A��ٽ���<�Q��vU-֢z2�F�����R��6��Ȋ��@�c� �<�]J���d�ƽ���f��E�漄1���i�=uݸ�J�2D�_ �)�� u����՜i�弇�R�&SNJ��hs�������+��6Tޒv��9x��^��{��ص�F�E�8�t���2�7�^K��]RN��83d�������o%�d>�[�ܜ��[��:��(��{n����c�X�7���pnRY�7c%N��oWa8.�z������ge�9Ezê[7FvG����!�k����6@���p��ޙZ�o(�����FX\�Z*�)�;r���|��B��vZ�YWZx��9�����]p#��n��V���2�u㱑�pn��� {D���R�7G�+dn�F���pe�t`wZՋ9�g,5�_]����ىYWO7�4����sm�-nQ�A�K{�]:ڔ������YeB�kS�X4<Z4����i.�<�!Cb0��L)hE6�kd���:��i�'痡lh7�C��;Ƹ��<�Rx%m;�@K�����O�m!���#���d��Xk狡��rU��q��j�'��`ivɉCf�|�rW
��ՎљD���u}u\���M���.��D�9��g�Z�q�mc_��.�7S,�G��7ME[ t0fkTV�\ۗ8�k&
��r�f��
�T:`�Z�ê;=cB�C阤�v���b''s -_���Y{��>)�r�4��{NSC�X�V�y���8.����0��v��v�-6���^�!G��hwvO��*.�L��Զ������1f�7��B(���ź�1-,9��Y�DM��Px�z8���;;�i��s����2��Q�,���v��0�u�KWp�U��V���+�j���|��^Է["æ���uWK�tgv��!����XUن�m��$�7�1��]��ugud}�����c��}���$u��c�ܩ�������/��s��G��j�<o��.�<�X{�-�.��8*lո
@�k���K�.צ�)���EN��)r����p�;�$����	/��3s{E����Y�G�GL��N��vޚ�rC���4ŅO{rf��)��t��j���Mi���d9��;�1�\�YԆ���ކ�����;��^�2�X�7J������;��󷕍���]wqCV꾬��,>KsIL
�y�D[\r�Ń��h��y�6�k1����:6�1���n��؎Tf���9z4�7�;i��� �N�*�E���T���ϻ�f��û�^��)�� z�����5K3LDMQDTEM4Q�$���R�&�X��$��"�i����*��"�)��*$���TLT�̔QQ)D�5����&j�����&���j�h"Jhj��
 ��"��bj����"�¢J#X�K̓4�MDQJ�E%4�P�Q@QDE�ELSHL�D4�PD�E%4Ĺ�PU%AKM4D%Q�SSA!TRPP4UPPD�@QM%%4��R�UDCK�PPLSBULHT��VBeTEEMA1�5�*	���@c�IE$�ADI1CAE%TD�DCR�ӐS04�]�MD�L0A��4-R�I�AE�DQR44QSPD�V�"*f!����(�fJ����������Iے}������i떬A�,��7��kv%��B���U�S�9�n�����۩��ž~8rw`�W3U�����w���FN�د���GP��V]?.�w�����M���T�q�Ʉ�L���g�t�����������x�`�z3���xOB�� �f�q ��dC%W7= s��a���M�=��_
�Ap�Ĳ�HĲ�d� )���<5{gOMn� ��Q%ٲ���qf�Qfp�P�����~�d^�'�����>9�N�@�\����vO=�62P1����#�ӯ��<�"ٞ�^���l/�t&nS5��`p_Jw;��O��Rr��E*��,9�����}
]�����7��5���,#��An��۞ܞjOxT�O�[M��zNR��.N�@���6�ӎ]�t�y�T��e,�~t)X�t+塣�q�H��L����Ӆ�e�Y#YK�jf2�"r�JjX����XP���d�U���V��(�<ò~o�T��VjE1rfڋSnN�D>!�x��n�"q�|�v:��G��T��U��B����_QDi�����ç��;�r���"��)S�E�Yc�=>��U� �XO��;t���.Y�yll�����z�Zc1��wW�a+��;�-�?1�h����N;�����&��p}���O�߽��3��[�Ҷ�x����ԋ�Ѥ�벶Y8�E\ѵ[S+,1C%��u[y�S�����@˽��'�,�9Qf��Ҥ���(���-�v}������{��~���W{��m�T{�?W��N��p��_�$�̛E�nj����i���l>t^�Ưs,,gd�Ŵ�&:�mH���!���B(4]�,ŧ�q'DYx���65=�+�L��h���6f����ƣ"]�0v�E�g�I�	���s��fY�h��K�6�5���\5�u�ᕝ{I�
{k/C�m�׶E;�e��ȼMG��v��b���W��_u5���C{��mpmd9\�j�g�b�n@�t��N����?C�=6��r*�f��֧�n��l�9�|�R�_����'�j��$k��;����\d��%�I�['���u+cp��ٴ�]���q��FA��2ǲb���hR�T�SP]�ƯuEê��~�������Z��;��o2]�4͗0y�@�m�7����2�b�%�(�T����l��WΠ)YW�fsjiKE�g[� �4�rC�b_��ۃH��v��T�c	�S�i�ͷ&gW5��:2nr%�g9ٲ�X��H�DS;��`�>�T��}�!�G�����w})T���Sv���^R�e\U�!��I�M��n���M� 	�r,V���WjhS}[��q�ǰ�(:�*|���¬�U�����r�`WoQ�(u��8��2�jZ�}JE�q�f��yQ9�T��|����E�κ�/C�@4)���$�}�~����
���ݏ�2��}�^F���f�}~p�|��F�Ð��R򟫨У�vS����}�]ٜM�Ŭ2��PYs��Ғƹm;	N�R�X�C�Y��i5�O��P���Q�a�]I��K^�8��e6�N��%Qa^Y��j�����^���sۇ�p���>~�B���2)��Ee��M53AkC8�-���mv���
�\u��Z����_�h�N�{�}͗-��i�2���9�z[+�`��38#���O탛r̶�h��J������I.%ڶ�5-�Y���w.��3�=Y۪{*W���k�g2H�x!@x!0���~Ɇd��f�r�
&$�Sw^#��g3u�W-yӇ�<Rv�u�e�@�lk�[:y}a�q�ǴLB|aB6��`�n�����@�1Hw�~�D�-2^J#��i��q�<S���f�B,��̔�x�64�痉$S��73#��������y� v5�ջ*��W��^�U�B�#^i��t�:b��=z�/*N*��L�W�w6�}���W쫇�UF5�-m^Ԥ-|.�"��J�J��}�똨s�G�wfK����oB�XխK�ʛ|�渝9�0��G%֕L\�U�]q��-('%���SUn_g�/_��~2Pu�k״*��o��;F�Pc�pE�FifYx+BM[�]]�s2U^��&��-�Q������O��\j8)œ,�$=�A��d��)���ʿ��?R��ƴ�C��ig+��KsW����~&Behȕ��xZ��k�|��E�M�p�Mn�9��y�*q��x��=o��6-�/�0���>�S�@?!)���Nhn<qA�o�x��}E�nU��];�.�l�=}ǎz��>��О�|��By�hH�5���M
��L�f�1,��D�/2�d]ye�%I��qOw0���։�b�Ct�!}�psj_UR�5�z�'��
(,��!dRt��F�X�ʖ���0i�3׿8zh�
����<eo32���)*�g�۶�����YIΡF��w�5ٕ]/G"��_���X&��ߍ2W�U���I�� o??�"������g0c�>54ň,�vk���`[N��w�U_�E���Uj�w=,�̆MFd�ܚ���?H�ݥ4�\:��x	��ul"=Ú~�٦�}TZ�\%Z��^�I�=QP��˝�>�2�q�[7������郔:Cp8t!�����d�6�׷:m��*�n[A�|�����K�1��D���f:Xgb\3P�`<h�^@��|/{P���������qa�փ���Z_��v��1����+���S��-ӵ d>��	�P��ï�D�9�4�]'X��<��0��1�֥Vy��������$ć2�R(��$JY.��ښn�gG*����2%:H0��y�|��.ئ���\g^t�~4�߃2����� �zK�$@:Kϰ�b��!�c�����4>�>Ě��[��mN��;O����Q�&CɶǺ	Ŝ��i�K���Q��?h�ֿV��lU������7=�ƶ���2�?_N¬�}'M�mV0zK@���R]����v�|�k2 ��m�hۼJ��ũ��@s�<����FFS�S��ɛj��m�a�U��	�!Uᦂ!�k\k�k��݆��ȃ�?��j��_��Mw�X5�/�yq��X�+���q���%�;EhƧ��̋���n�X�6��k���gP=�Bޭ�z��-f
F�"Xd���l64tlK��X���7�J����̃� ���%�{H�2�JT��#��{gO4��A��Ivl�����ʼ=Mҵ�C
^�iO�$����It���t��^IRkg�m|��\�ȫw*��%�d�������b�n�0���0�}%�WuIؼ�)7H��Kc�|�5��)*�=��7��y�i�����:��&46���I�
�g�6��LZr�2�K�}~�cʼ��j�(��5�f�,�/����	u��y�ōF�~�5*�mM�K�)����DZ���ׁ��>�m>��}C�e9�Ѻ�b���Wnx��LD�8�H�f㤶��f�/���D&'^��`�F�Z�L˅\��EqB`pl�K��s�^����q[�vk&���n�0�r��>a�H`�Y؆���mt�u��\�~;(���!�t��41f��ڼ&Y���tL.zc���v�ь��~`�������\����Z�7<�ټ�HT_M�ɬ������$Ɨ�9����@+�A��l��wf��^p�C����;E�v�����Í9Hvw'��
4,��Ë>2�@��W_�W4��Xs�{�&ц�������C�Y��ķ��e~��X���k��~��N��i� H�v���_�9j�0p`&�M&US��DZ��¤�u�Z�f��hu�oE;�`����넛U+D�C�{�w;��,�
LՖ�ݗ6�Ɗ�D�א��h��xr�GE�S������l�`����Y8�P��c՛އ��Ma���kmj��x]�)�d!���|W>�ݜi���2i��rx9uU�x���I�75�Pd��m�s@�eY���zw��$`�����{����Vd��W�s�]*���j��^A��ʂF���c��eEÚ��P,�=��k	m��-l��ڨ䝵�a�;o�5�nvv��ҫ���2��~Q8���C<-��u*8M���,�j��EU�)�q��4��h2]Z*�dGt��Ŏzu���ѝJ:XT�P�Ep�����3V��Y���SY=��=��T܅����q���nv'��$5������UUY���b�P�b]V�D��OFAV,~����; vu��ѐ��?B���LZ|�F�+�I�2�lQp��.z�뻦ˇUe#+1c:"z�,�^���;���{$�6�0pИ/�bS�Hеj�'�\�*���cnW>mV�9���3���B�gb���9�˲��l���L�1����Џa�Ź�fj�:�
��f�xa{�  �c;��`�=�~jeyƝ�Ӌ�m�uT1he�>B%�y)�%�1��+K���<��~g�`�ԃ��"��z������5�Lų��y����vJl�a&���#�)=XJK����<;�@܇ǐ���^a	��^�Jg&u,��ٽ ��]Es�YB͹��.�TXR��^�?t7�J�-X�B�i��]���iY\����>y�y��cL���smv��B��'�Z�9/LUG5��X�d�gG&���j:�����rڃJ��H�`�#�٣��>5�f[]�XsW�Ԩ��K�FGBu.^۔F�NeC�[��d����@^��z�Τȗx�`<h����߯*Y�u~�n��-�|�W4;}9v���gfфe`��$g��D ��%� ��e�/N{A
J�s	�a#�3�Y/~K��.
5LNyp�W�e;�F^JBLy���"�y�k�a{R'Y�5������s��;��0^6�E36֗r�$�rV�AΜs`�l{[��#.ݮLC�x�cC�[9yחx#DawhO�,F��"[0�N/�%��騙�,�y�;[�;��� ܌>����eF&�(lg�`L�\F}$*=rɖޝ��l~W��5�m{��>̎!���}�r�9�M�ۦ���u]�T��&ue7J�h+`�|�w�2�Ҷr���*B׼0�*��+�U�b�9���9~�2����BC�q�I�v�����&�����s��d�ӵ-�O�م&{&BeBѡI�upGe�F����S[����Czw^�������Qm)ė�`$$vW�i�y�?!)���&@�0��k���4ܼKs�3ު.W�O/8Mq)P�ث|����z��x[@N�|��By�c@#���C���*�z��9yb�I�Q,���tS*	*L+��|��a=k�H.͗�.v�����V+��9L��ִ��7�]�vEL/�Ԣ�tS*MC7���NZ��kÇ��E*\;�㗜���,rf�B4Bn��[�v�60�wqOK�"��X	Ab�?+���%<�܈��_�+H��{�/%���)�O��{�΍^JU��5�v:����M8��bv���z3���=�k�~6٫�{��3����(	��Pm.�������(�P��͸L�R�q��Վ�k��[�0�M
au6�0�*���QOx����9�0�l0r��!�Bvh��Sl9"��F_���]Z��ݞ�����h�����7��f=ˡ��8x`8��5������zC�z�;4گ��[+�k
��t5���I��Of�I��gK�����=��s�L�TWW*+�,ǘv�M��ۏ�s��/�.��"�p�CWu��+^z�,r�M�3�@�f5���3��t^�<��u�_H͙�7 ɼ�ݴ2ӻ5�8N\����vI/ş�_A"�&+�tE����GD�ǐ}a���n[1���D�i����K�����Fk��h1������'��pZ�Ӵ��o�P���x//g:��SL�v.����h�iiAW��z^[��=c���ӻ�������� ���s��|kVO �q�K��C3���g^W�F��g����A��Nn�}<��3m�)�;�	2�-���(�=W�*f�]�}�����9��K்��h�(�Ⱦ����J�`��v+�H�sl��籝X�o���  ŷ��(�0�ј�oV�^��'Kw��g��l��=�Yͷ_��t�5� �0W ű���
&,؏:"�V���˓���5�!��ҾK[��W�,ᗄP83D�rV<�'��nE�d���r�y󝩣�EI�]J���#*u��,vs�˦��S�2���n2:����ͬ���׽�@��֯:��&%�{���Y�J�]�|j/l���qw��q&�7��'syvjBa0R4�����%:O��Jt��H�jd#������א���[Q�g�)���ϫ�H�f֘JY��]p�lpGuI��Rr��E*��,����@�r�<uɚ�U.�G��4[2�<�:m��ۣry���R� [�����O��~b�ȹ=[F�.����+��^[�h4�A���D0>O���Us�geO��-�ګ���4�Pb�,O�qh�����[��~����O�K�@��E/~�U�����Ӥ���E١�ńٹZ琺��k�.���֙6�~W>�j��5�ݛu�6�����nj�-�t"��ě��M�v�r]W�UL�0�ό��'����/͠�XH�u5�
���.d|��3��xI
��=5��M��]����}>;I8)�KC��	���1�^�1�]w{��{H��R�3��Y�	�D��6ԍd���s��4"�3Eڀ&Y�w�ޞ_Nޞ_O�o������ǇǗ���o)���ϋX����7mdT5��؍���e�$�q�l�w[���E	h�"��_=T,�,VU������}�3&;۰��L�j^R���Zf��os���ȗ��-ή�/i�:�yt���[4����>[��V�ęFp�7�z3��x#��U�K��a��J��L���]aਖ਼ò����#��ðI+;�f�+�u�9�:�H2oU��ȟVD�)cP���њ��Ynln(\u-�S'^Ǯ�)�"`��c���;%�ѧ�Xل5}ղ0��ʢ�����j�joQ�U�p{�!ur2.��snT�����;{4��]���.�qV�f�Cƪ�KBY|�ޝ���㮗oT*ܨ�̦�V��G	2��8�gXN魮ZQT�t������*J�<����Ӊ�"F/���DMV�����F�*^^#�mUn����/�9�_Q֩1�m�p�.�M����'8�f��]���^�cZ��j6�1^�|3��<x��x���T�g,U�O��G>��f,�� �Ri�i!�ݳ!���$:�#'m]���3�>�*Ռ�ig�9gb������f�q�a�1M&���Ik�e�L'�,�S��u}��d�V��P�T��ظ�ZB�b���3�&�D�
�Tm]��\��N5q�90&8q����S.�&V�+-�1Q����[��n���^��Eru�0U\{�,��Ϩ,�0f��ߝ+���y���8�"O�E��v�#jvͱL�q_;�QE�*]u�lt(={�a�s7_�q��3)F�5paD,A8�r�ï2*��hxZ�W:��T��4�
��U�-�V����S�˴����HvVتw��a\V%m[�A��t�4�I%T�.��0�*Ʈf���N�93R�k7���#�(�B��Sz���� Q��|�"Dtr�;�ŷI�Ѥ�]2�Y;�F�5T,������Lp��G3�faü�b�Q�R�tU+��":�d��c�R�S��T�UC�(D\��cӪ��q,c�~Q;��m�C����gE.�Y�b��&I�i��:��\��y�H�{����������Ӽ�b�"�ģ�n2^RFg<���ܲ��dΦ�N:�Q�Q��W;�Y
��J�J�Cx�a汱▎i=���j�e���f�
�4霾3�j�C��f�/3\��	ɘ�����s�a��n��bg������Ƅc��a�$����f�����_�qQ=|Ս����,a��.��ת.\�j9�=#Z�*b�s�q��AIO��G�_hN���j-�W�&u<Pԫ�V�G���<)�r:��5��5�n�h!RN����a|kpet�:����;	��&C���滩^�TRh��6���Ԃ9����D��:>���(��lj�t6*��8�X
�PNNb/`Ҝ|j'/{K�"��6A�9R�3/�mɺ��0@KᬗRX}�!H�I���e<��6�4�( @0�d�W� H �H6�-��3? �R���<�)��$��j�{�*��

)��H�(���	
�*)�i�%(i�i�b�������Z�)���������
�h"�����������$�V��f����"`hh
�ʢ��b�)�d�&����)"�(�������(J)h(�$�JJ)�(��((
(���Z�Y�**�b
b��ZR�
h����Jb����
h��"(��*!�h"X�*""$�#"�X�*������QELP�A5AAUEIAI4ҕUPM%5E14�TEIE4E�5U1)E�k1�i�*�
�"F����* (��h))*��F���)���
���i]3���Qγ2/<�7��ε뮳w�\V����i�{�^�v6���u�S˸�$a��]]�-\:6�9��4�;��9y��7v��4+��A5h�A"�,�gsR*E��v?��¯�鼝�Ѷ�q.9�&!(R'�m�t{�,�4	���Uc��5=��l1M��&]���?4S���`���aql�ߦ�}]����Վ��;���ީe��fb�T ڑ�g͋e����=;Ń'�$�t�uq�^����yap0��`5�!?5�׭@�T5��v>5eFc	�c 3S��3'�h�cۛ���[v!���(LN�O�αj��۝V��w�i�jT+L��%��[Dj��c�+/+��W�Sʡ��x��Pe��L$�;���Gd���L�ۘ��##�Ik���Ku��)$}�c߀Ǧ�W����ށ �4� �D9�m˷x5�C��T�U�z�g���έ�gWSEiݩ����L�`��;=<0���� H�!?C�9��C)��VP�����]E����'e�U8���d] �4�iy@��f�~|� A�בCw9��e�[�@�ے���9�H�N����R�J���
�����I�(,wɀɆ	<;���>C�ˇ����<u��r����af���M���v��b�Í�yhi;�+NH֛�4^g;3O�5��6jj���m��7<�H�`�b�s�m1 D���%�<����s�G����Oq�UI��
�OS�9ljq�	-�kh�E^W���5G55Ti3�1b��5[|It?9��c��QI̓YB�8�Ī,(,��5j�X�}njp�w\���yYtuwT����"�3�<�p��秤sm{����`u+���Jװ�zK���Q�H��7g.o^o3��(�|��7D��h�R�����9��66e�����jR
m����{��{tݗp���ƺx=Rf�C�KsP���6��K�g2�w���x��a�nY�|�n�2%D�3fV^l�m��Z�1<�^�.z̻I�Ƈ@�r�5���"��iy�2�F�7}ݸ���k�oB-܊�a���0�	3W���O#7[�0��f���T~{��й��V������G0e���W=���{kݍf��JA��/E\�+��5xdv=�C�:���8cSS��.=�Y�"9�x�Z�D]�'��Ʈ�9R���JB���2"�Ф��p�i�g�i�?�V/�]���
�*5�j��/)���\C���֕s�-�@?)�{<�	d����z�5m�(�n͡��Oe=��cռ55���b�S�/��HvO�j������%�#�'Y$+zˇ�\ǃ�l�wlh��޵1)���BGz�U��b���^ŕ{�y������F�?td����%�_"/�Z��w�5����XW��tt���r���f���Y�^d�b(�59ʶ�� };Y��p��T�\��4M���l��bS��$��k�J��l�=lz7Sݾ;����=I�$m
��;�0���ߙ��ve.�~�bT�{�BN�1��:N�1�e^ԩ0�?E�{����}iٳGMv.���5f��uЗA�Ɓ/�;�Sc;4�t��I�tS�a��r����5�/:9b��&2r�)d�f-"�Ʀn��B�N�M��tE�洠���T?5�~L�.6��SvM[j��a��E��p�G��[Z�p�n�٤��M�-GNл�2���b�;1��ˑ�+;k8�֙�B1��i��<{r<@B5�Ha��k�zvi�X����%Z�d���QR;��h���_k�\'ytTq{���}<�'2���0s�!�?���.���d�6��v�\���J��p���E��In,�/k�gӯ@��c��A��d�fq��}��l˙�S��P�e�7UZr��ad�s���m��$�X/�����'�`Z"�7Pwe��~�v������sMb�$���D������2�@ݬ`���$=uos#�T>�/>�[�l�::t��0ŏ�{�J5�T�#�u^<u�cEY�zi}l9�1�OԸ��[s��}�D��|81@V��Q&E[��ɧ���鄷����ff�}O��r	C(9�|�+�Υ�i-ù]��v�+/
Upv>j@�M�7-�m->�_��)���^�=�+���4�/��%T�+%sqF��m^�Yۊ���,�4S�cC>xX���'縴��T�y�rfڵ%L�;��|17�Qԩ�+$������ga����X����3g�=���.�,8����\zdSl	j�f�uw.�}�|��<��d��Jt�[�v�-��ջ3��X�auC"�Gf���3j6�H�ٴ��u��r�h~��&%�{#4��*AGc�W��=5��*�l�\����[��wdA	<f���#q���_�2OnbS��R)�$�0��1Ċ�;-����)�.�ڛShǜ@�f��=,�!�2ۇ`�^�;��I> �a�_�KsVqQ*}��wy�&nqK���z|�<l[�G��M�1��w$Iz�R�#�)s��`s�v�L�W��/ͭ>^<^�V��	<���P��E��sL9�D<2ׯmt�r��|ȁ�د8ц���)Y��h�)z�Q��c8�I�wi��3��r#�0t^D>7��<�o�C����CY� *�v�bӉK�eю�����6�'���ˣL.W�"��a|�8(��fP�ҧp$j��+ZL��wU�S*�%���e]V��өn��Ț��d�nF����nl;]��\s�Q��rY�Cu��U�oJ�*�VW���ކ�2Q��`A��0%�F����I�,���`+�@�Y��-ݚ=�����,�Wj'\��{sOD�M^Ʉ!�]�	�@6׻ML�0�ό�׉��Q�֑϶�!ݶ�6�DN��d�����\�2��pDs�t�^�6���i��!���C��LW3N���+0β��w�i�ʕR��k�w5�8Bgh��XR%c��s�� ��v�&�p�S���3�E�Jf�C�c��E�s�:��.���h�q͑0��t[j~��>Zh5Z�sBԘ���ƿN�&hZed� ܺ�}kO\�o�C6�%�縶w��3��^A��Xn/�׍��B�"U�Ũ��A�+��{6ʽ�-�<����'ۢd>��7�uͫq_w�����D\:2���T$��]�mH�V��g���ss�e�3�y��	s���3"�"qĈx�l1��Dd.z~�c�0�Z2%w�QaM1
��4�w��x��y�0u�^�婟�yY�'h�q#��)��?Bd^�ħ[��{�CR���Q��/r�:�'z:����w2ӬԍhNN?L�LqR�?'YW(\��1m-������BH�.�}>%�}�����w��C��m\�\��ʹ������	�btn2���w��3��0�2����ylS��⿳œ�_��[w_���l�	�mC��$=�d��bnܻpi��W@�ԩu�r�:~{��p.qM�)=y"h7=s�w�xa9�!#a�~��G;�mS�;oos���LR�N�&r^Ys��4�iyz'�C�mx�L�A���4�Dd�v&L�S������C_:���P�`�&@�yc�	?y(,u)vû4������!�=t��(�t�`C��=1w	�>��l�P5�N��T�,��5j�X�֠B�D��v:/Қu.x�`���t�r��	��'dk*�i�i�,q�G�kߒ�^ڶ0?'��jΗ�WF�9£\^�`�݉-\�����5�69�@|O#&�Pܮ`���@ڵ�)�oM7w��n�Go�]N�(��j[��@���g2�n��t��#-ώԳ*x�|���.��3Om�]���iRa��ov:�LȐtE��:3���,���P�N����ts�I��?��׻K�M6'/L�1�WaN�3"��Gs����G.�tE���<7P����W���IN�E��5ŨN?e����e-�S�O�z��$ ��(�ň�ܚ:��Ψ�[��'$�;3��.��8�S�&���PEQ��|����H��A9e��6���B�ICf��m)�p����BD���jI�n��s�T`��vyf9�z�ڒ�w�v�z.7��T^=�����rC�W9�>*�!C��4���M�q�4�ў,�,����򭈗3��� 8<{�O�.��ઁ=Cr���(ˠ�Z��]�u��6����	���J7�V/���T^���p�HƑ��i�]�T�r�N԰�5_UN�M��=u�ڭ����j�ӕ���o]ȩ��l�p�n\�V�Ĩg�\iP���r�x�H��wçL�y*
R�}����i�\�Ϊ~*_9�7*m�4�[G���F_)�R�0�-� �Uy��[)��y]�������s{fk,h�z@�IO�5�M����&or��'6j�v�9V�;�i�9����ܘ���ΕB�ckcuV�7�}Z�t@ə�	鬚��`rm������9Z6k��V�x�bY�Z��w.}X��<������M�P�W�?	��z-��lꮙO����w�b��[qdI���Mk1�Fa}:oTu{b����=?���x�|1�roն���_I�>O݁�A�r���E=ؖ`pӳ�#/'c���8�
w}>���#�Y�����M*䮫&]��#���_h��݉��{��;Z�^��fN����jK��55�N:�T.�����#����}�i�.���d�3A��׽����l5��v�&8���ͣ�f����t%_�o�)̅i쯮��R��V�Y�M}�����=ѳ�/�uBrϗ�ʤ�N��GoG��
Q�3�66q-Ѻ��RJAh+O4�̱��\?v4�L�^�~=Փa�"��d3�w���UyF�����Go�l�w�.���=�֕�=S@���++gb�d5X�!	�rg��r-*��vYċ��[w[vȍ�_��J��Ii6���.��������ۢ�Y�+�V�c�l��R(��Pd��@�d�sNg� ��U2��b�xa�=��T!D��p�|ځTL�A#*�#2۽
�b��'|ܵڋ�ʸm��91��	�n;NKjDs���J�I*{}&i�>M]�ً��� G���q�
Y�`�N���aÜ%ib�\5g�;�,��ߛ,]eGLW�<���9��G ��� �[�[����R���T���Y��v3P=x�*£e��uΨ6�V5g���1G�t=զ��R����'ˌq�IAW�T3P�{�6�oD�U}�h��N !p!~
2�U�6wJJۗ|s{���U��ב3Y�}��p�l�ۯ �{���,l�3Z�]q�wsF������F"d��)��Yϓ��]�������oO���?��P{(�ާ��ɞ>�fM�����+�F�e��,!?�A�x���eQh��%=��*��gMl�4��7r]国4(5C'5����rW�q]Y?���T�����r��";�w*rW&�z	�3��C5�A��|��2y{]�z��9�7��7f!��od.��t�=��ʢAؗ�l�tl�n�7��KN~p��Y~�S�_���z��t9?~��}N���W���Y��%sUp���cT�Z|tQ�c���/�<$�6�lN5@�:��ɩ��U݁֒AD`���i`�3����/HYoO��|��_�W��v>b�%G�%��Uw��Ʉ�B<���{)Wg,RS��@�gk"��(�>�D�Y�q�����kJ��
�RXO@�d�s��;b��ܔF�K!��Tws��$��S���w��^N|"���nj���D�N*W5{7�w6ި|'|g��HHK�
�S��H-��ߧ��fb�+$ֹ}7�b���F���S7�!�JX}|A�QR�#�'�G<Ʃ̮������^d�?QMв0B�r _Z5�|�B��K��='K�Kf���q���ksw!��>駁4�.�s	|6֍)q���B�iM��\�VY�`}�:LU��Ry��* �ċq��!F�w�<�8��yTz�9��zy���1H�n�)6vک�b^���x������3=\���r�|[}�%Q�\l6�+K������a-TUu�ۚ������yalW��u���bUVYtI�J�]�0�R����5�oR���]�����n!�8ݓ�Kz��%Q�6z�jAgq�
�K��[0.���f��Y�r�FK����a�K��'{�x��d�خ}���=>�g����o�>>>>>><������ݻv���ߝg���}ʑ�^:�l���d�CZz�_wd�K(핬n�Y�A�-�h]v��(�讅���a��&�u�#�Ylټ���t��y�|�Gw� j
OUT΄gb�GD��Rʑ[�,ً�E�V��0}E��R��e�Ԭ��u��(�Wε�k.��z��D�=k:�C:�f6�3��z����k.��<^�3�,x6��hNc%<��h��:f�]x*�t�e����5�kF�I�c!��eEY��J��Br�řY���[5�1�;��>	i�{�-7ϫ��p�N�f����g�4*;�Ց�k�Tɍ��Y������N㾷�fF�]ly"�J��\��S�kV��g�F��<�i��Z�U�X���C��}%|\�[}��U�]E�2�لS��<����c��-E�3l)�T�<����Sҍ�J��ٳw��iy�k�1�b�ed���pv�N�7�JC�)����&Pws��%�]�m��PSa��Ěm�P�Z���eh�Z6�v3��%�Iշ�NE�t*�Z�KY��	�Y:\Yh�*�:�L��ͅ��H8L�vI��\T'�bo��ɧa�7;v�.�v��f�ܮ�iB1��oi.��{Ev ����
��%+��J�n���hdڼ�"�=��u�+OOi4��6jx7�6���� �k�{�����T�A�xȆ�;�{�䮊�v��N��h��J*�:�:�$2�^b��4���\7!oP��{�st��hj���p';s̘6h�j�`�c�Wy����47o�i�D׏�6�L�*�^Adpʹ��e�F0ܥ�N��b��:������eK�ۢ~v��࿻+]�1V��ݵG^9ȝ�Uۚ19е�R�&2f>
J�6E�ŉ���i�_�����{�vڑ�c�EbN��Y�FVZwJ��Rf�2ͮ�'!�uhe��kZ)�E㢊��l�.������ͮ�����6K�U��FX��ݹW��%��Q�6�)��v:Q^�p�'چ�Q��6|ފR�Z.p�:�Y���y��;;58d�����5E%�V�v1����x�zIg��T���w��yΞ��`�ok�Vk�}u&�ǂ���"�*�`E�њ	�]�y "��6N�5r��;�sB{+�/wN��h��5���ʁ��NՌ����1&Z�Ei�\�6����u7i�}�t+h�8�ۛ	���Ħ{)�{P9�T�+)���Ĩve��QSΛ:J��-W�����p�ʚ�^���������g.��x�3Ӂ���jZx
�۩\5�G_]���S�`�[KB�����z���T�&eQ,�vձ��)��uҽ����l�'x��[��%r��;���'ԩ���Y�]l9�t�;��bI�|u�=w��� �*�J��hi�j��*��
i��hbih
(�E�ӘaPQUAE%D��R5��AH�CKCCUPU�%4�%EIESIABRT�!P�UMQ	T�\��-QT�RRU$HRPRD�4k ��h��"J)(h����� �
F��ih����^' ���)�(�)�&�h"�����������(�j+$2P���������&� ���J
hfh��"��"��f*�a��������hh
H����j�)���0r��jj��!)h
�����J��(�� ���)��h(������� �)���3��*�$���"!��(�
��VTEJ��4�QEKHRIE��(X�̖����Ji,�ʛ1&������|��|�W���޸f`H���'N��[���ܧ�}.�u�a�Y��m�ͺ�J�И��}���.�t5z5�u�;����[�*�;غ{���6z��|�9����(�@u��ܬ�����c楙z��k��ζ�z3��;V6�!�q�|�c�3j�4�`��9;M����ty�c�q}ʁ2D�c�1���s#M���� e��]]4�Z�[Ƿ�c�7��#���J�;�@H�r?{�D��<�:˟�����F�Ig��}w�Υ
#�Yj�{5u׻��Hy�q��*"|4�k�D��Z�Eu�I�Κ{��!�2Dow&�K��\\�+laA8n�L#^VJc][�:K���ݯ[y��ԋ�u>�b*Ea�8N,J�dJ��溟u=g�#3Q�-U�������Ϫ�u�L6���E�qέ�
�����Ga� ���O%JR��r6�G���u�{CU?[�L�a�w��w7�D�&��l�V�T�I$���R���^v�sp�m�	X���"~�{r��~f�Lo�"߮��.�~�̤6���db��������9.��Z�s��뙱~�\]�qUh2*̕]���^�r� �]�UY]$λ���U5�8�+<Z{O9幅�is�2Y��7`R(+��-�{	M�4�%�8,����l�k���ݞJ�	\~n�!gjk{�M��3ݍ�k�^`�M�S�A�>����l��kc�z�F�O\�����M�R���9..��fv=j�;@mo0�� ?�>AU��G�nL�o,N��R~{�x)�Ra ��'w|mt�i����gC{����6uT�\<ٷ��mn<.�3���.K8$MMyT�U�O�7�G �qw]T�q-&����E��go]X�U
��q�d�o5�;�v�1�hX����<�M�'��+A���LH��9� d���M�b=^/7dIm��n��5��~*�����;�����Ty�٭�J���첽JBBAR���}�9���6^��M�R�?H�g��L�a��B:�����b)?eV���sP��W�+� Z�V��ܖ{*j�jg������x�7}u?Vh����)ht�'�K��yb��Q�I4���i��V��Tv^��S��^�A��3ٚ�,$*u��J�}�@����h�w�%��Y��I������(�r�f��u�b]���T3[��'[����pf�!��R���7�ȹ/�T*�0�~���ݶ�j��Ԩ��$e-	i͵"�l��7aM2!�����c�-ף�.�eB�5;�,�PT��'�P�&���v�2y���ȅͻ�!3s�4�p�j|��:Hʡ
�o�f�����0n�f�ꭹP�3�[�T�q���t��#R���\���197��1�v�5חs�$�\zv��}�� ��\!�,�՞���Io�1%��`�F�f��h����rF�.�pϛ1�m��B؂�v	#��^5�5��q/�g���s���1�IM�rug>Ol����1�As�խ�p�,U��M'k����3�o��Ď���]ڱ�����\yآ�.�:�u�s1fr�U,�����=Ф�'*�����w��3"�i��5]v�LB'�z�'�}�ւX.<#�$
�6�ˋ]�?-K�yN�����ks���S(U޻���ڦZ6��m�on�a�}tE�mMc˭�4�r8�VC�T�m�_XB�?���]	C*)�}�yK�q�jպo���v�8�=��g�k#�;Cl�.oEn�����Y�X8���i�ʖ��tٷ1���"���w��* $1zé�y�� �y�[!l�8�q}��[.*un2zA-����l�;���gE~ɕ`p���)���v��7;�ֈʗ��i~��cL6��b��h@�vI,tI��1� b�	4>�We<5FU�.�{]�ۤqY���<H�����9m�zs�X0�ڣ5�*�޽�����8�77���H�� �T��²V�ul:N�1���!*6�]��p�(��^���2b�jKo�=EJ(�)u��٫wbcvmwu]�H�f`�
���֙�u��
�E�E�v���t	Gnt�z� �>\��c����������U�ْ:i�M3�B�.}	���K�|��3qbu�:6�7&ȭD�c��\�k��ܷSِ$[����%���
��ٿ���ʘ�X��.I��C�ҵ#r�Z*\߳���<���ٌxE�b�5	���a�����9��������dm��J[0��Z�С������!͛�
��Np�����AҺYI�KZX�3:�ǧ�����c���c-�en̳��u��foa �Knk��fr}>�\MF�f]0c��)#^�s�(S��þ��^�MrV��y\m�)Z_K��*	��wH��������I�����(~�.���:��{����]+�h%�>�W���8�DdNp���0 ��a�v@u��6e*�2,�U{�rY�g�bS^�Ȟ�RFL�:B�e���f�l0K�;V��T�`/5�K�p�"��5�����;ԯʺ<z��St�m�oPq��Wd;l�ú�}ų]���u�K��R��9^==ѳ�p�6�`����F=G��z�e;o�g�*w��t?$fDL��%�v
�4�:I6��B6t�(����$��ԏ8��ތ�&�p��k��9	o8&��en���p�滋x{>��5煨��[sۗ�1������'���.��5�vm&��^����@!(��ɩ���ȹ��V�o�����?������AW,w52�$�n��T�-�.��7N\63�v7y���:K� M��Vy]����w��Wf����X��\f˪��'QE�����Y�$����Sz����snjԇwLgT\!9v;�ʑॏ�֊���9W�:��-�77zP���R-��F+�ohWu��,������B�*�1�FHS9ŕ�&�c_Ѡ�S�k����^ґ�at#s�s�s5l��M���+U\ܬ]o�Ϯ�DZ�"}xz|�B�к�<�)U>�첱4��S뗐�&����ݰ� �ȅ���F����l�I\�|�ܠ���01�ߓ��k��:�S�hl���t-vy+F�C�T���"{����n.8��{#��~��]��H�[;�&��畓��ݕz�BMt���:f�s�)rx�g��Wy`�ǟ ����:�'��S�b�9�f�����hۉ'v|mq��Ά���z_#���^�l�����/�_w[�H�d9�U��m����T�E��O�7�Ctw]�����Xw�����8�����5��o6�Q���;b:Cl�����w$n��ʑ�B����'X����@�ժ�*�(/WqÖ���/�:��e��Lu����f�>OH�{,�:u��1�����L���^�]����8�p�~|�]/9wU��*I�.��M,�g2j�u��kW]�^�_;m���錢čgCF����V+�Ъ���f6ۊ�re�Yiՙ!d���G�tg��d�ƍQֽ�p/؊�����ˇ}x��F���
��{�ѱ�� <�$?2��-Xij�i��Ū.E�m�t�fͺ�j�!�!F�UyF�cZ#5T����X0���}�WRV�"���Z���������^�&��k�e�o���c��}y�̓��y����jHO��2M%^H�Nm��e������u��ND�F�[|{7�iTȍ�U��Ԃ��(*Np֨�d�朡W�^=���Ohv���9��d���{�+�Fp�:�\-�ځD�<2�)c3�P"��g����܈�)[�V�w�r%�7�v.�6�G9&��r�+v�bs�.��V��뎺s>����� �+M�7���OPfl�/"Z!]'���h������2<���-��6� �ǜ���O���o�!���!�:r.��Ѧ�_�Ǜ�o<��{��{Ď�i��r��L�V�qۻ�]�J���ՁcY���!�+1~�<�����FfW��+��m.�x�f���z���ۃ�kA>b�t�Vn'��_)�du{���J��,0�=})�9�)&����ҽ�����ei�9 �xc-�"��?{)�Yљ{Ãf�f���ٽ�I�Sᳳ�;�Z��IOx��X�a�mg�eS��.��qs❬�y��9ӱ�Ҩ�rr��>>Y�f��5#;�l+{�y6�u����ü��Tǜd���4��]@ՔOuE�I�D�+X�Bb�f_�{�1�@[a�zw�H~�v��; �3.�}��"^�Ae�ߧ�߽q;3���C>�g��3��Ib�j�]���u�ы7[M@�I�h���A%��;��]� ��=�v��Z�g�s�w�i�R�N�}�R��I_9?A�(/�����������w��k�9��NA������W��y|H� �T���Ee-�z��X�" ������3*��q�P�U=g��_�:����+}��QX����U�g��˶��A���Q*�eV<��u�6��l� �.�-J�E��)P&�oF���I�U�6v����m7�_.�ia]7��\�5��Y���gK�I'[�՚v�#lv����mR^�t6R��6mD��nmU��m93����{�����烿V��.����ӽ�ao��)��c�n�Y�t���Tz�:i�M2�("�!`�C��;�ϲe̩͞v��!������s	�|�9���\�-�@!y��ŝ\Ofѷ���o��ͯ@���L{�
6ܑV�)"t6��w_�-�v��?��\�%I��hB��� �mI�|Z=�%Q�\l6�>Z_g�M���O��Cr�<|���$'���t��!�0�Y��پJ�Ӌ�ܥ�~��|e��h�=�I�d�Dwm~WC���a�}[��*��q���-MoJ��5�H��W����{,2�HC6p�#;Wi�\��n�y��#O;WuuY'	P=Cg�M��Dx9���}oT�y\��#�9�����V�H�Zm�tl��4� ǈ`8�7��Ď�g�t-MH�Y*+������f��R�Ũ���C��K���������mt�	"'�h��u:Y��bR�*U�&9��m�U���|h�q-{���).�����{�T�H�I�V��*�u�/J���*���M��8��������]��$��˱�=�M������\�$H��	{��}�ܑ�ИX��k2��;xos�%�A�x4�F]{�ٖ����#�"}Ĳ�!���t�}[�sMe��v�$��$bg�b "�Uy,���u��f_�B���W�����\���i�7SH����x��W��ty��O��T���	��?�o<�8scW������#��}J�]Q��yޥC*�є:��B�
	C�!�y�
��E�wb�{͞�#�H7^�IU�*�#r��M9�U��i�f���5h�V?l�ݑ��w3���.������y%	Kd��i���5\��9W���Y��pW�?+�b#o��JJ��	-�Or$�?-Ys
J΃5ُ0:^η�Q�䶄�Q��+�>��X�"��ۖh[ww��uٛՏ3Yם|@=|��0�Hn&5l�t�:߻��oo�n�oo�n������������������ɯ�8���ؾ���3ڦr���:&���&�u���<�k�bQf��yc��bÉ�B�4PC/�����{\s'�.@hWjis;z���1���E�.1۪�@�+HX��j�*��F�:����'!���u��է9kJ��ڲ��%���,1#���xD���O�����2w.b��њ��\�[Y��7%�塗��b�v��:��Nbv:4��Bw[������噜��J�D��tQ��"�S.��1�RΚ�\b
��4�����<��r���r�w$�i9z5H.ׄ�Uϸ�:�"�X�0�Φ2��)��)��,�Q�81�j�2��<�]��!��W]��>f��8���`���:ÄL �j����fu��;���K]�ِv�!�7Mh�"JS�+f�u�K;)i�+���}}���j�{�9���M�f��LYC�B��.t3Q�G����=N[��׼��w]`Q(K�]b�a]#�XN�Ò�h���/�E���9�7��(��K�I�o�x���ȫ���h�v��j�
�k�e�"�rS֕#�h�Gb����9��JC{��/k�� ��T,\_C6�j�v�X��YX�w�k��#�j%<(l9�l��㽚&��:�j��k!���;�@����!��t�mE���@�u�t���cª(��S�%���a��<A��4�g�{�,�Aow�h;[EbN�ݤѴ�-ś|s4i%om�w�&^<�M؂��f�G�\���٦�k��_ҕ�m]�rA\J�Ż��i=n����Q�y��uu��\g/0�:��0�8:�Ov��aX˷�z�H�ju٠�G����v��t��v�r�A�T�����w_2)gʸ<o���,�вِlnu�7b�
g�(hr�5�Цց��b�ٴZ��fлA�̬�u�چ�Ü�O,���˨��<3l�΋MIM��t�q�F�0f;��Dϰ�mNwK32���kD�v�����b%f�Բvإ+ꝦCL�Z��,�� �Q�vM�t�aӥx��=�w�he魸�u��)hY�r�uY]k6R�����Π�hj��NC���۽�T�KAidN{°R��7 ���0>4�?�%҅[��V[�n����aY`��@�������~�����w�v�.� �a�9�-˽m��ol��,���L�J��˺��6rbӅw\�lr��$����+UY/���曮[�#Zf�mok#$ZC�GLM<�[�J�ռ�Q�rw�o�k��5��]A�/Z�uu]����M��c��r��s�r�5��V����.	ݦ�ɹގ���
�KỤ̃4���;�J���ܸ��i������K��p�՛��L�k9>I�쪈n������3�,�F��:.-����C+C]�[R=�GrU�۬5>꒗k��/;:M6���*X�:�M��J#BD.8�����Ե��UZMSlF�L:$�F��4�γZl�Z�y�s���JJ�(���p�������()J(J((
i!�Ȃ�)���*��)(�����)�)"�"JR����((�I������Z(���)ih��� R�%�q0�PSH��U	AA@D4B����PP�a�R��J�č9&ATR�- SIT�M4�Д�UT$@%4�D���(Z)J�j�
ZJ��Ԙ�KIB�4RR��DP��#CХ�J�� ���)I��!J��*�J�(�Z(���RP�S��{��6zֵ�n{���ל]�Ta���S�;�D�b̬,���]���z/��Ig:���og�e��E��1��V�4({��h��I�:t��4i'/��v�k����{��}��%r~Ќ����
ot �d?��m���
�q��&��%--�Q�W�	��k�Qan l���z(�v�O�:k���}���k���>��46g���@�[IS^T��r2���}����d������cj�PR6F���Z��>��:K���bj�4^@i֨j��OYs�S!����0l�2��-����3�;���hf��?�4��~�
��SϮ��L	�<+46q*��������M[T�n槼�t����`�1���߶��h�nItu���ՠ��h�{����33��a���h��(:-��#b�ϲY�c�	���3�{4n����ZDʜ�;e{Jla"=��@��5��f��t�6Z\3�6`jٸ۶��y��3����+b�'Q	�҃$�Zpz��}~�DyG\�3z��)�K?O�U0/lv6��f郸�ǣzk�N깖�0�TE�H�|[��w~�̀�A�j*�שXs�W;*X��u�VV�w�`u���A[|;��;��>��[7�oIZC���Tv!7+�N8��f����EH:iDAh�Ȫ�����y���x7����B�U:��L"�@̣���q�]�����̎7�s��υ[?��ȩ�V�p�ž���fb-u}���Ӊ[�71��}�WW�IU �}r�N�"�!O�FSjJ��a0^՜�ٴ{^����E'�1$�m�O.=}���?��p��AP.���Դ����؉�lqg��ռٶ��hb\C32偕ǖs��]������瓌�:����yc���
���힞�v:���}gɔ�]ڱ�0q;8�s7���ӷ]V���y�$��y��\dlΪ�4X���JU��ѥS�>q��t��e�oe�A�`�ϣTł�c��F�NJ�/�KX��͹yg;!�CUj��ݲ2��m�H�0!t�F�B�ó��}�8xY��OC_Wvi�T"���4sl����<�C���N:��w�1�p]�~�1 �=��d��u��2�_QlQ%�Wd��0��+�Z��Q�Q���}Ֆ��3^��P ̺��� �Z}}4tN�moTs@��i�U ڒIؘ�@����-����,��XHN��7�D��2��Ĳ���Z�)H���Oj�S�2a�v8Op�$��tQ���2�0�v�ߊ�]�=�3���^�e��x� Di�崗��:��xg��]91Ҩ�H=\w��`����
 =�'�����h��/���R�r���$��Dؗz����}�Of���k�ꧪf�VLT�R[^����0�\��gMT��ry�+m��s��Ya�s�gV4��:���#�գQ�����U����c��׬"��a�=G����T@9�=4�Xo�$ Jt.�P�Գuۣ��Y����E��$l1��"��5A��[���>o�gic�����c[���n���+nZcv7���Eg��HJ�Hڛ�U9��!��ŕ��k����95��E����jU���*��\oͩ-/��b�y���zj�7I��y�^k,*B9a��]��P�J�.�R��}ι�;&�m��K�K7LJfɒ�8I�',҇8w{bèf���zz���N��w�H�v2��'���Z���0�����*�K�f��^��YŦ����WGs2�_e��#���l���9+��s��O(j�N��flf��)R�o��h�N�jtU����U����q��xs������2U�g�r���zU�f������Nw$W4�����=��=�����l�+�;U*�0Z��V�
53xLu�U�1����䓧(��V����VΨ�bG�ͭ�����`�̣�Iucd�P,��)Qԍ�9G�$���i�^6��������\y�aj������v-�J^x6�$lك#�mq�d���$�yP3&�#���\Ú�<6�C�0�'`���xT_+�wM��5w
�O6��Oiv�8�{�l}6*=�訉��B�Y������u�܌�Cٕ�/�2V~2&��k�?r$��K?�g^�H��A({�1��,*UB3��9���-W�=��,�U*3�I�Ưf⛚u=,�)�A�M8æ�o��.3l.�j$!G4ף"i
�wܒ�0�B7 �܁SNdƯW��A�wS*����LE��+0fiUK(�)��=�$\�݁3k�=Z�T�\z��'��*li΢�W�Gs�6�?/�K@�an%�>��,��r>�ᣖG��h\z)����b�cK�ᡎm�NF����k�	`��U��h��p�ȳN�G�:�&�!��Wln���w����G���
���~�����]�nAH=��J�R�S�^�S1�N�.�Y��:kn]�i�>�'�Ȃ��ۆ��|�[J��{�ب;Ľ���v�d��J@>^ש�ߧ���
��V����W���ըܪ��gCEl�ag{;{k{̛c�)�A�P~[����R������)'\���c<LH&��	 .O�Ł��+���\�W��/��H��6?k~4��hӋEr��(¼1�'vA��XV�!�N���Bשa���D��K�1�]�2����Ua��ɻ�Q�Sc�E����01[�5J�oSd��Qy��Cdnnt�V�>�Q�Lv<��vU�y婩�.��
���u@���S��[h��d���؏q~�Xݦ!OlnS=K�l��\)�Aޅ#�Y�������³[8�n� ��#\��ޙlC|����u���[�Eܬ��CW*��f�H��':0��k���G^��)�d��R9��yZ��Y;h]O.Ǆ�(2v(2S\}�3V�oj��pFM{�����W�c���|��x���UcҖ�v7O��z˒,�mP���qK�S���ݪ��ކޝ��Y<$�i��2*)�}��������K�d69���۵=ӽ���u�緑*��ȴW{mP��`��S������r_�>��^�dʓ��sȡ"� �I#mӌᵑl���6ͽ�'^r���]����$���^�.2G���()�(2OZ���X+�E���Mnw����
a����иj�N�CjP&Q�Z�պ�п\'Y��t���;���~�O�AEH�nػ+]Z�Wo���(���Z�=k�����U*	%T�p:�ԁ�N�������D�n᣽���3�̊V�
���Ķɐ	��l\#u��B�Ꞙ�ǭMX�v��³�xFw��&߬
���*j	u�-�u��h��ɯ�C�i�z���<�1'[����==]�g�kbz�S^	wH��,چ(�k(;���a�K۶3��N���7�V�[~���4�Z5e���.��xخA�6��=�F�gQ=�jH�e�N��'ڳv���)�:�+f�f��t1��+⃊�o��c{k.(���xWX�����>]mWKL>���嚍�G�*Bw2��~o��#@s��;��I�A�ʮ��^��D-���ͭ���6kR��Ӵ�=f��	��7RbW�(�U�kB��A��O���"�Ӭlo��{��~�kd-����qpb&{25	��4x� �ʢA�&:Nٞ�ǝ�h�|
Ӫ�������H��X}���,�~��d��D��Sa�0���;�v�:k2*���Փ{�=�d<�$IDG��G-�P������h6���1G,�7�}�����v��E��p��ܑ?����>*��M�i-|1���=����Z�ٴ&gH�o���,*	S�OP����:�Ѱ��u�kp��{�фiK�l��(�z�]H��W�w��Ʈ�F�lNut5��cïNG���<fO�i�i�=^PE�_��5�i�m�g�:������W�t��/���:I�V3o��9�׳���p^^���Vϓ�L�:w� �Ӧ���F�J"@���S��7c�k;��:�IAc��!Û�E(�����rA;3-�Զ�Y�/Q�uR.���4��{tr�*,��^IL�}����{ҕ�EH0MS�)��GfH��ϒ=F��ʢ�la�S�t�B�F�$G$���J��-���q��;�!�'�Y����ޮ��p# :="��2����(�.%�*8�;�v.�b���~C2v|�0��q�.�]�c�{�.���b��;����2�ܾZI�d���C��dy���V��b��T�:p�|�a���I��nγ�wĪY�f���7�8	`�l�֏0�
�M1�����fn��k�Y���^t�B�Y@��J{@=Cz[�|�G4�0׽CZ"S��x{��*h[�m���D��E7E�FH�p��(�t�D���m�q���NS�*�82�q&�H+~��ԎfgKX�5�����W뵿<��$
}���ጧ�$#DG�H7ýޞQ�'gS���`��2�n���vB�Y��cx��`op�Jk���E)�.�*�t�����5	Fl�ݠ�U[+ ��b·*�XfD�+�F��*��I�(��R��V�.懭��v�jY�]-��O��74v��7���b���0(/4�Y�V���|n9�����w�g�P��K��a ,�zJ}�⮺F�5��?��M����r��3������?D�/mH觍�zЂMw�/��9��΍Ñy�da��Qҗ^�
��K�|���	&���g����i�=���r�{w�iu'ι�rx{ڂ����:?2{6���~�~1�F�_��s�c�#�ܾ�V"�t� �����Wr�w�
7*�%U.M��Dd�\w�#0J=��F��t��(�7�������9�f*����]�t�i�v�+g��u������Vմ��5�@����h��/�mҤ,��},[a�:8n&5n�9���p��.hi���'8�0��(=�*��~r��Ǹ�~�f:=���{�6���*d�K_Yk{7f����Y4��w.�7�	��k��m������p�A�ך�%��]�r�1���e�i6��\+����)��uY R	ZF�]L��P�=�\fpk;Pj2�ahx��6T+��!�]_	{(V(��w����i�ܲߺ�v̓G^�n�n�W9.�C2$��u��ժf.��d���B���2��3;[��R�Y<�pH��7��"�<ˬ�n�h�#U\Bx@�����o�#ss�k��φ�w)��l���<��U[����2v���X���j���F홌e�[�����c�!���x��s������|��!��d;�`F��J����0V��vfj�z���Q)�R"A ƞh�Qח��;�\��cww�y��m2ڍk�l��qwD<��4V��-����s#%��1��1��E��/h
rE��ۙI�z��)f��U�6m!�J;��]�'��w\��w���П3�0%�%�!�����:���<��R�I��=��o.*M�1wۺ��cݡ����OP(G[��w��m@�Sq͔]K��x�w�����;=Psƨ�d�o[)�g��'"��q��z6N�O�۷����������������{��^طX%OnAQJZ��wcm��D�c��v��l��8�����o���R��_�.ən�K+����h�W4�}�w'�w6<�lu�d�¯2��N���>ڳ'���J=�o{M�E�5ۦ���\4^�������w���_�,�-��	MC�3����/n�(��z���<6�^�]B��* �Y�Kma˭�"%��LL��Wi��f��Uea��c���Ү�8n�w�32��:B,��5�M�-�/BH�ÑP����tfa��v7��Z� ��;fWԼu���<J�7��u:T�3�\����.ť�WY���
��7v4��V��K��Ф���h�y�T�G��	��t6��[{��m͑pǪ�V�b�|�o�6��-�/��-�l��\��x�.�6�+3w!W�儦I���'M�z 23�,�.2�]����������[�iZ��=��@0���)훲��_ ��a
S�g���.�'�nv�f�t\HۃQ٤�%R�%j�W2>�MQ�����w!�ݫ
R+�T�Wp��4qS�+N�j�J:�s��8�Q�S&���T�{�/7��j�í�OP��Z��K�7Wy����B��m�j�!�v��)ꦠ;%�hB��nvI2��|�ʝ�FH���c(`����U��:�8g����{f��'�_�ʎNŸ��f��#J��IfV�@BF�ղj�f�S:��X��`h��A� +��Z�*��������׏R{G���'�tR®[+���N__qbj�}09�N�&���W��}�EGfPAS���ޕČ�up�r�s+��65ѽ�Ɨ�nZQe�87T���Vfz�)���Z7&���`�Ysx��f8e(vV�	���&|2(��O��7$TV��(�n��z�t��'/�dLVe�)V��&��c��/n�M�fZ#�f�{�a���.��k�'t����շ��w����䛼ȼ5�"������CH^�͖M��/�ͻ��}Nsf��w�kz���1��hgb6^Fq��p�S���wV����ح���̽$��
q,W_�e��}+M,�u�n�voQ��B�W�E[��
����]]�Nv{��}�f�H6m.��i�7e2�t�n�[�Nt�S��A�h�:���h�B�B��.�h��Y�Qh6�����U.��HEZ�v���F��*��nK�i����-IUo�,mcH����w�=\��װ��|s�R.�̛�٥�i��������aH*L���F���cy�@�$��&2s9�3��Ԅ已��v=4���XΥ�Y!����,���<|��ܜSm�\�]SzF֋̱&01⡥96��X5�a(f��#r[n����v�M9஦�R֞z��YI��6RrS.j��;��<��<y����Z�ij���(h�!���* ��
JF�� ����B�3&J�%

(X�b�R�)"8�V��(L�$(h5�U#TP�P�rh��JP���j���9-4TPP�AAB�PP4�9j5jF�2JA� �*��D�C	�JL�Z�()
uB� ��@�5MP��k��P�C�'�
R�9.B�)�P�d%&I�9':�P��ŕE%�2�2�"��۬�z������Q㷛��#9Z+I}�WCm��l�1'�A�N������{��V���{�_]�����3���2�f��+����u�gW�bN�&���A$���Ǉ]:�.6X1.�����ryD�Ƥ��af���zZ;��~n\h6ɐO.�N��6�_��8�[::��1�v"n�p`��[>�;m͊���d�&Q@�{]���E{q&Kh��l���7�7X�V*em����3ֶ'�%4�uV35��
Z���mj�Ơ�ݐ�o��� p����#fuP�4X���ϲ�mQ�۲3i��wfI!��vvV̋^�`�|�oE�ǿ{fš�w�:lܹd�;!�W���w"�:YH�U;��w�7�8.��1Q�+�)l��p�#�l�o�_eP$�c}�eOPc�9���N͵%>TV^���v04m��+� ������d��tQ�b����������r�r�v�
!��|�S�G=�`fY �"AN4�g��󔝍϶�4[�� �.t{���*U��q�t)]);,��K����\ V���Gx��΍a,����E�2�I�r;��Rj1C2WZ�
�޼G�m�,]D�9ɚ�J��v�b�J���,2*Ļa���i�_wqw^B�őo���c�%0f0�hצj��`ff�� h(,��fCd�*��4l�z�h����F��B�k�J�OW�͞���i�vZ��`�޷Vp�f���E�OA"����D��L�yd��&�*s]CC�1�g�;��:y98� ��xQ�.yN�-��駁4�<�՚�Y��g����H��z/l�z|��6�T�R�j��)ܷC:��^zٮ}G6F���z��Ho�H\�m�=��7aJ/��>��"]�A���Y����9�f�-� !�:������l�*������Q�\[-����k�hl�'��d��+Z���OKvAYa�.u�:��bR���WR&�����"�����'���|���q�k�Y}[ճ%)Qt};ڮ���s�=�� x򠳸�*ݟކ2�9��޿?'��Z�5����,�C7bʽ#jT�5�E]�H��>�ؑ��oS`���H��Zs3�u�4���r��U�j<���)�k�.��xEr�/��S�s�e��w�6�e8�(��8�� �/ov"�/d5ߢ��n�m�)p-7]���G��B��P�4Zsy{�}�'�r�ٺ�ҧU*�J�Y^'���;#;��|ɹE�I�ok�gw7lm�L�­��q��}�Hד�������7�/�q;L��"j�ޮ^�GpU��D�b~��e�������&H$�L��U�9����M�^��b�F+~�t1tY��E��I���-��P� �~�y�������A%�Z��9́yB���S�����r�5��/�.�;�~,�y�"����������M~W��7��:��4��0R���g^�)9�w�-�������Y���AJ�]M���%��i���O�D���92����(���dd*��Z2�Ќa۹����j#���j5"]����~��V��9��?�xi��܂ �'QC3;0��a5-�����wr�x�ʹ�n�����#$Ey#��:��BI�~U+8y����#)�7.a�0O�ά��	"�/���@d�؉1׀�*Ic$��Y��71��}�;�[��h,d�{��wjǗ��o��]�z��p�z���|:��/��\��2�M��w�㞱����Ww)�8f�%.+	t�^���՜���ݟq'�������tV��l0�cs�1�ݲ�Q��h�*�'�Xn�!gouv ŷ�!�,:�g���k�٭�^gH���J�i4x�ؑ�GRD�.O�����aty��m�˸|U�����卵��>GnĮ�յ@�b@W�'�wd��4�#X3ƈ�Юʚ'OT�s1�y9C��1����*C�Y�y-��55�V�{L��>�j�9�}{�"b��F��qXb7����ԩ��l4"n��~�nԱ�.�"���
'�?���ӄ��_������A `>٘�Y;��6�2��'@�=�ߜ��(�q?�G��Kw�~����vt+�`F�ya�9�i��tk`�l���ݮ�����e���K�$�y��Q��OӐ�vA�Q���5Yok���;��լ��������wD<��5�	�"�+)k˜�yj��3�W;dZ�j����j�m�s���Ul���,�1y��?#�=ӱU*55��ν����R��աި&a�M�x�P*�*��y)�r�z3��z���ˮ�ޠ�D4Z`�[����ܜ�:t�PT��8���	���Zs�d�;WC�"@�v�pfŕ�@�p����͕�#RBk�2AaIPH�;.b��^����ɽgú� ����D�E�������~ff���PRֻ)�LA��Ǽ�g$�n�����T^M�:�A���#�`��5j��f�6�d��k�,�4�y��V�佥�t$eP�f|v�F�uV���
v@��d�1]��)�>L��Γ��_]?K�o8~��>��1�JW)R��UA���u:\@"�eT��h���L�C>��[��y�� ��]7���%�ˍtGD�pyepσf<yu�<�S0��VyFM^A�
�2�@���ۅ"�4m�����-՜���ܿS;�g0��&y�kj�~a�ސ"�tv�3ֶ:�R^�u/1ks1*㻉��]|�Y�[U��2�{3���X4��G8��v%.EEL��7p�"s��-��� ��m0|��F�8(�vO��
g+kdY��!	�a8^��Cq�lL8]�WU,ɿ*C^#TΚ��b�P֞ʕ��H2� ]�s,�X���8�\,�^QW��miFkimK\4�X/�@���­Z��X�,;��u�ݎ
��{[����7���T�ߪ��ޱ��;gOQ��̞���:�/�+��U;��N�m��a�a�����%4u��Uk�W�G)��['��S��d��l�Pc��;�kPg2��oj��Ȱ��"���F�w";�A�2G�㠒�tQ������Q���}zxmM�/b,�ED�<r�>գctǐ���)	��F�E
�����';��2�si�Ur�3��(���G�]fVZ$u]V��l1��I�{�j騛ч�k��p��"�̍V�zYł�P�S�zp{�OM]W�)ٽ��2ՙ�F�B�X
*U�1ꗇ9��WV �:���;=��;6���U��ÈU�J5w7�3��p�l޼ޯ\#�m�\y!�%F�E�R��dh�p6��.�$T�&�ϔ��!��zn���Y֧6���(�@$��!G��Dm�n�F�rIXn���UC�,��}M|�l3k��kۉ��UAץ���9��خ�}�Ud����}Ty{}O�b�ga�ǋYۙ���zH�ih�j�J��b�Ph�0Ѥ����t�s��;W]wG���>�{(�IK�6ީ�Go��/h;`��U���M��g�n��Qv�ۘ�d^\���(���I�Zhj��n��A���nx<fU���(�&��[�ng�3����w0���:_OG`a��P+/��s���g�3]��ָ[ZOS�ٝ�k*����J��b,�C����`��oe��W��r���\����}{�3��Oo~����a��H��Ⱦ����Y�����,,�ƥ���J����VQ=Ԕ�������ɑ�f�oʹ��evwSew��G�@[>�2��)O�g��wF������ə����=�2���c�?�#x���	f�V�4L��H�ﵛJ+'{�L	��3t�U��� _E�
�Ef"�v�M�XM��c���;�@��܈�%�����O�����B�=%^m�*%��c��<��2r���*G,�@�b!�o*#O&��RE<l3�����6�����L�u��R8�5C'tk峐Y��Z��^��^���v��n�l�t,���B���દ��>�
Cs\t�?�᫆�%i�d�>ʈ�\6���SR�"J��9��9����{o'wb��ۖ�і��Y;���l{�S[�.ٜ^�m�;8Aƫ��sNT�C$���rⰔ�����$��ϗ���4��&˚,�'�ыxT��h�k�8O��U�ȁ�B��*���ʫ�ɻ������ͭ���S[��޿�h��5����V!|�]��
��]��[k����>�v��w�/�Ms��|^�͢0C�"2@�%�b#o��g�Ĩ݀�h�(k���0z��H$�A��@k�S�pEHtV���"�.M��m+���/�d��������J�#H�n�+;dw_K��H!�6�Mcj>�'��ǩ�g���B+s�貛}>8�$Y��%r~�g���\<�Em�+����ѵ�raF|��ٟWu��mQ(ąxbx��6�{��U>^��L��v����8�g� 0*<��O�l�tʟ?u���H��y�]{��b�Ɲ:l�ټ�y8��*�0@ߠ
��F����Z��/��S-66����C��:���o�y;5�a�%�c%�>֫N�Fӊ+�c�V�n10���F��>|��@RS��V����ͬm /b��:�]qn�[�aC���Wm2��sCv�FEt�ۖ��Rw/B�w�T��ԥI���.����5�7�߷h � t���g9�����e���2�U>�wB�Ɯ�{�_����2$o�c�t�)���$�?x���Y�klM_��O"?\�5_M^:��a������H:y�v
26)���i�k�ekGWh�5�A�!�U.�MG^Q�]�=�MhO��YI�_Yq�x��s^`�8[Yh޲y�㙙�D�FY�lp4�H�==@nEΤ�r�Gb[�<�h��%z?Y*7ƽ�������d~\G�Y;��B.3Q
�rw0�U'f���6K����o6i���G�.%��`���s��uRU�^�]��pI�0ٛ��j\��$i:������H�g�SP�.�0��c=�Q=�i���ʐ�b nQ�7A4J�A$����7�֖��[�*���_vUgoL�n�Ȁ�le2R/y��%�ˈ�o'�s�@�{!>���..E���U�S���V�7������Y�}P�ؠt�?^�Ǌ������!g�8C�k�V�ڒ(�NtPgȐ`�>�����_I0g����4z
�Y�z��C�ނ���F���f«Z�`w����p���Y52��lm�.ے�i��KZ��S�����?O���d���jh�:X*�4�[-eW�p�1횼��ɸ~#d��>~�0�+�#z}���l��8<.{:��>һ�	��G,�KC�i�p�iQEz�>4x�mp�o�S�3�:���2�M@�ªj���n��x��zhPj�N�X1�8ު��qt��j7S�RxGW�ٛ�:��P/�;��_��n�;A�7�7�CM܄�[��n�;�=�MrRڭ���i��7�/�J�A�_��E�3��A�������Ƃ`�����D���g�ڹE+�t�dњ�{���LnU�%2�u�Q�Y&���˛�)��#%�hQE���ڴlәd>$d�c�dap!���=94�hV�P�F9�3�w�����ѩ���� 	�/�_�<��x�l���x���M4tVA�6�D5�H%��g߻���_��~㿇� �
��TD_�y@�@D_��C�SѬ�pe�fE�eY�f�VdY�a�f�dY�fQ� � �F`X`Y�f�e�fU�FdY�a�fQ�eY�fU�e�f��eY�	�f�Fe�fQ�� �eY�f�`Y�f�E�Fe`Y�fE�`Y�fE�E�FeY�	�f�`Y�f�� �`Y�fU�FdY�	�a�fE�V`Y�f�V`Y�f '�yD�	�fQ�dY�f�dY�	�f�f�dY�f�aY�f��paY�f�V`Y�f�a�dY�fE�V`Y�f &�F`&E� �V`Y�fD�C`Y�f &D�aY�fE�Fd�f�^YdY�f�dL$�A�d�fE�`�f�F`�f�`�f�aBa��@Br@�`	�&E ��WUY� &VeUxǉҪ�*�2�ª�(0�� "�2�� NA� 
�2��
�0 �  L��ʪ̪����UY� &UVaUfUVe 	�`Y�fA��f�`Y�fQ�`e�u��H��0,��"�2�ʳ�N̋0,��̋0,³*� ~����s�:���F�I�PQJ�?ga-˳\�0о]�>=������s6<��s��;Ȕ����g����T 9���������=�� ��������O�/�O����� _��}Ῑ��M$��:�4�{����3����>�
���DXTII!eTBD�P XUV$ �U�UX  �� $ R ��H��<���,��~��<QhP� � f d(^.]�����xP�~\@@IH9dqԧY�|��������s�=���* 
��؇�O��}i�Q ~J�����!����~$ �
���밁@^�����i��p���x��� ���|��<>�@p
�����j���
���3��I��9|n������d��)hJ���0����j���]3�:
L]���G����>���<v�ﰓ��ʠ ��uA���L@� �����v��O6�%QPW�0>xr���|����br��
�2�ɡ/P,�R�����9�>�o��(Q�2M�%V�Ķ�%���UITiZ��(k@*J��H�aDHT�BQkl�T(հ��E���Q,e!�-��^�:ѭ[dҚ��������Jؠ��3��kfʊ��m��i3-�P(fe42ʌ�m��2��Z�[M-i�vͶeM� �V͢�kUl�mhKm�26d�$%��*fY��Ef��ڪ��V�6��jm�c5i��l�B*��Cm�1��6�F����j��  ����Y�pg@[؜�W5�kMuT�;k�٪	ۺ��Wm���uu�r��'9\�:���� ��׼-Coi���W��K��g��T6t��	���+,��c[%��  Xz(P�B��([��t�B�2hhP�z�"�
(P�{����(P���m���[�4�e��o{�����i�滵iGUۖm��MSEk׻��S7����wGm�ʻ�t%���Tb�-m��&[k|  ��t%����Ez��^����fq���l�v�mR�bk��j�)v�{u�;۽�f;�v��۹wgsf��ֆ��6�;Tݻ�H��C��w���ݸ��fi[$�IUmS2UW�  Ϟ�h�iۭ��v�S�;�ۇBۍ�[Q�4�pwYKr;�_{��h�8�5�q�hn�q�+����Ѫ�h�Zhms��h �nMT��b2!B�5m�   Ǻ�
=��WUZ�[�� 5լ��T��mv����lv*�tUn]���.u�h6(�Ut��#I��,��a��՛[�  �����;��QTh��Үڨ\�E4�\�P�d�wQڣVƓmm֕2�Ҁ�X�4�廕]VP�4նJ�U��ѫU�MU��  �Wl�+���T��c#�wS����#�� i�U�d@��Ӫ�E;e-��@J�oxǔ�cJ��a����mIk%[Y��%K�>  �}(��S��y�S;��Ҩ�[;^��R���e�֑n�g�P�lN�*Q:�k�7���F��E���P�׷����d�OJP�Z�a��mUkf��|  9��P$�+�޸z$�����t�\�K�@/`ѽ%ܩ%!R�F:HZ���[5E+q��EI;h+�ٻ�U5�^����^��B����ԉ�4��e�  s{�*�+��9�J�;݈F��r;ʶ��
��R�0'<����U%�z���PPo^�� 5�n�w�PU��X<�R "��JUi 4 E=��)*�2�)�1	JJ�F LE?i)Q@ h �o!���� $�JH�R�  1���?��I�O���.���{�
��0�C���!�3e��{�������}U�}��g������ڵ���[[mm�[mZ�ݭ��m�筶�m����[_�����;��V����ȹ.�J��16U�j�X�uj��ڈ�U/f�.� dlY�:�M3���y�fҭ,KW��h��1��p]J3e��h����y[�M	���8��5rS�`K�m�&1c�yp�n��xRtLFM�'�)c�c2�항bͦ�4(��Z �M��6f ��H7��|&��H��⦑Z0	wIʂ:���l��*�b@�c �U���,�v�4HL�3ǹ�j��ҵ�Pӈ�F+B�b^�&�$��˻$��D!�ɣ�˫��.F����Aor�%���;ۼj�L���jp	Fk9n�r��T�K��ɨ^�IA�Kn��ݔ�`�y����FR�b��6M�����dcEh�S`�"43�՘����*���M�:�.\�+���[��+ddRūH�K+dU��/F��I1�{���&Ry�6v(�Rm�C�6��U����Hط��imU;Z+HT��o
UCj1��U�[K*gi��u�*ų��@V�ᩣn9�]\�o���c1bk6YZ1�֭`T�c��su2Zn1�B�*v��Ѣ%�"�ݝ�nʚR;��L�u,`���Ki:5sK��N�U��*�v�<N�E���ɕ��	t�r�\������h�դ�=-�H�U����^[���5��$b�T<��\,�!��Ң�Mې�UF�Ln��Z7sw%Q��(�Kd��c��e������}y�롛�`łlYW�n&�?��ʒ��#z^��[I��S��8��uw�w�M��K����cK���*�2J�U�b�FU:�z2J3���Y��r�|В�ab˼h묉�2��D�
�ݘ�M�q���]Yq庼���1.md�kd9>ѻF�+qHe
�Yڊ��6L����j��ܛ�4��3.ވ��Vjc-��N����d�R�;�R�ʢKIP���6��nK�`Չ��;Rd��D��La�(��b�@��YǠ�I��M`y�0f����H����	��FKm%{J;�Z�5�b�Y4.�TsR֐�#MX@l˒1a,�|�%�������\a��#�@����o>7�$2�յu
��*l�7p�gW�^+���R����qP������2�%Z���׫3-Մ�¢���^ +r�^K��EwlV;�0��K�!B�uԳv[Ѣ�J���-��Q��a$vУH?��%�T�p����
�,3���f:�ݹ���K0�y�n/�`�6��"������
�e���cr��u≰�v1a��дe\SH�ZWi�V�'�r1*�	JM�Uw1&�'�odi�u���6�奧�!ɺ��$@]�@++ْ�KS��>���H�f�2��9Wkܷ{h`��9N���5{u�0�q��M��h�{����*˽��F�V��+�)�kyF�i�J���8.���4�wsʣ.�t+	ګ��/�'Sn�h�M�*
�-����[�m� �7�e�`�S�[3T����[�LQ�J����ƍJ�Y"9G?)��Wj����X�DTui�V��赫in�y{�cD�����w[�s,;дC��O@u�!Rؐ8���bՒb�+1P�h�X�Z�LS���*�
�{�f<oZ롔�F����J,[��P���� n���]j�0��,jj��\��ƋX�8DI�(��&�5���N�)ff�������uqV�L��0dܰ�5OM���=���b� X��A��.�,����iv�U�{��QLne�3I��"����@�D�E�Z]e!(3���R�������?��e�H�A���B�ٰ�������Ei����D\�Ы܇k ���T�B��.Lz��t��F��S��]�t��l��r�L��@�жi�)�c5����A���Jn�S6G.��ո6Jl,�q`�ȵ��Hڙ.6�+B�e2 'U ,��=Բ���qÊV��܌H�I�h%�u(�fnc-�4*)}����&��,U�y�-�Zf�Z�х��X��\Qe���mԩ��.�b��j�Z��(J#.�͑1��(i���;m�-Ʋ�Ö�f�rۡ�H(�&�f;��7>�mlN�m�	�e4٭�Pə6\E|��j�ųH�,��lf𒶉��a�/qbт�A>l�V�T��&'"Q����D��s)Q� /W��*bZ+)���@�2da��.�i�1�RS3�-�f�Ku���+�dѬR��J`�7m|���n�VS�*���ī���Ce��R�/�H���)b�T�i���-X��X��֑c�L����1��՜��.OX�f	���dbuce-g�m��Ŵ��[f$�dJua[�[�����l�F;�V7J�q�΄N����pڭ�E��]�տ$A����ڽ����P��;I�S�MmԲ�$�!�{w.�Q�ڕ�e�(hT���+�E+�XK�WZJ���|���i��(���!-�{M2�;Bf/��MT�%D�M�PpP�t��Oh���ql��M�C�9�Y�H�7]�l�P��$+��SxH[d�nK��f\Cr�
�*�AEl�.��^�."��'-'��V�iõ�)���,�/�r�g��%0�U��Y���/Aצ�R]��+�5�T7*�j�nlՇVthƕdù����jGyO%ZE<{�t�������Q���l�S�M�3T[�m2+e�P\�.谈n���Y5��c#0�
k�h����1'+]J�V	`MCZzj��aw�e�4��n[g5�u�d�X�I�75�f�9C,�u�	F�b����/	�`2C3	�13PK*���x�M:ӕ��6rG*ݗ�[��+z��:�a6,L�+5��jb�_������^$qӛ�i�p:��86�K��ԑ���6��XK�O;|�[���
K�_4��c���,����0,EA�`*�V]�M&�*�Y��^�
{�u�n�BIYQ:�j�*�e�Xmf��Y�m3�E�&�S�Eus^0�`��YN^��;�jL5�23m�s���[���㗕(eI1m�WlG�r�0���L�
���b��1�(�^^ejz©VB5�^\9JM��Rƭ�T��=�>��aԔ�V;ܧ�"De-Ư�.�	��K���/6�V���P5�C�g*��Na��
'ZU�l1����P�q�ŕ��U&�ȴCr5��(�	�V��Y�ݭٴ���f��a��9rmU���̅�R�]@�Vٙ�1�EJ�ji�[e(�Շ1,�-��|�J8԰Ҽͭ��]1���V�e�L��\���0f8��ͨ��U���LUi��f�s�oNR�����
���
�M�͐�(��'v��r��̬���5�/V�њ�aY���㖯l�K�K+NnK�zS�((d!�tMo}$6D�Q˫��$(��˨�Sӻp)�"͛[k
��hV]�p�,�5r�/s=%V��&5H�:S�Zr��sPAvΌN+�/vVbY�fÆ@�2kU#�P�NIY�K�2�n�!�2��n�Rh3^1{gl�"�T�gQ���6m�r�mK�h]� B��Jk��KG�ufVA�!���.V]����e��EY��f�@�ou!(Pw.=�.���a67
ff����P唱Rj����iI:t�nhYt�7��۶�^;��=U���a�1���E�7NM�fl�h.�-�9`��UJ�j:�����l�͎�W������U�ڊ�=�Nj��I@�����ٹB��m�	�i��׫Z�.i�a`��B	��-���ͼ̇�[m�.�h������r�c`� ��&,�������Ů�ۭ�oPs ��vt+)f�nk���ub�7�v�����@5�)���fԭ�S%^�IśB�d�Ck5S1*e)�x,nk��6��a�[;�nh*�\Ź�;�i�P��j���{x� Lz�`��Y!��t��P]sH�F���d�0k+���ا*i�sj� Z�77(�gn��P

�6�=�d���͌.�1�ǆ��h����)Mݤ`��.Sg#W��j�̢%Э+)[�2U��&DaF�!����Qܷ@Ht��y���bطK�[����Vd�fP�IV��6*bYF��*&�mji�Wo$�
-��Z*޷H�"��� l�u��ʁ`��E�e��ou�%��%��]�J6�OtEɳWĕ2����m"Nݩ-̣m�%4nʒ�̒-�v�n4���l�ӽE)�Ɂ�IH*�ҸMfL{iQ�+5��YGݩik8t�P�FQ��bї����tR�h�؞M���C�0֋��kv�{�:�܏�R�K��.m4�8f:����t[�m㚥��h�"�)O^� +jh��Vp����逝�y�de&�rkS7R_f�nֱ�L�&r�B�4�����<mҬ4iE(p!S%/zn]�Gx4ԅZ45 �IKuɼ
p��`0�̧��{51뽈����"V���mI���բ��ɧ �{OK̥��HfZ�1��M��!҆5+n�U�
B
*��`�T��,��3#�`��H���Ƣ�j��L�ѓmk��B����� ��x�el��eF�W�R�&�$�Լm����h��]�`��80��M��MCu3q1*Uu�LF��))6,F3f�V�b!6��
H�5*	�����9u��!}���;��Jr��.���3ie�U����� ��(--Ø6�����Q�;·]�6E+(��J̳Kt
�1��˙[��:܉^�T
k;e�U�#��������V�`��X��IP@����ǳse�i�6͜�mY痟j��{�� 	kfM������ǆDf���Q�Bpӎ���6R�x�jaX���G�Tu���dJj�*�8��շ ���Y��:�U]TfbC]Z��Y�.�N�m�f�*b����*^��o1E��RR�-�D��w�8NQ�٥��( ���r�1	3\Y����/7/U�J�Y�@�]Z�\�v �	�����6֍�������v֢2����K�z�f���
��`��lP�i淏]����ʻ�.���yj�F����Ie)W-��Kù{ӈf�/`׈l���dj��T%�4��/	㫵Tk\�ջ5`ڂf�/l�Y��;�f�7�Lqf���*L�KU�v�]����c9������51e���\j�'��iV`-����2"����cE�W��,3ҵ3 ��9Y�SIR�H@�uЪϣ��t�sSb�PWt��n�G4�WQYwfR_Oe�֗%���a��~V���	��{5��r*��"Jr�&ȬIJ���1	����їpݡj}`�V�\V2�(3�D\Ln��ܓ1-�Fֳ6�G.�U�ui5r�=�Q�eˌܰ�����{�Z�Qq�2R2��uހJ��oT��U5!� ڵ�eQ�X�1�&�Y��Dn�4��P�@����
��-;�z������Ч�*��Ҋ�)V����:��%�3L�)� *	��S�C��mңW.�s��^�N�2�sN��FBU�Q*X��l
0��^=� T �ݼ�[YN�u�V�QKH'Wm�k��3kuiN�TL6ebzkHr4v�h�"�و1ew'W�����8�dŦ�f۾�u����
Pk*a���G!�[��Pjչ -�qK�&�,���e^4��T,ti������m��Ec!�;����sF�foΐ�WA��i�V���!�[x*�E�X�Բp��d�W��j/e��+Z�UD�t�Һ-���v�vi�A��҃���D�^-�(!��I��^S܂j�Si31Y"S"(Ǘ�.�#f�!pɓV\�Q6ul���\D�� ��� T� ���z�!L�z�C�#�2��ݧE��J=Clո��F<ú��)�;A����T`�&c� ��Xf���vs%)�݅(�u���;{ ���mB��Ut�,�X(��M,�*䡎QR��yZ��0ko��gR�юٲKz�D\�M�r��#.T�C	����y�Y^�M��*�m"uP8�o�e��Y���h��9�� ������L��OfU�W�u�V&�*:�WC` zu[�]�=	.�,d�e�v�1�1bʲ��˲�.l��v���j�Z�:d��|���@�/��n��OAs%hj�\�m�	�'xb�4�Q��̫�3�K���S�&���Km�f�n����V*�֬*ͤ�R����Dw+T�g[B��j �[��xƻw��i�`�zE丢v��ec��2��̗��U$�CI��ۚ7V挕۽�{�K�J���k��WEg�hZ&eT�ި�&VՒk2GQ���N�K���ѡ������y��z>���HP�j�m��Jqc�zI����J���K��/Cp}x�@̵���i7Z��7�L�o�p�����V�zs%�w{N
e'�&���D��r�P�=	%A��ku^Cgu\?LҌt���ђ��R	���ƠH��U��F�e�ڻW�֍�A�
�����6�U>Ld��V���eF鬩��z��$�VM&���\JB������@�a�Y�(fL�(Xx�фiM҄�V4*�ȁ@M+V&]��Eu-GGNfƪ+�y�8��<Ő�4θ��YD2���@:'bP<&I��廕yW7 Rh���^�[M���&�+��a�E��ĭ���wz�X����&�ӢVq��QTYs%$홬��Y��z�gIz�9�钲�t�b�X �u��KP���I��ôʼ\ή��DѺ4e�_i�O!FylL��!+OoU�����6K��"�r�MNc;���~�(C>��ϫOe#�V|b��:�e��7Q����3�.+(r���V��ɳv��q���Ԧ�Nc�%����3�>�q<�X뜝{�f�,�x�9˟�<�k��/�ة��v�"^;�G�����odr-�:�9:��ebSsa�ۃF�J��PqR�w;Iǔkn�!찦ɪ��ݍ�	��]�k~�w\y�ʑ�O���4��e�+�oz����]������Gi�����uwxa�����e<k����t�P3����'���h��nZF`FL�D�s_Q���c�@Iw������guQ��+���̀=��iD�� ����Ƹ�F��C[���9�ձQwW����Ka����#d'��^��u���O ����v*ogMG����e�=�2�T�rS;�� S�;��-��b�������ETx0�V��W�{R�јF'�w}����Z �"mޞ%��@����(�`Y�U��q��8㑍�q5��|K�'Kז�)r��4�j��j�Ѽ��#fi6���0Xr#f�Vc���hl�.���9O�GH}���*:�ׂ<����n��fb�U��;��j�i0j��]f�.Z(J�C\��gg��N4���:��:��z��+*��HeC���H�0�F9����vU�&Ό�d����:��������k1䨏	p,<7:G�-n�\�2��r�2_e�:oIPL��+�{+�u9{Dkؖ@��Qf�Ep!�[�#/l���2;ԢN�B�n��[��H)c�W�v��8�s3gv��e�U}���85�	��ow*=���� ��s��ĉj@���uN����h_���<�d�<_�S�\���䴭�ܭ���=+��!%�-l�C7VJ���x�����[��N�Y�+�,脅��k���J�2�-R���Zo[n�����&�c����B���ܢ���kx�{3�����B �s��#Za�⎄�u�sn��+z�qM�}Y*i�o������3 jܬ, �df`���C�Bw+SU�բ�e����'6�4P#r�>A�.��$,��iN�Z&'V�SyX�{4�ɐ>�N�L�V��D-���V��ٚ`cz�m"Ƌ �I�+�Ʃ���HEO���t*�hoT9ƭ��tTɭ���͒��`��X��qĘ��I+��Y���	��t�$�e���w8�o9I�5���i��p��	(�ov�Th&�,W��%]�v����c�&�kp��Ë]%Gv���r����{��h�GtNxk$F���k7��n��M%[S��wJ(k�p���0��X��a�zJ��	g|3����{��F��ɑu58ve��9)�䷖{y�����q�ioÒqn�fol��S��0�ֳ�s�[���s&�Q�:us:�t���Dr`��+*���Ҁ�0�*�oEq�6��>�������5V�\ӥyZ΃%�k�Su�&�[ ��L�U�Sj�P��[�ŷ,�jH���.��NC�D�:�=�\c�,�֫����I.�u�Z��.o��Az�F`�3�f�tU�Yܰ�(f_�4<��v�R=��e���Yne���Ȕ�X�z�2-):��s�M�gh�{��M���s����gGIy&�n�C�q���:���m�l|{]f��V���T�k�e��ˬz'^f�Yt�%s�'�8�99�����7W�*`˚�V╷�(œ\V�Z���GBR�F�X��*|��'$46��Z��r����<�RYG����5y5(��@�m�?ouڏ��y3.Dr:��%w&H0�:<�=�7���sm��oH~���xf�ٱ��\6����f�]<���@���
�M���o57t��.���*�#p٘����)�Sj��%w���{$�TR�,��ј%����,�o׷�N��D[T\�9f��^�)� Ku��}�6]�o%����흗�i��;XR�9� ���{��WG+w�I��ԩc<��u�d�9�F��͕�b�f!ܰ�F���H-���;o��}ɺ�9P%n�	RY2����7c���3I��ҋ��+�w��O����iIg}Զ�G�<���Fw5q4��+B|FN�����Bx޾�@9��*݄i��θ3&"�Μd�
=��l\d̜�q�2�Q�l�%�-�sd *�.ᵼ�39��]���4�nZU��:>f�[�b�e[�d��]\��pS�3f��{��mt���/�Wrå�n�m3�.�
��V���0�Tm��ň���]R�-� -��6[�,M��[s�l� ��{ݿ,��k-���+lwI��j���L��2��u�F���b�=���� :��X9�:Y],C!$GzjN�C���9�"�N��c׮I�,ξ�v����t$�`�w;!rdmv�� N�:୰5��z��-���4b�^�3^�V��gs���۶HR�r�����|�8�w�A'�C#�f�(���.�V�̆���t����|�\�734;�������pQ�Ύ[:��;s���=|�T4�xS�U��VW�KJY�Ms���\~U��C���S���Ӫ���Q�3�N��&�7��u�Yhkj	`�pcH2�86�
���E��ۨ��lK���+a�Sy����N���q5�d�[m�� ��ݽ��Ɉg
�x�L��-��<��ˌb�E��eV];�k��&�<��5x�v��uRY�bK�Ր=���Ì������W�KH��ۣܥZ�(:�4�s3T{-A�7�`�Qe!�ɵ��&S�2$�}�1;M��x_�K�}o��A1��w%���f
S�p��0T�7;B'W-��m��N��1�y�9R�N͍i�Bl�]E�O��-��U�F0��;��U�X���ε�^���Tǉ[15X<�1���P�t)��h�I_��+�P�L�w)�}���t���]V�rJ�yL{�;J�jp����'�!M����#;oKjq
��Ep�ƓT�}�`I�m>³��LC�:���M�q��8l�f�\7)sF�e�y���@�HiPֳ����-h]�1�����WN�M�����1a{����NrRli-����i��W>��c�,�s;FX�X���ˬlq��_��Ɂt�y���^�e0.9��y��l���I7זldX ����4Q� 4��!H)��9�c\�\#��ԥ���yG:p���^�#O�H.Z�k/ô/u��+�1F��w��eIq^����և�M�;V�M���)�C�I�e��',�{z���*��ųt��mn��cK�"��^ӯL�A/.���p�LR<ż�ɵ�l}u�gQ#{�dJ(n���4+��mDh@N=6��xYf�S ݛ��ʡ���J�S4�:Tr%���;r�.�;����ٮ�f���W"˾�=�v1��R|�1��Z�h��Zy_M���� �����]9�r�Rl��Jt��nVw`�V��j��6�3t�K�vڱB�z�m�§S�:( e�t���[Cz|\7�(7᳕��R��o��y�9�.u�L�	�o��6qR�A�S�ȍ.κ�.����Rj����Sa�߷����)�WST���oa틌�����֖V<l����ˉ��˨S���@�R�u!���%vQ#" ���p�]�ř��Q�Qҕv�ʘ+��� C�X�	�� ې�|�S��մ*�oF��(U�"� �A����Ȗ�'�27T+���+�t�[|rpE���t��.0�+9���¶>�C���qK8��W�F�u�I�M�ίdpjT�:���]-u���S�&i�2�MI���Y/,ϗdV��:iU�+q^cZ�[g2�H{4�4`���xƍō
FZ�,��&�:��m��yr�2zqN������b����I�H�^.T]�Qh�VR[vZ����Z�Xt�[:&l霅�e��D�LU�5�e�So�$N�yB�J&ř������g"��&��vi���3�m���A�<�n����������*�ڳ�Ef�Ydf n���;���hdC6���̻�VTj1y)���
DvK�0�W��î�v��t��;s�2s�C�gG�٘���yN�O:ҫ��Lܗ��Z�m����=�Ƈn$S%��Ӗ�m#K����u�7�fto��[w���_Q딮t�-�;(g4�f�Թ��7q�� U�ݘx�@rаjcOP�]��p�� �*;��f�}��hƢz+�+T�X*�^�lZ����E�b�\5�{��ʬ�^�ݩ:54S�;�=m�b7@����&s ��!ћ�m�]��O�^��Y�WX��ah8��t��z�ԕ���M �s,e��9��	�T��gE҆���E�v�f�Ƅ�����Q�tj�\���> �[��U��_�6���c��b}�9�y=ۣ��n�%˲��t�Yz�}#�Ԗeu��T2�tŇ��E���=�b�aքk������N�H��\�c\@.�-��U��8Th���T��t����Ͳ�.����vm	˷���Z�i&�sܺ1}O������U�|^l��627�]o�L�t.*�:l�*)���e�Lvq��2uu�\3�2:.���Dt�`i>y,�e��q:�S�W����x��*���X�D�kq|#W�`h 4�]�q���]��Ce>��V䥋2ׯ�n-y��M��w�U�T�͛�yK#	dWq���{�r��9�8��:��/Jj1חeѠ��q�5SaNɇ�mF���+W�5���]%V�N��5ү��t�Vճ�Lp]�:��� 8K�Ԩ�F��Qk)�4wS���1سH����Ȗ	hҮ|���+�W�d�ۓ`��5̫%�+���{M����d6�Q�wi��Zn�.#�sM�n�9[8�Ҵ��=Kd�ב�<=Y���E�|���IdPM:5/���
�k6�B���Í��k'q�������c�Y�+Zyɦ!:�BotΣn�<��+��mLt+9p���f���-�@0毢A��=/:��f�6u���r�vB�Y�X��aD%�}{�DwOiC)����M���p�y�Z� �Sn�2� ���c$:�-��o*{|�ە�����uj�"oEou+��KÄ�:0wf�3#<\&��[y�m�cF�Q�II�x#m�0�M����*�t��opFͼ����фc��]�|Ua�Z��4h�͉m+l!&���jR�)�6�,�S�����`R<�3d�]��Ke�cI�N}@:{䗻(�۳R�5����F�]�&cs�&���v�r�۴Vpf�m����[��8�l0�*��
\0�2ec��ۊ��.d��٫���G��U��rV�4=qQ9�ـR�y�ˣW�t�7B��#hYz�c]u�3�C�������I��.�[+\f0L��h>r��e(��s֔p�N�<U���1gA�l�W(-Ύ�1\t�seD�}�1n��d).�+BJ�/eI�-[:�F��.��Oxٔ��w�5���b�͛ ���"�ȩ+��z��H��c��1���7Q�}�ju��R՝������fq��1�Uf[�tn���Bx1������p!�z���'��qTڔ�*�͎�����C��\k��8�k�.�w^!��6�R| w����[���3�1&�<���y��	Ҏ�&�aa�VTH��b�iđ8a�J�bײ�ƹ�M���6�Rވ)��rT��J�W1��/��Tښ_'5���J���O�n�����B����p��7�M��m`�KVg,��۬����m'Q�5��*�.��~�L�˂�����8�˱���꓄9K y<��ݳ"��=�Տ��Y2\����=�ݘ��*W :G �|�3�����t�Ē�;Y�t�����u5Z��*�@]�l]������o�����ҳ�-�vW3����U��>B 9Iwfٓk*]3Kn�yYCOWc�(�Ȩ
� WmAз�7N�N�D��,��d6�~;�=Zg{77��r�Y;�%Ct{��*l�c���j��X<���W|���:c��p�4�x��˝D�Rj�]oX� S��Ld�ѽ ��#�Gn>����d��᧦���w�A+[��;�!�Autn�u����V��Id�r��&���3��k��mq�ԍ;޾� N���
�N���}�1��]�2QF���'�6�2.���]Z�J+��������e�U%��ˊ���B�?����fj%��p�j�\Y �.t�W"��&�e@f�{�iu�(F�BU����hmZ^.�&ڹP�bIS!V�RܽՉ��=�&��R9�u*����yיsO&�#���]��C�k��$�*v[�r���N��$�J�3V�����ϥ4��e�7h��<NX�Ko6Bj���]ݻΟ���{��+/��i�]�F��$�x�ଘ��$�Εiz�	�md(Yꉌ��M�r��ȸ(�? _Ky�r�wʵ*�#�gu���es^�N�S �
I�}�*��U-��V1d�Or��g��39��[��p:Q�q��,gP�1��^^��p���ٵ�P7&�Y8s,�x��}R�Ў�tծ��V��ح���S��f��+p�[.-q���ѹYd6�m��bb�DA��iBk��W����Et��K�D��T���rS�1:V�|��XN�(7�f��Z��muXީJi��4'u�Z��b7N��W9��Lp��[��,�$��-�`�n��/&��6V�rel���$����#MH$�d��L�9w�$N�ﾯ��������G�}�G���y��4(�{5����Q��a�Qi1�[�otne�xQ{�n�nd��>:�0�n�[γ���f�H��x���跻��s��Rۅ�F���}���-�I>�6�ڮOsB��ko��`ܢ�2�6�k��v`��=�Ӏu�8,jw��3�͹�B4�d�ةsVoq�  ��b�F8u�fj�����Gʖq�_�a�������;��Ьgrԏ9��m�N����R��`ի�v$��v��|RJ�+z�';5����ee��lT8�B�꭮��$��|Aۘ��ͤMы���"��5|4ॹ�c'�i�V^V9I�b�O�����ڄ��1o	�qZ:�n�D��em�@�3w}��Mʗe�WPj��n{��n��ë�ի��7ge�q��Z"�Mu��E"9)��{2I3�e�R�H�.]�6y�ï�Sg@�펱���]��.U�V�ZP�O�n� m�C:J��K�9)ua��ma-��W��mdq�.���5�P����,sM���Y�a*��%��mC}�0u֩cjw,�ھ���7�v�S���C���u !�0�w��k�_ӆ�h8�5��H��1hàV�H-�T��
���x��&X�����������W,t���k�S�y�5��"�d:�NUz&�2YT:�1P,ɇW}���p4��`���=��]�t�I@�h)��mK}p�+4Ǐd�߂/�6�t�����V)nP�WuG*(�ǚ2���tjE�B ��S�Z5��U�ns��%+�[c����*#�Vq�Qz .e:ݻ�
��X_cfWf��ݷ+�A�����������\lm�|h1�R�$�dH�N��lnʆ�n۴SD�+�����9�8k�� `��L�-���\��VKŧ�a��&{���㲎	�J��݊�fT1	U{��a5�&��p�R�t��v��U���8kKCⲢ\v,x��t���!v6JeGN�iKj��"������L���i�м'u���3b�{K��v3S�hl��O�&�i
�䮬1%H��uu��R�++i��׺����ւ�t �[���͌foC���ݺ<����»{2��l�^u���Dڲ6h_k�A1�+�*�M�R����V:J�%t��%��34R[�������f�p��6�����'<��dƵ(�Q�a?^Z�[�_f#J́��1�Z�������us�R�l�.�N@{EC�K��V�{.57�졪"�b�14w�j��Ħ�ӧSIi����MҧBއZ��T�k�c5���*�������Y� ��1d--ᓩ��[Z��TWn���` {2�-�v����j��WH]�V��h|�lQ��v�ms��1�_.�\(���g6�����p��j�4'��ޡ���>��T����u��닔r��;4dJ���5�yr
t�b�6��i����(�r��^s�)bZ� �k7���Sw �7ת#)�r���郄͆��:�!%����;j=ˎ����z���R�H]��!�+'	�� |s��T��ǭ(*^���K�ס����<ڕ�&��W�5-�V� �G��q����B2f���!h*J�i�/+]��T|mo)v�Y�X�qe���	赻"ܽ��Y�2����S��[C`M�^3z��'M�hC{���"� !��5j�E�0L�Q�r%p�@�����aM�o��WN����xLWC]v��r�꼏����c���p�Uc��0�j�!��`���c&<X�� �A����m �o3���T��,�wʯ�gv�5`��.��
�Vi�il����K����E�'�%�"WEh�;���m���t_%��$}�#{�Ƞ���3�^g�����w�Rz��|�y�G����K��V�Y�rF�v}�,�62�X�ظ�սNȌ���y$oU����+n?���H��ѽ��T{v4�S�r��*���6�� ��ۨfG5q��1�iU�&�K�ڳ&wJ�b�2�2�m�'u!Ϟ\���k�u5�	�y��$�������1Q�B��=�c my[i�][C�\�h����P⬣%��˛��X�U¤�-���j�h��3q��
9��l*�9�#S���������yM]�4�ņsi"g<�s;(ɉrov�;e�}��(��0��P�oU�:I����rgVb�v���E�0��g>�דB&N'�������٧1�QP!C*�5���tXɴR��J�4o�0��;l�`p8&,y�Es8j�A�С���[�;L�3���w�꾭��]��3�oT�OG����-R�ʘ��\H����|�{DiZ���m^�m�@�5т뵩�F�K�*�Y���Ȫ;�ڀ��&��f���� gJr:��vfN]��Tܶ�/4nШ�4�:]18�Pq7K6o[ٗ�E^�H�A;�b���J2��ړ���h;�-fHͦ��ԩ�K��46�󷒢{FYW�eD�v�J�͡�MZ��\�4�)s�� 롅�M�giҥy�l<{��)Ӌlckjo��u��{X�����2��0����#�M_a���
�.��t��	�^�@���6��ެ���x̸���2�%U�3�ܒb�M�QQ��Xf6�%Ɓ�-ɑϬ���'�n
���ƩY���R������(v�h�\�j�Pw��l���N��9G]�$ȣG��y�L��%�q����.I[��k���w�5�S�J����a��r�`*gV���eb�ڵ�����E�[��-��w���1�
�僋V���L�Of���fJ��Ѐ�u�4x�77W$�g1�5����.V7v�i���0��F�hhc�r`��S��5�m>�x������9=̼Ur�KOjsߍ>Z��1[�n���U��	�nR��4+)��;���r����uc�,gcQ�ހڽ�ٶIKv�;�����+!}s�@�*m�i	1E��0�u�f���G�j�u9H���Ů��aݬ���J���ѼY�WY-�����B�ɼ�PJ4�_}����v��c�'���/�;Xٺ,���� �G��Ǳ�
+L�Ee�D�
sGh�;5!&�tU��@o�j��,ՐǹFf���@�Եe���i"tJ}l�t�
V�M	�^&-���q�0f@��fm��jf�#k0�f8�vn֙>7�9y`��n�S-��Q5"�6��$�6����l���6vkjh���5��:h�s���ҩĝ�܋\��iJ��ʏ6��A�l�ڎ*7�åY&	I}с�ʶ8���K��x���4ծ�1�Z���S�c��N4���%ؙ;�72ʓ�1�fi��8�[�7{�,�it���tݍw]bC�RŮ� �Ug .>���̑��z�r�7{W-.'Z���Q��Q�i�������h��fk�����%m���ީa�݊7���{J��  �y>����)W�m<������ڹԎN���4��Ϋ������8;n�c�X���G�qY�6l�u���ؑ�$���/z���z��bn�}t�D:��˝B�r����bgacGfAcUӆ�厜��?(�m�-�{��J��+l>��KG0ze�U}��9:It�@<.e�Ұ���76�ܥ��eԃ��$��S�4�s��٧���6�~�����Jު��t�_Q���;S�D��v|���A��)�opCO4�U�/�
E�Gqa�ͬ�n���fs���l`�tjN��w=�C^�j���<�/�[4�hSW�%.�tz�����-��䶠���ʐڦG۹������J�*MJ��wJ��X`����4��Q�g�!@0��T��@�������A�*�P�����luv`� �%��t�:BF[1�R��3[�e�i��{@�q���gf����E�?\��J�[P�û�-�Di{���lP����^&�e
쬲��d����5[�ؖj>5���C�b��kŰR���)��%d��vbކ��u�E��B�
���ձ�-5x`|7gy+.r�`\���.�K8XA
;�?�(P��9ReZQ���1ޗ�6f}����IbM�J��B�׏�k�X`;�U��:�4�Sj� g7f��fJ1�i�@������N�P��[�Va׹BO�n ��:cQ��Uٕ�̷3�ͫ�j�l'�&��U���1�3@��H���w|�I;�*Z�?^E}i�	������(n�E-��f��I�z�Obe[�������֋c�S^d!ܺ�g\��g��k�h��Ӵ��,}��8F��(:���WD5��iJ���i���bT����݅]i���TeN�CzA�!*u��2���q��=³�Z)��k�-h�X����^�̙ �S�̚�)6��Kw+`�c�òɂ�Wo
�k�ki�U�x��i�)Ø{R�J�p�`��
kWA�қ�Z�>{�n���Z�(��KH�FYx9�T	G)�V����ًh��Y�8��n�˺�Y�7!��'�tj^�3>��ɯE��_�v�W#n����f�c�@^���Hz�nR�Ww���(6�]M�Yp,���6���h#�y�� ��0��2���R�e�;ŵ�S�fX�t�+U����ӫk2���,��j֌��H����U����Q�"Q�}��%<�W
�7#��*��-���ej�E7[N�������1.�4S�9��E��\J��"��X1KU���gb3G!]�pڴ�ݚ��K$[ML����u ,ޖ�쮝8��N�S֊�s�v$��̉��]�����}��N������j�����q/w��֡���5vk'N��AU�J-�v��i���-e�MƑ��U����lrb���6�w�+r%�� ���0K�_m�'Gj�K�v��P[ua :,ՑQ�s��z.��dJ�yL�ǒn`K"�޸)L-�-p�4tO�-=}]��[�I�Oi�U�X��rC�R�	p��n����0[-�ێ���[ة�D�.�����.�n�G����c,mk;�Z];u$�ZwΗ�;v��։A ��h��#-�7�����>\�E^��$0(;U�Cz�ŚI`Ž��%{�E�v]�ݑ�Ӛ
+�LL"�$���7i�
���52���AVmG�+S�>�*+����N�]#r�+�v��by�R�9р�O�����Qu�՜������ZY���P0��-��3u�9�/]cF�$��31M�|�&�)j�1�h�<��%�A��ܟ)���ؐg*o
�C�]4�b�%��˅c���n�Ba���2�	�7�+�P޼�Ō�y\���ԑ0{�nN����s	��7��Nâ)�a'��F��J�{@Һ���JS����b�&=�\��s���������;)��ևJ̕%ˣ�����(VN�1E�o���͔8R�)घ;R*��0J{��^)@�w4j
��K�-QYR�a��!Sv[�@��ފ��mmn��9� ���P���%�Ի�X�F~m��%2^[��Zv��x�`4�2�B�+b}�{*j�r�mꌮ!��ntW���T�G<��/�&���9��H�,�u-wjr�u3���C��]�n��x���&�A�uq6:��C^�Dh��vʽ�a�ER¸7�2��C�>�f�ws5�ݺ�r�c=BF�ep7RT��,;G*;�������}���l݂g���dlׁ�,e޺�ًk+'ܮ�)��36^��-X��pI�F�&|�H���n:20;a��J���QM�L�]̃��8�@�ƕ�X�a���N��W��M<�X՗.T����D����%�C-�;9gܛu��)u��',�_}���y��YW���QL�w�7b�B��7)�I�x�5�����0ٽO��Z�|��^u���ְX�h��V3f���I�g��:휦�D�}��9�����-��Y4�[�z���0�l��T��Q���j��yc��ͥa��9��Iǹ�(�>(`�]WU;�׎��ӹ�ι\*0��]�[r���t�}�eJ�b����QFe�:�*�c*���$��S��\YNV��lP��/�����7,�V���9�f�I�-jF�v�A��5���eԳ��]˦0Ͱ�P�k�J���%��9�xt7A���u��w��5-Z#:��*d��}jbm�L<{�0�h��a���o{T�k��QD���S팙z-6��1_Rz�iR�wAD��Q9��u9��%7���ָ��Q8�k����pQ�ݖ��2�q:�������N�*��v1��1�ka���� #���7%���!*�eD\�H�F�!o[�-�v�p��8T�6s��xm,��Sl��b�"[�Ҵ��`슺��|ݶ+au�m�S��Jn����d^f�s_��g	q�Ni�\�e�vgX\�ԛ����R�alMq��؆-�o��0�:���.W	0d��Eު]�ZJ*�O�/���j:X�{�ZelH-p�@�lG�6���m���Z�� 7{�YhV`9��N��>�4���� �[�Osd�5u�
TѸ�.��7�t2ҫ��Q'y���n����\��P�n�;o�.�{ݏi�J��E�f���2��Ŧ�������^��j[�t5�C�ص��:v,ۺ5�3��l�Stit!	���_B>���<��Ҙ���}uػn��c
a��tq��w`W�G��:�K�]�\�PAWI^b��e5�"��.��킲�rя⻫8Yȅ��'*���(�
|$����^�|�-M 8;q�ڬ�%$��߫������ﶯ�Q������ΉE��qD�Œ]�Yx�)C�g�b5g0P��A��)����Rpo3�f�ZN���_O��/S�#]���;��Gr��I:-p�Kd�sAC�
uc��ƺ�:N)�w��@�D�oiv�}�����n�8se��C:ac�^�2��&[��� ��ޥYs��̵�hJsjΣ�Y�y�u\4��:�F�ƥ�L������e֊Oq�S�Oflt�A�Șe-IpNBEX���n��z)������ꐮ��v:�O��a�2�(_H����\f-�)�T���'ײ���ܯl�woZ7%��C�dh�Rss��~'a� ��&Ju��f��:l���چ�Z̟%��Cn�e$��.螥k2���]\z�9�]?�v�W\�H�)��K��8��F���coF�᲏
ܘe����>�NF��M(�N���u< ���#oz����kgwץ�JS�W(�j�JG���5�Дfu�����m0�BU��գ�v�3��m��E��jT�f��6G{j��'A�����t-7o
�ݚ�5��ra/b;R$�GF��NL]��\�j%�	�vj�H��kR�8�뾰���s�)+���ʻ�Z��b����\�1<8�L&�6n�h[��@���P��|�_	A�1���PK3>���n�.������_�޿ezWw-s�ͮnr�m��\��b�\�wb����k�s���\���1����wpY*�q�۔<n��ݽ*��dm�u�鱈�E�,QHn�n���a�u�5��[�t�67-9ۺ�\�ѱ��N��D/:�1ndԘ��*L�\�\�v�����.sF����cAs�]�%Њs��z��b�w �˳Qn^���*=.[�4˝˧;;����#r☋����.��wwu�b3"6��XѶ,;����E˙ ��������Ơwzx�āF��H�4��^#�I"��� �S�=w6*��g�(�{�(���p�24��2_n�&�q)RH��(��*<��u�nP���C'J�~uہ�R�3J������i�_}0�����E��� lZ��T;VYB�Zv�
��u�:2� p�x_�ޕ3���Y���#�V�E8ҳn���b ���8��*Zc�AX�b�9d4���G��s�g%qZۅ|���>����_ѥl�_��nP���+k�^�i8MCe0��q��K^޽X�Uiݮ��s\$�vjw_�Q�P���D�T|a#'�k}+Vڐ_f�o�IA���i�Q��C�\1.u����:�c*�p�`ʑY@S�y����V�\��CE��8r��\	�V���+N��3�\��_��Zu�Ƣ�KѶ���v���3��:7� `�g������CR*܈}�{�ڿ?
��7@�Tmx�^��/���	�/���X���'	�A�_TI�ƠhP���W:zxf��#3m]ƪy�*["�[�h��T��ŢP�j��ip������
9S�=U+�ҕ�8J�U��u�9Ie���ڏ�u� R+~��� `�:y���BѸ2��D�4�Ҽ�b���K���w0�@o�}��O����]*��8SAM�U�9������f��$�VEL�٥^�+�]���4�:*u̜���ιfv��"ȃ86_hW��8*g&M���Kr�P9V�ܶ�Nm.��;:
ἹԜ�N gV��z��
�?8J�8�B�_K,p��k���9U��~ʇ0�*�%���%���y��D�ҙ��#�!@`��C9)9�FtED-uÆ:j��sK��q/]D����=��'�7k �W��R5X���"�:L\KU�g�py��b]P�W��&���uR��Ӕ��;��e��L�б\H��:�Da#�Vӣqґ��W�����U�7LT��"���b�K{T,��B5�� �����~T�F/��x5<q�M�ǽ[�aR�>H��;�i�	��AnS&Kn@֡��\b�3��<#"����J�m����
���zWU�-����k��5��;u^��=�Y���-WL|��k�4q,���s���R_��W��<5<3�{eL�!��g��UO8s��X�<�` ���k��b�'y����a\T��P8v� t^��.!g��뙋�43K���vD-[��(P���&�7]xNc�u���_*�u���;� -�s!֫��I�J���=�A՘����hR����u9��-j�\�5��#ݻy�ٵ�m�����w�J)G3 @��=�s�0���Z?y,r��J骖$bʻ��5e��VP2CP�ި12�[c,�nwN�V7gV:t1NsA<<���*��K�$0ŧs	�N��ⱝ�cu(��e��𦊺���࿲-F��0^R]�����7�CP���*��Y�@��v�9����Ȳ\n�Evۿ�V_ͷQ�of�ี$�5@;� �w�O��.D�[!�魡�Mu�P&76~�5���e�l�ySw��W�C��.�"��:w��-_�okӗG�1\=Wz����_���t���l}p�:C1�v�W��3�|(G�)����5���}웛8�ŒW��@�H������%���p��cZ�h���f��i�N3r����N�rT����F�Bs�PS����2���R��q��n_�j烃�Iz�6K'���0�NTF��7�:�'���
U������'��P��}I��7.vN�%�^��n�|�WN�Y��n�lA�2J�$�w�`<"��0�-�@�ޫ~�q�F�ü���f2��rm�����q���k@�Sh�_AV���լ�%�=��Gw�t�g��N�#D���ž���:!��d��Iٓ'1��j2+e�j8�zl!p� �� �:��m�V]�o9Rw*��(;hW� {j�!�u��H��n��8+���%%�}�%<��'����c�����i�[�0�2XYI�֥k�|վ����o[n����ˎ�]�N���]��]IE���>�Ւ�wgt?�V4@BQm����ZMμSK߳�@�4�yT�ar��/�[�����e��%�U
��\�7�M�iѦǼxW
mU���|{��.��zƌE������N�2��k���鬧<���Ju�b�G�\Tï;hS�'(X�t��+��h�T�`�����V�*�gB�2��G�=y�I�y������G?z=�膶�4���?�j%����P�V��ıj�ҭ붔��8�޸Y���NэG��w9�<"��
�G߉��ν6��}[ǎY\���bZw�	7#zF8P�4y�
�t�Y]�)��)�a����t�=��Sƺ���q�-�(��xFN��������r�t7)��u���3�~�co6�\��<l��}�T�v`R~�2g�����7h}�=T#��X>e����k1ܔa����f�euD���t��UzG�1 (�}~b�� j�n���ȏ�C��fo��q���}�Ҍ8j{�"i�lhm�\��A.� z'%0�P4$U�ڱ�nOX���c0TzF���#h���5�ɜ;��}c�.s;Q'cܼ�y"����z�ɵuh�Lgk��l*��(�I8��4\�|���-3aN=��Zu�jԥ�^rʱ�hȗ=hp� �{���#ζ�vTP!sX�禺VbѶp���W&a�Yc���x���;� Tu����^O�r@�U(�c��A�_^-o�G�-\�Rٴ[�]z���yt��.�0��h㙌M���uLȥ$A�0�9{�B
��^h�ܼ�5���jh]oT1��s���aZG����y�x�����'��˚��N�;�N�@���GPʂ�^��~#7Lb��R�L��R�l��&h�	�]Iv��ެq:�D����@��Ǣ�}�0�Yu���\)v�?	U��솫+��cfާ���ԞBd�����&+��&߉�@��Q�Ƶ�qc�J�+�q9�c��Wy;ׄ+���o�y�.����˸�5�8I�C��򨛦3贫E�kHaӾz���7r���R7���L<1p���5}�UiLZ"�(J\��r�3E�\f�^��
Z�tt��=G�,2r�i[�d1����.u����:�aU-�(n��2J(�ݞw�*�;�ۅW5��] Ō	�V���ӿ��d�F��c�鳊D�p�(���+��O��ɺ��ܝ!�U���}SsD����P\!̻����k�Xp�ѫ��]���ǁ�!mf�4\[���0W]�0��#ֶ��',iL�K�[�v�j�w&-$��eZfí����ZU������+�P^NMT����4t�v�K������@$�+�
��\�>
���#b���g:ԭ�I�S��ߢ%���Qx�\6�ʛm���N�'�Q\�hסcGP(��U�(�,sw�X�����w^��,p�_�n1KT�d�h��&8p$�%�!��<k�U�7�x�ф�{m��:�-3���_rv��K/L`�1�θB��E\`�L�u[GxViY�$�=���[*��fw��?O9c�k]�v9�Ү3�S�B
����Fn�/��|r�n�r��.���;�g��ߑ�_-uÆC��������u�M�w�Y�#�il�7�}��:>7��'�CCCf��S�3nLp{��b��\�&���&�
9(�����;����ܰ�έ,�T�F��+iѺ�H��r��|��Ռ��@����zc�l:(��\�؝�� ��� �������;Ř�T{^
9���O2n�uo]�v��תl�ݷ��j���)�&�@sbdo�J�U�P�e=�L���R�p�P��a�w2�+�y�Y��"J�<:Y�%�,u�w2.Z�9�^���⅔❏�6���q���X�ȫr�<E��J.�Jݓ��Z��<��� ��%;�u��W��na�F��J��Ja^��Ķva�٣-��J�QM���m��ɥs'X�(�^�+�G���{o�dk��5n\��w�n8�3��� tdL��xr��j�fQ�4&a��_u��b�͔��a����Fjt8���_�w��f���f�+S�t�iOFO<\3��ٟ��*a�/��@
���1q�8��7\�u���')�Ϋ����u�
#��7���jpg��6k'�N�
� �wY1g�.AUis����Fq,��ݛ��p��{\/�ȵu�>&�K����U?7�CU�/ٳ,��"v_u�眮�c�B&�9�_m���e�ۇQ��ԜjI0Q8:73��}��.I#�{�'��l��]@�����W��Ls��۔��n��F�(鋬��b���Sj+�[��y�݁�|*��(�T�k�3H,�폮Hf9���6�l�l-���bgqg[�e�� ���z�΁��pvc��}�7�$[�c�5�ь}'Sܻz�mm�k�K-mD��N�s�"
�>��Yb�Pg��/=�u��#���pN{�a�*���슕�HzU��V�[�x�$�t�Tm;���d��W(f���fk�n��͜���qo\ŚLe�p/F�y��{,�1Y|K#�N��^W$XFA��*���ٸ���X���Ի��	�a+��0Q�`	n�ʗ�wv�C3�
���&^C=U��Bo�j�7�pYJd�������� �Zi\^!?g��p��XڤОX��.��?=ݮg!���C���|6 �)�W�R��`<"i�f�4i�g	n��]��_nE�#�?����7���k�ɸ��8C�q����Sh�� �����W\ngr�t&V��!˘�"�,�Zb�V��Ha�0�N̛Nb5�5���7=͔���_jo��<�a:��Πf�^�\����M������݇Bx_��x���M��t����Q:��8C�ULƁyx������?:��o�P����E��Sl+g]�7��85���(,=�HeGm
���W���#2붔^���AP=���<��)H��z������ ToOۂ���O��h|�ko��K��G�JQ,"�\d�)T���J�9最1��Q���!T�2�أ�\6���[��U��\����e�^�c�s�';����`�S��9�G��!���`(ن#a��X9�:L�������1q�ӧY�q%���v3B.��u�X���QU����&e�,̔Vi�ˮ9Q�*��qeNAKԹ�4��*��Gt�2�
�0�߸^��+L�*�g�3�R��9�&o*���җ�Y�g����8e�Z�CD�0+}'l�uY����eYX�f���$�*oWE�vu�}E��X�az�â���"�UVua`�_ �9b9����w��U�ɲ�n(��a����cP�Y�+UQ�����4�7T�H��Ghmތ��a�_>�>�m���W۝��'d[�}���7J։t-\>$󢾢=sew-�^2��_8�n��X�/g��dL�:ĦȂ��8?&�������Ɏ� z&� �*�4w[�����O�{X���0��V=�=ǔ�1�s��ꇎ�eÚFj�": ���4�g(|raK"��kJw��KW��R�b3��q���\;!S��d�-LX����uLȥ2Q���s{�f*]!�����z�ε�z�f�r���cqa۞m5���E��J�f��CnN*xT,uUۡ&N�P��|e�v&a8=f2N�&��W���VC�Q��T�{ +�R6Ч��6Ktl�+�Q�O��œ� �Znʊ�OX�z�m}�j]eG��Z�ƚ�r#0 �-�r]j�tٻ��O 86X_|���u���Yj,ײ����B��;J"�]'Y�^�Ҷkċ�ڴ}�t��v<��K�:��� R�crb�Q7�X�O���hV�f4T�]������etW�����lN̽<��`��!'FF�_a%+W{���3��sI��"�*v^�U��qE10&�v��j��ǃ9g�	,}�goN����vlF�'w�S��h}��]�	��t�2�����s��ݻ�k�*����n+i"x�ˌ�w��0�Ť�WQ�UQ�Ah��?!�E�]}^��iw�n�3�b�OP���\G�gG.;iQ��C����Q�n�ods�F��/ncd�cƁ��%�.8����_
��VV��`x]���(*N�
]&v�,A���\���}V���ѵ������v|JVg� h�e��U��J:dDRRE���T{P��;�G���Y독u�/8<&R��nF]�$験̂��!���b�\O&d����w��WR���������f.Z�8����&&8�Iډ�ߞT������{��У-`��}4��_"�	�\��h�^���mCθ@
�*��uw~�阮�|���@RE�9�3[?wت��N~�X�a�Z�#�s��Y�~�sB/�܈Ӷ{��[���qŪQj�3IO59Ќ��k��_1xP��q#���gh�}�E���ʲXݬ�Y��Qw0�%}l5���:�MG�.��&�;+yn2�]��J��tyG������P�W_�:ܮB�������-�O����u��ry�Y�3jj�4S��8h�]Q�P̂��i�,�U���v���+m%]�R��ra|xR�l�����3F�co�N=��r�66�2��'�:A���/Bm�Z;V��;Go]D���+���;�cWe�X��C��uz��:�j-p��K_�|"���{�YX6[��C�8z�������ZݘH�Ж�@����ռY��xMn�j6��t��<�Xr�N���x��i^�Yh�y�����8��#�M��΋6��շ1��Y�u�4�����l�yX7V-ѭc=�IZ=��r�?3Wg�u�^oi�x���X�W��32P��0�wm�YHrM�:u��cG�.p.��d��*eFv���t�1����xļ��g �L���p1�S:�P��F�����C���W�.� cїȗ�g-�YjK_ek�չ�a
���]V�5�����hP��]ؔ7����it�9'%�&n'�(0.��Y,��,����S�ثV۩�-C�6W5*<JV^`>r�49u�C�)�T�9��Y�0���;�9Y��C6�c)��=N���̛KX����;�RŸ�=�+�ב�o2�u+�Qϐɜ�(��t�D��>1ؼU���Z���׺R�*���T�L )�"m�V�9�K5n��e�:޶���V���8�I5��nn�å�p5#f� ���a��CE'��|�Y�E�b"f��|��\�D�a�a���ih�_�\T�"��!O-�,պ�jQ���pL8�	lr��R7I��n����"Aͤ��\<�i�c�JO���3v�ζ�&%���hқ~��<1�e�^a��"�ν�ҡt#��zs����&�<�<��mu��L�����؍ͩ�]��wu���J����v���*m=�J��*�J�N�w�b��*�Rn��qXD_aڗL�S�T�r�*f�{�us!�e*ޱ�t�ң��ϥG���m-�����;S����b�1t�Y��9�ǭ[9��L����ۣZ@�qS4T�E1ūrP�Q�\w�;zlL:<�S�dy�z���R��Bt�
b�n���7�K�����]-�bn3vEp�Zz*�S�GZ;E��(�<�lr�N����	�,�Yܭq쉭�&M{;)�Wn+�ZMn<��WA����ʝ��#O�@U>hMީc7�y�\YL%�i^�hl=����>B��S����h�R�E�Su�&�-��+��C'][z"-�1��Z̛�w�B��"R��*�0�b�Ŭ����'p$��n\�%�\��Z9p-��v�|5q�u37�MgF�09���)6�!iû�(�`V����.�q�	*H��eG�yXg7�ڡ!����p��Ts���樥P�b��>� ��>�(���Ё;��,l$�vB�-�r�$��f4h0�s���r�F((��wn#�����QFJ/1�%4o���"$��8bԈIz��$"`�2&̈�w1�����Bo�8��@wuIAA�Mr�DDw]�w\�;��.�E�M %y�=u�D���E�1�v�w9��oO+�4���Ѕ<�%�z�Ѥ�˦wk�]�N��犹�<����wv�]���F�S�[��v"����wt^+���p�@wq$\�+��n\�ℊ'�ĵݻ������0������W:E��K�v�]�ňM�-���k���u�m��z����o�������y(�qmv��+a2�'tL�:��l��|hb�71����w`�Vι�Ў渜�[���Ὑ"���^�/<���-�_����ק�x����\�+Ž{��cs}|W�u��������׿��羷�W�}o�}��:�-?z������ѹ�*�\�/����`���""�ˌ��ٛ���"��x����1o������������m������}_�F���u��c{k�w^E�|������u�o����_��ߋŽ{��/�x��������h ��>!u$��q�͵�k
}Db��������m�_>��~7���o���y���ssn����y�E�����|��~|�zW��_��zU��ƍ&�ܷ��xܽ���k����~+�����SJ�я\d���lw�o`pG�"��+�_����~j���oߟ>����Z~�>��_�x�j��ߞz�����M�}��}^��>�}��~-��m�{����x�[�������x��z_�w����E����j�������p���}�o���o_;om�����[����}W~��o?�ۛ���������/գ|k����W�_�j�h�_�}z؊��W����ͽ}����~�~�_��߫Ư�}�}������IrT=�lZ��5q���DHۿ���_������_���7��*��+˯����ۗ��+�ͼ^
����k��ϭ�w�ߞ�?z�7���|����׵�Z7����[~w[��7��}�����������vfV��e�'�czm��k�}����~/K������o�Ƽ_����y^��|k������^->u�x��6�_���x����o�w��7���ͻ���ME������^��'L}�#��m�2ϼt����
��'�����Ϻ�W��ƍ���/M�ۖ�/������^�����~/���Kw�[ڼo��W�_���/KF���x���_�A�=u��K��~z��z������}�Z��(�������և��2n���+y>���G�"�󹏨~��x�������z�������W������7�{m�~��ڽvޛ����׋}o-�]���o�~�n^7���om��1�>�DH� l?DhT���5���z���lE~/j��y��^�������>��>��x����7������[�~���h/���_�ϾW�x��u�߿~y_�|mͿ?��z_�ޞ7�n��+Ǎ�^��o�G�D�~�>����46��ݭ�Itac�Bq���z�7��wX=G��P<�L�|��j횵X�{y�6��I�V�I"sjV�2�]��օ��`�mƫ�;��������<����V9h�.���2*��YWr;�]+����P8]�t���r!̬���o`{����+�k�#���H���^����<���ߚ����ߋE�_�|�M��yھ�����ſW���7���������_�E{o�;�+Ư^���X�{m�mo��_��rտgh���}��#���8��B|����W�^u�o��6��������o��U�����签*�/��k�Ž��߱��C}�*�C�b#�d�~����F���x�B�U{G�>B"D} @"
ߪ�}�u����^/U�⯋��wy���x�_�yW���׍~�|�W���}m���/��ەz]��瞶��>���}�s�����>�#��J�+���׿~��~����w��[��<[�}��^O}k�ſ��z���Z7�_�Ƽ|W����������->v����>-��m��_��yc{��y���y��Z2|nz��"0G�,Ǡ���cv�/^jngm�������>����+�1\>������߾_�|W=��y�}��k��+������_�:�7���uz��x��*����w[��?���ܴW�u��W�6�}�zb(|�!�H���[Η`:���^�R]����ih���F�Dn��B4W����V�|k�m��������>����_}z��~7��y��߾}m���sr������-���u�zm�ϝoj�����_7��^4nm�w���������w��{Ԕ,���"GЇ�G��sB>�D��[���x���W����W/��W�ߞ�o��ޕ�W�߾z[ڹo���}��^��o��x���<�_���5��|��A���+�Gƾ���c��{n�O4W��}�?>�~{����_�O�������o�nU�μ�|noM�����|W{�����ͽ-�-��{��<�\�V���M�x�WϞ_��Z��^+����zTEp�s?X��i��#�/i٪c}Q!�꥿��O_����~�-��o��Ϋ���m����W�F�W��y�����������ۛ�z�y���}m��W����|W?�~|����Z-�\��>���~��\߷?W�I?}�B(G��s���}5Mv�g:���ϵ��wu�x�?���m�G��k����6�:���/�{h�^-��k�޼��������ս?���_�����>�m{��W���m߯^}c�
�>���
��X�� �eW�ND���[�]^�{s�[#��E�nz��ُ��̯Ehw-�a\��ۜ����o2nŶ�)ץ����֫��+p0�ܚ�� t#K8M��R��zc�cWka�����8ҭP��D��`��R\����@�;�Epi��ϻ��{�.m�箷����˛��*����}��zhߍ�_��_��~5��+���^+�������\����\����-�޿;���x������ �4Dh�.)-���[x]�c��}6�N�>��>�"=�YL}����>��UZ�}�x���ν-�������V�W����_�_��ۖ���o���z[������y�ž7��~^u�^���G�}�����C�f�7zG��o�pc_����=7־/��^/����z^��=_����|���{}[���/>��yh��;o=��}��|W��^�������{W��{��_���۽�_DH�}�G٣���?@]5��T�ժ>������^�������w��o����s�������v�^ץ�?����ۻ�����7��*����K{���}m�u����_��}k��y���~����>��W��b"D}��ޱ���j�/7����x�<k���ݳ���>/����W�����u��ͼ[���:�����~^������ǟ:����}W�~��_��﾿4nm�Ͽ�5���k�\>��}">b<"DG����=(e]�֗��=�����޵������+�����~o��_��oM�^5�_���\������?|�����W���~u�K��o���\�=�����_�~�����w�W�xF�}�Y]��aʇ�Zfwٜz;�����\�f�ۛ��w�~W��+�������?F��[����k�^���7��v�^��~^�x��x׏��yޖ�b"���ŧ��������������x���������{ײ��������{���羷�^-������_[x7�_���/�^._<~������oJ��~�:���[�����������76���K��U�|m��_1����r����쐝^,ѓ{P;�����[}������7��׋����|_�F�_�z��^/j��~����o�s�_�����^���k���~*���[��W���x����M�y��z��+�ͽ��b'�<]^8��]�u+o��DE�}�[�����F��~]�������p�]�ʹo���W���~���s{W������W�}^-?�������[�_��*�5�W5��}W�����_z�_���>���px�C(B��s&��m#�Q'�r�-޻��=��ւ�zl�\���������b�F_7�;5�з)lK[nR�2��ݔK�㲍�O~�V�*f۾s4�[���������Ⱥ_@��H��]�5b�7� H�m�Ik�ve7��/���|m�}��~+���������oʽz�Ͻ��s׾���6������x��w����׿[�����_~{����wε���ןV��k���k�w�k����V>��t_�7�D�~ͮ�5W�V�b}��~/j�Zz��}��7���(�/���k��{�����u�۾��+�����׶�����_��._[~��z�or�U����m���")���E=�o��w�f }"���/?ݷ��oM�wm������Z7��w^�ί��7��W��kžy��(��Z�������տ��hߗ��^��_��W�z��x7չ�k�{���_�O�\� �ەq>�>���G��K�|�D1}�~�������-���깹�}�U�_~��o��Ϳ�}���y濕�߭�_�����4nW��oK}^/��������ο�z��\������~+�_ȑ�ڢ�b�m���Z�����G��>�o�y�>z��k�\߿ݿ�i��|���~���o��}_�s\��6�����~+�����ϞW�~���[�]�ͽ/M����|]6�ܽy߭�-�]����<�I��i=.9Z:=�����o]|~-�]��_�����oo��_����}k��������Z�\A���q)�Q��Ҙ�&4ExP��M��D0�,a(����c�hNNqS�~�(2s�P�d1�:�p�d��_{ٶ�E䦹����:W�8i8+��z_�h	Q��b���N�-_ <	��ZfF+N�nQU&cn�4�L�'Xҏ���O,w�������I��v�s>�,�t�jC쮙2g�R$��|�.ͩ��n�J{m��]pc�r����������tW?�#^��umb�y�F<�&]��g���J������mK��� ����s�3X�Ӕ �0���S4Q�6��(K;����Aa���|g���3m���.b�Ǐ����0������]H*��:u�n�')	J���F�o�t�l���Ӵ�����܋7�Co������U��w��dqt�ƈa�ʄ�҆���p��N���`��X���G��q�T�f�BT�C��gQB��T��RY|cD1�:��m`�<]NX��W{Z�.�mu���t�3cg���Uc8���_9c���v��r4��������y�9}�&ʩ�R�
�ơA:2�ZH���N�#:"����5[9��7ىS�f�S�z����Sľ���6�UB(w?��i)�P���b��\�e0V���kU;�N���|���WF�Å=H���c%�8�����C_��&,�zd�<�'L,�7۞�zr��T�:��:�5�n��� p�c �UJL�J& ��z~�Wם��kI�c7z�;�3A��nK�p���5$u�L�-�Zf�p�$�8��Eq���N�c޵7E{��W�~Usq�9���Uv�����R��̚�-ˀv۽�7�/��!���gj\��lʹ7&p� '��1�xX��a4�e��"ǃ���*�����Wy�7�l�[�{�~~
�z��<���Bx�*��u=c{T©�8JyWC�29�R����5+x �+ܚ��p�Y$j� T�����-ӝqŖ����ow���U0$���+����*J�V�5z����7��9^Y���t��B��=p0��د����?x]��#�^/��#���]C�D-5����Uu|��+��B�[z���7����B��wo�*���5k�%�&+��6��I�X�t�:����'�����hK������་Q�<L��auEk������Y���)+{��d5R�������ɦ��}�[��V_�j��rp(I5�.U�)��d�f�|��8O	�2�R���t	��~Q�X-�^�nS+>����7t ��GO*��
�}b�}OȃΊ�*
�iG<rf4��'!s�>|�i�u]
.���,2w^Ow��]��mL����c+�@�HgUHnz�/_����>9�[�P�+}Js�28=�v0�ʕB���F>}�f	��ZM���E����P��g�OV�ZW��Qˆ.�>;��!��ق6��!5
d�����|JU��Ǒ�+Ry�x��q5��b~�j�r�_9���s���ͻ�-�(�W�R��t�C��� ����	S���D�z�5�̏����!.w S�g;GHP�Km"�gxu�-�"աY���t��Nc���z�J�K2��q�]�\��C5�Wo�t&J'���чՆ=�l�ז���MF�1��%X.�6u�օ�ob����Wt��CCG?�t�n�1��[�m�pb��2^D#Z|��"9�]�gR67�ԃ��V�a��e�5�j*�A՟	��=�}]Έw�1P�vd�'1�ch;�P�{��&-��-�'���/�@�#5�ǦyB��w�{��7Ǭ�!�j�qv7'��#f\B��	L��7݆�#�p�Ք��|{���.����^�2��x�.�9�v2�����B�����½�jj�/��b�X�F���)�2�(�Y�5��~�V���Ʀ�!������j�τ�xM��|���Tq���Z�xxjU��vú���7w��5�G몸�-��Aو��B��e��F5�m_��s�@�������3m�h���t��gF:	}旙�uMy�E�upt5ׅ?r�X9N�+*xFii�u!��v�ր:kV�`��*GEx[�V�M/
ky�*5����
x17i�jv���K&j���bC}Y1ߧ�VG�`�v���eG��R�X�E7B�3u�I�#��}���J���ئ�3zL=B�x���=��]Fev�dSPe^L������+�['c�+v��)N��o�f�YY���i�޾�����R�#m ��ݭ��bC2��kz�H��r5IKA��BDInd}|��Q2�jcª��Y�͞x�"j�	 ��m���wW܀����F	� ـ~�W�*e`24���һ����8�*l��~	˳�Ԗc^�=ꑷ���@�c��<��x1;3�����kt�o/���Ckf�q�m\U��{���c��7$GT<w#/�4���d�V����&椺ܾShތ�,���-�>B���\9K��?�͖�C���{(���9��deؼ}�0���0�?(�FĞ}4.�T1��2�g�ٿ5���,�W�Bd���Qsڴs��&{�/���+��	T���M�Wr���wR�|��:�*�sn�(_<{���M�?8���VC2�� E������*ʊ�][�"+f�0\k�/���ug��9e��e���\���Sr������K'���-�nl7��l�R���_3����e����1�����N�N}��M��*���x{.�\+@�Ŗ�n�� 4��of��~ut�\WS�x���*/+��c�EF�D��:��)�C�_#��ZRH�W��u���؆���u5#�.�4u�'2`�8��T/��-�"F߻]�i.xiw�w�.�Y�����7��Z&d�J��;[﭅9c�Յ�gWJ�M��3�	š�s"/�C�
���{�	X���`����P-������'DM_M��DD}������d�t�G	���0�ᓁ?��~Vtx���\��W��\�§���zꦍ���m�7�Sǭp8��vn3�|k�ßq�$�:�<-��+��p9w���S2�O�s����G��?��������ڞX�>%�Z<��v�M��b�w"8;↼9��1�r����rED<�J{b�1
��;"r�_M��]�$�h�W?����\u��������{e��C`5����.���;P���c{�����P$�4 �I��Է�ڋRk6� �u2�1q�0Q�P�5��8Ԗ_�gD<�{T��%�X����7Π��g\l@������H��f�t��EZ�#�s���uyJ�]_J��|��v�D��୤N�J H�W�v��js�FtEB�\8d:j�{c!��#E�\�&�}`pv�6��������C��P�ai4g�g)�P{s�.����/e���o�CW\�!�ۻ��9t��"�%�8���k�0Y���Di#bVӢ�nh��1�wL2���g77H��U���tO�v5��2����OIpݱN�JcAjĤ�ͬ��g5��j�il�{/c}�.�S�G��)E�H���_gpi)I��8g%Sb����k�j�m�|{CL�'�1��ɏ՝[�Ӌ�9��}U_U�"}�K��Ȫ�W��
��U��m�����q�s|�qq? Gx���� ��������	�w�2�ei�I��p��*ԦL����>f�TC��s��WP�*�a��7�˂W}E�
C��?/�{��pv_v��:�0�\�ɶ\�Ŕ�}Sof���s�vx�Gt��`�0�>|a�}��Ne���(xgr���ٲ�H�]�4��G�!R���U���x,\+ʘ]V'1ѿ�BC]>W^¾�=��vG|�ys�o/�'�d�NՏUB��T�^)�����ϸ�7��0��0{�Ř,1py����[����~驷��1�	�cVGI���(F-�IW�{P_��N��0e��e��|�w�WM�n�5�J�M�)�h�.�Xd��O2��|�"��m���Ӓte=�zب[�R͸�9$��	�qS/�.+�b���\t��0xn�ʖ����>�N�S�I��y��Q��`����:���Q���q���S	������:C}BӘ�S�	��� ^X���r��#NӴ�pDY(�U����,Ѱ�ߵu4dy�Tv���r�u�'FS��w]e��H 㴙�R4.'��(��}Vw�92MWQ�wy�YQL�P
*����x޼7��K�E�Ɣʒە������:Mګ2f�����s[G+5M�*]t��7u[�n��r�b.:
2ev�=|�+e�YR�lw:�R�(��zvf�-:滻����M��1�u%�ɽr���ͺ�IWi�绻Ұ1�G���Z�Z�����Xb�@��mGo)saI3k���d�B.��K�9�n2��Y{�ݶ�e3�&�s{ٸ9R5d�u�h|�n$�:
Z�s1-�wL�e���;�2qb�jU乲q�7M�gf�eTĴ�P^Rp� T�e]t�#7]�ʴ�d}���\
)�w�R���&�D�-U�sG�C��2�n.+J�`L�]����V�,fʕ�-!Օ�feZun�һnV֘)�V8�;]Iy@�銭�I��u���pXp�N���:�:i;��a`m�Dou�3�U����8a���F�4�oZ3��)�d���&��sXV.X�,e܎�PilႯ���`ӝ���Ը�ݸ(�dt�J�QQ�#�1�kue �YP+������Z�
�#�����X�6�7�WJ�Z�e�hc�<�k�x�i��j��{Fs��K��lk�Y��O�A`��&�ga�k����V������V�˙�w[к_rAy�I�*��h�������:�Ĥ��e��cp͍X+�x8(�0�μ��*�r�ۺzi^+�$�|a���y1�/���m���0���ł���r�u)F����a��/���XE�i`��=�.v��r��Aݓ�2�߰GH<�N�"�ٖ��13:D�4�	��V+1�W���d���!�k��9�N��������J�;0e�0�d��u�JS���5��8�;
�&��޺����ex0�{��c�1���cu�P�����1nZ
�['>[�����c�S��(�]���Ks��p�
��� �]�l2�Pk����q�v�ޱ*��>��Y{9.�o�(�Ot%�P,�ǈ\ۖ$¨�+����7Vk-lt�\O)Kbh�������`7�ă�,�ݤM�4i�a@����p�Z�Z;ԡe���$k%5�]d�3W�܊�0�\F[F�S�ZY�n�>:U�,�+ǃj\ha��b�a����9�#Y6�y��f�C�gͰ����5S�U��k���p5�yS�ٛM�e
��8S]�r��Z�3�F=�g�!�H��V��1I�AjN��Y�Ǌ9�9^ThŽ��d� Ř/Yg�h�|�K�f�q�W<���R�����F</U�4�zek�Ӭ�+GWU��f �,j���Wi����yEb�#��u�aml��f�f���]{B�$ns	���(�ȸ�λ��P�
����dF������$^u������j0���;�J2]�A�yƺ;�6���GKƮ0�ÝԚD�N�S EEΑ;��2`�.��ܝр���9&�]�I�iNr�$P����7/�&D7w2`Gws���wvv�n�C60BL�΃�q.��D�nphb��]+��t�ʼ��<]wq
u��̘�I�<�/:�!@�&�J\�)D���%�wWJM���'�ݎ���L���r�h�$`��sĲo;�s�5��wh9В" Js��ؘ��ME;�!�����t�W�
]����\��wsg����aA�DQyܨ��9FM�%�p���<��<��k+�
p]�t�dVm@��&BHԳfJ���L�x����ԙ
*�Yn>eo:�4�˅�����Z�9��#�� �x���kA�f|��:e|Vq��*<I��\�d$?�:�C<�/O���!����qY�f��+�l؃�&��Y�yT�κ�<p}^����������jx�P����:k1i۷���-'�7]�Z�q���;�n��^�#���S\@�������Э����S�)�nm,��)�^��~�4��}P���|�tCg�`-��;��� F-���{B�+��ܼ�$�Ճ�K�`5x�828�\@�2���&�nc�0ɶK�F�	�[���W ��7�rDnm#d��f`��;X0Č�(v���ZW9!��d�w*2k�A��8�-8����Q~�]Y��~����
���lF���=ߐ����SB&�����s+��d�6{��<l}��h��U����|{��2��2��g��b�{˯V�S�C�VX�ꘋ��3+"X�t׽t��MX�8�c|Y�U���(�n��\;�R� �%)b�E{,-s���IWˍƫ�;G����u�K�U�񍞩�l����H}.�.J}��V�=CF`&C[�?3�]��B�c���R�㸎cs1�{���E�D���M~�h�쾛������!.U��WHet�m�#qmO�1h�[�쭑4l_.t���*��̄�\���J�MT�׈3]՟�磌�y{d����vx\k�gf!����?kj�⩮e��F5����η��	>���ɻ^Ѯ�5��#�.�ь%�%���R�>�;(cj����`�S��K2�}ޕ�h���1Z����kSq��P!��p�$� ␏(���,��wK��Ε��7ʥ%qB�p�Z=��Xg8�.ʔn�>L����@l7����ʫ���u'�S<#��W�!�c.�o�������D���hf �}��5�=���ƽ�-�G=�˸�n{g��
T��CRY���k#��bC%ss�! z-ۖn�7�v�������0$Z١�y[Wq�{��;N7$G<u"�!�����sy�W�[�o�����d �}2�"v�����Ce2�d3�-��ة�f0�h�C��ʰ�;N%Ff�<�۾�4��R��Ѿ(?���u�}դ��$��q\�܄e�nx}��[/:a󚔶�]�3�9�}�"a=��T0�v!��~ګ/�W�;���"�믫@L��K4C��lYS�W�jkl�-EkLxQ�9�:�5O)uz�`Ӕx���֮���v,��`-�	 ��0��V�(�x�Әn>nfg=O$��]��d�u�c'�rU�Z�~�j�z���:p+ CyJv��>!�ѭ�lV���u�6��o������ʹ�����dA�T1��ɪd�fX�(��%:�"x�v��d-7�ED��y��}��5kz0�N7��\����\����Sr���ڱ��?t�z��i��Ҽۇ�eKI�[NUƱvXAh��j ����e�ruؼ���l!�Ȑ��1'�}1���n��!"�+ GGU�����Bx�oJg:�}�L<1i8�els��������[�x�2��6pEE�Ɍ�0���.t�#��ΏV��<�J��ׅW��h�@�n9��Z�/6Й���4�Xq�F����Ѷe#2�׵}r�Ŕ����t�18H+A�-�߯j��x.���!���ɬ,]�JVg��E��0��7U�*�W�S�Y��T>��mI�u)�LW]/8<&R���˵ĝ/�g���ҵE��=�}x�)��O����Pz)�K8�zs�!���ۆ�\�LvD�h�ɫ��\{S&,��z�\]&z�T��a���(�"�	\���jK:#!{ٷPxGp�:]h���u���S��U�n;�EWU�Aە%��a�~��qu�z��й�,%�5�[�Uw$�w��8!x�]԰����63�	����K�F�%/�(��4s�6*d�gy��G-����F�X�wx4��}�WՓdK�=y��{�6��&	@Gfr l�~�UX�;u��9c�k]�A�=�Ηn&�"�C8)��sB�%����F@0�-$<��/�������qC�m4��n���/N�7]���t���~\hqP�΂�i)��A��ɳeYy�OG��8�;ꤶ���6��.�1l�M6�@���Dc������N��S�=��׵s��x=J�Q���1P�
���T2[s��� h|j|�Y�<O�6���W�dk'{��{3E���֙�Ρ���A�'��p��"�Jdɸ���>f�U|v�5oSv�f{�,��O�돭}F^�C���a�׽A\B<ܨ��n�\�~�
����e��o�m-�8&��׶nznZh�����9�0-|��s/�&���7\;����Fy�ۇܐ�]3��y��'v����3z��d4�����I��5��=Wm�m���wh 㷪�fY�g�f/���3=��Q5a��'1Ѻ�G��~�o��
�%�4�B�`� v����՚��fo�t�y2�#KRw�Y��5Z�o�$務'6��6�z���2���/}I�.<���X�k��6q�!��-g0cZ:�4��G5�u9����v���J����Z�s���ő�'bq�c���_}UU�ٞ��g����_�1:�׮���4^��R�]tFHUӞ���j4�y\�t(�ʵ[�t�k�6hq쩸� �f��mPG�sj�����}����|c5��"�[�9H��c�{Wr$+�� ��
�U���L����T	�Z��p5���e�nS*cj���m<�ۏ�2vVK�Xx`����u�\¸?�J9�1�.��!}�^`�қ�k׬�W�;�t�#���`i�ڸ}�q�� P�|I���!!��R��t�'�2:}]�E	��	_n(Jԩ��T��m�>5���8e��P/��κ��C��_R��10g>��v��v�<���4!�p�}�k�r�459O��t�of�uHM)����-�,�s8���Sǯ���|4|%M��N�{�	�8�B��BN�,��P�k�m�npA�ꝵD��F�Ι�4 "T]ԁ�\OJ�c�f3A�]����8C�q��w
���������\MH���Lՠ~�MzR;}F����؜G���J�E��߳��.�����0Ґ:�w��)�M�s�w�0*Vj�G6����$�����y)���8�-���O8ܩ�i��EЎ�aܭ�J����ٚ��iQ��b�Γ�16�լ\�S\I�a�Żʆ[�Dm���=]n�X��j/�U��U|ͼ���	8�����b�b�����Y�O�P�1�u�Ǧy�jZvzu�@��8�p�Ω;��J�D6C�l�	q�p}_k�6��TN��>��=��Z68S��6wv�����_�
g��%�N1:��b��ىWR"��r����D��X9�˛%�CGZ�qN�73#�l�o6ձ ;'R��U0s��Е�o����Nw{�hn''��<a�*���*��T�d�4�m�WI�g���eGv���u7$
Ws؞t8���ɚ���×�_�Q?B|�����='�Xچ"��2��&c3qf&�ɞ&��W��:�<�O
�^���j�B^�>��*e�;�^͹3U�'��s]5�6�o�ۣ��6S;.t.fs�?�c\n�Z�?w�*>Ґ���Į���V*�yF����S�+n�v���|&ˇ�C����鹹��.O�?Q���6����Z�jY�T�`:��}�GG�BL��#ז��{cCn������`ƪz�_ �뙾Ud��Z�G��q-�*L��}s�Q����R� ����:��[��{D�w}�"�:r�C#%ufS�Q�oU&U)t;���@k���|$]t[�E��invP�GS�KY�����Ӹe�ElՊ���r�b��i�3Ov�G(_�">���k����W���ЌP���4N=}��Õ��vW���L��>nH���;���:�W]�vi_��F\�Seq� �P/%Q�|#Je�!�j�p�.�0��h�{y6��.5	�����x0I��Ԫ'\�2%��F���C��C�a�����I�C6���۫e�4y�=׼ώ|��^/�\��p�Gh��ڠ�tB��#lwE����z�N���̐k������Q�%,���`sϨ��&�Z8����.��*Rx�[�suu4��<;�9�it�ڿ�n��鎄�\��, �7,-���K'��ǧ�+��������K���^�M�,�	ilz�y��ԓٜ�˿�o�>��؊���s�v�.'y.�=F��mxK���:�o�.�}	�6.����aه�N+YSu:1�*r�O8��M���D��}�eFqb(7�Fr2pu�Mc??�����|��Ê�d����
懥��m;�Sx��t��
�q^\h	�B����pϕ���u�	�0kz�
�t[��,V��;z��\��X�Fk�d��W�����c�82 �Zm���P%n�J�;�ھ^7�����EXS?�����z�kf�s����Ǥ�Oww�Ch�ZE�:v.�����Lf2��(^���o�G�G�7�5Q}�,� z�o���ӿ�r�Υ_f����_��S����$��^�
�|���W���w_�����u��R�,�uP����gNӔ#�c�[���kp�n� @+]�W�!�lN����̷�>�����X����޻��]=1�v���f.Z�;"r�u�u�.Z�毥֭����a�	*���&uC�Q�7�`�_"�	\��膤��ƈc*WP۹�E�}�56V�ډU|U�65�@BI@H��f��G��U����}5�5��Ő���.k�7�PN$��#J����aQ$���b��T@^_�R�]���:�f���Z�c�bW2�Xp���p�ic[��^y��G���C��vPZM%<�:�k�I�חܞ�w���&�F+}p���S�Æc&�u�\<wF1��{�<t�Z���t���:tv�gk�_�T>B�/�U�m��� w�uٙ����8
��	���~��*�'��4v~�=����l����{\&��R�2[r��b��WQvJ��XY��i��v������@��F� ��2�D�hm��O�)��'<�Gx�\�K�V&�&[2�[�2n�\�Ј*���wfNn��^`+!��^�[��cU�KO��hq=]a?�Y�72_�c����W,�I�{�.�5��z�^�k�ﾪ�����k���c��)���u:���1�c�50��������ݮ:����k��91�|���.Y? =Q�V�jѿ1��(����b�Tk�����	�����u�F���̐���������N���j���W&L�7��Hk����}6��PT9g����ښ<���<�-g����c��xq���WR.�Q;�*h#\��K;J�K�!�>�����*cED̶O`�@	�Jȸ��H����&;���c���DP`	�:���ݠ��O�
x*�"ts��5�wN���h��v\@,2i��_l[��V_��
ovلF=D�omOop�Lz�b�|.�Q&�>�Z:�iz*�9�b�k���t�f.���9R"��m�ZK-!��$ߞЭ@�
�0|��˲�pUw�|e=��u�;�/�5*�OA�c1��s���U=���R�`3�ں�³��A��fQ\		MHbS����U]sI�;�U��qZ����m4c>}'[��p�S`\�j�訪�\���J��$W�Ϣn��ܣ���%�U�j68%�+3��3��Y�੖�����N�k��g��p�Y�����ʙWt;@��Ӧ��ga��lI��vV;oE���wdy��0��h_��6�}�ƚ_� S1�)L]w��ﾪ��o����ݭ(������T-}qN]GS����t���hZ��d�������Zxb�^���W`0�|9J����`O�ơo
��'I����9��[u�$�Wn�j�f��ŴoiQ"��'��N� �g�T��:7GJf��1�u�6�����xǰ%����ON�/5`��c�5�T9�H��`i�;X*%L1"�KhV�f!���`x:Җ{�w�O*�@"�Ԃ7DE�x�G#�4B_�C�ӫ�U��/ax,�'G���mk��❉�v���܋	��i�`<l}��ƁuZ�Lt1WKt�s���Cv2��r��2f>g���=>���OP�q�����щ�fVK�nb�GUԈ���*Q����7|�ξ���>�^(��һ�*�}�����@/�I�F6�M����Qߊ�e���F�4D�����7F,uO�m)�h���;j:�L�H��
�Dl/�G�{g���hK�^��O֍A7�a��e����8/湏E�upZ��T�W�lQ+��9����R%n՞{u�,�G] FU��󝱜�p-�9� �=7
�i���'��S���-��_I�b�p!�Ó{�hJ��v���V!;��ǃݚ)��<NGJl�y��1��^����U�l̘WRC`&q�+�Nj��h-T;2�^l��	}̬��k��L�٨b@��[%�͔Q�}ݑIuN�[7LmTpLU۷�0��H������[���ެkX4�c�Y���86\S��yaU�S]/8�搓�e�pu�T1蔃y�%{N;~�hۤ1�>�B1�ڌ��Gk*�:���G�H��Uz+�+Jc�\���n\�Kz��Z$j
�G�si��yq�q�ъ���Q�&��j���rX��1�7��43@[���v��Y���!�Ǳ��g+���<�wA6�_S$(pW�+U=�ܙW�%�VŜoE�����Gb��1b�6Fm��)Y�j��R8;N��z��'f�̸4$�:�����I)� sn&P��l��L�.�fԗ2=�qA�c�-%|�'wu,���k)Lw]L�
�BGl�*��n�+ģ��Pj�$H�`ѫ�WT�S8�Ù(�Ny���j�J�<�f�Y�a5�RK�g#�����2u�u�4o��3k(�4�}o�tC�v�.ޒ�y��Wil�t�ջS�uX��HQw��쑙��M���1���I�M�"l-����M�Q5Q[���(wV����fj�=euBQy��=��uǶ�K�I�$��ư*[����mP�7�ۙ���U͒��mo%���Y@����,��Rf�whCD�ˢ]�Ζ�f���d�R�VAYlyBn�j�۰�c��`�Ql!�>��U�+4�M�����J2��쭊c���)�5����΅�I��}��FֻrV��}��Bz�h��
�n��fI���j u>��*o2a�o�G�tW8�q�Q�ki�̻Yb9ϑK�7�ÍgM�p�J�c�+U�����>U�^M���a]���I�X���[n��dޫ"�m���*ܶs�z�f$���Vz�]�,�X���0�|�g.��V�7Z����4s����ز-�2��a���wq%4���݃���*u�71�h��q �laD̵$�&*Y��Cj\�ֲA�Y�F��5z��/0����D��ޝ�Hgv��ܹ��	�ע�r���8�6�zqݔ�VV	��?�	z��ݵ���hpS��k��?/s�s��WT�Z�5;���3�n˔���31C��d�uq4hv�õ�a}d�.HM�����w;�vQ
���n𬎥ҵs��:���[`�gb�Yo�w1Q���t �30�W6e8��!��.q�W���ܖbgyk2͇w(X�z����X7��wv�gh7������t1ɲ�i��bv����[3_W*#)u�tʶ1am8�\�4�{U��ч�*-�YG�;&�혙̃�"�U�¤�݌e"LE���&\.��DDh���wb��˜ut�]/y����.[�))�W�\�$�!�+9s6��r�y<n���J�# i<���N�<��ĢI2ɓ4�L�A�" ���9��,e�pE���G8N]��BF&l���5����S"&SH<v�R��]����I�&��B4\����u0h�L
dH���ɦ�)$�ݓ ��ɦ�r��wq	��4�2Q��y�����!�r�K)�HSH���I�N��nq"��p�ˡ%	��ۢD�,Q�	�"��]��rDwn�E1$�u@�R`�>�{��3{���9:hae.B��KC��K�@��ϻgC�L��.<`�r�X���:�1��n\��(�,�QW��}����|U�s�]e씴�E*h��y���1zp4!��u %��O����pL�k�[qs��6{}=��C���,GCr��\aY:�q�4j���⨨�[�|��T���m��g-�ޢ���;����	�2�{D=�����GGl�Ƹ@j�b�����9�p�K6��+=��^Ge�J6)l���gZ��m���{�#T�ʩ��^�C/F*�L�� >��<��_	-��![WfY��&�mx���ڥ'^z������}wH��=)�HK�DC/2.U��e�g�<7�;l�q=T�ȫ���}��NOY}3"��Q:�Y��(�U?*$LI��B�C��L��w����[��aw\��\n��C�����J�k�R�'�Rr	�j����ui��������P/jU��X��
���z�Ԓ�K�e��>�# ]�DR����
�a/v��w�td%��8�8�L�Js�ل6�j��s�c>MUɸ��Sr���ڱ����{�9�&@��tnU���e�3hŕ}���Vy$����C���%ׯQ~5zK%���>�TxoߝT��(ߋ�Q��<�a�\�D��\K��ql�K@J��δ��3��M$Ƹ��q��=�h��F�:�^w:}i�����#]iWx�j�Q���興���j��XU���8����Z|ǠpW\�Q�
�'w�"5:��!�Ž���B�T�I+}�p#� �J�F�*mp�C��&錞����)�����;1Q�.D\X���J�I�<�Lw#�!��*�j3MG`��PWJ�.�,�>���Ǹ�^ m���>��zw�l�N�`ԣ� ���n�og;�b�o*t� ]�B`W���v���Л�w�+�{}[��w8�@v��dg�ӿ�˦��R��M�{\/{jxݖJW~�w�V
�rZ��5Zy���8g���@��\nH��{�?/
��G�,Mi!��4ϟb�ֽ��QXg	4\�f�ʯ�L>448���/`���HÉj��Z�E�-�iI���A�^�ƁE�`�K~��S(��u�PBD�.V��RY|gD��+Awϓ�[Fl%��,�EX6��&O31�#�}���n��t\��M��6�{�ξ�"���#�s��g�ߜ��IF�����ai"��5;�1K-ԡ4�K{ ��:�o��s��#cs�ql���U���0�kl�?d4�\��A�ә���)���Z��4����tW�ڙw}6h�p2\�碅v�])3�Z7�l�&�P��t�M<�ې*�O�na��*�wq|�=W-��/\	ɝ'q�UU�W���w�=��u��K�*j��g4���q7��O���G���@�&�e�n�)n�;ie*.����b��\�&���&.����h��,�N���ۉH,����s�_`�a�D*�9�T>����b�|�F_*�MCn��� p�c ܚ&T�ɧFR서ܐ�L�,����ǧ�/k	�Q��\n{&��R�2X�74/Ҳ�[Ji�6'4=����Ւr���\)���ǝ4�}���^�Wϣ�ڍ>^�z��?D�]6vч	OȚ�r����l��a�@m#]�𺃕�0*�|��do�y�R�j���z^M�卉��,x:�/l��w��]3�ᪧ�?��W���?����p��C�/ܗ;��N#Kvx-� ��U\#,�3��3�r�^y�&�~f �cMK9�\'oNKv�X��.u�	)���@	�Jȸ�u�����q�j�E��ᘶ0uO>f�}�+Y�H�V��%p�UGK�Fx�>#��4��/�-��)�յ����*V[��G��M���=�Ǯ��3\����V� �&�_Si�H��s+N͖(�(��VpSB!�Y[B���hfS�mn�]�������-��1�OH7Lؕ͘��6�E�9\.r��艝g�p.kSH��oC�M��9������s�����tT��Ӽ�x�{��(�á3�\T�鋊�@�Z��傢�M��Υ���]n�QI\T*��t�V}M���^�U�0�$��¸:J9�}�QR!]��\���Y�9a�u1�_˺���r���0�m\>�3��P(G	�c��
�S�'"�e*^v����W
Z%=ܢ��s��ߨ�ˑ��>�#8��ժ���t>�ı�b����QfV옸۠*	��Y�5�
Z��Ӹ�����!��Cق6��!6/�/_;k���tʑ���. q������7��\^�	�8���~I�E��,��.���Jx��ֿ��t<�ʉ��E���$OB��
j�x�ME����
N�o���R��܈���u;U�V*ƓxL�W+�C��Tt��OTV3�SH����b�V�h�<:���7i��#��5&)4�ɴ�#]��+O���������k��	*���"���}����FVm��P���.9;��g��5������e�ц�a�g�"��'�l�lXIV��!M�pԁn-g.b͋��aVs��ړ�3�V��4��[<�%+GT`�M���3:=��nU=�͂�L���+��3H�o�-�V�R��p	n���L���u�;O��Y�w��}�}�}�ST�R�c�|>�a|5�w^}�lh�5e��*�"�:�Ȗ,5�0㶅A���]����x�D�3��b�t��.��*��������K2%LCG9�A�;��"r��ivt_W���m�ծ膾�z4�'���%������q�g8p �ȹ��H�ռߣђ�(3��ߛ���Y���y9ip��:���yE(��;}����0y�>e+�2b�8Ζ�"�&�yT��)^�AU׮��^傄������|�O%/&�k�G�w�c�վ��v��L�S�g�s�W˲�� F�A�3��b�Ǘy�O�2����th!�Z��[�
!�c�;������.O�Y�m�,f�,mA�ظ������)���os(�Q�~��xZ%����!�{�#hM.ǙR�1��zM�qr����s�yo��r�"�����cx��ڸ���=��L���Ul�{n�Q`�/���e�2��8�K�
S��)�!@C8����!����i�O����%��"�#�ۊ��_�j�WmB�k��j-��C�[�^�5����NR��Ĭb fs\%����;�a�>p�	'�uL��9�v\K��V���7���ȨK���,�E�Z��^���}\�A�L��q(�p�W�:�m���꯾��NwNr+���1�ΞG>�3"��Q;p�P|���"���A�1���xn�Nt���؞��v��id�}:>�O��1�VY�c%1?F*U\eI�1��X=2�6��<]�Œ�˞�[#�#.��D0��?T$����e��>dV ���)}�\]��w�@R��O��\>��R��Y�,����:B;�:Uro 0�`a}�Ճ�'�� w�G��y���n���>�C�{*����=�j��;���r*�غz�+�±m�Ώ#�G��;�=�fW�����~�BN_[�U{�1��'�����q��H���^2[��;��Rw��o;݊�2�s�ީ8���nZ���_+��Wk����sy_�g���}p�f�kם�9���M_���j����>�^�}[���$�%p1���L�*��Ķ��Wf���Vv��;����2�E���1Es��Me_YY���TN�j4��1�Oy���/���z����f�G������X�|o��/��k�u.S���:/E<e��;��R�.J�z��L�.�֗r���R���e���"��֥gɑ}&nw%/o����u]�tf	p�V�8��%Ԕ���N�K|�-��e���$�Q������興���[ȗu��Nz)���yԗ�:�*Z�\io-�o/���]��%�t�uZH3�i����t(9����D��{�eTɇ>�y=���pր�/�֞�uA��p�y�n�:���}��b]}6򔃳==��׭CzR���;؞5�\gS�r��Q�����`�0�A�c�������YV'�9�_u��l���C�sa�2�S�V瘻��u��:��H�+��i��No=�G-�4�2�;�q���æn~�"C(xypfg��H@Sl����Wmx�V�kxc����;�q�
�ް''o��3}<5�F�Q�WރhwX��n'V�پ��;�5E7g^���kY�Ρ9@�ݍw��F�#���<��̯��o(�Ď��+}���{������U��3M@��UF�7Z�H��1��e8Nf�U�;Œ�,_[�͞�{�I󜚳o�4D壟���\>��c!o�rWd�%f�q�T����j͹u��:FVsA������e���Ӆ��x7�R���z�鮣[�n6:d�!J��J�:Rk��������z�t���\�3������J^�bq�f���Uɗ87>;�o�G�����h��ۯ�/_ݪ+h�h���j�f޽ꌫ6�(����[j�AM�↡��k��ʉ)��Q�v$>l(���\���/tjf添��\$�PCy>
��e|]�޸�<uCQ�9lT5��&�M8������,���l���h9�:�K�P�+$W����F
^o
���u���zy���Ѩ�ZzP�>U'�����v^c���֎ȿFV�ן����[���On �T(w1o��.!�C|J/���o�.Y�~�眲�u-�)��Z�gφu<�
RA'l7h�)�:b��ӫ�&��ߨ���¢�Y�#����܅���x���%d.8��r�vT�_��P�Kgk�uB�P�J���8�TJŵ��i�T+�8�j���O	��E_V����2�]h�5^�����|#�5�.�o1�M��'�P1����̺���z��ӌ��3�@����qG�J�Z���`J�����g�m#����2u���ݫ:ۅ��U3�}�D[��N<$��j[��.<�2e�'��.4��=�y;�G���jS�٪�%��E�f�V�0���>�����%�=�V�1Y�Z�6v��nLc�M���{z�Uv8��ԟQI0zq��G"u��!�-m@w�j2��
�L�ȹ��\��{�7�Q���`϶z�[p3c�V�#X��5e�PWE�]�%vX��:��]K_o<��o���'��cj!���uM�oO'�1���u��d�j�f:�|V������/����ѷ��c�[¬K��Tz���������U79R{î b���^�����=0�y	Su�+������O_��L��nw����qU��o�2K���!�R��j�{+��p3Po�
Z{r����\�,�=m�	�[)̘��8���8˵׽nVBQ�T[aXJ�6�\��f�k3>|ލ�F@��xuY�R���N�5Ǘ/�{�%�K�Wq6^m]���m��d!�h �#�.'@��EӬ}o{*Q����ť�:��m(��B�Ɏ���	�{XJ��;n�
�f���Sz�N��0_4�Q��1͑v�(���W�U_m���Js�]K= ��D�ډ�e_��+��\=������d�xzӌ�����]��������D���K�T�j���އ�^�B�����X�VJڣ0����dJ'�*�I6,�3̲��s�:���J�:��Nw8��:�x�2�"}݅�-SY��7w�1I	r_4�LbW3u�58��֘���!�3�!Lt��h'�H�"�T��5W�Q��qz�8�R���6��j�e�v�0����H�v����ͷ�U�|�Ok]�jZ��9l���ڸ�n� �>�I&�2�]��0��n윆�I�i7FgT��	8r{s7�٫is�i�5i�-��yZ6��k��[jfN	<������@����'���[U�5�I�K}I�Ks�.����?FK�MB�V���ڮxn�X���f*����B��<��5��t���;j�v�4ۄəH�\Ј��ul��m9�g�M/���*��b�3��7��aL� ��[��e��9{��6�C�K���o-XV_/Vʓ[�]���y�}h��e�����6`b���c�]L:�$��;[]8s�7�!Bm�1�!}�P�n�0n<XI���r���`�A��hE��Ws����L��F�b<�J�qj����^k)nn�� �D�Uӕ&ŵ51�]PK���{M�|��msJcL�oOn���Cf��P�Ŝ;�]Y�70\u婌�|�GYJ�k��n+��f]�$�6��ۯ� �2�d�kWh�V�µΗt+�VN������\������m IŹ�Q�5�+u�5���M�)vZA@|�%�tE�p+�&N.�7;q�H�ф�ɳf50LR��l1��us��<�+3��V��+K��r@�Y���]@�򮝺G�VTZ;���t}O�s�$�$�^�稏	�+3a�G�������i�wboZ�F7�e�w26e�'7r����1t�M�r��n�kV�n���]Wy�P=�N�WfbQv���ŗ �1N��-�X5�	�tFk��eJ�H�����;�eI�|w�)����X!:l^�Ǽs���"4�bn��-�Z�<j�b�55�A�2krW͎[�V���Y���J'g�,�)�;�%e;�-�i
.(�/���\�r�WN�̡�+�a/�wi�t%a����alr=�anu>D��)ŭW9Ǝ��h	�]�;�n\Q����^*�d�7%����C�"�n��e�P�WzB�x%�d�wQAb��jt
��޼�@�`v�Z�ɽ�n�4p�ofޖ�k�n���K� ���v��!�.ٸ�9zT-�59¥
܃E��{�WM���%3Af�r��i�E� <�p=j�f��5���Cw�O@���woV*��,����&�/��Fp��}j4��]N���;cWژW����0����ѓK�{��B�<�}w�	�
ԣ�L:�p�b��U�]�7wa���j�;�Iұ�R5h$7�S�D�c���#0Q�pu�o4��/*&-�ꃰ�B^ ��[sm���˧��b�_`�Õb ��և�m�Sr���ټ�HAy�B�r���wY�@[˴�_q�Ӡ�'>����!���;a�=<���ť��5��ئf4\g��ʀ���NRr��RcHi[��Ʃ�-�]]*�-�������ʐ+x���#&kɱJ9GV݃nnW-vVT=>���$9�86e;�7'W4D���A���Ŭ벩��9��A�3+��	W�w6Ų�V����àfL��h+��LK���g��V�<��nh^E��U(<�ºoh��BFt�C��v0me�rN�S�5���kS�x�������۔�^���ܜЃ�9�V$�XN���^��]��S̓�� >� _   �I�n\�]'�Ԣ�2$�d�2�rb�@�bdRK��\�$̔&%��%4 -+�60��HB�",B2T��C$$�IR��!��uݒ�m�y�^v�$&L�k�����]$#&b4�F��ܢw\@�L�	�;�Xȃw]DC&��CQntI�P(�'94�+�������q$&k��c9��0�q�I�a�d�r�HX(ĝ��H�Hf��F�9F;��4�wgu]1$.�͹�L�ۍ 4���\���F$�Lɋ�3A1�1(SfNt�F�FI�ȅ��u�
�A�Fdafex�x�!�a�\���waH�b;��Icq�r����2b�E�f�ҡ��Y�E�����S;~�:I3v�x�n�l��2j]�6֫[��5({%Z�j��}�}���^rN3w�NX÷�q�g��r���L�Y�ET{�BN_[�I��:����㶟�WhowC�Ɲ��lg�/=���S{6Z2V�rNݭ��{�'��#]�gON:�J��1D�$ʞl)~��-�O����ƣA�b�ޞ����N\�8�'��uBWe������7�M4_=���q�s�e	�aK��S�="�u�QH��S ���u@T�R�-���7�/i:�y�c�[�rKL�	ܧ�n=�jtm�]��J~p\�xD�&��q�@22U��m�7ۣ�C���y�l�T(t�Ϥ�0;���#i�ʧ.les��3�!s6��D)}�ֵ����y�{���1���xr�c0U�Q�D���Z���_jת�B9�����I|�k����_<gYg>D(�i�����щ�՟n0���MN�{�#��o�I�l��c[{��Ya<h����b�	�o�ۿ�Vg��y)<�r�2��{� ���A�͌͠0x���|���fM��}���G�tx���� �󑠫���d<�c��wf��E�\Np黋��HG�:��OL|��ĥ�6�Չ7���e�wk�'O�}��Y��z�dު}ŗ\h���W���6��������`�Sp�$ӧ�IJ���=ck��`rѱ=�oO�.:_���ʏ��ͱd�8N�o;kk��9����k�n,�"���}������g���=�5o,�❜{�{|�m�p�D[p6���ʟg��ڨI�_Wt�W������ˢ�W��g�{�{V�){bq�f�X�re��$d��^�Fg����q�=T:���,�ڢkw)���|�9���vg��822�^b�0��ܪ&�+�)���c�!G�62%���x���vc\��^d�tS������X;�.xꆣr�ca&����o5�^^�p�҆gj�9�M����L��p�uTI}S������{�ϡ4�u�秕ԭc������m>���
�kC̗h�B����XX��u��nE�#�k78dM��R�wA;��鞕�o����R���ז���<�i�^Y]�0;�Ֆ7�N=ʱ�3Q�]\�y[���6��F���gK��s.8�>�ͭf�tw_f��LYQ�{���\�����v�7#9uoM�)X�T�k����է��i�j$u���!J,k��"�^Vcls{�p��#q'������5S�kZ��9��)A�산�WOk73GQj����ԕ7���X��B��Q_r�:�1�|K����)�&��]ē8l�#��0���u��o�I���u)O�˾L��M�����P홈D.���/�MO.ݎM�mK���j�Ht%�s"r��l���T�J;���
�6w���bzvcǼu^m��s��B}F�$�M�>�r']�1�l�Z	Jz�#�-Qr���\�!,�9�j�5�.�W�Ѵឆ��yU�rp���Un���T<:��F�=�����U��+g��׵m"��U���ۼ��!:Z�ƣVY�'\GU��ld�J�b6��b��:�VOmP��j�}������ ֟�����D�n�����R;u���{s���;�H\�v��b�N� ��_$�6`V��'b��Q�a�h�:�4����x�<9&[׏�r%���}��Yz�E<�NB�x�(�����y�#J�����ڋ�}��3�I�:�N��%C���i�7]�P]��؍��=����w�7���n�5�Z�BN���$�>Q�W�~��Ge?_v	��a�a���T+�h�Z޸ֻ��/��Cϛ������OUgaڊc���CʹTۊ޷P�V��]է���'��'�5c]+ا����O�_>��g��ZQ�\:nf�cy�S�8`�3��V_T�2�Z�c[�zˇ��i�#�����ެl�F�H���? >Udz��dG!����EY���9HqwW�թ'�3`����S������A������sڙ�Mm-���߷�:�Tn�^�$/[�q�s�Bﻳ��KE�M`�$NOjۋ�Ev'�^5z�N=�}jZV�kX�ਆ��r̢�t����싽�of�0�;mb����2�=��5l������;�}U�:y{ڶ����G�^�5������Wv�3o���a��iwGiХ�+k1#j{����ze�RJ��~�H���Rq�9X�[rw0�l�km�q`�gq��*'i�2�m�Dw˦��)�ʊ6�7Q.����v��6'�TZ.ͺ�}����u7�D��ͷ!ɷ�Wܝ|��IߒL;eƴ.1�r��y��t����̛$8��T]��=��յ���Tk�Nn�wr��+�~Oˎ����~������َ�E��Işj�n�\�3�y>�(�14�z8���;m�s�Y�E�φb����E�h���e,�X�hAhx��9��[�g3��z�f�r�t�ɖ�8H�1w���/��M�[\��۵��JC-k���&�����Ϳ��d���31A#Ld�[2K��,�q�����ʉ.X��
��R)-��vm�����= 7��{P[�w�ɕA�
g�ǫ��	_�e���=��)���$ܳ��皋�@��F��Gec�D?U������RR�0���.�B��qn�MH}�/�j�KO���@���ق��Ȅ�T�F��ű�s׎D��n�C�����Z�tK��9�L#���������b;g��<F�9#���*�
��ЦWfAd�L$U�ls�˸ྈq�C��q�$�0[a×��7�F�7FgH��g1ҖC /U�\���0�`�����2��kY�[#�j*Z�o꯳�t����71�Ѹ��km�{P�ٴ�P���p	n�hQ?z@�-�}Ng=3�g�>}�/tϷՑ׳�yw0�)�d��^��:wnL�錊V�x��-}̴�9�[��Y�#G��=�O�3*F�o�������w��[�Ri&_p�0e��7����^]����&f_g�T@>U@Z��mw&�|��.g�8;F.�gz$�N�am海K޽��,��bz�h��n?"��V8y�A�sR��듼�*5m0k��k@�k�&9�[��=�(ހ��O̳WZ�l��mmj�*��kڅ�j㓭�����ʭx5zڽ���ƃ[�V�~�{����Vq����H�x�kY�uF<�4j��9M5Tw214I�7�AN`f*�m�G�^��TV4���q	j�Syʚ�.�b�e墒y8Wr�d�Ƕ�īk��99��gE�������$
��.2��b/ �+W_N�lҫ&'.��%���������5�G� :+�Ӑ��ծ�b{�k�,X�+v5L������u�����u���ipPA��"xTɬ����{=�O�� e~��_v	��`>Us�Sp1D�bB�<���иG앮S��G��)�ƞ�'��,�[�j����鶽SG׿AK8�m^>żR�ٙ��Z[��E���Z��u��5|g�oZ>���X<*8����Iu�@��oR�l;[m>�i��og��U 4(k+
҆�8V��x��e8��S�ͽ����z�i����P��{�!�v�ь���mA��`K���!1��T��B��P�<���|/]��
��ޣ�½\{����4q�ڣi��0��Z#y��G:�Z�j��-�tt�jfi�Y�[�}��*,���7(��Ho�(H��~�W9��y:�45ONk����ܚ���Le�m�T;f~��dϭX�<�q��[x��Qk4�rM�;�)���2�O�m�j�����_G�_��:�.�����˹��u,�G�ޣ�$0g<��V<��:eN!��Q|ܩ5{�V�s=^��y>���iW����ܩ�{#XS>���Z���s���)k�f��d�Ò�BC�{��	ۙ��]WuAP܋�����Cn��-��E����2��t��ެ͟*of���\�O���&Bn5�9�ȞC]d&~9@���T����g�a�y]���U����Qi�4ہ��*;���r5+x���ʹ�Cv�ݡ���+�k��{{4�//�#�5_G�<粶���Js��/U�n��SD��ʄ���U��:��<���CV��i���s�����ӝ~n):�����u�7_w�`ub����Oxv; v��[��7;Z��wk��Ë��ng��ފ��5�o�W�3o���:�+�o�7�'������&㕌qщ���6/�i�]y�'��;�1�[�� ��[��]�o�UԞ��;�����\&�\�}potT�r�m�f�^VvY2�)���H<�OuDN�*�Z�q[ˇ�������0��{i�.eO	JٽU��@Dz�Nt�t�l��ϵ:��§e&��t��ɚ��e:�R|h�S�v5*�Ŭz���7b[cq�yf��DՊD;2�:�T��]u�F8��:�ǣ����븞uG�l	wE��wl8B�=�]�ܰ���
�[[�G���M�N�vY�s�U�/�a�ɛ}Я6�"o艹�z��qA��ö�qʅ)T
�>¾I�Ԓ[Y�p�ŮuV���Ia��i��%U7/��l����s�oa�3�S�wI�-��VmoY��@E�7�k���:�8�qTC��-&/ZL�����3�=!*�J	�1-�\�&ھ��S���-��QsW��a1q��{Y:��֜�)�p�gU�8�ꁶ;\����N� ����$�w�.5�X�UË���wq:�Q"=^�����=�:��k5gB��MQ)w�c�P]�7���1���k�fg�vF���he�K̩ȼ�8�o���	u���9��!?}����f�-�;m�s�Y�H����So3F:s4ā� X��r�Ǫt����U�'pT���kZ�ocͨUf��)�b���n���[O�]+GGf9�ڈ����Q1�;�S<�ȗ���͸�{Օgnי��e�O��n��_&�=�I��C���t�Xד�m���A�q=��)	R�K��h[�i+��Ͻ8�x���H�ۭ�i}�Vo��I�yMP�s{D�2�j��e�:S{���/t�}�s�u?�o��W��i�3yR�9O�|�.���ĵ?}Bi���t�Q�=��Q�%�2��$��5>��.Sk5<<���F���UEp�A�Q�'T%p6Z��6)�7�=Z�E����<�2���{��Zr�����ʾ����P-T�h%���I��{5rmV�����m�}KO����^[r�u	C��D�3��`�[�0�\�ɷ��<�����y�<���>��_�dJ��#+�l��S��Z�(8{���|i��KZ����<gyw?��'j��Z���L�'_֜����Cy,�s��އ-+g5�7�+�x�κ"���Ž����#%}�?@�O=����qKxf�$Ҹ�_l+ƶ���;.�3��5#��1-�H�"�T�D�ryvV�w'_C�6�/I�aM�_d���v:SfK��
�eƻC���nZ��Z�"㛏����S-��Z�W�^�E�s�L�PWT��؍oYf�W'��6P-P^�|)�������H��W����÷;N:fE��"�f�mY̩N�'�y� ��ܰ9�U��▫h�'�o3t��FA��۽�jB
��Z;DD���N�����������[O+E��(�����N�N6󤇲�wr5�Ƿ�ŋ��Z�r5������^��� 24�sh�f�d�w�f��YMM��xA�z�w2��QvrD9u�+7uYna�YU�\��3��̨r��Sf��H�����]"��*�ʵٯ�� #]�՝��ir��p'��l	GJ�v���Ds�K��0�a�7v໫4�p���Iܒ:��>���5����+ق���H\x��jb�ͳ�#��q3���QK��뱙�6��[3�p�e����T�l�ea5n�*�����o�Ω�s3�@�w2�*��R���n���;��ٸI��1mN�`��Γ�Ƨ#��F�����v�vfF嫶�����n�>[�o������P�C-�i��L+J�p���)C؏Qj��&舭J핻x������݉W�}3�%��������j;:�,v�b���p��fn��D�B��84�A��#vg�v3��]҇dc
qWdR彖���4/����S�D��u��r�:D_T���y⇌�|��ڰkr����}��o5�bLQ�U^�(Tػ��'qh��C�" ��B�u<1�|]Z�4%d�.iu�g��"$):�"�td�.��@����qâelx����n}н�Ej}�q{�}ǐFPӘz�Ia��n^��1�N�z���4����X+�a�[f��O�B{uD��Y�GC[�vd�kY�&TH佂�iB*���w�3�����R�:_�lG�S�
����
�ו���`5�&&�W<�� q֘�<%
�<��6��َ�!|��lS2Ҧf�2��9*��(L}Շ�����']t�!��EWv�8($����X�Έ��cM�CE�I�{�ӆ��+L��]v��tMt�Lj�l�}�d�5i��T��*;@��T;#%�eo39	k��7eK�x�֭u^��ݚ�`9��
��zn���vCq跩�R �!i�ML�r>n�}5'Z�v���8�N�$�3�:��	�&Y;�چ����������V�ݓ�@m��Gأ?GW���=xJ��[{�W�4irt� \ gi�7���R�n�Ys�R�i�7ٜ�i��ڣ��Ӄ4��
�t۲����ef�*l1e9��$���P�Kn泇Ν|�u�����(*�[f�]�0�}N�rw���i��P���WP��.LF�0]E[5J�\��;����I� �f(� ���p�{M19W���H��aRh�槺��8�uc�s�ٙ����I�$��Xq��v����ܦ+�*�P��2l�P�Ch��#�"JH��ш��~7X#,���iJLc3H��n6��B$D3$�s��0��&i��M"c4&"QX��"��]a��jI�*h�`���!$�P���n,�I%430$�W7%4�L �I	��d�L����L
��DPʔ�2P�QF�AcDQ�D��A	���d�#2D`�2#bA�T�(D`��q��̘�fh�:�AA#"�/�d1�,�S��LC$�J@���Ibl��Bf�T �|�&���9�'q�i�q��w���1�ZaG{�]�Q3�b/U�U�Y��8�f���0��n\	�c+{�;K����W��s^�7����θMQ�I�M��p��k�'�C�Z�t�ھ�_xU��'s��}ny�W�iuZ�N���j-�P�UF�7�/[�֧-��[�4y!����.�Z���e��Sѷ���=�){q�Ƶ�k���z��6�o��8�RN��;�sXv�?�m��X2����cN���p��SY<�G>뚾������V�ƽUL�[�"����V�*���꽝�2K'tw��-��]�{uޗ��_7=9:���a�O�`�t�T����^���Z�w+�,�y��cX�B���>���s6��o:ɇ[�5U�����NC�WrI�U��q+`*Z�\lS��_ͯ=>�z55��d�U��D�q9ՕɾqO&�]ׇ����u	��e�{�zv]=jOn�9����ǳ�7y��Fڠ�`t��;���_��E�*[(�z�{�{Dߘ	n���:��)��l�sb������Y>(]�c]ҾZ՜�\��:z+�s�ږP�u�Jnk���=�u�Xi���~���n^�&�c�Q�
�������:h�pQ�Q��26]h܃���f*�g{�88��)��6�n�.�g���wﾙ޵���[Q(סO*�˂�	h��5�A�"�9^>l�!�� Y>9��,�;9��]�*3�����JC▊��� �Sަ��c��/wy�9��;��{홄B���᠔��d뵼-!<�%�1�m�羹&}��*�[|�gw�9�	��v��-�y�u�84ٲ|�C�By�*qO��˘u	���q���tE�gIr����6�_]�|�<��b���?���q���[Q���tjӆi�r�Jm`�j-�a�_���b����!W�"����ʈ�Z�>�{_^ջ�)z��ԙ��%"�h��*a��'s��f�8d_<�b��}_IX2�S�P�Yq�mvjCwzd��.z�9߽�N��������U���/��-��u{��ZY�t�?�tM���)�l�y��q�{&�g1�r�W�VY=��+�R�~e��*�k��M�1�2������S��][�w)p%%.�]�N�CeoT�Q�5>/�.r��s�y��"�4�<"��dY��Ea�C�J�FGwV����voe�r�t��v�+�pr�N��t�L(�U�c�y�Gsn����SĦ��;Y�<B��u@��>lC��c�O)��'���)߇ֽ�nl��Z��c�|G�*JA��/>�uŖ�|_=�j�;����v�6^��<�7�oB�wh�$5a���l#�ٓo[ˇ�����4Lob����-\$\���|ocES�ETz���T�t��ϟ�",֋}u�no7����O0k�w"� ��q��JU���邾I���ȘΤR�[ޞ�='Nw�]��*7�y����P񜯜�0�S�w��c21�kj�ϋU�˻"��{�Þ}ojI��kX��m��r̢�F_���ۋhg,q�@rSq:��D"�=��\��L�
����t�Z�2�T�͙�o�i���Q|Yp9��6��56�j��|�Od��nu	�v���Ĝ���;�CtE�1�
�� �̸��{W����l󎏽C;0�#�ߟJ'ehq+�&��VuA]���{�cȻ48m\*9姪1�����1ǅ�˚P�W�@�X'cK��2T\TY���{��g;�\��c�Uk#"<�Z����:r9�[���R�̳J��~$�[��PՂ'��GggR��~��2v�S�j�l��n�q��q�ѝtEƱ�T�꪿Hgg�K͏�0�";'{��ܱN�fMc��o�N�,��7�\��k?}C1��duNpM���/m��Uvt�[�Ԇ��Q{I�R��q�g��uUOL\�j���,��W3�*'i��<��=]yb���Ss�y�QՍ;�3͂��7Y������%}�z2Q8��}���:{��}(��K�T�$���ͱ4fwm���g���^����;_W�u|U�:�%�Tꄮ�W
,�5Is��8}�y������ެrM���5kGg�.ѯ����\�L<����o+�]�U�z����->�{�(t�f
��|����w��NFr���j��B�SP�=|ǁcy�o�iT�~y�������s����U�D�ĝ�*�q-�e���k]�/]�h�t+i��%�Gh'4�ܽwpҎ#rm(�S��Xl��.+���� z�rQ����(wN�b�i��-}�J#VԹ�s�HU�ecG�Ś?��a�4kJ��2�<ܭ��^�U4u��w6���o����0,C��nu"�;���rS�e�)Ubݜ��o�f]��_50a�ފ��fB9�_k/�ō���[��R"y�~�3v�Ȱ~�{����}:����[�ji70R�lV�pl�zƪ�p[����C�T"�@K>�j'�m_���
±n�[c������j>M�w��p�A�,�h؞�ZhE�qX�Z���k{ճ��h+%����s�p��Qi0j!������F�#�3V��
:}����dvQ��N3^����Zp�Cn�7�Q��+�7�{�lӷcR*Gt���Z�	5_H�N�3���~}��s�^�<�Y:���M�L��Ag=����,wXo�&�Ԟ����v�^2�L�^:1����t�o��'U8J��Ǜ]Vn��ʃ4ߡw(��UΥ̙`�Ķ|�o���N�ڒ�ކ���=ꌱ��1�EZc�y�*�2��y^33Z�N*^,�
Kzu؇��5�,���`P�ǫ�x9d_f�!�6�:�
Y)p%�"���-�Ф��&�s�5{ �?��^O�U���!c��W{+{%��Ȯs�i���XV�AK�}����n;�OiXz�;{�"����h�9�JMwU�_{��
�6)�n�Z}q+sm=Ua���;��z'$w�˼O������r{*yC������C��\6��J�Y����h��/1=�nz�v��05uD��dq���_�CYqC�m=��e��U���	
�T1�?v����~�K�#���Ke�bkr�Q����#���t$m���2�,|��?���b�o5B���k�?=��:�&o{y��7=�����;!`��B�s T&wIt�|*On	6�{Y�������J�k��ڇl�B!qK�Sh�y�����k�{�w���z�N���K�6�6-��3�0�t���w���}�55Sc�xE깦�����4����I1I��p�|ev�w]%�i�[�6H$�퐪`�̸��q����6�����Ѷ�b�'��q��m���	١б)v�U�O�/�ml)P��]�	}$Ӓ-�ӧ��ˮ���5�7a)+�A�;�t�<�:����f$�W1�l�nq�� �A����fB�E������|��Ej�b��e�i���-��:����w��o�'�$�YDf~��-�)�L����}�_7�r�b�l���.�l��yhL�S��k���j�Ӌ�ʃ>�e�Iٟ-�?s�Cީ;-��;�D���5};����4����p\��I�Y��~��än�.��j�tZ�7	�Lz,��w\�ߞr�ж�����$��3͌�z����{��g*5�PVt��Q/����Rm���g*$�}cLv&+�6O:Wf�'�z���F�����:�o��r`{V��{�)R:������%��kp�d���uJ��"5v{a�l�� �=`�h�?��s��W[ɶ��s�(�_T`��kY�K�2��K�q{��U�.�W}~O>!�m;��R�0!H={d�gs�N�U�۽���C���Z���C�;��T�s,��e���߃Λ@=�9���.�|��=�lgTC�r�r�PS�}�Ld�{��ѹ(�C1�������>AV����[��>���Q�^�*z�w��Pn�E�y����i�N,�K]Ȼ��ոsEΗ�,�6�̠iwI�Jq����v*;�cceL����{��r7�<ny/1+����{\�=*�}��>Nem���b/U{��v��ZJ�v��m����=X�Ce��+`bŶ��x�q�#U�����Z٨�\�гFW˛V���!�c�Η=������n��۔E"���X�ϭ��(��\w'P�	�Z�r޾�ۖ�ǯ�T<�X���w�9��:��
���ݛ�Q|s������k���|��%F�e��31�Ș��0+r�����7̸�rV�%���+\����v������N���N�lm7�Z��F����n准�R����׎'�*'���n�[����$�Zϵ��w�h���g�����Pvz�g?�8��>��ˎ�X�D�ů��4��{)oR躾ӎ�JW�7�UG]�f�d�>��:��-�%�@b]Y>y��x�ϩ5�{�����f����x.)צ�kҙ�旔ogML^�
�wR�j����p�����6" �ј(�H.L������ 5:Ԩ����j�{1
�;||2.�ѓ4�j�c��{��N��l�͖Mg�2N�(�JH��⻉ָ(wR��ٕ��n�(\���oR3\�:�mDr��ݝ�ޞo�'o�n��)����w��s"�1��*b	zdcg�'�Unȥ6�t\�b�ow�^���n�����7�C�#�%Fc������yꜹ�,���*�H�j�ky�������7�n�P(p�ORCT��n�/)�Ę4����{�b3_wܩ��Ӕ�,kV�Χ��@��f����Uv��vrT��P�_'?~	h���X��Ǯ}�[y{cD�5��U�u���Qq`��:ȿ��߻� 9����^�[�eg�mD=��/O�����77ýy�ob��1��{� ��yvʺ�_K�8�������u���ᴟ3P��헮���R�l���M�ݮ�{�&��C7z�6Z��m������I0k��kB�]�?G!�	��}�窷��\��
���o[��ի����է�����a�f�ML�+m�!�vNY�4L�!K��>=a�tT@�'xj����`���J�l<(#�~��clgR� ���H���,9��=Ykv�;��}9B]E,�Q��'��X�ur�4e�����	����f�K
��2T)U^Ѿ���͸7�sd�!�s�c3�^eGV=��S��{	K��;���ژ�͒�z#=p;�1�6Z�%�7�A�V���;���o�2�*m1+L���a�ΚNu��z��tԾy��̨*�B�ܞcy;��������U�y���K����{�c'��τڴ�xe߳s��R'@�??Wv%��
���ቆ���k�[�p���:����>D���k��M��17�bh�Ƹ}�z- ���O�[�9#�큕��4m����w�d�|�*��Α���Oso.����z����ܻ1Wv�WGK��=A/���(�A������5��΄�}0���r�[/�C[�v�W���d�k�%�B���Z~�5�����m�]�>M[���t��z�q��y��e�B�︆�t}zV�y�?:Қ]-�Ĉ��7}k�[�<#qa���>�K/�t?N���V��N%�d�hT5�v�=��;{լ�E�!��Ӯ�'J�8r�Rtn��`�q�[��r�o,�w`�\�w��L�m��s�3�Lv����+:;��cq}��kC6F�5X��M��({��nP@.�&粔�_[�{[�o�`_w��lR]KN�ܳ��e-M��H�����.0tX� �s��X��'[��$�7s�Z3q8��Uc��K\����9v��hJR��n;�K���)j�1�1��8,]ܡ��l���7G����p�rC�t�r�C�,��]|^��c9V��װG�B��Y2�s!���Hդa����@�3hV7j�r��W��Z����GK�W��Ӱj��� ��\k(ے���Ï2��a�g����[�{H�i��Om�(�Ÿ��$�Yg�7�c;��~���]`�����r�G/���/�+�N�*�7�%7%_[@Li�^W/tot�ǽ��F����V�	�
C���kK���1�Α_c��X��9�S+U��QKcSE�U��zF7�3���t�"x��yԯN���M[�Q	��jo ��ѶJ��-��	��q-�˩v�H�kmu���e�;�� AI�����JR��ѭ�b��<�0���XzӉh[�M��ܙڕ�ol�A�v%
��Z�F��~[�{(��ss�{���Vƚ��T�	����+*�l��LM̰#j9�7wQ��bcHs��7���{�ev�t Ce�M�=��7�љhs�n������w�Rz7:��&��Q�6X�����ƹ�G�}��չ׺��hV��]`M	���'%�\��M�cU,�S������3�M�z1Q{�A�F�,@c}��2�(Z�5�t�=WE��6�����7��Y��H�θ�O'w��vte�A>��J���*�������~Ʊ�v];DH�J���=�+�\�Gm˜Nu(.n�u�[�gf_-��]�+�=+��9��ߍ�joh�*��=J�U.)r���ɱ�Xj�M9FXyW�'J��eqT���8�43V��x�vS��e����f��6�6�R��]�a,C�PE<C�g]jfrXf��m<�<�)c�r��| :��}3+N�YȜ���KNP��!JY��]{Ǟ��F���9\�\���.�d�h�n�!�yj�=DMd-�b��w�:��"q��#����t00�[��S:�-!mk1�\�qU�E�W+x�\�gq�3W0h���&���]�j訪XDp�;��[�f����;3���+�cQ�|ػ����"��s��Sz�vZ��G��i�]�}�N�Vr�u�釭�Z2�&�i�H�gt]�tGչ��;zܽ" �9��s������D��˒ȼ���%�k_DE���:��%N�eF�������gn+��c͓a!-$�f��y��P�	#�L�z�*2.WC4h4%L��V !H$�LHF Q�	�QDB0��(���� �c 
ƍ2��0^.R3��
K,�$��d0W.[��2�,F�1�0 h���Ja��\��6A6H�6,�P&M�d���)C�DL��Za��ę2���(Md�]ݱlQ��o"2X�
1Y)B��,@i"�E��Ԕ�ђ56�Q��TA�13b��� �>� P��^p�9_0�p|�]�w4����Ƴ��5�5�r�F��d�r��8^ف���8-K3��{OM�~��v��t�;�?¾���ݛS����S���&����cbz�D)���<�;9�n�ުxةT��A|f.�=����xeB\�|�8¶:�ȫV�k�S.�/����JM�:�ks��}u�k��u��}'~I1I��7VP;��*�>������Q"=U�
�߮a�v�~Y����N{�3�+�q��S�I�&c[���U}���:E�����6����u��Ѭz����Nm��!$�z�ޯ�ꓳ�]Ma�*r������i�v����c�6P������yp�ֵ�����(�}�w%z���J�l�̳��ZXtu㞞���*;M�M͂��7���bf 8?j}�.��N�p=��o��2:�9R\>���1���q-=��vhެ4�e������s3� �g�l��OF�Aw0�o�'T%{E�*!bXC��w�i�+��P4A��m\�\�5���JjK�1��mˮ��j���w�T���~줯 �f�c;o�_���W�;a��_��2���
���qou�"�S�u�ǐל��D9Γ��Ȑ{_�cs+���[�������UZN�'<��g�?��]Mh'�|C�Qaz��Y�|��������iwMM��	e�{_6�Y��:y `(0�}'��آ�f�?��װ3[�M��3�&��m�k睕�(���>���o_cm�E�WW�U=������6�>�r��Kkb��3��Oʂj���`�r��gl}r_9�i�|*�n��{�^�ݯ���-&/_7�+���0�Ѱw53�Q�`{�/�JPڱA�����T�є��l��Ȝ��skzwv������t8ő0��Gj�_!k9�q�nzW��Θ����9�4߱��M�/sx+�eƻ�r%Pxd�<���-�\�9p��Y��-�;}�^)��ݝi�5�4ۍw��6/ V�|��$�x4���L��/�סG=�eBھ���m�'�c�_k�u�w\eLT<��p�@��l�������1}�� gk�3�")�ld�/�E�S��w�,?Y�=F˾k�\��BS	�� ��ׁ�}4f���a�΄~��|fJ�kL��Q����j7���/���ܘ�Z�_Z��]C���2�k��)�a}�b)[�z6�5:���PԼ��q�f�X�Y�6����,ԗ�v�ތ�'\,�Z���T�c/�D�4�!L�/���n��	�|��	o��~w�3��L��3�]�W{&�*K}p1E�A8�a������>vo��)�z�s�=l��c��E:�W�Uy-�"����9͹���B���)��_m;����<�7�����7F��e_+޷+`*Z�^���o�Oz��P�@k4�lP�}sd3ȼ�u���3�[1�I�m���<)�[pm"�	�c'��(eF���`��?���N�zj���=�3�6S��m�`Y�͞��Iت���N����f��E{V��t������XyRf�|�z�;��NI��4?w�ϼl1l���W�A�Z������'�=W�P9�k @_t�g�oH
qe���(�����"�ɡJd�����#b��5���^>���y�7)�X�eX��co&���d�N��%�6\mS�p��.��7j�VI��ѷ�q1E��}�
s�7�;�w�Ohh�^���%�,X6�3W;��zM�|�~�u�-�m�T;fa��=�0��V�4�ڑQ�z*��J)v�_$�"���s4������D�C�܀y�`�E�M$339�	�����M]j��Yй�I����q����dm�й���cԭ�<��p+�@ۘ�ݘq���[P��_'F���m��#oow7sz�C��'�va����g��Ե���{V�)z�^jՂ��(We��ɞ<�Lq^��1Wz%��Z��%��T$�o�GK����7�������<(@[�d��ٿg!�t���Z��"�ν:U����,����㋱���c�'�0�6�}m���ٷg+��
�okl�Qery�z��9Xx�*\qщ�����B-�S�sЊ�+}��%"a�C�����Ӄ� ��I}S��r�ፊ���m=Q/�|.���:f����݇Kϸ�٣����9ϲ[>�ҕO.�2qXf�Nc�$6�.5۫�}��9Ae��>Sy��N�X:��z�r�)��׉%�'f>tȩ�� �U},֠9^RZ�\�̛�up�R�֔�d����e�yD��F�����!��##�Z�jG,{����v{3ry�']{��I������1O�:��t]B������P����s��J����H;���=��d8�w?�1O�$�I
�5����8���c:�,78��|��\#��>lg<f��(��w8���J�c3wt�y���O0<��ov�B���9�1�5�v��(Z�Xo�=��n��v��hv���鮧�q��K�_C/��q�l�ۄ�k�=�#�#3�Q|Yt8ڸ/\�].ٸ�N���:���I��FD�'�t�*6��Ð�q�l�
ڀ�`�̹�{W���<ko�t\�auҶ��S+���j!��!��^1�t��>��=�ݑy�Y�O�aY4ש<X���b��q�W��'[q��5��IeV�7�v�-u�u��]aVڭ�!��N_��'S�*���e*���˷�l�y����G<�r�c~�\���r�kv\�h��!�t��:���ͧ�t�L-��k�vgr��c�oT7e����謥W"q�ϳzYo�W }��㾁VhI;�˛���Β��XȥsV�gK���v4�1����Iky?eV���*^ZN5��C���k�H�1w�.����5V��]�������q}gz�~jQ��}= ~��sR�3����Ks�Y1_c�M�v|=���#gP��(�I��W6O�u]9�T�'+�iS�ժ���E1�@ؾ>,)R;E�^�ps�;�.���L1=��;��&�?=���Ւ��l9�y�QR�=ӛ����u�s�zh�[�_r�zˇ��Ĵ����@����+��nb^Mt��&��Lֿ��?a�e_�WG��g'��Z�<眶��U(w|�=�P�*&�[Z��;�7�5v���:},�����|/y�9QR�7�&�t�s]�t�j�O�jLoE|7��5�����M�^]^�W�U����������3�K���;��y�\�������>�|d��{��Ԥ�cO�E�r�H�*$�;N��=ٚ@h�7ψr�*�㩪GM�lG/�UhoC�I �U�q�Q�]p��C���`��-딭p�sS����3	���r�"�O�x�]��o.���-R&_�|0ɉg[�GXs���ؖ�w��q���t�"�W��CA��q�*n{y��]'���^�l��$j|�ˍw�)D�r?���$�y|�	dw�ܛ�3ԜK�D���m�4
�vDơ����I�.ok m��� �ճ��GE�ou�^oW�Wm]G\F���Ĳ-�����с�p���n�B���\<�wO�����7�6�+��zt_ԝq=�oS��u���~�ޗ��TI�M�.ܛ�~�FZ��x�<�6�M��	W��t��#�&��.�ϗ[ ^�ׂ��z��g罹�W	7w~�-&�O�jhf�g�FUԎ��F�Gګ��at��5З��~���s;��֐�4�x��&<�2K�"��-��m���օꝓ�s�P��&^��T)��*=I�����;�~ox��~P/���}����>:��s�����e�[��zt]�$�(zk� �MV{j�����2�b�:�p��a�q�x��Gšm����������e��Z1�;�S
��e�;�X���[[W�j��7b�(e#�R�R��/�w!�,���n�թ�ڟ�ÁWA7��n���{�ձ��N�Ň����OF��̣Nょm�)���U� ��x`m>9�t$��]�ԱH��n�vz�S)oW9�s;�S�� �t���S�^92��v��5�����3�{��e|�T<u����ؚ�UJzjq�~�;>(�x\�5�(����D��;))�^������GG���y���Qf5�7���zd�>k�t��S�w�P���Pf	-����b��m���0,��p���4�<��[to�=
v�=�O%{}R:�T�ә.P 7:}$O��p1ţ�5܄��$zh[���;/]�s�6ٙ�_ku�/�J��_3��)�Y�S6��$��;�G��C
����.�J�u�y
�:�xv�̿�ry����0����+ޘ�5�z~��vw�xF�ܬ����y֪ϡ�)��-�NV���Q���]ɋ�߬ɸ~�@�11�������XVs�EO<�8�E�8>����X���T�q+�༈ަ:ڻ��~��o������9�5h={�N:G�@5�Y����RGK%T�}p't¿�պn��弯Å�u��$:����7ui{��y�_$�3/>N��vg�#j���G����TܽO ���bEVr�Q��aLx����K��VFpu��^0�-��������Fc�sl1O`�Q�T��>� \���h�*L�2��݆lզ�`��8w�H�Y�L�n�d�ӽ:���y��f�^���^Ůg@'u�vp,y]|M�B��%�p�͏mU�S��>�lgު�i9�sS���_��8_��$���t��L�4}:�^W���/���%Ά�����詗ĳ�g�+WuC��u��S�L,߶V	��^��B�@����(�-��j����}��2º�����<�i`$5߁��:^>��f���,��Y�(��-��V�K�4�]�P� 7|3����~ =
':}ã�4g�����ܦ{'�l�|"�w���s����n�?v\�C��̣|�+��ֵG�.��t�~���{t\x7M=��Es;�G��TB����q��ࢉG!IU�p'��P��2�Y�˸���Uv<�����	_J��q^U֐��!��y#�D5�|�:g���l�<��KCu�O�_��0���n��@O_��٫��gyM��~Wq���q�Ln����N��3<���`{F�@��=�Q�W�m���W���V�cNh~K�V��͝�_K����|2qM���e��"p��}u�������=&1F��>jh*r�uC3���+#�W��G��ώzg|Kk�,���~i���t��F����/ڹpg��qJ�u�7i5���,�̵)���6KN��yU�����t��Rkk\!����ޤx�9Ǖʃx�M���T�m6&X�{l�*ֺRU3��������]N���f�ē��+	��,>ޅ���ݣ��_�̣���=1���}>��.Z�J��Ǔ�<�T�5������W����z��B3�w�#��@����z����\�K��9H�V�����1fL�8��W�B��m���z@�����}��Ջ��ԃQ
|J�p>7g��n���:L��M{7��!���},ޟ%>�yח!�]�ϵ��������or��7Ń�Yc�1���C���+�6�KV�u���U�?0�-���8bs��9c�����u,�p<�g����@��~ԥ�E��#?/�^Ώ]NQ�T��;�����G��^��+�̬�z�oz/$G��ܬ9���ߡ�q�M���*|n<Q;�fT	���Zn��Yi�������Ut�9Eno��g�h=�\�ɔ'؍��p�9�H^���v|J@ó�z��z��tx:�B���.=�އ�+3M'jd�y��T�<�Z'+�.ʑ�r�<jJ�2�џ#�z'jY�k�}�oyNy�8}ܮ���W��O���P���μNW`�*�K�%�����x��5Ӟ���K=�)Q�23{Ʋ�P�]�V,XSz�0�ٔ��6j���(��n{�	��sn�G܌� �3�k��0i]W!�t���I՚yU�(�X�c�����8zɀ�Nl7Ä(�m,N6v;0���wl��FŰ�2o^�ю����M��+0��4�#Y^S[����K/�i9�&o�w1�AS�ꗵer�\�zjEq/��-�
uIم�a�S�.PL>�8S�����Yj�w=���-�z,��u�gu*d�!̛���K����e���5��+JǑ�4���R����«oai�O"�h��	];[J�L;Y��zc��q�=�n�EA��nt�ؕem��7�+��	7(�2�:k��-m$�R*�3�s�_!��Pɤ[��L�2f�=�(w"vmX���88a=A�v��՞���9Jj:��u6f�_'Z��b(�(�:��@D����c]{z�ki�]Va��**����Y$KU,��� z<�Xx��e:�Z&V�Ϡ����n�5	����*Wƙ륶]�Ƭ��J52=���fGG���(�].�ɷ]��gGM� Gh5��p�8//9Dd�scNr�ﻴ���[.��� ��.�hu�v\��yd������L�el��9-+��aIb�˦k�|1�{C�VϤ��C�F�C.������"�<	_B�Bd��r��)��N�U��Si�j�kf��=�"�6���XfI��W�_�h�\�b�Yȯ�/I{m���t#'.�z��w�ὼ��O���t�n��
#H��Hv�J:��r�ֳ~֔����A��h��Vj�}[a�Z���r52A�\u���xI6���,�v��$�U��R�N�����˗h�9gwZfX�jd�ݘBݲi��.kYJ���Z�����ǥa�Zt���-����l�r�u�q2ոuP�I�qeC�r2�)y�(�e��8�/��w�d�W�zrJ
�*;��{����lQYf=a�p�rňKY4��E)Q��W�,L�l���(�lu���4��#]Y���l 5��'v
�z�ʽ�3,hR��)���!�$dӦju�����Z�Ԕ�5�w�V����/	�]r�L:
u�3]7x�l��8`s�@�\��4��>��wmԮ]��siź���c**G�F�ux��7w���YQ�r4p{2�}v+�UϢю�5�h;�J螠z���[ǥN�0ɳ�lA���wO֊h�����L�,֫���)ں�Њ�$x6[T���Ī=ۻ[����m��{d/k�G�QTļE`մ^�MB�:���hdP!�_ w	��L<[����/������LlV6g:%��X� �.�=ˈ�5�re�[*g*e)îӆ����Q[�/��������_�~��=��-���m��(��C�k�JS$�&D͏��FJ�r(�;�h�zr�$�Ѣ��,W��h؂6wt1b6,��I���]�Q1B%������	��(��\A��ʍF�e�nPs�e�5r��u�i"I1P��$Q�G��2����r�Thؓ#W7#d�1�I�.�\�G��)y�����^���Zf��Ѡ����d��ѝ���sL�Q2�Uˉ�I%cP빼p,sn��ɋ�+�+�p����N�A�wQ%��m:^.[�qF1�-˗-�Ȃ6��N�����<��wN1?�Z��L�⋥���؊��]2�|h�2�=U:��^k�}����:��s{.�U��b8Ԕ���"s1E��ͫ?�����,b˩�t�kN���r���kj;<+�dxW��F�0I�fL3��Y��x���!#9�x��>���_�
����������'F�N��;{��|lY�[�9(�c�c��|���Pd�}$\A�^s�΅q�h!���3ӽ~��!������W=@Z���}�7q<}.bu�,�" 7���䌜=����ͱ��0��yJ(���x��JWF�cЧ�����������s>�Pl��"e�z����k�æ�5�ө��݇;��סi�HTu�?+����� }�> o�5�T;�&j�s� �b���%��}�)%���K&��t�A���Tv�P���ǘSn}�w&}8�'p�9���u�r][��ej��h�|���S�:'WW��ܞ��51���Ϋ_˜K"��P�**1���5�;{�®h��Pp��G��s�y�����ZN��������%y׻#>���y�6�zZ�|'ǹ5�N�п@W�灇��p��<Nc��w�B�;�����փ���*/|��b䊏1�;c�(Q�P�j��\�P��#H�����x,Ċكn(35���B�l���ƾ�er���j.��]�b�39���3��+X��GV_Y�ۏPz]!l9�ۍ�|&���ו���+�V�{gp­��L��8�V�SQ�ө��@�-r_l�s�!pG�>�<��*�>��O �|u���c����'�Z�2b��6�r�Qv�j��Fw+"��<ܙs�{��pX�օƩDeQ`o�A=b`��C��O�؅8��K3��X�v�q�G���0��W��C�<T�9����B�s��(��Eq f#�mA���m~Y�V��@�c.�{LWӎ|�f}���a���cK釛 �
my&�fW[���vA�<H+�P
G�J��г*Y�v��[^�C��?u�F��l�s�[+j%8Y�3�ñr|jd��"@Ғ��z�'��_	���S��:=^��Ӗvw2=��(%�+T�=�m!:\����H�Tf	��q7�x��j5��7�D�t���	�%s7�*����=��RM���H��S_9�� s��D�u�ؓs�ߵS��[���V�'�����ap�y��U��\2V�߆}����ә%�$�W��tGdO���xӐzwc�9~��<�{#Ca��p�i�M��1l��w�W�?q�����Ƿ�gٛ&��$F��8]i�6t�����mc@r�"�U�Z<��Z��_m=7�8��\�>C����P���ר�EJ��5&k^E�5��H2\4oU�.��4$�F�P�r�k1
�֬.w_a<N�Щv���L�Ǻ���U�V���)���¦�Ч�fc�t��S�4//Ը�|�>-zH�~Wrb��2o�������EW�����k�|��z!T�0���z�L�Z2�׸�oSp��2!?]�����0��s׻�S<��2��|��,w�d���쯼R�.R���se�z�МZ���{1���v6���z�|r5���:�ٟ-���x>�b�j�ey��Z�3orX`��f����(����n3�߆:����7Q�Ns��ׯs��+���X8s~�xI~\��L;�O����w��zgED��,#������c�؞-����7\��Y+�q���)����y�x*����~�3��S�:$�G���e����7�K�����~+)���Ը��)f�[��ļA�~�1�[S�qQ)\�ʈx�u3�n+�\w��C}^_�z�7o����S3��SK��'|ZB�ӳ���D����T�P5���� H��(C&��&~8������qwUM�=�B[;��#�q�[�NOp.J4�$�3��reP�&�U2������j��Loq_�}�l��[�Lc~K�u����|	ۨ���-�$I�Nݣ����
����7�*�?/E��]��C���R��xƌ�˷�R�y���k��0'�L��DfL�3Wz�Y1t��:qѤ�<��"�۸j.ћڤo7(L��@�6�uQ.��>!�Ǆy��{UH�uL;�l�P��5X&抿\.
�o2=��������u�>����ܺ���kd!�ӣ���W�H,��>��(_NpXi�{cu\xa�D�"~�T��>�c�Σo�!�}M�zVSࡓ�
��Pq	d���y����n��U�&G�S'M:��c�����n��l3>��+#�W��Dz|���GaZĸz}S`�x��c {֪&��'�L���/��r�[5�%Lz�����*.Zqjz]����s�F��G�z�/#�|{��*��R��C�=s/�t�}[+Ǭg��m���W-{�;���==ݕ��?:�8� z}�`ihd�ד ��>%P8���^����g����Μ���ϙ�;���ˇ�C~���@zNz�o��X��f��
8YEO��60�s��%۽�9��@������6�W��;����w,ϰ�C~����*�~��muӅ�n�a�x��#w{��Ѓ�{�>�·qS�t\T��;�����Ꭹ{<׫�F0}�!!�����dgY�VQZ:p��Yr��j��w����-���8'.ЈUr�7�ȥ�J����s�K'�����:��w=��%͛ob��/FH��'Ru�V�Bi{���GBq=�,d�V�ʴ�o+��Xo�Gv���S=
��x�Q�m�N�<Nf��yB|��Zn*]��-v�d-l��mgo$���XzX,��w�O"���K���L<�U#q\��\tHQMQվY�j�O+�1�����l�s��c��z��F���*F�\�O��ASzN�P���g'�o/i=�t(���TuǱ�B��V򣞛�����=����X$�~�}�\
{���✚ݯ`���%���]K.�Эi߸��R|_�I��j�z��-w�����C+F*�O�UP����c]o�}��!W�Z�S����^��Kd/	�k'n�s��?���KMs���@�F�>-��A�^s�΄�ԇ��-���o+�Fb��[�n����A�N�Q4̖i����+��g�Gڙ�׭3�,Ѯ�f��d$�.ɖEDws�e΀�+�
m�{��Pf8�NǇ��G�A� �(����r���ZRQOxu=u�}{�_om2)�;�����ցP�,� ��${����E�����M:�C��V�䉳F`7o�"�ٮc��D;|����,�%�*� �h�l�c�w���ǎ����'�f���ԗ��92o��+8[��Ҕ�h�Y��|�%��sT�w*Pl�5�ё�'��])�o��4c��ErBQ���c�*���s�2���7���q������*!�P�f�W���2jov�61d��dd�9-v��Gч���\��V�����|n��y	��dk�W��g��J@��y(�]v��v7.�����HǉT2c��ևu>Ӣ�:�{zX��U�y׻!TqՁ��ӯ)b�G�!R�9Ħ��}��.�N��3�'tú����փ�����'�G��+�o���Y�yf��8ٝ����s�v�>�21�������Nc�u�Uܫ�D��z'���9�9J��gnz�k�K6���^�*@
���dZ����:�]8ۮ	{i�vO\\��6�^�|c��v�{g�n�	���GG���Ǻ���)��*u�\Kڅ��o�/��~y`��s٨�}Ű�^���^ʒ^�9�Îv9�u�r�)�4/��cn_T=���u�)^���~�W+�p��=�o�����& ��J��2��v��\5����=,e��h�
*�]����t��Y�K��o��0�G�%���#N�Jr>^j��_�M;�S�iA�̳���~V�Y�.Zs����أ5�nn �0�����ƖL'xv#��$�p��������N���Y:Ϗ��׆���[���ul���Z�!cB=alz�U �22o�̺MWi�wf� ���E4q.����*u3��	��(J�7�=�SelyQү�m!:\���.K([a���A�^/g�B�Av�m*]��{1i�N��u����#��!��{}R:�T��9��D ����E&�N��d��>WY�K��#�؁ꅢ�7�
��u�.!��69+��+�Ȇm�1ā�9&��:��.��{~z��䉈�t�\R�#÷���G�
��U�;�e�0-����y�'ˢw���w'��s�3�:�T�{ƅ�[�ƒ��5�#���L[o�d�s�5�>�o�z���X���zu�
'�]���z�d��>�-m�Ȋ�^�y�LsUV��� �3�o��WM��Gr��o�z|��{4X��ԃQ>%Pɇ�␍��)��x�Z>�(�������o�S�/8̫���2�_˜����x!��a��u��r���.�{���7_��rZA�JS����X��+��ğ��iFT�Ayys��i�;Y��?�W-�.n�u-��t��+�l��$���#�������c�<��Fm��������x��_�4��������&W-Lz���fŜJ���Q.�Q.�wӹ�.��'A4�*g:�i�ۜA���
�5s���U�!Q��4���frA��9=�VK�>�P9l�w��K �&�ZQ�N�t�w}�7+(c�9��ܣ�,Sc�R���{�Z?w#�m(1������趼��Y��`(�^����g��z�+6��'3�����^��낶�XX���2��,I>G~�tx;�a��|���>���^�5ܴ�(_��yW�Y^�<����Lk��g�GEW�W?��q�-�W�5+��%m���Ss�!{�����w#�D{�޶=�''��rQA�V�A1����5^fN�瘖iVw�П]T��j:z��|W|�G�
kd�o�Tðl�J@R_�(\���[����F{v}�xg����g���j9���]n���Ln���:>U�3�����/yݝE�.Rս2��W�,�A,��q>�p7�����s��R��^��dG�z�ω�2>ӣ'�T^+�3���g~�3���)?F�A��Q*����B�g��J��E�Oz�ԕ0��Ch����k��,�o��L��&2�1*�'��^��c��z���]5�BTǽ}�>c�{7<�.��v�T�Բ_�g�w���*���K'�����TT���3c�߿A��$w���yOhlV���7T;2WZ�0m#.T���k'�WH�PC����M���ߤ%O�Á�L�&�u�����f/y�nT#��|�t�/�4Zn����X���<��&���\���c$����+��d[����ewiJ��7js�W5�&�+�����ײ�C󫓏��{��8�ڱ�ɐv��@�|eŹy�^���ћw':|��ӨT*9��_f���򮣭�]�����s�0s[ܱ����_f2=:z5o�H�H:}�C�gB��cn'g�1ו��<e���q�X�'�9�&��T��brk;]��~�Ӈ��j�����_�E_�`W�a���]L
����ȇT���~�d�z5`g'۫�$N���Ozk�.1�h��W%
��Z;�>E����u.���8<���pS˥V�z�I>S�;���<�\OJ�!��յ<o�>% a��3�}2�o��]���E���{i���}2!z g��p�y��Sy^�<�᰻*F�\�O���h�f���x���w��J��Pq��P�����vuTu��.����\?)Ȋ��9\���zn�ү:�{�;y����Nz&P�N��L�K��Ԟ��^��;z�zC��-kjh�a�2�gP۾��d�e�`�p@^�,	
W���l����|s��B�>�0s}�h�H�?A��G.���v��?��T�GQ,�h���>�R�!"M 3�p	R���zv�������y�<l� 
�-��f^�mT�5]���56�X#�����{Jj9�1��M48�X�X�v���ι\tÊ"��I5ց����Jʑ@��y��ۏU3�%� ��ž�.J�ߙ�	��SK��lu`��^��"��ѿX�V�l{Ը�i��}�?h�{�|p'\�ţ�e���n����id�+=��G
�����˝�0W��nsޯ���1�}2��ٿ�I�2=�{+���yWod9�e\v�s����V��"�r��G�x��k@��t��,�#6��ͻ��y�Wgդq��U��%x�J_��mǱ��ɸ�/���� o�3Tr�qBzv��y�Qf���̔a"΍�s��ZpN=�_F�>7^\<��wƗ�Q�G��V)������B��U���JT)���Q�����������vl~��x?	�ɐ��������]�<��g��H�+��U�E�W3gC'3��/P���+�d��rM(V�e��^@�_n�ڻ|�}@Go+c�>��zy��gփǓ��W'�Zx���tm4���b�9��j݉ܔ�=��I�B> Zj�p�y�9�:�]8ۮ�нS�z�|JQ<!�uE��)�����j�ʱ��r��0>:H��k:�҂ӯ /w�C� �A����؍�z�������.�˦ʷ\{F��/.w@����[�@���ʵ��oS�3l|��f�S����Y���.�`�c��Z�(�K��g'/�������[�T>����b��T��U1H�^8���\v��ZH������W"���6t��c���JC�],�>���\;�f�`�͎��^p�Ub����]Žz����|v=W�Z<��J:��*�smc��s2H�\��K 43;n��D���G����	O+���sj��(؟u�Z�u:�89��j�M*�d�����ޱ�l��G.�ksW�mG$�Y<�O+�-�C�D\��֧>�Ɂ��*��9)�K��UX/f�Iv;���
�-��p)��g[�"ӭV��'^ӂ�]a��,g�pw^��c��o(C�ru�a��W��繇S�\�̖n Hޭ�e����x�"�	�'ayZ^�bu��t�q_ b�{N] �pÀ��2���j��F}ic�jstB�h��kq
���t'bmu�\e�Ѭ&'���t�ή�W��j,��>[�^��'sQ�ɮt�����$(NSz�����bg�9Ք���m���ڈg��V������<VQ��o�mh��EJ[��7�:6�K.�5�)tWK��4�F���}w6L�s��^KH����f��{�4�VT�h���h�b��Pǝ�ձ'���buv��"��qܕa)�P�:�Nb��Yu�'�ë�
?uvH�1$e(��]3&�-��ۂ��c��a�hiʝ��]*�e�1jӽw�R��M-�,U+;#ͻ�m�"�*��A�P�+)ޢ@ט�*���_SU�x�����ۣB�����N.�ZȈ��wN�̛�ʝ����ŕ�Z"v��f��aV�O���{����'�%�M�x�T;[�+�ۼ�T�c����t%�ţ84�Kq�+p���T�T)�O'��F�'!є35;Xhk#�$����A�-%��yC5Q����4�讳�^�Z�q��TOD�*��Z����y.G���qtnFw:�*�$}�h#��:�e��'���PR�����^��FnN�uԎ��ݒm�a�6.�d2��(
�CM�_:�S��N��9I�5��3��n���u��!�1Qв8�IԺ��5�s�3tu���T�TN�=3k�Q�q��z`�ɿ�,�A�l�(��)P�!���rI� zq�1��om	R�u�t
l&3W��닩�}���s(��VK��I�*�7&f���?`��_�yY�Y %_D�Aκ��9�V:^�c3����ԟ5��ůW]ϴ3R�"�'6�'M��<�'�"�F9eл���}��KW5\�b@�,pںc)}+��c����]��#Y6nLRРhY@38�,0]w�+�*j&й��g}6rf�NN�����0��#�*;q��Ӛw7�c�  +� �_P�w�9\��t��]$��F���o;�d����6��\�&����IW7+�ȍ]ݴI�]�sh��E���]݋�����w�E;�sUͨ�$ۚR2湃E�nr�E��EȊɌ�Iz�;��(�m˻�;�l�ě3N�cs��ݦ��"���F��i.WM<둼UȠ�b����%Η-�w+�K�we��<�\ܓ]�ח<�h�Q�%��4Xƣ��N�;�9\��5��v<wG[��\��\�����*�q6�9�wuI�����.W-r��m�9�9��q�￿-^�L��jW+:G��cD���UY�W��������ѝ;��+t��q�ʹ+�v��&1�8���GuXҵw_-�V=?�˨W�H�@�*��r���Xx��Q�uĽ�YmV������)�����Wl���� �'C�<=u3�1W:;�Xy���o�m��?9ފwT���o7|��뇞��q��>7��� y:�R��Y�,���X�k���_'�]����j�q��V#������}�;�p7���F�P,��vRS��Q>��\��{X�2wR���7>�#�z�y��̯)8yG���7�P�\�k�D a��-�'֗��V�mffv��,�Z�L-���i���_/F/���Pӓ쨇3�k�2\� �l�;;��Fx����jg��i����w��5|�F�����X	���M��z��`�lD�xT�{�����%�u�&[�*�SG���y����%��l���)��czٹ�n�t�y�M�����Ƹ��Q�Ǟ|:�TD��n��J��$y?+�1G���~������{��n�c�baD�v���ex�2�ތ�u�7���K�}*-?��ٽfIQ�A��}9+����u���^�jzf��T�[(�&lӺ�**��m���mYJ9�����V��d���r��Җ,]Ⱦ���WS�}�W^�طb$����og��/pr��c=�3�ǊY��}P�����Ĕ�r�;F�V�v�#s�O�!��܋�=��������E���ԃ_GO�U�}bwL)��JlT�.�(^��t��j�t��u1�ѝy~�W����C�^}����6���D���G�S�~�2�n+�k'2�X=In;�S���ϴ�8�}�q�n���	�n����wPz�^��\䜑E:�R�={�����<_�e�:W�M̡�sF}�G�5>�vxΰ�R�cm���9�Y�3r�)ά�E�D�,��ɖ-�:v�|2�<�O�踩t<��F��=��/k���L�M�.�ե��;�ע���O�g�Z���05tc ,I>Fu�e1ޫ��z��}�<u��on���mT��
�܏z���s�{p���'B����c��v{�2���du�z�O�����y����?F�e���=�ף=�}��#ڽ�c�rrx+�%%l�ދ�J������%<b��%4\s��v��3���j:z��nu���q������w �+�s���w7���fҿ 2��%09R�t�^|�k�GKى�r�t\q)���1ۓ�p�爀}:�fo��G����z&�dd�	4w2  �:
�b��w6�w��l@.��b4�r����
�,�98 ˝�ݥ9!�t�,.ԫ)gmNU�7>}x���\@��V����J��#����'];�t���4�+�\v��v����&!��a��P��]1�p7��~,n�:��>T�dt��l����z8Ԉ�{.E�,L�vÅ��x�sw��fE9�ʓ�I%yMV�x���=�������{Mz����W}-]�X��z�>�����1�7��I��e��*��e����3yk����k���:��*����-~�h�{�+�ۯ���f�@��Ol!���]iع&|��Xw:w��s���z��o潷�����?P�z��1�A���S�Vh���Q,[{�,�ف�^8ߝK��*;��,��/&�;�̡i�O����o.�r߅�R��^go�@�Uϲfw�
tk��N�wՕᲥ�b��^OL=��_��'�ݐ��*'�.���f�'��*����^��S3e�Q3���·qS�tIS���]L
������N`L�ӽ�!��gm�}J���c{�Z�(�ʝ(2s7�0��."�kMԺ�b�c{��ڏ1:o1�Sع]�����dz=k��r"�Oǲ�!�s����j���07h� ��>��X�c�7u��rw\�۟�f����?.Fb%CpiXDʗ._�6�2�՗NUM����ڹ�K�Bu�^V=�Xqa�ey�E�R�{�9������xy�����G1�+"3�w^�D:�&���=oQ䮉�Y�E�;k\e�U����mvƶ	P�I���y���؀��Ԅ(�臇Z�q~�<�ԇ�/�+���,��䮙�ɗ���:.��ؔ��u�܃�.��p8��vuTu�� ����9^u�r�/v�1���6����W�L�`���L��ǳ詖��]K.�Ц�{O����9�>=J�*�"m@�w�O�V�J�,�A�E�6�( 5Pe�!J���c>�w[���!W�Zk󩀲�{j�Gv3�	Ƒ�Rt��o�'n=T�;%�P@H*<[�"�J��gB�X\�_����3=u����w���ͧ���������i�[���G��C�	�T���~;59w�ɼ�]�ڌ�ˊ�2����^�dh������>�8<O������9�L�Ce�Z�̫��n��.�d��+e���r�����	�����Hg�5�{"�Թ2��r)��}�
��>�tx����o�p�J��le�=�����$;r�L���@w�>'Lz����X%��Grd�ޘG��9,u���w�JӢ���^oS�p�����w��d!&�aY�Y�H[�l�	:Uzb�XFmZ_��H��G�=X5,Y�9J���Խ�2�T��p�#��y�*���{F�|O�9��
����Dj�7e��-Rp����̋~\/���X|���E]�j��E:�,�����!U
���lX.ܕ�9��6<��N	W����P3ߞ3������Y��E{�KAz�6�pXX���<�Vgނ{�h}�z�S�nuI��*}��F��;��;�`��^�������uM��qd�Q��jNn=y�Ǽo��]������ T^�߆:�R`��X��5��N��\�^���:�E���]�i��<�^.����@~%t@�`
�ݑp�y�2�1l��G?��нS�{��������^n*ϙ<
��Tés:*"p���.=Й`dC�<T�9�/f-H�[���m(]����A�=c�ܖ=��$�>�u3�1S�>k��5����SRh��d�XiJfk-���S�ڎ��Lh��ߤ��X�b�U/Y�,��;ub��ӫ������]o�������J��Q��y�{T�v.J4��(�����n�x�c�*>z{�Y:���ۉYo��-���_�{!�jtN��N�ع,�"�0��P�%o�Y�������+�������0�v=��r���,�	��@8i��W��{�b8����3�U�x>��P�7U_*+u
n�,s2���!�4�b��1IA��
�,���f�U�š|�˫/n�J��0� ��Y#$wj����ִL�]Y�vMq�)��͢e�
)g��nw+��n���v��ttZ.��P�1�|�;�v��=$LJt��>G�c8��1��[g��x�OV�~�����~���op�#s���>S$�"O3����YJ�<;b��P�}0���L�l�� ��x����).�T�.x��pzm*g���/\����NV��J���Dy�!'w>�4�%�W�9�pPrD+Y ��eǱ�G	�]���������v"K[z'\�M�_P�Q��T���5k�;��UcG'U#я�=3~��ֽ�,_����[�ɇ�wL%Y����mR{}���z�b�����W?���Su��g��{�F�P���x��45^T���d�	��fC�1Y�y]��}�=�8��Tz�+�TI- ���y�������h���3��;�=k��\C'/y�~ђ���w�D�J�T���4z�G�b��}.ix����N���w#�N?B�7�w��gbw�����^���U���AmL���	�
O��ڗC�F�_w�]�(É���]�ast�^��'g�mĽ�Y�WժN
��ݨ�s�pw��%��A�O�W�z^j�X�*�"�ԍ��� �+v	��^G��+%���Bg���2�-tY��2ĭ�z���u+��*Tǻ?xׂш����L���+�Y8]���3������o��gS�`gk7����P����V�:ܶ���A�����c5�-%�N��Z̈�1�	W���z�7#ާ�+ԇ��1P�*Q��<?U0�A��ձ�ۯ^jR3�V�G�S���߲�,���E��l'�y�����f�{b@�q����/�������J��{��J\\y�y1upw�U�GWeD��=M�>+�$=>�j�p�x��5�KL��z^N����x�>�d�$ .u�c�g��k�E����k�.�Glj�oHdT�u�C�b��ѓv����0s�؂��>�/�n���X�Σ>T�c�[f'��f��躜���j�9��k�I�|ۨ8�`��7d�uG�G��п��^=���yomc4���E<̮��������&z~��?h.OX����Oa��}Dt�B���ُwQ�^�&��������R=��>���ϙ��*���,���d>2i�Mϣ��h	�16����齔2��(��޸|m�m�c�x�@zo�z�d3�b���ԃ�ôʒ�:��aއ�Y�{����jzR��B���*����C~���@zNz�
s퍿>ێ�j����0�%����/T��9�����sx=^��jy�5շ1�E��j�O&��s�Z���ru�C.f��S��fA�.�s�n�y�h<�P�_�~�zR�3~B�R�=��,ޣ�ڣ�r��o����~[+�f�t"\�N}��me�ֶ�f�)N��G��ݙ���h䰬l�wY^qJ��>�<�}y]P��,C��+�1�ԛ��~��T��s�7w\~�{��<m��Nlχ�ӡ��9GEԪ�N��g{=��Ϧ�V�>)o!'}<���׫�Y�X��J���Z8��c�b<^��Dٔ3bI���*^���緣���:x��'�#�]?�0�����'}KT���`M�&]�\�=��p�p��c�I�y��(�莇���m����������_.ʑ��Q\$���v��v*�@	�ă�Q�Q8\xp�Ϊ��e�h:��*9�}/���V�kv��*�3{g9����%N~�\	1��(T;��n|3�Yu,�sB����G���UlQF&x���� ׇ����3��� -��~
W��å��k�������=cёN�˱ǧ_��pg^�`C˹�G�F_{}q;�a�,� %�@>-����:�gºw,��n�C^����W�g�7ѽ���C�;�1y/�~nw �i����p����	�c"#5r�Cj��deP/��5\e	mK��v��T���s뙈�@��f�%,�x��U�К��Ε�K:P*s'u��Y�F�d�,k�P��T�ٰ��V�Y����X����{}���'�⊺�(���Y��q"����i�� m͜2����$�Δ����yєw����Q����8_;���.tl�l�yӘ:'&Ӌ�Q9u�v
��YY����ѺSᵽP�TC�&��}�J�Ƽ �c5�u����h8bWM{n's$z�ϔ�|*�񿊜>��S��v�%/��^ۏcU^7���9U�OJ���gs�5��
�}�T*<}�&��<zjJcӁ�T�:'_W��ާ��ˇn��׈��u>��u�Ff���ˏnnB�М<<J�_�kC��i�p��Ր_�������Ws��v�o�o���xd?W�#_�o�8�U��7עŻʜ7��ۃ0�Ў�d��	�0�j�".R�Przxϟ_��ׂu^��z���걼r9���W'�Q��K;q�^NE��d���f*Y#�:|}�qYU��_�Q����"�T�rr)�j��m�����"�,�g�~�l��L���$q� �%�UU*�W�����mJge�&yv�X���Fy��⼈�^����3� ��f���	A릗�T��>R�?;�}^���C�*���}v5"���Ba�u�Lu	L\׶j��P�\Ȧ�v;�.x�x+��L��ߞ�H��v*k���F��Y��,޻'��;8�d@i�H&)�b���Y\8oB; Ζz>+u꺌G�7�A��i��e��T�\]�'s�.�t꒳xQ͛˓j%�a��o�}P����,�q �,ȱqR�x�̩fX�k��*��	Y�u-
�4��C��8�Q����������0{�<7@�� ����X�׳V�OZ��Y>N�%\S�p�q�~�}^eo�Tt�l�8yӨw�,� yS�o][>=7��FVl����nP���0�Wcډ�/o}qT���RMǷ�#�=T��_3Ã��w�uL�F��.|���$9�zKG۰F討��¯��w�l0���uT�2��\�=��/2�g��8���Z;��6zH���B��T�����!Q�j�&��O ��N�Mn{\,�݄���%�h�d�E������t�,����q��*|oo��ݙ��r�	o\���Uϝ+�eǱ��&O�]���2`d���1_D��������P�Å{۹�=ij�>vo�X�CWx��w"��zg�> �B�h�w�����>0����,���ZDgeD�B#�)_�4�<�9_�μ����_�x�{��x�{ؘ|�2����8���m�g�_��%��䭡0M��0�1�
�j�L.a���b��>�T��)�uò�����xZ��Q�F�:s%���ʴᛓ{�
XqX�����Ѭƹ�b�**u�.��������;�:��*.7-c(��o�|�B����*�%X��>����k+��Z�y���.qE2�S�*���D��-�tK��7,��*J61���z�(�q�8����iԭ��3����Fك �2�)D��Y�$c3�]<����w�hk2�3S��Lzh;/:���kL���"��p��N�{Z���צ���ՠ@ㄍ��a��<�|��!R������`��m��x��EAov���7�PRD'I _vGE�$V�b�`�z���O4.ц�߬:�R��H���~��~��J>.Nv ��jPU�{� j�Њ��̧:eq^T�T��]E�+�1c	�]����_q�ފbo6��e0kD�L�a�)RǛ3v�����'wJ�Q�,<ܨ�+7�l
���T3n`tq�C�f���u���v#�f9ܹ[��u�RAt�&)�Q1��xX�&|a��}:QUz��ʊ	�<y9�W^�sI���*��Yeڀ�T	�b;���*I''i��'{�z�^t��a�ΤL�Bn��̱CaMt�v��v��U����xpNdӧ��'��l��e��B�Fܣ8�eb��
�q�D�Z�O�]W�А�ò��.�"���ڽ�7_K=�����Ώ%[vܕr��C�>qr���`=�y�k��2��YN��㎜�u�E�-j[���dLPX�^��]g����j�#D.�W�Ge�V�Y�4��]��<5Z'6�-��D���:)�*`ۅ|��[S,B��Q�`����\V��D�c�q��s0g� ��L�C�su����*ԛR��(v�e�w1|�S��K���:�Au'��1�$zx��$-�[֣K�i�w
�2a�x�Z�{��`���ZOP�w[g����i Q'���un4�_.���\;t��i]hQč���M�Q�ip\�e8k�����Ł�;VB��L��U�FS3���k����]Ѕ.Y2k��1����k�8nR���t�j�n���n����k���
��b�т�s���u��4&9�?.2�vpX�Y1���w/
Č��-`�2a�[�[4#�x,r�T4��h6�A:x���	�2�;xc�K�����%1�e�D�yN�j�0)M蝦��AV_L��5<�w���2��u#���uX9��EWmt�r�w��D�h:�a:j�쵸��ڻuAn�j��;�D����ĭ�;�ͭʈ�,��ԫ5kN�ݾUݺ��6�Ja,��[�]�r'D�������B��t�f�;�i(�"p7u��u��9�vY���y�1/������_޿��",Pk�s{]�Q�C�s�9r�\��9��F1���!�n��͹N��8b���n��wG ��nW+��s�w�779s��4����ݓ;��5˕���n�b�\ڍ����v�	\�"�GwG.�np9�;���\��*9�p���9�(��t܊屸����9]
3��&Ƣ��ܨ�M�y5�G776��b�4SιQ�ݴr��9awj��oK���-J+�sr,��\�خ[��[��.k��sם�'*wh��*(��M�A����\�F�\�*-sscF���q�;�Q�x��x���Y�^��w9y緧LME�Fd��4�����c�JS[؅lrX��'>����<�]�u-�J�wK^�V�,�N���gt�E�r��C�Gt��{�6��ݨW�e4n�Z���^OK��L�@\wLgiΓp��H�V�Ӿ����ŸV0Y��Du�I����AP� 2��73���u���=���q��\���#���������n,m��B}�ߓW����W3�x�8�e��x,��Q�u.���,�zk�ճ��HO�U�j�L�`=��@���?�SW/�u�"�Z������G��� =+��òc�H3�:���K�;��xr�7��B��W����yש,3�b�eJ7C�0s������z=s���}hY���������k,B�{ՁG�¸y#�)��<l綢=Dhf��[�6t'��M����$�1�=:�tex���2:�*&�:z�����<�T=U#`���x{:��򳒤y�@6NӐ���X���Ke�>���*�^�ZG!���9�}�w���=��\X>:kͻ���f��,҂U>�&%��lt�7`9�n*C���'��}�y���TC����ࡓ�
��A�UxȨs%�U0ݎ�&$�)�t�/�?����ˤ�5���2���0F�V�:���Bu�?���ք���/�T����t5y��c��{����r�Y5��_,cJ����b�����,x��f�{@�Ӝ�:M��wdzL"�<�8���t�p<K�-\Q��5�5%V�d��Y�H�������~W�Ǐ���wĿ	����D�\��az
�2��r,�}{s����m��v�����馥�8�'dx_���E�n�O�<g�w��n4
~ːQd�l�b�]Ms�z�Jږ}H8sse!q���p����C^����W'�J���q�C;V2�������mw��yW6} �d����5�_K��B�����^MLws�A�s��==��lK}��w�US��u���kط,x{&o����¸����Օ�J��x��n��tuk��G9�唖b�!<�ϯLz!'̽���q����fp�㓛3���l�w9GE�J����X�5^�X��nnۻ|�}@{;�C�^���9�m��,��Y��((��%�W/Gyߨt12R�[���]��J��T���k�R�o�F|�z�Ez��dS��y;ꅪN
��t��0�;�C�R��˺�����]B���F{��lȎ�j�og����1�^�<D�p��|��C홭z�ۛˠϔ� hdo	fD��T����_vuTu�� ö�7��ȼ��x��J�FLSX�:�e�@\B)=���ĭ�}DLOwi䮡�����tơ��e7���[��\�5����Iw�"\����3�=�2e����l����b���k.,�(���x䊑�z{��qf�I�xZ�K��Y46��;�-AS����NW@6O��,z�&X<����t,��o�n�U�4��B����8���+��+����\{U��m�������`HR�f�-�5��MboY�:>��>�����+ʺ�ѐ�޶�x�<�����S0�g�����I�z6Տy�H�U�ݮn�D�_K�3�[�Zgޯ;cYO؛��*>i����p����1�Y>.q�0���j����ͫ��&=7��7�����j5�VF���팏O���&���p�\L@�&7��y֩RQ
o��X6�����:�@�����Bc<��I���R��^ w��F[��j���AR�<ݞ��/ ?K|���f�*pTK��W��z�%/��^ۯ���� ��Xr��
&?q{?)���l�WH����Ç�$a���.�����i�:��-}�O��>�R9�Mi�b0U�����$��wve&�YÏ��*��lT``lǬ�l"��^��1�f��U;�uժ���������u��ȍ~�ޗޚ�o�E�W3gC'0^�]@b����o���t��R}�S�N�v2e�y�Vkr��jJ���f���U��=������'�CN��;ۇnJ���C6ęs��GP���d�w5P\�|�)f	��c�g5��ϻ�5������S�5b{�����1Wgq͎�d���B��q���.� ��;��u^����x�^��Uo�\������<�����&8��A�7&D��`nyK Tbnȿ�O7'"�F����瑄������i��������0���91��tWӇ�υ�.=Й`>�/��^N��I�M"�^� ���qLZ�p~ȱ�&4�~uA(<��ʶ���c3����8ip �'���d��JO��L��P���G��7�� �A���X��T�WE
��r�i���n0�.ZgӇ�m�X�O���<����u�y�{��;%�|ITe���x[��j5��n�8,����G���)�^����^�p�~��ў}^elyQү�HN�.a��˽w�9G�����t$3��@���O*D����f�Q}�QK��3��Sg<���|�ч(���К��}W�z��#�O���� '5���\��h�t:�E��7�l�w��}ռ�z�R�y�0���ѭ��l�$�����zH/҅J���P���!Q�0׻����?Z�|7�y�f#��@�1o��j�{9�b���I�Խ��T�����v^R�(�To��NSm݇�Dy����Ɗ�׎��2�N_:�dR���]�P�oX�<�[zz�ݵ�}Q�N�A�ڳW�X3ejݚ�e�r[�C�+����jc�!��H�p��;�}��h�d�E��L/`��Y�];�F�_8���<K���A��o=�";��!�.=��b�av8��fX�a��Fo�)aL1!�e�_�Ν���N^��oSp���T��?P�����/^
�ڐx���Y��B���Ս>S�u�����q.R�{՛~.3�/�>n��u�G����x�{�V6Y��c�]�|׀W�珤w��;�؀�é�z����<����lt̴��sR.{4)��� ���s���o
�QS����f=�����a�x<�D��Wz��a�^��sP�*��.�Lq�{�F�g��C@q:V���1���U��[�:v�e��3�I��.���_�ï��jP!*X��<��ߨ��@�!����ȯS�Y���|�|�\jڞ4<J@�p�2��8o�����eZ��,>���e�zh5}^_�z�7ޗ��+ԇ��0��Q��;\.5�{=wJ59��zAɰ@�>����;S���n��!�a<#�7;�A����ͭ��e��0E��ZbW����7�L5}�%C���^��v�ƶWM{�t-%�-����p���OE�O� ȕ�k{��fM�]��4�#�	��x^�Z˶�j���,���0�n��@�nB\��X�QǼ��̿����3`�Q눣-���'��ڊR��}�'�{>�Q��i�!��6��y�.ޥ���W�_�uH;�� ��@n��:[/>}V5�~Wz�ic�eO�nb����o� 2��q�BQ:>T̳5diA��Q�p7�����s������^�SYK5(�����:��l���2qM����X>����H���#��)��W+Ζ�ʧ9��}��츾�E�!�a�{���j�~�+>9��wĿ	����D�#.OX�����-`5��V�dT���I�}/Ԩ�{f�*���y;#���]ȿ�u�}�3�;��7?e�9��@S�/�1F�V���S�'`�fܔ��-������Z����M__:��W����[�������O{<��d�!�ڔ�����PF��.R
�a�;�_μ�x߮�����T��e&{qw�g���O����?nX����,,�����W�7/ʧg�0��i� �C�o1���E�X@�|�N1�������Ǎ�8n����g�����+��o�6m��i.!��6�A�5Z�c�A`$� �j��ʗ�N��ڐi���<!�y�����J7}������w	�i
_82�5���h;J���C���_heY��#cL�a���b����8�U���}X�& �
��W.	Ӛާ�ӭF�Moi�{��0*#s�#�̯_�W��Y�XYc��
h�h��c�ood�ɼ�lը��՝�sH�r��B�o�F;^��^�������H_ڶ���!�����@��L$^b>����Xj�G��R3�@n6dG(ݐ��s���1�^�<�C��3�kL�u�8�zC��ʑ닖I�R|�U���� ���C_�{NG�O�����J�mj��[�k������NW`�*��z�X�0�[���R��;ub�*����V;k$�-��8�#�`���5�A�S�F�<��& )^3��6+��]ݹ���1{��a��b��Z3�>��v;�4�������Lø%�P@HwwT�{�0��]��S�̿.r@G9�y�Ю!��=>tÏN��bnw ��u9sx�5�	�!�����c5g��	d��Jt��#�_C5���8\7�ldG�ԉ����{��p�';7҅�ǛQ����;��z'�g�>�B��D����n��z�T?LTjj�%{ޤ�A���FS�ZcE��gj�N���&E�7�xz�u����DZ�P�H]��@�JǙ{2���C��ni��ذ��p:��w�3�+�;k2
���u&l��sWVo �j[�:�mwu=zIf����b}&YRs��{m��-50�L��ȳc@r�`����i���JL��Y<+�2�j����^�gXT7!���Cੇ��/:�{��s��I0�E|۟{��bE�^1?�.�~X=uMv���K~�0���m�|N�K/�3oJr�̫�ˍ�U�-s�d[<sr:04��E�}8���
.7��7j���s�볧܎}�����!���{�25��z^�z���\͞��ݘ�#Ȉ�?K�m�u�E�O�Ǯ+)�Z�.� ������K���X�9�2��9���f)�Nz��m��G���'v��{��eV���~%g�i�+vE��nNDS���fn�k痖�{�R�s_�/����G$�\�%�����B�L�<\"4���x�-�5�5U��*��'�J�E���ȯ+��m�YӒt]�I�.����4�r�s�+��L�L��1�ڢ�e>ܖ��0��X>�m��g���a��7�te���������|�̱�w�ӓ>+�y��][ެ>y�(ۿU�����p�!�c}�|w�U}���4Oѡ�6l�#+�l���"�ܬ3�V�6K�dI�<.���E���K,Af2�5��:>�0)��~n��u��F�}�rt�ޚ�\k��F��Y�ߪ��[Ys���I��Lz�[�s]!�͈��i�|��;,���Y����犔y.�5*�2U�*�0WE��\9	�����H[g7�`��n����/>E����6���B���9�<Ss.�=�=��VϘ��0z<�`����0��	����M|���8�z17;�j�3����\�����8'�zd��@r<H��끿�KG۰F�>B�n��E?��1~,w�9cgU^���}�)��n=�_~��I-�ԶnI�HUҦ��_�hP�P��E*k��B]�2=+����2S�	^���=1��az�u`�s�4+bOO3T���-���5��O��ר�\?+�1p���6�>��Ȇj6+�a�jd�a��B���UvΗ�� �R�D2����+'�U��_�ڻ��B~����=3��D/f���e��,�e����)�����X��
���T}�ܹ_�����ng�q�C2�Ճ��s�{N���;�Z�זpI�+ʑ���;dfL>��#qS/I�q�y������h�9�ʱs��C���y�8�z9ܥS}���rN_O�Шu�0��s8*>�u���#��l�_O�^-��'�;]��M�u��s���*�b�38x[�+��zga����SFeELP�ә0QI�ὐ���'n�j��K�ٙ�u�x���6�FP�o,�ZSf�ZS�M����i4�:Թ�ا�m��3D��A4����c*��9�#�'�w�=s�Vzy������ޛɝ��͙c+�3�]O��	��S�]%�Ѿ]�}�|T�������r"�O�e5q���|�^���CĤ)x�ro8�ϳµV�x�0�評�ⓡ��z�<�o����/9~W�1����=���1�'G�t_4Vʵ��*�� O�-s�$���r�
�V��,��z�d{���s�u�z��Z=u�^1��������U*��o�\�5"�>��Á0|��FX뎷q>6���\:w�9�'�z6���hg��ٙ�l��,���%R6�Tÿ��UB���I`Hn��`���^Z:^�M*4�#
���Y�j�u�q�ތ��3a�Gʙ�zdiA��Q�p7�����l��1�"��M.�^�-	�ٙ/�q��E�2����6�T9��#�'d�q�A�ό���Z6������=sBV�3�����5~dz|�����-}�Q�)ۨ��e���ϔ����߻+�~���1Sʕ˖�k"�u�����z��~�����y�����ƶڵ���[mZ��km�[o�u�խ�V�V�����V�����V�����V�����V���km�[o�+m�[o���խ��5�խ��j��o�k[ko+m�[o����m�筶�m�뭶�m�筶�m�魶�m�뭶�m�孶�m���j�����e5�u�� =� ?�s2}p#�|y�!R��J�Q*�P�)""�R��%RIQ
���R��(U*P)(�J���R*��� J�UH�%��!U(=bl��kJ*�R*�ATtAUB�Q@��
)��-��Q�l)U!�n��T)_m*$֯a�H��*�lPTHP�J)RD�$*�*Q)%UD�EJD!RI%E[�	*J
AJ��P�%DERU	� 8��yvn���cwE �k����Ezwb�ny�^�%���U�{j�����UM�7�k�(�5]�f�֪*�a��Q{o�5��
�C֏cU@�U� ��͟s@<j�RU��c�^�W&������� �㣠4t  sŀ = �= h�ttM�׀ �EQ�}�L�4Q�Ѣ��V:4hѢ�4Q۶Ol��kJQE/  �4}��S皔BU�X�=��{oyUZ���^n���w�ѭ^�uTR�w�{ڶ�����@i���]�k����@�H$�
�S�  -ǻ7֣�Y����{��Z7��o[���TN��hX�p�V��v��m�*��m�ew�ٓ�O2wy�{oy��U��u趪��*��J�H��4�G�  w�]�}�hz��I뮎����#v<�]��[��{��y������Nww������RzWk�'n{ݞ\�������������*���靣cn^���]��Ǯ����%֥BE*B@�� ���nw[���ou�����ohz��Y��{��g^�j84�;����U�Y{��o/wN��/n4u<�׻ݻ�U���{o]6��{oe�%i���v�]�o9R�i6ԠHD�*�  6>���ͽ�=����/wtR�꺍�ד�n��J֍�ӝ�#���)^��yⷫҶ�;c�:��O/^��Uoe{��;ۯ���ݽ��v��oE��(6u����ة�H��$PT� �כa}�TzO^�:�`Cu��ֺ�[i{��=���W�;��{{�zv��o-� 5M�ݞ�ǧ�h�ݱky+���m�j��.����Sz=]����y	%*���$�#M� ;��}ޔn�z��{�2�����s��{�z���;^�������o!���o.�����4\Ξ���s�{������f���n׽��c�ڮ���G^Eov���k�xzP�))D��E
R� ^��m���㻷Tv��;��\��z�����{���=�:���yk�V����l�v[έgG�s��=��׮�v��N�z��r��漏A���)�4��JT @��a%)Ph  ��deR��  "��	J��@� ��'��UT�L�����IF��4�O����U�U�����"�_��-���6�Ts�ןu߮�{�_{�뮽��}B* ������+�QE?���+�AW�PTAY@QN��V���������Ⱂ�����6�%�)ۓm�m�.��i;ڔ*�Vb"��p���Z6��*�h�ܹC��]��T�?F�Y@J��xU�yE�ȫr�\ƌgh|�.;A���;�B�y�)�h,�&����0oI[�EKf^��m�
���Ҧ㫭�LZ�َ�*k!�Zڿ��ᑶ�EAR��EYr��N�ˣs.����)��%���DRP�1P�x��n�:���@��v��nq��ܲ����DAt~��8���Tr䶦�NY�5���e<��t�-q^3F�c6�$<�Y.�1X�r�1�)h�.��Ze��^��hŬP�o�X�H��2�۵��n����h�ʽ���ek�l:wFdtqȭ'�����Σ��-чh�G!ʇ*m��A��u��$e�j���bHe\Vh�7�4��h�6��A�-�Q���@��ܖŇt��pV���!D\�4��5�v;z��ܽQ&�xaN�D9M���86���7�WVFM��(�Z�Ѝ�Dٕ�5�v�u���z)ݔ�C��*�f�)�N\�Ax�uy-���r�]��m����N���4�F.��o���]���������ڠ/"!�]�&�U�6f1�1�y��ҹA�ǹt�n=r��L̲�'@Ii� �XiN%%���ۥRӖf7�@m!�I��S�Х�b�*�q�:q@n���Y�KD�:�WMQ�6VF�n
�YwL��A���CØ?�JIư���$k�`oV���3�"�T�w
 'nm�Ԏ�W�@��#KiP�J�L�;���Ê�ј5Lzʔ����;c{@�Z���T�e1<[�+iAR�T �C@w��OmAP]k��ۀ��f������i-��a����p ���$p�/�)���5�a����œC
ۤ�)��pdW�\2��X��x��6ـ�LB��t�A
m�M��ݖT�3-TL�{��]1��0�wwH�GX��@3EZ�@��r� )�.����ߖVI�m�����⳯e��sm�SK>b��04�y����Kv��ޫ1MB0*IG����[�sK�Un��Q=3Ja�Im=1�,k2-+\>����f��[(lT&�$Ø�����Z���.|��µ(�U�*jF��Eꈭ9tڡ�����óS ��x���N;oX(�1��d��q����gHjµy��{��h�[��
oH������eᗛ*CelR�(D��p)��m�b'"i�k�M�ߴsP��Ã�f=Z%��ImUޥYv�F�y�9p*��som� *7��f�,��.�sP̥t]���K��\�$r�i�w���QK��fF�`4m�o34͕E��>���(���K-u�6�@Ѥ3�F�+e �K�,���.�Ԇ�}��sV�GI��ג�HUWD
�in����j���¯��7K���7�T6�͚���a�	���,�%�
5e1e��(�@6��skv���"���@�dtN�ⷳ�+CKE:�M���N��Vv<���� T:a7P���sIk�B� &;Y������Ǥ��� �#7H\���Ŏ���� ���ց�I���+{��a�NI�Ke#��cY6�r㻴2�FcF��N�۲�Ȋy��Ķ�ƅ����j�8���PÍ�*��vD�d��5s�aiu�A�2�Ò�LB���[3q(�jId�m����T(�X�Vr�[N��69f�L�t���AhV�|j��u�T2�7�)=I�2e={W��4��I����Ԑ��8O���M��c�Xu��6�fdN��1d�j��n^%�Z�K1�mmZ�YZN�(.�J�]<��*Qd0B(�&�H#k��z�5YWt)�[����VB;0�m���j9�cWX����1PI���IRr��b9.�����<����$��j�˃al�u��^7o%f	��������d(՝VUb�Z�,a �����y��h�)��,]�9A�/RW͗-�,�Ș�J����BV�!;#���5��U�N"�h|[�XH�R����R2܍eb�JfmS��t�PW�Uc�J�a����b�%��A��{���SH�B5tR��*��(+[BM�w�A�Q���#nɣT$�$���L�f��m�e޼@�j�lo%CsD��
'\��7Rm���mݔ��5R��{wkFP!Z"P����1��F!�5x��m�J^#Mà��r@�{���7�2GL:Ln�ܕ�o�ꂴ�!qI/XU��j�ܰ��Bk,^��(��Xa�۱r���T1�ۼĨ��LB(+5��莭�i#^U�� ���1�!&%K��t&3~�D�X�B��������/#-���I��jƣi�{a���Ս��;Y��4^ĉ�z�Rހ����Zz��rm��L���S���y4£;����߅�d�ٔ��V��AZ��O�ebJ}	'6έ�)n����I4b�+)lS�/#�CY!զp�A�tޢx	K1ޚ�.��C�V 6��dm�̶ٹhЦ	V�Pz�(U7P�ZXyZ%<Z��~�H�U��t�um���O65��ݓ)]�={q�\�LmZw�̧gU�2�5� 6�����d:W.�9z��T&ܳaAp�f;��5E5����Xͯ������5#�%�M&�G����Sӻ2f�h��m��߬�tM;�(j�m`��#%�eɺX@��}7jAiM���7l�q��g(�0kA��4Fe�)%ȃ:)EV�g$�!bҒ-�:�̭���Ո����p�ǥu�-h!.MScu�J8N=(̽Tͪ�{��H3N^�Ԛ�x��^V��Αv�T5����f��]e=�b8S�֍�7� �&%�n�K�G�T�%�[�VI5�"���R��C�J�`�V��Tۡc@jۗp����}ӑ�$���X�	�l'�{���p��³Iڧ7[,K�#nkZ�Ś�s���55
���h�.������TT�-�6(��0�ʁ��8�]����>*c���E���@�@q�J�����('0�4�kBL;��oT�RVI`Ջ{r��M��0����� ++W����/@[cNK�دPov�v.�3vSV2�m;�c-V/�6� C^J-=�%sEIm��(���%c�!�Q�96CZ1̋f0TYm����J���wJ�v[RV藕��(&է�Ú%�F�����hШ�n���k/h�b՝tm�++(4���kr-2�B�ɿY�e޻8�j�c��Qۏ(a"�1u���������������-�&m�]�/i���Y��R�K+.��юڔ�hB%QK*�����5 ���$�	ʌ��\��f�(�7��25����r��,���I����<�)i�e�5y%����U���	�õ��4ڬ����P��"����n���$a�\9z揮�a>�%������b0��4��C4�b�5%�t�T[S("�����Y��GF����u�d��f�hl�˂6���=��A)�-R[īI���傘t]{`��POBX]�[i`̆�T[�#���QW*�[.��/h�E[$h����>
���=y��C!�$f`�B9X�ⷪӲ�&�%!3lږ�}�y��*��J���#�Yt+�Oi;��)'G/gұP�3(8�`�&�,EJ�[�V֬�d5w8M�X5�@�O~�6n��@�mb� WX�B��%)w.���V���$D�kj ���[���2�*�f�tSǭ����:т�a�ח�%�V%aŗ�:+Mi�w�0���/3C�(`�*�ɦ�]*p��eغ+P�3AH�6Ag�խW���q<�X�m�u�_̀��T�e�����+��5`�!��hN��/*	��b��q#B=7�CNr�ܛ8��("��`���U*ʷ�6��Kje�I��(XD�e]ڭz�u��[v
ˎM�b@D�hE�6��SC/53�\�n8��t�Xh;a�.�a{�P�)@
��)m��a�v�ͥr��M"�f���GD9l�8^�t��]J��ƌb�[Q���[�j]f�K"u�������B-�ayoN5�2�7u�b;c`KlYi7e*�A��h�♛���b�#���4���x[4�7X��XkXv�ڸv��ʴf	hpM1��s���Fe14�`��ՠ�]-DT�2�[zѵBՌLP��r�rG��K��̱�S�5���b �d�һ����ڼ�8�j2�A�Y��ŗ&�3%̐��Z�!�l������:+x�1d-T�ʳ�X ¶��aތ�WMP�e�ZL"���cYr��|2��1�ۄ�5��ȥܣ�{BjvT�)5K
b��J�ьn�x���d��PD+F��ƩmH�	Wl��k�wrA[��3�A#����8uWu{X�
f�w����2ը܆U�Xku%#��k/����ө��Fd�-��hD*�˽��q�A8�6D��X0�W%�
i �YQQ�ۥ�����-P����E���y����:Ղ��XB��V���[Z��u�-Jj���Ø� ��j�~t^c�&č��,f	g�6�?H�wx�n;��S4�ٷp�>#G��MF]-e�	]�	�Ӈ#D;Ѷ��0�q�X�Y-U���Df��6b�,)�ڀ��J(c��+q]˷r��B+��N���#	oX���U���e��aP��"���V����,2K	N��6y#d�z�[&Kܼz�*llK��v�+La̅VX	l�p�Zwǈ XP(�(��qӶ�]�Ŷ�1���j�=��%��͒�ԫ�L��Э����X��ں�"=�4�%�s�)�AQ���śzt��g*ͫ�2�^ZՐTl����R���L�2숥<��k��/c����V]� �S;�IyP�]�@��M�n�Nը�9H�B��dݖhb(oл4��VӀ+F��7��w����"��ݙ��b���[���[��AM���0��V��KMW{u�D�b�c�PÑ���0$�#�ˎ=wEaق�ѿ7)-ŭ
��!/;Eǖv�j�/!�Gڂ��`R�̻DҦF�ـ�V�Q<Ùm��k1��R0/�ܽCEؘ��Q�桱�� D��۷�ݚ
��{Z3��u�1�?]�e�Ob�1f�����Z���tjYD۸5�-Y@bhV���/fɏ6V��ҝ�3mŅ�@S�n��hٴ��	�I��˧wK��(C�mb`kʸZ�^��m$BҘ�E�F�Cn�0�n��x�%�+
�k�eGƥl�,���YV��D�^�DP�.[8pM��(ĭ�Yl�gt=��"-/3n���-E-��5��kSgL>&ѮV��b���8rd���T�kJ���۴V���n�+�̔�eb�|EEh�j�r�bl�9�	$��(謼6�Z�f�����v����G+1*���T�y����G�) Hd5d�GT�u�t��U�$Mw)�c�Mh��ڂ-� ��A5E_�cdB����Ȑ&�ؕL�%�[Q9�\���J�I��-"��6F5yh`�P��.`: H�b�34
�Iaf�:�GQ���F���,J)�r�i+�T��t&��P͓F�fIz��$#B��3%�^�Qe��ja� ZP��[�5p�Vm�1]��ͽ�`�Vj�r�F�,=�Z����&K�Zs e�5Fm�G��yv�ȇK����ӕ��z��˹/+oE��n�N�D�!��*���Ȳ�#!k�e:�<,���Z8PΣ�t��1��ț�����%��tAssd$��;1�KDj���ʸ��MlN��N9�ǒ�aIM�4�r��弰α���xw��qŷ�Y�-4�l�M��!F�m�f��gfaC�Q��97�Q�[�s.�*	/��j<¦�f5]L3[&nl�:������3�ԏ01�˒p
��U�����j�Ǖe�'6�N��r�Cw�ŉ�Y�VH֍��bwP���[�cw��^�a����F����٣��W�]�Y!ִ���Bޖp\�L'U�j�˽WZIX����QM��׹�qOZ�,5C�,\
4�"��OA5�4Tz0��d'wl:S�;hӡ�҅��gFǺ��E<��sPC#��3q0u�����	6/i�hW%���wm�4ޡ�w!�m��5����)�wT��J,܅z4i��Q�����2�Gj��o-!y&���%�]=�R�{6M��R�f�Q�Qyl��W�� �$�uf���0S�R�И��.6ʸ�X.f���ۤ#�=Š���p n�zD�4<�j,Jj���b�K����� ���L�Ks��pm��^�t�*�:(�Q����g��u�:, i���T�8G�M�ѼJ������n4�b��@�EaxS��Ʒ�2��h�ZMM-�	�[�����0�`�f�=�6��mm2��q-��5uSVښ��<#6�*����J
�#��Ђ��]˦�&CԌ�3{GVL�������:�&V �b�Bo��"�a���,�#HB��;�t���M�x�OS����(:Q�*��[K0���+0�6�03;7K^ԋZۧ�()WX����7�d%��Q��e<���8zl�~r�`���� �F�8é�����7w%�GA� ����)�ln8j4���Qf'��`��Ĵ#V����j��Q	��I��c睎�2w_�ztOf��&[�¹F�E�]Pq��G/H����o|��^s���U�%gK��n�whp�j�.ͲM��ΓdɼGT�¹����!����b�*��+��n�[v��R������z[/hQbb��JBo��v�<�N]fV�Yd�Heխ�3]p��е5a;[�N�}���\fe]���D���Cx �B#3o��P�G�@��Ա>�a��4B]�]�
�Wst���ƛr�%��g��s�ʓr��:��pr&m)�7	�f0شJ	���1][\����:�eA�M�lę�r���
p�y�V��|xn*��P�|%1w ��������^�W��*�Q���볲��5�ƕ�!bݺ��6��]}����� ,fJ�c�-��+}�t7��+����*:Y��񸣼N�%uk�ȫ6�J��i����G7��Tw��M<�\�,�6�7� ��gGJ�)���kuܷ#�E�kr��ɩ�sEPe��N��xy�^�N�o�棨jJy|eռ����q՘q�Vx,O�i-��ȸ�me�6�swn�Z�4$t9���p��Uloy���փ˱^���w˪�4%��0��ovu(������˸q���j=����\�����&xl�."C)eJ}�m�)�Er�0޷�Z��Q5�����p��4�9Wj_G�R����V���A,��f�%�������F!5���W���ѱ`IXmW՘�F���j'{���L�)T�Z����ZQ�yx%��^�h���a�2�滃7 <u�ER��;��@;P@v�t�0]gY[;N<ܢb��]�k�uK�Q��J���K�����J��A�·-�k�,��Kqު��K������Yu��iB�f).��E;"�`�2Л����Ln�q�Q�w��v��f�TWnS+��U�����wt�;wr�9��〫�+�Wc�0-��')e�"��lԫn��h�F�]��3�QV`!�b�z���U�M=e��x�^�3�A�����q�`����R+1�v�w�mPܷi�.��Q�Ѵ
�19�fCc�]����d�F��i�oY��\���{t����̴�{�k��駕���ʣ����K�2�i+=�@��v�����E�%MR��:�_SZ�yW2��U��Է�r7v��Qޙu��
`��sTǍ!J�]�m��*�7�$@3������`����WJ�^��3㺣E(>�%��9\_m��<
��l!b9��}��ˇ�"ZP�M;l��8��Y���3d�d�]��)>�� 6K/��ߕs.��dj���ڥig��6R��r�V�p��+e)�c;�]��s/�y@�/q��'	Y��]�[�4�Uc�8o'nß2�L M����*L�(7�GitZ8����>A+�	�C/~�:�Ve'������q<(T��+��A]�%�F#�ΰ,���oe�u���ʭ�Z)����WT�v)�Oyvs'o�Њ��7��ҕ��l�B�Ef:WiڝX���M{���Zh�B�1��۵���������b�^��2U���tVw
��VT�/)_'�U Llѽ��ۑ��̐}f���vY�VJ�(
�s����v�.�3"�o�����44��"Z��Jp���±�b�疯�
��m�rT{1wE��El�0+{��.�<�c��v���Z/9X�z3�5ԭZ���[�r�G��s��yo/���,�_bfb`0�;[/z�w&�wv
6���V��{���*Fx�$�Gt��GC
	]�m�χ�M;��W�W_q�����K�mf�ap�	�ݗ�3,���}I]��;U)�8�<�H�]�@걡}���:�N=S��oZ3�me˸׍�a�����
����4�-��wN��3����yZ��ӆG��@&@joj��~1�z�̵F��;�e�D%��KF���{Q�/��B	NE9�U�kMB��:�Xnv�	�|�r�.�!gnm	��&�X7{2����rќ%�M�+׌h�̻���$z���P��V�;M०Rڂ���ͤ;1��;�Y��e-�AZ���M"�^]_q�+f���(vj�jV^�s&HN
U�Iwr|tR8���:۴�F +��@�k�#2�c�,��?��bڸ�]��7Y[B(Z(H��-�:���k'
����oY/��꒱���!w�������&���,P�R���Lܭ�B�������B��'5��=G� a��8d����`��g��Y��Uu�}dم��[%���W�ۺ9��h=�z��s:�Wvڊ�b[������R�N�S;ڲ���A��p�A�e�6n]*Eb!p�.���̲����s��B����-s�rST����Аi�tN�9];f	�n�PXe[��iU}�í</����t���$�=���]F�b���X	u�'��"�n�*�pv�/�{Ǳ�7LgWՀn����U�X+F>Cal�N�\7�Iy���D	�)K��؇��g�K��#���-��ZC� 䑙sQ�4~����ocݬ��$ma��]o.�E���\k�ԭ���XY1�@Zs_R��*or�y�pcz�5׷R�9��X����
Yۓ7WhQ�t�>Vqd�A�Z7��C���#�3	�so߸�.�B�b'*f>�5�[��-xE�,�}�V�oH�_�m+�1Kdo�#�+�R� Hd[G�A������NF�}m�i-���/c
���<t,<N(o���5}��L;*��f5�eJ��:��,`�^F.�%w�@��j��vl�r�uEw�7�*D��Z`�z���b��^����*N*n|��Fa:�WPqޥ6����c���YA�ιAB�w��
/���'U\������m`���TP��v�������i8�]��;�C�f�ʜv�������N����ik����B*�㻒�Zk[����sm����خ��.*�&ֶ��6U��a��fc��.͔L��f������Զ�]� ,	Z�U�{{��"O���F��J��b,��V�̣�/��'j�PS��������;���P9ϳL鳮+r��۾�U���e2��%���'S*i 1�.*�$)p{�:�rS�]{h̻t/�仨;��í]Z{�/��!�9s�x�p�lv�jg�n�Ԉ����l���'rt,��W�tޙuƸ�F��Q#�+ )�LBdqgv}��� q��D�ΌeYm����H��A@�d2vs�:����K�dX��qs�1dG�o%(5��/�`�TtP���q���E��i��v�9į���8z+c6�9V7�uТ�_N<�W�t��Y��������P?�cݡ��E��ѱ�V�lA��V
,���J�5X����Zkƍ���eR0����l�9���гmƄ��+s�-Zи4�s6�}u��,T�(���PP,�Ӷ�+���Y�ǁ����r�Ew)�R��䮏t�3-ᗨc��mJ�U �(!��^�h�Oy�;*ż��n1۱J�������{M{��Lk �N���ѽTu�]��j����Ѵ
a_�v���y��c�ZM]Zk6�b��f�p��xl������W7�0v���=��*�����f��ɽ��%��bueqX���sg
�c����P������R�WY��ڡHe�rh��Z�J[[/=��[�t�:�WJ�.
�9���=���r�9�Js�
I讋K���iȎ�e�ݘ���t
\-��o(}B���tF-]���V�:7���w1�Q�Ƿ�p�
�ßp4�R�\=Yk
�m#������"�=�9>�z���t�u���۱�L��Î������if���-�pW�ǪF
�N"B-��P@��[��ԮD�!�a�v�z��'�����Ӷ��o��;��Fj���gPP/�M�S��3D�ihW���71�l�gv�=�䳫i��ZH�l.�WJ�5mfmkz�Vjו�(b��T7MӾ�*w �A�k-ۭ����/�K�G�;2w�B�$lf�h�����+����gM�5!-*��Z�c�>����k5;��"֦CF���Lk,����b��F����A�s�!�ܳ5�ݸB��N�d�d��(Y��ܹ\l�y,ѩb��HS�dhAr���l�
��������8�c�s�oWeˋJO\�㚧k}��WWd�`*eGd)�r�"�O�z�Z!c!o#��,�����{�ة��ON:��Y�)��T�<��k(+z�5�Wq����SN��V[����)\GAѽ�6*\������q�V�p����e���KL�*��L'����Z8��Q���B���Ո��γ&��qy������"�������y��:�/LWW[�b��Q��Y���8Bo�2���A\O:XO�+�٣��R잼J�zӅ�3�>c�.չۏ9��!�y��hS��{*mp���\)`�ܖ����h�	�$�B��U�d����5�v7W��;nc�����l�Z���
MIMH�å�/�U�çc���]�:d���L7���� �:IYם��44<�8X��c�D�7��� �O��5���t��t�s��=4�hלx�Xk8��V��E w�;8��]�9�����;���ǀḩ#W{S��CL��Qʊ3�9��2�r��n<��KB���ٯ�{�q7�}��/�\�Ah_F�`�<ȃ�18û��d����j��Ɋv���*۹���L�.f��w�;�kG��٫�����c'a}AاVxgϹ�#�Ȕ�Ш��d�o�Uf3�ȓ�XνX�ͯe� �I4��F��dl�q�Y�`*�h���N���qM���R]'�]�!(���73�u�L�8W:`�E�}�m:�j����4'Y����o<%]�F�3%��Tt�a�n�y�o���W� C��V�7t�:q'�F��u[=�l'��0�q�q����ޥ�QҮ̕��/����
���K�ݞ��KG}b�+��T[��j��9(si��u9���y���v�xCh&I�H����)c�ȝ�m��F�ÔK��M��rX�W�y���݌�еѡ�U�mN�s��GZռyjhNʷ�=�+�v�&�(IK:���n�����`�}�=�������9�x��$L}�d:�Cyw��I�&du3Co�y��gd�@��u���,�����2iT�y�E؆�4\w�*@
�g��k-WcL��Sh�*Y�y��5�1�[K8i��>�7.��ԟe�I�6�]���kos��O��s2��{e*�U���υs���E�a���2��$�<:.Uq����x�Yl(�����r5�s.*B}�z�:���.�
��'��>����P�ۊ�&��R�)�2���_6�9�}�0������Z�Ԑi�@��39ﭵ��/t���v��F�v�Z��b�մ�u�R�ڼ�J�넥�kI��f\���W�^m��TH#C �Wx���f�Q�B����}�E��!�Vk�
`i�z3 �����.e�df��gtT�R)F	]\"��x�F��Gp�}����*�/.\׫���Ѓ#�HۭwY�ս�������ӡm.�nĔ��yg���9
�cwJ�r[B�#��S0�OS� [����̨��6'm��묢%ݮ�zSl�z�����LҼf���Õ�����t��7C2��Nl�˽q�ػ'ƛ�U6�Yǭܾ2�r���@��+὘{��;IWp��׋��$�\J͒	[4�
�W+"0
U�7�أk+N�m(L��GHh�go�dK�t�[�`���9�s�֝���"yݢo�띭��m��\��R��X�=V��V ��κ,,*';P0�4ݾſ�v�	�h���kr�"�nc�hR�W[#/����m�7�>��wU'zօm�y��$�)��Q+	�uq���%�6�闤��j|t���W��j��mS	��V��g֘���n�t�g>޲-y�����d��͠s���Ñ�7G�����y%;��E�a]�6���7hz�h�.P�6�_w#F��]g,@�x�tow��NU`�q��)�OY��u޵�D�қ��m�6��p\oAٷas�ǃ`_opSC��^�P�=��U�4kH�D�pB���2wE��1!��A���Us����Q��gOa}`rLWj��9|JX�̩;;��[�;T5��˕`t������BkgTf�Z�������_gJd\rX�O.mf�/�
�97Ҭ�VB�pT��.�\�^��sZ���OC�k�m��#�8׎��vh�tI�f��9��9�-zhN���ݸ9�\Q_�<�YL�W`����3�[A���݋���Izm�"���gqC�:�K�}A^A]X����z6 E3)T�a�;��s���ޠQ�zFejͲk��/ �b(`��h9OrH�ȉ��Z�6����� $
q�J=���3����>}�'@o2$���cr���/ju��1?��qb���}y�WQ�,��$x�R4�b��6��|r�t���eE�2��%��`�H����V�7�C�>� �aG|��y�Uݾm�)������ �h������2�^)8���w�78��{x:0��Ts;Y|{�v��ǽ�T��l̮u;f*ٯ��޶���Z���x/�t�i
Ǽ�u�յ"��nV�� s��b�Z;�˦ɇO]�]K]K��:����HGL)ټ���Ν��r�}�#��gT»N\���Az,���WB�u�f$1^�QE3+y�y��7�|T������N��� �37�ګ�E?�W}}�Z���9μ�ޚ��Zx*�Z�JCeӇW'����D�,#��0P�{%�Ns��'\���(h�g�ǔB�Nd��]�՝p4̾}/gv��3}f�e���[�E!ݱwM2���5,
����������v�����FT��\�/�x
@b�|j(7���
�����N[ٕ��[��Rʊ�4s����+K�.k�b�Z�.�V*KYu5�
Ѯη|�":�4u-����f�^�#e����͆䘰J�>K)k1�1Pi�C9qO�S�XA�"��B�i�3+6�,���8�ړ��k���������z][��g�*H��Vˠ�*��l����<�6�9��Km�����z�k�C��;��p�ܧ(iQ��qf��Lʜ���T�xm�ʉ�y-���rƗ��W�t-�И�cȅ'
x��QyJ��K�Ġ��8b�3YVᳰ�f��j�#Bj�ö��HvU��S���N�w�)ރ�3;[!�CU�J����KL׊�o&JH��X�D�gV䮬�<W.���e,U��ӵ'����d�)_v%1����
�o.�0��3JD�:�;��P����e�I�����W&״򅭖e�Fc��(P$#���L9X�e-'W�I��j=>��@H�B��i����8������Ҙ�l�aP��;�w(]����9ט�����K��r8��^�����i�S��. K�置��Xɚ��.��R���|'i��=�x6���ȾB�5��u���f�Z���G*å�ytP�{x�s��T�ڕ�)�po��Di��NbW�nim_<��Z�K��C�s�]����ذ����Mʔ�@^����WZ��Z1��w��E9W�m�T�P&I�$fe�bv�--P@w>�:D�k^p"�gKǷs�������o�Y]Z�F��`[��ٛ����t��[ԯ�Y����"Y���6�쬳�����.�*y&]9��Zy�qd16�]�_��:b��O��b��X�%�	]MF�p�cd��0i#C{6�ԭ���oR�u�mr�zd� ige����V"�5u������'��{�U����T-Pf�fSz�V)x�-��m�f�7(��j�¥n�؝��+�[{�(oC��c�qќX��ЮՐ�i6d���=9ЉLa���5�U�c��+y��Ί�ŘP;�[�XT9<y;�_^�eA��\��Jp}�+}���,���w�1����t��h�Qݓ�=�����t�f`����:^�������+1�:���O2�D-b�q�i�^n@�aV� ��sj�l.�vf.���aV�7�j�4ay�ئ�x�����]C�j%���en��i���M��v�&�]%�$7�,�w=e,6I7�ͫx9*��J�5E�*��x�'�ﳷ3���B\ـ�p�WyI��rGG��c��r1M���Q54��)P!��3�.�d�Iyi���$F���e�p9:��D�ZR�2�뮥L]�׼쏀�%��Ĺ�J[\N|T��ʴҼ����Ǵ��ǩ�Y��=�w�]f]'Kc�t{��YϹ,\ڒn��a,pt�]�Ά���F"���c�h�챫�b3Y�eL��cEǇvp�pugp���w-�����ǒܫp�c{m�L��dU��r%5	�lm�A2��o%`�(<�'�/�j���Wݎ�1�*�1��K�*��]�Bi�:��Zۆ}�EA�ۼy�xG8��\ʽ��)cE���R�ӓ��co��WhYs�4q��Ԓ�`�"Zʣ�GnnZʈ淔���ƝIOv�r���[���a�%!(67`��Ih�6�5`�"Ж�hk�ΕJ[�b�o>����2mb��{o����q*{a�M|�ivqR]V]��4*�b��s]��A�kv�T��R7S�VѶ$4N�����c7q5ʱ عV �1����]x�_f��[k�a��)�	���}�VK3q+�;��Ћ�=6p̍��[�X`��q����)�^b��Eڞ,�h`Sl�N�9p���Mv���\�\��V&hO��tZ��r�� n��	��L�G-�"j)Lvj��(^��#�-�rpSonƔ`�0գjS��C��:��M��k�I�����rF��X�Uұf����5E�#���#n�a��L��۩⮀�M�J,ӷAޱH�oz�5�,��Rdj��n ��tFi�l�ot*H��q��1��M��0�xy0Бu��YG�K�m^�N>�Z�q�	��8��i�ۣ�9����;p}gvANa����[/Fjr�����'^+Rr|���H���
��/��i��{XHu�=a�{�|!��"Avy�����+Eòu6��լ/���`��Yҭ�S1`3� R�r��0�/1`��3K����kN^���Y�R-�n�!j�z��o��Y�O]�mkt�M�Ж���{R�.�8�zf	�n�8,���*��(��t;�s�ժ����=�$���M��JU��x �����i &��mJR.��><r��Ǯ��#l�K�Zd^^޽�,���$
��X���n��hTW5�O,!�6P��t���F��Kq�pl����W,S,N%Ǥ��ЖA*����Zz���x�[L���COR���6�Ϝ �E�m�k<�z�C2�G��1!RМU�>j[�E���<�����}����>d�E��:\�o��V�}�Fq���6(.��.�f*�Go��ԝ�8�����{]]�
os&�N[�*��ʓ����Kxi}٬ 5�vɱYP����J���+��
��ؗ���PWA��2p���ik�je��a{Y�><��#�]+�XuύL��M<������n�9H�}�z�842�%�]������PS�u�BH:�rM�k4MF>��j��D�0��e�m�V��'�zּ"Գ�qs�$��v��ݐ��+A�C��{��W�*@;{@�4�4�V�L;�=�!�����5��Y�����{@n��sȳ�㝢�Mj�;�7�y�dM,��n�ڽ�2���\�����W�Ulq�f
��S��9Y}��p�G{+Q�N��̮�����IŶ�g<�*�]�bQ�4�_V��
�jk�Ģ� 's
cg/�
'��1[���h�u��|�,-zNv��%wtX���N��M�A�+3����Hc�9��H�����!ĺ>���l�Sgd�C�V�^LiU�X1��{�0�@z��G������9=�q�+Ssr�4�2�b"�[���7֣�	�@�f�D�Ƣ�жv:�v�Pd1�&r̬��si�l�O��N��Rc�G�m&��)J��I�V�1�-P�~܊T
�u�ͷ+�]=V�}�����=�ɮX�}|��#T{7���oum'7��1�r��flە;ٍ��%b�N�}�w�,��;h+ݖ�]J;]�_]�e��fn��P����Ȇ��\PdUxU\� ��y}��vs��ҩZ��������Y��AkX�q�΃`�U��kf>�&��Q�=�s����F��E���{�+�<H(kmwh܁���ם�D�RۆZ�G)���z��x��,rm�&#�u;E���?�`���>�k:do���rw�vT�	�[ѝ#o,��gf]HvM�V��;t�l���R�H۵794.$j��"����wC��0��+{@�kg]sf՚r�.���K҆ FK�ᙊ�:H@�}�a�s��+�O7����%�z���1�߹L�o.lc�^nJH��clHx���Nt�ޠ�V��V]+�LhWO$d����՚8E\{���:uq�0iz^�<�c��sb͑�/Ht�y� ,!�����{6^)K{����n@�C+�p�D�'k�hbޏ�Mb��]נXx�#���]ռ���Y����q��(�gla�����E��݃/����m�뱬�[[�gc9r1�6Q<�f��k���`�HRd_up����AR8	Mi��@>u�q�.�+"�
]��M׹9e�
z׹�)ۤ2�e̚�b�l�Ko�Uf��z�D��u�l%'u�cO*�̤��r5m���$���vMy�!��li6KYR��'ٸ9��%�ۼ'�1� �(hɖ���DlV�7��`�}�+����$��>�)`Ac�%`��cd���o��QBwY��0��(��ʢ�u��pm�ue��5�M-�Rs�J%�Y.P�Zv�7�"��&��envv�g�v4�	�w)��Â�Rv�1�[�]5Ϫ�֍1�s�y}o������Һ.�GxF�ɡg3
H�9%ӫ�s�P놮��l�;T��|0U�L�(Rw*�j�\R0�[�m��Kq���욻�vu���=�o�`�/��Rhm�CCm�5�V]&y�n��<2�^\����Y��<������,�#J���70�k����c��
2�o(`��&�e�4�a\��:v�:���p�2���ݜ��º�]�;;)�0�km!eNti��ғy�Zfh	�&A�4��.X:$��#������S�Q��^
��fW=�|+.ވ�I`�x�hbw��P�jQZ�np���w�2��,Ya��� ʺ]MX��;��>�����::�CV)4���ޱ��w��,k���+��xksM,+���[hH*�]��S�X��t[ā���T���eԓ�����K&��nԮ�o�)�tf�'Ҕf��KGvZTku\�J�p*au��qwjv���҅�����b���������.Q�G� ��d7�S��I��2��)�5��ۗY��}��;���n`%��ᓝ[��|�rz�cީ��(�jC�jt��pJ�Oh(�Q�r�lzv�ھ�m^��(�ĺ��u����waYjk�~5x&-� ��pGX��=��f�=�m�ی0�8_܌�)]��Hl�c%(�#3�{,��z�tE�FY�5>[Y��AF��@�i�۵�h$� .md��əRJ�cOh.x ��!#S�7�2��fYO/@z�yAwv-�)�ku�ݣͰ/ln^g"v�'�e�D�p>�X��/.���ֵ�}ʱ�ν״��n�@M��Z�NJ�c=�:x�������4{���y�问��gKp�k^��B0���t#
�[�C�YS�Q�"�K�:�r]���b���U'f
�K롰S9d}�A�؅%��Ǽp��iԮ7����嬇r���[�[C^�;A<t�^�]�����7]m�x���u�6�tb�dՕͧ�Gӳf����,T9��ʎ��ƅY�jb���"��4M]�{���u�&��0�I�����ЫL����):㰺(��g]�m��+����MsNAk4Q*���Ŏ�e�8��4��;F�P2���m���gR��g.�l6�lws����q���f�ef��5�)ou�ѓy���Y*��ְ�E��X��Ǯ^}�q���Wj���ڊ�,p��4}
����]G���^(�3��:�(����v����nʶ�M�| ���sH�J_v�t�i=�vS&�V�j9�fMZ�{T��m�ՏW<�M�z�;G�o��������S=wN�O��<�ggb�Qc�&C��0��k	ͣ�#�e���_]u�a�yiXgb)�_u �YӅ�Z�ҥ��ʓw<�ݛ�eI2��"�U�e/�3J�+�u9�zհTE
�g�Rm\�+�,+C�|�4]#y�3'Т2�)�I7W"������ux�!Qڔl���-Dĝ���ޗԻķ;R.�
Թʆ��p!���������u�a�ht>ᵴLVʽ�sY�Tn�����E[��x2���1�T%:W��:����lt:�{Z�`���}�Y�;ھ�@�T��k��"kK�+F�n+Bdj��W���kb�Ρ�X���XC��T�_�٥_[�N�˭8�A�#���|�KF� ����(-q�:�|�����"2���S���a|V��V�y&��Թv�Ґx�jڃo�������Ul H��ӡ�wx�Z�</�7r`�0:WC��O�&M���M�PY����kS�-��듎7�B�9�M�[�����\������(�1���1�<�+P��鵝ۗG��
ɡ����&���Jׄ �p�0�v���ō9�{>�[U}u�;hTצM8V�s~����s[Ū�<(�8�G3R�ه��r����ȣBIٮ�MѲ�����\2�5#=�-ޘ�n]ڝ�5V�X^�f���;E 6�η�x���V��Q��)Y[�ؒ_]@!_2���w�lֱ�%��ݠx�5T����Ц.�hzgw4�Q��2b�%�_q�3&=��)����)pl��"����s��2�J�����KŦ�N�4��WΥL��C�HZfܶ���$+�#��z�gVQj��a^5N����*�X���G�GAN��١'Y�v.d!o����//�ùF��.\�ּnݐ:�������֝�M#���}�!S��ov�Z�k��`��_q�;p�l�E�9t*�Zd1��WZ0�<hr�r��WׇX��-� 9ɰ+�	 �Ct9��Y���z5[��ukf�s�x��m'���d��̠)[�7y�5*ō�ԭ_e��_a��Hj�R�@��{У��}e��MJ�e���F�W
�Ú�0�4o�����J��]����0T&&K|�����\���jב���5�[�6��V�&Sےe���岰
:p�e�7��8���eV2�H1��3�Y7��>�ᑕ����;s�[�쐹5q�����/JK��N	�@�p'Du[ɹ����ز>a��ε(t�;��֝�2E!nR'�(�˝-$r�hE�*������﾿�|y��;� {$P<w�u|qu-&�O�����[��E�U��7�������bbd��ږ���P�ec�m����m����{�-����v-���ݝ�wPܐ�a�ib؃��F���N �����ͣ���b�U�V�]��Z��N�ml��ոT�ipW5�n�T4R�r�:���X�r1:3��Ҵ��v+�7�Z���D�w-7��^uJcq�����G9���U�-��T�u�N�\m̮��k��A�7k�	Kz1���z �R�@651�ǭ��]���,k�8��x2q��[7� tyf	�.��EK�s�-��]�ʶ��Kb]h�WyDh��ļ��U��S)�h�~W�����)�>��OWiM+^�=�b]:9Yh��ڕ֬�צ -p��y2\Es��Vf�^iD4��ޝ���ҹ�p�k=E�� ��xsV$4}A彴��qP�g��నS���s^�[z.@u�._Ȅ�w2l���'&�/���Bv�w�����+�ݱv�C��^K�h�@`��,L����:��-�S���^g۔-�QbJ�#�e,�uyh�t�t{��@H![��C����Yt��'DJ�ǰTVt�W��V�G���gX8��g�5��%��^�f�_h��V�R�R�`��������3�i�})vl挵f�ЬV\]ײn��#xc�N���u�BR�d� ҙeH�H�#C@�f
䩒!Y*Rd�BP���H%@Y�8J�!��
P�
44�.N@P!����d�9	�fP�J�%9C�d�H�d!I�M��R�.Jd- �4IY �Bd����Y��9)�	A�a8@EPD��P�_| ;�}���rӜ�&�7i���s�L@NtW�.�Δ������4���e��8LȆr]X�W���]U9G7�)���}[��������ҭ֍	�j ZxkI�OV���{��칡;4FM�=Ŏ�5��&;�Q�#�2�\����J���T�*�o}�Xu�EJ�统&�^4�﫤�]���L��y��,�*L��|@�l� ����W���R�zx�@*YG�e���)'���:����D�<��ϡA�T�[�n���/��۴�\]��+lB���!�W�e,+OU��Yq~#��ϵ���B3����x�o6nwS�z����������1�JT�A~�W��V%�ʙֳ�P��yVVl�7��<��ݡ��aL�\J��&VVSi�R-߃?{����hGfJe�H�����|+�O�>��Nz�v*�L���0k=��j�>W�4�*�²rꫴ����	4�d�����z���x^SE-���ӎ��5���=�Q���Zl�4;���j��4�����+�2��Tv�WN�j�}�-�N�'}V����U�7���7hY�������[}W��u@�Zr��V����G+E���J�q�<�/g�Ɏ����e�b�6�[�S:i*;O�����+����IE�J��a��u���O.-�bX�XugP8-�K˔1C\��U���;����2��SF.�K,ah���p�K��U����u�	U�bf� �6��m�C�n���j���]X\Y.���WՇl�<$9Ww�Y"����^�i�Qg��5{�Z���w39�x| �rp�b��Z��t�$:�<9tX���5�hq�p��{�k�}��6�\��]<���?(ϰ��BK�Zx�@qa�G�??�v��I<^u6=%�uUO(+C9hn�������38/}�<5t)��t(S�B!5���j���Ǟ����$w>��9g'f��j9u��^f��70��0."+��A�Z��[���� ��bP@
5��U���U%O���
C�Xg2��D*��#�C�v����t3ɬ���@�Tw��eM�ѩ�B��Y�r9VXدb�b��z�B�t�$�+L�}=�w����!Eb^�)��e8�ЪbPe?Y񇮨�u�s�+�-*�ǋtX�!�,�����9�tD�����]Aԗ�p��!����h����G�K^e�#�#���.ps�A̫�:�z��n����xIWQ����6�]���B�0�O~[wE\�ې�]�h\��w�`��|PĔ� +�w��)�l֎)��M�/.O��W����{��17�;�@b�klN����L��i-_1ΐ��U'�U���C��R�8��N��M����:��=>��L�W��UBL�U�:_w���!��O�6�(���Y�s�z�m;�WƵ�y`����e
q�G���N��e�	P�]r��ݒS��1ux{A���C�]i�T�_`I��[�KS*ژ|=A���(�K+���͆�gu���k8W^����*�p�;fmܦJ���UX�^r�W{���e7�����2c꽙�}��C=}�f䫅LL?��=��Ė�J~`l����w2�oy�/c��O����e{l��R����Q�Z�PL�_]��Px��ƫK�#3���jԉ�]NKk$��H>&ɩ��n!���p=i�둱Z �]K�J���ita{����=����*��`ϩ���K�{e����Y��q���h�Hg�!nн��Aѧz�E+�h��˫�k"�|�SO��^Ե\)}'4�/��"�^�!G��;\�C���=;f���@��H
��Q��
OO� s��0OD`��z�˔�Ɂ���`.^X��w݌�Y���j�����A�7@�'���t�v�o3C�/�1�`��yL�U�����t!�HN�vS�Y+������4h�\��e�ɗA�M��a��[6��[ڙ��-\� &�̼ד0Q�E��gLFQO*>{+gt�z=���r��|"+�*�[	�I�gE�a8P��V�����2���)M���ͬ����nq������}<&�����$�t��}r�U��؁��J��
�;���8t��2����Ln�ԖEmNX�_<J�Uw�%��Q������"ه�\ǻ��e��V�;8W��mWwDAU�`���� �UY��3x"2m��ʯtŗ���H���:ȇ�o��?->���<k�D�4�J/���2������[��6H�����l�Uƍ���o��҅a�
�C��vy�n=*
5s����.7o\�j]]9�ZL��(;����t@��:a=�m]���0m?vd��;�����מ�����.�;���M%]�|�g��=�,�T���~}n�X�֕xM5"X��{=��V5��Ț�������~��zr��8q�/<p�P���s�h����@�\&;�d��&������2C�2*j��s����6��8_��X���ת�X�<���=M��M2���\#�`�s��;]�Fg�f�����w�m�cA��[����3�.�-����yݍ�W���|�Gvw
I�:��O\�"b�;�����v�R���\U���69���uN�,�{��,��N���$��}��:�V��ޏ.���X#6��f��=�ǢrΚ��5�+}��>.p#�ް�x?�?�U��]m���o�p����O���7F��R��^�3jl�x:�x�b�k����u��_,E[[�d��8�S7{R%�x��V�\��ǝL���N����i���b/�=�>1{�E,�"_EN�F��Ut�v���w0��5:�|g.�������dO[��82nB#���e�T6-nNO��I�V������͓ϩ��$���mҩ�_97�3��N^/sv캛��f�{��,��v��*�9=�c>V��L�om8Ḳs!e ��q�4L^xs��&���7���GG3ƕ>�y�ٺ���L���5Z:,S>�E�3��V��Y��A�x�.�#y�rMj���
A���і��|t�����U�zϜ7ƣ�.�b��>�{�_m�Ӆ�h��>"��Q���H��ܠ5՗�&@�i(���B�2��\;M�u:	��nUY�������W)�M�f��&�t�`Eh�]M;ʅ� ���Pi<���>�}���)�\>N:Ϣ/iĖ)��u���R���ٗ	Rhۿߗ��˞p6�~^�ܳ�'��O~���J�!1�#��O����S�U�;�W}�\�������G9\g;V�j��;��zTϕռ��uJQ�BJ]��O\_:e3'�gl���ޤr��s�m���wO���)Sj��������]Wc�}�R<!�q��K�/8w��J����O�k�Ի �������u��˭���33�@���:zo[�riO��8{fI��u>�2��w[`WS�\^�]w	sE���B�����ѝ}����zL����v������ˠCځ��W�G�!X3kb�Wҍy�;�O:gټg���)^R����ʄmw����)<��*V1���F����cd��o;i���{����^��K; /�Z^k�ڭ�3XЅ!ߌ^�vI�e����rS�p��Z�X{�ܿz��ʍX}�Q��X�	s��WvA;�6J1�.�60��xrJ�2��}]A����)c�l�]�RCn�z�������Nn�Nm���Ǣ���~�뗔=�x-�[Q����S$1�G�u�D�}���k��_o�M�_L����,/e�i�^�-�����U�F(�J�"k8�[�U>~��Cz����D7�kI��iv����H�C���v<���=Ҫ�pU��!{]в�4^Ll&fcά���-4��L��b�X����.:�!{Dt���[�l��gE?or�B}�|
ae���竳T�[��cs	�Y��m�.zx�=FyF��>��e-J��}�<�>�vT7�3�[ 7�S�����X.�c6>�Φ��=)��=C"Y�4l�t�)�ь{��.�pb��Mvo�Ƿ:��_��L�M�@q�kUu;kϼ��lV�K����G��Y��.bV�s龍��B)ƺu���VإRg��}j��]�I`��WK�+�du�y���W��e.;������n,9�ʒ^�~~T��կ�t����o�b�J>�w�q]#h	���W7N�
�I�l��"m�{-�w�_s�
�Gv�!��j�M���k
#��ڜ��o�C^h��<�)x٭�La;�N���[O���3�����Y�bD~j[3o �x���K�N�|�SI%;\gn=���Ǣ�zӗn*��6�w#�w����v���m�i*񦏊O�Gc��Z=��pU8��uAu�g�<�5��i�N���e�߇����K*�xt⎛�i��L�m
�gǟ#N-����l�c��{���[
 5���3�W�A�3��
�K��1���N�on�ao�j�{��쬼��ދ���tx;�����W��r�i|��2���;{/��T�U��i[�7{�k�́����H��Ub9T6�@�NV:j�������mά���=涏1���<������ݰ��*�8*�n0�j��\=�TU��Yh��"���؍�yp� �T-�)��hU�P��`J�좦T9�ԑ�O�{Ơ��]�q�3�+0y���yG�o'Y{������	�D����IG���·�X�����y�H(x�n� ��4���8C+�m�B��_���!{��蠢5m���)v@n;�|Z{����@��|�Y<�J�"�c�ٖ��WZI�v�y�RGub����*�L6S��u!������H���I{�r<��I����l�V����q�[��'V�x�3R�j�覒~z%���0��1��1���+�%V�K^j��{xM���/:��|���D�!�d�}'�s�����[��h9%�e��~��3��ᩯoZ�/��uA���
���EΙAȏ�m���UyJP���d���&���!苶�'Y�ޮ���=4F��{�νSϊ4O+�#�3MN�w,m�	WC[D�Ur�W[a=��%K���OSٝ�O5��v�OSc�}�v+x:��\���uY@,i���:YkWqiM��3�{03N��#�*����6i�
	�F5��	�&M黔���-y}�&lR�r�*���У�p/9�[��ܧ��=��`��Y}+$-ez_oN�j<����EՕ~�����q�P!��g��mtq�75�ɆOd���^���cQ���dY��[�J���a�/���	�H֦8�m߳���x�xi=ץvb�!�=�2��ja[v�5�We�X�ag��&p�u`mm����L�<��"]�ȵ��T��Ar���kz�5�{�<-��{� �\��������b)fz��%=�[QJ�[|��w=�k�i��U����^\w��hwl$wJ�	��t��/�ɝ�۳_.=:�pHr��N���E�ly���d�Z�܏��w�*�f�W�,8��Cw�u^|gJ��=V��E��B�x�e{���>ѻ������N3���8���g���/�P}Z�>�N��o�W[Ҝ[��k�������3�����9چ5��;�6Wz���ql}w��G�����΋�[�\��<��=*8�U����"�^�f�μJ�L�	������[T}lN��$�����s��E���w`��/�D��2�c��Ί�uC�4}mQ;����:���x䐻Oi��ƴb��>s~��ܪ'����uccD�Ur�}E��aX-����w�ֺ��Ts�����%���Y�^�f��F%2�۽�����ÖY���j;�wPd�҉Ÿ�b����+!O��h㸬,��c�9��Q���J�i��ś{p*�Aq�ܓ%�Җ��r����Ed��*�����9R�U��]R��k9xI��B��k7	���)\�r�u�]�Yr��il�Q�t�Y׀�j���҆�?+�!��D�]4H���kT2ӥ�Cj!y�b���"o��/g]p7�V�7�������mZ�ݑ��#]r��8p��{q���q<�� ��4���h��h�c�J���E١9X;f��8��%ͻ�;w#\h�r��îv/ڦ�ra�9�+v>\%��"Q����1��2�绔���������vZ��~�^5�z�`8D�]��,�����-k�&i������N���D�Rr�%��Q�j^��]�)h#�g���uv5�L�V�6�![Vj3Q:��c� �����Y�1^Sid�����]<U���u��J�mt�i�":�f�RI�nJVl�
�`7T�=��j����*ļюR�E��{b�S���e�+K�n�͇�4���M�N���iM���PE�z�B�9np;�2�Ua�������So*ã3�����H�v�#����V�o��a<���=����g�@�:s7�R��={�:����ZMj�U���{0?���[oPP��n`cw�t�1r��j<a\����e�睘���N^ڡIj�
�d��O]�U��'\�<H�,���:�oD0n��s#�b1�e���u���hC�.P����v&qoj�T8j�b�1���z�z*VR'�U�t��n��`���b%��pld��U��.rf�;�Ι���VR�5:�g˴#���Й�9;��3Q:���m� �Ř�tZ���]����o��j�WJ[}i���ۢv�t��ں�����^����KkM�rD"ń�n�9t$qvPW<�o��Rul��������k�Z�����c��n��\G�N�of.�d��{��x�
�qE�m�Պ���Lۧ�@�����c����yz�1\�y�z�'p�bJѴ�.D���#�d�����-ɕ٭s
���7��Sw�zÒqm=ˇ �u��_�Z��q�8(XVvZU�Q�2�-�l�@ME�IGU�(�l»yS�0�K8�˼ѕ��}Ow��s&T#��h�j2o�����ߖ�$��;R�*�i�U��h��i�N�>��]r�������k-W[��θ.2���.��6+�����W��^g7N6; ���D78_\<���s��dC)�n�:�:~Ԗ��wc�R�\��R�^��t������}��}���<���i
j��)�*JZ(��
 �)*����(�3��JL� �(B3ʀ(R����� j�����2L�H�(�J��JZ)(��
F*R��i��2)(��$ZhJh�2!�2

F���(�����)
�i*�b�"��j �
�(�����L�B��!������))L�
��((h)��@��i
Jl��((��HP�P��C�e�2����R���m7D��"�sY��Z:���yܞ7}�؜�o{_�J��ִ�����錽}vr�֮`s���ο>O��K�T�س�9�N�TCm�۪X�7��1������)�`n�[��'N�gx��q�}I�
�Z&\<�ݩ�$s��ܳ^��;E>͗����e�f�\�Mǝ�R.��91��>��X/|��"��ҁ�v*t���ۥ���6M��6�����^dQ>����fê>K����wU�몜�_[���!���Π穧ܞkW��6rw����q}���ޜ��'&���� 5�v*/e�o�N"�U�����s;��py>��I�c�z:�[�4^h����"(��Rsݝ�������(��'nC�t���m�2B�����3�4Y׽���k|g;�9s��{L�K�b�/��pU���B���{�lw���M�04�؍�x���N;�%�\^���E8�ŏO%�n{�#�yyG0���<=N-�d��]hH�:ƅ68��rAWgU�t������B���Ծ����ٯU�X%!���<���ܩQ�����kdK��;����9�W!q;
�F��ϟW6ڕ�: ,�n1���E�,(��\�?�:I��J���j�+�r��9l����-#��֩嫵.�x���o%�n��y�G!�l������O{{|�<�yE���C�`�th������B]v�h�ڢv2Mj�ݎݗ�h�ꑇ�ͩ��|fʜ=��UE�	��W�yr"{ݯ\���{�g����V�{N�3o#�%�Nɕ�E�#���ݱ�D�e\�1�aȾ'���_u����9�l�M{Z��8���m�\���ů'kY�����O�q}���η���4�\��n�x�L��-Y�-uk�^�we��J�S�hQ���|�9t��O϶o�"�+5�w��)C9<����+Ťw�i�H��Kڊ��@�8]�k�{mo�v�Ǻ�l�)wS��*�~�ϗ�{���r�c���:Lq	}���Ս!��2�XD�ۭ�k��o�'n:݆sÇ�%�R:O.z0f����^�_
�0����f%{�,gc�A22�ؤ���N�V�(v�ٕ�,�L�ή����z��r�3���蛬G����g�/���S6�\�j.�yNr�k!�|�W8�~���=^��t��۰�9��%=
��k�W�0�/�x�=���Uq7�
"�J-���*�����K�)�>V<�MH���O�o���u�����F`Џg�
�q��Z�!���Vb/*Υ핫w���}�MjmaX�4^+)�@�+#C7���Lz���O=�3����G�)�{^G�Uޒk�JߴE����M�N!ύ���& ��oN�[��1��e-�bW��{Z�M@��O��a~�#����Z��Qq���t�㜘ɳB�Bt�6[�u�z�����>�P�z�J���l/���EΙA�鵊�b��Έ֕?tt�u�U]t�]0{��lB����bbDDږ��g�k�T�e�o�/����)rv[�i�Z�W����U����UO|��YgK��,z1߁���羭h���M�:Y�;�ݨ����i�rUۘ�ףt��(<#;����h*�w0��E��?Bko��srR(�7SU�{�uv�D���;ImG��2�tY](��4�a��Ώy�l�}��#x=ܔ8�W�Ƣ��Y�[���Oo����Mo.��cS����r�5�nam��Y}�p7�/�5�/�Nȹ�0�p�f|�;w@9~��:,�����ΰ��B��i����l����x��t�W���#$�er�F�z�OH�$��[����gm�u�`�6`|�2�3=o\���M~Hz�e�^��+�ЏV�������x-폵��v�멟Hc3�ŋ��wۻ����i���D�s�nc5S����`�_e��t~�仔����a�]�����z�g�k��'A�;�J�KT�~������\+�>����x��`�:������>�	Cܾ�G�]���z\���A�����^���N�ܧ��܇�w7���{I�~�6�����*���߯���d�:=�AJ�~�z9/�R�P�' �����yן��u��R����^G���/w���kӭ}���������k���>��Ԟ������'����?K�+��B� �xr
G�=<ގK������>�Aپie�^��^���;�yj_e�{��2��u���}�}��߼��6��e�9�Od|�OGxC����{=Kɠ;?y��K�+^�A�=7�<��|�7�%�d���~�í�%�[�{�������h��s�]��k�C}�;��{���N|w3�+�e'ՐK�%���@S�Hm�b�5 �0wRqI�䃗�E�Wʮ�Gr�G
�s�ҭ3��u�q�W6+�u��:�^�@����&ʸTK\9ۺS�_uY���5���im��P�g��0�TT>���_��l������w/��u��|���X��?��Y�w/G�i}�r�2{{�w ����+�����w�ᮆN��ژ����}��Ҽ>���k��_iw+�ֺ��H~=���C��X��^GN�܏�d~:������r^AK����p�r:��w~���7���s.���;"�Y8���W�8f�}/ג;��{��]b��?b�Jo0<���n�b�G�w:�R������~����7/#$7���{խ^���w�3^��^����>�G^b�/�s����^IoI��~�g>�����s�.�~�����	�`y9.憐�K��XjW�7{��Oߧz�0t��ֽ��R�}���u_��ђ{����'>ҙ/$�s�^��z��sH}n��ZGs������ǆ�ira?f?A��
M{��p��<_����%���	@��C��}��C���'#��.���仼��޴K�y��>�B���^��_]��9n����4.�z9ޓ$y'��y�{�������sﻷ�］냐P<����'��<���=h�~�qԟf+���������=�����H��z�{������/�~�s��s����_�������~�~~���^yւ����C�P:�7K�����?OA�ܾ��t����~i7&_K�;9�����?��G�n������ξ�^��ޟ�����_a���h~���i�}hA�s�+�?o�.FH��ɒ�/�`�����b;������!仃~��?���<���s_��s����_~��׼=���N>}��7+�{���>�vs�L����O[����s��y����^�srd�]�u�]����_�M������u��>�w�����K=D�ǲT[t�I��Y;s�V_��eĬ�R7:@�Bhnhf�[�����ѩ�-o5�]\�P��ٺ�q�;��̒�[s6�R���?å�Jg�����W����L�k����d|��|z���bP�Tó�Y��v�5;���<����ܻ���iJ�=I���FI���rNH�9�C�(O]�IA�}���愡���P�������+���^]�xk�8w��<�~�~��>��w����bn_e?����{����!���p{�rW#$���)\�ޞC�(N����;���;>愡�ϝi�#�{:9��{���[�Y�w�s��;�;���������ykr��GGx�K�O�}��9/p�O��OR�k�h_ �{�����w��q��<惹7/��g�����/�_i|A����몧}��)�}�_�ޗ.��_��b=�C�����<����M��>�G�Լ�����?K�-y�z��p��r:��}��ߟ�����u�_w��W���8u/�����rr_oa�x���/�y�{����%�.�X��!�z�;��2:��nG���'�w�����y����m~�>�<�m��:��{�{������s[�����ލ˿q����w{�sHy#�����/p����M���Υ�z�>��E*��AT}�����M^���o�������2a�<�I��.�'��p����<��ϴr]�H�o��$�ܾu�r�]k�.K����K��F�O'��������}�7��Z���ÿ�����W�<��=����Z�=���w�����2zߚ 9��ϱ^Iٽh仼��y���y��K��Z�K�{)�����w��~�s�~����~�����:�n2_a�y��?K��Xj�nz����+���7.�$=<ކ�����{�2^A�}�縏�y���z�~X�/a�s�<���Z�u�\��9��prW��X�'���>�!����K��XjG�w?�>�п]~�r]��voZ%ܼ�����R�>�����_|�}o���N�f��� �_�Y@i�e[����Iƴ�]�p�ɭmL�cG'bŞ'�ê�I�¯��R�u-���(��g5��	ć�����+&+�S�����q��ĹW"fIwY:W^v�l��Ǯ	E
n�7�`�Ak��r�����y�W��'��y����/A���+�~7�K�P>��d;��������ъ������Gs�������ރ�������ώ�s��ߝ}���^��������׷��/P�����K�?�u��?���zi]��ع��?A��2\��M��xh�w�ߌϫ�}�޿������|��?~�#���{�w.�����?J�n��GR�#�ٽh�I�a�iyK�?�ι�yR�δ.��o�.FB��7K�d������߿�����p����������w��^���=�#�9�4%{/Pt}yr�~��<��,5.��C�|�R~��)�0A��#�&����i�.G<�5s�u�<�Ǟ�ߟ{�a�|��q���//���Gr��W��^A��Е�z��}��rr�ޞI�]��4~�pP�s�L�p�}�¾���_�e*�bz�?߄w����R��w���?}�������=�������w)��w��.��ﴇ��{�ﳐ�9ϛ�ɥr?oj������{��E?t;��'���o�q(<���9��R��o��~���\�ߏ�Z_.��u�r��Gp~�r�����ɸ|z�HyK�;����DU���"�m�?��v����.G����@�}�=ù}�����)<���Z�W���z\������FI�^�GP~�r>�ޏ#����^���i��/z~�#�#�\�}�p�q�����7��R>O�ǐ�rS���?K瘻�4��/G���^Kט>Y/��:u��y/QѬw?}��(�����ڂ���������p���=ޏ��}������C�+����y&oG�^������Ju�4n^K��>=o@y�݆���MS�_`#���
)�����=�~��le�F���9��Ҫ�9���Ө��Y��űd��/	���;�}+^�o�*��ݝ��,�"/R/o4.�h�W(��WL%� ʼ��(b��y�cI�i�1���Wd��/��D.�f"`rr�g����Wt��\s5��������=���:��/���:��i]�h7/ ����7/##a�ZGrrN�oG#���g�y/�b=���r�]���\���Wۧ9�^~��{��������k�w秿���9/r���I�:5�y����#�u��(_z�7/#!<��&C�wo�#�9'F���Ҽ�����?��]g|3��w�{�u���+���u�ܮ�u��}���2]����bI��Z�J��:br
G���7�$=|ޒ�������y'����{ι�]]���{�;�����ԯrp�t/�������δ�+��w�K�{	�1<��pR~��9�f�~�q��NG�_����
����s�&�S��?���w�K�|���iL���޽����/g;��K�;�d���y�!|����H����w'�0O`ܼ�'����~��/���߶����η���9'������w�h<���y��G%�G��h��=�Խ��C����vs�#�u/C��9#�?���({�D}��D}�������~���&�x;ů�C�_���W�7?��ݒ�G��}/=�;޴rW��3x~��>�G.C�>�x�/#�~����S�u\�U@}��U~�z����=��t��dw�}��y�r�!���y/߰����_g�p9jWq���R���u�������'%w�3O�w'��旑���*��5���_���u����^�U��x{ނ�������]>���~���kr�//֤w�x{��e仓�hJܽA��w#��:�4wC��>�T<�O�SQ~S�׍Z���u�P���&A���O[ށ�����~���K��<�?b���!�X;��|�]~�仔���a�]��}���x>��Q�}��I��R��_����
o�>)�W���0ů=,�8�^j�ع���=�U�-����p���b6��w2>�M��⏳4����t���;L��7��.P�zu�Љ�v���燸��A�Dm.ZRbݪ.;����־s2�ci󾮑н��$�k����������߽����\�����C�G[ގ���F���ܾ�I�}�	C促}h�+�:��.]���-/;�2����ϱ:�r�u���_��5����sW;��/��vw�����<w�!�u/ ��䏒doAJ�s���AHt���>�A��4%���?+�z>�K�r���#�伎�ߛ�˿u�X6ZK#[����߾���p��~5P}_H�;�G�ԿI�|:�HyK�+`���<������r��y��w��w�ie�_z�ay����3(?f��_�H����!���XC�}�
��%�'�=�����y����R�h�y��K�+����9[ޞGR�Oo���w��5�K�W����f��/�O=�}S��]|��E�!ԾHy�C�}�u�{;���䯑���!���A�w/��i}�r�2{{�w �[���W��?u���}_�!���}����v��J��߯�x������:旒�]�K��!���!��`>G�yk��&G��J�ޭ%��}�!�;�"���,�����V���]㽕_!_w&{���w%�7.��y�t}#�����]ޚ�K�{)�0<���n�X���]�F�ԯ�r:?`n
G���~o�T����~Mj��������G~����#�y�2^I���r��vf��O�˹|�֕��^~�܏џ�r!=3��w4?��=���I�}F]�è�.���1��!U�V>=�J�p=���^FHu�t@r^{��>ҙ/$�s�^��z����[��y���}��u��_cz��}�������Y�>�/�3#��j����>�JC�<���W�~��X�G�_����ܻ���z�y.���H}��z��^��^�ހ�{��|�w���?<��9�ӟ��B��P3�}�{��w0����Wt����^`v��x�Zz��k���ԬȹU�,X'��+(��)՛�)r�B���;:�a���}��0'��H(E(cg��",��b'x&��6���36��@:0����O��
1��8��}�w{�1aq��g�2GR�hr
O��K�)?�}��zt`�C��O����z���n���G��;���K�U%�}�����_�4Mo��o��w.�ç�w��}��?\z�B�:���)^A������Ò�2_��>�p�=1��~��r�.�~i7&_K��_������~�����I�_�?O�J�g�>�ԏ�/4{/P�ٽ�y=K���:�<��y�+�<�Z\���7&K�d��p���t~�w/���4��+����S����V��,~�s�|��I��y#���4w'%w�3G�w��&A�|��w�)�=��w���!�X�߹�2_��:�.��ߴTgߖ�����\���g����}�� xue�^A��J�=I���FI���9#�����;���|�Pn_`��`�=ÿ��p��.u��@<�^{2S�!�ػ��uo�t������#��p��w)��=�Kܜ��ﴇ�Լ����\������)\�ޞC�(N��=ù}����hh
�E}���k�S����:j���W�>��b��/w=Ť��]�I�^�#��:�r���G��{�rxu��z�s]��оA�:}ގAJ�~�z9.�%��Lp7����o�����'������xQ	�w�=��^�{��K��z\���y��{����X��y��M��}ޏc�y!���/�u/ �?{�^���]���?�C��_�?)��^����9�4n]�Ju�4��}��Ǜ�K��u��C�0|�_��:�#��z��c�_##�u��7#���I��UT�y~�`>[�p��.Iw��.����Ap���y ���rz����G%߸�~sF�份�îi$|�yޗ%��~�]I�<u�y?��t���+�U�����%�Ю�F���m�_��ȗV����e�%�Z���1t��צ�F8����n��|�Z9X���Jc��y�1 8������J�TB�H������a�}�&s�"�cj.7X/���W�F�4�ju�s�Vs�l��/D�n��ꔲ�Z1���];XШ[v5wv^�W=�"��;�H4	i���d�{,?.E�1��cfs��dP�� n�N\�4����¯ b��liص@>D��ۖ����oD��ӤnY��ս/jgx�+�u���±��ȶ���fU����k��f�P�-5N�Xw�_P�O��]�-�7M��ڢ��u̖g$��5�V��~׻�>KO���b����o�v��A��]R]nb#����9;�2	+Z������Z�������L�T-v��(��K�+y���k$�64-��"�2�,؇fNg�Z�V����.��H��-0�w�47C[��y�ֆ���v�wmZi^��q�*��rj�F!��=�;�� �M�WN<9p�W���a搭V�fEÆC�|8�����(�	��xiKܫqP7w�S��*�Ҿ�o��$�ohlax��b���!ǵq��Zm�ޠMg-d5Qk넣a�0p���N�:m����P<0��a��T]M�Z��(D�ЬܭsF�4����v/�_7WM��ݴ��ִM^��D�:�n���}؝����X���-_G��K�v[��A�stzȯ��O@�ZSaѭZ���nƵ�mh���b�yM�s�U�Q����d#u۝jhw���^��K�L{�\��޻-�P;�5�a��Og�E	˫/\�P<t��6%�;�[{Z[�X�0���ݻ|�M�Op7��CA�
��P�)*K�Y,u����6�<7� )7D���+S�� �X.v�Zd��r����;E)Bw6�,4b9Fɍ\���/s5(J��N]�f�Vz�Gl���*[�������\U�q��-���lq�gIm��c�� �pJq�����[&!��0��حf�Հr��ot˥��+� oP�S,.�i󵅚u�+h��[sΝ+�n^��/:,�'8�˫Xm`fc�>��ǫ�����y9j筶�5�;e8�闗�; ����Gf�����ĕ��k5�\͎gM��1�ƅ�ٕ�v���X���,��%�}n�6�I+�m�U�D1p9XU��{��]��KVR=W�c�
��e�N����}�r��dn���|O;��="�n0zZ��+ؕ	Y�L���Ӏ[�%<�*�r�Klӧ�q��oSw��^�/���䔞�%[��D݈\9�[G:9f��|��}\�)j�.L��VF*�sq����eF�]_�_!8qd�����QR��1}	1U�}��?mq9��u�w�/6�wf	:ѾQS�=����� ���f!AMD�I��SCY�C��D5@P4-4QMKKAACLFJd�PQ�E�&f�e�b䡑��d�IE%QT5YFXf1RD-P��%UU@�1�@d9�DMMSY��PL4DP�5Q�Y�UA�a4P1%afE!fY�UD�a���bUPXM�STMTL�AVX�TTQfMUST�FT�SE%E$EAMQ5PQC�M5T���TSEPDEMe�ALUEE��D5TTE������u���}�ee9w��y�9�G�W�A��һ8D�]k=���ͥ�t'`�`,���6�ַ�m^U�=�����3JnN{Ͽ��
�y����
��4�%�d��t���9?�y'���K����[��ۗ�x����]ir^MV�
�t/���_�>�?~ܫ*~s55���?OR�u����_�>�����7/#$:��r�2w�4&@r�ޞ}��M��wp�/�>������}�W�}��Y�{��w�߯�})��_����)���2_!���p~�qӬ5�����ҿ]~�n]�Hu��4����vs�)����=�K���o��^��ܳ���~�]�������+��x}և%w�~���~�7&C�)?f	����kH�������br]��z�փ�w// ��iJ���R����[����[�krgN7#��;kx:��
��[�� ��Bhn.y�cX�ws�od��$73�Y����xAty��w֌��޽���&�윛Ӷz��<����Z�\�J*n�U�p�����n!��<�\�:��=9�������z\���B"�o�݄Ʒ�j�g�ƪ�؋��µzO}Қ݀lr<�m��@��
�Of��>��}�^�
,��#U4<>zQ�IE�ݰ��*����V�W^��tX��Vʁ��*S_;*����@������ٷ�'WU��N�z�h�<�m$�=��]���/�.Z�׋�w0�I��V� ��Nn��[����
�sDXRWoq&�s�<���Ԉ������h�;�!ʑ���+<�o1�a�����:�wc�O6x�{X
�˝����6��hܺ�-�{i��ml	���>�8�d��/d/h�
�)���Vg��9\ys�',����8yA�d^��8|�u4��;�qف*كܳ죖��C����LKk�T}���<�@��L��an:`�;m��5I+j��<�5��7���l9�7�˨��GK����ҫ�"q�^W{%����wϩ��� ����>���'GPp.�l'�:[L���v�}Sܗ�k�޽�s`�_5�6�����D�W+��u&]��.���똸d�k���z'K�v6¦,Vǃ������,���v�ϡ���_�c����WӪX�L"�C��TCo�b����k��|}~"�F�
�@���\F�g[��i�_>��s*)��|�;�اUS�8~	T|;w�[�(.��qo�.�i��C:�C�A)U��b%}��[wΑ�(��5sc;37� ������Xku���v����Z�|jl%uK�w�\��Y�s�G��s�6�N;�wA�)Z��e�.���d;��u;}��~�������t�<�����ѭk���͙��Z��3}2.W%�ùa-�~%j�(*2�!G�=:����6��V��u;OP�z�@��n����V����+P	��6�R����Y�*�.�n���9����N7�2NQǫ�c���λ�[ǕQl=W�㿹.(|8�g]�yy�Ow<�6��I
�:NSкo-��h����4��j���=�>xzn�|Q��v�;�k>�Ys�H^�V�ec,��w����;�9t�,��0����^�c�)��X�u�"���n�y�Ye��<�n���z|�{��Y�z)��<Tc��/�������U�����o=�U�P3�Y�Us�e5K���3�Z�z�yڮ�����do�����>�loJ�=�{+/x[T}q|_�+P�����^�l�S�{���^)]2N���O��vy�5���ӗ$#<�{B�ݛ��Y����+�컁���uml>玏H����Ƿ;��L�>�,1���;�n���<���Gc�D��tZ�e1�}�%>��5(�a���=���ц�JR�u߰�ټ}�] v��� ���u�(�p|?}�"�����7��W�ōχ�k��h�����|W?a�r����/�O�z�%g�Tnt�s�Bu.�&>��?R�(��xzA�,%(���x��7�t'в��=2.�R��D����}2��w��#�Ѳ�9�۽^��j�ƺ.=�:�E�8�Ӻ��8Y��X쪚��n߃��{k�bWX�[�U�|�t\�;���fy֏@s�m�$���}&�b�]x�%�5MإU�Ag�#Oml-����z���;��}����-!�z�k�/��MU2����9���{�ס���;R�-��}+]rU9�����/�R�NMU2�x���OZ}8-���ZZ�\���u}�LݕZܞ�&1���g@�<���wf����!	q��e^�<9$��(�ݹ�Ҫ�pS���:u���}x7MUa�Y@��4ݚ��p���`$`&����'\�V�^�KF�U�:NB�G���q�4��哔B�������Vh�s.��}�euΜ�H��L.�F8�Qw��R�ѱ��X�;��j�l�j���E�M<c�����et!^'꯾���Fd�HߩR�	��~��SG��;�J�����읮P��WJ. ���Ԯ�o����ͮi,S�4u��Vg��8����5�h�,�S�im�p��z���#�m�}��G݃��J��ٙ��G��vU�Sgn��iNl=[I�z8���s�
8��3+8�[�+��N�ߝ�/adq���<�v��Z�r�+>z�9��F��9��;�l�үw�����5��>�A쫔kPp,�l �K�t/ѮBu-9�Q|�*3��S��e��WZ>�o�	|a����&(�r��!�?'�69ݍ��ٺ������S��C��d�U__q�6����\컑Vn�r��Sl�o�m{o{zj��o�v+x:��/�s���t$�"��-�pgc�\�4%��9��&_{02��<7�Us�����"*y��M��r~�RѬ��me���-���ҎW���4ڻ��G�y�`���h5�'�릺�z��_E�I""�~84�稝f߳N�	�whWq���ݽ���s��ق+��]���=X:k�]�zw̽�ּ�8�y�ͨ������������\g�������S;4��O϶z\���)���\�J��m ���ԕ�I��u�%�k�]��O7/ ��u�������Hnv�o��p0:G��í�/#�ͩ�N몛*/Ϭ��R8:���㑙�c�Y�nގ����n�L'~��T���ҍ�`��]�	��Uvq�+��\�����T��l=�w�x�y��[+;�]�O-Q��E::=��|�s��B��cU��L���V`�0a��e-�=��IVÓk�$��i��/T��Y�N:�Z���M)L:��p�T^���y�e��Pnާ��r�h=<�8�s�kt�ܿd�4�NQ��*���q4�=�t��B:_w�����Ӗ����,�\����zR�v�Ã/��m\Fp�N���U�����P��9�T�j���A����w�daʗ|�ںͨ�	8�c�7x\w�e�y#��y�u�Γ2���������b�Kz=o1u�����솆4ܷ�w2R�*Б�{�&ZK.>d����u��$b��R��G8"k����9@�!�+����������?7�MF��v\�Ά�ʵ~�3�߇�J��j~�I�z�����-�szw�${C&{C�6p{ݟ=���v6�e��ޣ������gf�ݵ��Vv�6uG3z,����|�n�oI�m,��p�v�sI����
d�!��?SO��7��2LY3�x�.���w��dOO�-We]uX�C�Χc�Mu3����!���t=���}��Z�=�������l���ׂ���g�r1��Q�������|�oZ���;�u;�@�K*�5�U����GcO��RM٬��$sf^��ʑ��?[%=Oo�.*����Q{�_U�������!A>v�ø�$�HҪӓ�$�3����+yo>�E�Bڥvo{ޤ��gV�i3�ͲL1�ǽv�*�.h�.t��2����l5�f����лj���Bd5�7��uγ)l�� m�=D�5�{�B�{�)on��f�n��:d�x��"#n�.�}�\����^��D:��Z,6���Q�Q�їՉU�4���79J(����7J�I;�[��Y}��ޞZ�`r���y~�������T�6�fo�^,����%\|3V0_)���㬈���lx�h\�d$��KK�"���n�S>8�q�`���cs��w�j��[>��Н9�Qo��)�V;h�H��%�]��.��<^�n�3wۗd��N�y֫�� �zTq��<,Z��m|}qQ|/��/����7�^ꋟ){1�k�[Ø��|\�3'����/9�(m��|}ls�D�df�x���0^��=+VER۝�9�8{��>E��
��}vӝ<��78h���F�_`�n�5&��.׆Nfus�w��o���9H�Gy��,_ye��l�<9�u�uƝN�����Dޠ�6�K���_�1�OT��{P]Κ*{>�}��:�V�Ա���{�OT�;{;���s�Z�4(�]颹����e�1g��ǹR��F�N��3�]�MlX%\���YN=ԡ��5�sl�Y���S�c�λ��c�E�r����1���j��q%XEN;z�-�Y}Irʥa�YY�����:�%�2�)��:�o �a��'k�����^>���	*T|����}UU_gDzl	H
4������q�3\��}2n}w�@�8]:٨��Q��h���|�Ǻ�����Hc�椯 ܛ�Cq�U_m.��J�87J��[s�.��=�hk7eV�'�LcG@{!�*�vV��v�Z�}�v#Egi�?t��ǽې��T��q���x�6/oӬ��oŬ��������Ƌ����̬��w����Ik;���+s�;�I%_�cw�8�<��捗��e=�q��%�i�t��R�v�A|\r΄㨲%�G�٥%V�lJ����A�V�y�@�:�d��ա��@o\�/n=*8��3+8�wN��ud��#�ϯN�٪y��t��9S��=s<�Aї9���_s��\�ǽ!w���M�0�����{�����NQ��sU.9пF��#ǟN�b��k0љH6]Cmo5+p��7�����Q/���@?P�$9�������j:"�)�
ld�9�
u���}}f�0h'���-9)%\���f���A�؎�voL�Ὤ�a��]���a����3_Zk����:Θʢ���YU�߾������K�o�������R*(m�<_��֪���l/:��D��L�������r�U흘�NQ�v6����y����u���z���yW�z�z�-G�֕ť;��ů��8C�*�6�أ��ut9�\������x�O�{=���DF�w�s��Hl��S�vУ[�7oV�s��*�;��f���ݷ�>إ������b.L�/~��w)Gs�x�����O�ʪÅ��j��ٰ��m������d���v�3<���f'm��(������P�\s�e����E�<�7eTr>1�F�{�����}5N�^R�]��Ʃ����G��$����x��z�!�ص&����꩏EX�lg���t
�˝��hFy�G���AVze���K�p�U�Q�oM�mT�.uI�WJ����'��)_&s��eA\�jFd���s�[�@�M4p]Z���*�5�K�I��hwvr�F����v����1�6̾\��1z{fV˗ӹ�I��{6.@o+�ͳ�;��e	5d�C-�4�>�@.pmޜ��� �&�؃�[V�1��:�!4n���C� �FsHHK�Ъ��79+��WvΊ�%	�xv�P�\���˚��X[�v␁D0�����8�vu�M Ptx�CEb�#躟̱FmD����<+݇��~y��s9t�(��U��iV9�����Q�����q�;pW�lt:�٢���V�@��z��47�n�^�+62��\3�(�)(�8.\�:0m��VV��m8�]]&7������\o���l�t�f��L�g�و���A�#��MZl�)�`]�����sfJ X!�5��3��J�]����ј�u�&���.�g����RiΩ�!%%�k4s �o7�j�w`<���6ݐ��೰����:�න��M�ʚ���]\��;Zn�<��P��ά���)_k͚%ÌRnJ4�n'�s>h,�d��	�����E�-'�K��Kqvl&����4�ٮ�tv����{��Q
ͦ�񎁗�����g��I
���^ �ٸ�<���E�K�;Q�X�{���N��Y���iWK=W�!�sh���{�1hSSyl\]ܑ�q���|���%[���Z���\%{=t�y���p�X�:O-�y]����ד��ό]�ѕ)�A��O�ԤaS����/�6<e;y�M���톆�M��9´�BV�O����U�#�y�Wwf����9D������mc͏G�nhⷮ��puD�&��.�dU�n2vl<_mhw5}�jܙ�|8�J>:����U�DR��0'��w�U04�r�j�R����v���pxw�����v3Y��)6_�O�s&�f�99j�k#OV��yO�\띾��n���׶Y�����c\mä.*f�d���5��aN�#n<Nj� ��m�f��M"�u�f�@��͙˴W0�:m-�p>�St�tbl�K�b���i�K�D6��\"�.L};�[i��Ct�i�ֺbc�K,�t3j����_fv}$����F�k�iJU�4)�xz�|�����S�rU��5��J�x�}7E�_�J������C���/�����'t�z�+�#S�Ia�xM�N�X��'
��搦�c���qdۭ;��Xd��M]��V��=��zu�$7�ؽP��k���60���ڮ=�u��&���]}\�:軑�P�Oz� vP}���#�j����D���un�v2��W>��{gN:��4k�ܓd�|,�4�U2���.�"�;э��B���"��Y}S��&4����#ҙh��,����2�>�v���ú�[ݗc]Y6�o)��Q��so$ו��;'Nر��B�9H�D9v��|��w�a�ϳ�t���2"��j���#,�Z�̨�)��`��j**��*"`�"�*����*���������(�J�����f���
��"��B���*�"*��*��&j�*�"��I���j��(j�"�i��J�J
(��"a��3	���*i����rr2��bZ
�"',"�"��(���(�)�!�&!�"���"i*&h�

�������̓"J����"h���&f*����$�&(b���������bZ�(�)&�� ��
����	�)�
��'���"��+#22&&j�����0�b*"H������)j��#3�Jb����Ǜ�=����_��ǽu������x7�:���g8��ק��vEJ�yK�*vr}4җ����8���=�ݤ���۶j >����9]�˥Z���{��
Λ�l1z�}��D^�s�>��53����]���
;E��;at=�Q����ju�풳�ވ�����Ӛ-�(�s�piy{����-�0%W��� �Uc�Ϲk�F��1�B!纹=����n��;z<-'�;|��Ã/��lx�Q�.���8;��^Z�,�;�vuÝn�;�!RLB:MW.h��������eq7��Z����s�,΅v:��Z?M�l͆��=���v6ǃ����4,��\1��/���n�|:ܧ��Ӫ\;��x�)�	����v��1��ϖ�5͝��e�Q����:�����NϢ�p���Mb��z�Kv|}kn�ȷ��Y��]|��K\�gMb.�kʻ���#ꊈ˻h)=�.��׳�9i\S��c��zu��ͅ��lO�~i��`���:"8H-_&#.���(��R�G4ݱ�5�oJ3�G�A���w[5��c�P-�\����f�����fe�m�w�9�<:�<�[�Z���n���a�u�9�24zH���ʢӣ���l��k�������՞�YY%l�-~�������p���G��(�K����ʊj�eK��?k.��j���c���u.�ͩ{�l�G����7��d|'��SюMτ70j��Í��������h��"��ީٞ��>U��~�I��/������ec;�S|�VL+p����)g��<�I��F7�ָ+��/h��)�&�"�tX����׺�����iO=
Ì�q��X���ϓ��Y�w��M�>�&�Ů5>׻�w��x����������L2��[��3W��y�n��F���o�?j��}���H��'`.��L�,O�!F�)��6�+�������}�ގ=�Ƞ���m\E�+����_���Sݽ���4w�o��S��8�yi�ή��U�Ot�Rv�ٵm';1j�׊�:_�8�XVER�s��6�R�O�vR^o�H�.�i��.4Wqh�^�<�����U��҂y�����Ax���y�^- �u�vp�e��f�y���s����wHGE��e8\x7��+���������m.A�SέGXOdy�0��X��=|u�z�[���U}����z��]�_����F��a�-�	�5N�C���9�����V��os:t�i�>��ڇB6�:Ѯ
��_*���Jwk][�y�f[{��d+Ӻ�-ORo�}0HE*��|+�.볦���Í�<�^�z��Ӓ/,�~��ι/o�NI�n�*� �S��J��y (�����nhN�Y�k�G5�T�����%���)�e;����
��ƈIg=�%�f�9����-�z;0>u0H�(o��p1�?�*��Ѧ���nT�r��	��v"������]Ku[�nB�N������6�7�z5O>ݛZ9g>F��43y�ΐ�X����@�W�pQ�+���"�)�������D�/h����h��T��-�������<C1d]霰���Kxw��ڡ\�;�O�m�}!{]ߴ���u���ٕm}����*0:���w!�}�c��6*����2����b���n^W�S�u��4��v-"�Z���W�I�\j­��^x�X�������\o9nWH=��b�V2{���ܝ#��ܶ��Xb��܅������d���78���UUWذo_�����<���1���g������J^�؁�RY�L�)��a�v����[�-��)���q�r�K�����LN�g{[NЌ3����h�1��ps�qL���>q�}_�>:��mL�v���+�R���p.tmp(�U:�Ԗ��Ϻ�K��v�Y
����ݩ������m6Ǆ��[_�U��m�f\��*�S�8Թ�dI��u�g����7���dmpzFO3��ŕ��$��	f	�H3y��Z[��kY��؜w��)V�s��\�s��l�4���Y��n#�4� �n}'3�$��=��w��n�u-��
N޽��I��Py���}�ޘ��ж^�b��r�o5�_�����剶�ʤ�5�Atzu��ͅ��V��q�?t�����l
їQ����eX֔�GS�#ڜ�Fiͱ�{�{����&�	r���.ﲮ�t�X��f[ֺjj̾�p�vix��ن�g.�^o'�*)N��1Q�l���n	]-&��m��R�U�}��^Z�#�yس�bC��=I=�,�[���������Ν9�51ʿy/�:�b/e��V�H����~��=Y����i(�]��`^�Ξ��������=zQ�J.��:Į�����0��u�O�����7��{Y�+ys/B���<�MŌ��랋��j5��p��C5d:�ָ+�H^��t
�)�X��w�7�%�E9�����٥g�5�� ^������D^뛥":��Ŝ6������ԏ@��g�e5K#�8�0~��{Ҝ�M�]��5�g�{&-wO��[3��R���)����`�Tc9k���;�yy#Y�q�̆T�Q�K�[y>���R�7��mU\����89R�Jz�G����7�c�z���^nQs�'���\�ClxF�[UD�\z7�=e�C'N��� ��g˄�ͩĺ�k�>�k#k��92��oj��9arF�;��p,U�/�P�����о8:K�WZ�;6J0l��; �|rކ�T|����/��{0-�т����.t�zt�8��c3+{����}����(��\r��<p'4K�}��q߾����7�7�7�usΪ/�o\u��5|'T�!�y3{;�)�}2����"v#vf�����B��ANL��c:��Ѧ�$NϢ�p�!����XbS�=��.횗����Q�]|+��}��r��ƫ�TYjm�I^h��]���BY�C˖'�*vУ�p�ӭ[۬�Z�V�/j�mCG����	7^��Ӭruދ�"�ܞ@@� Q�]���-����&K�5Y�.Kj���Ϭ����;��:�������\Y.�خĵ��_��l�ۢ9�j�����I����B�{6�w��C��O�b��0�D.���eR��2U�m`�BԖ�u�܅벌� *41z>����G��}��s���E]AT���&��]�=������SG�����G�QF��T�I�
��<x=���:,{;��Y^*���m��}��U5�GGx�Zv'�vv���.x:�������g�ڠ������7^{��7��Ԟ�������@:�beo�,\c[�[ťt���Ċ�
�v���V�,�Z�n�tD�)����q�um�k���=��w6:
�¨l�?�a����h<��?���/��X�։������u>]���\8�K�}_W�F=�i��78���[(xg�m�^�Wi�wᒺ�!�}�)-�y��u�MH=�[/4y)5�V�LT�?O^������н9�����Pxe^�����1���0��؋֊�]����"�^@�P��0��5�}�����SO���*]s���~���B�{h��i��&�xt��L����@7��$&مS3�L���\b��d�{C�l�[�w��Q>�i48ω�=AQہ�x=�)�!#6j���S������/>FOl=����I�N�}�x�*�s�L\���tO�/��f]_��ci���}pVw���猖����g>-��r��Q_	a�C~��3�]BP��y�ʺ���徬j�jVJj��㏽ w�B^���K�$��c���OF��[�@V�ق ̧$�k�b���������c�UvQ�'��:!��_�#�"�:\E����<�^7��*>I�Ƿ�r���w~i�L��R��o��h�'���W�z`�Wc*Bl��I�\c/ "*�[ v`0,�;e_o&R�Ȁ<SU����:W��}�3Fڰ��X�WkvSqH�{��\df��Z�TD���	���c�����I��&�W���2�.a�G0;Y7� ���,��;��{$����=�U.�]a���F���U}��<*�M'�H�_\���Y:?iC�_�����4��L�C��x�>dR������^~����C8�?�%Q��R�a��*�V�/��.�9�tD}�g""�%髻��wX�p^o[�� -�q:��f�t�i^�����n��J2�U������Wl�\����ׄ[�B�8����s0i��T�i���$]�鰪|uߨ��]�����"�$%`�Fj���8�97��c�0{޲��E��EN#��\������v����Y�U��� 7��		|�S���O��n��L��;o������t��|.���VD`2�Q ��:�YS�SH;�zc�a%�	������2����];���>E��2�[�u�-�G�	��*ofR��8����GǓ�Hm��6�1{�&\>��x�:.���d��Dxe���&����{���âF:]iz����yV�
=]����9U2��U#�`��xTTH�dm܂�r�o�m�H���=c7Wbn�CN��;�+:�]cjJ����Ӌ�=μTq���rrkt��+
5p���5t%��勭�$����@ep�n����9 ���P$&r�;�g��ˡٵ��m9��dM�7��w��| Sp�1�s���/�d=�B���$6`t�{)ys�x尜�#���XɆ�Ѷ7�M�齭ns~|�z� ���$no�Fp��/�3,H��q��"U�r��؇��;�{��'y��	^vx�w�3�t`��n����s�Q(5�}s��&����/B9m�HC��>�����+r���x�7��d�`kR����D5�@n��Õ(�7]r��7�ւ�|���h�Ŋ�*�.��K8-�)r�旅��0׆��j?��T�+��M��ql�ogg޾vS6�$�� �v)�]�]5�sć�7~JCYn��&��3k�]f2�������݉�$���Q=^y(���UNU�&}�`c�����!�bkժ��K~��i�Ay���#�֯ �x㽤����5ծ*�s\�Ey�d�	��9� Ыf? c;�=���α3}�nL�Lw�A�����#r��&T�{��u�#�/���Tw��f�՜L�:^�:*S1��YQ��ӦH����
��)�F�-�&&}q!Y��%ћ��5ቿ	Y�V�����e�3t���ks�e��n�@�PT@>�48T�լM6ND���Sa�Ze�[��D�ChZ��0^:�8���g1e�,�Z*
�.��gqr�:ݶ���H����.t��Bf}-^8Ș7���[vYS�W���JSӭ	�ϋ�_�O��c�}h��8K�#����+�����P�����z����Lk�����[�i���w7m��+���*���b8�:>U��P�j^h]�,yI��akF�&6-�r����ڜ`�qW��P��b�ʲ8��2p�	̕���G%��m��C���9ơ��v��n.��=���0�
�¯���f��JE��/f�/�a��j��<�v+�$�9A�34���aS��a�7��p*b��nvS����s�]�D�@�MƐ�Tҧ�W�:,�=r���f=0^�����^=k^L�3�J���5BX�x����a*��f�L����X8�{�Q1����wT�ͪT��:�vD������
v�
:��$t<��c���,��S�q�g^�[+2@��"�û>ҕ��xA�S��� (ֻ<	}3l��b�00���gV�L=t8����v;�}�2���i�B�� 0mt��TĄ��6��{ ��[�K'.����<�1���&�;M�xn}��8�G[��Qi�ܘM���ێc��VK��a�=�\�4�;ׇ����e�l�`*��<�!���R!%0`-�� ��c� �8�I�U���q_f&�u\��Q/��Y�n�b��{K��"�Vj����c��.zo�תعW�,t��l�id.�\�o
��j��wǸ�v�fJ]uA\͚��#*�|�W��o�=KA}��]3U�+�ǘ�3g�H95�c}��J�@��� cN7�p͖�����*ΝW����rk���q����<{4SS;>�<O[�6��׮����r*v��kӇ-JuW˄�ڹM�9P-�pVi�ҳw=��qDj��Q G0+[��(�BȚ-�g�o��:��~yV�t53��{�76�%����M�g[!d
�D�+�
I��r��Ec�Ec�1��Wr<Z|ٜ���Wcʠs7a����b�4�1SW�ޭ ]�Ƀa;�3h���7�]&�$2�֜�Y}0�W��Ik�Q�ɒ�]��R�ӄ�Ј	V�nL��m�z� c�YR�+���8N,�6�<������[}���@�V���.�ۏ�x���]�bd�	�ĥ�y�s�8s�۾�1+8�d�	]��wм%�Ξ$-N|()-]�sC��JS�ծ�u%Xu+��+��8�� �@�SV�;�.�G�P�_]b�T�FEi���wq�/$X�y
�{���zp���ެU��.Mg)��W�#2�=�[ǝ�e��ª����=�X�G���6�����U�m��������]�ea���K�Ηo��h*i�D �+���Ab���x�7gsl�I�p�67�s�O���d��wi���}��̺7�E��&,�f��Jם�i�o��X��}]r�]�ٗjGr�J��ԒFe-k3"���ܡ�0��;VC�1a�v2%ɷ��a|�*���%�38c�*��_����.*��pϵ�����u��;d�}��8R�"�/���=?^�� �Y �y�7�t�:�˧��ҍ׍iQBr"��kr^*��C�^w9�U�"��l,#� ��{�Nx��f���n;���V
:G?�ky�~m�h۫|�4r]�@Tջ�"T�r3䲚7�����Y+c�u� 8c;��Hu[	1�8�"�v�V��ޭ<�\P���2�ƒ��<���v&�8",�5�b���]r��*����F
9����b,�6.X���B�"`��:w�Ds�,�ch�y=�9��f��N,\+�'[�T�N<�����I�):��Nr�sk�D�����kn�侊�9��M��&��h��E�	�Z��.Ru��]�ɔt9���k��}����Q1ۗ0@�0������w;b�kGm�|�ռql֐,��V��y�i"�y��O�R���[�"5��~�����}���
"�
)"jb*b�b��*��(����"h���d�(f���h��"��"&��)�*���h�)*��"h(���a��fj��&����j!��`����j*���������������
**��
e�(���j�Jj��"�
j���� ���b������"����&��
*jb��*�����I�����*Hh�(�J(�����B�B�b
h�����"�����*��d��"��*"J���!����H���Ji(�)�b�* ��	�h)�"������b����*H�����������
J�&��0r��`����h��&�
b*����j "�'7ٮ�v~=����z|\��uNE�.��E�j�%�Y��}�����c���z��X�v����O�f�?3���/E�W� >�gkn�wvw�IcW�N�-��w(3;�Q%IpQRf:T�{@h���5ڪ���S}0%%���3U2���ua^�¯{�<�xj0f�@k�tv�U*��v�,�,�N��M��W{g���}5U���R���<ݦC<<#i(����A��ץ�Oy�����jc� R�x���r��W{�L��F��e��`p�.��3���n��$x3T�G��TE?s�*��9�E9��,<*u�5٪��n���ʼ��M�ǹ����ub폭�`��K�2���2��&U�0�x8^�GpW�Ԣ���*����ϷC�zO�G�3ў��ӵi�x����u(/��xÍ|�.\�\O��q�nRU����'�K��t�=x=S��:f}w�C�]��(���. u��9Ol�je6jn��^��m_��m�A�.���c�*��x�A��	[.��}6ȇ��}�Ws�(��G�=�d�9g�u����_D.�Q�^D�=@����-��5�ϷdQv{����镛��w�dr�*��s�M�>��z����A��Y=8��{�ቱ�S$����2���usP����S�6�z�D�j�ׯ,-��������ޥaԵ�G�Rts7��W�4Y��ݪCM.��iz���Y���u��1ò<ش�%�_��\+5����
�������_]�B�:*�/L@X������?e����h����;�^�S�Z)|�~�yH�+��*�,� 6/
�Z�Ţ]>}8����WR|�>�qڊtA�	~L�ʖ<��Iqr�elB�#W�m�;o��f:\�vD��Wq7B����d�>A���ɔ��)V�	�� ����t6�vv��Qa��=�X�j g��/�7/�Y4���B�U�pewDI_����S��*�i�%�b狅n��z���*�%O;Ȇ�Fa0����1%k2�3�!c<����nmd��o��;H+� F��g��
S�U2������˥�u���2z���.!���Jj��O�.�ap�	�kR��<#*|�3��Rյ�1Z�|�10n�{���D�L��GK�U�;��Ϲi"R;���-U�q�<�q2ro��pp૎�Er�E�G�-|�{Ӓ�0�-�2�����3�¥��z����00�����m_>��X�w<��K�u�U���*Ŋ��:�;;�ͽu�P���]��*�_�
-7o3�0�*#Kg��î�g�b�#{5�'���6q;!�=f��x^<�"����Po��m��|��g
o�G�(Dwqʰ�ǇR�˩N��e>o�15s�z~�懲�Ƴ����EN��om����l�\�Uc@_`��z� �bg���d8�%�X���)��km?{�̮4�c5^��aT+E_g��tM��
��$J��^�//	�Ȏ���r[_D�!2��S�ޙ�)��,�|.�B��kg����AQ{�	�W��3[gͿI�\�ڋ&o��Ӱ���U��G�������#�H����N�h�{>�C7e��M��������`g��G���Q-��[;�enr�<롿V��B��o�w��ȁInɜ�g+�� #j�#+|�#�酞�ǫ>��Ǆ���~>���+a��ܣ��=�"W���
=u �dU�Y��]�N(X?^3cpm��qL�Z���"��/%e+zU���9`e����#�(+o�k�A��es���[Ȏ%�^�~���"�f�r�!����>�ۏ|��6V��w�6��˂�L����$�ֱ|��	����xX��/S��<�^�����)���n�j\<�i�$��0W�݊��`
�(��{N5d:Vz�?$�c��ǵ��oRn�� }��\*3f�8u�����H����4�^3�񳛵��gX���c8m]l�V��r�uv�B�l��Z�`�����������zA�m�+vy�}����|k��R�� ��·�}�^�ڸ��U}Pz��vAϳ<?������~�{��1PnU�': 5QB�]i�e�%��F��QN��f�q��(�Z]��;m�KNt΋��#��ت�c'w��nέNc��T��x'�u��&Tλ�)�:��80"���&(e�b{�����y���v�Y[�F�S���V���"aҙ��HE퉣����Ern�{ۯ:�����FN��{�-鈔U"nYB��l{����Z���Ymz��3��/"����PL�3f�s�G׵����"�P>7�6�?�*�8#Xy�����D�1���b�7j�O{N�y;ҕxM({{˃ʼDpTt\6jҰy%ו'H��-׻݃��n�Q�5ޭ�!9ơ�#�^�ܥ��zG:"=$4
��YB��ܦuMOP�%��/�ꐡwbh5�~���md1�l��&xԭ�z,�����2S�KZ��MB�D����!�����Ϯ�V4���j"�^̽em >�^�Z�0��9V��9���T7�D���c�୼,���*�#Ce]L�e�WU�C�WV�A�GS���ʜh΢��Ht�;l��~�ֽ��`E�k¾����c�Tã��Eq���h3rj۫�����7��;�e4�Uo|�[�3���3����Pc�L�N�hh�`��}ulEYl��lW�q�!�[Ƥ�n=�Jg�t��Um`�ڗU<�B�Q��G�мKG|v%�P��6p���\�"�����e�];*7R�+������;��`W�X����5^^�]�Jᜃ���2��sR���޷��̩�(�
��|#։��+s�s*R�e�Z/��I�冏s�8�#�|�h�3��C�Z�n�pz� mwgם�*�v\�l�M({»gw��́��K�j�ܳ�-����-�ǽ�L�{����� ��Te+������W�˛Q�n*k�œ��L�%��.�=�Zi,R6�;V2%�ݺi!�wU�k�;�7��]�	K����x�૽�fW�Z.x~Ƀk�w�qu�p��fr��(Z���?f�Nz�֧�����;U���`��1�� �k׊_#~ͯ<��z�#;�б�����1����E�
�y�2w��zx*��U���c8����i�(=��zu^"�wS��6�{��|Q�}w/z�U���{��WS�ۥ���K��x��U��봄~�p̯];���0;�g�WY6q�w�,fA���u9 :G91{\,�/q� ަ���;R��5�xm�C3{�.K�q�����z��<Yv�X���x� [�T�Ӡ��xÍ|�V�:�~>�8��*��	�CPG�Ö��R�*�
�]h����>1%�ҟ�b���p3��q��*�nXz&fg����{��s
�L��ֿ���d�g�ґZ:S�c�{�H9ba�i4�zy�n���m�\�r#'՛��d5̠�Ъ!u���ʿ�d�\1]�r=g����G�w���@L��/��W��2�_�<�`�.�+�E�N�Ы�)п���8JZ��W^Wv�y�kT�����ɾ�W)6%��'4��s���tL9U+>���z#�*!���5os��� 	�6*5u̪��UL�>g�ʎek�T��i�K��C�(���w��Yԯz�kS7�]b�"��K�%PJ�Iє�����S�X$0�*�*�Σ�j���d\�҄�7J�^Y&�Y��a���#҇�>�B�O`�J��w@���;�r�Q[��|݁[A9c�|�*y]�C
��ª��-Y�Ղl�b//`�֨z�tg�-Ն�SWWZ���#[ݏ6�3�`�Ʒ�>�
�g,�rc;X��9���)8��ʒB�f���u��� �S,<=[Z��ꕷ]n&(]�:�>0Z��h�X���e�/�4/;h�7��B9o^n������YT|��W��{�Sσ����Vɀ�d���y�u�U�͚��KΥ�!I=|�)-��=��s�-��ʹ}vL�
�j�q|�{>8r�r�+Z���0Wt�^>�6Ns ^̗�3�(�5�h�.�-U��3���OM�c�~�8pj���j�i���).�#��%B'e���|R}L����AHs��v6��W�_;��Ȏ�S5�ړϛ^�g����6*ª�e� ���s�
��!�	UX��G�ע�:���\��a�S���������
���1]���U_Bh�p�G"�����yv־&}�__��ʞf��cj1{�>�p*���|.��I�U����1fǊW*�2{2�ghm��(Hx��-����DSʴR�Wq|�#dH������_��my�wo,����6C!��`�s|���Jτ\��0������E�=��=۫��'�*y��1��5�5��&�թ���,:��I�䎩r����Aov&���ݽ�,���Rsl�з��Ӗu��$���og%y�c�
�溮����k!y�A5��2Q�G�M��z��bv�/EZ*�q�i�s�"��h�����s�Rƌ%�Om�k�;̮wF�*�Hݙb�.�=v.��s*ե��Kc����8"�.�纝aƳ׵�^};%]�4>ʿiU��]6羉A��������ޏ�J\�#����4��ߦU�_S�E�s�*���%/r�/r��?q�?����=[��W���]�Rc�`���\�e]ET�j��/���Wpudc�w;��&�W��C��xi�dr��`E.T���F�PV�X8�Xx4\^�聯a[p�۬Ԍ�+|�{�-)��m}�(�����[�s�E�Oݘ��������5~֫�୏i�e��ދ!||�uk�����)QY�u/�Dz����q䥙N��g{�6�n�c�1�*M��߮.�-�����J����� �۰/��s���nt穁��xK\�ߙ[�5M,F�|~�ӯ���y�t&�Go�E�Y�fϳg�S�f����HVgͦ��:.�Է�|&Y��	�&���®��]v�s{إ��Z�BP�\'7-���Gu�5�5^�����"��+ċF�M����2���D��S�>a]�X�|W�(p|��K��ڝ�O��m�����y�p�o��h�P��z�vO0�orS�����w^���5�3�t��yDվ[p�bw�5�}Q�Fr����ԣ��i��	q�Jq��t�oc��E�1:�'V�t_m<���R��G�c	[�xq:���ĪwxeM�����z,\�7s�����^I>�u/�U���	�;��j"
sn���kӅҐ����������XU/�3y���x�@����%^i!X��eP�~1�l���⯦�t�nd�������{��)TB�SH��z��,E�ݽ��P�?�y����Ȯ����/{V�<��pAȰ?SHп��0*���˫b,�L������y@�yr>�ZM��=��B�k�ho�
�j�B��B�-��ܬ�b�U��]��/ͱ��;<2lE�ʎ*ג��܇k2����ҜWT0
����5ӺT���n��|�,���w��RT��討��p]�� �8bV�)'Ɛ�ǋ7�ɣ�Z�}�h�XD!�2��|����(:��~}[�(��K���L�@R���j�M��[���=�	�Pe?Y�@�>"��0�fE���?I��VK2KuH�!7���eq����h�y�3m� %ql<3^㰔��Է��5�e.OA��9g�o���qt�$�nOVnD�:�F��ʔ�8�i�+/�+��=���ő�B��:�@�/i�:����mګY���2ƅ��B֜mK�H�GK��]$�hj�U���%S9�߸�#��@^i��b���<��Z�<A�Y�s��w�k�!c�/��y� R�C��w�bE6����s�N��`������N����6ǩ���f�=��gb�~��TBq�Q
X���v�Hk�[�M�m���Ъz�9�$[�����6���ނ�C�?_T�}苬��zr�����������nG)��xf	^�h<��F�R���C�[�<aw��Pq���N�W��]�^�=��f�cU�����h��p.8��LQu�p�@l{f���u�H�ʝ.h�������(^�Sk2��<LL��r�=��! �W��H+IKN���jů�Fc�]�s�`�����`W�U��V8N�<}��$�;���\���ɘ��g�5o�w�($'`��Y�ƓREK=3��B�4S���{)��!kW�b=*ōx:u�<���r�b^��Ni�(��D�E`A>����7	��l*�o}�"��i;ӳ,��΃M,]���%|*���F���[�>���/���
�%z�X��.�7���+nL�/,��f+e�0b*��t�x�j��]�;<:m� ��&���c��;YG\%���.�ĞpO��t�P�f�Ũ���Y���ZŌ�v�݉�Bd2RO]Ie���ts�J�i�R����Hd:�|B�����8���-G�Lk�B~�of��+�w��joX����C)�Ա@���o.N��_-<������� _>LR�?�d)Wҭ�32>��wcF?n7��YE�����E����'�:t2<�풰sˤ �H���N���+d�x��:�igf-�ú���9��ġ��9f=�JMQ�p��X�>��a��37V<r�������J�;�Q�8`I�.����)��A�˲�B2��3��9�CU�Ι(���>�X)w[]�,m�G�`|Q����1��X��o6�]�4���Z���i��X����_V�����eDx�9խpKXv������,�%�l��rK�NԲ�Mv�ǉQ�~�v*��e@��RƇ���y{S/�V�&&�&b�cN@+:���݄���[��J�kL�&�۫[$�wm�@�� �T�*�)��G�xⱹ=v~�ʺ����p��=s��w���֖.�PQL�է������3�Ʉ�8:;YD	��m[;�[k^�G-5[�fB�Ԫ�[F�b�����4�6��l�K�1�W�5�����;���O�Ý�#�ޔWD��]�wOt�+�ड़�1���E���P�^ZU;IG(�2����>�{����R��G�b�_M�*��QR�`�0�G�7�Wj��S��<*�;�G��;����GS6��:�Č/vTI���଻���"K��J�.\s1�>��nN���f�B��Vw�ȷwV8����	��K{��C	��q)�[�P�G�n<�w2��}�H��tɊ%z3ka�6��E�Ֆ�]��c�=�}��-XT���h�|h�
�z�M�7<�����M���X�]�SX�����2��d�N�͆������w��s+y���"ۓ�*>o3K�0����8R����Eحou/P�iotՐj�m�YXrp&�Ì��������R��+��Վ�h�H��|e\8��^]ڭ����)��Tq�2����h�����I��+�*0�'-Ϣ�g����^�����f�]ӏ�e��T:5��J1Y�w�Q�)��uh�X�,�K\^.xbP�,�tK^F�b�wXK|>.i�&���:��:�}�/vW-�&v�wr'ƞ�����6tpůGQ���mD��v%]����V#����+,\.�/�x.\���X�9y��a�wk�j�3���ʜh.�/��odʗ��"9¹*(��Zպ[	�v��m6��{\5P1�F��+* 8��|> ���U-DER�ATUUM#EC34Ԕ�PQK�P1$IIEPU5I2�T�2D4�E�4R�SESJT�+Q��1MP�
QME$�-P�U%SAAMD�Dy&QU UQ�L@PFfRPD��4�P%%STQDKBP4D�P�PS�D%PC�J�5KQCUEDAM$KMUQSACTP1����D�T�4Q��5IACT�AL�T��LHQE�T4PMCCMS_UTPWS�����u�D���˃a��3��YM�I��֝bh�	I �<ZZ�嘭U��ۼ�x�q�ys�'O{,���~dr�� ��@���p�r ��:xgw�����c7�K���m�/��9��$�յ2R�u�"��x�~�g´Z��v�����Qm��ez��ϛ�
{ym`��g�U8����d�����r�U���#!~�hC��*�x���n�6�N��{s���y� �c~qYA����7]6��Gк^Z/-�uV�qΈ�K~��'c�ֿ@;� ��X���K`�疪ew����u2h�$"���}~�v��b�}0��[c'�f�>h;
�k�+Չ�}F|�?Oo�W�u��o�ӑ�O�-aj��ޤ���q?����E��,Us��)V�?x�X�7ʆΦ6���pmme@�P����v���ܦO��\����(��� ?^���-�Bt�Z�����η���J��v����U����K�����/x��������e��R�_�b���������y	�T�������U�]B��Y�3.�EYn���RN���[�����R����A��sBxJ=Y���A�)��w+j�,�E����,�	h��74NWʦ{XB��l�(-�u�ޡ����V�[֏W$���e��g�Ǜ���WQ�S� �%E��e����=Nm�ԩ�����k����H�u_2rj���vT�7&�Q��14�8i�
�:��/�p���N�G�N�4�RZ8*����o�aO*�Q������T�#��"8�վY}����q����'��_��M�.���چo�z��$�U+\��0���a�>ayX�|r]��7շ�Q=l V�>!��C������Q����=X+c��Ne<���˰��sL5ݰs�P7䩣>��&�W;0�WlFr��o�Pն6;��VqX3�Cި���,�����ɯ�hW�oqh����>�WM<D]s�%�ߒ���Q����!kwo��dc;�h�t6s�@�P��x�ch*r�S*�*x�5z��E���{=@]�Y쓸v�lk<2}ڽƠ����Ϸl�\<�� g�|F|`�[��eW�������-m�muj�S�����t̻p�~��l���Q*�� !|���*ޓ���n*��|�J�MWr�"�3��Vn�E袅����(JG:���|��f��Iϵ�TW�s�~��{.�ws4� ���Yb���85��m#B�=�\b�m]Ԛ�=v�Z�c�������氛%6؝����ܷ5��W[�T6�i����;W�2P7؏C(�`���F� x/X[u�i�f�i������65೚c�tނYmڿ|��u�[H3�R�R�x�hR�}ꂐ�yB�w�2����~nC}�ݺ��$\J�_����Y-�L���J����0zyu��������M�c1��W�]�|�A���wCyx/��{�"+��d��
cEY旱mn�v��OioGǋ���)}X̄�׺��*B;����M�5�~Dx*tn-��cːpl�m��9b�v7�c�}�MA��-�s���V����^�����z8%����a��sk��ѐ��0/	�v�VUʺ�[|!+��2m�9�b3T}e/^W�`Δ��T�*�J���8��`�����y��f%����pM�X���e�㥾򝧽���q̐*b��[�ioY�<9tX�AUu�v�C��oE):u��w�n�s*�c�������٠��0#��ʺ�&�Ī`dڑ>��x 
��J��vf�?M�@�I�]H�OV fe`�:�X�C�h^$/_���m�-��ݡcCt�׽��4�nŵ�](���뵯ֳw5&�Z�\W\}/��_{�V�=G@򻱧��6���oڎ�jm8��l͹����ñHx^'A�G6p����j�!�%�ؖ�3M�ŻF��	�V�>��Y-.h/;����y��!�{�G5ƅ沑��p5Y�M��YU��/2��}�ʘ���yNv(-�⫭�N��9C�S��<	�*�Wo)�u�rtTD�3]>�&3�\K(�ć����ϧ�����ą�Ya��ʤt_��˃�su��3�*$��%�DF�Ƽ���ͮ�y���n��ʑ�}1(2������X�����JOG��=*��F����dk�҆�_M⻕Vv���b�Ie�}��tϚ�^��uX����P��c����ۙ�&�?m@^ឤ(�����Uy� R��\;�sn���#�!x�bc�\>��g�#�>��*{���\xV�cW�A+˗���C�<��2�.��*;�ל�x[� ��.\���֓x���RX�Vn:�Y{Ai�A�uD��.��ed�J�*7����є��ż0���Uj�h�s��^]���]]V�tV��r��ª��S���(�I�7ڸ>}9�h�g�3���LW�����ayWz$��ݗ ���wMy��S�����Ѣ�jWfGȭ��C�Z�����L�7e���0Xw�Gs����2֫����i��/0����o{�Xx;u������iQ�zS|p��Z٧6p/�t"��gBV��"`΢�����[`���{��CI�W��s�}np������ϼz�$Lw��^�ƹ}wCM�O����ߩD���=�ˡ�6,i���d��]�}6Ȋ��y��������UQ�TlW���� 6i{��\s�9w��G[�xd�v����/w��%:�2�_� ԅQBXy���o�n��	�z��.����R��/.�����i����/T�Z��搹.w��1�ո�m����<�~Y��<���� Z;Q���Vl*�Q�:�������c̆+{;|��m˙��:�ӳ���>��3�pD	��%}v�u�B�ۭ��������B5W��P#~p�{r=;�k֐�>�t�����xM1)��ll�]���,���gՐ�Ú=���{A��\�R���pgwY&	>�'C)�����ϊ��S��"K���`��GZ5vg�j�5z�;�0]O����o��S}�\@jq0x>�`yS�U���:'������|76h�YS��"�.#1��;�x�ιN�낈�8���p=': )}T<.���&m����[R��=I˓")�&ks1>�ut���yO���R�9���(��ѓt�t�*�F��u}u;7X�j�b������мl���lC|�&j�y�K]}�"�=4'4\��oQU�!�xh�*��˝�6t��yy�)�a�)�h�ӂ�o�r�!,���J��/�����=�2�����d�鞫W�`�/dO������O��.W��]^2�1}w��w��P���
�n������x<��Ye�'����r5�]�u�}��?�=�t�)5t�+�.X�����w�-���^�&|���a�%_\�j�PqM>�i���!���m��g<b=�jϷ���^������#�����j��s�����m����2�쬵ƴ;��?Ul������&Y�n#����T����㤽��\���Ϋ������}�_O,�1з��J�w�q<{<�y2��%�h�\�Q*y\�2s��a������@����_lu��:z3�ݭohv2V�"а.���E
��Q�4��~:]�/N���K���ŀvv��0k�\���IJ��]��,kVh_;0�WlFM+�x�x��~Q��xf.Aݴ�=y-[�V���l��ɗ��x�";ܼE_��If����c�Y�'��^�a[�X�|�;�c؂u����p������b�ZY�W4�V�Ӵoqn��k���

�l���M�k��cX0T���Z���c[Q��g[9WWJ�Ye�Ê~uh-=����u�j\ɛd�pqy����^��`�������ys��ݚ#%{P�b3-\���"=C&\�U�T�j���O���f�zhNo(�����a�^q�;�y��n�"B�����0J~]Е��������js�0�@*S�{⬸ubRO}��u��Y��t�%}�
�r��&�?^>�w�'��+lJ(X��#Sն�l��q\��Okw��zX^�k��8S����;�S��=����9M�ۚ�F���f�?z�-�۬��&T����Pݧ�t�c3F�Qf��7{��w�q��x� �j֬�ϩ�x+������~(�^͑�3pK]����P�nx�2%.P8G�\�&UH��g�����v��Rޘ���O�_Y���w��Q]���X�?%�C=j���)�X̄�׺���S�;Ù'zv�
k��*W蝧B�
|�����.��a�|�*;tʺt(�J��˽M���A�U��~s��̰�.J���� ��]^.��+���ch/��]r��!>dC�"
���%��3�7�C�p��օ�>$�Q��
�ۜ�z��	��t,��^s��r�mպ����K&��뫥�1VmX`^�.b�+p�<�L5p���j��W:j��o(���y�ν܍�W��#�s�}(iC���[b�^�9T��m!�P��$�N^���w���H���/�q<4JP-�#�P���Z=)�+_��u��>@tZ���Ll2k�y쁏�P��̜1J!u��t��C�	���if�b�����+]�mbp!���Y�og�u`��TTY���T���@�.�L�8��g>0��V��{�8�N���n��K����%��#z����pp�I��z�'��M�+j+�H	.��gM;�5�L��b�|9g'f�f������y�;������������7�mN��ސ+��F�'� (�_Y�ybT����a���Q>��'�`��^�kr�o_�Ip�ޝ�?<�lo��Z5����YC�l-�S��й����<d����w	觲[�����z�}@��&)s��V8�ЪbPg��|fUu�X,0�)���I�|F�dp���0Ιn]s�	:"J�d�ET��U%�:O�Xҫc~�>��YG�K	�=oS�b�cΏ���б3�?7;VB<xxMq v�� R��}���w�T��>=�}m�j����r�nH�_!�sV�:`���ÌK�gc,��r��Vm���H�Nnp��Ik�����=ǤT���V����T���ԇ-�i�H��Z�bf������S�g/���q�9ۍ�Z�������nq�ˏۑf�ϲR�|F��AOL�oZ�o�
��xFW��n�Gz:�	�]�;_��+˽$t�}�c�V�&}w�s.*ҫ1W�t3�5���^���X+��[7�\i�"�;Ħc-����;*!��Y�]W���z�&%J5��.�޲�9M|���ϡ#}�����Z�ە%���8���:�V�0��,�8���J~`*� H��OI��=p�����3�m�T3�Jrߎ�aV���5wCM�O��ϖ�8����`�<�ej�����ܦ�A=����DGDvjxɹ԰	cx��i���Z,�%��ʙ,Q�ܭ����������_�T9s=(��7��{��@N�U��_�&�*��w���mox�E�d�����z;�R��.��=�uu�b�Xʦ��}/T�Z��摥�2d^��,]ow�T��h�;f�=c%n  T�X� `����o��8�3'��K�dv<6˾���{��Z�޾ë�c�0g�*��3�Y*��?1���A�� �[�n�r�)��8�f��~�6�5*�pC}Q�y�ϫ]���P�Ҙt���B�*B$z�ki����V-��F��X�E:��[�%����!h�M0zL�B���Y1�}��J�}Ϛ�Q�'�U�]��'U������MU�����I�;��E���ː���JK>,.�J`�SĒ�Y��a���R���Å��	Y�c�8�;a�L�v8�;�$���):NX��|U<J�e�Xޣ<o!]J�owaW�������}�\J�XJ�e�?�����4t�U�8�IE�6�XUO-T�O�ѭ�x�>����%t���'�_/C�Ұ���?wٷ�1�<V�(��� A��Q�W�9}�=� bo��{�i��k]��1҄,3��C������
{�~��L�S۸���t���Ӟ�#�m�:�mxiu+ٖY��e .��*LvjPR;��Y���e\�=|�[Y�-z[���,2^F��;�=\8`�0ݽ�ՏC>\�S�R�-�(g�`/6t\�dZ=��Z�����qe:r��wQ�4�(�6����s�f��S[9�Ό�^��}��>մ@�ĉV��'*j����s7&���2��Κ�-� �N������o'��X� �~JP��2�OE�7Ӱ���h�7zΎڹ���t7�tj{��<;i�)ui��6P��7�d��6c8)ހ��-`�Ǌ��%_VM��G
+0AP4u�mN�[�zuIݘ��n���nDp	�7QË���B��oU�����ݠ��ߋTn�w���	��=�,!o�79��nQ=K`v��NfA29�ٱ��j�Y&wV���,>F`�e�������d��kO:�c	��O��+�5��B��{�ԡ�B�xq�O�d���%�ڼ�P�+.�X�>~k�q_֓��b��a%�x�Ak���a˼�:���N�r[Fب>7��V�som��Jj�ݲi��|��(�YTS�Y9R;S�Mb��ȸ<An�\Uq:3m��Un�՞U/i{���S@h�~K�1�˺�_�Q���ڼ�hZ�' ��a�r��5��cz�D���fJ�f�t��Y�uvw��ș5x�8�R"LU3��Slcss����B�s�z��>5p��v�*��Y�xA4�N�Kh*aSg���k�ص	!]{yzu0����M���k�a��:�k�u#��7m����Z�ug4伻�B �[�Xcb�b�΢Q�}[ں�D���v����0�]s�FB�E���-��ȨAP����:�ܸv-ݭ��O/���^�Ŕ�Q#F��j�P� �X{�J�����Yzͼ��_��D�z�]�r�N�ڰ�6	�UKV�?\h^��ia�uy,�Q@�>�K(gQ�*Cfhz�k���Q���}���^�W��bw��F���,��eh��1��=��-L��}/����ۉ�n�pMwu�9v��F���S9�*�K�^Ӕ���7j��SPPQ�~cQ����u�X�:hᶯC�a�Q��i��@]�MR9ڷ�yy�(!�Ov���D-\|6�Z;.<��Y1>f��u��.�Y'��.=��KxZ��gC�5�����]��YiȻ�$���N*"��Z��%!wm�lm�ruض79�^g�Πb���C���IYt��y(�T��4��&�17�%�:}� �:]t�m<8_i�o�WcS�5��ݷ�']G�Vִz��\��c:�]Y*�԰�V�kP�Y�5�]ænD��e����Z��B�/��=��ٱ���Օz�o��pc���H�*w�N������LK��j4���v��H���Dk�q����2����ƺ8$q�_K�\}�v4;[�;Z6�j���2d�Y�1��3�U���/��O/��?V\�I��8V���Rp���K�յxp��c[�~o�8�d��a=P��!.��ʉ��՜͚r	����vd���~��>���fWS���ىH�u���;M�����;*n�BY}�3���!
�]f�ݒ*�&�_�6�T(�l�g^J��VSn'�]s5����������9�g��i*�u9�M�tՒeuҮ0c-�nW\=�}�ޡ���PU4�fP,�!KM,DEДIKMURT�I-"QE�IAUJUD�D�Ӑd��E5E)IH�M%R�4�U0���QQPE$U%#AM)TP�ҔU MU+E-TM)T�%$ITIJPPDPRMU��P��Ҵ�TT@P4MQII��QBU%$K�5@SQIKAET��H�R�PP�BD�-R҅4IB�TE04�UA@SJ��R%SE���MIO}@U}@_|y)�W��Q�:9�m��[j�$8�G�D��.�������nf��aɕ!Y�_̋�½�t���7����V�S���t��������E���Ċ�R�Wg'����.����V���\����=Y���Ǥ�����e�Ac��G�9��< +���Mr�����^�uʓW~�y���yd�~{�1-�}W(?BG���T՚��%]�ʫ��]-⩎�ٵ�xFV���,�
�0<έ~_\9�~������9.���s¬s�*��b��9J�]-��O{̽�N/�8z}ڨ�~�68N.ձ��Rc�F�Pɗ)�uS�I���]�y�ҭl���w�ğGq��:��=q����A��^V�"&UK�ʆ� g�pY�������
Nz���K�<�Fé���h<�}g��!�HG�<Ր��z+;��z��Cc!AО�ʺ=���4J�{��/��<��&k@h�D57lE��nu�R9ש/���E�m0�V�C�qg��f�7wC-բ����>�@0<�� ���Z��O��2��ҙ>�k1�#2��}�>�Dtk���Ru����t\LeB��!t��L~��#](�-�K��y�%�6D�de��w����]Vq�5�[���v�4�n�D�=�F�5V�)�EmԆ���V��O�P�m�sG���8k�����o�ɇ'h�rR;�[5�I��O}���^'w)��.�%�@<��d|�^��V�H���{�ϋ��(6V����HG�r�]�O���B:.�Է�	��e�&�<���3jOf�wt�]�^��Hb\ʪΫBP��.�����`�F���#��gd��p���ou1��?R�-C�Y�i|z뉩B�P�P��l3����ڜ`f]`˺өnb��Aq������s�yA
�8ή��Y��J�]r���O���p�^���lU��~��I��f����N�����X:,�<E�Ė�"En��
ۃ�c�=�$����J<	����|G��eN
�����H�G��J����S���{�������:ߛ��ǰ�ܾ~��0p��gO.g�}B� T�D��O(g��<��^~���y������.߭��g-mš�1�H�OV f3�+�j�iйJiĳ�it�#�
1��H�{j���Y�Y�*lE�ʎ*��y�9��������jdЃs.�^p��Mb���YU++*��xfC��Ƿ��f��H�Q
K�iӓ:h�^�)��^�O@��]���n�^h��W��^�Kܐ�P�:y��#���*Yt��ʕcsos�G���첞���V���;iu1$�ww:��d�f���T���/47V5u��q�}$���}OT�B��3��ٜ�o���Z�MI5О���C�^m�f���Ą"��G���]�c~ͼ�U&߁�O�B��u��{�k8�'"�
����A���@h_LJ��ό���]Pa]y��VLXX�G(;����cÇ��;�$���TUH�А�6No����߄��>�j�у�WF��'$�v��c��@Jƽ+9^?S���� W��
_I��>���s�ʢB���;oU�:M���+����j�/��W�d>��U����c����Y���;\��r=͝����A�}��?TRߪ&rݚn�n�������������ka��؝mL:;���k.O�H�ǵ&�������دJQxxez°��&:%��R^K��T�`U�X8xW%S_O_=���&?a�a��������{�b�+��P/�l���l�xF�L��������5e���>���3I�	��'���
�������i�|L�*��k5�c�E���=y;�JM �p������T�"/��y����N�r��V��2�xdv�oB_�ӺYGOYW1� ��]ZL��S�	2�\�r&ݮ�ͮ5��3XOG�,�n�R�<�dU�����ok��M�&f*�T|1Yn7{$x>����|o3thDzЛXn�s��]�-��2,����.Z}d�Ѻ�H츮!�K��q�uKk��9��9��c��}@�Ҭ���,cQM>�^�+Ӭ�ef�_�*���8A~�Eŗm�}�݃�9Z��W�(]ᆍsW�XSMM>��{-W
Rs��;��5�=)^:�`�����J&���CV2@B�>F��+7���3�g�)��a��ΧR��IJ�g��dR�[��<�G�EQbT�dt%��+�����(�7>�����g�(��u��ʋ&S�)V��K(�g�*�rz�2�=		��]�#g;��͙ҵ����H�82��$���B���T�E:���Z�v��Z ���+�zp/�ɺ�ݺɀ{ê��Z̾���G+�"��,���Al ��XV��̬�W&�8����%F�|�#�0-�,��{ګ�-�a���z��@�8�q����Q��gN�z{'����X�mK1Z�~ ��u�wԴ�ROv��9�_k�~&^�m���kK�'��b�@�}��W�ٔ��.�{2�1[�D�a.yxu�~�G�&�Z5d�|;�XF<p�j���<]��7�p�'jS	g�o�Ԛ8<�8AhJ�k�����n�J1��i�uot��oM�(;sje%f����/0d��^b���{Wɾ�h��b�=+Sb�Ⱥ�L=�c��b�L����\�n�p�_`���p��w)��;���/sFٱV�-q6<�.X�5�b~O��mo�k/t	��v� u{lL�Wg��ќ�t<�CJ��P���; ֏[�O��u����y�-�װ�W��WКY��%�(x��&��w���r�\��r����Y��y���0�Pກ
vZ��ּJP�c,��=y5�,:����Mmת�j���/�W_Fu��>���Q�r�'�4H�e(�v}��'(o�}U� ��r]���N�֌��w�z��5}�v��DpU�/��ExѮQ�4�r��5�J��zyjj@�$=W�2�˞{���
��Gi�[
��B�ل��u��:r�����{1��=�A�Xɶ&��=�O����]��8&\D!p�b�M�F��6�k�6����;za��fWlt�ED5�@l8����7�0Dz�L�)Tʺ��u�`O�y���FJ��R��/�_3�����4ǟXy{�dHPc�6�@{�WK�<M�ΙІ��S"9Y���98���
��Y�mZ���iT#�z�)��[�2�`o#Q�Hp�X�s_��$9��i���ӫOm	�;4�L��d���[�i�R;�Պ��!�Ձ�cN��I��.IYy���Y��*�;�9E�v_t]V���e�p�����U��U܆��VB��Y�0{��fO]=�2�	�4{�ڑ��<��7jޓ��U,0���Mm���n���n�$�S�����MԚ���W8��{�I�$�gE����*���N䡔2�f�#�)o�F� z���N�ܼ��9ԡ���)�h>��c:.%�:N�O��7��~��e��X��^�7�γLò��6kc��ҙ��!��O�D�{>�Q�N���-�Bf��ʼ�y���˪�쏳ݩ7e0���VZ��P�T=��r�-����?~�G֮{W�#OV�~��4w��X�K�#�v�P��k�u�}t�Q�"�3�[�U�b*�y;ҩ�Q����M.�F�k���nޏJQ��`>�K��Uh��k}�[�2!�{/�[Vna{͖�\��F
��b}FE�׾�.��3�^�;e����.��v+�ȣ���4nT|q��`F3���l��v��T��pT�K��#��*��W��VZ�uz��P�3k2��e�Y�i�MFYq��65S�	S��-:J�P�]#Xݕ�$BCj�3K�IK�VPtrl��COhX��=Aux-k���8�P�(�"ý�o|-ְ��͢�}���:%�+�t��ٽ�f9	�u���V�13fm�7R�;Oz��	ú_IG��U�W4�cJ��g��9��C��,
+�9��1P�R�$hozߦz�(���=�5�L�)R��.'��°J���2f3���L�	Kh��9���w��.�4(T�.GC��ձ�-��)G<x�:x>�-'[�g����b�Q���W��ZA�uGٕ��y��`1�������wOK��>�u�p����L�|k���Oz��Z��)<�q����u��G��U�6nco�Dm�r�]�F=�4̵�����2�wvQ%T�&c���s��A��g�gX��c��K���|�ߩ]��Cl�9�͐J�5-���)�������_p��Z�:���]3��Q��u���=>�6����L� ��'��Zd:<<&��;��I��=�1��e�t���N�躹)��Ѓ�X��{j^��6�
zd>��W�r�\(xeyǄ-�y|���6g?:\���Rc�;�9n�7hB}
2�Ob�+�]��[��q1%�2�-���=��X���4�*�T�ʔ���Κ֬�-y~q�Ӧ�$�2�`�^Z�x�>O�+�,��Ŕ���mEˠ����� �v�-�4Y`k��kSI}[[)һ�1���u7L�:7���m�.f3$u��#�EӼ-u)�+����c����_���|~Q䡨d�J���R����w��n�2Tf��«Fx-oA�[�ۇ'��<g��nfA����������ʤ��u��=��Ė�+�����ٱ��S���a�F-�՛`H=��N��z{j0�Y�	�j�'��LNM�B�]C#�����U�}~�R��=y�{�@�,E�6�SS�����pN���u�w�'�$���x?{�
�	d� 3j��J�,cQM>�x�*��k!t��`��t�#z_�V{Fy�������h�8.mM�W���@Ff]]s��,m4��ꗪ{-W
X�Y�J�.�b���l�������{��3ꘀ�L� ���NVoM��\�摯�~�zucǫF��ɑ��ǙBK��E)T�2��*�[	�r�m�}C��m<��_�7��S&�p��K#�z�qCGfE�)��FIe�.�����L�M���~6_ ��yw�lmL~�{�*�]��i��83�"JT):%�[A}NX�T�*om��hJ��x�M�����YH����Y��Bɨ�wj��|��͒�`�fa��P���2 ,�Z��'�@����i��-���lO�!��_�c`R���r[N�.R��Y����%{)��c�ɽ\s-]u�9H��M�2��7Z�_��:>l�焘=�Q�.�/ī�eȸ`��s%�f��� )� ��y��m���*�&�oHߩ���9��TZ�J��XX�Љ��ex�r��Z�5$"w��=Ǔ����p�U��s��,��K6��[�n�(B�<��խ^��ޒ���"�S�ǫ����7L.���4�ʛ��v�\8*���gLWz�W}L�|��.<��=�ڮ	�y*}�r���<~�		 �S����� ty츾
�^Rnq�1_����թ�tW kSژ�-Q�uS�U{Ɛ���{lL�S�PqM>�p�*z*�pg���p���������3�8���UYr��`�	td%�5AK��eOU3rm���➌w��[u�5gRp_�g�?�^V���F�f|���|1�K�`�ꝄE<�Dø-��Ϳ=q:�N�D{�ם�׍��$Gt\�����ܻ��<d��&���d�|�Ss���Ȟ�4L��2�^���a�dpڈX�s�@��+G&��Ml2�kӨ]���N~X�,���t�tM/v�s3l��r���Ʌ&b��f _��}\�{G�%
Ǽ���;��c�'�0�[M��N�[�v��F�+����3�ߕ�[��(���6�l�.�0��.��ܧmp�G��%m^.c��>�}��-錿�f�������+}3+��?a5f��s�	UWlFD��nl�؞�c߽�c�fJ\+��׿;��m��Pk>��F��T��4�|��9�ʺmY�׹vԹtz_
G���޿Ov��OJJ^�DN����,Fs�@��)1ޣG�D`��@�"�z��۵�`A�^$��W	�����(9}�^�Lz��������/l��!3��k��������4j�݊�S�.�Q�>���ϒ��{��C�7|+3�e�4@�;�CYC�}��{�˰ؕ��n��;U����a�zD8�u�9�H�O���b��tGqF�5�;:���'�%9��΋�*��2�ت�x4�)J���j�#r���΁�F�d~e���ʠ݄�==�})��{��xb:.&2�d�.�x�����G�ʻ��C�$�$[�s�3���W�p_ҡ��HG�r��
I�u���/{��<4t�A�l���Z�t��C�@7��	u��H/�}�e��ip��LL�s0o�5OM?������a�ΰ§Z]sZ�
������B;�Y�C3aGqU�+-ti�1�&�;pM�_%���֦�2v����&򵦂�u�|�;2��\��d�%���P�E�*��7z���HQ(㨸L��Ve��Gi��V�:�ꅖo��ə�fa:#�T,$U�{s�N�$h��.�'oM��-�R���e.�֥u\l-�sb(�6�κ�&T�V��S��S⚡d���t%�.��sԎE5IV7pm�Y3�zm�"�;;1,�uk;Y�W�z�Q�p�u1\�M�[���S�=�n�R
򅁷��t�V7��$9�ؒ%��T�GK�S��EHroR���h�WW���F���鼦������Vȫz&��Wv��ob�����:��mc�5�'6(T��V�Dh0z��:Z8��`�u�%N���pA�|-'B���E7p�dq�%j�Cם�7S��C�]\ySuf;J�ƈ�f�WR�(���1&�utY9�a+UۧsQC �CL��D�p̭�_sm�ȎJ�6b�\e2�],��<�	ޚՀ$$�ٙ��x��y�|>e������;���o������c��>m7A��_3�Z qA�YN�_iu��h�fS��n��$I��h*ꭝ���W�xVC�5���̍�����R��lN�6�[��n�&�R�Ws�UŻ�ZSI�e��}f���Շo+�W]�j��b����M�,�F^�C#QI���`�v�tw���9G���4s�q�Z{�[V:V$��4�;2wgk��ڷ�.GG��&e]�����;���ڊ�Xw�6�du�AL��(�㕄�tz�CS�t-�PGʅo5J�=�:Z;RV���:&��a�{qN)ۣ�d�D8�o2P�[�Fh�3�U�Kg^+��q�xR��ۣ�������o<���2H>�8��S������I59�t��j��`��E��Y/�Bރ)j���gNZ�Z�{𳎗H �T������� �Tz���a��1שwB�u�@�� �>��2��F�����I����P���y龡-�,+�^�[L��:8 /V�=+{�����L�U���k�t_Rk7�{��w2_VUm��[KJ��wV�![b���&�+8u����2�fm��9��*ʡ9��O�*Ґ�L�9���x����m]Z��K���in�@9+H�����k��� ���Z��p�=a���^n�r���]t��
�����Rr�b��*z�-���G;;lm�p���nV� fT���sĠ*h���F�a���׮����mm��Zvũr�B�L;ò�,e�ᶨj�eX\���x1�p-�e��2oC�j_]_|S|�ۂƇ��'k���q���;	��O�!0�,�(�TL�icݻ]vv�뺍+���;tm����n���^�����E��ob[y��y�]��Ͽk�g������~BR�H�4�4�4"�-�BЍR�"ĔA@P�4@QM 4�KI�FQ#M)E!E4@�P�!QBQJ#AM�IDM4�H�KE �IHRҴ	CAJ�+B99"Ҵ%@4Б(R�4� P4
� ��U Rd��RPPP� �A@�R9E��@P)H�b4@}����N�l�>�Hfsu�E�DTr��cOq�/t�MnD����qJW<Mj�xg`�6�f٧����H�[�s"y�ws=fǝo�_���9gQ��q�ӡGP�P��]�bb��9���:�;vvGw��N�v2���Ţ4Y��=�}>EV�mgVTߦu��ʍ徕ڡ�n�^|{������ _:����jp5��3�x/��Y8H_�w�o)���*��W^y��#�+���s�5�f�T�0���0��N
���B�U4����#����,���7ϻ�^I�޳�����ʄ<�ׁk��=+�"�Us>��4T T�׵TV����F�&���M	��t�nh�7-�����~X7�r��)���38"[E��w�,>��;\q�Jѕ�BXb���G3�WV�*��,�6Yf�qV�R��VW��F1^Ro>U�;ReS�V�@9(6e���@
:��*�ˇ�U%O���
C���_��T�
���~������+�x�w���H-��]A��$ �a\+Y���5.b�v�^��W��v[�V�TI�IpQU&c��Xg���+�;	�'�`V	�{��׈M<b�ܬə��fDsͺg����,1-���.�LN]kC�3\��CD��*���ݏ�4�������^u����ym����gQ�멜3�Wd���������|�o�~!0�[y�af=���.he�էw��M��9��3��{��:�~ӵ��Ok)ϣά�%�T��ê��Td�t7�/�}�ƕ������>q����(���i�U,������qGE�<�@��@H��#sJ�z���p���\ޙQM�-hBpX�Y�{Do	t�{�|^�=KT�=�Ņ�˯��E�q�=N>^�N��p��RC�;�9n��ݠ��e�Zr��.���l2���������wӭ5چʶ�
l�����E��0��d��wpi9(׭�rc����\�Z6�	[�x��|�UnfA�P�����LW�ւ�Wm�Y:-��׽GJ6�����M����n�ΰ#ن	Ƨ��Q�Z�PL�UwCJ/ճ��i���dw�[���2���yf�w.�wr'�
��OvMΥ�>��F�]����.�;t����N�%�����x=�V�c)���}/T��CY~�ʬ�[�$�\c�v����[u_L�5SHЫ)к'��uu�}��c>i���g�tKה�fWb[��G�U,d+k�����8�m��I"�v����Ҧ�}zOuk�՗�tN�!L���vq���ܤ�O޲���	Q�`E���9����Wq2���0��5�$���W���l��I�8��].�1hCok���|����;��[��i[L������(C��_2/d6�:,�����_; �\#WN��S�j�8��g�z�$�*}��d�&Gg���*K�y(�C�U�$eWK,�X�����Gȸ��lԉ6c�C�G�/�e?���Zj�T)V�	��r�iyE�S,�5����*����Q��>4{uի�/�(z��(>�*��ۡ�Y��{��;q.m�V��ޫ��N.�ր�_�U��i���ωu���9�Uk�f� �^we/Awݮ�޼ww�S.��ڇ�!](2=2`ZB�<3�~Y����ܭ�{�L�:J�(��{�c��ʱ~=!x�<~�B�,��f�Wk|O�n�+�ߒd�^f�.x}���J<�s��+�q�C(xy�d�M�c�nq��K?fF	�ζ���B�Ց-�B_"+�t�o��d�3o�A����3+���S��һףF
�>��V��<�k�m�lnI���6�c��p���W ��be����8��T4�z}Y6eu��.�g�s�����u�����+͕�1������PU�s�\�32x�H��P�٠��{�\U�h"	���ެ]��ƞ��b��4/^�U%��Ư�Gw1T�df�N-'�{�y_WE7��6��&��6�R��N�|�r��U��I�_t8i�N���[��o>�e�.}g<b��
˔/�[����L��C��r��6���X�4�������E�6�[�l\8�t��p*��j<�Y�ߨhcd����l�D
��h�����������u!�������9U2��#�����$W3r��rx����1�F��Ε�Β���:��������ULDpQ�0��F�p�rr*�&�m����y�燅/ݿ�a|ۇ��7�#�=�!���*�&�оva!v�7\nvd�t|e�׸ttU��U<�wNm�D��}W1hʠܳ�_Ep�e��Ћe��Й�.��E����By�������ܨ����)�#9s�
Lo����d#=�ϣ͖��f�ܼ͡ �!_��I��}V�YIA��r�c������"?���ڥ���<fn��u�X���U.��E�5}.�@��uU������O��⧵��쐲��Ui˘���o���TL�y��bá��[�s�QAH���X�	gj�ᗗ�𱜲{�ʎb�kjR3�ߗ�Ń���W��(�fX�W�\���k���)�5��yι����[Rѓ��,gdh�wI�4z�|�Ǽ��睄��-v�m;L��-?+������*v��N�5{� �:Z=e�Gt�3���<
��wsx*P�C��Qs�L�A�|3��H
��2�ت�{查*4<�҂f�(���Z�&��W��'ҭMeVw�6��u���)G{C>�)W��d��~���:4-�PN����Y��A���;H�}q�?����śRz���P�&e��^(�}�~�_t�D��O>z#O�a����i�Y�I+��)
���{K��'p���'��^�Y�u���M��55�^��z���T�Z�,�4��⪮�
5�E(ev�a�N�p�����ͱ��豇oYbK��2����|��2���W*!v�blm����q�Uo&9��s^�;�x�p�:��..f�8]{�����Q�,�	GP'�;�U��!��m{s.����PFCɶa���ʕ�R�M�LT�k}M#���3�}��~��o6M�֑3I��^�7��u�����g�=+�"�U"�~G�T���ߥ:C�ug�>Z�
*�Пq�]z�yulL,�����塻�)�1��������\'�0SH,$�r��4��m�\�{q�2��ثF^rS9�ȃ�Kz�Z�n�@�j��]��M����|_e���
a��9v�Y�{V��[?{��L�?m\IygbX�ҝ/R�el�J�FG<�u�׽��̍_vG*LB[�G�X̼I�i\�.t0ȯM~�}AЯ.T(Vp>&R;�e*\5�r�e�js��$�s���svJ}�{�wϴ�a��`\FT��T��A (�����S���9}��t�.�S̋����}�2�>�!Iy?B�����A�����1]�U�6+�e�3��B���<e���Z�Bͼ��S�D���t7�,3Վ 4/�%}O�|d6�RY�9��z|�o�v�V%"��L*����4��`��*��TT������=���,��b����f��� �˴�mek6�^g��c~�Ռ�Q��k�U��ǂ���kY�K��QXp6=��p�$g�늸*�[fCټ�J�.^?z���ds5e�)v,��o�K'n�'EWg�{��m�C�	��%~�����p:��b�����+ڗtf�Ip��	����*_?J{�y(m�A}^��:�	���3藆pe��j��!1�ڮǮa	�ڱ��Y���p�s22ߋ�F`��b�+ʪ�~�g����e�+�v�1�B��o*ɋU�g��������ef_�P��F�;M	���v�t�Ҥ\�:�`V'�����u��ᚱ\PX�c��#'/V���R�G�N�дAi���ү�����1Պ���V{yV��������8ֱ9򷹚���o10��%c��}�\ /�:�l��W��508��ڌ*�s���=J<���W���<�ܨY��}[�Y���{�JBFVʺ�9���L����BX��Z�U�}]C��>���x.��b�]ɔ;Ϭ�����SQM0�ଛdV�7^+��c������2��9e,�X��i���p�B�fe]]sX�1���ջ������ᖵort�u��'4�d�0���c2��D�; ��5t�Q4YSU���>�K��
��3'�V�KY����Zs�.a䢁�e\GBY;i<�k�wus�ne�搧g�:T��y��t9Qd�~�R�%�v��U8��\ W����Y0�d���9���-�j�҇����82��$ӆ�P��^�Fj�iʙ*���i�D�ۖ���>����C�n{%����E.�Ӄ���w;���iw�z��w=O��s�qW�[ &�42��-WJ�M��ei𭤞��^b0����P�.R�d{巯|Cְ��qM\��(H�k{��O,a�������W��C�G�@�ſD��eD�}����vΛ�V^�Ev���津#�.)��V9bP�:"����C�mR�/���h=F��|Z��t�M��Es	=t�x���M�U^\�m�k;G�����
��� A��耫��ʠ�z]�N�M�,���oMt��Y�󸭇�Pq�}�6x��*����5�r[�s����O�#���P��K��iʘ��/zG}Mvd�f�P�ު�r�̯3%�F��;_c�ü|+�Hv�{������7�ͭ&g�-X������'c������.N�|9���(��=��1OX��o�غRYղ�����=e�길��_݂�$ey܄�T�9TWB��'���o|Χ|%t�re��W���q/���̤���w���c��!`ƚ@�8�r�1k����E�U��f�����92��Q"8#��O
h�\�Q*�����9���WL�e�'��ˬ�3_��j���F�D`ƅ�u�2(hb=Ӝ��>�^�J~~���O����T��|y�����ɗ�Q�I[���hО*��c�L�Ngv�[\��	'i�X;C�M����TJg�1hʠܼ�0�iR�A�G��IسC����r�9���S���1ĦbYX�ե��/�×q�!nt�[���sZ�Z[�g�3#�X/���[`c�K=���=֖�iWo:�O���(%Y��O�%3d��R�S�6�<Q���_�f��e�[Z�[ΆVU��F���"��wYT���*!��aϙb2b�;D>�S�Ô{Mtln�5ϕf�*|���S��k+X�$��+�7���i�t�ㆩ����`�WY���{�'r�hC'�6���ž A��v*����!���zkw���B�>��jx��t{2.*y�+#o(�U�P��/�ʷ��t@j��_qi�/v���*����(�͵�ۜ���X����,N�D �x2P��9��+EDz�_t�4jۃF
���2f�ԍ{-on�]�6�?Q�\f+��Xҕ�j0V	��y��=���;�t��tA�R~�sE[��y�mb.��~Y���ʈf&�4�FR��!���eH��g�j0)d�=k��0zFU�E�s�v�=Fc��^��a�_��tSg�YT߼\�Lu	�c=	A�uJ=����tq���_rE�N��������\����X��!�:�/��⮝
:�R�jIӺv���o�?w����8ʽEV��2�T�^����dp��pBv� �
�!o��c3�#[2�FÂ��__]kc]�S�˦*�8�	?Y�n��W/�cfr5��&z���ӻc9��֤ح��5,�׃���0u���}(�~EZ��8�oR�]���Rg*,�����	�]��%���r½0q�ts�ȜC�c����(���!�>��@��paqs5���ݟL�8g֪���Ƽ�8�vwB��حƟcē��+�O����g��Y�<�&9�ϧLR�!u�Ʊs�<�����n����Dٔ]�ԁbC�tX��i��>͸�ӭ�2��������f�d�����z��G ��Е���طS��F��T�o)p쇨�2]�������"�Z�BC�~�!2�}G����S�t(V�a9Vy�˫c��Y�����Il�ynQ��4����nR[�X�y�;������ʘ�ܩ�
�t)�	ckxM̮��ox���I4<���	d'�}\�3�Q̢����B���ZYR���@�6��xj�f����g{�diomk˃�gԎ��w!gt�$�.
*��t1��9`xmTĠ��ai"���{��[w����`V!�\������:A�|$��Rq�m�R,�=8d�gk���,�Q;���G�L�LU�V�����yO7;V2<xxEZ� g�S�g�'n�6])�fkvg ��4]9l༓H\�x,�-0��l���> ��|��a�(,Q&3���9�yn��ݬ����6�׽�1|Ǆ~Q�,���Tܦ�ߴsŕ�2��	�qqg1�8�Ż��o�Tu�_1M��S�Q����*�����t����l�S,M��� :�o��og2NX�<�,�.��jK ������ZkdF-�`Y�<l �E�i���7�U,�#GL�ϰ�9�sz�њ�@\���1`��� �-���92��Y;�'A	���邝�o.O��㷪��"
@��͈V�<��:���e+�;8d�F҇6�ŋ����v;��u���*��i*�ƅ��JO{/_\K&�.������t8E�]�K�غ�!��68N�H�A�d�M>�x.�ݥP�)���@���α4�]�z�y��w��R�NX,>�h�ց
��6��S��_g܍�6V�S�[��ڸ��:��������,����7لH&(i�6:�u�eԤ��hN��w81S^�C8�H�\\]�D�TY��o��a��c�
�����w�Z�.��D�pֹF��!ԋ�/>)�,[��ȋ�9S��}��_i�ޥD��������tS�X����`{5R8�hk�~��ߚ�یn�Xp�5�ɦ�A�7�{&ٶ��q*�60w�cX�C����.t�������ː��,�	gu&����yٯ�ص˞��Al��ˈ絝
��C$�4T�t�z�,�1�am=\��e�".�� s�ڂ& :����l�.V"#E�ܳM��J�R��vN6+�c�������s��;u�M`�`�.Q��YMV,�Vjc��@v�3�Р'���u0�SU(X�;g�kx����7}'�(��t1"�(�}v��G6�n��]�h<��*����A�4�j�쫽�h��Ve$�wg&�,�`�+�Y��m��u��	�V�@�/BE��y���m)O`?m>���F�F�x��zcY�&��ܴ:���z�Z9(\u��N]ٝ.i������o4O�mK@�Ny�������V%,3�1Z2F�u��y��Y�Dm���j�Z��Ϲ힊ă���;�P�F�P�8�\ۍ��^^֜D��[D�ʕ�s�c���U�cIh�nX��m��JH��:t%�W,��Ib�.ؒ��5�F��\zs܀�~"�4��hN�Ub[EY�R���7EIFs��Y*P5~	ll��b����W�AR�ɬ�	�Ɔ֞�䜁��\�P��0fDW*׳u��[Ѡݔ�Ҭ��ٲ�j*]y�!/"9h��z���v]�:s�z���ßZɡ]��o)<{d�Y;�n*U*v�U�,>U;9�X�f�ޔs~%*�:��d�%a��U%5�ݝƥn;u/� �{\N*Re�uь��xs�7�BX�{��/��
����|R��R4 HP��B�R��Д��E#�P�CBҁH4�RR�B�	B1#HД�H�)E4A@U4�4�U!JQܹ&J9 �����JTf �PR@Ѝ@U#���B�-.C�(*d�&H�����～^�W�ƆN�Ec���H�y)��Qጞ�(G���:��t�8JA�(��Ń!F�Q��V��ɍ2��l��tj���V?};$̯F�!<`L�n�
eUq�FC��X%&^sP��� 7�C��z<��p�VWwf���a}:�j�nj�t��ۼ�+��/��L��z��e������n�i&* �Fe^������NW�PV�E��^��;И��Xϲ�X��@�Hыjf��~�&>���N�x�a�p�s2W\OO�F`��b�+ʭ�t�`�$�ܽ����l�%a�I/����`������'���*�}S�!I�{�|G�"|/l��͓�z��U���D�Ɣ����b/��������=b���3����`��N�fUc|�ud�<+���7��+h���SO�ꂽ��=���=�T�i���Nil���t��=xg��ET�#SHЫ���f5�~�Ȱ�Cn�t��`GW�>3�W{��C��4�L�ؾ�"ʩY]^N�wyWR�Q��P�I��ELC�y�XA�@�����}�!����Be	.#�ς�R�"+�U��:a����m7��:g2�νU���Xt�٨^��F �A}���;@�e_�T�����݈:̂v|���ۆg*R� �vpt��}�o��[��"�4h�CQ���w���FW.b�&��u�]�À�vڒ���z�����j�X�/���J��z4��g]{�׭����|�9�G�E�)��FIe�2�è���Mk^�K�Ht���z �hH�g�,���Z�b�J�t����*�T):
��/�Nvߕ�g�w<<M�~�)КD?��u툓�G�Z��x�p��\2�NC7|�)S�]�/f����`[u� .b�t��X��yx28^�B2`ZB�<1-�_�t�	м<����3���[^��Jyƈ��s�
���3��-�%3��VB2u�HSz�/s���B�J����ez���r��<y��ɾLwm�Â��Y��G�>��s��j|�0����ߨ�u�r���k�u�*C�nfW��J��A�v���˶�P�%�Ni�R��r��Y��w�ȝ.���݂�#>z�@^�-Ŕ�A�4�ɇ�T�h����NxcoA^O٫�l���e��K�F���y�0���w���OG�BV�������߫^d�w�2m��7�����g׈���t��K����r�
L�}��ɥ6�Y�|��x݊�/�L���na�*r�8R�e7��w�PԎ�/�F�ɟ<ۄ%g.�u�k��,���	�M����H��;B����h���Z�-p��!������D�ͥLA%��ٸ��{�{z�t����Z`�����ƣ�\�c�M>���N��oSȰmJo���q���G*��|t\�
~&�pɈ
�}#�`�Eg�����b	��S8���,M��S��Ϧ^���X�1�D,d�]j�[}�<�v�y�yϫ�eO e���r�p�ǙӞ��0�ID�Qo����#"��~�[��im���﯑�ZX=���K4�m�9���e�Ţ���f�!M�t���zT�u���M^�B����B륐�V��(9W�Q}�@l8����t�Ԑ�s缂���<=eП<�)Tʺ�Y&����[�]��^�PWZ���W���a~ɯ�9�#eV�;�� ��e �H�<�U���9������F>̼={/���7Z���g�݉���JWt�%W�HlgР�/��zOK��w����=z��q{E�{'��O3bI�q�/�G�����<�΋�*��2��T�/M�~������L�P/}j�6�o�7+
�eM=�}(�hf�0#�~�L�+��b0�Ek�S�b�;��@����n�Ct���P+�H���l�U�9�s]A�GU�}y�j{����_�D�+�\n��ǲ�k�`��%�
���:qۇML��U"ꀍ�[��m
=���jp�v*�:Cw��sf}��,���|�Z�/S��,mq�έ�c�-�k���m5�ǥ���&�ʥ�B<�xL��]��RH��3\�;7�'DL݋�����	��e|�T9g�$X��)
ΫA���.�WN��{r�'��o�mN�cǵ!�ڧ��Ѩ��유�F|�Z���A��X�Aq��+=[�ڹ6��Fy��9�b�������U�7���ype"4]Q��=),gӯK��L��.��4����&�v�=B}lX�{P�}�u*n��\\\�z�p��g�1���;2�vC�y��f��ù���+��I�s�k��>��a�|��x�8*b�g�T�>���'�����Ny#��% xHM&�H<��?ϋ�9��OJꋞ7ev��T�����~�}��Na�DF *K�Ct�2�=n�X�P��ћt?��5�������
���}����<{��s3�R�=AP�uN�P�Z��H�x�c{��,�wv�^I�|�2�p����Yf�NU��;�������Epze�à�*�`�6�w�Յ�W�j��b����Ycm&޼�N�)09w|�y�䳇ƕ-(��27&�+�y��^_ ~��G�1r�2�ǸJj��Ե����o�
���=ޥ'<���@��tm�gov͕1���:��r��=g4���+��1q"��܍H�ur먂��ʩ���9�B�/!��R|}�1�>�*����c�u�B�H_�����k����;0Y�s־w+±;U����wL�J�ࢤ�t2���S����ݺ!,˛�ڷ;�K�����GX��!���W������}�%k����S��}�����OYο>M�|O�����	��Z��4��e"ȼ�@=�_�{�TB��T�O�;;jj��&ݏ���jq�vT�HSkƚЄ�X{*[#xl�{���>���[�R�����u�}�B��R�q����n�Tw����cF�69
w�61zۨ��Vu��|9�b+�5��ʥ�������`zsѨ+}Jb�G��b꼦��� �dB�Ló��e��Þ�.K�J����m���s���[��C�c�!Q�V�Xt	�6��T��Ü�`��%S���"�k'���w,}�. u��8��0N5)���5��{ǻ�`�ez=v)��|Kg*��dTH<��!#+e]O������=��Q������6���=OuX@�P�_U����Y�t��8l�i���mc~x^f+w�B*�Oǯ��k5s��b��!�;��<��黻��n�IϘ�Fl�WYx���m^�r���&�9�if�qɲ�ZpfY��f>�ż�Y�m(�v
%Z��χ/p�4����>����	�] 6�o��m1���d�{����q.�[~���x�.2�'��p��[�#B�p�B��fU]]s����>r+�v����4x�Jj.�Ϯ7-W
Rs��).aNy1�,7����d:��w5ngljo�Y�c*�xX��d�A�:��=}������2���)J����a��[S��-����S�J��]e
co}p~��3��t2�T��J�g�XGigiH�{Р-e�Z�NQa��=�U�� d�����v�֔=�D��,��qonk�F�g):��r�5�BV��[A�0�wOkm�x=��-yh�J�g�)v�h��tU���YV1)��s�ȅ�|z��S+����
�XO-Tʮ�>4�|f)���Z|+�=ln�{- �[�6W�D��u�怗+k�5����>�'�=��]PՋ���K6��[�&Q�n&��O��N�fǇ�0%��H7�μ�VÔ̡��-�=��u��Â����=oG]�z�#��:�x�L����i���1U���'Iv��z�E|C�մ#F��zL����GWoG�B��.}������{���us�b�A��[��9d�\�0U��!y�7�6�PI�����ۄ��R�ۭ��`�\\�s<`��un��'>=���(��R��d�2�f�g�w� B߆��!��\�%N�M��/ͻ���Z�^Ű.J��Qy{/��j��z
�h�d#^��W��ʷS��ַ����׽4�_�x9�@̈́r��ˡZ)qR6Ϣ��_�u[�%s���MW$�ZO�K�X�[|s��P���L��w��귥�V�^:G��_w���d��ެm�d�jދ3�Z�&V�}�N�"�U��/Wq�υ�b$vĈ�����]�]����{49��k�]�)4��'�����}S���<�";�|�VG	`�ؘ�˛����e>3��a�6���S�H�7�s8[�̺ٶ=����eS~n���­>�=��nhF����J�B�n�%U���,U���;�6ߢPk>��bє��o���@-�O�t}z����ʀfޟ�3�`s�*��e%*�*!�� 6�X��V�ݜ阮ά>R�G���^g�,De��L����$�ֱ|J�z<�~z�����ź-��̰5]���ۨE�8���� =U�N42��\u�k��Y��#�)�����%x�JN������U�i{iS���Y�ƺ�~��%oJ�ϴ, ����ݝ�^Sܺ�JI�:�a�o9[��3bFD�G�����oCl:7Ľޛ�kܙ�x5q�D<�^Ci�2����	@�Gp���Uʽ�
b�eX^����oT�(������O%}�Xt��%����\F蝇�/zy��E�.�f�Vxx#n��*{Cw���L�p`�|�,�L,i��h��ͽ���J��鎵9��T�Я�..�t���)G{C�0"p�{9l���ܭ������t<�}�z��f��x+ҏ��k��[\0L/��������ǫ�^�~��P���M��H�]C�%��i`)oJ7��e��Mm�z����U���5�����{�|L��J�p���
;���m�ϭg�Rz-C�uUE�q�Jb
�"��0����S�×�f�!ʽEV��1T��]��v�tQ�����<��W׃^�٭�ri�2���������>dC}7�U:�_3N�p��d�c������S��o8��6���C�t��,HI<&��\���C4�&�O�>U+���`��eohAEz������a4��`g�r����iU�;W݃x]f�z�<+uҼFL�ly����� S�c/��$U�؍K��@�����+�
T���L���W+�ۙ��m\�>��Xр�v���-��ql{;0��W�2km+�,v��ya��aV�6p����@�p��bc�ZT�k(�'6�������_���$��Ŏ��}�-�B�_h�
����zx�AQ�a�ձ�l��n�]��=���-��:���Q96ZO��������8/dO)ۺ(��\$�g���䨾{����\-�N�����k*8�_�^f��70��0.#*b�ry  �u��|����R����?>�yis����2o����G2�U%�4�P�������Pj��,i�7��[�M�v�C�������+�]��T)؁'�\�}�p�������+��6"���n�ߑ�Vi���=u@�utz\�	-*�u+��;�x������P�:�%<��s��* ݮ,��g��zW"Q�m�c#Ǯ�}{�<G\�7�ʪ�R��L�v~±̍ivm���Sj��v+	�HE6���	g�
C���א{+���\{זHV�y�^=���o��R�q�r��vK���Vۼ���f/�,L)FR�w~���Y��+޶�Ey{n��`���J�����}]z&@,:�qu+�)⬮��gfv/n�*e��K���+�U��!�a�U�F�t�sup�����sy��P�N�F%��޻hZ���VE�@�|�I�G�;fchgL�ځ��ޔ���ڣT���h������ka�{lN��|�Nz<�5��Q��U��PI�Hq9��ؐ��%l�KF�R��*���G��/�=V�de�#0oq��8ޭ�\��j�R�*��a�u؋>�%��-@_`� Y�`�=�
�g�8]N����7������w!���U��L�Wt4��d9WփϬ���A�4�$f�ba���9,/�7n-��|i@���Y���U!6�t����tUi<)\>�"�t����Y�(4+�v'�{W���w��������HU�K�e���HШ4WPD�)u��Ձ��U������j�4����x�T�Pk�/P�9�i2/bc�DYU+>���B%��k|PŽ��k<�|@p�(����z|"9�Y�'���a�fCԢ�r��� ��gxE�[ն&`�/��J���(S��p|�s��O(�d>�t���6�4��c���*҆m���v�謓ce��&�d�k>��f�WH��M 1��1yNi1���m�G��{�F����Ϲ��*�m�zځ�v�E�J�Դ�,d���j)JdϪ|z�����Q�4[V@��
r_WK|ӗݺ]�&	/y�p��[R��RU������_����7rL�=R�u<zw�Wv�,<��\5�e%�(ʙt�x�>:#�%��_u�7l�wV:>�z4w18Rŕ�AQ
ШT����]��v�\����B����������m]s�5�jXɝ�w(3x��,�\�ԫؿ��2bu�m}�P�������Ջ}{V�Q�۩I`�8�%�ׂ�$3δ'~c�|�-H�.�G�ܙd�O�g��5�)����5[Ε�=�x.ѵ��2�6�s�q��:�LDH�"j+9^���Tc.���O0D}6�L��=d������.Gܱo59�����B�OK���4/�L �A��m�3�&S�L4��iժ�YʘC��{�Z��Ճ��y[.���qnGȧ����_����Ӣ��Q��c��|a��L�S{��|0�B����VH�}:go4̝�/�F�\SV�V%����=fus�t*�o7�<+#WX��% �0딺n�Qq�[R.y�.�.�(��}x�l㕼-��a �S�qPy�Xt��]ä� s_X<m<����BLވ��wVn	3�K^���/���:4��J�M#*���白�X5�O���"�jl:�	��'9Y�^�Ŏ͹��f�_vWc�)N�:b���Q2`���s'���l,��σ5��vnS��1��yw�r��ù�:��5H�Td�%��(pͥ��.��8W�dt��Y��P��Dn�Uҩ�8mad2u����:�E��Cv��I�Ӹ�b��g8pH��d�W1���z�gV\�s�J�KS����Mέ�5t	�iD`��y�M�.7�4�&Q���C���:1&r��j��mE�;��U�[ǩe�0��y���Aͥ1L�+���!=J�w��2��]>6DI�ef�唨��k+��ާҴ:ٚ�v�(^"L;$�Yw���Y����
�B���S�Q�jZ}���N�\,S���v��7y�e�9եt�n��O7WY��V6Pu��Vp���M�s��[���\t`���q�j��Mh���B�V�t���Zzj�C&[���K)Q�J�Q�itq���;�˼�L:=�b�'L<�;Վ�a�p��AYV0�&�d&�R�������u�Dl�8�u�}&]Ը���޺�R%���f\V�|F�fe<g�[[/k2���(�kv�3�O'�ڭ�}��X�ˈ�(�����r�س��:$.�&$;����g�����y��Ɠ���i�i�H����n듹�͜��oI���wC�vV�F+V(j`�7'KT�Rwo��rU�1#.*�%�����z���}��#Z���$hZQ��ZA)hJ���Z����F�A�i �h�(J��L�)J�2���ZV��J�j�h�2J�"J ��h�J(�
D�)ZR��3�)B��$C!)r��2ZL�F��iJJS'$��$�)2rQ2&�� ȪJh�ĪP�2r(��
D�fh������V��}w�G�&�n�av�Ջ��c���k$�)��,�}7x�[3k�Im��%��ɪ�or�7V&1��̛d����;�q��o1U���dV�p�>x�<�"K
���Ur�{}����)[��<s�;J���kݑ>��Nh�� 58��������TZ���o��?6 �
���	Q�g��Nx@�`/�f�>�;����^J/8����r��������<�9��>�ww�]"'9�/Vd��KO
Դ�)f�1{`�s��s�f�u�e:t���ܒ�"^ҭZ�s�����g�x}.��>K��5(+>��ᰯ��C8��r[���DVU�d�g�O�}˧v�n|y츨+�yH!��Y�L%�j��/�\�e=\ l��މ��x>{��X�s➍��ǾBx8^�=i�8xW
�UY�3>���_e������{����b����=�L��b�����PPs�N��M�#�\˃��4���
�-U�����.�[i�8zv�ۡ�}B3����N�"�U�/Wq�>���#�:.P��bu�ya��U�{�'�o6��ω��ܻ�Ld��|X�Ꝅ@���!���p_�Dh��n�7s�l�*�)٨Z��ZF��2��|ՐC����������/Wx�)x�z�Lf�M|S����Tb�]@��r�.�E�su�@M�)�(N"�+D��v,�n�+̺�
����mI%M䲰Ea]�Ѫo=�}P��qn���Ѭ��g�@�4k�Tz�5\�=!��ן�Ӭ`��G�Er�����Y~�W�ȳ�����n�>���F���|J���]*��T�ӛo�(5�\��O��ӗ�=���'��[gz��WM�49�=V���(9{���k�[�����b�m�M�mSӽq|�Lw�0Dz�L�**5�Mn�|J�|"ϒ��ʖ�fo*���o>!����Xyy[�!B��d�Ao����[�]Е��j�N��_�-D���D��{������b��B�>�DԞ4�<���Pt�oIϺ 5,0�.]c$��oYƯ���p�[��Ԓ�P��ר������gEacN$�=y��z�U�z��ۮ���#��2�TC��g�\��(۬	i2�u������k�_`��Q��\<.�����q�=L}&/���/}e�x+��[O��ǥ��И_*���nA7)\�����ǫO]�0'�ׁQ������-���d�,�x�6=�������U�ۇ��4��PX�Z����|���:��Z֐�5��4��2��ғL�o9��&q'R#e�Ҝ���z[45R���`���$<��GU�\�g�mq}�Ķ�i2��d���ʓ�����K�N{������,�L�#Oo�� �X��9+�Tt:��&V�be��7Ѫzk=��rr�������l�4��ԝy�����a�c�V��У�jt3�\��bs��*�׃ܼ�<��Dp���{[Ľ�������/��=�V�JEW�?���U��%}^v!�*n�9�3^�.��]���:-��jȲ�c�S���W��Tv�!�C�w�b���I�X��x�Ӭ§�d��lm���6t�}�;|=�T,�SH�G��J���ˢ�U� �T�k)ߓ�~��N�\�vN�%���ʟ�*��9�T� Twf����J=l3E���ɜ�v��\�=�c9�S�k52���񐞬@�g���A۱B���p�Vy�]뗆���j�����������b,�TqV�R��na��t�̰�A�v��ȃ��DE�@+�
i���6�9{�^�|	��Q
�����������3��)N}�*󹓙��|�ՁR�G�Y�b����ym����B��I��FF���,SX��:�:�Q5����������w[�S������e��u5��F��z:3�w;�C��˂���|V��.��|֧/��CDOy��~�$�ܻ����S�9� {J�ZE��+{����c�r�v�ֺE�[��n3Lٜ�N"����ѿ	֍�M@Tpbo��}wy,v����wDIE��e-�z�ӻ�����[A|��:O���+q(�qY���eR[����m�ܭ���WN��|D��k�� ��tv��o�O<p�8,�(�Dv|-ǥʴ��c�|�s,+���~.i�Ծ٪���>���t�i����N��@nj�t�n�����o�\D��������r�U���U{�V�p�y{R�Dr�q���J�b�M�R\��rU^�T����xf	^�h<��Fƒ���t�.��aʦ�p�s2W\OO����gm�.ܒ�fF߼|��LW�ւa}�e�`|eRKG�?0�� sP���G��F����4���#*t�����lb>aV��3M]��d��_Z*��x�A�4�$h~���b�\ӛ�v{;i�a��!���y����pN��k�b�]��|K�!f���U�y�z_'�;O+~��w���{���~���x�.2��颾�dj���WT8S��u����,b�t8a�)J�f������]���Ѯ��|�孾�t���Y�s2����K��N��+������).�k�w}�j��;��i)��G!:���sւ�3�T]�͝�atwi��gT� _]ՙ��c�D����s��Ҕy�Q[�?jט�K��yn��MM>�z�׵-W
��f%�*}<�ɖ���M����5�Z� ;�ʩ�f���A��,H|����fK����&Gg���*K��N�^�>�E��nT�Ovf�õ�}[�p/�"��Y*��*�1���8?|�ppc�uL�,������ov�	��m`�"ϪSj���L�M�Du�T��R%�}�������0NӚh�a�{�������I���e2���%�[AS�<U<J�WyX_u�_o�*`�>p{�{��l�{;�ؕ��>��� �Q�6��
�Xh�yE�
��JƇ��(:
�α�T�uN(��_A0��[c'�6��N�m{����C��9�W��Pa��t�w;�؆�� ���3�q��·�!�;>af�S���*N[��MX�ѻ�|�}Ȉ��-_�W֐@���I_VK����:��
�����T}u�n� ��f5=-�Ӟ��c޹��F�aU�-tJǡ���0l!�p� ��N������t8z/�J��3Z������g`�A��N@�`(�t.��Ղ	{RizM��ݺ��XDo6�ެ9�A�w��d4��%��$����w����.�E�xu:��T�E���_}���|�mv�M�3o������8�4Ⱥ�w�]�綟cCeƲ������Ӆ�S�U�~t�x�s�G�+�P��Z��g�W'��t_M�zL�P�=5	��M�61z�}2���x�:.���|�8��( gut��
���ur��WU�7�;�yV�3��w��.e��쎪�ү�8�^�u�ѭ{�񾢅OȑO����W'����,M�N� S��z�V�/:U�q���iV�jNz����6C��X]�a#F�5Gl�۞�/����,Vͱ�3yb"OZVci�P�� ��uP8��@"���ޡ���%]�ʺ,U�-⩳Nzܻa@x함T7��'���t��'�t���?\�Hb�0�ʺmY����d�����RPr�*!�d!�d�oח�߸{�p����qʋФ�x��2�^��ϣ$ҬഗK��<���������=w�%}�^�Pzu����!B��@ʐ[�0���b�T��!�xp�K˸�3�1��ݘ�fy}�t!S�vzΊN��Q+�$63�Pt�U� �mۋ���t�	㖅`�Xmp�n����Y�q���AR�H�[������Sj�����F�W���i��=u�[r�����t�np�e�RUַ��z�k��D�%]�f��U���vn���Gc�����-݇��uW7K�f��ޕ�Wg2#�fb�n��E&/��=r��1_W��Ȳ;�Q��������������,�Zw�x����tC��Y1�B
��j��
��sǩ��ҕ�4`��n�u@ckh��]�#���۬pْ.%}�:N}L~-b5������cҪ������հ�-и�;#�~*$�]=�^ٮ�$+�w5���3%���zs�:J�*�
A������{r[�G��Y���w���~�)V3!/��4�9�;ᑨ���'(;��G�z-CY�kB�߷=мy�W��z�$h��~�����qV���y;Ґw0*"ob�X��ܪO��t���bA��Y��U^TWo�!fƊUr��u�	_W��aʩ�D�u��3W��v��=B�F�K<�|�*~��xxE���>!��xʤ��F��u\�`��ס�}��0�X9R� ���YӇ/v_�ʜ1K�֦�ҏY�<9tX��i�ҧ�E�<i8�V��/��ɕ
���_^�NYJ+�)+l�P�����0W�ǭ��WV�Ίzc�,�s{x?��)�ӯ}x���y�/!�4�/��IF@U�w>���:��!P�����h�w/n�,�m��R,�:�X�b�:���U����t0�t�a� ����*U��V`\x菏㭁V��> �L��L��&d}�sż��܉�ټ$���AZ3������1�=�fpw<�
�4(Vp>&nӗ�S�v'�^�r sYH���K�`��x����?et�R�}��������b�fXC�=���ŧ��]����`�u�}e��%S���>�u�r8����~��y	*�^��t�����S�_4՚ў���,"��G�y�����?w!gt�$���(�����,��z.~y��t%Wu�z�D�1(2��Ϗ�ڀ��81��?��%�ã��]w`��*�r{;���s�H�=+hmwm:
�K�t�t��n%?Y����f�+�t��W��"�w�pL9?m@^�x��� 
Rbz�_q��*�O<p�9gA$}~�)���ɝ�f�ׄeqUƵ�y`������|��aW�%�QC���ݖ��W�M^{Ӓk�N�gUYj�W�`o����?uE��G++��P�ޔF{�'.f��Y���$��^:4J��W�1��=����z�l����<|y|��3 -{�����2k��_�ګ�����$��(0_M����k
x��4�<��l���mv.�Kc]��1΃�fa��|��U���I��c�Vavp��:��J�v��V�ѧ���LS�s$p�{�Z��\���]\�Z���e��d�9s�z�)��sA'+ϵ���c3��{Պ��*���=),����G��| ����r�&�yJW�>���o���ǡ��	��U��L�UwCH&C꾴Y�)D��O]J�@�\�f-���p�++�Q٩�ɹ԰K�Rj�L���t]�:����
�x�g�.+m%��p�5���J�,erji��PW�9o<��	ư'U.�*e���Х��V�_�����9X��>%�yuu�b�`ƚ�}/T�Z����`��"�*e���'y�
,�س�#�x�|ݐ��o�"�C���r9�Y�'���~L�^Z��t6j��\��w=��ς�4A>����!o��I�Z���/�ho�2���
ex'��8�v=����ҕhϛ���8�q���$�$<>�墓������}:�4�Jyns�����	D�$0<�'C>�ȭ���YuѺ���$�u�}e�-�����د�;S�n1�U�Y�����3�a�A�� �uH-��,*yj�rЅr����yB&�ܺ�yBGu�˛S�Ρ*u!��c��7%��F62�ce$-ejQ��w�tؾ�[�ɎW��sV�v5Y��
yPU���9�����9;�I�̓���L�(��^gt�+Re��[�1U��Aa��.	���.��|�yw6�ʊt�W�n��ķ�Y���w+kٯ%�����WD ��u�>���Z\�d�y���+|<�2sH(��Ym$ɮ��!K^��5��j�w��Nź�y�^��#ɩ�h��4:c2�1]�)��O��+�}�*�u��{f)-N]j�˷����s^w�u��U��;���ü|+����['�#�U��q�����s�X;y�{v(}<��a�'+�e�����邜=��&̮�l��E7T����©e��6z�f�p���\�Fv���`��sm��g*���ZG�#�t�r�.9v�io��S�Ҭ�d�I�aP�Y*����9O*� {}�����#����3]��k�z��!p^�D�M?\��c/�5�Φ���+\��0��{+0n���U)kUuуNz�K�fC��p}��4��~:]�-���L�U[n��+�����$���Ǌ<����=u����ִhh�	��c�=���{���濂* ��Q� ����"�
���+�PTA_���
�qW������AQ�ED��
�+�TA]����"�
� ���삢
��W�DTA_���
��W� ��� ����1AY&SY��J5{߀rY��=�ݐ?���a�{�^�P���JE"�"�T�B���UH��%IJ��IU*��%T��)H�%"�!IE�Fa�$P)H�B! ��)EB*RR���$ITZa"��T�" �IB�DA@���ilB���!
P���(�h��UPIEJ��R$�"*)UP��$�UT�J"�BQRJ�"ybIR��  ����2 -0
��R�J�j�+P���*��T�Vk*�-FV�%Y Y!TTA	T'  Z�4t���Ve�P��
���V�C6��R���F���Ɇ(�eP(Q��4TA-�`�kI6(@2�UB�Y�2�pТ�
ή�P�(c�� E �Crw
B� �@.�p� �� Pw(P
(�h`�*�a�Ek*��5CmUV����Z�����TD�����f�6�)��J,6֪ !�$�U�U���Z��T*���SV�lU�@(��B���J�QEJ��D*�݃+k`l�eh�jl��h[dUUC���ص m�����+MR����@U6�M`��Md%U*P(a ��@ժ�
�e
Щ�Y�Z��� ,��ƴ����(�٘ ����jm���a����Ɣ�)	�J� �Q�TQj0k@�[Y������jU�ڀ�B� 4+S@� -���6"R*Q%Uk)IF� 2�@�s`�Jf1AE6��IF�` %4a�@
�L��VhU�� �TPT)k ���  f�����U�ր�iD)�0�ml0 �2 &��КLT�X �I�(��SU�*�   ���6L �1@��� Պ` !J�Z15�	� �L
kk)J�@H �  51�ʔ��@1�� b)�IJ��4���a4��&O!M�F���2  �  ���T��� �� 4 (�"12L&��z(ڞ���h�jA&�@ʕ2SG�i�b  2��Py�^A1�R_}���	Fm���( A,@�ů;���i�������! !5������ w������@���8>�Lj�k���1�?���A��C`����� �aDd�I !8�2PH
t�6�8���q�@���Ƿ���
 #��t^P%��@��5��lc#G}��A�Y,��E�����)�*����y�]�n
9X(�j��B�Zl�mL��;��#e�-*楛���[�(d�s]k�
2��bڡV�����	m���[Y�-�����	�"�	���v�Zi6 �aj�����-'-j��� ��)K�,�Ւ�5Ԉ�ŕ��H�>�ȷ�� cI��w���7Oj�(zlRn�Z	��ed�U��YIR0�mKO6��=Z��+�VA��.�Qi�Y-��d��sr��n8a2�	CS�c�z͜b��ƙYm]�`���a����UoA������
��!��]7��<{��s1V�sdT)ܘ�{Z6�z�][��C�����,�� �P���E�i�7r%RY�3u�����Ha����؍�N2�Q��*��h^��pPLY/i;x^CfP�(2�uH���(��1;O+
�Z��ұS�Tn3�R��\٘�7�~h��);$<�HɄ�Z�;�S�MEgM��Ā�'�ݸu�:w0�L4�y����c������9�)흧�抶���Bmkr�\�x�U�LO?���'��;�{�s-Jn��m1��m-TBJ���y�I>�"��J��P����/2ҕ��۲]��i�b�S���^�u"����M�u6a��[��L���&:E*2cׄM9�f�%�̊�@�Ղ-��eaT�N
���G�*20��[J�b�����Q�:P���û[Z�D��mn�XV��0IE�=02�V�1��E^I���]�Xw1�31�a�4��sq%��p�cZ�ONiۗN�]醬M��`8�]����ӻ�Z��LX��o.�j�v�Ч�3��f��Ռ
Y�o4nD�̶ʃ�E�N̞bNCE�t@��B�t�6����v��t��n��)����fI�R���J	������\�5 ⫤'m[�/AI��5M��+h@���+h^ܻ��n�N刈!m�	��?�*��P�1n<!c��ª�Q��xR�'�Er/Y�@L�֎x#�MxN��1�*+�� ���pRTM���>�^�mX����\,�t�q(�2�e�����<�,�r�ovJ� �� �#4�&�O�A�yxm�Q�����N�$�U���fVRm^��΍tҊ�fۥ�.�K�f�?MZ�u�@�c[xvB���N�o°]�)4��� -{q4BXG y)�״3"�l�� ��� v]�j+j��:a����n�ȳ�M:Ya	LX����ͫ;���A6���Q�ڰ	�6�ե���	�
A��6�4���+M��r���ۥ�����S�D�^6��� Q�6*]�������eG6��6�l
ՂeX���@� ռ��Ӆ[,��7Z�����/&ְذ���Gv)�{T%���=)��GP۰�m�eؽ� `�+wf�{D-ST>��P�ռF�c[�.Y��bT����@ZV�u�ڹ3 $*�!��E�nQ�:%�A+j�*üӘ̖>�GGwU��8ېV�eJ;�q㶔��,\���Xe_�kB�P�#Yw� ]�ȅ�z���(]��a�>˱شĬHkTL�[2ְ��v��J^Q�H)�n삖�ܦ�eo� TFc�*��m�1���p�إ��UsO#4�v�i��ů6Md��5t]mLe��
Lb���21A��[z���X9ur����p �%ŏ)&i�F��Y5e��k2;*եZ, �9��'a���34��#�Ԫ%^�� VY�Q�Z�fO	{h�r�Fխ���r:`^�Jܸ��pHt��`�p�����]�ˑ:��̄T���h�yn=���8��5�#)fd�X���-���h͕��NL�u��\v�2�1͙[I�4#�<��
6��֎���J�\*��:F��s�2�ZՈ���z�At�үb"�"��v�T���2��\�c�K�9{��q�n\j�M��jY�{C,��]��i�ӫfTn�r��ݽ����z��xh��{ ��T0]d :c�WYfmBE��R�`qkV�ZrF�.�L���=�&��rkWF�P�T��Y[Z��Edɂ]d��.^�5��
�q˧Dg�鵲�"�dN�:�=�,�dуZˡHb^ZQZElx�n���r�X�-5Q�3%�i/��\A[3N�kb_��ð8�0]eV��G�-SF�jν̩��łm�C`�J�wObر�A�FRV����ܚ�N,F��°�)f��v#yB�ª�n�XU�� �W�I��hU�.0H ��%;�.��L؇L4%��҆b:�7����8�,Ź6T�h�SZ���IQt�K�ⱆ���-�d,�TS�h�ɇY�;���̹)%Am�Ec�-:�(kn��ab��x����Ojmj9j�kp*8c��������-�7-\�:9.��Mc���B;��fY�b����	�Dm�Ōۭ��"�����u���1'�1��3��1�Œ�`Pmb�[ӥP�Xo�RW�)I��b�+�k!R�(�6a$C��Grn�
�;��ܵ���������#V�D�>���fkY�E)��9�G@�C.cv;�� ��#n��O2����	l	VR�yZ̏ ����ŭ�m��V<�j٠��ݰ��!��і�LsU�v�v�h�Rn�ǎF>G&��Wb@��ؼ��!��C�6�����@�lŨ:v�l����lj�I{,�LOh0 9x��7E%%	r�nV�^�
�=�k]@�ZJҳ`\a�%���b1����&jx��z������>�L�60���l�d#3Wyx���n&L����6���u�������� .И`ֲ3Vh�Yąнx�E�֮��oЉ�7�|�KtQ.������vh��������p+�	��hP�*Q���=��y�F�B
`T&���M!FQ�qb8�tR���q��b��cn�V�F4+k2�6����@jhnk+m�U��:X5���VH�S1�x��U���c4Ӽ�z�`���"���f^K[��x������;m+ɿM̀����{1�x����w>5���EQׯb݆˔�r���/ �);UwRfhe+�Z1�0��z�n]�n'$��`��lZ�b��TVۺZIGPw2����N�V32V��c�t #����,-4�^�y$��[Wy2�m�rS�b�D�[��YeӲ1� �[���S'1*p�;�o	�Y1Ȳ�&�ۺ`R��)�<��f���Y��]�)	��:�b��yr�+q�؂b���!�m8�TY��`�6&c�lކwst�ԎM���o%*B�4^(Rkhwv鵮�"�ɚ��z14�c0 Fk4��u�'�97EAI�Yn��(P:�/Z�Z�W�-�eͲ�ZHJ�w�H�U�Q�O/[E�m��"!U��xӍ�*�ɉK�Қ,��)T:w(Y�/*m�1��[#�xU�Q�ƃ���C�l���X6��SJýHU�R{�M�.������/t*��(�4q�hf|��
�e�eS��	v�%��ޖjl!���ʻLԠ5A��<���"	�(&N�HTɺO둭tL:
TZ#/oQ�:�;W[�ALV��+fKͫ�P�B|*,R)k�EmC��^��h�vVҳ�W[�d
�!�� [���ͷwOW�P�R�LwzX�ul:i�'m�FSR�A�N�K�ŵ��&���t���1�Q�3.���t㠳Nw���OL,��`	w����(��ԁGl�YV��ivav�����dn�H��K�5P:q⧅�TZmءM*��p̩.� ���ڒ��a=���n��M�U�"m�e�q}v�+r�.�h?�U���lq�+XS���"�C�4�9���v�fkp���T�S��CE�!J��)��eϯ�G.ۺ5�F�շJ�ax���7(�KHw��Ie`�}��²^3
%�:�b@��N��)S[0Vg�,6�7-���!B%N�Zo4�Zp�5 4l�a�����5��V9(m�x��"�����SRPY�Щ���(-����Y���ۘ�����Ct�ܱ�R�ZHܹL3��~��eK���A���8�S��t�#���[P�V�&��-	�#�^Kը^�VM��
a�:��raz���.��B#фˁ�	B��`:����m�ΥX1^�f�퉕r;h���l���b���l��QW�aV5�t3�'�,��� ��%Y.���{�EB��]!lZ3�AAR��e����L�n���eXF�WHn9�
��.\Z5?����
��{Fm]�l8�T�F��،Fe�J�ZN�8Խ�$F�h��dڙJ����ne�۬ �j�Q�hҘw��ȝ�Z�{g��h]�lN���ƈ��Y.��f��/p{��Lr��.���Z1�7D ��: zU��ݮ�����]j��Fޒjd.�7-"#͖���m}[6���TJ]ddT I�:�ñ����鸷`��
@�	Զ���.iŸ#]�����^�
�Ti�8���m^<i����D����Z�W�0��Kڔ�룸��vXة�h���GK�����ƭE(e�hPcf����{>�&RPއ������(+�*ʻ���k����'A;��Ģ�:V6��:Y��ʃn��腪)I�&-p��;!P" Ɲ�n�1�e,`����LA6���R�4)U�Xo�M�Gbʁ-�mv��[�,�+s3`����cJ�\���G0L8#x�bm���fd�|	4�S�4��\���Ҏ��-3"��ef'R��CQ���D��j�@Zp��r���kH���׆��Aѷx�ɸ�Q�z5�ʅ�v��V@��c1n衷�rmA[E���U�
T*�Z�����W�Zj�yR��Ϟ�Q��{��R�aۤ��7�wO�ыC�|�+��C2��ز�cv��I��R���� N��(Il�m�8�ݦwCu.���v�&�o��]CE̠��B�"�.�&�d��㤕
SA�m���ol�L1x�/�*Ʉ�c5Tȱ�(VU�f��f���QmZ��+E@�5D7��o2��jn�DUq��sh���N��iF���5��j���Z�EL  ���Zڻue���E���]^�
�H���~��`�\;vi�u��M)�k6v͚3 ɷ�͑'���������J�pUБ��m�im���8�ZK{���Ik��P�"�D�x�N�ô��eTZ��b��#DG ��K`S*�(��E��0�����-tu(%Ht`��ɛ%H7*��*�`ĝ�	�-�f��]��X��{6�!^mE�nk�+n��6�n"���8�Z��Z(^#Mf�*��9Y+jܣ��Z�W-��{v�F�<��^�J[Z��X�U�($�a��e�Tݵ��%F�n��Ҩ$�[:DWh��1Y٨e]j��T���mU�l��+ݦ���U#k��8�6�R�b�Y&S.�����h�ֆ�[��,�2��M�)�
���r2J�[R�T�I��m%�h�r�l͏�="�r�z�ī)�H]`V�*�+%�л�Nύ�mSh�0�i��WV�CS�)��LU�7�Q��E�	k'%T��:�f�t�*HF��R�CV�Ҧhں�sf��4�;���'�E�n��V60���ফ4cڛ�Г>Ui�z�W�+L&t���u�F�F���tXGZ�M<ˬ��a���ئ?��چJ@�Wpɂh�2�\�['. ��� � @�@�Z5裶4�r��h��ExS�DJ��V&7H��GP�N`�$*۸�][��	�I�����g���Ύ���?r??\�mD������e��O��~߼�����^��֩��ќ��r�p�9�{��}ٝ.�%���Zbc����{���1������h�oL�Pb葷�p�;�����M�Q`�#�|�7�e�� o9[tZ�ˈ1����x��|���c�t�\��F�mp�[�v��һz����H#[�*�΅iq�����U�4�_r�jelf�DB��띢����r���O�5f_\�ʌ��̐ȄKn¾��'s��ɒ�|:�䜟.�l�|ч61��e��������qF�sq��*����u��%9�ޗ��E���
T� 7)fV+Jξ}���r��/�6TYJlt���T'��ʘ���&5�>�kq���Ƭ�h}&���"�a�m�P��r�����8bӏn-�|RJ
Cx��'�Ļ!F.���w2$Hz]8�S<��%,�r�њ�:W,�սt�5g��᧝������"yՁGAí:V��J�Џ��k!����\�d����+�(�!˷�K���̊�r���а�S%�ȴ�]�/iig��\o��+��Y��a��v�(s��+k"��V���Z6��u�hV���K>��\ܲ��N-:1h�u�5#+�����­)�a`�MJ5�� Y,���Tՙ.mu�hel˷5�Dm͏�"<nrh��٧�}��G/�9��s����X-��n�[Lخ)c��;j��\�m��A7$����Փ��k�]�q���->n�Vb��J��P��3l56�';!��5�[��w4�6�7���<����K�m]�ݡT�Or+X8yT��5�������kH�yB�s �.�֞'�GJd�w���Z�+�Hn��}x7�5�ޅ��8Շ������zމ�WDue]��Ή��*C:��m���;�[4)9j��+�ui�g�7��՚�ɀ8�H��6N�b��^���Wӏu��L�x�ߗ^bn��U�5�:��=-��W�b��r��;��8��X&]q=���ϳMJ�]�:b�B���>*�;��rꗗ��'��X *�\�nپ�ۺ��4� ����rwU���<ܱ�Aħm�z�[�A%��]>�s�bw놄�fP>�������;��v���?�l������B�H�3����	��Y���^i����4�x�d鴷fj��9 �]*��)��%���u+�%��|��^����nE��bX�2�q����Z
��.���X|���mI�׏�~�ƫ�a ��w�SI1�x�`'�T�`a�}X�����Λ�ؒ�j�%e�(�A�k�R%�Ѱht�wde��2���j�mM��>��0-�7���-՗k`=h1���uz jd���A×��	�"�Rڇ��0oq1}F���6l�U�����̶N)YC+1L\p�Y�>��4�@}�W���vq´�t����u���X�E\N�}��I�R�fapL��R�5����.�5�p%N�
��wH�Z��B��jʫ޹w��S��:U�t���0fhsX�!�{~�>����{uQ3�M��m���DvtY�m�h�u���y��_e�%k$.1Һ�K@��g"g[xv\�x����w���s}���ue��p7qTVޗR�Nܙ�t+[ިu2x��gZ��	K��l���#� �j��u�I֯5I؆���b�f��0d��G�hn;T�Ȧs��������Z�]��������k��}��r9�0�$OqG�ْ�6�+D?���n�ŋ<�-A�JW>�r�����Y̚񡑳n�խy���f�3��N*�+�w6W.Lp�,1Wgw8:kSȚ�|��Π7Z��LzVE`w}]\�_ �4�bwG.���6�!�R��s�r�Wâ;Q���b�.̛��c�e��]n�&2^I�5�����;o�#�`{�� 
<j�X�����n�'u�V��J����ا.�u`��6� j��w���Ώ^��j��z�p�O�.bOo-G0q��}�vKg­�p�ይ���P1ۼ�Yi���"�Ț��"u�pN��;,��s���Z����U��V�(rXNK9�fv��)����J��1�T;�&^��� GgTB�*�B�7��<w�o�U��3I�	�&�vt��T+��F�l0 ��R��.[h��ϵ.vd��찲=�i�G,����nm��E}�{%��S�8�u�M�vEٶ�_p��Ӎc��W[P�+�'��bB_tɱ�Z�᮷L'ݫ��h�����m�h7܅mY�gUีdu�÷V�kz���YsVᮔձ.�ժ�4��o/@��&Z����J����O�.����m^�4�����"��7�v�
J�+!�j�W8�F�����]�ٵ�έe�ĜD�q=҅��R�rq��q=ډ�Y��I*��e"3�wMj�ܴ���n�0靊�d.l������F4�{�a53��f��]��J��=����ݜJ԰	.���'5�"�*edW� tf���4F�S)\<;�;-\)B�8��w7mV2�]-���O��~A^�]p�z��Ay5(�v.��R�ڕ�%D���ڦ���O~Ib=S8�ů7h�Ԙ�����7���W��)�v�n6�5]�.��E��D:MWα��ʼ���\s{.���A0 �|F��7ݗzD��#�V7�yw�B�:@����⛻)9L��QT�u���j>�eN��ia	n9���d���$�(�k�փ�x��zD���D�Xw�����)��*V4�`�t�{YçLNJ��S�m�j�P��f��];ӊ�4_q8���e1�W���ap},l/:�>8^�Z�L��(@�ήb�R�=��W��f�1/I7���ڒ"�!4�V+i^�q�R���n��k�>�c��*����1�]Әd�.�B��yy���e74Y�k�s��%��7-N)�5^ť_#�n%8#L�з�*[���k��˅f�t#فf`b+_m��Qƙl�) �E��@7J#���l��Fu�����2�e�B@��Kw��{}y�(ĭ�*W��lh�gCGI��wR{��=C=e�hnl��2�151�j��.�5�Ϋ�e��bhXVV� �[KYΚIB�vt$N�f1]�rX6�T�e�*[�
�[ʑ��ݙ�>k.��/n����u}�����;I����&�l�g,S���o��[�[������dS[b���ފ<����t�������*W1揷+���L�2`��*Թz9v9\Z�	��e#�	�ʆ��e�|wc����bb˝���%�U���2E��o��*���k
��c
t�J������4�P�A�|�-ඈ(��iԥ�vָ��/2��u\=����X�G3T����o^q�k#�>�ח�'V��4'����JYg-m�N�G��_�eA9#������X�y��
�1�=ѐN��|� �����n��{�IC���=���6�-r�)g��ܴ{�L4{�F�������tk�[j�5�vu��_�8uE$9�p�X�Πz�)+�����%�o�&!H��dܮ�秵�M�F2Y�C�'��-�6gr�G0�k�κ��XJ�g�� Tݕ8;��c4Y=�[՝Ͼܭ�ޡ���3�=Ki��`B�K�F��%�
G�ͣ*T�7��خ�u��"�n����MyՏ� Q!���D>癫��
̍���p	Dك����W���Ws�j=о�k�0>��^������l�v򯸒.����br�u��>q��-<�$s���Z8�J���̗�\y*�E͌��+�պ(c���F)n:8�7�ޛ�ș������Z���>]I��6il��ҬðΉS'�r#,ú0a�BGq�N��2��E��-=�]��ړND��̃X���z���]g����G^�Z�rB��}�,c�I%ܮ���un�lw8)���җM�Y�U�Y������̻d�J�ܴ$iv�J��t�����j��j�Y��
���#���L�Ǜ5�X��p�C�,A���A'4{&�l��r��5�]4�lM�R�����n����9̬��.P�����
//�⬲�]z��^�Ɯ����cj��N1M
�B�۽*ݮ���ZhGqj���O�:tr��St|�.���0zQy��ʹ������N�j]'qЪ=�|���oï����l`N���a������IfQ�wi�a�l��6)wC*ra)���ovB���)�Wbn�n��Ƶt�23��9GrXv�/�h�b��i��3���zR��:�/�ti��0H�<u�����fZ�o[gVN�\���Ō�cM�x[�b9$�u���]��`�U���=�U͔�W�b�p��YȬ\0M�%���M)M��|�9���X3N�1]���)q���L=�F�P�k��;f���%���S.���C��SU�[��㪞�ss,��,J���i�%�����]�;��9J[��Ji�z�J��ˬ�9Ҳ+¸gRtf���;Ź�%1Q�g� Z�Y/���mn�6+sLܕ
���5Ϝ�lυf���!b�%��)��x�9�W��e��{�y҃�X�8��CJ��}�r;�V���7+r�x�W[��Θh�Kz�ٺ�gh��*b��"tʒ��E�������|�u����M]:�����t�n�]�����z`]31���g2s*�r�/U�!�ϙc�w��Q�.�Sj����,��mN8��_R���8��k�U%��t��4em��t�F��\%�N��_R�ٶ����;`e(��S��(�U��,�G�CT[/+�o�h���i�"�2`Lk�ݼK������g����)�e���"�J��̗\h
�k�;�U�_��J�S8��S�q������ܓ���j�+��"[���'#g�]��u8bm1����b��v�}u��7�*����u�q�ef��*��Er��#��72��J�Y�M��l2�c��ܥ�TQ޷;J���!ىn!��uذܮ��w����#��X��]}�^�^�Ӓ>'��C���,pe�k��`�ePy��%Ggh�}y���>�V�u��T�.eA�iRw�Z黀�2]c[q�R�sf�j]9��0�i������7N��]�u�����jGX��f֮A�}W��ق·�d�Y�:��\����[��º�Oy#�El���g<*���h�U��Iv�ԸU��)�}իb��՜�����d�\�Ԅ�&p�CF;= v�-��R�J�M�ŋK�h����l��r����Ƅ.��S��\#��T8�&*��3��H�K�rCjq7�{j�*���gaZ#쳜f�n%��T��Hi�;fb��;�Cƻx#�w
5�x-�e%��lN��v�gV���R�n�RvXRv5f��L��Lowx������w+�o�P^�R��,u��V���.͋��M{_]�::�T�������w3�k���gW[o\�]������2wpm��Z�g;P�re�+���8_env�̩W�2�.�q�;���9�s�TK>}�;�}ݧ.�2���qS�f���E�'sIbI-�˵DbP���Iwd�����
Ը����s��2ޝ�Hd�o�݀u�w�B]��QN띷��ӹ���I$�I$�I$�I$�.�J9-zG�����%�h��5����1�.�w]�B��r٨�w�tWAx�vLu�����wN��8U+�Id��άZ6M����֜�a/(�:�D���زE��e�=۴��*^��)Q�it��2��4h��%E״�m��� )�F���^��t^����B��-\i���rн4�ޕ�uT�wb��T0c<�'[ϊw��#����Y)`�#�ô����l��e�N�7���?��ص�jՎE�_�1�1�A[���
 �v�EA�CN��"a��T G}��a������?{_���W#}2�
b��A�gr\�ʎd�G�^�=�(]=yRLT�RgW8- qD��2���]˥m�V|peK�?�&�]��H�C�e;�\�9�-�KX�2g]f�wN�T�L^G1]mҬ9V j�5�aW�'uv��a�2����p�[z:u̥�u�;3B)vE'�RQ�Vt˦��bpP����e�a�:Z]=���
?e�9�gw6B^�k��R;X�ʻ|8'ڸ�������e���7��}hj�(�4���+ܣ-Tq�}�{�y�n�.��͒��)+��l��e8.���m^2�5����ѫv]�3��l�MB*Oj�}��8����R�yv�]-Є�����q�*C�+�7�ww2�mP�Ț�+� ܼ0MJn�"�5��Q��3�c��Ȼ�F�T��
��/���Y�2��u�f�W��
��2t��.�:�\���ۚ���+,<�Ŗz�ÝjԘu�\#��޻������7��Kl=�������Q�"%�:j�ia��ͱ���3�7(���K�,��f�ؒn�T��gY�z�k����hA.� gUd���u+3���h[��&�h�paq�1ϧeӕy
s�oE�\t]��{d��솲�G:dJ��9�:��[V�Y���D:�R!�9yʵ�Ք[:�
Yq�E�<����;T\��3���Ь�]��p7ו7+��E�h�V�wx���돺�Aj_V�J�^V0sXdŠP����ِC��V��K��*��*��.�r*���g>Z�I�]�U��I�@�xŰȼ�!I�5 ��K#ZGi����1�+����U���Lر�$��򶻍�J��b�)ruV�>m@ŋFkF�;p4��y�j2�P9��0�372����z�R�#�8���8w25�B�8-�ܪc�VK�Q����Ԇ�hS�)V@(���M�z�ؠ˹{bV7�&Q̌�	��,E�)�:�g'�Rڳ���D��πM*O]�F��Mxc�t��`Q� �ʴޅtڶ�i�/lܱ̻\��1��Q�3;���N�)�1r5t�T����ԥN��to�a<�KFV,\r��Brm�ҠP�F�n����w�&��2��^��"j_`J�M������<� ���|��V�rP�e9�X��c5s�v7L�MT�7��sH{k��� �,
#.ٳ��×� 
#sH�R��z�mt�Le�]�Ha�%���:y�X���6�xqI�qu&T��V���V-w *�
�9�������5I�����Ժeݮ�N��V��R�9&�Wnn��B[����RL��0	��[�����T9�B��ɽ�o)�(f�D.��ڐұ2"�w>��īegt�q�Ywl��0�soPs��k9��0Zwh_G{*��~���ɲX��P����L_L���EmT�T��)}w���;�i�\��t��[%�w^RH�oִ	QqIoZ�s2�r�P�9��}L�
�W�I�-�ڛ��`:ʹ�9��r�َ�Q�n�iV�+6˵����-�ŷg�����m*�q�boc�.�u7�<���#6��L�{�������gmq2qB��u�$�
�����vaodM���u��˻)�[���'y.3a�
�:>�=ؒ"�h�t4K�7[�u}����Ǖ��6�s`,�ۜ�Ī��Z�z�%�ErgĴ�W�����eN��Sd�$(�3�{[��k����M��B���E�A�67��䛶r��i]K��u+X�RG�ւ.gKOe�i��u�cEIx-7��V�m��]���ں���iED����u���0R%Ǔ�hڳq�"���u���zv2���Eq-a�5� �}�d�#�a������D�l�3��xhni"�]��l�.��;� R.�@�kw;%$��^��d�݊�r���x�ѩ�M�YĨpMV����m2;.���>�2���̾�U#@�`��ct�	���]9�;�i�x�U2�kGF����Yߔa����cZt��x��.�������B41�Z&­�#6oD\�y�wL�-����鵉���]Ak*<��a]T��wX��6;S�� ��oR������jT�t5�؀;0rF� ��E��X[x(̠SK㵟p�U�[Kol�]6�Ӻ���b��dS��R�tuT�}f��P���4�%��1�5��5�̸���$ٗխM{4�v����Ĩ��'��;��#�����-��Sv�ҧ&a����I*���K>�(�5�έUk���ƌ��M����f|͘��RG�־��0�$��V+VgoM*�܇>!�c
�ѧy��q�l9C$BV�%�^��%��_`��A.�����R"��`�,B�����i��O�܆W��VZM]��wR�F��������8��v�fՃ�H��'�՛�����(>��ڭ�]����R춢�8xê��-�\��-<�����u��=ָ�.���yN(TP�Wim ����	4�˺j�BzByb��u��.�I�s�����ͦ�b��]��;[��}��\��c��kGo'����ky���al�ͭ�B9n����=�싁��*��0r����O!�iP&�:�y{�X�*�a��þ�g��Dl�uc9��s�	uJ��ʝٗ�q�V�O���o/�ZwMQ�w��A�<�+�]����VX���Q�E󽇾
V��Š�é��u�'�^ྥ]����[ѣWV5���XZYZ�e�G0�ͼLu5ہ�-Ôp;��;�/��6��ϣ�[wz�ҳ�G#�d�%jb�T�S��%���`e�l���^�/,�<�07�OU���S���ï���h�X���#��-uĪ�t;��u�<7F��}D��ۀ���,n@a=���R>�͜�]�t�i4Ώ���ӵ�M�0}f�CfZE�Ѯ�U-t.�\�깃:��XMu2�U���Y!`�&��hݱKh�R������\����3Ne��t=�`�9�=I�����fN���M�ga5�qf���i���)��
n5C����\1>u�)g^�b��W1R.�l"D�I�1D� ��H]o���srT��\Vng��lOX�a�B�aU��z��M�8@-��*S�t���P`�(Y�e�Xk487�ذ�Q3o�K�:��1�|����b�t+�J��nm���b1)�ԗP�}�P��WN�Duϫo�2�*������Hm����n';;"��v�f8�O�:�-N����(v�,��S�d׎#�c8��ԃ�p.�oum��E �q�Q�rs'\�Y3��Qך�o�l��iP����+0�9q%�b�u�J�[��SlQͫ���wgpT;�w:_+9\.��0�� �
��K$��Tn��ō�t���	���3*K�\!�שdɒ��+-�*=ۊƩW1wS�l��	��#:�oL��Y�-���ע=����4N�Xc!~�9k�9K-JPv8:�zP���JZё��WJT7�ؽM�P��Ŧ�L��&�]��|;�̪[����5��� ���D�jr���5�}��m�WS!|�9#ے%xW/�O@��˵x��� PvmQ�:'h���(q�4W2�ͽN�b��r�bem�Yb0�d��m�K�@;���=�c�z�ܐ�Y�=T1�)�8eL.�g*J{�\��C(�|^A�ʉ����|v�v̡ǈ�Fj��e��(|:*n��@�,ܢ٬w�q}����e�e�'��Zvx�ҋn��#S�P�{�d#t�Wm�\�����ǲ@w�PP\����L�AeBK����v��s�9�7���яI�H�Uru�7�-C�g�9Rw5E%A\��aM,�Ǵ��ǐ�eZR�0��!wI�%���6�qnq�̚�Ҽ���m�楕˩ۆd�l�sL�ۤ38��sN�wS7�E��,k�,��N�r�t�=4Ur�":*㽢���+vӺ,Nw|��ymMr���S���{�a�b�]�X;1�k�`*�<��̛ r.�t�����d6��0\�k)Mټ+G3�*f!δ��)$�]�[%�aĘn�ǫ�-,����K,���^�ڼ-��([C`�Gsx;��ES���b�lJ�E�y�%F5P�/�m���j��6��:r�����;4�j;���5� �G��XѺ>뷭3�(��Nbai�s�gn*�#����P���,DI4�7�bj�J�t�*9-_*"%ӹ#�,�^�d�wmK�E�tt��v*���V��}�1����,J�s/�^�vGH�5�I'����h�GGL����a�GQ]`U0���[�T&53�cue���y@)ܤ�;x�
]lj��6���gG���:�q���ׄ���N��e��YGze���Nl�������}��1^v1�1w����H*,�W��VM���t%)���l�R�GLh�
n��l
��]~���,���7�8�-�sH�9iGMo6��}�X\�W��3BF�s��x��]�Y���zVǮl1�C��gd�۵�a�R���9�;ʴ��Ӳ��*|B��7��.�������%�J�ɽ#)
��B'͎-(4��gb���zv̮����e+%fQ���+i�v�_��f=�*ld�����n!V�2�pHFź+�.r5I
;2�ۜ��\5r�+��V�-�n�$���欮ų]ސx�sY�(sX��)i�[�-�(<�vDF4�W$,S�:������!Y��b�{����i�{F��ʗ��n����0ϣ֠��1/����λ��<��/��(V�Te�be�#�F�(� �P�*w���wï���
0��<��+y�E���>��i}W��u/�l��|��}��U{ w۱��l�Ue����gP�f��#oH3�S���Y�f�r[�@�Պ�ML��ֹ��{��>�u4�m��/��5�tQ��љ/B܊D�o.�>���%�Rqvi2�ib�w���+%��.��2]��X�eqY�r5nC�5��L�,��7`�le�[��>8*��U���Z���Fq��n.�Y�{�Z/��G@�d]l[�rjS1�#!��[�'h� I��%Ȃ��	�ٝw��VP��r��)KH�m:˦�z&�>����S�6�Ȗl8"� =sa���'�>	�N.�gu̬ΙMd�"�fSŷv�7���/;��#t+;���[�wJ�Ւ����3�7�]�:���k38���ް�@���䓡rS�⊨�\yt���{n�ko+.W@�[h�4�Q�i;�mq�d���غ��t�A�CU��G��Vi�o���]"�n�/;)�QE)pv.1�/���Jѻ��yD݉����e!���,��[X�n�l*֚RC�w;7�v�$1r�����j���L��0%�.��,Z4�&)}z�m����3ܜ�6f������a��\�J� �`B�7"Ң���  lV_o+Q9�Z�#��ۼ݇����άT|	����C���
v�F^;Z�Ylӭt]�YȗMM]e�"��Qw(�f���
�:���ڻʽ�9` �=n�e�W���KV�k���УW���\TTݘ�9y�W=W�FL�uy��]�U�t'X����0^�3h΅Z��w��g=����Xց�3��9����'/*r&;{�z��T(�K��W9]I�g�̜��G��P�i��[5>u�����i����6�i.[-�u��jy�)cI�L�S5�h�&:k(�z{x9n�y��=[V
�-���݈U�{]ܴ%�[N�u;�ϏY�c�ư<���WF�js�Ys���;�~��?d��"��p;��0}w�o��	FDL���r��(� $�ͨ�?�����u�m�7��B�.����Υ�##��[1�ax1�q��x8��Ϡb��dʂ��neY,ty�ԝt2���;M��j� 4o�\�M���C؃�Y�U�7+�U��9%ĵ�y)S�HvG*�7vY��H۾XH���r�s��A�֒���/�S6������U�	��Aze�Y��,�������a�yO;�V��i�5�������5A��r��G��Q�>�fl��2l?��V���XXy&��g��:��Ͳ��A����n0Nh��#k�)bC�����6R<o��5� u��$��	4���X��(R�Ω���o��nY���L�q*�@�{�2�E��M`r�!f@PÖ�HN�oɇb����}|�}Э9�^�sR�sd�������y���;q*�Ø8;���q���2�Y��u3�ѣD��7O
�.;rJk68J�yՏ��ۏ3j:��*|��0�Yu�>�v���,e5J�ޥ�B�����$�����������e<�<N�GE,��R�Ӳ�o-��D�J�m"�]�MR��]G�Srt�� �^v��G\�՛�ڢ�Z���kR�D[ib-eZ��c��1�Z�l�,m����+��+%VVF[
��+DИ�,��)SL*,�`�+��Ud>fe�*M�E5��(VN��HUZ�Rc*	�����U@XT��!U�$U �RET�)�"�Y؅B,#��E�� ,�c
�"������V��X#REF� �4��$���$�֢�E�R�X��BV
[b���)#�Y"�P+���O�{����s�}�5���|<^^���
��;�(#�^����*�ٗ�n43����ͳ���N0����
�}R��,>��W����
t�r���l�����{��F0��(�r��+��7P���#$g�W�T��h��G�]�ꖽS�ˍ��T�r��i�+��>�o�Vώ"D=G�1�M�M�����g'�X�����B��1�g#L��rǮU�[��U\V��c"�4L��P�W::/C�"v��r�V,
���uG8�������g:)��@m��3�Ns�Պ�o	w\��mB�C��d�Jp.��l�y
���������z�WӪ���*��9���'n��$g�{Ѱ�����N�K�B�mI�l�l7BnʱX��箞���Y����C6�߹����YU����	V%қ�-����%�x���d���;��Z"~��`)�@f�e��%ղ�*���a�v/]�q\�Q��)����
��$}[��
�9���ݻ���ii��\x�(5^@~����QnG+F�u�t����ݧsWH�E[}�A�����8�!�[ٮ����O�;�*��6�ȷ�.����x������m�Λ6�G4�X͉.#�N�3���-ԪX�)� �0Z}ו����.z��ܭ�>W�P�J�),B�7��	Z����L�v��8�u�k_\�oC��r1{��+.��O���ej���Q�=w��]�Z��N�J䄪Q �KCjyЖ�Ե�����no(3G�m*���z���I	@����޺�(��4�uk�K�e����Yۦ�+�<=��!8�H�k��9�[ֵ�c���W2D.gR9̻	�}/��sb�(��}�B�s������g]>;V�����')�ޮ��je�e��:ʷ���pJ�J�B�+3UYy#O���ݠ-C~���R����6�_66�WG�n1�{X��ƍ��ɝ�n�Aխ��L����͊o\��z4YL��n�g��Mr!@b���ӳ�U��w������6@ю�������4t�m��Rt2�A�"t�}g9�c�1�v)��U48*���M�E�v��*$Ä��b�+��oy�Qv�Q����؃�aWc�yPKx�{&R���[�'���>�c��B��k���./0�18.�N�F�����hօ���2��/���V8�-��f�ב",���e��h1Bh�b-�b�U���.!�*��e�vo�OE�2���5�T�.�Ae{E(�Q���4��β��)�[.e��ŭlD�j^���$e�opW	ikI�x*"ce΅�Ӎ�\y�:s�6���\2�B^�{3o9d	�8�|�u[�:���	j;����0���g�Z3ˮ;'�v�)�w/�!�6�5E�oEp펃�d!�mg\��pws+�Wݐ��g\ib�o�%u�Q%Nv�עM��v�%5�EL�;�z���CZ&V������;�,�MP8�gN��#���H�uk���L�Z��r|�r{
�IT�Hr�!­�̇�fz8f'T�]��-�+������92����YP;*�&��1Y���ƤE�q!�j�t��4`�8踫M=��0/�SP$q#T's�;��΍��_H�.�v���;�nHڌ��^)�-˦O�ұ=�1�q$kJ��Ӫ)wZ��W��)@:3w�$�_e��C,�r��g%Z�*WQ�L�bwP�W��:�]���k\^9�����^ㇲ����]B�ޭqd]�@![�f�[/Sp�����6��м�F�Do-1}Q9;a+����m�t��;Tň�t,R�8ʜ�y\_.��y{��{�u=uD2��J_F�&g�3�N����t]k�z��%��;�G�6u�DvR������Ε���7���{s/n>�m;�Z�PO���y{�Y�mmVj��傞m�;��ks��䢹��f���%��������a�`煮m�҅uਏ�c�Z쯕"�l�;+^��{�T&2����\e��d�K���=�qj�Ϩ	�#�ܪؒ�=���P��M(!Jr�l(�B�o��P�2Tc�]� *؞��0�\���1�1+�ꀟt�
::2��<:mʾ�79��"�ܶrk6�wX��Cw=��F�S�EPQ�<�#𣰰Z9��s�77g�cb�N���$���	�����>��C�EPZ},���3�����GFƹ0�Vvq�v�3��lj������T�>���F��×T��b����f�ԧT�sPFda�1�軕_�Й� �p�h��kHY����mz�h��߂�/kZ�����l�L@�':)żN�H�C����dQ�t	��9�1�V��I��X:w`�F�T�t�������E�{�����r.(c�t�FܺsUٕ!S]��f"Z���ߐ²�x��R��:t���m�	���n��OL���̜m���Y��U���X��wj���ɓ�_b�n���BknY�����M��!7��ƕ:�m�#�ͻu6�t}�u>�������X]�qQ�ݫ���w� y^��c߁��:�<�/i��g���(��#!��"�L���B��b�ѠC��;��wR����L�1�O���Q��F
}X�Rs��D�/g�ڦ!�2voI꒍_������mhy�]fU_��Ú�+�*�YI�D�W�e��T����C��w{V��!�UѺV��s�<���)[���S�mX�=suʯz#��T7~�_N4Eg�Ub�FF\��y�H~��cc����O��� Dd_M>�2fb�P`p��������=z_j[����s�jn6)����͝ƅ)�Xe��6�R%F�U
v!G\�䌓ӱ�NeJ*����m�*�,c��<��[2f���Х�\{Us�o�	qV�v<.�P̐wt"2�f����l���D�c+*�J�S�F�F9B6ds��^��� =I��ƺ�F��坙���{Cv�}���Е��R]�d�@�pjq����z�xS6\}�3j�N���;��\��u�tԂ�kz�1/���;pq[�y4�7�h��5f��u�}ƸQ��/����JG..�v	ۣ��܇���3�[�q	��b\vMA�U")`�< )�=	c�|m�3������YŎ[��<"×rr��]�ʾ�b�ܟ[d�Zt$)Q6:��Td���@�b=�3�\�܅�Ft��!\��.9�`��d��	b��s��հ&�2�jFC�	��&+��Qz%�W���	ת����L8�+$�gs��6j���>�>�h��"��
�27>�v�Q�n\�, �\.�kR�#?r���AunM^ӃR}�P$![���s`���Uph׻4n����2�<5�(x_E]Zh~V)����%�d��<����a��:0ea>�Y��X�8N
����+gc ��'�k�z�3�ö��R5|]*�Ϙ���*�3���8�1�
T1W[}Y�;�>�B���W#V���u^K��+YpY���/ZY�\(��S�0MD\�.�!p4:�L򞶏E���+r��*�}�y;��!+�(�]�3�v�5̩�GF-)+mx��c�m��Ti��H?����v�ٛV�����s�$W@9�L��I����g%G��qh�&�1�Z�롡M�QL�����.�m-��S7����n���;�s�t*���<���F��8+n�V=�º����D����9ԕԮC�龳Vb�vH4T��*>��j����K��f�K��Q�i�yKd��z�y�Dw6V��kE�@`7[K��V��
z��aP�D��kZ<c���r�Tު�!��	g�N���A�b=���m�6��j^[�����8櫩ěG��l�
S�뛱�Bu�*/��ʕbf�h���W��4�;�2 B��\j���p(l�tYtܫ��7�8)���$�^c���J�|�*��KP�C�	�=�5ҳQ|Vu��~b�Y��1ߏ��"��ageٜ���}�j=g����:TH��Mh^��{�⾇�ϼh.���[����Żfcv[t�L���+d��	�U����
�l�8�B��3mz���:�?e�Y*���P�TFy*�
�F��m*K��e�?>	|�k0�y�*ݵuP V"��^8�=�9N���Z����%vV�$�iq� ���d������;����ݙ��h���7�J�2�:��6t�>��S;�T���hYv����w4wR�0^�r�̋��,L��z�(5,�6ez�]Ss�{HB $�Ș .�ګ���Ȝӏ�n_h�W�D4!�:��^4�g��U�6��9��j�LW�Q��\.�����H%�:��b���:�X37-��PӴ�49L�QU��o;i��v;�ޞ�vj��\zT�+^������
����<-t܅������:do�޽�N������N��h�T*#��Vч3��^r���_t�0w<cc]�\��g :t��d�K���򮉠G���\�k�����{�1��bv-�R�l(���;
�Qn{��dQU�$.�	�ޮ�㜥4.��(~�("*�P�����jxtە}@m{s#[�T�9�iB�X�]�=c#_��1
,F̨s!G�Ǚ��*�����	N�S�i��!�VI'�''�,�&:>���;�>�.8��>| +�m�=��{����-#,���:�f��D�lT;,�9Ð�fj������f����U�.ա������_*�����kq��r�d���ac#��Z�4�/)��"n�rg��غ��O(�x]gh|v������e��.���?[.:����u�
�'���ӱ�\`#b�qv]AԦ- �5
�-�vd���:���Rɪr����#�3�<�
DM����}8y�&�Xޜw���o/���e�)q^��=`'~$	p��uV �U�F}�&30w�����Jb�D�l[��ZDQ�78�(9�&[�'s��r.'��C�]Ԣ��X�u��U4��dl`�$ԑO>9�Ҟ�Y�j���� ���
+�9OSB���1�[�V��#j�xPQ@FFCv	�E�������!�us }7vz�ƅW�ʗޛ�Ŀs�S�s�J�?G�/�`��U�'?�c��fDv����Nk��?��e��\�l!���ߋ���P��ˬ���\D�َ;^[Ngt�jz�2����U�{�iܷ�K!X�Y�Wu���Mt�o��ۊ�e3�{{lR?
�Z���r�͟2�Kͱ��WA��?��	��G��q�g�*��ٻ��5�S��j�j#�:ƯCb�N���ȧ��>��tm�ҦV^T�`�Kr���0�"��g0�����zt���@Ӥh����+�1��Ggq��=;U���{r�;b=Ӹg*��F�;Vz�#��M�6�J��un�vbisd�7���BS��]jK6���#B쏵��0���Q���!W�-a���T�@mH� ���ފ8�L���Σ�wsɉ��fVX�墥ZT�3zJͬ)	��	�9ٸ/�]������۹{�]�;J��in��Y��>Uu��rً	B�r�,pd��Ih�!���d=3ڥZ�h�&K�B޵K���f�.�f�d32E�&�����K�vAr�9���^�c �\�}}oCMc�ܡtK+MfN#k�n��\&�5�t��w��ק.m��w
�_���#R�o����SiX��@Ȼh�\����o�`�L�mĒ���C� U�L�L&&rWK�5>��J�}�3��|Mj�]׷�vdP�pċlbp�%��k���.ҽ+
3z�Ȭ�c�e����R {Z�oA\���:3w�/'���-���)��+i��_�B��#!؁�f��(vP>a��=���0����P_�i���=S;��ɽm��s��d�P�h	*뻯�+l9ٛ�~�}���� @x~�!�6ໞ���yz�4��?š�0k������M�2����ep��v�unR\:.�:OU�<��:wQa���D~(M�j��M������s#B�RR��%ԃt8�K�1e���7�z����#����}}Y
�ҳ('( ���,ww)5��7�pjȪ۝�ٯ��)+��*���hq�V�vXVx��We�k�yח�*���nd�ȵ�p{àd8�cWk3/��4�'�,2�}˱����v��@:��\���4�3�s��%�6��cI�C{��������3ͮ���$�����Zy,\�j�ۼ�o)�7_�p�� *'m�]���y��?����T&	���ժ��|ᧃ�y*ӑ삃��;Ks7�J�+P����m�goj�<��%�"v���]�w�L4*s���w��f92�S-���4�X�Q_<M�P���fvZ�/�B:�L�74Ռ3����Ԩ,yM.
�n��EZ�λA��� �Ū��hP��^�(�`�sl�x�ᗘ\�.U�}:n��E�����As�L�S0��g2�Wsx.��)f��r賻{���eԂ���cqq��-,Φ����0�ɗ�����T�`T<edY�LJ�"�aE��H����YH�"��((��e@R,��`���Ђ�)b��VAH)
�I��ȳ�, �YJ�
�ëdY �X�EXA`�A@$)�+-��EUa$Y"�`#
��A���1�((��L�$r��YD��P��AB((���EX�X#�VhaX,X*�,���UU��*& Ud�
ì��A��P�Ud,���AQ�E���CV@R(�XvMc���=F`N�V.!���q��������ODI#ݘj�n��g|���A��X��rN��G��+���=��#�y���#��@� KL�vzEt�5T|����h9�~�u�|�����x��.�>=��q�#����(���d�����\l꽉u��I����j�}v�GoI���2���=k��rs�#}���=��g���d����5�|�S�	:Q1��]V�*H"=���P�Y�<.Z��C�y��O9æ��pPyM�
)ut2�߸��¹q�5%R"������U���\����������SJ_��p������W@����˭�����+���0�@�����ݝ�x�>�B@��Ll׍�E؇Mȱ�h�#:�a2���7q�2��S+vu�F�ڡ��𳂍֮��W�*!Ӟ|#���|焜���eje�,�S�T��l�]�*P�������oKE��D���s�h�E���Q�m�Y��hDh�S1iP<��&��iA�<B�".�񛀇����yW����g,t-�lo1w�@2:�*2b��F�c�N�P�;(�j�0�U}|qz�����4̫������gr��LD�<Ε�K"�$���L�+8i	WK:��;��Y�gfcjLΛ��Ψ�����������t��
}��'j)P��C�_,v{�,��_���lWR<<*8ދVP1���A��TxШ�^��{{GC�7jB��a0}�,�:����y���T[A|��}v��6�l�t�R���|�lb��çCj��j(M�r����94:�|g���z-M��Jxo�������9�[���@�Pu�tIR}R*��nk ���]��v���Ѹ�|u�ze{��(^��O-��J��U��R��CC�W�}g��o�����П9���2q:Y�p:�+̌j�7K%�:2�\��׸W�0l[��22�,w� ����V�cE��׻�ѳ9���C��sA�W#���R��
�<��s���Q��xS^�]{MH�2���a�dl0�lʌj����f�kN��`蘗��Y0^�¸��Q�b��}s��7P��`�;w�Jo0����7���G/��]��P�\ ���"V�a���|O���5!g1Q��4[�p� Њ�3,��[��2:��#�gb�l�}"��W;M:�uzq��������cF�&�X�Zn-�-a�V�����M�@��n���	
@�ƺVj ��{"�[�$�dԱQ]Ap�U�oZ
�E�Q��S�|ӫzTH��Bk�ixR�p^��x�����̚T-ק��[H��`G�UZ3��N"8@j'�"��0G��ク��v�\Cq�Wx[�~䈫�]5�+����**�JtB^� �Mp�]�F�sɩ޶��4
ca������d��C�]d�6����3�VD��[����e��{�GF�":��4��4�ڱ�W}+�����u5A�z��$�=��R}�*�S�T�5�^Q�C�&�dUpͲ�b�*�z�;����I�^��$<w;{S>�SJ �myT��xNK�/���N��n�U)SO}'u�kB�u���b!��{�3�J�����G��R��
�#�Is�5A>��C��t;�[l�e�P�~	q�=�WD׈�7A��zEf9��A�E�͡9��u4v
�e�#�,i0�m^3a��u�r�*B���֜��} ݃���/
UE]DS;���Vcaf�fUH�sr��l�2U��)q޳�:m���<{O$�jp�X�73s�S���ڟ}2�P���'!G)pʎ>��i�C��	�<j�lHOG&y�z���n��C�>�B��\tt<Z��*���.�L��\}+���k����z�C�xO�:�:+�ٕd(��̃�vUO�w�Y�]�#�:m�ȸ�n*"Ţ��h����>�*�\������ewc�;�����i3\4f�ô�p<�$"O�z(o�b�L9p.��X�tI���C�7Ò����+נ`��scU���>����� �p]Y��\��^�Χѿ7=�_�]�����0GL�x>����gÇ��%(1ʲ*�N:���\���W�S"���v�5�L�>�78�(>Ω2�'s�P�Y@]+�Cϯ޽�6Q�U������Eu�H������O+�Y����wK��[�o{XKC{���n5|!ƞѮ�_@�cj{���C5Y���tsI[�5+����Uޫ-L�wt�E7+��w-��C)��k��tZ]x7Z�W�f�I�=��-OF�Y���5������\(!D	b�Wb24�ߎΧ�yU��`��y���+xb�
:3N]Z�UՕ�)�"?���}ʕV�d�/��)Ϲ�%e�x�d��C��
�xA�gq��v��~`ec�VS�Gs��;j[�!�aco`�%zF`��8�#e�1낟&J�C��&9N����Hq^���U�ho����t5��{O�<5(��6��Z؃�)*B�f�#�d\j��l��ȇxjǫ����V����M�|��9|	��R��Bt
�44�Gg���dj[�@�nR��D������ؚG�5�1Dmz(ّ�l(>�AE�Nx9��2r��o��o!R�����;$�u���JW:���8-�J��ګ����Z5���l�W\=�:����B�J&8�eeU�Pj|�F9B7fB�_��c{��:��t��U'9HQ�q�g-߸��¿K�ɨ)T�������i���͖�g�D\�'�h�4��9�ꮁu`��wL�O��r?����y3j�O��iΧ0<#��p^Ν��V��s���m�W��H)j�m2çy79�7��0��5��"�%o�J�������0^�૓*LO�_v'�웖���e��x�
��i�f�����P2Xzh�z)w,��j{�Zď��k�Jq�y��_.�=z�y��:�f��n�|�
�T�Ga�Cf-H�͌��ϣ����MH����LP6ʋ%�SD����b��:�����U�i�R���E�������]>J{��Ө�����Qy�#]w���t��#W";�T��YeL\/k�7԰P{�Eӗ�<|�	9V��c��v%M;(p^ۮ�t kg<���N�N�]҄c%T�0�Y�v���hĥ��邥R<:*D���P��j���k�Z;n�hńTS���YRj�7ɚ��h�*4�Q8�ӕ�8�/��[B�Hգ�� �eQET8�&�qx��^��#��tPF/x����ʭ*��	��y��Iٝ#'�RG��X�W��f
����/�Q�W��YE�t�!��[��k!U��!�F�F�C�筋�0�ןk�no�6\\Nub��]�`Z��*�EJ��r5[Cۯ����v���ؙ~�I������k|��0���:6�t��V D!n�� �6-�����P]��K��G����i�LCkϭ�4fu.Y����o���C}�>����G\ѓ�ݛ�R�rp�iA|P�+�^�{(>R�����t�W�4Gp���$te*�؜�^��nu���=��9\ġ�:�"��deE�|'�
�B\�>�[^y,�pX8L�B�u]e^>������ρ���$^��^[=ʭ�M���:ٕ,�:gt%��,|��횖�TMm8��%�F��^��6�:0�nU�p{�9[H�VѸ뷚y�R*J����Tߓ�"�<'�Dk���@������ش�V�5\�yE�̒���X�@�
	�>�'$GB�ܨMh��3��`�m�F��:�AJ���j����a�x�pfP��kə��z&���M����L�_u��i��H�Ou�u>)կ	���s!w-��+y���+p$�n�C�p�������̯Qt
"�no{HB�%VD�s׫�.��&�_�����R����դY�b�z�w}+�/��=Bic�2W�;�6���q�h�7&Mĭ�]C��]'[ЎX�㧊_E�/;��鶫�6��&B�v���v����k���l���x��� ȷ���[
M:\���[ۡ����� �-��g��2�'d̩GDӷ��Q\�rcL��JCu�����6��P���.��m�Ƀ�q�c���G2�ɢ���Lw��Ϩ}�a��C���=�/����#��f}H��k�u�� �lCo�}[���g�Y��q��q�T����c��)*pl��x��𐣶7"/w�]>Dev.q	�R�.�ȟdtf��M���.!�됖֙�tJ���.�.���'/�b�2}Be�B�5�|眸6Tq��~�v+d��4�M����j�B�
�ix��`;F�Ҫ<k��ѡ�z��C�K�@l�]�Oz��ƒS�"��/��3�X�F����B4��C"�(�d�GaKLl�D���K{7��d�mXnFG��LlmM1=���\t�[�ʋ���3�DL�|�����x���qr��v����B�::�ӱ]0���T)0�f,3�fnSC��޺ ������xJ��@�בؙ� �p��G~�ֱ��0����yޘ ���!G2��]B}$��7�|y�(*:�����I�3���9�Gp�ͧIW5n˘����k��w�l.zb̑��!2m��Ꜣgn.[W�d����X��&j�ή���ٖ�0tC���x�7T�Ίqow�D�Pຫ�*�w7dS�{��QQ�q!�5��`5
j�"�����AAΩ2�'s��ɾS�cug$33�y싊J�Ӭ����U�
��Y!	*y�A���Ne!+�Qr�h�P�={�f���""��j�U�5����
A<((�>ȡwW�r��!�OJ7��5����P�V*�n*��pL��4�+�Br��Q��
X�ۼj�NW](��':6�G�%�r�u�h���U�o��a�J��e�f]�!|����ckxW��Z��X�8=B�W	XlV3��X:3]�+�w,��s29�1��X�J3f)���.Eԅ@��Gȸ�+Cg̺Ȯ�Q�X|k�f�]�sTM��*
�i�H����ht���}s�+�@i�Gh�].����&��C�yO��>W������Q傖Jנ��_
)*������ F�]w�����y�(\SI���oq3���,��m�:h+޽�b��	�U�̳�t�&��x�ߌ5��\}��{Gr�q��d����K���Mo �_f��\�T��+��w7��љiD���N'sT�p:[�O)��c L�
����C�
�Y8�c�r��]k��S��vW�۩(_&�p篭Ō�
�y��t�[�}���P��|4���4r��ב��F�	?T�E*��\�ɿ�(���3�������\vMAJ�BY�U�y��\��k'NÏ��l�Vh�H��u�A_��Go~9�h|�����$Ͻm^c�*4�x V�>���%��^�� �S���'\Ŭ=u<�'�j��.�����A�D�ԠNJ2��~^k���ְ�>���`ȓ�^T��~�S���Rh�9�}ΆT���~�7��/Ƹ�,l��mQ���|�:�|���t�]���%3	H�չ5ciA��Vy
���%����帘��0��`����J�h~4�����uJ: 5��
}��'>�ɗc�=�_���8C��&��fI��R⁗���O�ז�\`���F ��d|i��J>�F���J���*��	,�>
��ㆭ�6� �,䆻8v�nl�]��.j��S���siV���BN�A�zVRD��%���Ѣ���O�޴xE��ȭ�9���7� �]���뎯,�%��V���x�Qi��[�
�hQ���+�Z���Ԡ�|�^�ɼ��/Skⷼ#������]�����j�@5e�p^��\O[h�b-�KQ��#���T�/�x���qnQ�S:��q�U�X���l�]��HQ9]բ�Vt�eq��s}&�mJ��X1�U�\q���ebcSB�_��A;��۱C
NL��^6#3�ӭ���*�,B��w	����nы5=5)*a{S5>v�c�c�`
��ܴXW��8����z�N1�y����s\Y��S��ho�P&rU`��@ޝJ;�2���ܣa�^�Ƥ��a�,��N>��z'mjCfe.���.ʙjL��C&�Γ{�/�nX�vnk�t���Y�i�%}gJ.��C]՘��n��Z�����0��39��溱�L�3�'V%�k��,�,��.A|(�e�N�����ӓh����ߖ��9u$.��r����
��H��e�J	��w�2�M������3�0��\���2�	��&{3k6����\'Bj��8������ȑ?��u�+���
�"�sj��g+�P�}��[t��Z���X\�y%P5����L�BNCf����W=�4����A�n�G]Y��i־�n]��+�E��'M��5(�I	QH��{g��P.Tq�a�t]�zHͅ*��Մ�7� k���.x;TE�s`�D3UhV���}�d�ɪe,f����m�;-\�e�����2���\ӡ��7B�h�)d�;�.��F�r�3�X���S�J5����a���s6^9[�:�S���3�����;�x��{&�-��o�;�Ŵyl�;���q�̣��a ���p3�u$��{�K	V�+&5xj;�/��9wn^ڨ�w9ԩ4	�qU)*��9�+��AN�%��2���a�L�ԭ���
�£�+�P�s�]9t�����3 �dB7n(y��b�qM4�ΚNr �������󣗽���n����eg�U�Đf�ۍj7���u�*���i��lp��Y#�j�T����U�v�E޾'7/��:�5�siDm�*�ի%8��V�aH����x�a��e�9��s��Z�]_e���'�q������H�A@�
��,R(i*����"�I1��X� � �@Y*�1���dAk$+,*Ri�A�
H�H@]!& )b�+	R
@8�!����Iz�%d�� �%d��� X�J�0��
Ԓj�4�H* :�d��R�E*R>���럞ѻ��e�|�z��uv�;:��+��}�t-�����ΞUԝ�_�a���^*���<eb俫�s&�6����j+���:(]�)�0VS�U�g�D� ^�"��s�6ɭ���觫���aB����.O��57M��[�����p*��c!�о�=��H��0�:�y:خ�d����T�	�u[�������S0��$�ol^O@�6���b��l���_<�K8�EX��T�㟙��O��:�7��<��o�Ϲ�Agʒ�<�b)��	���Y:噻6��Xm�@�*C�O7VL@QN3��`m� ���9̝&�=s����!�
�ɭ�O��ި�G�1P\'����(��|���|��P9h��YR�Z�4��B�S��I�gS��t�0��;k���C�l�Ì1��x���P�����<Ld��s��$���&���P��Ů���G�{Ʒ ��>aY8{Tr�Y�MsX��X�)6�8�=�ϩ
��~��3i����t��TY�[�4�tz`���@��>��"�U=I���-��m��0���9�C�:g��b�����
��lěB�;�墁Xz¦�H�<d��iѫ (��k9�H)4���Ԟ2�HVx�0�{�@��_8<��K�Nub�.�"t��z��oF�ֽox{B��vs��l<Ն$�t�i ���t���S�)1'�T6��=d�6�f T�N�֦�*�q�л�p�P����Uw���@����� 1>d�P;�xt���'���;�Af�+�u�d>�AI�Pĝ+*�����*��M��1״P�8¢�FP����1��V������݉�F�vu_Mx��0��ɨ�@���D�(��1�RmՂsJX�]�h���v����r��{���M!C�с�#ը�*3��Ma�B`����9�d�RWO�8v-�ܻx�d�U��r�(�������Kq�}���'��'l*%C]}�Ӵ��;�ERWLw�Z&!Y�Ng0�o�L8°��6��q�-1UH=��I�1�k�,3�B���y�")�������|�D	�p* 1+4���>B���vʆ���i ���X�I�@��.�q
��d�~����8���I1
ɹ����P+�i@�+�%E�s/��g/�o�Ͼ�e��b��sv)���I�����/��q0ީ>N&3L����ĝ�LE �5ˌhT���&�L9�C�hx�H,�Y�X�(��^؃1�-������� P=0=P
�=� ׶z�֬;��T��k��l�Mمd�Ă�e���퓎n�ά4���'S�7����Y+欜����*M�*L�w�^�3�����_y���B��Y��:@�*Az/�|ϐ�<aQC�RcT�}�� �a�b�Ͱ�%N�(�ǉ�La����J�'z�I;B���N���xLxtxLz��J�K�#Wѹ�M8b;�x��U�:�I'��ǳ߰8ï�
�s|���퇬�1'�ـ��&!�+��Ă�YS'�S�i �C��b�&�c&>&'��&=n}��ۓ�^LL���ӟ%;��E��*s�`I��l/(�V���i��*<�'̚@Qv�Շ���{�ެ�2�@�t��}��'ɏ=�1�$���b)&���ϳ���˫κ�ߞ�yl�+��t&0�,1;���Ag-& (�xʇT�!�ް���2oT��� x��5a�Y�J��sZ��� xF �P�Q�\R�P噿|#~���s�y��$���Ws�>S���XbcY9�R�X�jʆ�H�HV::� x���ˌ��C����
�3�w�$�8��;E�<& ��%�{y7��ʦ���zb�zɌ��i<I]!�I�����:�V��Z�qR>�Y&�T�B��e�>a~�+�wC�|�0�6���+:a��6�!.�!��)O�"���B�d=]u�mWM':���8^Z�Oh���6���h��;�%�ם�J0h@:��m[׻=�k���S�7����x=#�h�$�D��0�}t�N�˖wn<�aE72d�7\/�� �9�9�����G�`~O�ΐ�1H>�{��t�a�>�d�t��+:�f�
�>���
ϙ.�V� m+�O�k�d���쓉�Ag�;����{��s�}��J�ud��NN���}��'O��v�YĜq�]�=C
;�C��VN��>�t��_P\@�*AO��1 ��XbIR|��Ivzɒ�7|ߟo�t��\���{�c	�'l�	��6��!��<dۧӯ��ěgG����$�;��L����aOh��*�<`}׾o��=��{��;��͜뒲��1��fR�����C��݇aw��,�
���W��L�xC�%zK����
�3�\���0�a�7�i�m �Zq��C}�u��S4s�\��}�O�%H)/>Ⱥa�֮݁�V|�Ì�1;ꁌ�8����	��ɮ�ɤ8�C��IX�I��y���q
��O�!�Aa�:�aSh'��}�U��󿺖$��c�� 	�|�(�0 �a��(��J�����bAu�Cެ���CΩ4°�Rh;�N�4���Βv�H)זN:`�B���z�@G��H��j�����}�k�y�J��kS�IR=�E�V�/�A��0��=Xm�@�+հ<�|�Y�Y18��:�I�;d�w��t�a��d�t��O��}oY���=��ɧ�N�8y̚H)=T�{Β�*j}��� i+�����=C�;��$�{�*CVu�E�aX,�*$��=�Qp<" ��E�HYY���tn��c�$�
�y�I�[��O~��Ѷ��i��V�P�܁������׶0��<��tö|��L��w����bbk�)1 ����qd�Z�ۚ�'年V]������=큱�B %I�+:��I�;�CI�
����H?Q@��;��H%v�}��H��J���`i�'��9q'Hy�N�z��P4ö�7�����[�}�]�G���b9Z3c�u��yo���z;]��[ԭ=	�?�G���;�l�����g�ip�O���"��o�i��w�g��y¡)�D�tr�m9X���(��㻺�J��#����j�}�ҖdM������\����*�����M%E!���=k�:5@��&0w̆ z�Ӻc>T�O- ��������*A�ϙ��x����s�$=�|�_y����3*�ֺ�F'�( Ǽb����q
����u�B�������餂�j�ɧ�Ne1%H)6��d�A��X|�T���c=f��m;9̝"�Xq�:�y�{���y϶[�M���n��xäY�
��Ci�I^�l�� (�P�cX'hW�h�s\��}a��i:�3�J���f) �NP�8���� "���(���ͻ�^��hS���&0�;����Θx�9��B��S������hc���X�I�=�� |�&!]uG�&�YQaS�'�C�Y<9t������1T���{�R����w���*(b.�8���*M!�Y=Of}���L9��t8�4�Y�}�`q�'�Qd��%`v��:.a�&3^���H�aѫgʒ�<�
�<:47�����L�L}�!���:��$�vaRvyN�Im�I�[ΐS��8��d$�6��Y�)
���y̝;d�T���f�+�&��(
Aas���i�3��3ϸk�*�H9d���U
���ְ�ϙ�1��E �ﯲOP���^�8�f�W|�!�J�:�'H
(|��O�
�l�9��>�ѡ�0��:���U�|�v����ScƐ1C��&3�Jɢ�U �)��Vm���SH�L�1�rͦ�:`򘇨TR<̓�T8�C��y&��V,�4�t:@�*N'2+=�!��_̥�M�2=�>�@ Dp���t� T;�hi �6�0�
��{�k%E�2TR(��q1�I�*哮�ϩ
æK�h�N&$�Rz�M%E��5��������l��C�m`�'=�$P;L�������Y̲c;T�&Ң�P�}>��m
�r��'5a�CI��2��(�>��� �� L�C��-��D�ջ:n��Or5�v��>���]	e��� ��:�&#6p�[N��$�OjZ���%�n�׽��򩪋�}|�b���+P��V�ճc����s�=��v�hڗ\��M%"�U�o�#��������NV;﷬��N��HT?�a�:��d�{̚f2W�Ne7��
AOw��:H<���
��)���Hg�,*)���a��!�1�0�Dy�Q񘼟�<��R��g� �0RU��2b�:�OL
�Ol�|ɼ�@�*°�F�f��i��Xj�M*�M�&�z�a����a�4�Ώ��i��Γ;�gw׻�w�\�����OP�
��2zʆ�hc���X��w�a��R?P��,����.0�
�@�^}����f}��+
ɟw�N�Y*,�'{�t���ɉ���ۤ�y�{��|�v�z�e�;���!Xt�{c�N&�k2z��v�c%`q�5nЩ����L9�@�+�|�+0󬆑H(m=���v�ǀ����o�3O~�6���ǽf|.<W��$�:Hj٧�1E+q ���aY9��
��c�N�M0�
�+�O{�Z����mYRs����x(�`y,�G�����v��8m1 ��x�7�������t�!�����a�E�{C<J�0�ۦ�1E<E%q�P�2���q��̓ά�XT��<"<�ޘo��#ۮ>Q�~Ĕ��Ԫ�Xs�I�>q���鯩
æm3c�C��i ���C�����|��'��i>LE �d�\E8�;J���P�u�&$�T�Xi�N2o�}��<�c��<w����&��t�ـi��*O�|�x�Qf���� (�d�t{��AI��w�d8ιHV�<�>�'����g�>q'IQ���k2�|B��7׽f��v�̖s�9w��*<υ@c8�+��&"�P�}��OP��eݛd�6�Ϯ�;J����ՓS���{H)>y�4�d��R�d>a_5�i�5×�.�;�ӭ���ߧ������x�\C��:��P2Z)6��˭Xa�Y�v��>gS�`t�0��:�����C��;��E:>�,4��T>gg�����L@\������^����)0ղ�Oq��.�H߆W�'��^��L �y���F�jK���ց�<��=Q"�m���g��\\�js����1WV���f+��a3��J!?��v3��Gp]���f����r���5���鋏0?� bzɬ�!�l1��+'ʍ�|��ްU �-�I�q�׹}HVΎ�æf�ߔ��>B�.}�{�� } ��ou��5c�V�|H;�T�9�g��1�^�9��3�Y1�Qa�*c7f�m
����E���MM�)�*,�tj�H
/���aR
M!��'��Q�1�u=Lt|.>���jJ%���{�Ĝ��ͤ�ĝ���Ă��_C|��� �C�s�퇚�ĝ��I��4n�E �}E&$�
���e��Nj�i�uf�*T��O�e=��+�������� D��$ۉ���'l����SL>a^2w�k�w,�%zN�̇��H):7�$�YP>K�B��B�2m1 ��h��q�E#�����_g5��o�o<����o��|§hx�uzH6����2q�@Ĩh��&�����ݪ(z��`h�޴LB����a�P4Ì+�d�6�Y��4����t�	���������#��<�W��HV�tSL<g:5LgL6���T\`VOP���4�ud��dY�m� i�ˤ�B���1;��%E��T�:�y�T+&���_Q@����Vu���������J9{77Z> t�%E���M (���S
LN���'l��+Ѫ0�T�N&3ά��z�N��"�X뙦�*A��'I�r���&�6�����,��~}F��m��As�@ Dx�р;IRb:<��l���X;��J��9f�*�ZVOH,��N�8��=�Xi��+�O<�$x�n3�}��������x5�eo[*n��;o��t��9�05�!Xx��oy��R
�N3�4��TP�y�&�z¦����Βv��TY�ĩ�)+��&0�5f"��+�N�X`{ 	�}����`̧�8K���òo��Xv³�Xz������ *�=�$�g{�����B�پgl�v��|���AgL=LCHW��$Jʟ"�Ct+,��g߿Q��h�6���|@'��ho3�"R�������p1�9"aۢ�>�UΡ��-�7A1�4[[���u"�vW.���v�7�/�TO�'W_M�ب�փ}	�yW:`+l�UU{Ԏ����� {��T���2W��0N���vOκ�Xi�Mu����Xv��E�흦 |��%G�s�O�:@Qv�Շ�����ެ�2�@���L<a���6��큌�&8��1�n�������1���X��v�`h��݆'gT���>z�0�@QdזbIRz�yH?Y�&�O�̜a��Xvs��:��� ���@Q�dT��jM5t����HR�4�i�'Nwf�1��+�4���Ag�8j�k&�Au�$ڲ��|�+�γH%`uˌ��C�xL����s����lLwT�M�v�P;X&�ba�<��|���`t��i5OƹQ�ѡǯ�\hvEt/ �����=�6�������r�z�д�ip��*�Uxp�^�*k�f:�1J�;�qK-�ܸ[>��&:;:��J���O3i7!Gֽ���'[�q�Έ���&ţ��'ہ�"�p��K��B����^�����}*�: �AF�nxj��w*:��;gDϭ`�9�YѬ�J\���!����Js��9�{^����L@�9�.L���g�Ԫ��!y
6.d���XC�
�G�*+m*���LL}w�\��$`�^z�1zsR�g+���`���-�ᵏ�v�6L��G�o�iG0�V{ ���Gqʇ�jޮܸ�O��ᙼ��w�e���m��F�����)��fe��}[�^�;مY�Ļ�{�{��P�Z\��a��[Ѕ]��xS��'��0ō
�<����eEE�
r/^��3Z5�H;4�1��r""�h5	Od�O�&��#�FFCsݛ��(�u>�&��4���9X���9AT�qR��,K���)�M���9���\s��yw��}��ا�U�
�����h/�G�����,�rrL�[�=���hc��V��U���8W	H�X��Х�ן0��5'zq?d5�կ8�o��w�K|�o�b0X7��/H\��'�/�!Q�D��^��+��;槗(������3���f�2�llg4T����@@���,]Bl� ���m�)�sb���r)�`�i��=��V�,ՠ�V~�4|0��S(��JB����t���ӱ�Nm8��'xxA\��%VU�N[��VG=�;�1=z 9���A�j�a���(���t�[����o��5!m;�f�0D�7p�<FX��3v��nZE� �;����Ǭi"\o�+�i@M�yuഃɴN�=�AHr�����w��w����=]��r<2�&b-�N}��S*�������m�yMbj�\��<�~���Q�Z�;���}!׮��j�r}N�G�T߲m�QK���ϵ���|fqn����qbO2�mMC�ژ��‏P��e4�Py`�<=㵜�TD�r���i@ț���,�#�>��9��Ү\8Z%�āe��IC��]�:��6m�o=N,\�-��v�
�_Y��(�t�a҄NG@�՛�.b3T-��yB�dL?^�ؽ���S̈́��h�I�"�kD�}�_N��w=��^�q�)߾�چ^9��@xw;�U*�ՖT�������Y۔����_��(L�>��Wl�<��	�V֝ l6)�t5�LL	�2Ri뻝�T�rfk�4WEzg2P�H�*g�G��V�z~��s*� ��}�Cˣ��&���X�vG�����H������*{�i5Yp�{Ky��!�p5n<|�9��C��n�8����Eb��_�`8u�{Q��a{(e�oj�\6��,դ��S&�uzF%��	|8� �JG�'pZ�<鶪��z���P\�]���.��pFh>��u�U���Jꑮ7gS�@UmQ�R�6�u�:��`q���{<<��F�B�Ԙ�ѱp�2�]�z-N�O8�N�+�W��t4D���#��@�M�t���c��R��\�C����r!���e���ԫ�Ls8�dɨ�}��82.b�gL�B,���!�7K�tp�+�4Gpl���u�]�ڧ��XФ**��d���^� exUp�r8�p0\�566m��$n�f�SԂ%oS��\���!�U�q|�Q�6�nח�hWx��Au1�T^X*zb���6��ɍ��Â���8��H�F�C��v�%�
5v��-H����5fR��1��E@̞�Uw��ޒќhV����@��QC��.�ĈV���[����`���J�Z=
�Ǳ����xM[�~ddD�I\�=eòE��$C��p(�܁�8/L�r�&\��5�y��5����û��	;B�����\lT�ȣ�T�8�;����F{ߡ�/�0w���p�@4%�E�Ӓ���,we���6��v���}V�J�kQ�I����1����drm��g�].����*���1t_q��w�9�]��CU�����҈*v��J���[m�Ϋڈ�烕gXYs�}�d�x�hW�Xn��Ϡ\��+|hwJ���r��Ҧ*�v_	:�6]h����٣V��3!��68�:r�X埤M����S�T4����,�|��BM�����_u���=�C�u>uS��Z���Lv����!��xP�E^��C�vC���a��j���wRm��E�3�cʇ&K�3�`1�����JG�o�s�@n�6��(v���Tv,�кR35}���㠮ݍB쇖[��m>:���V�fD'Z�`P��V�[kF�e;���{څ���Z͞�\Ḯ��K��α����X}Q��ͫ�Cβ:m��GF���45H.�{���nV�j��������4z6@[�}K��ܹB<:a)���H�t� 
�vR�{uQXFI�ڒ���zqJ1vÊ��U�FҊ�Wm�v5O�Wn�X���`��c-�pE�2���>�=z��``3��4�������Ρ�X�:-اr�����+�%�� 9:����d	�X/R`j��뱹|����G	m�gU�c>6�Ɓ����<����\(Npv��(��]@�cnfJ��(:(�b4��ۘi��v��$�h�X�K%��_	څ���v�촺���+��1�^��i�r�.t6�%<��iɍ�m���᪵gbyB�+Tԧ��[EH3)��V�X������x���70�*I����]��ͣn�r���/Y}��dv�N��(�r�m)�(��賻
�����`�+4E��V�ˤ�^�$ �I���E%s�+SK�{�ht��3>��bW��@��]s�E.�7+y���+(>`#�T�M�W[�q�j�n�N���c���r=��R��2/jf|;~t�=�!;������v�(b�ZY)�*o�QR���ޛ����a	N�,�W���E��+BA�֐�Jf��	�U��efg9/r�[Q��`u�W�E�B�1"�9Nu�y�!uǮ��v�8���Bh���[p�O9�)v�*r=]Xi��6"xK3���P������(�^�Z�Jx��v�͛�w��s�s�i�)Y]�t)����'j-VGf�Y�6�$c̣�򁾮��jڝMt|��'s��˺���ܣҜ"�Hu.y��9�]M��g�g�k��Y�Œ.���" �[H[dX��V=�d�ZT��!��&!R,�RE�I
��`Q��d4�B�CIY������5C2ʂ�Xd���im�)1��)Xi!*�aed��@�&"�9V�
�V�����f�f��!m�V�H�d1*XJ!��D"�C�H�"8�
��M$1�E@P42Ud�@�"�Ԑ1�*,�CL��������g>��ӎ�@��Ol��eU󧯠��k�t-�3eam�+}�f`��RhI+������}U� ����xF���>��h�U��6�����\�K��U�79��g\(��i��4)�u�1�wl8��P: ȱ7V�`5���#!�ʞT.+�L�V���S�S��U=���6�u
_p�A��R.�=|���;�Ej�7=�*6��M������;e����ڦ+X��*�}�жw$�̗�s��%.�`�W�,�"��((��_`���c�3�LC�C+��ŽCu�b�L�b}>�!�@������s^��r5*��> :e�R!`ai0��Z�����]Zgzv%�C+��!"G�C�r�dt>��k�on�q;|�bB��V~�|J�s��dQ
�'��le}C�P@P㣠s��d�ڹF�RNd=���h�������S����A| 0/��tk���;=jg��u�Dǟ���}[��~���76r�U�"c��k��}���a�yO��}�ݎ�{����
؉����`]�����|��� �7a{ֻ���<ګ��ݾ���s�������B�{Hܭ�R��a��,��N�H7�����e'�hv�[��ݷū0܌�7,b��ׇ�����w�LF����k"x�\�(9!��شv��ý��!@���C&��.id�l=�Ɏ�T��)v!�PFNCscڨt]�Tt3O�#�V>˃g��㶬�U��*���䅞�|�������ޟ�����P{��u>��o��3^��E�Q�#ƕn���FS���y��)��	�S]ϹE]���u&u�G'LG�
�rh�T
2:&���ݍvp+6!̳}�O�1ض*β(���ޠ���墆%]�]>��R+��:��;/��ϡ�y\�z}����pޘ���ؼr��p����X���[\��'��T8�)jX�!K���
�%��>�VP_\��Vk��*�#3���k�s���,:�����T*�"3��L�
UP����­�������oR\����V0_��6
����"��7"��Č� lb�D+$���^��fACJ�����K�^�PV�f.۫�*"a�v�|���W[c{b�=D�D��\�u��Κ�w�|�}�HE^m;
�3�R(�'c�G�}w���J�v�"mL��u}g���  A��7�ws�j>�!�/6��{�tW^?�H.�xZ����Qwa7�O?x�͍|�4w�G`�]/U��ۏ���Y�DE�� V0dljY<�0�#Eʀ�P�.BrrON��D$bdu�����#2gTF�]����i��!��:��#iڋ�Uy��t�[����![��aU�ZKP�ت��z���9L����߲m�QJvp	߻��ОcN^(���I�gYA��D.<+���N�^T�,p��ɗّ�bR���]���`���~�y��F��p�h���H�.j*�*��=x{Z��00l�ة@v!\ا�b�u�S螥h`eA##{1���ɇ�U���D'��L���gT�siר&���A"�kD�"תZ67C����Hi阭�lU�����b�Mʱ�"%3�^][�K�(S�.����̴<X��d�On+�jN����������h���o�ױ;�#��̡`fu��1Yɘ�[��X�Y����y0�F��1K�:�LL��̌��uf� �]�������j�R�[� x{�M��uӽApH�
2��O��JNt�x.�e��9Q�ws�l'sxx��rw��J�}	��Œ���n��M��)FT���h��;$�yGf��n��X��W��Le_�Wھ�*��<+^�1���ϧދ�BA�"����JUyx�}�]�Y��U5B���P�KCAӭ�����*�����F� ����\\Z�NF��`bu�]u�A�����`��7[��eԊ�j�"�"���}�[�nm6\\NudXJ�����ö�hI�v֭b�!� ���II#�P3��!�7I�tP�+̦�qn)A��m
ÙžM��:�eI;^�^@�*�E9]8랆�`��L)��:�}	��/��� s����*WD�p��|0@Nh
���q�2w!NC�Κ�Z����ci�;'[2��њi�h_i���t��&q���0R�꼢q*��<��{��]Fy�;A.��&�c̥��x��1��w�'ޢ�����a���5��][܎�v�F�n���sz�KO�;}-Mw�{�.:�뽤!Q���`�Z6iܮ�	��0�w)������)C��/O@����g��nˊRr�X��J� �F���A�\����i����5�����["��6�^��y9�#�����ub:H����"J��o��E\
.X$C��ʁG)��G�*�L�r�&\&T���U�Ri�^����{�%J6
����ةH�/��E�*NK���T;\��{6r�� �D?'X!�O�u��"H�W�..��M��x�
q�{��54�Qu���F�)VDƩ�5���!@�"�+Md;�n��'��yR/�<�n��ͯ����4��y��'b�����]B�_p�,Ks�qдwn"��0u4�.9���}|\lX�CH�F����谝�����i��oFJ69q��FS������7�	�����h�^��ٯ���c���vS�!�穪k�q�9s48O�@pD�nje�z�ʌ"�jJ{�o���:�l��^��W	�2͞?M���툩�X/������7Pؽ��$R�7�*�>|���سL�A�t��&5t�T��Ahئ�{�6�N �b��׌C��m�5�)�jb���֣��E�Pn�oe�������N/�beIw���f��%��J����y�Ҿ�4)�9p)���+\W!
��.B�����L��\��8��V�X
�X0:N��'�B��8�Ǳ�n��r��GEFC�'��m �S���jn]\R��و����VR�0����Cw�0�26<�q���yh����!����	�Ӭ��}h�y��=��re�o�_��q��P�e� ��(9!����&ţ��>�銶�bdj`�^u��oR({�`�
q
TmH�-P!�Q���noڨt]ʎ�R>>M�prl�u����w[}uC�X�R��䅟��v~���eY����ɨY�kz�m���ʎ�d��9*(�����@ڃs��F�S��N����q��lb��O�v(��Qz�yO�!V4$k��wX��6>��'1��EC�dQI�ސ��""�-�vJ���C�5PgR�^�j�xb3��rx�֏��]��dԩ�p{T���%t�4S��>GP���ΣDwh�g���U�������6� ����%��\!��*&ގ�qd��c7�ỗ�j����4�ȡ=�57�����,�즜�6>6$�����S��<��>�uQ�_T<ʲ����#e��j->INw!:6e���+�b�S���(��S����+�vGoP�zM16��J��RK�۠��u{&�3���NI�Dex�ghR��k�b�}�C����릞�����V�e,ՇC�eL��{
�є���<�bnw��*M���*�r!摑�뢺��'�����b��P�y�s޺��9�z����3��$WK#Q�.=�M��U��Mt�U��� ��k�^x{��u�+�`P=C�@Nw�'�nz"�12:�۽�p��*���QOU���p2e���W�P�BdtW���l��	j>}-ʄ���ea��:���=�5�XӂѦ>���.�o�^_'��eY�!E�[�T�u���=��5/;��l����<�Uq864��N�v�����b�(����=�[6���q�;~{��&\��D�Af���i��ޔVBƇ�ŏ�۹]�qr�,!*>�� �+1m�u��%q ]�T�T�pNJ�RV��p.�`��w����,۳G9w� ��w4������6����Xd&w'��9�	���|>��"�т��3����~Эe�XS����u8�d+��>����~�\t{:��ȶt�m��yD�ā��&+����̜�nS��{�k��^�@�0A�so�ϼa��ۙ���C '>��b��r��Dz����vU`���C����}6i�pjH�"�N@�P��Wh�ĩ.jf�n���Tz�T�3��9��u�AI�c�������M��<�l��u����2֓��C�^�v�LJ�TAZ�R���t�z�_��\?S�=��,�����X�.�EA���Q��h��qy"�Љڇ>�
v���#���m��'�?ء}C��d籣�jpAr)�����^CY�]�E��N?7龡@W�PΓ�Q�Ud75�B��W�7b��O��|갸�=F�w���冺�����S���&Lk����ʣ��C��Aa>�I���MV|x��R�iZ3�M$�\��g2�����NwZ1��)��Hiy/1��֭`T��+�*�qPU;-�<]bs�}�UU|$�z��\�,W��U���Kt�[B|��*�q��C��5
�u>T&B�gza��ȶ�=��G�Vz$teIN��
�@ʪ���\랆����=�R�(�9���lV�ȴ$c�*d��ҭ�W�\$uyׄ�Nkյ�'';�c�D�nru�ҋ�NT:��t�fA��#��7�F�C��Q�}k<�o�;=��%¥,e�qfF츥!Ƅ��u�����"�������C^�W����
#:�5���!l��6�oWC�����N�D7W=BK�MJ|�vĈjD`� ��'~$C���Ssb=�W�0ܾ	�G��1�!�O3Z��������\l�9�
3Ų(��T��੨�O�u��e�����;`\c���-��@�/���(�wJ>~T�M����R,U�gr5�l
|KٽT*���"`�U�h(��tEȃ%�w
����a��3W3�	��Ŭ�z�r��Wլ�+g�+�ҜM��I޵���q�D)����Ϡ���#�\�i��h���5<See��%i��Z�웦S���k��Xw,^��ȫ�ى��/�#�,��!�rw^bj~��  R�����1Q�̌�|���P��c��_ʄ�PT�y`I�O�*�vO[�_l�[�6�q����(6r�bq��@O���7��Be���Y5�I6��psy�Ec��2�Cu3�ɠ*T�}Q@��"�DfH��O���U�	�s�w�I-�q�k�5�qI����'���GB�>�֨W�grT�����h���<�f����~�CrE�Ϗ��N�^����z�cW̪"
��lK�Ǎ W\�6\q��`'aA��7�Ua:Հ�����ZҪLw��w��뱎\l(6Y�ا=�@<T�F�l�SLRدD�DlQ<؛��,�R�����9
��Qh�?���}?g�����r�P��L�3\e��sGwYM;�^~�O�+�å.vd�:21�=Y����w
�Lp;m�b�DmHnD�d���s\R2TC���&Ǽfr�����zD��#��(��a.n�ː��3�Cc	Q�,������V�l�H�{w\i�e��$�� ���8�(�[�aU�)F���@�ݕ/{T��/P5b�Qi��i�oh�us�W��M��*���W�	JSX��_)�K!yp�6
1�����g�8���z��w����"W�Wx��J�.Em�+�H�=�9�/c�w3i:r�n����Gd�L�!��n���[�Y[��Zu�R�|����Dv�-��ˑ������{@Cw��joQ���84�������W8>����KE.���w��eފl�r"��n:�1 ��!����������6���iB�0��u���A9t�����e�c�F���Z�3�J_X��Yh��r�)R�s4�j��}�N��S�E�>�<<�d�Cw�����)���_x�惷���IFUD;w����k�V]�Q�A�����{�1$c��KH��������+�r�]ٹ�����ŖL �[՚���W<�[���ʽ]��*�������s.�oY���}�*G3Ŭj�tF�w�N��}�eӽ�[��: X�&F&�Q�]��c�Ƹ�/f��g^G]]�rCLV�8Ξ� �@:	1(r����M{-���r�/1b����[���y1'�3�R���:\bާ��.��'���Knᆗc��+���O�5���o��@�Tk&f�]�%˚�9��4�Cr�tcE�ث��@.���mU���^�9m_���߷�\�MD��Ԓ(�i�w���S������j� �ݧ�Cp"�iZ���� �լ�IѺ�N�>�|؆����`Zh��-��&���JumA�m���1��9`����SgVT�uxV�a��9������[�����u^��0ٵ+*�1������iw�Q�sWn�кj��f��4�V���xR�oW�u�8�QĻ4wuj�+�Vv�p׺��G�m��YI����K��՝L��aն�ƭFo6��,�4��7�+X��j�`br���t{+�pI�!ᅃ��єv�[�]	���Q�Z�"�\�4o=`gx�%���%P��zdz��/��؇t4����H,�Ӥ
4�1�]WH�8��{��,DLn��_`���.䧀40�g�`��ƣն�,'1j5���\XD���dԷḪ��ɢ'%�\�v���>��Et]��	�0E �]Y��ܮ��C���:S�m�S��kY{ju�w>(�狏$��%i%�r�W(ʌ��(�����=}��w�u����t�T4��L�!*(��
�b�d+�!��*�Xd�Bc�L���J��1��2B�X
6�H-dHJ�E��I�VM0*I+%t� 听X��Y+�!S��T�5!*J�M8��
��1eH�bȰ��P�V"Aq�
M3H,��D��
���C�_[�T�{�h�MV��;ۡr���f�`��}�����H+���%��҆�6f��]�J+��_}�}U�sq�<ct_�K/!g3�� XR�pOBʨ�pjc��W��Mɀ�5�38�<ɦ�R�q�X�[�7~0㌸s6#�P��FL9P}GNGg�C��P��Ӛ�IF��f�3�"]����A��&[��Rk�>�BVyTYK�Txѵ��߯g�����z��(}�[���uȈ�����ɫ��Lg��
� ��c��F���p�m���*���~����1��ߣ�p��f>�^�ƙ�:-ǯE?:f�O����L�@�>qT��e�̑�~d�r^<˵�����կ�_���*�K,<�P��j�].���ǽ"�� J1֌��.��9�П1hX�����y�܋���eM.�'D�ݘ�9MȱS��k$�9�����ޔ�m~���[-��.�!�Kα��:访{�j��A(�XY�N	�۽�6\
3��(]"����v�ϣ�#�X��K����v��n��7��ְ�.B+H+��[2��.8��0���W��Đ�V	��L�h�{�Z�-���6pX\�4�+�X����Y�W0d�9:���`���<F��ݫ��{��3�w�j������ k����s�y�*�rL�1��_UWݶ�ɞ�Q��ѣ�vSU�
��V��]���� �##�g U,��a@��Op�K9��E��{FЩ�"!�"۵+mg?��{�p�/Vi�p N��QcI�rf-���M���T� dN�FӤ"���A��{��]m���,�j0Vw o�:�}~��ٕr�\�%S
j�s���ɧ@��"�Ce�[|��j�=/�����gr}a�r�9��G��zquq��Hf[���l�ʲ,t��JέrB���F��(��ctQ:�(h%��l�
=�#���.*�e��Ω��9
!��sV#�f�	��9J|�I�m����_�j�{��
��ס��R���w+��OLY�m�<?F���r��{F���b�+��m��Nt})H"桹�`���r+��v1{He{���Rv����h�e�, ]�
!������$\�#�i�P{>�E�T��Z�1 K�<ͯ��,�z�3,e��ñ*55o��K|�5�|�xMk�p�.ut�%�L��Ǖ�����l��iHܫ�𫬁Ն�W�F��߀xxr��3͚�xk�T+���S�v�L_ 毁��[�<|g)�ǳxí��m���gF�Y� [�b*{�G�6U�Έq{"�Љ�>��9��/�����G
J]:땆�*���.��9�OE��kyװ0'W�{��\�8F:Ghh�<-�r��.n�T7d�ȝ��ʁ�e{��v��vˈ9+���i����U5��>T�LS�>�t)�"�!��aZ�	�gA����õ��6����i��o�ڄ�K6.�;�}�$!k�\"�r Y�["�E��)�@ƙ�����(i�\�Nz
�S�<�N�~u��	��t�UM��5R�w:�Q,g`e��]%K<݅u�4��f�@�B�H��^�y_z����)�;Sw�)�yО��
�^�=��qeP�6�d`k�ʛR wj��r��nGc咴�\1��Y�I�P�Q�'��P�s�GC4��Ϩ�@� ,U�ҵns�ͥZ��ڱ�x�\[[�t�l)�1[�5C�կ#{��$ݎ'%�\ר�����D��}=�y̵㜩u&���G�WPȲ��W�`�i�U�[��U�������ŀ�:9�Yz2�����L��N�NЅ# G�)@����H�4.T
)��G�)g�e�tg�Ot����5oC7���U��/(�+)x"V�@��Kb���+��USE��7r����i�Cr�{>�)_��(�R���y`�FY͖�܅]�h��N�]%i���zG@���s5W��*��t�g,ƥ��
�z�æos��;��:�d23ȶ����z���_g�'b����ުf�pz�Ɲ�j��b�`0�ۙ�q]��23��r3F�f���*��Q�Z��f񈷶����SP�r�C�S��<F�A?y��v�<U�m_I��+3z�nx�$*Q�~���.u}&�t��Q�*�U�
�}�u�B�_C�/wJ�W�]���}���N��.>!�..]���9�����"�PP��9HG�9�j���e��-8I����Nt���ځ�;��9�T2+lq�'cc=�ʕ��Q�^�i�lgz7��r;�9���s�u[��,�y�7������nO)��|�B>3q�E�*Z�*S �f(\�;[�����5��s����o^pS�Z`���11橃!�}hhcz�'fj�*�(����x�^��.�r�J�
�\lWOd�Mb�2:���ĺ��u��z)o�'.Rq��d�쯘?gB�z��Pt�8��F����]_Ґ����}�cV&'ǖ:�8��36��O�z}>P���	e@��QpJBTts�v�GTgGx�Y�v��lI�1��
�"���L9�"�VI�4E�:
��nc�H˜�N_>y���Qѣۃ3y����X5�@pC��Y�*s��w�nN>� R�|x6��9q�.-�`�9P��raʂ(�ȑ3=�v߳/�[���l8(c�yT���gT�m29:b<�P�rh�Tx���HE��u�{g;�z���k8�,\���CSrީ��DEr�AJ�&�T��J�B�.��/����aH'�(lT��o�������g(*��!-����/��;Վq6[�c8V��+E7&� ~�8�Q�T���8@�i{�w�a���T[Z�=d�ְR�����s�Ўs����\�I�H��!V��~D=�w��  �˓���YQ�Wm�l�yw��#x�R�ܣCu��x>�0�rr,r��N-�}��������f�����q�욼g4��J�5j�xR&x�	H�/���6�V$�Q��&��d�!�@���!y���T��D�q�mA�-�B*�����gL��s�:SCL� �<�z�D7 �α���V�D�C���ɨ��p���Q�^C�N�@�>Ƞ�*	R��-�n<a�V)�=��䠭��{��7�YX��	��(]l
��.Br�J��Q\�h�-����8ϳl��y+��0�C� l�p�2������l��d��}����xN�]��S]�alj�bV��b=��DF��X?gƱyu +�g�W�����d����=H�n��ё��u��~N��&�áA�r!W�q:;Zx|�!�"P��r1��u���tp��3�����d�M�BEx*P� (q�E獵����g��Dixx?P墝]Z��ծC�A��G9�O�8�u,���ǗwI� B�����.ټ.N�س��x`�M�vWp��7W����W���m0�����xu7���pv��+ɕ���.]$@d�nan�B��P��Wg���?2�v��ւu�a��{�U��hZ���,P'�;�dq���EA��.,p�3�3�y:
!�A�=mwc�gW(�&�?)3�=`�rEIR��d���T��ewP�qo���H��N�f�C��>t1��5��#�F�����TJ��f�I��Ʒf2�ZI�Ï[�����/Ң!\�R�_Bs9D_�G�{K�nυJFxڦ5kʜD��:Ҧ�m����H#/�ʞk�Z;bc*�QO��J\-ա��*q���Z��d�3+��]N÷^���0�+���Q��W�:!�승�a�����|�B�*|DJ�YN�`5�V�tl L��==�S�����1�SO�vr��kf�FM��A���*ECu[�d���P8��r-ڌs5�rv9�D&�����_�y��{$tx0>wHPnfQ��5�@s��1�҆H�-�j:��6�W�
�a�	�,��H�ʒ�ؔ>F�u]<̕~����}��ݔ��%�n�e,%���׮�r؍>[��]H]�U�R9����S[�+�:*����t���.��<P��Y�i�W���ht¨���oldwk_]�#{MŢ��6���|����SJ��Q6��oo}� �cm�u��R��ٵ �B��27��E��%Vԡ�GS����{)E_Vtn��+eҥE��<v��nY��(<�fA���o� u�����lA"���ݍ���x;�Uy��A1հ���=dnˊB�������Ĭ7��#>��#�=��P���t0��f�rTz�eA�8��
�x2��5�i�}6��Y��5}&)C��CE]-�}�P�c�h)�"W�y^� e�su��kX[S����½u⾥��.�����%i�S
Kt*#��l�x�ou��h*Z�f�(	�b5�B���44R��y`��ܖxe{�8����o	ge��zh�:eRs�z�P�0~}�������L2�O^4����eg��J:v&�T���`f�m3�#)�g(:�n���v(*}���9v�������r��pJ�"�\`��s
��W�X�QƘ�9��y���>�3T�G5���2�fMz�[��]%wFݲ�iзE2�h�̒<A�w��̩펙atT����*b����d�glL�|��S����(1�ׄ�������8�j��{)=؟	�|h�t�cA�R�pG�R�w着�>/Oz�]�`�e��L���V�?.$x.�����ؼ��h(#\+X����z���g���zv���`���02���P��WKsP�vx�[����M�Le}Vg�:e�ˡ�;9�����$e�C�FJ(:��lSJ[w�T&:hWO9���
��8s=Nʡ�[��:����w�;ԫ\�F��W!�UѰ�J�
�\lWOp� �1[�~�nO��o;�/�xu��e�s�S_/|�̸�b7*�9
=g�Q�]t4-��V�!��ݴ&'��x�i%�,5��<���	��:f��W���
P�"�s�Jz�aA�e\���$V�����H�R����η��j-��ý�� �J�^R��ޑ*a�A"�e�9
�u���֜N\Y���EԨ�|)��v�ǜjTN	�YU.&#�;�,>��(c���$Z�V��\*[7�)I���'~$K���䮃�TW��j���@����/3�i��jE���W՚�#Çm�Nc��<���-Ɲ�^�ǻ��V�oDs�da��'��.nɺ:aޚN�u�Ύ�K�H<+��7��������`LQS櫜3���M9�.X£�>���j�8���_�/��')G����T�o�A:b<\�"��Q5��rww����A��u����/��#)���0�*�P���Q��/,�����9x�����E_
+�.$���U�vT��� uf��Q�T��ï9�k�ŵGf���CD���)�59 ��yĂQ��o�NPY��[q�D���whж�ƶ���,9���Z�^���Bw'�%=b��C��ޭ�k��
U*��׸�C�ٯ{)[����a
�u��j�&��l��ݾ/_N5�G�D�$<筣��C�#!']�0�2$�tipr�f�1����P�pEm(>��g��P�E)g�ȶ�qX���{�P��{���)M@��""hezwN���`YT:���X�<!w{�1r�6n灋�����/�{�Gd� l�{�С2�
#�S�m�!��Lf�W��r$�g�0O�"�:63�M��۶Z*���ڻzN�w|c�B�Q�Ysep�����aה9���+�N�n�L�|C��n�X���os�ҭ�x`�5+)��b�{!���9���璷e��Gl�L�z
ˠ�F6�"�ӫ�;��:'Z�비��^�D܍��ט� �U��Q�IGf��,����ing\a��x��.OF�hאH�9 ����>�y\��x�P�+�PZʢ��ZA�@�V}�0	*�&��9�뮭��C$�������v��&bxS��U��X���]S���G��[�_QQ�Y.�N��)Gu���#s�ܜ������G}u�@�(�s�Q��ݧ3%髬�)'fS�[�i�׻�U�$:6�;[����d���)��ª;{�`��+��^J����h�x�r��]��*�'b�z��n���,_uhN�v�p�<�*mf+ukuhX�����b�׳��Ί�c�M��p��Ыy��R�%q���.]�m�#���t;�uKa�B+�Li�6�(bb�q�Wr(�t&k�!*c(s;r��M�!��������Sq+�Cde�^�(l���a,�����O���o�qڼ+�T��ǭq,Ŵ�H��'Q���` N��Tޑf~�J��v�ΣF�ZT2ʹ�1/c�IHn��Ե�)� �3睆A��p?Yt#�b
]�fEVҖ���Kds��|���Y�j��\c����{|�b�׏%r�-���I֝�5W4%+*��ـ�WՕ	�h�G��.�^r�f����銳\��Zwk)5�t�2Wy2vެ�&�;�z릫T,6���&M|=�ͭO��s����6)6�f�9��޴yeC��M�o��GQ�<U�{QL2���� �72��BOqO�ސ^�̝J�S-^ý���HN��+D*hވ�n�[ׂE�Zq���8��7x�j4jB�v����R�f��듚�Ay��hn��w�7���W��>�jt�lI`�x��l���g��Q+4Y�A�2z�бu5m�x�w�:���h|&&1��l:[�~�D��s7�,#$ת����8RU�yQ�O�1M4�O�̇�+üQ�C��B�n�ܹ΃�ݪt�N�n�����nɹYGM�A`�@��+��^qV��ݡ�u8�"v�Hk�͢��u�`<D���&p�;�zm�)�]]��K�8�̡�ζ���gq���>&w.��5r���V�T[Fu�X�F�y��w�M��!���Ccq�*H�iV�*T2��t� �Ld1�P�-�\��̸�f$1�X(d�c��J�3T��M$-bbB��X�Q`��JEb+Sf0#L�E�T"���4�$�a�"(.!XUPP*@���\b�T1(�²�`��I1�Z�2c4�IH�X,�Mf�fU���QƩEEB�Lb3MEFj��c�l�q�9׹�4w���_u�~���5�2����d�^'V (��^)���a�[���s��(��ׇ֯�rqW��1W޾��*;�-L�g����Ѧ*�ύb���
����|"U��	B���Σ�2�m�q~.�[w�+�	��̡�H��T>�5�x��KS�T��x�c5c,rޙR)�t�\WKs֫�]YVu�>n��W��!J�:�i�3�%�J�,-Q�ǳg��sy.S�8`�pέrB���F�X"����9�t>�+=g M�JH�p��EA�e���0��t_b�t*�9�b���x���횱"�tG��>�R\�220n|riI̧r� �S�w#�}ܷ��ܪc����ܚ����	�7&iKs��j��z9E�ռK5#]d>���cV���TDO���k��u��.���� .υo��o�h��N��PQ�aO@��%t���Na�tY��P��}c�Y֧D��s��<�gRw�Cu�6*r8�G�r�̮X7�G�L�͝��+����%Q�}S������$�L쩢�p����䃐R��b�,Os��:�v�{�.q��Rf�Y#��!� )�Wv���򗞯Md����x'R��]�l W�'ғ,�69��ii4�tZ��sW$�q��}UF"���z�P�Hi�P:b�����T�*����5��
�
>>ҵ|�N�LF���4����(��ʕmĊ#޶�V�8,����"*:l���c3�J;J(LP{�n�*q�P�f��H��3����F�h�.�9� {�)l�a��(w��=��Z/����+�VO���׌V���|�Vc����!B��Ē砩�9S�2	7�0U�9Z��k�����X�N&�(���r� ݅�fF�|n��ED�s��9scU�*�;��q��<^��A":�iu��F츲�k�N�$L�i�Y�Թb��*��Kr l�[�ؠ��~5�9J<D=�#��T,��w^�U��%=X���lR������.$B�'�DE��P�P(����pt�M�<�K2km�����۹��mӅ2�7ᨴs(�9G��آ����? E�1
+�"�m�N�ճ�l��۪�
]t�"���7m�d��]�ى8�7��+�6�
r��.5��)�i���t6����6����ŵ����KZkL#PsH��DGvAAޜ��ʪ�s��X��&:�}�I%Ar:�i����'�X��Z)A!�+���vTs�{�v\6����
�p+*��ޠ��,%X"`��V!G���륌՜��P��P}YX��F�f�@�ϫ%��B�q���q�;z*u_7˲�+L��u�b9M�R.
�NC̥������+V��3������z�]bn� �J�gԦ�\U���`d���<���M��Cy!z1���.�,'���8�����!>�((�L�8d(/�"�ok���&��xƈ�령նψtˋ�T�v��{G1,e
2e�|�W�L������ �a�@Q�f����\OKZ���]�^�h�o�ʬ,ՠ�C�]�&t�,��Q=#��B��eB��.,l�����nG7@�~g^L������ըZU��^�Q��EJ�!_��̨����e��+�%9u��/8����N���L�hm�<�O^�<s)J�#*�T�+�{z.�v`9�.u��%1���<[�/-���4��}�����n��p�,��1�����Djxw.A���k�T�bV��������a����NO��nؘ����'���#P��g]"���W��ۻH�F�eOY�b�����F܄�D���E���~��@{���5y�/`TB�;f�{�j�=�G���Z"<4x�83��:G����i>YVDV�{���v�)��l�ʼLu.��L@�':�[���s>^J�o7G��f��7�������A)����:z7<j��	�p����(9�&[��PN�� ���&,�we�B�
�;���!\��38���"�[��z��B ���M�g-�q$�g��&�W�k�)��ắ\��;*ˋ�]��<ż��`S0þ�ض���yP344O�D�8*rS�J>�}��V��s]ǧzB���o:�|kaYW���J�5j�xULې��'q�szK�s{��R)�P��5�
͊�M�x=�PX�5[Q]��Y�~�~Hs�^B�@�yL�{C+6"��X���>����Y���`���I�A���Xu��Ez�W�0N��n�7�;��o`nm�Jc��e�yD�_*�1���ɓx�َ�)wc��vwy�����R��OG,MM��+�����vB��\�]NC"��bG9�����.��lg����r(�#�
	��w�+��)ptpEm("�P3��T(��[N�{F��˽Y�s�u�檪���*�
������-��48U���C��NW�S�Z|3{e�כ	1{
�{(km���C��
XJ��H��J���������Ӳ1��DU�;=ː4c�|�S�P���k�{&Ԩʐ`dH�H�����ӻw0w�Kȣ�)|z}ŝS~ɷ!E���ua�}���áA�"}Y]TF`���&W�z�#���lj�N�||�=j�ՀU�S;��l����#b�Xт<3���S��.�s�A�٫�Qw��Fuk����챞����K��i3Zr�(���/T��"@r^2��O#:��+&p�a��adu:����DtGX��MX��fo�D�'�)��S��U�����*H�A�G�ѴFR�ee癛QxV�U��:��������n�C1��=q�������0'��qΌϴ龂�րʙ@9�+�շoV:�H�t�����Hv��.�������uY�ۊY����\�b��Ӑ������%�ұJ�\}�lح�c�;�7r�c�L/��Q��[����~�qת ��'���s�F���X�֪�w6w���lQO�q-��}^@�x�(�)�oW�V�X�7u&#.-�Q����ۙ���ϰ�!W�09�Q�e^l���].��r6�����K.����Y�r�q^�t�.�.�OXzz-O{��I��/�H鮬�v*o)���W
̢��R*���#'�j�(�6i�k��H��gN;e���ЕwI�jvf�`�4}�>F���~�^k��pL��C�s;d�t�u8�y�]}+e�Z-�[K�F��g���B^�t���AO09�= ��JS�6�B����i�������z|�� ���W,[���JL%�^R5L�Q7|\g����nY�݅s����K؊�����z��NK��)Wt�6�8����ir{W��H����`s���J���pX�>��e���Ki�_�UH:��'����%��M,G;����m@�șӃ30ѩ�+���؅p�Dқ̓)T�W��R�x{e��s�bo�/��<8W�e�Ճ���
ݗ�k���N5�0��5�'*1�w�*@o�`��N�O����ʂ0N9eߣ�I���Z}�{,�QƗ_����K��A�]��d���D9�
ڨ�q��a��y-���>��B��˃2�2�(j��:%D֊q=9���Zf�G!�kz�a�	F�����=9�Dt
��'s�!�O�c���\j�����/�E�]��U�&0Met1Sy$Z�M�8F��ޠ�T�X"`�U�i3\ȫJ'��w��#��G@y1s�EegK�YFa�>��"���� I�{"�����x�0�;$�d\Я(����XNC9�F���yTea�3�OKZ�qz�[iT�>����xi�A�Zi��kʬ|x�G��_��a��꾫JQ�����D:;����ń�_B�g�����'�\((�Rܓ+L�y��d��G�Yb��mu_uX�<�o���.����L�	�������ի彂2;�+����!�h�XEC��>c)���"���7�泽�ԃ��xEk�mv�d�� t���Tt��Ɣ�UV��ҟ7\d/�k�Fe��u~m���m�G>�3�;���2]*)���;h7�a\)�LA6:��p��ɮ�z��'a��������Sj�'1�7{ڱ֬B�"^
��"� U>
v���;��w�D*��=�<Ò{K&�V���O���d��#H���y��l�<���J�s���:ub��;�(���
����bDLj�f��o���EP�D��\l(�n�[R��'E�.%$���O�=��#T��
�
��%�V
�.)��Ps��y���9��P躱J:��9:� P�pOB����=Ω�jz��
n�aM^'Ы��Ɉ�:\�;�"\uˋ�T'��T��\�#q���
��Ԟ�m5Qv�>�����Ω2�drt�z3��ݨz��Ŝ�����4׮�
T*ǂF�����?M���x�f�;�أ�w�@���<�c��!$e�5���-\sdܹԍ��s39q�����4���-<�� ��~o-|�/�����e]�q�l��T�I�̓z�НR�����it��Tt���5��u-�ƥs�B�o~z�^������ ��ɫ��+X�Oh����';���d��.�Ԙ�T�bJr1n� )T�[ӑz����@�։�V�nH��X�8�ѣ�L�e�;�?��^2v���X_*�*�K,<�	U�j�]/
=W�^�	��)AY͒��B�*t���'�R�kh/�ج�[:�J��X�/ʭ'"`Ө�G�̆v�A	PXʃ"2Z��T�"=sCH���<���R��nA��lE��S��77ۮ���m��#���x<�[L�a{��uѥ��k"�ݠ���1gb7n����"qG�'�����Kg: ���4}���8)q���v�ڱ���-Z���R��d�9��۽�bvHV"F�׸m
�B28E�;�sg��U�RF�;�����o����{!��^}-��t.��c�R�*A��>�H�(F��&,,�=���v���^���M�
,�a����{�	��Р��8%�r1�n쬹1^���C��l =ڑe�o7UC�V��L¹�ݾ�k�`bV����Y���7uZoq
<�|�����2��j`�y������vٷ.V�d�Y�Q�k0�����#��b���S\���/��}�h;����@����%�s���]R!�L�O��r��+bU��2��+���b�b��j�A�٫�Qa�@у)�9ծC��W5�H(ή�P{���`�����'ڼ(�yp�jƊ�Go����mECF2n�Lm�<�������TH犔i�J���7K�H^5��C�??D*[�Y^pb�2u������.�ej�8*�Dw������.�FVұ@-��RVf��׮9E��$A��ӨP��Uէ��E�k��y�"�h������/������H�.q.���W��5�i�|���h/8Od�&w���/Z~����te,Y	;>�\=B��Z�
���޵�1���ܼ�i�e,����2!����}(�-Z�=m`�5���EQo���^0��y楨fZ��bȡ�:�'W�{=^����7�P݂v��`Oa��W5��P7�u�.�����%q���j�B�[V*:��K��M�`U��H�mZ.���4uFA��'��b;�8�:d�Yu�#�=�f��.�
�jEo83�����ӌjB��Fȷ]oѐ�L��&�[��f��J����SCe2��z�mB�������֙L�$Cs�|4ͽ��p�*�����9"w�U)�E�b;��np���Gҕ�|J��L_).�Ѥ.���SnD`T�kz�"�k�;�YMv�s�.Q�<:�:ܽp��s�2\	(h�x��9�U>M����#@��;�Ǻ��AJ�����t�V�0�i^�afܶJ��k�2�)hY�	P-.5�qk�z���u5v��M��sn-�U�d귵�}�m�	����E]������6��)��ou�yPehz����a�E��pW�V;-cU�h©����Vu5n�����`��N���_3�))A�t+�d�����B=���.�ܧ�=�F� ��mZۧBwbw���!�-�J�Q,Ֆ�n�s����7{���U�t�R��mn3Q\�x� >���u�B>x�́W�צ�k}x��n���)۳�pJ��,l;ޖy$^�Y�ƍњ{C���>�y�����VM��ڈCW-ͣ���R�©m�>b����A�E����ݱ4<Yj���U88uZ�w����&�f a�R��X*��5U�����aKYo��Z��Nl����{u�C�����LE�K䫎�f���^C�ls�qĂ{��P�n���	X�B�,X4a�k��^6p�hCĵ���@�Qw[8qg��]�ʔ��r��[��-[2�G��֟m_P��u=��|+2�Ny�U�wI�j�FB�r��)�9�K.�F�L%R�#`f�M��<��d�[���%F$')�]�����j���'�ǌ�h��!��Vb����g��;���%���`%ҝ���t�{���Ӊ��4eY��ʺ�WI������k��c�u@1p�V:ê��v�f���q���s9'�`�2jB��gfԱFT<�7Ab7����K�����G���p�[�
g&�5�r̭�si��y�K�/���1&SRK�]Dw�����2p5&�Ķȋ:�����ՉK�F[�r:2��V"+}�{���2��ڣH]����b¶���uu��'y�n����]v^�T�G��!���X���bK���F�+0�ؠVܩ���i�u�[�i:eAH�R�I�,Pir��(Us
I���L�����XV(��&!Y*Tl���^ڊ)����V�"��*�,������$U�,X,*�X
��4*Lj�`�T"�J�YM6
(�"�dQEL�.�U���aZ(��E#iZ��V�)Hێ ,�E����&Z1jȪ1UU�Ȱ˧�"��TX1�l*[Z,�Q�U�mKh�2ƥj)m��H�jQ��Eﯼ��s3��:��/�{onGl�=�Y��%��J�{ ÜMh囃&��z�Hܘw��+�G������$Ś��2����ܲ�C�ά�	Wt���@�@P����s��O��]9�szk_w��Jj��tV�^e5jy��^�ѕ*6'���l6��U}��i䧹�CD~�b(t�E�q=-NAr3��Cs ����p��ɞ9���c\���M�~�O�ؐ��u(�|\,���\���
�fFMˮ:�)�����]�R� q�ഊ��q?d>��~Z6���൭|ՠ��DTUbv�,�V���u��wySaH�>�}t�k��;\>t=����h�M�Ï��n�p�s$���Y5�����V#�D�jDH+�W�c%�P�;����w��4¥} ���2$�g\ùx�q�7�j����/W�I
0�v�:�o��kLDl��E\�S�.
���P��;���!G��^�.�2���5,|�P����k�cM�n�4!@��nw��#�Q��t�󯝢W��fur\�u=�=S�K�p���^��S4_e����ms˻z={t)�,��k&C�=e����#;�Q%u� ���2��Ң��މf��pܕ������j��
�����^N�"�)k���S-4��\M|#��4O@���pEec���72��l���B3��F�YzI�sx��r��跕p,j��OP3>p��z�\`���J2-��Af<��VWr@~����$ʋ�;w��d���D�x�$x-K�f��<{��ϐ��s���P�;C�P����G#@O���=���A���>9++�c�p/9>�|f�Q	�R̎����#Z����L��t7'c �2�z%��cv��ĉ)#ӻ���@��ꌟT�!£4(9Nz�&�^�@�NÂWE��}ӌ��w%bb�
�-�D�l`�q�P�"%�.,l���6�/f`�yNcK���I՘�\��v�?^z6c'b�xF̅`:
=@�*?��>B��A�Ƃ�&��]�ZLB~�m{����^DLo��4�+�7���#fG<�Tt����k�OTT?d���㣜��z��C^/*![ìU������ %ߢ��m��<�^�gdWY�wE�sFA�S�ab�<�L9G���Įn�.H����k�b.�n$��������=������G�lxm��\kw]�h�3{s��F�;�F�Y1ut��������5�I�#6g���'!9���E�Ҏ�i��ru�:>R�D�J��3|�0�gG1U*L9T�|��W�e�)q�>���1�L��f�m��]�Vh��@y0����!�Ó�'������Re�N�La����m���#�A�ᠸ dtP��Y�� c.*��+%�-]Oo��Z����1��DE�CU�5}^��q�!��\
��t��/��bt""������)=�7]�z���n�0-UC�]��sJ�r�J���U����F�>{�-S�5��w�7�s��uKgvG�f�vR��*!������1Ф�}�7�^��wm��u�,��h߯����b���Wy���ؼt2���T@�'�`f[q�9���<�����h�_<����M���լ���\�SY|m���^D�{��c�w�8�K���Sst��=y ^�!릗SF_.i�Ѝ�;����b�1�}��SpV��5˝�M��wXUa��)�k��j���+���F���$�e幽ݛ��B��4Z�-rf=��˱����2��C���3����ū� ���i��r�DyEʯ��~�H�y�J�:A�;��l�ֶ�Li}�S�k��k�e+�%:�Z%g{59̋4��ɶ�K϶ޢ5[��GZ���BW(�2F�D�E�-�bhF�9�W",�VV�-��G�)ApjfLcv�i�y�dn��s��"�k��nv-��]�W���d�q�Ks��m�5�R�@��x5R5��'H-vv�rU�nn���z���v�����>�b�@�Q#Q��A�8��m��Z^'�Tf���.ʌ��h4$P�:�>�x�Vk�"y�)������1ג�NQ�Y�ҋ	h]u�V�}B2�fz����}�W�bz��^�;���j�9A9��/yR������"6 ���a�hl�⾵�d�K�3o�p�a�F�,�lSʆ���|�d�$�WW�|���k�l�	���oQY��Z�af�h����X���W����LM�1���u1�Ԏ�y����i~�_�V�".�X�t.����'����;a�]���oЮ�6 ���K)S�ݛt[�B�W)}�OW��njU��1��n��]��]�Q��VI{Y�Ђl����<%l�&,����u��vn'}]�A��D�7~��_=��gTƫr����Y<�ͫv�n3�-���"���H�Y���a�:����P3�&�j�B�y4���c�}�V����t-��c����7\��q�3޵<�M~����ƭ��.O8�I�n!��%:����ΰ[u~m.��:�ȍ�.�_1G!��'�O��l�� Um	h�ո^�Vѽ�;<t���L]���O��]�g%z�ݾ���El�D�y��7��e��0l��׵�7p<P��T�xeuܖ�rڹ}hOFuYn�q:u�QCP���\��5u<��8%5r���.9P����oM�.�D֮��Ie8���w�X�X���^�B��]��P�۪�_h��Wu�������^Ncz�#^�؄����c�}����F��Y��.WgG�ߓU�2��k�uU^	�أ	��l��܂B�^�A���q�9�M�q-���9��5F��(���B��Cj��iaM��*�M��(rz*�;������:�ʿRif��a�f}(�	�n���ߋn��.��o�s7�/h�9��'3�G�`DXn�ݕ~�wj�j���Ñ�:_55%��2w�o>:����q���R�)Tf��1|�,3����Gԗ���3y�ϓ�?�^ɰ���:[�5#?J��S�9la֚��6C����R�؍�V<�t�P�X���N w�3�>��W3�Sm�Q^B�8�x�f�물�/M[\]p�w9Wc��,���Z�9�L���9]<@{m�m=�����;�z:�@������1���9�v=���1ǈ��ku����):5K�8�;����sM�UJ��畷�7.^ק��`���L�v���6"#�îl4�hE���ڷp�Q��ћ@O�RJ(k'm���YȢo_!��=L�O��Oj䄪Q�F�'��'�휻5�ˮsqY��>=4����R�t��)���:�		H�4T�I�EI�j5�2�e9�L-Df6uw]Y\ϥ��v��Q
)fYn�������WF�nBp4�W�6�`�YΚ}N_[`N,�G�EUle��hWUn*���Ee�U��4��\�̊J.��I�Y�gc��8��M��L�
F��k*򭹣�dIR�d�4�����F�-mΩ�ઇU6٣b�_+���D��y�̷�z��t�8�{c�m�	�
�Cy՘���9&��K�~�/�;���R�����,c���#�������3h���[Xe���ev���ڲ���z�9Ο��e�}�[�s+���q��ᝤ�%bf[���g����*f�y����燂�O/]�P��}J|J�u�lo	�����_-�s��XS�d�s��-�Xb�?1n�7�ج�:�B�_9�x�m^*��5����5���]UM��hYJ�Y�x.d<�(VΞ靀܄>�Ujׯ:8��*V0��n'�ב�PyCE*��a���J�]����9\
���B�׈�i��t.���#.���xX:������u������J��@�1�-�a���؞0�t�3�/.%u��\�U�6���7	-j;J��c/������h��tY֮��+\����"1��w���^wsb����.S;r�s��݂���2fs*7��N9�(M���VnU��P<���8��=�b�h��;���uNe���ɿjJ���V�Ŏ�<�5��y��Y�c��v�<��ͻ�R4�s�Ro(��m^�<+T���;�<�"f$S6�����8��>��.�D�9a���l墷�p��B�;).}��i8�}���r�*�WYN�P$r���N��>f�*�zw�F��,Qɦ�CA�$V�����OƮ�F*wb���p�l7��5մ�>ކ�ZZ�ܢ5T�	�fk �E��q�%�9���� z�����!>+.WU��jjK�-�,��}8��/ް�Fy�wj��M��_R�DL͎�j�@�D�{2������b������/F*͚=�k�o���2�s�窱X�J�WY%�Y��9�!�z����-Mqy&w��]�2�ezG	Qr�zM�U2zGfN�:�I��s�#+��w�[.s�.��b���DF������L!�ı>��arjƮ�@�IXt���X�et=F����R�n�H�m�n�E�����f㵆�f $�ߋ���2�6<8�����`�yo����z����:�
[�������Q�Mŧ�
"��X�9�S�4�鰽Q�W$�l�������6'�籋Ȱo�҆��݂뚽/��bq�ۍ��\����ї8-�!!���<��y�5��[u��Ddl#Я/�9����m�Z��<c����F�jZ&;T�)�D�]�ќ�kI��)��V���g$����o�z���S�����K��Y���4�g<[�
\���	���]
�N)��7/�:�����(t��9�pe"3��a5Bn(X�r�$�9�^_A	��w(h\�����7�c���M��7.�S�U�L��[N.�a���T4c�Yoũ�YTr�#y�̜�
�����h$)bܭQ�WT'1��*��ŷT��0�\��iN�ų`�)�{f���Qc6��Gҕ���Ƴϻ�ᣢ��QѤ����`���~�x
�]d��if`� ��m�֤��|��B
(���k4�ӽ�{��8�WIp��)1g}�T���+Ns�nuluu$�7�p=
*vr7z[W�^Q
��!w�{+M>&Kx5�p��7����SY�C��}J���,�e�	*<۽��g�f�[;uf܋6��\������)D�ѭ����t	
��wU�e���T����®t��1vP)%zh�v�tޖ-L����GʻV�&_^�=�/�J���3]Z0�\�P�[�
}x�茎�y3��P�ǅ3΂�ٺ��#���p���|�:50���«C�βv�v�:eNrޭUьƘ�l�[ȱ]�r�H����:)���fn����"i�v�w�#J<�(���[{x���$]W���|~.gV0�����x6�%�;G�I�7҆bwբAe�]���繵�ȝ�@��:���Q�+G�9�Q��u.T��4�I�����lx������ǰ�u_`t���d\��_4 �������Zy,P�5�j�#آ=X��I�����[O:.b��������F��u1�G�k�jc�u�ϭp���!������أ��犧7.���v^I�p�=j��M��2�ݫ�o=�C^=MZV���|NF��u�Ȓ�p�X+)ؔ(`�.�%�;\$�ٳˎ�,��H>�5fN�3�tt�X27u���8oo.�Vos�Ƹ���N�6�{Om
��w87206�+[(�2�4-�)Tl��uW���6�]�Q���k��R����I���F��rd���kMN�o.�WH�rqS�֒/`qЩr�R&�5o���Y�81U��ٙ�#���3|J'"՞��ރ�ץ���/u!ߺ�5b����a5)`l�6E5Y�3�K���ܣ7����fn���qK�ޤ��#U���.�X�c�M�`�i�\$d�rkIcL��f3v+;�J��v��=��E]W7q|��Q��Ts��S ��!ں��[���:�F��YPT�G�9{��ZZt���ڮ�M�x�e�ח�R3����q���w;��{pq��%w+L,�2��?ҏ�90��+@Ȁe�g	�2��*����q�hL�j]���=ӽh��v���4�;Rس���Z;>9ҋ���~�$P	Tѓ�����oz���5��p�8{��giV�)f8z��b��{��_\�&��s���Q�%�U�ݞW�"�V���AZ\�C��^z����g[�*�#mE��T[j����q����������UU��֪��DE�T1F�X��̴`����(�5h�X(,�VE�"+ڰF*1b��b�,cb����V(�#����FbPTDEA-*�Q�nZ���(�#hQUԦ��1PQ���j�b��F,q�R�*�[�c�X�EQ*Q��(��R*��YV"$XŘ��UA`���A������Eb��5�"Ŋ�Lj�2�J[�R�e�F1-��EĪ���QX�ص�b-J��2�(5!TGMTQU���f5D�^����W�4�>q�svbʾ�|���,b��C��G1	d�]�"��p���u�l��d�<��w��<<4���)�ۿ�nP�4��yq�Vc����$0J�|�²�i55Own�Nc��R�^�P��K���r��F;[��l&v� �X�N2R��3�|2��E�˦�f�u�5�R���8�Vvfo�ה]w0�Qޠ�O�'�j�B'��2h#�v���s��~��|�9-�5|ȕ�Ƶ�r�<�e�\�wr���#օc�s�-�v!ܢ#"|4f���M(����NIA���䑎���/��o����ܧ�5r����Hhl*���X;y�]��{���+�՗�@OV>�ԠHJ!짞���r���C5̸n�Ćcz�ܕ�=������K�Ɓ�xf�؇�꜀�d`nčT$l��"x2V�2�T37�4��g���>�����+��M�o�9�Z"�Yt�U�U�5äW^�,�#�X��Ƴ2�#1�խti�n��3����uu�\�-�:���79c;�>�Ffl��soC�Z���i^2[ob�[�����W#$~�V��߶�;���ks�Prv'�m��8�sN�n�.Al^ɤ9"���ЧFtK��yVܦ��'1���x8��ٮ2�����9`��r}����ኄ�jU���Z�p�]k��=Z�L�5����� ���޷%�N7���'��ГzUҒzȺOw��(�->�{*�^�	i�6.���V42���T��������c��q'�`�=اz��~��+3h����`��x��lҔ6t�������$Αz�W�q�.s�p'���$PyCE*�t�x�q!Y=�N���ڴ��e��f��_I���b��^���QBތ��pt�妯�x�M+һP���X���)��е�kfcdŇ�U�Şk���jϭ��E�W�Z������n�I]bC�'��i�d�ګ���ԅ�hs���������{�Rl�ᷓ�����v.�!=�22%m�h�u6wn�:Fm��r������~���+FB�����j:��p�>�cY+�O���"����6���~�oE�u��/U-s�7�S�W�ٓ���2�Mc�[��}��_��O��Ӏw�*��-�+��@RA]�݌���m�����Us������*�� �&ގ�]$2�mUWv�(�wEn��D�K�)ء����	�����.(�WE�]U���~ѵB�v��rE{M�U-W���x�ZZ1����M>���k�
�2��:J$%�t�Q�S�#��ܲꣳ��(G�6���.�J��oz���H+.sZ�t�I�ygZ��~$7���>u2R���X}��ڣM���u@�S\oU���_<�p�ǳ5�'���X>u��1o -�0�u֬�	�wU��Л�э�a���KR�M���67]��w]n��9�����;WT���9τB4n��$�ͮ<�E�BȊv�j�"�N�M���\׬+;��Dۅ��y�u%XaGFWe�ū�7��9&0��oy����窱_t,R�8ʺ�1��qWfiخ���\�n�|.�����aA������͉�V�E�Գ���yJ�.w;�FW"V�2�s���[:u�N�+'��t���u(Mf׌���j�B�&�r���GFͬM��g!J��q>ѹBxlp)M>�u�^��P���Ks{�%��՘옵�=hS��Gz�^O`���W�0dr����V�]0����|d��>��im#U�%�93`[���꺪��gS+Y	�+�P����*W��Hhja�k�'�?}�	3�#Wu�.f__'cBp'��a�4�.S
�T����󑝒�g�r�:v��i�9>��Q�*�]h�,���o�]e�AE��N��͘�]Y�Xe�Gp�]�a�W:���Ѽ��ڭ_rw�����n#32s��]�򠋩1�֨je8�?R��ޮ|�����,й�E�@EFNk���.����rub�u;
��ڐ��4p�1�9�M�N(�،5M�Չ���\m�x%SZP3�^Xn�SE�De7��v/��5,��k[�BZ�5�r��hUC���������C��}��5մ���P=�:�پGj���M�����uBWti|�M����w�؄�<�yq��u�Z8��y�E'>��H�����d�en�C+�W���R��z������щz:�"��b�0B��N2[��r��U�E�˦�����%���6�w6���ls]K66�Ά�N!@�P3>i�X��B�U�GA��d�D#}��a[����m�D���z^ׄ�z���OUY�Mt���M��<�Q�sh��Q�dHћS��N��k 5���7�e^y���v�$���{:��M.��;KǳUd
�t�;�s���1f�ð��O��.:�3��5|��B)��%w�����8�� t�9��:4P�*Wc$�8
�溜�F�KM��0�*F�}�5�=��?s�u���S�ѝ	T�"7�3X\��;��1��%θ�ej8^��]ά�|����JP/�u�Mڄ�����L��D��s#Wu�.}//�[݂]*��]�����Y�`��k����M��Fs.�Ѽ7��&Zz������w�t����u�&�ʼ��@{�p��9��P���+[i�l9"�����V��o���4�n����;�;2X�3k^�oC��H墀]�$j��
��1C�=��J���ő�rkX��7���8�GlOZ�7���T.(�5U٠�\��}��R��sK�]�����;�Ns��xM�E3��]����Ots��T�f'��`M��
ʢ�x�w���r���3) x{~��^�ވ&�Θv�m��GR�YV���	��ƙ��{�{`s ��A{�x�b����5�r�z��ɕ��[c:oFP������Iܠ�� ɢ�l}۬���zv���R��lv�:�q��Mv��EX��,�X*Ͻ㋍�JSX���V%B�.��5��[q�y�=�7�>��t8�^ϵ�}�Z�n�����u���{I�e��0��Z�􌺐���y�V��L �u���j��:�x�pmc�}��66;2��(���u���4dp w"�+qzۄ������dD�z��ؾIk�6�)��"�ރ�m���+\���̸]N6nq����(�k[�$'���#U��nv�m����MV.�J7��.��0V���͜��	JG�H֤m�G���Ôn�;4�'U����ص[�Z&_Zdg(�Q>[P{�=�G6�fu�nh�l鮞av�M���Ƙ������V�Z��P��v�����t�1��w��@���Y,�=@}|$}�-	��3���^�m��O�����1��p��K��x�3}7%���Kb�8�/2��&+��9����&L��m-��o'�VE	�剩��q=NuwVu���+{�|p��Kw��J%-�ӹ[�����%��xĩ��ؼ�\��(]�Ң.�޴4r7��꠵}���ªs*��3�O���n�v��Ad`ZG]�Y��B��c�<cٞ�"����fUͺ�o2g8���c��L�4�ԋx����7����������wV)F:Y�QX��z+nz��^6���<��A��k�fC�v>������,��2�Eñ���lc�9\�E�-��;-.���Q�y�D(���Q�����b��>��G�V�I+�]��g�Y}�S��hɋ���<7!���>ji�]sV4�J���[�ː��r4��W%FN����zQ�
����S𺻹�C�g��q޽�Hgil��w��!6���j>ۺSJ��d�:m�����{�K��	�+��gz��ȹi���rs@^֡��H�Ѯ�.V�JZ�ᜆǯ�����r�h��di���s+�jPf�R;���E�����uO����Uj�ӱ3qV�=4�=Dazk�]g?w����}]���>��]�5;�67��t���H��7ڻ��s�ǵ<�D�:�>Wйab��J�8�����qQ������i�����ӵ��''����lh���7<@�K:%�\w]�����.�9C	�dۊ�SZhΉw�M�jhʬ���m�a���w�4�.Qwwk!#ܰMjܭQ�P�j��7'4W[}���-aBvΨ���j��u�纾��2e��t�l�謳A�ق+3.��P��:�@�h��)�NNt~�/��y�������Y42���B���N��3WTS�|2�)��jo=�y�4��X+��@mZ�{xr�J�l-0�Wv֛�D֌ʎ�E�q�d��eL��z��xc��`f�r�Vh��h�U���{�+n8��^����i��{A(����'0^�P���J��5�,�ک�O!����kO.�]T�q:�)М��R�g+��*�&��s����l_jBek^��k�f�й�B�w��vi��R����Wj�gX���n8���[c�(nX�����()l-�õ�jRN��.y<�Ӝ�㹵l3+c#Fm�O�s��]�t<��1�{����_:g���G�r�8��	T��r�;[h�nK;�+���G`NuԴ{V�z�w:���Տ�d��īNN�k�1Y�g�0��VT�C�v�v�W8���W+scK9�	��c�)(�H�ʽ#\���M�KM���d_>Z��e�f�lW(��D�j's�:��&)�K�s��Qf�:�F��U�آ�OSA�9"���Ф�4�O�۸�	���"w'�wqn��\m���,4��`2em���Pʵ�
���������ͽe&#��7YaL����
|ST��q����3=��K' ��6�v���/���[) '�9�.u�H+��8�El�m��@��y8�6� �v�/7,�z�JPs�֬�N��uֺp酴7nд�
�ܤ��U����q�`oC�ۙp� *�3���f��*iz�#r��Wp�*�� PZ�p=צ�T�ChE�`��ľ#�nĵ.��O�Ko�ٗ��Z��aS�l�����-��+�N��wC�kp����<ՒT���i�O����a�EL75�T�!��q���uAE���Z��jP�ReHL.:WY��Xu�V�4�M�����k�u�«Gg.
⿑�����Y]����o(c�oA�
y�{�㽥�y��ֆ�����ǉ���`�
B�`}f�ݩ�[�R�J�-2G*t�m��\wS�u��Ѯ4�٩xmb,��xf
L�Ԫ�T�U�1>멝��7wf��];�O�Q�@}�����:��Gk5B��^XwRD��%�blE�YE��+�\Xm�m����}K�c��x��iXFJ��3AN�H��K�r@�D�5|!��j�V�d��!v�}W��.ڋn��P�����x�;w��){Z.�Pl�7R|�J=.d�F�f�9�G��a�9a\?/�쁝�5W�p���ہu9ö��넰2�b��GR�Ʈ�7EV�2��tPNon[ش[�Us�̫�q����H�ftA<롙�}�رR�w�;>�E�LUƵҷC�k[��SXG^nP�)��y�!x5��y���D0�+�U�C�+�7���S�Q���˵��؛����ʯu��;*�"�X{�ld�z�m2Rte��Y�[J��3z���)�u��k���i�R���.%jkNV�&�,`�#��Cl<�L���G���<u�2=�L4f�aM�w�]��ϳ���WC&n��6.��ԯ;�>���
�V@��c字�kԠ;�Le����fH�ļ��EImnEG����v{X��fX2��Ў_+�!�y��pC��9-�o�]�9L��i��)�j�<Syljںo�W�-��w�j@3���ק���3�nқ7�
))5Cp'g��n�Z��_-V��}� ���l�7�U�gW(X�3���[r��b𜗘��g7 io#��]��r�v���>���Ϥ/���O�Flp��Kկ�}��C�AX�g���[�Q��Vڙi&+
�-�[���UZ¢Ѭm����T����-�1�Rت[)Y��F��b�AX��1"0bR����r�" ��5��"���Q��,*TPh�DUZ�N&+��ũkU����-��h��h�f�,�r*���2��d�sF�r�(�m��(�,�,F�F,TE�˖�L�aq�E�"��"���T-���)q�5+b��Ed-(��ڬY1+��cPQJ�U��iֲ[bł�ŊEXQ�*[kh�)QDU`��acFءU�U�!m��
V�m���,�e�J0���YL�k#mm�PYR�ڵ#l1��a*"�VR�*�RT�a�@��1m����ZЩl�VV�J�j�F���B��ny:=7`�J2W���oW��ڇ�t��b�[�_Hd��%x��:�{��>�#Ǘ]�U�ӳ��r��m�[	E��9)�Q��L��W���R�:�k������%:���\��~�H���k�u�3�v����a#��"�;%o��-x�N>Br(l��tfS����o7xO��w����Rn&��:p�.I���?k��,�����U�YT[(���+3�+�V7�n��8�4�lw�F�4<�"-�8�b�=�&�Þ��$���$?k��"ی��	��P�J�'r�G�	�JL��NWsJ���OSl�y؂���P�G�]�����.I�}Q!��c�pMpҸ���qmc�}����F�S�l�>����X#���!oW�h�֣�����_��TY	8��^�3�3�Df�HK���V�i�Wb���(�iSb�>���{u0�偫�`�ss�k3w�fڦ��]-V;4�7o�g^&�=,����=�Gq�so��Φ.qΧ��fһ�ݲ��6�MdQ��0,���C�]�J8�uEn,�H.E��ϱ���${ڃ唖2��Ю��sJ���Sk��QM<=���S�)O�5�זͱ}7N�iwB��X���/Q��o<Z0��F�r�E�zM\g��'��Ȟ�n�I�4s��ѵ{���A�$P���"�j������	U�κ���R�DoCJ--
��C����۽)����a*�F�u�݊���^.��Ϸ�k\d>�E�{�.���w'UN�=��Y�v��r��J[4�B��M�n8����Wc�7�fz��Y����g��-7,�옖/g��$�>N��v��|�Y�����'�\�(6��E!���[܉D�`V����2��@�8��A���x̅;�T^���tymA{^�X��T��ۛ�1�Y���B˝�o�6�tx!�)���Og"���֩oL��c�'*��zv),*����Ώ�I-ܼ�@� �r�&�7��qǯ��ϥc!�D� J��Ӛ�!̢�E�rH;������[ԅ	x%E�,��Ň� ڷ~e��{x ���zz��ӽK�O��+�8:Σ8��ڻP�:��F�j�������yةM`�y�=³�mQ�j�s��{gC4gFa��lR<�1���|�Z�%�Z^��O(�"����ҵp��Y�Tu1���]�V�E�����<}����u��*�k�e�bV�	3�i��uekOmv���}�J�v6�c��ԇg��~� �!j����w�\����O'�@��ڙ�=��d��	����oJѝ�Mpk3qt��x\s[�!x���,hq:����
|[�
 c��N���s���`r��0�N�;�:��xˊ�����fuXWqd|���8lA�����R#2�I��Z�e�'U�����3��*v�MYQ�e՚A�r��P����x�|ʤ��6�ܾI�u5z����Y}�� ���{�Ι�U�s���չ�Ȥ�s���5����>�Br��O�S���s���;�:�T�'���ֱ��򙴺��oV�!�vv,���U�{����<�˕���]���P{���㮵��Vnmq$��O���n�!����X�ÙU��2��p����y;�u]㑸}�Q�^�/4���jVv���IQ}�::K0W���=�fv0:��sss��R͍.t7S��26a�Gc�m�m���Oi��)���[��;�hnP��<n.���q}͞'1o]s��dbqŵn�;�J�:L�����L��7��/}C�y�i���.���i}�x�W%*�����V�r��sl*�5]����o�S��{9�g-��^&pG�Bw�F�͸�ܩs*��A�)U�o�:�A�H���(|��c�CE��&w.�b�_\ˬ�9ҭ��c�2mwR=ӆ#���9*v��aB��Z��U���)N^E�op;���f�O$�o,�;R����Czg!��z�cdj��q�pd�uCDÊ�����ŉYj�YA8	A��������a�*�N�7��X���z]��"_[pG(��U�?j��v�@��[��'<�I|:ო��}��z��$P�s^Ф:Pu��P��������}Xf�����B�Q<�.�85T��s#�4���h�~B�[飗o��G�����ε�`��5�wm�R��]��Ku�kG,�U�r	V}t���0��7��X�ֵ�.�k��XW��M�J��܌��?z�TM+�ת�Ǩ�+0osC��]<��n3uF�}��{H��x�عӭ�m�ɢu�9=��n�
�C\U�˜��	���Hw�)g�0�zJm{i�s��V���U�]tyq=�x�ha	������J�s�+H�G�)�z(�-��yۼ"�����G[GUu�/��rpљ�sD\�lr����"�%ȭ��2-��8!�e�ͤuD�����������9C撽���Zm��Y����U�+n�u�Ҕ\�P/u�vk���R��@��q�j�}n�c0j{�
UUo��F��2����-�Z��GwU��b�@���a`s�Gђ7�-	��z+Z�/T����Ɂ�g%�4������7��ƮR�K�� �L��K�ӌq�6n�_5U�WZ��t��M<=���S�)H���zȭ3���t�ѯ��ȃˆv�y��2��#9@�r��,.����e�n>,.�NvA�8�8�6��v���^8&�ur�j%-R�����"��ib�X[��8U��7����ӹ1�����s(�SC�΋��Uܝo˔>�ۍ�7�+�&�Ǥ�9��C�;C��|�E*U����0Т�E�W7}'m�讙�Bኼ:�r����H��<�X1�ΉC��J�+�7��ԥv^���ٰn��9��)i:�n�bw��=L�|�`�U�l�[ܣ�qwb���$�@.ܓ��hU\2b�/�Ǆ�@����$�oOnLo�Ƿ�iőz-+�6�ƹb�{(%����{|�V&��5>�k	�"��b���X�u��}Uc�!��z�}52���ÝG��*�$��]��<�A����w��7̋i���o����	�n�oP��Ŵ/�6��[����'jJ��9����(nX�� k:��ͫ��:#�hgJ��u���{;�t�؇�ElO�nB~��}š;��u�gL7�J�Cw�!>�p�P���Jo�!uZ�cA�RV>U�f=2�t�skf��uO=�t��w"_&�#6cj��Z���]����S�Z��B�ۮ���� S��U�^6��֫�����8驑/���t���;�:�t)|���Y�r҆hX��@��si�5d��s;��K7�h8:�]�}��u�m��9�,ug+gEC\%vb��ؔ����ͻ91{%�}�G�_ �$@����z��cdj��cJ��q5G3���;���5;>�nS8�l��DgC-�!�%B��ƒ\ƮS$P�sZN�#o���ܜ��\��^V­��E]ݨ�䡆�d9�^#ve:RǑw=�nd��i	ɶ���b���do1C��X&��rH���G�Q�N�_�#���%�7u���u!~�ֶ��$vh��%�O\Ec�zU,cL1`�S��ӌ�e��4�[�xk+^7�9�Wi��v�]m���G�5~�9�w���[5=3���nK��8�*����5���#���J��7`R�g/�Φ�3��Z1�,�cq�q�y��R��B�Cu8�x�?�ծ.�lTڀ���"��Gl�דy#c.}��	Z@�-<G2Bt�S���V��0<���6��ǖ�X��j�<�M�k�qXy��;��9�YK�e��_^�Qu�����a�I5��w�=7O:p�V��;�1�$ �'u��:�ϫ<��{����o)�������������.WW@R���������,�8��a�����R��y=�u�����FT���ʁ��|��������Ʈ^�ճ��dfɾ�͇�w1�3� _�ZSʄ�@���겻�Y}��Tl�vS�ҝ35٩	;��w$�8��z�VCU`C՘٪"`N��]��]��R�+/��	���G+5Б�}Oj��r�R��q�檸��WbE�����lW(��'U4�ب�l�0OZ���2t�U3�D��9	��H��潡?G(k�Ч)�����գw9}N��N�^]�0ňzDNm�U�؅2�*��|�v��*�98�{a�r���g�١��S��ՏI2n�k^4�+;=��,��{����uy⫪ k���rg��y)/!2���=����k��)���PK�97�N��1|(2z���osnd53y�չ�X@ݷE��GS�ժ�|�iތ���Vr%���Q8P�'0���U�����پ��=xVtW���X�-�e_����$`�\�*�*�lu\���\\1��z+Km(2-��sz����x�*��"t<���-��UN(�����s����y1'���E��f���yAቱ,[���D����kU1)��@�SM+�L�,�{��*��%1�Y;M���?O<�%>�,2Ԅ�xV�=i5�J�5�Ƹ��rf�u#�������O+�6'�41�����խ]��l���Էi��Uoc�a�����r�d���'S�u��,Уnc׋&�ּI��<�}�S�)�,hΥ�{P|��D�u2ԇE�9Zz�=F��ew]YN�����S�!)��༤$m*�
�����Qwgt��3�;���� [��V�0(�ӹka�oRRtW��6�-ǻ��ʼ7Z�r� ��ָ�X��{S�!�n�M��_^2��5�^`'�G���Q25{0�{��-+�����6�)� ����Q���Խcr���>N.O)d[�6C�v��Ժ{�I��JT��Z���ι��Pۜ:�HjI��i���M���7�NU�/�g].�v��ʴ��}��1[�La]�[�8���Y]jC����l9[Mkr��M���R��Y�sl:V���>U!�Z��U2w4�[���;���&���,��Gu8
[6���9oaY-m^X	%Mؔ�QR��cua;��)0H�j�� �p�5;�Y��`7�`���ʲA�������>���c�T���W�F�d�7�Υ&��F�>J�����h1�h� ˷Xe��yȃ2=��Pˡ�Z�[�f��9��*�z��QT��c�-)�s��K	�E�mi{	�u�1@%��+q��X��f5��@�u������J���yՔWz����z��ʭ_"�ʵ�+�/z��*�K�:�6�`N�\
���x�B8��N�\����`������5+�ܳB��w�q[�c[�\N7��z���]��kk�h�xݰ"��4�u�
�r��Gd�b���
fb	���ü���ƺ�J�)�Ь�v::�b�8q�>Ё�%��X�����.�A���[ƍW:돭nܲe=����j�ǹ*oL�Y�u_	��[�8���J�^�}Kr5��ѹ���T��m� K�ԧ�Wen���%���P�r�������"��uw�R&��涴S�~�=[nt�k)f��kViU|����3����4�Jso��D��N������v���Q*������Y��Ktvv��Vc�"�}���񂩤���Y�J��%m�V��g8UX�V��Z�QRn�=�J�
�3���-ֈ��F�j�q��W9b�� Ԙ�(��񾧳��-�a�ϷMYWV��Jֈ�P�ʉ���6�Z������T�JP�/���][c���_��>�P��rA�D�m��9"�"��
��`ɐ�-��&�]Dv�5�w���0�;N������D������R��U�}n&�!�of�7z�\!8�:���x���Bь��<9�:w_k��Z
��=�p�v����ˮ<�:tK��ݜW<�������[��Ɣ��B��5B6�t�C�W� ����*
E�J��V(,R)Z#l��1	�4�Pr�dkcl+U%jTcR�b�,DE��P�AH,Z���*Th�U���B�#h�J5�ƣ���d�V
�m��ذmA��-,��m���VE�
ܥc�R�U�Z�f.P\[AJ�fQpTUXTeˌ���e��jJ�&10j�e�5B��Q`,3B�*���j
B��[,�V
�Q�[&��Q���t�����T�����ej���Q)b��iZ\�d��-�,q�1���F�Qm�Z�����,�-��,QkPFض�¶�\n �-k
�6�ŭ�V�bVX�ʉ�Lb�4�*!R�mb����pʂ�J�W0̑�m��Im�Jܦ3,�!PRc1��jc"��&%I��V&\eE1�aYm��[F�VF"�UAL�+��.��)DY��j�R��E��`�IPշ}j-\x���w!|�i�%����Y&���>�Bd�RU�v�є�vwujo&9����Q���&��Os���ά[BŴs������N�P4���kW	C^T���N)���W����h1���;��6�����`#��\Jł�KsG
�t�oC7��PGMm"w�9C�a���G]Mp�����U�ڧ*�9�L�V�5KW5F߱�C<VE.ܓ�΅7�&.ړ�*{��~��o����Q�Beּ��K��ɞbl,���v�=]��R�ڹ\y��y�ZY�F�Gyi	����}T}ae..�-�Y/2�;�1Bi��qu�np;|���U����f��`+;.)����M�����O�9�	u�nw�\�-��M�Ȁ���nhέq{�����/r��[(n@nġY�g(>mN�S�(�2�������O�����Ӹ�+�U���<�
|��sL�U�,�&�pd���0�
�/��E�2���:w�f=K��{(�{w�Ti��-�c�cxk]�����;�x��u}q��pIe�w!U��[�V�c���[�r�����v�.*Ҍ�-�Ws�Σ�Rnƕ�jX�j|W%�������\3���k��	�Z�()a�γ��6�kf��;�x���d�������!�3=���@KD��YOt
��VV���5���n�	OG]=�%�W��_���ѭ���Q������s�kw^�9]����HU�[��~B,oT�}!ߎ*����<�L�̱
�#k����7P�.H��潡F�#Oe �$_d�sC�|�;r�F������[A����{B�ѝSO�"����r����e����B�!ܨ�45���͆���/"����߾�²�;;��u)�F13�؆{��&��O)�U%��
T-��{��uwnt�#�|A�����V��:��=�Pb�b�X̴���[������a���me��G�
�N�bO���,�f��8�۩w�*��3'bӶ	�x�j\$�n�:�<�w#���[PR��Nyb�Q<��R�i<���<E���YՈ�Z��"���u8<�*��]P-��+TQ���\�斡���7�����O�;�h{�8hS�
�r��C�
nxI�ǥ�˦˜��溕�ؚ���8u�1R/z,YNW3Ɠ�Os�ܮdj�ۍ<�nV��"�I�����:k�iL���b{U� ]&}��}�#�>m[��T���j\�Y�:�8Hm�`�cT�G�����u��ܧ�g]�����D�������]��z���e=T�]P�k�u1���ljE���}�@J�.� ���ʖ��=D���*"շu95�;�I4ŵ�VW8x{|�'҉9T�u#o��S��LmtozG���:��D��щ�K��ԛ��� �W�-��d�Z�ĈV��דr���nuwS	�Wib�pѴv��ۉ�Ѻ���`Y��'=ܢ���P�.�N�o|̭����p�A4�3'UV�wOQ:s�+Y��kpd��e�M/��lW�D�Q��j9��ܶ�,���n�I��#��z���s0TKDKF���%r�a�q;}��(Zs@隶�ބ���h�}
���7��wjZU::x[�6�����-�Gu!�=R%N��/iƺ�y��oC
�a��d�D�u^��	�*^ J���V�a�n�hg+(�C͕�Wϲ�دj���a��K+(*ۦR�p��4;l�.�Nk�c}yl�S��hyx*ҋ��;9��d�.tx�N���k8H<���_�l�9ٸ��y�&+��QR��e	�)МU��Xi���e�ۋ���[�n.����'��W��#��N�-��jƕ�j�I_cʵS�)���a"��{�w�����c�a'Tcϛ�C.�B}������z��ƙ6�S��g�v����--l��L+ܳ����+�1�(gd��#��d����U�iV�����[��&�Ù�f�OC����E:�s�˕�9���~��,�V�T�/�`�+�o��֣{�'����Edqwܘ���CDkQ�c�!+�Dd��Ϛ�q�	 �'J�F��n�Q�W\�,R��!=�q���.�j���랋]�"�f�UP�6y�]Ʃ>Vu���|��GtD/�ܝo:�e��Xc9PgX������o -/��cR�����.�(]�V@}�>��	�f��SGѳ��۴����t�p���V�K��ɶ>U֫�䮲Anh�Tq��8r]Bf�K7������#ӹDk��E�4��W�j��Z����"pc�ę�;[+�@�dX�$�Q���\2�]��q�*�nR����QΚ�����QtZ� ��f�)�+�e�N/��;'aݾ�6ݩD+fvYԑ"��{V��6��pt�`�k 8P��j=|@j.8]av�e���!�ܘvC�]��9z�����
gM[�Lt��:8의�rLR���Z�'��&��J�W#�����]����p����ZBef�;Uy��z�;�-��̗��	DN18����3�����\�kqx���q�:�]��2��Gk^lM�s�8�Qs�;2�޹c����>�xfj��\�e��k�-��$7R��q��;�*DB��nk��`���k���>�^7�yؔ���	XkX�y"&��7�#׏^�t�^��jC�-�Ư��A��^��G��Wޞ��?p�Yj��ΰzۦ�^kf�T�uO_l:jmE��n�<���r1*�����^�Wn��
�B{�{)�=�y�fu�Y�v����9�F���`�ή�]��!8+�7�]nVZ�a8!��H����X�^���umԋ�3P+u�%�s$9W�y ����g������,�����A"5	ʾ�v������5gsЯ�Q�+����%�oqe��oMm,�S`�p��˸U5�Ap���7ev��ZzNj�
�F,�����q���n(j3�Ghr"v�B�\�>��a�Y���{7�o3�݄�|A�7���B��(���U�������x�;<���:���*r�ѐ��xq���S��/�Vu���JZ�?{�*����u[�;��Q�J�;ؒ��[����b�1F�ew�/a����eW)�Y!)�9i�uc���w�z���WK���
���AWL��օ�-���/HoV�k��/"x;�*�)���ai����w�!���u�z�n[�77���3bh\�n�p�u@�f�c���.0���dj��9�W�[��tAۗk:���B�b��(HZ�H�hev��#�!�m�J�n+sqǮ����\�/t�kJ暴=4Z�֟�M@B}�I���͆a���E�t�p[6�����s[���F����q0�X��`��5"�����I�:��^��=�3��Y� 0lb��X2��FWZ����B�.�
����І߄�|�ǚ>��v]����Xgz�OHՍ��rm�ے;�DF�%����ڮ�+����l�ɵ��6N�%�7��������e	h��!������Uj|꺩��ڻ�p+����x��F�U#^̇�.����ܦ4k�d�.#R9̻�h�K�v��(�r����{3N�n�|�B�'6�&v*����>ΊnӐ��$_´�^5x�w�
S/�nۚV��*ۚLնϷ�
J*�Fz{g(��2�+8=ܹJgW%�|���qI��y�w����q�!{D>q.�p�Y;�����®���k�+��ґ��o�su][���%m8��E�qy�-V�{�>޽�]g"�_�6K�L �\�5�)�3i�Ԇ�[��ܲ��� �d�Y�q��@��C/���π�ٜ�|�_L����[��Y=:�ot�4��ħZ�=m�b����l��UFY���V���1�*w25�p
9�:��}Aj~5
���u]�ȝ+aA��Y���z�:�v$����}�qV�e�vjy;��� �v7^&
���`N:;�g)������Zm�n��>����Mb:;���#�2�7���'dR֓]�+��3ۤ��+����l^�o��m/�Y��Jc��X%y�[�w�K�T�;͠h����	kQ�>��Q�f�O��{+�P��jǛS���f/x�z��r[�Oa[�=м�{f����7Q���Zcr��u�=C���n�q�:O/���N�ټ��ٝ�k%k2Fh� �!�X����oFc	E��8���y�8�W;�|���l�Y^�����hڽ��sA�u�etL�(��T�i�����С�dR�"L�!w�Ѵ���� ����[��n���p�=Ს���^� �/��#[�0W�wW-Ξ��|`庛B^�	QZ�
���E��%mLŸ�������j���j��,�Qcb��4�]d��p����i����(��cm�BZ-f��(FX�xi�(�eM�gm���vc���.���c��q�v�j3Zpͣ�;.�Oc��c1�w�y���^Oj�f�m8��-5K�U6�Y��㘷:��E�m��B�-�u9�ͺ�O�2���FoiL�Ԭɠ�^��K8c�Rfg��t�5������R���C�)�Ԛ��7igy!R�������ؚ�(�okz�s��v�<�����F�lv�N��e�v_���>���C+;�!�ou�UN�ڲ7��v��Ս]Z�d&�r����Q[8nP�6�j�#\t�!�H��"뒽;�3� %֮�1��#�����x���D�R�PUU�A�H BcO���$ ���#� źSф�=��f��/�{������']�؛�b?�3�5�xjCL�		!�̅��
���P�Ɇ�3ȅB�+8�{�]%Q � b3��M�6a\���<�����"gd��?�B?��3E����I�~�<�2gᇲ��ϸ��<��@p����y[ۂ� � ��>��"�\WD�@0-��E@~ax�#��!%hu���s"Cp�?��CҤ�<�@�}�m^��F$����u=����:�H �ƪP/"��S�B����ưҡT#B�%JB$��\=�,�5״��9%�*=�`�-D�R@� �OOӢ��}�����jt�#�n�����V�D�
�%�@�W��b�l*��?b����R�&���v]����w�jI����.��j�k���u�+�CIq��=�����_���&\F@k�2��(��)�c���y!��B��'���$��T���d��ȶ�ǋTصS�����3
d�6����to5��C���0���0���eT����P�p���C2%ـ�0�G� �����B?S�I"m(7h=�!���у� &eU�%�� 	;��qX �dɃ��D?�zO�� FR��F�!i�,��|f�"�jJ��	�M��'}�{���$Ț��K�1�?�S�D GKpv��Gy�&�7� 1pGC���Z��a=~C��F��B|GHC�C�
 ��Cj�]#�
��'V!���	�H4�Mj]�ے`~~�U�7eu�#b��Bd�^]��0H� �2��v1�C����6!���Қ���C1;��҅�Ն����
)H�!�́������e`�榒�#/i���i�s�s�
 #n�%�v�s��Ɂu�$�C��4��Md9_�ӷ�\���U��
B* #��h�� ��h� ��u�������	5�d\B���D9ҕ,&i�
B�J',L�q����w$S�	�� �