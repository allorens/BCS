BZh91AY&SYQ� �ߔpyg����߰����  `^���@(�*�!�}= P   _�z��s�R�)�   ;{�^pm@2h���G�J*����Q@�{3U�4 � =9 � �l`䓅�� ��  �P�m�p �
��� n���6� 2��G��{��         @ T��4�UR�F�0����bdaL��~��*Q@ �     Oh�%5H` F   �  j~��jJ�	��&FL ��0 A 	��4&�mQ�zF�ѓ'���ɴ�"OJ�$z�h�@  7_tww��o���y�҂���)���T4Q� C����2����6T1�����~_��ݓ���������4dP,�j~2�1U����E@P�I�"s�K������"Ȁ�s�z�Qt|x�����K���o�ϖ�����/�-�F:oe�&�P�2D�9Q�zE���I�ӣ��FM�,�<��2$��q7ḜM���'Q��gg�}�3����n��`�e��,�]ɝ������Z�.E>���y,��ivœr2�l�8�3����U�>�:��xP�6��������/��j��N���"�}9��x�����M�F�{��D}̗:S5�S*��)�t��TD�o*�<�܎D���D<��,�eQ��,����=�7qDr#��T�Ȗ����tͲ���A="f�N2M �H7�r#qD�0�,�����U�d1�N�BT��y)��JD�v$�+V=8;#8p� �%�f����r��7�Np��`�xd���<X���E�7�zg
ȍ���]U��jԭ��u��j�Exr�&�'�����I0ò'�'G�M�L�a5���nRm�I��#Ȉ���t4�A��Q�C/�����,�7mU�ٶx�'$�{��εZ�:q�/%�*�f	�L��U��^x�Dj`����M`9�������n6�����<���[�޷�VhhXii�p�6�ҕ������=�a������!o[ۡޗ�p�n���<>:�2L�&k5z�BS	�Ih�6m�/��Y��6�"p�0�3i���ãD�Y�va�e��-�D˗z�:�I��()�������	��S�լ���ǩ��?���PXhh2	r#:WE�"]D�%v%1)�zj{�w�oOE�d;e�z^��Y׬�C�z����v	�c�J���ȸ�*�vm���t��Y��n�U�q��/[�u�LZ/-0��f,��-�!�3T�>����V���x�'��f�+5��&,��
�kSL�"70{���V��:})+̬�+����%�zm��c+�9�T%���z�޾�����z��7�І<&Ұ���oz]��Z_�����҂�w	��Y,P�w|l&���QY�VE"H�o�B�.�_�9�'|PGђz%{��Q��"�w�u��9qnO��"��=*a��_ļ1w����8��dƧ������^B���΢�#%\&��xp���3�܅������a�;mSq���{+�8�ׄ��k_�+��P��qc��d�3"�^�:��VIEdz�����fZ��S<ME��0�{�L<o"�t��;P˅�QU��������ܯ{/^[Y@>���$e��>4�6���4��G�V�,s�Fw�7ݚY�t�כR��4�]����x�<x�/������J�t ��F�c�͓h,��z����7!Ѵ�k�#��(nˬ�t��~����QE�*0<@ٗ���ZR�=�J]l�o�Fi�.��(�L-���*�ջʑ��U��N=p�I��T��V��*�<��Iڌ�}��A�Ia����2�,�&\k��[��<t�Θ�%�Y^��M4��~OOX��4�(��4��r�+�����=$�Pܒɷ����L�<l|â�s��Κz�Qŝ��|P�*5���<B�c��dz:���0'_z�^����:P� ��]w�ce?���,��Y�����e���U3�]����^zV7�kҀc:iҍ������:� ��ýi�g@��>�C����/D�Pm���<`R�۬*4+��[u��rv8e����ʝ]x��*lT�P�Y:>�M%g���y<�鑯W�Ts��v��\�]~ h�6x�]o��
:�3ӾZ�]�Y��Ǆ�J�4��xe�3�U���@0�vHx����Q�މWSP��xe�e�@t4��<x�V�<��(�! �����:Qf�=mt�Q����e#�ϛ��n Re\���Ww�vmd�0(�R�4��Q�O��B�Y��:޷#�"t�T�Hs�Y�nd�4�q �����fW����-(�G�}��IYget!���t��>!������Lo'|�����/*h� I��'�Yvdϰov�f�j����t����}�s݇�}���6�����×Mǉ�H�4M���^����V�AKك�FN�C�q�C]=�a�L�1hNc÷	�]gX�B��� ̮t����k�a�k<dMgXN�i��W���!w�`s�W�@V��h3 C�5��*�F�mg�4�uÈ-1ǖIj��g�c\#BM�,V'1�k�Ţj�-ʤ�ק4���s���&U����T$�`�>W�ۂɮ-$1:��Mb3q���i�cFuD;bƋe���< ��D��~9��Ѯ�� ��*8�UH
>Fޅ|�C�Dj45!�*�����|�8��E�odL��8�����v�[n�(��.|Έ��t�y/��jA��{<�~���>�����t�]XƧ��;!�����?���1UU�UqiZ�V*���^>f�Sp��9d�*7��߼�������+UJ���"���� IR��nn��|�7U5U�/�����*�����T��Uz�UW��拕q�sJfV�2R8�1 Ђ�^���U_,UZ_"�U����V�U��\I�M7�*%)��K�t�0ы��W����U괪�,V����mU�W��4BjM
�jCD��	�J祚�F�o�1��^*���Wj�Ջ�{�Uz��W��[��&-$���0DU1�x�;�mUx�j���V���UUťUz��P4n�Mj��U*k��8 �� ���%�Lc������U�U^*ڮ������*�����։4�$�$��1%qfsb*0��q��g!�D�̔�b��GWOj�"���I��������t���x�!D>C�Ģ��l��@D��"�AD�6%�,bp��8N	�:!�'����"x�ӂpJ����q���훆�RL�o�IJ�$�B�A�Ö[u���"��hWFլ�$�j�:�N��V�mYT�X�*Ơ5[�q(���UKP�rJ�S�Z�P��H�5en�*D���V
�ӄZ�`�j'ƤiÒVX宜�NG�&��9*o���ځ��
 �*�V�N q��'Y���ڱ���jRd��0i¢��`�cE(�m�EV��t'T�q��"��CT�p�BQ:RVZ�H�r�I[D�
�d�jD��Bʔ�+B��uK�� J0ebn��#=إ��ӑ����[Ƃx,x�Mik�μ�2�얣��DW88��
Eb�EF��-�QâY�N�!�TV�v��c�)Gk���k�^����B���TU��M9�A6���� �,�li��5���$�M��VQ:�!��֘��u��*d�Ɛ4�D�5h���I�$��	 ��u��U]��%�+Qґ�V6�t���N�V�+n��*�����[cBT�u�J�&�e�1�%T�펫"n�&�A����	Km���ӥ�P��EP;�7��2q��
[)-B�p��D&���Zr&*�8Ȭ/"%N�'A
 P������s3331%�����$��ffff�@ffffh5�����F������9�s��I�	:t�����Ui�3)���z.�=���j�4&
�K1Hy�m=�t�rյ����r�V��fD=8Oʪ�x^�ƍ��3����aur�=H3X��b�\b�g�=���7Q�C6�|���v�I���]�u�F�i�<�\K]�@��7N&���P�`:4��V�?�����e}�v���E�yuJ�	P�<8];?*E��Ęo<��c������6�p���B)������^��R��j�+N/�up�T�EI����ч*�n�>81A��[����S�߆�{�GҎ���5Z�Q�e8v�� ���2J$�Q��b���qͶ��"�����Χ��;ܠ���WIM�D��fO4QUW�*�H��2fn>lY5�@xj���D/�9�j+$���I�y�_�|�Ƣ�����m���O���:�g3���V{r�6�?+�_'+���IaE���[��5���u�j꒩}���DI���\)=��.ir�N#��w�IFp(�uI�b��-[c��O�-���|	G�Ƭ�}���]��b��i�q��MY�h��0�N�XQϔ�b_'��>g�o���|�E�P�K+���ZԋE|���&���AAG,��]�U9�w�LbК���.���o��4��Β��5+$f��x7ɫ��!8�K"�
z�F+0X}���I#��e
��m�n";V@*Qjj���e�sNYH��-�s4����JT�҈���n�D�J,��Q��J���;m��<�����$@�6|C8B�l�=��iDi�IӦ�C4�i���3Hf��C�I��
4��G���?����0va<�p�p����O�њi���4z|G������I�r3��B�'�<�/����'_e�{̌O��׎~�藞F�o^v�3�s�q1X¦�ET\gء�_Y��0?w�>T燪̈B^7n�t/)?fVa� ���<@�<�	|I O�xA	y�(B(�e�K���|"]
Y�5�aCS�B�a�+��}�#�(K�H�+� ��\i����p�ī�����|�	œ��PՓ�4v*�r�N���}:9b��0$i�O�8AE�f���B��a��A�ˇ4�&�rL*G���# 	�0�#" �f&�~���Z�^�-Z���NJƔ����8a2�N�j=���m�a�|�a�<9��Թ}z~���R�k�ʣ2�'\9���	��ff�:�3�a���&�d���ig�uX��WU!Y���F�[��̳�Ȋ2�o�'.�C����'��f�����[���p�,dC��֒�����_�0�]4��v'�s���C�N�G'Vr�b_4���ݾ���0Z�F#4!B���#H!���n�$�idXd6���؂���+����Rf]��c��`��&̇��lA2�i�Ρ�)8�5�0!xI$���^'9H�4KK>�R���>0���?X-�	�,��4��`q�SƜp�b8���|Φ���PQw�HTh�wa����N�0�N��5`u~�4��XQa�|���O.f`Y�l��`��LqAc��OR(r���*z��c�D�,��bg�k!���9@ـ9Ɉ��pb�U��
L�T��1bibLR�!Y82���a�.��M]�e��%�~��`����x�2�84/+��4�l�,����
�g^�,k�#A�fu�G����@xi�%��\�7HR0<�&SC�&�Q	D.Y��L2���2Ȑ�-R�]*,�F�p)j�oTq±��1�Po 1�B�7��-��w�iY*�	HE�
!Ie�LI�Qa��I�&D��8[1��2p�b��-4ؼ|Q�uU�:2b�t���!A-G��A"jAh[��"E�5H��\�\,�C�J>L��	<�D|5Ž����������l9#G҈����1�<@� c�?���Q��>:iR=:Af��4'F�#H#M"�P��(z=�H"���!�<<p� ��<?��H���=G�߇8FE�F��9�S��;8E�����\�}{[�"�r��Ȼ���/{t{��|yv*��y�Ez�]���i���!ٍr�Ղ"�*$t�4�6I4��.��:� ��,��Rt��̮��鎓o�����A?eß/����">���D��2��"Kr�/��ia�+�А$A P �/ (!/!B�!J��Z�-읔�}p�q�M��d?"�..�c��M��j���F���=�v�v��fXD�T���>�|����U�r���oY^qy۽tV�o�qƤ�yQt�Z�E�,x�q�,�D"�J�<Hv�yw�:ݙ9;L���*��uM��ѹT���FW3As͈������Z�YPȋ�klT�+i�ʼ~���KV��&�4�[��"�}"�j�
)@CTIyJ�^=b�׉@q�V��	�+�<�-�g0��W�NXY����ͤ�uB:����A޻D����X�@uub�(�؈.bG2ՆZ�Ͳ��@\(	ū����12�8i&��� ��&�w+0��@Zj	��í-��!�F|�Rh�#":���.ab���՟T78�	dG�MiGI,�೽:7�1+L�+�r' �����"�<�W�_&�_���k�����h��رB�����:��U�G�:�ԭU�K���
�s���EM��v��(�)�;�\1a|"iĢ��%"��ծ�'�x��^\,5yyLB�A$ry0�tP�I�([����F�	�\ѝ�KV/�����$�ޮ ���嶞���,��6>� n�T��SU!��m*�J���Xp��A?,_*	�խcn�>G��Xt^��,c饚Q�/�;�X���,$hi�@���U4�&&�L��?�������.C!���_��yY��4�L%�+"�À�z�v�8���''),ai^0XÅ��[��6.�q���>��\L0T+^!��w� �(�+R�#���Ҏ�B��s_���'*)P	QSQ�(Pu(�0���~>^�5{Խ=V�R1a�PGT	�˲�����&��u���[��pR�����0m�X�<�>��'�Y�I8k��0�������(��G%|H�8���'��)����ux�Y��d� H�f{�,�8i�$DF�!��􁐘����iDx������<���a0i�t�zQ4aK"� ���p=,�d<#����:x��H���ޏ�n��H��8E�G%h�9�K�z���s9�h���L�w�zڪ"�N��Ȉ�6v~��>�eH�[~��B@��Ɛc� �� X�c ,iB�B�*ҵ	yK�}���10�q�P~u��F��Q��+X�g�xa�i�v@"ubD�$-RsKŁc8-(��$��ɻ��0X-]j��,2I���>�i7q�#�v�>^\R+hl";�J��40����5�|I���O�bo�I�P���X�z�%�׭ם�{wm�+b�`�(m��Kvr��M˓�|*P�9�s�U��AÁ�9)P�u��'D\��_*
:��7p���&�!��c�%68��ˊJZ3�I��쉒�wX@E�O�p�ލ6O�{��~���D���\ߵqo-*��3�&��v�MIO�O��m�z�m*z�Pt��A�c����2;�؏Kc�'8�tV�V#�z�=i�e��
��������a�4Ho�p�z�_9P��R@b������|Q��p��JgXq�*D#�A޶�C\(%R��H�I��UѨ$��*DMJ�]�G�B� $���+�:p�g� ���M�d!���Ȱ���y���-��&��R�^aN7,�U���r�D;	Nu%���.�u�(�3�ZrZ�W�Y�NP~Z�
�Q~P�~ ����x9g(�C0,����p�Ko��VwyC]$�"���'x��:�IP2~��C�E٪�PJdb���J��67+`���P���1K�{����QQ(] >h8�Sܑg,ms�w�*���x�2#C�	�������<k�n1qyy45(ŋ#���J�CE�Q���ŔP��ߍ�62�fx#�|���Rqg�B����T,�I��1X���R�NL"��4��W��d�Vs����$H�l�i�>�!��oM'G�N�M:N��Q�6i4�:L?�4Yó�Y�<:�$�2����y�$��><O�h�?O���o�p~,�t�nG���k�̪��>ͫ����|�)S]�/��M�e��t*�Jʋ��v�UL=���r]���Z�V��٥t[��'6y��zw�6QT�(�2kkutX�Wj����U�Ki��*�CqF�
�R�M��:�t���(��U�� ,~       X�5j�U!ZV�!{<�"dQ�5Ma�q�T3 m��A3�Td��u�*@��eE2y�L�ܱu�(s���D������ļ̳s|���*� �[l�Ո�v�Sd@�n�W���5$8u��a���\�!��Nc�I3-�&��^�/�B��iCʧݥuM�d\(x�"�ɕM��4i�d2կJ����%/���>1W�P|�/��#�|����b���.%É��M��q<��W�,��8��:3g���߬�H�#V�,�rqQܙ�Å�{�;F���j>XsfD ��� n�L
��Ih����U��I�`Y^A��F{ziUT�j������*0���Z����,�I��m�5Ht�IY�ҍ�ZS]8a���8��S8���]ԭ8I�N���F}���f� ���[q�sZ���~Y�Rb���_8��p��c�d*�5�+�|��Ezt�Ĝ6�aO���Ln!�":"j�޻�����Up_�;;]�I�#�J�yG_9ً�c���x�\R��>�;V5f���)|{�U��(X�>MK����(|�8��L�iP�I�I00,�P��8�x"��}�~ep����R��E�� �hƍT��{�Iҙ�qXN�t�e.�pkzJ�����㦒|(��L7.b!�����Ap�$�ޢ�+�'��1}fth|�+:��С����7�t��"W:ZXyd����P�A�$�p-M���*RR����s؁�DG�2֣�ՠ���>��V+ ��a��YQ)���	L���#,�h��20��/�?��DϾ���ȫ���q���YL�fT���Bܳ����	D�>R�Ƶm��(�{$�b�!v��2j�l�Z��ɻ�����fB0���:I����ZɢTMق1J;�>Va�������)|qM3��A��e����x:=IAꮫ]��#qr�V�rl7#�$@�6?��G�z3�N�M#N��'M#F�h٤3H4z|Q�2ʖ�tii:�i$xxr���8G���O�4����zx�'���D��Di3�n���t]�[}�n��a3�b�Һ�R�uZdE�^�*��g˛�]��f:�&/�~�  /��  )      	�Z�%io�Q�ͧ�B����VQ�
~~3�W_�G�2Y)T�Q�Q���
����E�Ō��7���p�K�U�(oc���Ǒު(.��7u���qP��p�;�Ѣ�X��(�&b6����s�J8p�ԋ>Ä����T��S�J��#�g����#����Bb�[N��$���[��5��~�Pq}�v�ܵ���J�O5����	$�����YK���/a����!H�D7�ِ�3��8qB���c��:	�؇h�[+�*F��+�����q��qAߚ0���{��yB���>Zx�L�g�t�#�L��#;�`�(����LdLE���'g,�m�j���J�����Ln	���Ȋ3������"��A�U���3�IQ���:I���![<{�uBX�p�ll:�L�̵s�ժL��uYҕT�P���4�ˈ�Yj�$���(遈��\�D�n�꺪�����ƺ���YK5�X3*�U�Wd2��L���c����UHݬE�^�Y�s�yZ��u�V�."���jzX՝X����I]���."l���W�3�Ҹ�"�ig���<��0`g������ţD|�NM�����㖚��cܲ)`������*�_?T�Ig��b�J��X�3y�2�X"�gT�#����h���P�-P ���3��W�g�/q>4��>T�|p�F�:�������3������Br����yqXw���c���F��='�8��^�p����#�z=P��4�gQ�SkQ߅j���"G�H z6>4~���&�h��4�i|i894#F�!�F�[�I��H���Q�h�z5��c��|#�Äx��$��=����?O�����Gx�EGD�E�]�*�琢?��xˬNłeqԜːe���b�}�/��¹�����O� +&l�Ȁ��[޽B���1S�������f;�����gݼ����ޕm�0y{������办x�eQ�h��AE��|��iO�4�{M�  ,    % H  	�Jҫ���x�'LN|�lRW/��n��JT�8J���#r���Aw�αo�[C�Px���D����"�B}ʫo�X\�e�R<���-Ve����o�L���;T�'�B|�\�s5�n��=@LY��]�����l���e�76�f<��U�=�w,�6��EUZ��w䐡��;��P�CN���U��"| �&�])A�ɯ�/��x�kE���������h���q�}L��.z�3�K3����i3�da`}"WQ�B��m���Q��MO����C�(�����ߔ���Ƶ`�m:\����i�g�6)�1å*Ƥ�E#�<"̟C:�g��1*��D8����q	�!��J�ͅƸ���1�3N�dH�$V�2a�L��M�6���s
���'���X�R|lq�qc��F{DGt��˓��@�<`Y>�����nɅxE���s�H�K�*�a[��V���G!�H���,]X�3��c�SP��|Ǆ
G�RnQT\F)��uBxTL8�:�:�|`�0���CC��p��{�Q)!c7�"���J<�R_	p�͆l�%S����܎�Έ�3�>�h��[g���;᷻3E�����1�850�d�L�����&ӏ|A3<6�>TR'5k���>�����M��es)�4����q����*:�ז�����)`o�Zx�=�:��r(X���/C�ɍ0��+W�ߟ:p���=�2���6!��HgR]팷�����n\�p��帲�0U����\�����)�cL�Eb>D�F.����ALf{��E�}��<�Q�M��g��⣱�ז5K]��J��j�j��yp��+b��i����G�W���u}�V+����Ȳ��?�����gHc��I�H������|i894#F�!�F�D�AF�N�F������ѭ(���<>�y��'��G��ў<G����4}8G����� ��CS���k�LdXݪ������	��2�qq6��GZ��:��1����ǻ�s�+t�^L���}��%�   `      �B!ZV�Ju��!�ӧc���_�:4T�Y��h���㖛GS5a9�e�il���"%�D�d����uJӽM��g����*9D�������v����JGqvxa'
(�N��O�2&g��+i���po��+F<��<}��^��c�q8���G����Gt�46�*��9�ϱ��o����;F+E*D'���e���^;h�h��a�XY��t�˷��ȃ���V/-��yq3�Q"�,�Ӓb>V���Y��Q�����8V�Rx4�g�A�ʧV�����U�pA�^'8��D+Fj���lˁ�T�wT.�#�Z%�-PZ(�84�:�,�dp�8Li�8�����������
$�,mv!�#��H���CGӃ[���lD/���X���������`��᫨�K;�qG�8��R�/O��^��O�``�)��}�a��߫���S;�n�#ݭ��J�)��n�Mj*M<՞>��Gz�[6�"O���]<����:T�lM�d��&�r���`�qW�(���~m�� n)>'v" �,��
�FY��*<p��	h��j�)Q�0�8Rg˜Y��Z���V~L|��o�4��{��k↵�OV��g�ys��m���n;*R�7���J'��CVv�!�����G �е7�
ɲ��G8b����.�A�m�68r�|e��~_%U�S��OMyf��P^-�5^�(����O��òNK���ل@�f��g�1�~4�t�xi:t�M���f��#M"M ��$�4�(�F�J����0g�<O�������4�����4}:G�<��D�����ɞ��l���O�/?Zo�K��\+;.�Uڍ?I���ec��[�uN}����Sۤ�Z�e��w�7\�'Զײ�c��g�������Y�{w߮�)2��S��맾ͮ��Z�����i��6�(�r)'"q)����51sY/���=��          4!B�k�^�y��Ma� U�5�M#�b�	�rff+�i��q53,���Խyp^�TS�<U�k:J�rSuwu�{A�u��n_M��;.,]����j��o�/�T�ߪ�0�V\Pv��=��y�u�E)����c�E�۝�޼�YU$rFڅv@��/�^����� x�cR�H2���ȹ��#-w�5� חCx������Wb��|��gŪ]G5|�x(աѴ�I'��Z\(�}F9�̅��#��Qэ4J���y��!gy�����.9�����׃T/�P�Ĺ��A����i�h�������uZm?����|Z�y=G[r|q|��(�mp��"�/
4�0,����p��H�|dx��q�i�ֶ�|=q��|�Z�"��F4ы�"�8�E." �M �g�'��r�wR9D��2G�&����lW�3�"��cu�&�Yc�FU�o�*T7*	]Myb��ں��^�ghX�ᯧ��t��,�|t,��g��P�GW�X�+'�<qQ�^3�R��m���q�ը��Ē>�4b5p�h��j��Ĝ ��ϑ$TÁ�r���R1��,#�L�q(B�֯iF����ȍ�ǥ˗,���3����G��Q��y�yY���Z�Dז�i�}���'���B�Ө�cM��tD�X���=�F�O��U����S��AO�9�.�QZT�~I�\��8&��hO��IS��Qx����pC^����x��k��{;.�=�G$9��^��Ȥb_((6�Ũ�cOs�Է��y��~�~̑��y��B8���5}�b�Y��
>���u5!m:觪F��es�:6�9����Dl6��1���(�3��
><@Ϗ��:>�%���C�p�"AblK6P�BlNp�Âp���4��O�>>>4�O�0�� �Jw�n�#g'�ְ��V�$���}�q'�N���Wg,�9M\��E<ʢ�����B}Y��F�V5��5XTd��®t�d P          �R�*U�A3*[���mR<�%_��:�\S���R��T�m��NR)VyQj�/���.�0o�J���$�(�1��'̦�m]\)z
�����>R�k��l�hJ��J�8�����yR�(���'&x��ӊ(�J��~��i��nIV��Ce'��7+<����(,�F�8�"g�Dn�ϸ�#Uj�Iզ5㒺���W.o�߈��yus�ի��i'B�>G^����8�N����,��p����=&�8eK�5�b!���4[�:t�N������?���H�ˈg�	NHm���>X�E����-\[lm��妘t����ճ��.��cWT��!���������cy�-WV#�R�B��E��
<��L�Ox(�G�g��#�w�n�e[rnk̙v�1�Vڴlj]R�.�L��q	�nʣ�u�Mj��J���F����ˁ<��?-���m�t�^\<�p�L
STAs�Y�.dgU�]է�}?�Ua�TL�Gի��Qn��p�K
9����j�/�\X��̱���0�/����3*���l��,GW���YD���%M"�l&B�?��,��_r2��L65J��/Ķ�R�s�A�O��.��1p)�(��u`�j��ې�)���� ���CI]�QUS  ����O�|���'�9��ɦ�8������F�hM�DM� ు�����D�k��Π8��h
��
V�`ԁHo	 `��F	! ���6�FB	$ ��B��X! ��B$ �	!`�� `��	$`��B	$ H�@�P��@�D�D�V	B	 � � � ���	X%%`���P��T��P��P�P�3�r$�H�@0H�JH�	I�\,�JA(A)���0`���BA	��HA�4��i1PАi���$�C�JA!�L#B� ������03!�\PD�f,A0��p��� �@@A�����" �& & � ��H"ds8h)������$��("H�("�H����`X��	�f`"	� � �&`��X�8	 ���$��&�"a	!���$�a�$��"�@�����&��Hb%��&�f�$��"a	H	�`I�a�Ba��"	!���Hb& ��d�"`�� �!�0B��0$�L	0�P��P L4$��0$0D3
L$�@�P��2022�8R ��R
JVHB	B	BR		B	RYJI%`� � ��B	%�LBJRR`�	`��$ ��B�*r���`�<u�K.�'
`M�	�o\�0� Ĉ�*�5T���	�������N;����>����.�����o3��ۗq���yy���^��zy{Q�x�i�z�o��ǯ�5��0{z4΁ty��ä����ܟ��~��:'�����gO�"�(��}n01���?b�Q�9������&(����?�N��m{�����⑰=�&t:4_���/0�8~��a���G�@���O�|�?��*S!�����e��=@2�!d�H=����Ra0�M�� \8�mÃ���x'a��g�Cӕ�4�c$H��o\�S^AL��dA�-  &(@5�@�,��0 rQ0�L*1()@H+�揵Br�m��&3�>����8���q�t�y�"4	A �D4  Pm��g���~'�����{	���~snI���O��p<�b9t�`���y���A�~�a��g��!�@P�y8lW�ǹn߱w~�5��OC�|�&���7婎>3�w>f�y{����Q�	'�t�s�|��:���o?M��}H�(tv'��r��~kG��c��='.F��n��=P�����(
�+?���o�0{,�Z�s>cc�nj�N��HS�|�u`QE��pv�\�$X{y	����a���aA!���*B1 �0��BO������쉍��j�C9'0je~��T�'	x	�0��=��*�z�~�j7�z�"���{�D�D�;^�Oo^���>g�Ϡ|G��?�)޹�����bz'p������ ��)�0G��������'$��A҃��I_��C�*
� RR�J��`�8�?��N'}=i�|��u�H�#��y��BF���_ɡ�Uhh`ȸ�������C����1} �<tC���d����.�vA3����"���G�c��:�4L&0�:R9=@�a�2�1z�=��Oo3w�sSt�o��ꩀu�#��ӈ�W���!Q�ɟp;Ws�;���~��;N"�/Xv&��9h�}X]�=��0�狿�?i�2>4�2�0�.������.�p� ���