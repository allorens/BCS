BZh91AY&SY���֜߀`qg���c� ����bA��  |>
�P�(UR�֤��QQJD�-eITց4�-�l������m�PT�T�R���5��bKl[�R}�v�mIV�Q%��ihm���5��J�F�ZͲ�CTԢ��Y5��"-m�`Ԅm�ja�SfD#b��m�H��m�d�d��ϻ׵����m�Q�b�i�&�6RY�(R�[j��(�[f�M-�����R���M#V�Dm[d�����0�֪X�U�����մ�X����k,�le!�   |7Z��� 8m��9-��$�qU�;�h����k�(.��:�m�4dmUU��j�uk�T]���EHմe�-�%�A#�  ;u��4nS��m��  1�t-�s�@)��K v�wcM�PuL�6�� @v�uA��7]� %S[lB�k��  �= �G4�@�p�u@ 9�۠��t� �]�GT��� 1��@�.�\ �[���N��)��c*m�-�
�S'�  {  ��z�@����hc������t4���҆�:;�� � ݓ� ��X� �w;]�U t��)h5Z�iU��P�[U  7o  Юݧt� qc��t���(Z�SJ�75������j��uܻ84 �Z���:�B��+��A��V�֣6��Ykf�Z���   n��R�u.��:�g�$n. @�����:9f�Ҋ��ۥq@�۪pA�sv\�P)�r� n]��L)�)��i[m���R�   r� Pi��M:P7����Vt 4iwS��:��h�r��� ��뺠f�An� ���:��@�f;�@�Y�liBѶaO   ��  3@ w\ w[9�@ݳ��0�w*`� ��+@h7v\ w�U �ٖkh�U�Cj2���'�   �� ��-� ��
P��  c wa�
wv]@ ;I� X�4Pe�p�A�j�Jj�j�,ՙ�ѣ�  ǀ =��  ]I� �� 4�W  m�p 
��� h���A1@ wt���     ��M��)B0� �ѐ0�a�{A�RT�0     ��BR�        j��	J�h 2h     *��&� ѵ      �JP�T1&e&�14ѡ�FG��� � �|������2!#�k���E� >>=�o���|?g�y�����6�?�6�lm����m����m��6ߑ���#�?��~��������!����lm����U__��m��6��!����m�N�1�������?o�b���8�� �����;|c�`�8�?�<`@���z �0�p� z  ��M�z6@��� z �6��;=l�v0z op�=�@��=����	��@����o�6N�{l7�8�`��pd�=`1�@�`��ǠM���Ǡ@�lz60o@��6�0�z��4	���@�= ��q��m��� ��o�8ǠL�	���O��i�_/��#�^O���g����Cz�	R-�-�t����QLT�,V��S���O��nb�-�UWiЪ5C�A�hX�9��n��Af��s��c��l9���QULh��rV�kV&]2۳MM��Uz�Q��\�t#��2��Ӑ����TV���m��x���Y�0��a�S�KK�6ޙug�A37Y*A6յn�ZU��܆KgU�M�HdV�U��$Vѽ')��aa51��Ǣ�[�r���7CH�-�L �\�D��>�:��iAN��]���{F�r��X>KA*U��)����=���n����gu}�J�V�M`w��%[�_Ⱥ�'�圵dL��Ikb���������J{L��i2��wM��K�2���Juu��!1��,ܺ���h�p���0�ӆ��P��(1�ʂ���p�0JJ�a�Wy���8C�Q"ƭp<�(��b��3zjjU��h�K]]���rY���st�{5Ayz���v�U⚢�P�s&���ldLw����z�8���6rn�4)l���Y�c���ع{f�I�_e����۲ƛ��P�
#�*%�b��T�۷d��1p��C6+hf�H�69��*�7Xc�^ N��T�n�2tXU��`ZP�S�+�eޚ�0��s�q�"��e}����YMT��c�(4;En��q�I��v5��@!;��
��ܨ���7�U��<�nЖ�ϋx� ��#�!���)��ja�Eѵ�,�7�!�Mh�YuP�a�a��
�B���!8�\P�d�Cs^V3��)(S7�]��q]�J!����oqW��F�����2ȶmKN�K�	��L�-^�d��Vq86lB��(���6Y�!���\ܧd��{.�d�X]�A���$�@7�&�z�¡K˃0)n�ic�Mf�Ì��̘\ә�)A��a%1��5w���Ek:��t�дA�+v2��g	�z1e�&8�)�4KJ�ى��Œ�&����XӚ����<������	�)����C{zp�y�{�ؖMs7� ��,��[nT:��/��FV�O5��X҈��I��zN�x�Mm`�nXѫ-�i¥�WY��H�d���0��lf]QŇJ�%PT�~:E��+��t pPz��Ցx�4���j�P��,n�U#VY�*Lst�����'fP���[cjh�(�5Ȉ�mqG��9�APlv�%T,V��5�c�.�-�o(]l'*�5�� ����p�Wh��?N�M
�s �6�Z!��d4we-����͛OB(�����̤�E5E��#"=r�I�85֙+"�Y�Q����,�̓HԢ��hDʔ�ژ�0.�����kN�ޚ�cf���m3t�
����3�u�9څy0I�K���44V�j�U��6�����R�K*	�hH%�d�x�L�),�������A��V�jGGʵ�I�ń]�9�'WC^���)#*�M�ٽ1܈�c(�[�˲V�h���&��b��� ��j]m���,�c�L�t!!���74�^;[ �⸌`����^��u.��X-�n��')�K�x�- a{��z�R�J�6�Y{����,ʫ���WY�R�wRk�Z�vF�T�J�^
9
F��5ktʵnZ�enHrM lGv�:�M�{�޲3X�.[���(�5c�/rV�5�x���$�c'�aC���w-������*F1 r�5y�'c8��*�L��d���{F\��mn�R���ZqȂǐ⼏+i).\˙���Ә�|�y�F����aG-wd1�D�����	��ݱD�aV�(�����ޡ��;�T)o�TA�Q�P�%K��f�s3U���֨+eP��53I�"���7@�Фߦ�nK�(�%�
�j8�#]n 974e�P��a��:���g.XT�
�m�K�[�pj�6�H������kk{w�k��a�X�;Y&#4fح�[E�q=�W�C桎/��"��o/sm%6���T�GV]�vlٰ/�z��T)�+�p�.�R�(?�bp�آuk�m^�֊[�[�6Ί��l�ZC���;ldb��Y�C\ I���Ӗ4�KU�ݳ��H��Q#x�RaP��v�䱻$PQ��p��WO旉�ڷ4��(����%Ce��Z�U�7;U�.�30���WBӬ��2�KY�a��5[�8����˴Ci�yV�(��b�L�m�F���	�7UԚ�F�Yd���=�![JȖF^���=�ݜK.���������̺�DX.�h,�%:�7[���:5�U�(o�areCw&�H&P9�*���W
d,�q�Gl����]��FQ!�,Nꎝտfna�`TΫuP,�:�zq�Z���0ȱ�ChA�9�s*�ۘ�Mʓh�F�7���6�z+Xm1����tՙ`�X��[�n�ʹ�e�6R�^�T��3���0-궆�D�]��.�*Z��,^
�kX�Ǘ4@n2��)�Pa�CF+?�Y�(驭�#�X��&�Kh��-��r��f&�I���둒�-�V��:eE��A"\�U��cT�ln��y����fv "mkݘ�c�h*,ͽ��7;��G��t�7PÄSI���g\�����I�WWX&,F^�+s2�[��h�L��ֶ��He
A�(6�欨^��P8�m�!�?��hZwm���[�J蚔��V�$Ks0mH�Aw��x���L�`[4��U�e9V��l	6��r�&ڙ(��Ӡ+�v�gk-n={3t7�2�sF��732�Ұ��o1u��WY����Xn��顬U0n��##���ǒe;�ӯt㩻R;�`l�ˢ
,��[˵����L(w��:*�Û��=u�БS3u��Ӳ�5��۫�Kgl��{��P�W�M�X��'2傑�l�DR3��[ɤ^�cY�V�6ti�fۃ-� �6���cJ�3�;h/뉭�ҳab�ލN����Q���L�B�ܙ��b�^����4̂�M ��^mՔ!�ieRY����Kv�-�x����Kz�+�9���đO��l�[w���n� +;x`�͹,����^"˖7^���'&e�ڃ�dS���LZA�jUq��P$��x]�W��T7`�:�b�|�fz�a9f��nh?Y3Ls/���d�Z��(X:��$ĳ1�$+	\���q����9O%X6Ô�̩D�7���X���m�_K�N�n�ǋo5cå+�"�]fQu�b	��TS7�mX�R[	�A�I��)�ř5�m�t��B�B��ΒΜ9�2�AL��0ֿ�ܲ��j�t��A`#+C��[�@V���v�*-�t�D8�L8(���hn�)��h��!+>f�12��d�Z�J�j�@����QŠ:gJ�-xٹr�Ѧ��k�M��Y�m%�7O���.�:jӺEc��S,�.�L��Y���-^�a��,�D6���8m�b$��x�S �w[
KVY"���e1�P�θ�
��y+�m��Z��|n=�7)�a���Ҷ�V��5y#%��Y.a��t��6�*�5��57$h��z��Zf�Kw�cHݧy-ksH�˔��XE��7h�PI�+35{���a
X�0�W������e	V�*�ǓE�����~�� �,��Rh�ڗ1i��KZ��u"e�i�'� %�7p�!�Gr̺�m�u�LS��r���t��*f�Jڗ*ن��NJב�A��
��=,����r�phӟ\cb�T/k2�қ�J`%�;�����5�Ԛܐm�X�pY5�|&#�I����3Cl�5f���z��{�ɩs2=^��B|(��u0,7)�v�:r�3���I1^���U�%'Be�0��oXŠeJ���"̫�w[z��'��e��+]�L�n����,@�V]t�Z�0�nf�~��H�V�/�E�́�{o0��]��h�0v]	��sI�cٶ�X��jU73�.dV0��Yl�ՠVX�w*��t��t2��T�����4�4n�ʗ �,��2�6q	]�YY���F�P�vLn�L�&,�����$� :dw)ɷ��{Q�_%Y����٬w�"���H�w�(�@6R�f���k[-^�K�46t,��Ř���^�7�&F�,E���ǎ]�[�*�&�QAe��9�ī$z/N���F����WW���cdi`("��e�?���Z��]�;l$v����ܔ�N�sJr�jx3r�j��N��9{@�C��A���+eV1��-
����CГ}����٘A�٫* 0J�9aZ1�Ʊ�\�Cq9)-�ZbN�Ӽ�&��{5K/.;QM�K���Y/C6����yy�����az4�ᗕ��1c44�W��GwUi
`.�A�b�^D�6�r�ٯl��Rd�����ǒ���sHl��^ ��bj����O^X�1��=Ź�]J)�ik6����˨KXEf��� ���z54�/�1b�i�s�$mE��Up++\�p��qE/��큶�
�NVn0A,b����u���n�kl��-�V콟TUX�$��a���V��mXn�����f�m\���$*�g6f�2Re��ҏG��S�$����x_����(��M��Y�΀JxF&�)i�-Vl(�P���WZ��.�n�nd��W4�,Q��4��� �ԥৗ��e�u�r�w)��11jS���"*��3o��U���ٰ���e�`���U�F�|5�T劊��G���梪7����ՉqPt�M��t�6V^�Y��е/0j�Kp�c&�)P:`�
!�QL(���ȷ�h���/$�4u�bn܄�[��L��a�Nύ����
��ˢF%A�q�ʭ;E�M�N8i���8h��mӭZ��V�hkt6���MN�����{��Q�n�w�]C,Z�(7{z�F���=�Q��)���������w����PA)����:
΋��S#;l��`1�MJ��n�$�聛W�E��Uk���]���ïJ��n�cʇ_��g0h�"e;����	%�޷2���IVF��u����t����c�����vY���g)�r�B7����=�v��kU:��0�d,E�8������{��]'V[9��I����̃Xp�H���L�Z�x��υO��ͥ�T�v�J�t����X�t��{��	ԭ�WX��)��r+2#w��fd�f7E�c�u��7H=�gX���B
e7$;�]Qe,0���fU�X%��ٍ�f����0�i��ؔ5���_�����֝sE�є��d�.iE��6i�5�q� V�
2�f��>M��Z����p6aR	PP*� 0:j�v״0�JD�j�ʆ�%� �MЧ�k����b֕%�%n�k��u�,Rb��ڙq�.d�I����EoН�m�1�]��qP��u���uL�T&��f^懢QG.Qe'��fcs3��n���-Ab-��w�N�e�����5E�,�*��Ť6ȳ#�.�C��^ڴdʽ�6F4����(A��ZAͼX6�n�H�%��VI�^M��8�Տ+//]�qém�u6���/���rXYK1��Qʿ��3�r���"��fH����il���J���-�5����l�A��7X�ij�X��;P�B��ʨ�L��.]��sRz��F]�y@*׎,6�B�\�/�9�ͧ�L^Q֬�*�1{�h��;�:��ۛg,^jc�X����&]�J�yS���/S�)�fn�؅څ�,_��߭��ýKQLV�A1��:��6�R{�|,1�
����>@�L7J��+J�V2����Z:�.���y��8;�m��������}O��ܷ3lQo����ԛ��,��72�3W��Z	�QZ��z�M��l�.�D�kye�Ƕ��c��J��s�Pźt�K�Xa�Y��E���e�(�ܙM�ʏrJ٨�Z�y���t��f��GcD�������h�m�z�9�h���,ɹ����&PՒU��92#�'�%6�Ŏ���X�MB+v�����+1=�Ln"kO*1�6�m=�Aya��L��m3r�c���L��f^�N�մ�L"��E]�6M�+/&|[̵K�=X�_;�����UH�Y�Ý4f���45�o�ᯩ�5�Ƴ���K%�A�q틲�45Cj�]ͧ�e����܄��@p��ao [�j�Z���� �,��eb��d��r�O^˄���Y)<{��5�GXX����6�b�wf��N�Y[Ytw4��rm�æ;�N�wsJ왲�`�5X�BMM.�k����\^m�v���.��WC���I�KUy�
Lj4uXTʲp�#z�V=�ս�*��a��&���S�k0�!�PGSYEK�Ӧ��[0��w�^ �ж!xe���kLyL��J���wf�`쁗7��q�B���߶�fi�yi�2M�X�m����ݽ)�v)J�kF���L	����]�"��ܻX��-��rb5 v��q��(��&av��T0,H�ُeeVVl���9��֖�ta�h;�#][���
ýM�Ot*N<S�/lT0�x�
1U����z�A#5��cB�3v��r�E��2oKD
��z�ce$��8sb©466p�*�	��V�փ�mMq�1�R�����z�,Ǳ�. ��V�Zե���ܳ/b�M�U�,J
�Q� ��Ӊc������ߋ:[�o2�}(�hǡ6�Z`��V��l��'v �Yॗ{EU��.o0�)Q<��j�+�	Wa�σ��w����{�$(�1a�*ʒ�t�ud8���!��)F!������T��*�������1�v< ֽ.,6a�LhP�Bq���J�8NO�{~�5W������>�`S���#��ѵ���Owq>ž��K0-m
���gHm
=��v3�n{̷d��\�j��swvC��8�"�p�JR72�6 ����W���B�q����Z�c�v�{ވ��~�RB��T��^G�9۬S]��AV.�{L;I\�y(j�W�:�q3n<��gwR�jÑNm@�;q�ֱ뤫Gnj��5w���0o�ؗewd�����)Ψ��a��G X��ͰwzoHJs7����삢���r�:�oN�v/��W6�'�l9�	���#�Î�! �p��c��^,�ޕ�N�o.�[#]^wv���k��*�עX{3��A�mՆt��Km�f�PI�F�S;h�t��å�h��huEyd<��݄Թ�bAα�l}{�l����<N��Q�V[&7a�M���z����n�J(��.x��D�)j�;2"�8V�e��6�Un�ۂޭ�$]qڣ �qx!��+������uэt ʴ�v�%�O�2Lcv����à��]C�ai\b�����e6*�V
9 lI[*ru[�ܙ°�a6P��e-�ö�ͫ�*Xa�v%cB���of^d�\se�Gm��E�j���$�n6��q�f�4q��M���i:����yv�2�U��]@3G�N(����� ٣Ñ�ԗW�]NӱP Rwi�Weݸ:iżIqq�!���}�0&�re1X�K���\��^�<7\v�`�ѧ���\6���[����������u�t��s���Ua*��X�F��J�C+2�Ð-B����	6���������}}*�˪f�:h�]`x�,G�!%L�s��M�5E���V#F�d�2o"�˺����ur��%c�nT۠�B��js��)��u��j률X^PVˏ��bt�������[ɺC�^�f�F�ee}�N}P������Rjt��n��m�Nsj�Y���j���m���[���f9[8�LA�1��Uǽ��I3Xȱ�u��\��T�j��&u�3k(�?l$R:.ͩ
��҂a�q2����ۮ39d6�C%�w��%�okmpn�]|�ޥr�̛H-zwՖt2�d�_9��p�x�#w�m�1HD��E[�I�V�p��U�޷B��\�k���0��^��9�`q��דf2fN���ǋ7gnfM�5��c��WKR�5�j�����ydpʠf�ͧT��Voss��\Fʘ���6m�{�F$��^��S��)�˹\E��62�7�Y�a��p{xRN XE��r];���k�|:9��"v��loBi��3u��*Z˰kdl<�Le�}-��\l'ۨ��g�eGE��i�y�lE/����&�����5�"ͳziV�zp���k\��S뮩غZ=�ls��e�l����t���YfK�|2{۠�o�LP^�tq�~V3�.$��gN�|�=�������0+�}��G�Fݲ!�t{ghl�����j�(]�(���p:}��,��dtٔ+^��k}�nB�c���`h;��]�����w8�:��"����wDR}� o���Y��ȕ�[L�5���չ�e�$�E���\I6g^�4z��}�)�\���a��_f��X��5�E59B>��N;o����ΧM�5մ-T�o)���`��w�����GvI���:���;Rb�uJ�}�G3�(X�ڧ+�1+L��P١�ꅋ�w,�aw�ϜL޲௷��S�6�E�Z;!��Kh�!|���-�J10�	e��`%4���k%ի77p�m.��W7M�z�Mj�I3\)q�6ʕ���,S|�e���N�n�H�f��f�vF�B��=7dQF5����T�wA�RR��j���ˮ��r�T�bl�d�ޣ��	*�t'���)t���Z�%꾈�V�A�qcg�d�8��F��K�B���_r�uZ��P:z�N	q<���rZ�GSVP�u$�� R��뵕�Kد�s��q=�!�k����I��nV����2��x�j�����*du��J��{�1᯦������Ti7�F������c�L�4!�₻Q���C-�Y
j�[<��H*ذԂn;(b�����;2ًk3AM�ې��`j��v���%��@UŠ�p�E�2�ƕ���T9��㮒��2�=<�D�����WFd�\�ێK��!�3-hbS��H��u�:>Q��{�F4�ޥ�QP:K�P���nh�qR�٭!��^��H~�7ܥ��S}��:k��T��*�.
� W�;oS5�g1t4��l�MCH%A�K ��0#���G�Vh��l��͒�Q�	u\7meT���v��:���6XZ���V3A��u^C��{e��!�q���}Ղv�u��^=�H�O)a�zꟜ,�9�M��9�h�1������ѬP7��J�C5m�&T�ХNc9�7VnU�T1�b	��
�}�h��c��뙫_e�4S��3�7�;�aBt�ʲ��Ӥ'+��R-JlfM�����������S��#W�fʐD��iv�E�Ov�q%�T���v�ިouW��~�"�Ȇy�ǉ�u�-���wvfO���Cu���5m[�5�>ԃ���#�b��j�+\u@�+��[]�s;p�f9,�Y������8T��'A/[�p�wm�;�W%��O������`�n��ש2��mn%h4�-�V��'�+'>dڙ1���󧣟���5�Cz���\x�,��q�'6�>�)��鹘���I���sUZTM��P�ܪ�w�#򕎖�՚�"=@���ؤ{e�j���=�G�X���s���s��
CzٰA�[��G213S��r��aY͕��N��&�y�r��v'�ˣ��Lu�KF;�k����촭���!�(tKlU�5�S��-�"��-S7}����8�������A4��2Yl��8Y=�p�Sp��&� ��8�+�i��d�+��}���7��|2�"���ne]�M�v�#@����wn�ӵ���r�u�qP��"@բnu�'�Z��v�5�����ݼRC��R�;��t[c2h٣A�u��ȋ������vy��Y�j�c/�<�e����;$<4�5�Y����fh�iw���CWd���vd�����ǍU-t����	}f�J�;�6�Cs%[���'�S�bg5wY�^�kx���S��'*�쨪WT�!�����ʤfv���C��P��)&L��AD�t,�]�g&��S�s#�u}��U��o�V1˵��7�lt�t�M3&-�]J�i�»�v�
��Κ�]��I�ԋeC�B\-��n:�m2"��t�v��r-ɷ'P�t��P����8�:mW\��u�x��zN�X�j��o.�E-��W'e�O�Φ�,��f����PR���ɲz�i��)Z/��N-)$�)m��2�Y�YC�0J<��Jq8X4i���ǖ^-٭�7�pX.|y`�4=�F�u��o<�`3��ΤPX������;�y�R�R��������v6�C��/��.�0֩�m5Ճ��!EY+�ʱ7����.�5s�98�;�U�	z�ו0�̕\6���̐�'`EUǯZ��(E�WE�5�^B$�ip�x�w����$Ư:)j���k(L�%�Ѣ�ok�3�B��Ŗ����V��>��c��F�כ��r]��d��rYv8:u�bAOW��ִ��f���ԏ|d[��B�a8���Y��ݳ�^��y�Z��{�11���QC����)�%�k�ճ;���6-�3Vt�����&
3���Xk+pm;��_Aۓ��h�eg0�6�̋x�Dp,T�Ч�hq��h��@z�tf���;Q��N�Sˬf5R�)�ֶ�4D�c��,��[ƍe��d��W�C^�I���s���4��޵�ڃ��*b?j�gZ@��;��Z�(oj��4�qy�B�uθ�s7��F��ht�d%����n#TT�nL�W�.�Z����4^=�-��s"@�,���q�z=���������w����ı��	n�3�ˡ�֙�gy�Vh;�h|�i;�)1�C�E�նz��\L���M�$��.���۲f��y ���s�G����0� jw_)Ij����ދedv+����yaRund�pE:���Z������ej͖b�޼�qnU�W��@CQ��t��n��OT��s��q��[:�o8�#��)�������ْ�]�3h��4Z�F��b�D͜�Ɠ}�&�$�@H�.v��,| ���T
����\�����m�bv�<v\I{��eap۬Y�ce�7����A[���hP���S�[�����̼�*TmPѰٶ�:���]���y�m����wJ��g�Hz�KLULİ��/,:�I^+�ݶ�Y�Z��+�S.��x���:-*��ã�oR��u�Ī�T�Z3�.�`Nn���j�t_@��,�7l7�d���8�e-m��΋�ٱ_m�]I�{�L=X1��Xz����@��R�0��l�W��m�SED`�e�d�,T�%!��7, nd��ʵ��]����;O5�sZ찺K���#�f�A�5l��*V M��ޣv&Gp޾81iN�<� Z��;{)�Rc�w)���&�����\�3z�*�0P{n��_v8����F��e,.������f�-Н�������tr�rbua�YD��C1Y�X�ҋ�u��K�K�.�������j�6JNv;�5R���p���U�PUg�}��-�'Wc�ʝ5$�q�}B����QR۰����Ɠ�����-ԃ��ױ��-��;Ȝ��+m@ ���f[��-�����`2e2H�����
�r�1$

�\���B��;x���9w�<[|���wY�	�(��Y8����<r��Km�6ix��K��5ӢW؆b�ٮGh�I6m:��P���{��R�8��A��y��ݜ{���
�pD�2Q�ޱ.�/T쳥�j�|��p�Q��x�x�mKC;�s��⭟w5��;Q�����P[3Lp�y��4�����Ԕ��-h����]g*r�M�Qmp�uN�<��Y�F	N�L�jj7��a����*%�BT�p����9�{��ٺO����zjudЯ����rH.j�+r�O��"R��֙M�`�����}�e��;7�9�B�D�7M�Tܬw&t�eˣ�s]�9�OKGAҫyp׋Z˖�we�9I�Eo5*hq�K':��^����'4�IWV�3�2��U�%��1UH�TAլj��3�l���,*�w3{A0�k[�E=f��\-��5�
��Ӆێ�gM��gu�\���J��ʒCG���/ywEՉ�˶I]d+�Y�=�2�`Ǩ�V�7շ]F�t7K#�i���[,�K):�	�	��c[ڑ�/`�u�����\]n��Nm�(���Gmr�Z���R�ʷ���>��3�A�b�
k�t�۷7����Ç�˘�|X�r�M]ĵ����,�c�U����@�|jF)8�Z�ң�=�BW�>ۘ�ǋ$�D�+tq�Pu-��Q�V�W[�,�����ܖ�1S�R�xV�G����37�<��ȏT�J����t�:�m��l�<˷2�Z�K�Y$[ó�0
��Dd�� �*��z���7�IR��kx���3qD�\��xL7�&EЄa��ܕ�&�][yi���e+��g1����M�
ɭ�/��q�2;���+CG�;
.�G�J��|%7�H�:i	�H����Pέ��%�IvZ�݂�ͬ����܅)zK=o�9�诉��ENw&�z6�k����Y��}�\-�Q�j�D���hʰ�"�cf݉�]�@弶�8�Z����w�W��ʕ|��N�nZ�TUu�]ݎ��*AŲ'>�wѫt�(_b�]6��S��Jɥ��>.F�c4�*�R�ѡ�{\�B��K����8_�:{
N��qQ��W`��,ݼ����w�w<�&�Ŋ�9���#��Z����!�c��Yƺ�a�an�X�����XZ,˭{pȯ����u��j�t^��w���lY[����V���Fm9�Ƃ�6�(Q:�ھ�ξX�gN]W���.�jCr������o4���70�D�l�w��p�B�M��� WRX1�tX�g g�q��n w0��g��(�FK�CCy]0ix��� �y�v���h�wvN{p�zCA��+6�қ*'g���ѝ�B�>��96�[U���U�0�5����C^���I+9��i��0"���xÂ��l�η�Qf�޼˹kG2���e�lu��v`K�.�u/��di�՗r��;%ܵ"���������;7��=��w?�̊��+9S�VK<*�Z{r�l�IZ�ڨh�ȫs6n��s�˝G��5Ѓ��Ș'����"-���	��2Y����T���hV��b�+fb�'q6u��@�;�Gd�s�>Z*\z�EŎm���n�mTlkɄaڊ+��[eS�BvH�oe2�4d�	���B��-�#��o�|��GT��C��jT8�t5�[�7W}��vV�����ϒ�9�I��ֲT9�Gw��rd�:���xn����@.o6d�gcz����!{��l܋�z%��'��
9JgA��{T�>���l��ή�`xd ]gM;�ʊܫ�7�f�|��y��\��r�]��.0����-�{t}����.kF<Δ�%�O��v�4�n^4c��D��g��g)��Sd��m�.f�;���E\7:�a܃tr���I0�K����Z����\ݸ�s�2k��vp�tF.�����s�A0H�{։�Z`��ۼ[��v>�
��5	7���8P�k�����eH���N-əiД�]6'.��s��5����#�����d A� �HN)>dD<i�/�B����,���Ŋ4�HA��TZTA0�FQBH8�4ajZ������ڻ�ώ���m��6�w������� ��}�~ϯ��� ��������}{ lo�������%�K��L� Y(H�E�&b��XDbh�tjQ:��f����[�o����ٜ1ղ�S��'�	��9[��Bν��;�O^��q�u*�̈́2����ͩݣ�_��q�E�K2�
ʊbE�I�٣���ShRڌA4��]��׼7�}dY"�=I��.��'X'I�dn��J�P2���K��9��	mr�����
�OY"X�=�p����=K5f���:C�����yJ��s���$���3��R�֊�K'��W5)U�+#4sV��wY�02�v톅��^�b�;��CB�|�5���4���G`]l^4����[I�S.q_B�U��/:�`�I�����;8i���[���QܕA�¹���>���[��AF)��;{\F�[[�1�M�}n�|���ۈ����x�F�wWT��������J�7��
�!�>��y�/��V��Y�j�}b��z��в�q��-tQ�rs Ҹ�us�jQ(_��z{ll�]���!2��ݚ&`y6���B��
���5�L�f٠�e�+[�Ċ��N:� ��d��T�۷L��nl#s�Wn��s���HĐT744Px�x����x+�Vw�h+��������m����3����q���YTj�ޓOgo��qchRt���1	�6���9�tf�Ү��\�0�8��*�:v[���j��[6�2(=�,��f�	�R��i-�j��؃%[�Yn�Wc�8�f�S�8�ہ5�2)�^SUr:�>۱���&k��,SD9�E�yA�D����S�x�X�4yY��Żm*�Ʒf�ǩ�I������AX�h�K��FU�ηӂ��|�{%[[�ib<�7��w��6����ghU�De�-z3�1��2C�d��S,�,b��덜��Fd5&ţ����>�w|�ȋ�ꋐ6�C;�-+�kcT0��Xu������.�k�ݜ�N�����O^U�5gbO�li��1�"�	����zb���:����Vi��ػǭ8��L��3a�f�|!Ĩ�a��#���U�E�{&j�Ɔ�A�*�$�Zt'e܇�ݘ��*I�m�uA�6س���4a�J��ޮ{	Z�Spl;{���7-1��,Z �7,эG4�<��8%�c��fs,�6:�s������B�W�O{p��qU�,�������a�D)!=��H�}��z���A(���k�n�a��v�����9��Bk���{ئ�Nu���Fu��[N�e�V�--U�Y�{��o��Tq�\؁;#��)��p��#^�2�kg(��z��hn��J܁�v˃�u��ח�+^9��P���d����[��ɇ�M��N��,0L�,.K��>���XGd�x^�4%R`�c�Ӹ�V0#��[̭设Gn��yn�QaA�٭-iM|�zT�]��CKGT�����R�%��rUGp��p1ED7Fm��m��g9
54��\��]&9�N��ϸ:7mn!(��� Q���O�c]"��:X�öv"���B��+f#�Kb@�0R��|��˳���/�:��4#��x�i\�Z�V�E��a��J�U7me2&ứȎ����\�8����\]Se^�������=`�����_ɳ;�dGj��'6d���6��(���Iuu��t:Wx��(�0J1U9�.p�s�+�"�5��"������t�K�l��W_`�w�U�y�N]Ⱦ{|�t��]�}k#ܕ��jN�k�j�(`Ed��ݐ�ݤGWya��sCO11�q"� �KT�{��2V�sN��(���u�WP�r�-�u�bQ�#�b]���:rS�ѝ��Z��(V�fZ�w����F��.�m]��d"�[U��μ��Xғ��s>��O���9���3J�&nh�7��$�`3/���^�d�onvL����3Y�7��и��TJ�M4��4ט�2Vlwܪ�E��O,�)6"Z�W2��<۽��>R���`�j�{��/^�S7���M�Donu�Z]�	{�rm��˚]U��a�f�΍O����p#7C��J�IZ��]�/-f�m�VM�X����aǲ���8�]��yW�N56��f������Y҅�c`�U�jV̗�9.
巴{oAe�K)�k�y�#�{�}��]��$*�Om�eҷX0�ˮҎ�pJp��&�$ʝ�[F�ԷV����y����$ss%�YnI���j=�S��r��*�J�a(�nE�Czܡ��wrޒ¹��Uќ`�+D���}��"bs�z����;�r�̔/Z��b�15my�a����BԪ��kt�^��:�* n�=(�I.���i�� ��h�b�E�w��1��]U��$#L�*�)�b�O(�v�۰�T�X�!e!� �p���2��DѬηXܜM����*螞��u�Z"����PU����(�*�CG	�	p]��>!��3f������h��V�!�Β*��Y�#��f�z��ab�j�	q�`�>ː8��{α�T8h��1�v���bd1\X+�R��p�s�/�cD'���О���9a�.�C�D��+۽}��kfw(;_T�`\X�G+�ܤh�/궴q�S,gӴ��
I=����qaܒ���eJ7��uH��Y|�x����mؽ�fY{�n��"�2%�/��\�Q`<{�4����z�`�ﷃB�D�c�uѽ�u�ӣ�o
n���/:�B�ų�\D��&�Փ����f�J���=;\<xh9ղ�&m�i+vm��7�)���z7)��Cuw=�i�D��@�!��Y���ܭp�S�f=H���+��o��͝.���8��:�F��D��N��s�pC�h��`��[|��Y;@�:_������dc�I�7K� �[ׯ��c2=�n�EG{��۟!�r��h���D����R*�ty���0R�e��HA��ʚ%#4]���h�FF>}�&���L�b]�7��=�0!�@��{�2&��*��S��([�;1�RQ���e��7n]����:*u!M��F��+��1U,�'	=1K52�+���m.�- �'���Q`�fȇ1�m���d��5���JGkf��{3����U]��V*�>!����"*�N��QkS�x��Y�l���Gh:�U::x�Vp�����0��x��-�H�v�68]S�B�%��������b��Nׄ��G��tľ&�g�k]9�!K��e�F����*�e�Dz�2�ˋ������2e@t����W
�z���_�h+����9xz�`��'CV�)��c(�V֟��]48�eq��%���+�t��{����;�B�w$�:^��ޕ����:�tQt ΂��h��d���֊X�_B�AY:�PJ�eX33�&�R�%7u3�ct {-�Ftp����u��[pka�%J�q;=�v�wwQ<㗕b�m�L��D�����f�f�0�8:Z�z��Cf�m���AS�M�]��ΏY��.���O�����-��m=#T����w6������.v�KB�Otq��s�qa�CB9m`�ܘ��%��+)_3����H��xb��8��U��UW�*6-9l��"j���o������I��)��Y��2$�y��]�jɼF�fYz��56e��@�Q^\T����K��z��K"��'3���oA��NT��)ψ�[�_aԕ��BU�B�rӺ��˵F�J>�moV>ٔ��դ�q)fr�L��b����˝5Ɩu��p�±�;LО�-�̮��*u9��Gq�dӣ�8��Y`.Üw�w)J5TWۉoX��-b͠�#D:і�F� �}�����Y�%g]��	}.��e���a��´�`g��խ����V�SMe�E�I)�]t.�|s*ڹA��1̷�o�7OP�U�����^�L�41y�N����[�u٤�/�u��˞�UR�N�r0��rt嗘�֍��WT�B�Y���Nެw��'$�TsQ�l4��`��Vl�S-k	��
�E�VK:;��K��e�Ϛd,ג��@�/d�t��]l5��WՃ	��:ޝʻ��ė;�}0`�.}�/���c��&�<q�
�-��.SPKKt�`ĺ�J�#�v�ʺ�b��g����7��u�T5�7�If�p��`�y�GB<�_v����c49��x�ps��u�_�]h1�J�]I��i�c�l>5���M�4WZJ�a������h�@�̋VQ�H��8��6�)h�WM��o˾�L��-�su�����`�6�A7WfE�]�OO(u�o2���L����P�S���zJ��7%fa	i�}}��:/�j�-�Jm��ffY5�>Z�8�0TL*��^^`���ü�ʻ��k>�M���msUي ��ƺ�Y�vXО��tY��E���DU0�/V����]8qɫh�r�L]kqv�T-m�:&RNs�je @dGY��뾺͋"�ܧ}%�wV��^�#ɢ�r�<SA��}�t�1N��9�tV���g��6޼8D�@�DU���P�WY���H�̚mL���&��`\C�N	7Ϩa/dS�zw;����M�:;2�n�Js��l�w�޹�u���V�	*���ˮ���i��̝[/y�r�z�LH�l�WAV+N�q�Wc�ɤ��&7�,�����_NdMl:9�e��{��M �����X��!�����ͬM����Zu��'$�^�I�\l����o���H�&�"*�Nf|r�� �������mR�t(q�횝a�6�S\*J:m�ٹ3\�B�&wl�^4�)������r��vmn��IcpnXc8����< ���E.Bb�,�n��M��V��4.�����Κ��-�2��k�����1�̪H\���?e��n]��@�m<�Q�]��܆L�K���\���e��5��l4t��nf�w`�,Z���X�(��V�8%�#�8$ic-kK^�6f�8(+j��J3�1\���B2�Z�[``,����G)���>Tq�҃����
�n�l��Te+���1�*��a�o��oR礘)�����	ӕK������<�	5׌��{6`�۹*j妭�[b2&����CY�59#��z``��2�l�����׎sr]6�c1�H� .��{�*���7�'��<s�d��97#{xQ�Y�k�h��@q|	�;#1v�6�=���{N���2��"|��ܝ`�(���I�Y75wS�H렓LCri�B�2mg#at/:ڮ��>ݼ�V�_v�dَ�T�1�fd�V���Tii�%V���Y(�t�c�*�mӤ7��Zk������YOH�wg:�[Y'�Q��nɜ�ؼ��v�o19�U��%����5k�5������.tz���ڐYYG	�o:�d�����f�:+:��y����.-��d��궉�V���_	=���Zv=�ʓ{u+k�|�u>��%����V2ihE�d �5Iա�u�� �7��3^���v��j�׆N¶�R�{ci����R�m݄6�:�ۏ8y��S��L�RոR�(�Ye���7�B�p�9݇3bd[tԊ�C�rq�:���N���ӭ�}B�=��}�)2�	^�bf;��U9���F��A��y[P���ݲmC('2�+�P&�y4���U�P���nnN�&���{HP�ΥVF2�*���Q�X��J�-y�]$��ѷP5՛f]N�^�.�nE;r7��9"��+���y-� ��w$�7.�.��C82�!5�!or���n�,���X �A��Ed�y�^ob�������Az;U�ﻊ�8Bѓ�hak�r�Ҳ����%j�k.Uyv	�VL�MW���xE�{L�检3΂0]�]v0I� �����8�Vpɻ"^ϲ������*�/a[P�KH��(]r��׹���x�Y"��U2_ot��T�V�uUwy�ĝ褋�#a��e��D*wu�S=aԃX�������gr�T�d��0]�˥Ɣ�*˧ưī^6��F��<��[5�S{��5�`����4FK4����fJ��pq�@�����V�9#k��!�����R�eھ��tN�̓x�o��l�������
y5��I�F[���)��&qd�?#|�����f^fP�#EwL�T�q�|n���7+i�z�d[���|�T�q}Z�ڵ�����g;����I�U!����}y>�mT��Vf��8��ιl>x��@�,Z�%����p�ˤۧ��ϔ��Z��Ժ� ��*�rY�+E:8���v��}y܌���+�r5�6\���ʜ�]��#�H�Ww|3�bPF�1�HU5t�����/n�2��f蹹��N���f�j�w:"\9��B�`.�ΗDW>7:�:I�������B��yZӝcH������z�,����&-��sn^�h�C��%
h4���݈K�N�����jDx�6��If�<v��i��Tp^�mU�C7��igI}�R+�DYƭ���m̝w8������$�o#!̸Q9C��>Q��B�a���;&�[u�ҹ�,cb9K�' ��}f�:)��S�ڑ���k&,jK��[Ξa��+F�NǄI�|�%lK<���a�r��fN��vS��������T�A�K���V��>�O.D�3q���=�&�c5���ɧF���!�/p+�Ә�e-t�-������;��0:��e`UU;[�/y���aJ���u�-�{(n݋��n��h�1âh�W�.s��mIF\�w(�_Qb8�˼bmWV�n��z�࿱Qխp���c �����kw��>��;�����6��o������g������~>��>������/���q�|����ww�K�)����r���p[~�}ϳe.]$8Tv�9��J���q��8`٫�fq���i��I��&V9E��O׺� @-dXmf��78�ELĹ�K�w�����*�����+�ČR���� ���.5��Y�.����+h�-:��3\�+%D���z:�|:�Ե�Q�7��n�����m�W(,ޒ]uɲ�ZN]F��lha�0�e��]d�9��X.�h�]�fʸk��6A{�ڂ=��v�J�ki%�Z��(ū��e��p���n�DbxpM�i���`�p�.�P'�y'�w��zGn>�����C��vX�d���c"L��FK����]�Z^�혮�-%k۰s� 纒*����}S'�/Me�u���mv�@�ۺ�kh���c)=�4}`�킯�����p.s�}1��r�Ů�����]�bsrS]��{��JЍ���gX���Ϊ�4�t�v�ˠ��݃�N�Be��0�s�"$:�b�%�Ƶ�&��r�__+s���Ɋ5�~�]�ANė��8�=S[n`�wK���Wn�ȧMw�J��nVkm�(�����^7��MJK����̙��o]���\Un#�0�q�y�����W>/i6�mVӵY�RAB:x�4=�v�6�nv1Җ� ��ιΆo(z�{r�o.�T����t���R�����S�[���s:]�o�$y#�'M7�o�;����$���E(�nǜ=swqsd�x|绗��_:�����<�eGݔȜ�N&I���K�p�g����:�R��ZS��H�5j�"�q5ys��)�NL�D�.���9r���s������+��RT�ݧ��E�(:l�a��r���N����u��ȋ�Pp��7'Y{��BvAz�e�K��.Uz%&&g�9�S�9_U����yI2�'#�D�b�p.QI��r�.]�".FWny�z'4��\
�ä�a
����]!�p��/;�o:ĲI�D�kː9�	QY�ˎ�s�<(���!�ԋ����S��o:�;�˗U���"�����ٯ�ڡ��rs*agH�]r.*TAt��u��prJ\p�n�C��\NҢ�2B�8��'��s%<�Ф�E�8���6�B(I��{�<9,y�t�p�����Dy9�1B"��T��{�t��+E�UI�h�O rNGs�Ps�%W]�(��tL*<�R���Ԋ#�;�z��RQ�Y��=I��,C�B4.C�;V��Ւ�r�.���Y7zWT�D*��@����n՛�Pkn|���$���UG�)��ڶ߭Y�g�����ǲGX�i��M��vie�5�zc�O)���<<ӛ�o>���u��/�9y���l��D�2��ե���lyV��@��AU�#n+��� ���T#�蒸������^��9�ټ9D�Ž��6'�`��B��E�C��Z�+�z���v�Y�6Lt�������<��L��6 ����>y΂��ԲJ%Ƴ|+Cw��<�G5f�{g{��{ �:y�y2�40��<��K:L��]�Y�eJ�=��.֮�qvOI����@��X���ܽ1q�{�F�
�=v��>O��h�]ưZ����p��E�%��W�p3�� X���:�(K}˗��r��n�d�#oضֶ���~>���~�҂��z�b�״�A�z��vߺ��ύw��B��;��Ч��	�	9���琿[4��ޱ)l�\˃�n����=S��U�ǮV�@�q!1�%�Y���KAq�\��R�["���Ȧ������e��"��Je���3��̥%�I�zE��7u:+P衳{J�Q�
��٪^����w5�=鮱}Z��%���k�U��AX���_1��3�5~�><Կe[Ճ�y��D�C�R�wG�B,�͵�޼Sǒ�o|^A[�z�Zy0�N>���=G�1ߑ����W�/|�2v�zf��Ȼ�݈���<�1��g{����oo�;ҍD/�*і�moH�<�=kF���â����[`H{>>AZ�6��X�jF�QJ�Z�}�p�t�ޓ��`+�� ߒϫ�C܂���
�%iU�v� W���GV)�@���GH_�8�cS�>�t2����R{�W=��?*���x���h!���0v�K�x��efOf���/"E�bh��"���V�z��y.��~:T���W��ru'��Eq��˔G@�A	T�2����*���}��.6j]LÝz�Ҭ֒��(u^�t�lz����.;� ��s�r�[�v��v��y��c�kUj��mtQh��6�g�Pmh[�׮xe����)�U�����phзz��0+�U��w�úcKd�ݓ�3(.��{Dj�7�2��
�;��.�>\�V��n��=u������<�ڍ�o��Z���X�X=0L�x9�{~=S���<����)��BT�w��*	R{������L������z��7��v{��~���n���9�ʚ;cΪ�m������A�����u��ٿ�����.��*�#}�U�'�<��v���G�;�V�g�����X��nMo��݆�9E3��.Ǽ���<���q`炛�t`���u}��XF�zu��R�z：wr�E�o����F����J��؎����I�(�k�_�PAk�~[��?hN������� �l�Cf;�1��z�z�����m.��@}+�i�W�~�o���퀩 s�����jg��[��4����ޅ���������D/7G���{���p+l�ښzz���<���Z�v׬6�pC����TV{���D���z��G7��!#�a�^:xT��Z mq�opWlcDڂ뷔������{�0�Xx�P���l�c�����1�7����	r=|��+v�dz�(5Wݠ(ĺC�CC/�g��Ωף6mխ\Un-c��7%�z�z��o��+�wQ��q
�*%vG�f��I�� ����v~GI�K#� �AJGQ��B	s�6�Fң^]�c�%^lM켸+5h���N���v��(���L�U���j�I`3IbG�����rV����}C�^Uu�j5+�.�ᣬ�c�h��z�(�+���\Nm��Ùsf�m��B˽�
Zl!��ï���L���g�|�=�����3h��=�@��M͗���+�;�O�";���<�M��U��{���3�m3�۾&I����]�]�����D�6ȼd{Z���7�'��+�rO�ߍF��Ҏݫ�IB|���IM˃<����������?{��^��%}H�km^X�-�y{>(�ϩ``���
���w�I�}7ϓ���{98�O�Z�"zg֩�k� ��A�{�'���*�l�g�����37u]�A�c���x�t��t�:������J�_F�G�߷w��#�	E�ɵ�S�Z�h��ۺ�87&�D�i_u���!IW5vŻ��`�i�&�a��&n#�r���tZ��S�fuK�7D�w���lp��ѱv:�}/�U�.M{��,���tB��B(�{}^��68�(�}��PWV�lv%{.�{J�����T��|�UX�J�>���K�R��m�r�����jt�s����-�=�V��[�؊���9}�T�'���'�*���߻>/PU����	��ݗ��A�a>�����a(g�]u�q�l`J
���wmW��vþ9�z���~|���������l��#�{�&���'���Hº���K��\���[�������-S��k��}����>ݏ����GO0���ZmJ�H��RF�RB�H�]��ό�XQ��o����w�D�s��ZY��^�������U��b5�n��$�ʻ-_���:��/���n�����}=<��}Ð�X>�w_t���<�K��!�WB�a6�ޛW���=�d�X����X�Q{�u�"��t�!��0aǻP/i�B��c�����F��������&�U�5\`YzSh%�	��<�v`Xg/������nl˵�����s�2K3 ˕������)�(�-OkZ�=��}J�,�Ӯ�/�֚���#�uLwv�A��&���Y��+��Q�:����(�����*_<u.�R-7c�͓�"�Eb�z����z�-�Q���_�~�y6���+̢��Da~���T<0-�"�^*אy7�����h�m�R��"����΃�A�BnB���:����Ի=�OzJ�ΎG]�|{g�����m�W��Ϛ�&
�C����j�ĂnG�T�֏R����%=ǯ���pg�S�]��Lz*_���D:h7�e�w�)o�K�?b_�>Pmc ���M�9$
�<�M||3�S٬��͜���Ϥ>�[����g�
�,���ش�6;���KJ��ILP�g��'��,JӨ�
E���x߻���J�����p諮�����|�[��#�Y[�:w�{���N���Dǽ��*�+}�h�/x��?v��=\ÞK���@�ݭV8�
�Е�l�џ)�ս�(��{��z��Gg�p(�=�t�d`k�Ө����}�;��J������y���LLTZshms�`J<���^lvm�am�坶r����q��3`�,i�#:��no3a�Y�3/�Vr{��ӵ9M9V3b~Amh���RB����5V�ϣս�!I���U�Y��z�H�!YY�Of���^D�z��#D�V���l�*v�m�g��R�Z�e��o�F����;ލ�z��ǖ�º��R�<������;6���(�^�
�*({�%�m��3ɼN��7��N�x���$�A����@��{�k������"���)�/��Ծ�߲�s�x��O��J�w��u�ߞ���y����x7���7<g�2��S��G��=�x�>����T|����2�?o�2T������a�qd��19ʷ�?yͽ�=�9e�}@@�r��a�k�3�c���z��f�>䩬k�uU͇�SWŕ��b�����Ώ�zh|Gb>����_���㶩
�#cR��)�maP}a*+�/|pGD~Q]�+��<��iוf�R$j[���L5U�ݾ,�d��wp} l_^Nn���*�u�B+�`W���v�	�y�*���+Es�s#���"�ۓ���o�2�C.�Uw�3x�.^�*lŏ�[ۢ!���a���:z8�#��b�*'�J��v��t�K�:o�����W��Fo��ZAO���oW��Kex�!@�}yy=��g6{��H2{�)9�ߎ�w� ��{������3�%�4�w��Y��7��c���Ad˜|����fA������ɴ�jں�s(���9���׬�
����[�
�	Db�w�/ ��Tl�سٶ6�N��E�+~囔�Oә�_��aɐ{x���9�i#���f�voU���1Hw�����^�<^�ߗF�� Z����z�Y�K8�YY�Oe{����=K<5/K-�w�$lx?�FX�����1C��ZfB*��RxZ�vDz3��N�f�#��O�v��!�v�`�w\iaQ���R��e]���G��$��7t���::X"�y�t�P���U�{�}�.7�z��T
l�t5<�d�k1�7��eD����1FE�J�V���׈l(�X�ۡ�/Y��#�9�2۸\^kV�.��<��	�˝��5��d�!u8�E-�½��}Z��EG)v^�G˯������P�L�㮎��d3���q;F��g
����&�Z�~����|'��DO��D�l� �C�{X^�y}�gٱ�3_,ۭ%xͪ��(z�J>���1w�^��{�[���}��3���=]���YT�#X6�w�,���^�Q9(�� ���(y����K�W�H�����>����x��JD�]z��ԥ��i�T��֐���~�^�B�:�A
<��gel$��u�M�4G����lY�Gw�\�
[W�ٶ����z����:Q�i[ޜ؀������c��n�ߋ�ﵻ�s���^��3���]c��K�zx���rξvA]%vJ��(��Bx�
�Z��E�Y�p��!�Kp��G;��ｍ{aH�R���'��m������8����M�Ȱ��	�U��]5%�{D�xW�j���|�}^���)X�mb�ܒP�{����\�ߨ]�2��$GF�]u�rw����"
 w��!�]����WiH�ó�r=�!�Z��<�T�l���fe�+�{����[07`�y����[����D�Q0ړb�%M��ƃ)��W��:�M��=�WG9I�vuG1��*�H����63h�=��6��HX�"��]G!�8f��vmH��eI½^����7�JͥAmJCD����n4�;�7��9D{}�Eՙ�j
h���E�:���;���P#P*Wu{v*.�Y�>�č�B�#
��v��H��M��WGX=f�"(a��Ñ��;&Nsu͞η/�m�.׭�g�`���k��l�z¨EH�M����6���崞���>��5v��tΑn�'���7/Fy�v7���2�N�Y׽ސ���eC�*��b�~X:�,��c�/aD�}y^J�:��������|��k�l����\��>��tG��^�z�b���i�����]�;5���oR~��"��[���EKA_1(��]6�y�]����{^}\��s|j������D2c�R����F `,� �@g����<9C�N>�$kҭͭi��WgUn����b�!�����|���Z�7�2&O>ڨEj甕�ܛ9���uv�l������Fx���{1=H����C�)��q��%o>|K×x�Т�n�5rV�7s"�N�$h5Y��M��;�Y��2Nt�
f���΃�F��eI:�R�z����m��M�N\Դ6mÝ;TO,����+]�Uo���sD��ױ�W�u�4�]|ܝ0}	3\��ZdԱT��Kװ؜����oԣ�POo[@;��ݜ���Y#]��{��W¥ͣIj��6R�uX�;��0����V�>�[B+�b����Yy�w�a�Z5��b�׻̀��q��W8��]����fo���A;�l��X낂�=�J���ՎׄY��1�g���5w��WY�C�/��-�0gofo^��SM�l*���]w�kL�M-��"���̈́��H���Z�1rZ�7k�m�a3Mgc�х���Q���.���B�nY��7BV��1n�Bx���U�.�/quQi��0��2{R��I��v될��	?G��9�SVN�*�@uT�av{�����^�G�.:վ�� $���[������7p�bf��]AȐ�.�^[�T�l����ZV��[����㫄�|M���3�FeL=��E�u�r+ҩ��w/x���s����X�S�������q��۲��z�m��@؝��';�����;��^grV;��+�AgWOt%r,8���M��$��ʚ�έ��vM�j1D.���㡋ł�������������G�1�8�q�����$�]����F�/�f�Zb}�ͳ�	��\f�wVJ����
�3�
�� ����Sq��2�����g>�4�yrd5m�ܲ'�^��	<����m.T��(ή�γhN��4.GK���pn����d�r��k1f5����Wwy�(��gJem����gh�	�ۨ�׺LHi���A٪P�Թ����`��<(�^<xj��3Kw���Xv�6�Y7d�ưs�6�p+Y&��;ʩb�}�Z3d[���\%�����g(>�Ǔ8����Ѣ�=�4g5#f��C5�\�4�>P�bѫ����Gt	�E/�Ҿ���t]=����qX3U�k�	9�6>�5�t�R�^t��%�4m�gC�e���;YT�5��3�cq��(��3�݌f@��P���`X�Ie�%*͇��oeȞ��u����vf&�թ�o�M\��땪���%Ũ��W����w��9ŁMCk�O/,��慛��bہ�6Λ�jcv3lԚ�������;չu��5U*H���n���a�եj��2˚�UT{ץ�� _e���-�W4`̆��N���rbI���P���Cr�tN��f����pX���̮U�M,T+!�{Y��v\����7z���A�ջ̙��U����Jj���o]�1�Ľ�Yj���Ǖ)�8�J�]q���7c�}�(((|Ŗ���Z�d���"̈�<�Je�h��e^�S�U�ܣ:T�VʉR�E���na0�RW����C�R�I"�\�Dt��*
rH�͑�r��S��$�ҹȎ9b�Q���;�D;�qۚ�GHA$)��:Dd�#%��5՗N�8J�T��-\D��*���&f��Q)X�I�U�� ����n��݅�Er�Ii:���R끝W�u�X�I�&r�
��/%P�kj����蕐��^BPR`Z�%�)!Q;*SL�wi���H����.k�y!r�V�s�H��ꐇ(�Oq݁����"*�-C��u�\(�%i�nK���S%��XQEs�r���l��#�Sp���J�pq���i��$>d(}W�4�jꁃ�*�c������T�p��	��pJTkw �%�L�C;d}n�tU�˓c��tʇ��Z4hd�Ƽ>�����^�Qڳ'���-y,���O�)Ć9���?_U|2�����DE/e���J��ii��.<6v�����N�m��	���p�����U"lo�\�{j������!�{5�)�3���
�2׳�*}9v7g�>{���������jØ��/T	���#����Ba��u�y�*`�#b��)I���0z�t�����Ÿ���^N�vt���A�A����>��S�|���������k}�U��E�lNu�;����o*K�Q�j=���c�%5���z`\{�UN����AJ�A���7<��0��h{�NDmQ���"���	�ņ,k�g$չnT�9O�\&��r�p�VԼ5��p�b|ύ���R��u��,�!`]s�z�̋��|���`дC�0%:��a���
R#u�c#�b��� Q����OGwݖD7��:<��/K�s���%�6�Y��<��\�/�V�w ��@���`U�U�7�؀���R���5ρ�^A�����T�� H����B����f���ٳ/Wj��{�j�3��+�H�Ź3{h����{;9��J�V�mJE�O�6��[S�kK�nӾ5�O?oG��e��tF�a����J+�h� tF��w.���T{ըX�g�p�n�腇�s�ۜ��̤��a�5n+H����eI��*6g#�
�f(�4>_A31J6pa��,d �.�鹾��������4roz}�l��Dc�� ු^8൦���<��e�����?�T:p	�t?N�o��Xc���ؙ�����I�73y��uY�zv�� ��Q��.�3*|Ǌ�G���-���P^-�(�$z\`S�dIkN3���W�oW�̴?D���&+C�*��V�}c��pI��6��N��bw0�ˣ2#�8���ᷗ��Q����ٯu
�Є����l����ѭ����_N�,��V*c}tخ���it3}~y!��f|-i�U�Z����0y����R�xg����]���g~�"�.�c�Os���d��q�7�b15~��u�<��Y_��'��1�`�(6=�d~v�T��6}��#(��BWE1 .`R��`*�sѿ.��>L�p*0ǣ=��+dDo�:�ұ���|�w�v��r\� �#+��wI���H�}&���*m�^k=y�F��q��pOro��eٶk�����r����\Zw������Z�.eY
��4wr�u͝aI��`5;����#��X�l���Vyb��R�j=tm���
Ԋc�
�:�(`�y�uFl)�6lm�����H�Yŷ�>w�ْ����EU�N�V�?X?7��LlR;o��*̉ʂ?*?��_Z��\,�_5�����4�S4��z����o�15)�G��w٨z��`i��xo���'���R��}t�3�B8iW1`�x���4&�{yDw��� �tG��ıy�w��Kߨީɟl�����*Prp��H�|8y=��3�������n�|��.���l��r����f,r�7��D���_1#�n�&p�c���.4!9�CV��W'��ɣ�`~�f�����;P��ʁa�L�Q�O��O����gw�Z3~����G+��E�ec��=�V�V�F��<P0f�+�y�-����3�&@�#]�QV���5[�Ņ�{gJ�	c	�Qt88r�����t� �F�N���cE�JFtY��I��؇�::���/D���D�_D ��P�)X/�a�|{����e;�Ό�uH�-f�z���,��@ǐ���8�J�L�*_p���v�߯�0ܽ ��7��P1�7��<���q�q]����;,wQk�l,��Q'�y�4<��ai����0��R�B��7���전t��Lgk������ �n��6�^�����꒿ȟV.�S�=�ޣ����}+iqe��b��8U�[�Ӻ�vDǈU��m&Ʋq��Nwe� ��9��M�qep�=���.�z;���1���7~�1�"�O�i		)�b-�l������ұ3(k���H?~D�ˢT��9�[�=�iQ��L��+�v!��K��Sbj3�L9�߬1���E���q��mK�Y�n�!�3^^~�����r:���$�ٍz/�����~�W��x���cs��"M���X��Н7
�⳷�׿tS�~7��������$�n=�Xp����1!%f����o�>�ɨܝ��a�Ň"П`������>tc��Ÿ]�;ٛF}��xy�|đ����ڀ���a�0��ƭ��+8���|���-��Ǉ�tǁ^_����S��U�yԚ3�xc�-�^����2j�K�r�����K�̜���~��x�\%g�Jw��S
���'�ͅ��.��Կ����T
�J���R'"s�YTP��/1�{��J#��h�	]�{-X�F/;7$U�Lo�҅��U&3�"�K�w׵t���Ax�۸k���&��+�\z,S��v^9z��G������s�k�e^��L�#����I�Y��r�۹�N��-�W�RK�΍vh��w��N�FJ6��5�e��ݷoޭ����CZd�F��F�J[�s�6�w�T�%�r�b됰M���ں�p�H��
�-;��h�x�ʊ�P�l�}"���,YAg�Ud��H� ����9=RxW�g�,?�x��o�����_��Nm7�1F��o:|Y��|��t�F�~���w3�/9Y�쨂� JJ���4&����c���f;����ܛ�Z�T�6�M"c�}��t��e_��ϊ�1�.�'�<�}<�<<���(�՞P?^�6�����|�$�s�����k� (;
��$��w�U�Z�Y
00�����J�7�K�ʝ0� �����Gk|�A̇Vm�����%{��Wݞ��p�lN|�Pb�h�E������YRv<-�4.�=�n���>�l�8a<�%���\_J/���.t5�Hۂ��9��z�� ��1�5j�J+�pA؉��x�㩃�W����)i��S�3���g�2e�`���� }w�ϙo2g�u�#����R�=��P�:�����	�u�Ϣ�W�����*�
�V��g�t?~��蝾�`D{֥����\n.�pf5�A�Bh�w�t<7��c}8�lҜ>�a���U�~�a�,M��xb{#�P�{�JGS:Kd�A�*j��j���n��F;�#fw�
�t5�Q��;��MJ�9�G3��L*�|��p,�z?�ܓ�u���綞o���s�^�g���s���6	��u��pJ#!]�WIX�;IT��+&[V���w|��$n}��qB�I�&�ڍ��t�=��N�ep�v.�q˼�.��hlrF�{�6���0�?²���`��l�I@^9�>UV�3Bᐚ�r�p�ڗU�AM��|ƌ�����=q����S�2q�s�V9O�lb}f�ӧ&eT_z�֡OOSۗ��}=bl
!_T�N;e���1N���b��878]k��!I�1� ɣ�ߎ�!9��\����ϑ��V��6 W�/���@��MC�'=y~�xc_0Ub1�4;������QDEݾ���4�[�ế}�bV{�$o��C�9�@A����y}�F��(���u�(m��r,u���`�^Y��+NLo���z;���	��"v}��� �=�Yvq��ǲ��r��#�zo%��r����D�pU��:Q����a��Oh����;�dAkf��UGy�O��A!���[
,T�y�tɞ���Qϼ��~�� 4��sfp�Q�p�UX&o;x�h���_	�Q1:'�0�
�]]/J����pI���qd'z�1;�q\9�ګ��������o{	��/�uzn'�	�(Ϙ��4�����/����ՙ<���\��0	臍b����F4��M�g[���9�^f�k>�C��۹d7v���pѭS��U��ϰ>n�;���v�αhatJΜ\�\�$��	��,�� �KtwU3֞���H�W>Ӑ���W�Xj5fm:���̻�\(��]�ts(����_����w�����\����`����$���_���S���넪^b�OӇ��n5�֘��ǝ2$g���8�߭����'=װ�#"\���B����p�:�F&!�/WGo#
�N�O�Ł����у�0�t��t.f�'����Ͻ��+6�F���������磼��%���V���Xf3���Q��p�2�=��ܧ�cwj�쭏O"T��C-E{��N1�Jp>??�Л���#_nDxA�?5�4�ߕU�zk����;���o�In_���>�D������i�#�P�v����s	ǎ���k(�=q��t�,nct{[��
+�F�N3횁c��W�1^�(98r�
s�*b7�˿[�Uxw��QS^[��J��ঁ��1c�.�3xQ�3H�E$36*P�g�.
F�e`�K��m��f���S���1h��0/[3q�j�joBw�P�5�P-�L�P>����'���if�b�T��^���d�q�#!zMͩ-g�jߥZ��<P0/9�b���7:��r��[>��:�������G
J�z�<�HA����;�墓�ۛcR�3{���B���{����p�����vYG�pP���|�N����ǩsu2�s]�I��aWq��s�]#��包W�1���r�5�f
��dЕ�j\z�Tf���}�g���|!;)T� G�Ѷ K���ÖvX5����Ӡ'IN�ۤ�vr�"��0�l�ץ�X9.���w�N��c�@��} PC���Dy��70��Pg�x��z^�C�=��{^z�������.����gT:hw1�^4
�A|<®�W�U�'o�0ܲj ��w�*%;�W}ԹGe�s��Z�ϊ���®�/��ϨsW��TI���I��O��T�Gu$ �z�琵��"�:����a!8�!�U�r����.��B��;7Z�F�m����� ��C��,f}y^���z���ؚ��)�4߬1�4�����*^��vq�ؽ�68��jG�h�-P���-�}�r�ֲ�a.�����<~�[�x�������ŕ�� d��|�����`~7YR��dM~c�c���X�г1��_C{}� �N7�*Ç���4��=��jΡz{:�L��߆��=�v=�uP�V��R�����E�>Ⱥ���`�يY�A�՞���\n��F5��R���Ph������v��ԉ�C�_��ȃ��uv���8�U�jIk���B-�k;�s)f�UҮ�&}R���B̸���W��dz�G��K�=�7��5�!]9��-��5��+X���4CJ��`��_:L\�!z	C�ǭ��l֠r��]�]m��S�w�%�yA%�yd�V��Мvk�=·*:I��m��I;o���� ;�;�Ԑ��~~�>��ӗ���R��y�k�Ma��wn���}=��#۹��>�ə��g9E� l|�1�P��j�3``^�r�{�-�~k!�ώT�Q�Q�":j֩!�غWnC�:��x5������>9aB���ו��k]���Z�ƧJmT����w+v��99;��a��1�%�T'�|�@�D�v^9j�`(ԽcO�}�� aY9���ۥ��m��^!W9�3���_�"�b��D�����9���y�=v�w@��s>�Hw�ό��;s�ը��� J�'�>,&?�P4u~3��H��9��f���v�MA��?��8�tr}�_��Į�b�BS�&���Bk�5,��^1Ƚ����'��#ә.�K����GX�iI�
��'>*(g��ϗ	�Q㢦��uL~�h�쮝��y��ˤ���27hP�w�k�zZI`�}������N(1b��\g�xz~�C��wK�
;:�4z!tf����𞊏�!�qb�����{�R6��'�D�g�׎C����`=�Q��k3T��9S�#oѕ�Z�Nni��eP�x�g�u�uxFZ[X�����K8z+ªx��H��=���j������dI�x+w���Q�R��e
Gfégim�Z�^K�hWb�=��=�������jۗ�b��Cda�ާ��﾿ZA�{o<=���D�׮p���7Z)�ń8�S&Z�*}9v7g�~�	�/�o�j�8��q{l���΀�>^^�9�9�Ui���
I�0!e�a~��>���[���ߨ�$T��n�A1 -B��J؇��9vk`}�#[���[髝�L��ip��ؤc��I4P�%��1����a����ڼ��<X�v���0ؗ62�K�L�����NE��6�M��?²�BhU�/�6���V�S4� ͌���Q�1e�zϟV`��bO�����EQ)��".���U���ݷ$*�r������c�ƯfsZ�@�;�a��9|)c�l��d1�x?���v�ڜPοF)�'s����\g�������¨��F}�M��9��Y��HО @�@Wы(SP��� �Ǣ~��T���qJ﫟G1ԌՌV=�
�g�g`�U�1F�&0h/���SJxko�Ur��.c}}���~3f�X�J}�2}Mg�ySsѬ�ɷ��yU�_�����(W������4��a;���E��`
����9db�2��T��B|�=4��{�J�R��޵�0�6�)��{1^#nq����	�$fbi�q��u`�m���;�O��˼���y�K<E-�	Zi�(�aƯ;A�����[W}��wc-�E�y|�gM;N����Q���R\���y��7�mR�xE��ct 5�9C;>s�����7�s8ث.jumh_@��c��;n�r6�I}I+F��f
��ͮ���||�t�oh>�=[V����Uv�SB�<������e�0�ed ���8��m������onu�*���W!ɔ>4ށʸ�[fam��z�j�Z�b�nvG��z����9!�P�Q6��K*p��ȕ�97Z鋖��>���4�f�3�n󱠕�IP���{�m5���F����88��#u�O;{�5��S[�1�s�%O����9r�J@㻆H�)�pC}*��ƫ��(itž�a�H�]͘��˶{V��Yx�B��uTN�7�~�c��slg:��!K]�K�(]�A��<���k�����^e�.ے�mM0V�mc�yc��5�#}���L��M
����7��!c��Ey�]�7P�;f��e���cʉ9g���l��Q�x�G�E��m]wA��!%��[U0�i��j�����ϜgpǷ�iUL-{(,�F�F.�P�̏�;GK圆�I�1�}Ɲg0Y:��3��]NOjd<p_g]��6;s&�8�+���mT\�%���x͠�'�nM�E,\G��Ɯ�Z�y}���Y�ޑ@�ULg�5�_�3|���()���]]���Z�P�bI��7�N�*��/+o���1f��c�9!D��V�O	�{��X:iՂ���б�W.*7���wO��m���7U/��c6��Wi�:A6S��k��K^<Е���֗x��t,��{�����#Ԙ{h����=x79ќ�o��$�
�T��R'�Ou��������ߌN���k��%
Q�����e��XQ�i}5�:����'KW&��9u��̛9N��ʸk0G��Е�ա�&��+�$G��{�)�t3���jCo��&>���� u1�bڽ@�w������ݬa�$n�z�܍KL��#Qs��0�racE��=!o���Lg@S�|�-j�G�7[�K�i��%�U�8���mY�H8(��䠧��V�eG�<���=To��l>���2���I��AF��Ց�H�ۭE(��Y.]ۢ���I��H̜(��>0p=����H��]K|f���sE��ʴ�\u�gzr��J�q^=aC�ݠ�PhNA,�j=�3:��P�{[-�44>��d��r7@�k����,�X���y����v��D�_k}�3����>5����H�s.\�5�.�Y�'el=k2Rb�A}��ێem뒞��Ss9iNwk^�~7Ւ�&���%�u5�\�|x$�'Q8;��RO�s���G��s�����_���	Vr�(��ٮ�琇*�
��s���0��� ��T��,�	'(��xusp�������y��BI��*qd�d�ܛ�)-���@�����9q�B�n'����r�TG]�s�N{�*��D�QWU��J�ԅ��d��'9�����( �EQ5s��������ruNҠH�p�Ws�$�8�n�^r�Fd��:�	�Bd�RY�z�;��!���e*J�!�<D�u���Y�"��/utN�c�F��rL�w<,���B{�N���]U�9Չ�V�wvnf$�#�g1�]��*s��]P�����7Yt�O&k=�<��p�T&d�q�{�+�G�k���y�0�gY؄��������J�!;��J���y�3�B�[�5+'%��a���NJ�S�{�wo��333�>|>KVoj�܁*f#et�>YP�+ȗnϡWC��k��XaG`��pT��7����M�o�

�?�Lk�9P�ז�w�3�X܅�CW�����n�Gn�ֲ�����ѓ�)�Pwںd��l�0=:&GD��"�Lx)Q�t�+E�����8$��qe;�06y��s/p�N<�eI�{��h̋�j� ���αs,@��c�/-�~�~� l/o�H�|Z�}w^���h�>�����]�w(�`3i�cw�b0��ltc���]B�w�B��
����ݱO�:�Z �3r��Fz1�.�7�`yRbF�b`o��bj��T��K��� �+ư��"^��wz������K�]3;�^v�_Vz3�0�B�a�����9�Tv}쭩K���e�r%l=d�b!�T�U�Lp��1��
�39&����U 1��V-�b�������~�Z�1�Ǳ��m~�xS=??�?Л����ۑ���&�7:��˱�x�@!�^���~��=�L0���]{�>��Y�G�a
�]KbE���M�!4��� n�}7}�W~�u�b0��jˏ.		��4�ڽ�cS�(0`��mD��{E��
����13c6��r]� ��o+�'���z�'�ݚ!s�
QcS�e�F*rit�t:]/�ӫ;F��i7k��%*>����e��uo\���Z �%0\��}&��zg�^���?T7�lc�3A`UF�LG�j���b}�JI�):��w��I�C��r�ٖ6��ɋ�i�h.���4X�1c�U����ę����bC3��%��q��\;�Wz�9E���+�=���B��7���!;P���C�d�\VQx�"��j���+�����C�'f�z��
�9Xe���U�������f�+�}��	��?1u��_��Z��f轑,�(p��b�Q!K��r��<�c�O�9���NR��Q��vS��z�?+S�w�*�(��)��@���D��b�	���� ��o��Y뼋�%x���Vv��rg�7s�˅�4<��V�\�
D��j�dתa�~�ui�Ǩ�����fc�Aa�łD|�Z�ϊ���*��xNB?sW���}�y���W�ׯ0w��V�����Ͻ��s>���vۆ�	ȁ�N�5ʂ"K��?�7Qk�l35�P�:�B��WeyU���{�ڮ�`��3�wd:�{�^W�v4�38;��5�L9oh1��?�C���]W�1^��1+�[�B=�ov�D�v!zr'�~5dxh�WW��W�:N�"�{�,jՄd(�ING��MAu�u!���Ȁ��z�+#�K�#sh;IV�d���u+2*8�F��x�f^�˘gi&p*
�y�j�l�+ػ��K�* > z�N
�%�W;Rz�&�W@�H�_����m�ՠ_eǣa��]LC~���oU�~wN�c�\�{5�ȗ�@��YS�9�L����׍��NF������6��A-ǀ6_O�gc�w��5�ǣR���+���E�(��TQcÝ��'신�v��G�w�L���{��qE*�^Ô+��&��[����tW�}8:{�Nsg�6 ?NԷ�+��:Л�Qz�ׯo��UQc�����)MM\5/�d<�5�I�20N�Ӝ�<���~�:�����R�����9`�!y
�V9�Վ\-��߀3Y |r��TrVN�"�t�<�f�^���W���
N1/�"LV�QLQ��,8K�Ů��23��S�L'&�X�aó����h<D0w��Ll
�`S�	�_:%A��t.��/���K�3�O�a]�+�fvAW�~iTN�>3����~��Td�="G1F����"_Iϯ�#����Bps����u�׊̫���̻])�S�+���*��bH@1EM���q�j�gʪj'�b���'��������i����[��Ȱ
��#1�q��p�s]N�'��R����(v�JS���|�P��-�3e���A��}2��PxR����/��4;#��TrΈ�ǔ��a�AI]q�Sfӣb�K)c��l�x���}��J�|j�t9�S�����P���J��Ӆ]���n!b�0�*T'*J�u���ɮ�n>�WR���,�کrp�cM�$)���EP}EV|�M|tT�w�O���y��$���^���Y�4�T�����V!/�vz��]6'�Xh�F[b�4�y{;��Txy�x�5Iv6~cj��pz�$�1Q�z�X����~k�:��8Q��yX��b�2�=#3c1�I���������U�Zf}����������F1��5���,�\��_On���us�R����q�6�1�~��������������'�#��x�şl~��g&h]�d�	#��\ŪϬ�-Ǵ@*؇5��:���v/&���L����y��8��_u���C��.�Bq���W��&�r
���W	Y��ϣ��s^z�TGz�tB�0�g�K�xv�������z��{�	5n[�3NR��x����r�]�8�H�z��?��Գ?mQ6i:���"|\�w�̌��<n|V9N@�gށ��-�ХaI�p�،[��Y����,��Vz�4��ys*`��]�3�ܛ��)[Ƌ��T�nwB#
��}>BƘE�D����:�nUp�쓳�((=�۳���<cX��Z�XR+t�Yu�6kY6XG��J�Հ���2������5p�hX~� �W��{�(\�O߇��s��ʼ����z��`^����P����F)�'s�ɉ��`Mn�*��y�w���l֩o�̈́����y�#bO��~��ŁR��c�����FE]�LVv������&/n������U'���>��*nf4����	��m��'�s�7GM��`�+^X����F�nLh�S֥�����HNP�Lh��L����v��=�OH$9���8f�aK3��3�<�K� ��]Ӡ�go֫`S�'�m�싛�}x���
b�ʁ<'�X�
4T�yN}R�x�s���CW��ڤ��=Q]s=��썽���Zk�V�)�|Qx??����/�t7�ę>^8�/<�����ih�����Ɇ����ap�S������.f��Q_p�<�ۛm����-�.�g�^��t\�����ԔA=o�H�S'~�#J�6:1ό��,c&hx*c�+�1j7+StD���rx�Q�����,^z���՝rؐ�X�7�b04���tN�g�lK�3�?�Thkw�]�ŗ�+l�7#W��� t;���̱%q<Y����;.��h�e�n+8	ߕ��wu�dY\��wOY!�"���U�
�ӉS���~�+A���Of@C��yF�u�K�=��K��NG��ř� y��S*�dʣ�"�����1����}��৖�Wi$���¼���N@=y�߯�=8�z4�Ü�B�gɜ�NGg�|��JFD{q�t1�`׏>�O��"'��P��V�Gleb��}}3��39&����
�r�y��i�n�2<L� �*���A�=���nS�k�5��q�|�\F����0w�`����	4�-a^�gs�+'�t?iBH��=<�+�y��ݮ��}9��G�,!Xc_� ��꾄��37������;)��R�<�1Z�G?��p��f�9L�=�K��L��ь?��ၯ˝�mLjo#7ئ���P�9
X�\<�LY�[s�w�Կ)���b�b��sEܣ AU��'��/	_��7��H����N�js啎V����G�8�/[3q��ڛН�X�e@��b&s՞����m�{O&��ˑ=�8��9Xe��`ղ�t�Iڀ��0�q�@�]�9�VIڌ�ՄU�I�A�^pǧdM}�"B�n���:p��yX�e�� �Ѝ����3�uf�����L�;�FF#��b�)H��_DO�������tG�{f��xG��,{�,3.VR��ܑ��imӼ��\[���Wf���ԒV�0�b�R6�[���w�ޒ페�I�[3��iM�]p3Z ���-��S�|�(S�W�J,Д\�3	K*V�z-۸xm�Y��M�����\ʥ�bYOi�����͐C}�����}��	�L��=K�����Aw���L_�yp����W�%��*���{k�/h�Z������&w��{(Ø�8���y��(UZ��U�N U�E����D������C�`����7�K�گ��ow�!�
�,�8Oo����@�z����a!8t�h�E�¶���k%k����[O��2G�Ua���Ќ�k�Y��v4�#8;��5��8߬�hm�Ѿ^�zUa^�g� p��]mK�Y@xS�Z%9�z�K#6�j���g�]�ҺX�'���L`�t�D���C��gP_�ޘE��c]���8�21�s���_e���(�YO}3��*�����0ՏC�k9�l���t����FF���­���xE�l]����g��@������?���f!!N
jܽN���v�{���s�g�*���{=���:��f���Y�<��0�5�iw���n_���j_��Y>Mc��Ma��wn���"�)�.lT�0A��?�6�=2�'>)X<��x5c������5-����>9P`	��sb��[��j~V-�=wߵ!���S~X%�{��+�t�r��᩹Stft��"Dn�:ؾR�U+��=C��+:�t>[8��=�ϳc�E.��Q>4��G��-V}�Y�G4��;���hE�R�g7�H'P���H�&v�;�������r�0���^�����D�PaTG���)�Ö,�����d��WZ�`�ԭ�eK^^T��먶5Z�p�T�]"}�+�P%�D�=}����'���׭置�X\����0�UL����9u�W)w��9��2�$I�81F����N_^G<���dF]���*ٽ�]�lїP��\��4�)�3�,cV�>~ۈ�9W��$hM(��yӾ:�-��I_Y��p�z���Y�O-�G'�U�~�]�]��*�
���;��D{�nEw���=�Ŀ�+Tة�>s]2d��b#��RB����;P*��\+!G��bF`�yi��.�=��s�*�xA��!>r&�j���Ki,�wg�:��bp'����T	uSw�Q�����eT?����kt�V8S���3�����ߖٯt��G(ω�?-��XT][�\�d��[05�ϰ U*�=����7�Qg�F���0Tɖ���ӓ�o}���1=9����s֭�JQ�a���Gk�b��
9�����ӛ4��ɚ�xH�`���.��#�/uH��/m�^�6RB6����ӑ���F�b�-��3Q��k1�'�l��`3��Dw[b�p��Tz�[�B�ΰR�0�׃A
p�9�;h���bM����q�:X{�s�I��\s٢>�v��o��R
�pK8z�i}3M�*��H�_T��}���<R���TN��!��(m�g�8����{~*؇��9ߞ�g6}��4�c�+E	>���._*�C�[��r�XxK�pȻ��W��,9ӟ�"\��᧋n�*�ϡג71��N�YxŢMOs�NK�LՎ��Vf#�"�@x}C���	5n[�*�r��p�׾��nL��d�q�b{��G��;f2}[R���Dl]7q��D<]s��̋q�s�+�
�ӧ�F�*���
�,]��J��=?O}9�1_B��$xߣ��g�f#�1o���h�z�L=t�R�rZ̈́�9��Y��^Fğ���tb�JF�4���xWE]�r���Cص/ٷ�w��}MM���
��g�L�U�1F�&�O�c:Mx����ce�|�9Z��B��c<8�rc|��԰+�����'(k���[�NK���o�9=ކ`��
�,͊�R\�*� y`��@�]ӥ�;E��ov�|W����\'�7L;P"~"\M|�8Q1��>��s���G>���-�� 8 �����������ѣso��9�2���1g����ذfeY좬 ��S�������Z(*f�	�m���Jz]>���Wh�+�^wx��c��q2]�f:F�f��Eg]7@g�ׅ�z���IG�!��_�W����x���}��}�����[_�b�9z�T}Lx�$X����(��}��E��������o�,s�{�ӑ������e�v��j��`N��g~|���^Y�)i���"_�����_�ߊs:��i \��k���+�����Eg+Ja:�b;��^́Ӭ/�(��`��i*A�N_��o��hw����fO�=a�z���6$/Kὤ!���'=װ��6(S�!쪪O��z�u �@�b�a?�+�1l���]Ӱ���	u齅Ƙsѫ��:�T.L�n:^�,�ް����*��{+jVȈ`��E[����c��8�^�g�b�~*���N��N.��DN��=�g�9B��;�f(�lx��X6�bT}���;����z�;N:.L����b������]�Yf���Z��&�kwi���u����)�G�,!^��čt�:�Opz�8���x&$Q>�u���!����ŀ�,��4&b����XѽS�g�5���1>��J��fX��ܭ8��E�>�)ϼ�\,�LY�[s�]�5/�)�b��X�]xf�ę���h�2/�w�`��^޽h�
l�V�M�����3img��@!ٻh���R/]�ng!l��0_rwo���!C4r�D�A��+z<z�w�dL�A���eSDۯKm�'��5T0�jl՚6��S!�\,�ƺT$)C�^|�sd�#�l��{Y�qn�ٗ@���|1+ �V�"h�gxuݜ���ч
����J�O��j��g���eN�fk�[ck)��l�p�dwÔ)�vq�%���qֽ��[�z���J�����f)�Vsi
k�Gu:�|UÍS�2�s{�*�C��X�FR��v6��Nb����8�VZuA��κz��#H؏��$m�;�5m�&4/e�j}R���ق�=���Q�e>�5��2TJ�����
�Ĩr������|\8�gQv3b�4�7-��q���W�ũ��c�4B��yR����2�!�>����Iơe+u��{ lcq������C�T��`��#�-�4i���C��0��������nNʹ�
a'�}Y�s��X^h��.�!T��!9uk#����Yo�ƶ
���M}�p��0X�9�+q��N�����Q�����ˏMiuѡ���7�P�����A�}p�a�4s٨�Q�w��-��6���rJ�x��CZ�&�3�7�n.!K �d�֕�d;8\�ok��`n��v�CQ��	�a#�\�X�N�Yjr���[�\�X��S�cy�Y#G'.Xv�q�qP�hʵ����=�&�s�Ln��4������B��H
#��s=��c����bN�s�jc��Qq)H4��q+���꽃��zwT�+I[���T̺ݗl��6�,��9�f��mo��r��68�|K���}O��}���<k��Cכk3s��ww����^T�Mզ��K4k��Z�{f��g5�NF�]g¢�w�J!�3s���`��F(.�Z',O�)��5�����YE�Oi�����49��,��[�[R�U�;�G�$�Y��ܮ=,���Ÿ�2��(��{���4�Q�X���ջF)��e�n��7V���]�<�k�:�ی����J7]Q��1���1���
����e�dT�xy�~��sD̦7���\ң�\�1n�M����ot��������x8h^�81�˼�ͳ�O8��E���^ֲn!g(v�F�-j's�q�t	r�@�A����,m��ܑ��ةdO�T�Gt`�t�Й�Kɧ�f�lZ�ֆ��Z�w��kך]n�]��$���Z��	�մ���V3E�v�i�Cy���58Ry���k��w|���۫�M8U��D���CY颇vku�b2��7�*���r�r�����Y�+������@�=qAW/��}��b�h
��k�9󘭳���@λ%�˱)9�o)M=U���o�h��CM����1W˟oa� '���k��5� �.f7�ϳ!X��M���؏��09N%�I8:�%AAs\��-J��)t��F����ȧ<��Ғ�PC$�rr)s@��᫊�����/�(�wrۡN�N��	�H��W<�sȲ�<���<�9J	��n�Q�5nWHã�����n �8,���ww
tE�ܓ�vzU�eS����s�<��P�(�ibn�N&�8�:�I��BB-se���p�;��J���II�24q-Օ\����+ԫȹr��h�����l�������u'=�a��-]��t5H�-0�%K��dUz9�t��'R��<�Ι���*�:�E�%U��D��Bs܈��*�DN`�;��Фs�S��bẅu�ݙ繃��p­��a"R:�U�Q藪�J԰�Y&���s�?��jTX��WlV�2r��F����
��T�r�U�f�;���_t����'�Z�S7Kζ�ݑ�t6��y�)p��>'����}�I0�ܔ�H��D��!  !L���+V{-����fn5e56�,5�P=O�בH��K��t9��1�OMȓ�pv�(*p�a��,�Z�]#Rv�/��f�T5;�v*�sw����^:���`�쉡� C�f OA����X1�,�]��j�8�*��^��Ȯ�|e�EN��-�R1�c�*¡@"�����1"<�z��y`��N׌�]��Qʠa�x�f�������<�Q���*0D�|�\�|B�5���yR��|	x��w>�����7+A7o�ؠ4�8s뻥����B6��~���뾯i;Ǜ�x��AC_
�����@W�W]z~��P�χ+		ϓ��Xh�E���G;���X�\�Avf����D�è]��k�V{����ӱ�����lMF�a�{A�b>*��u0����f�ݧ�1��.0��8k"hxS������f�|3lƭ�q���?J��d���U��c{�D]�2#[>��BX����K���tS��p��?hb��]�j@�x�&:{`(��5W���A��f�%�����V�c�:��7���iq�9�:u:S__5,Τb�@IŅ3Z�p�PF����0+���cF�L2��j��Mj��5��wh�(��\'��{�h�|rD�v�`������Zd��F��bM��Rp���;�_�|>���S��)����G����JÇ��s������Ͻ9�Qd�LS
�-ȴ'��W+�?le��uy[��
�,b�����f �NSV��v�8���v�{�Ξ�Ӝ>�|e׍�$9>{+��z���zX>b}�\�@�i�+>���r���R��|��$�ŝ��*�ި�:=��I��VK����=uN3��!g�BżՎf��c�K�j_�3Y�#M�8�殇8ļO�V?����O���TX�<��>|�8Xp�m�]�df|����wT�9����(�qS����]NmT��"�M.�=p+��8��DWA��x����,M׼�c�WF>sۓ����Wy�sx�s]*�c�L��2�$O M	1J�_T�}$K.�c>ȗ�ǟ�]+щ�}�6�o=6�u:Jv�q�Q��n ��*��X���*���3�o}�_��T�G�C��MK���d/Rx�o�������x���n!b�0�o���k�:�}fJ��``�C>���>3��*NwX��4Ԓ!Wք��7��p���z��$�[������"�X�U��x��`Xm�f��H�mjچZ�L��n���c�e�".%ʧ��6�tx΃�\΢�f����eX@NH1��9HS5�/;��$���_:�QpB��]��Qջ�˰�*�/�.��jf��؍�(W�  ����5��X��u�{ELz��f��W�'�E�����ޖ��`��~��x�lNn���|�/i�u��㠗0}�03�����UeK�E\U|�(��ǩD��7=���N�#�]�Ij��\����}w}ܢ)u	����O4��_�\��U�>0��~�Z���~o��m�?����m���y�r��`)<����<u�6װN{���W���������Ǽ�[��y���"�A�������g:[}Y��,[�LC�5��.�l��pl��)�G�u�S���`����T𫀽�v}�"���	4Ñ�W��ڼ����Y��;L^o��x7�=���6h�/ԭ'S��2��{"��x}���3�jܷ>UV�w�f�ɘ�`�Z+�ݿWKZ��7�lo�v�d���`5�ATF��w��dC���=T�ENDOs��y_.�u�랷��QS�ey��V)o�A���0%:�6~�}9�b��B�v�"C��E�C�/�eI�,ǔ�]�_�����.��~�̈́������
���6"�\F4} G���1n�˼vz�t��=>Xm�-=��6��G.�����/p����t)���26/�r�V%{��gNyH%��P���.}<�ÐG��r�g^�	�(gB]p�����@�op�٠=��F[2��{*K��i���]:@���| ���x��nO�.G��WN��א|U�b�36��c�T�tL�L�
�f(�D����_�Ψ�[>{�R�c�9阃(���^����+��6ܘ߇���z1����#��y���X>�U�R��/fb-��>�W�KST�KS�*�|y`ע]�!WC��(�ݣ����;a��e������X_N��z�8�8?(����.s����{xμc5��~��*�<�������prG��|�DȠ�O	11��X���Z/�t6LP�A@ײy�;S�ęo�����1�'s/��̋p�Rb�h���ɖ LX#iF�~�B�!퇩�c��e��}�8�/�{�&��*��r��1;�1Һ���rb�i��L���:J+3r��Y��#�f��M��5>�����j�Ă��q��[����=���~�`�p+ۡ#$Qsè��q�XD$�-��?,ף��՞�2ßA�u0�5иD-�fg�s8y�?�~��{k�mm[���\��Z����c����Y��M1��U����B�>d^�5ݾ/�='���;���mY9����V#=���,���nm�4�	:�a�N��x��Y�ۍ��s��2k�Glv*̩�\�a�DI� O![W.�y�T#�XU�NGrn�۔����M$�˺g���| ��z����/ �L��k=1@���ߣVԺ���
���2l5��;��n�~�!�K�=��GtS�-F×N8�����MXƞbr6z��>��f�{�W�a�#~��l��z�����Ix!0z��֮`�vᨐஊ��V���>٨=: ���囩����C:�9a�9�B�槓}���{K�S@ǿJ�ߞl9�j:=����V&�սS�N@"n`GC�!t�1ώV9Z��1h��1zٛ�ն�ބ�B�!'�����<f�~�f?̏�Zi�sX��/C�A�S��2�g�j�%Z��$�@��ĦU^�w�B�VZU3�2>�1����>�M}��ZA��� ���aS����������۔�wV�g���c=!�zZt��h�IH�΋1�tL�"�C&�'�Vň12�d&.*�5�^5rz�'���o��z_����v �\(�hk�N��aX��*�}V�ڱ,k�NZ�wx�@��)�50�S�A�/b��9���jw0�s���/�¶��k�G:���}�D��ҹ��]��Y[�\S+�DW<'�\��jV�D믑}���OvH�OWTy�v��W��	v8 keL%�]�"��mf#}��3y�}||���d�mL����J�x{ 6��2u�'��*�Ù�D^ ���>�����| ��G�P�=3b�W����M����o��7�Z��}��Bq:E���w���Nך���M� �2�z�f��"#�Ȧ'���j]�{�cOS3�-��!z�s63����e_s�H�z���,nl��ȴ����*�?Ņ�����/�lƭ�q���Xn�r2~s�N;��.�9���1F������E��Ȝ5�3뎚��U��Á�������l9��oDJ�.b�\(��q�8k[��v��Ѝ�N}�͚�;�
�^z�qWy��߷�Ic�O
��a�>"/��f0Ib�-
jܴ�@p�^��C�`u�p�3�!$s%��>�u���"�9� *�<P�,x`=�Xݷ/�j�~&~���[��3��ގ3��������";*��D�P��#�T�39��By�V9����ˁ��.��	�lz<�E�Z������}�q$_��~.̃�'|���T���|�̌�\O�}�m�T���}҅��3r٭R�D�j4�zr.D�]Bz�
�Ё.:,
"�v^)pL[��[f��D6j�fQ*c�ݵ��FC��Z��Y�����(J�����G�S���H��ڎ�33b�Vÿ�;����w~��1�&�I�걏V跖�}I9�K"
��;Wk�}����W�(v_��g;�EI\Ԉ��;��;��|��F��ie�������`�M�����z1�&_�a�
}���Y�)�0>
�_+��~���I���O�c���q߯!��[�[��_S�����nm�P�*#���*±;kU{ڲO�����k�H�%���͊�R��z�;ӝ�{i<p�C���_��¨��]���UJ�FA��+��Q�^���0NP����jj�+Z�������ˇ���w�wې=�i�o�{W��8]��ՁCg(${�8���cB�!b�ީ�}^�o�`�}���֯��W�ʫ��q>�pJ�C(�E�����:�*Nz�&�����(��+a�߅��N�ՐA�N��O�ܽ}w�j �����DV�p'�cV�D��^��7�Q}7Z(�ņ86_B3�6������,Fv?l����-z�џx2��|͑5ߠ(���	�V���͚f���k�xxΪ�~�wh�$1��'L�_����t����X�ҭ�q�kw�u�@Fseb����~��\o�Ç�(�s=4��d����C��W{.l6>� ��!���FI��U�s�6�!�ڻ��eZ
���tO�+wܽ5��t�.=u�oG"��F������c����e�~������zsEfؘ�5�3�w7�oa��#�7��i�����%��N�"���ֺ�ݙS<�,���#h�G9ӻ�bY�mlWQ��M|����Od�S���L�������&��������}N>�p�h��-�a�������I�g���\&klm�'յ/��PU�-�GxvY�T�s�F)���;"�}$�~T����������r������ΙZ+���}��a����8㱴z���*�w�o���v!?�_����+����.��~̈́����o U�lI��@^��-ȍ�k����G|�a����X7W΃����x�1��ڛϵ��U8tL��}3�p*ɘ;������uprmLL��m��uTC���2�,����K=�m�1��Zٽ��
�2�l����{�?���N���ޭ��w�T�$�B
�����ʃ=�X5��]�)�{9{;�w�j;���o������7��Zk�[a}Ph�"h\S���N�����=��~=-�q,j��O���& ��Bqa�|�Q�H����Dȣ5\(��J,U���A�����<�7��7�c��o���~�����9�jaC.��\'��7�K:����O=�1�l~�u���疛��{ZO8;�^m��a�̞4n���d��O������^Xv.�m�@��}�[�7=��k��)s>j�Y9�\	PPJ-
ژwn��.G�тIk	V�Y��tv�mb�<x$}0Z����%(�ˢ�rݿ����k����^B�"?�:�˞�����	��{ڲ"���Lbw�bUQ�=�>3{4�m5���U�=R����xa?�;�_��}O���g}�F*lH��LC�o��`M_�xV�9�b���A��{	��Ĺ1s8�C������`:��ھ��g�i�=��08�%
^46v�4:P�k`.Y�Tv}�ʗﶄD��m�j\p��0v�z����ǫ�y��N\q�wZ���٬R�y��<�#;~�+j^�D���(�ʨ�-�'3Z�)D`�'�xQ�i�!J��LӔ�M`ׯ19�����ا��}A`�^��DBv�t��Y�����Y�!��LB����]�_����)��=3|k�M<Uc�	\n���~7{�i�+|�~��~C�z,T���1A=��p�SɃ��8��j_�S@Ǚ�����b؃n���S�����R�鿤O��,PjpT�	N|VZ��1o�8����`ն����QÂn�m*��+"}��/	���31�;.D�:�	P`!�S��a��g�jߥZ�,���5�����J��J��vhR����ֺ 7�d������|�>n�QV�z�.��.a��9'B�[ġ5�9���ћm���%aZ��82�D��#ǌP�'0�j�.]��cUmr����&HR\�p&>W0Y�����Ir
⯹��u�w��x�N}��OP �㧨���y�>���.'\y㭹�.��o��A��Q�R���)��-�R1�c�V�@"~��:�ana�3Sd�F�և�b����������;�����F3C\�*հ#*q�8���zţ�Q��5�H,N��MS�U��)�OL�W�����D{w�f{C����	tn�G����
'������лA����/����ϻ����w����x.:B�h��{��B��|o����={N��l<�f�t���t-��"ovے/+�;�fs��lMD��
z��a�U����]m�6_?XC
Y�l�ˏu�/����J܋�{5K�f5vS��|7�i�{|��ߪ
�/�a�vN��������Cx���7�6�*V}Ց4�8�_�҇ۘ��i�͉)�'��N-L0<mCZ/���b�{J��K�o9�v��{��x�1,[O���5��g�������a�,��Ĝ������������8EM[��ڀ���n��鹿#�P��p#���%[�R�o_��7�h�å9�-��M�%��̚;��YY/֕>w�����r�SV��v���݁P�j����j�S�u�T����і����f������/Fh�z=�c�pp���ݍի�7�ܗG���ȟ�u��;�j�vQэN���<Z#�i�����2�N�b�����P�9�ܕ�0.�/�Ve�;�J��6/�EM�m���]�F��e���y�ݜ�ɘ�m�Zi̙�V��V�:�JgR؍muې��	�iͧlA.�q�8n�k�p)%U/>)��F(�S����Lcg9����ηvHAc{s�m*�|-�d�$D��ٯ8���I����smh�Ec[�M{��vhh$$�����mՆc���۱��,kW,�h�r���ve����bG�9��ۄ�)�$uIn�H��*�ػR�b�9��|�N�\��vk����驲�+gجt溨Ʌq��$�T��v��L��&T���O)�Y��0Ѫ:�q������U-yq���܏�Q����5�W�XG+��/m��`�����3���1��i�k;$�w�q��q�%S���P�}6
�p�x8u-�#ocTmK�ƅ�}4R�+��Nkq40w�iB�7�����u�22��-��j^�%��+���n���f�\` �gi�ǧ[�C�7�A*۶��K����^�k*�Ǘ��;r�Y@�Ọ�='	ĶŬĬU�f�/��,c\@AY���q7�r��zV3	��m]6wNt���F�z�O�:ݨ9���eYO�l,�q��c���`}Ɔ��	E���R�Amb�U���}.������XQPQS�sȘ�^gǔ�â�u]�pݫ�����;�z}�le+��9s#���D����6��PkVK��ru
�)f�l�0I�,�s8z�U�D��m�Ȫ�F\��s���[��9�6C�[��/�;s|;t;d����m�jQX�Lԩ�c�u�����>h>��NB��Z��^L��˹C��qv��5GH������޶6;x;^m�a�.�E�U�yp̖2v
����x��EF�r��\�F�8f& �\@L�}9M\8�;��Iɰ�v��5m�i��f��or�y��)2�'`r����uح��a�h�?SM�ub�+[(MF*��7���5�ǬC:��f���)�K��j�t#��fc��j��r���Cx��3W9,�����7�xN�3� �J�u�)М��=���B��çH"d�a�3�����[�$x����q���|F�X�������"CF�c����ӛӠ�jVo7���Z����K::��kv��R�]}�T��>'�q���L�6�-X$���S;%��5YBfm��;��tb��6FE�)v������m�l<}	m��AHv�ٮ����D%��˿ǻr�b���P=eG#x*��4|�|���NV��R�GUgM�wJt����Q&�f��B�����A���Tn�u���rp���W5�e���V"N���e!i$�D��#2��2 �����,�0��*��B[,$J��+B���bhSL��<�BD�HIV$��2��Q$�E�jrDİ+��W)E�Dsd��8�B���TRI8�'���hq9��z���	a�]*�R��HU�	]��崴�8j&��u�E�	I�������q�°�<�R���'tE
�2��P�UVbHa"jR]�47R��:�9t�dE�i�R�M�Њ��<��I�q��jr��n(�[(T�9:�ŭ2��8D�I�a蚣Uv~����.�zxz��E�<zmswq�ii�6�e:"T'R�7h��sZ��ӳ��+����
}����k��!�������[��VÌ�S�����w�%�?Yu�u���aU�������JB}��pi�4����5pԿA������P��xN2�2fm<���Y�0N�Ӟ��`�G�U8ɹBy�j�3`��ˁ�v�ޛ1�b�����s%��Z��K����ϦDtБ9è�E�"�t.]��#VE�_
�n��3�F�Ԍ���xns�U�LhN�,��U&09"WH������4�a�LE�KTv|kO��l�r�J�ݹpg���'���&U�<�?P�8�dM�$W�Q��z&��g���w��S�b�1j��8�a�7����o�9Jr�cV�
��{ql	^��go�8`^���=�� C�P�)���aI���Ox�B4�8Z!������=Vʻ0�L�1,53�s��N�Ӯ#�ޭӠ"�?0���yF�,�~][�Du�6��1�*�ПY~�4��Ne����=~�!��L��xVB�:*a���bT
p�)*������X!Y��.k���S.{.����I����ʋZ-} �鮯���Eχ��g�1��Oa��W���*�{`�M��4�Xrkd���߶�ur����f���w�αr�=͢Y¶�	[�ГOj�J�]еn��G61%p���RP@���8�U�Y�����{��G;zv�f)(�S�Vi*��١�Z�5�Aّ�z�����rI�� �'�ԏd��������+��<����W߽<�W��,�-3��_X|a���}��$�d�e����֡���l������|}w��[Ȏк؇���M{�vy�gx���d�'��j���\#L~1�M�
����}lz�t��������U�0kw�]��
�0iͻދM	����cӖթܟL�d{�j޹�؜�a	�e�!�W�/Z�p�i�L"snY�=[O����2rv<gbT��ٚ�§��1. �,!cM�/7�q=3�s7�{jm>4�*ˣ'eLєٱ��5�66�و��K�5��U�-�Gu��r�|lX�����C��0���ȱ�X���UX�0hZ!�3��s��}=@��A�+���ŝW������(�w� �<�ъty;���pns��\��6�.� 3y��"�Z�!��s^F_�� ��p6�/��뫂d����V�����`éO�L�L�+�˲g���s�7=�fb������C���Ί�RV��^��2
K=�m�1�y�[7 x=���^�q���WU9]X�5WULUL�gV\�O(�ªm�����!]�Z���d����+L�&�=�i�f���+��t���/jhv>��P?5m^��U�����V��f�D<:�v`a��;��(���;�]�#/c�RY�����ݾջ=��W�?}�z� �����+��K`RT�1�ԛ�3���7��p	��fؗ�g���Y��q�f���n��=�~����s ��qO��>05�<�Mk�ۯ�|JX3NM��+=��e�:��#W?�������q�)�2LO	11���D�ݠ�଺��9���8���og���aN��*u;�Ȳ�̋]Fx?�(��:���_�쟤�8�x�!�<6�//-9^���	Թ+��z�+�r��0���g�+���Ѯh�qZ��}��"��Aw�m���BП@�7����^z�ç�:3Λ3��b7��?Qv`=��!���]�n�ؗ��:�o�X�0��68~��?���=C����՞�i�=����+���ψ������иXQ�D⣳��emJ϶�CF�*Ը�2�Lg���ᥒS�3O�L�<�;,K�#�;�U�_��mݘ��9[R�}�����nx�E�R�����^gr"j��0ƛ�b߭A��N�
�ܽ�����br6z��;���/�Vf��[M���������{�Yզ���u�o����.�vF��)��P���M��{�}6�(��vc9��ΠK�rt��N6�Ut�oN��������;!��l��J	��谪�2���^�u2����/+�0���P68�t��ay��v����|��]�����?T�K|4�BcJ��'8~SA�f([�L�E�:�W���nxk&$����1�P���4T���9a9�B���SɃ��8{K�'�c�åS.=�Q">ڄW�oR���"}���!ɹ�)@Y��,p3��7ϳk�e������Q�u3���Ͱ��<�L��4��K��ó���Ǽ��ї�=�Q��f]����������g�y�x�`͘Wn�)��c$O@�OA��OA�
\#��%Py��7(s	��V�.�H!~���b�%#:,�|�D��@��G3lu�32�7v�{�"�C'��W0����x�f��ө���<��C45�|�DJ*3�U����U��&����4e	���
���t}~���Q�/b����1�\���Wu6xM\�0b׽g�Ǐ�}a�)�b�������4<��a����q �z�	��a!9���a�zʩ}��b��p���i����v*��a��"�g��υ�{�cOS3�3t�o}�F������[�#���6^�`ސ���L�4mm�^J���s\�z�LyM	ƪ\�&�c����5S�of��o1e��+�ѱ�*�A@\�
e۾rhP�x9�69n��/t�l:�d�\�b�UVjj�v�m��oz]�ZR�V�����9��o�)˹���~2&��� �>o�i_��]���Լ5�5�J܋��٪Y����^/O�����>������s���)X}+��k������$�@���PED�b�tl�v��/*���w�AJH�0�;�*��q�-Ǵ�kx1��>�����8�(��Y���V��_�����`�iC2-	�t�� �ю�Ÿ[�-:P:*� �{Ԫ��YO+�w�} ���mSW^��ޡ��B��dC8�Ǫ��T���:�K�#�{z��x�z:X��c���b�l��ۥ<#��Dz��p�9HBϼ��y�Ϝ+]��c�ȣ�];����u|��`6r�-�����*G%FL���L:��]N��H��U	��z�X���ʗpy#֦E�����&5:P�>�k�~B ������Q�Ҧ��{�*���>�l����w�/�u�w���<W9��&U۰L���)NȚ�H�X�ze>�GE�V{Q�	`c���}"K��}y�Y�Cw�6�t�Jv�ڥ?e�x��zP�/�����	�M�M�e?�5�'c��E�G�U���ߎI	Qi���޹7Y���*V�M9����un�kn!�A�sM�v�X}:��u1�}1�|ث땒L�B�/o�a}P���W�,�(�*���;q�bO�9�	�}\���:���}�{ޏֹ��l	��,@�"o�)���c���f;}]�[Ԟ8[�O�����9�//����g�擔��SP�v�;�0�����BxKS�7��:/�\�����ǲ�f/��>���Ԯ+�}�ي�
���
�PpL�3S<��yHڷz�E�{���:&�d�3e���s�1�A~x�uN5M�ϓ�[G*-O���ʓ�z�%�QQ�z�zc�>/$�g����s�gKk\�f�@�yK��2߰1�Z�cz��}�@ol�s�;�g�ڢ�<W,�/{��}xz�X���ez���8���-�G.�!��ߠ(�0h�oޖ;��h��z���x�ჼ�� 3�I��6��"G��%9�z��=o:{}Y��b�x�b!��9�ʣ+�8�;����H#huul��������?W�d�(����͆����a	y�i�!�{���o�Ӻȑ���p�71��#W	�Y�����-�?� �����%x]�G���,!-?g;����\�?N(��tR�,�S�U�[�62�8��;f1c��W?�dُ��N�?o���;��|\i~�u�6�����Eo�+�
Ɉ��x��]#�(� ������i�YصU�����|��+w���
^~�"e��C����%�$��:1��LNn�;3]��Tz�ޝ9�@q+��j�"�k����0v��C]4#*I�>����u"�Y��W}Q��3����v�E��7*fܦ:��a�c>^�㠫�����n�R?�]�Rz���P_9�N���F9߇����pnK�sɹ���`�W���r��{�v��h}^˱�%&ቶ W@ۀ��a�#@뫆g~9���|^����t:I�:&{��"|�Z��x؜h�1u3���I=(��cЅܠh�]���z��B�K=ƛ���0|"3	
�=�ͫ���j~��T��k��٬�D�Tة�������y`����1s��g�mz�8��c0�:�/N�Q���O:�^[a}Ph��A�x����|Q��*؎���~��,��U�0�%3�,��~�� =	Ň��b�l���%8��5�A�G�$5[O������b����C���g���aN��`'��tfE��s�7�KOrf߻���(��E��ze�*+�ыyl���o�vW�7�{ڲ#�Y�Ҙ����i]B�gާ5-�>;K�D<�5K�ٯg]0WK��r����/�O�K�y��bF/S��q����f�ȏfgu��з�3q��H�Ժ��OEF��ڄ�һ�(�(:,\�**�`��˙��[��uT�)5��W.#}w�����������::mv��M�fa%5	����n�o��=��b�ޭҏ��8���su{��M�t�O�S��#������=�mgg�
��b���T�cb\ٜ��
��xSs�=Ӑ^v����G*1��VܯG�tE��A���4���B�&obyQ��z�*W�Ј�á�&��S�-O=>���@�~\(R��%R�%M�k��=�<�!�V�A����U_˒�ߟ�0f�5&m���q�]51��0A�81�O7:�����z���+�`X>��}=9W�E��ob1�=/G�0Né$H��"7�XҮb�8����f�9L�#��"�֣|_n�B�=Onb=�PPa��mJN|r�Ý�\n}��şe�8]d5.��&,uMܟ%]�>7ƈ��B�(��.�3y�Q�3r'�HHff�g�+�{b֫p/�쪔(�����֔E��=7m�6��BϚ����'�,V�����_�F���U����zܫQå�m��%��Խ#M⁬хv����=��"�Bz��b�OΊ������}��A�1�,8X��ײ����)�S�NR��txyXK�y�e�����x�.����Y��9�.��,E�҇ud�aҘ��ҳ����fl��{s�2^��pb��u䀇�B���*��\p�aqv��hn�v-��c�v�9���ԓ����'��ޔ��N������и��7����Ⱦ��{�daabV��΍��z���� ���Et��єb�	NV_\����#ɼD3y�~�;����\(��45̑Q�H�^p&g�~u�<�w�O�T&0k	��?�{k�z�����>^���SU�L��X��Vq}��=ZF�Ө{¶=��lI�鹗�y���H����0��t$]��O:���3�����K��O���_:AF�<�V��W�P�u���P���"�g���I��Z��G5^Ĩ�x���ⷿ������5�Ö�����d��u�-�vQ�є?~��տ� �/�B�����צS�6�j�}�����uu1�������z�*VY1�j��g�I���A����Y���c7Нu��L[�o��p�[��t[>����I�{MZ�uJ���h���{��c��c���r-	���>ϐ���ٌ�ŸZ���N�ja�]fj`���Ҽ��g#���:8�o�z³���O�$ ��E/JϬ#vܽ�U�Ƹ4����j{��]q��$J�f;��d<	�p3�5�F	ݺs�:="¸�L���|*EV/�J;(R���i:1�<�/]�gh���{�����oXי�.? 1���Ց����zv����ԉ�<&uk;F�Cs��a��&L3�6v��ސ옺�!�U�HIM���e>cCZ1��9Dٵ�A�J��_|&sӪ"F�fa�qD�7��M��	��)kޒGw�=$����W�J�j�t�38�����j_���x��Aϕ�:vD�S�=�N��M,��Yy睷��E��b�1����<S#������&4'J3j�ÁR'@]Bz�W�7&3L�o�����u��N; 9x�+�����`��'��5�2�F<��3�)�x#u6L���.�'8Rr��W@ۀ��%t���9��qF��o= �OҜ�9shъ��YZ��O}9�ch� �눷��`K�� D�hM|�7S.'�1ޟ}�7��;p�:9>��ERӺj%˲t�s�n?���]�f {��V��S�`���'������򿦵�v��
���ˊ&$:�W�\Tv܏���S=_Z���|T���n���\�1*�"�[�Ss��Л��%���3|��Q�d��,����S��8�Pb��f-���5��8W�Y��ey�uS���/0F3��>��[ӯ��O<��^��o�j�H��z��} ���m�k|]艷�s�d��Kȗ����u�c/���/�2}U��o";~]lC���F&��d  (
 ��@o#�]��s:nR�W=h�%�cPUnvf��0h���έ�b���9���.��\4��4se�iZ ���Le�/o��
�F��S�������wF�o,O�+D�H�#,3�ι�#����%���zq�S��W�Wl�b�v�c�x�w�^���"�.�=t�����d�ل����uk>t5K���C�Q���õj�m�ܺI�ܒ̄*�����h�,93nʻ���K{t�{�.H	�������* e	N�r=��t8�f\���ЙO;��sluH[�3$4�C�M�j0�nH���W��-������7�X���E���K:M�7F�ޙk�I���ŝ��4G=���Kf�
U��䛆�w3j�]�w�|��xs5�Vd����S�E��Bj��oK9�$�5��^"]E����-����q:e�s��t���3�����,�HHF��Pi�12�2�b�}3+V���gn""���/{+�V���R��ٗx,��B��Ѓ���U����"�6l\6�u�ۓs�R�0C��.�j�-��=H,[�8�<'�˗.���[���_aJ��5R�Y�e¨�W�5�� �̵|q+�j���v�mrS�NZ]���K6���GHw���rq�,v����ݬ�Z��0o"�l�+�t��.�g��J��jtt��033��u�ձ�^�;yv"l���b��V�H�:�Gj���%<ҵ��E�Cs�'uA���q,3���q
��5����<[�YS�-����Y��x����l!]�e,�8!����f�]�4֥�W;�Ϲ�X�Ř����X\�E��q�ߚ��V�g���6���z�<;%��B�λ�T�Ew܌ኵlE�DE@��$��+]�(���9敍��^�3�����R���fA�t���^X�;`:�:�Sf�&�6��X%w����8eөJ�������ʳg[�n�4�S�Į�3cֺ�ۉ�]�j���>�C�te`q�E��zhsigm�;��b���n��bdv��u��ڇe�]@T���Ll����S�M%zf���4�,�����ޣZz��N�*��C1^*w&fƩ�;�iK|�<��Qd5ׯpEm�+���b!�yx�����,�o�R��9�X��a���:ط�]�t� ;I+��W�Z�8I�ٖJ���w�����":���<�4�3ei������9��w(��9]�8�;�W@��w�_-�"��cEZ�|)��Ӊ��XuK���5�¥ݎ��U����Ix�Gy�h��ic2 ���:;����5�pr��;�2op^��W�ysfE�h�т�+E5�"邭�s���B��}����
X2�N}{1@V�v3eCv��5��=}�n9a���ۻ�`��N�EMb��f�;Qi3�\�%�z�f�|�H�r��y�^i-d�#��]�$�~���?o����:N��=n���(��6�瑭�"�Ⱥ�E���;��Z��sD����dQUR������K�+T�q�''#uʺ뙝 �z�uK�e�MVD��⹑��y���(�D-H��Μ��w!
�^�]�,�k������69���R��|#β��vG1�nP��w"�L(�ͤ�皎�h��Y�sΑ�8��n��]��=�*�B�M�T膈\�s=�r�=�(��$(���u=<ȝX�U�˔9��wYz!W*�ȼ��+��eT"�r�0��^E��I��M��|/�����wfV�xÕ�yJ/P�Q*�H��'Ĳø�O<��Ee$k\��Ku(̋�jA&ʽC̝��x3��]*s�����QU8����!��˲�' �'u*.R����{���Tv]weό���xqR�QSP�q��yw�����G�y���g*L�&��%Ҋ"yʞ�����W]��c�ʎ�D�E����ά�ȶK\Xv���^�����ȃ�཮�$	Y�9������nͨ���| ����b?���#�o��M�걢K��_�E;�צ�\X�ҭ�q2��*��ͤaK��ޗ�X��0#[�϶sf�����|á�p�\�lN|}�υy�K=~��Fk4]\ՖA��}W	ζ�!�x���Q��`3�.o'fh
�v
�S�R�>~��Tެ����2Ea3����2������ld<	��l�}s��M~� Ǚ6m��]~�o[ST}���1�C��]!������s"�����Uc�����0%^S�}_Og��_i�o�t x5�ᢾ�%C� �VŹ_y;���\s����%�'X� �E�FS����%O��ipg����z���~��>1�CZg�,Y(�/n����k�Ъ`{sMǦ�d�N�s~��{5���d���f*��L�����G��t�r���(���Xn�{�Wh�t�73k{����zL0ٵ�z9��R��"w>�A�<D�]�:�ytPg�<�Qt�Ea�Y���z�q�as֠,���t�����a�S�'�8*`Ϲ�V��x/���ݓq�?s����?���rT��]EsL��SΟ�.c�ӂ˷�K����YM�f|o����vxJ�:�
�/:��(+R��Z��T������Y&�a!Q�u�{�r�N������c.#4XFV��.���Z76fҺЦGA#ê	���$'��}��J�/\�;����+��R��܅���ӊ�7X�>rG�����U����������IOΤ�Lh��U�����������/q������]p�gȊ��4+n�J�y�Sp]:#ƈ!tfk��3\$TPCi������7�;+�W��"+9ZS�C^~�Eϩ�Ց���ͧP�ύ�\]'�{GP��~A�XF)r��'-�����M������q~ݔ�(]�#a�~�#>)_�p{�a�lK�3�hT=�-Ͼ�����7m�����^W�j���>{҇O�zPR��\,�3������=s�+�hDO�:cEZ�V�P;ca8�u�=�7eZ�`xڇ+Ԍ�b���-�ش����oч+j^mz'�X�����y;��棏j���|�S��'�=޹��A��M8nT�9d&�O������t��-�W���9��M�U=�}����O�~�HH��HCϴ�BcJ��'8~
h8O~lc����C�Fe�Ϗ�����^���M@�<�躔�����T.�s��[s�=��m�?x�ik�5�H�'ݙ���:	v%�C�U�(,hւ��9N�ͱ��n �Oq�g����9F@ �cc(�)!b�����M���kW���8�P��Q=kQZHσe5��f�|��u�!������ze�P�)2�͓�r�Sn���|�65{е�6~�w��ং���Ŏ�����F$́"}@ftT����V��{#���J�M�3�9�E+�S0=��M��f�N�&��53pUz|$NGX�.�T/iLǅ�foٕ���)�Q��)�{��t�Г�>�l»w�;�+����h- �����N�^���>7��޳��*�6��a�`<�k�.�H:!�}:��cm�R1�c�)nb	���?y�;E� u�'�
} �y�\���@1�M�[�3y�~N�3�<�Q��;�Ҟ�<�i�������ع�:_p�&{d���n^�q������V�muu��%i��ǲ��,������F~v�g��Y_���}�y���P5?,"������D�E��}��^���|���"iu���"�h�E����MB��!��"�����gKX��aQ��=pMwvK0����ʑ����b�0���1��F�\�59R�Ʋ'�T;���i�gb���pא!�H`�9�/�lƭ�q����3(�P~�Z�dNq�@ڛ�Pe���3c�^#��@��S���m�J:�U=�O9�WDԨ&x�׺v���N���`���3T���Y�ؚUuj�)|tޫH���\�ʩ����l.�9ph;�����#�z���uҭ���d�\�#�%�����̫d��Ě���qAq*$��)C�.�,z�[�F�W�pc��rtn%bԱl��"�)�~3��J�����ALw����zsf��v&)�����z.�c�� �юX�B��-zG?t�'��0����s�{m���pnׯ}8Ozh��L؀�;R؟e��E,iY񓬬�����a��h��2�ϔMAR��xX�d��"7*���VDz�S�̛�!g`�B�V���53ئl/V)p�j[�d<�T
�J���BD�S�=͘&J�r5==^4�e�e�{-��23���\���B�mT����4����gW;�	#���2A!���z,R��ݗ�^���
3�vГ�s��W��8��SG����-߯�Qw��?h|hC����N����(�z7���&��w��)۔�|.`mB�Y��3̦����� K����A�4�6*c���^�����d3Iㅽ�|_�2k&�M��+"�t���Ӆݘ]��V��V�!P�)����)���.L y�I}K�}���p87�%7�������R�[	�^��1�w����������P�7.b�K�V�Qn^���he�ѥ�}VŰ��ږ��	�/���*h�ҳ��M�h�Kj_7�ˬzC-�����vmM	K�׽�8��G��QG�`[й���|>�s�Ԟ������[s�D:�МE��Y������GܚU�|�Cy���
��m��'ݯ2X��9k�,�{� �s��bs��Pa�uS�g�������\I�B�3���z�GH$�b��ga���jtY����q��IǑ�/[������Z�{׮]GJ�;3q�J��u$���Zg�(S���>���2e�d����F2�Dv��!��~���/9�����?u�w{����ߜ�6ig��L��64CS�z�a�����՟qb�l��>2e8�O�F�@�^���]Vd�V�=9��y4e��隗C��p���Ϗ����)�"�a�w� Ҙ<��c�g�U�s�6�!�x����GgцvੈU����+��(���g9����y{�qT^@[�A�z\��-ʙ�-ld<Mc����c'յ/��`{�ޫ�uv���g��p��b��BWLB��0���Ȱ8���ʫ��61g��0��v{���"Nܼ����1'5}:��F��},Q�ϻ,�8��1N���b�ˎr\��sa)�!���G"�-��?>9{.�0��juߣ93�S�t^c���m%v]�#&'�NW����@b��(e�x��~�4��L1�,<�meV�=#��w(�	�٧�o����nW�|���c{a\��Eh�3����ax`�|����燻�����Fd$!�����bM��@v :1u(@�Ɇg�� ����?x�P����ZK��ido����eK��σ�L�73tL
	]���ý�R��|�;�z��0o1!�=>����*��~�cXj��Ə5kf]~�?�T��k��٬�������G���ЅxZ�{�i�������1�pj�.��B���ҍ����b��?X8=ȃZ�_t{�~X����w�j�6�����C��}8-T��b��� �^G����Xg<�c�=.0: H^�'3a�|f	�!}��&(`U�5+�C�0��`Z���<e}ޗ�k�񃖑����4"���z�C��h=2����{ a�~3�������釭{>�f_��O��(ͩ�[/ǣ��N	�1b�����6t�,�-?�6
I�0y�?����Ō՟l�멺�n�4y~VϹO]]������-�!����x��GP�K�3�h4=c�u�;�{59�o���{�z�ڣ'��\Ū�C	�>����R$��%|����W��ڕ�B!}�~b�4�=�?U����2��y)ڟ��Oطz��6z�puH"7���qpsݴ�z�R��͵o�"�#y�b|�VjY��2N�L��;n�h��6?�R���;s�k*I�c��*��n$���l��Q�p�H=wC-��(B��+��W�2[���$k>��� �Z�j��/,���O߹NF~�2�Lc���^�f�g�V9z�`ǯ1@���~���mK��{�-���{�ܸ٘7^^Q��G�B�_#.�*�~5�<4�WꔥO��T�U�i���R0pN��_n�dH>�~����Gz��z�b��}V�E�R��c����i��"����N<p��p��{��Ke�1�Lez��lw���`{F�LG�j���躔�tS�yP�y����>��fS����"��W��7���4_���u�ʣf��>�Hfo� �ώV9[X3on�1[�T�<�9R�1�z�?[3q�j�joS��WSzg�t�	p}G���a���(_i1���y;sjKy��R�Iـ��0�F<���Z!��(Ri���%�^���{!Lc'!E�
��`�a�\:~�C�~��%;-�R03��<g6dCW�O_����8��	�Rc>�>R���}��(0&�-�o=/�'s۟j��0*��Tl�Z��r���p�zFzz0D��\�
D��j�d������A���>��7�~�U�誐��	�=���>��]Gdn�VU=�G��n��� ;9顮���[_����~�<���L�;l@�e����7*��W���:����m�7�2�[ȥV	�"�幢�:�+4-��F9i^a�t�7��+�B���(�)�.W��� ���֑�q]�Ó����®�,.����S�¡w��^S1N}{+a�=��@�;��W~�1��]?	��		ϓ��[F�-p����f�`�
E[�G�C�u�sj�_�(��׽.��a�����bj0/SS�sK>�^�q��jY�����w�(�G<����@c�u�����3lƽ��.=]�+��x��b���q�@v�mC�ty<����A|y�J}Y@�Q�<.�_޺f1�oE���4L[�Н�5�����=��gz~�9e��6�쁈����χ�6j/읉�a����Z�R>ϐ��F8Ib�*�����%^�`Ж�p�6��g�6�8���w���Ozi�l�f���R؟d]�A�`0�̏p�h�/����*&��c�ϻ�<A�5�+��*��9d�3%�c��z7�\��_�ky���Bފ��S'�n\:n|r��T�TdȎ��D�_��^��ݽ��{�S��u��,,8X��1o�9�������&�	����\�����
B��́���z&l9Fd�xq�����nڃp5��R�{8��U���d��X��#S��&�=�?^�~9a�'���#y�z�Y��Y,��z�ż�s8���`�ZB�SR�e7-�ܗ�s��#�w]84d�)/,r8Mrǥq%���/���8[�^A�&!�������(��'�{���W[F���O��?Y2�݄�i�ՉX����!���ܿN���a<�G?�A~��\;�����o=f�M{&gފ(�;/��T��&v������� J��� țQSb�:\_���N�7����O������}�=���Мy>ү���Wf@�ۄ�������'��-������5��Ut/_���~5�@�3��m��`k���Ы�Bs⢁��>�²a�S
����ĨU���ޚ�����x������n��W�X!_�=��.���-������UeI���5��1f��Y<�bLT>�X˭��E�ޝ^G(�O<���p��R$��e��f�if,�I�\�G��?�<��+4Q�����ܕח����F2�Dr�b�;���ޚ"�h�
��^@�`�c��T����|��r�K2���,_24㟴�u��������³�0��>�.�pf5�hC�n��xo�3�k}8�����X��?1�#�dP~��y��/�2�W�4�D.�,Aa8[�9z;.�<t3|K�͸w#EZ�u<{��;Y۷h�	�����������`��G#�B�E@R�A���B��8졡5U����I4�i���v����iͼ�j!�k��닞� ��:�n}�ik�N�װ"��߇����ՠ�A�*j�W��<X�tU�F;��vf��C�LzC�*I��wˎQf�#��t�,~�X>�g$չn|���ߙ����8��;f2}[R�šsZ`���==�����2b6q>��<]s��ndq�m�
��D�`9�:���&��v���秩��z~�?�V����	q��dA�<oъw��ō��u�K���Y���^�Z��'7X��������
F���`.��Ŋ����f|z���7�v�:�/+j4���]�#�m�
N|�8�� ګ���ע`Pc�|lL�C����e�b�5�EDvp�emZ�,,
��F�Jӓ�Z��Y�0?T��k��٬����A�I}�4s0ܧx��z�����c�P�c�\:p	�]ӥ�;E��
;��
�6@���󀪠RU��mw��$5�r:�s��&{<^
8���UpN,>nmG$z\7Cۉ�c3"�ɼyj�`H~��8V�������z��c��pI����x
�SU�( �4``��wj�t�Yw�I��q5��*IN�r7�:d�L�;�s���.
ʽ�����j�F%�����U�5��5i�Qt�*�&���`���K�N4ȡ�N�Yb'A�5��z�#��λ�׮��),[��qd�n�V2�fɦ�!��s�r>�u��1@���̥��}�[�Bn��L�9���)��vnâ$7NL�꿬�r�j)���s]Q�J�&٬�#�*;��E�s�}.�;�z��x�/��f��/�����L'�7�� ��|t�G�hcx�*�Q�X�R��8,�ҧ�dg�7��n�|���\��)n�9Q�WC˕wN�d�Ҙ�S�-<������$�Ap���8A|v��ˆ�ӹhK���|���W�;�v}��WRZyZ��V���p���`8���r��]ٓ�n<Idj������P$LY�k7�c���#����QF�^���30{��YU7���
��w�;gxt�"J`4e�NW�ں߶�<C!�.0b��
c��V�\�F�u��"���"k��aGYB��,����;�x�8���CeZ�:��$J2�m�O)�>��;p�c���BL�t�Gm�[�ϭ�9L�!dj�k�U=�e	�kRx�uh��H�c|G+���^jZ��1�C���bi��c��ڰ�v�W9�,|�x�o�Kޮ���N_�b3��cv�b`�g5+]k9\Oh��sִSy0��;$�d^Cg���u�$y*Π���YvM!���VJ��gs=ßmEtí���+b��,α��-�85�H��p�VF�}5V	��j���]�\x��:��ΰ܋�M��7��5yKkt��wRj���uB���R&�L�ɴE[6�b�W,]ZΤ,Pk.��h�j��y��Cm��p�td}���<�M}�8��WQWm-u�l�K{�����:Vy�Ó�{�+A�`�Z�e�A��t�w���Ɏ�-��z��b��V��#�u��bn�d���\r�tg���E��o8��������r���F�l)�St١�ޣ���?�F����90ޔ�wW,w�G����{		S���<X;Jax\�R�t�}��EDup�S�5n����{L� A���;�$l�DŶ��MZm�q/f����]��{iam�1c�Up����e�7���3�Yw؎�I���JWr�[f��.g%��'��le��@WF��Z��P?<�\��U|4�2�]:�m���G�j�WUAƳ���m�-��6��w0���;[Vn�G!]�Li�Ǡ������)@�s;n�wB:�vɝ�h���Դ9w�C�P��7"����[�uM�̉���yt��m4aR�UŘ[�ĳ��*���r�]��a�Vb��ܛ\�Q6��IWrXr.���en�D�:�nW�RW�e����"����l#���++l΃��k�oS;RuǸ�և�k0i�P�j�f8ZYb}����(�p�����'n��YU�U}���_PO�|yU2�7�9�J�ˮ���W�ۼn���:�8�y�P��;Hp�Qf|ql�ۛ��q��B4K����DPUùb*�{��֑w	>yw�w(��r�0�j-�]j�g�Zj)MqO+T��T�;���ΔGΚ�����rp�s�R�hQEI!WL�������n�LJM�R�+�K��VEE�EjGQy����FaGN�<;J	��xt��Z���
�ue��!Fft�R�[���R9jQf|8�.�,�O'��dN9%���0�M#�����9�Uz��{���n	o��� �^�<��X�d�W��l�*�{�;#��Jl�Й�+5e�y�<�*���5J�bw	=R��j�i����מdL�hJA\�8�;�;B/qM]>0��̱�ÄV��
�Qκ������f����_�8��.ςGqܾCk*�x�9��)�����T�ȩBڬ�*�C�6��/7I�vb�qҗܪ�!�ͅEo<��m͓M#2e�\3G=˲�J$�bSN�:�.�Pռ+pU����{,팫KB����֊	��뉕�.�ۄB���s^��Ċ�6�^^[r�f�e_{VDTܱ]����ݻ�ӹ��X�uy+��3�s�B��u�ѮLVM/u����%��]Z�_�Oϲ�䶅���=kT[1�a��L���8-�،M_�pu�?Hȟ��ɚ_���{�-�����+�£��{��	�Ł�՞��L9���Ü�]�����Gg�뜩^B"}[��3V�,��t��D�c�EZ��"��c>�}
'����b��Yr������[{�݋�͌��z#��W��T���k�c�t�#r.���T����2�!U[��&�kQ�"���ĭ��� nO6+�]���,�u\�� X�
�]KbGT��i��"����	ǎ��`�s�q�g�({1��j�e�V���>٨�P��EԠ���)��B��O���6�1��v��n��?P��ٜ��a)j&@�y����'��2�U�~�,�Rs���xnB����5���g�b��g����`ն�����X�󚙈��|���U��T�{�͛��{1���������Vܘ���_���$ ^G@�ڗc9F,�~��w�z���K����n�2u��՜�Zw6q8u�kνj9�W+g4\�������N:��e.u1-w�]p�M|4j(�3=�P���HAW\fJ���Xwۦ;�������G��*���ŕ�R��F��
�]#Rv�c��6��@�;�z0�Ș�~�r������.�'��m��Ŋ
�<̓yX�e��3O�~N����IH��x��ˁ7[BhQ�w�C���?N��d�@B~��c�Ĉ��}s�Z�c����o=.M��{�OG��=�����~����u�jx?	V=�Fg>!P���8��v�߅������3�1&Ǻ"�����Q.;/���.�3��ب��B��ŕ�������f)Ϡ*S��Uu���:�z�s��I1�!k�ޝbk�D��1�h�E���~�%��2*�����E�_���-?1��d1E{�^W�v4�#=�ؚ���8��1���FϮ\x�i���U5��sC;�)I3_������T/����{5M\�Y"���]�!u1��b���}8�3�f�No��.4��zl��*^Ț���
�Ѿ��G�:(�Cz/���|i�q��;�O�; c�d*��fzX�m1ޖ/`�ߺ}�Q�'bb�U�aȴ'¤6<}�!|���8a���B�	���B���{?ѱ�sz]�C�y&�1�<�𢔥7n�)��j��|S��5�G)�@�Fp�om~�!Qw��."(Q��x��7[��F��
<�U4Uv�r��r<�[u�/̬�n(#{�434�<m9h�gb�{}��TԶ��t�[K�`iK#�d�H��G�xg��Z���@q�;O�/�^�F�M9����Ď��Kb|*Bo�9��w����}S��Ha�0U�r���R�d2�����$�Ĉ�{x���(�;���vt����vS��X��j�3`��ˁ�����d<��ʃ�*Y*"t���}�;]�xz������,J��XP�.�Z<�̌�����r`��Bf�I�� 2����ޞ�;3�1�%�1P��~x K���t�r�e���]�w���s�k�e_\�z��Qi��/��;~���x���8�}|����Lv��b�b��H��k��gl=���@��=�.��zn��-�
�9���b�_�?]Bw��>�<9��(����^���������$�w[�����s�~���~*��IUF���V��V�!P�)����y׫/��W��G3�n�̩r��xL�i���?R���e}�u��(|pu���8�vQ$V�e��Om��^G�@cD�dX�w�v���ׂX!X�g�;��'������j���	�~ۜk�oe���.S�崺� S�n�#:9śj�qٲ��������*B�M˥l&��"���y��L��J��V����(ͭ�E�7:(sv�A�oy-y�,�
G��eO�j��z��I���@h^�9k��3u��`У��|�&�i��gl.:�V�Tu/�Y�u��u���[�n_���Zg[6:��Ȋ��P'����ak9*�V��]м�n����P�-35B���`��OR�]}FH>��g6�#��}fnat��.���U�0R�	�u��٧��L��D
u6�����7|MŜ!D��e���f�Tq�<�?1}�ձ3�n�˳[t��9�Jv=3�t=~p�n�)cپ�/R"����<U�'��A��
@^C�ߛW��<X�v���3�;N���d�B�Fc޼N8����?U��8"�@'�A>�g$չn|U�lиe5�64Q�1^�WN�þ��Y0��.F$��T��������n#�vY�T�|5[�m�rUV9O�lbv
A��Y�y��;��A5�(J��j*�/(V����J㳆Ys�������z��4:X��$���{�F�*3�1A)|�X8��
�Q��pY��P�@t����=�ܯ�%��o0�5ߎ^��w�ϣ�;jo�
��eǦA��b��D��:���I3u0��O�녟���l5� I��Y%f���+r�=09��q'J�r�bk�S�/�����>�N�I��o�L��U��]�NΛ�/�"���*d)�b#zԹmN)�̔��-�b�k;�~b*���^fl����ΙWY�H���M'�l�s�^��Y���mɍ�V�oq��*�=��fb:��B`Sr�ϻq���s�ןC��LzY�eC�Ϗ,�ӀOЫ��J5���U�0)���0Odj���/D:	u�$p!����0S���Q�9�S��Q��܅�CW���X}�7X�;��!����I����O�8���<	�_�ա��?���
�~Og�/)�'�<k6,���^������K����ܲ#|W���<b�i��h�U�r�Y�A�^&��j�:vc�o/gSs�w��"�6��u��4j�l�k�3{4�u����[����jn�n8�S�����g�秎䞍.eVt`�Č^�!��lF|��D�����Y_��I1c�`����P�9-�����\��n������H��F4Þ�]L9ϵиY�g=���x{+jV�H�Ӧ!GLV��Z&�<Yy��4*�U�G�Eչ�����Y��M1ӠX��|�c��>�N#�:c �ۈO�n� ����c�[R�mz&��]S�q�t��z������N�3N\O;z/n�?@�a�4�\�q�nγ�Y�߲��4��v��d|m��guE[����ۭU�����ݨN�t�S	��D�-=ձ�Ji�+!bF�a��״���۵���<U�Ż7��7�5�-��F��T�kh�@��.� �����Bκۛ0�P.��"�d�iW�?�~���A�0�~��lo�~}}	��Үc��w��xlD��(]��ՙ�1��Pރ61�&V���>٨��(0�z/��9a:ux�8�hxf���F��>�P��	��' ���5�C2��/�3;^�1&`FG�uU]�L>�i��c�/fm\NQdE���+�=��⁘�l�Ƭ���v�c]�C�j�+(�{�W�ŦI��Ϣ��U��2�,�P�zFpI⁚͘W�tS�'�M?y��ׯѩ���7�����%��< ��\(�(*p�̓yX�e��a�}:�%;��/Xy'f?3;��ɐǎ�P���A�D�:�]	���`�@1�݅H�c���J�̫����/��b�����F���:"U��\�|B�<�)7���G���\Ç�����UGoa�Z��[����|U�N��,.ϫ�b��L~b@4<�zN��TdF(�,�1�jQϧ O��"�'"z���T܄!�Ѻ�¶�����(��U�Q��d_�*"E_m[��b��r׋�h��t6ꅈ��(����t�	�v�L7p�L�zJ��>=[y�D���(ffvP�Dg|:�y�آng^{k�;;�t������^��w�6/�Y5���������179\�Ǘ����z�OL�T���\�$?@�@��^������=\�fs��Q��Ü�?Xc>ig�{^�q�n��6�b5�O�HI�v���YC�t
�%H�{׊z�0��.=˰�uu1��/w�����X�����#�l|�P_�e�>5������>���0�t7^���X���P��y~�-�k(*��c�����*���ߺsӛ5�N��0�bÑj�zD]����*�6驉!���؋����(��`�����󚾗��Pc��n�]{�Ξ�Ӝ�g�4 �!�l
����5{�ݫק�~{��er���/��g�	�n_���j_��Yk�Xdd��9��r����	7��כY�焸�UY� �HG����Ԩ�����B�P��уPR���{i�T��qɁ��:.����{/+s"�^xnsUk��	��L�_^z"�'/�fW���m��@��| J��"z�e◫/�`�]�w�+�Uΐ��!;0/��[�U������?P�8�dMzA�X�k�/����s�j2 ���66�d�J�q��Ӗ�Qe=8�k��2(�GF�#���F�;P�y9ț����k Cn'�]g,v��J�����	�pExЊ�kB����ۏr��m�*_Ƚ��=�n���O��eN����Y�v�����_!7�m�\ث��r��$׸�U�w��]��N��ܬrc^�'hs�O�
��'���(����K��ׂ�W�?{��r�(�S�ՐX���tW����]�8׶�>�;O��<<�^��&�\M=|�������K3��K���cA���*�В�A�V}ap��tT��J�U�Ǣ���ν���x��闢r}�Y�4�T�N�[&���s�RTHA�r�Ց�5�[��!��%�����ʝ�U��"�\[�S���|�y�V׶��,���LE��fQZ���F,Y�p�K �<�v�u�3
v`�??�Tɖ��J�NT;$Ö��j̍�q�׵�zʨ���qٴ!��~��^�8��Ϣ�i��ɚ𑱢��_�En�u��ˈ	�GΕ!(s���Ϭ����U�3[�s��@���:8���D����Պ&��7��y���gJ�!��.l4%��Ey��M0�e�!��m^C׋n����1�.}�k�RX��[�O^{�'�?L��hu��3�t`,��,!`�ќ�M[��ʪܶh\3�kl|2ӝ�{�w�]���7��dW��>I9ח�[���X
dԪ� A���LΧ�T�B�Ҿ�pn����KE��"î�A�d�W�z�9�H��P\�(P;��Uc��Q��
�gwLw���e[F45)�b�ۤ�E���:�������k�5�wÌA�Ő���/~���6,Rw��hB��������nے���w��_b��ڻ���B��1��W�ǧ��}�O�(S��";�oY�S��c�˖"�]F�3�j���f�f�K~sa)梁,�@�hI�+���L do]\3%��ꤽ�3�^yJ�O?��?�/n������U%:&qϦGy4�sc��;�ܱ2?+>�ǔ���tq�*:o6�Z����b��F��m�1�j���������G�gG�1u@��VW�/2@�{皻H$9��/ ꨃ+%��3��^˷ �*�~��;E/���)aSڳ�^�I�s����3΢��G��r_yet>��OX�����_�q{�j$j���}�F�QCxo��C�Q p1#��OVW�7�	��}�{���r�yg,�&�*��Q��
3K�+5��z�XU_p�_][oh�b}�N������u������\�z߄�E!'�XD�}���}q�M���s�M
���~C?�	�k�T�Qp��wms�k����ǽ���p���ؖM3����0��s]����u{'�=R!���0A�Y��z@(�_K[�^���u�� ��#��d{���z�o$�8�_m��&VΗ�m��[$q"��ȹʧ��ʯ^v���l"�ö���G�����n:M�5��Q��so<����<5W�^�3W�ϧ��|���;Xg�#�Sp�������!x�>=�+�8��{b*����W��,=ϊ��/W�y�g8cY�u���f�ٽDPf��4Kc����rm��������z/W	Cs<�}�R��>�v}��z�٠�u��|�^�W�/$;��;7�䂪4g�V���2�f)�ǐ��b7%_Kzg3'��z"�$G�{o���*:�]�o5����w���7�c��������-?�44Cs����~/��CV����l����ōV �6��ۨq��Tex�w�����I���m}z/��
�J>���^k%V}o����NDLM!:\'�=:)����k�k���G�+f[�`���� ,�@<��[�~����;;73�j1�[S-���吘x2�s]#3�C����7�4��oU%��2X�����s��#���'��wf�oX�_RnS2�IGMeC���W���Q���w���c���s8Y��Y:��u�Ȟ���M>�YԦ�My��}կ���G-NU��q�M5��[i�Ӹ�EJ��ݧ�D�)E��O
*V:���͝�/S�.�u�*$y��c���"�}DzY6�¤/�����ܵ�d�6�X!Wi�/���*��Z�n�	u����t��Q���x�k3K��e����b��&b�=����9*fR[α}}�]:U�V�i�<DN�ٝ�P¸�̴�F5��y��s�vo���&�p��**����3 �K�)c:.vgG:n�;�)��1)�Q}`MF��Xw��@�o$#v�E�L��WݶF!1��W+���z;�eե��d���a�*��`�\�t*��֓�w1>M�X�	�mk�-{�.=t^�d�r���eu;)������d��d՚��%%����қb98Eݑ��m�����q�T����]�X�؀�)�(���^nP9��u�/m���:ܽ�{4��*b����52�L]Q�`��ٰ��;��}�.�NQT�o^�pi�P�ί���cz�V�гvr�*�@]&(��׷�
S)�q�[�k�Ԅ�ˊ�����w�0Y�T�z���w����o���wl���QU�}o��|����1�E�A�~���� ��Y���-���Ն��M�ëE�lޔ��6��I�h�#z+��xůk�[r�N�Ӄ�.|�1�����vr��z5�C�S�c1;%m��b�f�".���l��m�^X��#��U��VH�VIuz���y�%�;\���;\8�չ��#�ِ7]6�����4��b��3h'�7���P�ͩnp��,!޺�x@u&3�e��0�g�����1s��G�ۛ&J�.���b�E���,J:�K+�c���7�Zׂ�5��'���K_*�f��.Ki�v���e�S3����K6�C"f�|�l�C�������p�!��L�pus�˖�fe��!dl��x*`�k(l}�eE�!Nd���ݞ�]�Ż ��o�˖t18"Z�m�4�z1�n����͸��su�k�ҳ��U���o
�{MQc��x��P�B�VS;���<N*v�?��������֧u&Oq׻��r[�J�x�޹]�J`�;A�Ơ<!�[`���`�E�	XwxD[Wu�������Fgl1M�g$���+ʫ���G)�Y�����vn�B)���k;FNUQ�T�,n��x�c:�u;��9Sa�ݖ��<�ݬ�4��5�jw���iΣ�e�>�h�
��+[)e(rv!yҷ.��}Ws$u1����y��Z��_'���nC�����YtR�W#�l�S�"<*s�r�<�ֲ�� �����,�����.BS��u�J��	"�h�G��yǌ��<�.�ҵ=�W���ԧwu6��.u�\9gĴ$1I�O'J�%TM/=�Meh�p��8��%�%��9n�:���%�)�����g#�J9^u���	�^��g�#ś��;s�G$x��ʊ��GDΒ���	��S��"T��
9��t���=�Ȝ�\�E
���&_h���DJ$^wv�*�o�Ȏ� �ľ�w*����B�$����p���EL�u��VVBM�K����.x��s\:��B'�ǞG!f��;;]���I$���� �=J(����UR���;�z!UQD��x�'3�r�h$�TL�D3P�y��7B�D�9�+��I
��t�r���-*9$�y�RqN�NG��Uw$��
�&����\J��燘;��3��&���{aZċ��*Xs�\�%��I�@,�
"��ݷ��=㻮N�� ����q��c��o
�t��<Sw.�]&I��*�)�Ch��K��"2�����ٳZ����s�W���8
���(��kk���H��FB[��w�l�r�m�v�#���+o�q狾Z!W�T���j���*2��z�C�gz0�7�LE�_o��5ieR�Pt����-�}P�^���\�Nyei�"/��'/=Ȓ��O�$���њ��Y+�S"���s�Ǽ�y����lN{�m^��G��<��ej�p�GOݳ6��Z�t�T��Ӆmd���4'CB~�z׾~�������j�GK�}����p:�z��Uܿj'����o%�\0��U�l���o+�zbxJ쾼�wn2UƤ�����sO3\�����=��y*�bX[@?Zؚ��:p�;X��e(�)h1�+��F%��"�;O0Of���y�4�X�`��;}��9G�yE o��g'`�m�����`S�8n7%���c<�7��=�~�ԌDP��X&�\� ��>�&�by3�2�.51U�Q�i��[ G���GέE�����Ir��X�=$���1͉>K%q��,���5��t��Y�AE�΁,�j�]Ndp���a����Ɵ��	'O �Z0mIi�Ap�O�v�OAx��6��/_g��vgDڴ���e�߫�+���?`�������/���Ë��<p>�[q��ݘ�U�ݪ��ݚC	�]H�GP���>�$q�:�<�ޥ�K��
�d\�ʙ]�`���� ������+ z�
��	��_<�וޑO]���OZ�5����'N�H����Ͼ���Yc��c�`�$A�U�Y�f��h�Ѿ�8m7��5o�Jh��׼]l��eu��S�]v��g�7��H1��M-Y�z;���JD#H���ቪ���gc�&����D>��WQ>�:�Z����#}��شዌ�[���̈�ޏ5>�=_nܭ����M�THa���k{G{�����%Ҙ��u,��\��7�珟�)L^�ﺲU��ރvn�vׅZ��}`ĳvgߢ�?��6��CRţkq~�1V�N\9��TPl�P�-c����IDmZMZ�;�Joh�4�w���v�ItLgKƱ^`v��Kޱ����I���u���j"�z��[o/�������3�2#;^�>�l�yi��q�Q<���X�E�����1��Ը{0/ �V�Mlp�c�����4-�DǦ���=gb�v9��T�v�qFv|���S�V�_kG7�m��y���{�O�>��G���M�\����%�xU���-�b���zv�.TO�ӗ�'�����a\}��ΐ��6s��ϾB�4��ShĤB珳ԭ���xJ�̙��5ݷ{�?�nJ���Cr[u������q����A�����$�̟n]���伇�=�0�(>����Z�_WF��uX��h�z�,��%��I�1���u`#�,��}(r��q��ؾ~�yL��,�v�_z��}��g���O�bd�g�mT��8�
yױ�^;��H�R1x�#P�߇�5��I��_d�����L�B0s��:C5!�;�JL�y�[�����)g����+1yn-)-XO@�#&Y��f���L��u����D�u%L�Wτ0�V��͝�d��6m���g��C��@��YL9:� v��X#�À������o�.��fwwS�p��䳐��Su�v8	q}:����>���p�ǁ�1��!{惉a���X+���S���#m�#���Pb�߼������)m_y;Y�c�}4W�i�����.ox����ϝe�R����G��q��2�-Y*��D���ᦾ���o��u�c�|�$���C�׽�M�H'�y>��Z�[*�\hS�7^�4ly�����SmA������ߙ�Y">>m��y�a�b�L�o��^˝��4�F�o��z����ӻm��9�վ,��v�c��3踆��^��j]��_m��O��/D���+���V�yM!�}��ø��0G���AZy�3��y.�b@��Hh����;_ȓ�b0����Oh^�WsVY:�Ja5���'���e�>��=��p2�T+���������(�-o�4�A�i�s�8lF����c�wt,�GY��x���&��c0��h��sU���m�w{�\��F��W�)�MXb[�z^&�U5)M��8byոƮ�UC�ݓY���<�<1�<�I0ɜ;�U�8���������-��˷��zw���TC
�:�S��\-��G"��E|������	�����P;m�}�Ze��1�r� �]nqZ|�L�޼��䤂A_h{�,'f�%YG�[�^f�5I�~G����iR��sϵ��쀅�}�XSEg޻/�,�}����U�%��3���W�^��ZQ��Ɯ����?q�ڞG���}-��2����jg����Wg{��[b�L�>*�1�$y����)���+G�vM��Q���I�7��+lq���V� �$�o��*ǘ�s�_��/������U�M����hYPvʩ>��-�c� �So1Ͻ7�W�}����K^
��[� ���	��$��ذѕ�o'���#��G��gU� ���p�uR�M�}�A�o��6��`�z�(������1�hv�8{���Y&���45CC~�z׾�����|���PˣO31U�wz3�y�/��]A��Mߧ�-ɲ�^(��w"�V�&G>R�lڽ��9Bv�x����`Q;g	[��Ǖ
�.Z�'���[�U6�u��RM�Q��i��v*t�\�7���͒�in�=�2��VqP�����e�!'�j}*�/[�wP����H ��cb�m�\���Ic�%��%l�#�<��y퉻���9�8���bY�7Ķ��g�gqvo��U���������m�^n�W��=��.V�$\Ѳy�?#Aa��`5mhI5���{6�{e�l>��L��^½�{{��0'X"P;�!C8�&�z��{j�E<��лL����q���3�1'���3A��4M��z)�'�u�˶�����k?���q���q>X��P����97���#���e��k58�Z��_j.�P(��F�r��ܞ����T�j�.��M@}BH��I�|oR��y<���k��=���W{������}k�Ư?�l	�.�U!�=�7T�����6�l�^�9)k�Y}������[��r�/�11ӏ��;����R<���;�	M�׹�~u�=�U���N�6݅�����F�%��<2ua��ؒ�Y�t�酩Ul�Ƽ���RZ�Z��Cҟ^C�Kr��T�ÒTޡ��u|���R
���a�mܺ�{�щ������o���fCy]9*m���Mergi���@j��G-\�D����g�h��̒��FD�Кz�W�������������4.*ԸUm�����$a4���1���yP�z��|������>-��"c�]b����=���d,�oMw�;Y/���5h��~�f��o��yęi���לSfz���J�.-�~b�S�{�VJ���F�L7 h{��� �����l�fJ�kϕz�I�`>a^-o^��c���]����j#yv�a��m�y<P4�1���W����S�5k�������dY�q�3���<T��4C�ǁ��$N����O>*��ռvVGި0o�^r�[�����ǒ�ٱ"�m:clE4�B��GSk@3I,���똓��������>a�Y�p؍�V9PCr[�C��Н�����}f��ܽ���d]�v���ZM��d��G�=��l ۸'�65�XѺ��oW�y�լp���ly�E��$Mh+o7�^�'�M���ej���x;)V��N}|;XpݻӇLtgr�+���'W����fZџ<H���Me)c� �LO�ܳn��-����V���Äh�㠶�qI;/�j7�fB���%����X�{�y�}n��`��<�f��f_UC1#t����g�\��]����ҽ|����X�,�OP'�}I��y��#�?X�����.	g���C��fO�r�q�ϥ/fro�Y9T���74��%k�Wy��{�G���Ծ��T�j̓��,x��\������H�S�pD�W���jb�J�`}b��JB�/WC�T��揢�,��ʐ��P������������[����D�'��^��͉ս�fikGb76f: �_$f�7��П�)���J��W,��n����u�;o�UbX�;p%��]����#��<��Vɱ�	�O�ns����>��`��C�]}�Y�5�*���]]~M���!�b�;�����:==(�U��D�x����H���t
�W���^sx+�|Xzu�'kx���8�_�����}�*ݝ�W�\����܆T�(�ni3�L�r��Ѯ��S��n����Lȵ.$4��P|�4�k{��25Tٱu>uw�c�)Zȝ"�m5�}4�h����[��*��C;���"h��v:�UmC��-�V��O���{P��z�������B��E-$g���� ��=�R&�gh��В/3����e�>�Y���At��Sb�`���b�\/}tq��b�A8���)��&��VVd��}�Ͻ�z�����ڻ��b�Q���b��.��<���J�֒0�l6�&Q�gѹ+��������S�s}�7�S���z]����w���>f;�]gϘ��u"�j�o�2r"��05��M���^��-�/3X���&#�-��ĺ6�.">�Kɀ�����@=_Iea�-VZ�ҏ�	e���AG�)���r����eV�rǟ� Oz�Ƅ0[\�gǖ7�-��_�{�����w����N=�����X!�(�8Б��������@��j��W���}�����ܢ�����W��X>c̡��U�ٍ���ѻ�w߁��1Ë��`�%�6KH��GrX�u�D�knh�c�u�8螘G;�h�K� ��h�E����!�]�,��3E#+y�k:�<�:'I���z{pX��^�#a�Ȟ�b[Dj�ݻ9��Z3����L��' �=�h���'�Aؚ���(e��èi�aAV����S:��V�	��u0���vl��{aX���.�4��v����k��'�C�m�a�${�s��]���b�����R�
"�}����� e�^{��^��y���+XSIZ�HP�D�`��Z[�<� ��?��@x%C��^�=�ֲ�����S�ޚ�ɚ��G�E�g3�2���mcg���k��������&�}h���8/
��%tQ���2B��y���gH�u�����ؐ�Ӧr"K�T]�_��I}c��hX��/��Aa� �5�"�i���lw�Z1S�]�F �4�`�c�rH��B��!C8���m�i�u��p0ϣ�6n�����pg�)Gd���"�BKg �z)�؜gRO�ƚ���s��*�9�DI{���*�6C�� d�ǪH}�Z�ֳS���,�����1�G�y�>0+��kܪՃ��L}T�
��w�a����f��SB���mVӒ�*.�:��GP(�4�35'r�ӷYʾA�<ڷH:�Ë�*
v�P��S�2��tx���м��_w����<B(��z��/�ա����s�-&�ӝ9Gy�b��1�s��.����nPX�%�0���K �5�m�Ջ�{�w����Y�UC����#���kn��ZJ����M�o6�gf#xк0�x���ݝt r,��P!Q׻`%�QJ�J�F���%V���9�Ԡwr�ѽ��� �z����C�E������&�N��+��M��r�Y�V�T�4Q�0�U�$Ѿ9�6{u�&�]���c�n-�e�VQ����[#7��q�8��퍬P1B�o^�6�r���j�T�Tz�;/.�b�骈]8�����<�\���Iv�>��Dv��y!�|���J3�;�{f�e]�2�WT�՚,SS�I�Ch��;����,@sKcS�ȕ��+&^�1צ���!Yt��}���%q��f.� 2Ő�0Xk���l�w��P������&+�v�;e�S��>A��g�\��d�-��,��
;�ZF�� n����4�)��61���hf`��`�qއE,�ཛྷ�Z��z�tO�����v�,�sk�x�u��7R۬B��@�e�ȓ�K/�f;�RZ�Q1��[W��0p�;���N:���^��u����#�f��ܺ�i�\;ا��3jK�i;��#upj٣W�Vg��6��Rz/:�ĥ�8Ј��X5n;^��k
[l̔�s˨+��{�;��1��Vst�7�b�an��v�6�8B���"���p��(L�9���]�w
�zQ�a�:�t2v�T�E��B��P�-�����4�86�]��X�n�j�ǌr'���lJ��]L-v�e����ԉ������F�ܽ�N!�\_ΜGZ���^�n�j�h��Vs"e}Zz�����֞g��0iHp�Ҏd�(�-�V�,v��P��[�5Q�����c��c/$���Y��
�I�/�;��V�<���b�ik��OG;[��o/�9aP�++�$��:n��aR������d��T��5M�;�d'5���Me`��	[�e��*�)���ox�/p����lhǞ��qL����z�*����1��ؗ�-&�]t�=2p�J2�aq�.�kLo>a�Z�F�#�T�e)�R�b��盓�����LMW�[�T��xgE���d��(�bl�;:�/D��V�/L����<T�
��y(pج�/N�1^m���@�9��Mj���.�@�e�kCݼ���U�����n)�*̘\ᔘ�3��[/5����ź�*�U개B�d��|�o`�낓�P��"�ٗb,FP�gLz�gs���8ܽ=�����L��n��Ϻ�}sn�A+�.=k'j�Pe��S���3S��F���M3L���
6.�ŏVES߾��9'Ȱ��4Ћ$��L������+�r#�a�^�� �*�;��P䗩�>0��$�u�P�8� S��L!2
����VsZu=��� ������8�� �*��.E(=1�T<�!�wH
�HO�P�Y�>A>!(���2��B�u۝e�u�8AW�IΝ7q�� ���*+�2�l�D89���D:҉�O�<�cnL��uV�Y�Ww0��˒�ӑD�u9TRy�\�.�A�ʼ�*�$+�\�B�iUu`�u��H���Y\筋�9иmN����
�G*.U�PN��n�EWx���_r�<o�
VUSy^%B�aJ��!wE�Ey�**):r&y�9	�dʢ�O8��;�ʊ�"��s<�9U�'��!8�ȫ�a|c��T��I!�L�
-����r�.U"��V��f�J��Q۫�C�L�$�uu�.�\s�dNeG<� �?���ڡeh���Q����FA�W:��Fb����TJ�{R//��£��e���p�R�O{�uI�C��C�9���(���	��?v>x���	/����)�i2��W!tv�M@}BH��I�^�t`���zO����ݖ�䖛�ف6��g��e��Z���z
����X�y^��q�#�n���Ib�%-x/����o�e�_c�d����ۜ��ٯ^j�=�"�}R>)߬w���)���� ����Tl.��u��/���r�Ww%������~T>��Y^��=�zZ8!C>*�z��u�}s�o��������3����P<�^.������ym©��a{2r�n����:���u���ӠvVI��*�ƪ��kz(�bQ��͛��>�|{޳w�& Փ�{9�?1��1Y�vVJ�����0ې�u�uz'��}��������[�^��Ŷ=���b��������O���o;\nr�w�d�!���ޱ�-�~�W_�üjҮ����{��$PUu��u�Vo��è-�5BH�}A�^y�2ڮ;m/Mw���c_��nt��i��V;��"��q9�Jq���e��ovgM�v�9��>��S�v4�j�ݦ�
!���m
c{N��Xm+�bȲs&�PZ�d]����)�)�99V���z<;�M{[`�!�N���)nHm_����>���T��F��Q��z�s�w��{n�G�4����lGSkޅ5�;K;����{�J��y'�4�8n7%�ܤ
m}-����'^T}]���i�4:�ў���h3h��<���>V#ޞ�Xcs�LO]���]�Z�I�� ��ֶ����W��Q����^2��$ߙ����Xȓ"�s{wu�W ��ktuv"mN�ݲk(��+��5x�*L�Ϥ���o>�zgݴ.t��I ��������xmb�Kك�}�k'+ ���.�UT��z2#�]:)��W��;�@����y[�I����>ʐ|�r����o55;��﫬��pA�~�k>��X+���Sܻ��	��0Ϯ׫�Ƕ�H�\�p��n���k���/���4�:�뿋'�f�f�2���x\�����Y��p豙y*���L����&M��X�a�x
��9�/�iۙ@ً� ��(UpC��|����Qx;6*����i��i�[�����t��v�n��Z(����jt�A�zᲓ��+�D�;���0�v��>�T5����q��䌮��J��-�M��'-��
�vNV���_z���
[شw?{P�rH'�y5����W8S}�n􎑗E�2Gu��
X9��oVG��ɰ�y�m��ؼ�olUh��VK=+w�p�p��e��C�	�ޯ{��?ŝ�?�/!ŵp �[Vz�z��}������Q�=���U`y�������7U�n1"n.���Au��x�ϕ��o��vlM\����׮M��������2��BǮM��i�Mc�����;�.ϽB�uJ�;�����gs�=A��8����ii���6�2�	8lT�J��o��c��~k����`�6�U��A�.�}����9�+A�|�w��{�.}�C7�[�\���Bz���@�T�^������k�J;��ɺݺ���{�n8�h}xL�W���w�C��d��X�]Wozl��*�.\�{1���ojs�+$R�m�8v�;1�25�����*��;{W��R4ւ�]�Y�y\�=6k�VH�ˤ�;Lݬ�YB5�T��J�`���b)z�N��I�w����K�b�b�wC� ˟�����
�}(�	����1|�m"o���.]_w�k����kpu��=����Bj�r=Go�`-j�n����Pd�||r/aD�߭�l�*�-?Gq�쌪�Of�{�Ժ��S�y/&py6����t
����D*
�������L�C��P�Ǡ�ah�SOVW���;�iҸ�Bʃ�
����Vf����\�����h!(/��TOT���ij��4I���M�`6%�8�&���<;~�n��ڕ�1_VI���G��5h��o~��aߏ3`w6%�ɍV�0L��ʓ�!u�������c�Y.�7����{�W�7�qw��s�r��T�}���>a��i�����{y+�00��Rs���(-x����1?M`�Q�,u0�96�[����.�m\�6< v|" ؘ����s���'+��ǈ�׫�*j¼�����N@��ޗ�]�&u�	���올��3fU�9�f�P�ĕH�0�ꢻ �:=�q$�ҼHE+gǕ��c�1-�Ӭ�y�rS��K���5����ܦ��AI�l�i�ӆ*��E$0�̂�p�e �o��׆o�۝�Q���f!������7a}A�BCފA�{8�&�z���":��Mux�ˍ���R�1ݵm�9����@��i�h.^�w��gZNB��b�[z�}��̟n86l�����q�$0ǨI�u��.���N����PʎvJ(���7	�_Y�a9	O̩7�W"�]������8���]^���Q�ez����v`I�����}k��Z���z�Wv��]�E��ׯ�ｉ%���)[8(�y)k�Y}�4���R���$�����~�7�_J���ߨl!�u	�����V�M���{C��`*���M;�3CH�#<\�>��!W��~AĎP��Y^���(���Ͼ�m��V��U�4�fmoҶ网Z�u;<1X8!��XJ���SOVWj�����ʭ��e�n��n���ڼ|9'�����7��{Շ%7Uz^i�}��C��jIɿ7��,��e�̞��ԭ�V`;LlϯGM����:�
QVH+�s�7��m+�e���Li�:�oh�Z�@O<������O�Z�׹���'$�l֧\�x�Im��﹚l��<�MwՒo�)��_]-me
ڇi���Жd�wd�g�W��M���-`	����1���Y*�\N�Sw�����f�5�Fw�#N�u�vpW�slx��~ŭ�k�~�v6�\�/����ϻٞ�V*�.�G����=^�1K���!Ň�g�ZU��k#ꭀy��Z�"�Bg�9��y� !�_h���E������&U7O!�1W�$�*J�_Z�m�������oU���6�SO�!_"��+��;��DqWsV}=؂�)s�Bi�'�ܗc�7�:��!Ȉ��z��f�uB��k��	ZoL�+GM���#�q�OX���v�TC�H�胕�5���Q�V�h��*�o��^�$����?^J��繷r�~�mZa=�y�L�H(h�T�_U��W}W��bd��X�&�]/
����۷�쭜���Ah��}uz{5�'Uj0�v����3������ Ɣ�~�S�׻���s�xh5�h��m��7��g�"̹�yԵ{�.P��O$�!b�w���fuf�B���4,U���|�0e<�ދ���s�9_D��^NW������}���Ԣ����6�B[~��>r��0���:ږ�o�IT�~�`�P���c�Ƥ6��g�;�8���������Dg�}��]��_%�3�d�]���;��>�jO���}_�M�S9��GV{t�QKD.��'�������@�OÁ��{\B��ӕ ��_�/���������}�O)#�y Q��֜�^��j�# z��>�w�R>4Hvǆ�]_�<���J�r��j�!ɠ�N���U?��z��w�3;z�D.�^�X#�lG޻#]	�j��f��m��y�a�bV��9Z�G�]Gn�_g�_9�4n4;�������][~-�^ֈ��=sÖ�+��"�s�t�,$}ܚ�l��蕛TE���߸��C����'�����JB�>%+�i����.�Y����F�!���Uy&�7�A��e��k��T�b�����a��%7��|�:�X�D�6��7[Q���&e㳨z��JTi �o���B���C�Lc����si��h���q��ђm��Ra�o���s�}�c\�sf7Vɺ�iwo�Z�+:�=w�4�`�鑸��%��H��dg�KO\smj�o>M;TV`��1�d�|}��a���R#���G��p�S�; �Ɛ��-����ep�Z�a�w}e�������c�A��׆��-�@�T��N+��v�ߺ[NG��u��7d_^QmG 4�\LA�l�ɦ���s᥼^f��!��kB�G޼�G���ܞ����]��'��� ?T�ヮ�U�'[����>��J�W}]�_y"��d����nq�;�%�L�=�����Wz����ܮ�i������?aD��m+gWO��Cx*�W�.*�����r��*L-���דiC7�9V��]-Y����-��Yo����uu)(&��駽��	_�=Y̬ZA¦z�Sű��Q��f��5�w�)�����������kA �����I	� �N�_���^�����p��o�{�Y]C�.����5���C���d�1N�'֫����v(=~��^�W����!e�e{��g��0�k���.�1*�'mc�i�R��+���ka�#���E趞Y�w.j���tX�,��(m]5���x��wCqs��[���7���cL ��cU	�o+��tg�w�ߥZ�`׬י3���(.+Z��jw�����	���ַ0���G��ٻ޽�zQ72z�5�ķ�0�=�m�E���DǴ��Nh�a�O����O˷<��N�χ>+z�x��k��Y�}��r���<���Md�_)��h+Η���>C5p�|�	��i�O/��-_�m\��Wb�[�}��Tw❏�7뒇�E7cB��_��o@SMO����pI8�����Ax��I�q�*�HC/�->��C��t18��[��ي�L�ۏr4��d��gz ڰ����(�2G�1?A�=|��D�y�r��\P�{f�w�ι��V'Gx���A�����t:_�?�!�>A���w!�72
_z�
�����,Ռ^rWw|��Ͻd/�O�W�'�J�����k�v���b<���S�(��P*�g�ҋ��\#��7��]�EF��;�ٓjq2�)cf��9*8]�\g�|3ʎ��l ��,�wa_���jM��=��[t�{���ny�mm���{�#�Q���F�;�)�0Κ�Qtw]����v�e���d
��P��W]u��6��^��	����]J�V���J.�6�IS7G�>�? �}#�_�c�c�q���,������DE��b���;���Eo`���8�a��N���Q�����v���KJE��^�'���z�To�j�����	���M=Y]��������lZ���'J��Z���%��H4��g���;Y&�Q!��0�������0f�ѫ���g?gOb����!6<JX�����{�{K:�=C�04���V6`��Z6~��G@�vϧ}ɱgXV��&�=�Ǭ)���{%�������S�nQC�X�=+K^��n�=︰��ütdDf�MH�����*���n�=�ko'�&$0��
/��;�u����K�.pMYb�$I����6��f�.;{.�lH����zC� P�
pl\��g�i��'ӣp[����4��*��+y�&�,�ҏK=%���#ٽ4���d�)�R�9�x"۬��O�KCp�����0^�-�zFV��j��1�.j��P��V[t�a�u�felsc�B�q�#1v�����������1�=w�Iy-�ڻ�X��%�Ug
/Ƽ��ݶ�J�[�#�WQ7�]�vl��/�ӭ�Nf9B짵H�Qb�n�/���klϥ�-��A�*������{t�3��ٓ��o���!5�G�7(��,$y�_h�5I|��7�.��<�n�$dX,�Ѿ�s;�통I���2����g![j�]���
,c��Қ�`BH#�.L��Q��_u6�܉+[nޚug�V�%9��2���,wp �qIw����ȬrH_u��Ewe�R�
�+���)1�l����u[�7�g4�0�*چ�\w%S.i�����}�����i��Rj���=\�T�_t�Ppy���YB�2��o0a����9�K���<�o��$Ӿ����Eg)������H�nL��(�ut�,l�;i俬u���ۮS�Rqj"�ռ��������_+.bĊ'��kM�b#5�Ң�tn���lm��i���P�Uϖ�c���m�eE�I*3w:!ء��U��PA2�W�%?'���xqi�7[=1uwVԴ&HHv�!�����X�$c�Az3�"{"y�x���0ml�*匍�H��Tv����kcLv']E͡�'����Z�7L��i֩���,;5ZХU���	@�-��L	��Y�!\3p�xil$���p-�*�#�+z+0p���jr*�5��c.�#)���9�1�v��s��
գJv����w_�C���1�j����-���B�&�:�t낵�uG8�ώ��"8����<⾻Z�Ӥ�Id�ƹ1�\6��L	�Uh�ÍGTU'H]s�F����8�;��N��;�E+Yr�q��xi����jVjxGUv��G�����Y�EX��fv������La�dY櫴���T�����B�� }S���mw ^�A���U�|h�9l핶89�r���'j��LB��F����m��6�P�����������2\�7)VZ��6�Hl�Iڧnf����*�;%����:�X�Uہ�1���a�x�*�Q̪�)��;3�(:]����^ޱR�s%���>ɒt\+X����ս�<��:p����GP�ˡ�-��M}Wp�T���e"�}�kU�D�ޮ�M�K��B��TPr�$i�e*VVno_׽*�.G�E�e)<�oy�n����2�l
���Ҙ�X����ݤ�jN�a���[zl��,y�����p�̘��qu�v��	w#*n
`�п�a|����n��(^r��"K��$�����C���K����v���<�.�c���5P�L�	�>�j���Na9oD�%�u8��J�Nr~��
�.UU�J'�N�r�l�\�"��Dz.�{tU9��*�09ז9\�s���G�J9�! �EqD1Ux�#�A��D�3�ӆ���eQsAW'"�J�.˹$�B/$�蓞�UR�LJ��(�.r"
����ʲL2�.�8yĶZ�<⑒ZI��95ZT�eT��aT��f	�(�3�	g�2��!*.\�ԋ�܇8�j𧩙�F�\�r�jpN�����B)x�F��\�i��I2����*�^q�**�Fa|��]܎9�1ͼO;ǲ9T\*̎B�{�Tr�HPp�Ufd
�.r����$�:IP�g��U�$�S#�Y,((�!�]�\UP����WyO<��.]w,�)����g�����d��P�j٥Đ�%��dQp�x�D$��H/u�+Ը{�Sl���)t�ma���t�oݜ���sΧ�%�wU�ss0�k����*��%#waku mL�Ǔ��S�ur�=r��Y�k���d�;r���A�-�5s����Z���^^��U&��COZ�i���+:mX	s8����x٢(;}S���o<�(8���7��������/n;�����t���Tmǩ_�ў|��� t����w�]�k(�K� �걅�Y�dQ빝�����<�_�0,
�U�u ��Y]U���&%�g��镛7�=7��F�ws�)����>��q��ߍ�w���F�{6W����};}��Z��̤M���pA���}�>i�;7���d�5��=ew��$Oк�N���k�pC�Q#��*]��uj�{G��a��M-�(�Y ��_r�,q�VQ�\1X9	�zm]��U�l����]���ַ�{ڄ�rHXM
��\+��/2cI5;X��DP�ƛ�{�+ Q��f�C��(�]��j�uiKFkmĝ9��Ю��J[jB���e���M�,�p�*�v�҃u�'�,��Q���3�{�F�+� *���u�B�+S2J4h�.�4�_q�Q���̻�JKY�G2��!�	r~���p���1E��U�;˼��?/0��Led����X��HNz��!��_g��s�f������/��沺��"Eגc��)܎Ԩ���؀\B������v�U�@`1,=�+��B�܉3�7���� �rIp�{�����|��`]�5s��$0���6jiU������>��'��;WX͵�)��L�+2w���nE+OF���M{�#��@�^��$��D,!��m=���2�2D�5�7NUz�sw�0g�)�K���&w�zU����7��(�Q�M���ꃦ1u��1��������? ��I��ڰ��-�`!(_VL׵VO.fb�������W}�uO����	��:�8��9�d蹽��w$��m��d�ϭ�Z��;@�@�9Pv���^��;]�i;�{q���[�1C1���=�%�O�VD�:�,ЧBY���]�=oFy��]�פ�P;m�ƛl	�YB�J�����8���р�ר�SO�V�w(���fA��%��u�z��X�8Z숫�ܽ�:�c�\:��,��C޲"#><p=��F|V��m`����>~ϊ'�J�gW�^��؊����q�=hHN�c�����b��U�ƺ�>Z�z}B����?j��.f�P�4U��
�'��M�_�$9���Bʃ�Tz�T}=���I���a�K</ly����W��,���kI��Srf"1���tg�Uk�;��u���F|�tT�0Ư�^7�]��S���jo��}avn��u��>��ԸM�J��,"\X�c3s��'������8�w��t�������r+���˓}��v�U�Ϣ���o%uFwW/�9�tfS½vx�#��;��&��C���x>�s�Ǯϯ�sY2��,]t��<=�E{���ú$p;_?Z�E6,a����|餋e�"��M����O������G{�z��;�U��H�D|�d����1@iN�F�u}s&6�zk�{zz/�q�>�k�#��C�w�u�*�D<��A��ꊬ=I5�6I�nMi`�0R�u����1WmSiK�|1��`����/F���	�5ۭt!�4)W4أ(;�%n�đ}� �+p�wP�&�Y���/�5*K�bP4z���ߪ�]{�����������/��->��C��w���O]g�ҍ(uR����מ��=��~�	�B�� d��?9��^�y�
1Ugo޲E��v�=�x���|�sM'�y����큥�ڏDE߰tz�Nw�c��dNE��U.�׬��]��MU��+�ֽ8��}h���i/�m���M�c��{�����ri�I8�ro���YX-�"dx�Wg�g.�ׇ���!����0P*��o�8�~�}��9��]��@M�v�!#�~vz���B;��W�ڬW����(����u��^u1�}���;X
��J���Q�:a�s��i��*�S�~2}�?v��娥oރO���ش��g���;�$ߢ�X�gX�q��Y��N���C���Bߎ���w��ĥ���)��c�Ւ���
���i���~�f]u����p�vbQT���+��UM�Y��H��=ȍAڢ��J�@G��2��8-ʹ�����RK(�ٸ(U��q�0�(��$G���<�w��љ�;Ӫ��߭�\"=�^�n�8:�C��R���W[0�Դ�cd���eN��I�L�xCY�߀��g��ɱgXV����B
�usgr�>�;�\�0=����{����{�X~-���Z{���Z�������m��<����E��~�,.��7��zDfN('����Û�<��mѯټ�]�{�
\��Zx�3�N�L��r;���xS���Cҍ�I#�N�E\u��.�M4e��.��������(��@��fƗM���.�S��`cϛ:p|�=�xaA��˞���\ x4`u,'c��i��Ǿ�m�v�Nz���L�QT}�U�K����==X�⎠�>��(#r��lέ�K�:���-�P]EN_H����z��٥��D��7�\~ʾ��iZ�K�h�=7� ����iA\Wgy#�U�ӧ�=��hC�Hq����C�0��9���"WĚ$n^�NĦ�ʯ�n��M������Q)��i-�~>�\��@`�bK���=��4�_h�A溪	�lX.�Y��]n�k,���q����1x1��7���{���e�̝=�_�sw����yG��I�v�ݒ}}�j�F���?g�����:����� ��-�N�KV�n���~�b�����9�����J��vtF��s�O��0;����=�h��%a���h$զ�Qc�����s�1�X;����=B�$T�^Of��w/{P�@䐴�Ƨ��7*�ԁ0w��M��Ӓ_Pc	�֦�����m��7��J���.}�!u����/�$g�h�<9�7��ip���]�P��J���ڳPLA� ��ؼ����|�谎�����1ۃE(u%y��aыgw';��Q8h���)�y���5-6�_<��}`ɼ��ٚ��r��J���wj��_�{l9�{H��W\rm(��M;
�̝��j���?k*��͍�?Ym#�K����HoR�HC
��M- �i�n1ܽޟ����j�v�����*9�z�O��˾���D�]���z�wp�f�����B��(�g2(_}��2��N��t�6�b�6�s�A���5x�����q�I���A�<e���Rd�e��;�C!U2s�P�&�j�f��,ISwt0Ѫ]_2_Hd�?h��2�2]�O'�-���zU��S�m��y�^�c�^��ǽ�F�O����w�n���~�!���{�^����/.�ag��1F����y�V1cX&�v>uO�� t�~���p�0��s,�l�f��6�;l�g-Gل��Y*��ps��	�@C����W	���w�n�|A�b�������Ϟ�D��m&lp��"oNl���>���*�a;��~������am�i+ �mg���U�ƺd�r��9�6�� ����� �Dz>��M{L���W�̬Z7��u���Vf�>�;�Z����͎{.�5.�]�+��]%<ˇ���09���win������3K�+`i�*�ƪx����_���ȿxƚ��cl��$lw&&�֬�A��c�Y=1``'f;�O�
���` ̸R��Mgw�?��K��H�S%�s�vސ~2�)����疓肶�Y�ܺ�N�ĺ�ۺ��~���p�iz*��߅=Sz�k2��f�%�p�kY�jk�T^]��Yv��{:�3���c�[Q��E6c�( ���jߪ�v֮M�y������c��J�B��f�W�Յ�<�1'��{e��7��U�����ϵ�n�f�z�_�x{ŉ�9�d�1ޜ�6�]�ؐ��k�Sb�����Κ���X���1ѷ��<�V��]��o�ȟ�떇���a
�)��Q[�'}h����.��v�����ՔS�gѹ.�D�2���d>*{h1���>G܂�����@v��	���^4����-\!��/��[�,C�ޒs��}�(�^��y��|58�����sКVʒ�J��C�s�c�~B�mv>��������>�Wm��zNى2�|����=Z\/�a߱[����nl�'�Ǉ/����u��v�I՟ro���ة�ݮ��nc����3�:��r�w�P*����mJ|H��ѧ�vciLgH���9���Nnۥ3�k���	�P��B�cU�Ù�ڋ�}gj�5�S����Vbt��e���n��U�rn���ognT�J� [��vt+�f6��e9W��i�a�Wor���h�oD�wfɆ���\�r�|i�M�z����'�]���\b~�bBP��u�~���譈����ޏ�q��~���C6����a�Y�̍v��`�pX�jg�{�,�x�G���M���?|�;����,'�g����c�$�ިŤ�0=�����֩/I:E/�7nZo��z��w��ĥ���iNz�z!њ����o�z;�~���O�aȩ�jh������ذu�a-l,��2�5���8��	u�v�d 7ج�0=��%C��bwͯ���Xz�ą��7���W��yQ�=�>G}m��<�������n�*����������<�b�����m[�f�.ͱ�e�Ɗ
C�1L�dE�+0A����>�&��Li�(�G6�J($��M<�9@�K�P�ED[��/8��Ǟ�=�;�S�P����j���M��2�M�	s8�� PJ̈]v������n8�7X.�ĳ���`��V7��;�N�V�����8|��]�g;����p�<�&�t����5{��7\�oT���E�9�ثy�s���w�mu�����*�s�(`x����2�<O>yD'Z��)�~�ٗ���-�x���;���!_�\�{���4���m�����v�o�0�G끝Q�v� ����t�Ph@�­��{�Qs��.������4+t������_����v��3���;cX�|�	euW?X���)@�����-]�k�������~��p,h����Bk(q���:�@^{��w�Sr�QC{���\��(��H��9����5V�]�}�G^�^��B_>�)C� �u�4r[z���+}��8!��E��U^fz}P�w���I��ԛ�H:��Oty{�&L�V������b�hge�/T�@��4��f��w*��69$7�Ѫ�Ů���[�	!'���ޚ��p�w�D�Tƪ{��g����� ����أl���Ww��$+	j	�^���S�l%Bs/��������>�� � �cm> 6��������m���q۵�c�s�x<�` �w p!�l ���q�l � A�`�<�`ݓ@�l,m� ��m�	�6� ��d m�A��d'�m�q��cm�q��l����&�m��q��m��!�ڃ���l�  ����;l��  ��d 	��A��  L �m��� �  �m�6� �  ��d�l�m�@ :�;m�A��d ��A��8 �l�m�v&2m��`�!�����6�ö���t�[�w�~���6�e�m�2�� ���|�z��_G�����/���������������������LG��߬տ��_/>��}�6��o���?M����������m�����m�c���{A�'���۱���cm����ǯ���{��1�����������xb���>�����l��l )����b�����`pcm�� � pg y��6߇����7��`�(
��
�����~���}�^�oݏ6�3����#�=~�`�����c�����o���~��~?���/�oc�� �cm��v��o�����o�6��}�cm�l}�������X6���V?P����6�#	�>��k��=��:�ŇӋ�}�����!�<��ǀ�g�#�i�������cm�}��7�Q����g��>����>~�����}XM��Ϗ��m����>b~Ƕ��o�Ǟ��}�<�����y����u��}����y�1��|�xM�����cm��G�-�~�X��z�q��O����Ϥ޾�X�����,v>���0lm��/������ql}&���
�2�Ȑ<t�t������9�>�>o�($�lɦ� �hh�E �M5H�
4Q@� ICCA� 
e�h���
h �Jh)A�[F�G��U��f�J��M-63[5l�S6��mZ�U��6m���E����Z��Mf--�Zklb5j�Sj�aP��Y�kK&M�h���;-���͖�`f�Z���m����l�mm���XI��mi�ɖ�LMj�m��&Q�[m$�ZB�T�%iR�e��؛hղ�R��1�m[F��  ���v�鹺Z*�v��֙�w[h�3r�5��]g[��C���g� :v\��:�v]-�(r:\����Ns��a�ӠOu��Zj���˹�2���Yk|   ;uǶ26�!BE����ZW��l4m����x�3�6hdd]������}��T�Гw>�K:4.��:]�w`[�Sw'ctۉv���ֵ�um�[�5�ٶ�ƺk�iZ��L�e��f�P6�iK|   �x[i��^��{
�la����+��T�5�]p���]��u�R�:�Zsv��:S�l�.��ݪe�Ӧݷ@]��Ҭ�u��T�V�4�Ed�ʫH�K6[j�   l�Ψ�r��ãFu,t���w]�-��)�Y]�;�롻-vnU:ܧwM9bws���ηsJ�f���8
[n���΁�:u��`�٤ƴ�6�S4��   9ު�q�]f�-Ʒj��t����tW9��X���S���5�
`�uۮ�K�Z]j��ۭ�`4�t����6KkE�4
�[x   m׀E֎Ӷ��@+�]�
.T�U*�ӳ����jwWuA��F�֮���Ѷ�H�7V�
wi٭CM�L�l��[e�iJ�f�m��  {�ӥK���i�V��]��A����(�h:ζ����q޵Uv=jܭ;�������n�т���"�t��J�ۧ�M�f�J+��[Pb�-l�4��  '_}}��V7�{�
����U$�;�m�wJ�EB�z���ġ���
����^��u��]�F�AA=1���^z�Il��y*�G��+ʡ����uVcSm��  ��(J�K�R-�������g��^Ĥ�j<��= ��L�{�R�Mj�íݴ@����J�t�;���':���w{SVf�Cj�l���f�J�   Nw���s�x��i��� 
{�\�TP���ٹ�P �of�(t������x�IR%�.�B)R��n��)�{�C��B|��*��  "�Ѧ)IR�h0�Oi�ԥSS@ ��%%R4#MhE?&�mU*   e*
�4  f������D�c����t���}�]"��1.^]F���A��!�b�}_W�U}_}�o�/��66m��6���i��cm��c`���1��d�cm��?|����@ջ�5�`��7N�2�[0�,%Gl��Ke���@[�wW	a"�[�W�@��X�Si�B�	[w���*ʍ,ie��� 7+�k-���y�٩���e�	�-v��R����r��u�5��K��"ˏ�rbV%4m�u1[�r�$�P������O��
��B��X��г@J��==j�=���[O��٭nI�-$T+3i�-�3R�{%#��Yt)�ʻ��a���,=T���i��`&��)Wk�8�JZI|I#C8��ƛ�b%젥�RJ��Mn�cm�G\�_)a�Nˣ�Z���m�[ugo,�y�9�A#�����ʱ@j�ds֚n�������ګ:H��8l+u�k��|���ZPz���U�)�W	Rx5��ڱ�Clɴک�Ywj�t�
���ww�uc B�XeM�mXx!j�i���5�O��@;�E۳���Z��У��n�����nQ����c�9H�U�JD5�R�M���^�Êm�8<��K7�L[�Sj����*�a�]67r��1;���-V�E���VK��:�m�m����2�$�&�t s`2��V�I�R�)n���3)%��:OȘ��V�YM^c1æ@���3+t�l#G!bN"�d���4�FR��fb����\[[��1l��z�n,j�͙fۘ���O���Rӧ2�mJ�aT�m��-� 4k�zUZڳ3n-B�(]e�`�])]���zI)��3y��?�$q���:���_���@�TÔe`�3��Z��*ne��i-y�nZ5a�
9M�'iՖ��i�ݼu�1cZ�i��VH��vkE:&��5P�Oj{l1�´d���6f��DRI������ �k�oV`��aq�N��l��9���x�!,K�(�ݘ���u�R:,���iݫ�{���u$���K�0,�'���-�Xn��R#U��EkCV7x&�j�YA���CuSwDfc[Y�!43�CU���3t����Y�4+��4�����A2���D�\�	�
Weʙ�˹H�5eA��B, c�0:�M��u�ըn���6��-X�ύ�Ͳ6�`�F��%u�,�,.�Xn���5����v�w2�`��m2�Z\��`Ks[G�S)m\�5��=[�r�����sN��xqEw��MФ#W����uMyru��&��T�f��&�: 6/��/i	��Fl���%H�Xd�V��Tl�Jқ��Hd�z�7�ײ����u���F�B���hlEi�%`�Aa"k1�ޖ��ΏR+�Yc����kKѐܢ��Й�fa��- ۴��&�륊�CF�tN�@0b���1a�[ɣ4��j(��6��H<��DP�Vlt�T�1Q5)]�M��i�he��q�N�^쳙f]�@��B�j�%Pc�4�����|��w2_m�z�5�Š�m#u���LSʱ�0�%VP��8jb�fPEI��Փw%��4K����Geŋ-�5��m!��,��jmf�Q�aa��.�C0z�w��GN=F����n�uEk����zKO���m �Ͱ�MF���ي*�*�2�*ݵL�6¤H6�ahM�X�6J����3KGp$���;�`����/ia���� �΃L3G/�'�u�� ���yN�J���\� un��5��BK���T-+3V�PV��2��Z����=�qt���N�i�l���4��x4��)���ᬼ�x�^�9`\��rE`Ү�$���Z/u���U��|���zMl�^K#4Q���y���^9n̄7kF$^���5upk.�#�iH$�;�S��Հ�0�RG�0���̠�f<Uֺ4���W��߮��(:+3.#��[�Fv�%����;��͊�����KeIzz��%5�n�ە�8���ګ,=�Ʊ�9���ԡSX�L�r
V�ճ�:���Ӎ�tz"���e<�k���z�H��n��6Y�7�)��ҥ;�Q�b��f,3&h)����S����u0��SŐ�h
��Y�G*`;��������ڵ�AV�d���n1E�$r��u�/盈V�����4�7F�^jt�B�c�E�5���ͼ�72�DS�FY4�Ԟ]c	��VuVI�Uʗ�T����ւ �R�2��Y``��2j�r�:݁�F4��{z���/�,�i������#u���"�D�`����$�p��J�]���.�m֜�!ݻ�K��@6�i�C$��Vfmj]n���]�u���jV�*iBl�F��M��P���=Me<�� ��+7b����Kok6�k�+�n鱥Vgrd"P).ݔ�{�xZ���pՊ��]̪Ժ��H�Ӷ0�Vaw�6��*�t�j���I!��
��_�-G����E�֙�B�S$Wins?߮ݔ�mdVZ;M:�c��T푟bʵmnh�J�SC��Kٸ!�$�;�uC�o�6�S�k��8�XP����6j-ma���������u�y7�iƶ���`��d�)��7���uYV�����XD,f8�B���[�m형*'���ն�6O-Y
.��j���M˰�<G�u�F�K����YC�uY7e#G(nYD]�n��q��[u�7���k�r�F��������:��x�%��CZ;�%6�7x)��kOvfjxR[N���Ef�d�]��imlĆmd$%83�su�{gp�%��w[{,ܖ`�K(C�����]<�X�֜�%ͧPS�;yf:�ww"�`۠�էK�3a[Jؠ�������e�0�-�+%ޱc ˏs.'1`�B�5�`tS��~��V��`�5��Y�ڂ�(�BK��v0��܄m�MғI\�,Sˡ�*�^����0���f �*�ү��X2�Z��ZT��umV�֪E���-[hY�a�u��re���lOQ��r����<��5��}m#��qO����W���)��T�I���9(M�dt�[�T�]�R���&���<;�룷T!,�hm����
-�5j�GH��P�2��s7Y��"J�8[����_m�:�.�F��&*��i\[u>K+@XH�g�70��i|�����
�QT��f��n<X��u��!v��/�d�4�5�\U�4��V�_#�o��4��J����ݭN�i��6J}��/R��"��x	.J܃&�=��}�[Z(ְ��L�2��ť�)�(�{�,�w&����H��dPYZV�n�5��oCU4�;�{���X��>{��߱
K�by3��WE#D�v��cj|���T���u��d���W[s�tK?,�t�J`�j�/ͬ�5����J��%25��}��ҭ��,�����(����2�v6�0���Of��mU�]� N������Wؘ�۠��O��;�(�g+D�+� �Z��0ȵJ��6��Ņ:W,�����Q���:�n��-��S���a�`���@�V��3v�6�^�F�l���Ö� p��kt�T7H!����g%�j��S�aRU�1cv�����U�B�U���ט�[n�.�V�Ȼ�:��t++iGj��m�8N�I���䎎Ò���6C�ʎ���N�EP�Y���֛� ���e�^]�-駏X߄sl�pe��%w��FΘ)��Z7e&�e#Xڍ	e��s��8�y��B��:ɺ�sC��0����h�(V՚j��mk�+8]���#�
��֎�hrH��h��m���%�Mf/���vW`�j+u;����Y�� k�d�a�H ��j�̫�R1J�c5��+���e%�V	4��JP�4*X�*�ZwL���fQ���I��P�ئ��������b6�t��u{x*E�f��Y�-B.�X���oM^�Ze9��<�D���4��R�TձDF^3��Z��:h�n� �HV����b���fhJC�c�(�(PvV<ݢ���Aي�m�fTr�<��*�h��U�r��[�b�q�/*��Z��cm̈�k4��J���=U�sf�Wu�B_Z2����[tfb�R餕�����()��݃Y�2D,D0�S��ēF�$Y3�fVB�F��1C���ʱ�eʹ��=��cDе3K3sVa�x�xv�JT�R�WJ��0��l��X�l[���B�o�գt��w�gAh����\Y�T��H77f�Vc#08NlQ�1b�����j� YR�P����u���
�NV��U(6��'Y����znȬǑ�`Gm�"q�գK:��HT6�V��)��;x�I���YKbzopRصYy���˴��kwkj$��5�wn�-��W1yM�EKa/�p9W�j奺0�//o�h���z�zZ��i�%�me�O[�hYa±7v/&ՊT��R���ciRfݬ�wt�/--�
*�%�Vkb]�\����l��5{�P`����t��cڸ�l�n��I蠅a�����CT2�Ku֞�$��@�m��z��h��)@�⺀;�5Ҭi��vM���3*M��h��m��t^�8��v�����yj��OZ�k8�^�n����k4[H�ל�2�%iᮙ� %�U��.�:+m�[�7&�w��xn��b4q�/l-��ePc(�{m� F-jF�ͷ/_�сe0�摻1/�h��U�K֑�Y��E�����Eh4��R��&8�H����#vEf���pK��h�d
��G$��C4T�m]�7�kks,��0�X�V�𰥇��ʽ�t�oAm4^�$�b軶O�c�7V^coͅB�Ӑ^׶����$�a�ؚ��L�1�v-�i���7��1T��.�è4�Cf]�n5`"ppP�y�]bYW���x�Ygc[�P{�.�RaȎ�6�h���ٛHQ߅��/XXD����̨��V����kjh;��N��Yh��"��"������*ԑ;&D�j#��:n��M�	гyM>B�f�A�*rnj�Pn�$��[����Yn���܃(Y��;a��E���+oM��LM�o2v�'32��jF�R��X4�y�M���.�{����n!�x��5�EJ! �Y$b��K��4�����j�ob��qkp�Ķ�&Z��]�T�VB��X�K�MH@�e�ÙX�Űfڏ,<��M#��gAٹgo7M,��5t#r��AL�7j���Д1i6��Xm�4�2��ԗ��4bk>9��4Դ�B��r�U�/Mx⼣�a��g��T�&0�̺�V���eҫ�%L� �񘨜��gը���Ŏ��W�Y�����m#7D+b��J��E���Sa��g8�	�$���|����v%@%y����SD#fEvFbK��:+-w5��o�qӁAH�k����Sш��'z�����G�N�x��k�����=l�·���fk��*���^,u�+�K�ٱ^h�e�BɆ��i�.^,:�{P�{Nn��E ��l�)���l$�Zm�[k2+����#0`Sѹ-i)ŭ���nw�J��y�Z�Uԭ!��}N��^�a#��ܒ�G��n'ER(I����T(�6��A=x��m&nnMw�1|�=���n^��	��Rݘ�Ѹ^��/hjog�SG,�#Y|	��Leh�+.�n}���N6��P�F�"�8V�+��!n$��[�vq��8��i�$���;�H&8��u+A��Ҋl�2�,$��2�ɤ�z��\�\QB����+�t+ade�+E)7퍸“����X�Z�^�D�:u��~�ӻ�[�kqV EcY�ፌ<K5������Z*!m��SS8����y�k"� ��ͭ�����)A�B,1|P�=ۡ���f� .A�ykk��f�W���U[�3HG��4�U-0�ŭ�f�����36
�)Mm<!!�K�]2ihz� ��Y��YCf��M	�mVk����(e��"���R�j@��4Ӌ$t&�7#)n����ek� ��ݼBTl�Sx5i;Yq�`[��&�{��Eҡ(Ǳۀ�E�W���m<�І�Y����a*ne**KX6��zskn�a�81(eEt�b�u��ص6C��dej;�Ee^A���AI�*Ѐ� ��Y��.�vra"���xM��VgEn�{7D܏jbR��]m��J$[��76U�ՑZ��6�s������;���tu���L���`�*��utXW�V����T��gRVS!�Di<��u ھ_0Eh�[g�f��S R�Y4*�*J �� p���u>G�e�+\����ZBφh֩ZՅ��c=�
͢�N�y*5k���weh�U�M"��غ�� ����F�F�̼���;g[՗��n�7q��-��� ��7M�v�ϳ6J4U��re��]k�(��{� ��՞�S����5�C�+;4�Э�9X��,�,X��� {o�%J�%��J�(ⴶC2�5+h�R���7Ĥ�ZC ��Z�f�N����t��V�tm�����sx䫺j�Ģ�nnUG��u4p��KS���u��DLմ�k͖�ٷ#Ȇl0�^(^�;���>'&܂�"�Ѽ5<�Ł�gh��Q��ͽ�k/�#V�_uX)�w���m��M�%�ĩ��4�+����K3�t!ISV/@�Ȏ�bn�-TY�k��}]aR�zI}d��X�8�b2���${���6X��R����%6v-bFʼE�>2-��iʻ#j�A�Y��2���)���4�í�xF�5���٫�h�nj5qz���qM��)�L�Nʹɛ�3���塋��ޖďa�4\���*f���.�C&�m4nP�S��N�j�ƾ�k5�_T:ذ�ޥ�3���M�R�\��W��N܎���p^�k�iSgp�i	Q���4^.���/.�y�Qc�M�����\i:<�,KU؇�ĉ��7Ӱ]��-G~�f�(d-p��)�~BRҝ
Yi�r�3�1�P�Y�8�lp%�.d�7�3������F&�M��VcO�"NMyfZ�[9yP�\+;Q�.���+恦�8�]g[46]k:����y�9{�jxf�t�*E�Uo.�V泊���J� Yu�C:v���`�+�L��l�[�Ef�ˉ�m�9xhS����u��=�L�Z��.��8�؀�.u<�8��P��h�ԑ���4VWkx�id)vM�N�Q�9��tI-�L����Y��ʘp��[F�J6��^]�]�[x���Џ]�ॉ�>�t��h@�YKV��6KO�V.bnWR�V[����ԁg#r���i>���h�c�p���58���y&n�]�_�i��#�r��
��D�s;�;g)f�@�p�c���ӌ��1��L*z�m��.*��97nf�p�F\�j�R��w�ɝ�v;q��T�\<F�2��9"xD��T����Mf����Ōx:��U��	�O�����O�|��.�ZX�j�Jm$o�"@�4�׵}F.�V�������QL�=�z��oSսO"�]���]3@7���g����{�m
�>���u�Y��)�1v�hz;���A�qwz*Q�����s�#�T��1�5�Ķ���΁s9ٮ��O�;+��c���[�I�Bɢ�rtI�!�"��������.
��0�;/(N|
�����u=C9�ٻt5��]�C��Z�:���K!�d o�����{�Ӂi)v�,���s���s/k�'F��:��6�"ݦ�ysU���m0v�*B)h��v�j7n��lJ��h<���X�{v�R�ut���^��GK9}���F��p>z�mPF�Zј����mfp�v�|~�``%�{;/L���c��>�>��m�Y�]�oL<&
ǻM�k��&�hzI�5h�"[���XU���u�`T\�m֩�BFY�f�g%;��^X����ݑr�T�;�os�y����N�+�C<M.b�yy
�.�Yw}��e�c�m���[@:�Bcwi����5�V��D*�|��ɧ�aZ�e5jQڗF�Э�([��J6ᬺ����eV���O�L
 �n�8]����>؎PQ�*`�S�EҢ�1^c/I�d�d\sU�"�t^�#�f�ЛC+*<�Q�lll3s/E�����>O������j4t�$��l1����G�a����@��:��(
�z^s��Q�� �tk8Rё�Ml��rL,��6� 1�����e�Mwך^9X�*�n��|�S�]V����c��ܣ�lnw�/R���U�3t�}Y֚x4Ѫ�8�9��y�:L[7�H�Ki���g�ѸL����=%�▵����0bŵ+�@��[��y��Z��;4ʗ�f��:9��.�p�N*	�hQV�ݡ4��m��O`�;O�̫F\:����u���BN
�H<UՂ�eƹ����Ŝ1�ʽ��m�*8�I��曄TK]9g֑�f���n�'��n@jq�Q �K����P�}�Ooa).l��s�]%���M��!Ć�%�q�Օ�j�	
����
���ܡ6RS1�dˍL4���,{.&�
ȶEգ��Rmʒ(M��f�=5;�uy|]��:)����eZ��܁O��Z�A�Ν��q^%Z;�X�oip���N��u���s��ce�J&t{N/$«n�|����E����yR�n���������|����l�Y��v�)KT[_fQ�*_
���a�׍�gE�0�����ЊH�gNl.�3i�3���5��+\�[���ꍦ���zQ���-x1�}�s��t�-�*�!cJÜ��5Vʦ��R�`ޮ9v�(b�aI*m��XB����7�ݍ�R���>nfRJ^�[%���C(7K]��l�[�/��Z�^M	'�~]:�.<�[p�YO�6�K�H������@��t���%��w0���en�\R8c36Eֽ+���X�J*N<(d���,K���9Q��b�s^��i�f˭r� b���r=�K�}5���a(��n�#)u�U�4�]Y�Z}���t����[Eڏ�3ջ)�J�qܮ̃e��r�3r�3�>��=��/���5GW`�$�%�cC�5b�	�sT�&ڛ
���7��ΔW[ڧJQ:�^;H�fe��ن�і��y�-�C��VZ��cc�.�h��\*��ˋAO��t�V ����NV;���0>B�Q��;��ֵ�7�C�ګ
އ�r��0��Ek�2�v|�ۄv���<X7E͛��e�!Q�:?̰��3;@���U$��Zr��ػr*
�πLӫ�t��-�OeN��P�R�n�'C$T��ފ`y����ƫU�[J,K$w��:$��Zʼ��E}��#�6�'x��i�㊣����/N؈��,��"Iʿ�-��;\�:Jďou�9�8K���Ԩ�N��-."�z�F�4n��N���׺�9َ0�o����y}�5�[#�.\��=*�L�Y�ky�<N�"��4�c�zP�-��VKm�Ay��F���t����]ڇ�F��9L�5����V�J��K�,�Yg�-Wf��<k"�a�uR���=ܦ$���#^/;�K<��%�f���^A��F���Kt�#���U�f���ǠhZVm��kt�<,vU�̖{"���� zq�|��T�*�4StS���9c���8��W×a
��`��C�6(�����)��i�j��xړ���QD���|c	��O�;c��JҺM�Z1���:�}�J��"��ȷ��ƛ]6B��쬃Mit�r�J��׃v���\����)�"i�S%�)�rn��Ɇle�l���FP��z>xc����6�}PC����̖�vVa}i�XOAU�����	N�rͤ���7��ĬQ�<'Q����j�l��oFFE�w:Y#{��7iU˂CRQ�8��,�긆Ίj���V���.�n�%I�K%憺�b�8����w����ұW\5��9Ɠ�䁦:�[�>��\�po*�!g#Y��S�
��VW^A}؝:�Y���|v"{C�mVŰ���
���~�T.\�^�Z<!6a
�恰��$7����ʄ��ˌ�WWg�hl��^�,��Hu�N�dS�}|�z���i�Y\w�GDq�YV�T�n���l��X�HޭYNY6�YLm��&�H���}7���P�le[��r�٩�
-Vķ�vqn�,��k�+z�Ȉb��gu
�8Z�w�E�	�d��)�5+�h�U��n�f�^.�]�F�$k��s �l�U��νoE]��͘Xe@6�)�_;�7�lO�5ڀ#%n��N!cgDی]�Q�H�nec�J���>�B	�����Vګ���B�!�p�#��i�{6h�Ʋ���ԅӬ�O;] �v����Y3"�ԙ{65�+t�GFn�}Q�
����҈E)R�{vWK=�3z�e�!>:��E֦��R��̻���+���Nr�Z*e�l�UZ��VN1w�}bJ�w������"��ܝ{x��L�gM�x�� �J���"�oU쩦�eT� �2�Z��ufD3����D��67�+(ڄ3}u�o�giE�,>�Q}�<���q��rĂ�줵<tnQoSs��WP���F�_�	Ek�&�w\ԼS���u
��3�:��v彩'r�Ws+j*�u��r������D ��Vj�4��-�gt�]�B>S����jT^�'۪����{��TX�e�R�Y����Wf=�]ˬy�9��fVn��1�Ӽ��1C�9K��7�1�JP����i��a �Gx�9�Fua��TEk�|�r��K,
;Y�l��.q۴�
�*T۫���Yt�ǒ��wJWi���(%g���ċLe���vN��˞ժ�,�* R�+��!^�\m�{K�id�%8(S	^��ZQD��b�7�k����z���nW�ܕ�$��������)Y�ru�Y��{m�2���X�E�r��#�[�oyj(K��	����/H����ar�J���SCv���\V��X.��G]ER�c5���#�u��9}@a�R���ӱ�r�1^�N��6h�]�,;q��n%��K�VL����W_]�('�rh��l܉ޓ��c�c7[Z�.�g���d
˧�8Ě5�LJ�*�]<�]o4mB;%cA(�v!R�[]��10�rg,�n�D!�F��5����Nc�JΖVî��KyN�P�!XI�h�nvEB�d�b����J�5Фv1b���}���{G@�������!�`�J,�ۨ�^��0�7x���Z5q�ndח:��.*��Ǝ*<����Z��4V*��?�ݗ��ZkUJ0˺��%+Uff�g��v##vgV�,i��}�O�N�*ʘ٭��F$.Mh�Q1�BV�0�P������5��-���-0�(��V�\�8��:�R@p���}Y����t�M%R���E�*r����ϬS,�/8cݕv��Dd:�_5f���!�-P�o�p����ĭ��8�6�!z1��C1qmq��섇��ԍ-S�p�ˍ��5��;�	(���f1��θz�����n��)�����d�k5֦�ͤ�7y���Θ��c6��%��e�f��\HW)tz����m�]{����!%wr�V�f>(mt�u�ع��:��/U���d.��r�ھ������L�Cyw�Z�x���h��-F���}�H�M�����폜/�ӭ6��=���;c��fb[V��ʱe;����pP��>��6n���y���ŝ��=�p�����ΫN�F��o��%k7J��;3��ty���#g,�\*C�;%���ŋ�6Rل�r��A�Q���
|`��^��a3.�w+dT��3�$�B]�Җ9-<�w�����ᠷeFer��=�QmY��>J��Gߗh��j՛�6؝�.���NB2]�aj����Hgr��D7%eY��l��,h�)���\krtTɧ �_�Nd���W��J�kKΠzM��亐3�nj�c�ݐ�|��y±ݻU�A��Vl�f���[;�y�m�Sz��dY�g`R�`�<��	�+u��7j�c�{qh��BeR4.��J��)Ԁ
�����]����6�x���Y�vJyN�om���,���Gv����j\���8q�a�;fv7vk)���:솾%k�FM��J%gw�\�̩��܆��v��0���%X�U��U�"Sug|� �ˌ)�{n�gsF�3Y����eWN�F�y/wr:��˦�v��;�
�,Xv$��Q�+j�#G�MMLS�D��U����,�����SWWd��|�4�|��j�k�hL秈Nɻ�R*}�P��X�bp����ǳ,eIQaR/G~^�Wp���t?u>��ޠ�!��3���f%�����g9&�+m��wkޜ*�Z���8gX���(\"��*�&ƺڕ� �t�msn���ϓD	0wٶE'��k�铣1)���A����~�����s���}9ˣ��ZE\�]�T.�]��-ȼ�v��9t�"�/o^��=�M��$OC�e���և6�M������@���x􄂭�z����[QSځ^U���[�^k���WYź(r�h�YL�6�N���մv�9��L��1��f�6�e����H�n�ĕ,ƃ�\Q�-̔���3��%a��D\��UF]&=Vh^-�j;Iο��S���qu ��@�N�3DYx(N�M�*���ۃa�>.m�
���C�,�u4�m�z����:�9�]]���ٛ�h�R
<��m�M[���P�-c�����[��t�6�7�ca=u1�nW<\�e�Ia�7{PUر�T�%���7dg�B����vK.�U��5��iT���-�
Ʒ�y*��:��sE��h�Sq:��}1�^��I���R������R��6��Y��Q��d;��dI����%WT$8�U�v��y��%l ���1�?�̙�lW����g��*�)F�����Zݍ��t�=N��e�7NKu)�F��ʦ��μ���4p��fEHfU��ś�f�Ơ5p�Y��tu^Y��t���͢�^ �" �ݜ�-̖/���8(����:��1�45@�ƅ�-{���Bdg3�2w4B�tZ2=����F���ܠpW,x��c�)�Q��쭫a#�Y���%�PzN�''Ja]�[yKuT�"���G:ɸ� �%{��.t�� Ջ�fVT���2J΋�����=R�e�:����u`�/Uql����o�̨�>��8�_s8��H�{�����X��+�2o,!9�LO;ro��^tQ>�N֬�ks1KAǘ ,�복�Z@����I�1��Rr1��M&��$1�v�)M�FX,RU�v]�:�i��rq#G�JUN��e�:9Y��N�fQ�G���aU���yA՞���.Nx���L��to@���b����3��9:���B�g�R쑗�X���1cv���x���y�������f�ʑW�2�a���ժЋ�ÊTr��eA��]��z��)���K��.�nw)p���xh��uT{��O�4#�v+�3r,���oU(��ٕv��Y(;����h��+,e���a9�uxUcH�50[C�Ν��Y��>��tMf4�}���^>|�����ll���cm���G�����
���N2�[�t�r��Z٪t���qU\H�m+�Ȅ�����j��R�ǤLwj�3�rs1J�CIsYd�p��p�{�m������Z�s�+m�����ɭ�C�r�ֵ�2�Z�����c�R� �����b��V�����B�v����"���2U��n�7o:NW(���}jF�m��2�Q���Hcu
�wY��T%*���� 功=1�ecٝSE�u��,�!y�R��C]]@�ˬX'XifJỠ���.�λXC˅��X%�L���áN�*l�5
�##U8o�R����U���\���M��R��[�s^��VZ�	��Fwo���ީ@V�Gh�,nR�]�Zp��(=�~S骝f�IF�**�vc������hw80X�W�U��9C��B����v�v8a-f��nm��TU;A0�IV���݀����Ėb�d�&4k�#���,�S�Eo׽Hq��׬ieJ3�^4�}����9��u]EF^ŀ�qc+�.��[�o�,Ok�Z��ہ�8�w��o�PExI5ȥi)gVpCgG5K|��E��r
7�$I�N��86���Qk�͇�n���++�7+V�X���C�xF��],�[�e�����n��SiQթ��y�q��u�F�b�j���9�(�Yh�� �h�� ΍��#�f-v�*��_V��(�捱N���ȝ��J�$���p���Q�lr���K�$��);@�Sw�!ϟX̐r��K�PJ�jP_\M��v��%Z�O��D�)�mkO����}�L̗�aY,J���\Mf"�ʜ�����WٙyHڊ3%�+W�V�Y2�!�Ë&�y��W.&ڕә��kV�ŋ@���4�3�"���/5V�0gR�cK�9'G(�eE��)��0_K�%�������!�m�|��Ijv+t���6�a���/�x7}�k�k2 u�ZJ�k��t��M��_"��H���|֊�]b�;mXz�ruu��k]����F.�](��&�桐�Je���t���{����+�G�"�1jΚ0�u��i�q��C	ܷWN�Pnp��wF��i��
��e��qK�V��hbG+9��lҜ�L���(��2;�C�$(e|I��;w>`ن�$�<ˤo�`�qL�0:�k^7-�̻�f��.�p�,��"���Wԥ�]2/T���9EB!\d4S�Q�;��r�l3�TH�֨�1C�Z����B�@��Eõ5m��`�)K�&Ƞ.��H����L6�;���L�(.	m�V��<ޏz����*Ldo6/5^�����kZ!�.� �C��6q�Cgٸ7��
M[Ѱμ��@m�.ͽ��vХ�hɁۼ�ֶ�Ȩ_+VQ�9V�!YҺ����PYc1YpG�]Y�J� ���N���\a��E^m�bل�{>�=鷀��:�iib�V��ĻQ�X�;.EyU�֩�sn��4�j��D���Uc��*$�T���6�3�|T�+��P$�w
�|`�����魱��K4&��9�`Vm��!I�̲�g����-�����[
|!��줷��d���ՃWK-�t5ٹl&^j%�A�3��k�Y�8�ȚWG�k�Xv@����Ond1ۭ�oZ��5�����Z��u��:_L��?NYK�ʦ���(��a���D²���q6��G���Ig��+_7'nL�шqp9�󔫊��\���ZM�s��vTӉcDVP��E]�<=�)�t����YҀ��`�1������b�=�޽����6F�F�Q�6U��k v_C���c��+�㠱v��`�)H��պl�� S�
z��W�~ٮ3�B�˭]`�6h���+�M�a���՛�l�F0����3��Á���<��f��,v���Rˀ���{x��˅t��*�h	��LJ����%t'�"5��>8v�_Zy	�{3V7����Dø��R�d6���D�H�^Sig�U,�����es}���l�{[�٣r�*5�Iwُ�����ॸ���T\���%;r`��ؓ��j����ukr/�`�KFx9�wp��5�M׻T����q���(f=Z�"e�s���lA�w����\:�f��'��Y�֞�����c<��m'[�P��HGڈ&�#�V�o6�{v.�W��a������7Tzm�W"�(ںLN����$e>7�D^X诖�&V��nĬ�6����H:�8ɮ��V=W\ѻ��(��zZH[N�kmc9j��}
]�\���R���]`u.*�8\}ϙ����i�٦-�f�AR��0|���|�_f���GL��KPb��9��6�WeM��2u�]�L��¸�ut���h��r�J�s1^I��e.�wE����2��<��NE��-t�Y�*>�w�,�����v��$��lP���\]Ըz��b�|;��Jͭŉkt^ƹ�#��0SR��H��V�6���������]��τs��Y�:�3g��V֏�o��jH�FM�\�:�^#�QQ굡]�}���eqQ�[[��)ѣx۷�v�=�f�R#�����+��V� �c(��`B]�Zf��̹�f�S�'6�9�m#�-�8u�f�F6�B]�:�)�Tk0�WMK����&p�������@�-S�(�ef
6�)hb�2�ʜ����
��+{��eN�%��1�0�2��3�ۣS��+����/��h�J6��'�ڙu0��ى)Օ�d�K�ͫY�� �+Wn�
��"`*;�v5t1G�F�q�+��f��^r�[�O�j7���J��t�q=�>�bQ�Ȱɑ�7Opvv>��+0���E�1�n0�c�̪46n`�D���G	(�U�<� �ctm�6���p�h��L$�u������_pX'�<�i�1�{�q��]aI'��޾��i��2�$�wG]�G����x.����>�Rjս��Ut�4V1ԝCx|$J�Q
t3�Ch�GQ�w9˄�;x� �6�\2�n�ܫ#I�ɔx�4��ۊ�2E��np��ηl��zb�V�g7���T�����G�H�m������;�Ѵ����i�V��Ko����D�ɮyi ��iDv$ҕ��J�r�1ݴ�j���4��WM"#D��;�ۓ�Ӧ ��&���h`S�]F����F���������Dk�$f�7/�K��v��i2�D3�5�"f�E�k���u�t���g;�t�V">�P)Bv�o���따��X+��,�d�n%�q92�$a'
�3[T(U�9u�����j��)W�w8c��.6���F�uiSO+9NsY�i��7��y0@��yL��P�1b=�g7����u� BY��j� �K��]���p<���ӌ��kY�(F"QKP82 ��/���������ӥ\L�Ლy[T/ra��o%��(�TT���{9PPQӽ�n��hmdb���:�wK�t\p��{��t����������V���j���R�k�M[�ԍ��r�|�ByK2 h�zB�/���H�'��(���t��<#���]�j���y��;�K��Y@�l�f�X�����L�f�S��S� :��Tڌ{���x�m�(7I�Y��N��lQU��r�{��W�J{�C�͑t)k��:=���@8���T��{@���}ط���W�u&e!]�f�ݠ��� J�x��=�V��K�X�>jjG���5�i�,a�ٜ��룹a�>���S�Mp�n��J֜��ݷt�0齍tCR��=P�l-a��.�m��D��]��h���hԚ8�ޚHԧ���Y��>(�²�V]����J!�����&
�hl��`؇�AG8�d�v�f�P��Z�ßcgf���X&Ĕ�\��1f�
54�W&�VŸS���x��{>G��� ����8'`��Rbm����_0��R�]�B���J�P7�zb۹E����X����M���U�-�m�z4e�(��b�����/Jy4�/�o i�1�X��۵-"d�(��fi,7��n���:���f�S�.�ᵷ;�����T�K;R�3Z1#F�����f�wyO�VaΫ�Q���`w�:�3�鸧fb�gp�1��(3�9Y�Z�~��q��8�op�&u]�G&��
mTՉ�nh���O�=�;��:�"�Rv��ѡ�c@�0e�=Rl{X���wM՚�X�%�$Y��q�G��->�<��·y�᳓8��� ���U�Du�E<M�p����.���M��pMhDXv&GnT�v�x��V�ij�D�E<�;�j��V��Y.#�eK\j��7��x�:xѵ�5,<98�.��pn�U�x��k��BW��8�i�x�D��+�R�U��5 � �\t&nj��&���a'v�1n�9+0�1MA��.�ͩ�XB3/�����7�B��9�IP��0�$�
���y�XTN�F��VȖ�ŵ��-�D5�Y��v^��t������@;� �(,bY٧.]�stW^L��M����L!�5#rZ��m��[���F�1,e��$y��銦^E�s�"u�wIн�t�F6zX؜�4��J�>��Z���n��B��ڎg-M�О��31#��2�ka��,ʱ�[�r#H��0�������Z���<�!41x�/�5���[��m�9x��0AQ5�M��������ٓߞS��EZ@qX��0�}	�*xen��
Ս�
�n�QN
�"��9HրR	�hW�u�qp�y;��5�dV%����#zovK�,�An�ر��1�ۊV*�qZPf���#���ݤ3:߄���R���̶�j�P��׼ٺ��v4����ٔ:U�wY���G9�.��vd�+/s{
i�$�d�|T
���� �G�5�te�p٨�D�)#a�ւ���ʳ����%�)���U�hj���px�x�����`2���@%&����Ӡ�͋�b�K�ĦZ���|;R����ī��uq
����Q��b:1�Z����L�՛$�x^d����՘$3-��i�<�m���[�P|iΧ���n�YV�*ಸ`�ܳ����g'V�qv�&�.tJWy	't�]K����ֱ�;.+�F���T���%�Ɵs�W�/x�MVs�,+AUa�t��KVS|�q�Ż�C�
�b�k�v�&�5aN�
�k������rk���dF�w�N9ʠ9������Lm̔/yƷV�R�e��[�#�z�J.�t@ ǀ�f��ۋB֘�������.�+/eoۨ����`��r�O�f��E��vEJ\5+�y����C/�&b?k,��W)��#nq}�kλe ���V�J�m�n�(--눷��x����ʧ���c-ӝ���u�]�s �P�̝KXCs���A��6�9�f� Wfe��\5b�,[��)����&=��L�͠<� �=�U��^F��(2Τ�wz� �J
z��OM4�-B�SR�gT[E�e�Ф�L;����wk�鍚�x.n�f��L�tF͡x��6MkF���]��ZQcJ!j`}��\����@!W�� �eث�FcK��Jc�f�\��^n�,�ڗK��}�xs�m�9��$�#dpܽ�[�T5Ɖ��i�k��E��~���v��t�A�*��w���۝�0t���g%H���-���;z;���I�(m�� YGy���MM�n�ӗs]�
�;S�֥w)���k��Mهx[[��(ݿ�M`�W�i��y,�G�����2���Z�O١��N��f�\�aҎn_���]�2�,
wz����t�U"ۙ���+wi��QO��efL ����r�]Ż�j�����5k��k�A[���\�ӥ*Y-owol�Z�Z�WRwK����lW���k�X�b�x���-�^��h�f�>KZ�>UXG��+1�������%Y�F��
��\$�i��[�'���c�����=�.���Y�}�P��[9��q��\c�a[uʈ�6q��u�/�'��JԜK`E��rV��S{�/�f�c	��{�fk�K G{+���E@� Ƭr��f̍������|@��R�-��g�ƅ)f��!�r��b,[ �<։X�7yȅdٝ/�5��Q��kB�۵c�U�F�h̥�}L�Ø�Z���!�a�κ�'ѡ}�8N��N����*B�����n�a��Kc��
�V#�4�P��o'JՌ�sx�M8�(��Z�6Q������+���9�MMW���Qb|���:ۉ�dѓ� �,Z]&�282�+Ӭ�FC+2.lXM��lҺ�2֖NЮ��M7�5Ζ9�;QXd^7iqe�Ë�y�j�nP�-2��Q�.�#a��+�/_uŲ��#e��j�I��\�7s96N�F3!e���5y�GJ���}Z^X��tܣ(���F�����K5�%3��"llF�<��$��VlHFƻF�	�Tq�w;�ݛ8�`){N��hA6oG[������%JF�4ѽѢ�X��sR�l��m�����m�P��y�n=���[���X���P�+�"�~�˕n0g]�W���%Ͷ�B��
��cO7t�ϮE�l��l9���OhR��X�&��Jڟ 6U���cP�eĕ2�۲>�(��ّ����&�\�/�춭��V�ֲpf�U�d��Ϯ>����k���OAo����t��7�YYy��*�I�����sD����j�Ap'u����#&����)3�v;��A����\�Sf�t�]��	�SN��f���k��qkիe��q��<S[yY�%��t���?�W�W�U}_}�}�'�_O6�TVd1�6� �ؐ�;++�u����lm8�"��gw���S�92⮗�Ӧ��Y�5ӣ#3��@�w�ۺMKt��w�U�q�T�� 5�3Eb���B��-��_]]k�N�����F��EAw�-�����ryxv#93ݩ4rA�w��Sl�µ'� �ݕ�̱�j��a�e�Z�9��2���Q����ss�3٫��N�Qt�1���[�&/Ӫ�<��o!���_pʸ!_�U��wƬb�K*�b5tJ��*Ō<Y��k��U���u2�k�f��R�5g}�ܬpײ��Nl�6 �ua�gW)��}rPw|�%����`;�ɩ H�'���\a_KG,��t��=�J=9�fՋ��<)� ��m�'m��x.���OM�e�]v�RƓ->��1EH�;<oL�Yy�̾Y��%��'�6��г�P)�����K���!�y͇M�A<7�m�"7�ZC8.�@D?��Q#C���b{�A�bΓ��b�K7ک��%�`�9ۖ��&�$���R�6<A���e��'!�r�L9M��)�B݋8��3f=���G;Q^��2)[N��/C�hu`�Լ������T'<�Hi`����:ܺ�J�ۺ5�e�ylX�i�!�uDS6�n^OG�X}�:�:G�&9���mu�����U����(�E^�ꃨ9�Z.��HR��'��1P�[��-(��U��rC"QD�D�IR��S��j&L7W,�C��L��,.Qt��AZ[!*�:A���D��a�JsTY�/q�!EV�ܬ�wEc�gS�G�'5\���䈩V�1Q��9I̱2B�M"�CBE�*h�s��ʊ�^��v�B�]Zif��Aq�J��K$5]�$��J�B��r�Ι��
�D���Naa*�h�
�����a��N�
%P��P�TJA2@�f9����V�d��fay��4-D�H"q�n��U
���I#W":T�"�VT�g#F��$���H�"����*��`a{���;���:{�9Z�ny�'w]��ANG%:��I��]M�aIJ����H��W��a�uf�HG���#��}y��ʍλ[XlU�.f���g��ޮ�tӨ�eX��j�Wò��za�<��cb��ʮSo��a ������C�v������:J��]Q��n4-�f���f�I�.�}ce��qb��XY����s�j�LLW3��^폢�m�>-�ג@�
����E(�*�I��1�y�)�_Ui}΀fc��+�O�6tG��ׯh,�ʭ���V|2�[�L*.�7\�Y����#���t�/����
f�3��p���\iz�R���D��/�ù�Y��g1ή�ᑱ�o����$�D��n5��yӨb/Χ܄��wM�w3�B0`���*G���3�Z01	�O*��T���`LE�i��;�T�܅u�@�8�M�!���֓�,��ߞl8��,�����:!W�X�5��@%�]���l���S�b
�b����@5$�Kr��c?M9��� 4�2���#�`@���t���G"�[���I��n�ڠ���q�y��ܫZ#���iT(v�2�������)���r���I.��q�S"�/�ĻR	��!��Qo�Q[�l5�@bI@O�O39c�f��b�^�#q�Rgק���]R=�]5�k�j�L�HtL�p��i�~��5����&%,w�)�.��w|���q��nC��:�^�Y���K�Fʫ��%^�&u�p�ls�Ρˈ���]�sb��fEy��_�ू�z�����䑖μ��l<>qʫQȦ�Ƌg��=v��r4��/��W
�A��PN6����Yzs�.^䝛OH�5�Hj^�[�9AN�;�-���{(n{��q7��0Y�eu-�+������n�x.&��s��k��S��XQɫC<[�O�����^ O4mV��~����e�͡R��V}�5d��~���)�J��F�j5)����ؤf��^ߧ�Zl 4_�lK�P�?h#�Y��{^5S�Y��8k41�������+����Ʋ���M���݊�I��(F�0���|5�h�j�=Ԧ[���z(ZBߏ�Z�.N��/>�9=q��7���3�B���Vr��;F���� �����\/ԕ^��p���^��1���:}���!#]xuFU��f�ln���G:6�3���5xgݕa�Z����CA��@�0�FY�g�f/���-�����1���כ�gw�A�(�ۃ0��j�^���q3)��H`	����a�c,��i��vL���P��x]5q����G!�e,�@u�B=��1e�������TF�0�2O3�[;��u�T iu�<���f�e�̙w�o��/L��2�n�ȓo��?B�v�X�(㙙4d��i1�����s"�P9k��v�a!�{�� {Wxn.7$�����滣�8�~���VֈO�]%�A�S>��o�W�ޯ09\�u��NB/���tQ.�W���p�g�h����u|�4���%��m�5Avqyn�O�3#�F̞��/x]z7���4�`ۘ�6��Vyۿm��0h�|�u�\|2l�C���V��"��TrQ�R��kS�=��j"�M\>�6ϫp*Å�c#t6R�T�a'A���G	U0[�󄋉R��yM�r0�Ø�p���N���{n�9�}:1���C�� ��I�G2�"�p�O�&廎���-U[Rm*q��wu�T1%i�-��%T��x��A�2���?&7��wnɯ/W:ە�٦|yk�w=�.Nh����6�؃1�$�"JDBg�TGT�:7Ț�,C3E0�b�0�מs��a�I��O
WR�\�%��5M)���	�q�`bɺ���Jاuب�S7$F��0�T�:��i�
�ӳFۘ�jh�vd����(��c���"�V���mU�K�Y�sMʗyY������!!,��ua��R�'Gs�)�&�mC��������\9��5�W��glB{yt7cy#M�f�Zm��b'R���*b��׋���=(�T�k��!M-]�vѻ�5�s�e<���"�Ok�N�zo �ck]ߐ���E��[,�o�S��0��|"�Kq�UL�z�ԛAn���T<+��_���k�jy�"ֺ�T���t�Ԧ��C�)SԶE��!���������+��h��WJ�s��i"ϯ�=�#=��{�C�q�<Cf7�F<�v��U�?�D[��uC�U�[yw�*�S�<g��v��%Y�:�)ʤ��w��<e���_r��h5u�)��`a�̖�^O�����:KS�u�օf�ҡ�t��0�W)L�r�g�Ƹ���1Q����½/��5��x8�I���O��,D��2uPediuadiu�*<�:B-�T��3�c�0�]�t6��w�=�'N��3�4p�x��G���n?*<�UB9{�w��0��c��x��i,��i�z�q5}�@0~���~ Dg�C�ڔ��WpY�����
T��M 17{��n����6��iΈ��ss�! z-�G�<�i���N{�asǸN��%�(��)F;:��5��J�؇�7�j�jV[�.��G-8����`0C�L�Ŵm�K��v�}W%\i�SWB��}+:�K0���W�Y��ks���9����}��YfT��%�7֋�H[�+��ɹ��=̧Щ�tdԕ���S)F�lK���#v��-�#<W��"�>Dm.�𴍩&�
�J���l/=z��@=)\�M��uLȨS%)��S�dA��&�//1W׻�Zs� /�Y�iZ�Cr����\��C ���R%t:��*�f�l��27�K)�=����̥ב�86�V{���徊C�g��S%烖���C �ɩ�Z�J�/���-�"%%�@2���un��m�1�q�p�Tj{lcj���W���f^57��;���[�H�`i�]�á�?Qx�C��,�1����cCSx�WA���x{��w��]�\�]8({L�VL���!�e��*���[P�諻�0M#��^�;��E�-��m���L�҆Bu\��wpx��C`�`�� �R��:��\n6�za{��y�y��~�tBv�#�sݐ�:uE��Gq:�ݝY�1�Γ���f57P-��#pS�1�`G2�We^��T���	�N�21Zw�~uM�ȅ{�C�l��5��ܝ7��O�[=�;��ý�I�?`��)5��)�:gp��֓����,��'
��n��ݲSs.�<l�`v8뗶0$���Ep��Xb��8f�6Z���P���(	�2����k�͑m���pm��������!��;Э��-�N��<K@�����6X�5��@%��Xl���瀬�'���c��{^�B�B;(p�s�ʙ�r�:k�y�2���%Y� �Q�]�m,]d11Uk���ŭJ���\����f/���ᥭ|�Pp$�%�/����o�1�O���Wt��Y}xw�\��\�BjV��s����gz�\!pM#*�������|�T��ဝ���Kckl�Q���E�u�P[<0_=v���#O^K�sB�RQ�Hѷ֕tL`w s����i��D-$i-����Nx`�m_�;�Cq:�'�8^��&��̆��%���s�R|�*�8:L\�}s����ɪ@5<L]˖2�����竀B�q�8+W!y �#Gd�����\�z�+�јƭNP�ᇲ�ڞ�e�≒�] VL�Ѱʓ7�O� �����K��Wxi ��ƃ��~h9�-�E�%(�qp�m�51#�d�&��n����p�$�t�=5㒄T,(�n5�l�ں>�� 9��l>��QT�����j��L�Kq�#�OnR��}��=�5�F�-3즨ː���}�~F���EU����oQ9dr��h�6+�(��Nێ��a�	V���2<�QW�7�7x��O�Qr�"�[h����%cި&H���g��Zt6��]]B�$�ч��Nۙ��QV�zhA^ͻ�50�N���IO<p�IWa�9�W[����1��矦VTjt�,����ʱB���˲���\��IN��:4��g�A�0�63� +q�1p����'\�^e���e�͎bJ�ImN�E��[��W��ݳ0��j�{&4S'��� �������\��*�`�[�_rޛ��^ϱ��R����TVv
ˀz���Ŵ�>'A�1�znp�.�cu�T7@��pi4��_k��
���c�a�66-I&$��Pq"GG�}�èqƳzQA#�㪈��|�4�`��g�9l��;w�OJ�E]>D��=�m�b5�"���QP@P�\=Q����T�S{���p煸��GSU{�m�!������gS�6�^$����$���+�Ⱦ���⺂��
,X�r���#�����:���{G4��lA�z����������G��6�=���'�ޗJ׽u��<R��)�/��0U-�0���Sn���BCÇ*�����2a��m;��#�X6T�ĢU����|�*�<�_�t�ם�]ׇ���W'y�M��gNM���BWE;���7�3���}M�{�����vC���kÎ�M�+Ω	�2T��x�5X4�F<�^|���V�V�e��r��W�r��C6!����n����$�g Ԥl� ���u ŨE�r�y�Q�=�:۱ � ���u�7	�p�.<\�%�`�4�d!NA��z�ֱJjRɚ��O��`��/�i�ޗ��S���I�iѣ��F��*�'eْz�f�`
�N��mjjf��ϔF.'\h�N�zo �ck]ߐ�$��\B,3M�vׯ��$MS���m�w^C����@C��ԃ](�P2aˠ�O��e��
���`ꡏ��7��Ҭӊ��Ú��Yk�.�:,�q,+���G.����
��U�QUak�0r����<<2�{s/�X����J���L��2���\����z+��"륃�(;#�eV]鯴P'j]A�Er�j�A\N�"�u *�e�-�/C�4�u�+�_�p�/��y$�(�ަ+Bty��'���m���6e�zf��R�`��Ψ5�7mVq��`p���^G7�#՝�X�U�Lp�ET۬�).�j�g�i('�jnm���)��R�Mz4!�m[��չz��K��V`��]a1ǅ�w
|>!_f]0�Y��{2�
���y2c�ek��'w�׋{[�ic�su��R�u���ԩ�������l��I,FD렊��Q�׀x���fS�� =Y{��w�H�gg�����1�!Wu�C�x`�2�j'�����rD�vUC�^��@��AJ��o\��	�j��I����d��rx�ITg�Cb]���wԡ4<�!�#�J�B߯й�w��$&�l�RypR�e����=�/�hLq =G��ʼ)�����nc;6殞��+B��]��n&X�6\��<��m��i�2��8�D� ބ����X[X��26�39Ǆ`Cx�b�����c	�)�X��m���~(q'���(�7(
��F��u�P��&KJhu9�3����>����[VY�b�*�z9s���[;�$;�Ԁ�gIUf�=�*$�rf���ԃ֪C�gϚ�K08��㴂�*X-�Ē�5@$�^�a)�"c�'`���܏R�W�aHԺߩO#��A���{=���3��[�j��� 1M�K�[V!��O@��,���w�p�H=�t|9���V�#��<���Xn����9kËVC*u�&f��ѻ�.RҚ�K��&��p�;��ͪ�j�HPR�&��� �fZ���=I5Ee8��g�5y�N��2�-�kju�TkoXv���-Bi>)��̣;*�)s+�}&�����*��[�j�rU��vlB�����:Ҝ�6=��iY3�abM�p2|�m��ks a���m�<ú�a>��O��l�ү�L���{u�EO��eo!�Q�F��U��7���./fʞ�a�0bJ���'G�Ԁ�Ʋr����n�wgV����`77����ܴ�f�(�`�a���
���%Hv`LZv����;�s-��SyW�w8ʜ��#5��x���b��l�>%���'{&uH���������"b�̍�G�=<��SYLB�u������mԌ��:H� ��}�W���	�����J�u��y=������X�,�w��J��S��Q1��N����	ŭ����H쌑�v/Htm1V���xm��r�d2��>cj�\!d�*��t������C1ּ��]��)�f㌴}x�����Ơ�x`�z�#̌:�2X�S�B�9�f^T(_[qu���M�@n��"bL=$V��S���Nx`�m_�;�Cr��D{�uI�&v�Y��|���B���'��X���qs.�Π��O0�{��yq�t
`�eê�<F٢�U�B��9ia��)�����rp����Վ��k�C>�˽B���炙i.�Ct�&[�+f�|�ݮP�9���Z���8�����c�Y��=ؘ��U��Nk����
�)bOJIe��}sFۊ�6���S��ui)K��]�	r���}��ܦEݪ9�r�Y2	�^�t[��G��y��U�և\(uK!m"Tvژq�����PwٸE��Y�7��U89Xά�H7��㓵WZӎu�`��>�t��{���MnF��r�E�N�L��.X�_w3-�O�����
�-���P�hFGgK�N<���cL�bĥ/�Ne� 5�\e
���!�)�Vځ�yZJ��%jģ�4t�yy ��fe�4���̥���ai��.]��]��������XQ?�(7���17V���"b]G�!:��c��:��J��9�ݛF-YٷLfҠ�!�)j׫���Rf��{K���Y1s)R�v,���1Ŏ�qmu��/�j�e�l�:���}��c��ul:�5��k.�i�,Iݼ�=+���ڌ�y�@���$O@d�Y�m��k�'/R��,[aQ�1X����e �u9����G��Z�Vޘw3�hóY�,WM_dH�a���

07v`�w�d��c����.�8p-�������6c����Ԟ_��Z�Ao�S�4P�)��ݗ��`�W3��H�]�ث�K��$?eہ�����X"����hj���d�O]�6d���9&���˾��^���Cе��t��;���fZ�F�5�Y�"yP˹0�mTE�`�^�Q�[�lgwf�b�[���;�k��m�C[6��|��g0�8��s�S\�3i\-vS0T���qʉhd��K~�վl��%�f��u���<���Z������ϰ��)�a�sl���-jT�M&vT�(f�w%���|a{(0X�����.��_q���Lܵ��kB�)f.V�E>v�^�Ϯ�n:�F��1�K��e[ƺ�d)��/5En���j'5t����>z�G].�Kr+T�j�X�ֹ��tc�Dˋ	��:���/e���@�_E7�^;F�Ui���-��Y*��L�$��с8�5׍,|B�kc
�{[c�0���xj�Y��d����h`-����Mޅ<
�4�YY)-�B�7�*��1����{�A`犊�zIˢM\�&�v﮹�R��t��9Ȧ�V�}٧�f܁"�f3�f6�&����w���J�I���{N;����t�sf�UӎK��њ��Q���Ј���=2�&˖�R.3��=�r���E^,N�K���5wt��״�V�A��:8j��4w��p*2�����9β$��3n�\V�XSgz_�u���'UudQ ��D��]+)>���I#�� �+wh�h�����JC�H�*�N\p�*�z�T��C����'C���*DID���j��HԬ�O<���h������j�Ir2BBR$���Q	2 Ȭ��v[�k��U�s�<�	]wC
��J0�
���QF��뗜�s֨!g���Qd�"V.륫�y+���Q�(��r�4/7*̥R��wB�-e'#�ezA���	K�VJJ"r"J��NA;����SRV��\�t�-j�j\�G��c�7u�{��Y�����Pj���EQ�P�s<�']�2-wr31U9��T�����.y�b��#L�1Ee$�C��G7Ow]�se;�rD�܋��U"�#�=�D�]i���P�uqSWG
n�\\�;(���TT�w@��;���i�"%RQS*�R�Ze��F�3�ZZ�D�*y~;����B�.e�:i�t�U�9� {٩@��� R��e���]�]�����kŉ�˕|_O���QT�b�Tu�}�_�T��W�*RU$©�[�E	>���
��������ۓ����������|��������~�yL>�뷣��^s������y�c�" Lb�sd�?l�SPX��) +��y|E}�����;���xw�[��O���]�<��7�r��<r��~�ϝ����F'x�>��ǔ���ro�`�}O�$G�P���@ {� ��k�d=A
�&�%%�[����""�z1�c�p�s������]���~L��&���������zBI�P�����z��x@����۝��S�s��>���AV*�W��U~[�#�̋�ih�b� �����"�H���"����ޏ��x����Uǭ����7�'��F��'>]����m�<��I����{}&����������_/	��ϼ�P���ޡA��T�>�?X3��?��wӝ;Ӵ��������;�����>�}B�o���N����=����yL.�������ӏO�90��wl�����>�����y��ϴ��/��}�?|���U!F{�N�f��v�|���ʓ���~C�a�\z�xW;H������o���'��~C��ۓ��߾Ǆ�P��޽��࿣�;���1�,G���5��#�|�>�s@� �����[10EZ���x���\s��^#��'�)�7�r�q��S�r{C߭�
�녟��ra�ǟ<yL��۷!뻃�N��u�������o�N��'���|�ߐ�������p����ʛɞ	�������~������o����.�oi�;ݏ����[�zO(xMz��w�9܇���q�0����O����®��	���wA�c~C����� �������V�Qd1c-�9w��^���}C�|�A#�1���߼vS����x�?x�]��|HOG����ݧ�hw�o�v�����ߐ��[Ńþ��y�z<;�yL.��L1>�"$}./L;�]5����:����vQC�!����(��|�O�nNv����m��on�~��I�S��=w��ra���~�ʻ���=^��zv�󿝯G�7�<<��ʓ�#�D��1�{alj�����Z�ʛU�U��[��]��zw�����ï�숃{�Է��Q��ONU�B���|2�Y�/�n7y�w�JC\fI�G�R<��+�pN�+2g�z�y(m�ak�Hֈ��r�����خ5�r�������X<-�n�޾��J����}�ǟ6�_)�0����뷔��]��������}��<;�����O�9?&�N}�݃ÿ'��S���?!�0��޺��Ǵ9��|��e�}"}��O2r���������8����;�}�X=�)�{@?��q��+�}�1���p����>������� �����oN��P���>}�n����ѕ~5;`\��=J���h}���S�A�	7����nC���y�[�ԜN<]���oτ����"���"GќhD!@���z)�>��.�vߝ;Ӵ�g�ݿ�����G�9����n���}��-V>�B<G�H7��{���1;�<���}O)��_T�Î~�ɼ�
��㧟�
�I篯��_nܜ��ww����7��_{yL.��y?���o�zL>#��{��T5�/'��?���>����{��<��o�;ۏq�7�'�'z���Ǆ����xOc�;��<[s�< |IӴ��9�G�i0�'�b({��dǸ��b�H��{F�ؗ�Nf��N��)V��=��4#��C��|���rS
?~�x~���;}����e������x�<���������7�����$ܞ�G����|��d���_�;����i5������O+����pͣ_F�����#�D;�������{/��ÿ!�܇�{������>��;����M�	7�$�@w��P���|q��N!��E�G�D鏢A}�$}����T<>3���º�!+��!B=��������i���;ô����;巷s�����]��o������ߓz?x��q��������?'��C���q� (��?>��y}8*�.�6�*a��w��xp��!��"D~>@s���~��W����Vﱽ!ɇϏ�O�ޕ�ݧw�S�~v�yޓ���o�O�o'�޼�
o�O�����F>�>�����$��!�G�,Ǜ��7��h^~���8|��H"}�]��L/�|�������o�����NL.��{/{C��R�������������e��|�ň�b�G�������G�D�^�����?A�^)�T]E�`|l`T����0[�VXy�r�5���	J�3E&t�?
�眕����cH�f���� 8\����yp�.^�u:)��~�Fs��f_L�Oon����$f_D���wt#�z��͕�����),�_{���=�n�,A��lǒo����@��ϝ�p�ô����SÏ%q����}NNC�ǚ�Q����OGG�=����x�����R}ԭ|�TDW�*�q��_Zj�J�y��K��я�DH��Z���"#��d��"�pB>B3�s#� 3��"}���	��I�Ǥ���i7���;s�yq��}B�o�r�	7�yy�1���1�#�x�J������KuL������q����ǟ���}Nq��9?�{�<+��=}�����󂭿���]�����ܝ������w�����=&O����{C�<�?�ӷ+��x�)���P������ye��b��+�3�h?y��X�|LP� z ��[����X��A��ȟ�c�!Ѫc����o���x˿;J���ɾ����������ߓ�O���=�'&{Old3��!���Å�L8��-��~>{�����˾��q�r���L�S�~�X���'zq䣼[۷&���/<xv���]���	;}{�o������N����~����t�>O�݉?'�>� ����G�C"#��}��K/"o�O<��o�#AX��$��!��B�q����þ��=�r���{|n��~���x;��o(Rw�߮<��)�>��!&�m��߾I��#��?W������t�S�Vf.�L�3J�}���ޱ�<��jb,F��[{O��*�S~w��8��F'{~V=>s�';y�nw��㟮�ׄ®�)�~O�s��V<�����=�w1b= z~>���Ƨ/W�=U����}}OW�*��� +�Ի_�\5����>��~v�w�_���|v�y��=�xM�O�`�U����`�˷'|�|yӵ[~~'�� 9�>���c��|@��rgG�����,��F�}w_4*��7�ߧ������?�x7���]�=x���$���9����~8�C�x1�L����ݷ�Iޝ��o�ܛ�}����p/��$���x���_�����'�jԆU]�f�^C�>���G�#G�p�]&�{���|Nq�į�}�$���r�~q�|�N������7�?!�90�v�s�����~�<+��'~���yL=�=~�)���������x��Y�ߤH���p�1d��yoS��U'[��f1ԤgJ1�uߌ�Wt>���֐ Wжw�x3ۉ��6�^����[:L�(=�Z9�M�[��I�)X�L�4>qIt{SXCBr��d��Q�:����[RuX��6��+uW������\q��W�����oO�~:�P�W�>�&�$X�����<;˴��m�<ߝ;����o	�!~��|���SzwϾ��o�_#_o��>\s��8���]�����!�v�)�£k~T��y� ���	���Â���m��^M��<��'��z�����ra|�Ƿk�os��>�oc�+��׿�P>���������}�����! >�"��A�g;�~�v7�=��(Dh��H����/��;�[{~��e0�Ӵ�P��s��y�c�}�9��]tbw��㿎��o��]�c�	��9�������xO����0��L��<�>t!u_w�@;X��W��!�h��G���m�ռ�roA~����HO߻�o�I;{{��}��.��!���y��t�����rs��y�r��S�ry��M��bw�������|Nv�S�ـ�jV@���Ȫ���zG�Ds�ߝ��/���=�;Ͽ�ސ�~Q��TF���""5��,z��)�=�c�a_v�~��yM�	7�/��o	�ޓJԇoΓ�קo	���0��a����앓��fj�Ͻ�����Szw�=<���c�|�������9�����ÿ8�����߯P��U����ǁC�{C���}��ɏ.��M�����c�zL.���?ѽ��Fb@��2c�"$|S�X��bF���qϯ�>}���~㝹]��єi'�<V�|;��M�޼��/��p)��p}B~�rw�=|�yw�j��{����&~v�x�~|9w�i_��<���`�{O�}��/z���ztQ�H��&�۸�r�u,qB�1#�0��`�P�"$o���+������pxL?`�Q'�n@��������ϫ{v�?��}Cˡ�Œ"/&��fE���_ OɌ�;�����kH���~H��ܻqB%�3��
�e��QZ��8����U�D�*ۄs���DnE���xW_��ŏ�U6�uk�:H�9�\�:r��d�75�~������G��bBz�4=�����
��W暋ݞ�#�o�x5�z0���\�[�+^�)v�͓)j-4u�c%[���\.��)��8	��{��̜Ogt��7���0�aQ�r��Q{��z�?G���ˏH68��c�~���7��\�Ԥ �h���۸yU=1�V��f-Ҧ7"&�GX6LLG	:JD����2�h���������>��u,�{*�jf��B�o�s���|�վ�@	Eh6���[n�Xx�9Z���<���3��}jg���$tXq��Gc����S�_�H���L��Vߣ�JmL�T�4����� �ZH���a��놌���:�C*�RБO�e��M����~|���,�b��TT'I���q�1��)�]���ll(����i����O����jpJ�r!A�F�vH�����u�G�K���J}�m5ýcwL�j�R\&�y/�� U��)��w��1}�a0T
�#����#{a���u����7�߮!�R+�'�4nt7�Cc�Y����$0�c�,�i\�G��;p�!c�J��}l^x�zk]���BN��>�9=x��󬢊���p�5Նl���g��T-T�T`��p[�\L\n��h`b���FB�HBѺ��z�e�^�� sq���N���юwS�&�L�
�(T��uf����1��7	�m�JQ�#Y�s�C�/jʘ�a�_t2�+7%X��<��q��B�j��d�ti�,�7]���ԕ|tq�#Zin<���s���o��TI}��f o���U�5�}=;_�?}4�'�+:!9�����\��i�'����u�{q�00]-J�5*'���py+�G��`|1�PW�~ʹ�U%�e�%�uPʌ���6��wķ�]��PgqG7K@@݋�F+�l��>Ū{���RևW���<O�]%�YZ�XT:����L�(�������וK��eP
�a�PԦ_k��
�1�n����nN
D��NX���;�ro[����ep�T��s�!k�,X/�`2��'-��v��pb�����[V��~��|��Z�*h�RA@�. !
��u�5�%�SF�lz��!�X���NަE_�k�޿y�5eR��a���P��\�d�B�%]�����o8H(�a8<���j�%U��o:�U�k�a�c����B�rQ��|
 T�I�G2�����=�n��#G��H�Q�u���WO��:4�f ��	�2T�q1�)V���3P:ޛ	�S�5�>�7��x�>5�N�!��Ճ�� |�QU&x�k��ŀvuw��y���^�۞���{�˽�
R�$9oY�����%�3��%��ޤ	u&T����kѦ�7������]6yk�y�B3��V��_�5Ŧk]�t�]��ż�eJ�������[};����q��;������}مc��ϝ]]��n�-�´�t�tq1{�]n��s���/`�I:Lfr��{��]X�g��}E*{QX<k����ػM������;4n!���]
cV��ިyrQ��l�5�.0�pf*quƌ�T�'�����_KU'�7��ղ����
i?�o�"K�o/6>Y�hX��V�n���s�
���`��錸4� ��:�tL{�pU���1xX:i����D`D�
ʈ;�
�k-�7��z��3ոR��">��t�;���9����/T�s��G;�9wX5�"��l��*�c�����Mh�{|�qU�l�L�%�#b-5l��Y8(b:��n���F,^H:�:P��|{�8��s(e	�umR�� Ҡ��,%�a���)�C�l�A�1��,�Q�1�ź��|�-0��:k�8C��.��B$� ꐏ`sC��^�r�Hݠ�=P���gz��j�͔����s�R�F����>���-j'��� ��k$J�{+Z�ܣ�u�</���5=�0�ë���ʙ�����:[�A��	騸�<"S�U�ӂ�;o��UP2`|�ÐX�+��6����C���.Ge9�Vm+Tx��<0wR���B�f�<-���7
���[�J
�ӕ�=�C��BFm��"B-�W?}U�����cq�U���p�c1�9;��sS����ci� �3��%ޣ��C�����oۘ:r��������>a�w�����z26����,����IAĪ�z�c[��N�@tH��s*�Ս㔚��X�=�1�r�#j۲3�q[�*ɚ�#���klJ��y���2�v��JU��(Gx!�qt�މN�1�ޔ�f,jn��鶤S�=� ����Yh7��1Y��d���:��DĞ}4/�֪�
Xv_g.�uz���Cŷ�ܭ�nc��&*hԷ�^h�%S��N���]��il\>�upr�Nޱ��E�س%� �f��=�H��1��XL����BЇ������+��3ՄT��/L��
eX|����v����r����ƏY�(�Ltݤab,���{�.�0:2���p�U{���S̴v9Lm���\�y.w�ߌǡ_�|��Z#�b�&܁���t�d�5ۊ9���8>��{�v0��x5�~u3+�K��<zy�;���*���&�kz��!�X��s�<�S�﫩]MA��Qi�A,��X�7d2��ْ̕�Z(f�&�Bnu�P,�X�k�
�{�|5].T�8/��v=�XϺ֚n+�x�Zv�t�
��ٱ���YP�4��uxĝ�w��vN��)'���/�{������:M*�@�ф��1��"��ϮON�u 7�a:uC�h�%tH��[��HI�������V���h_AWm��/*��%�̭�7~��0&"Ӵ̎%	�ˌ�5b�Ao���^?_f8;���	�Z�ۈm�=ύ��]��"��*?xFTP�n�gP����;Ċ����w,G)u�����z{n�eIӾ�̂���AJOV`{�9�s��]���xH:q��]]=84C.#�f.*cr&�G\d��@��:��vu�nS�ʺ`�m�;�!F=�Bir��#��_��6�T ��7�ͮ��GS==+��=]B�^��y��)\b��r)�����ﯸ�O!�!MM�.�V�5�.<��!ׅI�Q�@��!i#I�<#�;�ڿtl��.xm`3��vG��O&fa��[ ��h j����C�t΂�iR�q��A생oBn�b�P8x��]��t��hg�t��;� �V�&�!A�F�,��o�-5oY�F�bԭr�e�Y7�J[KG^��N�����g4>C
�dފ��B�2��r��ٌ��W�;a¤*U��ݳV`/�*�˫���3zq�I���k��}&=�����U�ܤOt�W],��<�� �/�Ѻ<Z%J��fӼ��t��hU�QZf��{ޏo_2�Z]��k��~CZ3�T94���C4�-|����t�}0L�`��ʸ�s6�	��o�����Hu��z���惮�<K-�[ʠ�Y&^fML�m�]���[}&�#��c�ڹf��և������
ޚ�k��X��F2O���u@�	ۑ���Gr��ƪ{�F).Xg
�5�aViW��9�j�W]jc���}�r��3%N#�okx����Bu��eY��g_h�n��g�ʰب�5�rՎU�˻�-��5*���:g���W�Ӭ�Bu��3#0���b�ԋ���Q��Ϟs;wɻ��Z2���Md�]���H�Ŵ�HTa�Y��K櫄_��tT^�I��/&V�vT��<�j��ԿG����.H�fUHn:@a��jS/�_�A��1��f��ó�^dRH
���MIZ��ͫ�a��S����DE-u�~���]��岲!ۿn�*R�<�V�yT��J�gb^Zd!̢A�x�mW]3�}�Q��1@�tǻ�����4.������X�-����).�1�i��o�4��ʾ࢖��km�~�M��~�d���<���]A|��j�MK��(g��nևQX]���ܔ�k��o�׆����@��]��p)v2�h� .�=x��k��7��j�&v��:�6��Y%`[��ѯ����Wd�!���۴uH"�-D�5�f:v��0��d�i�7�ϭ͌�"wj/��v�kr�JWdsw5|$�u����-��36�M��C��Ŗ���2�]V����0M����fb��v`�5R�&�B��M_cs��=ub��T�y�9ԡ�Z�u��IY���F��R�v��H�}��|��vfV�;�;��в��o��R��z�(W)�~P��ws�ݧ�5�nN�f�2�A*��+�28X�Aۻ�+P
�^gOn�E��a�f��۷�|����đ��ˠo� �X�
<m�+6�-q�(gf.�m
/v�	8��ֲ�X{�ӗTR���F2��ͷ1�@#n1�2*$�YՈ����]h���m�]QR��G��dj�2�����8f�F�en�okiO�6����E�Z$M���t���=
}�WQ7��=s�*��]:����a�Yd�i��HgV�Z,4h+gj휠�w��d;�� �K�D�T)tnR9&|E�%�Ay���}ZN�{_j��"WY}��:s:Zx��QoQQ��d��)��ݛl� �G^�H��M�0�J��iҸY����9AȹHO8��*�v���iG�!wEY�0��Xr���f���%訮�Z�/��%D9�뭿i�v�{Բ 5�Ȟٱ�\i>ua���+e�|�#d?�[ì4I�����ۡе1_VU���e&��	0�����A�4�"�'S:�v�M�y+Vuqw,�]���㵨-���k�#z�⳺�8�9M���h^�אҋ#1,�:��nu�wzͻ�&�68�6��&gR��M�wi�]S�̖���Y�{m��0�6�m����1y����5Ⱥ��jt��p����[���u$���-���
�q�c9��Pa8ܡ�[�Ρwԝ1z�V���"��lYz�	���&�+ӭQcg-��֊3	�<R\p��w78��d����MJU�pa]v�
 �A�/m����z&H�ds��Ǚ�R�4�����s��9�S���>���I����s(R"�7z�����<{���2cU�䜀y���x�e�Ĳ�7�r�e/�����f�&�2��s��S���7�WV7��T\�ID���:�Y���r![)] ��e��qt�������5뒽of����8��Ex����9:J�n��d�X��T�0���9Ǵ!	�N)�i`��*�Sr��h\�x��%]t�jU�$���iQ�0ͱ���\�""��Ss	�j6���6�zp�t���'uN�-k���o�|8�|�8y�
)@�ͅi��RDiz�:眴KQ(%K��K1wnxR�YV�R*�����H�*B:Ujj·"͈X�kLم֮�/%B��fHs�<-AV�
�+5,�D���e��)3P��e�AC��=�KLT��ˢF�ub�˥�B���M+TtvyԌSMSU�Du�<*WWURC�(r(�!%RJ�$�B�E)�s��.$�9^U�b�zB�����Q-	"9�jbj	)�ID[ �(�H��в�GE��T�EV�S�W(tA3-D�J��52�%��,�hi�Ufeв��H� ��JT�
�j���b��G0�U-K22�V�Er$1+0�R�ĵ�)R��'��]H��"��RR�u�Z�"�a9h��$:a��A溸���*�1@��[��ER���ZZk�z�i�Ŕ�r��J��D���
|P�E
5oyml#�7a<���Y�`�3Yd��b\ٮ��q,-�2+&t���+s�7�k3fU��+��Hn��gg=��U�}����P'G��j�j�W�p��1#�I�2���̋����*�/�����m�ڳf�wz7�wE�\�k"�t9�*U
��F����@	�J���G2���Eb��O��井yH�U�ܷq�˺|u9Ѥ�s e:�&�L�.8R���4olr�]�:�_g�)�n�.�En��o�\k��N�8\���w6�U�W�؃1�$�=n��t
��h�����P���& #4���T�:7`t�n4�1�˭ѸNc�1p\�%�*�9MV-���7���fC�08���w��x��4��l]����l�1�杚=@9u(Ƀ�h�m-�Uwb`z�u�K�x������Y�Ҿ�7��+��^'�aV7�1�[-�E_G>�gs�Z��9A�q��Cr�1��u������UҎ��+�*��!��zK�a^�U��=.;u���1��Ü��]k� ��wR#&����B[S>�q^��t�|�^4������[7���@!�N|�Q��������
�x0����I�N�}}���\�^[�x�#Q<\n���+"�Be�n�'U�Y�+�JX}���<wv��`�r��`����)
�ɮ�m)�p�X��u�"\��]q��Z0��Yjf�GL;4Ґ��ٍ@�:=��)S ���59m������a�9�AZC��d�D��3��ܪ�=��B{��?�ۃW�=ܻ�!��+i>*�qy�Ԡ�~��À�zϺ��Yё��#fXW�a��S,	^;��M�v'ݴl{5VF-�r=�#��F*0�8|�>؃(]:P�
��Tꠊ�.�,��^F��֊.3m]v�H8���Ͼ�V�}��"��Q��U�n?,�����߉P�{`�Uܦ��ܶf���y^�|&��@-N��86(�=�UA�A�ĝ��<�!���䟯��|�~Zo���qE�����r��t�~��Fڪ�����_�w�lz
�*ϥe��l�k�lu�L!a�x��q�M\M�e��p\���#j۲2�摔_=�-L�]닷�є�2˒.S�
��L��5���d�m��&��s��`���Hj�ө�*�Җ�\�]3�C�)H��6H�<�h_Z�cr<��>�q�\�OB����pO=n��/D�Xt����2����� ����A*��
p�j�����a��_��_+�[�r��i�rn�;��)��w�:I[���a��Fdc�o�B� ��<�2Σ���[a���go��`$ζ�%:���!(��ט��d�7�g��	�[��Y�T���=�e�>��ۛl���J�}P����D{��z&��uZR��vH��ö���S%烖���8���;�ȕՂ����:s�-�4��ImF��Ek{l6����Sr���Պτ���?v��Q���naw<��r���؊��窦�͎�vX�{:�\�`s���� ��J��<���p]�O8�_��X+G��ܮ%C�ƙ�0�o'�h��3J�W2��A����Yљs�/��H���Ɍ��0��������ψ���ΤF�Yg�:�"�Y�ܺVc�餈9E?s��ռb��+E�0�0��:+��NT����x�ߘs�=:p������x���q��d���#��Um�z�hT���^P:+��$Z�%�p�Q�.�ï��,8��z�{d�����w,G:���h�_� ���[@�Ħ��� �׎�c:���a�Whױ+�Y��Ӑ4C.1�6b�*crn�u�6O�C�û���iAjږ��y��0;j:㮘�1�fD�����!���eDZۇz�^ͣٶ{(^�5���**�6J�wѓB�U�}���Mq�:�1ZtUbէZ�������+�xn�)rٽ�mgq��x�D�J�ީ�&J���u*��4����;ӛG�[T���ѹ���*�'C��@v�%��3���}Ҟ�qW���������U�W�U|n��Χ��,7�B��#�39�R>�UZ�Su�E���=v��8�-�S��W#8k�OU�S�,{+�c�s�4x�D	25�H�g�d�r�E���V�54z���7<�Z]S;��)�&Ҩ8_��� #�	T	�`���;� ��'u�B�����Oݷ`�mZ�DńMCS�TCf�*]z���.�-g.Ѧ�-V�X�WEù�z��0�Z5�Óɺ�^C4�-UR�5(�gw;�`����UG���δ;>:�Ts^�{�3��q����pڨ�K'�4m�@s�{v3ˏ�%:��R�=�j��4�t}/o��Z�����PW�6�����&ȇ��'�F�%�UU�\�ø:��Z8P=�^3YVtP�-WK
�sJ���r�&.7e{401X����	i�V\z�&�o��6�!\�gDeX�^�8M! H�ϽW�*un�y@KV���Z�)D��;��:�ڎq��<j��p���}�]��s�r�pw���]�J��lg�J�pu8����Z*2x,)���!A��T�^fm�(V-=�s��m �M�œ��ፌ�R�'��:��sً7�
��@k-�2�	ar_sK�q庸�`�p�-�o�ќ�ku(Լ5*�Fރ�X�/�W�U}�,�H�e���Nq(����O$g��6M�9�-�櫄u��bB%��\9§����R�Y�Q�
�������  d�<��/�+/�nߝGE�^� �ƕFs{�C���~3 ��gC���S�H�����4�`ۘ�7�岽#�.��w&j������V�$�Eߓ��0��(�S��@@bԣ~/m<�S�[޿
� ����#t8���;+����� ��j���|��Ę�+�T�H]TJ����n��W��bP�}�cP�D��ү,hb��,��k"�s��p�*U
(�pzH�wyBM@i��f��cd{��ݮ�U�1�����8YwO�M�+�7�:�H���}���I��˵�9V�ޠ����F"��0�1�9�J�u�<˰�������L����EV�H����@j������4�W��3zx������'1�����.��آg`mVaf�6ܥ�8S[3!ᙎq�`�H��i�ޕ��:���(5Qט�W��|�g���3b�U(x4f����}U'G�Z`�����o.q��Bl'��T���Ө)�߬*3+n�v0��wJlՈ�D3N̉tj�ƺ^����Ҁ�sn�[����[F'��8<&s+9]�v��,��Dz=�d�e�Oz�Qg��ʫe�4��LL�_k�}f��\h��OM玆5�)�ՙrf�ho*�����]�A��y�`�=x��<O��*�an���`��8��y�NUf	�����2�X�uLB�!���b���~�u"*0�r�gCF!]WpL����A?ov>u~O.C�jcD`��L�n�[z�o�ך7��\~��]���ڙ*LS�;㝷[IB�+�j�v;��N��� 1�T�T��U\�'<(b:��h=�Td��m�R��.߾���GY����X���TF�;:2*Nl�
��1�e�E�eٺ�&���&_a�7?M�+�l�����u�gJ$�:�"�4����o�#A�+"�o<N��7>�^�LE�r��u���1P�*Q�0l����Y�w^�&��ɠ�X�M��� ���ܻ�ȧzZ�t�N��ܵ�]FUy��j,�'�A�Np�]�z��4�u�����,���*xy��e����#*�(Og-���dѬ�����b����楚��)Ր*%�Pۛ�J��c�� =�ȗۛ�ƅ,oIË�=Hb;F�謓*%qb}�T{7:�b���a�
�"��W@�;{s��,_Tb�;ؒr�-�>7��k��\kO���XU����a`�T�_}��}_8J�#��JWc.~��`��^��x����M\M̱�C0�a��ڋn�͹�83|�]�f�����_L�"aA�K�&"R�2���+W�N�1�ޔ�n���	x�S�sաEY��:�dR�)M����ᨄ��L_��׆�^��~�A�(4��yG��n�;�h~<ݖ@�D����?r�u�MOQ�h�F]��&*��Ɂ:w7%�v2�qᏻ�B�����S%�r�ב^�S�"8"w M�����4U�0ޱ7Dkʺ��75��\�;�GF���y�WF�c !^nX^ymX�g�c����%��i=Ւ7K����-��zZ-�S+ۓb;���ޅ΀t�#M�mC��ŋ���5�쓓j��_)�p)�z�o���X#�^�@ ���Z0���=(g���Vm<���בhI��kkz
S|_���iD�Q��d�S3�|�u�O��5Z�z���g����q<9F��-��]^�m���b��ۈ�
1�\�C�LOJ<��V��>[t�$�a9�[�蹪ηټd�ԃu}\;1:��2�ɬ�@{X����m��hb��dؕ�ێ�xr��j���*W8�4Dz3�o����K�%.ɒҢ�!j��wV��
���<�+G�:�5:�f�f�3Wkrk�i��}U_}��B5*{�;�w��h����׉��ß66,�/Y�� �g���ԫNa��X}�5�N�C��]���P�8�����%6���~����r�?�M��3ĝ"���EC�.�vz��k>��8�j2�5�]��.������pه*XΉ��a�E[�/@��̧=� {�V�+�D�J�����P�;�f�6hMD.V��s��㑧�j�`,��6V���e4�ޣع��J08&���F��@b`����f�4�G׊�Y��ǽ��J�7�?7��8�c�ϔ�lzL�����W
���@	6��Wi"�)�}s�f7����bN�zRG�_�ĕ�ý�7��o�:n K>�F=@����iR�q���|@�<���ҧ��Z�:�z����T���"b���W�`���5¼���ӹD������}O�"l��)��%~b��Q��C�P���,��UR�#�S���Q��E��Tȟ�i�X�Ch<�[צ�*@�6"��#����^���4�n��Lk�q�k)�X����M�0�k�+{�XC�V�S��EtMD��	vsqn8(�q�����j&�^�ZAُDYۗ�n��9�_�/m&D�	�u`Ń �hFNi9cw��[VU����8��< ���Fk�p�u�G�9G,q���}_}W��	�y�W#�3IF4�,F�1aTjև�g�m_�5�ƧI�`�7�nJ|MҦ�k�7�O4��0OOn�F���C�V�4��].��үa�t�8Mn�{���cz���D��W=(p��uw:u;�]G�?^�eY���Aֈ����a�IW���M!�kJ�^�݇{�{ϣP�S�W��0�#,�3��3̌��K>ʣ�d�� 	S��9z���՚Y�l�-��9yP��L�"VD���y#<�a�n<�ضo��q�:*/g$�.�紡���E�n��<�@�pQ;e��Q�j��h�r(%�O2�z���ﰈ���^�9��%
4:srtS$��XugBڙu1�\����ˣK�Ø�'/�b������0���p��e���;WA��X�2]���Z�'��u͜�Q�FƣȄ�pg�,��<hs����6:�̂�Gi5p� ����b�U�1��*�<���U�p\������X^�G Թ�Y�c9ܴaF�u��l�SO��|��/�PI��7˅�(
��j{�$g�<nVcG~���
�'�^E�'�^n*��������B�8!-��R��r+��$q� �nڔ�7h�W�Bm�Ol�0�v^vϴ���|��S���R�E=�e@�WSۧ���=�2���>%�(;��UU��Og|�x���~�#�Y�{�F'�q-�p�.���N�q8�zꐚ�*v�lF�e�oyҾQ``�8x%<ƙ\V�	��\k���G ������������9ۚ4���E!�̓hߍJf��<"��qѱ�2��1�˭�L�c$���8�͞�Mo���`74�dR04���~X
0Č�i���F�R�����E�d�z9�j&n�f�f+=9�|�&&J����Y��F-����n���1���g+��.X�l�h|��E��[,�lz}��A��O��*3W���X��V)$=�bJ��g���}�Ƌ����9�#���<����Yy�G.�U*�B]F�Ż�9�p�,�P�&��"Lh��)���ax�L�'^h�{��z�A�T�������F�4�To���� *6&;��ihts;�@�nUg�z/]��=��i㎐,>����������������.�_GZ߬����r�=rV��]
��&i^�g@M�zHI��_��|��Qk�1Ա���HR�jᎍ�`t���i�چ]rÑ�VF�J�Wf������1֧���q��n*ٻ[)P!�Wy��yζ,;tΙKy�Ël�2�-7����kZs�)�����봘9}NLyz�#3Q�"XZ��!�D&�q��`�wOq������J�U��Z�ї�n8z��k*X���ɍ龹���$�7u��-�\I�Y�۾��Y���i4�����5o�N�Cԩd\��+i�_�^Ӏ(�1���5��]J����Ze�x��s�k6����[���Y�>�phz�7z�;�2���j�oBm��d��"nl�,�aq��L�[���*�na��Wd�F�`9Xi�.R�۾ic���Vs�$�bV��N��Ý����g�r�rAth�u�9�2>�H��`;8b%�̽�v�!�ԠY��7wEK����*�|fjJ�G�'e.�D,rwW�h�tD��7p.���{��{i׬�h\�rn9"�-S���ϗ:Iaʅn�K^7B�[���b�h��hT@�Y����LX�r�K4�f1o�ujj�K�0>3ڳt���yy�N���Y+J�uՠ>�,��C��e9��|��:G�c�.�s-[�w�	RxR��3�Y��Do�hr��s����Ttp��V�<P4��$E�Qv�G,�M���o� fh�ʃ}+�y�����]�JS^l}�Ɇ`����Y�Q������O�	��y�섖��j*�9�70ǽ��\&J�v�R�w4jj �ٍ�*O�Ƶ&̾b����ެY�m%vb
��hE���ٕ��K2�e�lr)����Ɔ�'f��fr��(�\T	w��ȌuǨ�+��:�Pƶ�gY��n�'���_"��,Q��C�2A�ڢ:���8���m)u���2ؓ�^�X�&�"��2v0|9;�,⣐u��o�oiϒR���B���?Ml=�R�<n��f���7t��'t�j_=�-�4kr[���:���M��q�k-�)�۔@����������]R��-��1Hx�m#���6K�'m�NU�k..V���L�v��q,Vd�1���sg�R�դx�'<4�� &�(&��r�}�|i�$�)Q��hs�Wd�j�d4�[��Te�W��DK��n=�bTe�1ZљNY�-Y)�\�0���8�+cJ�hu�h>�{�:����k�hKre�+"-��ӽ7��S�qޮ��:��U�ŵ���!&���X�b|�EK�ʵ���/�y�T�T��͝L��F��p���ݞ�\�t{.8֮��/�H��'q�����w�����RH�pN%�Æ�"�r1�I���ė
Bq��K+%-�]�����4�o�)3�[��#���!}�%�Tͣ�06�}V�	U���V��W�zM���E�
! H�E��ɤs�3�ܩD�ʐ�,)H�W"T��븕�[�9�\#F��wH�*��,�J�(��BT�DV	ӗ��.Uz�U!K%#9�h��(BR���Y!w=Ҩ��P��["�Ґ�#���T���!��W(΁TAE*QQ��U��Ԑ�WIL#(�@��օ̬�Wdr(�&�ٔ�J�UZ�s4��A��aҲ�l��IB�DtR��(��L�S5�2�U4VEr��E(��+i֒�kLΡ)*��DFT��Ar�2��L�hP&��1��	.H�%A�͉e�P��#*J9elJ1a*���\"
U�K�F�kH��r
��%,����G"죝#J��ZY)Es�a��\BL�%"9�J�QL(��f�	P�gP�P(���B" Ԋ����>ۿ�������;�	C]����k�G>Y�`�l��M��8֎��ċd�Xܔ:�Q�r�(9��v�ɰ菬v�ꪪ��qӄ��y�����vx>��RG��mp�p�\+��\-�+O�
t������HGP����A>X�mX�z���L�vT�Z��q��2�3`�303����Ֆ��x|;G��2JI6w��q�؅����	�3���;��q�6��� wLx�L�%��[,�W\O����ڗ�tj��̇��)v\s��m�:i�}Dm�Uy]<�5Ձ��X��(�M� .�e�1!"�1U��)��S,w�1�S F��ۆ/�]T��PWom5���	ÚFY ���8�D�"})W�{L�P�o�]\;"S��Fߙ��gޥ�}^�`�8��5�	���������P|��VZ���A�1��C�Ψ;��w�v��m�jw9���-�dՖp��Js��*�
��N�	����I��ӻ{ym��ю]s�%��
�Z�X}S�橒����z�f��(���d-/UIu�7)��'m���{s+��El���ݸb+S�c"Utn2ܰ4�[V!��P�W��_�:�t�qu k���蛖�+7�H��Rm��)�
9�x��6���]��J�z�Ʊ�X	�Y�QAj�Y/0>�ZɄ�PC������$̵�K��@qμ���ym'�\Z�Y�v���l��Zv<x�e�(����T�q��ok]��_}��TF�Y�������T;��Z���*�ʴn*N�z}��>Z�0v�}�%�c;IĪW=i�P��ٜj�K�vD/��g�.[�L9"���Ӓ�i�Z�Oˇ���s�y�obzy*��
VۀR���A\���ʰu�_S�,dd���2�4���M^��=0�{��⯹�q�~��sB�*�2���%��҅z�X���Ϥ<]�kV���&-�L��V��_�SgUO�
���r�M�,�Z��u�3b����x'V����5\��:��-�*Jn{bS�]pcrr�=�R3�=:��E^V�=��Yd�H�A���֫���J�/
��Y~�pً�J�݌�S;F�7{g�k:��:)�d��,v�e>���_]!^)��x6hMjV�w��~c��"�[I\FF�mE�X����\!pM"��x� u�Ze#�UZ�E7^)�ĵ������Ӎ�s�E���h�s����,{�+�4x�D	2#]��Z��-���Ab$��]80�]�jc{ǯ[V�ioLH�҇���#�]r��a��XIl�Y�D�������P�$��3t�t6K͢�m��H�e��ɮ���կ�E�Q�NJ��@�b����x����~� 2pR�c-ͬ�{ޏDGVc��K�H�>��CFD���졩��=��0Y�D#�@ %I��˩�.��,s�΄y�T\+��ہTj�W`��MZ[�LXb�&���*��=�r�Z�arԌ�ۅ�� ��Q�)������j6�*�&���癦 �h��q�T�q������ۈ�TP��7��_#��;�j����V�O+�ͪ��y�DҷSkٺ5
|OS�}���ܞh��(�3�H���'p��W[�C�Z�.�e�x,�3o��{��?%>r{�8���=�a���B�t��?��a��(MC�����m�Q���I�s.z�m��59�et�V��5�Þư��s6���m���Z�s2pg�(�����T�d�@�� �n:�-gQ�N����;i��G�rɧ���E�ܲ/3��j�hLe�z��F���L�@`
O��~W0�6�ضn9���:��0_Jg��4�:�>]��L:,�0�d���Wtg�CG�] �e���+Uאۈ�bkPVRZ����z�� fv���p{Ա��t�Y��m�z�����W9��Op��A�&�b�cx�N�V��ȫ��'�嬇7�R�[w�V3�*���k�bir.���(��.+�:�[��˓<ڜ�J��K�n�,fj���g+��}U��U�[%3'��&1}�M�ܜnI0~:�6�L\Er�"��ו�t���S���l��K	?,u`ko'����!�+�ƙ��ؗu~�����>�9ۺi4�n\�1k��q`�������̂�Gk��]zaW���@��Ę�P2y *�����~��v�鴨�����B��i�u����y��h6\qԿ��2�ꉇyꂺ)��^�����e���*�KyW�Tb}q7��.����uÉ��0W�R�(d���ܭ�Jm�8y�u�/�A�V�ǺU�ɕ�>�N�8\���AyX#Y�Ը�Y�N(��>�M�<I<����& #�)�k�ѻT"��	�N��j�nH��`a��z�Z�>�˧v��w���>I�W�R���<k���
)�B�w�{n��YXG &���5�Z4�wz�>��O��W���OP���@.�W�\h�NJ�z ��8��v��g��W~B�wt-��������ζ�b�|�*鳚hul���9�:5-�	MKj2&�t��4;�*��efq�W��K��+���è�tBH�6��K�D���Ԥ8k��h^>��0�3��A�R��Q=�b���Z�a�����b7ֹ���Kv�j[qF���k1��r�q+%��;^K�Ν�㹕������c9y�m�����qp��?C/����Z�3]�Ń��"��H�s|���h�]l�����a27f;���9cD`�)�������g�:�F���).����(p������}�0E���K�>8�V]��T�|J8vb-5L3��K�ofe��E�����),����:oK�^�X'��x�a/��[��r��ٖi��Ό���7��J��~ܗŃ����\cv�Vq��`��7�2Yګ��W�=t|9D���U�v��|�H��z�<���S����������1�9��Rw[O��������cb�r��c;l5uN�С岕؅����	�2��n�=7S����:��͸/-)J2�:�Ϡ�àTm�Ef��,ߨ�>�)SÞ�!�یt. ~�=���{&S|��G�����d�� �N���*𧦻�g&2T�Ws,w�1�N7AC���6J1ۚޫ&�YniD�"�����.��zWx���C3��	]7W=yYN������h��h��=�M�{��$���;eB��VQS��?j�`}Aun��.���Ty�H��$mi1eK�)f�Fv��T���*(��r��u� U�����H����P��j��Za�n֍9�RS���s9B��¢�a���z#��VٝM�f�a������1�*!7Pr�S2*�JoƧ�Ƣ��D�|��'�KݹL{�f�.���)���s�a�mYg<LZ%\:��� ��u���2��h�N�����Q����)�Rz�i�z��~֮C��}Q�2^,s���<Q:t�J�f������ʝi�f�oњ*��ۄ#S�c��WF�c !M�KX�l��g�1����o	���>tۥ��~(��:���8+�U.�t�9�X��w����0����d<$���-��ZC��%�F��F�	c�ꊱ��L�`1�7���F��b�g��\Ns.���I��"��h3��C`�a�L�*_��x�*$�>���������蒯Ci_@8K^B��1W泎���$YO��֞�\|P����|�.�o�\��Y��K��a��Ӵ̌�i߅êl�+�n�F�k1�pwf�����+�[[�S%���-�b��V���.�z�1�"�Jn{|�~�\ܜ��3ol��U/de0�l���N+����Cv���&EA[J�EӞs�A�ΏQ�/"xz���yH�g|Dշux���N�kR�Ԁ��mh��Lh[5���6�����jj��i>z�ۻ]�%�R�kazQxK7��1�(��I�#������%������D���E�$�Q%3PeW�ѵ0䫃�AF�+�Y���!�v�1T�]]�]bg[�p�)��h����pV�łN�L�&�}t�1x�5�BkR���s������a��o�ś����mZ�,�E\@6�  6�?(d���t�^���K��P���&}7})#�����N/~�A����W
�D�D	�̅H�i!T�VM*.�R������[ͮu\4d���졹	�q8�A��%�L#�S}��L�b��M^�Zm]��mq�y�=L�;���҇��s�eʂ�"b�1a^jp
V�%L�*��zœ�YN���{�U��P?8_�"jTs�r��į�V�j6Ҩrkɺ�^C4�+o$X��"�Ji����iG :�Ex����,�����骞:��"�O�y�{�k. |���d��Ś�zs���,�w���v5d�Uq��qp������V�>8�>�����3 j���T�kU�ܣj��}>rz��&Ư�Y��a}���HT�W�����A`1�Ԇ0_�mAڧw{�Zc�]����S���cy�������һ)��d�\�c�����ȴ`' �߶9�����
+.k��S+��n�gj�8�o�r�|�$Y�6������,��{H���r��GWU���{�f�z_������fuR���\L}䧂�"�Οd.j
�[���X�0籬:8��~�ZA��L�e��/=�{�V����/_ 2��
9�Zu����#v}1n�E��_2
�m�j�欜�[�ў:]�.&e�VI1i��1\�dߜ���C�Z����i�/�t�����U�b4�gIᖗ���Թ~�f�qU4t�q,�k��_*F��2ϕ�Ȝ�\ik���<�n��{7'Ź V|_��mŨ����E����[a����d�*\-В����d���ߓ���v��f+L�q��E) �x���[��k�7S���OϬN�	�GZ��f(歏_�ä3 ���C�3l��$�������`�W-��s���΢��5~�tKzh���9�]���|mY�]A�DJ��[O|��*�{��BZ+Kk0-��'Ƽ[��ny=�V��3�2+CĖ�Qj�OsWZ��/H������s�z���M(o}�/j�77[ ��b	2��l��uq���i�Ǧ׽��%���dJ�$4�W���ap�t���J I��q�P�B�^��b����I�Ns�HS���/
n�;9oV��w���l�\;Y:�<�Sp��Q��l�,�DīG��s��}��U�XF���sz�*Fm�¤g��P%(�pS��]��9<|n�gnGb�.bT3M�]ft����;a�+�Q5��@<�\��jmvӥR��j��ub��Z��.��������bjq�Tf�"y�kj����� T�t��͎.T��|��u�k�W������lmu��b�&1����O��m��oяK���H~_}<��Gs���c�^��z��t^1ƺ��q���-Γ��9��5������눕�*;S���x�'��w'te�:�v$��kkB������;�Gַ�7Yq{����}i�����]�kh$��~O���~�?�YG�v�_v�s �Vӭ�	P�M��l�Wk2��#qe��}�9^ӓ޳�����?T/
#�e����g��W��J͔3]9]^��!�S����\�z���x�M��|�ͬ��{[.���EbW����{�.�ן_Fo�/!��H��Tۚ��#x��a�*�J�i.f��]V���y/n>�7�B�&s͘�����å@I��#x�I�[Z)��a����VV;�cVΠ;�	�������v��jE,���P?{��Dz��K[����Q�;=u�JT�8��CYq��i��:
�BB�Hv�w��j�h+�r��I_�Puޚ)<��m�-���\\����oQ�ֵp���1Aw�����$�3��'���mӥ��[�%gy�����b^��z��o��2�
{���▊�Қ̀����[�ʜ𻣆^0�(��;7�w�d�)62���tts��OE��x�]{3K[[:9��p9*�|s�5hL;A_��(�!�3��U����-�*Җ�������7��{Z.��T�4ø�;���-s�.��|zŰshu�[�~�Ķ�7V�jz�U4��n5񩛨��P��}f'mF��{�B/ȋϜ��|����o�
?)I�j�,���44^n;�I�����=�}�LL�S��Êh����Vc���}�;IO/��{�n,�RM]������'���h���ݭ{z,�+�7r�((K�՜��]�"�g3WTo�iE� f��X��iU����L����l3�֐�c�P��,�s^أ�VV��� \�r*8�oS�H.�
l��b�W8�~�#��T�ĩ�����{�,�wA����N.mૻu�l�Cr����Yy��̫�&"���w�=eH;�!�,�;r��n<oZ+v�Sk��5Q!�WF��u��̥t�z��y�����a�n� �ZUe���9o���t�BM��qǣj�a�4l��[nL9������-}ڦ�0([��)zE��%AX�
l�l�{p��@U�#5��3�v�7b�"&\�AN�o�<�����ݫ-�+J�č�"���r�T��X	��oz��X����@n�\=XD�X�W2��D�ɕ�Rst���J�j۫wFm����
�3�|H�D�XJ��wq�s1�h%.��+��eeb\z�^C�u�]�����F.M����rb�EU�d�
�ʬS����ο��6��>��|���*\:�m���hu�:Q�6���V=�K�EZ[쀁b
�ޡ��'Y���^-�߈`$���Ȝ�#��X�*�nȤB�QG o#sZͺ��oe��)eX(�=K�g�d��5Q��b�m<WR�n)��St�o�x�.�q�b7��.�4�#۽יNKw'3�>uҷ�k4�
�R5��zk��r�8���*�`871굔�V<4���h�v��׸$�b-H���AY ��;����Gr�)-w��0�,w�%.�,U��
5--�$mtnkK��A}��R�qCwF�r�ۘ�]5t1,Sw4M�vc��
���{0�e���I�e\̻\��S����-�WO6G�ք���&��]�5�s�i�۫��.�bvf�L���_C��Ýk�*c�o�-�k�Q�X��T��?��=�P���e���zT9|�)V����q�Mk��w]u��<���C�����ˉ�U���!4Vj�j�wBzU�`�Plܼ����1K��)i��ڙq��|���p��p�3*];n&��U�<}�ʮgTO&ޡ��1AwK*���e+�?6��j�ͬ��9ۚ�kaĝ	���d�j��yѾ9&	X����+Np�FE�RF��$��՛�x�2�	�
u�+�2QS��ެ��(t�^��#y���q�O$vTZ�[����E̭���޴z�3OB�̳��x����@������(�u*�*��������@�ًCb��vk!��gU��<!\�>�b��jopē�%8�*�F(��Tս�	H+!�Y�����i��R��z�Z�]�Ҧs���mG�������j�<̑�}���$��U�@]�{��t-Auf�=
J wZSJ�{���س=�S*Cq^v��e�22�s�f�*#�v�¾���{��.�*,aˣ��X�,�µ�]ZE��]����NY���ڣwþ|ʏ�L�r�"��dF� ������bQPjQDj�8E�%K%
Ĺ�Xt�D
&UE��Ȫ���S�r����Ԣ�:�#�,���H�����EVX�Q��9ȬS:Q#�0�Q�IF�U�2"(�C�&��IR(�E������-�T(��
��PU��#gB��kU3��5�.Y���V���Ujg�Z��,�R��D͜�#��T}E�ug���N9�I��C�����9���!'t�ԋXYW�+�zVS�^i-S"=9F��QjQ,�J	��Qy�"����Ws�SԹT�G��4H���u�ZI�\�0��G:Dg��"'=� ��!rs���EG��z�"V�'EԊ)V��*
����EC��5��9�Ȫ3�I�J ��Dz&��Ȁ���'�Gu(򤨩0!]���	'��wv��%BNt"�͞(�ʈ��=�砐r=�r��#�t��j��n����i��N@o_jS76������c���;v�����>��p�\��\V�3�bڶ�Zj,|��ꯪ��R�Q߽�P���-�{;���7ŧ� ����V�5�����S5PL��y-Wh\v��Iڕ�_�G��������m�*^��Y�CD�<��<��/i\IP��qi�T�2G�{uT[���[��|���V�I�Q���W �Q��juBZ������N�W/�ԥ} )��8��l��Yؔ-�G�����DmK�u�{�~��[��^���`Ń�q���V�j���V���؁C���T�l��1Pu����[��0F1��s���[��O���*��n%B�Oy��s:P6����^���9��wQ��/�5ٮ3j-���*�����c*�����{
��K�k��Ci �V�'�*�P��}�t�]dG�oo��ӽjwٞ+�vW,�b�|�s��a��������У��,6�6��n�@��7�JI�A�R�����a���Y�s�[�]���VY��2\��[���?"w�=m�]�V8
��i��9fo��s%�t�4.;���1$��ʔ�6ﺊ���E���6Qǻ)�ۣ0��?{���W�K��>AY�7B�8�e뚎��7ܞ�s|�9���WMg<ۼ�sT*l�I-0���0��l�k���7�+c�mjx�+�M��X�3"Of�j�Tˎ��n5���dLr>���S��q:���rn�:�6{e�o��;�5���u�p�1��w3��z1�.Һbu9[���6+���D���{X�ƾܬ|�ޅ���t6��3���b��ZCŞ9+�&|���پ����5|��LF[�~S/QO_k���7�L�[�����ҽG1�^*��Q=��&aq1i�T�Û�>3Y=k�Vľ!o.����(��~<!�L��n+�����	��D�����E����ؚ��rwB��Dv�˵��>������.���Y<�3�5��5��b���3C���Zm��Ol������y�޼t�<ٸ�k�E:�g�]ߝ<�lq��\�ρ��)ЎmǷR�k��.r=9,JV��p7�C�.�.�=��R�A�S[:�`t��(�/,Δq���_G1۶���t3��[�ae�%�]� ˩�����˦n��b�+?�����'i�Y8ӌ̹ϣ��ԵF����k������Έ4�@������X��Y��{Ou�é���^*��4Ryq�x�f���ඪd�zl�~7��6��T��,z/�ϋ�9�<�B�����o�>��D*�-+�V�y(��#�41!�Amԕ�T$W�G���F;i�Hu�m7E`�X^k[֦�:�8n�b#1�?m^I����Ɨ[�ԕP�p ��\���zj!7��@v�U��l�Z�{=�Z>�^��D[���f	^�+6���ֶ]C}S\�M��~W5���Z3*������(��w9�o��v�K)F�����p���X�MClmu�8��u眆�+{<��=
�Q���ߨd�5�?>��%�|��<�^�c=�h)-��\����G6N}�e�u�2��@�Tf�AZ/�7�����\̷Qiy��#�5?��b���c�&�)؃��O�X�h+.��l�>��$�b�`,�/kD��ƺ��Qňe�# Щ�����c���cTĨ]���gQ&�^�M�kj>��)�εQ��"�2X�[B;�ّk�l�N�3�WY!l�ص�qG��G� ���k\�*k��C*?^O|�׹�ʂ�bت'j�w��ī/��{���F�oo�V����[�Z���u�۳��eAW?X�9�;Vo��*vi�,U���躷ac㮰�+��6/Λ�=��W��r�GG�՚��㘻|<h�f/O,M��5<�-WF����m��_=��g���puHt�\_X�ډ���9յ=*��)J؎-��ը�SO�l�߲u]�c;��m�P��
0��(ݤ�)�%�!'{����O2��mh�И���U�����)J���邏���rG�S9<��<����_73�;�_(֮wq�m�܄�6���8�S���n��3O �Y���:�ʮH���p[J�;Գ��
�leC�P��R��Z�m��%4��yD�+���_n<)c����|r��5�h;A:��(��!����2���|:Y� mڔ��`M��0H�������(VL�7J�d�%m�V�5r-�lY}Oּ1j�{V��=ޓ:��˶T�3]An����	e�san�oS.��f�vn����9�'؋혥�Q�b�j�9��ն:Rn�-T�=.{�d1S�U����N���fR�܍��oMz�v��y=h�����a���+vɚ��m�N`�������ZF��w�~ZR�'��U5){��+f��ë_c<jO.ܯx��}f*�|��Q��~[K����e3۔��ؖ9�;}@�1��g{�%{9?+�^Y�G�r��jq����N��VH���Sұ�v����N:���fg3���S-?��8AR��=��zCÂ�F�����ž��~���v�6-�-ns676m�ʎC3v��Cs���y�C�2XOj%�i
��Zi��T�[�U۷�z���c%gEu*�ur�}4��a���A�^�u5:�+��X��y�oq�iVƭQO{+�ƾ���^�]m3jam���p5/mK�q]!$V�k*	.6�lRt^�2���Y:k�[�����
1��A^|�i'x�5�lf���Hs�2nk F5��Gzmy,���״�V�G��j�R�<��_����ib�񺾝�vr�5"��6]^ښ�4�ͣ]b��by����jMo*+�a�0����ٶ�|�6
��.�r�������+,��^5ow�bCo7���}�}�|�L��/L��?Ri��z#]�h��~%e�O�<�Jm�lu�*]46N���Ӯ��ʵ\K|j}�����m��)P��;��/�4feqwm�X���yh����,�Op%�
����-�{�,����!�v��o�>(U�n��f�is�Ub㜚Pք�;B9.E�ؘ����+��ui�@?*ߦ��X[��^�o�?`�R��mB��Q����L�~��z��(��CfN:��"��/�KqX׋v��jx w�����n9uM,�&�q��eN�"y��,��n�U�ݰ��+dd�
�X���m{QQI��o��ʩ�/O�Y�8�?9~�S�2��sS)#.�'�����p��n��X�9�녯��t7(�B�c]�����+=�
Λ=Z�PN��f�בZ?w(��|���S���η],��93�r�-n�<D'ē�� &XH���ĝs:Ȗ���{���(0��6W��y��uF��7��v�	�m5l��,ͮ���p+���0���XU�WZ�BsiK��<;^^J�:��7���\�G���]*��,<�%��7���U��W�s�����h#%�hE�_��gU`L+��m4��Rlm<YW�ݰ��h"�4�]��wV�Q�� 򠫐w�i�קT5~����Mzfk1Ղ��jF�q���C���_n�ν���ك����(��G��d��M��ߩ��4���C��Zm��OD�v��@l�����t�6-��#��ٞ��˭�{o��5��b|����P�v�5Q��1^\���E��{wMƖ��*�[�PRy|��q�O8�fH�&�y�5q�of˵в�
��8�	h�i�"ެO�o��;}�ܵJ�a��l	��;��f槪 ���C�e��	H`��V��2ެ\s#Za��ʹ��-E-�c��Y���m�Y��5q*��q�JT4��Qt�"\�u(z�XV��Ֆ����Q�.;��{�9��p����D��8�f���p�+P&���,�@�R�k��Ջ+�Y_�L�L�6:�+y޿P6��% �]z��>��k��v��i�d�e��Pm��jݗ�Y��Vn��5(�1;eςU��}��Y�ͨ�h�<Z�H����IS,�r��㠟]VH@�߽옧��P-����gm^���u�MG4��n5�+��tD�j�r��V�5[�==L���U�m=͉���u�I�ז8SM���0r���ƳwS*�ԵD8�E��@�u^e�.}��kr��s�ֵÞ�N%�=��iR��#�"�s��A[kֻ��U�6�ĭqڞ���ET��e���3�-��)�M�律�����1�]~q�b-U`��ޞ�Ġ<De�R��,J�7�љ=�?{z#=4�>�����p���k����ښ͠��w����Q��
X�b��Sٛ
�b��:|=&�Mo�꙳����	��t�CW�ҿalS��_�o�_=��61��/2Y���'J�3�]�꾛����Kҕ+��ކ��-%�$Tu9��ϒ�ј��P(.`pQ��Tm)��k=�I�f�T�~�XZ��y����p�w��A޻�˻��,H�^�����Y�q�p��k=�:���vQ�eS겵<�xs5Ν�)W��tx�Z�2\ӵb�G_7���5Գdol���l�8��Kpv�dS{�.�ԍzPJ�-q��q��*�ű)@u�f����ݪՁp�����%�<���U�5^F;*�I����w*O_�	!���r/�O8�,���I�&~�|��ڋleD9Fa���%�R��`rS�n�"Z�(W��=!�����I�4� ;԰<�P�^r��!u	J'�i�D%�ƮK��~�B�>�-�.���^��9sJ|:As�*Q���:D��VpߥjS��X׶�|"��|�'=>MP�T�4ø�0���-E藬_sP�$��9�/h;r�s�������߽BEL����.��I��x����Y�Oԙ��K�^?[ϬŵW��-�AN{��5<��}K^�B��'k4su��o�q�U7�����MyfV����U�ƭ������g;��s �<歊礓~YIߔ�Ս�5��u{/&9ٺ�C2��5�0��NyM:\��{_O%o��s�]>|y �b�n�osm��&�b��"��VQ�ʹ��rk�b��}'⢘��t�~�饨a��Y�e��>뉗Հ������Ǖ9b�e����ӷ��u��}�W;WD�J%�=��랢ѽ9gtO����$�4��jӈ�0�����	��J���D{޹��q|ѱ��ۘ���ݒ��6-4ͪM��t�ڮ݇��-�y��f�-[ܭ�U8�vr�C�.����u'T%��E��ޜ��3�m8��W��JA��<��َ�9QL�s ��.V�t�Q�R���K�G�!-e*��4s���\C���oPb*��=Dzv��'�3B[M�CԷ�{��L$��'.K�i�놶�-�E�Z%(���}%B��Fe<X)Im=*�͢��5~�Z�%�5�ˈ�v{\f�[c*!�U�;@�u=��iX7g_]��mv(��t�\F��g�ޯb}���;չOt[b�N-�-ݗ;��~T�y�s��b��ͥ��T�b?9��A�^V+���J[��c;�=�1yP�#1�9*�	Z棩v�rk���hW��q����+5W�2�u�����)D�r �Am���=��e�Z$���6k���I܃���qm�����$֙&�v���t[Z�J�m90n�"�ݪ���p�a]�&�I�8T�&��B˗���#��'P�qڋ/6������]�s����ȭ���4��6F�иӆ���V�P�\쓷	iL�;9�6���0������A(�-�D|�����̶N�RnU�f�0������"��^F@�}W�׬�k>�B��:�m>)닚�k��`0^J��W��ѰM�xX����q���[�t3J9Y,X>*�qR��Cv�-�N	3>��\�����z+������Wozdy#&r������$iK��0��W��c�Ʊ�-��!�X:�;�z-]7o(�&�H���}�҉!EԋMX�$��?^e��V]����.���Xu�ڰ +�h�ıa'i� l�*=�]]ָ�*�A�l�L����7�h�#]B��2��՛[��8>�ΤV#�A�;k�L��h�bm-����I�A�mN�����c�4Y2q��f��m�X2����!X�Hl��֑��P��"���t-j��u�)�HLk�xֳ�*�A5f��8���ћ2S��z�E���AD@��������N�8n
�3N՘^Z[���v[ؖ�ʄGk b��#AwGa?=ˡ�y��GSv�y�'k2�=��[�8�R>��E���w����z��ڽ��� T	�ַ��gU��}��j�HA�v%��έD+ȶ�Q${2�%��2܆S��N^Kw�|l�gnj\���\���yr�b��I���JZ��Qݨ[;Z��4;�e�C�
b]�,�l�aat�j�FFc�6��S���t��mbn�EwRe�к�Or����>�;R���VPu��4w�j��y�4��C,V���Ca���ܭ��j�玀W��\���yS׍\�y�wW�U�V��4�q̲�Ek���_V*@�#fl�ڕn<�\�/�@4�Tz�z�u�1f�r��-|љ�i[�C�}��X�/��L��v�M�{$�]\\��� s�+)�Q�L�O���D��ۚ�8,4,w-#��c�]�=��ͧJ�P,cK�ƴi���[�EnC}gdH@D��@kV�k��$ђ�&�:�6�ح+�!4�e�����F�混w���Yq��,�'��J���3�{}3�(ث���)�@��-#{[�Q:����x���k���]u�Ӛ�Lc)c������m`��v��^Ĥ�D�C�P�̵쨯�n�xW�/��@3�p����l���2pٔ:��-Q���Tl9v���Do#�(���I�/������-H�[uoȾ9��B�
G���o9FVخ�v�N�+Ar�������O����˺F�Vl闘�
3j̟-ŷ�5���vr	�9V�g`Y7��WI�8�R�\wL��Xu2ue�*�[Zo� �P`�h�]��Ua�.�.s��) ���B�u͑Hp�2@�5i�q�\��s�ą���K�]�76�gt,�q��RfR���J9ㆢWw)�3ZuhQrQ�QR�\9UU�R�(�dʤȑh�TP�)D����,�9wn�Qt�L�uB
*Ia��Efi���K\�J�Ar�Z��N\.�Ddb���(��E�,�"�S't�M8t�fʢ(���&�HIEs���tP�)I��#�O%ԮQEU
��A�t���Zi���+�b��t�#�"N�"�!:ָ�0�閦H��;���H٢f
��=S���a��EG*"��UUJ�MC0̜��:^eQvET�a�D�&�eG ��L���X�Wr�����̮���hQ�**�iDD�@\R�	�ʈ��EDU\��3��U
]�p�Tֶk[��8J��ݲd2��}D�ښ�����Gw�E��9S}% }�$���4��`��oJ�����֯�m�<$����t0���Y�My7�N�#��赹��5No��H���*2��S���e�����{Q�դ�k�=���;�Tk}[E�fC��f��~�%Pef\�ứ�nV;�9}p��Y���\��� U�Tr^B|�F�v��<�f2m�Z6���c-�S/Q�'�t*��y���w´Iǜ�����n��s��C�{'v$�!����O�ɧ�w�2�A-����n'��oy?D�2��#�_��V�[�ͬR�<��+muwW	d�rt6��T�h�I��v�\��w���9(�<�\ʯ-ۡ�_9;^^�קS��r�g���د<e�o�'�kf#��U 6ҩ�D��6�w'���vOS�X�6UzR�Z���f8YК{f����4K��|��f�N�7��B�Z��.F�JJ�Pe�!'n9�]��3p1L�1����3B����$���3e��L��q��+���7,��"h*�j�VT�ZQMۧ�7�l ���s�l�G(9��tCM���N]�5j���Mf[9�'[)L���o�t�:��v�آ���Ļ��JŶ���*�Tx��.Y��U�U�7Ў�=�����9T
�|o�Z4sW�oTb|h���ÓW�'7Nn��Jn�s�le9E ��)���+�`[�18[�sj�f^�3�G%c4��yXw����oЉ�Aw1��{�X������k����Ƨ!������.r���vøWP@��?p U�'�r���b��Wn^�D�v�����]y���i�m�>W],��۸�}�޹�6��4-�=T�}����_�^ֺē��X�Klf�QV�g6��H:[�B.Y�(��3:��ˉ�ϲ;���c�r�p�BegE�96ķg�%���J~N�ҹ�F�#��uᘨ;�+F\v�}Y�07�R�H���|9�zUӎ��g!>k���דߠ/�O�ӫ0� q��In�,7�ƫ�.��b�N9Jl[�[i���ٷe��[f�Dl��S{�A�i�,C����X:�i+g��R˵�e�E���N/&��}���jwX������5�,�Z�Wu��\��m�kIN�ә�k�I�ϡ���*,��U۳���,r�3p�ʌXˑ�b��&=ɽ1�m�<�`I�q��u4�_5`��U���m� od�����J��X�b�7�SZF�Ԩ�Z�z�T���%+.��@-�Թ��	\it�#b��k/ɷ�/���+�n�EU����J�vr��%��jz]��¯JT�7|�5�+��rR����\u�{^�B)8���f��P�`v�����AԷ������gH �>Q�n%��O���-/�R��Lw�O���В�Qd�	��յu*�V���R:�N�4[�o��ڋlc(�"{�12+4�W���\���셝kwM+��R�v562���]��#:���A��w<�v���-)��|�"n���CZ�Wƃ�)<@�s�r��e��Zh�sWK�o��ִ]C}S\���ڸ�k�=��s[�a'���\����;��p����Q)��
��F�������m���b�rs�v��kzi��g��9[97����=�Y�u;�����ͧz�#��:��s�V��f���u92]]9�b��ɝ�G���M��Y�'׻�b���L�:�]C���y�6�UmvI�`$IE�k������N���:�S;�
~�6�]�ʝvG1���@���{���\� ��q�%$�r;*'��--�اz�"�c�s:��F ��g�boO �]H�ka���Ӟ�7u����L�X��[�����5��1YG�U�r�9��v�L�eĝᷜ�-��Sb���u��.B1U�3ʆ��-���NG�i��*� .U�[q%CXR|�O$���5ҙMQm��c�#����m�
�(����U�5o�ͪ�*B������Y{L�Hj�}�O\�>��ķ�~5���eڷ�a��n{!�^\���L�sǯ8��E��;���co��h[41T�5Q�4=9���ٖay=���f>T:�[�^Ԟ޸ko��m_�Dl�{o*��}菼<OoZ�;\ܗ�P�Z5_+�Z�[�P[��mj�q�Q��󔷌M�#�p8E2s&�{��_&qTA�2�J�*:'38����������f��{ݿ\]�gV1m��[V�]m�W{9;,Tw���J�cOgV_K@���`�W*�h�9-lh�C�R�BY�F5{NB�)�ˣ�k�7'����"�O�����^��fx-�O�6�:����C�5������W�M��aq����	L ���\�-U�����س(^C��4�'��A�d�Y�_�[��&<�A�)F�+\������S����I<��� � �8؞�ͪm�w�\kW
Q3�l��xu��/�.r�Z7��h�犳i��ڍo�j��g1)����c]�1�t����OnŽ3�P+��O�����^��k�$떸s����s8��*�h�f���i�MGޚmz��WrT2w��h�=�,�w�_\-|�Dk���dʪ��d:ԭ�=�d�>�m��-��Ў�ꅖ��^#+a�|j]���g%�iOWx�׹K�#]-�B,�t9��Ĕ¼.��[T7���`ڣ�[��?{z"�4���~�~���u'�p&X�=��n�,K������U_Ju,�w)f��^����a�LD�$�7��j�F�������P�7E��m,}�D�*����t�
�̾���[x_%�����܎��e��_>��J��W
��x�\����V�:}<+&���N���]9r���p���x��p�u۷����k*���͑:�۵M{��u�2��M?*�5)Q�+�-�x˞���l�#V4C��Yt{~���7^��P�A���ڞ��E��5��u��SO65췶��M�+:���-�`t� w3Q�%�C���sƸ,�qnn�o����{���I�>8�Z(.�삠�%��O5���1>'�9.�B�w��R��6��Tn��l��lR��X����9z�:�����.�\�=.#wNTsiXw��y������B'��Ər����h���dۛ\q˖�{wn�1�ʎ\�7�æړ 󖇷Z)����3[Nxduۑ�����M�ڸ�[Q��P�T�G4��n5ߕ�UI5Fl�<;(���r!�hr/v\]�u<���\�؄�MB�
a �<�m@S�"��ԩ�5i�d�b��� ��C���F����4�g}��dC�Va��ݩZV� �L㕶@W#"������Ӳ��4�ͮ������ں:����׏�JY��Z��f�E*Ű�)�^�M�7w�ևSc�v�C��l�т-	7�[?R9�!x��>�4�|Fy�Yӽ��r���Q�M��S2Y�{�n)���=x���̭���]�m����W�m����C���U�ؓ�[T8��K���r�9����}�#u�fTq�#�Ȑs�3"�FCkYyWx�N��
�M8�)�_x��zw*�������Ƙ+*�z������
�Ku�T5�����M�����Қ��i�;R{i���' �u��r���sS����`l;���`�,��,O-u@W
�Ϛ��IѾ_vَ���G����Z���9���ż�aN� S+l�ob�\�t=M<�5�B�O :b
�򊍤��1P�o����0�Y�K�;��=�Þ�Ҽ���ڷ�K|(t��O���u��ٺ��]����	wnV��?K|C}����'�ؽ�P
���t㙡ʰ,	�����p�>�ˣ�_X[~����Q���+���o=�]3����<��t���n`�;-�
�-!\�ٵUEH�v)EJ�:���au�
���ޝ����[;�'����bX೘�#���-��˖_Y��d�t_B[nee5&Jnr��U��Wߺ6�	���,�y�6/\�%\��׽�79;�0�|��W��@���ҹ�@M�>9\���p�������m%���t8���9�@ے��E���ִ]C}��Ԛ�`�E�1<M����e�}k���'�^9j�#~7���(�痝��4Nqնy��u��]S^X�Kn1��T�'���2�#i��0�,�x2B���ok_s[[�}~��u�k�=x�k�q��bb���6/r�K{,�ݧ-�+pf�w���r��S/Vy����u{/'��*8�D��`RR��z'z}C{>���"�䗩�����RSb�b��1p=�r��Q'�c#efkx����ʂ�C�Q�[q%CW�.'֚eJldv�k�7�Fe�c�˚Yxg����i�~�"ʱ�����l�!�5�Y6��ٌګs�է�)�o �*;*C.��
}��z�$�)���L-�om�M�W}YJ܏��Av���K����C�b��{ʎ���cYZd�圲��rd���K�n�R�!po!ɦ^��I���������:�0�j3�A��'��5r���}���v���XsV�wE:�KJ8��K�$�qݴ�4���5���)���bNGP���^ݯ3dd݋c�]8���[�Z���m�8[Qo�٥6�m�O�<�/zZ{�G�� ��,U���7���k��m�8����ɉ��=�7��B̉���1PR�Q���Y݉��m(u�.����c�;ySt����PTp�Q�;\@���y��y�j�b��cG�Z|���.3�Ry�ӑ��0��2<�A��k��dM�,�y�6My���ޞ��ً�[պq��4���q��d(��CfN�u��-���0FJ��.T��;{��=����Cj��g14��w
�}���;%Z���U艪m�R�t�mk���s��^k�sKRu���23b�ͮqY���+ו����c�a��1V���	�րۆ`���O��c�q�u��Jo[�q����x]0�@�RUwgW��ʒ�{�QO��]�J����Q���*�jβ�sVR���u�w1��LU�����Fl�iZ��4�u��!ދ��`ټ"qKpo���U��1�x�̹��o۩��c�^�q��s�vT�߼k� 4���I���Y� ��[w�v�5����m�}+*��yx��)�`~�(��x���H��ڑ���:�p�����3��O\q��.�%�;bg5CN��ظ�M�7٫�v�������4"ʱ�N�=[%�7^D�>Y�b��\�w�*F�DsM�;o��f���9^���K�r���N.\�*�����9]��OY~M��t�٭5�4�V8�����J%t�S�/��[�<i�&�I�j�������Uި�ѽΚGT7���[�35ʠP\��������*�[�PRxo�dh�z�����u�X���{�������!�
c��/%�cO5�o��-Q�IsFq�J7h�=������m�eD)�%!�R��!-�M���ФY��H��ܠ)���������u)=D-K�3(�)�m��Z4Ѯ����ܝƦjQ��j�;z�4,��j�L�0�T"�9�� �љp���:�!b1@�o*'�2.���V��A!�hU��ԯ��N�kyM�I�Tt�e�����6�fg>��Q8�^i�z=w�`Z%�����S5���4�҄L�b��)G6�� �j��YԈ�on�ʴI�hA*#��*�k�*esa�V�	5�[,�t携���fJ���X�*��>p5�-���77Y	�ֆ�]�K�,�����<ʷ�-Dk`X�i0G��vm�Q�zW9��I��d�`l��S��Y�U��Y�R��I/���]³k*t���[Ű$��dL� �u��n��҃9'5��+��S`�&!H�pv�CfR�RK]�T�B��}v�8v����z�ж�B!]d����Ue��+y���8��a�����W�&�`�V�/*P�]ˉ+�j��ڀ��v��ΠU��l��V�-�2C�wY���}���{|��fN�vV%��w���S�+uM�� �l���dՋ�:��ev3&��i	�kp*T��l�[�"� � H���l$36�����x��4��>��t�F������n�G&]�<�T���{���ފ=���a�L�o�k
�[E������"h���nC
� �Z�'�yC��9�v��(�VJ�>��|u<���/Oe�b����@ڜl��۝�^�tC�Y׊�ヷ����1�唗�yu�\o%՛8�����S�͊�YC���T]�o$�A+o��1��X��� fV�����p̮��;Y�u�B��݀X� 8�(n�5ka��k�������U���ڧ�i���V.�Y�/�f�jL��A��w�F3����UÆ�5)����4������c%��Ю���u=RS`�1]eW_�����O�oC:$�v%�{:�O����{,uE�f�������w���Np��(X�N�|nv
�"]0P��JX�<fVtB���U6�kz��R�eZ|��B��[lst/B}h��o/�6V	N�ڏ]Eqn�3�f���J隒����]G"*�,����x�}8�@�st7m�t\�p[ݶx+X�H�i"I��M�8����
��)�x��
M<�e�X�94���H�.�<u�;� ��dw�n#eI�����'Wj�|����2-��Tݼܼ�a��]��C�38r�9�] R�R�S�O��d���E��0;�:��S˙x���|�"�Ӱ��|;��Zr+h|8�pk0u,�]�Q��
��S1n�{���L�G ��i5�"r�^�	�v��&GRoSX�F��(���:g7�Wڡ�����aj�ࢳ]��Y2���85�+�w]�Hl�V�m��)��-����ڐr)˺��o��XU�� �(P |MH��L�UZʫ���@ŗ+�9�	�9��5*�U��Q�F�Et�	-"��ʰڴ2KZ�QU�d&�E%�NIG(���+��
��Q����t2YED���,���V�:r�"rs�\�QBeI����"�.S���r�#���^�B��tnqȪ�ݗ��u��*�kwB
e�J�ws�2�<����zlMiC�财#E�HDUs��i;�,�"=B��wRr]�R�Zehyݦ�Q�z \�8��Dj��Ĉ�\륞{�8G��E����-٘W�r�8b$	����p�v��Q�D�tB�"����:��(��"���U\���s��՜�O>.��ٜ��z2w���%9�3�G	��n������֓k�
W�H㣉��Ւ�[+%v>�~D�36�U����֣3��]��#sF>9\�V�y��Uό{(.�^�ߝ����,	����@vN�vf���1��\�5�?l;W�Q0�n�n��j�K؞��M�X׿[8"���5���S���y�mS�bk͸�nF�wUb����8�k��$��H����qv�N��~�{Z���ql���x�����ͧ�.�Ȣx+3�z�W\�;"b10-mΣ/2�<��F��dw-�l�=�S*�b��������{��mo�eR�k���&X�#OgKI[��!n�JԵ�5pOܒܞh������"��W:�iDo��l�&5:١��kuOms��ҿI�:���ӋR��m�k��vݜ�qk�͹-��ǹ��(m@Z�Um�P��p�b�&���z��%bp&Ȭr^��j���W�,q���|w��[R�uBW]+�د<d��'8���g �D-�{�9��|5�˅'L�]��E���~�G��F�C(QV������1��\�dq`���p�X-�r�l���vK�	�C�i�mt�i_bM3E-�k�Qj�ժw ��C��S�'
"*�`i]L��o SK�^v�Hݓ�m1�ԛc`Q��Y�D=����=�a�[�<u��L���q	6�}a	���2m�}Iyx�m&�٭�������/i%���R��sV^�"pK����w��=5U?W��u�S$?Y���ݕBSd��Ht����Zu�d?3�^:�)���u�o�!8ͫlc(�!%���8��������]��+$W�H9;��{]m�M+��R�0TBleߺN�Y'1M0���yt*.4�T%:}5��s�7^��*9sW��>�ع9��r�J+;��*�q���l�νn|V����;ɨ֋�K����i�3���Uz�_�Z
�q�����'�وmG���q�9�l��V��+9�?���{%^�Rs]��ɪ�X�Kn1�ʝvG1Ϊ��mq�����t�u9��zT�$��]��j7*���X�N��c]Tkb�4w¯
�u��荿i����T�Y�ft С�tf�33J��
��؍a���c4�&L��-ѫ{Uؤ5��'D���3��ˍ8Jݵ����1ǩ���:&[��LT� ���V���)H���]R��ͻ�soG��\�Z������$цpq�?�S�ܤ��e�l���uF^_c�Y��*�D\>�`^����e� X�@�co9D�e�v�Scj�ô�^��=R�OPL�M*�NtŻ9\�`Ua�9��^�Lz����턓�/���0���~[<�T֑��Eh��~{B���iԝP��m�[�w<��S<{�b������bor���������̏R�T;��X�G���(q����),�Q�X�+��_���z��{~5�B�rw�U��}C��nzba��Q�/�z�^��ףR{q᭸�j�-�4�ӳ�Oe8{�'=��6�
q��\������w-������l1�[��$���{��q�={o>7�=b�H�[�.�}<��zN�}�aҽ�Y��+��Գ�M��%�*-��������Պ�5l~]W9�&�>X�m;��p��,�ɜ5B��[�����P��#��	���;�C�;ZޣS[Sٜ��v��02�M۬��;�{�v�1���b�JfC�ד:v�J�e��*_VJ��ⷊ�:��Q�!�T�uh�Z������3\vg7�r��S�[�����+�\MCW<lHol|&�6�� �'��J�NF�����q��K��Co���y\B�L���0@�嵻Pj��.��}�������y����j�����M��Ds|��a�*<	�8t�ںBm0�B���ݹ�ή3^�I9ֵÞ�FKu�nճي9����"�Y���[����˞\7u5�X�#��D���<�hGq�y��))�7��;�'-+~w�70����9N7�k���w�tС��b^��?jF�\��ir���4���W[�갸��o^Ku�ѐ�/�x/�����sW��ܾ�Hl��4"OB%���Bd�FmA�<���jj:�%z\,��$޺oS�ݷ}1{g&n[И�0�*;���9�� �Q�.j'\X�+�بx�M��t��k=Lf��(Q�W�)�=�z-����;���}=�7���7�����|� {E���4����"��b:�i�+�e)��z�˛0���w�=��}hS���9̼�����1�u!�[;���vu�ZΔ��lR57�^���8�cz��L��tmN����[wD�����7��<���Pb�Q�=.��)I���޸k��X��؈��(W��3��Q�m��0:`�>�״��Rޕׅgp8���G��F&�[�\�������������ފ��ݡ���U���̕���ԁ�ku�w@v�S�m��r����S��Cº�F�*��{g�g��26�g;�����>�޷�l5q*��q˴
�g�Ջi�Jc��QԻv95��r�<�����\eR|����� ����'p:�sSk���w�2���MDsLL�Xb�v�X-��ʓ��&�r�Y�~��Ѥ�l������8a���	��0�M�J%�W����P�U-g2.����c22���:w���T�^2N!s{�����M����Þ��v6���k�u�C"��n!-*�{�B���:����f̤�<�U's�-����)+i��8�Dp���ںX��Zct`x	�����*�I�ƍ�x��m,ydx�U�� ��m�l�+75�m�2��iIm3�S˙�t�i��=}JY|!m�w.����̣go;�:��>Ӝ����'Pǭ���p�^��O���B�:��_�-�wYє7&'����W�ުpډ�����u�Qi��6�ͅ��Ժx��[I��?>P7,�Ur��Dꭸ�����$�����Yaؾ�$[}${c��fg��/�P�>UmK���	_��W���眖�UW�2������;�M�3Y��AYT����)�ʣjz\���u
�3K������{���q�T[���!�t�pQ�:�h�~Y��6w���op��s��*~zw�S�p�(�k��eyJT(t�����e�+[��ҽ��w_<S�ҟ��t:}���6�߭���3��U�tV��e�%�����łS�ZSY�oTb�ۂ�Wޥ�����K��߶8�����
�#��������]K���c��\Ј�G}I�X�|7w%�fZ^֥.<�+t�F��%�B_:I7��/n����2�_��-P-iMӷ��]fw,�� �`KRm\8���'�Ou��;"����;X��w_d�gnP	���m�"R�U�JA�˕��0�u������X�J���y�: ^F���g2׾�}l�Йe9j������GcXi9�[�t�3[)r��y]w�ɗ�0�7�FBtD�j���kU�o؄y��$�[�����t�Պ���P�q����5��O����y��'��`��d3��h'��h(��m.��9�f/W����B�؉Õ�+�='��9�j�k�xfh6��ѝ��nRv�^�����C�/��n#Ȑ^ӭ�{�Nd����m��f]e��co9F[��S)��"��2����x�i�X�bιU3���٠�'}���\skj?`������S�C���<\ǼgZ��K�W��G�#
�QW>Um:��,y\���^!SS�9+�;N�&&�C���_=�{8�7�j�<�@r[�Ἄ�k7t�T�K�,��O--���o/}p�=�/c�1T�xyq��R�LX1�XIM>G7�˘�]ʝf�Zaè�K��/2ҧB]�,�Ĳ��A�FqR����eb"��c���*P����'�W�M5�c����ݣ5����z����@+��v���D�C�Αj��,+�`+\�,����m��W�U��JQ@s=óvKO�Pu-�Ԟv�kq�η�v֌�pls�Y�OB�p(d�y��P`w3ZRX�K|j}���ͷY���"h+���Z�E'�l�)l

{����KE�� -�O��W�_��7Ntk[�U��k�ݳQm�e����h0y��m.{\���-J���](�e>�Q=/�Nsi(��p�P��¤g�.X4Nԝ�Z��ݧ҅eK�U��k��֎�%�j|�n5��R���4MHռ**i]r%�%�4����˳k��Mħ��{Ѯ��w�[�h��~9��}"�)^��P>qKp_��eU����X�G~��/*�V�s��Þ�[2.Po�n�=˳M�k�R���:B{s>�f�3��k�1o����O.{��nV=��T�2�1��lK6�mO4�sZ�gF\Ϲٺ�!�����+���v��F��i�Wp`kͩ�����ۣ����ռ՛����3ӓ̌*��u��n��pN�ۭ��9r&7�[��]�L��c�O�#��f:�.��[�)d�b浝@�*�׹z�Π�m�ҽ�R���;4���{�t-3�t���t��)�b�VqoV뤓X�����}<�?jH�|A�r���U����w������2������Zi�U͇6�c��㥐�_�cn����W^������.geC��.F�{�os���=��H]���em��KZ�H�� N��[R�ꀷ؝-�a����܀Fv��cr>�g�̨��U��W+j����y��ܓFҞ�A��Z��n��u���uD�5���Ol�T(t�0:J�;��)+�_�~#��so�~���Ӽ�k�輧v�Y~�O��Z4�<��w �s^D�r�n�{{�K]#μf�G�ۘ��������^��>��z��茧+���d+�Gt�˥z�S�T��g��7}y�s�Zi���8��cO�l�������a-M��##�fGґ�<��W�ϥ|o'�51��:"g�����������m���0��,�sl��L�M+~�țѹ����ē�Y�[��])F��Q�i����m�{-=�yg�rf�\���x^�VH�b��A�ٴ�5�A�X��G=�[)���%�V�4gQ7 -�����Ӈ��t�X�>�G9lWP�BJ��|��ufR�u�Aۆ�1���Ҕ}
ʶ�M"����/�J�=��7��5�o���u!�o�H:�nb��/�����tu��5KEK�l�7��`	�}u ���0���c=�_q����u�8#d�Ҿ��͡;U4v����v��T�Gc@r���٨��:ԃ��y ��51G��N��Ǖ�P&�����2�8�k���������	��o�րk�x�A�JE뛓xx"��؛�?6�6�wff��e|�}Yi*}��l�5��z��)OK���|�\G�4�����;_����p�-��N2V��;�k��~0���㣒V�|�b�x���_ܹ���9�Ϫ=��X"�R5��_�B���ڞ~l����c����t�W�Z�7�\�}xS�4���L�VdaۦlN
�q׾��5G��1�y�F�3�!�?EC+��}j��?���ty������\`����4��{}�2���w��i��N�ۛZ��S�QG�:T�eD��gȷf:3ҫ2�6�Hpl�]�q�~����Y�F�`>7�:�vM��X��T�I`/y��F���s�P��^�`���ǧf9�|��$5y�i���x���:�Ǜ1#�_i:��͸��+,.���IxU��X�*ڰ�e��m�$jX�aGB��@��+֜��ȫ���L[��	*��t�a{���0�Ԭ��}�%��\���Պ�)ZSs�s�b�M��oS�ި�n�X]��$���$i\.f�{lwt�c�۩��O�Bp˶Eފ��m�7�v��i�g*�wq�ym.� i�h�7M�"���M͝�7ő%�Ni�g3k���i��@���"���)����e�Wy#ʆ��X�P�����W����r�i�Y��
�مͼ��5���f�WX���uw��vVe[΁���CLuҋ�!�?���/��r�^iF�����7�K]����ҕ>�]N��ud���`���5b2�y)�Y��Ȼ4�N�[R��J|����:2�T��뵔/A�:n!���]��̫�[Lұr^] \����� �fd+�}t�v4^El	a�u��SN�q�')��$�$zM��3FrЃ�R��K7��n���7�<YC���%Kk�Y�EֽD��F��L4ST7����3wh��P��3���R��Պ�̔�U�*�Y��T���:����e�p���*�M;1��kn�/�n9���k��`��Wϋ�h��+(C�2���8q��+���M�eu�/ukx-7^�)]�o�C��7:�;JF۲k�	nwh4m��U�V��;�x�]G�j3����,b�Ҍ���o�];q�v#M�5*�\�@�c��Υ*@��	���]��ڽZ]�5�qYm橝Eq��l���V���؜Y���F<��u��B���Eo�sY]�����uR�R��F��fݸ�L͌��zw�e��ںk�,�ٮ��D��OMgXB���&�)�ISEa�P:Y|�f}��lB7��酴Uͭ-�\��OsnWQV(�c5 ԙIe�.�Ľ��{%�T%!VM�)(��Ym�h��;��]�9y��N�Lɽn�<tX��gEAe:�:i���l�_b���vp���Y6��@�h�U��[+Jɹ/��{y���M�ljς��L�9�6����p��Rp�]���n��0bc�%rKtK6x�&���0�#l����V����K.�u����^ZzTD
���t�g����cr�cƺ��8���v|�mWRM�kv��h,7�P'R�7Ls�gH�{n��Q�e˨7X��T\N��9]��9�.�wk<���.ݶqF#4���� �ʶ�ɏ�:_ͪ?i��A�q�N��A��B���e�S]ÔNH-�b;3����I�T�M]f��GD���5�N!�Z6��9WZ�/�J^U���l�$��X@��Bx������s>ks��j�m�ӽVJ��:���η�*k� �U������$ ��EE�]rN�I�K��/RAq���v�Q�nzѪJ�^w9�g*��e(��-A��'D.�QRg�L��B�K����F���X��܇M���2�<�-�纻t�J�y:�G�K���,�:�Q�5���PU8Q��y9�W4h���S�����Q�g��Z7"��:�p��wK�(�yz	Ner㈧��8Q�;3G
��F^y7!Μ���n��9��BnE���q*�*�%uZy1ʓ̝�Z:�W#F�]��9dEW�D��s�绞�!$�"���C��T�/P���\]�C2sqf�Pj���J�T胳g42RRCuʹ�I�D���:��{�&��']':N�F��;��bd��E����g<S���#�Ċ-R���|EQ�%@U����GV�T��#h
�hz�=�e��Zw���Kyc4�H�'Q`�L*U��о]���1�xI�k��a��w������g��H�P�ډ��u<7���{M�c���ϕ���/���d�96�#�s��[ί|��pg�L���e���:���9�}-׼b�u�9�a�mA����#�;�UvC�2̟�Z"bK}$_�]|�
�Z�8g�_����u�p�\��rk'�I�F�?��;'�\7�}Q,��
�n+�TU��~��\�M�Q]�Hq�G��J�:~�5�%|>�����]DږOP2�r�y�?�Mg��Um�?e�P�P~�b��������\+��#^|�.�4��l��܃^R��Fe�?N[�l���Dv�c�(�6�GQ�?wO�o��q�D7�H�c@r5�m�㲨(��d��,K�����`|`�rI��w�3���wO��w��Gc����;o.'��1���M\F;�;Pբ�^���{g�ə��B(��d�� l������t���\nW\1|�ۋ��y���@~���L^B�%ns[_p/�u�b��S��'3L�4'0�J�a�`��z� �-�������%�K~�N�D��;|�ͣ�V�t�Uɭ�����q��8��o��ۣ�Q�pE����[(o2�u�f�h����k
U�C�p�ĕE�=ILm�j�b�)o��3-ӝ�8��&�M���&��r�3$�[�(u)��:U}}Ʀ�k�V�e%p��"G�i�.=KY��6�n����L�����A�xk��P�)m��t��iz^I
���gs�u�`| q�gz�r<ܞ�t�zn:�p����YӒv�r����ў�p� ��OXk*r>˹_!WeҠk?GK���i�O'�{��9���?SqkB�����Q]$�>x��]�th��|�#�4<	��P�Ԗ����G�Go*ii�zK.�c�Ϛ�Xvs=�4�Z��������cj>`���]�	�-/��φEu"̷(N�&08�v��#��P�䄝�.�������f�c������x	�}�2+f{�n3�hv��	����x#И�ʯ"�bm3o<�W��n;�i뇿\N���C�%��D�����뉾�_��G"L�򩆾ָ�6g��e(̧�����\��9﹭ME��ʆ�D�C�.kȀ٨=$L����KT�ގ�&�^���r��p�|G#q�#Q����l��7��j+}�\g��� ��u�v�a\x���4��k�!�j��O�q�������ow��Pܿ�����V�t�������VMW4�IK�
����k���,��｜,o{��n��������86�h3t��k��,���x�bE������K�J
��B�u�yH��VY�n��͚Y;O_�0��k:�<�c��4tr�P^lNX/��lM��%t����9?A����g���V:|m)z}�*��H�vy�G�p1�z�r�E��;�5=�%{�G�KfI��������g�-�֋����f���Uc�y��dlŋ����Gdފ�k��b�u?+(�jl��x��\�za��N��'H��>��ǌ:w�J�bkXk���]�y/x�kC�{>֨5r���ԋ��'0�8su}	]=>���w�zV8���aI����Y�ͪ������̧�B��B��gmp�ϧ$�`��]���)=n��DޔV>5ݔ�l���$��g%�Q|���GY�y�6#Ϫ=�Wȱ1[�^{� ��U졳���6�s>�L���]Jb�k�}7�,v,�.e�t[;νQ�����Y��~���>��v�ME9 ���@3��m$ѥ����v�,�x���8���ȸoSQI��#ߪj;�Ds^��=FXOʘ��U��Zʂ��&��r#zN3����w��t/ ����H=?M�P��F�����a���}&�g��*��Z��s'5�;�#bot�V�B�������ĺu~�I{�f�_�A�2WI3����f�١k�/wiey�;�Y�d%%�f�=E��K�"QҴ��:��R
�WɇF�,K��m]P���W(P�;�>z;"%U�ao*���$��������D����<O�����E�"2�9&�e�B �Ԗ���+��q&���N�x��>g��x����-�x�i��㞭��#*�2��x��lo)��ӗ�c���뗾���"}-���E�χN��w����:�1{M��.s	�� ���B�X��n|�G��$ڑ&�Q�s�49Zw�)c�ߕ��M_�a��񨟮��絻!Η�%�[�_ܢ�KML�'r�y��}fOjhҾ^�W�\6��u!�y�WK\(ɬ�<�j��n�F�2�����	ﮤ�OPɎ�Eڅ9ޭӋg�ڻ�÷��h	���n���#�F��Y^��#_v4*�n�f�=r��ε ��%�lv���(���B���TN}�~Uo�:��^��*��I��k@5�v��"��ɺ�`�{Q𐶅���c3��b�^�c>Xw5���������7��>rg�?I^J��_]���~�����>�3��n���*|���N��2�9��*�,�ȩU�S�3�(���_.t��t�������6���0�7rTT�׷7�l��p�s�ݽ��T,�\��^L��+\�f��\�����l#�-)ò�[Y��掕���ג���=��.�ҳ� W��1�u�+C�z�L9�O]�6�׿qɏ��R��qa� ʽ�L�2K��)�m�ۚ�37W��H=��N��M鏳��p�'v̱���r����İ=c�71I��
n����>���R�K����xn���(Q{jp�Ŀl���3��F�M�[���d��WҸ�=���z��;�����~�~�N�ۛZ����$�#��>Q�mӱ��<��o�v]N�U;G_��:k���:��iᷲY�ti�~��&+pu�d�^�K�K �wx��!��v�-P�z�:�Oǅ�ԋ5	����]O���rڋ~�2�:WyT��ܷ���7"�}�=W��|p@|��Ci�Zg���S�3�tK�n��]���dYɑ���-N�4��>s���A}T̊��d�J	TA���-��~�u�;��qա�%��̨S9�NQn�����Z޵?b?;�ߓuCMD�'��LwA�`�G�S�/pra�ֈg���d\�lg�M��ǟ+c ��"~�N\�|p.�n<����2<�}mB�����c�bUx�z�&�H���{��ΜO�Q�j5�L7�H���ɂ�L���`O:�Dzx�
�in�P��T�_� �����z�����ouA9���}�# �Ŏ����یJ*j��/�#���CQUJ�f͵:�V���C�ڢ	d1�w��$y)��q�GyQ�U�p�1R@�pN	!��/gE39���u����.VO�B�%J�{Nt��b�e�Y����.Û��md��h�n��_o=�v�U#Q���|�@k���.�Oj���s������ʺS�%_h:C:�g\u���=\����)��m]B�'��1�����߮����kõ��e��FF�{�G�O̬3��d���±��ߦ�>:2��OwKv�u��$���eG�����W���{��%?f�y�V
����ʜ7œ�~3��	Z�6W�n3���X
ޣO�i2S�-����^��8Ի��ϝ-eg�U�㝳�>��(2s�e��C�[u�����\���z���n`v8�Z ���G����n�M�W����Z�ܜ��d��ė��	F����՛%}��\wζ�^���n6]Ttc�O�O2�"�s.~U��9\*NIъc���f'�|�(��+�	ڇq�T�b�_9�ލ-<7d������]P�U�'��Q>3sگo����e�A�3�H/ǅF��2+�jj��ou1���w�ܭ��$��/����5c������fهp.J5
*2����"�e�9����Ԅ��׊�i�[����b���@���u�:pU�u�ն�u.�OQ�DU�~��7�q�5��0 �A�$EN��f: �#od�����$,u"���MByHh_c��[x]����Q���Q�lj�T��� J�u�[[��V՞��C�O6*�s7�����}]ѱ7�o�ɭ��O�u�Q6v!�Q�*O����Ɋ��ߣ�W��t��8@�x��5v�vLw�K�"�w��微]��֍&ے/~i�J�Ң<@�(��ʽ���e��}�q�F�t~��u��5�Ѩ��:�7�mxl�\�3�����=2��;�����ǳo�c�F҅��8���R
�Ի�Q�zy��_]ަ�e��{��_M�}��nN:U�!������C�0�e(?]P���,+��M�^�﷞�;�����:(ѳ�Q���u��V|��?T���5�2J��2a���
�o��_�yy���Ln��p�����_#��Ypf�����Cn��9�`�y�,�Sf����P��Q�f����ۧ�ܔ7�;"�W9��C=���q�I����ݭP:k.PQ�jE�FO�Q��#2c�E�,i��!��v�{4�T�*w��x� �-���y�)�P�s����£>���
X:v��L��h��������l��6^Ui��3̞7��p��b�N����R���Ϫ$��}����/Η��*����,-�9�S��L����37>4�b�U+4FU�+0��:W,s*�/2n�ܨ�Mm�[QqXul�G:]�4-��q^H]�L��;�R�(��9݊��1��A�O:�u�[4������ɴCHw[��w4����>��]q�}� ���6�g��:=q���V�A��d��-0m:��~������6V�VY�%�Fs�0���8j(��|g��:x\m$ѥ���9�xZ`��ul�摊��ә����{˙��P���
7-N���5A�bK��Q��^Nn�jm��sT����;��L۱���Ή|s��y�l}�&�
�ǃ$���(~U�s�5�����5L��{1�8�UA�I�����xn#�_�ƀ�5��ʎK�@D�F������|%� ^,������ �����/��r��z�Է^���������m{W���o��xv*�F�,�[m�#��ѰG�}�<�A�2��n�<��Up��ٌ��u�t�:��;~���K��n���K�O�J$Y��6H�����g#��\��䭈�&+=;�X5����s?Gd�j.��HQ���1�_	�0�'�4j!\�Q��wڰFW�!A�Q%/?zkuȠ�}�HTG��&��偎����jg��b������=���(�y��͙�=t��c)���l�כ���ׁ�'��4�D^FFa��ݵ��Gz6c�Z-�
<��`�<�ƶ]�ZT�����5̷�ۣZ�w��HJ7ܩfvӗm��v�̛�C�k�t��I���ޭWβ6��[�ޕ	�3��&��ak7NRR��R������c���#]�ʾn�k�(/�:Ԃ�x����jG��.hδ�������O�GՖ��)h�wܧ�=�u���{\���c�])�����n����[8������Q��Yl\*���9��o����L����+�󾻃�|����?@w��Q��2�Ϲ�����;�7�9Q2����t;���:2�W�o�*1��>���?m�kSY�,C�9O4�m���z�[��9���@/O�땧aO `��{5)���ae䛢^n'���q��7�6v��^��bk)M��<K�c�lΨQ�����~�һĺ�y� �b���-A0;<1!�����0�Z�c=6�(�ڐ�G�8TI�*��3�E��+��1��i�W��SG�)�Wѝ�Q��x����,�^:���������Q)�,j��������Pr�:}�h@��Q�����u"̷0r#������a�G[�FM\�_BS��n��}+G�N@�p�*2����j4�E�W]��S�������������[.�{���8^��� E}3>"���tV��R�v��~ک�N�D�G[��&�OB�IZ���:�����l� l�{gX�ڐ��GI�z�<R�(��ŧ������n�%�0��I��ݼ�Kc����8_!�ot��g�l�ԊWh)�*g)_j�M>"9"� $=�33}���oz��4����yA*����-��~韑�
tu�j���/�ݏ��} x\u��{*�^��>�ح��9��su4�J�2x�����&&'�j5������b]m�M�����۞��E���R(=|��mx�68�����TOO�_zc�OI��B	���܄[*���9����k�wjh���_�����H����M�q�c ,�4�{��ue�ٰ�'5`��|r��z{Mo=�w�}T�vK�|�@k�ʡ����&��r>�Qxޡ�s'�S�?�_@��i=:'{Ɏ͗����=�u\a>�+�+~�(S�.��k��V�/R)���H���3g��f��3-���/���=ġ��9�X�	��y�:�y�ɺ_�M�6!D/����d���4'0�5/���Г�!��qpI+��脵��u_[�̬mP�7���Qnԅ<M�1�n�>�q�[8��������.�;¸|�ԏuO7&�(�>~��kE�8������7}�fxz�¥�(K<�j*'"Ӌ���^zsѾ���XJHv�1���&i@�Va5̃�֗�qJ[�7��$^;�B�Ƙy�a��+��@>�|hwkHF%����3�s5�ɢg5�+�=.G���P�XnK�9C��u&]��]G���>�ٛZ�\j�3}���-1Z���2����%���(a�;,��6��w%��7n�+pb�`=��; ���2h:����h�;�p�e��.0P�ǉI�"��:�ڴ�	W:d���ع9�!RQx�nq}g�)��sg+y �wn���6�-�Ue�dR�r���ٲ@�f�v���9��!=P8(�X�0*���T��b�F���h�0�c4�t�<rn�u�(��ǈ�XC� ��A|�m�1Z�F�⻭�9�xݩY�����|���-G� c���mryF�}��VpSYLYE�������Y۫.���u� ��fU�	@�U��6�k�J�>��h�٢�N�vV&*	N̕�A�{N!�+����U�L��`DV����ݨ�d�a~�^B���dtJ��3�5��҅��x�;�^�CoYB�Z@K�1].���I�3��DdW�'�,b��V�ج�n�K���(֚2��#Gdj�=�5����f���װ��.�k�腶�ZF.���ٜ_&n����0B/p��g�}y}���/wP̽�q(����&��͒�LR��Z=ܝ�2^�ɐ����ںf�U�(��	��/0�~�+�[��������+��V�W;/6B��^�W���NUݝ����ݮB�3?�n(����!� <ڃt,��Y:�<��� ���	���8�s��P��v����IK�х=ħa5��0uխ��||��{�w-���=���D�a^]e�e-^j���[̚4��m�GfDR�����i� ��`���FIn�.�2h��3]��G��4P���9�-I$��+�U�&���.^��� 2�]�rgY��5��bǹ�	U���,��K�t��"�Y����]���e�-b���r���5��1���P�:�T���\��&^u���b�c�W�d��2+o�Z�\�͙��̨U��38�eޮ7n�K#SQp����܆\�Ҩ�y]��XU����N�9ת���wk-�Z���VoRf������dd��i����]]ԛ�jۧ9"ё��6��"���S�V�F|xV%u�:L��'���O7��lDp�\�ܧH)3]��k&X3C���O$GN�;�q&6\��aC&7#�Q�,.��z���-�j�����y݆(�m]�À2$y�^;��1r)�o2��_%�R�T��o`�豲%�oslb�5�ue4D;�۸'+˽Q��6�����jfuŠ��Y�Ǹ��L�r�@�++
��= �2*��VMF9�+8��z��!��`[��9�{SNc6x����䡅H���z��ݹ|wf,��z'�K��r���T�˜��p����`S��a�GCe듐[M"��Q+����$���H��/Q<�Js�':�$��w\S�h�!��*�,����B=L����;�fTn��K���м��;����S��8N���%'B���^fa�ҏwr)�i^�xA�^(�Yx纅��zG0�etw[���2�����'u��7Rr\��V���{��,���J'G#бs�79J��*�IDGwu'JU��Z��y�I
ЧS�)��5"�U������G$���BtB+�=B��9:Q��k�˨�[��r(/X���K�ٴ�2(���=���ݥI��ʎb*%��8;�<;��ȝYU33�;�Q�Q������xz�գ�åAD�ou]p��Ne�44��88�Y�} �A�wۣ�*5݃��L���9�ڶe��z<�?1�-Fri#�-�����Q�d�>�e�;��z_�^�Z5�k;s2�1d�S��B�t�yL�pL<���1g��kT:����Yt}�[>�q��)qn'X���]���`�(~���z��|ȱ�*��K.��q���p6l*�%��Q���T'AǶC9^�Tv�A�f��(� |��|
_L���m�k���]�Z���2v{%�U�J7^	�k����ew�0��0l��~%�"ʼg���rTWH���
�Ϋ?(�w}�k|&3������~��֟��i5�#*Pg�'Ң4����o7��z��V��5������Z/a�j+Z5i�]�˝�.�O��������L�z�b���O7�_a���_A�"e�¨�.��{���?^�SF��~%���x�F��^V�m�y\��׫��?Jə
<x�Pfa��@��(gЯ�����1���T�{����\��7h۾��2�/ޟ�r�X&#��d�=a�����*g����֨����q9)���&�y��KYr���;X6�b|�GB��"��=̶����Z���[�ȅ\��}�n�;�����aj]P�ble���'��*���� c�RZ[-V��p�!�����Y|�R�fR%_%��R�xub���bfF&]Nh�ʯ_���ꨮƇ)�nx�j�:ԌK�c�ُzS��3U}���q,��={�;�uxp�ܬ�/�'�}�}q�P8iܠ�<�H��'��y����x����}"i&9e/�>��H�\O�S�e�S�'�3��G�Mǝ(ʌ��F��9Yw�]俩�Ϭ̭�g�J��t�;g�*aTOeޜ�%�Q����V?��2!���Mé�;qϪ=�%�=��"�Q\1^f���]&�{'�T����'F*5r��e�V�5�\����²�ћM��y�%#���F������@��
�����4�2��x�~Ls{��KމW7�2}�!����Le�M�_Δ<�'E�s�� ���y���r&���'�T�}C��7�#��Њ��X���F4m}θ=7SAIҢ4�'Q��/Oٻ�~�9��-1z�7S�{PY�&��j"{���/�w����ߑQ�%è%��H�S&&�Ou�����H��r�t�_Lf���ꉩn��qͳ�9�pmE�Da�wP�麉���w�nB�D]ܗj��Ԧ���3}1P^u�A�ݦ�^~�K��⹜�7�ŭ���8L}�\-o����7��/7����F��Ӫ����Uӱ4q���3h��5bh,U�)��V5$��#nR��]�wTs{��d����C���'��77���=�yoc��?��AF������Q�h7e|~�+��F�'��`}Z��>E�2u$�w�<���K�Qk����#ߕ��޺��G�(9|��4zx:�~�P#�n�י�ⷱ�+�hFkTQ�%}Td	t�EB,��0���aD���D+�Tk�=�Yw�6*�?z5�c��}R8s�Ho�&M7,wQbyҐWޞ'`Gi�.�m֏A�g�\�!�T��O���;�)��Q�g<��R5�c@rm00�PQ֤<K|��#��o�xR����:w�r�����^�ܫ���i��k@5��S;�e��L�Yo��uF����k���&���x�7>0�{*���{I�~��kr����k�?J����e�+��F�%�䶷�/�Ո���;�F��c�x~��WG��|�	��O ����FuO���o�k�=��٩v�6�3��v��Xa}n�����T����V�= >�O�;�R����X|�?w:`ۤ��S�w�bk)M��Ľ�3������=F*P��/�����@��\K������S��˯6B1��6>V�����c%v�
���/Qʺ������ITX6�nu>�5!����j��5�,�U����J�o"_ޖT�s��Sֵu�{] r��3���O����ԡ�mOX��Z�ފ̘�N�w���|� 5�F���DzK����3�8Lh:gĝ%�+�\�c��ʘ���]�������G֮k��S��n�ǋO���e�����s��������p�z��M_�އ����$��Q��^��yԋ4�PW{��9��d3�0�-��Z�M���v���}�Sh��f�A�FX�i����9��!5�xA/<[�U����bqy�����0��i�T滋��rY�P@J�~�&K}$_L��`S��I���f����~�ǃ������{\/�s�MsuD4�J�2x����'I��:��Q�~�~�)����t��0��\5?ܲݯ�|�pω}�sc��f����D���2<��И�{2�Vx�[��l�5b5�������?�ݩ�Q�ɂ��� c��`LG$A���K\B���*�mx�R�5?a8>��6T�/�A���+˥��yP�F��X�k��_��6�+
����{�Br>��dɥ0�����p+미����~£]���'��0����hR5}Pk6 F�D�Q��	�kj<���l��\2�t]0�ZP-�t�,�|\��3��q�q!�OMN���*���L4�1VMp�ޅ6��iuEES|'hp�Q��B,t9K�r���9�̛ۭD�F82=�}4�PD5�v�鰚�gߪ��ЊjM�xg�d�c�d�W���"��OwK}oFu�9��C����+�N(}����s^g��}��O�)����<�wLTL�}��]�����~��qx�씫�S@���{q��c���8��e}���;�:�RG�vuC�����n�*�ƍ�^�^yIƸO*�ڙ��xS (����7'�t���y�hީ�XjM��/N���W�p*�y��6���.c�]T�D-�@|oe���,��}<�܇w���Q��W�&-\X��~��ǉB�C�)���_S�N���1�MLT,�>>�(v,8y%�fb��#r'�.n�}^�J��e���g��F�E2A�X>���]+�dR�,ߢ��~䝧��U�Q�v�O)Ǣ��͏&-�����}�3lÊ%D�`H)}2/�[s�g%o�C�do-]|~N"s询wm	/�`�����#Zu����鍄N�G�F~�O��3F>��2��u�#����3ٟ2�|s��x���Z|w���}�#)�c�'�n1�'P����$,Q�j�3LduKr��Z?����R�F��7�3i묬s)q"��q�CUp��5��}G�߽���*��.��M��˷�7�)T��	�(�	'����u��u��xfE��� (��œ�Um�9�,��{�ْiR��&Gg%J�G�n���&"[�.:���C��oZ5p����������+-��K�:�cm��Y�$��̿��� ���J���BR�7����G��ѯ���Y��s��$��!N}��ihw=V�NfG�����P6h)S�X��7�������|RB���>2k��<�0��}E�.�����.����'T������c!g�f��z�lF˜}����X�5!}#���b�먮Ƈ)����v�j��2/��*c��N��A��V��5�~	�Y�|z��ۍ��V�e1q��փ>�j��N�v�]FO���c�G��Y�����t��?	E�-N�rp��g���w�'�3��y����ߣ-`���{}�	C�~��k���N�`��U���u�u��'̟7=E��b��>e�p�s��b���}�6B�Ɣ��-��8�'r��T�BgG�6����d�����͠���5ǈ��w=������e}����3~j�a^ڜ(2=�g��gO
���4�����e����{r�=�+G�Nh�o��m�lmZ�*a,����o�o�m�ZV��=	7�����k^wVf���=N��t���ե^U�ջ������P�`�.+�U/��:餮X�]#��.�e�z��3�e��*�K��F�@��h�oG}e�v�i���#�q������e�M�_��C���1Q�����<?�A�L{��������5�gzSk�;��Fhr?��G_�u����.1�;j9���jtz�.J4�$����J�HѕU�Ӯ��*��0*6����,�&��j{��9�n1�;M[�#*9.wMªu=>�ȥ^}�|M� wK�����5�{�\g+�S�\M�~��#��?�i�{��ß��"���ݤ�p��z>�fj>��"�~�&[��1<��(j���cW�����t�{��ַ�K�~.wI��zꙑ^S%}"L7�����SB������s����������ھ��CR��r9ǻkÅ�o�Y�.o�놢�Lr� /�<N�1�	�0�{SF���N������9��>���٧�\:�5�Hb��R|�.�X�,Ls� ��<N�Giߥ!>��*�OV��ɮ�/2��"6����Q�>��ŷʑ�ƀ�M�K��T�R��Qu�;ݟ=X������~��~:�gűկ=�9��kN�߽Ϋ��;Z�N:�9�,>��.N)vI+"o^_oN�)#���^F�Nu0�D��n���vo&���wu\hm
��_P����h�[�=Y%wtU�[P�VX��W,(��r����]�<č�mj}�裙��+���ֺv�^��uW@=.Ia�����܂�#�2�g-K���aX�������.�:n3g��^P��=,]�*F���,�Oì$��T'���_]���zv���#���~�37GT��N�ypg�Jb����U��곉����:Y�n9���L/�ڜ5�������k���u@B��t����w>�n`v?�+}\̎\��t�3�p�3ؠy1�,x��
�a�&5��銩���V���ssѮ:��^�u�uB:�tC���s���N�ۈ�Z˲�i�,%�\l��qn*�IG�IG�̯���g���^H5��Q��>{%���Pߦ�rcn����{|�k^z<�S�h�P�N��~�;T�=ԋ4�T'������3�F��r�@����ݫ�+/�\>�6˿`�J*2���|f��[,dk��z�����R�&�S�p��v2-(��w�>��W�=�ug�\����w�J	Q����-��q�+�;+6����߶njW/�W$�'��׆��.]�p��I�������	eh 7Bx��Dw9l�?n��-d����h�T�fV���]�Nr �,���g*�0��x���DL8��j�8���@Rk5ђvXR��6�7@k���zU�)����/sw�Ǔ����R�^� �Q��v��88섖�+���-ڍN�XnĬϳw�:��8�P(/����PG^�]}�"�D{�W���K���M>�GS���,����7fm뜙�|�l�Q���I9��תxd�mG3_7�FTwz�<��x|㕁�*9�M�ܳS�/}8w��(O���S�lgԽ�o~2�ǽ=���T;�$�vO�(�������X>�{7o��_}�b��y2iL2��%��luB��:/��b�3S�_k���T܌чA6��8�G�^g���К>����V���f�F%�1ޡ�T���I�'�]�?|�o�^E����	wyYr;m+{����5�{\�wج ���ٯ�ʃ1�M��v����A2��##aZ��O�k�����n|��|���9�y��5Ct��dW�<Ne'q�%�߲�s����g���O*��Цy��������_�S��jb�'~���W���Qp�}�_�kV������P������Vʀ��c�N�R��wP�Z&���˿�&�|�E���\�ܜNI:�g���3��#i&�*�<k��zZ`߮o�-��ݝ��z�ǐ�3O7��x��Bo���h%;�Fn��t�����P�G�0u(��=���р�pY�F��복h��qY*
���%��>�AR|�K��n^�S���DW=&��˶g_��ҁ&4�[��_R����'��^(n;˰�2�?��0��>�q�\u�(ݹ �x�ȱ��J�㖲�-�Q�O7~������Z�8�K�mxh�����G�>�z
f;EIF�����$��,㢽�QQ]����P�k[s�wP]��g	�o�ѐ�����F�0�D<^���(�Rx���ұK��~�����h ����[2�^dqQ�9��'�-��.Z~;�pa>��_4�MP�,���.���v��R��.H)���Z?l9�E{Z5i�m�����:~��z��2����R��+��B��4�I_�S����D�%��*�]4xnx�3X�Tm}��4vj��9�M3s�����ŭ"|F�u�`OJ�
<x�׌�/���s�X�q��T��?�����̻$��e��"�F�j���s��e���X.���ǉس�%م�ֻ8}U���6>����}!N �+U�����6���p��uHWcC���ܰv�X(k��t�~P2a���b����gor{��L�}YkNz��Zԯ�������~7��e{�p�Ak�"��v{�]h��n�VTܻ�F$-7M&���.v`T6_]�;|:��*C[	(�䙛��G�_3q���g5VS��xH��2�;+jG��kdǚt��*��8ω���pSt��w�ս�l���>��+\5�߀Ÿj���b	՘��!c2J�O������B��7�H�h�WN��{�?��`aܗI	�!���c���ۡ�f�~�BE��ϑ�;��#�j��^."�n<5�}v�K��Υ�T�\S5�m�p㏞�kE��pkq�r�Gd81�B�ڕ�{NUќ0j65��q�B�9��oqkR4;N��9
]�����ukڏ>X��<�mb�ι�3C�9gT��qP]�)�� �m�\/7)ِdP���Q�8E��e2��7{B�+x��_84kWtM>[B��8|��7��1v%Lub���!i�������x��{���Y�t궉oNՉ�w����}aJM6L�}����;����Q[n��L ��k���U`��֝�ɠ�S��g3�-:+lǊWj���"^�yZ�H�,挛Lq��i��7V�4)��.c4澹�N�w3���b5RG|� 9�s�Y+/b��ΖU��q������� �i���|d�p�z��B��:J�����ڀ�c�š�.]�z��)h�_b�i:��]y��^�V8��϶���}y��<��U��JV�����A�Wf^���Ev)�i=�J�:ņ����q��f�^�b��2�Ħ���b�:O
Ý��J�O��g.�β8i���&��a�0������{%t̤Dd�����}f聁��-�<M��s���˦	Jl��ǒ���"
��}��qՕ!E�.�eܠ�(�Y�k�h�y������n$�V�tl�W5�)˽��	��N+jNmdi�T�T,�bs�rn���r[ˉGo(+ ���ƃ2�&Su��E�2d��1;��쭗����m)����i��C��j�̹�Ws@X���
L����I+�=
w72��Er!�0u�.�t&��/���%mk��=�'��'t(�u���w^Ac6�%��Vg��{j�\��3gRu&��GV�h��Ӷ�P��9����«S��q�ϲC-�ї>��j��_;�R��o���@z��Q�9��iż����Ӝ\�}3D�±XZl��6¾9�@�����u2�۵6w�1��!q�y��͎@�J��uqB-	����w9�"��A�6�-� ��Ķ9���s�n��;@Z�W���9٧�v�:��u ]�B�k�V�V^D�+�'�{�RdS����a��Uj�#��1�y���:8ϝ�W�� TTI1v�����m^u��@x��-�ҹe��P�A�XK(B�\qi���9�o7�gV�U£0�$�j��!��#�oV9M;�:I��[Ē�S"&6�rQ����.��t����ۼ��ZJH���W��T�Y��Zz����]�X���ؑ
�z;�;�^n[�b'"u$�(�t�u�+��y�#�'B�vkHN%������r�wY���;���r��=���]���"*sn���Ge����\�$;��UF�n�*��R$���=�y�yKB�ֺ%W%C:uC��7p���,�s��79e����"��ˮ���Js1����H��瓸*����ʹz��NC���.j�Z*��X�E�K-H<��c�n����ҏ7p�M�n�wV��zuq��#���ii�͊*.R	;��C�I����8�H2�%�T��JC!<�2�w$*!6D�hU�4
�H�C�**TL�ӕg��̈́W)u<�u̈́DJE)�N�!����ȼ��P��B ��B#�d�et*��G,Yܬ(�B��B�9m
�jW-H�I,*9�Z҉6�R�(IdF�0YG�f���(����G�HQ�@��6ܷ��tOx�}�	�uؓ��l�s��*:�e5�)�B�gkӲ�N�j�%�.l�I�ؕ9|Ѕ���a�h���X�s��Ki��>����u)<�nW�����3�j<�oΔ^�u��ދ��4�S��Fl䜵,;e���J���g̟9=}ϩ�q�y��W�)��B����߅�e�4�}�_��w	g�g\΍��N���2�L�Wi��er�	c�!�#�1�&�w�y?!��{���n&��uz�v�_�+�S����FxZt𭤚=��uO����
�vn�����8�uPwy0E[��e�sM�[�����i�mL��Q�N�1̋���ݖ�X�����ׅ���k��)ڃԻ��w�jǞ�|r��h�k��蚝�'�oµ�.�y�i�g�����ǠO�uh�������-��n�ӑ�9��@zTgʈ�א:���g�[T��o�g�]	�ρ�u��w�X��|���F����S�\M��ZG"ӌ�K�~ϰ�	��2��=C�<��QqM35diA����-��e�X��s�޵Htd+̧PnyG3Q�G�/31o]�5��S��'c��9M&d.�-M����Q%|���+�Q��gs`����vTJ	}W�R���8�1sc����Е���7y���ѭs�*�W�y Y=�U�w^��_:��k��۴�9��kk�S�6��#vD0�L�k	�����q6�YF�ݞ��3���0)5�����sk�G�H8�{P�J9P�ͬV_G��s�Y�&�3�����"�|\��b�t��x���y�	�0n���5�}�)b}��4��w�5�,<~R8?��R�ɒ���q��S �)d��F��
�~ߑ�0�U��0��kt�Ծ:�v��j7���*F���9St���;X�e��C�ͦd}s��-C���Q?P8;������u�}�"�Z?#���7�yp���v�>��k��gs���Z�2��ykq���z���{e�:���uK�t�oK��vڸ���ğ�����o~�gW}H���_�������5�fpߑ�����?�Z=6�Όk��2ׯ<I�⛤w>	%|[��!����9]k<���Y�3�Ӱ�'tw�~E��}�]Eqjw$�>`{+�w�����+�Q|뙑}\�:M����o�t+�S����/y�`֙�
����G��Ţ���i#�-����u���"�O7;��0�ӯ6�֋����s��X^�.uN'�%}#~��If�%�k�UG��]y x�guTv�.Ϟ�g��C~��(M�Ւ�/����ܮԥZÎ��Z�)ʳ,����-���I<O��F�I����QƁjc�^:�YonN��hMO�Ӷ�h�0 ��L��6�j,t���t��돰�X2�l���1��]�gb�ul���i��p��5��wyI�o�~:��D�K�Q3�L�_F��,\Fu"̷(NDw�����`���@�,JZy�׶�n��]#�׍\>�} �(�B�ʼe�!J������5-�{;��976W֔�Q��	�W_	�����F��Ͼ�;U3�\�k�	Q���-������d�U�F�3�g65�eθ:;^=�K}\,�����6ڃgbj&��,����ĕW���v�k:>�c��h�G\�_o���z�H�~O�la��D����ɿ������c�v�x�$�Y({!>�ivM�dW�Iڹ"�qo��f��Q���h��ͯ��� c���"\�f�kݗ/��|�ɕ<K�3<�M�=���Z�;F�ޞӼ�Co�#�f6�ϊ�W>�s/���"Qo�}֐�.�J��}*����R��:'{Ɋ��OI45�vQ�ч2%�3�]����\&��@뚓qz���ĸ����TJO�Wn�[z���NM���;k�%�(/�j�1~i���3��=�}�P>��a����Qx�ʃ1�ctc�eU��as��Y��ͭT��k�&�ãF3I��uwQ5Q�N1X����rƭ7����B��Y�q�!oI�"��iIL8��\�ïj�1@���1�ub��l���Q�sjr	�}�-7+�kE�;�۩Gq�v%�,fw_L��3Kt�+�A��=L����rN���5�{�P�9gŻR-�~�uU;�{v܎�R𝿠�v��{��EL��=q�0����_T�rn(�ٿ>^���.��َ3^�JS���9'n�co�.ʃ:�ښH�-�����-��ƙ4ܿ��;>�%ۡtl�X)|qC:�Z��M������ܜ�9$��jΎ�2��|�����q]W��fݲ�^��f������7��C�|f���ed��e�0ȱq�J���&���u-v������1�g.P���S/�p��hq���l�3B����d�(3�]֗�f80K�x|�z�C�3��q��_&�D��{�`��<O��5��k��t�:u(�LO�o�ס����Թv(�@��� �Ȏ����b��o_ʢj%�_�����Foe�NM��񼁝����K��>��9�\�3�\�۰G#zѨ�����ޖ�q�Y��������=�΁����\gĒ�;��8��/�B�]4xv�2�7�Tn�Fߓ����S���ܶ�Qٱ����a��;����jG�����2��ȼ��Z�k>P>;�j��o���@>۩��%lζ���b�$����*]���,��hY��\�$]����"�@�Tz,���詻�f��1��D �X�V�E|G6ht��GC-��a�֑f��x��Ͳ_M�zfG�x�3u��e
�_/i��	��^��~��P�����ҩ�������F���p5�r�'eђW��f;r�1?!���X�Dc��W�ϧ�t�4���ݖ3��p�i!��hr��僵�a�jAY<K�]�/���.��o�ޅpR0��M;�9��~[������꯼n;Z�^:�t�;����_��-.�w^xg��~�'6<�A�P�+��pT����=<���c��'�3��G�Ja��IlaE��	:�}�Y�y�]xy��W��Ôz��8:���6�|��z�|��{�%�n%H�4���6]�d���v���z�<�J�.�pW��9_L�&tz��N��=!����>�"WZTQ{�����8�t�,��l��W�7o���S���/�xZ�gO��=R/�d�U���ڜ�
������t�ތ-0E�s���6}q�����i��>7Y'�N:��'��PʝZ��x}g�3I��%��u�Pz�w]�ՏC�/�^4m}θ=7S���l�Bؼ��@v�U�Ї7q�t����]�V��1�]�e� ��)Z���g~�StP��q�,��{,'pK�.!.�9w;��U'����X�b}��+C�\<�8�qS��P�ӧsj�^J�Ed/�j�\[.�n;�s궱��uN����x�����FI@��R������uTj{Q5=��ߜ�ӷ���
e�m;�]{f��uo=\+��UH;�l�P���An��l���r7��ꉩn��Q��nd�N�\��f��n���aڋn����2�d*="�'�"e��x�c��Fۏ�>��vn1��ٚ�ޡx�s��q�.���9��}���i3!t��MASѲEğ?Jf���m�S�z;t���zxu}�?T���w��[�C5�����?G.R�^&0�w�_����=�/5���~]�lÜ���+���\o��_T�+��T�y�d�X�,Ls� ��յ�C�X��ߪ�'&㧵5?a9�27����圈Y=�j�v�����b��H�v4*��`i~�)b�wESYq�r���y�p�T�^�,�^�l��]_Wi��h���������=��?����%��O9;t�K�j�u�
4���}<*�
�Άg+ᚮ�'�{z_��_Ρ8����+F�6'{�{ެ>���V�c>旙}�T^�Y�����G㳷3��CgC�������1�Q�����&4����*mV�5)�j٪��J�|��Wi5��n��՞�����4jw�)Z�mbY�î�G�J�Uz$n�G(�R����C�	N��U�6��N�,s��f�c�v�M$�w��@��eθ�����86_��4���v�yX���*�	�ZS�}��G�?��~��w�����L[��9<NeD���c�d��v�]����GCOUq�<��
��3#�4��t�;qԼ7M�\�W����-U��i�����ԣ�'�f�j:��uH��Z�CHGXm���s�������z,n���˜ɾ�[�y�t�Hڈ�d�+�-�}1ڌ�{����G{KO��K=��̢wW�o��	��Z��M��������pV���	=S<���{���E��ڡ=#z'�c�"yx��J��ǯ;O�h�͑���#�3�p�e�@6
4���,	��|f㌶X�͚��϶�wn��Q���_�up��n�0\y���r0�}m�����v.K5���De�~�_j��/�~7�Ύ[ŝ�!��[��g��сķ��˽��s[��[u|�Q+��WDҙ�;�&t�Ϸ��(`n��(��j�떋��9޵�4Z;c�R'���p2~f�5hR�_k'�b|���_�:O(�ds5��"e�h�z��u_�Q�־*7�ɣ�mx�p�u��*�C�G�:��(>��P���7�@t���t�	W�Nd��sB�A�U$���%��$��!'�[�o&�<�WCnf�]v�l�̺��lc���n��w�!Ӑ�dtZr�Vua�A��F�>ɤ�	�]+e^刭r�&Z w8�`9�&|x���k�鰢'��U�R���J_�m�Ҿ���&M�����,�rG4��E����]̟���s�h9��W�踅��b��5,�V�G�p�9U�������/���~�tu�� u�I���f�a�Z1ޡ�M��u�/��;������׼�;q��u��V/�?\\Fs^g��j��F+/��M�M�] ���5�ޱu��F��*���qU���U��F�`
�ϕ��լʇ�/���X�9�<[�i,��/#���+��������^-T;�-��jg�=�Xo�;�q�<ܛt�;g��ߗ�����e��[���kd����£:rN��'�ۉ����B���wF�\����@u@ƙ7�D�'+S��g^������2���\w}��{:rN��$�����Ύ��I���o#��5�'���g���6�k�^�K.Ϣ9�g��>���H�F����`�c]�+{�A��g��lởf�eݵ��z��_B|�N�L`�|-��;\�����f:�\�i�*;�횛�����Gj��JR�>��olK�<RQ1���՘k;%���p�$��LQZ̓�Tm�fS��Ƚw�bǷ��o5�FvEL��ۓZ��U����&c�aY��C�,��3:vR�b[��b�镘�f��,���]�e��	M�h$������:����~Nr5�A��w�ED�:�q���F�0�C��8zza��j?W�7�V���}[�(_?F�挰�5���3�{0r���ꉨ��~�~;�pa/ݣ�:e�y8�}0wս]�.�L�?}2T� 6h�$L�\�h��G#zѨ����V �wB�'��mѴ~�����\�3^S$������D�K���WM���p�8�啤�}�R��.-������'���K�V�����x�c��VD��(/��^x���;߱?*K�.�9�|�.>��i��ԆߒF6#ϝi�p5�r�_��]q�1�U�ͰF��5��N�k=���?��z�b�]��7SZ�p��T�}���4ܰw�BFuL�x�>��T=�:����vN��7���<�Ͼ^��~��2զy��o�����:�t�U�z͓f����E��5�9;-H���v�	���P�*��GK�x�/��m_�����nCg�v;�|��f�X��/���JTe�f�����Q�.pu*˾9S+�Q\�1���'ኜ��4;��ڶ��N�v�һږ�V�s��(���l���
�܇r�H� ��c�:c[�e�d�3�:��>�e)x����^R��5�hp'���(��&��º�ja���>�f��J�����e�.:�s:fZ�wi�f����_>�N�����z�'@=I�������}Q�_��Qe��2l�D��tz��N����5U�k̍�̝��;���=��L�������˙`�Γgn:�Q�|��^ڜ5G�~�<.�����.r��^�x�ԗ#K�=��a�8x��g��x=i��ڟ�ÿ����kb�_���C+|P�2�܉���Fhy|}殺�[���/�c�;=��k2�V��_g��tG��J����^����_�Q��z�����7�Q=���/�|�n��f/��$�;F��Z�01���Dm��0��U) |��K���-����#�O�q)��`:8\.-tgx��,�ޗ�#�F��茧+���� "�~�&[����������ke�t���/ȸ��᥵�c����\�\�Aʆ�2GL���1�QQ��7��+�]�����(y\�c����E�{�Lp��~��f���Qp:zd
����M��܂9�	�y#=��n1=fl��d��y�UZ�73!�5L���T���6m��ll��c6��66m�c`���6��l����1����������o�6���6m���1��ll�F������l��1�cm�1��o��6m���1��������6��������PVI��JlD�����` �������^���UEJ�UB��T��PU*D*�U*��*�A*T�*�@%J���T��$JRRR���U*� *����G�*���PR�(�(����v;�%	WZ� (��*T�ETB������UE!kDJQ(�+Xۡ�5��)"J�%U*AJ(�I�UTJ"T*�**QB��(%J��*��J�D�J�E���E*%)
�P$�R�HT��E+�  Lw���[S����%*�;���l`���N�]eӺ�e��Z�WZw[57C��d��wnST����Uf�9��h�:5v+X�wJT RBv�)(��׀  {Ъz�e�[�p�̣�����tV����rpQE4Q��� 4� <b�4tGi  h  ���(
 ( î�����F����R{5U"[b)M����O^   9� ���We�zL��enk3�������g��u�a;QQ��=�^�[*�{�ֆ�ծ��KE�,4�]�h�L���Wm�%*!R*I�V��  ���mUs���t�9UT�ꛥvn�U��9j����P飗2��$���e��u�j(�һ�vjw([u��*�D�TJ�T�Qlh"7�  g���:�w\�
Kj����]16�v]nCu��v�W7]�[uv��]Vr)Z˹��6�mv\�\t�;:�A�U�m�-���n�sjkmi�GiR�R6�UT�"�C�  w��R�m�ەYԕPҚ���mbYJs��m�Y���n�II3�f��e�U�U��mmrS�v�SY6�r�:��g6����gDvw+$��JH�J��H�  ����j��[���՝���v�#�v�-r��i�+��YY��nY�J�ݶs��.��[]��jT��9��u��'�Snu�.˺v��볝�r"QID�	A���    ؽ�4�5)[���ꥻ��:�ɲ�vSw]ݚ�!Lr���b��p�ve;��s�۱$6eq��wF�ݻ\b�u�k�wX�Mٚ*��2�֚��R��	J"IT�   6���k��us�gn��s�����kv�fu��u�C'uU�Z��m-wsE۴���mnV�-���U7�v���6���U9Y�d.r��[#�U)PH
���T���  0�V�qΕ]��Wwsr]��۶&�-N�l�v��ep3�%��eۆs��r�Rs��,��A�vv�Ԯ�m�sV�Gk�e:j%����j8��� 5Oh�l�J�L���$�E  T��OP  E?�P� �?"c*�� �	4�=U"��zjM���B�&z��2���p�����Q�P�{�}�gﵭ��׾y���_�	!I����$�@$$?�B��P$�	'�!$ I@$$;�����~�3���~Z��f-��!�W����H)��(�1�+hn���Z^������.�N-���.�`Al��"���S��iG0m�V�t7�p]�.��ܨ�UEW@��f^�0�	{vu ��d�MV%M���LM�i�p֓�-�ifQ��'t�&ja7WWlG�^Y�iZnim��	��YqܣiPp)GG�C(�ɛs.�#��  ��W�R�e���%e��X-L�ŶWY�$����h`%-5i�r�n�{��oVT�Q
;+��̱��b	
�Q���ky���H����-�L5y���ҋ�Q��:vv�U\�!m�amH��y�z6�7����.KMd2v��Ͱ݌Y���`���ɣ6��n��nc2�XR	U�,��Qd1�eXi���ea�Tpaتµn�f�W�ض�� �V���1�v\K�0�j��Bn�{d5�����f�Y"��eހIf�O/rEWF��۵a�J�VfCZ�hc��Y��m+��� 2�,��jZ�U7nָ�Yu���VV:u!��E9{kq�v�y��SG1�:�5�H��{�H'V�a]���Z�*2�R��c��5Uى[ugjnFI�ƨN]nj�	&0LMd���d��ζj+*�9�٦l�j�\i�N�ݻ�+f�%��̻��ږ�Y��G&�h�.Fj�^l�i���X e\-mk��QT����5	q�k~ P�����K]�n�!u�iX@*C���Yyi��t&������W(]h.�����x�q����/Y�N�l�q����W�1cy��dX����P��S�J]F�����D��PEC����0y��0k��]�\E�Z&�W��#@к���ԑe�˃i	*�`1Zjj
���t��yl�S��(��j�(��Lk�
��P90����ע�`��Pѕ�dɢ�{tb� ����9�a�[+L�wCrXض8�V(��fM���j�v���;I���K��T���[d��C6���Dh��pe`�wV��0�V��X�QŁ�����bo	Q,aޡrv��Z)�$�cG]�[��Y˲ �^eBCT��fm�g�%n��7�,��!�Ä[)�d1���v]�v+m%%)e��� �Ѫ�"�q��2K�M؛[�E��$6�
Zӥh]��E��T�� � �mk��YxcN◺�FRћF�ٷ��غ��հ -�5`U��2��4���!j:�J�n��i5��t�d�{V�왘b��1}�E9$iD�Y�f��\dwu��F��ׂ�C-P�h�w��XU+�6��FcIz�X��LK¾�`HX������Yk�5"�ȬK��`v�f՗/5=B�ĕc�e�ƫm�Kl�u���o�;��1(�g�ͺ�"'q�T�CH�XWy�ph��o0-�d�b�]"�ctF�	ݭz�`z��2��wŚ7#?^�9(�E��j�U����E���_��P[�+E�L7	!�KV��W���n��l6Ց�27W� :�:���M�u��[��h,7%l���J�0ْ�p��n>�2�k7T�7q���e����+%��W-k�j�hJ-o�{��
X�BS��%\�E����V2��LM��E��ӆ����[��U�P"�j�ږf���
�i*��w�6���m�],�$vY�����Ď�k��\בݔ�MKsV��M�9��̩����c�;�7�a��ֵ�%�3[ʹ �0�6b
�KG��B�L��hKwJ��(�[��%�N�wP7D�vv��I���H�bU����=ڛak"f#jb�V��Q	*f�u-eG���D������S�[�m�r�Z�Esq�4��Ѫ�:AT�+E��s�/f�K�!	��/�#d2�K��unS�D~���f��2��&�(�y�d�������h���DXˑ�6*!���AVe��Sܧ���
e��d���*��7{�M�Պ�L�M���J��lg)L�����å��н'o/'�VS���X-���0�r%p�9����Su�LP����F��@�[B��CCJ��hVe��c��9�bxcC� ���3l�=���z�Hi�Ma�u����J�t�tg#���m���9yL�lR�ګ�*��V�)YW �Cb���$ɰ�ܕtݻ4D�ZH���o(�F�}0 �I��"�+3�6���Q�6)��� ׵�ur5�J��	�ffC*Rz�a���v3���)��7�̣�b��{fC++#�
tsvȘ-�4�ri��b�e3HE�n���,)n�F�Oh�E<�ڽ��;ԅ���50�wp��l����92��M`ӯ@b��h#2�NGACz��!CNk�
���M9�@T�+]qTo�y���<�VJ�4�[��+�by�&@��&K�thIy�i�����H����81�ʵ(4ӎ���m���-K�^L�hC�M����϶�.��@�l	T��kj��mŴ���KNj�kOh&$�Z�l��kd٬1
эKͶ��*%k^-�1Yx����E�Qv�v�+!t��0�F�ܶ� �`D�܆�^�	�����ll�"�U��+T�͒�p�Mv�n8�f��;��G��]4�A���4S3\Yfޅ�G1�N��y�»P�t���D�K%�m��� �rh�5a�0��	��h"AJ�Jc�$ 6�X%,5��cѹ���(���[&�B��S��k�/j�Sj �Ê7JK�3i2Q;K17��{[1V��Ĵ���U�[�s��n-���mc�׳�
4�b�h�;�E��@b7%��M�&�5h�7
H���F1-0����W��8�7 ��퀕����ս��[�HB@Ś��<̚���R���a��2�b�U�Xm=�4\M̥i�5�^@�l�J7��g�ɳXHvH���f�n�^!X�����"����<6,a���)�X�B05�+	�n����%+^l�Z�w(�VX:��$/B ��[4��k�u���o�C6���Gh���VP`*۹�V����a���kT�&���L���9��ܕ���Ao1���HC�G�X���%���z����a�n�[�YGU��]�R�3�tRZ�cT̫PTӪ�Tu� 9&j������ز�)�'���
��0�`�FV=�j1ec#1�WSô��n��Wq=a �c�ݼW��j��w�e
�Գ6�L�l�6�������r��e�XDʺAؔ�tӋm�Pko���.��	3~V�L5�H�e��š�#�(Y4Q�V��]�Nn�ɸ2�'
.a��
ɢ�,R(��.��6j �F�*���Y`ȣF�!6L��-f���q�]6v��x3i�c�ig#��<���N�^ҏUn�i����G5�WcrM��;���u,��Y�&� 4�t;�W�nU䥐^m%Pkxj#�Z��,��R�u5��zC��q�
��t~j��X���kv���]�v�ܖ�����ur�`�b5��%�B�}j�Uj�[1�:Xq�U����t>ʄP�ٺ)-еr�f�EZ�:͗ie����J��sU�������̢�!70�Z����Q�b0�rk[��	�l�N�ӭ��ì��)V+#o[����!`*gȾ��:�:i���l���Z�%h���# dZ�6e���t2غ��T�?�SS)��˫�r��#֘p(�VSu:`�Kz�!+nm���� �Ҟ̐T�S�u�����F*j �v�r�sCT�-�8*�+bZ/c����b|���+h���I��f<т��\����hw
���ѕlb߂�lD���� ���:u]a�q��������MkyN�H5X�а�芼IdP���[2��gs>�-�.�8(�����e\;���"�HmE����ad�_:� %���\�Y�a7T�s�u�V���|cP�Wjw�%��e�i�4���u{��z�6v�k(K��9�@�&#�Z�Y�����[jZA3E`F�1�̢f��ar���aů[/ujQ�ˉT�iEʳ�NT��4T��n!v�c�`1qcB���Z��^Wq�P�� �b�W(OP����M����fG�'����V@/ ��Y��h�.�U�V��ʙ��:�V|�ͽ60��E�i�2��K���-AI��ٲ�R{�N�XǏޫ��ܠ�ͅv����r�R��kQ�˺V����^Bl!�^�q���ΒK˳W��\�s�,�6�y/�N��[6�P����Pe����J܉��&�{&�1k$��E|�[Zɉ�Xò��@�7A&kE�f�ج䭸�ilVkU�-b��iî�]�Q��d�+������Z����+�E�`���ݳ[2���"��_6��ˀ��PL&D����h��f��m�ub`�0�;�T�emZэ�
��UXi�An��N����:�'bH��-�3�ˈM	O!%���݋n����*=z��,��h	y�c04$ �ݱNDg�ޱ2:��B��x���Sf���&.�䡿e�B?�f��ŕ����D�3kC�,R
cU?�!�KaWzF,���݋V�t�)��B����ٗF|37#Gp&�l%�$��>�f�P�&����2����f蔠&�V9zP���y�u�(����D��4��X��JÝK�4��=�۷f�oKB��hc�q'���[{���rA�)�A���d˰��hB�Ø�cTň��7J�U�4e�/N*,@�J�m˟S��`�mрP��)9�.˷v�:;�(�R!F�LP �l�k]L�K]Θ�xTr,R0$��]0�;Ք^�y{���e$K�d��U�MJb���ʗGZ�dٗ��" ��9Vt֙6��E���@��cp��n�ڽZ)��`(��̓V��5p�7&V�Z(Z���E�-�)�$2 �^�����>d�7oVa��D��1��^�vA�cUj�e&�6�q��c��Uma�*T�<إ,Jd��wr�T��խ���)咴ZP�M�[�	f�N���h䨮�=iIM�*�����X��ϯEH�ϖ�v]�ۑ^�5�Z�b̩��e-�H`�wIAFA�b�#���1��E��ݸkr�D������t^ê��o!T�^:sIt2\�p��Ԇ��2�Р�Ƌ9�%tR��jD,�H�зa3n�ψ6Vf+�DWB5KM6�`��)�F�k`�,GV�� �4�a�BW�ɷj�o*�]ʚ>)�aCuZ�γ,U��9�eKF�Y�HhǸa�w>���'��*V�X�%m��Z�.2��U��f��7*Z���x�9[sb�g^����b�[d�ˈm�چ$��55��Ab�=�*�Le��Y�s䖻�u�^����bn��VeG��N��ԺSn�U��6��L��i�ʬ	�K �j�Բ�UD��ؐ��g��+�wR*�.�u]YI���Sٸ��ف��2V�h�f�X�>�&J��nm&5���^����Y'Z�0�N��)���m�
&���a�Um�H��#/
V��e�gpH�6ճkfQ7
�
+A�"�������]n$WJ��H��*�PY���V��%5E6�Na[���"ًSC*9�h�q�Һt)}��W��.���Iv,ʭ������2��y �6�oV��8�"m ����H ��b֨i���/
�Gc��V��`Z0^=4�,�S����T�[����S̙Wyv��n�=R��XwY��ڏ6�efZ�V��&DY� ߢ'�`�`�v�ˡ*�ش��_k^a�ئ7�g79F����.����䛲��;6�d2�b�@cg5��[qG��/2�O��"ͣmک�+�!nk-:T��+֬!�Pt�wD��7j�����1�ܣ�uw�I.d}��-�(2�b1|%f�ϋ�[R3�3�8���E���*b��&f��e�� ���[�	��]Y�STCj���o�Pfj�l�O(){���!w%@U����Iށ��gpǬ���a��*b#�tX�H�){���ٲ�i��P]�j���t��b�(<*U�V	�FS�M����Ŋ�c�lMy6�a	a�zܖ6�2�S5�4;J�ѾaQ��>̊�R�v3j�K���b�����P"�9t�*p^:r�"	�2Q���jc5�+!��[�,]e�1)�5ӫL�t/�]djxٺ�AQ!�(����'ֶh=�q����34� ���y�t-��;�O�-��Y,�`*� �F!͹o��b�D�	o
ZfQr p�)��&��T0��6e�2]��F-9�L)@�g�棑�>�*M]*�Z�V`�]
��.[-���:Uo,���J,
���J�tf䢶U�,�D�N�p�ǈ������Zn�M��4�)}�����U y�����mj��7/0!��*��ĭ���>Bk��Q:L�����q����Z��m]^b�f^`@����:���\�mKg`��f��3EZm5X������1r޵d���a=�P�w�/e��n��7t�����Ҁ+���ط�ӈ��h���^�e*�[F����U�ݦ�`P�C0�q�m^&u���K6�%\AV���"¦��.�PZ�ɡe��GV6�ʰD��j�ݎ��˰�&�@؎����ۺ�hڡcUbY��P����%)l��S2�*ܭ�q�l;wq�@%j�d
6-ևl���L��F��:voU��Dku�w�R\��|�L��s�.�y ]�MT����W5�Q]JG/�F��<���gIks�"$��j��2�>w��_f�6�%��{�l��B�&��m��-e``Gq�cv�MJw����΃,<�_C�8�`�j`,�p�Q��St.�VQ}t��-�]&a5S�]Kw��%�3�.�4�QlR�8�D/�tF����ouY�V�C5�~�{$έ҃���W>����F�L&���Bh1�g\霊�v�J�7�e��keu&'n��K����kn��<9"��U��+{5�.[뮸��Ő�S����R>���pa
k���J����`��-�����k���'Z��r w��T�"߱���O�ra�[�-�
�fW)/��%r���6Wfa�N�hy�TJ�LZޛv�-�2�`4�Ļz���G�қ��1��r�a�즾���<U2e�\܉�8��]!��� �e���Ox�����(���7Y�m��xBT���;���b�a`'�"� �ݮ���m�	�ѝ'j�1c嶺�m����w2LYGP�f�)��q&�k���YyQ�;����|(�����Re
i#k3U��&2� �t�w�[��Fuq�;b�ޮ���u�S�]:F�[K�ߙ��U6vE�����Ѻ�ս� +c�TyCk�1ƞ��0ҡGV7�`�yv��Ha%�r����f�hot��i_y��U�u��G����:u)o��U�X�܋ģ�Z���9��l������bI+�7.J�wغ�2�J�N��*Di�#E����l�i�u�]�u�$�r�%Y�Е�N���[4ȉW���ʜó���\�em�5e�k4�V+������O-t����F�v�\8J��R����K�}�-V�;�꥗�7(E[��M5X�̖�r������ɫ��^@�B��M[�'�k7G}���)՚wu:y9�i³@�l���c�U�vQ�>��m����}s� ��_[9��[�guY	ud���Ȯ���3��3���}�>�������a�ݭ\�yd{��F�_W-Y�tƛ����w�!��1��:n��]�+ \�!Ѣ=��'��/�����p�}W�V�}V7�����ɬ
���!w;�'|��� "�6��w(;0�v��ް^��Y�Gt<yn)Y&3�$�mNʻ��.R�j���n�]u��y���ikL���ї܁�>B�jJ��L�� �p@�*��Z��[t%�i�E�8�;���/5�H]E�,�]˔�XO�����O^�%������h,뷯:>�u�ky#(��]���=N�U��+�[�1��<��胴������&�;�$�����E��	���˻#�) �K�U�y�/yY�e��3$�	�+�ų���+@�m( ��]F�Z�"�b�]�k�ٶ��WR�B��W,���
$��`�Q�ل*ī�U.�w�`42A3��b[�1���,�D]`U��� ;*�k	5-.���4��j�M7(�Gb����#�;�4�uy�ݫ6����J�D;ʼ�x'})f�6${-���Bvh~�{(q׷wz��m�ܔ��C�xɱ9�)-X���*��r�F�c� ���$�1:D0s+F�����t�pj�ة�0D(��JG7�M6K�0HNj�&ҡ�n��l��)�7�#�8�9�Yw��=�@��:�KmI������5F���h7w)���M\��R�֒i) �mbΡ�w��"�s7�}`b�Y�>r�,�2M���fJ�Ja'���e�I�H�9�lz������c{�=���[�p����E�lF�p0J�g�(�����磸v^���\:�ͤ$���x7fI�;�]�	����;&-u��c{]�i�J⫥8q��ܧI27��*�_b��P�>�Ffv2�O���p#�aA4tW^��]�*�GY����]�v�;Q�v�y�7�]���G���X�eHX'�ӯ��VG@Y��#���䘬�"�#�Zjsr�D���������I&�tfv��pfv�f�W9�(Mc)�b,��2wVx*���L=�{|5c�$���cw�vp�ա2�
���5.�WGrL��rWV��똨I���E��q]�U&�2c�.aj��Wh�x<�J����>6,me!�M��ߺ	�E6i���7Ƴ{;�w�N�͟t��CR����[�C��ȕ$�uw=@r�k[a;{��c�.��M���ۅ+����W���.� (��o1��aA��F�y�li�s;
���i?Kw�䕡�j�GC��)�(R/ ���d, �E��7�:v��ʐ�˔�J�L2
Wl�<T.mZ)��*�������m��������d���b�����r�e@�&��cB�iuc�U��1�C���+�I���\�WCӨ<�4J7i�rbV%&no�����Q?c6͍����{�*�Am%� ��)-�G]ܮ�Sk:���+����9�]�['�Q뮣se����V,���2Pnu,��TqN"�nbS�`��a�]w.��_tʹ�[��+�6���1)v�E[v7t�J��b��<�8��&wB�@�عŴ�fƣZ��(�uJ�7I�gi_���E��>؆���������Y]2ow;��Ӕ��Ѯe��k�z����)�y0��	�Y*$�p�D�WWW}���f��p����]�+pV��Z��wӮ��i�}&h�t��2¼�f������{fef��K����Ӌ.%�Ɔ�ۃ�[�u�7�C��x�����*t�\>��b�y��r�6�o��woi�d��������«�A�ܦ���y��6�	��y�M�V���v6�s3l�Rƣ"���eSͼĭ�o5�h�}&-V���[�)�*�S��u��J��Aկ��qk���"�~ʤ�C�۫����>��,Jo"#:/dv�^E��Ôܼ�K�LMwGDK�Z�	֝b
;�o���Fd��N�p��0f\�F��Rf��i��_$3Lh���������;��w��l3h��0�.�̖M_:8�s`N�e�+�	��I�j�s:�dqo9Fg]:����yW|�#M�X�'�ƕa���_�آ,��\����HV��1������9�f�$���	s�	%���Z����4	�*Z ��U�{r�T��O;��o68��o8!׷��w���53��{��"@/)��zv0V/�T6r���Wr�m�Ζ-�ڤ�GhE� �R��V�Ь��q���T�c�ƴ&�9��O)Ӗ��7.=e�u;Y�6�!��U<���vخ��������d�������K#�u�� <�'������ b:(w6�n���oM�:�uu���|�kD����r�u��wk�.�4	�\h�u�5�r7�P^	`�mI��nS��)�ڗ]\��a�b���d�2P���,Yh	@K�wiRa�l�KE�p��J1.�Sڰ\��f�H�O+p٣�]���K��̧����T�@��;#�k���t\�j�uot�|�M�̓AD��������&��k�ic������9�ed{ ˗�{5��J��tT��hwٻM;��$]u�a�>�fFh�e<���5���TJ�q�Z)t�uTe�Q�Bb�.Q�۝X�v�oPH��@l�������.��x�PݙJ�;�4�n�V y��c��tYھO���7�h��xkA����=l�M�p{E�����k�.��Y%O�z��{V멑f���m�6�rAXI�s�Z&��k��_u�tx� ��(#:G���:��s.�LD].`}}�_.� ] �\�M\y�j���k�&I����ᴶ�<��Pa�;4r�)-����H0i}���,����$�O�@�)t 5.�a��a:�+*��8p]����[Ox.��9˥��*$*GE�k)N��&ӽ�N�Yx����7{�T��fd��T1�UD�5)H�i3oYD��d3�[���Ne�8�q
�d��$V�"J�>��7ZN�T�ZT�9�n1q�Ͷv��S)�<�f�݂�d׹���E*�vQ�8��4cH:0o'Q�7-4�]X�6lh V�����ka�=�Nw� �����:esʹ�*u��D�.�l�G]��`rʑ��6R���Վ�9;k���qs�Ҏ�pZ�t7oun,¶��GeWgZ[ab��:��6we�Fn����S�����t�!��d�ܣt6�C��MS��#Si5�3m+LX�7�t�j�K��`���R�nS�aVFNm���⻆E��2�s�v�m����ll�[���ƪ%�ʽĕ.*�,��j�����OڍN�Lhnj�ٮ+��u$�Ʒ,v��XJ�J�N��Ǔ��-٩�eɼz��u`��W#U���L���րR��Ri�O�$�ޥ���Afߚ�����1X�VH,A�\/6��f9w��=+N^�VڠZڀG,\�����7`)69��U���9w�����2oXR�v���-+�g;���W�:L�}>9�mۇ;o]��L�ǯ1c��
S��2���F��g@����3,\u�P[�e4�oܑ�*����hju��7�!S8�x�+��[������۔u[�%�Ǧ�;9�����#<6pԭ��D����l��v|n��.���Nپ��{iА#75���+��T���\�J$i[�,�NuF�V��x+�x����IR�o!��,�������Zg,� �fܱR�V��n�0�Z�̙����|‭7������:v]�,l�37�	n�șU!�m�Yӄ�kn�Nq�y�u�����x�к�6�k�aG�J�W:"L�.��T�Z��@Ef�rð�Z�ݩ.U0.�s��V݈�o`�8X ������k�6�..�����,ucrY���c�\������f�u\�R�s��g�`�ed�2훩��ܭ,�N��kq�Ŝ�7C�#.��%w8 �먚8��֩"}5p��wrS��{�r�*%G����5�5�;#�+&�Ȟ����%:j{�e<q��ѫ��]YzUln�p�|U;R0ɺ��2,�qv��n.��'�r�4dI�$�X��W�9o	%�/�_D���	+����1��D��gj�+1p��5(gH��hx�y#��F�\2_¸�]�����<3K��#`>J�+L��<~/5�7w�E��EK��5�t� �{���6� .�	\��4�j�`޼S�כ��[}���H�qE�����(��{o,bws}'��Q�%�j�#�3�R�2�W;�;���f)�菟JS�a,^���.�养ی5d.�G��'uh�H�@���1�_|WW'g1�S:�u}،��(G�⥞��rޮ���v��,N��3�D����Ӵ6h�G!��w���gr)�I$���u�X��fnjcC��ټ�T=�w�b�P���q�z�	|�$�7yf�_p�ݱ�R�e�I��7^|�&�wi'�vU��b���F-�­C�Yy��k�3q����g&W$�1��Lg,�t�[�&c�Vf/�k�˸�Ѓ]����(�������W�o�F]��At�ϕ�#D��뿗`
5.�����1ʙdNE�n�b�*��:�T�y;K��kI����H�B�&�OCۈ�=�;�����O7}3sN�J��]1�h�l��:��L��=�Ђ�f6kH;uom�]�����J����|byYJ��oe3@�����G�".��n���%�8lZ�ZƮzyl�x�j0��jN�!>�����Y��*���7��`WԜ��ye���+�o	nF�h�i�آa���sy���୏@�Z�rɲ�Vʓ�ìvn*��yp���f�t�kn���L+F�y1�_To���R����j�(�4_u�Ц���91���M>�w���:���w�1k�I�E���>	tɖ���#�^�7�Em�8:���`a+.b��/�Y��xs"u�X�4/s���&�[�kR=S2*Ԝ�i	�hc�h`r�h�ó6�b̊we�r��;6�ݽ����N��z��0gL��b�.}������]ī�Re�3�۹��1E8Ďk���%�k��}�:��4e�t�݌��۴����!j��l4��C[fT(�Mᜡ)�;�B����X������gr͍EV��4^�����`$��݂S��`�A@5�t/9�J�n�V6�s�V�� ܽ�m���G�3���v�+�w��8um6��\��w�H�-��Hnv���2�7�Х%�v���0՚aԷ̗��޵�*�#:�9k(�[��,�j�grY�3(����9��.�����]���m��.�2ٰo��[�o̴�
��&s2>>#�h����T��<�7xq�x]��=��8�5��o0����3�B-	h��,��cp%��y*��H6yf[G��(��X*uL����g):��g{�_�H(�ؚ�0� NYű��j���]�yۏ��aE.��b+:J�z��s�.�v_'�� y�]�bg;��W�V�8媛i"47��goa���MK���	\��y��Di�%5]9J�:���eU�;�MZ�j�V��&��+�S�����^Y��p:�s����X�J�`�yf`n��^ԩٔ�je���oSFvfҳ[%�kȷ��b^�﫳I�^����@��W�3��DJ	}����a��7�����Ǯ�����)�sz�Z�i_ �ɣk�f�W�L���V���+%N]KupNY�ls=��C���NዱL싦�-X��jNVyd�h���u zs�ꛐ����@$$?�B�\�����}�i��E�/p,�8)Ok��H7�S��������
sreA���u=�]O�ƵN<�[;0���d�\��T����P�,+t_�P	f.('�G��%i�/)<���D7MK:��JD8�����K�,��yu۠�dC��WAr�E}��-��Z4m�w0f[� 9�z��]HgE+�d;�ٕ���r8�g��Xw���B��w��\�%W�٫�G/2Ҿ1�5%q	� iW5a4��B���{��c)j'��{�ڽD���N=�wgëU�oN`��ELڲ
n�=���k���)�;�Q��(�18��+U�pQ�;��7^�y��.Z�~�\܈Ѭ���&	J�;�����=9X�/&��J���a�C0[�}J���&����%gcOv�4��Ñ���t��.ʛ}t|�s�~�����I�Cd[����6Zv2^������Sw��7����kŚ�| ������v�p��}-o�ⱡ5�E�Ed��%�J����q�"�وL�7�&U�B�oE����8��,C�7�A*���5 �h˗,@Tܙ�>_ǅ^;G+Iv��F]�u�{���2iRm�N�íŽ�ܔ�\�xj�<Pqr�9�����J�gm���1q&��� �4��<��W��ne��s�Ǳ�J�:�Rv&p_gih���NК]ܛ�(�Yռ�ޮ4	���Uf6�bԀ�lY�:��R*�KJV�{}T�Zն�1eZ������WY
��o��;���ař.�w�	�~̏��Xۭ���Ï�g ��s�<�u���3:D������h�![s�A�ƴ�2<:bQt͘�[����QB��Tg��V\�]���R�ʕ��sN���T���*���gj]X]������؃�'�����k��V��ג����D�{|9M���uݺ�(l��)�x��'�iU���9:6����/���ʾZPb�2."��a�WsQZ���X�([�&Z2A��Qҡ0�kY�,,�áoۯv>��V���!m
z"�V�Y�*�{k��X���5��2&a�w�V*��T����;��]pOz�v&�)7��TŹ�����|��'R̴��g�&+�˚	���|���s6r:L��nWm�ŝ��iO��K���� �R���żG\����-����\7�Q��J˚�Y��W��e�]%�*b w�o>��weګ�5vi*��|X{D�t�϶�N�	�@I�������ܳ�Hڋ��l���ԕ�u:Y&�s�]L#�c0�|]�Q>��`s�8Ff�)�a�/Ji�w{����@@�ݔ.eeiWO� y�8Y����E�{:s�����TX��.�S71L8�Jge\���.:~L�$�j��h���#�C�������
��9$JRnо��V�n���|�b�%YJ����X*��ْ�C��z�,�n�`<�n>uC�%p{�7�fEL-wZ�5��o&���Wc]9^x�-�e������uߖ�P(;���ҽ�B���{�ݕ��jA��s^����X�bXwU`fTX�r.���-�dW	�g��]Q��qgd9*W`]'��;��P����.���j�\�'��-�(�9�	P��𪘦QF��u�Ӎ��a��xh�������9`U��7��yj�L�3(�����G%^�$��J4��P�d��'cK��Y��y.<�7R����LJ�m� aaba)mb��M�V�����<��s��\�� nw5�zM�p��U����ڇ2��9���������Fu<VAX�͟`���y��v`�8v���r�O�ބv�efvP<wW�ғ<E9O�d�����#�e,�N��&m�(_u���bFA�Y��a��7Q�Zi��iQ��rn���Ǿ�z*R
m`;��4.�N�Q�"k�����ѭ�^��S.�t���j-�R���nwU_>��.����K����}v`�%��w]-�kb�,�iy���N��nź�����;����C_ƛ�s᫱�>Pk��1\��qP��<n�j���git�S�����X�S5u�b:��Α�� RY�|!Ϭ	mVa�$��ŷm�h�Zn�w�9�B$�N�Px
��CV=�z���{r���DZ�#Wy��Yym��a�B,�Oo��ESbY�0n"��9�"[(c#�ӱV�k.̑h���)�P6/�<ʭ��m�s�.��ܶ�5m����A�wU���3hwٴ�aH*W*U7����l�d�n\��d�1��\Ѓ�,!��I�Eޗ���-G%w;��6��G`WmE�B�� ��t�|+��e�0~n$)�����ݍ��ٓKma�7��;��9���a�OkcX���_dN�L�g7TTft��W�p2l!<ojL�N��[{]+�V���#ά�x�ve�ƬGF����DZĳ�r#�K妊�B�V��`��2Hp��ŀv �J�-�D�p.j��H��Ҭ��-u�]�若ue��e���0�Oe)Wԍ*y�Yyj��&��u=뤳�y�a���H۩�o�L��A��^U�=��Cm-�r��׬\Q�f2WZ�e,���_e>�:c0�C�<���ε.�f�A_W>4�:�Ѡe�$&�+�})b�6���/�ɻ\q�.�S�L��L�]��3���-�"w,^�5���.�aP�� ��z �pϚ�df)�`+?
��+����a�R���ʎ���2GO�r{g�h;Z�^����>o���j�Q��Ԯ<��	�+:m�>T霡�܎�,j
�Jy2�J�$f6!���_U���P��mJE+�v伅�ڎ�+��J�l_R2�E��rMˈṚO�����r9��63��'}�3�N�l��qy�w�m�1���s�g��j��9��;���0��uݺ�fِ�{K�!P3�b��:�AT�_#�0���Ѧ��G����.�`Y�f��ug4�*�.r:��+�*�2vئ��ĥ�+���eO��ͭސ���At����Ɋd��|�L��u����e�#�s��[�X'|Rυ�u�+�`��Y\/uKu���C���ndK��)�c��k�t
0�k����^WWd8�h�3���y�ǴR�e��'P�2m��f;qЗR�$T�>�b�}��j��ܮa]��ν5���q�E�r�4o:՗f�������N�[�A:q*eYYl��'G5��I@��'m)�x����2��`ૺ˰)ۀp���g��y����j��2�����O�j�ȴ��,\=�.�Ⱥ�k0\�o���մm�%!�:>�o:���=�gMX��ԫ��Ը�9�����u�W��N�s6H�+�cB�<�m�!t���oR��|c�c��c�M!6C��],N�0I��D�xۖu���k��;���+ 3���``P�J�����=Jw|)9�b���O�I�����-��S�y��XS޳N��v���&>�O�A��B�Y���Wg6eJ\j���+H]��L�����R��ͬ�[}�nWXs��`e`92�q��t�V�[W�e�?u*ġo]�Y�sL�]�F��;�ۺJJ�\k�E��Μ�yO4+u��0}X��n�Poh���5D�8\����>G~�y��;�D���T"휏(h���,�� �24S�8��۩�]�C��$�h�U�1��ե�e�ƌ����Y�_|��x�C�R�Eul#ق�&"�k����w�;��FQ��8�t���n��7���x���>�Y3�n�u]�4�d�K��uM�EQ[���d����v�o)���
<d.�fఓ�X��e�j�D��@[�+U�y.�e҅^.�Z\��R�Lj�Ձ)�)�MV��Tʻ�N��s�3HL���-]�ѥb��F�5va�L,�܆6�g��^N"�*�h愘r���L��9tM�Y|7�k$�h-)�el�,�>�7�-u���;j]Sl��̂�ژ�q�K�/u�:�'�*���n�sٹY��j��z�%Y��|A�(��a}Z�Z�.��Dr�r�'�����o�������uԥ%o�e<��Q9v��+ef�wX����b�kz`"��T{6|�ݖSխ�|�F*7ʝ6e����2\	Pb��Z���&JջZ�0�L���qhN}f��2Su�ΩN�"��W�E=�^%�m�Z�k�a����� =*�F�㹚wWԩ��R1�ڐa� b�M�Z9
��+^��Tel��nce�]�${JA\d7��ڦ��� ���%<�DkIl��0w����œ�N������2�z'��;��g,L��;Ro�Kc�+Yt�zk/���|c���x��Ęhq!w`��G�tn���v�ڀ���6.��1]�,V��.��X����d�X�3/[�����_7�>�𮤳/V'4���ۘ��6'��p$M�JP&��gbW�b*�ޑ�'���vV9��Z5s�+K����3d���w��y[��2�q]������.�ੱxwz���k�g:��%��#�sW]Dl��r�gdEWZ�x�V%���6^�ts0�?�w,�(M��bϳ�&p�l���̄y��ZSg0�{�]�n`â��3/��1:� �Ux�v)ϖ��p�t��A��aӶ�J�E]KU� Pе�!��z��	YS�K�I<�w>��� R��@.͋Z=\a�͓}�դ�i�YN(�r�!F[�k���u	�}"�.xκ�}��ۼ�MڬK�C'��//��w�6�6Y�3l�C3��zLU���&�CuӨ���ᶪ����*x�u�ENtM��S�\a�j�폯!��Z��kC��S�[���)�g8u�x]�;;�0��
U�y#��%&�Z�(������u�0��'&�뭬�8EuIǜ��r�T�﹧��D����Q��d��C"!j,���K%��������̛l1�j
��\&Lk0nU�i��VR��b����i��:����I\�n�r+-���h�'q��G:��P��'ag̊�5yҶ��~�өt؆?��]wLF���H[��_%�oC.���`�v��^R��d֬�m�g7��9�o^����P{�]a�U��mەnrA�kU�]�=�����=K�Z�Se�Z�ux��R���;��9!����5f�rN�ċ�8���VP኶����]���M�PM�V��d�	�"Δ�(E��8���|�u�s}�q'-��W+dIXo��b��$]eB]����ĳy���Y�S�֩+q�����-`T>�e�jDBۣ�E:R��*2&�r�yس�*eYY�~�YNVQK9���d���}Vtw�y�k��λ�]�Z_n���e�dE<�{Yz���Xʺ����\�Cb�ݔ0᫨��:�ж�f�C4��mR�w��u�����)�$��SB����wˑ�jwt=�5d���!"կx�ff�-X��7�mڝ�F�W)k���U��ev-o���2�ѶHv�e�c8!�]*{J���I9�d��VS���m�E���˲�Zv�.��l�](�噎�@�*b��X�w,���e�G֯�0)���ܯ
lP��V{����B�����2��0�&��
̾�#����C�SY�f��Ҩ��QۚpsSp����*r��8�&`N��e'6X����4$a�@�\sL0p�R�Ӻ� 0�4f��
�"r�l�.� �/8F��J�|,�v��Uk@��6&'�r.T�L#n� ������}+s��w����w�[,[�5-�Fv���YfesWS�t��ptλ8q��#M���.�خ���X2�}:񞬴���i�nC]�j���i��N�P)�b�����d�B@��N����x�7t�y�����e�����ڮv���>;��֩H&�s�)�i`�r�f��=WQ��nl3�uj���"�qݤA"]��[8%
�/9V}����R�}>6��xW 1 �n���(wgZ:sla��"xԗE֚6B;AtT�-�'�W@gw΁3L۬3UN#��Ab�L���%e�Ts���Ybw@�F��SJ
���wg�,��R��e!a�
N,[Ռu��ܖ���JR2qẜ��8�DY��T$��=�
f1�z��|z�Nb�U9��Y� ����:fQr��	���e<|��ȕ���;Z�`$,�u��L��N��k������Զ���u�ق����"�4��v@�$ v�%��|��{���wz��J�4:����Բ�fn�>!�!Sv�d੝�8�Lqm���IfC;�5�������di�W���Z��W�o�/V�� b��3�����M���?Y�����:�R�D>m��n�`��N������#�t_,�b�.�!��/�����<�� N�m"4P��X9�IW�ۺ,��͸A�gN�"�=��໖z+Y�����[[t�aÉӫR�#��M䷰�%m>9cnӜ��>�6�͆h��`���a����_<�Z�1R�:k!���wjP=%:׽��5v�5B����Il'���F�����]8���@�����!��%M%�9��˺�<;�CW�GsV���,6!��e[]��T(LÉ|��\%J�Q��o��tP�hs��C!߲�v�v�#��r�\=Q�U����������sl���z�c����>�Y}��n��HF'%V�N��'X# k��%I0C|*�gM��"5ok�<A�gS��(�L��Ֆq��
VT�B�1�g�Q��ݝ��!�Ȱ�Y3J42}��Rޭ�ݴ�=�j�өاeh�U�J���uԠ��>���꯾�~�oe�b�Q}^e<�"3�7�늕����tmY[����"��7��xV���e]���;{��ju�;!�ٖ�E�J|�P��EJǴ�K=RoPX9s�6�s��Y��R���&^$��j󲶫0�vHJh��1����Ն���BZ��cU2L�;��D�;�K�{J�
��Z+�����ϏnV��]<��mu��T��V�[{ze�˝Mu]8
�x,�g*4�Q�<�
t{�w|%LS�C��P����M)�Q	��&�<�kzhbB�aƫEl�*���:��TJknY��f�ԍ�c[\��`�?��ƒ��)��'9�r�1[�Ш���C{@Yy��r�k��x�dh�+�>����y,]r9�b��p\�|.�V�j�W��0��g@��tX�׎����x�Ҳ���,�k�8VYG�V���5<�+T��"^�6ãV��Vv�׊m�B��
����Q�mN�Z8tW��5Эw����v�w�j��j��j�bI%	��f�y��2�rf�#��t��i�O�Y޾ˬ�P�e�$�o�Z�[��ɠ�v<�ke�ź��&�@\ٝ��/X�{�$t(R9�gt3�B���P�oDAt2��O-ܝ�q%ٚ��g_u�pO��]��we�̈�Ħ�O�l t �w�a}Vk�
�]q�	0��pJ��o@�q�o=ߛ�z�����FA`�i�+�Y�FE�T��%,*e�F)�A�ԥ��&5*ډXb
c�s(����"��Ƣ����\`X��3EE"�[i*�,Ds!��L@QTXV����5��j2(cX�Ԫ �����ĕ"�2�Z.5�(8Yq(�`�D�
`��H�b��U�ִf2�X��$��-3*����)�b�,��Qq��bV
fR+&[""���+�\B���(�lČE��ԬUV�aU�h�F�9Z1-�-��Gc*�ы�R��ZR�(����Z��U�#-%`�ԱIQb��4�X����-�h��E��j��ڢ��m��c-b
[UE�*ʕ"�JV�,1�,PƊiR����UJ�TTV$PX�ȿ���.���������߼R���-������+^wv�ܧ�N�^���G�.�{�*�[F���l�ifwr�ϔ̴TC���曀�t�NY�����f�o�ˡ�'ϓ�ҭ{��Q -<4�/���5���5gz�<��8���I�B�+�w>
g�J�<&�Ctx��s�Io�8���yَ�&gC�e��~�e�[�˨��P�EV�>pS�|�9@:�3c�4	T2��mre5����uZ#�[x&8F}�yl>�n�^腜�3��b`�pSԯM�EW?e�w}wJ��(�wüXB��Ȇ��Z��\/��ҋa��m�<O80�����vNP��Aߠ��]�u�k:�3�/*�3K')J.��>ҩ��fJ�v�#�iխʠ��Ļ������@����V5�O,9yU}�R��U��a�~�;��.��2\lﳲ�b0?^���Y�]���u�8��껅�,��R:)�흛�)o4	v�_W�L�O��<2%�\d�w:Xz��;��&.u�X9u/7��|���{�AKm�u�V���.禡��a��NP����9��h�'����x��tu�.s�dϑ%�\:�#�Y�x�<�볌XEgx-[(�[�\�q���������2��X���G���x�g`�z+S;�=�XŃ�uB1e1�����y�	�-�N)
��Z������/�,�W�v�ʊ�n�������8`ʋ���D�}�E����E�߰�f�P>b����s]�0���V|�����*�����w�3V�DI૳�ᠰpmG�`������M��W]m��Ϣ��rK��~\Ϥ]2�tO?m�P����a�r��v�Z�E�z�(X.�}�Ҭ~9:{N-�c��P�٥���_!z�����cӟ��L�k<��	"J�J�]L���Yx��O7|)6�WW��q<�ْ���ssk��^�Q����g�I��B���;��NU��w)��P{Zq���jJ��X�\�ݞ��Yd`�07�%�Όõ�Yơ��|����-o�u�ؼ7[�[�M��G�P�Rqu��ϷUH{�,��L\�C�!�~2J�=���]���bxy��bJ�uF#@p���<3�O�.��^k>2Vo�"YX�F�H�[k����:!K9���tZ��8t	�|�)ȑz���=.V�����oĤ���->O��,����S�q�X�8�d��Gރ)1Z;(��C�|q}�ۡG�wg��vmeP�	�0XW���tU���9�#�Ez���ۻ�<m@�W2*6�_�l�7���<w.t�)
�z%��8S�S���b=�s{.����U������=Chk\rI5Q�(ثH�̼_-���'z���בc�$�a��z�y�N�&;�\w����i���kBHߜ��+9f���R%g+yF�(+�%�����+�puz`ь�����꽏������_�2��Ȱ���{G��=��%���ʏ���aFX����:��A��A�L��Z�q=_;�}���=9.*��^s�6��|w�3 �5e��3�r�N,�����L�(8R7��qY�R���ꅼ�=���T�p�&��E�'�$�yo���y������s�]�nT�r��˗��}�w�F����'�uص�93m�:�Ĥ^�e��qg����C7�뻞��z�<�Y/�̚^b�҆˪���h�9�Ju_qB*������%�Ӹ�\<��{�S�<�Af��}Dr����A������ ���ʉ�T���0��4��<���.���|���=@�dxdS
�z�>�����.y=3��#���6cҲ.2L�N��sxs�h��%��x�5�JD�#��
+�s���7M؍���!]���
oϪ���'G�B���f!0&05C ��XǊtG5<�ac�!V�7�v�n+��W�V�����x
pc"�{�{�74w���Ԝ*�"U�H	|E���vj�:�QJ�7ʴAq4�k�4ZE����g68���JS/vnZ��]3���s�kn �2YH蒓I&GR����]O��8\�q��/:=E�k��qD��`�p՝��ƅ��Ք�H�,��q��0v\ñ;�=��n��h��gvU{��.�:�S1�A�$`7�S�]���i&lpS�B���e��r��=��|޽�~�
�R�h�ܧ���+���j�1�d)�w�P���/B������5^��6��;M����i�,/{qB0-�Ώ+�3K���삨���>3��Fe�#MJ�V�]��*��}�6��V��U�� u���\�$C����t=�:x���{Z\]��|`^n��v��ݔ0�X�7�J)�Y�D�a1yxu�~�Ցp�W�΁/���.���K��d=2�޷L�Q����^U+����])+���r>�1���<1r�m��ڐ�gh��1��f��]B��p31��!״��v��0����m� ������VĹ�s�9u^�%��)��0�I����w���=�1����v
��_yіZ~W^$��M�<:!Ѿ�ܩ�%���a�U�[N�T������j��ban����*ؼ�0�իU �����^Ú����-�i�ZW̛��)dQ)uD���X;�{7�*q.O��5C)�<~�w�XV`�9��V�-ǜ�
<�
j����m�zX����J�{v���L��c�g���cZ��o��6����ֈa����6v�Gc�5�^�h'�:�Ώ(���L�⩙���!zs�0�E��YXb�ҹ����R�������}���`��C��ԃߩ�MY򕇱M��L���I6��x�#��w(+Y�SUL�wH��(�LƴPL��q��9�<}B��Iw�eouZ��-�BfZ�ܼ� R�"�}��(����"���d�r���3�<�}պ{9�#����yar�e�X-���~�^}�:a��+�2��0X��H��o|���\�Or��b�ssLPWZ���'3.0b2����Ɨ�:�=բ�/>��x\mhx�.���46��*b�I����׼�s�A!�Y���U0�U�`�����)�礦-2c�^�r��u�C\����Mp�2���ߥ��o."�9��]������{y�r4h��잡+��ek����*a�IA�����4�u�|��z.�����a�e%c��&�(�E�C]����E[��S�18~�a@���3�0�!|f�-Ӆ�΂���Yݖ�6�6Q��5;�KV7��KerX�
J��핚�3y8a�(Y`����w]՝b�j���m�R	S\����O�c�z|*7}C>}-q2P�z�%�L�;{U��R��U���*3�Q�k�g�����-��P]c4����o,�E&e-y�8�#�o7.�NB����;�\37\O��z��}A��/��)i�p�e�����{z`~ ���Leg[�U��;3��	:�F//��kԶаP�V���.��b~��s��e�㜭)&�rM�w�qй�0w����FF���Ғ�}U�-b��5��:1E��ÿIY�L���g�[o�{�+�uۄ!:�w��:�X:,�<CG�eRKG�V��&���|�a�x��ʣޗwM��u@�W;|�`�׽��a�bY���Z�.�X�G���f[}V��{u�4�l�[Y�z�_�=!����=X�5������B�tD�_K�\����M�(g���{7�V�h/�.%=��֋��]��^�eW�DؗR�����̶sl�5���Vsȣ��(F��8,�Z-�g˲Y�w��#���L�^�.�"��4r��B%wۤz��y���V5�%���R�/,�N�71�[�<;��g&��d��ս��a#�81�9K �|���2��xpW�)Ӫ'^P�U�NY�Su�f {��5|�ыN� h�/Ze(���fnI�Za]��c����}O��^v���_S&�z|��EE��qV)H��8=��C�Ie��D.�9j���z0��N�X����1�j�1�y\���,ʔ�ZY�b�;.�S;�/j�{Ԣ�B��S�wz�buH�5�!d�.��i1I˦|��{>���L9{���+�-�����N�$_)����s��?P�1��R=cr�T����7j�ނ�v83[{�ռ�z��4�|�e�Q���] )ί8��[nka�k�勤9�vIGB��f��4nj�d���y�O�����>�J{ ��ŋi�C=�q_��37j��<�6�.<\-��wH�9���/�x�q������ž�}�[��U-m[÷0���-���g+{
�'ɸqV]vN��m��_���ϷrI��U�����SϖS'fV�wlv�W��f�}�k����t��ΈS���n۰��2X��{Ï8kH�^�'�l%���%X���U�6N9�]b���&̣��N�Gؘ��l���
�Ë�ёҗ�3�-��ʲ�
��i��w�L6�1��7��(��
��V��[�Az.���we��b ���4^*9o0�e�{�7=����5�5l�O;RsJuw`+��-��X}�=�	�6]�< >��]�������ޒ�{��]�<�[�Bﶵd�Ӟ=�����,�ǗcE��A���.k�����^��ȟ���7���"���/��g�ayu?���w׸�eh3�:u���nm{�!�j���k�.Xi�Qn���Y{�q)�!b��E�N_2�f�k�x�g_W�>nH�3#P�jp_�UwZ�\�X��+CWy3�#��N7�U�~�|˻�6#_t��L[��Xs+�t�w�gՕ��S�W!�nR��g3�9c�7�wD��CO�����Y�ug{�#~�>ٓ���%�R�y8T��ڙ��o����s��V��9��Ob�+u'D���g���k�9��s_eg��[��j`\�-�I��/��zs/���
�N�l�R?���ńm��"�{��r
�hp��`� >"����neu��z�A[J7mP{L���K6����.+-�c]��u:H��]�
oP��V�1�'J͒_,n���ѼiR���9�JTѡ3�6���A�Yaj��Е��"��i{�m;�P>�|��k����0�s+>O��vm�o�����to�T����z'�1���㦣��7w>�Mm����'��f�=�dׯcs�w-�q�+ON�����d\gj?j�aʗ�V��=�tUh���߶�@�lP��Ho�G-����͜}��*�8T���6���a�g���S����
�͛�$��W�&��s������Tv�j����gQ��v�8`����jUp�6�T����^P���5��;��A�sސ>�gZ"��,P:倇:�u���{a���g����%�m�O�{o#�Ԏ�ηE��0�\��)+��x.��SW�k�q��N	�=*D�bϣqz�_d�����uO��jB��O?i��ݗ�)E��Ǜ�@��C}�93���&*�un9Wu��v�Y�r
�f��;l�6_D-���|�Ή� �4�fU�f�-l�/j�;hM�z��Omp�V�xX��&'i=����WƏ���"k�-�kE^��i��B�[�fZ�pZ[/j7���Ps�:+�Y��ƥ���T��N��ח��Ξ`�q��5��umw�:+o�dp6�4����&y�UN��MG˗��zf���;�u��{r=���fW:,c����0�o.0��^/s�ߎ�����ɾ���8�$]fEd�����ޕyJ߻˝���-^�l� �_�/�<Z��^�T�>\uf�su�Vl~�c��X}����i�+)j����%��橺������+��GK�\�������H6ԑ��\u�N�j���GW�z�)��F�7� �@�.�]���{�b�\3�,'/6G�}5��3��YJ�Oyv�m�S���Y�����8нb�H7�C}��Nt#�n�U�|�C���'�ik�Or�������YN��V�h}|�1���������vn���v�ࣛ$�>�]�-��;G�cϒ׵*��nݚŗ[��K��Ie����CM�5�K2�Ha5����)����꘲�&��`rE.d���
<a���ĕb�����G�V���:ﻩԶx�;���F��t]̽��h=��:�g�5�S�J���Pͱ-�O�#Q�q:�^�A��7R��R���w~�'a�f��Q}%��j)"׺Qx]*�1�X��X��[=V�`cQ��Y:�8@�v���Ɠ���uP���u���7�:�mJ�ux���Ϟ;��NfT��7f*�E���2��G���z��]�R��:2�t՛���寋�ݭ��з�X�Q��詤ǜ#�E1�=^D-oqڬAxú���<��>-B�j*{�]WX4�5r/z�e@U你�n�^y4>�E��������-� B�ޡepj`z�u	������Dm����̍U��b��&�},�J�a}�>���z^j��_4�W ��C��DV2!�&գ4%O�+��y:�ny�ԏ�-�.�~'�h���J������7uy�VP��@+r��ri�ղj���]�^����͂I��6�q'iX%�Y���%������� `���LA��^�{NF��:�v%�#M�V���#�Zigq�WL�`]C�����g�s�G�3@��/qF��zќ�Js�݅��}6���m]�_u��ٮ5�<v���Y�%r�v��xJ@V�z����:�T��ȴLۊ���Ƚ�
�M���)�l��1R����0fY�e���&�J�''T���ɢ%l=��f�ol��N6M7�m�e�H[+6��y�i����Zm_[����I8��W|�K��t�|3���/�V���n�Ã)2���\����4�Lu���t�p�7���f�򏤓p�D'������N'[�@v��}��:�뭷���W�r�a�h�)uul�����⢺�ԉʮv~�dO!��B�0f,� ��X90~IX�hK]A���n�˹k��8�;��#k��5��
��(Yo��z�����t��veEy!�"�^��������Rҩ���9N����̺����:�Y��W8���dճH��Nr΍|�|���h=��X�N���Ǝ9e8�嗋��źxy�*�r���x�qͫ�_r��3t.|8���T��=tAqxS��r�ƸU�q}�N�eK��?_TAG�d��5;*
U���Ƶ+�f��S�^�.�Y"ހ�
�38^>y�^֢k-��i��:*�]{kp����������2j���|i��1׺�\���&7P��h�=uZ�ئ�mX|9l��2����{�s�^)�9����Kč�V)��.���];��Q�c�[W��v�Gh���x��O��uI�֨/0�!�3ka/���{�̩;���Ӥ�&Kmи�i�L�Z�r�#��9!�¹nvr�ٴ���wÃ�"�L�{������X*"��,t�)r�ȌE���m�ATX�0�X��9k��%q*�̵PDS-�0iX�P+*���DZ�UX�������TFҪ�J[c�r�m�̥2�TKh,����QITr�X�\�EA6�c*T1��VF)�b�DA*�F�q.R���
YF
���֕VJ��m.d2D+(�iV������P�+2��R�3Je0�k*�fa[,DUF
"�X�[���1+�f6�Tm�"��L�J�9J��YRَe�2���QbU�l�R4�k ���Y.eq"�UR��(�e0PQ�U��b6VَV�cXe�e�Y���˘��kX*(�,̪)W�30�E��c�[q�Hګ��m�kP���ʸ����˅b��71�*8։e����30�LZc0�2��-�3.e�Jc����)h�Q�Kp��%-�V�F-b*[X�)s�k�<�����.n�W/���aSy�
�����/B6wC��Ì;\E����.�9�q��u��"�y��ǁDd�ň-i�4�ו&�X�{�^����6Ҏ�pqa����)伷�~�1/?mkGo���|������v|�5hE�X�y2�ˡs�|�x�Q�Yը?\�.�{��@Cv<��&瞃7y7>�5��)��.��/s6�{cF�UOf�&������y�|��ص�:��7R�љ�oAaz[XY{�zu<-���N�aӲPl��M�Q��͘=�0uZ��U����L�M_A�C��om�����*~���,��؂�v7��ߚ�j�m���/>���1�p=�]���I�L����{ONF���J8q�^�����?9�y��P#�����]N�x�>����r�uc���#L�f��eiP�e�Q|��/9���/����n]�ܷw����~O���ۘg�|��\�'�z��I��p��{��E��z�>G�;�y֙�=泸��W�e�p��\r_���I������2��w6���K	�N�]l"�Ό�.�j�m���Q5�[T�,v���y�r�����]��y����E�Vfh'�!gG��e`�[�����s>l����e��^�{'���ǳKݣ<
�OkF\x�[�ޢ����]�H�O_�F+����J}[�_^�����|�<�;a|�ҧ������gl�c��:Kφэ�5*i�ٸ$���[�Vev�v�d����|f�]]����{B	���A7��@��C�:ö�YцIǻ�#>a{�kى���d����p�W�Xw�y�~�Oޗ�m��ՍU�Lo�o+����is���ty�_�͐�.o:��v���n�[t������D����0�v�c@�5��n�.mמ��UAvD}r�&�9�0o=ݸ9y�A���x�7�4��m�w�隆(�*w6+{T��y8�7}��q��I�k�.���=:��*:�]{�W5�5��u<�7ҥ��C}���>�_s���k�:z={ot:_Z�3#��L��coŴ~�&�!�95�NL��e��+���P�jj]�񕽊����v��R�~�� ���N'j�d���fu+�WWF�	P.�J��p4�C3kaUy.u΃k�cy�¾�xB�;Ң�+I'q3'b+�+��y��k�����j/7���o��$b&5��,9��X���N�߄E��^�Ci�( I�ū��ĵ?w�1��!zM�ۥK�msȪV7�y��M���g�W�/�{��w:z��{����dazx��ک��=H7�ʗ�+sj`\�-�I��!\���G[+�9^��}�%��iA'f�u�D��@���f,,˰�WQ����)��NS�����ٚ'�<�����j�:ϔs��f���N�պ�yv�Џ��B�E1��*	h_�໤�=�`.dC��q纽�³��nw
�Nf���{OT[\\9��/��ǘ�ߣ�N�Ǜ��u{t��+�S��֞�Ȭ�����il��_6o�bL�A(\���&�T�q�t`z�4���B����������is�6���6lc�]0�}�<�	���(;s��ɪ��̡���ݝ�	X3p�b�Z=���un��N��lm�����.�G&/�Le+��0�ۛ����&��՚�Νʢ=I'i}:���M�,�����}Vxu�U
Րk ��z���w��>Q�"�����8t�r��vG��H�v��_����u�l�6�ُ{1�_�����\�oM��5�#ki�_!��r~�{R�{���X��nU'������I<�D��bϣq{~�3��0L�yB�Z��P�G�x;����?uX������`t��Q���=��I��b��fR�u}��>��2�W�f5�V:��c�]1��XqF����*ǋ�{���K��{^c�P{-�U=r�ѿ��^O~�tH{��Ցtb���.�Y���Zj�s�3�z���{X}�ezc�����Ͼ�G���O;ہ�L����{�L�/'c�_s�������%t��-���'Ss,:��+w�<٣໿;Y�D�v���R�������N0�OO��&�:���p��:���è,'�{�u��P��<I��2����OY?Ou��� h0�X����+����<�>j�{:~�3�'�l������|Ξ~��M�5<�3L�b���M��N��}�$���Y���=gǼì�J���s�d��}�~h}���]8��ٟ�2O��s�������b���T�����5Kw�]i�z�n9W�ܴ��gJ�*5�bv��@յ�RTɃ6��=W�[�-�Zvb`���5VR�Bo;e^ʇ"(�s��S��;+���9�`ڬxfio�.�+�r��[����b�L��9I�R~d�je���d�k,�$�+?k�Ru	��2q�[�|�:��>��N���N��'�����N?0��^�cO{��u�Ͼ�����̞�s�N�̓l��A��+'X�I�R~I�je	�~d�Vq��
��� �Oƶ`u��,�9���N�����>�_\pC����sw��{S|^�FI���6��ԛd��a��l�~�Iē�Fk$�>d?����a�4d=O̜J��|�S���Aa*~n���ߨ��})��t���u����'�4ʝ9̐Y>a�S��q�9;��2m����&ߙ5�d�a6��d�'�š�+'�X!�N'�Qu��u(~H�ޛ�g�~:�E��]���������N%`h=��d��=�� �?r�>��'���i4���L��6ɨwY
�>O���T�$?[6����W�C��繚xP0fg{������8��;0�Oq?ẇSL����'Y/0<d�'}���ì�I4y���O?2y�0���&�';��M2k�_��������\���2���R��p|h'M��+'�,��N��&�q=Շ��8�s��~I���XO]��s'Y=a5��^2x����a?���T���_��m������#��&':w��q�k	PP�>�IY:�����M��'>Of��uğ q���:Æ��Y'!�ȫﶾ?هg�ݿ�VϿl�����m}<I���a6�2m�<9Bu�?N�d�C�5�T�'�+&Ҳy2��d��j~��`k�\I�N!��d�t>U����?%u���ixq���E��Lg�;9�<a�I�9p��Ğ�xs�̟ �P���~9�?2N$���*T��0��|@��'>d��Fj�}��W�k5vunAK�-��.ȴ)��������6l������Ǩ�KV���QQ�q����whRˁ�x}(��+p1ޢ^�	���ty���*��
�=��D�X�2�D��k��C���wx̱Wf:��,xk�������h��5B��_�=����w����OY=C�7���i��~βLJ����Xu���9ܚI���w ��OPY�n��ORs���q'���/�I�_R,�|I�'����W�}��}���������vM0������'̇�^d����I������r}��$Ĭ?N}�PY&?�ܝI���w'�8��V�:�䟧�����'��E������|�3�7u��_Rm�Bx���іd�>��?2q���x�d�N0��d��N1|��I�a�o��LO�s�m+!�w�d�+{�ٚ����{�s���y�=�l���$�&��.�u�i�,'ϩ4ʇO���X~a�g����'Ru'�y�q2u���z�_�}ߕ~�}��c�j��Ik�+-���3{���Ĭ�No�d��'��=d�����1��Oi=k'�N&��x�&��,�$�*~5�!�a5�̇�A@���M��N���=s2�_o�����y�y�����	Ğ���3I'�xoxq��XO��:����́�	��2J��z�La�=�!�?2u52�2Oh_�PC�g?	����.w��+?�>����>���z���l�d�Vt���:�2�g��>�ì�}I�'{z�z퓟��q�|�3Y%d���|���N3Yd=g�N'�}����Ӟ=�<ߚ��w��m���$��qC��J�ל�,:�Ԭ��A@���d�쓬<��@��O�<��I:�&����'���+�w뻇_�?k���{�����VN$�*C�1���SN��k�`q4�?:��8�ĬyH��'_߽���k�w�N2~d�h;d�'{�$�~I���`)���y�����]����+$�:s�IXx�)�'PX)��'R�a>I�����$����:��l����N2u�~�`T'�]Ϟ������}|�N~�s�ӹO�tۈع�m���#� sZ��\��o���m�O|G��}A���-����c9f�b�wHJܠ���\#��#�Xw���o9:��	�A`�t��.�'�t���]l'6;�:�Û��CV
�S�$�g���,�3g�W��,s����?�Uc�N0�\�Bu�d�s̅d�'�~�*
>�hT�AI��6���Mad�I��}�٦���`q���8��;�N�����K',��^�ێcȿ%���}��&�N��l�2~I��2N�<I���	�i�S�dY'��d�	��m
�Ԭ��(a�M�N u=>�>�����O�4Vy��5n��̟�*O��I�;���IǨx�4��	�ù�Y4��;ܓ��M���v���?u���C��d�*I���+&ҳ�Up���������]���0e~�^���x�9�Cܤ�'Xx{�!]�is'&ޡ�w$�$�Zc&�x����X~I�4r���~���q#�>5������e�Z�u�m_H�~_��%d���'���m��?P�������N�u�B�d�~�I1���'Xu�p�1��)�܂��z��r��OYa�����g�����ﯝ����<d���T�����d�'_z��I���k�d�!�^`x���'�v��M0��Τ�ʇ�ϲu�$���a���PC�����7�7�݌�{����?~vo�¡�'�ӖC�=d�oX~a8����_,��>�O_u5�Ì���ה4��C�טzβxÉ=>� |�g߫�/�|>t�7�+���;T��ߟ����
I�ӛ��N�Bo�i'=J���a�'��������$�R|��T&�Y?'�a�I���<��8�y�>O̝aԏ�y����Û�^�9�oo���'�=I�Ӛ�O�������3^�'Rq��ם��N2}��ӔY>d�}��&08ɣ�OZ��N���=}d�h0}����.�_]Z-�ԫ=�߼Gq��i��'g�É�N �yu�m$�����I��a��$���N��+!�i�N�|��z� ���ѿ2J����}���c�*��O��y��X�^��PR�v�.�,�z���³���w����7���ݬ�m�/Qok�bW�Z�l��Y��EE�'L@$�/�����e+�Y�%"��O�AU����\2��9�2�=�,�Ш�՚��@�?�Y:^���N�3��<�t���������7�}�{���6��?���I�T���1d��_d�&���6�:�<�Y	�ayN���>7�:ɿl'�;�O�Ry�̓l��5�����Z�[��r���x�}�VL`t9C�VO�6�d=Ld�=�l&Щ�k�PRO�ف�N�Hk�d�d�Tם�N0�N~î�'Xyy�Y9�'̙�=��9��Ͽ~�>�����6���׬�Ú�>d�o�J�䇖�Ԭ��B�6�q�̸�>C�����	��o!Ĝe`h��'Y;�=�H,�a�5��w���~����߾�>��f������O0�w�q�&�x�T�n�5;��d�3�?d�����Ԭ�Aa����u'���m'S�d:�d��f�I�V����}�wW��k�o7����d����t�rq�5��N2~d�?2i''{�	��&��	RO��s�IX����+'X)��'S�$�3��9�g{�ļ����������[���p�������xI�l����'ψx{�8��	�i׉4ɦM����'�?'��M��O�k	XN!�9�$�(L��B�u+&�3��~_Ǿo^�߽��_p�8��:Y'�6�Ӿ`q�����2w�N0����I��gp�'�&��ÏRx��uܓ��M���k�!�I���Y'w�t��{t�{���?}��s��PP�9|IRxʒ�u'Y9�����d��}C�$����d�v��4o�:�q�&w0�$�[1�l<@�s�'SL�Ag����������y���ק��Bx��w��XO~�Y%J�d��J�l������2u���a��>���'Y8��|��&�׿d�	���4��'s6S�{���3������g��y��x���C��(u��jr���~9�?2N0���*V��E�~X���'�?0�'a��<~I�'{>��u��;��]~��~�D�m�败D��wˁ�	�G�D�s�f��L�dU��`Y�����ʿOuĩ�Ӣo�s�Tv$I��ӷ�hQG���\�,�|�\V:��X+b���zH�gM�����>�y��kr�P¦�\6��|;�g-�צ�c:����ŉ8܆�������I��o����;`��O��7Hu'���5��I�ߙ%|d���H�w�O���8�<}MXi���y��!��_�w��g��^{�[C�P��}�o m4��<�y�l*>�Ad�?��m��wԜI�*n��O�=��I:����+�O��̄������F
������'��>��+�ߝ������>f�6é=�́�i��/��p��:�7N������ì�J��i&�zʇd�~�=I�@���_x���3|�ӻ���u�~k'̞%a6���+XOl����u	�<�3L�b���Y&��'P_>�z�P�y���I�<=�d�T&���:ɿ���v�u��L�g~�Sc����� h}��~�c'X�I����Y��M&�Y�I�V~����G��̜Ad�vM��N�g'���I�4g2u4�=g���:�]��}��ts�nۯw�L�>��n�d�'��t5�I�I��IY:�����?$�5�'������q��
���Y'�[0:��MN{��:����z�����o�9�}��sY��'zæw{d�a�N�q�'̞��a=~d��M���3Y%a�!��=ed�!�,�������2O��k��Aa*{���Y��Ipݘ�����W�*��Ӭ}I8����9�'X~��v��a�s ��M�wm�m��}�I�i���*O��YY8�'�l��'_�y��|s�:��y���zq�z����Y�L���8����`x��N�C߻�
?s�Rm��Nr��Ěd��2��&���d�'㟲J�����~ǔ��?����{���y�;*�h,;l�����6�i��̆�L��wC��|d>/0<d�'}���p�&�My���O?2wT���M;9�$�i�y��� ~���4Z����}�AC{��U�f8v�t��opȨ�6�����K��62_'7�����ڿk�B�B�9�4Wh/#�)��d��gT��u�˦�E:��VKF���M����K���N|C��0��<��:�7�,��>��1��X�I||>U����AB,���,��M��m'S��d7l���y�2u�'^����3�:��	��:��07��õR����vU��X��>g�?}��5I8��;�0I�?5��(O�$��J��P6��6�aa8��~5�C�$���{�!]�u����N<C9�]����:��*�ߊ���߾w��W���>d�OP<7�'Y�M�g��'P���u��N!�sY%J�g)��iY?I��o�5?XN03^�=q'Y8@3�8�KU,r�8����}��<G�~9�:�c8�]�0�$睸~d�OP<9܂��O�Y�Y!�'?S'y�2J�$÷�+&�+'>d��~/��wu�b`��vwg���+�@}�O2x���'P���x�L=���bVo�u�XOɮw&�q!���(q��kt�Rz��5��IĚ7�I|�N>uB�X�_���=�y�w�}U�Ν������	����:�~��'���0�Oa��٦N������ϰ�$����N �4s�=I�O����!�>�>2�����ȷ����k9o��>��9�I_z���e	��'FXu�x��<��'Ƽ���'�8���2��'�O���!����$��<���΁���£>�7�	�������f�a�&Ұ����~u��&�=d_�:����	��M3FP�	�:�e��a5�z��:��8}�I�4�ԡu���`��>���V6��U����]��>d�C�9��:����p<a�O��{;`z��'߽�c'�I�Y?2q5�ǩ4�e�d��O����0�l��>�@��.oL'D��~�R����2i�5�i6���u�I=C��a�N}a<;�d�'�{�2�'���d���������q
�z�d�e#���}�����9G�c��V�J#�2z�慫w�n���gUJ5|̰F���F��]9�u��TGsS/��t�YͷYSz��of@�Ӌk�%/���[
��6�PW����NV1�ʋ@��h�j���6�}�j_hXmfi+w�]�򈍙��ZJ,��n��v�8�H$�>f:�)<�|�P������E�S�ef�r�%� �w�qΓ��r�EJ��T�6r^"jM#6�U�XV�[g
��qQ��L�CH�~i�n���k��}���~��ܲ}�{F	�Yf`��{1l)'��Iа���)�w��Z\�*U�e�J;�oe[M��e[傡�R�GiR)��X�]]����\��I�x5>XK��bwa�$]����.��EW������b�\���9*i��\Аu���fӒ�%F�[����(JǮy�t�%t �������d�cΗ\����71��қ3�^�}���uv��*����@e��W�Be����}�}R��X]P�D�ٿ��E�!qR-�u��
�|Wr�_������nKT��V��4�ׯ�"���������K�C�03p�u���~�tSv-�uvkg����L�8�(S���u��n��|1�<��`�VZ�� �c�ޯ+-�E`ׂ���\��}e�m�e��$�y�:��3��c�`91�y�Y�I>���5ե�9;e=�Y
Bv֤�|��PPf��9l��pS�iV�4�1-c/A���:=:�
����D���ǡ�3�q@��+����o�y���.�cݛ�+�=�������}p?�b�,��뷰����rN
eq��r��M�xR�o)��S�����Β�;oU�y��r����E�y\�f����!�[���c#�=7):�F�r��6�k��]d�'s(s�� ��툚Jf���ym~ ��"�{�I7C�e�H)�Gq�4�=��be�u֣�e
��Ds�z#D���-vpG�X�N�8%K��S�V��b�&�-d�zs��s�����l�]�����[�F�4�@���nƝ�:�_tM�$��/WS���;;�#K�*�}Ǳ���B]Ɨa׫��^T��q*��H��3:�*gh�:�B]c鼲�^[t�ڑ�O�gyn�U��4'�L�Fa9�7�U�o�bɇ���E�=��<8�*]�u��0�c��Xv�	���o\���8kKwx1�w&|��DvudP�[�;�`;W
�O<�\%>�w��pu,,6Uh׵��r�g^��cN����N�����{�nns8��Fԕ��#�j�A�V���[���ڽV�wE�!GY��-�HZ�&�dlny��)����G7�jήa��;[���bͶ��u�z��g����ɀ����{�$.���ۻ���,"��j]@yE��Xɓ��c���S�HwTw��/Z���s0��*θ+}c0iQ�Y<�Y���J��m�{���jg4��k<|�7���껪.���ʴ�ێ)�V",EQD�D�iX�S�JZ�D��\��2��j�����B�Ekee`��-��TJ(�����TPZ���-�!Q-�%-��X(��1�1�J�\±��k(��!Z�EiV�(�Ȉ�m-q�--��kh��ZV��if9��[iQV�V%F�-B�Q���*�iKV��R�R�R�V���
�b����E�Eb��B�j�W2�Ej[YJZڔA2�j�*�ڭJ[hܵr��\�Km�V�D��ڪ��VT�*5��m�ʊ�!Vؖ���Tk(TkV5(�e�j5)kUEF֨�F��[)E��*�jU��ZVQ�ֵ���F�h��2�����)T�KiQ�ЫF�����m�,��Q,�)h��֍����1-ˎJ�7)Y�--�VՈ��m����h��V�Թ�cVR�1���eR�#S)��Dm�j�y���߿�����/�)�éo%�k�I ](5�u�V+�t��VK�w��#�d(�6�rɔ�g<��F���c�/�类�k�������~P�
I�<��m�X)8�Ԭ�&�u��f�N��.��&�R|��{�a>xɟ��d�?L�IY:���%d�����������:���\��{����{!��d��ˌ��>fr�ROu�P�'R�5�0��u+5�p���?w�;�$�/2�|����I:�&����'��\8��4�ϻ�~�w9��f��+�-R�x�l��Ch~d�je1$�3_k��I�ћ�q��Xy�Xu���{� �u�;�'?2s��d�'�������'���Ưz&�k?���0����2O����V2�N0�:��H|�Y:��1��N&��٤��7��'=�K�8���=�w�*�9�:�9<��v�ڿ{��߬`��|�}�~`z��'{a8�̛;�B�O��?d�	�Y�*N ��[&�q�����6����06�0�g����'_RJH�u�`�:��}���+���Λ�p�'�'9z�L��o�d�N2x�O��!6�2js̋$��k$�(L�͡Y:���P6Ì�Maa8����1�,��f>G��=Ƴ�|4���W߄��㯩8��9��痺�z;{��w���js��à����e��ey�sq?u:�Q��C�uٟy����<�C�����L��.<Xgt{����,	Ϋ�u���&s.�b;�I�2��ei{��8�%K�>�Ow�ۇQ��1���Gx������5���{��IY��*^#�;��i���NBz��'�#�uv�rs��d�֟/uw���fu�����`��H���6S�vT�������{w}�.��K�c���'�P�E���:�Y4�u�m�u�厫�T�Pkҳ���O����R��������S褺�y���z���ً�T�j�mn,v1lOo*k�����꟒�gK:������ޝ�o�U[�k88��O9���-f�y�2k-�����eVl��Ƕ�.86����经6��;�2_�2��pw-��S��K�}+��|2�@��K	��u�9�����v�J����F���G��Uה>���W�����|���[�\ȇڀq�U�Z'xqޅ��̲��fVi�q<
q�c/��ǘ�ߣ��r����f�"S�x%��]n��FvI}�:S��Y�8c<�%���U|��$����:��wK2k
�c�9�L��}�Ǻĳ����ǎ�a.v6��Ve��	�y]���Q.��Gɿy�c'��w% }�L�[��L_��6Vķ��[{�[��\����}�$�/oFs���k���N�)�A�����8�l���5>�u��i��K��q����y�Y�t#X0�f��)r�s�᳇wҦc���u�mv��b��N�� 
v��b��5[��fe���)�^��b⊣�qfn�ɺ�ٍK��'	�Mb8��V��N�v@7	�D=�$�v�t탹���iK�}��W�KY���vk�������3����d֌���2L�Y&r�bb�#�S���V`�� �0���t���.x�G'u����lW��,�8,�ٝ�3k��:��y]�6�In�Gٸ�*�.r���|_�UΛV��W=��V&��'1�;�v�M��^�o�~�ag��1��1W�����67Ƚ���b�p<6:e��'�3����@V�_gc�v���������xoN65�^N{���Yy,Ce�+������~�&>�wL�P�jk�o�Of�6@�g�\t�v�Ū�h�������G��lz0>>a����ٟx�m��g��f�ng���L`�a�!��w]��r�V�0�ߏ�eg�᫩,{�1c����Y���خ�Yk�wkSȴ�'>�By������Y�;3�g��X�� o۞u�N��R|���G&ŧT�c�R��׃�8♓�3�~�(.�_"�����t�H������<�gCd'�:.�ћF��GoU8S=���;v�Z;[��u.k��|H�H
��CyRꅋa��c�ȻU�m�W�W�Ul�C{�K%y׮�|�v:!N=�G����]xmG�� �D�Z0���w���P0Oga�pI�s��٧q�l�Y��D�vi�K����e?w:�%�K�G�;��nl�:�����%����]}k�+���ҳT�u�T����G?.����x���; S����ʻ��Ҩ˼Ux�#�i�=>�!f
���t������ߌ���s|{B&+�YjgGr0o=���^�v`h;yCΥW>�~��>hu�;gs�p�V�'�i�z1r��r_�	=b`vU�/*�zf�w�3�ҙÍU��\�Gv}�O0y�1��z�p_�7���'g�@��u�x7ّ�����UL�ח{�[�CW�K��08�5�dk>b��\��_Is�6�nτ��p'1f���Ƚ���GHÉ�8��}�dt7O�ej��٥ڰksR4��m#��W�*����!��*�Kʓyd+���d��+$�1p�{x��N�edfY~U�%�߮�뭷w���
[��>��ʬ|�ewP;�'U��/Y�ڷ�$�z��Q]ja��.�g�+���ǝտ�}�����6��F^���U-����V��[�/c{8>���+��Tso�X+����ݽ��#���/�>W� ]����k�b}	��hs��zk4�u�o�?���X��hr���q��~�i�m;�ay�{�n������ۖ��Q��<����ySVռn(��sMj^��/of_@_+-X�\�ǸHo�c��WN�l��^?`9S�{�b�J���)�'v�N�>�ω� �1y��LI\��#���y���k.�"��;�{�L;��+>��C��Z��ty��ę�K�<�+���.z�,�X����5nH^�vv�tv���|vBy��]���}�>}R��!��]����U�9�)�u� ��x�D/��y�9����J��u���]��ߎɛ=Up�s�Üj�Q�B.�����T����.��=i�|ַ"����T˧]�ȳ�-FS�F�����
.m#�S�,��|l{�b*7+��ܺ�������B�ߞ?SykZH������m��ێ	�&�ڡt�����M�l�մ���'B�gb
PVn�ӂ�D��9ܝwuC5���]�$�!������{�f�|�~�M����fl��r&o*�U����ۃ&xn�ۃ��,�{PWm{�y뮾�}3#_C}��~�����<�,�g{\���t�Sn����x݅��h�O0o��$hClf��QTx��o�g���Sk�& s}fvUM;���?v}��ʜ�&��.[�6xM�����Z���7OՃ��ys9R~ܞ��;�&��,AX
�3�y>�>��w�Q��Nuc�����sfr��+w���+{�e.MR��s�'o:yL�/]���G�8͏O=�7k��d�0q���9l�y��u��/�{ [� �����t����>�A�e��d��pιG���[�w��4.��z#�r����2uNP1�U���|e�`���+2��;*Z�h�+���`LIX�����f�������l&F�=�%G�;�N�� <����XӘ�sS�{�x�b�uȺ{�t�8{�U��jȟ�yF��V�Ӱ]��=Y����eRp������[���!���s�T�4��FjZ��g]oc#�Rˮ���������f�8����痿���Xo��1�up�~���b�)X�Z���3�{v�հ6:��9��>S��%������;������{�fo��}y�SK��;γy9�����|��+ޮ��1r�:�,�s���򬷙y�]�p��D�/�rj�����=�b�$j��;�;lЖ�����,�$�tBs�V��?gS`&瞃&�f,���$εc,�p�k3M��Սy�bW�d-g�Ϫ���틟����6eǳ��Om��t���7�O��� sjX������ʿ��yy6]��W��/=J�e�Ǣ��'g�(�6�8;� om���S�+-���;,�Z|A^���"�R����9��\�1���t�e��Ry��,\�޾֫�p���=���ڴ��?����=/~}�����ǧæ��Ɋ��]Y�	�g�n�er8�P��F�PScY1�r�yV�E��s���>+�T��^�]�z��g
�����F`�1�����D:ޝ�1Z��u۩�釐Ǘ��5�]������TVi��/Z����s"�ȁC�wV���f��� |>��޻�B�o{�+^� \��fܛyPv͖�6����=�}m��ZΩ�OU�~pˮ=՛>�u�e�y,z���2�@��K�^�F��ѫ��!Mu=nS7j�}ӽ����귇�3���ɫ�����٣�d��>CJm�ky��o7��k��~yaY��<+�����F�D�X�
82Y��ьV1���p�Ӂq�`���{���8c��S��i�3�j��ng�CϽ+t��ĆǠ���:3���]��R����(�gpN�n{����y�nh��}�I�A�[�����!�oh<��f�(��L���w��Y��;%�9֮���ꦜ�I�殭�qy���ƙ>��S��+w����Qx�@��������75��)����������9~��}=�󏗵���"���n�y߭�Bt�\��q�eBy��hK����*�-����G��>mh����4��� �� �+-K��4�j�t�Hf>����Ƹ	��@U��[B�5���X�U��6ݡ�s�s�2Ƿ��3��r��8:k�@>�ڦ��C6�>�.ҵ|�W+y�<�7�W6��|.��ﾪ���,Ű���������\�Z�rgI��tN|��IΪ���f��j��7ծ�q���{ƶ����`�ol|��r�{1ߦ�<�S�sҶ��.�>���ۙ�S͈����b�p<:f��%�C1|�dw��x�K�z��1�kp),bZ����~��H�_#T>���a;N���/���)ŭ�;Ҽy2�����Oau~���G���핃�~��o��y�#�}������^�1$IA���J�\���<�a}���[>ng��)�w�}��Ң�
�Oh�z�����)t��{�-�(�������9�����?O9�x�����ڷ���јߑn��=ĵ�����ά�]��v��=�t�RM���Ls$�o�����0�uۖ=\�%�ʀp?R���	�+��t�E�^uG�犖*p�<�иN�u��]���yWE^���A������Z�Ц�7��M��7;
HQ6�u"��j�:�j�P���j������R��J
9G =�a�D�U<�+�˩�ˢ!�Y��!����v�kE-�}R�p5uΞ���_� }���8��5�u����Yц3��K]��uasf��$�d3{�	�<{��Z�'��w8�ӫ�&W�Gh,Q�	�m�Հ�<��^�T��T�)�wi���8��ν��w��8���;_Do<9a~�u�q�ͮ��,�?ퟚ����j��<��d��:.ǁ���R�MЏ%��/l�ik��!�J�~ؾ-Ɓ��T�I+jIU,5%V�hu?�u�u{���k��j�Y��}oֽ=u��o�dk�o�8/ü(^Aw����N��0ZK���>�x������{d�]<؏I�s,��F,�[������ |'�>��s��r��UG�y�T�ٹ��=K�"4��T�ҫf��F|�]ы���l�;+�B�0��V�}��t�,(�S�V�CS����Ϻz�Q�K���s������
�}Otd����i�b�h������;��]�[����^��"\kf�����]�՚�pg+*�L�ǤV�V-��7�Fk�u�Z5VZO�5N���8&��;;h��=���(�)I�]Yke���-�&1����9(�t���5�3r�N��Z+)�Q�逹�<3���f���r=5}��e��vd��d���*��ΛO�C*����ڱ���e������ڢ�s*l�guL�ע�N��x�]�3��4h<GV�GJe�\*�6�|;��K:�*H	����C�¶����Ja����U���Jov;�KċN���8�� :�\|��t��\(��GeeՑ�%wbv�+�[�-�#��.����a�©���Uۈ9aZ��1P���H���ɀ��3{����ԋ��.��(�3��A�nՒ�*�-�l^-��i5c��n�Z9��k&k��b|e�<��δ�g}yt�ӛE����i�k����X�i�a�6�6Ƈ�X�z�]���y�Y�y��(�g�pZa�j�KPc��}��G)Wm޴�t�U(�w	��M.^F�	igLR��s��WU�G��{E��\���B .�7�5�we�# 9�T=|6��}�9���I�t�af�:l}]�Xs^��1�so9*�[�b�Su��㠳vhlT�V���d}|�Q3)��;����4��wZ���g:�l�e��W[�����y�:��A� �NF�CUu��; �7(rC+q`Uu:u���1;\WMN�����fj�b��BΫ���6�r;�"L�3�o��N$q7�*Y�|�v�]Ym���v�4p�$�G�D���n�^o�Pf��|�77U����E��jx{kR���6��t�.���Vwd{�1YѪ�����3�R��\DVe�ӄb��Oc�e�,�ьE���������/��1�5��f[�{��Ū�x9tԂ��y��F����j �x�(Ҹ)�>D���&+Rq�2q!f�˭����v����i�ZhL�
��]�]�/U��hbuE(X{�IC��F��j��q��2��^���\NV��;�r�sa��Vh�|(�BLo��ztέ��F�a����@����t���s`�������-s�rct�������Z��k]-�M�Avx�(q�.�.�1k����]��Dpe�8�+�;�ƽ�Tu.E�<��[��N�5d�`rCD;ګA�0�f��LU%&s�٫waUn��ȝ��˳��Wa��rFм� :�g;����yp>�k룧�SrY�������~����gU�j�kC
N�-�y�»t�n�Y�*!�^�%`���g����Z�n�媄k�f �����=N��]&%\�5��rş�Y��'|�r4{�ly�¨�k���ѻ�}�ي�_;�[�G��ռ�d���iY���n�]�<(� A?*D嶋Q�k�Q�*VѬ��m��j2�c`ԫq��c�ʖ��Z�U(�Qs1��JزV���Q��*X�e����J�J�aUV��J��KJ�EKn\0�J�Z�[kh�i���Ab���%LQqɉic)[-�F
(�҉c,i��Z�r��E-�2�JŨ-�R�iQD�Z�5��iT��&%KLr*ԵZ���+�-jJ���C��-E��8�,QB�̸�ZZ��J\pfZDd��q�Ek�3)�����Q�U)h\�KlfD���dV��T�
5X�D�\kQ��eC��0R-eZ�EZ�U��+E�Ae(���m�ڌ)F��j%R�UTR�Ke��r�j)Y*
T+DR�V�kV���X"�f(� �~�>$�!N��s�L�`��v)�;��WW�3H���ܷ/��[�B\9u yq���\z�=��m�V���C_����}��:vy��������:h�<��S#��5�Jc�כCo��?/^꽫��A,�Ѵ�u�{���/�|���� ^�0�j8��9۽�̦�W)L���ono5u��vg�[�c�S}t��o��>nZr�WO6�Z�[ۮ:�%���os����i��+�|6<ąC�w]���W�o$���Ǜ�q�t�B��x������}*��3;�v�c��ݵf=��%�\�9���GWe���}��We(�Նm`4�9���@��x��Zs����bNH	���Έ�H���&�J�'~��7g��P���_o?c��,��Y;=�xx��J��2d�nm�a<��7�^���R&�3F����ث(�b��v�yO�yԹ�c�:�Z�]:������u�>��+7'�T�=X#��m��Voj#Q�DE��)��b���+8�Р�<kxt�b8�G7��Kr�n�gfa�²Z�j`�}�V-5�9���R�Z�]�^zl7|�6ܹ�O<����x�4�[�/[G�e������j`��=���6~�������כ*w�{~tZ��g���XyT�u"�,���f��E��\Kյܵ����F�x$Q�m�����-����+-��Uc/0x�s�͗��M\��sK�[�w�I�c���t�e�T�̗X��r}��&���wY�t�d�K����{��5����ǧ�5�f$<)���5����R�@�xb�\��\�y{ ����ϵ�T�ڻ�$U<�'P5����v��ng�������6�A����xI��Y��Mg�<���F�V|��������|�Sڳ'���\5}ẇU
�vّR���=[�'/<6G��Ms�>�<�fP�4�eKO�w�\�(Z�ܼ��Ƌ~�C�0=����u:{�������zh�8cD:��cɽ����d���|᱌H}�:N��k�7����Ex�v�ÆmdX>�6�������7��T�T�7����k��t��ΐ�]v3���sa%|�SJ��o4ƽ�,�*Nw�����8��߯5�����VsZs����&>Q�ی�>4��dPvM�]�Y�b�k���b�������]������z�n�1�߁��_����ܺ��������:���7�E�%4ma�lw��^�(�>	�����x�@떇:�uծ��=�d�{�p��{��$���e���<̭����;�<e	t��s�#��S�ɹ�P�n`ATLW��s+�u?(q�lS=�.�h;�CY���A�L9����r�J�\���SM"�~���l�\�3593�zİ��-�57�J�|�9��}C#��{�g'w>�4�!vg�1̏���8/��yN鷡c�=X�c[�n9�y�"��:�_��^O�R���%��c��ѓ��y�n���6JW^n}.��ԧ��{�qIbZ����{���?@X;i��΃.\��S��M���������2_�|z[�>UN_�_�1� ��wz�5�����̯7�9��}^��K�������^>�\=���v;w�b{�=���f�ij�j�oFr��U�����ç2�6��[S����%�yʘ�7Z�
T��%�Sn�ӱ�Oe�]I�<���M�
���Gp ;1�݂-k;GX*�R��� �5 �k��|��u�>���P��W�;� >���Z#]%{w�/}����侒�e��结6��<�Z�9�����da���%�ϓ�>]��ss5~S�?n-ו<�Y��t������"^����������pr�9���:r�&���xc����sJv�i�˝�w�hrڔ~u:�ew^טu�Yr��|tM�Du��l��Kn՝��Cɓ�����α'�����	��͹L��P6KRsJuwd����b�h�_����?��Z���V��L^��^p�w-�Pd�;B.�;�zú�X��S�rʦ�H�V�h��vΞ�_&��z���X��b��A�vB�0�Wy�<�{ykY�ʝ.�3��a�.���� [�|f.B���:ԕ�l��Yeř훭�[���+�3ϯ ���y��]v`�}��m�A�;X�<��@c���ov�G�ƄN���N�1c�E<ƚf�n���R��rM�����r���e��5��v�{�JbX[W���fJT�r@�銭��L�a]>���ս������脠-�F�V:�V
�D��Y�2�oa�v��`�\������ZS�I�ms�j�=���duʟ��_����̺c6"+GHӒ�s��^~�e11�/�2��}d��'~������x�z{�2��}ּ�7�->;��W�~��q�����vgT�{Tϭ���v�]X6�~��I1�{>z�v����uc��:���!�������/>;ᴝ�~ ٭;3��[�&xB���o�<�s� Cؤpo��X�~�Zb(�Q�4��`޴��'v�.��B�;�۝ C��3Tq�Q�Ҷ�Q����R���~�u��*`Y,�9t�^���r��-�|��Cu���[Mx�����q�+�+2��;�eC8�׬W��Æ�Wc��F�e���tW��}��t�q��>�]�Y����d��~x�v�.�:ifR����5�`ȷ�65l$�3�xN=�,�GF�;vxx�e1'k��pI՝�����O�o�T���U��^̧��A�#Xv�vZ��1p;���;��='7��,gCݔ{"$NVM���˴���\]�%���J� Yn�2�d���J�b>�y�i
J�+�OX˵��w�]��d�Qg*�3��C�������ryK�������2뛯i�o�!��� ���L��N�O�׭��e����	�>��W����yv5�.M=���Ʋ�yc4O.[vۆ��]�_)G���mG�J�ϰ�ǗSϓs�L�ј�����_�l���c�owzc��ML�����^~�����]"|�ͦ*�t�ܼ���g���o�93���U�\�5]�B=�N�raK@��rM�֊��������Clc��3���[�ʩ؃�9��G^��_l���_ZRL�����E�u�Kb�M��-����{*��x��ټ���;N�c�}mn�L~�vE�Y��og�3({~�b��������F^�;9�'���<V�{h���՞������9(<K���
��6��8:���q�+��W�mG��0��������>�w��f��،ï^<�J�����Z��Xl�5(�}�X�92R x��v�Y�s�����̀0��Bq|�Rn�� Θ®���8a;J�ݷCy�>;��}[��medL��R;W���k�6>��ЎټU������W�75 �w�/������@o7J9��qE��o�eW��]�F�[sv���u���U��������#ٮn1~yaY��a�ae@bJ���َ��%gL��V�7E��׆Cy�S��q�����{�gGyz[�@���xۊ^�s���&C�+s��ĕ�(%��tݯjy*�̩|��6�J))1���!��G����ރ͛�&�)�u|����f��>��G{��pN���|�Ŋ��s��=�M9�*N폦i��~)ծW/��ߞ�|��i�r��2*�%� {�
���C�o��ѡf�p��E�����YK��t��sp9��{��]��n��aй�tDm�m�f�^��1�V�"��	צ7b���&p�_���˽z
B��)���������	w���1�7]�l�qF�6�8/�z�gaN+Ʊ,��#Ƃ�*�~iˑ����t�6�>���N՗
�O�{��y8�����+y#tf�sl����y3,B��,�zRȷB�,�����x��c���,Y�i��M]$P�:8�	7�nhU�U�ZQ<��nP���W�W�}Y�g����~�����=/������S7�׺Ix�0{�س����Jz����(?|��\�ʔ�����⏽��y7�O���R�"!����׽�y=V�}�`�����*Oٳ�����ض'�$�Z��N{c���c�
s��8��}�v��q���?Nܻb���Y�fHqvΙM�Rk���'�/��3��!�:��~����KѻV��/a�ux��Ƚ1{:��X{�p�1wH������q�y��ķ�G��(x=�+������*���S��a��(^�Ǹ8{#�K��z/g����^Yڎ�'^:�^P��z�V�)�r��J��]�N$|1��,�H�q�;�з���t�^ǻ�:}N枭}WQ\��3��
��G�*��d����'3ą��z�Wzy^o9���~�z �x��n�����[eEf�&a������H��ujy%}y[]n	& �2��W{���T�f��"<�]�x�'`��_�^�J�4�:m��ȠY	:��݇�)+�	�W<���6�|�8٤���`Ī
���Xu�I���B�=�Ar��
�S����7�}�۬>�-��Ok
t���  �Tx��\��/y?��Qp�$=9أ-n��Ҹ��e��ĳD��JiQ]�^;��"OckK]WN�*��CVڞ5
�ǅ��7$b2�d�E��y��/pk���I��PAn�3�t�+��(E}��a�3��t�2�śN�FC0���Չ�	�Nb,�����a&���2r��x�d����_k�\���UŒ��}N_��S�N�{��u1���\L�Z���}�	":<��w�1·Y\D��e�����vS^����֦���3�-�M�
|���C=�&����$]��
�y��(���G������t����K��@h��B���4�/�v³F&�z��2�7�ȅ�=�%	�zp��oG����8W��,�Q����>��p�<��^,�����3�\�_��<�/m,�p�ӾJ���`bW-�R��cF
�*������+e�2�����e�2���O���}/��q��	�t~�i�+���Y���Ur�Ȏ���#�� MF�c+7�ۆ�k��|w�ٺ�r�J�fć��&2���"z���SNX�9��^�
�Je��T�&�G{]k�\!
��lWk��(O�<���Z����fuA��uK��gp{��͌�xq���GK�Z���u��o\�Պ^�{��>R�3%CI�-�;��x��k�0��Ҹ�KH��ŗV����Cl#�N]���ΑR�񝂧{��f�i���x��6���Ԭn�!V}��,�,���;����g��4���w��{�Uy(�S-xe�e����9c5`�k;�y]#����xU;S�V��t
�;��Z�qm�V�M+�U��誥b3�à��B�V;���4�����l��+k�ݼ��t���$�/{�dU��l�|�՛(��x�f�?{յ�K9�=���Jk�\5��C�whi3�ȽA3;يX��yz������[Y&1��g�m;����ڞBZ��"S�@��Y]L�P�e��iL�Ɣu��W����:��[T|��S�_^�	ĺ�~���r�B��I#�:�|5�z�e��(�#le4Zc�v.�.OVk���s.힟��ӑC|���v���a�d����_�,�81,�}�q��C�������|�R�к��{����ҡ۞�0����3��.��Jf���W�w?.e�?Pzk��=���F�JG�<�t�VA��鑛�"���<N��芀��Y�I�R�V���X�E=�\P���o-N�7E���	�vn��:[[&Mc��Ͳ����&�G�'-]\���cb#3��v�S���e��ql>�'&u��F���<\�'	���qfu�U�Z���;.D"���)�EGl�f����D%�9��V�hy2hG�W%zP�fu��]qǼ�:�x��r\L��+U�ƜUG�T��u���I*�ൔ;u��x���$0�=7���xeIJ�l����%u\�Πڅe�sC%gK����-�9�G!�K�k��i����ܾ�(��Xq�l�푘������o1n,�x�G������#[�����j����NKrhY��tڴ��b��>	m�T$}�uEH�9VK��q���Z8���0�m�Y�R�a��j�boax��ܨz����^��Z���\z$![��V����k�'/U�뫢��]:�ᎎ�
$آT�&��}�N�*�Wuٕ�������E
��/ ��+�ձ��� �l��F�KΡ2�ʖ��Zv�;<	��\�+1����h��̦��7���"1���݊�X��0TG�D���]�ɏ����g��W�[=7�O�tזS�V4=˙��[�D�7]�us �xC��fMse_T.N�▫���u��j����I�B����YעY�As&��z�ΘH��O���j��5�G���h�SpoR�;xQ�E(�m�w7~fD-��������M�Wg��voS��p���0bO�݆a��PҺ!o1u��4qL���(�r���R)�;��f�u��r\��SE��!�O���i{&Ş����r�z�5��Ծ��7u�sz.��,�Zm"����V{m�C���vk�U�a�N�\���Z8c_n]�CW�Ji���H5�7�Wj�oJ=}C��j�_<�,@��7��1��(��6�cCVL�[Q\,��V�ȥ�};�m ��Β��qF��oy}%��/q�̕Ռ6q<xܾ�QSB��V4��o�	#�i��]F�����c�\�7�a\(^I�#���A�]��9�_.�MԼÕb�e&�qC��~�5�la=��3:�ɅDe�N�+^�W:�Ps�tHUp�W�3�GmI2�5HR�	U�ސMWPo`zWJ�2]�Ś���._e��):��=�)��&��,�>|-�����p`<$A�6�fD�n��9P{��싮����WM�Z����Eg-�z����eݷX��!2����#�o2�>nt��44
�u��{�u�:�9�V!�:��
u�;��$lp��ELVr��k*��ě��^X�k'K�.j��|ťG �c���R���K�eD��Z��r{�fލ�
�T�.��,��^v�_�[e��PGR�~i��1y�P�Ukµ��F6�m�V[b*��Q�6ڵ�[R�ե�ZZF,�YV�(�b��b*Q-����"�
�҈�*��%J�2�* �(�F��m��X1m���Aƈ�̭�,km�Zf\�U6���"²Q"ʪ�V�)LlX�iJ���`70�TPb�[*��kj5L�
#�`���1UQQF��Tkm(ZԴP+E��ZZ5��E��"�U����"(�mh���am�QK[Q�X����Qm�V��Ȉ,)i�imj��mQKh�)[Tk*[F�#[U ղ�
��QZ�UX�e��"Ԡ�QiAb[[V*�� ����X�V ��R�iQ��Tm��[b2���*�J�*T�"T���R��cmA���	-��R��V�)P[mT����2����A����+b*�+J�DU�5�+B��D����O:Q��L��Lv�	#37w
���>0����I��L�*��[��\U�Ke�{r������}���}��W����*��w+4�SG�:�q'�t.L��E�^w���Y��=�Ӌ������F�M@T�ꇄ�u.�,v}���;ҵ-pPO(h"�Ǜ�S��Q��˴ߏe@��Lfq�<���{gOM67�`2��/�u�o�C+ݽ��6�&RF���.X����>Հ
��� \�2�����`�e;uG3xT����_�[o1�����Ď�]��cgǼX�/�Љ~�Z��}z���B��4��#l�Ҷ���sE���r~)�3
�N���V��g��1߭�*ʇ��.79�(�Dn�{ޑF��L��x�M���&jxT!�a��C�9sWh�dk��dj��Y݋��Ų��_	�Y0�,�J���d��I�tL�{�b���Bx[˕c�9[�{β�i��΍jz�X�U�(���h�/@�Ox�u"G�~[^a�]�Wk*Q�:yl��^Z��a©Ao��*���� �%��C��B_8���9��0-��D��4�f���h%�2ľy[kJ���md��*���l���m��:~�h+�a�u+�L7��~I7վ��î�g؛C��͝���c��0=�&��36��3WR�2�*x���T�7�;��2���Wtx�� | �%���i��F�����o�9��Pv�OR2��P<D�	s]�P�w�B��g��[�Lj��.��y8�\�z���-�f.+f㤄ܪ��U�X,�T�uE��j��/�ы;v?ik�ӹ�*Cbpb�f6�zŤ=��)ˈ��%����Z.�Ea��:}z�F@o�� yKI�԰ʼ�p��5lu�FlA�9�i.��3��ڇ%�Y�������C��7�zL=B���km=޵����J�P�AVtyɩ3��JCpc�<%0i�wT������<�Ƀ|���kv��׸�F�"ld��?s9c��n�f�6�[$��P�Z�0vZ���TR��Z|({E�T�:�k����'9c|�+5u������}p7�8���3��\�t�j��*�z��F�E�j"��!'�r�7K��&�HJ߼���`�"K�;�[K�2���t�Չ3N�
�>���и#�2U��]�K��%/���)k�B���q!�e=.y��=��z	��2N{�Ȫ��-�F��]����.Z����S���Ƿ|u(@��Y����=��hU�G&�Lp܅g���R�Vܷ3��t!N���[�f�cߐ�o�/8��j%H>�oN|���uwo�	KXygB��+�U�V���)�Ō[	ط�r4<Mnqvy�E?�|��3!���q῾*����j���+J�=o���
�tL$��L�LB]���6 ��ϑ�=҉����Z4L>�5ק�3��`�ţl��VYV�p�Z��Nyz�t�ޱ��5-}��KE�������h}W�a��j��u&��o�<�����������y��6�E2��/�K�	:�(�|��#���G�����z�wu��̽�w�]ǚ�v��^Hb���	T�n�E	�к�{����O[#C�� �=g� �l�ӵ����
g�����B&�b9�E��7$zm�Hr5DfjB��V�WlkP�a"��f�]����E}��a�����җ^/������K�W���soH��Àr���4�,�x�d�����k�xk�@Sg�0��4�s�U�zS�ϧ��v߼7|w&���!�A��ZHWњ�I�2�뾊�:�B,�u¤��ز�XfOCc��n����8�~�mn
z���TC7�&��1"��%z�z���]Gm+�Q˕��� �����|u%!�����:tRm���+�GEn�f�yŔ6��/2i����"b_Xɔ0�U�$t{"���Kb1l��s�"�L��[Cl���O��<�Iugw.�M�߲�=����P6���w������s�!i���M�[�Jd{�zxR{p;,z�(p�F&�z�uN����*7+���+�\���V���|���m�!}�0q/��}���+�
�^+��^�q-
�c`-�_��k��R���.�j�)C�S��o��=��h�[����`����QZZm���~g'oW��2�!�;�B�85�~�i�V�ӄ����֏x����Ƨxm�)w��lV܇̎E�l���A�����Ϛ�,��Y���i��`���P�Nd�{�����U/>��&5�\��U43c����x�=S�����U��B9\���;P�*l�7�ޛI��xc�YA����P�����X{����
�����P�Ɩ^p�hr���f.\�@,��r�M-��76x�|f�����v��,'�EvK���y��e�Q���1%�Ҷ6)5����8�x�s^���J��Dg0���.Ys����b��K42��Cz���qq{�	����R���={�><֟��[ z�����G��1�M�Lm�-�ZAN=���w��V�=ݫ�l�b������^�zNӏ��u����u�}W�t\���#���5��P/iZG����[&�QO��h��5V����j��)�]Sjd�U�e�4*Xjsc�m��y��_ﾯ��#[�o�Pz�䊽�e�Yj��L��_j�W]L�P�fv�&-�(y��J�Lx��w�8�7y�S��^:nK�7�.yx��`�����q�s �9�޽y���y����\�Y�`n�#:L�Jr���5��P��Y0�6I��I���ʪ�`_ZpC�}��3�3�Qy6d*+����FܯD5L�J�lO]ԭm��h�eg���ή5���k��hu��/szR%���������Z������v�Ie����M`C�]ֱ]{fQ;ץ/|�T��rV��

�V\Rº�R�#ț�������/}g�'���me&X��O���u�cݯ��]���%���Zس�����#����,k5Xَ�Ub�}��2|����������K�������ga�X�����ٍCF�_{���[�فk��	W�1Ғ�f�?��]gw�΂�0�x:�g
U��¾�N���V�2���y({Gر���\�D��B��oE8�5�e���5�Rxא��\���L77�ƓӧK���*B��x:7�,5�Rz�����\�[��ܙ���)la�����&�5QZ�Sެ�1�v��ۡ���h�8 zOe+(�u�����r�y;�Z�=7]l�U������������b��K��\<K��t� �	�C
�AÁ��+As'�qt7�Pc��SP�pZ磼=��l���e(�Zi�����|/��V<�q�d+�Q�I�&ۼ�Ju�<x�{�G�=m����B��Ċ�@�%������(�b��K�pOq��M���ˬ^�Q���[ʮk��q�T�����Q}�\��j ��;-�Y��s�\u$���w�.3�ێ��][:�9No5���Ef�L�(X��X'��@��r��=����O`��C�q�I����<��h9[\&�\V��J$�z_��������I���.ψ��8���lW���ЏA���P�N)kG	P񒲧���t���t��6>Kte��4�4�X*�J�!�3t䧿7�����8�{`�u������-�:�] ���ꂚ�w���J�y�b��I�����r��Y�}��|h[�7��~^��)� �ݰg:$`7�)��Px;-bg�pST���7��kv���go�uſ&�*�)����sw��;�ȆL�\OY"�!�8�
xLC��y�øE��4�v!݃Nfg,�Ϝ{�4B������ز�)�
��o��;�.9[�J�=�+olV_*e��u���c����uv2��|>��)�DRl���|�]o����h��̶I���z�D;p���X^쫮M���<�M��m;�B	�ǹ`�V�A�&t����WY�4i
���P����hW)�H%��c�&�����ۨ�x�_$!�N�}cbUa߱�id�C��Pä���vä��zW:s��/���f&Q.�N\�K����6�s'�`�%����zL�y��/�}�o��|Ǌn�|`���%a��8T} si{�!�*�U`�n�W�\�J�{J��M��������O�J�(b�Xa��6������P[G�H������%\���V>��n��w���qσ�Q�j��\����?rM5�X�Е��z�j0��w����`��{}T���n�������*+5�3uaupR\�o[^�;]��b��}B�f�"�W�?��Qw����Nh](��mhc���>���}q��z�mt�藸0��-��aP�A^�� �a�:,�#q�G~�r��x���u��1�M�Ij=�i'}��<�p�#�»���
�բ@�k��NN��ʽ_;͏�,hm�t�X�����������xD��}#�yH�U�r���*�OpgV��*��� ���97,���Eȴ�/(t���?��c�ik�� V~;�r�֧��h�a@�$��T�k�#}ƃ����S�c:.,�z�
���W���t5����q���\`�|��A��"�$���')r����z�����#a#O�B���]o�y6�r����]�����C��뤐��v$�|.�!㵇r;��Y�	}#���
V�s��r�БB���h�x���uD3c�Mh� *�,�;�޵�.�q�ͽ��+�RkY����K�tB��]`�S�U��v�
�f�M��Ӛk�S�%y�Cc����u�(j�X�E�����B��`�_Ab�\L�!T�ĉ]�F����ۙ�Q����k���/��jF�l+J�X�)S:�*r��� ��{���3�{�X)��L}{q���՜��
8My���K����8>��{�M�E��@���q;�o�Y��_��su�69���;[��0�NB��P���WV����;mݬ�������vp���g�:��J��c���=�h�N�Z0�͚��Km��2��,���h���c��;��G_$���h �|���,�y:<;6���)�R+5���E�X��U�"9+�'���<K/�S��w��W�������b����H���L�Łʌ��N �5`�?4E�)�9�{f3w�	�+-
J���� �,	{^�*�8�_��:'����|����N5���l��FF���	O�[��xy{+@o�-F״�6�R�Pd,�A@������g����Y��懧�R��u��N�z�<��;<����g�m(�<d[T�{ZB�����p�}��� �����<�Fw�5j�j{���Ϝ%��v��H���./PL��~�K�S׸�p�۪��yn)}�rL�׋�>����Ȳ�!֯���@���D���e��3;)��gy2�6�z���qw,��e��SEĶ��«ՠ)���nDU!A�v(P#ί�5��'f�M�9��.����rL������B�K�Sޅ��U��kQ�P��Y0���$D�Vrow�"�x���ڝIe��@���>��+��]pr�!��+��pS<"�6p.�]����2��n,d���
�xDsǆ}fa���gC��!d��t/I�����C�Q��N�kWuI�u�"�%z��%4J>ϵS �􏃩w�c��U��f�bA�z��:;�3֘6��*6��Jj�z�ڶ�f䵏r�=M���.��9ȓ[��1�P#]�n���Ȭ�5}}b�e�s2��J׻|A؇�783.}�[����[�}V��L1��,%��{�I�D7��1�N4k�xW���Y)�;A�<�Es������5SV�d���xPY�?�α�K9N8�xgZ6w�U^*�)1�S���Cִe�q�!��1�����z�� ɜ� �S��|o<U�X��x�G�R���m�b�.�%����i�!WY�K=}_��Y���VW��4i�x��C�.�>Ƭ�q��&���ݯ��^[�%�q^��]�^���P'J\�g���+-��ŉ}>O޸7;���h�����m'���N.�&,AX��0�.Pp���V�\���N�Y��]:�{Y*Bq摮�����J6��D�>2�Z=� _�9��x�
ȌLA���s��wf��d�sk�~yt6�g����š,I��}r����5�%X���Bm����f�m��S�(�����B5e�4�{��C�Qi.I�N�\_�[�[#r�b�8��q�;9p�
g!�-��^�2u�Vrg?a�	Aڹ�FX�hG����B����=��S���ϨPƼy&ty����c�KE�#�Ӣg��/��I�`x{���%,mT��m{2��;h씟�bb<s7t��;�n�h���
J��f�v��2*j��m�w�=@ԵM�Qf:�6]����y:f�펋��-�j������sX���D�xb���:u�jre�z�f7�'�:{��:n��p�	�I��w(�����:W�#c���Y�!y>�$����Vs�Oq[7��H:��79Pf���owi�Z7ٗjWk��QA����̾��x(��(�T�*��Tۡ���/5��C��d]�s8lGy�e��ܡ�3�L��i;9Vj�]@�A��-b�s�32��� ��u�C�����yS�1oX@$�[���qh�h;}:�m��!�10�#zW�1R-=Q](3N��\|v�3S�V�(%r�>��$��0`s�3m�}�NDzM��f%J�f�;��:�`�aiXC�(�Z��I$`�5L���d��9ֶ����5�;�C�b��RM�O-�˨�	O^`�	�9�;93�EE��#<��p-=�.Rx^^������`�.��[XY� =A�]���ZV�&Nkͤ�.��fP<�,foX=������ERudX�����F��a��X�v'�"��ͱ��-�KyhQ���A�ę��Ӫ��\/�}-`��뮤/%u�v1i�]m���md�Mrj�8��y&��V�����J5*uػ�"�ɰc�f�b�9Պw�-�)%t��͋1Wp���*���w�(�j�S�Q���9��'NƋ�W�b���J(�M]5�L{�	��֨TX�9�f�6x�
�[�ve_4�Y�u��9V-�����_"kC�9{!���/����-C�itY@G�/m�Gr�v�/NfK��&�|�OLnCWZ��3JɈ��n�t5��s@"��#sZ�J�3���R��R��]�ۀ5S�f�#rkU,�D�x�b��[��fČ��U�A��W�y"�F�6�[p��kk�Ȭԋ�������Eb}�h�i�x����4��o
�p�*�j[�Irku;��vj�,��}XQ���RfW]�H۬�ԏJ݁�t�RU��\���i�J�U,�A��f�vW]�i��A�k7��Ʀ��Lq=�r^�fc�#���f�Au%dμ�x�j2_<��������Z�7mk=�E�ۜD��4ϳ�3s\J�[�ݱy:e�JhҏjTs]��`�h�+�.��b�Jnu�
pU�^ڌ0{	YO[���f�7��J��Fj���q�+f��7�Q�@��n�5��������O�j��uYt7|�.m�O'����Ґ��L�F��bꂻ:�j�Қ��Yg*���/��CL��ӐV��v��n\�=�R'��*#"&)�B��J��,�j,@+�M�����v��_*zy��A/���\,�TB2?���m^��gzvnw?T�gZP����l�����H==��:h�ٳ��e��������P��R�1R�j
VU�EF��e������DR�J��V�խQ+P+bҴ��kF�����1kZ���il��*�ڒڶ���F��ZԈ��"���ұ�Q�aV���-�UTb(*1TQQ��T�AD��Z�(���Z�%�ƨ�+T�,VҖVYR��F�DEAb��A�m�++T�[EE�ҕ��*�«Fڊ��Fҡm�Ԫ�
�Z4������KEJ�J�k��A�Q�m���Q�*�E�5�Y��֪�*Th��ITjUQTDkF�YU��Z�2��EAXň�T�ҡil��Yl6��ԥb�E�,R���5UQ*D�mR�������U�,���X�AJ2Y��*"��+B�Qj�X��UV6�U�|�\�g�~u��y
L>H���ۚ&̀�����w,*J�����s�͌�CuB�R����7X���s�2��+直��o��b
��?R$�x B��~ج5�د�y�#�1ia��Pr�<)���7�X.�u������d��K��H���i%�XC*��ۤ��G���S�t���6��o��L�{�^iQ��>	؞8�c��&�OJ�g�]f�=�ۄ299��ۻQ���pk�����T���&)|����Ӏ5��å�
���7���+ۗRf������9ȧ�jy/� �{2Į��'ʽ�޷�	Z|1�N�+m�5�f�joRf�^�ݲuo-����(��qp�V�1��1�@h�δY�OR��b�Z�A7֜g J�}�w���a/N��M�P���HJ�+h����Uaю[K�&\=�`N��ȴ}���ٞj�,��E�����0��s%kpWv�A���n$<+w#�}���-u��)���7��-�/�྆�]>J��������%_Y0�yu4�������H�,oY�S���9��D!��X�_Z�}C�-���zR+�U�,�|f�\���eN�ÓXj�TŴ�z���)����ʷ������,�I��>�e���"Q������Uf�f]�58WC�q�k�e��Gv��._E�J}����J�.Y�C��ӥ�Kt.т2�3|��7z��1b���WqY�u�O+�+̝���|Y�=�l��5����%�T.9�M������\fa�8Z��XZhCdu&�ڼ��-�^��7�9L���9.G)Yt�ϵ��=��UL��ƵFN��8��'��.��X���=����X7Gs{*���ς^#I#�h��+柎������BF9�t���c��:�~{��=���a���(���7�A.��Z�S~��J���07�Dݼ+'D�Hm��c{��v�õ
��@��(��3_X2��.�|]{LV��f��*����5�
bW=�8�V<l��x�RУ�)j��^n�i]:��T=�:�����i��i�3��mc�Gy@\R/T���g8(M-�L��}�I�u�@�d�me��ھ|. �X|���.�yY�C�&�^��R(\*�%��Q"@�f��A��.;髆B29k�vY �f{��&W���tHޞ������/uC�^������۹�Π�>,Ə��Y�҇ڴj�X�-��v�"��ħ�`��\L�r�Y���{-�]w��l�wlב��f0t�hve�O[�!�\�s��iJd��6Y�G�Y[��E�r^��'�S��8�h�\,-�;����Ś�au:��I�v�*�#��v(��I�t�j^6 M��zQ5�gK�e*i�����5Y����oy?~���+R��Q�S� ����`y1�*a�J��ᰡ�S��̕]�+G+����[�3q;��o�ڷ�E�m��Jƻ�Ã~ٍx��k�~�i�K���?N��m�CѼ���9/M��2��==�τX鯮fP�GDls;�)Rma�>���U�P�.��gY���)��<���W }\*i�p�<��V�U7�lv��w��ˌ���eTY,�s�K(�l�qߴ�@����P��X'���r��NX�X'��~�z�J�K�iM�i�<�'#�|��K�4P�;��,+�sM+�F)����c�jqd��d�����o{W�.��h�3Ꮾ�� vkC��>!��xϒ\=66):Z���P�8��� Ʈ�����y�:i�/v����H,2%7�@��ԋW
��u3�֕M0M"�'�rDzi���$���w��ϩ8�Vw�L���y��!����V+���̋����<c���5��%�;%C��ͧ��[J
�V�6%ԴMȊ�ȡCY\��������9Sa��r�Ό�_3�r�X=Wh-EE�4xڠgy�Z��8|8?K���-/������:X���7ax�)Vse
ٰ����՞���Sz#��6ƇG0������t��3<�)���#Nh�0l���z���Y�\k��������9��2S��%��Ydt�f%)��յ�kQ�P��&�ԷL�`��[��F�H�ԼR<�^�v��܊D���h]`r�!�1�p^����(?46l�^'���fV���ڳS>?r7��J��n��+�S߽���q'�dV�tA^�W椐�H)�}��ctb�<�0?F�:��N������u���i��vX��^��j��swZ��$�

�8r��K���}��Y�҈^#�aj�o'ہz�l^]Kޑdp��ʻŦ|<�����0�}<L��:��p���u�t��a>�!꽤<�1�;��[o��Hx�UzP�^�·:�@�垨�w++Ԁ�4�L�U_f�Ӥ��Sy��t����)�y,�"�XaU�WSi��Z7��d�bu-a�P�^k�F����_��^O������Z,y@�ف1��=�x2p.�&,AI��������:����U酉�N�]�.K�<�̮�0�'Ǳ,�Ih������k��(��]�o�^Nua��f�V'��y
�����f�^Bnr~��u#O}�ܳ�/�]�pnI�؞�|ty�0���hU��U���騡drk-�:m�������q�-�l{^0νT�:�0���d�42���K����gnӮ�R�z^~��j���n�?�̔�u���93m�T�	bLj�������������;7�wO</����F��՟k�m��hNVd�O���(�$�L	kS�9�f
������.-ԧL�r�&O3rP���.���ǧ+D�kiB��ԂfB[�Z�H]�S�交F�~]�B�vx�Pߛ�ɩ�1�,a�3LR��17/>��3��w��lkS���(�:D�q|BU�T�8��Ў��!�63Ne���~�x�͞I�3yؘ�S<m�T7��jJM$�K��W��5��QYśRf^[��>[L�M_�A`�C�����4I:$�OJ����~�X+��-t)�$䮛���=7�|��3���R�_�I�p�+ÌӍf�p�t�4�Ƀ|����Xޝ8VZ3w���2e{���|�/}�.�����já&��d�r�o��X��� �u�*����!˔�8��8v���n(F-����~E�.�S삮��q�J�/��T/�n�=g|v�����LiJ�d���l$���[9)A��F�09�uۿ\cmwT�%����qV�ӥ�kX��#X�5b� ��㲽�op�N�q�ɬD%e�-�3�w̚��)���Ǧ�xH3�خ��9g���+�;g�{�䗩��v�����X�����|W�k��J�WD�(B�!+�^�B��2�K�s9�^4�-��#�]O{b�~��n�@z�v�����x�r�{�b��]�'�5(�{f�ۮ�^��r~E��>w�<P�y)���`�*���9m���n�Gƪ�p�+a����v���/5���UTn��s��ze��.���=B��gp�,ߪ�#���[�]ε�B�ɥ�[���T#�bquظ�*rbz���_ t�����	AӼ�=<}W�yS�C]S�e<N��./��s�wb�w_DF;��AסyW����~5����	�C��˒�����e:��&����%z-�R��{�j6��v��]@��(��G�u�&��J#`�a��O�����<t/kx�^��|�^#��ּ�����z26u��&���5dU�	�v�2EJ�Ձ�]�=z�'����l.fx��q�g�mv�a�(	.".��aϢ�$��%����7��&�zH!�M�Dj��a4��Q��^�g3�]�s:S�X�:�G��Ea#��ma�[�t�g,G�x0�o�|Y�m��]�ξN���ԧV��������
w������eR�f��R��fŃ%-��d��w=��J�*��XZ1�&�{� t�;��ESg�WJz"�grP4�2+�b�뤐������V/ً�^����2}���+�u���^��"���U�K�=D�|ê��[u��>����8��J�2��p�[�[3�1��q�AWX0�l8)�]����EK캙~�쎋W|;��`3^��vv}Mp�2��/e�'�]�5���X���cY-Ua���?�.w�L���x�՞^�H*a��<r�����S_C����֯6$K�o0���@�[�xKظH<��P����%��;���^��ۆحĬ�p���~�eE�zj��ٮ�u���y�8�#���id�+�>���na�g����'��>40�x�`P[���HJ��B�eNf�i8��:m�D-a�By��jJ+��wo{v��`�+hu���E�uצ��(38S������W>�^㽓޾�P�;QO?{�ò�hᰴ�3�N���q`��.i�c����a��58��ϗ�#X��߯���Z��oF&\x����@���e��o9Z�dj���=[K�'����iN�Y�lgb������ �f�Q˂wR�K���ofkx�#��UXWK��s��K��y1:YVf�6��)ۣ��
jSP[���^pgՃ��f��I�~�U��F�ahG�����$�zllRt���Y�SQ�2;w�|(KW��Ne�tLn�Z�|g/H(2:Y�����,Q�p����Ҩ�e_b¦�����E��3���v���V|�kk5L�e��i�C�v�����_��˼�=�e�����'������ْ���rf�߮%���«���.nDWԅW.T(V���'Z����ˮ��1xI�G��]�n˅�K,��07�%)芭�8P�#�%C���P�6M��2;�2t�[�N�>6IΔ*�MN�v���!��Y�!�h]g�Z�=�1X���X]S%t���7d�6��Tė��i����?l)Y�����fkس9�
I���.;��0��>ݧ{�6��9�/��3�J�L���l鋬
�X���|K�K�-w�)��ʒ�	�xǭ�Z{��(9�a\���@8=���Y�X�C)1Z=�V��F�c-�g�q��=�;/o���xK���,u1��su�$�����V�U�_z�L�f_�K�h"z¾[/WU\�99KE:�b�J���Y�j�� ����
�:K3�B4�kW�j�uB��N�n��J�譇�"�
F5��A�U��٤WN���i�G�Tq�d�k�n��ھ���V-[�Qj�ٔI�U���D΢�[�]��;��s�����I�F3��xz�c���VW�}�4kd��<0�iz�[�[郠r���ʏ��}
2Ǐ���|���h�>3$����ð���u��<mL�g=�V�NwOէe�?a���GW�л��ܦN�`Ly;�a2���vc��ߝ�v��l��g�ݓ�sW
ΕM�
��a�tm�I`|bKG��@�s��E�c׾���^G�,��N���V�Bx��]�>6#^��:�Ę'-�J����&eN͖�WA5�y��~�dך�4���T�2hw\��`�лL�
��B�*'Ib�%�P֖NO���MPE��p���܈�+s'��7%߽"�[;��y����z"=���x� �b��t���~"��*|L�/�X�Z�%��N,�����B9��l��v�g�Y��|��;k�.v!�=���[Ȁ���|���x�m��Hs�P�x[5��������A3�G�P�暈C,�}%&��B:��B���ݣ��<3�ׂk�T��b�qوDL��r���%]M��<�
>�ȝ�z�����@t���c�&���W��#W�p���nq��Vʥ�C��x�[Q>�{�l��wo+���:o���N��m6r�]wR�D.���N��鵔�U���>z�`��͈=��Y���?f:Ol�`IH�J."�S4V���ۊ��{rfn�����*���K�R��$�8j��3N�]�t�\�ޥ���&�ޫ���3���|&U�V�nW��q�t�+�OW�%�S$�ܡ��U�ՙ*2Ϗnfc�[Ω�כZ��Y�)C�긇{6ǚ�Yi�L鏪G�u���O@5?j{�<�;�%�c���^ԳJ���.��!v�o#_f	Ly[F��U&_�/M���ҿ1ܽ��Mۄ��m�n�*������z}I_��3�X�ˇ�������t&>�^���qZ�h<R���y2�9��|�ٮ�1^�6Z蕇�x�-s��i���o>1Ӈs;G��>�Y&�:fz�� rޖ!���V�Ô=B��;��';�3^	yR�֗�IP�][2ǁ�i�*D���#��]姟�zz���r�[s�k�i3S�wi^�R���lF��G)Yt��b�OzeTj`�7JNǧ~���|/+0dn}0���Z��Cj�{
y�B�%�EP����Ь֧1n�n�K�N�,N��dL��E�[g��Ν�4/a��{KwN��9�<�-�x��,�d�r�c@�hnW�t��:�.c;l��t�Ը4�ћV�@���r��X�Ar4΀@�θܫ�u���ba��M�+,L��z�]t�k7*�"/l����h��ݧ���}dPTq�E���N��-h��Ҝ�,�S�Xnf�]��������7�dZf:K��(�ak+��mݍ�/I�+��z����xj⊕��ө;�Ϛ�z�{\U�׎�y��i�3�q:6_l��gk���w7qm��ʺX�ƺ�uz����>��o;�b���%A����u��:��[Yg�psk�C���ȴ&��l���9G$9f¬�[�k���8$PCM��J:M�ݴ%�;ye���.աҰ��R�vT��^17'�c5� 5��p4�pe�M���Gm@�m�sH�����$R������H*>����]7_g&)v�XA���
�R�ZfԢp(�lLG3���j	� j#+z�1o7S��b�ŭ�C�Ӡz��
�&#]Puոr�_$6���\��t�U�qw�Mʶ�@��V����0"�cy�S-Ke'U��"�Y�	����
���w'ٸՠ
@oZ�����(�����{Y��[ywO��v__`Y+:�ݢP���23E:���:�� �I��;�x�ɂ���]@8'5GZ��>�$��t��NT�r��(sᔷQ�?l5Ī���2-��5��A�S;�ѕ��h^f�)>L��hu�+����GK+gc0���[M����L��9�m�gIQ�� oCx�k{pR��K���TN����F�<4%j�r5�/f+���Ֆ�71v�ok��3л�\����u`Ȫ�(f�qW����ea}��u��T�@������t,^�onT�=�9���Nɴ�i�<�e5�P���eG�[ۯ���}O�O߳mtGg0V��,3uիZ�.ѫ��}����\�+m�v��*�sZ7B���@�`�E�_8"5؂�͎����+dk�OR�z;)���x���H��G��mӹ����\z��A�"T�{�5���[26�mK9e�B�����2��%�6�(욙G&���֬����V�W\������{oq����ƞ��He��G_���f�z6đ捡)EÆ��5]�5W7:-S� Ly��ʶ�h��cv����eM5�z�R�|,�&�w��n�b��(2�b*M|��,�ϸ�n-S�VK�Gi{��yA��*57(X��j�NK&eٜ��K;C8'h�Z^�uv�o�i�;:NH#���Ӭ�Ht[�Oiv�7w�I�S�u�º�q��)$/O$;F�y���*y���[$��?|� �JC�,b,b�Tm-�cDX�*�������Q��TD��-�TDU��[6�TQ�iQm�V�#H�E��-�*�����Z�[*���1�TF6��d�Z�E�TcQe��*"�m����Um����+Qj��b�,�E�e�S�*",F��A�QE�Ȣ��-�Jʂ�aW-��Q-��Zڪ��Z���T���+m��-b.5E��ZR�$�4���m�[QZё�EjY�UX��*���1QՆ&AX��"���q���AE��Q*�-�n8��ڪ�h�iV*[E-+*QAEm��YV�kR�ZUV�m*�H�Z��UQ�
Q��R�V�b�Q�E+)Z�lբ�T��KaR�*R�E�TA���6)[��F��hԡmkQUb1(�JPV�(�6��b�Dm�iZ����-�EX,R��#
���>��$� ������!��t��� �}RP8���2���5�p��.�J3ء���ɣ���,��3��-��/9�yޛ�:���]�kj�+@'�L ��yrC����*�M�E	��5�<����N�����'d��%iڒd��ᮬ*�t�6S0�A.��Z��b��(�w!W��9���ۛ5>zo�x�#��w(+Q!ȴ����va$����묦e�r�|I�>�y��z��Ao%8v�ͧ�iBK���RϾ�Pw�����E�t�~3%�ݳ��V���N�Y����f�|}��+�w�ih7�L�v(;�I���r'B{�W���þG���Wb�C��'�����H�p�h��8)�'�^���-ؓ�I�a��SS�Fn���I��4Tċ7��"=��ȴs�G���\��0�����g�a�;y������N�8�r��E�8="���}Mp�#�zS�^,�Q��ڀy-
�Rvv%�_B���=\���%U:�]��N�c��
�zRP\�p�pr����!�q����B�Q�2��T^���m3K�x�x6'�K��<S
�����u�S�a��fm*;���w�H��|�[٫%�6������������z6��A�ܱ1(D���6������#-j�P�c&Q@`p��x	�6�|�*�n�8�U�%-ݤJԻ����Gv�e���>��X��Q�hNL$�[=�y��tjW��K�i�Z,u���G����h�n5��~�8��ݒ�p����ySg�>���THj�հo�+�c}l�
s���eD+�ؐ���f�Cn�����>��j4g�M[H� y\+LU�y	O�r�[���y8ʧ,/�g�ɸ�0mֽ��Ǯ�K�}���S�Y���F�G�=�|A�,�:/�x�V��76x�F�˶
90��wy��u{o�-{TT������aٮ6��F�G�e$�zllRk_p,��XU�2�>�v�z�r��-�y�g+�P�$�Cmݠkz�b�\\^��	��\�n��խp����cǍ_-�r�����ӵ���8��d�
���Á�������D�	����xv�doqOuk7,^�Ϧ�&-�(y��3i��P�U;^^&Y��h�j뽱����oT�g���
��9fB��]�{%��,���t�Oz�U��P�"d>���|�~�����ǫ$Po��� :����_�Ř_���C盧
^��-A\b��i�3�𝓊�˺�F�͖���X��2N#�ek7fv^�v�0(���OwTv�u���4�-�|»WQ�=e�]y�D���6� O3w�$`�r��Lq�v�'�[[�B,]��i�ŋ(�X�hQb��%h�s�_>b�_m^!�g\��1��k�x;�C���;s�f<4�?v�}{�S�u� X7ʜ���~�)5�����RC�ߐ�g�\�x9�� ��2��`~��N�l�V�*ac��޽Y����p�0)��?rE�Ӫ߃�֙�ޗ�xs�¹�8V5�g)���Y�	�C)1W�t�s��?x�	��^W��n/^�wb���mL��@d�~ S�z=�o��u�vH"����D���-�Gw	��ONA}�Պ�!_WW��Hj��Y��r��K\h��c�X�Y�M��Hr؛g/p���ԥ�	�'���V_���S{B��k��v��x��%��^b�n�O��~� �K9��U��u���(q6��/ ����P`��Qj&j+�u�L��>j�6C��+L\�����#2��Z><N�Z=>{�bӖ�3����h����۲Lh��ƌ\�B�懦���o��U%�CamC��fgt2�z{��2r���Ii�ݬ��HM/KJ�uV1�.���ʥ8,�¬tP�����N�����p�*�UZ���*�W׌��e������Y��{�SE�Qk%�u�O��<n-�{iaۻ+0��m���؋)+������4�9���$���7�j����	�!X�O�l*�
��WL^��b����[��_)���t�#�Ѽ�]]��|�b�
�]��o��r�3rP��� ����sy������{��tW��<�
�J׌=>�FmR�"�����
.�x�c������kϔ��Xr=���՚�{.�^��*���ʓr?Q0�4Mr$�F��B�Ec�������{��a�y;�,�<�.���҇;��˕Ց�2��	d��_jTG�+��)_o�%]�����G��bS��H�D9�i9u��a��.��$ܖi�W/�ZR��u5m��.�Ц��w��酕K�2�ϙ�*�:�0��߮��e��N�l]3J�%o�=��H7ڶ���ϴ�K>�N&7��VOV>t#D��'G(s���oe,<��,�ݦ� ��:G!��ys�7#��y_���T���x��+O����l�N��{��;��X:��W*/���!v�'y���W�3�G�U3�� ��b6������Frq��<�o\�)[�aXN"���J��ˇ���"q���<�y���T��[��Cj�)�ޫ���#r�C(���n�S��Wn��3+��
�r�Q�C�V-���[�~�k͓���f�윀��g3m� O��fպ�b����j\AkzS{]�΍@� f���b9���7���-�o��t�{�0G�;��C��u.g�/d0W����'���{e���v�{;y�o-�&
揾�bo%3<9~��B��U�������"��䂧�CR��/w=��c��I`����^p�	��r�����3�v�}W_Er�q�>�p�:�w5��C�C��GRwJ������2Ұ1��n�&zPևI��d{ی{�M��j���ecS��G��G��PKHv��ǔHb��'K�S���	��d��u�HMO���S8��Eװ�W�騰�T���G�BA=�i����X/�����p�+�]R�3�q�GB�(+Q!ȧ�� jȫ�f�]���`�7L�ǧ��}SO��e�_x�p-3N�FX��h8mIqt��r!a�kPn�i9���;;��{ۉ������)�x���k̪l�*��Oa�u��X��eа�Xs��m�.�B�ķ�ɅoRA��,��w�Xά��t��5#���EV�.�
ᕧ��ם������+IS��i����}�f�����L,�
Nђ����<�ǚS[ �;v��Y����^�n��jUҏ��C��c��p�6��k��Ոg*����*�h1���`.ע�X������0V+�%g��>�:'S�Vͼs�:����h]@���1N���!5�P��n�^腜~R��73��S��5����,{]�b���L��XB��k�^����>��:��<o9w�Ō+{O"���%�Ntu�щI:7�|<�g��`y1�AL !=tW�fU���h��o=��:�쮀)�PW�T:Ac`�%�����zo}�QxZ�g�ʨ��ʧSh��u5���5%���\����X���dg��#�69���Gj�Y����Z�vy�Vpm����\<�������)/��/��8J��Qn%Ht��B��{���6߲��Tב˪{|rW�oB���YhXR�������zj�7��[��V�;f�Ec�ظ�~b��C�V��g�+֏MC=UFX�CH��0>�	�j���:x�V�Ϲ��m�mASe�v]�!}:�w��!�yGE��x��xϒU�X��dR�56��i���TG�8���uV1�;(S3����"����"�<\V>ex5B�=��=���+�(w�Y�t����G<�.���y^�ѣTP��Y28��ac�[}��`�Z�4�fR��oUv���D�7�G;��jR�c���f�D�^3*n���P��Ռup�D�M`�B1e��*AW-RH>����a}u����s1�8�έ�9*_a�k&��gԜ���ɚ"3�5�_+�6h{���\̭���RK��KL	��L��Ҟ�p�kl�x��^�«ճb]KD�ʵ���2�N�W1ìL9���hB��].k��ۮ��,�:=,�3�zbC�f�>��;��e�/���\�����5%�{>�d���$.�ZR=�����ȲJMy}�кB�f�1�k��Z�<�Ow��Wp��L���v��ه�<4�J�q��l�o��������-�ɰ^>~��	L�пb��L����`�����,S�"�}F�|5�'MgN{��H&�Tν���u��n�P�S��^�W�	���xj$_ Qtf.�c�����гN��ǜ|�|Gj�}���P���)��V$;�HSy���˱Ө���jP�iW!�)B��u�w�L�l��8��:���Q��E�Uy40UX�ܺt���E�ܬ˘<Q��j���K�]]C�M���|��Zsyx��ԁ����T�X����k4b��J��W&�4��G�*Y}���剕�}�U:�Z�Y�z���WD��o��5i+�]M���-����nNx�2͹�M@���֑BM�<S�l^�:�;:�{YB�U���7��]�\y��(�����Mw��.ʇݦ����ڨI����C���c�z�#���uq�2;���\>]-�ؙ��25Q�a�s�Y�/�+���%����)���_��`�\+�d���N�\w�=6'/|o���T�%	'w3zC�v
ɾ�ً�d����}J�y!4���J&���ϝ׏��kL����l��+Wm'7<{9H .�US'Uk.]�<��9H[�<j+�H���g)���ҵhC��b���,�dVM�@����[� �Eg�,y������>R��1�K;W#��Ɍ癌@��9{&[>�d�`O'�$�#Om�(tV=�Xx���Ob�k�
���}F{���w�� 3�����0���x�
�4�II��ڗ�㶰#��]���^Q�d���#{J�,�:éY� �������v�5n��$�Y/�-ѷ�*��=�/�2*}R�k9v�(���.�����˶��H�l3�/�u�T�ϻ$��6<lJ̼"e
�yI]��9�7"��V���P�U�_m�5R��%�ȲW�O9��zT����7*���]tHV���N��.yA����D�;&���!wO*Tp���X��@��:���H�{�`��H:�yv�i�n�*������X�n���!{�]�*���f���#T�M��E}�M���t����:D]~����ḡ�M7YC���k�/Q����1������.v�����P�*�	Hx+����u0�B�HJ��L��c�%����RC�_�w��o �s�f����R�Gǉ���%���h�F�A�s4s���gen�ڴ�nÉ9v3D�Y����[��l�s�,WD��7Y�dW���=��S�N)Q�	���AM��v!&�JfxS��0�oVD���^�3�����E�
X�F�g�S�C����a�.�L�Xb��p���.BV���NBy���\g˽@��G�7jX�Ǳ<=���^B�Xh3����*6�;��J�nl�2�,k@N�+>v�K��~Y椆�R�=�K�x�A@i-!�H��.Ů��W�31|�rR,�X�̥�u!>q��|�]�Y�������ĳD�:Q(CH*���X�o�!��7����/M8�%�����'�FM�P�g�8�^�}l|�Hǰ�{ղb��/�Ь��v��y��cq=b� Op�a��g�q���pi\��˝�2�������Q���ua������:�E[:����i&�w;��yƼUz��#��$g�K���r)�f�� hs���cA��+j���~*%�~�Z���o�u�b���&e��8sJ��"�}Â!a�Xj��e����=��Y�B�#I:`Ɩ�׮��rGZ��*z�x"�gb�:d��,N�׫1��������tYK�=YTK3���׼C�����o���!�׊|@�����g��5�f�Xά�j�;wA�*� ��,��됌	����7ґi�{��
qvL��·�h��`Ϲ�z���mY�(j6�_؇�z|��*������!����ySec�:�u������j i��hm'<Ϣ�gWT8to��E�ςV}<3�Uf�|=L�;"Wս3z[O�|d����.̨)K��Z�d�)�TGi�n\>�����oc�M��S}�Y�Լ�u���%\z=�.�:�����wC�#�|���_J��kwu��IT�,�K�:�(�j���S�ZE�=CM��^)���p�<��V�U���Y���f��a�ٗsS�=�����g*[Mj�0Ud�1�7�-
j&f�s�c6V�t�G����N���`Z���h����:�īLJY�oj_i�,28
{ěIw�zZ����o�{ө4���k�+ ��+e^9�&���˛�VNu^i,�_V`U;q� \�G�.��/%i�K�*�&��׷�D�3�Lu�*�X��;�Id�$��y3A�CfD(os�w���lsOM����'aSg�޹�"�����'���u<�Oumo7��e=`��4��]�cf%��xSH��}�����il��Ŵ	Tbٹ�${����	��.���� ��&���ް�+Ǐ���0��;Rq]Ի�i�!x��p������k&l����F�޽z��۬�G5�;�k�H�O��q@@�yN�z�(�S0ݷ�r�A�%���f*\���^�S�Mr��\�s89�y�"��3rI�\A���6̵��a�!�q��Nt�XB�fE8[}�g�7D�%�M�8�L��H�9�`�ueA7��E�(��u,�En䄢���]f�w���b�r�����[�{C��q�
IFu��'Q���F�<̤��jL${����',��\鈵�Z���F��z�1Ł���.���ڇn�H]V��(��O[��*��g��<�FO5^��G�sV�48v���LW[�S��u����ԡƁ�\8�� �sA�\@�+"��Mu�6�D|3Ur�4��%�%��"��B�tբ��]��(+�KgsD���;JnQ�D֑d}����ot.��c:w8��q���"��|�I}2���%��E��&���r�6�WAo8R�x��6;VoZ[���z��ø��un�e\�
է݅�.f>���-	�ymWKw)U�s��>�Z�K�B�Q�;uy���V&�V�����En�VNb�$����M7{f�P�]�pj��x)֮z޵�#��VS�r�&�! y�ut�1,�
�^wa�X��������U5Z���K�:�Qn�6k ٵ۸$Y����7kme>�@uBuG�_�ʾ�G��N�+QMST��8j�ќ�]���zC��fo��1 7{w��rQ�B��X�'i�o%�����PԪ�x�Q�C�z�����c�mnWb�U�ws$�P�7)��;N^��|�r�oq;J�{N�gl��'Ci-z��{F_W�7�bb�$\�y���,�Y�iXV]f��
z�����%�dPc����
�X]^v:���;��v���h�i�	�4�:��5�(�]���h&���̬�$�H݅R\Mq��]s�4��l�;�L�1�ZMo��	�#���:�S�|n���d�B�)w5\K�NLn����[t��1�,v�(!�����{�B���ns9qu�|�F��W��jsOR:�Rp��Vϵ�Q�+h��VV6�h�Mڊ�,\Z�"[DT�����TA��Ub�FѢ�iDH�QX���ikj�,�kAEEE�U�����*��jUJ�Z�-J���`�5�"�*�����U�J�h�1j-Y���\�-kJ��Z�e��"��¢�����R�����(�U�F�[
�K����%#YeJ�q�������F,DV�-h��[[lV&[����VcQX�E�"1��1�L�+�\�( �+Aa�kS%jJ��+*�
��P�EV��E����̲��V�f��Ir�ER�`������	��2�*�2��ܲ�ZZұc��,Ĩ�S%B�bҶ�W),U�,e2�Dʉ[k�[F�*���Vas*"��(�.d*�[j̈�Q#r�km���`��b�U����V��m�#�fb�ƅ9q3,�pb�k�TX�01��*X�U�q.-�Z"�-Z��b�)��� ��jZ�9�,c�T�I�S�e,X���Tk�.T��#����2��3)��$��?!]wOF���f�&Sm�\^h����y�iV�to��ޫk��HW}�j�6�MR���w�t:�|�\���&.��y��6΋��#���W��m�U��B�=����\�}a�ԛ�/d=��D����2%����
�b�yo\8t\����E����fǨb���0�w��^���c�ۑ��n�/@ݓ�˛N,�\МP��'�4��6��F�\dI!/�r���qvZ����ָ��u��[:������b'����x�9{���hk�G�oR,l/�e���Z�	&�̘g���0X;Oؕ"�4B-c��
p�`S���y����_+�(��A��.�@�xEN,��\���u3�1l�C̘r�����.^��lK�8k��bcNupɬM>���`�ChBƢV,�<�ۮ]r�B�,�3��ޘ������ye�|�u1��13�|�P��Y"��H]Դ���E/�]�k۷"�&s>u�=�s��1�y'��y���U��Q歡�j���}*�'��>��@�H��u�\�a�3�G���v�I��h����t�����t/�1^QkZ��]�����H�Z���d?l�Y͙`4o;C�N��]p�t0!ӈ��e�\$K�ך����*�0K��WV��m��N�u��S�����f��.���؋�M��Z�|�R�߶�eȦ��{4TU��tWϱݜ/U+Ш5Wux���N�2w"�ob+�+�7��3�e+�j���~�*hgzQ8࠹��c��jY�r�P�%A5�Ea�d~���bO��m�Zn��$.�v&k~�S誳]ʡO��{�߇9cܦ}�*^.���Y��鮻�FB�y�z`ь�K��=W�������NH1Z�����xuܧ�r��+��fD8O�c�^�:�
�u2��h�@wj^	�Ϻ8�cv�'[k�z���p��~���^����3�| Y�TkK{�3�KYz�C�����-4�'R�;�a�:*��M�
Ƙt����I`|B��(m��;=���q���o�Jd�4L�vJ1_�:��u�|�؜��t�aL���,�S}��.�͍�"�E�%X���^�DT5R);]f�ɿK
�{D4/���!�S��KZIԘ$�N
�.�-�YNT��e�3d��6��(A��z�e�s��Ҟ��W��	BZ��F�RQ�4�Q:m��u�7���}s�y�{Җ��0uJ�}�!���xLٕ�{Z�R}��Q��4(���)��j�Q���j�]z�S�"n�Vj8��o	�ڏH��j��:��j�Ֆt�ٷ�J�\�`!�[{��q��V��y�{�!�=�	ub��:��Vv1���Rn\�{��`�cs4�Nr��T��2J�O>�/��OD�z� ��Q�:��sm���W�*G��;��.M7���烘�bT/�Zޕ��xT7<iieWړ��<=��'Vs���9��T�ZWT�酕�:��8�U�U�����s������z�H]�c'p���2��ٱK�؍���z�^;ҩ&af|���Q#������;8$�L�g5�� yh�c��8��f[�	�.�_�0��}��u������k����g��2D�������+���ä5�_�e�P�P����%3��_Z�c�Ay����<:s������B �{	���u�e�~i_�Wn��B��	[;�+ݝ�)�v���y9H�ŧ�5��P��5�d�/��n�&�'ǉ�/R��4�Ns{�!�֥�km�b����t _{08W��C���N����<��<����73:X�j�;�M?�^+�ǽo���
q}��$�L��Xp�oT#�O]{��%4�[��A�˜A���&�k�x�޼���Z�i��ɰ ����e�.�n/��]Cʼ�[��w��n�ң����[�ռ�+�Ma\h��l`�t(.v2�rAL����E��ѕh�S�p��(�c�λ���]d���л�r"
��nK�b�'e���u���>���%s^���;����z-�G?��Z>�v�U���!��2sX�SޙUS+�.��>�m���OF" �'���0��}3u`(	:C$��}=�~��f�Dv=龻��)~�oӮf�z��yĈ�4.��we`��~֏E�t� �|�zӭ����c�P�-�����_(D;��� ����4G��j:��
���^u��<҉?G��m&��Qt�⋷)�"��`h�t��.V��śJ�9�	.".�K>�!a��W]v{�6��*��<�q+�P˪��:��{����EꞸ\5L�A���9��������{݄ EA��Bq\p'\e�]�V3�9s�'��m#,"��1*��Ykr{ݚ����i��\�U�!�dq�%��LV)3�T�_�o�.k��"�n�(�F�o��ohR�zh��0n�Ի	�j��XB�ke��^���l���r� �P�y�-�ۂ�����hc���X��r ��Ʀ�;Rؚ����^��u��,�n%�س{�5y�t��i�N���Tu�W�����h�Ef���.G;��t"��]�-4J�zNVls����� B뭎��{K�rZ�LO�_"�s��q:@B�׊����ɏ�P���K{�,
Ѿ���W��
��|�T�]�PW�T=�C\L����z�M�Vyn\+�+�C6�j��S���-�E{	
�ܼU<Y�R���iY�!���	�fP�GDls;�ك�.�;�탹�q��F��0�1+��KH�ł��h�X8x���o��B�J�n^����v��*tr��!'}Υ���ً��2<�Ex�m�tyV+O(�.�Cn��)���WƵ����g �y8K�r��-��Z<mi�bH̥CH��,+Re]��B��{����,�}؇�_0<�MN,�UsCӍ�v4�+O��6
�"À��y��ЧS�����PuݑWR����MX6Q6�� ��nAa�bY����ņV�U��ɹ]G�++x�����kJ�v!��_�8z�)8����¦�{����EGG&9��Z�npx}�E�R}��Cau2�(S3n2b2P�;r�r�҅«��Yٽk�Iӌ���ʻ\���^]sy�BW�V���f��N���TF�i�7u�lWv9�U�{�vG�b+�z�G���z�]Z����b�z��GP�S�GMX�g�S��N��ױm274@��GR�lV�ڳ�n��O�Z�u"����g"�;��u^���tH~��W*�B�и�7�q.�]r�B������`l�yH��T���9����<6}lZp5�>����+�D��u-*�.�_��f��r!�K��9u�t�8[�AX������FEq�+�|�xxJ�o���F��mU)kۍ�T��{�y��^��˳��6��$=�'>r��b�4��^�fJh�fn��MeL�5���{�GR��.��p߳;�^��֡���ɽpXV�Õ�jX9N[ɷc*��������c����YG{A��"��.�B��"gGg_�<��>�&��$�y�G+�nO�>Pzw^e@�j���j�-�"��$�φ�g�U�~��w�,ge����r��9�Fr�{~���"�j��bn̈p�Լ^ufǪ�"���)�#sr�}��2*^|sU�������-,��15�#s������Ա��n�#���{�[�#�c�bwL�y2R=1���)���]�F�¬ح�Q8*��V�����Z��.ǋEê���h�&�R��&Z�/�n����+��$��V�_^�Fl�˵]�t;�6F&n��ʲ�Ȝ�� �hLp���#����9q��2sY��-Aeg�.�:1�}���"��o=+�4kU�F�l����3X�RK�~��9x �rB�#'P����br��:�
�n�a��G�z����{A䶅��k�J�}o$&��&���uS���(s^"�6�p>�{"��DsY�c�Cl*#	<��-j%��e�+>�����p�϶O	;rb�o�%�pr���OT����"�P�fa4û"��^��X'�b�Ŏ�WS� �����Vl�o(���nͷ�;��0�ǘ0OK|��e��	�L6'�C�$�4��:��n�W^���i|�Jy��B=3���	.#�.W�`2���X��&��ƪ�'�C��ޞ��?�2��jB�=xYK�:��8�U�6��z��;G_:^,Z
쵫.M?@��JL�s��"����Yޥ�7��V�0�r��$x��1���k�봦)<ݓ��2,��VjW��Ƀ|��u`b��{L��tˣ��UW�)��^�ؓ����f���L�Ǐ��^�p�}��1�7�n(F-����������������Y�;~lv��a9S�@gof\�ݶ��'vX���[xvΉC�\�YP	�'S�e�G&`���Ê�=O�v��W��U9���;��+�Μ��x��k���t�-�.rY�+N� y�n�εf(U��q�{�������w�ЉC��5xR�v��}�-��f�+u�k[�xE�;��s֫�#������F��c~���UH�5�d�V��!R�L :��xx�����[�k62r�z{�i3�3q���1^��@ǳ�9v3@�J��p�-ͱ�^!���p��C^�����g�y-�\�-���
�v�$�&bj�3��(C;��05!׹:].ޡ��j+i�9I�K��7�8��R%K�[��N\p���뇪}7=JWF!�?��A!�jZ��W�rJ�u'b���zFǓ-+�*�]���.z���i�R�9�C+A����V�_Ef�]��M@I�$s]������S��N���GǕ�P:U@n\j�<3����Դl�������P�Ûq	���p����;Qu'�X�a�Y���{�uK���E5V�Y3��b4���v,��E�$���hu�]9�{s%y�m*nZ�Х�E҆a��P���X8w�7��l��YXV9Fӎ����j��ج�����LR�̬�/ѫROݝA_ю}Q%ZFM��ex���N֞�!�hs[X#�Q�t�#��X��z8qk�n��XKk�b6��.Z��qg,c]�!������W��A�v��E�ȵ.�:��=;ցƑ�`�P��������h�BD�R鞂+�v�]k苊�����Q�M�E����D���$[u|K�r��x�3p��z)y��T�Ư�M�GgwEV�7^�o!�C��ƈg�Q��A؂��L�_\�c�b���g$�k�U��ԧz��t=�
On5g�2�Â�����(��Gƻ�Y��Þhhbv$=x���.\���{���"{�%80��T������(ASMw��%����9�u����gZ����}~�6ϺV��X�c�ixd�k�ϦV�Q<�4Z�k��c��P=�S\u!���eҋ�]�ش�G���"8;צITFh�q�8U�pg��z}V�/��we�Px�_ݛ�
���W�z�`.���/$(o�P�gGx����)�L૴am�M�ȴ��A��c��~���Z�R�禮/R�B�t9_ե�*�K���J�L�ݷ�c�W���j �q�s�8K� ��O`��{��G�ҡ���})Z+��J���:~������w�֛W��LD|'f��
v1����0�t��R��������ΎV�1.4E����J6WU���E;I��is�Y�����E�mj��(wQA 0���[�(�Y��v��Ǔ��*�|^���z��R��`/k
t����~���5����e�0���V38�v%�k�m�ޓ���huG�'Xlz�WK\�7r����Z�����%��z6)X�A��bȉb�o���c^��,2.Y��<�n_jp�74�g��0�&�&��z�+���;ZU��� Z�=z���;�/��+������lR�=	�I>۴M(��_�)��M)�d�F��2��}N{H�������]gOt�<����y.���4P�t�B�j%b�5ޡL��=�)tY��!z���&N�o_甉��y��j�����b�%�,�l�t����N�u�=Z:ݙ{����Eħ���j��y�ht]�Y����1�����
�p��6c�H��]�t�onmz�����ɛ�H�\�x�LS����ܯVE�*9�"��K��4��;�U-2t���PL��)V�P��f��:�Z�zU%�\�a�nV5�f5;v��5��7�{�J�mO�f:_{l���lo��]��^S�[qxο4y3���j}�]��G�A-A:0R�9A_Q&��}��,��un���d���Y;�n��q�u��p:�Ϗs^!>*}���_t�f�ҷ��U�m'����\;q���'���˰[I�����yl���%h"�C-vQ�[4sTT&�sOww���v-��R��X�PE�����:���z!N���^a	u�ޥ�8.�&������rD-ϰH�<��
��32�އ;�D�,��5"Ik|�
ҏ�B�k�b|�t�˷U���d��ZQ��QY[��Q�Èp��Щ��Y�t/t�����v��y�a��[X�Tfs��%�w�3�u_V�-�ug��	8X;AJ��{�n|��`�e��m5}2�u���Q���ѡ�.�D]�j��!h�!ۧ3j�^���k���1�pYь:��e;��c�H𳦻4$�����O�Ķ��
P/@ܼ�R�f���ʱ}�t7�f|����(��F�'e�	���ъ?�n�u��g p򾹊���#Ը<�o.�k�R��9��ݔ�a�(Ⱦi͇]�wŜs�*�"h%�Ulg�ƪ�+��k6.}�9DGQ�
��9�.%��l0ڼ	��z��{���S4gڱ��;k.��C3&��^P�-��r$��ٷYwp��<1�V�C�;�\�����J���O����+�$6Z��n��y�a*��v����m�V��p+�3��\�Z�gQ���l����kIl����Pʧ7)bu��lk{҉�
�a���W:�m�-\f^��,�始�. ��G����u|x�����Tv�e��K�F�i{IrՆ%i;�.�g�1"���姗chݦ�U�Kvh�z�Yj5D�m�)�Ϋ�[�T��q£w�Ƭ޹L�F�+��y�w\�Jև*��|�A�5���k0�6�vP\��Z�ɕ�;�UI�:m���Kj�`���HTWqG�TR���mB;)�/��x7���I��r����MQ���%^�JN� ���F�$p�ƶm,֑͢�=o��ߕ`��y��E`�z�h�H�H:ջ��O�l��y>�����a;�ivodk>�knI)�t�@7-�S�(�SY����(���|�vև8�-\�3�Z�u4��f>��:X�\��o���V�E+�١��������gM�S�˗��goJ�ݓ)���^�&�T�
ږ����ב��G����M�
�f�]�)@�8�=�Q�C����(D�c�q	�P[��t���(].x�%L����ՙ�t<'Bv���M��dǳl�ۯ%^�� ��4|$��Ő֗�]�ެi>��Q��PQ�l�Y�{�VH%�̩N^c蹚`�t�+��$R�U�Emb�+�{w("��_J���u�V;EL��2���wW>�3��e�=�+��W�c�S�5.؟k0�4.�{�ye���Ը�Kmw'���"W%;�fWU���Q-̨��Q��jfP�2���-�R�1*
�c��r��j�X��fb�B��\2Z�q�7,p�
�ܶٙ�B�#m�,r�UV1��hc��"��Z��8�"���m�U��LkZ0ˎ
[fDEƩX���0U#YD\��B�Z8�q���[L���11�Sb�TEph5�*+��.7-�-�1��J�SV�-�+�(����E�&4D\eť0�S��hŭ���TK��eZ��R�����kGU[a����j�"�f[-�T��,�QA[LLH��"��*��[be��QF-�1s!�3˖�����2�Q��ڌ��S�i�f%��j��Z�e+E"�*V��m"�\l(�1(�q(��VَUj���ت6��Ym�r0s,1�)mŶ
%lJذS2���k(,DYZ*�*�)Z!K*"��b��*,dU-ƬET�E��h�Ɉ��*�m
(�T�=9�f��y{�A�+��cԷ^U���$L�լ.� c�;���|6��꾴�Pm���L�X���}YpF�b�:����gt`
���f��m��ڑp�ڼ�6�5�;jC��*.]{�^h��u2d�/�����Z���~�ym6x+z�9}f����|�}��e�v�	���]ᗝ��A�N�ǆ�ىԵ�~j��]�Yn;'X^�c�%��/g����A��s�S唉�4`���.��p��sއ>��]�J�k��a��VnWԁ���t2�{=Ӓ�����Ī],��	7��!Y�I��`k�ri{�i{k�J}��mB:}v)�2}yMY���(�b��$v'�}�������Ur�����i�!������TF�	rLv)����zߕ�
r�S.��N�T�ji�򲜙U�1��+3�ߏ�����Y�`0���1H��>�c�|-Wau퍼��Om螾�)w[�\���f��ieE/�M_V5uN�Uu\�$���{tf�H��B�s�{���ブ���[�b��c4�%�{7钲�!r���.Қ��V\�=�v
��1\2�;ܥN�����B�Q8�h�:��r�'���,�S{�^��0�l|���v �|�6�	Ж�N'�I�GB�6�����Lh�ـ^5�p �7����(^'Y@��FYF.^$Z���GV^Pq��F6�̲9���;�[�V�K�T#�_�q�{��z<��a�B�Aʻ
��Zp�B|�[l��gg{������i%C#1xT�"�V�#�lS].V_�ze���R��������k�g�~��z�ET �����"��L���e���.�
�>g�|�9�ޫ]Ҧ<w4�?q5�m�d�0����Z�����Q\��QO+x�B^k�6߅�y��]��[����%��{�^��n�%Vط��+�	�=��*7��3�̐�)��QB���]oS���2���}�-��0��@u����[˝
#������у@U�ϖ<t���AZ<�Ёf
��/%�=��t��u���R�nn�!�(�}��]��ū���K�"}W͘I�L����	��Q��u�t���ϪE��\��1����9](��"��gp�s:�+U��nK�b�'e��mzv���|'s�岥A9c�}^f��=P�\�҃?jM�T6{���7X��J]��q��\��ks^���'���;Yy����YP��k�O�ǯlm��5��nފdQ{��{���t�ק\q�/�ou�α,U��OXk!��������Z�R��9�S����
%m�m�ӝSps��'�oe�-���EtN��]��3=�w�K��cZ��o�Fi���G��v��@p%�;H�h�*m�^S�D���iD����%N��2S�J+�ʐ&y�=h�f��9҈μ#ƺ�pɉfX����5���S�A
�.ȅ̚a���}OH籭GB�(+C"�j�ӻ	��9�{Z�������UC"�ȭ���ST�u�={J���t)qt����y��Vu����ff�4,<k�	�N�w)�̇�:����=�ț^���K��ӷ��p�c^j���{�2��0X��i}���-s����^��\7�擮xM ��4�RiM�]z|b2��Ɖ�pS�Hg�"��&��v+��9[7�}|~o��Q9�(�����n�^腜~Q��*ab����x��|XC���!�x��cY=\k��nl޼w���j-�[�;h��8���=�`���-�M���9Zs}2������z�@��3�2Za^߭������+~�~���<���_l�g��b�5[ws���Tf䜠h�v���н�Cy�cU�KL�G���zlk|�̍V>|��k÷��ٽ�A��>�:�p0�]�����}��C���Rgk~�'\��������H=WF�ŪA%M��%��\|��<7ky
�yN�e�皝�U:}�˺��w�\��V�Z��vӥ�ǭ7�>���֏x���������]�m�PY*��Q����aB6�|}�;V�r�_id�*�P���l]\�8*,.$����������o�*w�w �a���wV�m3��p��/
[h�,���CH���
��ӛ0{z�;��X�2׆�f_��r�K��z{�ޯZ<mi�g���]��S6>�~DeAH_9/�v��>Q�����Q{�&jrq`�N��uԅ���+�ts�yc;�q5x:IҪ�.F��/UT/����]m���,�����Lc^��a���iެ�g�ݿVum�[�}��G��\dHgyݛb���x'�skA�q��~6���oy=�]N`���^Oɐ�q$8%���W%<�{�
f_e����p�kL�<�a\�6��,�[�27�>{�]㕵ؗRߦ�E
B���P�|��8,�<�[���%��ق�ڦ=�٥*�=i�=7�ڵ������5S�NE�>���K6l�t��}�7� 1P��GD)��ZQ��[��� E|s�����}2�w�gU���`�q��t�`��2ܲFxv�[�^���k1ѫ������-Y�re��k3.���܎o6pؗt���PCbֺû����M��:�#`Q�yr?�4�O{�5݉`�%\Vb��ȥ����5�·\��]"X�{c��Y��P���E����>a{�ג"��q�v�寳�+>ҼUOu�q�t�9P�����."��:pjL^���<��Z��~�52���\�x{3}��J�.���
Ö�4�y%�b�;���2�OsK&38��߄��l箊��C�;��9o�xl���5c�c�;�]����3w��ɧդ�9�ޕ�Y�oh=�>R${S��Z!+��ϼXG"�^��13+7���'�zpu���6t��?#�cud61�ȇ	�`LtJ�d�^u��]�}.�[�k������3���Ե�~j��k�F�׏��P�i�.{�$u�4�[M�/g ��2qc1p�b�aB�<�J����C:]�F��j��WSTN���6����b��vRXI-���K�U9!^�F+��� k��֐t5*�Ǜ���?A���t�z�X�[��k:�o��Q*��Bk`""��l",�g��ՠn:K:mp��x�v&l�x��0�b��T�r����֝\Nv�_&_
"�oGGW����ּS�¥�B��8V>��f���+O,i�]J�;]e����
|{v=�߬�n'[ΐ��ꋦ4ު�J�B����_��r3,lܵ(�9�9����{꩕�x�+�t����I��-�z�q~B�]��3����r~�d�z�͖߽C��5�Og3��[[Ke��VNۻ@��0I�P��,��j��"���Ͻ������..����z��ߌ��3�#�ʊ[E9��)�U+>�����H��C۵��Jَ>�S�(��!A��HpM#����B= �ZCߡ��d3�\���N�)]"�C���}��\uRį�C������/�M{�g�Rݎ�]�>r���ll�:�#��ws�����KF�4/k �d���x�R����du��p����w�R\�0����<L�<9m�oQ�\���UP�Xzp5���	.�p3O�X^Vϴ�K:�1�]��'[X-$M���K[�QS�;�ծ1�lHi�o�P�U���ä5��2���#d��;G�x��q�;�'�e&=\q�P�	czl�8���'�{�_���^��V&	�#"�;��]ޚ�Y���z�ܐ�~/y`�D��'/�Q_W�>���}������>�`S^�Ԗ�66no�2��EZ*k�Cd޶�k��V�&�R���VzI����UK��^�W{2� |��m�֪|E�q:�H���a�u��XNJ6gM�|��}�sh��Y���D�/�L�����C*���T.j|�9����˰k�ʎ���&(pߩ.�'�p�\|�/��P��n�{08P��r�9�%wSV`ו�k������ *�������GB|p�������χ����W�  ;ks��ߙ������1��v�1v��0��l೸b��u
��';�T�M����ai��V�A-ӡ��=�?_W���(Er��@�A�#�;�Cf��h���]U�����ݴm(�S/s_���cZ��|�)��%�<l��6�}�W������ɽ����t9ג��'Ք�n̄��Ҋ���An��u`� �x��_C�3/ܚ�ņh���_a}n)�{]���bF|��
�D9y�4��s_��i*���t�V*�� Y7�l?&\�z̕�w�6�r�J7�6FZ����<<��(Ϣ�W��
� |�ZW�:���� ��x��t"Bٹ�M�>x�ݎw�d¼�vv|j��|��PE�b���I
��\��u�]Vſ��A����OwVd�o]o��0��|	���D˾�i3��a��tH��χ5��Wz\���������Lx��ǕY�͗����Н�8,N�i�ҹ�۽k�eJ\�� �)�oR+*��V!M�4�g����Fa����{|H�n�-���5�^���\̺��e?EV�.���:���&�����b�9G�jף%e�U�YQ�����$��d]ozxR{q�<e��=K�P颋>�|�zAk����9|�|$��w�b˓7�[�����)q^vqG�`�W�蘥ӯ�[W�[�q�Ó�'���r����J����Zѹ[�ҩ���)S˳�������\L��_�\�7�X�g�gL�X��g���`VLk�Äן�붝R�cҭ��U����{�w�f�O�����<�����J!�'���[�ˇi��H�K~<*�i����CHp=́{��F�]��k�Lk:�[�W�t��B��wU�g:�h�a髋�R�@�9g�9hK#���6M��X(@��p��V�^a��NP�Υ��s�=�^[<��˷c�����{�Qn����䜏��í\�CH�M�
�5�tb���&g�|ȝDv��:�U95�ZW��k�W����d�^F�D��7���u��^��覬�D��k�1� eom��G���=G4�[;�N�G��)�b�~��r��͡M>������t�h��W���9v��(�ӹ�DU�LB`ԛΤ�X��b�j>c�im؜����A�	����΀clKF�p��\�۳ү/-Ҝac�j~���_>M|�#�Co�Z���� ���B�u3��X��zB�shH�������M}�/��Gq�{χeȳ��ڸ���O%���A:���1l�C̬β+i�·�܈�~]]#�V3U��5�ԴMƊ�6�_��D��5��3�ʃ�GT��گ�_�[r=M5�γ�K#���%��>j����(o��ҡ�tK8l�t����ī����N���^rL�A�%Z�8�߄�YHt�]`r�!ʻzy�x6��^��lx
ȳ�]�\gٹ;{�8�*B�G����pY�`��g�J�D,��˔/I�p�:'��bkf�g��W8p�F�J�Fϴ�O.J�~�f�ߺ�Z����+�,*i����x殄��7Y��>[uP�X~C)1[C��}j���nL�>�/C��xި�������N��6�ڬ�v�V��ci���#�@hh�v�r�גG��{�+C��rga�Y�SM�(uߏg�m٥��,�����i���c�%~2�`N����ƚ�ݝ��ה�������ZB8WP�[�n�ݔ����V�c�/G��J[{�@4�uwL�k�:X�a��1Wv�\_2 Z�.�\쏆ͺ��Ż��svfSܸ�T�O5��VK�CS����z;���6����"�W��q��Q`���gɌ�:��:��D}Z)��P�y({~ś[H<57��N[L�F��2�4�G�ܪ�\�:��رc�(0lu�P� �%+OL~=�.P󹃶��f.��'�缙ۭ~���^"�JK�Z=>}<M����4L�p(�$���ۂ��y��u`��C_��i����+د'I�
������49D����@zL�������s�{���U(��o��x�N5ܽ<hu�#M�&	>�x7��,h�f�Y�ׅv�6���'��޴��{q����|�����5�a�J��R;aݠE!�IsP�.ɽq�F�<��'��r�R&O�CΥ�C�9�V͘�������R�ETIt��sM����W9uKQ&Ϻ�X��ՂiF�'C1iD63J���^}.+,�����+]������RV���'��%µ+�)�3G]c��_u�]
��9WaW�BK�z��O7ڣ����E�#�`�-�5d���;3�墓�c��Þ>��x�3|�#�������7������R?��f�A,�{��;�|�3L�����!Φ%<.)��{����u�	e0��ɻi�q������T��{�鲦�W�v��ꙩ����ܷ�}��h�4]ͩS��7�BW>]�U�$Av-�������B��>�6�#e�ҥ�2GL����C�[�r�#�4'��7_�|q�P�R�[���f���w%Ե�װ$j]޷��fu���Rid�V��Z��,����7��rA�0�l*����d8���]��G���y�d���4C޴�S~�D����O��X�႘�5�^� ݘ�qbe�o|�d�p;Q 6+Ms���]���oC;F4h
���@��.��4:=;�J'��D�t@�y;;{8�>8�]+�dꛐ�7��ʫ@�At���%4���6��@fI��b�0�B��IvS�"�Av��f��$�ٚp��N	+w�4����%v�hqlYBf@
���9x��`��f��SVfu�*��xT���n��+��lli�u6쎹H�FX��gB��Ν���7��jԞ�P�����{���G�ɬRwh�v�N7�u�w�bV�zr��g1�5��V�fi4َ�U��R�\�xս���z~o��� ]E��b���.�빼Uj볔·k�u35���<�+I��	��aB�>d_��v��l�L�1`�7�m��L�O�i�TѲ�ݖɕ�r���^�Ê����h�r���ՙ�9��ޢ�F�^��T`�u7:��m^ ő9�Y��ޔu��_<�vkM͌��+��+�S쒅Ŋ��|[̜���^iPG��;;X���` ʻ�Dgv�wv;Ί��e6��j�oE���8�hb�6��RQ����u,Vy/�k�ï(ςc����#��_:Nɸ_|YŜh�oh�Ev�Ժu\�<��]}��Ntq�E������}�&�"~󲇄�C�Uv�w��!U���2ȃ�0n�>;��S���g[��+�	��� :��N�PaAX���Ja�=��{Q:�j��r�3ԙ�����v�|�����-���La�NۛV+�k9ғ� 2�7�ٵ�F��"������Zu"Kv�fU��b�+y�ۭK�A��Z��ݧ�u�����o��p�]�l2���ߗuiY;]5�����Efغ��u-��ec�:Ոi]��\�����G���>��[ZXJN]��-�Y�������\�U4��%�:c���J���ZU����зE|����\�-ƶ�5�֞9+Z=��/��r��
4�}xD7�e����ԓ�z�
3FV�j]9!�g� (^3X9��7�<j����u�j8��`����6������fV���l�����3��c="���܏)��u�xA,��lF�����9��v=�?<��]��S���B�]sE��WK�![[���D�2<������;5��P�UJ��������DmmUF1 ��5�aEfZ"V�cQ+*�B�ܦfd�""��6�)lX��b*	�E
��U-*$Q`���mb"�5E��6�)Db�["���U��J�b���b��--�(.fL��R�����Z%e�A�++)ԩ��LLeH�J�V(������2��J�X(�-�)kj �j�ҙh�-Z[QB�ƮP�&Z�[Ue*ܥ��P�V
�ʕ��WaY1���iƙh�*����YF(��T�-����c.f�fS+-h�VfE`�Z�%Eb��+(`��%`�2�q�-�e�,�3%AF��`e�B�.Q@�U�Leq�LJ�-��%�5b��*�X��"��-R
��-1�0��U*J��D��B�(B�q�����s�1��ܾN����C���{G��w|�j}u��G��z9�R�q[���.����	�����e'���y����wlW�wT4V34�k05ۄ�Y�4�d��Cp:�V�m֮�мY��T�1i�Y� �]�Y5���7!�I�����:C]~�L��^V=��.�߶[�y���!��/VZ�N'��4w�q�<��������>���yKt�^{^7<����ۭ�6-d/�����၏,
��k��훎��U�]���
o^H�J��Ȟ����%�dK���U����
�v7]r�fʅ������va�}M����vL�Y���%c���uQ���
�t�$��L�n�x���*���ɯ�!�2�x����V.�Y�~#����Z���W��0h_
q#B�k.[�B��w���𭴧��n�xL�{\c+91=P��z� t�� GRh��mZb2�4����8<~j��"��X�)��������C�)��`��k�OR=b]��֚���k�/8�tE���>�p��>�$1_4��e:���BF)���Wݷ�H-�_��Q~>Ҝ2��,�H�X}�o�t=.��<��í��^t���N�&��+W����)�y������e̻��>��$�՝y�Y�������^<04z��ۍ^�O7,����mm܁�u���/�{�G6�����7N���'���=��o>&}%,F��	qx6��i˘�J�ذOPy$x)r������f�J8�uEZ��ڂx�6:�C�(��3���a��˛OK�ZϪz��v���ve%��R;���,{����D] ��0�?Z��ZWN�w�.���'ﲉ�AG�B�z��^�z�����=�\Wf������E���߭$(6j��/�ku�Jy�k�pf���y=�%5��#jwYj���˨�FSB�j��
|��g(:��%�
�]�����{��泼��L�#b�L���H{�p?(�P�X�8-��2����H���H�����p�W�H��p�2�.��[��m�����q�&*R�Zy'�]
��;���ͺ��:��0?u�B���U���(*�b�%*x��P������(�yZ�����`�`z�c�e�x�>Kq�V=i�g�%}q���9֥3�����-%o���s�J&e 7��!}��>Z<�����,-*��."�&F*����g���ڋ�r�%�h�^	�dO-p�.@-|�h]9ݢ�n�3�g�.�����ԍ����s�Z}{�����­��G�^����/��tV����\j�#�W*.�ײVJ:�C�:�����g�!�5ij�Rbnwn>��`=yԶ
��.��+�w[J:ܭ�6J��D-ī��L�-�'u�L\2R����#�Կ4/�P
m�����i�E}p;`��b�Χs�9�c9d�z{/-��Z<M�z^у3���ѕ�8ͥ��8PU�,�5�C
�b�����àK�d/�[�� j�Μi��æ��:���@�:8��t�xĖ�M��GWp88Oa�� n>d�]�2Z�p������G{�Zp8,B-١��Z��ԋG�¬SkJ�x��X�kdI��ib~=�ЉC�ܳ!/���U���y`0�P�$�@��W%<�{�
f`��LAP~��_!�ɞ������P�0[��{n/R�Uz��.��MƊ�n�
ta*�3��FY���O����/i6�$���w@������Zr(o���v]�d�C�W����`F��{���X�`HM;�,�3�R%��I�E�q�+���������/}3u�0�g:=���4�Ȑ�|3�Jx�;3Vk>37Α;�yB*���8�eZ���ي�E;�F�޳�]����|��maj���]}�c����׳�[y������z��2gY�u���_�D:�v�����lГ�ה�s��ů��[���gtA������_Qӂ��i�kg[��ՙ�9fb��ٝBr��^;�M�='^R,@�W�9fJOl�j�aχ-�<�K��;5V��>��D�$�ޜ�m̹��ޡ`χ�+�L�>�8��̔�(�p����Zn�h·�u�|�c�:[][�0�/�vVu��w��
�5�i�/&:�X�2g�R0uD�
ka������Si�?�i�l���U�h���u���4����6�L���i�;�1��P��el�ܼ�y.8v��������S�� \OW���n}~�8v�lT���m�Ѭ�mE~]�n����&6RY���^'�0`\,1K�3\�����T'���ȹMV��V�ּ����gz��Ω0��,��K�>Ih�������T$��d+�Q��^��#:nL̨�׶���l=S����hSA�/��P�����S\�U��HM:�%N�e���e�4n��;���9��4K��h[�}�k��`TN�� �gȭ�sGF�;�T�n�y��>��ǖs����ܔ7~�ϔ�s9Q7������4)U�(Ɇ�lH�˫��F)�z�A�kp%�G1n�� �[�35c�l�pWM�4�u2:T*@K�n��t�<<�!X��Ǭ����s4+��,7X+�����8�P�f�,�QYs��79��K�%�gh�4�)2�6�UI�s��ؒ�4AK���-wc9,XןZ���}m��fnl�h`r=ܭf=+D�t��0�[7�K���]���a���H���D�˪�{c�b��B=��ZC���!�}�s�K���ys���pA�W����4��4�du,!����^�,���qD��Z�=
_x���� �|��wX|O���M�d�^+����o��[�v����/�2��q�Y��o%"�T��(����f�f�n]g���2`�m�Y�����&����O����6&��tU��x���h�d�����D;p��i�z��r�y���2t��۫�/�Bڃ}[�ˋJ�\��q� g�Լ:��^X�����fuk�ir�k���X=hˀ4fz��E>HJ���`�XP�0W�\�Ol�u܅]wJբ7g�}��ON2�A:`kR�c2�\��P�^�P����9��DT:�c]u�����}��S��;���b�]ګ�(l����9K�J�[�7�">�c�a&�͠�:��ˮ���v7uQ�Wx���ypX�IZ�F�R:x�{��+��^���}�%حd�Z�_V��\ژ!1��xkK$���z��7��-_H&���F�wR�t��;1w"/��T�FwM����ܺ�z:5�8����2���n�,��fη�^�;z��eZ�]�/�a�(ug ��b3���t�wn�W�z��lM�v�x�ziA���w���=�;��ֵ-C�+ֹ��+�j�`��ﳁQ
bH���uE9.u�"铃X�S�誦|�3+L��n��w������O�/*�������O�&�h���d�)ϗ4�C�S���P��sB���o~�[��oLJ
�۵p�7֏��8҈����]h?
s�V|�a�Y���0=�j9Z��'a��˞7� ��8�R��vT:��҉$�k~#}ƃ,����9�]_�*�u�M�g�{c���n���׎30���a�X���:E�b�B��]�םarv;׻�u���Ӯ�l�t�x���>=5�~�\5L�(e��(E	b������6k��n��f�٢�A�q���g�
}�����9ғ�{7���S�
���>G� �S�!��Pp�N�a����e����8Fk�[�;t�����3��L,V8-���\�+��w���Jmnݕ��i������)�@j�!���uЃ����L�
�\�����5a��\�*��աt};'�v;�K��Wj
����>�.]���mk�t+>��7-�;�x�Z��{C`��,�q������be(�w^I(�}�Y�;6��Y��]M�,�[��n�nŰ�s��C�0q+��b�g��+I�}�̦!�}���&>�L=��(��P7�S����z=W��t|��-��F�Iǆ\��Nx7�:�}��?/b� �62�&5�0�5����Mr��V��*�f�9/�u�k�1R!'&"E��w�H�����C^GD-�'���7.�xL�tu��1�Z��y��������m�19vr|:Xz��;��*bᒔdxv�{��pnVY���d�����mI�������1{�̱N�(p:�3�Nw�����C��w��{D�ڤh2�{�k�\�Ux��z��*E��aZ�V1ъ/d�0�98�ҫ�U|vVn}�j�+׮(��>������8��F�\dI.3Gz슿����Y�SVl�\^�������/���^y{��������hm�v�X=f�Ϩ�8U��gkJ�[�􊅂"7zoF�?F�Sۣ���+�w���]�/��,0�W"P�_\��.>�K�����1�]���Y�A�m,Wq<J�#CI�B��y��]A>����[rnP�ǗWR8��pI�\{���n��V��>���]%��g{�p���c<87�J�����g]$��Mn�w]HjKXz�,�螭Z� 1������ڢ�S#���-/Rm��_{Io��k3뛛]�[��*3���lK�ENаC:����t|�q�6Sz?i������x�K=�Ydt�aO{`j���C|�P�=d���zy�`���_����F�H�Jʂ�3�vh^���e��H��|�Cߢ�z�8*�Z?X${f{�y4o�c�^��,"�El-�Vf�z�^ޖ).r�Z��G4�s!u�-�|�EF��_K���d��Fxu��co��>�[��ʾu2��]F�6��i��v=�U��ov��p���`�r�����Y��%N��0�U�:g�ź�t���7�����i�je1�]��'|� �ޏ��x_�1�J�!��=▂�T�����9���Y
��W�����ά��Xd��6t�~G�&X�P��^]o�k�^c���¸5��LA`����.u��D��o�Jz(<7�����yi�\OT�P�-=��oe�r���)n� ��ax:�	��c,�^'.V.�f.Pp�Ȕ�����躞�*��-ŝ1wGgv�prE���)��r�6����%TM�ܮѨ'��h��E4E�{;n��6�ש�=Bh�������xUu��B�G�d�����KE^:Usz���X�6�A��۰	ٷ���mM�2�fu��xnWV�gc͕��jse,}��NJ�k��dm�Vn�i��>2�Z=>{��> d���\2U�"�OwxJ�}��,�?�k�Bqu����W����U��4,�S_r�V�Y�s+Z�G�<�R�1� \t*y��f�P�gںx����&+>�B�]�P���"\��n�Z����r9FK�j+�������T���X��X��vû@��nJ�&#nbx�ܤ̳C¡-Bņ��vE��Y��z�hc���h�1�[𛎔e\��q̄��fW^�X��A� ��ȁWC��,8s�oV�Ǵ�-�#�Ť9DZ!�p��UM\��s��s���	lٿ��o��HԔ�WT��_3��_��<,�!�Bs��o#�V`>���+�h����ѵ���z��˴��#�J-"�ն��[�԰T��{�t�v�oq���j�뤭�a~2��$xQ�v�%�}��>Y0o���uU����gKK����mI��nW�N-t��ϧ��LƉ�2O}��b{��X�Ͼ����\��wʥ���]'`r���m�K��'�����K}�;��K�=&�����їb�q���M���7�
�Vv6)�lfҁg�I�|�������SF�{3i3��$���0����i��/M�i�Z�qI��Yö��ֺ����VM� �Xm�S��Q���q��q��´��|��#�ťwϮGv���}P����'z_�_w����g�^���jP�{Z�B�}�	[������T���d�^��H��&��{��{b�b�����^R\0�����=B�"�^��S��n�5�X�����#�n���8��]�7lme]�:rڻڈ�����۵�Y�P�ʷ��J��벟�UT/����Mfc��C�iC`��s�B�Ϭ��3��o߉}&�zK��櫻F
�q55�p�.P��M�x�ok���k^����r��e�+��E;ۑ��~��R(f�=��ɖ�0���g��=,kP��N�� �����\-�y޺���^5� /��]�:+�Ċ�/'��)oN'�Sxz(H��4.�Wݷo���{�jH���[�G�4M}ΔF�+�$���Z9s)X{OPχ˵��uf������Ǫ2Z#�ϴmM��a���F��<���1Q�J�Z���{��B���IO� IO�@�$���$�0$�	&�IO�$ I?�	!I��B���IO���$��BH@�r��$�$�	'�	!I�IO�BH@��B��IO�BH@�p$�	'�$�	'��PVI��E�E=�Η��@���y�d���7ϓ��hG>�W�t���P�7���ϓ�|����4A�x��.Y��g����"'������pw���Z�oG{5Z�ֶ�S޺�r����o[��9���y��k^�v��׽��Y��     ����S��0!� � ��E?!�*�M0       �~��J�       T�@)U�       I�	�T�& 	��Mi4�2$D !���&j5�<��jL��� B?�#t�H@��X��B$� BH����@>��|��������gREA�M@  ��+$ �@1� XL��a���{s����\7�Wm� _ M��a�5�[ *��3�|�?;���zw�0~���*��v�Dݩ�mE.���kM)C�-2**M�_fV��H斝f�h2�X�
Wup���X�ǇE�D�vJ۬7�͒ɴ,e9�A��.DRJ[��^"[WN��!Q�+(5�7��E�᧠�7�^��8t�:/`�N�*��Yo2�&��j�L�ۙl�bD��t�"i�V�tq��-Mդq+�Ѳ*�5X�e�p#Y(nދ�Y�֒f�r�t��b��.<��2�Dx�c%�t%�g2#`�;{���;L��e=���4�
���
�3���)���S�XXYhK���Ӻ�z7mh،"�
�7�`[1�G4$*�-���kw)����wn�j%[��;a���
`�q��H�1�;� )�b��wf\٘!����\�VdV��k`��N��E��2��zv��J⨎�B I�eX�.^��Z��5�P�P`YBR�O�]⡪�ad�Tņ��f\�e�HXK��e���â3Pn�T�;Y5cqm���0��OH�r����]`1=W���`v��.�r�	kei��]�gNݢ�X�Ţ�����%���`����a��4z�����V��k5�e�)Jֺ��m[�0��KJ�"mJIF�,K��tS��-o���ʸ�/��ĝ���r���=CJݏ�t�h�������%��v��ʵ�9�vR=.$��"N�u�l:uhB�	��@U1*�
�0�e������gX����l���i�N&��9�s�z��Y�r��޻u�GVҝ�}��B�;��]��O[���ΤE7�T���un����5�/w`��[�M��h�W���-�8riw]λqL�}�]�2j���u��]�f2�%0�έ���%4�i��YА~;u�����H��OLf���X2��M�"u
{^wI�'"�]ކ�N� �2����E��PPuN�K��rY˻�l�\���k�'}z�vN���K��w5w�wus�r��df)|9.�ǜ��6��=��"�����	�$�����į��YWv�(R�]b�:�F+Ͷ�����d�}ըfF���]Έ���r�v6G"�ewJ�$@p��Uc�-���2c&Х���-���C�I7hg|3K��ˌ�W�s�&�n)��`��\UnX�y"PW�䈍��j�+�b�C��iu���9��;��n�|u���f��r�3�� ��1��T���):Ҹ��ē��� �;Ʊ��׭��TfK�j��C��V���ZK	2���IL?�S�A
�["I��[Ǌ�'T�����Nl�D�xB�-6���ېA��+f'HCP!m�Tl��l�_�]�6�(>�L�e�&�"J�C\1-
m��r^5P���kum4�)���@�ә�1�Zh��l ���%XK[`u����-���I�e��N�P"����6���@�a��&�6����Vn�PVy��T�*�L8�J�o#����
��G����L0@�
ebT�j��(�7�6@fO�-	Ż�3Mi�**���@`�D0鵊,5��:~ h����8g�i	�]�D�Aٶ3"��$#g� �v�Λ�\Oqچ��2Ű5f�?0ٲ�$�l��+��\(��x���'�G�J������d���L)Q��&���B�f�zQ0��n��N��'M��l�R�Fo�ۋT����'	42��0�	�QCGe,`�����l�kU�+�@
�qd��2��dd9�(ݥ�tVB�&p��b��4�- `��o܃H��C�f�cH�W�Y�u��{��w+�ӑ+�Q�5�[U���q��2���V�1�'Vwvq��t}�=��}�o9�u�w�<�Ad�Us��*��H��(|���s���D {쏹~�
=�(�-�>K�
���*3���}��f�@����y-1��Hv:�T%��Wo�Ub,'��	[���4�����z_��H�ef1S�9�e�p2:�$W��3�����u� �{!��k��]>H�r`b�P��fGlq :�A|��5�&���y�眝և@��n9��V�����$�	�ʁf��sZ�.l�En���^r�v3��Un�w]��L�X8Ŗ�&�E��'�Lb>	�В��yޕj�xl?e'Iꮼݰ���'����:��#�%�����-�yA�H��R��hU�Fz��	o�\�����]�*��޾���)�RW�z�3'3����
��'{���$��o0_2�U (�x��C	<@���,���;u��JI���ݬ��6<d�)�0�.�)0��T�f�I�e���<`�t۔���<�59��L���i�w���i6�\9��L'��+%C��2��m��xʚH��!�6�[�5��7��|��#�w40�l*n�LY_"$X,�T^�3H)��d�0�I�a��m��=L1�q`uæe�3�0�Rq�p��H(c���|B ��]}g^�s7y�V�=s�a�`;�0�F�z�<�i�O7@�i����Ƥ�
���he ���ۜ@�x�;�aY���u��2�N$�OS��4���.���6"����Y�>Y{���Xc>s'~���>
j���uI�R�I�9��Y3kqc�]HQo�v-H:���־`Y�BN�YQ�
���Ԋh��Ay�ۮۙ�ݓv��%�VFnJc6��x�X�BK"✤�0������Ŗ�:BQN��$�MM���S���' 
��V)b,X�d޾9�ߎ{ݹ����H,�1q�R�T�Lr�v�fP�Ay�C�`a�8&Y�uCI����S�>1.�e4�RT�C�S�V�I2�^2��s4�f��X$���� z;	��ۚ�D{SZ�������|d��5��?C���a�I��|�M'e0�W�s�d�4�Y�
��fc�0�>��̺fX{��I:�fݦ�0�`x�U��sE�-�baB�)��۽�e�������X�G�Km!��'6��BP�g	�QUl
9�<����&*���)�Z��m*r�LeK�h$Z�Y�9L�il ÞŴ�6�w��IlՄ[��q!�ݳ�hP�	l;u�H��Zk�v�#,�S��@��Q!A^ͯ�6U�/�a��	1d<�E@I�秥\���Q}�(ʡ��MYtg��N��������{��<����rr� GcX]@����J����0���l��WT�(�8c����ٛ5Mo
0�����5E��B�`h)���Xj[jAj�� �;��\O��ܻ����T�"�C[}
Y�FH����oMXB�I0��yڙ%�j�}�OUKTՍԟw33_2��F&u{��]=߅�q�d�YMy�M��L�����s貮�Ud�?���V�]wU�8�$�|�b�G��1
�b��xJqP$R�j�e	�֘�c]�^�ko_{S��.�˜���n�`����l^�/��M��r�B&bҵI҂��wM�K1&z�j��W';��٧��� �{�mX�DF0D#xX����(x |�ƈr��g'Qq�v��a��)�r�Vb�JaA"�0*9x��I$Ą�@�Hi�I�ϛ���|w���x�BI� ���g�BC�d q��@��/��-�)�A�_7�&��+%���!gj
m���vQ>��T=n��F�m��}�'���^�)G=�\TNu��I:��
7�S<�^���1o��j�eB�7�s�'�Z������w4�$ì��� x����4�Z���y��s-��vvk�}M��p1gN�k�*���
�J��ț'.�u�����ͳ�3Zm�,�Uٜh.��2-��׳Rˁ���rMa�+� ��*�+������¶��i�x�I���F;1gX��κ~�1ҭw9!�-���W_��i�ʅ:��5|��G�WX�����Z�
�e�j��@3��B$8U���ܵjZsf�gSєQA�:���7�����^~�G��|�.�	o�͎��l:�GO�޹�b�l�t�T�%D#'!E�A�}dԖ�ҋ��T�_t�:ge��IO��L�P�����C�cbg��J�%�)DD,��c'|ueo���
,R*��,DX �*�v+�k\؝�e��T+D�#Y�����r㺪��]J��}h=�s���״%����H�O����ެY�6�SxGD��8ޮ��SV7IYtd+Ke�n:�g�LV�h��)K�3r��A-���w����Qn�����}^�g8�U���(��N43�BSn��*6$�u�Wor�&����|A��zrv�y�[���p�v&2�5َ��^��R����K�l�u�2�e颧 ��껇Z�w5�ܱ�EU�F;���!�wg�ع���eH��TPU�EC�Տfb�!K+�l�TksK5%5|�c���|.��ɳS3-��������E��[J�<*��u�n���(��'1�f�u7�&6["���ݺ@c���M"(�C:�6Eνwy��� B��}���Ƥ�[�Ѭ�Y#����=��YL0�e�곩�����]�mb ��Z]���n�f7��R����h�ͲhY���AE7��uKQH��1�+ws��y�O��k�Sx����N�I�� �\B�pwcvH:�wgsTء:t�DT���A�)Eb���`X(����(��"c;��v�]����?3���eX��Ʈoz�ϴ�g�DCi{����Y;��E=�e��-lͫ�;��3�v}��v�E��.���=͸��z��e���\�oo*���ګ��33�Ku��h#�� $iܰ%���f�(et����ĴB�1y���y���Y踗�z��S�t��0�|�2�'�Fd$t��\ �����^������a�t^��Wt��&z��l+i����l���ͬ�5��H�p�(�u��1~p��L�:�®�
`�z���أ�o<0u7����y �z��v����Z'1>J�u᱋m��M�����ٶ��V������|���9Ĩ. �C2��(3#�;���<�,��S�f�2j�b�����y����`x}S1�a5t��Ht�¬��j���<N���q�L���B��333
i�奇�~�zZ�3V'b�.�%�yn�J�R�S_ν��ϫ�G)�r�aь�h��^L��I0������6�/U�*u�Ӹ�m�z��͜�5ӏr]�sAt�ϕ�V�]�W��H��n�$�u��V'�	�`�r�+@��aQQ,�W}�����T�mmE�҂��J�1'����B������������1ӣ��l:�4\Qp* ��G�]�DnV�v���!ֽ�|�j�s{�w.7�ة#��R�٥�a�u��Hu%�h@[&a:���q��h��3��  ��	��X@λ��LGN`�Q!SFэ&m�k�d	mWuk6^����*�8�Ǘ6�o���d�`e�56_P�*���\�e������w��w����<��Q.��Z�4���ouA�>�S*,N.r����H}1�5I)���x�v���O:�7�$�j�h[��fF/a�M��r�/ �ઢ��2��3���1|����m|��1���wh�G�"��:��yc]x��{�fc�g!EB=�6[Z9�UZ�0��"��%��iSJ�6b��Q71U��s��y���W;�11�R�+~$�S���tu��޵�G�6������6��F9��`��2��8?2i"���B����_i
��W���X�bJ���m�S��]�Z���x�y���`�M]��;O	YYV�*dXS{iwV����2R׹���s���6���.�����0�{�x���:�p�RQkB�� �e%8���us3���~S�O(T�Z��[BŌm%@��3ŃL����j���\[��A�eR�$�Un�ݔ�S�T���m���=V�U:����iC�]!C���+�9L��^|/��<liV���-��ȥ�
3l+iq\m�^q������a���}#N�!À�Q���"]&E� �4荎�&���q���N��#Շ��ѪXd�U��-�ې�D�
�.��e�HC ��R2a���6�+�/Z!��U]��]5!��]�҂�l�x��m�X1/T�J�ô6���O��vj�'���p�,ʆ�(���ub���[�>!u&-\*�84NH/.�)v�i70OD�T����']&҆���ی��r�4,�iG��Q���J4�mLkʫ��U�=^�<;J)�$r���7FRZ��`���*z^?���/�e>��{}9۳Vf�t"�&�x�я���:�1�⋓P�r��'��25AS�qZ|���c*e{nVݥ��K�ô��4�ꗈ�t�Z�L����6#�F|0�e)�ꅵ�R�E���cuZjۼu�)QԳ�s�%^;���ʫyg+aoH;C�t�q�c�p�ھ4	n6ܓ�.���p��bt�V��ꞯm�ט��RR�wi ��+Y*�2����ⶣ#5�^�8 /	I>|&
A���-aQ-,+X���R֊��b���+eaEUE��}��v�׺ӟ�欀��L�d��Ҥ();�3ɵZ����^��{��[��W\��^wt�5�Grh�$ͅ�,"�X�D�a֣F�2e�y���!�y���[�,V�7i1�n��.Or.��d��ąn$�4oL!4�b�ؗ�Z�T���u�x�.t������ژ�z*r��XulY�XY�n5�ه�� ��g��s��]�F��&�-9��ԟ"&�P`OuF�MP��I�%��M�H��-�#��X8@! �t�[��*�S���OS�u���-�["�+-b~T�1���dB�+�p�&��͈K�]�!l0O@_vf�u�S5���4Ƿo�Xf=%t.�m&>=kj�3��so�HV�C2�!��t��J��V�ҁn�:��[q!�>8o�"BV�'Ls��\�D��i^^���YэRBep9���8�e�Bp�����6}%EN��{"��s��Q�Iin�5��A�$p�Z'
8�C��[t��F�M��9����4��]v==���US:��d#w�ي;#!
q�F��T��c̸�����n�.cQ�$���t�����뚧bl8`$���vJ�گ�),K*'Xʴ�EZ.TM�q=40`�`�kb0V �*�ZԌH���""$��+AV("
�E��( (�cl��P��b�V"�TamQX� ����� ��D�m��n�"�J->WP��%���A�[-ۙmYq;�k�ed%��]w�U�brv���>���zf�����P�d�z�&�lwF� ��r�7��u_k
�DK
�JbD��'9
��h��,nҙ!�.՚�;}՞�h�m79&+���Zr�O���������0)�yDT%�s~:��㹗ޏ�w{/T��CV�QUeB�(
-������k(T�>^PfX��u����t�ܻ���G;N7(S��c�6������n<8��1����b�5l�+�M�:��9����.�dv:�
���"@]��B)iE��s� Db�e���gU}��s9ʞ6&ˣFz����M%�<]�pR:�<p��
��$�︖=Qz���\����cۚ�`��q��{Y9Vj�����r^����Q�A;�6]��ZxȆ�X��<捘�r�����\@bi�[>r��:�s�cg#��8HlƆ��5�Wn�Q�=z&����k�G6l�%���Y[UgBN޸�{ĩ��i�N�ӷ��������j�V]�f8Nm):��������s��IF+����z'q��0#&QB�U*@DR*�Z*�-��P�XT�a �ju��&.�I/&�!��D�^3:H�20`H��1A�ʹ�U���:y]�EM�O+7]X�ޒ8�S�;p��0�U� d�֨�50f�d���w�[G f��3���ॗ���������yޚ�3Sp��1@�v,Kiν��D�� %aQK)ꅭZ�� �ֳS+��N��f���ܣ�Ie��5T���	���U�y���NΓ�Y�F[��Eob9 ��oN�n�Z���~�[<��auP^ �K60�N�2�̒�p�����'�ϐ�h{J�Ny��:-�L$�-�q�OS�� �gi�A���}�������VS��p,�I�	(B��}	�%FF��l51�CHɕ��K"OW�Ѭ�4��/�ʉ��y_Q��;k��X N��@�FX��.�Lt�R5u�8�[��S.��_i��5 p� pdꚉ��9	r�݄$Z�[j��DaG��(S2B����M^:��ں&B ,M�K�%˘\e�]�RZ�DF'QH�ë�ˇ[��k�9��@���l�8m�6�o� K���@ ��`  FAH=�?)�P )$+�t�I}5P�lQ@`��R� �V s ๕e����<�mR�HQP�#�ka-  ���X=Oe�ҿl��d-�7���җ"��Aɹ	�J��ּ���cK�ͻ���IX�WV�K� #�Ky��׽?p!��u$�|���G&� G�.��	P�3����u@u�A�l�/J�>y�G��7�OQPߠr88z� �샤}�:�0m��E7cP*�R0��P���x����/i���ҔDGl�
�{NL^���/Ҝh�Z'���*@��<�_1����d�T@ ����D��:�ؖJ	"���L���pl<,-Y�֦g1 4Vf�n-�[Uw�f��J���o���j��m�J���ؔ�G��]�!o�{�� "��0���:#KoK���j�Ib�|��"V B�^�˳�n���7QlAT��8���I�"��<O`\k8� ��i0w���I�����+�
��6}�e�1��D��EA�w �������������6���#:@��� BШX�! ��Mr1�1`���.;��$iT�*\4�pX*:`N8�қ���B*�JPZ�s��!\V�/�@~% `�;v��<Q�  �O3zG�'�v�A�����/�#�`|�M���ĤB��hgHO�u���a�^\vM��(Gy��ۙr)�~$  �r[+���	&�R�! ������h J^���x)>ނ��fG�8�b-If��@�ߊV�.L,�r� ^�PH� K�t`W�<��+n(0w�[[��{��a�S`��*� G��T0�=ۄ�H�Bȼg;�j�4ؑ�u3X�8.�m��Q�*�;r@kI �St��I� nEϡ�]տRH F�7�
gdvvBV
�;%x�V��J�3R��ci.�3���hYlW/�.�p� ��ޖ