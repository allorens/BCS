BZh91AY&SYb]�$_�pyc����߰����  aF   �    @  (� �k�  P  (  R� P    _ zKkM�)��m��.<>� ���   �� ( ���;�۳vi�zn=�nt��eӹށ���m�	��i�_Ox����(z׬�������iRsd��]�Qh�(�[5Smvʮ�HK��PX������·G;=t��8sm�ut�k�݌Y�Sw�[-��8��*kޔ��y���L�P��y�����{nf
6�TG�����y5�ٻg3�o7�^vqsC�z�v��<���l� xJ���٫�f�<�T�Л5�9�sN�;�:ҙfԭC  �{ oTzۦ�kg��nz��ӷnt.ǻ=�tS�x��������c�nu�:;�z㞲݃�Un8s�Ǻ�-�Y��u�:��9���p��V����h[ooN�y�<��U��=�z�զ�r8u������tha��)�wsU��9���h                    0 H    J��LiR��1�	���C0 F��OЈ�U(�0&�F &� 0i�R��JQ��F&&LL 	���!���L�IM## 0F��&CA���M14$�@M4 @�d�L�'�di��S��@TPC)R�i�a4�F� L�0 Cpr;����B�1yQ8��n�����h!!��Q�A5����?h~�*�?�=�PTQ�rE*�����{(�U� ��� �`��)5�"TeG�V-QU!%��EEȣ���Y$�I$�H)�TT�q?J�����,;
�1;�Y��\k4����ƕ��<H�=	� c&ԒX�@�m
O4�$���CŃ�(kKFA��!�$d�����!�}#�wDQ#
GI��`�a0��Yek�ㅧ�aP�{
\BF>"	&\*$�L���!xc)+)T+�&?d(���S���8_y�^p�eㅆ�����*1�,��"L߼2�\&Y�dW�~4��НY)(p���H�g�r��L�i�J<�,G�bR2I��@�8[�9_hY2�&����@� D�( f����~g�8�S���i8p������+fa���#Q	�HǞ��,{p����j�X�D&H�+(LK�!�� cʄ�<x҆��2��I�bVQ�1�!T�1�Bg�,�Mߖ�ì��0c���P�&�i��M���E�H���C2�ǻ	�g�'(���3%�_I�����{
G�Cp�$c6P���!�8Hd��&P�9�<1�B�F2��aX�}�y�((`�И�`�zC2�
Ę�¶�bя|C$[����CĨmi�xPab��
F?)�%�H��F@���?�G��D�3-��N��
�~Lc��S�H��ʆ<Lf=#���O�E3=��fQ���n���;��3R=!�;��8�&�$c��2�S!�@�<�c��^� fId8T��11���0Ǆ@Ʋ���H`ͷi��њ����J`E���4V�VtG}'G�WF��A����v��t^�*B-j�ƺv�zt�u1���bD��E�_1��,SP�ʱ��c�_Y2���&1�c0��G����2�<?�g�T�cHf���4�1�T���#k�0��)&1���c0����1�.�d<��Ǌ�34�I����f��L����1�o!a#p�`����&P�[�dkT/���R��K��1�fJ��1��@���<��TA�
�X�Z�6�d$e� fi*���N�P�?��C f�1�x�L��x�D1�2�[��0c1�A��1J��3P�>&i#%���Z������f�Q���TP��j(�J.1��F�c(f%G�X�yb0��F<�YpCD��~_09P�`���](b<1�	�їp�1���*j c&d�3^(g�ZYl(`���p��(�&P�X��Ƭ�Ɍd�uG�pC��3Č��c,e�P�ǞQc0�Ψ���MDH�S����j ьnTX�$s�>`�mE�H�~Q3�����1�E��G>�g�aՐ���v��<��D�H�W�<L���"	&���C d�I9�g�y҆`�Z�C(o�,yJ<2�Y�8��B�DCz�:&l�^H�0�e$�C<?\&<�Lx�`��L3ބ�~�ǉ�DX��	��!�;q���o��{�0�1�ǉ�����CK���17-3K����ɿD2|����C4�ɚ1�QF�9ȇi)	0���ΐN�rJ�ްI֓�<W�:A��]:���_d�uV���]:�G�1�,h�������(g�z�L,g����6xc�C<ҷ��-N#L,��cĊ(p��v��7*,���|�x���j,��1�چlՐE|��)�Ѥ�$���r��z�d��X!�c"��C�ǲ�1��Ր1�Q��&�Y#<�C���1�}?&ZR2L(iP�I�[Q�T3i����2�x����҆]��3��c$ѓi���/ԣ��QB$2KJ�DYc,����@�8X�?3?DC$���C�Q"�2[Qy*��~�6���Ii#%D�t���5ڏ	��2�;qaC�'�њ=�CC0y�3W�����I�H��"2����I�c)���11!�1���c<c�2�f?Y,���b#��`��Q��.�3�(��7Dk �$����Ӆ���C���C1�* ���$c������J*S5&h�7	�a�1�L���g�(e���,��K�¡��"//<P̶E��D�k�0{j0Ӽ��}�V��T�#�0ogK�>d7����j �tI�D{R���g�S���K؊I.bԢ�Bd��Nb.�K؉4��2D"5)�(iC��;�_G�S趸=��k��M��Wii����Q}d�!G̪N�'Hv}'H\�*"R6����ci3M�Q�4f*4��������d&`�i������9I��2��!3Fit��}��A�c)�YC����T|�z��?���C��?b�����\/c��z���B�(c��cI`�j�&�"\�c�i��XI��B<1!�mx��ɐ3(e�Z��3Ir������cߕ�Ld?(c-҆h�t���Q�,u�(�
���R?�(d�j,<x��3�<���3[Q�(o�0yJ<2�I)�#���(�0?(z�RA�C�FL-�2�,�ʑ�~Lc���r��j�<S>P�T+����a/�a��>�Mѳ���7͍���|�7�'���4h�gH'q�0靤�g�{iC/�x��1���x�+F#�c�b���2�v��1�����<��Lg���.�V#�0i6D��A?P�3�_�2f��a#�K�$���*�Ȩ�(�ܤ�5�IO!x�ߕ�"d�����av3Y�°��0�<K(�p��̭c*�6�Rװ�c�&�O�BH`��Ǌ7P��zU�Qi1�p�bLƑ'�!�P�P?/��@ǵ
=be�
O�M��/�O2D11�aEg�P�6��H$f����/���S���$�FS�R2?��`��C_x���0�.��Y����A?���&A�P��c�I��*&���v�ؒr!BR��m����\�v�+O����u��o2�I>?�� Ͻ�������A��|2��g�,g'��Irwr���!ҞU���?�<i�����H3�%��=�L��}���\�����/�5���Qm�k�9���M]��(͹#�{2z�>�r�:}0 �����?5�gK���3ݞ�'��������޽��?}$�|L*������ޔ�ȟq7?L4�O�C���I����J���7z}����{���R����yBĔ-��NŹ�3ww�nJM�/��ҝ̘t����l!�� ˽�
<��xeŚ{>��7�م7�>�"�i�w�A��`˹3{4ɳ{�l��n!��$��27a���j���8��{0�7$Qn��w3�×)Ӌ�����f4#��2N*O���l31m��E���V���~cs�4��2�`OZS����}ո<�]�4�-�� c2�Ye3&���C�\�����ޗfɘ�x���N�*�����5u}�i�f�NK�>�ر�m}�8e�8����ge;Ӽ�m�� ��*��	vvs��k-�v�`Ye36q}Գ�f�{.+T,[Y=	igF�]�������,b�{�gw��*�}�}����|�ȿ~\�H'�E��d�K-q��nk�#'�H܃�^i� w���A��Uj���gL
=��5��{�L1��w{�fO����$�!�r��L3����f�bp�9�E�J5�h;#���A�$��� `�Y��}t���,��Na��->��a�%9vI/M��{^t:xJ�wf�l�'ݘCq���.f׮΍�	9Y��|�ܥ���}�����L;��+�c�
�s3��Ŝ�m����_d}��&��	�?��~���^��<?
+�;龨)����~7o��zOi��S���Y<����S��6o�!�ja~�&K���efn{�{�g�,�=o�v��B�W/ajly�c�%��G�����v������s�W��7��!��c�ɾ�j��އ�+�d����t�e���(�������2�@J�O�V)~0�W�\�c��;��Q�X'�e�w��:3����*<l<�aΔ�D�N�Fy�����q�ůi��fv�9I��z:���"��b��W�q�!��\�����t�_��sg���x�і菭զ���)�@�|Os�!�-�gY�2�mv�^/��(��cuiyB.A�~�/-A+�L1�9��Ttz4�Ÿe�t'����E��-@�]���8�uL���H���E����䭶��l�"��{������^c����Fݝ��FL�P����N�f6G�O|�.����X����]��M/���N�ϢCzǣ���ww;��pS_�k4�|0IF!�d"��nN�f�<���e٥�<��H}��կޗ2?��;�n�3��c��<]�d��s}��ޞ��PB��tnG�&���t�rBIIl��êg{w �Cy/L��}��[��Tnd���������k�ۃ�=�Q_Q�;��Ǳ��� ��c[�^�s���r��.��ֻ�L�b��tKGpc�[�k}������;�9c�ͫ�HǙ����x��k߾M�
;Kff'���Q������tZ�d���m���V���ۿf���_�#�3�;zZt���сO��2l-ǅ�d���t�1��`��l������.n̗~��{���y~�{�n2̛��X�5����骊����]y~usB���7����;����������5���Ϸ����K�ů�ݽ��Kh�{��w+�޵�����峂�����e�ϓ�G��=���ܝ��#w��!����U�s�ݔ��1�zVv|x,u?X���̐��͙��1P��w�2�*�ٙ���f��ҋ]���T�ϫ�f��?�ם��w�*�W�R�	��ь�g=���ݰ/��駻�6H|2M���ݒz}�0�����2��;��E��~�W��9ٗ^۰�=�k�w'a��1���_�w�@<r|<7֕	�߲ﴠo�_�:i,{�zt�۹ϝ��x���.�s�F�"N^�P����K��olp�d	qܻ6�}ެ�{���/�����3����÷w�9��ٕy+Q��mO��eo�H���K��{��O�>p��_/�^�ϱ�6N�Vc�۳frX�u3;{*�ޝ�|6?/ �s�:һ��Zg������ @���8���Ͷ�욤�,��A�= ��/�>%�+��<��5^7�J�?��wt������(�gJ}ѳ9����=r|?va�0���퇳i�I���$�(��}��gTo ��\�a�����Y�ö��cd0���݇wc��iJ�Q߃��=����b���-�2�M׋X ��������yO�햋��z��#!  <9����$�9!����};�9���$:=��U�~U�\�u=��R<����8��>�p�(v���n�O�1�+�� ��.d�o%Bb�xC�a�U|����:J��G(��AW��m���}٦0��;�^�,���vt��H�f{}0s�M��?�`u��5K���N�u�8
�R�{>�b��8����[<f\���|��4
Q�T�Jk�4Q��������3-�w�L���2��ߝ�Y�{�d$N�qcɤYv�G~��ݝ�u��M�<�6@2���~��͑��ϑ���qѷ!�ڼ���{��e��(�	'�^�ھ����%�>�H2d�isgfL03�{%�b��6��Gw �'%�����@*fd��{��<� I$����5����g�o2K����6�d �����M�7�8�پ���:<�x�w��܃����+ߝ��ӧ}�s\�Ǘ��3^��I)���i�v��ju7��愧�f{0��zr��rM���{�(��	�Hb�0}fid�^}v�Iv�LS�3�by�z�i�^f�?#"]�'N�vu<vL�)�K4k�x�M�0�U�;?�zɆʬmk����y!�*=0�Bw��X�����^�����z`b��x\�M���Ӵ��!	���/�Qjf��5\Ȼ�$]r�*�-I��ؕ�����c�Дʺ5�8�l����f[X���Ch5�4k��5u��k��v֗j���ٶ7Qз6�����R�ҷCL]Cg+q`���`5�vD��J�^ĚkB'R5�%�ޥ�w��ϵ���I�ݜy{���`ֺÑ�EX�h̒`T>��r��%j.���iD!a`�^Q���ͣfk�,u��Izh��XpO�w��KH*[J���B7�*ՖCn�5	5i`�V!��ޥ/Z�";Ws�[.�Ǝ���B6iL�"cm���ڬ��ʐ!f�+���c1t��֩6$��rh�bh�-c�k�_9L��X��y�Y� &إ�3��8�g\H[W)"qK�� X�Hi�_M�,r'6�&w/���p�kTQq]\�י�]�Q]]�I	Mx�n���b�ml��0f�5�E)(�U��J:����2�}�-̠M��K8��  6���
��LɠO7���}�湼�CeK�B� ��}I<�=-~ۭ}+{ܰ@6-��W��#�c-j��:�ĺ�&�Ժ���B�7v��W.B�h�n��d`��zބ�w���w�SS�u���9�4�]��;OB�#\�>��b-(�)���%��ҁ�֍^Zq�q0Ei $��FT����H�*��h`ܼL�V3��(�`	��Eq�' �-�I35�\�� �9�KD<��(D����Ǣ|r�W�s)\L�R�'��c
)0��_���� h�Ą)��>Yg��m��2���m٘_F��&�RG��U���:֋q>0D���Ӫ�$�S���F⋬d���L62�!��ޞԓ���ؤ�$��e���,q[�8���Vb�9H�{ac�Kk���K�C$��"&F@�D\�������hZ���g`��O���#��a�G���|qv�~�3L`�!��`^�UklBj˴����6���.�h�4(.䧒����4�4��+j��Gpϧy>�n4ii�K���xLMĩ1�_��Z�%к@���0��la^�NS�s�yj�㲰DPV٦�Hlۊ����x�B�D<J�����=�Oq�XEE/����G��?��?����۶�m�ޱ��m�M��x�6ۦ�~m�m������m�i��o��m�n[m�m�6�m�����m���m��ݶ��s||!�	�	-D�ԑ�a���lt�r�m�nm��m��m��۶ܶۦ�~m�M��Ȼ���6�m���m��6�n�r�n�m������6�o�m����m��$}RЅ�K`�E�����cm��7�۶ܶۦ�~nܷM����m��m��7��y���X�~m�m���m��m��z�m��-��ߛm�m�6��x��m��}�����}=ܻ��oX�m����m�n[m�m�6ܶ�vǭ6�m���y�����r�m����6��nm��m�����vۖ�m�n[m�|�7�s��9�5bеȑ�@�.!P$۴ۼyE`F0a �|�y�^� @9v��')��q4!��ac,g�P2�Q#	�0c�2FI��0f�h�C4��h�`�c��x�1�1c��	��1�3Fx��d1�H�����
�Í6��mU��8�������c�b�d`��d��1��b��i#4`��4��3x��4f�`��xg�H�!���3�1���� `��@��bD��N8��;$����9���bF����h��n\��bFb�k���ͭb�qT��&혓s�k����#���F�55�Y[ts��m�7L�&seD-���U�:�umn��L{޾�MM���)�!�Vɗn,�85ш\�f.�f%"���G6R%��#�G]
0�v6B<��\H��LYZD�+n`P�2a�$�JF�r�3;XCm�lk��d�̗@��i��ST��]�~}}�Yb�[-ӱ��\�̺����	B���ǳia4bؕ�1��DY{%u�#�Ԩ�:���L2Ǖ��k�a�X� L�vq�.��%� �B%�����j��p{ݝ@"d���n3���k
��mP)�6ۮ;g׳Ԧ�n�z��r�~6��7�E5��G{����P��k�z6��/�ԙ���~��z��SA\%�i~�|��b{��5��]WYe� �.�۪�(���1���\�kK��1�h�`�6�e���=`�{Y_����ǧ��eYjx���LJʦ"Gk Kr��X"�,$�&~+��-�Ŧ[�S-���ΗKA�Kv����V�]QԘ�.�+�m�d(0�MM��KWX���KM��8���f�z��M�,��5��i��.�.Ԙn��%��Q,�n�����c���\��[N-QkQ�\�H��M0[l��ʯ��.
jչ�֕�6۵�f��ٚkyv�q�B��u���mT+.�if�ݦ�%5/ϣ�{��3�6 6ͥ���^�֙���,�m�Ym]�hC����4��lLU�Ģ\�$ָ�im���.���c#��᧬�Q��Y��릖�T��Ʃ��Զ�iVVa�bXuҖ��[,PL�b�^U��&���nbR2�f��o$w��պ��e���ˢ�t%۵�]B�P��Ĺг:*Y\hL�\���M]5����蹾�v�{-�j��G��d��I��@w�e4�B��6�s�m����و�fv�j�F겶%���qI�XQ��Y%Vb(�f@��&Dc0�5��q�i�3d�%�2�fT��2Kt�fj�`&�n���γ[�T��뙵��k����e-�_}l���R��2X��Z�8�	��!rX;[�0�n�5�YKs�M,˙�ףf��%��i�t�P�5�A]���y�ٙ���˾�>�����333;�>���㻻��3333������������>� �q�i�1������i�����V����lrJՍY�J�Mn��v�՚�6m�����l��ًl5&� ��h	M3�v���	z���8	sYmW���6�	��Z��U�,���5�Xm���k�6��6l�k.Ś8�V-�̹ve����7�x"� j,6u�mAn(�vn�ଫ.��R�收�S��b�S[X@�T\��69�)���f)fa�'��I�1��8������9��(�&��S�d�\]Y5�&.W0;�MYV�:����e$�)�KZ�����_up�< v�#��`umR+D/P;UW��h�E�A�]��3r����3L����K|ѧ��d�C(MѳU�~�zL�)�*䖘Bf8�֋Ɏ�����7���փ�5,���Z��x�.���u�=<2�2FI��4e��?P}��Ptmp�Ԇ��0�~X|�6�i��ȶ�ŽD�M�e�Uh� ��v��&]�nX1��&,�%�q����K�CW��[F[=�O��k�����,�f����%0�(��+�F%dA��3M4c0f##$�O2�4($��2A��%O���'_��ɚ00����O�\'�i��.U�e���7sR�^M\�f>��T)l���)e��h�	��Lu4bZ};�[p�u��n��Bgڥ���mZ���3j1�mO#��|����0�K4ӆ3aC$c$d�i��Ν{	A+�QtA8�hM�P��h�ϟ�^2���[-.���$\o9���f�m֍G�cmkL�h�Z"�sG	&cU���k*��l�V�7Gy�$&��	Xh��(��8���	#���xe�1�c0f2F2FI��4e�����Ծ��������꽥b|v�g�4�S�}�׃'�F�ǹ�K1�VJ�֚��\x�Ƣd5�����X��V�(����+aF8�hd����$�:����:/��h�R�e��O��O���S���ګ�FU
#�R�ɶ�|�1�%SR�O³�DP�U�M��ꏄ7Ͼ6h�G�sK�"C�h������+���a���}D�4�hM�F�ƕ�Q�c괵�Xb%�+���[O�Q�D'm��+��GT�3�m�^=z��8�Ǭ�##$�O2�c�x��ȗ�e=�__��2�=gr��6n�2f#�`p��$��5c��7��>���F�	 Xѐ��8`J8��-��^]��k�rb6�a;&��aKXHV�E��̒����ٗ�I�/Q��!;F��)��r�)�����~hyc�-�>|���$�x��0f2F2FI��|��xY�%F��ƶ��ѵUҦ�`o[!tp���XeG��.����z��AoZZжҍ�wp�#d[yxԈl�u��6��a��2�'�P���e�ZZ��DE��I7�eF��X0�1f1�%{|s�孵1c��۫W/&ʾ�>�jQ�?}�Kc4c4f�FH�H�4�ƌ��TL1* ���K�D�����z|����N�̓N��`I.��.P2eV6G��
%$�ocZ��j�m�ˌG溺�Z�Ɇ���4}bM����Wyj�%X�K�R��]��6v����}#4�a�4f�FH�H�4�ƌ��M?�j
P*I|���(Q�(b��n������Ȏ��Ae|�5��	<�ca��_MX_�y���֭�|d�/&�t��T��R�UJP+cV�[9�f<,J�e��c"�|�&'�ԗ�14!o�M�o��k|m�i�?T��\=!��^���������"޼;��dS�k{�����řw:����G=ģO�S�G�MCzE,�����N�Z�cO�oZ�9�ꬬ0�h7��U��G	��(��F�ﲍ����:L�5Z�3p5�\k�q�ա5+.�X�ֵV��wѓճU�F���R?������4�F1�X�a$ce�_>m��*������m����IK+�6EFX%Y��Ӵq�����ƛ=����9���}���䯞�O1A|�S$�[U�,ɣq���ŁÕ�S��l�W����`�{�^��{�vf<L�?��8�$�4g��b�Q�ɐ��ǡ.=>4L������O��CD��GGL�#�#����i�1p�/�di�H��Ƒ��� ᑥ�G��p��qAҸ���4�\I�8�B��G�#�=+��q3��h���<���$�D�pQ�ѢX���_�	��>�x�x|>4O��8\qq$�$p.��q��^?g������I�a�&N!���g���i�1p�-�q<A\2,Z.0��F��œ�ǈ�qGJ�<q,���p�a.0�K�E�~"���~'��C�)O���6~&'�ó�x9Q��(����_�b���Af�������8�#"_���kPx!��v~�ng|w���vQmA����\�i�����߾��Y��^S0��}�b���vffff��>;����w333��;����ww33�����������;��q�q����8��,��:l��d�R>UTDD0X��T�5W���U��`�
��1d�������VR|�K�#4/m����|�Ő�T�TS,A���4�qIPMl�UX}�x|J"R�X�Cb-MF����z1�v�M�S��$�FO������lM�1$ʏ�6g�YT�,�Oј��ǚ�*{*2đ�WL�E���)���|��1�+SǄYA}��Q��7EW��&����M�`��"b,bRU!lb=Uh����,e��8�N<P�Y�\��u�VڥR},���Va�aױ���"��"���Kb`����lm�J'��F�U�o#�9�r`��1��F���j�p�q�g�s��:�T�8��,Ҫ�P�?J��l$�ɳʷ9��I�g�UV�~�Fx�ŉjX��1%Kbvu�*��o�CV52���[�֦�#�}Q>%"%�Th;��U4��C�%�~���sDQ�)ʢ���{n"}*i���5RaRL��)L/�U�-��SB`�!U��I2���8��,O�S����k��W�\~u��6��A�q�2�q��{�6�Н����d���h�4�
���"R%vdՊ�O�Ğ���yj�#�A�nfMi㢒qC���V5k$EĈ���Q7&����������R3X�{B��l��Y�f.���hO@�B}{i��λ��""���F߽�~�eD��)����gnH�sw>-���:�Σ	��Ϲ�w�m�|x��F!`檒���#ņ哬�ʫq`��}��dʧ�26Ğ�b#-�'�&UU�*4�3O
maȣBG����f2Ļ��c0���Ŭ�ԙ�`{G�$ʪ�<���M0j�
z�fR6��v��d77���Z�Mg�^}_f��B��|�E��4�T�g2��"�J�c�FU/\��d���X�x��&UU�����a��EJ��f�!�U~�=���"v$!1�&���\X�����ض���dp޲�V*��	U�'�RB��P��p�4�J�~�d���8Y�+O]|��_�xۓ�q�q'(c,gP������?L����UET݌�Ďy?<����ꍐ�Є�i�TMw�N�q$�4&�j��j��	
�%�m���,3g��u&����[��B^��� F����8�6p�F��VPg�n�*��KX5d�0k*�Tuو�Y&��-�RR�����[�؄!ZKQIY�Z��a��$�R�b�<XlDMq���[�CH(F�Lj�D�I1;�w!����!���e8'�UV&a�d�Wg,*��"�lY�ˌa�曲ɏm���J��%�i-���L�:�Y��=X�Zܲa�UX��hS��G���)A�j�+ @������?�Y�8�8��1�:x����W��p�UZD@�Ak(��n*��~Q��a7Sj�Ė'�bɶ"�}�1�L*ǿ��qa�UrJ0�a⚴��+Eʯ}�]����(!��D&UU����F*x��M,���DHq�_���-� �T-$!�:r@�	�b�C<�N%уV�3qH�_��	��\�p΍��1�"v��+?j�I$Ά*\1&*Yd�Ll�v�Ⲫ��o�g�^��|k�؎����J�okvQ�\�ȼ�E��V"��0�$�����������+D%T�J��������4C�q��;gݻ�i<�L��T["�e�!���#O���[z�����8�?:çq�2�q��s�?�}j��{�3f~������(̯B/ju�!t��(��R�����V F� q8|�J��a&i�d�Vj�.*�%Gܷ1͇cl�ڦ"����<4���*��Z(9�~����W�1����V��yq$�jWʉ���jW����I�x�*�JQ�/닉�OG��ʟE�F#U�♧'��?2�L�c�&"�,�S����Xc��)�ed�V*3�����CU-�kjbT��n"uF�ě�$�Uq#*U5d���LD�S
�Xʚ�f&�L)�ف�dj,NY:�[4�zXTX0��SRad�
aZ�%�#��h�?��q�q'(c,g~�=S��>�����D�B^�2f[���q��x�vH��1�0�E2��7��J�@lxE�C)������x�%��$v�\j�bV��ހ��{_Vz29��:ۃ�
س��ZY�����zxr�o�D��nW�}3)I2*���}����$2��g�hV�]��,�Rz�~�=S&ԛ�:��/+`f,�Rf<V#�,O�4��NE�TʛX3c1Q��a)E)bxj�p<|��]��Znǌ0��Z}�4�x�bQ�	[��![��D��R%���Y��X~���l�򧵵1�g�b��T��a�b*a,L���O��a�7*9,1g5c|��b�^Uli��_��І����5���=Po�]7��|S ?d}��� �s�D��X�5c.���Y��Q2�*@�����b}�"C��"X���D�b6tE�q�~?��q�q'(gM�<p���G엍�2��*�%���fU��E1��ʙ�aO�곈�%j�4'�D4	_�@��%4I���e�d�FV�d�q�7����x��e���J�$�sBJ����-|5VcT4�C��u��
فP��@��	�??l��F�VD����jf��[Z�L=��\��0TC�(h��5�"Bτ6!�aV&�HX��zEV3�YF���O�?E>Vaر���z��"��5�s�&7�`"s��ه���g�aƌ���,���� �8�Cc8ÿ/� � �:RH�O%N��K�F�S�a��=�%��
N&���I�}��)�F�*�+Ic1Bt������nnoV�x�q@C^~�I�prܜ�#l���w��|jK���abn��[�7��ޙ�U0��bq�'��_+��~��B%��r����%;VY��U3�y��e6��^���K,�k�,LHZ|YXv�J�g�eO�cj�[��	}e�T�W�۬�[U�)[��|�����?��q�q'(c,gw�?�W�U������ ���WS�?G猵^��LEO�̫U�|a�4@D!jr3�f7�ڲ7���$9�sy��ս]���c���M>*����)ȭ)�S
�]%|!�_���BB��	[�"
n�%U׋,��	bŸ�=�Ei��n2j��r2�_�v:ʔ"���D$�\����	F�6n��v�nS���~G�̜��f�����Eb�(�S(�uZ	E����&҂`�I�P���������K��<	���Q�a�0|Y<XH'���x�!0�a�����?�%��i��3�2<+8�.�i�2��ƑƑ�'M#ŐA� \i.8���q�p.(� �T"8
'�8�/���q���apG�Đ��&pt*8
dSD����=FŒ!�	��'�Ɖ���<>/ODG��\G%$p��<-8�e/�~?���q�g�gi�9�8�.6B\-8r��b��E�	��BV/BGU��#����־/I����~�ʞ�����<0��C���g�|0����8��٤q���_�w�H��1V�?�qY����MOqב7 *�ιA�j�k
�-�#�I5}�Cp�`���!�$�|�[���s��ηؤ�ǚ�X/�r�筵�(�|��Y�24&��~�D��$u��X�kkJ;2:.ƃ�����d��튉�[\Ǒ��(`��G�m���3��K���-[�~�`�Ҷ�Ft{�O�m}�9|bn��"��2�]Ջn�mT��d�0�*ndX@V6�i����N�{u�A�쮻rئ9�c��0�EvD�W��m�EV���?fU�Bz�
��7�~.����ۙL��sj�Tч
<D���}���U[�wxY��]Ya+���
�{� C�xT藏��h��N�b�dg�/�Tj�ʩ��6Vb��in���1Uh��*��T1QO�D���CK*g2A��{hK�kv�v�����,�V	�RmFôn�M�{&͛	qO�m�оn�Ǧ�݋CA8Kt�Xw�[�c��;1��;V6Y�F���IFi�*�olŭt���\g_���[��������m������9��yۻ���ɶ�{ۻ�����31���q�q'xc,gl�q�V����-iL,���m2��f�`)6�XSf��(4`��5��6�����b�V'���WD�*@�Ա�f��˵�M[b�`��~+}�U��a3�5Ib�(��N	�;2ƴ��+��VѶ}��yXbY��P�	f]
���l9]u(�� ��(跢�2�M�/��R��a{8��ȶ�h�sx�т�^qA���Ѵ����q�T���sG2a{UTBg�����~��n�{�3$��b�Tf�F5����^�%b.S�P��׻�Sr]�Ͽ��~%���T�n�!��A��e5!�u��������a�4b~j�]�S����6@���d�Ԭ���+�uX�y%Y{�rD*��8���߭���7#�,4�����<�m��xf��|��TZU�����W�/����z�%��%�$6h�Q�A*pp�?����g��e�L8ӎ�8����3�QĞ���Pw�1U�UQf�3D�������y=%��h�:]�6���|�B�!�9VM����F��ف��I��&��v:�F��feeO&2�O���,OQ�ծ	�9��09�澒-��q6��a\_�Ƞ�����i��|����\>=�̳3��!�:��G�^	F�l���R��6,0.��X`��[��a���?�Y�A��A�q'�2�q���mf���.�]5�UD>>�����H~��f7�����> j�ag�^S�h�|�9W�+��0 X@�˪�,���s�ʐ*p�L���W��k����<�����H]���`X�|��j���9^��Tl�#�_*��<�뿯�w,lٳ��F�G}[j׬͟G���z��~}�knm�����Xx����θ��W�(�J��~�~E��*�E,J��f��)�F�t�@ٕ2���~�׍!ʨ��G�W%��Y}=��.���aeͧ�/�ˬ���>/ã��Xr���Xk��Oѭ}ieo'T��X�O�M2�,���f��-�$�|eo��-܂r�В�d�	D��AK4B�ōʦXy�r���;cnF0�9;�e��:׍��Xq�����._52�=}�V_0����_��x��#�8��(c,g.^��ǩW�
\*�;�y�ڬ�U�PG����-�̖f�N^�,[-a��ܯZ��t0M�H.֡�zF�x�W�&L���RQ��I۽��  BY��o\�"�����˘������f'���/z�k#�>��f����$V�s����p"�	�r��^9gO����b�l\��<��?��6꺁��T�������W(ڮ�����,��0���nYe�,��u�i�x�Q�~ŬW����=}=e��V~^����:�}��E���NL� �_��m��@��qj��gM�P�=Ֆl�a��2��F�_�a��:���|q�u�Zt��c8�뮅�te�J�ʟ]�vgY׭��gC��?��|8��f���϶4ؔ���?�2�o}�y���]��ϡ���UTC+�r�VϨ��,�__�iA�w<�|��,$ߊ�\��0�0�_�<$p�9<;�8x���\�f�/��#
X���h��Æ��߬�^U�٢2&i��R�y�6ܬ/Ʃc�����D�ٕ�Y�:8W;�r����i��\WYjn~����Xz~~e�3�?~?�ƃ�8�$g�l�㆏���qUQiG��F��Ee{-�z�mL�'�rc
�q�%(ç<"=���ݴ`�;�+���?,X��ƚZ��rh��v���2B^TK��u���^Q����ߋ�H|?���M~�"��4h/�C�ƫ�ύ���X�lơm���z�,���\,����ab��0c�?}G8z�F��'�F�a�Ez�S�ng������z����<m����(�Fxe���.�E*��}�:�UU�z�Iwuta� �����7�x�׫TXe����w�5��&H�*�l�4v�e��f�ѧ�e���a����F�}��^�}s��y[���n�~�2y?;-MƦ�>��|�Ob�ב�];d���ѐ�t|n��lOP����0�!e�Y��3��<h1��(�Fxe��ws0��W�)yyr"�9%�ŋ7�%:iZI��^�I 쵞�p{�EN"�i74���J����J�¦X���}|�3XZ�L�s-��  ��넟Ͽe��[��X�<͌	����;3���~wݵ����Ъ>{��p)��n?�~��nD7��/wk�6D�2�=G���K�O~��ch����L���I��b�d]�s_r�_�4j�e؟�d�g��sdg��B
Q~�D5FE�Q�zg踎5����Q��<����b͇�~ ��?:f��#���e���N=m=�9��޽��k��?>a���O��Y�A�GqG3�,gn����1��;J���9D5񪰶��!�鼭�4aNk���*�<$���ä"�hь�;?G<��;W3^���2���xj�_���g�L�ZW��Y�1�k!�.��*H�p�E,h���6J=�~�ܸp��UXs��r��k�|>����.5��m��U�La�ϝg���,�A�d1q�A�Y�`��K��x�xp�>,����ŧ�x�é)�q���Ƒ�f)��T,?~?Bk�3��G��#EƑƓ�����0�OE���|Omk��|x�6O
�0�<ap�x��0�p�ҸDq�q-$�_.Gqv0���׈B�A.��<Bx����!<YO���g���q�q$.
#���p�\T.<a\\/���G��_�#�Õ��^<-d�i�1p�db\GG�3���ӈ��fB�,^:��i���Q�Y�q��a��\C���-��d<60<A<A
q#�##�Q�㈳N'
�ձ�m��}���֝���)��&�Kh����P���[�mM]�m��f���W�^�ř��us+K}2���3�J���h�|Ü�ӎ3�3�Z߄nO#<�=$|{�LI~mun�?ѻH[p�����7�ۻ����6�os�ww{�sm��ۻ��ܹ���������8Í8�N,��!�qGq�Ξ8i�EUD,�hY>���;�ڛ{2��<4��̲��r�<y<�)���a�6��`���o�F8�$�KK�.7Ə���}F�śR��������o�������~�m>m�oV��a�}1����V���6@�T�h���e���)���l�����|���Wu��<h鳧�<���B]_�EUQ	D7^y�F\��p�<2���j�q�f��ِ���j�mn~�0�6f9�.�P�k�>7V=?�~���Q���1�Y�GѦj3���sJ�|}�Q�{[rz��2�~��o�����l�AZ�?AMQ��Յ�]<s�h���OB����z��X~���a�d|�i���?`�8�ƃ�q�0�Ξ8sW.���c��̭
F�K�1Q�e�Ƙ�{�$��yB��Z�N�+i��Y��I���2H��J�j|mlR���֗;Z�Ω�7i��+�rPU�t q>�y޺UGӮ�.�����zm�I��)�7S��{�<���y=�f���Y���5���j�$YMp�h�颚����PB>��ѕa�7��v�[���i�iM>�Vߚjo�_�l�u���%z\��جͬ����Qg�^aV���m�<�7�G���֣,C��̵nb&ED��-�eݔ��zɇX`�5f?oXY�6�I&�,�FX�?2�b�qG:l���h� ���4��^Y-�j4� �R%-*�U�Pk�E���UE�[B� �"�ޙ�I�UTCS�]a��~녟�w���3���5�a���br�V~��H5��>����}�]��HQFC�h7D�1E��}���A���A-[)x^2)m-�-d��Ĳ��>�{.f�r%i^���MQ��Ҭ�D����U�Z�B|e|Y����?>e1�,/����m�?Q���3ҩNA����7���r�q�xÍ�~~~|���1�8����a���C1CV�j�F
�����������ݍ�l�,��/�`��m���lL�߽�����iyt��tp�.�ee	�ՠ��h�%'d�������i��|�#�S��q��ϧ
�2��|jKm�Rm6�XG�|HIda�3N,��!�qGp�,go�iL�T�{f�����"�M��8d^��(����� �=G�nI}GD<Bx�	���te`��u-y.Y�9��(��9J9g*����"�b�*��D����R�Br�|}W�ʰ�5��:�����X!�'��E}�FD�v�Z9P�Sm�����K,C�J6Y�,:$~Tޟ��?=-�����Xe��>~~q�4�3�(�e��߽����	>���/�q�Z��Y2ӭd��]�Oki9$�:�a��Y�ܯ��t��w����YB�ͻv���d�1�ֳU������Oc���@ !(�?^��I���:��w6�_�8�ۑ>���u���ߩ��p��ù̙��8��UW��<��?��G��J�%xH�v��p�� 4Y����>4l��,,�/pEW5GY��%����S���U�����4��XH"{�؃�hD>>��5�d�����4@��i��%����MiFK�r�e%��m�n$���hi��19�:��2���0ݛf8�O^2뎾u�zq��qG��q��UU#�I!FqUQ��)�5j�>5�aX7ʼ�'Z�������g�<j94d�´���ǉ��g̺����ݰ�~>���~����6���8*X���[`V���3�̩c9Z�,�c�уye�7]&�D����I?6s�lٺ ӄ( �ǉ8�~4�N,��!��(�,gw���]?@�$�B��Yni�J�����kmm��bs�������ҩ�z���=��e�J�χ�h�B{ZwvN^fL��_���cy-�оՍIJ}�F�8a�	]?J�h�����,�D�+F
%�RX~ ��]~5Z�z�H�'Ԧ�����V�\��/�̸���������ޜq]:0��FΞ8{�T$T⪢�->�.��� <h�s��!����/;0f^�l�/���-�RA���~�h�����3.��)g���m�'��]��Kg�8Cj�!7.w%l?Qtp��*7F�k��ԃ�)?Pܢ	qj�Q�{�$�r���	�0��"�OǊf����8&#�#'b�OqdY2�G�"E�Ĉ��OA�B����'E�#�ѓ���"�p��+��~:�b?F~J0�4�</B"��p���OG��∐��\xDp��8�(�0���q�q�q��x��'I�.�"x����ii��, ᠕�O�'�'�����H�H�p�.#ŜO�"�#=�4��~�I�����o�������.:��?�!��6R��'R\&.,�K��Hĸ�I��WV��x\���\x��Դ�t�<>�c�8Cŧ�O��E�᱂� � ���&�gHx�����x�|x��M�w2���Z:�QTF5�������#���\	�A�η@��f��Ď�sqb��W���dɌ\�q�&TF۶U�q�(d�2-̾�)��-Ȕm�
�` r��^A�׈��R�"�(Ȧ6fQx����g��B���\i�}:&�'0�}�p
��S"�d�31�,Q7Ǎ��d�'LJ��u���޷�U%k D�BQx��d����]1,mB\��t�������ثpp'f)d���bu�ۻ���˪:�o�&Ad�<�1cC��1��:�F�Pv�k'�_��_���{�D5qR%hEM�����Lz�w]�׳:E�Ř�E�E��w�vߛm��k��ºK%M�[���q�傁-��ih.�[Dj�
\h�m��]Z�L��C���Cct�}f`�Rx��镳W[�Ƕ	RG���f�����3[NO��B�G1�x���E�e��X�%�1����4�r�L��C"�1YI ��~�����ۻ����m��������ow;ww{���m��n��w�qĖq��,��!��(�,g��������,m-��f0f,k�� %��*5��arYvv��j���5=�7c�%�x5�n#�m�DwYm���]{WQkj��F]��f��A��%�*Ț��YVh�����3D@��kq�`�������Z��ND��;m/ Ec����.���.vJ�\���:�a���AI���hb���f��1��u`j�����������#mL	4z�%KIlo%-����s��s�Ѯ�g�>��g�b��Z}��Q���&�WA}�_���ힹ���1���f�o�_���<��ܛ+�ZF������a��鉗篞�X��<������G��=����]�5�l��&c�����C�_���:/���d��~ި�#�����HY������ḏe+c�$&����L�Q��͟Q����F�,֖?�I?AG�<"�4�ŜqƟ�<`1�c8��8e�3�:AЁd@��N*�!�?h�T_�en�C��$h�4%@�5u�}���J�Q�Q
n"��!����[�]�j�4}�t~����4���Ϙ�/,��Yj��(��������������f���r�r��~�wl����hN�q�i���sƞy��l���#��cF3���Ɵ�<`1�c8��8fΜ<p�r��d�ٕ�UTC�?-4;�����a�W�/�*)^+n��]8��<n2⧛�)�_a_��M�ō����<	��B���C�x�H�������ů��l���(����K6�f7g�l5����^uG��(�������H��FiG�q��b�?Q�,e�`��B&Z��*�!��Z�MlH~�8�/BBs�Brx>���6n�k�6��j�LĪo�8O����I�ŏc듻[VՌ<W���D%$�Ռ~��X9�|j���7G���a�Џ����l�i��錐�K��Ҝп/����(��elNj�SkV�/����:�|�m��q?�Ɵ�<`1�c$�8e����}�mbbD>j��7��$��R�Y�OY���L-���u����&�9Y�����2���d�Y�5���۔���Q8* 	J���>̏n?�Fvw%��P~���x.�gT����������M'��ߔ;$���0nflhO߫�P�?CkQ�����UL��ō�_=�b����0Y*s��:k��Ie��a��X�T��[�i���g��2��:?1�����t�������-�G���\�x����4����f��y5v3u1��g/��_(Q�D�`�?q��a��C'�8e���9��귮��N�oj�����)!�Yn�����ڰ�+�_�����e�V��.2����O^2v|����:�ݚ$���45�%P��ߺŒ��8A~k荜�!�(�D���-��L��0h�p2���V~�ʜ�Yq��cޮZ��xx���j�o�~�Twn�ą���"$��~0�0њ~0��!���0��gM�8���F�Q�)nG�Sj��v���Bi,�e�t����4a�6`'�u$�,�!�0�BQ�,�<�3]�-kc�fF���/^�ԅ�@�_A�c�hֵ��;F~6	��F�B�!p��nNՄ�k��Ut'�)i(��L��J�k�f�!�J:h�|?W�4�@��*�j���a�֯8���*�rݷ���ȭ�z�O��:i����2FqG��8þ	J�!t@��x~��x���>-����)����+F[Kf�ׄ���9Ő��b�t�W�[�M�,�Yi�=�4Ұ<G9G	��م�؈Jk���(�yw�`;WT&�8X@���n��f��s�筶SO��i�5o���ńYǊ,ќi�0�1�3�:l��+5�ʈZ]����i�l%&��J2��1�D�M�D����&w%`�Ƞm�1E�\���v���ҲpM7N>�\M�� BRw�u�ﻸ��j�rg?B�I���<W��=��+-�7ط�X�˗1?v,Y���s{mocA<����w�5ϣ�R2A�]��f���6~� 4BP�8a�ޖ^�Ր��%���:p�d���}�:�3��L�)eVM0�S���>fx�뇼�>�Y94���O�r�l�?��Oҏ@��e۶-�ɕ��E"���+v� w��ˣ�h� ���	8C����z�5���<Q�4јx�c�H�(�:h���Ĉ�UQ�7Gퟍ���H��1;�kF�(ٕW��u��KV+����*�e{�q���.X��X�¾�-ʦ���%Z�
��s��>�{�#?�15��>.��t4Y�[+B �M���c���12ba����1���n�-M0w�1�8[��ȱU�y�s6Y(��8c(јX�<2� ��0��� d�e2�2�4���#4��3��X�,��<x��(�8e��P�I�(c�H�xcC� `��!�!�PPQBAC1��x��21�g��P�`��c$e��c8�N8c8�4e�!�`���`�,c��,���2FS,g�X��i��b$�FH�!1�A�(c(�������s7=���z�d{���f�٫a)�Y�n�[��%�%��j7+3MT�elϽ��7��{=�'�}��ޏ7/]�eʱ���;}���Ƿ}ngk�vf���3~�7|6Sh^e�+'�{q߾��s�T�{��خ���I<�i���ݙ��~=�����}eESƞG��Խ�^q:�q�g�d�L�~�����~�j��ۣї��ty�1�Gg�f8�C�^��3~��׷G�Ȉ��n�-�I!�	ڿl����.����rI��~��߈�>�S�r�m��\DU�U�'u�_�=�OY��+v�K�8�۳�-�F�uy�%~�*�c��Un���ȧ�¸�N�����͙U�M'cu/=Sp�z� �Ѯ6}F����p��*��^�n�b��or�.��f���������?F�V��d����������m��������-��w;ww����ows�w{���,��8f����2FqG��8���>�� ͘BIOP��X�̯�$�;�@�?��Q<\Wc�g���ٕS�Wgb�K4Z��RD����E�UH�Or�CP���l�A��9G�4Y� ��L!�D!�Qk��D���F��ȱ����3i�o2�c����R*��WL;�F��̉f����Q��+,��ƞ���ϝz�Ӄ�H�(�3�W|zc�RS��� hIG�!Ĩ~����b�r"����!=G�'��Y����?5��נ�J�I,�镰�e�g�d:`@�^L������b�Q��	�J;BU�__���͉LOee��]Fg]�/�4}0�v>fm����a0�fc��~��ǭ8ӏ�?~0��!����8e������S�Q3�jt�#�˨�ȷF5X1̷S���Xu#5�R��ޏ�,�6&��jWj�;ZG���^�Rk�  !#��ِ��=��A=�9`[����T��Uk��xw$�UmMe�zrm�*�^���a�"�D��N��	����X������~�&t�M)�޹���g-��y=b2n8�2ܽ�����~ڣ�à�|�6��_��d��X��5o�����Nco���ѯ�!Z�G��w���C#/�t�䌉i���@�~�EP����(?Y�i�4�a�1d��c<q����i$�x���=CG�e�9��-��AN�e���p���ѿ��Ǒ�X+�0��d��kW�0���H�3�%U��zQ�����[5]�_$����A�_��&�$����q"�f]���$�X�J=F�|!����n4ٶ8a��v��J��a�e��fXS�mz�cQ�N���O��4�a�LC#8��X�,�KO�E�\�ER��{UTA>6}N��c/,k���,��~�����t��/�F��cm&��|�޻��������C�x���;!+ƨ~�u.�F�W�J���/)X6��d��r���T�lj����5���Ӭ�~-Y0לּ4ì�ه%�����ͮ�X����m�c�+ژq�ʞ2�1{���G�h����i���b�'�3<a�o|OoVĕ�	�+��S����~nם�չ޻��7�w� K�CA�/IvB�����ۿ�|�=�{ţ�vG � ������y��z�b?'���b�6Y*����&.l�������aa������:���"�0B��jy�ě?F|�fsk��l��ˈ˼���?<q��箾~zۏ�@�H�?1�q��-Ǫ�:a�!嫟+��H�8�X�yLU�bi��;�i�&�#c�H�RH�AU�S-du�I��m���̤@"���lN�=�*��Y%�Nh��  ���s����o4��g� L�-�l݌R���fk�Z�3�vq�'�b<H��xn���S��"�H�R��p�Ѣ��Q��S]�6�����Jr,~����}~������iQ]QcG3��th��h��	$���T���h��Tl7���|j��0��#���ɗ�$�E�����j�3��2��.�._z�uX�.���F�ٽR����	u^����"�8��Ɯa�2�,�g�:p��c�~�2H7�UF��G�O~�sq[/W-MuS������$d��Q�Q��)a�щ����d�ʄ����}�c��>�)�s��W��OTt��BX!��Y_�2�L!us.���Yf�9FW�,����~0M�x��""�����#<h#BH&��D�e���"$��?~4���1�t�ǎ�8x��,�E�I�U�{7;>��<??g�4o?�������ǜ]G��e�m��jO�{�O��	c_W�x�><T���^I7K���ܲKl�J4r�e��T 0�3����]T��LJO��;��g���`��o��˭�U��<a�EO~Ի���'tfn����i�xӆi���0dd�����8xᇫ$!�UTCu�>�2ӱY7wv��ϧ�n�E��~쯈~�;x���!��.�����J���+�_���\��ş1�96�}\�)�?Eo��m�2�����ڿ�ƣ���K[2~Sͫ���ڶ�G۷i��=L��I&�i��$�4f'�A�<3ĒQC C��`���0e�f3Fi���X3`�0fҲ�@�FA�q�8�8�H ��DP�!���0��1�4f`�����(((�����@�xC dc��<!�c0��3ǆ2�3�8��8ӌ0fњxf��3i&3
<H��f�1�c�H��0����"H1`���K�(c,g��[�_f8s좄��"���SEU@��;��*�m˲�������+�c�[ث��=��BǑg�i�o��2�.+_v�F�!�:����l�;aJ2k%A���;s��Nm�S
�#~7���#�SF��vL=l]�lr_d�d�֐ڔ�ͼy�X�ӻ�9rۙh��s\�n(񺤄�H�u�M<�R�:�����n�Ye{��w]h]do�>��'��P��%҉�K���\�)D\DR<dJ"���ǆ��Xh�����Ԏ\F�ʥO[�
�]������õD�r�c��WA��.�0���#�и��8��1��єl�%����iwǶQ��h�FɆ^�r81��Ȃ3KjWnv�[�Ï{մ�.��L�61�si�`�o���t�d��.&Ɓ(��k�5���ʜ�Ֆ��H�4:�\�;e��	��i�&>�ȅ99���ws�w{�����w{ww����oww�w{�����ws�w���0��8�N0��#$g��8x�+܌#�r�2����7��4���Z+T�� +���,&�;hL�Yf��[Z�&�#33k�@#�Nb�)pK\۬��HD�u����QItl�X��uV�F�FJ�Me�u����M�+xɄλv�M�3xڍ��M���T�6��bWX�9P�s.�ue�d%Y46.���-�.�jgYM�Z�������Lk�Y�q��G2��� Hklzue�8ߡ��k�Z�8c����H������[�g���,���y����~����z��s���b�q�����~�������l�ۑ����U��c��l�}8��Q�i��}H�G��'���J�r26��m�'���4�MJޢ�t2�a���n����p���f�:�NA���K%H5��o�o��UXJ!�$��h�&�?if�3N0f��I��q�x�gO/UO���=G�rH%�Ǿ�I6\�H.��ttmX�h?'�er��07UdR����6?��h�?}�4`���s�1Z��*eR�)Z�IX�|�Z��Gϵ2Uq�N���Z��-|�mRF�����I��Ad9�M�-A� �����e�q�ӌ� gş|x����K��ڪ�Q����Ú[+ev-|]~,�G�k��\�^�׬+�F��nF`s����l%�x8a���CuZH�MfkS��2~>����=BA�^k���˫,�J�;CI��vJ����y��V<^����YJeF�*�i|3��FO�v4Ҽym�ҝ�s�=��ﱂ�x��,�i���1�i&�iƜa�]��⪢T�3}�d��>6hN	�X�����L⋃9���w�\;:.lVV��>�l���X�Z����߇�h�@�J�?>Z�&N�Wϛ��[h��sE�TxL�V�� rR���������Fr��$���ӥ�&����Q��ǍI�
�,Na���?Y�8ӌ�&�iF�i�8gc ���-d��je�b������+������WZ#�[1 2��^ԅ���K�%�Z�<�\� �&%MZ�슄i[��0�MLB[�#���pL� %~����1���u�5�dn���}(eĐ�l����|�#�]��އ����E=^�}}ܷ1]�O
6��T�zA�	8�@d��BR�����$!�o�2��q��Z�V�WOf��K�Y|Qp|Y�5ѣ��	a����&�.�*����_QL�{��n}KQs#�!;�x'��d������`ʰX��[4�1���,�z�Ŝ1�q�0c$�M(�8Êj����#�2����&8���t�������3{����*�!Qugj�`���z-J��v����������mJޘqS�g��Ǒ����)��a{�id�wDg�,�%HO�W�]a��ݖA��0&c�[rK2���a�����MR~0 ��Y�v��w[� ~��~�tosE���&�[��~�ջn%i�^�g�ӌ�&�iF�q�q���U��0c�	6Xa9��]�cU��ũG�Ѕ�F��4����	H�~nvޮw?fVI1����o���1���bZ�8�eV�{U_ջs?1�~�|܈lO'?/��]�zS �#�˪���dзqn��	�-�B�pf�� ��dĆ�7adL����Uq����^���}��&���%v�j��3jY�4Qh�Sf\cu&y��]�G�G�~�`�v�Q6Q�z�n��BhN�vXԖ>�^�����:���^���>,��㇏<p	�EEE�j5�B��VIT�"�B��
�#T�@F��-S F�5�e�}��eS�9�ԫ7y�����'�s�-���v7Lr�	%^���Z���;%������,B���Q��{fc��ZQ��ʒI7F�E��j��ߚ}r�BZ����Xv�4&SG���u^?����,��F���8f�`��4�J4Î0�W|�y|�0�35�[�cYtxcЅ�����ǯ���@)�A1u ����MChUZ���3�t%��g� �wsFx�nľ��'哬xZͬD����0V�趬�ʭDFުRLCϔζ�W�W+�pt��W������S^^�.�{��G��o�Tȷ�t� ����{+nG�F�[^?�qΖ����>,Г2O{u��H'�;�$.�����?k�V&���a���gSP�7��2�~�/{8�9�*����84�em� ?�l�o��ׅ����]����>��J=fܪ�;}%���<��YƘqgf�`��4�J4Ï<r�iUi�3j4��|)��?vf{��a^Ev~_=��ܞ>S�3�,���T�ڴ֏�^�t�攳�W� �~I".=��]kX�4�c�:�-�n4�N+�R���.a�J�C�Y��	tp��O�{��	��I���Ɯ1[K�<H�2��(��!�1a#H�Qc,c0��3MfH���,f�am+<x�C�1�f�C4r�$��qx)8��+,��g��0��2
�Í4ҫF�8�¸ڙ c�3�B0c�H�4g����gq�8�fњxf���3i�3	<H�bc4�����&��	,C� ��Q�bd���2�Yc=x�?���֡#ː_xh�$�-�I�k!.�٤��z�o�\@-��W���*!�O\�q�KxH^�me�6q�s���Y(.a�*_�i�ѣEE�u�l���*s^�ʸ�9E��.n,��z��b���.�|�yY�ۻ��w{����{��ۻ����m���n�wwwy�������#Ŝq�3�3��&�|a��ǎ7b)�*�"r�&�����x�.>��e��vz��.f���OU��ݳ��8��%���MU���5�K"�QNX�a-N�u�����Y��3��9{e]�nO���Ϙσ�W� ���fj�v��X�/~Y~��TC�o���h���d�dP��A��$���8��`��4���<p�ݏ����ڪ�'+Փc�l�'*���?؛�����J:�)j���Ӎ�>��+9�%�?WHN,0DNT%����:C�=�s�If�~���7��&����aa���޻XpF��{tJ�u�߾��x��1��e^�7�G���(�N,�3�1�i&�i�a��F�$j�L@�fL�Q���K���ro�3b�1�S�����Ga�6W�-���@f]5�@,�Ik�TȆԩ�g~ _9rק���O,�C�d���~x��vg��HN�����M7K�f�gr�i�6L�A�z. �H1q�Qҍ��N�D�3�jH��~�5\?Cb|&�W�S�����٦����0���������^�
�m��Y>V�P�N������vK�,��T*��zO%�A�}B31��h����0��(��Y�gq�&�iF�<x��AҪ�&뤬,ݢ�Z�?�~W��媪�3�-k�K�Y��x[�is��)�U��5i��,V��M�eB���|'�*�O�E��?��ȝ��ZXb]��\��(�5Gbz0���t'��$BJ�<"B/�MU`�����KǕ�:��`��tt�	��0�K8c�`�I��Q�x����UZD��$��\�wwf��>'K�tl�	�U8���V���qq��~~e�m�c�陆�̬���Fb<8p5D�%��L�ڌ*�{��VZ}����k'H��(��!��z$,O��1�cO�����v=x���|��1�a�d��J4Î0�/'imĿoWx�p~�����7~�Md��6�{<e̮1�����ٿ���ҟ��E�Y=���\����q{����s�ѥ��6B	�:>��7�z 5mBK����TA�G�r�� �'�H���KN�C �˪�p��>n1�}��=G	BhN	���eǝ=u7&�0��ɗ�~��f��e�x�����N�~<Q�FX�1�a�d��J4Ï˫�=�N��8�C�i� T2g�sq��3O�Ϸ��6�^��{6�6�c9�T8����W�F٬.k	���U�O��[�֓_v�j��by���W��~����eJ��n���}k�ut�z���e���K�m���y4�q��mO���*�S��Y�*��t7C_��E�M��M�l��%y��6����W5cQ_��GCG�������g� ��=�*����'�Gq..۬>�'��<q��c-�e��|��8Ë�&�i�a�	|�I%iˡ������&�r�O-�|�k��o���n�j2�8m[f��?n�[hK!����ЏɆ�n�քD�.�%��)��wy�ˍ��D|l����QHBV^?�������z�}�g�J"#���� ��4��a�c8Ë�&�i�a�a���=�5fqUi舣g���ٕ�SU6pM��E��	��9.J�\�b���^}ǷZվN��f�+��Eꥭ����w�G.�ɫW-JUW˖f}w����c��q��B��uwJY�Tp��,��u��NQ�������ЇI��Q�X�4��gqc#$ҏ�<p�+n���U�q2_V�����xڽV��bn۾�ͫ���;��y�j�S'�������j���eF0��_�	�u���A5B|Y�,0DN�*��\�,φI�Hđ���D�T����|_��ᅉ�Wgj��Dއ���I�� D�\?���|YD�38��1X��#�C(D�2D0`�"�<1�����,c0e3M�h`��2����ǉ c�1���c�X��D0`�!�1�Bc�-�UӦ�WXWN�hѦ�Z�!�(C c$c�3Fh2D0`�!���2���X�`�7�gq�8��4њH��0f�6��$c�aC�1��K4����X� E��2�ee��fN;(�[�a2r�)�L��L���^�R�mZ��҄�k�����A�0���$6��ݦ�~��ޢ�[�Em&�͚G����YL��ʳz�g_W_�g]�z{�2XS�]cz:6�0b�gBRmuf�e��$��3�hs��WL�ɯN`.�!��ZA�0ws�h�,w��{_���k}YbprG$(������N���C`pTV[-u��n7��☝i��P���0�1�i��˙�0�v�6��_��߱�.�n7\�X��y���'�OX1���P�l��#Ou��\�.�y ׫�0x�ݪt����gL���3�"�է�Ui�kI`�]S��b�k�Xb�m��kP -�n��uP�ٛ]���SG�0ɶ�:�"��6��j�ɭ���b��Ȁ4�$�n�x"�e���*��۩������c�����T�(R8&O���p�>�f˫�b~�ǹ�������y��}������33/������y�����8��8ӎ0��,c$d�Q�<p�����ԐI�2�Dd��]�0����R��q��hJKu���u��uf�ݜGi��f=,<W��,� A���Jqn#6!3�g[]VF$�&�$!*]�&ղ�KZ��	�kRYa��[�;���t&��B�	�ũXe��;[��H2�\���R5��@;\\�k�\<@-�\����1�͒ɋ\�VY�!X����Rb#*tU�R
�R)bw\̈�&
0%��\�ƍ�F���[m���1�f�ְåX�π��:��-hN���--ՋVj3���������`��=s;D[S�tj�n,�'��q�*R��[ysTl�lK;I����ن��S��$��lL�j�n�����h��_��c�I%�Y�8$g��P����QgЯ��n�⎒�8��dp����%�e�ffs�x9U�7\F��Q$��H0���ь�<p�'�>z�]k��ݶ�*�G�]6����RBD1j^KP�����"�Ke˻�`ޒ��U���ψj��abn���.Qr�p�|?��U�B�_�n��'#QH ��|��P˿��4|gt#$��n�e�V��eX0ۖ���v|�1^��ǋ4g1�aǎ#$ҍ0gq�U�N�L�R6�h�L�>n�W#Êʻ2�-+�c��w��z}FϑГ:��Y^r�ݴ������&�0�.�C�}��ea�xM@�t�dE0!�ޤ��6"~/��ㆇ(M�~9�Y���{=r5Nuq�,i�va�u����3��h�q�8d����<p���$�%�ي�H�O|�Z�Q�ǌ���Y��Օw�3��6gr�.�[,���V�9Gv�Q�V	�R�M?f���~�n�����~[�����Mm����~0����WGF��s�ń��4CBv�0ZL��v7r��т~k��I]?<ɵ6�<ϝ���箾uf�3��Ë8d��M<`�8�b ��EVp��
S*t��!�+nl8�b_�������x�).v�k,���of��kρ� ��*��ؼ ��c��[��v���n,gUe�,�L�wV��K�E�m��כ&����>�գȭ��Ѿ_+��%*t��l�؛�����l9z�hʾqYqz��p� �xw	"Y�zt~��p����	�{��.�if��WTX�������%���,��IvJv��Y�è��*�c0d�e�fc8Ӌ8d��M<`�8ᮧӑ\�{�:\բ)6c�3���[٪��5cMgZ� T�U���<]X��un���,�p��J�6lHkݗ�B�.l�kA�_��z�m�=[�Y��b$a�q�B�D�"tp⡵D�yGՕ\��>��U��0ؙ+�{�1��#j�y����ۯ\0f�ь�N<p�&�x��q��j�H��*�>�������pL���H`��`��ƍ��؍b'�>���A3%��NRB6r�,O��Q?������^/~��BJ�<<J���)e-�Q�4%���HA2��>��l/�n����+Q�����T�T�a�WD�X䯧[z��^�q��8��[uŝ,���æ�<|�AmUi���٦�M6�ǲ~�i��j����n@Lp�.]��3���>4~�e�����-=V��a�c,�}�Ͷ+{����ah�"TLi?$QŇ�H�=J��qth�!�3R��Y��h�pK����BW���a�f�,fc4c8ӏ2FI��0e�<p_$n�O	l���!m���➹S��Z�0���5|*t�"�q��h��AqZŉ�]e�����(��蝩.�qKV��ԡ1aL@�O| !������~�\SV����BE����#����as�%?a��lS�7�qd�,���( �>���C�k�n�o~��ŉ�9VY\�zE�{�Q�^�|$0�X�f��\}źiU�߽nj1:��Y����lL����_�ꍈ��B� n&*��3��J�7��+�q��s/��۱�����κ��u��.2��o\x�Ϊ��m�NԢQ�te�&���|<d$��u���ͯ4ۊ�n�<�mǎ�#�t%��Ҏ���`�m8Y�������E����Kd
Յzє�.\�Ԭ����6X�8w�Jg6*�E'h��9��U�؟Xz��[�-����m�z馣_�=e�o���0��xg�P2�P�#<Ib,��P� e�f�F3Fxf�I`�C0e��Fad�(��d$�3��xd2D012`�x����(�e�q�p�[6m�V��x��}�P�@�H�1�f��d�`��C#$c<1�X�3Op�8�8fa4њH���3i����H�!�3Ɩ1���<1�@��1`�$��C<H�Q�,d�TdW���mm�I��e��}�ث�}?�){��N�gީU*��s�~�o����h�5�­�;���ܛ�S�4�U�G�Zw��y�����www[��̾����������������̾��Ŝq���4��I�Ϗ�:l��W�Ui>"��
���$�AcG�l�"z�ߖ�a��~^Н�G����RG2�a��osZ֌�pO�|4n�� �8��d�Ɉ��.<eߥ��X�[f|��;���t�E�`���\0��i�~4c0�q�$d�i�Fl���Q�U�M�e{(ѣbX�8oee:��������΁�����~�M~�˜�ǭ+�X��a�;��G�?tB�9Z,NX��N��o�_���m�	�7]0���Y^+O�35��a⚏���e�h�1�q�q#$�O2�8��h�5�D���� F�K	Rю�E��f��-�ډmi=�^�<⎪K5a��n+����F^͖٢�0���늫H��s�L5ɦ9վɷ�{�/c�>�쉡����wM�6�x'��V�U�>�mg^��#�a͝�o>�_rIG��؉�6hQq[ �%8��i^�{-;-q��ڳ���F�	�.��uZ%wz]	��g��?Q�2�r�٢��>���o.`�����7^�#�>�T7	�7���E8��4�F1�Î(�&�xіq��@��S*|�I|�g�U�Fhh捣�'���d�lN4&+��ÕO}��f�Y$��A���w[TѣBk�[������*�.�~��:F�jIj���-�Xz�SK��q�NҗU���ن�|׫^�7Xs����f�w ������6#��A�>�����<31�f�(�&�xіq�y�x�3J�H��QTw_�C7J~0��Λ+��C*�Cf�!�Y�%ؖ'��	MM�)vHZJnznѼ�fal�]A5��t��u#?���!d�1����J?Q�hDآ=��TM�LT(�,D��i|{�0�i�8c4Î(�&�xіq�'}+��%��y�G���U�U���\���(�UZD��g؛�؝2�����V	�Z-2e�eʅ������y2^�W�P����<��Q�6pG�+f�{$�f6#Hv��Fr�+*�U�ǵV��ב�a����{ؖ7r��O#&������mz�ś|�ΰ���_=u��pf�q�q#$�O2�;�+�J!)�|Q;������a\[-�?m�SBz���Jඬ0�~}���^�NN�Z�%�"*�4
eo)g���2���� -���q��!KɼU	U���g]��io�+FR�7#�}\����t�;��������^���_��Z�$���G�}��O��_�v�1�z:z��	t��ʛ��`��-��a��Y��"lM+�a�P�������Uz���E�D�,>���a��p��܍������A�*�K�5>(�Dcl~L��ljB'�k�����޶�+��r:���_N7��G'I8��h�p�3L8�8��4���M�<z�mUhk��mr��z\.�ؤ2�����=�Y��8_
�n�b�g�Z�T��U9)w��wa�2�D/�gFxj��%���y���]e}N��9}>�cL��>��lt�� ~���6{�fh�ц|/��2�8����qGIĚi�FY�t.��U��ޣa
>0ʤ�7�%ː+��WQ'�����V��A+X���V��CI�z},�U��s�t��M�|����-�ӗ��~7Bh���1�M�<d�{/��r��n1���q����1�nN>��LƘ
8��RH���<3M8ьf�~8��$�M4�,�'�ED����gV���GF���o��K!�h�i��h-��B�zMО����X��79�˵p���Tz��cO���s=��ۗJ|��O��2��(�ʩZ7V~��Pϙ(�Tr��Q��d/*�\��,�B� ;�0����T�a!NH�HI$�Eh��y��	�L���b�?9��ňfa��BFԈ��ciw��k�E�V�]7��U�-R�B)J������)aK�))K%)K%*RȥJ}�`�XRT���%(��(���R���)QK�JU,��X��Y)T�J��)K���JQb�
,��*��)KY)T�J����b�E)d�)b��b�KJR�)J���J�-)E�T��R�)�(����-)E�K��,QJT�R�U%��)K%)K%)K)JYIR��,��,�JYJ������R�J��JR�JR�Id��R��J���d��UJ�TU��V*��T����*�b�*�T�%T����d�*�R�UUQQUaU*ȪU�U*¬��1Ra*ȫ%R�*�Ud�
�QJ�U*�QV*���U���d�U��U��UR���R��R��EY*�aIUeR�UUEUX�TYT�%UX��%T�*�E���UV*�ET�U*��UX��Ud�����R������UV*��R�UU��I�X��Ud���UQb�U*�,�*�Ib��R�R�*�X��Y*�R�R�R�U*,*�XUU���T���TY*��T�%UUXUU���d�U��X�UEIb��UaT�%T�*�T�
�V*����TUX�U��X�U��U���0��%UX�U���U*,UU���Y*��R�TR�U*�T��J��QeUUY*�b�UVJ�E��U��R��J�VeE*�R��*�d��Ub��YU*�T�UJ�UQJ��U��UXU*�ʊUR�T����������UJ�U*�U)��Y�)V*�d�dU��X��V*�X��eRU��U���Y*�XUU��*¬UJ�QVUJ���dU�T�*�T�%Yb��EX��VJ��UEY*�Y*�Y**U���*©T�
��TY*�d�*�QVJ�X�
�U��U�R�UU�T�%EU�R��U*�UVUS*�
�UJ���aVR��R��TU���UEX�*�U*,*�aVR��dU����*�UV*�aVJ�Y*�UJ�T�J�U���R��VJ�Y*�XUJ�U�UE�-,T�RX�`�RK�����%�%�U�b*%RK���%���B��,Q*�X�%)%���%��U!b��P�}��Ib��H��,X�S{����`eF�0U,R�d���4b)T�J��U,R�YJ�b)JYJR�E��,Q��f)T�RX��X����KX�)d�)d�)aL(KX�R�QJR�aJ��U,R����JX�F"�K%*�JU,��U,���3�JR�*�YJX�F�R��)K%*�K%��&3�4f�))T�R�b�JRŌTaK�,R��JR�)Kr�b�K%*�R�*�JU2�����K�Y)JYJ�,��YJR�R�R�d��,��Y)JY)JR�)R��*R�X��U,QT�IE,��)T��R�*����*R�*�R��J����)T�JR�*RR�*�ڌE)K��F�K�X����U,R�JX�R�U,RU,�R�J�U,R�,�Qb�K)T�J�),�JX�)T��JXR�,RX��J���JXR��)E*��JR�(��T��T���)*R�(��QJR�*�)R��Y)JX��J���)JK�*�JU,R�,R��,E)d�)T�R��J���),R��,�)b���R�JJ���K%��R�)d��E�����K�,P���b�K�X�����T�&
Qb�IiJ,��TR��H����R�)R�%��X���K����JQb������R��JR����,R�,RU,QT�������)K�K�YJR�,��B��JR�*�(�X��,��������b���U,���JR�)(���K"���Y)JXR�Id�����R�)JY)JK�,��Y)T�K%,R�IT�R�d�R�*R�)K���J���K��R�)Ib�)d�)d�R�,��,����R�)T�R����R��R�JU,��,�Y)JY)*R�*R�*R�*R�,)d��,��,���)d�JX�E%�T��T��K(��R������,�JY)*�)T��)e)K)JTRU,R�b�K)T�R�e"�X�R�*�R�b�J(�J���,R�E%JU,��K%)J)R�)aIb�)b��,�)d��,�)e)K)JYJ��KYE��XR�b���R�T�R�E,R�d����b�K�Y)T�JR�%S8�*R�*�R�e,R�,R�e)K�X�)b�H�YJ��U,�R�U,��YJ��U,R�d�RYJ���X�R�U(�P�E��,��YJ)b��b���U,�)b�)e%)b�E��,R�e(��J���,R�e)K�IT�J����R��)QK�)e))b��R��R����K
T��(��,�T��J�ء`�E���f��ɭ��^��4&�q�( HH��F�,`�uRVě~�����e��>?��L\O� ������8����B��C��� B�uޅ }�|SSYG�]ָ&�����<��J(s>į���R�ؔ;�s��`hlQ�����W�>y�>Vܡ�" � d�sE}�PH@�B#�>�x��\x��C�0�%RAJ_'�l�At�gA�|X��6�:OZ��@j|�%�t!	A�1V�ׅ���-��]�����Nt�O��II�LO���5͆�!��"ySr��������!?�/a�������R@%j�r& F�D�&e���3P��XLԐ�PtET/��+�EQF0J�S`���;�.�ע�l�ZXt�� O�b�I�RH��H��D��& ���(U����X���\�9��w�Z%z\�9��]N�4A�b�p0(����y�|�����/�
"�(�:��E��ob�#�L_H��zN�1 �}�jbd�� 9���Q����L��/�����xV�;�i�<�'�p�E�tEH�}���W���ffbf>��w�T�6���TF��AQ�����"�Bw�y�'d�Z�s���y��pܮyB`���0�(A@�ѮB�$�lI,�X:	g@�(*4��`<X�l�xN X`b9��a��1?�R/�GĽpi���Ł�8�zX�d�K�d'�rUQ�τ�I�w� ��*�qAQ��0G�AX����ڄ9C�=Pg������d�X�;�yj	�=���ǀt�=�0y�ב,��(~O�~���QE� kQ<b@��.�J�h"�8���9�9���È�a�6��nSX��r{��2~@$�E#C��a����₄.�z��w!rA:z��bi�`̸��%���P����m�����������.����9�q���<V�/b��a������Z9I9�HQ���)@ߙ h}���f�� ��?�1O+g��LL���ш⛝fb" ��r�OU.>LJ��8�~]�=	#PP�t5�c�����)�0��