BZh91AY&SY��ܨ�i_�`q���b� ?���bG��   �u�[T��ZKi�*%�F��S[Z�H0�BA[�6j�T����UJ"֊ kDUm�4cZ���T�h�
��	��V��N�m(�jRf����CE��6A	S6$H�a�Ъ�l������ژQ������6���SSj���U�0VT+CZ�4�`��-6F�5V�v	vҶ�e����UPR1���V�%�1�$�-)[-j���֡Y++j�4ɛ5��MY5UMdm��5[m�!m6�Vն��̶�uRSSd�n   ���[�io���R���itt�ڳu��{��OF���ZMҰv��\bm@ƫ[���dU��Y��u�w�/ct7m7���m*��ԍ���6�J��   w�T�=0�{˞��K֊���<*����{�*�m*�ޏx�-n�W�^�N��YJ����DEk-��}��UOl�}Ϗ��R����|�|��m)��W�}�&�$����F�(�p   On��RT�ý��������}�|�*��w���ʡJ�|>x���
U=�>璩T�־���j(J�3����ҕ�}�h}������ϩ�>���R�^��M ���ղf�   ���ꊯm{���}}R�**|�}��R����U�zK�n�!n/��ȥS��Q�xO����W�}�
}���*�R�����|�/CJ�}�u�)V���T%Vڍh��6�5Z�a�   ����*
��[oy*�Jgw���/�_p^�P�����ʧ�	)��Wz��5"3�����_[�n�W��:zҚgm�対}T�*����aR���[lf,%�4Y�lkUm�f�P  �宅�����x����+�{}�ʾ�JR��sʔ*K�hp��"��wt:�)�^׽��J�Y���OMQ%+���z�wJ��Y��S����·T^2������ڃU>   1������y)EV��==�T�(F���҂�*���^ڒ.����jJ�S����kJ��Gp7.�ƞƊ�<��U:i�z^�y{i���[ڦ����U���V�|   ,��AB���ޔ5��
�
=�0 �W{�V���)ΒEG{�=��@�r�xڰ��Y�@wQ�T ��V��m�ƕ�P��lKBɾ   �ޮ��
��D�w���T�p��]�^9��v�'s�<UW�V�5s���u���t�k� �Iy��{�z�5��[� i�i�_(  ��	�S�����n�M]�^�5�Ҫ��ծ�
Q��C�Ps��+E^;���Ҭ�7%�]��s��|     �����J�&&`i�&#��ъR��hmF&�hi�aCA�~FBR�P�h��  ��B)� ���z5      ��L����  @ e)$���ڙ���CLM?�_������5��O��o7�������*�j����=޾|Og����y���m�m�����lm�ll`���clm�~�M�m�����z�'���q�������`�����;�����`�o����Y���L�1��6�?������c��b8�m6�m��hC&�mmD6�cBC��6��&4;m6��BhLd@q���Bm��hM�;m&�mƄ�C�`�C���L�ƄƄƇm��v�	��`!�hp#���Cb6!�Gm�퍂�؇m����!�Cm	��� C������`!���l�l&4 m�����m��`�m���l�� "`�C�`!!0!�l80&8�1lm��� c#�BcC�m� C� C��hC��hM�;�;�hChq�&��m	��C�І��a�!B`�	�m	�6� C�,�޽z��x�?���_��w���g��>�<&^]���.Mgc�Cˆ�� ��u�UhR�ϱ��Z�|a��n����͙�ͩ��G�wV\z>�v/�J��V'{�%ѱ�BSN@�q�x�8���L`$�n��z�]�mjyy��YU,7RP���	����p,q�z6�?^ٰ�t7o��oiQ�5_5Vk{p�kcu��jݡ�[M	��ˠ`xE�Ze�eh���\;JԱ����+���Y�T���VA���,��eTh\�I[&V��V!$R�j1`���Ŋ�y+�`��9TX��ݡ���VH]1�0��y�N�H�*�Z��id���=kw��#��`�=��!���f����B��3J%��:����ˤA�@*ɲ�:h2�wiKh�˙l���`b�mZH�q=�6K��~̠D�!̤���$9`��R��l,8%���r`���^ʦ�*�姀[�;��YA��^��/K4b�hY�0^�ԃ�0�+�P�ź/�:_Z,�4sP�Xj��+��pS�7�3�M��i�n�`')�I�sUx�^6����XX��±iW�~�Ld�ۖa��cxr֖�f&�t]İݿ������(G[�S�m-xfkE��_YŃ6��TU�-�n]e�uu*:G+P�!��+�L@�϶I��@�fF�I/EejYi-|�]��F�u۴Ѓf�B�Z-��ۗi:ߛ���6A{�7��T����)�xM���]e�� |�㎹�ƯU��37I�a��
��י�M����X�V��"F�<~��ua[����.���Mp8�M����v�x��V�4����^=���K�n-k��RF⚜J8F+B�r���X����CEb$6�9y�bwXk.b���%�[��U7����f�2��
�۵(�.
X3J��rC�ݸI�b�w��;-��j�x@�E!K0��d�X5K� ��w����h1��RR�l���c���Ѥ^h�,Ux)��ҝ��mc�2
�ѻ_��7�S�B�Ev,�c����$ggom\�(I W4�Ö����*V��l�̑b�ň����1�w\�����T5��k]�w(7�R�MH�)�e�#f�r5c���W����jN(��.��n���]���
���bڗO���$���kU�Ϟ�6�m�E5de�X	m�ͤƠ�L���9�[���T5Mς�`͸��rʳq}7�o@��2k�n����CN:.�����9���:�KŚ�m���o�C��B�"���k�̓��	X9������֍�n�mf��2��Bl���t�^'��vh 
V�d���\Y"
S�7�Y������8��J�f;(�ͻZ�2�`.l�{m���b��Z�ȫ(��ȣ�M�c��Mû��kuۆS����?eT��E�F�r��ɱۭ���)T�N�3#Z-��c���(�A�ǧ��P���7E�[�+)D��v���NL6�j��<ǯ!��e���l5���d�@��f�e3D�ZѺ2ȱQx��y���l">�uhv�����P8��FJ7n�Hu�b��k(��!�m���T"�z1��R%0"j�"�y��=���]��	�'�wb���QT�\������7a����"�b�TcI�͚�eP�P�G�=���ʇ5�2
w�r�v�Pݹn�A�o(��U��bULDp��V2{�q|���������6��w�C���aW
��s&�z��=���
�,��7Cy�:�9�ͨ���sj<�۱{��e��`?'�R��p����9��h%o�iR�}�L45��GL3^��Ė��� �����n�Y-� Uš�zD �M�{GKQ�D2�&��5��n-Z�T�U���+.b��/�KiHS�jZQ߱�u,�&M�Y��*�)6�%H!Ql�B��)��VZ;
kv�04����j^3,�����\��N^�!�d9n�������f
�7���m6�`��@c0�on��;����2��/��-[�-}��q�Ԕkh�݄�kpi�r�f%�$�UҏZ��Ե�f�7�Zpk��y3E��P�n7��<�����gպ�}��k	��崏`^�n��]1Ϯ�e����q�D�kp��)�|�����+8���E�tA�K7K�l��z���`v�\�a	��A:&�;J���p�R�`���Ȇ����Ѭ��mnb  �h@7J�$(�QK���d��씯n��4��n�-��R�$�W�]5c�t��]Â�lQTN����nB��,ʳT7p�sd57X;B�JnՆ�d���mѪ���H�2&Ѳ��B�5=5ͤ���8�8	��6�����qA�Ev+%0�,S��B��d�e�n�)�CikYV����T��ᬬ��� ͼm+[AD�i�c�4?�敀]�'5.�k�ZB 2:Ȕd��L�5E[T�V��JJ\sU�@�����&���곢eY���;����޸j�wV���!w��팅'�!��"ir�Ͳ��R���f���<YKv�(��M��*�L�,�sT,�b�ڛc)c�4�Ģ��:o6�(1"O�.�kw�j+�����/�)��"2;��4*�Yd����Еz�J̈��^m`b��/Su�L�U�W����|q�J����Q|ܳ���J,�ɴ�M0c�Kf�[�V�T)gt`��Lm
��ٶw`�6��;���0�T�+ZeԆ�d ��7�q7�c9�n�������V	�yp��U�ԛi���F"&�O2lH,�Z��:�;c"�X�Jj�.�3v���i�geMZ��ݪye!q��m5�nl\̬ǋu�{ug,���%��\v^-kS�P�k��pT���d�A�Wv+���Gh��2�8̍16ѳ%�otx��4�޼�*V񵸁\�,��,ޥ�,�c�{*L���a�?X�,�e�U㡱	&�%�Z 8�G�u�b����aSZ�&a����r���W���џGI�E*�w+]M�rv�$��ʧ����v`ŏZI�ً`c	�S!5�;��G�|�v��(����{g[z��DR{��NXǠKgm]�U4�!��e����f-��	���w��]*��v�&��֭���ٛv����|6Ҽ�-X9�d=yh�p�(r�a��U�Wl51n링HCZmA��f����4-mdG[�>)L�ӗJM�b�p^$Ԍ��77q���nV�`��,����\Q켅ۻ�5H���޼�v���L9`)j�lj�V�w��3*�94�ǳ1����@���y�
3/ L��&��&ģ��2+�D�M���ݕ�BI#S�k�h6�hs2蓒�e�-��mL��3n�E���b��j;��7�V��ҹ�q��{z�8n�[#��k���6�-A��f#O",`2��i�hT�MG|u�.��V%X�����wNs���ڰ�(41����^V-fևq�E����0��Qjy7r���FxZй�\�(b<����g;�m�,����
�5n�w��ޔۤ�sn���H&Hy���`�l���m]Gh;t2�C/-�ķq�yz�r��yR��Ń(y)���8S�-���`ϰ�����*4م��*�^f��Ho��,'�(2\{Z2��v��� g3�{Y4\$.�y{7n��dF-��A��4���0!L�0�b#q,д��[�Z�KcT.��0��V���1����sEH0ӼTsc�F80Et�՝�LEn��2�z����Nn��fjJ�\��R�#)�z��,ֱ�Ҫ�^�:�y��3tLPF,�oq-"��ƅ�𴁚潻c,Zq��О<�	CM����XKd7B�����j[�ee��7"��nf|ͻƂ^k��q^L��䱂�ڞ�!��Y�q�wf�J�):U��w�Xt/N�F�9oN�qv���5���rU�{`66�����	����d�8;�*����Q<�mY��_$6k�h7�]�YF�eȣ)��N!�n�x�Lj��jkK)�w�O��$�d�Ů�*�l{R��n-���([O��l9mBs1�[%j�F`�����^�-�F	�	ĖW6ȰK�p*�Of��D�b�j�Z�����9qb�(\x%�h�pd�e��o�˅B��i�ܵ�"(\�-ȥG�Y��dU�����0l��{���s#�0�����Y��l�j
8�e�nbX�7���6!��[�Vܒ��䄱`�e#Ƃ
kj�[Wq�n�aM�
#'��h_�MW��J��U��
�]���'����.h�U�n���s!���Ѥ��kcx2� �3�p�JR Ӕ�A,8
Wgu��M�U]���Q�Y)'���6]2����R*:o�l�a_8�ݩ&Vjv���JPx��em�)1��@��fѐ��}��H�c��di�_�!Z�D9��`[�>���ŇK%޺����虸;Vz��k��X�i�q�8�_P��N�駱��vZ�9**��ބ6�Oa'p�Uci���%uP���lB��2n&ӓw��kH�܋LM��gj�є=�-��]ne6�&d�n�A֭��[� �33�N�3��a[�䄔&���b\wL��j�%3�X@��M���̪�֕�S��m��3V�09� �M�RҮ��ӻMZ�b�%�"�W����]�5�v:����1�C��@�MP{�d�_v䘓R���!��ù"�B�mS)fIcX�v�A�7H�zff&���U�!uw��:Mp�U��l-���B�w�;����^��Y�L�X��^�FF�:$d��y.���iLo�]L�AK�U���m��pD2���K;����T���|���[zI�������0']�f$>9�jkvJ
S��d՘2��`��7x�����L�j�ɲ��gϢ� �oN�bۃ�qha�n�X���!��d��^����Z�s�	u��#X`�bZ&�� �Hu�<j�Z0-�olX/w@�TRQW��Q4�Om}��b���R���e�dT�̘Q�� ��[m|]����e��Z��q�g�X�O�� L�'hm�%�kn�i����m�S5��`ʴ�`�Φ嘃+�[z��4��ח�JA���jnb��ޭYdڛ�lC��6��T.�yj�����Z�ձ�-7\U���;b��B��ڃQmb�G&�z���͗��hF
M�%͘柝�!������{&�%ꦢ�f�e�RU�V�ˑ'A}mꁌ�C���1k����FP&�7j\�t�`�ͩ�^0]�N�Y����2��͢q��Ֆ�X��ר"45��A���M;����H�*D!/ Sy�,���;6N,.�庸�����^]k�V��41����i�[�`��f;q ڐ�q�ϐޕ!b���;t[��Ҩe�]3�K��U��^��@'���e@���(�����m�����w\[b�6]5����32����E�`�+`�L�����՝$�L��bֈ�[ͽQcNd��Ǒ��N�,�ѷY@Qn��45�{r�A�4v��2���u�����K(�p*���qݸ��u&vrM�e��̟L��ޭ��V�ǁ;�!��ǡ3�����u(7m
�Tc2���*h� L�]���B�4�v��2+۲N�n��Z�tB�o훒�u��\�X^�;Gª�L�C��]�hu(7bS����c�^6����zr��3U��&����s.��#sfm�ʰeڴn�T�xe'd�[�"f�f�����0����n��u)��Ŗ�S��1l�X/�i�Y��+b���k�3^��`��t$���I�Y��/��x�]:����wXf���9s%�lG0dӯ$	@�`ڙz��ֆ �d-��i�Kj�$^�R�Ū��3��N�Bkshn��[��x���Y����V�=�V��@	wZ&f��Qlz$�K�V[�6��b0�4�cp�ڂf�1�d��hd+n��fa���h��x�Z��&J��t���)f.�P|]a�w���(RO@�y/�EY߹&Tq���ٸPR�R�or	�p�ƞ��t$�q�w{j[[M	5�Z��[�3�ZX��q҃Ly�u�70�71��1�cwv���w��kLRQ'Çb����Q,kDǆ�f��/j����Lm�I�av�ػD��j{-�x�*�Œf�t`��Vj��{q9����yK���b�U�m�%��+McXڰS@+,Ǥ�wl©cv�E�����y�a�a8(�����CN��ὄ]�Z���
��Li�In����F�(-t&�F;����D^���Е�p�ܵ���BUc�q
�L�Z��u�C�W��I[݂f�q������Z��b�;��t��(LߒLnZ)����܋V[���1
�4���ì�B�8.ֲ��V�2'����YXFbM���w�3sF^=�0���YϲU�k�Y���*:���`��櫳2��d�P�kU�Ә�ؼư�GZ�ǌ˘�k����```�Z�J��S`��	���X�6�w�x�?�N��d�&ֽsl�,C�!��uUe�YZϵL�긬h�{t�>Xʫ�!ӗ`
v��U�]Ţ��K�z��=� �7x�:��F-�MM����Kr-ۼn��+Ge��RA2��li��+K�><�Shn�7B�Ba��P���sL�i��GN]I����n^����r	,-x�'&�{�y�n*�৐ZQ�Ϭ*y�-�oR�R~��}V�c�M1��@�u��DC�n��k��'H!�Yke�c���P��'L��ʋr���~[�懵sR�R-��˯%N�f����^~f�4�N�Tf��_bʠ�ӧ��oo9űB�E��$�U��Ec����@�ڕ,l	��~����������߾���=�����;�t��b*rYʏ�±�}L��M�D�8��NKs��0�����F�-�Y4����-�Tsw����AI�uY��NҼ�ù��yJ˩��\B�����Jbcel��^����d��):�b�`�(qP����i��eN��Y��SjR`32�CC,����d�J�4^+z�I�y�8h�8N�w�R�,޲�����W�_q#��R�9\P�ᏹ�9ԥ]�܊94��W|��(T�|��j�]�}R�Z7�B2u�m����ǥp3��������t8ܼk`�jV$wM�ٗc�Ix���)?�l��Q#�]�*VD���VWufM�ܮ?�����glεD����8dT�:�tJ���tb�T�� #ǀ��t���J�[j��Jº���<��}�u�{{�1�ř�n����!�yz�Vv��3ot�&j�#n���[z��"�ˎ���K2#��j!&�ܙ�(�s�x�$��gb��@�����-�֡X�3wzf�1�R���^��d�<����o�D�[]��1�ݻي<ц��j]}f�c�F*�l��j��;�t3��loh�$�@�5�+�͝�(S��'a,T���P7={�Z�}�6�ޠF|މ���þ40�/wj���J�4b�4J����rރs���J���G�J�\��(/�V�����r�)$NlA7�}C���h0o`	�W>�c7��֦��4�9�����b.���0�P�<Ry*Ĺ1�;�K���[�4�:��o�tn��kx�����Z�഻�;e���叢�3.'Yor��1��f�y�q�95F\���	5"ԙ��|Uc��˽��$wuѬ{9B��97���yr�����ȧJ�c-_u}u<�p��V��b윛�:]w�K���F�<�a��nXJ�T��\��4X,���~ň��*�T����T(3��f�.�&.�Ӝ֗�q�zX/w+8u�]\F�D�NB����)(sނ���g\��o����.�ƅ#C�g-��h'�;����ot�r����@��W+
��"�������3a�R�9s+Z�R��Ă�q_4t\�È�U��B�5�'f�����@�W*�$ʾ�۫��Z��+�x(Z�/	wǌM���큈7MMO�6��n^Õ'�~��,�S=w�|)��W�\[ɝ*��,��F��(��4��ԍ��^�=;�Q1gE|+��%l��GK6�顥{�W~5|L�g���I[�t�-�\k�hYb���R֮8�x�T�Kp�w��8��W�]oihr�T1�;;�U��ܚ%��-h��W���̤��;�Yg�N���&/j"�i��"��;�*�p��a^8niV �sJ��5�yk��*F�0|��שXqnj�]Si�EG/�=cN1tX;�'�.^t�/�]t�Xt5��1�g�X��>
� e���.	�YZ�C���&kF�L���Z�X�T`Q9�9*���E��ty҅����Me�̎����W`���g�3���{�� ���HW���i��X�>P�e�R
��5Y|��;�X��8���]�&릶���y���V��xrg7�
�kkp9��h�О橖���薄7�p��p��yB���JӀ���	��-�d�J�}���o������;�aY�f+@�W7���Y�pz^�<e���yS���\��%�}Pt1��ް�>gn���k0�lG�B�k�Fr�6���' ��Ǫ�����AϑŒ�5Wm\�TQ�JRI�Y��tM˥�G=�2��2
un�Ű��5Yo (<F��z���ɧ��Kv��S�v�������H=�[#�v�65L۬��-S$����\�%�
Sw�i�b`�{,�+���C�&%e�#�3��u_d��T���9���u��ZHu[j�;������L����;@@9��G:o
��p�嵹��Y������X���U�y�u<�n7*�ܜ��Θ�엃�h�'�BM�s�a����+�������ʂ[�N���Tᦡk6�.=:��-Q��A��܍�"�=s9�٬a���8�YvJ}Q��s�����gTڹ��Ꝕ�����(�g[<5���漎bwҏԕb�2�w���ѼY�ǽB�2�f$3�尝�sbJ�ݳ��o� �J1e�ˮ*�{6J=zV�j�U�]�3���U��Ѷ�<�f�y8���5gix*a�y�pt�'{m�t(���a
D7�mc�S̺��z��
�#���-ޑ��۟p����cNb;]L�u���l�ӳ�ڕւ��a�8����+y�ɲ��9�ӭ��5�2\ڛ�l°�ɦ!�]{�C��ќ�2Y�@�sq�*��WF@V�sM�AY��U�K��b�N}��1���h��m��k��wV�)sj���ĸ5)�0�ܴ�W>��H�Od�P�y[�`���sP�Ղ�)�z���MZ���q,�{��.|詷����|�g@gb:�Kf���N-1C�S�nqS�0�B�Ԣ������ݩ
�PSv��ţ�F��AY�����+r�ʸk�U��59Х��9t���i��N�����+^s�ʓ�P^V��wxil���t�M�R�0_iyܾ;�U��ܝ9	��U.�ڳ4\�ӍuR@��q5���y�*�Ώ�y��AJN/�G��v�Y�uP��'٣L��c�.��rʛ����A�V�)�ƺ��h�5��|u�K�V^����b�X��A���W5��ogl����K+���N���5����dr�]4��q���L�a�1
]\�*���b:$ڗs�6���xp�lD�oRMҌ��F]`� S�5ar�8���Ms�GM�� �N�<�c8�As�cU�9�ǖ��Z�ܒ�B���jL�\oM��t@�)�'fj�VA��q��n]hoy_q�]ho�.�VLz3�����PB��9�L�]��#Z�o��*h�p�`O��EH�f��XiHw�Mp�Χ�/~�����1�v�=F��Ϯ��̩*���7f��3���`c\�W�e�J��f��3�;���+��{8.���u*�铩��S:=0�u�0�`�Y�7/2aKH�vr�̩��rz��}Z��C��{Xi�W�o��$��YE	��=0�'e*�v�]�����EU��+Ff����U��3�U��kJVNc&,}b��F:�}s�ӬV$��KV-v|�]��jP�	\�f��0���P.�$��ų��h,6/VQ)�Ji�3���䐆L�Ϩ� ��ғ:��/u��J� z�fe�^�m���*VbU�܋c:�K��Uluļ�.:�@ke,��2PƖk�h�X�ݮ��tOhP uāV���4�.�a]�]���R��Q���<�K7pcwE���(iT��N�rM�x�u)Qa.��:�Du����n�A��7ZI�=�2Nݴ�7I\�"')�����ޜ5�6�z���є�����T_"e�ɹ����u�V�q㎛�%��n<���U�k��'i��.���TGp����4j㝣֘�v: ��8�*��|�U��b�����*��+�Q�r��m���V�$a���,0���\�;ݬ�^�":,%�s�r����8�
ۨ�ŦvL�gH5�����:g9�2�f�-h5ّ9;n�T���hMx�-c���)�E�V����lݼ]4q�(�h�х+���ꮝ�J��Ʒ�&.��8���"rc�4z]� ����.��T׻Թr��z�Z��A�L<80�&u�o�U��4.�,�.�� ʤ��l�Ykީ+��wR�X=��τ:Hg�}WA�e�=TQ�u�	7y|v�b�Y[�p��w�D��U�]��BU�!���;9�|��BA��]G̳4z);׭Z:�Y˻d�\Y�آ��LON@��J�e�r@��\֯�,7t�X��ቯ��V��C;I���{�:]0N���k�S쌬zN�D��6��GtEܴIdu�8Җ荾c6`�k%4�����D�a��L�vr�KI��y�}aa�m�	�|wX������4�-�[�d���b�e����z�HN��%�-���-0z�W�<ܒ���if�ZtEY�3��wzg.�r	bYڷWT�z���N��ƒ�lUyDR�Ē�vY���ؐ���>��u�D���A��f�6��r��p�y3s3U+�y�&�ѧ�ֲdq��{f���N����hq�N�v;�79.�ק�e޺��@���F�C�.�����U�rݝK[H��;�"��g>8��;�m&������
�>9T�/����BԸ/r1��X�Y�)�ئ��'p��6K�k���3�e7y�H�s\S�U�Ґ�]�*�����9�d��n����Zq�ԟnM�6j�ݱ����ʮ����91\<jں��P@W����#���H�Y�#�t25]��oњ���)���*���g5�(NvJ�M}�����]���6#%��>�:����f�n�=N�4��Sn��(��i���&�s�����x�z�r���y�V.S�|2��{N�]��,��v�j��ـ礤_gjc$hGx��)]7���S�h�;j�J�"J �����������WB�6�����	+���8����*Œ��H`9�{hP����[��͵�eU�wMvU��W����S���&e�4��;��ɸ��n5�m�x����:����ui��ZA �`h1�掮fS�y*(.��l�7�H;���tz�!O���s.���}[5��I�4X��7/Qq�ή�R���7]y�'>�X�S-�����჏h�)�q�yq�e��6Mv�
��'[���R�S��C=�G�Ǖ!�vw*õ��ŬW���u#k{Hy��t�A]K�������$���iq����@G��0V�"�-g}d]'9<yc��Ԩy�z73AȻ�R���&��E��pq���M��t�k��]��Ga;��0��δ�mH]M�ݑ��oS�J���9[Ⱦ-]m	MtS��s�;��sz���VƠ{c}fؖ���bHV8���[�G��;ǋNY�ȡ���3A�2��}��-T�#�|���-�#���������.fl|!˦����j�֥�"������E��������N�eC!Yٕ�!z�	��Z����%]0� +V�[뗴�Civ�(��^Yvy���
�c�96��*�|���X��I	d�/�Z{�0��ܗql)��"�o-�/$z􄕗J�bi�o�6+���p���t�c�0f�÷�hf.�2�;�X�@1�S}qM341��.�hwh�B�ۊ�{�Bc���\12F�`�54Y��-;�����6bڌ�,v��k����E�7u�wF�ǹ3#tbo�r��P���
��o�w2U
�[�E9A��d�Uo���YT�9���8��ƺ�O�E�Bn��:�/��qA�������!��2m�j'!L<�$������a2�#|N	Q��!�s-���q�i0LB�ֶ����b���.;�m`�#�q�c8ZG�kov(˶nK(b��o�;X��=I*��]{˩�;�����8om͛�ǊmK�!Q{@
M�w.;W�^cs�Q޷���E�g�X��{[�{"�8�)�nfC�9\�eԈ�&��Iu�u>��&��=PK��Em�Fu��4_k�F_�wA������fGY�
�*=�ـ�`��,{ſ ����5VVb(�^�q���)7��g���O���&���4pd��9�>������]JnD�V�=�+`ޡ;.�D�hS0�0�Y{&C�IW_8��0v�+�`倔�� � �[u�.����3E�63����G��Sj����>�fKW�&�l9�3g]?�i��'.���ePL-#�"���9�?-�pn���������PS�Ѡ�)��fb�w\�y�h�*CҲ�\�ݑ1ޚ�;�����Cw2�!���p�u����(��-C8i����y�y�_vbT1	+��f��W����̫�X�k��dy�;������;v�R�Zy��}��U^*�k7�::���I�C��NQ��Q-�ξ��序ӝj	Aǉw�%7�*�����b�6bk�
^f� b.�38q��@�\BFH�e;�Z��_)�53�N��P;�ڌuvv�<�fn�ܽ�6��
!˵<[�.�,�f�m���[uq��RMF�d�W�/o\��P��|'EJ��:`%'/)S7����k.�T����kT7OM�ɳCA��$C}J�Z��Eo�Z:=���1h��I[�
��{��\��ty�j�r2��\<x�6���I�����o7�R+"�M�ʙR�|�DzVg!\]:܌ϻ��Z%�@�[H����:�
(%f�w�D��������Jǻ��ƧK��I;��(��B�tv�d�wm�K����8����tV�S�m��Ԗ�ނ�t�ˌz�ɬj��2��88"�vҾ5,)ڝ�H�d3t�tyry�V�WKAդ�mKtЪsj�e�G%�N��T�/*9�[�+�%Q
W(��@Y�5J��v�7��%��դ
�$�ƅ��o�
���|u|�A�4e�LM#��{�iA�ۡ��;���&Q�K�oW<�t�ü3��a	�;��!6���+�;�t�k7q>�Tv5�@�7n�O�Z��R�y�R��M��+#�a.r�W�]o�y	8;��i��$�|y-������]*���n&�a��8���n�fJ
�=NV-Q�C%��\�$�M�Sa��<�P�&�3ޑ�ධj���4.�[���n��06vK�28����]�tJp�S�{w��aQ�pt����:媎^b�ap���ԗ\�j�Rgf���S.����#����蜭���v�[(��V�cyu��֩����R�>�t�P�R ��J"�
P��A(F�g������ӂ|�=�Re�IѤ�awB�&��hY-�ʝ"	L��R�1Ɯj"��@�w����w�ׯ���绯?р�6߱����� �������?�3���cc��������~���"�����]1�%`�O�N�Q��!�@Ś����7P#�S�:�(��\;����n$k�J�W�f��r�1]e�f�0�b����%�`WK:+��r�1��I��vQ�5\�uZSl<#��5F��n�A���r�ԑ�+�N]��q1���
���]B��ZOd��*f���a@�j�li0�d;�.m��Q4��y�����	F��M\N�;�����Ǧ���9����$��gp�2b�N�=֠FT��
&�wI�k��	���W�A��ms�5A2���P���J����U�VYަ�*�=Sz�CهD�ǣ�Z��g[�5�_R&~���)v�	�"]��ei�aɰ2^��.t3��u���$�fЪ��Jя ;ˤu���-� ������߁*���ږ���0ѩZv��WC������ƊD����P���f��׵-6�M�"�;�mT��o2s
��3\�]ݔ�:b�謤��.+Sy��u�K��u�4�U�=���s������x��z����f�yM��ZRfuk���7���'�Z�vmR�����U�r�N7���*�P �ͧ��qPu��,��u,:�{�G6tc ��D�̒-Е�Ggi�{S�q��MΨv�Ŧ�&�QF�Ԭ�Wm,��Qhs7Yy[t*N�La�Lh���3�u���c9T5�#�۩�u�k�Q�R�O���}G�G��G��}��'��q�8p�8p�8P�Ç �Ç
8p�ÂྛHC��(;��+���R�U�ov�@�F2��q�tpA��	�[3�(᠑8{��r��t�x����J��Wt�q̵����ӡ&�<�uu֗R��೮�)�a��7yB��l|.#��p<��t��VЌ��]|- �9LreG�Շͣ;�9f�X�F����8�$��gi��tx��A}b�O?�#D�oJ�,����k��))c�YR�/x���9�-���i��5�&���E:)f�P���٢�/TaY�~�.|���N���
]�9a�����|.b������+�#c�2�Ǳ}G��휈ӓ�؀�&���XX���7�W՝�ޥCIôuNm�6Z�<�*�+d�fC�m��EY�n��We��tH��&lae�D�ڼ�R`����gs�xLV��߮���S@\q�gu�;��ڹF�W6ë�W�d�D+�Kp����b|�@t�ϯb���t��W�8�n�൹���(��M�_ѨQ�����OS�ܵ����e/�5�]7�-5a̕��i<�IZ�mp3A�`��m#/��Pv�4�^L:�;��Y冮%y|�:�t���0儍�r��Y�7�_E�X�Zh#)����X	�S�]������t"��!zB%�5�غ�gC��7u��;Wj� ���9
�u�>Tdc�]`{������h[Z��
�Z��]�WmuڏM.�FQ�3�:��.5xO2�"3�À@���A8p�Ç4hІ�4 �h4hѣF�0p#�8p�Æ�p�Ç8p᛫`�O�{v��*@V]�o*�`���Z�uػd� "-�R�)L���]X ��:T�.��5d^�ѹ9]�
��f�����8ޠ�R���-���B �g�jh���Y�+h��k3n�Z�Vi�Ͳ���Vf�L8/p�"mr!�Xk\ɼ�<�+8�aG5��X���X'Z��a����5l�Wt�p2ˇ(\œj���o�9��\��7�iM$a��k݁�����Z[�d��C(��M�	&�օ�}R� :K�4gH�ӽ�ko�����l�+6��Ї�k�J�n��r��e���kG�IݸT��]i�u�;�A.��͊��H��7#Cv�R��Q� ��X�ި�M���[���Sg.��U�+8ޅN���Jh;�EԔ���4:�n8�7Oi,�0SW��e1:Z�X����.XN�u��ef��ĥ�l|���<M��c3gK&d����.��z%	�(+�[�5������$�]	�1��qN��M���!L��{,]��Lz��x�nw�i9��Jز����z���b��lD�!�{�\�u�X\gn �D����R��7����23^k558���wMP�vv(�ڨӸ�%�E^�
X����#�;Ī���s{]P�ٵ3o����K�bciݎ�Q���Y'S�ΙN��uCvӮ�Wyݴ/4B�N��HqB�땝��C��S+���X>��I�V��g�C�Ř����Sk #����W����;�Zz�Tl��]]��Wt��y��`���p�[�E�[�1�e_r����3������.�p���#��c�t�\	KH�l��[�=��&l�i�o5�Π�-LY�$Q�!��1Ż����d�Eךq�ұ�{fA�����
;��T<�Z�\�E��n������VM���"�����ݞu
+,sb�i��6_+��*%������U�s�Ȼ�OQN�n.}� cE���Q-�M�Rʝ.<l�َ�ec��x�BV&;�������H5[��Tҵ�痤�[���&�|��)}�0S��?��E��]�b�V(�̫��n�T�O����Lg@���(�#__k�oR���c-�0֔-����f�%4j�bp��F�|�N��{��'&�l1�U��Vו2�P��$�^���9�n�7�!��^��u��]�����.<2���mBc!�֦�J�QG��:А��	���k�<9�<V���
�ɝĮ�͂`�K�2���_�6r1�����Ѻa��X��Dx�j�Ǜ7[[�c���mLp>�|���5�4ݑ�Wv�B����kv�X��.3Ap�_u��s�^A�K#
���7�����'_h�.�M�Z�"}|�M��w��2�#��A۫��_.�ы*�	��N�,:�@�����zH�GY���!����+v}O5w;N�t�!��h4�G��f�9���R�9{,�#1���Us�wQ��b;��EкB�o0�F�^Y͋��Uy0GP$�V���ݴ�8)|><^�hi�s.�X0���4�����ݝgp6Jj���۽0��K�.17�ž�Y:�*,�5qE���Wsw�D�%D윲��[���k'���Z��%�Lk-J�:,J�p\�����ʳ�LVr�%l�� �+"�+d�DV�5x���J�1�Y�RpTS�	�u��Y܉s��4*J�����݇��G쨦��90��ۭ���I�tEfAAf9�dh08j�ԏ<��]6t�-oa&�>��M�c���K�1�>�����3Pq:��$Sו�����T���r���B$n�5��S�]��Z�������*#����Fhf�.�M:�Z�<�Nb��[�&�+;�0ON��l��Kk&˟TuaDg'�^c7S��cWJ��4���Zd��ܠ���.�(s�Wpe	p�H*8�ڙ}ǯZU����AG��-�R.���+c��9PϷ��V7t��5�w,u�3h�W��3���]�ٺ�d��,}B�6�fZY�pI�}v��5qyt��S;Qۓ��8-.�����f�iى��c��m�*>��a���4a:H��Q"��V�q���&�`ګ�U�	,ڝJ۫x��%��}3jy���w�1O������VQ�,r�����}2�S�|�PM&�OAt�<їԊw���M����#g�ɏ�Qp�s�J��d�'dyv���(o:�p�:��Ltua����ti��v7�:-�sN��A��F��4C}ƌOt⬺��5�� e����o�1���N4GU)�6�x&y�Ĵ;�Tq�s���A�g,�2�����d⠰U���;V��r��<%2���t_>Tf ^͛��6�goX=��1)��c;X���O�:�6���a}�g4"��rխ�n�hs"*���BV7t�Nw��Z9����3H
_<^�pF�p�
���O��U�m���Lů1�{�Lέ���֢���F��'�0����^/�v��؞�&tw!�Huͨ�j�[��j��s��i�rwP�28�K ��W�|��ytgwmcZR�≯8o��A)YR��Z���t����wk����9(A]�곂�o,����	�5rZ����:�j�HeEa�U>ɂ������Vo�9�K��;YU]'I�&��1�̪�Ñ�}X�pUN���dɔm��K�T�u�x�YsWs����פf��|����L��msq�#hH]�}[V�T�C>j���P��v�E�#	!wa��]$����9,���o.w�Gy(�Y7m���&���>f��t1��T`9�u�ۨ8�a�(]����K.�Vs�X�f�.�:&�[+pޮX��H!/A���.��/�Q.� �<��ǵ)e���ľ�n�WKEk�LEۚ6��C+
S�'U���G���p��w�;!Co[�*+e,������E&I�ϓ�V�%TD��ۓ^A�LS�oH1����1�li����a�Sfv�����5O^���y��.�,A���S3�UuՐ�n4r��r�c*|OLzҡ�vJ��/��훥�+�UH�&�f�3�����wA�!���^d��ԑU���vt�{_�U+�x)t����]�N���@�s�R8���`�z9�&��䙰TY��p�L����j�Tp�v�4N �q��Ce-�>3��Jn-�(vDܰe����7fd�Q�N���͋<w��C5]\�ĳ; �1{�A��)�*=�-'}{- v�7:��Q�q��n��/TF���#�j��ǁw4�M˹n,��K�fV=M�<l��xo��"P��:V��Ջ�5�כ�S&r��vv3ᇕ	��0g�]v*��b
v�Cf��c�YDUa6[?u�e��B;�$ۋ*'�Q�$����%I�zf�W-x����wN��Dr��Iot�@�����K憎�vnkX��{"6�nҦJ��������=6,<Z .����[L�[�}m��/x9S.��#÷���W�l�Y�x��5+n�$/ve'��<���V����wXJT�l�\��T�N��Y��	U��8-�T��Kp��J����V��Fno \���U�L��⫄3,˳�Z�:$�o{�*�hl|�<"�]��a*�h��(����ʜ�vo'�|D�0[�"0j���U�8�颥Ѕ�;##A��`������#��Ԭr3��)ݝ���u�C�{��&� @S]�n`&��j:� 8�ȱ�W43�i����,�#R��	��Be^�������-*C�pԸ�N�r��O���������uN<G�J�Th�'s�#S�^ @��n�ܜ��AśÁ���u$�Ǝ��|�%j����C>B�r�gr��{�:��ܔa�$9�Q4ȱ�ڜ%�aIfX�]-�KQ*�ܸVں-M��}o��&A\�
��g��V ^0n��i��0,C�c�aӂ��}kl���垰�.��WVl�1�7Kض.go��~r���9L���h����[Dfo:]{�[�	��N`��q�7T�jn�p�6��7n�#t��ϲ*f�ً�nm���b�M�bt*Z`�'ע�OwMN�W"�nʫ;���S��K&�^ł���qU�ST�t�wml�/WM�
���G�w�wdo��ޜq��;�g7���Zܨ����/��n��vɧ���9� ��H\���+�8�VM�ai�����ԡ�	r� �Ec�5\:���4	E�.����Pc�������λ�]��]7�CAݽ1�R�81���'�bs���+���ҎͰ��N���/�%�|Cm�X�4�';���o����9�X�X��=hC�3�[�8^Q���6WV'���`��g�+����i�-�Γ��
������2�Δ���Hv�����Gyo4��дq{�9@	���o�ڜELׂ���e�{(d�ǎEz̭����q}*�v�� 2ՓP�sL���fŘ�X�j�,��/^�9�H=���$m�V����������;��զ\������jm��ĭ�bD\��ut�6��f%VBkQ��9����~)e��3U,Zs)c��ge��e��y�Ce˗FYܽw�4n�j��V7�NBuwi�It0�Z
�m<��(w7|\���1wi|*��͏�\��C+���h�piz,�ݧB�#�^A�\�*�����A�^��O+�+o��{O:YԸoL��7/)��n��]��wX�]���C}�uZb�ݤM΄�r7t�i�e�O�A�<��Bf�R��Ncv�nK��3���9��s"�t��C�� N^��O�,Q;�^�q�DCo+N+�|�EM�q�q����Ŭ�n]L\T �^�5l(��Rm��¬�{�Kr�%�p��nl��t����l�\�+��C�6K�hv�ioTl����{��ޥh���;�٠s�i�����:6�6�E r�ߤ��f�i�O�bI=��7&]3ٯ(r�Jۊ�'7�-�7��#e��= J�n%��_*t�uưn�edȦ�z�����3�h�Q�%����:Kr�����CׇF��&-[���gq��G�z��؃%�(�Xw]c"��[��Aa���tx�[���`b��V�*��ۙ6��D�#ۋ&֛ťj9X�ك����/�mti�{�d�|�Դ�8�Q�7��v^��fI���on�Z�"��wqv͗�� XŽp�ܺ���ԩޡO�o\�-���2��G�бT�M��2��D��%�̣�XU��I�Ats�Ղ�U�eӵ���>ޛ��ϲ4nL(u(V��ΒYz`� ˛ѐU8��5&l�5*�*����f���8�����'q*a{T�4�A���j�TV��h�I1�e� �Ρ܄���w���u�̫°�G����˃�V�ˤ�)T���+"�/R�j�<wf��]+X���^&��i��v����#M8�L��ʁH(�R6:��w�Mݹ۽��IMK��_��&�6�������w��7��������~�x����4w�;���7��(se�t��n�N�3�;j�J[��b�S$uo���9��ɵ�@��+2TW}n�h�3���:��W�I���Q�Uó��|�UG�����:!��=С,����<쓇eΕ��j;�3*��)[��c1��K�#r��NY�>Q�J�uϯ'A���܊'���W���[8;@'z=�� �@_9}Vf�f��srV��K2�J��Kw�Շ( ���bzIޑ ��Po�\gq;�e�5�LM�7���qS"���w�h�
⛮j�v̬�jO�1'��eh�����i���.�'ax��Z.�
�Z�͢��k�׀��;S�a�"�s�=KtC�c!�Q�S�S�|�V'ۖ���3yKyN ����p��*Q�f����n͎{��RAԐ#*��:�k̶_3���l����ý�9��5���`��z2��X�3���
��x*9��`v�����H�]�Ԫ�������"�7z��X�e-(�+-�[�ّ/g�*.�b�kN��5�G��6�Nt�kI��srj3��CG[qf\�w�aj
�X+��ϒj�9�"F��.���rX=�����P
� N��s����dt%h��Z].�;���MCD���TB��T��L#r2E1��n6<����V��k��:��8�am�(�gN��6���a�N�%�����$�R$ P4����G�Ʈ n��xZ���zxꠁ�_�Q:��d���sB\���E\$p��]U���a���<y	�T�'���{��^�#���0Я=���S���y/�!Q��Ut�s�-]g�y�$<�d!<w�o<i9�k%Ǉ����{h�JaI���y�2qw)D�����<�H�=NR�=֘UT�[�V�M@��6���E(r-TB�7Q�\NP��rGwW)c�8�T�O$�6Yα��$ȱC$7W]ҽ�n����r �5�q<�)K�.nW��K˼�-�I�wtG���]x�g��Q��y�i�;�s:�z�G�U9:^����y�Q����!rܯw
�p�g�N�t��:j'����yx��ݡ�X�|�u'W�*$���X�JVa<t�V�ȹi�ZT�������\����qH�O3N�Hs�r;�<�o)O.E8gFZ�Ԧ�%�<l��P����D(����'];���w$�
R2��C���cʈ�Tu49�%&z8�Ud��$�Ɗ P߄gH��k�3-}KaT�8��s�:�ګN^�m!�f1�ng�k�](�-�y�P7R�&6N���v��q��_-�� �|�������P����#��{��@��s�{�f0J���-���>���uL_�R��o����������5s�%z���V��(]m���\p�����
�!w	�
Ѩw���	rR��1]�����j��7�o}���E��T6R�	`��+)�l{�w3�����xxv]���	�vzO{��X1�`�#^��p��p�_O(1���'�Z�q�ާ��{�^M�܋���z[5�-��=^����z���r^:-�ޑ{���&�y�ک�{�Hk�~�]�e���̻� ��0�N\s���%
���e_oi?w.�������s3n��]ee��^XV�ni�O0MX�W��*�r(������5#�t������	+o�B�|!I�N���~믽�+Gu!�j�r��uz�x��ܲ!��o���h��`J��S� 8�2�4��L��a��{6p���ѻ��q����z�	�'t�Ķ�m�B�ƾ+���}�z�k�ly��S\�H��nvY��9Wj��[��=j];�y@ɡ�F)H[H#a�l���<{��0��v��} q�a�����>ڹ�R��R�zm]5�?%K*�z2Jb��9t���FV*��N2:&:�4��c��tφyWL��%�˰��+��w�⤫���7�$�A�ˣ�Yٹ�����꠆tfn�[}�׷SZ�>���}��[^�kg��ޞ���Tȼ5B�r��G��}���۾�`���WY�e�+�7�!�9`?=k��~;`��v����[ll�%���}>@�OG�I��ԍmP��XGw����~���{nZ\�����H����G�p��/H{��gS��GUi�����QY�;ځ�%}��F�gm�5�U�����W	`��G��^w{֎�0"�'/K�3���g��y�X�{ͭ{f5��8;����`�^T�f+J��0� h�^��GZ�_�ݻ]ӟ��!S�ქ�#A,Sۣ�*�%Zș̳�W����X��M�`�71Y�-�.}��u��.	��`�u�!'���G�L��Ws��,6M��q�u�n�=VB8_N;E��|�w������ש��u[�3�.N:L�8�k�����9��9n*5��N>*���ͨ�'y�o(]�5@>]R�n���c#��jv�>���T����מ�E醽��~�y�����}OrA��>>�>����u%���]7u�:�/�2*���[��`͓�lJ	��7�Ӽ}˰d��p|ɮF�uR��1�s/C�;h�S}rU��X�ޟn5��nw�����+k&���c�4��-�]z�O��l��.����^�z�tz֥�u/��Sڼ�s|5�I��8�����m�Jh�HW�����ʊE� ��.����'"���GnNY}�^��W�������ν�>���@�rQ��Q�~�X���%�MK���*œΚ΢��p��I+��ߏ��B��h�nͅ�l���n�x��:c��3�e;(`J���UT5.���+F���W�x�Ws˺�Q*՚ѴL����̽�Wrj%C���#��C���7,�Ѯ��T߶�a�$^��8_R���������y��n���ʝ�gs��(~���tR�(���ol�:�0�1���vq>ۚz���9�u�Cbr쩊�^�.re��r��p�;\���ҽ^y)w�Po�01wu�mJ��]s���!�#���8��+V�g:<w�}�)�N_�� ��8s��+����W�]��G�{�<�?GRD��^�t��]�6����oˇ-N-~5�����#*4 2����ώѓ��ݒ������N��_z����?h��+�䨪,��w�>>�ړ}=�d��i�y�)�����.�'��ǩ�Ѫ��T�<�?2}6��"�Z�ռ�=��x+Y��۩�Y�=���v��5�y���@��������}�
z���km�b[�Nz�7���M#On��R��<R�Wb������y���0�����yR��c���'�k�.��j����x�9~��ڶ(���k}u�O�i��������Qg��gۚ��6��+�+��Fj����u^v �^U���fCJq`�U�a��r��:Q����hl��xT6��o](\}�|Ù��������޹:����vL�n��*_]}/a)匷M�o���-��f7����,lhαE�x�fL���UFUȚy��ݡV|r�ҽbW��1s�F��o�J��� ����իJ=��m��^E������f߳�h��S�]?*���Fؾ��ԥΤΜ��6g{��Tu׾�\�k�&뽢�@��Ĳ���Ev�S��JvV�:＆n� ��f���)���Mz��Prcޕ�Z8����"`�فzG�ϮUǞ�7�����c�^���\Osp�Q���p>��Hs���Wc%|E3���ԍmz��,?w%eu����\���Ҡ���Ų{7�������ƀ��R<<�xy��GRIt��t��m�����vgx=�Ukz�vB@���dp���_{Ԓ�"|�]�B�׊�.�9�=k�Ck}�*��U�jR��0��b��ߗ����m:�m���y9���ǽ-���������{|ǘ�!q����J��,�|*IC9��\���=�'1
��Ji���z�=g��ւo�ymM�cJR���p<�`si�5f�N}P�ĻY�J]F�ھ�T-wm6C�Y|:Xꍖ�����@�X��du�#�KL���]��i����%��wNe� �z�ީ�Vה��<5�|��<�^�e�V�릤������ݘ��*�ҳM{�_nza���vOL5�oپ����f��
�9qs�^�������Uey��Kʑ+�^�)J��^!(Ɗ+��2~������N�֋�g�����PP�ɷ��g�7�����r����^�����T��k�m\�WN��U�1t�k��C29[�%�����+wK��MU��є��;/��v��<Dw��ѝBi�h�m�������m>�C����ջ�lw$/�]�l���P궰���Le�^~Z��U�k�^:���k��=�^���zAy�|~y������֞o�b��{|��ʢU��c7oR�{�D�5$<@�AXˌMeg�!��ϟ�����)��ޭ:8���Ѵ�Uee��jDV�y��*>����@�:��mr�SgB�ۍh}H���]�o*�-xU͝Cc1�%{���x����<��9=oܖ�;A:�L{|�r����j����&�0tE�qP�A�\8d���Av��/��a�z��К��QI��*�g��v�J�:��8��<���k��n���+�/xA�8Z�їfK}�.H�n��w���r��u��L����
����u����y����SX�g�jB/�a򎤖�H�`(��a O��0ʱ�R�[�"�^r���6�H{�w��G�+��N�o=�S<羶|{љ6���J�"]���^Y[Kյ�*�w�2�[�U�N�������H�-�����}aC�o��z���W]3���)����g�ּ�b����{
����и��U�${e���tթNg�M�y���*��dS'n�a�g��D�����L�=II��{D&���_JbS�)zm;���lf�����z�:z�kƪ���N2�&3�[YT�[ϟ�J��^���l����?WTxe,��g�X���Tz�R�.�BAm�^����S�f�I>G�.8d��]��~j�y�_�}u�w�r�a��ä�Í���-	���.��;�]%�
�����|��,I�}��ut+�̾
�E�%vkR1O3�����V�*iN��29��F���Օu(��,�3vj���lY��Ea�8�ֳ��&�۫����`�#�U�㷫���G�s�{�
����z+|ٽ��^<0v���O�\�����[2��s<�w͎�����KfN{z���J��04�>w�(u�ªC&����ٿme�I}崤���擾���Wwc����Gs91�Y�l���Ƃ�wmUbIV�I���Ђ���A=vM��%O{��'���{�:!B�c�ܳ��E��f����Іj�b�ǐX{�"1u�J�/�_�U�������H{�϶C�}�W�׉��t!Cؽ`G�DGRE.)RW�>>�̻ܽ�G+����Nk��-�VW���%%��l<)�4�o�� �����/'q�cP��m����q�ʮ����cX#��r�	^e�P�Y�S�1���7Y^�2z:MA~�H�r���&t��ǈ;q�W�P�٦O���I��/)3�]��Pr���9Z��)�s����Lv��Uc&ɬ5i���ܷs�Gك�}�#�����uX�� ��H�iż���t�g��]4.��7�(5&i�y�N ӷ�]Nx�R$����1��ۼ�ܮ��/�JA��_ξ�9���)}���x~����zC��T=�!�W�L��}��/8�]b��ԸO�][9�� �
��ܺ����;\���F}\3z��tx�lQ�f�Y�A:���j����ʖ���}�]ąk�.�p�������_?C�x��[m����J��k+�\O��S�ޢ��OM�ӣ�d��L��%�}%/ k�����
Ǭ},{����Fr��r�̫D��&�_F4ev�^��쩯�AV�*�(���@`�_*����n��uE��ѫ2�vz�^yuz�ģ���HP]��1�ў��G�:�U�bWD����(����:�����BO ��.�c<T.�f�������c]�Kx��GV�-i^߉�S�x7�Ӝ�Yu�˽7Ɓ�]�ŵ�ۼ���>������^��*��Ի����#�,?w%`ֈW�{Ū9ҡ�N�0)��UG��W�2=���!g���Ƙv+��S��w�^mf��k�G0^~���\���5�Ƿ��-cz.���a{�G���S73m�\y�Y�b�;EHm��*Uԡ�^���d�-gL�=R���_��&H1�;{u͜Tn�fl��(�Z��ؼ<���^�� ����T�18�|"Sλ��s�ȶ�p�C���@k��a�_l��ꪞ�G��wm�g��o�y���o����{�5l���H}�+����J��	�C�(�MVmk�T��[��º߽�^��[>5ޖ�Ha�C�+�����Ҵ�4�{+�����	:�{�qk�s�/gy�پ~���8�]��e�d���}��+�����E�T��_��v�-߫��V�}O�=��l��n�����^��yèF�B�
A*����۽G��R��R?=�ޓN�o-`h�VF,5����/�?A޳��P��#<%����ޗ�7�3l���۫���[�ܱ?�چm\��_U*�����#^e�݊�v��:������)#ϳ5���p���}}|G�����q�͏������`?[��s��Q�MC�0��?�
m�n%��N�6��W�I�9�t���Ls��-A㜔�{�M;Ty�K�U���=�8��2��vS�*:#.(*��v`ɢ"�/H�R*�_���7�r�"��V�tjY @tn���|�����.�F�%�
���9˪�S]N�2w#��i�P��z	)V�.�����.�U�<��y��NH��f4�᳗݊��Dvխs��g'ܷ�����Siҋ���2fD�ʼ�Q�]�.xF�ǹ�}Xj�Bo*jYΒ��D�Q�L��"�3�0�
�ovdı�w2�5.�We�t|�{Q�L{v��~M����[R�Ӻ+o�oa	N��YB�nM��[����\1��ڗF�(�Z+B���\k���DPF%W��[�b��"�"}6�	+�U���I�YƝ3V�?�-;��ҥq6�Hf�D���Y�;
-�D'�)Q�o�PS�S�悟c]2��l5%,FyG�
�,j��E�g␜N�u#V$��4�3�2젰�����Zr�m\p�^X:Woyb�온^Rc19����z��;���:�/C���A�����S��,ܑ���0F�N`�ONÃ3�WS�Xַ�Wan�ؼ|7��sxkf٭s�Y�v.��B��e1����;�o*=�r��i ���-MQ'��e���~���o����n֋/�Ù�D���Ӗ�ͳ�r����;��N���d?�R"�i�'o>�ĶT�e]Ek���V0m�)��o�us��Q�M���[�aQך�D�)Z�yN�~�3ݵ�4tt��/e&����ݸz���`ue�*h8��碌�U�⩿��*�/7RW̝c"����7����:���{(\#,�.�j��ȱ��ճ**%�)e�[�	W���p"��6�3��/J˛Hkۦ�ʻ�{��C
�cj�r�[�j�Od�[���%\{ܻ���0��c�M;9b'�)��%]n}pљչ�Q�����V�V9&��oo�j➸�zap=�J���Cܦ�۽&���n���4�e��lXpP(��8�j̭0�I��}�u�@�_��n�첺�2��ڡP�����x����,����W�`��I��w1#7��a��.W^��^���{6��9���1E�\�F4n�u^8�>#�5\kBc���Ɖ����KE�����j�����@<D��RVo�,+VMI���7��-S�en�1�j-DM�j�osM����u �7��/,�9��p���T��x�k&u๽p���uY��]޳����lT}�v\��򴭾s��b3�9��ں���ZB½�]�h����d�"�T^*�s*�<�C�:���xJ��TQ�5g��O.�r�Gw��:�܋l��Ѡ�78�U.�ܢ�J9�e�U��m�#�v՗ј��L�M��3��I�ޫ��T��֫��w t&H��`�F�|�J���l�������߯��C�;�♘r͙ea=3�ZN�n�x�f���"Jts�
\۲$�H�v�����םDz>�G���D{��-S��B钦����Ug1	$�RN�w�Kª�(�0tǕ��*�<>����^�r�,��7B����$.�W6����T�������)" �6J&��;�DyGTx�-�I�"��P:��u*�RE9�ty�9I)���(H��J٫4.���rN�u=S/:W���"݉z,�(H�Ν8P�9:�HUҖj����wV��ң�s%u<Ύ���ɹВ�'+���tR�8��eJ�gO%�H�IC����^w�^xʜ�*�d���^�}3>
�Bʨ5!38���f0ܗVV�)bt>(��y�X��w��ND�D�)$�΋ĺ	�U�חU:SIZrztr�$��p��C�n����wX���)�Ξm'�.�\iR�b��]���b�<8O�OYf��î�c�����������ڲ8����+ON�K@WM�o�\pK����O��wv�Uܩ�	�թGf����7��3o��*�V�u:kT��"�=�=���߃a$}�<~��3P&6��0yg�e`>��Q���{��tPӐ�����Y�ĺ�z��1 ��n���1��r�i�W��\��;�s��{�zj.*'�T?�N,������~��#ͳ�G�j�!�w��ng�}K'�4&NdN��
��}��j'�cdx���*|d\���/���^�B�dD8>�Z�'-�/�zig��=Ye[�FDdf�����`՛'�riNF̰�gp�"�6'���|2�0V��MV���U��W�0�6���{yL7�Xng�����pK��xq�:gƉR98�%<bA�O��[����{���~�n�:!ܽ>:���6yK-�y�8���;�T�����G�o9,a\�*q������������\�w��u!u�n~�*������#������O�fj����u�S�|���}Ä��
Q�����{�`����B�q�>�X瞈v�6�4�lr�ص�ܶTچ;ܦm�;?
�t���G��9*a��ϣk��튯�>+�3i-w@�6���Q��y��؍(�v�ec߮�C):��d����:�%8���!ǧ��
�t�0	N�)�9}ٓ��n�8�H���j���}/DY�,�N���)Z��(1F]�����ʧ��v��3�VE�$�fR����I���3���1r_Չ�q��n7�����5� �F�x�zZ��/��a-N�~���G�V���]j�K�P���#+(��PwR��Ղ����C�}���{�_�\�:�u��[Eˁ��C��ol�=�3�k�9`�#|�����6s5��܏V^̘~۳kz�1����v�&4����/�9>���xغ���:*�.
���~��f��T=XuUUzoss���18���������w�4�e��Nl�N`���8��ҙ�^rF�FYI�ݸL5��B����n� �mprͷ/x��d���f~�3y�x��:�j�S���y�f˸�V�������3Kh\�"��V������A9���6*ze�c��Y�_��$<�B��bU�9�a��C"\�\��`T7D�l��jy�5硪����^���Lqb􋌂�0�ѪXr��a���=��7�*G�HD��`�����]�_�Ϗ�n3pq�QBLч��q�=>:����*��x5��K�`�k#�&���p'�Pw��)$vN!x�ݹ�T��dY�l������Z�L���tۻ3:m.݅=$�*�*��X�7X�����mj�&����+�w�z^fnl�I˾�9]zk7��I�䋓<ۈaukkG����'c|1�W����=3�>�{M~b��^��c7^�/r��}����=N��V��h�n�(��G>�4��z��:@���W������b<!�hJ��ң��r��A�0�	�j9��JȈ�����E;m�:t�tT	����%�D���wes�	��H��ۑRn�s�9��Ϗ��/}y��SC��������L���p��2WZvL�ʪ�z�O�veD������v�ic��Ǡ���}�u-�W���GS�y@)(���F̂�L�O��[���
��X�lLfK�}>���>UkӢ7~I��F>����N@�5@�{MV��{�>��d�ޮ���n�8����8�������V�#�৭��t��}��jAh��W1����Wh��[���1�2Y�	�"�tX�:��q�o��6B�v}��j"r�W�u�@�5g�O��:�C�����{��h��x��v�D6_n�F��t	�����sW|�F�>�{�^���E�
�] ĩ�O�J��<�N��-����x;���n%���w�f��PVR��9$?b��L�����=1���
m��v��`~+���9p����kmY�	�WV�E(E/3(�mh�b�Ѥ\�N}�	o]s�3�E��]�]�J4{w��EI��ʌEh]�qΧ�f^ַ���+}���t�X��^�7�,$$�A��Ϥ���CҼ~Q׈D�r 0�������dpX��?`�o�e�4��>��`���Ɇ}�u!��?F
Y���*���;��د���8'��;�:���)�r�3/�z�o���~��LC!�Rd�^� �"����� ͯv�of�G`0A�v.*ħr�j�ޝ��~7�V�;A+ƈ.nF���l�T�k�s0�[\��}EG��Pa�!�Ar-	��]�m��v:�)�-�_gb��Up�y�Xzy������j���TMY��������C�!�������rI�՗^�WsՓ7��#����t�«���ud&ˀ~t��r�G���	�.@I�zk:<"�w���&���Z]��c�c�/��U6;h�p0��/~������!R2���z7*ì}=�����eN�����D�j�����V��A!k=B��+gb�m8竑��D�bf|�lNGD�^�-�,M1��z=W�z�.Z�0yyx��e\��v��)�{v;B.�F��#���~���}l'��R��gsn���F	>O�Yy����m1�ܔ���|�R�Mw���$��1�+��mz��q�\��ig�E*�̾�(o8)�b���X��e\�ˉ∶r	�7�}��Z@m�$k��F���;;������e�nҲ���Q�&�J��������/��xُ<J���;g��~�D��\ uMף����z���񗸯��ۈ�d	J����`�F0���|c,�e��3�.�.�;_i�D��k��~�Qn���_+9���;�jb;|�A��B ��Cp:,6G+���� ��z�]c�q��"=a�<�HO�(-)Q��Z+!A���$���
�j֯n�
�M�ZLlČ��W���
��=&��?��t����O�SbO͊_�јQ�g��Q���b���q8�؏����K��Y�lԩNNG9�k=8�..:w���1[��u��>\�/%P�)l�g[*��/�e�A׋]/��]^_��Y�T���V��F6�"�۱b2{�2�	h�n��e����Y��o��	�XW��<J�@P-�����hNr|'
�ήo��3Dt2��/�nz'�w�'X��[��S�����ڪ�D��7�%0�m���j�E�lO����<D���9=Y�&���W~����#�w/�5�j�<e��UvN�A�spfv§�zTD���B�L�*k�BU_#��cj��A�ʗ��I�N�Q�Y���?;2o�c�&|5�Ї7E�[6��q���zk�m%Y��u��Z�ÏwJۂ/c��}�œ�o�Idл�d3��9�"�w#b-��]M�\���`�p]��=��O���" ���;a�rf �����=�_m�����r�쪷/X0�	��# ���?N�T�����,Z6e�u�i?�z�X�ۈg�ЄW�`-�R,��s
m�l����ޡ��y�w&q�������P���k��T����\{>7�8��c��[N:��ʱ�5�7ٙEgW�f��hd�v_ۮ,qJ��Ώ?�,��ˁ�5u�1����gy���1�������f�9���j�c�##��s[�œQ��/r|��W{�b�߸�z^{��u~�8'���اX1�oN�g(ܨ�j�M��/�n�' ډ���}ฏ�W_�/~yό���*��sn1ۂn��m8�y�.�����������>>;'��#ӪT��b�A�'ڮ����P��OF� x�)���Ȟ!x�!`՘F��!��EAs�%Ƕ:�\GB��`�@�#�O�{E>�$���\�?n�����Cy�qҽ��_ �� 7qҚ͋�C�O<�r���0��������D��/�R؟O�y��o�c��[�u�[��E=���Hf.%I��@ɖ��,�5���ǧlf�X���JY[��?'�X�l7����7��X-cDd�'�S+���::�{H~�m�1��#�H.��;Uv㆛�X�)K�|z��(��>As�*���1V����U�p�s���S���~|�z�;p��?C���7ϿϞ�￯^������aߦ?f�BRW1y>�rzo&���3Z��VB�\?��������N��Tj	��k���ћ;�AR�(H��W�$nMC���p����B�!r���3�P��bYӺ�3�=w�<���A�ßF��.�P�g>���Z�\ /ʑ�"#gW�~��9g��̐X�0U��}�L�~���}=LC���/ ֈ/.�e�h�L��b���L��K�����<W!l|�.��+�D��xeɍ�.6<��������j΅�f9	�º��tEK�"��f�H�U}�q��KbE�]|�>ژB;T!�Yp�����򈨆��Hb�=`� rH��R�Rfw&�X��1;9�l!��v!0��w�cڷ2l��w�����0x��N|9^CR�wʬ(#�ŏ��Y��W��}���V)x�K���E��tp�!׎��˭�@�a_�:�j��zf<:�[>�磼�<�K(��2ѳ$�����)`�K��n�1L&$\>8,��x�� Uk�3e@8�8�;ϜzE�)���V��j%�n�'�a-��f��_�p� @Y���f1���a�(�[�v��7�W��ͽ��IgjJi�"�Z���e�3�+��!,]CSxl���׭-�uY��׈ �H�ݸ��,uj�W4�{ɜ ����������+㾏����#����N�k�X���.:�O�E�]��G�U����z��S�Ԕ�c5�R:�k��AHG�]k�Qぺ$Q�Kl0$!h/�cWD�sd���{��l��zϥL-�üN��q��ɡ�->��.#5��Ld{�
g��_H�W�9�'�QڿLCe���o���}��
g��5��<�ٮ�J�;e򻨰�+#���*�O���|g�e����=�QD,�>�ב�4b�X����2��Lv�v5M�!lrKq�͑�LY��}oC��ͽ)΀Mg�#;Խ>��&���L9!���i����~,uԥ�;��oTGЍ�b���n���������B��"B��V�
S��>���<����,C_=�
�����1���_Q+�e��Ij��O���tjt���t\H�)�ܡ:c?�ڹQ��O1n7��ͩ�cB���M��<7��fX;/J�3>]{�س5g"b�AVE���t����}�����[�ޓz{�><��m_��v�8!�dd�z���,�|(�*AɆ��%�{�=s\X�`Y�_��љ�����*�0�PX{��.
F�R�Ά'
�/�~������+�}�U:��E4v���<�A������J����r�_V=6;������\iM�1�t�\���xi�'z�T���G~�{�>}��}|�����I��#���
D|�wf�x�l�1���~��J�{
�.��^��ˁ�����j�3��)�,������i�I��}θ��j٫l[�/�b�Z]M��r�5tԷF����x�{�Da�õ1e��~���yoa�`�GC����A^����xb�sс�P��3���C6!��}5Y��+�X��r /���b��G��\��@P~^^#3�W&��.d����S���A��ڻU�F�1h�/��>���p[�@���}��F=���6��J_�Ӌ~���s�e��z��,o�)�9��jݸ�!V@=="�L-�!��U�f=������^=�E��)�fW����q�bW��Oܮ��JH����?
�ׅ5,x�X�R;&y	���r��qj��_�B�#ޱ��Jx)��Op�ؒ����+!A#���ҵ����[�(����7��A�9dJ���Y�x__w�t������ɰ[1�k�w�O�pQ�;Y�[�~ьs٫MT�ʸ��^��6Ti��ns�g����A��1x��m��P�E��Of]�8Swۛ��*�E��^�H��s1>[��3g򽵫�N5�D�2���7Wt����z�`A�y�핗t�j�%�M��Iȯ�e�ˆ��9��-D��CV�3�Fk��ukSz��]x��V�h���e6����������D0��W.�q�pavˍ�Co���}�~y������<��S�2�]�i`�����~_����7�d"z��ߍ���H����)����f�@Py-"N����94��f���񛛟���� 7.��H�D�7-�p]�9��~���T�8@cV\�=7ݪ��Q���Q6�a�v
��w�yo��,��}�g�1���ަ�~O�Z+Y莖�|�\78>mY��2ˌ��՜�j��Ɖ�N�>�MP�ࣻ�tR�-�󪾘�*z(�a���4幅4�7�2e�FWe�c�T�����Wyn��{Q��r���f#=�����0���E�[��U)�u�����V��ʻ��b�
������T$���}@/
�u��j���*$u�&��a^�s��tA�۹�����q���Qc��Y�V���������G��#%L=5���Ѭd���*��g�6��o����B{^��卅r~J�K�&�s������#�@;��3�k��������m1Y:�6x�h�V�l�u���4�~C�鈿�Q1?P6�/�pq!�}�~_?�<���=y�T?
�"�0�V�}�dF�^���l֪�z*��i��4QR�4d�ik�[J'���7C�N*h�̩׶�=��)�'���; 2r�B��z.UL�A��N�\M�ȺH��	<�\��Y������z���\���x��wXn��w7)��Ӭ0=ˈ�����T�leY��
MQV6Q�5(�8	�ED�A!�f�ݵ�^��*���^X�s��"eN ���#��;�n��5��2�7u6~��ap)�6>��w�0�S��㧂�%kd���7����F3��:���ǥ�Wî�Yʓ�PP�x�����umM]�M<���e9�¦/�ܔU��$R���F�i��\��*S]@��%ݣGo;2[���c{T��a�#�H���LdǓ4ŕ�f�U�C��j�{H�����b85��	�c'$`إ��::�R$fS��RyCvu>�)l�h�Y�ӈ]�"��ݼ�/�W7��|���_սl�5ݛS:N���v�ђ�t����Z�O��w��q�!��[�B�AY�*����Zrs�˃fH�Ѳv�t��n��c���q*�P&�X�o�*xb�2'
���Cr�g���F��(X+��QՎ�.��"�Fu�vM�0�l�N�[�\0Vp�5�V�����X�)�ռ�Mf�E�x�ProT6A�: �ի�fi͗}_�۠��x�(ݡ�\۫�	*�O�ʹ�`�]�v�m�ٜ�bt�a4%8�U���W�	�]hZLY�x�G�%�뮪�F���ǇV�W�16�~���ר�a���&d=Y2h�ӺV֨�o"�*�̎���	�;B�p�i�a�E�4lvD�y!4�;
Δ`۷rt��[�B���x�7 7�a:vJ޺��t��t#������zu���ΝUx)�r;w�qa	���(˹�Y"0�^�U]��AP��[S���=�x˛xk������̆�Ԣ��������<�� ����h:�:W��q�J�33��9�x%!�+�=��`�a\��3{�P`��d�2@��G,� �')������(�m��+�� �Z�82�LVC��b��(7��@'lZ�n���1W���c/�3��e��b�ܢ�k��f.7�p|�̓�b-��^E�)�X���,��Q[�.�=ۇ��Ʊ���]�9{a�v:)�[AvU%\z��qN��zX+&�hS��Y�k�vr��A���C�R�S�Z�OC�9S"��j�憵K��m����OF-gu�hX�F����'V��S��;ݏC�Pc�1+����SFV�R�}J�����������2��g5���g�@��vV:xg �B�=E��u-�GT��t�7�%P���ʁ�l�DtkHMϻ+��,I��q�zð}|z�꘹5�)n3Z�s���J�,�䑜qLT��䘔i�������K�r.�����Ihr�����J�Fv¯%]�7�
6O<z��<�%���C����"*M'���tRI1��מv�9��'I9E-4r�\�L�dDi{}�G����w��TiĬ�>������r<ʲ��vQr���ns��)�3�;�9z䜤&��/G����{=ӏi/��Auq'�;�z�OlҴS5/��Ӫچ�É78���
.!M���jEJ����oG�3*���R�Wpzy}^*s���"z�vs�z#΅9��c�+�'��z�^��3IP5���yU����JstI��T���Nt�/Q)�I�ϕ������;�Ne��.���s�!�wyw�Xx��=y/�¤�\zt���H��y�|T��7z��!�=���(��;��k"�B�����¼*H�p<v�ܹ���R�n.+���: yc����o:-���T�O]�n{"%Ր��=<���j{=�C�E�ʋ'�ܹ|{��Z��u�)9Nr��>	�-Iw��3tw%����^���v�x㻹�U��;��oQ�(·=��'<���"��W�;�J�Bx<>yxW=r
=Nb���K�--6QuhkǄ����/}���j���y��/&}V��˫�**f��j��=+tjo2��o�2J�"6�4�չ&��F�P���ʿvߎ6��C`U
c)��q��
�n���}�}�W������y�F,���ә���t�����~���Z�3@[��3_l{��;�̏��og�
�����Zs���Z�����܄��0|ذ�~N��=}CƢ8n�F*{�m/44�:4	���к!�R��{+|lz��Dt�^�\[t\�x��J�pp������{%�z�)�`r&���l��"k�P��Kc�Se��7�'�V�_��!��w{�kx^�5m������s�ǃsP�xk�14r)���KG��
E+`U�^CSĩU���D�9����,?Q�#z�1K�ylG>U��?B��?i��ġhH��C~��t�{r�<�~����{<��r��ßFTÒиd&��T��*G��{���#0�͗��~b!ȴ�W���h��;o����鎖!����y��Ax�pE����=�~��x{���8�yR7F�܅����"�-��2�Ɖۗ:�6hR˭�rł0;��b�c��7�Ȫ�l���]�ꏲGq!��{H�ݾ�q��R���[�ɋk	��8ʁ!��Q'ߪ.ݾ�F�n�F<�t�fJ�"#¨pvoL����q�%al����9��H�9u�c�F1�lҟ3Y睳.r�k�ȗ�Ꙩ��3��[@񮔎f"d��l`�+B��Ҩ6�$'�ǿ��q���l)�0.�� D��v�91��.�&a��9q��o0�<��#�:���4�Y�+�$L�M@�����T��)��y:��<.��[����ۨ�JK�+�j^�4:,kQc��=6~��270C��}ъ8'k���2"����u�y��Ǡ��+rۓ�7jkƠXsS1ٝ���tq]�$��d�q?EF�23
�8y��xWW)�"�w2�}}�<>�aN`�A�*�.���N��k�> �"��u�b��Y����w�����=o�>n���pWa泌>�Ν�O_��P[��� p����g�'\����?���м݅p2;��!A]�ǶL�a�+<����y�و���
g�q���$���(`N��ܨ�����c��=J��V�%�s�}�Ҙ�J���Wu�L-"��!���=b���*^\��~Ң�߽�]~�G���m�$;�1Wu����#����xVC�5�"	6�b#�,��賞�͂�cE.�f���9�&��#��'ަ��TÒya��?E��>�����0TmԔ�Q�P��.��i8^�#oH{�^���V��;���nUk�.��
�#r�#W�>��G{Z�z�M77�#�'���5� "|��S�#�yVɢ��o��[ʔ��]���R�C�p�iaEwwW�#!�����u"��o2�����~<�<��F�8��"�928���Q�����
9����������������������|���yȝݲ��^�����'A��!7u��O�ؓ>�mO�ǡWN]9����1z
М}qa��Bt�5��	�I�{������mIj*�OOμ(������ĝS�(�e����l":�T��7+����˯����ت�:*��0���g�wK���[�&��a�)�Q�P�C�(����;�@��%ey�ʹ"m�_א�˷�ve��G)�˱���N�i^I��r"�`�Q�*����Y�ޢ-�s��d�\!��ŵ��{&ܸ捵/c��#Z3B�eF���ٍؖtxe{NwY�b	`���j����-��A�ge�{�/R	Z�\�U�z1�P�w�θ�gJ=�Z��o_6䞆(� �܁Ϗ��Tz.�W���YR��
���f�W5�ߪ�>�����s��Ƽ3��nK�/O� ��!|��1��Axw�g���j<��*�pM��f���i�<�8�;�yIN\�x�Av�8����@�A��1\ډP����*s�X�
�c�yW�5�W�LDռx�FZ,��ד�,8�Ƌ����H�ه���,�{KVՉ��P�	�3R�ٱq����{Ȝ������`�k3�L��um3�G��3�Xq֧�&i)��)�j�mg�!ͽX��7:f4��,�w��������|������}{|����G\��Gp�v����8q���׿�^�������?������#�;e��5�}�_�U��r��!v\B�*c���}��8X�,ED��v���ㅣ,��&4��H�ʹ�����>ҕ�/
�Q�L­��c����ig��=���>�}h8Ȑ�f����H�W��v�)SbKb���=��~9>�J��-�\����^F�9L4',�X�P٭�5ݲ�#2��&+��aȥ݃�ٻq���b7z�j�f���� �ՓZ}�h���`�;
eĪU⸛��{j��Sbs����?)4������76����@pSZD���s�fi��f�Hȯ�KScoo�������b�F]Ӧ�殹{��G*���15e�|ʽ�WVl��NM)�ٖ��E|c^�T��u�{��%��D���X`��z��ÐBUpܶ��V����'`���̗�G��:�qB&�:|����<%�ԣH��LF��h�_m��'�ܷ;*����2>M�<.>͙���o��ۦ���1�F#o��Q�\�#=���^���ө��r��N9���v� ɴ'vՠr�[e��,�y9_|��1yx-Q+���i�L�cPx�Zƫ~��0�~�b#���M�;*��2[���}2��K��out%<{*�i�L4�ξ�m��K�j�ֲ�mӌ1of�؇F��ҶY����?F�!�a@0���\ �"m�������}~~��}|��.��U�H���� V@���J��x�P��u��󪈨6'}�OwkޖA���|Z�r��g� �%:�(y�����v~��L�$xi�C���3�f��^.����K�s�q��^��Q~�іu��|6M�����9�}'�F���F#��p=�#<�x.�9�i �|��Э����Ƶk&�<�������j�@רP���{5��Zo�j�&O�ے C�m��Ӷ|�:s۝�N���*�=���>����D�4�D�]�cҦ�&b�k�xg0Y�B�k�)�F���>�+ܼ[��j��6,?z����du�D�睵syL���0�B��L��+tHR������^�n/��Q,��W�}r�]��}�����ۈQiR��Rzo&��$�P��EF��}-���7Ǫ���ό�<*�ٌyY�?�u�!;n`�5G���G"������#����h���y�U�7�*oȭ�Xm�ܖN_�g��v5�bGT�8-�&�bH�^C�_�M"�[���&�6���/�޼L*Q�XU������,vb��bT�u��췶�Úa#9\���P�+�tL�6���ֻ�z<��3R���Y�{ْ�1r̭ۨsP ˏ�L��6e�C}|v�ԉ�5�}��&�@0�K(����~���p ���p��Q�-3@�_�E{f�w^���O�o>�Q�#��s��,9A��Bh�$��h�U�����%T���o����:��ExPR�FTy{�xm�C�|�=1��ts䨿��Ai�{J���v�f��o��c��d0�eO��5b�}AҸ�?D��xeɍܸ����uw�}�;S������*�j����#e�Kf�H�U	�l�}#��0ؠ�����1�)�@��E���m�^���P�(��v�
���GX.HM"
W�O�;�P0Y�+�G�;*���=v��E��8z_��ǈz�E��m����������c(v��ς[L��Gp16�#2�>�����pB������`^.[O���'>ڄC^5���)ak3�NWW�/|YE�\+��t���:/���GŁU�H��$��=OgP,�ν�1�B��֑=�ބ����R������E^ �pZz�!llˎ������#�CR��������Y𾂅�fwS��̟C�K����Q�O_! �_P%1lH@�9���ړ¸2��`I��W��P/¦�յ�+�2+��"�V�Em>kJԴ��!U�V�}o5�t�wR�$d�{O~[0���uP��c���%�&ų1�:�*yz��v^�����:0@,���$|��;l��71aT�G�j�Ec���Y����]7�}���������dq�����m�>|��K������>��z��?s��C��ϸЃ܂'�h�
�p ��9�p���w*guv�~g�ް�>����*SJc�+�^����^��P�<da�S��o���س�Z����力��;��o��n�!4Gu����"~��bG`U�T�Q�k/�8l��ws!{u\��ݽ�"�'�M߳��yV���n�`�uɆ[�>فDߑ���
1��{��9Yk��U��h�?�U#~��p<(dJ��W�S�]Bs��C�X3��v��:eF�� ��Y�"��\�X͚�5+ȿb�N.$�&�	��C}9鍍�_]�x�B0���1�<���f5����q���#0.����rj,Ș�d8���A����b2ߧ�u�oe];W�����}�Z�%1nUn^�@p]�Fg�&��a�)�Q�d@vdMSi���BG�L���)c�$�A��(1}��c��z*�n^�FM� �=G�F�.ԵR{5��UOn�\?Q!-���Ɛ�W�Ų������ƍ�/c��:ј�:ܩ��ɥ"�����y��Y;�6m�e��9�b�`"f�Z-.�5��¬�o9B&ACl��ʭʌp���[�)L�ǎOK�~0���s�2�a4�'N�F��J��e��R��r�c����
�Thn��\F�N�_L��'6p�Ӫ������~ �)��6>�����>�;������r�H<�6�F�8o�c��=;�?n0V/R	Y�1V9趯�w����/��z(�E��d�8��A��۰�bPwg|?x��z�y��s)7�H��|v^ү<�����X�O��:��>���h��!��:�_/�/����1�uҷ�GV
�l��J'����|k�k�Ԛ��;����By��|�߁��T��E�t��c��5HǶHz�!�V˅�9�3�J��I�w�Wd�w�P�#�1y'��m��*�W���6Dp/�l�Ft�5�yG�B#6�t�	���9�b���7G�²S�T,�ЕT�6��/1Z���a�� 6�][�S�Ʒ��V! =�I	SbHlPcc�U�(JM�����k�2��0e���U�w����N.-��n����g���ǡwy���B��QT��2�{3��iw_ٸB�V�D�z����j,a�4|�N<�_�`����)���yW~���یN��tν�������dc���5�'�}x�윚g���#!P/�h���e!�7�P#$R�˔'}�"5S5%<LwH5f3�������7���+e���Af
G_U�=����X�4&��f����N�;pv�mD6��!8�t��ωګc$�#��e|c�jÇ6X�3�������>>���{��|�^|_'��ȣ��c�M��el.1�ߞ{/}����������^~k��/�@��?w1N3�+b�Yr�T#}�11���ļ�P�i�=^>D5����$[�U��".؎BW����=L9���s��f|�.3Wd�h���j`*&`����ڬ���0f_�=J<EU��i�.�{b��k���-�)L��Lq��t�J�\$����Щu��vZ��5=����¸���7qx���0���P��]�0�-��%M�QB�����3��z�GQP:�V)3�� *��a|�<���N��ɸ�5�ڋ�P�T�s<s�1�V�ڮ2O��s�a�JH�Qc���Z������lJ<4��n��8�:X�~���3e��cp?q���zڛ{C��{��Hs�;B�3:��A3u���#�)��6d��ڎ�C��*c%�2A�{�6#�v3;��Q�Z��y����7���ɘ�f���m
g�(��ݪ?�K�C��Ɲg�u9���.�G,�g���_�3�Ğ���O�~�'L�kA���r�<��N:'�r/������DO/[r����h�0�����j�ߞ�2qF�|������*��v(�����D�K��[�<CfF.���Ywo�}� ��Q�"ȝ�����Υ�]���@�_�h�U�Q�[;+/I��]�|�so>;g��o+��]��������<����&6D ��� >���9n��c7��m�dxq�EǻB�������`ņz)Jvz��2��Dt�U�ϹMJ�l�%�4�.�Ǟ��Zc�Dt=k��q�����"Ib��et_�ͷ/��Ց^�T��#ìi9��v�3�ͫ���3DwZS��!�=�֍Ŧ~O��^`m���k�z��gF�p��������svk�^�;j�ČR�8l��M^ĝ��3�2%�hq ���s���QQ�Q;ynw����;��7��@w�g�k�/u0�EZ���иi�؝�|�ħ�n<�����U�mNPk����"�B��
x��}��=��pki���b�%E��ȕ"^���i��A�����>ߦX:�� ���o�KX���������߈��c��ێ�cW������.����|Z�f2ker�;e������E3�v>��B�_�-��!�p^���%/g�ß�)�0�~v�/������8Lus��#�.��~*}�Ոa���
S
��Y��\�θ廳�:ƛzK�}z�E��m�9�W�ԽSC�Z�[W����x��I' ���sVP7N_��A�zn2�U�S�c���C���؋��sk>Tp��!�b��H�N
��O[��泂b��U��yU�p򋎫�r���k"�mH��l�������VV'#'��n���(���O�ll�R��r�f5�B�f�3V.H��N��L�Zb��*�������a���j�w�ǻq�ع�����|�,͝I�BoP<B�ȴ`(�/��]���fY�>���	R�������kj5�S"�{β4�@��o4�� �U��(����F'=�t(<�n�v�'�Q�z��H�x*���M�rDP�n�^`<2�v.��;ZRKvPn5�gv�$�5��GFNY�M��K��<v����v���F�=��n5A��u#h��T�X��XkT��������5�yp���%�MvvZ�T���Ȇv���:�a���M�+zc��Q-ڬ��S��F��v*��ۙY̻L3ے��bU�	����u�;�vɩ72�j��)���t@�[0�]����mm��UNw(�Y�K�h��s��MCu,��̬$�����cHhӫ�ڛ�\��ub,��V�n��٠�+�SN�RK)6�+w��j�j��q<���9Q�{A�kǶ*J�c��j�q^����@؜Pn����ƯdL�[�f�����т�ޗ���L�]Qd�C��W�MQa�1e[�����_��7y�(�Ӭ�qaGz�cv��O����!�8;�4������� ÷{F��>S�J�<u��_��[ř�b��}ǣ{O��k�0FFb�ʺt�#79a��61v�Q��F�|/"�����$w1C�i��+�kH��
r�Օ�tMr��v�C;#� �.Td��K��8ܹ8X:�ެ\�Q�f"���>�F��B®���*�E=#L�*��[n�#gc͓��l�s;�U��ޣ�|İ�t#�+S�8�{'���`�m;�j��};9d̺}���}F8�[b�)�z2��NN��C(�+�8�}�jgl��a��=���@.��!�s��9Q��V|�bia�:O]�.��87G.;�����̢jj���B{�d��z{�0`�VL��ኢP]���A�����y�𪎌72��w�8�VD����Qt�u��H:��qr� ��`�1�.�u�{p���9�kc0�A������orO)Q�����$�����E�㋗mј������A��ccK���M���d3��2���&W\���!c�����o5�,c�pO����76��	i�V0m8I7�l�؎�!�tNI��]ܬD�d�L��v0��,���w���e�=F�<v�G	�ݱY�>J�S���gb�gX��͞✜kQ�/(�O2�h��z�rt��EU�8t�i�4g$������m�_8�=2�V�z|�n[�ݫ2WsT��q���d��������t�s5�	�>$�=�;��!L�;��BZXI�LHȤE��}��g�ةȈ*���y������.Y&�J�}'+�a{}��c���=:i�IT'YNE!(���*R�����{=��S(/9���f&ft�
)Y�!D{����Z*�Ukhӡ	+	$�v.H��(!}D;��z�䡲��E<��<�e\�%U.Qe�Lzd��w���x�D<�۬Nz��r�%6'JK�9����zFJbTUPd�a�-�"ZfaU4���^H�q�'8\�
I8�XF`�ՒIAEό
]ܸTr����O�����/���9,��	֝���t�T(�qd�*�G�N]����QE2�έ���A��Qf�,�5�ҡCCY(Z����d�$	,-2�i�Ğ��kE@��T����2.�D�QQ�P���	#LY�H���w Řf-��heaΡ�:�'α��I9���E"A �JAFP����^Ǉ:ڛ���7c<��\FȖ�r��jQxl�B��Ete�o&�\W71�iw/�z��������޾~�G�ߞ��m��!�$| � ���ZZ��������O�$q��`�b�p	[o���nN|ݨG�j��b�ƛ�oL��M+~k1|LC�Ģd����d$o	��.�8F%4�A�L��}}څS^��Ko"�A�cmcT_�{"�����W�D�G�`O���Nltx����V�#��J҅ڙ9��Os�_2�䀹�`f��CZ/�A+U�
�!�OA�m��zb8�O(�
}�t��7t,!D��Cq�{/������/�c��=="I��	��{4�:/��a���V�lw_:���q�`^�P��{����>�6��ұ��*�|^�O���������[~��kp�Z���������
��MwPI�)�b/_I��T6=����(Ċ��2��s�F1HD0b#��#��[:=�Xj+q<>�M��¹0�~A�ھs£zo>S�w�R������y�G�r���)xR�ķ"�wN)~�ы/��!s��d��ỵ��ķ��G8���h�կ�%�[���Aћ5EJ�=�^��	��ؕ�?\���������iU�"�sEd��6*P��vؿߞN�w:L��u��y�.m���jOA���o���Π��W�ч~�{����=�Y2ym�(�;dnb��1\�*�u�7�:i�P���D��=��I�﵀7�NG��9����nVa�^��3��J'� ����| C�7߿g�;���}��{��}?���y��h�򡕤f��'퓓Q`��q��Ȟ�]8�v��\�'�u�f1�|~��뾂'��*�/�����~qz���)�Q�}6���5�e����``�]O�K".�'�(1`v������W���0�v�t��W��iX�����e^Y�nr���!���T�>��B��X�~[ ���\�ѷC��0�[�軾&��i�a�C��f9�O�ǁ"0��|4r��:��A�A{H)z�H�Z�\ߓT��^��
�W��b��~�w���9�v<A[��}���D�#|''�]����� ���q�����=�&��T��n�4��t���ÍP�@���6��"_��3[}&����O�0��r����A�*2;�} ���N�)˜�!��G�d	V�$p���3��w���\�Pg��Ɍ�e��u.~p�9�3�Wճ�]���U�&�U����N���o�76�D0��p�B�{��w�2DFHۗ�hG/�������S�����ؤ����_��׈a�c'�Ǎc�	Ԥ��M�q:�.��)�SC��	b�0�n��A��,뉗fI9音��'�[�9�}��T��op˾l�u��$8��ab���� ��6�.D˩��,f6'v�ne��{|������|G�]��wx���И���.1����_���������?>�o�߳��ϹI(h=_AK��k|;�#�������4�=N'*�%��v�g/]����bx��(�}j`��b�ciE����>�Y�ſ..:%^I}b��D�>��q��7k������c6�!��cϧ�k&�����F���0×oorQ���+ny���V32K�K�?�s�Ta����T�41�@pSZD���g�Ϩ��I4,Q8!FT7���Rq�vQ���R��XY9��N/}?n�.-*b,j˜e^�?.�� d��SN��9�8I̚t�}��2��1W���	�=���������0����Va�e�}.F�P�zv�t�4���yqe���J������"u��#����k��=V��Un^bڡY�(ɋ;�Qbb���E�;6���:�2,Sw��|!���`;mԃѸ}��I��;���>�.z��1�-�w�28w*�~9@U0���8�g�Do��q(u��WOlU������Q#�8�'�c�{�R~�Qc���Z��������d����~��#�>�lP�ڔzs�Zr�w/(pk���%�u�lN�nY�b4}c�42/ӆr�ϳ�yb�U�I�Μ���������R�ww��	[��� ��]ZmYrK�bp
��6�*ٷ����j��T��=�|���K��l~�0dp`����{>~>�l7�FH��]\v�3�a��z3>^����FC����qd�nr�1� ��t~�W�جr���(^��w�c�	�7\*f{��A�x�a����nT`֭d�y��w�b,ރ��6�_{	K^fMh���y�@���q�c���t��F<�nU�{8�_�Ͼ�tgyћN��*Z*�uu;������)�+�A��Y�r�tHz�P�o����w��}��3>��a�k׼�1��k����T<�����
/eh��n���YmРO�d����9�Ƙ�7Us�;��a�1'�k��`U�ax��8�
0Q�>�m��r���zr��+a-�w��a�^J��iU��Ҙ 'yA������c��y4�����OY3uZ����6
��J �.��<�A99����LC��bMM�𼚇�yI����_z����8X��+�sac22Va�ǽ��Ӌ��u0�E_&�&Wt�����&��f6aRyǼj�R;DDW�@�.=� �S���85��H��!���[�}�\)w귓.�����\6-�Uot�ܶ!���rd���犲�Y���vpҊ�CX%�7�vJj�C�U���Dһ3t��%ƺ	X7s���(�'i�r�ͣsG�7�{}�S�vz��Z�����4�@�\Of��ǅ|�{�^�{�����lm�B2 `������������{�Z�.�Ʋ:�ԾWH] �LE{�ُeɍa��z=�Ԭ5=����[�`ڸ�1�2���V�r3+�`_ݵ�L��`��\ n��&"��	(����{���m�xE��]Gu�p�lA)��M"J���P(`������\�W���ګȵ���?�p)��यP�d-f��i���W�ԽSC���X��zo�V�\|j�����n����I��ƈ�=snRGH+��V��Xi�,7jɃTf�:�����w�_�P�D�/�HKf��;����9I�zZ�`�V�#0$ʀl���s�s�띊�a�G���ێ�G�)���U��AC���y����Z8����������"���͓xߝiiH����N7INF|�5 ��;h��!A�!|ű(g�R�v�4^2]������=*A~z �9Vz^��q�L�( >��J�*����9�3M����ݝW��bj�����r��:�^Ҡ�Z�!+�^�+��^����^ڡ�x���u��mS1����õeA�?D�"�MN���[Xzs���;d]�/'�%d�y�!��fj�<��Aqk�u�w$�Kv�oCk��L�;k���Xt</nV>��}�C��[�;*�:��!�Y�E�gh���a���??}��w������co�@��~�������g�`о�tT�N�>�v��1�ݬBh��a!%:E�j��ٱ�S��z���TGd_��Qlr
x*�'�w�͏yVl,Oal\�e
��KmDS��q�G���{裒v/�H�3����["U����S�]�_��Dϧ7�vCv7�&�.W����u�nZv�"x{� XˣR��������u�S�/�����Gph�_(�璹{��M��-��V3�\�̭#2��N��Pc"a�&��/F?dĪ��a�<X']�~O�E�w�D��`�V�J��vٱ��{�p��<2p�wU�o��	c����*W��B�$v�/����{�*�n^�Mt�.��K=�xE�fu�S�꫇�Dg����$j��K�=>iD/E�d-.������Ѷ�������;$\�y�J�K��b��S�=6\�1L:�غ�N8�����`�<�e��^�����i�K9�]}�tw����D�P���P��+�zw��R�[�y�&����YC�+��d��'>�,Z�����'ϑ�{,�!WW,[#*��������ʜ?ne������T��cNpmz�� ��*�O����h�B�и`��g^���݃Wچjy�4թ����RA\��D�b���j0U�!N�]}��ɺ�}7���?���C��"l �_G}}89�
N������#0$ʩ!�wO�ӯ��h^��w!��;�?Su�e-��B�[�45��N=6c��*2�{���N�)˖Hv���F d	V�@�ȫ����Ǻ#ڶ7��~�X��[3�1�`�1�le��:��u|���_+87�v;|�;3�jM��
�v/h��y��x'�B3����(g|3$Dd��/������}��u���OC�TC�&s�gzb����*����9�T���z�"���9&������g�FUM�"D�����.٬X��Ӏ�*�'�Ї��՚��G�&�>J�X�j��[�Xk�����]��TJ{YѲZ�C�#Dc����j�H���|4���@�(�a�aG��fD��\W��+3����ܐ���و�j�!����~"H޼�س4��f};ڡ��X&�����ƃ�w������צ�߇s�q-�q��O�sʠ`�Uf{����Ǝ9u��l�t�K�ٚ�CoE\�.�bH����g���a�)U�s�6��.�SSr�=�4����__jP�B�&�]�����-��U��O#ڢ�:��}�� �nn#�nX8?'�
ӧk��F=����>�Sw:vWdW���G�ޅ${)��Zp�ʓZ��}{�PǪ�)�˄���Ƶ�S��-�s.L�%�^����f+�|}w��ߣm�C����o��+�������'1�\&(�{�5L�&C.0��#<"��dvń/��I�z��s��ϙ�ԟ��$]��ygmd�z��i��"x�Dd��È��)��?T��#���C+�0�bA�,���:�U��og35z����O�t}*����������X��'k�ɀ� L0�_	�T����؉܂}��k����c���1���N�	�9��%'�E�j�o˭�DW��W���O��]y���`N��C�����f��>�����O��w#!�l���&�HTfc�)��z1<��b���u�a�W{�������Q���p�+�(w[r�5�Y7n���b9ő��M�>�]z׻�{S�6��A���1�(O@����1����:s�s�)�j\�r�xw=G7ow��±~��t��_����>���~����ڠA�v
a8蟑Ⱦ>�(gy=8�9�q:vC��Os�ikdk����Aގk�4x�ϸ�$l2�aXk�T�g�h_]z����pe�]y��[=��#���E�n�����8�t�=����*�bү�
,=�բ-��=��g���U�����$���' �Go� G&=һ7�Gw�뎶����3ͥ��&�S����0��׎�eŷ@��=��vyu�6�C�SL	󹶥j������H=WBe�9j�������F��$jm>��ϫ������wמ�`�~�dq�c�?���:���q���GRǗ�엽���F"���C�TǆO��:o&�i�[���p�x��oOU��S����Z)5n��:	���ޣ�~�M���p٤!��p[�ql��f�n�/��y��*���P�й���G0���g�u8�Q�,9�ł�S�=���7���Q�E���A�5~T��"(4�q�L�ۜ�����׃NO�"�W������HA�~�T�����ϲ�<�R.���!t|�k�"���M�ub�E�G��*��)9t�d�ۛ��x��s�U[�ڰZ�r3+�c��)�*��^�W�'u���v��܉���@?�����}��,w\=�A�y`�)�B�J�I�grj�-+��j;��v���cP��L?�|=,񰂒�\2�j/��m�J�5-�4:/Z���)��[��N6.���$�$��Gt�J�'�4\�ybׂ�p	[o����m�emO�?E�����Y�Wy�K1��T�&#,�4A�ɀ\i!��ZgK��1b�^��I܈����.;�=�w����g��o�ݣ�r��]'��R'9��S�.+X;K|i�z��qORxdd�NWu���㋝N�>��UAk�ѵ�LzQ��U�H��"oA�"���ޠ�m��
�����у���H�V��%�����U���>�y��/eaMﯙ��u_C�o�o��i|�
��A�:y��(y~>���G����k�=^�hN�`��s��O��jx[;����|G�}bH��Xx�6'�CS�����zT!�.�J��^�~7�@~.A^l���_|��?������J�b�R���>R]��'����Ȏ�!\�K(��	1�oި� ��@)U���W�'�����
��M*�z�qȜ�{�OW�S��%���l#,�d��>��D.�p+۲;�
�A���8�ea6�}/6b�q��}�x��"!�hL����ΏyV����bl�z����מ�������K��f���c+�\�ʖyz
X] *�$+��qy�T�WV\����iz����$�[��>}^d��_k�!���L��'�y�ˣR�7�qQA�vb�����\�%�w���1�0���s�]GG���p�8dcD8??c}���'��QT�z�롩H,d���-�-�<�~��t=���~b/��}�W0\=��/v�8.�#'�rX��Q@����=$~H��~���{O�� ��]�`��ץ���yz/P��g2�:�?n��k��R���o�;�(���ԓJ�fډ�X��t�%�P��\pS�נ�r�[-_iі��v��ܑ��&��:;Q�Ў���˺A�w-���P�h��4�Z�]t�Զ�a�������fm��\?oޢ0�+�n�����)^6�f@Ge��颳���7-r+݆V{>A�*؂lZ���Z���7w����p��B�#�Xm���I��aEwG��|+�q�kf@kB+�:���$�N]�$O��y����cf�d��ʎ�R8�u��(���,��c['F����N�rWp�O^�vf<�\�Yw�E]$<f�J�rMЉ,�Y�'��i��}|�6.0��"|hs�ABw�2�
�{�v)/�V�c�� U$4G��ھf��� w���b�"1�[[-�����Τ�[���dt�U�d�%�Ъ�S���_���ə��g�+J`atJ��3��K�.쾔�۸).�߳ɶ����š����1lb����Eʖ�ȫ��FZ��}ݢ�A�[5˳�Zpu�=�v��T��e�nt*'0A�0��b֍�kj���ѹ�y K�5��L��L*5��n��y�vh�*\���|�z�wb�4Y*l+St�kqYJ�t(�.�*[�n(�2�p���L'pT��j�a�:�굍�usp
�Y>x��C[�Ոѷ-vse���PEs0���r�Mj�ui|ʕV�j��dvk;>_X)�XN_u�6���[�n���$Nu��; ��P�p����F�y�z�x�!7��]�ۍ�(��a�,k(9W^�1�v����@�q�I����7(���R�6�AR��d�5�hK]|M��`����C(⡍���9 �rU.���K�6E��/y�Kq�쥗�q��z't���Ew�l��CtK��T�~f&s+y\�!�]�q}7�
�7�j»�Y�&�8-p���q�Pc0`�fwh��W����(V<�YiD�	�&�x8(��B���b���|wJ�[���*��u���u�p���*��|;r�8TZk���"M}�.K�ƿ����֧Vm�V��S;�>���8w�ty2�s��^ru}��ם�6�.�+�7{����]\П��]�~��7��R۵�/G�f-��P�ON�]�g��.NVủ�!��ZK6r�[�僯��"T��N\�6Z$2�Uf>(l��_	�����ge�ï�FU�ұK�\
B�[��5���K�O-�=+xm�ѳ;�Yn�Zw�V���@���M�P.�N���k��dJW͉��V��F��^v�u����;w��d�֢﵃us22��\�6S]�y�$ԕ����2�Qj�u4�^q�v�9}���Q��V<+yL<sJ�G����Z�60�����#�S_Ab��2�M�ꝳ�z�:k`1��V_b�1�}�#(]�R�ڜ�~�4� �����7Lo#�ww]�z�Rr�D��C2��%QӚs*����>^9�{D�M�v�����!�����	{�l�-+ZhXh��*�R̒J3HQ#
��+��a�J�ڭ+8[�<=��g�U\zr�Br��.�W���\�	L��/�&�I��;���pUD�ݭ�t��<� �(�m�^���$3HS�(��L�+):Bwu�S�C��u�zrs�
T.�
#2rp���Iʼ��t4I:�=�s��t�@����9T�6�����C�v]��p"��"f���:�VY�y�yay��.x��8W�V|���E�(��:���q+�(�X�Wg��T����,�^{��)�ݐsP��ͻ�'#W��Щ�Fi�t�:�Z��\D
	9UQ]/1ޮ<���N$���8�U�D�$�/;�T�q��2���EJBnBᷜǉۋ"4��]�P��'�G�a721z�/�q�(lKPb�Ds����g���+���%Ԗ�`�k�֤aUs���/d|��y1�����www�]w����&�����������+�fɑ�1�dJ��PB�j?X�n^«��莣a�d��}^��N;�
���t�j�a��B�TF�S��O�iD/DطAiu7�E�g�I�{��T�inR��rV�
2�N8�G�H�qT�����$I�:�ر\+C�Ϭ�p���x/F+w>�ٓ�e���w��R��z��x�Ct���9�v<Ȓ
�@��Bq�!hY~z�S[ٛ�^_����qkmקZ7�=�x��L����s�wK���$M�L-�ދ��}��ڮ��wkI���r$��͘���{��[���%9s��=ۈ��U�%�[�V�xL}�������h4
г��cNīF3d�o^Bϩ2�`s\gq+��$r���;��OV?y�#���Tx�ݫc�Ј?ph0&�(�7��yC;�3$Dd��|v����s2�v!Jg����^BG��;�lG�F~`�t=��9�$�@X�5\o<�w����q��8�y+5�WO�PKͯ!'��,sFb~わ��%�w���A��1?1k�}*��;����3����O�b��IY��7��S�R+���]J�m����-�1��Je���/�}�ݐ3�-�'}�X��N���"weu�qބ9=Q�7� ��`�S�cx�*Ԩ29����fҭƷ"U�0֜1ÕNͫr�N�{m�������y���子	{��J�z=�W_�t��7^y�� �/3cL�Q8f
��yC�Xv��"�uǕEn���yJ��dب�=�Y�و�j�!�����X�o����O���z�O����a@��о�sL����+��d�q{��b\n|��5e�U�7y�\��A��>��뜇�X��+��d��P��B�A�X���Z�A�z�r
Upܶ�LB/��ܣfY����.���lz�P���y)�ap��mŊ@��'����˽��sDn����j�8�Kz������E|��c�ڤ^�����#{��C|1i�;ZvOV�i�U���4�5��!+v���.SB^�~��U�,�r���0�@S#}�9_��onl�d���6�x��{�󪅒��/�c�z!�!)��c�V`U����_��	�{Zw��A=�̭��������4*�\<���َ��=_�|e�N���1	œQ���̚^8��n�&�1���T��)������<��A�x�#�v3�����Zɿ4��)���fDdVe��>����s�<�_J�Y>�I~����!����٭`��9��C���lBj��3.iYO7�Y8r�b�Ե��̚��̛�,��<'[M�og�h��AmN�Q�p�aǑ���a�$HL��Gf�,3{~�^��W�^�~O�������~��"0~~xJ����~���B!�L�+�z�D���8�(��Ө�����Nȉ�OV�PrVj�=�{~j
��Wת��Oh��t�G>B������/����<f�?!c0h��o%\�����Z�#���}�bC�sbi�|$��ÍB�T4Wp~^'ͽ�@⾻r^����_r��(lf���=��q4�fQ5�$w`U��f��A=�J�gԒ��w�h�#�C�$)[�쪌���v~B�����1�z�z�p��L�T���s<CX��c��w+�-��BI`�&Gp����g����^��[mrby7^b:����R��uAK<��pT�AWMFzШ:g�>%C����l�9��x����
����G{��{~���=[{~��?m�/v��<��I�Wd�4�T�2�D�á�&�����Svߡ�/��:�EF�%'�L�J��m���ڱ��X�sZ �1�8�{q��delJG��b+a������*�km�S�=�hŎ�ѐ�:�6h�Yu�}�M8܃�W^CW�b�{qQ�~�y^��N��6�(+:m������q�Y�Be�x���T+���Īݎ�T�����T-h�zQam$0���v��{�a�I��z��Z��ьrˬ�z���jx
��Ǥ�������n��Y�>=s[�>�1s��D�[Y!�������߯��~�l��o��m�����߯��XN&3�G����ީ�#���,w\=�	���\��!`��6�(���}=s�oKe[J~�����a� q������Z�ô�rZ�Kjhty�K����8�C����
h^�a?��sdU8�����0�{��h�Y�:AX��J߭��uT����m��t��&߬���p��<�He�ѳ �q���q"cx����C�^��#U#����[�//iiH���*8FkW�K;�;�ic�AWځx-=���P�~>������.���}���oQ�`/�;B�V��:Jr�R85��S�e_ʄ	�_Dm�Qժ	��'�}0[���v}��y�Dw�m@�%��N:�e�n�'u
<��A+���u}�\
�>�T|t���cIbG�:@�)e�~��ˡ�1a{J�BUja*�[>��3���3
]�Ɔ��hԽ۹���{��*��$���������������7}�j��#�Y���*��ք��F�O]�0C�t���F��SEGxbX�&XU�,��nt��NFw��p�q���p�c��������4<�OL��1�y�}(�m����hse���.)��`��s$�		���U.����*�c���vM�O8RB�Z�f�7x.�&�ݸN�l�FFc=CV8��������v�3�\Y��fN	�!����E.��:��V5c�ϡ��}UU�`D��}?~��}}�~wĿ>�>�.G�&4�s�>� �Բ��l�E�����.��Ȑ����˿��)<���Ϋ��?���e�k����T�2� �	��$�� ^]G�q,K�B����yA�i���!�1R�я<���Nzcc�X��%a�Ƭ[���f׾��3Q�Vl]x�����E�U�OF���D�'D鋠�?v������Ay�p�[��7j�����3�b�f��Fei/<}�n��Eب�Q*#b�%�x,�-��಻�H̙�=b9Ltu-�M��(&,X�c%��KQ���.����m��z*è���@}=r�//E�eiu;$�d@b���e��������Y��qq�d*FT&DzhH�9���\)�6.�~�s&]�$�yz�w^�=ϸ�#�nvN�\��������;� ���Ϗ�� �Ƞ�����)���c�#�=>ϙ������F`�ʩ!�wK8�$=��%NH��P���c�����w7�ק��rC��_@�Õ��x8�w��~��T�a��ڂ�n#�u;��doQ�b;޻~��<$����dٹ�[&��H2#,a窮����"�c����	����A嵰הimxv8���k��_i��>���i�3�B�Ǵ�u�|4>�{���ؘ��J�����U��o@��$�)L܏�8Z��_�����|A�>W2�{��1�@�t G�:��
Jo�c�V�e�e��:�.~q������pǓ�xHg�H>�gf'JJ}}u���yD[P�#�����!�|hg�3��x��/�t�ٕV��e�7�=y���� �7n�T~��p��#:���!��SU����՝�݃1`-n	��U�r�#����|9�bHm���1j|2~��S���)Eű�������֢�:�\wc�q�i��Μ�|\t�3Db����j�H)��,�*7��W������)���h�y
Ы�`��仺����� ��و�V�3�;�Mi����r�7j��u޽���V�	'C�u���o�xg֏�7�_����8�|��5e�[�����&Wy]�0�<�骳�QZj,�?XS߾���;x�
߶#��!+:��:&�(���V�g�|�mFd������.2g��h9�����
�zf��n��p��q��o�۪*��u�gԼ�z*�I�*��`R�z������E�;gȽ?`C�h��[��V|S�F8��%�S�A�h#coę��K�](�}�	kEaցԧsdc�ҡt�s�[xp�陪uh�^�F�.�%���WW���à�����"{�U�[ǖa��q�Z���8���E�*#c{0��L��/ϧ���m�C���1��<�]����ߟ����w����=�R/���r��GX,���Wx�8�;�]�^xC
� e�wUZ��Ď�$��V#�q�4;����u����v�=��՘Y��jw�������辒�N�"��4�ECӓJc4n?lU�|g�܌�$��yg����1V��6�'D�YԳ����F�������3痑 �ܡ1ܺj=�n�g�wg�tb�!�Es-�Kˁ����S�n���g�Pt��`�F0�>�GNxnw�<�E�C(�ߩ�ճ~7�����q����K���Ο>����#܈/���
�}�|��~Z��z�� ж��o׾��3���D���!(j�ؠ�����tQq�Ɓ!iPp���#pgfq�k;��>�3c��|;����V��7t�y��q:�;�f���˝U&�i����Φ0� �F��]i��d�����#DwZS��!�<��V߂�*U}>w�ʾQ�Xf��}��kC�v���Hi�n|	����z����G���N�5�Yt܈���&I)S��v��F�-���o�I-}o���H�WR�����)�K�t ���5���<ۻ����}�߸�<���,h0@��:6B��W�*M�b�:Q!�7bX]��im-�0�s��ÁVk�(oi����?�� �A�1��q���?{U�I�^G6�D�蹓�P��M��@�zv�'�o��D����ĥ�ղib�_��gpLl����.	�蒫�v�ʔFP��@�.3#��c���}A̕jn����z��xe+b���x5��K�`��/`�5�B�b�*���G��N��2,���%��C��A�ɂ����:\5/�Un[j�t�)��p6ϡ8{[FNm��Ywn����>`�+"��^/�HB=�0�_j��ŗaPp���'��!tDU��F���8MNe\���{%��T	����hW89��a'�T.Z�E��nKTa�w��0��ܴD7"	���z��F1��c����8���ѣ�}�5���P�3���`GH+��K:#'ޜ��&�T����\}m�8p^��	ۇ��P<��E}�F��ʀ\l�����:���z�H�'L��+��̏V:�~b���*��~�O�|\��/�@��� �P �=��tN�Y��O��`ďlw`������gH�֥�ѩ���q�r_��	�c�K�>�$8jw��L���������:��c��Q����o�g�$�Tt��T���E�Q����wC��/U���|ǽ���'��ԓ�3�kŜ\Y�����J��q[R: ��\v��C��7�o5���
:-�N�[��'���Κ�q��.�w�?X?B`Gcm�������������������=�N$\	^�~��;�@�+͐����^�q���}C�-W]yJ��W���/1O�1�JpN �r���q�ཥ@JiLy+�^�ag9��SH�����14��<¨�rA�g&�h �]��Z��.LQ�����
��1��>��H��Ud�]J�=����V����c�C��h��B ��&جRn�s���NFM߲:�&�v��ʉ��wG]�ӛ;�j
���ya��H�K<\j>E�9at@�D/^flM��[�
�M_���iK�8ꧢ��Q迻\������C� �L��${���&��Q�f潤ԉӡMzw]�PȺȿ�пLu����"y�q�Pp���� ��3 ]{�S�U���rq��D�t�?��F���q�߀�A��?p��s�g��!U�y�v�8Kc��ĺiګ͈���S¹�>�W
6J�Ad�`�Dpg~ۄ8H��}#ve���p��c�r��e�S>�m(98��)�8:��{�U)�}��!#�E��=7��!�-�T���p�Ӟ;��tp�ò��e)�S�*!a6f�v����.�L�g�`�rR�YR���� paW��%\���y���B\ڄ�����R-�*5�+�ƒ-�=��h�)�KfZ�S~N�����4�q\rpӘ%u���6�"���=�ss�����G��������k����5S��;>����/DugZ3U#*�"=>�90�#�b��
W��I�G��Wz{s�||������ ��U ���'c������<Nǃ"H+q�}���қ��������2`�C6zZ��
��W&UK��PxGt��7��9"Oc�q>h��q��g8v�,Hb�8bW�/��|lǞq*2l�	u�5�5�jM:sу�^{�q(��jDj��u�<q�yҨ��D#��P�;����V#g�}5�9q�����֝.x�gjW'�E��ɏ�E�m��ߧ��T �q8�x�(��Y��b�V`Bi�YI���=���]��-l����$�����F�*a_�W2�(xN�V�ؽ0*�k�M
�2K���d�߄~DB>���)lO6(1|׌Hわ�1/#��
atL5y�}[�.��G]�����.��K���Awy���].o���yf�i��⠽�x��^���'�e�K�,H^��1dOޝ���&���m�G�w��؆@�yǿ{�U_����:��_�l��!�2Y�Q�o Og�:��J¥����qup���j���֨���rVF��8ZՅ�}�X̜iGf_E�m|�
X�+Ⱥ��Y�)8��)`R�eS88��VdF|��7����\�;;��7	"�C�P�Ի�(\�V�t]%����kw{0��,�Z�N�.7LN��Pt�T��_M���P�X�����s����m�sX��t�Fq�VV�J*y��"���سLnc;�ڕ���Ǭ����<p�L�4�L�ؕf��^����1����obze
U�����	���e]z�`����;kZ����sR:���]��3�b����}u���������:�;�f#�ƫ�T�Q�
�Ea��5$������W	钺GB�[�ҡ�J���</q�i�ꉅoz�s�0�aՆB��5�3���UV4K��6��yJ�X���T�m6s_+��w�"�:1�����_�X��=�BZ"[�۽+���wX죗��L;E�'�iVԼ�RӲ��WQ[������]��SoU�Q�j����}��=�ѻ�w��ܩ�Ji��"2&n+�%��%=�r�U$��r�W>��k�&���Q�U�4M4w0��T]M�v��ךhw��~Fm��G��VR�Y~4�:t�<�f���ǹkC܌X��S���A.���R�d�e�Q��L�M빔��L���<❯��4s�0���R��c���Z���x���/��c���%V��"��m3�9�2j�y)�X-���߉�K��b�y$�q�CWX��ʇy�û
�6e��ft�*q��7-���˧��i|rk1V�s����;01�+Ff��ԵӆʘzL;Ɲ�u������}
�gڅki��+���X�Ų��E���ꐎ�v��%�ri���-�˕qM�
E���)Ml�C$�˗���y��N[ʸEވ=i�f��*�E����������Nnt(VTmR��6��,5/�7k"������}�/b�w v0�=��%�yf7�u2�V1�����O
}1��×�^�M�y��Γ�Q��4�))��ͭ�y�a��Pdc��7�z7���z���\�Τ��5�B�N�¢ SX�ӫk�i��[��x[׏�b!�Vn޺�幇�Y����q:f;���Zn�6+ �:�ͩ�w�D���*��Eo�r8���֭5�d��R3��h�s4�'-�w�%�r�-	�'u/����V�Sss*QqY���q�Qsn���Uw��o]�0���֊�Ӯ8�P�õ�YtΊ��ŕ��`����\42a�xB	���YB;��.n��%W��4��v��Qݕu��-FE��O�� !ϻ&��WS�j�;|�����J��Z.��&���k��3}{!Ae^>
0.�ꗱ�����-�.�Iq��Au9�\}Z��+�o^.�O�&���e� �D��j�e
�,#*��܉�R5*4.D�����{=�ڭ}t*�ywy�x>M"T�w�w�"���V�.R�A,AH$�@�
*�h])ϝ��dAE�ZF�薗��!���y�⪛�G%J�HE�vi'@�J"#��U\�v��4
C3e��- �+wrnJa|eUU8�3ΛQ:T�R�Y�V����|�y����"��ռ�yp�R("*9y��^E�)�^]�M2)�<{4�0�hU!s�N_"<�����Eic��1�Of��g�]Љ�%[B����QȤ��ˤ�{U"��bXUS��Db��'0������:�x��R�unWs"��v;��KH�	�H2�)N`�s8E�����E*�K�K5����p��+K�1�'�?O{�������������sw�o�5���E]��^��M�Nh��oC]2p �si����{��]�w����������/�������l$��Zk&^�mN�}�5���D�d`�S�oo�;���?_t��JX�}m�W+��E���WVl��ri�;2Ñ����]�đ���z&�nW����*��q�[@�y�q�8��e�`�읂:r%�EBG'䧌E�%8�TL�]�>o
W5��&���K �[6yK-�G7���xڤ^��!�8�ڸ�V�h�;��J��m��"��E����7�<�����E���s���Oc�u���X�6~�Ex���E��w��������J��rn<�v9Q?
.1���u�6�����s�U��TOz�q籌Tt<�� +��iؤxi�����\�7���x�jl���w:/�RSW�uf;6jq�c��4_��G���d��� �Hup'�o�sȎ$�u:F��B�v*����<�љ<g
����c��ސ����3-}`?L�^�`F0v`�F0�>�GNHZ4�r��2=6��[�kt�0SW���җW׽�4v=��~��F6~�A�_pN:�d%~���[�����~*�E7�-� l�x��X;���xz��KZ��C�Y篅���V�{�n*Y�����R��Zw�7�5a�W0K�٪{�>�w,��ut���%��������H����M�K.�v�I޷��n�g��;#ތ�>� @����]����7�.cӫU����܅�p#��غ��5EAxd�*p!T/�5�CQs�٠�vb����r�F+�R���zFC��GM��EŷE�w��C��L�^�c��P�9������Et����$�!B�K�T�e��n2�X���g��J��9;�b"�c�D�bU>��늕�����8���<J�Й��p$�d5>��{z�ƹlH���g�K�ڹO�V�v��FC����or�9y5����g�I�dU�	�9+0�3��U�i���>7�D�v$:�>����Fk�vB��s�d;�Qk���=V�Aa�R()��-��Q�X��I>6V��[�y�}n:m>���1g���Ax�p�{"�ܽ�؜�w��l��O{�!����B�1"����s_m���:�6hR˦�}/͑U�ٸu��~�u=��V���}�����|�0�%��V�>��B�]E�\=�	����J'�� �w�}�b��*��M�P$`��>��\J<��o�P����ۦ��|bBy�3��츱h�=��cK7c� ��� qbZ/x��q�t�[^��v���^4x�\���Ȁ��__6�6�#
�P�l��|����[1(pG��gW���oi>���c�l�uΑ�TK-�=XڼO�XZ���;�8
x�B�����Й������;����{�������E�B��b�z�[��A�_0C�T��x�r� ��yI�.^��&��q��^�ij<��M�#M��n�"׊�!�LB�F̐n2DxBq�H8�1��Kbm	�R�٠|N�ε�δp������s�:��Ú�ײ�ƨ�}��+P �=*ޏ�MȢ��G-~S�ĳ6�(�#�c[���zR���;/N}�t��;��w���~S�eW<���O��m��[��;ម���T���%��m�E��7
*\M��~��"��B)_���>,mF�?9J��8����b��۳��=Uj`��/k���:�S�O{%�{���r�{�zG��4��Bg�2��p1y\>��D�qxo�ͫ��C+'�q�O��&�P���!�W0�$���y5�bX�&C
������W]�g(4å�;��Ǳ�=/,�7���f.`��ɇ'���4��y^2���YR��10+��r$jqp�?=�1ݑ�}���Ϥ:/���/�_��A�.v��bp��2�D���ܺ5*�`�Poy�M�/fh�k�������u(���("P#�Pg�2TW���yt�]��P�dK�=���ak����5��=���T�s�;�d�vv�F���J�1�˪�W�U�P{��D3y7�<K�YR���Ը�.���R�����)o�?�����<�4𹉡&p���Ɓ3U�n��=
y��R�ᡏ�.p2��������|��k��}�ݿd=�����5���~�%�aذ6����;�S�Ъ��lz;��Y p`�>.�\yn��d՟}�,�>l� �fQlN��9?v؛�~�L�_�������ejF�kg\u\s��GQ�@M�:gH�y&s��)�.BNӲxG�^O����r�7�ݕgv���M�P�j^��0��ј�Q#�.3�è��=��964�����ᙞ͟v@y�����Ak��E�w뗊��F7J�'c�2$��A�G:$�-J��>�[����p'aE��z�Եu�/�����<�|�n����~v�酶JK��9s���1]�-a8`5��rUǟ��#&2;g`��}8�%9s-鍣{3\C��p�ˈE�@�}b�j�o��h�Y��{5���~�r�^p�/�ڹ������&~,Oْ�#��A��B ���(`O��g��ڍdt�V�L{�/���ŗ$a�h{� ���Nsw��
��rIuQ��cB�j�mG�����N�����-����k���-�)��GmS���8�V��N�T,T,,��>�;���Y��s�5�0�$<X�6����hv����*#�M�1Z��;�s�̫ۖ����$���|���k��O�ݕ�+�!W֬E��ʏ�;( v
�V:�f��%@��'T��ᮉ����h��]{�篥j���Z��V!!���HJ�ؐǾё��ڳ�J#���Y�^�~�z�w�o�!�(zt��9��N-\G�ǽ��QgZ��O`�j�M��R�:
�w�^b�t�~3
�bxjq>���Z	�����Ǜw��V�3��y����A�ꂓ���Щ[�Ma����<J�
�|g뛟������}8����Ÿ����~Ĭz���ӵ�p{<�i؃7���U���d䜚Rrve�#s�p�a�$v��T{��]Y��D�9;��{�W�a�V0�}��4�O���󊤶�ǀ�PY�Q5#��W����(3�)�}��g�f�`]�!a����R�f�<��Odz��8�;屟T����Ǐ��]�ʂ��>�Q�:������W�`;mԋŖ�۔ǨZ`k*A�*�>��Fa}.A����z�}4��]���P�#��G��8��O�\c>�TλfGq���%m����.Ͻ`��3c�u�e���u7|T��RC=�zFG��r�����TN��JI��������m��"\���Q��SD�n+�7.ۅ9Z�NT+�m�`h����8�E=Y�؋ ��7��.�b�_g>{Qؾ�_W�~��R��O\��C��0+�rLp:~��ģ������\�6����P��ɩ
ʮ�&a��{��	���g�l��9I0��p`&1�tȩ�<�K���
x�<Rb�c�~��Mﰯyd��f�{����Zɼ����31���e�p;x�F0�3#ٺd�㺉�z�oZ�Q�ul�g�1ǫO�P{�=�y��Ǘ`_X�)��A���+iL���^�F=�6��f6Tn�i�ΐw~��du����A��{��3���� Uz	�Vr$�zS�v�T��$/NY�J��#�	0�k�ܳ�ܞ��'~Բ�P�J�vP�tf���A

[�7/��J��P��1~֔��χ�#	���}����.�{5`Qȭ>�L�]�H�(X�&C
�!*����@'/���z�Ɲ҃�M������ͤ!�<� ��bw�a�hddi�48��	� d��P�_l���¯�\�Ge��CJ�S��T�XYA�M^���]��~�YR�B!�#'u�w��E��[��/�@�����3x'���Í��>���h��Ļ��cP#�l�3�UO:�K��K���Čg~"��yө��&����z3���޽@�������NS��+Y�G5ڇ�mu%pQ^��f�\�\�]��^����t����#�� ?[Oڟv�i�D�����8��Zz|u1��r�ֈ/.�e�uɩo�Sھ���I�zff��Ҭ-?~��c��{ȿ�nc���j:��-�s��ܼ��#e��:��faoQ���>��Y��t�|���\J<��w�&8D���;�.�T'f3��w)��tG�
up�������tMq�7E@��Z�_\O��d��ڤp���&[�.U��m��wR\�֏���/���s��M
|葞�i��:lj���<#vO.Uiy��ooٷ~��zw�V�=�{�@%m���F��n�9��P,9�����fA�'����9>f��&���X��&3%��=>ϙ�1�Uk�3e@���������-,r�*�9���Xn�߶�~5��?X[�@�P�����q�����"1���Gb��Ӂ�Jr0i�5��<:���Q=�4�d�k�C44)O�P!+�sG�������d����G����N�"���"��Ly���A��ӓ���z�Ь>Ѓ��$�������
YGj�1���7{/� ֱ���t��~@�M�T��ÓM����h��T��PN2\�����6v[%����s.T����ȰP�2@��;�/���^pz%w��l;�Sw�H���{�.H��k9n-{��s�҃��擄����QR��s1/�N! z��a�rU�U*ꮮ���2�v7�.�1���'��E��Y���*la�S��|ef�{&���}�9͉��|*��t�q�Vp�<�$$��15����CҼTv�9	��U�l��=�o�dَ���Mԥ�lwf]=�Yӑ������Sbj*a�������~�l?�#���/��l�Wo���ad���s�נ��7���j�!�xAx+�$�u�	��[�jQ���ݚ��e�����b�~�)���@_LyW�����t<Ÿ�JÆq�<�^��V���L�W���0�_b����952&0pu�nE�:D]X��q?!;]�<ŸF8,^u��K���ފ:��x`��α�Z��l��^��#��Ͼl�$��E�o�(pg�p�G���mYq����kj�_ӉU�GU�r�Q�~	���:OH���s��E
�6���}�)e�ղ�#�=}��ڧ�-�ĉ�s���^e�})�c�z�\ǘT����a;�����QXZ��]��h^^�2��R�������V�4G��읮T��g���;� ���W'�^&j��9��&��t�T��k�m��"�0̾��twZ{�z����%_vvM"ek(�LK����0��
խf��	û��Ķ��:�NZڭ��lÛ;���2:jTA&�>���P�]��<9�B�t��D�춠zr���ElS�w73�ÆՑ���@� 9ڦ���_�E}�Ztح��]���?���x�}��&UI{]��|���u�mTٝ�N��m�%e�����
zP!`t��R%�x�1�q*2l�]O��7rE�M��M��>�.2�[qn���{R��:���AC�P_��$O�W�"�}��sD�41���K��T�Z�T�=�į���W}.ˈR
�0��B"~�>2��0ݝ��Qv"���ڿc[�=�6K�Du��S�*�В����ʏּ(�;EL%52~b\�5�*(v�ᾞ�̐�SS�i�^�"!X���u%*lI�sW1�)�������%ŴC�M˙=����uPٿ�����=�O���=��ƛ�w<ɣ�j'���T��ٵ6��W����/,�3ED�3�p��G'鹺+~&��Gm�Am��f�bU�����̗Hכ'jѓ��8��i����0��9?�8���4�/�W����_�H�Ȝ^����$���<��{9:9�9[�B��.s�U��xm{g6iNG�X�+l)���2��a��m8��s�"0Pލ�ȕ��-S��i�_wWe��_ƉY�U�M�rM "5't�^��}6�7�u�f�%Am=�ˌ��H��&!r?�;�IF��n��L8/.J�d�����3y��4��+��L��a������U��ki��Y���>�������:Ǉ�[���L90��7-���A�\f
���B��Rc&h)9_A��r}��~rf ����(1�� uK-�<��Odz��8���=v���͍�\VT2^���o�kK��,uD�]�ύ��\�v��H���s���Lu|5��ǰZ�ɛ�w�sWd���� *��A�ǂq����{N�uBo�s�K���(s}��7�5^�c�j��;g���;?@W��l�P�SM}���mn?lVK��,�M<=�Pj��כY/�e����<���l���)&+�1�7Ma�Q�2'KH{��9�d����>��Vm3��6��	���Q�R3v���7qF�$z�^�½C�n7S���W�w������Gy�xSe8F�����W׼��B��?_�ELwL������u	��e�^��D9�dVC�=���)������|B��G��flP~��q�˃��g�1����o}�<1�2�	����)�������2;ڈ��VT�+�Q��kC�~��f�tĬ;�m��_�#HF&1#��&��9�Zu"Xt:C�΅��^�T�zX#�J�E��܏��-�D\���l��[ۃ[}��4k�H���A���Is�욗q�6�#z=������n�X���;:�Y]f�
8j�v�H�bc�Nȡ�Y�� �Co�Th�Λ(���z�&p��+�tn«TU(>���V^�|�s��WS�V�̕fR7źj����W[������W��;GN+���C�Nl�z)�ߕ.6�S-]r�N�הfv�V)���AnRޑ�Zr��K+so�rn���GG�IY�94���쾤V�-ւ��&V~Ͱ��'�q�	�-ŷ5��j�ne-*u����Q<n���8m<��l��Lv(�y�
��YBn��13�x�$��t5�V��q����`hqS�2��HJ��E��ֻLZV�j,��8�;��d�4��L�I�	�IE};��z�X��v���vUo'�IS���<;S5�6t@]��d�����b����K�C��e^���U��b��p�v�H���jL��9���2M2�mYC{�R��X1d�L���i�9��S�}���U�h���_@]<;xؼ��Oq�q�D�-��:�vo !/r)H�ڈ�0*��}�]u��#>$��pvof��M{�����R��r4��/v=-�9�!�r)��롑��^���{�yfS�x��eں�p�ڏ.���8��SEiy��I����	�S��D��h.[p�t3#��%����s�Q�4S���>d"�f|6�Y';�b��SP��lt��xmoYJ80�آ��{9*��}�]�s&��j�JJ�w�^�ו��D�Rq|�V:������3��E��3R��h!&�j�Gv�q�g\q%O8��&���
�Bޫ��J���.]���u-ȷn�^��Ms&Y[��\"c].pDC��ޜf�Sf)��h��90\��F�m>�%�0��S.�'�O��-�Lf�w����+�{Ft��]-�vBai�`�=�eD�.� ��M��9�EeWrv���hq7=[�WVP4��ŉ�T�tL��|}�ߟp�����U���7���2f_Jj��zӾ� G>9�Tr�4��i��5͡s�^�n���f��ǔ��V(����כ��E�>u��O��&+0���_?�׮�<�B�U.�W�u�m�W9ƾ�J�J�*�9d�nTw��,�<Z��$2
�y��{+�����z���5���RQ��vgM��oMb�ݰ��͗F9�M��r���t������Y�j.$:s<���U6�2�5��p���y�9�o+�.`,�K9��hr�)�ݸ�Gc_#����4���S�1Е���$7�ڙ��]+h8�k$�i�.m�gnl.����R�T753dv9��:����qC��e\��.�S�%�-a	�NN�Vt=Һa� �y|����\�Ѐ����UH
�
l9��s���H ��B��E$0�da$E
��:�Z�:(���G��=��b"����I�fj�ӯ.EC��z�I<�:�E�κ&rYaT$��Y�g����>�"�L�3A9'J��=�=)OuڕfU�4�1T8RZzS�;��I�J9wfETJ�(�^����+���Ŭr�^t=7��]�q�
%��|�<��g%�����R@�r,��j�����K3�w�������3��=B�؏:�E#����<P�p�J�"+R���D.Q�WCRO���Nl�"%wiTI��h,�2��X�J�"�D��q(�I���B5]s�K�Tf�wO$µ/8��x��u�/��KT���,K��Ћ��[����u/��W	����^\��\*�R.�%D9˗�4�77!H(/t�f� ��Q�
>2�q�
�TK����>&��G3�Wb�2p9A:ԗ�+�Y��O"����K�׽��<%j�9&̜D���\�t�#�鉕��h��'�̍ӫe{$H�L��!��@����i�Z��K�G�<¬>f�~�J�B������|�;oc�+��Ỉ�	����z�|jV�զ���:���܌g�r)�3Ew�G�V9	��BUMC�cީ����K�?��%�aP%���3��Ԟ?P������#�*�V�m
��ē����Mϸ���r��ǂ_�4O�՝�ٝ���(�x/�r;��;��a�{Bᐚ>�!X���ω��G(DAW]!��|�7��x*�C?E���0�i���b���y�^2\>�ؑq����>J|�I^��x�}S휉b�t}_r鈯�ُ�&4m������7��:��[�z|3+6u�DT��-��n��P�U��#��0�"�J��?}�sE��u�qe�7>�Eu��#��ڽ|1pK�I�!e+�$L�M@��_0�lX(9�8�AN�]�~�M{�����;=����S�<zc�����}���2A��&a���܋��,�_e�������? ���?Ym���ڄZ��(��8]87x�6$�Y���(j��������� ��ȿ��wYgE݊���]a�aiEW0`���v*-��ap��Nn�U�\]x��-Suvn��E����:j�)i�j�8�ɵ�#���]��"�:ʑ��4����Sq�4�x%r�أ�2�6I�W�{�'�s�>�#� D���?>�?�U��E�=/>GŁU�H�&T����|����0O��Ș��ܲ����؄t%�\	�(�����6:<{Ȍy�xF�jxu��j+����=LI憛���p���2�G��b�[>�#���~����Q���*A^l��zϧ9�����[�ܺ��t!�Ҟ�K��{.�a��L�q���$������K(�}�������閧��ع���{�<�=V�w�$r�����d#��Px�%|�!3�_FY�s�{�N�Y���p�rJY�����4b�X����"���^a�њ��P����B�x�/�On��w�j�޾��$ȇ�C�w�fd��l���M�������4��`e}�.�u�/Ր�x�ɵA�ƝAr@_h9�H
��Zo�Y�ۨ1��2O���< ��l�B�9��e���~�̘�S?�?K��n��4]8���_L~�Cx/�㠁<Ÿ��+��N��|谂�Q�,����bOX皧�8��P�C����	�l"S��k!Vj��0�>���^���wGk��#*/n���X���\�Ć��!����������V̌��uժ�m�w��k�nZ��:�#�D�\��I��Wь��)�����9B�u�bĪf���;2�,�3�]0W2o����;�%/��5=����}�Ͻ��Ǌ�Ϗ`�m_����@q�-�U,���9e3�6L��[�#�>ջ�s�=��Kӹ}�a�nY��Wm�
j������p���#
L��b/�f���X�3��ˋήP/e�#��,[!iu6;h�p3捵.�W���}�Ǥ�a"0���#�%�F�U����a��#*!D𞇼l8D/ib�u �A�g��Cn�#��v�z9��ؘ*�����
���8�P�E���<l�x��//��&UI{]��}\�s�.,X��[k9Qc�]r��� ��!�l��_@��k=>�}v��t�tH�}A���%?R^]~�;�2ή�_2��Ԕ��<��Y��V@��� A5�-�b0���f�!�c^.�wvc��a:���9�3��W��O�E�A���"ah
�G"lxSS
/%NC������ѵ�r-T�K�O����J{*�ВB��Sh^�����iD�d�s؍e�%�n��0�rȐ�֚�x_X�ә���rl�k�1Î
?l�$�~p$5��翱��b�{���V��z˨,���^S�]�ە�D$Μgl���gJ�تZi��w{��C��o�GI�[h`�*><*{��qJ�S�%��W0��ۮ�����>�!؊�Iz�3jC��tg�:΋Y �]YaM����� G�}�*�.ylH0�N�U��W���Ra���zq.�����b(��j '�0�zk�C*v&�b�>��W$��/��Q8fУ�q>���ןV�Iڣ�و�Y'TX�a �ݭ��y��b5��yA���$��6NM2:ǉB�8�+_O��@lE��#U�/'��������:�/�n��n7lC��Ys��~��NN䜚R~�ٚa��*�=]ûhTo�3Y�{{1�xK�c��g����0���mU�A�\d���ӑ.lɛi�gSď>Ǜ��dO���pG nT!���i�T�َa\�_>�a��\d`�����9�������{�j˻v������j"��(��<o�2�s��mԋ�����E�P�P��N��+�N�)D��{�8^�����,_�
����|x'�%h����c�hv9Q=i��GLFk��΋y*�b+����ܑ���`U�#�W};l�p�1N�}p"���;;�K'VKENo������_)����rC~�|͒7Ô���`/��6D�LC;�}��۟�����-�%�NV+���
�����_�xh�;Q�Y�Cf5���7O��ۏFT��ܴűfW;cjۢ�;Ā���.�`�ٕ���6�b0Q�z�̷Q��H��$c�QB/�u�D����у]�W�vb���%�кt����O�h<�bic(����{�Y��m��b�O�̓!�;��ە�Zɼ����7qG�&b=� v�y8��{�zѣ�=�Ov�7�A�,T�JRY����"1���U�~�K���<��.���b�뵓�����i�UU��ͷ`�
�bB9�����D�^-�Z�^@y����ED���n^�]��b1[�ʹ���P����TLf�
�4�W�����q�a{QR��r�EƯq,�FoG�[�gˎ��6t���
�������J��R�.��q�z�g�ͯ]�L%���Ru��q�o�`��!�?sW1��.w��iX3:�!���^CS�sKj,e^��f�]c�Ň�;�ؐT�
e����I�}yd�;�fh`T7ꎕV*=�5��W|�p�=)�~�����a��}��r@{Bᐚ>�<��ǅ�R={am��;m�%�˽��H��"���g,����LC�Jm�CZ �� ǝ����]�ў�ܛ�7��\V�KX
������"��1�1�m8��u8l��,����ᦰ�h0�V�mO3����6��6u<\,�M�xV퐫�%׉1wEj����Co��<���=��G�C�ѧ&�#<(
��S��\�pv����E�kK����vMZ�v���fL99��G���w��s8�΂�QO�Y�kz��8KV��3�:p0�UpBǸb�Hd����#2����ȥ�q�F[NJ���1�6�(~�����E[딶Ϲ�oH���{���M"R�RD�ܚ�~B�V��R��#����dF��z�t��?��j/�ۓ���jZ��֢Ǌ��O��:d�P�!�#�{1�:/�����6{�Ȍ�˛��gH/��J�}7b�l�k��ܩt"by3�w���^�7�{��Ŀ������ZgK��ʭzF`I� ���v���S�'�>�\C�s8^�d����8cR%܈(J�b�ؐ�'���`��
tԼ#k���ܥ&.�uD�Wp�5��>����AX�f�/���}a�-�"���a��@�!y��Oz�W�M�%i�b^�̩c��D_���AuR~S�%*
�h�,�
YGj�1��b�۩x�e��s|����e�ʭL�!zO+��Gi�_r8d�c���B�7��9>��ut�W��=mT�2��=��8n�!4Gu������_5s�+!��eMTW�p����k����#�l�گ��Fd1���v�4�?[���zR�i���n�<dMއw)�a*={�{��؁3b�1��G�k����t�� EٷaD+�fޫ��}��=�nR9��u�(v\+N0O<��Z��L���Iy`�'U�SGi�n1"�*�*�ّ�}����F$��-V��K�y]�3��57Ø[F���>ԏտ����`{�����ӿ.e�.����V���u��0,���u�*��\o�k�{/M�G7A��ک�g]nm�� `G=9����,�9��5��v�/AZ���Į�(N�Ʋ��Ll{X�{~6��3�;F֍Z�-��s�/��ԏ0;f���>��G�A��Q!�<tT�Ǝ��{Y���rW�����g���s�;8�^���[��la˰������-�}�f���ҩ��Y���N�8Y��,?����I��B�����a��e�3�zA�t����cb)��ޓT-9y�jD��'�2�k�vąƕO�*����:�-�𮾎����!r�(/x��{�=lD�Bz+�
�=)
P��YW�%Ԃ��\�ث�р7J\�抓�A�7�����c�W��� /�} �dO	�v��R�#{B���reT���ț��p�u/!%;/��a)Y#=,)�_l�O@Y��%�x��f<��%FC�_~�N4�����XM���&$�eZb�t1��G������[+�1�0�9�e��dGOۆ��x,:�_,N&ė�:�[ڥ��P擮�l�Us�p�;�7�b)��>�m�:l�kX�Ӿ��0�gfbÿoikDRqk���{��W���iS��[=��gz��9JM�O'��Y��{z��P(p[�@F0���;�3Fr����y˼ՌǞ"��mߜs�ɬ	���A]��ʰD¿��	��3�g������'�F�����������N|�GO�X����S�
��%!!g�Q�����t���Q�/}��6�~�Q'�=ٸ� ��q�?)ٮ5�W�����:@�b�G�ɰ|�A�}&=}W��2�%�y�ʦ����F��/Bq1�ʍ7Y�V^���ˈ�{ڮ"�R��FV�u�=j��^�6j���$�2kN¢���0P��&'��N<�_�`����D��[�²T0���S�nNN}n#^�؆~�y�	�"N����94�}`�聐pKS{{x:�
au�zY�����l.��֓�q+b�˜�9ݪ��O��Q�Pa�.����F	2e�����o��Xv�/}a�+Y莖�%P.[�mY����3��� t�K�FYT{�+rw����~�~�H�8b,#�:�ۉ$��1�2��U���2M��^\EFi�Ip/�Lӛ�sh��:��L��[��5����e�Q
,�yP�s�={���'෯�D֣��TB�y����F!uwk��Q�t�22�^;i��:D͜��3�κ������ϖGw(j�y�9N���*a{1��N(�1"��]\R�d��꦳�;��.uP�OtF�Gk��Q?&�#2V�xd�v۩;�-Nʢ�3=�3���{��Ø��]����|��Y���U_G�*V���.v=ƇݎT�M�f5�M�����X�������Y�I��}7�g�jo�
�t���G����}<�_u
g�ҽ�6� ��z��G?w{b��_�w#!��kt��$oLxb�����.F�؉P���/Np�&s2�^Ϋ�p��v3����5�Y7���������H���A����	Ix�b��oWz��'\�GOt��Q�#��!�\D/?%�{��Z��2ƙ/<=m�D�ݭ��+D�~�4t���!��j�ZֹGSm��M����v�D��]u^]���DC����:45�ݵ��J���3Ҍu{���M��<��[�#����R�+��`ډaU�m�ךR�zG�f:�U����o38M�iL�cˢ��3Ւ��\H���c��B��o-j����[廾�u�]�Js�&u��f��4͢edCT��ދ85��n�]�:`���O, .�˃����P��c���J*��6I�w�Jpl2��R�&���A4��폋���a1f���M<E�����%YĤ�VvG���H�N̻���+�o[aL;���^3/@�ޏ+�{P�{�-i^�@�44��[�ޤ��o���3�V�l�סu�+Y�Y��7C��Gw{5f�|�q!�%���,jֈ�}q�<)[GZ��[K�;�}35�{3�*N�:�����*C��p�!6'*4,�Ɍ��;��v�7T�fd�u���W�]{��qG�I>�c�%�÷p�'>��>�ƪ+�mo���K�~Po4��:=:/	�ɫ���q��v����^=8,���҃�|�x�l�[�>Y��<�|��nl=�ޭ/g�}شd_���(f�ձEJ������0hvK����tv�HZ����7��.�w�
��|�~����Q��w������̫%v�����t�v�G�w�������{�3m*8&fpћ�o�o�'�<7;̇O|��o�GLQ������p�;�4"�%���Ui1B�n��KV��\i`��d�j��~�RMh�|V�q�����+}�hp�or��S�D҆%8�ս�v�y�T�Ap��ls�B���B�k�8-a+�\n�Z�+�\٭"�0� ������Hs�C6�Z�5��c6�\t.#�F��u#m^ږor][�t	�I��<���hܼS��W��v�c7����r���#j"�Vsy���W�Vɭ��],uu�9vbk,�{���ft�t�O�c�Ӫ�<i[U,͘2%�u���#mu�5���Ib^eb���h��8��tS��rG��b5�U�����X#Et̬�7N"^R)@�[���u�R�����RN��:��{�Ʃ+%�˫xmFFF'}��R6A���ƞ0���GI�+/ۼ\ڒٝ2'�V��:[Ϡ��gG��Tj􌴕�x�1u�9�S/n-ӴDQӴNP��:��<!~yg6���#��D��V����)���<y�l�y�0�ռ�L,]v9�>��<ol�{�gWC��+�9\�Y&�{6��Z��
A�W�b�͋v�^̚�B �����wwZ��iݢ;�A��ɉe��Wl�w�o\���VZ|��ݯ:;h��\�AF��=w�1M��G����
��j"�b0��iu4bS�ڜ/�$�(it:��V�LY�m�Ƙ�N�������\2NJ�'�.�/p�-��UG�:;�.*YK"[��95�k��+1�ץ_K6�|�xsi*�ơ,^!�"�A�jB�F�b�7oE�I����|�'�L.�l�p�g�����G-��er�]Cb;�KU���q  E�M��hJ�b��c3fi!,���.�������b�Rf�!�2o�m��q�U�U2��s�?v�:Y���G�f���9l�+��-���9�"�q��6��j��E����w8�77����^C����p7%�<&lY�f���5r�9�4v��r�t�!����g�"�`�A�@�3�\�zh^�}�YUb���^N�l���8κpt��d�+���6��y��a��3G(�L�ot)X�ZݼYo@��M�B P�86s�F���u�ݠ�:V�.��>Ы�T��{�w�SF*�n�[J^��.V�H�9fɛ�TfZ4����/6#�ӯEk绔�4��(n�v�*���Of$#P]h�!�U���6,�#�g�����^f�a$V�]f]��1�s���3bؕY��,	]<AWڑ$ņ��Z8��z8P1Z5��,��tȴ�ot[W���퉑�}s�(s��zi�#lVSr�E-�o݈6zŗ�Z�N����lT=t�C�;��Kd�@���.���K�4C2j�ɷ�!m��y #9o� 4()�4��U.Ӑ� �"0:�_���T������EV�%��.W8aɩt*�m�GzKx��P�Q孩C��4�I�8��9�˕�Z��q�2��/�'�G�블Uw]Ǟ���'��ED������<a8$�Z��z�%�w�Ǉ���{=�QD}����x|jF^�Q�wyB>J+u�BU�*���-S �;W� ��*�q��{=��#R{,4(���J.IV��P�5Cs�J�sȢ�� ��^�;���YVO&����x�E���=]Јsy��xs)�y�Q]�����:�Wf�|y|Tn����r�x���5�x��܂�\�Qyrr�*���$�$7��ȧ�x��|J���2J5��NF�;��KD���,�R���{���H��ܡ��J��u@�Ϗ]��H��*%#n-�2.W�'
��VtQ2zb����O/#��+��fC��K�q��*����U<��efG¹%QWsJ�9VI���|y��D�jn.�=CbE��Eʢ����Z)�B*�V�:ȵ�bN�K��O;�%�w=��]B��!pJԭ��,Q��/������
��
����޽�{CD�����GTpaf���^')l��l����]������vu�#9ZŐm��;~��Ǻ79R��:�+�,"!W}ࡏl|jw�}�*y�0j���s\ד��T4�Z�d��	
�Uֽ؈X!PU_���w��=ہ�!�9�b�X����-�iR	�9T�����^�0EpQ'�Gsl�����v�(3o�����ջ�M�䅋M�y�R�.���=W�vL���������z�c�|1?����������bl��P�s���d��t����k���F>�Y}q8�0'_N{|@��cͷ����[�����ú,�]�Tp��S��G�������?6kk�H���v9rZB��b�=��|/�|���2���r�U�ϘYA�E6	5�8����뛟_gs�z��`Ba��׾K�t�����ܗ#�wG#l��.���fE�e��Ȼ
+�B=��w[o!So>�Z��=9�.����~���4`踍\��_RК�"��'Uf�ǃi`+�9�M�ڝEb�jVpGv�Ûx�	�-�]W�J�CMG��Ö`��U��W�%��|�@(��CW6���vC��p�����S�5{9>Ofk�sc�a�PY�.�Ku����ü[�w�g-�@�s��x��lSX�ƒl,om|�'��c.te]���=��]�n�q� Bx?X��D/m�����꿏��É!����!S�,eH3:
�s�7#*j#�7�p6k�����>BU���ܬ;�k�#O�������0;���y	�c�~f��1��VU���9�w�-��@O�>)�h��P���=�����u>������v;�F6+#�oWřMq
}x{����+DGW(.n+/lz��[��"!�kض�{�uǯ�.0��)	�l�U�����xȰE�γW�V��aÚ�n��#��o>�@n�tRl[a��=~���6g��YJ�B���w��OLb˯Oߧ\��=�C2x$��g�$��}&��i����B�Q�`z������a���v���a��~��.�p�3q�����휨�;�,#[��_�J���j���_l��v8�*4��I�z�l�5T�K���W^���=�3/F�H��"J�/�Ŵ�����HIY�(Ғ�E��*=U�o+Ww� `�gm��\zԑ�ugz� ��=�&l��3#��x��;s�c���u�q��r�{�����k�3m�Y�~���e��B��d#�q�bl���a��_�3[^�����u����7�eX(lƇ;w���|hL�>�=ċ��1�;<��?X�0�J�-�g�i'��F������
๵����v�ﲟgʸe�4�l!C�uǩ��Ԓ�GwI��1;X�:4����0�&-�������%��W������m�������(�U�ۭH�%���}�b��v}p1�0�(?X��k�l�wT6��л���2����gJ���R/�=����Z��]�@���(yH�2���r�W6q�}�s����ҷ�Oj��?;?7����|����m�����饓��pE⑋,w�@�t
R��s|q�?Zt�����Ezxþ�ޓ�Y�û�~BBu��sα�{QeR|T����q�y�W�֩��,{�ͺ:68kyLv\���\uҶ�sx�)a�z�U�C��VT���e����UK��#Y@Lp�����ٌ�t����C8Vw6�c�-�\L�v�'�s��U�QY�l� nS�ƣWx`�,Z.��4F�{����>0˘*ӫ9���σ`��` �@a���G�X~����qS��ܞ�oD��6�є���$o����xc���<:'CT��~�^op�_��^/�~�5��ui�v�X	|�j�+��f�K
o�:��o�sy�����ؕ��\�w��	�/���E�Y+��
�$M���8����^��OS�vt���[����,�ƌ�1�����X�F����Q��{���p��kt����z���{��E�a5�`�U?LF��\�e����t{�/�h�@���;+,�����k�k��2�>��#WXW�Br��J6f�e�+�h�2�F
�:C.)�~��^��E�����ډ~R�Gԏ�D�^e4^����vܞ�ݡa�le�Zڹ��b�o���7��w�1���ɠ��Y�����4���eX��|b~��ŋ�����;�*~�u#�&��v+��J�ਦt�j�<"��'�>>�n�����yē�S��'G�C�k��)�i�.�|�Ð圵�.���[���M-��T�u|��'���yFI��zr���ΥS�ps�e��suҞ���i$��(���w��^L��n|��{a��o�'�vc##)�晿A��^Ƽ�;���5a�<9�]���oݭ����`��7��zn���q^���ᭉ�[z��΁=�%B�	o��̫%]������u~i���,=�j��&�+�`{`p�}��&��Z��Ȳ=������p�/�(��%yg����������Ԉ�_w�
)�uH֤p�_rZ��序�;M��f���\+o�u{���X!PU�D�����~�X_w��W(榮~����q�~��╡i�ʦ���yd���=��!ԕ�=���Α��+)�욷�;�W۸��rA6Ǉ5��Ҟ�Z"�u��[�c������ħ�^����볧���~�bl�D%�88�ՙ��0y^-�:'?\�9x���;�_PmZ��T�Κ3V�x�C���7���z���A�7�y^�Z#��q��I
Z�=��Gv���5B���E�"�W�j�\��gk�K/{�՜�ZV�A�޸����x䩪�X^pym�|�l׺�Z��l�*�|3*��`nN�wop�e��gf���H��ｽ�m9�Ov�l~�݂Q]|�~l��[=��.���)�Y�A^u��p�6�5l�XJ�m��eX�C^���÷�ӗtj���8�f_oH�����-���9��u4�6��H����vr#U�ڍ^��=>�����w��~���jY[ӻ-��lZ�����L��ڕ'P{����[��s��
�o��K�N�9�RO�����y�{E�V)��Ue�xwێEZ����\�BTd��������x�	�Ю��-E�ս���4���c������b�Z�<@��;5�U<��z�Y�9�Q��K��{��}K�򲏼��yd	�@����r���v���-��j)/j9욾�y��+�K_�.|Biw��=w�8t3U�Nd�tZ�,����'P�y����~�*]�}x{�����������<�F�����E<��p���mQ����˨\awn����b�݇D�,6N���J˷��6\YH;u��2�aŏ���'�>� �Y�m�E��+k��ư�eM�z"-���'���Oi��3�VAG�Z-�P���j[�.A��,�)a��b ���-����B�!0��Z��۠�ả����u�BAm��Ţ�U�|�];�ʹ�F{���A�`ְ_ S�>���w����6-�=�I�b�ج�7�w(�
�;ly�ؼz�{���W)]M�y◰���^����]���M��U����;��o��DP:]��2�\`��v.+0�����؁���������4�l=��͍9�+�kb���Z�6�zg{sK#�5�?8mï�OWxF�.�:3���5���y&Υ����ӑ�:<s��׊fvT:��)�v��ƪ
}�E�,vy�N?_��!+m�O��o�K/}��'�ȬGݹ��/���"hw�c2)�~�;Wh�m���!��ڻ�^z==�2Z�bV����W���c������f��vЏ2�ئ����0��o�`�X���;��E���.�b�4bѽ�x���-�wcJ��ι�Ԃi�C7�u��<7����"5� ��8�fX\O#N4�˱�L��>�����z��C�Mt� �N�<���,�oz��2?�z������!SW��YWHT�[����4$�*\�A�!hHZCB�,;{:�2h�i��;�~m���YV���)��j���[�]P5P:{���L�Sõ�f�q��_��H�}V?;-�X}�֪�lo�GV��{�Lu`$������= �]���JV^�;��}�]i�Cy�5Jo-銿Y����z�3����H%�u��E�'��>~ %�z�:����کy��������`n�,�âPj�{W�6����y~��^w�P^7��w���~{��ӥo���!��Q��z���#���\z<]5��U�<q��H������c�^_�FU�D�ª��k�}�6hYo5�웨�K�%ҁrVT��*Q�>�p�����f0F�w�c�3L+Ֆ��=�@�r�Ɣܽ�[m���ÿ�e�O�,f�����
�R�"�oo�km�����C�]�k���/Q^a��;��op��ی��nNY7U�{� �z��ngB4� \���+<S�n5c�B=��_�z,�Onr<#+N���9+om̝o�%i��"�J�ٸ��g�t1 =v<��qG���ok%�����Q�#�eڋ�F�vV9�FzN��o�*�WH�����m]�w ��1Lq�yد�ުRr\_�P=T!-��#C�or5������+�2��ɬ8�����U�Zw�of��f]������)�c�1@l����q���e��g������o��ݞ9NF�#nБ��ű\³X"朕O�M=U���A��+2{���Ou�4��<z�a�xk�{�,Q*�7:�ުFwƆ��:pmkO:�[Vݐ��Y��Ƶ��}:�ZG�9�Zfz�,��=Ȱ�0{�n���jw�h6|:ީ�y����V	���s;oJ�)l����}ޯ���~��j������>|�֌ �K.�����X��+a+�7���c�=|`{`_�{��!5~��=�\����B&m�]�ui����]��-[X:�DB��x(cݒ5���ù7!��v����W�������z��������VT�'���2�R�ú�����e��4�-��ٽ'T�N@�U�4�$R�:��LA�S��v*7��w	b������n������/	};v[�uoq��z�5Ep ��r�ʧ%��ks>���Oi��w����J����ɶ���5
���nh�1��v}�LNmY��B��q���كۭ��7�M�z��P��{�+bc��|��W�َ�G��9N�ɫ}[�U�!7ܐ����O�K�+2}�.k{���he�ɷn��<+�+��	�Y��~��6&�L*<��E^{��g�z������_����e�F���[�e���C4��*�u�{�k��_���7�2�b���fU��a�}������u�V��F��]s�rg�G �����g�k	�{7*�`9�ʓL_Z�s�l�[�9 ��R��X�k��4Du4B\�v�"X��;�:/�P���5Rǖvj�ͅ���į����{9ou��\-�����s��[��>�YF�v�'�Y�Fx��0R��{����	�S(eOs}/�Z�(HؤK+Dh�b�o
9}Uѽ�C�Ϡy�/��y?d�D�@Z��>͌���+�����MR6M^
):�_β�����^t|�F�Be���ň/��.�7�k�V��rS9��E���Z��٫D�P�$���J���溮��yǐ��FQW����!�w����'x�:zG,���Y]Sx���nh��[xV`��]	�gj�s���-�H=��:�8AB��	���a��F����}�*5f�rM�]���D۷7�;.W"{N�T����Wo<�dV�U+(�R���������ݤ%�J�ݔ_5s#F���;'�{����Ȏ�\���9���'5�'t�F��y/m�oNZt:a���sW=��m5���I/E���0sp�ȴ;�!�D���`�9!/�2
u1���6��U����!�ȭ+���ź$K�L���W�T��*�Ŗu.�6���C)Jɾ�nM��Nu�+f1 ��#�J�'�.��3�6����1v��A6ᣃW�pF�uӚWuu)tL2�fg�� ��- QV�}� �����Ŗ�P�gr5Q&y�YK��,ݻ��G��,����FL��k����ֈy/��u� u��YE���C9��:�W��!�iY;ۇ_�)�n��B:�%�����]/��՗��}E�C����:�i,%��B�7	uԛ�j�gb��hJ
`ܝg�@;A3V	Y֟tr�Ci���q9�ն(��ms��H�Ϻ(��,3���������}�}�i��-���,q�O@��gj�v�ӷ�>K�u3%������li�=�lE�s�c���te�˳�(��.>�
�E5�f�_�Lf�a��t�V乥F*Ɯ��s�.��u��#��W�Ne�J��^F��M���ko;_�Pn�kLU�:|��e�nӬq�{�t����o5��3%��˫9GP!ʃ*����hƣ�&;Y0,�j��Ҳ�t�_'�f\9��iȖīQ/��e���,⏨4&�����w|y�iiy�P��Y/s��h��"s��n㓩WN1�{(E��=]���,àD��O�`ͺ��lqJ����VWp���PFu�:���*`�Ir���Q⺭8�a����|�v.Eh��&C�\j��RoXUe�z�����f�eY�d�XsNwy��3g^��+*��A�������-l��4W.ӓv��������֍�;V���+�V�N-G�����Q�X�uJ�d���ƚ��J}F듰��1a�[�֌�.�Ʈ�]�,��F��k�G`�iB����q7�Ѥފ�b�����u\�ɧ�a޹zå/���j<��Gq��s�J��r�L����K���+7��F�Ԭ��H��O�u�q�W�`�3���z0��,V�CI����lK��g7�;��Ye�Ѵe�c)�ܡ>�>%��]��&^�X�.�]v����C-�,}|�8t)��F�r�}foE����Hgw\�]t�]��+�9������.[q�<��қr��t�̮�$���ݸ%�$$��ݖQ�����;��T
�ny�S�MijF|���s�XY�^e�V\�y��=�+�����g��TrG��Ǻ��D]ҽ۪@F):�W��zX�+6���D��{=�zg� �W��y�����IO/�	�Aϗ��(������]ܣےp�Uh9�n��9E�A�x��HU�q��r���9�����Я+�GR��Z�y�k�9;�V�������K7w��^>]'c����U���U/29��U�E^G������^Z㼼KId|���v�wHO<���U�X&�"�N���y���C��*s
,�udz�'�n;�q\�=����G��<�|Z��G�;,5W'=r��W<7ݒ�#�R�㺞E�����pꆼ�𐎢W���iN���y���y�a��I:���u�s*�"/^x]�e�ʌ�]��WSPw@�$Q@��(���͗?�U��jj�;����pn��_N�*}> n֝��_hy����p%��礽@�ڞVZ�S��2�.�ñ�͚���7��g{��_��y�M+�Q�T���@ɕu����d���yִ����w��*����y5O=�j�����ށ?1ޯ�C}����P�䂤��<?tJ˽�>W��k!.|Bi!�q���=þr:�D�^���ь�����/�{�v=���D����ׄw;��u���^��T�r��J�<'�]��Q����8�bk��ޱ���Tz�Z��qC-��ه�b&�����E巌XdCZ���ȧ]욶�ѫ��覩ʨ="�"���������wclK����P~b��+���l�{�:���D���|�.�E]�Ь�9����j��z:���#�A��֬'����QXV�v�*��!�e���Ӝ±�E�[�f�_�q�>ۺ�M�h�y��� �FRj��+�;��+Y#u��P�Ð����e�k��u�m>}K��:�g!��A�>"���v��t��i�-"Ho3��P;��w�zR�l��j�2f�x�}�o�CK���RT�ݞû�p�c�%��ɖ���"�$�ب��{�S�q�vy=�8f*G{�PV۝oM�Id�w:�5y[#�L�켙��㉮��gm��WV~Z~�lX������	�M�nm��?:2,�x��k��MJ���vһaW�&�ǅ��z��V�}��4����d\H^���b���g��$J*��Ǖ0�-�X��v;a0^kOm���6�y�ޕ}y���\�G�b�ܗ؆��㡆2��fxɖ�L�\旸}�|5ne�-����܋�{�_G�z�X]P5zA��:�h�X�������
1c͇w�~����k�=���?;oôO����=:�!��荊���h��lHj�wP����w�@�E�i w7����=�{���5�~���9>w�_@���r�j����E������������#ФWFV4�Ϟk�,��;�������f�Fc�A���'�ꌏ�(r�ŋ�Of,�����t�?��:�X}�!
�+$md<>�c�{E�ٓZ86���|Vp����5��)�Y�CTt��|�at���t��T��{ޕ�}����W����vVl�a�6�\��`�r�fl���B�:����-7Ѭ2��S	��.�V꓀���3]�]ds�u�s(��Z�Fj_�J��x/C*�p�|�/X:���aK�NdV�3��2���L�f�t�5w\��s�����I���!��;g�z�}��.�kϮ�=�.�:{;շ����ö��j*!W��I;�����|���:�����yAh�S����O�5�7����[È�5���}�n(mi��;�7w"���̻���`���Up�z���4s�2]t�ӛ�}|/Ϳ#�.�~V�|s����"E�>t�X�o�"�j���4NI��z�9u�`_{1\sm��M��.RW_ܗۻaS�}����o���3v���Hn���w �;<Vd��/���O�&�G_oцS�ė]��I���-��������3�����n�ϋ�����юt�j3,�ٺX�\�63����g�Ph��/��l���H����Ob������ݞ &�NR���
�OT�dؾ[�Cu���p��ӛPf�s�˚�WwX!I��b�˥Lýw�c�)gN��M��[��-���/���Sۥe�K'�#0v_*^F�Cũ�v-a�\ ǕJ�����j�+0j�أ5����k�q~������"+��VJ*�L�6�׽P{lm�OZYX{�}}m�����z�`�\� ��Bjs����N��7~�Rp܃��s�|��QS���/>e����Go׃�c7�bU��oL!��Z5؋���Z�w�͢��\+o�^���X!R���|V{t'�ڹ&᫼��al�����v�#�V���[|�t_xg��<�U��C���58��a͡���/Qָ��7q	�䅄�b{�q����IK3'�T�s�զOP��I����қ����@�l�qj�J�g�˳+�v�gW����p�w8�[ޣ/���}��[�g�{|u��8��n�ʽ�W&�}�:���n��l;,�O��ͷ�>=90C�ydV��lT�p6��{[����u��G0�M�T�q���m�����^y+�^~�l+�W��TU���v&��K��zD�;�j�}�$.|�O���ͫR�[[4VP�]�m���]�������)W��ÃՃ�s�1蝥�Xb�땺�0"7�e*&\v�1o �1ݙ]f[|�����j�����a���J oUܫ8��v"���o���(��dE{��k;_\sM�6C���|s�I�95YT�p�{�{{${t��? ���";Q���#v[u�u=�D]����7�CJ���c�����~��X~hh��u���;��I�@�Gq�zc�#�Ԛ�oꉹ<1��˰~�Qa�����K�H�U���ы͜㓻��u���O�ݍ���B��D����
�W_�|%9��t��i�-XA��j���]x�C��!&�缯����y�o^n,�&~�5]�/z�l<�C��?u���X��?&��3�H�[�����4�f"��ћ�?���{�Fc�q�~�(�)�*}xG�ߏ*�s�'��B���GR��Ψѕ�a��7����#�]�f���#�x.((B+�T��5<ùD^p�O�K�����ܾ�}ׯ]����\�y���Kq�Z���.�4L�ޗK%+ʄ,ĩ�ܧ�ZiY�=Z�%e'�Jz4J���نX�b;E��<57E�&L�����6��]!���9�E�T���*b��&������C���U>�P�b��&}�.��;����k�u{���N�WMx�t��4����<�;Av=Fz��~aU �+���_��}q�NQ��N{=�xw�.���(Q�5�<�|�E��
��f����@�F����\���CZ�ZR	e���/�cNs
�-��3���<?CQ�w5y���u	RH��/�C���c�6kk�sHI�<�jz/���̭�x�i0���?qv��1<hM�m���<�e+m�J^î��(h׻Lז.��O����PV�lE4���
�}�nU�5ՉZ8��h����$n�v@��.N�&ٍ�^.s�*�3潖w���r4CY>����j0�f�����G�r����t��C���������s�v|�E�am+�k�cn�H�x�V>�~�%��w+��4�������V���j�K�W��r��O�M�ow^ٚN��ߍ�E�v�Y.8T@��w�}EB%�����=0�Yp���R]*.�0n�N�Gf�zs��.��v�#J�6s�Y[��S]֔Ƨqb�ºԓG[e�꾢�ŕ�1��Rګ���M�qb�����˗л�MwJ��p��uTmG���1��������]��֊*��sv���\�^���tY�;gTSbzGH~�~��E��FjBj��oڋ!R|z󑮡�`�0'ցٛ㙄�����2C��`��b;}�}�o�?e*�2�����3�r���ګ���6��~y�!�ڣ���!�78�z��F�ch��{�F�mrϻ�R�V>]\/�rIB�k�T6�Ӏh�����`�d�V������}D/D����^���Bo�!i��у���˙��s�D���aI��het���6���1��:O�m�m�F&�X�k��4ok��Y��cB�:vju���f8���e�ξ'�O��joV������{��UG�ƪ�
��w��b�v�%谸�5r�TK+,��u�Xj�B��z�^�{=ïz�#�J��J�߂��fj�K�:C�O+�u���{�Y����,'�o�G�V�#`�!=n5�\�����e:\�L0u���1"ֈ�`�p��}���|:Z�L�Z���\c��Q��R3��M�|��;9
����Z*ʜÀ�s��,v6�TyHn����Ppv��kF�򴮽���9����xy��6Ciڤ��/�e���O*9�aS������'<�~�+�!�M����x����5����r�́�9U��l����a6����C��l��hv[e��^��=�
F�Td{GS���)����V��0/��ϧ��}������EX�)%�t^.:��L�}W�=�\����]1u�g��sq�~��Z�h��uW�1��w:�5�S�k��2z�'X���*:~��\����{צ7ޗkWm��:�ç�y�.�n�.#��%_} �^Rfh��+�_��#���>��rfy�^m=zWV��W�ȯ�WN���{�1�]W��WyhBED��_Mnx�������	��*�>1 �=�~ۑ>���Tdx��v�U8/Fi�v�Z��ջ�lw$+�����#O�����j��?�L�#���}����J�}r�9x�1��Z��ku'�%V(����,�wk>��}�����iE:�}O�y�Z�H)����rrr�4�D�Φs���]:�U�������%�t�b�Mq�O���Vo�Mf�����gB�y}�OMo�xrLb�.�g�t�y�ځ҄��}�;�<��x�W��M�wu��y��L�4=Q ���6�J��+j}�8�� 㜣���kԻ(�y7��j��]����,ʿ�q,ٍ��/z�l:Y'Ow�yN��7;=�\ڲ��
�,?���Ot����Jn�r|34�Z��BƤ�DRb���/���������M�{ ዚ�!*��8Vx�����1�tа���cn)�ڎ��ݖ��ٷ�;@�ˌ����p��'����.Vz>���������+���.���Ε=a��?j�c|y�������T�#���������z��~���}w���H>��j��{�����^�2���u�*�H'�40��5�lie�{���+�x����X�f����ް��@�ޏ�Y�"��"�ǒV�A|��6.��N*Ֆ�7����Ԇ��Bg�gEW~��l�԰���_`�4C
z�����˅Z�(X������y<��yx�k� �q��������^,���+�%ڝ��1���[̵3yD㙥����q��a�o�X�Z���f�>���Sl�{���~�v#���F��]�����j}�]3��w�x�s���S��kX+��=�^�~f��s�p���˿�XgiFa��e�G��|:%��>�{a��Q��m��#�g;�]~����ɷ8�X둼���U�"$za��D��޽l�}��i)]��W%85���M�a���8Pc���PC��ШJN&����&�w|V�-�Z^�q�~��P�G��'�sQ�.Ǩ�Qcn����������|����MI:���#��Ǜb�0��g��ō�r��Lv����n�����F�FH����x-y���sI�!�콝�F�G�R�-��
��1���,�X#�$O<����`N?X�0��ʌ�|&�Ћ��8�Jwچ_��h�j�����g"Bp��U��{�� %~1/5Hw�vf�%�����Wd��u@�C�n���ݔ�1�K�,A�E�a�Шk�7ќ�B�Y��>��mH�,�tK�z\Դ��pq�@�Yx#&p�O$�&�g��v� "0v7ʣ�W���a�H�tPALP�o��tô�:��f���:�k\�,�M�����zdBƸS�Z�;��+����]���� t����7�ܽ"۹s�Aj���4�����dp|/[���!�`K��h�[�2�0�
�Y�^��\/Q;�(\����ؙ��BK�1j�&g}z�ɺe�;7�j�<+��92��*�"��X��Y�5�J��He`�k�P���▘�"�7�3bF��+jo:���u�P̧�ҷ�+P���r)\ݠ\j{L��*�p%�-I�d�#�݁�ɛ��:�ؕ�

CQ��ie�+a�b�d�����6rɉf��Qho��l�u����Org��@i�W��|���z��G����=���ǊD��R���}���	j�n�E" ٸ3Gb�9t3H�j�I�|�p��:ȵ�DAԹ��˽��{�߼���2\�Ŏz�}I+����Ԫlq5�x���ZkqB�3���ft:so��J,n̩s+�3���W(�#�W�sA\��qw��e���\
s���aOq����:0_y{"��B��^Z�cH�ܪe�v�D��j7*�ak��q�v�hQ3Na9�AD�j{t/��(����vh���Gnu�k�ٺ�j�v��"OwV(�n�N�����i�s���B���M���t�6e��
��דrw��K����u���du�2�f�t�sQ�TK��2�d[�I�`�ۙ��V6k`�BS6&qٙ��7�^��J��e5�q6� 7��	�(h.��u�-��vnqP��e1�j��J�9��]rΤ�n���틎�K�7�B���ͽ��v��k�+�V/�:Q,	�n��NCɳZ�]��SΚԔ+1)OTܣ�Ӄ�-c�_^`�.���G���o�6NY՜��)��Ġ2& /:X�|ݛe:GG7�Jܥš�
\�:fN�����-΄dĞ$��G�Q�{�H�5,�Fq��N�X6��;�����[Щ	ocC9�]Y#6��:�O��WD�,"؎��_`�؝�K70�`�*��Q3&k�飕���g/����)b��z���a��9�o��v�r�X�Z�i���>˖���z� tr=�=�Ї�c�*fSGf�4c�@�׎��;��e�v_e� 곖�].������""�u��v���J���(�!�n�M�Ҳ�\Qm��J�wu����s����ӭ��3xT���cJj�&�.�F�Ԙ�p}2��d,q�nѽ�/0M���F��L=��*�R:�����Ѣ�B#|����n\�L�JXI�O!��;ph�%��-*V��e򋯣v>�F! ��!Uت��B��Jg;����(*����"-).�)v�'V;�<?� _"�j���ڻ�B� �K��V`t�5���s�)�/:���۷t�����{=��g�}�S^=ÔU�'�����-sqh���VEoK�E��h�	{���E�^����'#us\��1����C�;�H� �a�x��H9EV���3wv9�9Ⱦ>+�=�t��'�Ҩ9�-ݎ�99��$V����x�hO<��Z|�\�Ing�T�d��y�t�LҼJr.�ҹ|�k��sΨ��Bm�<M�\���\�V�x�(Ed^��>yGwǏw$*r͹��=JL���2sg4rt���㧕k��⩳tw��5�]*(�Q���Ȥ>w��&t�מ^x�ܪ��y{���TT��WOS�\u��ⴜu����wuE�:�|y�l#T�3��U�$��t\r�R;�5+>]�1w.�)��9���dtty���;�.Ov������֥B���V�~||��������J��=V�VK.:4����3�ɉmK��39�[`�q�Ɯɖ���;��#'��Is���\X�.o~���m�tf�sGRG�~M�|n^���BbY���`���X��񞉬G�|�8b܇�T���G>G���\���b7g����nj�ǵ��3�Xo�!m����]����۟wy믭�Ob��i)��Y"h�U-�E��t83��re�jw�m��Ńi�>�קdc�x�R���zU��bL��^(������+;��������op�j��<�4�Ҽu�����@�����	���{Qu�і	�3A����[?/�{�I�����Ӗ#��|��{Z�@�3ر��$��=ޱx�����.!L�۶��	Ұ�_X�_Ppl;�RaĊ��6�hG}�~�z�����V��c�r�Jk�
��Eړ.Mp�Ej��޿fm\r-��n���}Y�w\��	�/��,�Y�$�PÕ��TG�;(Q�Qd���,ai<y�x�E����+˯'�v�=��84��(����S���)E��Go�����+�� {��������$�cp�n@�q�Cq��UP���UN�q���YN���u���Yn��1��,/�� &H11dgF�;�4k��p3U��sA�]f5������͐�&mGY��ш�&:��7c��z�V:.v`�C�!�����O� W���f�X]�ksW]{�j	c��^��q3R��a��K&tD8��ي��~�5[�&���q�:�k��E_2B�ޫ�f]�< [ �(��3�����yz,Z]��!Cؽq��
[o�T�?N����]B�=�:߶�N���v7�(M��>���Wb"���������v�@��~ϻ�n�Y��k3cԣ�2��`�%>��C��?-s�"����O����p(zc��y���9z������x>���n_����\�~81���I�ß��Tߧ����eš��y�Y<��.�!�TD�l�gV�,���\�>�D3�X3�̄7^�F�+�?H�֫��5D� Vk3��Tp]0�MՇCE���kk�SҴ��ߖᆧ���s|;���Ӕy�9ʹ�[���Y��(�m�X*wu1m�P��iv��㕘�ۙ�������v�HV}�y#��umԉv�˵NA֮�E��\�z�[�!��n����Uif�lsGt�	�o��Ol.��K��e�`�F}d�����Q���^�Hpǅ4�@�m]v�ֹ��O˫l{���VfyNd��W��d��^b�D�h� h��m��yO��V�AdaF�f@�E�=�>��0Ҵ�<��?xb�4� m浃�j��8�4_R�ӄ̯l֭y~V8z�	������d��[�H1\�P���Y�kåX3�I��9�v��,]g�f�(�n�e�}�,g���f�Q?;�l�i��]�}����j���a��+YFƤ߳S�z���Y��.�AI���:}���+�
��.�=�؜��a�Ͳ1�d;Yk�=�(ш��QFll���oi�Kȟ�vR�Z%���P�����a��h���w�^��r8���lB������ʟA� ����E7c��r߻��Xk�}�7w��vv��@���ڷ���]���Eao��g
�}�T�_���f���ӳ2��`X�� Ԣr�����w(r󝼝u�>�=���S���U���ƭ����-�nN���MFM�:g�2�R�7]��3.�ٴ%$����^-�4.W&9��'k���g�_ц]�>4%������a�-1E�֧�м�U�Z��W�*��^r-<��c�_�Ǯ{��#�ۺ�Q��
����pϴ���k�������⟻z�:o�F>�|��ϩ}���ȶڲ|tw��+�у�*�":���	5Vj��/z�Ǽ�	罎C7)e(����o|a�ؠcDf93��2�uv#�s|SH�d(�fȟ�N�el��ՙ�h�����ǘ@���� �|r2�/K2��5y��>��Ȉ4<��w������6Dfl`�a�\��w#/�'1���ʓW�g4�}���وF;d|�[r��^X�DMLK��i�����4}��:��$�>�w�߇����M���у�~�=cj'�&��E��渭�U�Ӿ�����X�x�^���rD'�_5t�Mʛ�J�鳾�d��ʢ�I��w�Ѳ}H�n����(l\�����Rj�#�ӡ��BoB����u�UK٠��p��m�$�H���w}O�$ջ�Yd>��37����ም[�]&j���6y��o��92�7S�ͿeҞ�m�v��r��df)�D���}�s)��w������>m�y�c��$&�(y��C��I��M{���66�vuNV�����o�Z��u�}�11���y\͏�����Ә}��ͱ�e�">a� ��lK�?�s���@��Ε��7�;1$}|-��~g�շJ���f^�������i�]�UW<�y��򺮴�t��p��9$~���v���1ןvv<�PC�C�t"�[�h�y��vM��5�-c�T�So�ϐ�-�ψ	b�ݑw."���y؞���S��z�l�����W�)�>����2�Ŭ���������g��팞tˇP7�q����h���;]�ݏ�c���A�M3�[.��["f
Y�h�K��fQHh����W���򥅧%�t�vo��YIo���ޤ-:F���o���{�Bj��L�"Ou����=��9��\D|�}�mbr������0�eqcb�3��Nk%����u�OlM���oy�'9��c�),�]g������M�>UT,!,b<�}:wK��j�;�V���m�h*�,�J:�v�P�����S�����<�fۉ�*P�IN���t�_����̹��]���.4�ڹ>.�X���Q�o��~��Ta\�scy��޷���ָ�>����}iҰ�]��`F�b*=հ����y�"a|,z@��YMrC�r�K�Çp�c��������F���ל��ΌB�%HH�\�\�b�>����/�����4�D̐�UTS�9�1R��n�ܨ��A�0U�ư]�'ڷ[a_�WFk�����-9�����p�w��̾�����I���T��k�5�q�oݜ�Y�!����$�v�ɯE�ƍ\�����������Kٗ���f���}},<)5e+G�|�]��rlǲ�C�4)#\Y�s���+��W������Əe��O�~
[�ӿ�$cm�#��,��=�^��V{�In��Hg��v�;�-/�yn~w��ͯЋ��݇v��nC�Vm�����~%y�4m�'�IH�З�{��ݲ+[)!g�P���dμZC�,=�� ��qR�^G\.�	Mv�b8�]b-xr)!��	-�z�!6./-����-g��`[U;yϗ$-�����J��s�w@Mnc�'r��ۙ�L��Y���<�rxl�ޗ�PږĹ���N��U���Lefz�}�&앲��Q������	�p}�����lG��H���8e"�;���Ϙ��U�[���ix�F\_�"�Ǜ���NMt���}ճ���;-�'�ܹ�}΋>wF����n�wC��z{_e2��O��5)��`� _zտ2;Ȳ=]�K������#
�ߠ�*�ռL�T����c��~Rxo�NC����͢�ꃗ�c��d-��\oս~�~ɭ��h}�0C��,x4��W�H�X������5ҡ!ub��C�|��7��_v���%t�aH���϶�Z���=�{ƫܠ��{�l��y̏_Y���M���B�Xd�[�K��r���4Y�KUL�	˂<Jĺ������؟���;u�d��W���w�YqgLz߄�1����-,XF�Z8�G��+Z���8�6�O��R�E�k�ڞ��ЯH�&#Ԣ�|!<�4k>�����Դ����HP�K�J�q�6�[�x]�N嵷��6C��W�K<�P��ڕ�=
gP޻��d��Ǫm�%+l��S�������qJ�׎yo���}�W'��L;��"�iv2̫Bz��2O��N��;�B��O�e;`����mP�0󹶱�n�:���3�I�b�G���,�g�;;i��vj;__��;]Mg���� �}Å�u!�/^ZD���0��M{r��-��+��y����_�x��z��ڦ��X��g�$��x���.�4%�����;�n���|�3*��ˍG�fMwZO-<�G[�}����� ��P�z�ߚ��!�Yg6�G�����:�@u<S���@7ݍG5R�z==�"N@��#��v�t��Ç`��}y��[~&��j��/zGS���oJ�%x?Y��/o}Z+`pb�O�7P�~��ߟU=�uv#���5�����8�/xf��u�g^}�P�Og�v�jo��憎���M����{b�/��R�K������TU��Q�F�t��S�:�fS��Ur�6+����Yl�:��فmw>��s|(2S�Zҽ�6%w�.�S�l���Մ��55L�2� ��(9��>Qnf� ��Ն^tw�s ��|#v䅽��q �.�`���_H��z��T�w;<����p|�+���al���=Kȝ�VUj�ݚ���fj�����*������D~�44��r�M1j>{�1k5�fΛ޹������6��6�=�>�r1x�QdyO�y=�;��fߙ�vк}��}k���&ǽ��1c�x���NԥEOV�	©�M폆���-��1.Q��%�v��clI��[���]<'&&�=Oz8VV�<v��}�W�[�`�٭�w0���٩�'di���tgwn��+�wk+�o,ʰC��L[B�<�1U:�(�l����y�ޤ#0k�M�j�v�׎_�K9��W:�绝��Jg��wg�׾�
z�y���I'o�m��cr�9�I���`�{+]5�"���硼�(w[o>�|�z����%���&;����`��k�׌�q��z��B�;*+ρn�B�ý��R�u�6�f2��W�d�^E.�9��nrI8���zVY��ɜx嬎�}5��&�{���o �o_G��C���JG�����{�V�`�5�j�uC&�7�>N���n�t����'�������Z;��6�_<s�9��t���{9T��r[�n:��}�B�#&^����m���!m��7�A9rb=�t����i�%޽{f�Q^^(�_+��#�cz�(3�b�ݯU��kOw�w����i�������І���T��Np�1���b������m�%�|U'��>~?�����o|8��������gsi���13~�;K�G��\~w�;Ǽ�ǵ�!O��l>��[�v>�!�*�^�:���Us7Ion�.'���
����to]u���t��(�X�3�to�<So^�^#=�ފ������j������Wu���p�"�L�x�H�,������3��^*^}?>�h���C���Uu��]�'ڵ���z��=�`�JS�زP}��GoO��龣������׮������7��W�}c�(���`�k�C6����?��������[�(w����6 A�`M�	� A �"� ��p���;`� l z�f� �� DD��"�8 Acmc "�� �� A  A  A6�o+�8�l�  �m��;m�A6�d��G�F�l�� A��dm���;�Ѷ� �m�6� �m� �m�@ Lm�	�� � u��m�6� �m��� ���m�M���m�M���m�����  �m��8�l�m��;m�A6�dm�A�0 ����m�L� ���2x���� Glm��~�������������q��������1��������뾏�?G��o���|�����%���6����G��ݿ���F�6���=��o�?���cz?��?���y��m�lm���_Ӿ����z�M�����������8�������6��ll`�#�`�`;l ���m�A��g��gm�M��1��l�d�m����0� &M���m�6�dM��q��8�l�m�\cm���m�m���`���d`��������60m��aLc?��f�����|�?��`�o�?�i����o��������=m����?����'��<?[��m���{�6������y���0clm��m���7���|z>�m�lm�m���7l�o�&���([��c��f�'o�;�����c�w��o����~���?�����m�lm�����o���|���~���������7�!����am�m���������`�o�7�{�ݔ?����7���������_X<�7����r?��m�lm���>w��n7�[����ޏ�~���߸���A�ދv�o~��6�����~~�[�գ~��(+$�k63�I�l[0
 ��d��H�Ϟ     �� 
  h �      @    �     �S@;f�b%d+D�$5[B��,��R��6��Ե��m���T�� El�k1[a,��nM6Lֈ��Hƶ�[VPKY��Kme�V�k�E:R�MY�&ʋ0�֭m��֔եM
��fk[Emh���kcm6�i�d��֭�%eZ(�Z��*�fjm6�f�4���mmflm}۶�Km�mVS�  Ǭ-�F�k�����cG���һm�4���=zn�5m�zo5Z��n��.���
u��^����{�](�
��U�n�N���h,շ]۶�Qb�m`�F���f46��|  �Ǒ}�aF�P�B����xt}
44+�$��ռ>�
(}
cB��4��(P�B�>���uO��-�'���V��S��e=z]���{�kӝi)F��{�ݬzj����p7��`n����R3�����l̕�   �}�ѭ5�>�7���u����:ճ�Mle��݊q�c��[oCN��ڸk�:6�k��c�*�j��"�d:]X�ۼ��Z�Mzks��r;aAR���mm��V����d�3i�m�/�  s��h����u�Pk^��{�ojuɋں9^�㣻-��s��MNJ�¥�cOw6{�[ڶ�[��ה4���Uh�m�v�a֍iW.��j����iZk&Q3�  �ꢔeۈ�:[�:�E.�u (��^�����Ҋ���	*��W�	
�MU˸P��gZ�f�)l�5����`�|  � 6T�*�=3�M�e�F��w��UUT�uPJ�wgn�֨3�
*��d]��*��uw3mh��6��ʶ�f�C+IcQk|   }��R�Z����ۙ�]���nwu�	��U
+��4��Cgv�KQBu���@{����޼Z[jPَ��l5��Vo�  s�B��w�P ���� w�� �nˀ �� = � �hY@ ݳ���� @ڧ,���j����&խ�+-��  �| � ;��  ���`PN��U�@� �, h��
 {z�x ��w  �{�x:�GU,@ ;q���a�ͭ��B�5_   ��� ��� ��g  ��  n= n΃q0
 �ۆ�� ��@4��p��׶� �O��*��h�B)�)IR�h0�O`���S��F����*��� O
UF�(  e*
�� j~�~����Ʉ�~\��M���B2hl�-�i:YRꗢU��ye
�<<=�<=�VG�����6��m�m����6���6m���1�M��6=����������ӿ�HG0�ݦ�ׇMz>v��!�J���{l��E��+�@7�9{p����CuB��R{���(Y�ݫ� �Y��۳�EB�Q��ue6�Ӂt�\Bhж�([;��q�ĥ��SZ�E���n����Rvt]x�7U�{y9�M�{X���i���y�1�f��t�JF��
������s���'3�����v݊f�M�Wp5�/l��{u�Q�j@�[][�c׳xૂm�7Q�O`"�ʭ90��[�4�>���ǽ�gXV�{D'&���?nlj]̷]43Y=WC�VE�n�n����ˇ���:v!U�$�qm稸�1Cn�ӥ'�m�ˊ����	Hu���^�`nct��,�a��u��'f�-7�����i���8;���NQ��|�0�K_n��z�]X՛�ݻ�dVo7��K���xJp�ٮp/�s�,ݰa���d_sЏh����޵�^�T�֫��8&=�=����i�*����qe��E�V�	�$�J롤F�.��)�����r꽪�7;zVն�-\0c8Ej)���v,CdH���&K8�.��oZSb�7důH��GF�x2s���Z0�0,ޘs�M)�n�.�ݓ�|v`˫3Yx�RL$��AS�{�O�����u�|��uYF�Y~z��7�,v*%FM�exJ�)�^�Q�M��QC�/Z�reB��m�"i!�iη)ɇ���\F�2��3qk�f�ꨟ@�n����S1��ZjL0t�{�^�5���K:�v=�0� ��;F�
:��Pݹ��V��&��D�%t�3G��$(��W��YŽRX��B�g	a��wW�iSb���׀���{:�Mͺ�ֶ0c��i��7��5iwG6{��݌����С���$0:�ҫ[� �B�o�IDIvtl`��A,�!o	�@�����m�w	i��fƵێ�c:Wu�,���u�-o��p��q�W�d �����wcG;�a�w9:�^�aV��'91����9�H���� $����b�����vt5g�.kD�8&�6c� �-��� �v#�N�"�g7�ݳ[���w��6p��k5��8i�܏tN��k�%닰>�]#��E�b҆�7�=�>쪶0W�5� �K����VSN�z)�a�k�܃�` 5�n��}n	�b�&�jr�ՉX�@�.g;�ٻu��v�&k�6
d��P���!�;8r�*�,�s�C��$�qQubD�l	
+��
y��W7t��hj�f��d*	X���,{{8��^���ç�9��c9�{��2-c(���%j�$������L�ȇ!��sʎ�a�}�r���9d���Z�N�pHM6v[��C����	��ҋ�NA�:��D38�lK�����n���F��>ÚZ��7��8�vج�4���X;r����7����jY�M|�Yd}�N�N&��f�
}�>\z���fSz�rG��{�f�9Bg�.rۋ򘦈���>�:B�(���郆�uC�����z�Pj�.�X5>}L�0��������.�
�(V�i6��;�ɺ�E��|SQ�Q��V�{ͥ1Ż�
���H@�����& �cT�&�鳦�L1�ea!�o��w$�8�okwJO[NF�T![�"yN��p*������&��q1�D�Oc�~�:s�ǯ�4-���np z�\�I����/���%�����d��f�j��!����F�M}����E����S���y�*�������N%�B�5	O�g�7�3c�M������]��$�Bq<�Bs/r���zj�oh+wZ	�3�nvk�^�����p��,����G[��u��C�֮���d�X���ىNۦ�o+
��gg709�H�����,_ITZyZ�$�w:S�t׼w^�;��7�M���+�{�e�WӺ�R�u���-k���T��h�&���p;(9�jG�)È�X�I�ȳ��7��U� ��*$-�W86w#Ý;��UoN�A ����+zT0�ګD]Grj��R�1��EcWW�u�m��&���îhY�_!7�pgv�t�������X�1v�L4�"AC{MRr��P61��V{;�$��aK+�\�����<>�\8U�v��Ч��A2�n�7s��A�u)�a�� ��{�����ݓԴ�+xLG 0�iʸ��vc#���˻�6沇z;/6Щ�Ǝwmw�ݖ;�]��q�aZw7mZ3qذ%�7�z�cE�ʥ����L�n�+��M�TM1�l*�^4��B ���V�z����t}{��Ǯ�5�$���&tH���U�o�-�ӭJxu�ݪ}r�``Hb����|u�Q���c��($�=�[�3g�_
�h���s�=�>�~Y�h�V�$���*Q�#���	K����-�������	���4����%��P�I�^�s�s9��a직[�����7��+��`�>�쒨�Sf��ȳ��O�j�e�ĕgm畭���SA���pN�{by��g^[{�;!/��q��uS��6lz�:���+�N���[vBRе3�K�3�*�ͬj=�T�m��d�s��a��r�5�.U��M�Z)��d�Ŝ��pѽI˩N���03��o=���o�����źd�ET��f�!�6�>h�pF�k`���8��/Nn�ɍ-��9Û���}̫kǏw;�5�3�|
�����Ԁ'�����ʱ�/��}j��[Aդ˷�V�8�e�gI��|�;FN�R�L��zAZ8V�X�d���4�F�CC��-d.wvI��I1�-�ť��%�vh�pQh={�ݼ��:.�CsN�p��݅��+��#�.��'r� ����\��磉l{{t��Įb��J�����yswy�Ρ�6�Y��隫	�0�s]�<���Hq����S���9���i�=�]��`Dh���jA�l�1'�@�t�F�l�k�Ӵ�9-U��صlm4�� �˷V�r�Y� �\*�i�Cϵ���� n^W�˹^��Ʒ�p�W�5�����7Wm\�Xh[d��ݝ;�-{�Ѥ�l�ݚR�H�ƨ�׻�8�<���f�jF}���/[z�[Iq�r�Д�t향�GJU����Տ8���ƝӿQ��_vn9Kl�: �J��74�Mü��A�&��T� ]�rպ�����r� 9%��C��� ��ׯ��u�T��=���p���p���S��oHv�֗��N�7ZL��r������v,�3��T�v�_�
����f$RܴG��2$��"΀��X2��a����UI�8�����;GD��i.�K����O^܎�(��Nlq*6To	Y����Y���5�<]����-�!疜öp�s8_�.O�@��ś�Q�����6�'��#u���{���g��c3!/�mÂ���і�r�2uw�Ժ�¹�_a㝰5P���8�v=��T�^�T���}����i7ݺv��+���ۉ�a��	�L;ܫ)n����ֽ�Y�]/�vG,D��S6]��u|�]�}�N�[ywǸ~��wK<������Z6�n�kyB�s��>���j�� 򵳷�X�����Yoxۛ(S:�]�û{�(�)�Y�y�q`��,�[�;n�)ЏqoC�*�6izH�gL��9�%Kcr�bz9ح'�iZ_Ng���"����ץ;:9A���^��.Xw�������6>�zD���|V:�ۂذ�w^�h��o �EXj���|�����*ᩬ��u������^m�3�Lp׏4#�n���l(�n��i��G.븆�-ҜxRa��o���;�Yp��\zG��y���L8�R�Ӌ �kֹ�Ӳ�����NuL����@�f��E�yc^�V�Q3Y4a�X��; ά�;D����L�����;۴�8�mdd��&s�W�.�	y�C�:S�uI{�q���n�j��:�<lsv�;K�/c����R�}�cW5��-Y�Q�uط�.��v��So5�U�q�f�3�m�/i��k"oovނ�y'<� ��5�ΫZ�ค�����xI>Ri�\ȷ��7GYTԷ{upR>��9�߷`��O�Н|X��M����l�dql��2m�lU���k�9Q��-��nd4w���{�f]L,Sn���Ik���ٱ\4��rѠ(#�$��D���(y8��_
^3�2s�2�FL�n�f�bɜT�:�T�������w�f8�!��,��(f��#������v�����	tXr��(�W�VB��}���%�܈��W�oc�&��]�5�`�.�NQ��gR�k�{�%���P>��j�e���v)��"�92�8edx�����8w$��Pzgr��.[��n�f�n�!��
{�6��p�-R��\zg*
�X1<��F�wF����:y�ҋx�˚����z3p�T;�N����4��M�u.�l���mra�n�H,��u��^���|��(
j���P<�H1��v���2Dӫ�o{j�n��[0 �@3��:&6��7Ӵ��3ݠ�pB�y
�9��1�ֻ7;t���Ǽ*��4c�Y�p���y�MCq��MyR� {��n��e���T���b�j(�$��k�UV� �P��rZ����{�4;�a���V��$�wb�����NhYϕ:�>���>�/<q���)�K�sK"��{A�����	��}��R��]M�<���EZM���)2�6S^6q?o��ݢg��!;���%I�*u��I��br��^2�+k��Hn��z��A��ι�JB�\XOvB�ޛ9�]vӏI�\k��k^�Å��3X���۹;����P3�[�sLԹ��,�:�nR�N�/q�Ό�� l��-�� v�wo7 {GM]yi�Y�6�ձv|y�����7p/���b�u���K�h����'������R͓��hŏ{���p��v��t�j�^y�w�����1s@o-���s��]]��ͻ"8�7*i]��μ�Pf=n�}Ǚ&
�P�?��aܘ0L�j��H�f-cn�{w�N��'�[N�t7�[�x=�4,Z`�
��f��y[�����S;�<��4q���k��QQ!�B���Lc|���!��)m�uӐ=#������AT�ǒE��� Y4���.ی��;v,໧vw���*2�h�';�N�\$�)���A�VJOR�!�K��\�.zn�׻�Q��V��uX�U�����������8t��wS�w;m�H���U~[�0�@����;���几ɛ�����{�Gz��P#A{�7;Y�%�s�v��/�PNe����W�1ae����")� �w��ɛ�{;FG�%���P��ބ��
��dw�w�ɻ�q=���od�μp35�fN9�ܹ�7I�FQ�UӠ�
m�����C�5�Opi�g��\�tW��T���׎s��;����k�)��󏺰1�3�ݲ�AJ%�i\�������לz	��q;1���@��`'��m�-�;��W8�bn��Zpe
Lq��ÄWm�������Q��HK�D�O��C6��>��8�3���N����Z!��WVi�gX�!������N=Ci���7�2�g"�MW��WD�X�X��䚬���Z�P�Jtgn��7W��s�"��2'�N���S�@��j9l���;�gV<�0}W;���F�L��5Xܼ��WGk�<�:�|�E&y7wN5���{UQ9���;q�0�("��5^��|ܧ^90i#��3 >A\)\'(BZ6C��au-�@�a��%�����V�x�Suu�7n�zFve}l�f^�
�l�����n�kP��[^��nV���2���ۄv����q���ܵ=Ᏸ�o�h� uF	7��ν��fl�8Q܈Ϋ^ᏻ��6���J:��gv]5�c��̻';��\�5�Mn�r��e��L�m��1�<NamkA4ѧC���ytj	i<Q���ŋY٥B��G[ON�4� 4�l��{/�5��@I���5�����L�Y�5l������+7y���.���y^����osp'#=���Ad�oYJΛ$��Y��Z_=�.�EZ�~�݃��-�V�m�'�Ff�;��#;��-g���1��E|D�Ġ��n���'r�Z���,�V�%CqYFH�BJ��'P�7v��s�w~��4eJ@��k�uPʇ��^�m=���ndj+ؔ᡼����3�ߍ?,a��US6��cP1�W�hGP}g�Л�#s��M�V滺�<F��9:Yr�V�4�w5h罰v��T�3�a^PH�6�rJ)/;XN
��Kt�	9���T:�Y��8Üxn	���'+�&�eV�����Y����޼^T2	��^p��z�]+Q�8��!���\u��P_gU�&�lC���ck|r		ݚ{vu�GT�w��[E�p�3����`���2^�U���^ޚpՌ���#By��5%�3]y't��k@}ڇon9�FM-y�mݏB`ydow���K�oD�i�r-'	��J� 0C��`&�����r�2��IAά��o����!���k��:��Ɨ�mH�};H�r�Ś�W�֟�sH����cֲ��Fy����(�[�7ß�c�+�����2�o\q�n	��ؾz��ѳm�ɍd��V_P����mɷ� v�
�-�E�K����`���Zj���u��ԱWÕ�&g(�"��ͼ�ycHU%������H�o���d#Rj{�7���p�u����P�7���p�ċiq�Y�s�M;J��tv��P��;k(Z\��Ô�����k��Z:jr��sf���-�,Ǐ�r��::�7����k��Xj�r��w����Yԅ^���q(�������a1���;���b��"ʾ��=p�u4���r�<4�o�8f+���سT].�������&�际˧�őʕ����7wv��G7Ւq��c��Mœ��é���<ݛ��{���W�z�qY���B�qǋ'�F\'8�N�m�v��)�.�m�mamv�(����C0.u���wd	,s�� K�ڞﷱ�)E�Ug���[˪�W����p:j�@�ap�Y������B�I����]XQV֌��5D^��6ˡ�f�{�����b|1����r�����b��2��J��J�C�M��q.���f�S����om�NVl�����-2X�� :��LfA��\����j���7�h����]˥@�Y�1}�,�N�OY1ok:��7E����#��O���Ǯ\R���nOy�LM���s'N�ʴI�z�jG 5�4�R��7��M$�ԅ�A��enRk0J�`�vZF�Νɍi�����~�΅�
�������D-"^aNT���s���C�f���*h{ճ2��ڋ��d��`ѻ�/b�, Z74�&X�v��f@���
�Rp�Y>ƺ���)����u1����z�⼶f��>7/x��}�Ū�����P����f	����(���p[�e>5X��C�ޣ�W)�Ή����rR���]k�Cy�t��4l�ő��oI�1ٻ壡�����ϼ��BB�6���#��ݠH��j6<�����g����Ǌ�u^I���<��hÎ�mڵ�͘�%�]��u�eo�����]w�= ����ܔp��{���<f�k��_����V�����j�F�2FA���:O!���)�a����}���$�#̾M�ג����拺�.�d��W-t7|���i�<�%�3spW�2��Lԓ�!�0b��n$����1M�8�6�to��Vܫ�P ̺<���Y���,�-ɼ���zӾ��덜�B�d���	�V�-�ਫz�lc+%�d^��a��`x����3��`���
�>�n�B���I��R��]"��i�|)r�;��1�i��3���a�S��$~}8e|G=]HG���H,>&���y`������V@��b�D��m�/,۝���l�uiG�;6����:�;�e�v D�{�����6�f.� 8�a��f8��L��͉��ӗh6��Ǖn���t' .� \�@]Ûth�{p��Ɓ�4g�n#�}�n%�W�7i[�c�B�w�/%՛߷�!r�>}��ݗW+5�;��w�����]�r]�a��n�7F�o�<i�g�\��I%I��$e"�pǂub�C�=�TF3z�xsA��ISwx�7l��y�7σ}�wO@K_���M���}�r�D�X�J���Ġ�	�����#Dn��٤J�i�/��Z}�W��ɼ`)���=AR��Hd�|F��stK�aX��(�{�H�t(zP������ϐt�\��ؾ���3rȾ�;P~�"G"}��=�7 �k]-�]�~
W���BafPGֽS6��:F����{����\�ՋX����Ѭ��{�v��z��}v8ˣ�/�.�y���7\#n��o6X�X���|�k�zu)�ggF���Ϩ��޽%�P�P9�\��D�|�S���N�uhٹ\�ϋQof��:�`�x����q�l���G�F;�,!���̹��!��S!Vv�B�kU���/U��k���H���&bΤ4��Ƚ�c�ӵ��hz�P���"�R.��z�J݋6*j�F��L
�~���Əs7�y��������BwhO\��'�#��IPo>�ԝi�?;7�����ȣ{�+waKz�m4S32cTqv9)mqG�	NP_(p�?z/�_��~P�e=w�E�u۟ j�2�6�����T�6���h���R�#ƌ�v6�ӫ��q��-�Е*T��rY&A�zZ��f��ٗ�z�'O�]�t �ܫ�V{;��w���`<�S��i���n+�����"Z�g�YR����͚r{=����[�+3ِZC�ۗ�����]S�%I�����,�)��VS��a�;:k����c�܄�.]9��\��p9��"=�A���oR�m}��{w�n+Y{���T��f��.q�w��Exw8�D�ψ��Kg�6��YN��mR���rz�3��ӘĢ��v��x�����ޕ�VN� �îA�H����K*��4I�f�����GWt	�2Z���e��Լ�*�ÔoK�j@�B0�C���Kιh��ԗ9n[�)�ʦ�kss�ұ�-�X���=�����AP�ƿT&��K�\�1FϚo���A:�5Nm}/��V�`��iW7��QO]"`�y�!�;7*�D�Ǳ@�W�%����+���C�pB���qr`Ƿp(�re)ɺ�����</,U�$"ԯWnLpV܆���1V�
���B���sm
��/#Vw�Et,�tn� ����r����1	ʶF�:�r�Q�k�I��(eb�����������7]�Ɵ�z�w�"�g5@)��z�NT��6����pg�A�[�2=9Y\Gbβ���˘��BW$���5m�����Y��}� ��5��u� ��u1�ﾲ�x�~2 ��",ڌ�n�'�"_<�=X�j������wOE>x�d5%i�Z�P��C��6
.�	'��}C����=4�I� ��7;��Aۏ��\z��]F�>�G
�&i�!޼�Gq��xO��D�{ǹ�D��������qӱ��Ov�+k
V�5�,	L�LyEZ!���;��P�!��~ǅ�^�Px>�q+O�I��,�/{�kڈ������Un�;�ARy�u�B�K�o�
۱��h\:��"�9٦�G,���#1��ǐ���Gh��3vn�x ��V�I��O���oylc�>����԰�^z�.�݊j��t�H�[X���>�;�jk�mp��2B����$�<���ﺠgv�6a�a�a.�7�c�L�~���q��d�[���us��٣�s�)�|�Y�;_�{�l���}��ޤ��W�o�	�7{��i�A̶r'��d�������k��̏��RxnD�� �Q����1�A����'DoVhI��ݕi�Ç.�%s
�� Bz�ۚ��MgmjUĴns9�i���q�ݺd>�t�j�����v����Ɲ�.m[�)��,ڹY(��� M0;��o2���/2A��;�_\�o>�-����y�X�uY4?_�-8;VL��R�����n�6R��P��(�P�+�"�q-&`�y�n4I\f��6K�{{f8ĩP��zԚB5�y5ojْ�2�jh���E["�}����1���P���P�* �X],��㹣P����7.N���^��CA��A�f�*P��a���%*{[��^6��R��"+h���y���P��6��[����[�|�ݻ-���5���Vv�t�#V��� ���+��RyM
�W�%}��gT0b�\� p�G�� ���vi|�dh]V���Ȅ'b�tr���=�k��N����X�h�p���R2c+S�o���w��Z�7]��<��?j3e
�%�����GV
�ǂ���S�G!�%vֽj��!*��pWU��Gx��Ŧ�g�|�f��}Z�Dh����M+/����o8��6�t�s�S�P���C��l��fit����L��@7R�J�9B�ݾ�X���	���[��:�aP:�������*PуQ�D��[-�w����1M0���œ����T�E�k�9��f�ݢ�!{������?S�A����.�uD�N��J��� $�^�
/5i(��ޅ�j�Y$q[lQ�1C{f�W]�v�9��G���lt����6�PgFYvDM��PU�P�Q�#���a_�8�-ݐ��5G6��쪱����s��{$�41�w0G;|����gw'ֽ�V��ٔeG�7%�(�:�㧋}<�No+���H�<s�u)e��^����`�x��������Ge���;S����uƱ{�(#�ao��ޏO��m)�����GGn�M��j��
<���v0�2�ԑ]/%�S���F�ge�p�`Y�pNv�E��y��>Y�bf.��ū���
��a&�zWW]�����c�x,б]@J�������YFΕ�2윃���O�z�kKm$?�	�R��Z�v60ۛ�s��J;8�ZIb%�:���gp�wj�z.t�FK�I�X��SE}����9��K0m������ǀ�/rjYJ��>�]}M�˕*�^A��idew�^��V���R�D32��w�9`�׭����M�U�WJ���Oq�q���1��өV���ğfd�Cu�_nЉ�=��7�Ҡ}�V)g}��E��Z<�4�vn\憧��V�Y�t��>V��q+�v.ݢ>|��J�q�wy9q�s�u�Wq05fC��%<]W)��a�gj�f���:a9�7�8լ����;8��i��W��w���U���L�`�r]�7K��]��Ԝs�5��|_�6ԥv���c�N�&��:ؕ,9@�{Q���o�����(Z[W�p31�ot��$1�/��bW����K���W¯����qbec3����"�N�V���H.D��N4���'�U:��γV�1�Y���B�}�sd�Ҽ�7�[5�R�}I��W�԰���*�v����t��]�a0��ON9�퇫1�d�P�{��#�[��WX10`�%����G�qn�:лh7�]`�U��e���幮+D�9r9���X0���R%��Ll5)QӀe[��'h��473TF&��/q?�6�J�*��o�*���n
0�qh�����9�&�.�WwL�`U�S�<�0/Sj,�4��U�>�
Qk~�����d��L��[�z�DyԾ��\Z7�13�H��|ٷ"]��o,P��IL��Q�se1ݱԐ�ƥCm]t����Q\R�j(,��E�`q���u2wi=m��2j���{�A�g�l)7n.�>/�9m=[̯�Nk_�䑮v�1u���l�j�pc{՘2���C&�%6�{��fX����R�]�w؍�<x���� ���~C�[��}؃��b��*ܓ?g�r/G=��m˽;�;Ӹ�+9Q���
�HQ�]i]#�����Yi���ǈ��]���ɬP�5�e������ki��%#q#�]�<\f�7b:�N!x�2�7�3�/oE�py���
6�s9�nWj �<~��T�5��[/N���GK{�����˵�����|�/���	�u��v�}�붻S"��iV�q_w)!I���Y�g҉���~��z���
��Q��eS3*-�,Y����`��
�c��	��b��鲆	8a�5��vq�����F��vv&�����g���|��x�Մt�:��7�͍���:����s(��ﺝųQztX����Z��o& �S���<-PZ1�D���_0�ôE�ɽ���M�7m:z���Pǲ�L���.��d����d���o� �}���8���xn�r;{D��v�Y�v�y���+����㵽1%�31]��or�p;��P����]l� O����r"n�b��<xly���A	�HO�$]k4���3:�h��w��-����8P��eN��|j3<��e�5�Y�Xq&�d���ff���_p3��wWq�ص��&��q�;�c��K*2�H�*�dR)������>����M5EjgQ�6���!�lq�mK����jC>�˱�)D<�����	n�Y��t�i���q ��S�ɕv�7�TN�5����z����=d���3v���n[����3����;����+4��B�+9D�V�y�n����d!���.�\��� �2�J=L �^���8,-�p�Wv]�=��X�b��m_6�$��L��uʹ�� �'��wϷ^<Ǟ�"��Z����ʳ�&�j�i����[�X����4T��[���j�l�S	��eh���qH�k+���^�q��=~~��r��*T���j��q� �Wu��@�2�L�u\t�n�}�i��fv�4�l���+Z�h�z����:*7����-�Y�����/�"�����Y0oT��me�r8ޮ����Սd��[�Q�kDeO�@��g]�~�WykKq-�/�G���-�{���ᗳ��jj#]�`���Oz����2��n�����Ԇ� E�o.��ۺ�-F�¯����ʵ����s��:ۻ�Իč�N&�:"�ҽ�D��f�*��G�N�)Zj�VMm9c ����U3��p��f_�%NܺT~�p����5�F���=�3�W ���:�V��j��N��&2;j�́S���ή���s^	��rI����^=��w�ǃOG��㲕=�Z���\�x)\�}P%��	����|����ϟ��lll��1���������C�S[}DW��؃7.�`�5k�Ώ����6�ːۢC�z���)4^RWZE(*c���L���Ӏ�*��+��F�X�
� �R7�c����Wh��1��r\z"<juͨ�=��<�$L�s[��O}F%aK��@�Jb��k�򸍊{o�
�#�a�͕�n�s�,�J�������y95�{3�n]�t�"����&^�[�����Sxцoh�+su��Dc��(ܛ���
=pJATǨ�;3�˙ϋ����vK�fY���Z��+jI���hq|	��ö`�a@��]@"L���m��.�����0�fR��*�4�=��.s�^�/n���STg`����%L>0�I�z&'6��b���w{hwD���$ںt��O�R>���n�
0gb���y� �k)�ʞ�pptt;(���uְ�����+4S] �ܝ���P�����Z�)q"��Lޱt@�V�����v���[\�T�(36�5W	)чh��WwB=�����n�69����۔�s��r��5��ܣF��a�[5s62���	�%|���-�ɉ��ʱ�B�B���qʴ���v-���oid��0`Ui輰A��@\�"K 7k��r�8躛*PHK� e�T^���z�ݜ���T�k�+}]M̭Xo�u���H_tҚЉ�u�ڈ��*ǃo9w�u�.mT�A>���+wR�I���^ͨ�ho;OB�(�H{o�W��9k28�m�:����]а�S_d�>���^Db�Oa��wd�������N�I�`�������|�g���B{d#*3���d��C-�]����p��w3śq�x�{j�0F �f�d�)n��+!��(��������n��r�P���7ٻ�6�抹{SR�0K�Y��|����
�](8B�]����J��;��yȒ�
���d2�Աb}:�i��i��`Ui�%w�|dV:�<Ҷ���5�1���4͟%�_L���xB:�u���Nnҩ�n+Gbu�4z)_��5���<l+ؚ��?��a8+���+���2�\�A�*a4x�ͩX5�O:=�JT�<�y�#o�o�з1y�}[�K��W���J�[�ڍt�x���m�w]��f�sr���xt�	�V���VubL���Ѻ��W�=}�U�}��8�����];�����(��w�풜RJ ���A�(��9y�2��O&�J�u�,Üi�,|�C(�ޣR��֝�8*2��.���1i�噢��'V�ĝ5���1�:�d�o���:H��Vԕ�F�a�K�s}�&���_Cy�;Z����˩Y�9��!u� �xԽė��L�D�398�ݢ�Ϋeen�h+��d�ڶ�^���}�y�^9;5��G�[�Z'���KM�s��l��37uVb)�N�*c��.R�ti;a���No�G\�3f8E�O7xdh�a������F%�#/O�iz��9X	.����o�%I<��hm�	m��f�y���I����i�NR�=(fۈ����lu���*}�lwG�vG+�k����M�\�ޤ7��B�r
iAj�κȹ`)em�ۤj�˩��&=�g�v��hk�_ay܉�΃�G
v5��Ӕ]QMVo���R{��[�RCݵk�P�j�s�e.y}0�N���,%K�{%�d��Y���N��/2T�EK��.��t���(�ҳ4=����N��=y�`{wn�Yo'�l(�c����Y[�Z��I7��TJ�|��q0�:+��X��M����"�}Z3qMw{�$e���utEߴ�Ս*�Wo��=�ycF�"K{!PB=����x�zi�m�������t�v4;��
l:F4f#;J�';+]gxg�H��6w�:8�_n�ߥ�|rY���:��3$$��(���NҼ'�%)����:�b�y�w6�+E��s�(Ioc97��9�]��0'-�_�٪?�]�1��컾iXb��s�ܷ�gl�a�L&(S��L��7�lڄ��	���!gN����o+��׵Qi��t�+���ʖ���9m���,j:�$l0]��Or���"������kW��E3q���w:�ܘ��-X�(ѨY����9�vu��ؾ7j�g������ψdr�Ʉ��[��O���@���_�y�E�V�ʽ�n�3v�ɰ)���<������{Fw��XƠ��}��cGL8��컫_z�A����p��I���=�E��Zy7�v��٥f��:x�X� �Sn�ݖI;3�g�@��(�n�*\��*`a����*�T*���>Vx.���\NBz�^�#`֝c4����rV���_Ҿ�]!-�P��H;�_s$h�hT����}��T��bR��ֽw6q��>!^�0F����7�9�V2ˀD2���m��T�N��)���Η����Zq�ׂ�L��ɳ�K��y���u��O�R�AД��K���^�
cu��W��J�N���x��v,�A�<�]�N��f.��w�i���u�l3�]�Xf�B��l{��Yr���Mv�Fް�P��	d֥�yr�u0�H�I�+�
�2����n3vl�J�?F#4츓�YQע��l�5n{۾�-f��瑵�n ��d�dZ�/���ھ	Che���W�:/{5��w�X�*_v�(�����4���5�b\�ۓ���:=�ǧ^6���׫�Eh`�M9���:�QՅ%}�`���%�j��]�Ho#�S\r���)��|�@�����sY�0op�e���l��@1�Zf(vw��.�J��o1��"��Sr��l�|sh�
��1oD�7j��A��Ƶ|�e"���ؕ�}��c4Z8�	�u�5n�OO;���K�<�k�-����e"�&��4Qe�n��O�n.'���&C���ogO~;���dev�(�tmh�b#5kX7<W*/m��狘�����e�xd�}�nl[�9F&�͖��������գ���+�L=�9�}�>� �T���m�\]�f��؇D��V���j��w���U�۶��8x8=Ձ3ʋ�l\�e
��9�_s��U���b���vM�
�/��@���k��#pq��Aܕ?��5����A!2�>lJ�{�c;uf�K�iyX�M��%�K���mV��738�pO�v8"R�*:�������1�sBX�������u^YA�Z;�f��V^F�Ҏ�&1<z�
������n�u��~�]�]�]��ܚ�Q�IJ;*q�dP�`X�����&�\L����e�3S�Πt��E���S[ۣn�F��0#�N�i�
^-˥���m�6�.
���{�����jzS�f��.ۨ�Y���W�&�}����ָ��Njgri�ҚNv����ؖ^��͓�=ޤ#�+m7 ���s.��W{v�&��;����[���),���yˍ��b>c
J���`���;��&�e[�6�����e�>v�Ȳ�p��*�-�$j_gEX���v�N���L��m՝��C;Ĭx���gd2c�{��#}�XL�zǏDxQ���������a�('+k�34�G3�aW���7�i��pX+�WjJN=����g'�R(����	>�������3��(	D��!���yN���e��b��yycAރ��)�V�\��ęt��6����άo���r�cs���v"�\Mɘ,��
�n|�����]�{5>-�9����R^���>/Zi�r�%ۀˁۛX�:�9/���k��7 n�<�ESj���vx��J���.�fC�����̄���h�J���1EV�|�eQ�����IhδÓ�-�ԆN#��5��o��e�,��q�t��6n��6Y���/��a��e�[�=���Z0k�za��q{ �����,��r8:0)�2N������G��o}�!F%wQv=��X��*��4�������*km�o(bɚ��^�T�%H۩��7�Wc<�����yf��x�A�*d��	7;F��ѣ�^x-z�=��m�'k]\�=�i�Nn�#j�$p�{_b�Q�8�I�A�L�S@D�L�|��{����7�v���e\�h0Gd�M�8w�^����cשp�3Y���"	�B]Ekܗ;=���*Rr�kY�`g	{��,ʘ���q����4>m���L�G��dK�b�o��\�M��w�h���K�Hv!e�u:p����m��{L���/d��ƃφ8�Gt���� E�>��wJ�\������	�=�׶(��)Q{���H٦���� �ewt���`�;V��}��K���I���jI+��{bE����nW"��e�oM���L��^X8�>|����n!ϤjM���)��{��񵓃�:��(���v�dT�6��,�ᛂ���'��tWZQRFT�nԖB���/q��f��N@B�19�ˌp֑r�S;�{�P�y���@>w����+��X�矒�y!G_d��B�Sk#�4�t���J]z��Ei�û����{����!F�Ft#�ؒ�ͤ�2m���fYF�=�����tY��m�%e4[��@�.�C�w��ɞG�l��qO�G�W����eԭ�*������+�]1�=��ؘ-D�{5p��t,����r��X�Z����ʔwXj����}��7�xy��[i�3�$n�&�m�0�W��Z@P�;Н�������c
�X���a��/�NI�>�=uw !�K�N�^;Cj�)��$7Y�qa!Tɻ�?\�O<޺��aZT�VC��K��=��KW{SS��h{�=���M���������:
بk����C���j&9����W�x�7��@D���!݋�f�ȫS�+'2ݍ��To�ub���I{S�_����@o�f���=��>��/WF<Қ�y�޷�N³O.���f�]s���u���U�Wt=w@�;v��k7w8G*vA��b�[�d�Fi��Yp�:������s�4���PIl)f��6�,�)�(�nP`QGN+�#��9�{P��\�ޛ��؄��z]p<�{&�t%NJ�����k}�^�{=�=�"<Wm]gC�wM��;OD�-дF�	��ݛ5�Mj�s-��JAz:Sʑԗ���m�iZ��%�u+e�Cqꭠ7Ɋ�V�0Ya��7�z�sr!� ���[c�[Ս�i�uؾ��yEKڈ�V�;���6W3f0�V���$��"�s+y�q�maZ_lOw7���)$h�ֻk���1/A�t����Z��J�U�9��r�L�aå�l�]9�ɜ���[w/Fފ��]K�����y�y����k���	B��K|[8ɮe[�&_lšp�a�H��fI�pi���0�Mט.e��wNV��a��V�k�
o�	���!h�Kظǈ��C���fӵj�ϳ�?�w<�и�z)���`գA�\�h�ut������8�K�:V����v�b̕Ϣ����I�8u$ M��М����w]�RL�jlǿ�Wko��4�jD�����I�S�&6R!�� ��\�D����s�3G�I1:�V�^�펪";�0���y���&5���ڳ�Y�G�j؎ƫ�������sNŢ<)�M�<���P��s_s 5���������9���JK��._!������+��CnubUl���3E�&����ޖ���I��WGÔ�L�7�.��`+Ym./R� �q�Lee=}I�.}��qE�.E����f����s��Ozۺ\<=�]"�ɻ�m���R+8b�S�����ο	�T*ކm-�R��Se�x)�l�V��T�tt��F�ڛ{�z��mY��X�d.����<�]�t9�*�0��l�� �R�:�5�[��wݫw�ݳC��gt��H�*�$��p�Uuz��Šk�gR�gvc:��+�k�uGѵlĮ���fF�5Uқ���a�̢�f�d�����W70k��-�]
�k �,
M H�俒������/)�_[(r�׆&¨,�ܜv{0�X�x*����6u���G�J1p�\Sz�:R���f�i*��>�䏛ݯ`}<�L��>�ȷSZ.��lV�FN����x�CJ��	 � ��	\:��,5<Y���}J�s��([B3y�� ~==�}{r�M�B&
�;��pК���x��ov[O"�#�A]Y)�Ԇ�fՂoVM�]�I�!�]ы�mG~����g�(x�ãk5b��g��ԾN��<���}գ8��Ì
�B�s(Y�$wf��"u���4s����*���#��nP5���ͬ�-9�H16���o�4�3��޼�7ᾇ%b��[z�R��&���Ŝ���'��q�Po�!-s���7������b������N���:ֹ�v�v�{��i�%^����{��!�ɢ��i��]�w3:|Ӎ�s)�Dm
3R�%��[t�kh=�xܙ���G2Rj0k�	��z�K��w���TZ�r�w�+�%�k�ڭ�T<Q�>�}N"v�n__]v�sK�}z{� �z���*r��`��B�Af

ގͬ��N���OC�S����
՞�r�躷�@͜�q�+���-�n�n���yZ)΀���Mwa-/��s(�[δ2jM.��D.fe��hຜ*��Q�PS���K�¬7��T�EH�(mfǃ��y���U6�gvEFy>��!K���G�����gQQ�h(!��n�n�����*����xx{�x{�~��.��[ª*s�2�q�&��;J-c9�2�4����e������+���p>�,���a7�7^]�ޥQq�Ҷr���՗k�a�d�2�7�2���8GM�I���vޠh#�ޏO%���H֥�J��	n�Si�s�����.�+��Y`��͂y�N�^�c�y��[��b�����u`L\�]�{��^{�h���sG��X�ז>({S:��o���sͻ��޺�'�$Jh��XZC��)Է�(�����b{N�i�&pR}��+9���]�;�53���$�tDW�T���J�Y��p��K�g�'G����}sps��B�F>t����\��
�p%�s5%wi�p���\�Xie�VL�ּ�Z�3��-���{������ߠ���Pݭ��[_�-=>�T*眶��1f�ЪU`I;4�fu��\�gn	�~=�����)�kh���Փ�^K�M�%��R��cY���c�'[ġS%>��3��^��x�Ezv���c�'̦�]�c�S�	�aP�.w9�ʖ�E�C�c��.����X3wf���z�0���vΗ\#��o�ͳݒ��a�}��qT�T.��T��U�ǫoz�$V�����6#vUwWv�>j6��p�I&�#z��c�/�@���=�ެr={���j�d�P���5��P��̴��f�eDr1ۛ�}w�B����$�J�+��hAʕ�'$��F���xAl�Ny���*G�븑y3�T�-wU=J�(� ����v�unk�.!IĮS�E�����eUG�{�:����8�����R�չ�S�.Ua�v�E�Z9x�@�Dz4��X���U�N9$�Y��(�B�j�K�NU��Dk��Λ��M$�ң H(�wr;(������n����rԹT9%fy�F���p\�E�uhS���Ns!
��«�s����!ӑ*�N�wE	�Pp��u���B���(]ݹ^��$瞦a™�x��4�B��Q�=.e�jY�V�j��HW��+2""'S�s�tr�Eg'I%�A!U+\�9�p���ww	�����J��(�/\�T�(��W(�1��#��@
P�
}f\bd�}ݓ)$�y]�1w�X/R�2�*�Wj���Fm���"]��$faO����o#a�+bӅf�Ff��ﳙ�&t4D~�R�)���\U*��4Ӂ5#kp�uT�r����	5�7��y(�^��7�k�ĳ�\�<�����c�ﯸ��!���X�b�|��o���}��ewy���l}���zf%�j
�_Pu�Cѥc�-�O߄J�� �xi�!�����q�B-/�}|�Jヺ"�U�H[nm_�	*Tz֤* �N�[���,Psѹ�;-n�b���'m�0/Z�aKUE�K�gr!��L�LV��;ꂮɛެ�|7�O,c;�g^�_`u�A��,TRʽ2\��@����3#��w�M�ϕ�٦�W:F��+i�SQ�\�Y2]��K���`J��e?IiY
�CP"�	ݣ�2}'�)��s�)�V,�f��ķ���W���u~s�-IZG9o���	نJ��A��+���=0�D�X�c�p�s�t�6#��}p���t��ȹѐT�c�������LikP<���w�cZd��{��y�4�/:=v�v�˱W������#L��J��@�@� �.�T��x��Oe�d��X
�c���%���7�n�������Wi)d�j�w/s�M>�q���EP8�0��M��J���?�����:Q�ᒈ}!�n;���'�{�0�݋���Z�Ѥ�T����n�N��]���5��V+ׄ_@[w|��co�مrS����F:�g��i�0_�k���Iү�>�a[��]�LP����Z7j�v0��&7I�5;��Nx`�51zP����&����@�j��@�ٽ�kc9f�E0@݃���Ju�g�py�Tb�W`���2!ˤL1+V�]uJ���ڂw�%�YV��\H�#��ȍ$\��Q��H��_0���a�u��"t�j�h�j7��ԁ��0g S*L�J+���qzV�Q��3�/�F�`��Y{��ZҰ���������dɶ��C�d��%$��5c4��<d뷖�3|�&�����l]�Q��E���Pw�>=P���(�g�q���ӣP�a7`"�Xb2)_��t<�V��]:�h�d-8%t�1xPc$�A�O�25:�>�_��*9�N�N��.�Z\�vҝޜ��{��YUHklm�j��� */]CK�Fr�f.9������_fk�gbT8z������H���N����!��"{*4\L�d�6��!�8��$�٬�\��Wj�Cu1�U����,�-�����8Ew�w}�ȅՃ�)K��`u)$@�\��]��C�8�]W\r���ל9NVȪ#0��wW,�6!���d.�̮�hj��D�Arw��.p��i�����"�1po8��},�p�u���y���huW���'�.��YZ㧝T������] ��DrF�_Z���{m��2h���{\[��V�f�Σ���U���I�8{�	h�O[�U�[�m�9���>}���Gh*H�[?'t��-���ymt��%��+!b��[FPf_U��.z���� ��U�(�[�(�R��W:c�|!��;P���I� o{ٶ�4���'����t�d8�h�ۨ�t�p�p�X�~�}��C��`�kn�^�|� ѪO+N*�2�!��>$�-ش�!̬�
���D�q���S�w��9��zg/#�L�l�����{���	���t��e[��/M�������ĥ�
���˹��s:!���k��A��HOK9�U� J;���qYוa$@T�1������q3�\�c+��ܛ��8Cg-N�
iL�B�e?w�oM׹ؐ�^xU���Yp��P���.5��k�� �5&*N̔�F>�V1.̓\Q=Ѯ���UQ>�x:<<�a���8�ܞj}i6-��w_���S��
8�fk��>˚�YG��Kw�	���&��Eo1gD���y�]	3w(��j�ؚ���R�Vl��iM�:)\^��X{�l̡���3pm>X�Z��MʛպR���pq�i*R/�����_Gقڨ�qK�j6a���!rwr/�	��[,�Xf���nVV�U���Չgc�|]�� ��Rx����z�тh���S��fz�����_t�f6r_�z�24>�v�B�a�q�c����B���h�1�0v��6ձs���6+lD��t�Wk���&\%_v��\��lǳ��HA�O�|�έ�܁����]��?:�u���[f	�qW�l�d�1l��j��Y��+�k��8p�/_v�juX��{sR���Q\x8�T�����a�֧�`˖�(�\c6�Vq��`ᨁG�4}<�k]�X�ov/C�..U�Q��WӮ�+4���k��x��E{ݮ��(b�bb�U^��=�Ͻ�d���f������\෭��Ϭ��T*Wbn�c�0�=�f��"�)גe�B+�K���%��1rKJ����$V.��f���B�O���;q��Y��h�<b�>��}$gBo��d���ܝ#�xV��ά��P�^~m�蟓-�5n����p��<�:�T�u�ֽ��go=ܪ���->b�e*R����#B��Vè��U�l3g)�+���i��/�t�a�Y�,Z?�N[����mki��]qR,��E�e ���}�f�_2)N�b!]�G+�n�_5j���M��	������[!׽��߼Ƚ�p�Q E.�8��"�H�X����lO�P��R8ߙN�����θv|��g�{)�P��;pꙐ�b�n}��xSr�G+8ä��iJ]4%��3��<>�k��2�k�k��k�d�GV
r9J�ZN7��ֶ��Kxؼ%
YƜ��"�ޤ�D0��?SJ�-���Q�XP�
�3,JW�!Ϙ��訊_i��	��ʊ�պgL1���E|�屐ګ�����MU��m�ns����5:M��uĘ��^,c�<W��*rrb�q�Z�A�Ne+�`]y��TD�t���,2tE��w�#[���C�؇uCB�V*
����b�?���9JU<���V�Þ�UJ'�ޔ��[��
�xX�n�Y[�્�҄P4t"b� �J��;��ؽ��O�V�qT��rt"v��}z�C-T1���n�ogV�yS�"�Ö�f��'L���K�Y )pf����5�b*] ŌN�2%w���!�T��i�����g��4>Ω���U�%�zN��݊��#���]�:��Q����Ѭ�aA�=��;G�'��K4�������f�^K��W��^��n�s�7�}0��-��#V��(���U��h��Dp�*Ūm	��nobi.=��5�M���0I|tN���	�����:!Tf��j����DcrG<�n{	�<�uR\uS�y�˗�R��T�����0�O��IZ�5����z<�Kdyb2wT:�t�;�7ɾ���2L��E�4G�j0�Ҧ;"&�GX6LO	:�(�R��^�Mb��g�j���(V���-4&�v��5%��>!���tA4��@�� 1�J���qIF]�2u>�ns�Ԍ�fR?\c��qۯ���0\CZ�"�8yFKeEyTh�=u�����\,����yt�w�d�cY"�;-�݀�DV'\4c���/J��iT5���s��[�|��b�@��(��.�5�,����Ů�W`I�AC�H�����7�0�]���Ϻ+��W�`���Q�!��#gd��VӣWJG����|�F��D��#t����
8(�y��� �'/��P��C�*��Eq��<-��-7��O�h�=�6Ze���]$WQ�ݯ�j���)�%� k_=��Ւx�<��()�ƥ�y��u�j�8�2]�Ys���` ��>2�Ն�ܺ�]�
$��uϑqR�fc
-[���������+{F�K+f�����W��В�*�VV�ٯ�ܔ�T5��t]c�Fm�q����Y�/`�dzv����k�][h��G���suH����`�}��'z��t=4���drw|c5�̕q���YF�4�3��L ղ�fI:Hgul����i����*��(L8/��|M_٪]f�Kێ��-s�ތ�4+��׷!5�U[7�8[(�ۈ3�L�a\UT=0�sc:��]C�R���Y�W��q2��j-����X����>縃���wl��_����c�T��&eLi�rd��3��Q���]�Od*K��'�����$d�1�M��q������{w���W�����ϠX!If�ڥ�l�2���u�-��+��
Ϳ:�U���"M/����<0���M�!x��Ŋf7DE}�|�\�Y��J�����OO��j�YԊ���u�u����[�`؍K�Go��7�(\폮!�t�c��D&�a���'��S��ۉ�XD�8��O	~+�L������ۨ�-�	
K5�ь}'_U�.����'���8���t�:��f�}�� L�I9�|}���]//:�D�	A���`��;<�߮xm/ Шy�Eu��P���KT(
N�c�e�N�Z�B�͔s6�*�U]ll��e��t��K�H�ԧ7Ƭ�F�������Q��Q���`*�{z��N<XD��ɒ��0vT�/�V��2�&֚���9�Qr�橧�\4�g��J�1p�>ڡ&����y+ϋ�����~�"�Q�y���#�P�(��lY:���%���ꐐ%�����'B�]m���={�'|�
ߪ�O
N�w��`�V������#�D�H8hiE*�{)u�-�Q����Z�����"����/M����5&*N̛����w�%��Jiy�VH�:b����S��%�W���`�uF�^Q0ƾ���U!��7,&�����t]a�9�����ץ��^'��^�t��K�0�0W�6��bh��j��%!keu�Y��k�����������i�����q��dn�.��-��S1�4_l�x*�i�� ���WA���Ճ-�g��A��_�lg�#1��� ��ΎȈ��T�����:u��?Rt@�*�O�J�e��F-�����9��F0gy9t�k�}H�bk�����mFt8��	NA�aޙ�"��e��鲲bs��"��HX�-��3�ܑ3�-�r���L�Ʈ'�a�սs(7Z�yg�i���ݸ-���K�ݸ��th���[Ar��/R8AI�����ZХ8|�2�6b�z�����c*{얯I��^��P����O8qg.M=ܤc'h��%ė�:M�v��=r��G�+E��T>T�S[�!��J������g��pj�Rc�&pb��e�s=f�F��0~�d�R�=.{�6>U�v!`��F>c9�2V�뽙}r�x�<2HV��v��Mh�h��	3J��q�=�!�:�%��/O���ff�������5�ծq�B�u�=j�5��T%�=��O�`Tb�
zjC74�8�nK�u����y���Ea����՜3���+ð�7$GU�de��f��"'��=R舕U�>�Q,�R�n�],�ջ���4��c8�غ�v*vٌ6R,��	����3"��JNIEZ�r�bvs;��^_��:H���)�<��FXv��Mu��C�����d�u�1I�#��Fi璷.q�{� 78OW�f�=�+�:����*�z�w��ų�~iK%��Ys��8l�ǆ��Rs���0E.>'_�
M�}����N=U��n��\��ީ��.T�Iz�1+2$�Qi`*�����Pv~���~Zh�u�^փ�y ���uv&n�Z��<T(��K+uuBv�����o,`N��9�I�U�[haa������l��]�q>��ҙ�H �N)��υ�z��5�eZ(�-I�\rf��r�ΰ��t�锭oI^��je�OS�4�DT�Ч4�;4]I-vN-���
��U�:�9���ۿg�Cf׭��ZV*
��j��/��nGMe�"��^��k�)�Sd��ޔ�u:�#���es�����HŃf��QN���(��wJ<�w�V\��z��VY��ON���Z�c>����sl#�oZe�b��4Xg<X;��D�g��+>�ƀ�eV�T*q�t���j0<.�ŧi����r��]�p�h�9�^�[Z'�^�_{���v�ҾKvS���tB�;�Rj�P	`�v>����o7e�p��5���{����ï%��^X�]��˵	:]#�.���W��G����jV���&jV��ǯ��R�p��F���yx�ڇF��H?bҒ��P�:�G���%��ز��{y函�
�r���	\��椲��������i`�<k��Ƭo;]���W{��t����?\F*�g!ۯ���0[Z�"�8yd��T9�!ʎ��P��Ӻ�X��Ӆ@1���������8!F'\49j�b�����G�_&�ufz�|;-�M׻Ї,�▞�[�.�C���)�;����!u�s6�Z�S�+�����p�7ST����N5�=!��d*�7<k;��%�r�|�,�,�g-�W82��$��z�;�{��s��礬G}L�3�g(�x�U�^p�
&��@.vGI���U[8�����ܚ��6"��{�Sɲ�S� ��B�U�]���*�8rċ{������#IeѰ��QfB:sk�pch/�2ʗ�,*j�ۛn�klcBk�Wz�J&tN�pW�*:B�7w�6���T۴<���7A{M/�>&�t��[��x���4DܮZ3V^�7T�Z'U���]��<mY��n�6��Q��hmV�M�/;��bo�}x�-<���Ǡ�@q�l6^�������Iǡ."K��5���ɹ�k�#_S]mBu�t<�UjN+f���W���͓��]@�r�<H�Yܺ�tVpoe��������C��On����gh%���>�Xhv�A�Y3���%�j�����k�@췲>-'����$ȳNI�����f�BNʻ�%R�V.)t,>�b��u��:�qQ��oC��5�G�yB�n�Μ�r'��7h�1|��,ۼ��ܺ�K�ƪ�co�oZ��r�K�����8�@�f��	-U/���^.z��C�m�Ͷ��g{��(����Ӑ��z�
�3��.� ����n"	��������]����J$�{���	������$�!E��u�;;q�kqB6����nr<ڸ��Yv�Hc]�T��;��)7�FW=�_�Q�͎jVe̳�P*I�@�^:�0�B��O}�cp�=y�G�&k/�l��½�^�=���[M1���vuSܹƣ�}]|'��o���[e�	�����h��ț��S�f�꘎����e�{�=嬛���u��Mx�~^퍈ZV�b:��mub<3�v�0ɵ��e\(hռ;� 52�f���	��%���a��0��Π�<	Œ�_�T����;Y� l��xu�gAIp;�J����H����3X�-�{F������2Π�*��K�@`�����+Ռ����Rފ=j��ê��DJ�ݻ�\ze�f�'yd���꾠�K����3�a��*XVY�1���UJ�❽M퍉�tb���5�_s+�$Zi[�{�ҫ�x��gY��U�YZ��4�f��n7�C����gt���u�Rž��f8MZ6_dm��QVH^�nvl�}A'_L�ݯ�P��N��~�6�n�9�W�U�p≏s��e:�I����܍=�=���V�˦�&�k��B��f� Z�<}w�;On��L�S��v�]$jd��3I-�-��룛�e�#��K� ����|��S��-��u��:',O6�rZ1hf�Y�uum^8c0����&)�i�+��>�ۓ6�	�m�2a(�Î[��֝=Z�*T5,�A�N�I,�Cs�R�����T.EK2.D\�Un��J�!^H��V���up��Oq˗(��aUE��=pA�wB��rwip�ȋ�wSg��Qz�L���MN�^I�N\�wt�I[H�E!$z����H�Q�d�J=��r�I
�,0*����Ȯ:T�C%\������ZDEQ�.z%d,�R��2��U����Hp���*Ȉ����E�UA���j��<��r��E\.�9\�瓩�&U�b$S��Fa�):ʨ��Zr����ȋ���N]ݡAr=�JXY�z�y	\"��B��d�+�bТ�:Uz%��߯��y���)��ҵv^��9u)p��[�c�j���e�}��Z^U
p��x�u�˲Q�\7W*I�De1+Z�,�+¾�>C��K��1R�x�,r(I�~8�:�N��AN}�rra}o��������z?8�>;_�{>��0����}x]�Ј�D\C~��c�}�}�ʓ^7�q�ԧ݋h>�"01��"@����G�;rw��|���j���O���]�'
o��ߜr��~�ϓ�۷��N�}�ۏ)�7��޼�����}!�l78#� �#�&�ۚ�}7=�'��U�v�_x"��i����۝�����<���������7�'N��}}����I;��<�~���;��^y��;I����I��)��hk��$�dyJ $�ψ���uVF�ݽ�}5��/��"�DF��#˧�|C�޿}��|C�aW����)�	��z��>���'>����m�<��I���~��������}[rrnw������o��<�����C�>y��|����z�׋P��N��C�|D}��;y�m�ܮ��߃~w��o�^�{���7��?{���yL.���|����ǧ��_���Ǎ�P���?S��������M�zHg�N&}ֽ�z�����{�c�$��F�/�X} �>������>8�Q�]�� }O'xx���󿝤�y���/�nNT=��Ǆ�P��׿w����׽��;~~'�aw����yM����¸׸��\Nu/3ލW�%\yTVޑ�دE�}�����?��ǔ��9G����9=����	�]�ǂ��q��&��y�ǔ��=�r�����n�[���v����k����>\
o�H�����|�D��E���<f��f-�V��� z~��w��x��.�o������=���=[�zO(xMz��>A��P�r��G&}Cӹ����yL*�'��!�7�$ޏ8<}��N~�zR#����y�]��^hi.}oG��w?xBC�y���m��&��~�&W�oi��������Ą��X����8�z�����ù]��c�}w<�����`�奔�w����S�;�Z���F
>��{����>��חk�翇�m��(��=���~�����w~�n;rs��������~���^S
��k�}߼p|BL?��ޏ�yW|v��oW�𞝼<��k׮7�<<��đk�d{H�@^��7�{�#*�7c N�,ǈ+�X�vʟ!�d�#�s���/ّ�%\w����8�-	Wٻ����-�gh�n�{��ki��sb+۔6f��_VY�<���Y���s���?U	�����dq���o�%|/
��ͦZ�-�99�B���z�=F'}q���>m���a}q���ng.�������<���_�r�?8����9�������r|O��q�I���u�ˏhs��˽�&^�!Cꯤ~1�ħ��'Atԣ_�|q;N��˼���Ǉoo&�����׍��M���Í'�{o����bO��&�海�ޓ�����Dp�ml�Yy�"��.��1�P���|BC���F�99������N'.���7��oI������s�G�}�)�������zw�i�_|]��N��;���ohy�m�ܛ�ܞ~ʫ��O�����̜}|q�F��F��o��߸�F'ro矈xw��]��A�<8���A@QC�|w�^�
�I����7�۷'!���.��۾������aw�k����M�I��S���̙)�W1�Y�"�����h�N?�v�O)���������yM�	���ރ���HO����x������<[s�< y���M���(��&;t}��{v�7�����S�O���|JMl<w����ߟ/�W��)���{����߸��>���x���e���������˿���G�뷔�Н'��ǏQ�7'��xO���ߐ�O܁����t�&����.f�1KU�5��ᾆ"G���G��~�	�'��=�����`���~w ���'&zC��}���!�߿w���~BO_�p?�~C����ly@���>����7��o^��goi�|E{Ux�Qw�����r��}�"�}�����˿��'��x�:w�i�? =^�3��~��>���ߠ	h��ɯ�;�xw����߾������r���x@QC�~}}����V>Vŧ�*�罇9[��PB>�C�D��~��u�|�濐�]�:�}��L=�����ʻ��w�x����S󷷝�?�~;
o�O�o?�z�zL)��>��ޢ*P�G��.�=旽� �]d�����җ�Mb}���2�a��y�Q|��;I�����Pyw�k��M�����z���aw����x�����>#�l�Y��~�G���>���#�>�Z��y�������?�k��3����yS��&L�d�.4���oۭ�L���u�K�9sE��b-��Q���:B�j�����#}�Σ�g7H��3qM0��!5�;a�s�5z* �f7��O�>��WMौ��P6oe3������χ!$�/�qU'ҟv�)��/�}�$}T���|��<������~��]��}��9���=����\xq+�?�ro���8[�bw�?;�������]�������N��s����o
��D}� �ˉ�dsx䋪�����LG��q����ߞ����N?x�1'��7��o	�~�ǔ¿���z�?x7�<���yO�v�oq�<��ޜy=Ǆ�P���ܾ{�ro���z?!��19��V��7�ܳ�Z݊��X�������xw���s�O���
좇���}C���V�<}���ɹ�����n0���n��~����©�=�?�{C�<���Nܮ�v��8��9��H�Z���-�ٯ_�=�:��h��D��¸������v���1?�����ko�����{�xw�i7���x˿;J�����&��w�k��y��yw���뿎���raw�{OG�yO�>$H��X�h��%�L���bT������yC�����/���zǄ�;ӏ:��onܛ��v�S�w{��<$��������N�����Ǘ�Ӵ�?v$��\}q+�c��7�����|7V�jv6�M��0��������C��
~��?����q��c�Ą��㬦��!������ԝ�Ͼ<��	�>��HI�~�y>������a�ϣ���>��#�Á�`�=B�D���)��>ޝ;˿~���7!~���^U����矞,yCǸ������9���s�����t�aWe�Q�>!��X���yw��n~�ߞ�
#��G��x�Ie���Uq57��ZEp��ɅS���獼����&��px�����n=����O���}~�㷔܄�w��Sʸ�|�>]�;�����ڭ�?�y������>��� ��yD��3���v���s鼥��|�g�}��5#�aE�}����%߻��� |߼q�]�4�q����wA&_i������ rN�w��<��&�w����S�~�� ��BQ��w1�f�o��i�[�������.�i7��}}�\.I�����~Nq�į�}�$���9?�~x7�����>���zC�����o�=�þ������q�������)�&>��"Ǉ�H��i���s�.�]^v�γ��Px@�������������T~m���S���M��׸��3q;�,�����۲x������24�
��鵹����F�k@�;��+�z���,]�f,5���nr*��]��Xۼ
�c����E��舨H'�nZ���f`��A�h�,W����	�~XS�rnB@�x��~v����}~v�S���ӽ�hܛ��o����W�ۼ���Ǥߐ��$����_.9ߓ�~��;�����}�q���;��ʀoc#O�� �����{C���V��xw�s�5�'��z(��7��_>;�n����y����>;r�˽{����I����|zw;I�!?�����p(|���|���W2o�u�[�[�}Dhc�D������ÿ;U����S�;I��χ.�iP���&��s���x�N���w��~M��S��>��ǔ���9����c»�i���z��Ǥ��	2���ߡ�:X�EGm�^�\�iXd�C�G���>��ϫxv�ޏ���'N��@���xM�	'oo~���=��ޝ�<��O8\.��-�7����\�7����z?�x���=}��ސ����}(?7`�l���oG��������c�w������Ǵ'y�﷤<���~�����ې=��Ǉ�?>}|?Տ(I������o(I��������ޱҁ�!������7�
1�/L�=��
���yt?���D o�>2o�/Q��~��&��w���=��<;���=�=x���®ރ���(~O�9�࿏߼�1���ɹ����ݏI�0���׸<�F�� }IS˵ѬDH���=15ۓ�w�@�_��zbG�H]���2��$������&��/�o)��S��p|B~�rw�=|�����m�׿�>��aw�k�?x7�˗~v������9��������bw���<�o����fb}
;�B�|�H��~ݿ��ǔ���9޿[r�M?�?�90��AE����O���?���^��2�a� IK�^6~%�O}=�f�"O����ʹ��{���\��a8��Z�l�1꺇jej]���$�!_(E��	0w��ʈ�HN9��~�
���G�b�m_��K^|<;?�ݶ�˵
V��T��9-�du��)��.�G=����Ҽ�a����w��$�:�������EA��8���hwK�!���C�u{ݾ�:'�P������+��l�FC���;F��F�c�s�ҋ]!��ܨo���2��쪙W|;�0���q�R�b�⭙C.7�4�IY��M�fse�.����(�5�S ��C��CD0���&b�*c�[���6M*�']% �K�3����k
j��9��6dND>V��5%��4C����i@6����Ae*���
'O�����֟r���k9�}4�.�i���W�Kg�.F�!D���c���I�Q�@艓IO59�N���/���iCmF��Թ��*��-N779Ew��B�%�������A��
E>U�۔#��b�4r�m߭�s��V��샷a���&-��ɦ� �W.��+�>��D*S_���C׎Ռ�j�ۼ�;���{���p�C&�u��%�4!`t�I�(���Bf���u���0[�6��Ļz5r�9��z�q��}Zj��S&O6�yn�q�$�t�=3S�s�%��Sr�UR��_S�����������˅���񂽟x}�`�;�t}м�RG;��n��<gKf �0�`{CÂyO����l15O�59���k@��ѼϮc+�k�
Hʵ�;��3�*>���C�m\�jU�}��EiG���7��Z ~��5�����)غ���4��eM��b9�����pR�8��}\�`익���q�����9��-8��e����Q��J�a�����׷���#�`%�3��WUP��(�;Fu��bb2�5P������]n�k��֦���I���~�_*�[B�'vʩ��G�]�E��d���}*�C��q:w
��R�`� 8���3�s�q����N��8:�V#N��O�ZS��uٗ���hf�KyH�Oh��Y�g�BE�t�%�M5<��u���ͷQ�of��RI��X���=}���p2'�	`ۧ�Ī�+��|�k�����pܦVC�>�m�-�ּ�='�e�;`r��"��'�\F�o!򌖵h�b
�nt����t�c����c$ 
��6b�pq�Y�"�m����Y '���9�|�Hn�m�^^��C�^�\E���r�B�R:Zq�6�6������qԱh�_{��� FG��]�/��æ�Ư���s��u��IΉq��[���v�8��0��'�S�#\��^ym�೸�s�8�e;\�K�?c5����N�,��Nv����*؃=2O3f�"��ָ7.D�b��K�4��*�Ny�Rt3��h�Q֕�ݺ)>N���>����zgnَ���<�m�^�+�kx@=��w=�px�y�oR��'��{f�{���xe
�v�S�n:��.|�O;`�q�%��,^���7(Z��C�W�G6�l>{
 �	�b*\�:68�_�xƺ���hA��d��Z���̉1�Р��a�r^Bj����n'f8H����cx�=��5&*!��ɸ��#X}mo^����n��̽h��:�J�%bW��+�u�"ʽ}Jp��}w�	:�����{Q��]��5����"^�E�,��8a>ъ�\	�?W�.�WJ�o[64r���[:�6�B�'Nj�E�t��Ń�׍ �}m
xa8��lw���u.���AǷ�r>�T&�&�yz�N�T�~�/'��m�c>�!��n�h�s�����	�0E�@ٌ�U�6��:DoN�RWЗqT��Ϫe2Q�;1��`<�%ыgm�u�ӚhC�.s�<��G&e�o`R��L/ԗ�~��k��Mz�R4���f��2��)pk�f��8�9���|��RU���p��.��(]:P�C���+C�	@�_ �9B/*�2w�Vk8�Yzf�+�¯�:��B��G������^YVl}"���p.���J���Z��ts�J!���tֶE��Rk��2��W�H�*8�y�hT��9��fwum�r%{��-�z{��	�;�	8?#�e���?!/9`��7�k����f�\)GJi��il��%ٕ�\���z`�A=��yr���si�G�};��s�i)w�τ�p��z�}�n+}}��p,W�B]���p�ũ��j����p��Ț."���9t��5+����R��o[����D����.�7:o/.�j{-�9��P�p�Ҝc��)5q ��z�1�q�":��#-�#5�HHt=쬣��;�Oղ��E�߮�C=J2�5t0}�Fʏ��5`��x
�S��	�m{��&��,�~;�˃;��$g��k���U�=9P��Uj����]l!��,�`㕺�Fk�^�o��w��Dﾯ?�� 뗉�A*�]�i�:<�v�w��v�Y^m@@��Zbb�r���a�n�d��fX�+�9�#�'pH��3�aXk����׀b�_)�׫;��1�׽��Uro 0�`ak&���zY=P�M�]l8�D�97���}ԣ�>qH}��V�{n��'w�5:˝>�S#����W3�b���p���h�������L�c.���7�3y���*a�c��V󻂹i@Vsp䀺���"�τ븬��U�&̡cr�=zR��q�˴���E,�b�I�)b��B��{jw�&���9�j������i��rxRޞE^��������FN�ϫ}�J/ӗd<�t�r�@�f9J����P�J�[&ܑ�*?}}�Mڑ:��T��g�̢c(�8��G��R�!�<�ϲ�I���WE^)y_�梫������o=Җ�7Fo���y1�7�C@f2�B���>ʽ9�J����1��d��{�N��N��R��a���g�3��};��kM�Y��Y_XTuTuG|Z-�`I[L���u1u��$�L�E���Z~�*O7=��W.�1�����H˹D�$s9�U��Bﺟ�l�4�)���N�(H,��]�,��õn1p�W��^h`a�=��BT�D�~��Lvl��e��9 �b��u��`3��Bj+|r���4CQo����%��,
[b�GQ�[�v8z�B� 8g���)�mV�����P��lb}�w��ٞ
��Q�T�u�<2H�>��r���y�>hm�c��z-��y<�h������ͅ\X�Xw�����q7��0Y�!� $���_.��n�*���

xo��i�waS�� �}g��~�ˤL[1��P���q4as ��H��M~g}G<3<Fg^�C��CPl1��2Z�Im�Z'��r���R|��{5N�5�:
��&�ٛ���j���Ci	���B�P&yj��[�r��l�M�;�9Q�R��&E�>������K]wǡ�9���ʻ#� �k��9�eEqv�u�u��	_����"����f>6q�}�!_>B�yL2y�\�i�8_�������L@	����j���v넵�{	|'��:�l��z_��_֚�*-Jd�m��=���OX�P�]�K#�Ǐ���q�K��DP�aN�i�g_[4<=��˄~s��Q����C����f��N8:Uٜ�*�]Iґ��c�|X���xpO)�b��I����}��+�81l����͹�8�F����dБ��l�jԮ������CdD@�RZ���
��F	�{���zl���}}��љ����=�¥?f�@�Y�Uw�r��@�*�T}Ǳhqx���X�ݼ�"��vQ8�� M��HϩL6M�b-l���p����ܘ�(�2��XDK��-�[W�Ir�Ц�Ek��t�!#t��Yd�y��-��+s�3n!�p�ٹ8069�F';F�S�zݩ$���P&Pw[T�b�����`ۘ�6ܯ}��zY�Y�T�X���M�K}�f;X�]�XB��p<���[�|�nJ*����s��q]뻢#2�w��j��ʒ�GM[�n�aI�)L���:5'�%$=g:��=�*lG{�蜨%�	�wrǼ�[�M>��ѥG\��}F;SS��7s�̭�������n�̣r��kG
y�i�_i�oq��%��x�.�@��c��b�g=̝P>��G�9�y�	���X�+������mk��4s�L�ON�{c+Բ1��*jW�U����G'Ѝ;O��m2�v]1琢O��"�����u/9uԡ�qF���aSwiɴV��>7�v��i�ǭ�L�{��#A�a�L6��ϮuF��jY�F�{R����hĒCuv�:L���&c�e�>=B�`�����������߸�>a2��y�{(�GU��lm�/d�{/�����`��?嗾��*��u�3Uy{|�9��E���ʋ1��z����tf����C�¨��*�����"1���qͽ��{��3���Ôm���Jn>7�f���)/C⮔�j�R�{�WVD����Q���޹�YVP�Z�x�ϝ����G��ii(�-�kj��zյw��)��*/�7�ޮw� ��о�����K��<�X�P	�!@�E�4�Z�+������S�kE�\��'��=g�Y�p�4�fd�i\�
s����ɶ����Зx���XUr{Hr�X+�ݓ��ںm����c�FU��=���\�oӻM�,��:��^�V+��9o�۬���ۀ��0��H ���ejծn��լ]OV��)�0>�)���݇m�e�y�K&Bo��ݣ�@zź*������?9On�^:�1r��}׹!#���OC/$�mUј��t9���x� +��9�x�曤x�������rn�m�2n�}��W��ㄍ�����h�<�������H֒���3)�{O�tHv�o���9t:�74'�rd���Y���x���=�u+�dɎ���SǞ�$9��[�V��T՞��7s��.�U��9vQ1'�9ڸ�im�h�5�jT���ozRՌ�Z	���6���0�]nN����כ���T�1��ct�z������t��K�����sg-�<��i��j��n�B�.*ܲ����/6T��0/T'b�����W8�׊�޺�|�����Y���C<��o��k����g�i��Y�>��Uy�\C6�Y���
]Fޚ�ê#����܏��uEs�mԼR��E�V湠��~׎R_L�h�����9�h>�|��&[��%|n��#9�#����g��ι��Xm�H9�����348hDZ�wJ}G���YC�+J�R��eA���b�麙�����/j�Y���c"8g=��`�=�����HM��W7a���5Q��R�N-��7��"����羑
��)�;S��A�����&/]f�m���g�� S4 ��"��o��W]� ��aE�����Q���E(b�Ef�(4hL�T\�(̌R���$Aʢ9S*T�I,���"�: J$�"������U*�r2��PRdUkH���Y�TE.Y�Er��""���9Up���E¨��'hFi4 ���J�HUAp�e',.�QUD�TTE�NH������2
�hlU�2��R�'H�9r�p҄��g@�r

���u1iˡU��
��]38�bY�PUD
��#�,��GL9Tr�ʊ���*)3� fV�2Z�Tfd�G3SXQ\�D���qS�.DR@�*�������:�L��p�IPĨ�9�f�k@�.TQFE!DY�DjZk.\�S��DDRX�2��jf��5*5�UU�]�B%��)�&$N��UA�I$A� �HI"�%)1�&�c#QfD*9R9p�U$����{!�+�0FA��c2m_wn�EIJ��.V��G|�����bQr���������۬e�R���o�=���6�D��|Y'�P@�y!|�Ho��z���� �.�r6-�W��JA�����cI��|8.8�X�at>�r* ��6Ls+-�u�9��6�_<����h5􇙮�mӸ�����M��`�uHK�� �<>�v��!�ע��z���j�u����D��k��t��n��U�wT��N�!N6�r��X�t��x���4�Z���b/�`,E}=/���)��-vҒ�nc�0ɶK�Z��7�]\@����x�t̏x��U��:QW�\=�����p����Rb�N̙SA��N�����1�s��]��ҏb���
�1S��4dꧦ��Ϯ�A�'�yL�Տ�w�Oe5��j!�`�����Ԃ�B|�*�an��^y�)�%߉^�/���S��w[Z`�
&�:�"�8<����j ����"-J��9�h%�3sՋea�O��؉g$j�I��a����Vm�c ���7_4y��������0E�Ko�m��ڽQ:�&�U<�sGoLc�x򩸷����.~8����\0�r�+B�8qa�u3�Wf))���ۺu����l���d��j�o��Y�M����1<#�^�.(�ے�]�C~>���M�"��`:Q�����Ơ%Ԗ+V�T�������=�8:y2�|�9>���U�o9s�0��`d��Y9F-�����Ӛ��F��ar�����Az��x��T��_	���TtIRJ��ý3CG�`�t�S���YF&\s�5<6��:q1wD�O��i�p�PT�T�i��<)�-�C2��ؘ7���Wc�p�b��\�R��Sbk��g������;���Z���Q\෭���6>�_f�#b�g�'b��ܴ���0L��>W��0ŧ�C�N�zo蚝b��Z��O�Ť���JEv%�=�Z�g��K=��>7G�~��J����m��=�=Ȍ����'� �Vx��f�WLv��g,bPq�4ED3ʼUcx�+j��=������#��n��sH�by��1e��,��q{���aòE�u��)�#�g�WȅN�?�H�3#yS�l!�9����6��qA�$}���j!#�����:�ڇ�����]l ���[����ɑ�V{�b��4�g���b@:�	����a�j����F+z�=��UL�͗w�o�v+�ɠ��u}|�`��HpjT7�����i��bg��h�;�V�4o19K��4w1������4�7*�^O�}�,;��Cq�Lo��u𵘈�͇�qi�N[���Ҿ��	��-k���d�`ᳺ�6/M,];���ﾪ��p�+�`�f՜&����9��BsD�N�!i�G���u�3�2�U.{�-�c����"���cUrn"0���q&J�c%�
���G9q�JU��9�Z���U��C����m�pۤ�]�����,��b���$�y�&�=|��o&,B�*Xv2~d�B��x�\}�n�����{]T��D3|�͕�$�u=��ō�ᘰl�Ԅ�y�N��R��J����o�C-T1�5��9��3�,��991��{ƝdǢ
�j�^���;ӑR�.9�J�˙��k��:�����^~����7Rև��Z�+R�+�e+#c���I�]U�a�GOOv���(�p��;����䊇���m�b�.�1�����H˹D�$s
���n�U)���>>�㨧��&R��h�UP�:zr�a��=�LÕ/z��k�/�_���2��'����i��07j�]LC�44&�+|q�,�!���$S=X+-�&�4Pqe���<��Z9Zɏ��o3���\�T��V�z���;��Bl�/��wc��9~����E��
���u�n��^�r5�m�� 
��Wt�b�u�L��W��JU+k��Sg,H&n�	� ]8��ȴ�BF�:���������]7'����(��$��:y��2���mV�����QX���i�'��:7 �;�35X�S3K�`��E\5��bF�0֨�Na挆��F��}W1]o�{]�3S1?L��^�m4f�A����X����&����,���?�J:MZ�>f���HX�WG)][�w:�9N7n��T�:�!܅K�I;��9����+hꮓ��Cq����6h��ߥ���?��C%�<P�0�UR�<Q?(g�{�!�3ӥ&��G"�O�_V
���gh�oJ�i>����A�d�meڞ��7��n��;g ���]0svjO���+k��q:�ؼ�:�}yp�:�1����e�q�p��f�U�վ\��v+G�f�E)��F�IEa�o��j�5A�:͏~Q��&��Q����ad-N��<�T���s��;֕��.��{*�"�n�y����q�'����Ʒ	 {�C.m�n���L�+o�za���R�(l��<q��T������[鵾fz���x����c��,������=3ۢ��<�$:�)�	���+�|\�׽5^C�w��y��R���1�v�Vs�׺�5 �b�n-\���@e�C-ꡀKHp�{Q=y	j��xq��Z��l�����Vr#�G�|�o>���R���l��a�&�O$dR�l���Zٸ櫄s�W��
ߴ@=g�YUd�R��<�`�x��˨WM]ɸ������@+%�KG�z���+s�3nG/��\yޫ^2���$�����%�-K�1�\����:�F�`�C��7�r�],k�X�V5���̝Z�����+���� �0�
���ּr���T�.v���k��&��+ો�c��0��#�����a��,��X+3���H�ۨ��1}�n�4�k�$�!�����KF��N����R�W�(���*�r1J���Rs��Wkv[���_1Q��Ĺu9�S�U�88��*]y��$bu�*[1"�<{;�j�A����)�� O�Ʊq��r�NgD6s�s����V�Jl@�p��:Pu�"��hw������ �g�w�=+���ҙ��eD5��c�0ɴJP�3Bq��{H;��^l�=��H>44��w��<E^	Ք�b�[�ЏJ�P�f��!t�<Ï�u�T�$�C����+}\Ԟ�ڄ�T�HtɽĲ����n�*	���U�wF�)�����B3t�}.��d�{ec�t�N@��e�.Ggz퀵��U냲�`�Y��Ge�]%۱�(&D�z�Uys�V����K�}�m��9�<���71��1���<=�2~ڈي��]q�ꗆ��1���v�ռ:�j�҅���a��!��r�l}?d��x�>U:��?4��1|}�0��������i��[.#Ybڪ`V�<�o�*�r�}0ȊZ�ARs��z���/��ZܴR�㨲��ݜ�5S1�4v��͵l`!�n~h멃��^��L{]V�� g}�-e�d�.�,7�zr�]	�(�S=/��Œ�ų���f�:NV��>Ģz2:��cH��f8?f�b�L����:2*U���L�P��,g���D`>p>؁�>����w�WT����T��:`�e
kc̭>v :K�]� ]��ؙ��/;�ד�r��u���1Q��� F�����Ř�ثcC�φ�WS��J��GX6>�
��B����b��!�u���kG]G��	1��x3J������3zs��% ��qy��qE��.U�ֹ�����h�lG�
���R{�t��ίb�h�̽��]�JlZȻ(V���]	#W_5�C�޸�
��Ź�6����/b�D�z�:��2�kxЊw��.��aɻ����_͑+/�5z��k�$��v�����E3s9g0Y9��.Zq���;zy.{rS�7Cf�u�U_}���p�c2�@d��;0�h�ʵ43J�m\P,�s0�iϛ�#�-�#&��q���]����d���+�HK��<�y���%|(l�P���q���z;l�/e"�_Ym�T�ҫwe�:����>�FB$ȴ��cQ
��rb�}xmC��}�췎(�EE�]�yv�zr�7��Rݟ�L����E�(N��w�.�N�N�&l�1T&�ր��7�����w[]$$)�r��g��PҦK�e��>����u�L@X��;D9N(��Y;mvv���˧0����!�屉��7���健�ڱP���K'�Ƞ1��k�6��r�l#�~��r�)g����jI���N�r�>�c���1OI��8���{x��\+���t2~U�͆2⺗�7�3y���*a�c!��e\^˾�x���j��S�v`�U��%J�kRi��N��DT�He��K�\�z����*�4�w;S�ja2�ת��x/L�)�LV���C����tU@�{��=(��*��z�����HV[;9�L@D!�N�r���,+�i�gZ9���c�N�t��*;s1�fի3�Q�!G�}��+/�B���d�u1�:�vHh�\'i��DD7��椶J��s�4�+�<�%�V%7X��/f��N^Q;�ue���_W�U}��5�c��B��ꪽ�fF}M;�_�.�=����+��nT鸲�h��Ժ�jF�Պ�����E>�t���UC�1�"�O7=�_��K^|<;>X�]��˫P���*E�?e�ͷ�/��}Ec���P�Y���p�]r��a[{p���J��S�� �[O��[���Kf՚�a�(UD�C�=(C�44&�+|r���D1�6ՌQus[�5q��*�i�%�J��`$񠖒1g'en�n�V������,���i�p9�a��� �j4f���#%���sB�RQ���]�6�&�v���&辰���4q��y� E}~���}�x%�U�ĤWt��K��X	;�]�s�JG���
�r�x���K&�WO'pF
I�C"�D��1��Ѱ1Z���0�9��:��`wP$�o�.[
�q5��e�Go�����!Q�ʡ�Pۮ�U�� ���F�(��"���m������Gq/qFq@V�»�1 C��N��7�O����jS&M��q=���7��n���|'�YPW��`Ior�r�P�f�V�6�Lkd�86�@@�ؔ�w�En r������y��wC㗊̸��m9�t����4��j�yM9h�e��ï�@8����O��eM@�2���#z��Ղ�kұ���o��}U��	��6379�C�1d�َ=#
����V�>�Q���W�6���CN{���ަٗt�~�[�8l\}	�}^���U��U��@yP�S�*�C�p.���"_�e�!D���|�K�J�0j�Sk�##[��]|;&��w3g'3���EL̯!����χ�vt�k�1�N�^� V)�R�����b���9�}����� ة�_�h�S�y@#�k�����#?9�Q��fR%d	� �M<���$1�w��uΊ���1��_J�c�f��� K�f2,L�k_��v��4l��Z:������p�f��m�ל����΄��+�tXp�ܝWȓH�t�.����FE<�K��n`2������6�#�e��g����O�P�Oج��kE\ ���\B��,�_en���[�3������F�H=������d9���j��A��B�p�'��
��$/�� ��ʼ���p��ؚ��BCu,`k%�;����T��!-X��i�$.NDh_�Y���u
ۘ���s;i�t��K���9��v��
js�6�+�á
ơ��Q�tJ{�^�@�[��uw�������X;[Kr���������T"����]`TP�{a���⎝��P�n�;7nae��HO����>�����g7XQ>���/2��V'���p�s���s�I�g�����&"S�elŲ����r�+�4|h��]�ۡ}�^N/���'6S����&.��}�{:�jV;+V=����I�nKFɀl����\tn��L��xƺ����8C�(X�Bס;"�N)�ȷ�W��h�r~I*�U޺�k��p����Zo�ΈoŤ�ľ��T@�n��
s'�Í���l�cS`(�vd���?m��DN.��uK�{�\O3h��طu��`�{w���UL�2��!���m�B|�b���[��wW*�.iݷ�s��{Z�%^Y�<!s�޶4^����Sx�e(;ču2"�qu�Έ���\ro����f�Z,�w�V[FI����^m�cͷ_4y��͏�z*���x�������Y�^����ᾢ/���D�F,�o.��L�%��+�DJ�e�")��+�6����ƻ��t����W�x��]f�?���������Όj1����0��ۊ)�VS�V(����/y$g*!R7����Ym1]�<V����*X�����&33��-���_S=gt=�b�Kd)��"2�T�[k]�˕����-�fG��Pf��Bm��p�8N�1�^�S؃狅����缩�.{v��1R��D�m�F�LE8����Ա!�c�{�*�R�<7Ǔ\�������=l�n�ݫ|�p�j`Q�q
�x�U�j%���4�*ӷ~�8`u�ڄ�{:#����h�)p$�<�n��M�����c�Ue��ؗ'rw�s�*i��:��C�4���<t��f���z�o�����?l�s��y��ev/![�q;�PCa��$�����Z7�T������6�V��GU�)��T/D��/w��󇛋��#�8�k�a����Nn��^��t�Yy.jXmI�!g�*�ǔ��a#��l��I��%��o��N视��N�����J˽�!h���f��5�������s܉��I]�2��-}}���V�z����	�͡6���->��;��=Qu�/�Z�[(�ޭ�w*M��&�w�e�RH�Uكz�x�\�*��M��J�R�<��f���ғ�WWFi{�����sc��>KեG̴͜59���"���<9w%MƱ���C<q�x%3T��t�t�=��<\�3˨�sgK�3�/y:y�ʼD��y��]�8�e+}n�JV��,bW�S$��U��K��z@:E9�V��؂����sW`��#�D���vx�r^\N��5݁�u�%��%�:��M�ê;�A�r��5)�e�:k��*�ݨ������%��x��y>(�_k���9,�2��pC4d��e�����~����/��Z���Yski�2�� �H�w����K�B���d�b21�	�Fo���:܃C��;+j��t-'BѳOD\��Bw��j�D'���y�qm���]*7�6o�PSmV<��N�Γ*��[L6s��g:AK��bsbP�ܬ�Z�ޜ�������z ����NM��y8��]pQ5�b+_:ݸ�oR��(Mc R�V���e*n��.�G]�M�֩s;o���7�����Gn|�J��O�٫5�����>��I.kB�/%��P����,��x���\�ͮ�ٴ f�c� �)���I��7�O�h�C�H�F��[�F]s��w�g�& �Mn�z�MY}g��!�~�Z$���{���p�N)m�0W@9V_s��|^,oV�v�I��5����h���Ԯ������&��\��2T�I^Vַ����׷�,*,�.�����P���h�/j�DE�o�k��a��;B�WfjJ���J��:���� �]^J�y.�)M�OW!�˅���vnﰉ8 k�^��T���yi�
�Q԰]t��d������;�s��{��Mm�:�*w�fʜ�Y[X;�x�YB��.V�JTY"�I�bQFViK)L�+�Q�i��Q��Ѧ�gYL�B.PDA�ʬʤ�PQ�p�Q�p�Y��
(��	��%hQ���\��B�IM
*
�+8W-J��	8�*�EDUdiI�]���AQ"�шBg
�*ʪ���UΚv���Z�Z��9\*�B�d-
��EEE˳-�Y�&���jhb��-R*NQ���� L�Z�e�B�SC��!�$�]Ee�
ib\Ι!EG���*p��̺��	5)#��Qf(��p�HT.��*Y�P��Bs�J�"C(�Ve�9r$�fI(� �D�g"Ԫ�H�t���I)�PTr��"�hR��T��E\*�	R
ЫI$U�]��W9Y�P! A��9[fVU�5�'4����g��v&;l]f��:�y;#�IʄJ��>c&���,b4ރ GD��w�G��}��G�!4�S�}������⾚X�{`�u.�̨-���l��N��!�{$W���Qr[�ݛط	����__C���NS=���o�l.ʔn�0~L��z�5W�TA)�����eꞗl|�S����A�-��!��w��q5::���Ʊ j�e���쓝�/\��ú�V}��7^���xr��m����1��g�pY��w:��u�.�<�{�x�p� �j"J\�Za"�M��ڸ�Y�<�a���"5R��l�^��jb���晚�2����=R艔��Ce2��_��up�.�1%���9��SWH�{̃%;ޙ��(�?{Ύ��o��HȮ�_J�A�L-����V	�������n��O���rI?^^W��� [%s���U TGJ']��ta�H��)G~�P��]�]�j���X�S�
�|��.�?W�*d��fX����#�'tN	)8"�4k�ul$�ͺ�9�mf�1�[�j�N c�nXZɡ���8ݘoJ��Φ_����*�q��<��9/�g'I�R������-��_u3B�WX�:��9H�Q�9S���b{�Й��]̷YH]
�hɨ�$�E�q�Ť]��3����f�o]�	�=Y9g����ڦ���yV]�c�/\�x�n���(� t��}UU�U�7w�֫�\%���iA��_Nb��Wr��1���lG\$���jt�9��l����E��l�c�9���VL�b8�k�~�%��1U�����W��ʘxX�00�)u#���[��UjtN���g�j5	*TkRCO
TbJ����v��37|���O<��k�i<[�љ݌:c�8�6��Cuc{>�i�{�vA���T��ۛ�pN쮹��ǖ�Q�
�(G��3"Ru�R����4�B�ћs:h"_����*S���N{�B��e��T� �s�ܐ���s���bˮvD�}?v�H�)h���{����lT�5%��E[�lb[!aej�6�dn@�ON�ǵ	�P�SQ��(��&8p\6�����(2k��ixBs�q]HC�`3A�Bk���jK/��z���p�xϴ��j�u/����w %�J��`$�'I���i�O�ⵜv��e�;���r&�A0,ͥ�ވ�X�>�^UGT0��s>d*��?L]g˪��o)Z}��T�KP�ja���+��<zP#�`��y�.բ)�t�˸��ι5�re<��-����c�X(��g*���T0�S��*�.�F��O�آk#]A�T����U�C�r�ل�s�������0�-��������R�|�t�B.�P��M_��9�Ȇ븛�����~��=�:I���;z��S\���E�Jc�܀�1j�"��$ՠ˔L1+��������NlL�֤�v;]:����
R��WKG�!+���Lg)�Km��� �h���ui�ja��)�������@�*�Ǝ/Jۊ1"�W
E��S�����olj-JdɗC,��������O+�5���s'��!�*zD�N����㫩�_M}�.���%�!�wu�]�ˌ8J~d��T۬�ZV�zh!j�XU�:({��|M{U<٨t���0�.�R���`�
&�:�4T���i{~�so/���� J���*,��oU�-{P\��3l�Ǫ�,�����bsl�Cu��3"����6�_Ne��d�������7N�}��u���%<Lς� �Ob�x�>sU���\ΆS�i߯u�Fj2O0��#HY:/�%0������7�t�4o㮀@2��jy��n�ag��I���EB���7o����=�4^�����V�-�6��9�T�|�Cn��Ѥ�$�l�8���}q�C8-�&�V�S;�+r��L1�<c��܏��E&���K;I��J�:���]Ԩ��ܰ��e!A'�0^��z��0���}�}�}m�b��<�")?�y֋����qi�Q:&S�Nf.�QX�|�\�d�觃[��@Ö�
�ר�f�#t[�L�N������ӈ���
��k�^/�}�2dWs�[�yk�� _�ա���Ɓ�Y��;+��/G���\�´�s9���^VW!�?/X|�u�"}md�/��4�s��WS���\��_���}r3^�8(i*Wn1�C��m k<�O�b}q7�q���S��&ـ1�ꐗ۫G�$�H���Z���tV(}�D���[�eH���Ӈ�u}_$�#�9���;X9m=�2�KT�Εdt���f`؃=2K��#q�/SҸ���t�cx�����c�CD�c���JfC)Xu.��D���,~�Đp�Ҩ�]��:Ja���1q�+N�7���ث��o�%jօ�N�� 暓�vd�Bs��#��Y�O1���j��X2.���G
���I^|���Rʖ�ϻ�.wt!2�e4P��+�
%�Ʌ���u0�N�"Þ��f�jM����D���x�C�]]�<�װ�*$�����-ʚH�A���y�+V̪߫��z�d��u�2���b�ՙ��1�6����	�t��?l;�w�}��֊#�G���m��η�#'����菢#ﵷ���u�R������ÑJX��7�������Sblx���,/ƐU���EM�Ljc����2[�Jp
���P�-��cDh�����[���u�F��uf �4�/�*Çu8����ɂ.�|�%Y����ꬻӕ3�%�#b5l�\�&I���/Ճ���b��ӿ�����5���×IA��%�5��t#�R��=������}�S܎Mu%T!����N�(O��Y�*0�8hB�eAl�e
K��J�gc���\��B�q�U��]|<�����dS���1���nA�2�N�q������Ook
y�T��l|�+�
9����c-��ӿ���jtu��8��*�:����b\��������.6鲳U�n(�?T)T���If6����>�5����!F!lc�ˤ����ɏ�ɣ��U�N�MHe�v7�+j��=���1�@�G"ќ˼ټO8�/��̋�'� ���8��BR?�����eP�8���w'-�M��R���k�4r�:������_�]i������n�]jc/�<c'mҨ/"6-)�_MT: ��73���Æ��jR�@���G)ބ��D�h�ţ�xtSN�Z����.�LC^��I����C8p�c�\r^���Q;8�>����s�4�U�+�Ǡ�h㙌����^o�I�ik�Ƣ�rcM�Z|���/]��#�ߵ��{|����8?��e��F2U��)U WJ'hL�;�b�@*@�vi�fj��Ѩ).��1W�q��d1l��T�x̰9�W�
sD�N��g����j����n��3���B�gY]R�c�15W' 1�ܰ4��[V-`���k%#��nfr@���[_�� {c腑��s`ּ�{�|�R��Y�O��rOP\♀�)^սNʬ�����_����K,�6�����+t�c�T�O/��>�͛Ff_{���Eʌ;�I��"����ZP��
�7L&����b�.�yg�xx�K�jī-v<	��{���6�@;ͺ���ׅ\K�gq����[�*1�N�F ̯��!0!�C��v�j�!��-��+�2z@A�	�N�22�w�M�U?^�x�h���p�zr ߤ��1Y��\gy,��|��'�$xL�� >P9ݏ�7$T<�n{m��%�;>�����������/	&k^?#pr�>�����ε�b�V��69�]���>= n�������Q���"��b��]�ӹ��:��k�ab��u{yJ�5��9����z�������r�',�wj�I)�sD��5�ԣ/���G��L�Rroj�"(�'Pu�ꯪ��랧y�%��l��^��#ګ��yZ�(�Z��`�ON|4C-��fK͸���4��qi���+iq7Hu�d��	;S(	��u!\b��lЗʞ��p}x�-��\�s��a`�n==�4ϒ�[ �+x`D�a-$b�N����>ۈ�D+�M�N��G'.i�ǫ��=��������:ԝ+^�T�.��Ώ�	�HdhY �U����>�$e;+!�P�Q��z25\3�P��t��n�񿄳��0 {V.��-��jr�yԮ8��3��9]]F��0�Ů�pF
�&�\�j}�X<K�X�.�3��ίBSU�Ƈ��WS�X�1��K^�מ��b�|�F�r�d�6�lK h�5�T_�gJ�m^l��%��j���Ş_	��j��Y��S�����z���9�i1�tIH�)t����8�IUʡ��()��}����ο¯�m��Y�ȵ����hJ����
�~�k�
��P-m'J�'�crB��6k�oK�tQ���>���O7R�m�+�U�N>V��^��9�у���D��l��4���q���ʕ��*diF���@U�5Y)ܡѬ7;o���";���f�|��i���v	锖	���K���	(��!˴���w.�j���}}���6�v>��Dǳ�pv��-�}���p��~ѕb�}�pW�>�����so���vג��Ҍ�:�����A��`�u_�K�fq��b�9�Ӹ~�S"��'*)�-�ld��8J�aYg�}Q=�	)��� Zi܎�S�q���|�p�,b�U D�+��:f��E����ZS���\W;�7]1����%�̽a��ٮPܭG6���=��K�j���^�Gߑ&�Q<<�Z%����[�ȧ�O?���{��wuOw�§ ��ꨁ���缶����"��d,P#Z*�@\@,B;]r̾M��e˲b�i�yܣ��E�)�7L}��5��=��ۃMP����*/\����]�ݫK7��AJ/�G��=��%�4�<�kZ�|3��E-���g����X�&����_-pv�+᭬���#�_9}�[���EE�7PW�393 v��yqP�ȭ�����[#f:H`��P��0,���)&�����27s�g#��t�F)|m^��.�UN�b��w�~�O�X�w�e��"'h�]��~AT���uj�\��{y�3dx���%�S`��wKJZ����"Yv���\�����"�^�Į7��O����+�r���kȸ.O���_T}&�K������G���u"�]�R���'�n8�5n{k���穜�
5v���i� �㱰��a��R��Cg�y�m��yѭ��Ѹ����/yĔ��5�5��ZL�7��F�"~�6E���Z�F9Â��S���u��&�������潨]V�'SV�3P�Q�3�+"~�6�oY���֩o*�S��T��<��k��n�j^�'�t1ѣ�����Z�E���}�����=�&o�6��h��;S���pT�g֜lL�ju7"�&�T�J�\���я����]�}�w����*����=���Q?,i�s�NF�<O�������yzB���v��1їCz�o��#+�
/���w���m�&�Y�)>lީ��򾘽���hN�R�sye������#5��d��it����_ɧ�/����=�RN<�����+��Al��W�{��sǅ��9K��)D��^�7o�5Yv`���z��i��λkcp�ÃRrU��7q�Z�g�L���G�Q9��k���J7��i�7Ԗ��V��������ibRXz��u��E����%TP��:ю����������3�nxկ@7�=(����R�p9�����z�ɧ�kzFL�棶���g��lڳ��4I�!��I\b��zv!Jyp�kn!�z'*%p��1�1<��m�u
=��ax:�$��z�?ru������ٶ���5�%&�Fof8��u�/\�(��l�=b�����&����R��<��\a&��Χp�jLe������3�!u	J�h'�H�j�<pR�u�k�Ջ7���c�c�mk���gW ��_tC��ݥѻ��,�A�6���&�elo'O�t�Q���q�^'D\8��y�֘8̑M��z��D�!��[P��MQ�ឆ�k��c6�[K��]D8�:~��}S�t���?-���=��y�R�|���Ig����N�8���[�9�Z���m����|T���Ҟ��r��C��w�݂�w;��my��G�S�Q��"Q�g7{"�5tþ��O81ˠ]^��M�\�!�|�֓�6��ʦ���T�xia��ɱ�[Ѡkd}�oφ�Qa@���GJ��R}�����[�:��_vG��"��<�e}�H#�LwouDr[=��5!��k��*�ݛO�F�1m�#�]�cI����)�~z)#ǥŊ54ӏ�^�����F+���ccz��c�>�zĒMIl)\�vV����`2J<��
���b�`�]�1o�䀊C;D����er�Տv�uut�uc�sm�-!s��.d�f�o'w��aY�W[��#xpf*��;&�����<���Ɏu�y{P�3B�Xn�^X�s��8�FUb��@H!�sm9,�v���wOH�h쇖ֻ
�p�W ��n�D��N��'��ӛٍ����X�+su�&�i�Rʕ�9u���5�ڮ.�KE�v�u�<:^e[Pfoe���8��
;6]��L���+_Vk�:&�ۡ�L�g�����2���jݳJg=C>�QH�bc����3����$�z�3v�Q<l���Ӽ���ۋ١˞�#�>�>�{S����:T1�~%W�S�.��	�݇nL3��A�(�}�C���aЙ7�z�K���M�ǆ�!�������0�3���)���u��kaL�|�j��l�ݚ
��R���o5�p���ǻ�S��֍�i�s+�r�
[6�,<E���{��(	[��e��ۢ*���d\�T��VK��y���X��t3[�c|}&�c��I�b�S՜V��[��7/r�\�M�؎�bV��Ǒ�+8b[|�+nZvb���hur9������x�jys!�Y���}��b��/@��s�Č%m!�d�يF�DʽO���vqyxoǹ�_cA����{�UML%�u#��r��%��7�ɂ��{M��mV��y ,.�ǟ��ȃ�	[�E=����_0v���uX�3ge�j׼�Z�9�!�/Q�y?�6�K|�hۖQ��rvu��r�:��奭�)j��������gz~�}��hT8
x�O�o�ʹ�O���ï�q<�u��v�^:9I�T3xGI٩.U���!~p�r�w��tL�o�����6�)Jd2��,�ډe@��׵囦'/u����e#g@�je�>����3޷i��殫��,�S;���16�>�\����Ai����4Z�VE��-�u��
���J�hڑ[KK�pĲ�;�{4��u�wr��x�)�::z�3Jp�8��o���S!ފ�˨����9y���d�yײhͩ�B�1­�Lg�,�\k���N;i�kiE`sh#�Q'��%]�K��K#�d�ܺ�Dy��o�fp ��K���^%fǞ�^/L�����V�Tf�A��uw/A�lU�́uf�Uo8������6Ĝqt~��T���R�Je
��d$�Q�p����r&*QAL�.	�J�TL#��H��Uʢ�$���ԍ)I3"&�9ԥ��buȰ�fˑ�`RE�Yi"��CYT��W��-�r���L�DXYWJ�:R���,�ĮRr�IV��ؙp�B�&bq8f٭��VuD�乪Y'N�Z���e�AR�P�$���!`�l����,��z��I:Rʹ���Uʣ�r;p�TMY�TDP\��Q�a�҈���I�eP��"9W(�̙�0���!YU&*]�ܰ��P�J�&��*�
��M!5H�$�#R�.]2eș�Ȍ�B����b��4���Fu��(�1�Qj4*�N{�L��idQ����Z�_��_bQo�>!��+�[	��>�J�9��Y�!�	����q�(+�N��ε�����͘���諭��y��N>�F��"��/CT�����)��m)d螢a��>�W�Md�=t�z���D�9�8�i�\ظ�o[��Ҳ���d蝆jy�w}k)/5=5t)��:��%p1Ŧ��͋��)���r����o[����Ѻ�Ҳt�s}Cnb]_m:���	\t�6sx�����Ϻ��6�����ǌ���9u�z�5gg����yT첮+�*���kw�o�7e"z]qU������G�����[�#�#�P|���1Pe�;ԇXݞ��9l-]��)�����{W��om��ȟ7�Ԅ���#J�C�V��������Y}z����gT[c*�P(.��l'�*5OZ��՛���.���O�ܴ��[�����Ʋ�"BGK���Q��TI�UN�	�SS��p,U��RM+e�v�0��6�����vu#������vltXV����_�xK*�s�K�by�P���#����o��������<�5�Qv_x#����q߽}0���J�4�{X4�d{a�ϟm�:©#NT�9`�髪u-��uŭ%mY��Y
�2��*KJΐ�̵�������Y����x�;����D
�5<�j�:��Q˙��4�������T�U�7Rc5��;(��6`������Iŵ���oR]+��6�����sI%�J1�y{��뢯l�G�Go�Å���<�KވP9�[�����ᕌ�tz#����]��W�*�E�ί����kؕ�y��}��E�[�j^�'�f�Ys<��b�l�Z�[�����t,fe?��S6��ڢm�pT�g!�j�f��2֮ʤr8�Xڣ.o�7�2���΢{+nJaX�i�J�kA��G,��R��ל�n�M[v�/l�E0�*���:��Ӫ��`lnD�����s�{�M��q\���6�|�����5�v5�ŭ�=ͽw�!�L�y�ѥx���AV�s�5��}n��5��g�)�ED� u��W�a�3/P�������)�޴._�����	�pnm��V�`�K�l�������σq@��^z�z���["	��m;�Յ��i�͖m��jC�x�ĞJȸ�%��xX]Vx�ӵrN�X)T%��Τ�y�][Z����ݎ�s�_�}�UW�|�(��2�@��/JtW7��5�����OD���O0:�'�w�L9�iBA���^���x?+[E�KzQN�ֻ>|3��)C�P [͸���xsk;p��8K�ٓ`�OEi� -�����_s�;��EՁ�Y�X��.2Ewq��o�<g�SЦ_�	��M\/j�`자���Ǧ�|T�VnRq�u-#�)��N�@.��|4�MO.����"6Gt>`q��;Ła�//8��l��d�(���YV�������>J�sx�Cn��\�k�YO���0��;&&�]������O�����x��i�|�U�K2��oj�5j饩:���ᚆ�ޣ��9���P���Liv��;�|������<���{V�{q�����c��0>�z|�I#�pow�ٺ�2/�@�D���Jѷ��^�w�R�!����寘�;o.�u�u�do#Iu��lT���y����!;ނ�xftZ�Z`���&�����c�,Xqc\�K�� ��ӡ��&�V)���wփ�܊ǜ���6(v�=��Xd���'r8_�ǝif��kW��\�O�}U�UV#��{�qk=���^sF��̨.��TD��\���J��å<E�N�C��]^�������ovlŻ9Q�fW�\��}:�ml�(I��۬ǖ�q�
��7_al5ͅ��=y�+��/l��`�דI�MѦ�J]����.�h�����-WlW�Y&�\K���ڶE6y��"�n@J��%�܁��g���
�R�c�ǡ�x8M=�t�1'pɻ��hk.���9�@)��?�+��I^*�[�JSˆ�Z�m�p=)M���|
���g��C��}0Q�$�iIu����v�
)���C��(�_�=�t�׹���-��Q��
~ﻃR�QSYi�M���v���N�Sw������C;��cYg>D.��@вkL�K�ٕw��ou������>��|r��|�3�+yJ1?r�B�wC�pʋ��z�e����s����\�	�P�CoF�ۈx�P���䊞��L^�U���o��o���ѷf�E!#ѯ�[�)^�hp������V5�Ǐ�yԔ��u*'���/s5��\��ܐN��<��]�	�dnt~�>�菳�rT���mx��m����o�}	�i0��`���Wp�ݶ���)�*_��k>�T��y�^jڍOjOZp�Уx��5]�7h9�Ke�ɸ�p��VD���3�^EV(�񜷞vͽdf����cVL����ƺ7���b`Zꁘ��q���������{52_�;7����HnnD6V^.�m��]�gͦ�ք�gvu�{�K�Ė��=q1XӸ��lO���n�g!��N7[x�����Z�p+��VVܗF8�M2W6���Wf��� ��G�²	Ι;؝	r��X;���u�ө��	X�J�6*s{��B�4JH��=/���J�vc7�|��@�kW�\Dک���C/{y�1p"w�������'�����/����C�-�ב�d=eB�_����)�SG��͉���D���w#:衅��{A}$nb{�.B�+��rpO�\��I���<>�y@�h�i��t���1�����#s(��i��G(���xSÝ��:��w��If�ޘ��t�� ��j�!��K�RО�9����" ����AF�vy�kn��o��A���������t4dp�U�Ue�Jo\�{	X�ֻ�O���ı�_|�g[b��Q!\w����.Wi�⧹wѸ���P5�gb}��p�j�o�T[ci�<�d�o�g�[K���d&����U[�'�n)�s�V.8�I��?��-}�cU��c��Jv	hb�Ʋ�î3�t��_o����n{k�Zߜ~�g�X�kL]}��3�3�y2�U�!Mr;��?�&��lo-��r�*�=t�]7�a����i��ۍw*u��!��W�4so;J��.I�w5^eGE���r�}V�9ΌNX��w3��}�8������;V+>q��O�""7k������q��Y�vQ��f�\Л֌����[��aS����_L�ۉ+F�v���i�R����Y���B����A�z�����bA��3Eݩ������1�Bp�LneW[�7]6�������٢��1�]|)B��d�u�+O��9���Y�p!�g^�+����	E�朧��1V�6�+���W��xL(�<&�VKDd늱����_}�����T���Jn��}d�}�_�'vJa\@��d�h4�0��jri�Q��r��ê�B�+��gܸ�~77���D�S��p��畕[��yf�]4,\�"�j��f���ol�Rf9��S���=�X����λ�v����N�)�k/���I������H���s@��^��=��)N%N��vJTW7�C�X?�Ol�U�V|X��X'8���9t��s��n4��mR�Or��z3�e���g��݂����T9��꽵��򇾑_ �	���a�9}��>�÷ә2��^m����z��Ʈ��fa��)�����d�F0kc�6�G|�����jxwv���i���	���3(��R�	��M�<��MK�J�8}��|ߦ�;/���3;�a��R���6~:H����.=�m�O9�9���BT.(����x$�H//ޏ�Z�>^ J3GV���A���i@l��s���do��мE
�/�㝡)+6�m�4Q&�"��V�у���\�^��oZ�x&�絖����&�p�U}UU��z}��)3�K�zޮa���i0i7�A�DLr;>�a�n��ܧ]),��O�sWf\Nrڼյ���N��8f��7������i�۬��hCht���3}2�.|�y����j^�bp�v�d����o��2�7^X�+>�fU5ô�9W�o�d���>�V����g�y(q.���7'6�­g%v	kW�s���2;��G1�P]ǱSy{à3X.�s���{f	�{�.��Ļz�����ts"9�������z��dwv��v)w8����Ƶ͋�m�®͵}7�r��s���%���+Hǉ#�ׅ�XgkA��hr��
��i��/����oPnv:��䳵5���R:� � �0*��.����%*V9��z���{p���D���܇��p��b��T
1��*|���W�:�[�JS·W�Vj�� Um�eқ�j�mjx.�����,d�h�{����]�'t��)S�z/�Ɯ�w�OQ�k�]��ION�fZu͛�ʎ�T_Z���>Yon�r\���)���G:.�� R��f��ft���A��SL�R}��}�p�XZ�=6:��>j>��KE���=z���3SR{ŷ{�[l���춻��'����b�g63��le9FQ
c����)h ��S��b״�f��Y��_c��ZL^w8gp&�k�e��JX��8S�U��]�oPՈ ���Y�u��S\��������1�P�.*�k�o�����,h�y�6��I��Y���:O���i���)՘6��jT�3�^.f��tD�j0
��Յ�oQQ)���@}τ��e5����=���<���dO1��Vy��UV(��F۪`�j�r�]�$,4v��z��e\c����f���ڲf�gx���>���W��7��o�Y���ai�s�dF�����F��E4������7��з	��'Pۈ�q5�0�����n�osfݜ��L������;�����R��Ɛ:gB�����=�C;��2;�y�G���Z�sq��X7^t���`��o��6'0�o��Z}�å�$m�6:Ƀ��r���k��1%c���&�j��y�4����$��t��/.hς�������MFJ�x���DOemė_�LZi�����֫�vB�Nw-*���X��Y���]E\���6�I�	p�J1����N]�w(�WDw/T=�p��z>�rƸ���χ9�yWӲʞ!l-T�-�ш�Jwݨ�R&����S���}f��G_܀ق��|���ƣ:fm����\��GX6%��5	���Z�<��l�T(v?��J�͂�jd��0����������r�--k��Ϋle9J�}�yeet��2�ӿ�?��sX��kk2Ψ��n���չ�}���Z���D3=�s��Qhv��;�{����f�W=�b��M+e�uNU�Q�u.�b�3b�z���{r�q�����h%k����W�rt��S�/��Y��\�Q�Hs�q�\g�Q<��3���ڬ���nWz�w���ͫ5��`����_%&e��\�luݨ��j*4`�X��*��� ������[�	��k<��,~�w>U�Z���1�4�B!%;�a����(�E��q�{�6Q�t�%�A����/ ��kQ�6z'J|���sqo}{�f]=T�<g����}�y��hU����ݵG�JÚ�@��(LB��on�u2��w�ܺ��?d.���mW^�����4��Fˊ����w�\M9����J��%�w.�a�-ZM8����8i��
z�>� �Q�_UO���ҽ9 {<eh���N���q�j!;He�{�;���t�e �nlh2V��i	s#Yەw�p6P�%��\`'�f����'"����99G�xu>���mJ�4in��nv������yr7V�b]GiܵQ5Xw9cQ939�V-�/\�h	/9��y<�<���k��m:.؟n,�Q91m�����ɤ��cjgC6ʺ��p�f�Zs�1+UwmAMv�E
�8�u��ns	2űUwɊTM�ff������Ay1�Q�e��U�ҏ|�O�܃8cœ@�u��o�� 'D���8��}V�}�)2��:\K���*+�EZ�u����q�fulytJ��2�l��i�ٶ�&�#
���a[u+;�+g��ϸ��G~�w�Q�Y���_t���kI�ln�:�9��EƤ�C����xb�R��S����4t�M
�!��8�>�R뷾�M�Sʑ�WOyzy�ѕ�^z��0�y�gr��ZZE�9�3#6t�]C��Q����
a�����=;�������f�z+��{@�e<x�΃�.��Tkyv�:�xdV�sj�N��R}�n��)��í���d�1y|�
I��W��N<݌�s����$�c�Z�\×���W_EG��x�xU���pS��dr��H-��K̀��j+Ǘ���hw��;���i�}�5`R��\{1�!=��g�Ĭ�A�Zŧ�{d�4P6?�s��9l��-�(�_AٰQuV�HBQR��S�=����{F��y���s�u��ʬ;���.�@z����Y\��Gv���6����E�&1'η8���{�`��qԊ��ƤW���)�Ї��W�k��ZѸ��b��Ad� �]Jp��&��ˆkuf��S��A\�ϐ@qm�i�<���%�k�w�RY�vʃ��^]�L!Tt����,��o@� ��.�W��ޗ�]r4q�%J�6�����mӛ���D��`�QcE_;3���]���	Ip�c�ka�B���z�n�pc�H����)S�ZKSMK�Klv�����Ġ��B�̧5`��Zㇰ�|	~��q�F|k=ǍܶE��:�E�ig� ��Z��f�`}��j��?:��������U�@'�d���w���Hw0�L��MPpL��\��L-�\�i�����J=$��	�p_�8��H���ar�2�d�DL��$�9AA����r�3�(u�R�e$�R�$Y��PU�r���L�9���X��hҨ�5-��M1Yg)�VeZ�P�:qwK�:b�+b��g
�
�"��[Yr��N$�S.b�3�Ҋ��PsXP�P��D���Hp�A�R�,X��Ei�C�ӦF�L�i��c��\�+��DZgs8S���X]425N��BJ�I�®$Rl��rs�I�
.�2̊�3��2�БD�g��죝$�-@֪*N��Y]�8P�<��
f�%R�ww��dQDF�sI=�� �3�X���+�aYAF�����]��-Μ�k9�`Se4�\��<ء���wsȗ%�v	�If:8L��)rf�Ù�����۲��%��ﾣ�2F����o4�����6��&6�]���]�1�t����݇�qJ���=�}��JI��kڇ�j�:�N��F���b1Y��޼/TT��뤂YUZ�l��y���N����^Zx��������t�S;-�;{Ø1�[��#1Tͽ�+F�v���al���#e[�w����@����篬���3*
��OemĔ±�&�L�ۺӬ�Tk�4��^�a�V>��"o�����/�D쪰�^�k�KuO�F�3y�����1NαI�{��W�6��O׶r�)���:�8�Up���j]�/[[|OpW�y���<e��\:O���ݶzP{���{<�h�{�:QN��)I�\޾Zz��wƚz;�sؖ�$�ի<-�L��:\���oM)O.ֻ�SS��h�֍N��2�~�y�P��a��<^Y��wM�h�jWo|��B'u�t�v��bg$�s-�	֣���n����Y�:ek�>շ�G�T[N�k�nt�a�]R�X͎�L��+k�u�����M��=����:G
L��k|x�b�C{n!L��ªq�\l��H����NǨ���U��C��(>��Q�-���Y݋�xy�S��}9\�l�%���R����EE�6��3�!LGBP�AKE|5s�8/�t�o������I����z�gpT&�*30�]BR����@ET�[�^�V�/�7�|��z�ۛ��*�i���3�;��T�g�Cdx��Z
��-��(�K�������y��i��i0i7�dtFؘ�Ɇ�w�&��K���6��N <U��ݘq����[P��ZN��ӆjc\�:E�M3��ͭ9KR��]D=c� [ځ����̿��5�F�ڽ�m�t�gu�Q�gS�q�	�G5cj�����шd��C1TL�돤�qڝ>��{��1Z�p���r���֮9�ڏד�F�̨��G�T��#�{T�����|V��J�s���N��t����J���Y75/��W�`��T�ե�b�#��05��"�*{T�����4c�z���G�W^	cx�G��3O1Hz�v�C�pِe�|J�gl�	���ɯ��)}3�]`yЦ�\��Gj�tD��X%X��a)8;zk�#��O�(f�0ھ��_~��I��T�ϢuW_�z��F�5͋�m����]��s*��1`Cv��2+��;�~y�P�[���ˡ��x�M>�|�,��Nvm�4�t4��w.�������w�<��/b�¨��G7|�5�L\�[�B�wf]ݮ��p�����5x���x���(}~r�$�Hn[�1�%�=3W�1=jM)����yOE�)D����U&+�),"�qe@,�X3��t��4߫^�:��u�8�r���2��(�?w��XЩ��{SO��5�n�,א�#v�)i[9�g��
�����3���0Ω�k���*Wyj4ޗ���u��\�����l.y�b��P���ju��5�c�Èv:�rV����W��|�I�i0�rSxݾ�X��D�X1��E{�R�/>~��b*����������T����<��X�%�H���Wc�Q����V��r���G�ܕ�bWj�m�@�ا�`�"�w��4�.����8U�Q�v�0�bVmu^޾��c���J��&iW,�yM��F� r=Ԕ�2��'��5�$̩B�9v+*��{��y���}G�!`�.�%fH<\n�e��eLk�1��tF��=���Q�O(wX{p�OwRZ`�ڽ������U�;���p�/ձ;&."d�L�|ry�ع�lu�ju���T�y�s�f�Yy?s�u�f-u�9/if�_B�fS�[ꉛ���<��j��i��s`�y�7Y���(dl�#�PY��iy_0]������S�[q%CV1Ŧ���W6oE��W#��?؜m��W�_���W�ຠ���g�'.P5Ҹإ���WX�يB1"�;�M��uɫ�_>�{=�r��'��xLb�ꃟ�R�=�Q�@N���7��>�I��kz����P`>]\��MM+�|뷎��Z�Pu��|��>m������o�IP���|��jl,~H���ׇ;�	^�{�ä�]�|j�ı�_>�ضWVe����g䭆�1�g���>�=�6�'�lJ�[=�����#��;Ƴ4��X��&��������R�LvN裮*&(�NXp�u���e�)NF7��X�]�ؾ�R��� e���~���'\��/"I�.���'g)�8_�}���4g�1��`YՉ�ۖ���j܆�CO���n�5pT9F����o�<g�}B��n(��\0�9I�=��/c3=�59��F��c�8�%�0��(�	g�@��kk{�����������qû��Z"�no��q��d"���7*��վ��ș��y�[TVg8���E��q��P��MI贘4ۍv��]��-��N��\�]~]�)�*�{�|�5�ٮ�s��U��Fӹ�Vn��FN5�̫,�:羸eg�\6�7{V�{x�kZ�n��.l�n�&Q\ſ84���p�2���d�;�aZ6�D�XӲ��:�d�ʨ2�{b�eC��C��ҹ�Ӈ9}�N�8kVܔ±�$�f��}M'oF�3=e�),{a_zD���A5��tNϬ'����wӞ]�$#�qM�[���0�W�����oyyN�p�� c�N�u���ivO|1`��J���ك�X�$��vy�K��osn֏N\�#�ybJ���Z���v�l��]��XV�N�^Z<��>�..g�o����Vԕ�#	��:���#�V��m�Q�
����cZ��)����ӣ�]�^T�Hw��˥ˎ�:�7NN'�MD�br�kb�����-f�~k��%ӯxQ�#鉌{6]��0#��WXU�JTk�\��>e�k���	.`���yt��N+�����t$��]D���a�k��j����T�)�W�頭�ѕ��@��;��T	h��_|�b|O����I���m߆-��>���F�K�v����c�ڽ��p�{��.�ߴ/�EF�<�34�m%�9��;�7��:fQ��Uj�q��k˫�Oa���ƑRԙ��-܏�n�{�*�i���l>���&�Z=���k;�4���;^{7���}�s_D��崹�I�i0jq��C���%�a�	p�Pb����sF�\g��T[�{Ӥ��OW��=��v��y*��ޕ4�Zb	9��ɦ����;������Or2�-v���7���+ �7�d�kS˴rv���W��wknp�oS�9�|�Z�1���)@�ҍ+A���������S{w,XI�/��4m��=�������e�k��f�v4��y8�z����^����N���fu}2�.'�5����i�y�F5�	�ל�J�%k����v5Ѹ�f�A�}��fF����f�T�4�T�v��u>�%��s���8޵�Fz���#u�1�E܏b�;�d�P�gn͈ͧ��{�K��l8�
�8esb����n�tE�9_s���u�H��wcШ' �TD����.��V�5͂�ޅ]�p��RM�+r��ɾ���#N�wW�:�vY��	^�J�6)�kOce�(Q�W�`����Jپ�ݳ�H�P�ʰ���=����"��J�
R���s�fA�Z�S���]7��i�A����FQ���V�'dc����^uM�__v����{��0���Cڋ|2�������?	<9Ѻ��t�:�0��w��n1ֻ�S�/��gnCc:�-��Q�B�������ǧ�<zv;,P�[�/u
�z5�b���T�a�� �݊���o@n�9ۏ1����t\z���W(!��*(��"�44�����Q���q˅S�.d]�4��V�o^�)q҄6�kX)V�Zz ˖��s��6{_�R��{�zW�G�����+@:�h$�[ҡ�\�}B%{Pk2Ψ�]�p��l��X�M���,�Uu�C��5wr�^�
Pw��<��	��|r��j�|��-����1u���������LN���<�m�Z��m_���>A����ː��c� �	���؎��9����?'DO!�����D��u�Q-L��Ǳ$�=�!�=}�%ŷ���Q쉈�:E�����u��[f&�=��q���k9g�����m�pʿ��ڇs��b���*s˼J�_g�l��/:���2#����N��������Z�t:��Ɉ�f�F�t2�p�񵫇yy�3Ǻ��zeY/fn���v��i�S͌�����3k�B�V���z2sB�\;��	������'���p�����\�G�C���G�އU���⺧.ZK�te�v?�_�-�%������Ju7��Lq?��z5ӷ�b@���|=i^�}O��I�����-����E�׬N�_���*{�<�J{Yo����*�mJ�qZB��՘8gRr0K��1��(��J=A,��ZV;Υ(����/;���3��TqWf��NH��/6�4ϫ}=:������r�{ʁ�ꖯ��je���k���]�;AB\>�q��C��\C���t�	֪��9v�|ѥ�ԟ��O8�5.d�L�YN�-����m�C�|��%B�[��'|Z��pc�JW}����+�j�-�[Z�[���Ե��|3��{q}���#��bz��?���E{{�f|ub}��p�j�HU���wW�nq�����hm}Ҍ��]�YA<�k�Q��o�0|ۇ�C�I�x��ao����g�k"aR3�]�h�+\��kq�^�%o���ߋo�X=�rw�	�4���q��AR���6`�u���N&�JPcVR����wF�._=����=v��Q��q��eLF�"b9�������5I��jp6����N�uq�����N��8e^9N�b�zjv�do!\M݅�\W���c%�;�@؜��1�X���}��:���=�����9�߬O�t��m=k��p\�P����x�֒��m@�7j�DV��g����������	�����-ĳ�N�1WjWan�I�։Js9�_L(�l��+���sH�~��t���1��̸��ï5:��w�R��8ֲ���ڡB\��+/\+����n��w��Y3s;˰Ek�jVV�O_���֗��U���2���r21��J�VU�ͺ�3v=���{h�^z52�l7Y㼷O�قa�^�%�aD�Z���eg.%������uy��~�M�U������Tal5��ڸuٷ���c�n����}^��\לǈ�3=T�Q:�=��p5�P�5����I��kKn��X����on#t�Gg��A�}���u�Q)Q����կ�������!+���Eb��������;��)+�m_KziJy�s�nC�%�*�t�&4^�c��uE��[���P��П��y�q�&���i��N:����!��m�e���SC�ѓG��(��s�q7�9z�ޡ�v����x�`��t��.��<mgfj��.�s�9*2քl�_�sYٞ��gd��b��no���;k�v%;�A�p�CE_<��@򮈝���hӳ�q�Zr
t�o���M������<%-,Fhܳ݇*�בȞue�s��%���l
�u2r�ˑA�4��EXYqf�؇O�Q�CtV��0V�3���yAؑ,� ��૮�u���hq�V��
�t��Y2�. ˚�����VQ��+��.�rY����B�Փ��bӼ{}�Fqj㲹��ʪ�A5��bX���"����Ƴ�J��R����.��ΧR��h(����:66�E5�0V���3����Q�n�������作��5m;�:��^]�8�t,~)>�ԥ����I�0���uNJ��4�M�}���&搦�mӴ0|�x�SfsbУ̳�SU{��T�e1�j�}�ė��/ؚ�*�-��Y�/�2���6��!��}��>uK��׈*�VDy�����d��WYkf�73+��׊��6f�S�%�&tu��d��AH'T5ݼ����y�^��]1���Es��C8pe;,I	��غ�n>�u��������W��[ק#ߠ�;�G�r�Bs��ȿ�aL� ��ݥ"�wk�|cݏ\�+�p'��t]%W�pW2�^�y�8��	=1R��6�P٣UL�j�*ʸm[AX�n��[*,x��p��ܦSޕ�Y��C�"Н&"�g%�+���Z����)�JG��4�Ո��R���1f_ru�jk�s]���9A ܚ����C>.�?Ob���9�}=�+�r��O
N��	#fZ"�.Əu�V�S�IKk�I���=���B�H�_3�X�ĮPA��v��$O��(.@e���+r:�ϲi4�`����(�-����<լy���6��T���9����f�Y�Nm�����W�	�;��N|e�!��c��wD��G�.��权.,۫�ge�w�(�Ӥ��N�X��.��x}dLK4��΅.��j��sg7��c��Lj�S'@�>��WL�ѧl.Z��N@�zz����:$�7��Oe�Nټ�a�<����X5K��ۻ���#��:�tO:	�Pd3����PVe�0Z�&AB�����-iʓL�i��n�A}��a�9���u�HAsn
c$���X��������Mm8ȉު䖽=/q���&���9�����4�T�ݨ�wa�e�*mgJ��ˇ��W^Ӷ5�]r��z&Fb����H���v�Im#|#���.T1峨�0V�Z�r�J�u"T9�8���u�	����6�]ƥ�Y�&�`&�K�R�_�(��̋����q:	.���0L�:�s)�͝]e�9f���E�nJ�/N�ُF+A�cj��"Cݲv�w#�o�����|uO�����ϯ��]�X�d\�����F�R�\,��	2�?�ٻ�ˎV&QB��V�)3V�������re'��8ED����E�㎴�k���N�*ҡ	%���;��2̈�(MօCs�,Zy����V��Eg4T.Y�E&�O#B�72H����Y�Hu���"��+Y(Z ,Ъ�Y֭8R���&��V9;���Qg
�S�At���u���d;��Uf��P�j۝�Ls���t���s��!��8FIӚJ�5,�nI®GZ�����	3�u�-3��-J�,B&�rD(s�9
 n�Hb��9�
vG�" �p� ���((Ig((#�N{��"�hE�ww3��2��:j��K�U^l�Ωm�����(Q��g*I.EQ&�E��5ι����S=���s�L�L���$��|	'��S17"N��[�Sw�7.+}A_t�b��i�I������A���S���͌Ѝ�W�;x'6���3_��K�ދ��)�S3�X��I�l淐��M�WΙ@Fj�C���^�ü�8�_�.��8� rt��S\�Co��gv��Q=��Ǘ}X7�s^Bj��{����ͬ��W���0��4�`��h�veӭ�����\?��5ȁkh;��$�-�ڏzt����^gi���T'�)�Ɔ��=���to�VD�bE���X<k~����;������N�	���[=���*��ck�s1��b0/��fG�W���W
Ќ���O>�æ�2�<�����g�oZ��C}Y��F���=Ϳ1�^R��������]�ɯ�)o�8Xӎ+�.��kz�f-��,��J����/���4����X�~��ۉ.��8X�6oT��a�
�Pt�j�
u��Yڈ�QW0���k��	\F�J�6)�k9o��塽}�ps�1w1�:��q�#A��WNs�a,�X}|��ױ�{��8QJ1/�u�!��&�{2{���bnaM��`Ç�◜�]&ӕ!t�+��M�];'-���	��e��`[�swH¥hG.��&,�o7��.�S�a�R�'UHv�g�,��z.���������z5������R9�Q�Yʘ�����fR�7���C�M=��oTU�.١>��d���J���6A)��8Z�N�5[ƃX�,qo�R�����}0T'|ZR-}�7�ҥ���j ��x�9K�9}�����uE�1�C �F�f��gv���I��g.���&x�����YՋ�mKJ��sRc,oɱ�&�j�i�Yhw�U�	j�.����a6���)�j���Ξ�A�bg'��l�sy#_� ��l�Πm��jmv��'O�sU�󀨽�GusENa�C�2�]��BtD�r�"��e�ﰿ-���5��+���K���k�/s��Ri8��q��V�"��_��e�VՉ�$6^.~�k�ԦS���[�^��Ns�8ec���g�Vn�1�d�}s`X�k�;4ș@fN�F�!������,��������6���k�4�Ntj��;\\����w:}�S��)�����vs�e>]Z����}�ݶ���T`u:c0L��c�]�R�ih��ib��*jӕ���t�MMZf\��JSO����S5*-s������N�S���nu��^�{G�M�l�1��kQ���9��zY5�ތǑ3u�'���Q?V4���}/S������If�Ӻ��gd����s��W?��N�\qi�j2�VW�!��T���f�c�}5��N\���3.����ʐ�o(�֗�<c��Ջl�*��a�7�覚/������:��5���w��IЭ�it�Y�鱗�])��V5�z��>��'���܀��`G*�s2��s��Z尡��ڕ:�}�:��������y�o��rv�&��r{��a�~��S�jJ�mc-�e�ֹ��W��Yu9ъ4�n�Z=�!8ﻃRѵi�p�3�xzL�i_�g_c|D2R��-��-������BSA��sj�G�j����<��L���)"�N"m!�� ����Cr�Ƀ�C@7@��CLٙ�/����.]F����tTVT-#+o,;7�aK�Z.�����@�Ym���9�m��FJֽ�zbө��ɌG��cvX��~�����\t���v�m��b�Z"̮'\����[o+&[E�d 7Ԋ�����g����T��Qu �.
�6_]J�N%����;�sk�Yڧ�o�L��p�Х?r ���r���a&id�o+w��й�MQ��I�M�֮s�vA�[Њ��4���k�<T:�N���Δf��}V�#���N����GD�������E��|�.�Q��H��1TL�˞\:�S��zԽ�$�������'�(:b�4����Ύ��ټB�><�f*�f��IZ6�;W�Å~��`z�'
��WA����,�����u"���9��"uyÌ�^_��=GL��a��7��-�N&4����˷��޿�6b��U �Ҙ��f�u��erJ�B�N�5���`l5�c�ڷ]�;��8�S�&,��qO8�ZYݘ3��pF'J�kb����C����{рn��Xn�e�̶�}j�**̤��v�3y����2b���������n^b�d�7��F�ɯ��B��K��U�1��o���
��h[�Ja���c��,����Ej��vvt��8�+`��@�]��$ť�W�a/�+Q��.�ق�3-Ⱥ����uN���4'*��.�*�J����k5<�l�ݕ�s-n9�m�j��d���DiIZ�.�[�E=���a��=�)0l��*/W����v`�^�y��"������?<�`��{<�s,�N�Sw��r���}�����NQ�.?�5~�Ҍ�=��V^��O܊������,י�Wظ�BM+g5�2Ʀ�=����`v�`�@����ҕ��Njy��rj�ʆ�������z��.�9/��9b��%ñ� ��sk��]�q���0����4�1.Uq6i^G\UE��{Y4�ɍ��ê��7E^ޡ=Xg������'m�ݫk�cb]����7\3M��qQ�9�kjgT�̸�\�)ǆz[͵?e�!>x�u5�K��w�'/o�U㱵�r��v�e��~�g5�}�Hy�*w<����a}��7���÷��a���Z���i(z����t��{%��?%Zo^�L�T��ۼ��c���ʴ�LR�(�x�����	�뿵i�+x�%��pT�ۭ_���CSp���o��YZ�����䲳�*�fۓ˶)w9-��Z��v�oZ�t6�=y1�F�̫�G޵t�_�����u�2���3u�'���acN�+���{p�޿�6D��;u�13o�.oM7�2���u�S�(|�c�X[saKo�6qo�N:�i)��]�3j������v�����ʒ�O������uӶ�uD�%AK�a]?���/�ٽ��l� �g����q��!��oz�������o��AV���5��=�M=�5�B�O܀�+���v���E�=i�/��%k�A�{N��m�j-�ʅ�m�����x434����(�e���sV�7��r�����63�-���jb��k���V�{���fI��֧�71��g��
��#{x�������܇=������!�|%*��s鸞\�n���k�I�*rD:<i��x�K���d6�%Zy�4��o�O�:�G�?5���&h�㺓Mw���[U�Q�鸠�,Y����N������W�.�Cs}]�嗜���ܵ�:+Ly+ �SfF>�C�vu�F�	�y6�ԟ�bE�JÃ8Z	��Q��Cdul-s�k��y5�fs2E�K{��H�ٴi4�a�>�d��6ۀ�J��;�h�R�1;W~[0y3����3\z7�r�7��k��V�#��kU�*��[Y]�/)�*�{k�y�i?.Y�I�]�x�m;��5Y����7�hE�|�I��Nn�c��Yq<�u���E�'//䞵���*��q�9v��hVc�vn�ʃ�Fb&�2O1��+}O6;3�.{?sǗ�N�u�l]�Y��H���6���㛌������x��i:�.I�W��c�9�~�=�>��ꜳ�\q�=�;�vj�^U=ɒn��,���ٲ��p*%F�N6sx�����s�K>:��V�^�Zq���/���l�o�S�:jZ
��Q���շ���O��*��Y��7+	�o���q�e+��տm_���^�&�hp��O�^؞�OST�gr8��%����bf��:{�����C({�7�vF��վI��4oif��F�h�l�'��7y6EλkM�c��j6s�E�rYl췖�oW!6�"�t6��g&jQG ^����Ζ���%�Om�k^��o���Ǯ:���]s�)�	}�ݬ�wr[X�[���Ե�s<�lX�Wܹ�ecW��׫���j�=�t�`%�����7�3�`�0չ+���;I�5`9M�׹��lf�fQ
ch?A�~��>���Y��K�����t�m%����R�G]���;�D3��>��cR��m_�ۧ�er�j>m�vˍw��E\�����k1߰�ya9���}o�y�ڬ����\��&��L�����S�!z"�vwri��o��b�j�S��q:���f���j���n18g(�T�T��H)�I��=G�s?j�u� �Zꁘ�ye�k�����k�����Q�ы��|3"�7)z��ޞ�~��FY;�~�&mf?��#ݽ�L���.|�~��3��Ki���iVf�]ͣ�PH���Xk��Q%i:&���H�t�xV�EֽwnX�+�G�5ó�R�8�^�MQM�k5n|�z���ǩ��fȎ�S�<�RXg�T�Q��O�5z����[y/	�3r��gB�H�Ƞa�f�.^2�>Q�6�smѫ�3(������L9�h�݊]�Ka�@�f�%s`�y����ݽ�����d�)�[��n��]R��DN�j��F�\�*m�uٮ�t�V��J��νfʑ�z���o��c��Ƣu@X�������o���w�MX�Qm��V�|�Ʈ+V?�)�v�U06`���A�=}sk$ѵ���=ݏj�AD�+���c��>i4��?�v.J5�>$�3���o�[/]����������,X�ݤ�މ���>��2�����*#m�0�Qs��<���0[��k�(��زyu�ar�g�z��o_���z�i��;�����=�#��L�9�YPr�~cc�n1nwU�v0�G�%�p7���7C�F�Z5m��1�^�q��n�|�x��LGA�O�T�{�M�=�ND���D|�	NV�_,{ܨ����L_��g�=3�'�8�}��؟�
5}�N���^�rGkk)���{W�oc��;5�i��5��9�<Q��ƫ�AJ�J�@%��ߦU\^^"R/ih�k����R��A�Sn��q͕�ZF����H1*�y+1+SB��e�9L*�l�)�ov�n���f��㚚�RC�L4��2Dk�p=�U2k���0�bV�}^�u���T�5�#�?+��Ҧ����O�F+�\Ʃ�=�fS(^�\h��]H(�{`d��=s��=��z�z��^q���q9���w<�,2w�=�UѸ�z��߽���po�����/�G�H򻁳���S·���p�w]�v��&q�E��u��dG�W��k��s��=qˡ]��9���~9(zf�l������;;�{��7�N����W�K��w�s^��;�Ox���=�&��?��>�n�<�tc�t^~태��ś�φPs�L�QѱR��9e�������0eͳ��y�r��
��S����������ߖT��A�����w�2\��mxi��~k��v��l�xMf�w֫D��{�u�x�ul��v�W%��Lu(	�qx��o�΀o8��C�����/&�=;،��7��q�A�����'+�B�F�,�O�/Ƣ��<eI�{�R�޵�}ގ�m���}w�^Ӟ�>/s�d{��:�웮
�%"�*vKGӞc����2�Q��V0S��||)�Y�	c���Ы}g�ڦ�s��d[:j��uM�%�~�� ��);=�3p�Ҙ1�ת��}���GA�bgqs�Jg燣T÷@��%�Q�`厇��(�D�d���w��0S��QW7�����ǩ�,��nO1#�+�O]s����n� ��@��tpeu���������鸇6�1P��Sڷ��d��~���.תGC.�2Sn�f���,��n�aj��H�9."v�\�V�_H��YśpA��a[�u�� ��;M���o�ú@��w�F��|r���{�ח�hz����T��m�~�D��{�������;�Y�h���:�cc!}��\�x �w���5%tP��znGcѪ�	E�l�_�iv�<2� ��q�q"�"��f̄H��*�'0�n����C�7U��g)��|a����$�z;���;&�7cR�9��vr%-��K|�a}9��2��4c�0L����&��bVYS�vXxLү���(���ͽWq;�&"���� �N��ؖ�ã �5ؕM�p����z�Fv�W)IP�lu�1f���}��Æv�Z�����m�"������ιV]>�tv�ΔJ�%d|`��@z�-Y�򰥦iݎ�#h%���{���+��$&V7ji��
�i�)k̙V�CI�ո6��c�,��� ����}-cr��7;���#1����=f���]�F-�4����
�����6�q�y�)9�c��d��/�7{���M8Ϊ��Y����no�$Im�Ȕ�'0cA�@�<��P^QB3��jO��<�8�V���,hX��фu�z�	46H�7uo��{��T����X^]�^��t�=��1�Ҁɔ@�4*+�ya���Z2�e��W\�5K.�(�Ğ�:�|V>$�(���]�*9�<1���bA+j��'n��޵a�����ճ�+��p�f#hn�r*�H�<�oʅ^��{Y�.Q�ö���28w_o�5�Bcv�t��ڻ~B���on�X��gx��f�F�ޘN�Gi���>��Lc9*�?X�~UU�Mg8 -�.�XS<st��_M�e����&D�pf,�gt��~��Fz����bN6P��ەt쭠k6��qT� �r hX��q-���'�!��lR�^�d��1���|S��c���>h���ʘ0�\>��f�ٗ ���Q*6�}�]�9��2�f�a���T���]��le��븆3��M)�n�ͧ)�q&ݝ��oU\���SD�xsl��UK�*�R�s�v�,1ۻ�Dc�G����(�Q�`tv`{ʏP�]'�U�C�����k��j�e�3�5j�f�\��E����M�q�6��33��R<�s��f���G�d�\�l�����;�C�]v6�J�%�q +�>�P�C:!I>u�$��/"����X�5��Y�甖ZZ!�g�3Z�D�s�
]�dȋV�+Ejg����H�t���X��^�r�F\����3X���	Y�I�nE(�u�yT��J��"ҵOW4ҸQZGN	�P�(y��TC�2�$�"�̂�Q�trf���J�gKT�wG3���¨��W<��T�ۮ쪹�R�i	�d�p��(U�������ڢ�Ĩ(��%
�M�SJ"�Fh�'<�%eD��[EDs�Ț�I�B�%�"(�
�J�:����B#�ܪ��Љ�c�3h�t�1̜�QE�d��0�Λ2sܒ4M4�9�1dJY\ԣՑ���+�Zv{�)�;�^*ki�˔]/DĬ�����Ѧ���F���5�$���v���>'��*2bC��('��\�q��o�Ŗn����/�Yq��5��R��\�B*җa5�
0����n�>k���d��!P���s?W��� �y��W��n��NDy��|s�t��*#:�.��lW�(�a��F_:��h��&�9FUG�}��07��q�}��k��]zP����c=;�\}�p��z��������OoI���VxyI��L�5�U}DLIo��<���3�-j��:�<s��?m�L�S�E,S�W���[�'����N�X%��
�n��1?J�*2�G�|���h��rֶ2&+׀�/rXn�;����d�����#�@�t�O:	���Gܿ2�����Kw��ꭿn�.�=
��9
B��Uɿ��xdx׀�Z�]�(�xo�e���v�O��K�m���oG/>>�����^�׺������?P��z@�'�b��ċ��	W��K�Xi���b�9�U��:p+��><2���;�}��.D7�1���/7�pz�ՔB��>�|�}=�e{O�3��J��AF�fo����JϷ��\g[���u��Ȇ�]��~����TZ��O���\�p;�Y�\͞�΃0�P't�Ue^��U�{[ U���V6��3��M�Fj�F��NU�o_u`��<GO�9�4p(saJ=Z�v��XdNĳ/%$���1�o,Q�*5KD��_f���[r�.컷�wyЊ�� 
�]v#�9-�1J��69��P�5{<�d�:�lY��n�9m�V�T�H�=��)���~���[^��x�-�W�ԍ\�܀��Pʡ�-��R�44�u�fg�O����ك� z�FW�{�r�^G>�j�e����W2�/�K]J<��".��P����"���E9p=ㇽw7��W�W���P�S�Z��u¾�Ӓt]�$�qL�Y&ϭUb�������DR�s1Wz����V@�W�������_��[��ό�s�2Ovm�n��'���t��8Z$�,	�|���xo��{�b|�xh_yS����z�U���g�fx�g�Eg�ﾃ6�(�Q�P@򯌰&K� qm���֏e{ք��W�����>������_53ZӾ�ޣ�_��\>�0�\�P��Ku���^/v��kn,JU��?w��Z�_$�{�w�zv���z��n3ޢ:��z�Y%�|��ċ�W�����HS��;�8�=^]��=���Lc>��#Q�߭���@���;^��@�6���e��\�ʹ`�Lܫ6��ax�DMu`���&z�G)~7LTm�j�&���ȟH�8��9�=�O������x��=G�z����J�;eXT���[W.��快����v�u<k_�rߏ?':�8���ٚ����sZ�y3tH�W�v=�m��l(ޅ]��=��D��!x�d�ג;����T�:�U�:�����?�L�?���>4�^b���T��5��?;�1q��̟x��R�AW3��ŉ�{h���k�(�Q&X�ab�u�r�m�W�_��2��FuY+۞�cfkgs���=��}�,�ؑ���O��_�'tú�^�ϩ:@�޶<,����wZ�ݻ}V�a�����K�Do�C�/{�`�{�Az�E�d�t��7f�e����jԩ�w��z'��Gڽ@T^�߁s>�L����}1g(e��KS���It����7�$��;�^+����Ez���2�,��g�)��NE�d�9��g�n�*�9����ٺS��3���YY���&xe	��]^�����9�=>�O��ߝ/q�����\oh�u�Rv�U]���Su�=yS��Ԑz���g��^�q\�7��U���!}��6_��1~^��~�љ��5�^��gUmGw���]�(�Yd��,�S�J}9���n�H��,�vǲftѿ]]�Gyr9jA�!�p���#�p�l{�M�����#�J ��Ot�eߍ�3s5�'/}>�1o^��z.ћ��-�ZBP�A��+���	^ ]/j卺5{91B�A��ɴգg{���;�̜$��nv����3m|�_8��Ji-�������Od�q�&����cG4�μ���m<ɜ}}��v^T`��X�{��B�m���wz�o�����>�2�ʈ�o<���uL;˚D�$11�gwz��j�e棛��
����Tr7���o��H���ZT{ʸ�3޲:�4�ә��s��O.n��+��l�W�i ���:R>�ΣzѨ��M�~����Ǧ{I���_r�mq��=;�����FG�2S�&<�Q>�#BⓥǶ�=~�dmǚ�I��{�Ϗ�.\W������V�-��m��F��s2m�&az�J�����X�q�Rƾ�ǌ/G�S���]䃜�
�w:�����'q�{�RB�OPɇ�z�2Z�ӕ��z��y	�C�Lg�Y��{��i��=�u���?U�����S ��dШ�yR�O����ݨQuNZ0�z�ʱԫ�k_D�m�S�ϙ�}��^_�G�W��P�9�ʃ����w�ɼ�e���ܟl���9��s5��g��Y~G>��q<W����wϥ�{O���|S��=�oM�~I����#n���=�(uM}Z�/��իK�<��1R��=���[,
��yׯ��z�ǽB��������G�u"�c�3��{}(��ٲ�z�NiѬ=j�'���.��?`�.-H���Q��� �MV��sK5B"�$�7�1wH9,��'1׽�#IjP����U C�*Ij�b��96�Q�]������enT��*�OGr�X˻s�����?~{�Ӭ�֛��c* ��z��EK�<� mxq}~W�������x�=�wS�g�3އt��Ǌ�����qe��fa�=L]uW��W:�nN�%�t&��mג�x�	�F{���EǴO�܇�c�>�Znxj�F���<j$�2��jb��f���%�le�I�WPY���w"�{N{���Ͻ�G��9����pV��`�9���P�9[�g:��e��[�G[�^,f���>�TO:w�9�'��Ͻ�|{<���4���ٙ�4��h�����<���AmA����7�l��k��qߩ
�W�#��Z����m+��#"l�=���*��A�z���� ����K}$_ǝy��t+�Z�8dC�;bk���(�R�Fnw��bk���=�߽���^��	eD�n�
W�Q�Z>�ׇ����߽��<��8I���w���D���:<\�`�:w�'���G\�D��Q��r���2�s׏\�-�~�v��9y1^����y��>�� ;��	�~��\^'���^�r����b�x���z���ک��v�Ʈa��X/C*���;�N���=Hf1�S��O*.ý?NoC/L�{kK����~c�����>����Q�^�W���$qv)���SBhn�ۧ�iCCv#����e.��Z��vN[2��D��q@���)�>��x�����k�q�~wrq�@���z��<�}�'f/��da�hg���ӏ�B8;�g����xdWy_���>�Fu��ϛ����IO��\ʍ����ZᏻX�K���'�sه�/Ὸ��_�����*�<te'H��,y�u���^܋�7ڼ��y��Ա��͝untN{��{�`����3eqd��'t�qU�zs�^�S zWˠd���nu�ݵS:�z'i�`�z��d}�U��Yo}-ڽ\���1ԡ}�9��b��؎ׂLU{(3Z/+,v�8�0+=x����T�{�g���+�j�vD<��t䝢��=%�u99�9�f�{kT�.�~��Ew���9p9���8�O�Q���T?�=j�M�
]9'F]@Jz~��0�����k�L������S1u΋/��k�ޯi�t�i��K�Y�q�|���e��]�k�@64ܐz�3�$����+wG���z�MǓ�C������T���=��t�,5��sڎ�A��b�P���FX
^�z[s�>�����	��Y"0�{=QXY�y��ؾ�۾���w۞��;N႘-�K�������I��t��iv�O��}6vh�E_j��]R+Ȗ����I":��NV��F��c�1�p�� �
���(���S�(S�PvK���>����UT������~���عJA�p{������W����q�P��f� |L\Ku��+��Q��|�v]�B�+^���h>�����_�y����{~��'=�#}>��d���#��e�V�<<�k�����y��9�}�=Q�޴j6�[g#��@��k�ߝh�ٔK��z���J���"�d_h�H���T���Ϡ� �>�J��E����Tm������ȟ�_:�T�za�&�}j�ϟ\�x�<�̆,����T��Y�qX��o��/�0�������Y�1/鹥�s6�t�{�u>����h���6����d���1Q;�z'T���oW�\y]�aC���4~�`��r�*�I^��!��ޟ���B�^T�����Z�u��j%�����J��3:�E��n�]��P�g^_�C�W��k���x߲hR�T���Y;@��9����[�lq�}�����)y#}�x�{���:�R꽾���7�_нu{����9'/�,:�ą5�j$���;/a`S�g���eޜ���QώˁO|����d�s�Ͻ�q�Nq��gω�9��$�����E����ș�!i~G��O����%\{�l��89�3���6rOr�
��O�%��]�f3� ������>�Yo�j�[��#�n�h.ʤR���{#�6_nsVc食o��gWa�rٔ�ڔ��2�׺���	��� �w�
/Ж?U~�aۙc*�OK�·����z=>�{ŉe���=�UxU��~�}8�]ğC����4�;�����΁\|-����A��_�����̇�����Tiو.ͅ����Sރ5�+�*x��PQc�`�S]T�ӑk*���\}�=GwWwZ�v��A���w����l����l{�M�*�T�<'��(ʼn�C�y0	����N�V�>�{�븟����mӿiϼ���{��#g���p(�� �N{�Y��2M_�����C�z
��o����]G#��(�W�#���\}ワޢ7��d�n�~�B'y�/`Opye�|zH�����l���Q�������m����[g��Yǽ̈�L�Q۝��'=�ͣ"���	�,��xQ�Z�qA�޲6�V�~�J~}�"�����>�&x���~���H�Y=Bf��/��w���5q��!�A�o>mm
ik�v�,2|F-��������C��/�R|���>4}u��K�����̈J�ض�v,�r��͋ig1�޽y��v_[��/��hUj���K�2�t�YC�� ����U�n\Tg�G@�(|����e3�@U��Y>�Z��Z]�+��t�7�m�V �{"�n����8�
�Nb�O#�R��ɻ��]n�o
�����Fy3��\h����c�]~�=+޿�Y����d�����K]{��ot�^K�WB�g���}�Y�-��>μ��k��9��P�9�ʃ޺��l���Fu�[`��=�}�P�K'�>�.|=t{���(�'O}���g[��f}��D{��/";�p{���{*=y�UY�7y��ˏ��q��|F��P�P?N�qUYgFT��M��`=��/�L������Whο<����#Σz�4�;�ӼY;��X>��]�9R�<���&óK_S�lf�.]M��3�y�V��O��}�o�Û�t�J���ciBy�w��=��*`��^���w��(�x
|P����~��;��ǜ�����¾]�"C$�!x�tlH�ʆ<�������;'���F�w /W��O���\{��5::ݣ"}��r����K�M�O�' ��P����/����z��4��r<���9����q��~�$�_`�V�ȿ���O���lj�_�O��2�C5]w��J�^�"����3yw��Wю�v�����*ܛ��
p���n�оl��M�x��h�32\���G�㱍;{���^�V�T�W���yP��Ǎ��榔�+r[��ާ��\ha�X]�1��!�w��D�kT�r�>Z�|o9���{B(������6Le2ƣ^<s����ª�rY����"~��I���|���W��o�gzse��osϙ��}cޝ��Ͻ��&�~�������3%�p7P'�����7���7��W��sE>ʔ���r���}��#���lx�Q>�8>�U+����2�����m����{�_�V�>�^te�Go�޸���y1P�O��y��>�����@s$��N�LV�	��
��Ey���&}N
�|�E�������\y��IQ�|=&��P�A�k�c�y�m˽9���x���08��6�pz���<�x=�����yp����~���c|���پٽ��F�z��k����͟}��Lu�
f}�b��Jޖ={U_�5^@�h�L��W�7Z����Ok�}�{&�/����ƖN�0��'t�L�{NEJ��l���ct_�u-�kp��=���'���>��(�������ʑ_B,�˃0���T-��q�!�pQ��n�-��/$}S,{�� +��FS��IȯT>7��Gd<��t䝸�d�*ϰ����@�3�1�#6�ĭH�;�6�W���={Qt�������7; '��C�~*�L�ƍ�G�}hյYW|ኂ��-T����������h^4�t�ޢ'T�*1>��*.�r������\㒿?
b�hk)m	��ޗ�E����Ś�A���<z�is��錰n�×Y��)�͝	�wԉ׷�z��栎�j���)���C{-�;Y�*�J�%�s��,_[W�G������E�R;�?D���t���j��櫓A��2����O9*�z,�9n�	���Iw��Ǜ6Q̰.�/�����j�o���Q��E�w�kWۏ�v���)Q�#��H�9�q�~�o���e*�����W+��s����b�;�p����Sw�^�
�tr;���{x1�]�_B0���ۃ:M�������rv��H�G��eq�b���\V����da�y������>Kvp�����U��v�9ƀN��JM�T�A��^6�hY��b<4"�Η��W���p����O$Q�����f�s�x&��-u��e�c�|��]RG#�ܧ��g��=3���pi�u�s�	�@.����gm�6���ݾ7�y'Ԃ�rR�s��Wh����+*t@��RGJUIy��Z.�'̋�+�7�����h��l�s�N<��2������[��|41r��s�Ǯ7���*�^rk�|vl���]E�f$�<9Y�[��.�a��b	��׏yRf��9��%��\���gw5dӞ�<���u��'��V��B�n���m�32R�����G%1=�(���!��C+�9�VS��6i�4l��;e�u�&��Ц��� �[���ꋅ�bc�b���rO��$�.�0T�"�sQ��C�``�N������s1f[ODYr���!@�nު��8�WCxX�w��ݏ�g�2VyK3uh)�n�BB����Q6�U_ �����8�^�K�� �%�X,���9*K��p"'l��0�&/��wRw��S#�Yd^S�"�uF�c�GY����v��#���5Lk�tP����y�hSOX�S`������X�B-GX�e��1��n,�1e���*�k�(-h�D8w��]�����zM�f�{=��~*�y�7����Me��7(�� F�����4��yW��4����,,1kٰ�%�y��5{ۻ@�H]�S�
�������2�<�ɖ�Cۦb��s��m�a7O8۷�Y����q�k�ƥ7<y<���k�\�ܤ�����N�ծu���&��:ҵdɄX �[E���)�[[i�Zgc}wܗ_>��6,��94b�2���%,sTw1s�)'&c,ʕt�kܲ�gA���#h�8�Ē��!}���en����`��{��{O�:�v=���V̺�սES+�{����()��>�D����+�TT�D����S��J�J"���$���)2��R�r�nE�)�q��ݡ�l$ʢ�@�\�c�)"*��r9r;�'�,�9$&y婝;���/=��-MGtq:qLM2�W�Gs9l�\���Q�Q5e*�RQ�K*�J浗rY�:z��q.]�)�Ur�0�E���y���N+*�L��S�䨺)#�r+�&AaNW��jC�H��4*�����֑T���D(���t/7:9�(Y�z�y99��e���鲌ٮ����=��=wr<�Vz9�*�j��N$Aژ'�u�G���GEy^�f੢F�x]���(�u��ND^-�(�5�Gs"���^��T���"(�:*���NN�8� U{��,*.�z�W3Ԍ���wrv���"�*��

	%E�S&��c{|����w{9K��|��]�k.FJ��֢��N�QG,=�ʛ{@ˬt��6���䥨K� �:�R�y(�J��Y�e�)j�N�O�y�=�c}^&��9^>��C�^���z�ܧ�o2+�K|h�*��\�����E�$�|	�u�^���TQ��z�<�w����'��s�z_���OO��1>����8�3��o��ͳG!zH=Pe�ȱ�ԯ�UIg�����^��'�"�dn!������yI����\>���.J5� y���R�ȸ=-�}S�⍫Ή�nl�{ۋWi �	��z3��2�ʎ���uҨV.V��A�`'�����qhb�Rj5���׽���g�z��u�Tx����;^g���߽$o��PeL�< H��u�.��ɼ�מ�z%��q>���b��u�1�߭��x{�����7�Z|�ٙ�i�=�NZ����o�,w���zX��T���_������W�7�O�>>'�}Wa�V��m���x�6�ziLȨ��M��|:lT��X��o>�O��^���+�1�������rC<�𛖯R�D��'�{��s�V��>�$���0����Z��7��^*�^g��zv�GqI���:���q��B�0����(�� �o]�����/�P���O����.��<�\Mnz���)8���FRŚ��~�U_�6��<LZύ"�:�������P S/$���E�c&�U�vAM{2�	E��G#H�K��Kos�o�,4_|��=��^����`���F}���s��W^��P�-��ʊ�s�W5y���}�-z5[�u���U�9��P�y���ǲhW��R2�Y;@��԰o��C����ޞ]}芧|�T��x�.�
����}��Q�Tw��/]G\nV��NI̭[QRg�\N�YoAf�>�QL*�˽9�)���r\�u����9^���y�oE�w�
��ժ�w �������2Q�D�Bg�������C�rσ�>�~t�|�vzf%V����:���-3��߮7��#�vT� {���x�WUzL��?M��sr�Ⲫ���[��Q��'��=HnC�?���\�1]�S����=Fc�`�S]T���,�� �ۘ���s��`ߠם�X��z�/p�|���B?d����J�0�(��,���g6�Su����9ڂ�£�_��q>7^�\K�^���>g�=�G����6��0�R���PD�x��G�c����=�?+�`�����Q��F�+��W�#����}�Я����=�+��T�P«kgՄ�teZ�U��������/L�w����k2\��l�wNh���5���Ul�^��XP<�����Dt�SG�Oj*�[SIȫ��esU���A��4V�ڔ�E�n�r���c7x&`3XDk>X>{!��!����o`����L���<k�q$TJU���ex�n�:��Up߭��޶��m���d�oU��J��D���#L��s%��S�� �q�q\��{ac���Y~۸A�t�9����Zn�-��=������/�˙
d�	�^��c>���=�D���A�}�;�i/�<�^�.Y\?+�����?O��dC��/�R)d�|>#�0�Oi��{w���}���K���޸л�Lw�ߪ����^��6�hW��,�Tt���q��U��J{�U�Ϡ��>u�v��|�#�/��ˋ��^��@z\��*\{.��I�!��;��fjʿ"wޖ4rx(ӡ�V_�ĩ|O���o:�ǳ�s^��{��/-!�p���C����1S�w�w���Ņ�͝��*&X�Q��wU�teJ�ĭ,{��%w�Ǽ9���ys��}��V?V�?�5��I�҅m�qc�%����(dWz��� y�kSgi�n�O�ك�ם~?/W�W��+"�ǥs��+��'ɍ�V0���v��`�ȯ������m�/'h�qܔ�p�(2'cZ�4=���4D9�f���_C��u^���3�6�$2>�0���E���ܙ����e�H�L���^����4.�+�T�Cvt�]Nh��jn���!��,����^P������bT�-9����r����D��/�O�n���z�C����{g������ק��0Ƿ*�\��g��%\�_}F��՛w�v��>�9Q���>�P<k�n�/O���I�{�������!�'
���K��f՟"s��`�$�#�0�n�,k�>+���CN��<���9�>=��':���ʀ��o"�ў�=6��@�� �2��
|i��������O�]�:�����
|�^I%+)�H~���:V{�;�L�C�,�( %G�D�o�������l�����?{nT[96ڎ���w�G�z��z{I�~���~�TM3%�p7P'�����,��FVz@u�o�ާ��/ɝ�Q��\�׽lg�ԉ�DxΏq�Oʕ���(�P2����=v|��f��az��g���+��q��B}>��n��<k��C�]Qz0�EmQ���w��>��`|}zpT�V�������/��5��?;�8χ����P�}���Y=T��գ#3���:+�>��g�r��Nq]^��"���������^\,��w�'��O4�~hR=��NE����
34N)������t�E�<�;�|g�-�*������0b��Rʅi���J��y�6;E�������l��b_1��b��&�x��t���pl�3)+��|���rU�}z��/n�.@71�i�z�J\���H/����;�_��}�P;�Rt;3gt�}P2c�NuU���{6X�v�����;��un>���v�c���_zh_m`�ꙣzY;�f��;�	�����Л�1q뵾32��oT-��
�������2%ׯ��{վ+=걼s���{*E"�����{��w�>�\�t)�W����S(7�6� ����,�zK�T>6��GdC��YӒw���sgW��j��ǉ�5]B��T���@�9�C����>ex�]���/>����Edq�g�߸�.���Dy�#��"O:J�Mzַ�*����n�w��z�/�l�ay����>���e�x�-��ϓ:�j;�o�
)��`@�,g�ԯ�UIg���7�9�n�9mB�\�R�}���������\>�3lñrQ��ʌ�&K�"�=-���4�]���K�����~���_���W�z2��+|��W�z�a�J�E�����T��*�=賕������'�e#���F��\\z|��3�ޤ8��z����1Z�������cʸKK&����4p`�m����0m���W����{��AȢ����ϴ��mv�-�z�W�/X�Ε:��Y���u��ES��q����<s2�L�/j��MSS�.�}��b�kq>��۸J4��kw�UF�*�Z��W�-���N�0x�}��3��h�m��l�G�x{��'����=��D��t�mp0��l�x�<��}�X�3�l�2�xUҦ��/���Tm���oޟ"|l������0Ș}���X�J��7����s2���3���b�N�к�^�y�񸆽Q�Ԛ����2��[`�_&f|���td�\jphtd�B,���L>�>��vp߫�{��ۍ�˘eY�[�u%��W���p��]ȸ��������¬*5��Y�?Q�@�R[8|�4���.���k_D�m�����+��W^u^㑯�<e����ɡ_w��e�w�iɏxߌ���]r��3�Ϡ�=uY~G"�}�����o:��3�����;�r����n^��,�U^CTvD�{������<����QΏ]V]�x�Q�p)���K��ύ���sRW$9�y{ލ��\^{վ5�d΋��:v�X�<�uz��*]9ó��O���Juo�b��N'��ؾ{7�΃=)��z���|���jĮK����.3�O9�\�0(]�ӛ}�ښRp�Y����[���fԕL��1��%ה��[���M�Y*#�T��5v�mvbLm�v���˕Juָ���~ȉ~���8�޽r`wan5��Рr��qڷ���s딠�P��[��Nܝk���<VΜś�{ڻ	�g�*�"��=LnG�O�g����3|aụ�e�z��?2���wBs�^�p��e�=4�`�|��b�^��p�x�{��u����&��.J5�JN��9�Q_wi�&��=�1{X�8�����K��븟����\����=��#�n3ʈ�uL?Ff��v���Wݒ��<��@�G��7�l��V9�����z�i����>�8zmb�ٿ'=���6;���b��c2���>4��U}�"b[��t�7~u֩�^��O|��[�y�<�s�g��Ϗ�s=��{޸=~���-N����u1%yM��x��3�����ҽn�j��^<���H0��,��L�y���H���f������>y��s�g5n�Mf��޽���A��N���w"��x�g�����S �R��dy�K_���W�0���m��R~��n�NEl�ǯ>޸�����{ή�������i�{V*;�R
�N�x��Y�[�]���_�cQl-����r�|����>�}����9�@z\�`���F�����~���~�n���h��JYVs+%q��&��|1�زE�Ѵco����׏�v�[�%���F�&F'��n��kpf�ymw;�_R�����eѩN��iJ���L����@����cQt�����M��o��4.�B�+��f�F���G�ɜ��Q胒±���EV_��R��G>ޗ�y��=�K�����QH_ضw��^�ޥ����y��=�՚i������������g(�ڕ_�������snT�o����V=�h��ĩ�Vx��43z#�x�}��p�'v��<��>E��[W�vc��'�U��5ܣ����u�+�����Ȧ�~+���������ʝ4>]aᩛq�~����w{�v����.�~��uR}M��]�x7޲.=����e1�>�<4��K��lm��k��$_yQ��y��J��4H�>���z�iIt�Ag���z��#�'��{���ׂ�Vu����w��^��]��`~�%Ӗ	=_L�	T;�φ}����W�V&�w�9����7Z���D[�#����g=�p�>3~.��P@��aJ����X�S�*=~�+_یߋ^��Mly<|���}�G�ܯ�*�޸;�a�,҂U}DO�[�"�J��vG�|*Z���W.�'�+۽~3��lg�z����q7�����5�A'��x����t�������¾�贮ï�P'-e�j�o��y����`��^��:��^�,��������Y��>�Zf(�b�pI]b�
�{ ��c�X�K9�[N�n���c�}��*ā�Jvza߱է�`D7Hf=tQ�+Z��/�����j�Τ�X�5m��FQ�/a�b��d����R'���8v�&�R���̠>fj7�zm{c�Ԫތg�I���>W�p�m������M�ޤ�Ƽ �9�=�u/jU.��ͯ�X���"�~XL��n�Ł�s��9����/��^�g�Ux�/�����p��۸y�Ѧ_��v*8��5
c�M�:ǧ��\xesW�y��7�����:��]�����$,�-�%�Iy꠲}�T+=)ʡk���;d�="">�c):D����^`�ic@���y=���`�E{ﳮ�xg����ϵ���������
�3g>��홅�9����Y����՞ؤ�>��x�S +�;��u������5?oZ`������Y�/.��,�D�W�2�;G��2+�;�W��T��/׀���#)����Ez�N/:������i��\K�jSg�J�RQ�)6��ҁW�Uy��h��(x^�?5)��0��z�(�*+kg�j6�qS�w���p<�躸�<�J�%�����D��k�Xqޟ>�W�HB* ���\��5���
���V���2��o�14��OJ�m���*��r^��ue�5���6ޚC�@�FD�,���\��FKH+���E��n�o��]i�q#N�p���@"�8���Lv��{K�Xc~eޘ��jJ�Ty�y%Y�rϼ����[����B=�Q��$��� y3��W>9��*����"�yI�W��}�H>b}�lp�!�cr=�|z���{���ñrQ�GĔ�K�!����+�� q���gR��_O��Q>�~�=/Ճ�g���<��W�@鿝:�p.K(^�r�<6/0b�����b`|V�~�^/v��o�~W~�,C#ӵ�{cޤ8��z��U11~��<��ޝ�T=s�]��py� �>*H����c�Gؠ:�F�֍F�~��G�w��v=/U�m2�I�Y�Z��������w�_���I>GbO�l��2�RqJ�<;B��~�*6���K�Z�@��W�4KL�>�������%�9��=5f�M��s�4'�7�ʟ�8z�]2�u��B�'�g��ܘ�~~�&��}���	���&�OW�&X�a��k����	d�Ǿ�Qݝ��<7�(o���	��E�?P����O��X(Tkʐke��0�u�+KAV{�;B�7S����7�T����ȷ���8\Fu��g�u^��<eg�ʵ���Ϫ�����2z$#8�F#:��	�����K�v#��@xt���Y9����u�Gy���2�ڑ�XH�`�a�X���h�չB��մ�2��s�+P�� EXXxY�Jŗ��:���gf�Z|k����U�j�.�³'�E��S�����\�`
U��E�U%7ʸ\�<y�{=Ȭ�;�W���x�F�������-����[� ��R�7Y�F�)6�p�	�e>�.р�F`�������3��t"�9܁��v��.Ү��h\�(*�󐻝Ak�i]JrM'�[Ń�iM���D71����w(Z�O��<gN�c3�vTD4Uf�SP����ɾM+v-PSkCF����Oz[��wu��۲���3�u�A��G��۷g�r��<F,�CGmM��n��]$�S�uh9�y�B�:y7�'7��������қ�K�l��k����'mZ�-���k�K��fN:/vY�R;�;f���)��Ƿ����`�㻭��`I+yMyGvd����Y��b&�����o6t�˺�:�p���i.0��Ôq��Z,լ�Rqݹ�{H<_.U�ޛ���s�� vv�C�gx)�gy��C�SU׺�m6����z�=/��{~<�S�>��ݣן*XX%|qt�+{�ܘ�uC�p�M���z�٠HU�qkGJ��5(6�������l(d2r�K�@�BSS���\j��o��mJ��m���{0;Z�B��^b!.�U�/qa	f"���הeb�+.��x�� ��?߽Y]�����W�y�z8���`ig_fء�㽗)���lG͚]+���� ��IW;#���.����g])�"���%�$%���\�䳅{W������2��gn(��y���^v_)���]t���X�E��� �Y�֡�(�O#�݁���F��r����wB
��,]�c�n�HW5+�3n����v�9!�pH*i�Ɍ�7* �Ռb@��YVA��@(MӨ��r��̩�EQ�F�)�V"��F�ЩgV�qg:����4���,頌�ګ^p �"����#C�z>8��u��f�;q; E�Ch�b2��2�讲T1�J�)�wz��b�|<�{�,q�5���|l���Ҙ�!��F-fǕ�͙�7������k�w����@�+�z�	�3{9<�s	��<��tI����u�-��m�-VRzx5'�4��w�,o��r����V�1޲��ʾ��vlԭ[���z�J޴kABw�Y޴���Ժ-���#�%�RrŚ|�eŉu}�P���B�N�jY��ˌ���\2��!���Xx�t0&5�R�s�����xý���uZ�!�9t�G.w^�8���ł�jT�+/b��4�I�N��M�mѬI�H��A��δ3�-3m��)�y[�C��ź���P�����Q蓰��;�/��V���S���7��K��]Ȋ������ʗs��)�D���7�K;�㞡���9�*sqӞB����8E�z&����e�#�n{����VJ�Q���p%NG"��2�s�G3��̙�`�w]�Ȩ�:*f%ΙjjTUf�QEf\)u�*������뻻��r��p�R4MJ'DT�K�e���R���B#�f�8fy�r�Tw��ERy<L���jZDf�Wu������z�ҳ���9y��Ȳ.UQw$d[�z&�9$ʃ�):甫�Eݻ���9����f�N"���yz�	Q2;�e����A�L�GJ��"�]�M̧@���wnj�.Wԛ�ȩ$�����x
�W��@EUG.t�D#�繆����	���8E�c�Ap�����r�2�*�FQ�EJ��T��Z�D��wH�7j���)o��)1��ӂùc#�ܚ�r��N�� #֫�$�uЫX�/�w��ȳNU��� Ǣoq*�'@���w���Y_���=�pwj=qU��r*e�<rK��w�.�����;�r����[��H��G�}[S�t63�8�����5S�j�m&�vzDEL�ioȢ�����}.���U�K�J��Y����h>�w���Y���3�x�8�X�<���	.G���;>����k��m��3��i��ȯW�V|�\o9�c�;*t��Y>WX���>�n3�>X��%�.MWs��W��UX�|7��E�G��������@���R��d�����FٿxG��v<k1�-|����>c�N��Mz��v��8^�`Q��ϣ�D{���qț�
��D�+ۧ�n��1�;���Uy�x�=���x���|o����\����=��#�n#<��2��v�L��Gd�xs����� ��-ׁ�[/��.)�\M��i����*���]��&f�t�z�N�l��/;#mMx�9�Y�PB*�}DLKu����/��GZ�5�+޶�t�܃9�����u��zu_��L���ꃽ��KSf����D�^SBⓥ��}i�����\G�)����O�������A`�r�iv�o��%\�h�R�ݝ���>�$���K��}�(�����\�i�rl�]YϾ��S*T�"��K�����s�G6��ָ��㼹��Q�j���q�G �1a;��Ha����w%\�W�����������;�^G�6��ԁJY=_	�^����/����t���^��ѫΏ��<�o�>qN���w#�ω���ϝƉ����yg��y��Y�&�������&|VT)�;��z�z�񶽷��x�@z}��|�{V<���*��L���eo=���z|J����g���}�x�|��>�}����:� zT�1��yFU^�~���Q�A�G��T"�g/e��A�a\���7>�M��~.3��{v�uTmuG����Nun�g'�	L�+�w���Y�����|vv�&|?oֱ_�wOg�ɿ�?H�����9"�?�f�*���O����W�<{#ޫ�ռc=s:vd�٘y_	�,m��;p�C��tS݊^H�Rq���F?[�Mz�W��+��O�ӿYd�f}y�bϲ���O�垆}�U⚻�uޠ<��>�����q��Ol{)�<�������s�3�=5⫼��꧶�(�e/H�}r�(��|�|eT;�������f�5��y��W��O���\?)=qz0u��{Y��+��b�q��ꂯ��=�q�9ƴOg)��Iocqo�;��]��Q+��d���μ���O=����n�M�={6���A�)������t7o�����u�)�s���qrRt��p�J��"��U�����(4�`0�ܺ�G���)���@�.+<��&�p���>���`H�w�M��t|n��7�N��z��=����8�B���G0��)>=g���6˸�F�P@�2��
W��l����N{�ܜ]�ϯouv���
�uu�����؏):U�����L��%�P@J�>�'�-������Q~�~[-vo����N�^�Z3��lg�z����q9�T>�LKfK*�����5��qW����c̘���u����F�ֲF�o���O���������K���}���ot��^�9c�K����G2{�Q��>G�>�p�|��΄��M��z�>����FK�Z5�m�<4�^o#n��z�ɚ����񿊜/�ENJ��:�һ�P�URM�"�����e]v�ᾞ�ɓ����T7��d�)�T��:ǧ��\xesW�y��{�ʅ���"+��mԿ=���a����>W|c#}�I{�w��e����E�}8��iП��7�-�f�wb��%{U1����{�3�~��{ޫ\m`�P��8oK'v��0��ӭ��g���Ѣc0�����A����Vٕ| ,�N�n,@P�-9(�	Ppf_Ve�X��jj�����5�Y�����f��3i�Y�(���l���<�]p�,�ƞ���rXʊ�u�CPQ;��N���5>�KGC%��6�Jlu�1NeRG�T��{!u�{�^
%ׯ|gcޮ�x�V7�v�
��T������y�4{I������%ߌǰ�釱Kn��L��mxQ���"Y^���}+�tt��Lڬm��ڀ����phܝ��C=2���
{�Rz�\3�� �4��O�^>��9�Q7we��W��:���>��z��{!塜nN��I'�&P�@���1<�ѯ�a�t�S7���ʿ_����������"������<��7Ƒ�2�ےQ���X��W>.�m�FJ��,�Q��FV�	M�=C���{����;�vA��q�(������7�w�MK�ZK��A�s#�\���u�O����"��?^��>�2�����@�N�����l���p��q�K�u��t 3e�4�Vx:�G_�D��^X�zv��lG�Hq7�{�G>]�gT����U߇zD�=2zi5�D�u���h�w��5֍F�~��G�w��s"�k<O�^l���r�f�jo=@�=ՠWM�4�IL�-�=$L�Rt��ô)~7�B�e����*��2��._��U���@�}u�; �^������U�ʗ��w#*�ѻ�딃;[�X��	]��aKlۨVQR�7s6|zÐٝu1Q?K�n���7t�#���N.�k�ns켘�����
�DX�>k��
��P�5�Rﱴ� �c��"=�!��w��h�9�3"�g��30�p`��=�Bq��~��ڜ�M�	L�{wu5�G�}���p����Ǜ��6�>���K�?�4�j�R����5��B����'�[�nߺ%�����o7�ï�����\c�L������`�Q���d��[����y�mg쪯G?	���;�9JZ>{�Å�g^_�G�W��P񗑾������#U�)�!y�;�F��5�Nz���ݨwU��r�_�K�η~��=2����n�֝N)���-�K��;'}}��$����t헆~>��.��+Ģ�ˁQ|��6���v��i���1�^c�7�:��Q���%��~GN�%ᎂ\%�uz�����Hwgy�}&��ois�0}"�l�}Լ|W��+!ڸ�sh�FuC�>��}��P
x��W������w
֖�[R}M���q�Xy}^_�z��z_�?]!�f��B�F�OV��~Y^{��^͌o#�,��֋�U���E��>�o,C�޽�}�=�G����qϦ����2zdY%�L�LW�Y97̍��W�>��9�3�&�$��Δ֙(
�H�7L,Mj΄��ul�AIջh44�J��{R���h��s�6\vc�^���[0ª��ԩ�q
r�z%Yռ�Ӣ��5%�)��T*�:�҄�Q��+D*2I�.����-�Vy�,"Nz'ʘR�i��O���Q<�ߴ�y���I�K��b�������z3��_��z�d�� ��K��7�[/>�uc���Q*=^��AB��=�'[�h�s=��{�t�������4��9�YP+g�Dķ\�:_��=�#b{�.�ϻu�}�����c�:�.=3�M���_��dS�-+��{�C�
���c3	ߠJ��u�����{��Ϗz�ǹYq����O�������z�`L:u "��&��+�^��>�[��^��6c�n���VJ}7�X��vG��+�n|O�xπ�d;��u ���9�H��N{w��x|�p�>=���V�-���p���{o�#�utn1����{��8���q����z��S�S���ʐk�Ī���
�}�>�����}��m����v��T�O��V���^*��xN0���*_��W�^L�����9,+:�e�nE*h�sz_��dn�O
����^(Xh��=;5�P�~��ު�ߦ����|vv�g�������^���Mv߻�a_vЏ.�A��]�|� b��\�1�ҫ��a{@B���{3�4�T7R�hE0Un�D*V��J�8��ǽ���sM�5Lw���4�~淝���j=��8�2 Ֆ/W �6˶�0J]�FuM���j��
)u�Z=��x��^�^���#�"Z���Vx��43z:��g�gJ��f|)o�*m�_���.�:4=�Z9�J��^��ȗަ��^�X���?Cud�Ly�;����0�W�OZ�����5�P��U&{�Nz�C�����+ޝ��z�hxw�<>bz<%���R��1���Kf�bJ�9���C������Z�������{N{���I���A�~��aj�%�}�}	��� �n�+��T��OT�G�C��φk�>7^�X��7��U�\��<�R�JA�#��IG�s�t���}�f�v��( yT|e����-����ku�w��B�k�gke���ֆ���[Gc�N�q������LÊ%� �Q"���?S��dg+�>��CŹ#��^���_���lg��޶;ޞ�Tg�px�z�Q5�2Y]�ӯE����Ε߀����ΗG+�#���5�W#7�ldG�ԉ����|������}G<�N���sV=��D�ӄ��F�I��F�KG��~>LLoBj�&��� |�� u�m�nt_�n���g��v�� �w�fS�Lu�tѭ����Vc;��� �>�ȸg(r�8�]������JI�
��K,E�L60���As)vK�;c�ju���Q�TҨ���ٝl�L��gtW�;7�����>ȸ)A��WQ��r%� ��_���yuQ~'�%��8��Sr�vʎR��^�^�f*��ӷe�O����'ْ��Gt�'��yT�}�%eN��:ǧ���ǆEsW�~�Ѳ��$�n���Gr��|��c#_��%�o����Քt;3g4�}P2a��և���׷�ܗ�V��b|�����L��oSΪ����^�~����ϢJٸ�7�J}k��0e!W�F)����;2�;F}��0�Yo�EK��#U��x(�^�fwޮ�k�C4�l�ɶ:'�<��܉Y�Te���o�<N����4Z���-��S/ļ���F??d�e{�g��go	�p���~�����~�?�g����TFt䝿���D��Pg��]��M�WK��p��i�x��'}w��\�]�yez%���gs֮���˭���\9b:.�ȓ�(?:	p��o�1u΋)���ԯ���u��;Wa �����߶�����ޥP��f��#�e�rA�,	�"���|#���r�����e�O}o(��?U����~3�z���Q���q��3~0�\�j�%o'0�׿$�>w[��/�\���E
'.�0޾��b=�퉹�Q`�s����ȹ�f4ޢ+�Hm�J][���qΙ��R�]E�R���d����A����59���ĳ�6�-�Oe(���܃D=�r�Ͻ;�j嚱M�[���F�R8�"�����"ϥ78��'��{��G���tG�W�[Tt��� tۧP�e�t�"�D�R{�{pw��G���_��~�&�J�{�F�z��'��h(��y�z��E�5ϡ��>�����k��g��z����2}4��>�&%��lt�}�F�zѨ��M���F<|bL�e�{�����}̾>��eOtY1�y8�����(}�BƋ�oԅ_ԩ�ô)~2�\'�\׷S��^��W�B�$8�Dv��7���㞙��82�d$Y�3�V
�\�� �u��������5��/[�~�Ը�zH��w&.<߬ɷ���:�'��d�E���ɇѦ��V�l{R�	�[l��[z=�w��o"7�ï�����c�L�����¬*5�H+�Q�#���W�ZIŇ�K�1���S>�ñJ|�����8_�ח�u^�k�{�t��6/1����7W_���x�ȿl�v���l��;���#$�'O.��y���>�U���O�\z��V�h��yZ�{>���O����MT�j�u'���芙�Q2�J9��p7��7U�,�6>�O^b�������B�~��W��_���߱���kiZ�|s�s�8*�zV�m\�9���i���׻W/b_J{��>��~�_ؔ����1��e����� Hn����YEb�.�s-�fԭgX��:b �9�odW�b��p�76����fw��i��W�<{>���,U�k�KE������1�K��|�Y��W��6���}�;�LVϾ���ק��oΗ����{�c�q��:�b���M�d�Y�3c��6-�F��A��7���{�CxX�E*��-�e�>� o�����S�{�ߌϿ[���*�ө��<�p �(c�,�dl���I���φWU)s����v��8^�`Q���u��q���Xe0E�{�j.��{���_2�.�Ǡ)`du�
ֻ�����n;��2|�rҝ�x�ٽ�Y�s��=��C��^�#Tσ��H�<�d�%��<e��V9��q>]1��<.���5�^���s���{�t������g~�24��UO���끿�K�cko��!_�k]if�w�d���w�ý>��?�;��؏L���ꃽ���dT|�KSf���== �w���M�f��sC�S�^=��>��r�:���1��+>9����Tl	�ө:~��=�.��xv|5*�E�'��DJT��d��yʡ�ϕ��s$kJ�-��������,c`���X�����c`���������l��������6���6m��1�cm��c`������������o��6m��6�1�cm�1�?��1�6��l��c`���1��o��6m��1�cm��c`���c`����(+$�k**ʗ�:R��B ��������(/���EW�h	*������	
m�� +J5��(���mm(s��VUZ�@��Z��U�6,�32�-��6�����@m�l�R�Z���l���[[ko�G+e�h��X�ڢ-���kJ��E�Y�%)#U�_\�(��@ޯj*�ܪS�b�&t�����\b@���6�;��ZݛFWݧ��-�q5�[� o| �� w]�SA�/y�  �p  ��   N��^޸m��j��ش�1�e�T -�/mu��7q�h�6���z:/Oq���Q���n
{k�<��۴Z�V�,̴>h �tעo�.�㡫�����׷�N�PF�{޵ú�*�i�x�w��+�Y��%l؛S�@�Ϡ�ۍ���M�z��`z;w�{�=3���zkA��z��:���� �w�W*��T �� o�P�5c)n立s�������i�O{�����{�<�������WB�bSkя�����l_=����$��P7\�
c� �@w��cݍ)�`����H�bŦ�} 7�{aGI�n�C|n�C��.�7VdU�lK�Xκj�ă���sa��	P� ܂�ްfed�]�l.�ݰ�4,�e�r]���'m�iiO  �{&�9ۡ�l�m��)l�j�� �sunN�����I(�Q@ �P  E<)J��0 &   � �{C
TU       Ohɔ��        j��	JI&�4  d�   �E)�F�M�bL�2�OBi�4�bm4��A"@�M�����#5#@#W���;�~���<<<<9��߿w�w�����u� ���!C�HB ������!@	�@ ��)��S��	 _xIz�>}u�� �Q?��e����o��̇�a�I6 ]� k������ �Y ��!������0	b!� hBI,i���]��6~�ǿ����|ß��B��*��*�����B   T� ��$�H�HV@�T���� I+ �T$$�Y	 V�* T�H$�
� � 
� J��J�
�H��, -UUQUUQUUQUUQUUQUUU�����7���O<=]� ��!ú�&�*wg�	�7��I��ؘ)H�w���˝�6�wۻw�4;�Soj�`-���^�g��}Y�� K+k��kǶ���}Z��*���oEZ�4�j��^l�y����B�SM�'�5/J�ʠY
��+ZA�i���H�g)��ѐ3�l�;�-�Ӆ�
(���QaB#����Tr�[�sm2�URf�(���]�R̔Ӵ�3p>�Ȭ�K(�'>;��r/��/�(f譢��e�� �9��V�"`o��ְ�,�9���O�-b��=Ŧʫ�J��xf��F�W���4�c�wo>�RWe2w{z��&^���t,] %YU��pX�b�ͲL؎h�5��0,��nBj�zF�Me>OEzmYĵ��U��>�\e��UƷ�n�U�ln�5���1]��MCGt�X�Y�FY��K[��'�&ԫ���w��(0��oRy�tbÊ����Q�L���f�ۀ�N�F�Yp����Nq������(�r����pԶ�x�ִ��yz�-�񗊫u�Jw�`�����镡o3@�da���{)i���2�:\�i�C~85���8]�DBcK�g4�sk.�
�Ed��YPE�x�k�.��ܙ��X�91�v4n�j��Lb�܏~p����;�u���K%��0�g1���7���qX����ѥR�L�yU��G��M��!{U/�KȨ,5��ٺӅ�wwt	�[�
0a9��uPSI��;��q�T�WV�����*�=� ��;��+�Ϧ �ɚ�3Z�ذ�
���@`|���1[�]!�K��E���YsK�������=��2�ᦤк���Y���׊^U�wx�Q�bwH�f�FL��o
4��Y+J/�,f��A_#���A}�g��oH�Vkb�B�b��J���4r�n���f�hu[�V�f�çk���ax�%&p�F�`OR- l[���U��\7j�]V�uO1����P�5c���z��R��$��d�3�l��B)���)��G����X�T�F�=չ�-ţ�x���4��K$�^b;�7��Ô�J����0Z�,&�=���k���9N�2�ba�����,j&��/6�j���쬪��)�*��w0A��sv�1b���M�[��L��؇f�.G����2����xdV�M�;�OJfSeoլ
�
���v�m25ѿ���1�y���ie (�$u�VV*�#�>)�RP��Yh�r�'�W�~�X���q���\�6�Z��]嗵̩���}{���z��5���t����[jӢx�5k�g^-�m�`7CA#R&y-��ub��,��UHe��ڼZ�4/ц����ճ��	���(�43.'��J���;t�xVhQ�w�hͣ{eǳsU]��M�e���#[T����Sph��RET%f�7�I �"��,k:O���sl���-yg8����M`doQ֫o��U�RIV����5����zhlr�^1���Hٰ��M��]f���Jcn�Y�[),��3nfm �������\�Uu���q�z�+Y��Z�'� ��N-�Z�ǔ�7���L�e�a9������V,m��G�[�WYkNP�h�n����֮^�.�ݠ��a8m�C�35����"Z�ۗzp�J����K_^��ഓ���\�5��#5��+m0��3�r�*O�s�J��v�� +��
�l;�����/%lf2�94�4ʬuv�ڧ�#̧����T4c����l��v�9� C�N]KV��rdt��2]�vB�ռz��6�^��0#m��1�úM�z��̓uʷXItA��+^v|�噂���z����"���m +���8��D6����B�^;xwt��d���Q�����ʲ՛�W�)�U�Sˢ�eB`��)1�f�bCr�Gn�%��BF��Hi�C5S���ŀ�V�PHR�� ���ǚl�]��p,5���^=�^M��'D�[R��D��T�q-�L*2�fl�Lٚpcd��h��󷮴�4 ԓ|;WI-Ţ�rxM咩vY�{uclY1�2b�Ҷҕ%m��=i��b{u`��J��m��k��ܬ	uB:�i����P���ݻ�F�%��[oU1h}�@���g��Ѩ_rua}f��<t��F���{����-���_p�A�	�Rҩ��@�W>�AךH��2��T/���k�ו�Ov��!.���6&3Xx�t��;F�NZ�ՠ�d8n�����0��d˘�`�#�V�mY&�8��ݵ)�{_)W�a��ufGe�F-{hHN�`�cb:uu�.�1جwmV�6��7+�$X0oڙU/*��`˥���`���x+vLN�C����b�פ<�Q�6)����A�VT�5��Y����T1�3,0�]�pf�T6i�6�ok/&�	���ж�`N��%!��GqDj�nU���Mn�Dm������v���<q`��� �Α���5(+DZAM�G�gj
��S�����A-����ʶ׮���5�W`���7xmʸ��CqfÈa��6՛Zs��aۦjS��f&$:�7���s�l��Y�wN�f�݁c(<���˗�.$��V2d�p3�UXY�8]R
����~��w񼻭��{H���R86�,�ێ�G{-�d�Ouk��hvՎ��Ln^���Y��6;�VX)�qde=	�{|S�z7��[���`|{Q�@�]mSj:sY���1���P.�B��Ue��V^^ृ!'-�u"B�[�F@�wi�3���r�(c6e��Q��u�����Y��@�+�%ٖ�D����荻���،�%���W w���Kn����{���^SF5v���]�^i��r�%v��j��o�҄����m�5�"�G�r���,�W����N^���95Bd���j��A���XEiyZ�Y��aA�]�T�^E�/Q�ע���n�i��n�@�!�-�+jĥYUmĠ�,�a_c�ǀ�5�\����2cnJVYt����؂�8��/H����ڦ�M�����%�5��n�5T�]T�����n:��q�5����f��y����d�Y�s�gr[���sb�J+s�+|ҷ��Ր�|�o^@P��i�(�l
8�-b�+��l���m
E��9����C3�Y{m�sR��MO;��=VZ��c7]��Ы�E�sr:Kt`�+��n�gv��F��x�+sյ
pD�IgM�\Pm?�
'Q`;���kN�Ih�-�y/r����kLګJ��2Yt�tX0�]TTfV��[��D�<�{ϖ"�V����\񭴑��ծX�"�]<8��V�t��]�P�-jj�0�:���}�ҩ��_Ϙ˘2�-�IQ�yR4�=z%O%��(k־�蓴y�x��^f��-8���zTRb˹��:ƍ��WDl��
�����ATE<���^��v��}y\��E�(yv^e+z�kCDX��:C�ȕ����k4+.��p�R���2�	�6�����k�<�Y�J�V(���:��GC�5Y��5usq��0�իܼ̪>6�f�G�h��q���ta֭Dm��mEN"\��LFc$�s�z�b%�RFz���I��T?��'�+=>���~��wS��O �>w���Nϳ�T��O�q����:�w�Ǭ�=M����d�`-���:�ٙ&L�9��:��C{ʵ��$f.G�O��jM�z�![}��`&����,����f�P�8G�z�����t�ӕ��f��Ǩ�S�ҹ,�osDӔ�����5�6�����XWЪ��/)p%n��C�4��oM9���bB����֐ܝ��m"{A��/F-JIv�p�vq'�éÊ�Va����D-
Wۄλ0�����se�n�S��H�J����AfJ�*�<���"u�z˷
.�R��6�B���P��wɪ�\ݕ���pK*;dNӫ��lgڼO�	�̖B�I2��J�ny*�򔺐緛c �=��nW}n����@�%.coZ��>�wGRѦ��vdd�A��u>��$͂�)A�ͮ�Y-��`��Gpy��]QS���ź�E<os#���C���%b��e��:��vٌ��y6�w�r�Y�ĩD�)��E��:8T�]W-���I�ԡAtGХ��06�WB{LAe��uΉ���S͘���W�*L��ކpr��#�T/m�c����ȏ$�tt�Jw.M��f�V{I��ӗ\i�|̆�ﲗ'Ύ*I�͸k9�y��=F^���5�]��U�7�:�(D{L�YЮ�ژ����Ihty�yDP���շ\�ag^C��â�]�|L�~V�N��B�[�ٴ���q�]@`�/�e�b�1�8$�p�}��W���:om(��ĭY(�S."Ċ&~��w������Z�KR�풦��'�������L������`�_��jv/k'&l=t���&J:��}���עP��bm�ה1�6+@��W�.B��I�������v�����*�x�2 ��kǱX9]��L����.o��F�/,tX��.�w:��6�+u�L�z��=���5�MD��&0v�R���>��A��́sx�V!)i�1�p&���S7n�f����۸�s,U�>��,\�vv}̢�ZNV>O�&��
݄�t�2�\Q�t�����UM�?^`+���J͡rv#9���0�otKZS����+�3m���,�����7R��G31P�d�<�%wJu�9nu��ԡ�L��Z���r������r���U<�ӛ�`2Iٗ6�jDLe�-�!wǮ��7��:A#�r�q��UrҠʉޓ����͕ͮ�.�Ț�C>��5>.Q���{�]��EyW.#Z�.��y��[�`{�Hۑt��e�$<.�U�v9�!�	vp���R�땆�����\�ժ]
m��m��@^v�$嶾�'qyn�hթL�IQx�ʺ'3�~�f��^�ͼ�f���m3�]VjuP� �"dfkD�Iڛ�����7z�ͮ� q��8t���V"����(m�&l1�[��̢,D]�x�涒�$C0^̆�p�j�82��C�%Y�]�GF+��e* �6q�Zn��:2�+�4�4�B�#eıN��l]�����/T�ݧ�P6���T4��pe����^��,���7�f�ƺ���֠�6���i����OC/����ikV3�iV�i��� h�j��`��l��
ft�nc�8f���a)N�w֌)2�BJ�����KgQ�-b�n�˪���	��6����J�"�a��66�(Y��V�6�Ι�v������<37��(���Xd��ЍDӨ3�e+n�y�,�D�&KzD��m�t�[�����L�a�)uy��y����[�����z8�]J�B�؟o_r\]ٍ�J4:��ɵ�FȘm")j<\z����<�v,e��L��C�(3����ض��Mꚋ��݁
]��\&6��B����S�j(F�_w�M�e`�����E�@��g�\���F�Y�u0zQ��sS�4�ޝ�B:���S嗣�[,�����%Q�o��� ��6>�eOD�3s0-��/���w*��'U��+3D"�v���;�K�e�K�B͚�ɻ9���C�+�	d���Щ�8��p�&}�keU���h\������il�+���$
�fa�;U�y˽�ORi�׻�h�F�J�9Y�7sL&�3���{7_=z��b�ӝϪ�#�]}s+��6�;�F�32�2a��t��I��d��ͺ:͕�xPo*�.�أ�o4,<�X�Ҽ�Zz�;�j:_dU��,�a/�s���S�����u7ATS4��i����t��8��V����;ZN�֞��k=H�[[d��g����u�ux������f�H�(C�h��PN���	R���E+���/{Xh�p�dcP�dJ�t�T���l#�2�e�,kT=��"��,#O�� IY���=O���GX�י���]٢��ON@�SxZ�ѤfY2
�#v�X5e��S%�zFiƘ�E�ȜjgZ�M�r
�|U�t�ojJ��Yʖ�����+~:yj�LP���}��ّ\�0҃��$;����O���"W�aիm;�2�sqR��J�#>Ot)V&1��s������<�2���kKtR�]���nN5���ӗ�Wbvnp/C��8��������m�m���G~UtL���P6w={�۳��ݧ�A%
]��Ml������j�b�g,�sRQ�H�b�í������A�3~��6K/g2W!Ha�R	e``@��8��7vd��g�ٙ��zd(��Or�3�rt���t�

B��=f�b��s��d��Jh0
r����.�i��䜾AnK�R�������{��ݫj��ȾM�3K������{�=}]�VAu�(ְw�?�5h�(ث���{	i���	%�ǅ+��ZƆA�+�����@�AX���B]�Υ�򘜉Z��kLI�1��*(��3�o�$XLU[V+׳zޘ9�E�����Y$K��~C��,�0N&f��%	�5��a0��b��u��j�buuR;ң)q��)A˫g���y��Lm\����$=�2;�+<��I�Y��w��|sOT�"����S��B�9���J�ޣ�ɸ��YBcصv�("n|��$��aY�E��5vã�N�8���:Y�6)�#z��d�!2>���2��&���|+;�$���ݪ�
qԂ^9�!����u��lٚC���QP+|�c$�.>����m����Ս��D'���#��Κv(m��7
����E�l�=��3z��`d�u�r�W"��s�C4f'�9�T���y*�����#��3t��I:ð5�*r��ۻ�[ʲG:�H58Շn�a���ͼҙ������e�A�sn
�t����.dٶ�+����v������ɝl��#6�Wl�#�-��R��ӝ��r�iǤPWr��`�2���	WIZ��r�ǐto���2��Z����2��X��CӸʎ��u���a԰Qn�ˇw�N$2#���_vM�KM��с\�͋q�(٥|\x�pH�Z�����
'd2��������5��j໣�꾬A�ɴi�\z %ZOnMR��v3���J�8�Y�88>Lmp��`�f>�ftw���E��˫��__7�3u�<yVufN�}ٙ�����_�}����q���?����w���� �Kg�{�9����4@�w���=�RO�_��V��!����I�|O�3��=ޟ��?ﻟߒ�i�r����>wz~����|.�R��Zb�[;T�������&z�9˩^;�ٮ}�gU��M�g
�l]hΚ�s���a���t�����;t�%�	G�S���Gk���Vˡ��z�\ѸG 8�Ò� �aB����9��I�Yy��ͼ��Γ��7�]jҨ�o
�]>H	�%�w�*�����vJĖ�R�����irA�W�m>ɕ�jZ�n\����v�[��ݎ���fPYW��v�K��:łފ�.��P�Te*%We��C2�(]e �I\�k�tiP��.�rD�yR3t[��T<��}������h�wf��zԚf�%^�e�0���f˗�֍��mDUM!LW]G�v��� �T�).LI&I$�I2I$2I�I ���՜�`ٻ�8��ЬlSEPT[��NXOk6��9gm_�b�J��#1�s��b̙e)�-Н��T�b!B��bq�!��L��ktq�g,��b�&9+#���U�TN�t���<J��"��!�����a���5�:�\�Vh�����Sxp�&L���"�[[k��f���ot�ԕ�_Ke��c�;�>��Zt}	���;�+�LLp�*_E2Z+6��5F��*i�+�QŚ�Q�)j�m��b�JT�W��W��o�.��*)r�M˵w�W��z'b�Qb�8����`�]�*ͪ}:�ɽ��:��iOu�ZvL1���כ{Ho!	���Ż��3v�d�$��S*�a��'7��*g���T��K�V�WwjI$�R�I$��$�I2����x��B��"��N�-�2�ds�Jw_5z5;/RW�[X���IbSG-�gc6u=��'!��v�vpaJ�ڨ�Kd��P��+.3����$�����V��+�o�i-�ڔ�ԅ�N���-e�� ���tM6]�7�[�Q���I��e`�T�(�	ӹF��jT[�M�5���Z�l�CksV���Y�`�7%�:�<8&^LM�9+m�Y�_in_�ܡp	���溷�ܼx���Q��{��M�A+���ٝF����N,$<h�˷A����J�j4�D�偘R��
Ae�ڽ��yFr�{��=��ɇ&�\�ҡXհ>�0�[�z(�eލ9%BGi����%i����	�����gb�`��k$$f%C��:^lV���5�)j�fg���RNWY�T2�y*�����Ǣ��r�W&5�2�`I
��L��wJO�-ū4p�7f��H9�lk%r����Z���;pf*���aB,z	�s{U'+qX77�8І�k3���-;�o�UH��I��Yލ<8�7�M���;{�LT/��_1��8a��H�=N�="������TK:OTw�V�aЫcZ�oo2��A��h/�ߘ����ƣÚ�*�R]
�a=�xu�n��w� 9R�Ē��n��l�-:J�I)��z��Ȗ͡o�n<�Af�I��5:Z��Z��y�r����Z�=}&me�{ T�s��Kӱ
�s0.��B�l����q�-��zz}.���S�K,j]u�Z����[v6饑u���*��[��$�}�`7B�$���^Q�P������V.��F�M�9%a����7�L����
��Ų*���0�w@��/��7�Y
eu��NZPXe�g)�1iX�η%�؍�t�5�Y�����]Ҿ��u�j:�$[	A�W\Z�c���m$�#s��v�W��ٸ��9Ȓº�쬸�tG��C�#�ehՑ_p�B{s�:��cwMQ�Ł�`9j;.s��ʢ��������H]k�:��zcնo^�ێ�E)���Ԍэ�[�]Qv�s�GR�ݶ$�n7n�ҙf��Q�����7v*�ή@EL�GFH��:��\A����m�g��z`�u�P����4�J�3&��հ��BU��=�c٢��c�9�T�ka
�!�_�l\"ʪ]m	��Nkv��w���ָ��Y37Nu�.u�/�M8Zc�K�K9�E�F��ټIN�mj���4��D�]Cu%� �8s/�[Cnj[�m*n����c\�x�[�I
;ϭr��b��a'+m��{n�h��2�h�I��u+���\W���-��.��;�M���i$���x�<E�p��#���o����l&�b�9Ǔ�3�򾼫�Y41�4kP����^�du
�^+��}���bԙ�j��7I^+���oo4\I��l�!z�*��5�Ŗ���[o\r�9�P�Eẋ��G���4�];įw��M�ʻL�j3sZQ�� �aV1B�q�����j�a�{�>��)��'Cuw�*�F�l���'�ct&p>��|J�LV�m���	�l����J�7M�X��W�C
>wZ�N;�!�ۮY�u�ʷ���z���YCti�8�Y3�T�^w�"�8�	�(�9�z�����n��ѱV�,Z��3��jN�4G^2C���Hᴃ�e��-�OX8��]kJ�W�UC'd�4�[Ef�El�����4��r���0&�*V��	��Gjm��{"���ֵ��L+X���;jĠ�5�] ]�v�aKͺ|Ug+*��b+E� ۣy�.RX��w�ա���l��'�D�;��^#�)n�$t9��e,�R�ŕaR%��Y(���l$a�A&�{���*Cl70��쪩L��捧(�=bd���^V����;)T�T�4u
�aFx+8ﲛ[�ɺZO .���n*�D��2'�ܢ��;T���ۙN�����\�)�y���[�a�p�Ć��[m:j^��ٝ�g�U6:c��a{�͒L@�
�e#�/wXԐ�Y�mD%eY���RZ��v�)�9qY��BB�r]G-���SVMtq�ҙ����U������Ť��V��Y���Xc9��X��Ao$��:�!�g4�tK�ʧ��}!��aw�aW:$6���uA�,���f:��n��J��!�B�Y��.��I�F�#@iT�9C�j6k6�Ù�)�73�+����um)��m,�n�̥�N�0�+���b���]L��fYY���Ç���8b[��0�Gu�:=�^���|&�[VȢ30K�V�\�UmoapC��9���e^�]N��YtC��H�'��gX7�����
�e%(�h�ڠ��EP';���X�'�
}�@c̆�6B��Q�i�a���"�a���r����6t��d���w�Ďn��K���g:���h���(��kT��F�YH�V��g�5����ͩT�}��+�p�s�Fq�������f=�u��3�s�;����FϘ��h�i���f�9�����w�屩o��Cxgf�	t��h�[J��e�=���)���}��e�Pe}���1ڝ�U�E-���n�"z�Y�/ln��͔�b�Kd˾��vc������kF���3K��}��U��IT��JCM�С��]\��2\ȗW�hܓb_�2K�ZYq�^K&f�ƟY��mfv�,�$�v��t{��+L��˖�N|�*��&��-���a��mێ�R�1p<����Q�+�  ���H�z��0�Z:ܼ�8*�94���H�ݎ��2a�y�,�7k
� v�zzE�\;ȳq��F�[�=;[�܏��W��~�ߍ{��V~��a &�ě�B�4>��ƖA�3���s���|��z�{g����j����yx��Yz���=ۼފWa!����[�{�^���;d����a�9O��ޙ!1ۤp*�;�B�_F���YΨs)�L���ő*2=�5u��1mN=ٻ��K�3�$�
��b�b�X���yC��-����՘jOm�E&G���Se[N�~�4�Z���lT��5�W�M��I����V�d`�.,�ObWf�ɅY!��3��Y�2��	.C�(����1R���0�-�I�;7/WT�Ń�Js�����]��z��^ɵl�ގ,��P��#�-�7wSP�&r�v�t���N1hn��/v|�]��n>�H���v�{"��y.6�[+�BGV\�N=�b�	��9c\Tl�p�J���.ղkgw�bD}&"���l$��?Ram�nW��*�n��׿~�t��b����(�l��+FХSI~J���%�p��'D4����r�u�	�Z.h��h������*�Ůל�U��9P^s
e���lav0lۮ+[Jsc*s��Z7��-I��4Խ��sm�Z�TE��r���2!����^4�s�	��n[����
���k�.n��
�3�Z�UD����i�;�8rpn2�,�,�ۭEn۔�q9^$p)Qv�-���kȨ���r��C�k~��?�+�����o��\X�Ĩ\蕼	�Xe�����1�;﫪N0����s�^��A����~�����d6��ǁ�-F? W<�a+��͞�ㆴV7�!��&8av��e�xfq����Y��&�B�ªͶ�pyv@K�OQ�x4+2g�}��Qҝz���"��ʨ��r��y�i���#]FNnr���F��X�#�^�ëi�/Jd�@���8@3�E����]U=u�d>�R�5��f�k�l�'b�:q��R�Y�kIf35�|��� ��s�d�#��&3+2~hf�;�xAh�L>.�nkV�H��i}8D�!s�n�u�p�fYLT�c����������J9��T΍�������T�7!Ӛ3�� h���[�;4���_U��h��B3����}a;��/+�2ʾ�<�ݜ��)y��r�2a�c0Ȏ�⨶3HДU��dJw����bJȢ�Q���������.��#I]�Yj�t ���pЌ�
�Ԣw"nx�����v��8���2`]*�נ˺d�/J~r�K�3�������7��A �	�#[{�L��3�M]o0�V���1^�Q]ea6��m�9�ɛAĳk�p�@oG^��Lu��V�`;����i�%�۳x�r��u�%��m�qN�GC/�������N���N4��l�C�<~����v<���F���QV��YK���Vpx\vh|圯�sn:�aV��Vqj���z���֞z�G@�˹�"��Y��ӯ�����Q���I]q�N�_s��w�5�>9@����cE��6`�D��#Y��ሇx�vdJ��\��AU0�4d\�8:]�h�k�I)���g��l\�C�
n��¸��`�]���Mg�� >��6َV�Z1ת@A�b始$N����}W��1�l����i��&QGN�8��C��Z&wM�����F�D�7�C(�}+����ʫ���2OH�D��=<]m�w��f��f�U5)�j�o��^xJX-���J6<�����\#S�l(���z�\6�/�Y�n�Eq��L�1;F d�)E� e�;�u��U����P�~�ꘊ}XԆD���^���z�
"�2��7�8Y�K̓4d'�6v��j�m��nO^��|J�+)��5�kj�xK��x�[;e���X�*��JB~�3i�>�kOJ�P���������`����
۵+ysL�L���$����U��D�.c��f1
�	c��;��|�d���GWm7#b��w0j�_-��=�϶�e��y�J��=(�Ш�5Ѧ������X怰�g�?oL��r$�2�Oa�e�`��P��2k�D�� ��ɇ�o@{B�>�:{(� �h��U��j���j7%�¶q����t�����G�}0�xn������K�]ACis�G!~�'e�s6��G[Q{�h:�_c��3�
�v��Wn�y�~B)n3�8B��Fs�7�
b�Ҧ$�&s�va�W���c�˘��][��=�D�a�}�f�r�X�9[��!�X��W�Z%*�f[|�K��I8�%T���Dd#�Yuw�����u>N�=o8@3�Ƣ���]�ţ$�CYn4܃��t�+@d����ux/٧-Ч`��KT�d����v7��d0m�!73�3#aU���C�(W�Q����e���*�a3�I��S�}�F��7��V*E헝"�zy?A�c0�b6YL<��5u��GN��.^Y֩�k�	)6�F��&�Nr��sYt,D�8�aQ[T��7���O��;f��DK���g)���q��&2�Y���sf��@���H�S[��Cx$B�o6�LP5 9�q9qa�wɜ�R���r��.��.�.o�w:R7{8��	�'h��`څ�8����9�8؛�:E�AT�	#9�y4�m���о�n]��9�ь2+M��VK�������#�C-oτb��X觶�Ɯ����aYy^ؙni��&+a���cZ��-�[���5�d%�쉨��*�M<U� �Z���EA}o��KXj0��E�+��o�S����)�Q�n9<�&J��WG���*^��c�Zc�f'7�y�����S�Z�n뎻\Q�om^�sR��A!0��T�Q��-@�M�Y$}>���CS��43�,�۰��f�\NV��3�56��$.*N�݇ӫYJ��;7�T4���ta��L`�n�������+�Qm\H��4,�aP�rd�}��-E�o^pJFh��_��L+�OH��=�f#��[Ƹ�&���^�M6��Y҄8��S�]߶2�'�<t��Φ��=�3r5z��8�:��G���rpa�4�ܳ��r�e}���9J֒i�tc^Bu�EG��JU�zL�8{�C�PJ�U�d��(H�w�h���>m��&���w���񫘌]���]:��&�T���QP�ِ���p�n]h���c9�?0T�<z�&m;��-��}�0�����f�0C&�j��Lg�S�Y^�0�T6L�׈��>s3_s��/�J��W�����Rn���x�
�2*Y�HS�!��i3S�,�\�>iy{�&�i
��T,�rU�iE'��8#���Z'�/�Mњ\��=�ռ��`
���nr�WC�L��'p֣�O���O����߮3��_�J�("q���u��#�*�Z[)�7c�!l�rc��"�L�9/���kW=1k��+�+�9�v;�&4H��`��F�E��/z�i����o_{5��,���j\�������|�d���u�2��ƣ>����W�&�l\c��$s�V���z����Oqpb�{�G'J�D#}.7/�֋v=�L��ٍ��R{B˗�dތ�R�=Ƶ���L#5�x����[	%N����c�3�:km�K�l/e'�G��E�F2aU2v�1g.���3���w|~�t��~��zHp�) -�G���g�{���W���?�U�Um_]K�O�8Ь��_E0��'�+en�K���+����	��M�3D�N��l޽[M�-;bj�k����&���|����R���T�j�n�5���K��w҅:{�HK��'��D���4c��.�>�Z�
�/0m=�O^�"�cV\P!&.�x*�6I���Ǳ�����A��e�}Gv�7/�G[��i��j��Ƕ�N��ω��hٹO���0�a���Ff	zj&���o����Fq�sv;������\�S'[��,�{S��4�!�Jl5c�f�b2��E��3�9��3�H���-���E�a�Zh�qm2$�m���6� �C�n��v���8#�74��f>,�����l�r̵�K����O�kN���0+Փ���^���\�e&��JZ�qtѕw�f�=��`8�
�2�=	=�dRG�V�U8v�
�3����c��d�0:�nP[U�a���#t��o��Z�i\�==��NZB���!1-�p�
n�hg��[J�8�r]Ĉd�&U��-�ج*:�H����ģ�ݕ�D��^��;u�����Rh+.����)�S�bSx5�smQ����68�����ˑ���F���MS�%�I�/r�b��W�ESP�c����&'�5E�,��u�R���	� �/_A#)v��3���j���e��ll5m��-;�3x�I+j�&�M�Ƨ{��VE5lǻ�Y{��=t֮�irwu�-��/f��c����^8�֭�����rX�W��D�+���1������g�9kB*"��Z��)�V9�Kv�߮����EV��QJ�T-�sRks�Qj�+b�KS��X��Q�m+YYU�6��sNr�-5���P8�ƩY\عw9ǖpƎ���Z�ͺ��o0^r�ه�Q2Vƃb��7h��2Q/.�T�3��R���G���mb�ҭ��V'bѥ�L���	�F*��մ���s^]�m�B�ю�+jZ�m��]u��xcd�ە�ʲ���&mm�s�7.�[�m�9s�K8�
p�026���
XNva�����nvt�Uu��A�e"�	H;^qRl�9�茁�|^G�,gy�y��*��[N����r�"ػ�yok�r-��{��z���_�}^�e���0��O�������-�բ�٫KCJ����B�}�o�|����-{��Ty+s�� �`F`p�.����?x���>��^���E���_mz��V�'��(fG��4ƅ>��)㎼Atc�����*���V��e��&�mZw.o}�k�;1q�����pcc+V�3�9�2ֻ�����9{����_�o�:(��ϲV
�F��Ғ�e᭴R�E���E7W�[�i���Jr�Vr��T�B=�9rN�f�%8)i-���~��yz7��{�q�8e�A��"w�P��ϭ��{Z�f��fx}=g��k���:��o]w�<�x1�Fu��iA� �d�͟n'��ݚ<����܋����6�����o|�{����c`l�U��&�4���,Z�>���bV�R���A�>[%﮾ds��ì���uoôN��f���G�Pdk�z�*!���Ɏ�cܮA��X�4np/���T�k��[�u���=?!�M��-�)i�^|���np%$�>�{1#�l��Hd�ӌB�m��-�{=�/�j�ǖҴ7�˝�V��e:Ks9\@)8�e4�{���\#;C������3A�<}�_cOpW�b/!T�L�������;r;�%�b��m^IW�F���]'��g��d0��;�))��#�	s��E��Dy��Ze�P�ݟi�y�s��F��By|�?{�!ؖ�?+F>ƙ>`�6$������K�
u^�=�yw�����)1\�����o��X���ܸ}Q�����9Cձ%_�}j*/�=��f���D�,�-���~d��f<�����싡�:h	�c��0�Vm:��
h]h\0��P�,�l7����Yhdzoi��"��C:��ۨ�b�Gb;�Q���7Q�S�sЭ�M7�������s��f�\�w���gq�-f���բ|ϔ��=wQ�󡟕��=��}��c5��ꙃ4z�g�����X����*u�=vT^�]���C&=���;����ˢx/d��.$�o��w�]��н������XP6I�FB��a��h;�߼��f�U��@GE�?��s���k�i���Ж4�������\�}��/���T��l��%�õƀ�1��A̅�+h�iu���6|�s5�ʾ��
_Z��ƺ�S�q�1E��<�	q�0ِ�Z=����
hZ1,�<q8{�d�Y}�`o�4걑�Q���Y��rL�y�/��ظ6��neAï��G�C�N�2�����]M�y�rC+v;Ի��H}����]},_ԥ�P%,Cb2���,��H������.1��Ѝ4��� ��V�P��^�&�.�d�M*isЄ��%m��%��.3��/1f�����SH���*h'��V���w9~��y>���0���ʃ�J�[iKǭsI#]����H�6�6��
e�)�i���^���<���swb�-4��хANؕ4KA�Kmb-��Iy�q�� 8�0T�6KIK
g#}�W=�ʱ#z�h<�[H��
َ�A��Z�tM!q�и�v!&�<�W=z�:����3.�m�Ѝ��(i/8aM ��)��,�4��A�%--� �me@��l�Sg3��c��^�ˌ:��CH�ED	u�c��ZH�ҷm!��%�/�"���4#���S�zg^D��E�q�iX�a�lE4��4� ��
b�A� ,��pĩ��1��@K�b%�z;u��k9~�%�q�~�K[bJ�\aM%l)��h����p%mhR�l��1�)�7֐��L�_rg���L�ĉ-
�P#M"��H�Ĕ��n���5�K�*if��I��*�oﷸ9�w�Pq�~��@���4�6�S��#!�Qk92�{�u��oco/�f�}AC��(q����v��z���7=]���ݰ��	�H� �Z50����a�4�i1q�b]bס$E@�K09^TT�w��J����
�F��� ߠ���`�h��7����#bV�K1hj#�黽�s��󴖞ؔ�h\h0�i��cH�hR�98��F�	�h�
�J��l��h���s�����w.f�6ď4��n�K����
`�� ��f4*b��H�H��З[F�F��W_"{�y�W�1�y��8Ĭh6Ҷ��4$k��bR�+�*v�6 �1������b�����Ejߢ���Si��D1-0��,��4��1(�I[Kp+p�4n���B�Iq��i!�O&bk2��1�X��1L$S��R���;���B�,K������M�u�7	km�ɏ^>r/~��0������
b���6��÷4u��L?D$���m/0�I��<��.�4d4.5}���X�����:�;�%�m1KE�[iҶ�d<�u�a��J��j�y�����8�C,�摨��IG GXK�M �CJ��0ǌA���4�`�pc�,߶�KΖ�?�/�Q��;���ԫ_4r�0��c�#������_o��b��B����f��
�+)Л/rvd� +���BI�X�iDFʘ��1~X4cIq��$�9
�C�&Щ�m%�/3�	i�6��m!��%�J]��+;~�đsvĭ�M4+tк֚�a#��HR�� �D�PBLѐ�i+k�ru-���]�$C�!�\�����l�B^e�*|`�S��Ii6�����-���+z��U	KK��B; ��$q�k�������ј�SĀhZ`��4�i��:9�Ȼ�+=5�(`�B�K�L�Bƃ��cI[
b�� ���K�!��CaLE5�M+��y\���(1VBХ��\r��,bVצ�0��%,8T�\�bP�0ƒ6���b&+�}�����KCaL-�6�n`H�@�>03P��)�KH���W6�`����o��w=y�y�C%�Ќ�A�h�-�*imvt�T oЅփQ��۶[I�f0R�gu�Ƿ��;�Mq͂���{�-0���
X��-�1[BVҗm%M/4��U�+}h7�c �9ewy˙�з0K6�L��S�`A��H6ֻ
��=�V�q�z�$i��1)f�|ﾽ���2�[�3��E,����KUT���)�״�"�
�w�=y�)?+�R�h��M��H����i2�:�g5!F��FI
�BKe/�ퟢ&b.D��3��H�
i��@a�#ga�ѹ��k���5�u�[�.4�O�^�'y\�n}����	6��G�#�
Z�S<ĵ�h-��$K@٣p�֊h�����һ�.oGv��\�`ؗJ�X�Ǝ2+aLJ�<�ٗ-�kp�hA��1[H� Am^�Ǧ�?4��aP��1+~bJ�.0�ۀ�^���u���G�wTVyn�N�T�uE�Em/*񢷴��}W��Oh�x���O�բK�:�f���5�a��e���⧑� t��2��vTo�ϡ%$F:�MY�Ɔ^�����9�W�Y�B�`v���V�ÌY����6C��U�o:�f\�^��u�V�y`�6��>�oMy�~���e�gfD�\�zћtN8ok�{��#��<,(l��/���r��y*Q1=Вr�a1�=N/����|+�����0��W�3n�ܔ7Y+1G9b����`�$sh�`!��w"���:�k0�!c�>cB�z=b���̀5{w�e�y\"��R%��x�2{�/�˾��C� F<1��-^�d�l^���Z�l�Y����ѝd�s�\����e��D8�q�H��X���=�b�$�vqʛ:_�n����|�����9�-�����N�_�3d�#��H�\u�r��<���Q�el�#9��m���r��eQ�/m�4�i�r~��Y��x�N��W����.�.Y�m�i�9��i ����S�����Oߢ*M�\���M4���U���C�֌�����V]0��W.�{;{��V{���k^�V�=�l��a�}�+9�Q#eyz	�W��/�B�/����9��+�2SxK��(�~�o �����L��F�Π�Q a>��"X��ú��\f�UTe���8r'a�Hjm��j�M�\R�&#n�}� ��W[�I���������_$�1*SN:�ꏾ���;�^̰�>���GV,?�T7�5Ӥ/+6�9Fz��w7+Fu��P�i�ڱ��;N˜�أ�P�\�L�쒗K��͎�����9萣��"��܇j쉆o�cꬩ�}ƶ]2qvre�FvK�*���4o%mV`*�����{��UY���7�eH�^�&]nDZ����)���v����������fѻW �uL��!ҥ�`Z-�9y2T��˷J��1*�Q|� �n�zl-%��V9�,G��5'�wk;Z��]NJ�Vdm.63QR�aY�ӊ��x:���`��u_72��7{�d�!q%ڞ]r�l\hY=٤Z�zn!�X����BY��jua�l���5c.g����)��Tb$��q���\�	]�u��Yl�f:El0Z>�`�'�����j�����q���N�ERfˤ`) ���,�l�Љ��HĹ�fH�.sqL��)�%a���6����P���SH:!��v��϶�z�ot苌��M�g�H`�ҚӘ�v��7��t�`�b�M�hgJ���"�IT�-|�v!�Z��5$���E7��/D6�g�kgS,+Ww���+N_�;���P�7�n�t����]�r���H�DW����w$;1��˲ɤ�ݔ6�� �fJæa�sI���
RWr��5���=��ׯ2ֽ.*ς:�
F�<�9!
{2$�{��n�+y����
orI+j�-�ڐ��4�V�{����Msm,�qq��Q�Z�-Τ�'k;t�9+����O�������u�L����^T��E�QD�%H@_�Wb�&�N���)w�sq墴Ᲊ�4�M|AQ1
(���%�Ջٶ�<-���1�9͹���j�8W�a�f�]��mV��9c�^UEQ]��+�Zla9J"�����&s5�G[���Y�׎9v��2�Z�(��E�<�sZ1��i���w�ܼ^<�R��皼�5-e*V���m*�Ux���EFkc�UNR���ET�٩N<�Q�y�#S�]K^mĠĥ�
�sc`�։��n�S9Z���[�rU���kd�ռtN2���d������7���[!��;#�#����Q�ke	���cn��)/x���+�����	��r[��n��z���O}P}�m�@���ҳ�k�ӗ��8E�%���p��iM�|�z󮌃�P�f��x��}I���:��?43�C����7�qfX�$������{d��\:��՜i@���4�ymcl�Ǖ�[ںX����Z7�FE&õ�G�7�VYܓ;�9M堧�����Co�ʚ�C1�n�"�N�Spa��:�u�ʼљ��Պf��\X.}����J�Z���t�[�qۻ�vȑ�n�� ����JC��}g;'��ثK���p��t�{m��N��7?��n�c�x�����(1�UL��ӳY�U��nTY���
�D(ρ�:$����wxT��v�j�Ň�1�Xu-;�oS7��{�����qc�(�)&k�����Ic�
�m��T>Y�"��|g����@������Ud\�u�Mi��n�9�ү��_&��;��h �'ei;/w%H��,�l_=����g�(r��|̓HZi�W�3�uo����5�_{�Q+'��V�I�[�a͠�]�R���f����g�����|�f����1_�w�>����o�α��Z�ț���%3K4�Rl�����
���>���#�m/?&'�mL$���w}�]r9uw�_e�ã�G�(�z�ۊ���ҧa9� �5
cvcB���eXLJ�h��V�t������!.�]��fD��¨1����2a���A֎���;�(F"�p5�`��3���6�l��[RN�}����%����^^�\H(�V�����)|�pefչ��}���\-ZXą#m���qVCո�N^8�S���i��/F}&Z�oJ=;9���M���5P코���\=Z���<p��z���[(�[|8�^dBf��"WmΚ�f䃺''���~\G�3DG��K����o���x�����qu#=�!�Q�__(�u	��9HK����ޞe,��.��u�حO|�txm` �$��V���s�G��U��ȝ���{��*���/(>śQq�{v�3���� �<:&	rwV�S��j�m!�咈�2醠t쯉�9�nV������t���J�"��tfi�˪��dkf�M���07����J+�uW�ٙ��5��9{�mk��BGi���Z��mګ��9��q�l��Y�ʻCGh(\h���CjnqE�^�;Bf����쎹��;�_$|�m ]���0�����5h��Y7���"��M�8k"k��� �2�*L��m�� �rmm�
�/~���42vM��������}�m�bWjm���`�IO��-�3��V��hڴ���˷�p}�7Cbx]*��W���Y�TK$�Ro�5"9��q��SI�=�I�ޮ��I_�e/?;�������Ϛk�NM`�����)p�rQYAߧmt�,�U"+�¹/)c(g��1t�jzg�I0��A�Jw}[��W���in'c�U㸔m�.Z+.�.�rCH��ՙ�ճ�$�E�O�k�hM����]a��}��u�G��r=$ъ�|�\_�wa�
j�S���@�<njpkL*1�8WZ��ƶ�䝡=7��~6�{B%A2�ga�;�9�G����x|���Q��u�h�q�6��n�Wގ�ɾ�l�x}k=�����V����*��u"��A�!f���T^Y�1�u�9(V�����[u��D,��sǛ�+O��\��rU��'\:s�m��{�0Kގus�J�\5��5�<+��9Z�����Fʙ�ʹ��Zm6�"����S�n�*�*�9L��ާ����+�DG��>��">��^o�x��n�)�S{f���w�[��X	�.	D>��3YqE|�%�O0����[AN����-�	ݭ�X���00��<}P�!��N
=��e�8Kt�O�w~���m��*u�qRn񂊉w1�~� �Rs�]� �/�=���+2�x����F�(�ޑvcJ)�tp��S�u
�ex"��E\d7�zn���Ýo]G�|(���7��}��DƠ�X�#	f4'����!T���;���<����Q"홻�h�V�Z<�����{�x�����n��fJLm�b\�=Ηeo78v�xz)?j��I&�HE��e��Ͼ=0:��蹟o[ș��'��E�-&�3ޓZ{�q3YX��N���m��S����Ź���h���K��CöQ�,t�#��#R����F�=��lf0�{|"��N��0�'c���yY�3�E�c�|"�lg7��`�UBN���Z�y��g��b
�Cޘ��e��~���̪�ߏR,,�U���_�/=c�Q�-v�����nh��%�ol��p9]2v��b�z��|v�:�����E�q���s��&��W:��U�R����	��s�n�*i�۔��Z�)bR����n�(Z$Oq�2\-I'�G�$6�	N[�����Oe����kS$ў銈hK��Ԓ(.ɭɜ/~[ÔQ��,���o�N�8!�C�j��d��}w���n�����34.k��EI
ZHpB���q7hհ���eu�|J*���6%X̼��ȓ�e���p0�ǜ\7g�dV��P�ݘˊ��-���]���5rK�%+R�N��Et�٭#�����x��v���+��pgVФ��*��Eth\W[YNz��#�lL9�q��3(�|yR~���/���g�ШS�l{����,�u��u��rܗ4�����r�����}_~�W�]��W�|��}�D�~�����>�U0��;�Жu2�=�,�3�Rs�u���ك	;�)��/�ڄ���Y6닧���
_�(k�75��$�h��0y�uPڭD�u�eh���$l�<��$�{Q섈)�(ϵvD�p��daweu򦬺�(��5MP�f�mckS�CF�|P��q�L(&p13V!=|D�z��B��f��T��ֲ�L{d��=�ޞ��K��y����~�A��������j��cn�o�ã�Ɔ�Wɚ�M#*�7V��I���X�7i����������(P5&�V���3{bi�	�n�ɹQE7]�C.���xA&�F%�;�?W���g'��Σ�T��{��ٛ���ԡ<VT�Ko;Z�r.lt�k�tX�,���T�B�z�8�p���Gm����qjdosr��c��lX��__���
�}R��L���j�E,�o����IZ����m���2�h�v�s��'z�u��R2��R��iS Ey�tQ������e9��X�W�%����Hٚ�"��3�u/.E8��R�Y�uR�����s`�9�/��߉ܻЈ}R%��l���I��Vj-/�g
6���Z01�R���R���r�o�'�yr��+�_�J�$�(���f'�J<��J�����Ej���p^�ù��Gwb�V��������#RV�UḷO�;��creޞr��j�R�u�믳76&�|���(l4����.�_}u�Ĺ���(�Mm&�^���M6w�l��TD���=Uiɺ:�w��0ElUw��K�r۸���2���V���XZg>���mH\��:{�j�ٰ3cbrf8�/^^�.��>jU�5ؔ`]�TP��.h�ya����}���Y.v��s�ݰ�av�����S]!9��V�d}�:0�}����S]u�	On떪8�	{+���i�E��k�WU��2Y��Z&U�Tgfkw5ml��G1e�ޖ��T:lE� �{���V?�Y����V��3J[mZ�)���R�9i�����5ǫ���D�S�V�_0�*!��)�҉d�wm���U:�*[���^2���&-Q9�mZ��.2�ܷR�M��י�LѼ���j[m�J�s�Q��J�N3+Ûxr��x�/-1/���-������;^.�(�R���.Y�a(�ȸeJ<Lm�]Kh�U-�n��s[^k2�9Ɯ��r�]����8��F��YF��-���;gQV��q(��]s2a8�C��߷�_^qʣN��o��a�K�[�֔��N�1@YnO���˯����ﾊI��zz���P߅]��~��#�us�ڻ��,J�*���읠y��G$�|���b�C$+ٵ���묎�f����+�36���&�n�,����s�F�y��A��Ƽ�N���F>�2�v�ܓ%n�!�7�6C8W���&P�x���vϳ��w�J���t�r�6\OW$�q��b��-f�Q�Daz/!���1��H1����hն�wF�
�fs,�Ե0����>�T�}�>�	����;87�8M/:�X2����M)r��/3Ie	r�{0>\��-rokre��]\gf���8��;��>���ި����UW�K��G�?{S���|z�'cfT3�Jf4k�Q#�m$WQ�萝UEU��[[5xC+6��Tf'{�ս�Ks�`|PQ�o5ݣn����<Q�mh�����5Ό��uvXӶL\�7�8���K9�5��]��9�qʳP.��r�X���h�(r\!"���V&��H�a�3�Uf�i,g��|�(��}��,|� *�Q�R�V�{s�w�-��7�oF򚷒�q�N�8�p<h�#:U�t�cw�ӟ��F��*�#�j��2Қp���X�֣�6jm��=�l���O'��� +2�n�?�y��z�k�H+����{%��ĥ@�~u��]���of�␦���E�h�\����hrYuȈ���'��Gm#glg�t[�L�\e�5�sy�{n(j:��l;J������G�z=��aV�fG~x��x�� �]�.��7�hA;P�/y�ũ&6J ��N�ȃ"+J9`�U'��b�����&�6���́�ֺ��
iJ0��F�ֽ(�X�s�����;�PsN�݈b�[
����+��:u����Xj�Or��Wv딈d�┼���h'��mǵ5��j�Z���| >hI�$ V�y/�+��'#�
9g�}�(��� ·z��U��\�.*��<��#W%l�W�$
5�ǅ���tv����d�S~���z��=^�ҕ��m~�����a|{�̆����Z���Ār�(EF����U�Je�������ACWgz.W��c�I<J��g���)�S�h��RM�Qlb%U���E~�Y�2<g2��N���$��$��9�K�k� ������X��R�˛���#�xBr��c��v��H5d�.&��Uu��k3j߃�����q�҅w]�-�7w)�z&�,J�Vv� �UN���M=�w���|�0bHW���~[���}7]]��o��vr�b��[~�z=6�מ�>ނ�	��	a�[R�(������������D-�S;�\V��~5�h������	t�G�m� ��3$�ud��,:�f��
�Y�jt]<:���Ao�\��S͸1�4E�WB[uUvOG~0q�q�WT2Q� �52�A�T��X���k��lv�w!2���帾W�6x<Z/��FE7o7rkn��5�p��2���]��뻬�˲Tyj&��89J �r��Ud���{���X�+QC���M������>bI6�$˼��٭}�QGׯ]�$�_�O�$��*�V�-�+���c��P~��4��c+!b��j"�Y/�B��Ĵ"�/����H�ؘ<`�'T������z�e$�uЏ�;�*3�GOsU{�1���V�Q��.{�M6n����0q���"��5lr24�����qB�����!�=5k�S/�tM]�������"��3�7�^�������z�Exo��,�=�?/}����T�9�(�d �r;2�$�������,�wj�d5�La�� p���ڳ���Vs�V��N�F���:�ʙ��!|�!��B:����x��`��}w��:����q�����'���MYH���T�[Zhu�5P��@��qڒz±s���[(�4�r�7�i��Z�lmn��.�9�5��P5"�ѵ�U�NQ�ID�z�9��m��G�N�\�e�3?X������2�cV���oq��<0���|cu����v}�鵬l�$���^��>U�t��S�=�N��]{=t�)-��g|�;���VK�����v
�32�dh1na޻�)��^�Ik'j�u-�3e;7Y8�j1�=��N�.�{�>����|���_�a���j�_�bc��j���l��ڇ�A9X߫��?U��U��\���:*0Ok�U�#~�n�^q5@(w،�EO;I�y��b�<~�j�f�iu�;<�����0X{�^^��֕��!���޸�=���`��
��ڱ]Fd���t��{'���|GE��E�$v�8&="R�z>�|�������u��n���Q7��!E���7�泫��w����j�c�a�&=���D�8���ҽ��_�.��I��7�5m���"T��x=�w��Ö�dc/ު�����G�8%�z3��-�l�ZN�cQF�����]���{�z���M|�_0hI
﷕��3��>��z���<^�>�9�4Q�6���Xw��mfj�5 �a�Zx�	�w���E���V�,���॒��~/��#�XHB����y�.'F�{��^^��x1D�r�	z�)���L�U1%�݃�n��]�9b���u�,��oNR�Q����nv{�+�z'iƙ�N�3�������{KS�ޭ��fɚ}��;��x�z�H���K�)J�k�7�{����b���`��] �M�?z�7x{y���}�D_��T51�ፑ"{X�B��!�f�f���<=ώ�@֭!����C��c��w��w޸F:M�	�k����[%C�!Ƒ���f��Ρg��+�7e������]�
���Z���l�2N��曟���~��_6�!]�.�1�gǹ����sQqtū=�0;W�rt�e^���LU
=����(p�'�⸎ iכ��z��̞�o���%�9��_���<h�X#9"T����p6���V��2X�H���>��Z�,q�ۣp,��X�ǋ�,,{�a�N�`���a^������MgI#9#��^�`���tr�$���H;�|(]l
��_��Na�}U��{O��m�'�cM}��l���E�kQ#w_��z?uee^u#چiB���E��]�>`*���m���i@�ʍ�ʳ_?�}��'��O��`���� ��2���2�O��u��}xl�6b�ה�N6r�9�,{|���|�Y�7��ǚ�ޡ{\)	�`��|P�N�Ȋ=d��Ů����1ifli���Dc,�{�B$���أ�۩�w�e!7��&����g�Եaʩ�5Ȯ���kpa�:E0�uq, 
R�%�C���9�^�H��Z�Z9:���a����;����'ǣile���'��V  �x���G��7�Q�!�O�>���Dغ`���뽚�iZw^e��CNq�#��P
�]b}}�����}���@�\�sݮ�I#y��6~Ԝ�(2���=rj�U�,㕋2uM���.�D٠z����Knc!������$����9��<wzVWW�Ua��
ݦ�A$�[���_�U�1����K�zTJ�5֩��}��'.�bjV�2uV�RvY�'�:|�p]�L�����+�eu�n(n#�*nX1m(��-̬�^� �
�z���5��CC�w��\qY�Z�V�Ǝ�u�*|n����)6fTB��<�:����b&U�@V�j�����s�w3�{�&��+�*�n�.^og�Sj�j�l�������D0��Al_�{�����2����7z�B���d��!�ucz{�sӟ;�i�V�y}F�#.�2]Ý�e���G�3�Itu�'�;�Rv5	PL���p���`V�6��ݧԤ���@fZ��jv��ux$YY%7J;�HTj�-{�Z�W3����|��_^n}n�-�Զ�2�ܶ�"�w��n�J�=R��⨹�֖v���b����D���J�C1eee-�d�*V���Z�\=�f��B�Mk)v�0��d���gyEȌZ�f���<�xQUh���Q-�,-��1mu�L&�����r�D�&���]�qZVVWl�\�R)2g%���enU˩U�Y�]1�cR��n�c.6+v�DT2g�6��h�gL�2�5(��F(�Qu���2�W!�]J��(Q�i������ �w�7�ɲf��B�Z�!�^�,]�e7�n����	ؐS7��a�/Z����lk�H/y
��yP#O>S'�R-�waã�a$i�}'���CY/P����GLV��CeD��*s����q��@�)x�U�p�wK�ػ9�vw;8t�{�0��6}���m(����O!N�h{�ܻ�$k����_��N�	��� B�>,$+օ������_�":�r����a�C�ܾ����c�5[���(��0�:b�+�9v�Z���}t��wQ4�ل�z��\\Vp<l#-qSO4z�%��n]���v� ��ŀ����֒|~�Q��2���޿z����<E!��$�����$t�~b|����q�Ig=u�j��G멞[��œٮ�>,� �%����T�Kڰ�`u
�wd.���5¹[~���Ts�3U�K� DS���=�1ߍ�ɓ;�dB��5U&:����%�1֜�)����hp�S#��1�qٮ́|F,6I�;dw^����7���\B��6���6��,�~W��N���	=7��d����z��B\���J\Ԓ4��W�E�9��� ]+�T����Q^!-�>�mG�L�܃�<G�o�u-C٬ �ʈs�RE���]M>�%ΚSxB��2׉!;4�V��[�=�~����R⏫�c�Ic_���c��j��&��m^o�݈��N�5��C�}�.�ێ�~�7/�
�a%��O;����!����lq�2��>?���^/yf��gM�rel��l�MR�W7@ĺ��NX�No��ʀ�7`�R��T���)NxOA.�N�u�pբgs�Br�qn��PzD���������������{�l��v#����n�iӚ�<]+;&�i4{��:�O0���q��E�$f�91�R�GG뼙[^�Ϭ���C6|�ʨ�0�"�t�����:��S<h�ڂj�K��*�P��Ar�7�75��v/{٣h�Q�6}�8��0��jtѠ�%ﲔ���$�Ci�H6�x���B�ޛ��1
�9�'��/ۄx���F��A��hv�#a7�_����w�j��,���$�[�H�@�t�l���5Jqn<�b��7.��)��Q^R�yܚ]/಼߇;��{aK�8�ܴ�i��Ƹ&I�����t�W��R���.����O��:-	���[z��;*J�rTk���ܒƳ���`��P�֤�'N��g6�R^��� |�����eg�������ikp濠<t�<h�I�_UY8t���gu�/Z"��?���_�l���I���qT4�o�x�.Рl�ZB�i�#}�+�'h�e����C��n�:I���H�����q�Lsw���2�p<Z=���P�6�?Y�z��ё.ǭ�8X$+�0����{\k�C��3ʾV��{������ղ	k��ϯ���8��6z��`�#8Gu��|��+���3~T)�zq�^/�x�g�"}��W^��X��`�"����q��X��˛�<�����
�6b�-�����_bLCl/�s ��wm*n��Dš�0S�`'��m6;g�N��U�X΢��V��M$�7'6��m\��NE�\3DݧZ��4ވ�ɺ�m=�L��'?~��n����� �����~&��quQ�j�������L)��3uF�({ܟ���
�7#�������"E�z��wj;��Ɨ�}kM��i�<tѲ�#XB��E��u�]W{�B���2���iN_x��;ю�v%֡hZ5��C֣W<�i�&�h�A8�Z�>Y�*Ab:�]������F��+Hi���I�q�Q9��J,,�}\���ؘ�J���31Y�O�T��\���Z0s%�f������W,S�e�K|-���P^%#`�2��=�):y��u}Y���P�@EV?�l§^����\���12/�,�cǈ��<g�w��X�*�K=�RU��g$�G���7*,���NU�@vKs�b͜��+�yѱGe����5(�Ӝ;����?k謹n�M�.��.�������#pu�Qo__�B���������>P}�
Ww�Bϒ��Ƣ���W��n���v�����o���bA�ik�Mi3n�zy� ��r�쌘ً��;1��I9������0?Jd޺�U�Lp����}�h#�:I��T��ޒ��߆v6	��>4��-���a�b�b����ܿz�3���z��~��BiLoW���Y0f=�}u��j�T|Gj$�c�.�XcUKvy���Uw�=��4�"�� �'֑t���8��|��1J����;}�<��H��V�h^Ե_���)��ۼ^�Q(�S�b\��Ի�kڏ�=�O�Lw^���ڻ���8����6v�\�L�̻���R��qA�n-W�U�������u�zf��#�$6���U����u��	�/��\Y�̠�kDd��HS0�>N��ƈ��OP�~(�^a�i'�F1�U�����8I�;� 많Y�*�/�G��-%eN���/�h���V]��)���ۦ0�!j�7�=�L��z�X�y'�<N**��q�<ǋ�gz��U���x`"��#�������ÏH9a�dOB�~y���_@n��wX7��	Ŗ�q�}2�z�&�q�{�x�>.�j�E�C�8��ԭ���D(���>^>�8��+�MC��9\G����bu��Z&��Y�H��p�{e��r�֚ߍ?6=��y��{~�=)�'MLQ��V�f骓%z��D�v~9m��%w�[v�ε��;�h����Ơ\�j�dE�t�������뿒\�����53�^�Z����ƴ�\T~5UFMá0�9��"���b��,�D{Pt�'�q$m��<t�<�n]��t�4#�t���A_!�_�F�6������,���E�h�@��>l*)����-H�������7��ވ~�#�N�ƈ�H�3�)��;۳�q"!���W)�\�8A���w�R�>���{�K B<a�V����O�l�ȅ�=�G����w��b��Q��㤚?lM!�<��Lא㵜UT^�����|�����k�5����߯�uy�E���ֆ�l�H�����0�"5<��'0r�ݾW�1W�. \�:����:J�Q�2�#E�����WHmNrQZ�ժ�n�G[��E�gCӴ��fqjm7?)1b��eedlm�����8�5���p�����Vo�/]�I8���کq��־{2Ǯ8�}����1�����Һ�۝�����Ymy�Ha����S=8��Phk�KU8b���W3=�ff wsuQS4����|���Af��H!KR8ig|���e���W���a䆸���_.Ck[?dY�vA�����ܞ��A���-/�C��G�N,�1,#�<V���n�{��>�d�㜆�M>_S��ˏE��7��=�ٻH'�w�y�Mx�\EJb�=.�<��*�����v���_q�T^!đ�����D�M�C��{��A2mͳ�ݝ�UaQ�cI)�s�k���p`�������fۻ�++��	ǻ��L�.=�j�;ݤ�պ����U~?�����e�H�+G\��sSƵmcĐ�◍��pR��{�����k�y��FZ$>YH����B��[{�~����>�r��k'OТ��G�pF��U��D�r���#a�<�B�6a�B���?Y��3{���,Cf��K�1-�<p�\��B�MW�y�e�6b�d�a�n:fVz�rfc��7NrzDNJ��O�a������ml�bjA�(��Ɩ<:Ц��	�6t۫��b㙬YB����$��,�H����v��g�<TB���x���A�:I�"˿X'2������s���R�=k�����q�V]�����<l׽��}1��vN��GB��f�Ut�E'kZ��;(��Э�L��M���̬'�������i���Ǖ/"�
�9e7���d4h_��wyn���8�%z��W@�)(B���tЪ5��*�:�F��H����r`��6�->�&��%V�ŧg7�.���u^j7�/&D�@��	ّ�F�3�c��z���t�⥺`�T�:@H#9�h��X�{PM�Q\7�h��AVv�_�P�+X]��T}�����2mR�a�*��i¸v�,=���sz���Y�-��^��!G0�[1���2��F�^�q���F휰��X4kl'���Y�Eg-z{�u|��J�BS����a���l�sL��3WB�U���XH�%����/�G�1�A� =mA�V~n�*L��B�ި7G�Z��&GN���oe�9�}����mZ��-�6�	7!6�f���wԥ��$
�Q�3���r�EKIy�����o�A�����x��;�tJ
桢���c�i�$�*���r�;9L�
��3��ܵe�\��J<F��yk��<�<$�30nW|B�sC�F���V��Ve�v�,;��Oz���1�u|��D.����R�����1�FD�^v��ł�tCVj���hK}�����C̺����E�)�e���ì�E��i�к�{.��S�L�1��:\2)��U�;w-C�1�M�a�$S+.˃K.Q�r�=+��"����۾�>G��7�
W9�h�h5�r벊�O���q�m�U-�҉uζ�L!u���-��Ҷ�9֧7]u�J�EES�P���[m
�V�#�B�L�f�m�9��뮺鶬0RՕ���Y��̊�f� ��Fa�+�Muf��죶(ˮ˚PL�eV"FZԤ�f�f*lm]k*Q�m]kW��5��G0���݌�)�)�.�s�Kuu�WQJ�m��[m���[.�ˌ�ɑ��Xerݳ��5*Wj5�T3mDYE�,+R�WV�ڎƃm��2)��Du�����ʫ+��Bz�8��4�z�d6��Sw��ڨ�����L�����4�+����{ޕ֒��Fs;�_��O�1��}ͫ�j��̚���Cŏ!�</�!�V�@n\�'K��=�6�s��#�yQ�,�kf�j��rGcx`ȃ��\�Lw/��[DY�69��
���~�=U�oe6q!�D�#O�k�лTX��ts4z�:��T�­"�1�:p����Ej�,[��ro�ݛ�%�#�_aZ�����Q����xj��A��_�z:I����s�מ�(� %"5�6�5U�ݭ���I�[ȑƎ��\CJuܮ�\�l���ԳOj�K��P���EO��<v��5���q�=�������#���ȑ�ׅ������ V�-mB��������)-.��"4I�v�U|��;s��R�ÜC��d�8�Ǉ��2D���������K<<��{1�Q���Le�P���I��vl
�e�8���Z/�j�l3��
�Ø�s��ʯ��t��S�яە�ww�>#��Q�8�����p��Z�8��Ow��l�g����$�(h"��E��s�P�Y��}��p�b�?��črH?x��=���u����3�o0�g���լ!H�}k�#uJ�PL�y��R�g�d]F�����1�?'F��k5�[�Q��Hu~
߭��c-3E�9d����7�h�u/���xxz��K&��_��>�O�ǎ۫��|��){�m�O�|�� ]5�8�)���U��w!�O1���/���:���j�.���^�*�m�����
��v�V!����Q�ں��=�Y��h�#'9zV�۟!|�6�-�g�/$%��_�'P[栦V��[���#��:��f���C�O!��|t��H�
��*�#%��SW��=�/���g	WE����d�0>��~:�{���z�,���}h{4@�W̋4מao�����^T�h���؎�r��:<�����E����v#�i�����8߽�Ƶx�Z�+v\����_C	iچ��:|ظ�#HA�#�`��s^9~����k۬DCX�M¬�$g$m +��2>�ǒoo����F2c�+դ!ԅ����<<B\�*��~�֡I���\�p���B��Wo�e_|����k{v���F�=V��z��Ƣ:ra:�lݼ�yL����Ou̠�*�2�J��}%_j��VܭEu'n��-)���&�En�/*�� 滫��;���	�<֚6Y���k"�8�g��&$�>Hq�B�SW�?K<Ǐ����7/�����H����/��U��;��u���Ͷ�B������Uh!�������8��6���Wo�p��Xǋ��0jdV%�qBk�ո�e��o����E��xG����H�;ވ�76��9?�h D�(��P�?�k%� ������f5�y�0.�+j��̦6a�r��]Gܡk����4����2򑼧��_ �5���d2E��~��f��u�E�/�
�6���H�����g���P���/�X~4�$[����6ϯ}i�0^��$��{+P+̽��o;2R��XN�lu��suW..\�jfk|��{�e��<Þ�g��24�u���h+n�+�-LS.>>�Q'�ɬ7�1dQ	����ل�C��y&̪%_V+����	�l�XätA8/zG����)J�g�1d��gvD�I��X�W�1�_P�� k�깽�R�tp�m3�%���I�`J�J_�3�1�e��������3:5*�z����C%y������ƌ8|}���G,�1���J���_я���XC�G�W��+ˋם��Rp�񤆒FL	�6�$S�p�4���M�꼨�4�+P�K�<l��P�_alH'�n������ �dC������ޔ]s:o�
��*_��F��|S����
�����BdyB���Mz>����jR���궸�P๴*��Ρ��Q���K�{鯄���BAYy~���t�*$��_)�zl��|������q�����x�!�D���"G�Z���z��!R���!ě�*�w^���(:��T�Ȭ��.T��gL�x�T_�{VLLg�<l�aO�~S��+�Y��C�|�Kĸ�^B�=� �e�+�Uf��2��ي���!$&��J����)�C��i����� 3�]� �,!��ia�s��ˏ��qW���Z����O�:���:QI�`�F�",~3�->6G���YR�׏����TF7�#N �_yh{T��l�̭�Zh���CÖyx��2��Q$�Z�H�R�Q�+�,�c��]޼�UVTh�k��x5M����])�St6�f��M\��J��kF��72Rs����pK���b"gﾈ�/n��C{gY���gܭ�֚�o�y�O^�k��C����Q��=K�g)8������Ӥn,�rU�9F�^�c�B͜���ç�A�z�L�j��+�Ow{nI~�W"7�_�y����^Q3ƢvE��`����>茙qBeW�=0gfH�T�)��`�o�G��}�=S��ho>:I�����û��H�<��γ�q��>b;z�B�Z��7�|�ѥZ�{����;>�%������EP��������D)�JO2���GP4�U�NXLVv��B��3�{���j����g��������C�x���RX��8����#�	W�rR��+,3C8!Y�I.c�p�V8�[9,��蚅��
)U�O�fu���7�����)ɱ�(�ҫ���bY��̽K�N|i:�=F��)�Pj�n�$L��t̾ӥ�nYw��M�MA�&�����͚x/��̀vy����H�Z�PIKRp�mf����̤�,�C�=,��AM�+���}��R�x�E�NY ��=�5
�FP#�.���(�
ۧ�����4�m��$�7�a�F�������O���3o3tf�h���D�4y��3j8Ӝ�����ޣ|;Q		]k�6���HD�x\����J�kw��#u�Lx�.?c���j�CĐ��9wޫ���3�]8h�j��^#�p4x��['��*�}����j�ʞ
3���R�w5�M�us�;����})^���K��Ք���;ms@��g5)&R��FA�
�~��f>�����r5?��D�(��.�����%� �G��.{u��Ư䂸�z�@��D-�f+X�b��ٓ�~���_��.�X�Ĝ$� �i�Ő+�;�^���=\�V��}辢MםbC_=0��m��W�,:|�K��m+��4���kӲ�Ε��`��I��Q��Ѻ�:���hv�w�����l���ZG
�/���L&�p�ހq�t�FoJru�9ɍ��ٙ�"��iVҸ����1Mx��������T_���$���j��~Cn��g�T���v}�Y��5���S8I3��*�X|���;^b#\�c��KG��M�M��s^���3Ǎ��m`;��+��F�wtzj7�J�B 7�<���Ż5KΤsq�7��N߻>uS�L�|��m! �����z:�
����Q*�3�.���$�'�*������3�:Xp񴅍D�#O�V��}���U���A�ӈB,�H��!KN��i�U`�.�w/]{�?���H92x�~������oHF�
ZM׺�䙞��Q�1F�:s��:��_bf�Q����kۻ�\&ڣ�qG�Y''=�H񳥥�L"�釽J�{��0���"���!K���Ө���ޖ���}�$����	��?cXh�/�r���I��ށ҅��:�����w���6��G��>{Ȧ����#2�<D�.9Hw��k��1�'���'��#�L��X������U6[�5�FF��<�8�'kzR�Mڈ�귌��K��M����F�Ps���Ԩ^.���a.�ۧ+��FU�F�/u�3cei����+xA��^G�MS�k��+�V���8�:u���@62Y���2)�0��X�{W�����Q�ӔA 6P0����!�!���n���u�A#Y�lӯ~����߸�VU�}�&$�~����K�X�T�6������fe��f3.�@Ј9i�ӣ��_=�!�c��@댇P�C�e�x����ba�=j�ŊEdjL�(���m��H�u ;6b��n�d��$�7+Y�VJ��f;.6����]v����BGV_bg�5I����	얝+~\͡�W"��ݤ�d�1�u��o���NSH���*���Wq=-�=�F�c��P�����&mӾ�賚�w��+�-جd�{���G&���U��*�M���3�Fv�y/&��;O)]d��z@pEs!æ���*p�����۽R�U;H�ZS�$۪���:S>�yY����f���e���s�Zz����qcu�􂜽�nA;-c����R)x��s��xN,hf�KS�En(r�N�E�g���!�{6<+r���oƪb�GZ��=���4��ss�3�1{e�s�=L�ܰ�M��W���w����@×!r3/��)�.@��J���)�j9]s󹧤��ظN���ۋ�) �z�yO��lJ]���I���B���,D��kgv�F*2Ī��B�B���V�6�XT.����Gn����9��L�4kYYEjҔIU����]u�S�j���=Qk+]v(�feMn]��b�5�s-]f����b�-�L]G����&�ETP��bR��j��]M��ز�e:��mv�0�T��b���(b�d̩)r�暔�ŕ����vˍ���2,����J�Uu��D�-��������v�UrT.��
�ikCk�r6U"�lZU�p�0�6�a��ظ�C*\=�f���d	g�[��m<�]��)�z��=�}U���	�Ue��~dm!�!�0�-�?������M��8�罙�Z���񢈢M�4_��Qn����&֬`�j+Ss���6n��4����ϱ5�~�f���CK��ߘyg.,�Dn�I&���VfߪM�x��`��P�w��:��!b~���ͦ����g��o�<G�P�#L�˭��z�؅�v/��_7&�/���|��]�W�m��ʼߦ�w�D*_o+��B��59�9O)\�3��.�U{:�}@�ށ�<I��#�C��NT ����2�(���W�^K(�WA�Vܷ�b�U��`�e^��/NLX;��@8*;sV��Þ'�.��+n�谛ՓP,lczI��j�����̨ۇal5�כ��A^�)��
�G��������^��13diȇ�瘖�Y�2��g�g�/S�U���~�L#��-x�t�^���"إ��y+}��>fR8� �0j�b��9������������!���?���Ha��x�o�#�(��<�����&^�>��Ml�UJ�D�����PK�����"Λ�=k�N�E�*D�6t��k_�]��/η^��0��U��Q�����/Ꚃ_��%��d-���V�{��A�g��|G�$9������>cf�Y姅#2$g�S��B�����@%��"��[�[�6/`gB� �9?e������`���X��4�OW���}�F�UӋ{��L[]x�J{ւ��������M���up9���Й�)��
��o����ޞgbݝ�l%���U��{�_�|�@*��]�{�_^>�k�Q>k�q��M�U\�۽����ka�<��i&��4�0����3RJڒ�{���g鬝 �c����X���cǕ�M�y����s����S�
CX��(z>(����O��u��{�H�+����D���%:=<�Y����:�~�Y^�mj��;��ZB�\�l	��w͑�U�������_���!�x��0r�e���<��{~���A��*�c��Tb�7<����c���[�����D~�J�n������6Ե�B�Ha�D��We_��^�0Βf/�TX�l�!��@��dp��a�����+e�2�*�Qe���&d$կ`���y�z���Ж&������tkq��R�M���R$���R��_�?LDL��}���{�����D�ĎX��:�0ώ� �vi߅Cn���^=�@x�bZXHU����uJ�b:���k�YOe������N�6E`�$2��~Co��[vu�v��#�|�_�#N�:Eb$�c�?�g���77:��{���R�t��FFO�%�O�P�bEL���Σ1MBCjE����1s���R��ƅ��ZaӤT��f�r���1y��"�G�x�\�9",�2���R�L�_
����^����_�'�u��Q}�mCS3�0���D�>��^�hbf����;^���Q>��aG<B�N={�,Xw��H#P>�.I}}N����9�g�.������r�Z��>��x�Q|��EZ�Q��nWF�n���v�����t�{g��U�wC�I���c��&c��7
�'��u)J�6��E�JC�⢖xz�=oz�=�tPݡ���g�_0(�F(��~�H{+O'�ٛ]h�=oL��]-%���%ݬx��pк=�ה�^�O�ҡ��=�vDX��B��mBucz�����0�@z��:�^��"�1��GE؛JZ�Sd����[
�Xj�٩��&�CX(Q�H8������]{��솏��sM�K�_P�f�#�i �Y~*�۷����K�l�Z^y���șdj¤I4'�M}�[=��ݳ�
v�(40�9�9�6C���*��Oݵ~}�����x��i8��CM���u�^�IEꓥ��v,Wa����E:����m��%U¨�jV����*��pD�+2�	 �h�j�v��q�[՚^�L&��jTTlTP�'�u�']}���%ب�k1��8p>r	���vУ���y\9�S=�؁=����$������!��~\F+��ڧ��lc-"=!ߘb���9��j$�<�o���Unm��|e&j���C��GoA9���=(����ٳ�3�C鲠g�~6F�G ��s�Q���U�Ɛ��x���@*�'��������?V�uhg�9Z�V�%�W�!��`���u��46,x� J���*s{P�}�
4x�&c����VuU��t�B6|/�1kmN�"-a
D�Y���N\�W���1��:g���7nݼ���t8���i�q��H���ێm�uhE,��m��A<�����w�B�x�q6���G]��DWڞ~��#)ik5M@�����7U.���ԅ�$=�y�#�#��w��~C�sg�����G���xQG}�)w(�ǀ����!MX�r��*�O�n�����? �����}�+Q�濋N�&&���[�ż���*�/)˸�������l�F*�i�^��]+��=�Y�([c����J���F�χx�=�r�������2_���:E��bG�o�����!-"_pK���pυ<Ǟ�-qk�g�{�>J*�����x[$Y�J������<r({���OfCվ{]�=)��H_��"z�a6S�]f����i$,�(U�)�FqN�m���7�E>$R*_���qe{�V���'��kǆ|&K8��%�i��DޓW1��v�z�@y���'��޴Y�C���t_\X�,8�IƑ�QQyp$�k[�%�/��	��x�k6=�t��*,�C_����,��͸h�͝���9�����%�/۷��z��4�O��ɪ>���E��ǧ�
�33����$�8Z�S�1͜1����GJa5����5���G�ޕ���D<9�I�I
ɳ��r<��}3�?Xu��۽1�h�*,�f�~�?]+wJ}�.Q�ƈm�eq��j�Gj��L�m��!��ft�Ce���У��~:`��ό�ɑD����]���^���BC�i�q)i��i$�r�������<�},m��V�i�\��w~�lvxm^Wǎv {v���ҷd��v�J���U�)1��N���i�vK�S���R�~������B�,`�u/�j��:p��\w�Hŏ���%�A����HO����W��zQ�]�{~�^�j�Ő(K9�6���N�4�ؙg&Z8,)�X��\Ⱥ3�jL�R}�z�fI����V��84�B"�墐�Z���i�{ܻ
�0Ϗ�X��+;�
�
:h���8��/{~�.	v��ZD:K_Q�����BM���ݐT\�_W)�3�_$/9�O/���c�x��8��;�:{����Y ���#M4-��r����j|q>Hצ
�2���W��H�l(Q�H9�Rt/�(.��n/W*�W�oo� ����&K��h��A"um:3U�-�}��+��λ�\�iHTC�c8�������&EZP)zy���5�S�a����G1�]Z��
w�"��e�ʩ½�oc$Q�y圸���_���ݩ/;:�'�ݘ��1�SCֆ���W1��6C:E]Iz���ŃO�6����4�^!�4�C�4
"�=����^�Gy(hC��8}c�7&?X�O/�����h���i'�Z���B�Յ��;�н��oVzx����/P*�#	6p�da�p6_���Û����������B����P<V�㤜^>Z���5�,����"P�r^��X��=~b;zy�2��ͳ�s��DC�Y�>y�k��|e��.�?�?O��e�2	:_湅��I64F7T�E=�(��-�sE��]n�5�z>�nU�u�	��Y�n�Q��Ŋ'�\DEpo��̵�rⲷov�;�o��m�u��wL������WX�+��ܤ�`n���)����8�!��x7"k@w�7������#�����2��JT4p�Ll�df%�/2v�v>����B� +��X��ː�6	�f���R��aR�
6mQ��-*��0�n�1bCn���V�G'[��f��3�啨Í�Υ�κ�3s��U�KvKt,��S5�7����qsxEۖ��R#�ʩw|w��Y���K��Z�� l@m�kF�����gN��0wrR�^SD\���؟"��]O�����e�Jx�cv]��d���ú��e_��(�O)o0޸�`Nݻ��f��cx��lK1��n�P�x��:�-�^���&Z��A�dM�0ʚrfr��rg)�AU��ǆ��e�د�4�я�8���#EvW���`W̰vu�L�4��oq��+���\6��%d���녺�ETx���<��h�n���R S�LB�\8T�d�]��&�6�;���M����Fc���]�d��Z;D�:���:����b.��S�7q�&h�\]sWkL�m[6��H���Q��ݖK}�#V��2�v��7��]���L�9���G:�bL=�9�Sm�'+4�&�A>Ul�CV�F#'�&Nn�FJ���f�V��v9lb�x��+�0�ͮ�S�C�;��!�����uWuS>���h��Tc�E��w��]��uf�5+D�*�Q24������{ތc�
1�n�Tk`���Զ�*��6�\є�T�5Y]]���DK�UsjUu�-�iF�ڈ2ڣhVA.�G9.غ�9�2��u�n�E�͚溶�Q[lbT��ˢ����D�)Zݬ�ʅ��Da\ʺ�Q(���U�Ժ��9�)����T-����m�V�ͺъ�k��3�gx>>��c��=����跹s��w)Pç��1�9�#'�s�x�z|���9��&'j���S�V�hX������ή��7_ۘ<�+E�<�]:A:W�=���F�8���n����)%Z�i��>����E��qk�⶷{;;��w��?qٮ�Z�P�D5�)f��l�}��}�Dﭲ҇�����1��h�z��0�f�=���`��d�gMEK�S3e������AccP����&?2,����Iz�.0R�6�q�^��k�vt�G�It�"� oV�F�a�F�H�j�u��_a�8�HK��󻿫o��p�#R��o2��}ظ�/o�b�O/��z�W�\�k�{:!��_�Χh"��:���׀��L��e�Z'��[�=.�n5:��*�\�:of�&L����PZ�%����<J^�SL���m��W8C�Nv�����sS"j���w����%�{�HQ|N�7��7�M#�:�I�y9ӿ��>9w]g����
[*/i�ͽ���:Yr�'F�ᙋ��eH����Z8A�^��s;�3Q���櫓U;3/���kf���L����Ëť���[�k�W=;��A�8E�iQ�t���1��Vp�>ytT���L�l�7�-,�t�ϼ�ڲ(</��k��v����&֝h#��?#{�D+X}o=Yr���y����o#/[8c����B�^8K}	~��t��Nȅ��ܶ�z�����:���$�ڿo3����C�.�Zc%� P<��DMV�ɂ�E'���0=�������v^$p�$�MD�}�A�tnI�f��}w�x5��k��1a���r�R���@�=��o�.�G�������b$�Q���) ��gnn������GO��BǗ�g���b&��4w�6��֑j�M�8��|��X�龻�53`͹��o����[���ڂ)�<m�E?�QӇ��>1�r��->:|�(*��K|ZA��H�����y)>�����eo0�x�����h��a�?��M%Й.��}{7�>�&�G���%�,�˥h��W�f?B_^y9/�/@���DW��e˦��"��u,��;o��{E|�ҥ���s,R��P�C�����=Dn��g�:��'�5��I�:��Hq�+����1�do]��|��t��U͡2܍����'$2�c�E9��`���c"�Y��� �����*�v�W�U*~Nf�p�E}k��Qx~&����x��R��|{�nip�l�EJ�Z�A�*�إ7QP�O�`�]Ga�}��k�l'S���"r}KH�H�eQ���&�o�o��L:���sӳ	�9_P�����#?1�=Դ�(���A������]P��L���`��qg>װt��XC�E˶o^Itt���[�_Wc��o�6sK�0�B��
/�骾-����������c��G�����I�+��=�p�)��x�v�:�{6����\�1�:��4�N$^� E�[1���Á8��d��QrC���B��QǦ�ּ��CM���xv�3׮)����r�j׋G�<j�>>$��Fo@�yvP��Eq�ٻ���k��-^���a�a�e��5����>�ت�J4�<��A��;�8sN�Tv9NOn-^޾�3�9�_s^>��׶r.n���;���U�b8e�Zs���oj��i��K���6c��ztaO+�B�d�^�/_���W-���O;�]�"t�MFN�mbh�׻z�A��O*I�4�oL���uh&i�נ��T�F�=r�X������ū������Rٶ��d;�H��(���r�a��%I��7��R^6�/va�N�F8Pe�]��5kT]^�ʥo?e��x{R9G4����]M퐟Kz�':ޔ4QB�%�Vb�D��!XE	�ܙ�s�4MMY��.𳪬��Xq�5K��}���V-b�Z��P�!�2���4S�z�(�5 z�"�>���ͼ��S���5�k�֋��}��8�ik�j�+����SYj:��<�:{�1P��v\E�e���%:��t�S���F�fgM��֯*�L��r�s���I�4�aHt��I�ba�S��r�Vo4׫`��=T]G&ɥxO�����!!z�CIyn5a\;j{jbW�]qE����[���C��C���rt9�-*	aD=i�1?�D�뿾�qrʺr�-dXL��h�:
�:m����q��$C:��ME�F �a%0�G���O92���@;�o�W�2�n��r��ڪ�Ax�k�
O'zi>=n�	�ˍo���f8��V��7켫F�����քg��P���O�V}E�C���d�d�
¾b#�F�K�Yܮ�gs�LT�	`8�ڒm�ad�C��G�]ӱ�\���nEr8��'l�P�&������aD� �@�����i`DAԶTE��7�=U{��k�]$ݷ���!.M�t��QBN��P��#M}R�yw@n�e7^
zͅ؃�L�_[�m��G�מ��e>�vy�H6�}f/�����5��8�Yډ��\���*ZX���S����3�� T����,1�Uj7���l��KF��z3hZ%�)w����K�b��N�FZ��,sݦlJ�.��5us4a�jtWh��dwV�γ��{��u0a-��"��o3Y�9�	�nf��en�zJpj+Iï��ƥrk���cԼ̑���������2{�8�ر�E�l��S�睤�bB/��D�Y�u��3�=t<bk�0�8{�i��^w�	��(�(#��2{�U���&>�md��q(��N)��ܴ�2���7j��XY��i���ѭ�v�+F�n��N�@�9��U�$y�絸Ǒ�����e�@���skqW)�qЄV�����k�C���[O�#�P��x΅p�܄�c��U�xI�e�ޢ��]���y�´��3����Z��d�㜣i-�"��P|"y�Ғ��N'����6p:Ż�c&�	�qm&^�N8���b�bu}Pھ]��j;ی��ƣ��#nI�	|���p/@�����u	�a�Es��G|�.P�'Ef�A��\A�XtI�q0K���%��p�dj�d��.̒o�b��\Q�9�;���.�9��_P��ҎjaP�������>j��I7Պ`��M+��;��������#>jc3Y��7�1J$l��5h��1q��zd.�#�����3�蔕�h[C�j7�D��WHn���
h4�y�!���e
0�F��{t����{]aԾ���䒇;$q��c���<���52�3��֥�6�y�$HY�uc��ɹS�*{��vJ�Y0y�eغ���l�g�sBm��3���0����+��<�Q�n�7�s6�;,Ҿ�Ps}�fs����J�^�2�ڿ�8�K�ɜ��T��tk����*Y�x�@ޡ����G)p0#Z^���cY�W�E�	�R�x��hTq׏�ֱi�-�L	j՜W�˕x���/XX��,�c6b</3�����]�zJk$N��;��[ȋ��dK�{@����n�Z�7�q\�Ď.
4��v����T���4.@u��m���-g�c��xBb�E�W�����3����,@�Y�';���+��i����a������jz�h�7�zQ���']+y)�0Mu���L�+0�;52rL���)��=ה�a�E���q2�V��5��Z쐥����Aű�;s(�K	���t���C�*}��/1�{c�_Sv�ڥ�Yyč2�K�W�V3��QR�GA�b2P07+�U������7��س���n�k.a�]�_����M�P�+v�JH��Nz9|ZZ��,�Un�E鷳c�ƤŴ���ծ��b�6z^f��H���pW@;��~��������sr_��!���)�����y�q��՗�	�6櫬��zjFGc��1����e�9�/�C�2���t讍Z}���JL})iN�]r�[n�eR��֪�7w��맥�bҢ��l�n��Fژ��F����뮺N������\R�sR&��KL�֥
ͥb&K��&��l�K����Dh��i���\ki[nJ��k�*k��]UKc`֔�iGm��݊����뛔��D(����5�mZ[�EWk��u��f(�MT�ms-C&��S*6���lX����v�v)e��m�i��2ƨԦe)k��W6�SGZ���r�iq�kJ\��4]���楦�qrT�QwuU�|"I�m	���bTnܺ�Gnbï����v܍T�<�r��ӌ���h�&���o����gt;^�aC�C�f������w���qifp@��O�[���H��d����V�頖AU���RL1
me����93�<�T�7y�/��Dyr�}L�;��':�P9t"�,����YO��)��z���+�u[9@�ҥ�N�̞&G'���gΞ�]�-��g��/X%eE�d���W�G`omNC�_��눕�5�a��J�6�E��z����Գ��:Z��93��E�L�΁���i��Z�o�U�~^� ���9g�6<ƙ@�+/u)�t�P?{wa����%[R��O5u�J�8g������X��V�۳R,���=��o�*4�2*�'цe/&�u�O"������k�=��ݬ�tι9��uL��&�Z0A��&�k��f,�q�ZW�zj�[Ш����f��|�>#T檺íw���·�I�߰k���v�o��N�"�+�{�R��y%�P��%(�/���ә-�t�[Di�}��B��~����jS����D�Ѱ�ꍂ6������mVU��i��i��O��T�SW+�*�w�Q:��'ݻ0v@if���3x&�H	��nbq�<�n=�q=7��`��W/F�Qe�����]us]-�zyL���Ը����=���Ւ4�
֟��=�m/�d�n6�iS�½��s]z1*.po�8\�*M�G��T;!�FoR�$�L��մ���}��^)��}��W�*p.�����U�ۦL;��M���7�
���P���<N��,�U`Wj�9�}�������=j��U��l�s�Q�i���7�5��/��l��0�P����#�
݂'V��)T�d����(^����ug�Vb���Xa�;hB��Z�D]\�!Q>�do�=�v�j��5�1;��uj�^X	��6�y۞J-��r+�{�`�	4�"����b�SW��zm:vX��y�����}�'�@U���*�@V����8f�R�=��u���E�*821y��'>��C;�1,|�f���_,�.��So�G\�J$5�@XZ�p�'���FC��ė���ǛUv��j��t͝�I!���"*�V�\Գ��yxV��h�t�Dy/\�;��hZ�eB�z WB��3ٵ2<�fy�WD%,���*��x����&dyW��b�z��A��8��ڐLI�4���P��'c20��˔
4�W!��]חxD>��P�͈&�c�Ȭ�l��v�.�34"cS{��� �.0�z�h#lo�/�H�Yx�+��ő�0�����X�L.ѹŶ��Xfy�@�vx�� �����u:q���A���qv}�M^r	.�J�N#����Ȯ����ө"õ�1F%S�&�b����׎���*#��,9�U���t��XU�	�*��D���&d{\���&�0��U]mX.i�=�����+<+�+ǃL���������L[v����"S&�>�O$�oTnB|�)u�"��)�m]�v�ӞGC}�I}ғ�����_�m}r�{=zn�#���7׈�;zr�s*5�ߴ0q�VkM��v:��|�hf�f�K��r�I,��� j?XV����ew�=��x���ٍǍh�J�jΆ`(�f�B�r���Sc�����E�ze�*���&��ʹf��
��Ύs�Η6z���#�zY�u-a�i\��!]^�F(yZ6�h��b�]+��ͭ��&M�2��eJtɸ��A�G��9"��O&d����[�M8Ob�y��} ��T��Enp���R6����V����h�g����RF��������Ӳ6n6��z�7���������n�b����2��x#!���]堬
%���,;��`��y��ĩ[R�z����{\'����0𝍬4ր�uE���f9h��U����s�sq���-\
�5��4te�n�F��ϸ�d5����B5ۍ߰�G��UE���]R}{��j
�q�S!�ό.'=zs�d�apeb�;g�W~����X����h>��H��:+R6nG��Y�*�$Gf���i������4!�s��Y�	�%.��7V"��a��.ۓ���u}�Լrē�9J�U�����9�{
��Z�Y��J����u���MZ�iǴ����Wm_��0"�	�n7���Ox����f��˸�,�(�-����Ϛ�0��3�%�5��tf-}��$�5�V�8%R�>~�fj���9���7��I��S����I6/+|j�z�Z�"b�$���_q���ZOX
�6;��s�2�>v��E���g>�ً��=�r�"/��C:��^�*)���KhB��8*�,�h`5���1٩UL؛2.�	��5]���! �]�麾۴na��b�ʰ���cSp�r"�:JNB'#���u��)P�����=��Տr������ffpȹ��p�Jm7}�_j�ہ��ى,5�j-�P�Cũ�ӽ�}\�A�lS&��J�m��{kuߍf�at���Dd�����X&��fk�Pm?M u6��$��%��I����S���V�,�Xg��.�+D���nѨ����UO\y�7�b��Tt
�v�K�����ó�E�R���Si���Gx�_�y���+�\oTe�ћ|Wh�Stnl����3��}�Q���$>*���L��*��vy̩x&�3��q�m7-'S��g��0�&��G��(�z�omgՠ'�����Ic��p2��b^]�OT!|�3�a�\�U�O@:�4�|��T�r�>\�V���ZE���Ӈ8S?
�2ڻ9����G����ch�!:��S�|2^�������T�k�Q���ξ]೏j|ڲL�c�c����}�<��ЍPk$���?���.j��VԢy���Յ�F7�QP�x���͞�����S��S5W*
���D��u�Me���'�*�<|�Й�2���~����RK�w��IN0^�nU�jn�k��\��H�t��9&k�E�S&c�æK�3R�YJ�'I�ݺ��0eA�z��l�%�V��6����|�M�kFДɳe�=Z)m��Gl�lQ87T�j���ę�t���/SG�\:4�Y����v:ݠѷ'ܭZlJa��������nq�tN6 ��w�.;J����ߔN��қ��l��1��/j�Zɨ��,JX�	�M��f�Vc�휴y��/���i�lCΥ\|a���V7��qywn�f�־=�3`͇h�kGf�r+�:B�O!�5��Toc$�a�;R��U6�b�qԱKy����4�V��V@>ފ��(�6�=p����g�������v�i�bd����[�#�H,1�����)b����$��Z�E&N��Qʱ��:ږysѡ���KvSں�w#�Nnu�Za$��;���6ЌEW��4��s@T�$J�V��^^�!bp�j��&�7Sm��g4�79Y�Q\}4�5���*"���nh�{/��M!�t��W[�j=����՜�ur*�Yf�{�)��)	�x�*��`����h��@f/M��+����i5x�֩}��-bܘ�/�!9	�_�6�#�-\wi��ô�5rb=��e7��J�V8�՗r�N�n���՛E2�N�CZz'�Gi)۽���)�T���Ec��y��J�Wn(Uc�iϸ-K����x��^�5�[�mZj.l.�*]�2�+���L�7�n�u;YF�+�"2ػ-��r�)KK6sm���]t'n�K�Z�nM�m֦�L�sJZ��p���m�8u2<o(^&)�ش-�Q*���0�m�%�ح��囇2��ݶ���]x��A����V�\:і�yNs�����6��j��sKS��1+-��촮�˹g6�u1m�U���q�8py��
��ggk��F��7F��ƗR��Do6qʱf��ʩR�km�Z�0�Q�2�i�s<jZ�ۗ��(l�n�rSH��$�QE3�(�R�__���6+�n=��n'ִ��W�!�:x�2�RGI$n�TkM:�����b*e�����I�=�<9}�˯B�!/s�l]�G1�s��u�'tIϲ5��n���ڷ��諤��t�+�\M[l�������yX�P���ku����Fu����n�m�-�2���YI9z�j8��tM[��"���1,_{�4�ז��A���0;�=�aؖ�8�yqZ^:M��4#t� ��fO+Q_&�i�u�@':vn��nZ�B9�Ϡw*v���:�2�%ŕ��J��i�W>��A3F񂲌�y\���1��a]�N���O"�4دu�E��G�²'�6e�׷5��ֈio�ґ�����ۥ�[>�ËAD���R��ߦ�E��61�:�i�g�鹟3��w�7@����3����j-��j��eu�t�VL僽�SEu���x��$�
tyL�ar �r7e���c�"p�f.����lf��%��
��켳��8a<E��Y�Db9q%�YX����)��L�C�xО(�=;�b�~�ׯ����=�7�ѪsG,�o]��b���"������wă7��I��f.)�@X�ǈ�6d���}{d�8�7��
䕭R�����8=MUN���N��k��>3�U4�)GFr�$!j�E����n���l���0�ؾ�t_Sj
��T�P��u�q1��9��q�i�U�;ijH��<�Ԉ߰FT"gv�.�,���{Ϯ)�s���eyt�E֕k��u����8������ %��x�
�hV�r��������Gd�cJ�.o ��	��O���[��xL.;�8 (�6૽y�W��8ǖ�p�V{b��¤� ^8�T����=��w�7_��4��B��;�7�c���Е�`�f'_Y��庪�E8Eq�}I��V��Q��ϭσ�l�ſ�@�Q�#`a�T��g7���={k/3τ
&,���ᜥ^wF��*�c::]�If)}΋S44��?�u\74?yjx�2M��Z�y�X�<���
ꙣn���*��^M>�>�J�rg��]tH+��z�n�Nx�']2.�)Mh��`����S}y�&_!`����x�06�og��flG
����Wg_/�+������}Rf�2�o5ӗ��g3[�7�f0�l��}v�b63����p<
�j(c��t�� ���![ڨ�IW�tQ&���9��b�d�b��T�[W#n�F���ݼ�t���r����08@E�X����3��[(�{�U3`���7\iS�b������OA.�EA�n�r2��p�aag�N�֔=+^�uM8`����}B� ��خ�t��(�>;��#Ƿg��r�T�v�vZ���\��U��6a����oP���X���Z3��kY�\��$u�_���K��q��;�bv'$^ǘs�`�c�ZB�H����w9�;�,8H�T7��cj�#2�e.�����ÛP�nG+W�����߅�΍"w%�M3ϐ/g�8����}\���)���V��[c��f*�^��µŴ�����w�y��h��؆u�ֆ]G- �luj��Ҋ���{s����R�gb��O9S}��DN!���MǴ���j�j�o�����s���ߗ�_'S�y�df�Z�������2莠z��2�8쮌��S��B�`E�%����ۜ^Ck$�0�bd෽�f��dB�ٗ/w����[s�9��`U���h�u�aJ��d���9Oo��&�]X�;�vJ�]M�{�nC+v;Թ�k�����r����V�0��$U�/�у?��y��dj���uv^��	�[����V��dB7�j����́O�mް/T0k�T	�5�����3.2��Uƺ껌K�B1r����׼�[8y�1���%��Y{
ڧ��=�Y��O\c���~����"y��kgv�$� �P�J�W=����I�+S���,ٖmŵ�s��1�`��,2c1��V�Tv�J��Ε�úg#�F^�jIV�n��7�������1�s�ZC�;O�8N��3���eFh���Ge
=�v	��b��SA�gW�(Aϱj@Ռ�[�)w�z��a�t+I�,�Eخ�Ż���ǅ��~U�T�uǟxK�f�+L�n��gQ7]��<��	��s�֊G;�3�j	����	��ۍ��o�L�w><��9��F�q)f��`륛Q�ud;1��6`���-��cA7=[�>������ȧ&e�Z���Lz�����S���Z��Ɍy�{u⣗�}��D0̆�,�;�ױ�
������i�33����=���J�y�����R�Ԥ=�/Do��I�b�u#w�䦼��ntU4�4�MdNNxLA�w�s-4�U��w|J��ϑ�=N,W�m;5}�2�4�5ɜ��%�z��0z�SQ�CI>{���7��<�8)��%�������Y�7������<Me��Ef"E����.u��3m@ΡQ��7[���6`�Bw���r	sW�C�f�ؑW
f�k(8�Ե�'�zj#���X�jo�O��=V���%6���ԕo�ܦ{��QOճ��"v�� �~�D�M�����Yͅ�ڱ�z�kVqӥ�L��u�3R�n�/H{x(	}�^�J��]a7�@�Q�Y8h��]���n���E��z�f���͔L�j�b���W8:-S��@���L����ђc��F�
`p �%�>��7��G�[`*%Čk�)C��3\ёp���"�&W �SH$(apk[�;�X�eZ���8��A�x�X�*�,}��𾫃F��d���.�U�u����^&H���SǠ���	z��(Kq��������`���%�տ?MV�-��ZX8���Qˮ�������>G�~��b�>�����(V����h	B@� �S�~��BI'����I$��OPr��F΃��D�`�Y�w41�N��pz��g&�5'n��h�hj��LF�!B @R��$�R���:`�`!* �@�JR�����A�f�Ü���@����6�������c��g@�0lbb�
#"�EQEDQEQE ��b)����gX�� ��pj��n? }��B�r�y=��,�I$�)	Z��t#�:�U�=y�뿬=F��
����z��C�u'c�z�@�v�&�x?�eHL�Z�TỆ�<��a&h4Z8��@E) @ �=_�}�S��� R��%$��|d�I$��;�=  '�@d�a1>@{��y���(��0����A�����?���C���������@|䑧�� �=�����0|�#<����P~�i�I?my��+@���?�hx��0�������6�����c��-��x���}!{��}�>��K�~�����$�I���Y�;z�@�q��Y��ڀbI$���:�Ay�%H�	���^�;�N��pv>g����A�g�����s�$�I=�Y

@�I
$�IZ2 ��O��>p=����z�y�hO�?�!���w�Y�D��0�r�p=�����~�I���;���?�g��������_����"JI c풀�@�%��=�Gȇ�!��Hy��
~�U<�����H`�}D��|�}��w�Ϭ>1}}Н1!���/q�!��1�}ӹ����O�<<C�B \���	�	zϧ��?��o`<O��O�	@�}?�l���$$ �B �2~��=�ѐ���H{��~��-��*�v�#@����#���I:'P=�D=`ipS�RF�H|��b� BM�%�~���	�{�����c��o$g��Q-�H:��I9ױ$Hrߒϴ�&I�]��sf�%0n�a��@�
Y�}^�}g���(��y /b?��$���D=~��$���(>����}�`{�o���{@�>P���N|Hp$>�|$�9@���~��zС>������@�C̈́�>p����ӣ���0=P����JB ���c�q��@" ���l����_�����@�a?N��}��3�?���=	�y�}ߟ�id���!��ÿ��~��c;�����s���$���o��S� xs���~��1��rx9������_��>>�Y؞$Ǩ����>��� ��ć��n��O(c��<�(p<���ð0<D?Wp�?�������{O!I���aXx|�z'b ya���`�?����=�#$I$�����}�`?_����BC���{��yϯ�$I$���P}�zA'rv0��ʓ���= �?`u�C�6�w�� �?e| ��p@���$�_L�?�.�p� k�%