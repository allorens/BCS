BZh91AY&SY����.߀`q���"� ����bB}�           '��� 
*���@ PQ UT� �@  P 
$ P"4 P 
�� @ �e��2�(3U�4ֵ���6����C�l4Q��j�CC@�ղ��)��V�R��UF�b�=P t�t�m.���p	�+�F�p��R��� : @   �Z4��	(��R�� ��j�  s� (c�G�`A�1'h��5Sl��l(4Z3Rv�a��[m��
���i���n�AM��v�4��!*� I* ���@1��M �6���j�x�*y�����ڝ���m��vWJ�h�C�)B�z:\�f�i��r����v:-ֽ����oN�G��=��w�����)@6�$}�U@w���aҴ�-K�{W`W�um�<ޒ�[�k��Q� {G{��}]��ۧ}����� �����5�Cw#��>��v�T�Q�5��X���{�_y��j�% ҩ��E�R��������*��˷���^�5t{���A[j�׾_�j>�� z+�o��]�T�h^��}��l���>^z ك�]���OZtۭ���د]� �XiAJ4U
���JP ����u��-��o �V�n����l�Ҵ��{޼^�А�����݁�r�ӷv�NA�E�=�����Zù]v��M]���1�;wt�n��8R��+��9R���5XԚ1})J �����̻w&�Ӯ��:nֻ��Tt�:g]:]��no{��H���[jv�m�j{���S{49�ݩz���g���v��v�
�ݨ4$)!�m�m��R��o��B��6�ݫE���j�c-;�UХ.S�y�m�h{�׼k� -����Z��Xvջ���
��N4R��ʠP�3I��	^>�P[���9hj�NmF㓆�F��օ���R�kmݱ�@�-E�ޭ�U4c�8�T����kTU�����7]�AJ��@dm�A+[ϥT��}о�i[����M ;Gu)B�1R	;��pP,���R���)Q��Gh
�]u8�]��\%:�QV��*2U �>	���������#�Sk�\t��5GVX�罗�����Z�Q^tN;MZŹOx�+���`)*x�  (T�R��!@)  j`�J�� �� �x���#   �� �����      �))*dz��2b  M �'�RJ{R       D�Q�RI=!�Sɡ� d�zO��?������_�O��L�������Wj�gua�7��o��ˇ��&U�>ʠ�?`���H�*~
��� �����#������o?�T U����I'�Ђ ���*t Q|�?���~��LO���ؖĶ%�-�lKb[ؖ���-��-�-�lKb��hm�al1-�lb�ض�b[ؚb��6Ŷ%��m�lK`�ؖ��-�m�lb[����-�l�`�ؖĶ%�-�lKb[al`�lKb[ؖĶ%�h-�LK`��6���-�lm�`[ؖĶ�m�lKb[�i-�lM0m�l`�ؖĦ�KcLtĶ�����m�1�%�4Ķ%�m�lKb[�鍰)�lb��6���-��#ؖ��%�m�l`���m�lKb[ؖ��%�#m%�-�l`��6Ķ%���m���-�lKb[��`[L`[ؖ���m�m���lKb[�6���-�l�`��6���-�lKa6���m�l`�L-�LH�Klb�����m���-�lK`[ؖ頶0-�lK`[�Ķ%�-�clm�lKb[�Ķ�m�le�#�Ķ�-�lb[����bi�lK`[�Ķ�-�l#��ؖ��%�-��-�l`i�Ƙ���6Ķ�-�lm�lclM6�Sؖ�ؖ��6Ķ%�m�l
b[)�:b��
6�F�(�`�lPm�����`#lm���6�F�$b�lm����"6�؈�bl��(6�ب�b#l m�-�A�
6�
`lTm���(�[`+lPm���� ��LF؀�blTm���� 6�Fآ� �1����6�F��b�lPm���#`�lm����
��F�� b����`�lm���6�؂S �"6�GLTm���T� ��ؠ�b��[ b�lU-�-�T���F�� b�lm��`l t���KblDm��E� :cli���Q�"��F�(� [blm���1��� 6�F؂�b#�[`lDm���Q�
6�ب�[`%��Qm���� �� �"��F��-�$blDm���Q�
6�� � �-�Lm�-��6��"�[`���[ Z`+lDm���Q� �E� �[`�lEt�؀��*�[`�lAm���� ZblEm���H�F� � � ��LR�)L`�؅�m�l
al`�lb[ؖŶ��!lCLb�-����Ķ�-�lb[ؖ���Ķ�-�l`[�6����F�-�lb[ؖ���-�lKe��b[ؖ���m��-�la�6ƘĶ�-�lb[ؖ��6�[LK`[�6Ķ�-�l-�b[ؖĶ!lؖŶ[1m�l[b[�6�����lb[ؖ���-�cl�`�ؖ��%�-�lKb[�4���-�lb��6��`�ؖ��%�m�lf��Ŧ�m�lb[���-�LK`��6Ķ%�-�lc�ؖĶ�-�l[`[�Sb[LKb[�6��%�-�ldb[�6Ķ%�-�����G{��z����{^�?v��ɿ7/��&�X�Ò�4Ƶ4U�v�W�E�Q,��c�Wre�;��=��_����U�[W'�ό�;H����p'w���;8����;cQL\��OuF�u�,�5�U.��G^hWJѩ��l�Zq�}�b�����f]'�ʪD!ܧ�Ͳ
W!�RͰ��zc�:��5����n��,�+�y�.�<RՅV m�8�sUr�)G�I�lNA��[��le4����M�
�+5�z�a3j����0�^4"��(�D�Y ��۳��lJ�
�˙��qTթ���`H�N�\��!uNŨT�Eʪ0�(-���,ɖ��A��Z�{U�h��C+f���T^*�GT4W�E#-=�\Q/j��wKM#����-��%��ǗW��!��
/��~6wq�%dBJ�9��-���hm�aaB�n�P�`���{�nGDn��|�fCE���]K�F���]���*���$�̼r,e�[!*�0֌�Y�o`����6V&*�ȥC*�7&����2�V�M�1�,*f��	8��2��j��ܦ�����iF�j�SE�}���M�'N��I왻kp�Z��jb�a����2�7�=ˡ��Me����n����!�٬Lؓ)Sfm����1XxP�d�$z�	r��Cc5N��im�9��X����a���\"0�R^D�ar�MfEgP�yu�1���g^�S56�MdЭ���ys#B�7D�l[�S�M�UN�no�B���V��`�%�b�9�2�HʷWb��y��2g��T1dWn;����Vj����;IL���A�z�M9�5m͵�Ee��˜��V�`)�͕Nr�AR�V��m��ܼui���Z�+^�MQ��a�)�"���T�F�%6�U�=˫U�@=����5��ݭ��[q�]�v5�J�H�/]1w�.����J�D1W��FV�2�C#�e�7��F��-�s�^��
���������H���Fe����M��;vp�&�me�^E�Wb����Q����.�t�9�+�Z����R��i(�	䌳�� ӅiƭK�EĨ:�m-{�`�cئ�o��L<��㪜��K��(�T8&^Z���ҫ$?A�/i��qS�&Z����[[A���MʒX �mD]�`5���2��v]���j�5�[@�J�H��,vk�!;��T�E�\eͰosH����ǲ�e���[s8��v�M@8�:f�&�����{��[�{%����:��fT�v71�����V`��k���"J��>9��B��61h1�1,	M�5&���A�.�mD!Dm�m�2��׫)"iRp<-両�"�\K�v�T{$BAמ�Wf�I<���0��%Y�N�䐧�D�`�0]�y,�*�YdD�3؝!/-�4�Ciėj�e���R�ʨ���w��$ij��Yxi�W�-\��따��M�p�Fʵ�ܰA"j���ưDe]A�Գp��7V*��ge� g�t�v�\�ot����[r)�d����
m(������c��y�����#'&�Jb��V8i%c`��W �.i%�Ly�v�%Xӈ߳qk��+t֌�b
��:��tl���vLi\��&O*|��+"a�m �e����S7VQ�ͷwM�̦0���t/k`�mb��g���8�q82�N��ڧ�oq��[�5$�Th+�n�7F0$���kUb�%y{�\wF�v�(�W�$n�҂ق5��U+^�Z꟪��Jk�5��/��"�e�%���<�ˊy����L��7hv�\�I%k\G��f�]�6����V%YiIt����(ͽ�аp<ul]i�T3�X��^��]�V!�;�n�5OݧYf��2hz캙,�T*�ʎ�g�U�E���m��Y�M��z�E���x�j�l�,f��PRĉ�۽�z᭪�X!���6m%��V���Yiܧr�f�EX�:�	��M��*�pm2՝�H����˻��J��q����u�U�(ܙOc����Q���Wq���]F�.�).UNy��3z␘�c�enEY�Y#TB��6��f
��r s.C������D%�.=��63CD/DA�^�B[ʻ%��$�a��U,p�#(�q;N=���&��:�fX�GQ8�"�+�s1s����6D�"�������yLL�2�+Oh�����s�p̨q^#F�dKP��/V��0���h����jK�5��ݩKffԹSRզ�T[P�5B�ۇ&0�1��ʛO(�BY%n�b��øc4�ɕDiЌ���"���ySj�Mࡖl;*&Bx�&���5H6ܬ��,Z��Ɋ�f��Ki��.]��X�V���h������E �6�+��܍��df��y� 6�"Z�8*^%%e)Yn0��o-�b�^8�Jj�I���H���NB����,�h��-ۨ�u��T��Q��tV�ִ�JdB�Js�I�-��jp������L�*������&X�c�Q�t-G�����c��
���+7)+Gqӱ�ˮn���)�j��6ѕy.�(#D�2�3�^H��*�6�Y~�ob��Zᙒ����6�����jn�"�D�&�L��J��w-�;����ۃ;XK�V�
�YK\�)ӁxD�s���0�@f�[B���jZ���S���Z���44]�L0�j�vg1JS�!1a2�V1�4K9s3L��^IE*���hdV4
���sNQ�� �܆AX%ӻR���4�	�ڦ�-1J�v�6H5Z�*�'R�	ɛ/�dP�X���L��p���ud_�KH+�e]fd�U@�h��YV(�v^ձj�pe������A*Y�RФ�Mf�����X�S}G6�,6�ܼ�B�9r�ҙ�2��Gq�ԍV6w,�V��u)��M�<���֥��c�L�^G!�7w�Qj�]�j]�͊�f���)���-iOw5hMX�����ސ4��+M��*:��9��{�����c��]5=�Y�o:��	� o%��(Zb�f��.�"���L��o��-�@5t��KZ�E��ui�z7Y0@���hVQ��)���T���])�*Y��u�l�cp8���#�Xr�F�t��&��J�Q1f��(��mY-U��x{�a�`�#�q��"���cr�wY���7�W7n��z�Ъ�.ӋrXˡ�����r�@�@���a��n�6�֘�V	Bd�+j���dzY��1�n����ךTi�,�\LT��(9�XAx�U�!b{�A�%�r�5b�cBa����|Ud#Р�VM�R�ܦ++fd˻�-�U�l�AMU�&����U��H����b^;�`n�Q�L*�z4��Ż8١�J����4��r�/E��ckvh�EEd�Y�v��Tw��n��L�S&�6�Vfi��o*X8�
am�d�cjLpZ�2�	J�Y�r��DU�1�J3b�F����-��d��yk1���Fe^�.��u�iڼr�%�6P���2��J�����źF:8����Z��V��c�NRY����8K�BX�ڹ�M�V�i�t���'WB�ڣA�xs4�XHR�^�tޡ;�v�\��ʊ:tF���V�T�6��O2ڹ(Cy�&�ͼL�Y0�7���V��Gn<.�˫:ݍ�ԥ�[9(Y�M,���НĜa��j���$�h1N��W�$�N��nD��љ�3�浱�J��ww.LǐЖ�r��_\'F��8�)8p,�qyM&� ��5�C[0뻭�b{n�Un)u
e��`�a�/e�WiTFM�YK3m�SU�]˰�̠�-�ݗ��m!P�SB��)D��B���!L�թ���A�]�0 �b(�SY"��\�!P�B�Bѭ�*�n$�0�Ǔi:��{Ygk-첷j�ݠ�%Q�қ��u�PbQLgp�a#p5el����W5�U��{%\n�Ww�+V]e<��yw�r��b�E��l�%�.�lZ^Hƛ4����V5�3\.�Zl,J,���h֚]S���M�M]���ղ�d�-SFX�F̣���C!;�x�y(�[S��l�M�tӚ/[��F�"�� ��]S��	$�%��M+�7y���T�u#����b�SWOh꣬�Yv0��FI&e���eb������l�؂V$�6Ҽb��4�0B�ƖU^;H�9�ӣf�Z���o]�Sr���Vn���*�rʬ��r32@��=�m]��k�3r���z��fe�[�׉�=�L�İ#�*!���/Q�/��ѣ1k������8T�KXd�+	#eee���^0η����Ul�wh,V�wL���� ���[��uX\�01d��9�cK��`P�2�����If�Ov�G*�h�i��;�㲐ۻ�ٸnds.ꪮ�k��34;FYT�9[cs\���a&��LDɑ��6��a8Fb.�,Q1�����N.�8$;̈��i�K ��S�hb+
�M�dU�՛f�ե�P*B����[���N#lU�7Q�m��Tu��V��ܕ��vn�{�`���G��J���
v᣻{��n�c�YqK&^����BM�*�a˚v����V٪�X����b��I�y�nctj�1�N�[Z�Q��7.\��bEk0�׭*/F��ln�WLJ�v�[��r�v�lѯ��d������њ/^�b]m�mU"��Sy��˕���^j�v��n���0�h:��r�Y^�,�5�I�G�U�A�1-[wL�P���m����ͳO�.\����:8�`�{X�-��{u1Z���v��b̩����̛H
�N:�{�Y�:lL7L��K����CT��[-���N0JP���SR�`��Q����C|�6.�eI�c>{N�"�2���xs�`����gN+�*�K�Mՠ���<�/TӶ%��ګ'.�V�Gr��fGmmCM%�WkIb�Ѹ-2��hk�>ͬZ��ي�;�r-����dz
��[�9�V^�;#��`k)<d�u&&ӛy6`BD`���(b�!Ѵ��`1j�S����a��v���Z��B���d������*���.L.fS�Pn�E*{f��m��o�����E�Y�Ff�Hm��n��6��u�[�F�!��P�1�]f�E�2�	�&��+!b�Vի��g�Ö�V����ЁY�i���LԘq�T-1�T-ÒC.e,�7��$�.�����t��4[�J���3wT�˰��E^tl5���Z'q��U��;6`�#�e�j��)5i�K��Ի+D���y$;��ml�
��.�)��F�58t[������A��Z��L�{�mMїT1%jd�x����ณ�j�H�[T֚�𵀼�6\���j��]��r�J�si�o1��U�c�2��S����XֻݍK.���Dm�J�ՂIձ�Fm�FܬY�,�kR�D�p;�D5���N���E]�`@�f�K�ҕeܢ�i�a��������kƨ��k
\�d-����� D`��Xz�Ĥ��e���xZ�t�j��VȽ�t�2�8�%,�1�W�x�Oo0�%�Z��0L4Qi�&'��ǰ͹I\:����f*2�M+˔2l�oV�)��.q����a���A�<z��Tkvܚ�u�Д����U���j��kh�mБ��&�X�ܳP����y�Sٍ���;YUwfk{J�56n�,)0�HDT�J��]�����`S.�T�n�h�bڷ�5Z�����c�*D�ҁ�]2j�Zb��eS���T�z�m�5z��yY�QU�Ь�/.��/����-ܻ�n-ٙmɡ�������w#ţ*�R�iff��~�Y�,̅�5O
a�;̽��ny���˰���6MA��Gn����J�xm�c��kիp�oU�j'F�@�<�S �i�㷍MFUD[Vr,'M�չ{o%e�d��l9+6]��V+��Z3`�@ٟ��Y�j5g�Fb��u �9Z$,����k�y���qB;Ցuw�f��q%�mW���R��Z�YR�W�j���B%G�*���&�(�ا����VU�h��*�U�u��^�m�.6�%%Qe�\2UP�v"�*��]��U���unfuԥ�;)ڡD)�-D�,J�z��]���T���-�1>�&��&�Q+���\K��[����f��ܹ'�;G*�F����p��l%�^%�R��/��U�IĩbW;�eY圭'�*�������2�q*OS�T��h��g,����\�-�9m��Wg�bʖ��:Ζ��v�m϶�E�u����n�&+�*;r�b�W�M�4��W������dQ*J��6ܣ��v(���+��+�v^ы(��+'"<��i�Qh�]5�u�С�7���شfG+�r�om�;ݨԧ'.Հ�V�jj�L噣&�:�"�]��u�]���e�6q*X��V�魌�|�%�,���P�iX9X2)R���RҠr�Q�1v+�x�,!�iacU��J��@�I(դZ@�\Eĺ�eE��&�j�+����ZV������փ5*Q��ʪ�qD��Ubcd'-�ҡR�����H{�-K�YT
C�Z����}ɗ���N���kGV�5$���rX�R�h�Z[���%�%Z�ZOiKJ�)�]j��J҈�y:P�r�N䪎����bV�����Ojt��y�W^ {�����1��ZxE,a�n�;�(���Ε�fQ�Ԗ������Q'��-��Od8�bI��%ڧ+���y�*l���Y┗*JM�e+��*�@�'i,�*I��U�s);OT�h&���zs�D�Pd
mh9���T���9H�ʨ����� ȥ椊Z���{��m�z�c\,k�u�J�%@���b�;����"��Z�iOqRD��)<i:�-j�f�˰_Kf��Q��X935\ԋO��q(`o��7q��$U�՝ݭ�e���Ě@��I&��ڑIS/.UnV�.R:����n�5�+�����R1TKQ�qjX�r��uJ��ٗ���S�
�Ǻ{wx�z���j�)������P�~������_�̻5:a�k��z&���ɔ�[}39������sF�n@���cY��w��v6��nZ%�Kd�F�Ղ�Y��l��-I�
ifQ�ꓓzH�}4B���+)�!p�v��At�1n_���6Fq���=3�u����k!d�|���GE��OqW�a��Z.��3t]Yufj�B�˅���ۗA�*"�6��CcsfnZ�����^�-7�Wj��WX��tr�c�`���[B�UN�,���&j2�^m[��@p�7Z8ķ�,��X��iEl`�0U�W;���AK�u_N�:*���z2�v�1�v-]mAEx��Z�:�F8�e���6���)��Ruq��)۷;�TÛj�<w2^̺@D�3�;�)���5j<[�c2A���㚑e#���%fV ��7����S��%�!aׂ%Zz�SVmf����<�ۍo�s.�v�FwM��Y��\��I7H��0ȸPd@��R���1�b2�mͶ��0��	��F����۽�8��U�+,����\)<��
���D�
}��}��A\�|�Wh��&K�^'��Q�u�Ң�A)Υ�����Y� kq*�}�Ct�Ԏ)TT�F��Vg+�n���+���y�R�+4;°r���`��-ނ�d��M"�b�K/	�y�=,`<��u*c���u��d��d���;�Z!c��z�X�:�ui��e)�"��\��EΪ]5M,��1�ʼ�ww0�̈N6Ҩ�H�F�s���_�)`@��|�e^'(WxN�z��ۧ	pE`�;��'�晅,�qT�	ڝ�-��h\YzQz����gV奷vF0�居�)�!����IDU��]�mՠ�N���?U;�#�;�u:�TvZm�EM&[Щ�t�z'"��bۓ	C[��5Q��\ݺ�Or9Ng��ں2(�Td�!��)��H�me���Y8LL��ˉ��Y�,Mh5���Xr�eV;���njY�0��h��N7[̐�l[c����|2RIo�i�Ji*a;To�iحwR�����<W$-G�+�ʧn�c����I�l�͇�T|�z��(4n�N�:"��҅b��z'Br ��c:�\W�Z�z5|������L�cS�I�v^0g>X��00�9�/r|��R�xX���s��VcO(���P0���R��z��{�伺�1J����t�&Bڸ�F�7��6�����¨[�e�ْ�I����ӼޤP;[�6�����}Ht5zk�Iy+I*��!]����Ò	�iE��]��}��6\�-mr�7�Uƍ뙅uAL5=��ӽ]��"(A���U�8�`޴�Xvv�y�:��s��Z(�̛���N ��$V�lA˂mV�B��p��j�){I�����/ff3�^C���^	�t�zڋJ�.�u����t�ns�]�v��Kױ�6�Tk�q7�5U*�78��z��ٽY�s�Ky��낭�UZd���^���(�%fv)7����×J����Ak�lN����wX�0�r�+��B���-Y��ԮV�J���"���@�c%E����Wzѫ�2m�.�.�|�F�ۆ�*�d�r��֫*, �vK�b3&�#��ٌ��_9�Ps�O�Vzڭ������Bpٹ̲����s�[��^�`觍�7S/i,f����t���36\�͵Քi9�E�y9-=�����L�R�e�P����w����H�z�����C�轢��*v:ټ0,jӚ�,%5P�j��7�#���f�nʙv�Wx�tn���C�K*��-;��Wv)��E7�vX��&��̐V�vM��P ��a�=�+S��]����s�,��O�]���)��9��I�k-�b�B,��ҕ@?8tL�.�-,ǕJrMCH�e��+���� ن껠�f�õ�� ��`]hb���U�t����jʺ��ݕ���Zl˳1��;i1�A8t����VQ�5i���F�݌Pe>�R���Έ,�g u���,����a���4t�Oq3�e�\}�sywO�>�%��:�3o�m�.���W:>ٕ��fH�ġ�l��O���o'f5(�bKIb���
��N�����D���GvY&6v�Z9��,�w*�Cuә��'nUcl^�rP�[�&r��Ӝ�����0&v�Mr�YF�b���j��\�:�zDb�w8��\}�a�Ζ��as١,��=�M90�d�	�m]�7J���B:��
A���	=���Q�I�}	�9�fa��nIpλN1��eU�g�F;�۲2�-+���mPq���뽗tJ)7�#�����q�x
Hwp�<�]�y�Ha=��fm�S�K�ެ����*�f����vZ�����F>�j��E[��B�2B+���ǝY�򻇎�̄!jL�V�w�;�*-6Naۀi��Z�a���!���xޘ�b��:B�w3$ch:��tbFE��k�7�z�n��RU60t��n�T�p��}�\��Ol���7��iM����������f����u\)'��.��V;s����(����R�h��2*��}o�4MV>�j�h�h�%��0�JOJ�j�D��i�-�x���-Ԃ�Q¶�i��P�I�k�	�殧]Sڭ���w�\n��fJ�	˨D���8��.��5dv=�A{�!��I)�ա��n媽Y_AOL�j�(Y�Ӫͪ�Po*��5P���ze;w�2rcq謧;&���"�vC��=Mg\&fё�ۇC�c�+	NΤC�wq�h�j�)��=]Q��u�:yw#�t`,�3Y���˓&YҞ�Ԩգ9��cf��Ĳ�:��|T�QP*��%rɂ�&�ܺ��1\C�f��FG��R�Nt.�]���Lf�����W8���Pgl��t9,wb�VgA��o(ۧ��B�ٕ�G1A3:��.Q��N���Uv��Yoku�'��C���z��X�)l��V�;�����>ҹp֗ikpp�����8�2�ͽ�5I���We횓(��ʹ��|R4��a�f_F�;���(ss
R9��0�nJ����V;k5}b���)��̇��`��[�If��ZOj��wP�����w�,yV:VJ�ޙsl����w	u�A2kp�C3�����l㽍5Bz�ʋe+t�n���u�ez̼ûX������c�S{
̼F�QO
Ac��q[6�g\��ilo�4�͢���^m<�:�M�U0��W�W
���x��.���U���N�gpۦ�۱y�:%0�jo�Πc$էj�;�7��I�n���(���Cw�3���6���4�nc�hr,���dR���$n0�9r��al��e^�RA�F��{r�Ά�i�وڶ���L��&܇I��[.�fu���'U�v��L�l�ٵ�(m�.g-U�9��:2f$FVR���u+pj<�6��ʙ[i��I�[�]U�W��k0D�]0�7���HyG*_!���{����U��[��0�FZOn�f;T��3T7l���Lf�,uy�����{6+�k�Ua�km�����p�B��iˣ;�u0�E�-��ҫN"�2��<�OϠĝE��w;G+���6%���ם]��Ot�>�n�ⷻ��T2���,��tv�l:ڕ�X�q���ŷ�OK[�T�w݀��J �n>�R��UU#:Mxzɾ���p�y.ح��5��ohlsxos�������/���o4�fٶ�Gv��P�M�B����l�j�rH�W�=��NqU2q�q&�×Om��QM���f#����.ݓcGX�0��朦)N��@΄Y=»^>E>�w�^k{Yo^i7�*u�7<��U �v�EO"k^��u��-�&�������L֪�۷��4�?��ܷ��n����.�����&���'ڗP��ڦ�Gw[7v�����u�=�K��X��est�����kwƔ��C�b��m�xr�|uV��a
����!p�\#Lib�RʐS�/��i�I]}��Ԭ�{�gn�m��Ɍ$3���z]9l�;u41IG%�[B�o&+ӍmN�xaņ���+x��S��pFWWe����HX��'LEF�V��(��r�4��j�7��Q��ce��5Y���B���W�X���6�;����2{v昶�R^�;�53%fVҫ�\�G��]��]�	�D��,N�P�TM=�ᐥ�Y� �[3^��U��.�:�7�$����·.�bpE��Ө����}T�X��$��ːf�T�
��o/���m�鲯l=X��ݹ�DR��T�-eKn���<�Y�^}�Omjt.�j9V^���n�=��/�]��:�3�Z�{��"�`���l��P��X� ��90r��/jZ3R�؏Z�։��a�Ȼj��b�}���b�X�s��o�3V�����3.�6T��&FV+�V]��.[��8���r��yw	FB�X�U��c:��o=�]�yH�t�Z;j�,c��XZ0p<��p�ww|����n=�\n[T����<5�6]i�mm�p֙rٲCb�\6��1I�Zf�a����]�����Y�010T�D��̼��f���,Χ��ERމ��pէN�hCIJ����ŕE�:�&����S��I�=5�;����\3��(4�7:]����Kzț{3�=����!(7n�eS����;.�K.�g^N޼бoyM!�U�[{�0T�SC�*j�E�p����GV:++}��3�{���A�vH�b���n_\�i>W�W��W^&��ڰM�oIni����V�*˶K��)T������_�}ٚ&Ao�u~+"�*�f�vi�vk�`������d.�,��t�qB͉PrF�Rf���0W�1�j�q�]o�z�Z�y*�8�Y���b�!%����ܵ�kX�A;��c�ױe�3ԟZ�[ޣ���Ҭ��+��`zV�s�(t�"���o�#o�
��������Yd�!a�{p���b�X^Ѵ�[nٗs5^�[˵���a�v�d���F[e�MP�jm�!vj�A�o�9�8�Sh�K�R�B����Mtv�k7����c�u{� �#
$Vֻ2`w�j�rڡj�q�#�aè!M��Uڨ��x3
��HYz�'�c7^R�{��ҭ�lG>sWl�'*�ej���,��S�:{��|�o;zSY/���Z��]����sU΅��̜']���7�7T���B�\�Y}/yjt���W{��=��/[p�W�ۇι�74�2-��QyY���h7�
�eݭn+��N�Ն0�(�12I�ؘgUތ�ސ.��Z���/3���K	�2�Hڛs���e�1í㾦n��ُ̼V�6���1S�-�U����dKKs#s��UH=����lή��`�ٽ}ͩ	�mP�MN�6A�(��Dwr���42u��{���,9V-ܫ�&�� 걈�%6/S��Rr���B�L�	����7E����o�{)e������­���nuI��Eև9fi3�f��Cхg z�л�VwJ��B�N�J���z�Nskm���^P�m+�㛂v%b�2��p"z����z;t�=E%�耐�S�H����k1�{��:�1P����
M��P;L��7��s�b��ˢ[،@�uD�$惉]S�kt�h�X�&�5����je)�`���s�g-��D��2���BV��FC��[���NQB��_l)�U�]7����ҷv�X�CfyV)d*�켪�vo9�'t��+E��qi�[ɗU��.�:s��H���M��Zk)���ļ�qv���_v��-e�����Խ�oiǼ��/��B������uVҍͧ;�<i�N▸r��ZtK�]��%� �걚�Ne"pjWw�JYZb�I�kV�杽�]1�j=���o��T��0�u8U���R�G�l���t8��Z����T���뮯{7�Yʈ��^���ȣ��h��8�Iy��׶��L���TfC|o�g	.슊��jp��Tb�y2��ˁ0��pSq[Y9�o)U$�u%���u;�l�,k���(�vZvr�o���x�/{���a�K�f��8`�R��6�m��p���D7X�� �<R|<�T|=��>�P��������A6^ԝo2ʰ>>l`N��T�(� J�(����؟�ޭ�t�5�5�xi�F�O��>$Jlx@����ֆ���,�F��}�&vOv"o��ϐ!G�P}���Ζjc*�!j�(��L��D�C�[�̤	�=���t�"|�#4��v��th���xk~P���)���#ʢ�sTn{�|B֑��t���'�$0��Ŕ�����ǆ�'~_ i��OBi���}m�T���X���=�� =f���.�D��µ=J���U�ҡլ��"%�MA�'d��B����x �}�]W|DI�~�Ƒ���<Ԣ����`�ͻ����)FH�1Y%D:׼<�M��'gopC���z�K4@����NR��3�������$�C�ڡ<כ�_�@�y���C��Q�T*5�*������P�3�	�}}z)���A����_���������tOe�C'�@K����ɻ�x\�V�gs�p�so���):�2׻�_\iq��`�+L�Qn��v�}I[]��2:�H����'PJ��+2V�ٹ��y�j&��2��Fv�;�R�^K����p%�O�κ(�C�zx�����ìu[1UC)�ʜo$�ՙS&s2�2�[�yْ�5Y��M��ڜ�ױ�k�Xv�A6.�i'	���p��ւ�I�mM�<5�0[�6t�6�y�҅��t�hu�y+;4Wsc��ّ�ªN�m<R�m��F��/1󻥇��ih\�;v���+Uq�\��u��y˟�*JC�����U���|�8�Bep�;بE�k��Y��\Fa����gu<ۛ��K^��Bn^6g\���T:�4uҹkrsgj�U[Y,��7<�"R[��ɵ縘[k<��^���7��Z,���U�r;�).פo>uK��>����"�,�^6�]��mmv��͏-��esb\��[��Ȏ��6L�6^��BBWu �Oue���T��l��&�ۍR�8ЩY�E�v|�����:a�3:���j�.v���v̭ڇE!h��jΗ�ɹ����%�n�L�q�JL�k�Y/xY1'��,�}թmQ6Յ��8��Y�f�*�fN���}}q�Nݼq�v��8�8�8�8��q�q�q��t�8�n4�8��<t�8㏮8�6�;v�����n8�>8�8�8��qƜq�q�n8�8�<q�8��8㏮8�q�|q�m�q�q�q�q�q�q�8�1�uX]�����pS�%W��(.Z�.Ɇ͌]c�6��A�[�V�zBZZ�9��m�}-N{�ުћ;��jĴ�
��ͥ���D 
Qa�8�]u]�=���l�ڪ��$H*����1L%J�(�c 7��u!#;v��n蔒�rv�I��Pt��&E��5Ȟ�!�s��{Ó� dcY|��'����we��|m>�1��,��27tǗ�)C-� ��Y�0�W����)��-iK2iљ�s,��"WZ���F��"���y��U�+a��a3��v�0쨏y�A'"oxe]a
��Â���;;z���(6b�����]�p�����yڂ���Wr�U�Js5�r�>�6}|��\��r���o�^Y��g�n�FĴl�V�;��7oa��!��b�fb�n�	l]�kU ��A��u��\�o� �Ǥ�3Bk����3���:7 B�=��u)�Gk���M�0w(��a+˳\�CoD�n�GX�ht����c���J霬Ӄ�W��w˜՘�ݐE���9YP�o���UJT�,��j�wU[�l��Wk��b=+�`]���ӯ���nk�in�`�(Ŗ��6�� g;��U{ݼ��Ȳ���je��ky���2űN�i,s��uC��7}�ԫdu)��@�y���C��5�Þs�/���<ߞ�q�n�m�q��q�q�qێ1�q�qノ8�8�c�8�8��:q�q�\q�N8�8��]�۷nݸ��8��q�q�q�q�q�qƜq�q�n8�8��q�q�q�8�q�q�n8Ӄ�8�>�㎜s���{�^�p�Gj���#��܌h���Wse��
����{sFd�A�iʣq"n4B��J8�/���93��ˆ�Ǚf������[��`r�%�kk�9){�֚݌܋�H�y6��c�l��ʟl�3-E��c/y���ߠx�p��{+x�6���&�b���.��ڮ�Ӛ]Yo8�S�ə*�/GC���b�4iHI�w �xҵR��S�q�p�����2j�q�gt�f��:�IDng�1�rl
�J�؉���2�(�Y�P�¡�`򷖤���^e&N�v֋r�8��O�sV]�T�$�@zzD�ê��sSY�2�a{*��w�4h���Ti9��T����FHUyx�Lz�5C���ñ�w�OP8��t������z/��i���Ne;껫�Mu�51S���X'\�T�����ɦ��a�+"�U���������F�%2����{ah=�b��C�Զ���j�6�r��MU�%f�m8�nf[�)�5�VL�Ud�6F<���M{�g�B�)v�, �	/����]�M�d����/���E�8�!9F>��R���gn�[�0YB��0]^��S���6����<��V�)CN���)�Bf:��wR5�<�a�O.�{#m�۷qێ;q��N8�6�8��8�q�}q�q�q���q�q�q�8�8�8��8�8�۱۷nݸ�<q�8�8��q�q�q��t�8�n8�>8�8�8��q�q�q��8�8���q�qǎ1�q�=��^m,v�4��s|�J�Nѧ���0�Ns��4�J�P�ۣ$U��j{.n68-!�F����5̺�̱���YP�iӰ&ʽ(��3fe�9�F��C���I*�*8����ĭ�0�-�T��9d�3�;z^V�\L�Q�u�q����+]n�*��7��"�
{4\zm��i��gDU��a���1/ԁVN�Xք4����"�FM��x��,a�1����O�[�S���iW9T� B�H��8��'ole%�Ĳ.�q-Etn�W�i"/l�)?Mq��9x��9[�t`s#��ۼ=���y���o�3]�����и���ԋ��r#��	ZFg=�����}��c��m�[�a7.P.\�����f,+,�k+���]C.死�i<p�D3lӪ�'�,Rg,�vS�T��T�`W,��M��5K��	i�W����r]�@�|r���9=k���+�]�FMIRqQ�J� \6��m>}[7r�+o\}uX�Kw�D5���^Ԭ���ؗp	�!4��F^@M�6v2|<�4eS�~�Gg:���8o2�m�5���qS�uU��A���&u z��ӝ�$��}{�p�o_]h��S��#p�v.2�d<q�ST�N�ƕT�LɹuػB�1^ctNk��G��y��/=H�����qǎ1�q�}q�8��8���8ێ8㍸�8��4�8�;q�8�8�<q�8�8��v�nݸ�;pq�q�q�q�q�8�q�q��t�8�n8�>8�8�8��q�8�8��8ӎ8�8���8�	½�<�W�h��������Y�8�zx8�x����#��r!��6�Z�M\곁׬��mX�jǇd�F�ޮj�sqvTA�)eg^pkwr�dE�cg�;Ue񫨋f�^5|�z���� �髎���U�}F]�v�aB�2nrLS��\�vr�;{c7�Խyu}�+v��Y�)�	�����Ę2�Z6��U}�-�#Z=W�h�uJ0�;Y�3�oc�]
�A,3��IƑ���B�R����r���㫐�}pC�{����)���!�]+�i\��6�xT�y^�K�U�yK�e掷wٜ�{&��(��b�����:>�E�8�/ܚg��4$|�^-a�z]������SPy�|<1$Y�J���6������vPҷq�wo	k�5		�R�ZD���#O9��rFk,뾼�3I�����H��VWohܵ�����w��V�6��uWky�@N^E�]9G)�+.���[/k�kF2�� ��̦͕��m3��{�Go�]V�1������@��VEg�.���1I��(�D:}J�
Ђ��v����k�������Ri�sȰ�$���y�&P���[�����\�`�޻;5�5O��Z��Ԉ��^;�U�pj�+�$�:��w.F�D"C�m���ʙ�ȉ����夢v�W<r��M�zo�GN��I�OG�_K�&�ɢ�F.7�s,�P�Ӡ���,�| �����k��Vku���ڼyqwY�R����Ւ&k#��	oy8�	�~WL��v��nE�zh�R�q����y6��-nhb��=��p�r�k��}$��8(�m����"����S�U	ۛ$��S""aZ�Su���Q8��dV�;�{v曩�H���_�P���:H��7&gcU	N�Ă��&��_���Y8iݗ�fn^#�]Y�m]2�֛�@}�n�DMe��
��+ͭ�.�l��9��@�+����ń�[ٔ5)cd��;�2�2�a�Cw�A��1�����m���xu�^ZjV���u�V9_l�a�u�S��#�<X� �7~��Ә1:���Vd��	;�t߭���uJ�*x�r��*���]�7Hm�Y��[���d�KW]:� "��w�w��kĩ�M�ח��Vsj�`˚�,�ԬAֽ�M�G]��X.Ӯ���,�l�gT�a�I�wX�R���.¥ 5��9:v(��1�]D�.�g*8�ph�Z�0o>�,3��������|-[�`◬�D�TR�^,<�(���..�i����W��uw!�3x���4ޞޥ��yTGUĕS]��fEORU���+ϕ�R���0%�i~z!У�)]�&U��}3
�i�ݛ�NH��vвK���N����Lef�,�
�C�U����N�pmjP2d��3om�Aּ	�hYٖ�*j+x*��ˬ6 �ɆқWU\�� 낄�]�z�h�O$���o{�q�[��rf�=�w���s|ٽ>��3N�Ka8��{�T��wY Y�B9�];��cCA�����h�-S׈Xaܼ��֞��ݪ�� ����o8�D:�����5Jex�[�RA,\h���fp�Y�tܖe�&�L>���<Zw.�0��9�=J���ڄX΃r��}XY�O+�>��M�Xk`r�i�ӓH=s)�ֺ�S5��K�5�$���V�6ܬ�H��_�����C�N�a9��x�{�U�,��;�yH�b�V��pR/c��t�0���̗�P��x<��s)�M�i+�W�hf\9�MR�<.�+�IЦz�BqB��A���
u$�O�Rj��z W'i5�yi]�r=ve ��+i]Ъ9;�RE�/Zb����B���o�]��]�28̣[����gX��Y���CD�J
���c����(Ae�u�c#�t{!j�'���v�3gUb���U<���gNI)��ٜ�9�(��IA@�ʖ���n��q1F��A�X,+Ǹ}˫�"�����&�_fncSs��7sy��"t����er��yZ��Q���H�Z���b����u�έ�E]A��jxd���6���qD��okV�8GhAb
�eM��@y�9f۲f�vv���AS��v����������S�$V����qȅʥ[Ky�L<(u�]T�;6��wp�Gj�yT�Q��5�Ϟt�����Ǎ����Y��r��J�ᇨ�/�93_�i��0񧲉�'�]2��x�8�����T�_oi�/���j\���Ǡ�=ы��q��]��m�3�՜<���|7fmeU"Mm���՘s���1�Q�=�8�T�oUÝ�0�m��*t],�ۈ�N�P��zuY�cΣp�;Bd�f�z2҇1䆤�5�5����Y�^+N�ɻ����U� �J��Sn�Y�r���:�E�iFm2���`��o����16j{C�k�lz�!�zw�y��.��E��5����JVP���GۣB�ފ�I�&[�M�sf:�'!�7\�j�֊��D:s���s2�j�=r��;�m���-}	K�<���.�˳ZCaouY�OioQ���6��#( 6p�.eia|g2h���l939<������z�$<���`�eD々:�f�NLR{	9j�Z���B���=�1eEZ�I�E|���kpFv���L;J>o��Y:ì�W�<���HA�C{wWdmX4ꢕ�t��M�WW3��a�y;x���{_Sa�J����������W!�|�e{02���Ml�)��s;��f֫���%����*mlkH�C�����[��<f��L5Oj\(w.��q��l}b�j��j�jI�j���S�͐�
���:��K2��7p��K�}����WM�[O]MO'�ѽ�{*�ʱ��7v�呃
ړ�I��+��HT���1��ش��+�,���n�6qu�x�I��Z�����.�^]ܪ�U�y�K���P�L)�g1���O	ĺ)t��o.Z�+�h�c���!�:��T	��RG6�i7M���֊&C�M����
�.�)��(�2:/CŦ���fX]�K'n���œ�rK�ے��c{T�I��uD�d�a�N��wz�M�����VT�.&�n6{F�=�~5��oQh�'W��f�m�g�Z;���DV����:�Y���{z��&@���3SE$��q�1��Y��Gsr� ��F�
s�MC ��7�571��q��徧�y{mnZ��2눩�ö�i_Z���}K'\j�J�]b��spWvb��Vr���Vk�uZ��f�R
�;;�~�sR��h�:jU:��M�T�7�r��(��zw ��P�¶�gD�����o�M>�ۊ��Vj:�:K��uf�t5W��b���ȣĖXƹ/�슪&�ANF����u�ʗM��H���'��}3N�o
��U��Q���t�=���J�1Q�=�o�l�\��[�H����ako2�z��2����ѩ`�/m�*�g��1-D�%�.�Ѳ�r�F�#�`�\U��i*���}��N��l$�9����R)t�[�%nV#�Ыf5ni���U�5�㸚������+���:�lH/��Lx	���z�.B�Ͳ��[�Ֆ69:����4RԻT/�]��h��W����W���Mٓ�b��2��	��9�U�n�9�`�a핔��oXK*e��7+eL�oKR�;��턝)W�ˋ%�Z3�[n6�OY��yW;�=;��Fw��J�ۻ�����j��s7"���.��^g��L6�Bi@��v��a��+��ZXI�5����Y�g�ά���������[n���Mں��U���v���1�ˏ,u��;%M�%�Ŝ�J!b���X�lPwH�
���V�x\���Vlƥ$�*�{U[�0�͊)�'lg���c� *����7����޿t?���?{�ߞ�R���6�t�$�e !?�T]P��
(8�^`��q��4M�P&i6 .�0�A��B��5%P�B�gɪ�(	�2g��P/�uT�i�M#����B\&%)r�z2�B���!Іt���.��b
���	��Q4�1��H[A�(��J�t�SUU)[��$�y
UFL���MB!m�(�*��Z�R'�*�nSL
"UB�B@��!!Hw���1[τ­>D*��8o>{8z��1�zhѳ��5i�{��j�{+�MK�&-��ĪN͓*]��%n�v��/��[P`�e�{&J����6������r�ɋ<�tr���x��z�Ce
98Ȗl��Xݸ[�*�[�������,͇8������֪b����!��91vk&�`nQp���*¹����`�Vr��]�*�;qDO�w��^�թok�Α�bva���#ŏF��U�ll��n�Un%����q�z�](�x��7y�I���:[4���N����U�z��K��[�:��7�s]�Zojժ�mM�w2T-eu�o��2��T�D�U��^�,���0�_]��� �����b�o�z�9U*=�w�j������w^▕�#W�-Z��ud�5O�6-�:#�j[]A�VL��چb҂\�o-�9tt���jh�!6��"�.�*^'wiT��nf*�\��iI@ŻzpÅj��m�3K�+emm�-Ԛ�jܳ��|-�bB�[Bkq鯶��Xsv̺FAhe,��z��PN��t��u��l3UpS[�Y�"�horU�J,�'א���6]��Q����R(��8�N��VL�Jz���?"�!�`��(9T�J�4�E�D�A�#dD�p��P$���Ɲ�j6v���bH�p�(Y)��kĸ��$���!0�4bLKQ�#-FL��%�ƌ"b)��D �`�E0[��eBrUB�4���K-E�Q&�䌏>�'w�Ͱ�o�9
!&I�(6���cm/h"j&� 0��#R��M�d(���1��d���jK�O�B8�[~J��]#P��Z�>��D&�
�UJ�к@�$A��U@�-�F2��t.Q�H�D
��4�#!J�0F�)EM�L1�[$��1��2ÎQI�PY)��kĸ�\J6�N$$������	&9@���
x�K�a%���P�!A�N�B�")�l���-U8E,5�J�&���X�A�! M�T2>M@�22��uLi�����nݻv�۷c��űW,m\���msZ�#ӎ>8�nݻv������ jd��"j�i�\q۷nݻv������I��=���wk�ɔ�i"��gwASh�#2t��z�Ǐ�v�۷nݸ�z�2B@#YZ0}���p[L�f-��$S�n��5$D�-Ͷ6,�Im^-rɂ��FLRA�h�1�J$���<��ӵ]\�1wqZ ��E^.��y���5��@����4 B��و�@ߝ��i�r�0�-�c1ㄜ���c^��6�nr�Ҽ��y�Qj�P���5$[�K�ҕ�EQQ^+ڮ�Ʒ���׊J���\��c�ʹ[�W
�W+ok\����(*������צ�����i�.
��eHڍO�j�T�A�h����29?x|&����q�Mp�
�����h��l�.�L��Vi����f���ݥ9J턱e���"�*��16�#A0�I"H&DM&٩DWέhP$8��$���$��rS@�]UR0�Q�IMHϘ ��6��L$!e�FJ� �0 '��$tE����J�'�`�V�[qB�HGI�@��<"ھ�+8t뭶ً�g�'즟�7?ݯ�d�{٘��a��e)�8V��4��O�c������r���*S�Z{���xXN���{��Pq&�r6}�x���g��z��K9�{CaN��3�ϟ0Wu}��y����M>�WQ��c#��t������̞�U���BMñ˫5�|gݔ��{�[��_V��M�)&���-���$Bn����ܮ�+�����g`-|/TS֪��X����_S0w�B��8p��`�*]��d�_T󺟰�}h�sy���j�p�'Y��U�u���8ɉ&�@ߚ9tE<_L1�!J�����[۱�*�'��$��д7��nu�Yr7|FO�%R���c���D�{���G=��N���բ�:&:&�%+���^��HS���zf�֛F�efc"2g�l̛��-4m<�.��m�o[v3d���fØ��9���m+4�����qlʝ[�ΐx�D��;��t͞��Y���J�闩^��6������k{e�y��
p �E���͉Zo�Y�t�7�9���a2�%ַ��l���yˀ����p�4��s���geos����}����"_Y3H�v}�ȗ`Q�_!�*@xj�1vj��W\�4���l'�]\�4��������4�ul��I*�.������ޓC���l>��zhC�����5����;�˵�d��PV,�ᑏ]��a� ���(k�Gf�J��s��r�碶��<TfSou�.F��nU�����G�Q��bEeKU������c%��Y\qk��+���r?�c��)��tt|�|���^�=�ތ�q��g#-#���ޭ�wrϜ��5Ci dwmFg�+�.u�%�n`\I�j
��_9��![��&ퟣ`�'w������r�#8��j#قt7�Ϧ+�[�aKD��+�7�b�Ѹ��ܾP�U�t���	Mq�ed���j��tm2�]۽@L~�-�<YΪ�d7}L��@�u�%>W���łr�7Ծvc�EZ2p�̼p�4-��ah��)�.b^	�4�u�-b	�6 ���tA���u���E����9ˈ����7jΘ���҅;��y��1"�hfY2�ңxz�b�8��|�5ՍDc�[mN����7(����b8��F�y�zt�u	0} ����������/�Ի����<ʺ�n����+�t�N��w�*r6�5)���M��#w�6,��̦��7��A�����r�W˖_Af%|���k).��=vʻ�~\�����=;1 �kE�&�#��M�oqk���j�}@>�o�q��l*�Z-Y�B���P���T�۽�k�t��DGڬw(��)�i/�T��7�v�Frx�%�%:�w�Ͷ�Jj��.����H�}��$v0�(5�v"H�$�vwT���Bu��K�;�Rkr�@NE�Ө8z#��Q�5� V�Րݴ���I^m�+�S���m���rv�ٺ�k ���\J���jEE����%J90hh0n7(�!"p��V��lJ�ܝeI�q���|��N]�&��de�l�Id�^�gB���Sce=�CN�6����-֦�[!E��M�ƺ���ʹvDp����wYP)M�5{�`�81���ᔾ���/��z�ݢm]�p�W�`fD�y)�:������w�Y/����y���b�n�wg���v�-1mG^�ȩ|��G	:��z�BP�>ޑ�Z�C�YB�¨]ݢ>ϭT������F�X���}[R�������a�.W�0���u�r�7�b�������{�!�]�9���vVQ�`�~U�;*z�nQ��u�K˲B���M�9/�a�4%�(!���o������ile}D4'���Χ\��v!��I��4�>�_��:�Y���$��F����S�������:����7�G�ʗ[u����U��mi�/}�f���l��}���	���փ���V����PyF�i�+�WLD�jsm�޴-�5Uz�f�Rk+%8U�]�jp�Mc�-M�����p]�.�QNYok5�!X�}O�
�A+B�ܵqU7n�RD���i�^G��M�ҝ�K�u��6#�h�z���x���ʑ��V�Z��Y��n����1v��oq®�4�6��� t5c�����)� >�#0��L�˷���c���f��~/x�=�5qb��GWƌ X{1 r���S
U}dA��:����{Uv���2,�J����8]�M*yH�<�>]b�Z���rȓ7n~?y�����HMu}����C{������9��Zuó�0.��ڻ�{'�Pl�ml1�hf}yO 72�MG�]��\�9��L�>�&�����h���y������Grw4����ޠ�N�S��8���n������{]w;xT=`�b�ݛ��n��KݰC���_Xپ{t;�f|�ץW'w�1D1�J�z{��M�;}��6�\���C*{`�˻��S�ڴ�/;���Uͬ��)���k� ȃ�+��
���YzZ��"�rs�iCr����c65���!u�r�������n��l��Ivgb�R��p�|b���;xks1]�1��..ᕖ�(�?E�im,N�dh��}�ޓ,����mյ�sk��yTy$N|ۤ�s#Y�� ci�a�qw���86�PyRw�>n�'7�Ϻ�A�L-�ɷٽ*�.��Pu5�#���縟9�\�|�����"]����[��9�f��PP� ����S7�*��`��ϛ���u�)�,�h�q�1����{XW�C�#z����\e����'��؄�޲���U�ET��jE�}�>���	%67<���ko�����/.�k�8I�㗺��U�^%��?j"ұf%�:9��c�n�d�����Hw?��H��j|�?gd��&Pȼ3r�mD}<*��KB�Zs��-Ti�����uyof��tF�]�g͹��!�{1�p�F�U;�t�\uj��HS 1��yUV��[����ov������i�{����+�AU�$`N��P�n�v��Vw��s�*�$I�Z��P��>Q��u��8�TT�U�و������d�����"��6��5u�-a�KF����:�|�iG��qX�\�9|������'p�F��V�1+!�޷�3E����V�N���Ûa�̕������v�� gY�(^�҅]Wu���MMGPc�O��J�<�@�3����t
��:���.�׉樼�l�����=��;�[�JXr:ZRA���`G^�f�����x�H���u|��
_ ��vtf
;Kry@w�e�a¤��;E˝������7�����q�>�>�o����X�6��.�SI�Q��W�	��8��1L|�}���P��KWU���GJ��I���	_WI�콄K��<w�z�}#�=0��*{��Y�~�>���\շ����R7'�<%@sC������<��Tz��4$��8���X˳/%��ޭ���s���rC��ñ7�0X*~���'2�8���W�v;���6�v)�Ӻ�=�&���ƃ�4 ���r�c4�q�Mc��8>�9\�gm=��?`N��5Md���?'j�*��Ϙ�,l�bkP�U�?d�u6fEm����g��WM��}3��^U7�;�o�ڛ��{G.��u��Q41��&
6���;p(+I[;��i��#I�QA��;�2D�b�'�9ok�ծo)w�g�{"�_f��h�k/i��9�X
�{۪n�]]CD?�udl�o����~��lJ��>�/v\����Q?V���Bi�����[�SA��op��`��3-v�'��bAU�i��Vcg�@t7;8.米�W&�g�i��N�u�����)��W��q�}8;��̸ƒ<�Wv��r�$�giC�e���W�e\�wݗ��$p辅�اYx����5v�?&��y�C�W!ՕCm:�Q?R/��Ih���͓���G*����T}͞�f;������n�.�M����oy�S�ĹVxP�m},r���W��T��A���`�����o�[έrx1���47X{�ܯ�L*�겢��\�16jgm��n��Ea��ڴ}f�*>��c��[9x�MVH��ܑ�=�x�Z�$�dH�{�y˙*%f9��8��x�k6�n�$d��t�۽�4k=W��v�ѱ�����]+�I�ڂ7�6Vv�F-�~��LL��ތR�*ݬ���/"�]Z���S�8wa&�*{�CY�R�IK�b�xOp�38��URE�(DB��@��rfg�3�|��NOL-����ryoe��3(���s��ó!�ض��D�.��="�{[��k _�<m��,��Å��QRh����|��O@/���w֩0,6�c�~{�ε|�e�.�����Þ�q��j,�=����_CT��B�Op����rU�ٺv�"�Pw`��yۻ��6�́���;1�?E}c�:����Z�S����G[<�̻e
\5�D^�ض����H"���x��<ۍ}f�Mn���3����\�/�Z�pIb�`����04	��\��@15�ӎoR���W���8X\�|]Y*��&`	!��We������aUoΚ������F���1i�ȩf�vG^ѯ���)af���h�:P=�DͰ�oh5Y�ύ��;o�No�]U�]�P"{�Tܣs��xͭ��T"�s����n�<5������%PR�|)7Gs�eɏk5K��J�3v�d[ݫ�5����\���X!uku�����Xj�:[E4�
�UrY��W �7+IΆ��e5��Y����r��>��r��2���Ӊ������"7dv��n �᳛˽ۖ��\b��fA9'�b�u��Ԅ0�-�@#!G�u�X��^�Q�,�Y���L5ӟ)�!���Pd�$��U9�q�>sp�VZ��E���gY�S�Q	;���34���5�ρͯmxv�O�4�s�}}z\n�o���0+8W:�J�'������*Oug��VWE��'_A�޲�(����"����O���\�|�;W�cx�X��Q�B�F$B�.0Ϡ3�H�v*��ꮡ$�)�����R��DV�ƾ���wW�h_�p��y��$nZ��I���W<�l��}Ilc������_�SYA؅QB�`�>�O�ʙf�T=�Zy�ӌ\����Af�!J��6c���F4>>��|z1!D�Bro��.���މ�qvQnuep�Xh]h��D�%j��T���s�c�c{�
�%����[0�Ĕ�9l��1ɖ���c����������#�*���E�a&
��VK��'`�1
ܫ�,�"��K0h́&(�"U^-H+�=:b{:TVTL�j����Ĭ].ѽ0#d��k/ei���x��a*ʪ�O���e�I{�Q��j��Y�3ku����(�w�WQ"b�W_@\�(��/vi=�b�TXI�惥B��Ն�uۍSX䧹)�-��vۈ�����\����U�y!��=��w�'�[�L���ڋ�[�&2V&�"��[h�16=W4��T�$�+;l��t�+jfN[��G�WZ����Ll:$%0�m��[EsXn�%�u����6�k�
�ok�P�T�nc�
�������v#���r��bࠪ�}���og:�ɹ���a�P�ʈj7�7;O,}�e�޽�-˺;!n��C�{��-�͢�1���U�3F����l<8���Y����j�,Ѭ-w�������`Te�-�]c�]�X����X7hf^9��oݹWݜ% ]��ӍX�5�;D��W.[���2������o�]�z�G;���V�������F.�w�̪쎹�0r���+�qUU��{�����A��U�	&����kzn�K8�%���Hr�j��H���WV������Euϔk�/8�GV5%��!�������b6d*�̖u��g#���a	�æ��-	V�'�k��ٗ��Q�&���٨�f�N���ׯ���󭛴�Y�r|�����W��k���v�x��Zi�E���;�i��WQ9v]�o���R�P�4-j�����)�lrZ�:�0ܵ�mR7Dm�;n�����+:��
��uQ�	��t.eZO�VJ��,l0~-n�S��HGq9�XZ�R_80h�h�ͳ(b��1[�d^�}~�UR��C�"�7���B��*3���c�� bq��4�����،k�(L7���
�.`ڻ��������M����r�wW�J�g�k�������*��X��x�;[­�K)�Y"��4^:e�a	h�7����TV
R�Z�^Z���N�0�G�:���wM��|qL9�E��eQ�Փ��!R��rmk��4W=�+xqj���9�{R�ަZ���H ���:����Ju׎W�f��t�^@nj���UMf�����N�K)u��Y�xF��ul�n�>�uN�[�3	�Ð�T��l�iO����7�FA�[mꍂ�s4����)�����{W]pَ����v��(H�3��ٳ]�uU�Ju��ܸ��T��5U29bc�u_�~�Ѐ	����@Td�R1�o�ݸ�۷n�<x�ǣ� �H!$��B+	 ���^�q��v�۷n߻��o�o���[d1���Gƞ�|z���nݻv��ף��������y"��v��	�j�F6��ׯ^<x�۷n�����Z2��-Q�ЍnVỸѰZ�WM�QQo���;�EIETTlQ���~��6#�Q�b1�LѴk�oNQ��v� L���'�~��cgu\4G�1��I'�O� x��=��XoGsu��ʗ�C����tp�n�<�ܵX��
�&v���ܡ��Y}����g�Ns^��T�	�����5�s�{��� �
Un ��8�������Z�bQ�/G�����	�}����p:���h8,��g�7B^���H������ �P�.b�?	v�
Y����*�1���aX�_�c�y/&o� -���(�7Ҁ�ֶ��4�3��SאE���lm9oCy��
hZ�xU�ʂSl3����J�WY�{H�f�|и���/}ㅸ:
]�+�� _�@�H?; �#��%5��kx~����/)xz�qꚠ����7z�1���t�
+�p��q=	����&����텏���u��z�� -�ne�#Q�X��$��\�^^Q����Μ�9�DP��L��t��)����ޭ�R� �����	�Fc�1	�E�?D�VT�b�IB`)�t��^��oC*ˠia�|f�	t�;�'+��ql�@^����n/8j��}�� ���&*ۤSx�*y�5�1G�����5����_߽�f��JU���A���5�x���A?qk=P@�9p+O�F��r��y�-*)�.�)���@���v� 3&��PF�h���25����^p��s�����WOYC��O���zmǇ����G�|ݘ2t��v�C>On:*���׭���T/��uv�;�$/E�{�b^�u#�5۔D>R�g�V�t�պ�)oU愮V3�8g6�����77^'ww���[Cog%�"��9P�Q�A܍W��2JyG�p#�c9]�����s� ﴜ����9���$���(����a�$;���	�W�C6�	��U3��T�r��9{�ׯ�nb,��q@���@��UH����6!4a\����%��������˦ײf7yx�� �{��Ԙ���<k��u�;�%1ߣ^���2��z}�!�g`�ў��E��MҤY{XgY�����}߇�&S4@Gr�"'��fcugZO�y:�a�?�f�\ź��^øB�yކ�\�����e�����:�	���>�vo����%q���V��2'c��ߪk�I!1��TWJq���|�o| ���}p�fȓ�A[���
������@��b���5��s`�J��\��U�nJ��~.#��'�lig�;��W��@6:�	��rϲ����)J>nׄs��1��\q��h�<�K�g>�,�����x�����^M��m���L��
w�
x`|N�Lf=������ ������ڏ!�{m�,�h��-���#�
����{aӧ�E:�1�_��3��2�!�t�D�i�=ၣ���;Ƹ�l�d.g��{|@�� ��Ĵ��^����~~��0}�;�.-ER���s)8`+0kb�2���RgA1QTܔ��p;A(�2I�Y�"�@�]�4LD/ :���}Q]�l�
�fL=����\����\/����R��\mc�;r.�n�+���uH_��+���������")�s�>��5�س/$R;�T]�
��E���?��M0SnQ����#��>�w�>�9��*c{�2!7s�'p)PU
Jx�1�/G�yn6q~"�X*��	�od����ڈp>���	ޕI�. USpZѼ���=��s��  �q��
�p��X~��i�۸���e� ,��u�-�!��W��<Y��	�R��ƺi�ý3*���`n�1M��y�<��s@�= V� �:�OΈ�B���L�=/��7l4Dq]��܌��-����W�۷�/g<0j��T�K l-5;��}�b'ø��fa����� $zV.���xsi��/WO�gF������]<�l}���sIzw�4F�3awn���� �x@�-���~��y�g���a�j�b@�OB�)��ze*�</��g�Vv��!�Զ��7� S&��	�#�@8� >'�vd޹��&�ԫì�{���>���1yuҶ� =����%�|��	j�]6@^�Q@��	BG<@���~��b�}n5֩-���IM�P-�cQÐc3��������2̩��`@:"���g0���s˺�aZ���d!*Y�V���׽��"��
��i~fU-���,���ꃵ5Z�4�M�7�0c��j$�.� ��+^gt�RMt�Q���Iwзo��!!���/2>*����~���mr02��h�3�t��T��T%�=�����a�M��`F1��������]�� H|������ϔt���@��ה��z.�	��|��T?���P�9*y�җ������������]\$��/a7�P+��F���ަM�;��}Y�&��u��9��J���c��B�¾��t1Q�)���� Y@;��[W�X!ʳ���=ӝ���6!��pe]����_���>�$�v^�� �|�7���4�L���L�)��q|�^^�l>4�һ��s^�{״G���_��i�v�\�L&<�^�������R�y��s6r�A��ts3j���9��]<�5zT|���i�Osߋ�:p$Sۼ	�aAp$�T�I�����ʡ2�U���vNHX�_b͌]��g�-U K�1,����5��� ���`k�L[��h��6>��@1�?m9Mϟ���xc`nC��ïc���yN�.U(��p(��5G�WN���$��@�ڌ��)�������|4T�?D(5 ��z����Nߚ�%��:�/I�� -�ǹzc���� �3�`���=�[�� �4dL�9����!�:����{ƅ�FO�`��b-�GtU�5��U9{�ټ'ƣ5��o�wO05D9*��;�%��x�����E��,VTz��Y:q��aG,iT1+ʫ3.	���_X��jW&1��W|T}�h�F oz����(I՜�U�#��3z���W����� ޼{=������a���� ~��-O��G:����>�8׏���$K'���a��c����%�nh�q�n����Ň��_�kjO����@�Ø����,h��h��=_: ~���X�Ռ�^gs5�C�_�/��/�G|�y� ���Ok �g��v��0 sQyӾ\&r(HhS�`�7�{^��N�Y3�·����G�6ǖ�oҴ9�� ��S��ߐ��hdT�kø����{�i�Vev��l�W��]ŭ2
NJC��b���Փ���l!�ٰy�������i�}���x��*߫�%�y�[0{s�oiP^��v���hP�a� �ץ�ލ���}W]B�y\E}�u��kf=&����f�vήj$/{����p!�k�<X���8�k{Y�-���{ij\��*�e���sT�m�xw`/��v�x
/��L��u����o�|gF<%޽aŴzÀKȋ�Ky5�&�y=��*�QB]��OW��6��_la�%�%��6��}��B�i�����������Xa$�[3��r��{i�
����o�bY'I@��4)�A?c�q����i0 ��.�n9ki]���>89�����j��ˊbC�S�	7��.���XoEs�Dm�W�#����[3����]��D��J��|��r��S+$�'4�32X%*�QS;Ys:�8H��v��}M_r���s.�%�\z�
���c?���<�����K]��{��!0a�h�Ts{|b�[��h�oJp}N�IRkk6=�'�.`7i<(L�sU�Kw1��� q ��X�sյ:��מb���}*Qtb P�w�*����%o�&�t�:�^ T?K�=����
 ��_������>�Л� �����jb����1	>!�I���{�����灉G���s���;�Z�`*7�E��\�$�k<�4ϓ���щq'�1��� ����́�a���7'ԇ����f�ׄ��� >>�_���τ����Fĩ���|Cަ�>����c�S�X�x��W#������.p��O� M�{�=�b#fn��YB��1���-�Ԋ��6�5<��N��Q��n��~P��:gѰ��m�2�גg�J����e)�3-�	�=�]���,���'��i�	;4k�	�ܴ/taɱ.�Q�
��V��s�{�@А�(��_�7������ǆx�7������������z:����^<̬  �G��Ph���Z?��A��Pa���� Mj�t���S�B��czi�x���Ȍ�?T;�Tmh�̬�i������L��rr�F�m	�J֌�ꠈ #� a�t@a���ѩS���w�1hF[Ul#��]���)�nÊ��n:��"�>+��*�[O��N�NK3��J4��|<|@?����z��}���4�]��j�T��b�ϼ �@�/Ῐ�@�.3%�������sd�;@�c�e�o�[#�p=3��42\�-*��������l^?��C&�%rI"���˜S;y6{����xG�Γ�Y;���G��Ӻu���R�#ӓ��N��.��l��d	`�ʊ�z�𛘨�A��f�z�m%U��
O��n�>[��uZ�k� vh�[_��3�<�w�������ZB=�Y6{$��3�TM�x_�<�> ��:�,��~I�#!�|��"j}*�� �[�DK�VR�T�v���T�u�������%�N8�u���N4��t�z ��őqb�SQ���^�ҩ2�Zc�%<������_W�����j�ȮzG�מvj�]����i�I��0��-�2��7�Wsñx�d7�w�Ɋ�:oZ���\�6�zk��������h�}��7p��C����vOX��^3��nZdK��v̞xj�r��/��,V���& H�חq���9a�IH��&���4 ��5���_��������RX[��f�ְMm����h��f_�ѐ�<���6S�F P�FE#)wL�MT�f`�u��/���6^߭��$�\C��f!����6j^w�����˃��"#P��n�LܬxQj%-���E�^2]��6�ؚ���iU�4�4�,B��q�%��>0#�0h�|�|�uΝ����#��ߘ9`����]H�3�E&0K�v:�PK�B~`ru�t;D�f=k�$ =�cYcۿO����7I`*���\����Ԩu��u脎Gggk0I�}��������>a@ߨ[.Ï��`�P+����h��~��i�kn}�A�E�{��tp���0���мۆ1��1)�W���	�4E1��l�@����!�님�C!�ȇC�bz�t%�����8�E�^D�NQ�r=�{�7����O���Q3ց?�-�^e���ȅ�i����"�3˄#�c�M���{h��^Z�a�%s�d��U>m���Bn��{�Ġ�M>4^�&�)����V�?h_r�����0;<./�}cc�b;8��һ��~Q�ҭی"//�o���a�}O| cF����jaدf�^q;�J`618���ig�ju�&����ݼ�PX�R�
��=��#J$�F���k�)�b2���oeW4�	�c��k�j@z�DK ��ux�0MP��k���z�΃�[��qV���l8I�W>�K:�uJV���;iD����'j��� �ru��s�Q�"#\-f{R��ga���ognZAew�ڪd	��2 1��1�Ċ3��b����m]6�z0�6n6�
�yc)��lIL�`Z�(�8�X��w�Y)�ؑ9��n�Y�|/�}�>��4��R��	�g�hq�HDֻ�g�}�>�S:���,S��}6�@�}i��E����\8�a��˩N�z�y��������3��f�Py���<9���ʥYϾ�caw��~��|t%�ufD(��8����(��@H��9��0l��w�J��I�O���q�O�S�%t�~bH��N�jr�3�ђ������)��T�sP��0�]T�5�����#Ê���a�8���Sz�]Uө�x�������<��q�W4��E��TA��X#d���ى9�O�s?�VvyWk��V��Y����w��1%�[�{)ԯ9��F&*#7X �D�b��.�O8;& �pG��ex.}��������E1B7j<�Y�>o)����ڑ<��r+#hO�C�*ބ�{�dԬ��p'*<*�P`H%�s��a��졽�o��3^�}���&���𼎆ܞ]�\�@{���6�)��%Ȳ�7�9b�ǽ��D���4����y=���v��-����rֲ$�'�ɠ����>,�g�7���i�3MB\�OU	Į��õ�R�������&�+�Ts_}fd��w)mП�6����luZ*XAekw���7��KYv�l���O�����A��C��M�3C.F�y����8\�]L-*���1k���>�r�������Nmε)j��V�Q��:켛+ô���yySMIM4SAR$���7>{��|����q���k/^/6����V#�aϓ�T����)�v(.�Y���P�z������]	�/�x�`Z�����9��ɳCh(�b,t9����%鳿�Y�'������s�� <�L�<�}=B ���<2ǂ�S�`y�@��И�`HlD��ۙ�؉���޼����;2���׷�l��֟lB	�1,��Ji��Q�T���|�9�=�;��/�r����+Bá� =C!/	��]F0��MBǓ���x.��ƒ4��׾6/�����.��f=*���}*L?[�@���;W�:�\k7Ӯ�F���k�wM��s{�S�T\Mjv;1u6�L�@{p��`YQi���=�l#�(�"m	�~܀���.ۏ̥�!;M}R�un�R������{��M'y�m�a=��y��B
���A�<2���D��1�𒢓B�+�L\C�S�����P�r�����.�c����<æ�5S�T�����bЋy+�"�gв���qKcy�y�ϤU#^{Z��Ѻ���rc(Ij���糧��kޙ�^��.Dd\�A˷y.��gѨ����:�:L0��ՙ��$�넝ݙKL�B��є4�v����V�1��&.`j�8��Q���c)=�$-���I��הk.u�c�:�)�xU�ݪ�̘�7��gj�7�����t�s���H%�"�T�.���y��Fʾ�We��V��ZGʆ+0��{��dUA݀�F���r��u���%f�Zp�K���b�;Wr������oo-��L�8�.��ul���F�~�e(����)�k�FZE��A�p�G�xP����\��<SbU�د6=B�ͳ;�
�Nn�3n"��S:����ԆK���˗�ז���R�4�pZ��B��j+#\�s�����!D��5��6��T&��e�n���J�)^�Y	c0%WLk�����6k�c�$�c�0�e�N�l�FgnګWS�%/;��]�5��-tZ�Hj��;�N�Y�{;j	-�]&�3�b��qd: ��v��ݚ����QM��k��}2��*��if=���/:�h�§P�g&��٢�bEJ�2���B�r�|���q���V'	W;X5�C�3�uL˫�|��X.��ܫ�u!�U5�&���Jʴ�b����v.g5�N���nr	 wKog�a�ı�Ѧ�B�����ԥ�Sn��[Gf�q�䈖����)wavA+��|�:y	)kz��D5�F�
��N��b.B���q�{q�a�h�$�{n��Օz��(t�},�i��et�������s�q<K���֤�����y:�0�w37xF`��aE�����X�g�&�i�Qi����Kx]1T�ES)�$]����Gd��>��[�j1�����M���V�U�u%W���Q8��{.��"a�Jv�oc�נꖶa��,�9��M�[`�k���s[杉���N�T�vi'������ͼ#R�+���W�e��2�A�UX%M�-W��a�%b��kRw�!V���+K�Y7��ԧû�f[��q��uz��	�X�z�Κbkp�>���9�ga�](�N�,��;�hT.�#ٗ�G]��T���{�'}�m�5�r�}(�Jk��z��0hv����nqoU�@,e,z�.J6�:���vآ�k���f��C-nD��7tP�#Q�͜w�`CU������"26YP�jb�I{T�%u���Q�5��g�pFjb5xb�����<����hTґ�y1el���˅˼���ԭ�����"��0�!;&ԓ�Ƽ���'B[	F%�@�@�V��5�.��p���&�f>$�{�`����|iu!�q��V6>�T4.�ݦ�����m%���.�:n���p��)V�WK�R��#��k{s���A$�Ÿ��ʊ���\�ޗը���BF1�����x��Ǐ�~o��k�F�A�̃��nh���3v��o�����<x��Ǐ�2�!$$��	#�& ZL�.Ili�q��x��Ǐ=z��- R&��F'���EL��I:i��8�ǯo{����{�����Ƿ �J� >u���wPD[ӫ�ݔ�HiE��
B�����ی�:�4d�)3ӊdP�%a�HW+���"Cc�ѯ���1�x�(��	��ɀ$���4%��	&g.���WD�Ws�n�0L߫�BF0I0�珑�<z���r6bI�C!�$~"
l�O�`��s�b&��U���
ě�3��X��ծ;�ѹ����r&Jݦ�=���ȉt��iߊ���#3 )����&��P���F9�8㑨!ed�"� �M�C�)�Q3\�T�ER�NP�F�h�q0āD�eb�P�.��7\n�]�v�۹-J����	A�w�4��U�TU���s�v�{�g��K���^��n^w��r����߁���xbٖgtO0��G������@(�ܟ��So�IN �^�9�U�^���}B�p�1gv�_,�y���tK�$t�&���E�Q�#=�7[�g��/��5�;���7���v���gunn`J��/��lw<Ƀ�9��]��&:j�#N��T�rf�m"?o�h��Ȭ{���"L~g��\xt���9��e�q����n��m��D�+8�W��Pi�F]�'־p(r�����,>b��ջ9�\��Ğ%vgn䐸�j�!qLn��7*dԓ�}�u/�'ug�d3����,(�+&��{�z���N���C��vn3t\�Gsz|k�^�	� �iF���c����9dGrtl��rtV��� ����=s�&��1�����䴄r+������״�z*s����]Bqf'��xן�!(T�������c�n�ވ���Q�Oj���R�;Z�we!J6Qqw c	܋h5ӌ��u�xTa�q�{�]-�� /*u�r���\i�E<֢��V{A�yMݗS��:�1����P���v[�D�������d�=f�f^������F_���7�T�s&�>O�*���X�6ؗ�RM˫�0�F�I��g�J�n,���D�-�9)�8�5�"����h*Hi�)��+i� �

Y���Wk=�s�;(���h��W�>�����w @AF4�T����oqSU�g�{xwq��ۆ]�f4��,y��>b��<�~m�����
jw�ؿ	:|��k�H�7��>�iĞ;��5�k��k�$��:�C��ơ����0ٍx�f�D�q[��N��hB���d�k{�ES��C\�y\V�(�مZ��3~�W�)>57rs
��>=����掻�p��p|e����n�&2�2)W���q^'�k�PK�"� T��y'�z��0�/��I���ϟ
���sƤF��4A>t���O<�v�Dn�&I�ef�����ܤ�=v���}�|~0���|Q^ ������~�fKү�9��|��,�n�@���	�nǠL:"����3�g=;��hS�����N�&O{U��+�s�<%N����"r�Ӻ���|x����+bÚɨ�~�1!�^9����0O(s�7�}�����*�p�(��s��/`׌XK$!�ϛn2���-t��cέ������>DTtF�����%?�b��ብ��%��1{ʒ��t7�AY_Y��{-�'�z';��ȯy���30p�ﶚ���4U��qͽ{j�qyw�Q���ܦ�=C���B��Iu��:�',싍��{���i* ƚZ�F���
F�Q�""� ,���\��>|�+G#]�d���^Y��#�@A�8{���Dn*�#>�Pe��4��hlM����͇*ɽ�s#9^8t,�0�.b��^Y��@�������R|eY��	��
�==u���T�]�F:���_ݸ�P���A}����p��F���%�$H�pf�fO{�L�𳣳܋4�H�M'Y�&��`FNc�S ��!��i�8�����r gX*���I�p�l�.��t��}���3��zP�KέI�¼��)�ٕ)�<��浙�Z�|��s!�y�Lk
i���'�+�5���T��9�b����v9l�}�Q��<�d�HA��T0�i�c�,S�R:�/�^zd3��PI�/O���e��PL���b�=�����2Xm	���l�:'������� ��oRw�A~ˈ���E���[���������π�A���U31�N�Q��^ ���p���<����U�O��]M�E�8��X"zN�����yN1T�8�����
$�b��$S�߿'n�O��(C���J�5[d���i�Cr���wz�)=ZF,�f��r��OF��Bj& Nru��~�5𙷈��Fe;���A6��"KS��q+Z��F����N�o.��zo"5�{S2*�|x���'0�r���-:�
�� G�R�h��Ti�P���H� ��ߧϝ>k|~;`���nlF��1�S�3�������L;T"$ �K]��j�-m®6˨{d^��_7 3fnJO�^=-m��A�O>hMC�7碦'y罾��|n^�]o6s8m�4�`{a��q"$��C�cW��c�9�[i�t��,>z���ې�;$��u���(�[P�Cf�O�$I�tИ�?{҅Bp����[ү�c��_����<�Ǎ����[��E�����,���P =ŧ7'��t2��~���i�ԝ�ǖ���ۍ���)8;a�jq����p)�=aŴX|F(FG�@���u�9�#�q���7��S��DJk�2bD��WN��O�� �o [�3 �P�e칽�ͭ�YaC	B }�W�mAqZbY'��
i��F�R�O;�sS:}0����u�dNJ���`,wW^�s	�qt&6��K�o�����oJxLK�E@�䑤���q�7=>�B�s����Wޘ6&<�zF5IR'���(�`��u�oJ���b��Ӫ$-�#�#/�mv{����΀�u��w.j��!�����UgT��F+�8p8˗!�x��D&B��y��F��/��P�K����G�ϻA	���Y<V菹�y�5}t�m��gnmn�c��aH�ﭼ��*n�b0�n��,Q���C����~�J��i)���hU*�jm�Z���TUcX����L�⮓z6��r^	��ک�A;U����T����cN`�9¯�U�9���S�y���
3�%�㮥��=z��8�|��<���r ���c9���G4�瑧bXg��?��:�E8���]���ӌs6D�jO<7��La�Λ��]�s�;W�}y|���\�
��$E9վ��BdJ{��`F�&�S��kz��c��x(���J�W��sH�}������ C�s���c�}�l֑��>�{�G��ߖ����Gç�?Uy?Cw�Ѭ����S�
�8Bv�v�ƝݚDL�)�T>5��.|�q_�b{��%�@�Dw܄��Q�|���s�r�3������;�ggZ ���=B&}��]B��V!J�`��U*�r�9�W}��}ڢ]{L3&�`�4�	C��;���I��3�1�?�*j���*��7�ƛ]��6f#��Ňн�'�a�yt�y��֞���+(O����T<%�����oV�$�+1���ԥ��	��ȫm�djq|�7ZN2�k	)"�m�����s�� �eZb�@{�Y�K�*�������U���:��2m��|nq�@�Q�I�E[��F�|j�Q
�SH�ɟ�O��.`?�����H�3��ܸV3s^�"7��誡�U����.�s%���Ô��Ɯ
�(�tqaw�ZVU)�n"<������/Y��ҏ�	X�2�I�-��u[��kf��Z�$D�4�AIRy}�9]���|(Dc�=Ϯ�ۂ��Ս .��[�NV@�4Q�g �S���6C���M���������k=a��F�/���,��V�w�+�?cAz���H�˯-�l�%n�� r&&#�#˕�W9Sb���l�SzB�#(L$�n�G6g�~U�nWWLQ�ٱ���V9j��8� �RS����7"�T:q�!��:N&�T�����OW1�-��ﳽ�*S�ͼ�7�֑<� Я>�s�]<~�a����G����\���%�J���h����'Զ��^Ԥ��)�x��3��`�Ņέ�|��)���Rg3޺YV����y����Љ���,A3�忟�̉�Τ«��y�<�fe�T4���{��k��V�#����xva�0~lD@���/)�������E�Z��3t�{��&�-�5�"BU����0����X0d|n	�?0�
ƶg�Ȥ�\���Ӓf�TL��ܟM]�����N�0������`0 y����y�]G<��0�/Z���|t2:c�(r�*{3Sx��&�N��e֗�C�a��zn��D�j�41�4p���������`ٵK	m�#4PF�pe��ܳ��*V�9P��sL7�U�t76�1N�ü'-�'r���2������$�v�/<�� ��1��*"�i�D��"	hJ����Ȭ��(ȀȂ*���|�!�W_?�����=�;@��vb���f�ƈL!�2ߑھO0r�VJ�Lg=�6�us�16�L3z��\H��-�{�[9y�K� ��'�ť��1���lx�%K7��*MYu��������Ϲ��hvf�I�w��6k�����'���?���"�ȯ���I�[�d'� P�wF��r�������
���mj�u1]�Y��T̃9}\B���&��7ĉ�@�-��#l*��z�)��=��{�O�Ӌ	��}+7�>��Lȟf���s�J1#�Y&C� P����W��,,K�j���4�SաSZ �>^� �����w8N$��<:Y���y ���ГK�D]�S����1x��s~tfD����J`���Ux]���,�cЋ�t 2m����j ����b��k�xS �ͨO�ϳbs��%�{���%L9�+�5�Bw�l¸2^�Y�W��ȱ�Ɇ@��A`Za�2=e��y�ހ(�L,r�E�x�4ޠ�oM��@�w��������I_�Q�5K�U��id�T
��h�$��I�>PpI������B�6�][�hD��������'aUD� ��rF��F�����}V��w�W(��W�ʐ}���M��*�#|N��n�c�Y<ok�r�f�Z��\o����=�����嵒��ۭr�ڍj)�usmE�5�nݵ�[h֬Z��ml[Fբ�H���
$�(v��_>|�������w�ޚ1�^"Sm�����D���'q=�z^�ŧ�Y���:��4�ȕE�&�-j]�`��g�S(p�m����p OG�:Fy�AɟF�r1X��
�vu�D��%2	�y��ѳg��ܿ/�&Y�9�J���"|�����,��, �j�	��}������aC���eA/r��0yD��ض;�9C�y����+R�mSi��;23���~�������S����=�{8"a�ʄB�p��0 [E/$����A��S�O��!����B�s�:��1Ƀ��voOgk�0񫿾�3��WG;�Dų������x�� �y���,��Ak)%�v��#�Ɨ/��/wYS7f�vC�H芇U�,��W�ZP���M^J0S�=���]�'t�t�B\�Vb|��;Jw���PZՎ�wO3a3�Sg��+v�ėa>��!�0��7b�fk�+2�wr�㿏��	M�-A#��g�Ƕu t��D8am@Xt\���D����Yf�P�W�I0a���ڛ�H�ǌw`R�6�_8\�2���9�ȷ�,}wsu�z	6ŹS�(L��G>�_S����u���gee6���F��A���RN��Z�>�^v7����9�t}���y��u�\�k��Ё��<>  `��iZ�Ȫ2 F� ���i�j(!h@* �
�� �  �!"0B ����z;���U�e���z���f�b����T���͑x�����ez���%5ޙA�,x��u�׫|��x/V���FC�1fG*@�B���?S�ε��U���S���%�tɦO����n�fL$=�О�w���*��Hk�qs>=�q��Cc<�ο�T�a�8O�{;�%���0%�on6�N��c&�'��v�ƶQ�"VEÚ�G���(�JzG�{9!�z�_裐^J���Ie;�e�9�5��W#<Û�LYz��׶
`���M����N�D�UƙUgGR��,��v^�n��LZ�G-O"�}��F�;4ø�4tמi���F�eV�gK���OZ�J���LKeZ�BԮx�2z*;��㸏�x�S�0<d)I>�F{b�k٣ԧ� 8� �d����n�5߻�'�]<^l+�@�Z�q �٨>��u��p�����uN%�~@������(<��P�PloX�9�!�yN���c�?f[��R���	�7H����,�q�.�;l�`��� 鹪�.��E�"�Rp���D���g�MU�8K�$̛ԡޙR�u��Ԛ��}2e�Cw:��s����b�^c��bj�v ��5 hX.C�gr��ޞ9�	���[m?��$��O
n�o`��Ld�U���n�lF�nV3k���)������˥J�ʵS���Ib����Tu��"#�j# �H*G�ЂTH�@@@#M �@�4
TFDj��-EU�j�֊�ׇ���k�f���z���o�1����#���#��q^�a2��=0%C'|ϯo�Ȯzr�5�:[�/�ǘ<L�B�o�'J�$���0�yB�<�ce��S=�e��W��XaQū~y��Hdy��К�l��VzBC7�Ӷ75'��o
�C6�ޗ|�O	��i9aC��-�d�zf��m3��Rq`gAYr�{��/�C1��e��v�9Zb����E�_�("��Av��TEy۞n뙶�����~��+�H�W�ZΉ�o�d.�ǥ3]��l�y�D��tt�����1s�����g񳅋��y���x�UlI���>9;�4�17���k�#�����-Ԡ�O�-�
��&y���If��Ր����D�W>Ɩ�Z�˖��(bTz�AN-�-���B�a>ip�Н'C,���M?���7��^v���]�d������\hS�W=#1�{vxz�5�,mk�;}~{�<���*` ^mט	n��N�}RS��Ⱥ��e����yܿ2�'+`mTי�|Æ,�>2�;�j�V���UM֠y��u�r��P�����i&Uk5�]S�f�9t��eS��3n��l�Q��6���T4SL�s{`U��0�t	��N���Ob0a/]���*m���V,͙J����N�sXb̭�3Xb�]Q�6>0N2�4gVu�m^'X�Y�:9�9s�t52-�gt�9E�Qf>�f�"����wX��@me_\��.��Yq{��7�'/rljX�<�����K��Sʬ�t�*�ս[��db��i�s��²�%�/7��^�l�7f�����FxU��ot���e��m�ݓ�,Z!'XPn���}Ӳ��Z�r��V��F���w8R��oNΚW3�L�AȺ�z-�mY�w�.3Z��ee��*�lwa�\!�0�ͭof�s����ڗn�-a(�63:��o�׽.�_�ȩ\��aZ�q�n,�啈�u���V�����e7��6�+54/��ٴ���l���j^�0s�QWnoN�.�V�쒲�X�ҡ��W�[x:pw+s	�=�u�S�ܵ��5*5ۻ���TVd��`��o���
��=��m��k�7x,��*�ul�e��z�����y��u�%�8v��0�*���vR��e\��
����dL��z�4���%qý��|,��QEW]��x�P�o��i�i���(O�?c|�gض��b⼽��[�B�����qY�10TޯW`�8��jXּZ)�1��Xp��ꗸx��R��g��$<8$�*�ex�2�MZ7]Tt�cA��m0��G-qVM&��τf�:��B{\�NVΖ/[�8�\�F}�X�T�&�[8F��yO�Î�d��P�}��x�]����u㇄�ow�M�,��ӔkU$nKtv�w��2�RJ�9|�=�}��]>�b\�U�2�µ�v	�,l%Hv��z۵,u tlu�ͥ=q�+�S�ƝYҪQ
�x8݋|x[xy�u���P�3&J��'Kz-)��:4K�30D��HؼP�a^Ú��Z��Tc͙�K�y�ʢM�[E�D#IY�Cs5]q��+���Y&��VZ�"w�6��Z��Ŭ&7ws!��U/�s�1#�AEqѡ{�(W\��M.��bk��T(#'�� ��v�B�n��p��dS�U+�^��l�cD�Ì�Iݵ:�5�P�?�i�Ѵ�B�D�;Fh�k�-۹���<��ƕ遊[8�T�\.�!�̥d��n�
�X,�A8��M��$�Q��j���-S��a	ě��)��4�,(%�VIãV�Gr�b��ZU4乏����{{v����R,���X�X�$T�P��1Y�VE�j��e�[{��0�s�^��r�A4���[(�7�L���lAPSFda�1��/")f��C�T��B�TET�@�c�v7�Cj�J�i�OqD?���~=hw\�Qd4�P̢@^�܄�	 @��}v�Ǐx��Ǐ=z��L)��ivĦ��l�B'uuz�f۷�����=x��Ǐ=z����2u0��ü���b�Ȓ��dj-H�:iӎ8��}�{����{����J%��J=ҹ#2�]�OJ�$RI!#t��8��׏o{������"Td�i�DF0$(�h"�݉U��2��wb,(|n�\P�iO�,�0���6N둈 |n�l�)�$A��d�(!b��f�l�f���N R�z�0�I! �;��Q#4D�Q�D���瞽~w���FQ,�1�N�U��:���UK�R�cP/BYd��r6���ۜ��&R����V:�ѷ}9VM	@2 �#��ٿ��W*+Q�5Tݺ�nm�ݻZ�mi�uV�+X�֊���lj��k3� ����#
q;���;~`p|�z,p��ӯ�N���k�$�ν��z}(���O%r¢n�7���n�据�Z��×�p���bD�M���]d����.+}�QaB�O1�r�TY�ێ���f��&(u�3X�s�֟'��D�4-5��4 C��z����3�.�Hڈ�({�e��Yn��_�������.�ȒW�>��Cɛ���B�D�,~�1���9	�%�w�{��w�ϯԅ�P����O�X��'��~&�7��%�<<����A��0���]m��}/���Ր�	��8%�>\~6�b��c�^'="A�ǜS9|�R[m���^�{��Z!�2�xSCע+��R��kD '(�D��v7��G.����Vͱ3.LBY��5ՙ�<�)@'�6E��%Ͻi��C7y�-z��BKܩ��f~��sI۸f�^dbm�PS#^Y�
S�)��3P%���_yz�º�Z�S�z�����:nw/|�~Ƈ���1Y��0��)��
L8�yOl�����uܿU�N��.�q8-�14�/ɼ��-,��WTJ��nS�Ϡ���*U��}n��®�5͑���<B.���MUVS�Lo3
Vh�7nbp�S���P�n,ʝ�t]��δ��UW* 0f֒����ݡv��A�W� Wo٥ �� ƚ��",����B��i���2" ��xa��|��&���v����#�R�]���h.|Ǧ��C��u��O�l!���uO%��z�Iz�/��}��G���2P�ݏ�)�j���o�=k���Rb}7������K���h���@�`�57[��>��f}����<HSި�4Q�KM�����͏��)���5���\���}��2��B�_f�a��Ӧ��]`�Ls�A�6�a:w9�q�F7]5p���M  ���&���M��[泂�z m��A��	�4�V�^����l"�0Yr3���h`>�h�G�:l`&���Mt�,
pT��ѣZz=V�n������^~CQK}}/���8C��cg��Rc�{`l-7��G?0��������%n�wc�YE�k*dKl�]�q{�W=�l�* ��U1�t�xt�`0d:]_e��Vk�Wj���L�0I�]ƽ�V�<j|��}:�_�Ͼ5�i�A����y&�ݪO�:&x���a?�ܑ㜲#��-��e��-���,Hq�x״����y�Q�û���F��pCxP�A���O�\��t����]�8b��ޫ��b*��T�'g4�nJ��5͓^]�n��i�m��K/*�Ҏ]�������{��U�ҷM�(�s�孍�73z=�����H��iA��iD�2v�sV�۪�-�ڣXִ� ȀH�*C��z��Q�.#z�^On�L���J�P�R-|� ]<�i?x���`n���_����d&��'�b�y]oi��ѱ�+���[�V|�n�/*Y��G�x옷([�|���˝xg��h�q͞���=K�=e��Ԟ,��5gF�]W�)�\E�C�l��W�v)Ě���馓l�H�소Ni���}�u��t��t-�oOy�>B��`[R;A��^����|g�*��x��[ON�#��rΎZs��_ІE�ͯnW��	M{�ex2jY^�����yi���\E�z6Kfm���5k�>6GW�,�H�S"S�`����o�/��$��B2.>C�=�Ȣ�\mu���U�KP��Z�(�P�&�N�htW�Zଅ���1ӟBd_�ཾ�6hU�棫� �O��'}���+/��>YhPꋇ\�� ��cT������XJ���p��d��EFmE��a�h�Y�2��7��������E�\Ú�1e��<�l!��%7_���5��~�m�;���Z|B��d;!��_��~D'��8��m�a~��"�S, �����x)�rɄ&� ҊM�^�vn������e��"��VM���;b�&��Df+�4Cƺr&�!Lv�]���J�U�őDn�`D��qO:ѧuou��D���a��b���[v�V��.4���q��-NU.��*��vy������Os�7�s��7�*��� ��hE��V涛�WJ�&�U7n�nh�cj-�Ҩ�-�� $�	�$�d���g~W��u����xd^��[��С}�(�M��_u�	��@/�5흃d�����Z�r��n��`�]B�3wD_�u։�-O�<՞�̺8��� j�e�Y\�R-��{�\�m��7�\S0d~aI�C�t^���M���n���Z�8���DR9�}���[Z��z��q�Єhb �
�L<�ڨ�r���d�Ж��aQ�xo9S^�R�i��@q��u���QSC��
J߯�2@�આ��x�Z_���25N �Ь�B�LJza�y���0��oP���]"]�`�:.B���KB�ev��l���>�޽��Z�{=r�ef�/E@A��K�mjO�ͼ��f�W��*���*��u��{��
�M�O~��SC)t�e�p�9kK&�P+�h5͛e��H�6ڴ�7�ֲ�f�3!��׹��7�Ǆ��0|Ǧ����I��!NB�Ǣo%ⵛJ�۾L��
���6�E�T?P��P70D�\`;>S���R���GL�����Q�̋�ǘ�z��֞Xh�D�u���Ӓ��4$�j���L�̒���ngN\k��UqH�3KG39��3y{��D��ױ��l�
�M㴊F�	��G/mk��s�t��$ޭ\UL����n���P#�ҕ 	�4;��v�j��֭\֢�{�ޣd�Ja]�kh�f�R��D̖�� cWQp�Ol���(2.�0��fi�0�ܬDg�<�s*����>L-�<�+(*�%8�2q��5�{�Z�ƀ��l����5�/2
�J�uR�܆ƶ��y�>k�In �̕�y^�W���A�Nc߭�[������A�5�Tr��(B�P�_��|��kz��׵<�=~�6ȯC`m�ZF.i@��>��D��G�MZ";c�<:���ێ���Q�h_P�O���lrך������'I����zݰy0��s�}�a���>�!l>����zu��Kץ�:��o7_G�U:U�K{���=t�V�����Ux,\El3��D��D�B��no
p�[�J�g�0��P֧#���y�|>7L��F㑋����*��{�����ث��6A#�dp�{HyN�-�rxnE%!Y��<:o��2���d�#� 6���K�3��Y݁�)��¯t�g�,Hwۭx���D�n˳�U��i��3f��d�I�oD��a��E0 ��cC�[9}��U^������1H֋{�N���H���l�}9�G�K++?:�ݙ�s��eD3�} �{HUj�bj���@:�@t%�A	'F*(���iK¡^��J�vΠ�.p�e��k�SQ9�ջ�X{u'�f�Ů��cy�9Z����H�4СM4�d�4�EI!�dA�@�u��o����;U�?1������d(���@�H@U�J2�����8���5�SR�̽4Sj"X$>���mtg(��qqp�i�p̄��y;�݊==}[����۸;S/6$����k�_9�V��S�~�����!��<�X����Sf�wn�Z��_F��F�`٣6oP�W��,�Lp��l7�1P�^Yµ�&�O".=A��}�{q�g�o^������+�8��K]�d�b�)�Wj�蛸A�q&�3G�K �dZOx���WU�Y6miw�s��"�5�Ȃ�4ħEB`��EP�Ȼ�F�������lܕIj�*��x4��4��[��q����gٱ��x�)�j�bQ�����=�=Jqc�5˪��3�DK�����G0�v���]!H����]0�ʥQy��z�0��Չ���(n�J9j͑!����Q�r!6צ6��7ҝ�g]eE9���yQo٨9���tF7�m�K����L?2a`��h�C���zQ_/��\
K1	U6�D/hB4oW�W�TڛY4�D�̪����M��r�q��i;5�ʇm�����׫�*l+~�×{ɓ�s�z�xBȌ!���}�9oηj����[!ʪ���]��r���3J��Quk�CQ+;�p"�����S7���(�wUQ����S��_��Q�ƚR���+v�ch4U��F��������w�/)L&���6��R�wSVF��$��l��+6�2�P>D~��wdW�F
2�*5�P*�s�q��}�ٚP���_T���v���s�GՇ��hQN޵2��>}�N�&��d>��C�~r'�P�2Y�Y@�{�r���aMU,%�X���y�d����o\��u�*��g����w�T��.�64��\uZ��{C�b��f콇x��_��=���D���� �?[������sRJɞ����1QS���=��C��DW����v��}C���q1*l��|i�Y4�Q�L'��\��;H(�m�uc����պ`w�5��<p8��̨~��Ԙ4�i���'�z�����w�ޛ�eS�<5V�G�j�Vd�w��C��QhO^��W�KL�P��C� i!@��R�8�9��R�Xc�J�Qo�c��ȶ���&��P��ʇ��`Z��x퇍�O�c�zE;�&�#)��c'�2g�5�[/`}�|�G�=�+�|�)�L ɈY^�����I��7S/k�x���y���S�����6͈�1�V@R,�W5�A8��ܝ#�F��-Ѫ!:>1�������1�Z�+Q��MU�I7�;&�S��UUe
z��%YZ"'�29ܭ��k�w�c��)0*�,�|a����Y��<�-x&���{��%ް\+�����"bL9F�dE��;��E��1�ݺYW¯$���?MT	4Ѕ4ҕ45	$YBk���9���o_	k�Y���PR����W�]���+�M�8�Bb^tw0Y/P���b��k�~=��`KZ(�kgۏ�p�<��cސ�ƃ>?[�#ۦ,ur�.���SYڋ�V�Ѿ��(׊�a�^&,������	��t[�#�>���ȶ����f�m���M:�u��;�YK������sN.iz%���l5p5��&f��~Ua�3�p�!�vI�m�z�U�\�fc�*;���{b%�C�,��pK/cV���c��4�Լæ&���u^� ��~��r���x��W>�9��ԛj��o%�A�[؆��*��$A�� �bH�گ�>_�/�4�>���u@\F�ӥ�&�`�h�Y��Yw}��[�|�+b��~C'dT0g���Ani�>2/R�&̌M6c�i���{�'���#�|̅9�aD�4��䨴�O�ۦ�_������<��4(�`�˞&s�cݪ�y���R�*�6<Z�^��b�����f� hz�q�(�3�`�#Č�[r���2L<b�1�rn#�g RO �jڌ��׮Ee#٤�(������Ȣ�(yx.�λ�LR{h�T$�rSr�S��Z�c���-,�茋�x�1N:��T�\���Ĥ��f$���Y��q�<{�G��w櫢����症�����v��Wnֹa�-�@׼�](N���[���Mz��쫣Bk6Qz@A�ܺ]��֞��q&r^�D�F�}��={��"<(e����d�t��QEsN��|�8�!�d1V"4���%�V��ko�Hf6(d(�zD�詆����B�=o+�ғ�`���b���e�р�	��$�")
i^k=1�o[O�⦿j�����A�r��,�_����b!��v����䆘�\�P�����;�W���%�#��՜{��Y���w��Y
�N��ѽ��^��T�q�9C!\k&���ι�z"m0����*�UސH�d�s�o�Q���LP}\�A�
9����Q.�n�-���2ͅI�s�2�s@��
�B��Wf�xa7���7sU��EۖrH�֘t���s�8�RwS������7��x`�HM�Z5�m��M�b����s*3������?��?%E�Y-�*~:�D�^! ��bJ��.��m��rl���"�=�/ܵ�w�%^����{y�T	�J�ϣМ�s}>�6�v�	��)�d�S�+��}N��{{ȩ|��Ѱ�3�sI�j2�{)�Ȑ��� ��mޕ2mU�m��16G6����i��b�X=U�� �[&r.�UfF�ջI9G���3;1Pm�o*�)����oj�(����M����������hi���eH$�(o���w�>jwW�,�{:z� �����\�l!r�1�@��㪗�,�ޢ�	� c*<4���y�{�鐢��5�	�X�T��*+��ܳ��mv�L�0��G᫋Ϸ���
�;�#�T-_� ��xL��R�����:�_��׳�H�����1=�̎���{I������xf̬���H�)�<B�70�S�ע!���v'�>�zԑ�"G`�=$�gdt�=z��Vј��êyw�
y�w>y�����<�\@ϴ�EA9~��Zؕf5:ˬ��L�6�t9��h9�yev��/�>b~
�G��ߓ2�7j˫r�y�n�λi�NҬW�M6�i�d����!
��^i��u.�
���9�=���I��Kʴ�%�w�{^k��S�F�(<5i܁L����'�ë������T9ז{B'�m6sGI���Y�`�|�s�cn!��f�)�Ɛ$&�� ���7p���M(f���)��*�#M�E�`8��q�aO�jO��Dsf�'H)�jo*b'-ׇ���x ��/Z�Պ�C�[m#��#���94^��t��t�d�e�k{T.�U.����6�z�r	Ҿ����e�g�_�bT*�������;��{O���w^��H��˱����Tf�w�ެ�x�v�Y�Qa�rMu��˟jq�W9�՘r����,�ЗP^��|%5[w�u�D�_p銹�3�z#}
��Z������5��TȈ$�X�Y#���F�7q ���wO�H�Z�YuO�Y��sA簺��&!���zvp���jE\Kr����Ʋ=�YNK0��y��\�������8y�#霹����ΜR	�/1[f�5�	m��7��Y��5)�/.��YI�fL�qP4��i&���P�D&���4�aܖ��{8����ռ���Gn���iZ��+�<�pf�������)s�,���+�k����y���%��M��Xsw�*��b�CfEz�Bn���wLF���X9Y�PE�`N��XחN�m�NXےu3G.3i�
-���w���n�����z���P*��A�+V6��g�0���pι��� �K.��%z�%������Q猚���6����^'�.^�H�ZjNmY���ڏ_v��:�4����	�خ�)���ì$LT3j�*��\s�W0;U�^�S;T�s1f+��F��k�]N��0��7�e�$�/y��f]�@�����(�mK!����K�}�éZ#�2��.zt"�]O�6��f�jͨh�˽��`1�j���fɘ���%�6b3��&)�媠��vE���t�.�*z���{TFQ�'O'yr��Dm�2��2�tj9ks�]5rKIռ���5��H��Th���n��X{ee)��Q`�W�6�;��%$��'R��GB�C��B7e����[�*ڃ'6�U�q/{-ר=����rxA��ܠ�὾|\�OAy��M�h���\¡��Wd�5��p#���N�Wfؔ\%�%���W�b���ˣ���RؽvLo-�!�o�
�*��3�D��G;��q(�#i9s���{m�Q��c�f��3n�e&��Q�V�.�l]2҈���6�t0MԆ�[��Uu��i���j�ݶ�rKXJ(���w���nv����[Q�������e=w�f��}֑��Tu�����^\kjP�/�����P������aN07ٞ��^Ї���d����dt�,h���9�S}�.�+��[3K}�+L�d`����B*pn��b��djC�v�WZ���51vT�W����J���YVݼE���GQ�1ݼS�MG�M��Q��f̎�Ω(��/_CAծv�ba�kzw1��ےj��{XIl1FY�S��H\�{����߿?~WƘ�(��Q�)6
6"�b�H1�}q�Ǐ��<x����$�|�k�$$��/��2h�D�A���ӧq�<z��Ǜ�������!,_��d��n@ABb�E*2!q�v�Ǐ^<x��ǯ\{S�i�(bAQ$ى���F��?���q�����׏<x��ש��:ݐT"!"cA�u�	�I)�!��1Kκ�&CdH��F|n�D���R�1a�DE&M�˗g�\"T��&��$ɩ�"ACQI�$фьY,l��$������3��@�L�*d��"j��%E@��ǁ�c)ĜJD�HXi�u�4�4�JQ&'	��a�b�p4��Iז$��°���;�i�x�A������"q��l�9&�r�,d����|�M%�=w��R�$6����`�#NG�(�2y�݂ca����m�HhG�Kn	A�HIٔ�iHJ�L�\����0�h�Q&�p�"d�R������u������I#M��0ff}_/���.��m��g�����u��:����֓�ￔU/�Z�$�c��^�
8��e�Y�G�fQs��,S�yc���;T��y[ͣY���w���UtX�:S>"�e:/u����No��3�F�^V��Y�OҚ>{/�ҏ���5t��A(ׇ��E	�>)
��Ю6��a�R����.��e��IE������a���	�e{��б�;_����&��~�t���Hq��g�ܠ&9����+x�0�jE(�c����,t��2/���r�4z��l�����������)xn؁�7k�V�bJqޢ��Y���l�@�̀�Ai��F�ͬ�^$�}�x@�
W��E��Q���о�&\R�G�����W�U������q����t-2�T	��n�CF? �;�w�8�xtx:�ߡ���z]��2��f��E�G<zY9��3��E�O�D�Z^fK渏:��6{��<�|%���Xh�IM�c��	���L�%�$6P�j5�*J��ג:�m�����,�����q���T?c�:��ǃ_�����d���'_P.L\�~b��P�n��@�D�n�45[��\=Ӑ�:0:��T0�C�oSҐ�#\V��N�ٺ�9k�ʛ����n�.�.:�j7�*%��Xr0����to���7C�K��6w�,{�Eq�ӝ�/��W����1� �����<����7�8���f�z
߲�#_ ,p!u"�;�qt��b�1a��ԗ�05>_��˨Z��w�<��Q��.��;R�]�C ��`[@H������{gZ��؇0��q�rtF330fC!׬8t�7ι�ё�/��s��q��9D�L��x��a���Z �N����چ�x�f��a�؈�@Y`��z!	Q���[�ƶ1N����2�l�Y*Z�6D����s�9zkw��\\:afo�A�ɼ�\��GTymާR�>�o;5�Zu�1&%"��F�[X�ɖ�{�U��ŵz�"�.�Sj������=�����7�,��q%R��D r��E��sq1e��<���̂�aF黌��3\�xa�
�w��UJ:nnc��8�����O��"=aŕ���j�I0"��fB��"�Ʀ޵����<_�!g�T&{�R�^�|EP����̈Ne䨎�M��ڧ�<6�9�0�����no�u�C�;��<��t�hL��T��Kk��5����Y��������Uk�� �����uԵ�3]=�]\s��C��n�7�Tt�[6�JhA�IT�?(u(��l�QMJ���l�c�^|0&��'ez�Xg������lff�7.�7�7ޞ�cq�S�A��]7)���ZdVS���j�"/��5M0#(�$���N���Ϛ�^V���y��4���{]�83�y��Bo������pd�fF��7j����"�0n�%��U)��r�n%�hC��d��?ǩP�z|��z����؟
t�i"��s�o:W\r�~�a~�����Hg.����H_&Q�+ϤQ�����E��'���x	�*��Lbhd�Ǿ�#y�aۘ��;�����o9�Rk-������?��c�?��j@����Q~�#r�q�z����f�/EB���K��ִ�-3<"�Q�N�� /^)\�>x�`Tz@Bq�K�a��ꠥ��#A��#T�;���]��]\v���1�X21��b_�IO`���~��v��
�?s,���w[8��Hr���Vt�c#�T	tFy��ǉ����q"�*��;G���L|�s�|��K��rB�X�]�.�����vo/x���ǯv�s(Wʊ��i_ݎ��|�4��AŘ^[��E�c����̬�����`h�TccND&\�:"[ŕ��'PV�5�͐�\�>_mY���3�^��U��dn��#b�dco����B��w/�tc%G����JWA�5׆�9s�s��\��Q"z�p7:�X��|�A�U	$�7nj�c*L��r6.�e�tN���d*T�6�]�:�wJ}��
P��Υ�xP�{+�fG�B����XČs榽��g��>�+>^������7}0�>lҩ0=�	���}9����.��x떻�O�]�<�j� ���!ҿG_�@#�F8���x�rP�T����J {��vG�����c��S�7���'�H;rb���p;��D��l��C���vě� �����˭�u���
V�/T�W�~^�D��q�Q$w����?��28_��TL7�T�ڥ�(�$����pP*}�XZ��,�}J�����G=;Ƹ`��5�>���n���d�B��ƺ�uަ.(Ҷ�PK�X�b�å�j�G�'>"
�{8$�W��۷'N�9�&�)�_����(��Ot�y�!�W�Jc���r�mA��~��;2�H���}^����`8���q�����Ar1Ǘ#6k��'�������m�m���?Uy�_�YZ�(��|�:|�j~WH'e~�!"U�.^A��f�Gɍ?M��k��T�~�
�Pkn�?}�*$�0`���+��.}�U	�(8f�N�''��"���]F U�T%�K�60U�O��	����8�����=ۖ�gK��r���:
v3u|c=)� �q����x{f���_X2�V:�Fd�Խfb�}�)˫��07]РN�Ҩ�B��b��N����rU���#�1�ܲ��|�s���>�Wݢ�!��tBS�u��W���xv�q��B�԰w��t�:b��)��4���`D]�6e����[Kww;����G}�N<������"J��~۬��9�M`�bYd[bD�x��z���râ˥�	�|m�$;gg��a��	��*��v�=����o��6����e'��	�s�i�����V�b��P� �O6��u��q)�gEH���8u�=I�q᪳E�χݫ�e"��"��W�ߞH����g��]��t���bMlJ>n�E�K�em����楚�S�3�E��y��``\�&���]!_Aw���P8."����M4`mϑ��c�,���-�sh*0q�S�mxw����@~�a·ޢ���*4uʸhp3���$�нCJ�]�Gc�]O~��,��b�8�\W�P�$\C�g�&6�����y{2��ﰨ���2&���6*Qj��*��b����*�s�q͢��I��|S G�?�RQ�=����>�ýc��zߚ	}�dj,�����7��@X�W�ܧK产
�FFk;a7���܍�{c���/_Fu+R��KS"���#O��W*���b��a�{�j��t�ii>�k���DP&��Chb����"ޱX��Gv�2�k-�P�:2��\
�B����:�Ԙ�oN�ʛ�XA�޲�^H�@~����>>>:��}%�\�C�ن�@`��`BL�v�Mb� �㛎*��`s�Z��H����l5BE��K�my���#{S�x_�����L�?�(ֳ���_�P�@^[�4���T��o/_0�m{6�#8��� ���]���-��:�D>3��A��`t\<(�1��v���zġQ��2�P��a��W�A"�G������"}m�]C�~#?o���T��Dլ����0���T�Zz9��.�Mf�a<�AOC�>ٲ���髊8d���G�u��s�q�s,f֡�,�!���zM?w��L�!缆��%��D	S�P\�u�ދ݆�5����x��`��9����	w^���,>)�q���Z���zg<���-����Ş���m��۲8ҥ8m�!Ž[��=����Z��o��T@4�,��QaUp��yW\)Lu�Ɩv�O�L�w�/��ۢX�)P�
;&1�r�cD=R�������R�����*ȍ��t΅��DJ$_1�9t6 �WC��.��ƂF�;[��"@�x�u��`[L%#����2���?T���SV���3��v��:�0oB����/�n����N�仼Xj�A���tb	���ո��̃��H)�8��ъ�@�cZ��9�o{���Nh�f��w��cf��i�ȥ���Vp�[᪨�<f�ª6�c�a������'}�=�'h����"ԗx���I>xL��l].4�C�'�?FB8T�������Z7��x����������o쌭��/���v|���2��sP�R:�uz��N�җ�9	F-�]�-��h1�!��8�xn���W�1�1 �{^ؔQ>=0�y���Y�6�+t^On�&�P���c�~��t.�K��$W�\+����u�H�� [����g_Ȅ;d;3;��|A\�T��q=���:B@�lA=�!��ȹ����hF\�1�K8=��)00�1��ǧ�^2��M+喽�$vƳ�tR����~�E����Gr\cK�����6�����4½Šv׉���r��@�9�^ p�h��[������a�O�Ë9��f^� �͚�,oo�5y�+�p=s�S>�k쭉��Xr6��g�*v, �x|�ߜ}9��+���,�U�P��K�@A�ܺ]��Nt�jɕ;�dG��Ǻ"�R��L���gVAQg���(��s�<��O�:���Ԙs��m̉$�t%�ʐ�4ڒ�#g>�]��s�7*��ZcJ�K�B��Ք��%X�L8eӚ��Jg�5��?|}b�H���>!I7yC��U[���:t��u!������5
SX���nT�)�����ܸ��-��-�.�sB����Y�� ?x�����7�|���b��C�n����ܤ4�;)���,�ё���O��?�>���5r�(�K�L]�	,?y��lT�V8���	�,�ic�w��7�b��m����>B�_�MH�_7�D �����$-�~��EGG�R�tI�,T)_�W0�[ߌ��t�Cߩ���>BC�M��)�c=E_n/��
B5�7�CY"���G�������0
$0e�-MR�q��7���8��E�N]��� �G��*��K���Q'�H���}3eRc��d�s�0�F ƅi���ޝv�%��n%�t��i�c���P��˚����-@+z������yd]Wri:���ё�m��7�Ƀ�Q�����;L�YT�:�J�� 3>��
�}"v����ȫF�n���Cgb���4�}ێ�@�,k�}L�ި�q��7�H�R�y�?�3��7E�G#��r|�@��k�E*,*�����,�	�bb�l(�8A8E������5�h��V�k��3O�&)��?�H��'��;�*.���U�p�v:el9��d@��^s��LT�&V��D��Z6�]{ܚ�J��I�x�U��3��1�K�|�o��qvԆ��g������Pꃥ�-oK&�$-C
/��ͤ���n��U3��D��m6���]�-U@c�NZ�L��%�:���増�������q.�u:>���{�v\�Aݖ�RL���	_x��я�+⧒)~�*pZ�)��L�D�'hC�N���c�4�c�~U��䷲���^b 	 �|�ߚ�t����ٖ�ql<�����Ra\bS�0�q�5d^ζ�Bi�MDi�n�Ai-�`[:y��(4>��}�*Y�?��	�3��i.ۊ슼�L׵k���ћ.�p�>w1�NF���n�<`���|����g�@?ڙ��St���=�n�i
��x33*dtn���A1>�>o��ӛq�Թ��"�K�E�iA�qR�7կ��2����#k�=F�m�K���0��y�7���9t:��R$��]MO �"r�7��$�PR�,b��v�t��ɳ$7��H�צ̙+2#�ag(P=�T�ݘ�i�V����F%���4hm%ĵȈʟ�W,��=>y�A�[��i:��S�E�d�*UM��m>��?���������W;D�L����"�m���f=9�(�#;n��|�շ/���̗>��F)��&�<���s	�\9��-�0�����xLhcAt���NP}W���"j�N�
hPX����֑����]X�x�<cUa���i|^Z��ݟfqp"<(Y��4}�W�?�Ճ���N�NA�q����-�2+]�̓��W�S�^TCM�{Wef�f4�TSw:�"'g��y��o7���s,�9�K�b����@J.�7E1��W����v���ty��	�Ә VӶ�jxGw2�B۳�FQ�u��r���I��yt��G2apCu�E<_,�g��M�@�9^[��MOV<@w�l[2Q�ټ�)�kM�4.�ƕ�{��C�����@���@P�%����;jʤ��H��W���K`�]X��wU�,�F�WS��W9O�E�Ҹ���ȇ�0$�(�\�.�_�b��a��0g#�G�r^a�]4���ٱ���<��D�&��i���]+Z������μzIڑ-�νa�tU��3�:��5�~U��z�/��s�SLɟ*�H�x���#o���@iH���e{z��g�J<n�4����~`��f�����ۈ��s�����>[_[t�.CdZ�a9� �DC�S0��F/P�6C}���,'��Nf�F��3�����K(rՏS	�� ��
W��(o�Q��;0y/�٧zLꘃ��Ƚ�`��ݸ����!6h�H.�]O�~��
�~��UB��e�Jq�j�H�SD{�'���L_WX=.��vgE˳;	d��w-��(�*�����y/1�TyFB�f#u���n��:�P9���Z���U���ճ��S����U7�sz�h-�x��.���yBѳ�q��+��E]��j�L���-�V��f�yX�p%;�K��8m!���]�-�x_F�5��crv�L���wv�PS��a��_a���=��*^ރT�1"l�R�%�Z�u7(n�Ҫ��i+��14���Qz��:k~�q{sl_:[��,�V��ǳ�N��Re`.������l �e8�1��r깉F(��ay��S5������Nj� ����S�|+Bg�����D�O'v��l�T���*���P*�\��J���uBXǞW.��C����{(ίfl\��s���ɕ�a�6h�X�Y@�=���P��Z����r���(��=�˄-�J�-��3�
����7z���+�ׇ�]қeH���h��)�5���6�帶-�Wd����GK=�f@���z�v��b�[��r.qF�f���{E�aR�nN$�̥1���/5�F��E��ԃ�A̸�x�ܷsSE�oy}0p?I�#+��*�q-Ҋ�a�T�ДA�+����|^�e��k���I�J��;��J�Z̆�±-�&3���UZ9sw�/A��O�fk�{�%*k�5w�;���3u�Mg{�`�*ա�����\X�¡��:N9�^;52N����2���7#�4D]9�Ƥ�����tEC��rc(Nk��rmE�㌉2%
��^^����3tdi�d<�����e'�{�.�jbEM����Rݴ����́m�}5&��$�J�è�X6��-5��us�A,�_:��� �2�_^vsE�UPSi�3F��q^��Rl�C��WWX4��9��S���Ün,�ff�ٗ�c���8q�ӱ�:F&��J�,�7��O6��Ţ��}����{�qf�|u5.!��8U`�W[M��'�z�9�2�ң�lڗ1Zsrh�@�Y�b�>lʫ��U��8w:	h�B2X���^bj0v��*i���q�Y�K���@6�V�C����y���m��֪�[�zes��ӓ%���ܰ��]���DV�K2�/]^i۽�X���9�Ո�f����utx>�U*Uކ�)f�K5*������u�[#un���D�3p�i#Hq���h��?��J��C(Ԫ�45���j��ye�'Bl�j�q���&W�Öi�����Uw[zd
��"��.���֣��{�H`�D��'q��m�c	Y����ɭue��	���nV�,�n|�+C�,*@������`�����ˢ���K���B/q�Α��� �˽l�S�i�eeC�e�w��]i�5�A+5Z�URL������6�;x��J����+�9㕛.�OG�%A��3@��	H�
� H��>�z���ow��{����}�~�5P�B4@_��Q�@����CPi�qǏ=x�{����}�k�M��O}�DZ">���.�YI	$@�@�4�ێ8�Ǐ�}�{������H��&9\"1�F"�C&�"�(2 G��q�x��׏<x�����F5�`�%�V؍$h*Hэ��3�Z��i+��k{n���4�(�bƨ�6��1cZ7��j�Ƌ�]Q���ƍ)��TDh#[�w\S#�MF���*�6�zmr�^x��:����;V��J�L�FEj�y������J,є��.*ڨ"5�*h+p.����զq;xЭy�k�������1��瓙��t�!]�W��ܭd��*a�@�Lʏ�=,�{����ދ�����U�4��0���P�*�3�h�=���bw��o�������2�s�<��� �q9wG��$��Nk
w�/�m/`�5N�ҍ
�(��Ɓ�l������`@Y��,L&M&���X��*������g14jx#�G�_�"���Kw�&�w6����>�t:C;�i�;S��Ӿ����w3%�i�:��
��N�w�RN]�6����ŗ���U-1i�.*���Vu
GG��0���E���Z��}ő��Q�C)������#kk��K9������P���2���D��턡3�P�s��<2���z%���yX�]H�X̐�î��QHwl�Ԙ"��n��J�_$��I��Yd}�m�W�L5��͇��bY��w�C���Q���+jl\DHh�q�2/�����*��6�s���S��!��$��wf;�5w����3�	N���gՙ�F:P؝a3��8{�_%�Xk��}X��̂���n�y31���E1=!�U7R�K��[8���o\�]!�d?N�}���Ү�Z�;�6 i�[m^~�R����R[~�lD��R�b)ü����x����omf3154Uc�uA�a��+*��gbc�V$	�qr}���P3߼|�o7�����ˍ�Uj쨗�/B�b�v�C���s�@�B�F��i��q�t1'"L_F]?T��0�f���:�ߞE�f�o[r��ce���H��\�0�� �fw�n:z��.=����������o�ߖc����-�S~/31r���Ǟ�M�oT&d[�gG]�iE��a;csW:���L}c�U	dL9g���� #��,�Ӄ9ιNm[ꍎ�]�T����"~��y(��b����!܍`����'�W��¢�gZL��ͨ�=�eI�a��WFNF6k�O� D��	�z1�������j� xz�6~*Ԅ�I�4�n�=�k��m�����ё)����ޅ.^�����2)Dv:��
b�1B�۾��c�8�y��E-�B���S	T�cKȷ#�	���M���N��	�qqHɌq�B��}���VF�]Ҷޒ���Z9d��L3e�3�����{3e7�1�����y_Rn/7&58Yt��/�-�e��y3۰#��K3�'o��pscdT{��WO�T�w5a������g"j���1�BYL^W��:��]��Ty$svL���=�޾Tz�o{'!���Q=78ln8�7{����<(�]��k�8��'.����T3Q9x&ۛ�P�R,M��In�#I�"U$އv`Vڒ�9G~:����=�}G��GڇH�B�N��q�3J��{�9�F�]i)ܫKF�[[�s�eqsH���zs���;�BW�X�9Ϯ'��zŲ-7����3���7���Xr�:xjnQ{	AcK�A�4��1�Q!�������.��+I�����w&1j-��:�qq[�Q!|��@}��z��/�C8kaDN@ ��3m�2m��O0z>�����`��,*�T�<\P'�k��4'��ڷT&d��pw�c�`�Z�{���'q	�(/~IA��h��櫘'��J�_���+����[�~l��g���k��mzv��l��Ǡ�łhW��A�b!���˅����nڢ·�K��I���WY��2�f�_.��;���ŕ򃟜j~0ƅ�)�<��訶G=����2�2m�b�=�;���,#�
z�7����c��^)�3X@���f`E�O4��1�D�򻇻s���ϜBs}N�.U@#OL���R�6�5t���E4H��!�ip�|�rn��wn=�}ry*�Ay?x�P7� ���@���p��e���9�!"\4�6c.��;�$X;����ӏf�̕��4E�c����KZ��Zڂ��c{��zaq��;(a�&2�V�`igR�Pʻ��R!m��â�L��W2���oD�goF��a�5�֍���H��V��������&�>`��/�r�֨D$}��>>>>>>2����<l�:�	�A��=	q)�0k'�<k���I�{d&K�Oح�u���;>��p����n�J�B��q�p�g�	ŘhB�-�� DTx���[`�"y����>�'eB{O�����eʙ��xX����eeso��c��c��Ƚ��O>��k�"���im�9��U{yu>��%�{���4
4��>�O@@+��-"�c�-�zO�<I�4�������	��5Q��q�.�<ܪ:M�E1�-�@��-A�6�zd�K\������Z�<�����%C����B��~n|3��^��pJ}%��0���SH���I�m�op]�[c!��Mn�>4%	��@��S�N�|�y�w�\���Q�ްܱ�AżD#���zZv����
0<DsW�S�V܉P󞘖�M,�z7k�P�R��%�^3.�wy�eE1��[���W@ߔ[��1�|�'�����h�~��OtG�?Pݼrh��&�ڕ�2�����f�ƾ+����j���&���q���vO��s��g=f�'�Mͼ#�dѤtFOM�w���l�J^��wx��sCQԋ��uR�p+S4���$��M�
a���.n�D�o���uQ@�zp�j����v�J�c�*r�,�U;��¯SƩ�Y�D�x�y��^�a�5«X�c}g����Ĺ���޳���3g~s<zZ{�o��z�^�
<-z�E�Ny���q�Լs4�!��~Yo-�ֽ�/��CX�K׉�=N�_E���a��%�[[�a1����l-[/H��vM��Kպ�.�O� �l	N����ߐOYє��z�Um{�A~�8�^S�<`�iiBzD�ħ0�~|����*�C-�YT�Vb��2���O�x%yQ�"��-z�CҞ�oVE���N�,8�[�d_=�Ql	��."V5����Gguț��v�t/����� ;��8���~��=!�&�U3����1^!P�+YI_��Z�8�|��m�M�hp<;��y�IM2�dNڞ�ֱ�l���!�l���BF���Y�����[�f;zAxL���.���[�$���#c��}��tz�Bޚ���^3 
zy�\9���<x�1��"a�1��={=1���N]��t��������b�ө�`��E�=��1<>6y��bo�t'ǫҽ,�a���5�Z13�|矸̧�e#���c93�d-�L^<�[�1�Rg�x�\���k!m�S��cVFU�_Fŉ��abD���&F��`2f���j�w�N}S�r�do;"�X��X�e�p��N��ƭh����siYT��(���
�ą=������y��`���WFNɆ7��r�4| ��.��!����_K��	�[h^����2���c2�����}�5.��u� OFT��>�d�S4�L���䧚�{�M_��ρz�5n�e���v������%8\W�t��_�,}UC��C
��i��T�����&�\X����S�u�1c��(>�ï��d_���F��o�!����0�9�]����uZ��z(��_����A�^�ߐ�8_���Ɔ�ua͍q�}�G�n%鋅0�8ȉo�r��<		�'F�&&q�:�ǩ�m?V�5�U���9{��?��W>=�bD��h1���[FT�C�l��	=C�Zsyz��C6IwXvߧ�*�6e)�q޺כ� �Ƀ� >�6)���N�z?cE0�����2��-Ӵ-D�V/d�&�i�Ԍ�Zb��:k,���!�^M2�tgO=^�w�Xt�D=���h��m���/d�r~/m�:i�fLk��p(�c���sc`�;@A@�k�/He��R�/�G�e�w@�f��gT4�Փh��ެ7�xN�ߥa���׶mr�T������^��ݕX���w��F+�Nc���m�&'����Ѧ�Vp�3��+x:��)C�6;��wO[x,��Y�˺�jʭ_��1�`��{�e�׽���ܦva��+����ctBXS(���'9;Vt�Z����ƹ&*̉&gXK/�ƯuE���J^Z��DYGD��,hT#�ѱ�.�5;zE����4�o�3�߇DJzE*
�IN-6j�v\�yF��7w���p�p0>��kh4g_��;W�礧�2�Tk��0 b_c�E��G� d�S�o*֏o�:K��3�����]A���+������i'ʘs�e~�N�|�v��������nwf�r6��)�u�_�H-Z�H�2�\���Ң�Y��� �/ǰ�'U_Y�1��l���H×:�Q�<��f�?�ZPX��P�3���{|w�F����be>i1���1f|.f�]N�ߵ��}�+�^ɯ�5y�Y=��Q�"�����Jlwn����l�����1�楮d��0'��`�%�?0ӹj8��N�T���˜J<���Υ{��Q`��� ����}/�0̮�-��*[�m��ׂ5n���Sk��I�9\�e��Az�#g�����x�	� �o�&�y�f��T@a2UHF��^zeԥh��|�g�OӲ�h:q��FQg��T�:�b;ř�T7p��k�bOE.���sV.z�)�Љ�n7:�h[���g-j���eJ����J:�����on>�E���]x�9��5u^^�y|�J%��1�SL����|gnqH�3O�f�&zD3Ya�i��1e�Z;�5=���Tj~VB�S��nF2����B�1֙��\[D��%���xA�#`}��N�=X�	@~1ޠ?��;��ގ��t�3�3��s�|\SU�4U�O-W��諐�{��E�-�\��Uܐ��w6[W�����;��=A�q���ш�Ԋ���F5{6��d�,�c���5��,tK� ʊ�د��e�ئ|-��6H��%��`ޡ)�LȬT)>)c�j��`咸_� ����~��P����qM�J��)F69���L5�sk�Xz� ͭ�F�]�';���k�:���<�	�%"�2s��=5�ؐ��2/�逓��g����MՊY8-.�9ܼ�Jg����r5E1(�aϱ\��cвH�#�Y�PI�bc$$�lg���6��6d��ފN���-�]`�LVϺ�q���>w�ޛ�d���p���]ӣz\P���ؽ01�N04�jV;K��pw.z�G�ߥ��$���}eɄ
������� �f�P7^+���3*rYp���т7:s��%�Ȩ���˙:�Qu�51q��`��)_Z��o|��ˈ6�i�3yU)�G��d]����LN�6r� va��w:�T�c���.ȗ��ӧ�a�d3�m�gvJ~1�c3����~swr�p�Z�H\?_�_�Q!Y�ܲ@�Ɵ/�>#L�F��*���X�C��r��~�B�����f����w��� G�8t����q뤱����O�/Υ�����˶�������ΡT{�U"�K#+$cF��;��x�*&n<eo`Z�M� ��w�vv����c��N=��mF`��G�������/����a��疨CS���z�\�$���q��8�����lO����eoW��4�Ew�6�]M�O@$ ��Xs[���;��W��=���E�����Y^�]�GomA�08��L��YP��#�%;�znW_0�(�w�顟İi�gb�#*�����)�!K���+|��ut���{�����O�\<t��3B=��3�(W����c�jټ9����-�jT+ݐC+����[_��ojv։��(��Ї�� ��1��
!�~/��,:O>��M��'n|i�=30x����3l�/v�)j^=(��������נ1U������F��6`p��׎��q}O�Rb�߁Vs�6T��:1\����Tc^v7K��;�/�Lo���ٖNf�a0K+���[�,�|C��w���O&s^�b��$�h�(n�լJS͋Z��7Z�����W�W
��im���i�����@>���`��N�py$�{^�Ԣ8I��s�L���d�"��Uo�\�ΞE=���H0�{;Ҳnh�\��^�<��0XG�@�5�^�fS��]YS�lm+���|+��6���C�Tq�f����y�-���~5�+�b�\�OH����w�RN]���"���g9�����ww����B�t����@#�<��tݓf�Ay�]�ߙ��8����\�'ɫ��2tr/��2{��6��tB��]���~oM|9�?�T�����X����М�i���r]�V�s��eἆ����Os�}w���5��X�t0uϾ���b(o��Ԛ�Kz�q�Lg���(E�k��"���T�Nl��^B}�a73-e܎�}7����dG:֔�$!�X���G�,,����k���&/�+VX׍83��ty�:��Q`V��ϲhqn�&��b��E��N�����rM�`�:�d:قx��Ϊ�=�|��/F��0�o6�<ç{�?!�!�~��-[<�yZw5�f~�EC�\���]����q�b
�ۡH�J+w6z�[#[��"5�E��[���.�3�
��:��R���(���J���BJ�ۗ+i�v�䊼n"5�Z1Q�Z�!������v��5���5��0��=˭Nu�.�FW��޷��>-î�����v�m�Tw΢��;��J����ءo����ԝ<�p,�m���))���S�j�9�U����_J=*ԕ�tL���ꂟT�G��]*�;[�9��Y���}�Ttkj�uau����Q�4Є^��]`����ʴޝy,2s�ڶ��-]ڴf&���
���/3v��փ��w{�C(;���#��W>7{-�,q��@��V�Vn�&t�%�uA�E�[1vfd�uW��en�0����_!���ړ�g������x-5��ބN��E���ifc��i=��kc�.b�}���XńT�Z�7êl��.щ#�곓8!2^�BX)��N"��3�L$��R���Sj3)���Mh�*�p�[7�kUd���bve]��,�QꝽ�(��̍Ct�M��T�r������8i���-�f�7u��u��x�Ӳ���Z��#���J���W�:��V�]�`_���+Z��v$�f�;j�$�,�Q)f�n���ܚ���Ow�#nm��#W.�׍�-�w�,��5P2{kGF��ن�¥���QfƦI�b�mݩ�OP�D×���&H�6�O*�vnlY{,'��#N�n煫��P�{�Q�ƳTCL\ƃq��urZS��2�5�ə�g&�4s��fi{/0�	��6�5�Ĩ�U�%Hg�/�T7�(����j�\ewi��z�>��y�Y�.�lQ�vtNK1��ꎌ���qs�U�Q�G���5���˻�{��=nk�3��rT�qBNu9�8L;�XnI,۪�E�ѲC"��r�7��Ot�t��V��ɕ¨�0V�/�k�ŶL�X�^�:�y32�����	�Z�F^Y���ݺ���y���9U�s�Ė�S+jZ&SA����Ɇ�����gZ�����7\<C�7^#�Y+�Ɣ��y8ܺ��̭���Yw[�1�G�80W��r��$Ry۪eS������W�Q��Qz�v�K!��6���g2rP �aK�/C���B�L��+��^�|�p�rɖ����k���NZ7���f!u�6�����99��dD�T'��Kao,�;�-���FΦA��H�t�h�/��o%<���.�ZR������Zgq��ͬ=]9���)���Q���`]�(�u��iĶY�1� V��1�[9O�rS������Af+Xܽ(��X��A��0��D,��Yrj�2�zuP��[��pV���UQ`��8Xt��U��,	��S:��XT�9A2�B{� ����V�si-F�
K�m���<x�����Ǐ^�{�6�h���jJ�%*,�PDc׭��<x��׏<z���)p�5K�D$I* ����ƛ��z�7��{x��ǯ<x���{R�� D�bƤ�E�r�[��)Q�]6��<x��׏<z��`�W,X�mcQlmi������\�Z1]�Q��4�r�X׮�)54Dm��[so+wj#X�Ɗ~�C�\�kF�QQ�5�[�oэ���^Q��lhI�Z�]���Ţ�+k�\ j��P1�X"d.�b$�SU(�N���nYnBZ��Hq�+B+B��u�������U1E��f��޹Lo!%bIp�oe��F:���G��\����y^�V�	d4j�U!y3@���Ȃ-��D�UzOGq4�I�J)�h�.P��2�v�	[xߚ�BH�H���w���z�t�˻��ӗW��̣��}�3��U�����<��{%(����P�lBR��z`̓��_A��p���K�#}���$D��p�K'��iZu�Q5;����O�U�A���Й��R��j7��w6lf�z7�>��U���
BTD����^R�a��o���<Ex�&���f��*>T�v�����.�J�׭�	�|^<��zb]blv�q�ճ�F�Q���,��Ѣ�^8��j�9�5�lƩ9W��C��U�-���	جb�0�b �O�w
yo=H�%e[��s�T
J�nr�����{����,,6�Ь�-�J�Q��sy����]Aʽ��[��t-nG��zd��.3CU9�3 r.�#b�*T'���A�m���Ū��|]�|��ϟ	��[ν~�F���8;,�n�zim���};wb��vGr�M�eS��x�Wf��t��:Nչ�v��}�� �*:��\2�عbRmQ�8"��̞=@l"֗fO���!��Av̞�scߍ���TLtY��`��;����8�$����V��wT�3yU�^\l��Y�m��E�ۧ���ȷa^q�,�噹�V�1��e��F�O��2��śe�){������7�8�1�_3�u�=^�U�D��\��q!n�#۝L�ˤj/2�0QZX(����(�8��Od���z�B�C�IL�Kx-�_�n�� ۮ�,�I�"oH�ށٖ�X�Ё��[��Tab��a�ؾ��ٛ��'r4��^�v��c<�=1pG�I�#��f�U3/���I��}UYֻ�� �H�)���89c��'LN��ĥ:s�9P�4�^�����ہ	�{���Ɛǘ؜h~��:+%�,����l��9�)�D���:XU���H�JG*#O?���gZ�솖{ܔ�2`Gjwݫyծ�I�
P2ف�|�ꇸ�pq�����$� �e����ؼ��Q,�6}�~�����ǅ���R����x*���
��}�Mx?}\ٹm�5�j��>��8�(��H�g0e��lJ�YZ��-��4�;ho����W�}82��zu�Yn��0v���Eh�RTmT
�T2������J U!�gva�r�2ڌ��J�I�Ȧ�![ǫ�P��Z�[�~'v��ٶ-Fe�kbr�je!b�q�o#[�ڤ�r%�~ �����~?��b�H�j��'�ѱ�D��ʄ������Dщ߈�d{.�-�o<���9����G|�@�%炭F�q��ő�gʹ����J�Z�ѷ��־�X�r~]|[z��F����Y�>>��Z��w��,�����v�q��doC��t��F�� C�T��{�o�}-�j!Tż�k}L�їڬ���6�vC������H�r�t{�`wxU�.`��l�"��*�2���k��0މ����I�!9I��^�h��$�t�ՙ3��l�8��3r2�kc�GW��,5]���Oo}.<�UN���s���fw����ր���*�b \H5��=~�������W�m��0*(OBt3ѵ��]�NM2)���������R��/Fʘ[͆���HP݀��lN+�X���3gĒ;l?����mx136�����w�P�ܼS3���j&��s2����Z'K3lnЅ��o�\�܇�':��(r�J�� t^D��'��Od]XǊ/�q�����*�5tM��[��.�UT7��1�V�E�+t�J���hՉ��/�y�}�����y����ڵ�]9Y7X��P���w(o�Yrh[	�較����jK�{���ݞ��N������yz�{x��g:T�v����h���"�c����m�Λ�M��3ffD�ۥ�q:ٴ���
� �2��8�>�Vǚ��Դ/���n��HjB�pc�?�.S�m��*�+<�Ʉ{tN��Sܺ<�i~�Z�jY��2��(��pS��Ap��n��ٴїJ߉��D��1�}F�Z�+�
Y:=M��qTi"����`|{�mT���<�Q%��<3�gTZ���B	�c�-/X��������`�nT<�J���9W����᭡U�����p�-�,�����h��S��F�3P&�Q�[罝e����ݭA!����:����f:6E�����>DXƫ��v�$�v�7���#Wr�x3�}@O��S����z+yw:WŝܳJ�f�씖I7��f�up��::��Q5p���yq�lͳ�KS+^�ټ���iػ#Ѱ��h�(Hjk1hMU�άh�����r�P�����G�=�e
ӹgVB:c��qs�f,�!u�P�w�^�w��MkO�1�~��w�+��U��ɓ���v�6MѬ�Y)ө�G	�z)�2qݛ'cX[�s���U��[�Ux�B��>/0!��ї٥�6�k$�)=�CWH/��G�q�#K�5��+�C�]b:��3��,)�>ǫӤo�'��hO�y�?����/yc�|�P�a�i��5n{y��e�(4�'���8���kĒz=���Z���l��"���[*�<��˶�/�����B���<6*��'�@E/r���^�<ۆ���D?V�L.�2#N�r�G��8��`_ @����������m6�f��r�po��	)��\"�V�u��҆�ku�%�����*�ܖ���z��t󗫨�*�FfK_v3FɳI�'R8��̌���5�A��UwzX��Zk���]CJ�ܝ,m���%וX���� �����M���9Wv3������m��1�{�m~��l@���Z�%Md�G��@C�9c�̵N���5�jEB��;O��(�J�֬�mJfW%�֠A�¨��������[����R���"YSռ�$��C7T�޲��v�uSI��s���֏x{[35�>����c�o�w��̱���������O�-΁�ۻ˱(�p�WC-]�2�빙a��>�J��$�0�.s|�ng�l	��'oTx�m{����l�Q1��ye�
���QI�̅��'���.�4���R��W� HuV�F��"��I�'�n6kyU��+��w/Hd6�1/w*dk�_�dߺP�;�}�=�xUj�=�j���k���>�f�w���y�z汧�X!�Tz-�t�[��0�������=ԮJ�z��<��+T�qGM]��f
}��8��U	�� j5.ٻ�����������{><}�u.��2"@dƑ�x�4 .�B���P�t�\X8��*�2��nx�@:�z���x3=ڑf���� �o�)!��^כ_)���$�<�pTys�KBg� ѢF��n�w������ܢ�q��`�b�KO)� t���]�X���qj����%U�4s���r�����`�wsyX���g�����̐vmX����^��e���Ә��3#��]��Z>��cƩ���r�s;;��k�D�߃+�=o}ꚺ��U�D���<';KM���>*��q��OI���T�ǀ!�0C�=ܻ��.��{��7\�<��|!��r����^/)��c�Gǻ#'d+J}m|ߞ��TM���<���Y[�U=����mג*i�ղ
����Ʌdxꈘ#ϗ�mF�[1*;%�|�QH���*�*�i�	�xp��~���]9ts��j���g%��K�Oq�'x5ӭ�d�˪y���X3�5�>2C]E�4��_>�w�I�%ZR��j>�toa|}�d�\�sP=5�
�N�v�-�0��6�{��Ɨu����N'e���c֎e�`�^�0|������08y�l;��ۗ��0���3�gH��-��Y}�`y5<�o|�쇾u����2Yh��9>V)�3�Vn��K�����]UK.6�СnmO|~���m*
���L!��P��L�=�S�!�*�"#Ѓ
E($Gt5i�C�s���2��Û[.��_4F�S4����7W�ۭͫj�]jś��7,ۗ�'��0Kob������y��o;����v��P���^�/�;�^H���+D�ϲ�φ��:�8�F�u5��j����0_+��4*�)�<��)���I�f�^a��h�J�܉Oe-ׄ���="ܯ*���-���4���"E��@�Y>�������c�r�؍�^.�*�S9�� rK˽�mFj� ����
��TCq��E@�x�J��������#QU�oQ�aW=����PqN$ə����7r���x+[�/א�X}'��zѯ�.@vU�d��,(Lk�Ouo9y�������uO��N"��nG��	���g/}�k��8g<���b��룠��Ԁ҂�px����{<�@�Y�$b\]�;WkT��uHA���l�>9�ЉF
S�>j�S�0��X׾c�o]�.���c#�ßi�ڰ^��
:��`׎T8�����x���k����Y�釴+NT�Bts]x�MԤ���7�
Y{�����;m����������Y����Er�N�Vd�ך�%�V���K%WQ
��%�Y������!��3��F;���;E���L�	p��6�v����R�^o7�����dP8E	"��[b����{���ifIn��N�n�� �FQ�t�GC��׼�З�s�ً�÷[����j���;�Q��0��l�f<xm������ֺ�N���li��7��jeO�\0d��q!/u�3z����X��(c�F��!^�����ٻfU�J1x��*�3����Ճ�[�r�ىc@���<]�-η7����O7f��	y��S�ا=���M�ޓ+Vn���/�b�T�qc0�W NR�r�Ѫjt�ۣ_Nsvϖ��� �a��F!٪#�WdV��{��u�Ѐ��Υ�ϲk�v� ��d�T_l����gi���``M��3������8z3�%^��*���Y-��f;��	��n���s����)��m��:�[N�K�:`�m�'����Gv�$��~#C�h�-�C��� !F@�ᇍ�Sk"����>~���ޘ���&�\�r9&�[�����'7-���#\�:a����ǘ��G�t�i񯾂�_P�N�)t3wSE����2�:���F*�s�����4>��r�p�5����7��
�D�pmL��^�������D���I��xƅ<!���T|*���{~�+�Wr�U��W_��m�`L#X	kΞ���2�=T�eH�p��#������=�^H��ҮQ�z��ݲg����qb;��&��}�8�Vd�2��_H3U��dp7��{M�D�M3�3ʺ��H��E	W�]���J_���k}�X�᜗G?���b����o>`�o����U�+���,N�du�6sq����7-�J��G��N��6O�{�2~O~��c&Ëq�in�>�'�7É��}���]<�L�#Ux����������-���=���b�St3�Mj5|y�Q�.�y�3lz7�3-7�J�e��|��a�[.ՊeԈ=�MP�]Uk��.��N�x�#o-�e��Ͷ2W*1�x�dz�"_�wk�~�������o��t�V���t��&�I�u�j��O���Tm�;�:�U����֢c�U���yW}L�]����P�Q��£�Sz�q�:qD�܌��h�N�o��t,�R:s�!\�o0��N�-�D�,�}�?\�	g\ne���_t�'ld�w�_*��gҨ;��Eu�W�Z�l�9�h�7Ϊ��p:�݋F5���NN,Jꔝ�|)�`�:�[)�;!3F'+6Kf�	���W���y9��S*v�Q�����E.�_T��ݻԍ��J�Ee!�ŝ�����u +���6�ej���
\�F�Em�Z����3�Zu�7xz�7/"y1�<r���w�7�:������o�Ӿ��si.�Ʊ�;0��7�l�d�v��.�%ɑ������l�˭�`�v3'J�Q�8u�6sM��<w"P�ԥ�2uܻ��J��5�zl���TmڲD��ӌ9Y2�(�B��P)<�*�n�k��/�E�ᗻ}[���;{��Ù��v���cn�4���[:"[ec�$�i�{���N�aQx�ĺX�Z��α��XFR���e��Т��r�c������7rqZ���q��\�!A�Ѻ)¸4�n�2i��Ԓ��:n½Wv���1)kn��m�!�`�-bG2�Sۑ�p����ι�X��ⱚ���o��;~[g(ȱev��ɯX�}mYӅ$7�Z)�1-�ǳ���LĽ<C*�z)�C���N�^�fOgE��%�/ѐx���� �h�[b���4���#&Ų�;�?]��Vى�S%�[ʝF�o{ȫ��򬮁��ݝ�K���w���o&��e"J�uJ���ħ4����\aэ�q�Qc��r'���Zb� ���wGO2޻�G�n��FE��f��;��0%��t!�]\OU�on�"AC�w[,�9e�V���f:�8ڽlK�9�
�"�G�V�	y�T���z{pm+G��L�Y)���\�"�묀�gI΂���q�(C��$�[�H򡹯v��j�n���!�*c42�/Y4�+��UU���x��N�N�J{�L�뭳�0ѵ�7����`�p�ڙR��Х�m�ĉx��q�eӉT��"g���]��YP�gGfV�4�_hB�VřT�מ��U�\�0�(c�;������h^1�~�{�Ӄ��5IϤ<�43��Wm��.�W �ý֮�A����j�f��h���.�<�5�eUXF�{Ca��Z6�=�zy�g^)\	Я&[(��0�^�o�S0��e�b�+��S����Ξْ�Np��S���d�X�Tn��E�Iq/v"��<��J��<vW`(��ޕ����M�2G����e��4���i\��8f�%2�n�����*�0�̱�Vp;b�n)dM��{�֎y�|�Cd��	PD{�@B�BDdR8���ێ<x��<x����	@$P*�U��9UEQ���q�<x��׏=z��BMQ�5�Ū1��@$%JX����q�Ǐ=x������U�X�W��X4Z�}x�,h�����n�oqǏ<x��Ǐ^� ;DMU͵�_Z��x�65����[r��Qm���[r��F�-�WM�ݶ�͢�Ƣ�[�W�^5�Ѩ��j��6��W7��m�>�.����*�
�.��{��CH{��|	[vr�mM�Yb���.VM�݅T�he�&���	v[�;�t8�l���^��lީ�y�r�O<�ŀ�����似@>K��~� .;�����[�~��-YX��/���dP¼�k����&s�E�,�ى���^�O�Z���q������yК:��^���;Y��F�9�Cg�..����l,��ئ�mR�\���Q��Ɖ�Q�x�Ӟ�'��y�<�ø2���O�$q��5�=��T�<�U�c��v�������:�� �&�jn��f}վ\+;u�z�����){O_
�f��{憫@-�>d��13Y���큊z�UYy�i��0[�
;VV���q.�e�!���=G+KE���>;�y���բ(��K�DOd����s5l�@�cd[,?tt�ݬ�Ҙ݌�p� 3�"2�ּ���7���UB/�z�M#_�h��ǪiR|1�3ӯ��� �ls�U�{�ϵ��{��r+2)��5	ͪ����M�ۧc,�e]^��H\��X�����N�����Z�\z�f^��G8�^n���g+
V겖D��ł6��F�`�rtҚ]������͙Y:��=�#�W�@]�r|;ms��r_.UvY%��������\���)����~�5���Ƚ���qh͞J�*E[wz��ި����zf.����tTl��-q� �p��^�]8ck�o���q�܅��(i��.W,��:i�7S�����>9n�Tc�0��3�c�f�V*X=ɹ.�^�f�Z�	�OLe��$�\��7fy���G�.2"3d5&�����N��n}C��Eh�������1u쥻�`C�s�L.n3G� ��w�_���B��:ڳ����=;'��A��b�Ȭ1q8�q��������]#���\�~�O|"�wz6�W�W�n��8�Lz�E�ם���r�����ī4#�w[]]�ü\a��J�_g�x�r�'4���3�	\�ꝱ!\�0T�(E]���Ϡ\W@s![�q{�7�VGm\.�!��O�ngb���,��D��"���1�%���QJ�3W&�m����I띭�J]��._N�Ӏ�wZd��J�U�I<�ySq��8'
yA+�eG�j�)��=f�E;��R�U5N�zh`���(�
^$r-Daî�o&kVc�*�F�HPsKu2Ɔ�w0&���>>>>>>�6�u�6}��T��_3�L	�$���'�4�jN����ämH���ٸ�wΰD��qav��ǻ��B#Nl"�}
��^���U~҂��GO�G�.%��8��y�Z/h��$H���f�b����{�JU�q�Nn�:y�e����ަϜ�Q�GK���G 'G�^9W��(�3f�8dd+�Y;��_A��݈����e���@6�웂�����7�%[T�5�=[�؝���ݜA�O�&�}n�� O+�??��;����D�҂�+���o1�Y�D�yr�2��-l��+��<ֆHDoA���"$���r�tm�N^�z��8��n<g�k�i�"Z���>xUU�7���aD��{�<�l�G��}���J��A��0^̊�[S\�`���M�������Ȃ5��rɕ�-UO�;�g�lx*+�{е�	�}U`K�a�/��6S�Ҳ����d����r��]Urб⭪���ͺ��n[D�cws�h�EP�NJ�{-�Ո|O��`����^��4 ��'�G����Y)��U˱�!���Y=�յA���U39Q��I���f�=�~�������!��l=d[q^A�=��5PB�Ð�u�o6A�A�dML�dLn^$�2pn��Jz�yi��]�]����s�J����v7/a�f���2�}wA�ͨ�rlR��3��Q?xT���{�A9yݏok6�^�j��f�J"=�Ze����;<�������F���)C�;���$�y��7׀u�)Q<P��T+ٷ���_�5S�&`�������vC�Jj}���kՙ�9���د�z�i�Hx�4a�qс@��@̏}S�g.,/K@w�
�����j�q4�ϸlC�������nB���K��LA�P_�씰f��X�I��W�M	��.�Mj����ƂIK�5Ov�ۙ��J�v�H�@.�BV�!�;��O�K��^�ǯ_��ר�\d6�
���g�����DR������9��=�ӲU�����KZ��v9�D��!������PJ��,���^���j~~7���.׏k�nM�J�뙬�#K�.�2i씅����ǐ\
�Go���u�M�u���k݈�H/~�����}o$���0$���u��bqX��.�>��c�ʱ��D^��J�+���0���C�CV]�>�F�����my�vlz�1Ԋ�C�I7��v1m;<��,_]�^�\v3Ӫ��{O��VX����#���z(�EX��o׽:���ҡ�m��/پy`�?bŊ�_�����[��s.��r�8��i_�/���V��r�">�ς� ^�؅��=��R���V���x�Ng+ܣ$��؉��!�@�=�@~/t<{�|�zj��ﺘ�"^�fm"I]�)��m���9�c�֋Z�м5Բ�#˰uHVc��S��⮞/;�$oc~�@��D;<�SV��r5�0��f��Xِ|T/uLR�ϷsyծK��L�A$�ީU�OIΘeBd4ِb�#XK���%>{��n�2��k��Ϝg����̃�
"ґSY��i_n�,z���ֹy��՜Pf��խ�7oJJ��s�&��̳��j�V!#�0��e6cw������w���xM=�s�ێUg`fYz�f��ۡڭU܇;䞙����s�y��������?� �'sv�yjni��T/T�?W�0����k.2���˾��O_V��`����d����)�����vx^3���������ZY[=�K����*$F�`�&��zˢ�q)T"��.�Y_����f�k=��ۮl���蠹
)H��{�E��e|�Ub���p}�_e��j��c�Ǽ��p̜�|"�87��a�aH\�W���J5䛨�-��^���hh�Q�}�Ѷ�����Ú8O�ंv��cV�9�P��zh�n�u��N�y�������Gqw�J5����_C�>���>��N	�m���CʼE�̞��#�����+����dK1>O��G��kdǴ��\\�����d9�[�g�&�M�3r1z�gO�0��B��յ&�WP`��R�;�����8��+�bOD5>�]`��٪�@������ΠK��Z��)j�Y��2�T؜%�ʘs���U�k�e�O7afD[��V�׼y*�P�j<p�y�Dzx�|�DCcDӗm�tJ��85[�+�(G/�Yr��kݴl�O~�c)eѪDUͳ���N_��z�zf�ل-��1�`Ql�u�fEuGlRQjJ�Z�+b!��#37f�5�\L���z/����`˥��&����>�o4�v��Wj��klB]�����؁���r�}�
�z;ؕ�+���Kq��L�EI+ܕ,�e��I�w����م� x-��{�BS�@>�{ј����3�,w�Ú�}�,np�j��f�M�v�p�|R���u���X�o�N���"fLߑ�;�w����F��֛��h�q|�RC���(܉D)�F^׳3�jø���r�f���W>��)Yۯ݉�Ex��g��v�Q�k^vW"5oj�x��#�xgI4�*W�&Y���%�׳4��}<�/��q�#�f����J��h��}��=̩��	��ض����fh�#��˱x�4�Vө��ǝ&�p�&�Z/y�Hκ�n�R7v�oC��%����qi��כ1�q���}����;�}�]`OٰXɛP���.�^\nO�/��ӭ$Ĉ�f-�������x1+��*���`���6�$�t$�:꤇�	�"�Ɉ��[�ٜ7'�{��m1�
ݦ�'Y����	�eܵ�r��N�"�X���Q�S+]4	�4�����>���V�C���yz�m�R��4�,�n��Rst5��|�)�0���{ō1���H����_��M<���Wr�|���\��~�Xgñ�'-GH�bb�{����ڢ�ʞ_v��cx��.�(UYn�y�K^�nX�xsX�<�E�#��FDmǨ��Ӻ9�m �q~'(a��pK�Y����2��߮ԩ1�w�3͞��:�v�~�^����H�p�t�ᇵ��Pp�GL��3���i>uf��-������Þ� *��rMwZ*& ����"���l-�î�&��
����d9����C�C�ڊ[(u���"��ӽGT��X���s��LFe��k�.�)îA�X>����Y�f/��,��*��p�W)��ofy�/�����l�Ův<�����@�]>�uʫo8
N�$��N��4mYݨ��K���Ď�R�P��V��ka��r�f��+ю��L�}�%{��X��bUp�Tŗ���FpT�:ꌬqP�ݞ�wt���*��u-�t�S,*��T�]�g
��������.S['}����~?>�{���ӛ��׮T�e��U� �t�H�[�n��P� ѝk�����uSܓ�]���O�8��u`N	�tB�s	V{���ܺL5+X�]��G�O�ћ�/�9�q��]t�{$Z��iF��S�eM�,��i���y��)!�&A\d6N�S�z�{L��Ģӌo�ף���� �}s�1r(S[~���O�Ѝ[j2�x�R2v�љ{q�-]�☦�td�G�|8�ÛI�q>�D
�|y��i	w;ר�Ѳ0������ﮢG��@f'�0IT �e��yr�+��N���5�{�en�]L�R:�=�϶��!��t��E�F�f��b�����]{ϛ(�sy�?*N�[F���
�t�1LN1�:;9�l`���h�ȿv}��s��m�L�u��r�p�#�xK.Z�E���}�WHOUf����H�9RqbVWi��Y����R�6|ش>ǰG�3P$ql��R��f.Ml�	r�ݜ.��$lAo4wI��ԓ/v���98:�+v�9��UV��gq�f>��߼||�o7�Փ&wLU"��IO;F�z�T�F���$uϧ�t����L�Y �3���=�} ��oC�Ҹ�Gpcյ5�r&���ĵ)쎗h���-Sfo40�1��}��B�ozJfXg���U����J46�ɟ>q��u�n>��Mz,�ݝF/}��`�ug�F¥	���j��K��ϗs�����:�+z������fï��ʁ�M����(��Z���~R3TL�l~�ˮÔtt��IPX�(����K�m��0��E*hԵYIVP$~�x��t���>�6����t�BT8��B*���F�*ݩ������]C����4�2�1I���o��8��b��<Uj�=�l�8�ѹ.�ܬRp���`��'��k���]�QZ,E4�ƨꬱ�P�3�h�=]��h�Z<�VH�����5ɐ�
v��g2jN���E���(�������U,d[ض����A�䨪i�ak*q;P�l@z�����l�gM�Es��ɸ�t�{���V�sZZ6�#Vr%*�����>������3J�n��غ��|��������5��`�Tz�,Q=T�}҆�j:ΡW��5�j��n�Ͱ�=۩�b��d��{����޹�V��n�A�,]nSv��Y9�2��[��,�iZ�]�m�� �SCu	��r�^LC��otVFV��d��S�y��V�WrU�`2���bl�!����[K�$�������$<L_m��h�ɭMzjUP�k$�=�(_��̣:���5gcx^m���st𐎼����n�,�%%b�Xj8��vc���V*J��/
��HX%�sNf٪�d^\���|m����sv�ZD�/mP����Ց���6�kyb��Cn^6����7�5�ch�;h�/$Ӌ��l�m�5R5��6U���/�"��r��w@Ĕ�:.���]^�A)�5�xm�vi�Sh;zEF�\�BU36�JQ���Q��>����M\��ݧ���+ӛ/�&<��{F�E��ι�L�j�s������F�j���9���x�٫ͩh�UBΒ
�n��N�5/T�*�aHdTw7�r��B���J����c	OW-�!}�+ko�Y1���Nʆ�X�Q왪�{�ڭ��z':q�ti��if��:h���˟O�VË�f}��!u����dmS�s_���5u�s*oi�`����(F�)��1������ٔr��aRմ�3b�n�+N�H���N�,���+V��e*�e<'&i	ղ�¨鯂�Hhx�l��0�W���V+h�s*ŝ�Z��.��t×{,��ڏT^�xs7*��`Λ��p�sy�*�.���o�Ċ�r	�ǓM*Ƴ������:*j�a�]T'��}y��g)�5�MV��"���g
f旰5tLs���7]�{.�0Nc7��5���#WX�n쬈R,|��#yy/;�)2׸VY�$�J�[ըm;��A纫ն���$@�¬�|p�p��`�i�8m��\�F�ø�"Jݖ�hv�����ɩuj��.��N�����]�1l����vy����Y��]��O�`��^+8�uM�&����k�3Q��*�FRU�u�9��륣z����^�����V��Cx���p�;�����+Ոē�E=��VI�:��H�@W�$f��8�n���/��V�í�#"Αr�WP (!C��b�0�b��ѥYY��ٺ�
�JK�)��B���ڹĜ8v�A�ԄdI�%<n��^�,GEI�*���[��&L�c5�X߷��T�	 <��QR�T�J��^�QcO�<q۷nݿgnߏw����cFыcj4kD�A���Dco^�>��۷n޻v�ׯA�dA�����T�R�Eh6ѫ��QlcQ�������v����o^�zv5*m\���Z�ţo��5�j�=m���v�۷n޻z����4j�n��ֺm�nW6
��6ܶ�F�-,�m�Ŋ�5ʶ-������U�mզ��m�x�b�zmt�ZM�Q[�܂�m��sh��F屮V���m~5��x�ܶ܉=�j(HȪJ��{&��M\���Tȓ2�ㅰ�q7"	4�Y0DL8�BD�=����^��a�4�Y�Y8��Ī�2o��\�T�:j�1;.�ڬ&�:�F�h�6�b�h_ا�E�d"#�t
l�h��P����j&�e4��0A�&�e� A�XT�EW�$�� `)z8�&5[z5��&ޱ�`F7�=�Og<���f�&ֻ�ۥs��.[�C:j�2�V\]�����{���y��������$���{�������XU3��y�u��v�{�4���Vf�o�R.}KK�[�������ҷ��t�J�n�:eZs��u1��y�~�"20���(��e�p��P�iDI���vjՌ�rl_P�BG?]���+��#�O��A��D�N��Q�=�pQ ���1���逮�]��w��7�r'��Hg]��]�����d3��z=�^��`Fߠz�Ŏ���VJS���'T��=���ǻ�؈U�����9ͥ-�t���V��]�wen�8����$�B�/��>ا3��9� ��Z� 7#p�&�.:b���u�m���@r�a�x�����mψ��}܌�h��4$)^�Ww!0��M�f�!n�w�Y��	�K�9�,����x�e�\�G�㋆S�o6�)M����K��*H2[��b��v�ݵ��0E�U9�1R���=�-��������7;y�;�����XR[݅���ɒ$�a;B�����%Ú��͢gL�p�wK��m.5�Z�I���/왹�ߏz�P��*���F�4yb����Y�JJ;ʭ[���.��v��A{{4���ȫg����ohZ-l����u�pZ���Id>S9������؁�]�SK{�n:���i�D���@>��5v�v�s7�˗E�vs/+TOYtU6�OY�&�[1��nWB�WtC4�egTh�1����b�?�i�d�[F`���Wq�W�[��7!wst5�vr��/�~2��5cL�`/1�6�FV�y�.������v��Ј[��{ު�&8��8}`��`P��</^���9�L��SK@ރ*�j�sԶcV@�޵$���"����6i0m�p�ϣn����z�{��p�Y��x�>Mi`?W���ͱ���� ����=�����(8"��D5�,�=���޻�x�+�y��\��!��q��}���ET��<��	ZO.����	���d�67�/�%�h���ǘ�I:RU�mB\�[��i�:�eɃF7
���QWK��֜��%�;�X�5��:@C'o)=��*j��pb"��4�E��Щ����-����a�k9�<w;��5���=��������ҹ^,�Y1�b�fza���k��u��p��on�C3�;��4�=����4�]���dXx>xҽQV��ow6�nq҈��Z<9m��<OV5���K0���T4?F�y��DB��g��U���I]�� QΝLp�u;1w�օ6i��l5��
�;V��&��#�**�-���z��<&)D���[�5��/MB�,��f��
����\wv��ɼO�E��^�WۥyZ�@A�\{0ĿM2��	?c��ˀ���v&��"��GB�K:�+|��ƨ�S��u=�E�j�4��a؏-"�gN�#U.]z�v��,�7zOB�25�a��f��9�ZVe;'ٹ���n�����=[<�L�6Q���[ �6��E���Fj0Aa�f8 "�D.�F6M��򭫌ǹ�Og]�5�޲����%���λ�g#���3��ɮF�؇'�Qʹ����S0�n�5���_:W�3
a�H�1���nZ��uR�$�Y)
��'d�Ɩ��w����GkTݐf����r�^��<p�a,am��V�����&�����y��o=a��ķvB��R�����\��^Ng�k�t1�����N-U'�Q�n�bz�&���m�W���6�8#6�
3rщ{C��n5��?ou]4r����i��Nz�]Q峳�����x;��{��������WנN@J9b�K��M֘������2��K\�؄�";1�゘��ά���\�Q괔p(��� ���f�F)7��ឣ6��]�М!}
�EZ40e^Nio��';
C�3��6qi�RTC��]ٚ�g�ys}�Ꙅơ�IO�3�rn�z|�۾�`��b�{ zcW9k%;S���`�迵o��M*����P�u�6%�b�j����	��Kl��t}j�׼�Ǻ�/,ȹ�2�_�!vE@�ɇ֝�I�9���:�q=�
�8��B�=��=y74�V���Q��n���m�3�5(y.�(�w�����ڶ���6�\8v,.	)KW)Y��v	�}rُ'8yCr�U��u'*�\����+ھ�p��&^
Gd��Otu��� ���^lK6S]Vgi�u�Q�&���x:��%���������u�yOs�F�"�5�K�Q�p�v$E
��nՌ�e�^>��ahRï�����F�� ����8Q�pH����"��/g�k\c�$hy�������*�N����پ�04���Y���ׂ{�Wod�>&P�r�O����oIZ��0�F��k]�'Z(���l�m뿣Ы�;C� xh��OV��T�7�/�U6��V����8�>�͉�uX(�\_��m�����o�֩�ƽ�w�Tia�Eq�Y>�Y���(���s��@��i������K*M��K����f��>��=������0��379��Յ�s\�#l�Z׾��A��E�t��}�䢏�>�A�\�uBȎ�\4�TUP��coCa)�����y�0z�L
�v���*�����6y�en4i�@@E)@��>�W{�O��~�
dB_����eP��Ѹ�k�wp�Z���#��1q	N�m�2ܢ�fi�Sxi���5���q�Ż�H���6��u]���m��u-�۴nna��r�F㾫̈́C�)f���H&+k/!cB+gF %8�=��㬗��n�&ˈ���������y\�5X��\��fB�}��΃����9Km�u9�H6�D]q5�����`4��^���'��&<ll��r����0�8�ك[��rf��P��B��T�:S�!K�G��ZsmM���%�����3�]n	~ULD��{�=��Y3@Z���AJ��{#��sM==V+z,�y9%��>Ϩ1QB� ¿,��|i�������"81���r8v\đ��rjƫs5l��5>�Vh�Q;~���w�`t������"+��i����S��339/V7<`H1�	C��M��>u� >�Z���"�nk�(���q��=#�{��l��a��͙�T�!�;�N��7�4	r"�EȷȚ��\�3�mr��`Z���X=��̲x-�mڗ�\<��Fz`�1LA�Rg����6�μ;���'�1^�}{yT숇C���pM�!�I�2 [O]	׶�l�%�Z�L��b%�j��Y�>��G�򯅏�U0G��z���r��NA�0������b#`{Wfl�꽮&Z��Ac�muq�"�4h���{�=&ߌc�;���ܮ�;���1�4�`�?��;��kϗ�<Jy����?y��N���a�5�!����G�[J)���#�(wC���',�X�Ӵ�v�<�y.�?]�ᡰ���N�i߂6l�P�F�Ϙ8�0�� ��Ѐ�k8,�����捾��<[ah�ݲO@:z�:q2�z~>�.2=)gT٦x.�Tm�w 0W�/��9<0�C��WP�k�2�y^�*�kM�mX�g6��cC��Sϥu=Z5|⮸@�'AS�4�`�փ�c.���R1��ӕ�&�p����E0k�{�5諚�
�ڽ�R���U-3��v�(��:zy[��KX2(%Q�n{=�N�Q��7~8Gl\���7v�e���\K�;�	�����V���-��oM�����|U��2lɨ:����gM<KX@�ba'"̪��Q1^�.��t��#l����N*�����1oƢ��t�e8�u�|�'�l��Znd�En���dה�Nv��/v��Q�4��˭�Û8c���BZ%�M�[�gwq��<ڷ���J�N5�zލUF��7����#ɟeo|����4?�2g��Xǂ��%!���Z}�N�U(1��KR�ʷ]�12;۾4�0lZ�W8���ƹ)sA�Wl�:�E]����}���w��ȅ>���zHY��
��+�«�+g�2���&"3ub�1�o;a,t��.�����1�sP3�<����ݙ����2|B&T�W��ؓ�ץ_r}c��X��`�oʄ �<���AR ��E&�+*�t�U^�I��[\�?g����ǒ���������
`w��؜�Z^��1��s�l:V��T�4���-(��i�ӫ8�J"W@[9����3yݢ��W#�2M�6Vx�����6<��Դ��>��c���팳��b�"��|���O{7;�dp0!�p�{^�L
�H��t�� ���@�[S�;�T�e^����P�vX@�	�i��$A����܏�	���������T��J�Պ�vu�Y�Z�u�j��!�"�)ނ��r���N��D�V;V����B=5��UQ��y\몓y�%��q���I�V�2oQ��#J���Y�y&�7co��L�������Ւ=��������V�W5����ߖuJ��>J��"S����R���~����E1�.���#�YjI�c��wM�o*�Qy�4My��Ҥ�-z,h����MQ?`lj�"��r�a�睢�k6#��|�ޘӋ(^����{E囉s�l\Z)F�̓�H�Ә�>!��7�|�׎%>6d����ȩ�;tv�L�D���;�+��h�ȼܿ(ńH�����gBUĤ�y~l�L�yS����"�Ld�0&��+ �̄�w��7�-�{D:�&i�'7����C�2��'�}q���N�����!�A\�KV*闛H��[X��Ǡ�W���;��!�x��oy�l58A;pY"5n�6�'���Z�H�T���i���TS��}�7��˾���v�#ʽl{&�FS�nrx���zc�Q�˞h��Eq�hϐ�p;"���g�P�����\o��+���j�{4Bm��-�YVb�OCXvua�ˌ�fox������+���.�9�j���bۭ,J�P������������Nн
Y;m��4�ԭ���N�9��M]��UL�G�㗜y�݆
��}9U�d����������{��ۜӯ0�
2����M*}=>~�u%i���G�f��*7z���gU�ǆ��by�q�c���X��C����S���#��Y��'��{���2͘!�&}�#A��z�����/5QN}C(z�%������>�^����vt�����煆���$]iuK�#]\C�+w�i���9p��WUʌ�r`xD�jK���@U�k(����z)I�[zjTH�������@v��ȣ�I�taX/=�Ӫc�a��9;BY�u�l���jl�8Z���B&�{�g���j���vw��|ǜ��=�ύ�V��DAJ�݃I���<�$�x��fu��޼���)�B:�,X�{~�U���+����WOqk�d�tb B��߶^kX�m0s`\ V���aA~ʌ�;m��&��4�]�ڜ��T�����r[us*�!Ъ�+K4X�כpC��g"j3p;�j�vС�n��vil�����S4�gkn�Z��]U�d�: �T��m\���Ǆ�鮿oG���f��cjp�^لD�U)�anN�*HJISsW/G
�0�%,���Wx���Wxo����V˹���Ow��9�7�r�R��ܓRS��xu�m��"���6ؗ�ո�	1�7`7�w(�A�IT�[�2�ѽ���'e��.�{92Nȝv;�L^����r�<۫k�����]�N��UjKqk[[ĩ�~X8��<�|:�ty�i��ͧ(So=�fM��	�v�>[��jf������*�M54T��a�.�L5t�����vwQ��w�-�ɕq>�Km�/ej�\&������&ݷ�,S4��K���tN�n�ʸ5�GK�UM�sv䪆�����8���{)Up�6q�=�і�c)�k��_3/Z.X�Uymn���-��g&�_
,_[�j����R��5�ťwg�6��քR؄&P��[�2��Όt`�b��N��7�iI���K=G4�7X�0�h�����R;nWmʤ��".�*��T���^���f��z�q��2�Gkd����ʝ'�;en���`�n�C��q�A��e;�KSH�c�MM�RJ1�mQ%�0�\[\��ʬ���z2T�u��N%c]��; M���VH7:���e�k��QU�Z�}���%��b��Sm�=@��8Y�D\�t
�_!�I�Z����
��a7��d1���Z7�b��5��"��b���٤n���Ҥb�W��wvm�N�C �Ma�}���\�eUW�=��'��d��2����n<Wu�v�<o[���y��*�Y�W]�8]ʂ&��]-	��Rʰ6C������	N��75��C���nS.6j��L��Bf-�#�AS�9�Zʘ1i��7�[��rw�d�䄫[)���'Pm�ͣ�Wg$d��Jw�d�55�mr���*�{��
e1gkx�KC̣�ͷuWY�"�! ��NvqF��{�wY+o�<@��g��-c�*�f��|��7�(З�U�M:3iX�ѫ�u�Q��uhuTׅ���ěZ4HoYr���Q�p���[�J&�ћ��i�&�W�������!�F|�n�W[�oU�s�4����v�S[\�X(CwB���k:!��M^n�YuACݜk-����3"���Ҏ�{w)������Pn=��m�#7���J\�4�KyD�Z�����b�bׇܶ;]CWJ��W&n���r�귳�b���)YW6��>n�]�9HM�����)�T�a��V�������z��u;s6r}^���Q���~&K�w�άRP�3L�Z��>����$ O���	"%E)�n<}q۷nݻ~;q�׽�ȏ":���d�:�]P�R�2)Q
z�����nݻv�뷯^� �������
�H:"�T=|z���nݻv���ׯ^�n/`�E���⎠��A��޽v�۷nݻz�ׯB��Ʊ�W՞v�Ut�sZ�m�rܬW5\�;�^sƺom⹭�Q^5����+sF�ͫ�5��+\���v�ͷ���~+��<zh��x�H��5�
 ����q
��� y�nQ�.T���D@M�Q"����ٓY��Q���X`�댧���(3�^VYz�a=�
���.:����E#p�ܴdt���+�0�s3S�	
~1�c�{�L�3�?�O����g+AJ�$UP}��S����g�U��|z�e��'��P�i|[6@��I_��m��ǗW��3���%b}b�O�3���"}�2Xhh��5��@���6r�+�ŭo|�ݱ��[�{�Tr�"O������#����T�j׮(�����a�)sؚ�{�ҕ���"$�\i�={ ����P�H���x��Ӛ���Wj�ܐϡ�����<����A���x'��N9�kڰ\�+��Ƀ3v�9}�|�������B��>Z!Q� _@cΧ����i<�_-Q�Z�]�k�1��~ƫ������mw>E��j'�pʙ�h����-���ku'W|b�T�xat|]s��;�@5p�Gx��9��F����a��aX>��.�[\O&��a������́� =�%�5���g�U��ڶn۶��-^��=�z��s�R�c���GI*��uG>�k-�����bM��}:�)6�T^p��K^՝$�]JmJ*�p�hɳD1o�aU2��޷7C�mV)Gn�1�,]H�|��ژ���B��x�o�x������t�2��x�/��[���@B�]��W3Y뀳�[�_O����a�(+.�݈�+׽Qz�w��HM{�[.=Ch���ns�ԫ��"n�����*�v3WU�<�C���S�I�=Mt��Z
�9����+��h����}��z��ohꡝ�Ea�л���OM<D���=�*L��z��޽�����m֑6������<%^))sƚ�`�������{X���1�K�1��߂�+xEg�l$o�JN+�y�z�ǖ%yy�[�#)_'�,n��n����`Z<�20�y�c��+�Σ��F����^'ү���3<;k˄�u�����g�1ND�	¢_��s�Dm��[�I�p��K����q�o�>��F��3�:1�)�����nv�����?v����%cک�H� �|xe"1^�&'*v���)5P�`��e�Z�e=��y�0��G�ۆ�%I��nEm��U�9�t��ѓ��%�,��G�3��̂ȂXWm���F�j����J���5g�k=���y�u��y+�h^\���w���rܧ�`=��#���||||||}��aw-m�̓�w���Ch��:RM'%�1n���5Z��L����W�{�XB�l��t{@ʭ�o+[3�w�Ǝ6����<y�Mw+Ի���i��ݧ�\�#E�����nv�Y$�}��F𰃊�ޠ�T�P��)��:�Z*����r"��Ӟ؍��wp����εڐO��:��Q�w�\z�2���ꦀ�U��=[dk���x�cԐ$���|��,Ǟ��d���&��*'렫uU�/�]��#Q	�Z�Xռ�����	��x�������5q������k����A採�ov����Ju�h��ޖ;L݋��r ]@u*�{�ী�(�P�Oaٮk��z�q:��s�=x��K�u6�F׬�]�хdG�dc��3�*����>E��F�G�$?]��n�g
�rc<�,O	��t��I/3�N����I�vH���V�ؚ�6���9[���b�To���/�죴v�)T8ş��wu꽆	�
��W_��Vf�Ւ�A1KV�v��[�5�tƓ���4u~6[G��ms�(�k���gk�u�+��k �����?7����z�8�v�������$���z�e��s8T�ٰ��Jx�#����E��&��o1���`��JD��Q��3 *�x��)����qJ��j=�"��d���ȥ��lN�.{(�\]ߺ�!�7�f�q���)�f�\������Q+��*�qE�԰>���6�A�j1�(��C�������쫘S�혌�BsԤ>�^�Y�Q^T��]^kɌ��Ц�������%�W�?��q��Q�q]*C����9�[t��C�-���%%�dH'վ�����\�Tpu���{�}�CՎ4Zĺ��'�q�{�r�հL�Q��p���hV�@�<7]�tLǟ�z:o�ؕK��}�	eV�j�葺�;�;�8���O��i�H~�I�"٦�������|�TUɫ��"�O+ �>
� ��Q�����I�*Z�1��l&j|pi�6��VP�U�Ǔ��z���c�u[��4)�*瘢s9�Q�h�up�����p��=�v��w'm��YmM�N�rحA�vZ�V�x$+�K��f2�y��Q�X��z�%[�cǺ���<�߲�澼Oc�Xp��^�x�O�m��h�G[a�G�U3���j5����#Qx=�4>�;�c���9�|<p{���I����c7��H��L�'x.�2E�=�U�<�!-��ϯҟf;M:��&��xgG_	It�IB�1WU��O�*���s�^��<�Ż�U^j���b�ȇ�މ1ϧ�k�IV
�0�*H~�6ަ24���i�L��#)*�l�;p�%t��hҒ|�K��Y��y�>l����u��	�^�~<)���.C<�UY��⧔�)�ŭl����sD�ܿ^��3��[��F)-��n�:L􈅲#�Ek�ӫ��0<#��C5�0���8�:���(gmP���s..�>���Χ�]^�.�LO4�:��|�q���]n]3���ހ��(Ѝ�%E�޴�=����)��X��֕��fQL�7�s޻�.m�P�r��0n�t[y��X�K�80Gf��Zƅ����y�f��Oe]Ѫ�I��1U���s/k�n���ן�����65#I���E����9:S�:ɛ�"��=n��=��*�^V�j��1�c��|�u��n��l���i�>o2��V�X �}c$��ѵW��DC�}Q��#�R-H�B��-�ϲIo7a:A� ����*��<�t����]1f�<( ƺ�"���fWQ��2p�N3{�wl9^w�����l���N�p��RB|,�
��F�*�sI��7�fv�"(��Oh�qi�qU�ʻ{>����6��BLD]�qY~��u��ǶQ&h钪��"�Y��lVmg/l�q� �/���a�s��f1C�w;F�(,+XYSY��Q�	:�]<9�,�C�Z+�FXk�vΕO�v�����d�
���fK��i��藋�<�E��ͽ����[K	vaiD.�΁DJ���N>�V%.x�y��z!�Ņ2*���Y;��9V�� Ɉə���~�cX��%c��G��u���)^�l�?tz�c90'T��3���\y��wi5n�}�ZN�)�i�ل�B�����1��*��?Q�(�"��w5�K��V1����U�㕊kcj�r�㹊뀂u�Y���uǺ�[��W��^�η�������V��w���"HY;,+�m%p"��/����<��O�Ď�X'�^���V��q���.*��Yp:RƝ:}I����G{ܜ�Hs�+����;2�ǝ׺�^��N���&�hke�ݝ	�J��p1��T��m78a� >{Ud��ܳ���s�7����#
����ʭiy+vR�t�M���/��FJi��\��;�!�2�4�Y�.>�_������쟼l����Tw3�H?R��k�:ַ��r;c�;`85�d^ǖ�/m�z��Giu��e�e7aM�w�.pg�
���Q#�����0�������t�#������zo;��l�K�;M���x�g|�£B-q�y��H�wƎ��*�-F%�p�}x�f1�מ;�k�6�����;�
��g��7�|x��Z��b�����b���Fʌ�1���߸�D�=�dz?w/,���vz�]��꼲z��+7}8�*d{#�j��Kmv��ҚD�ᓶv���©&����z��V�(���֕�'�:�˱ݩu�*�ɵe؋��.\ׂN��_;}/5>*�z��1�c��;�p���+���:�i�q�UoL�'��^Y��.bs����<�Nf�IV��"Aq��<�:��L����*Y^�W`��y\h>,k��h$�r��dl��sr���z�@�#��3�*�홉���p�U� �L��7�@;w;L`	SǣÜ$m��sD�Gr;9TN靋�֦<����.����7*��uG�}40:��<�~�к��M�zx��C��+vG4�ϴ������Xr������6;��[��sB�@����<�/w��GS�yQ=i�v�jΝ��z����P� �:� wlު�V��1V����&����1L��w�4j��l��o���w���;�Ki��y���	�Q��Fb�t����zM(�l�O���A�����wY&@���ݯWQ���C\l��U/31��(h�%]��|�"dt��.ɮ���|�BGh-���]�9gaܭ��6�8~���a�G�����W����:��~���ʱ�U�\3wq�ج�����L۷��j�U�y8BS�^���d���0wl�����4y��Q�c ��^�S r�t����5��Ԧ��Ƿ�]����|~�n}�>s�-٤���:�>;����!���"B��5�pEK*�n�"��^h�X]M�rL���������;��?�&����u161�������Fj��n�9jK\��s�I\̈�u�c�.|:��K^ �bGp�Ƒ����F_mE.FMÜ����hc,�2�4�UL�Y�p�+��Ki;�&ʍ<u�a��{c����@=�^���5���˴���/s��*�^�ݪ��}��B޻�))J6:�kŞ�:ӚX'��W@�v���K�[
K0<�At���⌄��|�ڧR7���H�m�Hs�DilS�M�o9K|ּܸ���'k��⻩�rep�9o��UY��)�� M@��*��`��R���;���E�Nuo).��լ��ݏxnu�1o��mJ�Cbk��u�w��ꔮ�g%�R��u��dJf����\��i��b� �oA�����Z��0/ZJ�q{W��x�w�2�0�yW8�lN��b�ǧG�����A��x�HN�uW^�UNb�1z�̩k�!k�텱]"�L֭p��c�<K��ޝف�ᙙAW��x�vm�ַ�o��Q�肦��d(ۆ�L?f#&d����8�N�i
��=���#h0+�ل��m�O�A�ߵ��w���q_>k�����:�_H�1��3���ȭS=H�0g��m�HI��j[\�&���ڢ\t��5@b�5>Kb��YT}��Í#"t�8g��ѳ��p9!����=Y5�k2�ѝH�Ȇ���O�}��ц<�C�#Hc���է��TU�*x��5�ju�/��'B���#_l��.�Q��^*(
�F�ߢYK����њ�KizO���<0�E�}�|��g9;z�<�����_�G�
��PPG�?����Ҩ(#?w��@�Pyj F"��,c*�Q����e�-iY��5+i��m1�6����b�L��Q���,��,e[1c-i��̶ًU�L�kf1f�J�,��S%���2em�ԭ�55�e2fem1��Z�fS)��fcV�1��efe1�*ٓ+Lf��Ɍ�Yc,�mL��V�ReVf�b�k2Y3[K2ڥem+56���e�1c+i�)�+i�MM�,�j�ŕY�2՘ԭ�f���J�m+-��e��i����5Yb��jm2�����eVb�V�X�f��1�ZVj�R���պ�k1�k+5���VWJ�j3[-E�XQ��E��_(�����VZ���VU���Y[++ee�����ee����ʲ�������Vj���YVV[ef�`���6b���*�͵T���+6�R��� ���S�H����U+-�R�֪V[j�`("�@b���
�+*�J�کYkU+-Z�eZ�Y�����R��T���]ڷj�J�Z�Y�����R���Vmj�0@ 1Dּ�yZ����֥eZVZ�f�+6���Ҳ���تA�H 0T���Vm�Y��em1�-i5�"j1��Hu��f֕����ҳV��
� 1D��YV��ZV[ib��V`HQ"1�s�(n���� 	UV1�O��W_����?�o��?����?�{������>�����	��G�J�����=���Ƞ���� ������UD_1��� ��G����?\_柼���?�ڊ *�������������W�o�&��?�?���+�~��A��}؂*���J���Z��5*�J��jl���jR֛eZi����6ͭ4�R���MZZ��ZU��miSV��D� H#H�",Q�i��T����Ki[M��R�[Mm*�eZm*�ڕ���S[+iJ���6ʴ��-��ڕi�i��T��6��Zk6�V�M�6�ZSm���i[F֒�J�kM-Y-hզ��-b�J�5���Lְ�?�DQ
���)
5��֓m�5����U�j�[L��Z������%��~��?�*
Ƞ"� �H (�_������H�~�`������ *�~���u���~�8pH���G��=a�x�}߰� ���P���u���9��V"�
��ă�}�UDZ��:�"� ��
~��(?���=	���_������, �PV~d?�ߟqPW���{�{��?�����������`}O��A����PW��?�?��
�
��oC����$O�~����	A����~��|��s�������{?$��X}��nׯ�ί�ETE���}
}�TE��/�{������	���e5���HQ� ?�s2}p#��<�!J��
{b��6�l�)6�m����EA�Z
�M�m�j�T���4�e��*�KJ�BQT�%E��Mm�ڭZ��hV��lhf�%m�km��f�H��m-b�Y*J��Dʲ�f�bխ��%��j�ԫ4��!�4�2�mi�UMV66VIf�ݴz{�Y�E6��-�*��٦�Zֳ4ڬj�em�RP�H�Y4h�m��m���kZ�LY�X��6m53���l�V�����Y*mKb�i����ۻa�����gv� �Ϸ�kʌe��7m=WwA��omZ�Kz����Rj�[w�OSj�Wr��yևO{�����
vջ�édպvf��w�
�q�Ot�u�@g{U�]w*z���
4��π 6��СC�СB�w�{�P��hP�B��z�
 �P�Cяv�M�����e��<�z���,��r�z]�u�w\Ҕ.ހ�v�K{,��:tt��ooT��ȶ޻jf��Օ����kM1��  ���V�r��s�W���ݗ����-=��ӽݱ�SU�vݷ]n�ۮ�sN@׸�n�������Ǽ�Z퇧�vU�8���@�n��K�U�K�w����u� �jPci�KM��5�>  �P�,z�]}�=5��qJ4Q�tpqV۪۵���mۣ�V�V��j�5Gn� ��4�ӱ�nZ��ݼ�limb�zݤŶYmA��� s�m��hQ�ݝu����U�]Nm��Z���;�C�9�:����T�]��ں����n�r�p(���U�9ݵZ�7�R�Z[f���ViTV�  �}�uV�7v����WAʖ�����5��N��ȪvoL�0	���p�+Z��q��T�(�4:���`gT�4�X�,UTfm�Zπ 6�  q��� t8on�= ��p  zu�X  ]����]�j�א�W  �=��<�@�8�����
��m&�l3j�6�Z�� �� ����@ �x� (P7r\ =�j��  n�  5� u& �a�p  �� �7�/le�ll���m����� ���  Nu�� ;��  e�Ѻ]��h :a�� �:8�p  �\ z 7{m�t ���@��6�����f�*Z6�����熀 {��  �y����=��� ގ�=i�or�  sww4= n�� �  ���^�= | �~@e)RF�FA��1JJ�1 ��d%*I�@ �!��)F  &��*� R!6�Rh  �O����u�+��I_�,�+��'�љ2�c�K�����G����y�?Y�����h(�����W?��D O�ADE���(��� �~��>�+�ʿ���
rZ��;,eI/(��Xu (*�7e���`x���h(+�5��4��Xh�a̼�S(d�F��E��o@^�UGu�d͒$n ��S~U� )dT��h���R�K��jVB(S:n��TB]m�o.Pv�K09WG]��#f*�,8�BS�Q��������W�n#E`ɻa�h�f#�Q�d��U�db��J���C�ݠ۷2�ث�;�I\q�ÿJ��̉�zm�ػ`�/A��f�����N���k{�Өf9��5b-c	���]�R�B��gB7��(m]  {ĵ4B���p��� ������,E��Yy��̻���Jar��^=�a�.���N-�+;���L׿,�ǷfS��t��u�6e����<,�]�@m��nn,Z��i��˪��0�l��/��B�W*k{%ۤ��B��;��[L�wt���5�Eee��jTW���VˀC��ѡn�쳲ܼ�&*\�����Z��^�w��jM�&���Q�� L��^�
�E�<g쿥�62���)��Hɻ�����I����h�!�"]
XH�͹s��]�2���O�-�Ў�)�y�&����K�4��O$EkYL:U���b;��J���L{Z�e�C��*Ί$���9}�kOL��e'�m�8�U]˵i�%:8L7Y#uyx��k�'f���Z�2V^�c�a	�n�R
n!t�B��ƛ�T.�a��$)�ݵ�N8�c̐ ���ffI$��j�ӹmYa��VՑ������l��L*4Xm�w��ͷ�f|v�ͤkT�L��]�{L����wm��B�ѩQZw��y&� �e-�t���kvV����%�t�bu��KV�iRh4hzP�����Yf�\:7 )�ѥ%*�5��GVU$�]1j�VF��%�u�-�.��;#Z5w�&�q�Rt��3����XK�Dz��K�Z�ݱ�sg͗u�`��]�ل�c`�*ُ������F�I�R{a��8e�AJܬr�w��3 {J2u�����sdi��"��oe�Mv����ٶ���K�*��u�L�/�Ͼ=u���6�􀸽F��U|˭k�ê?tX�w6��ɍͽH���U [V,��vS��ݦ�@r�m��4, �3$-�=��-Ghm���ʅmV^Z�F�k
ڵ��Xl��&/��we�{��ݑX�@YG���bV��R�5�spZ�һ�����#�J"�]������w����QU۷A�F��]f�Aah[H��P��e�^�J�����WzU��L�k��I�b�]h��x����(ZGY��@֐�[A���Tm�wy-��(
Mղ�ݼ�JN:�e镶�\�kO)�sVt0��:�H=�oD�]�V�4����rK S���-QZ�V��Z�h��A�x��(��f���A�{7�$���i��r*X�D������{p�ass(@�W�dC4��جlv�*;���͸��u�ZP��3e6���t�f��M�{tA�ssp
�u�Iu�q�j�Tڰ��CnY9K�K�s3�2����V�H���j����,��q�˺�U�͕6V�Pj�yJ�EU�tсli9g,R�V$;cF˭����Қ"}�(Z��e��#+�.:4��2X��k�C���Ҏ��rX�w`{�:4��xw����7n�X�)��m��Dw
�T�S���־���w�G�a#rS7[�c�f�˗��%ӺN�y.�0��}�'l*a����ͤ.<=R¤2K��mm�2���m�ub��(��<�F�єo.�&>��i�sM�k�L�ƥL ���hT"�k�mGj��eI���i��τ��(䧪�6[����)�̛�6*�����r��
 �e\ٲᴆPd���Fa�����D�2yMݖ7M�m'���%*hϭ����F&/7t�9��
޼{7�0i����Vs,��}]�\�]�o�uh(��R<��Q٠Y�a"��{�fK��@m��W������W)!0�N@s$��w�+FӴ���t�}e��۩��'ơ4�`�;"�P�H�� ���d�p��yTX�b3/T�u�e�[�3���X�1����4�����G�h2Ĕ0i." ��w�c[�xI��+dj�n�bDu�j��9*I�b�Olh����ެ�V�
K2+��c��h�ml����ZT�u{+c�.逫m}I2��2��J~Zjc�B,
���8.�,x������-��2�`�l[sF�!`.��Z��溕�Qt3 ��ڌ䛠�i���MtA��Jt��y�����

ln��:�ٌ���'�;+5��ٲ�U�:WCVP�lY�m�2L����W����rQv�6�d���l'0F`�����[z�9�H�!���n�7jL�/dFN�f@�k≯�Vn<��[�j��tu+.��'%�7d���3B�l����W%�� ݋ńXGr-c��(@���PG�,���u���YM�+q�V2,��X��&�1���
B��nY�Z	Ix���p���%Lc]ͷq�ǃS�^��[P��d|�I�RV��b��!�*f5QR���W�<n�4����dw�GdIg-�d�ƍX���3i�-��ke�lˏ3FH�\�LG�aRȲ-�Pc�ܩ�2�9���:o���cUp�W�V�m7vVRb�@���t]�n협w5�Z�I��ьݪ���f��U��K.�v>C.,�WR�Z%��tr�\��8���`�����N��r�^�gi�v+]#�&����ެfn�<��-{Im=qyEHK�R���fef�Fr]�t0<ͬ&��S�;{�3)�Ђ�[t����h:�)E�I��,Ӭ�Yu�V�ŹHG.�\N��ef��j�����}-���-ʍT��j��)i�&612��t!����m�B�qh��r�s�}N���t�U�{�g*��(�`�x��&,0�������,��읿��D.S��=�0TaJ̀�&�v�1Q��0+��6Q5��H=�;U��D��O1��F]�q���DZ���N���l�=צS!i&m���x�:r�\bm��a�l���a��iV�w`�awi[-R��ڟ�L��2���u4���+\l�,PZ�Y��Lqm���b��4BJ��$i:yp!Y�Hsr�r��)̣/���5l�0�N�r���O�xv�� +�:��e��f���-6�YU!�Fl��Qj��uXXF�O�^X�o)9X��HF��&�5�.U�y5���ux椭뿞)n���љ�Er�[hU�-7 �J��V���Aq����y���w6���%��{R��1d�hI�_� ��Od�i�a��>w�NVd܎K�jXs�����T0�Z/1�*l"�ɒ���,,("�뺁@$��P���>X[Gxc�t�S#2����٨G{�ɗz Ѩ�.����r��Z�չ�+;�<�i=d�Dw�μ�KZӋC9�X�xu��[���*qn��Ml��[��,e%�'N@�W#�B�uM&������Q�(Cz5���5Xb+c�,���V��(-V��XՇm�6�\�)#�(�O\�p�]��hm�c�.��sEZGL'�Xٿ'NSoN�H�Y�[%�M��!m]捫-��*�r�o��1������r���f#-�%)���j,H=Q�v<�w�m��Rj*N��m%��RB��2� �qnM�1j
��u�7�c�l�/N'��!�{X��H�t��RE[XO���X�7�j���Ou���:3O^�;y���Z��u�ʍ�Y!�,�Gz�C&�tU%Iu��k�g�5�0�i��Y.��TUL���D
�uw�� �J/�UBSeUfE�Ս�\�A��[FU�(y�����j�v�*�Y�y��Z5����$4w��@�t`�T�fE��a�li��Z9��,��h]�'p�&�Ea��D��^^��k��I�r|s:���|�(��a��[��
|��	A�K�� #��O,�k���I�n����p̖��ʉgʉɇ�
�Skp��$+h�w&j��^д-92^��^ۅ�|��j���XsL[#r��mK˘�(v�&L��Ap�ѰV���@`&R#�7X9Y�@k���Yu5�z��ε�,����J�RJ��Fpx��&��mG��e�zΖ����b�5�{@}�q�
bE2�� �4�ܚ��$m��-%2��@�H���b���l���+R����˙Z��1���w�J�!C�׍��&D��f��,�w�l�Q�>�vP�
N�Х^�^бrq�&Č��QH���M���8�f�G��J�iF�ʁ�͎�ŻW[v�X��Q;�kC2�;���D<	@e��&l��J��]����[ۻKse)K�o,�Ȣ�ЂCQ��QR�"�f|V��Ō���^�t�f��^*�|��M	Y��������a�S�N����
����/A*̊I�%�4�вDƖ6����u%��F^ͱ�j����Ɇ���;V����*mȂ�A�<N[=�{u��&��l�uaͽ�D�k�,�M7�xك1X
k7p���I.cқ:��������	0�������ᘫ�D�ư)k�T�M�!AS������F��4��=�R��ݽ�.�1\h�ӕ�3h��02�7#ouCC5�5����U6m+!݇$�W��q��d7uQ�^%d�	��Riu��*��+-He5��	�y��)��~��6�@t�����%�4�`i���*�p@����^v�F�5�P�W�T7(d�NP��d��DS��K�K�� �D��k�Q؋p$��de��j� ji�^�AVl`Ҋ�spG3 8X��KM
Zv����d���j�,4�!�th<YC6`4(܇�� x5�nSݙHY�X�5`=;d�a���(�{�#��f�ǫe��w%���	.o�%!-F˩G �����L��W��1� ֧��J8�gL�M�
��f)�1�+D�3&&�l˄K+�M�%8,�Q�z�7eہ�ǘ���8M�n��Ɂؘ�ڕ �wVR��b��R0��p��f䲳,8�\l^��b�k��̽p��.X��u2YNm�L���
4]�K3oSkq�l���2[1Ez��v��s]�TM�Ǹ!�[v�*�����)���W�s6��D9j�,�QD���W֒r͕k/[ӎ�0v�,u���5����Cj��9��U�,k1m��m��� �f��U+ʶ�@���6#��4�m�8��w��"ɷ>�ؑ��h�m�zf��5�����q;�S�f�YF��:V>x�P�C0���e
�IjUt�m�#�FU���WN9,:v��hdƯ5F�>LY��f�dJ�̙-�i�y�We)X%�Ak[z�O$N��8���_[�d�Iw��c.�ѡ+��KcR;v�s��|8��
T�`�1�h1�ȖՉ���J��E�\��kkM���h�%fPm�H�4ë)3`�n��!��ۧ[V6Δ�M�su������V�.<Vwr�&�(]f��V$*�r�ƥ5Y&kR�	�!�J����@#�����U&�����v5g]$r˩V4�v���f�HB�;��n4�D�rշXz���Y��{��&��7ZVݧ|��I4��(��iS���3s^��XI8�밥d݌����q��n3���$�%9�M�R6Q�,!�h��F���F�*\aYjGQu�{j�+*���i-���m��滽�tƜ����L�j����G![�	���6���XM�e'7B����&�Ch;�7�A�d�\Re,f��5s�o��D;7v8�
�>TӶ]�;L��Y�N��J�l5s2��e&��(�J��/30L��<�*�Y4k7up<A[ZsS�yXw��a2��X+�j�p��H��Ğ�R��3s0�9 ~F�����&�t�ZsVX��B��q!n�hz��j5J�[�gnm�⩌T��&�A�y� ֝Ϸo7[z��5&����ǧi
j/s 5���ڌ�Cc6l˪A2!S^j*ά0'O5��˻C�&e[L�2C��Z�-�V��4F=��}iamC�r��!�<�� ��(VlkHx"ߢ���u�u�7N�b�a�Ѷ�`�U�ä���%d�ӻ�n���o4A��;��iÇv��D�+,U�Pa�j�77wrK·d���Л*@R�[fķW��*���wEf �����[Q�uwH@�<�'J�1�2��]l����eZ��r�N���kO�\\��k�e��+�.����ԙ�M':�m�`JḤ���[�Xt�I�-lߢ@���A���#)=*H�*�K7d�`���oQ;p�*U9�ح�c��4��웈�bTշYKg#����V��VCL�5�Sv[�`�x�J���X�w^��p���&d:�Xp8ŭ�G�����M+GƂ�p�h�E�9�f�ǬV^k�`W�|Rd�<���ù�h�.Žy!���%(�oh흖��eU�VʧW���k������ьm���v�!�#w�jbN�%VE��V�t"�)2ٛu�m����k�f]��4�(�(�l��Zy�
�跱n��GM�Rd�V�:hf�eZ���U��0l)�B�Cy�C -��'3n�2BnŨ@�d��T����K�zAO2�mJ��˺I=��yLP+v���զ��Z%�����SI{��m<��6S�m�E�&�.{�o�9�+\Jc���6�i��ŕ����J���e��_3n鯭�ꚤk"��;���+TԜw�c_[�R1.�k_l�B���f "�Jzܹb�y�7�'ڱ�)�Ơ��]&��{�_�ϲ���hY/ek��'";I��]�k�atz!"|�n��V��+�]�*��zp���i��S��%M��Ww�@� ����a)�&�Kw�mv:�Z�����l�a%�om�+y�lM[����ľ�޾�E�l<ʚ�mX��I�үpV���)01�&��n�Rlμ[�a��6T��999�rj�R��õV�nљ��@���k0����تQ��0�:�j�KB��\h2H����#b��s�CL��c�8;�mT��ؙ����J[�3QG�dm�E$�.Tr�/���h��/v"�J�W��lWr���݀JW���^Q��c0q�Yw��p�O3U�"u��zUn"�����Ӯy׼$̦��Ђ�\�VQz�5݆+�SF��h���{�+"3����[49��:9}Ca��{qw4H���{��9&/Aݗ��D��Y"=��oR|�yϻ��f@�r���x�I�[|��Gʻ��0kh�z+v�]��.�G̥]n���� �#���o+t�����ڊγ`��.<p��A�Y-۬�2��̇�B�P霝�s-n�3qU��H�0)f��M:��w���/�mc�4`ݽ�dU���E�1O���)Y���v8'2m[R�;+�^|��H�5e)�M�؏�b�U��Y�snJ�ԡ�K���bZsEc#����e�:��_ {4\�h�Jξ���E�y;M�w�T�î�a<M�P�� s췛��}}vA0��$[JY!�ywǊ���r��u�+�Bq��9-�ή҅�y�D0O�ԕ
buN�Y���K�̂.r�m3c��S8���3-vi}�W`d�w�Nr>�q���C��o��z����[yw;@����)�,S���4��T��^:t��@������+h��R��ܨ��g��p$#$��4�i�����_gM܍Cf[��9B�oTT�J�-ʱY1t��ؾ;�bA�
�)�Lj�4�h����5nYkF�U��]��s�t���RwÜ&�Sr��W+"#F'BV3���}�RGKA]�m����4O8il��%�ۢQ�.����s< ���7��{���+.�瘚�n����8v%NV����b��W*��V�Cu�rgήb �J�'�o&���Җ���>���C([l��5Wn�f�6�uj˳�g���L�z�a�����OJZlv�Y|��w#�@J˾D�{��q�.qsP�ٗe4�K�em0���X}QJQ��m*;�}�%�hMg�'E�A�8.륝5��3VR)���|�γs��G�(���7���,4�%u�Kg+�C�:�5�-��8&��L���Ϫ�X�d'Oi����-���f����P��C,���#M��.L(�����Nh��AF:�o�E�|��0$1RM�I�����y��p�*�Y�q��#������3�]V���,���ت����ֺ��Q�_ڕ�
�ˬ�(	�:!�v�B�U�]��3B0ݥ�7 ��b_|���z�����;�HE��g:�Ό�\*�ޱ�/E���9y�4�$��f���]�S{�z��eY��=�-3��7Xg��k]�=�mϓ7�z"�_��޵�-#�*��l4{���jJwA�4.��Մ�;�
�@Q���r���� ���qQ|�3Fu;�v6@���'+��N�kb�z�WX�S�8��҉ �CG3+k�X�1��c@=��Eu����ʗ�PjY��s���.�XS0l�{���3��z�K8��T�����/��Q�H+^̍�z���̽�,�ic�b\]�Ǽ.��i�T�t]ys)lK�5�*qh��ۡ�//eKX��P��w&"OMR�r��(>C��
�+_LW k8�`�Q
X^���Q�P��3uZ5�b����j����6�hʽ}���N�֕�gF�I�D�dmեp)��v&�U}&�jB�YJMaCMN�����<Wu��&턕��/P�#{i
ņ'.����wjӫe�0M��O�g�<��%�z�]�nSכoz�g.
�h�.՜���,�ܸ�Pf�/![6�ղ^ޕu��Y[�N�y����Zfdy��$�\sm��/6�X�\���4�2�k�� ������ݔaʠ? �w��T��IY�Fx�%�W�C��*=��w;����h��wa�EM�A\��02�۸x�Ҳ�@q�|��#2��x���_&˹.�@=�QZ���Tً1N��8Ʀ:�sQǃq&lC��;&5]2fɗjs!�QIz�8�u��kGe��]B��T�v�xʌ}�m���t��nO���{1��Y�ʒ����Yw���pz*�B}��y�[Ó�,���[<��5�B���Un��ܛ�zsɣ�T�ʵe\n��B���zFM>hn+�\s�p��gc�Kc��}�["Ѫ�o���i�̮�ƮwAW'n_Y����fu�l��hmќ%F�5�����sT��ƕ��.�t�J1Q|I���;g-ø˴�7Lv����r��BnE�rt��T��j�s������\ٲ��5�:�:�|F<�&T��[��GӮC>��)qaVw�E��0b��.3^�;��a-�ۛ��43�A�/��C���>�szBō<�[���V��ۜ�W^E\(iY�K(+ӭ\�b�����j�,�h��͓��F�[}]����f�K�Z?�����O`��Gs�he�������W���r�W�u���M`9��Jl��V�лw�ޛ�7,��H����n�8!������8�X \��B�-�xEp��b��t!u��\Me�
���-�^�y;o+���`��UՐ�G�¾j;As�K[C���Mغ<��Y�L�E7Zb�e�%2tut�}NN`�7����<Ut^�B�#����P�:(gc�l�	5�\��>E��J4(��ܛf��4���z�:]�c X;m��k���=��id�&\����g@0�5��	G6��.CFk�;_T�3�L�[�tn�u������i��܄���!��eZ���k�g0��;q�Oq���:;e��)��\�X5�{�x���y�����#ϓ��j*�r�S�x�ω\Nf��&�
�3���`��(I�[�L���u������B�j��A���9��Zd57uV�ɺa�aT;��EZ����ܮ���{reY{t���kt�vԳ	+���i��A=���w�)i�R�Z��u+.s��ju�	G����;�b7)>�.�H�:��mgorTeP }��f�-2ʬ`���y�<��	'�e��p߱n��q��f|�'	��nfW-ڔB/3h)0u#���(dҒ�ox�,�wWƝv� �Ӑ��K����p)t������ku�5K1���qu8m˷z�N��4����ĨaT޼J���uyc4�,6y�C���c�9�s	=N�nU�<�byڑ�`���J�w���i�[ɹ1��j�D�����=%���-����C�u�C�[i�&��v�7�����U�R�B��v��?��+&)��\�A�!X	�]N����v��>�9���ٌ��t�V릷��+��OGa�m�,��d�N��cs;,�*�nuU� �3J��@�zX��߶�N�������њx4�k�b�ren��ݓOq�W J����	[��Q�j�a�	m>�"��F�Q�Sk"�y�A�Z��gU�F�E�iTgvΰ���d�{$�P��C�'}��`���f�9�����.ŗ�?����vFЋ&��fe�!��LX̕*��bT�2Z����s�s�g\���w,^%u�֟t�#gt�W^iu�bۆ�n��ͩ�i��Ѱ�|�Xb[1>V��~�Mu��G��e�Ui��36��ʊ��B�aP��2m���u>�����Ω3��B��Tл�@0�!����f��J qyg��ܠ@�<:�t�u�/�.@Zf���)Kj���{{����ب�����baz,��,`�Z��j��׷#&��T���b��@�ޥC]��y��*�� 4l����GR�gx��Q�˼fw}����gB�̊�������*B*�Ĭ��3e�)�W��IP�뮒�ڔ�(�NW+(K�n���5�:�.����״"yc9��ˉ�1q)_N��I"�<<�H��M�>�a˭E�gy�9p�[�|f�N,�����,�|[� <������@�muJ��2��KBǼe8��:�7��*�;HD���8�h8���u�n�v�s�Sa��A5�l�b�;�͗�2��v�vFԻ�h�F�����XEbS�X��񎍹�4U��ٍN���7��yO���v��ĂtM�
y�b�\�u�(�Wk�k���[��A̰�B�r=
p,{��S��ݼT�H������y�
�x�+��X��N���)�ܘWK��������r�/�eښ�nJ��U��\ݹH� :"�w�Qv�ݙLj�m����A������2�P���輭��"[��hP��2\;!ӷ�i�F;�+�|��z���Ĕ%�f���L���æ�+zȕr�kS�+Q����+6^���;�e�r�n�05Ѻ&p*
�]dw;�=и�\SD��8R��W
P��h�fM�֔��?��ﲄ//m�.@��3�,H4�f��[�����N3�C��BNdU/$52�e�*�BLޢ��Z�m���JJS�H��:�
9R�!�kx�[@n�W(L]lwm�Z�2�UG6���E9h�����.ĝ��S���笞3���5Lj�q�蜘�VX�j�.Y�a�ׁ��T���|&Ye�/fI�.����0(�ֶ����V =��j����yv��wPd_*}}5�� �*�W++�s��%�#uhN�n�m2p��1:�DH�g�9v]*�3���g.'s]d0���K�O[��"���Rf��R�ۆ�K���a�R.��YN��``�z���yv�}svlSN'��<�	���v=����k�E�V���\7@�5,�\gJpf����K��T��E���M�ےg]Ͼ�ל����!��㊷�C�y !���b{��0vEo
Ŏĕ4��3�V����YǖUgm�z�\��n���mALN�He�!�iʱ[ɗp�\�R�sr]�,� �g,!b�*tG�l��WE�h�2��=�EZ]���K����Q��� ��Ʋ��ի;��Q��#j i�r�5����t�ЎD��+P`T侵g+�ӥх�n:�����t���txބl�����)�-vt��vPW�^�.�sN�]]�<����=�:�͞J���j�B)*����<X앎�wb��Z�w�_=ZiT�l����s�|,ua��紞ƭM��Τ���e��ju����k1.;}&��ZPVT��;L��`�֝ޙx�(��J�������J�,肳��a��}�pb���X�r�`��O�֭��U����7�`�E�n^*
��vSb~2zz�����>޾��(�@{7/D��v�^u�����Q@̛N������g��[Lǋwx��k��͸�F� ����m쌓���־�Ϻ���vވ �!�*ļ�Y����-g[�]pH�7�����).Op�D%�Ƨ\�n�Iz��N�G��)B�����p�Y���fM��֦F�P���-���t��KT�:*�v�e)�s�G�����c(@a�l`�]W9���;A6�VQ�-6�Ik�z�IN�k�]qA�l�uŢb)̷��r4#3Wj}���=�Yz�<υ�Φ�r�ǚ�)<��1����ƺ���X�M+�I�h4�D�������5�0EzV@�ҵ�� �7�t��B>�EH�ِ1�,U�-�p��ϴ%�n�W�k2�蔢%�J��%@���x��{=��i��9�%v'��XY6�_e�v�! P��k����4�g.�;K�J=7��n�����B���x��<�'b���}�y��gxl��V���ـ�' �U���^ը��V�t���]]ή�G�p���@�rΞ�(k���x�m�܊躵
���G�7�90$蚷��u�P�u��7�nH\�Vn���v�-vB�e᤮�u����MNe���B�#{�uk�F^ŋ*C�u�y�$����ݧ��e7µ&�u7�k��
CM�̟9$�,��Qo���E�Ǒ��yx1���H�C[F�o�Ky��e�Y��[��J{y���vm��������C[�nT�Bт)�.N�` Au�*V���v��a�a�����B�O#���V��i�Xf�=�r����5��O,��4s%�Q���[�5�z�d�:A�A�&^l10��j��j�����f��d��u&�8{'"wU���}���e��8��)��l�wDWS���P��k�2�XΏ�0AvU�8��LT�6�W��qυ�Tzd�� 3`��@��v:�3{�����mP�QZ]���F3GNM�BH�U��V�m]�3�o`�:�⒏1����`1r�1��s2���4��%aeX�e&,�P��2f>��B�n�6�M�AW�9�>�T�m����:�J��מ[��G1��Rk��� I��sD�&�e;]�״�[g�Ӑ�gfN>�ۑPhV��z�]l\iU�H��9�����`�����n)�2%�_Qy,�S������c V�s+�=TF���S��� �/)��;��j�=z��Xw�%��xnMk!��Ԭ���'v=}��0żt�0qMI@�br��t���q?L�[��zY������ 
��������6��{��Z�u5AL-EK�>��l�1��]�N�`?e^�(��	K%e,ǘ�W0w\q�N����-��Y�fp�����<pm<9��
�r�uha���&�<��p����:��}[��]Z��[�0lU�./F֧�\�sZ��5Ɛ|��|����E�y�!]LT{[(��o�ՙL���x'i[�+d���uj¢O������+�U��G�9^��.-Pl��_=*�95�����ݪ��9gZZ[��`��K�r�q&�`w#�%j�l� ��3&|�<�%ɯe<([���4*;�Yv�)o"�gP�6���ut�\�	\�5vP҅����[��=�;
�[��S���b͠&5�������[���,���{j����-�V@S*���
ߎ�� �����P�c���S����lM���2ї�t�Y�c�n%�)+2�=�o\��2���U�_%}LY�@�@n�ёn�֋u��ʻy{G8w-��� Q��)��@�f\ˆ�Y��eg[��`e�5B"��ܝ�E�p;�@���#e�`>�sR�kT��ZU�E�w�2nS	5멁�>)��#6u�դ��PIR�^m�V��ٗ.�����������P��2�ʘ#j7��1}��fR�[*Gtܳ�ltqޗ&�OL�Da�%�j�.[/��VD<�e��sn��Ž{�mE9�q��w���&i%�F� ;Eu(�}Y�bz�C �ʀKEvRZ�B�&���3X�c"�]��so5���5Ѓa�2Q2X�qCBo-Wdt��KR�Z�ޔ*�	�N�V�ﰱ)o=Ph�\x�&���\�/Eӻ]���ݔ1Gؗ O��V^�ђ��A.^��u��kx1M�d>���	1r�sk�9���*�1v��y�U�#��i��x. ��y�c����mZn�Bh�1����3(;Eh���:��v����rv�솕B�lG�Zb�b����	եQm��ά]	��*�˅c����eu]��3��&Ǹ:�L�O`�y�8\���r��x��"S��[C�jv2������fNMh�;e�X��v���:=(�.��hn����ۮ���̬��`�qH$��m�Z��z^�{����^Ч�������n�����-�6�?l��:����a<���kX�K�w�VVeM]�ǰ�&z��mC-�ܶ���`�ٖ���[}O��ϛ�[��ϱ�'O��i�p ��d��kRŬ:�]G��}�+�ɠe����Ei�h��VSOLc9ꗻ�v}���#�,�L�ӆ�[���܍oQ��d�aƹZ��qt��E�W�f�Ff�V(�H�e�ކ����T����5x-w�bi� � hӭ������*��� �"&����ך.��G9�QKM˵|����&���Ts����)��\kzT�Q��:x5��.Kq�y@�'�Gi+�C��ٮ-�D8��]p�t\Sq�2���1J�J*,\�#d�[,���h������ d�@�֜7mds��譖��#��D���b��ɸPRj�m=�f��
�r9�̠��.�S�[����|��H�2^_��.�G���B�OU�d�b�H��z@���n[ׅ�Dbܰ�Ik�y3��`��y��I��L�NbX�h�gM涳5����I�H��հL���V
��ݵVm�Ί���*��6�qv��hΛEU̓7靏��yI�n�KN�i&�u��������}��g���/EJBWla��U����J�C$T+-�Ы�2��D�̺����N�n���%��p$!Ý�"'ݮ��l�'��pLu�k��:��*�"	"�s`��p�e��M{�0Ĵr��:n*�ylWش�W��׉:0o'��R�2K�q<͎Q����z��*���#�OG[V��R��'7��1}�*�f�����=ÕW�\ֳm�!D)��WZ�"��WR*���7`S0�VV30,���s�g�y���X�"��^mnɎ7�7:��c�\�
]�Z7ؕ	pλ�Ē���ɢjQ�Des�p ݜ�ve���{LU�tȀ�Xs�rp�9;:�9 ��*��]��:]�`�n�l�w��7':��=P�Ma���}��K0�j5ϵ6� �;�K�!Y{�ݦ����l�1�����9&G�{csZ��Y"�l����4y��ROG��ve^��kc�\�4�=�c���`	���͠�,҅���d�Ľ�m����m`9�w�ce\U܌�"rĺ&�@��2\�G�>ՖA*IL+��+����D��-uYU��9iE���]�ru���3k���*���٫yX���Mr�u92o�*�Z�؍nI�Y�qCwuHĥ��r{B�tr\r�>��A�u+D5y�1,_Z�#ô/�%ٻQӉ��`ѝy/
��\0�N�։Ŏ�QR\f���ڼW,��wNRHQ�.��S���1�B�Jռ'el�iΔu��()�����<����V8u6l��U����Ye�Ѽ�'b쬝�B�i�r�^ǡ�+m��pQH��P�OF��We9m�kMf�+X
���%��Q
���2�Ug�����׼�rN�e�ؕ]��&�O�vi����[F�6m�5��Ί�[{�]���h���T^�R>�޳��0����)�g�qĶ��':�X�f�칎e4y�.'4����$�\$��wf�ޥ@ek��Aѩ8�V���9.��-�U�_CBo��ϰ���P˶�!,QQ��$5��Ftcb�R�Y��j���.��&%��܊���<
����Rk[��d4٭�z⚈�4�\�r���Ŵ�T��}K�JdX�2�� ��t��]�ui�嵺y��RsV�KR��]������l���k��S&����iCj�Z��O�"0d��+�7�Y��I�[7nq4��1��/�j��0a���1f����w�� �\ ��hKW��}O�B�u�WS�L7G�t�g���k��t�+B
��]�����.鸮������uj<]�����ո���=���3k	�['v�y#���q��k�i��Ӱ��[۶���;��V�����!;t�e���7qnD�ܣaPY�znoV�Mܵ��
��Eu�i2�7Z�����#yes�م|�+x*�$�]>F�\_`ɗG8������iӮ&X]���7�d�dQV9ΙF<N�`ϔ��<�TVXң��hr���j�Ʌn���V��'�����!뙔�r��pH��4]��V�&��ģ�0�]��=��Eagc;3i<���ݻ5�U�zB�[���zA]o�R�B@uݘ��B�U�i��S��Z�r�+6�8�!]��U�i��l 8)A�op�X�+u�j��� �|�#���m��n�]:;0G+[p�G �z��f�M���=�d�u�]X��R���AYf�"�<�ygE�p�30]�ǆ}�ةl4�=��嘻��x�7����N4f>��dz��w�潌R7��z#<� �G9Siҹ{{q��Ȅ$lܖ�a��>�nd�]�u��.�d<Ps6�j��{�.���I�ҕ��xl���,�mJ�P��w9�ju3mD��d���i�ٵ���FG�L�Z��)�ʋA�z�Y�U�Du�t2wˌ4{ȼ�9t:�Ob�O��A�R� 
��ι��5}\��S�)����ap�<z�6�Č�]��x��V֚8�&9Ǖڌ
nYR�;�.>0���+Dg�7��N�ˬ�n��&7S,t��4�Z��
���H�Ğ�JW��V�s����mAۦ�n9�E�%h�P{��|�Ru-}��7p��e���w+�m���<�\��6뮮T!��9ɗ;�>Vu���+�D9,�����*6j��^�v���w��#!�9cN��G�t��-7�֒[��%u��E���0�s+��i�05vu�� ۫�P��s���W��VE���-���w���G>oo����
��!-��ʴ{z��!X ]���*�>vm^!s��BS�����j~����z�r���Z��3I�*� �pȷ��<�JIBo�#�d�+$�'6^�& vW4.Ҕs	.s��7\x����V���	�`İȨQ���Mu�/���V�j��G�]>¦Sr@+:�1������R�tp��E�C ��41�PCNM�[PM3Jw����2�&�㜅^S�ڭS��s�A�F���Vp�B����p������'Mn^�IF��㓇Н��J튝��ғPT���UCi��Pc+# ;�f]ɕ�(F1�B�W���M1�Ǻ��6@�4�.�r�[�TќmJ,�6P/y��R۶٩�wP}CN=�������t��-˗�MRڳ�r��W���3 �XGWe�����ۻ�8���m����{8��UW�>�v�;5��C�;�73��b2�k��h��������3����z�c9n�kM�B���*��]�U)gA�vػ��1�N�@=��#s�4�]lk�[b�
�(�wa>��05�5��R��:��W�rNU�E�C�s���k�&m0`Һ� vao2�,�/F�g]EP����H�,W �)
_q�pq�;�����lG9����t>Ů]��Q��]���up��=G��g�I�Yߖʁ��0a�.M݇��.��ذoIN�Hzb�(bT���
ʿ��ݗ֍^�{ ێ��+���:v��	%�+X=x���ھ�D���0o\z"��xF@�m�s7Bs:N���)Ư�;���m���F�i�N
z�]�0u�O[u��J��-]Y5N��so�6ݵi^��We�Ħ��r��?ZǪ� �>��u�ܹ����p�⸺m,���l��	A@���뾦�АncU�K`D�d�o�j�Y��F�X�JC[!���s%�������Ov��a������ե`���%��R�7��F*����L�R�@�7���A�4)u�4�#%R�L�f�B�.g��]���OGA⵽n�Vu8主%�9[R��R��F�Tz�˴�/({p�Daneڕ;�nkh'B���������sA��ٿf=1� �i�R������܍u�ܵ|�
��I	u��\kM`�@Ų�5�Wn�Ҩd&mXy�q���Lf��ײ�w�sWgmj"q���Voy�b�RN;�tUe��m�QqiŒ��"ݣM�tL�Y��C,J��-t���i�,a�=�Y������!��J���)�4^��DQ9]��dUJ_]*0No���]h ���Q���q��>���5g�@�q��iV�}��AN�X�S�W�V3fKB	PV��wD*O2m�%�_`]\��d�w}�r��@��gX�\K����Ղc\[2u&�vہ(�R�ɵb���b�4Ѿ��Fq�W��^�oBs[R�����XØ\�~�U4�e�U^Vc:�V���wR��#��΂���E���'0J����sA������L�E����L��'^Yj ��s�B�V�ІQљ�<�b�0�ӏ���*�}�0�
1�����@��IQ4���,�5�l��`S���K��x�M�;�[w1���6C��n�a���C;(ѵ���<�bJrJ�}�o��n���F���G��T]�9��X3x�1��c5�Ѐ�}�J�萇t�v�0�]-ǧ�3i�c���.u����m����
������ut�:0E��1�D��g��iCne���EL��ӰTD�l��Zaݔ>� ��_5�j��:�Y{/^��zP.wl�q��kFtk$�W���[9`�V��m�Ȭ��0�&�:,<FU�j�#qD�X�wwݪIf��u���[������u0���$z3I������'n��k�U���w�c�M��B.�k��"㫆�,���CD�E}7%_=���f+t��f�*�i�׹�����g9��P���D�6��o�z�\YQA��(�s�D��ogpֈ�X8R�B�9�fՇ3��b���i�*Ӑl�EtA���}��sGK̍�7C�u�Q��y���"�8��r^���9�U0m�-R�ʒ����{2�u�S�e*p��S:������qi����vf����fuyWݕi'��)�Iz��ټ���yOf��X�T&#�db��Q�6#7om�T����p�௶�;)��+A1����,嬊&�t:T���Ƌ2K�� ���`U�U}-���o�T�%�8���tu���]b��D��6�[�֟�R]Zq�i�<�j�4[�fQ�'pC�W#l�m�r��pQ�6Hk"�R�fۥ����a�"����y*[�Q�-�+������PmV�6��:��7��v��Q�P���4E9*��C�F�a��V=1�WY����`�Sh΃���KL��ĳ�j��ą4�4�sT�f���]��f�g���ɤ?�E��}��gm�C�x���3ױ�=�E���Km�ªfp�YB����oi\�eGeVn^�� �ʼ��(#��4�Sp�.Q(�����2?��`�#qSdu��r�U���OhM�æ��K%����נ^���h��
o&��:*3Kb5�D7�x�V��Uu��n���l�(���!��A×h�)bw]��H�9���)*�Q斲�a�3�������!/y�:ۓY���G�����4l�¯�}��.b�*5	�'�=�tr��0�c6#��/�[�a�{��y1[˫)����a5/� ����uZ ��;IO������N�G Z>�b����EN8ˁ����Pa����7-�؟a{w�M/13謝�N�yk�ħuV?3{���{��~b�s�w����dJn3PQ�+�N�S���g!�w��M�0�8S��-�fM=-�.�4�����´�hJ�[j�WKMq�"�E�Y���0������0(��ۀѤ��������îxn^�E��n�"!�q]�\�û��������9\���{W[�tɼ�˲+%)�]�kV:�x3�<�}��v&�Z**ԝ�)2�@^m���o�j�,U�U[�@q�M�re��Z/:�!��izA���VI��렖��+����1qE��٢�k4�z����(;Q�-�LL��d�2�P�wl	{A���I�9OJ�}\�΅,��5��Y�<%��靕�]B)�=�:�A���5��NC*.��,isTz��[����-�2Ť�E[e./�����N�AY��]^�Up\5Jg+�A�Y±�Zd�}��֊P�M\�&�
���&Ko��*q��K��69cyU���R�ܖ��ϓ���h����g��]�=��ȶ�ԯ�7JI*}�$3���K�o;`��y�o��9b��L�^%���zn��V���;o����B�[72�s�ymhp�:�wLg��k`1]"���+$�me����=]Y�2���. Rx�e7>^����MQ�s4`6��L����j6%��u�!ѫj��k;\EJ������^s���L�]���g�?yȽ�BR�IB�R-&B(���&H�.A���.H��B�)�H�f`��B- �4M.@RT�H�T�,M՘d�5�f��E,BRQIBDD���CFf)KE4JL�4�LĹ2P�!�U���UU`a*�HD�ѓ�PR8T8NBYcA�f9@4ђ9)KCAE4�K@��FFFEfaAf!����Df%VfP�cI�!BӖKCD�G�|&Ƀ7s�Z�2�6݅���:��_'�F`{��h����I���֟p傺��dk1ir���˹Il�;��1?�Qv��Đ�F��n���̹eٮ\��J�tt�vп�������0iZ�#8o�� �V�ʳC��\
��v�dS�zvs
����[���s�.k<�R���v_��I��}���p1�#j�z�l��������u�$�'�(B�UF\=z�`lz�<~?7���^�vk��׏��^W����~��X�ׄT1`��+�0�ay	.�Ihp���Vvx5خ��k��ɵ��N���sL��5kLX�ɜ7��N7Wb����]����E#����ԥ+{�"�y��1�F3��{�`�-v])05>�J�9=��m�j.��f~�?�@��R�L� 7��sI�1qk"b�q�233m�Ӄ����v�Z>�	0�{�����5�]P����ó�<�f��噮�-�v�8&������3-S�xb��5������u�M!?��]�c���P���ME��F[�oNr��ӟi����M��L�(�RAN�0:x�3�nu��
PTb��o��S�}�y����Xð���tI!9[�C*�T�h�BЩ,,����.NC�ZUȨ℁e�`ȑ�J;0e;���8uu.��h���2󺷝��"h1ú�M�/̼�l����r��|NyƠ����}��l.\25��ɎfS���s�ida�:>�sBcr��P@�r�v�m���@� p\�SP���։
WW�c���q7�7pt�©O�7pZys=8Յ���V��(�HR��w����ա��+��h�n��ۗ\g��r�z�lC�슳"C q a�)��kDa.���^QhmC�^�b�a ���7��5F��uh@�B�Ȅ��7U�皫�Et.�:�G��;��C��iZd˫҉f���q�f�/+��D�E2h�&�xh�O��V�,}���ɏ��	�֛�m�X�!1fq)���)<��nٵt�ٵuT|y���yۆ���s��
� ��R]�����>'�ν�ܴ�4ӳu��V��(��a�Aާ���C�''qZm�ۜ*��d^�,�=8ry�7K3L�y����@�k��Ӄ�._���i\`:��M�(̌��3I�
1���*;�}��HИa2aUЎ��LDw��P����������˛�"�۟�3M�(�xj�wv�*�T�hcJ,sD:�r^��#�w"��W>�iM�n���h�X�����Rhx΃z��z,�����K�����ԴiF���l�G����k�,.�s�|�
5��ܾ�3�hc]��#��u/�H��s����X*Y ��-���C.��>��r�2�����TC��)��ܝD8U_!�S1��B=U�)�t��<��֗�T&�y���ꧮ����Q'@A�1�lc�y"�q�;>�eZw	��0���,���o��ƺ�P3<
��K�u<��вhB�鏭�t�d;M���MP|~�¥�U�q!^��c}Y�A�RP��*�TC�Ү%��J��|�Z1c��ۘ�p����sN�	Rw{�	u=��k���r��h*<�
�.R73�
�i���J�7/�Mk�'�#�9�&	�����<�}�O6ؚN�\�  ��>�`�P(l�z���ѳ���{�����V����u�r��nvF�;�4�$�+�J� �����+KV�;��/����6v�v������&8C��Jσ������t����k��7���t�nH��n�F�`|w;�C�<*LRI�g>.b5�U� T5�䆦At��q�9e��<�����n�#�~O[U�sg9�%�rbɵʡ��zmȆ�TAM��Rv#	ꓡ oCw��
xguI� j�X�m���c�3�:z��)W_ugX�VOR�B��3yTY��h��6���ICB`�|8�����-}��G�SǙ�Z�w��]ȴX
e2����Z��Gނ��9bW�i�_��;U�\>�ɝ��^K%�Di�7�7S\�k�Y�k��zm�R���ބ1j�O&)�hS�DI������r�AP\;�u#���4h��	�b�j.R=E��P���������mA��5t?iUF(9�˼.���'
C�;5(�����P6!�<�Y�5ȁ���_N���xԆ�:���\%x��`�͹��A��z׽sa��!�������}�뙁���elT؍ۄ�x���p?P��0.���H7,������p[��5�.�bc�*����O2�d;��K�T��1�çU�1C|V���$��U���CeG��^��H�L�Dn�f��C/ �`<䶚����sb�]�	�Z7��<Z4���FR�BELG>��D?����ůA��B��2��R�Mn�5~���7�ޤ;"^��A�R R���@��@a"�p5�WrO��
`�AwY���.��tҾn� �s3n��r�/%�Zq�Q�+us��\ʼZ�Z�@��w�V��(�H�ۮ�񇅣L���L=:f�Ddt�c3���,�O7�}Ի$�Hd�
.c=�r����hNԲ�Y-�7e	�p(��W�w	ǩ8\��k��"U���L�\c��rm|�܌��uh�g��qD���J�e���j�����}������8���δ<t�敥3#�����hZ��F�P@���X'2:Tgf�z��1����Ja�P����N�C>rՖs�c4����uZ�qgK:�Wr�s��#�*��{M'���N�_�s��!7\K�X�u]UE�FP#M�v2zOXݿ��G��v�F�O���]�t�xbu��R��e���v�^S���'�>���݋�G���M(��j����񨃳a��պ���+�Qmgm����˒s�	�n���Ӑ�����@���\k��7~Th�����>P8����9��1�k������=��\x�~O+�Q���\�F��'�j$L71`�o��F��4u#��y������E����@��o'Z�F��Rߚ��.�L�3N9��6�*\���}�@�
�
�t0?���ߗ����pg�������*N�N�r,<��6p�Oh#,M����;Oޕ�!����=v��o�M%�u���kQ�A���17^�j��ʓ�9v����
�;�[�k��N�I���LfaΥ�\��Ծ�����淞ڡNlx �-k�t�^^,Z��t�Õ��8.�!��T]��#g|6��ύ�
��\@��� ����缙F��Nz+|���M?U�I�w��Z��b����F����#g�恻IgdϨ�*�2.�v1Ea��&�(���~a��w	�����ϥm�ԫ�Ď�Դ��u��S�z�����:�FǦ��H�[1(�s�����^�!��2~aEq�帍�P8����F�b�i�t�ԣ�=VӘ��f7�%_�J`���<�ë'��I�1��K6o�< >	t%��%��A� 7�� C Q�O�� "b/�h�j�_�<v�� w�h SJ���첫b��;Ѧ�~qf5�q����`j,��#��MZ��0���k��S]�^
_�z�dB^�z�m���V��tHҨ��e�3B��\��ЭTJ7�i�N����CmFIo�0V@u��!
!;���u1`�\j ��%m1R_�1�I��U��w�P*�2;fkQiq��亢EDr�ɢ��5����~���c�T�ׇ�,3\ۍ����3^�x6\Q��W���UՐ�:;(Vɜ&mtnv�@y\�y;w�fbV��}�Ό7�=i�s��o�+�NZ-�����#�FF}�(�ZC�3��|�u�+T��5>8-�ô���Y�6ڮoDvXXq�y&�\/nu.�C6��C��ؗa��z�������N�L\c��5������r,ݯ��]�V���Q��^Y��څd�\0GY���1��"��O�59 �f��9��&���yp�S 3:z�s��I��}�$5쪵^�t8@eԾ��+�u9�ycL��ܼv}�n�8�z�NwY��?-�Bw,�<@$FT�=��J�`"x�k�g��:��I+
�Ɲ8���@q0�>�ok�s���=��5|p�ivEk�o��j�\�nT�Q|z:bJ�z֗:�t�9�\�ȅU�1��G�VI��x���:��!.���m�1Ƨw�����AɎc@�<�eѸNS)ү��*� �<H<EcWU6��co:^*����x:K^��Ԝ����������t�a`3��j��S��u����U*WC��h#���`�(]L�3Ý%x$tB�c���Z1��qe�[�����P�#�$=��5�;jY��r��h#��g˸��/�?���N����T�Artvsh�Op�ufgyC5�`�׀��J�i��%O����������Gq3���,�ܥ/�����۲��X�ElՐ1w&��μ�)��IJ<�!f3[YN�l�j�`��<"n��f[���%$DԇY��d��I�8!��ə[y+8�k��F���e9���uR�� B`}���tP��1�U�����2P�*%�~T�t��ad��b��uv��]�Yz݊N�R'�����O*�f���
�.��`oչ��ĳ�z��L=��[G!��b˜D��
��١p�$Tt���:�!�i�F���z��*��na��1X[5��!Z�&)$����T\Rt,�rf�;5�Y�ź�w�̓�r;h��/��f�{.�\K��� �?g;����_Ȱ�Bk�Ed�|U	K�h�cN{;�ə��j�����:�5^�Ad?]/)�<!���*�YB�ՈJ���ԩ!��_9s�u�/�r�9j���{�HV}�1��C�]<~�l�
���AE�S5�l�̉�����	K�C�2^���=�b����E��PFZ���qÓ�:��xz�`⢴G�:�Q�z��&˄b&�j�T�2q��~����X��X2�#ip�9	R��ij���ܬ��n�=T�3�B$S�<j���x��~���H��y�a��]9C�gZ|}��*¥�2L������\e��q	2����^���w@M����m�\�
5����:EB푓���Y���<����VS�#ˮ<��2�	@*Hd@'����=pF^�1�����k����g"�[����#CVG�.3��.��(
�ꢼ-����q1N�!ǣ�ъ��y�#>w)�ϩ��}��B��^b���������������|g�����)H�PAdn�dk��}1���)�b�j����a]-�l>�*κ�r�D�@�b<ǟ�e,�B��/�(4~Os"���-��[��x��;�#��M�=�C�^���L�)��/���Cø�T>����j�8���q7Y�7�\s\���������
ߺ���$��^�=su��m��X��ـ�l������M����ƈ���\;�f����xr����[��6 �of��Ja����t|�:AWQE��M���Uēk��R�	��5U[�O�����"�i�����VIr��~�uĸ��݃sk����Ԓ�=8ɀn����[�5�rO����N�G��S5���}���W�ٍ�WXo�"믤�X`��9`ix����C<7)n����~�N�a^�a�5���=�C"�5&���N����|����{F&�fc��Cs~,�рRI�&
����T	�>��� d�"{�4��T,�*�;)����	{��u����nn���:�$�Z���&ջ'�gq��x�!¬����N��˹2�s������[[BZ�&ځQ��f͈��U��s����̇3�1&꼨
Ћ\5�B/��Κl�Y�s',��������N��ѯ�//�ޘ|b�k��s�uLOdN���Q�o ���^��g�`J,~Ӓ]o׸�;SֵBc����+���x>oz��k�e-j֘���2��
5;fyF�����*�B�<���>^`�%��GO4�:��y��MG{յѾ_9�=|�JzĶ�E��b=O���QJ@}ci�"�
 A��-���q�C�=o�@"��)��s<0f���b���j�I�	�6|;v���6�mT]��8�����@U([P���Bf�Ln*��z�l��<	=S:�}P����փ��2���iR��"�5�1(�B�oNDs��ӑ��6�5pŕ6��:%�����̮4����-Yu�?�K�mLI1��RU�(1�㞻H�9z�'��_'P�;Ύ�cD߲�ջ<�n��� o��_�� �=��/�y�C�G��Pnw��������q~_>�
��
��uk�����t�V�Ca���8�1�M�%vM|h��w���q/:�Kf�Qx���E��u\6�!�[���DJ��e-"�{}�A�-:'9��ݲR�w��I�2�Y�g,�S��{k�yć�f�a���������ݮ�!�;r��'�.��Zf��v�ݴ!K�LY*�[��o�!���a�k�V�u�5�O+�Mծ�9қ�|�lJS��=��j����֮m7�	%���`�t�� Ω��e���.彳r��P�!H9�k������o�4^(�ꀻh���,��<00������r�%��Wdh,R^p��,�r���R�W|� sb �t�H�u6b.\��5�7��ҥu���D��M��V
�:]p{L�$x��f�]p����d AwM�����8,b�۵��P��j� �Ro�Y�/� 8I\��i:���w��ڛyW�ɻ�&��#Vmm!����]��ܾKjn]n5�Ʉ�S_S#Y	?]�%nX��F3d�9j◷�����ަG1s�+ɣe�(��Lqn�E1���ub�ώ0� �v1ŗ�N�8�B��(q�M{{�G��o7�o�1��C�Ⱦ٬8����(t�K�&��v̱�Sꡳ%f�*Q�N���y�' )F<��},�d���/��oAo�0���|��K��x���{"���{OӇ+ɷwwo��+�8�XG���n�M����������w3��$���/7yn��uT�,ƫq@<ogp��\��Y�r �>=��t�F��;�ٙ@�)M�u�ky�Yh�9WZ���ĝ_s��ͱ��mU�5���l�Ǧ����E��ZԬ���6n�y�f���+W�3�ܸK0�fE�Kxmn+����>�MD�ʂB�;bt�ށ�@qe��N�\���AE�h�=�ɫ&n�D��pH0�[��H�ٜӲ�Ǜ��lh�[��w}r����,���+0ʾ��Y�p��*Kf}*�J�9�����f�ޮ�[�-5p\��.��~�+�P^���>~��Ww¦I�!n����7:E���p��' {��l��+ Vv��
}Y�1v�AfA�������6�A�i�K/�˩��R��EF���/r���
j�-��e���ΡRz���VwF�[2L��Z���Y	봳��X�M
۳F7ujQ�g83�����h��)�{ȩ����Q�7�ov�gi:厤�f��bQ��s3��/��m�uiN4!��|n����Hcd�P�{C�1����Y�[�&���[Yu��k�Y��s#yoz���#[�d�F��2�J��Ö�]�,���l�������e�7Fj��tR&��ܶM� .��J��̀��)�d�N(�7���Ã����r���i���\�`�o{���έ��N��ɔ13�)�$Py�t���i�֭�Qt�����=�?[3302h()h����J0�
b�b������S%�2r
)J���
���$���̧%"F"��$)���2Ci��(

*!ʄ�


JZ����,�(rh� 2)��)
�J*�'*h��h���i
�F �"h�j����ʀ(ȧ	������ʁ����3)c0+&������F��f*"���)&

X���2h�������k#	� �(��ƨ)���
f��¨)��j�*�J�*���"ij�)��(
�����C/�T�o�������d�a�K���*���3_E��� U�˛FM�׽NS�pɛ��7��Y�ޛv��"�:HV����_P �F��]i:��p�G�q5�A�yf-9?^��0�FK�rް�1z���:��<�>��v�.a�^���өr��׼�k˹�7��Bl�?/k:.Tw�7~��1��D��r ˹u����:���c��Z��Jz��oI��ˑ�>᪀�!��5�k1֧n���:�a�5gX�G�j?C����%S�$i���ǋ^n���DF�1�9ζ5�n]K�ϵ�u>˚��|ϵ����\�e�s@d=����}����'Pwδ�C�ոK�K�/=�Sְ�&�B�z�G���ΰ����5�J������	u�0}B#�"��������~�OG�~�j:��N�s݇P����k|��F����>��I�d{}y�hz��O^�M]bO����9�n_cq�R���GR�^y?'��Nz:'&a�Ro�w�R�Σ}��:��z�ۨ|�:ǿ1w?C�ԝ?��o��%<��}��:�ơ+��okE#Pjz��]��NN���0:��d�G�f�;��D]T1�\[��sq}��w�� !s�� �%�$�0�O���ѣe���.GOX<��K�j���&��y/�ތ�����z�~��!)��>����j2���n�9d;��=Z1A���{�x��(G�8��G��h���7��<9��Q�5����%S�fj�O �%�;:�p��캃���d�.k ���9?K�w���������yk�'Q���Ư���omR�#s��8C��(@|s�7=K�.�a���i�N�B��Ǹ�:�p�x>�nA�����j�A���X}'����w���Pg�?A���w�#$�2=���h��
�36��8��������߽lz���.��4C�g����|�p����'���.I���>G_�w:�{Na�|�Z��3��x���jz����%>���ܛ�ѩ�ͨ�������m��_���@G ��؆�ŧ'����22_}���u����U˟�湠�B_��<���K��}�\���wj}�<;�F�K�j��X���e����~��]�H穟c����㛨Y4a���8wWd��L�)��~���kg���Ӿt.{]�ƹ4�s�f6[ܒ�v�$��U;�R��j�T�8������N�5} wv�t��U?��+`�*Z��ɫ͖ӥܤ��E�޾X��8���F�l,�=�(��G�>�Y����xEBWoXr]�.^�ON���C�C�w��u	f!ֽ��:���}Q��}�7<���r<��#�J��c]I���}�����K��p�{�}���z�>�~e�>I���5�rN��c��6kK��#�ozC�����������my t��&G!�琔C}�:�C�b#�l�����˘��=U�<��uw�9=I��%���<� �~���\�'PFI�|�}{.�9����������Þ����9���.@n3�u��ӓ�=��~�"�~���GՏ=����o��6��z�7O�P�}�0L�C嫧�h;���J~�3���M�#P���'-B_�i��5��PF��w<�.���n�%���c�Ub��f���c��$�%�{:q�x���.I�7���>��S�O�ϴu���y����:�.�����Fs���ϴu����|�S��b���y�R��F��0:�������D�B>�7�ğT��wjf��%��׾���%=G$�}���y�Pw����䜃R�����C\�K�5���:�%�aϳ�z��d��ޓ��L�q��7�V��e׸u.�P����kW�}� }���W�:��샋=��e��&��L���j��j��㘆��=�A��l5���u�=���'#R?o[��2�����~`�F�E�&�;��#�ϴ��K��>ޢ(G�(}GǮ���Ǣ�{��Y�X��py���}�����r��F�}��˕/#=��u>y��y?Z����vo��=�~�$�w�������MOѨ<u��pP~���z��'0W
��&���l:��^��#�@dd|y����}�.���w���:s~��BZ��r|�'#q��Z���bP���o����J���sK�u�'Ӛ�k���q�u�]��ݙ��l��@h��O���5	Hue���%�P�`ts�O.�q�5��gq�Jy�k�������;���5'oX��C_G�;?a�#'�s��˨FN?��ߟ��ѿj��wnOR�t�S�6R�^i��q�z6��%2=�%�����;G���2�vr�L� �����3i�әj�J�@;\��.p�c��J]�qԗ}�5Ж��guJ���O/���]m�aSKl�>���HU��f�Խ�ԉD{�󨎣%��Xg��OR�}���}�jw.T���ɹ2����7�Q�=���w�d�������%<��'��Oѩ{z�U'�d>A�}�u��Q:9�{W� ��c�"$G����{��2O3{�j9y.�;�>��W؆w��Pu��Y�y�'��|�!���GD���$��7�f�|�WF����}�F����d�o߳�ޙ˙�ܕ��y��}P}�����(}���+RjF����Z(5�����_b��[���r@dg��/ө��.���hz��*���?i:��5���y��������j^�O~}�ןu�_g�~�ϳ��~5�~�����e�a�n�(|������ט&]�X{.����;?`�~�3g?u�c!*��_kp���,Û���}�I��~����J��p����p�����c�����!�ןp�zy��g�rԜ�S�b��d5�r:5��c'�:�5�K��.ΰ�]��!ON���������4����o���	NK�A�7���5'�eO���w#���{��w��sdTK3x:	?������誒"4A�j��y�A�{���5'ReI�d>ߵ�	s�5�֍���#'��7&���u'gX�7C��_9���!�g������.O�{�_���F�|�g6��*oe$A8��# }�����}���c>��<��wR?O�Wa�i<��pL�^kI�jy����}�Q�5>�:��U-Q�{�.bw���.C��K����]{w���^V���yF8��DP�� _)�����5��k0亩�O�>��FG���v��G������7���wR?~�5w.�\�?��K�����t� ��.f��W���C�u՞Y�u)���@��M�~�+�R�2��-Oq�5~����S��5�m5��j�a���˒~�\����`d5�>��/P������:�K�1#�|h�ŕ��ν���ƭMN�Yhp;�|.(D-;δ<��M�ZS1������h*5fv{ك+_��V�	����t��˃%ֻ�ƏpI����<jPv=:g��n��2ʣПM�S��ɸ�fĨ��[�H�ڛ{��t`�;�Ν�KF�"��P'&�PV, �͡r��&_ڔS�+]�����	��:
R�2:�U�� ݾ혬��@������0�\�WN��Drv��'h.j0���t6(i��g�W^�}��ӽi�n�DwX@Q�G�uL��Xxz�8p��TB�ꔇswaw5�(�����)�W�]97qD��2�:]�l׆'��Wn�2�`Ї�l.�7�U �*�7x0EBr���আYqf��C%X?>4vl;���ә|w\ı�q�Y˫��?vS����0n�����ޜ�ޠ������CR��*�UF�	��~�_�*1�p\�1�y�}�}|kq ({�v�����k\W3�ꘞȝ&!�����4a�-+�>��0�&�Ơ�-M?T��s
kd!���}q�ֳ��S)����d�+�ޑG�*N(W��rP��WB�O�ڸ]��"�V�z-�zP�@F���ᚤ�q�|���V1ϒqk�Kѝ���#A}aU�����k��l�W����w<�9��,�Ji\��W�s����]C�F�����ǩ�n��H���9����^6Nv�S0\�]���hA���孭r��I��j+qfަ-�]�+J���3-�N
��4j�JV��1Ӫ˕݋�ek�7���f��O3�*�j�al8*�̗�sP�'u�7������*�ҧ*�{��K��1=�۳�85gN��J�eOn�}Uo�}��N�3
%�cqV��J�LH�I���k8�O���}�[�t���r1��B*$�H�#��-v��s��Ӛ~cjW\6�φΉE@ ���G]�ʩ�2��{H 	�<��.�c���*���Pc��i�r4�����~r2��;ԶJT��ո�V�dk��Qs���k��z'�@�WδH��K�![�{�\%�Id:Y�!�ٽ%�냦�S����5���|$* �։���pB�A�5\�>�'xu�*6�VnR0�0��7ZëyfD�*8��4���\s.�7����Lff�T�JF|�禡��T94ۮ�Z"��`�U�ܣV.�}�Yy�:��H����&��_�2�}��x-������#��S&��n��h��-U�=3feE������/�������{��
�����������F�����PS*��^�W~L��������@�B*�aTб>�SƝV18f�镕[�`ݭ�q��ٝ~�n�f��i��wDI��z����CA�ꙵ5VgS�uѡ"��3��^�c�T@��T�
�M7�c�qa��M��3�i�q:�ԕ����
$7�tŝԴV��F�4:�]�n�����Vd���M����=,I�\��IJ�y�֠dH���T?l�d5��{M�x�vvheWq� ]X�v�\���z�s�jhR���zF��j�sU���_Ř%#̞�.t��=2�M�n�� w�-�0��0�>����E����NI�G	���a����{�\�XD�7�hOh29٧��T��#�� *��x���|�YL��p�=U�xgגx��K����˩��.�c}�J����U��1���P"Ytz��t�����͐;UyxyG:��;�|�c����.g���K�9��(�,}�=�̂�g^�ShU�X���Ċ��aNh͔'�#@R�c�3��z��O>������,D���:�C���Cu[�a����
c��I۸y��G)3 % R=�L���%kX�`njm�b�KS�N�n_5��e9���uR�� "4QJ�jq[({0�զ�4fz^�\&ФǺ6~?L��r����mԌU4"\)�%
��=6��ҫ��+(�LSǝM��VV��soqq�#=yl˼�D%�b��c�s,�9dB��6��$��|��Os�j����d9,���c71�
�[8�gJˇ{uW1"ohۡ
�L��*�8T���*s�,��tW&�r�`����Z{�t�7��	�m�)�5� `��)1m�L��p
��­�@|{�*���Ϝ�pb˜D����W�b�h�o�8%L��>��)��W�"mjc*��pA�8L4�����J��O
�	'e����ת���w�H�zj|�:�NnK]mz��Ȼڦ�f�%���4�e�����\"������m
]�2ߛ9�n-�3��<���`kO�=��t/�GXj�_�d?Z򐺢�=��i�����?l�����%R��IU�Z�3J!�Ps�p�Њ����&P��w��������٫�0:�s�7��bC���W���;;�N��-�S��=��AŃf6	|dz�6�+�9ߺ�t�.��Ầg�DA����k�>γp�W�kk��c0ƇH��*tjK��n���V;�eq�g�[8-��G������񁊝�V�؍ۚi����k(��8�Z�h�1��(�b;�� �C)�(�{`d�}�U���bk��.3 s�{[t��Z�oeq��C����0���2��1pD�L����sc�^�>�<'����ؠ�u2t�j��(�Ujլ��i��@Ll���*%}��ٝ��G�����..i\�^��?R;�V®�!>���n�\N���L1M�NۅF���\5!r�z0�&�����p<�Pe���2d��k����;�ҥcj]�r�f-@IE��0L6��J��V8�c.# �"����J��L��1���e-$$M�{�f�*�p�k�q�uE������k��n9��HvD����%Z�)#��s*��&��E��a:s��>b�f���h奷fQ�7�\s\�P�܌�uh�g���dc�6���[�6�s a� d��@0�����o�hy-�f �+|�Ƌn`��=7ܳ#o�W��{+����ac�m��D
�5P<�h])�2�:�t|����rՖbd�~rC�iŝ��;+����nU�>�ޗ�:��Ӿi����t~�G�3�+8K���\��GZ�3yk�=W��j*K'��%`r�ב��&!:c���~FO��F[��=fٯW�<ɺl�t�7�z8C�.�C����L�0�FE�.,���*��Ǝ͇�V�@]�$m�w)���6G���B�7���;��wzs�΀toጁP�P��]��s G=�^ ��nc��Uv�V��w��_ȀA[�t�����W���_�}�o�C������{խ�5��#eOu{*�۵أ��cwB�t�ݕ4��7&$f��Z��5�z�i�A|L]��&�u��ȓW�%E�o��Oe>J=���:lA�f�s���XҢ����:֠���+̏����h��ꪯ'�}�ُ�2`��9jY�P��jx�t�Bc��Wd!���}i:�q��+�MQ�&Q�|$�q� ��~1�9�w�U�v��x+�x&T+��P�:�R�N:k��\��9�KzUQ��'_w���ֺ�����Lp`�@z�aJUF��TW	����� CG��y���?
����F�Om����hFa&�qpg�������\;����{%�p5�[T��� �|��f.Z�7*���ғV
�v u�z�5,2V���9�w�@b�C�����ȡP��ӟs��ӣ�3�5p��T�-X�܌�78�u݁��h�.��T<�����f����_)A��]�w��=-T�詛�K��p�zG��(F��q����E@\ GT�O(|�D��R���v�)1J����ܨ5��F?���o�:nR����4���0�Q5��v.X��U�fP�)����bPG����a|ф�� sN⑑!
�0�PH�%:�0�a��;�j�W� sG<�ȇ�����׻�V�=�jw�!Cd��y�ŧVoi�h��V��iG��J���:�����A4�v�Fܭ��鱌��a�'6Q���{G�;��_0*�r�^'S �B=B��Ko�*��Q�U���o��.�Μ����:��%�1�S"O�~�1}���*�&��\��CXB���]��o<��WC���z"�.�zOb���MO<���$�`���=�l���۠9�u�WO�n�v]�YH���l,5�Ŭ`�|u����\�.Ûn�9;�1q�~D�r�N�6���
2��_{�ɋ�wX�(B*�:
��0�ਥ8�hB��\F�>�se�͌];ԫ����H���%qZZ̩��������1�=�sr���K��VF�������с�g�/z7(�h½ٓ�{���ed��?:V�FNz���^v���{����s ��6UT0.��r��f�>KV
0p|~̜ז>yH�ګr�q�S��S�l�`�h�luʶ��	��\��U_!�3��!�Ud�N��y�v�M�w�7Z�8�����L�L_Ԥ1���P*"Ytn���~E �w�� �|��7���e�q���G�BA�Ep��P�(�mzr�SB�5�\C��DNNWP*pj£Kn玣.l�����)����D7�O�3�/���M8��ߛ�r5�K�W��坶�2���|Yޒ�ى��et��خZ@�m!�����PX/����=�xJ�ވ3�{_��)!k[�v����ftV�=��il��F�ܙv�N �C�!�֎7z9��J[�[@Ws�� eb:�x"W�D+#VtJ�� ,jy�;F\m�Mgm��Oh�:@��P٨B9q�yH�6ou�j��C[֟�0Ď�K\Y���G2�s��-c*�F*
���l"�Y}Qp:U�y��TC.��JC�`�e��h�諒R��͆�+�����Q�2AX��Y�E�N=A�zl�[���gPZ]�[�K��15�ME��b����5R��Z��7۬@��;7�y�1��)>'*�.�u�s�;B�#�%c:�9l����΢���0�����g�[կ9O�3�>Q���Ss�s��Ȩub�n���q3���j���7!]�Ƿ�@��SO����1���R���2H#G��i9"�K�69����$���(6���y���t/-*ʺF�R˨�-���ƶ���&d,#a���cƧ7�/��ż�m빰	/���&�U���n��⮮�K =J&a�/=ݳ�Q��̧�$�B8�0�;7�@�9�--� mv��p�a�J�%:�g&�	�Bc�F�Q�F��븝%8����C6�E�`��\�6�Ԣ�F<�v�"�����m�dR<,^k����$Ek�Vy2�A-�WP��V�ܾ�y4?�{G}�+�z�d:�Z��pQ�턪�������`�{oث@8��Y����&k����u�h��,�ͫ	(0s�؝i�2# �G�;1�E3Y�]=Jdb��&,�Vm�rA��}�Xu:�[b[��Qr��I�N��+]�n�;�m�^cN`lS84�`̚��~�M����P��4wGB�F.�P��D�k��`.�;sd�)(��	Y����a�ﷻicu|2�;���]]Y*E�*[ӷ��������d�w�q(֓4"���ѽL��owU�=��w	�)�fWWi-�tw����Ŏ��u�{{��"�ٞH=����Ea��P�
�Q������;�]������4&�N��a���[��!�Mu�R�}��˳�B�M�"c$����T,&��F���Y5w�Jz0Z�\[{��������V�*#K!���jF��'r���`�B�Wemu.L�ΆG����-��O�/�NՊ�yC�f&&,��*)�7��Y����qm-�-�.�'q��²U��m=�h�5�%۶�&�Ƞ��mcP:�}�����n�y�ԫyg���0*�,ky�B�1�U���1�QVE�f�ȍws�������'���={2�î���V�r�6�I�S�v� ����N, *B��(-c��eU�8�DE��D��DdaD�AA�DQYd�fa�UMQP4�EaSMQINNMAIMffa�0DR�PLQ1QVYTD���QQE�E-�TTE�ST4L�QDMUID�E�RY�8�QEIAM&f1ME1U,ES1TQ94SM$�$AET�5IQ%UQ0STLdd�0�@�UU2�DUFYTd�PQSQEUAYIURDMMPC4EQEMD�EQ0PDP�_B���..�ށ�L���v�F7G2M��5�o�ڄ����k#l��W���I�4Э�Y���6/0�a�j;/��������3Cr��U��ک�]E���c'�F���w�g;D�, ��Q����,��lG�t�r���(8�ٌd3�ƃg�*��mJ6>�ʊ����0��/�拮�%aom��ϐ�ͨ�Nㅩ�|wS�5��1�1�>�k�� pC��1�W�{
Pw���_���ޫʌoF��{$��	�lm܍��Ո�`��Ōsh�5�Y9ZԳ�4J��;��v��aϐ��]ms1��.q���ջw�g<1��c�^m�I���^U���p�i���H���F�rN�;��|h�q���o,I�k�9T�t��l2s^G9/��f�v]K5�=�H�}��~��~� ���kx�-jFWr����r��)��}��U{�H��5]���~>1�g�{ �J�,��3��0&`��v+��x���<�]Wy1S����1�6=�P��0.�1�{�,��{u��lݗa��X_��b vW�:���1]��f��{j��Έ8a�z�v5�fl�ԆΧ.������71�]�}�x�FtIѡSo���5"�W��<M�܄}�i�-�,��oo$��嬭�ɍ!ã�����)�sd=ObBJ�\��=���f}Ү��=@%W��h�YY���ˬNK������\w�/��mP�5��UUUU/�����1��V����D�b+��^�N�����tϱdW����m��_^`^�͢�p�z#�?x����>C�^��A�E�<hw�|g��rH��WE�����#���׼j�,b���i�uOɊiHG��A�DW ou�X*7q����"WiB��{>�\/�jkn�Ѐ*i��EG���W+���5��ԅz��t��pU�C!%V��a�t�������W:��帄��a�FU��p��~��}�+�m�7�WEL�/�r~��^=������HvK���i�%_Ф�Rp�Ӂ�na횣��»^\�>����QFQL�Z[q ��yc��� F�u"�բ�J��)ێ���I���"�0��g��@�c����u��Kvٌ&��)���މ����|h�n;����x��٧���D
�5P3ژ�|��(p�Qh��ӽh!+�"�}W�t�[&�Y1��I��̺��U4��t�	A.8�rj��I�����wfQ��z�S8��mHr�^]nRm�Vk�yK/� ��e�n�ו����,����/������@[����=_˗�X��zTVǶ�YΙ�aL+y��}��sKEd���ڜ��]W՝�3*wV`m�N����v�����ﾏ��@�.6�b[#�����uļX�W��L},©�+�@v��jZ}f��),�X}B�c�Y�
zaf��3�����w��K���\`O�T2U�?>>��WM������m�[�ɺ�C�Qt7L֓� �Ko]����{� �U��y�b]䣮��,3��;���6�
��	P���ۂ#�&7ǫ#��Y����+���T��S�T���5�v���h���L/�j
�E?�O���E�/�{ep<��{6�g�%��[c N=|+�k�:�vM��b�N��o��� �at�]��M�|�-hJż=ܮ�U�cu�q��z�[R��)��Sǃ�|sƒk��؍���FR��Ê$L:�W�x;ι�����u��7>��=Yr:� 0�Hk��Y�y���V��ȾM���2�8�
�? ��p�������[|7&�}���
����	=�=΢$ADxN0Q�L��>�y?p�����9�z���oϓ���4Wu5��$��2�kC7+UW�S��$1;0�S΍��n��k�<�̺I�������E➙�X�`�=�ݘ�wp{��0�0�
�[ݖ��x����έ/re�	J�"K��_>�9��,S���J�÷�������b��%�\�ܫ=�t�m$A hE��Vҩ�S��./��H��*7F�j����+w�T��_�(}�ʡ�w�ܩf�9Q�A� g�{@�W<� �}Φ���m\��RW�8���']��cwM��S�'0Y@@k~� h�)P��Pk�[Y��7��?DÆ��Vй~�OC/�ٕ��4a5�n��V�*�Ȑ�Dq�#����F�:�B�y}� �ї��1?p���P�9T95ۮ�Z!��߁�w=j�P��\����v���8�l����ޟ�<��i���}\����R�4o��� :�6LV�N�����	���o���X�F�h�2>U��ק�Ȇ�g�Ns��]���U5Ѭd��fd8�Z�;��'_ܮ�o �4PP�d���5�`���<(��~�ܵ~��$��#�x�Uvy�|��4�-�@�qZZ̩���I�1}��릫к0�T�/�T�F�� y�P�������SܬR��ٗ��^�	5a9���l�����wu�WMt{�0e%WSR
�׼z�;���%�.�FZ�����Z4񫊹�r�q�G�VP�(Jy'�
q��h�f���*Ņ�=,�����������q\�j}�M'�b������w׷ ��!�$V�6�:����5ɞ)J��V(�����W���T�0���/z����u������>�USc��Ok�[Y\-��ɋ�G	��=�7����Ν�){�-�A�X�X]�ƣ��"s�d(U_!�3���d�y�]����9��]��	�M��^#��0[�%���^���GxJ���Pq�W�B�Fnf<��F�V��R^���R��`9�s�r���W��_)ȵ4!F�c��ڠ���Qʁ9���gjW�
����7pu�I��Z�}iW����2�v2�w��A���ऐ����	AhŲ��84����������J��v�3��VӋҥ���uIp�h`;�-�5���N��;|�US�cQ��c2�����  �@�`�Y�+�e0ou9�k/��@����V|&��"�"���ϋ��[u#;�ub'L#q�SW�˩�Ȯ�ԗF!���l� �H���/A|hf�
��[G>s1���(��B���ZQ��+J��ގ�b$�I���r�PC��aL�t�\��I����tQw)���{\:�����HS�������u�K(]����sC���Lu5ti���D�yOq�S3�jUb��w��R<:�h�Zb�P��}�/:5S/q���B��+hj���;�!3#+�J�s��^x�</<#��S��J�5��������O�=����A��*���:�u�b�ݏ��r_GT٦�]@�\����!r#�^c��Ō�����%_ �+��L�', �)��F���u�#��U��,���=�}�:���c���ٽ]�dB��*,Ք/�Ո�Z�3V�(9ٿ��Q�.�EC�$��<Ã:�~��2fǫ��EW�zޛ�#al��� ;:��!���LW?�x=�"�����zꜬ��W��KѾ`�$��ʛ�¤�)�a���Os\t<;�{3�*��i�<@�^��kG��[�|�fb�$��X�~敳���������/9�AW�7N��z&#r�$���H���b��@t��n���8x/+!�]�{���~ױ/5���ָUy� 8�s̱Y�]�1��锐�i��m��Sh�Ъ*>�C-��8�Z�{5�X����[��&�r�����epL��1��k���_d�LbO�ِ�P�1N��n�x4s�r~��:�9����:�{҆�����8J��G�Όڕn���9BMُ<Q����{5eU����G��W�k�ӽ=��<`��9�jb���S۽Vz�9VD�\�3�G\�����,�r9H�����oT�Z�6u��qw"��Q�ȦwH�bDxC�A^�r�p[�&P�}��;�8�L^�;��l	�k�Q>�4\[RYM#h�7>�͝ F�[vF"64��Q���IHQ���z�E�
�=���s�ꁩ�_���u��:vـ/J�u%g���Ş|c�����"i]z�=��w`�U7w =D
� �ژ\k���ţ�J�6��+��F��q���U�<���&1���a�;��SN���	X� ��C�TV����4"�1�n��n���X�9u�b9��uļX�W��L}E]�ZQ>��:��~�T���f��ZTzz��B��B?f��3���xx0Be���2,8��U�sq�G�\%Q|�6�]_�⢞�T��;��,gݳb���.t�c6�n�s�ִ`>�Y��a�W�vswPz���X��(��a8^������>1p��s/�n�Z�f��5;�n_�w^��ĉ��,_L^��:`d������\���\`���yX�P���<��ݽ:��sL��j֘�"P��@IQU�U
��V����xI�]��]�k�4�܎V���#������+3N��˝���p晸\fՕ(�^'�W=u����c��E8ة�4��.�-��^&����G�ջ&�:u�L���A��Z�Slw%YN�L73F��g]�l}�z���[+^K�,q�Y�Q~���������v\��bw���;��Tc=����������;�Dhg����y8ȸ6�"q2_</L�끵����ʹ��r�j��pѹ�s����ˑ�Q�hS��G4^�t�}�j��ӼB���ӟ��-�agÝ����1t���yc�y!��>�U���L�^��$F��I�%�T��)� ����u\bQ���ޜ�rzr4�����s�O.;�Amꆬ�M��6�d���� �4B(w*֕O��?���� *�m�$QMC;7�HUm�n��=��װ�C�ne�P@�Qx	�a &�>��P��Fp�� gsP��ťz$8U������t��n�鉕?&`��� h�)P��(��j�pn1c���as�1�Q�!ɪA��FcF��y�O�OJpuЖ��POue)������lz�[�G�K�����L���P��n��ֆ���)ݰ|h��̆�ώv��s��P"��Gc�vJy���$�`���y���a��Fԁ���zD]36]�U�;�p�Q����K<*=���LUp�8�bՓ���BU�骂��,u�Gb����w�2��תi�ɚ[d%���J�b�t�q�����'��/���q�:���:�=���j+���������ݧ{p\���
��x����������[���12;��/��lj�(������|~����]�L��Nx����ht3�p)E�WO��%^#!�F���X�������PuѯC�)�N���eL
���4./�b��*F���[p�: ��0�ۄ�+M�[�8q�$�����
���Ƭz,\]G�ZA��,S�����2�|��jhD�{�����_s�V*<u�2N�<�Y`�)=~Ͻ�)^�Lk*]ا�g�Ւ���ӟ'��.��=��0n�vF��~����ޙd � Ȱ�<�(�>5T.7�s#!U|��L�읩tu�԰�Kѝ�}a�=���FtO�tvSK�U���*�C:�Q�K.�y7���.�MuUj���z���=>��
>7N"tW��pt�p_������\����j�p��7V��J�����:c0���Cނ�͔2|fF���cC?j����q�o�m�FRQ��Ӊ��5�Kyq���=��q�N���T|��'c1���N8��	�0*�[YK���s\��z���RC����V�e�V�{3���^е�
�\{O���`{cV�5$��hJ�%���*wF�0-;�4� ��-Z�P�]�a��­m�"��X˻�)+�ytJ+�H�n���� �pw��ۉ~��������}���@��K͞S��w\#��8�vͩ��D��/F$��p]��!�k1�7���an�n��KJ�P�Æ��nU��P���R3�\�J$��}�9t�ҵ�E�L�ΧOu��N5�_����(���;��<:�b圗��tuCZ=�Mt����/�C��tf�|Z|�],�������¸��c�Q��D�V�ѕ�naN�Z��Z�H<������8�خU59m�>��*#\\5D�
[KkkE�3,l\v�^��ow]�VU���[k\9���m��qfrьGT\����I��W?U���}���آ�/*q�����=W[��e����{$�l��&�9��H7i��MK[�.t�ޫ����}�q[�!Ȏz7h4�/?tڋ�#�N��^q�Xs��5](�΁Us~��m郓�hp%��ʤ;%�Uǋ���{�F��2Pw�J�$)�rήrP�������c�1���B/���|K��4��=�%�v�C]a\X�b�n���8����!I��
S���[�pc*4�^�c-U���$�S-˹����f��I.�Ͷ��S�ˡv\hH�(��ݗ�G:��rU�E�*m��}-�[���#�n���v�m�̉�N���2;��Ȑ�q�v�+Y���e�a�m:乓cw��gp=�)�-.ø�a�Ѽ<��gŻO��ɦӱiMWQخ���
NEV�"���u5�����N��`�`�[w�>�9;2�f��TV��@�L5����E*�rn^&�İsW�4�ZRG"�����	���u�P޽��xч��r�M��OxWQ)ղ.��Ӂ�;S��a��՗#��2�u�����*Q�R��M*ؠ���i�Oc��*�cX�8�d���6���u��<ib�v��i&�ZѶ{}u���:0q�];tδ���3�:��H�"e���kr�l#Bc{�˪E�LKL겴��!P�j��a��q�,v�Mr��7�'��P��4Э�A���wy���M4���cP�+Nh��G0�2K�ɒ��OD�:�L����h����q�!s�{U���-xҍe�[�kw��]`|���IV���]o**j��DU���<(��Ýw;����@K��&�F��&2h,��[ܕӴ6���LY��q�cn�;�]���rT�|ux6�Ws�����G}5��Ĳ�{F�[�-�$�6n�q�'*��(�����g���̣^�GT�Ѩ�m��oB��gc&�����]o���.4v��V�Mf��;9���`�x�)- ��p�k�^u���H�e�лBm�+|��ut0��jµHоEPW �#əi�`�ֵ�k@�øT��6��k6�/���]��P���5�FQ���9H�I���ɒe�=-Bwf�K*���	r��H�����dLP�͚�G�ņF_<6���4R���y�9|�^W�udEs��9dnP[��4�@,oW.��]͋�w'u�����Hj��G���S�bژ2g*meh|��`��-0d���N����V<Ǵ��+�h���mK���s�<>�c�nZ�s�ʏ�Yf���p�C(	t�r�*N�����[�ͱ�x'H��k�EmGƶ���yW�A
�c�]���x,0�k�j����d Tq��� �p��vc6�$I��^b�ُg|�1���̰*��0����y�{���5>ZF4Q*�.�����Dl!�ѝ��"�w�4��z0��˒���c�&��E�loZ��h^� ��"��k,7"Ց��<S��
�\��'���M�K�I;�#��]�O���B��3Y��J����{9���(�S::e.S\O88�n�T� T(P�
��(�(� ��"���I(
��"��3")������j*hj������b��� ����I�"�"�*Zj*��&���i"L�*������"���!�h���*�(�b��b���"�J*���%�$���#"�ʌ"����"J+3+3
�B��&J�i�������**� �*�b)�����J��&�%�ifi��
�*�(*��(��"������$�"���!����"��
���h(�I&�f�rrb�0h&l��,�(��!��f����	�*)h)(��*�*h(�&(�
j�������o��{H��6�����!1��\�VDxVe�Ĉ"���;fki_K�볖un�3�j���v���<�dD�}6���">�蹌�T�&�Kc�J�����<[�)����w4Յ6���%F^ʢ��H�CdC�T�>��Wa����>v�\K綧95s��W�W@�fxr;UNzr��毶\�ň��5���e��>����Y�6�Z�!=EXꀠ<�����1i�D��.z�L�vsz�X��C�[���h��c..�8�J-v�8;��	"97��+��5�z�3��ߑ�iX8�S�<���}�|���*�_r�1�_o>�o��rқ-8��{�o\�t�g�M]��n��Lg���߻r�V���{<�v�䵴���wf�ՈQ�py�d-C��&�|��EC�sJe�}�.��V�ۙ�<���EBR�:mpW}JZ}��l%�S|5��'LQV�G�X�3�N]m)K���&����5�c5���ֹ�I��aMָ�o�����G�\�=�U��Y��o�)��1��#�_(*B#���Y�\2oUѫ�S{E�'��0��Y�Z�BJ�xZH�B�����;B��n�6n-۷��� YF	)P7���t�E��B��dV���R,R����|x�¸�x8\�}_W�����QK������k������j}����^��z�-o����a�tf7ofG��n��U��k�Z�%����ǒo}�,7���ګc~Y�VO'�c�ī�l�h]j�']'캥�K���U�<� �ky@�]��^���^͟{v]{$1�]Q檇��0J���m@��u��>w�0��{�,l~�U3���^�6}ڮ��y��P�|�m!�gW�+g��L��:oo�Ok�����Ux���ZF��myNߗ#����b@ŷj-��9�w0m}'��G%����'�P���떞�2f6�bm��37��Y������"��ht挎��+W*ikyz�CnȬ?&6�v�\��n=k�ʶ�l���)���¾*����ܮ�.�],�s�U���&w�k}�/:"��黁�]B����(���	�f�m����4k���6�Ƃ�ݜ�>��I�iK���<f̾�[��E/r!�!�{�~ޚ�>�=��V�2���`�jjS#�x&��U��)���K�� [�i2(ø�L�Dm*����T}֩KK!�m=Zj�^19^.�]&��{���U��_}]����e)��>���B���'�*�Q�M'%�B������wx�[GB�񼗶�}��-��*�&����|�M�3.r!L�K�Z�-VeL��#�zzf�O]!V��V�B{�U}˜�o��vťIj��.ݝ����6��s}:��mL�6�ϳ~��T��o�=O^(K�s_w�Q���e�c
�w��*g�>�rWf\�����괻!�E^n�@�M9�U�y��\\C��n�CS������tb�u���K���T��k^
�ulOv-�z�k\oJ��ᚷL��s�f���"�Fb�u�y��T/%��29��O���8�V>���q�+�'��K��{���������Ww�����i7�nr���Վ;=�*yũx�"�놳�P%
n��i����s�Õ��oeA�YG2%C��8TLo>p�Y�C4ߙڿ'Wpf����M�NA���䙔�����7tݒ�yҠ�݄�>W1<�9�;:t�M������|pQ)%.�	�s�o��S'Tf][뮁�=BTξ�s���TK;�攲k,��
m�_i5�h>T��Ks*^�y��k�U�}_|��y���9�,kU�花�\@:�}��u��1Ew�d�3	����&P�.��/�ڜ�mas�v���<��%�u@X.Ԇ 7ܧX�J��w�(k/=������«�\!TVW�a���߄�dT���Lp�y9�])J�P�sd5V�M�|����4ͩW���w��EW�ug�����kr����ۉ�uC�r��)c�[/��������$5�g�R�>S�\X�JR��,԰<��\�&�d�Y�,ds�!��z�թD?GB�О��˷�^j�+�?J��q�[*���	^���0]�	��*�N��Ц\�q�mO�k�]�_Ӽq>�X���\�<�M�n�8�O���h7�������������dq��=7G���5��>�����*Zy;���k�X��|��w޸��B��m��9ç���D���B�k��'nLv8v�賎P�.WKt�u��bgg]����R��-�e���l���V�T�4��G'!O�C�̦���c�w�tM�mC]Xb�;yl)xl֎`#�X"NyI�1��(ޙ-K����wܺw����WՋ4�/E�~����{�4�eoi���[k\9�yNv۝��k..���q�tWrٗ���,�	%�$��Z���\�W��yp��v�\�r����+_Y�8����_��4�{iM�T��Tb��ה5O1�gfM��	�::�ܴ����"�{|�����9U~sj��nJ�߫V��)���q�F4��-�K9=�i��i�SՇ��wQW?����0e���C�l�P�r=��+��*�k���o�9��k'�+��+���p�m�	�U�S
���SЕF)J5���e�O�Z{eg+�F�2W���BV��g ��m}'�}%�rf;9�p�/�����-�l	�ڢyT��{d^Bjs�Zps����H�sFw�q
�GƜ^���^������{���>]T����4���}:���gz��&4���K;)ۋz$�ةй���<��_��/x�Ǘ�O�������|lR�Wo���pX宻��k%7��1>���p�ʊ����9D-������Y#}�{H�%z,9]����\1:� ��f\|i�C�U�kB[(Y�߾��艜��'"�^z <Oq=�m�s.T)����t��9�ԭx�;63�W �Ԛ)-�S[��$Ҷ_p!P�ȧ4��#�]B8]ڮ�h^T;���;����&�Lgqu	s�M�w���ħLTAV˪�Z��^a��Nz\�u�Nԕ�5���X�5��J�,�&�q��)��T�������������|aaV6�n>�;ث�cZaOն�Ù��#M#��ى��9�=�c��X[����g:^�t�:��4�]q=v&�5/�V%��֣���:��we[�3(����鷥`�[�Ť�wp�n��P:+�X/�I�r���eC�×�,�U��2����FA �-VgC���g�y(��@���Z��������k'�*�b5��Ŗi������݂{�e��Z�ь�G��F���!�}n�v�!���	Q�����`���X�Ï�1�R#(ș\z�=6�	S�0%�9Rj��lv��N�77�.�"�u�mJ}\�q�̟ud���>�K<ۈ��2B��%&ʥ;M�Ǝ�����oR����L��i�i��ڼuЯz��Gt=! e���e{ﾈ��5�9z�Lov�OǺ`U%�DJ�U�Z��&-BM5�c��u��2�ay/1�c�<����p6��挍/N��\�ݾ�xuC ��vy�0�Q��N!�{P�{e[q�V�@8m:
�vR2xK��#"Ǣly��
{g
V�-k�\fվ���7_8�*rV���o�ĠW�����+��1i�=5
Wu���!=�_[c)�)�NK_5_P��WP�m�m����L�w�[1}�RM+�g5�pWɼ�e�;9D�!�DffEнX���rЍ��n%ne�Nb�J�\�|�x��*D.xy>�[#)�[�Α͹���������־����zbu��wÝN��XE��j
�����(�a\O����_�����G�e��bu���$�t���<��y��8�է�n�o>���Ź3}/3%�4g����{z�K���x�s)�5��`$j�8��t�m�~��.:�`���*kH=@�z�T�D�L8i��ww�I��z9�PY}ܪG�ɵd$�t����x֝�G���ԓ���B�Cr8���q�i5�z���r�w�׫X��Y�興���32�4��U�d�YV���{��4��qu٧�Ɂo�B���c�
��|�έO`���++U�t��|�;}.v��W��t̱5<j��Y��@����Q78[��v>w�S�/�/by�t+�'�:���sa��K�Y��`�
�ol�ʕ�t�����?'�%q��gk��Rؽ7���S�:m���XSk����ګ��+G���ѽ�K>�=�V{��+	KM>���mNuCk���8>��~��=�2�r�̹����z\���_F���Ἴp������ej����3G��MБ�J�(]%	OO1�NJu��j�,4�<�p��c���^�M��*l�mss��u�s�n�7���Jʍ�攮�-�rq�O��n-�{d
��S{��쥻��,�9������O<7�3=!�r��s){���Ko�	қ(�JpKH&�������%�7���g{�e:�Q�*=�5�$��@\�Z��;��t�ϵ��wvP��c"�ЙV��r\�QC�����J[�f��t:%K�YV�l�˸�]W����@p����j�'j��������Rg�����G��j�%{*�D�m=ِ:�\{WH}o�7"�W�|�H�54m��B�7*6�ce��<A_��Jt櫒�t�C�˗LXg$K}�-���y��ҩ.���w��
�������>��7)���kΡjyOa���,�,W�Gk�i*��c�5	��@Sz�>j��*�_��sױL
��swi��.�fT�{q�2�w:��k�4��;�o�|D�S;+�V��j�tO��ʉX2�9�ej����q�����w]D�����j���~K<r��̣���R�[�K�G�~��~,�޸���c�����ƫ�"�{���wju�o���;rW�RN��
�'-P�_)�U��:ЎS����ґ��^S�.ă��/��Z����q����f����p1���˛��i���
r?�݊[�FN�zoٺ�z���/Q��R�Nr܏%tM�6b�*nV�W�n1ˮJ�J��FF&��CҲh���R�Ά��t��R�1nP���s��dt�T�R/{���<�ό9�.��]]�e0�ES5p��RV�d��Ԗ٬2z�_;�z�g�����ݹ���#>g;��d�5�M�J�kw���>-<ⳔWf,�q���E��5���)��`.D%�_+W&{9��n8xckeX�S���%!t�2�����܆�@��iT�NR��ہ1�k��M�����B�kw%�i�s)l���o�4�J'��amvrqz:`C�;�zU%�8��Z�n��[���le:�5
d��v����o�
:�LK�IY�f��8��١lri\2�;��
��E9�4�\��ق*Q��22��/�sw��5x侹���;�����Bo���7�+�劮�u<�p}�:ܻ-�_���$�sj�#5�J�B�bk��k5p�]d�7��6�w�Vn��q=/�]��ߚ��vy<�S]��l��}}ٳ����MHJ�3��\��������b��y�+W���N�m.U��ǵb�A*,�8U�y���+j&Jd�c��6.�A�O��=*|M�(�@r���&/p���b��9F� z�$���t˛�^ѕ̆���+�����n%d����s�HWmel���7��[[0�w�5����"�7�K�m8�'��Ve�t�R�܃�Ji��L��2%n�^���FhKz�o���P�6���s����Y��cp���(�K�F5�f�kaa�f-�R���k��h��_�c�	ِ����&Z�̇2jڛN���Rq�$�'{�$���J̢��r�r� �C{1$���b	�;kV���&�&���]��wˍ�0N^Tհ|�q1����D'W;c�K�W��dQ���y\�ʸ�F	�9+�*5���Ұ�K�Q�Z w ӹ�hSal�"^\"m�4ը�[�؏gƝ��{ې��Nk�p������n��6�n����2@�����cɘG�NMJ�W�U�l���6k�Tu첥omYF���[ï8HE
�@\�Q�h�Aջ�&iE��g$�ʰښy��[�[#��$����Uo9�Û3[�kr� ��@�yӣ�������!�DE��l��5�n�!�Hj�k� |�z��l���{{�.4k"�Do��Ǽ�:�e�9QZ頭�RT5��׹�{`{K[���-�A�7){��7*��{�W$�+D�2�����k���;�X�Ӻ�t\��1L=@�:�rC��{c;o)�ԫrr^��f�1�L�u���%F�S��'E��\��K*���-�إ�@TU�(��l��*T��iQ�0���fong��-]wp)* p'���F��>�Qq���ňX}�!������(ûz�fgWo�r�<T:�����oد!zޝ@��K�	
���,H�U����۝��|�N���
��1��	�W+y�]�*�^�r]p�j����,ԁ�o&���s�[5̩u��,��{F`�d�kK�F��|�m1D(���×��;�nRYDߤ��R�j��'�Vjᔱ�0����f�3��%�������>���X��B�o��YZhe�W�=��y�x[�m��r(��ӳ�KK�kw�-J�h����J���|�3�h-qS��뤕�i���h����	�8�)ˌSb��2�E�={��P�q=!)bhG�n��>�v�
∎p��i�U�ڊ츯m��VKjk�-��}qk�J�:��NY��� ���S1��'�L�WXoWtXl��WArw9n��@�E���RV3��Ea%�m���2�k΍�ty����'���S������wZ���X�F�l�t�XROi|e9Mdp��kL�[i������J�
3�M�&�\�Q��v�k��s�h_[��S��{] e��F�Qާ��qLrP������͛���\�;���M��?L�
mc�u5Yݮ�rN�(�>��C�>5Fbd4ME%A@SJ�IM4�E0D$AI!0�!��a�4��P�ED�d���P�SUACAT��%PRd15HUP�DVf14PD4�-��4ٙPPQE-11UQd&I��4)�%%%D�%M499E�AKYQTEE%S@�����CUP�RaeIA��-4�I��PSE-S3�EH14�d��PR���Q��MULP�TAHTAE!A�IE��T%%4�M,T�5DT$HUԳD1%D��dP�U�&>��Y�����l��fU�\��+הj'���ސ��
���97�����g�J�љZ���J��_��*�����}�`�O#s�"R��������{.v�{-����� f*�{�ڭZ\%`S��6�Kyou_L�����ٲ�۲��!��K��P�>!�t�>���b����J>��矨�z����ިƲyI�a��Fɝ�I�L��� 7D~kQGT���T�Ք�~�w���{ZR
��uAL�
Z��\����e�5�p[�)��mJ���&-BO�/�$���5�*���qG�5���thC����P���������+�r�� Z)�Age��i�AY�4�9Cyx��&��m�|7
���);�p�'"��Y��f�-q���N�M}��\sֻ#\f���eBt���.���!�O�Ar����*�g�������V�'�*�P��'%��Ȭ�������S|���0������b�J��i\3��@{�7p��ƉQGv�����fd!�k�64py:�-�@�2nH���=W�X�W�o��j N�����v���sw�o�*�:�;F�5��e�=j�4�J�je��'wP/m3uz��lki�[x��/0�봞�
hq�{y3����E���W�T���:=�;�� ����b}5+s.s�UDr�-���Z�̙��Y�$�G�t�6�>W���tk����^��gb���茘+r�tm�̃��dV-.#[bi7����[=p)�m\ٗ���uO33}ݶ�3J��:y�J��ZYNh3�&��59Z��a�01m@�B]7�5D�a�VS��{��&��_t���N�t��Bs��a���6�ݫ̙]ݰ��I��{X[������[ڡy��Ӟ~>y�^\T�Đ8����=i�7�]��#�9�<�b���|�y��)z�)��͝�b�qs��C�C8<�u�zu�Hq�A%��6�yC��ϧV���u5{�m�7�9�$�[�{j����M��pgM�sj��%5+F��e��kU�p��p��������n�Wͬ.x{�yNW�[�i쪑77F�C����g=&�?q���N�1��Fu��ІU�3��k0�`�榹�g�<P�Z�voy(w�6��([¥�yd�T��޺S�e�ñFD�嗼��0�GL��'K��Y����Օ3��t�d�&��=�ޫ���WE���:tpU�����%_{�R���8o.1��m=����ª ������]v;͇ۨ����w�S���m�c���brމ��逴���6��î!}�lPo�
�[��wZ8�r���o]�L�uwOtl[W���vp�����K�B6�%5>ʉ}E��I��`��w-f���������*93���|�J��B������E�5�I��ӣ�T ��d�S��Z�8I7l���;�N��Ц\���֨���3l����]/d����ԥ�}9�]B]SQ�0���;
�8�>��i�5ʏ�k���Iz����/.%vMF,��x�%SK9�Mƻ
n�}G��v�s��/�]����X��ꗱl�T�{tU��������輤����E�(�9��	9�y�.���w����}�$���0��Ur�?���Z�s$%�u��"DS� y�U�,���Dān!�g5�����X�V�C����$�Ҳ��ž90�3�sR�,��z�RW���"��g��zu*�TT�;P�C$���)Z�I�;.��vE�S6�ȳ%��v=<kC��ΛƸ���3۞��u� �7Χ)D�Gt��_��l���et�3D��D��b�r��Z��&������]�N�p��L�o�q�$(l���/�o�s��_��������$�l��ҹ�-=N�v�Ψz�˧bAϔ��j���lNʙ��v�R�TwP�}p1D�|���v�\K���{=;"��f'vM�OV����
ډ=��}�+�ㆭcO�Zz��]9���+	����G�D�wo>��� �8���S�����[�2VŚ���yYF��|���oWhV�i��ܤ��CJ����RXr�E�(�cm�Ϥ��W��3�t�k}�/:�P꒰�_r�B_o>��M��u����sG�y�I�v򿔴�ެ�=�Qm���T�S%W|�Dn�`�J�K��/�.'V�.����4�|;c~M�T9�4�\�D:��&ȦA���7�gv�f&�=n�N���J��x,�+=޹:,�3kMmJ͛h���Q^ܨu]���Wr�v��$/NL��
A�E'D�/\����1�ol,��L�#����2�J��0��%�`�Gu
�Ԭ7�G%9G%�}U��<���=�aw�[:+�]��gyd��t�|���\ea��e���Y�9����mU]��;�'Jܚ��j1d�k�|��M�Y�jX6O9�}`���#�=C����UM������G�X���b���l�cI5�U�N0ˤ���n���9���79Z�S�:E���b/,�� «����P�=.7w|�K��M��})CQd�~�3���v�>%��>ޘ�k*�T�P�Ғ���c3c>�Z�:e`��;�r��!�eD=�9ka�q�U��A(r1��*�b�T��DJC��Z��/�_�^����ޜ��N�$l8ٹ���$��v3t7ڹG���t3������|�Py��`��YR�Cw�rbw,�og�ݽ�(�=;Α�k�s���o�]�u�s)�V�Dԫ������~��#���|#�v�*�7��g���2_e*�ߺ�{W=�l�e� Òt��Q_G�I�,7h�V�����6$J�(��1����M��,�� ��ߚ�s��Kin��*Km��s6\�K��q8<"�cHkNn��G�;(+nTz����Gz�a�������.ꃭ`�/�oR��\�[ﾺ�u��qn:eO�yq�ˈ�j������Z�6;��|���7�u'� ��3��,������)O.9�]��6�����/Wܞ\��D[tK}�ƶ��v$5�l-�禾R��[��=�V��uJlb�۬�ʮV���[[�_��["4�J&Ʈ���JI���o�����d�V߮���/����OV��ѳ%�GH�P�0�[�p��ҹs���?�owX�鳼�L�r�v���S	��s_q�d-r^ܯ�e�ƘK�z�=����P֐��'	*5�1-���\Lk�����O�j��Νi�Pj�g�z]�Mx�$��ӆL�}�r�'��#_&��59Z��a��m�ʻe�u+�w����|���D���^v޼���]��|�Ú�L��s�f�sZ#�%�{���Y�}��a}BIt$��n�������̝f��?<�*�/uz4��څ�չ�u����^�%��[�.u�V��k7O�	�2�B��N[YN-s{�C�6`���,�>u�Yn\�[T6����j��)��W¹�uԑ<ݺ�^AIN�ާ��o�e�-5u��++�m�nC*)zy.�&̥Om���pG�1�������u�h�|:u�j_�|6�Q���:�K}]ŜB������o�������='7!n��!�]���m���������Tp���'��V{[{ыuG�j���S�<�֛n�
�7Fo<�S�]V�U��P��ja�m���77�i�ľ{p�:�maw\L�=b�a�d�sq {U�JD�[
�(���5o�q�{��М�\&�\R�;$��W�r$[��4L0�H�{��%��Jy|᭿��ڷ�!O1�	��;�Ku#�k��*��Cb�Q!�RVV�sJWt+}�%��
��fO#�n�=�ѿ'=��>r�T�֧�TJ�J/OW>�3_GT�_^�B�f8X`�m��uNj&`�O.=��-�����:�4XYf�-�),���BmsW�/����pħ^\O��#��e�D�Sz�b�묙*Lz�Dn9ʆH�N�'/&R�إ2B�g��#�t���\��g��e��p]M��R�ה�����H�j���tj.��o0���[�ʙ����md��rC��{�p��dX�Pd��w�|�3�3&�];]5ý�
؅��Mӝ�Z�Ջ��{'�7��<�ē�v9&���q0�TO�[6����f}4:銽�'�=dܜG������U59M�>
l=����X.��!�Փ��k��%f�7�Y����vz��v�����Iђ���s����N�2��{|��WҰe��ŝ�Ar&Yd�/wS��}�Q?�˞~��������̨>����+��&�ʚ��f��9t�v9C�x��P��p���-�Os���_s�|���q�8��\��Ts��q�z���?v>����9��O9��CwEM�w R�䕊J)`�YGrzT��1E���3�׵��]x����^H�'�I�I����"�"�g:G��N��]������Yx���.��m�pL���#�ޠ��k�������r���d���[����i'Ӆ��y@,X�f9��w�]x6�Q���	M���I8�Ɔ�6y���kr�'�S4'@��:PG��ѯ9��D�z�T�gD�T$��{��h�t\��O~tv�vl��8���f}�\̧�]����SSu"P��,N�fN��w<�.�nvGt˳���ur>��)�s�����u��|���;��iTI��Ή�.�J9���6�^�PR��:[˄��ȍq�Qm��uI\��/�I�1(�7�.�g��Qy�}-
ε.�篜��<չ	�WΩ�$���v��w#,�ׯ.1��5+�B��Ъi_̾�<b�M�1����A6D{�@��Ųr]���K�Mĭ���;��K��&�;��c4�����������}Z��!����&�SɬY1��%F*�^j����K�rh�ı*��%�Q��qP����W�m�OfTD�sX��i('g�]�h���2�Rq�V�p�|���nr�����t���P�U��Ģ�l��En�`��vfu�o�r���oK�Z㝽�:�����W��������'/6F�+�<���eb�oU����ֵ���}�P�C=���]���K��Rl�~ۙ�,�uk-}|OQ�ɷ�(ma��rv�d.�����L��N��x�5�:��rz�=�۩ť]eM��I�PD�Ȝ�4�AN�{���*����`coV�T�
�7b�oX�ay��f�Q�݆�Y�<lD�nd�� n�\�]����Kc��Ë�
^���5�v�є�ò�Ɣ�Gt�Չ��>�������v?��uK�ҳ�7�=KgF�D�c�u�Nv�v�iwc�Ov�K�oa��E����h�5�9�j�\t��]댺9\ý+�VgC��i�t�"��k�x��n�.�ux���R��
���;�5�ky���8{P�{m��p�\�;���k�bEn8�(�a���"O5B��JS�x���o�Rtݍ�Єӻ��%�F��hT�A�ۮ �����l-�禔���,}��{����t��[�ọD�5R��_w�O�#L�`,j�-��Ҫ!&�����P/kr��,�� ]�w/�S)�O���:�t
���D{n�y\ҙ{(�	��mB�=�����[�¸w�W	�Ӟ�F͕�j_d��v/�ZC�4�á(&_���RS�dA�U�Y2�u����`�6��1���4Z|1��H�t'� w��a�Z��vW>'�*}[�[JJ�]�-C�}�.�a[ŕ���Pn��z�֪ڔP�Z���3u�&.��
���	�Y�݃Wk�,Ĉ��*aU9�\q��-�O+�%�;��t5�kd�m���U>�7�{�[�Qısb�|^�U ���&��.��JTn���Yg0�/�as���25���|�����[�s��ޖn�[�����k)��wR����kFu���<��f�d��RB��!�G��7�H���oa�ľ=O���v����cmӤ��ܠO܍�N�$�+`@2�X�Yktɴ*�۹�WU����)'� ֙ǭq�8�gJL!�ށ�Ж�,�M�F6b��h�G��TCr��H��t�s���1&�����m�}����L��N�r�ǽ%>��v��+��-����ϵʛ�e�޽�d铠)pu7����.�][Q������/+5���k��ĩ5��_`<T�p���s�o��wg���F�It����ñ7*�A�7:K��{Ec U�!��ǣl:T#�(g,�d��C\�7	(ڊm�a�LwQ���ٮmo������y��-�n�����X �j�aƑ��uߝ�04�۽ڿ��8s�R�C|�e"�R�BKE`���Ѫ�N<�[l�p�OLw�
k��-�idm�&.��E���9S�CWI���*V�r���l����Աi�����j蒥�*���w<�؛��5��\|��Z����R��7��3-0L��1X��]����-��q�[G5V���5�d����S��.2�T��B�^B����0�����ٜ��=��t�ee��HDR�jWE�nb;�w[\�w��&v-�/f��th�ĦCՕ�g�Y���ZIq)^�a�vQ#.v���*�3;)��dCQ���#1�
ի��Q[l�B�`a��59�*Ū�x�2͆��{S����c�A��ib�*�E"��W��}sV��QU�\T)�E��.M��0ɺ��"�tk-D��!k��-K��H���5.�Fp(��{46p_e�7���[�Ab+6�7ә�A���{z��͚�W��ݸ!|������D.�	,�tf�'Wn�m�y���peL���Ҹ�G4/�C���+����U3dn��'ʷ:sѡ�2#��A���7���U]����,${T��n([.&���R�ʲ�ZH�a�b�7ӳAzir=9*̀d�M����a�*a���g�ml�\���}(r����HM�$�ˮ�V3�m�s�5B�C�tw�<u�t�Q!T�,ķz�����F�V2�X%ۜq�+DY*�N�u-�\x5<��wTt�lEK�ޢ�9�e�G5�����A�iM���E �Nt)'��N;���}��MD-�+JP]XPRQE1!BPPSFY1D1%%T�RPdd�!KSP��Ҕ���P�0R��HP҅#T՘�-M+T�4%D�HSEUI�4RP�B�E4�MU-ST4�%
D#CCBQM�A�HRUHSIU-JR�P�UKM,IE��CHU-QMRҔ�R��"D��E3!CEQEPU- P�R�LԴ SDB�4��CEMD45TR%,D�B�P�EIAT�
RR�����*����Y2���;ד.��G�biu@)T����C�h�0�J5�5n��*о��ëqRˮj�W�E�-�A����\Mu=�,)��k��LO6�]�q1�*%�g�_FS" �����=����=�#����]Zp�nkS��.%�Q:�u�T��b��};VOYKk'v��B���7�F/W���3��׳U�E�6��<ٳ��p�bO]'�=���뗜�R�'Φ�[9#Lh���E�=��j�|�_t�=�K<���̔��n�Q����r\�J�H���M�<�Î�����}3��$�<�9��򖺽��g����2��I���[��0�nQ��"3^��x��=4;����]�٨��g��1�/\s��K��d�\q1|�sp�}r���maw�r����:�Ȑ�5b�X�����P䔽�>�BeLp�z�z��t�}@�szQZ��X���C�Q%*���+:�<���[��V��j<�Q��^y[&M7�ՅK�k����<��d�mG�z76�'��]�';�X�w���/|�{���;�I�{��lj:F���v��]�j�cJ���!�=������<�����s���7�	�.�|�wp��9
��RZ�;vw�l�5	�x�HNz�5�@6�BR5H���}e�/����Hi�#_��ܺIf�C�Ay'�6s	㛞�Vk���C�SI�u��&4��F����#�Rt�q�.�탫�(ĳ��n��K"��8�\�)���.�ls�=ٺ-cntV\-t�)���>���#�52�;��q�O�Ӛ�2�\>�g����i����Ok�5�j%�M}��qT�T�rL;�7�+��8������0�[���wǳ�y:$�ƨ�$/z)�>�x�%R�ÞMƺ͝T"�+g�28�A������k��c����S��Y�6�w��N�:a�o����ˣ�y�׫=���o���S=�{11o��\7~�t_d�So+�X2�9�\�ڄ`�[���
�c=/q�C�s����[7�`fv|$�MLo��.Etw��|�k�\�V�>��k�R��?Q���ؑ�.�חpF�\���g�z��!y��qc�L[���x��O�kb& �-�=۝Q�!�C1)H�nm�I�3�-yh�I�9�ȭ���4K�:q��n�߻X��M�KI�	� [H�7��ŕ*�+ܡ���qL�4��S��-4�:�d>�C���Ja����1n:ok���~���O>�iJx�U�89KGp������e�R��ϔ 7�p;n'��T.�/��/�7)�|��[V{��-�G�{�m���uݼ�G�g�D��*9V)J���c��'�g4�L!5<[��'���{h���p��ς���ͬmV8j�c=HU�ڞ�2*[εkz�����jr���n�Ӄ�wӑ�"@���$ݯ#�1<���65�9X�ԻGK�Z�g��6���U{vJ�S�2�-[l���m��T}��?�S}7��-v�pj�OtW���U���ܑ��J+U�{�o+]�~9�BY.%kˀ�c�B��L>@x�&���E���Z��`%UR�s;5�>��׮jV��bs��R\�M�k-%��9�ex�:���r:�Ýf��t�m�9�����5�Ɓ����L����>r� �Zۮ���>Y�u����&��8O���� 겝K<�Ӎ]�LPǝtr��e���z��,���2<|�J瘯��N8�*��0a�:��
�C�61��'�V)�ĶF��I@N4q(I�U�ɽ	kq��N;�#xm#s,�C����ƻ
o\T5L�O�i�OfTJ�4�Zi����^P�`��!�{5���%v�����o>�j����1Nu;�-���|9�t�'ʌ}9uj����q��˝���QY�>1R�WS�#�n��٧\'��Rڬ)mc���P��<ł�|�\����d��N8�v*(M,+ޭ�������2�	9�X�xG�FgAQ��ũz�jMI\O�Y]m�kg}�y�oa�N�����yF���3�a�n\nX��P�`룗��iv�j��æ������λ�q����>�N9��[˃��p�V�5}	;M>r�qWػ
�x���b���]����,�Vs��SP����p�_���&��Vݍ �����Ţ�<��-����굓JSˎz�k��zmD'MԊL���Ǖ�v1{�
L�T�de[ϰ0:�l*�܅��,ɛo�T�\�S��]+2�����+���U5�wB�C�:5؞��F�3�򓏊&�:s�\Ԩ&R���eZ��n�y���h�������ES�ڵ�ה�uL]8�^S»kI����}y&�|��p���_)]�c��Ot`x�C&����Rr'CԷ��ɞ��M��z|���w���-	'�з��is���������h�\�[��y���d�!v���O���ςg��_]�g':T;{���H�w)i��<a¨�銅6済��[�"�n!Ok}��j
u
��N-4�z���I�I��mƻ
�c\TKV�5W�}�ͩwt�l���k� �yq�&�NuZ�����M�ڈjr�\\V�.���2�c��@��+�&��-t�?����n�c��y]S����l�5���Ro�$��y�U9�we}f:���:�k��{T`Cb:��k�ŮGW.F�����n�wf�`�tz�g5k��uN�qwX!�xp�ݕ���.��L�R��w��gS�ö�fQW?�Q���cj1�&������
h�Ů��s�>��pywا�"��q�FU1�h��F���7�jze�M�ncn(� �X�m���c]�u^����� ��Re�.���ң��v���(��-�U�˓��kt�K�pl�ЅS+ޢ�Od�۝kx�T�)ȫ���q���$G'�3�o�S�:m��wx�	���P��Hm0�\����2W_�1D����i�ľ{js���졝�Y1`�)��;�+@N���'��_+�r�kun�P��i�̾<s�)���iJ��:��.��s`�|�K>���),5
S��i����R���@���s|�*v�q�C*9Swp��-��BQ!�RVV�rc�p!�lp��M@�=���=�e[�J=��u���'�+��YV�y��]w����U��cp�M9I@y�d�)62�S��L�_t����ٽ�%(2:���ڗ6y�ڗ:�/���B߹sW����:����%�ULѶ�v����o=��&�Q�|$x#9�ry�V��5�0���c�����hY�Μ��F�3le(LmEC�|twFPYwҞNC�5��nl�W��ҝ$�E՝A���۴�E[2W��*ݵ��v�˙��������ȲV��:���M��R�x�}uZ���4
�:�=]�#V�t���Va"]`���b;iy����>���nWG��{�r��UX��1����%�{.��i�R��ܫ�w�η ��So3;���u�E�����C��N�I�>�ض���=ݵ�N�?)��L����z��H]	�j'�m8֡�<�:�ƅ�z�-c1T�ʉX3~�3�H�@�..�C@���pzV\$�]�9g��s޶o~^��=�v�+0�f�|¾�)�{ŞY=[����c��:�Ģ>繇m`�!�:���|.g{����׽�hۉ�]X��ظW�/�"����n{��{�n���q�^�|'��}4C�g]K��P�0��QZ��;O�ld�7�8Ȳy����4�KO�o|*�>{����^�'eF19�^{����|�7ϮZ{���T��;���#ӗ�a����%B,��U�D��w�C[x���Y�^7���_r���~��}lG[��6֕��p��ᘡ������ٮ3j��R�_rh�3���Z��A!YJ��z6��e#�h×��M�Y���:�ZI�9D�y]��h��S$�Pk��t*{�"��>4����ʬ���$xvX���]�o�㶮J��6�J㷠+���P�Y|i�ו/-�Y\"7w[����l�[L�q��o>i-3� ���Nۭ�Cv��NWAl���p��g'�-�z��4�Tj1(�T�i���l��0�+]��t�hT�J���x�5cԧZ�!W]w-��á��{5���x���R�ٹf�t�Usbl���A@&�K����y�Ύ_!�(�p���l�G�voՓݛӾ�J��H��Noh�1�5�o�㒩��g14��wMָ��j�V)�D�{/ZH����Y�z��k�v:r���V�7�]k}iラ���V[��*�䦯��t:_E�'�:��ø.ۺ�J7���-q��s��=���l����ڦ�ݷ˽&7<dBN����_mt�X|�y�������y=��2m��5������o�1�d����c���u��:������+,3��hɊzNl�'?(Cu��h��1�������` Tt+�}ԅ�}6ⵉp�<`�D�tԙ �~����ǝq;��.�1��/v��Ml�c�+D�&�a��*hݽ�G�����sgN��RiǬa��3B�;*����^n��C�EwSۗ{��S"N:k���)��jDf]M�%N��r�6�>!ȝL)�NRg���f��"��j��=u�t�WL�����%���7b���ju�Nt8����u����I�i���uB��yAU��T�V����'��/x	�aU���L�J���kyq�ˈ�i4��*۸�e�򜻭��=�[��4Oݡ��_I�j�ΩO/���������L0�GsəW�I{��k5�=��̪
�\�'���/�l��C钘9d�=v�Z�$C�����5�oʓ���H�0����-��*��J���̜��Ԩ�Y�Z\���ȯ���7�&�ˏj�T��Yp<)bKH����:Rғ�#�|[\羆�a��
�a:b�M��!u|6�\��:�!�R��D��j�t���Q�7X{˨�$��6�]�W�*%�g��;o�t�8�I=;���tW:*�o�Vs�_Zp�no�N����-�5YBz��
����u���H��'��Rx\v�d���c�Ѭ�hV��c�&�,"�EvI����/Gf�J� 	o1M��w]ɣse�I���	\�z-en�ݚٔ{rL�ƭ}�UZ��G]7�L�)^���p��"1'�+ovu#���'!��&��Q�Q*��v}W�P�u�*V=�Փ�eZ�/9k�-�3ݗ@��\���9(�N��;_%�n���GC3��m.��;����e�8�X��%-R�K�7˝��s��=�n��V�%�y���I�t��^�uت�fv�/���Z�c�fyy������]��ݴ!�M�n���3tF��%bT����=I�s��(�~~�2Dk'�5<���S�?i���Nú�j����k�yT��л~/�l_ ��&��9Np`�j�1���r��]�����$hʦ/�H̟�Ԇ�w�x3}���P����[�Y;PMS����ޠ��^�mK6�$��3O�C��-����[{q7�~ӳ���E�1~�]���U�Ӟj�|n1�#_��<�t�p� ���x	��@��̂��T��{.a�^�ΨR��^�N��|\���4������T�5��B|\ ��:�R��G��d������RoO�čP
H~Q�\����55�(��Yjm��v�=q�ֹqf�]r��5!��
!��܍N�G�y}s7"H3�F��ЀEN�ͬ�W��=U�����ca7�6��E�{���Q۷3��t��p&h�� ގ�\:EP��w*=�H�CP��ub�S2�G���]�]�#L��bʴ�BqF(�˥�e��^���[Ӄ:G[�26�����f룇GrNQK2���N�Yȸu�ZЩ
�g}���T�g3���U=�:3�YLf��ӗM��W)L����[	�=�ʗ��޴�RQ�/�n�Fem$�YnVuĨH�5����b��=�N�U�[X�`D>;�7/r<*����r��)S(��֙]q:l�Fo:�Q�/����YV𱓱�˧aD�	��ñ|"z�ʆ��S�����2[�y}��b�6ҝ�g.n�<�im-X,Sv�&rufΤ�e�T��X�5Т����2��t-L�Ӎ��l��6�-����*�'.g1R�fu�U'��a׶�>{9q���5"N���{$�$���)
*�+�vs9������DR��Z�j�I����*�w��c�u���4�,m�����j�O�j
�e�yYfi�(�%�vR]��0�l-fh	O	��´�ј�-���ƅQ��e(co���S��PoQ��:�R�t��ۍGҌ��&d�$�έ&m�҉�D�]����w�^Ch�v:���2��׮�A+�Ǻ�ke5t��6��$e�˥�^�>�6��x=T'��^;��[�'7v�rEw|�	G&WM�V�F��1�O�#y�^��˸�7\e�h9�δW��˔�-[u�-b�k�p��kn��Xd��v����w�ԍLK�;�0.	�������Ҏ?��ޢ����W�^����wu�ś��e�0ZF�����iY�0w�e���AHl���ŭ��V:�6M������(���5�>t�bG�����5werY#��s�d�]O�@�Q��	}ԗs����1R�β]�Ӗݧ� �8C��ş,�7�o�X���k/.��v�ۂ�W�e�w���c����3,H�P�'���0�M���Os@S��fBV�SQ�C�3�yn8���mw6��!�����ܴ��Z�+n���B�v���O��r���wZsl��.�)�Rb����{Vk��!mJc�����&��	c�����#4%�}��NXc�:�U{��Z�B�ͮ��R�4���ҕ"醻w�F�_L��蘢�OC&���ԛ&��y�t�Y2䝈��>yʗr��Q��S�sT&���3��Cn�	��jm#ľ[���m��C� �붲�f��P��V1�k{$��U�L�� �yF���m��.��������ʷ�H��W!w�!-�W���4�fe���!�@��\�����7��]w`���Ia� 'n���3&*���.�Q�ڒ
�R�݇�THR�JQ@�E%M%M��%R�AT�HD-	@DHQB�R�4�K@ELAH�4�ST�P�	TД%-
4�%MTPU	P�UIM+M	4KH�*�RJ�P�H�ДP�P�A@��!CBR�E5T�!M!�$T4�P�%R-P-!J�HSBR4��STP���H4�4��JPP�P�HСB�R%R�+J�H�"Х-R4� ��Hg��y��;�:�]�a[pD;��Ox�f�����;#�梊���� �<��/|K�n�m��Y*Wc�N��FLZԲR��%��3Q��<u�l��u6Y��o޸;~�����U$4:�r��6�<W�������懩�gr�Kz�i�x!�O����u���b���&_���t�ֈ{{М�_����$.��c>�u:2ɭ�c���a�UA5>%������|`	�C�o+����]����RmDu�Әz(���xuw��1�WG�}��f����x��\�u歁��2/{ї��&eX6;8�W�t��^�q����/-�f��Elv�9ɔ���ۻG>}��o�u�]��C�ΎLߔ�Q��·VW���z���/,��xF_��CKs�I������ǲ%M{L'���L�;�~���NxΜ��A�ۙ�~��P��>�9���\�������t�v��`O�~�3�T�@�^�g=������v�OdOT׽��9�s�ٞX�G�+}c��KE���,���m0%k���y{ c�������66B2�Tc����f���PŞc�����Y�R�3|g�ת��rWj�������:^���	�~�`7�)/��d�Y�RٛR|4r�΋��$#P��\�M�O]܏BcS�gg~�F�=}���Xr��/B����\ J�8n:���qO%#�s�
}(wV7]zy�-u5�����5˖<�ّ���9۔�xQ<n�gc.�D�+zV��Ȥ�¿z���\���)���a��B�"Y�R�M$|���3q����Y�����uY�ٝ�:�Vf����#�ۛ��9^u��/m�:vK�r�%W�<yL<��nbm�W�����{z�zO��G�hMv�ߎw�x�9��G�_�\>�>���������A�Ѻ�q�btI�t\�8[ԧ�]��m�b���M�E�Z&�;CFB}�h���z�޸;z�ه�=�>)I�E��{����<�<��2�>��K��Z�h�r�!��؇��&�=냥�U��S+��P�E��:qƛ�E{�5><.�Hs�s�/��"�Kz�a�*A�<K���� m�^m	����N�i>�j��U����Uz���d�� s��E�ڸڇ���9�t*0�Ϩ�����*K�E�
�W��� ~��;.��1p�O�]�:���;����/�^�3�ٵ�o�:�>�}6��ꨯ���4m��{>�e�w�a��`���s�t��l_�,b���o�ntV�:�����ь}�Q��ϠO\?]��3f��I1�
�������]�c�v;�H�sv�z��i0�K+9�I^�]<��V���iI��p�-ћ���% hmE����o�&u��Z�Õpk/�umL���p���Z�1�P�;v<Y����'s�mar%:��i��A1�6�`�����%-�d�^�������,�9�l��˼r�u}�Ӟ�3��p��Ma��f9�d/���$�٘J�lVW��E9�v�i�&+=��|���8�yzn|ğ`�~����R���w������v�nC�'tvG��QYU���XV�de2����D�R31�q;+ψ�c|�}�y�}�9��=�4GY,F�*��Q^���F�S��W�˫L���wo{J�|�g�T$�x���q��z��v/n1~�[%�$�Q2¡3��9ޜт�����~EzG9�}4���Q��|}G>~��N�ڋ�GYZe�jH*aOA�s��zVz����|/ꞮU)9ϡ��uo��2;��cr7�<zߝǸ9��ox�uSR\��[	��X珙�O��,"EArٸ�����/�Oף�����<h_����I���T(��	º�GxvԲ���A������Y�|k�{�&�5�z껣L�s7l/J���>;�^�M��ު�+_���l�<�$q��u�K���0��������߽�8��ڭNG����	w�;n��~i��	�O��=�����M�Dի���9�^��m,`���w;�w��z¬��|*'�c�Ҧ6
v1�8�_J;+�s����jʃ�}0�Qa5|zoNW[r�nn�mA�9oBQ�B�ͫ��zgx��~>��n�z���j��T�.Ijl�:~ԅ`��4��7e>�����k�Zj�G�>D�����s`l?U��n��F�S$5E�4�H�7�ϼ�{�R�M�xи�+M^����!��Ra�o�h�{����2*;�,��z5���a}�η/�%x\�t���m�ȯO��챵����r.�����������~�>��]-���Ga��FT
K.d�1��a����7E��du1������J��m��Vs��3��~�\�'�5�ua�NCsC��=ܑ��D��py��P�'��xNŹ�J�v�حp�-B��K��B��i9ׂ��*�
Y���G���s~S��ۉ����C����<��8��@;�f���}�;'O���1ڕ�ϝM/1׫�V�m�X�8�����ǲt�̱�����ݝ����'���p~�tx])	MƖ�.�W/Z񁎽~�[�W������s۔m�x��^��qK���}�L|/���\�k��$SOC�l��Ϡk��1���~<�H{��ڧC�ϻ�^���Nm����2�6"xm�5���[�{SZ�[c'ƽ�h���,�1ݑ����E��k��t5�,I�G�{:�fec�����ȶ�u��pTz'YO��ۓ'`��&�f��k�5w��Z{z9G�X6-Ro�|f*t����]�؞%�3��J.�f�{�f4eSJG~���Ԇ�����p�x�W����$Y�ߨ��37���V����y����Q%���0|��l�L��r�ۉ�rr��33{.��x�w�ϓ��Oo�i_g���~�Ӳ[ 羓�L�Kg�>����aWe����g��m�Z�ZG>.w�q�~�������f������2m���u�z3�ݼqm��
�<*������[f2����ӺM�z�����h9��O4ヱ5꽟m�{5xψ��@�:A~SB����@>
�[�CmW���g�x�j�2�؞����b�O�!9�G(��q^��4��L��p'��}>��d���ԮC��������S˫/D��k@�{ ��wDr����J�"6�:%�n��/�j������ۃ�gT����5�ʻ��nD�yQ���@z���d42��F\
�βfU�6���w^��qE��S����|�Fǯ�}A��#�y�ݣ�����j|+_�F�I����TAF�O�������͕�����O�EW5�Ӣ/��
��p�/�BϽ�����el�("_�^G�ǆ��۶�%!���^��h��W�5�Ҧօ����B�҈>����2u���[��X��8լk��u�4Aq�P��>[�a�SzAkF����Ci��RE s;��T�ƿu�ۋ���Z���&o��B~����W��~�}��~��8�H;;��2�V[�'vu�:��]�B���NQ�qJQ;��o�~�2Ryz��xϏr��֘7�wy�y��c=����~�}:N���YP%#�VMi�@����hr���1�y�\�tbz���Q�������5}�:j�N�\Ɵy��J���$��w�n)�F̏�
�ފ�Ϣ$:�w����5�yHydz�ϝe'�o��u~�@"Y��8��䏑M'@L���Q>�����M���aϵ��{���~S��^�K�A���.���_L�ʡŮ9�����U����'ܠ��/���}1���/�>��_�[�~ӝ�/�o�x���W�����gAe�4#x:P�=�Y�|��}��,�}�>򘺙oӑm։�N�џ'޶��zF���z��Ǯ�|YGU�NMEs����[��* �@�[ Q�^SX_b����W��=�Lk��Vɀ���&��zb�����?��ܺwUk��C��  _A^��q_lif�%�H�˻������1k��|z4��%�e��K3/��PM���V
3��~���m6�˵:O-rqs*t��m����B�m��ʚ��Y:j+��ZE[K'h�7t��\�`�wZJ���(×��NA�ZƶJ���b7k2�f-�TLLC��r2w:�G5���w�H+���듡�p߫@�׮+a�W�n�Z 9�}^�t_��j� 4`��nb�c}���5#�^�������@����@u�W��~��zf/�2|�q�_N
�)�|�	]�6=�5V(K��e�A���*=p���-��h�{ޠ;��uCn;�0���9��F��B��L���ʷ�3�S�:."���\l�MF�ˇ���h�C�Ez�Ƕ|'���m�z���7�yL��=>�}}K7|IQ�7#'{ꕧE�zt�҇��0�W�FC�P^���5�]�ty������K'���լbkϛl�w1B��o�x�������:��L1Y�ˬ�F�g�oB)1z��6�/u��GL_��P]{$h:�	��]���s��xP��x ?���m�=J�j�X��D�]�t�#Ϋ�|�a�i甂�:�+>��P��eᯌ�B��R6�v\M�w�1�v;����0>���.��N���~�\{�ey\w/m��o���$��e������ee[��oGG����%9�S��6�k���@��>>���_��[��dAu��+L�|�c����8v�+:#��#���-;�Ƥc^)�.d-�揬��+����1�'\|y%�Ԃ�ʎu�Y�S�:*.�5+fb�b��Qy6$�᭾���v�\:��q
T��.��jb���R��-��2b�4�Q���bTh�2e
��2^��˂J+���,	�3�K�6*���<��{<4w���?��<z��q���$rɧ���5Ϥf����ږmItg��"EA��n*e�n�H�����ϗ��ʱK�WB��V�V�Ͷ�S���}�'M����������3Kt �Ut	�ƣ�^��J���4��s$�䈤��=v�����Hq7�����*���}, <����P(t�>�*|{љQ���V�8�}��C�O�����������?z���U�պ���©-H vx�� 1���T��N��{��ѹ ��\j�j�G�>D��>��>�� ~��#]ez�U��,��}��՛�՗�-�mX��-�ZkKÿwz�w������7�O�w��ȯZ��[�]�rǴNt66��O���A��al5kݏ�����d����1�r�܋{��{�
8J�ge�7�;�@��}�"��ܣ*|�\�W��wL9�����Ɗ���a)S7M9�'/����zו�Gy���=V==8�4:�����TIڀpy;�Ⲽ�4����{��}����̒~��yy�К�G��nf��R�5{zȒE���7�	J�r��lT���|t�Ǒ�V��c{#���ܩ�~=���.�9O���R ��U�5=Y�p�U��<���\G�7Գ�ݖ�Ò��w%��s�5>����E��eNr仿ރ�e1US�r!��^9��W�,�wf����N�N�D��Gӡ�����q�"��ML��	�U��21���T	Z�Ǳ���ϧ|yC��%�*�5g�3��Ӿ�o��G{�'�u��L��\�JCSq��*��G/Z����������a�mPa˹�U
}��ovzY��p�ve�����S>F��eF�Q����_�c�?�汐o%q0O�w�;	y��E��n�ʏ�t��I
y���x'�.�{ׁS~����}��n�V�� �o�z��[���9/i���������c�-�$w�N�6|��|@�����)w�}����nG��o�q�j�?]�z8����<�n�.�q��s}~�dR�;Z�U~�}F|w�{n*�t�#����:�#O{}R3��V�?L���pB.��>�*��s��jw9�����楊ϠƱupx��ٌ���l��};��?z�����`fS���qll���ޯ.�M$���H�4%��� �*�oY�W��z|����/8�Twь7=r�� rj(�f�V�b�w�i�A�6�B	Hm(�]`j�M[J`/d3.�P�qEիi䳜�L*�b��]�T�հ���U�[�uǒ��Ր���)o.�����59]Ɵa���u`v�0tTy)؍�z�ή��rj?�������=�TmL���'��K���-l����J�0ڪ�1�S�(��{|]�n�������)�.�Ty��M�$����TK��9_���C�6�k}n��l]i�ɹ���Ǜutm�U�_���fE�������l>6vp;�V��Y��������oyǻ}4]�G�i��/.D%�rz��mO�oC����ΎLߔ�Q����+��uro��`l�W�b^�����g������)���}Y[M�#�W|ӿ��g��?V����s�t��tW�-���t���
S�Pmi�5�gE��/����/�����>�E�,�o-ۦc޿V��?)�	~�c�{�>(a9���T	�,\VMi�r�����Z�.W��Fz.OO���~�3�ތ��[���|���{r�Y�R�0��A��w^�F��F̏Y��ņ�}��^��yow�Nmԧ��3���u/zk~�W��z��Yh\{�nB˔IF���hd���F~��%�yX�K%��(�L�����Y;��9����#}p��+μ;"^�>;%��P$�x�O��Ѡ������,�}M
\b����}i��j#3?nے*J#�����Wx��^�U�C�j}�
E���Fm�[y(����"	6���K�ǚ��m���
�ʙH�%,�3.�k�#��nt븅N��wjAE���*�8���s�2]�7��G�P���Q_^A|N6�5(�u���V�wD\�=�t.���Ε�ү��/�S���n�)qgN-����g�fY�xa���Ң�Uk4�0V�������O@�5ǻv�nq�7�T�:�� D0�܍��]���9����tk\���U�o���A���i��B+�"�{⑛�9�M_Id܏sM��`ѫ��]n�����u��r�Z7�[௳*
-�9kd��v��3�����y���^Acv+�Z�*��;��6J��J�B��vL���*�ȵ���`(�r�Mr�G(�v�v,�:Z���i�'�Lbm�{]Ǣ���;-^��v�b]ѧZw�}/���(��a:\޳t����ҡ{�̙#��V��qb��(��-<�[��1R�;��r�a:��yw��f�u�-������}ˎN�d�.Ԋ>z�X��F̧$�Բ�^��"��t�sԌ�����%��u�AJ�v�GOl�-��o=[�;%����኎������2v�cHP'��L� V�����۝Z=�M^4�n]Vz��Zz�/�U�<ZP���o��`��'[���$�ti��bAw-wD*���y�P�i֨U�`����	�e��:����{X�������s��U�h�5 Tt�;rT�ޞ�Y�NT�IutF�L��/2w9���j+IR�n�v����;M$� L�ݢ�c}.���������|�� ��8��oQtM��u)�S���@��j[2�ïM������;k�t�c�f4w .*�,i�����"������hS�W<�x*�D�%�����7����
bS��xJ$��]�kkNC����*ҔĜ�����
�<�t؉K-̷�P��W�f�ƖM���Dz6ti��2{��\���q���Q����Ⱦ��"K�Bs�I1Y�A'V�ܴ��M������r9�0Ώhl*������be���si�l�l����_r&�]��:��雃kC���Ǯ��a@tT4c�!�UV�	�U9���B�ʩX�Cg�������H�	��^l�$���:��sPc9r9��y���s):�gVF�A٬oP�W�U��B�q����4&��mG]��T��t�=}7l��s�*4���n�����v����V����Y� [��!���q{�F+*ʊ��򣼓����+,�T��6#����ݤ�p�n���� 7�+
�N�"��N���g�o:�ʃ)9Ō����c쮾�N\z��&z��I�O3>^�Z8�k�����w�����v&�N�)�᩻I�*��ʵ}F>��=�=��������r���*��
)ZF��*��"
U"h
 ���J@�����)�B��*���D���JP���(�)F�)"R���*��*���(�(�hJ��i�JQ�JhJV�����
����F��i
�J��"h�(����(J$(B�
D����bj���
��
����"fB��"�������(
)JF�����
i��������n�ׇ�����#ɼ�q
Χ�H�#9u�f�nɗ+���]�l!�;��7ԕ�u��\��:�hC��av�W�=5�&9p�Q���~ȿ�Uy��sL��>w�9�/�o�x��{U��>���G�Ym�Q�F3��X�e�9��w���`rsS)�rۭp��2!>��w�#O\g�pw��y90�h&*�r#��x�F��/@��P@N��1 �@W���V/_�y���z��ز{�W�'*�Vgt�;~�'����p���[��f�� p��]F���t-�!���U��9�����\V���}�u�^@���6���.>�_�*��W�P$�@x��Q�/��{��*w�4]J�t�z�Y�B��\y�����HG����
~��7.��S��?�3���BeW�>/?R��JX��Q�!^�������mǲwtm�F��P�s#;�,�)��S�2;(��mC���n��@���R���ׅ\l�5����/]���Ez���@��~���w1f�#����,�>��p�|,Οc�OW�&��֏I��Nt�҇�7.�1���#>}�ҹ/z5{#��@�#�sp��]�^��-�T��)$�Z'tÿ�+�n��������	n߻�J[���̉*�'��	��:���Pwm,Bޓ�WB���0;���R�P�E����6G�a���f�W����~%N/��Q��U��n�ǩ-g���
�����HUJ��l�u�i���n��C t����f��#7��z�N��2h�̱|��\���}Tק�d{zW���ݨ|�����5��KuM��^i;�S;D�#~��U��TT�b����B�U�S��H,��B��:�+.p�6��xA�YE��S�ސ���
�؏���$F�v�P����o�ˏx����;�{���:�(dZ�J2�_5����F�gi]>�P�	����Ģ��|S�Q��|}G����+��֢݅79�l���r�����L�XH=�3�H).�RU>NrMW��g���!�cr7�<y�
ݏz���<���u���O�o�.��Gö���D�Fx	�R$̒���D�������L�L�]B����s[~�;��i���!:n����>6Ȁ�|f:�n��ҼUg�	��'�y@�xǤ	��3~���'��{Ϝ�y���&��z��]�p�U>� sĎ2[�X����797��/YM
�v�^�Lr5��;��m���;��;�Z����.=U~5p�K�-J;��@�K�6��7���x�ݯ
�����}�Q��C����ǽ>D�����X?U��䗊韦z=]��MWc�8�)�,�X�:I����\.�C�(Q�{pl�&B�Ը1V�B��5�	®�s\��;�d©���h���{������ISa}7�:hO �p��Y�Y��89|)TJ�����oo�����n\�v�r�k:��"짩�4&V����mM��(��$.��`��46+Ҵ��5�w��p����o�h�@�G���;Sf�B��V7m�G��B��JJ�1���K[z%�a��ckU�9z�ES�2�j��f���R��é�R���o"������2TQ��'tú�n��/O���
�Y䴌N�z�{ǫG=�!R�`�U^㏽CƳ�Cӳ��4:��rFyI'8F�;�r|�V㜋�q�*�g��G���k轾�UU�'!��^9U^:�7��~��`]1XA�pk+�EVR�B��cg��� ��:�7�D�q���[�q�=��>����	g�w�ߺwfx5w��\<���gb�<Q�L��&P늕GD�<���p9z���_�Vײ��aZ�g��=�ۥ�m��!_��8�}g	H.��}3�n��U��Y]����W���K�Z�=qc+�U��(7��S���#�۟���y2������U>	�[�4<��i�M]��iϢ^�O�z��H�z�z}���ږXD��c�O�ʡ�-��)�vۊ$�Լ�w��Lט�9�V3�Y���.N��ʵ,���v{���.M{u����bW�j�5�\��B�����)
#�Ϛ�Jn��s�Q�7���ps�L�@]�U�}e�.
�l<�C�b^:"&��J���Q��V#�m=��gE[����Q�z����n&�U����<�_���n=��m��w��;%ېrG QѺ��^g1]՝�Ӱw�=._�є}�[ʊ�t�#����;�4�Ƿ�#n#�V�?L��&�[d͑=�EE\n�A�b<4� o�{����B�ƣW���ف��l��Su�_��S'<�D�z.}�h{�U>=$�.� t���N{�pKz�vڿ2=>V|v����^�tЃ/L���@�<�w��d
������Mz�!�=F2_W��k&�6X��R�u�{�$����Ԏ�����z�K����Q`k���������8#Y��i���-�N��[��ڽ��=�O��P}����a�5E=����}Ƚ�F\
�:əV����,������m���g�sǸ�q���7/.=����}��\{n�+���u��ɛ�* �4��g�8g�sy��Is����%���s�
�ҋ0�T״�'����UxOg���N��j�j�Ο���2Sޛ3�Ϥ�����NI�(��Q����vC�����̝�}��R��
�T+d�f�a�Kofn�� ne0�e,N����Ӈ�k�w���lA�b�h'�=�V�hz�7r&�u�Vb���\�2���\���c�Z^����!Ξ|y�8�l�t�=�m=��b놼��-ܘ����Y���z{��O�i�}�sŌ'3`�<��X��ɭ2�Y,]�Ge|�J�(_��'��B��K}ʩ�K�]`�8���ǹ��4,���<5z��z�d�Zf7j$lM9�)�z#�g�UX�/zkc�^Y�Có�Yh\G���,�D�j$�k�*��{^��v��>�܎�4�}�d8��]Sz��|G���B}2Ա�ep^�Ӳ]�@���>HU��nT,�K�{��u��򘺗K�-�37��~��#��q���\{U��>���}1Z�z�Ӯ��ԍ�}�R�[���7�x	��@��$��=�h��N�џ'޶��zF�����W�)�q�^�
;1��D+������p@N�2L��J��X�^��;`Љ^o�S�k�*���n�{���:\M����~���[��f��+��n(�>�v�-��L�}�z�cb�@Z���zB�߯�>���>��%�Ӏw���W��Sh�-�G/��}xDr��W��'vJ�w�eםG�Ԍ������ޤ�z� �C�_��ˬ��Z�>S1ܠN����8j����&PS��
ʎ�|��3j�mP���Wl�2��޳~��y�H�x��V�x����k�01�]ڽZ��TN�������O�U4��Ү��@E�̾C�s��n�5h�5BK��c�̮�h
��T�ݚu�Ǔ�X��+�R��7����T>m�ѷ��M��@w�:��ޡ�C�'�l1t	��Oe�jUn�*}�_ç���ߢ�ׅ_�/M}����/]���Ez��{g�'�����}Jwj��ϫ�]�o�g��f����Ta�(�����t]9�wJ�.�1�ʼ�/ފ�z��=�[u���8�)�q�k}�+��۷8|�'0�(�a�O��8d�����𜻉�Ⱦ�(k���]`>�:������b<�h�v���p��3||��Ui��Ҧ�G�����W��(�;'���v�d�x���|�_��Y�y�~�[%Q�P͙x\��eQ{6��]/2=�Z���U�tT�Ɵ@U��@rr�}O�eǼVW��v/v1G���C�2���LX��Y M�^Ŵ�sĕ�|2��qS)L_��'/����L��|}G!�_��:�n�8�"j�=w���2��~�}����i�D���,eJ�&O�����uq��3�!�c^{kk�D�V����\��w�N�vAu�1��g�eX<��"���u2��[y�Dͼ����3ƺ⇔�lAAa�:î7��Ҷ�Kk71q[x�MңC���]b-�P;�\�Q�@�ړ��P������&C2gS��ө�[>) aqkcV�T�r�C9�qG]8�2�+�t'm
���a�������z9fVnڕ�3��%NM�6���������'��ޑ�W���/��/�mO��2 'Pf:��
�ҼUG��W�/�����yAql��q7�,C�y���&��z��US��U>��@r �F�F�]���s}��w�"�#���.3���r=3�}�=���?z���W�V�K,�FY~���W���5�N@}z��/��_�b�P�5~�q�O�>9����|`J��ð)��z�������#�z����#��uX����	�Xkce��Q5U&97�4uu�*��C��q��b��5�o=�7}�lW*@���������c"Z��,�tl���j�����Sjo����P%�e׷{�2��#�w�T���	��ȭ7ތ�Ys%\�}p'tø�V���wBz,_J�EG�oj�*Ї�3�-�T���P��U�OK�绒3�I9���6wj��k��vz�M�Ȫ��[����ӣ��ۗ�ኪ���w��*�
Y���NI�p8�������=1[�D��߹�u�Zd$J8=-��I��K�x��jN��������nQ����Ĵ�H�*�޸�� g�n޴�T�%t�!�͍�E�:��W��oHY4��
�׫c`��
�t������z���Ԍ��99k§=���r�넄`o����%5άcW��4d9�x|��v7I���-9Y.e���J7����l�;s<2��\T�:.��)�,���^��z��!�~7MX~,��Z���%ފ�G;���nQ�8JVe��g�S>FY���C���
��e`�>��ѰMc��� �B��'<�z�H{��j1�<���r3F��b�����O�|ˌ+��~�q~��A��{׃>|'��o�u��Ǹ����ɖ\2�.��@�>U�>��(�.�{Xr�9[��2KϢ߶�o�N��x�9׾�=��ڪF���~�9%�s[N�¼<o�}�F>[~�=;j2��2��~ʇq��p���c��{�ꑝ�����o����+�쬌�<[�g����d��@�y�P��ƾ�W���ٌ>޶ΟN���� �s~���~��ѳ���wwŋ��!$&��x�x�����m��T����2�}��!znzꚋ�	2n�x��Y.��ߟ��n��F�L�Չ�1Q/��n(��W�ǧ!���g�`o�A}��V$�0�����x�G��� �0
��.�W�y~��'��먯��n��w1J�Q���YK��h��,^�y���N��R��9N�Vhŕ�g��Z@�]�x������.1I>�)ppmv�s�`�ؕw-!���ժJ4��&_f.�#�0�1�<�8��3O0/��}%�ξ�W:<D�cW=�5��^ž̓�~L���8����߆6����P����}��ˈ�F\
󬙕p��r���ǎ{�.-Ft��cռ�=C=[^�Q���>�/MF���Ľv�|����j|+_�F�:93j�� c�7>�S�K6�AG�A�ѱ�C��Cn*}��Ҽj/o�D��i���/}U�=�t��y���u��J�l����x�_�?ҼA�Ή�P6t;���:%����~��vC
�<��ɪ����&\c�ԆW/R>�5▵kL\{�nx�3���A�yQ|�Y5��)�WL	�%��ze&�c{�%b�z%%쁎�����X;�����������0���u�r��Wo�G�p���Z;JQ`'�ꠇhr�=�4�X}�]����:�B��!QD�z$�{7d�#,O��ѱ>�8�Q�����e��w��r#}#�������^u��/m��t�����eT{��v)o���G�GI)�lT��9ni��n��>�H�|s��Hg���힇�^�o��
����v���G�YP O���k�|����~��n�MçhhO}O��]#������x̡5���� �+� ykҰ>�S�.��b1e��]��b�*C)�s\��$U����~E�mg����M��V�.E�M'��#��nl}��A�q˘�n�Q�!��ʷ��K�jƃ@4��&�����b��g�g$���q�F�\�Ww������ t�-�(��)����������x���[�O���"��hg1��i>�z���W�+a�Գh�A��W�����p�)��WWU�7����.%�5vH�OΘ�sĿ@���7���/�~ȫ�U^��d����m�C��x�ϕ�޺>���ڿ����Fa�6��}�J�z� �`u�?Ux�U���U��ad���Uyv�.�).��>96+�j�U�O��:��m�m�Q_=��h߽���T6�X����J�=o�n����!��d{�u�ON|nPV:pz�V���*�6^�Uuyz��ފ����\I��l���k��� N��T0͛jI*0�[kC�����I��CەV�z��˳�{�X�W�Z��}�?���N����ʋ-�Pex��1�a�e{��9�w2R�]ý�=VM[�T8@Fw���T�A���ӝ��˧�ݻr7!Γ�pf��P����",aF���2W���}wī�@	[�d\�R��7�v��Y綅ǹ��Ys����B�:�o�*�`ڸ&`{�3�D�3ͧ��a�5H�f�8��ӫ���`c�z�2�%ܰ�V�l�B�%Zj�]�{=��'HF�BW'v�t�~Ǔ�L�-�6���{+�t�
e�)���ZN��:����y0�����i����s�~yS�&كLj�M�fl��m�I_4`��{n#����WQjiwK��h��U�aG�aN�t������c��Vf�ad�6�:x����<�	2��O*\��u�
%A�3P��Zr�7����HЍ�o��v^�3-���w^N�b*�R���׸.��:OS�W���<�R����㕯��vZ
剴kp�p��BV��fr<;:}j��
���}�<*7m�JbLm���;�\�V����/�Cԩ�a�f��{.����◷��]�*�Ӄ�Ě'��{��b��m�j��j��nnV�H�Ƿ�p�v�K�t����0��Mޱ[������כ쭮K��<��w�F�#Mʍ=b��p�����h�f��wqw<�L��'�'�Sl���̬�L�]-J{i��-��˦�J�Bl�G؏f�\�F�\�B�"��a'WQ�;m"T8^7����ׅ6��o`H���wj`FT��+�����_9(���(=���wv�*��WU�T�wwM�3��#�yy)N��F3�Ǟ)��-�����K��i��I_����3���^��;�a�wS����|���"��v���S�|�sr�W�rQթ�^vTݮhp�f�}����h�wa��X,Z�ݝ��`�r��ܬc�����R��Ӣ�h���k�ʓYR]���kK�BZ�{z4>�`�f9��j5���ܧM3�]�6��@��{P1��E�s&�ia�í�o�9��
5y���y��cԔ�-�Ɩf�c4mdt�6��kY� �=��EH�ͮ8�G�����	e65�޸�iӍdS���3Z	�ZQ�w� bu�!�������xk.P͈&��w�N����U��¬.R�^M��yR�L�t3�Uk��f�J���'I=�,�J����gdYٔ����&Sۆd�C�Y:��NW6�'݋���R�#�u�k]ÂhH�c�,��}���ʬv1`P���>����2�o�V:
�gj��$,ҋ��F5�S�7�e��)+C0�3Y����9�ƒ�qH3���9��M�B\c����\��2NX�鯺��j�;��kp:�m�yi����us2�gjH.A*�,SpN�����[�7�GH�]t�1
z��Y�H4����ޏla�w���.�����T��^e�E�q�e��8dG��ɀ�Υ>9��blhK�V��\�8��n�N��J�57Yg��'�3����4�+���m��-I�׊���u�ع��s��ͅ!9\ʨѽMV�źN�������t��E1]R����'K��^��w:��b�Sb�]E>���RYu�����((J�h(R��R�$"�����hZF�$J
��JQ����F �*�hR��J
Q*�
)ib@�����!)(R��
�2�%2b
(�)��JU�
) 2\�'%�� �\����h22��i
 2�,��B���i
��P�)"H�(�'$
��
F� 2����(
�+c�����K�V�)
uݡ�S&Ʃ�v̵fr�zkh��䜄��7Rj�P:�!�O���ʍ�����W��������UO����q��F�@W'K�����O��wн�Ÿ���k�i����8��l�={$�_L���I��r���^.;��1�Ϗ����c=ե���f��ޛ��г�)�F�T�2�"A@� �.�RU>Nq��u>�xh�aMΔ'�U15'7=�؜����{�<zߝǻ��dږXD����H����u2���w;0�"�s2߆�)y	-��Z=��=�'|�~��ڟ�D��t	�� �>��=1������(��{�+Ƹ���c|k�^�rՠ�s��{b=�C���doz�ا���̀<��(nǵT
HV{�N�Y~|{�x�]w�a���a�~��zgx��O���{נ_ު�������<7�T�=�Cީ/��$�t�I|pf�/���&��o�z|��Ϗ�|O���'��,�P�.�V���ͿP�D���Tn�\�.{Ƅ��5����wz�w	��0�;oϲ���վ�������>��.<��6*;�,�Q��+>1���k+}N}��e��{��z�����B��\ـ�3�N<���㒋��|�֢qEG�XIR���$\3�/U�
�_�Th� Iuֳ�e�-ͷ>j�lIh�]��y)]��뵶���w42ѠP]�keŪ�!���z���`�}c�ed]Z�-Lܕ�����BO/�����Ѡnm:�Hݥ�{��܋{��ߧ�O_�Eiu��]��G�j��,�^_�Cۿ�Ӏ� ���5��ݾ�.��CE}{y~�W���P��X����{�#3ʉ;@��6i�:��`����\��ў�)W����;��5�}lgʪ��ׂ���Q_�����Gnd��T�55�S����N����<AG};�3��+*����F��|�=Φ��};���n��ixR�d�����{��^�|����b�:v�e����'�tm9Si`*��Dr�����_�nQ�����.�y2�^ˎ�n����=�F���A�2��ē�v)�eF�T�ImM�y��E��5
�9��p��VC�?>�=�֣�۟��*��y2�������?h��߫�������5���]��~����;���~���9/i����%���x�� �f�O!���Ͼ��<�[{q7��J�s�#}@{���U#m�������/��/Nfqm��c�:��w����G�P(t��2��=�n��s��|W��F���o�F�H��xfb��^���ﻂҍSΧ�i&+a�UeQ�aGN��v��|��O"��wxu��wm7��'�rԥ��+�[�e�2ޖ�k��WE�̝S�t��f�isp��ܨ�}�%!�:��ɀWF6��X��C��[Z�v��ȞǁFߪ�zU	�"�"d��@��҅p/�b�����0Ϸ��]��gц�9�����FV枇;~�'�kWUU3C]UK*Ip�:A^SB��x�D����_�,�>�Tzy��QZ��G���e���wļ�ꌁO�늷S^��!��b�_W��Qkf��,ձ����]΃v�?B}r��Wt-7^'���3� ;����y��J�#�z�	����^��Fob����+N�ya��ڸڇ��{o�utn���\?_����9��ތ�u�2�c;�]W�no���n��)��t�t�Q��q�/Mn^\<��v�>��>ڟ
އ�ڽ|R�:��{66i](�o�����|rPWgG�++�n*^���Ҽkr���J��O�;�����\�l���w>��ﴶo�=�� ���3�*�����:6��'oe���cݺT�\w@�ۼ��Ի}Щ������Wa�neN�C:N�0��.�kM�9��f7}ۻf�ʃ����.��n�q<������+Ճ��{�Ho��"��)_�f3����H*
��"�ZS�)$!Mz�.�"hZ�f��&�Ɍ=[��^��2����/=�;1."��1W4Wv��M۝ӮN!���Ov���*jʬ�g9j;�F�a�s\�H�^V�H_*ܮ��d{x��y�ڋu��n~�f��5�v�v=1F��l�AO~�?��H	Xڠ�ϴ������Mo�����]����/�{rIG���̘��>�c��s��q��G�����&o]Sz��>�H�{���9^u��/mB ��<�Ҷ=	��i=�s���g���C��nb�}I��sL�Ʒ~��#��{����lW�b�f:ǈ� �%нg�}}]o��p���J��ڙOӖ�h��Ӵ4m${�WY�]h%n�^hH/�3�C�W�O�8�L�� s� ���^SP��e_ym�Ϡ]o�+o�Z^����z�2=;��lC�.&�=냧�^��&e����8Y^��:�yI4f%�g�m��k�^�d�-�;c#��D�>�%�Ӏtz��p��(Z=dw)ao���n�o�mx#�^�Qh�lǼqq�o����ǽ�@����X?]��Jn�����ne���<�f5_�$dWF+{�E]O�v���c{�p�wtm�F����qݔ�Fd糳�=�5����*E%X�ύς��NIZpK���j��y�۬Q�Wx��͊���3�M�����<�Z�'�e��[���G��pazƮ�sX�zme�e'��v>ڰsrWmAЫ���)}ЍA�r�fޗ�(L�o=��D�����-�k��)�)�6\l��'NC�^�p4IP�O���s6�w�ƥ���9+8_j\��G�7.�u#;�,����U@Ɇ�gC���Γ����&V�TF{�sɑ)z�w��!��w��g�ϛ�>��b�����c0n�i���{6_&����������s�^�i� =Y�~��z|�yzs�hy)߼��\y�r�U{	��ȱ�o��eL������o�ʙ��<�WL0��"�z���u^�;�m �<�пs���)��(O�%�����ɢ<IC�/A�Q��*�n(�F�O�*��NW������ϫ�� �ܫ��w���ѵ>���ղX�RIU2¨<�L�L\S���Ϧ�^@�T
�~���#k'�Ƥ���)W�ܪ�cn	��G}�'p���{�r��4�q�c�|��J�/��r��u[��(�Ƞ�3Uom�O�yб���H��yT=�[�Ͼ�,�(���,�Ų��wz���f��F.�w�k�ׂG�{ס{g���P���Bp�C����k_����UJw3��Q~��d��Ӱw�{�r�Ud	�q���*��X�C��#��RMǷ�#�=wlU��U>��cR���]����%�A/�76�Kz^.>��^�'��*�N�a���ϙa^k�kkI�3X����"{G׽��;�ȥ�oR�#��e(uj�\��დN��5�,=g�du������uj7����p�z���{�@j�zJ�.�F�$| ���z�P�|}Ya�\j�߭����>���{����w|z�>�Wt����.�vi�̔=�'�o�@���
���΀_�F.55^����'���l�v	��'�7��f���
�V��+�n�\�.{ƅ�zV���������>�2(�s�삷7̉���/z̛�z}�c#b;�,�Qy^���yX��-m�}��zϡ҅�;7�.�/.���rwr/羠�n��O_�Ei��e@����J�s��;�(qޒu���10�3�=^�>�9�ݝ^*���Ȅ���"z��^z�zz_���=ܑ��D�4�YQU�}uu��-�]�W^����,��nR!��l;�.vy�L�h[u�|�|+������*C�����v7�r��>�=�:���Xh���+*��^%�.�:�s���C�Wx�B����R>�o��T6%`��˜[��X����J�j:v�/t�����^#�)U����.�w���w��9}P��(�|��]���;^*}u��|�_���9p���,e@3ŋ��#t�2�	��Mȱb }C��բ��V�.��y�������X����s �R�N��4G�uo�Jmd�qYm��C,�G{�R�(��lM"�최nC��L�|����\�
W]"��C���t�B�*�5��0Jj�A�:u��P�u��ډ��IU�P������LW�~��҇�C��b��>9Q%G ʦU���eO���;�G�S�-�D��F�'���@��z�������ɖX�K�����ҽK=y��9�\Q�#q2��Ϣ�ۉr��{��s��o�q�����w��><&G�z=Tp׳l^�l���@�<�z�TKf��/��eEs�i�x�+��{�lF�!P1���(
+���+���T%� "�zu���B�Ƣ1upn}M��㹥��n{ol|[�(�&�׹�As�M�~�;~��fe��RCW�:A^SB����>
y1���"3.�c�s�{"�B�n�<2=>V|r�|K�ꌁP�~��u5�7�!�=F2_W���g��k����6�W~V���U�\�m]иM׉�x��� �~����6���}�rIx��vK�Jyw{�G�o+�r�Gj�������m�ѿ����\?_���he�z2�tsi��>������:��T̯Dct����N�آ�����ܼ�x����ޠ=F��^ʻ�_��ed(�ٖ��̜Z���+Ɇ�hd��h�YT�`fid��n;[p��]����,�����v����mK|�5�H�_��|a9�T��8m,�q���6�
���;+�X֗�Kj�d�KT�wso�Nm���W���qW�{�޷�����h�I9���	�ɛ�J�(��a\@��6��:o�+ƣr��⩯q�!��'���_S��sٛQ�g�r�b{#����~�9�:s����'�[�������;q���ѥCȲ��f��po�8���U/du��r#ޚ�K|�i��v��0��3 �&�ᘕ�MX�lH��df+��}|^u�Oݪ�"�5쁎�����ct�{�H^���9p����&|�|��S��9��ւ�C�:�D�&G�/����Mz������-��܅�V8�ޱ*�u�r������>�A��G��RBE4����2Í��q�C+���9^u���q�h�U��IYٞv�uϴ/B3��	+�x	T9%����&r-�37��N}ޑ����}�� �0ܸڜ&Rں��S7�q�G��]�[��3��p����!�>nb����9�h��G]��]I���h��x,z�_���Tg�pv�wl��ڟ��:�2@l�8�)�Q�{�{�.�v�g�|����k�1ם��}�lv�Wq7�\>��E93,�D@j�� pϢ&_�t2��Wq�B%E�f�=�c��Y]����r�`ܸ�Mc�����Q�+�Rch���Ϯ�s/b��m%��;�g�b9�;�1(B��^�Y�Yl�V~.+۾�f)��G�6�nG{�`�Qt���=
`6���yU�
������f��� ��!x�s���k�	�������#�^��>��~t����>��%�Ӏw���Nf}RU�sN=㯱�k=���Y���M3�$q��J��2j2������W�7�z�>������K;*iru�=�>s��!���}����G�X�^�C�kߎ�z^���m�Je�ex�2�~$dI�H=����u��PێT0�����A��Q�Ǥ�8:�ׅ^��Q���u��{��5�]p��t���^vc���7�@������w�a�q�$�a�Z�i��Nt������y��ayh���v��C>J��ȇޠ�>�>5�ډ��Sg��$n�A��9�%�E�e�;{zrI��~%.�f�El��� LEg��3�T�A���ӟyM%;��V��v��܇:N���5��dOm��#<&�4*�����n�n��M�l�q���֮����xo�ｴ���C�Dl�ýS=�=�������}d�@���aʙT+�*�a����gL6V��c}F= W��J�K�]������IAE������L�L\S��-��Y]@ᜫW��>��竵l�F���f�6z�r��YTgS�:�kS6�n���n9��V��&�aȴ|�6\��'rH=�"8�^��y�<8���Y�N�$�3���u�[o)E���o*�ۈ��[%?b坕nB�p	�v��`�Y2��}�*��A6�t�?�ޕ�+��fQ7�{q([�!�ϑ�M0�=�T�9���L^�f�j��xZ�>���_����xno�x���=�>.�C��R��<ITg����0v�(7���{o�4�����O�g�{-�4H�Oף>^�3پ����Bp����gö�R")>z�,7��jڶ�t��>��х��=늷Mb��_{�����H��ݱ^Y���PB@[i�#z��~���5��@Wč3*�S>���b�ߩ��sJD=���.$Ǳn������ޟ�{�E��X�_UT�$�R :%T�>��\j�j�7��ڿ| ���JM�L�}�S���`�^1��+�n�\�.{ƅ��3_d�4}�^\r�}p�*�m�Z�C�n�L6�D/����9����@���+�n�*�OY��k��+٪م������Ja�3^�1����U!C�Pu6�>��������̕a�{�c��zA���3T��|��"�;^�#�{z#���u���}�5O���ߊ��~����5�u���6�?fl�/�i�}A�%vd�-�K�٫���P'*<`t9����\�3P������V���CN�b}��vwRIP���*m�����œ;&�\�q�Ө�7��%uΣJ}Ѧ�Iw�v2�VR0���-�H�t�A|!�k`aJ��&k�]���ap$�+��y$!]��/���j촹&"і)Y����7$ڑUmj�]�	�W*V�+ CKr��Ǌ�@8��sS�� �{����AZ�K�$���p?�9W��%%�:�+#�w
�^�u�'1����%�j[�3Z���U��&�\%p��	�J�\`��B�Bpa��$��ά�
Z�k���T�}�1��L�VzA�(fI���q�����)
f��m!��`�__;�"�0�nuБ�P��G9Z9*5��$�T�u�BaQq��t᎗*�.����+�M�pw5T�p� n�9VU���-�D�lP��Ͳ���P��T�de���z�����v*�BP&�Y��d��۫#��OK;]�k��n�������2*y�j���r�&[;V5E��d�u��9�w)0xm�h��v�j�[4�R�����vfuZJ���W�r��T~���yV�*Gn8nsP�N�]��n��a\ŷM���1���W���/�� �QHJy�(�_%�����dF_1!�[�y����\�8º�1M�̎m���4Mh��Jp��u���"�K�I��z,����u���Y��8�:�s���IX�D��P-�]\y����Ró�7.����l�5x���r�Hj�
��2���,��:<Sh�;�U�Vb	�&�l��i����P��I,�co�ȫN1� :�U�ÝMR��Igt}�q�sfIM�
�v���/F�s~mp��k��y;$��傺��H&��v�)P��m��5����|��0��S)�Y����W��0� �7i*&Ϟ]hvECZj��՜+h܊��n�e������S�}����)s��%Yǯ�x�I�ĺ{sY��2T=&��4rI�N��rd��U�r�wKcC�ɬML�Y.�4fhQt'N�ewK�L��6^6G�Nវ�}��Y�RܷB���K�����7¤xPڹ�ǲ��t���*^)�+0.��5����r[G�-R��ᔨ���av��sl�,n,P�e�@�Ke����7���솵���__hG���ԗg}:��&ʛ�}�NSWHsܥ�(�q��wݕ��ad���7H��n�B7m�Ύ��:����D�1�l�/x������C*�Gت���8���\X����P��K�Ј���`M�(.��fmc�s��1���3�L�#zt�m���n���x1��k��L�S�M��TM�U>e�G��5�D��F-�1h,3)L���)7�]��v���-Ȯ��Uv1ٽ�DQJ�t�	B�P&@d�`P�Y�&A�����!Jd�H�b+�#BRf* �&HІH�#Y"98EQM 4J�҆@� *��&CC�4��J�f!�&K��)M-������CJ��HЦ@"ҙ@���K_�,����6�+#�e۬<�i��)��&�t��3s���c7��6:��]��)�d�1�oV˾�ʥ��<�rRK�O�/��� ��2�Ϋ)
�>�p��W�n_Z
f}�����
HXƠaW�sD^绌��Ǘ��N�t�Ô_�����ʮ7W���\<�T�d]�H޹�Ss;���J�s���L��F{�?�%�ﾋ
�W�஧�t_��yM�`tר��a�%����n�\��w�{��x��u�����\wc����ڲ�}p��P��x�D�|��B����٭���×|Ut(�����k��?_��?S�Y�CݎkQ��y�Ⱥ<I���>>O�+<���]��g��h�T�fB������^��O���T{��z�������,�1�Z�3�Ң�����"L����ۣ<�����sj�x��9��}@{��UF�oE}}��=��#�]���:K��H9���L0$zR7Fx���t��x�;S֯ݻ;;��yޒ�oÎ�ꑞ�u~6�:'�����&@��@��<'~i���yj C��W����-ĽB�{tǏ�߆C���ꃞ��UK7��	P��0�g� ����=��f9?>�IZ51�&B�O�M��j�d�4�s:���~�)�c����Y)�^g�X`�SN�r����vػ�|vo�6Dw���t��&Me��1L�o9�<��B�c���.5�0SUr��!e��9�RѮup4��{�DpݭQ'����Y���aǧ�ώDN���ꌁ_?_�)ɟQ�2CW�	���q�r�Z��g"Vs'��}W�j�g�V�r"��ts�|ǧ�o�����y�zI�>����S�J�ʔ�s���L���KU�������zk��lgͺ�6�|=O��4�40��y�g��]@s�:j�67"���	����vpz�n��(�>����^\4�U��G�ᱪ�(���w�]�J����TADa����]z�6�*^�����ܺ�hbl/�H�;e'�yY�w�R���UxOg߿\L~�5�>9����?��:*$��Q�Nm�`�N�/.���7��@�����c>�N�'��W�5�Ǖ�1�̩��fa�	�*%��l��xu���r9W{4���+�@J�Z\J��@ȇU��{Ճ��Ԇ��R*���ӟ-�Y���Ft�����=1~�U��� 5cj<� o'Kޚ�exyg޻B6�{-��T��<|����|���C���>"��Ji>�������TV9�c���x�
L-����m��Q�KWY`WPS\f�.�-���\�C�8+d�q�y��*��Q�l�	�x�)�4��v��Y[wR�4�Lc����8�F���vѨ]�/�k��-O*��J�]����,+�Y�x���r�SV-���٢�['�nu�K�p41���KuzbQ���r8�i�^�i����_�lv��E����܆v�W��|}�G�Y`���j�sJ�M���7br^���pR�	�t�|�z�=�0��@ʇ�a���S�n	ј�[ mݏ��c����tR�Y��k��V/_�-Z^��������z�鿽wQ5�R��"I�s�d�,a7q���{i��=�J⽂a�F.�\7�ldzg�}�ӣĿzp�U�"��}�xOVxR5SXWR�W�j���}�$�6H�'Ν�/���0�qq�i�z����HG�<7��{B�O�k�6�B9�w��%�y�nRS'�� ��
��oK�_oz��6���ƾ��M�KO�7�[Sk�G��� :����"���N�ldI�8.��¯e�=1��\���W��[��Z�*�?Bn�E��E:6�>�=q�Co�CW��U�}ckC������y_��k,V�yn�ٯ}�C�*�xoܫ�#>}�7�f��+���Sgb<���yc`%c�&�>��͍���w�{;��A���V�'^��ב��qW�o�g���S3����Zg9(M����0�v�]�6���R��8���Wv��k�ν+����SC���b�Ltt�8�F�.�Of�H�_^�ެQ��{
�+-[��1�j����J���/#j���[
e��ח�#�h{�D{��_��r5��ɩ�9��;���3�h�%/���ț��qG�'�� �[�p�x���|�c��A(�gi�͝����}�.�G,�Np�#d��2�ў�W�_D��o�.V�@TB^��n'�	�8�-�8hM/G#ҝF��b�ζJd"�aA<��QNC4�k�s�����}��HJ�{;�/3��w�Ϗ����>��t)��~r��9����t��X��U!��ow�=��vϷwy W���4�W������P��y�{���.e�P<y��4�K���y넧�1���fI�ע��/�Oסx��o�x���'M�_�=�#ܗ{y�������p1p=ޠ(���Mv{�n��2�y߽�F����vz��M�=a^�1?���Z���������K��@�+������~��G�w�f����Z�6�4�xN�qP�n�����UX�[��,\*���G�	����r �Q��CHnOvNM_�� �z��~��gbM�ۨ���=�`�d�H��e�mr�Z�����xM�Y�����g^:��Z3�cM�T��z�[����8Jq���mZ�cm�k��a�I곌B`�*U����W[�/k�C��(�2�߶�5]c9�vԆ�tb�2�,��Q����l�}Ӭ��V ���[^X�3|�ꉌ�yOŋfaMg�y@��fe�;���3���;�5w&.~�/ޟ@�`u�B���6�yP����r�����fT��JZ{��p�5�/ѝ���/UHP��M����;ތ���\�]��HLD�y{�W|��O�pF�9g>��>���{yqGw��q��x��jǫ����Q�3�G-���S°�������Uc�@j�[_�'��d��+Ʒ/��U^�����6��v�����-����[�^���NI�3�Z�iя�73�4��yk9�=���<�ǽ�s�ag\3�~z�Ğ^\@�ʝ?ë����g���Y��,#�F�s��ߩ��ȧ%�h�U����矴�@{��r���^�ⶽ��բ;ڲ֙L�w]�_��4���DWOߩ(Y:�U�x�+�V6h%�;��N?S�Y�W�vC��c�yR:�y�=R'��'@�j�{�[�>�.�.*g��QA;�]�a��z�do�|��o�=����9���~�u�t+<�f�YB���[]Eu:`���1�S�%fG_Rz.e�S���T�3N0�5����o\��|�����7�|���5�k�m�Tz���9\�F8���K9��f�O�8M�&"v�U��o�C���Yo�S,�WD���r�d���{8����َ�}FR7S>�"���Z��9�<����.qOy�"�N�x��RO�=m�.	�|� ���_�L	���Q�+�-{n&�Ӵ=��mk"�Íձ�T&��Ǵ���i뇾�z�ٸ~���_D�0��=��nZz��|��V�X�k�>q�{G{�J�����?N�6�냾��fe� >���l�V1"�H.5:��k�2�F�;6�iz��}E�A�ꌁ_?_�*�u5�6�Hi\�·h�����f�-���y��7|�j�|=Z�Ȋ��]��x�d@���@wD?]�>��wu��d�=���չ~�(wO�]EO��_�}㕓������]�>n��q���Z%]#S�0�kQY���.�z�%X4=����w^��t^�ͪ�����2��x�خ�[�{݉]b`:>�楉돓�ޑ�5�TAF���T�
�+��R��7W��w�{��0��1r"Rq��zk�c�R���UxOdG���Mxώ~rN�����N�������b����ի�/������*,Le�^+=L��1��7�>��R�w,�Ζ<��\���m���%��Wt㛠�=}u�D[�������W�Yk���n%y��K��3�#�Ue���ff���X�T�gu�gtsz�����_!��NG};nb��3Q���^�:�_vCO�B~�g#ޚ�Kʻ{s*C�p�ˈ3/+Sr�~,��풶]������p����H�J��@�U���`�9�u!{��H�u�\w�^n_��$�zǰѕQ��*�o� y_�k�z]_G'Kޚ�exyz�g�{�ό�c,+U����\ï�� �h9�l�SI"�N�����x<���!��"y��ut�m��[hL�����I���нj�K˔	(���C��e)���ԙve����w�s�+0)W�j=;���NG����C=o��݅�x�>�:7I��$)@�|�����Ϗ�īw����>��*�*}^�Ը�;�4��y\�~��d@�����5(U���U8*v�%jv� Qo���>Q��	�@<�!�ӺO�޸:o�n⟌ό�X�*���6�U�,@��@�8z@�%����1vHa?:c��YpΌ'�ޭRc+r1:Gs׹]7�����^��3
+�H|��<}��)��3-��'ָ�;�M_��ޔ��Ch\�,��6�^�g-�7l3���c��C��f,��8]�U�U�Os�ba��̧�����ӿa�}�Py��J?wH�ʚM��]�I�b1�MJ��la��d�˄v�X&I�Eml7,&�'P,��t�C)=�ྣ-�aw�a~���9��y���_$}���`�/��5�v������Ѱkq�Ѵ}h��4���ue�h��~��@��"���H��M��a����Eo�Ҝ���xW��=A��!����WQ�������S�o���u#7�C���U@ه�6�9�<xG�	�~�Q�q���-6&�Ӿ��ڍ˼g�ʼ�1��z���6�v?\W;��3�(.pc_�v;���*/�v�������qWYI�s���1�_E����]`=�u���)����wV�>o�]=�\��qϻ�7��Gz�;�f����ՕZn��*��`	�o��d���2W��O��"h�{S議��'�Z��py�����.ml��s����e�=P��U����y�.�.�ڸ�Ʃv���E�W���R���*��VS��s��
=ζJy%s,d��Tϔ��S�ԇ���Q��M�ʁܶ��=���:���|}E?K�Y^W���j7��/L�� ��>
�E��{��^��}f|�O���Y�������Y4�޿��Ϸ�<z��q���Q�����%��s��P�7=$��Q��5�Mjn��F��tP�����݈H�ʩ2�h�<�XM�݉�����k�ػ$�s�]��;�}����M��7#�m<��6���22�2�<����-M�p�2��Le�zk\��@6�h������t���Ak�L���
�=3�n�X^�o4H��?^�^��=��=�'|�~��}���ɟzt�	���h�v���D�1�.�@���=7��\U�kg'��~�5�nYKE�ċ���T���w~q���� 澒8�n�G⫄�㋺���$w��f�&nm�c�����2��{Z�~�}��URX�RZ���:B�!WR��n@>F�W�A�G��A�Ba5�F�}�6��9�"|G�2Z����h\C��Q�S$542\����ÏJ�m�
�a-�x�z��J�z�M]Ɇߨ�����Q�O�,�Q��6�c��l=>���QS+�Uv����&=y��>+tl���ף�wr�C�P�>���a�E�	��Svꠈ`^�E��V칒�𹆏׋�C�R~C�t�֬�;�R~��S�P��ՏWNÜ�������w�zONo�o�LeȻj�*��Ѹ;�ⲽ���t��W�F����g�r�Q�.'>s�GW>fv���|�W�,�ݚ=윓���-�Ә��ꛙҚE�aM�3� 媞
��z�%�5F�q���f����F��m^Ӛ��@M��T�iN��y;�%)w��_]X�3�}G;�H��k�om�aM)��6�練�H�����}L�{�v���,��f��
�n`��ɻ�J`R��G�QR�&83ɗ�ŧ����++R��]��*�C�ϧ|S�Twd>���N����͉�2��T�۾�oU�^x�fz����ş���=�dT�x��u�~+k�qݑ���1q�{r�% X�#�g;��S����C��g�"��(�P}��xV�)���R�sZ�_��۔{��=D���[��&3l}\����1���:�T�F��w��0�{׃7�>gs}LydEz��{��]�V�&�ު���ට��D�t��C��,T��L庨+U{�|G��ۚ���7��
��iz���^߇�%��@	�}'���A��l�Q�_�[{q>^�yD?�i�����Ԉ������Z<�ë�둷�e��������:Cu���B��C1:�Glf����]��K����ٌ>޷�a�{���z�磌Ɔ�:��mA�� t&;ƺ�:��Nۭ+=SC�WO��¨[�CO��/�����M���6��Q[��+����9�O���=�����@Q�'8��=5=5��$�8]wy�������W��� DW��Q_� Q_�ADEqAR *�� �"����DW�DE���DW��Q_��������
"+����@DW�DE�
"+�@Q_��`(���(�������)��Y2y���9,����������0�� �� �J(P���) 
�JP
 P� PU ��*��IE�)T�JP�
E��TTU*�� ��E$9��"URJ��R��PT*	QT*B�"�R)*%U,؈��`�d�32��`�1��,��Z2�6�h��«X�f($
(�� l(��m��a   n�(  ��  h u�Q(��UR�`��kEQ��T]��*
��ScT(kPU"�S&k *66i�-�P�%Q .�jZ��IR��R�gv�Q
��m����Jc1R+5j�*LL٢��+MZf�J�*�8s�%��RL١���E%� )�*BKeZf��̔�[V��F�*E�-��� \�J��2���dd�*32��MjA��2��U�KQJ��J�A��I�e4�(�*%Q�j�%Jf�R$��+Y�ڙ�T�����Y��kFR�&�E�`��mEJ�IT�G �(L�Q�U��lU)�UR���P�fJ��D��TD�G  v)T�Km R�$�1��C)mb�&k6b��)6�J�QP�p9J'!�FA�--���(�ʦc(���2�TISw��@ M�b�)�� �hd� i���
R��hh�M�h��4�ɓF�� �0F`��T�dCCF@�M44�I & '�h'�i��z����h�$iD0�T��	�14�0� '�+u����ۥe�e�u��Ƿ,3ʱ[L4ө���l"ΐ�"Oʒ�0��N��I\�?J|�j\D�V1~��~2����`j��F*U1�$AQeDj�H�eD^*���
!$A�#��.6َ#��?7.-PD�5rI�E�K�{��,Q��-d����鎋=��,��?����]C��e��S*�xZrZP)�qUrѐ�k�NL7�v0�-X�1lĥDou<�z��\��KMJ1J�'�w�iiuݧû�=�%J�8�&l����fΩ�۫ǻ�T&�L��J��A�s(�1��r��ܷU[���'v1���9��j�i��շ�ST���+1��K�)e�׺�mb�Y��{h�i��n���4�V���-�N� �U���ݭ��I�K�]�`��,��{Tۥ[oh;�7�����e�i��;m���נ�E ��6Pks!�x�<"*�j�j�X�(���ä���B-�M�������,�j-̉�B5iIo&�P7���Hͭ��\ܩ(R�v���Q=�q�d2�y.�U���p��Ybȅ��Y��3r�-I��P�6k$�_Lnݫu.�ZY�aT��l�J���^�6{�4Y;e�^˨�<��H�l�w(�꬙�7�de��[�/s�)[��d;6I��mٛ���5�l�4<U�+ӽ`�n��x��O{��%�q�V�EC*�C�0�(<w�j9��EVQ
��H�T�w�a�%V:q
aU�������Qwk3(�-f]�S\�d����F���:F�]�i"����d�B�h,}�7��p��$��ڙ�N��*��՝I�9R�9[JeV㢍�&�U����*?U#�h:���j�R���0�"�+�R��U������f+��u.�څf��Y�I�Ws#�]G~;i�D��*��%��Yz�E��M
��$*ò�cB�jĕ�P=��Tp��+F٠���v�-yIQ���U��Fi�M��B��5)
��Gc)΢���ޒ+[�!k��GRÇ,awU�r��/S9Vʕ���6�A�ifF�[U�Y�M�J��f�Φ.���s�����Ą�ձiw5<�-��)��I�*֩U�[v��1۩v2f�ʪ����iؓ�P5�jY�gAn�'Z33c��tU�
76���w�>Ux6�<A:��r�9�Qv+V�J���1��n�m&Z��6���w�: M=0��9B��xC�(��I�N�-X��É�.���Ѭ&��qDc?�k͏S��X�w�i�ޔ������
;�9	��8�^n*mŹz�	O*����-]��fm��/N]���3�n��*�TjG3�5˵+hehɚ�I�stfl��o.?�R�!�I
٧J�a&M���h^�:�V�(ΔN�kF�S�nhGt9&���;h[��;�DP�����e�a���L�;��-]� DX���1"yR^�95�ɺ.,�3��9L��8+�L�Q�T�5�e�Rxع��6j[���UJ���1�����[x���h�Zo���z����u(��b�Y��a:Ǳ��*n�f�X�L^%7�j�j�.�)���'��40v�*�u'���%o#�h�t��B,�f��.�̋o/(G(�U`*M�p��o^<L�E�F�㢷/q�
�CՙV՟[w-P�;����ɴf��A����N��иekok���F�9�u�1j<��Qfk���x���)�����#�L;�{���8Yy�5&<Eʳu#Xn�mk�V�V`[z[��kN������k�4ȾJ��Í�->�R�{yg3T��0�ņ�j���2�%eH�&	Vk!tJћ�#ۼ��g]vup�Mڦ~���V3�n����ιV4�2��齰:J�A�.,�T�]��:�9�;z��^֑��X X*R�ԱҮ:����Tuv����9த��Kh丑��o/��UԚS��+��l���q��Z�q|��A���.�:�tR�ݽ5dE��޽0�y_���K�/��*��mݴQ�{��7Ő�=b�#c�YwX7HT��q��r2��Ԫ�eb.����W."d�"m�yX�!���6��
�*�6q���m^L�8�-��L<$a���(����Rwv���j1u�l9k��JV[	�k�8ٙ�f-�pcɴ�:�!wk^����B�R�pV��dڤmL�[�ZrZ��Qժ�X�.�\���I�N�	�JyY�tLWR���զj���E�aN�c+*<{v��Wwb؊���H7Nۂ�kYV�z��P�J��E�їWtV�!�cf�f34T[�ʭP��f��˔�sv����
i'^Z�ۻQf��kD�OR-�wuQ���mz^��t'Y�>��yX��,�=�͜ט�����U[b:�t­8�3yh���z;hs�G�R�&�V軛�rBm�ެA�;��A:@��Um1Iu��ә(+��Sm��G��F庚.�Ó�hj����Y.�B���ãur�W�k�d����E�ı�t.��
��8��&��ۖ�]LF*x�L�Y��^���ୄ�kd�/w3�		�-W���e��d�Е��"��
���;z*�E�wP2�!�5�
a�x�K%�UH�kj�Zz���/0eՑz���w��i�L;�7jJ���a�D����M^ރ@���Vd�l4&�Ш�6���.���K���}OT��m�PEa���wDʱZTv�hP�������t�<vM��P�C(�H�Wn� ��MU�9{���n[ڪ��ҥ��ݣ�����=�ȍ�y�vbbJق�b�
��r��s,���B�ٚ��T0��b�٧��1c�qKXD����T�eY���	ܴ5��w���X�䵔7Z'�7���U�8h;cj���������k*���LK�5U��ږ�<ne�+e�̡����)�daʳA�ձ7$ ��CzM�`Zr�FFBܗ5D�����AD�YN�6mmbm�Tj�ּ8��ͻ����5�Vjj�ҬՋOcb�/]�gq�Ғ�Ӄnݱ�[�͏^@�c.X�4D��jU�w5}���(m�f��Qª�_ؓu70M[�M�K��i���h��v�>���n٢VY�S���ke]���ͽG���Z�w�����R�dVa֜�X���te/���7�Vӧ��+Ԉ%X�p���Vm��d�r�9b�ؤ���4����`��x��?��AM�ϭ����!/\52MU�K/]V�tTo��3�v��ݶ�$2��e�J�uQKS���e��(����7Q޽R��Ǭ3��)�2�/2�ک�m:�J��wl�lRB�J�
ۧ�+,n�Kf�+F%FV��QT�l�ܕz7�j���sv��T�s&�9F���O
�+k4\�x�:�W���Ʀ-�_%FV���\Y�����6p��8*��%GJV�B���#a��{� ad�%3ZU=stK�*za�W,a9r&��8j0t%LY1f�֡�don��WR�jh�Q�f�P�$����a�1:Gy]����U���q�Hu���8Y�M�ِ��)�nn��ʔ��:3 �Fcn�%�mn��/VX��A�2��V(��\	�PD�ni���3V/���	+qÛ���je��0c���^�9�l�DL��*	Gs)��)S[\�#ö��=�F�eG�=E*Z#�4��=c	4��J�A1Ka^[u��B#&�'še��}@�=֒d5C6sp�M˽Z��;�>���k��j��h���ַ�m���$�y"�O<{{��n�fCl�*'t4�:�)d��e!n�^�/oIK!�f���'Xp<�mCf�w5UϬl�xNb�Yv1T!�%U�*�f����K�m��2*q�R��[ܢ�Y�����;��#v����V�]��|��޴����ӡ��|M����[��Y��Wi�$��sH���V^�7DRF]T��x��L�f�n���#�lo�d���!r�T&:����ȏҪ��t3x�-�1�Pk�.dˣ��Q(j�U��Z�n3N��oi�e��[�b�j�D6������.�t$�(��c^Br,��eim�Z��3h��Q'�ja	:
���!�i]�.�u#�I�"�C՚*�ٳ*y\�y�3�{�ozC���O�k?柮��8�%>�J���mp�{��T�L�h݅�������n�4�1��#y�).����AÆ�ܛs0ᤈK�b��[��p�"ۦ�"P*��Cڢua�9yЎ�+�9�5f}:V(	���g"r5[4n�����E�DWN�I�Ь(hw���q�R�&��Z�YF���꺚n2��a0��Zl�f�!�ӻ�]� �/H�F�a�p�q������u�Ǫ-�K%��dT�Jq�W�o]��f���.��F����]>a[UW{z�V�x����������^!Y+#�_[Ue�v�5�vs̛�f���vn�m50]���u�\7�f�+p�ΰ�/�	7	�٭�Q�:�	� [��RD9�����Y-qZ&���8�kV���>u	<�O��ï7M��U��=}y��tJ)d�Y���&V7۩e�쎻,�lu�'f�o�B�D��®iTU�]L�vQlq�[xB�*��n�2��VI�=�Q�V�0�R�� �0oRۈl����!+��f�`�4f�*�'2;��U�:b�m���SkNW��31�!��[S�jⱳ�كMK"k׼P7]XZm�
�sr�C����D8��6�-t��� �����j����t��>p��K;|o�Qk>����\tnF�Let�vgk�Ʈ�Ʈ�3;7Ib�:]h�o%��"�)O�	�5a�r�3�dپ�Nk��f��np�%s\ɴ�MK@)Y��wu}��уV�\a*1�j��qVayJ�ެkJ��D������/y;Y�;�b��wK�&`��bA�c6�F�����j��uz���R��̃B�L7:*E����.ʘB�U��+��Z��bÕ�(�q�ra:��:Y��Ќ*u*�ts8$�n�<t�*�.@��.����I����N������$1�G$Ʊ쵢�gwt� �����ZI��[��5)6���F-�Wv@x�ٱDQ�V�T"�m��.�v+�L�7$]n�[�vA�^�(����PѻP��۶75]�R\֯���\��,�g���眕ʷ�8�<=�K�ge.�}Cm[��J���������C��!��Fa�b橨u^�4`���E��b���g<���+�̖X0��}��.Si�bȅ�ޫ��k�����bt�gm�)CD��TG�M�uL���tU޳+hL�����ed�P	�z���W�F�0yՋ�+����:��ʸ��DnĪ�"נ��8���9�+ϗK_k�O]bx�qR��ҁ���5��&E
����l�T�!���;	Ǉ(+���_�R�N.�:ڕk��Œz�%�ds�h1�gA\��Cґ�
Y�v��{�v}�TW�m;�:�z�������)��m`۪�YL�mtN։Y&�.��	gx`&�M�c�q
�,۬0�����A��v����}�6���T+D���e�{U�Z\��^l�μ�R��*��mb+n���q��+R��:�&��VdMZ�!��z6��Cۺ���ɰ�o�7��y���j|��z�=�nk��6e8s��mf��G8(Gd�G5��u��j�1؟H2d�!˥�pc�w��4�#
B7r�{��6�Cz��oT���j_oڪV>�t'f_G�>$<'e�v�,ꗘY����:W3X��ݩ�g�"�R��`�ec�7H�
���L'M��[�U����N�KPkR+;��/Vq��Kr��<�q�6�U�ݨ2N�Zn�r�9wZ����:7�
Vl�V�;���۬3��8=n豴*�P���e �����t����Ǫ�<�9��wr���,ފV҃{3h�b��pf���e�Ap�%$i���E�.{i�2�~����;����]f���{����$��t(P�(��s�J+�Y��-(} �,����hne\z�jT�Ǻ�;Bs���Kt�} r-3�T�1;ۧq
�2gp]�Q�C���@������U��9��4.[�!ɓ�J��D��yR�J�u���+(�K���5-c� > �t� ڝ�V�u����J�%���iw�	�v�E����{�"�-m-�G�m�s #�
PoM���m"���5YqY�ք쐀���sPї1��j������kG;LD��v��S9��B�N�@`lX7B��ZpJ8��ZA�d���+��Cݯ�D]���f�DL;2����w4ܝeЂ�`��`��8�N�aُ�+�C#Z}0�YK:'� }�Q�ȗyiE��G��uyϳ�v����V�e�i���)!�Q�#79���:���i.Ŭ�+��,�_ذ�ۗ8�A�y˙�I�P>z��]�mv�R�+�&y��bd�>���*���c����n�x��m+tX�t��M买sA��uӒ�jI�.���vm�>z@���K]��դ�+X;}��D�XwUp���W1S^fR��Ȑ&v��z�ҼJj�,CH��xr��֑Oosx(�Y�3V2���z���s��k��N��k�w��U:gL��.��u�@��N=��j	s�Y��5@.M�G\���V6�a�{�iw3���{�m/6{m�D{�t@Ĺ
�IV5@z�m1K�Ι��(i�ᖩ��8kda�^gێ=w��*��bߺ�r������Vԩr�y��N�w]j��u�7gt��+�TcH33Q�����ᕻ��2��e���&�7Q��.S��7�������nH�˩:�HT]�wd��A�$q�/��!�,&�9�TE��J^��w��SN��KM�QQ.�[%��]��+XW>�Ł�37�7}QT3�S���ќ*�蛙mn]���|㺃) �AFz䓛���ƒ�n��g�Ƕ~K�u��)=�-o32�S�����i6��SsWܤ���R�|�+O��2��|dXVX��7Rh���d����f8�(V]]>��#V|�i�y��ggMҳ�<èu�gl&�%m��̭�Dj��������V#u�i�C6Z��^�=��9�
sH�e�;P��.�����������
Z�4)�D����Zɤ93wz���t���$lG����(�L���|B�%^ԃΣ0 �]��κ*U)���[�c��䳛����;�q�f��j"N������V�^&"�ߘ��\����bV�u�y���r\�i�-�����n�n��D�ٶ�ڻg���CiJ�Y��k/-q$�G/qErB;r���\��Q�̈ř��g[3�!��w�nA���i�R��q�c��v�ja�V��T⨸n�M^��s�*c�K(�.�zB�J�xEiv�����ȸktWF��-���H�3\:��J�}ˎ��)䒾��A���:*�
T[ړ"m�Q���b�S\�e*���j��R86;�;d5��_]V�~��f���G:���BK���6�Տ���6��.��Y��v�uXs3C�ӷ��@�[`Ʈ���0͵/y�6��2b�f�n���p��v<�c3���n^f���9�s�<�j�^��$Ю*3��[Dp�%��n�)�tG>��]2Bb���u�����%tju0��	m��AG!&=�iٌ@3�'<��V�$ᷥ�Δ�B7eJ2�J� 9$�$�I$�D�I$�I$�I$�I$�E$�I�Vh��l�r�!9|���[s3�w56F/1�n,�D����2n����Ʈ�.���,���:��-�S��.�TbP��$�a��iW.8㾆��/h�`��SEq5����לpݖFa�ó��9��N�rҷ:�Tu0�aeFfo.�f]�D.�&ӫ�+��ݬR����f�:�e�n���`�����Wq���O�!9�'�Iv�3Q'��䳊����S��C���\�zϤ5=�7J��_q]9�#�gTוɎ�!��Fn�,�gm�u:�d֨P)��n*W6�fF��7o�ٵ.��0�<]�8�J�I�_ܝ��ȑv��8w�7Հ$��//�蔆ۆ��+^ء)Hc7#���>~S~�ٲ�7�݆��"D�+dS/�	"A�-WI��mR�<Q�� ?@���>��?�s�����?/|�~}���ۃ�{���q�^�#���j=�M�;R��aIEӨ5[��x;]��*�켛�}dɣ��"~dQ�����;��{� +����!��1*���F�����h'��r\�<��.Ȇ�b更F��c���1�c��R������t"��a�����a����,�t�1Ջ��8�f�q][��KS�r^�ݏ:�Wf�[ߌː�S�e���b��R��z�:�x�҆b�+���^���T3c(i�J'+�W+2I���L8���0�v�cڤq�S��A�x��!�ty�g�\�0�����)5�$�=:��;U��ތnMX�;��2��_Wc��2���gwQ�)$����2)�����_0eP��y�ri�T�6�m�yHr�é�ÎN�ty,�NV'�^j�a�����W��8T�͵�N��\Շ�G�ѧz��򗙸�F���ɜ4]Z�δ���c���36;ú�b��N)�b}o�\Ƨ݄c*��s.��)1�Du�f�����}W)P���ium*��T�nժ��0������k1�MSt��&���P�R������tԂ�4PyϕS"]�gwr[3�|�WG̬�aK��91a�z����4�~x���-�CH mDl_7u��[��&���i}
uh���X�7Mղhn���ʵ
�S�3r7:YK��\m�s�wS����9���u��_@��@ݍ��7)��aҗ/:�j�׸��{� ����ؼ��\���r��ZdԬ��vP�Q+z�e����f���+7�Avш'U}��䪗���q-�j1�&��4qiÝUq��3VmG�r�I�nlޗ���T۶�K�D"��Aw;�vY�ӫuF�2�YDr=Q��Z�o~շR�l��:qY�uח@�T��$t9��8J���㮵R�;�Z%���A�GݿIwb�dh�����ĻM�c�'\�[kQ�i�p"� �q�K��1Z�,���Vd�yi��ܪ�����Q���Μf�M\�7�8k. V��s0�a4�5���{�wT�a���4k���+��,�z�0�
��]��l��9U�]��wq{�{�,w����,��p6%j��:�elf�Դv�����i(��y/��L4Z��ce���WӔ1��C�Sf�l�$+s�UC*V�:y4�?]�.]-����igۢWA��$��֕����IÅ�B��f���^���;���R�ĉl7�f�0�e�ˀA���+�+D赜�u��L͎�_V[���y��|n���ZCJ�jsu;V��)6a�l�Q��*^�#{��M���.�����j�8�{@ӦX�|I�9��ooj�K$U[�Q�L7liŕ�M���c��]�NĀ�5��Օ0����X
ՙn̉�j�V	k�eqWs���/��-캎� pH�4����d��R&�n���3���Sͽ��8+�3JԲ�nP���F�0S�SZk!m5�<2Q�Ut6��������߫U��'V��%�u��N��GbB��;��U�-�̤am��b�M�Y>���5̾�gˤn�NX�۩n�v,�"%g\�^T��T��w$��&^Ir,=y�"��)�,����Z�S
������6W�d�.�PƟvSҖV��6o��o6���>t�������j�p��"s�)��lA�	$�����6S�XB������L��F[�����/�Ks;hӗ[O�\��QLa�ڹ(�5�t�z�����0��iR��t)k5d�YƂ��n��bKɼ��,�r%\#	Y�vq�a�Q�P��@f�u� h���}��Vu����^S�)1W�%V�+�N5��.N�z�D�dkULjwb�Q���)
ڡG\ӵjmqSS�ܣ�3��VBk��{��]���Q��P�B��5P�0�[Z�9�ۖpè1������2LY�����m�-%�j���u�.T�Vǅё:N����Nە���۝�,ZDc�P.�5�D���bь,e�~�l0��*�@�nVn���$�*��$�e,�VZ�ʷ%��C��.���^)XUL"��vf���Ȥ�؝\V��Eqxx�N��gj��]�p��D��=�	zN�T�Y:��t7�՜��[XE
��sg*����FE�����Y���&KoM5�tN_0�v�f��ʮ[�)�,:k��)g1��Vq�]�����2 �de%�I&r[+/����tp���
(��J̥��<a�ZU�,V�bþ�=yDc۾��V�%b�.d/kv���b���8(!b
xy��pK\_]��!>u#��]���P�>��S�!`��@�@�:.���=��YQ|�T��;Q��
��[�U9�M� I��}��.��+�"�e��nH_8w-92��*n�xX�y�8���m6�Z�ڄ�奋LU���p[�&�E��T�v�%14�y:,N�Y�ՉŇMUf҂!wl�ES�ˡU4k	�1T6Q�ۇa��n͒�obYHt�;'T�m�C͌JT��&��X�X�':��.'q����S"ڙҶ�Wt­�5ZL/����+�����.�*s�w]��⼽�]�S�q0�?�;�{�()96T��[����L˚&:�H��UR��/m���$�pT��v���6!�ޝ��r�R�j��Ţ��u�s�������3َ��ʉ�ΏVL��M�Vm��+[�][�o��f[�WoQ5�O(���-�y��f��Ea^��5�t�r�w
U��+%5w�<ٯ]F�r��ռ��5n3K�ooJ��i]��S�Pi�6�L�v#6�oQ�r�X�WwPuK�o���mv�;U�G��dڃ��״�u�Ei�T"�H�p�t��mdUS��:�Y���������u�l���t�*���/G]+1�d�GP�V1�R-���dt	�f�!	���Gv'��!�ʤ��r��F�>�wM���n9a�J=b_M����K�����mNņg	�C��0f�<��Ȼ�ھ��瓛�z�m.-��T�\{,�tk	DR�0%�F6.�;����Ӹ^)Z���ԑ�|�����}l*O���緉ʪ%ؕ��l�ie6�Bƅ-֞0�^����v�F�a��t��b�.F���u�{�I$�]\�#����oUL�+�L�,E��[y)���º��x��� Nɽ%��f�7ky�%����kK��]c��V2�X�W>��-��v�M>g���=��UH&�S����R�U#HM5�SV��vxt���z������ʅ\l����]"�E*lD;�0��6u�/f�����Iܥ��.�����U�S�Ǯ��ҟ9���"�K*6]VY�kJ3\I{�+X'>9]֚ߐ!��@b5|⃷E�zw�Q�6��k\�> �X7F��c��
XBö�T�/k,�U9H.�]ͫ�N��t�yJ�*���aJ�']i��o7�T����ƣ��|�l;\��M#װ�U۸b���U�f��R��rյ��k�MM즰�ԥ��v͵�st�9�C��)=�K����% ���Sn}�ı"軬����\�,j{%L:��f�[��
�ta̠�.�
y�KD��1���,��+�N�/�HX.��S̜��*}t�]�r��[�M3�W6�C �"����n=���b��Tt�x��D	.�h$+U��$e3�n$�uO����dt�ٓLd!�V
��Z�N�v�U��3��T��)ׂ��w��n.k*��4JK�˫�����xՂ@����ޥNgX�ҡ��$��#q��+kr��n���Ծ��m��r�>�3��8*ie,���mP�� yUpT5f���+J���}
�x�]�o(j�e&,ƨ�yZ�郻�H�F��q,���9�3j����ӻ�� ��j0��/�yw�����ZS4x�Tb�4�o`UC���WUA��ծ�d[���.��Y�^a�o��1����ˏsLV��O� ��XE�	�0t�=�0KW�V�g�_����`���}Z�i�[o_t�r�e&̌l%a���Uܼؖ�}YN>���H�f�d����3:������#cm1���C��{[�XȄ(�ssfaGa�p&
���w]���xxޚ� \��g��sμ�Nw-��n��\��;�	��á�2���7qXS�vfƒ��Gk�4�9����X#�_
.�}4]�=��>���'�'�J��V&m6���)UTV�˶�.�yꔬ�u*9uN�ˮ
�����[t���o��B�|nu�{�d�U&��@�1��p�S9��$�ɶv]ҋq]^:b�rv�4��2�����͛�g�:�8Mq�WJ�d����u�Ɣt%:]\xµ؝��V�N͑9xT�$�{h	��Ͱa�s���r��쭘��e���n���g˅Q�Z�� �j�bȥe��-E�@��PU��b�2�d�a�TX���\5�LYX�ҋ
�D��F.-²���1q�pڸ�\c��s@�����!�\%}J��QVEE��-L��ĭ1ZX��Qdqn�0p��ŕ�e*&\8Z��Qŋ.R�K%F�,��b�qMφ�_�b����nr���M�¥���x:^�omn�GHU	˕�h�Kq}�lY�.�>������r7~W�#.��AJ����%'q!넯e�[��T�;�TNmYZ�����St[��F�UQ�lB��޽�1�=v�L�s�P��v:	wv��j����/EɋY�V�����;��au}�b�@��9��2�/Zr$��wڲ��n{x��s 9��߽A�=^�I��٪��,޳�� �96����կO=�kD�u�S�4���y�{�/֯N;{�i�+ķZ%�O\7zs@�F��/�6�X��,H650�#��7�
�	W�'��������{��ۨQ����;)�GB&i��ui��sm1�B�6�r����Jq$L�ÕŁ,>�u{�VV�i�N���Ѥ�-�؎yA�Kݸ���ƶn�d�G�D���& ���@A���0�)=�9-��'�ktl��js���X�Z=9r��Ok���N�KA�=�Y���|ɮyf��Y�hb�h�+�	���t����i�m{]^�8=f�6�d��hF�W���3�i��;X�-�#�_f���J���m��#���eU���+x3t�w,N/fGM�P����֑��̒�|�`�
O���"|������gf.����7��ƀmɜ%"���0�S�r�6��s9�ލb[g��Өgiת�:��!����sQ���׵f5N6cc�����+�"��ݶYƐ���Kw�:U�9QX�am$e�v��~�{D��hu0i�Ǳ�
��7����.��x�7�,��m���y��ܭ��U��=\Ŏ��m2W(v�c��-N*'���~�|�}{s2-�j������o+*�&�JFCg���K���:)�F���՛pʯb�u@�|�p�L�C�V<�x,w�ؽ���x�[Ma?��#yJA�м;�=��7�P���J5Sj[T�h�[�]vږ����gU�08z���Â�.	2!@3�����X�v6�2�1;�knZR;;,���nh{pi�a�2��إEn�����V��y7f~�zN�c|�RTE�a�tO���9޵���g��������O
]t":�����F��n^դ�ww��T�.�z�َ�%�S��]�H���;��'�2���Ъx��3w���ڸ[�܈��q�Y��=�+s�yH�;�k�a�[ɛ��������	�j��q�4UzЇ�����nf{�'����3��0/^�=9Mީ��Y���D�%�D��*�_9�m|"��yu�wY�[�����l�Bu]p�go)*k-�Ý�_��������s1�����l&I��F}C*.�M}��[�?D*��'%f���t����w�+�����8�wu#�GbPx�Q�V]�~rA��/{:�m�xv�j|�1\����9������׊��yͮ(��Z}(�������)��jU�RZ]L�)�(D�>%��"{*H麄^�"�.*�7ʂ���ͼ)���8ǝ��d<�#PYSՂJ��B�|;ý�AWY�����u�g^�!�n]�rC5V���Z{��K4YN��-+�}!�3�G��_Tז4�,OʶU�b�)ʚʰ5j�Ryf���j�2!pDz��/�x"�F�K[��ɽ��G��9s�Տ��u�����0��	��w�v/�EVRק����s9^[��2���ک�l�9�Q�⧨p�z��I�z{n]M)����ק0F����<G��X��C�Oe=��Sx��u�8��Y�MM>+���9I!=y��L����沆��_<Y�Y3� �Ֆ�b�_:O1��ʯ���{��E��T!v�q�'X���G�na��f1�ӱIR�"4�uַ��.�y.����C0s[��]EEWIG�8fdũ�ѲV����;��N=|O��u/�x������y�Z�Ŧ늊ℛ0���ӧ���w����=Y]�}��s-5W�ff��ܛ�_�����TP�*�Q�ya�湏r��NX�}P��� nTBf���A&�f���{Պ@pW�`����W�J
x$�y\����y����&��v�>E�u�*6�ո�8����跶�ĸ�ǎ�0��T��ކۉ5}��z����ߪ.=�e�V�E-���Zɫ/fM�\�{^x�b6;u�ߧgJ�����}�Y������k���~���Ex�2��z�3�8PC�)*�Y2K��]�L�"�AӶ)궦x_�|.Tr��'��گxlv�*�eQ��*m��v��J��]���_Q|����)#v^�FoU��o+*�5�rNR��'fn����XV�AݬL�;����#CU�--�xc�Y`�1�=�^vȂcd&ZU�Z/,uA�'.���mY����nI���j�YGj�:Xu����k�� V(��������Lm�Bz��7��>;x!�\T��/\�u���E��P�1��C�������JG�'�W�}���m7�u��k�JOI�H�����F�U��b79͞/�͸���d�O�\n����˟3�YT�sK�*>CV��3U�Ia=FN�V��1�rma�<jWW\��Fj�`�����L��95����Q��K£ї|z%�8|}C����ya�o ��� �1�^]������GIma39+_a�T��A.f+�F��+%fC�n�X:h��b����	��TYK�y
8f��/���*���ٽ�ܮ�Et$(������|��Pr^$[��B�xl����2�K�Ec�ש��B� Xˠ����p�XR��g�M�oPj�eWO;���I.�)�!�Y��֫�c1���>R<��N���l���^���W.�$�]�7���쪝���*�wn��&�x�8�S���E�{����k����.B��۲����;�]_�/�?iq�Ѣ�W�;��DC���~��/1C��ҚsOV�}g��(E�v���{y�Yh�I��١������9:��.듥+��r���^}8X1��Â�x�����q ���{
��~������f�*4���z��7�AŨ��UtV%Yi���77ve�ӟ|�ޚ��\<�1�����p{]�}�ձ`D�Ö�A��;�|]�⣛��/j�8���n{����z#�>��O�/!=���S.3FW�vӗ$�c���am�e"U+��|�u�Pi���Ti�	��nm�l�)�����:�;�+������Wiv�V
�k"q_j�$T��Y����Q��D̩��2����`۲huv�0w@�}**�������+��]��Y8���|o��u�sҩ+W��lf��9��l:��ڤ�����J�jSs9��h��E���J�&�s�5ԓ�rV���gmԭ��g�sJ^u��_��b������w�<�烨�Fk��AM������æ�ͧ�#�x���Ʀ�\26Y�@W��8�IL��~Ρ+-&�Cv+�5�ԩ����ʾ*�j�ry��U�w��Fİ��i����.Sr�>��33S��.�JmIX�H��úV�&�JaU����
���5�H��kT��E=Y �Ղ��}6R8����Re�##w�K�_ʿ�2��.{7<7�P-�yWi�,�kE�NnXB��oj��`�]��vL�P`zDz7yp�MVǕ�����<VѬ�g�e&&��i���0����V�,mW_;�i�[��
̈��x�G�����y6i9��en�v��䆩G쩓u$�O8�f�sa������z��x���i&��D��})���0Whȅ��b�$��p��tl�;oU㣖�%��{É�ΘM�a�K���[��v3a�5�r[G(Yߤ��\D�*�V�Cqي�EP��wkecYT�V���󉗭��k�)��I�7-�����қ�jW$9�Lݽԛa_|���{���ց�P�S�+�`8�_VvE()��P���7,�y"��^Ҹ��y��)ؗDa�8��˫��nɤ�ˏ�������M̀��p[Kj��rS.��q� �#��i`�f-�iX�-A6�3���ba���|��QPX�����[3�m1b`��,����Q�J1k�(���1*TV*x��������3kUX��0TUUa�`��A(�A1j"�*�*��G4�"��T��X(�*/���n���i�㭙>�����j���^6nBwoKy.�hWw��L]��35�z�o�omE�ŋ�Qj�aԪ$�Q�3%��u.1�z��V=�Pf$Ao�(�ۍq;����(=�cf��5Kj�7P����XIvp�i�6E��BקK�F5O�/n$ǽ���i�ʷ;7=9�����F�Ki���ے�&T8����캍��y*��ȓ�+��F��us�r�I��O/؅�˶L#�C��$.�̱���UԆ~T�FF��3�r�,\j�K���7��}��kz+�q膪�b��|+r΀��1I�]�s���TZ�����?�8gS�k��@�ob�X��8h�U��vnW��[W+�^ə����#2f��EdW�yh�7�~�˄�Oj�=�?BF��>�y���Ԟ>�Èt�!<"��|O|9+��Tm��܃-M:���Z ����_!nqǖ��;%��)�IӋ��o��e^�������V�SI u�y��UH�%�
�흜��n��6So=�g!HuX>��y}BxlHy�<���x�{�4G��:���pu�4�^�<|��ړ-2��E���mq�O6�s|���	���MіI|FO]9QL�]�"�U*�J��IG��	۝{7DV���H�U�9nP2�����y�o+��Q��+�iӻ�Y�f\�VN��M9c9A܀qXe�&��rC�y?RY[,o{��I��m/���J�U�ĝ��.W��XlG)�rI���ʭ�.�½yu���'��	��ͩ�֌G���eYN�W��V��w)��Z���Y=���\[�S����T���,j��}�*��G��^��1�������Tsw�C7�⥽}Gu��:\�BE��]���P����y4���j�5��cz+�>��=�I��}�Ϸ��ֻ�d�����<x���@0w�	��X|�@>I=`y-�$�L$��i��>��d��{(�����[�,�v��z�#�\$�,CmL�'ߓ}�^g۵<�����a/�e�ߘ4Y}�a�u�����;�N5�p��r�H�o�}_ |�~��C餞�0��d�d�x��i��J�z����!�6��O��ϗ[�=�/!�@�2|��;� if�XM2|�I�ԓ]��N�z��6��C�C�
I�zw�j�w9����J��p��d�!�CL�2u���8�S��!�XBq8�z�$�Ր6�<�$6�������}�ɦI�(I�iBgX,����u���C�<~a�l'����ɤ�I�P��]x}�<��{��+$�=� �I���	�a4��i��=�����{f�'Xd���q	����7�s���sy��3��>Cl��$/{�
I�I>@=I�O�0��=;a�	���W��}�
u�0�9�=��{��=d���C�
d4Πd�VI���'��`|�L�2u>�	�>P�� t�^������;�������+*Մ�8�q�ćXM$�d�i�!��8�9��L�`b�O�e�g�u������w�w^rCl�}��I:��a	��6��8�*y�:�fm���l�d���m�}����k��|�i=r���$�3�HS�Bu'̅d4�RO�;d���`(Lj̤�	��6��7���_;����ﻟI���\��h)�2l��ڽ�B}}����R�U��W�o��{�L�K��}.�#Ja�!�nr�[Z�{lN�EF��E*Yz��ǽ>�ϣ�1���I��%�S��!�&T���!�Co�����2L���t��n����k�@��I9���&�3����NRz��O��2L��{d�5C���:��!�'�6�o.��_{�wZ�u x� i��z��M�wvIԞ:��x���HO�!�a���S'(g�Vj!�z ��K��R�{�J��1���=�0� �����L&�XI��'��i�kvHx!�6���a0�SL�Hu/���̻�}��Cu��:v��8�g�!�&�q�dO��'�&|� q'�8�4�;�Bq!�J�k��q�����rC��d�d����P� q��&��!�M0ה�I�M'|��hY0ya�I�.M9���o>wz��	�<d4ö�z�RORu<7d������d���z�8ï��&�7��N>�����q�����OS���
g��,�@1�I4��J�c�!�c6�m�ͲI��<�!�����~�x��{�u�:|�$��!=p�VNv�Y'P��0H`d�d�P4��m��&�&�qa�'��5�;�X��kN�0:�N�t�$:&�M�y>�0�|�i�{�dn�RO0��I�%L��t��>��W��3�"�:��δ&�ȚY�*�5˙�*�ۍ�À `�xT�`�ݧ)m4�3�Y�DY��9D�c�l���N�m\�f�GZ��w���o�Ʒ���6�m�aԕ�!�iL1퓌�ܶacV
d6��m&9`H��P��@�<����Ww��ݓ�O=N��l��I�<���!�/%JÉ!���$6���8�i ��O;f��s��	��]Ϟ�zߜ$2��&�4�z�/��'������gY�x�$�$�����l���=�s|�����H)0��,�d�=�d�>d�����2�=͒OS�&�i����4�(u�Rq�s�Kn��������s�a�I���L{�%d��M$�`i&_X
�}�!�i�2�3�'�u���~_'ε�;������ ar��C� m'��<d�'9IyI��I��I>`,�$�*g�$su̙�������z��R@�|��	�O���H��l!��P>d�O5@6�ǿRO&������iޝ��s߹׳� ��P:�c7�6�<d4�Y�hORq��{>�6�u��O�m��x�\Đ�����~�c>�����)��s�I�@8���$�a���OXq	���7�8�4�?SL�I3���=t��g߷��^��y���d�|�q�i��y=�>C��d�a��a����!���!�M0�q�;�/jk9q�wYts7ӛ����-=�Ur�����:���9d�Xq�s���� q��uCl�eȢ&�^�w��T��a�ʵŕoD��Z4�]:(��n����,������Ì�����H`4��&`iX�I�O�&�@6�3�@��hy�uƝ�\�:�����H0�N�M$�́ēl'��&M�m�c�bCHL�hi �����,��L��6�m�D�^6�q1s�G���b2}��u���,�N��|3@0ɤ��<��$6�`,�}@��ε�������w���!�s��m�3Cl�d:ΰ8��HhŒ'P�`y>���a3�Hm���@��!�<�7�{����l���	�
���'��Hf��W�&|�����d�	XC!��3:�6�9�㏞����u�@2���XN�m �Rm�L&qBLv�_RM!�!�&Y"�!��2L�����s�_1�w�]�Cl'}�d�)�Iԏ)!�O�6��RO�=J�i���x�>���:��� P��>��w8�~���AOS�C)�>`,8�Xm���B��$�$�&�>`}l6��OS��:��N��7�����yl�!��I�����>|�7��W,�x���q뢫:;�k`��Ϸ#�V��Le3Q���X��k���-��g�����K3��B�8+�5��T���n}�s&�dދ�)f%ԓ�H�V���}�����#��@5x�b��T�5�#EY�Z�1Ug*�V�$����4K�%�f^��DuW{���p��8��cVG�LoE%l�d���A4���Fo���TٷϯT}��������z��U��l��x0�F1�~?����'\=@�J��K��1��f;^�t���c���ˮCk37S`��K|�p��d����)�]��3s����Uhj�w���!���ݾm>95�k-:�p#�:�Y��U�2�$�"���"�ʻn��y����;sjڥβ4Nf�;.���4%�+l�����Nu��)�����-�VC��G��g�٤�1����KO�G~�lh�
�!��IG����t۞9���<�ٗk��CR����WB�Ƨ�5/no�bw��I�7�$f�]��Ȳvz���
gE	�j��4r�v��͉�[�(V��b�Ѯ%�{oo� �5j�6z�O>o���7^�ͽ���΃!~	'�p=׷1�.罼M�^g��x5\�8)4Ji0��+�k=�UՐ�t�Qz�����[�������*���bʑ�G�ߔ+޿oՕ.�'��(g'}\57Uۇ�:�X��J"������2PC~׿�[T�e7��K��r'���q��2��4�lEճ"K$�Kl����D{���ms������%��ڈ�8+Km�S���^Խ����h���!��\	��Y�j�cN�g3��] ��2�YB�t���c������a��{9�d�q��rhM�^�Cw�q+e�����#x���iV���Rj��O�v���b��sh�Y�N�L�-CiJ�rG#���R�Z��F)�n��#Ҍ���y���xn%gw݅��t�%�=����o�����w�t�#M�\�l�/��+�������߾�@����3,��]Q~8z�|�����.f�I�:ܖ�y��7ދ��[9=o��5�¢��e���<[\v��Lͷ�����q��u���f��x��r<�ʭC����{3���!WC�G�E���w7\ɝ���ʮK��$r;u�+�=�ZQR>���3�L�ob=��Uz�si����У�Vm�Ɇ\���Z�ľRwC%J�E܉�t���q�Uh�i΋eM�n���=���Z��g'���\tDqW["�oVT��F���'��F��d�+�2c��2]vUv4��v룎���B7���	t�X�\�:�7����yy�:iӯ�R���+���ՖE^}]Ak"PD5�U�	��\��ӌ�����t���j�6�k��/J�]k����h��eۋy��>�D\�Rz6���Խ����'�������a,D�p���Z�n�	�7��}n'�
2��3����*���p�Q݁�{ݫUi����|�닖ǌ��q���@LuZ`o�nwWy�'r�g��#�n�Z�W�٨�z���ܙِ%����B|;3��4?�����;���,��Ժ�#�ۻ��ӝ@~�Op6-[ْiw�]�8Ą��KO�GV<��y����uf ���߳Q0�^��7/��t�Ƹo�Jɕ��̳v�\���ϥ)�BV��]N.������������e����fj���.L��v��چ���ɱ��!ܶ��v�YQ�}'V�*Aد�'�Y����ͨ�7�G,�ډ�]��ƨ�e�{{�d����5�u�̘�o��P}vJX�n	��P��i�$d��G.NqQA^��� ��!v7[�d؅�Wk��&3t���}���hꠌ(�Dbv�eJ���v�U"Ȫ��ыPDA@	(��1��AU"�DE��1�((�PU�X����b�E���FEY���TE`�ADUD`��)b"(��("Ȋ�TŢ�RC,�b�,��)Qb���TH�'�o������y���n���錾OOU��[S#�XM^��Hى�雽\J�G��De,)��]��N�~�����C����*I�>��_@�Ku��n��^��u�i�<�b�j�]j�A���4҆�(>>��8�7�4�Ú�*G�rWN�Պ�'SYE��k�}��s�D	,K3U����o�/V�*��4�Q9tZ�U�к[M䇰n�7��4&��9�2&GT�2x�4��t*�M��2�v��`Tm0l�{�*�r��aM�"���zL����p�#p���B���R;<�+�{>�MX�g��������.,r�񙃸�6�uV�1uF��b�7uxl_�o�������1��j'�\�bw.��,�Px��oaݤ#s��ﾪ�������+���H/�i�����뇅��TQ�uJ!yҧr#N���Ҋ��3��w�S�+���:�K�t3xV�<S�>Ѡ���I�|;�״�&�����7���nj079�Q.��u<ά�p�n�z�cN �c9�}��~<EE��W�J��/(��wth�Δ�y�8GZ^��cjT�괛,TV�R�r5����.�GB��m��co_X�bϼ��4-��������y�]m��ܝ{I=Y
ѓm�&�9y�4���Ǣ���
�d�����|�yg��.�P���2�^em�k��2��e�ժ	�G�k4����DE���w��<&7���k���M�7H�n�붳��+��!��h��~<�~۳:��b���Nf��%X�Z�+v)ϟ����~I53e��,^�����+:��Qv�"<��
"p�u��]V�<(���8��~^O�'(w���ʮ���T�i�u"�MKS�$�4�y]Z�210c�|�\u�a¹(}d\c=�l�hꋵN}��쬔�k�b���l�ۨ��^�u�"��v3���;w4�.q�6z��Y�s�5
b{-}��e��(�1��
껌��ӮAB�i>�=7�,��U����������(kjJ�{̝�	MH#)�5�_�EJ�gsNN�4�}��UU��&�Z�"�S���dnem��-*�-H<p�*�Yv�Rxc7�����F9#M*·V�Hҕ��B�����{kܠ�'bRcC�J$��^DR���{*G��T(ѥ����w�=b���e���3�����^�p�R;�i�Rۧ�0��&�IK�~>�$N����쪫L�Nw�d4[7�|�vM\�s
{��wX���ϯy7�P���jw���=�_#l�k.�:Ҩ�ov���q�Y%��vz�2�9y{ ɡ���d�H7�b�1��`o�S�>�Kġ���M�`J�v�6����S܎����"�y{38B���^f��l}�{ޏV4�*+�g�ݵ����oJ��]��8����:��YL�Cfp��)��y��ҏm�8��!Ҩ�:^ց~	饚��|r��/Ĉ#��h:��[��P�-�`F������+V`y|�x�C�@{��O���Q��<��Vs0�Ǚ!<�M�΁dr��ImeZ�-5���1`�7�	*>2�"
~�;jnU#;4���5揾(��3��ʴ(��F��%5"��>��o�lv&��M^��ƴ��٭=z�\�E��UNE��{b�z��+8�U���@�7��0��&^d�:���X����f\�7��
�nV�W������G��S�)lM��S��do)�>�^���&��4��>s�>�TjK�~�t�ΜַF@�hc���SZ�@ܙܷ!M�/V��8�V��p[�]ĸ��8:θ�"ᮗD�Տ7���{۞�&���@�Qv�;��-<-�@1m�0#���,�'�N�jd�&� �㫷�z#����2���m]�%���ڎm�����v#zշk$Z�pP���+���ܲ���^>~oT
|���{�j��=���0=z���W�ʆ�U^�U�,�x���;e�| �y�jhQD�����a#]�z�iW�@��rXU��W��{�n��Q����WJO����z=-ޖ����G��4"���o�.�6���}���+�g�g{G#s����yD�gz���%�|O�z*�@���#��_�f�#��Ї��^�ǮpA�ڮd�t_�2��e'�A��5b��؉���^���"p�&��W�̘�I�������SC==��j�nŋ��1��u�*k�k��n�\��Oɰ���
Y���S{I�]l;���[�?>�1��
�Y��V	�v���ּm]�Jbg���uC�4�����H��̾[��Zyԗ���2��k�nU�U�M�.� ���	rTi�L�b��i�"�
�r_z=�y}��y������/��+tb�wt��XO"*��u:���n�9<���fv�t�T����郭�w^��=[�8��(+gҴ��m���r��Z��Mխ��~��@W�.�����6#U
O4�_��U��Q��Z_G�x��4�_���6oY���<�C�g��<�J�����<�W��;Y=��:[��j'��{��A�W�t� /|=�9#�Y�xȻ�>�<p=k���n���M��<�����;�c&�z�:�Y�:�K���X�����l�O)�[(�X��r��ƜY�P�תR[�*��2*�u�z#��EV��C������-פpR���\%���(N.9�J4�4q�쵳�x0 �X��5����ڝ�b1dMt���t��Ii4����a՜TfY��e�fZ�z�-LA{B�Q�{��pH3k�\lT�u�g��Lt��Çf'x�n	����+^�D�βu��;�� ӮC�����r������I�{��4���eޯ��������.�:��wp²&3A��g9��k6qP|u&+���LՊ��,s�1x������k�	����׺�.mԧ��^�)�V��4�,�Lq,|�;нj�h���Z��v���4�"ڱ[�Y�H;�\ ��Wވ��z��m�����I�G=Q����F���6k%�|g�G�j���w�(�X��-�~� ����i#�h\�J�{��s����;�xt�ABR�Crޜ3��6�QȜю{z7�������b>�9�;.j���LY���ɛܯ����W�K��qS190؅P!�@F����;���9*L�B�������5�BO����"u�>#���G���11}W���e��,a�����6U�ߗ��@��C�K16T3��WB����fS�Y+kh����.���h�/���L��F�C(�~N��Β~�W��j5�nئ:�\ﱗ��h�3�L�#��Ω�4�q
T�ڏ~��C�\�hL!S��g�I&n���Шpum�.�՜���e5�6��=�Vvd�Ouu.�e_;�����,���5��1W;�(�}�L�z���]6��8�ںGS�t���R[����6ջ�u`gM��ё0;�<�d�cC����q�7�^����&�i�iV���^���S�|���j'q�$d�{y:�V��{�Q͐W֪^r��^���6q]x�G^x��^��St�� ��]�(�L���rRb������Xe����v������NW�����)ͣz�Ã��gQ�o�jՑ8$�|¦�lB�J����&���&u�=��u��U���n�u�,��͊��*EJê�)�u�o.Jwk�� ��A3�=��j��c�V�v�"�%gQ�{BGq��o%f*�Q0)��˾� K]Fu�����t�TF�pjR�����c编e�T�*(ir貥��۹�����UOޠΛsw�Tz��mm���j��J��؝̹y|�6!���ܢn�r
�O��)��o��E�-��2+C\��+��gS]��L�e�O��gR(��}��ݲY��qwm3b� ne<� �Uj*soh�.�nڦ�QXeu�iۂ
9�x�]�/�q�{��J��Y��ޫ�\��+��I6Udæ�ԋlnf�m�*�t�2�+�펮�v�𻪕�T{�*����L�)a�q�Z��=��ӝ�VH���-�nC��S�x��N7~.#�s��%��m�>�E�Xn�*�M�Xڭ!�776�Чaf-Β�$�L����_v^k�cYE+J��n��aʸ�չ*(��:]3C�����q�)��jdh�ڐQ����U�*u��}�Ϛߗ�����j]�u��<=QBDDd>J��g��b���`��Y���b��ȉ"(�+�E�**ᕂ����J�iX(�)�@PR

�`VQD`�0PAT��0�XCL�* U�"���2ʑ�P��k&RQ� ,P�I��dX�S,��X��`
@Lca�dF�,R
��m�xo��w�߮s|�<NlR��.�S�V$��;�$��ґ+��G�v��9�j�?j5��Q)Q����ȟ��$p�<O6&�$��b�!@�k5��tA������]6��w(v�=�4vz��)i�>~bL/虳[�7/{s��s��j�D�X>yO|���3�+-�q V�i��j}*]�^s�j��kzޟP����>��G�0����ܻ������^��d3v�B�b�x��|�d�kӅ"�r��i߯z�Q�5�������j9��j#&3<�������]ϓ�����psx�BB#Ue�h\���a�2��8��3�1;/�@�T�]/6�����Z*��+��#qsZGxSFg)_�!�Y:\�8���'�.~��FSR�9��<y.��6V��ܪQ��ݬ��a���L:��?xgZ�a��q�F,�ZVʾ�U��*�+��7#y�c.7?U}UQ�-��'�*c��B
T�AU�M�@A�bcI�\�j�$�u�h���0y���ֆ�7��d�_*Xm����3��c�kYQ���6�uq�%��u\("!NȞ�"+���1Ƭ�N�E�>J�z��AK�sZKH4�#fxQ�vӲ�Y���L9�=V#�"����=c�ž"̬�\�������ش�@�|E�H��ǐDO-2�9*�YЉ��u�}�^ͩ�W^�b�^�ڃ&��cј�#!�ى���$z5z�y"̾a�^=�:}�G�o�8���s5oc�M�<]8�#��
b5-�'�Ǧj�8E�)�~�]'���>Hy�~.y��K�)qg�Us��X�n��Q����˷�,:{�vf��^�����6
^	������ȅ�>0){(�&$1�#��b�X��p��A�v�Q1�����T۷-��(��꯫�5�)��b��b���.�e35���*᫊��h�1�m�]��<VS�!T{��B��P.c`m�1�>=SӸ�*a�	�i[}=/�9�"�w�B6j ɨ3M	����N֚mn�h�班 �T�Qi�X]��:p�q���쪋��3= ]=0��t���-Z�	�5JaLdOL��WK^�(�3�1g�`a���ǫϚ<�p�x��>a3�[re{���VG*�oM������d��S�j���gC*{T�(��R� ��C��,$�����Mh� ���[t)�
֚����l�%ȋ����Ԧ�GNnE٘���!�	� �⑤vy����y9t�5�,��~�L��WNO�>�ݑE���Ĝ�tnj���U�A;*��b8�=�ׇ�<�/\�X>cZ�sO]ĩ�9��wH�FG�l�c�HJ�����Ⱥ�I/��DnW�u�{�Y����d�G�㼑�W%V0wNy��;k�qE5u�+�^�	�:
c��kI6x魧�yI{Z�蜞:�[C~�P��C���s��I���1��y�z���ʜzn���$>V]�!����� C2��)r,ݡ����<��Ʋ}3`An��3��HwW|;��=\p��r��R�S�Z��0g ��g�0�(F�e�=�w�;��xS��DU�)N�6zp���:m���Uu-c����a$�hw�Z�g�J����D囬1M����A���_Uot�|--�1�<Gr$2����E�,9�0y9{���AZ���L̏r�1!�̝b;>#��<~c�B%���,�������%)�s�*�Tb�����%^�߼pQ�ٻ	�q���2 ����ι���e�ˌ+g$�T��2�y/�=�j񖳻�	ى�}��x���~_W���N��͹8�,GM��S�=p�K�d {Gh���.���8Yq�;^>��17�f�R�\�,	33�H��lD���ݳ�z�� �^U���N?i41��Ɠ�p"�(����c��6�o�+>׵8]���Db戙S
_�M<�\�$O� ��4�1��<2�5hi�P�����Vn{�Uݪ�Qx�l���Kƈ��<5b�ehs� �e���=�!��FA����3�+-�]�[��dl���ǧ�{Je�9�u�AK�e�T��#��"�F�A�Y���}Ο�!�>�4���(���K!�^�13��*t�u��9d���+��yy��*�OD�u`�W']:q��De�+2�InS)m���>�G��}��y��ޏG��,|�ة�*3�]A�]8�9����f��c`��.h,�"MzF1!�͜H	�����V�9���X��Y���;�eA��Xn�Y��6��L��ua����S�V����{=O�q���)�<�#���mk'K��U��r�� �c���MH�6�J��l%��VIkQ����Ueu�P#���=��deH��UU�Ʀj8{�	f���t�pv��S
�bX�uY�"���d#\��*��zc'']R�UД�DԒ�C��QrV�Uf�wK\1��>8F���׎D�R�]FBq$��޲��I�ٌ�q&vTıo���R���L����z�f�{3���rRހ�i�ǇS��}LM��{L�<�j�R�h;�H��qc�,s0����Q�s^�2�'�k+M��&���ȷ?W�U|�.{�a��o�d��=����5~�ڃ&��cu���q�*iΗ����QA~ʎ�U77���J�Tt�ʏ��Å��i�e]m��i�K���><l�U�%s��Zt���Q����z���V�6Q$_����>4p�9K�?nmt�
s�E�rk��ƋCa�	�.`��s��5��b�����6#d���f�]���H��9������UOHB�Q=��긞e�
zZ\r2�WI��,��pldu�u��U}y��<���xr/���ՆƬ?aͭy]�k�����sg�KL��ßth��R��0�'���
�h�a-3��w��R㧫�CC���Z�s���Yްt�&+�&6B�pl�������DL�x��õ����pj�.�3;ǑӪ��ZͲ�p��b�R[e�'ﾯ��L�ۓa���Lg�N��&�Q��Z�p�{},��g�a!8l��z\i���<�|�lА��-���[�5 �0�6x���a���A���2��6b�y�'rr�޴��Ĉ5�&�E%��d� �y��a,9^¿C�����ŧfT�ر�9��3���RP����I�ɵ��.?$<|xЕ �VFALx�!�M�:ki�C�b=J�'fo��dByB�x�<r�҅���{�'y�]�=F�����׳~�ED�0_����Ij���m��_��"�\�K�垨�Y7@[�1�jf�դNpr�GQ�&o�)�r8������8�`�q+���K�N��f5�Z}N�t�V��I����;ת_��]�N��,o��-aw
�����1ɭp�588�I�������''�����Mu߇�V�Κ"�qu��oN=�m�5�j�z^f�j,�#�y��mi�k��i���1&���K#��ZJ	K�.c� @�BhP�2zWC�~�XsyZs��k5F[ae�׽Qt�wv)=Wv:���;>0��c�����_�g���Ɍ>�q����1��x����� �U*ڬ�=�J@�.d��0�Kޣ*�Ҿ\v�����64����=w���/�@��!�t��q�6���O�oQ��̗~��a��֟J��Fj��	��+S�3�S&i�AYww���ҙ\v��-�:�Q�W��/��|��qO1QE7�(�M`�>(mCc��f���y	Χ��X�)ޝ�;�5�PR��@��7゙�F��<I���Ǵkj�h�r����j���ڛS
�G����\)�E�ңs�_Wխ޴�>���C���/����:��
6z��,z�3{l��M�9��Y��c�
0u��&��@�]9�>]3ݳ�T�f��M�W��8����(��EW�w���uy��Q/�3�3x��~�짴/�E���h�m]����ORZ���c�A`�!��^�3��@y��F�����Z�h4I�N�٤�GlV\t����C/j/r��6�+$٤��(5ǉՇ�^J}��'��	�4�U*������t-U����ۻ*��Ԛ��f9�WO�H�^aK��&å*l��*' ��3fa.��=y�_A#baR����\0g�#�o��Kh�Xw�R�<�=��V-R5�5q�P'�pSͽ�q�ڕ2�6�0l&-��l��_%�p.�c���В��6���߹�#�ˌSm�r��09�B�m�EN�u��;)�/^�V�j�l��l��W0�v!��w�a.v��_XBa�ur���(�O�DI�D��\ ���eN����j�RRh^rbvm"������z��X��nI�'���¹r����pa�U����/�$M��Y�m){Ϋ��J����g�$m{����^�I��aN���E�L��p��ѻE�yr��]�|�ۊ�ޕ
�hȍ�����94�=|L��Yۗ�a��lpNeõ'WDo.峹�1���bA��̀��^���u�˧{��/[����I�=N�s�H�C�s�k��A�㵀rÎ�3o�Sm��5�y�!�6?��ӹq���դ/*��S�Eun��e�[���]E�\��F�=w�|෤G������f75�LƯh�M��Z��e�D��}}t���rg}2}&t�ťk���C��]�[!d��x��ꍙ�En,�����Q]�GY��3*.T�3�n�X���+�ɖ'Y5���:nf�R�CZ6�S:��l;:tZ�$�4|h�ٳ.�7�9���l��1r��w�)V�FZ����Z��u% ���9}�_5�qՍ1>�zL�»m��Hgʅp�n$67gO\�)1�ě�D��ϸ�R�K�n�M�0�٪og�8z�2{����}ot��V�O3 g,�Y�����S�㩆^j��ܑI/u���!�S ���9r��L��Z��Б�u��|=n���� ,TPP�6�p��#�U��V(�"��d�H��T�
a%a"��敐D$T�VR�Ȥ�XE!�¦RUB,p��ɋ`�E�Xe����A((D@2�Q$U��2�Va*EF
�B�(e�R,
�~�^��\��巇�c>{�{X�^�C���x�p�:mu	��E�<����B:�Sd���P����\e��DK�h�J
�B�=t�j�y\��0t�`��i����RJ��*:s*��&��'ML8�(0"�J�=1���Íx�虡Hx��D�εo�{�ez��G���� U�!ڔ�/�r0f����k4QOJ�q������ɡ��rn�WmA��W F�|��Vt��DHj�)�ԋ2��=z������Қ���*�6��i/�9�şi^*2��G�ɇ=w��3�2a�$;����e,: U�W0��}c2z'$˙��Xz/^�ǐ��-2�X��B�ZIv?��Օ֛�Ov�H�/�i�� �Nbf3�}��u
⪤�Ө�8�?Z����p]eU-��*1�W���0�!5�TB�4n�TUۗ��pt��L����^�ܝ�ʫr�jR���1����Ѣ1���������+�)YȰ�������Pt�>B�	Qa!W�q���U�z�#�����t���ӳ�xa��+x7+]V�;�4�9�1
�mLʚ�c��Πv.����^���N�[e��}S<:}$��C0_�2�И�t��¥8�Q+���=���`1D���� �ُ���ĵ�g�⇣ڽ�S3�:Z�4ٳ��`�H�֗z�����N-4G�,B�w���sD�j�.%N�2���������*�}�N���>��� �aFV����5��J�>�Eb�伻h�w.�6���i�&D���!Lo	�AJ�
JI��yw3�aG�Y��n:��j֗*A�ddC��֒U�:o�G�����=y.���'{5`"���g�\�OM���EP�Hm���BlB��o�C�W��g�!�pU�q��#ss-jDJΑtO/��m��T���`؊(��)�x�s���;�:���3�QaÆz�.&�����Hc��U0th(�����MO+��*�G�gW٪!F�zq��C��gx�'կL�yqӚ�kW���4����-#޴��U������bl%�,>�SӦR
Д��1���Ͻ�*G{z�7�nB�'`	� �):�hSQy�g,x1��)̝���i���2gc���Aa�i�I�Gz�ݣ��yM�͆b��6Fw=#	>�Hw#'.�\ܩyԥ�W���Gt�}�T����^k�1X���������u�,]���@��9\� �
*+P���i�B=�<ygc�Qisy�m阴Bv��+d��Ql(gsˎ���Ow��<yh�oh#���n���Y���4ިsv�)%�F�H�u��Ut���Bo1qK�D%��Vtt�:����"U;s"L�
z`�$�ώ��;�A�8�=�p�;�5�ҫ�(�+�����q��v��T�T������V��w|��:�JTG�
�c�Wg����O�һ6D��
��<��L�և��d�3x����z��D�B��0�JZh��xYF�jU,]�]�eW��	��# �5�2mj�o	"'x��h഻�Du�d���.:��)x��h��ں$��QJ�0#f*�`��#B����zg٬Q�V:"�Z�{o�.,
�"Z�Q җB;n�O����ȍ�U�)�Sҕ�K�H���ݭ�&�V$��6r6�ܨ�1��CSں�B���v��ގ4�<��h����J.�&T-ʅ�1���[������ڴs5%XQL��c�DL�6�>iZ�������D���UϚ{�����,^��φN��1;'!TT�S�z��3�����s�����S�Hm�pA���Z��k��]����><'���||x��,45����x�{��k1�k3�l�/>J����_S��x�=��G۝Y�;���͓ڀ�D���=Z�yYEGV�O7�����p2	��O�6G>�ޞ�p]/洖�|q̝�dY��΅�Z�0�U���ǎ��@�|p�L��r�w�����������/�6����J��?W�+{�y�J�'z<9<�Y����Ũvw_�����[e[���sZ��o�,]1��f_0�q鮎������:����+*��wf�,��2��%��ߩU�,�u�M߲�ل-&e1r㩖�ϱ��>2�)niI$(rmMMt�Y����a\��{���[{���2pĿ���>> V��îz}�N���t�m�Vg'�e�PTY$z=.k��1=�MO�TuH��L�)q�gD��5�-2qa�B��Ob*���������uc�E�8�Lq���L�Ƈ��*� ��q���v�kKp�t�O�`�ǎ�6x�ƫ��"�0��Y���\d5�����SE�|���"�v���{����q���=R�x���<�V���a��姓�3a�zdFҟGK0#hf`��[#�%әbc1�����ٍࢍCbMj��e%��!�r�(��g��vj�e�Y���"F��ǐ���gM޼3>�1V����ԇ{�Qqݏkn�j)�Iv���`�u �:;��hw�i�3#a>���N�;\�������Wrb����%����Z1�վgSK!�޽�"��2T��(j�UT<�)�ټ��{X����Z��O����JD��̑3����59e1tN`��2��_�M9�SQb-S�S5�t��)u�T�e���i#BY=*��C�Ηh��c���$��zOy�˕'���<2��9C��!E�<����U��g��
%�({���,����,8x�[���Aq0�������!6`Q��(��2�Ø���"�t�;�I辺��̧�^��X��x�%0��Ͱ�pB�NL�{U=5�@�0g ���k�Β��0��ڋw3H)2��0RZ����ό�bᵵv���gXlgĐ|�r�Zj�V����j[���5�_�V��`�]������˃4��P����2�8j�w�`�6��9�;ƫ7"Ù�R|�{f^������ϩ���Zj�E��s�{.���d�����5ic�A�'�Gr$\P�髍S�W�oz��F�Y�L��o>;�:IY�Hs�ج����v��	���4}v���!��"� �5��c'�M�͊��}U���̃K�{�4ݦG=C���'�B�g�G=U�ۆ4�6���� y��GK��,	3���u�;Q<ҿ[E�|�AU�%*��ƠUt�����+�_����D�Dm,>8o��;V��m�B.n`�5���N�Í�f�6[oG�hPڇj�oENh�'��t�qa�s]�=�,���T��4��f#"'�ܘn�^Q�U3s���}~ze���r��گ�C}�C�����@��f�M�DU��VA��Vˣl�*�k=l ����6+���*�uu�au�ml�)g$�^���SO-�+U#�U�m�;dç��Xy�`�2(��ݝ�=�W1{F~����|=�����2�ʔ�F��Y��գ�z�\�3b��x�	���Xo�|�Y
��*�S�g�֞�������F1����^��1���R;�82j"�e7}7"v�t��F�x�BB:����S�9jg�|�{g1C�|��]6>�f��l�/���1Fkwatܸ��d�ӕ;���Fm��k*�G��xX��|�YX�P"z�:f�^_:+�:Q�Ǐx����`��K��b^5 A��c"��{gْ���1R��8@�O[Z)[���Ռ�����i^�3)�s��X��QQ�^�TɨE�S<+t���y�GH�G�ޞ�WB���5���!�tD�c^\mK����ޠGP�����x*j�N3d�G������u�=�w�w�{W���&�p�T�N煀NH�n��˗��\���D؊��1Q	b����ǎC�!����綛D�/Z�ִp��
��c҉2�a���S5�x{�䮤�L����?`�[����Lٺ�F��+�h�@�oq�P�W�y�������"ym!�H�\���ƲL����8j|���o�8��=c��`�z���z_:��+�^]6��U���T�,�TY$l���2�I��
T<�^���w���3|�f��_#Z���Ň�0�ZI���u�1��{��9:ʸ���}OUji�sr&6]�\ƺP�6�b/�3zY��,������ǎ��x����>�,��V��.�}T�"��#�/>'V�*agN�j����F�OΛ���׬e�R�f��
�CcR�;.Ʀf��Ov����T�����Xa��5�a
��6)/���I� o1�n8n���;���sOk{ݤ�B�(�>�#�/-I]��Մ�\�c2��u����r�k:X$��ŵlLo�}��g;�N����̻|����،�K]:�@ɻE-+ق!.�:�`�#������G���g��A�Ti��\�Z��sR5�a��w^m=e}�^e�ˋ+"x]�q��Sm>έ,Тc������[�V�ݚk�ws7�ݨ�#�VWvgQ��2�N�!kPX��U�����1*2���>a*���Wf�pCZ��F�^L�UU�u�v[�y�q�:4���q�����VᎢ˕��j����m�R�u$�Qg�#�-2�6%��l�ܾ���	o����XĖ��m�Z�R�_F�[��W�v���ez�U�.!�j�7r_]#W�1�V�'x��+�F^"�Kz�I^CXg���rU"-о�W�3�0�*��Ψ�ZWNaH^���H�������܌�\��9�k��s1�f�{���'&f����oU�mꆞ��rWB
[
W�T�nƟ,=���0� �uY��gE#[8{M��[�!B�h^�4��h�Q���en�c�̛heǇ�Kn�)Ͱ�e��ug8Un��}{��YE�.����p��e�HK�|�s5�:��m��MZ�B��L�i���j3S<�έ�Z�>=*�<�v¤ꫦ6V�er�Ms����F�z�u�q �}��:�s�5����k�Q��H�̚�d��h��wa�#��Sw��ڔ�X%>�kr~߾�`
0YE��� T )v�,d"�(ȡ1�%���d%L�� �X�H��P�$����.),*���+�X�5�R���,0�**�,P*Q�Z�Y�&B� T�p"�T-������KnRB(*�C)Y��L�RJ�&�d�E!�����o��ϱϾ�5�Ʒ��=��i�޶k�'�#��TqE�R�K���z�z�c���l�Od��5� �홸M�1�x{F�a���{�a��������a���5J�����C�sٌ��Yޙl�F��K���%�b�6@;��mC�u�x�=�,����D�8tא����,^�LϕF���ՖV�g�.���u�&%N�2����˂�����Te�go��C���miF�'u�3���9�Z�-,�� �Sض�µY:Qd?,<B�d�Gƽ=%�y���֍�=am[$x���cƈ��8��%?`��ٛ�O�C�u<>"�-�QK+$`�.{�l�n�Rz��X�s$C��kN3���@ �� f�<Gd��������Nn�G�|V?���9t�]&�3���9WU�O���7����Ч��ǝ.�V^��o������ҋ3W �$���Ϫ{}��6��?�Gd?�-�}�A�q@F���j�A��i.�ҡr��p�q}Fo&���NoU=4��c��{�wT���x�>#K�ɮ\vSӦ
BȔ�����s]Ѥ���._]y����Ĉ��`@u��geM^Q��\�`�>g;���d�j�C��:p�8�����D��"���ȳ�π�q�r.�a�E��0��'�fg���*�;UR\�2;�z��'��e�4�cر����Xc5���Ò3f�8ǆ���-ޙ+��b�4!�9ʼ�^�s�k�۴�rVЕ֨\����g->lqc��_B���:!ة�n�GP◈�~�Ϧ��欢s��OAb�yW M�@��ƭ���4ygz�q۵���j%,���T:�͊1u������N%^��mC�L���y�+U��)N�Oʧ^��U��,���[��M, go�@�ަ���S&k�@�R�&z%O^Q�LA�t#pd�:Ĺ���Bf��t'g� Xچ���;��C<R�VoYk���!(c�C���!R����A��ķ���<p�x*T�
{D*ꩻʈZA}Qs�U�i�C}u}�uؔ"X�	WK�3�n�����u߄�~(MH ����gޤ#Q�F���[W��cOr�y������l�:��çdN�d�hʡ�F'�b�n��]S*2��K.��S�z��+�����$ekg#`_��{l��M>}Օ6�*�`��E��'�+, ��7U�ݹ�a�&֜�������Nw�"�C|�^�!�Lꮬ�q�?��� R��jҶ�F���#�}��Y�B]}�<�#��l+�����mL��wyl��t�W�4�".��6ꍉ����S*j���VX��AJ��&
T��w{�u$�C�6���#֫��R�/��0��<��*�-]���i}�ؾ���DJ�2��]�%�b2Ȯ]�k&��MV�q�p2#H'	��8E�=�����L��>��ݴ�]�-�>:Eb:�7��<p���,T�u��yמ��p�Bߞ�k����<x����jR��W�x﷊p�^xeW6o-!��ς{w��횒�x��'�h��t�)�T��W�f*#a�D崆X�f|�=�����:�^z���|�̼�a'ťc�'�a�^,�H�ڨj)N����j����33r�nlѢ�#�^����)a�B��,�sg�
�X��]MH�̈́:co�Y�.�� �ib��Zb��ﳙS��׹'M>X�vCgf����9'��D)Oy��{�Q�];\w��я���U���#�����X���4�Z����g�#ߥ�ʩ�y�9s2���
zڸ���}KU)��)r&���9��-]��\�!N�ix��^A�<T\jt�CS�(qw/o�7�:X��K�!y=k��2�)Ḵ���Wg����<��?a�!�5˚b\e��x�<n�Ge���Ӫ�4��|a�&���3X1�+]n2d���+�6&)D��*\�cb�ABg3�dӹ�����g�$y������`S3w��B:�%�/�ׇz���\1<ww���'�F�f$W���Nh\X�O?��y��ۣ���ӌ��/�y}1V<�.TīzQ�B���ƲC��5[�ʗ�]�6�,����8����]�+A�\̠�M�2>��ԯ��/k�V�!��J�Ě|�Z��I;��]�)/�/y�e<����V����+�Z�ɑ51LB��'��t[���Ś��z#K�h��㲙#�mi�����q�Vy��{3�ś$�.8`�<3� C�H�Ac��0ώX=R�������L;�����c�,��q@���r���v�ew�ݟV�G����[�ߵ	帥Ҹ9A��z-��m��+�%�̻?q�b��J��e�Dϕz7�^_�7���q�!�<Q�O;t��,��0�R�����n�?vp�B��`�7
r$A�8�9k�辬Y=}�S���D��{Xt�5ic��Aa�����,[.����Z*�,�w��L�[ӌ��'5a$q�z��+h�9,�5ٵ&J{RR4�cыmZ�ڕr�0�[󜱫�����+͡�<�eB���t�F�0��̱���t��08�ɑ��%����mgL������<h+�;4��x��D��V����#�RU��쉊�X�0�:EL9R�@GI����9\�J�!���7E
p�ٝ�m��N��d͘
y�*^�i�d.��_y�ń]�aڞ��*�2f&T�3b�Z�Yn��}s:&vS����xW�l��l�Q}}�Z�S�E�l����]QLZ>S�	Ɏ�
������3 ���~����~���ֹ��V�]c��_��%F )C=�S�aGMzޘ-xٔ���ڨj쨹]7-����wJ�%�
�k�"BVg�]<=1�|����>�uob�L���.�g����$H�+�c��#x��{��ęz��	9vIBD��dS<J�w�6�DRq/r��Y";^B�Q���U�N�C>d�)0x�d�PGV�br�S[1�ǄV�9���{ݭ�_>�,�?<�����!d���ctb|�P�'E��>��CF���dL�L �Hc��>^�c~N��qy\�G�Σ,k�U��g@�]{�K_4�8N��@˙#��m)v7����0NT�� m�bO���E5D�"|j[~UI�~\x�(�Cup]po��X�L��15l�t\)��mW�}����z�6�<o6i�g[{ș��8m�hW���z���ˑ�5�n�kcz�EG	 ۨsQ"zj��飆ϠoOT�=P����Y3=���G�I�����X�u?6:x��+�෻�q��/ ˌzm�\��ޥ)�~#�p45q����*�(m+ּ�C�`���s��܀�s�W��q�Rϋi��ܼ�+1�ag��p�.i�NJ��stV���3��L#��|�FE��W��O8�^���W��RrD�ed�u�"d��h�+M]]V�,�>ڎ�uc$_�&����?6a��Lw�Z_z��v9J;����p��ħ��Q�pÚ���xv�LŐ�.D���Zgݏ�j�.�l�
�-!�^�5���\��%�&�_�;���<�_��&�z�F�Ce��̼W���{ݮ�̴=�cd�W1�"��j�By�sr& �=�Q:(I����SV'�����G�<i3Q[2��oyO�|�H�kDX\��Xa�T�Ν�?:�/7m�}� �OՅ��>#O�ۗ4��ݧ�:<=0iݕ��꿡��ц_���E&��u�&���5�#�&�Kba�@�S=�8���e5�-WfwZ�"�͡w;����[�9��|�V�b��2D^l�⽩�O<F�b���(���T�>���W���:�Jn8T��@!	�A��� ��e��HB8�;~�{]G��g�v��Ӟ�*cL����ej:y>,��� {�Z�DaS�)�
�0h\^�y�?���O1�ұ�yFL���]����!�S�Ȟ�P����;�R�qDLË2+��ia����w馾���!<���6W�:���	���,{��O��*��v8wW��#�Dޅ��M:7�۔I^Xtͧ�yqiN(TAd��w}��q�T��<w��ڶ�({*}t�3ok'��V0Lt��M�����".����k���a�Ο>�.�&v�g��5Y���d�CY3as�&x�8�Ϋ�X��p��Ś�U1���S���&�$��ٻ�����},�j�ˤeX�;7�{q��9J8�Z��umCm](���ͼ��{n�<��P���Ž�oy�¡���e�U��R��A���	�W}lA�
o��+��+�HV<��BL��f���tr��7�;.%�Hv[�I4��]��r>C7����0������ǂ�t�ub�Nn�ַ6��b����M����E}�Ћ)P�[p��{�j918k��vB��ZHGo-R�����;fC�h���r�F}�:�:ޠo�L��Ⱦ�FA�WSC��
S��o�"뼻���}�~Qۥ��kwvU+4��2�Av�%�W��y1Z��[#�vR���|#Ѕ�������V��������2f�as+w8�#��i�|l^���G_�X�9�J��(g4.Vՙ Ù�r�YkX��pZV���e呮?���\g�r�B�'�g��M'ϩM����.J�Y��NL�X�����c��{,j��L]fU�e��%Զ4�]�-�H)����k�/��8�[�,�[��.t�����
�fi�@�^m��MNk��НXr)bm9]kA�Z�rɠ�ɕdᏍ�&�-6Vc�<��ۺ�ϮB��Zrv.�F�U6ebꕂ>]�
-E"��BZ���:�2�*���.���݃�9�4�v�������ם	�j0*����9<�$ڳ-�ژ���&���Ij����3���B�B1mAX/Wl]+V5Y�JRvU�gi�*x��o�aLq�5�m��-@�n�]�qT�ڏ�w
R,����A�+����*ɕk�imJ7;m����aH�׋�/�]}�]�RAHE�+lX��e��@\2
@PY"�*�
Ab$X�+���,�E"ԨQ*J��
��)}�b1I0�mHV�
I+V�Q�V�E&\8T-,AI*T�ł�I� (B�`�YX�VUXVJ1�E��U����+i#j��E�Q�m��F�++!P����JQT�D�-�!X���*
����(��~�����wTه�բ�c�h�mqiV�2�=6$�d
�M�������c�#�$(��[B��O��zt�P2W�2O9 �9ڜvZ�n|���"�ZD%�?-��14�o;wsh��M,��'��+:5ic��XC��/�j��Y���m	��=:��	�e#}�8ä�Ն�f�s3ٛ����T��G��x�ƈ�!ݏ"� �a�1��i���S�l�0f�WNۯ
6�B���S���n��8!aԈg�`cH���C�=.i�_(�����L���b������9� ���3>s�YI;�]BR�)\�0E��w��ْ��My���f�<pނ��[�O�n[��i�{ez2b�TTk�SHL�O 'E��ɣhz��f�����V�m?��̑�]C���u��DN��ڜ���2CkMI:V}�m�gK�}Y9��%�t)7@�����vsl8����B������ޮ%}�esk5͡S��ߩ���+�7��S<F�KJ97�ھ����(پ��Z��̔�C��A�K�g9���GK�n.w�Q3P�.L�et�����6����_>�b�e+9_�>�i~$0�?1�|Bj�N2{&�*X]�;l��s�!`�e�ه�z`���,�Zz�c"�}���t���z*�7Xy��^�2��;�Q�V���]����"ﴜu6C��(dO�V\v�ʠ�X�"����g���wY�[�r%�.�@��̓]/6����u
��PbV��z(��{w�i�;H�;�8}-�9|�4<��Qk�'J�G1���WK�F��Q5l�tY��n�e�}p�ݜsj����7�w��OwAW�.�;�5�L����z��ܜr�r�����MM&j�k�2�>xch���Hv]�B7?�Fy���s�í��Q8~��a���
}pe��{�;�բݘ�!eEGUE1(;�SQ"zd�d����w�)Iէ^<f4v2����_P��ʎ��
b�I�2�X醛�GYdx�R(��႐�ǥ;|G��t��@�!o
�ے�#ԧ(��ǐV���P����D͏�D4f,��Ҍ�v[vc���d�l	��6au���e{7�0{IB���u����=��@���.S��4�����Ł
ћ��d�@�p�2�XHs��{p����Wۦ����:7�����ƱV�W���ˆ�eK�e����;цp�=��"�ѫ��\*S�ݹ�YsV������T5�YX��*S��if�<��*���r�`�M���G�^چ�!U�uYvˬ�tzN�	*�q�5��6;f�JIhkJ_G��<�g�>����T+���F0�^Q�yNT����9Z1g��T�����o�B�	Q$Uף!����t�C�L/V��>�ߵ�9�~0��ç�0��i�b\��/�&T6z�M��0��[�	�j�ܩ�p�o��CƢ7<j�Y��syxZ�׮�9x�&p��̖5i�;�]Zm_"r���j.�ڋ��eN�MTQ0g��C�&�aϤ\j:��d���K�<�^4�S�!K������/Zy�=�HM�|�;Vo����Ϯ�.T��2'�G"������2�c$ 9}���V��[�'~�t�q�YO1�l�L^	�
�ͱKs��&[�����Sa�T[�.O�[ʤ�z+�e_x�.{1�	MC�VŪ��E�]W|�X��qΙ��
C�f˹Y�VD�VJ���֟��}u�n�l㨯�U|�k_Lw�Q�HE�3;.L�x|E�؅��]-�KTd����s^;�:`��*���Zo�Zjd��c�,�Zu'7AQ(9��ə7[0�7B"0x{�\;^�VsY@���?�>"�\��R��5x�(��VGIZ��+)��0f�+�t�ɯ�q�ON�6�Y�{��֎��f��������tV�Y�H���Š�ҋ�|h:^�7�N{�<�B������2g�6x@��Si"t@B
��\`r�;���9*L�*��I����=w5���v^lۇ�cY=�6�Ρ1�B1��"⁘� �ep��%�{��h�\n�?�h�P�kL���E v�7֮4Ga�2���{�>V����,7�T��ʎ�ͺ���'�η���yV�ϭ��R�]��Y�{(�+�s )5W�ff���U����/?�6�z_L��˿n2c���i���f��jbw���֭=ζv^�ɮ�ꤘ��oUB�#�n�� �^R�xH��[�|�4�e���g�g:�L��)[ �eqڶȣC;��o���~�Q	J��*�z�eغ��e��f����O����oENh����1��b`�_eK����g�̤�_���ڬWc6}kƈ�ٔ��]��p��i:��hsX��{>�V�� 5��k�It�����է9���ɮRѮ����F�ЄF�M!�{���G�?N���Іyq��~UY,��zp��Q����C��(���o3j�Ѻۇ�֯iX(��1�g���򎪏��x662�$NNh������K�RΩ��}���lk:��Y�ەB�fNe>"M���[țf�d��2��{rO�W��I��d��M�TG�6}ª:���+˼��X����E�'�S��]ە�� fbzK���:_m)wxz��+�M=�{�����<��;F�iegP�Dɜ�ڊ�=Y#�ʕ;[�sP]�g.rW�A���-�R�L�@A�bc"�S���>�&��p�s
^�xq�,b�}K�B��YT�͆�� ҭC��Q��qe'W�t���o��)d��28�-d^1Vh�&L�j8�!>:F�^UQ<^o�fu����1E�:z&o�C�iV��������n���ŵ�dÚ��^31l-3�S��_W٬��*y�
��{�y<��7���0�[$o��#`O-�c3Tv��l-P�i����TN���UJFH����L}Ek$��׳c���A��=�fɣ�����KKn� �\��5a���	I���������_Np��ÔEɖ�I�޸����6��5=�+o�'��A���EF*2�� l]J0٦��H��>%-��{��3K�������;�aNp$GA8EʻLol�F�\]/.�E3/���˿�:�����M�JbVi���߰���4�X��8`~a���Դ�S��͟L7dUz��u�n�|"���>x���������1k�D���T���y�}��k� @��?a�!,y�FLJʍ���JeM�0��ΐh@�J�t��tD�I���'
|��=��Y�C�/�.��邁�PR&�i��M�z���L�7�Ö#�lY�G�al?�4��C�g�.�0yS�l��Ń$JӜgh,�K�����D��[�ح�wp:�H���U=���!w�d��8��il>}QQ�K%b�K�G��Dmc��:31rg�}]6�S�O�nkE?0�.:t44�ۼ�u�/�k$C������9�Fb�څ1R��]ӽ���p�}秶�P+�R;V���`^�碈�ڌ��G���U윦)e5�j��G�>d#��F7�z���<vM0����ςK2��OO��*��|�I�r��y淵ʳC�Lc��7�i&LΔz1V:g�# ��CN>2�"~��v��9Z�$ba��cT�Ʌ\��s��沐9L���v/�7����݌�5R��vp�IF*#I������n��������:�;��N�����\����2֢"�+W�%���F.�W�G�=yh��߽y�g
��ab�E��۽�FO5$�%�M��E��r/\�Bw��&�t�ۚ�y�o��G7���H�ktO�~q5k4�3\��^��a_w��÷��1�ۉa%Oi�ʕ��d�y�v:�R#@(.�P˚{s�NƑۓ�"��sq����gq�*ۨfA�]��=yk�1{�"�2��=�w���<�G,�)�pvyaH���ڬ�����}[��ܻ��h�o8ٚu��Q�#EY1�Ms�ʷ�J�&�����;����eҰua/�<���2��mWf���]J��D������t6�]D��O���UF�=1"�5��Y�y�%%9+.k���v;�I��RF�����>H5ʰ�X{�N����*�w��vv,�MD����J��wںfm��T�J;ɝx��p.�m�W��U�g.���Ŏ�WR�-�M�Z���?����`��E����b�5y��T�>�̒6���;h:���c�Dd՚��7t�S��}�&�yr�r��om��V-��f��lE���J7m!�m�}�3{���ӹ���i����g	[�q��ouãy�Ɉ]��J���oM�#��t=wx��8R�w0�]Tһe���,h�W#4�r�|�K�œn������73�Y[CC�K�9>�YUpv"Rw*��}���Y�D�Y���؅V�&��	�e��m�g��n�K��G��WnX̼��	d ��[܇k2J�`;��"��)|���u{(܅\Cz�AR���kF ��4����g�5�Vk�q���x������om3����`N��ofk�b�n��7�h�U۪��+���Z���s�aw����h�VK�����Wd���ˣ�S{Z{��$�.���IVc�
n��8�(b�;���E�֞q�vV�U���:��K-`�&D�T��U� �Ct��(���Yh+ ���n�O�
ci-�{1�t^=�5�_F�NX1+&�ꤧI�p�T���2�]:�;�a��0��Bd�\�E*=���rE.�`H�ff(+eh��K2�QJ�j��ܬz�n�����<���	��`ڍaP����Db�Y��[U�j)DFҒ�B�����X��%
�V�mTm����k0Ő�Z ����Q�X�&1�����P
ʅ-+m+-�>C	�d�e
��Z#��ҪF�b-�APE��VҪT�\ �X��ieh��a0*T���LZ�b�QAlT�*��Ҩ����)YZ�m�*�m(���T�#P���A���m�T(�P��X�"���q@�P��"����$�⒊�Tj
�lrn�����Z���ȶ��.�G�q�u}f>�W�{�����gf�Bۯ,5��e�����([�)�|j#l����MN�k7���sDK����N!Ew� j�{�w7��^���mU(��'�^m���T�Z��{�Z2�;p)np�ίj�p��.3A�3[�d�(
��td#��y���uNZF��1����s�ą�Z��ωW��N8m�����]ڶY�i^�g���5:�*����
��]o���V9:)-Sn�ɋm����I�霶�_����Ƈ�W�9P�E���j���"����\ex7+T�i&�"��64�^��GF�9�v,�he ��JH���a���pr�N}y}��GDŞ�K���2�q�^e�l�Շ�z��E�3q�:1�o'������
��t��z:��C�uj�Qou���J�6;G^����K6y��{
Y��u�%�n��3[��"��OQY\V�τp�����We��������N����⫧��������z���y�0���߽
:�N�@�k�nr�ékk���lZ;�m��M�*��r���.ډ�9���S��i��S��Ʋ��Hz���*�����e�9������"�������q��<ݧ��Kf�s�Fo6e��+{�n,�X4��ki90#k�����w]�Z��E!���8��wX�<;-i�~�O�_W��2�YA��=���h���Zٽ�&��h�R5��.,��6�-N�q;�MqI�])�-���f����Nw}^��·,"=	�)�'~sţ�V��7�+�Z�+YNq��֌�;y=��}&4�ϓ�CѪ�Q�r���ʖUwn>��3��Nl����ܠ��-���g��w�[
]�C�v���V��~	��u^�u��2��u�sR����+{u�f�򁥫���M�=`P�^\\YS���|�#ջ����bw*-Җ��JI�t19��/���cZ�9Vh~&9ǆ����Ti�<�=1�	�r�`�I�4���P/7� ñ��Aؓ��`Y���3z��N>ba�V��0��3ޗp}�~�_�O�5�9ѧ]��"q��j��u���N��x�j�q�w�b�]Y�k�:.2�j;�+N����,`附���%�	�tA�ܙ�{ ��/V��ի��͗���kX�ЅK�r��J���9<s�{ͪKzįSO��m��#k�.�P�⻉gZ���9Kr�xצ_PG�}}��g�wL���Y#H,�ۘ�a �um��\i�O�)jl��e��P��2H9>2�j�R���b��K�_S��q�U"�qv��W�Tr��J��v��jė'jѡ���vI��^Fɞ�Oxo��l�:�Cic����y��K�̽d���-T�����F䛶6t��t�
��<�"������ݜ����杣[�����G#f���'��si1��̭u��������sL	vx�9&:�ځ���+:�j|��yOt����cle����<��u<W�]t}�/~�nU���] �4�m޺��ב��0�:O�~����V:	WW79d!�nXSl�}�^�I����ک�O���_J���h1ò@�Ԍ����LomL3���{��
�+����[K��L��ʎ�9�Z���k�tg� �*�q8��:G�9�Ui�^�d��:�m��*�Yq�Dt��+U_l�׵	=續�/mw���.kk�)S ϔٜv�5�N��+k��B���mǛ�SV@[~�U(�[�7㢗�+��6�[�=u=�����א!Qt��;Xgo
gԴ�����b�1�k���y���k�D�Κ�$<a�~(�{�@�<��YS�����1��h���3Y�3h���EȨvR�ozV]Ɲܤ��yvv_Q�\1�ӵU'���ò�vM�..W!{D�"�"�����Ӗ�n������aҞp�Ν���yt���Ԏ�U^���8@u@��f�O{�%S� ���n5}�g1p�Y��v����
���9�A6L���[5*�����pS�i�E-�m��Fƃ�ʧ��U�ou�Eg@u=UxC�'��Sn��|2�V�!���H��u�m�j���D��S��dD��x�c�wU�Ξz(��͸Űm՛�,̇L	����u��3���q5Gm��
aS���Z�-0d����܌^:�
�8�k��^c4}w�r���D�2�����l�S4H%]]��ު$b�7�)�a�-�7��:�O>tS�2����$̗�l�� �/0{�
��lQKTSZ&8�Kq�����eonׁ��u���|�vՒb�/��������w���i�`���ݍ�oW�b�>���-���ˉ۽:���3����tD���Su�3��Zee�j�����X`�jo�v���u�'���z��SOC3:��2_��f-/��߆R�#��ׄ��ә�+k���^�1�P�%�;��^����y�3�M%Hy�Kj+���uaΕµ��f���]pJ���u�����}��uj�����[
[-]%�[��f�@/nMWs$K-�Kl�\�"�7�yD�ډf:�CO;�Tl��[�su5�����e��GT��:܀R������h�3�g�"꜈i'�]AN6�y>�ة�^|����o�4�+-�<�0":&�F2:��$&�f���Oy2#M!$���Y�B(��(���o,����*1��YU��.�;�X�H.���F����߶}4��s��R���n�%s��K�W�4D� ��ם6ݲ��qo��79Y+.&���8����Ǌ��O�޷Sj��k��L��7�]�]*��z[�:r���f�(QAZlC�R�	kT�6#�[e3`H��1N�����s�I)�lSQVB]�D_gC&�rMtmtoHth���+��R�n�Y�y{�k��+���f?gz�Y9�uG'�8�X;׳��c;�fR#l|z��a�≽k��z��^We7D�N�����t�4'�\缞���H�n��@��ɺ�l�' )պ�I*VGBc�#�~3z��0S]��� ��[�PAj�<D1׮{`iz�T���	�e0f{���D�����P�7�(�!̨�Z;ݸ���I�������Ë���]#G�6k�mB��d�[X�(K:N���܍󒤭��WP�n�H"j�^�P��HMH��)��d�Dr�\��/�ڪs�Ausjsd��zb�R�o�ٜ���s�}����+���Re�L�}�7坃SE�鍻�>�2���Й{\!:�� �RG�h�F2�v�, *��b�FZYD�����g
�ش�9\d����Fk�7(����E:�����n4�[����]ԡ�]��U%�紕к�p��.��Ο0�RY�۳�
�����VZ�.K{����j��n�#v�(ӵ�t�����Y�����ͫ�`WkW�ut�K�$�Wl	���Ǥ�K�O\�E0��P�7J����M��f�Q3(K�2mޜV厳��v9X2�P�9Z����d���{R�-��y��q�`<+8Aʈ�+}6�ZfN��[SBUSzT��çNT�U�a۹�b+�z�������6��}��z��=��ڵ��rl�؎�)����*�Ai=����hyM�*�s�T���Q߉�p=���na�Qe�V�Ï���Fpʾ[N���K�Ѫ���5%ۤu%�݆�n�1Ck��m��Cb�a��RZLj���J��@����ducݦDhvė_p��Ր�l�V����-�a�DS�|��xТ*��n(��sbgl�oQN��������3��^}6�we$Fa���h���"*:;y�� �B�G!Ⱥ��N���֋�39�B����}л���U8���	�ByVzX����ٸj���)�5�6��@[�fȜ̔��õ��C�_�^��ݗ`�&�c�\�I��VgʋR��EQm" ��X(�6����Qc։eDUAA�Jэ�F%e�Rڈ�O�0�EQ��F1UF+%��VVQ0�U+%A��c-��������1EU��E����bb���+,X���T�m(�1�dQ
1EV���F
��qAKDŪ� �	V0͢��	�Q&Q�KEX�(,A#���,X,"�E�|p��Ţyh(��`��0�AC-b��V"E����X��`�[J�1l�L0��@� D
0����M6o�F�,mgn�rͼV3�����t��*٫HF���i�Cz��R,gR�]gy�RNYr�]�1�8�,T����}kEw��-��o;Q;Tt���c�O_5y6�"������jzhb��QOH�9wq^nϬ瞶8��yP��ӍuЫ�HV�r��=+���t���SO���>k�y�0� ��z�43����T�ԩ��<�c���w��X��4(u�
��u/D\xv�����zִR[K=�x�k�&�Z-B{l5��ޢy:>�	��OU�j_Y��a�y*��I]�L{�n�T�Ke��ȱ���.��F@F��{�uv
q�qn^���v�(ȵ�����R��*�qq�.�X��W�F�v�]�jka��67)�Qnv��ő1��w/Wu�]����"\"3�m����#����_����3����w�.Tf�Vbģ0�੫���<�E>#*{m��QռYx9oK�4��[��9N�@mY]d��P�
��aЌ1���Xmq��I�A��_ud,B
՘�J�����.�ޣ[������[�7h"�wƻ�j�?e�aW�������ʫ���;m�on�J�� �����CZ��ƶ�%Ws�L'��Vv�}@Ӈ&��V��jdV�u�P����o��Uq�2��v�����s&H����S���D/�ʲ�6ʼ��
?n쨺�p�+�\k05ي�[��^Ȅ�-q;�EgV��!�F��RI�Pu`���3(ž�O^����Ov��V��O��t�mI1�X��2�ƾ����6��lG�pD�S�l�ۨqB�^��'YQ�=�*�Oʋ��D�:��Q�^�>�9^��1Ed�K�.��P����db�]E٫�Q}g�5���̝5�QO2ޘ�wS��լdb`ĳ��A�P7Ku��޾��zs2�d��Z����m�?Q��,Qtм�����t1hq��3k&K������+-k�{aD[�ɠt1���ii˜$�C�����W�}t�bGc{b�����*��U��8r�z�P
���_x�y*��'�eI�2n�d�WR�
���]��V��؎Rݺ����*Xy�H��Q��ȴ��Fgh�3u��(,�M��Rٺ���Xȍ[^�M#�����zx9�v�>�pz>"�,�@1��4q�et��B6�e���d^>����@]�<7U�G��u˳��PsS�O��h� �ku�iqا�*˽f�oޛ�~8�&��t>����֭���XWU�7nl��\o^b�S���i�d���}�YÂ]eku҇n�]3`[�̾��N�&��V�9�2����1�Rc��	��'�r��ՙ{�F!�GA5Ǵ��]D��Q���e����]3n�A����˼)���,��0iۋ��`_>O��[/xB07��G.������;[O[kS��x�A�ZR�;Y�L�d��5������Y�ܡ���oP�L�,�#h�b�_�C�C�l�d^v�����ʠ=���'�b"P\+�_Ex=���T%z�O%������b�`�*>���\�A�؎r�;�3^yJ��ÒmV�Q�0���}"ߡ�an��7Ob�Oa���xe:�Kh�������X5�Um��u��=�P?y��1����zo}4*k���^)���}\���L�5�Q}�|Ju]�{����UE��8k����KB�q6<�B)�Y���F�2��[l�N.	˔b�:mG��3�)����P��=���$Ͼȥ9V���܇*���kQ�{tWp}+/r9
��4�aʊ6��0W�����U{`��F�,����A�{�ꞏ%
�"o�X���b�!�j�ʒt;�E�Ơ�r�5[G��>��M�]J�A����ƪ�.�}f뛾5����}h׃�J�U�HBov��Y�JHrѭ5:�-��{$#6D�Ӱ	?vͳ�彝�rhVծ<2W�:�Q��%�@��A��#`��w]����o����[�k��lU/N��Q�ܣNnw0g���4�*�Ϸ���D��*^�Kx�ڢ�%iknV`��bP[��Q~
�>��xj��i���M�9��?I5<槗#k�:�K�6�n�����^��cy�f����={��z�δ���q�{�g�{`��u��4n9H/�w����ǚ}IVDt�^�O6�ȼ;u=ɣ2��9NX}A����M����Ӯ�f.b�ך�����J�k����XޓS�������u�E�W.��8[�ڸF,0I�d��oM���*l�NN�qs:]�a�yz(�k�~����G�i���M+�CU�ȋB���Ў��-���]ɵ}ic���n�Z�N�Y����^w�����F&�sS�ْ������s�K��D:t�8{b��ܥ�� �Cޠ}y��*y�=;`{Ti}e��5������ࢧ;i��w�{+;����O��Mۂ�ח��RE�gx�����%;��^J�c#V�A��A��3jGK���<n�
�}��3�d�9jٸ7T��HQݥ2�.j8`��1�+����8�b�k�A��k {Si5V"��E�s�H�z�x���#\�7���pQeT����N}Fyt�%�E
	�Y̏;�6y����^��-CWV�A%�%F�)x?zt��P�m��%�R�Ǜ.����QOb]���-ThƠ,��7���O�/k��{�-��6����;,�b�C"��Uu��\��O'��<l��9^�Y�{�MF�����g�a\���:����F��VV�/�w `�X0�� Ù�v��ɱE-|SZ:`\�*�M�ʐ��k�-t���0:�G\�C7�eVfz
"�T������IY��I��g�wr�p��]*�T:���}���,��qG9NH��p��q�L�htcO�נ� ���-)<K����޿����)_�ۯB\�����E�9�V%�|+�_EaY�'*����f�Ou3M�3��܇� �j�v�W<�;��L�=�8��(3JY�~�{:�͇X�=�3F�"�9V�/��\�}��^u���+!�s �P/����%9M�Z�5���l/Av��2ZnP�U_�f;kCO; N���$�Z[����4���t^����t�(���>��?��̸��%fԩ>�u�V
r���:7�����.q�gei��LQ��*%Y�u=:��+$�c��n�Q���j5���F�Xs�b��!���bOq�{mn�j*�ԺWc��|��Inm�6�t�gf-����xE�ed�m��TJ��U�&�����&���n_2,˵n����͓(�������sIv�q��hjŘm,�ױ�;�mF���h� ��Hk�c�"f���׊х�6��&ʻIT���X{�>��9��-M���p��)VT�$쩊Ғڷ|���'�k�,�1Pל��G)�͋���B�o���'�iTQK�ƞ[y���;�ͨumT�U�5(�ÂJ���)�D�}q�G��H��ǋnbU7�7j�&A+��h��m)Ux�;L*6���&�kX�x��]�|��LriTYj�x�}�kq/\1��m���N��i�?�Vw�)֬רVM�H7+�-�ay��H��E��̛��J�kl�iw 4���eI��X�Q�;f�5Ƶ�)���NVfG�or�nĲ�dt�ΪIbvӛ[@�9iԡ�Ɩ`G;E̬�����QZ�}��c�举�,W;��>�od����zUu5�ԭ��fnfi��'
�,<s�-\ܱ*����ܐܫ�����di�$֝�X�QM+�����)�=:��V3�ڇ �s����v㜊7�n��GU[R񇽔B՗���I������1[2�57h�Ի0)����\�lT/u��)����W��Ǌ]*B\H��gN�%���V�j '�ܸ�\���&��7��;6D�,�Wp_7/�)Vy�4��)�{e��줃��-M���߾����7UYr����
"-[k��ȊT�0�Rٔ`�����֋+���
�`�C�QŦX��k1�R��Y���`ł��R��+��E�VaW��*((��[k��#�5��*��LV�+��J��V�f1���c�U0���B�C�0��S�R�*��&-����"�͖\`¢T0�)m0*8�p��-�.�W�R�=X������ܗ�\87WPT�9/h��i��o4a�QF��*��H�晁�$�ɽ�C�:�l㮃#F����w#���C\��GnE;|����1���7�*��5���܊�N�v�|�$�y
�j��n�W#�I{�N��KF\B�']"=YB#]�k�Uo���{������V��x��:�6�<�e*�|Q+�Z͒�,9�Ѩl��=� �Mk�o��79\������nl�/'�gPN�K5���W9
*h�y��f�RYW2o.⟞SSڳ}^�i;^fB{�r܎v���״�חF�<tg��z
�v���{.oi�a�5s���Ð��Қ��$�f�j�{N�Iξ�Z�7-��(��$)��4;���eG'�"��^�#63�}؈c*�-��7�h�G;=W=����yQ�U��z�{j&1�+F��gE9y�!�p���LvGg9�7��F��+¥V�ג4E7�"p��H�n����.�����Vd�B��s�c�IRmY<N�m[�w�'u���Ȏ����0�n��{W4���,/��N�j�!;v���W���>���z���%�w�Q��X������0y��;c�E.���:���f�F����.�C�7;e���3���-o��D;��=��,x7Exa{{N��k�3V� ЗgW8�5fR5q���[�}�+��Rei��o�(�h�����l;5�����\�Ń�1���j�|��6�m��w�<�o���zi�TA�]͐}��M��m��=U��Ͻ�+���i�s\v�,<<�+Dmmf�r2Qı��9bU�){� �2�na�K�7�Q�a�U��>��mC��Zh�'k���_C�s�ȵ�ESՓ�f.�PWS��n�fWF�2�V�h��o�ǰsyى�w�!�ɱ�M����v�d"Y�=(Ou׋W�o4M�ف���K,�N�zpb�cx�1ǎ��B
���<����9�o^��'vB9� ��.B���.���S�T�r�38�ү`��Rpd�]��)��¶
��\��zi'�>s��LU����ZDv�\W
w��I��g��
����7[E=�2�b�ȍqw�ů�qI��*�67�}J���)��S�+u��n��]<}m��^�h�S8��S(<���w7p�śƖe3{z�h���!�
�z�o�jU}�X��hW�S��G-��9lq� ItУ
df�ޗ��Y][ʰ���5j�[�ז׊ovw���lg�Y]�P�j��7P%�]Va��2�;o�M9��z���U�o-�H�ٿM��3^�[�뽛N�&TR��[���-��3�������n+�I@i%��sq,A:o^v�}�8�^�"��9�Mk=;��^����J�A�����em*(�t�V�o��I����y�7����j�>��tn䁹I�S�<x���:��,15�=�`F^�ݷ7�ѽ���y�V���6=�х��A'J��:7H�P��W}V���d�#��i�t��ѓ�ش-l��1ơ'�2*A�۫��jaD��*�����s�j�C"��U�u�Fs��N���yl��A~�M_W��Җ�\����oV3�u��6(�J�Z�Hټ����q�HuԵ�)=�{�C���
�0�hj�f���]��9���q��f��[�!$�w�f�A��g�{~��J���PD|ݮ�5�+h��=�F�*i�^�s�v�6��CުץP���|T�8�藆�yp�Rr��9~��N����u�Y��X���m"�%Q8"w*u��J�8EgSn�w��*���W���܌����7֌��ZzӞ�_J܃�w��ɮ����9t�cV�7���WҳSK���k��t��T��M�B�;�'[�Y�;�
ǹ��5��K�D㵾�.��C�:	�6oVoQ$*V�A؝�BoW.�F�VW��+�7Z�)&��|�>���7�����-j���ӎ���̵�h������7&ty�Z�=��SxH����!�~���wj�4J9���Џ��)I���,����)�B���.��p=��f�*0ً=�u���`�㏕ݮI-Yu�hN�9i=��;�Ӽ�g���ߩr<8Ȭb5�j��Q]Ǳ�y�U.K��zvn1����D���&��~�"R�γ������/.�[d�zY���#�Ѭ��������qt����@ǖ{ҴAMø����1=��t����t7";V2�.\����x���C}m���y`eZ�Yn�H��]A�����T�g�m_m,�Ij����XB�"�z��kR)9��W1$��jyi��cDNN�c9����,�%Kh�<c98{���&ݚQ0�U���*�,�{�j�Y.��R���V<^�R���.:��N�B��"0���},��v����B�To�V�a�\��왻χ��>Dc�0��~VB�pGA&�OmfW;jN�b���Z�Ӻ��}=�3:��ks�*�I��I	�ݗI���J���=拌�%��(���x��
0Ƣ0WT�F.J��ӛNmp>�E�~����H𾭓��DT�W�e�SҦҹ)ߊ�Z4�����w����h�݃ ���5�a�`� .n�Ԏp
�192���@��V�F9Su�#�9z���7��eSZ���糈�W/nw4TAŕ��Imhu�f�L�5
���3�ΰ���ɼ;���ӷ�X�<I�(*1p��#��My�̯�rC���+�LFM�y��<D�L۰����p��Ȧ�'r�<b�J�S4Ye���+�l�^��1�X�wѮ�W�w�V��uA:J�]���2$�i�z�&�=6�����߸�V�v=��L/Wo�P�R�	���CRN{*�,N�>�n�2c��1e�<�j9iP��r�n^�C@��z,���Q=V�L^�-�}Pz��i���m�\�p����c0J�6����y�8�b9Ɡ3{��M�J��^u��諬�����K@��6��3���{�e��c4��덫��L����}Wj�V-�tAz�%ƥI�>�|�o-��'ot��dmz��f�<�ϩ���9j�h��QR��(�Y^�^q���4^T=���OnϬ{g��iT:d��j���KS���ӽɊ~`,��z�W@��u�W�bx�����$��݋S�~cd���~��������MQl%���H���!������)�*V��UA��[�����"_�MPD�6Z>���2<���/vW/�����
���{�	�x'ic$�E	! 
B@Y		 �$��'�g�y�����b�,ĉ�B�)C��C��e�u�2�b�[e����"%V�Ή���1���a�F�q.hl5�E���I��
/9�ౣf~�3��C�C0h)I��V�'ߝ
��C��9���D�?�5��m��wI��a%$�:�"D�RgH��(����w�/�XtFՎG�'�=�b���sO�v�i�bv��d�gw����G�o�γ�IJPٌ����H�H���S#9rY��]F�1EjG�f+�E�8a���I(ǫ��Nu(�;mz���dS)e깩>,V�$AM�Zk���k��=L?���L�!! �?����M��i1KK�bmY��k�1��i�pd7lOكk�H�t�%*����#��Lx���M���bץJ�<-5&&��Q�n����,C�����}O���?Q��f���h��<��Tּ8�R72w��GHo�ݓ϶�̸Yt�H�������u�ҫ�&$��~��n/�I�e�;�oi�����ک(�9z��=G��ѡ��u)��n����#�I"
)s�H��>���ME1}tNuiUdq\a��%��$�Ȧ�bč�C�7^�FC����(��/.��$���7J��$����i1L�$qr2����2��%������{��B����5L�8�i.U|����HD�5˞g[�ű#���"D�^O�������씟Gߵ>�k_�|X��ޜrGO1�M�,��vR���������G�=����T�>[cH���ւ$A��8c��\Uz�k,���ڍ"��D�-'�/��~��}������i�g.܏G�zћ!���x����*R����c�r�>�Pt���FFn�5�������sK�i����v젉_����a���su���Q����)��n�M�*����6�Ϸ+qъ0�Ǳ1H��TJH��'����(�D���/'	����"$A�'[�8E&I���;����+"�4�s���������*�(�;��:lmD��g?���)���X