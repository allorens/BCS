BZh91AY&SYጳ��߀@q����� ����b@�h   {�_d�6jֵVe
ҚlŶ*j�
diTj�հHM0US!l�D �$����i��KX�U%)��6֒�l�R���E�kM���I���i,�eSj��A[e *�[m��R�PJj��Z�ڂ���ж�[L�U��kT��j��f�ET
���Ԏl�b44�IV�l��I���ZҦZ3Zٵ�Ͷ6&���Z�̫[3ZmhҴ�٘-P�[A��M��[f��V�Ռʙ��s�ĀJ�l�>   7/���5�֧j���[��j�0.��J)��%:��+�
v�v���a��5�k�Z�Wm-:��b��v��UO��fM�)�$jkShچ̔W�   ����A@`�Ҩ���v�: F��@ c(� :1�U(��we ۧ9� t�6]� �Rt�:���H���2E�+L$�R���   ��y�/m0 ��t� P��{ނ�c�����A@6��T s���@t ��y�z  �����P ��{ީ@ 6��KT٭["BH��� ��  �yw� �zyǞ��Cם��f��t�e׽��5��[�� �u\  ':��m�� �ޣt t����Ckd�ْ������ Yx(A�uV����ʩ ܜJ
R�v� 7]h�@Q۱�i@R�� 
m������8 큦������Ji��ٕ6�� �^ :R�NN�t]��wlܠ ���n��9w6�Ӧ]wZ� �;P�t4 nWphPtuY�
 �+D��i�j�f2"R�[x <��n��@� �۵�;� ���4 �w@�9Η
@��ۀ )gkw@
Ԭ  m"�E�*��VTh֪�  �� � ��h m�ᡠ�� ���t��� ���h�8;��P�¨ v�m�6͊�����MM4�/   ^��0 ڕ� (`t˃@�c].vp k�� �軀 �6����Tl�ʶfŠM��   <T��� :\����A��U ��À t۴���\ bh��h >�   JEUA��2�*�� �`#  !��{M�%J��  @ "�����j�  �  ���~%*��       E ��z��L�hM�d��h�ɴ#�z�(��H��O(�~�'���#M9�96�l"V�r�:SkVS�E�����2�ҷm9^jB寮�>K�Y��Te@T��������￳Z�[l���V���Z�m���W�,����� H8��H�:~_ᚧԶ�mm��� ���UV��m��6�6�ֶߏ�_�?���<ڿ�m_9�L�Lֿ|���V�̶��j�-�2��*���j���V�����׹i���׹Z�6�r��V��׹�{�W�Z�-�m�Z�5�sZ�6�sj�5�r��m�r����ֽ�י�{�׹m{��r��V��k��~s^��V��k�5�sm{���m{�׹m|��j��{��sU�V�Z�5^�k�ڽ�|eor��m^���Z��׹Z��ܵ{��sU�W�[{��r��j��kܭm��Z��Ul͵���վ�[V�͵���k[�*������6�����{����V�ͪ�-j�浭�Z��ʵor�k{�Z��խ�U��ʶ��k_yU[ܭkv[Z��j��V��m�os[V�*��ͭ��kU~r�׹[j��իܶ��3U��5�osV�{�mW������󕶷��[{��[ܫm�ͭ��V�ߌ��or���-U�*�ܶگsUU�mmW��U{�[m�jگskj��ososZ�ڽͫܭ{�W�Z�6�r��Z��W�{��r��Z��W�Z�+^���[^�[�ֽ;����{�יZ�+^���V��k�ս�kܯ�Z��k�ֽ͵�r��+^��m�so�7�� �oE�?�K j�36�����^ElLjq���-�N���n�����%U=���j������
�Qj�nq�l���~W���́-��땴n�zKYE�-���F�Ԍ�{�Qz�[�`���6�M��[*��A����"Y�T���t!͔Pa�q�ɩ�d-�5�Kr��Tuzr�����-	E!��Z1V`�e�ӈ����A(3p�4U��R� �,�h����sM�*�4�x���td�jff�`�eIA���ӪZi˫��z���0C��i��P�Y��ķ,�-�IY�cG/���L�o,ЬU��W�d�kJ��Bn�HRC#d��&�J;:�S���ޫ�4i_:K��	iլ��s��jgQ�{A�yf�Q���-��q����]^A5F�M�&/��n1�n8+/1;V9��a�j^�2��y���Z���m<�}��JAH��H p3�B�[
��ȬݰA횔�����/7n��Q�mD�JL���]�\��7��/�:v����]�SA���̊Z�4������V�W�S�c#̕�w���.<�[g*<�,�GS�EZ��Wt��f�/��U�-U�X�-b�G5�����7��R�mtH�QZ�=
�5X�m�\Z_6���}j�o{�ޠ������V����d�8�#�)�Q�Nmm��ߎ �h��;��^%r���t-1�)������mխ�N��-�{w]#nQ��|�ˊ��]k��fn��, ����P˳��E���H`�S4jY��o�tI��˽f$�;�>J�`	����a�b��}[�vЦ�j-X��[ۃ(=��6�P�?f=p�Ʀ.�p˰
��SQ��-}U
BM۰沯E�����Z����	�,��r�\6�nS�ۘ������M,�RZ�)+�Ʋ�,����/��w(+X5i�%�qT����¼٬�60�@�J8lK� ��⹷c�~�,!���F�=�Su���W���1Ób�������M�.��ʛF`�ۨm�R�I�ArF!ڣ�^���+�a���j<���{6���KLGC�5�����m=�B��D�rbЕ��e�dL�*bY#*[�v��tql�E=;g!6)2�Q�R�uX�zw��g�j�b���� +֎Rt)i����&��%8�K�����v�	#S���k7a�e��Cb��֊�% Dsj ��RK6�s�+*J�.��dA7�����4j�bB%�u{��9�X�*n��s3�F��MG ��*Ĳ� Z��#�Mm6"�mɨ�e�^�ٔ$*� �f֛baf����moz�=ʷʛd�CY��B	Cle�ږT�`�v�f��X���%X��Ա&��ݩ�X8��r�=d隠�fl�Ǹ�]�`��J�vp���H5���mf.�K]�7�i���N�Z��L��]@���˸��A�n�<�m�ޡ k\mJ���@n��َ捠cě�KƷVr9/kVu����vRy37tR�:��	+Y��;�����ҵ�1�a�W�j�lU-I��ʃ0����
�Tn�+Q*6nMCz�����Z5��x����z�*��t'yt��x������G��ś;R�A^�8�w����*#]�S�%�v���Y��ݾ���el�����O2-�N����%�6`,aKJyl���*�N�k/�R�n�G����r��9V�����J f���Z�X(-Ƽ1��.��v͗�d�6t1�Ɛ�����Jd��WMf(�Y� @V�tk$Umf�"*�]0�hWc%� �0`]sF��̭���@C�DA��ƽ����'�W-�uy�OB�"�ح̬f¨�hD�Z�hbP�Ѡ( ct�+mԴ��{P��r������uzj7�O��l��'6�DKB��.�A�W���)YVre9Y�Q;�su���t=����5bh���iř��X�@������P�Y�73n�
Qi�+\�)��&e&V����jҘ,f:9.�)�B!�ql�Wh�G]p���ن���f��k+Je��|�В��V���Lnw�&���^3���j�N=S��pM�A�o�c��G6�����7�J�S�H�p=���V�(�q��Q��"t���-�T�5�Q�/*̄ZHVǻ4!{��M�aZ�S)HQ�kq ��j3��aQV
Р,I�X@����ۥ�����ZqM)�T��ikĐN�עi@�oF�n��q��	|�n���ך�s�0ئ�WW����B�*�V�;�y�`Px��Vl Pe��E����n��S��enF���E�_00*��Se�L��2�\���k�[I�1��OR��@���gVS�C��fy��2���i@�F��G���1�"�I�u�n��Zf��7	�\�(�0ͼ*�B��X'B��f=ۻnfMЬ�2�d�¡@[�b���Kj%)�����#�-'�m�b{A��2Lݙ��C����+��������=��\�Lf`-��!n�k/YR��V�
+ZE]O��7��l�i=�11xC�k>ô.Սw���x����e��h� �R�'�a�{�j�Rn�9	�52X�KdWL����)��GKr�aK�_m]!(��Vt2|��J�F àef���(ݭݶ�T�.�s7GcV��m��u Nˬl����n7o�̷¬��BdK?$N52�� ��t�x&�Pp��V���\���
���7�V��I�2�"��`��Y��3\��C/�b���F4�x��ʹ��gH��x��f���!�V'��v����)I�9y{lL���S�'P熺�=?"(,a��=��#�,Q�U�
��Y��cgdڹ�Du����X�k���!�Xlm�8�+ql��o�4�{%�˰�:����)]��$h;�f*��I����pI������f-��0f�J�>N�J�<n�*�Ab��Ʉر7 f���IQb���Fkݶa��P;�N򵌙��TB�٭�^�4�֪e���*juO��U*�^�kZ�mIW�jV�hU��/�x��a�;&�F�<+�z�+ ;#ܺ�@�d-�i/p����Ɗ�*�j0�\;$v�W	�N�Bxq��)%Ag��Qѣ��nڨ]d0% So�Σ\���)�4��Ūz�o������hq��DWc�(�����v��YT�u��Ս��j�U�!Ѱ=�<��ʓ6*15��d�L�5,Åmkb��  ���շQ�:�X�y���aG������'���9eMŢ	��׻W�����%����
j����3rA����[���kD;1|c�.��Su�6�y(�n��{ �A1/�N�uR�;�B&
7�������i�e�o��0@$��B��$��Y�]��Ѽb2��P����8��3&�y	�#w����цn��F�.������ ��P�X��C=N�M�$x���P�8)�7�\�6;٫�E�����ܒ`4�A��k�f��1�ظռ��q���]7�"׵7 ��A�k�a#@f��ɕ��hXhQ��^�r!�!����ta�o��6N�@�5�ս�5�:V�]Cr��QI���a�aT�܄��u�b-j�O��t;6����hk'3p��P$-��^3�6�km�u����S=z��]�e��wF7�p�\�����뒡ѐZ����عn,����Spe�N�h��K8�j�OU7��.�K&�I��̬�6 ��9�bu��AIZ�mTg��]�w)��)ɚ��2�M�wU(��Pr��2^e�D��si>֫d�*�1�Y?1l�ź)�\��A��b3��ÁMy�U�6�l-�f���i$�}z��P�Vf��eI�0��]�V�n�^��cr�!�6Ԓ�:q���Ңuy�#7.Z��҉ƶ���j��V�1Dr��/�.T��`�J�V�X-�����W��<��:�3K�`�"����e��#v�ث:fTz�23r�#�� �u�Fa�֢���nJ���Fn�2U ��j�`�]=Qڼq��H�Yv6�`d
�:��\Wu���v,�ܖ"Ze�#%MyH֖�e��<;�Pv���J
�6�(bHP��'r14]hM^%�BIܭ�v��и�b[o,o��Q̹�H�&���V.X0Q���jí�-e!�@���w.��p?��m:.LK%�j�rּ�ZM�n���E�;."B¹.,ֈ�JF�3��4�ܱ�!ro��e��A�́+܁j�í;r��V٤�P��R��� SC:#*Zv3/m�P����b�ZZz&4��$QV� ǒ<uX��6ݺ���ce���\{ָZ�h�X� �4�����Q�KP�ȹ3��R�f���vn1���&G�GYWf!�!�u��`�fw0H6����Wo^
7�E<�N��WY.��.dF	��#J0�#�oMY/ +0�m��7��Xь��1b%͊��d��Kɡ���/V#*�eZbT�ǈEy�җM�5��X��ܛV�ٔC���֚і�[���2�2��r�g�ջ��y,�e�M{��R	�����My��2��ZjՇn�H0Dl�^��v���wU?E	�L����UB��p��\`��E�gfɘ��[��ʂ\xm���b���w2đb���;�y��%�k01E�Z�<G�(� ���1E�-p�D���U�,;��� dˆk� V^'�b��L��2�el�V�F�ݬ�i���h�T.�U�l�{.��@�0��mㄡ7F�%[����y�!y�ٕj-�0��yz`2`�)m� ,_��1�G8�<5�6x�]1�n��z��^�.�Y���`w�d��CsQ��6L����ГE��D�um�f�^��4���е=ξ�2�+64ag+`Jd��K��}ƆcU��woq��h�N���ph�ԞS�ѹ����ʂIW�M�P �\�2��cS+VF�ӏiͰFYH�����m��27u-�ɢ\h������D4�[�Ҵ�ZW�s�a��X[��3pm[��U���)kɏu���m�b"���%Dpf�PQ�ޜN�6G=�V��Q�MkR��L�PB�s����2��1
������Ʒ��7r��.l�u�Zݘe�
B�X4I55�l�ܬf$�w&E�kw%-�)kW�y����[���b�G���;�U�����M��Y'_�^#	�.n52l�2X�Nh��L��`���2����Z��3,�Xtܚ� m,*i@�1�%[U�����Ir[b�.�r����<T�C"ޚ���f*�&��i��V����s	s2��M[0<�u� Z�6�e@�c͸�7�қOX*+��\�$�
��z�o`;Xr�P�˨�B�ڸ�h���kw5�z��P��2�X{��uv�YM����U�v-S+u�:�Kzp)�Z.���f���Y��{zF�e� �	=����{��Ē��Ձ���Iި��snF�,A��tsnk�cۭ���/�B��&)�NC��VG�4m�"+�[jޒ4'��hhh�L3�[��F��w�7��0� �Wt��M^�f�j�
c5wX��^��߶(��80��fZ�%��"�c�bc8�=/빦���z��aEŨƄ�Ex�G2U��q���4VPN� E����ĬHLL�EC��H���m�krAafiu4Ď���w��h��j���e-�ehJ`ٶ��WNcߖ#i-�l�2i�V��ѶMCkt"AVUƹ�WұUm���fSN�8\��	1<cm,����[���m.���_�PEb������3��$�PPCD�FҊ�L������2��vZš[���
#-��D��ܥ���$4�/vSK@�]6]KV~lV5Cd��yWGcL�ԤÆ��]�K]2�elY�w^��9D�v���onጸ��;$��)��f:�i��ܻ�&,&� (��^���6��nd�J0�D�c�r ulPi��2�(F����e@�qMy�hB��jU��ֵab2�h3�j����Ƌ&X ˹�b�u��%e,ķ	��"ZV��2�;R�ޚ/"Г_m0���������m81�m�Z���z��,,�&��7�i�^�r�$u�����������a,;d��z��me%R�3՗��q'�AYy�b���f$�V�Σ�n;�jl�se��%gv��5�qӧ�mm�@\�sA�n�7*�r�h3.�Y�a�c�+�Y.-뢞k���Ҽ=gF�')�HecL�ZNkF��EI�T ����j����M���j�$�����Dv���I���}��X,'�*���?3���t,�p�1[1mwN�Ү�_Qr�X�m�|6��*V(���ˁ��n�CwVe��Vi"F%;�=o��l:{L[4r��;V����b�"�х���c���m��K7�1#�|-S��f�m�bв�ƙAՈA�:&\�;���b��+t-7�T�F�2��`��U�� ¬����6��؅]"wi�1.n�ܲ�֠��G,n:��*���}KN�$���1��L��t�{�Z��Xd���jt[{THK!?]���T�ZԨfhaX�����P�1�1k&��xL����;|���pp�K�"ƻ���v΍"�]��t�i�@�n�W�W6���]�`�Xxh�6Y��K2�-�Z�,tVl7]�<��� ���H��[͈2��p��Q;5Wc�#ݼ��S���v�a�)�yn 4��f���fqz�]0t`ȞY42�	˽���k�u�+#�K�=�;m־\�Z&��s[���-]��\=p�x�%�&��,�j������a+2���4��Ӳ��b����ת�N�0Ʊ��+����偽����6�>��|�z�'�~��@�C�����ڲy�n{��zk�T��F�����y1�Ԗ8J�.��q�jM�z1
��<x�l[��Q���5)7��m��7E[�v'=�ԭ��iX��{�&��F�v��c�U��r��N�SF�s�J:�u��R[�U꼇̰���q�,PU}>��ҭ.lW}-���;���n[�p^��	\@q^B%+��di��ǋ�n�7b�V�B!7gd����XX�b.��r�N��-̕���qy�k�yd�D�O}�.�*�骅���v�&9�++��4+nZ��s(��Fp66V>�ܖc�o��aw<�qv	f���5*3����[����:�lb̙u�e���˜�f�/{7
f�JQ��kE�f��azH�T��ԉ\���V� �զM�c5c��5�����ږFk��!��ҢQ#��+�U�*b�����9���P9�:7-�Lx���{��Еh�h�x�c@��ެ脾�c��vf����H��`��NW[�N�;]�qaVc��Ь�K�+����#�1�T������N�yG����6�.X��*>�D	�!�Z�^�9����پ�l֣f�ډ�F���G@�|���+�9�ceve�y��,�ٜ�M+6M5�A'�Vo[.B]k��eIؚ�����G����)�XA���f��G5ӂ�)��P>���<�2Pe�]�]���'���O 9��:�=�mr�5N�$*&��Eern�U>��(���1[�w�w�]��:���Ȱ�S7�:T,�]\�����!����ƱJ�6$���7����BoGz�p�u���V�rч�,�v���*hKk!�;T���/I��5��� ��^���^�t�T�6�u��|#*����!C',�2�/>9��[\���T�b�|[�A�����h���v_�^����(��r&f��Aǳ��(��'9���t�r�v�'b�#@�L�%[���~a����fR�S���!��)b���O:'���^
h���
�9���-�}��x3qS!�f��*���;1���m_-擬q+�E}q���+l��B�(���=�敆 �4#`�fI����]-����7��/m���S���5؊N�����-�le��7���;M��&�t�ׂ���:̻���j�M@�iG9L�ׇK�ǖ�h�]Ä���`�+��brS�d���vƿ�&>���<jrf�WỴ���l�<Qm��OT���)��]�ɺU�^�Ad0��:��/����$A�A��cj�JS4�l3mM9)T,����F���vѤW=Zz}�L��&�Iyxl�.�̺�4W3���WFփ��#�-̓��a�RL$f�Å��)�e�����;�j$���֋A�;;���]�t,rD�h�z��u�N��	E�q^n�Xj����3�qES�n�~W�LrV ى�n+�VM��

�oU���o�u�<%	ڎdХr���T9�=���,�I:q;�v٦^�G�"'o���ΐ���yp6��ʄ�0뫨`J��7��������2}�U::۱⽘!8�*WN�q��D�H� .�e(�*[�3QC�CV��Xq��(�"1c|r�5��N�Ŵ���b��;j�GK��<��b��ڨԢݼ$�Jf�zuqhRR�÷���:`�K�飛)^.1v^�RaHwr�k	��o��^m��Xm�p*���ۗ����u��7;U�f�������ź�Xm��-O*h2�W]�����#�"��j�0�B�1VR��7OA+����=��x�Hi�Nvg#S���5&���=�з��k��ͭ����}S�d�T�S�g�uQ:��\�� *��{}(b<L������b�c�A-!e�c��Q�&"�W7��R�"V)`j� �ܲ.T�;Ha�̹i ��f���D*R��
�ú�rQ�ʱ6�������"x8����z����Yv��G�7�n"� qws��uqM�e���bq�85����i�7]�6X�zؙAgv�;�Z��Ю54�q�7��:�{�M�^���ka�2�.�ɪ�v���2��cڅ ���e���WP�Z��G�f�>]!�qi.Zk�Lr�R��y�r�ⰲM�Kl�j�XfV�(������,�Z)��"����|M�p�U1��j�˶�E]&h�B����Of�l��;�����2W%Q��,	Z�,�m�EG����v�$R���r�q�N-̷�ҵgCwd*�{�I����:e�z#�I7Fmn��y�l!r��Уƽ���w�����)�f��$Sa�jxvZf�x��ػ�m�Ȏ�;�.����5,�k�Vu ŠZ�q��(�a�����fYjw�L����J�*�9��]p/s��w������y��I9�����Ӎ�7=<�����.Y��9\�)h1��.��e]c��1��ک%傶uoF�10V�
�k�\\��Б��c���d1q����M�d#:bٖ�6E�IM`�L���O�!�8K�.�o�+�:"�d��kB���nh5q<��L�6�%]��m�*��M�8������}YW$��{s
��[_2y%��r*���5���N(�+y��LE��Aqf�Z�bޝ�2ڝvAK�ؖ5G:�b�L�n���%,�qn�⻿�J����h*	^2�VZK#�`���� ��V�A�o��
j�W"�O0@ɧ�6*\��茭/��&[��&4���I%��^;�n(�f4�^h^%�-�R�������ۗ6��@�qp�֤�۩b�a���}/��Vse[����H�]��gk��:<3���w8�wj��I
���-�����$�at�Ÿ��5�3rmg4�&�*Y��7�ɤ���MtAd�l��2�W���V#(v�M����[��䙶w�!�6�l=A���gP�4rt�7Ӷ��3^���:5����qIB�<�^Onb�Yϯ�K]�+M��5��כ�V�U�.�dL��6<.�ִk+��@V=�"����\]��2�G��^(���_x����;���'S ��uu]Y��J�j�XkT&6[��R�v��k���}������.9�V�n��E5�9�������6}բ�2�J�umr�]�/h���N�Jb���r�c��U0�(���ۧ��!��1��n��-��<���&�{X�y)\������	��q<�i�̅3kB�ڽ1���
5�RWXd@T��Ihe���hh�5�mm��eт��ˠK
����f�f�s��o;劈���\77�BmX�+k��Σ-Hlݦ��[.a�e�ն��Ž�o�����Ƒ6r�x��c�����m��nwK��0ݍy�uLZi]���uiK;�)��[���8�{]����m���3�z�<��.r�mZ�W.�i��ٚc�Q�t���i�@���+�
��˩�v��i.��v�;ة�6Yx���Lǌ�͸��kހַOQV���T�;nV�u�ph���4�in��V��64f�f�@S��a�+6�*')GV[�D�.�r�B1�c�]>	rgDF��y7�!׵��_S�8̅��Ed�,,���2����[\�g{ �i+#pk��\�D���m�>���|���.HV�b|1��fe��%���`���.�u
�b�d�j��ySl�o�Ā�<����(ְ�t�ڷ��J��K0 ���v�s�]N�մ�.��$�e����H�S:��Vs� ��j
qd�%��F��/�_Vp���{,<C���N�����:r��	� ��2�U��|Q�4#��

	�������M�]\����o����x2���2zK�Ue�7�Ƀ��B����D��.J���\��6�;å���6�.�\��u��1]��T����&V�jB��+ǎ^�A7#��a�	�ں�8{��n'
q�S��D?�����s���ڏ.��s]��!�!�r[�$��A"���Y�ݏ����oh�
��p���|������݊]�˝1��o-��u�΂��2Ԃ�V�3��%�O�nT{��g/��Iˠ{�|颳xÜa;�#�m��I�9��t�6n��&�sOلd�U�8�V�q�+^��dR��,�p-Fj��	�1�Y+[�k�n|�VbH}`SFu�.�)`�]}u�d�R�����Y��̎�W��b�M
&	�{��nv�%f�2�P��βd�U=ᵩ�����+��N�{���F�Sˆ>���H�h�r����x(���5�ڧY����ȡ�s[�7���\2�5՝�.
�]؝�����.��:m�f�q#�}G�o%���R7}�6=j	̽�cbB��n����Avg1c]L�v��ҩ1NJ23wU���b�()j�-���OdJ��x,rUnʱϻow�3v�j����{��ʴ��QЗ�oX��*�&	�śL�hйԔ��n�8�R��-���8�b��%G���۞�����z���)a	�9�={y�zlrB�����뜵�݀������+�=lh��*�ae@�baE@�{WWS�T�w�U��pW{YԠ�u�"n��F�Cd��#�q��tz�"��6p�V�<��mNuJ�_dw�p��Vͨ�>w�Z]Kt֖>yڅ�^���,ɶfZ���nl��rŸXA�)U��P�7f���֏`�B"��q%He�Bۮ���C��-��C˥�۳� 
{j�wX��v�G�ځ[F�նhi�Ԕu�a�y��-�Hc�JM�֪�o�!�n�_��5���P�SQZ�����e�����O�m]Ϛ�)Ѿ�^⬘�sq� ��ƚ�|F(/�dʆJ�~����!l����%�i���ћ!٘�n�>(9Ŧn��Y�y��gt�2��_-$�,;W��Iq�!��DkS�����]�z3�.�͎}P�ɄĨ�4S'NhT�)L�s�Â\��6��+�˕��r���sq�2C�+�c�s�#ge��Aؠ�.�m�'�z�s�CIv��,շ��g>}}KDZj�7K��#>Xw����xb�Y4 Bٸ�y~��7kA�A��}k74Ʀ�ú�o�h��f�g���D�])�x�S��
��c�.�m1�.�[�A�v�/��+�:
M>=�Լ�mj�޻]���^(6�[:]G-e�w��U㦈�xl%9
K��X#;n]!S6����p���S��(Wh���NZo���4��\r̀�;gz9!�����-Z��!���èK���_U/��U��m�rj����[|�nIb�U�n��5,;e�	.'=]�|���(&�;;F��AgR���+�u�k��6N�R1�Y���7"�{�/s0{v0:M^fj����sd�X/[6d�C5V`�+R�X�%�4���.�ڨ	B�m�{
���}�4N5���Q�m7���g(��z��/�d�w�{V�Ls@6���{��Ϫ���q�{���ˠ��Ơ�{���Fi����ޚ�WY�_I]�7�95il5k0�J�8�G�2�˻��u��Xʳ����&=�ʔR��\ ��VH�љw��ti�s���ڽ��t��Kͬ�]�`;�����V-���7c6+���GJalt�k4-j42��BcwJ֨�ӻ��V�������}�8,�����ra-�Y�P�49���s��
0��=��~��X��v2��I|�� �f�5Y��ɮ#D��3��܇Z��͏q>�%A����L��[׹.�s�Ƞ�M}�n�}��v�xL��p��y�1�XW���o.t���&���`�Up���t���J#��.�t�S�"�^kZ#̘�ަ��W����#Q%�}���y�3)�oRS�0��J�(�Æٻ��8�pJ���Zv�SW�S�. �["W*�]�g7��r�2h����Ft{V�u�y��	�0�6�ȬYJ���e �����K=;u���1tD�yR:�V,*l��Y�ݹ���R�їJ����x���ym��2�_P��]�:f
%:��M�PP����Z��6��:XK�y��̺����W-6y�	0�y* ��+m�3��hsƕ��6�4�r�<�y�Ga;6P��0������*g��t��,Na��;��a��������Rsq;�&ާ�[
؃��%p�l==�XgK*�SKj%Yc�e����\����v� 8L� ݃'�%��X���'n_5�ӼT�b&�+�hWn*7"�k��vw"Wrg�����e1c��N���,jW*YY��[A"v}{����m�r��V��jd�}*y��Ft�0<�upv��v�vv�.���ى��LQ(\�j���5�|�Y(�)�Q�5r�+��ͷҝF������\�)é�aF�V9�1�#6�J%G���=�S�ǵ;z�ޫ�R6�#pܒs�ڴ�5�y���)̱�;0mu
�D�C����Ԥ�;ފ�E4_���5����ڤ�9:Z\#Y��V�u�O&O��W�q�/��u9G[��P�R�}A��N�N=#�\��|_�k�2e�q���9�`+|	�隟�����fq����~�]�-Ӑ�IC����:C7_R����z�[��v�H���;�Bw�r�ʹ��6Gz��
���l�����B��i�:/�j+�we�b=o��ۍ9s���a�/�eg&���vD����w�Xs�oNNI$�����y�8�c�ə��d�`W�B�r�,D^;t�b�pC^Uz�87#�؂��T��LU^����Y,ZL��T���G�|D��ƛR�-#@��bJ�!(���r8J RMZЃ�,������ 0��b$Ki��-�eę�����W{�*D���;C�p�� ��}�Ȋ�˼��DD ݎ�#M۰��t��Q��ǰ�;�4�ǖ5��"��*�Xs��H%���&X6cw�f������S�kK�����Zٲ�$�V^��3�Njd��J�\�b+7�ֳgK�y�M`�� �����a��Ϧ6�a�9�c�M�}�@��D=I��:j����
���q��͗�P��5����9�r�$�ߏk)�p��7%c�7��Xxvl�����3N��OPyM�'��>ѥ�uMo��	�?EفҾ��7�[&	8,�_5��-us��ޛ�0S���Wg.�}����Y��.�Sj��sSn
�.�}B���Y�+��
C��s|��"��E����Ï5M�cϴ�{f��+)�&����P(��]r�!Rx�)��\\�/;RX�X\�v�w��a�2��.*�:�5�}C��uf���	�y�VQc��[�UWU�
T�܎���@9|��g�{�Y[f`����l�C;���Bi�5��n��='�$3wvĜ��ʒ����[�w*ɵ����0.�f6�^ �Z̶nZ�F�V�"X8M]�:�M{�m�'_<���;RX��0������Q�:�a/$�މ�{b�%r�����Į�w�m5E�n3x�o��V�Q�ַ����݆�K�]�|�Έ�+0�銓;:;;8;L�'�����=���w�l�RG���}7��T�g��Í�L�$=l
Oz$�V|��3v�1�bxDY��l�����Ў.��m\U����J��Sv���T��ٚr,�:����hV���ڵV�� 	-�2[��v a�9+��OC�Ʋ����s�_�
�2_I��&*<췯%y�����&����n�p�c�w<��X.�`��(M��L�4��8[ݧT��x;��P��#'��B���ԕ�d���<�3�b��v��0��Wj��R���b^F�X/+R�`�"�:�U��J{��2Lb��]�)�f������#��'3��&h��:�!kY�Vw)\�OϦ1��uAF�`��G�mZ��>ɔa��
���;�D(b������|��������
��.�dP���r)�c�X7���	l��]v���9�t�ݤnݼH�Sj7��:q�ٺ��x�G 1���z�ћ��ɦL���Y�呷q�{��k��.��:��)7
v�+�3zH���X�.��TӜ�
Z�}f �Y]�zS�����g2E��Lq�pQ�J��80ɠ�ox��8��AR	�ޒ�J���p�6�nЊnP��L��{����l�b�qTf��,�5�<IgU��VP#�4&Ы�ID*����Xˍ�J�e}Ƿ���̭�]��0@ q��ɗ���&�v75��
�ؕOo�4C�7S4�7k
�����	Zҷn���٨is$��P"j�RF+:ã:�[[��ښU.F(�/pN���f<�2��+5����%����n\C�3Ћ����vgc��S9	�_ �f�1�w��H�m.Z-�2����N�j��]դ���O�w�{~I�QD�)�p�Q�0�VD��qСA����5k.RPAΥ����
�/4>�\��vB�q}B�,���67Dw֏j"��?=��Q#Zǡ�i�E�v�4c.&�� ��>�gCx$Kj=p[L�Mk%k3:������#�rj�7��ܣ�7��!�]��ޖ$�alz;q����)ލYɒ]V$��.B���]�t�T�nSMRѸ#np�N�A�w����t5u��נ�c�וH��:��u�l	�:�p]��Ξ�SA�x%����Gw�����N���P���L�%&bn�u��M��4<�K˄�Q�}���3ct��<D���vD�^� �\��:�f�B#�9����Y��	�Uk�1}��Wai+d]���ca��)��<T1a*w*�v>+]�P�)ز������Wcu��Q:o�baI��'X%P��v�ѓ:^2�]D较�`�WG����"�k\!�j��pռY�����$D��P"p�yX	��]��>�+3At�A�S�[��_)��8������5�u���w*k��Ptȴ�$���ʛu�f��p/�r���j.��S{CY��V��=bxtѝ�.���&��ۃAz�c�9�X�e	�Δ̵����KFJ5ɚ{Pc�����O5��|p]	��^����[��h.�]�,�L��������&Rub�stIs!�3 �-��=D:�lʚ�Zo����v��^T�-Q�2�*5�7a���q�曮[�S *�O�&�6�H~.����=���V����Ck$�i7 �Ɏ�ɠ��e�dX�!]�'Np��Z���لwUѣ
���d���hl��6wƩ�jH)Wn@iK�	��H�F�6��ؑ����e�n[9�:�E�cF,�y�y���bҀ�]���PdW��3"�f^m-�+�uwS�(������T.�Rl����D'(������q�}Jb�4�Y�Wgw6x� �y�(�k�l�Yj��OWܧj��eV*V*<��nv�Jm�� ڱ�J�"�m�ă�`7�D�Zt�B��`mu)�����X�]{+V�'��u�9);�D�!CsZ�u���݅{����K5��i��:��7q�3�j�Sβ��UNT՘-Gn���1@4:���g	|�z)>��E�5��g:Ʃ�u���֝����+]8�<�}��0i�8m=�[˟�p���oUpa*4��p�m������0v��U���=�'O��i+�3�*h<���N��tTNt뺢Zx�l��AJ�q�xm��a^�	�pqU�~�vV�˰��P<���P�b�>e���x�u��%�XXP�/���t8���c�9�m�V��q�������������a�3~�P|܂����е}��J�.YV.iR����1��ٸz�ȯv�A�v�R��7w[�bH�J�?�}���ffFm��t˼�g3�t�!�:P��r�ԎjWtE�H��*�I��B�o)���B���R}���ܔE�.�q4�Z�8�qBdح�ra�7���u��90�nA���J&}Xi�j��ް���pj�g3yY)��7jm����M��T$�n�Jr��Y7c�M��V�� ���*M����!��	������ù&|��2vv���L�<Τ/���[���\�)��6�5�� � !}�@��Y�n87�7X]�X��l�b����z��t��:��r�k[�K����A���j@̀�[�󳅹�^�{�qӨ$K]\4j�]���GJc�b*���k&�_ q�R PӺp��n��䑶���̴M�9u�t��2W2*s�mv�u�f��@N���bn��z��J|T�v��D�b��tUr|��,���M���cj2!.WK�R�[4*=�o��퇂���U�\ ���"�[�y���ӭz��Q�b�a�amǵ��J�]n���;��Y`�v��^�\�� �#�\����q��ӌ�KZP^N1)�$�
E�R���c6qK�tJVc'��hu�V��,d���II��]��-CM<���U�u�ʭ�¥KS�q�nA�j��=(k$�.��89l]17�[�S����c�՗���B��z��A�e�7/!�되^��/Ii�%)��p����{Py}��A���.����T�0�}X�wC��q>Ɛ)�����A�G�Z��\��,�7fE���.�G{� SCw]�����A	p�,��#�c���E�c��հ�ö��́ԨY�^u��C��cІ5���m�
rۺ�f�ţy�:��+��\h��;3�ʑ<\��k�Z�Fm��n)�4�ퟃ��`�'��1�McK���n�T�sMV{�g.y�{oP�}���n���ձ��g��i�5̊�HL����F�����I��]�<��;6
h�I�Mv�g~�$���V�{Y(څh8�gM��aj�27�ϰ�tF�J\�d�Fj}xQ���K.=�̲�f�<�e�o�`�Θ�f����:%�vȕ}����M�ݼ��|����=������Z驦r��H3������؞�(腭**2��Z�V��;�V:h�2��f��&��oҭت�ow@nc˧C��VfI�͈�r��s�;*��ǽ�������n̠/���t���=*n"ff�*��2a��H<ڶ!���@��X	W{u�ݣn��)R�����_.�$���N%�+�L��D����s����	}��{��k� ^կp�	:X_*�vA
/i�2����ǭǹ�CG�u��f�#$�-���hل��ו96����ʦ�Q��nQ;���W8�� YA:0���}k�i��aT�w4�]�H�C�#T���]xݴk\��;�h�����uH&����(� he�MY=L���׮��~ͧ��C ×V�B
�_Ru��69�(���|a�c�ٴ�����p���hV�����z��O1��!�A!���`�{h���6��ض����֗S Z�=_8w�X8i�6v���C���j<%���S��O
ff9K��P��;�{��F�om(;���kSqWYA�O�TA#گ盫��D�����ga���-�X2u��8E\n�h�D�Ф"�+wa�ƤC�$��U�Mz�],���	�
�*�7p̴�#/hD��U(��5i�4�g~IU�̠�l���[k&�ݩ��Zw�72�B�©�B�*Н�U;P�7/A�8�@=�ߔ��V��䯍�S'o��=f'oE��ɽ3��zr�2����$�$���Wn¾m�ᔕ��WR�:������f���Ű���4��5�2v!*%l;;��F��N
���́,9���M�U����G�|�W�L��87eu�И��X�����S��;M�E`�*;ṧ�s�ﴍָ�B��C���̊��o��{n	9�w�� ڱ�[�,�T�tgS�gqv��Хm���MKC(n�eax�w��0�!�.�����hm:��,�p��D�\�vPYۊ�9�h�F�m��q��WOvpx,�X+ !B���=u}��+F�4��,� ���զs�w���)b'��ŝ����)>����E
�!^�c�̤W��'�fә��K�ʂ�����k�Gi�,�1uK*i�A�.Q18�B�a3��ۥ���N#���Nce��Ǖa_E�eN�sl�����r=�w��"/�ى��7)����m�PP)i&��xR+�,�Now:d�.��V�ÿu[�3\���f`b�:ɽ���Z�ݛF�"�J�{���\l�{{mfX��� �T�3Y�.��,N�u͋�8��������\��p�Fu��`�^-��qsv���Jo
��xѥL�ni�b�F�:�Z�݇�ⱞ�5ǽ��EQ�	��LrP��JA�Y���b�N�u/����5��;K�e�۠
%�t]�͇mk�/3-gK�Qǘ�"�t��Ci�����z:5:��l�dgb��!�uurV;*���k묮��]%�7I�[D�ȴ�
z6��<�/n��Iܣ((m�Z���غ1I��zx�R���o���2��&���
�UJ�R�3�s,�k),�ߦb)qWL�T늁mK��mf>�+*i�Pǻ"ׯ���O�
;��7Q��WZ�pR#�F�]s{d�Q�c	�b<���3�8:�t�)Qʸ����{��ڌ}�u��U�A�����I^ʼƣ�*��S�ӊ��+wo�����f��@�d�,���f^���@�ᾦ�UN�$'>�eA�EVE�����Bn�Ǩ�4L��k�1��;��P@v�	x�Rט@2q�Bb���o�5���e�(tx�?#e�n	Zk� P�h�;r�6cǧ�c!勢m�|����i��·�z<�QZ ��iV-�{M幬Y�zl�vaH�V8�Sw)�ju�A�9\:��#�
��A�u��Eo\4D�*�0���Wg�]�U4q��W��v����:��K��m�fs�]'xN�f���΋��3PR����\#JPQ��M09��|�QY���Խ-vc��Hu2.H"D�y�-Or���w^����U���(�V���X����y�������k4[J]=�������-����h��ص�Gk/�;Kej�Wۗ����*�S�H�`��*��X����� �lw\c^�:�q�:&�L7���}�4�l2n��+D./hs!�F��<�ڈ��Y��$�c/ꣷZ��(ՙjde�J+Z:h��,��x��u%4�0ZЍ�4�����:n\�^�G��(��eAۥ��n��]��y���T�VR'l��*�h ��2fS��$hvV��}�X*���Å�!ՃN	�< ���C��V��t���7[����<b���O��'܊��4��aݺ�yH��"�R�÷��f
U)�f��&B��?���f�I-�U5���g����A�XS�������{���*��(��E����E�;.��6
F:,�֪�Q�;���Ѿ\�E�`�JN��j�y�P���tS���2�Lv�V����ą��z�z�b)�4�0:a_&�b�I|#�N!Y�C+�[��z��0'�YY�9,�74mZ�F}�y��a�:�<����NS�u�v]A֗N���n	#B��y�*2��)w(�`������z�Q̱c����;2핻��N���;Q#��r��r�ד�[�<���v��Q���	T�}z!W(��4�T�o:�s[n�d�dM�����"�/�lo*h}�3W
�'��aͲ^��TM՜�
U��[�t�b���0*�+������z�}��3���/�f͛6lٳw��9l8_*2�NQJJ)&?(��l�b����H��|��z��]����r%�1mq��X�F;Mv]���}�&��؇eN�ێ���b[VT�[d�	圁�E�1:Xy��b����D��6�8�cr��2k:7��� wY[�F�_f��������j�XDwCh��p�5bY�="��QN�Z�lF@z<�Ry%[�}B��ɮd�._E���w��F)�¥	O/��u��`ڹ+R�jJ�;���okI���0`��u����Ô�y\&�)RR�C�`u�c�6�{���hڵo�V�PV�Vle۽&G�W^�a����&jwR\��Kݫ��=t�jkh�W��ژ@�;���f�X�{ºD�3 ��+ˑ&���t]Js��i�P���`�j�˥���\y�F)�ۇ1�wXُMdz�dg�T���;k"u��6�Z^��Z�Y�-�L3������q�
8:�6��j�:�g����;eq2��M[p,N�5#+[}b�$�����e,�%3d��!���.��}���]��m�`��3_���3""�*��A��#�Vq��C�Ι��}�'i �r=ͪ����ౝ"�Ø����4��V{t+.5���]��qs��9�[��^�����Y�p{kQ}�plC����E�(��'S�sNhs7õp�$KMv7[)+3�͹�Lf��/��|݋��ҔAH�@� ��eF�AB�HƜ����Q�4Zau8�c��7x��ӮX�u�+��ۜ����]������<X�/:�˶M�q�7��j1h��0�c%wr��6�ADF�q#L��yܱcc��͝�Es��F4E��/�"��,h�h���E�,�4�d��H<�#d�
/'ur���#`0Q��)& U�؆c0I�1���ў;c!A	�34����P�Fٻ�,b"	�\�w\6J$LX��.Q�E���2ch��t�+�L�sr�h�t��wm�t��i����\�.����Z�F1I�k�Ѡ5w]sWLDXwk�ݴE�v�clsk�2��kE;�r�)�s�	F"*4j*4�Q@l.]"�;s���O:�k���Q4cww:c/�Tx到|:�ߛJ��8�;��8o{�V^F�6j0��U1�Ó��$S��\7���X,�oN�|y�a�A��@/2p���Z:Co�*�ګy�U�ᮐ�E!X����Z���f�Ei�n^����^|sTo�x���x%a��{Փ>� �x6�ѳ5�]������y*)l��)?viC��y������Q���k�1ę8�׷�2ۢ͞�9G7zr���5>����rE�8���T��ݫ������q����ow��������ƭ�?^�!YR�({�9QWJ�l��@Tb1����{�Ξ�:fQ�ޝ�z�d�n��a���p�,�?@k�G�ՙ��E�{4������m H6v$
4v��Hy�L0q�������f+�8m��*���]�G�kΓJs�{��{[?{��u�5u�~4n`�qt��<1{�Z~ٶ��Z�~gޛ��?��8�/nRtu�K���C�>Y�{�s/8_A|��g�//O��{�|-�ߜΟP�&-��{��{N���T����ܷi�b��X��U�UER����'�8~�1�DoH����Qz5��+kM�N]{%�Nh�T<6d�9��x�YQ���̉����y��3o^%P�N���"��:�S{�;�Fy]�R�sY�@�=�&�Y�\u�u,R�L�j5�~�k5��6	cQ'w���n�;�/��vS�5�������{�
g�Qռm�wgv�^�Ñ$�'��Z���D���t�VV��w¦��,����=���[��tDp��l���f��26)��v9��͗Y���p�Ã��uxAV��v�^���a$m{�� ݙ�4�O�%���k<��7&��n��=��λ��4H�r�x�A�fK��}��2�����3y_�5���IF.A�;�(�Ӣ��g�Y�9�V}�J#��1��T��x�x����X�vr~����z�͜r��+`�輺���_�k�,vw�;l�t�����xdS�3�W�>�����Hp��2�*�w�Լ��Wz7GV�4y�`��7I�c^L��{������3�Id�s,�m�(�8*V���dަ�77��Vt`[�R/���/8�+��9O]*$G��l^]����s�/�#94P\����w�{��OW����ǘm��)�p�CIV�'I���[1�L�x�ч NF�-є�9�"�4��tjm.͎�l��5��̔�� �O�0t���_�u��h�����f�ȥz��M&{tϺ��s�Ǿa� 0&F�9ۍ���*�|y��tI;���>���?z�k{�~�,�Dx7c�R�UywM�Q�Y��j�N�S�z�/��n��e�1�5�k�
&�O�N1s(�c>?p�����܂���]ln��Y6)�R�G3i���E��2�G�vXc`:��_q��+)�kg��	k�;Ճg�}Ϥ���z�{��	�:$�A�]�ݱQT�xP&�2�1z�EV,d�bS�T�����e.8甆���y�e��X��z��S�#ٳ��_��K����ɍ핅H���w��[���� �B��2�c������ʕ���n/���Ͻ��}RK(���j���~��Ê9����˼{nc6�\�w%��ѓ�o,k�������͊������q��P,�KL�z��c��=#��]6�K]S���5�n�٩��l�tZO�S�j�u���M����!��C��\�畝�'��Gi䝗;�t�1Xy^c�QNG�v7Z뙶�T��9�,�R�r�~��M���y��r%����PbA�'��m���ә�oW۷����r��I8`�3� ���sV��s~T���m5��|_�u�
�/��p��`�+�Hm$�9���h�l��s��ݩ�{���iy��CέJ�k�Y��y���\�������m���Z����_�|{6.�u<A��ä_A�+�G\�5��b�{�ӓq��Ҽ�1�Ȃ���ٵr�}��I`�٬g�ri��O�o}p��X����\a}(K���g�w {�	m�^@`v s�����~�+�2Ok�f���?˞��}�=�}�þՕ��E�Х��)<�������S��!���~�'U��x�5<f�7����Q��=cg�7@�V\�[D���5cm 2{��=�z�������G��=��y����]^��Qȴ^��9}�dB���8��U�<�݅^�-���{��4�R�,{���
�	��v��~0D+�T�}���[�o%B%n�/#5�\��2����Nz��|d}wyKI&���ćj�����������pPI��,���;[�:v+*K*�I$�{˵7��#�+�տ?����Y�ŕ��'{�"t.d�N[����H'��|x��ߩ��V�~�O}c� ~�rʝ
��N{�h.>����Ƴ��g��ON��W�U#��[��DU���C���;ۻ=Er�t�J����ޮ�㽢$#���>=�*���?�3c�f�J�n��-=3s$k3��D��z�/����ɢ{Fm����|8LΝ�A�v��u��=��r��Ll��9CI3�fI����y��l�xMVaq��f��>����>W5U���"	�,V��r	���$˾; }�ȩ�M$�ۋ�Bo��C���z�^��k���ռ�k����ڝ��������I�m���!�����mk?^��K*Wh���*�Y��T�}�K6s�3���R�<Zڞ>����;g@ϣ�����`>v�}[���K��Ut
r�,�a�^���_]l	��a/�fl�� ]:��z��1b�Ք�_^���]��b��SK:��&7{�WM���Զ%�n
	ˀ#q,Inw<y�T�7��6L����#����z��y�؈�2�!���J�uڢ�3�]������i[ޝ�ݨ��j����8��]
���N̹O��͗-��o�@�c��f���i�@k��;�����׳�=��m{oW�VL��^�S.��Oq{~o��7>ӧ7ēRD��f�<���n�;{|Ѳ����O��9A�n@v���О�<����%�2r�3�F��S�mz��*�K
�,.��y��an��2�+c�����Ϝ�깊�ޖ�ȗe>�t9j����eNEy�ߜ\��[a���\��N�q�輳�D�oS��R3]�=R��1n{��
r�-�}�%�A]�#*���ǯ/�N�t�do��S�5��g	D!�ݳfa�^�Y�bcAƪ�����s����A�n̂{��������֓J>��Y��t9��{F�z��6M�3x���޸�َ�:+�H���/�6ύ�:f�)m���W����`#l�<)7���oٖ��onᐛ}.^��rRIp"r��Ъ��F��*�U��tM�f�g0#z`���H1� �q�ݺo�m��]�Z�����.Dq�r3˥+5�j+k��NH���d����y���M?H�g �X�s���C��&<z�U��5�V�ݍ� �h���ͯq2h�l¬m1�&�]x��!�7�r�#���6�=�t=���������I����g�����*�gۿJU� ߹��՝�k�4�1dlރŻ`���O�d�J�Z6��Ј���$�'�ԽU��.W#�S�s˧�*w����xH~󁭬�=�E�K�yoT��ٷ�#☞<�Tx%<��|w����wܦo	W����w�;���ˠ�ǩ<���y��������>.�`����\���fSSy��������ۥ��NS��������
�O�w��9Ň<9�W����T��]Y�5o>��r�"��RE��\NSq�� l����}�OPc�x��S��o��j�����=P��X��vW]���0�L���=���˱�ߒ	���z��ҰX�y�V@[�"m�;�ˊc} ���g]\[H�Uz��0X�K	�5��:qt��p�}��}�	�BޡR�k�t��77�|*��Qe���6�]s�Җɹ�Źx�\��er�;ۉ{ۉ�Nx�p�.\��E['���++cݞ-��9"��8"��Mz6��@�@��5ݵu�OQ��E�����Í�pyB�G�|켾�-c�|E�j��S��yd�M˸�*��z�np͜��w��������,�P�,w&�l�PDn5�I�lv��$���wQ'�� �~�N�H����[����S���J�x���n����v��~4�&�8�铕s�;֨K�.�}'�6�x��m`�p��b�p�Zxi'y��q�&8ξP��̢��3�v9����S�^��u/�uy�u*�-L���z{j�32]=>��m� �����1�/ga�����t��W`�Fj�ʆ��x������_xb��>�=���~�L.�TzM�yu��y`���~�ֻ~�]O7�S\�buY�����u��B[��ƭ]�i6C���j"l�0��)��j�<��{��o�O�,B7n���Tlۨ�c��C_'�y߳���qȪU�8�\8L;ٍ���� i�G��˒U탻S��S��u*,�K����o�۸]�;��A1vz7�C^�������~��o���}����!�l��G�����<��ϋ��UX��T����=��[BNݧ=*���|W��on���&�������ɆGDw�_u�9�g�(�7r@��4�z�{�n�x�}:��Wn���6����'1�I�0�#����;8_��ޖ�J��P��0g�=��EҰ7�ڹ�]z���hz�f���9M�u����g,/�M]�v�Ik���\T_Sۊ��䲧"�0��nhL[8�N۔�����9�;��a�s��Hӭ�$�ا����l�@"�ݓƘ޻�{��ͼ�,�m��k8�����:��4F�x���?3b��Ɩo֨.��7��X�<eIun����<f��?)�8�^>ܞ���I�}[�En��u���.]�LE��c ���G�,�����sI=�w���Z��
�y�̍Yn��~F	+���=d�8��r�걫���0�~���]lF�wj�ϋo.�|�W�6�~w��u}���я�͕+�J�{DӋ�Հej���蜈t��Ӻ�C�o3��U`ႶL���+���n��U����
=$8�ѨJ�#�t';�Rq��,��iџφUJG=�\�	�,V��5�&�<{��6�:����ރ]�v�z���%����u���p�h�V�zkğs��v������f)�W��c�����Z�H�$��'f7�q�6C��3��ud��j���||	�rMx��7�&A�}����n���<(X@��Bj�+�+٫�=���i0����_�gb}F�׸���9t"���V�i+�<��;�Y�*�}uF r/dFI/���S�z�zV��5� �4���{=!��}��*���f��a^0ã_#z7�ӓs�:r�'��Ǝ�н�j@���~�ob��U{m�?�;�7��0����(M�~���26�#�fi���v���wޙ�{�����s%[�c�}��������EH��f��Z��Q�P7����8o6���+��A�6q,�pfX�4S��W�.Nm��۷n�?���_J�݈�g:��*�y{Ǹ�p�}S�[��ۙ�Ur�,�bk�t]�:!&�����7�-Q�HS*i��TA�;�$5�ŝUy�0���ﯬGI�����w�����d���O�e'������LΎ�Y؂�%�fc%� �n���Jf䗥��+�n��5�6��Iөq�U��B���N��ٔfG:��4�wgU�E��w'N�ח��i�Msv��)!���c}y3��P�Ⓚ��o�]Dw�ngTo��77C\���h�.'�kN.��i
%�GK7��S���s!��f1(�Θ�=�]��[)��R{��[v4R��f�X��W�Th\�"�M@�y�2><�e߱�C
�*]���C���׭[{�>��Гn�u� c�p��-/�%Jgud:^�p���+�tӪn�wK�h�/�S�{ݺ,T����չW�&�֧�*T��cT𦮻(���0���94�;�E�᛭�Th뾖�#)�KDV���{���S����um�Z�3�W5QG�qP5��w�����8����O]KVѝc��۬V������I�S�f_&Iǌ�{��0������m���5Zs�^Z\��8ԡ�6M�K�2��DOq��[��
�숆^�@Q׺��䙒��v�ar�޽����2f)�C]�P'0wzc�}��n
����F u��h�5�:��5"�;]�=�:i⺽/��[nեY�n�[-��uә��{�2	��P����G,�g�QM�H���T�V���~�r�z��[�zx�M�3:�u�NzH2�|\喋�1�c�&V��j��� �y���V��1;�)��D��.\J���]IJ��w��挟d��z�]�Q�N
F��s(�r6��Y���v�^�b�.T4-i1�;`�r�pҺ�Բ��롥v�3���$��lX�s�]��%�-=�`q5����`��1�s)��v�+/[�
�S���C�Hk-�둌�D:�ո�����Yp��'���W�PG�oxl�I�U�Ll��c���Y�%R�=hpŖ>A���mڪ�%��>ߚ�rt��i�jn�6N}M'V���X�N��v��v�U�ȓkjuN,[8�*�:O����X���䩡��W��e�� ���;:�fr Ǎ\�:`;·-�{���ց�vF��������&���h��p��IIv��*k�3,c�EԬ_]d�P`�9:�u�GGL6�/(�ΛE�v���p�M�� �js��׻rcʴbz�{�,�I���h���#�?v��|j5\��yI�>�Qu!XX�n�S:Hާ������G��1�bg��u�.�Αm��u<V�m���'�P�E�F�u�K7m�	:V�L3�����(�2����q�V��L�Kc��XҎ0�o=ݺ�g�{ZX������5Υ��-��;GpN�~�}���4�Ѩ�u�����a�?=���h����q�,ZK\����.��t�"��4EE�|.���|��:�#���w]��<U͌a$�x���4�.�̛<�ʹ\A��]"��;��h�;�@%��<�.n[ι4���!�\��&�Lb#f%��+t���F1\9�H�spe�ncG9$�ۻ���6NTm�%s�I�P넨����<���t��'v�y׍�:�]�Eto�(��x��<���$��[���r�wm��:���8�wv��;�[���^9�^w-���^:ÆJ�yy��t�Q�]c�\�<�׎Bu�V7���m�uDl���u�$4����m�S���5y�<K�����r��9��t�5ۻ��K�[����F�urN�����M�S�������K��q�wu;���]u�uڻ���� r2n���E�ۻ�۾���p���k��pL�s6�}�M���<�V��vSqY�L�mb�]:I ƚ�O���]�"G�.�S���}�Ƭ�4n9s�z0�2����Qb �z�M].ŰS�@؊��Xl_،��t⻗Ot��bx?*���B߈5g|�*�^��C�7=D��XK(!C��p��I��Mi�6Y�x�w=.�����f�R�>L3���#)�Lz9��g��������d��-8ݻq��h��h��_N��V�z�߰8��a�yp=<)Uc�j+�'x�MM���Gl�
T� �1��N��@;�~ ���9>ׄ~瘫�@U��g�
N�+�d$E��!��`�0�����8ѧ��t��w.d�C\$��$��)Q������l��Sۼ	H
$�67�m3p�
��m4��gV0(b4H�$��	�~��ƩNc7��]oǂ�musg��t�[���в�"8�1��ɛ�z)K0Y�`��)��)?9�NV{�E*h��<�Yp&���s4P����jO�a s�G�?�ڝ���M)�
�c����ܢ���'�K���r7c����U�1������4�$#!�CƯ1��G4Ñn&67�����7g)Ƣ��=����v�w<tx��׶�;��`-��J%�v��;R�O[������wE�p\挵���R��+ZS��6���2����T�G<ة�]�46���T���ܳ�y[�6*:�9y���hi��3��6�I���6��t���B�˝ɶ�i����J]j��f�R�0��ybC����K"Ø��r���ީ�+�_�O�1��z�k^6Q1Dn��c�V(��l}�;�Z���y�Q�A��lia�=����8-�<��~~�wc�umzxt+�n�O�W���a0�c��t���8����#�̂���~��+��R�Zgji�y�t`u�����%�uCs�g�v�pB1,iN���ԟ��j/a���ML>Ќ�x���9���Ԉ�v�\��&;���H�P~|9�'G����-��s��k,�D��Ӭ�{Q�� �uo6�c��qn9��Y=x*�i�i���ξ��^��m�Y`�;
;3�.n{��˘�e�@�ƿˋ��f�G�py@~jݞ�Uʹ�u�v+X��vc8��������q��X��bz1�f�2��l�瞝����0BO0��L{_j�*K��f;9���O���EcW���t�P%������Á��D|�/�U��*��� ?%�j[t�&e�����18�=���^Ƀ���2��Q]�-��)�xR���
j򨶟wEæ���;=Qx+(e���>Z��sz:q�8��
�Ntp�y)�� bv-��0|��ժ�H��v�+���l0�p/p< 	cq�Z�v�<�;Xb��S��}/�V`�o"��݉S �՚��<M���-܁���F+�!�g��q�-oʀ� +�wo��[4��3��У%��K�N���f�]	����2Oc�"S��F��2S�o����j;q�Û�9KX*1m	�A>7�H"1�C�H��P�nwf�b�ñ�sҤ�	�)�0��q����Ǎ=�Dc���qӅٲ�XѐA�C���OH-�/��2�eS���7��+�nN���u��ᾙ�����ʖ8=�;�,GC���-y���@OE'-�vof��f:���PF�
�R��,�E�~*GjO�û4 v_^�>�H`���&��͍^����!�[��v�u;��O],`ۊ�8�,(,��5j�X~�џq���*�G��yj�3}_�Z<�۾t$檞�͵�hZ�R��[.��a(%�T�aH��`:q�l�����ʤ9hw�*�fpA�� >5�f[C:�{|���zU�6t�=�i����MŇ��t[M����̬����gR<dK��ǴBa����:;���0��b+*}��W7]]�e�e�qɈ���s�-���˼ �@��ݡ=�ݛ�d_�I�Uk#&)*G�5ģ4ۍ�l�䀩�w�`\��N����,��˵�����+E+�6iW�_on�a[��)�6T�]p��j��Mٮ8D!�ڏ��m͑T���'w+�!d1����Fel"c��C��+T�����YU�lD�����4��o��zN�s�P��yP4	�Ht� �˥�A�ʇD��p�c�	��Y�ՕO��:c6N��#��i��Z{l�:���(<���r��MW���������0G��降��Kիf�6`�=[�����&�����S�_�)	�Z����P�~,��u��ޜo���N�m�N��콻W����/\M!64�	�v]�ŲY3��Jm�R*
N�q��:�4�<���C��9�C����{gh �ҜI�&B@���|���L�ӹ�{p��k�c���&\D��R��]�7�衯��V��,y�H>T�о�3��]1����4�S�-�f��ȩ��!<k��}�ʒT�P}��绘N��	�DB`����t���mdl�(����{�;B�y9�0��J.��ʖ���:��;�׀���n�u�#�S�����P��S�9�a��S��jv]j-?1NX��a��'���Ƽ��A�䦣H��A�<a��-1�5�6$��&m�j�r��@u�����Wq�z?�[�V1Ȼ/,�+	r~E���B��Nۮ�{���l�3�s[I�
��zF᫵MjF��p�:��w@9䭐�㛧"0�;@�j��.w'�v�a����W���:,ҌP�SY��g��s�W\`����c{��g&g���}���(�f�� ���c㇀L?4�����8uO�;4ڬOQkep�ɱ�])���������C��;ID�����v���u,�C��?t^���؇mtӓۏW�6ɼz�캉,����"{{z;yKj�(4��z-���5�,�.�G�@����Z�+jj� =�5D�eb��<D�9�p�u�nr�Hv��%���=$:)�I��tE�n���:%�r���9�C�w9TM�B��ތ`�%�k��f�Yƃ�6����P�r��9u;H/���6"���Uȱ�{\���so+4˾�Z�t$E��8(-"ۓ�=c�푭ٸi�kݒXK(!\���oS�y�Q�M�UW�������d-��K�<X�ii�>>K���O=^��Pԕ3u���2oC�i�L�+X��S��^'k��[l'$>cz,��o�K��-���\zy���S�������sO0X6;�˘����!v�Rڒ�Z�X��߄��a@�f=n}y/B���(#Kx,�2�\-MY�E���C��nw �\�Y'���+Ti5�F��sS:|�R�x��ŵ�_��A��#	��V�����\n 3�ӻ�3.���^��t��D-g;"�x�0��c(@8�4Ш�7��5�1��֝b7.f\��"����P�V~�of�R
�����V�X��<�NSp�N���bwz�g���x���0BM�1٪��4|/����:O�"S�P%�$i ����^|��M�8���mh�J�+��{��|~��½���6p>�����2�ăԩ'b���Il��-k�v7�\��i����ѣu�#n��~^a��#���Bm���u鶢��K��M���-?'�ކ�g`íh�����zε�N��G�/.�aO����?>?���yɚ�ӮQ����U,�Fn�!{�[�n\��e���F6��%�*��ćy4�xQ~�@B�@@�'���Λ���1���Nʶ�_eoNi�F�c]�����M�])�*��+]�N����G�� ����c�e4�-Z���������:}�g*�Ν0���X�n��j�5�@��OP�n��oV��yb��]|�{�ׄ�^�֡�m�mC'��T#�����`�����TAmO��0�兩��J�7f�Z�3��`�gh@�i���cc�Y"7�?<��vf��v,N���e�˴�%��].�Z�p�砞m�����.9�&u~Ӎ��z=זi�o���_�?�/�7�֖r���k�X�Z)|!��9�e���/æv�3o�_�i��61�v��?,��>�Z���.�>�y\n��N�5V�:�e&���ެ{�.�Ã�}��U���4v���I�8�&_q���h���P��{���>��v��p�k�#٢�KS�Ȅ��maL�O��������biDYViM���f`���À�S���0�Mm_�R��l�<��O�>�����~�gs�߰�]~�8h����;����s����<,t7��RFw.6q�T2�"��=;�.2�BN�
�	�w�%��x�9c�y~d;�~�:��繵J��!?5�� ���X�]X�F;%���f�J�X^n-m5u"���2��Eڽ=:Ųs�D/Z��P'V�P��R儶��8�LWb/�窻͜��Y���\��Ђހ���R���Et� ?Bd�����"��z�s@⃳4�:)'��[zXb���.^OF7� �����!�z�@f!��˴�4�2ow��]d��9ޯ+7���8�j���+^�$�78\
�o'F@����B~�'�^���M��}��-UWM8N6�+�<��NȪ�פ���E�/��������H.+�AY���܀y�8���qC�f��*S�՞� �
�%�]ȜX���0��e�/EAbQچ_�w�E�B��yE�zw��#����Ш'lB S$�'��ՃWB͹��.��Q`�t�!]s	�{�����Ϗϟ{�ǯq����� �N�{L��hJ����;��m�A��#ĳ)>��e�́ᙈ�m�c�?���6U�Hk�\>>�@[�aaL�����h����7#�}�ͻ�Pj�^���>X�@kK�wB0��F������YM#c���1������o����U���"9��55���5=#�k�ƅ�P��peҵ�(%�T�G�>Z��s�KSld���wБw����!fpF�4���xmK2��XsV���.��d �����ή�$�T{�;e��kΙs�/���}�"]����C�m�Xʖd�^��sz����T=:��l�7N���R�0'�5yv�rb����W1ey@5D� �hy�S���h��G�ؼ�4�o��K��vבh<�ސHzJ<�]���eC�m�y�����>[��/?#��$�LBRή�^\!�u�ME��X̓�@f�A���+$ ��5=˦����U��e�9ϸ�6�,gR"�G\���S���j�U-�ZT��`� ʅ��Jң���W~,�vK�e`�V�f�\�^����¦*k��3��5������9�~��Kfa��t)��)	�y�:�r��1gF�#5f���ݲ�s�KhY�}�o"���1m>N$��p��/��5�`5�\��#�R9�F��;��k���;�/
�>�"������xO����,v��$�/ ����E�H�!>17��\�wo���g(�=r�9%l�V�D�em�ja���t3�����MִSK��-dC�bO���Yjv�\���|x��@ul�����5u��l`�X-c�	�"��u�&9-r}�E��;�3iVn\�K\�?~{��{��ܩq<��,�{$g��r�V��E�3�.�����)���kd��ްz�h����39��ͱ��/�	�A��"U4��<�L�\�{�)�����K�f�\1�y��U3Y�6ϤK��k@�f,�>6��	�7Az�j�w@⮚��Z~k�%��ga����_i'���P��sd�Zï	��G�[Y�>�d��u)�m�r��Raվ��?�Z�C���]ڌ~���멆�8Cu�f����\ff�hA`��z>k�N�6��Z�\%X����:����9rj�nr�u⠗�{��β���Űr`0c�������rb�TY{�}�pJ-�Y��ǥ�s.��(�|��}8�8���f:Xgc&7���!��kd���e�f_-��Oٰ��>�1�!�qh����zb�mv$�w�.����+v�3�CN 5��=4�-�v3],�A�l�/���hO.�i/��yl&�Z�y!v1G����S�<�w|v�Ӭ斔6;["�=�g�F�f�i�v�J� ���<-��-�;3V6�a��^�Q��L��v��H͉\�VQ�nmL�7RV�S��jw9�
��U(\�]��*ʉ�,���O:w\=x�/�����C�凞2�x����/C㽧��2�N'B9��j���m]�GkJn�������x  �^�J0�
��<���颞Ƽ�ň-,�t����sbj}<��ٜmIK6��9��T:��uw����TW��	;A�ٳ��cռ*�����=a�y�\zxR��	?���N	��u��L�Ww/$P�m��MAb�O~�Ӭ=�෫x/V��q�+6u\<��ڞ2v����q�0�VL��<��'9D�O~)M2���k�2�m�6,+� ���˷,F�����G!Q)ٶ���_	M�����'�b%9�R)��&����V�]���R�Rc��;�GY�׈~��`llp�:�2��
l�wR�_�'+=Ͼ�m�L�Ʋ#k#������.��$���0��{/~P���a��H���M�'g�ugM��v�
��-�n�%�l��LV]s��]�e﹠t������@�߉XtG���9+��j���緝�R5�73C��Vgm@�săr1�^�Lw=R�fA��E�>(����ܠh�]���ɖS�-.h*�Y��xE��R)����ƻ��)?2���G���l��n��;��hߍ���}o��߭������[�}o���[������pyK���G�V�a���`X���1&�F��{&�7@�y,�G�������Lcs��m؀b�)��c�O�ݗ���u�+C2\R�%�+��p�H�)9Z�"�����R�w�K�'�� [�S7���]�+a��ù�;!�s]��y��h���xu;9a=]�)��ZN^�A�>�r'�����U��W ��.�\��Lڶ��0s4w�����ꫩ�ܼ��,ж��ps�2� ;���cq�fJ.%xz>8҇]P�k�uh)���I݂Ke7ζi�2],W��[)v��u�k�ʕ�[״�(E�)ND��W-��w��yPQ�@���R��g':�֝d
�u���A꺏�%vej{$�/�\�76X�l�Ɔ���vr<�R�6��/h؅g��׷�n�[�|/yP�/pD��^��ee�u��R��Mg���Z��t�2���L�V;3�lݥ8�Q�nm�պ�(�U�[w\d�n,�o�G�u�h4!�Ӹ�T�����^^�-�a�#K�Vc���ph���4�nY�i��6���e,C#5�P��/z!7BH�t~� 'a��Ш@ߝ��dj�qf��\1���fIV��7���� ]��*nʃEo<�X�6D�7�Jل\u��]:��qB'��.�ٷ�2����P��u('�]i�}�6�$bY�����wDQ��}�c.�1|���e�<��v������-X��Ҫ�(�����s�Q],¤.�>��S�jr��6Ҏ�+Y@�Ϊ�V$�tF5�(�Y�U�6�Æ��y�ws��a[�I�j���_ r-|q���s��>1䫩y�E����I���|4@ޥ���:�NdI+4m�N���EEo����b:�����q�� �E ��ֶi��R�.�����c�wEQ���҄֗^:�lA�b��md�zê$B��vS�zU�e�7�)����t�7�,mk��e���G�}F�I֪9�p���䋾! q��Iq�����Zh9-���p����;L���}dn0��-��[e�/�u�o_p�v�s���� �l��� {�r��څ�B�t]hM�;Z��pɻ1=�EG��َÈ��qg� .))5蝧!kmnK���[��� �y1@��@��M��a�i���B��-��7P\�kd.��H��w���a����_F�i���ؕ��@+�Y�_|�(�bFi.sN�Dn:ǜV�:�������MpL�-�;�n����0M�Yk0A.��'}�Ȁ��E�YWZ�ۚ�����Z\)�4��K��[(>f��;����'i6ޭ!��d��c�	�\�p��X�:5�5J�}W�M�j-�ּZh�jS�1M���7�m�&��}�})��5y�8��?�v�.�OT���m��������9j��]<�������8L.u��c-�����X֌{��Τ;R(A����@��Ww�����_����,�.�p�Hر��%+���-�UȨf75�$C"�%��4j�AI�nm]c����9��(�wKE�t���wu&�K��%9�nk�4cU�żkƢ��4���ļ�ͪ4�v���u�j*5c`�ѱd�b���b�E�Q��7"�Q[�Lk���hأ^-��k�X���Ib��cd�;�Kc�sAQd��-�|5́o��ZD#b�I#b�Acb�\�XMDX��	��Igu���Rb(Ѧ��T��ԕa����bŠ�-��b��b&�X�%�F1��5h�4I����??�~/��ϥ惬��d�˺��R��ZXv�����5{�z�����0=p�m�]4M�&R�.��β��u�:�/������V������wׯn������~��~9'�=Ϲ�E.u)����yt���Es����Rx��l��Ɩn��Z`�@zgA�&vֲ�.���i'�df�+4��TQh�Ȼx5 ��YHA��̅��q/��� �������,ӿ߹͡��6��𷃳��L.{uJ��pb[$����_���li��I�2��o�?ߗ�0�f��Ũ@2b���Vs��gF�I�W)��A)�A���i�֞����)�<0(F0��ȹQ�fŔj�J��_j7�ix��kbt��92j+%��ҳ]�یY_��I1c�b<��s3��h���-]_���"��[-��֞6�X�]P%�]6Ϧ;%��y��?o���c��g!�ݞ��+��p��x�k�d�'*W=�B���E'V���a-ea�"���HU���o���vmk+��uB��?7���5ץ�'j���o�1j�~��=�)�I�3�j�_�6�宽����"mT���6�@�hUӍ��i�2��bo��W�賧c/Ȁ�b���(Y��w�U���~�� ��2���nm~���ix��y��뉃I�"ᒸ�)�i�i���u�6��ë�)��sp�+�[$t�Ơ��d����6�{jn�d���S]�I�k
�o�}�J���q��쁣����+2����Վ�p�{����xxf�vF/�;g��߃�_<�/I@؎�/@;�0яl�!�B~�= �깋Ƥ�
.��,U�3qb�F��L$���6Ⱥ���+yרu��M���Y˰kj+��9VY�D�֊�UoX1�c��m�S�X�GLT�[��
�,�熠�����vL0A<;�@����W3xc��$�n��x=�kB`���&����tf�Q����\]�TX,��4Uְ�݇�{ͷ�1�oE�'����ᤸu.3��y�&�e��ƕB��J�a�Jװ��֧��MBe%����m|�������I�;��ft69�@|Nva�n��,9�� �5gw�u:�I�7Oq���p�ͻʩ�;�ZT�5�e轆r`C��t#m��T�$��`8�ͤsř�W�����N�^*$�q�n��f]��c�)��yw@���p����&!Zw)p}g���XG�<w���D0/�
k��	��yt�L��m�lg�*�!`y�t�sI��R"ˉ�:^%��3as�l$Z�O��d8Ƽ��.�}�J�j��Jz�\\�lV��o��K[��s\�|�J �h'���ΪO��e���D�ST�fE�'���67�k]��g�L,����i�)��sjU	ƥr1�U��pxu�t�z���mھ���2uKF�H��M��w�S���a�����x � �����u.&Y�G����?�Xr\L]��5��2�[�)������$a������hۛ��sG.�-��T?W�)������G;J��J��KsWA�@���$�������E�ĿVY��,l�����(-QE�_����'��k�!�h0�2,-�9s��a]��f��ڋė�0�&0��vd�>����F����(8Z��|D�[L�4�=�����!��剚��BF�CA|��(��v �#���x�I)L9�/�<�軘O��Qd��Xػ������t��DS�S���a%P�I�NE'L�E��L�-5�c���ԩ꺮SU���e��wN�P̙�?7g��&5��Q�)�Ox⮗�Qi���,voO]�I�lx��=�"9N�߭�?��O�����`��pZ�����.��I�`[,܊#��z,�f��O7�-M�����H����3��8~�4#����u�c�[�fKS)��=yi��h������O0���TWJ����q�N�p�(�~����/Ǿ?v�V����A��/2���&(�`"UX�m�v��z�kx�p�8�޻ϴ�������H�(,u�u�Ũ�
`[�^Q�P��*Qs9.�VN�V0��m�K���U�ymC�5��D�r��X��[>Xwe�1ƶa���H�`�f�+�꯾�����+j�mm�լU�����ʊ��m3i|&)��Rca�u>_)�����ۄ�ʁG����_0�6���5-}�w`O��<ے�������7ҋ��1�!�����1^:��u�v8�\e!nB�mܬ4�S���	L 丑�e�^��<h9���
^��S8CG.�g��c����|nY5���H����mo�*��<1��՟ߕ}9�+��C�}������������ʝv.~u��Dp@�N����`��6�ӯ,�g������/\���W�L&�ޞ��b���������������W�c	�	�#��͜OX�o
�H�x�����G����F�����y�ܭv�[�X2��	BSm�R�&��i=���Oܳ�
�j
X�����7y�٬ח.%��2́C�2��ݑa�j���Y')D�>Ti5ߢ6�����p�}��={F�6��yӝ�a�
�O�ق^B�H"�	}�N�ሔ��H�5�����;���T��w"w��R�9��Ty����JY��g�*e�)��N���I��Rr���~�Z���K�t6c���ۗ��ns�-5JV�J�q�td�|�23�h��w�hv=�{�,�&\��y46��맖/]k-�F�'K,�?�o����]���0w���U���Z�m�v3+%1ɬ�p*�6\=�=��4��3���j����o���)�Z 	h�����Ԟ�7�o�Oc3k�����F�>G�d0�a!�"mN�p~��X�O~¥�0�_t�}v��S�(���E�\��?�%�qy^��D����'��C��5��:z�mS-N�u�{e[��k�b���nr>��~}ʿ,K�&8�c^C��:X?s�J�A'���[]o0�֙�u	��z`K�k��O�V�6�b����r���;_I�@�1x��罶�W���X)��!ؾ���~}�2)s�L:��X��=8e�X���n}�Nc��^��de�ت����P��`|g�D5����u�s�����I��23L�����w����>���Tz:�sSp��I�$&S ��F�������6{��E�z��t���R�L�a�tmfoT�]v��3�˶�/�� :"��<����.����<��D�N�L�m�U U5rɒ��eS'����Gy�yy.]LҌ.vJ-�e�˴�����x46E;��`L��Z��*+r税�����W>��حj���M@��P	�z���dgO<��|�;�Xbe�BX�*�[�n3�X��'�~c֮�T@�
��P<>s�vT�K�{:/v�"���d�ͱ�N�g�.U�q��h�`e>[um?u5��ص�̈́�,��MblL�ho"����r��<�]�`F�}c4���'vM�������?� <�� ��� �r�QjV9�������܂�^m�oA	��� ��@�5亱�����g��Ҥ3��mM���W��ʸ�^�\eLO;H=:ɲs��B��Ru���)�o�dZ{حw!n<�su�a����R��sB��<G�Ao'0�w/	;^�7�^�1db)�x�)f��
íֺ�r�Ob2��J��2S��ٶ�ȶ�C�� �Ɛ:a ‎�_2|fɝ�ֹY���Qjd��{�c7�ǝ%}Z�<�d��I}H��<��L��~�����]�K��x��u��s9G@��t�~����NT��~�6Ⱥ,�f�'f��ߙ����gnC�o4⛬�-���a	�P�sƼ����F��aVas�+�\�RX�GjHO���o=bQ-C��vv��p��e��.㛋�<�j�YcV�*�
:y�_�ְ۩�Q�.�w(������p}en�!�>mng���͹�E.u+u�˥k���]�0"ȍ��ɽ/oK5l��K�8@�y���r\0��g���ږe��E�1�{B�=3���j��TZR��u�j��Cr�}˨*��2mQ;��bU�z�e�-2���T�?)�M�P�@�ә�&|�\��mɤV���]Suᖅ�]��ǜ#7@�+�w�F�7I疓�vB3��@�e�U`�L��!�P�???_|���뾿m���5�EV�kRZ��b�j߯��_�����������C��������r�ƥ��8��3���<�`h�a7���Q�p��yr���wS7��]�@ÔXP�]�w�=��m��D����¼�(����6;s+y�vX�a�K7v��Cͺa@d��rޗa޼�A�z!�pCi�vG[*�xcp�:�9Qzݼ�wi��Z�@�>��|���&���683a ��B謐�"k����1�:�9����4ιes�S<x`�aÔ�b�h���Ʈ�2�[R���:Rt^�,�����G7�l^>B��R�<r���gA�c`�-�G;-�d�mT�3��NTO3F�hU�o,PH�4*�����ߏNk�ǫxi�=�� b�0�2`$#��̩��vR���.��W�c��BS+/��	�g\dR�����xO���x��c�R�/�M��~��l1a����^�8Я�zA锝g��E�{�)�$�0�ؾqOw0�6����w�Winژ�8����m�Xo=	�!�{�*̧so)��J�X��P\k./�����+��4����3��N:���=�E���j�4�\�
;b�E�m�x��m|VjI�
�U�Z4��=�y�v��	�h��z{[5Í���.��vp9�pF�[5t�4B;7�C&�$�4�2����oH�Gz�������o�y����|��|y�m�~���ѵ%m�V�Q������}��G_E�/-����� ]��Ꞑ���t(��I�UU��-E��c�������5*�S�N���-I�-Iĸx`>�����kO�p�5��f���6��'(^J�
!;r�����7=!���:����WC��S���|p�3`8������ ���6Q����<늑���t������TgV0��V�����{�Ү��k����0j���Dqs&�����<ج�P�l�>�C�t�c~��1�Q��~�>�zfy��3,3��`3u���!�9Lf�;���<�t!z)>��چO՛!�gޛ�Ezt=7��@q��LZ��q�Ű��Wӝ�'j�������%�c�a  ��LI�׹��t��2mc/^徔�ܦ���-�M�Z����ۄ2��5v'eO���b*hdK< ������{d���^=���>��L��I��"����zNٛ9;��J'(h�L�p��I�m�k�<�->ABi���11�箎��Z�z2��Bޮ�Vˑ�f�eU哌$g�B76u=cռ*r�|*pG�SH��y��S���,w1�l��h�3��ut�l��F2��� om:΅�5�Z�g�.��59�cg��W��]���M����	]H�,�Z�\��l���J`˗�sn	���T�J��/~ ��WL���iq�OV�fg;���F5"����߳Z�-�EU������ןaKZW��G�ʮa�{Q^�7���c��ɫ��x]�A��{i���-�ߢf-Cב�4�>[�F򧮠�T���#H{�F�*�tB	�Q,���YF�]�m�2PY5�۬�j�Ɍ���}�������A��D�}��_<%���%	�~1���"��;�8��ə����K����c!�����G�
Y���JY�D��ʱK0�e;�=J��?���p|��k��7"-g��E�WQ�,9�y�K�`!����5������Ζh����Y��E�Ffl�ǎ�ؼ�슎m���Z~X�A/Aqy^��A��������/,,�3�^�ᷣuW0T�]Iɦ��#Z�`a�^)d�c/^J;�������61����p�rڵa�PA��'�P�n�	�άԊcB	�k�Ro?5��M�J�b��l��wf�X��o�rլ�4p�D�a���V��I���z���Yƅ��1�שּׂ�#���5�nj2<��`ҕ����o�����B�C���`�r�Bb���_6���xg�e'�Fi��?�mt'��܈%o��g�@���m��������v<�"2/�{�AfC��zZ��oY�(A���m�s���d�8�<�r�m�֣��vK�I��r��I���:�]�T4�2��Q���F����i�]��(N��-u�<���[[o�m�[m��-G�t����ws!��QI�'�nZ��HqEA��E���q����lo�ߗ@��&{n3]�y��o�mN�B��j��!>3��!�
�����@l'� ��q�>���T�y�bZ�a��͵Ͻ�q����� ��W�z�2q�(�A�F\��_�r���l����z������26�]BG`N���zj��o۱Z����~���΃kw��A���z�͜e�)�=�y���w2���K�X��xH�<!�C�<�17!.j+������	���	c@%Ռ���o�j�n����CT[�!u�.2��X�N29��N�l�\��,t9E'O6���۪�Z��_h���v��/��L)��ƣQpꀸ�v�	[�f�gI��p��ŞDj싡�K�(�U�wź�j��x��R�jª)���l'�-�P�����&6e\��t'�3��Y��d��o��W��X�Mj��Qz�D���ON�����}��dH��8�.��k�\��p���׸�N5�.�g@�T,�v90�֣6Ⱥ�^4�iyC�f��;��ﾶ��ݾw��ߝ������[�������[�{���dUd{��*x�PiDB<ӻ��D\�b�
�u;�6V�L��J�8ࡻ�(l���ŽtQ�(�ώN�iJ��o��	x��ʔڰi�z-qwVE\"��V;;����렭�A90�Y�/[|�9z�*{}�n���CE�R�wo��y�V���P��B�τب��H�f�<���s���f��F���������(ڰ��m�/x	�A�V�L�����CE�n2�@C��9'���<o~�ֹ���V���n�Xx:#��	����M�cct����|��m�j��NS��v$�X.�->�Dj�4;�_${�E9�t1��t���5	Ze���C����S��ot&�8y1�s\�;�4,h�pS�{��-m�Ɍ�C����=���ht��m��b��;���Դ=ci��[<�!����/��J��N��FF"�7 ��k��έ����~m��"�v��g���'l��YY.�on4������/B�c�.�FEB��ا�g!��R˻���w�y�awQ��T⳴e���@�ۗ��aVt	�H�re�r�|;h�͸�˸��nC>3�����E���.�kB�j��	��{ױ�k���)�8�[��� :��h6��V\ER��4	@�4ݏ��s�+3��XFj��@4J�a�J�]�isZp&�+R��xzT��E��U�>�� nҘ+W'v���7ƪ��oji�@��g\�����9M�qQ:M�F� R�y�ۺ�pQynSwS{z�v��=~n�b��c��8��
[[*p�϶�ԧ[isͩ3���Pn��8�R�;	�.��}�Bm6*h�v�mʜZ�.��iC/{E;��#���ή��N}r��%s�Z�Veo\ӧˡ����7t�S��5��N�����e�y� ��l�*"�0Â�J@]f�]��r�;%9�g9��`���٤�#������8��	7Y��s(�N\�>s!���
<(\� ����L����+&p���P?�}8X����:���+Z�U��_f��ИΙ��.O��!t����uj�/��^8䈓�ǘ5NM�8��#w�a��ܒ�p����f�I�#����O:��zN0�vS܀头=�瀼�l�f:]��Ҵ��sCE�\�7��z,�BU��ʕ9�O]e��䮛�6:����kO1LpL�s�����x�](�o �x�J���6���L��]Z�R�4����6�]�\�5��l�t��;n��Z��~ېhٮ�0���D3���r��@^5�$�i\K�Bd����2�;��ʈk��i�m�#������xYri��X����n]8�n��]�-ꊳX�u:tE�=�(=�[���.����z����,M=ۥ�ȝ+#Rr=۫-�@�A8��
QA/��B
f:X�䧷��H�wF���Wب,��ܐ�:�}�TQ��clQ���BQb��cDRAP�Ɋ4lIj��Q��b�&DV���hœ�ƍ%4��EɌ�(�uṟo'1�U�IF�j�X��PY2b���j6�QDk&�%ADj4Y(��Z6�lQl��Qj�dƴE�EID�r�EK�����сyDL៳�.�����3l��
�1\��w���n܇,3��۵É�bR{Yۓ�r�b���~��+h��j��Vص�Y6�*�m��ZJ�7��� �V�����:�3�=OE'7&�Q�4�UY��Ae�/EAb|��0����S�ls�:�f��]ٔ�><��y�u� ����u~5t,�d닾*�
:y�E݌����O�	M���[)���R{p�3������@0���m��B��Ԭq�TA-�s6U�����X����%���|^ù�`0��f�69��s@mK2�J���c2ѻ�:w�5C����]5��ݢ�q�`9�8��3��w��!0��
�*��Jf�4N�wd)ǽ�f:���ۤa�,(q�.��2����f]�ly�3��k˼���K7C2��7�qΝ�`t&C�:���¶nq���N��쇝���� ��].�pE����t�_bd��T���5�z�3w�8���q^����5�my���] ��㐁z+$ �|F&���SN#�=}�]N4����=nZ��â��x#�Xd�\]��5�w�ʩljR��ج���G'�~��F�H�T��D��^��2㦽B�YS����?B�=-�d�Gj�3�j�]��m˳�}�j�n�7+pS�֒.h�x<�G\��7���d,P��e�<2�u�oR[|�c�2�6X�ӝY��:{���|v�/�vM�K��t��YqH+Ӳ�}������1���4�j�ņT�˩�w���P������ ?|  ����F�ՓV��Yk3x 0��o-\��mw�ߞP��m�!2X�J�o*�v��z�o>����֜I�����WkcX|×%�w�HC{CM�%��	L�<'<
��5EQl����~Ǆ��o��enJ��1-S�L��X"�U�/Bz�/�x�BN��K"�9�RJ�
}��!<�K-�����tWd�©��[��
����OAk�D�Ve;�yN��<�k�@�gJ络Õ.�olء����@$���*,p���>|����	�a�p�wmN�z7E5�����Ք_r5n����^*)��0���p��g�#�`鵦8F�T��u`I�`[p-Q�J�y�]|��fu!��#\f-l꯮��y�8�}/n<;`8��s,����(c�ă����.��uo�*z��V�T�Mm����z¹Z�T�Ob�sJ��m���4�� �z�w!�3`��N����`O���kr�6a�q�z)���ܙE���N=q��v嘗����䆚�&.-�~�h3!`<p���5�{j?P͐�/�u��Q^��;(q���yk[Q`����i�>H���̗��KǚnZ�y]�ǌ�V���x���[�M~SwN%ޙ-���6տK	�@�փbZ*;5�5��D�@�w9���e_qk�N�t�^�}\��� ��j^<Թ���$n�-KĆd6z䘲fud���}w�}��U&�em��F�4�#h�b�TԶ�|^5��������oPo?�B,[��*%�L ��ĩ��;��4�ͬ`��r���i���R��YY�>M���C��.�iO��ӱk"Y�! ��z��:�~��w�I�-3x���~����1F�Jf��3�%��R]�����\��t��.,����+E�.�M3V�/	��[�Tof�t
�Ƣ��n���*���	�$v��l�|i�����[<�wu��4���nr�EG�X`��XÍ�Ezw���c��ɩb�O~�Ӭ(�f=zޭ�SU��LkT6Ҽ�R�:qs���B%��L�C���"�@U�C�N+�K"�
SL�ʍ&���L��#1w�3��~����?Z8���Pg��B^W�A��%�����)�X��d�_A���'�P��;<�ϗ��.P�����!)fڝ��a�`��w�o��ӲrSى��-Ә�r��E[E�5х�>G�e�[S�	��g�s�N�4F5Dd�mI�Y�����t�O�Bn��9E��<�]qx˦�D���-�X(�z���2K'B�_S��<���[u�r��ǳg1����M�f��e:��9��7�r��1���3cxE��P*1+�3�9s�0LCf�7r�{i:Uf�����A�N������gC�2��G3i峘U����E��i��]� #���$�����٥����4*1TQ���&��K�___��{�?_���\k��"Yk؝��7�kZ��/d�c/C��ܫ�ćO��H��
 �:�b�^]�{��λF��/0{O>xa�zg�W:���P�w�6՚e'�-2m��Ky�?i7h=�?~�Y6��_���O@.ʨ`�0:aI��]��~}��B�(L8�V�=��6�j�&<�-�?vk{���Z���5V�?��X+�(zѮsk�c�xW��^VB��5?Ƿ��=�[�yMO/��G�^��3�}gk��L,sbvF�QL�T�0m�/���Ϝ�c����0_杻�Yǒ=�ߗI�6��e���g����E��9\a�ؽx_�w��������m{{=G���kˡ���Zz�m�׶E;�S꼓q=���w9�SI��R��<��^��ϕ؜j�	J��[(5yq�g�f�2��-Bp�ʥ�Sjj]3��;�hU)e"�$�	
�`�k(%��޷��'��׭@�;��)��� k�����<�ԋ:�8��2��ց6=��>��ʎr0�4�42B箈A��y�m�:v+��nk-�v�%_������W\u4�3���	���b^w��Y2JP�[b�����Oy]�8T��������H��X�A��U��^ڒt��X����E@�N�R��5oM�ʝ��VS�3��P��R��]2Rki���OE]��OI�c�~����mI�TU����m�$�*�\��F^���TXSP[s�\�G��,��|�/X��P]����:k�ɼ���0n�u�^
 ���(�Nl�B��U��ѳl'�-�W�N7�H"1� ���]uةgSEewF�Vf��h˴�I�0, ?���K�&��Y
���.�T\T-��9��Y���p������zG�\C-U;�I��\��9��฽����R�<��n[M��rL+P����Ay���S����F��aU�2��,�E�,y'����b&��qgN���`���ve�)aTh�JJ�;��'��󎧥'\_%��35��5�A����o������_��Wai�V��0~OO�Zy�LrzG6��R�z~����j.0�{�Ѻ�8�z7��=2U��pO5��d�`�#������V���|�����5U����T�sW���k��E�Է5�e���Ɂ���}�Q�9<�nC)����A�)?h�f���v�r�
�]��e۱Ɉvâ-�Ƙ>=���~���$�|���
���B���ހ@�Ft�������T�$���9��-�=���CA��;*��mm����a��Uؘ����ZkUEɥs���u�3G,V�����Իz7�ؠ3�����s�1^�f�h4�����$��K:�:���V?�����M�bجm�_O����������~?^wy|8����y�F��#�y�L��쇜d���r�v~�a�sZ)e�����q6��A@fp0t	�\H��I�j/��l.z̈́��t�y��!e��Ә�'+��ehh=TD�iW�E�S��T׹B�����ܯ'ەPᚗ%���<TI� S�|Ju�����{ cV��$�����똨s@Uk�jv���t��?�h>Ezv���Kv��E��뗫��Xљ��^0�׏�v�Ԅʷ
OaWm�zs^�=[�S[; ^���[�:��v��lB0=!0���{�O���PJee�S� �LW�B�ѓ�������&f$�MYh��ع�	��hp2����8#E�I锝`cȺ�ye�IRa��%�T)7o�ػv��K��.��@����Ϟ���"Uz�'�E�N�<��nQu�Mؠ���JЙ4x��6�wf�lCT7'2��6�y��B
��8Bn�OHLkУ~�I�T�2F]LJZ_�f���鬯r�t��ְT4I���\<x�a���:W��9���_e����,F�j���Ybo�N�:Gѐ.tIj2F���3S����_c�/�wK����Pom�����֭��#��t�����ܳvh�Hj^vv��U�J���44r����h�U2��sJ��ۜZ��'"�u4�خ�,|^ؔ�q�d�xy�LѢO���
��>���`�<��o �b�}
oT���+`[�Nл�z���wA�
��di/N��a�t�ė���F\;VSF]�Pڬ'��'f�lt��]	V0�]+^�)%� �Ү��k��?OH`�6���g�z�R�I[��� �H�����&���B/z���)���� r�N=fy�p�ze��ˍ镢!���UÖ�pP��0d!�{��mC'����~��=$=qh�{b�YKY�k����<W8��������;t��]��9aC�q D���X���g�9��!���μ��ʳʧ:�T�^%�h��u#<�Z�R�u�����3���V�=OE��2]hL��K��=��{{:���GN�4�$�4�PB�Iw7�i�y����yg��-((U��j�r`ʉ�F)���8���y�׳8ڊ�m91K'&���@f�'�1��t�w5�Xm��nD�[9�Q��Wh��2��.=$PUX�Q^�o)��J�8SI�J����w��oC����YP�/r�����;��b�h�a��D:�F�%W7;��h�Y�R�d����Ȯd�w �V��,v��g�p��K4�R	�)w��u0��Ҿ;*��or�u��qìYo����Mo;R =��X����V�+{��c+G�R����@���[������b�ٛ2㵦,�t���Ǯ�a렚10ѷBgw����}�����0����@�J�+������=��휼�ۼH02TIvl�xL��F�I/C�%:NVwZh5|��5�,�왞�F^�R)��F�[X�<͏P�=��٭��m����0Gic5u	��h�W�;�c5p�Uե�:�NW4	+'�kz0�c���L0 �y�t�X���SE�����(a�j���e�NBn���-?,	����:��Q����=/7����L�g����͇X��q"gf�K���7X�U�w�Qx��5�����>;���MuAa�z)*��P��hɓ֥��F@2��y�n~5=B�՚�Lh&��L$��::���>B��4�S�?c�2����#,h`�S�4��n��|��|�O�����x�~}��BՇR�u1��$0i�Ѭ�i�EvNs��f���5Z����#��>��t1k����.��s���:���3�<��{�̧Zw�9q��L�
	4ew�q���׍}�a �2�.(������v��K�ʲ'i�.�Cv��9���?<�Ρ<bK��b��1��|tE���6�k�"]�`��A�m��>\�*�Oל.��%57�ծ����w��OQk��b֧�+j������BI��>���%��3��[&Ћ/q���I��گ�����ΫJ4뛊rZs2�֬P=	#bZ.]�����;��u�l[�o�iHS�
<��"��!]ө�� 7@�$@D	�9a��9fff�2��DŔ�;:�[��=�>�^Z�i�oI�d���F]���i�m�N;���N.h͌ͧz=��uB�M�L��S��}]��\�專q^92b�m�Fu��"Or����9�X�p-����;Ń$S�f<��D܂r^m�.��X;'�R����u�{1v�V�v�܆%X� c��eEÚ��'V"K���v�Ӭ��L.t�PS��4��R��/ �ʴ;�����^u��%Tc�)�nM�uEê�D�(2�u/	;v12'���7ku3r-��1	�{1���R*��b6m��ȶ�C���F7+K�;c����d�P���(�!�������]�ʔ˃	��%�$Ma��*	e�A���Ӯ�`߰vLm~��,>2�k�t��ʗm*Rz�f�X^4���m����9-�R~�Z{7���vkg�N�<���"��z��N`ԉ:3Ɠ
�Y����L�ӛ��2E��z�����~��:ؼ-���`v5�����6?�|�/��"��8���<���u��yX!�բn��]�E���}��W��j\�Gz��-3d	9�q3/o��OwU\��ڧCi���ʔ3z3GH�܃�mR��Y��2_v��٬��X�t��-=2|e�{Sxpv���J�m%J,j��Z~�j=5���S�.� ���_���<qB�t�o�0���cJ�X&�����>�}��-<P��}����y}ULMu����9
�zs]+ϓ����X���maTs�#[=�{�WHa��� ���c8�=�[��v�KD��`�a�{jY��Ja��R�l2�{�ӕƥ���e轆s ȗx�r�����}A���t$E���6���,�:އn�9E�q�.�aۭ���i:"ئ`U�Mu���{+��P�!��������j�!�a��W�nq���vyC�{L�C�Piut`��F�/�D�WbvB�E�O�ݛ������e��d��&���j�s�Fĵ!�%�U~�����2㏺md��q�8��h��t������`���IïfM'�&�Z�muHĮ��.^�c��mAޮ�Z�F|;�k��:6��+J��zޜa71P潱L��!66rݴ�,�59�H�kF����6��T�79�7��ʖ*����B���y�kGX��?ΑY<�^/{�h~�T�P}�L#}^οӅIb�Be��JrT&	��U���t<=��O�������}��o�����x�'ՙ�[&�%���]�����Q��,�J�k��'��x���^ι�9�oeZ6�����8�[�k��c����t�]Aa��:�Џmź�n#pl�&hW��T�V_S׵y�N�����L�V�Y2�E__��g+A{˚�*ٛ�<FQ�����&e��7{}�6_F�b1J�N��������WȐ��;6�V�-s�'rΎ���f�N%NLup�¹dJ�n���IC7�o�e]���}�x�^�����mV񡏈w:.�u��[��v6�mvB�2"��!<�^<1���}��f�vua*e�Rp�'>���h1;�wg]I�Bm�\U�����y��Q��+�6�:[eKUN����c��,��i���U���jT�n�F*a5��cfM�����Қqq���X;��Y�S&b��sC坏5m�D�+E�lҊ�A
Z���&�Kl=�������0żw)'���E����Y��K�d�nf��~,�=�h����jSZ�3y�Fo��Du/���B���R��es��%;ǹ��E�;G2�jVd�*����^	�J-�[	�\�Y�z]Z��ouΠ��g`@��F�n�0a�O�i�n���z��#o��*��:-Ͳ���h}����l !T��-�R�������5�t�b�e���\p��]	�73Qt:��zu{�Y���x|�]�k�8ᥤB��䃤��Q%��}�9�<46-ved�;ov����+���n�q�5V�&���^�U�-�s�Į�x�`�jtw�sw�ō�j�K�Q���',�G$OY�:�6�'p'}��1���%���ՍB�ע�IUoA��N�eGkk^޺$�4��D�.���=��Ȕ�!�<�z��of�AD\$J�5Av
�Y�!gF�M|uη�%�L�t�Gu�M�䙫z�]��P
�G͡��;G���z�f��|#;��Ur�Qq]��X-�"����%�i�얒p4j	�+x^>
��v5,�2��
S��W0Cs��Q�96�c��+�٭(o�8$��}Q�kq��78�^=�:���^N�4M���u��Y��hʕ�+�ԞZ��V�ܣ�w25-��ۀ5�zH�� �i��>*2�!g�<�yU�Ws����H���N���n��׌>��vu�xS=w�&�V�T���å!���k5���j��5�֞�ݧԹE�w�}:�*���A;ٺ�6�S�!Sv�p�؆�.�q髲�k���]ʝ�y���9�*�Y�J���b�8Ae�S__�4��Κ	�Yj����kG�Ӊm[�7�^
@��+��Jjwh/���jۤ�1ݹTӦ֩�{cf��,��ƶW7A0o��ʡP���oV�ڈ���m�kA��tk8m���aY�'t�vi�+6oăew3�l�S��OX4s����J���FR��q�΅F�cq�^3aaU̫�<(�A#�	�Q���Q4���߇����m3Do�\�cXŢ-,��F�ÛQ����3Fѱ�6�E���X�6�ݱyݼ���cC-ȗv���cmͺ\�Z.Z7"�	�W���x5���(�Q��coђ��lYKy�\�E��B`"�kƹbЅ	�*񮑪)XƯ6�Z�U�^y�DH��@_'�qx�,���sM�^)Q^cB�u;E4�yݼa���o�X�$�¦�6��^M���NVrHW&`�czWd���<�E���>U����G/���X�O�o��!Ŵ�������D��^��):��%�u��L�/_vR��{J�$�段,�ZqOw1�Z��!C6;��==>���$J��iޖ�'�÷-�,C!�V�-��Υ6�������W��x�������̜3��uOHL�8bD�`茌�k��E㫶/	w�5��;�N'-�W�.��I�S'�?o����LY�>�U��_�EB��B)��-s��ܡ*m��r+}�Q���;�ի���@�^�>��aö�M �f��с��e���:��mo���+��r�X���RK�<�����
=Y����Y��0�d0e`<	;�k�XɆmǽ�]Rc�GS��N��披��w��2��/�>�mB��;d�g�����v�z/�چOٰ�}}(�Xc�TW6��L�����t{y�^t7�EzFhvx�Xh�s�?�x�4,�	�w�k�Ig[�pk��׺ц-e�ngN�,!���I�#�S����H؊��ȖxBKO��-0��9�y�s�|ǆt�쬊����u�ڻ�\�bvVhz`�t�?h�TK�S�"���=�0��۽دZTyC���4��e�S��y�+��wx���������t�U������Õ�d�L�VG��9Ԕ<��ae���_�Gx���Ls�]\����������on���\�[�7��;�T9��73MvI`h%���=\R~�xiזx���N�v{�g��@�ᙰ�,Dn���eO���Kׯfq���S7Y�A�yd����z͜O�4�b��_&�9��`Η{]�[�cG�:.���,�c�mE{x�M��Pd�Jx[�o�~C�ʢ�w3�xǹ��8~��+�J����2#���"�J�nwA8��%�~��6S\�"�o1أݴi� �Rk���ƯΞ�o��!@�]�*^W�A�K�FQ��l��^��N�ގ�E���65H�4F�?��n8�T���@1�M���'^��h�`�d�b�{k���l��y����	Q�_���g<�5�XsQ����}�l#�!S���;a�b��B�[����E4��aR�'!7K׹E��<�^���uyt���V���ve�Jz�9��B[�?a���5������(�r�j�Qx�H�2��w=y>;��ب�۪q��_��������|&-����
|��<���=B���ԊcPMc]锟�֙6�^iˎ��b]md�z�j���zxQ��5�$ɫ�9��n Do+�{nh�r���8�I������S�F��᣹��n�v5)gC/(�lpr�������[�F�>�㚑+�{I�j-��a�ΩL���N&	����JѨ�x��Wܟ����~�7����	�ʒ'sᬂ��1�����	���8ȥ�u)�N����w�sj_F�-V�gնEsP/��:�;t�0e�qO���ϚӞ[���u��j؁s���S��Q�Dj���,8����ℿ���	��и�X??5�{���[����!N=�= ����s�N�G~�D|g���	���~U�Z~��%�ǜ��ƽ�����T�O�//m��.Ϭd,lc<:�Y�8���oO�,�yްoI�j�Kլ�܌�H�Ɓj;�Ŗ��#[�,���5�׮E;���'�^Bu��Ʋ�5���q7�`.����A�q��z�9�2w׏r�fa_sGZ,��q��l�瞝�'x!'�������ʊƥ�B~e]g�Ֆ5�9N���s�ڤK�`KjI��g�_[%�eǃ3�P.��q����c1ܺ�lSP�nb��GN�v�΅��u�yN����ʨ����8�/P�.1��-�����N�ܾ������}��Z]��K6�PX�;�Eш���T-Z�)�ߣf�v=4~�g���'��	�NvVZsV	z�bj�01,�j`��l'ie=<+;y���2󁎱_K]i樂�{2i��E�>.��՗u �C]����M���X}�Tҩ ��2V��m�o\࠷�	n�����=ɌӋQ�ec�WI��<k�'wT0چ_i�iN�̛�?���a��m������C��cC*�Y�i�]�M*L���_��Qz�D�78_7=�岌�~M7����[�	osB��A~���0%��.�T��a�E�g�W��;:�кs\��T�Ivng�N�p����z��Rs�I�)��B^���'��WWF�of�zC�?W߽�ȟ�H���(�ð��|�������Z�H� �e��B������z�΋�mƠ��t��u�]�+A=@������y�>�~h<y�\�Xf�4�b�I�Z�7�c��2�Z�PK�)~a��N�5~��?�G���f��qQ���{-d =�4T�u�m��jR�l2�{��s��so�@�����M�q3�D�D��w��"����|�&��XP�~_�oDz9E��Q)بv�t�vښ|b�k��U��{�A��\g	���\gג��O������Sۘ{ ޤC���2	ћ[e�=Z�������r�����hze�&���π��B,�|�Il�x��0|+���_��X2WuP>Pm9�*qN�.�.n50t�!�3��++^t�xރ;�H���?x���B���D��]�N@��5�^b�����D]��or�]���h�{7$��LݫR\W��\��w�Y.�8�:�V3h�h�KGA�����%�5M��� ���1��ƈmq���{�pנ�HA>j{�M�1�Ʌ~��x�, Xu�Q�����6����}_�����1�T�5�.{aV�D��Tw},D��D<���g��&֜�ԟP8�|oA�;�����d����J`6�HL�b�I�Wm�Ӻ��z��Тb�4�\���f!��kRcJq:!�C�x����O5t!)���O�T�	�B*���)c;���魸W����5zױ0�i?�Wڽ஄Lp�8N��r ��b[��R��S��f��X�3�_d�j��1u��+�w0�[Zvk�D&��'��5�"D��I�E�;wa���M�Q����Θ�+ͱ,h�T`Ӗf�a��G�PTͭq�vBd5�S�r檦6�T�ېE��w^X����Z~k*t�~jN%Ýp���``鵘ч-/,����S�0Zاf�����ݥ��F���sV��sז@���rwsLz�H���1Z��7�a	�G�Ü~�OM7k��_��a<�V��`��yO;
�Y�<�26��~��ߎ3)X�>P
���Ȗk�Q%~��x45���2B��`�O{�����Br�-�iaY:��t/���f���2��Ah9�u�j�%N���!��[�ˡ� n�Y��H�YK$���kU�ԥ�vKP��+��{G^�N�;f��yI=Ѿ^�����5a�`P��D;k���f�z��V �Lm�u>X�ӎe�h�]�L�� �<��=]�=��9,Ƽ��;)0����?[sVylG���#�_O�]C����5�]f�f���O�C��������<"��X�c����Se�v3].�=�&�f�7�w���(��J�C����F}����n���|���|bsۊ3���z�� Cd��iﻤkp��L�C�K��CyIwy��)��6p��-�>��r�p��x1t��FS��O�=�E�{RT��㲃*'&H�����1i�$bc�tkr�3��<ȧx�!ŵ�%�Eǧ�U�����Jm�R�&�,SI����N�~Ɇg���x+<�֋
�n��[�=o��02F�1 ���� ��J�j�q�J'vl]��&�v"�n�䦘ڢ�	)-���񿙄�x�O��@��K/�������\��&�;nwQ�ADI}/��.&���Li#I��F��6=C�������Y���KU�.u�4���O�յAq�Y�N���e?��F����m�+�qȣ�@g�	ja~)%�V"-to�
��q&�ͷ���z	��"���U�gn�j∛�]k�9����l�t��q��I�\�b��a�e�eu@�ٖ��.��öCvf��4NWtj��a�a�jK��*R~[�I���"�����х��<�!�[�XkEȻ��m�<5M���b���鶢�.�ft?'�����%�o)^]4��ꙶZ�����Ӣ�[M�~a�0P�a�s��lK.{�4�c9V���(�R��]'�w�ۉ����%��x1���Ã�$7����?CѬ{���e�;���\��H�5�5ߴ�O��-hrvi�3sTv�[��n���F}S,r��i�k ��~������	�r��4- _!ޙ���R���Otn�Ó(-��9t���y�����=B�z3�C�<	�L>���[U�z�����}��X���9*�e'�23L8��z�j/�ܱj�����Tw�9�l�D���C!�m�\H�+zC��ÝBk��v�ŷ�c����/C�mߋS���@rU�E�_�����!߁��"c���N6ۜ�輳L�[�yڂS��W#.�)��l*�*�������{���i��RO1  !���"�髟W^lV����G���b���D:[_��̓�y'ګp^����oX�q>��*FMs���NE.tƞU.ʘ���gg	,&+) ���",ڭ�+��%ʯf��hJ�f���g���@[J۝��P���f��R�p�ʇE[JW���*WVY{q#��E��S���FrC/R�4�����=�s,�9������=f�2��-��s�{�`fI�1�z&�c*+�0��i=)��nD^h��D��J8�j������v>5eEÚ��'B�Iq�1<���SF_h�1��z����� .c9��k���Z�B��,%�T[l����D�s:���+h��y��R�څ�p��,Z�!2O~1��$����V)]��0ɶ;"�u����u�Я�=����8���p�i�:��c`�W��Co���i�)� �b��E��4
��mc[4���7����z��lݮ�A���	� �cH�A?T��ʽeS���)=Z3l���R2��n+!��zjr�t������������6�� "�^W��k�9���OE'7���9�4�R�W�9��N�E�eʝ�i��s��`%���F�ɤK�b������Ǽ��̓�u#�C*�7y�|w�~<�c?��=�.�)QaK:y�z�(�a!=�}49Z	�@���Zx	�O����y~�.�&��;�Xe��vBm�3�V�V8��V������Q�P�l���0�?�����e���NS3�t�Ѻ*�޼}�� Y)f�:M��I�vk6�Y5,W4J+M�xG(�i�}�X =��E:]��`�Y/v�lf�60�mvY�n�5�O&<���U�u�����eX8��[{7���@�2M��%���M�;�j%u𬚹�a+{�P��~�� :��R̶�mՅ*�t�=�i���R��z��C*�y.0��9���9ت#��zU"]�@r����~��,�:��v�9%�8�s��v�v�4�Ǟ�m5@���=�\���쫄[u(˔�L~bM<����a�����DR��z��'�^J\���eG�g�p�v�Rx���ca�{�m�����`L����!'�"���K���ym�ؓw�z���Sv>�ydr砖HB�5�q���1p�)�=�����C������q5]9�Q�!m:��j�eT�5FB�ve^��)X	Q��VUKM=L34Vg����+�$���vں����l�#��-�b�mT�5t)��HL�)�3'��"��u�l��v�HsF\]�i~쳕ֻ�[��b�0�2`$&��CH�S�]Je~/��R�&�l�H��5h]3��+�o���9�I��c�!Ŵ'H>B^	�_H�5�=2��*��ejDn�Nj:�=��M�A<Suy%I�>��{����k�H.͖"�BzcXD�Q���$��\�
���I@9����&�#���|*U�<��$�������EW��V_�<��y�Z=�W�����l�gs�U�z�T�s���V��oZ�Iv��0�N����[�˺崮��t��Fج���*��ݛ�4��w�t3'���ߋξ0���]ctS%�a��`Ӗf�a��@AC64��	���LT��r0�Ed��)��t+lb��*�qWKը���9cg���,!ã�g�#Ǣb`�'�F���b7���ƈ�����Q�Lh�r�ك=�Fc�ꊺ�B�z4��8xP5���e��gz�H�`|��>��zvi�_�����J��.���A/t�J9��3;��Ӿ4zi�ڢ1]i���ql$�`��:��^�;k��d�6���M�r�1	�^�03��`)�-�V�n����D̖�w%�P�Q�����&4?�H�Y��{�f��W �]�:ܴ)-��?�����h�1^:��{�C��zA���\LJ�.pm��֘��e/��]?o}e�|
��6q�60Hz���=N�_E��b*�dK<!���ո�4Ryq�J��1xhu,��=	�{��זe�Od���P�%�<�M���6��I4S�:~��L�J�v{
��?=0<yK�������[`ԕ3q�A�Y8�2G$;����z}�^�w����{���o�����\i����V+[�*:C7��yke���]ϝ���Ќn�&)�f��Ʒ�M�����'}��VZ�r��UE6��s%�m�F{�7�V�x��9_&��W�Q��ݽTWP�yu��V���n�ŵ��W@I�(�y��;�PmMG���Qz�0�l�N��N��fNc��%��OF�E�R���S����4�Gr�+Q���CY�حi��7��d��F��NK�؈�K�/D�!L��S���T��W˪�ɜ��L��X%����4�#ȴ�SۇRB�̝]q	��][��6��T�8kf�G��I����z���M���K��I��yN&CA�ٕlݢ�mu������6�_쮵����C���H��7��
��SP糯��3����싡�s>�jwL�)��ۛ/����Z��L�眳�7��	����ec8gRźևL�A�!5��-+gM*�x�J#/7hu4R"N�wC��s���l�/Aԯ\�;�L��:��:tR�{����>u��Ո�h�)�{�U�������u�tW7D�L��`�4/C��j�НFb�(��l&>�j��U�T��'������Oqs+�.�2WZ�K�0���;��n�v��C'�r7qu+e&Ζ�pt>����`����y�W:J����r^�@L�]���su\��"qj�|�ے�����RM"	XCltX�WZ+N��ep�b]C{�S�C�,�XࣆmJ֜!��6�����:���OH���p�'�4�ix���;�tD����vA[M��J����Ack-����]$��&���ZI�j4��f�s��K�gkd�U�v&��كfͲ��5�Y�Z��:Su���
C��Z�Q����s(VC�X�Z카����X.�/�]����p`6)RyY�p�剔xq�@� /��J��꼍�6ֹe��M��|3���ꛚ5a�/��+'(�f��nа�SJ[�,؝y,s��Y_x�A��P)'�z9���m�S)�`�`��b7]����,YOv��9yl�vG?������.�,�FsW@�r����a����#P٩Cև'on;<z+�p	�VŔ�\��a��r[x��^mB�/�%[��!8�*�o�4$݃!�t�$]�]Z"���[˧�MM���Gym�0���h��j���������{ovEWpL�^^i�Ť���H��N,0�2-�6�tFU�{�ӽ���[��[onAn�<c�Dί�ܗƇm�+]�E��Ocݜ�	�6%-�O�t��K$��s��v"
��*�Hs7�3LM���:������4�;����Y�7e
�G��ˬƷu��-�5z�a��Hm3;f���Y9Ƞ ��E���J\�x]���*[����"��b��r�_M���wu`]
�lv�"���DG����Cb�����[s\��O;sk��H���W-�r�nm��wh3�ƹ��X��k��n�ɴQt�ck���k��n����r-sn��h�9N������N�����QnX���E���sj5����U�s\ۦ�����Q�mµͻ��l��k��m�\��sF*�Z�^y��mN�75ͺuݢ�w;W1H�Q�����o��裡�`�UI^�^hx��i��Y��P�-V��E��Z\g�����..ɝ�䘠�,�Tke,�gd�M��M�9K=���xdڣ"��0�������ª�	^�W���ټ���7�֞���l��U���*�Д�X{��oV�^�n��x(#K�DC�]������}��2y�����M�j���D�\b[y�4��Mw��D8�`?��W^U���3�+���FM>�M�»]��7B��^1�'�b%9�X�F�[_�['��b2rWG�f��jZθ�#%Uv�e*c c�f+Ӳ�m{:Y��2���I>y�Rr�sȣKh��$gS��y����\�������O��0G�9���Cv�鶤��K�ۦ�����)�����+"�r��{4�=�,d�a�x��Ñ�&6%�=��n��Z�xe�Y#X��Ц�|���pe����c�Z�~w!��R,kc��:r�4.�	�+�_��Ơ�ƻ��~�솥:b�f�]���i�6�t�Џ���o����̂�ฆ<yO�֯�O���<���M�vؙ�K'k������<�����|�O�l�W5��� uv�vCC�'����{��ޡlQ+�lC�\)�7{����ݩ@�v�lN�w���XM�T�_8���3�{fN�ׇ���c[�H9��얍�=�;�����Wc���}��D�s;�ZP�T�wLw�u�A;��J��K�v��^&�lP��Ipf)����:��w�������,j_����uC'�ʄua��d��aŜm�1\�_��j�;�Ѿ��}]�6r�kwJ�����섌�i0q��H�J��?>2'@�4]�ñmc�ĝe�p�[�t3Ԩ��9�RG,׍W"]�C�d-�<:N��q������m�W'���dhT�ǰm��Ǩyi�n���/��V�}῁�~f�^)�����E�j���3b���a ���r+z�we�3g'uPid8��j$γ�?�cW�*I��0?ߔ�5����8�7Fv�_L�ή�6�#����	��	cA.�g�c��^��]�C� �d�Iq�5�{E��m��e���V��+3ͭY1���2׾QIխT)_�QaM^nq�_0��uy�J�5"�9%�vYQ�����eK�j��D��LZ��	�{"S�)P�j���������̏+ۻnʳ}r��P���HB1�C�O��A������0�T�(1�����Yu�t>��蹚��}�K���
B:q=y�-ᄍ�|k�9	��= ��\C-�����OS���F��Ʈ	&��0eaZ���u�u���������{E%N�����Y��9��mW?�k�.�^��K�ގ�&�5��z���KE��}��[&�����HS�+�u�ָ����C[����[)��p9���[�3��#n�=���]N����2bvdQ���^�Wz�mƙ���s^��^e��n�������[P8Z��r����I�ɺM��`��U3�U�ѥ���&;^ye�/V
��s^GjO�û4���`�۬7H�	��G�5���ظ9�櫷(	WB�����U�<ƭ]k	�OvMr��A�O^ӱ����V�4�΄��v�qNX���C8е~"F8�d��V������PXI��^��ܫ�Ŕ��7]-�ͪo7�M��@�3:�)��9�e�v�jO���X���(����nY�`��bb���n_t;�{�6D�ǐ04g�0���~�eK2N�z]�p�8ėi�ku�V��z��Y��u�ܝ�j�v�tE�P��^F����yF��-�����D~�狺g"��a�S�M�9H�'6�˥�A�ʺ&���fq���B,�����Uv��`�ょ��V���y�T�CkO�"M=�G=y,��&|�q�髦.W�)� ���f"�Iq�ڎ���p'.��{��j7�R��7���gaT-e
II��zq���*ǟء0�=����	�y�F����{�2�r��"�EZ����'u	⊮��]j��6��C��N�gF�U�y�n�[��A
���h��.�sST7nS�2-�j��(�����2�A�ټ��}��e�m��i�����W��r���j��������?�~F�d��U-�]Jm�R%�D��	]�.�sֽC�Qp.�s2���qF��t�4-aE��g�~0G���A}_x/��W��ȳ�sj���[T�:����Q�خ��l5��"�d�=k�<'�|w�!ŴH>T����D��צM&&_5��|űѝH��b[�z�n��*L)�/�P{��������q	��r�X��,��
�n������+"���J.��U妡��`Ӗ��^<�� ����q�R�n^�as:�FuLv0Z� �,�J��w�5��W/^����,J�0���p��}���T�v�U5m1�q�!�p�fn`�Ҽ>���|n��N���s'(_&����]�X㘝�$�#��^z)��vm�5;�Bn��+`��9�����j���(��t��h�ҵ�(%�<�0���C��~�]}KF��((��:C��H�/"��NL3n=^��+�I���zn��։[��Vgq{=�t��5x�f4b�;0�����u�Z��z�}�����Q�y�N�I��hkoQ�e��,���u-:ukq�R
4F�����s�A����Y׏��GE#ъ��z����G�P�lC�U�"	�rw^���j1���۝���+Eӻ�"�S6vU,�����i�VZČ����FT[Ha�ͅ9vU�>����\J�Q���~,����C��Zey���������9����$*"�>�jw�E�V���lND,�Sх���s�8��$=qhO�b�)�cb*Ն���	�����I�ǞE_�f�Z��5g|�s�W�ܾ4�3�L�;'�	e+��p���t5���	��=ڝ景�][�҇�l�����-b�|�=�/fq�jJ����A�,�`�������&*ɞ���~���y���"���kKߢ����V0Ke��7���a6f��Η;]cV��V����}+��<#}�1U�����Y�~c&�"!�.�]L;�n��kw�9M����.�c��d^�R�e~Ti5��=�s�:y��x��K�dh�އ)<bTӗH��X��BG	��E����D�7�R)��&�}���#=�����:[/٢+v��Pb�̄R�n�=<W��0�޳)�N�T�烘��g��Q���ه5�.`�X�R�#3B1��y�0�a�	���G6קg�u鶤�T;t\&��9E�+�%��G����At�5���\;��zGkT��{��l}/Si�J�u]�ވ��u�/ ��� �-"�6 æWKѿ�������S6�@JlfV#jw�w�
�������[�*wEض.0�oNL"�h�.#�r�cvS{�G6�>��/ϼ��'����_SM�>�~��lkH�!�c�.|�4�yʵ���Qx�+�CoM��G�x8��/H�S���@T?yċ��t!w-��g�'P�_�y�1���#0w�B�����g!A�x�r���Z�&ެR�@U2͕�n���A_x.!�.�_���\�5��>	ܛͷY�����_Xe0�c����m�QG�ݺ��P�n�`ա��'[�bw��~ܢ�P�W�n���?�n}��B:��N�3L+�@���ͥ�[���?��{�xs�������c%�cG>1Ƿ�>�*>���}�<�z:�w�<lZG����J�x��	�͹Z� �:�oP � �E�5��N����}�����¨g�	�:������V��ϼ��w���wr���Q�i���E<,�-�D�P|aoql�ؚ��u��kU���jxuu�rea}����6��Y$5y#:�@f�2��-�<�ӽ��``��a��X��N%nk��5ޯ�4�ITV2.�}na����ӌw�.Á�5��* ��ʧ�?L��J	���W�=4Q:������.WB�j&m]���r4r�yc�=뤩�|��j(ju�UW����1��4XV��*r )!�A�w-O+�����:H�5}إ��&L� �5H���,���\��K��Z�����7�<i�Y���\W�bq�@�nl�<��2׾QI��j�Jª,)�m�5��uQ\ky�
�٭�cS\:i�3�������k�f��T�g���'��)��)P��JqF\�k��+����w&��r�04��)��zG�vH8��!�},�4�|o�G5)L�(�y\Tl	�Nf+�Nh���B1֮4�N���n8��i�9	�:츆DYT�fP�L��Z�Rs�/��I��)�����-/#N��s>� ��`��C���S�I�Ȝ����|U��+j�;e+��aV�s�r˔^��������cV��_�V���z�j��,U���N�'��GC�8�¼���ի�a>OvZ��n �b{0t���c��f~3M�A8� �����n�=#�k8е~u+u��Z��^��G0�.�:ԲL����z`WE���˲ Z�0V#��-^��\[R̶�m��)P7�]5�~�ә����$�mx��ǲd�K��V��ڱ��w�\=Ƀ����;0̹�l;iÔX7���h��^5b�;Ot�\.-�D#����=�Sշb�[�r��;��@�8_p�˩j齁T�G��*�R����;��w�����9*}P0z����"��S�k"�![.Ŵ�)4��Ⱦ����[�u��sH��Q���3���0o`�A	�^.���������ݽ����"��������kγ��;}#�<���#C�}�<��s�����Ւ�Դ�ro�G1?��u:�i��8!��e��ze��mᎸf����ˈL��6�n��i{����َv�ME����֛��Z�dΕ�CQ5�>�������E7{3%�x��C�OXE��p��k���L�[jP���A�,��%G�>�[�Q�-b:�KVḅ}�Պ�t9��u� �6r�#���2Y3�à�M��&Eb�I�,3���L�W���0����=^��³�/�����1m!8�!�C�x��|���B�v�ױ�g��i��e�R��EP�Ȼ|����z��!��d���^	�_<�^t�E��eP���v�����S'\��YX9�PI�&�|����ʔ��~h�����:['��\L6dR˶�T�5pb�p�;B�y"���E��M�L�ux��,�^|�ݢT��Pd����|�a�63�rڧ�sn��I�Q�=/֢��_�PX�]&��q.|�8�mHQ0�Z�Џ%�FHyF�m�#[|s#�!�}��+8D��mO֟դH/��:��Tl{��>�q��1S�mD�=����JY)��sշB�p�}��R�}��4T��������f΄�7�#�goKw)�ת���DHvr�?���x���������x�1i���'f��f��'(_&�����H�~�Nq���Ex]7�Ɩ��t�k-�@p�_�vi�X�����*��="�^2�����[��]/t��`�����PQ�T(>�TQ���"C���V6�1����3[���W���-��K�0�N<fy��,ƌXgb\3P�`<{D"��y���8��<�%ٚ)f�\6��5����;m���c�C�B���'��iA��RH�W+%}���Mrb�A�������p'�
&�k؝��+��$f��KP������\M;N>�H��T?"��S��̵�/�]fYפE���g��=OE��yfY���,��9IwL^۹���z��s/{g^����Դ�P�a�������/8�|�/d	ƯjJ�����fWB�&�]+r����VÙ{R�^͜N{����EC�am���+U��`���4ۨ�7�Н���x����o-�Ɔ�@,SI�J���ј�-��վ;�
H��� ���mΒ9�٠�#K�O(o�esܕ�[G�-��xkOz�;켇n5i�̗o.�k~3�8�GZ���چ��uE��oE��CQ�m�f�11����kR����SZ�Gf�[}�����CS)D�X̝`M*�p6n���yhY�c���M[�Mw����<=�N��ugv�>
v�PȄ��ȹ	��dB�I��R��r��)J�py�����jx���ʇ�@���Ԅ�&z p�/����S��b%9�R)�y#I��n9�>Eá*vE��L�1�3VȵLi���	��e��N�8a�-e;�iRO�9�NVyV�a��R٨���;5�E=}K�Ә��l!#��M���n�鶢��K��mO��Z~Y�m���2�̈́;���oGa��Cuբ�
�z���#��G��W���+�Q�߫Z���T���{�S:��E���N�4�6ˠ�w='�q�b]�=���!��n�!�?��	�!�岩o�:���~�]9�s#���ʒ��֙5qt�w��Գm{��ٺz3��fXHA�t�'�㴲�\ҁj����L���z>�r�j�Ja����GcӇƢ��u��Hwn�`�v΋�L2J�����c�uB1���r؞������hGVI��Fi�-���*y���[��j�ds�O7�f���U!�C��v{L�G9e�ڑ�����	�q�.�8˱n���{<}>�g�������=��o����"�7<6�����g9��s�9*�Y#F<�4��Y�Ð䩉u��h�d[D9Pý.&�j�B��h4��@�:vs�9j�jN7ʑf��eВ�������'.3�~�0�J�������/J�Ժ���rly����u#�;p��x��ݕtБ�p#�I���D޺���: �J�Y�!���y�v���֗� y��#2�a���.u�i��j7�	J�����X����4�{p<#}h�7TƩ��[�t@�*y�ٗ��u�WMt���;%��+Eby��7>���^���:�jC'�&a'�K[�c�۬٩��e��+�h�Hf:C��.#�`�r�^������=��eE]���w���8����1�yI+T�.��.�a�[a"z�eF;��uII-Z5fJy�t�K7xp��zed�GY4uWN�-VhZ�y�&f��6*X6��t��e� ��b�S�|HЪ��F�|�ɵ/�GJ&��W-��pAN�yY]l)]��fV�!J1ݝ2�
�yT�pv	��W���N<�������wC��ݑ�{�4:$�#{j�p��#-s��=�W]��p�+Ver����0V(^2�M/Wk�آ�̊Yp����Y[;�k�h����?.0�Tv)gd/����zum{%d���aVӛ~I@m ��9I�H��l^�I�,���l��v�p�l+��ݮe�=j�-Q��3&J����$��tf
j�'P�z�J��g30����n��*wp17�n�l3�~r��(�V/{ۛ)�������0��d�����\_�y�n�{հg5v^$���3_[je:���^C��S���1���v�ͮ�y�I�����^¸5z(���_�*K�l��]���i��8�d����_�O0�	.�P+���Y����r�7�l��fm.��H\�3FZ�C���$qD	]Fɚ�-��QйWٗ�jA*ÂoUs�u���ln��b@���^Q����G���U��ܩ���i�����7��T�5�3�oG�,�	�����`�+H�o���W����{��&�l^r��ve�\�^*,9r%_e�t���Ч�(�}x�vN��+�q��������"S]�tvR{$<�-��dq< ֵ�XT�5�����=ϪQ7v䂅�N'�SfK�g|%*�Z%׋wU��*����a�G��
w!���y�c�\���2�hm?�]�(���s��bɒ����mEJ=�����y��7��1^6;Vr�[Y�,C��]
ځT}!�7V��nSۼ��#�����f�h�E�N&��V�E:Y����1q��TA��ۜ��Q���O��Z|���E�˸��"��4s��4K�;s.��(��I����͹ҳ��oy���a���w^v���s:r2R{��5���д)��PV� O�A6�o����W6��m˻���7-r������t�.�9�l��ِ�66#J-깹E���A'8AF�`�1��wW�@�$�1��W ��r(��q�9�6]�$�r�d�Ĺ:�"#s�wvM�渙 �r�6����u9�_�ۉD$�rHr�s��b��Q�t�kD��F���4wn��ӻ���Ѭ�n�$"B\��b,��w:��N㤻��R�� ������	W��G��骽�WC��,m�\{�+B�8k���sm��[���:8�q�c-=��cN>��o$%��{�z*|���_�xH��Ӝ�<��8[?=�"��E<v��3��[�dH��S������M{n�uIz#}�j�2~�{�c���gCa�}o�i�����}���T�������WIm�5mq�Mvl<�],��ޮ�V�t(���IA#:�Y���dgO<���0BNNrЂb���]1�]�ղ����^!� V5�B~k;'��%�%լ����=���E@%��^Rk�,�/٬?Ώ����6�'�t���\��2ױ�M��j�(�*��ۜf�;�R/=�Y��K/�WC�,�$Ao'0�w鄝��f�"�SsW�!2Of"S�*���|�n�:�66�m��.w�"����K"��oD�0Bq�z �Dlʅ�f!���]�M*L�.h��$���^,� އ�@����$�78^���H܁!�B~�= ��\C*M�)h�f�s�g�ޝ��"���*���1L����>��Pml�T�\W(VX���|׃w?X��ţe��y}��z���r��
�f<7,�E��*K i�q��?�H�8n��? /{���ߝ:��pO����%l�i�*@t5ul��w �K��+���l�W����Werj�#I��ji�{�ɹ�HDMi\S#o$2���x�:�P,xv�Z�gs���jn֭���+	,\0b�{Bbʽ�>�w�i)�Y�E�Z�&����n�k87WS�~{�9|�t�����"2OBz+�\��e�q[�Qa^Y��jº�	���`��UY<���-����:��>���4��1�OH���q�i�+q�l,u䠗��*�a9zp85-T`�m�͵|�.d-�;�p�3���9ݩf[]�XsaJA,�k��Vɭ��y�㻞��Uww'l�3Yyt/@��d����0���~��fI��;u�LaMZ�4��f��_N�)`���#.ݏD̻Hls�[9}��� N���О�Mq��E�٪�్Ɯ�\�P*����9�A!�rR+�;�R0zó���L�P&�y��^'lF�z4;�[b;A���<8^��:�&���65�^B!��~	d�)^iN��b�ֳi(^͖���/���{ �{=�BWI���ԪR[�e[XK�-��@X�㰃*�̡Jң���◪ʠ�]�_V^����/P�@�3��cH�1�H��`a�ѳ����so���|�&Ro\y�w��T��j�U���(W:�гј�1��E=�� b�|�I�ǂBo��5�e��[Y��6�I�Y�U�z'��=C��<��溄B����f�a��X��"�gJ��D��tU�x\�gs,�e�Վ�E���=؞�=k9�4���r^��G^�U5������'��oFo�����!��I޹�ALԮ�y��[�7rRVbw7wS,p�o)(��������nK����ބU�9�C_q�=z��C�h	��K�B^\��-�6r�VON��uٺ!yvקܦRu�1�d]`爧Q�&�_8��s	�k�H.͑���ˤF�LNt_en=�Q�8��sŹ���D���N�E'L|����s�.�Zj���0mvW�����,{�gZ%��Z�-ً(B5�;�!3٩O��wGt�Qi���,it�~g�ч��&��L��6{���\:�d�8�1���"8G6P�I�ɛ`Z��/��VGs��x��-�����x��Ur�Z��r�B5�O�tz�Z�ڷ��Z�X�c	�(���p�E\����5n�T�O`R�i�wL��L�l�����<;���,��^�W�,����w�u�1B3��ߙG?�2�O�ܘ�c��\ņv2g�`<��5ft C'ޮi��Պe���d�Y��o���c�C���\b�'DS��%z]_��w�E�tE?Jk��s�F�
!!�\<��;^�Kx�|����\��Š<z��@<�R�~?O�|=��9x��Ĵ�����Ԥ{�L�Q�u ���,=!ߛә��*�m��t����ﵼ02n��Vx$\�qX��BR�6ӭ�9^��f�=u��I�Sr�P�j��E_<��}$Ѣ��W��L�ϐ�4|��hC�W��_bdQ��Λ��ka��\K>��C3�2ND�^=��ݚ1��i��,
W ���-�]d>.�x��ܪ��\��:��.�)�j�;�����9󧔽bT�r�{&���w!���6w����9�E���s���x���j;A�ٳ��cռ*�H�|-�2.���V0I��r3j*WE�z����ή�^$�Z�� ɱb�O~�Ӭ+ǣ1���x�
N�\��9Ww-9p�w�޴0�VL����C�N+�K"���%&SW����t�On�$f�$��Q�yL��X�<S�f�wpѬ
�!	e���9w��	j�R�����Y�ʶWZ��u�f�D�If�ѩW��qCo�:a�rvx2��m�N�L�I��Rr�sȣ�Y�7[��t�W,aL���?�|�Â�Ȅ�S{՝R�^�¥�="̦�}���:2��>�j�;/|�y���;�M0���������s���e�Q-��p�I��;/bj��9��lfr���^(,��e�~�Mn�y�ݱ흁����p쟍�=�;`��h�&F��w̆V�0/L߄7s�3qԞ�ܕ�W;]��)�����(iźJ�'�_��n���U��ĹO�"_���Il~�}Y$�(cd<�Y{AWv����[��t�@�6"�v�ų����qer웕	ٰ��W�ϵ�k�0�:�-i5'sf�t��f���-�A5�v4�O̴���)O�6Nj����AC�q�?~C�WvѦu�9�>�	�Їkt������q�VJa��5�=�E�>�2�͠�`H���!`ޖ��Om��}���B�< �i��^�چO��hGVI��Fi�x��+��4�2�3V�	ݍ����~e�{��<!��0(,���ڑ�����8hM3Eؐ�X�x��~����O���_�Gγ��<"]� �E�5��N��S�nho>��/�[���/^��(��LӦ3��	N2@r2� [�Zz�o`K��{a�ql��Vӡ.'���^3.�՛KƐ��Ka �BX��ALgY�6q��l�����������ĜSm��*)s����0(.�V����e�ϟ�B����A=,�,R��}1��ՕgJ霭i5{���+�<C���\e	��i�dݳ��n���Rt�H�UQaL��m.3^�B9�]��vmkT�C�{g���C��5ИI���e��殈L��xNw�흧8愷4��f^��؏c/���\yk�դ�3!�J��7/o�+�:�J���8���B���&��.2�!m�=�	e���Zv��p
[[��*���a�K^�Heƃ�z)�3��Wt́Ҧ���q���^��"5KG(d�s�26Q�2K��)ږ�Ы��$�!� ���?�_B|ވ��~��5�uޣ[/xb�9�Gl���1W�"�Œ&A}��>w�xa;�  �c;��zA�m����ٸ릑y�+i�3qb�F�<��)=#��� �-+�������f�~|���k��%��E�L�Xǝ��ᷝzv)?\�Хxi0��+��\��eIc^GjJxwf��|{WEE�)��m�A�v�jb�m/S�\�ě�fÙ8��gG1�ְ���>��
�6�+f�^������1��q��)`�8.����ʹq�o�`B��:�t�{J	{m�6�R�VĶ�n���8�z���_�������%ᯌ,��[Q�ol��Q��tc�ʞ��g���Wջ>�p��-R��@��^�9����z��L!�6߬eK2N���_1lXr�k:���K�9ӬQ%ڸ˷c��i:"ϫ�����~bO�<�7�x[�U�jgJ��l{��r[{7��^=��L�CׂPn]��-�tM�1���*�ߏں��Υ�3ߌW�nM�P<z�;M2h����ük)J�$C2�v-���p��Le!iJra���,_uޛ��ltksv�o��m����B�e�V5��#b�k������.[��#�]v�ͨ�$υ�2�7�QІ�-�W�Δ�Mō8�Ñي��V�w��<Y7�})�+7�k������c���C�O����aߩg]C�|LE����E���]����g!��Xr\L]���Ʈ�9R���!k�;2��B���3��1��@��sG+.3�$\�5ڡV<�p5�m�Ͽl���������M��E3���6Mh���3ۈCJM
�=�,�f>�z���Ol�@Ųa}��$':�CD��z�CJ�Br�o7!G]��.d�'Xߓħ6
��5B*��E��e�'�|w��2A�r�`�swr��k�V�ta�"���^��):�1,���L�%I�k�8ǻ�OC_I�ٚ9���_�ݪ�C�(/��n��*s�o��+���������n�cY�6}���y,٦���F��uփ;��(fM"4G7W��&8jD��I�Q�=/I�>� �,^�!g4;��c�4�oW+��B�K�������k?���E�ɛ`Z���w�Q�S/��)�_D�f�ګ}����H�����*A�Ƈ�=#����]Bl���Ije^!�D�j��%��}����XɯA�d�y�{����_��|���Q��@s/�X�YF/<���b��ES�u�������Ġ��Y�u�3=2Fg1uur��nu�ݭ�^r�����`����T0�Xֳ�YV�Z�h�l>r�2Ӝ���X���װ
�^��?6�]K6׺-����p�G���E��ORl�a�,�?]�m.�)���I�������qɈ��w%������g:f��ε����64>����8�^�����l��Cm�E��Ǥ���:�q���L[�;��G{Kݛ���6ꧭC��G�9.'�=6^����Ksr��D��ӭ:�R&��1Y�f'��k�J��$ߥ���#m��:�nm�|L�rj��2z���Gwvh>y� ��;�vZ�<���rk�==^���)ˍ͉���2��7�Y�q�KR:���SsN�e�X7k�ᗬ�޶�O���D�fs�Z�ޞ�]��$�;x��d�ә�d�x���v4ɷ."�X#H�l�B��xM���C��E)T�ɫ��Y	h��^��K���gA�;�eyg�W*�|D��G:KG<.¥pH�=s�x�X���]s�y�v�C��f}��P̡��+շ^N�V-�My�nN�2J�~���A{���*�!]S��.9Vm���7q���2�x����y��$������GX�8m�}�Gd��o_}�yƮ�;���Xv�D���&� �&��HA��+F;�^ݢ0;�l��B��z��ۻ�F�CW�S��|��Hu��7����=�).�O�^"��^X�����7��?S��1��lB��[�r�68��:�.'2w7"��Pzs��~�[ν�UI��,ǘ-b7�F���\'���UǶ:���q=�U�'�A��k�w.��.�F�dy�a�9!ߩţ{q2��ס����c$�{eQ���P����Y�SF�yUxF0�a�Q���ܖ�飖�pb�����G7dޚT䮠�VPG���j8���׹�s�x˵d����#�X�qù���+K᲏и����B�[@����
���&*�?l���W�*e��FY՛�Iԯ����0�'FN�w��5���n᩾����I<�㢌����C: h����Ed����#q�)�wu�oFj^�8"I<%+"t�E,�^�26Y��b[�큎�c�CЩe[�ڴ�d����c ���3��]G������.�qf��W_j1R;�%�B_��E��;._���^�ex����̎WǟA�RqSb'�[*&��Ґ�k[� $��܎]��ĮsE;�����/�:ə�	�$5̑ ��ÿ�&��߫�^H*Ȑ�i�婵n�����~��9,e�d�sQ��D��c�B�D�*�L\��-��A�mI�%��z�غMP�9���7�g+�u�����A��� ����hd��΂���Q�H1s={�~8�Qv"��<��뵨Y����Ϫ���n��o��[#\��Lo^�^��݇Mu�m���L��Q�k��l���g[w���.}B��A֨{vx�-B�6�2��lf�gs�1H�noI�����R�w �G��٪�q#��U`����KP㚧�Z- ܥ4��e���;=-�����:���v�[�oM������a�:�)VW<���F��Gv:N�Ü��|��T�Z�V��̗&�Խ�0M���pGO*j�����W�w��wT>ʛ�7�����2�{9�p�O���
2#Om�J�+�e� ~�o����z���o�����{}��/h�n^^�x������ܬ�yP;s���`1m;��,R0c-"���F���g4|O]^�=�I�N˴��gc�m�t�`��F�C+�ʒĩ�^����_��_�=˧u�Egq��ʷ�O;,>����ч���f���1��[���6U��K�j]J��]ܛ�r����NH`#���}��>�o�n�!�h�>~���"912�T���t�.�e�Ñ�M�zx��!ڶdXh��W��zӝ��f��nJ���
�e���k�B���7[KRmnM�m���W��z�4S��׵���5��TDmr�e˜��*�s�Շ�z̹��e6�H�-�k�yP�����G0��2��E��-��&�o�-9��t=�$د�AA�;�ND�[&�6���]�����q�4Ҕ�{d���v�n�)�2�n�:�c�Ǯ�Yu�P��[��M��ɅT
�&x�+������I;k����7�����2w�uqB��}�2<8�n��|�Y��m����qa�a>�hF��h��v�Dԫ��f��;���A�rQ>��S����]�+R��(�!�]��c��W���-xt��������C��ugm�0����R�㙛W;�7��7~+�u�w�
\���
�7�Q�-�1� ]ȫ�<�9M�X�uز�D$<���t��	ĺ�3c�f^�d��V��'ͨ��*���GG���KUq�f��&�3�wݍ>A�ã ��F��������Z��͎�F�:������� h���/�{�0'�s9Kz�1kڨe xe�𭘻�e�����g9Y2&j�S����.\d����עR],_`���l�)֛9���f�S�z��/q�N�W��L*�3�R�T��v�|^�1܈�ҫ�w2��K�є�M.��b��c�-�Y-��W:)����cuZ�I(�J�ai�A�¨����3�0���Զ���Һ�IB�%��ӓ��'K��D���9i���YgeLXf��7nGu����q6�G�\̲�m�AI-W�se�A�.�XG{n-5������(K�ғ��fQ�SV���u*�с�!��0F���S����gH���ٽ��!��� ���rW���H4����Y&�Z݅�%��R��I���-/U��#�x	�l����"�5j���o�r��h޸���Z�T7}WɢK��=�Z�}#�O!�p��k�ޮ��7%<�0־�ѾQ�em�LBm`��ss6�����)���nff��X(��W�dj��@��I�ю[�[�P�-@�>��h�T����Y�@7�{��J����6�TzA|�R����X�
w}�s�>4�4�ͺ]@�L���pQ�G�v��]�L�٦ukarU`Nt"N�փ�nsõ�p��:�����栭=ej��f;��홸��})�7N�*9�`�j2�/[�VP;�QDf�D"@ɦ0AI4wgt �WM����˺�wvi32fb�5�$��	C﹍���s&�wt�ɝ�&Df'8�svN��� �����	�d��]u�E/y���
�R#L�	M�\�y�2"�A��^NE';9�&�b�E�pB�H�9�';��&QFe��0)`HHs���2�Lɗ���� h�p��y�A����b��P@fbx�nt���K��$��H&�gw)��t��_̤�'+�
d�`ľr�b3����4(��B����^}� &>���4=���MdR޼�:̲)t���|E�!㙝����e���N�x�qΚ�U�����BН����wVt[�f�Q�рz�Ϻ�t�h�!��#9-�Y#p�"���4�����у�(�Z.@ލ�Tt�b]��l���%�	��zo��Fg:s���ױ}|��[ky��
�4�]� b��l�қ���0�i��^(���]����N�D���\�゗<�����5�m���P��v]��46+�X��J<�d�M]vnh{���"�"F�M�GY,��kI�˾�흍��*)�zYǬj�5����l�楫;�PZ�-���ƭ3���v�{�t�:ӛjni̍�p����8H[�VLtK5��i��Q����ݼ#;��B죷u�j�u�FT2Be]V�Wjf��vѬ�"��u��:|]�Þq)B*���}��uV��tz��;�Vz�m��n�Ǳ.�2l`�����x��&I%6�c]:<L���k���q�'�S����a�ݭ�tV;�]9wmJ�AyƜP���Vw{H ������:�����/������m̫!m��96�#r��阩��n�Iv���fJj��و87e^�����챂��.��;)����!٫\W&��ه�0d�^� Ȳ!M�:�~)\:�g>޿g�m�q��w^��@M��d ��o"�jN�M2mlQ�����(J���?���kn�w��ߋ�:�-�7�-�?��+#��NV�而CD;�(�;�p�ɝ�����&����yS�`�3���zcgV"���V����ͥ��w�u��|�Er�"jkҶ����w��9��LlS����d��3ƛ�z5�H�Tk�Q�vn�ҧ('l4��౦dt��Oe���0�}����=�`�x�ѵ��M6��^�ݒN$�����D���[5\;b��b��f�x�������>��dY�|}��tF]�]�}:)'���C? �B�6�G^Q���D�B��:sK�i5�f�vT�	�If��W�6�}R�c�<�Q结^����x�03D=�7O����('e�N�U�s��p�m�w��[~�T��}Z<�òy�{��e�p~���8B�4R<Q�h��z_rhk�/��:���ӕAq�t���ts+mL�,iJ܊����њ����WW{�&�;�-��M�.7X/ef\�G6I���:tp� ��8�3mH4�vY�`�z�7Y)�;�Q��_�f���㣡����.v�����{�-�Q
U�5�qQ�ɹ�2����K��F؜��Է���z���W1�!v�7g]�B<
R�)�ު�\���ٖ{2�E��1t�~A
��l�L�?
�C��_ �F�G@��0�YuqM�3��X���gW5uA�>ِ�OӪ^t���Y|
���<�jYS�9�ю���g:���y���Q�#1�t��Do������gD� �Wx�v/9���'J	��o>��Ry�0-��oJ��Sw��m�z3T�O꜡g���<���h��]��0q��o&&a�����\�t�(��t�Ҩ�79�-�����P�����t�u%�;s$��H�y��ݒ/M&�]�1յ�{�l}�|�����$p�����m��ow���勹�0�����o(Gg8R�]1v���j+�9��N	�
��s������JЕ��n����צ-J΢kp��HiYN��9r8;@0��4��A�wH2��x4��}+M
K [��;�_�;/��w*��;�J�5�-d#�ᡲ��}�e�=*�7[$��'�U�V��Uww5��I�]#�2���9��/*���X�`;z6.���7?rܸ��p��[��p�?z\�=/ʏ�L��K���H7X�"��}@���۷���Tz�Љ�<�4�w�,��Nse�������2y۪�r5�	%�:�7'3cdv�	�d%��yjm[�x��~f��=9����'�����R���L\�!m��mI�%��� >s��܊j�x#W]n���p`5���{��9^�%3>��!w1
���M]�=`ܴ�5�eY�['�ft�*��藡4΁�PEϡ!�+V�dH��Ȯ}��Mz%�$�k�]�n��ȼoQIH8��[��fHYa�1�-WaC-I1̛���RsH!�%���"��T�L�V�U9�f8@��YCs�����Y-y"���O��>�xn6�����8�ﴘ�M��{���O@���M��l��&5�uE��6�i�o�=]1Q�qU�f=�G6�Rk\;�d�������ZFpclu������s�cw(͗�O���
+��T��8>������-��őת�M�*]+��t�i}�vzXe���Ԣ��M����>��O���r�OP�Ux��t�%�>:]Z�~�M��cu���mnnm.k��MpÝ�d]�Q��ʠћ=u@o.T��8a�V趶�s�����J��K
�y�l�⺽Z�gU�J�S&��g"`ƴ��oi�Vcs�ϸ�R�]�lG��tqC�y�3��뻐g2.�7��6cuoNӢow�إ�.w�{6�8�|�=\3�ʗ۳9�i��"�l���d
������s�#�Oi�8:G4[,f�Wo*�#�j��@�����XO{y�/,��I"RHO.h8*��zಓ�Eѫ1;:����h�!j zJDm]u����"$u��l��3-tö3���8����
�2��F�P��J�K����φ$V�G��]�l�Y�%�/#[�1I�V��I�ڿ�%���!�V�ċ���=�ٕ���9�L���;�2��ΛyV72����.s�-SK�ع��.�6]�v�n��u7)��nV��]jښ��pL���	����=w����Ln�Нн����m����lyY�N'�"��.���]V�{a�A*rp;����E0�e��f���ή�><Fa)#�Juמ;wQ.f����%`�{�>���5wW4����.���\�H��<�)��]C�I�R�U�L�M4�L���znk�ަ�����5�Uz�![��IXc�)$��Ϸ��Kǿu���-6d����s�Q�SUGWm;�H�z�h�J�ic�UȖg&?`�	���O��{�u�
���G�����,���םrhYM �ت�x~mn�z�w<v��#{�"�⌮/Ҍ� u�<���i�l�*����ylms����}گ^�gFgVw��o:4��k�Ƙ?����s�p��d����aJ�-��.�yV�`� ��֔��D�Д��r2����+{Y����sr���'Y��"5�'׽F���݆�)�9D�I�:Cl��ʃ�����y���*�^d��4�/p�:v1ng�����%f�}�Œe�X9���Fk���0F�+�*������4g�UqmʃU�r�8����R�op�rghMU�3B�J��<�^D�;�}MjCJ S���4�U{o$��B�n� .��S��;���
�� ?Y��{&��ϳ��z�n�c�����O"����g'�8�"�3�vT{0��]����b@�H�q�0:�5��:�<fQ�͵��v
R6)�; ����G^Q�JN1s�}|̣P{3�w�A��#Bq�W�r->���.��-`����T�TV�����[n��w6�Tof�(%$'���Ҥ���ڛaN�En�7p7�.��m�B�����9^���ڊ��׹ �+��w̛�r�C���*��:[��w���p�s��Sp�u�+�#�)T����57��>L;�=^ˮ��;7����U���b)�X8p�PY�#Pg������J���2s�ư���*��e?T�2��E�A���Z9H�7�jM��׿�����/cfj���z.��3�k �A;[�!l��� w���V���������d=N�����M=��=~&��=��,�:F����^=�1��b��p��w-N:5~U��g���]C��t� ]�֙�'w��Q�A�oZ*�3���9#B����\�ޗ������k��&<�ަ��~Ύ�ީ������b(��B��/�s_%d��n���{2��D�!���A�s�1!+Y���G�\��H�]�?v/ �7v5ϤhF:����}�1�
0�5z��r��&�<4�*�ztӅ��je/s4��Q}۹�w01�R	X
2#�&�ҧ%u �VW���S[�!�9盟��#s��ƃ�|� ��Υ�/:��(�V��p�36w7��Y�ޔ�n�GH;FGPc��@�2�c$�SŲo���7YL]�S�k�&VF�˼��e?d��w�eO�O4gƘ��g� `�@
��x�M��b߭��*���DH�	�~�ϯ>~]�4y:���3�qKnM�����7��E(z��5ux�V�@�VD��E\��yy��7]�q]f��_E��s0ˆ=�꧀��=C&.B䶀� �6���e��^x����Os&+y�B�%Z�(*Ǜ�؏���U�wyŌ)��\��!Ve�ڱY��o�r����#��w��*�z���������o͚nּ��t����p���5���h�qY��Rj�ܓ�5�>eݗ�b�q��N�}X���A����1�JS��^M�^������z���Y�ŷ��WO9�tPw��I��~����=�)ߡ�kϑ�Tv� y9b�
2jl���2)��6L�ޓ1�u��G���3�Q(���[��=ّ!d:B󦟺����eh���Ѹ9_G����rEsAԉ���`*��c�9�����&ʱӒA3B�/G�;��P�YM�*]+��]��@;=WV�˻g�_����ܗް�0�R�;���f���*�qtR�:
�m}�Ս#eǢ=��̘ܖ&�߫r�zZ˨.�����B6J�4dY>9w�(�Ig:v�6;�	�X��m���T��T���u0q����������8褃h�d���s���{�cw��;�^��J�tyt��n����gm,៝�+uwJ���~��;��0�k̺oK�{z6}�lѰ�<G���;H��#���32F�y�5���{��W�w�Q�����m�ͫ��3���سB]���vi��3���u�Ѷ$yV�^��j�TwP��39�95���3��|u������ȓ����b]�Ԗ�v���,�=uCy�{���f����%	_�|3M�i��Z�׸��-�#�@���6�{.G5i��uRm���;��iW�/��輳�$��I	�ͦ&(�c���q���^�ׁ�a������,Ǟ��ں���^�a����vO����f���=G�>��}Ħ�yj@见��C� !({�40�4�9t��G���:Ù���8�G��wt�%�3m\K��%�!OA���؇tvә�ѷw�p�kw:O���PҒ�,R�d����s>�gh�哃5��L'kù�FR��np�|zG:
F���8��B*���e��ѕ�p�6�:^�3n'��`�´fr�W V����0�ƱQ�IDL3��$ba�r�WU��9��Yy�����pEC���;�H�QM v�*�+��P��n":1�eo^[v��׳gvA���d�)�� n'њ�:���=c����������=��g����{�|ވ��;a�6�߮Nӵ��e0�#C�7y5���W��K��v���v�.��5\�k�k�
�(�Wp�*@JIN��\+���-��w>T��Ǐ5�IqW"���1�]�F*-2�<��r��7h�}r��%c�W��]�-M�ťn�+v�٢�Յ�.�0���'9������Z���X��DeL�d�e;u�Le[ ����G��
XP�h�|�y�u�5u�H�;��5:��H��Jr+)�l�	���.�n�rƝΣcfGǷ�S!��by>�{�@����-��A^b2�I�	g��meJzF��c�G_!ê�LR�[9۶ĳY���'��;�y��f�Ɔ��)�7e)6I}�F�<�K�ZCvF��"�r�c2�B�֊�G`�����WRյ���
�M���$��2�Lc0͋&�K��S�r+J���4�U�0����wF�����4^�ݦgqQbQ^Bz!fc���h���z��k� 1(�Yk���Ѕ7����wR�Du]i��ޓ��t]tAd�b�����Cvs���彔T۽��R�"Y��4�������	�N�}zk�e�Q�[lp���#�:��T�C�ja��Yl)�C�`�B��c�zU�R��%h3�3u�G-$B9́jj��Y\�/ym2ueMc9)��Y@\��tb�e���#�Ё<�Xr-v:�f��)��JxJV����w2j�of;�U�Ί����)K�bU�YD�2�vwn@Q�ܪuL>Y�-��-e�Q� ��/b�Nͥ�X�{��50�9�TXhl��SkU`�6��A�Q�Pmm��[�HWZ���'	ܛ]*�}G���6�|a���j1;ɔq�/�aj�E�ef4���C�˵ �j+�y�"ǒ�=E��'��:<�Gyi�|Y3P]�~�燣,�]�:��ME�:���Zq�gs�I�i�A���tJ�3��8)��A ;��x��W 8�����25Nܜ��(E7s�����w�ҁ�/a�j�����'��`|�f�Q���zj�����Xq�2�ʹ��&�l�е��/�T��I�YO�4���nC�9t��Y�I�_ a�2��-;����F�8�c�GRs��^f�%-�;3����Fgr����y�LQ�*9�Ơ�QT��
(N};9��9�0�Z;W[Q���T���5}�C�R+��5�+����oիh����ޕ�����4m��'���u+��Q3��{�(��#�=����R��Vh������[���]>N�Ap�V'�î�,>744pYܷ���`��O=��	�E�{Q�@[\�+�X�%D�/Pb�-�і��p�K�u���md勤���m��lu�84)���5V�Tz�v{v@v�E[4��`�����l����{�)�ݺ�K�A3jm�Ї9�jV�P�,�䊠�r�X^�4����_J�Q��J"
7I�w|�||�����w?��`�Ez��$"l���.�3 ��ɮWf̊�wp���e�먡(��H�(���Ⴛ����,wuΞwTID��HSI��6�'9`$�w���G74�w2bG��v�Dɜ� �W
#�9��\�S.�vB�4�`4�]�<��4��v0n\Ė2Jy�h��.��]H !��\�nd�;�(�X�4�H�"W5������ٚ�<�BSs��BnnQde$3,9ғλ�@��<th�4�h � �r�Hѯ;���(�]���vDd���h�;��Te�v&9��H&��t�I�bRl.n1�%2i+�����Ȏ�$�uvR��	d�\�6I%�.�%i���C�3�ۮ��o��q>�C��p�r0%�W�]m���9���|����q���[�\�$U�1�h-����b�;B��(��U�;7��=�?�֕h�!q~F�㭾���l��i�猦T���Oa��Ξ�Eݕ@�^U�D����Iv�n6������RR@֦�D9��a�d���= ?u�����[�n�S�0.v��F��#O��w��}�%�i^g�u/}���_�[o}{ԩ���n��NQ1�hř��"��3��ݛb����z�'ѭB�0�fFHY7��o���9q�x�gY|�衻�Ee���b|�ss����Ҩ6û�;��cxVh�J���}f3y�K�˅��Tٺ��g�[�J��O��XCf	�����}���g�X^Q�#��׵���%�r-����S���c���̞�4-��3�}�O��|�"T�a��8��ֆ���Z<��ͥR�vY�}.GwNm�&d�aZ�����PU�Pɍ���$���w����v<\X��Y���	����8J�[?����s�Þ����.����(��o	gk����v��R7���[1,<3��8]Kߕ�5B�����MULN�N�gf�\%���G�cu
4zi:&x�L�cD��������D���B�����{&�^wToe�W^�t���V�ڤ\-���T9J4R�Wow�̴u�ݘ=��XEu\�
�3V��"�C��G�F|ڑ��£Z�����E�+{rf{���Q�QUA�����i@"�ΐ��
�r��Ȏ5Yu�Sض3y�3���'^�]D�47��ǿh�Ab��Z^����xEFa1��Ftl�-QQ�W"}Y��;%w7z��֗0��)��F���C�*Dl�U��S5�^A���+�v>�-�붅�Oc�ѕ�2cV�J�������lꮓF���W���w��ic0��2�`&��O��HgџT��y��7�8���ـ^�U�%uZ��)w8�W=<�����h�'�l��0�� ��#��1�x>�����3]O�w����$�vO�;G�1��q����W���_g����MOumz��%s����*�x��%WR\����J���]Q�o�6L�����'K�n���J�Fg
<�[��&�KB������c���p��R.�X�0��W�X�ͮK�T�W�:)CJ9�"Ki9���G�oB�����^�\8�5����f�*7�{�UO�3��e�f�i�y��7��2�4�e=7�}����E<=�18�x�7xo5E�7�		u��Z��r��*g�l�'�Q�i�l�>& h*��蚺�xvBԁ��G�%YWu�n��<6T�pams�{3N���q��A�X�⚪; ��hdŮ+:��/�Ǧn�H��4w�kh�ܫ��c��D��,�� �߄ �Ѭ���7J�6�x����8���L�`�ΉzL�NE�$,q7/SW[/"�Y���w5�M���|r�y�H������Mr�n[��̐���Lh�kQ/.Tf�lT���Y���z��t"m�"���&[+EK�"*���%\�[9��@����ٍ~|�]���r�.�\c^��./�&:F�U�-�N����tz�a$#X����#"�OW������R/���g ���e�Ԝ��hؗ��]�޾�n��umX���YܵQ�U��k)��<��+u8�P�N8����֭̴�O��|Dۖ/�ף�P��#�����x�J׬0sq2�oe�Fu@�eL���!���؂��К8\<"<%��{��d��{������]1u��sq������:r���l��sH�P���F�J\���u]n{���	h�s�jie�1��SA����T��5�����szOu+����6z��ӣ���ƽE0�s-���E��K<.��r��(��y�M״���l��f��0Gw��+��5�4��31�5ۻ��J���x&�l�\t2D��u��;��W6�n���ڢ9k���m@��ѡx�����bt�%$�f7B�L�{Ւ�tO5v3z0I�_$L��Jc�iLu]m��W/z���� )Z�1-�=�[8��{�ܚ�<��3��r	X{�5��c�lӈ��:o�U�oV�U�?��Z�WK��k�X.i̍�!N("��uۅ��&���e�z��g��&#8���<�R�J��O��<tq�޳��~9'��!=�G�X0�Q�9הv�B�oY�"fP��^h��&�Bҷ[p����s�����:]Z{r�+�#a��tP��Y���~<�)�:�1R��+d-$7�1)�]In���l&�&;�޲l���}\�5Su�Ses�7�Y[��壣,jޜ��k
%����9��:[k�P�"T�֍"+������:
F�]ĤD"���vLӗ{馛��G^�r�)���x
�0�S�"������0�(-�9�D�<m�>I��]p���O���k��rVקx)���QM�VT[����m�q?-���M�~��Q��ݶ:��̛�0���Lf�Ψ-F͇�ܦ3�3��f���6�\MVD�;��S.u���X�1�B������.���l���[S��[^�r��/*�A;��k���lC\u����5�.Y�4`~8,:N-'�僦L�u�Җג&��qtR}��C�%'��{���w���8	�e�	L&r��n�m�r���&;+d�auz[E�;�['M���CTL�s9�}�>�$��|���:�5��E�{[����G���
A�]#�6�@w`E�Q�F�T3[@>B*R��
�mX؆9x��+.)�m�v��͇k3Nm�%�����Ҙ�I�^�6��g�����L�
��nfm!�!������n�u�����+�9�`�C����1���vC��V�-��ff��~@"+k���si�Ǯޢ����o��v�wyBp�I�iց�(��?NC:�B�<��;��h�ȧ�����ϫ6����tDO��K�r-u��=�K�љSI���H|'��ca`bы�nj�н������6�$u����.��Q��K��e�Xމ_{(�t��I��XU��&6}�B��$Ҏ'if魧g46�c�]�u�u���"��&��!\�\#˵[��t
�R�g��*����7Z�}#��^>'�y���
��d'"��誽 _#���������M�᝹�O<gWJ�ESl��R4��t�>pE�2$N�loY�4p����$Z���.45����{�c��nB�&���+�|�j{�B]qf�#��9\Z<+�Q�T{�O���4w�R\��f;^��^W&�����Y�f��}+�ꞡ|�Erדi���c��wJ�5沢U�۸���.��E[�����uw=�޶�vX��K�ĕ;��L��O�5s��
������b�gk��6���N�u*s���;���t4���y*�'���V�Ƿ���9�2��n��q[�P���qo^<�ֻ) Dʋf�c���D��
�X��z�<�0>^]@9�"6uP�4X�����)�ޚ� ��"N�m�}=U�6E%L��f���ݗ�V�9+���
2�þ���,�5f7:l�q�T�I������B�؍���d]���v�<ҡ�N�n��~ ��W���ݒ�hϺ���F{��[ރ��l���ٜ��x���l��$o6��A�G���!��T>!��G#���P��{ <-���l��DN���q�ܲ�Ad��^��b=�yU�G^=A��)@{�j&��jԁ�qUO4�UhZ��g�69=4X,�],�qAt���"l�����.�^mݤ�}0�-�����~����֓�Ok�Y�
�X� ;�����VH��=�b2:�qGNmwv�p�D��plɯ�T����i�=�����燍���p�+:���M߱�r�f�P�6a����#+��:�3��C� ����)���+;�h�X�n��߾����LF��xC޶Z�IOUK|l�GN������-vv.)Y��m#n�7�[iS�^]nF�Q�G��y���<5��<�@L�.��\��p����K�~���E�% ���R7-���*59��b�Rn����]A���B7B�g��v�&�ܑW�*R&CeotD�:<]�����GTӤ(�d<x��GM�B�h7).�čt�)Q<�ǣ7gW5u<��3.2
}	l����E����Rmg�y��fF�|Պ߲t��Q�<w�'a�v6Cv	�V���N\,i�7��^ә�箼1�M�ܩgq�U�*�g��78oCvo�X��`�(�C�M�3�ŅJ���r5j��R�+�t��n����6����O2�GpmXˋ��2���˦�3�oF׫݇a���s�F��ш<*4��^�Yn���kz*���5�r*��ź� ��NE����pnxS�m�����x�:	�p�/
��f��n�^Y�I!Ǐ���8�k��5~�D"��>�\[�*Ŵ5Yv��+��>�^�O��e[�R�;�\t�{J�n�#s��lY5�n�g`�'�ق[�1m+��u}p�E����d����5󚞱r�\����|m�t�:&�ٍn��je�e�ms�Y9�:^k3J���$AL�����{��w�k����kC��b#�0��Ƹ���ݧy�.���<9��~ܵ�"�t�dN�MyK:;�	a/,ǐ�{� 3�l{��;�-��s�y�;�>�R��:�WK�i��>��3���^�|l�*p�e�õ�A�;q��g&#��,���f�FĞ����M?_��~�ɡ��+�;8�?O�o�5����s!!�D��t�j��8��B*��н/u��=y�r�&[��@W[�då\��2zRK�L���W�j�y��t��I�׊`}gy7Q��N�XT"<�Jٝ��P(��w��&���8���=�O}9�Ԑk���)gf�m�-� ��������8�v������*(}eʑ\��U>�UǺN��e��[`0��)5���Nl"'_��=�������s;˞M��ɵ�Xn3z�u���4[չl��y�ݭ��yu��wp|;�;Y�
sQs�F���VPY���R�n��©����8��ױ�y�J������ڟAH罣,��Ȗ��Ǵ�L�ۚ��h��(��*����u�諕��&_�Sޱã�X�v�b]M�B�t�M��z��h�qRo��&j�Κ�L���״��䉩�f`Y۲3e���ή�y9��r��	��1�@f~�BP�R����W�MV�n½��g^x���OD�%LO�6`���Vx����:G��Fl��/K����Kmy���9Iǡk�?����O:>U6�������xVj7����x�b�{s3qw=�q��PR#G1�:��(��?O��+���-OҎ�q��Ş��(�^��]c9�WHD�;�W��'�j�W�Ndd��aqs�Tm��Z��$S�U���3RCz���iPH�O�mS[k��w�{G,���2����=ܪ�*�Ll���$�J;�ƾ���`wʻ�i��5u�^��>�qQ�(1�?]�<!v�u���[B�#2q�"(+�7.�:$�&z����W��M[8��Tâ�^� �w����yx�{=��g����y{��+�z�� �[��p/<T"�1����켥}2>�A��V�v��s���1����j�a�X�N�j�����J��u�[��d�FIm���|zFvt�gV��p�4S9RpsD`P�i��m��;&m�0IK��\�՗3�so(eX��4�c�n�l!�N9QT�	!�Vi�n��{��b��|�yoFV�9nA:��j9b�Y(�+Lƺ�$:SGT�T���3Ug)���5j�Fӵ�̱��]/5�����&5��o�3���Hd���c�9q+��\�%lpͱj�Oi��׭3:�6�t}����}�^Ma��6s.XQ��,��cv�@�67{�{�c���3C#u]�P�(���:v�܊�gS��jJ���8�K�ԭS�6�ҚZ���x.��י��\�>�U��%.Qó.��R=��ڹ���%�kzA����4�6�xF-HZ�.�i��rjO���n�Y5�V�5�y��% $��BK9u]��s��Э�v&��*���.oh��o�~���?3 _]��hǩ�P�7�&�xT�d,�'U��
����3�9]�Z.[�X\h���y��,�L�zE�Y��V,�7���%�N5����]���	;��I�]�e��0Ҿ|u9|�L+
ѳ�[�'�;��M^�aY��t�zG#\qj��Biѻc3B"A�y1� �M�x� ��3H���P��T��}\e	Қ����gr̖��P.�N�|D���.:g,
f�j��g<�x��y�eG��p=���'h��]�gy�%\�t4��d��J/�mAԴ����ʋ��������ǯ�Mb]���q��0�'�to�v��/Z�Ϧ��A�fཡY�fm)A���l�5�ѱp:�N�.���[ז�\�41N������b�hu.a��	�&e���Y��p�3i�8~�P΄���'%���##�T�R��5���{Kw&�N�q>b���ٟމ�\kzV�n7��z�OE)����'�9��*d��A��n�C��lջZ:�&
up^3�{�;����7�0͸�#�@�B�[�
���fY�-WfGP�m��e�x���kRe�S��u�9s[�tҾ�;U+?K����8���EkAC�µ{S�eH�C�P;��*�aR�Mܬ����T��x��;��Xp�:䲮mv���/r�hK���v��sES��<x��@O}�D��v�;���j!�:
=w��,���f̩4_-�l!M�+>�q�֍��46��w��ce�H�+;r����A�E�����-͚�vrdSM�qwsU��״��7ۜ��]�4E�։��vm�WC��`@;͈�3�ɭ]��e,Y5�����=�-��",����&K��fC��{�q��N���L2���L=+�r����N��T��zv�`W�����q &O��K��"����IJ0�L���n��2$II��"k�rLZ�sb�����]��t1B�ȉI�F]�	b��9ȃ���-�;@��$���n��7���&Z&��vk���B7wTE!����Q�y�Dm�Qd1Ad�.��c@�����])(2k����H��i8sy�	��"�w��xܦ'�v�"�wt�F�cDW�fb��WI�p4wv+�wF�㮇]�j��I���+��#���GwI�n�uǗn)s�8�̂"K<�<��K+�����D���/;��o*"񻺮g;�񋆎�J6�I �1�k��,r�oȷ��;������;������LQ�����\ɱs�wU�ݳ��W��d�^uy�A�e��W'�\����y�)�&���+�:���wv<yy��.�:㻦�y�/���v�Cwg\�W�)Qy�]r$�r����=BA�|p�sC�F�<�8���٬�iMW�V��a��'~c�#ޭ��oR��v�gTv]n����j�y����QS�>�{��N���zr�T�ъ�����(�1�:�,B�h��IXn\hk�I<��{�{�gyK=�Y��ѱ�t�p��Z��篠�rh�rW�7��Wϰ�_$vJ�΂'�Pw�2bcr���+�n��F����������&ϓ�
O���P����e8�@S�v�@C6��<dFΪ�4k�NU?~��ɨ 7��\91z7��o�y�z��C$m0�@f�Cz_�+L��+��*_qxFv�����?}W��P���q�è7w�|B��G���]®J�0'����lz�|�87��|OPc��rn���h�=���FƆ����F�"�C��������X��f̍1�y��'�,��f��2ݴ"k��[�/�]p��G��x�כGsL^Y�{�ܒ�˛=�|��]x�&��0�Bn����>ab�pץa��G	�F�E 7�{ɲ�oX��/.Lw�a�ˬ) �\P*���f���շY�%z����ֺ��t��a��_V����ke-<�JU���"ekA�!�'t�q��Nq{�)U�S�j��z��H�s�:�mN��~� ��DFݢ�76/�ԁ8��^��*+2{�[����V�G�N�pCm�����x��\�9�T�6��1�y�{��	:�=�5�X�X��3��Wa�7	P"^yp�s�����D��z���H)�,��䉳A�U@�䎚y��.׆y�M0�*.�G>�M��O��+4G�{u�H��E% ���JF庞ƺ�YVe֋�Ӛ��v<0\1�
�|�\`v]�"��a2D�L>Lm:����Y�3�;�j�`�S����H�#��ʡe46�R�ұ�{I��8�oy���<W�8ݬ{ub��lvᄸ@�n�9�S�/���e���wjܸ+r/���=Y�W�!q{�;��]���z�d��"�ݵ^����]i�ٽ3�<|wn���^Y�eN�W��l��7�0����8m���\������@�u�j��WY��\���樉�
�&�����ΙV��A��9Eq~�J�o�w��s�}z_o	�+5XR	��g�&xj7#��l7����\l�V��jJ��ե+'%*dG2^�{/|j��3�^PWZC/��vnv�ָStJ��ѝ�����u�^ 3�*�ϵj��=ԡv���MѾ����:VV��tӏG;㍄�@�����nr�'�]7��7�g�ٹY��r%�Wf��;\;I�-��9O�������6V�<c���t������kM�W;��xD蝐
���C g�E�xTj2���yfq�.��Ƕ̥}ʧ�l�=�D��hqェ^_�Fs ^��"N�7=�%^]��<�J �ޏ��o�j���ϽdO��k�X:)�a��t{�$]�V���ͅ��5��\�9qrKl�
Uڐ�c^R�sNv�n�!1���r�s�vW
��n<����U영�B�������NݰkSFjd̝��׳��\��{��r�Y'+А��"E���AO�B��R��m��\��M轙��]Q��Dn��x
�#3�0��5�8�����M���G`0:L�#2���~�g��K��d�g�еv9e�

ڼӗF��m�X�@`MV��ѹn?�����Ś4Rh�0�Sn�<�S�wF+s�&�OwV�)h�_�n8��۽gW>(`�'.��?S����jn�آݶ.�*b�gM'|X��)#Y�E3���'�͕��ԍo8"��[Bw��d#�����ۮe�^L�v��1��+*�V9�J����X�ǃ
A	�pX�!���{����MgO*+�nv��kbF�:�$�/�����_W]���}�5Q{������T�{/ ��gW�ivr���W�	�6M��r�8k�Ɍ��"r]��RR&N��WL��~�M���P�Ƅ��e-����Fi��e�9��H��x5���G�>�5I�||�q�,5N��ܽ�Z��v:.N^�[�>oOn�=�T�0g�lGHm���4s:�휀���W������ xa�W�4~q�i8M?ؿ"�'�t�E�Pgp�	�h��Y�3	�`��b)�jN��T��4����0i$qc��y~�����9+��q����GFS��`G9�[B6��?������$r-W*��Ns��;�"e���C�������O��.^���f�E�X�r��*�3${�yz�vg�WU�~��TaIyoz�wǘs�U0��>���k���B�/�v��5��L�0c��Lu�/x9���z�g�GRu�Ýc0��Z��J��w;B楕j�8%�,�����Ѯ.��& h.�����2}�!=ht�*�z���~��٫Z�v��O���)��ކ�A\z�&��`*Ĳs��-���΍�k��Oh�}Ųo���W56�ðg�����Eyh���}p�5��Mٻ�y���Z�������)B০Aʹ��u"���yA0�Т�H�&_ch����n���I�9��qT��U�ڏ�u�� �|wc02��wf��T��i�V�|Z4�J�r�Z��K��=�@l�vOv�dv*
F�F�/��
�����>ɣ�%5ʗ+O�_�^kb��yQ%[�4��v�߾�{��@�9�#euz:����f�k�6��a�����U�3��[�72Х� �mhfߘ�\dFΪ�^V���i�KM�co��f�&�эΒ4���XP��`��#6<F�8(�we{�	�Qf{zh,��P���ș��O�1�P���c��K[�9S���N+�m��r,�2�CV��P���޽NW6���R��y��S��+��ۖ�yk������e�5�jb_��Х֢�8�.��DD������� �����ϰaB\�ݽ�޻����~4j�{������=A�{|�.�EVՈ�f���X�-S֣m{�-�_-�e�;+�u��;Fz�ʐ��k��ț��/�����4.RJ����F28�7�L��E���k�,#=w=�U<(v6T3��D!j<𔍊�lf��DN��!"1�O<;A�=�Y��u��]�D��J-�}��xQk�f%�S��;+R���P�~�訣��o�wdAz�H�o8� Uџj�Re���PI���&�MMTS�n��ܼ5:������� Ԛ	v���Oh,�+�b�\ɐ ����z{]w��n*���!^Hɳ&��o'�4�馑r�̴�9Ӭ��*K4!0�>b���[:�%`�#^))1�]�]�k�1��f�S�x�W��7l#*
C�.}B�/�\_�����c��J��|��F�q��������ʹ˥��X|v�e>l�.�ޕ��uX��Swl��1��;1��;U��*��c�jc�	��|z�_����D�l���AZ��Ԡ(f,��U��\+�q�f���i�C	U싦5�_���n1����Oۍm��p���6S�r�`DRMv��WN�� 5͌��S�����G_!QLM�[�3)��������(�_��W��?y�,3=� V�r~F��e�s��f�5ӧ���^rC����wO��
?� 0�`����{�slI�YUۢ�N�ͪ��E����è򠳸�Z�W{9�������;�j(VS�6u���A��I3�Ŧ��*t�@ի	��P6���B���ty�w܃�e�g���:	F�׋��F_r,�n�����M(���,9-�6.������S�@��`E�/��$%7��Z���$��\zt��k���l��v	�T睴 \h��Q�y(��u��ݾ��3䝶�9�_�������N�JC�6��^_�_3��,�$�a�T��`ف�i�;9�+_Vm�$
�l��HEò�'O&���tS�m��C�<�|�좠&�~U݆�[+����Sz	eЬ���ի3WN��k:�X�f^�^2
r��_8���Ȏ�4ń�wG4|���N��#-X��Y�w�+��U�N��{~S(s��^�L���7�:�/�5V�滽"�hǝoKU�8���D��vJ�r�����9
��'��:���ԅݍ ^Z�\ӝ!���Ĝ�l�{Ք���z<�}$Q�J�c8�x�����}.+gqv�7Tw:6+��S�V���-�d�Wa���΂�P�XE�g��~�s۽��(�m.^��P|����i�YDft�¸���X����6[GA�P��`�mui�Xg��)��T�ѭ�T:+cx(P�ݜ�Q5�$����y��)\W��J�����-��AP�Te�]��ꧺ��S^�3_(a��S@6�4�����j2�u��Mg]��`Ѳ�W�ߖ酦C�Fʪ�������,��;�mq��Q�Z�_Bܸm��zFs���`S�b6uWL�Rԉ���l�L���=}G��*A���|�C���0b3ے/z�9Z�>������om��BX�8�e���w��;��ȊG��n�Kx��h�u�;4�e���tEʙ�EA՗�2ˠ�M��
���y��;:G�V��S�.)�mV��T�1�����j�ܦ��S`���smV��E>��5Z��	[.��$Hlޘ�;��?��������9n���yL���L�慆������]n�ƣ~u���^e�x��/��x�>����g����	�bRm޹jV�w��9�~9vDooVklP���f 1"�e���@�u���+n=��=^TA�����.��הo��tDX���Z�E�
�QݪO^͟F�w�����t�K?�tG�"�����{#RBz��m.h�P������~N��Z���S��Q�U������u�fIS�.8o��s֥�����uI��5���I�����葮:�AU��.Ռ�מ�'��;;#zn緷�����E)G��-���u5l��@
���(�lMسY=w7f�+���EB��Db&�n\h��*�x����G��]B�7��aLL�d�/c�E���4���g>��+BR/�@�)!ˉ��O.=e_�El]N��_V�i�Ŵ�"�lΧ��72�{WC�n��m�d�����[JŘ�	�Ͷ��RX0>��p��Ɔr�W�k,�~�A�]���+8h�����v�gs,�����(��'%p����'^�ݕ��ǵpe�1Nc����Wt��T�R��p�l�ä_B�
���Ȅ�n�lktonf�ނy����Pn�����}��S�|�}\��nڱ�V����1��?yŽ�o�R������}��f��q�FΪ%�E0�CI�*i�nR����Oq�ޞ�T2}��=f�#z���wf�c{f�m�38�5��wZ���3� �����ޑ����򺹨���m��:�zmq��۞�'�u����=A��'�+�pS���ٓ�ߢ�ሁ+��}��s�+��l�/�ka�;��;��M�j�|e�78D��5M��>!D���R6*ѱ�b�ȉ�<1�o���8�z���ov���wv�,�@e��Z+���Q�=�+��ˡ�>Z��F���,�;��������C���T-�ʄ�2Je9V��Q���JH�*���-k[ko���o��ֵ�����������ߋ���ںͬͶf�el�ٕ�+fm�5�-��l�ٕ�-fm�6�*�kf[fV�+fUL�����̶��fmfkfV�*�[fkfV̭��������̵K+fV̭���[2�e�f�elʲ�ٕS+fV̪������fV̭�UL�̪����̪���W�V�*̵��Y�Y��+��٫3Vf��Y��+e�fZ�ՙ�3[3VeY�ٖ�*�5fZ�ՙ�3Vf�f�f�ͫ~;y�o�Z�6�lͶ�2�Z��+UL�U2�T�Z��ک��S+UM���n�j�kj�kZ�[j���L�UL����U2ڪg6�m���o6�lͶ�3j�e��3j�f�m���f��3m���m�r������m�ٖ�lʪ�Z����fm�ٛm�e�����lʪ�V�f[m�6�lʪ�m�ٕ[3[3m��ճ+fUL��[3U3[2�f�em�o�lͶelͶel�lͶel�ٕ�sv�2�el�ٕ�5o3nͶf�el�U��r��u��m[mX��j��m�1�K'�۝�tK���xJ�_?g��N��#��	1#�%'��a�gb���A���s�mmZ�|�iZ����������Vj�o���M���_�������km����e{���iD�=i`�~���\zC�rD��VD�[&���m���U����l����m���m�R����U)��Ym��im��YUTզ��[*���USR�m�6�lҪ�����Z�-6����:�t�o������z��mkmlmkh�Qj�����@O��ד@���
��ۻ�UEfR<��y˔�����g <��cջ�~/�ו��km�����M?�����j����V�m���n��������k����mZ�|�
�V��j�����Wk���]_��@��^A�	o�P�4%l	��W���kl��￶�:�����u��km��Ԕ��G9}������j�3O��;��n��m�����r���o��[o�W��p���r+�&lH.����ݐ4�_�}}S_������[o�~f�����������yYrsO�Y�����VA��PEe�o���	!�?��e5���� i!}� ?�s2}p#��<xU�����
R� ���	*	UQ P"J�IRH�!*A*D�T$T)*��J�����*�%T� ̒�IH����D�EHٔT����	))(R�UR"I)E)��J��R��(!H�HP��:�@ATJ����*�D��@��(Q$$�UH��TD)(T�J
BB�B�J)"���!B���@*���  Ys-��֋Zm@٨iL�j i���ѭ0-(ڭ�P�$��m*�X�6j����(*�kY��PЅ@�T�JE }CB�CBC��ywE
(P���Xth4444444;�Xz=
�{6�ͱ�@�{u٬�!`f�֩Em(�mtu�5&j���0�T�CV��D�[hT�U < �4)=jVۂ�հ�m��eP�Md͕j�٥ 
X1Zi�P��j6kc5����fփ��IV٭���ɣl�QU���J	TIB+�ܠ
�F5��-T�
��Mm�J��`!�ιR��jV�eU& �i-�R�Zi-T-mUe �V�H����*�JP�� ں��(�V�Zej�Pkj�UF�45+fѣj���hkb���Y��Q�2�(UU�֬ -�UJ�Q%P��(p  Z�j�h�
�6�5���Umm	f��d���А)j��
�`T�  3T�P(0�AUP�UQ
*��  @��,�PD���l�B��F�Xj��.�kZ�ca1��UJn����)Kn��EE�Q*�
�HE$H�RO  ��[2��(mÌHJ�\r
����t��j.9n��R��wAΚ�)PwUwR�F�6�u.S��s��ZJ@'v�ΔI��ܑ*%RE*��*U(�<  O*��+��J���]���)EMgpwi)(�ҵ:(!S���J�۩�wU����7IE)�]��)U;ug"J ��%���RQT�  ��R�%)��XU!F�s�)�����t2J�ps�)B���wnڅQn���T*�]7)"UUN�ʉM5*��\t�H-3�O��*P)�IIT�2F��T�Pѐ  "��	J� @T��L5T�   B��P�$ UF" �A
A�'Z���9�pV��d���{�Z�w�wg~k���j
�+ߝ�׹��APE|QTS��T_�APE���+��)���g����ʿ�8n�'�GF�z��6j
�>U�\Jm�v.f�B�9j�+/v�����C*m �_��(�5tsu�xe	p보�T��]�d�fݫj)e֪�(]Z.&#��j��I�6�/�E�&P�BO� ��3q�a^8�d��&��l��[�N}�2�K�Ԑ�>��
�dj�inZa�eH�CY`H�%2Nܻr��!�԰�ڽ�0�Qf��޼��ĭ�#T�D�l���h��W�&�l��a ��8�4���tK�H����k�r�	kC���R��A�tӣ�D��?�`�C���=�������k
����do*�1	�a����m��Z$z��[%����\�{ MK�$V�x2_�E*)��^�^B�]X
�$ݻ�O!���B��4(b֨}���r�anY��-Cxq��(u�sg�!%SHn�ێ��wN�]6��I+l��&ݶ4���Yy4 mңan-.��eʚ�$c5jj_[һmd-r*�jwlYσ�!�)HY�Sx�f�m��;����a퍨CO#��&�ю��ɱ^��ĩ@)\�B�|�i����{�vI%�C�@ǎ�fou�(] ҥ)麽B�� �2]	v�ޡ0,�ͩO0K�G�ؠ�b:�Kbуb�m˦~V)m���/wS2Ȗ�ldJ�������[��o�V�ca�R�V�C�q8��o�w��|��r��"A����a*�阩Y	]K�be�n�9������
_j��eŮQʚ&�OIEE!Ӄ����RJ�A[/Kn�ah9$��$�7�T,���-�&� ]�"����g$:���[M��j4��XR�6���v���R���&c�"�֖�;xU�e�6`��8+74�5Ў DT��n#W{�1�p`�1����|��4He?�jzb�A/sma��72+�@���[�1
wN��)� �f
X�Vc�s]7r�-vFҔD�U�(<_^SH��ue��`E��Tњ�46� F=^�X���g�����֛��XW�f����]��i���@�qY�ԙ��Y�3v�˥s��=�ed��N������GinQ��b�Rqܘ@0�4����:8�dr�Vy�%�N��	F���UZ��{�XyD���;�J��E�3��|6��ej�)n�iR�ۊ�I�YNQ��q�@-EnU�h�mޙ�ֶ�k��ff"T]H��Wfd�N�wmʔe:�JǢ]��{����mu�"�Z�EÂ���7����@�$1��s"���D��2�J��1���2�x�^%��w[���ճY"�n���V�Ϸ(^ n^��r���mcV�^,�1k��d@���ȁIn�;��FPɥ�3 ��c�ޚD$�.�ԫh�6&2(�Um��	���x�@ �ׇ����#V��^K�ӣR��+v�`
�vl;������u������\b��G)��っu���3/-�/F�e[����f��)^��!�@�$�}���ܻ6bw򫼗��.�.Jw/j�eEW���H�`]e�A*62�a$�f�H�B��{��������fh�l�V�p��\ӡ��$ш,�`ݷ�(��h�36[������˹��8��V�iLc*�jk�v�8�-�(�8���+wRڅ�&h�0]����R��ʕ���mn�t6;�U2��ݬ�Kk4	򫡪�{��ЪJ�8-VIH�Y���L^>�����e��fְ��zR��l�0�^�E'LiO@T�����t���q��5c]��&a�L�AX�㺻˺U��(�%�.�1	�!j����,�ID]Gt
�b�eޒ�Z��cՎT7kwnU�Thnh�Jj&`bC��Xhnf$��z6^`��,ʻ�&�LԷG
"��8��-��������7ͨD�0)&�Z���kd��q%E��q;3NDб^��"�.���(tb�Ջ�V�G)Z8�	Ow�mmS�0V�b�jUx��֘����x�-�6���(��T̚�����*�L!
ǢH��E@���t!Ǜ-)�'b�3�[i�(��Ӆ�-��Vk�# 6V�c1=Z�ɏe�s)�HF�rc��[�.����˩����m�G�uĠ�:1fa3D4d�(dەr:�������U�j�!)�O7K2֡U/�- ^4��@�֥"bZ"�4q|��dp^l3e���H�ר#���6�h�����Z���Un�ǯ"�f�Y-�6���"ϠچkA���h�L��������Dx����b��pi7j�H��;���8�ɕ0��QIQܤ��?�n$25iڋ%�b�ҝ�:^�(V����cr�r���5�ג�w��6���KŅ��5lݍ7S�Ң�n
7L4Me���t��jS��6�wl�7m'58,�f��%2�[�E��+�VP[��;�'�h=[`Î��:Y56Δ��H�$oTX��2��Y��i$8�$Ӕ2��i��0�R�#����ن������W�����MR�H]����h{�i`�֦cH.��I�p�e䤆�qP_2�_]��o~���Y�e]5D%��7lc[e� Q̴�/5�	���P�Yȩ#Zҷvv��.)z޺`�ra��	��Q��^�6�ݨ�L��F�0 *}J�J{f㩖MA�7E�.��Pd̴i��&��PV]`�)//V�A�v^�Y�i1╩Q�wI��c��1�f֊O�m�X�,5�� ��)<ae����ı��l���J�X3>ے��%��y��A�ѻ��l�<�ԧJW�^�bEu�d��ر��QU�
n�"�u�BX�&nHiR�˭��$6��[-��q��I�̕cs����Y�A��)��{bW�U���L*aAm��j��R�-�HnmD�cfNYk�^�F�1ٰ�w�Ff$"��c(�[A.8��w�y���%��4���i�:2��%P%f�^R�aĠ)(�2�,�knT{n�85ʺݨ��-�AE�����N�ʶ�d��bs4��=ciˬkfQi���R�Q�y)lO(R˛��urfR�f�g��X�5n�b4�kF�h��,6��3Y�<A��xt[�ZZ��c6�ise�'I����1La�c���q*�.�����[�e�4�/4��^�MǷ��,%Iȝ���d�
���%�l�4��Y9FJ�`m$nZ!(2�zr���	Ѭ
�&�hYa֟�j�S>]FM!xD(���ef�Y�.�	���HҎɇ&�t-J�"R���[�oK+`�@�mͣ��:'!�U'2�6bC$��̴Jئ����ډ���Fћ.�P5XnTj��X���e�ӗ�<#GB~��D��ǫ*|��++S�x1*H��	�BWs(���GЬ�w�a��x��X��JC�p�AW}�X�	��,17*ǂkKH �ґ�vL�n���]��)�_EP/,L
��ѡGv����G\S�(V��N���]6U
�ln�H�;e�)�l�7���v�[�s2�t ݇��塖��c�*ea��b�Ib	ɐ�A��wCK.��Ǹ�n�� m�J��%����Z7�ID-h��E�{MU�j���ri �`�@7J-5���]�-H*�`��ۭl�Җ��"81��k{#�b���Z��^Zt!,�17J�Jg^A�w�
U���V�A�@�qU�71��,Zz��̱��R�d)�N����U�)l�جx)�j�Ɗ��%ˣ,h�1Z"a��_=/\�e��gV���un5�j���;%=&�(n��WZ ��B��e[z��-��h/`��uy��F������6a�mEYj�AB�2��,��L8⨴�*�n�8�m�0.Kh���D��*� fB��c�v��M�ԡ�%�[4m���&�Z�+֒�+V����]b�c �tm֋4M�8�'v�a�׬G̗��r���0ual�oe^��Z*�������r�P�F�,ԩ��#��e�,0Sݢ�l��$�	2�U4�.����I����fѴ�]�)$��fJңeJ�����Z��R4]������7F��j����J
Z�6���ee֗�R9���`�B�]$��i������K
���wm]i�ªB�5��J�"p HLbV��p�`�����r�(&��J(�-i���N�ٌ]�7M�)�u���f�M0flYr�Q�P��!���ܫ*5�[�PYi��a��J*]mҙ#�F��1(�r���:����"��&5C ��I
�%���PL
�-
�V̄����;A�1fhoV�ǅ:��ī��������UՆ�3�Mō����`�2�1 �i�n�èڌ�KDD�St��n���4�i-�,DoR��f�¢�S�o��f�scr�5+R��a�I=mڍ$H׻�D���[���cG�:�J�R}G&�N���㈠�vm Ƙ��A���I��4�ڀ4�WE��z�\`dL��D�F�Lh�Vm��k/X�[6T�Y^���:�*���.Q�ՃsT��Tł�ӡ*2�!�>]�h�!��2PE�a�t�+6��HQJbAa݀��Gf�2U�����㧁A�N�+[$�lJ����9M� �v+/��dUbn�!�T6��(G�`K�u����h�Œ�h	10�.R�ӵ��V��[X��&VXmܔ6�j�6�WVм�3`�y��:l
K^�̘�׆]���*ѹD���Z	{b��t�X�XF�X�*bFR5��S��A�2��u��:�F�Y�hl�+#Ӊ��LffKV��ˊޥ]��Eê�� �8Yۘ�c�◁'�uP�aw����JSwX�6�ȷ+h�����m�sf*N�Fk�[�cT�,̄�a:��2�8�pXL�+�Q̛�&:� ��4�Iv�e4 U�-)R�E&^�R�+�jJ�%4�21)��,�������\glE.�]m�-�Lc��5m���J���% Z�Z"��-��0d�]�3hh��]1��M�cqR;Lm��dB~9�O�B�,B���Z�P�2��ú�"n�{$:��� ���d^h͵�'6נ��rA�-p NӍZx���u����pk�A�
��՘�Tkq�`�����3bk��w���1 uA���oNժ˧O
]d�(�eM͖[�rA��l�0b�6�9����2%��NP�yt�1[b_4��e��P�e�c%պ�qƳ.�R��)�mh�Y(Pۀ"p�WJ��I�&)[�u-�Yd#�kvaUz/�pE��B'Wz�h(�laM�7��M3+V%��k]:F��wl՚����v��2��bKkl�x fU�H֛3XВrZX��驛N��n��+h�nڎ��жT"�"�U�)�nb�U<����7e���r�9�%�n��c� �n���rn�U� �n FV�2�cԥm�M�XxrRV�鱷�h�����̙I|�٣.@�I(B�f��03�G���t.�ݢB�u�*���ݗ��U���呪���K�+ ,lG,�t��n���.d��ۡt�Ӵ�n��+u٫�,=,����t�@;��ݫ��^�b�*��J�ܻ�US@T�k{[��"mX�����Ox6%7B�S+���H+7Y4K���գ��lӗM	tV��e:ڛku�U���!{�c��yd�!�f�]��B�7n���rH2���f�	��v�[GNi�uJ��$���585n��1Rj�Z�t�ہ8~��B���ffz���Ǣ��m*�� �=��$2��]��u��5���:1�F��	��r�KYW�6�)Wf��!cen��ù�֕��@��ON�J�-bf큕��(^T#Bo�����`Zçuqx��\y��	
����Hj��D�/7M:h�ݛ�E�fI�3���T۸.[coc
��h��)��[�P����fA�%S����U��跑l�Y�]弭0��UWV�Z�DR�ۛJ�e�1�1�d���U���z5��іf�g	�nh�Q9���ڻm��w��XK ��湦��:��Km$�
�(p3c �o^^K��ƪF�u���x,V +6�K�U�v�m�j���@�1���/� ��'���ꩁ�H�[�n��on��ǅ�p�/T�mAC�G�L��=yCU���J�0��E[��t�$v�(���(�n���+�$hr��{�e���Er^!i�Y�R���u�	nQ�opY��`����������H�5ɷJ��^� �GJ������*PʘmQ0����bB�F븅 �.�U,N�\{�mʲX J�+m��4X�5#�]���E^*����=g$Q6Bu0�10�h,��J�cmƯ1[�Q� +l�D�d�j��T]���˱ԉ5�P
2��F�<�{n�'98���9��<��{YE�jgS7kUEja��v�Nާ��6f���^�u5���8�f�)�3c�gLv1SU����N[��nI	j
�\t�<��v��.�~�ݻkFXV��4�
`��K\�?k�#X�%ˤ����($���mmjw//wiۉ^Ѐ�f�F�ן]��Qx�i�,��x/mVJSd�` ����2|eR�<�,�j�mZWj��(��隶[&"t�(ִ-,U{kJ�p���� �if"m�V��%
iM�&&.�Ӻ��AK��vJ�3D1(o�՗�J�63^������Ž6f(=��K
��Աu/L*~OLK�BQY�c��skX/+M�h�e����x%��y���_h�R����qҺX��	aE�Xܭ���m�[�hi�1�ab�i�,�t@��
Z�'�i�s��iR����:�\�z�[�'e����  �#��M��;6ͩ�d'gһ���I�˥�(
{���7�����S�1D֝x�q�ՅZgeop�a�&��nAao2F��S��\��*����s�ku�WP�\�!�u`q�Q����8C��S�֊����en�դ� �9l�Uw���E�>F�j��cGR��ou0gh��N�����E��D5v���Œ�t.�gwN���
GC�XlZB�36�yI������1�k(bv�U�F,�e���bd�"� �8%L��p��&鳟Y�w�n�ɼ�X��o�&����@,�ky�5�0�sMY��K�X*�5�'�����z:�h�\6��jf�rHh�4Z
:��SuQܬ;��Rt2^U�Υ�o$��,��,BXO���tQ�.�%Y*����ۏ$����ݤ`��zŶ�B4��Ε}o6<W|V���7_���H>�tp��o	m�p��I/��v.9KgU������fR	b�L��{�AH�a֒[�_�Ne]����j�����Y��){��y�|���d�c���uzC׭^���ާ�����JWwrx̸5VZ�����.`�,b��RۺA���������wE��1Nuu��ԸA�v�R�^[��htPڶ�֤oU����ۼH��и㕝�����y�t3Kt�Qv�zT��tZ�<�J�����[�ݦ����z�p���;FnA����[(@FLCҌ��26H�����n�@��gl'xP�kNs�iXd�_$ƙ�sZj"U��,�F���x���;[s��C
H�9'!�U)(�3j�O
Z/��=�>/�n�b��e|\/��{C�8Q�����tC�4�ц�t���5�Alt �2�H��G��w(�L�}r�Ε�&�dCUi��l}¹��`�̈!�@�67{,�h	W�)�Q��������Ɏ�͈򩯪X�<f��8��<���m.�	�f^"}D=ɿa�©��v�
�k��U�y��n�b���pRVe����L�N�J��������;��Ǭ�m�̸O
2�'6kxw1� �Nrょ�w+3�]�l�MSQ�����>�X���F�(�߬h����Jܼ�qe��A-J�� ݠZ�뙘ɻ?^�V���*�%�rsy٪Rnb@�<x�vS�\9��Wc�tV�Z̵e-Qt
C��jX��xȻ�J�[=�\{r�aMrk=Pń������`�;���`-�����/O)��I[:c�U�J7pÒ�{��CUo-u�qg�-�&%#QM�ɰ��c_m�p������O:_a�V��`�S굃
X��٪�4�
9O��#"T%J�ɴաr�}L�
�s3(`�6>P�]�k���;��Q������H�Ba��	F�ܽq�ƎN��	>��� Vy�ђ�<v�+.�T��ag��k��:�޷� �Avw�0p�n�j��:y|�,��fRc{l�
TJ%��w4Y��]�P��dm˔��:�鲯Mcj+������w;丰�� ��x�bC��b����=]�t�<��l��-���0��(Cj���7x��I��@�n���c�zT���$���X�-�M8M)GE��7�
�X��5lyH��{!wV�ҭV;!��$���O���w2i�o|�`Ïb�	*�n���5���u����f���@*�ٗ���ab�X�f��+K��+����z�Q͡k���]B�T���,D�K*F^TS��z�.�)���]k�V�uT�w��x�Y8��M˨��r�^J��^m7��+i������S'&]�!!]���`FH��^�`l%=4��̀P;��^��C9���š�;=�[p+��B��:���wP��N�oc�8c��^�t7"�)�56�9��u	��Q�*�tKp��d����κ���*�1�]�Vm�C�Y�%���fP#��`��+�Tz��y�t��M[�X�X��Mbq��|�V�7��o�N�Ƣ[a۫�6w��Me(�u��.��t����Y9��xJ�O�y�B8����7�#].�����,��&hL ����j F�Kr��&H���9���w*͕0�����`�	��JV��'�A��By��/k�ȧ���2���xa�%�S ��S��ükr� ���{ʝ�����:J�d�i���^ ���N*��L]`hd�=Ѵ*<��g9�lb��?;0�aŇ����1U��%V�xq�7x��%��E�4�"�.J�"
Ue������GS���X]Z��u���f�pS3jv��E���1s�B���l+P*�8z���Uov.��6��t�5��@�vW!tnh��)t3��
ҕӮ��xm^w`��ȵ�؉�i�����*�x�b{k�Մ�kھj��W�&p�9���97F�6�;q@#hZ��έ�R�up�^ulX����݊ʺn��O����g���|7wv:��5��.��t9z�t[F��\)����7t>�+i�ޢ�I�u�EH�u���iVPM;Z.���J��a��p(�vi��T��*�p��憾ʻ�Bimt�G�ly���c�;�^�YIHc��\٬�O[�ݭ�����n�l7�=bݮէ��[҉�U�����#�bb]&��g{��ka��WE��wP`�=�����0M��qe��C~a�*�r��vZ,�\j�Fi:F���z�����A��1I�-b-RY��ִ��u����ܕIƱ����s$5�3�d�h`���KQ��7(ʻ��fu*��9�2��Z6����k o�v|�;�j�7mv17�[��:��K"���˳��i�;��&��ޕ��w\���h)���C� �xih2Pʳ�"�ZX8���՝{�)��A.2�v�\q�I�$�:�t���Ώa��-K޾��B��Q1w�D��s�;�M���]��d�]s�k���q�n��A��+$�̋����r��Q�2�S]z�;H��9Zn�o6�PO�N� I]�[�˫��I>�{�����9�-}��D�LSJ��F�]6�ZIԦ�S�5!�G�дn�{4er��f�)�ꛥ�n�ffF�_�|��g����������Q���J���	cMC����6j�KO��H^PY��N�t$.���H�7������#{G�|;�a�v���FޕY�c]���������S�u�"�>��}��ھ���[�v��$�Ծ
�6�wyN��te��q�Ԣ�\��ܷKG���lBt��7�����Ga�8�M�;�,R���+r�����)خUk�j��ܝ!�7�9��(�	W�q,��i���7�����5c:��R�nmY;B�7ܝL�(��n��6�� ���XBhWƷ��['+�<T�8�%
i],Ꝫ�t�J���}����<4�k�O�2��PJ:���|�>i�2�
X7�kE�*�t{�C�2���ڧ��.�����Ԓ�mm��q��X(�R�e�	۝o淆Ɂ˂���L���قڻ��Q�W��p-�{)p��o2H�G���E����B-����b�O�b�-.��ֺ^܆��;1p�S�O�J�]h��2[2���4;k�V�n�Q�ͣ��9e��̸�`��N�׆csx^�h�L�K�y%�B�R���h�4���l�`uHRy��,�k�L��Qs�:�y�)יӰ�ޮ��7�H|��e�{/OZ-4��޹5|��s����4�<��Q�&�ne_fSsu�v.�����ƆRun��ᮎ
�[���=�����7l��d�iU�l����y̦O|iAW�u�"ĻU7�l[tj�(�W�E9�E���/lBw�U��1���n�μ��2_qI����=ރ� f���ظ��	�Ƙ��d�αb����#WB@�MVn��
�cɆm3�ͥ\{���,�̌\�J���D��G��GF�5��wD&4����9|$��"�(Vs�9o������r����J���/_*�_�j�s����
]b�Ε��&��=��ȋ�Y��t�J�Q;��L�p�i@d���>�(+�G��YXg��Q[Ft
�k�ֲr��V4�9w/Dk�Ogo� �)e������8d[q�U�p�ٻϴ�nr���W�¯�����:��k���%�į�+s��M�)�:�kNhw��" gJ�ZH�9���H(m��I�^S�Ct�[���d���0p��\��z���`����6F��vڮ�v�L��V7+��<�)���tL:�Y:�nT�{}c�X���)��|���yM���>��~�5� ��:[�`s Ƽ��e���b�����Ce\��2�L}]1�y��*��^=O�>�c�n��%:�^��uż�N������*����]�ǘ�0�ڻ�k�]Z4�4��t~�ۼ_�f�Ƨ�h��<�5�-U��j��B��:�j�%
�}ئ̧`\/@�u&�lB�_T���3���<�sbwP�Źl�ړ�s�'Wt[c���Xg)3˛�����m�[bI7k���2����O.L���f^"ͼPk����A���dP�7g.�B��K���'n��\|��9J}����o�!�;���b���Y;�n3+UMS���2����y���6}rO^Kݢ�æu�E�W�ݼL��]r5��J��j�5mF� zk�R�m�bƥ:䯸�y�˾�V����+I�Z��r�o��/;Г�Tr\��� ���|����z(g���I�
��杆1i���)Z�6r��7\��I����J��}�t5������o�[U���E�ٔ��̈*]��ڷd�j�;��Ц)�Á�شj�*��+yg[Ёׯ<� �%�n��+[�G�f�S�N�%=���9�9��[���K��za��/U-�]su�Թ�/5�ľwAdj�Ѝ���Z.rz�4�l�sv�]����_v8Db��j�'X�v�8'_q�iL�u֒M��b��zX�Cn�a�GP��-�;��\�CQcU��d�J�D���@��ehV�ͣ՜�N�Z��&}2���E�d�}�̫�6;�'�8T�͹�C���t��5�]���9���+�iY�ˮ���۹�-g��t�{P]v��zR�qnZ�����|�t�ESJ�h��,-�*���C�5����%��v�d��|��5ʆ8is�޶�Z�cȧM�춮M4.���/l7�ٛ��_f\]�	z�������p���:w/\�Lrf��v_pȷWu�����əg_j�ն���*s�7V�
lmCt�\��ݐ�q����ሉܳ����������v��	D�ۧV������Ie+��Etd����e�N���V٫����ĳ��1u�Xl��q<vo���ӌ4�	f�t[��qQ��<�i�7[CsK��Ӓd��#�(o��w�noLaa��"����߲Ǎ�H$I5�f,�'|��Y�Z#SP�.��nwo���RA�m��∬���36NN*p�c�Al=ǻ���P��Ե���s�|�,ވ��v2ڶL3)��r#�*�uwK�ѵz��_..�=z����1YRS��ګ/�ZP�D�eru�p�R�)�ŕ��=�2���'٧Q�~��p�!�t�1u�6]�7f� �S_PU�m�@j��7�v0�"�(mwb颋�*Ծ��%���t3oW7h��os�-��Jl.ڡL%wۉ���[��9���W-��y}�����u:��2d�B����&H���e
6x�귨�{�˵�nĻ
������n���t�i��l:6�ت�Y�/�^�c�*p���"X^�Ѝon�����8c�����QWr�"'�:�V�30vlt�8ʷOz�2";4[�vo�|T��h�A�+.|��
�%Қ!	�y�xﱯ1mwF}ݚ���� �*���W���톏̱�h��gp���Ä\f�S�h<���*�:/A�fT��2�%���,�ur�X�wcj��xS`���E�F���[�%\ѵ�Iki:g��ԯ@|��*}�{��	k�s����9;cE����τՈp\iWa���[.��qÈ\	�֥A6[;q��7�k6��`��E%�Y�
q�y�7�r,�Q�d�y���Kpi�*<в�&0WV6�;N�h���A�7�ˣz����8�v��X�b�W���1Es^w�Z��4��f��P�:�m�G�Y��v�Zw{��5��]3� �B�%r���nN(>���aK�t�D��u����-Ps9�쮣���K]WK��ܮv��p�kpg'Cf�n�cQ=%gu)V`�
��r�1�ƳNgh}|#��X��u�YO36��t��$`@u<Ady���w|�V-�%4�13������w ��@KE ���.���5E�5�e���M;6.�XL�a�\�Hs�nW9յ�z�Zv���=K� vzp���"��i�l��Κ������[cR��֪~���n�a�m��4���w�_X����[nhu9����U�K�]�T��Ir���sW�o����36u�N�����y�AuFG+JHStF�k�MJRU�nH�7}�}V��Z��7�0v�Y���a]��$��=��,�{���V����q�֒O���hSַc���R�Y��G6h��]b�4�YXG��M�q+l�J�;��c�����o�$o�k�d��L�A����BAu�W4:L����h�N�A%[��2$�5ֳ�+\���]D_V"P�Ʒݹh�a���7.t�/Tsv��jt�����w.gj���$�,nN%^�^��~y��5�]~���EQO�PEW�g:�,�O�b�xm&��[4�?
��D'4�l���Ҕ:��x��SE^Rֹ�//���c������gPbwڒ�C2��c�q�W�͂x�i�ok��3D���hv�T��:���K�_L�����8���s��m�M��s��z�KN���a���m�w� k��C�T�λ�ʜt�T����Jn7�f�����6�%Z���n�`b�ڻ��a����D�u��G�@;|�q=�}����S�5.��j.�����ESmL�P�BX�gcG�AI;�28*|]k��`�j��1����[H���P�9������m�AP��3k����mB�\��%��	�S�c.�;u�)�U���|�a���"�fͩ��7W;�C@&�U�q��$�wU�q�� e���@:�z�:�h20��֤L��ji��wVJ��]꼈�m���V�6ow��U�=&��0=��ˊ��ΛO�Z4�6�ΛD�3�K�8 ���^��y��bI���C6ԁ%�횛w��Ws�"�8�7(�R���M�6e֧��wl5������굵މ�ᵹ6�����-�fl<Ù��p��X�6G�n�'_}���� ���5-�j�Ҹ�4�Hr��2�g�R%�Ԃ��p�ѝʑ�f���js�Y�)rM��EI��L5��z��S9�(�1�wW}���EtVWY[DN�ϛ�Z�P�=`!�2e�1��ONT'�4��3����܃@��dT�5��u������,*�9�K�% hQZ/%��Mo�'%N�	���6l�Ey��Q�`[P�gy��wZ@���&���2����m#yI�#���ٶq��+x>�0b�w���:����Y;g��{�X��2�gTi��V,,L��U5�7�!���3R
P�⤹L�j�|]��|�J�3���}q�B�bX�p��-�׳#�5+F�T�o+�{({z��t���kJ�&N�q��u�����1�`�[;o��1N�������xJ�k!ˆ���r=�)L�h�dЫ*�QI0�ZQ[-���G�_}�oT��p4X�/�3��I�W�Xr���}bҬy!�|�ԋŜ^�ϑ/o%j���n�Oz��|�(�s+o|E��N�{;l<U,T�事!�Xj]��j����v�����^�c�MnE���l��4���l�Kc��.�t��]�׶�y���۲J��^F������T������|a(��52��S�,�6da����X�����(j���^��s�A��G{8�����t�R/�� ԲXG�*ɕx��J�Tg�v7X�zqN����Qٹzy74��l�E���/a��$����%�\���D�v��G�2�������J|iu	���}��;�i��Nwl�v��.g/�W[׊���1rO^\vy�����٢�]2;Õ&��3UA�N���s��
x]��v*��U`���*���^ާ��|m������o��l �R%a��ݝ�0�ύ���k���-@���2��]G�:�*v��%�ݷJ�Qd��qۮV�;r�<�X�;�qM��@l�O�E:Ϋ��]�cp�0�����ݺW�MjX9�\����|ރtei��:�Y[5V��S1��gװ�t�
�,��p=�
��Q�1r�a	dp�]�fq�͛�d]�B�s�$�v7�OgZk��^!V5�Q4��XڭK0��3by�8� TJu����Μ�6��8�şh�v됹���V�֡˵RS_s�O�ژ�QXե���-������0��ٵ��1�s��o@Ԩl����'Au΀o���E�X����p��iF�����b���]r\�:���UQ!D�!�v*�3Z�ө}�\TR�h�YQ6Ee^��"���:֛�)��-e=��ĞT�u�}�GE�H}%���O3LU��G`[���=cj`P�f\[���mvݹV�y�K�[�4>yF�wE�q��a���TX"{M��e�/o�}IA0���}��@�Fq�GD�����)t��w�Z��tAc��Y��^a�ؕW�xwd�(Z{FK��%�XρL�+&띸�i��W1WIZ��<N�T�6�I��M̊�ޮ��=��E�D�R�к��"�u�]
���R��4t��=(#�R�Gmؐ3HB�˽��W�cpm.L-�xe�5�s]�[��Hu��3ݱ��ԫ��m�m�
ѮF��vU�A�Xy�׽:�ed8Wκ�p�*�sȅ��y����n�М�nj߇e�n��5�0t���43 ���X:��
�Jr��ZV]g�R}�~�n�I�H{e���g`��5�K�֍�S\;J�Dd�0���Y�6�L���S� �K�ۙ��]=;��*^�4Y6-��6a}��'V�Q�(t���b���oaQ�g�h�]��c*m,�܂�"gZU����{��u(vKND��J�:�DKޫč�+7�>��N�]+e^S5�F�*��%]��yw�y
�c�.�YX���xM�����I�Y+'�O"��ԭ��o���o1�X�[��)�h���!�k�MR�DGݎ[�jv��:+Q�5��5rSЄ�n8��p1�cn�̷j���\��A�\�Gj��fWn�rpՙPC� ��Y�v
/!q�@r޵�
���z�����E�8_<O�w�!��d�Vr7j�V�JC�ֻQb��i���Խ�wmc�#\���O��/+s!1�2���P��u[�O]%�u�{֫�3v�s��kO�)�k�c<ѹ
ި.�\TEI��Z;��T�fv�A��
�;>|��>V����R\����^�r�F]��̾} �3�4�4��L�m��S}�����[v�_[�j]5O8�ba�#�j=���2��]|�^�A�j��]LD��[-&����M^v��v4 4Ӕ�i@�[�!I4������2mMt2톨P�>:��qG:C�0eH�] 2�\<:��AJkx�OU+Wز�m�+��y��V��wJ�c�Q���\weˈ���X�T�]
ӕ4��
��K��ۼڬ8Fi�����_H�e� ]�ELG�%�=wP�S�B���	1Օc� S���)	���s��� �<����&ڕ�+�]l@�Q�N.�C����;in�8�;N���V��1u݆o�M�iƦ(C�W��p��kw�ZQ�Q�[�Կ��Cy���l݁R,� 3ɂ�ܕn����*� h��=3!r�QtJ�Ce���x�����U�`ͦ-�0ސhm���jf�x�N�B۳c����;���!-B���mʕ#`�����E^�]�`��R8í���F��԰�̡�4����j�/�Q�Y��g
�?�܁�/TV�z��b^y��r�J�P��5Y2��4�R1ͮ�Aį��z&�e*�N��aj�)��U��2|A�joF]�b'%ꬦ�ee>�f���M}	�Dꊖ���wnݘ�ǯKۭ� �Z�J�j��H�ͣC��ǅ=�ܙf>����u��gV�t+�q�ۂP�G.�hN6�w6��m'�1�l�g-�o)��l����pv���,�
�����8���#�۷��QM�{2	N΢�pf����D�_p��A{:v)����̧`d�VaU�HY1^\" T�8��'`���顐��D��n�|l��<�]�tE7�eN�WNmZ��^ء���0��V��\	Huv[�\/n�Ѩ�6ķ5ǣE�XjT�P*j��
k�V�1��>ܸ,՚�(�[�z�����p֎ʂ�����a P8�|u�sq4�CZ&[���w2�Z�}�-)��Q�hWޙ�g����f������me����6��#f��I�L*����b�;��9�y�)l�\�r����q/n��H),�gw�:1�T�9�5��s �kzhQD�J����V�!ZM�,��H����ʺ�5/%��y�`�oq���趱7�]0q�a����ʛr,1ӑl����ݛ�	���T6��uwk$�&>=x��̘�H ����/6(ά����߯+)*��{6�n1LJN�W���'^��f}�s2�ܷ�z/e��Wt��r�r�Rܹ6]>� +[�F��0=%Y[Wxf�R���[T���7��2�X��!BиH7��#���P�d�n)�@�ς�v�մu˄��Um���-}�ׄ�����*�`-�Wƍj`_=����%(�vB]W�('����J����t�h�����ʽ4��7H����:�f�C�g��Ti�Ǻ�)���:���p�ʺm3/�wV�n26b=QӉ[����"��U�͍Ю��ބq�X�r��9�2ZoA|p�R��x>΁U��V���� Y7ي�%$� �o��|j欜�A���_<V���5󩡈�1ش��}Z��-��N�|V��J�9�> ���6g!�{�m*��_X]�H�.T���SES����Jh�];.җۗ)4/�-�F�ik���T��νM���C39RU'!O��+sM�2��f6��8��l��-�p$���ҳ3�Afm7W�e3�%��P<+aT4y�g׵(�]hUPs=|�Wc�n�N��R���}[{�A;�wIF�m�(��*�5a��&E蹔�YO-ͬ�PX������a�#EA����,�9m*����7��f� �]]khڒ��P�M�p⫢8qX��,R�T.���G[5�<O}�)vHE�,\cSR�����n��ݣ��8H���4�[ᕺ��嵭;ة�TA��+U��Ѕ�RN�Q+���a�ep�z]Y@۱�H,�B;G%X�4�Z6����"���u�Nu9��ܹ����0�Z �)H۪ز���w�|�3�HGg,3�y��7���lhZ�ʵ��q<��n����@-㰳
��o�E;Ҧ��^:�]����Iջy	��Aj�������*M�T��1���E�R��Me�<w��R��lmv��r�+Y��*��aS�w}w�+t��śQ��P�B���ej	�i���T2�p�Q#I������m�Ѝ���2����!	[��实p�6�q;�{���8���'[�R5}��l��g��#7�yAJ�]�q�VŻ5C�iU�i�ew:��f>ޜo����zQH�ovԉS��̏B8�a4	�IV\�  S�'�h懝��vؤ�R������fe��|�-�Ԟo0̼�$�DDj\3��9$,�{f쥚喲�}�/`5t�Q�1��M0�6L�Q���3{��5`��^��y��3�L�gZ�)��{��oE��o�R�-�
�v���s�Z�[k �,R�%�5"��eǲ�*B�*�Xb��m�f���/��R���j�.����W��>���%��o罯:�Cj�XN7���U�	�X���/_ݷR�N�sL����صƝ�]����:�ͧwD����ں�����������[I�.�������I�ƘL5Ԣ����/c���`�Y�Z8k�2��˹�kL�ӧP�]��I��!���Yױm��=]�d�'|��C�B���	
���T�p����v�s��]a�����Rʼ ��V�T�V=Gf!���1�nZ$���ʒ�Ûe˦jhv̉��2%��ul¹Pt�k�79��[�D���÷#�$q5mwm�3�9��t
 n�Y���0+���ڕF�N+�F&L��u���ܬB�|�Y\��wPk�+_>��6�΂,1uwV�����:q�(vS��m܁�b����zi��ݖ�ϩ���sp�-u3.�˩v�	e��r7� �:�]Nq	kS�ޭ��Zp�윛��-��PmJ��S�ST���������-v��F���rjx��ҚA���X�n���^��|LUh$�NL��	Ht!�˾�r�YZ���j毯쮑.n�q�m�r�u�om+Brz80��n�T��EXv�7�3N��Li�ŷ��Onr5a�� �8�7�����,A���'P]���A�7��Gr��Z �Okd�Ed��V��[(˘��b1F����B*��lfѭ앥����B�bS�f��ֹqzD�Ӽ9��P�y��{�V�������F8s���q�ٗ���!\j�Y�8X�ܾ��=������R T˫��s��$�4S�ų��X��v�tN�7�f�L��;����v;Goo:Y�#\P������i�ܻ�x����Ck^>��ZU�7CTl��U����1�3\�(��H�eIQW�>j��:��q�U�R��I�J�4oDt�J�^V-L,K����0�wM�3%lv�v2
�qUa��iu����H�}@J�w�w�sT��ޭ���b֤�X��ǣ+F�e��M���¡Tr��3WVTF믍v��ewau	��f�y��s.n�d_#�u��Jz��FTw1sYQ��Yx(�&p�w��ϳ�Y8��B������m#�VGRT�
!�n���`٦r��F�"7�.�PK�`�b��=�)fEy��K[sM���T�l_M��j���C���z��^ǔCT���w������*��҇t��u�'7]n��,�� ���>�|�l�˗k.�q#� X�b}�,js#6n�ݮ<�\��"Ŷ�P� ����-��5H;��G?8w����J}a���)-�ü��6�6`n��cq[��.o{u�V����E�v*#�W$r\yC7��a�諟S���*(h9N��� �CD�R��/o� ���ӻCm�W���tx �mWF��te*\ |{�㒚��&���.�Da�[�2̓�M��s���ks^ m��Aeܖ9Q �}�- +�..�����􃔂�Ÿ.��j]:ŋk�~��諭������
�=뷩9�>Y>�շtTxw�o�gB�1�������P�����6T.T���h�����9�yH>Ғ�
p�v����Zu���3�b2�Q��%٣���wFR�����]���)Ҁ�^e>����롌����.�$̧�n�d��W�e�����0'��"Սˤ^��s�n��,Mvq�.������K�Q&�#�Ջ�]�R��E�
���`nQ96jF���ֵ��e�*�q��M��٣��\��nw��ʊ.�ۓ���u)�b�X�els�n�(��z3%�������Uc�k ��ګ�[q�s��F��B��f���R���z+=i4;�z+t�ϗn��aC'@V&(�ļ|�l0�Z���{K�Ȫf�0B#w(.�$�J�!��r�Ͷ����(�r�(Nl�ښ2{.���6�=p���M�ɵ�E�,t��;;y*���U�m�@D�օ��)JW͵Ϳ���%�a�0���+k���Q3�F"�L�~�OSKxxm�MǴ��_\����F4{������;hr��{��Nb����Wf���I��5�ҹa���v5(���	����\	|�-���X��nݴs2zT��[׵j��l�2�+�/p�ڕ.�M'�j���m�|���s�rK�5�����b���˂����b�Q]O/��sB��VSW�u{�;��sg�~��T1AE'Y�Y&H�P4��Hѐd	�KB�-ED�Uad���FJTM-6fH	��9D�4)C�d-4�RRR��E��T�CJ�C���,�R�%14PRPSM+�AB4�,B�dd�#QU+Q�BP4�@�%�E �4DT�@�4RPR4��RR% R%!@1�P UT*P44��PD-4P�T�B�#%)JP��RA@UKAJU-"R�	J�*U PƗ�]��7�7�]��I��UhƵu_�)�� ��/{��ȭ8T3�Ή�ǜ#k������tB�c�E��ܚP�z�}�k{I9��tE�6J��]T�c�7L�5yq�*;�\\B]R+�h���u��1�;⎦ކ��&�6��b��L�l}�o��}���t���J����>([����Z����o���2Grt�:(}�����f�1$ܡ�Z��(�.}�����P�s>���`������ٕ�(���\]<k!z��b��Q�Pa?��GPdjY�6sXw�����ˌ�`V�YgΩ��үn>w�܊��+W��uvN��v ��΂]���)�E��l�4�.��fF|�;�\C�l�+����q�s���E�&ܕ����̃�e����b`���2s�@%���crEZ������Q5V�O1;x�!�,X�(�Y��r��NH����5a&;9\,���lʋ{�fz2��Ii�3�|l�>58P�g�E���aR�$�D�C�}uH��E�8��L�>3`O;���v\�iq�C/�F���y�\h�� 1$�$t�3�φyz���&�s�.�x�)��;�+���˼ڱF���)\,��E�c��{rV�슙�TԬ�b{\p��%j+5!�8�%vp\.dg$;�������$�oLr-��YS��w��T���������{[z��-���-}�V����q�u�7��W��������]�v9���q����0�s.�� n�81���s��v����4AH��g���3�19ᠷ���P�N���z�'M�g�e^�W0xI��Ι��`���2��Y1?KU�z�py
c9.�&��D��O]H�j�j��eT���C�`;��0Y���#Gd��[N��u�G�#���C�6����	�>G�u�R����N�}�x�q�s|�u����a��=�Å���fj�/�n��.�0P؆K���z�buɣɺ�3�b��V�㩛\)�< ����g%7�i %��U�E������f��חw|c!���(Nkw�n8�3���F�s)]�L��wfއ�h�cQ�Q��I���a�l����ʟdd.t������{{S�q,�x����ʓ�9��3�@�1�SMA,`9�Hێ��8��'\�4df�q��c3l8��&�)'��ǎ�K ���o�ݿn�fS'�"H@���*0�2%i���d�kdF�-C�t�`>��|y�J&Z���V�8mSյ�յ��u	�%Zh�W�VKwX�%n� �I�%˫����y��ב�F�v�0z���f�����P��q5a	�Ds���}Dӫ�W+d�
�����;�:��5j�5���-�@��r�v|;�T8�Kł�G�F�9qV�ճ�3+b��'×�<|&ǥD���]��\F9L�ߞ_�uÞ�mօ���'"M*'G�KJ�ߚ�{��8�9˕��|�^+�&Zu򿴺`�+�r�X���q��<tA�T���e ��#�Tr�R�&6�EU�\r�(��ĉ��폵Ô-A`#�	�EC��W�R�-y��w&I�9BI4�́ ��q�0��S�;yʖ0[YMϵ���c��lU4r��P�V��d�z���:jД�f	N���eb�Oj%�-�p������e��r���	T�K�[0FT*�%T��@����J��L�/w�#x����Y���.���Z[J�U�\���w6��@�8 �I\D��D �g�WT�:6^�1�bx�R�8t�q�,�1h��'���'1��.m��W)� �(�[�C]��B��L���Z��X��������7��R<&Ls�F�nb5���]Dl�2Mq@Aؽ�~�O��x1Mb{U��0����u�������-X�ə��$N��wL]7a'�&es�Bۻ�eV�x1}��Z�>��b��1�
�M�r!Q%8��w=�$�];D�5���b�b��Gx;a�f��S*#��rQ+��t�|�k��]������"*�w�0d�xk��Cj]���$�� �s<ܰ	��8>���j�\%�=��f�,|��>Ŗ=؀�k*J��v$C�!�o[.0Ֆ/�ULB�!�לI��wu.�t�vR΋�H�p��n�H�L�`�#1W(���-U��*�Wxʤ�>���8��ksPK�ܮ]5��3��*�"�LM��Tw���`���6�Ui{ģ<s�^����͜�9M���n��L�bE���j���?:1�9���gZ�>����#�^�~A���a:����,��1�S,�t��\cv�Vq��`�C��`�k��P��
��Ph��>c�^8:��> �C�"Ӗ�c��� �񋓖/���}��Q��`bZ����0t�~�g�=LmL�9���TB�v!dqn�g��a�����6B��v��j\�ț����L{��.K<%l��F�$VDj���(?b���~�q<�;�1��;�νS�[�����f1��[�#T����� }5%0��+�Ս�]���Y��_H&^S��f¤͞IY��MTH]�Ѻ���;)m�F>E4ڛ|���/9Wi��NFV���V�}��;0�wW;O/��a��l�&X��]p�n/f�..���z�L�NbaFtq��6��ss�t��y�OPv���%�#n	���܌�sH�Dr@�U[Di��� �/���n�j�]��F�Q�iVP��k/zxoD�m�ω�-�X������3"��Jl���҅�h6�<���a�OuoU�#����ɮ�2Þer�a�����ŢU�_B�1+MΕF�40V$x�z�>�&\@����Oa�499w+�M�RZ�Cٟ�sT�y�Y��w8K�sP�z壢4�����Gi�򢾕պr6��ͨB9s�c!�WD]I���:��ǹ���^���#�b��zY=�M��u�onW���ƅ[ ��[�o�;����K0Bo]ޜ�s�9ʬ0}��z�O�+��
�\6|-}�g����|� ���ڙ����2 �>���ڿ��=1q��2������i�b��p��u��7��������u9G����H
��k!�2��`P?W{M�0�R������??P���-޸�������[���q;2������
���uM��W_n�S:��iX�(�iޞ��ʬd-��u�8���kJV���A��V���v���8^r��y_f-�E24H橇�-�7���:��f�.yz�
�B�0��/1�)bZw�(I|�߆m�U�����1���m���w2t�v����XoUĈ�P������?T:Op?1(�αx4^N`w]V�H>��*Ԧ竕oY_-N^Js�����1�2�G��йp�w��W?����V��S���p�Xᐶ6�Z��V^��Yx�1r�1�9Z:��c��ș@C酝uH���Q��%ޝƱ�00�BD�n�d2����O:� )��Ǡ ���dlv��G_P���\��2�L�~��Uk9�Su����9봎󑧬�?eC�B|*J<�9��d_��������BF�Ify)݄g�W؝p�ڿ���e�N��5��X�M��G�5���h�׳��<R?!BY�G	�Ky�2�b�����0rj�P[�LP��2��I�}]W]��q�lPD����-c��0Y���G�l�9r���_0��Ť'�,D"-q��{��r/9p;�pǸՀ���S�\O��Gx�:�G��r��^�3(�Za���fW<+�wK�����Ď���4Sr�.�>1����y3k�1�`�M�]�m����L�ޫ�,�G�әv�H2(��ce ƺ�V��ќ.���,�0c��ǃ4m�������[�O��y�6�&U���R=ǳ�[��Z�6+5s�ߚs!-[��\4hA�j�=��7a�{p����Ħ�͘Ziu��I�i����ɨy(N�7{f��3���0_
v7S�"��&Ξ{\��Sn�F֫I���A��401qʟdd.t��>���eX��Ϻ��yHt�ywJ�J�ܢ��;�g�0�ʘzj �0� �Cq�Nu�h\��u�o�l[ə�d$��/K쟦��E�GK'v�������e2{"$� �\�@Jg_j�}����8����G�q��^,�����]dU���H̭���J��R���C��x_k.��	e�_')�nW�}Ძ�EfO:Ц(��9i��%��e;Ȥħ�8=��μ��T�c��Dit���ea�岲��ext`���� ��͡��3�F�\�-���b�*��뒏+��:�1�k�Hf|X�j��}m��&��U�m�u�J�$��<���E��$o���
,?��hƲ,탩���G8Y���c���BK�U���|>���)�v�̄k���Ė�8p�\�IN�"i���6�<�B8����Kh��V4߷սh����_+�g��O|9n��c5^9�v3£�C�@��ʔk^ۂ��x1�ݖ�t�w �v̠��i���M�8�I�%�=�z���V.Jt��u��[�h�j�Mwe�Š��w�����X0�W�Q���#�@�|�����d��2����}��ro����`���8!�̓�Cn�s���W�R� �����Aa:�5kT�r�ٔ���cj9u�)��"��/!��3#!d��;{���uENd�����R�"���^���C�<*LW$��l�cBkz�yÇ��޺c�����,o�.��P��`�4�^�V%[��gv��I�дXf���L�Y����Ö:����Yґ���RF�'�dÔD�:��S��졤z�N����]�'P�=a9��	�5�{aAYk=c��@��0�:�_;~���gJe��m�� �����Z�2^)��:��5u��ޘ"��l�dx��u�ͧN�!k?*~}~Q\��fb&�뇟*��' P�v�W�_M�"���d�r�dV�9��d��:�G|���:$�J��`+�P�Ts��W���/��M��T�l!����9���	�ܪ�Osf�0֩��8����ւ���T�8�k;��ǩQN�i��V�ƺQ�w��N�B����\<.�g����X՛U�L��Қ��Y-���)�t* (�vgf4b�����ˮ\��H4�O3,k���=�d�N<��ϩ�]�G@�8%���"��.�-~�C�"�9l�����u�'ݒ�����Lei�{�(ݘ4|ѳ=H^�WS��]���T!pn�b�\ ֵ�:O�b�m��׵��@��ns���rx�ITg�?�ԤV*������zph[bgTo�E���|+%U���g�Z*����'^��:E�qa"����W��p�>��cr+L��s,w�1�z�#i��ⳒR�h�:�^d`�[kG�=��켚��M|�P��cx�����c	�-���ۘ��T̊�L��������%SxU�3�V�EI�sB��C�,;s�쯹u��|[VY�&-���4T^��,:�r��*��:N�	W��4�EȻM)��{=���~楒�.�����|�M�U�n [Έ���'(�n���]�0�ELl�f�!�[Y8k!ғ{j5rԏOQa2ܰ4�.ho���K'��auF���ͳ�}��N�2>��7�푲��y���:��}w�R� 擩�>9���n=�Mr�yΖ����IJ{��ɻ�f�pJ��'Dd�rڴ�����o��Bܱ��-��XQ��Q�	S%6����˾���K/b��>*@Q�w^W�����F&s�W��hk'm���ޕ�@uӂ������_�9f��~X�K�ٳ���z'+�{7$�I��~����ey�?O{g�:�Y�S�6��)t;�}�Vv�jj�pt�}g,m�NQ��N�';e�F�YdC�WB���w�܊��*ܨ�[Ϭ���/�\���vh�t�m8��E��	��_3#��Sg^ν�W�2�t�ϱW6������r�Df�N��>% ~�d腥���j�K#��X���:;�oޜd6Z�����Hr]g�������[��s踓��#�.���F�ÓZa�F��/�Z\Ԏ��v���˼�q�Sӑ��^;��9R�w�u�e	�Zxq��!�u��׺������V�`�53Fu��E�_F�o�}�C/�F��םP�A6����x�t��jƹ�*i�͋ҥ�R!� 1r���-���UZ�E7_���㞻H�#�������C�90N�mu�W7��Oj�Qqp@�P]2ai#I�:#�΍.��@w�Ƨ;�����:ތ�cڑٹ�fVLHҕ��r��ܮlJ����M�@��VnAYjE��p���0&�ɈV��Y��YW5-\��G�|�k:߮��E�+��r��ә��JX��^ɘ�[���3���En�駣Y�hu!�D�0Iޞ��|��N�Gj�"�� F"���J�=���ˉ<і;��\��G�$T�#x(1שu`�*�wN.B�|� ��Øi��)���8濥���ò�2Z,h����uu�Ӻ��S��Ȓ5�nmfL��Ƚ��������v7�E�\�̶����'x-(Kt�8� ���}���F�p�g��s2�P�aS�\7���������f�n� =�c����HZ��0?r��ޏ�j�N�s6����77th9��=pR}V�5|�J!�3�񹋢W/��*����dsu��]��Ԡ+���֢8ݎ�@�6to	���WҤ�ː<�n��|�O8�89#���u�͹�@��lm��`岴��zU��p��S:m2 �u��;�B2�J�zhR��J}uݹw}Wx /�9�U���Q�t"�k���Z����:n�oE�CuC��U��k��f�Vh�of�˭*�.wm�����]��2�X�X+u)�Q�`a���bn�Fn�8mx�[w3�7�n�jW�B�#'��]2�yb��<y*�ψ0�H��D���{��F�=�a�w's�1sT��%�/^�7҈�C4�wh��Mŉ���2�aut�ΘK{\��m-�v��e-�a�b)QSO�`}�"�L��)��JYd˳L��s
�W_:V��vp���h��Ö?�vKY˛ɣ�h����r�j�Q��W܇I�Ӭ��X
˴^q�����S�K8��K��q�%'0�;w�L����R,��e�OQ��.�IX��<�zR,���eM�g�lv�*�-c.n@��7���2�K�T�Lde�Y�Չ�>�s7�]y�9��z�i���Fw[ꏝ�l�|��W�8K���4��[�R!�^ܗj>�*s�ʍ�+:��[]wۢG���$��ul1�(wc�������:���}}�i2n\�c�]{`��vv��.�k�(gu�(�ɦE[쫔�����7lXtSj�5ۭ΅c�����Y5'6$���#�~sr�Y]P+']���仺�ξ;՝\ӛ!�-�`Xx�A,߱�5!v���
�Gw|���H�Ј�/q]�[�͋�����:���2,���O(��*pO��|���v����*\���Fj���x"Lm\�Q��̢5�D���WW������[�w,р��w'�5Y�4t�	s��S�}I���h�,У|��vvo:�*��ں��S��J/Ę��z�u�~�&�k�����kf��|�sx������N�z�;���n�m����K���F+�H5.�`X���R	�e�\�;8�%Cn�]�R�wgz����:7���ځ�*!
j�)
���Jh���(F��i�&�
J�r �(F�*�
J$���
@�31�X�)hi�r*j�@(hF���)��$�(�
U�(��r!(�
B�(����)B� 2fZ��
)�������G$r�
�H�&(E������hh(iZh�(������#�>�*��rt.M�<�x�V����'=�q��]��!&57�n��:�����q�|��|>8󷵁�2,N\OV`�N�n<�ؗx���R�)ܝƿ����5	Tl�QA��5�f`�<���n�]F�+Q�1w�Pjǽ�wQ��?��/0�^Ͻ�t��2:=��_�����e�Eu�ψ�Y�9N��e�@{.�U�9Pe亍p���N��s1����%;��bZ�婧�:sT��`j�Xy.��d�h�N����������5���=�]� ��|F^	ʄl�9�:3�7�R��&A�%��7���r�_~ϣs乬~��5���9.y�v��C��������;�S�=�@}jԔ��K���OZ��7R�u�G����� U{�yɽ�^B���T]3{;�8d�s�<������Cs�Χ�ﹷ�;��N�s�P������� �j�]]�sK��L�#ۗ��~���2^�q�~��jN�sp�٩v�b��  ��Hy��{6g��*O#ϭ����\�˝c�ؾN�B�����?A���X���R}�����S���������BW�{��������.��2wy�惻�{�Hv{���}�h���e�v�w�f��ٰʊ+J���Q��9�~�p��y%��.@{G��j{�#�{�r�%�j���MC�r_����?`�<�;O~���~��������?Z�~��=�*"> }8FS�xw?IbiU�m`����|w:�;�2����:���5g�:��Rj<���Z�U?I��_���/����\�%����2K�������?A��矹��P� ��җ�8�#�&>PD8q�)��}&�8�i�/� �Ș�D|��T|�>G��1;�U!OS��7�ΰ}=���N��;֍�S��WN���P�N��5�2�ރ`�F�a�f@}&I��k��<�י���8f�n�Z��|���":�} 3��F��Û�B_��|��{ͿK���w�'s��\���������d?N�C�3���Cs�?�NF���$>��}֫�U�*���ӥ�c#R��&Ϲ���_= }�F�#�mO��	��٭sc���5/�c��������������z`�K�<��`uS�.����w.�O�s��?A�R�5Q�b�`ːb��s߹�g:�;�钭�Ĺ�<�X������)�D����kJ�/^/_�X{�����f,}EQ�<���+o<8���R+u����o�:f�V0�~���"�]6��YSN���JS�Z��4�W@��μ������v��H��ŕ�����>�lT��(N~��L��G�>����u�/.�p��^��f�M=~��^�(~���é乬C�sY9�Q�?�Wg9�7<�I��?<�G �����5ԞA�����kQ캈�}iS7�St"}VeU�sV��|c돵�w-����7�z7/���^ǯ;ڹ{��5#�����_���i(�a�{~�(=��l>�G��A�	w�w<x�N
��ZU�6��}��Q�0:�!��`��A����pFI�o5���yn���_K�jO}����r^��6~�e��5�iy9=˓�s�?�똿N�S{�7���*��������b`}p�E�	��Z�~��~��)���5&���?��������n��޳��z��Q�,���������i��e΃���}��KxG�����:}�[Wowo�lD}Q��>\����S�}�C�{.�]��bnA��똝G_`�;���7�]_F�:�NK�������!(5�>���\�g��n~�d�r,��k��8g}�'�\�v����\��D|�\|&�m��J������K��4��C\�K�ƹ�?GS�\���/p�NGg17��u���կ�}�VF���֧#$�%�}�����=�5�=�;;V�]10&> �Ԩd�Pyy�{�!��N���=�dj� ���v�<��ԇ��C� ��\���j5r?kI���2:��w���;�:�Bj�|�N��y����{:o5c���} ?���T}r���D���˗���������.��Z�߽�í`�<����y'S��%u��>��ܚ��Ps�:�� ��zg�����`�h�;%;ϻ��;���չu��2k^bp���)��1׸=��K��g��S�\��u��:�K��?�I��^K��h���2��iz���2x}�ms3�(
�t7BF��ɿG���=���p�.f�Gks�\���q9��ܹ�����5&��:������KXy�j�xrߤ�����&���k�쟼�Gp��%��g[{�D}�GƸ]�v��Cb����AN�{�Q�[ɧ�5^�룞����xL�N��T/ho�=�u\�����L��ǯTu�K�C��a�Z�c$&���D;P��%k��[k��NQ�e�<,z��Y�%g��� ���B��ƦGy�v��ى��\;�ﾉߧRASԫ�}�q#�#�ܽQ ��bl����FOr��-]�Ԕ�\�~a��:�reI��P��A�N�3]��>���dy��J~�����~�R��N�O�d?��ur�5���3�ѹ8��7f��x�� ��'}� 8�?9��5�C��w�採*�/Ѯ�}���-���N��.C��9%���'O�n��b��WZ����H��1�Zc�#�>���.�53�����y{�����5!�]ks�9�W�j?'���h��ߴ{P�1}��=O�!��u��hL��b��;����*�c��M�����0��r������j^�O|ўs����g�ȡ�.f�T�h���� ��2B��#�P�=��W�������}/Y���n5��乘?_>k���\��y���05<�5��w�:�G$�{?�u���%>G������BZ������g_���8xn+����>����F��z ����k��:5��c'�:3o%�<�.��F��3$)��?A�d�Z���sԹ��y��%%9.]w���GR}&T�}���9�ه�i��_OnF*����?�������pw��J:�=���;��ԝ��j��2-�Ƅ����5{.�>��:�rn=�����������_��������uͯ#��\�6u��4<��:]W�V�����# }�������P��_#��k�����jԝA�0L�o��ܚ�cR���MF����J����G�j���'S��:���������\�������0k�^�푾c� (��}�K��{�P�>�y�%�O�v�掠22>��Wg<��C�2�~�q�������Ժ�{�u�nr\�^^��P?K���f[�y.T9��/H�0�]z��;��D����>��'��MF�����Ƶ�&G�y�9��n����A���5�~�N~�׸�O��9����]C������fHV�q(5/�����1���j�U`��a��5��:>����?_����!����}�cRrL������j��ݏ^��>��soprF�/γOpy:�O�j?k�u'�2N��r�-����a�ur]@n��y���e~�|'�)�Բ��{eM�鼦dTw;���ٴ���YIZ��jP���N�r0m�;�8��KK��h��==�6 4+$�
0��S��(z�MXִ�.������*[��q	�޴6�qt�S"<se� \���He��ͻ��/着���;��?��'Q��z�9;�P�~�����:� 7�5�}/���\���/��/''��P��/�߻r�(O^�����g�&G�\�!��MO#R~ִ��##�ŗ��g�GV����7��{�U-h:����>˩�uy�c��%<��0߸?��%k0�\����;�K���]T�{|�A�ё�{9���ː���{��7SA�m{��r=6���)2�c}W��5�/=ӹ�\�_._�ֲ����o���u.T�P��O�tf:�	��y&�u�����)��{&��?A�<|�I��C��n?y�P>����yX�y�6�w�\��}<��mz���=��l59.s2�����22_-s?kI���r���RRS�o�w#Q�=��3U!C�y����'����'��2��w�2/H�kX�v����`���Ϲ<����>A����bn��������/�}��������~��:�$���?[��N��J�c��h?Gp�C����K�����e��_g#n���1Q�.&zw�;�e� �o�'�����<���3�	�[��}�&���z{���NF�������U/o{(9A�K�sbn|��c��uBS�1�y��� �G�j�`��&>�"ւk��1ӌcO�g����Ժ���h�#�9���?��~�γw�z�T�� ��u��Kvy�xgުWF:�G�:��=��mG��ŭ�6/�Z�wJ�Ʀİ�$�U��i�t�ve�,p
oM�B��ޟ(B/��9Z{|�I�n��2a~���~�qަ�?�{�ύ���v�b��m�,�.�D95Ʊ�q�\�
S�;[�ݮRC���S�g��R��>��8]#�/����"kʺeq��"A�89�Qe��:��ԨlΘCY��=���E���^m_���Y��0g*gT�ٍb�{t���w�9��I ~�ջ��=ws���{g��|+�Z�g�&���������׸��V��Vx��J����z���#舏�QFΦ��(�l�;�Y��ӣ��w�r��蓮�@�}`�����/"��Jq=w[�0������ʇ���a?��><�e���p��[�63{���#]��|ʊ��l��΃����UZ�;u��ų���i�r4��~�맶��]�P�����:ĺ�U^�Ӱ K~*��0��[3�N�tGB�\8g�ڿ�;�c{'k��D�˷#-��Ka���}��JX`^?p��}Z@�tIo��>���{+�_ol�,S�/7�I��zGy.�W`wJ&,"ju�\<w 3�����]딏V-��^r�a]�8�jE}��<B�/�N�ɤ�p/>f�E��Rf�Q?L@!3G��#Su&�\�i�T��F_�����{���O���H���4m7@s�r�_�OG�e�MVrx�-s�V���ê���{l^F�-5�.$���C��ɧ���{f(��[��}t�1_f����E"�n�1�TxpW�j���ݔ��r����F���z7��U��x�Z욡�V��c(�u���jz���J�v���h��j�;N��ie-��c<Q��څ�%����k�<y�mߢv��g>�0̛
��8���WS��(.a��ƅ�@yv��S����{��7�sR��č¬�w3���R��}�w{�]{�{���OM��ͭ��Ϻ�#
L< !`�� ��P�C���l�Y}(�	�;�Ap�1�^�f�aSY�	*�q9���.�����QXtR�� ��lay+X�6 ?�6�FD+�l��?b��Dm��b��X�8��ǵ'y���k`q�z<Η �4\u�CF�fXWK,�E2�<���s³'�hU���+�ȓA�Xy��k��oG���1<��#z�G��4���?�ƗL�,Vn[+>v��1Z@�C�s����4 �u�A�Xcfz����(�+��5��_������Źj�Nr��&˵�׸��1����_��x�=�dq0��]Aw�p�J�0L�{�fG�3E��ݝZ�<�5�D9�U��s�]>�����TUpUG��2���|_�!���ͤ0ˈrU�O8�;=�;��>;��&���ꐔIS�@Ć>	N�z�R�v�P���	���±���=�_rr�؄�W6
J��eL��٩H����N/WMSז6넬P�5�cԶ�w%�5�@�g*{:S�q�6Θ]AC��x�`ҋ�!;��{S�
���ΨM�% �1�j���1���,�ġn���O[B��ͺ�{z��!�ih����C�:���rqɐ�6uYW�!Uڋ�ܭ}'ﾪ����-;�_(N4����FT�tn�l��ck�[���i��� �)��u���p�q�s=��>)T�T1�kU1"���.;�i�Έv�I��I٣m�F���U0u�;9�k�ah�F�s�Q/��-}���ӥ��ķ��]�b�5uW�o�;�}�/�h����h۪ܥ�JE�/���	��8>�yRDl�e!]($>u�ā�:�����,*���3�٨ѵYy�f�(CZ�3]���Vz4)�g��@��2��:�i�UN��t�����p�l`���fU���a#��W�{��GJ�Gag��Q*�{ip��]�M�+v���'�V�i��SȔr6f"��C�T�d�b���O�}�ab�X�N���,��4E��{[���Q2t���j�Ό��PjsfX
�MCQ�S,�t��5�7@=����#�q��ݰgL8�`�P���+�?�XxR'¯�|��.�(�?�j!��")��'*y��>�!�K����ptE]��w�+_	U��~WBC�:��
���|��B��ʓ�n�]z o��ܢ�����r�)�~!9v��#���P���@:���t����v�4���w̚ �Ꮶ��WO�܌sȹfG7w$�V�dlZ�X6�Qߖ��U��R�]��\�ּ� tv�|3�iݛ]��`]����#����q}o[���=�&�~`vJ�O��&�l�Dt�<I�EW��\i���2�	��!��6|RϤ^P�O)��Q:xr9�f6� ��ީ+�����Z��G�t�W򆁬�����W�(C��6]�ڱ�e5Q+�c���L1�S Fs�r2��#5�@��仗;����Hz��'�1=��2�B3�cx�-���)�f2	�-��06�&���[tlgD���S|ʪ2=Q#��k�D*G{S�s��>�<>����[VY��F���v*������>I]�|$\���n����Q��MEܮ17ԃ�����7�C��3�saR9�M�IOԔ�y�,yDE�?'PDON�!i��WV�Ͼۘaṟw�[��7%�1l�8EN�����Q	��7��@b�9`ix�U��c�������jʹk)���Ѻ�.^��cS�UE��Z-JcE^�B�����r��>��]�&ob1U�§������v��p�}k>�rY���bT��3��]�^b���xs�Y��ee��v�}@D�UX��V	���0q�(�y}t�_fx�>Ή�<�)�N��z�p��'k��k�j
�R]Y�GGl�ݥ��XC?\�g����E���?*�	�!6p�C���6���5�)A�w�3����c[�{����^��G���E�״����TQ�p���
NI� ON_ݴ���Ʋ�T���S��5`[]v�q�=�l�+���b�eN� �a�>(U\��J�b��+�d�� c�Y��.prϯ�7\W���<q����`�<O�|W�5ұx4^N`wr�w��IA���8Y�ϊ��|�ܑl��W�+¶Uy�j?�ۑ�s踓�����8�65�w��<�F�h���-k�����ӑ��c�l�t��5::�N�H�J8��
�vX|�\��T�A�)��2�	�ԭ��C/K�?!�:� )�L�ؾ�sơ\f�N�t���4I<���f�L�~�3����}5����i�r4��ݖb��M�v�=7�j?Ob�X�G�� n�"��F}�<�������Z��[W���0:�&�fM�%�t��� 5�Ʊ�.48� w:	�K|���lU��u���zw��3��������.�=��ٷ|ݠ�O�P�\6�@�x�$@f;>���"�~g)�����[�����um*�p�z�s�<a.�s���s_�˕]ۥS��;�'Yc�QC�X4Cy&JD��z�j���i�t��Q�a�8i���%Z��}{P���4,S�
���<Q��V���x/�������U}�f�m�,�;^�]��|�
����ri7\�i�4\B1�L*�&j:Q?H!3;J�.�1`�j.�8n,�������v��K�i>���R+咙4m7@sb�Zj�8[/$���zǽ֖�EL���1�t���Ҿ��/v]��u�;�1�>����J���M�i��+��ٳP��c0U�Ϭ�zP�|�y{�*���͔���O��Wa�Wr��}e�B��\�Ȧ�|�i���[�;�s���a\T���R u͢�/{+a��@��w�`(�q	�3�1�o���В�q9���#ܾ�QX��i������8�
xՓ��! &��3�s��ֲy�荣��ܘQE�F�9 ����L�^J��s=���\��w�toh�l�
�%�Mr�������3�3Ǝ�ٹ8��3�X���*G�0�bg��S���T	��N�W�����ۖ��v�ϸ���a�����up�g�أ��|�8����mW]3��E�s&�S�>��ä.z������]�������M��ǲ]D�j�&��04t� �W�HBt��ѥy�f��Ψ��]�Q��-��{��=)����W�_ ����
m�B�����t��mWY�d���M���X0�j"���k;;v�c2�i����������݈etQ�[b	�%��{R�q������,=v����k�Iv.�}yH�:�k�<�촶�R-��X�+�o���F�q��x����Z�ZL��g�h�x�\0u�=�T��_4v�E�t��%r���WN�Ѯ]�iC��и�6�}�_a������5���Yz�V�ԣ��z�� �P4 ��Ov�����x�'�����Y�[���'�_NC��]J�1M|E*�<{6�׺	���k\�9uA�^u��ݧ�=FCjvZ�/T��[J+�2������`�-<
��^_<����ή��7��l�9���;{&ݜ�%dB��<ܖX:�f�WT��[��S�Y�k��CSb��=��vt��k��ʱk�L,�ΉZ��p�T{gp���b�Ua[�f43F��ɔG,��=���r��7���Iجr�/w�|�X�!�|��o5Q�f�TL�K�N�`^d�;,(�W.R�5[�׼��k��G�VspIl�n8t���)r��W�ʕ*6.sx˸��[Lb����0���V#�axK�cb�(֬�5"���v\}��s�Ah��[)����B��Ҿ�d�uσ��J��������C���ۋ����#0C;#zpu+�9غ�n[S=|�0�n_f��w��-��rj�|�utҫu�kV]83�����˵���v�
;��*YǞ�z7��8�bCeͰ�'�(:����dn��Q�F�Q��\C���t.�(;�ݚ{�Ջ�s���Q�T7�dp��͗gl�WQڛd�C��1���e�Oo_�lh�ӹ�����q�S�Y�o5�m����G���wO�D�ܡ���V�5"{�T����[j�:yfA��4�4�kpX]�t�#�{��P�w];�j�pK; �.ܩ3��t�gF����(�B!ᢠ��o��7�yʣJ���%%��.�&��c���t��=kX]�5�!ק���U�0q5x�Y*�q>�k�6o[Qa��S�5�ij^���KEN�n�!�����1�3:�W|��ʏS+5�L�EX��-L+���˘V��l�+S^����0|KR�a�oUf����IQ�s�j�OZz�������$���ԼڏQ�{�M���wt�dӓ�;M�d��_r�=t*��ȿ�J�������]2K]t2�[���3z]�Jaw��s��o�����V��vMNǥtWu���oN�i1����C9�˳fr����X���ʂ�C&�e��i��͝܌�O�]n�w�Q�<�F��[��SQ�qܮBM���)\wwz��ݐ���wb%/hѦ�g����^��{���o���(J
(@����&�
R�����dĕAUMSEL�-�4�P̴Ҕ�,M�M UPұRYdT��RД�PE"QQ�d�E,DC@̥%@U	MRQIT-%R4�P�	M%-,@�!BQBPД�Jd9UH�ER�JD)BPSHд�P�R�%-4Х"DUH�aHQE����>�ʷ��뽬���}��91q=Ģ�'v3�6�n��}��ݝ������i��d�_V���2V�ӊ��^�;k�W�U�}��k5�k��$9��\wdA�G�#��d����'�{�Ⱦ����������AdnR������z�KxXor�1��a�sT�:|"<X���⫂=�	���뙮`@�e֓���v�
~��>����8R��s�IofʇT�ҙ*k���U�UقU@q���ͪ�I^��\G�V�I�V�9�!�
��p۽�ࢪ�"{Lm��ݿ6%̚s��g�M ~�����_�e3p7������Bs!����/�&izrp\�0��̛7�m$��)W�v�x!p��57Wa��dzW���ow�e��Z�P���ۥU�`R�(R=�$�0�8<~����Uվ~���U�ݲ}�^z$��WSِ��]m�%mr��a�-9`�����8|NT5��f����϶.�ro
�-.U�i=Z7Q(i��D��Ӫb�֯��MC1"~�u"+
'0o����v��^B�z��w��X��$���g����c><s7	���DՏ�U���������Mb�o�J��������#�n�Aύ�)	�[��dZ�rE�����S}ʺ�r�粘;�e+L�;�*\��'w8B�j�ڻ��Q§>V�*��˾���K���'�eK�Ĺ��zV�f�r+���0��������ꯗR=[�߻��#�X��j�`��D��l�D��뇟*��' P�v�M����Uv�����{�P��[�³h��7>K�	}��o��ms���a�|�2��wM��.��ٓ��g��z!e�-]��vElXX�R�z���_:P�%�ͥA��Յ����=��{
:����Rr���'	z=�*i��m�Ŋ�}�:V��7����s���`����Z�Kc.�Bq�;ё�&ˈ�@-�������b�񯸢J�?A�%]c;�hu��{��ת��u�K7�l�_����!�����>�H^�s�N�@j򣝺�g$uɩ�l��eH�sEa���mX�9�&�&�X�7L1�q96����=���OX{|�mn��7='E*θ�DL�_
�2�B1�4���d�o X�=����7g���,\nks�V�J{[�A֤}�#�X�BG}����1�K���*>���2V��Q�����<Sk��L_���J����N�J�҂�4�E�H�M)Y�����U�B��Ԟ༲Lڃc�k�ޓ/��=s��Z��o����L�{��g�ާ1ݕ����8�bՀ(�{wmK�N��6Of��v�A�'[�9a�s��'I�K���M�w$���w��n}2���r33ԑ�9��tz\�uw*�/���G�Df`�^�nv��g���2^|�5���A<Q;_!i��u`��=�5����	2�0l����\��ϛUtoጀ�|��4��r�\��=,�����m�#S�.�>|�
�A!G$/�'p��=��+�0V����s��_���Wsa���.^��r����;8�Ǒ�h[�d����F�Rgx����ey�5=��ݬz{� (ԏ�P���9<��0Y�Y�5n�ׇ*�j�F���Z|M��@Tn5��:�p�sњ�pC�ή�˙�z���UX�ά��! U`�i�Vn����8Heu�ɢq׫,Ȫ"����V���ӿ���;�tf]yma�C����}'s�LT��[�-r��]��4��bԯ� �iWc끍�jSs�򘎿�W7&����Q'NĞg*�fw97(L���U󍩎�P#�2�UB���z~a�:��/�*crn�u�6Ld���,��q*zی�IH$�6��B���a��0a���[��3����+�[q� m0�����8����+��/v�+5��ͼ;��-ek��X�2�ޠ��w�!�`vu�3����:����6�b��h��DW�,�`Q��A|�r��u�ʗ������z����s�Sg2]�;�RRlgP�Rd�=�EO+]�DG����n��5�I�.����f�`������O37��H�x���N~����㞻H�]ܢ��uC��{<���P����Y�~�SB�%�v�]1&�*6g�����]p��նl�W�7����;�u�W��,n']���q:n���q��i����[�϶*���w�}qYJK9wɝH��kn �I5h�
5�n�x�$@f; �#@��m��g��x\�2����j��1P�
�Ja���p/>f�E�1�*�o�OW������ke%���v���|3���;|X�8��5v��'��jbG,�ɣp��9����jzj+bF��x�]/�N�Z�j�$��Ҥa���7�",\Ϭ�y\�M;\��L�>�	��=��W�ۑ��+������&V�aVf�W�*�V8W��u[9�1y���١a������j0�v+�켺�-J�r����#W�k�+�T�x��E}�ٮ�5^���41�z�Eփ��o�s��ŷP�������=�^��a������ГW�(��:=�U�B��C>c�<�nĴ7H�}V:�Ͳӗ��ͣ�u��
������6xD��e�V<jG⌠����=B�z<�d���\�H���-#.ax�l��vr����P�9^�o���jR5S��������
�Z5��,���^�`�:����|
�9�W��B�G�̮'�"H`���&k�O���o��gT�h�g��µK��کfi�?z��Pɵ<N���b72²Yd�)L�ח�p�n�:�3ep�]���\WCz������&����	`������l��Wޯ��,��Xn��W�K��R�Oo,7������f) ������� |+����n��<etT�����av��a1�Yw����V9�`3�	���g��/�$�|e �9���G��u�nE� �-�!��W�c�P�x�a�YM�r0���85
�B�%C�3IJ���B9��vz��^tM����Tb}q%��]>;��&���e	�2T� #�A��LYp���sP��UJ��=��"7�|��}_rt�؆�/+����T�T�����@�ďJ�U�x��L `4xEuJ�v8�f�����tz��\6�tN+���xsv[�y�whۙC�7�J��k��r�C�p��]�.tC���1�`5J
�6��>U3r�B��:���WU�8[�R�52�u�f���M�:&�]M�,i�@�w-Yl!6���Z�����|��r���t�'\����3Jm�s1���G��l;�l�ɲY�6�u��f�J�]Χ9�E�xX��N�B�UUU}��s=ϖ��>CAb�w��v�y~��2~���62�=5�l�j�����9}��f|����Z,3M� ���8>�yR}����� N���^$&�|VX�vM����ꝰ����BƌE��ULE��A��,,A��hS����7Ƶ{�a�T緼&�Z�h(T-Bq]O��"�v�g6������|Ѹj�'.?e���R�Dx�8̋֫���s>L��^�&+�u���l�sfb&/�\52�d�Cۄ���¹#j���oO�?d	��f4V�8r��b�����ߡ�ms�x���ׅ?�˙`��vU�y	�w^ͭPњӯ�\cvk�4��l�\+���
�>u�PEg�]XTސHѝ`�Y�Ҡ�Y�Or��!	�g��p|q���R��C@V*��x������ƹ�*z���(������5N�C�[��&��@-N�xL��.O�*��}����幮-0�ȵ�����1��S��h��u�K7���R��>�!�یt�=ꑓ������������w����1x�LͺMj;gm��%����l����h
\Q���u�7���:%W��\ X&y\���*oX�lyEVA]1�c�LPK����b�[�4b���/�ft96�u%���꽥��-���Wh���ۧԲP��u��9�dٗ�o������ꪣ�M"a�u�� ���P�Z)��݉�ӯ�ҔR�q���9	���܌sC&��F!ov���#ҙ ��eǚ�B�wW�AL��1�j!oWȔ�M�h�s�GR �b�Ǯ.F���TNZ�fB$�:j~U6H����}j��ς�~>�&�9=f��d���N�r��ݽ�x�OI�}���\��z��a*�@��:�pyR.�K��Ш[���#�u��bF�՝DppT�Q�S%�,y�yQ>�����C�����e�{mV��J��Fy�ȏW�[��f�u��1ͪ�7���r�Xx~�K'�.���cn�p�;ε}v\Aɰ��U�v����JcE^�W�ޜ�s�r����F�YS�V?G�9���/;�^���j�`F/���(�.}�����s�Fx�{2����l��7� y7�yfF�cN�v(�_��~.���&2� �ᓁI�?g�x�s�P��C�/�x��p��1R)݄#��p�Xݽw���,9\h�UpUB����q;3�����M� ��w��˽>H�|�Τ���X���Q�0��jmu��a�_b��3�ul'n9��҉��:���MC	#���;[�F��5N�3g�4�(tu��!�_WG��ᾤ�5(����Z^l���A7��mX�Ľ>�9��{����h�`| ��+��a9����#>V��/�T��W_n��\�ܩ�YD��.	�	���[��\�7J�7��"���������1�"�.����V��z<0���F�ȸ���ai�`�ivJx[��d?\��8!���]�Ȏ.��0�c�lÕ,gM֎�6&QyS�V�v�r�B|��xpz�e�?�}uH��)��C,P�K|Ğ���
����[�;3��aM3�Ƃ��ɮ;�G#���
�����i��׊�Y�n��-�2�8���B���B�E
�f�L>��^-�W]v�h�� n��!|�vb[�Y��B���t��'k�{cy�lA���|=1p܄븛z�'M��~�����@J�N�YY=�DO׽����.��0���o�ڶF�}p
�ա�[�LXb�&�u�O�~��>5���K-s�uY�nc�;��(��9}]F�۔�Vr����Te�P��&�x�0�F0	UJL���a�s��W^b�V'� �����%�`���l��zW��_�ڨ�_,�ɣi��y��4�3��wD�ʓ��;�\��wS��q0��j��+߳6�7Y;z9�p�ň�M�k�H��/X��1�|Mvc�R��O沇�����ւ�XZ��0�c��8�*ڍ��;ź�au��٫�r��u��GeΡ����~����>�����,-����$�b�:����mm�����.�Wa}��	'U��M�Z��X\:�u���HO����ȗ�0�PU�ʳ���yJ�hW�W�k���_��}*��������m�������1��|v��P��[Vf'2��7f�SU�>�ڙu���n�<P�h�r�� ��u_��:��y�J�&3���U=j�s!U�s��>���D�{��G/�ӓ*�2{$� ���$g��&���f㚮}s���h�/Vo���s#vX燷��K�Kl���k���ت��V%���||K�)���<���s�7M\3��m�}<��M�
�+-	&���%��do�GR�&-9���L�,V���=ylx��%^Ʋs�9��Ba��g��u�KB��~DtW �
����?�<�H�ʆsm�F���Rz�͔>q�!���7�\�~�#��d��(	�{�e��]���'�/�W�񲽼�4*�o�Yb��<��g��a�s*al���tUp�Y|�xZ��O��y[Hl�9��q!��5�Ef�l��&���X��
�,t��t;b�dK&ԞR��6�Gr�W)^�Cw��$͙�P�x3���]^A���]��c6���C�r� ����n��:x�ʾ�2�Fz^v)���gZ�lq=ݑ>�_UU}SL��OT���W}Ì��ٜ���-�p����N�q6�`��T���d���i��:8�Ni�Z9� q�G�m oL�/vH��P��}_rt���6p���X ֢� i�#7�#VV�W\�ȃ$�v\���l����\tn�L��1�����`�û;��l��k��l��v�ީ�'��av�S� �*�U��v˕x ���V��2�]�1]mNo�}em���R()1K�.��w�5�ْr8�z�O�@�1R�ҳK{|�����^���w�Q��w����h��Cr�&��8>�ו �d�Y�����kOxd�AA�tgr����=EZ�7�&��*�"ֺ��/
#<�2P���.a���:nvC��ok�����+�q�����9�N�h����N~��xvǙ�@��r���J��9�T`�q,1POYgU����[�x�ؕR���o�|B��\k۔ȵt�r�#��^�\�����8�[X{�lܤ�[�	}��8.��cܯ�0���۰��֔���*�	n#ǋ5�l�a�;�m(�2a�V��>Rih�M���=�Y�x�\���rwJ�b|���@�x+��~�=m'���Y�ծ�"33��kH�������$.�tOG��ޫ�98���e��	�,b�t��4��Ie\W)�]g�BT^ke��mG�;��=P�m�N�{��D���:Տ3�Y��1oayt�h�l��� vu6P6��9���l2n*����ҠX�ʹ���crVLRr���ϯc[�5��*>/�rnQ�"������8���gT.wJ�}˝�*&�d٤`J�˫���m����[O�W���ń!�S�P�)pE>�ۯY}.����|�u�D�������V�u�G�*0��Jܙ��י'8擲�����%�J��;���ǵx��vj}{O�+�W$�N�8�s�M{6������+'�#��ۧڗ7��u0e���뻱ѭ�*�\
f�#̗���mw^v�A��J6 �4�Z�/��7k�f�oz���תtcn)�XeW:\��YVdްIXv�uQ6���
ԡ"��𠂲Po{_�Be4wf�}0��vյۇ�Z2,��J�v��� �vz�*��nW?��cl.xY\�G�Z���V�Ln��27�K}�ts���#�Q�FA{wWK�٩�ro��;� B�j�����Y�(]54�>o i���p��k|;Vt�^�]�mJ��Ftn�u�8b��:3x��j��������5����`;��]esc�ۏ����И����r8s)�����L�����[�m��g3���x,���W5�]�tN`�34R7w�����#��&�&�"Gn�vk�����u�-s�6}���Rj��sx����=��	 i�������6�y�V�f�P�`7S��kz���J\�t!��W�:���PX�0<��(�p���vp�O�oZ4�v;�8���\��re�&J�|������Z�[S�ոzZU�A�3�YG���j��ۙ(�v�;�VG����*gwK�����/ ���0�R���-���a]�r$�JR�Yͽ��v"��BAӽ4(���]�d��4{�Y;Ru����䅷b���K-E�8�|��fW9��c���Z����)ص#sj��۝�ܬuf�^�N��7�8����b� �.�k:��=�5��I^c�m�t����cV�GG:oG�Q1�C{s�f��]��F.��']kQ�Ɗ��U�­_*0�U�hMB�Y� �����T�yU�M�S�/���/��ݝ���� 闗��m)vH���Mj�;��t6f�uns{��T;p��h��om]� ~��Q]%p�y�����G����kK��gV$9�Ioz�	��$�i�!�.7�B��[:z��a7�w��`-5��������;o�u1�:Cs�6f�v*ɻ����]{�~�������RP4�A�5TÒ�9�VI��H�H�-���PP�	H�	�Pd�JJ��d9Vf#��d�VIH�%%"VC��R���% 1)Y�F@dP���A@SH�#M��!�dM��JRAIJR�` �ݗ�b��[�W�%`��vx�i�����։�	�N�B����a��Vl;�Q�JʺAl�r��=�����p����������⚺A�:A�?���*/MfNw���`6X�����< h�EFҠ��n�T�w.��̷��������
����9L���D�1P�*Q�C@V��QZ�bK�6�o�5yyXѣ�JX�?*�N�B�-ތ�\L1�������:;E���SW��m�,����س�?�#�.�-uTK1/'��*΢�x���L��U_+�L�QS÷��P$�쿤��_i��[43�Rj�ne��eL1�S F1��ۦ$��N��>F:zF>��5� ���dK�'�J�e2�d|�o�<4�I^�G�]�m�n�Ug0��������~(:�r����1���%l�^��O��W%ñ�֧l}n��amYg	�D��f���J�k�NЙ�pz�dI�䨛{q!�C�j%[J�9�K�\Ƶr��?s�d��5�P�*i�q�(v�ގ�ۺ�H�Cqd���.6��ݨb:=�2Utn2	�KȄr�\��kr.k�{���uڱ+6쮅���jih�V�x��k�͞�+��o2����Uɳ��t�vu�i;Z�sQm�,�-륎�VpC-etՙN�vJ+��6�@C�ި	VJW�ħ�F�j^v�ܦ	��]����*��%uH���q����n��1��2e���������m�X�\�g	�+>96:�+�t���P�Ɗ��pB���.t�9l}�����gkU4��J�/��Մ3&m��"^�r���a�Z0�@ �w��<~=�OL%͘1�P�ۍP�#�Ҿ<��w���YZEA���#��68x�7�)�? / ��{�o�0���\x*j���>�A��N��u:�gНX�Ϻ��Tcʜ2��l��W��P�8�C,o�[��h	㇡�^���@O֝�21Zw�^o�9}ه������W�9�Z"fK�0�hͪ�q�#�9�Rv���}�ݏ����nu|򘎸�U��ɺ�c��FY�n��u�����r����$��=����W�a�����W\qt�柘y���	Ҧ7�m�ݍ��d��"x�k����@�iY�IƖ�^��ebx�e�,P��J�d2����B�/�c'eMm՞�lb������d�*Ǡ ���<��H�x����ۯ��>�xp;7S�ԗ-<,<z�̌:-��ØB@�(����F�	�r�6`��/�n۫:%�3w2�a88�S�q��`��F��NWIet��!W�1���U�b�ˢ*�E�W��kea����K���f�ۛ�ox�,��)�;���:D1t���e�{;>�{�`[�p�������D6���Ѿb�of;�wd�""#���x���#֝pᒚ����7��^�����#� %Bt�9M_�F�ҽ�HD����L23트-ς��.�rj��&,"i�Z�wP`�U��YܳA�5Njv��n�}�Y�"gv��떏VBW����J�ɨM��`E�q��5��U��w8���Ez+'��.�O��[X(H�r����6����1#�Jdh�6�Kst��1�~~��Y��l��&��j�*�WB�
�s���?5}��'��mt(��dj_��k3��ϻgF!󟔗�	͆�l�qzg�:E�.�J���
��{Xh�DC�{��y�I�Rй��dа�r��s��'��G6����@�g�{>�����wԬ3َ��پ�	؋��A������8��Нs1CSCt���1n�E�.'0���$"��6����۬��G}_M�`�'�H`	��\�F+�l�~<�zc�z�ý�j�-=�x�Z5�|N��YtV:ٳ�fV�U�3&XVK,��)������Ͼj�]䘓��u�)�Y�9 o&A��P��*�ѩ&��RR*[8h\����:BX��e�z�ekN��cJ��	�<9�j�Į����Оqyz�>�ڄN���k�#���B5���rB�'`곴+q��⽍T�pދ��Oo��}_W7�+"S޵f���Ѱ�I4�u�t�ߚ���F���ݡ��7f2O�])�;�k��@ü\.�E:u���?q��E) �A��
�����<n*Υ��$��n�{���{qb\[v���!�X�j���~�#��d��(	�{��}���[�=S��� ��V��)lDi�uYϴԬ���X.�뭔"">Z��˥y�9�t;�ƅL펄�`�T��n��!��F'�Kw�|s��M��`��uHKg�]�t-�Y*v5;�%K�,�4���Z��L�/w�"7�|���NR* ��������-��Q��V�J����8�8 �$�"O��& ���:J�:8�f��1��.�E#U'��;xj;u�u,Sp�Pe)����g)� ��C
)V�}C]���LH�(v����it&��X�Ws�A5�S;xGYBd�杚7�F�F��6^8"z0�����Q�3nT�L��g"��sMq�1����I�дXf��`_G9��}�*A��Y=C&>yy4���k�{�P{��vr|�:O���n	Գ�x�o>�ef>���������H�7��@�0�rτ����^
�`�sD��UֱN}M��n�(�0m���52�%v��R�����;õ������v1�7:����󻝀\<�l����U}�aݎ�������N�a�۞�#z�тh��ʩ���kc��^4��F�ei���(���5���ys=V�oj[�E+�}�3ћ}lA%ۙN~\\CWQ93����7��
s'9s��X�z`������(>����*q����@����k,����jiQ����zs�):u�fl�f���+�Շ[�l�K������8�=˱/ݎ�;�Np�k7���Gx�2�ϝ�g�q��U�b��e��^�x:
6�ʸXD$L}7*��}t,�Ҫ�φ��
�P���3��>�3|b�]�(Ѐ#Gɚ}|a>�C;8xv��Zc�ת�����.��&��@-�N�zL����dQcQ�~���NR�9�/��D���f:��Y��Y�Ogꂕ<9�9��:i{�#�4��;x��K��=��h�� Ԑ��
a��	�j��Ϸ�ư�g�A|+�9�At�H�N�	\����r2��3Jdq�䈻����<*�f��Z3:䮕���t������Q�GMA�y�=җ>=���C�c���ELɅz^�y�nj�m
b�wY{�{�Y�{�x�2�IJ����6�)�o�\kt�T�q�	H��f-�cCmeH�����T���\^�I8.ݶ���t��%�]z�VWE�T_%����iY�W�[]|�����-.cSn�r�S2*�JD��i#bO>�Ja��)�So�b���.m��Z'��R���S"ڲ��W�5�L*U��LsP'��UFt�Y�)X0�,�*K���boz�z�Ha@}S�}�S%�,j(���"/�'r4�]V�uv���=�0s���-����sEu�����{lgͪ�1���D',/ʰ�{6�&��4�ðzy�<���	W�a|����Y΃�we;,�uS�K=�~ٝ��u��6��J�=���z�܃�)��+@��ص�:Q�\��Iӝҙ��m_��9���0�}}-b]Ѹa��E5U�k4�#���>8:|ճ�O���*oϼ��ub��ܣi �'��}�\1�u�N�wgVq�W�k�@]�\%
�����b R��4�QV���5������\̎{��仍����:,�-�2��}�n�tOu�q�`��0�#� 0E��B��ڠϸ�����䊋R���yLGJ�z<2�Q�!���W�����3@f]xd���á���e��D籉��3�-t�LY����Tl'o�w5;�.�܎$_��4�E�3c9R`I�+.m2�%��Gv���e��3��G��\Y�����:�� ���\��G���dެ��i�ꪬ<V�p����G	<}'��2���jaɨ�
F�j���qt���~a����W��iߗf��L�=�Ą�'��1���N�L�$>�WuH��)��|�&�ԭ�^|���f��=�h�g4���V��&�V�ƺ ����΂���Uk;��c/8�5�����E�Wq�Fg�sB�RQ���]2ai#B�����vJ��c��8�FxEDbuÆD����e�M�=�����~�:o��0�����E�'������"�K��簱,�j94� 7�ä5���j���ޢwiwQ|h�
�A+\�u.ٸ�N�!�s�ք��W�C&���ܼ�F��4��Ct��7>(�nv����څ�]�j�ظ�����7C�G�0���d��\.��xD�0-m@v�'�-uѺ�Z ��f�t�U�ڝ,�q���-p�ڀ��yn���㪳�m.��$���h�l��ض_�Kεh�ڴl�e�W.��J�T�b;$���9����O��L~/�\�56���g�o�]����kJ��u��޷DL��V��#��*'Q�F�v�	�2q��$Uf_�G`��fվ�]1c����[���r�=����ݾGM���0g�kui񝞆����}����Ouu��'����o*dҼAC�|�^�X/"3�O�o�����|յ[����۪�
��Y�E�w�I�yϒ��ꠎ\}�qP��?�Q1|���Rl[�[s]�Y�{�y����s������\+�9��5�7�J���`lr�s��5S�4uuB�ٿ?W�k~{�B�޻yT'����^�ߗ{y%(��a.5�K+�����8�cm�t�	܎�=T�Т�>US��A�`@tB�A��2.�u������son5�Yc���i�j�P��I_U_k��1��_HD�VY�5�ƨ����H|���|Ry|����T)J�Up=���B����_M	���i�����o��
�nD'�)�9���b���o��$�dZ�}o/��/�#w�� ~)h�+�b;Է��&��z�0���I=z�5�V)㩋��QJ=i���#�CٹZ�nd�N*uvHw8��0.�W?[پ�6��"�I�_B�t:vK�. �r��[���l\���&�!}-���oa�}���s"5}'-c�ݷ�#yǣv�D���­X�sw�,��UP�=�B��)�C�vvE+fa�
X4�MGR���;�r���-�Tkq�ż�体��R�
0��n%R&y���VV�ӽN��3�?��s��t�>�yr��"�U�֟T�G$��͸�h�k�/�فkaӮؘظ��6�U��
�Kp�>��sVr�p����c�5�_s��df��1��ٰͅ�����r�Ulf:���]O_do=��{��p���w:4+�,�v��6�mVg$�IN3H��f#o��X2�S��k�%�=	�U*b��oDT��!��[6s�/w#}�w�]��*���=��V�q�B��ĩ�ӆ�󔡝�e�s~�{�?B�[=imP�V᧾�pu{�`��TV79m���:�q��-
�i�n���Wn�+��d6�k=��Z6l�z��3/�K�إ��i����yUw�߭jsרẸg�е��y����w^l9�H�+ s(���Dt]D@5�JW%/�k
�u9���mJ��nF��w��v��j�8N|��������V��v�\�bP���/4����k���G�K�8_]#2��N*u��h��bǲ�3R�����V���Hi��+�����ʝ�u�T�R���^8o.#-������Q����(v�h����Y�%v��(\�xR]�-��ߊO/�5���R�6s���u���V��w���w˧�I��)%��ҟ��t�8+fc0���fv5Uy��f�f���W�t��V��d#�7��B���+p$kf�ǛV�Y��f��3�]_	J����}:���؞��K���ƫV�.t��Wܹ�o�Q�6�b�!R3Q����N"P�9Gn+"��g����y��\�oy�֋�o�k�i�p�w�L'dd���oa�����9�����/#��/s/)���յ���U4�Ú�7Oټ���8�^9�,����'�H^?\��U��_b����w���]%�X�u5f[A#�Ӯ;lmG<��h~��Y�Is���v����꧝g�k�(F�l{�o�n^$�ݥ��-Uu ���wQ��h�G��i�$[ثXM�����z�(*�>�1u/�;��Y���]��^��
��BOj-Y����h�Lu�{]\�.��q5�K��W���6R�{8��֩F�_�\y�����N�R6��Omv�v�:�rᆛ�J|��
�Xdn]\��u�%�}�V����cDR�i�dRo�\��c)u�{�9 ̙�pZ1�pO�|r�u��w,�s�o]���b�Ҳ���)I�3v�Â�{{O^��[K:�"
тumkjU�T�{�C@�s��s�,�Z;�8�\@�c��rKj��ۺ�
�vlR�2��W�qˏ�&�o�m�%���l�Xl���Q���������AS��y���q��&n�<-�Sjf� u�17Û��6s;I#�n[��hQ֭MBm���ðd�+��k�;Jw@�8ꎂ�Z&�PN��'yE
v�TZq����"���f�h俬�݉��PadXS�[A�����pw{3�{�~��8N�5yYzԠ���U�%)�WVD"S2�NFS��1�F��K,���)��u���3d-Ztv�[�Ͷ�_�e uA\��Y�1���9�ħ`�F�3V���W�.�[ďR�jp�
b;���t�'i-�)hL�Z��}�?�_f\�h��
��54@��/�W/������C:�ou���2����@�-�ھ�C�{���Fd*dv�	���d[�oB��u�: y+/��X�UA̾�S[�C���N���/��T0�~Ǜ!F�Ŝ@��4�K�qS��[]L�ϖE��4���足B��\�n�έ�ɼ8��R���[��ՠ�WS�w�)ɭ�u�z�ub0U����M�>����B:T�v)����1��Z���(_	i�p}w���8sT����գ{�3XZ��w��,�E�r+H.��6��̠.;�u'�gv�ԫVJ��ֵ�^�˸J}���97��tt�9�
k�`6A�7��>��v�(u�սDq����'2���byE��w����Lft��=��٩ޫY�&���mj�2�=[[ a������n�1J��u0JqN�_LF�]���>��{0Ln�)�u�1(���,N$͖Uu�A��q��Q�\��㣂	m��Sw�V��]�kR�(>x�#��[��N�tY�V>��pn�Y���f�w�&��1��@�[˷�q.��wBW*��Y0V
]{��q״v��[�]�]Lp�/
�ڳ���o(,�H��r��R��
YQt�8���/� 2�s�.��+{6��]-ؔ��q����8Ӎ�;����@��F�2L�Ё���ݮ�W���O�z��R�e�@@Wsu���"�-�4�L�_v����&IL�c+�����T�me	V�O���z��{b�V���Z�_�������O��5��d儥AK���KK��K�dѓ�I���8A�Ca�Ra-�-%d�VcN��K�9��Hنf4�4d.f�(Q��ef8E$M���P�Y�L��ـdĭ%�-11ffYURS��Y�U�fEU%PdeNHa1���5QKC��Y�4Fea&a�ɑa�`dQ1R�RfefNYPUՒQI�$��5B�4> ��Vf=�3����}3�r���Pov�Yxiʼ���V����+��9��{v�,�l�Cp���-�vG￪��V�U�OS��ߣ&^�7��9u}��֡�E<��~É�]�f��i�L��W��k��O�o��ÜZ��8����g+�̢�Eom�N?�r�rUҼ�w�-�K��l_.f�Rl_Λۅ]�j�~��� ��	�eXݴ{�m	L�������iBW�Ҍlu���;O��u�`��͓�g�����b�ߩ��>��<�j\�+aj�q�����4�<t%
�]M����q���oP������ʶ�'�R��ө���e&�m�q���FCȮ]�f�q���j"�-�IT@���>
(w3ZRZ��rp�ps�k��]����g\*}5�O���]��6����}������T|$�lwj�tno,gѹ�۾4"��Gz����i\z�>��C�m�R!)[V�NBݣ����㥬�K�@��S���,䷆TriXo���
������Mg�t�^�����qn8n��r;����It*[w��a���� ���!�*J�6�_dO� �	�tgkU۽n���#�N�4�����eY��{i��l��w���l�*.��o����d�]5S<��J����x@x.�}�u�{�#�p�,�h%��]�qܝ>Ci.r���U�@�Kd&��[�]�S
�x:�X�m\9C�Ó�9ϧ��l��,��;)�Z�J\[LKn1���Tk�'����;Uه�ņ��f�/EZ���/����f�7[k\9���m7���g��L]P3��7d��U���w�	{DϡRCs{�#r��/yk�k>}Gr��;7X�el��M�@O<�ݧ�o��O`��O[�L�G>����3+�F�RZ�J.mZT�M�1���p;���SaQ1|���Rl_αmF���+�J�o��aǾ��j�d6߇[��_�_m:���_�\*�-�űr;�7�ɮ�[��NG�?}퍚�E������`ꭩsQ���:�d\����m�o'�.�Y�����[����C�����m��|�C����dz�f�o׆,��'�6�k�2��;.�e������X����Vt�Q�ǣrX'ܝ�>�<ylW�f��ܷ�F���Ob'��՗t���Ω�8�u�R4���j�=�{�坉�+3f���R�vE��ޠ��Y$3-�}YRo8:�UƸqո�93*r��S/�M�j�}��6��k`P���cNm��N^E�&���HY�y�'q�:�Of�O.9�]�k�לoT�&d�Tl�`���u���Ah���b��'ƾ-�B����j&dl�3��]nM��&��:tq�R1-���2ި��6�5�H��u	f*����E�v�K�~J��öf��CA)��u.���"y����L[�f�u�KM�w����H��6~�y����������;u|s��[#o���v�Z��\æ���bzq�Ѹ����ŭy���n*�r�qwK�Qd��r�l�[5�'SK9�m����Uk���9@۳
�[�+.Ocּ�қ�D����T瞗��v{n�s׎����$����n�iH�����J3;���ښ���p�^3���DĻ5�Z���]��l�]��������I���w7�[C��X����Ęk�4���oNw2��`������d;5��n�J�d�ޕ9.]�bʁ�����t��q�j��	����ɥB���Gqn�:�G�k��\�y�Hd���js ��d�ALZ���u��q��ܜ'o�h[������T<k���[y?\Wԝ�ug�sϖ��"1E��jU��	䃇Z�5�����6��히�X���{0�q���_U��¡`lo4ظt��ʻv�WʦCk��scgͲ�	���OG�:�aS�Թ��P��t�ፊ�P�\&�[��J/�:akG��*�6ʓr�������uFԹw�e)R�7o7��gCi�)U}H��4��9ɉ
���VԤ��u�w�᭮Y�����:f�ֽ]�)�T\�3�ond��(/�cBI|���%>;:��۪g;E譍Ԓ��Ic��6�3��D.��>,���)��C��1=��e�r�u���6������k <�P�9P�D.��ho�'|�2�dy2��Bnѩ}Z��m���Ж��p��9
����D �5����O2���q��+�6:�n���.\OXe򮽫:��*䮗7���Wv<�- �?�;�T_v�`�V��]Z���b�=W�5�h-�>�����K�-�Ȭ��u�k�m���5�֦�U�bl ;�3����Yf���Y�h�){+�����MC��;]��Y���.�l�o'Z�u�}S\��q��[���J+���ŞgK����*�\v:����۫W<}�����tX�7��\�����q��dd5���7��As�'2��#���#bj���{��ԫ��
z���o+���7���t.�Ҟ���c��͢	Vny8���Bz�8��=����O������ϧu���8|L�ql_��]ײ<����}�[��k�)�lc�]q	������6��ߵk��p�\�Ҷ��������*oх��.eJl/�'�
�v��{l����Ù��42�U�ԞqLjW ꭧSQ��+��X��DZM�;�J�W~w6,�Ս/>��Fxl�l��Ϗ9�yTmK��iAT��^�4��i���)㬻��/�]�}˭�}f��P���Tʶ�'��=WS��ѽ������&\��+��5����I=<SK�| ̓��OS)CO'K�I�ҬŐ�;�@���
�p�dˏ]��6���wE�n�F'E_g�/6�[�-'��,"o{3X�A�D6��Bٗ0BF�WJ�E��[�G��k;Z�ܹv�ۍp��F8[o�q���g�A̝�΅ªb����X���V��}!����5ٮ3i�9P�*�ALw���/9�|؝���i�7lV瘎�b}���w�s��C�m�aD��"�\,�T�p���S�[�0K[;+�t��o��ҿ�|�v�;����vj��t���9
�|Y�X��ٵ7��'{ӭw?e/5�����!yϩn͡O�=иR���S����&�Nr��ȫ<(kx���WL�A��)���M|�15	��q�k�9�i׷�D����!ǲ����~4} �Q=1bپi:ծ���mCyU��k�T�-��x�/�W���V>Z��٤����;=Ի�=��D�G2x�N�=�GhV�k�lE��~e�6��߯<�.3�O�o�����|���n�o鸹��/} c�
�r��o.��
�÷�v���LV޴:�e;��ox��*�,%6f�p��:�������F_N�4�()S2Sos�W��bR��B�ȴkI�(�u�n��������21Y�֮����'^GǙw����V�p�K�$�C�G�;JZZ8��p!d	Lv˙�I�7k*B�W	53@�
J����I�/*�!o���P��X��.�v��wy�|�"j;�U���7T���\cM�C���v�ؽ���܃��ڗ?;�dRGu��W�Zt�Kb��5���S��l�������e�(����bc啻�e�c[=q�u�_*U5�����Yq��ͧ�m����3�D������ǻ;.��B�c��T����_<k�\f��zuJ��ڀ���J�q�LH�����Z.4��9�.�=����Ƭ�u�V����֡*�A�c9P���-�s̈Gz���d�U{�e�t���Wʜm�wc[y�ȄB��h��}=+�,�cLp�%[��X]�cM�5��� ;a�7�1�lw)?����N��i�Û z�������]�i�ӏ4�"(8�mo��V�Sz0�r��^�x[Yb������ �t�����{�f�9�q��Jh<�/L��Y�y������ʇ[˴��������Pa�)�cg�fpy�Ur�rgH�9��k6��i�sB��7�q���0�����by�����y:���}��v��I�{;��Z6�9�R{9�:U���J�[P3U��c���՞/zg�w.}��\m�mUZPr*j����[�R�ָs�E�����'5�������M�v�Z�3������r�c�m5���������k�AL��ջ����[Tsՙ�o���.���Ss�{ìS���
c�2�̈́��rm�	֮�Mwun۳��esa��k�h��3�yV��r �n���z���+�l9o;�]�j�ol�DR�.��omL7�m����T��K�K�c��k/�����=�[QN�+�XZrvh���m�S�5Q� wΫ��ʥJ����7���cNh���a���Of�1�\[P(9�@pQP*��Id+��=�)<C�� 3Bw��m���"�M�:�^֚�,��B�B�%�gh���џ4Ւ+1�:L��ʘM�lZ��d#p"�������nk���p�d������q��O��%��@�b�Է� а��lPnT��	�6��!xM��k�/�-v3�H�wej^����볺�u�Ϥ�!&+JJ���fJ+�ہ��D�+��"�����nBq�O���3�]�v���dfos"D�s3�6��1�մu��Пt*����Cl�C�P
�R��03b�n�#ųY�	F�^Mew=����2��5a��=}�4����EיQ������G��0*�۟��5t�f�����������w�s�D䅵��Eo_uRGvQـ{k��-�ϲ���۫W<}��x�H��zɬ��N�.��Z*�����=�уȪ���NL� !�^���u�q�uз�,���Z����Zڞ[�> ����M���>[S��T6�OT^��a�nx����p�^�7�>���VOw�֖��9�z_/gv^cq�B�i��T	�2�TN[���u����T���`ǰ��g�U(��*��2���-k|�(V]5�����՘���qc�u'cΨB�K����wrC:�R�f��:^��^�ɹw8�������ԭ��5D=�xe�s �����s��tӫ���]o��gزH��K����<8l�9����Yt'E��v����*`Q�ع�)��w���7'�N�j��ÜC˯7�9����@�?������a[S�=ΈoE ���s)�t	���}C^}����`�O��Xז.��|�؛W���ps0;4L4:����O5�[�)�ޯ��@hQA�ڔ�IU}��imT���x���S�����F�ko�p���-�ID���LAQ�=nּ�Ypw��j��JJ��Z�>t�k��g;kV�ͧ��D9J���&㌚��<�xT4�4������3�#�-�aޭ�Ot<f�A�Z�{UGnVu��Fd��2c>j~[5K���j�[�94�o��1s��RnJ���(�7H8���[3�,�|
T4+\�����M�fj��봍Y2^�IRR��0�!�иR��Cd�-�ۮ{/��s�[����>�87K��D��3�u�M������
N,W.�÷�KWn�^�pd���ݮk���]!T�<ۥ�qP��Ю'`�噜�c���C�;6m���5�w�:J��wr���,jqӳ8���nwgB����3p��s����oQkiL(Ó�������t�MY`�.϶A9�t�>=��9�n}w��G�c�S��XXM��%	r�=�8f!Z�u3.���X9*�;���K[G�8'M�#i^'�z"��tņ��keQTl����r`�Wۂ0�̧��|��Ph�f�k�>���8�w`��O�>Qd9X4k�wmc�r�=]MC��^�`�#m�s�p!ؖ�E�;-Z�!K�;9��t��]W����ɻ�YK�V%�ĪW������v_��T5z�;;n�S�-�ýR@���+y�X�$˦T��v��l�K�����X��gs8�MZ�e�E�Qj�o6ŝj�] ����4�I���B�CxD��U��vXVe�e#��6�	�R�&	��z����iH���]ýë�me_σ��+��B�#��v�8�q�cLI��7S.�Vd}J�9L]�������S�q5{b�uoWO�g�X���s~�n��� ��6eu6(��pa���U=��<qk�Sg������--ܱh`u��r�;�����M�c���=��e�yT�z2�jS��'>�f�m��5�]�w{��Eܶ��\���š�v���������*_<;`�ʻ�����iQSw���-#2IB�
�Z<��"j�p�̈ET�'6�A5v=�� ���V� �u��YY=M�����C�_#�����xu!\r}������{���2^+��깖�A=�Ө�+]b���t��j;\��˼�on�8���0*:{�m;��o�:
j�u���k[Z��"eI���\n�u�v]ާ��Nh7�¨݌M���_E@�|{B��vѼ�X��T�V��$wu�W0�2�{m�Dn��*���Ɓ}f=�;H��aoV6�	�u��W��2�YN�����Xw�e���5G����9�{�3]���9ڊK�_1��.3��b�K5��]�y���L��3&QRT3��zXg泵�a�წ'�3���^^P���\�sk8�4t�3�Θ��ĕ�ˢ��X��y����u�w��fw���Ժ�`��v�tkQw+g7g:�fZ���Z��U������
А�r���W�X�8e���($JK`!���]^��d��۸,��##�K��0��Y����>YOn��ӵ��f�M��6���ŕ�r=.P��ǧ�KcUyםH�����k'GS�u��o��S�YX)k��bT@�h�<�!Vn.L�L��f�}y��5
}�捾���>�:���Y�]�7"��o�Iv8�K�]`������UV�L��4dc�EL�Jf�NVR�J�U��ad��EQ��dD�dQI1T�Ee�YaP�V4�1R�ba�T�fd4SUAQ,QfdDQM16a�LDUQfc�TfY�UQELFa��ST�DLDD�C9�UfbA5U1fT�E1��M�1I���Y�RS��EUTFS���YQFa�%94�Mc�ĕfefe4��Fa�Q%SUY�P�fc��e��D��Y2EYTUYLIDQDUSDL�U�Q�T�EE�e�L�KD�`�DD�Ewut5�����䛷�r�i���B�����m�uG��m�2�K�����g�'��:�"|h�Y��}˸Y\*�R;�d�a];���޸MT�LO&�]�:�C4_m@v��5uG��c��9Ʒ�e�m��n�]6�s��sm@�o*�ẍc����6[�������lRA�Uqv��ʎ��n3S�ܫw���q�dC�=�sl�5X-]!���w=i%RJy�0kφc��{P%`�����B�z�D'�F��"e��jfy 7�\oW�f�L����zr�-��\4�VQ�/�N2.�դ��R�;%�-�k�oе2\=.�J��~i�c��|:F�EJ��s����)4޺o\�c��M�o��wʁ��n�xڕ�R�~���XR��Au�ҽ-��-�Yp�|�=�[=�z��o�]��:�-�3���^�������+�%*g57���k/-���6�>�ۅ��dR;��_CV��F`
OA�w	����N��|Ryq���F���ͼS}̒#]ݖ^�\�2,v�SWf���%�^�1K__uފА;[��9˝)����6�M�(NX�,���ͩ�+L��ۅ����Ky��Di6ܜ�]�@�[qI�.	Rt+{��d@�R;�:WLF�]W���תu��^ͼ`�iI��*p~�~��g���h���b݉��t��-�V�㛽}ٝ�U^k�)c8�8�S�S�-�s̄w�<��3�:�Ŭ�ǡ�x.�.p�x`�m�S�g�D.��h��L�ZaN����N�q(Z��58{�i.f�|:a�P�R���8����*y�h���yg'Wu0<9<8�c�ǵ��M�MsLM|ۍv��ƻ"l:���gu����t/�'u��O*\�ٗ�S{7�iuZI���9����f���Mb���h�[��D�?{QiM��[��~��������?����'OY��}�T���ߡ�~ ��Tg�ט����.;S�="A|d_nXn+��,�I�����˨�9�K����9�4�"S�H�B���p�U�aQi�D�A��WZk��fݜ�.�Ńܻ�@�iX���sw2˲+j�� �=�׎��\.�Y.�?k�Vx9�����;���(��@ld��a
ٞ�dg��v��@{L���M�ٌ�ݫ�����W-�#1=�S-l5����V��R\�A�=Uݬ�t	����k��9x��Db|JXX�:eN�w;��z�W���c�l(t�ڮݸW��휆��e�Ll_�j:sM�m6*����R涔%z]+�cb��e��}n��� �~�Cr�+���bu�YU� 6KP9^��x��Z�7��{�y<s��}���k�9�7����e��P�N�{��!]P���Q�gF"�ZFb�J���n�<p�ㅝ��8�[�LwϦ
�b�JKC���S���c �����8θ����S�
�nBq���(�"�}�?HΙys]bl�jm�7zh>:�!��wQM+��06��9fQ�ȳզ�ij���i��J�,�棩��	����\Ҁ�3h+�r:���u`�1���|�>�l��X��y8�qO�S�֋o�y�f���:�˩�k^�v�;�`�UN"��o>�ν�sIg<��մ��5D�Ɲ��m�ڊ��L�r�EzNmr�9���\=y�(���É�;O��n�F�ܹt�b��)Ҩr���ptS>2�����V�{D�d�z��(P�CYj��r������7��f���|�J�Ղ�Oy=�W܍���wQn� ��Dn9�R)K��M|ۍw�k�3�赸2��^e}8��*�n���Y�Ú��%�ijg��k<�^�>�S�> �Ϯe������#{Ĝ:�ü�rd������ǲ^�q��Ϩ�e�:5z�`�:�h	ۇ�̥X�[�ﬗ�qm㖌}X���L�c!֮���ۍ�#n�L<���N��<Ɓ=������*^����x�M�t����ΐ�>>�S�R����jo!���;Y�����}]�
�_	�%���rK�ũ�0\��t5�w�L��>��Xד�Q�V[R��П���U��|�Jyc����|�=�{s']�B�Ӕ���6��Y��l����ѪN"���T�k�I�Ƹko-���_
�>�=�0'�Z%�55Y�C8���)�ΟHo�y�]�k�ڇ��|�-[���,<}Fk"�+�a��62�t�r[��)�2�롓ubR�]���+��ܮ�ͽ�V\X�tI5��Ǒ�䉩V���&����&����KtV�9�MYم����ܹ���^R��]��)\��㔈���j0��N�kr���e����v��م��ĺ�迳�KkF�j�ި��� ���w�q=�	:|ta�O9�ݹ�Z�1���%����H�O=����s�R�ɤ���NG]]�U��joE���sy��E����s]K�n>�Oq���B�n��-�ԫl[���|-�u����1�t6/�e�7!C�M��qY�v�R���_ػis�ڙ剉�Mƴ�z�2���N�s��m'�#���9�Q9��ugB�ē���E�V��[����Q�+�"׷]�S./%c�k��ZSk"[7��O��֟Ns��9�}G��{2W�G+v���h��3*
S1TD�ڈ�e�(��|���l���a�
3s`N�ӄ���Ml�ٷf�̢�`>F�d	Lu�Q��qwJ7GfS�;2�z�bB���;o��يd6�z]�׏���wx�f�^��nF�f���5U�A]���t�g���+��T!�F��̓v��g�!��Yu������e�v�uj��-駯RW�Y�1�9�<����)�a�LN��Cl��y��gT�f�烄2j����-���pt���¡TalrM�v�[�ݷ}7�r���d��7�U�^tT�a�V>�sQJ�N��lW�ᬸm�r��Έ�<ס�ѐ�~��{����{=*��R��M�j�8[_6����*�:fë�5�W��bz_�`t�T�0wsR�Of�O9�[Y�ਓQ�����trYQ���G8��()�L�Z/O5�������uqx���3���UCq�{�|{�o�<�?�ʫ���[��Qћ:l�,J�8㱍��4����06�5�3�!t��29�eP�ރ�VY�|��K�ջ�S��6�K�M�j��Cs�ml
��R�d��W��gu�E���ymF�[}3��M��h�t��J :'�u���fO.s��yUf:�~�,�,+�y�G2�c�8'���T7�'J�(��;���q�	BWc2�&��K��6�T`���8Q<�0�pu�B5�ۆ۷�N��S���f�E�4��}Ɏ��t-��f��t1:�w}D0��:,�w՘�L�#���&KG�
��xo}7�Xk2n.)S�������y�~��y��Sy��x�j�<�*;t�p*�;2�OR�k�z�!^6��1������V�ma���[�2���3ZW�6ӈ�M�)���j��u�^LsF�̯����^�q�pT�$PxYgء���Q��Ϣo�;�L�Ü[�&���m�̎c0�cb�nuE�ɜN��31�R��*���0�*9�Ö�v��9��щ��6��=SRu�1����:�6��ʄ��.��lW֡����p����o0��xX�}E�c<���@�:Ƶ<l�e�sm��/�
��V��r���ы���4�V�H�@j*�*ڔ�+���eO,�k�޵0�e��\'m�ж�q��JQ#���T���f�u�K`��ˮׁ�Mmj�������ۉ�m<g+�(�"���)P�]�Q�x 9ɇi��F`����M�y���}:�����obm��������-Lc�i�ɝ����)�X��ux���C��x_��~~x��nQty�R�D���9�ޞ��J���2:��ժ��n��y��h!z��έ��󱎊�^6��+:�o��n�!�RuA~��As�Gz�wYM+��,�<��7�Y!dU�zM�FL��p	��;�%����:n���\��o��f�Egm�� v!��s�eK�疇d)����������v��j5��������˅k��J���O�q
G�h\d'dO!�
��4R����6��f׳+�5���z�:�X��&�]�u���6)b}_D�̣5	+iww�i�)��EɯϿ=/T��R����}���*����2�I���жAT�{m���{mOV>O<�:o�ֶx�g���T�/�4=�Ed���E���OQ����c�#a��iv�Tآ���u �u����>�;6u��-��^��)ڳ����PU��79_	P��¢{2�6*�Ԛlv��u�i�|^e����U2o�����X�Ӭ}]ƘɘU���8=R�bp��U�@s�r����#���ή�����!0_'Ń���GMŵ��Gx��������1���w.ܻG�s�&8�s;���}��UξVƼܓ����xh�a0.���A�\zV4��5����o��'&���x�@;���J;���=���܇i����{l�Rf9�U�.@��ך^���ŗܺ�+�mc�����yo[�t�_Ʒ�>:y�TddL�=�V_%��5�㹍5Y%w:T:u5���\5��8[V�h��P�3sa΢�.�ƦW�B��9���b�|���o���]��6�x�S8t�gk`n�:��[O�e���ߒ�	-���3�����iXw�w�3��#\#5ԓ�j9T����,�"��F�����\��_-��j��P`TI��z����J�T.C�hSo"��0�=P
U�����]��TZ��֭�C�ý��Z�1��|�M�vˌv�D¤L��l��us!���&���`�p�O=�r㩽��{_.z�!�R�1<��v�����6���&�_m��q���U�]'+2�q뫍յ�Nqc�.>��m7���ٻ��y�Q+��Z�Ҕ�*J���2��	���y�B�n���z�߼��̘���E��{G<�w[v�G�ceV$���<�`ڑ�ϯd���/�Jܦ�b��
�!��B.3WCy�ؚ���D�nU�z������+��ή���Y�M,K�V9H�{����_�Q/2��h����[�^�|��=���e��a��P�w,!-	i��eQ��<��fr��|�!��u�WI�SV�C��E�.I��ݽ��پB�
������X��hn,�r\�v���=�ߦN�=�3;�0���� ���w��ے��m�]�q����ip�b�&�!�|�5�L^�ʊ@n����b'F�s˂X�M@�eN�}������hlu�ko\����l�2�ܦ[���Z����88����ڞ�u�B�SQ�ۍp�^8[gx3˫u-B
�M/Ӆg7�c���T�}U�N�jC�Of���3@[ֲ���K�����|�6�q�R�

{��T�Z4sWЎ��k;L>�6��=��]��<�\@v�q=�P�eD.�,��)hq�Vjc/��s�V/�}�9H
iӼEN��D.M.V��C�ٕ��yBLApԪS����,��pޚw�X5�Z�k&:��W[��5)��%�ج`yP�m��4�a��U�J�ꀻ��M,r�>p����]�w�vJ6��0z�s"#�ް9�~qf��M����N+�R��C�&5ֲ儇Zx�e]K�6���V�t��+�ʜ�l�@���ʹ�N�����4�J[G�3F�s���^��Tn�
n�8/&K9����ޥÃ�DXnPz��P�7�%���+����΅Z���Z�k�]�8������KTj��s���c{�R�ϣޡ[�ܜY�٫�fSBr�(�v�V:>����S���٘�2P�Z�d�Y�$�)im��WԦ�����M�2=��&�UI�r��ݝ��3�z[\-�b7W�_6�lk~�N�����/�iP ��$j��6�Ӄ��SNև�1���g����ᥜ��M�08��3.����Qj�M�Y!-�ýu��vs�ʔ���]��7�5���=wa�����Ч)���oF����2ʺ�$�oa9�(^�[��@�.�HV�i��Ks>{5o=6{�Z�EoS�Y�k��U���P�r�o�b}y�L�"�M^�ЩSF�GS�z�f\Ӳi�`�� l�C!6��V�GX9z@h��	�$6̺���)�q�=z��L1���1f�
ᴬwfwR����x+AKw�K��jy������Q�c��y���NgF�eN�Z꿍G��FF]��|���a|��F��8%j��Վ
��+9l�.	m-��+�Lr�/���x��IVekO�.�����/�Yyi���F9��V��Wѽ���e�� 9�Q��%u]1��s_N��]�&���Z	 O�`̽���w��0�:t����X5�믟 ��i�\�n]�v	 ��A�f^0�]I(����:�<�k�76�h+1)]Lui�۳3id84�AIU��̓��zuL�ʘ�\��}�¬0�ih/R��34��VR�4�k� ��i�w!ᕆ�՛qs�+��*�ب9Nb����N��Ոht�,L3}��s�P�'�7��]�y�5>�P��7S�^��T�gVr��u�2�5�5�x�S����n���gkX�*���ص$:�
I�lKTJβ����iv`�2�+y�����`�-�t������1J�>ĸ�#͠Lt��mn*��X�c�*Ř�������ɻC����c���
97<)��)�^w����̶���siDq�%w*������3�%S�:�s4���������VӊM�O2��U.��=}�d��tw;�����LRf�̱2l����YB�K�.Dy��r�+j]N�P#J�eP�z�q̋�
��rVG}��b�6�ws���-�mB&�m֎��Ijެ�Sl�S�M�5�Zw�b6�փ
��T��+��wb�t�m�}�&�A#�w=x͘�}���j(*(*�����"��2��b��0Ĉ��**"�f"���,������b���
�I��&"���(��(��&!�"
���*��(j����i�����(��"���(�&�X���*)�j����0�"�����"*���$���
����*)��
��+3�)���b	(�*�b����**J(i�&��(� �hb �
fi���"��i&()h�&��H��h����(�����$*%���
*�`�`��*�"���(�����*�)h�h�"���,�32�  ������fJ(bj(�j��)��2���3)���&*����5���߆t��Wz�������Z0'��kx>�R4�Ve��rr���p�V�I��.�V��q��ڒ󔭧�����
ד-s�}o���맼7�JbP�����N٘D.���ѳ3��4�F�����y�YIn�G���\�7��l;F�J�8SB�XaM�=X����7����r����o-��2��昚mƳ�6u�I&��F]c�)�n��6`_mrTIgyd��������TwXv�T���o�K��T�Qr�ߧ��i��j�)��Jg?8睝h�~�=4��d����{bL����^�W�����M �˭e��X�&�;\��v��;(�Ά{�c�u��s�2�sŽ�.����h�1w��,�y���V3�șV�x16��q�D�>w�Sa�-O�v�۳��pn�ӝ<�ؗCV���VP�g�~mum��^��˚�z����Q&s&�k���=��x7G��s�Սy?��w^�J�cb�-CX�ٸ�(Él�����븅r���e�Rw�!vj*s�&�����s�Ա����6�>�U��g0��b��i�dR�\l�s)3�vɋ�<M��@f���3��=*v���#θ�E���{Y)厌7��ݛ��N������Xi��p*��Gz�9\�o�=���#"n��=��;��ƵbGmn����A{ǱU�1�}���S�5���i���P���?APC�_mJK�lM��Sf�yf�X��S��ˎp��ж�q�R�H����;�i
^1��NU�kwƃ�-��mo\�Ƌ}���N3j!�9_C�f
���Á��'Ŝ�d�G>�ۃ@�����gZ��Ϲ�w�`y���s/Ք�G���L�ކa�3�E�Y��.���M��˚_�=(H7�wۮVh]�1eR��)f�;P:ps�o�z<.w�����N+]K�+~I��s���iRS\��ˌw�JvD�!�c�ߎi��<:��ձAj�F���{�����o&�yc�4��w�Tk�9�[��h��ҩk�=[���Vw��N]Eꆧ{Y�~�f���ڞ[�> �>�3���m��Z�ř�կK��0��䘏?� /��q:�{��Խ����$��G��9��Ď�>�F�A&���|eDÊ��F��E�]c�V��Vd�X5��2�.���<"�7���B�jv����۬4���ZVfr\Ծt�|�n:�����:��F��:�����'�)���7�C�;Yx*�a�̺w�n뫒UD��3+�`f*����_b��|��6�Ղ��םlA�ڮ�����B��WÎ}~��qm^uz:���|�X��k7[\�� ܿT��lo���!m}�~�8��o�N���$Ԇ�ԑ{�'������-�o���>�u�nl�����0{�7�KW�����ܔ����U�h��k�z[��������}މq�|-��5�.e��i0�7YR��R��!ө��'��X�mE�[pi#d�r�Y����7K��)��bs5�%x�]����o���]�/#�m�XV�^-w�c�ۍ���}�"~ih��_|��F'�p[K[��ɗ2CʋF�+o3�*��|�E|���,�"��%#A<�vT��P�U�u��������u��Y�溋48�m�AHs^���n�so�6�2S�B��#���[s%2��E�/,g��ŷV=�/��ˋ4���
��\W)�u�)�zۋhPflκT��"L���"Q�kh�SV�Y�>�T�D5u��kѤ�\�pV-�6��@v�n�~v̢�P)F��͍U�/�]M�s�kW)(⽕��ϐڈK��o�až�r%R&~�6bOX�S���Ӗ�]Jp�Y.
͚�ճq���s�ڙ剉��k@�:��w�i��Wy�������*�D��o?ao��wӻ�'ݞ�'=�3����V�1vD�e�o0�k"�P�U�*:����S��*��)}�����Q�L��ﯶ�?}&��G3������=Ir���r�T��?mߨ�vD�{�;��ĩ�J�->i��ݽ�F���
��l�(�GvѦ��lm�p��Ƽ*&->�O.������E��z�����k�\��W�LVљ�C��í����5q�¨�خI�ϝ���m�^�ʔڷ�ûqu��.t����9��.vTi�(�ب�e��\:O��՗Jf��qCT�fC�j�Nj�HJ6�kõˉ����k�����ws"����r��U��y�%̷0�W������ׯ0�T��{Xj�K �.���v����,�i�e��s�ns}7�;�Ybq�R[�t��'�K_K�r,[�	���t���.�+e�_Rf ��Tn�������ͧ��/��W#V�D���᭘�}����P(w0; �#�N:�Of���c��%�	t������Kz�c��\^;�iJU

c�|�h�ϭ�d�Ei�gg���}ٌ)�奔��S���C�oa�3�=�S�`�ӌ�\��fy��~��ߪܕp}Kxm}�V�x`m�lC�f����µ������;}Vl��7�w�o4f��&�;�;a�7��ـ�?��om�[�U2`�F�x羺]�q���S.��昜�����Uk�wڗ������K��!}�1|'c��mݮ��I�߫���f�]��Mx>!��@����i%]�\�e��k�wZ��:`Z�B�z9X�=�TW�ҹ5,y]�'ï�vU�o9k�=x�mCyUu��Cd\��\�-}ޓ}�y2�/To�+��%�Ơ��ZNf^��>��%[���HT�q��z�]�;3*�e�;��N�X�nl���4���T�[��Z�p����Stf������7��Z��0�k�M��>L�)�.�ʬ�;��kq�vͥ9oDˁ��Gr����F��ֶx�fy�����G�׳��`���:����A��B�;��]�M�W�w�E����D��u�;�7���^����@��zЩI'������e07Um*ہ*�����lW$طM��`�W��k��5:.�*nM8�c��\�����F҄��.���æT��n�k=��A��}:{'���*�h�9���'X���b;qx��e��[�����Yx��i����P��
{�2�L둁��hw���Ѫ^ۢ���1�ˎpֽ:vTB������N1���`��UnC�~�Y�w�Z�%>4[�V�s��6��9P�8�z���T�N�Ok�8����KZ*4����_Fs�)�z�<�7����w^��[��i�d�:C��E{5���|Y��y�#���Xx�=��Ih{+��$��wc�ҥ+��������U��:f��&�R��\���wKt)E)��˻F=RR���Ӛ��¥r�.���L�׽}�g5����p���3;�=��J%���̠�\xÖ�n�)�/;�u4[v[i�ݼ.��Q�{Ӱ��W/~�U��%�j�:���5Իgy<5p���\��p��1z�5�E�bS\�����@�9�rV�'�Nt�y�Q�be�u��n8׊�K�j#�9M�>F�]��h=���ך�W���1燼9�W����k&�}���-p��O���u2�`�~��M�\^JǾ���a�U7��u5�O�y��sO�⽛V���Ϋ������Ys��G���~��]�������c����no`PΛ��Gx�~�wv��?��C�](��c�v��I��YN��;$t���}�"�i6/�?[�nd��/�Cn�!�z����G:Lj��7g���x�E�	�g�z����={�c+���?x.@8�Ґ,�L�ÎHa�'e���Uv�Z��m�t�	��A��;��h��)@�������C=�vomD����IK#���F����o�VŃ6�=�Ph{��ד~w|��F$�NZ�M�^�;���v� ��%ݴ��\%��8�`l�(�w+&�T�q2�n��x��a���$�r�09�=)��SQ7{}A�ҥt*�П>,ocٶ������e�][R��PT�T�o7�᪋p�>Yv�gͅ��NeU�����������iIb��^�AI�;kc'3*��;6n2{�Ww-���$U{s)��.����4�Y���b|�f���4��=����
���{��x�T9����SP}$��R���S�	�5N�{s���Y{n��u�|s���/ˠ�������ә'�|fR#I	�'�+��I���(�wE�&��9�vy���������ȟ��φ�!��+�6�dR,��Q!S�m�w$�r���=�̓�|hoޭ]�xf����=oj�5�s�#=��G���u��'k�;�.U��k_#$�'TzF���Nyz(V�exwSm]�c!�]���P�N���t����/O��c�VG�Dm�⢆;S'P�����&��mM��^WC�u�pr�^Z�ˆ.}=4�մ�:Z�w�Os��zڨ8i�T/��Lz��j�P>�Ay<5�S�M���DL�=�9DK����c!&Ѧ[��R�AGY�V�j��P_n.t5��Z'EZKf)�=��EhK�m-��i�z{9�'��J��uъ�9��R����n��w��5�>�%ҏG�^�ow+�m���ѓ���N��d�����45�6nC�w�ӎ���߹�����!t.���O�l�7Bg�Qr;ѧy޴W��,���Ք�;�>�5-��lϠV&�.�e���;Л�K!Vq�D��r|o�E�s�Q5ׂP��?Q}�\��_��!����s.#j˧���\yԶs�}qݐ����wp�2���6�pO���.|X�z�3��.<2�h��\���:�˃=����i��=�z3������b��^�4�V�T�A{Lǀ�3^�Y�����ެU�`�z*S�n����z�1����}�Ǹ�Ӓ5Rp���8�24D�^��N��>�����,Tp�W�k����.�o���o�����m���d�q {��JBU�k��B*�����^��q�/���B��	�-���=>gp�9���L_��:�Ae@���wL�R�WW��yB,�}9��oL�|7Y�E���I�gS�e��-�=�|��]���h`k<���#ʸ2�}���j�Ƿ�e�_�Y��P��g� �q��P�n�4����`��yVڸ&�����7_,sX313x+\G]5-�U�f�U��Sm<�{4'h1No��ރ�15h�Q����/O���ڳ�!��fu;X�W�^��ɽ��d[��f�z����|)Y��|��%���V�Nl�1�܅��^,�o���X��ZY8�d>�Obhתr��N�h�u0�oj�VR�E@��o9��^��ĸ�(�C7�ԃ�Y=_@0��T�})L�~W��~竿g���Z����o����F�ڈj�ӈ�Z��(c�0V�'TGa����%�x�ڍ0��s�e�3Nƺǖr�����W�W٭<>�D5��o����4��_\�(��{�qnv��,�EZ�G(~����1K�l�^�f��h?}�S�5���T'n#���H�����G��"�Ϲ�nF�������p�b6n:������5��z#���������,����di��6�������R1�;*x�N홋�}���_4�=�;�^�-7��>Ԓ�����2�\(7����ph�����;�/H���O�Q�^Q��(�֚h�W(���>��}蒆�M9�úzD�ڕw&a�n_�Ú�{�VÌ*r/s�a �l�'Y@�!��T���̯tP[p�E=��������uA�9~:��z������s�r�+�l���[�_����]D���ǩv�ԭv�9��~Ĵ��vYc,�:���p��v���z�!*:�uuJ�ڻL+����^Ԭyӈ��Abl����b.O��z]����Y}�c��l��iڔ��µ�u|W �=���q�u\�2J����ڵ\(��i=p!S+�1�˸�S5`f%�`�K�1U��u}�:0;��m��f]�&m�L�lq�'���e�7-1b��G��qe��l�>�m�Y+f��Qwm�d�}�";K��nb�ʭ�Tz^u��������v��[����6tاwLk7J��ǭՅc;!ob�PaK�<�l�[C�[Pۮ�@�gV�Z��[h�ɶ{�HB����l ?����3��I)\vg*�Ɋ��kͥ�䯀n��ѕ�sG�g2(�	�͵yZl�:�<��%9�7� �!K!�n���I�SB���k.\�8m���]�㵅h����cW7>J�����W��utdF&c��T��K�,��C����-�4W�{mlM��R$|j�ɚ\�H�9S4uwɸ�K�kD�Y�Y2��U��2Ԯ+6����D������^��Sg3�`XCl壓�%X�ŭ�Rc�U��e��qЕ*n�2AQ�S�������8�4m�e�f�	�P��7�hN؆��\���]�T�uʗq�;6�'l `�JH%C]�����5]�۔����J�
\PU�E��9wuu�K���,Ȱ���hi��r��ݳ|pn���Z��ۉk�e�)NH藲��g1�Vwv ���/T`�Q�%p���cTX+.�]u���k��yծ"��[�Sz����1��>��Ծ�Ngr������T	��y�� ��1�|�;xV) ���a΁��3ѕO�xzc�9���Z򊁞,]h<��j���w;��˘p�"uc:�N���]n���
S�ุkn���������+J¬�;/.40��L�Yع�
��/��l��x�bʏo��y���A�Q�P�c��F/[�Hoz����S'V���V�>#Sc��D����7�M��/N|��w[�$���*T�>�����F ��ܪbݎ1���$	N�v#��
�	Jq0,6���B��n ��A+;��%f�Y�R{yٖ��â����Ku�4-�Nw����W0Ӿ�i�̗J���~ɪE�����ڷQ��`�fo�Z:����Jo��X"��T����G�	�ZJ�i��=�1�[*�73h�ン��V�h�֥`Vk�#�����etu�yh��V!fG��6(�H�d#dTEv�q�lV�wav��Z��O+1�jcj��m �n�c�/u���E+`��u�6$�z��}:|(�.����p�(���ym=u���r��꣹�VK�o)<��!���Mc�R������أϡ*�ԭP
�����2�n�rv�l�ނ�Y��qQ�K/U�a�(L�Q�᝴�1�8�N�ݫ�Z�ؙg�3U!QIS�EQM%UHU4�DHRQ�4�c�AHSQQAH�PPP�E��E#E�E--SA4Q�5CT��1$I�d44�4�%1BQ�4	��U$IY#@��L�HSCQLEUUP�@U0Qe�QKEUSD�.FEPR�UAUMAIM�DSCA0QY�SUT!U1Q1�9P�QLT�3RTTI�HEK�`ELDM%SCEIFY��IQAD��D�5CU$A3$KTY�A�4SIMM1QfES@QAU�4�DMQQ,M-d%4P45��~��]�<��;����^�b��p�f�z��o5�{guB�w6��U��9԰Pk�N��,oO��6�s��'�n���sI��b�b�RO���ԥ���BVwS��s�9���{UF3l���`LsS�7j7߬y"��U� �!OQ�y�2]g�;�[��C{η��b�Pv�M���q>�qG�U�o��{��8W�pA���tDĖ�H�|��#::�z�C>��l_SU)�Q��+/Wc��3�d���6k�M	\d�ZGr8H�ֱ*{KˎC�yF=�ժ��dyg��2s#Ig'c�:�/#�p2o�zt
�n�]r^K`(w��T}��2���x ��V�"#��7]���X�,y�Ax�4�N�)�E�*�R0dd�7N��}83�7&s�>�Wy���u����C�T�m�xk������᣿sh�|�]����d����l�fmﳪr��ފ�����<���C��}��8�̞�ؼ����;���"-k�Q��� ��]�7�y�ҿ)2ϼt��1�f�ږ��mr�s�f.���q��熷1�wU��yO�9��*������o�Ne)�Vt�����B&�&�٠
��߾ܮ��~{N��h����w�0g)��W�@tZ|ܠ�:c�-�����j�DM��Sa�$0�h͹�i��zM�ƮxL�6�nd�j����ʢ���&��X�êe�פ�mԢ!����Ǫ��_-�n�E��U �Z�Ck{KAs�w�*<�Br�/ޱ�{f��ͪ���3Ӑ��������dw���Ch/%f��m��p�3�B���7��P�"�6�1ﺧ���H;45���}+�}Ӓv�'�D�X3s��;�{wz��a���P<�t�*�q�)L���?~�q����R��:/�rI�qz%���~�M�F?h֢�L�^IZ�k�'gmʍᅧftu�l����2���5'b˿x����� ��n�Q�?��W�J�n�X������ޏK=!��7#�_����m���h/Gp5�7��� 5�X
^��=�>����`��W�߅-����oV�{�e?Y��r��>(r�6�T�k���F~?y��o�^/w�j9��\�ty����z7�ܰ���c��'�,sYM;jb�4���;+Dn�2b��Y�qZ&�)���c����c��͉�λ����ϋ��4uq�3<I9gt�!�a��ʏVŖa�x�].��-��/7��<��Y�ˍ��o�m��թ���Ěs���꺞��`���Z+
����V�=��>k˗ZYO�+S|>�wR��+ݏx��/O�xUa�����⮐��*��5�b�o��:6���y�|y`��c�l.�3�&�#��Wq=�wn7��f]�����۔:����}��m���"��2j��eESO
�j�=�C���Z��F������E�z͝��H��l֬���l�%x�6<Fv�xb���_�j��gu1��ކ2��-yaY�+�ո�)�U>��@��\TP�ja���*Ge}vF�	��[Sp�ו�����%�������!�$��桝��Pp�3��1��mA����u/'�z!��x�.2F��ǖM�i�uoiǹ$�lsC_K�#�.�Ew�$�,9�2��$�ޚ��3��&k�3��1Ʀhě�l�s:!��hDs(��r����Y
��F'~��D�Y����J=H�*��ޙC+�3��GZ�#'�N�.e�m�N�̸�l纲�f�[��+���9�c���XC~Sƀ�σ���,_��U�=NC=��U���N{���?�[|v2�)R�珳#����2�̃6G���}G�8�2I{L_]R�J������9�'��\�~>����v��^�X��'���@z�޶=��}#P�'
q|dh���jwN���IV������p]#`X�bYYգ��L �[+�B�l�"�/̟vNYJ�e����3��j���<ӂ��R��ս'��e�wz3�;���"�dȺRAtx��<V�0:%���%���GV��s���ˮ� ���;�{�ce�}4q��0�}F?����}<����/�x[Q��꘺�7��%}��SG����!j*�h����X3�au�2�~�C4���_	n�O�=>gp�9��v�b�+������h=d�VKi\ø��K �1?N] tx�b�g��ʣ���m��>ο3�\ݓ_6�\���<v���	�[5�ZFa��7s@!�����f1l�;�#,z����M_�\?yY��lc:�'~�l��ܢ��z&.�1�E��"dk��M��=��^��3W�c���q�1�n��e�Gޣ����;�C�i�A���f� ~��Qd�zT]EK��9S��K�_(�g��p7f������3w�[�R5��CT9ӈ��8�TV;H�/��l{H�g�]r�F�L�q?P}��*�E��+O�:�������Hl��7�QcK��W�.����w�yj�;���yy�8�"���R��=�١�[A�r���|5��������f/�/EC��G����Jpfn�:�<}>�13�ś�����jd߀�]~{A��\���N�۞�����=�o�����R�_t�|�[�w'��nQ��gF�nڻ�:foo�@�f� 'S��6�	�]���p9&`���dC���Sqk��4��U��|s��>�����OP����lgA��.�`*�V�Ǻ9e���E����oh[m�N�}�F+�YS���|N��fP�"­��>+�C�)�!�u��G����Ld.����(����?q��/�z��%�^�XeC�t���_�k�O�~��U���6u��xY���O����}�#<_�;�:�i����R6��x�I^5�C���б��(9���T����(��R�xоuC����}na��h7�¼�Í�����,z,,�@�~�=K��r�͊s������R�k�MT*�;����0�a���8�C�L��z�!F���U��n�J�H:}�b/Q��u���=ǣݔ�� �[Rݡ�>O}m�uf?_MX�VG\�{���1���uW�YP HzH!-�t���fx+��A�y�6mEr3�)�L//{)��{�S���%���M�i�(q��"px��^��}r��lQ�D��;�C���
��h��/�`�ؽ�c>>�"_�3��[sq��}�.ghA��4rLL�&�}q�$�K�WX>�Ǝ�wx�[���ބ.��Mnv��qo��h���xQ�~-z7Ӣ�3���������ԋ>X�1���H���l�@�w{P�q��:��ne`�)�Ϸ�:l�T�(�Բ*��H򞭻{�O	��;}.S�;>�T��D������7y��.nҵ	cp�;dM��ӻ:h��z�+w3]�����k��2��:�������z~Gg�G�f��]�(?7�H��d�_sj#E%0��;����2;�I���zno%�f}��l)���i�qZ��/�^�Օ	&����y<��F�N������xM��K��ߌ�����#���j�K����� ��7���K�֫���R��Tއ�y��y��S���3UD��Dǀ��>7Y;�����0��ӭqu�)��*Xf��}�׏��y^�c��^}�V;�Y�~��iK'v��<#�a�e+0v	t�وn�mÜu�q�]���ǇT�rZ��s�k屾�,��I��d�m̼7)���񮪙����p��ʤk����L��m2kzy���C�ֵ�հ���7�|��<x_��(l���ʑ�'},u	��3�޷B\�ݍTw���ך�]�峾���}�=�n�Y�)&�=��O���$�(	ȱuҺ�ȵ�Y����W����;��cn��	�ea�zY��C$��;��g�J(x��`H)zd_L��5�A�ǯ����(L0���:=r�kR9l/�Щqi^#�uU��l�7��/9T��':�B�}�����n��G ���:�֦��Y��)�	��A�dV!��^s�m�Ѩd�R��:��\��M���y{J�k���j[��:/���J�jp]��m��?��l��Qg)�؛6��;�\�iʌ��n��%x���T))k<_��_�5����	s�}��ey�~�M�}R6�TĲK� �>��χn���Y�G�[u�ׯO�QX���{6$^�]����͂�\���猲Ih����&Y�驡�{h�`{E��13��*I���g���a���ѯ���Y��%�O�=��Nn䙇��l�:o?ͤ�m~)W�|9�kӌ��W-½��s�����DW���D���6ԑ�<{s5橫�x#Ց"�/�I��r��;*%��=�W\��3m]�av�w��]�}���m���,���|�j��������j`������_Dݑ�Wf�����'�/MJs���R�ɵ��K�z1^[�^F��39���p�3�c��\�6����n�C��+��V��ܚ�_�J�,�A�l�9�+��:��9��9���s�8�d�.`u���r�x9�Ģ7��E�K��
ޅ7q��o(��ѳ�6T�%ٟ@��Q�{�������p�|�8����;��6*ZE�x������Bֲ�Qj�[�!��]6���r��!��9q!+�nĎu�K��n�OMV�DQk�؀�q;���l�\{�ѤhTD���tE��+�);r{S9)3��f�}G�n���0�K'L]��c�JL�]/���m^vޗ��ip�f�%���zuӳ�K��+��
����)���/�]{ǜxgk̕����ye��:3�K�Ոӽ����x[�V�	[����<^}��a�i�x��]tʐ���V__>�ь��j�+=t���1P�*Q�,F##�@ή�)-N|7�By�M�p̋=3睼���vS�Y�W�l��b6�n�	��hD���ĝFG��U���k�7{W#�J}���^�/ѹT��yAP��v}�a�煵�iީ��TÁD��H�n����1�a��Xی��1T�,��}��������N��3�o�Ŝ������W��W~�3Ǌ��֣۵L��EKF��>�<�؆g��ʐY�m�����;ӠlDw,��/˪��z�o�|cO�j���'�A��(�#>��2*:�s9�,7�Df�V�/ltV�[=�n�s����)��d#|K�5�ۨ�Y=�&az������7�-t�)c�"]�7�����)lۘ�~�T���L��r�-��4=���
R��d>#�0_Na�B}�p�n�o�͎ʰv���̧Y���SX%��l���G�"���GCLXg��#N��k'N��m�'t���vDr�}�-n;\����#6�>���gNN��D���3P=�r72wj�eY<G��켼Б�A)�������or�8waVr�
].��X�ka��v���O����]ӏ7ʑ�s����T��1ژ+e��A�vͬ[�;�>�����s�k�����{�����҅��U�ݍD5��-���TW�]��Qٓ��3�._Ff���#��9חEꗄ����h��Ô��xkkY�{T's^U-ֿdL�>���o�g�͝99�g��i���(�4��;�X��,�uO��xx�x7�Ƚ]���=��՜w��3ؽ�y�͝�O���� "|�
�k�|i�y��ͺ�C���<�%�26���u�u(n�gB�;�l�%��3�ue:�Nm���/�Lש�;'�<�=��=U�"ۣ�nr���{�VÌ�K!}��1uSĜ*N���y����_�L磇wG�b�R�S�,��U��Zv}���z�����'��xO�F�D�]�c;Sv�2�W�<�k�$ۙ�D��YIk���R�Zr�grv_���>����{C����@i�q��YK�Hׁ�|j6і�+�x�jw�[�����{�h�W�ё
K����=ɚ�wO��͌����AC�k���g���Rӱ�n�n��� �l��.l��}�D�]����d�ϛ���j�@����1Z|���}`�y/��t-r��)��Rb�#l[��ꃢ��3d�4]n,�9q��(QIԮ�;�����v�S0�e@%}D�I2��w�g����AW@y>���>�l���f:����o��%�B|p4Д8�f�����+��z�G��Z�p�*�ѓ�ލh���-���:a�z�>�7N6�DP~t%}�.gj�q��b��Z�6��>��S�>�>�W<�W*�����ۆ����z�>��|��E�î���;~�ݺ�����ʐ}g�'|&�\*�-�枳�����h��J<��[褠��C�oˑ�s�ח}[�u2}������\8ԭ:'_W���|o�n7�1���Ez�����h�G�Ӂ��_q�=/'�P�T��A�P2a�����T�N�V���c϶�G�e�Wv�3���U��W��}�����F����TN\�Lxk��'ް�hDݐ�++�n:�t?0���n�J�R���7�I:aL��g�Լ^G�X�9�d��T��,��a�S�~��Y�{��*�2�XYS�N��)�B�m��LxuO7%�w:�r3*n;�d�MЩ�\Z Dy������01��Pz��L�;u���v�Щu��Q�uӝ��<�Ȯv���n`�+�VΊ�h��ћ[��o�t%��5�q���u]3]
�Չض��o,l ����Es�4��O�	��*DoF$3d�Q6��B�Q�g\�|z��s�[}��X�Qgm��2���CW���̼�*�%�@�+|�������G�
��p^���[��W�e�ibG�_�c��9�j���n+���n�E8g;����ە`݀�7w�
.�hP��7z>U�ĭ�� �5�ZجA��c�L�ʂ�/Q��6�+(�3r�	��F%2'W`�oj�W�������k7o`���Ba�EȪ[6XSv'�E$�Y�;��t*!+9]�L�/:�0��ʄ(�����)V1%�9X��W�^���f
x��B���u0e;�X����&WufwV�0�]]#\�lЩ�FLW9����0�[n���Vk��X�t�v1�5�ga劷M��
�R�����wO}��l� w��n�����0�2>u'�� 	u��ܰ(5�����J�ok,��a3E��m<U��릲�&�\�-b�ؾ�x��`ƺ����,�[*�"�c�0K�:���.����+*wB�ǝ����Qi�P�Ď�y�f[\��
_@ƌ�֬�;&��R�V��u�����o!�`t!�M.���t��v�V�C�(�vu��!]n��)���;��]����zqD�&�|X�*�o:���Eã�&��w�K�gwp� w)r�V�U_}*,T�z���^n�9o�뤭��/�h�� mp����y�q��?<�u������~�U����E���c��a��]+�Ы-⮬@��ed�Ienn�(-�c�ޗdk�sj�o]���O�z�HD��:cP���C�y-7���u�dW�����q�1LhZ�5�Sx�7\�9��F��E�&��S�F��y���wZ�t�oyJ�Oo�vy<2���lq�yA%��θg�'4Z���;�����S�͙�WHʘ1����sFr�SYAȊu	��Ⱦ�@�����VUw@[�/��Pw`Rh�s;r��/4QLc�Q#6A��9�;�������7�l���٤�ڇ%�TV��s?M�7����Y�{r�g+z�=�ȱs4\�b��T�^]��Ko'�(ʤ�n��5�Օ�B�+u/2�-9-����.�R+#���	m�i.|ԣ�5#��wY;2g�j]k�P��e|5Z�ڈ��i�v#�Cm*yx��Ԯ�h|�e�s��u�tz�L��LYa�O{�0e;�������\�\5y&>���D��.0�S�/x���L�ǡ�;�AQ� )H�Z7��U�%�f���)FrW6x1�?`��Y�*�m��v��d|��ӗ[��VVJ�vÍ �Cf�v��rMB�=��!����wlV�d���|;*i�B��)&bh*�"���Z
JZ����ih(����Z*"j���()("����$����)j&��
(i�������"!����)����JJZ��j*��*i���h�����)
brLjJJ�"�(�JfH�hi2ơ��b(	�
)b�"� �������JJ���b���22�j$�(
 ��)"B���Z32S(��(�&*�)J���i�()

Z
)�)�����������!"�
��	�������
(JR�
h�h���i"
fL��(��r2�ƢZ
2S"�J�(
)"F$�����ȪZib�
h("h���
i
h
)j�!��v��*�i��ޙ��x���K�׊�0��M>�ɛ�V���9\�vu�|J�I&e���Q��\ᔳ5�.uw���C&�{��T����q�Y9�<��~���[C3ߑ�F��T��l���szQu9��R}�$�9��2�jE��'���Tw�����3�:�Μ]�NMu�>�s�BB�b��k�a��$�,	ȱG]+���Y�n�U�����RW��ҥ���x�H]��5� ۸�^0��F��%Q��)zd_L����@�TB��=u��.3�B�'[����V��i�l�8yӨv.K5�Ua���q5��������;�F!���$^�ob����=���9��u�Sz��d�8��;�I%�z�G�m(Ύ�#�=yL�2�z�Ƣ��ƴ�m�f��xj��n�"�����m�m���8�nq\�rs{�WzIt}�8�H��
��i���<��e�2��y����z�F�fKĽ5�7y�j�㸆�̊��31�aV
�s�42��5�ʟ~�_{��7��s�V߷{)-�L����1�H�.���x�Q��"_�Bym��s�4��9D�[�p�e�r�;0�:������-���m�������j��o�˶.��یN	�{{�yy's��6G��pߪ�.Ҥ�u����;��c���U�N�����ʴ�gJ�ЛEe(��wp^�yuu7�{� �z��InҨD\o"�q!�L�����H��;�_�?}��#�l��y����j`�����;.&썤����Ǯ�T����K�ѥv;�<���m8Ȭ��8ޙx}�c����zfFG{*F^�'h�%�4t���.MN����)���T�&π���{+iǀ䓾���45��>�&�Ł�}'�L���y Kw�v}�������*n:���_['ML��k��K�d�q���p�#מ���d��Î���#��L�rt�>�&x+�Yᆝ9�}�eӃ�<˃Z;�ڡ��ڙ��Yln�Xq�2��g�{H^�)�B���g��U�7�[�������-��>�U��zj:ʋ�^�+}��]�M�����5�!��:k�<I��̠g�����?�Z,�c�ݸ)�,��,��;�X�1��P���\zؖ�ۘ����Y6tw�%E�UA�p2h�������lYLS)w���@�_:yAT�~Ӑ�#�{#}@>7�U#nS��]��x	s����;�^ UϤ���H�2�x��r9��&�޴�9��9�8�	ۗ=Bx��t���1�l��C��+h"�����H��/Kބ~���n�����37󉾒�]d�AƵ��qsadv]>̢�f��f��cW�I)�Z�3\:fw^�r���3i@�HN��A^��6�M��[����<�wl����ܭ�rGZ��ӛs�"w��ު�C�g�?�e�6�e�K�s��~,kQO� �%��1����wx�#��}�<�)�[%f!>`rL�!�'�h��#���eEmr�r�ç�F,����{d�~���Xر⟬��ӌ��5�ۨ�R��1��s�!=��C�=�)�{�(��k���`���1��LlW=�Q������~�`�� �)d�@2>ʍ�Ґ���1�%1��~.���l������})mD5�8�/x�TV;SK%L���qۥ�D+���-��[�/���t+�WR�7�=����C�;�V}��C]>�ߐ9_7~�ٳ�\�(�v�۞�U��e����A����ڋ�����]m'�����}��<�ϴ����W��j�Z��R���m�16���+N��K77Q3���·'$��4��;�����G��ne��32�7ю������Y��V$�`�K��`��د�������
t��cc��t��O�a)���~�31�ծ�|�6s�Kc0������<K�����3�v�|NC�F�h�"�%?���le��!�Jr����'%ye^K�[�|�� ���j\~������u{�Q\I�N���hp��:s-a���}w˻�*ɘ`����\�to��z[56m�eb��6�r[
Cz��M��?�=s�(I��w��.1�iG*����V�<����E��Oz��K#��K!nyL]
�$�"�l�K�#ҽ��pΤ_�Z������R�x��U��Zv}���z��L���s呻���Ł?≕?N?�����g�$F��t���)f�t�B����0��v�8�+��
r��E_����1��cq��z��lT �2��W���e��}}K�M���-��Ƿ��yB"'oB5e����g�R�xs�x�n�����@%�D�o��%y�&g��8u�Y�·���i�<T�`��z���������%�B|s��<V���p�r�]D9x܈�w���s;�����u��,#B~t��%���ɿ��W?:�e��3����d,��s�V�=x��E�u;�j�{Ѕ�v�F��ԁ�x׀�f�
��93J�]4��ʋ��Ӯ���`̻4��!/��ͣ����5����R5�\�%ڈ�*j��� �ϳޤ����GG�2^L2����=8���������^���U�A�2,�MMr�y1�T���a<���L[�ր��
@ԗ�7rW�&����]\����+gG���eT�B�ܥuo_ e�x��$��pɘ�f>��{�a�Jގe������+���wV�U�À�����G:�N6εc�Z�n:�͓,8wQ�9lk��X]��0�uG�v�^����;��@�7���U���٢��$��uם�C��v5���r�z!��|j�wFF�"n���y<7����й��U�v��`;����nyS��jٞs�u�U��g�!��1���n���w̂��������0�+4
�d����~��T�r|�y9���+�gNI���Un#x-��{�Ta9E��:��ڤq��.7���&�ޞe�8�!v��CҹN4�k=�/!�Y>��U�I�2�9ᔓR(er�鯯���-84<�3�c��!���g�+�Vv��8��t7`�(m�EE�H=FX�b��u�J���
���y������h����f������zߝǸ���P��(�2;�[s8<�0�*�Ϯ��q^m{WQ`��~�Q@O7W�]��lcQg+�kbt�s�%�D@�0ĥ�A��W��.�Ī�oVD��L�]�3M�&������'�9�œ�ژ�itJ2zs z~���E+i˃n�����Zl.������g�C���ٷ/h�I�J�.��7DZr��7\�Q���YX3y�����x�W�Kr���=��NL���B��:ɳ*;2�b �5�u� ����Jrq	�fjC��]������k;4Š�tb�ǒ7�b�z� 9���k�5�^�w��ٱ"���/���[6]���^��]��T�'���R�-#.�I�4T�4I��KkaV��9cL�4l(��z���|���݆|56����nv����?iv�A����UߧÝ��=�B��.5�ʟ���G���	/lѧGsٷ�w����EnX�~⇖K�Pd��2a���-m`��u�5h{�j93���F���d�����\d{[�Q]mCR�q�k��Ev�
�d�H�zaK�,v*��&�{/��r���EQ�/�v�FFZ��>�I���P��Pl���CT���e���L�rȧ�O4cֲ�FrG�����C��H�����R�o:��`䓾���}>�	�����a�D�����.g�]�۲���r�ٺ�g|Pf��6l�d�=3����.e��S|p��B$���=3�V�y�l��c�.����W~GO���KGJ���:�r�g�-�B4�x��+�gR��~�u�����ƤU�\)C��#��\c+�g�S>��n�.��\f�����F�H&��ݔ�x�B_h�h7VD�9��T;[�zJ��t���ۯ��E�\�g��Z�첵k$♧q@�����WWF�r����b��Ϋ��yi���o���nSwҐ�A���>�bgeL-ؕ�z�"�K��N�mf,��Nԯ+�ꇓ�a�G����|�l=��kCs�t�Yd��0�AR��&��
�Y<��<�K�������@���\[���Ge?[�9<��(��(sY_�`x�ۭQob��� ��w�}T4��[�a��s���Q�U#nS�B>b�]Ϸ�-h��W���� SRP���Z��c��~Ws�ZG"��\w��8�ă{mht<d��[[���#%�Sɮ3]2* El���n��2�X݆g��|��/�ف>}���c�
�7�ޫ�ԩݖ\ݓZ�	�i30�d��I�u2W��T�x���΍��1����}��*��~�훦c����G�oh��}8�y�Q�9�E��&az��b����g��;�R�5Nc��so������c�q@7�J+_&K��."߾�C�s�H(�{`���ǥFSٱwO��,������8�/(<5��y�T���CT9ӈ���ʢ�ژ!��s��r�y�J��_���:=���*w�ܾ>�c6{}�P��U��v5�O���=�^��^�*�����Uz��=��"\o(M��Ek4���S�0��tŖ��J�6�w!���:REe(d���*g�gH6�aX>,�-��/�H��S��!n���9����:��Q}b���m��;58�I�+�+�C],�7��{*��7��<�����?����ٜ���(�,-����VW��+����ٓ��˭��L�"_������H^�\�#N���]���,~fl�����|?F�r���ү��}��
3�s��&େ}�׌t?�%���K8�5Q��^��~Sf��&�Q/OE�ZVZ���Ą�K����.z�td��:�f=ծ�:M��R��>�NG��l�%��ZNs�
�:ʙ���tv��k��E�r�}�0�����t�s���s���M��27��*ĝZ�f�23�$�,I�(�6�ʔ��\O���{Nϭ�3�m�{��8�Y^��Y9�J�D�ޚ̵	z*��l�I�3�=C�L�K��R�:j�P�O��3�}�{�6Ϥ�W�'fԯ{��=����k�]�q�`�_( yW�X��2�c5�w�W�HJ�7�&��NgMkٽ��"�#�$�������=~�\N�z��v.K4���|}DLIo����W�ﴋ��^��<z�v7ؽh!�K�쮌����iۡ6k�����w(�$x �����7^��2�#�G҅�:�?{������� 4�!X��Ż�ݫ�\;�6���c_$XḭD��k��g�7���;}�z�`f�CQ���))�}\S�������Y���*���ã�띅$���u��� q�:b|ַF�DJ}����9̾��9��h���>�"}�3��q��D:hM�˙�g<��g�8����'j���<B��D�uz���������1����6��̧��\BJu���~Uv��j�kv�̙u6M��cME��W
�KY�|3g���yA��ԙ��<ɢ}��Y3U$�k�.k.q���uC�ɓ��*h��Ӂ�T�:.���^Gu>-VT88_�`�d��=�"_�ht�*�e��s���z')��40�3�XY:�d�WkC������Ň�Cs��,�Y�^�`~�Wz�����ޠ�/b<���Z�(Z��ƅ�����־���ɍ�X<g-�-��ިJ��|i�{�����<9'X���ֳ�|�3�ӑ�S1^<N��m��Gi2����z�|q�Լ��N�;�)�B��~��y�=�t���|�7jr8 ��>5=�z>^��!���z_�z����0������(haw�]2o��w�6y7hm�z�ٿ?*ė9��~����ߔŁ�=�	�(z�<��z�/�З7�VO���+�k}��W{31ʊ�Js7K�wߣ�=�u<[䮵��ͰIj��=q�z�A[(��#Xaf�:Y1���*o�(�g1z�xu�:cR��;2+*�����:�1ۛ�!N�m
�8�o���Q�9Z�Govd�G]���mV�%!}w��.�{��|8�>jS+#��<� ��{�v��e�0�b���g�V�.�����mM��%��6����w.��1��/�[Q�(s�<�!ع(�#�J�`��T~\&G��Z���X�V�L�;�p�K~����V�ޡ������t�����DolQ�Uǌ��l[�ɓB�sK�P�5|�����4�ON_��FA�S�X������>�����+�yU�\� nO��H����G۬�r6�
����o���al������('�-ڛ���[:8�@Fٝ$�����f�I��ԅ_��ö��~�*95^�}�X�g�>��^Οc&Ͼ*q�f�
snfE"�M|fF��^�=8ʊ�r�+�f�á]�FW��U��wg]�9�c����[,E�P�/�ICO�=#���~!}=�W��q1�<�G.�z�e�u��
b�8�j�:=��W[P��n\A��늋��� ��*,�����!��Z���v�8�Α��l�ʝ���m8��T�`�I�s�p��p�~��Ǭ}���n��7��$:j�e�j����;x�u���̤q�|�%m�{k���ӭ@Ik��� �o[��4����dm�[7�gE( �&���Ǎ��U���2�LA�u�u����X׵���2I�ʱ��mg�>Ht���,貺0h�>�\�� �H�hrޖ�m��o��K������#J G�����ںC.;y�3]�1�;���!�)���y��,�S�89��7)�krrG9��AVwb��v�s,=_+�-�8��_)r�����J�w*��R�qͭg�i�[׮�k^Q͜(�Zu�f�RP��ڇ(cl�9���<*���3;�����/����-�gCb��Eq�����F�K�}`��#��������3p�ѹ�;dT�hu2Tv3�����v1'�@���[kn�>C7w[�r�r��Ǵ1Z������=usoa���۷0%)��QV
���ˆ��ݝ��9�I6��j�U��r*�J$;��jl��l���b�չ��3N����J�y�)crV�4)�])ڬ�H� T���u��Q�N��|DxJ�%�ET�;;�ec�X��}1�M�ͭJ�%p#���{��d�jn�l�Ֆ�۩���.���c�ٴ��-N�Ph�SF^h];���|yL`�ܤ�p
�[�p�H(�f�ȳ�¹Q�k�r�jھX-)�����T���N���GsX���!�؋K�qyX#�6m��Y>���#����{sou����^��L��4Ev
����i��8���t��(�WuF���=3��ѫ�^�t�q�I��.C�R�l<��87k;$���Ee��u˻�Qe
���1w��(F�n��_t����2:��D���o)a�&�uǝ����kyb�ڈ�D$�>�Ƶ+�������*���Ҷ��=��}����]N�X�V����/,�Zs���u���v��la�]Oݪ{7m��e��2\��\��j�U��k�k⃩-^��j3r�����ǘ�ʱ[ɑ��Fa�*�B�a��"�+�&F����(f��>\p4ep�I`əD�p1�n�Ⱥ�"�&6ҏṀD
磙+��K�=�ΐ�h��Z�,u䙶خ��iWB������t���c�+T�>��{3�խ�S�괫/E�R����F@Ն,�J+��|���-�8���Ou�4�J��w �V���ĦH�u��^t������H��]��X�g�v��U���]�nU�굹3�^�S5���Rv�ŝ�!6j�& *��:�v�gEF)ϔ?b�U+.�t�Qs�>��u�wx:-t��p��ݡƏf�1:K���'��:53j2fQ��vq�K89�ek�i��������˔�c}�J7�'ma8d+{��V�����\�3��i���Y�+\��1I������:���b�Th��|�U���lؘ37v���T���}�5CIHW�0�����ih���h�"����hb�" ������(h��
�����
bih�i*�`��bJ�����1
��$r@�Z��)�ir�(���Jh
)���H��c1ɉ����j%����l�2h�)�R��*�h$J����J@�J!�B�hJJb$2��h
h��
P��(2\��Z*�hhhR�2$(�hB����, 2ɤ��h)H�*�
h��
(b)�h�
��"�)�

Ji�"
h�
,�J�bB�)ZJF�!�!���(��h"T��(j��������X��i��Z
��+�@���/2ż�P��x�U��1�/6d��nЩ$[u�ڵ����r��{�Zi�3`��v�jJ��m,2��`�(����������h|n�����K�l����}�S�䓾������ϩ	�O�N=!Z��y����9�9��4�#�C�ʮ6jW�GI�=�h?K�d�5�6�Z���R2�N.	)�q�o+���Yư�&t\/Iӷ��Bg�����xIr<�F��w��Gt!�֟+.�������l�C�qݎ�����A���c*�.+)&��o��Իg���2z��x�ʣ�,��Ǹ9���i��t�{�5�-�)�Tx����R��N����Ԟĥ�s��:��������˩@�Kuq�b[7�mDv6��F�6*N�\�\��Nq��[���q�rI���u��������PU=���s�=mDvv�F��-��T���O�{9�`�
���>����Ԗ��q����c��ohM-��4���Y^Y[��s���^�J����\��4̲Ae@��"e��o��7Y�F�*A_��P�DN�d��;�v����=�~t��svM|ۨ���U�"�s%��S�I%yMV�x�z�?10��܌��vgH�gܪ1�m��_ [�4i�֥4$�N@n)I���݅q����}֘�Ps���ࡸ�HO��ݛ��N�^*�f�n`�s��_v��+�*J��#�N��\W��s��/�A����}9�/W,��;8r���])��z�[�A�� ��Y�k�����n�iK'��/_�'��{�m�3��O�x��x�E�NvJ�٫���0�C{T�_K%��."߸��G:S�g�½D���zo��6��?g~���s[	��	�����8��*F�[QP�N#詠��v=v*on���5صK�x�=�ql)s�{�||��)|o��ˆߪ�����S��3�����&�3`�H�;��ܱ|^���O�F�K
�·qY^p�v��fO3C.���(L�[Hĩ�&3o/��bU����Ez<��z��Y���������Йq�����>F���M�h���D`�g�����;�<ꟳ�﮹��47{�8�g��M�,��3(O�b���c�'�',*��ja`�#��i�/oV�1�ծ�:M���[����_g�٠(�/k��DS.�Nc��cX�/�8��䑼�Q�(�E�F+�<�=�=��]�����p��ӥE�E��Y��OLy��$�Rq�gPt2�4heOD��ᅧg���=~�7��[�5{��V�D�>���Pf�z{�|�ǽ�]�_�����{Mޭ�%�ۡ8$+��啥���������{VF=�x���o\������r���xR�<�w*}Bռ�$*of$p2��G��8�q��w�PJDsnN7z�#5)���-����HD�h�r���}_)`��2����C��n|6]O��MT*�O	}��]Z��*��{.(ݟw�3�U��3���liAʌ�!�9e��k��ej���vNwL�>��{�x�Q.uӋ�~k���1g(;t&��LÊ%��A*>�&K}$s@�c��Hc��Ϫ|�F1��S����_�2[���~������&�v�M�4%2Y��@o��nj1i���m��r�rLz"o+��m�Gݡ�s�|������ޭ%���q4�Y�=��ܠ�ؘ,��W���52��1�5��1"{GQ�6�6�3A�B����ͭ���)�E�xA�����w�sg'�z�+�4��R�ΖN���F�K��W�KǨ�)|nyA��#(��lqޗ~>�{{��J��g��ؾ>ٓJa�5%���JӃ~����y���߮l��s�F�2�����|갏v0�4�D�7WF��3����G�vЋWJ]��*�5fpʨӯ˃���
�}��)a�;n�xdBt��ñ��=oUD�Z�(Z��Ƭ�7t�t��-�R�U2`��wWFNe���e�BiwN5|���ZDOy!L�Mە�s�{�M�C�g��d�aę��_=�����YԷ2�os�爹>i���8�6t:��r}�#���86[�z/�\����o,�1���uN��Κ}/w�We�}�;B�+/7L����B��پ�%΃�i���c�����Ox��V;�Y�~��w�*	����?I�^��Z���"�crGZ�Vh-����"�k�Ǿ�nO�!o'_NF[�g�M{nĖt�p�v�����;\�Pۉ�a�3�6��R42��>>�&\u|,�ɭ��^k:��]=;����v_���c�r�!v�s���Z8%O"N�K��T��U���
\�zo���`��=(��q�6�x�[�.چzϛ����P{�f��eҸ�7�z"`�=���4�V;h�wI�2s����m�l���B��ӌ�a�G�[Qǭ��{�ߌ;%<I@�3T�u	��j�*�V�jC\�̏GL��5�A��~�QB{�\{��㷍E��������8"x�=��?M�l�^x'��/#���@�D�}2�z�Ƣ��\M���Ϡ��#��\8����j��&����X��d�q�q,
�9(1�P=&'��\�h�u��F�!Q�	��#���Ƙ��x�~3X)U�J���^�'�_�{V��<f�̒ѳRٳ�D�/ԅZ�h�e��y�6��NDq�iGR��
=��)�)t�[�;��V�-�l5[t��Ӽ�L��c�\O�Mo(.�sݢ��R�>���������Q�g�L�B��:K�̕Z~.�u�ؔ��X}T�C��[����w�B5c�E�s&��S�^n�P�e�����0H�RJ��b��Yȃ���&��snfB�际��*�Q.{ƅ���q�3��z��u�{��^�٘��=�DP�Ί-�"ގ(y}��d�4�8�zGeD��e�:ڻ<��T�s'Tu�˰׬ySO
�b���W�uJ:��S�ˈ9Z�qQC���Y;{���5�_�=��ѣkf��+��vC���x^���"������=>�j����.���d�����mY�}�O�?FΓ���������O��{<�em8�䓾���}>�R�fL��e][K�}�4�߾�))�9������N�q�eW%x�9s<!k�=Ug[32I��P��{k:ra�XڛӞ�P���aC��f�ɳu��G��������x<�����-��u��
n=ye��?DmG-�Ƶ̸>w^���ڸ��u��u��߬�|�b���� V�>R-ݚU^�ٳ��֨g������Zpb�����4��:[=񚂷���H���w����Q�1�a"���U�X��}�'���P;�in�f�'�;�������9s�N /+��_�뿕����^�YG�:x� �A6��ƫ��vgcÞ�~�#%�1�6�E56��������g		Y���\�Z��>Y/u(v�\�v���s�r垢b9Q��B���Y|�
`�ۺdM���}F��<v�4��Kw�U���Nz�f��g���N0�?���z����_��[�i^#�u���|M�6�A WMR�x����#���d�@I��x�-����#���&��=���=�u�����\@"��%v�����<��#;�L�$r�>�s��q����3<��G��n�f璉��Y�X��omG��t����˛�i�BrU~o�Aג>�U�A���~���ui6�u�{Ӳ+��E�i�9={��t7��t{���g������<!ur��'�L��v�LMC�7��=����r�f�s$1=k�T�d������0�IF|�/���}TE��LUw�sWDw���z}.���/�3��@���.������v����T�[�������4s^W]�T�ѓ�JG)��{v���N�>��,�m���6�axw���>����]�9Mtc1x$��Y�$;��cs����Q��3V2\(�z6����������N��M�]�]�1��{jMaX���{X�I��������O_��4��g
99�>�·u9GG�3�ϝ
�%�MS�۾ԘJ��T��^�*\ž���vr���nD�۳ҰV�*�T�̠�LťS"���W�Ō�Si%&Z��,��{ ��E4,C�� E탻�9���N��}gk���+ Aз�,<#;�u�Np�|��ll�3�����,q?l��_��8�%����g��3=��B��<<f�W��v�nznO��0g���o�,z�kM�� ��bv�dc���I���[���g��l��{8�t�)���Վ�\̍�r��ڤk�Q�(<�0����:���VÌ�ɻ��������t���藐���ʩ�N�O�L<����X�_:�k���r5�2��`Ȑ�{�
Y�^�����/�gT��NW`�)Ol�G�C��n|7�S���Ч6��Ęv=��;���-�;>��H�|s��z��j�}�gp(T <��X���-�:�.���^A�D��cڽ�-aas[By֍��|_zF��o�'}2�>%��A$Z0xS�vڄ٬�5���٩0���N�3�\k���D�����5?Wq7��Л4�BP�'��ڭ��{*�3jˬ8t���:�@�&
�ts��>�s����5��e���C�GM�q�\�H�yu�J�:Z����g&n�f9&&^&��=�j�͉c{iɡͭ��#�9�a��5*�zs�o���\t,죂��+j
��W�:�����YJe���zR}����B�j�^�$��!R���Ro�Ηu�;1A&n��8[of�v&���yh<n�s{hw0���Ήr�\���o�(�3�"�4Mt��������}(����A<�;w�,ɼ4�-�"�߸��pB������xW�e��gЧ�\*�-g�l��(:}v�k6���E:;�νӯ�`{��(�m��g.����2k�0ʚ9,tx�{R��R��qT3.�ez-1i3UGۄ���]]��갎�%���q��lavg��\2a�����љU0������wU�ֳF��ۦOwJ}�z<1:��}��yꨜ��z-~S�_Y�n�޷�^2�5e�;~��7�)�����V��~r�"���Òu����k=��Tf���ߜ���M:��It���ωݳ0��J��eV��Կ�M0Bֽ�<:���ԏ;��Թ�3U�f��������gX��3��ݹ�KL�4g���ꑯ���>>&\uYi��7� �t��i���ec]���qK�.+Ԫ7x��^����ē�&v3��2�jEe��\Y�τ\�d���U�-�Z�<�3�|���:�|f�����rA�2��|���r}���K��8��=�Q����"�}��B�i�Ű�c��6���3L��'J��:��YYl
���O�,��Qi��]���]�=���մ�ڇ*.t����D�y�m������n2h��G���f{�^Vޣ�@׮�>�����:E��O^��f�zu�ܲGVqnj�k�����uG�f�Ḙ[��.
`f��|0���/4�G��K˝�HߦE��~��wP}���[�`���1����6k�!�-G(���.N[];bwr�3���/Q��%��hdβ�~f����Q*'�X�|^W���Ѥ��N�	����vs��'}��d��v�D��=5��>�&%��x��C5��&7�?[g`��,��ѵ���~�ԫקt�����^��~3�d����͞���^�]�#/L�)�c�n;�/#��uy�]4hs����%���]31_"�M�^��K���Ձ��o�Q���\�s���;�k9��A��Dk�:ܱ��/�_����'zGd��]�z��W�M��Σ��_���i���xf.��ګ���T��mCR�q��~���v������H�v�91���&\l��;�R�Ҩ�>��+��q�y~	�����2���zT9��3j�N.������%�#/����ݨwY^DIzN�R�n3�_�:�������8��F)�J��׌�d�����Ws�>���C��ӡ�L��5+ģ�2�t}� n��*zS�FQ�g�׷�:j��m��l�ٕ#�Y6,�n�V��*���qn��j�c�VP"���-@t�<J��,*��W�J��Kkl����-�v����Wqέ��u��H����LT�iݮz�=;��K�Ң�#�tB��<I��LL�7��aڛ���ݩ����7}|ϝM��|�f�^¼_�n(rl�}3��9YI�Ȅ�Ǫ�Zɧz}R�"�tm�⮏d��莫.�ֹ���l�-Q�������VY>Ve��7,p5�X���9�@�����5�&�}���*;l���pk��4�� �l<��ݶ���+���'K[��R{�w��n�,�-��I�;U"{>��T���X��O�w#}@>~�=�\�ۼ��|.����˸N*K*�z�z�P�]@{z�f�<��{����\���ݎ9C��f�h�t�;O�Z�F�*��6JD�;%�?���l���c��~Wq�WN��X^�X[�n{����_�ê=��q����s �_(!_O���[����c\ޡZfor�����z����t�c�y�q���7d�П9�f;�$}�Qj��CY%]ڧYKr�`<W���c��R��b|r�t�o5�����3\Ok(xB��%�ђ>�����ED��P����p&��ݗG~˖�k9T:֮C�H�橒�9`j��?}����
�+� ��+��*� �"��EA��*����"��EA��W�T_�PE�
�+�
�+�*�`��+��T_ꂠ��4W��"�� �R�/��"��"��b��L��x)�Tg� � ���{ϻ ����u<�>(��TT��H��R�I�4Ց� I��-0RP�%!�٦�ٲ�ͳ}k��L�ڵmI���e�m���IB��4kA�]����=ޤ���SSLA���B��V�Ġ�a���X�j�K5H��wO5[�>�:z.j�wc�E�an�	f��ƒ�����]��4{�*�Q-��H��ow8��u΄[d5��{�  (  k   L���rti� ���Y;�k�;� �P���Ŭu�AC���D
�Lъ��v[��B�F��5��Z�R��x͔@��t�7Z��ͅf�mX���͢١�Vc4��[x=�^�o\+Ѝ���C6*�M� 6�X���4:�dk���v:zҊ5�Ӷ�͵��0x�]{f�^�()�w�*l�Z�fà���F�]w45�Q٪F� �V�:ڳV�mYmU�-��l)���c�h��$$u�eY����۹Ѡ����-��� �;(���m$P+<  �R�v�g�J��wf�鶺���
5n�º�փ�����&�Y`ւ���� 	J�6��9�"�
�)U'Fӹ��F.H�ֱi;eC���0i�X(�b�k�9(����ݎP�*�]�;a��  @ Lb�$��F�@a h ��{C
T���FC  ���?�ɩ*�4 4      j��	J�OS 	�  M0�# �RDЀMi�����'�f���F��P�J��  LL� LL s�\��;}��;r�-t��Ҳ[V�g�$����,�$�u�:K �H�@\��Z}j\����n��S��?���F�~�n*"�(���$�TYCa,��x�2J"��H�9���m��ȧ�ӧ��O�ȉ :�m�r������T��A�&'����pT?Sp��,/�7���W��C�j����8� n�%��y���S6f��Eil�ZX0ތ{KFm8���D�:<�q��Wl����Jt=ڀa�<�Os�o]�7)Z5HY��N�C�V͗J���Ñ��ܵ���P�.h%ؒ��M��E#��%�ւ����$�-Ю\F�I�+Ȏ�fLdn�fL<\T��$��(��I*�\��
<��j��b�E��� ����B�!<��R�[�1���3c@���	p�^w���z��tU�S�NV.�]�(l�k���Զ�s�uR�]R�;P�B�;1��"�6ܳ�3hUM�P[�I�w��6�8��o3K��<�1���5[�O*�����v�@��
s�3���t���Qr]��VE���gB�lc�ÎpK.�ks-�r����EP�ۼ��j�	fXa�SC@�ڊQZ������9�[8L)�+�(�X�^�W��X�o�rs/dX���� �s�[SttY��UV4C��J#*�ö1^�Z�YJ���Y��U��J[��6D�2X�*�m�4V�%�/e��l��@;���m���]��Tɰ"���ۂA�X�
�^ڻ�����nF*K$œ�����[q�4���6�n�z#�]��S�3r=����x�Cr��CUMP�+#x�U��B Ӈ)$�)!��U�1٫i#��,Ց��Q�.�Cd�\F�.���{J���T��b�-ʹ�l SJ�"�L��9y�W�y0qF��ĚD���lRn�5s�R?��f\�nMo
��a�z^�{��n���{G6�$��^�ɩGbϰL�i��Y�%A�
vi{;��+KBk�/&f���f��S�S܎�,���s���V��+�ī�;nn�!�tf�0U�Q-���v�P�ڀ�Gk5P�z�#�O�8�Wb�#�ֲ��q�|�]�^���5C�&��ps�1K����:l(��&�7m�'vT6Q�7Y��p`4.�(�[X7��탕���>������beDN�T�����-�m�(�"i�Zz�Ym�61R�dW	)K����F���gqc��82�召�pf�]�~U3!�+�;S}��ӣ .��\�9Z*�0Gv��V�sC��KI8����<��s wR+��5f��
��Q�Fj�J?Q�@��,ᰥcȵpL�����-��VEl��C,L�k+���$�L�q��k^�y�̝�f���ah�!IK1ZY6�ő�+��J�#E��@�vȰdu�Av�Y����*`���U���l��c%��s)��n2��S�'�u�h�v���WM��r����[��"_Ń�[��D�[5g0��m�mÙM�ʥ�%����q`�w9�x���b��i�H��w[v^\e�}^���cf�X�V�$��2��#� �Թ��~�J�N1-�.�5A�3U�&���]��F�V������:���&>V��;��ۉL|2̢�n*Д�Ȟ�eS��NX�лJ�;��T��,�z�2��q�45ٺѸ����^�Xu�����S��hoN&��̪G�ސ�p�C<���o\!U��E�	!75n$�0�8^��z�_�-���Vr��Sz�8&�s;��Cg.$MӖTM��ݒqP��Ĉ�-8��OFm\�C{
�̴6N���(������0����X��fL�M������	��Q��.�0�O/J�PL$���)����{���sf�0&p��MeI)��^��l\�tٲ:�i��#5���H錮�[�/v�Yd6T��r�ˈp��{��z��g�Lv1ב}+=�>�-�ݧ[�M��.���K�s+TjS�S^��5cǝ���jޤ?�k����6i�oV��`"m%���n������ђV��I1vq����v��&H����Q;�oqz�	�7����ĝG�ݽ[mltq�!LSD��Z�t�]Z�X�ۻ\
��{-��S�Ȗ��R�����Uf�)�m7V�m'tN$��y!��Y�݇IT9�t��˓wB����Y[H����TV\�$��j;N�?fӪY�k�6�1�YX�T:+3mIX2E�,4�9�@��t^]YZ�LGo1�o$ļНKg[�d+��_�_����T�˴��I�*.9��q�eI���U��U�.o�y��R�Q[�v�Q���-�I�v�i�%)�{l��D� ׎I�&�z5��+�����v+ywMI���m˹�8���q���ih����&*F=;�co�jۯw�f���Y��5�v�dD�O�s����x��Y)S�a�w�FΦ��Da�*�6��&�y3�L���m[��+�6�n(:�3@�t��ΫX��;��qg\t�͌��tpq[7�V���
4b�Zu.ob*N��#����k�5;�PD�̋>P�ؔ2��V��On��2��V`In	�r�+ȇ\�I4�6��(�rä�͜3oS�B�J��`����)f��Z����g:��Ÿ����t3[V�e�.��nީ�%�F"j��:ީGiɡ~#����4��z��v䚛���qj�h��5��R!CX��3y�ZyKkVP�ņe��巕	2gM��m��v��2�<9d�j�VE�4e�ci��W�0�m5�h*Ff2&�kif�J�bNA(jQ�9Ya�U��|��9L��Υ�֯e
0��SrU �T7��sX���fj��eV�Z"� ;�Z��]�gS���`1��{F�r�)F={,CR�Z?f�M����98�my�$�Pk�W]c	�	Ӷ���F�.;'[u�m����·r�3�ݭEVESp	�����8�\��
���*��w�F>^]6�q��7��[����`ռIZz���:�"�W7�=:b���o+�k2�{��P7��⳱[����2�2J���_g\�$ZV�&��Z$�mԹAx�w'1i�Ӵ�ݙ���]�BHT�J5��[�%e�7E�d�	!be��������а4�y3:�2����r��:��J�UjjP���@y���R?�}�Ч.�&�S�ojU����vs��ok�����6U��g�ٽ�h�)����Z�B��t�B��y�4](�i:�N��s�����:bu:u�n�t4�	�4Q�x���&	�+�!R'M��2Q�2�u���$�E�V����:vh7��Å�n
I��*�њ�AQ�xA�j�֥�cUwX�����Ta�5�B��rq/;�T٪u�.��7Y���ت!$W!���b�cv�<�6ED����-��c�"�}���h���!j��m�l9L�o�b],���H��3�[��0-�#��J�C"�y�UF�a��������,���t��0٩�����{��C��5JyV��w���V��YH�����
HnU�n����l�"ve_�^Adٗ��w7i�!�!s4�M��i�/$+<s:B5!��N�$J�B��t��*��%�g�g����YZ
�3�,n�áI[���%P�z����;ePgH�Q�
*�Q��X��έ|a���e�/}r߽'���֝~+)�*��i�/;h����߶�B�Z���F�b��:�U�u���tRLA�z��ə�.�9Ϯr�5������]�f���A*#R�Y:�����P���d���5ܮ�����R�dN������7�5�������c�$���
��+m(V�~�r����%9��:�����\�	�:5P�d��c�b��Ė��W�����_�^�,&���	���5VZ�t�}5Q�<�Y�G�zf���TE���>CH�z�N�܆�Ӯ빜�#t������Lr�V8�����F��1�폞�j[V,"#w�Ԧ/��{�JT^X8�ז����;��ޜ�1�t"�؏])\4���ԧu�s�h�[���y5KN t���_(j�7�P��`��.�j�zQ����>��|���5�5�i��$������ۮ�;��U�a\n1���%��w�6!�5PH�E�	��t�z��&��ɣ��Ztt�I�����3��^�l|�LC}g{V��Xݜ#b��\�K��Z��ޡ�.����{BP��R��O�ޔl�Q�Z�@ϗGK:�J�k�QڼqY� "��y�Z�maJ�_uc�	to�5D^2X;��eDr�i��+-��*�wfV�J9z�KPI�	ݪ�a<kd�, s����t�#wg��ݽ�gUj�Y��@���۽r�F�w=��'��!�/
�J9)l�]��=��}K.��L��X�d�M7,r�T�+^��i�c�L�^Nw�G1�w��q�Q���پ��C�0�=8���,��j��f�N:�;)V�Ȍ��ܴ%n���F�$��S]�lO��Ҟ�R(�-�x@T��D�1���"�Z��o����8����{j�p��q�u�lS2pT��ԛ��m+�H�e��۲���&��.|u�x�
}���x6�=�,=��s���ʼv̼�\�wT9rgX�j��2m����3�);CJg.}�Ȥ]�v�\�Ă-뻶�9gf�53Zf���W�r����Mr�x��-6�{�4h�3\�@v�J�u��f�&��J����^L����^���ʊr��3:b ]�:T2;h|�T�΍dĬBw2��I�RS\r9yY[��a�y��5�)يv�< 8&�R��תT����o��V�y�͵�cgc��q����#�E�a˗ǙB8��G/f�|��6| ��;�߄��h�M�F��Zȑ�7�_D�G& �q�S�ݪ�Gr&h��:��V/�����Q�i�H#���*�Fjm��;�{�X
��o�.w���sg�N$�:�����`c�v�;2�f�Gh>�z�������V�QѴ7r�.w�OE�*�{o;^>�`���"�*������bg�یu����Ԅ�Da��^=Z�Y�m�ׇ}��@�@���ܓz���3!�����G;m��3�E&6&6�,���W�z�v#9xhţ`�Hq��+)��LHMp��7�5V9j�u��t��Ƶ�1���ټȑ+s��m��"�>�T��wD���Nn��6��/�RF[Ÿ6��rk�f����`�̟'s��~��"1��EY�.9]��Pa@��m�v�f�+��pt!܃��zB�i��� [�v8W]�R�8�v�����=�J�����=�Ë�U�5�nZi�i{�L?*�iޥ�V!��0Ѳh˹y�	]�G7���@�&+ �dƪ�Z�b��T�#AH�y�6����7Ѭז�-��ό<� h$��Z�ܵ��/S��j�賘L���n슪:���.��*�Js&��o�3�GV-A&ha�+ �(8`vu�d�9�������4���T��[D�q��P�u�z�ɼR;ў)]����qe�6uo�k���wW���U�Sv³�;�Ewqk��8zU^��G��������"�^��D'1C��X-U�����7��	&c�ͼ�P�au��b��u�Ivv�QoJִհ3��o)��n�ٚ4�ى:��&Dɩ�
<�U11���� /w�����w�2��w�Ãn�%�V2����c3�^��C���r�Si�D�M�=V�����Θ�ae���.�r6�K/�foK_"	:�P
���y�~]�]�X��+Ե�[/�`��wHU�{�Q���S��r��q.�C����!�6���s�a�5Pʤ�.-�M���-d��aӾc�W5�n�lr�$�Af����).�ݿ�gygB&�Y��}�V�㚤K=|;oޓz#Q�7����SLkX6L�svr���W;�t��L��J�����;w2��+p�I!S�A�<Gw"����f�u�,m�_t��6d|��q��o���(X�SNgO+��ȶ���,�ɪF��� Yf�k�}�2ޱ����u7���۶#�lz۵�to����jZx�9���	"����sY"�tV5��4�C��'���0gIyR�7Y�A��P��T�l�X���+��Q��u���h.��ge��bP������}.�c��Y�A��U���
�ˮ�ī����vʠZ��=����xd�&$A���Rd6�e[(��×��\o�F�a�Kn_V���Rv�jWJ��=�%���c[G�`���8Cj�þ�� ���RC�:�����[�H�2��l��pB�f��2���/�Y/Kt���	��H���^�PkSoG���>U'/�t�9*J�
6K���N���A�TnF�2�~	L��9j�x�ᳰL�cV�#��n�G$�%�2����Y��ūfOV�M.n��j�݋������;�hCyVrr���3�n�w��{Z�;�P��LL}�wWR������n�����U��r2�;"C��f�=�q{���Ӿ�շ޻���\LTY�H�˕Yͮ�mb����Fq�v]�]p�d}�:Z�GUZ�v�c�)P�����fŰS�����4��v�%�}I^�(j
�l�D�{bkޗ{՟7Ӣ:�ڙG��FF}0�Gf��|��|�+�Ԥ�z�^�O7�]�Ss�ٝ�|��v��9&�7F�Z����L^������X��'6r��y�H#j�tϮ��|�M%��B��������Aӥ}�ĿE���l;Y�L�O�L�;sU鵎��ɛžN����h>�vL�n�Dd��-����V��XT�wy�й!�ە�Ye���Kݒ%Odfd�=3b�"��br`M%&eNI$�I$�I$�$�I$�I$�I$�I$�L��䙆8�����]%�A��\���Nt]�3de,��3��ԓ�"�LeGߍ��Vw�E�A�i�,���seE�8��:�Bއ�h[M��γoyȶ�9�4z/w,;��37�Cz���O?C���C�Y�ugRy�n
3u�X0��ߟO��-?�"O��=|X+�r�V�Дq���t�A������(�ۈ����Q�ˠ2݂&(�d3tp뫡(����8]�M�2�% s3;�ڪ�!���fv���v�t�G�Gn.��hvwś��FG`�V,f^/�a:���tl�e�Ύ�3�����	6#{��[�UK�;$9�[6"6�;:�o�m����B�>�&����8�9'U�:��mXF�p��w^�q;Վ=�:��e������2���7Ltڿz�뒞~d)�<STBr�q���Pt��`9��A.-�Z�R��%�N�+��9}�5%�Z����������O	�����ώ�*_�"I ��W�	@�ˤ�ڍ�7)j��d�$���/�E���tP ʟ���n�=�7P"��(���^'y�7���,�;�c,�,K%7����v��R��ڢ*�W�R\�i�o�so�|{d�SVB����&[ffcUT�#u�i<"���`���iF��)U	�I�6�l�-�\��MyC@��~Vַ�''�����4v���k���c��b��!�Ku>i�UK�n�|�Q={�RyNN�ؘ�E[�3�Q}�);Vl�
��Zs:�%U�NUݪl]S,�!�Pqٽ>��Y�YF(fҙ��[��x�����n=Y�C��ǶxI��s]q�rdVRaZXI�(�x�	SyEt�b��J8�nC>��S���:�Á�����Wb���p��i�Kղ
��2fy��%0�6��R���f`#�F�1�H��Ö��`���H�<:��q��I��ok����7�2Q=u��:��"=��J�z��V1k&���F�f+V9�E@����b�^P��bZ�*������_z��5�+		����o\�%c\V�+F���\"�@Y!��ⓚ�Y��ea����Y�$�F'Ƶ���,X0r��,���yV��k�}�MǏŌ`X�:����fRq��h٪��E�rT���)x���MK�v���}�F77r�����[��ǀgY��~���fR�y��%��tS�<Xr��M�`�Ҭ��
�ڼf�ΐdO�kq)HJ�Q��6c!�zt�w�T/z&y\�0��1�.��'�]o��X���WT`�Am`�ɚ�y��GIfdT�Y&8[!��*gY�
��"7����}�i뺾���F�w�s��r����7V'gu�H�6�`�����Yd�cqV�7�/7O2_������9���v�^�� �Ow*1���D�$�C1���mB2�}{6�\���.�>/�bo.EY�Mj��Għ�}���a��-��n�-%��MB�t���,:ɈY����N]L�1WJ�C��g�NU^Zv$��?�%l�=+c�ٺv~�\�����hy.����e��
=�»�l\�)���Ѷ�*YfU P5�V��k�w!�@�y*�>S��9���!�(��3�^��V�W�$-�2���/��(�g����#�]M�AkHx:]>��jt\�S�.m��J|Em�4�0��ӏ�ԡ@�iː��l��[����S�lPUE)܆Z!&2N�۸R��y5Mitpۘyse嵸jM��w1K�6n��Z�]�Qdq`�A�X.�|�DNY����!\1ee�YyN#��_ْ���+w�lAs���ё/m����]m�����Ӻم`��(*g7�g��R�� ��t�)���fW���d���0�<]8 ��q۩+��2*3X��n��A�8��d	'�+�m��M+������%�����ZNG��s^��NfP<�Q�l��{sC6zUʊ�ic������{]|�t��$��?u�������?L���!Ӆ�c:cL�e�V�mo�7�\[��k�����]B�M�Zь��ê0B,�o{ĕC�&.�9u�e�U/��:߄{A�V˝��,S�L�\7o	i�4PxT&�Hu,��Q�!�,#u#`�+�KoP����#>U�Sʲ¼3�Mp��|ql9&��/2�6h\Cqk.��ϯY�g���(��a9th����6Ѫ���E�i�hۦ�4"�s�'�Ě���۔;Ddᚿhc�'N�EÍ{���F$y��ȅ��C�z���F��X
����°�4sǦ�-/�Z�J�[%U,��j��é|bn�a��QǠ1$�3��T��g=е����aO���|!qZ��1�
��%�B�h�Ӊ�p�DBpUA�K#�ޫ�ʹsk��֙�C*�Bl�UNRI�HP�u)�tBm��cv����v�4Cd�Uvƍʻ �M3��T!2��*W�+O{t�TC�#���UJⶰ�|��ӦQe�4��&̫}��7p�A���y۟v��z[�R&7e�7�D�M"�;0�2bϊW��� �m�yPP/��{��C
9B�"-,9Zkj��'�P:�b�}�l�{,��d���4�L���O���62vH�]�N�CL5r�uu*�Bm��@��;,4�X~GXaL˚,3����%�N*��RYw����X�=�}�BC�#�N�DF.M��E��*���dVUIN`��A�,T0�p�uuU���S��>�YD���PZ�3,�]��N,Pռ�cB:��hI+ݏ7���������m��1�*�$ݜ����X��]��!+PL%�DgE}�%l.�����%u�IJ�T����T�����c�s�j�&���R�ER��â�&Μs,;��Y�7��Êa�%쮋e�\��R�̄&lʬ����iyo!i�%9i�KdTV:2�$�:sYx�x:�R1Wݎ��Qט̘\���h�D��Qu�eUE酏�r�o�L����+5�,	(�kL��a*Wȝ�J�AU�AERV�@<\!+|ar�h��]b�|�n�ag��v�+8ͩ��j!0�}���{ �V�ZfG�[�nF�T�T)ړZ$���r2��/db�A8�A6�4�̭Գ�b�N�b�g:���KJ�R�6�Ʋ�	��kh@�hGNcybކ�\Bb�ܪR���l�.O�K0����U�xZ��o��r��V?�P��Ή���(h���m}ט���jJ(E�s��J��2�[I?�kD�K�����R�$�lQ������F�����dƐ�u�Xz$�+A�v9Y�d�WR[�]+/p w��,>��Hc竰���%I�H�v���o&D�3S]�I��\"����ԋ��L��7��R��1����yB���n�R��]d�b�ς�Nǚަsu�	�=!�I��׸�����/������;���S���f�����0�Y�䬼I�2��nl �i!��V�-�~��������8,w#y/\K}Ow���}���e���l�+�x�,�O�-���%����22�J#'@9u�V��ג���0u/
�P ����b$�s��_WȌ�t��)�5]7򿌾7tpд:��P�6��#�!���d� �;�` ֔fE���*RPIU��b�,Mp[[�GJMqͱ������:]��%Fsozt1��#�O�m��p$�5x����7�$�{�������3	�U��#y|(:T�!L�(�+�j&�j���X��Q{p� �s��k{��M�J�t����:�<9%��{�R]��42��,��RZJ;V�Ja�C!n���F��`�m*����	\/ ϐVZHL[��r`�G��=Qѭ�d�"!�h94��];�)�ٳNL�GcsP�ςKg6���;��ud� �<ΰ���H���vRq�{��P��$.��.���.��x����*���^*%V�)���\�؜��	GЌ1��S�k���&M�e8k;i���̵g%@��غ��B"r#�ަ�X���[7W �Ϧ'sw��e�5�2�l�c{�c<��+oNI �E�_߁� #���p��(��,���C.����1�.M���D�0IEF���6����0���w[d�������=M�.��f��Y3qU"�WՒ4���ѳ&U���v
�U�o}��mt|�f���yL�X�\�@�D�Ɨ��+�´������s�v����}��B�)uj~���V���Z��U�y��b�oF���3L�V�����������s"���v��gX�OTX����չÞ�ܟb%o,�d���J�_V���I��0ڦ/-/=/��t3��#�$�g1Ev/�,�Bd��R���A}B��>ǮVJ�_A���k-��[X�l���
{�'°�1^��˾ a��kA����1{�<{�ݍ?����Ό�I���?x���}��?">�'��B,�U"Ł�X*�Ba�Z�+%@��*a
��� �
B(()!4�A@XH
E���P���J��$*T0��2�D4��P�`QX"
(Ab��T��f�,���%�ATP�����0�*2,�ʒe%fm�b
�g���گ��Ϭ��H�r9�]���	؎�4�\w>��a�(ҝ�)&�T:3���_W�~�{��k ��wܲ��zrﵦ�K+_	J<x��1���w5����P~�#2�H	�iqC�1��̜��P��˟]`&ᴣhل��'�{w\�e�[�=4`T<�[D���_3{�c�v�
Z>���Ϝ��`=<Vg�ꂨڋS��t#�%�"����,�w�~7�J�靇:��;�_�o-B�q։�
�1�b��	.�g�K���B^��'Q��f��y�Bx��~����C'�s:'���J�wφ�������۶��4�v(���HFv�&��w��ʏ�obI����#}%k��*N�D���N�ѶV#j�E�m�6	���ⴷ{�쭌�a&��^��u�]�Ç$�����P��Hr:�c�+{e�}�]o�n�TH�����:d���:�ZbݜS'HL�9{�����k����F�m�����TOm󛌾a�J(��6�^�/���ߜ`�	_\�wC܆`��u�W�K����$vB3�q��.�z׷�[E����:����AsW�4g
�7�Cn�iX��#�c1�d�ܽ��m���)k�Hg84��գ)�����EH�V��y�Cs]8݉'N�&��J9ޥ�&�������N��Z�`S<�N��[��W�������7fH.�d9ǜZѰ9��c<�c�w����E��3�1Ԍ�U���+-�R�)�JO ���Gs��Df�&�?7=�]������#���h��e��Nb,B�?���}]���6�DT�c�f��AdGc��)6��gy����n���(ݕ���$��Zw��B�R���o0j7���$�w��y֮��	D}kt/.�
�z��f��l�!}�m���sq�cN���ot�Lz������E� #	e�c!��X���Sfl�oF\i�m9#i%�@���߭Vk��~��� u�>v������Q��S��nc漷ΐ��>��M�UeyoX��}��Z��3]����LU��c��g�TNk���(�gS1��ؽ�1�D��U�qUvn͛qÍM h�n:`�q�i��{�u�W*U�x��4����ue�`��� E��P�4�1u1��8�N缛����힓����ϊ�W�-jQf�pm��k�e���C
V�ӷǾ������߼$���*s��Ʉ�f��o!�)�q��x' �3a��H�)��<Ř��6�;+ef�iyk��(f�f�9\�#"�)���vj][�۲G!{��٭� ��SYC���[Z����@S�]zW	�m��OO,�Ce[�r�P1�]�=��c���q�%�ꥷ���B�?�6�4�SACx&�c;)ۯa���!��⹠{-n�Z�ÌZ��w�������YqJ9��B[�V�z��m證]��8A+��u�{�7����-	�#���f���֤\$�QE�x��ts��6��t:d��l��::���d�#Dn�Cs�]Cz{wo�Dv	���q���9�a��W�VKQ�ڏ`�7x���q�I�ٟ_�:8�ڀk2B��+ї9G�of���soՒnu�w}��们fʹB���:f�j�{�/������{�\�#c��h��I��M��_���ld牨��b��C�n�5[��=j�����_����K{F�I\�M��u��(�&bf0�:��8��&Ɛ��;fh�bզ��;}�yP��kd6"[0�7����ھ��~�(���,�d}�U�x�8l�dl*��^$9e�n�8�n[��ܭ0S�&�8��c�ܬ�)���R87�B�K�>q�w���L�^~�I�����iX��Ɔ�&S\�`��U�^j�^�*�
B��	�R�n�1:8���⟳�ia��L�Md�U�Ԋ�������	���7��"H�z�����N���F�QF�YM��n7q"+�s̪����u����S�Um0\ʾV:������+��[}��gK2[�4�FJ�<��*����{T�K�)�����s���i��Xe�w��#C.���Q�%Q�=7>]qڗrT� %x��W^�^�Q�dKr��-���׶!�W%Љt�@�h^���֫����s�5H@�oG [��~�.b� �M��+7����h��mƙ�)�$֚d�<�*ko��K�mN�Ik$��Ӽ3���2��T�����2�x�X��ފ�:�Lhk�T �NFw�(��ISA�1�6e?z�y���3���K�ߋйs��yr�F���&㠛�/�m�`�e�u�pf*���39q���%Њ�h�M���]MSX��SJ�ܺY�4 ٨�5Z����� +1�e���G�%4�G��*e6�X���;�<>+=^�N����P-&���2�<pgul�i�#P�+��з/Y��C%���6�{9�̒�s}MPY쨣�T��rթ"����%}��O����0���gl��]r`6Փ�4;��OB[8hFq�
vD��LV�Å��t^��I�˞����蜳U-��f*¸��#��8f��wM�<ˣ���1�@��I�қ'bU\���(�pvv�
x8o��O��|�NK��Zʫ"�\_��9#�-�����cx�G|�Ur�
^͟^�k���~�e+$.v0�h�EE.�Ov�Љ�a\�Õ�`�>a�x���;@I�
�Z�{M\P��wh��Z����aɹ��7��NJ#�ۙb(�{�^��X�`^��6#ފy������U}\�`��u���1_2�H��q"��`��(t�
�W|�Ex��ʮ��uԩ���
_(�\����t��yZ����D��ZV��x�JC&�oK�*����.�+�f�����z�������?ol
�;$��ѱ6��䔲���DT)��r���U&Q��,#�yv�wν��@(�Z��n)�j��%��iLg�׹ӗ{=�wZ�4~L�a����o�ot��C��m��E졶�nwM6�n���"�so$Y`�D�-Z���y���%��"�k���#*UK8z�\Q�*��:�NYc��]6q�6�ݽ޶y�yn�ky�(�Rn�jZڨк�F�nu4L�ȵ�,⮎��S;)j���UÁ��[�P��ٕ�hzK��H���齾�d#�ӎ�pgԝ���,�T�IZ���«(d!C�3�ȹ���&��\����L�k&wu]G�[yhB��;L�:�8a��7{F�A�r&[�eԂ��e����w+^��0�:�b��Y}8:"k�h�o�K*��b�����wZi=YQ��A�x�Lr7�G)>�
٢�r��q1Y���l�����C���dU�¢-.y���,����u*0�^��:]m�����^�^��\}�^���F���Z�ⶪ��b3q�n�&hN�4k��2lm�e�9����P|G;h��9Źm�DR�T�'˻2̀�F��u�kJh����Q|0~���K�[�=T��ފ����
�ofu��LK���o�o�@��wkMTo.f�gv;�;+p�g��6.�zoL�q�[#h��z4�e*ʞKݾ8͍w�,�$G׃�y��MF~u)�ީ4���y`�J�x��}��Eڛ�,�ɫ3MݩZ �j�Go�K���D2f���δ�l�V����[�j\À����+��NUMAXf���\�{Z~Ĵ���%��l	Y	�-�.6[\d�aq'yZ�؈��\6���M����T�c��B���Y��_d�����0>��	+ �PE���孤����$Qb��0)E�(�X,�a�b�"�$�2�0�VEY&Vd���őd*�IL�$�`�X,��
ʅHV�"�E��)�,�Ȱ�B�d�HH(�D	Y��Ȋ�E^-o��rU�Wo�?zh̥PnJ��V����§<���OWR�h��h�?��>�3�ؘunEj��q�r8��)��R?s�3vG�u�>~����>�㦾���_ke�e������ ��q;���x�{n����L<	q9r�31�b����s�Q��b�3qB��ֽ��N�i��/ٹ��+�Uaԑn'#Y{7�0;#!���zwyY��Z��_�U�����t>�<e��˗K��E�5vUYj�#5�тlZ�ť�8X�f�{
��=ي������O5��ϻ��!y+�o�=�[�	=�k^��,�ST|���^V��wSJ��G�O��i��I���U��w*���[�FR�$���I'`��^Gd�^������F��w\ky�{!r�DY��R2VV��Ty��585��V�E���C��v��k{2ȅ���z�����|�~�k�d�?�oqř��m��|Vob�yY���㘦�qBVBMf��f�zr�&�mfs�`�0YQ%�=��nf�����]��:��WLF>�����hG�ez��u	�$�J
�<X��b� ���XÁR;���קA����0d���6�x"���8����g�>��۷�oܥ�;����������5��ˡ�1��ڍ�LRI�\��9'+&E�?1k�*�{'U��1Tto��/��"C|�:j���3�q0��q8ܖ�k��mcbL�l���s&�|TnQ��p�Zɲ�y+�p���g���ؓ��<�.�x��;*�9Z�j��۾�)���	����/�r��SC�Bl܉!��:�瞄��
A�&��9.j.�aX7�/J$����"�Ynm=eYNOJ��)Q���6��%���^q�M�s������T���V,z�\��w#��%h11ur��g/�vH
��(@���ʾ���㺓Hy�%�VvVe�De�u9�c�tD���I��rq|̒~Q>��L|�49��Ӏ7�}�f�;]�c�$oK�ޙp���M��<�p�}�������ȿ_<��Z��G����F�o�{<x�p�b�L�
n�2��4�e�#R���;3��B���6e�u��Ȼ�dO/t:�R>��^���H�}�8�&'�&����}<��u�y��v��C�Ԁ��S)�!�`(z�Rm��n���I�{�O��I2�o�5�d�s�st��!4�l��I2�P�M��!�a'
 d�RM�c�E ���<������2M3㔆И�<fR��̆ܤ�C�l��4�{M�&7`q$+'�����*�ίw�Y�%͗��2�i����T�����qyX��_.�?�=�_�9����V�m���۝����(�z�]&�q�o#�y/�G�8`i���z?:��5>���$�HN�S�ChL����5�'�u	�)hz²L3I��<߹�������,�d��$�&����Lf��|�Y�@S���c�2h�	��Bz��1��s���>�yΒ��8��|r���d�ɴ��L�ϖE	���e��`����&P�@Ɯo�{�}�w�|�>=�Xu�I6��M��N>2e��I�	�C6��Pn�|�Ŧ�&��p��ﱋ�o���{�C��hi��:��!��Y=a���@�݁��	�o d&��&�["�z�;׿sw��߾�����S��L2N���C��2}�=�B���&�=@���ROS��q =Ͼ�<����{�>�Ć��+!�
I�$�I��$*d��C��O��yHu����VP�q���kzz��<�{�㤞':�B�Hq	�"�qԛ`{J�`�"�m�d>B|�6�
��	�����y�}�0� m&ن�l��u�u$�O)�
�Y1�I�-��'��݇�`͐]2������>�9���L�a�HpN��@���Y��!�L�Hq���}aP�d����e
��������Of#U��8X���R�^�Mz�]������]_�&*�L��l������!|�;��j���UԻ��K�����o� �I�?��CH�a�N2M2��P�!�z�m���$���E���1lsl�#�"���yL5Q3!�ٗI�'3x�*Vaά�Ci�XI6�Rq&�P��s�>���y���$�|a8��hCS�'Y��	�`e�d4j�>a�i8�*x�B��Xq����k�c:��pl�'���ĕ��d��i��� �d���i>a8��B��$�a����q�>��=�Z��q��!�d�=d�Ԑ�jȤ�O�N=`yi��=Hm��͆̚C��1��<��y��@�aRL!���!�l�~d�I=�$��u�RO��z�4�3�$7�u�����η���:���l�КBz��=aR�S�a:��u��p�q���	�9�!�e��ּ���o��Cl�)'sv��zì��8���1<���x�k�$��L�z�]�!�ߝ����{���z���<I+��ēhq�ILXm��1�OXu	�VC�N�����ɻԓ�$�z��;��W�>�����l�Ų,�I���d���a$��8�5���'�P��	�Iě����O��~��|��w���H\��a��ݦ�w}��6m����]�FqN��Q�DfJn:xFoF��o;���$l��"I��}�}@y{�����x�$�{@?N�M&�d���!�M[	��'�=O�*�Z@�ACi'X=5xw�}�{�I<|I<I��'�a=fY2�d=Bx͡P�z�l��O����_u�{Ϸ��&$;i/�RO�!�O�&��d�I8�!��"�Y)��`g�q��]ey��Ϸ�L�m6�V�0�e����q�b�0ӨN02}`a�Ǵ&��!�@�a;�_}���5�~����$��M�i�}�	�L8�qR�����Y'�V��8��6�q�[����..����݀x���a>dP6���'RO���CW)&��,��Lj�$��b}d�����r`��޾����P�	�Aa�'�XC�!�YN�@�CS������|�:��|�ѫ� ������s�w|�M$�;�q�6�����Cl:�2g��K���	�a�I���l��x�!6�}������<���r�e���N����d:�$�$�$�&޲N2kvE$�c�'_|���h���sߺB��v�L���x��u� |��@�<g!�P8�1)&�!�Rm�'��^�s��=q��]�}�1'X�u��/���ڂ�ٷ��\Ӊ��_�.f2(L�/�s%�;=��./�i��@�E-�W��/m>��$��l��ܒ�z=興���4�<M00�zʟ�r�
b��3;@��OXm�Щ~Y�!��x��'^�&k>���Y�{���a6���"�\Y���u�)��I1�pd2`)�l'�8�=�Xb{N�w��>�<�=��y��}� �'�d�$���$/�%B|�{I0�P��u�ԓ�6`,��'Y�����;���2\	������O[�[,��`��U��l�N~Z��r��}b����{O���p�}�-�*y����]b9p.p�ǘS.��`�:T�jE������c"[rv1� Tƣp���AXA��u��1a̋+�2��B���Ҭ���$x��vzlh�b��g��|}�HÉ�o*�O������U���$���U�5��R����7�^]�c0�WM%���U�g��m^#���!Gs�q_�G�=��x9�i~�~*}I���HuG�4|U�u{pl�J���J����1����|F��J ��$�H]dft*v�b����&K��$��P9���i�v�F�η﻾n�<��������!]�f��`�P)��������0���$�Y(&�V�֠�ld�
��r�\��~t�Y'�C�Uǂ�;�᱓����Wx��~�2R�&zE�5<�ˀj�7@uu�D��ܷs�(]4S|+xu])7��UQiH�=Ye�F}y�-~��`��u���Q�nh�7�<�M�����Tiv�_.�{�U�����娠�`D��W�z=�̶[���!{C���� cY<�����ylm����1��>�7\��v�>_�����OF��j���騦ڞJXe�%���:\P18&�w��m̛ƊP��(쇉��A7Ƥu����in u�eU�Zvfz7[U�J�V�$�`�7p��l,��`�j��$��͔v��U�=g6�¬dO]�fv^n�������;�,�r; �q:�W����ٴ,"]U��Pj���J�U���zD9��Dk͗N6�g�8�+volO�:��a�	
g`�m\DnR��M�ʥ�ɣ[��=F�Q�1m��&]r�3&��f�Wˍ�Y���5X�-R�V�v/d���-�U�W�߲*u:&<��\2��qJ��	B��w�F����~�~ǁg��*���o�����Ŷ���=�cw2fH�y1����Y2�#��[�������]�\����܃�M^Ekmf�W0a��BQ�.�WK2 )m�z��,l�)E�`�A��uC׹vo%_�7(� �Kaֹi<h�/zKT9ѧs{~�%�c0m3���Vַ��ﲍ*����#u�E��q�eQE>0S����R�|͏��Ҙꚉ	=4��>���������߻����t@!�v��d�D�=�E^�,ԕ�Wۗ.�Tѵ�6�F�
Xi�[�����}0B|gf������Zcg"&[�7�N-�U~�&ݻ�,:�N&N�z��!J�Ê�*V`4��)+�[��s���/c.M��@�m�k;��i+�d�8���
^I	O8`��csh���t�� �Ad�����G1�pFdi�ٹ�������r�Ê�0����:�[vu�s6!Fm`���V��bHj���#J�t��:�Cf�s�JȲ,!m���s˚�*��ܥ }��ܢ�{g�n
�0�ƟSU�cVt&JX6��R������tuF�!}V��"��Glj��Y�L e8�.�u�*���@�O�Yj��zH�k��ò�2��^�{:;��*���B��S��=.4��BRc������k��~z<^W�11�R�+��-�)d���b,FE�W�p����o�a���mmIX(,ͪ\bb҅lT+Օ�+e(QEFږ�(���E�b��Qb��X�!�qaJQ���iU��V�"T(�T[i���Z����Pe�h�F,U��6��Q[E�%�*ԭB�"T
�FڭKͤ�V�F�,Q�+
��%Tm�B�[J��QEU���.s�`�j�1�U��*�iZ$��R��A���S&�e��[��u�6��/6�A:��g�����h���Dz=�h�_|���*�7�����bЎ�1�h˚�C��-���ttb�b�"�n�s��ٱ1�S��A\F����9B`�])�yO}�[X�Ğ����J�c��!���9U9� �����Ce}�����M�����;�Dr�
ʫ���-З��%�G����o|rUaA�%y;��Tb�;������{�&m�c6Nu;�'|ckC[�N�r#�TQ��Q��D�*$�U_&0��Qk�f1�|!�C������*o��ϑT_�a��6�:~��sPR��V_zˑ*�q��U�|��b�Y�fO�9i��TDD{���m����xdث��*y}��Q���u�6����^��o|_�{��c�&/PC.�yJ��B���c۾��޴�M߹ӞN����}�7Z�H�8�gv�Z�z:���А�&�9�nk&�v�i@�զ�Vs�J�:ޱ���px�vEè��
gsY3.�Z��V�8�ډ�Ao����!�����&4b�V�^�"�N���bҢ�r�2���d/uB��bo:��1 G�}�+��='aWb��7S�So2���֛�}X�7�_�x�Tl��%s\�P��bC5^nN���{����6�UZU�	/�{ޏG�/m=�?L�I�;�J���Fn��a�yA���G:�1q�F�����T{�|o�u��"�
��c,�4�裸���	�r��n\x\-A�v��������Zu
vBC���2���Z�k7����E��A�v��`�@1���̃\� e�x*�v�U�����:��'!���{Y�}y�����T�w^�z����r3α���V��R�k��j���AM�Mi0�t]l�Ti O���,�qSg*��t��h���9}-�_�|8��`
�����¾68��J���WZ��ݑrQ38���z"n�ۘ���^0�9VLl� �L���W=pr�t^6�.÷#c%�q*C'��'w"�Y�� ڿv��7���jEw6�s�v�ѡt�M�	�V�*(Vۛ�d󁺦pO@����?��R�ʅy�h�����[pLu#K�cG2:SL��H3�a,��uF��y�]��&��_c0N�OQ1��ɦ4�U���
Y�Q�M�e�L茢������*�y�*u��d�_��������tlI��7~:�i�S�<�z凩~��⼸�I�˲9��m�ʊS�b�;	md,J��TZ�)�cVOrF{���Xe�c}�蛵�g�e�0fm�,�ţ�"W�����%^lO%6�Ө�!�o�b�r�,a�ci�_{
t`o��yr*	��[%�)Z��%�]�K|Mθ�D�����nF�lgD̔�IB~ݸ�Ń��aC4"�n,����s�H�<z��Xm"����W`>6Ƈ�|!r�=2$�Mtf��n����eQ�Α�cC�����r�0B7�R<�k�E;ӽ�ۣ9%������ӕ��{�*�;P�����K���x
f�
�ÿ5��ڱ��aĺ��w"Q�0��P�Ih/��z5�ˍ����7�ڃ�]r�	R]��?<J�=y����F�3t�l5 ]���a�֗W}������A��`4��
'#�;��N��ͱ��<�Cɘ�Y��xz���-q���N*����:M���V��AȖ����4tB�A��t��:�E�x��]>Z����s��l�,��{q%g������:���x�C�bj.�dZu^jfD�*{&�{���ӯ����l٪́}5z2��v�Wz��Bx���>l���&�r��XV%GK�ysה�m����`��,�s/�1T��9�&_$��Dz#o���}WdC�{���%f)�]LkqX��,\
T�M�
������/������<���k,�>U����*�64�o��/mUJ�BBo:��7�;+g#2�Xh��v[0�5m���ZT�l�wh���i�p"QRm��΄�2xi-�Zũ���D�U�W�p�$��)*Ӊȭ��_�m��yOb�<�(������N�$:���lq'�E�wta,��0�39݉iY��V��uXy�b�Cg
�)�[/�G���&���$�d�9���)r�tw��8}b��]����g�7���8�L��9��s������ji�w�s�7�iv�����Fn������W-��7�����qowf!�2v׳�x^��o��ߺ��b���\rG}���)�ɮ;���)ȼp!J5cu*��IY�x�-k��u�<&��%��(�v�8��!a������e>K�먝&���%�k�l��9���ē-�dr��d�-k���.�s��ooq�!ȩ��Z�,ؘ����A'HX~���8w�Nі�)���$��ҷ��ˍG'�y�a+0*h�n��nw������{�,��4e��0�q�pޜ�;XYd�Y!�&r���r~W�}��h-�?i�[�][Iâa��z�l�<�����fkj%+�0bn0�	������\�wC�M��x�[W��OԿ}�>X}��R�݃o:��;Ւ�u2��j����|��>�صA6�OՏàʣ�e���p\%׽�����Y��dY㴗s����|�Y2e���ְ��U���0��6�(K5��zvN�l"Ի���N�g,��yw*�XV:;
��1c�2�m^���f���ӈ�ȡ7#CQ�uʻ�q���ѣ��M[��-����T̩�#xe��w*���	/�ޏz�M�k�m;���������q���o["������%:$��R���#$P��.�Y���cR,�&�~����λ�Gz�]�
ޟ��Tg��KSZ���av��9����M�3�]�m��Q�K`���5��:���y��O�\�k���1��ܮ���܏AM��ǖ��o��rm���ə�j^T�ڊƵ���fOE���"��H�G<���}�f}�*�+��2�n�O���^U��Z	�5���^�r����__k��F	�7�0�����q�����C.��7��#�kV9V	���z��4��Ku��hH9��}p���|�$1��&�&~���Xs��5�|^?<�_��>ŷws�%��y���'�L�/&���:�)P��/{��m
���<��d�koK膂�{@��M�҉֐�F��;�k��@L�2i�p�@6��3�LZf�\%�|q#��n<âF���:�z���p�a��D�Üۖ�Q� �W*cnSۚ�L��V���=�{c\�_��L<yf�n����lǜͲ���{I�&:�lb8�WF�+2�v2�[�up�I�o�>��_,�8Z}��M�-v%
�h��5ɚ�}�����x�.WwNM橡d��FU�̣�+�vtU٫�&wS5�f`��	��v���%�a�aP�W���1&^�b�̧(f�C���M��7���ݛj=~���Ϲf��/\���s��\�m��ݔ&s=s�?�NSɹ�OP&�Mz�t�Ov�#�ν���[ɻ�J m�+{�fM/ul7�57��:=�&�#4@�Y�J��|ߢF1���A����P�����2V�N��;z�`W`ƖA%�;{Ecl�yX��P��G��Pd��ꢾ�G7��ܞ�5��-S��F�Ww6�u�v��E���ܓ�i�Ĺ�$��|�٥ ]��
ԑ,��c�y�TH��t5tC��{v
@���vi:�v�b��֔�������QX�F�*z�Y1j�Y�ƨ��,0¤b#"��a8e�U���*�b� �b�UAEAVr�b���UX�PTT�e��U�=�닿�s�����IK������:RA���"�����"#�e�eI?�SZ�GU]�J�GԲ�0������M�r�U�b�ڃ�1��L�9��攝Q�9$<Y�O"9�{H���؉�P �i���v��O@�Z��l0̐���U��酸wl�����w�QعAF��Q�W,�[V`#�ֲ4���vS�������E�Q��T+D5��{l׻M����m\bR�����5����f�V�j(�Y������`��P\��u���8��[)�g�5��g�:~N������DYh�<�:���Ԩ=�~���Q�<.�����`�3L�t�'EÊ_{��Gg�<��!wE�cL��aT�7�>��$�M�j����1���".�F�<Qvׄ�Z��*���֎n u�U-N�tY�j��]^�n�\�o8B&�S.�3^�:��t�$��������Z[�\�8ü�]��K aU��\�H�ȱƫ5���E%�T6�CP/��_$���9�<z��,;Sy�*�+qV��]��Dn&4�w_[81��#$l�Sl��^��dя�:�]2�Wf�繃d�BGp��
�uM�v7M.�zk
��^Ls�����C�i������x�aM�Ο�����tRUz�]��D���L�Fx�r(к)5�P�=��h6u��bo�d���E�ͮ���\�'���۸�$�����э$A;���Q�h�jD�c;Zh��f��հ�C���mANf�;�>��^��u*c}��S}~��D��룺���q	g�+�?%M�f���ީ˝�o�MY� ��y����h�/�W�!,��G<���J^�$<e������ʱ)I��U�/k"ZP�5'GfS|*Έ��f��F�fv�c�R�R=�j���U( �G���;ͷGU��)_��M�us|zz(�������C$��7"����'��2�%���*��ҽ�2�c�*5Ќ|f5�o.�R"��/��_d�/n����+�MlU���#wu|�A� �xȚ��g-��w�l<�Q�5��Ӹ��p��"uT���;�g�����c:�Ēbp����Y;Y�XD�#j�-	y���C�0�8w9n����z�,��-��k8�}�{�L��dܝ�������v�v�������/�<w�3κN��D���Z���j)q�]ݛ�Ē�
�*C��Dz ���O�)>7��f![�Z<�][��K��5:�NE{"Pw�5V*l@wۺx�F���aW���r4ʍ�n/����W׎*N7у��S�Ӻ�7�'o�٪O��j�,F���oK:+c��t����c��U�b�g������Y���Έ�ʝ9o����kH�)qp]��b�X�f���ᳫ�50�{���ad��J�A�g�'�6��M3��n�f!���&��M�;'��_"�ڴ&Y�F�z=��^��,�A���.yv�j�q}��T�X^f^+�rrlb5�$8�	�\�h�[�Wވ���\�[����f(�^�MTiۇ��63-JCq��s �݂ge.Mp�ްt5{gt�5�	�� �j� �;����u�g���O_�﮲�b�^�Zd������X7"�{����:�~�i+���EeE^���li�s����k��ꝁ����7��pS�A�]�n�f+�}����Z��������`��ä2]�d��ѧJO�%�1q�6+�e�7���u^��Hi�C��+;�JUˌ%��m^�P��f���{���A+�ٴ�mM-h�������{'aO�.h�!p�W��DE�%4�>�*+�Q�i���\w�W� |҉��8�f�RI!
j�Lì���{���bk��#�	���v�-��CV����n�ȳQz"�Y�&�u�|��m��U'�]t?rj�{��OX~�qI�������$�9��C9#�����z�������!�vzƎ�~G�N�����G4��y�N)��~\T�&�Y�F,,Z%Fϋ�������׾Y�9�>�:��,��\�wV�#�-�g\����LC�7XXfR��y���g8*S��7��Iؼ�����"oS���zrY�y#�a�*��wXECu��F+��{5�ZMը��]"��Fj6I���=#�m��3?C۩���&�91�!GƼ��m����W����D�=�����{R�=�XM8�����{d��=���8\x���O�~����A�xC?1��u����4�k�y
��O��r6m,>�}�[��ο��SL���
�K�O�h"�9�ԝb����:D�t�i0��i����=ʅ![��7�:s}��(�XE/:*s��y�6v�&�͊P��ޗל��R�`�z�C��A�m����ف ieL|Y~��LcNgO�GA�/&Ϟ"r��#�ڽ�{��/��(�v�W�E�dx�ш��A��+bD����7�Q5��'WIŚ�3wՍ~5����\�8��/Nm)x"6����ܧ�E��䮁͌($.J��WжQ�8��{�c�晇�u@�i��\��a���0��DQ&�N���f{shX#�$�-cN0��xtE��j��W�_�}�~>�h��0�O��L6���6vzt�<�M��	a{�a�B�$����ځ6,��t0�����co)0.�º�N��b�L�9�oi�_�N�0��#�2��&&���=1�#Ђ�����Oz,1λ�^U�?t@����A�_CI?h�����{�{�r���0�U�s�@�] �g���%���{<�8/������ �����r	����ot���z,>�@��6xX��C��Ls�{}]z뼳D��2ċ�쐣J��Y�n��2�͜�4��y�ĵS0K�:�W�L�+V��f��O ���;!����I)?>{���~�a�W �Ԭ�>�[_���*����E6c\��U6�;�"��� �򠭂�@r+ܭ��vfw��'�Ggھ�C��񣸾���9��vP�k��~�#�L0x���JCK�N&\��1^�[*3�/;�}�.C���
��t��m�^yU�շB�����i&g��6Iػ����T�K�~������sdC9{PIKRp�D��qr��ê<�[3}�XeD��SCڑ�� #<�THk�����k}�R�&/"�4p�"��h�ǈd����}��CI����_S���ֆ�k�5>�D�bV��x�_�=������J��8��;��&i?k�}e�~�t��VCU�y�����1�4a��x������w���@Q�"R����3l�(E�\�.9֎Ue��]��(��h�Q�L��`����#�X\e'{bȹu��V���"h<��U��-V/�Dj��V���Y{�k;-��ebt"+L�����{�������W(4=��=4.��-Ƚ}h��{�≝}�Կp{��Q�r�]�o��/_o�Ԣ9t��&�S��Q��o�=;���X8���x�;P��;a�F�����_b�b�Α�J�.̣r�ZG%-ޘ����w�(��(�7(��W}�r�f��zXy)EV�O�C�	*¸��_#�q�5�1hNw@c�^-�㫽�F|K�����6�%���ύɮ���W���dZW����{��u��~m�>;�i��L�e���0�V��Zx�t�V�f�S���yMu��=Ψh��Z�qn"Y�f �M��v�؊�i�mt�%�36��ê�Y�z����-*bgm�EWIK�Uv��沫��ag�4)���.��2�|ZǸi����S�\��|na3�0p�o���d��^��C,y�R��CL&�� �:';.m�{ǯ�	�RjIp�� ��!nT���~�[�+�e���Y�Z5|r��7Z��T�QU���e\Ys��ݸ[��e\|���6Нd#r��[!]њs0�!m�RF�rԊmap���tWun����B��gpW�4^_�*�U�Lg�7t=�9�r~H�"�Vv����]Ҭ������-�V��
�ʪ
��R�(Ԩ*�A�h�B��1�����"��0QuK��%�լF��p�D�z6� ������{�	���FJ��f�^GWr�tF����f¤�k�;�g��Q��6C�W�k�*��v��yP�4�j(�����h��_y0����1�����K�P4��v��r�|Q�^ �[�qă�藍�D�#p��`�f�wg��#�#���l��)_i�
���*�m���،��9��<�ٯTԛ=�04ۙ��2�����0�`KU��f�<Gp_\]�cW>�������˃QW�
L����Tj��������/�~27�~�>dU1�p�ܴ�Ś8<@����N���f�Z�WHi�kh#��?`j�I����=��V8�!�LR�e�HC���䎝�O��"/�=����zP�֍OjM;�W��}�N��������N܂!�}i�u�������6�{ԅ��Wwr$-�(��� �1�o1x���q�v�e}Oڦ���ݽ{�U�=����iT�C��22.���va���[~3u�~��k���-���ei~��|�hj���?m]���u��}�`b*.�<��Ϗ�6����U7��ER����"Θ���<*]FK��JԷs�ɇ�a�<~�_@w�;���q�|}�^�.���4�l�S�r�ļb�e�1���]���q��Wʞ������ּQ����O���i�F�>�K��{_�:٦�2�T?V�~�O�k�f�~�U��w��)��䆛:hF�#"|F\��v�箴��iWf��F@)���	�;OڥMP5[�E`�Ỗ�O�y��v�"��.���Q�m��I�WOV���c6HE}�ᬶU��?|�$�!�⢹x�1��Y�(WwW���C�|Y@G����$:����8��6����?�c9W�/{�P兜+W�EY�B)!y���Ur~�]�
�\+�T�7��+��(P�9t}���+��y�Nl�u�"�A�b��)3�SWN�L���ۚ�d�AkV4G���~шV�>�23
l�wSb�����GL&�z�6ok�����s[�!�z�#r��Ը�t�T�%z�F��	A��4���������H�b�4���*�t�ؓK�D�sn�=��)Q�x�D?�q�1�#� "����v��~��`�j1��������$}PWY�u#�\�9�joۥ^��}Ԉ'b��$�Q�Ij�b���G���������:#I?
k���U�gr7o��E������<�s�@�1�M�/�{�%uf��y>"���r��Pz�`ed��7T<������Ը�㚼kQ(�&��xX��C��B���]��I����LYw7=1q�+0j���@ώ�\�o=r�<��Z�6X�����R^�F�<���+�ǼQ�dt������^�K�b��������<��0�$!m��F���)mٕ���1^�����\N�yy>\�z���u�ŀ��#G����s�*���ޠ<GbI�l�$^ke�b�����՛�����k�t��^,}^P��Ѯ���'c�l�Dq�V�1J�:��$��J���Ci�V��w`�.f$VpI⾈�l�X�B�0�*��HQԇ6Vw�S\G��>��Ҷ���7ß��~_.Ck[,�HYc��6_�}u���Ii��,Ze	KN�l��Ȱ�!�V�X߰�?_�uC�=�P�i9����`�<z�x�����wnf2~h�Q���Rˈ��X����/�Ӟ����1D�>�"G2[����d�K������%��{C4p��u}��nc�!E�K�Ϣgj�3_q��;w�xk��x���+�1[$.K���;��﷓G҃/��w�>�̙�DԐo۱P,ۖ)�� ݦ������S"�[0��<x���<����h7sS�^3�}���\��
�p��R�#6��!�SN���2��nv�٦�@󑃧	Js�m�qr(�����y/Ȋ��ͦ'ceO�Tff�/�1�r��AW>��C�0�G5ѫz�V���0��O��0�2���xЊ�)qg�:QK&c���]��{�)k�D�4<:Ц�����3eS��7|w2��"�O�R촉sU$1�����u�o�{�"��^8o�`q�t�d�0��p�{{����>_>{��1�o��b��]��p��rv�����>��<�C�5����+H��z����9	��y��oKu�f��TL��������(r�N��$̻���Dg/8�V�֐��xϐt�h�[CHJ��}�}���"F�ł/�j��{P��C���Х쁷�o�\#qC�/bT)�ͤf� B!M�t��x��Sz�v$���2�:���#�I�}&������H��&��ˊN~}��7��
Ɗz¥����ƢxƯ��OŤg9!FL�^�v/�'�ZҎW���i|0�g \���sf�o��4f����ؙq	��h�5��ӟ_.�W��#��k�(��v���|������\Aڝ��/�}L�(E�漗�qB��5�g��b��F����{�Ƈ�l��������׆b�K�_�}����~9N6~�xApp9O��v`!�B�$g�u��7<�ꌝ���"ύL{ʾ#H�A9�o����V��Qm��w\��c�i�M��=��[~���D���@�:I��OK�Pȳ#* �fb��tg��7;\%ye��U�����ѳ�S&�*Ly�����ߗ��j�Z��o���!�{+L��A\v�7�B�K�>(���_o6ʎ����J��mT��)����.�m�V��5؉�r��_je���aR$��ƒ���}�����Y�^h!���l��H�&����Z|��M��yY�͙��xj8�Fi��N�E�@GF���RԼ������nO?\@��:�5�E{�c)v$3��.S�����C�u��dLN+�244�@�(̙Sa���^3W���6cd1#څWE�+�W�ۢ��8�C���D��D���I��x��sg���JA��E��#�Ĭ�C��eC�>%zyq<W�ED��Ms����S�.R�_�%YR�L5g�~�zsT#�~��b_��B���_�՞�Y������}��}j*BL�էY�yH�P�&`�05)����)f���觚���@�@����go�_!Ƈ�<Օpo�-Jɒ�`�T���aߔ�HT6�M��I�90��qY�ͦO��7.��,/1��lG��4�n�{���I����Ƚ�c�'!D��U�1!�U31��Vx=rս��ݸ�V�/�%�RA
Z�c���}��G�;x��*{����]������x�E:���Aj�G���s����b�}4�8�eF# �����M�y����K@��H�^�a�iM_P���<�\x�<B)�����7~��J �Z�ގ�
S�Ȉډum�\�<a@�Ĝ��*%e�AR$ag�V�'���C�ɽ7�Z4��BMt��/ͻD��1D{:�S�yx#�@V��5G�Jt6K&o�Wv$�7�'3���\���*�\{�_���M6�O�u��:e׻���<ZA��K�ϓ{&G�ٛY�6E���ψ�\(��h��R���yu�)5������Tt�����>�q��5�
;z����G�o H����s��!��H��dO(E��f�<x�?3��je��^f�Y%Ğ":c W,�)RTgΙj�Ѝ�N�+.+jdٽ���<�����g����Ä���Y��uT��-K_J$0�8���kI7�u�=�����ԡ�����i�f;$��ƁH���#�a>k�X�N���^��`qߎ�@�,�Uֹ�
�o���L<7��V�J�}/���RM	�^���ӭ������ɭ�1�rd|ntV�S��o-F�Jp-�q�J��3�n���*�qҾ�s�[��X�����v6�+���>9[�?9|s�y�qE���Y���"��I���@mY8�h�32+�EyJ�%z�X\��hê��vRpY�0G�c'��2tR��LoA}��[Q�w��i�zK���া�VE�m�/�=���Ժ�V�WG��監[@]b�sM��5������v��5�Y]ϩL���6Z3��$1�L]��*��&m�Թ1����E������*�ޣR]��X
J5��5�QN�m�҆h�+���D����T�z��T�\�h¨��E�#��֖|!@cG�y7�i�)O%d�E���&R��'Wk�K�6�~�<T�p��\�2���1fY����X�\+�^�]ueVl�s��$ƞ��6���_H���^����=7����ʃ2��u.ӑŧH�]ކ>0f޵G^���BQB�k1u�{sie�B�z��_u�~��^~��u䝰k���BgO�v�Ko�Zm�y8����a����MZ�4�5D�� ^�vؘ�R�~sE����r�t�r�OU���K�/�N�%�;��:�V��зC7EI���0r�5=�ƀ�C��}|�nf-��mn�4���}�˰����%���bS�L�
t
Zc�
J���yW�w�7��D%&i�Q���,�V
�x-�{;T�T�͋��Dd1�\��8��8��`͑�v�֩v4�X���P�g�r�g�nK�*t��@�R�h)��8�\7���j�-k�`0��F�r�R�X1�u��
��V��h��(�-qJ�ҴkE�[F�a�st�f��j-���T��YPKJ#[�W�9j�j0�1J-h��SR���1CD �Q)�#�.���ý~*T�f�Vv�ؠhI��<�=�n���i�ց���u�<m�B/�c�������Z��C���h�����!h��������EE�X|`����}��v�\�)1��c�8.��t ��8� �b�J=��{�O�q|��x?�h�7��ԵV}�eoZ�_��6�gU�F4V!)i�9qz��P��dl[��Е��;��b�^�QB����ƀ������,5Y>��+���	i�_)��,��A��V��ZN��\˿{��!D뷼�j֘��Ɏʅ=�5��^�aQFa
R��c}��G����S�3�k�x����z����&;��5~�D�V�6��n�p��<�����]g�VMyGv��#Q��r���� 	ձN1NpF\Ho�)�y0�'��5�>��U�=x��0�P+z��E%��He���>��\ٓ�kW}��;��7e�ӏ�����Y�����2X�~2��!�.\�u�[0f��f��0$$�.=�!�#Kh[�1ˏ�����^�5w�sv��{ۛ~,���MB�2�$���î�L<�3�KB�5�^ɋt�&
���G��A���cC��$(�|��g�9a�,��e�P�D��o�	�	P�m������Ә��w$E�#ڂ��YBΟ8���ۛ��+��G��C�q�Q<��!��4!��d���w�P����Uz��O�bQy�&l�ŌC\q��/t����G��|�cDCC�'������X�U�{�sr�Z�:*{�O����>����?|g��^mܾ�9��A:T�K͎�Dtf�]bGŴ٣r��v-�$=ʭ*@rK�Q�m�3��g���GM��6V��/!���/�w��݈{q��y}Ʒ���6(����S�i��;k�޾��e!��Go���]�"E�5G��]��؅
�T�Fva��1������N�].�nu�U�r��E���AV��	j�g���8ϼ����귺g�s~��'$bC�?k����R}�>85x��JJMV�{�,���TXQ�� �Щٔt*��wC!�}ڃ�q����@7��"m�gI#+�- Y�7;�o5��*c�ikVH�Z���m���\Zߚ�yt��T�.� ����daC��{�uM������yf�:f������ef�9��R��w#4F(�goe)Di�q卆c=;b �9JK�?d���[�?�e[e��/�!O���R�š�x�e�FE�TH��]N��p�h$��}�Bv���{n%\9R� #�_hϲv}�3���G_D%!z�a��A�j]��J�y�Y��;�GS�����(�0��/�-�l*s�o[W��zK'�zb\+8t�'Vq^��c�H8��m�%ٻ/Jl��;y;0��쩅-D�J��@�Y�ސZ����Kv~WU�VOKq��U{�L���/fźc;�����?�B�ޑq�&�E�"�}ZǏޫ���#���_w�,o!�Ia%�
��ʘ�U�h뀖����̭�~��nyц��za�QY�w{Eت�,{=%�1G�p�x(��AJ1
�ݪ��j��)8&!�SVmȁ�1��!ݙ�+!-��ă}YxivjKJE}%6�LG|�}9�BZ��?Q�>5�Ǉj0��W�}դ��Mi��E��i�V;$�4�Ю+�)���i>���:!mx��I?P����x�����D$��B�Ɵ�i�Ϸ"�g���7o�P}�����*/ȔE���<F\���;���ů�3������Ƽ,Z�j
�%�Y��a�j��yv�e�gw�O��J8GyiI�H�:B��8��;]�������/W�����#N4E�����l��n�������sӮ�ߍL���^�v�B`�N0K�� ��C���`��oJ.��夵�nj)b��x����I�U��^^�
e,�;�In��Uk-v�w�^��o�ؔ�����>��o�a��o]57���R������6�&~ϧ�2	�R��9���M5�����l�3ٸ�{�=���>:B�N={�H�"�*#�B��v�fĭ�mtt���<�&���.#Ƃ�EO0��l��ٻ�����S�(���������'(����}�Y�TG�a.?��*��X�,,�L}�`ٯ��c�G�Yl
�>]���7�xݬ��Z[UP��W�݄BH��p�-�s��\}�s��C��̆�M�x�ʎ�C��P�P�p$BX�DK�*k��C�����K�h�AU��1Yw�#M�F��*�p�����a�㼇�g.5?n�_R$��|`�z
�>y�#��<3�����s)Q�������p&s��@��o��vތ6v����jkV��*�Klΐ�+��.��I}�!ͽ��1���!�Z�ml�:EjWʬ�����_�/7\:�L4t��\CH�T
d1�f1�B��ޣ���3��P��(T��f#j�}�9�qܞf��u����#�|Tf�ƅ��+�������+�g�'�������8~�4�5��r����Qz�^�\#���P�:��J�8jf �L��}*��DA���4��s�ǟ1�����.���%fS����u���ذ� �EFÕ~�hR���#ON��u�vw��F�>�*Z�������/�^��N�������H�,�v���o��}�>-8g�:���k��8�Y�[�&]v���-c���f���6s�8�v���:�YvDf��,M{��Ƿd�57�WށZ�m����;��:ٸ���u
n���Ÿ�F���b�_����Y�q����X�M�U�0$3����[�vv�P$s����Ya� +��^�h�ᕵ��x=7�a��1!贍���7@��@Q�]ۛ�=
���+�t��q�ƈ���:h�e�3O1�8����8G ���l餆Z��bI��Ǘ���!5�0�{�r�7c8E�x/�"Q;��!z�a˼3��|�y���la>U�x���A}H���~������U�T��o"=z���<E}H[�Ҳ����+6׶�=Qύ�}�ᔇ�i�k�y�����"�������Z���}|�pV�ZX��V���I��g�P�m�Zޗ�H�x�;�`�}��Op�cI�*
�Y��A$.��ѼD����x{��=�z}�����D���S�����L� ��\�S|��q~�ÝO���\2dl0D���6a�V��5������/���~,1�8I�(:c����z�ܭ�`�[�m?w��Q&�g�c���\B�%t���nx�p��W0�BZ����+�X��~���V�&�y�~����p���>��0�!<z~��e�O���ﯼ��"bGO�0�x���Mx��0�#I�M��g�;޼� �i&D�-[���=k��<v��y�L�xJ9�/�-.�(F�#������u�=!Zm_m�w�9���.:D�<�dYמ08����wz|%�jM�Uħ;NF	BO���6�Xţ'4w2b�zMխ=�-��9�L�}���gEG�L�jT��֔v.�gt��ČeN�E%���ͷ���P�]��W=0UxxԔ*�"ΐ�W7��r�;8a��3�1K�Ŧ�Ilb�����/j�+Fx��W�����C|5�TB�<h�5�Kg�ʐje\MA�c�JV�g���E�a �"�_q\��ִ�s�-'����mg��x�(vA�-/�:�ӅC�۩��_eW��d�G�4�L	��EQ��"L�e�\:َƐtN�k�!���,��(E�A5�q'*����H#B�^j�~�xE��~�C+�ȫZ`!ņ�E�-�������P�ǤAK�b?���ݬo�XYµ}nU6}�7�{/�t,P���b˿!,�ǘ�׋�uxX���D��k7(�kF�\l]m�N�^�XY��˃�ݺ��˅õ,��A�2�����m��t�+��;�����}]:��#�%:�J��&Z�}g���p,EY.��Y���P�4F�9��y���Y�x����۸�t��t�`���X_�*�4��&Ă��6�qj�Sї����j<ԀB�;΅�� �(��P��[h�Nee������b̺҂�-��d���n�E��Y۸��k�ǚ�cYܣ�0�=�յj6�N���W�^(ӫ�++$�wR�t�w��JQ�sM�S6&[놅�
�_����0�jŮ���員�GN��Őx��ـ�f�w��=M��,*�Ɠ�;/�kp���V��}6��9��Wqm��r��뙸����Hy�oAY]|�����f������A�cAm��AD���s��-��g+Vf��w��Y�O`�Q�NO��T��1��"�Ζﱉ1x���7/���>x���SF�����[�g���Ue%W����'vsY�L��O-�՗J�T�]twX����i�������i�n/z��V�To�u�էZVV��:o5G�:i	�%Iȃ�o��~:��Q�9..a��QV�Ot<�ӛ6':w8Ƭ�QJ燼�/CV��ә�U�i~�D��X�Pfݞ\�-:&��.nV�$�]�ȋQ���"\����u& �s����U�OnT����f�j!n���5���U o%�5+P&����d��1�Ɩ��P�VG	(�f���1��VQj-PY�
#3�k!S��b4�T����WĢ���-�Y��ACX�Rڠ�e�)Z�%h�ch�b�X��J�ܫ�*\cYn�1��"�K��˅2�p���L�&�)���Z��ELk&�_J@�	/�_|�U���hf�6�%,��b��.��V��7�tp�X8y��-����B�����3�0�����yq�U�!��/�.�y�~��븻��EB�6�E��!,��u���p���p������uF�������ih/�FZ�۽�z^��~HiR�����9qej�"ILZ�Q���T�q�5u`IuS�	m��iP���4�՛��~�-�>��1��q0����Ӹ���9�Rܫ�AG��}���侶�ç�y�
�'NnbA���r�EÙ�Bʜ���/V�+��@�c��$�ܧ����:�`
�A�Hsa�\B��j�s�5��ژ鹎5��X�2%7���~؉��y:����Mw�Õ�$��vq���R"U���ͩ�����-�'p� ��LW�%���r�]��w��#�rvι-%�� �(�ꤚ�{�ۏ�E�11ʆ�ke�fd�/<�W����� ~ɬF��o�CX��=w=!z+��ܱ�� ̤ya Utj�\vvs��)�}-J��?`Ӧ�}�y���E�7�*�*ͨRj����k+C�z�h����KH�yc���<.�Qy���G��)A���V�PDZ¤M�n��Kh/yڅ��nT���QG�R��(B�0+����l|��r�8ćE�o/��5��Oc�ڝ��ȇ0�T9b���uJv\����Kw�o/I�+|��7.���@��$e+��È�Mx�]��~����U���vC�����ܽB���6昌u^ Н�*�=�xt���0f`~��ʎ���cS��%�����N��Z��.<W�ވ�=x[h�t�sI���J���� �1s_�����o��:�ԇ�XF�J�"F=-�~Ǵ&{��אa�=9��Ha��^+c*�Ya��+�������l}(	rֆac��k��\(1\��S�Y��G�O(����
��({���N��ܨ�ʪ�"�J�n���O��^$���!����|مO];�V�7w����^# _x�ߊ��K	,r	�`�Ɩ�������B;���v1��-��n�rf`�yY��u\6��&Q���)q૜x�j����x�~듵[���l�=�gę��h�w��Y<z`"�Y�j��'%�9wS�q�d˒-ʛ�z�?{ޚ��э�X����孒��]ewKaI��;��⪴��8���xi���i����S������.D��!K&���=�;���'�"x����������=��W�?U����h�z�~�ܰ�'�7d!��;pb�1b�0���.Vf6|�U0�ɞ�QB�e�xI�s��}�d�����|)q��]����Cy}5V�t�g�&N�����w��*������4�Z~��	��g��=�1sXA��x�H��-8`�㤞j�(+�)ru�����X���w��^�5n�|�����j���'�GXE\���3�Y%�ӟ�:��@be����s�T��}�e�i�>qC�ǯy@�񳦣b��zɰW{g��|p�ԣ��Ma��c>󽠧�����c�֧��U
L�O5�VGH��盙�Y�y{ҷ��q{[�ŧӴ����<u����1����!k�r�CHGR���8���g��̾�Y�C4}e_�`�������5�U]�Z$OzX���)i1}<�:}��yag��;뽾��Ϫʇ��������;#��x�>6z��J�{��/��>A8D�D\�lx���^�齻�냆*���MD$�#A�$CM�ezx��<
�1S�K���\��ҳxV�r�p�kx��]{���V��&hR��g.,����(�K�Φ=��^{]Q$L@��Ɩx�Er�y�iEU��H�|�����d��X�J�φPbk#�����Ջ�(J�쵎ɕ�b�-S��:9���O_t�������1޾�b����ʑ���Yح;0����]2�7�B�K�6T��������6F���C���7��a�� �>���6i�%<l[_�hA��߼r�G2
guƅk~c���2gw��ځ6A�~>#IAa���4��t���>oPτ�~����ꞜcF<�,����"G��u�?lB�}��_{��ե`��0����S���10Uz�r�h����N�ow$��~�OK(��.4FZE�m�S���C�����N��ʛ�4ϖ�Z_>5����<>��㻑ۼ��{цx^�����XC<��Fچ�Ɔ��w���މ�����~��z��d�FrN�=b1��ǫ;s��f����0�w�}��o
�"-tI&�Vt��{A���v_����ӑ�}�a}3��w��>Ƿ@�|��"D
W�ٗF�,sٚz�T�ך�ɽ0�ؐ�In����F=ԙ}�cf�`^�����)�!1o)�)hv����֕%�Aô5��8�C�O�z��Zb<��r��o�|ﯳ�9,�C^�%�
^.�ۉ�Ǐ��j���г�4<՟"^44k|P��'Z��r�oH��|~~����.`��30'�"K˹�ʎ�s��5�3)Q�w�v�r>]5�$ᚂ�Y�=���U���B�c�V9$��E�:EZ8�Ha��p����w����|F8��ƇS���-+m�k�q�{W�7��wwh>�E�x�V���妊9���;��*�Y��I ���7.����C5o�"��4�rۦ2��xs�#���M�(�󫒞_G�m��	��A=�w$Ñ	~5�-�vpy�ϖ�*���Y�<�䘞ι�?,Oݗ�_����ޏDG�5c�m�H�ڏ�:��e�ǋ�>:�K��la��*��E�+*b �U]�Z�ß=�r&g�2�rr��c.�.\��[/iI�ͧ7�#���K����p>���펾��3����qY��z�Y	��T�������z�$���E�tm�+�P��=,E�gd���r������D9���#KKI"���A��G����r��8�/=~����{����70'�&*���1�u���7,�Z���?��X�V�a�:hj
�%s��1�V�9��ǘ��Fv\󮺁
��L��� ���DQ^~�g��]�x_�i�#HC��q�[Ip��/}w+��g���M��$��&y�iTt� ������9l�6��mJ���ا�7{/;�n�:��3k�6^kO(�P�oq_G�މ�m���.���n.k(��)�U4�66��1*d�(#�q��k�?T��	Pt�!�r~P�֔}���<7׷����%�!�
��Y�N�����N�Yj<��W;}�2�����Gx��N��D�8{�9�go-��j�6S_!�`�ǹU ��Υ��x�lYު��n�*�G�xk��>��`�þa�V��΅=/�	/{+{;��{觔X�b�1����\��o���,5c�=�ۺ�!�_B$��:qQ51�;�x�%Nʗ�&o����~T#�����F�ι�t���R Yͧ�`
���nR6QI�a�P��"=�{7Q�6sw�����;����L9|��r���x͐f"�,�2�m�6e.�b������v���h�,�K霧<ؒ�BrE$j����+8㼿��m!@6:�\�����9��fT9���UEKM�r�Q3��xE_7�(�r���I���2�'}�g��DJ�7�.�]��]�7���ϖ�L�J�f��C�i15�D8�)�}������l�>�x`�k-zT�!L5��"�m���V������<�G?b�}�S�+�-�Yz�	,�)^�1�6j']��I��K�i�-�2��P��$�m��מ�օj�a�W!�)Ș��I5����{{���&+>��C�`�G���Z���e�Ù�J��^ߺ�V�#���e9���xْ���8���_I�hE�M^d\wX�Uu*�:^����ٿ�7�7�%]Ly��j�s��Զ�<Fɟd#�[�0�%�v�,t��O�p���3>�J&I�eY"��opP��«��-
�K�M���L�bh��{��01!�8.z虯�{�3|��g)~6�1 ���̔�mA��h"è�c���{�A�!L�}������h������=�[��{	OJxAA����?w�M��5�Kp8�>�@��H�ｴ��4Jo��wh��g2��L����oF�Rh������R����4�v�Pf�9�[7��Oe��P���02̙�
!e��
s��Dv1H�g���*]�%���6n mcG/��Q�ӆu���;��pZꪃ��-+{F�͓\4�:W552S�\N_�ĺ�I ���%B�7�\���l�Y�4L�9zq=��:�"�{>��j;�)�)�V���.?�T�QbeǙ����6#�X��;x�ogʶ���؂��N�Wfn����l��0��c�)%_Yg� Nw���;��N��œ^�"cM3��O/	�b�����|cq�[#���<����9���ǺZ^�.�ڳ����|���.�P=�(�fQ��V�+��1/��l_eh�
Q��'i����t��]I�:8G�ôәd;�W.,,�Ђ�d8znMnR�!STbXu����yң�L�n�gJ��3t�3D�e��-v>M'�<Ǐ��6������y.Q9�L�'QM�X�[Ƅ�m�F�G:���5Kk��������*�9e�=�~:H�-���A\X&����%�(��	1�cƮ1**��Q0�f�dh�L���KlU0�X���-��r13J�b�-�ue`�+��mid�Fa+�+�R�hn-\1p��Ų��j�Uk+m�b��3�ήQL�DQ�╘cB��Z[h-j���ᨪ����m��QDŨ���Ì2�F�L!H&��,�+iX֪��*��V�0U�E#(�T�8�-&0T@m��1�1��f�2�A`+�qJ�,ūD0�AH�Q����X��QQ���`IP��eh����"a�E�kjV,�����VjTLZ�ł�&-M8�E�E�4���e��+��Dsi����V�b�8L.R�,�0g8��l[j"�D �A>��`��7"u~��Z�]u��^�iԫ����n9J�c��꯻��{o� �s�
��� i B��:���m��s�{N0H;����� �R�XC:���k��e>8���J�_���x�M9��b����T��8�Z����y)W����c�X#M]���MW�V�k��&�GS�XH�xO�uQ��V��#M����vR!�N�뜞e���
�8	wf��
���3�q���R�`���!����Y~�{��^"����U�!�k��K���+H��U�36���:YDd\x�B� x�$m,�!4����������ɻ��)��ڧ����M�Q�1�%��屜*�2�� V�pMw
n���l���������ߺOQ��voG
�>c��C��>��<g�!fi��F�W!Y��s�.�ԪMm'F�ҝ�g9 �rpd本ST_m��^$�%�!�i'�C���u4��<�]M��a��ǉ!H�_5��3�ǥZ�<�K��u7/<t�^��LUj/?��A<��L�G���w<R�KD���\M�~�lTuò��~��C��9m�X�˝��ݸ'lü�#ő�K҇}�	a���MxV��k9qj.\*3l��6�3P��e��'���'�ҽ��1��v�����O��F��
��P�]�i����-[ӵ�a�$�/�Eg��A�Y��cےV�\��H�,��66�����:
z\^:t�i�������:�����d�0$*��d5�ܨ�yBx �D]�Ud�8����rNR�-dtܵ���U:�#}5@'Q�������sA�\���m]��H���:(��&��#�������7����i��4��O����<�������d���Q�4*b�*fi�O�j����t'�(��p��]+;�Mg�<�x���8�w趥矽���#Դ���#��f�t����T��.4M��xvw�}%��@a��1�5�qi�G���Ly�K����̫�^�k<9�P��҃��C�zC?`���<AǞwEyg�ٵE�8j�-i4�b�p�oO��M8hn�����{y�h��+�'���,b'yu�G����M�9^���<;d��S/�F�P�ǹB+PgR����kJM�V��6<�`w���
۱\y��]ʈ���'�#8��s��YK/I�b�����ZM5ʩ�^�Inh���ޥ�f��wM���]��I��})��w!4�2n�����D�&��>%4u�x\��Q�n;#���I�7_B����;�}�D��"��1��W�M�y�oS��� �M�yui��Uc.����]2�yO���$����Hf��ɯ��4f��:$ToK�'n��G�
a�e!��J�����p�_�7͈M�1�Q�5bзH�N�}�cu��s����љ|�#3����x��_I�ؘѪ�Ɨ3Z�\l�8���#�F��v+ga#9_�)��Zh����у����������'��py'��z�{G�&C�תе]����e��o "���Ҧ�dD��Bq$-a��U���t��1Y��=A�%���e�zt��;��37�xa��[�� ����p�WG�-�$�6*3$�Q�x]u���H-�k9�Y�+���sW��E*�Q�|�ռ_&�:��Z��;�eܗ�G�=>,�֚�l��/l�Zg&��q�MV���X˱j29�X���q�p��Q�vs�i��\%��M�[��BF�kU��|�~���.ULh�E���Ux �O]�E��x"�� �p������3���k����_kKL�:,uN;
�jBr̹�[�쵛$�� ��"�I)?��c�`�'q��ɥ��Ȓ����6��w��]��{��Z������N��y�J�������78�usQՐ�:���v8����9%�YP�~*��=�3ч�UTq�R<���_	��#o��/�:�����b�5�=�6睪�D�f-��1��썦�t�����Ee������7���bY�J��ہs�qD����sx����wOg��з;�-(�޸Z���9���%����z���a�����4N,iDRd��F�jL̴�|���o>��,9QLy���:���M��NJJ��"s�{�UdU��?g*=��.����^8�8g$�SѨ+����gy�>�ѫ7y�AÞ\��EP��I5�v�9��Z	��p���Α~��j'9شP;\�h�����"��oMz�O%�[�T/�R�(u�\�T1��f���5A�(k�f�D��3W����"���U�@���w�<�>t���ڲ�;����	�3B4���F}ё�IS}�	��Jk��ۯ��/�j'.�	Ǹ��/sP;�
�0\���u�J�Q[�j��'5�mV�O���y��Ȣ���E�=�-��y�V֒�Y�Mc�̝�������Ih�q�:�w��Q�CҶ�l�Ú�p=W�|�tW��S�G�����ͫ���/֜Z�7~�O��p�{��i)|��r)�fi냳�4yj:�N=	X:e8zF�UᒍlC�C_�lIu�Gޙv�0�!�nȷQ��1avmPG+�5{��0� Ҙ�����7.M�^T�����@��Z��;5� ��Aqy��4��T�5��f�M��{t<����p��ܶ-7diR�G/f�k�̽l�/}�w-1�:4C�������|xֳ�޵��}����=�����7��K��6.�+TI8].�9jQ�$�R����$נ�8�63�:;c�׸-i����7E��|�2/�<�u���ؔqb:Llh�b�t�X/���D?	��Ŕ����a
F��7�:�WD��c�a��iv1�k��̃\�e�b�h*v�Ѹ�޸8Y{����/2'������i���X�Y�ˉu)����uHX��oZ�sFy�����AN^;�
�I�A��<.c Ju��>W�ˀOP����^��q=�A��f�V��{�KY+0`�ηd�7��:S\وے�㶑��Y�i�p�M�PJjE�:�I' ��$'5����^ɺ���5�����j��F�[��}�8�T�5�pE
�̼��rhЕ���V�+����#�hB0OdH���d����`;���!�m�g�e(3�"��%ɷ��`V�)�n]�Q��j�J;�~�˛򸩍��Sj	���Zm]� ���'�� �����{RSi��m�^�!����N��u�љ<�)�v\�m����u1����6��Z�+²X���26��O��4f��o8qs�}wj�ӊ�ױ�ԯ��9)_�S���.��+��[���ӻÐm�n+i������@����N�߄��(�Y�x�����Zv��B(��\����>�q�8�A�.b�q+uL����w��� z�����3M8���{_U{4e.s��^���\�㬳u!u���e=�vf�VBj H�)���s&�tX�V��<�I�u�p���c�t/v\[s�\;�pe^����n�\���#9���U��7&<V��9{Ԇh�X�7n�BT�T�2�b��T+��'94��Mm[/M<��d�æ��=��bG�H��3��E�췭�«@�&N�n�m�
A8���:"tv��/5�a�0\R�i�&�nm-���ּ��=\o�n׸�!\��L��h�ۀl�+H����91�]�p�]*g&�*���n�3D�םR��nΩS���'C�_�����]�KՅ�YsrtV�Kg5:3��`լ���|���mf\�;�P�A&I=�z�2�WO+�yV����|����"��;��~�H��شĭY�(r�v+�hu��;���/Է\Z�ӕՁTw����,���M���g�
�7�y�IM��o�K�X��v��ҽ��Ż�B.vJ���A��Z-�c�:j[ꋥ�q�.�k8f	'dDM��ٴ5��e���flN�2��+cݤ�R4-����#�&>m$�DJN�s��Et64Ukέ�Φt���_Y/�7H,���QX�{���9�mENU��
)hX.�ᥲU"����YY�Qe��[
�ĉ1h�A�H�Ɇ)0�����"�3JE]&�J�&U����V,����f��+E���.l
ł�UAAVE�E���Bk�L$�M8p��VEV�Db�0�P
C���a�"�I"�X�V���L0��E�T0�PX�S!��e!FH)sI0*AAIZ�*J�#dXE�H��)u����}���d�Ϟ���^���	C�rٲB��"��8�G�W�#�o��)�=!d�׎'Y��F�|�����6�s��W��_NKO/6��*]ꠒ�ĩNE���K�	ow6nu�#�`"DjK!�)��\�UF�V�n�۸�����Zǂ�y����^�c{��ㄛ�U�<k+��Xm�ʚ.��	�4=�*ar�=2$�MV��c�V�3�$��?=.�Yʷ\v�#�N�]:.�12��:�}]ϐ��h���1�"��M��o�����Y=ژD���������ʸF��R�/����0�vj�E�W�]N9�j�R0#q�D���gK�[״h�;g�b*��T���s$9�3bR�G>��/�^����+jQ�U��oZ���`5�K��U�����6�f�E�v̸���Q1���;�MU�vfp����1��I}���� �������<ح�V�f+��9c��ɛ�g-�i.7�:���z[^�j�=�dǜ^�k�ٹ����댓vfv�^���$�N�(�ξ��N�QC��DnV�>���3P������>uD>�N��^� �u��l�uS��0x��thu��$�1�iG	ƕC�70�|��;����޽W4��9{q;�f�gSu󧺶+�b��%3�IH#�%N M���74���2����O{�p�n�t���5�VVp�y4�<����J���#2*67�|��˹�l��'SX�B�؉�9�HEYKu�:r�x�pk�p0��cj#)���wk�l�Ԩu:&(W}X���-Ց�rn��%�⯌l^�wX_�8-z�7�>oj8k��P'G�d_n��c�=��;�:0�`G���A�M�|�"M�A���s:��nN;���U�ٕu����Od��rՒ����s��UY�:b�S6�9,T2[(���G����N�'��k�JD�1�+'�!��.\ޕ �4�^�Ʈ��q:�\�y�dry�-��{�]kS�{i��[ڻ*���SV�DT.�s� %5g��11��Vc`,��WU֐|ZE�mZ�Xqq��g��[{=�/,�5VF��K�S����%`kj�E�7��k��j�29d�#(�)��5�� �yQ�1��&�&qO@Ș޸sE��.F��=֕4�2�Kzvﻄ1�$�5�'j�&���]
֭uߨ�'DƴԬ=�i�t�i���o(;Jt5������s� g9H���ɨ��2���
��q�r�ְ�fҴ�]���]�$��QVٸ����<�_f�/�7v�2^K��^EϢ��B�j��	�![��W\��u��ޔ�fl�V;��Z|���IM�d^�S�B����t#*Ro'�c�J����g���4+uGA���fńC���vh���.�Z�ƽ�˜�$��D*������a$#�/����d<�e�Q7�f���N�ԖC��v�Q�#/*�J��ҫ>�*1�!�s�r\���;�Ӿ���]P�3v�{�__��J'�ޥ���������wKA�3*��zXH�eh5ei=7����`�2��>�T�Onm�]ኤ�q�f'��Ć�D�$z�+��#(�Je��#�L�B����f�i�[. �s�A����b�8��O�d����a�����s�� �
<捵�[�yo�������+<��E�L�;��f��u9�F��u�&6����z�D�j-��S��m7�LB�mOo��r�S�7v�o������OAR�<����+�b��
�\N����Ňv{-�\��Z�V��ǟH
�	�GI*c*�D5\<+.˨�Wò��W]��B���wd ���j��bC���ĺ+���\��p�(��,s���,�L�D�.�ykWb0�����Zf��J��,?9�&�Tv�F��z�p���rŇ���/��4�@=`�tc�Дf3�Jn�iI���UO��2kMđ��GQrؽ��Z��՗�Y+��$8�8Vـ��6�-��'g����N�2ܬ�+��#>�y�V1K���N.۝ns]D��m6"w�dfԻ���-;�sV�X0K�яQZv�z���{�9]ބ[��n�~mo�p^Q�wӉ}g�#1c���k.��"�GO:t�v�B�J�3���k_��S@����^8�n��n���7��N��b0������G*�]}<j�r'B���{7(g1���ŵק����Ԏ�T2�M��e�P�aUI[�a���m��1]n��ORK7����S�]g��!Q�Qh$�b��D�9�5�ۿj���o)�#���m� ��u:mX4�����c2��v�,c�(��ز�D��/���kKa�q���"u"��ƹ}����sT�ط�ﾼ�b��"�U��Y��d����bU��W�x�T�!�� H�tE8�`����f��%�}u{3��9�]�oY(�s--'T��Bi{���*^H��#\��Q�bR)9�;|���B�yޏ�0芾������:�Ё�g�G����M@�f
�X�d���we�Gd��|.�a�vO�T����'	��}��{��N@��\eF#p��+x�ܭ�6��}���wA�}W����
�X�kRq��d�v�Sq���f�-V��]Uۉ�G��/U��ʰ�<������g��mu�#�efҌ�8��7�4�[Y[�T������VI�����w����2YH6_��������Y��Q޽TI���1�oU���ٶ�^m��F[��k��8����L�3T�&�ns�L/7��_���3:$ͪ�I.��]�ı8��X�<�`"sRY��lo-�}��h��.��B�`�,i#��PmM<�C��#UGqۚ�aF���|�\�1\�"�%r�D��]������R;�Vy��B�Y�r֠3�-�n�4���|�o�E�Zz�6�o�8��*�j+v��K���Uh�h#�99~��K����pJ"��	���{y�L� ��Ɍ���}��f5��������x<��O�����,���@_u�y����cI垹3��^��xT���$��gf�&�����bfӋ����CV�ɒ�'��AȺ��:fN;k��-���F���>4r��{�{�9�mj����T��FŞ���K�����w����=�ǎ�|\[���@�.1�j��c=:�+]���B�4z�Ъ��r,��:�6�թxS/gu�b�;�K���ĝR��2���s֫(��v��<�.(./���fƱ�V吊��+��	��s^�4;V$����Mޑ	F����W�㭥N����J >6`����9�x��&t�G)6�
  7����װQ3v��W94�3c���\A�����+6s1���,l�E�eб��W�ά&���1�L3Fj��/�Σ�i����$a�>��2��E�Ȧo<�<'�S{}/�Y�I��m��<������g*"�̮5ھ�f.�5i�㸔ڈA�hL�����OY�ۧ˞5�������9���.S_�f���r^a�A�;O����v˓�WM�]�.	��?:�]#��;��V�
AP	_[�R;PLJu�;qSQ%�d�g����{;���wn6=�T�wJg���ՙsFE�����l����^�ި��*�[�W����ĸytw��������t[��uA�F)�\|��ô�j'A@k{W8�أ	�6��I"e���.�zgGx`�jv��e!�u�ۑu����7�x��C3z%���>��ĕ�,�B��!PY��,���R)*�C��E`c4�	H�
 �`
E����)	Psd�R(��I��TAI"��E�$�d�U�X��aP��I�H�,�Ab�Ŋ��� �DaP2�`,H(Ad� �	�JŒ
E��Re�RLR�`�E@��D ���e
�EAd��g��v���Y��GNͤ�kVy���7�]X���I���m&�m����ЪQ�� b�
`�>��Wb��S�:�yX������{����@3Z���Fw���g�&Oc*ߍo>����v��N�M��h�#��y�W�kWju�`lq��h��\�Aq�91G�j�����+[H���*�p"�dH��wN�ݗ��%0�u�l ��=<O ��4��k�1��3��;Q7'VLG�sh���P�KM�}}Lfk�~
��߻_�Y�aq����Vr�h���UY��M�g3�;��a�(���jl�\:�ۓ��Rz3	�J8Fw#Jr��8�r��ܫ�[�}�_v_7{r3荍��5�����hBeoN�X�z�q�]�����a`"�uO[� ܚ.M�1m�3�Z��r������$��iuB��ܦO"�ts�o��I(���;j/i|�7N.��U�-�a5"FQ�[%]�P�0��ߘ���X&�><~�S8s�8��
��>��y��9��Ý�3�н�Y�fĖ�eb뛌[k�su�Mo��[I�۶q��rluF���Ko#5_Y����S�-	������� S���a��	EV��^�{W��U�U�C/�'�
�۲�(	ۋ��:T�5d�c�:]�C#Mt�2��T��q�U�ޮl���(��N����s�6�,<���=۹&㝬����y�Ý�-�!$��~��
���Ҿ�]�� �ۈ�HR$�)���N:KK�{�p���뵶E�,��>��J������e �:���/\���5m�Tj/�h�EfA��r|�L=5/A���]jQ�:\QO�Q1���j�ĝ�\��=Py{����A�o��Q���vt.#>�j�)�o�����h�-e�{K[{)
�s35^.�^t�[i��Q5�XNݙmK�03�x�d��H!�����J��T���/bx6x㻭S�kx�ܖ�p�Wϡ�v���j�ط�/bM���I<�S���3ӻ<oc�h����>����y|Eu� ���X��&'��G|����R���d������2{�{
�|f+W$0:�֔�;���ϻ�wأ˫R��U��m���G��xN��:���S�'��W���,�rt�hMv�)i0�d��I��9�����4SRo1YR�Ǆj�=��������x]�O^c8*u.w��Y�,�gܭ	m��'Y�ˡ�w�n_l�1�{��
َ�k�9�͉I��L��t�����*�����j��zRvRaי�ֲ&��K���5i�-���y���eOz�;զ�����8ۿ2�[��`���u˼����J�J��W��~�+��\Z5�N"a�</!�ޝ=�)�"�	�(�ޞu���^�6�	s�;ΔB��jסU�ɐ
x�R�i�OE5zT
v\幹�跠�,����3'ٓiO7���Z�؉
�z�1슎a"�."�vU`����ü0�2���T�t�N�\6)�y|x�T:�X����)OM����I:2�Ju��po�8���Տm�֫��;���I�1W��T����U}�P�"�i�F8�a����uPé
�gh�|P�U�7/����׭�[}���/&���T�|�*xƅ0_k(VoV��ʴ�bm�Zf��]S �5�M�̓y�v޴O8��yu]<+����F�Ȕ�s��t�Ki��gD��w%�Z!������@zi��c$.��/RD6\>㷞���]�iFѳ��q���p�Ǹwd���w���ֿ!K�VE�A�V�j�Ku���z�*R���oZ�c����,�G9�F�}%g)���br1�{�^(j�xc�𓭴�u-<�C�}����7��y��_kxB��z�z����W���)�~�b�v��|S����T��N5f��<k��#-���In*��:��Q�;ĊO_�"�V�����6������c'�/�9�]ķlۡ�i���{Դ�R�+�g�ԧ}¯m��Jآ��"�ݽL�4aX���H�*V\�h*ɽ�Z5���!��3�*.�B�}l��4zK�r;um-%�uݗ
�:j��ͭ�zo�b�pr�~j��`���o�L�,������]�tG8�T��2e�.)|#I''Dɒx�tf�a�>đ4�o��E=��Z׫M��n��S��mo]I�y�����(�:ZLX�sS}M���a��&꯷��<j�κ�7�ϑ[jdd�LLfl�xk�:�Mݪny0��\�.��GK���Ze�Ě8.�*t��'�� WzN�|nC5��wd�f�d��{e�%D�.4�7*���W�$�����Pn�NZ������5Y��}��k����4�3���z���I7}S�4B(x#�nqԲ}q5k:z����$��/T�/�U͉c�d������h�vH�sqȔNu�G�l��yqǅ����[��,I6B�r{�;��I�3;�-o�[u�s�-�p�(i\����$®В�3����Ǒ�)���u�X��H�Kӯ}pX�-Ax�N��'-nZz��.���f�����²��N����-�]�|��O.o,�&����
�:̂�Ϯ8%��ˎ�R���i	
���������0��5�1ѐ��Bza7e�3V_�����h���rJ}��ㅨ0�JV���Vt���Oū��ڤ���P~�7�]�:�|�WR/�@����lK�9�24�\Y�r�3YR	��"�	�eTZT�F�5���[��_
p�:[	C�r-�H��k_t�]��F��
+�NŸr
��)nĽ�ǫ��'�zSϷλ$��y>�/�4r��s�� j�'�x	�;��A���4� V[����x-^��P��ZL ��쌌Y����q��F��X{�g����E^IU���r��Vо����6�-q��|��z�T�*��t\��h�s_a��u��[��,T��Ec�z���y:<H�zUT��jJ�UUT�|Z�@/Vt�DI ��"ɰ� ��iQJ��qfE��;��m�hʳ������1�-�m��ZRI�$�/i$�H�UH(�o}ɍz{��'����
C�"z����'����Y�WHb1�ۭt�R�D�b��������m�f|s�|Ѻ˚���e)s90�ג�βQ|�5d�ݮ�Yi�e��.Բɜٺ��I�TXU�7m�cI���I �~m�vvɭ�D��0턒��&���*��]��������'�=H�ag���v���0v�J���"H��G��[��z����.h{�"�#�2R4�%�����F[��E��,�������r��T(ҽ�,x`�%�+��%$�N-6JLk{]�^��f�2"HQ뫧nRI��UU!�4���f�T-r�:>����������1@8I���*��������c��-����Db-zT��}������8H���>��na�:>ag�?��?#����������>+Ù�#�7z?Dw�Ï���
q3���cB>=�z�|Y�zN�U�����p/�I�3�;�ω���@8��IEk���%{Os~V�K�O�Xm����ʖ���$B�\����$������ZUY���%��$�̦�E�4f�rfc��ETQI�^]\����T�*���I��RG7Y������b�%�����g������6M0ɬ�U��#�f�$l���t{�:�v$�+��I�JI(�8��R}������M��Sh��qN�\���s�{+%~/E(�����n;���|{�/��e��"��@:�3�8�W �^�Z� ����+�D�I���yZ˿s쏰�u��:{��o�B]��^�Q���੬S��%JQr^��tpPǗ�<}�����#j�'�����kx�66�Lp��p̉ ��GZ3���N����-ݞ��в�M��q�U�Q�f��۞�#(,{�	��ʉP�@?�*I�/<�Ǘ4l�Gey�7)�c��$��:���)3L��q��d��%fY&���/�<o|3��*�(�;����77�n�O�.�p�!�u�