BZh91AY&SYVl���߀`q���"� ����bJ��               �r(�QPQT���j��T�T �
-��)KZ�(�HP� TKCPEkZ� �����iR�l��R�(�^`�Ruf
D�đEB�RT�M�P���J�HUIJDQ*4a* QB��*m�R�*��S�T�DJ�T*��{��$�!p1EN* F�H��v)��U]�A[�[�
�X���eJ�����B��E(&ثLQ(�)U��u�QP���NM���(
 ;�t�u5Om��ծ���t펹ب��{�!G�<����miS{�[�[�2�M�j��M����5��R{޽kT�����\Bۥ��T��U%T7��  o;w�J�E[5_|�OAm
���yӮMjU����zU�IV�{�UU�T������J����v*��J��[����K�ox�������'��Ҫ�KV�H�%D�l(ɪ(����(;-��J�[��o}���*B��Kץ)�ER����B�R�����ǅUT����ݷ���UOl-�}��J�ZR���|���j�[Ծ���W֗��7�j�T�_M��	 �T��Z����(4�y�}@^�+ݳ�z�5R���y=�ղ�Ӝ�x5UR�i�O;΃UJ��M�޽4}kmR�O}|UUP=���P�W�/���UAT��;�ԕ�٧q٤��K`0��$�]ۏ�)@�t���A���W���r�y֑UR�0�*�u���OJ�YJ���T�*�x�xj��{1�G��EP%��y֪Z�J�[��ԭS�ER%RR���T+��(����}2U��z�QU�K��{j����m�hA�{�J��K�zw��Ӿ{J()�v���A��a���@�UJPDJ��z�R�� {��%�K��n�p)T��F�9���2^Ӻ��EQjXR���c�(1���(P{��
��JU@��*UI*��E
���@;sn%B��v^x4 \Xz���0�(۞���G��.(lƝ�l\��L�TM��!JJF��V�J���>�P;{�)9��P86��w":PN��K�[qJɦ���I�ۭ��CN8��:���u n̪�� I7� r�6ԡ���@+�zk{�	�K��gm�
�K �r��� ��u(�g�(f�� >h        ����J@� h  ��1%*J��� 4` �L���@h�   � $�* �4     i�(d01�i�4�T~�SH4#A��(��S�I�O�0���W�p>W�Q+����4��")}�g+�<ݳ���*����*���� 
*~�QAW��
��:�_��_�?計*��|���:D~�|	S��E�������?�t��g����1�c8�8�c�q�c�1�cǷ�61�8�1�c�1�cǆ1��8Ǎ��1���1�8�1�c�64�1��8�1�c1�c�1�cLc8�1�c�1�qǆ1��1�c�1�c�	�g�1�c�1���c�lc�3�cx���1�c�1�blg�lc�1����q��1�c��1����1�8��0`�3�cc�3�c�7m�c=1�cc�1�c�lg�1��q�lc��L��1����c�3�c�1��8��;c�1�c1�ǆ1����1�c8�7���c�1�cƛ�1�c��1�c�ǆ1�c8�3��c�3�1�c1�cƙ�1�c�q�c�1���:c�q��c�q�n��1���1��c�ƛ�1�g�1�n��1���q�c�1�c��c�3��1���1�c�q�c��q��1�g�1�g<q�g<q��g>3��8��cc8Ɍ�8Ɍc
c �*c*c"c�	�����������^22�0	���)�(c � � tˌ#����c
cc*c �!�	���D��A��T�D�T��C�&02�2&0�����������	��0� c*c*c
c
c"c"c�c
c�&0�0'L��)�)�)�����"c#0�8��ʘ��ʘ�8Ș�v�c
c�ȘȘ����8����8ʘ�Ș����8���c
c �"v�ȘȘʘ�����c!2&2&2�2�0&0&2�0L)�����)�)�	�!�)�����	�)�c �q�1�1�1�1�1�1�eq�1�1�q�q�1�1�1�1��CSC�T�P�D�D�D���P�8��8ʘ�2�2&02�2����ȝ0&20�0&0&0�2&2&0�1�1�1�1�<`LaLd`L`LeLaLdfP�E������T��S�a&Q�T�1�q�1�1�����1�1�1�1�1����c c �cc*cc
c*cL�2&0�2'l	���	�)�!����2SCCCC���T�1�q�1�1�1����"c*c
c � �
c�!2���0�02&2&2&2&2eq�1�q�1�|`da\aN�1�q�q�{ddaLeeLe�1�xʸ�8�����8����"�i�a\aCE�W�e�N�T�aD�D1�La�LaGQ�q�&Q�P1�q�q�q�q�q��SS@�Q�A�f�T�T��T�����q�q�q�|a\eLa\dza1�q�q�{eLa\a@��`eN�GG&���G�q�q�1�q�q�` ��� 1�d\a�I�q�q�aC ����xʘȸ�>2�2.0�L`e\daOSC���8�3�1���1�c�Lc8�1�c1��g�1�c��x�3��1�c�	�g�1��p`��c1��1�i�`�1�`�1�g�c�1�1��3�v���g�1�gƙ�1�g�1�blg�g�1�ǎ1�c8�1�N<q�c�q��x��3�c>0c8�3���3�1�cc7��q��q�g<q��q�g�q�gc�q�`�1���1�g�q�c����3�8�0c�3���1��1�g��1�`�1�c�q�c��1�`�q�c1�n��1�g�1�c�c8�3��1�c8�3�c��ct�3��=�c��0c8��c8���3��3�cLc8�1��3�c=<1����q�g��1�g�g�q�|x�<g�q�`�1���g�q�`�1�1�g�q�gq�cc�q��g�q�`�1��`�1��<l`�8����L���l�62c2�m���t���0c�61�c=��c�0c��c�1�c�3�c�7�<61�c�3�c��c�1�����1���M���1�c8�7�1��c鱌c�g�1�o�8�1�c�3�cLc8�3�c�63�c���:c��q�c��g�1�c�1pL9����N-Qw����Zi�����l#���X��	�H1���کX�TF 2��I���	�0°m�u��I��Tӊ�HkIktIwGU
��6e"�#f����t캷�[G.�(4�+)���U`r4F�:�Ό����S�/F�A�p8%�"�����8Yfj��-�ݘ�E�p���t�;�BR��B�{m�x��2ID��t�:Na�y)�n�aq���O���.�S��7��q�R��9/��SP���F�r��b���,��1���OCc0��S}2��\�Ŗ!����V�ZB$jB%�Cue6�`��d����x�ǧ�%�D�7�)�mCmTE��Ź&G�U��މEU��:�*�r�q Y���b�%q;��,n�Y�X���6.^Pʬ��nVۏ2�r04qM6����F9��Q��X]��):���L�6�m\��ol�( F[j�SZ��7L<[0Pj�lM�HJSj�m8�^4�X�wٱ��������p�ז�(&h�"b�re��&ՋK Dnks(����U�3D���"�y�0KҶޫ�Z��tS%ط���f���m���\�2�"[���Gw�eۆ�˘)������Tuޕ��뻉Sy��x��:�9��<�LE�F�"e"��Y&Ɖ��S��Mό
�����͎�I�VLY�^�6��T�;���$M��Щ���ӈ�e�/C2��C�V�Rd�ԅ�f�7B);�n�쨷U&��b:�u�OM͞�۪l�݌�^�WFA�iނL�>@�t\5��Q�%��.�S�,�{�Xܤ�l*�ɛq�
�����6���R�#B�FV�Z3\
=�u�w2��D a����U�f�Ek�"��]��c��a*�X�,��A_z�K^a��R=G.��f��V���VÃwV��X�&;r*��Z�Uj�6N�z`ǵ2\���'�.`wIʕX��V���73ܛKC�b�V��$Z#��˘�=�N�6�SpQ�&�Ӓݨ�%������

�PR�;"��IV�*Q�{EBLځ���4�*W��NYf�{`���1:d⣹��Y��_�Mn�=��;y@�&n`ܛ�J�l!D�Ec�2�6�Aa���٨��85iT�M�,�H���:�6����&�W,7�\�cn9$�7TPѵ�^G2��i[���s
���)�^f�\�ś�T�$aLӘ�����,Ƭ�nj���	�	aЪ$�1&%�j��m���P{���Дo�cj����#~4m��=w��ԣ��E��m1�2`�_-f����[	�6�IY���Ԟ�����4l6���[�U=Ȳf��;6GV2*�eJL��dI �"�%޺�Ǎn2�ge]��"wsK�K�yb��Di��d=V7�ua*J�n3���Z`�FW.�ݏt=v��ю^��Vѐ����7�F	ZS6���ױ�T��im	��U&�[Tުg/�]��$�2�T;�u��4��{�\�,�"ؐam�7w�B�&P��ae�[EY,#�Hn��VXy �oQs1�,��ʟP <X&��[�El���.%Ybc�b��Y!�w��fLպ�Y���E�N��Ē�Ħ0���("��^��aت:$-�VK���q�iԬ�*ܽ�E4����tT��2�ۃhV�*�[ge�)��#�����E�k 9b�#!�ad�*�T��H�Us\Ɲ"$�1�:�d���!-^�K
�s\�G�ߖ(��p:�nn@�oFrm���Ӭل�;I5�H�m���Jcs,Zs-�EU�F�d~�LLؒ8d�t2+t5b��6f�{�rU�\Nn\^m&��[�T���U�L^�Z-R#Z!Z���.�1Z4�6GV�Y-���)(Re��+ߌ�;՛��VwM�DA1��p�w!�R�\.��Je�$hl�-���{�n5�+R�%{H^,̌ϔO���(��HQ����`R::f�QV�L���f�w�t�k��l�j�Ҽ���HN���7tj�z�u���m�J9���h��՝�Q	Q�g����3�(���f�e�#KV�q���f�Z��$d ��Tc]	M����^�R�Հ>3+HZ�9^;�Uxmr���m]��0Yp�ى��4�JE*�'d6Z%-�����\-*��9�P�n�#�C-�-Xk.�݂v�e����j��*VPtط�&X����c{DY�S7km�[�S�[��r����^Ø,��f
a���,�;OC��f� �;N������2l���n�-�wEM,)6tQ@�a��
U����Y�C��Zz,�ON�vA;Pciim�%1��F�Ef�s.	+Uk�����r+s6��(Lwv�T
!F�%RL�KٗbY��Su���89l��B��9�������MG1���r�9�2-̙X �_تһz��!���j��� ��j���n�2�چR�N�B�i�};&�$�����y͇��b�i3e�O0,֌ו��A�kEm���1^V�Q��G�i���U6�\6%�5�V��a�!Y�����Z+]�N���A�m�B�i7K]��eX�&1{�-�i�&GMø�s��.܈�V��!ݔX5ۧ6�����*�i�)6��{r���˔0�;"f	�@ŤU����)fV]a��o�`b]L.4V�ae�t*R�ڦ�M'L�Ed���D���~v��ɡʖ"G�w������Ge�	`o��Ŷ����tݗ
܇<���"�ڠt�*���l4t*>� xn�HQ�U��,�z��m̖m�mܩ���V��R]�m44#خ*eۼ��5�qY�N�&�Y���ӭr�
��8�r$�77\���}`7p������D�;`�!5$�&��X�1�Ft��ث�Z$b�Z4[8�X2�Og�ܐ��m�v���UT��0�3UR��5V���k� mXu��]D	�0Y��=q����pf^-�j�f�[�Х�tr`"��3!�f�1���.d����� �v.���V�(9�tƧ�L��e�7�J�䅽ɂ�h�)�d�����ģ��f�~׻����b�c�v�
1&��qm���C6�H�i�K�J��v�u��2*f��9�\�w+fȯwYj�ג�l�*]�+�wF+Ӥ�ܥ��]9GT]4��f��ȼ۵�E������H�ݮ�](�5jf���ų}�bpB�\�2QIJ���a:4��gwl��خ�OE,n�Ga�[t���>� ����4���w��w���voFŲl�rklB�mU�N�Q'�(^R�5nc��[9r˴�'K5�Q�J�ō0X�)x�ކռT��gEAC#��mR���[U�cWNT��)�RF٭�Z�$xwe*�h`wWQ��K��潛q�{B�refڒ�֪e���jL�w����JѨ^���7~��M
�]�g7\����o,2c�C�_K-�RL�{i���nX��cF�jT�N�-�&��P�by�ss,��
�Ș�B��j��i<���U��U1Ww.*&�1�
TM��.�a ��<��KfR��.��b�۸��4�Q�y�Y��*
{�l���i�N�f�إ�Y���$͑L�C���gd���-*�[�s�r�tf�І&�w�û�HdP���H�En�Yi��d�ܳb�LԪf�m�J�!7��37	j��%l[�g ��� �TC%̦q�/S8��f7���C%"�w�q�Y�g,V�I�3K��"��B+K]�i9S�q� ���`9�G��31��ٛhd���eV�R�,a������(��'Sw�W@�E�"�`U����"Q٬L;�#KV��Y
��v����0�p�Q٭��������yVPS�\$�J�ܬ�kyV�(�������(�@�N�T�2�۽���,7�uӭtpǏ@�w˃U�Ǫ���+8܆���yM�f�Zf���5$��ͷ��6�;u����� �kp�SX������O�D��\�6��<���4���tr<۶�׭�
D��두y�W!���Ԟ[1���ꕏvL#�s6�ud��Y�T����Uhy�Of��â��P�W����鄪Sh
"btB��ebu$�gw(3��̀��k3r�H�"S��"���1��\7�f��ʴ��zɷt��WljЗW#�[�ˆ��GH(c#X�-���e��rN��6�F���I�i��U!�!.�S�Ԡ�^cVr�'i���f骛f(��l܈�e�k
��4iZˢZ�y1AFY��hR�͝,l���̣�S�p,���r�%(`�GK���0m�j�༑�5j0�!X�T��kY�p�W���� ��K�4P��Z�oj<S�r6������R:��&���	U��e�Q���X8ʃ z�Ea��A�R���5jղ����ْ��:��L�olֆ�n�H����2U#�dZ�8��V�$�Y�m����6�n\�GoF敊�@��i�l��kC��K�řv+J�Ԑw$:�!9bb׸�óoSK8)`0�mr��hvM�!�
k*����ŵ���x��b�K��1�e�\�-I�f���W��2
�/8��UF�n@j��OK�ʦu��W1)����cuەC�%�(P�c#P���m������*�mn�2�,r�Xҡz��*� gT!�ۉ3I+-�;NB��TF!wb�7ZU� d��*��!F�'��m)7좡��Bfr�U�^nR&��Ջզ�CI��PR��M�r�M�!����Ysi9��j�df�������Z�Ҧ��*6�M�;��u%ָ�I��qA��(6m��I���V}�IQI�C��/��*ZCW�t+E�<:�*�M;�Jڸm�W2�*�M9f�H�[�b����b�,W��w���f�a�i\�-�ر=��"��,�b��Ѫ�Q8���K����S� �D6�Yik�۸w^�b��S$��N<Q�0��8f��h�4d��Q-ઑ��ʵ�ݝ�{���0]X����sbh�@B�"�@@�cE����*���B4��%G1`4-6غ	P�v}�b�Ęx�];�ܚ0����A/��e�Y4u;�Sn	�*�d���1�U�t�kC��0ܹ�tc�B��
���^A.k�Ki-"L[w�j�0�U�m,��8�V�
x�.ˬ6d�EZ�LU����3彖E�ODm*x}��WBy*m]=���c9��(Yoml���J���)��knK��JZͪ��ʆ��q���F<�;xb4b�;45���o-g����I�ct�C*썚B�yc3���x�nɉ��C"F��dj
����MsB������P�Oc��W`���V���:��Ã�7Mh�fU�i�g5ށ7I;�:�Z}�'ɉ�囼��	"Ԯ�Սn:��O���8�rާ�i�F�uŃ�RZ��������
ܻX6��d�����q�}�8q��b�F'>����5i*F��c.�ʷ��em{��WUog�:��{������C���+|25��ܮ1k��Ѹ���E]
�J P�-}˦�ѻbn��vU�ʵ�&G�'a�ˑ�N9��./8�� 2�ɰc�{���������ʺ6ћ`г�ܠ%���2f�wGq�wQ5ۚ�2�B�jg9���{)�)u�cj���bqK;i.g�y��͵6�/��PACY\�enf�[M;��q['CE��j�F���+;��:��īc��H2����Z��8H2�4#o��@�kt�bՅiOj^mX��N�\9����#�Mu�nUJHJ�J��`�F�o��ؠ����f��׶�|��R�YV��ܼQvЯYfa���+U�8Ťum礮��v��Ƃ**jԫh=��!�r?�Ђu�󈨇V9f���`�����i�lUTd�ۜ�J�e���ԥ\m���g�j��o�Kuan�J�C]��[[������R	�Ѡ��IgGj�mZ�ɗm>�T%���(�8zWW]V�sqѱDv1��^�mR�6
�����R}����Ƃ�Rb��Վ���vD���b#JA0Q�w�)�Y�N�#���UN�8���a�_;���u�|�
�7Y���F�:�}F�W���M\�veWdcr���싶��V9��B�&��o��m!�s������gw=�B��ݣ)���eX-�{����njYJ��F��A�+,�ư;p�t����r�xU���:�
���;$`�� ��U��L�+V,xvF�+ ��l�Ltpݶ>��㜫\�Kq�}_mj_o4�uu�=Hވ-]-�v��.B�ܻϦ��~���7�2Ս��a8]$ͽTÿz��Z�t�3vӃ;���K���ӺӁ�륤wt	�P��F.��]��&b����
��
ec�w`l|
�+t�M���n���.��ʺ�5I�(�݀j�n�t��ͫ���!����nv�s=���&�$�f�Vgc�[�����@�S��s��^*j����x�ho��.���E|�μi��ܴ�U�,���'hbQP]�wvX�-�I:S�,�+H*���ʼ��R��!:s���\˛%�r�P��i�����H��db��
����D�v�N�!D=��%	��ˁӶ�&�T)R�믧 ���[Dp�Y�:��s˒r��Y�Wa_$���+�2�Yȩ��Ē0�O	4�G�0Cx~���E���n�(:GUv�\4-U�Sx��q� ��Y�\v�:����I�	q��=-)7tBb�9h��z؄%RC�E�YN������]5�l�A�����s�B���.l*���V@����N�ǵ�,�/+]�,�'d	���1�1�ƒg���Ms5z��%�U��BQ�:�$յQ��8�g���O�J�"�]H�b隈Sj��}�c�-p����屎�[KV�N"s��F:x塧Ma��j&�[�K��v�vJ�	c��UW���Iv{���
���.�8��Z�5B]2)�8�G5��ٷZκb�K��'w*əq�}C��,	��y~@?��a�z~�6���$[4E�&���1�j�*�t.��ړ2����L���a�:V,�]�;��؏�:̔�C�c�8gt��ڋ��!��^�͞��Q���'�.��'�A�p���%�m�o5��EC�ɶ���D��M���i��T{�v��ih*��m��ņR!�##z�:�ܪ�zۛR���%A�;\��P��l�dXB��^_qYje�g
�|�tYW�Q!Y%��ԮэeV蝓[�k읓�J����*n}�R�#\&R�4Yy��ڝ;�9��aW�SscF�za�N�Oq8�g�U���W�y��p�C���x��_L��aj�]�_:�Ա.����]��ԙ�]�c����ѷx-�,���5+<8���ۡo�������2�����m�S�ĩg׵�����9��y�C	>-�S�F軶kpj
4+���
�S�}y�۴8d��M��������T����[6������Er
t��8R���љ=-�f+��E��]� 
c[՗�P�И������=��AX�@d�E��pc���TT+�7-����y�!ކSn�ou��*^���vB��׼�Νc'c�A"������d�f�(�%�v�S��pv.uS�&�Jh�J�P*�X4��l��xom��^E������ݖj<�{����oN�PKoD�R�v7ꨱ��7i:;�UX�ub�w}��o�B�'V�.Vƅ\�M��J՜M��8Ź�Ջ[��
�K���N�^�3����SJB��Ѡ�M�\!�v����hkh�gdoO>n��4[�n�^��$*�os:�h����\�p�v��,1\�#�Ϸ���*��-��
�IϠ��6��kZ���C�C4Pc��z�ƌt�E�X������7+������7	9��U��0���{՛:���"��۪�AN����r#|3n�7�f��u��7��):�X�i�BG(~\/��{��v�M���d��L:�8�!�b���Ӄ��d��R�R�f5}�CN&�\��C!��q���U��*���6f��1�uuޱ�A�ڬ�W#ð�z���k�r���L��<ܕ[6��$�Wg_'C���?oN}n�#Ց�#�C�g ���׷�N�I{CL�Z�����JTWM�������J'�0%�_tV���GM�<!T��i���6�w�{�݉�w�@�t�;��,�d��+��B��S
U9��Jn��Q��Z�j��Z%��݇{o�V��_W7�<�C8�v	�+r���6)N��;Tm���>ʙ�$�=UlX����'�J�����d3|�v�Ś[���'��2��7[��������RR�Y/���P���
Q�|����u;;y�s�jf��ԭ��4orHg4����0;�	/��,vM��ŏ��e�sj;�k�RKkrJ�n�_aщ��\���.��m�>�[t��eϙ�_09)P&:VnM��j�
Ͳ�)�=yAU����f���|���Z�:.jE�nH_d�4ꃉ��k�<.׳�w���܊#�U�ۥ�c1�l�����3£��zUфE��ږ`��6b�A����W����oY��"3�3��p���6yTw�8w8ww�Ee�V��ܵ]�i��l�2_V��4d����8MR���XGɧ�H������'t8��֛�2+�������*F�!
2&���d��(>����#v�{u萯�;o,Ǳ�g�%nVз�[;	�p�as씴��}{#�E�:eT�e⫫E�|��U>�Ә�֡o�]�M�t@�Ln���f�o��[#8k���6��/��7�����r�އ�`z�SJ�a�Vd�Vѵx�����b���㳶�/N9��P�&t3.T��br�}ˁ���AIo�k7��������p�"'Iތ���q%J;��x*s���2�A� )����N���2m�c�x�V�+�˫�W)�: �{uݺ���9���#˷v�X��7y�t�.C�G�r\bq+��x��ivT�.i�S�x[z(�/�'��ŉBrںo�{�%��ܬcm<왚�˅�5 '��UF� ���4��uu
����������[�ҮjtkzY�_w��D/]���`��Md����]���_-��gf�
*[�Lh�3wj�D��ܸ�vi���>��l��f��Wያ,]�In�wm�Q�S8$�΀��^<k�t��t7�¼���S����d��pr�5Y`�.�R��C5�c����^qw:h4�ԍ��h��0���O����+�S��gj8���s�i��q���N���bI;	�g�t�oy�yQ�,h�ա�{$�6��xnV�4W�}p.�ؙjU�O���/k�7����H���Gj�)�6,e]�7��q�5>�*�r�j採�Z:�W`w99V��i��b�����hm>^�Ѽ��XQ���V-�;m�=9��lX�͖�Yu�r��*e��YIʱ��B�9N'�U,$G[W��N��c��2��b8�u^�idO����a���\���^M��B���]l�2�N���EǶ����)L^���S�ݾ��',��o�p��s��oJ��['0`j�`�6��eK�q4jotKfᓪ`�U�V���eqJ�q��1f�F�_M��[J�m�x���8�u��FӻҺ
ߛ���R�8PF>�,jMv�ʃJ7��;h*V���[?6���%}����ͫ�x���o����݃���۵�oc�Ww���K�˫��ZHh*���>�ׄ�!�P�aw`YywyP.I�LS훯A�ƹ!9#u����d�6���	@�V]�e���n+�g�է|�N�[9{����*��B�L3��z���m�_=�L�U�����{'������ym�([K�Ψ���q�pXȥ�٨솶�i�v�X�l�v�&u��t��U���Gx��X�L� 9N���텊�H��C�ڊ�26cs�h�0�R�3܋|�f�kU�kE�������C����go�*�WT�bN�F�mR:�B�+�{��n��ʜU��V���Kt�2�-��2��C��+mj�5�})r�P��A�M>}���Ӹ��CBƷX�o`�޺����|�{!�{���P��u��`O�T�3��I�T�7n��H)q�5+w�fT�>Y��6�5��F�����z�S�%wUr�s�$���r����Qfї��s�wN|�=���<�}î����.�V�vj��t���q�T�\R�kЗ�*�ya���؉�;-w�˕�]���`�B���ܰ�~M,iǴPs�i���>Ϋ��ǡ�t���p;��O���70c�� �����25�+O�a��3/��u�z��׼��v�eb/�� ��F�v��Wc��wU��k�X=�.�t�!�1���0r�8N˝�`޴F��.�z�l"U�{YFv�Z!���M���vrZ|8�̤�0t_r�|�W��W�Ս�/:�7gBڙ���3[k�7���ђ9!���t&��o0�j�H-��(�&�ew��gk�։E�����^:5�n)�v��t����Z�'�Z�� �ʗ��
���	�`.�:��r.y���k����V�k��6S�|��Ry����x��Z���R������c
Ә�fS�&L��^��f��b��+(`.�a]��CY}zՈU�^wj㩧���сj�����2�[�Ba����\���;dd�t���3��):LK{H5Ⱥ��n����ubV��)�UJ�6��{��!�ݖ����Bv�����I�,��_f��M6���9��}�cN8��v�Gs�\3t<w��G�*�p��t[��wr5Y$H\e'uz3U�
V�w[�!�/ZM۹��6����U��N��-w5��Y��W��ל���X˻8 9Uˌo`����GWk�N��R����2��qR�9^�d��M"�K�A���3<�%����G�8�k�g{��Pwz����T���Z��:)�o>��-,$"���e�s�V��;�o�%U��Qi>;2�j��)�kC����k�grU{I�t8�Ә8�x�@��`�,��Yϴ���_>����b���7��rY���v1���@")���5��q"�%cV�r�>ݙ��;֪!��tl"�s30i��:�n��r��	^��&�yCeݹYY�.�"D;�9�
��f�a�W��ap�ߝ�����Y��<�lNT����r:k�Vi��y�H�;�TK�4/�[2�+$��L(���%�*�6E/�>�3�g>�&��m��%]3NgV��ݳk��1dU�ӱtt&̦�:Μ�6Ҝ���yi��\����.�:��אP�\˸7{��a��R�rx�o.�+�}u�3ld�P�ÖOXy���l#���%�n�ˏS��r[Z7]�N�F���:K����u�����Ltb����#7�\$��r����U��[n�0�j�b�wo�;Nv壊�voW��t���8���g��WM�)��&4�-9�wg!W�d|o�5>׹Y	���B�V�4֐��c�d����ډ��&A<�Kۢ�gKX5Q5(��:̗ȐZ=��N'o;#�N{2���.�r=���kM����WE(qC˹��
P-�iڷ���hv��V�o�3��r��­G�R��_�j�:���ѽ�鶻�T2r$���c}l�U;�c�m��|g}qU�n��1ڲ�H�mD�",U�.�U���<�ۖ�淓+�b�:�7o �f��_t#C���Չ&ylKCXW}�떮�R��u�3��\�M����\�quA�V��VR��j�iK/����W&�$%kTiG�Q�J�Z�צ���=FT/zҫwk�P|�^����C<�3�ؐ��y�9ۮ�JIw5�7��� ,>o����#g1�{)�E���}�\���T���}rI�u�i�t�n���nA�P�2v��wP]H[[��7������i�黹��ng]Ѩ���\���:�S�dG-�}�\��p*�j�p��L�giC�d�u�ܵS۷-V<<��;yٽ�?��^�ƹp�bn����!ӄXY��:�uɓC\ks`�{���45)�;�k����Z�;���R��Jt+�<����qu�}�(���%�Y�3$�;�:Mζ�I��vA0w��$;/ ����p=r�{V\�1�s�]�Ď�7q�D��]�ݱ�۾%^t�A^aҡo.�����U���E��y�E�>��+�����Lا*�|����91y�8��y��Ӯ37��S^.b�����'���^����8I�, `���^a(9ِ
�~��A��Z�ꍡL&p��yV�,�1�.��wf$'�):UM�DS�(!b�dq���{J�S	�~��Q�*sD���떹���J[m۾�6�^cnn�
f�*!rD���Pڠ��|�Ke�j�i�oh�XAN�A%��e:���ɁV��kB�H�H��H0�&&��bNm��֘JvL�K�O�2��H�uA�2(6����Bm��9!`و��4KuK�ϲ6�+�#����U��%�CN@nS�S�-�8Ĥ	1)���e�����,�ue!�z&c�.�#Q(�A�q������ۭ�%�NЖ�%�b�]�B�XAB��5q�K��cm���PI2�6���Rv�ʃ*�L&�%��9�aЧ2[.R��B�E��'���6�̧��fX,QsM�b�4�n]"�.��r�����3/���h�"��"��O$je��H)�[�V�T�Q0�P8�|�%�ě��?*>/L�D��.i�����&�n�R�T��n�V	ۄ��I8F �eq��'�
4�-�RقPbS#�$��8��OA;�U����q̹0wHк��	��v��R#
sE�������b3R2��)c���t�
7�H��F��D�2Ȕ���q����yCS#�:%͔Ŷ�K�ؓ- ��&�?$W!"�tBH�����n$[x�̫2���LTŦ�p�:��@��MofQ�փt:�?e
Qi��l�eUi��B��a6,.\�@�$Z7M����I�����3m�Ҙ�P�PzD���Y̚�e�NЖ�%�,�kI]5��Bü�)�F"QJ��Щ�U
Cc4쪓�0h+���!L��{�'lJC
�SD�kd�S;-
�����k��t�ꗫ ��Va}!�U�A�L�M�hч�m43m�P�B��.�d�G�q�e�(-��j�%�HPB'��rb%���k0��A%����Y�f�ڵII�h�5N�.���-�����R�h̤�Y����	)�Lj�9�A*�A�)�H��@�Mh���6�(2�$&CnI�B�� ���(3|��%���UR�őwX	��D�B�W�m
����*Pa����hf.�fq�b��r�79������g�~��* ����&��W傟�� �*��7��P{�����k��u��r?U���?^|�Zu=�h��+f2��l��B�(�[�a4ha��vJ���̍��m�q�1kX�'fv��f"$�	ŒQ�vպ�� �¨�uZ��5BY�z�_=f2]����7�L�l��5�O$�ƵVk���<�:��	ɪ�/�(��c���g,X�U:�h���`�boN�b|W�'a�5IH��z:��sgx�1I>#�f��˕ovgcRuC0�kj���v�^���w"�\%+�/�o�Y�;�6��Mz�^jћx�u���B�q��ʚ#
��WJ��¦nI����d�f�<�&SM����f�9p^hΰ���lFZǳ]�g]�wjT��Uo�])brc��3yoY2ܳZW�3;:�y[���:}z�����duqA��P���tz�~W�]��X��<+��\����d��� :�Φh1C/a�ܣ�������X���:�l�M��̝DH�%n,s�tPoo[G�<!��x����J�-��}ֻ�p1v�0	)��hK�k���o�v�@������rs'm��>�xsk�-�C`�����L������뮽��uק]u�]q�Y�]u�]u��뮺뮺뮎�뮺뮿]gG]u�]u��]u�_u�^�u�]{u�]u��]u��]u�\u�u�]u�]u�u�^:뮺㮿]f{u�]{u�]u��Y�]u�]u�Y�]u����������~��㮺�ۮ���뮺�u������_�뮺뮸뮿4�(�@��a)D�iɸ��w��po�23G�H5d*�3�q�r�wne�U�W�o���Nfk��v�aJ���l�A�$��!URSwo?��zk�n��<�:w���6 �maϲ�xl ���+`���e@U�RH9e摝]���
�}��]qx 1���D�ȉ[Li!�~�n�2�f�rH�v�Sp"��ٮ���9�׋ݲ]`��>�SL�G{xph�r\�'��Qx�����U��{�uz����Y�ES��t���Y������5zu�!s��W
�3���2��/�bN=�9v\4�����Z<{�Ǯ ��L8�6YUNv,��H�����>Q�Tr�f�����n�\��=nN�Ҁ���ye������	\#�m�3m����K^}�W<k�w{�e7.]�e)��D�, im������wM��,�uH#�qb��rJ�''�I�<,@�R�Ŗ�b%I�W�" M-�{��.��j�[h6�7�#7�cm#`��(�爓n�]K'&�a�DsJ��U@ [Mъi�t���Ͱ�k$�,cL?{ޜ����P��X����u�^X֭�����l0���!���-�^�sVĎ�4���\�����Rg19
}O9cg�애��#{eYA�=�*��������{~8��u�뮽:뮺�뮺�3���뮺�:�u�]u�㮳��뮺�����]u��u�]u�uק]u�]|u�]{u�]u��]u��]uק]u�]u�κ�N�뮺��뮺믎���^:뮽:뮺뎎�뮿_����������]q�]zu�^:뮺������Ƿ뎎�뮺��]|�w�`DaJ�u�ܪ��q�F��bE��+�����
�^�wC�=n�:r�+T2�#i��Z�[�Gir�)+�t+NZ�d�m۲@��Lq�B�]w� Ih���	�7m�P���3����$�3+mU��C-"5�bg�el�x�C�F��@����j[��8��M\@��\Q�a�6��qC�q���$	ĥo��m�f�F���k%��#y��DH�a�ʌ�j��sknX��.�@��`�7j�n�1M:�JFf�tkz�4�� �22Tu���=%q���[e�ɒ�v6=�o�%�+�Iߞ���9�8�+�Q��m��Ln�+x��E�#¹@A�t��W^֬���Z� ��K�CC4V����*�끆���`��иK*D�m����D.l"�q[�Z�c*T�9���)�}�o�6��rj3n��J|�t�q 	��j�嬹'�1�y����ڝUo�ʹ[S0-�ek)Z�k׭pjr��w�����$�|1]V'Z�{�Q�'qP���(��N
�m͏}[{��e.����/9ZC`z�]�vR�e�T�e���c_Q5Z��ihW��]�ɀt0q�rW�w>;U;ft�{�&v�g����z�l�9v��lU�^�]���W&j�ֆ�YL�&�~�+Kovb��y'i�}:g7�ǒ�J��wZȆ�G��iM<l��b�h;ő��St.���ia�W(e�.�#���ok��>���u�㮼u�]u�\u�^�u�]{u�]u��]u���]u׷u׎�뮺�����]u�]u�]u�]~�κ뮺��]x뮺믎��n�뮽�뮺��뮺�ۮ�믃���뮺���^:뮺�뮺���뮺�~�_����~�]u�_����]u׷]u�믏���n8�뮺뮺�gC\�N�C���XY�՗ҭ#�վ𺺜���}w��c���뭡b��=�*�p�;Ta�³�V]C�/5E���@�Ӎ��L��u�����r�Q���j��SI�#xWSN�ڥ�0=���m�G���E�&��*v�ʏ9�TȂ����π�p��`��)=�"��%�0j�����R^}�v| j�KuW3L�{���h
�<m�yD'Uj���۾�:���7�h �e�)��^ ;����#V��TK}�_$E�M3@}�մ8)4>��q;�2u�=t����Wq�ʆV� y��ΰ�9V��s���no��CIt�#R�<�Z��iW%����.���Kj�Q1(�,����U5����G���+r�Q�t��N�7��Z�ju���o�WK@ڭ7��6�ǽ�L�
ں@h}��,V��c�����4����Z�fӦL�x�;��]�v�4�f�󮔻����]'7�\(\�l6Ղ�'k^}w����|�`��b����c[�;I����O��˫:4���)�]�f�v�/i�.�gI�!<p;]}}���G5
����dtը�Usw��ヘ�U5�ވP����GF�룮�뮺���^:뮺�:�N�뮽�뮺�뮺�ۮ����뮺��G]u�]u�]tu�]u�]u��:뮺뮿u㮺뮾:뮽�:뮺�㮺���뮺뮺�뮺믎��n���]u��~��~��~�_��㮺�:뮺�뮺믏����8뮼z::::::2RX6�����X�y�Xf��N���U���u���.nP�gE��:�n��{\�&�*�fg*�M��}w��*V�4���)2ƛbep��J�Wʶ���݌q�X=��U�1���h��h4:F摗כ�j�j%��s@�rNtO*��l^ss6ew;R>�IHq�mu(�W>ʡ2.s��'J	�v�ob�Q�#�O����R+����3�X�rK�e��W*{2�M>$c{r�ܵ)�[�9�ݧ�)�T�7jK]ʛ��͵@;��������f2_v�X���w�r�R§>SԎN
�%�Ռ��a������R5[n����2�P&��x��sӺ�1����77�� �!�t�'0g���sYpf��B6:�ܚ�P"8Of��˙o^��(m뫓��=�R�Y�
�V�єl��
sE@X��7�.�[W̔ �w�Z���u�m35u˶r�N����X6(��6��j#���L��v���/����vA�]b�.��\3/D[�[Qws��S�/&ٝ�ji
���yp/���jvl�|5�x��b�������}6��7�5��!6.mS�YT�dtL(������_���뮺뮿]g]u�]u�㮼u�]u�\u�^�u�]u��]u����]u�\u�^:뮺��]g]u�]u�룮��u�u�_����뮺㮺��뮺뮸뮽���]u�]u��뮺뮸뮽:뮽:����|~�_�ק뮺�::��]x�뮾>=�_~=�뮵��{���w���h,�]�Kv3�c1oWΘ+g�d
����Eܲ��t�ƹ��]�v�fX�+c�ie�R����Ǝ�	*$Jh�W��Y��C�Z���U�
�������uY����a�n��-K����r��+H8��k�>y)Գ�b��D]Ҩ�d�aD�͡{�L�r�!�p��7��B�Nn@�t9��Z�e�nc=�ݖ���B�`��#ٽKcw�wv4��W��y���&��֐��[��@�f��;����֋L+]�;���'W:��{�x�rÏ7h>���ʦ݃ʉ��mmf�:�ƈ�c}���D<�.�j��ꡋ���5O4��:�Yٛip�D2�I�LC�������M^G�Ŗ�
��	Ծf�bSE�=�vX��t��7Ϧ�SݽuB���nn�,���5o2��H"Pֱ�����~��صZ)��`�}h*8^f���;����7�2����fB��B��k�r+�@���Qhg	w�u��:��Zȼ�r�M u�8�2�*�u-���OG��rqwfXM�v�r�u�o!3F�lŪ�����5J�ҁ�	o�)�<�<|q��u��뮺��뮺뮺�tu�]u�]u�G]u�]u�㮼u�]u�\u�^�u��]u��]u׷]u�_u׎�뮺���]x뮺뮿u�]u�_���Ӯ�ۮ�뮺�:뮽:뮺뎎�뮺��]x뮺�ۯ������~�_�n�뮾::뮺�:���������n��ۮ�:뮹�o̯��+;�7^�I����0�՛A%^��\1��"�do�}�bKe�-L�׎�%�y'V���b��
�2�V�n��oZ����%v��%ޚX�1�ߤ�bmq�x��,����~.E���
�,�B�I%r�sF�z�x{�3fgn�
G-m�e�+�Z۹�V��r�<�a� ���Y�{i��9�ݣI����#b�	�FW0�L��M�*�.�;\�� ���t����OAR�.���z5���t�3j�\�R '�;he�D�0��"q���:�Ԗ���fn,J{�����U��5�*��%��q:�H��<}z��0�]�����]�T+C���p�9E�[�6w���h�RV��0���ub��q��3*�V��4�B�[5����dK� #���M[]�f[;RBSү�����ڳ��Rq����m���&�:Y�������\�oB˦�0{n�}�(&ھt�4*�6��ZY���]2f(���gp��I����m�
�\2nBmR�/����ܹE�_W2i<$��Q���߽d}\��n1�+`����^ԕ�Ҕ��ۮ������T�=�Eƈ���[onɽ6Q��3|��8�f+L�$��.ww
u;��+�p���Y��[P�۰�`�d"%����@�T��D�7F�;̳�/�	�+h�*i�}VV������b���E��1�KAg`�,ݚe�'D��5zE�P
a�.�����:/$��Bns��7^�FSt�*���d=�e�K63HXw�tN� �Ò��Z/�b��}O��;,���\��uz�Z����(^=KYw�:�}�V1�q`��Os2��L�4B�r�J�O�0�0^����t���3�5ur���=��wob�GTT3gf��Cve��I.�,�W|��3S�H__tipj��y���:�ڼcy�i���J��6�9��H���ʼ��FF���-�ܚeN'��m;����ޙut�P�ܛ�5o7bF6ڝ�zЭ�\i�.���ۃgWo�������a�y��$G�#6/�_V|�ɗBn󎷓�d�W�v%xՂ+�ϥhhiCd�"�#;ٷ:�S�BAn^�֍:��la��c�aC�(��)#��oe���.���ʚr���<7{�ۙB��|���8]i�$�t�]��in���hr��{\�N��,�edoy�f���f��[Q%��UvP']9�-<��*�ꕛnܬ��]�԰ʌ�0���f��v'T&�V<�m0�6n�(Kq.i:X0M�����T��$�}x,6�;g���@V��v�W��Ԗ]q�@�3wvne�v�}xYj�ͧ$�Ä�' ���M�)53�7ʑ�����d����/����������v��K�c�F'n��'ܞH:uRU�A���L���C��C���d9Y��p���>0鷌�oi��=���t���z��f��-���;���lᭁ�e�+�����JPbh��K�}W[gX.�k��I�n5��ہ-�,����|+l!*��u�>˧r��R�Gw}���e&M���t��ij㽳J����#��8��/m̔v�^qC]��e.�ɻ�k�r���ܝN���j �)�si�V�SE��O)聒m�르��XYQv+�V^Κ��a`�#w�햋4�յ@%Y���\;&:�X���aޜb�d��i��]C#/�d���uPm%���0��$��7\^u��tp����2���
����+��M�QS�a������ch��i����n�e[�+���7�+Ы1!wl�0�k�+�=9�w:j��8����̀��y��άt��j�;
�.��,ԝ�V���xeZԶ�|,N�/:`a����P��5Mrfkݥ܄��F����aI�
�ж�︲�Ҁc�﬌���T�MX�L�l�qWjRՌc�uZ�.k���艭��+��êL����;�(m	����v���BdG���+6�.�R��J`p�(��o%b�za94Tk��.�pܦ��)(9e�{$�2����yw���:�_`V��i8� �o�w�v��gu.��f]s��dY6Y�Q�a�n�YR��c�,�����i_e�Ș��"�[��zUb�]�h8^i`auadVvJA���jYv�Sl��ĵ���{�v\���7ͬ��sk��_d �圩�W}�9.�s.�2*+-���v�:P�E��"C�t��w�K@�x���ڄ/�u�'Ai�N��l���7�c���t�#h"�J�k*�i"��DGd����*�Tgw3[����
"
��������߻�;�������g����PRY�tdg�Ze���S)E	�w��:ff5+�����\�cW[��v�ے&J	K�\�3�I'�*:�\�tHT����L2�v+u��Z�U�vAQ��dk�8��AQ���T��1��Ź�l�ȑ�v"��ݝ�Z9f9J�8����AIX�̻U�u��)ᗛ��a�	�nu��w|�BnF�l-|�̢V��f��=�:;�F]]�um��q��YB&��-)�"� n㛱���k&�ˎ����p궨M�#7B�E@��7k�G��u���SzZ��m�!���&����uAۢ�z��h�q�f���I��q�Q�,u�y��0�eh� `��ͻo��@�ɘ�ժ䑷���0`� 룴^s��j^�f��42�!�]!�+M��y+9�R����L�r�$=��^�#UE�+ˡ��I�,`#+Se�=�(�]Kk��i}y�r���!�S&vJqfI�͔2�ԛu�|��ڻ�*�t=(RYW�r�}D%Rڛ��&�wq-���* \r�a�Ǩ�"�ȖU��:ܖZ��r��8��P%��6\��W%��6����Yslu۝7��A�V��
��Y��/�l�����\vV�UO��nV#^�4�H�i2�2�r�ӠZ�&P���U��U���I���c�](��)�����b�n��e�Mңsn��\ѹ����]�]�3lUGq�n��v�+����sK��n�N�J�'�eҕQ�ѯ"�	Zà�! ġ@̻��FM%Qy�Z�E ��;I�{!���)��-3Hr\ܥ�z"�QaYX�����j¤mγ#R���Si+Ƿ���������u�g��~��h>�r��+!���W�bQ���@�������Q�(AaH4EH�SB4%E*�5By!ɤ��J���XHH
L�9;�͛5����ϯ��C�����	�8Ad ����Ĺd�h��d�P*,��B0�n+�q.e+�D��h�
�)"�d�� �&'���K�E Q�+ 遛��Yqv�R�(���M�sRJ��k"8�6�q[���"c��^��O�^�����G�_Y���*�����˕(Z[-�7\��h[� ���R�DJ���*�̸�d�
(�Q)�r����s)�qH̛>�M�6l��=�ϣI�|�~\^������.���k0u�u��5�V�����2�q�((�#,�����ۏ���믬�g��{��a�VR���C�Z[q��l5�*�D�Mlc2l�}96lٳ��<�O�f�z�Cܣ�m��b��[N�������"n_m5�Srb�6��d��3�Y�6�m*��"�UVѭy�1-J�(R��b�E�r���T�T1�K}̇6�Z��q��*j�9C���1\F��&
�EV�SLj����,s�1YZ�l�gM�XP�A��"��n��ai���*�{���X�z�nK�;آ�C�x���3�J���`Yo���]�r�WHYi�*f\���p�*�
�iB(SI��]�7(�f��V��o}��$A�f�>!݆A$���O����5V�j+edYf���\y-ь��RXյ܍��c�.�����Uޙ؈w������./�%�Ծ���\����Uϳ0m�sN'�[Y�9q5²GN}����,�u~9H�F�z_?r�H�9I��Vײ�{�M�x�2$)����Y�g��jm�/8�χG��{��_S���k�Z|>w�T����B�:Ƽ x�W�D����=�g���{��:�����0�w�;�i�{�x@/�[��wY�W�{L�=��7O7�3�%�ci��O��f���O����J�Rz�v�r��g�Ͻ⤕^�|�QN��-�[�,�)��__i(��)��֤O_��ǨԟNȳ�r���a�[�m���}�5�^ҵ�����=�건���9�Ws��;#����{���BQW���
\��U�}�[��h��O_[��$Ò+��+�Y�+wN�f��[���I�6��>F�록�{�|��n���^�2hW�~1a��Q.ѝ¡=oQ!UwQ�Hwv	 ������۹�0�d\�^d��)� H��G����{���z��ނ���D΢<f@{}7>k-CW��2.��[��^�ޓQ��MN!Q1��b��
`�\+����t(?z��.v��p�s��^�>[�US)�zF�5����$�P,iN�k��|���bu=zg�ʽ�Iڪ]z�0pW�s�T���j�Osr�+Mr�\r>��R>>*]�=Y�vs�ϸH��:�L�~�/��TOVC��h���J] ����� ��ل^����s:o���V�y�NQ�����faH�^F���)�K��=
+�{�*���EmO��ս{��ǜx歺�����Wn����H�4
���;��iح�k��E*��?�y���y�ٱ��B���nw]���h�#ԇ t6�DUs���n�=�w�|j�ɞ���9�[�*!��c��w��<(b�Ļ���^5�k����C.n_q����)rSh�ٶ��w����u��z{ſ?zM;e�Î7��i�R����>Y��V��T�b.h[��y�L�:�uv�=eWHh*���ې"*��J��}��x�=�y��9o[�غ@�����C�o�����{�S$��9�W��ٷY����z�/,j�X��e��|��ӽ�Ѹ`�w�m�	g���`��^�Q�9�%��,/��ڦ}�������^M��I�Uݩ�`�N.>�-M�Z��j��o��{��I�^��d&׻>������>7�i@�ЦV�R ��z��ߢ�wr��<�Q����Eh�TODg�l�צ������̖��?(���g����8�7���hg<8n���	�lVwb���t-y������R��os���*s�[�i�\��b�`J�
z�ֻ�ky�u��i���'���+����u?n�w�A�쓻�X_��!�o���"�A9�=�]�T����	�b:�t�>�PPǅ�w=��#|��s��w7UtMUN�a4d�&w[cA{Z��հOD�V���}*t�u�m���{�o����|����e5���F	Z�y�(�N��n����xw�n9��q�ӧ�*��0����n�Q��]��&*�WI�	�lgڣ]7���u�ԕ"������{�z3�\:�����<P Q��"R��w����3;�E���Н�U:^�N���[yoϱ��`�u�Q��Y�D�aO{/g3�'�S�yoR6��r��(Y��8��!Ȯ���"����T��d:��{�ˬ���r�e��H*zN�ޣ�-���9�^���V�<��B��,�V}=�_��������Rh��{�)��c�7
�m��}��;�����'�+W;M�MGdbA��(��$A����^��e����i��m��~�>���]x�T��W��yAeJ���矷� �ylϾ�>�3j�w�S�
���t������x�黽�׺/�����(�Ԥ\�t;��aFHѪ��F&�1�o��i��<���*׻�D|���ӵ��cݒ���Bn?o]9�Hv���-��2�
߻��'�I�]uG��g/���~�Ŗ>8�O��X��l��P:/��`#je�7�I����X�b�˦t��[��0��]C�'��uI��%q����W�;�=�ݺA;o\��C*S�q^]�t�NZA�qF��JD6іٲ/�w&�ηsH�H��`�o���{���I�(D_�1�s�2E���~ܾڡk}="S�r�}�|���7�s���y+��G`jg�'��J���j�e��;��L��gez�r�ϘS\��<�����7ݮ�>~�mw�gMͼvEݷ6���l�&E;��H$�xpq����I��ֻ�ѕ��Md����k�����~��B��0�}�z��7I�jOa����|1�r9�u�^�o��V�c�ٙ�{����p�edo`��K����iC�s�w����w�AA�*�J{5ɰUF��Q��u������z���7+��u%�'���U���U��e9�Hh��}g(ty����ۛ���{��{�z��8SHjd��D��kLӾ�0��7ٗ��۴�,�a��|�]�|=K/!K8t����띒���t��|�x�;�)���~	?����.�C�~�=|����Ҩ���ULֵ��}#��P���vg'�vwK��	��]_W��H�0��^YM�|�p[�	ҹ�}΋��2��5\������c]N��H7�:�Ө��t�)k3{����}���E.	���Dh"Xy�k�ݟ���w����ݻ^���c��".��jt����zM�-���t���,������6���~{h�3�������E��=�Mzj̷�|��5�}�=@�4+<y��M�puմd�,|� ��;>��'���,����35�p���p*�����p3�x���5��cn�>��"d�s;j|L��U���UCx;ݯo������H{P�dmI��t4�0�_���W)w+��b�{&��"�n�xv���y<��,�U<��� 5�Yxif��<�{{��y�&������[�U����y��x�̜�y�d0=��zq�N���܊m�2�h���N����M�U�К�F��N��2/��vc��ߙ'�Ă� $���]�ޟ<}�����4JA����|�v^�6�2�}Ɣ��&���)U���
��n^ɝCB���
�N�x�7�����Ƽ�c</�m����5q:o�j�	�J�_J��`����b��w��#@���>=��޽
*�8�ny�ۖ�q�,� �@C{�;y��z'÷ŏu$�I��)�;�UM,�A ����m����m�tͼy�0�Y@�����ޒ0�z"G�j��9; ���*���ھ����9Ǳ��yY���ڡLJ��]�w�U�G@Ϯv*�/���d��%{ۛ�~�ܮ���Ga�^���ɸ�_ofD��������D׶�{{o���I��}s��*xNN�d��ϫ�]�]�<k}�ϑ�b��w��c�^Z��ܛ� 1>��..�=y��.�y�p9�����S������s�r�ٝ��#.$6C,���]�r�po��W��nh�Yد���Hƾ�C�ÑC0d����v���=c%��f(=Z�1�=~(xT��UWY��������4�1e��@�w�&���y�B�Og=���[���7%b�y��vUv.�L�Ao�<��K��ܝ{l�S7��Yb�ː:x+sr���C<�gzE�C�y����3}��UD��r��Z��ދ�>���5��:��:য��Qh-�W)�Zs��Wv�uj��������e��9vlt�t�$x�<T���}�]��.����îs�6
�X�Nv����ߤV�y!y��Obn?|��>����1� �>����0��\p�l����߼��,2ZɡY���뢋Om�l��b#�Ǵ:���]�c������x)��O�8൛ʕV�r���㣍#^��$��0�$�N�r��q}�T@��4MM;�Ӏ�F��[�%��dH�9�G����P��W^_��8���#�#�Ã�uH|
�*E��T\���f��_a%��d��䧴^�mw�k ��uq擨��[��F����{����p n���.���W>����q�a'e��%^���Tzߦ�a5�g�ݴ.t����.����{�o����������c���N�ym g���ݱ�4n}~A��rt�t�G~a=>��s��(i)���n,I��N�9�J������|�6���b<}��go{z5²b��p�N��rB�ːQ@USo!��[�.���IN��)u�7�����g��s���7�K����j��3,��c�,��_^�s:Ii�ye̆��CF��HU����)#9y�wr���o3wN�"�B$" �m6���&�]�p���`��݅��4h�wW_����ג������pB֫Q�ǻ��Ә����[� Z�̍���wW��ؠ'�*���O��>���w-�]o<;�aE����M��_L�i�����۞��Ӛ'Y�@bo��;���z�cc8��&��;�zoj��]nuҎ
sƲ�Y��8s-?{��vG�����Î{h��;�W(�Haz��k)��U�/f`�y=~�8׶�w})�����X���+�����p��r�?go���^�^���4RT
�k�:p��˷��z?&}4x�{z���R}�VP��3��yԬ��}����A_�Gg8:�.�s�˂���\p����h#- uo�e�_���gC�U�Ѱ=Q~ѿ����]<��?y���I�^s��_!^}�{2*����*����Eg�Z�b�^=D��.U�|�("4����T�g���u�Y���n����P3�F
��Y�Hn�r�-�h>��
�k�����Q�rV��	/U���-�-�E#wK��7�lS)��Q7�Ídl�1˖mt/e�yi)��@�`�l���'Yp⪎�
s��{��ը�$v��M��wA���}��$�]��`o��*�|��� �/'�9���1}(͚Vvq���&O[�wV�軛�������/B��>�=\̇�6� �S�����5��� ��^&�@n���&�����<�~����wH�e�۴,���0b�	�y^�3���vo�n�����f��]"]��ٗ�I����U�ʽ��ޥ�s�^�gY�t0H x�9���3�ސ	嬶�m���.A�c���|b�eyW�|���r�>�M/$���x�Q拏C�e�"v)����Wr�ǉ�}ṺI=���O^OoO,�"��H�W��4��ėC����.Şq�{7������v��e�Q�i%�\�WL>�Ck`��>�p�'w��xx��Q���3�Q���M�r��]kte/�Nܤ�t�FfLx��:[0>��w����%G,TB+k��#��f��u�Pl=��M���ZQ˺�TFU�-j.�p^%�_��B��Q<���[8H���.4���T��$��uAԙD|& ƭTꗩ�:����f]�U3H<B��{�|w�6PU���k�����x4s�֎�n�a,��;Ww>�;9q��u��nEs��y�s��)泔�t��pU�ǻ����UߟZgﰎ�X��ϑ�ip�������h�'L�Iar�L�xe�I�&��{��i79�PEe��j�Op)��/VG��b�Y}���M�����ڻ�'E����ܜ����\�u�g�;E
�ʻ��	B:�oe��&WL�gop�ܗ��`^�C��gD� Q�L�6���?��<n��.wh�vy���ۿ\;sÖM��,x��V�բq��PtV2u����ݦᏠ��{�X�EٓR���1veTJ�A��t�`��-]�gtn����J���Fm-���ǅJ'�t�W|�:5v���/;TO�l=��+�����p\�n�X�+vS���8�-�4)��Y�W�6�uw��W�H�<j����b{��4\ �k�m'Kv�f�d%�A��Z��Ln4Ŕ���z��%PL�a6�a+�g���;��d��W�v+j��e�d#�
f�\ �%|l��OX���BT���C2'�މ�b���Yʙuz��4�ٖ�a5//T� �4��w����)I�w�w���w���RKm�����Ԯ����$j�w�|��K1?�'���:󺳬�Uھ�f7Z˰R�ن�3(�q��EsC� �w�s]�w��'����/y��l7�{�U��ם�u������)Ȟ�܏7��̎����zHz�R�V�j�Zٽ��w�Z�[
�"<K���9���Z"��)k���Co��M�Cu=E�PfMɪ7������I���{��W��,�
XW���â8S���T�V�2��b��X�e#��t�v.��Z�6�G���.��3��pX�N��dU)�ꢵ
vT	�Z�˲�*�jӲ�\�e�4�;�9rd�α�/��l'��j[�FBr���Z��[���[�e�]")n	+�1��(�&Rj����E�H9,{B�����b2,����|􎽛q�G�9Y�VJ�uRwe�C��mڶb��:vWL2��M���T�gw�C��U^Ue�]וއ�d�@F��c� �lĴ=�.5������ʨQ_����\����Y���ɳf͟Oc>�O�f�y��TL�~ڸ�㌕�nW���Z��H�ye���*ê5H�(�YTK1�e|}||{{{{p~���3��?MOc�s�J��cR�*�[G2��1D�`�M�ш1�d���ٳfω��}>�Y�#=��,����*��K�\E'h`�U��N�"���78�e�:���6l��=�Oc>�d���ט�H|2q)K+�\>.Aq��l�p���r5�̫A[eE�c2rl�rlٳg��{=�g�#��(��_����˹+
YJ�*4����6��E󛇏0���-�1D���Y��u996l��=�Oe���3Ͼy�K�6��AE9K�{
�%mm�k�I����H�C�{J&���cJJ�5+�YX)@X*x3pٕF��Q��kT�.���\���^4GVإ-u��x�SX��2��Ƞ,��6��u�G�F(�E�Т)��V��W�c@�Q�	AF�OS/3��oe�W�+y՗�>�=���K��ڕ�kO:�9u�P���1�IWn;�C+�wI^��}�0��x�0��֎����"��b�rǗ���q��ޡ�w�������f�3��k�=A���Y���R������(���E�i�r�}�� �1�3$Fz�Á�t(�1`N����{^���x������彃� 8��/�O�(9R�`�n����E��p�= 	N�voj(Ն�@�#r�2��Y��2ݹ1����KBu*�
P���D9B'cnl&@���0�0�\,�r�Qlfޣ��5���η$2��@r�1�A�|6�(��b®Kx?�\Om��?s؇����r@�S�r�W�\��e2������������ֳ���$��܁-�9exV(���^[P����N�K\���LE�K�W���8�*��9���LQ�1pPb��~/�ؿL�^��uW�N����?u O[s�ʨ�nP���<��y�^�3�1l�&iY��|��$f�Q��@_� @�M嶧��kQY ����B�7����_�~�y�4=L���M-�*�S�X�K�|���C���W�%8��zj�w��~����ؒ��6�5Q<���˟BVP�W@�4cxO� \:��A�F9�ΐW�̀r|=��ʅ�[oob���J�h��3t�)L�����6_L�����uXS�|+3�{��Bs�Y|�{W��i��e�nc���ꔝ���#;4/�\h�x���u�v:ボ����qo_V㖪l�������	(,3�	�<'��E;��>oYﾁk�w����j�0�/��ょ�(�>L�BP��|C1���	n���r~��6�PY�׼6���_�|D�F�=�Ѕ�\�1X�p@dd��`OsLB9��x~���q~� {~����
*�l�� �D
�?A��NA>Ǥ�Y�1>���W����($�9�`q,�����3^�b}�\���!�1����YK�n(���#cɼ'۱��`��[L�wf��咨i� SW��i�7�%w�t��&^cyvD�r���;�^��O��P���ruI���CH}s�x�<0= >�8��7��ˠ]�i�K�ה"��0��T�ӆӸ�ʀ� N 3�/��&ѨV@���|쁔Pc��4X����״�NG�������F�0�|T.Xy���;0Vb;�(��o4��\_+5���']r����}��&=�>�۽�VbO�_(=�-<�&/�x���1dQ����8�����Aע��^�K�� ;���@��P�%��6a��]�r�i�� z�h7*����[�U���A`&X@�U� �W�0=�(
<@��;��WX�V�k��uƷ��Q��l�9��؛RT;�����7j��'0@1Ƕn�^S׭l�P�L�ڼo�:m{:�|�f��M+�"���3$>,3KT�>l�c��I��$�@0�2%�3�F��H�v7��JZ�%�Uq�sd��*#��ͬY�#ޏzֹ���4.��i�WY�7����p��˖m����]6��q�h�m���\��tsM���Yc+,ee���n����y���
%��0���!+�DV����q@�'\�0.f�����_\��n�s�mؙ�:�ݚ�}�K*�7�p�;u4ml��k��0���g���PM q魀�i����'-��M�(�=��KP�@�������=���;�{XCHC��l�9�ϟAc4���O��r���v~�����'�$��$��:�p:`!�>'w�A�c썽�1U�+��B Ҵ�����������G��F��{��v5K�k�IN���0�L�2`i��+_�ӀZ���{(�/�K�G���60����?~���%@?x�����609��L�7�2K{�Q��`4���`i�=��b� bH��LM-��^q-kk��������)��x	$��X�w��@��~�Q�H �P3�x���`ik(*��� L�%b�L�Z�3Z9���>� �=r��@fq���(���g����a����m;Vr���(�u�:�-qnj���O���߹�?�������/A��
D�&�ǐ?=i{�98��91=��n)��EM-iN��y	�8�y@'�cL�DƗ̉���[�Q��	�
�w�y�����ߓX�LWEM�f]�F���+EV��M'~yok��a��R�a�r4n�f�v�y6@&���E��W-���}�:�K(��Ⱥb�f_ #�C6���7�_e���;f,� .?s����ߥ��L�#,�1��`���w���ݟg���@\zm0+��q���<@��(U�ŏ.�O�}w8�g�!F'��N�R��e��sz��}�����	o�Qt$����tǧzh�.k���L�����M:ƽ<���F������{̯#wc[ö�C���><t�!<�X7��
�T7���v.&�^�՚-�k���x��܋35Y&�ڢ8��1>#���G�sƟ:S�nh���!t����c����G�[s���mH�ٔ���<�ūhK\��M#|ťDS]�2r��ٻ�%?c�[�غ�fְ�,�j�!�[�jyP�)	Q�!�r�1�qx�v^��H7�|������!�34R�Ih����Ŀ�Ys��S*�YX¹B��H����7�؈	����j�q-���Yp#r���+��W���ݾ�H0�a
��Wӭi�A�S���ʭjM̙���c-�������B��33�PU��\��\�����������g�}�Cw'y3t6��w��ii��v���Ŷ��������i�k��q���M���oͭȀ�:ͯ�p�؆}z�le]�>�����q�U�zDS��w�+��� �L�s�^��9$y��NNu vW	x+�aX�d��%u6b�t��K�T��n�/z�݈ըQ)�ݹ|m�XX�L����������$bF$c(��v��>�����=Ҭ����\�P+A��%��W�U����KO,wƹ�q}I��E9ъ���/U�9WbƊP�Ʃ���A'pk	�$w��U*yn��-Y��*&��讴�1�	;���m���[o?��8����s� *G�n!�������8���r���:IU3c����O�S��3�@X#���,��o�/zd��vg���RX5%�%O���kاF���9A�a��~Ռx	>�TeF��<��8XK�O���˗6��R�YR��<U0�a��I}l��p��(l��ϟ������{2わT���Z}������������g7����/�)x�p���7�&��fa˳�^Lk�2|���B��gL�[Y[���U�OCד0M�����@l�/�]��<Ģ��� �Hx���E�Z��������f���l�8E���uo���u��΃�@
9��fBeZ���(�m��CXZ��*�H�@t:����UI`G�w��~]�j��� �:X!L����-�~>�*��x=�!�Ez�Uz~,/8�
����я�an���#����w�Kчr�uj�4�G���)���I���	s*�Q������!�@% 1���ݛ�4����W˄�#+(��P*��!N��ooc&�d���ɼ�<C6S��� ��o>��y1#�e��"W�_�����'�>(V�өѝ@�I3�Z�_���Hd{�M��|�W�ޯ�%h>���ʜ�lO+y�/d=�21H�w!�>30���=;�]}��黱H���x�8����t"W�pY�ɛs�@�pd������Q?��|P�}p͒.)�D�4���j�|�o���5��-�~�|����mO4��A28r�ͷ�L���+!�^���r����"a��T�n��iSе�D���$���/v�O�P~��DV��"���3&-���d)�5�5zY��<�.s�j;����Q�ѭw�gy�Lk��r��5bC`-+�R}�&�M�k(}�^��~'Э�aQ,��o������ C�����#����
���9��kl*+v��+�-aK����Jo�@W�^�v-~��0���Y �	��<���if�`�;���n��@�Q������+��1��~���2{Xu��c�z.X_-X�F���Gj��ϧ�H��O��+��)���a [�z��	 <�b�6zo�H�󞅰�j|e=����4��Kwט�N:���Q���Ɲ�+s]�Z����w������a���9����jh;"`�,c	�r�+�[<�'�J�᳆=���ݖ��p�I�7�c�.�'UY/�1v媖:k;_H#J�C��˔J��i��	�%�
�~J�%�l9{H��2���d����|+H]+~�4�vy%$/�△��<Z��S������ߖ��
}������O;��?c�睚t9fFX=4׶.:`���!b���n��8,[��e���G�T�~�c��[X|Q����XF@��x����C�X�����-����o{;jM.ɴ-z#[�n	�ve��>פl�rjׁE�^X��lZ��V��"�$������Q0eٽ�J
2���gf
�Q+������I�t;k�Ia^*�)������0���7�O.��qK�jM�;�׵=�wԮ���L�1m~�tX���@¤ثH��	��Z��*	���&B͋�f|�]��b����iwSߖ0~��#px���~�%��RLe4�Փ�r�F:�tf5:he���}^V�G�Jk&+�D5m0��R�p���3:�D􄽅�]�|�w�Zl��738�=�8���vJj������u
0#�{��
��L�*�:�|���m��y�Z�."j�={]�VR�l�I� c
�ڙni：�36=�N^��_.��_�cF�V�Fb�F���Z�������S�pA��(lf�2�OU����"ߧ�� ��kHg��#�-�D�-"}
�;]�kᝃ^��%0m���*tf<�>Uc:r)�����}&����(�����7mؚ7��a�W�4�Ԅ � �/�A&��~��������gM�Q!�ɳ�X�a>7�Qk;�h���yn�����҅�����ݼg����g_�8�KވWB*�~g�foө�Y=l����D���ѵ���d�y�l^�}���i������C���MC<�=8�d'�w������!Y�Ⱥ}h� �r�:Y�xC%��柆�=��3�:��%y!��k�J���a|�e�'y��bK�
����6C3'�=�5`ѰGr�״[l�P�������,_;)��~���?E�����Uz(��%άcÍ��ߚ�qv�J����H4�;���y�~]�3?G��k{�B	3n�N�ޭ��J`���逤��#�dS^�����<�x`?p�0JF-d�g���Ќ ��T�Ŕ�"�X��um����Ɉ�} R�^��4[�A���(bC�ܠ�S���l�D�F3|~�a�t�M�0jp������ζ��G���'�M"Fu�h2��J��K�.�i����v܇h�t�M[�&�=s��r����\[)�Sz���W��p\��D<�ݙf�R�4@�|����"ȋ�w�^v��VSq��R��Z�v����GGΙ��s:��ǿjw���"E�v�{�U��"`�O���v�CTѮ�o)�K]��e=�HqƫK0�/�O�R��Nv��ye�[�w�μNv]K�K�z~#�!H�ei$ĖT��>I�a���bA�ipnhS-��ns�m��q��Qm�5�#6n(U˸i�Xtm^���4�li�-�R�+��ϡ���|�1:�ԧ�����[s�w��º�l=�q�^�8�uSXd%nk=���K�y��H�gB<2�Rw���?�[��>�w�$�}oⅥ� �(��v�r���M5�T2x!��k̴AQ��8V����O���"౯Z�>*N�s�%He�١̝���L�۾�D��_�R�/��/����x�+L���yr�o�I�Qm���'��k�r|�]?��������<��G��?;�>f����	�Ƃ�Y-����`  	i.��\r�ϑ�:Vh��TL��ݬy�������1ʑsV+ޞ23��\ -L�c�Pw.���SM#��&)��"�Mmz�uÿ*��=Z���Q&����1�gѦe����ώ�qk�YJ��XxȢ�:�����&�y��C��T18x���8Ŝ4]�C;����ֈ��K��Jx��%C��Ʒ��d;���- ly@�j��=t�J��oU�mo�VT1����hyp���ޝ�d�Z��L�r\G�{��v,�����`��%!m���FL��_���jZط�/�����=G�P���t\��)�Gt6��Dav�\��ܛ5 7-�Qwt�gV���bm���/'p�};���|�4n���R$Hče"A�$A f'<=�{��~u	��Wť���dq�Vr���~�v{���@�@]�X����:VgԘ�t�c>߽��"G��A1�w]/..pc}��pkH�
�Ho�*Nӣ$���\�Eb2$6;�#8�tR�c��M
xH�y痩���mȓʞD��6�r��ɧ�M$���(w�����)�Uy>�kn�?)���!�e߾[Ng�gt&���1�]��s�.����u.*������'�
T���~��l�����kJ����N0Ǖ���A�c݊)��=��2�G�J��'�,�ꂤT��I��f�q{	�q�L�P��%kWA��y��}�G�/|`��K'%�۰!�G��9��{OI��`t����K#��lzy�ݔՌj�h�c-j��n��75����Q���Nb4T@6^7e_�
>P�C���t����A2���to��xoT��^�}�;0\�DnzY��� DbO��)R�m���]/Ă�=��팘���͎3��{!�7�3�rֿ��V~_H��?B�ɸ�la ϖ4 � @���[��^c4�%����Y�܏oV���O)>��wG�V���e��sN�3����v.��I��]V��L�dE%���X7�l��(�������t���B,���}��9�z�Αz����� �'���=�`�ݺ,��Y�u2U<жC��Ee��i�U�� �&��}A�pt�3�K��M���2e��n���@���r��2_*Xz�]q �쮙S.�Y,1}�����d����<�p��6�Twe�4ZAJ�F�m���R�<Ԓ3���+��:��Y@q��!s��2��d�|�{.!AZ��\"��D�u|�NG-ͥ�F��DF���{�5|[��x��O�9�VF;���:c�r��2C^���C�W}����U�1}
1�<ZZ�^ג[bvQ;�(��T�����䪞�)h{2�勖#",��v�]��t·��4o�������i�w����TeT1J��]�8:(��§:���3ifB*_uR���Wp0�x���u[��
<czip�+L�3;X#F�:"�����ܕ�Z�jX]u��MGC�P<:���'�M���I3��E�#�k5ӝ�ff�͕��,��2��x�a��ksz�oKi��¯��)�<�vfEڻ��[�-6�����&I��Vy�h����^Z����@��b�ӳ-Ŋ�Hi
�%
!ks�Ý<h��u�V�md�-H#�z���[DS�.3���: F��Ei}�Q��G�+��F���������:�>U���b����B���*k!̻7�K��U8���!k�J����@ș�.�T�����Ze7J�[�"�n�7�Yr������˩-QNK�ܖ	��;��u��2�O�������;@��-��ĳ��q�%���k+�_U2�e_����:��R��|�e��s�8�!�x���}h�ŇT�芠i�P�`EK�C��lڰ攺3���OqS�hvRWfW-��Wa��M��Av�t��s��I��ފ�B�ӿU�Ǐ}S.�ʎF�K��������r��ѹa������[�]�S��cv�ʂgPb�tD?L��F��c\�״N��;�)X�\9���7O�e�P[]R�pR���%��/d�)kbAу6�o]�K9�&>6\ѨD��yԔ�Y	�e&.��9vr��Y	l�q���❎�/b�KH.ze���g��s|/�+Ѫ�;�[�ZH�� I�Mӷ���V-�ou���2��[�v�XX6�{q����Zz�ۛ"�{��^��-|�-����(��z��Kɴ�rt.b�me�+qpٚd�&���S���e"5��7�b[����⊴�=�Rgj஭�rw��-ᕐc��\��T:m,m��O*�-�C��#X�4:�����nZ��h�f㽊����꡽�u�O����������O��iU��.l��<�Ɲ�bЅA�R��}>��չ4�U*(טt�
�)�D�mAn*	'�)��5*4�F)ڪ)�t]|��h��A�ѬI��5@�M0h�E_շ	�B�TQ��+�Q2��U��GMU���itͦ��\�7)�1.u��1`����EJ����W�����!A�U�0b��"]z�DB�x[�q:�7��YbG�%��n-*1�}lS^�ہ�b��%�V�Ш��W���fM�O�'&͛='�����}���W䪉mK����
;j���ElJZ���QYiS�:�2l�}:��6l�Og��Y�g�}K�ɓ)�VE3)1m�ڂ���?!���Z�+�IEEƶ�a=�������"jg��O������G���Y�g�Z_��5�.-�媨�Z�Ҷ���eV'HJ�G)q��ԍ���Y�����u998�]}x�gOY�����y�1����VU������|��;�j���<z{}~8���������x�;��
ʖ��
�jb
w.�,A���.Z#eoe��(���e�O�S�ӏ��������x�;�y<����BQ�KV�[ �/���5��)���Uq�����b���8`ui�����pQb���Ud�-j(w�bJ�Z�[C�LN�F��bTplrԪ�f���m�J�ۖ��b(�j(+��n<K����[B(���]J����P�V3[5
�@'�$P��!qh0TZKV��͝/j�]�Y�Lι.�h�X��S�ҶC*c���b����%|���+ͮ٘��.[��Ԗ��e3)��W-s��dH�	:���+
D ���I9�v��χ��{�^vI�E�.|!� �4���ֵ��� �͙����R���/�s��#XC[�t;6��X65O�0YC��%d�4�r���Y�Cg�6+�K�L�6I ����X��ʣ�S��Q��0��I!{��t�����\>d���H�����ڛ]hY��飥-�T
��~w���qM�Y%�2���\!�l90��)D L,1qRk�I;�YZ�^a��q!q���x�|������I'�.����X�+�{	� f�i"�x鴧Ѯ�"YҀLt�2����(�t���f���U����}Wd��>���g�_|����K�#�c�髕��s����A��cD ��I�X�YIL�qml��3h-���_�=������(e����D
�B$�Wƍ���2A^_z$u���]鶄�o�8�8MG��I�HkO�R�"��ޢ�}@S�ӳDw�m mp(���'�}r&w�C���Y�1$Y�IL�Г�����������Ѻ_l��O8��^~m��{vS�Ѻ<�?�:({G�e��m�_�ȼ{�)P����6n��Ӈ�/�x���1�݌�2��_t��IF�u|�|�K�� �c������v�*˹��x�%�e^�변��2U��\Si��{ΐk:�*畼���U��\��Q��0��h�( N�۾����>���D�����Z�x�^�w4L\�׷��P���MX�J&k1V���߼����o��Y�"�)HR<NB�aNA��=�*z�:佰�/�dy��-=yfe}ǚ��R,�
2����=�2D�~�vi��
��x��c-�=�ư�I�yd\�w��'��60�����B�c�XX�5������Ap��r�ksyu���%Jc�!��Sޟ�
Ort���L�.�j��%U8pӭ,��^u�u�փ�vu�\���gL�p�Z��A>��)����'k�XQ������gXv�6㗓M�*�,g;e����由Ęii�	m�c���n>]V�$g�KS��M�Q� ���^�osV:��gɨl�9\#�']�0`&�s)בIƸ�i�x���S12���r��� ��*�l����z�D��K<0�����i�È��{��G���QS�tj���E3* ����JC��w*����k�{W5x�<�����.�ί@��5�P%�=zTC0*D�Y��G�C }@{�Ct��:ٜ��>��W�=Z�i�5쑣w���"Ө��faMa�̼S�P<Kl�`y̓#k��鿼޲��3O��;��W�*68ɶf�����i�
��7�M�vff�?t�<��5���+�Y��(��\f-x��5J�C4����VF�d�v�1�`=�g{��ggN�F[Z6��C�I��^,,�H!$K([�%V`�YܠF�+]�)2b�1e<�t���G����0�3�͔��-�p����hkӊ��`��-�J� ��" "%��qIy=�C
�(� �f"" ﯻ�~��Ć��4�z.X;$�� ��]b�^>ˑ�i�h�Æ���&	����?+9�{[��v7��r_��L���s�ۧ��٨���.7��N7y��m�B$xm�3)y��_�"�G�[?r``C\_m6��F)"��b���6�4��h��`S���M�?{Wú���P��X���?�����0/�(ۣ�c ��Q2�K���v�J˴���~���<|���~'��َ����HTM�DSv�)0,�6*E��&���_L�O^��e�V0��g'"<�y�+��ӗ|�����hU�z��P��������u�T5O/N�w�954r�N/W�u^.q��B����?Z��a��:�N��r�c؃8��]>���P-��Wn�j��<��k�.~t��]'��A�����_�.������KiTyO���>�h$��j�'2�ZeG2эN5y��/~��謁���L�t��̉�4;x[;B^}��33)�Q�ƾ�{2Ӗ'p��p�<�;�TD�l�R%��87��:�n�2 �����m�E��J�	�� Л�!dy��j��ӭy����/���ւ�㿍۞��;��:�ÝOCy��N����ӺL���d��1�xN��8F��4����$�3(�"���[ٽ=�f� �+�l�gNS�<ɹ�\�6^9�����JHή�׹w�c����*�!�a�~d����!'�o��>�ޜ����_��4o�Pp����l��S$/'�=3�7"c�Z��u�>+�M���e�m9�1�K��'��E��"`cJ��W`qFm��pD���) \x"s�����}Jo��f��Cs�s�Q��2-�h� U�Kfb���������1Br>��N}Cdk\
8k�,&z=��KL��������ޔ�c�`���R�u���~a�rP�}��d\K+�n�F�܌@�c��>4~���������D`"���>�2�CT��Rfr��~�T׍tҜJ�y11�؈�M%k) s�]���K_�/�����L���@#���X�~�a�
�"w�ק�N�[{|�D�z���D��	b��`?���@*�(z�%�\�zF�=�m��+�@,�|��߾�As����v�Y�,���� zj��q������u�g��9���g�\��0L��E���Y����,c��_�!��KSf�7J�Z㸮>SˈΘjm�S����W]�Wtm��Ґ�VY�-����΍�����f���ь' ޞ״���s[�-���q.`���b��Ow)Ν��&��ls�%C�Z��D%�?1���;�N��qd�$`Q������Y�BY��n�v|L�(ى�)ו�o0;��jm�O�p��9��<�C�eY*�\wF��XS�;�,��+�S"I��KyR}�,R�l*��fL"5��dh6�	
j���۩n��a\��~E!�dBP���§�R�� |ˬ묖�?z�׋3���y.[I4�4��@	�x�R
n(�+�H�^엊��İ7�Mr�7�dǠ�%�-e�&��c�P S����i���u����F���6 z��e	��D�`0���{4�#X�`��D9!?HuO��:����
:N)�n�	�v@���WT�V�eG�{�Ђ�N�}��ja%�QM�~+Ow��z(L+nꕭ� 1���
y�H��_�u��J��~�z{���O���YcZ�6*d;hb�����q=��koLs;-]�D>2��+���9	яv|�5����m�i���[s�ά�Z��x΄�(�Ez�@�����˅`R�����q��Iů�M5�;��`��˃X�����_�E�3�룷Ă0D���`�񶒞��pi��X@��y�+���o�~��^�m{�� ���I}
o�<���Ly�Y�zC�"���Xz��3�^��{��̤�`-?Or:�jU0I�N�����N�/Je&f~�^B�G�6�_)�|�0��`3g�Ew�޺�Ɩ��"L����Y`�����ff����#P�_�į(�7<���B�o҉�x.'��*"$n�b��:��GZ�!۝Sv��Z/�u�ym�֛�v�}���*s���n�
n���s�"�x�4I�t�m�oǽzu����o6��z�K2���3��SA�Q�1h��.o���n��4[�G&-JN9c_1��+�#��'}7s�7389���5�
D$��9 !�d�UM��R�Ⓩ�\V=�^�X@f���NO����Q�ƚC�A`b���z�ϒSޛo^c�ơ�u�އN�/w���1�J���Xc�5�A>�u�9�L*�F�Z�I�n��v�MC3��^,���ߘI����3� )SJ�·�)L 9I����-L��r@�"��W��ý>��Y�t�`�0�r�A.�����N�1�����f6��{�H <K��-��{�7��΅�F�,";��Jc O���}�~�A��)�3,\w�;*����8����=,�>t��y�48�5��+{jR��$2�4x�t�8ل����.�����F�}�j/�����3}G���o�6P�|�i}�Ͱ� 	��������� C�v�0j���E6�2��5�N��
F ��:v���0�4�����#��,���q����SߥsY�3��Ԥ����mn�gX+�����i�J9q������P���P�������>�hS�`_�u��=�|כ~�Ou�y�Թ��鴁l��^ͮ"~������Dۏt�<ey�kL|Yg�y<b����m+�0�dM�!�Z� ���K�H��m�ѽ�C�;��n�݌�|p�oeά1;��SεB���ˏ�ӴǏv�'�=��A�;�2�M1��;!�O�ݔ�f��.�M��c/zr���?Ǽ x�� �`���Qa�^P)@Đd	���p���߳���d�f�K03�����M�����aT��
��(��Y��g�����5�}��ל�z	8Lb�?��Y�|nh�lcܽ�g)8W@fM����頄�:H���/^�˩v�F�Vzoӆm�ŕ0@CyaM���A��j��D\��p���9�=��W/i��z�9���B��XN)4\%���bc�P<�'�* ����[RA�e��D���]{��2�a>&�E�L9tO�7�V��xT-=�)���7���ӽ��\�Y
c����l��k��ڟ4����z�[���\�3׆��!5+�4�јL���28�S������>�=	�Y��u!xa�@M�� ��Ri�c�%fR�fW}6j� >w��>��#�5_Q4s^�����d|"��dZC�8f���=;��]Ս��wB�f����b�����WjL��^����k,koz��>�]����}{�M���P���9��_�ե���J��ʁu���F�O	�ޤ����L�?s'��(zı=Mb�U�>�Ҁѹ�x�
b�v��׌�*r}����M
���_~�٘��^W?_d��z��;+�t�@��gl�%�	�	��D&���
<�fJ骜���_*@��X*�HU�yQAZ>�O�>S��w�-	[��H]���ޣ�^v�s��J},��v7������`%�Q���+ꯏ���䄃��B 9	ܝ����u*Q��@tH��D@�`��ﶕ���A���i�+L��.%����RD�2.[:��{ă���G'��=s�G_i�>�#IX��{�E�[��V�?s�#�}���")��6�W�J�ޢ�Dm"���;<��4�"$UgW=�<q�-��0�"H�F8�<�7�#yH�ϰ�O�"�C���G��J8�H�D�QE�޷1@��S�12�ӕ�v�5!�-��S�8�P[[U���>�v5����	�:, �`@J9:��ˈS�i"�B�떖�6]L�f����+�XW�#�{�q����>�;�=��6q�u�,^��� 	-^��	&:&&Nya�%h8��F8��Y�����p�q=^�;���>O�M|���d7ԇ�?�ّ�DA�s��WޘH���,8}�3��#gID��8վ���yv�(ۭ�Wև��cϐ�d�#�~�E�[*V���!�b�l	C���'=��Q�`8��gT���>���5N�����B�g���|E�~T-�D�J�J8n �=��MTY��h[0�-���L��}\��fd3�Aj���9�_�dz��yH��*�=�`SY�p��-gu��\D@��ՁL��y���C1U�A6�Z%��(��p�ʛ�f�d�ܝW�:�r�N)��^tK���wz�:B�6B �f3X"N�A�ڹ7k��,����>+��⺴�Q�\|��޷|���R�a�Irk��u�:hЖ��j�i�z�e
J��
���7uo7ng���������2�P�0��p`!�H�H�R�R	��d�܆����\h�h�g��&f�.��s��OC��$�k��g�<UB�m�2��h��>�z�	�_���y_=b����J�������ӏ�=��K�fi-���2��$J�!����3�/w~�w�܁�8���?��zˆг��	���<�c��r�y�Z4-�X���v���]���Dr���8ɛ��ϰa&Jl�dc^p\+���X���o��K���Q��[�%�d���Td�.���s�sy櫭�o#�7/@�0EQ!Y3������I �`I7lQU21�s�f��q]��ckכy�^S�h'̚}Ie�=�!�xN�� M�V��l��n���B^|��'��9G�i��d�^�����;�zFíu�K	��|hO=�^��AE%��!�Hl���C�R��`2���xn�,ލChKx��L1p��{ʣ��~4'�l�ĐW�Փ>��quD�ª6�^+���;�w'�u��`����I�:��/�{��Ҡ_ޑU�K	�{r�C�#�^&u����<������/��@�Fq�O���N�$}%{��dn,���6TJ��H�����-���5���5k\'k�ʄ��37�IO�2Y�:�[����u�E��G9���O�˜���ln�&��L���E@�i��MC�u�ٯ�3��]`���M�+o;����j�4@΋O�N���-��]K����/�w3/�غnf�u�Ɖ�q��� i  80�C�Bu �0C0� ?�  �0P�	RC����v�N���D|�$��f	���-�B��;�tZ�lk�܆í��]��'�B���)���e�zdC�P�<I�hLL/?6=��ne �eʫ���WU��,�L͍��#����[�v�Y�׸п�vD�Up�:@8X[�� �*WҾ/I���J���E��<��|݃�Q�^pŏ!��.'�`(p�q�9�/�p|�V�����4G�@,���詐��>	z��G�B�Y&�~�p6}������w��ލ�ooI�F���/^��BT���#$���� _y�}*T)$���t�	������^|�<c-'�~�׳��}A��:_� 7z<m7�%������o��Zv`��D���%�yW�w T	9Ӿ�#�۬ 0����Gч��U��d��r��~�G�)�-'e��M3y�e�rY�!����7��zkԧ���~��������_�����<T���R��^w�w����%yߛ�٣c~�hy�&�4p�[%�qZ�}�7��������X����i]�3�C��=�DlD����G��#[9�S��N[ۚ#��FW7c���;w.���a�x׏[��Q®�,����,��d�FܴuKА�)}�ө`F��ذ����(��i��,r.ի���i��Sf"@s,5��0���Аùw=�V4v�j�ѡ4kv�|#��.�n�+u�l��C1S����Zu�%xfr���~ �Xq��\�Ǝؕ�ͮ��vE����e�7��v�;�����\�'s���ꉤ�u���[�R�|%>�����V#ڙضr# H��;e�ȣ�e��o>���&�B69պ������y�N��ջ�����N+t�{����Yp��gQAÍ�]�����(֬�v-J�r���:�u�(m��(6�9Mn�	��zY�`�+�2P}3U[xp��
��-'[��gT�wx����T����^�u�����(նy��6N�#���N���t
P�{�ʸ�WRM���97c�
n���R�k�Y�;�[ �a]���uAs��ȗz3�W
�Yk�����n�����F�M$���	��c>��x��垠��lX�n����u�5�ҭ$���v-�U���Q�`��뜸����v�+���2k��[ݑ6vKnE%ի��O+DWy����0�Ʋv3�'�M���h��%s��rٿXz�#�*.�fC�-�e5�8�A¸\�靝^�'��t�+��s�q�b�/��8�b�(�d��j�pV9����Tj��t27x���3^���n���T.K�k0lE{�٥f87<�R�mK�Z(m�9�93��DjMV�9�2�X��
n�9�f�'`+����7�2U�vШ���)��r)'PB�d�*����F}�;�-;Y��ɑ�`��wv��OzF�x땪I^q�VTB'��SR��vb'���m�B��m�Z�=7.Ib.5׸Cc&������x�(brڨl�;C����GZ�`v̘���E==r�5:k�{�|�^��S��/����mT�s:��ڮ+/Q��a��3m��^��f�%t#E�us8]��+B�^��PR|8kr������ˋ�,��QP��I#Wd�8��&sU�:�i�ٕ����j�}ǂ̸�z�f�05e��(S�qսVt7��ǕԚg��ʍݠe��«��WԴ]cэ�$�ι��LND�)xy�B�-�9f��u��kz���q�2�l�rU�1�γB����5����t|W6.�_v���|]��H �Z���i*kQ��m��z0��N�q�,L��W-r���ɳ���㏏������x�;�QU^��0���YGXW�8�5�ڊ�Q\�A\��W)RW����������8������g����7��
�%#�s.�EC)f%�Ա���su1*ml��mF��==>���>>>������Y羰���/hYu���R��-��Mj��D���2�ޟ_q�������Ǐ���֩�FB,�O���iq��p�+m^P��UZTX2̙6}9;�N�''��}>�Yg��|/�����{���*V*�
"�ܫ��J`TUc*q%2�,ɓ�QQ�qqQQ��B�
6{|�G���P�(���QUU��h�J,c�1����y�\EG[>c1:L�)R�r�#�UT�� b`���x�+2�h^ZJM2�"e���^���������$X�7�������īMrbQQV"#m%AD��Ex�D�pR�� t�]8���776`݆t��3rn�X���x^�ݻϡ�.c��K돳����qt6-��ڕ��A �*��a�C�peD�e �'ENJd*�C���^�#V_�d����c������Ssiy5 &U��sDHh���U9�&{S�3њ�a��˷��oW��ӹ�)���"a�S�0*�#�Tk�X�s���-U�M���q�=���ؼ��%�"���dn��*#��"�c��wO��H�"g���MON�yJ/��G�W%/�[�^��<�M�-*y��(�:�`o��6i�����e���9��Vl"HL?�4���	�z�E�>�tZ��P��RE�; �X�֎ALx?�.@��o}M)vw�gq��3�� �!�r|~y19�%�ԇ�OD��u'�z$`�X��� H�p�Ł�ЕN����Ѭ��.ݩ�7z����c�H��7����>)Nx�K4Z���A���J^�ϯJ _��g疄ϟ�T#�;�Z�s�k�͚ƈ/�3td��_#Ԁ O?��I}�yE��v��_��Bܦw���c�M�ؒψ�L�������<JO���O��
 5:�����a�ͅ�7�|h˿��aP�'���r��b��X��o�6�ŔEk>I+�z�;��{u7��F�ula�W�f)x+�J
��C�S�|B�"|���Ae�ª��V3R_�͓�FgT|���W��o�1]�����6rgY��},�jkξ�y�E�`�`��!�t2�e���{��s�]��r�ow���<a�PML>o8ב���ۯQ�VXHB{�<VІ���ɮ��a곔rét�O���Z�h����k���{���� ޛ0O��e��_�Q����Z=�&�~�8��Qh�#�B��?����1�X፽N��]zd��G��+��i�y�X���=���b��_@��V�$|���q28���UR���^��=���۴;��l:�f�	����������f�a��~�����ć"S�k�����Z��yttP1�x5����ʂ��TǠ����2���������]|G�r�p��:W"h|�j���d��������kc��=r��s1�(����-I�񋒬�_��a?6l�dmʡ��2)m�j�-"�I`-�O��=އJ1x�i�&Ѭ��^�T������{���Q�-�������T3nl�����.�Ư}q��zp�x܉� ��!b�0d�GLf�V�-+��K/;��Q���=�~[����,��(�&������������F~[�nvC�x�"&��vʙc��S�ԃv#ƍ�c ���굲�%�IRb�k
2�:*ӣ����.瀎���N+z��C��|�;�X���|r-�{;��CL{��|e���]����٩f toE)#���GG�w�5W����~�R�6��&�d�i0�V
�]@�	4��f��6D�.��V��  	 @��B��	��/�x2�C($2�!W���*��ei��>Ο�n@�Z�L�<S$�8t��zA��%��|��<}1�1
#�9獝�r�}w��GH�{qżƲ�����"gf �d0HG뒉�O8XZ�rѾ��#�_����k��82� �1��f�\� b�7���@#�������xH-���OSz}& M DűTj⹝I���WEi	���) .�)����X�H���=<j���6�8�}q�w��O,��hC�p��\��Y�`�G��L(�f�o��w���6�Xj*�e`˥������ ����.bX\8�y��τ�O<���rC}����I��-?w��F)�0���M���H����R��2��1�ʉ���f���)����e�[�i*��e���o�!���k��V|���7^N��d�]�l��,�kj���8�=���Aۖ�#F�3���������<���l� 8q��OJ��E�_1��7���	M�Ә�3����3)aM�Qm�;��2ǽC�9!��Q�'l#S栁j@vB�FΗ�{��ϰx��W홲Ȧ{����p��7�#�i�̡�q�7��V8U��:�h�T���X����=#�V,#ݹ�:ҽ�M���^X�v�α����[�6���M*�Զ�OaΒ��	֧���=��s����2P�ʬ2��]
q�e@� ���߾��{��/1�7�x}Pǣ�A�Z�}�gܝ[����G,p����)�5)z��B�^�\�;;�0���g�9k�R&�E��
0���	�Q�� ��C��Ȧ�Re�ȝ��+rX�r�����lF7���;��D*����&�ߧ��e����{�cg���Vi��,^C��G"P�d��T�\pJ4|j��y�%�̳ۑי9�(�W�%��8�L�X�:<| ��-��@#��ņ���ȟr���a�w��-ڜ�a���m��Z��K[����Y+�	����p�E��C9A���Ż�J�����3���+M}���M��F���C�{�� stD�UP��AB�����k��&�Oڌ����MH���z����H���w�"X�x?#捏���o;>����ᪧ��=}em���񃨨Gc_˺d��_|�)SB��] "�{�3?/
�������'��0ؔ=Xӧ�.Ǉp㦇��*Z�sM�([���2��Ң}�Zꂙ�b��\?S�s4~ˊC���wó�wCo�p��C6�.�T�]��k��T*��38�D`�Ћx�,�U�K2.�H+��I���lF�W�3s���n��ux�lK�nZ�V{�#٥쎶��;�L�4%��L��\����a�d@�6T���QLY�ϟ9���������ٝ���k���mt��P�5a���;��L �տ����&r���!�k��q�����uO�ݔ:��s^,��Q���U�U��]����m<�ne"���Izje��}ϗ�@G��_���,�TE�z�ĳ0�#���a�~sM���U�Kw��l��������c_�Bid�ot�WT���9���Ck�ȅZ�m(/� �1�N����e���[��������c�L;c�b� �K���86� )�0 �jR;�|����C���u��+��&&C��@U���5�E�.qF����ܼB�����>�����7ʎ�� ��7EC?�C��\T��G�{+��:I��m��
[���xe����;�<l��@S	����9��� ?�x���>�o�t*��:����bԡO7��J�t����ޑ��Έ�G�W�o#L��0UW��S�ST��hW�5
eg�7������Q��ҏ!�\�Ts�	��&�	
4�-.>��='�s�,�Y
F�킬�:�m4�P�ەa��Vl֑d��|��x$�X޼�����Q﵍�/��)��_q��x�p��]#Wv+p�'k_z���[�X��g:	\E�d���ی�ݎ1���e�b��R�W�;J�'P۱�{��DD2�a �`�	"Fa$�����u��%�71��yal��ܓ�IVJ���5��Ũ?#7k
l��
���B�b���er�n0|�غ�]!^�1PR��CWX�VP�0�����?nk�N�-g��]�� �H�H�p��!�����/ʢ��5#t�E��� ��������ŏc��N+�,��1�|vy� �z�D�':AƐ=fl�T,/�L�!�D����ѿoþ���?�A�<>c���3�c=�.���RbuZTa�V?|j��u�dk��~����9/��}"xaDq�i���[$�<�@wN7��,�U+eĽk��i�Au��5��T}9��Z� ��"d���T�hq����^�ǥ��w��7X嵬.
��;��,TZtxm=C����േ<X�<D�0M���?yު�<��n�����\����-޳���L�ꏽ8�\+Q/B < N�����5��l�k�~��P��r:��s�y��{�L���r�����44��Z����҉5���7W���{��^ �Iܫݬ��k�uQ�M��tV���ERm̝R�.:3������u R �a����}W�-i�8J�8��l��OLѫ��ݾ��~v�w~U�+!���OJ\q�}\�_Y9���e��,�m2��F�i��U1��A�
C�u0�B$`#$a$������<�����.���ư�o~�3���sr�:T	{�k		��# g>�Y�fC������z��[Y؆�{"O��G�sc��񰨿)N$H�.F�0�kכ1�ծ{.]�F�=���������C՝4j�����滲,���l�XZp\���=*F.�.50a+� �����y3���Uɽb>�ݙ�����j�v���]�Fc{�o�{�J�M�x�s�2��*�|��5�A���R��c���;-���a�nz_�?>�nA��Ж}[�tR���t�q��ݚ�^Ng\2��ڳ�ow�d�L�ǢAC���R� 0���C�L�Q&SN��7��Jik�d�#�Դ���T9w{��?9�s�;���r'} &'U}�h��|��J������XF��N'�(IfY�r�~�Pb�����C���yDή>�l�3��^>� �>��~9���KK9x4��N�Q��ߔ����|EEY��|�H���w	u/Ҽ�WR��<|����í.���N
(�6��ż��h�j�ku�����CA��Kǔ�IIAH� wɂ4��F���9�}]�n���v�#���Vf7�6K����-���K���9���mX�ӻ87�fb�@��D?�y�C��2,2t��!Ԉ�Di �)wkS���rrG8lx��@��W�m!�6ʿ
�</��xOv���{�=t��<���#܆���30Čb�����_Pd8�&���O�h$x������#�`w�*^�Y�&�yoq���푡}S�~�X��W7/@�z����;Xo�W��aİ<��'�Y���-���b���p����.~h.��	��e��a%�l�f8iRV5�;]����M;�,x���8\��9�N�O3�xm
�K�}�n|S�Q�����b�twn�٬�=�������5�C4����^ה��{Q�/�ϨܦM@�,���EGn|>v
�D����>�dt6CaYA�-Q }���>H8h������y��柋�cU.�E���-�e�Ǝ��_F}y:@��5hd��8�$��II _�/�D�_F:����!�6��w��o(�u��)s�9�Xi]������A��q�-�N|��s",ۮ2���#qe��^���tbY�Q�P(j��զ�:f�	�W����K�>�w�e�\�x�/2�DęM��.��E�T�,yC�(kS>)�n��˻I����a_��}����ͩaQ0�dh�^v�WlV �]�M��:�U��c�Ξ>R�`�����=/�Z{�s��a޻{��Ӟy߿���"�d��$FS�/�� �HxN��Ҏűc�>���r�&�}�
?GF�2�S��c���"�jȶ�,��/���P����ϻ~��[^�E�^�l�kNj�}��W�3І�B��:G��w�ө߭<V��ϼ���}0y?7-M�H�B� �>�X��л�p��+��|Q��p3b����ms]�ѥ�CvL�D-�ٰ���Z�f����ޜ�����2E}��R�|3,-�M�K�������ɺ��}�H���xČ��k�#�ѫO=-0sM�6���ٜ���q��a�E�r���u�{ZXc3.֊oF����W&��-Hnv��U��Q�ni"�Jl�#>x`���#
��{�ya���Qm;QT}��c��V9+I$���,
P���y +�&7��ئE�%9������!�I�K��[��d��_Ѩ])
�.W�0��/c�p#��Y2T&���	f0�XT$�����P�p�0۬]�ukn�`���D>ڇ+SHsrC��)��>;�>��]"Ft$��m|���s<'�U17ei1���~�ﺹ����Z��&�[�}ے��(s�@F�b�C9ݱ+!!�u����
�w���Z'!\�VvRVFq�7�Gu�r��������Y�|�3�nN֤����O
�?��aea�a���x0�3�{��xFr�*�HQ�,>/�U>�0�*:r���#�70�.^�v�q�*���j��m�����c*������i���;�������/}bWi_}�o�ī�3��.������'�<ޜ@)[TW��TqC[ =�كn��6�`�W_Vs+F�����	��ʳ�0�zek��WqT�yp��0 �zD�0؊Wq{±mss�R��/?�.���ʄ��LZ������I#:iA�N(�M�O{�D|DFW��f��D��@�S�&w�vWѭ\79>�;_�^�~1��ZWHux�/;��}�G<J�ܱ���� 2=b���> �%�+h�����fMM��T�>�Z�u��Q� 5����'�_A�G�p�<����cz�Ƣs�zS�A��"৔;AwD����5���X���H�<����>�gC�f!4�ry����6�򤕩	
(k\��U4��;�V*n�1L�%�l�A0�ް�Z��P�����ow*�*�TK���������v>��B����7U�wӻy�A�5'L�M]����V��u��fԠp�����
��M�Ո�qa�$��V�&�^���nf��bJ�}X𺩹�L	z��&�����p�xLe0���6�h�|�s�`�ObUѲC�-����:���z��f<+璶����i��E�r4��(�]�S��&[�L�ӻҁ�[Ձu�hdG��;!���J�_����B�L7j���b��v�����/{2�:e�tx�c�+(7+��;����O�m
~�}jZ�Mql�v-�pي(�(&v3vR� 8�m����O��1�"�8�4vժP����wwul�r��ժݙzGBB�wlFp���A�3CX�
��UJ��yBVr%u-fh7��p9Jzr�eV>jpQə��~�/X���s>�]��vm�M��`�JY����w�i�ѱ,��-��ʙ��5ꡇ�ڤT�7[|��/��D˼�Q3�|��awML@�c!.�!����+ (;�v��sSS�o-u��h�xۖ0����q��Y]Y�z��Yb�2�W;�8tGI'i���VH_N�b+����ls�[�9d�5+4��.)s!���4� ���b���z��P���&f�XS�Ч�Q��Ƌ�8$.�t{��0#�{��]��� �U
8/��T ������r�FVS�`WHUa��v�w���ܭ��U�F��vj�-7Gx��Р����b�oW]bz޽��)Pǡ�H�k�t4xR�������9���]0�Zܼ��(�(C+��e�D�\����H����Zyu*�l���#ϰ��g9B�+�urh����b��|f�;(�P;{mVgV����&-��	�)�,�P��S�q�lm�a�YG		����ַ��Pe�e����^��}X�rped@˙ݰR��{dY/Z���*��օJ��r���o�d9؀����~�����Ťdf�_/���xh����s���N<�u�9&^�k��q�\I�m9�{	12��r���MU���uʱI�����v o��l%@άT],��{`˭��!�i���*�v�!�vj�{�8_���@�0��,��'#U�'�_���Uʜ�t':׷��YU!���wn�b�v�r�Ӌ7"BU�4&�y:���t�̎�����_�f>ě{�q>���*��+f��!�}8�9뷷�[i��ܶ����ŋ�Lkd�[d����o,ɮŘ;	�t�$kB�i`�Tۦ�Ay��밥S"ƍ��x�\w�o.[�;��;;i�yƗNY�Dek糊��k�_RR�ۣ�'n��,�w�."{ܨ���*UQ�yCP�\I�[a�)R�_US�K�Fj�6hn0!qU6
F�*S�%D%6�I#A$�Mj�F�*lRt]Pq��d��J�b�T�5X�HT�W�k�L��r�ni��W��UyZB�`�ʹ.�ɺ4�,�h��S9!T�d�Z��	yydݥp�!��0N��:.�*��XT.�����N6� "&� ���%����|9���fWn붻��1oy�EA��c^f�RW�Ķ����ŋ�*9h���ٌ�1��2d����㏏����׏?Y���n��y՘�U��b(�3[~sR���CkC���z��:j�c�Ƿ��\q����������:�{q$A�mG�W+l\��Rڢ�mA.\��˹�bc�+S�rx�������8��_Y��?Y߾�%b%j(���p��`�-�`����h6۸V.Tz�<ﮊg���o���㏏���ϯ��#�>��So�R*�LK+U++��:b[��e���Z�ҹ��k`�j���'�g'''�������c>�3��>�1��&�w1T�µ-�.YE1����(��LJ>��m���/3^�y��������8����>�g�>�1Z0m+>h�Q���>SM��uZTkj(web�X�v%���[u��0-b&9rcm�lYs0UL��h��1���E#UE�&Z����3p�m1fZѢ����̦6��[lY�Qws&Z�X�O0�mә�t��jQ�(��9j��V�y�t���_-�J�iKZ�V��<�Lj:�FQ.[�e6e�LLp0�����vr��ޮ�
J>A���[ nYLr}h�d���u6�);�[}��W�ݣ�ǰ����:�/z��8w'*�t�}�y����C��֥���MB��U�U���f9����)�-3�7s�M���i�4�e�?������0NՐ��0��aO�=@��ؑ�˕�
F2�A�@��5+�����D4�UW�<\U���b���N�P��f��]����+]wm��wFC�`5٤M��Ao�C�2��d���ڙe%Ld��}��|�C�"�)���5�+N�Y^�V�}�rzz�����3����(���)�6{ö��4�K��ؼ�y��p�1ێ��t�G���tJ:�K�̔J����ៗĂ�ϑ+���5�����׾2�[b�%�7{�M�.O��$����Z��${ZI�vP&~�5�	9О���\e2��N�(���f�55[%�q��6��E�^�����*c^ݔ˧��P����+�:�'�y����{=4�	��@��mR]��H�z�a��1�_�c�a�:B/�
���#�:�W�Z��c���D�9(���r�4�>�՞��B�	�i�B����5P��<xr�m����l��zD�{/m�֢��|b��: �eFd�~��9��\�<��^Q�X��a'Hhސ9�PG��d{��cϘF��+��?t�E��n|���_l�J�]t�W��W�������'���M��v�L��S,T.��{0��K�V�Q�S��.���n5m8��6����nA}��4B�v'�{S}��{��P�����"Fd*H������ߟ!�����ղ0񵁎�O�[�cT�C�I0�Y�LI��2��3֩}�3y�w>��ϴ����A�����H�3Dq�#��~|.ͽŖ�I�t�����6`���f�O�fz������駖>e�>�Q��~�0ω2}@���'��Ԉ��8�����t��z�^��TF���a�w�.z��Q��?~L��`��ƪg�Ӆ��mz����>��ݨC:q�g�:�̠^b>�5/J_(cL�!��'';��?@�"OGϻF��uY~K>�^S�Vc�b�0�&�d�A���/-M0zO������B;��Z�.�ky�V�a!�130�N���F�+���,��:��Sm��n\��q��aQ�9q�p�Xl v�ǗY��;Xg��v�̏eiU�����I�p0��$�Z;+��Od�i�]�Kg;����;:c��f�0�P	��<�ԻH��ӱ\��Oƶ�rq�+͹��6�>��-�цд��,����`�n�:B����yl�d�v	QЋl�T�L��ɓMmu1y�ƃo�Y��A��p�:�1�eU��ڼ7��X����/im�A�:7�i819��(4-sݼ�N�u�kz�<�Ӿw,0�saӑy��BN��#�e�e&��Kd��������s�|��7����	?��H�$H$`���H�����I�3��?߿~Ϸ����<Z�J�iY7�%�輶�
���p�c�L0�k�sQ�V��t�R��t;��>�i!��:�lm����P�+�+1������)w����a���72�D6�l��<����["�E8>�/&X(������6oI��UC�ݫϊBW��G1����7I�28
���{�>r����_s��i�5�{��(�>�>������%qG>�>ޯ3q�+-C�H$1�Gʟ�a�;�얎ߜ,RjE'��8����n�V�n�sT�ͺ�w{&"�Ʋ�"&~�"C�~�O�Te�$�D�/Z�x��9f���m��-)�w�J�k�d��iN��dgM��'UZj.X5�-m�3��؞t��DU���� ᾵b��V��O����]�0|�Hn��
����(�$���9�i��fJ`e�y/�d��؜Ra>j�a���Q�p��!��JL����2<��`<�:��u9aJLH�	���?r(�q\1Vܶy����]�׶u�a�R�D�x����{V�0RuII�½[`��[�<��ڜdU�IՃ1`>����5���ʈ0Y?D���{���s�Q<���΋F���)�d��������S���&vJةWm�.�v�iמs�Ox�����-����)2���
FFI>I�������~���R��u���tW����񳥄��y�	��V�X��k2���s�kE�=�L�cU\���Ю�p���z�6�!��n�������{RSռ�����,]F��̹uZ������F��
 �N=������b���ã�$L 8>ZX��
~�~�X4
��e��^�����.Rᘓ�d6#M�i�ZoJ�o50�ߣm�L�D`���LG�^����r���˹�m)��F������E����F2�< u�
7��ޥ�}��2Iuض0�@��Z�L�6W8����1�wD8��8t���`Ҁ���5��p{~��k�>s�/-�0޼JE�laQl:ON35�yŏS0�v�n��jƭmw���+��~e�S��<D�7�*n-}�}��Ӌ���}&tm����m���͡���c
���Laa}�3e C���~,V"�b���ШT�<��L�5^9o��#蟷g��d��EZچ���'a�"aNs������=w����OW��w3�^�b�J��zz^<褽�|P���I�+: \8�2����In,������N�*;�u�)������f����(m�IHd�C�K�0tݛ�����CԈ��G������9S7���ln����hSs��C�@
o.	-+AIa6�.d�!�$���*f�δ��^&!�#"H� ���'$L%�0��+'�����?g��.V̃,6\ʙGH�|���?	}�UA7�kZZ�F����!q1ED��f��Ţv� {�B��S��އ�	^�Ѕg>H+�y�"��h�yʅ�W�L�R��G���|�Z�Ɩ]6��K�t]��`#9O��
P���}�&;�-�T��-�/j�L�шavǖ�q,J��}r����c�u�����d�C�7��A��{��WͯD� ��LP�/ƽ~��$u3	��vI������~�c�/���>�>8H<�c��"����Q6���!��-�&�f�@]�R7���4@��d�������6H&i��-��+ا�qrr׭D�Ud*�F���銀��>>�~�Qk��4���e�Sx�B��I��%��=�X���	�[M�0�|t�pO�}���#��_�u�qB!�;�&b��7�B�Hy�׋��}��9�;����&<�&?�y���k���mj�Qg�2k�f[m@���X+%��@P��3�a��*F>�����q {�����5��_��C:�#7�EJ��Χ���Z�E�{˷ޫ��I�-�t@��˪�5�f��
s��"��Nd�>�N�`&k��׭�}V[θg'm�=��:�J�F4�RI��S��0��W:���h`!�"�1*O�Wՠ�ߐ�O�'=�����b5"禍��V�����ͺ������EYZ�'����P��Dg8DS8z��lk��@P���&1/�;ى�=l̆5Cb��E���K�J�2�^��zcy��/�	%�lw�"�ϐ�c�|���7(¨�jʳװ�����Z��H��]��>5��1�d4q�f�\���"�3��鞀j'Cr�r�oB�|��̦E���)�7�&�,��	آA_*��	� �������u{�`����:�SV~�c���E���a�lk��h����{��a���yv��4�Ȥ�$f��0��?#��Y�}�bi��S�:G�9b!|]����-�.��	Ǵ��߽՟":�5�y�O�@��.m�/�G�G��@ŏ�h��E�b4�E����W�A��,�v���dM�����/%F��W!5�jνIRv��9Y��d�~�/����zcg�Mڿ�xYo?uj�q(��)���g������f9��5z享e�֝�ÖC]h�zb|�^�)Bf�5\	59�e�����=;�l�'3z!���~�����Lt���tVo-c�s��7�)�ZT���*�6�8���\'s�����M���*\���{�[Y`���\�B�"V,�@HČH��,'����^r��C|5�{r=z��̊�B����bށ�����ٝ<�X�V9Ut��ϭ����N9����k��AyO�ޱ�^	�Z졽p)��?1u[m6�Z�6���!��A�E�� 
�>5<����Z�[�9	t�8ј�]@q3
۹���Fe|�W�$9&�8�B@a�B1�"y��z�.��2ou}�.���yԃ)���W�\�I/�,6�m6[D��,v�`���|�p�[�|��OL�k�Х-#��+��{�0��J�wݑ1���li�]�|�~�>Շy{Osâ�F�p�N�:C��Af_G��3�V�����}�a3
Vc�]"N�G�7#dSS�=@knNF��Q�Ay�����o��w �����ڨj��rDl�џ�@��b�1����i���� �����!�vNp�ösh����2�������Ƞ��E�o�,RnK�.軆�^��Z����Kҙ�?
�����
����g��5�T;J����7�UC��E�'�s��R6����ie��Im��c69�ҽU��b�,�Q�U���)Ζn2�K��z�N;Y��^���~�%�@��߉lПЍ?LW6D�q͕��_&�PJ����]�i�R	�*�Y
sP��2S+l��t(u�P���}
)�DP�)�%��"D�RR$B��;�i���TNz����皗��m{�,�*���yT��,ա���7�G�#���(u�`��=��>��v�y�4ʹ9�-�㴉�A�n��+ԗ�A\\d��}}9�5��S��̤IRĹc�GZ@h(��C���'�/�a��j�Шa8����tnT4)P{J���=�i��W�G<�i���������0�*sZ�چ!�gz��!�A��85`��?'�������k�C���ۓ�`caށϖ��H��j8�N[���7*ӽ�/~���[��#}lK�S�䢣ϔ��6�<��y1�顖�*r��ߨ�=���ukyn�P�d:u�/�y{�3D�a�5���G8f2��zf�]C<S�T,�iu}�^��lNӎ&�_Ac���Jo�-�2����L��	����Iī��\v:�W��{�6\H�S�i��u�5"H�A��1ޚ:w�$�Qlgdy�*�Oʺy^{V��/Oхaz�ʳdM�Q���S���渴c�m����Ȑ���/�3ғ]�)f�!��Ob��Z)�ٮ���s.�:��<�����.����[͗.ZQX��9)���EsPf `d�j��� ]e
�+U~t�F�՛�U��%�=|�ݷh3�V�M��g#c�����K.M	���F�-1v�;�J�$�U�es箹��k�Z�f���/7*;��h�Z�$C��A&�k"D�|��a�}�<����ۿ���)L8�#Z�_�_�y�jOHy%�>�aʆ�Q�n}!YR1�<��&
�Zޚ�G�ɜL
��x̺<�߫�t��Kp�*~#��O�MB�*�rތ%��x���*�QQ�xwP��wP��4+���x|��S(�Y�41a�ϧZ]�5���UK��g^��m��k���-G����ԓ"�k���؟N�����vǦiD-�3�re,�u��d�Y�\I΂4Vzc��%r���L��ƘJ�OA��OCj�dO����v�N�v�7qh`([�NCha�v��[�*X$нD�j���/�:4��s��$�iōL�"��_�K�9�ߝT�2�lePa1�l�r����qX6�O'K�3.�s��kv1���m��?�.� ��Zo��5�������Gnu֩���k������*@DRlv!��{v�SȟyJ�`R��*��=�
a!1Zç|�3��k�0i�8Z+�3O����,�T��2�EYy��AyA@�m���OA�u"�tS)�{l\��cl�C��i�x΅c���Y{׽$'��7v^��r��nn�����b�u�?'j��9����WGw_2�Xn��F/��M�s-�¦��*_M�$'��6��o#�-rY$�5`��Mi�Yy�< �y� ��Il)"����}���������~a]����R)Mߜ��W���O��mϘ�*ڌOsOT�{�K�mL[�X9;Æg�q~���3�ڔ����*<��e{=P¼�[�� h���I:+��I�md��N���Hy��.���ߨV�)N�q�6���bm�r��j�Y�~��,6�K�=�ٴ�[dZ�-4�K[���/���P��.��u�}M�}����0�b߃_�'���=V"���<��7��Zߒm�#Im*��N5=dvΠ5{2u�x܉�A�rI�i��Ⱥ{оOC^�ȃ��Q{O.q�x�5�IӪ:7<�A �ť�T��^�5Ǣ"Ԋ�+��C�O)c Z���&ϔ	|�.�)�=/�wr��S3[w�hǣb�)��=!�����gБ�Ni��nŵ�jO�>��Ss�~hg�d��9~�p@�c��0v�:D�u/���iq��L�<�#�����?	�h:��w��gޱ�X�5���p/Q#����1 o����P~U�D�!�/?>щ�:ec34��*�/����~B�w�{v�$�K����W�&U���E�G��S�6��b�ζ��G��S(�JVvm��B�r���G*h,>�ӥ+mͼ�Nކ:S\�f��ٙW\��-��|�:�����t�6��*Rw�>ė,���P��o�j�OM�%ƃ��َ��5�4ƞj��\=%�oi�c)\vxID7�nu��z�z�����"�3�`����s)>ʸ�K46,z��E��wx��,?YU���ٴ�>�2,Z��{t��{P�����7P孙SrO(=��'o�M��k7'����f��N&��UY�̞O%����5-��J�����G(�}WM>"ҩ,�%듰��"�铛��J�oН�.�Q"_�v�����v�����J�w*��S�T��m��saڍ��ݹb�|������=�eg��m{x���t�otGV���ץ_j��;�C�o]�eeк
��yd�*�ۂr�ŗ2H*VsWu(��sT{'b���[|	]��o�����i�h.�g���de�JN�>;���t����+�:�e����^uRжW-�ո*�^vQ&pCHgeQyv(?AIZ�Z�����^��gou�Y��
ۤv�Jx�Y|��0��<;��T�k(�n�=�*�ہ9��~W��j䝗Y�L279���f�4q��q���6^<Mp��2��B:/:��c�_��v��CE,� [�x)Q��t;)Q9�9u�V����S�����z�7S�t�,r1�cu�hAN7�:p-T��3L=��t��CY�a��3 �W�Ϊ�ps���r�хN���,[��U����9���|�]͗aU��
�u�#�6AAh��*��_vפe�,�/_IGn�u����y�m� �K���ΠEۢ��J#l�гgoV��ӯ�"໔��o/`:5,���J�pg���$�;C�tyv���Z��GNl�i.�sʆI��5��8�����Ut� d���kIci���M��Z�r�lgb�ëU-�A�o%e�lܼ���\�غ�� v�БF;��X���-��/E�]�MVu�ʢ�S�h�B���&����z�Hʌv����]���n]H}ZkRD�v[�;�È��i���˪�iGk
+7�����&�UӜ�[�:v*��=*PQ��`�yz�h4�h{%���1�p(T+7�D�O���CʅI�|p�%�gr$������������h�VK�j��5����`�l�<e˓{�t�\	`�$������2��G�`���s+��@pt������еfZ�%��֩Ւ����3&8*�&͜���ΧS��y=��X��>�F{Z�~��U����V��(�V�#m�S��-F��u�/����ŵ�1�3�O�o����|~������V���UQ�#9i��Th�hԝ5>�"����J؈���h���Q\�X3�&ϧ����㏣��}x��~{�{p��|�`���5;3��1���h��t*`&Z帖Ҷ�O����<ɢ�ᔸ�T[�c��l������8���}g׌�g};��9r8�ޜd��QKiZ�@e�F5-���RZ�mV]Ɂ���Uj"
bU:��6�O,�ɳ�������?_Y��}�#�s�<+�E`ԭZ�UJŵjE��,�JiVT�nY��8�	�S===��>>>?\q�}u���w�V*z�kyn-��UWBL�U���צ��"�����`���娢#1mb�L�AJ���*s��~��J�(�b�"�UUzi�{h���`�Qbm�x�"�X�m`�Y�ŵj�����X�k���`��S�1ćIUU����QX�A���[e����l#��Ң�B&��Ǯ�n�ot�q�ʎo@�9�� R�.�E��૧�k�c�<u���T��O��D� �!Ė��H�Y#�~����s/���O�_v@LN�V�y9Q4)�#�L<^ /����k
��ƺ��I�8��'i�2��v��������X����>a����MS�����µ���܍̲�VO	�~"kU��zr&���?��? �a�yד�-�b�V�w\!�3�F�6c�y�U7�#���J3�F��[���93EQ�}��,�ﳏn��m�	!~|�����G�'�r���=WվlX�oo.��w��ң�U
09�Vx����wL�T&h��i*���L�&��{d&�J�٬m�`�3deB�421+�Y�C_�̆�aTcH��ØsT�˴�YT+'=*\��'���L���f���݇V����/�F�Ǚ�o;C�Z�|�	p
1����ͨ�D�L_�
�1��R�N����U���Y�b����7�����ZXC�h��/ye8�ra�K�Sn7,lሩ�)�z���wN�dvtK�Iq�҉�g�=�E����~����ݽ����c/ށSc_f��.�4�R����'t�r�U�V^؇�Sw��Upcj�)P��*M���,Թ�]�2�4�(1v[ԫ����.�j/s'C���:8�o�3��%u��M���������$�
F$@�����?~��� �yO"=�y"Ft�,Qa�1��Νl�����`���/�\��5Wo�ʻÀ�ې7S�?��cK�T("���
c��zD� �'C�XZp�هo<�h	Rm�D�F���^J}�!�v��kcT��N.�׊�e�A����d�	�ZU�X�-��9����̇OzC~xF�R�.�T�a #-�O��kKl�K2�+Q������_t����_r��!'��1�8�_U}P�
{��z�q�\�u��ca���}�ω�8C%n������%�u�-��7�ʴ�,�����`�Ӛ���k{{�T]NZX.�-�gmb�c*D��诌p�Kj@��e��a�R��4�S�Ly�aM�:o)�Q.1V�A�g`��i�y���0����� �&����vr�i$b-s���L�-A��Vm��`��Ҭ�l^�y^|㾚�
O:�N�"64ǇmBl���X��9.X��<�{>�4��$[�yv+���v�,SV�&��j6"r]�.;l���ڛ}ց�j޼G������:���v[<���9�NZ�"�ctr�E[Z�a\�Q2ϖZ�H4�x��iaa-[Sַ�q�F;S��gcCgU�@�ٖ'5wh2���Ϥ�j�I�� =8Sj�݅�4[DY#�:���K�ws۔�1�h�e�,�1o2�������H�D!$ ��L;Ջ'쿳%{~��ʁR�6B��8bN���_\����#�Y@/�Y�RC-̈�x��
�mOR���C��gЙ%�S�(��x���H�Jce��1�ݽ�G
Z"x���gi�{VH�~�l}\f�X~�A�ʄ+�����r-0��펎4�"zƽ�ڒ�m��������="uA�_���닾���[��������{m�1Zq�5��g���=��d}U3ʢT��>"/�t7$���:�Ifm�E\k,���z�Mz�ߑ��c��b�@|B<o��|gOl���-q0	��;7l��V���a�$/��2>���s��ع&BG3�;����#�b��9�ػ�=�8��<�=�Z~1؇X�^<z��2��]5$��X�q��M�7�T���V����۷��~d[WߕG��d�M"���_C��ӟ,8%����Ѐ�Q�W�5��� 5_u/��5z�w�^g�ޫ��5+�����c2]�fӛ��;t�߈�yuw�jK֝@���Oof���e���V`�A���	��)U�BT�7E`_���(��rm�D �	 #N=s�{�6� �r�y�	�z�]<�WP������^7��󽡄n�V`�;��#��#�$bF�"@�������_��w!�����0*x߳ל}�%eA�u�T�i��Y!�>��(���|��|-���iAR�|{z�O��z�c8����3[N�uq���Eܙ��#+�i�����RuL����x��maw°�M�4�7]�;壖=�g�R��zCh4�O9���Eԟ\Y��dw*����,t�hݽy�>�{Mtug�`<Ԗ���B8:�3_طp�0�$�=˯j8��~�Ü�KMpv~u�>���~�@�$L�`��C���l���år�?fO%���˒#���q����z�_o��l36���E:oD����.p��?s�UGN��ż=��iw䏧_ՆdJ�+(8t�!��t�n��2���B�_���?3O>�R �h�����v!�7�R��]X~ٵ䱷\^�텞��յՋR���Xۗ�h|��gi��t�t*�t;�>�զ�^��7���ha��%K�g��7��p���r���wj�V����'����8�Ԗg�G��X�oo��t��Ē�SbS� ~Y�'摐�# �O�g��~������gu߫�����]���#�I���.C�gn�#Q�{/q(̏��#L��弢��l������n�^�ׁ��ц7ށ��.�3o9�[�Wm\��-��_�2�{f�k~H�<��.Ft��IR�d�)�o��=|I�m�����=�D�a����5q�XDh5�n�HL+1�#Z2G����ң�ߒ;'=,�F ��wcɆۀ��}@UN_,�ar�����W����U��~�����ye�0J	�ܱ�	�����]T>�Vp�카ۧ;"��è��Egz�"���l5O����5��L-�����-�B��D*4���`���f�d�wQ��U<,x�e��nҥJ\p��Iv������^�~��렊�;�[=�xw�U�9�N�h�W,#���3QA��}^�^ڶ����Y>�4�[�ܽ�W�M��{p\�D��fٵ9�V��I�UY�]��T-���늧9.�0�Yke��d�2w��� �@Dq�3�8ܦNf���{���<��ӝ5��hU�&s���Qus���LZ��e���X��wٷo�Mt��U��͂�� ~cD ���80r�� �rۡ��i�wZ��gЭG?�E\t�&4gz[�{����>x�^a��?E�W�����M��j���]���	}vȪ���9Q�=It[��"![&�`�а�Y��":b[)���RƐO�s�=���� ��`ѿAV�|��� �}���a�N�1�\��9;����w�W�N�i�m����v�mj8f&�ڛ���^��`TsԹY�6��l�pz��q�㉃򐟪�/7E��mf�т��~��
�iS�c�=r�&�]���E
���t	��g8�R�{0��5�������fv)6s&r.��&��.�L�6z{b=\�>+
'��7��ӛ�����S�s�LP����	�⣫��Cl�hn�q4o��lt����t/:���^z	�G�@Ds6��
�g2,��q�A��'�����Ӎ�2ѵ���6��s��|U�\ZH�~Ըυ�W���C�O��b�=^�C�v˖�!���mϱD���Fڜ��g9W1�=�l=Bf�ޮ�b�9�ݏr�,f)�tjq�ޮ�}Ӹ�Ӯ��+��ݝ�(�-ЦT�Z�0��vd����e��z��f�ܺZ�	�#"F$`��@B���@9�7�g�喙�����4o2�O�/\_q�X�����c=I[�2/��1,,'���噜@K��]|y��{�4��u�%�v�E���^>B}���O���/��1wW�5_q�.���Ů�x�~��[�O�6o���C�\
���L�Y��\���譿B��j�zR����~�xj��`�xB�b�
��Vc��A��?�H�[�2|�����cedcp޵%l��Ir:�b�L��e���P��̷�:U�r��mO_�XO��c*ʧ̞��{���f�[
-:�>M�9m�J����j�vl��b��rir�����,��ت̀��5�*�{�\��!5%��0S��(��#z}����%�wU?Y`��,ފ�toq^�/&���cy�rP*\; �����+
Os{���o�_���#{&.��=�˥d�p*b�f�(��u��9�n!*��S]ƻjh����& �	B&$�����`�b���h��]]ڝ���0���9Wm^쫝
R���E�	�%��ky{������������wWZ�ޯ7�k��;^�I4&|m���e��f�H���)�ƪ���ztFv���dx�x^8)��x���r�k;��.A�ʥX�y�xM>H^�WvR��(�o�����}�yu8r.F���Q�tˡ;��7�&����Uo��8��@ё���,vR�0�����yx�<�5��|5����p��J��_=����=�Gon8FF��dǣz�cd��bǽqV����F�|�_������@��J��K����R@Iq��"L��S�³��3h[hъ��z�1�Қ���*�K�`�W�Di�d��z�d�j�Hrǁ��D����9���<��O�8#n,��&9��;�o�,�k�2R���J��귳�&��la��Ƶ�M�w�@�S �ҵ�V��im ��.���rl0�����L乿�>�.[�W�tT�ص��&p�Ѩ��m`s��Mk��_	ɕ�d��������>�+gz :V��rI�RF��wB�]��N�E�GG�S�껻eʵrqGǙh���I�� D �����}Gۈ2x�x���S�Qt
g��fB�
����W����-Z������ZY�.�Y����:��0�NKvi)#�t��KUv+��q8ڈ�}z�7���c8�܏;ߖ�^�'ۃ�՘����*�x�>��P��e�Z�o��׭ˆ���];%�j�i.�1�r�k��S��4�����2��뛛��>��`ݟ=CD��
�P]���BCތ)=gW�T�0�@l7#
��]���7Y��]X7��84w$����ŝ���.�}7!�����mWb&�S��"���P�ό�+�7���M�N�v�_U5ob".��o���K�
�Jw�PUxWt砑�CƊ�{*�SQYl��;[G>6�i븱{���iѽ������N���d���lO���=�+&�Y��	�h_��1���X8��:��,���m8}�%�ǯ8�Gh�Ў[�ڝ��.+���9�R�A� 	/otp��X�PK6� '�[v�n+�Jn��N��b�T����̽}�q�MR�W�e�3�{ޖ�,N�f���7�
��9*����q�N��O�̆��6���m������jӓUu����g�MG�s::��:`rV���q4ض��m(r�$E�p"[tf�7]��N��A��.HMKJ
S%2[�Q�_���VMzE�@�ݔ�7'�r[|�y��v���7o�k���U-n3Uϟ�*����I<�c�.��U��fH�q�S;����{lG�k6M�����o[�BO9�E>����V�q�z_MA��\�#�˯��ϱ��b�����`��
�^S�@��\�~�u}X��`L��7������!�����ۊ����ya7w����̌�RY���fVkٍQz5��ޖ�iH������4ե��[>������aZð:)�_�:"�����BL���X�a$������>�r|��a��E`�S0c�8"��OL �x=D@� u]+�~�BW_m��|�:*�v�{�7��S��_V�T�;b�U�m�]+#�\K�LW[����X*�Y��zN�z
WX���M>4��H�3	�c�v�U�Ӕ���=�wT2�	TFJ.l�G'q�R���v�	]ش����ʉe>oS��
}V�@���R�t��$ �!�,�,U�pd����]�;.���p���y۲��@�T�w٧%�X�y��j3W�S\��ܨh�A4�#��<���2úڝ:��}r�q�I���f��W���Q����u ��"�gƷ{BY6A���z��A+G!e�i��ˠ�MLy5���'�%c+0#�^W�Y�@�ę�]b=�vz�ٝ��G�WtM��ؕU���e�L�������
��A�:v`z^�3�)\ԻVDKq�.�\^p[�R���U�qu7����Eꖮ�jќ���5������m��k<%!�i;z��N�'�j`��>�[}/з���������Gj��7�t��N��ܮ[�U���ݓTS�m��Վ ���&<���6Xh(�$�ܸ�qS8\n��Z�-
;T���yl�u�cVm�T����@����x��*�ƪ+0��5(eu�H���K��uA���!ջ�b� ��{"�r�M��pa(��*��F�f�'VH�/6�:�)kU�@��e+Cq�h���\�75�s�:֙1M#�a��[�aZ�B#|�^a�i�3�m��vZr�ʎ|34��G7a��KPs�5+TY�m��/o(�ݷ(9dn��3�����܀S�܋o�؂�pA*�.��=�ܻE�<�lm��	4��RǴܻ΄�D���Lh�/��6�\KDz��}���n�uβ��enQn��ŴgR�܈�*3���)�dH��otFx�nc��0��9�}�n��sl�M���bF�r�ή[}�L6Hv�2���)i��oWt���u�e����Y[o��>={��C���O����"e]�іn��|������S�T�(i�k�pk�}}��m��Gc�G�	!��-�&�M�����(�C�����תC���Ue����s_ct�k!�ћڞ���6	*���o6���[��)��{F����+뼧v�ٱݽ�X�f�wwl1���yβ�z]a����c�������Rm	e�WF�	ܳ�w�֍�*������+n��;qC�V�p3%�4tձ�뿗�vO���q��w�X��&�V�w5��d}�a��Y��i���l�b�%[*�e� ��f��G�sm�@6�n����ݶn���f㹛�v��R�A�!7E�Tb��tR�%G�fT5r�2M{�,�E4lд�NR�`�E��4V�(�H�H܆�Q��I��($CaשmY(�J�p�Wʌ��B����D��#JP�h�KF'"�5��Jq!DUP(H�IS���Z=��ED�)��dE��Dܡ�ޚ�o-ygm����������㏣��Ϯ3�QT��R�UQ�D��Z�V�Q�m�EX�X��1q�-�����������㏣�����~�Z�~Ib�|u�h�lT���m��bTh�,���������������}=*=��!>h��5EL�
q��N����j���.Ss2"��ǧ���������}u���|t�iE�r@qeJ�;hykmAR�EƱ8ъ"�5�c������������}��Ϯ3��5�"$Pc"�6H���Ze����X�E��E�c6�('ǧ׷�������}}f}|g}���kg�t��֊�Z"*��k�d�F+hw�*��K�U�p�Q�U�VҊ�v�c�-++YZ"���K�N�QQ���|��0��j��\K��V*���3���1v���`�=Z��*�E(ъ#��䘢ŶTz)�[&�`�-u��<�f�Y�g7i���Q�g�N}��!ԥt}�n�R��93�<�o�o�wK��v����<�ݝ�����W�޳�I����0b���-Go2U�ix���q"�*�#M��=�ǘl ���mv�v�JFH��ł�/r_��6v�_�^������3�"=-�tN�Ǣ/uk��k8�����;����*�ū���	�a�F7c�����=cA�0��٭��5~�QӰ�2�V�ޛ��s����_Y �<�&�*/�����ơoR�gn>4�nW�FM@�vÚ7	�*�6eWFFȃ���k!��s$Fz��.FwdG�h�4�����)���E�g�^,�P)��=��݃�:��ձ�(�wٳ�n�n��]�a���\��[נOt��+Uw>^�ݕ�j-z�zx��t]�\�?��T��x3�l�,R�N���$���x�w��-	��I���%��;���]]~�}5����q&}U!�����9�v	̩��T���2|�»�{<��J�nͭ��JF=�c�&7�5Q��G��FG� ��w��f�C
[���3�J�2!�ڬ{,���P��\㛮YF�v�Vzk!��;TSh�vnT��'5$̺�U�ΣӴ��J����'Wv%ӐΰL�/�9�?�G�n��o�{�V�	��Zu�z<�-dG�vSc��s��Ng����A�ܒE�i��I�_���������G���b�ݥ���lUK�t�즼��Z��r��D���6G������o�s�]�/t����~Ҫ_�7F۶��HϣW��)@{���,�|�͎��'˥,��U���5㙒�6��K���@Z����I[D�옻��.c3���VO�Ǹ�/!��m�2A��ܯ����G�񖽦�<���Lio��{����@/bbf88߯]\C��`5U���۝�m�f�5��9������(�<�̎�N��Zse^�h�0�W�d��V7�2��z=1�"gWg�g
c�x�g���4UF�}��?$��Cw����S%#3���"��*����`U�������/�r�K�5i~��U(��y��iv�^�r������uoz�e��n����K���*�=��������. �b�^�ˬ�\�n�9�ͼ��:�qn�Lt�__l��+��������2+�;��m�	�A F���ǳ9��}s|G�7�*��VSP���0Z*��A�g���Z<��vM���Wp=9���ҷ
5e���Ww�1�x�����*�	h"��#��ܶ	f�hj"��.�ց3����w�R�Xɢ�zr�IL�\d�4co����d����ݺWt+��Iu�	�5�3��Hݲrxy^��ڣE�A*���q>S�&�Z�B���`������V��۹�)���xz���[xdI׿JJpo}�6�Y�mr�<���Oi=x��"7Xf�+;��]]+� s���	���Yǽ�0�'�z�E[Z+!#uۍ�˱�ϵ����$斉`��'ƛӵ�^���Z�{�)#�w�z}U�/k��w��+�ʉ���w֟�J��i�4��#���F϶
�~��Ό�/�2a/F��Tt��(�u7��h�bq���fcP�� :Z��҈}5R��lsF�������z� �u�/m�0�G3}Z}~�/8�r�
��)b������x��:�l���o.�����q��}��˔�������c+���CFu��%�� �@�۝��{��"���x�V�X��ޫ�0��|�d���:r�8��O�L��IεIݓ��g=׿T��k��H���eXɨ��x��%��^���ٖN����D��G��g�y]p>a�5�
&7��TJ���#uL����k���2_I��y*�����-st���֟�!ٝ�u`s��T����Ç�ƭRi�:��٠�2��;�Mɽ���^�2}1�3���0/;�jY=h�O��XX'���{bkP`�r��I*����ъM꓎���t�gt��	t��D_�j�c�3��Sxo�΍�eҦ}�5[�7[��z@��C'�bw\v��$^��g�������c�eC]���+!��]zbN^9��,6�ϡl9����%���Š!�ZF33��3�Y��F�o[|U�%�h��ޯxKa���d���0��s����^��޳�a0����^�o��U�D�z��S~��䆍���������W��Gk9����[�]�������n�혡"���"/�c~���}�_����Ow-Ǹܐ�[׋R�s��Cj�.���>Ck�[�M����V�i"e�ܵuD��+��$�T�]�iZ4i�̥o0͖)j�z��7Nd���&\����1vi�U�����$��q��M�ȝ�;>��g���I�F�zed��3;P�C�mK�7B~�q�U������G�zrbgط�����2c�C�i��AÑ^�� ��h﷭����O`���cy�0>4�N�{P/y]������3Ww,�B�#ښ�~N*A`�x"��E����tY�Nt�T�b��H�����rW@�P�h�cʆ�0��s6N�ML��3�g�����aa��ww
��e5��Z������qe1�+��>+$,�h	bg��s쟐�����Q#�$�������>] �{&�<�Tz�I��Z��x���މ*�Jm
�'���ts	���>=o�k�F��l��y���̝����:$�mK��^�ȩ�\]�W7�=�$l^S��V{W�����ɸ���G���h�.X�j�a!�U�3��u�����M5\�{���倿'�Q�/�-���9���]�p�5˯d����;��e��x�md��6�=��E	.��y�	���� �TC08�j�=���g�ӵ3>�7*s�m�������4��3�RJu�WS�,a!�\,oV���]����ʁ>HH�~W7�Qm����E^Z���Sʹ��;��7�1vKa�����#p��q׺r��]�a��hg]���'���j��n�|K��1�&�bM�5VNBR,�yR�����ɩ���{&�T���e���[��(OIޛ�h=�w�ɔ�%�+�݊�3��[z��+�b�ռ�-�1�B�_?>�4���)tDu�]������}��L�nB]��Sn[\'a���s�������mi�ˎe.��A�B�r���t�>�7Z�6�,��^C(�{>�ݡ'��%_y���rR}�!��Q݊]����N/aQRp�v�&7��b]�U��(~�V�� ��v������7|L��}L��l�Z�tD���Aq"�0KyU��6�<���:%�H����~�xY�n�|�nV���46��5�m�fO���{�J�h��c�-{��|���n�'�"{�e��vD1˄`|;����ʚ��
�y�
�6�+��x�)��� �<)Q�N����`����4U����" ��뭽��/F|�L�FlY�v�{{�Z�d����F���w�oo:Á�6���^��۩�3��"3�����!��]�+k.2K�]<����\d�)��}�%����td����$
's����ψ��@�#�nu�|����^Îx���'W��Z�S�&`�5�|pݲ�ԌW��o.`��uJ�!���BJ�����{)m���i�A���L�k�!�ύ�۾x�#��<���޷}��5���==���F���Q�t�3�`2g���H�dd��𘷮�Y0�k���W1c���nH\ìf"㫫0uT�դ]��7�:s{j�X�$ۅ���ڥR�(ɕ�����Bj�l!6���O^Av{$G9|����Í���"�g~�JD�C]cx & N������OiY~��>>�U�O�f�Q���Nt˶�U�����0(%K��	���-}Zm9t�燹�=��f�9�Y����hbS�팙�8����πk�,Í1׌ɗ��e8ov��^���F����v���]w�]^4�J�Ma�on���r�}�^Z�{��>ŀo_�y�t�EH[�X{��xENs?�����>��3��s�*�ܨ^���K���b���
��@'N�Ϸف�3�<��t�*�6Q,��Ͼ�y{�#A�eN��0+7�=����`��9e����tvzz{��-3/C1Y׋$P��ޙ������*�T$ZY��ݭ��u�]4萆ދ�W�M�BF�vL�s["5),���_W{)�m?��[���-��+ѹ��m�}v��D~x�T/��L$$U�d�6uVX����5�4|��}��{e��&	�C[O��D�z�<*MM�"w�75�{+K߭�3���O~v�j��>�PX��|�����K�z�j�R�L���6�Lߤ�+fs���_u��C<�U��y�����c��g]��w���
;���;�[>��d���{�=ȉ ��j��8�T5�2Luz��z��z�'�$ ̯{4Y�����#��&�e_�{.5M<l�քQ��BL�iUr�f���@\�0H�Jۃn��"@�D�f��ܠHhߺ�6��¡��f��Y�j��nJf���T�m��&Y���O�f��r�m75�?�RbJ�$�A�tHL�xt��(�IA�l�&���>d�qƼ���`�ھ{��V�0v5����9�Ox��]����i���oƩ9�[�z�*�C��Xy;dy�/�滼�v.�O-����{�^?���lЀ�j����89��g3u�7��z,6e��K�p�,9����r��{�f�U����Ǭ��x��{+7\����olu>%kzC���� �����R@�Fb��"�H�5�:N҄�7��hN����#j´u�at�>� �]bk�ј���v�dVi����$;n�M3�G��û�L�B�+���ޑ]�̆�e����SH���n��p��׉��Ѹ*��[�w"��G�aW�K8�r�re�Cץt�i�=0�l��i��j�9�@��k� @�'�~�s��j�z�R2�{}R��`�����~����aO�[��
�x&���*}/g���-n�p��8�8����`���cF���V�Y�ng��+�c���t�S���9Gڇ��k��.��*#7�7׫����]���$�l�W�J�kheF��V��s74�Vm���a1۽�">��0���z;y�ж|Cz��D��+��?�^~���+ϝ�
���l����;�w\��^��o��0�I���m�U�8�M;:���ݫb��/��]�����p��c�e�_c�z�Ň�U�>�a�#z��{l+�4m���2�N�&�A�om'��<����`�������F+�����ZS
��56N�~nBQ�wEҳ1��np�����
U�J��P�h�#
��,�!�����Z�[ٵ��y�bHA�,��wxvxog��Nc�ή�'�Ҽ��lf�
��7rn��.��m ��6����֒R:e��'��d��Bdg����:<��$U^�Nȧ���X*�
+�-/�*��^B7"�u�Sٝ<����x�.�ȉ����u�t^rN������>C�f"��D�"�S��i�����[i��el3A|��^u%�	��;&�m�)�\/5��&��t5��a��pZ��-��W��]H�a��Vq�v;���&N���qc���jG�����ub���Z�,��A/����}�B��k}��Jv�$�>J�,QJubt��]u��̋jR�D���������YU_j�zfd�gf���H�i���v,Q�LAݾ޼�y�xq�Չ��Pa�������ٺ���z:���Qw�//o�1�A}
:	��*�>�c�=Xx3�J*�;6�o��wʱ�$cF�F�k�[�3�2��k��1O��#Z��tF�G%9gW(�5���W-�f"������k���/���&��Ǘ�b�l<+��b�0�!]���|�[�y+��쥷�3]څE�um*iF:I�k9��YSEn�D�l��ܺ� \�&�ɣy�4�oS�}��ꩽT}�f^�,�������Y��tєiU=���(ԇ���0ޙ�i�䬹��)�-�.�uӸ����R�jc����0����!Y�h��+�r{�'��Rm��r�Zj=z^b9tq�E̡}�0#�+3�/���7|���J��F{)�a�4v�d#��iw�R�Hsv�jI�$['n�E�4-��ԓUR$e嗈W��kS2�&V�5�D�����eM�5��bZ�U�/�b�\ܳ�BQt;�c0󛝸n��ϵ�&c.��F�ٜr1��j�����h ����ha��&evqvp�i���E�r�c;��U��s�w�57h��m�զ�n��ՓV��|����W^/�a�ʱ����ۧ��8q@�!���r�D�ci[\��1�=� ͻ�{�U��r޽3睭T�/jKﰱ3���|��m%&!B�N	���y��aPM�Rv�L��M�l�yw�_[���u��2�WbWm�a�:[�$��vs�VAQ�/�t�Ρ�};xF�h1D]Q�c��}\�|OS�M���[�rhA�\$���pO�\�ը����Y�jR�\�䵵.�M�U,$�-���$�"�n4�/n�Ttu�u�ܿ�S��d�������pM+���ă�ܙ��B5�m�+	v��9��]Bz�5i�"��Yz��+5��Y@�T�iZ���8�.��	������"��8�h���7u��@�ə3b�cP�\��_q��/����u뢵L|�o,�\�-�q�l�a2��.
\K�}[�#��bɎ�sw��=�a��=��α�M֜e�]aK���ٚ�c�ݙC%-��]��*mX�V�Pcү:a�C��qt���G���93y�q:��m)ҳt���Ť-�ty�u���v��
^�n,��W���%�lwk]}������p�f%z2���(��:r�[������<��������1��"#�X)4�UPUEB�SE%��,��ٳf͜�����1�NFz|1^�`�B�չI̢�QEUQ6�dS��֢Q��}}{{{{{~��>������d��~qPFDb���H������+R�x�ۙA�}:�6lٳ���ϣ��gވ|�������J�EU�FZQ�1T|�T����lٳf�gS�x�3��:��8��������ڱF�����DUB�V�A�l�lٳf����}=�gӑ�C����T�Z+ܵ`(.%�J��YU��B=>>������_G_Y�_�n�b�Y�
�����h�*�R�B�X��b"���xY(�aPY�X�򲲢�=�2�PX"�Zr���X��c�MH�Ab�J(,DQb*�E��"�¤�X��QUQSl�(��l���x��@m[R��.�,r���ѡ$|	ń�s,)���l����n��:[��O��`��<9�p�ػ�_)q�����&Z�1��.�W�DE^���g���=��f3F]�#ه�Y؇PD��0���p�_4Hta����'w+6v;�r4��}���d1�4�}��a�[�4���Үg�3�=C4�-Í��z������<�ш�����-�nꬼ`}]C%NY�{�*��`s���c�9L��~�����S:2M�o^ܖ�R�$}���ݦ$?o�P��U�ў�#C�V�;3�I�b�j=�rW{����{���	�z���H�+���Z�,�9��O=���izv��lSz�W�]l��W�<E��f�K	܁vIuD6R(S�0)]�`�7��$\Ֆ�Th�at޺TX���̞b_ksV�p�V��y�o��	�U>�g���&�;ߴ-���U�����������T7Q-��_o/M�l�݅���t�$u-���B�<��s��=Z�q�"0��6��P��EK��;|� R�NJi:�;����<3��@�>N(K�p��e��Tv�>��7T���.�ԝ]r!��;/
��ÝGJ�����ofI�i�*V����k	v��2 ��O��w��S������L1t��o���.]��k�Y���a�"|�I���울�c�W��A�<�QӸ�-(�jn��Ӌ���쇶hqML&s���ζe�[2�l�q����~oZj�"8� ���o�_��y��x-�7s�J=3�Eﴞ��^�q���z/�(���D��=4��\��VM�	i,s���_�٥�M�9U���
�]��k��pҨ�]��N��9��ٖ��ێ��1ci\��P	�����`�gӻUmv�	uZ�˺�0Ȏ͛�a�Fg}{����m�$�YA��L���A�,���*}�1�g� ��̼����Խ��ey�^1��n.͊����b��:s��xk�R���wvp�,Tg�Q�c��#}�ź�Ti$A��x���	�0���as����k/ Gty��
O1�	c����<���iܙ��-l�4��Y�Y�sZ��Iϕc��1Ve��r��z5\����L��>
Ο
IjT&�v��JX@��څ��Pϡ���Z}J�|$��N��Gp9�p���>E��}2[;,9ۦ8��U�tU2f���d�]}�S���t�}zy���z��bT���B�}T�$5)��m�u��nr���ۮk�7�@�-15���{ξϽ���-�� �t��p��ב��=/�
`5K��Zh}��b!l(��6s���ˠ4l�y� g3���fs�~�xXK�O����r������#.%��#7�	���S�ol{I�jM+j�[^K�\̙k�8�������,bI"�΅��8�>��D���ѹ
7��;2��PZ�ζU]w�c�M�`&�.����)��]XW���qQuD�?"'�f(��ԓ[���s �u����!/�X�_VJa9������_���I�/�n҈^w����6�0f�Oe��1��A�¢��eZ���ϝ��h�Ïٹ�7��g�d��l6Mʨ*1E;*DW�b��O�=S�3;D����S�`��U�	�c�7䴓^)��oq��̴�k�ut�����|���K=U�]�q�6o.Y�!Ѯ�w����|X4x�C�=�pl�sZ�ȡ��
�( ��l�2�"��<����dfr.�!�WTΥ*�����6l����ȟe���w�R%[���}�:����eӝn�T���+�ںx�O3�HC�S�����nE�vKW!c�{<�.�So��|4�V��'C���}Inp��z^_w��Ǜ�|�N�]�"��d[;[}�]yq�o_L+��9�]>������P�<7�z?#H�;`@��Q=g���j-��oc��l��Gz�ў�=9�~��F�T��=��s�9\�7M�6�'��.Z�j�������<C���eq��C��NdC��>��io_2�&5����5Y0.���s/Hb0��Y�L<Cu�S,y���NƸvv��;!�%������ 3R��O��|7�<A*�!� �x���'+O�^�,'"+ՕoV�lbe�2&CDܛP+�^!�r��,�-�Ǻ�*�H%bU+Ӗ��l#UV��i;��R��E-��k �;���o��ecy�I*R�za4�ם����vb.A$�:�͒�E&o��f��F�dr�Ս���h@�r����������!^���ꭼ���V]�(���nf��!���8@�_[8�ul�VK����$v�����:��4��[FJ�*U� 2����`�y�/�]��[�<ҾF��C'zGBܮ��)^s�;����8�"�Nmr�nр�T���=��KK�ɣ)J[���U��\���~�(��oV�/;��}�-�s�z@��g|�u-]���A�Xܖ�\v���w�@>��/s��R|lTl�)�\�3��Vw��@�F����t�PiuI�&�9R�
�;~���}�F�2�`n掯Tj���i�3�n�5yWLu�S��ĩe�n¨t8�p0�G0h�_�s|�Xr$nR�Ng&�&i��{%����}FC�P`͌��e�40W�zA�g�wq�R�J�8��"ע�P2��ne��|����_"w�	^������eZ۞ӌ���X:Tk��=���]���j[e��3��}��-�s��6V){J!��5pَ����U��l]� �\��I�a)b��k���Dec�Y�/�N��DەN�z�Ʋw~��W�|Td*K�=���tߝ=P)������^���'��up�Yw#����m��:��5�r���G�4�<ͼ�z�_���%H$�9�~��ގx~����u�`I�Ru�/�b��e0���D�y�E�@��wʜ����C8Ĕ�z6���)�ϘC�]�F��>������Me�Ϟ�p��h�H� }>���&�VӆϹ�X�Z�{МL����@��s�z�+a��R&�W��^����j�_J�Y�a�R�8�8������9������'sw�qw��.��0�5�~�gL�ï��g���57�
���^�-�����ʵ�G��j+\���6�V�z^#���޼���Jc��U��}A3%2HJ7���%w�:y#s
�+[/s�yr�/h�����~���87�t�4,ю�b�6������6v�	n_?<@�HV+i���`v���Tv�;�����Ci��Y��L�DYS�{`a�ŧ)�|��߱Q��qr�z{���qWl3[u����Y�J����7:v�ˢ��8n̈�pf�v�`��^�Q�D#<Ax�l;SQ�n�2	
�Y!�mQ�üJ����:v.}���j=�T��y��WfN��]��Ż��d�z��,�e���eel�6@���ݹ�@��+,�Q#)	�)��uB�HӪ,Ӣ�B5
a�(�e�Q| ��ڵ�>��ﷶ��AR\�)$
��iܐ���9M�Rڌ�^�|����3�8����=��s.�ˌ�dW���<�E�n�1�Uꐤ����0�
M�݁����ң�.����}ze�����ۇ�x��.DY�϶ifIm���e����;�����3�^�ί>�aw㞱}���|�k�O�)�����B�b�c���1�/�CvYa��k����66��4-�QT�uM/v��*��@]�3��pqg�����{^=Pٗz#�(��ef�J���P�U~�5�d2�x׉wgg�W��D��g�V��y{�C�t�;�j��{u�AA�J��T����eW���G{M;[������J	W��u�{ְU�/m�W��1�,���;��4ӽ�f�V����٣]#�ԕWs)'gfok��o*�����弿O�nBȐp��W�Dx�)[�`=ka���7��A�E�7��Gh����g�p��1Ѽ�i�O;J�@���(��.�{�S��y�0��ڛ��wJ�۸��Q�3g^�W`_<֝��1�ܜ�j�'������ �Hs���u?�ٛCF=/�� ��	���&�W��4������ڟV�M���O������,�Gܯ�kf9u�;s��f�L���s�V^�-�z��:�ym3����DP�P� �gdmt\���Kd3w�pk�S�o���/��x�=f����O7����q�=cqȾjS���;�f'oJ�r}p��ŮVd޴DL��y{G�% ��Ӟ4}�\�_�y��)�Q��TçZgC<�wf�MM�q��fSR���>u#�z����n���l|���*+���voo���7��[�ףNrƮ���5��Y)�������.
�D�[Ճ]5�J}�^>Ǡ��-y�I�~�t�9A��2,; s��B��K�������� �y�9X�T=�~�.d��9���������b�����|�u�p�<����4$Y-)�ڻVU�#YkrPʔ�(�n��.Ư+Gv�{������)�Ȫ*�g^�v���Wqz]�8�W���(���7|����W���0A�fj����6�"�9/�]��+�辙�1=�3i�@�u�O=#0���vtw4�������a���w!���]S�a���!UN+����n�}���m�꯱��FU ށ�m����}5Ng7$���j��ZM�(�]*BWk��i���ӎ�#��ީ�!�~���!; l�
�0�^�G=��X�ޟj�D糔J|z�tu_�늕y�c���(�B����g+��}��KĞwx����9�}���p�Ӓ��}���Մr&�z;�ý��(�wm���X4l��{�F<jsj|M�����c�5�7��z/�>;"�U��9s����|����=w���3��d�M�s������]�,D霺�ꎡ6�&8ǕW#p����;�:��q��`�9���Cee\�׺�	�f�߳�
� ^u�ƚ-���fz��{&罋9{
���V�y�!$�*T=[��uc��{���MV�j���ؗ�8#Ȫ.�����O��۾s�)}f���NlL1�����X�'���Ч;�ݾ����}}��KpqH?\0���/��D��������G>�N�c9�]��s]FC� ���7�l�,,���тg�X�ׇ�~�8R�L�u���C���"�&`�ջ��<�-��k�������f����1�_�GR��8*�ݐ����eQ�]�f�{��̉�﭅4����y��}�Y�=/ IO��nອ�ʢ��^��x7g^�:�S�������r�����@�/�kiP*כ�MxZ���m�.�� �ʡ�[\yY(�Ȍ����
�<.�ق�f-%�Ϗ���x���ʌ��x�aW�y�~���^����N4���쿘��dK8C ��y���.�)v��Wk(�oO;W�pm����܂�T�����\Num��o�	�w��VPa��߰�9J��R�Ǜ�e�K�)͠[x��$���0�w��������y��m�:꽡���'�^���]�aGi�A��wmt��Bq-�zdYW�;y4��(�غ�U�سo�AAp�Ӭ<�WM����;i�l�O"�u�w#�Wj<�jhb�]ڦpu^�{w	�',�P�"o��Q�8�n�Q,՜=��i?_8�gt�)�0�F��������R���lm��-�ՈU��B��
��Oz��*��y�vv�\n*�fd���\V8�sI��uM��e��"�T��=�|sh�q���e�Q��,w�4غ�J�Wr�[!oe��]f��-f$b���ܹk�y�˩"��D��o%e�<���\��Y�3f�e>��Uj8�F�Y��+.��-��Io*�yR�ӡ��CP�����h˺�Yb��u�f�fu���]YP�=��c�y�ڿ[�Uo/۴`�CiM���Z
һ���|tfm���Q�K6UҎ[?`<(*_R���Tooh�(�*���ν��e��u�;��#�u޴:��j;� �+͏I׺f�����űJ/.oUeX�[�O&���S$�撨c�I%.�j#���r�S9X�;)�y'V��]Ah�Tƒ
�&�� ���Kd��}!�5�5GS��ZȆ%��"��&�v\��f��m+x��r+���é��~�x*e�N7�ٛ�틜�y!�K�w�y�_ڣ[�]T9:j�J�2��	d2"�h<P��[7)���,�В*$E���JI�(��D؂J��X�6��d�c�Ԁ���ںFԑhV�{��VX��N�Y�]�6L4�sr�k{E�/�v\�2���3֘v�&�s7)K��o*�v �g�dN��)�%�
�y.�X���u�Y��:�����V;���=zT��]��f�3�kNֽ��U���Y�M�8	���T�z�{r�!(��E�g\�Xl�v�;��I���j^X�.��qU�ӮFpo{#r��ݫ�mNu+��YB�l7T$j�w�c�a��9nu
��u䄭3l�[�U��9�9͏�ا"�[t[�3qꉂ+Swr�:�Ŕ����=��n�vV5�!j���ϑ�p�h�A��M�
�]�P�eN#m�d����5��y�H�Ա�㨐�*Vu�R^YT`���|�p:˷��U��Y�'�J\�-v3qr�C�,���r�l��&�˗4��v�{��B^��n���C׻[�k�8���2��}x�{�fn�/w�mJ�S[FFۙU#��gGTяT��Pᮛ��n^�7��v�c�Cz����waE��������i����i����,���ţ]o#��]��Ǉ9]��\-��p���hH��E[����4]�f�
ðK�#�e�U"�5�&d)%��ʉ
$��GŲ�
p�����@�Z���LQ� �0�P��d��u:�5�'&��l׫jFb��/d�L��]��%,H��c���%I�"�3G2�����_��EGiG��QQEuJ(#�*DAH�,��{{{{{{7���O�ϯ��|i�g�r�X �YE�X�5��ZT��PQ��%�>�5�������>��>�3���������P�jV�P��gMb�r��س����0[kgӓf͛6y;���c6|O��4DEƈ�W�Qgys�_]�X�UQUYZ\�Qg�-l��ٳf͞���}͟���*�l*�f)11\zk�T{	2���̤�{n�^>>�������~>���=����T����4��Ac���`��|Sn��x���{{{{{~��_Z3'�ϾC�=�c�j�fbͷ��q'�
(���㹊�����E�,5�l�.Zl��5H�c^�Mkm.g6k"����SiF�c*wk f���*J!�Lb��AdXVT��hb��(�+Sónd��͚��FQo�n�}يB���^�d�#S��vL!M%t�{�ữ��5y���=5c�M�S[�C�����*W�5�VT�8�(�))Fnҏ+�sZ��*o�
�Ü�2zg(����HH�(��9� |����֑�3�_����r�^�؜��8/��`m��ML�]�U9�����Ս�|W"��˯=\�^,V�O�(���Oo�ع��x�Ed�{.�ɚ���O�!/c^^����^�j̟C��t��;/���Хy�ۅL��.jʧ�1/��հ�[��SA�׌ǰu�?�g������uu��,܉9���oRe#]�z��ϗ�i�QT���Y=s�U��W�� ���`��wE��6u�n��)S(��y\q���������u"Lz����~'j/�s�X���o��)�Rb����}��U�_6;��55�e旲��K�};�/�l�h�v��y����E�B��j�~7�q�L#�a�ϳ��i��XZ:\mq�̩=# ��&g�:�g7,q^CN6�.F�G7VU�Ƀ;���i��0�r *��}y}D�u��t��6�{g%�/�aȔ�o���%6�͂6���D;Ϊ���ܼ�,|7��d홷u�	���j�ѽ#=��k;�F���Q����W|�z�}9�G��@8���wlt���aN\5�jSq��4�@Dl����75�.;{N�L[/Y��\��i?8�|�;�~���W��P��W��ήpi���
���zN��O�]�_)�̗�b���a;��/H>��\��Z�<ǲ�=�����W���R�vJ���8����od�����(��k�fO��6��p�>p��YܠJ7��q�1�9�bS����m^g�&��1���l
6Ѝ{�9+oH���a�-�_�)����3o7�`�&	H��33��?����0�a�};	a�����XBT�1�:��ݞ|���w�u���q��`���L�Xjʭ��t�[��k^�k����h��V�8՚7n|��컦/T���M�CL7	�:&7`���������'���0m��́2�+'�/��']�E�xS5�$��>�����Ϲl�j����}��k4�5���(K�z�@
5���lVP����O�-/u��7�$�.�Qe��;r�W��hUy<�]��^�u�e'aHZ��d%�y�.���C A" �͓�9�G^v�;e�C0f��&}L�#�g�2�氱���zø)u����k2;�;��
�7��ީm$�Z}��h�4ٛ'���l�_`� pm���S�)5k<7��ӻ������c��.("����9Ղ�i�noSFC�y1@0�h5�]�9��{��p�_�pfz�u���S�މ�6��f��=D���A%bl�jR͆^�5�rk)k������Z��.��BX��ݭ�f�S}�@�kw0�^j�Vغ�vjׯ(�^M��\��:MV�ט�g�;��WuB�9�X��54D�H�8�Ow�غ�o�,ⅽ��Æ[g����2k�^�B���lU�v���ǰ��s`���7�6vM� v�7�q����y!J�\��x��E��ʜ�~��5�$8X�v����K�iמǎ�{Ow5��R��k�����v�hKz�,yx�u�V�]2�R��x$ĺnUz���-!4��LA��
��t�/[|V\������}b��D�4M��ӸĐ���maQ��g����n�{���x""v�s��ה�4���9��㳌�>{���zit��S\��SM5�bi�$w�Pu���W��,�@�m�5��u	�y�|�|����	�>�����R0M"�d���?WH�# Y��ٟ]{�/�
���V��R"�~��	�;	��.�c_�8+3#�3��V{J�yR�K���.w���b*�Y4�z�{j�%���۪cSi��uk��y��R�{)����EM�y�4~��i��n�V���^èV���e���1�{�ֵu��x�گ=�t�W�����Xo^�l�ǳ�v�ӳ쟪l��t�f�^�}V\g�&�]���g��\�%5Ӷ���r_�f�*q���
+�z4��E�9��o����=�}I[F���s�����ꀹFrě}�(�.i�}P�ٵ�Фo�&ޱHq.�cd���R�w0���R��\���_e��[��O��xV��U��[�k�9(\�Hm�;V�(����a#��oU�}}�6�.����PggVN3t��wq�q�\��*�-Ep��͠���;<���¼���
�iʺuhF4��ڨ�1�ӵ�
-���_D@� �*�Uy=�sݏy�F�ӧ%:E����^O����a��L$Y���]�q_�DR�xŷ?G-���vQ�6�X�h1�m�k���,�t/{��k���w�qǁ���3Y�y�o\����n/{�ps��6���B|���}��3�7�j����σ#]:���R���h�;�c׃�Lv�����Ij]\'�`�&�]���0�z*f�Y���Q�!�﫭H��N�� ��)n̒�p�O�.�NS4�4Q{Ǻ�ͅ�v�+���QKd��J$�w�ǅ �A����9�c�ׄ��Z89�����
>�������Ҍ�oM�����>*�	���sSx��3;3�ݙ��w׬r$i�3�L{UAd}�~F~�ߺ�е�,��[�`�c1n��L���[�,,���fʟ���o�K��5~qf:S)�����H�X}��53T/�\7x9�E�Ē�-J�WA�d���W{ZD��%Ї8P$��y*��`�J������O'u�;sӜ"q{e62������Rf��#�5 q�l�%X@^˦�o��_x � �k�֩Y�=����>�	Lzt_0��^~�>��i�gV[k
kj���y���º���Nϗ�H��d�ѐi�����txC�ּC����z����_y���{�q���@�Z3��*B�a�f�m'̲���@��>�^�������u�z���;{`�k��鮮�s)�^�s&�w�+I ��A���C�\5�ک��.-+t��cxn`{N�ψ���w����=��7���\�LF��^3�)?m�ud�23�����{ߒ�9cղѾ1��1p�B"�6�Vp�� Y9xHޫ��B�B��+�0��+:�F�F$��#��%0[	\<���WR��U���v��T.m�n�^�CP���h�{�uwù@�o+�mD��yA�oF�-	�`�/_c��8�������-nzVPke�}��S����0����8��'s3�>\NN
y�������$��G����I�e�
�ܩܳXQ��7�s"x���m�V ����/1s��)���Z.�ʃ�$�o��r����:���L���t�#Q��l�M�'��ú��� ������v:~vY8/>Ʌ�=�(�2$�p֗x�_>�5?�y׬$��n߾�JF>k��2��o")���ZU^һ�q��¾��ӝ��XL����ðq�$h��綼�t�8�R.R獇��MU�׍�Fdi��J�U�=!�\i�>���{�ػ�O��j�Z����}Ǹ�8cC��D̠fNO��u}0�{�����_jL���vg7��å��vGu���Mys�$,�e�dlm\k��w�����T�o�|�p�����3��e��y�9���oxz	z4�D�R-�����ǘ�K�a�*��5��/vs��v�}ڢ*�н�i�fUT�
n3�=�,;I�J��f+��l0��HۢC)�����n��g���11дs�b��i]��P!�Y����z+U���*���\9�t���m�����9������X���jG���ڙbJ�ۅI�o:��*�x�w5��J�&|��hx�@kL�D�` �E�hs|sw�,[{�*��g>���wΝ�ׂ*˴+��d���sV�'�RR��$���)����,�������6�UB� ����`��r������U:T`�á���#�c�v��;��֑�"��J�uS���S�5�gd���I���D�"���Ƚ�n��;��rEF��Y�t�E�n�Ss��R��ud��6�(���0�\�y�
�qu	n���z8�Ȇ���| ��ꌲI4�Jy���g��!��oD����P�ђ��gEয়U�i���S�_`����=�h2��
��ޓ��gv�5d�wɬ|�=��Q�ir�s)W������4�,���Z���I;����e�Dw�����P��V�L NG�K�i���K܊3BD�Zjy�{%�:�Lߧ�0�
_S��ߟ�em�Kꇗj|s3�1U�ޞ́<11^���
���pZ���ג�tk��P�p�F�ko/6C�/x�ޖ������c��O���z�u"��&ܩ�cH�^�V1�S�ܥ�ИRuM�4�YN�MT7�(!�;t�\��uL�p:}�R��O/��,�6��)���إf�b�C+��p��&y�7B��؀���f�Qt�4S�Ah��UM�%j���DA�GOzMk�{���S)RD�v�}�w�*�!v��;}O��lY�w>.%� ��Ҟpo1M�[W��j���]�5[V�*��"���������E�I��+��c�.u��u�ӁL7c\�> <F�^VYބǲ�R�r�W���Z��2F�w�^�~&��^�ڼ�]x�����0c=�m���:8�a.���'��f�3Ќ謱YW�];��2�w~k�e�����y>8OfС�/t�[���{��ﳜq��k���39f$�x�l3����}BVn������+����cs���\w� ���uC�I���9~�>����	S��$�9l��d�8��nDnV_������������׵=ӓ�r�	�D�n���c��6�R���̓��p����j�ek���H}>��W���V0�jH��ۍE��W��]��z����j�^���f�yȚ����ǺǀͶ�3�����N=�E�ɂ�e]�g)�T\���֥ɣ�*]kɽ6�\�5�y1%r��:��;�(^AA+�]�%�˚,t�I���<� G��}��]u��`9>&�`ǭD	|͠R�vUyˎ��ix�`}�*���N�o�]T��H�w��P��衏��0�50�k��;m�n#��4��6�/|���z6�кM|���e��v{�ʵӑ �<�:�l-�G*�ֽ�nB�-�h��(�`=�>I��ְ^kc���*�n��~���~��Xȝ��
�}�[�ʲ�6��!nH�����aXC�F|�1�H�9�i��k���p�kB/��v��l�ҖH! �CH�<���f�mN*�}��+A��5�4ӯ,��C��=��2Dy�a�(��MT��kn�DHh�L<��b�۸�L�07��P�e��kv�}��ɐ�CQ��{{EJO�i�MM����sK�Y�WPd������LTڠ3�S������ʰ1[2��g��zY~T�!W��V��]���oV��	��]Y2*�T3H�q<:�0�������d������
'^I�aR�#C�Jp���|�1��r�C��;��G�P��l;K*t/6��!Y�5��9|:M#��%�9��z�{z�u
x����\Ԏ!�*��8Ҍ�}��X��1���x�,)[O6����W�
����W�NA��dn1RI�i�2�o�7k�T�j���U�B'��ά���a��V����>���E����I�lP6�4�q�t�4�:�L�W�2��c'��9�.A��_nVk��M�x�o.���ȯ��Ynve)l�I�!�|�vj��r�[�	ҦTr�u���K�Jvh��"��f	E�ef|��[AwU�	�,��-����[�l�38�����b�'6(՞[��SG�H��ՃV�cX�^7��êIؐ��N��N=��_UWA��0��W5���f�|+�g�f�hC]�zm���P��ѮL��/v�f<��s�P��D���0�x"��k�b���,�4��%�����.� ?tt�S���9�V����otN#�Ŏ"{I�ZZ��r��z��,aj1�t0Jp����n���$�w����33�ۆNt�rrc�#EJ�;ʯ��!ƨ��G֢�d���@�\M��d�Y�Q�����\�s��%tm��k!GoCq֤��98�ŕ��Y!]Ɍ�_D��J�^�M%�WjK�6��GH\'����|_��$q�������@�/w����CI�\٩�V�-�=*l$�d�����Dl�����S���4~mA�j^[�;�+�WT���jWkbq�4ٶ�/�䔤$��h�Z.e}�jnTr�eB]K��u.��Wb��ҭ0)�r������BOE�:[�@�g�at�}�ɴ�`�۸�o�W��]o����g�5�mGw7��),F�i�����9u(C������jv�h5�sB���I\;�n;k����[��V��2��CoR=��Y|�ñ��O�����b�GZ����C�7��Tk4:���ڮ&�L�<��	�ݮ)ڨ���i͊�p�
�"�΍����a1��O.����)TQS�[��J�����Z��+6�@G,޼XL�b�gl��7)q	`YmT�/{S�΀�����:�x������}L�4a�j���ړ��vV=�Y(����]جR}S��^�G�w��z�Ѻ�+0�F��;.J��ଣM�qǗL�'�k/eh����Ю�#�/�J�ĺ��l��F�b��y�@��� �("���0� �l,�!G#,���ٳf͝���c>'�g���z�<ITQ��q�>g��Z��IPR����eC��U���'���f͛<�ϥ���M�O>;q>u���H�����X9eB�
�m��bc%#,���lٳf���c='�g��D�O��T��*�ypc� ܥ���{�Azem���CR���r}96lٳg��챞���QDOR�E�U�|�$ĬR�J�<���٫+*E��H�6}96lٳg��������U��dkQ�|�U\/�b|�
�
xʞ5'����xFY���ٳf͞ϧ��zO��=����1�K~�è/��:k1 �P1�h)"+�=��`�Ƣ�1�V�Q���L�(�0���΋�8����F�P6�Qar�\���b�\@�)�*#(��a��F@ Z��0	$T7;���G���fm�Hd��[R��Pz�No�6s�]�:��:��,���-��Ot�#�E��" �! �}����ɇT�^j�[��W,~��#��:;�O�(<���KGCJ��g'�d����T!��{��[>�~�C�)z6.1����gSҍl:^�^bmfUhq$��rg� �F��0�+�D�yPmF@��z-�vZo�z�Hjx�lIN�R+f�$��ׯ]�vX���g�e?/,��YUb��q8f���e�|H=��O��<tW�7GN�W�؞f���pح�ǃ���@쬘�*����J�׈�w�u}Dc߮+��t�ﱚ3,��jCsL�̩Ӱq� ��_p?�\+��Xbl�0��'p�蛼����;3&Ii�z�c�"�t�ڨ37*[��G`�e���уe��d e[Y�n�����P��G��
�����/���U���gq������$Z��d����٢��lդbۖȅ�RR���s���W�#4堗�YI]2j��ѝ}7=��o�z	��=w�vG������oj��g���+TŊv��ָs�6����V�O��F�0�T������Ʈ��;���?� ��� ���?w���=_��u,L�ǦX+�»�`�ncn��	G�-վ���ֶwM��n{�wSԂ�|$5�D\M�ޯDk㧝[�&yڡU��I	�ݸZ_���nf�Ms��}�0�����F����Վ!X�M�#l��������z��Ovf�l��I�S>��I??}Y�<&h�f�r�a��}�1/^���{=��`��ּ�r'v�]�l��<�^�S���'Yzo�f2����=֑o"+)%T%��И��d{�����c+r�?q�U�h��W���\>���d�\�ؘλ�8sY��s�0��퍦�߽Y��w�p8���B$��Z�U�Kk�'L�����Q�O� �e��k���a��/�Y5K���X�}��f}�9mo���N��fĎ��{�"S�:S�|N�)\�MI�b�Xb���%��s}W�d�|�ެ9<Ō�]�K/�i������r�!�S�}h�B�Jz���4�J�]̺��,����D����>��ͳ��^r촥��΍�^�xtC��ň�]�fd���>�i��;v�`��5sg:�bE&1���L;��JQ�D�!�&�tW�f�UƋ�UB�͹w/3%�֏��@�÷9{ڼ����t�^��^��T�~�G-]v����{d6oRk�ٺ����a�=1�"#�=�ސ1#�rT��T�lֶY�4�;S����xm�����5m��#γ���׹���ce]�cs3�޾��E�yD��C���B����k-��k�B�RY�M�bz6�|���F�[=t��2gג&%�6sY6�����Vc ��Ӏ��mV�a��W�8?*>��O��l�Xx�[�v�]�y
�sM�a��~"�yQ��9�W��>h0Bq�d����v'�2*+}em�Wr�7�/p��u��-S��@Lzg}l� C.3݇��\�S���ƙƸ'<m�d4C3��{p�����U���sW��9&���M��>!F%�����n���0j��J�~���L}#@� �-��}��w����aL�sG:����'���
�%�4ס�8��Me4��XcR��R���A�j�ݓMF��g�&�]��y����l��'^r8ݱ}|��w��/��Ыs&�Ee�]6[��t`֕	-��\���x�!�� y�z�θ=��5�Ŭ�^�~Yw#��[�?{Zj��Z7�7,��ϗ��qO�^����ܤ�0e�C�=j��������j��E�Q�;���l�<��O4����+&-KR�nzx����Pk�~S��5�\����y�8���Ty����>(�����'���5(n̚x�sŢ0n�z��z��v*��sfe0�P8�&��j�#�Q~�j�e�sh�Q{{�K6�F��~��k^�I]>~�9���a�J��U�K�U���w�3��5y�
� �x�5[������`���Z�a��܎�Y+�ڹ��G�׮F�����D�%����2kC��tW�/`�?���o�������;�^��:�:
a�,.��XG/i��}r�_�^<:�Y����o�u\^�8C�Ə{d�K9j�;S�\n;y?5��^e;Eq'��#vFq
7�6�nF2EM�w�1�2͠��A �m�J��D#�=ܪ�;5����E����gns��e�hvvp�z4�{Xo��Q�2���v|<�	d*���=����Ț�4���w�v�ޞ����Z���V�?�[VMu��C��N�|�=������z�MT���J�7��p�R&����1��qK}���=֘������	MBm�Ǿ��H�Q�-���vͧ��ds�Y~�
���y�Y���`X��x�cUP/����jɒ7���*�6*}a��4��s�c����� <���UT�rˆfaPP�~sރ-瘼�WL{L��ꪳB��|#����ŮB�P)� ��73�w^�[uÕ\,>ڍ��w����:ɨ�5�=[�,�Y�ˀ�o�2R���G�n�@�o#b�������C=�(o*�US̆}a�4縊�h�Z��n�	H��Z�[¶9?vu�ˢ3�2m��66�|���ϑ�Y^�����LD���GjΩzH���df�Rߝ��H��8����׉��gq�kP�D�UU��劣�l�������U��k��kk{�׫���ӥ�O�E�p^�@^*�p�&l�6���;����V�Tv�-E�����gt��v���X��
��<�{��6��/3'���T��BHBX5��4t4��{������]O�>5�Ʒ�A�w��~䭎y�:!��st��~k����}�v�EO������ۥk-��	�dQ�u��F1�;�f�۰�y_U�l��F�M��וNg)��Ӟ��l����k�>��������f;�wD���sGd�*�0�����u����/^�:��/":�=�[�|C�L�k�^�7�� �DD>9������H�O�Qf4�B�����^��ک�5o�$���ʏf1��}n�y��Bq�!�}�>1���S�i��[���(�3��_kO{4�r���3��-��A���\o�nu�n�e�UQGCn������$mZ/C�Ƴ��s�]8�S������z� �Coj�5��tƪ��g5(E��B+W����8�+{��*k�r�6)��\~����A���Ӈ7�ԓ)泯(��mYɣ�EN�����}C}�n�ՠ�ӡ�s���L�D�I�[�Ƽ	&�&V��v�xw�q��ڝI]�񅩨U���>��8+-���|ΰ�3텙;�<Sh3����&���R�L��SwM�p����\g/6��MH�8u{m2����Gՙ�Ϋ��H%e	�����|�בx�R�.�c�f\��p�r�Y;\�q��./��V�(�=�b2k-���{Ӯc3
�� {��LH���A?u�Vy�E^�Gg=�25!��#�$�ۺWmyo�3o\h�u�_;�襃]�\cCT]ʷ�R�@��Ql��M��oJ�Ĥ1�fQ�3����3D�����0��YT��9b��	[}2���w1y��.^>�@��k7�k�;SVL�ei��"O_G�|f#6@����I�*���Lq�N�tN&�j֫��m�)��wp���d��������FA���A�w��1��չѸ\_��@6C,X�F`)�u�2-Y���Ss1Sʌ�;�1"<i���=<�6�]np&�VdB*��ɺU��Wm�ɧ��k�n����'��Q��8�`�� ���\�Ǩn�D�(^��v\�/>��M���~P�/2zƩyA����:���W*
��q-k:Sm�*w\鞝]�-�9*�0��M���F�Q>�<�f���T�j�]��_U�`Hg���ש���a4]L�_'v��6��k���F�wl�h���2 �"`�E=�N�z:��yD���3��C�'Z{6�Ϳ�uz�O�|i���zyߘ��偬���
&:�k!��=9������E����	N�D���[U;VsHC�z�J`UӸ�!�s���6*ڴ�����ڗ����̴�=��.ğX�q5 �(��mN�܎�/���Q����f�*|cOz�zOg�5Mr��c}���S݊�l�3�3�oX7<ȝ�g�T��f*^�K�dq�Uqy��a�ީ�^R��]r���̞�ý�y�'%�(9L�
�dV�o-´�i_�`VY�2J�#5���F�jE�,3U��Řޥg��Jӂ�hV6�l^�QK5붚at��(���8-�Y2����"�R�<V�<�}���8Û�T�>�8N^��5��rg�`v�$̴%b�����W��]�k!{���|���zA�3e�N��`!R��x�9&m��5�v^�R�ͯ���U�7�0n�eYmX �O"���Q
|��
�5�e��0���vܴQ>w�n�����;&���Yy���n<�dye�)L�;���z��Ͱ���8�Y�N��d �Á�Z{:�9��*cw5��i�ff�oh+��,5ud�ڭ�UWY��5m�p��jYc�b�� ��I�S���\��Rjq϶���g����
�^l={���/9`�t����>la����*`>�i��W�x���cE�걽u��+����e��%>����-@�-Q-P$[���A�z�q�vQ1�F%M�8fzz}��o�.�9��� �6����ʐ��]���va��F��}j�Z̗��0^��u{���ߟP�,���8e�/S��-���|����"�����4S�;��^Bj'|y���M�9:yܷ�n�4<��9�ʶ��	�Zy�y��/*���*b^���>\m�*d��\��!l[wq}�q�����x�d�����Q�]2�*�W�qmж�z�۫Y�.���u������- ��}�U�O{�Ϻ��(s�	�"��G:�Qf�%g;p`�^>.IDzD�L����G�]�6P��t7����ُ,e[�k$��.v)�:�N�m�=���U5r�p�E"�);�%'(�y�}�{�y��\��ۖo�uYxe33sV�ݥ��xUq�������j���*UQ*�Z�K�>��7�Q�s�rk�a��f�;�lW]3�Kj%��Q��ݜ0v�

S��r{��g��v��s����ٗ��LƑ,�b����������E�d�2v��c��Q.{�/V�m�bp���rO���[�£�*w���j��m��n����=ļ���`��_�8J>*�mխ�+�@{���zݱ�JWIPO��V�I���Φ5B�����`j��d�������}g���Qʛ�\j�]��4�~���H��-��׮X2Y�
]ʸ�;���n=�r��.�gTk��k=����w��eO�XT�޴���76KDV��\���q^22X�k`�<�燜����<���������?r��q�U����������N(��� �
s�z0HtF	��v���@��@�"����� !"�! !��*�J�H�! !  	(��x��@ �� BD�B%�T BUΰ{� BT^��!
$@��!
"@��"@"�!"����@ 0! ���)�$J��!�@�
!��@"u�t"�y��BU �	A A�P B@� �:�q T�U�Q��	E��E�	Q��e����X����X�X��X�q8 ��"������"��(²#H,!
0!=u�t���������������� ��*@��@�s�!�R$ �	�  B�$V$V$V @��q�<��O� �A����:��?�,���|����������P�����O�������������?���_���o���AA��*"
��o��ȁ�?�?���������� ��/������@s����O��_���`s�������UA�)B� (@(QF�V� �Ai)TJh�R�Y�D�V�h�X�bQ�V�ii��bE�X�h�bE�EiH�`�fE�X�ZE�X X�fQ�Q�V�a�b�$Y B� �E�  )V	V�e%�e ZU�XV%YE�VRE�X�b  V$Y`Z�V�X�a	dX�`��bU�VP�heY�FVU�%XH$X�dH`eY�dH`D XeE�$X$ XdX �a%eYdYRQ� �`XYV	ID�`�d�`Y�fU��Q� X%Y�h YeX XdYQ��a�e�d�` &��E�e�`�d�`�eYVI X!ZE� �FT%X�`�b��h�`�`�aI�X�d�iFD�i�d�iU� X�X�h�	B��ZAae��XIE�V�h�`�ZDJDJQ��"F�UOޒ ��E
T�UJ@E)N �p��ڟ��*P"(P
@(�������?��~aA����t�|�<� �
���~������X'�������c��i���¢ ��������~��QDP� ��h~���A��?p���
���Ӂ����0�(P�H_�y�0�>���������߫��Z� ���P��@���~����?P ? ���xp| �
����b� �����?LC�����N��.����=����$���TD|L�����'?�v��A�o���&������l��h"//���������qܟ�����)��C����,�0(���1�_>�)BB�ъBJ�UDQ&��KYU�UIRQJH��@��J��R�(�����	R��JU
�B��i[2��d�VhI&ȴ�Q��ь��-Z�6�ف�a�&��j4�*��*V�Z�љj���Zmhґ��5����ce(������=�mfڶ�m�4�j��SS6²4�mm��kUelZ��KV�U��a,m��j؂�-IVf�+%�FmV�ԵJ�Z��&�H-��m��ZѢ��x  vv���m���nN嶵�¦]���l5B�+T��ji�۪T�4+:W.�jіe�c2�٥.Y֭��Z���XM5�4]n6դ�ն��R�*6ִ�cV1kmZ�ڷ� �BD�
=
�:(P�B�
;q�D=�Y���֭N��Ńp�UUٚ�����[+6�Jev�J@]���v6�K[e�iV��R�v�PE�cZwض*�Z�D�PJȚ��  ,w�j�"it[s*ڵ�mn�;v�����E��ԡU�Zs�+1 �@�U�h��m���A�h��n�ClS6�[j�e�HѬ�[� n�4�-����U��4խL�U��+u N��]���4��.��1JD���b�ց��T��#����1�٬��Hj�Sm�  ��V��Ӫ��b����[mۢ��n��Z�U�n��Z�]2:[kqu̶�j읅tЫ1l����,Ͷ�06���у�  v^��2N�:��J�ΚdR�� � �0  � ��T`��F  �ۀTF��  �[jʵ�J�Fʆ�����x  � ��:  9� �g  
X��  �,�  5:� :V��  �s� 9�`P�ӛlҤ%Zٴ��l(���  �� ��]��� L냠h;�� � :�
 �N]4���  Zr� � �@;8  dS�M4R�kj,�lT�  �^ -�  n��  #0  ���  8Հ hX  ]�  �� ȷ6p ��Z�F��[F�*��(���  � ( {������  �\�  lL  (� 6:� d`  ;8  	�� 
��@4�* d ��a%%HF�4�d��	�&i��~%)P�  "������ڀ 	*ʨ@� �����~���m���~���^�1�7�m~;�C�l&��\���=�o{�����ϝ��
���@?�AQ�r��+��
������_������K���T��V��Sܔ��)
�b̵���k��6�l���Q�ۡ3X�JN���ԳLX���A*jY;�����U	��6�i��,`�6A���nmţ3q*��[������T��Y5����V�Q�S�AY[�%��q�.��4)��J�Fż�y*T$axDN��f��U-fYA��<I��Q�����Q��)P�U�F� �(��1���Gn�E�ʔ,;��Qn��pS.\��4Y(c�at÷;kLw0K�h]�9�&c>t��r��pU�&�F���uG,0�Y*U���l�x2R�(����4 -T@��Q'��H�T�-�O	�]A>��(Kq�����U4V͙��R��Zhd�suK�.�æ�ᣥ< ��_�]F�^˧��tV&��>��\��Et��<���c6��m��x�R2m㘥*E�M��6�Zd�f�ی�ĝ]�2�ۢ,D��%S����gV����؊��86���/]�F��Yunb��i�Z�l$�K݋L��Jxz4z@P�,���X��YV���#��F��,Ӂ)y�l�L�
-�Gr�6n�%����A��j
��D�!.&�f3���d�[Jd�PF�n����:�D%6m� 6��Qk]hŴ�)��`^���W)�rnFӣ(a�w�l�YZ����(i�`Fn��vH[-j�R�A��zeL8Q�cs)���j�;�6�q�u�p�T�*��'x��&���!V2�]�A��Ip�������f�T0���a�� �Jt��[��3j������l&`Ac1���_���&Z؋wO��e,{nk�2��:A��-�����Yy$���*fb�ʊ�I[tB��ZKv����V��S26�@EMc;T�Y�ƫPn��1��-Ye=�,u��*���CT �w��6�Q�K,�'�
�!����j���.�4���L�d:�i]M�ǉ���� �B��n�V)AF��[�i�&[�qd����0�+\�6�1,��z�����Ԡ\�6���62ʶCGB̻:o��70KQ�i!Y Ǆ�Z�� ��NS��;2hM�hd�{`�y�m�̨�h0��L�X�s�ē�+�d�9�S��8-'�W�YI�Yd�x¹�Fu7h��8���K�Ӗ@wX���� �ͺ�wIݠ�,��ne���N�d��-Q��F��ɣf�`f�+F�����hc �i�����^U�b�<[�5�N��!L�FE����h�aSF���>ɒއ�9�0i���e�uv�bU'µQe*�74�mbwy�b�+8��m��9��1�;WiӰ�Л�/��QD�6R�Նf�pkЪ��SJ4��u�t���3U=���u���e�qc����G�%�e��b�:l���Б��jRɖ�¥[���H��Y�Fm9HR�]Ƕ(�jn�eb7�������b��"��4��к"3R��`ռ����8SH�NÉj��Q����]@�`��KG�^����t�I�jS5xo۱Jz�� l�):u/>X@�i틎�����8�M�ţ,��k6�m! �'V��t��n�f�z�
\�֚g���r���1f�XIf�]�����I�d�f5[2�Aֶ�v,-O����f�W�����P�t8���T{u[qM�ؖD�t����rn*�T��P܂+ڷy�C����Ƅ��NӘ4�hMaXǫ7p[P�4ƺD:��
@����m���wE��v#{E�4���8��Z5���3�MB�&�ѻT+*f`�`�@�)+"�L�7m��J�P�X]�w��p��z�Sl4h;�����oz\�����`�٬��m��b:YGɈ��b�f����W� H�^A�ȩڻ�h���[P�!�6e�*᠙m�e��%%�	�%gZ����ECY���1cz_�/mk�A�.Y`h��r䲱�-*i�1^���א��w�Am�v��P{r[ҩ�X��6��I[�0Mh�	�\��9`i�Ә��zF�B�Vq��Ƕ�b��P���"ڏ7E�t(YT�Cub�O6;.���Z QVûR���\(��rAS%���xt8 5��l�xʢ�,`V'�K�L���<�U%�vQ��՟]3�M�1Q����j{���r�2�l�E�A$��WI�XMBF�&#%�0X�qRִ�sI1bݱZ�4�q���#r����qH*ج:�WE�t7B�%�"��#0��V-�Hi<��CnѠ&�鐎��Յzk*R���7���7�Uꥤ������T*H�\mbY�%34�x�Vf��`flZU���lJ^��:]�@��IB�gN��=��M�8�ڥP��f�P
;�S�ٹ�Bic��q��w#N�2l��Fa:Q�	QJ�t�i�5����)�{�Z�Ntb�E/JԱ
i���9��F�*��(B���im�Oj��B!�h�j����m�D�]��1Ӭa��v�mAa���J��&m� aR?E�KD�W��``d�{wa��N�����w����0j��8�:�f����z��� �e�E:z�ۯ\� Y�J�
��h� �B�85o�gN"X	�.�m̩e���0n��d�`���m��8s5�3P�*����݀X�Ɩ��n9�[��yDYi���E�J��R�r�9�A��q����WCiQJ���&�D�[�+��kO
�i����]�p|�-㍵�D�^�iw0K�1:6Yh5D��$w&d�p5�{6�8��/]Ňq̛�FP`����
S f^��H�Nێ��L�0�I�9��6v9!�l�W�y���mŇo+(�R5L5�YZ�T�:��!��I�����u�D�����	�+<�h�ӏk���k�����N�63(G�"	o0�{��okmcḑX��:>�v���c/E��_lA͔SQ�Os��z��X����e�ASKF,��(h��ȯm� X��(e�r��Z�Q�����b�se*�فJ/K֩�pR� m�2&�����}�՗��Z�4Pԩ�q`{��5PX�zU��x��c�Mj�Z��=	wJ򘙁^հȖ�V��6�d_nfQ��r�������xr�K�Y ^�r�F�RS3�1�u�tl�*�������M��:��yE��5i�x��7 *6���Q�[J�B�w `]Ҳ% �ֺ���Ջ]����+-KR4&�#�b����`,�ĻL�jj��Mu�V����B@4/b��ƔK��"�%�*�0L���q,�r�l�Nɫa��
U�ɴ��T-����^ǖ�f��lR1:�ܛ�A��5��wQ� TA@N�D-��ߙ�ӓ",Tt��3Yj�'[������r����1Ǭ]�t�+�(ԽڡGl`2@���LMMX7Q2�(eq
�8	i���D5fjʆ�L����(L����fr �����̖"Г���)֛��(չ�F��jެ��Ui�֫V�r����/��1]��mr�l�]Ҿ�5<ה�e��I��b��'[UW{mƫYn�x����4����w�4Y�qG4�.�x�ÂKF�eM�-�Z�5�g+M"t�e��g��Z�XyW�<
A��f�R	���F���w%D�L��gtEc^�k6�����"��1x��X`3���4*�M����5lV�%x�J��a ��F���&��L�����L�ܶ4�Yg5*�ef�K2a��0�E�We�n�u4/�H���Fij�L�\���W���ƅ���5YT�JX�2IS ��i�v&h��[xw]7����x��-�YWOuA*D�/�m��a��(�n�H-���9y,,8rDF�b�Rxt��^԰LŐ�M����n!Xa#uC����36u��(��=�Z��Nn���I�$6���y�L�fc��%�+%m�,�A����6�M��,��X�4�$����q��s(������nVJq]���R���2�1���V$����ʓj��SDƢۋ)&�$7�0��&ӛ*�}�%�%�*
���fZ�7���7bחKf7�%YP#^Lؖ���$0L�� /	��1����e�܈�2���FY��,"�U;M)BE�F^Ӳ�y!
�=��d���GxLA	b�����Ɔ�J���e�^%L�v2<v�*\M�5�e��Ŋbη�H��c��,�	i��3,�<m�:Ku�
�k��z@��M�d��,)��V.���U���3MZ�l����`�% <��*͡t�&\N�TwK6�X�(��woQ�E�Y�3C52Y�o2�P6���^��F����Ņ+2RiA�âH�����G� Ɇ�e^0S"�8�6j�٠�S�r�,�Vx=+4V%]\̡YJR�A6��v�Q
23�74�9�>Ő�O����̑P[vO$ځmԭ,��/j���k��i"���mG2k�6+�//�ǰ�X�HO.P{m�9���'��,�d<��1�p=
m�c=�n��&"���0��bm�ybS��i�3��bڲޥn$M�y�T�=��w(�%<o5ϰ��"���P��0��t�DYIe u)V��j�i��Y��6�a��Sdkh\lJJ��-�r�D&��i�����& ��	+UrԲ�� �F�����f!Z2;q���R쒆�w"�"֬'[��gr�Swfcl���oM��t�%0�=�GӳAeժ8�-VwJ���6	ո�Xe+rLo�I�fn�T����V���^Z���H7Sa)�VA�#�q�ΰX���S[��a8���Z,��-lVCM�$V��̦�H�6� 1Qz�����C	���.�^'��y�{.F�;rk�n��^�X�����!3HK�qX�,-7錇[��`&� ���7YJ��w�P��suf��*��&/d�飺�Ѳ�E^[�U��cIIF�R�iȶTV����5-mp��];g�ԯ>M�l*ʺ	1Ee����ZRV�a�>��/I����fU�W#Z��>�a%�� �÷`n�U�ؕ�*՜u���
hkZVe�t v�&X���-_&�ktZ�Em[Ucd�m�+���;�xt-2�8��"�6Ukh^]�$襹�$��Y�Ğ
,͇qaR{`�3Pܩ��X�E��e:����E�b�:��j�YZ����<+G˽y	��Z�)�أ��E-Y*��m�q�ݠ�%���Q��}�c��f�	ޡ��V����٧[ˣ�+j��-3�ؒ�ӣ)q�F�JZ�.��YW�+M�x͸0^�m5z�k���1������eY7�Q7X�&sEH˼��d9.lZDS^����ug�oT�p&��ōe�3V�c�cmUު�v�m���"d�ݻ��9��6�"J��I\36;2��Y[)��Rx̌:�.��x h�F*�ݭE��&�Mr[�X�ܥx�6��]F�;&�k2<T �+�%�	�I�a'M&�9(�e��B������A�/.��M*@0a�&T4V��t�]��:cj�M�y��Œ�Eb����G7Q�7��t��"��m	4��`B"�ʛ�w�୥Ȱ��wZ�Vu�J=k-�2[ }4o%�#�9d�M3��K4B�Î)y�(�&M-j?9h��
�!R��V�*�N�j��C
�k*ܱI"m�њ�q��l�E�m��J��(݁��W+s�I5��N��ɿYP:�fJ`Ì���C������pS/FL�0W�*�͍�B�`-��s!n&sv��yu�h쏡/
E���B�F�o(�{��j%#@�ŉZJ���G%�T��i�VQ���te�dm*�Щ�hx^��j��ʌ)%"M���#b:�.�� ;�Vm^1��kV��.���E��a8���c��Z	m9��Sr�ۚ,S۠�GR2�0�B�J��#����7�5���$�B��z-�B���d��P[�����=�;N��Z��55j��W�wKyC.�i�v�Vք�ډ�!q�ݭ��=���*� YL^V�V�lA1�̴-7��3�@2�����II�N��D<י�E��Ӻvb���1�WX7�y%d�j
��&\����Z��j'��i[v�
":�����F��ę�]c)25PSH(bY�,��U/s[[gV]i���X���3E�tF"�Y��BA����uLhETk�e�V َE31m����*�D�#���X)��E��M5X�L�B����fP���mǈ'������i�V��.�0e��㢐 &�͇r�Y&/��2�ʸ���;*D嚳qV��˕d��[t�����EX��+ �n^�T_[�0e恻%1r�s�XL?j�ed�0�ۡ�[�,'U��Yt
JT�+yJ��j�m�Y��7���F� �i	n՗�KU`�c�t4벲�nmF\MӸ�껋t9"yrĤ#q��Ň2�n�6$�G]5H�a#��&�ܺEk)�t�S.�t'1T���y�M����t��rf^ 1f�,
-CR�ͤq`�h�`�#)���n%��[W�̼Ȧ���be�9j�Y�$=$~�Xq�N�W糗bm��K5�T�c����&(i_���q��K1��=B��V��Ř�"�N۴���B�^���'�Os�KZp�j�U^��F�7y4�Fj۷3[�h�6P{Ud<ڸh�oJ�J]=� (L��ü��Op;$3���0"։h���ⱸӧgi��7#��0QM-�[�kj 츱�e�1q�v��/1C^0�ӏlҙj�L����&T�s�"Y��6�I�N��*�B�
���8xf��>T�ؕ;aV�(V�;��sM��A�C���F(N�����&����_{'R�R��<���NV�5�1%�R>�-
л^'t:�6�4���M�e��\���;&�Z���ےuoyKߛY2�E��s��@_���9�|uQ�<�ď,`h�)/}CF':�O�U��wONE^C���0�9��홢T6�M�����A.�Zk02�
K6�f�C(U�*�|�^<���-7�RVA�8�����U��ν�7$�%�mP����nSrw��v�L��+��YO��������0e-����:�����K��9�3v�vMmVЬ�&M2�Ԝ���i���h}�V�Ļ��5KȳF�з����
v�d�j�{�l��Q;��x��Z���U���"�]�Vf����V��=xZ�:�)�V.�#�$Y�tyr���4�k����e�j-��,<h�1�ܺ/���✭1�la��)�ӽK8)K.�0���B��Kc]X���7H�tX�=�[��;�v�D���(OX���?-+R��<������:��3�e�E�6�����3B��t�m���۹�5GA�Yp(9��[z��_f l�D�\���Ԧު-T]��7��c�m}�!�<"3F⠮��(��wyn��J�<P9�/bC;�ZSD ��Ke��c?B�CSKC{�Q��]�"Oss^L��ҠE��3��3S5EyE��͞��f�]w$K��yS%6�y�D�`�a�����j�����:�
���0�[-.7����o�"�S�78١�+mY_f]t�k��//��ׁ+��$�ŕw�zk�: �>#�I��j��f���������y���q��Q͛\#Y�;`3׼��%J�_gN��aC��j�=��akDʮz���x��oy^��|������t���{O��7.�	E���[ǆ0`���qY�z�C.R�a2��sw����y�m{(SFp���t�7���?7&��n�ˑ��0k��(�Kψ�m1�q��1�n�8���G&�kR�Tǃx��#9�ˋw�㾲�������4	%�J�m�y�=v�7���V%��K�M���v��W4�bn�@�6���v�{�����6�3���>�\��y-����lkT������ѽP�}�[�p�}�vm-��܁���4��V@�䐖��kt4U��G;[72��fls\���ٮ�G2���[��-�&��KeL��;�O61�ݪA.�b��)�h� N�5�v(�a�x��iL�n��	Ws]��7���ٗʍf��y;1���,�>H��ȕ���{Y+�PM�AGԻo������RdYjma��*�s9j��8��Ș��?�]	��$;��G��*���$��S�iv���-��"��,�����Ҙ'^r���R�F~��N��p�v��G��J{)u�8���[Q�.��$�:�w)�v��|����u�� ��;�$�곊K�l��U��2к���&�)���^'�8�ګ+��\3+�elZBӫvGrkއ��8c�`���d$�\�c��r7�2��6�������s�8צ$\����İf�3sh��jv���o��]c;	h=�T3N�+�<|��F�C�8�ag��}<����&!��$�[wl���҇U���tﭸ��
��f��Qvj��2����y= ���u�;�֥��CrXF�J�����$;���=S9z]��@�i�:Adl�tL�G:HY-�������H�֔�;��{.>n��є�(��@q�-�ly�L].�~8%x�[�\���'wj�OCA�&�LXG�Ǡމ���-�X�Y,.$)�Uu�����U�U�P� �'�&�C}K�ٰc�;�n]���RKu��f�rỚ���z��Hmḓ���ī�B'S����iݚ��h�W���
͝x���n!x{:޵s�txV�6hN���1OB�+�,�Nr�unP��o��ƙ�BOʋ멐�62P<��8��is�WA�|Y����o�ᒶ�P�:�u�*�)l[WQ��*�0�1Dr]������y�; K4�`�羴M�ݺI�� Bg�w�L�f�3X�9��D�)wnz����Ӏz�ʗң�����jNIF�L J�N�'�]٫n>��yyV�1�&|Z��-�{mԘ�w�$zw�U��������L�r���ϵo���ud<{�V2�pa@mtf����؂�nnnP)��6�����y.Y�h�d��d�ٗ�M���D8�>a̼%�z�&q��3#�C7�X��qn)���xT��i��]�����F���j"o,���ޱ�f��� �������Q1��:O+��1t�ۋn+����[��-��|4���Ҧ>����4)n�(R\��b𲆛���yJ���}b}G.C���鎚�:fZg���9L�(�0G�:�ow�6�un��B���o��Ԅ,�EX5D/'ҲD�!E�7;�s����YVp�^^b5kE1�ʹWhCF�\b��+ u���=V�{{��.H�4�\V��Ź.����tȃ6�kY��Y����{��[�(��9�z���*yt8�wbn�T��vd�ĳ�\'G��j05wC ���;Q�
<*4wI��庺��K����]M���Fbc����Y�ܢ�7b���\�s�th�\��������Psw�\&%���`�mE��9�bDj␹d(��u4IKն+���J��9M :�ݩ��WZz�vX����(�y�Yˁ���E쾔�\@�̪WH}�g��{TQ�7#�=��\+��<-��o�v=��m�%+ǁ�i�|6][��X���KmP9c��F>�:Uiw+SC��y=.�B�z�/�g�@�4�������|2Y���ƛ���R;�`[�:�����u���/��(6k/T��b"m�Em��%d��}/�؏�Wa����N[�2��p��f�#.Ȼa�����#Fp�B�� �ٕ}î�jīu,��LB�rс#Th|�V�ܯj��I]�\��/nccRU�+�:���XЩ�nVٻ`�}��6�6K�-(�9Zg0VC��(<��
A̛�%i�9�	��N���Y� �ԥ�'��4ќ�2�AG�u�5�e��źke�$��p��0Q+{��Wmn�q�#��z΢��V��˭೪V�`&�_'o))�B�s�=�}�B�ۡq*�otZ��mV�O���uK�=�=�	J2�"R2��ˊ�����ur[w2J�;���D7��5����a�X(V�@��0��q9�z1�a�W�c�ג�zw$Ma��D0 �A��*�w�A����r���y��-;5{�j�Q⋖�wj�M1�PJ�oP�n)�S7M��Nw�9�.�z1�*]v*C�������'�(�]'ZW[��"��ge,�b�蕌�-�d]6�X�U
��������Uz�BG���^_�!���U/%�m��'.���\��=��D��f&x�ǁ�l����Ƕ�;7�v��vt��Z��
��7K�[Eo7ivK�*���r���5��LqXB���+����V�LM��Mc��u��ۼ��x֞c�!�S��gN�[ar=�S�<]��gRؘMZ�Ҏ��/����Q4[x'V,���0�ڻ��d�v�X�CM��֣�����D�f���T.ٶ*ճx����̧ϷԖr��/�7w[�Qċ���ݪ}�r�����T�U�۴��욤�F�XyI��p-�歙��n���Y�c��7�G�y<��nf-�B��=у��3�7�M���5l{���\SxN�lf��r���,Y�|�sd���FvwӲε3m��v*K�0YE#@_*jz��0��fO��u�R���rE=u36���a�����b<��/ke��`��+]�%KPV��@�ᡶfR��gE[6_:c;f$��N\�`
�C.��vZ4Ci�&��yQ+�!���H,�h�Y2S.��c��p
�WtO���h����|���6�y�����vXݕ
�>�h��AE����C�a۩yR�Z����*W1�rc-'1Wa�{ܦ�[bz&0f.89�p]r�Q�P�?ӆ��hf<�Hv7�m����jJ�1�z�|5����@ �P� Y�@\�6i.��Ǵ,s��Q��wػ�d�Z	�>�sv��������.Q��9 �� ����`�b�琺'0�H����އ^���B,�÷��P�4�Ñ��T�(��O��@�v#��:���H6��8�����R�7�3N<�ҿd��ƙ��\p@;rI=��*ע�`;(�w�[��_���<%IE�	�uU���u�s6�Gմ�[����s)�sjk�.��}ZzP	�Ŗn�vM�TÒ�	�%���EE@����Lk��AkU'*��V�9v!7��.�Ɗ�3�բ��ӊ`�zC>�8����u��<�ϡ��Sk�^�V!σ�)��V����ōL&vCqX�o�����mHm��dB������3�\tP���♒������m�����S��L��ta�~cG�����y����A�Ǭ�'��6�m��z�8X� ��W	��I�*�}�3IB�Nr�K��M\9yI<�L�ϭڮX�wj��emVʵ��
$�ProIȯ�s�^}ܥ�T���׎��H��2r�7�+Rjb]I�ТV����u�ǜ�jƌ���0%:��]Ia��CU	2PǍ��ԋS�O \��$p�w�"�9f��H+���V��[���-����Ч[ʷ�i����7�j�� ��es��<_8��UC���t�Z�u�E}8hwYO@��V�ә���R�|Ŵ%�w�`u ��'��.�3�J.��td��y�j��-�9aX�tǎ�[��(�vX�m�)��±��܆'{ҝp���*�hfg�:竵+��7��֠1l��/�v���˵4��`\��Z/���A���f���r̠/�d܎*�
��140�����X�8�e�k�Ĩdc��(�]���R�5��Z�B��&�Ƿ
SsWZ�+*r�"P�Mt��2+-n��:q�o�1tw�qd@^��Q�86��}���5����(R��2�m��'N	�͔�̫���FT��'�\��9��Q��������9��c%�o��v^����/;�d���޾%F1�ni�i\mj��8�� �)����^RΕ9n����1��J7N�Z���`+���}M_P���@�Lc������h��Y���T������W�X�Lke<R���-im�/��e���2�W͓��aW�M�f�GH#u���gI�K�]63FVC��`�n�bݚ�ՙڕu�˨���,���ٮC�^�ʚr;\SLW�k���;�[�4Au��&p�ŝ��32�<�-ق�r��_-e�˛[Z��Z�w=��iV�$����}v���lw� �vyx����������ptH㹺��d��峡�9���3m�|+� �����;֩>7�_yyu���*R��q%K�2���L�Q�9{����']�ݕ���2���V�\+�`���T�L��<�[�؇��U9z�=2#��J�zFm�}�h+�t_r�`ī�Fnk�pv�&=�4΃Խ��V��\��=�6,U��OM^����].��S����&Z�m��5���4�M��B}�b�+�MX:62���{~��<�Pަ�93o���e�k1Ү�䭪|�:����nkXudF+2��%�ZD�k}��1�.Tl��}<A���6���}��y�_z��=ݚ_+<�ӌ��]i`�r�),r�;j=yh����V��>z�̢j��xz����o� ��G���iHmL�%_<[N��ȭܭ�h�*r���������:�I�a�h�d���&Sj���ז��+���r�jl�%,j�:N��Q��z�Ч��1�S�L�jK��w+��ru�ʸZ��0����c�Eޫ��� �g�v�Q6/b�!]V����n�Μ�f3 ��Ր�(���C�v�j���=�W�`̱�:A`�r��f��w��_a�<d4vȕc��I��T�֢tL��Od]IKZQ��ޡ�YI�ى��Y�x�5�Ɩ(T�fR��u�VpdK�/
��w�{N��v��+�C�����9*.B�09`[ru�ۦS��k��!y�oY6����iU�
u���:h�\��Y�%��D]AR��s��c޺:x��)�߷.�z�����0*� f �i�u199E�}p�\�YK�1X�2��ڛ�d������T��h��&M�&�;]`G4{�%:dG=|�Zт����&���\DV��*,a�6f"z�k�l$�w+:Q�S1�9�R�[�I�Yp�m��'o;�7�o��ıoԯpμ<Y.K1]��Ɔz��w�4μ��ؠ�i�f��&^	�؄��:8��*�Vv42���WkmoVe=�J��Gkv�lǦD3.�f���Ի�sL[��g>h�r�dyZm�ϕ��В!�����h.^.�,�v�k�5�#%S��7j}b�Ԭ9�	k��hq4����@�B+r�y�g�y�`�/�<��>�Ο�i�}�����}��Tah^v^ E};r�}����c�mθGm�m�X3y ���>��0*Ř��=�s�������|]V����]�I-g]]�g[��~w�7��]&�
��g�S=�u��KY۷��uSF,���k~�x9���sS�������+����2-���N��e���^�[��C���MR�v��&)�`�����)(��E>�W��Ǫ褄k��%m�܉؃�ٛ�o *���+��=����Ǯ����z�׿���#��_�.ɋSnm�d11�fo0�}ׄ�Z�[�WEi��nƌa��_ ��GK��n$�r�݉�o=5�5s�;��ΨI���Dfms��U��.�#��]�K��DN�X�*��	�w^aF��yzl�ky.=ڛ=v̙��B�*����/��)=��`8�\wk0��F�
I�c�y�E��7n�{_p��UǱ���:�������ZA��s%
 %�^��v˝�Q�uu+`�n��؆"n�1��)������w���9\u|4 �c`��&}Ոu�Sq��]��K#�ޭ�wR���i|'������o{e����m�כك�$0�1`O: ��+�Kb�4�Zo
� 7nO��[��NUۡ*�H���<�?��Mr�K^N G8���<�����2�9�6� �� 8�YE6��ػ��s|t+Gh˵�
�<8���l�]@�Uz�%vmE�tbm:D���M��k%ś� �(E�dV8�%�+n�2��e^�����Ge�Z,V����@ʅ0�@���{�)[u�$Δ���yK�r�5$$ab+����1Pa���5;ǯ��{n�bSԠʉg
�|��g.j���ͫ
T˳��4���֪ga�oRaWۢ1�)Q���2�Q�slRݶ��* BזmjZ�J�ؼHۢ��l$n��B�t�%fe��Ɲ���g�2gU���n�V5),�tY��ynV�R�d���g{b��I]^i��\^�J��i�g�޼���U֝�& �6��Y֠<Ыub�� �A$:�룅�-R	nл�zx:v���@E�q��P��.�|���[)���.+}��������@�϶��"[�����e��΢��H�r�de��$Nַp\DwŌW�r�Z�L"�\`
�h���c��Q��]�0��m��:w��e<�f��:��[�b��Fu��e�mo�1�9�O�ɕ�9��,�S������w�Ɠ���H8�
�j�
�f%���Ռ��N��bt��Q�oC��M��mfQ�.�=������;S��F�5��Ry�n���Z�KZM��ڙ�Xɛ��wSv���V�P�[�S�]�����Ȁ�]�u��]@��ɏ�.��wἐͶ�b��̌m`Yu."�e0vF+�*��!�e�j�Ql��N8�S����j��ȕ���Ж�w\����򹡻�Z�W����ޚ2e�y��Z��o`<����Y���V����;sK�_J��ppUOt�H�۽OR�C��U��[��N�Uv]���<��p��\�2�+W0�еe�jlty[�9�v�OH��P$�[!u�U�M#���⁻��p���Utі�سM�]Z�����S�;�� Y���5ܲ�i�Q�6�I�t@�P������ϳ������I�D��@t7�)��-w���z_W-��n�R��{g�.�}絘=_-0}�-�g����Vi��ޓ)
�p����T[Y�KCMK���⫩Y�Kmebu��G�qݥ+E���PiT-�d��js������ZM�x��µN�׮��?�R��
�k�k� �C9�cqd�1�*m|��+�֎�;F��keY�ݝ��*T}� �wU-�2鯰�z��\v��%b"��OT��\D%;v
g���x�15�D��*	��"���Սsø�"Aê��jQS8r���C��%�@n ���\��}]>��~j����tH;��7����mXR���J��l��ޱ����Łiݷ8��֬�:$W�>6����s����#�Z"�nͮ�D+��g	���5N�:]Xr� �����u�i*ܫ,�;��6�.��;u��ř1dU��9��2�V�М�j'��2��˘�Eq|K�y�ȍf��T����gS�i�zK�}��M4���1:���� �0l�-1pU8$�,�'V�%-�$(���JG���n����vLQ���h�+�	0&N�j�)�����if'��AIa$ X�S]�pv���RDw%�ٳp��%��[J��Ly�c��y{B�j��Rw}h��Z��4o*��P�4e�T�6l��\6h��z�NV�b�`����Xچ�ۨ�h"��OZXw�].�����������/]�J��g�Ռ,Jl���q��}�o*�"��^��}�h�'�]N��
PS=2��=(8yR�.e�wݝ,<�M�F�m��.<+q��j�%�4H�=�V���Uڭ�$�������bS����*q��dA#�I�ٝV���s֍�pѸ����~�V<2[�j�1+����T6u����5tv��G5���1���p���/�#��흫���-��n���j%L�مuO��Aǒ��3
��̳BrY��.��R�E���"W0�8���f�8�ȲwFsbڈ���k�<\�4ٴ�UЙf[��uvǚ��*�����pq�x��������'����:���ζ�=��)����]=�4}"�Ϛ9�E��l��b-�wr��f�|��l�vaY&���`'�p��c>����{�\� i[Z�X��VN���8�6��)Y������S-�G)�@ۼ��&�JU��to��{\s�f�1R���U�,�����ɽv����]^�K,&Պ�7tE�6*;#�1��ʀ���F{T����D�w8N��oi��2�SCWTa&�Qӕc,\�a�2�IH�ozmk��[Ƣ���8��`�v�B�D(�:��З��0N�j
U�_��-�6��VZ��y���-A��n����^�(�%���'n�3ræ��ވ�u���ɺ�O����Zy�Mh�܌�:��X�l�xȗM�Hf��pM�ҷ��3,7��*�9�*>U�z�yw�n���`ff,��XB��%#P��2�SE�l�8QE;j.�͠��2���w�`�;��V�g:J4�`T=#��ռ�y�K��ڕ�r���ϳ��Z�q�꽈ћn�g'6�f�"�M{���R��绽��n��N�M�1D�]�û'����Jx�Ŕ"�3�b��ω��;�z���^1w����r���5j�&�S�X��8�fh�p��d��VR�<�#�i�kg\\����;Q"lb�3UX��������)�wU�)�Jx��7t+>�{�3IӆA�&2&����o����W.}����[����Rw�J�x�
7HH�gM<oaY�%~�ܦ�&̆�Ǿ�R�PE���wV�SY�d�S1�N�e�` ��+��Ѝ�<B�q�݈+쉵�;�b܀�� ��ٖ�T�&�Jl��3�m��Z�e`hmƵna���l����Pp��u��K睽��;[V�~��0{����}��q�E����f�qf��`Rg��x�pV����5���Y�-;��`y��}���7R��-3(�Q�+�����XX3K�Ъ�c�XF��*o���k!^p�7I\����U���Y�\��Z7���4&Zr�D�Q�+���lF(���Ʈ�-�m��{�O
Ct5AĈC*]�u��x>ͻ���F���G3�Rq��}���U���!_�@�l�{5<���-�ܟQ�o�z�d����PMy���n�}��C�S}m����8ޖo�n����7��fl���ܻ����؍$��<��^�K����'[m��+FU��@i���j6��X*p�����������(��̀�ݨ����ݣ'��v� mLb4��n�;����\6�X��4�X���l�bU;T�Md��V�5�g��%w`����t�ͷ��t�+|�� U59�o:��eX�zuq�u;�I�)ܥ���CkL����tE=f�,��Ν�к�7o�l�\v�m�U��Ք�#L���u�7x�^��
p����Ԋ6A9eU�-��/��j��z��+Gfph�F�k�ef
t��d�wd�Mx�d��CH+A�����y�^�O�sN>�2�0J�׳LD���i��V)��4H���ZL����Gf�{��oV[q<T[;t)�s�i���Ze>�Qš�al��uebŎ��RN�j�J����˥򆥜��}N\���p��l��b 6��á�B���g5�݇�l�
�����9*�jY�wR�,?)}Q#F�Ί����C�ȅv)l].���-R ;B�n�[O���o���/uGL�'�WWcA.ڒi�.�ܳ���H�x#�pY�MS�On%��6�Dpxx�;���bO{o�2,�dhz⛝2��y^�<���$+^]����q\il�U���ar�<ӕ�R� ��wF �hG�n�&;�������qv�c7�ɀe��o�5��oN;��aK�%;D8d]�-�f)�:{+Eډ9�@S��_p�ҏb���Ѯ�o�SyMƥ��GW3R=��ܬ�4��L<ܖ��N��a��۳�uw.�]w��F7�uɛ"����WN��%0$��z�^��j,��JsFX�Shfr$�|�J�G��U�Qu�!b4�E���nu[�$y/�2�1
��FG���X!��1�O\
p&�2���}��.���V��(�\�e�oV��:�g���	yj�d��/]:,�[6���J�H��-d�5s������n�!��SyV�zƧ��4؁�q�Y�ur�q.y��	ZJ��oKl�Р�3���[�(
H :�,$���B��N�ݬM8>e+��:�{f|C�ʳ�vm��,	Q���1sa+�d��2�gl�,��m��ī�h_I�NÒ{�n]Ņ�P=�ש�
4x��3͵�]�a�]�m^�#���ȶ���x;�SZ���hh� r��[_���]U���%�Q��!��3���kf0��+XsU�����k�勸͕�|2�e��a�Rw1�'=+k�_�zpw�|�9u��!b7�"���j����������{kj�{o|oh����*~�n^�E�:�u���a�]{�zk��J�H9�Q�9��:��[�gi�i5�b�Ѭ��ƭ��]$\\���
���"��/4"mdW��@eI�OEE]��)*թЧ����];��P���	ƺ��f��ʬf7��jpPTP��]w%��ۆ�J�g[WQ�÷bc�!b�죘8��S}��kZ:���Hfp�<(tS�z��\|����O��Z
�0F���9���V�[����d�xa@K��Y��Cu������kS�7:6�֊�k���oh<Ӈ��{��� ��Q�e%�;����C)Ky��f��)*�U ��Ƚ5nrX�����#��yȼ��2������+��_b� ��rC9.�P�{qe�.�uy��JN��:tk[/bN���!i�ՅQ��V�]o�IZ����<��X��ܡ��buz�[��T�B{��.��>�Y��,���,C��&��k�@$/}3���a���]j�sܷ�r����a�0�=�iݣ�p���p�R�&WΦ��� mfΔ)�:o/H���1�mV8^�V��ͮ��W��|���.n�ݏk	��j7�rKB�20�ݗ֮���яjw�sˈ��g7�6���!$)Q1��r�.��P+��W#od��,�v&l����C�R��2��L���]LR����b�*����o���:J��.4���wmt��5m����,�|T��	���{א
�E�2�h<�Sw;WT���c8�n����֑�V�����T�rQ*�<��ܠ6�w���aP�K�Q����x��x+�R�|��wpI9�o��O�+w�������6Z�uma��x0 ��>���u�g���7���eK�owい��̋)�4F��5c�����4�u����72�V+319���	>5{O�Qߘ���U+���c�$��0���q�r�W-|��z����%�5��>6v�}�	TV��+7��"ǻ�NG��][��DY�֐��Wz� /����%�%��x�se5��s�Y)��T���ԥA]f����l@a���]�v���h�%Ǎ�l��;X�v� �kvmDa�	���]ny�-dNiY��fV8jZH[Cs����{Js�O-��i�7;S��pb-�
���|���Ѵ�4��K�6H��@joDE�x�PJ�;惙u�
�'*�|����I\[=��EL���WK���5��Ik|;e.�;,�ؘ�%��Qy��T9W>�̜�ΙB�-E�9�uk˩gf�=�t�5��]�{E+;�/W«�Ԧ����Jt�\hmՑ	�~p[�d*xPN��ޒU��^�Ł���(Lǯ��ե�(�����z�Ŗ������ʻ5d�x�f`�P.�:�E�}��o*vhSO-\,|Gik%d�u�Ҵm�[Ou��Ը�hx����O�y&�;Ҕ}qiU)���0�Ĝ�w��q�jb�/�*�ٞt��s���&{u.�B�oO91S�k����\F�/L���9q0���/���o����X�����x�A8����i��p�S�WW9+g��(�o���%��y�Ѹ��}n �R��{w������	�{��$>�+�6=�,F{��ס�[�ꉸ\s�步]�V���4/0_lU)r�j��>1SqgJP �>Z���+�sbc5WG�}�������pf���\�IOUjG����%�n�2����u'�6V:E�˶ :�d�G:�qQ�䡮�7io.�z򑬋Y�9�g���61�j�rh%qn�@�Ո��Y.�хd����t/~L���M����ہ�7���o{������v��;g��*�&��C\1�+���6�p޼vwY;8r��T��f.�¹�)X/z_fQ[��y���"�p�U���tՠE|�}�Xj��
[|���tU:����w},��j���l�ls����Q$s@�$mk+VR��Z�y��a�XB$d�il��z��</]�{e�,ꒅ�u	;��@{7���>ٛȮL;�'p 2ܤ�.���J�P��H��JF�L�F��a�xT6���1��m�e�DYTe	�ԝ�I��ﱆ%�E����n�cSص`��`-d���	v��ƍe_[�А��&���hc˫��:��(ְ���=�<�Nc1lB�VN|/�t��f_ �K��E���{�	i���;�.� ����x��ܨ$��b���es��z��)L=�w�f�jb�SQ;��z��0]��y��j���I�s�7��������r�%�Ɗ��¡��.��`ʨer�7�Tt-�*2 ��Ğp���4S�I�o8�]��jzO��oOi"����# `�4��\M�������҃�Ԛyx�@\gw
��w�
��&��}�Y��}�վܷR��t�WZ��=��r+\=V2nT��Fi�׹dl�O 14�:��]�;�)�ڐ1��j�!_u�N��^��ű�,[5���W9e�s�m���ۖ�)?�=Qm��B�Ѡ�tn�J�5ݺF�Bhh�j�LU��]MUlPt�@WE:M8��@R:Z]Rm�R[]a��z7cE�	Ć���`��nƐ��A�
:x�ݬ��(�:�j���5ӻДj���{����)ѤНwa�[!ѭF�-V��K��n��:��Iѭj���J"=�]d4�N�����a������Ӡ�i)�8������SmEM�4��hlj�x��N�.�t�{d�5F��ۣ�C���ɻ��-q�tu�h�kUO]W�+�
������J�Gl���z_>����?�7�%�Gz�*��+|�+�6Vn��n�M�4(�{$�i��� ��¯����ĝ�7j���&1����`�n.���˪��;GL4�.���,�bZ��5��h��1`(���t3٣[RKuɫ��&`� ���<��.ϻ���k�#�"Ǡ_F򠻮����LC�a*N����FJ�p-e
 �� U�ȩOX����7>������Y��c�j��Y�j���+�;,|Yc��c"� �� !i`O�X�-w[�2�����o6���'�i��m������F���R�N�vg�t��ڞ��i]O+4J����\Y��9������U�GK2�z�+âŅe����p�O��
�Lٰ�(�?��6깰�[�w�k���)t^���=W�k�GY�^۷�χ /���9�_��氲R�nE�,�$�Ï�K4��)e��u��/��ê������~0u���n�<�����VP��m��e@E�b�����8a��`�DАqD`�Ϛ�4��~"�;=YO��T�}�P[��m��m�s5�7�]��8�R������-yk�=k�zy�$E6��LB�*�0`��\E���y5��{沴Z��7 �%mc2D8n�=�%�Uc&�ss=���Y}�-n��[P�v�[6ݦ�୞��n��;.[r?q3 ��0Ƨ5�l�͘�]����8�Y�Z��r$��{OM^pwyG_cN��rs\8�fW�M���\h�	'�4ڝa�*��8�
��/2�_@7����E�G�\���O�V��Ǽ�ﻝx �[�K^�N���V�f�v��J�B�r�ρ֞���s\���O�ǽ���������7r�V����[���3yh�^�E��I꒝j�0I�2�wr��.(�	n��JȘ�_gZ��Ln/\�(��X��W:���'���]9͜����w�ݮ�̎�����#|���J�d�c��R��SK��1;Gw$Z��tQ%Y�q�E�I5��NC6�.!�T:@3����ɾ5�������r뇯��9k�y.��9��z�;[6�����]��b8�0V��[P��,���cfv�&�-�V�+�U
r��uSS6�吤Z٬�P͏���jq��.#�P�`��0�B|�j�#=���p��b�n��5AZB�VW1����;hAڱ�!>&t��dJ�mQ�����"���t@OzA;f��匿E�����k��g�R�C�<뻡���jU���Y^�->�͘p����-&#M���)��h�r�;�ݜV]*>�.z�=>bG%�YׁE���"�=���9���xn�P2z���-X﯀�7Q��6�'k"yɭ+��=Ʀ.ɴ����C�]��O��޼����.q�\��܂�6��V����m�
P�6��U��Xj}��q��-y�5�x�㺣�鎫\>���V;�������!�D�\+���v�Xz���±�y�#���Vc�V�S�k}ǭ➢���]�,��*3%����'q>�ʵ�ڮ���ΙƬWq�y۰v�~�dW�I4�-�El���S�@����V�k�]����<t-O>ğ�fJ����-�\�~3�j��Oo�:�&�s�A���3վ��[�,J�J�D�o�1�{M1=��־]����]��<�������][s��1Vz�̽R����T�U�^��üv�.�<�øց9x]늹�E��Ѻ�[�-��*��Ks� j�>Mr����t4!}��wr����	,6�P�������Si��fV��8Y�:C��q����O8*|*qН��#)\�R�Q�O{}�Xŋۚ�k��X+B��ۮ�������F�T�v�t��:8C��x���2�LL�B�
�6�����|v���<�*�~���Z~d�{��]v�D�]�;گ��@�C>~�U��*�w��+�a���3�y;�d�}bM�����}�jD�9%]`I��2|q�¶�ˣ���5��W�`ٔSt%M�<��k�7u�\8t��jΜ4!��do��˙��l���}p��n
�.dXbz�!4�����^��)�����{�O�'�!Pƶ�V���_>EP�@qB�w���?l��vxRx��B=�Dx �ڜK�Al��j^��m�ww!�}@�v�S\���P�Z��%u�"�Պ*�w����}�V�6�Lڤ�DеDP}ǁz����q�Q��n/1!M=E��Ώ�.��z��ťY��{]v�W����͐6Ӻ+�\PhJ�D�Z�.Z��
�(]��e�٤��i�VnAS���B��|�ZxJ����7o��GV��Y�\@�;戮�z��}�XV���oW:���s�1S���Lh{&F�L�]Y�f�3)�e>�%��eOR��� ��6�{r������e�%~2��
�3��_���}�o�ߘ^h�S/�`�<�g�����������N���.���$o��ԸS�L>P�{�>��i��QpZ�(ЁS�B�d�I�}�x�7��j�^�*�C7��Q�^H�F�;3�ߧ��/�e�-,[]`Q�/����lԞ\-7��o=&R�3V ����w:#H*k�ۧ��l#O.�X���$~�/��3C�'Omo��������ӆ��殚�����_]������팭Cd��;(�{�j�SJ������4��z��eob��b�}R����L��;�P�{��)�rh��E��������e!�Q6�>}��8e�i�-Vlf�܅��,5��W�\[�lP�L��
i]��'�I�Z�{v}]��ٙ����߻Ey�؞�;m�zce�"�m�y�t6�l�&���J���+�-gmٯn6~2������Q뫒4KYC�H7Y�������u�8�F��6*-�6��v�v�3�N��zҡ]t��={Qf�&��W�*CM��}�{��&N� �*�#�T� �h�E���z.~5�mfC��
�
7n-ZP�Q��w�ޝX[��웗�(��uӀ� �9uA./MS)��z���O�AX��/p{�n�e/W�61����M4�S9F={�B���,A��K���r�ŋB�j��+a��k�A�� �r���C�3G�]�ȸ��S!��X1�Cҳ9h�؛ �VL1F���c��j��7|�(��.�> 6�P��v!cR�Q!`�����M솖�y�50�����4����K��fɎ�s4�������hܶI�ٝuJp(Z.�=��d���W�l{�r,<w*`YeuI��?hN�fv�!t�b��5���`�w�y����Ϯ1���;ؗ��↝(d��E^��^�j÷�y�z^�K}���׍+{�����*�@/�s����մ��w7��� p��<{��iC^�(-xʻ��7��������j�lu�@�[u�Dj{��ײ�?{:����G�+��h��gL�c#�<�+ۦ�#Z@C�6ʫ�} r;YOy/�v�JW��x��s�=�����u�(z�U��Y�� ;\���v�S]�k��~�щ�S�ǉ�/�����+�[�v�D
	'�4ڝa�u[>�a��)�՞�ʣ��&��\{���}2�o�S��W[� ��ʵ�j=�7����z��hf���z�Kʍ�xZ�D�t��~p�Yo��R���U����fo#vRʖ6�篡���x6��'��nV�RH��AZ]ra0<�{�Le�uS�:�ʹ^��hݏU=�v��3z^ͥ�օ����tV:�����R��w��"W!��ꭺu�h�QP�W���v_FCj�N��D-�	�3sD���2<(��bus-���W.3*� 9��F�k{r,1*�9���vb�鋮>o;£��&k�v��+Ec����%°W���p΅$�ɽSt�[ސ]��Ѷ=8�01;�N�nKu�<��h�ͮ#2v. ۮzo�*�3�bx-�B���"��/f�1*������
�6#��:����&R��M;x���/7P���y���{G��o���
�u�ϕB}�ǳ&H����k�m0�f���s"Æ��[~��M;�[��E"��N�!;V�[	d�`.u�N��XFmyh������/��o��b��J�^���ʸx*�ǃ�R<C�U�}a��ة�;�:�V�v!\=^V�}݂0�!z��]zά˟KU;P�:���ƀ���VY쾚��Vb۬�j{v0:2�s������xp�]�r��1W�<z���R��H����֗�n��wzvL�s���&aL��mԦ4<���!mAe(/B��H؎���/<i�y�zh~{��yo��x���0Ӭ?m�����]�HFk�˼�������p5�Z�O�*]ѧo���$��]��h�^��P :uc�k���ٹnvT'�
���_�@)<F�9X������58�>��}e�V�puᾼpwZi�S��M^�u�scMy��J�׼���'+�=W����y��sU]�墮������ip����BZ֏p��i���lG���xb{��А@9�}�f��u#���3݋U*�1}6iJwK,08�P)Ztޮ�/��6�|�؂���hKNݛk�M��IR�p��P�$��	rw�.���}���M��do��a��<7ݶx���c�S|(�w��fR�;��N��<�j�������o��޷Hg�i��@�N��ph��]b�h?��䥪��Y�Jw�#'���(�,�$�ˋF����*BjrP�+!���������b�ع�Pm����=v'&����g�M������I��H�,~�°V��Gǧ�����</�*��ߖVK�A�z�:�m���Dޑ�F�-��3q�Z�B��![1��h�����j�zIK��2��(:/�9���S\=�Y.��Z-^�f,���֕�}P��OB#�p���GYn�<J��;�w*��{�:�y��)&�;3�i?Fm�<+���aְ�:�Lg���n�I56�%D��a]���s`����t� �����J��~E�t��dI�ԞՖT��y�ߪfb��D6��
�Mĉ]f<a��*˸�֞7�K��;���ߟ��>L�#ssN.鴳���T�֐m;��i�+���uZ5bx���y��������uo�ۺ���b��r�ٕ~C9h�\�R���yP���|�����+�?���/¥5;ފ[�r]e�:�jjj&<��^��^J���	XV�,�JDT��s�m�rryz���xܽK��n�����)	[ `]���l��a���x��Kʷs�7���r9]N|yp����ڷ2�_l9��bt���x9c9ݑM���"������~@_b#��޻���tj�y�4����	�V���8m�KSҼ��&�:�L�6�*:xs(mD��U�\�!��������0��ZwY��p>+�������v}�gYz6��M����^�R�����.p z焙�t-�ֻ��U�kɳ$�ݘ�/zo_��d���z��yw��+��d�
�Ƕ�gf+�b/O d��<�c�N�Jљ4T��y�z���)����.���g��Ȧyk���3����d^OY���~�e���V<)úrK@J3g0��nB�Cp����2���	q��"�)�V����9;�]﫷��^lt��́9|r/q�����ƽ���c���쪑W�C�y�ᛉ���Y�4��:;5�c�PA]�����ovt(5�(�{��F��ջ�qf�o\�=�:�UO������7ܱѬ��8p��\)g��vu<
EX�L"�;�[S�ƻ Cj��uߣ%�u����23�3-"���}�/{�?�׻��.�Y���կ���
��[��%��h�2Щ�s]5K�!�f�̇��Ֆ9�)���{V]s��P������{��1�<��R�O.P��-�r��2�n���1�HA��9`��u��5l����\�5|����D�^���yb��-�-�����/^��R��5��7�������\@�^"���|es�� .�3>�RI�x8�5*n|�Z��`����:Ȝ�DYu�}��A[l���S9F������2KC�gXZ'�����k{�$J�W�	���e$:Z�g��[�?J��U�c����ضh0���;�'kum��Fd�|��pϨڼ>,+.�xQx�lx�5���
��1�ڭJ��fSZ���7����Y����{ !�����=�R�U&F�)E� 3����)WY�%�nV��Z�0���漪��ܴ0�{u�=�Zt��h�^�U���I)�����}��yGr�Cw�P2΄3L�S��,�,Ft�hïB����g\��B�oĉ�Nk����f-�.|����y����@v³_ ���6qڒv�y\e��Q��9���O;0���"�m�	�ݹ�� ��3S�`R�q��g��%gJ�u8~4º�La�l����K����g�V=�X�O� �m� Fw�C�k�=�6nG��]a�X	�z'M�Q�[�!��.8i8�+y8�r��{z:�����%J�Jk5�GS�:���:�ĳ�^�ܛ�>ު]���'�y���E����;G;�X��T@:�ɹ&NH >*�� Ibuu0���tW�-³�&N͔�|�i�|�lh����D����٫jU�k.��-	��ICW����+�엊4�!B���`�-Jp����?w������Lo�1+�Au���IS�����le*�n��	��Yl�SK+����r���F��1/}ǅ���Zq+P����ũS�Kj���%g��ʭJ����-ɥ<ڮ�n�>I�'��=#;4Tɕ}�Ս Jz�N��cQo!�ˑ����z"}Fҙ�4�v6j��/yR�¼}w�nq�;t�CU�VȬj`aݛM�{v �r�Ghjlgq�s�'t���wX1d�1
/*�.���ҁX��o�ņ�:B�� �͇��Y�sO8o�"�^,|#�QLN���R��ϥŕڟ53��Vq�\jKc+w�-*�!F��$E{�6�������,7/=�݆p��={{}C6:�Q�v�c�A|z��Ɓ�n$�!9Y��yM	�l<�Uн}��1�1���V��u)�;�Q	M�xqa�^Y�a����;wV���lZ����7��hV�\��7��d�?gp�[ڴ�bڒ�y,e��BKXr_Z��ta�}+&�uGj��u6�8�T��n�� ������{��1u�J��&<'�٫��p;o����o����F�J���V�J�d���������#�%Tś��#�-�W��.+ǉ���v`Fk�ފ5b�3w��w"
ȳ�h�ۥ��)=���0�s;��y�n1�2��e�#� �0t�ZYZ�S��8���ݻ}C�����)���@��x���w�	m�o ��^.s�f��f���8��{�^������2�U���#�M�5+�e��1p��^��������
���p��� ��n��~5�wզ��� S��s���5�@��+-��eu���4%<$��s嵓��$���A�T�5U�z���g�Qnc�̺(Z\Ѽ�s�'ҕ�S��MR��[6�i�-�J�[{��w]��hMb�jm���(R˻���Ɏh�+\���휴jM�g���w�w����v(N�E�i���]'R��S�2@���N���$>�b=@�ߵ�T��s���n79+���8-t4m�F�
-m`S�X�g^�������2��p���3Z���+��.ݮ���C/��]�D�\�p�����,��y�#���|�;w��U�)'��q���+���NQF1)�<=�ou#�y����&��b1�`δ�O |����:��l����R��c��#�j�ˋ��M���q���:���Z�D�cUӑ�<F�,:�ɴ����:�=�or�%���4��پ>�f ��ʄ�o������7Ð����Lpf_Wn�����'jQȯ�����1Զ�PY����$7uꇐ��zܹz��3z���U�o]�'��'d��*wpUv��4�MDjv�1P�;b"��N�Lwu	I�1J�cv�h�6�i4j*���Q=8;h��Z��N���IT��J5lhM�"""�"����-`��j��-mP�&j�b�l]۳]qV�QM5Em�[���f ���q���v:�u�q���b&�X�h�F"������Ѫj'u�m��(n1�mAl�c`���Z�5]��M�4WX"��1:"�6
�[:u�-�D�P�$A��Y�Ɖ�����TWX�N4cZ���bͨѶ�lQM3�h��tV-6Ѫc�z�L�E0i�F�Ƶ�F���  �$h���ޕ�ӭ�=�Nѵݹ`Ig]��F��vfb�ݦ��AJ[�}ތ��u�/�H:�}W�������OQ��x��u�<�U�X���z��px��+A�>G����<Ɛ�k��珳�P4��PI��}���{�O�t�!��.��46�y�6B��
K��߽^}��߽�q�x��uC�f��}K�x�'ĺ}���~��	O��|�O��u@{تB��������C��C^���=����h}�����G�3`f�~�!�� ���K7n&�hrv���[ޠ��7�"�ނ�������<C�|�����ѧ���'�~��i<�<'_|d:>�s���u�Cz���K�
��g���t�����<��y���qj���ϰk��kF�O6X���� �9���Ǹ3���>s�4y��O1�:�4���w����x�Iׯ�ܿ�̺t��o\> =F��g�z��}��_Ch��4�=zCy��e�@t����*�jc.k��Z��6�8���Hnn�Q�ܾ.����/�|�����z�����c�%?d�?���/��x��Gw!�_�������������<�h�}�����t���`��z����jz%Q܌�����y���x��=ƾ��=�}s��:�z=����G�z<���{�~�?2t?�׹|�cǝ��w��>$�������h~�P�����y�
�,ᕾ��R�m����4VflO5� `:�߯��4x���v��g�������%P�G���q������S��^���c�? �׈<���4���?��0�h�gĞ���
�;va���]����$J�,M���(:������Ǚ�.���oG��~D�R���߇A��^$�����I�x��~��ǘJC������|�P�O��q�ph|��u�O�t/56̃�����ti�C�oel��C�#A���|Ϛ���u���>a��?Kޛ�t�I�:<�~�����I��}ǘ�/˪_O�|a����:���:������)�?_��0��043i��z�Y�j��XN�4�g����{�~ꐈ|_'���_`+A�����<�h�����A�����`?F�>ɣ��`��5����&������{�0t:�%�i�π4x��;�����_�}F��x���Pu5�� ]��@wIt����Q��*��X��P��u�F�Sń��5�#�I=�;�S^h�b��tq��g���,�q�)`�WFl�Om	�fWV&���O:�[O�U�=u����Ղ��Z���R�Qf*Z$�8ի3���r�Y�bp��.K��y����u1x�;����'��$�� ����|��!+��e��T����+�����>ǨJ����?�~�#^�z���~A�|A����z���|����t����+��
_�y��x���ȧI��7SQa��1���������Gz�R����|�azrt>��>C��O�|��=�J��'1�? ����x��>��}��u;`��a�v�{vN�����{oC�<GBW���]!��A��pש~�O���z������������@y��y<O�>ä��x��?`��~��x��:��;�4>%���?O��G���z�uڌ�t��Y}_6�3@ohc^�����O��0�ۿ|�c�%?׷�
<K����~�$C�}�g�BW�
�߼��>A�F���'���O�:_G��<C�'���t��Bﶁ��4�-tJ]�V��{G�5?��?���|�_��Ͽ�z���w����?�����~Ϗ�'A�=��t�o��'�x���������t%z�<q�=GBV������y�4f������"ny��҃���З�������0���������?��}���4���߾p:Ph�~����}@}�>�ߏܞc�4?cϾ�ĚM}����f������z|��zG�{�3 ��+y��T�S��E�U�y|����}�4��ڽI�}�kǬ�O���׈=G��!)���y��GH}����A�����t����z�=�OP#K�}}���?o�������̃x�Ep�=����D�Eu��f�ϭ�~A�Q�?y��A����}~�z��R�A�G�������h~���x�����!��>���|���<BW���|~�����t?��޾�}M�3D� �n �7���r���d@t��~��~��zy�����|�i�>!�hq�^{�$�S�>}d� ��G��� >ƃ�G�~�hA���/�;�C����ށ�<�8@o9�uRF
K$^�n�-O��?�R����?z�BP���O���	Z}�?�+�`������y�0��~��~~���A�Дy}d�> � �<����4�|A��<�}���ϹT}�U�D|й;�)B�e���%�m���%�Z��br�j��5Szh�x���r�O'�h�&��=D���!�L�yF
���`dd5�����fᐾ������W��'�*��"���s��Bm�=��C6V�#���O��z��y�U�C�����M&����ǎ4!�}��u���C��t���݄�'�����������CO���/�Ϟ��=BS��'��?�8�������!�ᘵVI��P4�1�Q���y��@�`fp����,y�362{#������q�ӪC�}��|���k�{>���P��?�������y�O���/˯o�><!G�3���.�a�X�1�4Vp|�l7!^T^Y������${�E�y��ȸ��x���@h>��͏�ݠ� g�t?��C%Q"mT-BQcY"�U��8�3�w�^�W�7���
��!�SO ��j��k<��i�Oa��m<4�X"���u�Z��Gkkݛ~+ �}KP}+�:��ᕘ��|���G�+_ 8!�S�y�:���s�Q�\�����qm�9���A�>�5V6y�6]q�Pq+��v4Lډ�m��U���Q�xT-�ҩ�
+J���J�X�Y5��č9.�������\�y\��.o:M�9���Y�0�-O���qA6,�5(#{�u�<�)]�x񪊰��Ce�Ms��%�6r�m۩��[L�&m�"�?=8���{����`�]L_$J͚���)F^Nk����]K`A��V������--����0��R�S����L�89���y~�����UuՁ�5�}��f���&�y���9L�yW�q\,��$���8��e�sS�FPحd�eY�؆�|O��o��|���3��$���,y���6d4�q�JI�u�5i��^�,r��	_�
Mڧh7�x�B�zb^�'�!y�,Nk諧{&��9��F��V�.ߋ���e���b�i�<p�u������LJ��^V)䡜q��%���f��F0y�i��xy��0���^���w�jyL��{���z�9�w�.L�P
Y]�8���Y������xc���-ٺ&�.�U��kJ{j[|Z*Gs������< h�j�_\W_����6�x�v��f\H5���a�w�Ia��w��lFy:W����Y=�0؜G]8zd �8̙~]�\�qjfn!*Q�����<?Jl�A�E�x�õ��}��,񩠣-���-��,Aid��n�ܪg�k�Y���L��i-2U��A����μ/�UK�yyJ�&1)`l�)</�R�7qF+�=��f+E�璼!�xx_�
˾^^.V�����:z��S`�)��m�wܢ�E�Ǩ��(�la_�8�=���^Ok�-�W]��{뻦��d�>w�Z�ۛii����q��7��S�m�+�o�]�C{u��8-��k϶�������nӈ�F�
`#�H=}�{*/g�*�岭[�üOQ�A�D�mg+S�����z"p(�<u"N	qރ��w��-�`����o����,���`�T���v{dι��V��]����/�V���`��TzU}�b�O�736���X��bv�c�t!ZgS���X ��}k����v�<\�e@ih}��isZ�<�����>�+����t�⽅f�A�N�!8�R�0G%\]�֮�E����ʉ���Z��^u*��%��
K`Yo��}*�K:^cs�����%���ŉۺ05����{�v�,�k W�_yj��[Dm���7�}���yP6���:K|.��`'6&[B��*}4}�c��X+�������%]��]E��j�p�B+��.��O��t�i��%����ܷt8^���Le�*�<>9��=�J�[�q�)4�,D�
m�7�8���+��,Y"�)���!�S Ѥ�NQ���*U�!����1��Du��U�qTļ�Lf��d�dxQ�LN��e������~�� ΀;L����#hX�!�z"�,��<Z*
�g`��Q�Z���Qb��Q�!�=�
]�G�r�*dj �H����KO&��<_N[���z��0&���h��YB��:+؇�>�iKݾԩ��o���ǋMk=�V:ӼF���( 1t2�����MR�G���P���WA�Rѹ@Ԑ�������f��#�+Q�p��M(�uٷn�<n����P��K����u�4�S:�>�w[�t�ǥ�6�A9�1��P�ֽ����$�S�r�+���f���^7(�d�Wr��r|�V��B�����f�u���~�օ���@�#}WR2HLՑd�Hd4�������:��z�,̟O�Շg�q)��II2�-r��F�`3�"=N��t���6��i��t-a�U��3�4.y���޸76,��o<�N��{����Y����ah�"Y�a�:�(8��/V��b��bq;1J�SC#:UT��|y=3X�|�e~�b��>��������AeZ��Ws��
���z"�OC�׻�j�Vq������:���V����Z��f?�Wj�����W�{��]n����K�]P��N#���ѡ���L�͵f�-�s:�S�}��������Q���)3�ƭ����5�"�0!�bh��j��sU]�EJ��O���
Н����1Kkl��W���!�~Q���O\����� <ū�u���2�����Z�L��-^=�iy��-z�[b|�-GC-2�=eS���}���VPƅ�`�E3�赁��2����/S=sfh��ݜ���AB�/�4{xK��}O^������>V�R+��C��f���� g:��,�in�[]S�R�b�p1Rӎச�t��6u�R]�T�`>Y���tc�����*Ńqq�^�nޝ��W���*a��E��>��]?i���l$��;L�ve*e9��jZXF�Y��YCԺ�ȝ��m-�y��
��קO��s�5t+�Uf,�c�C��>{S�l���JR5�'�wgej1��/q��KEd�["ê�Rr�̺��5�^m=)Jk0x�a��a;���(J,��t�`h
X(�;m�!�l�o&oeל�~u"�_�xW��(If����I�K���wn�B�Q���V��F� ?��1��r�-[�Eܶ�]Bs��n�H�
�q�n��8:Z$�6L�I�~ �;j�AW��H��b<a��;Fb�ȶCڬ!�Izj��s1��L�^UfY�����i���S��H����$5y*�֪��2]N2�Yb����.h'۠�Q�P�{���,7YaCw�3�}��_suJ�/O*Z�|�?-�g,��w���3|(ǅN�E�Ye�&d��;
 k�v�.ʢl�Wn�+H���앯��>��j-���՜�����r)賅��s�F�7F�� �W�/�
�X��e���}c�yêG�����~��/�Bְpu
�쏖 0�Q_���o�ڥ����!�:��U������v�9`�v_�w�@wԏ�j���G����2���-����G�"��⎊	��b[�'N�z�⦴�I0�3x4�;.j1u�Bd��!6�n���s�������
���5fF���񇼕e_�#�!�iz6��>R�q�����W_INQ#x�{��d�C2���oHP�>�S�Lo���|�xMv&�Y�~d>���1V�Wm�xK�b���0f����{x�yK�2����q�gh�Yd2̶�A�i�ۈg�t�u���s����}h����WK�s�ь�� �*��N㲍m��8�+��n���]h�P[�g_vu��{7wy����*^㇐x�عX� ��g���i=��W�w���13����g�*�v��A{��YU����(V{���R�ڱ�c>�5��j�p��[�t ���43KC�6�lWv�	�`���s�]� �Zj�w��+$��Z�)�����iT>����yW)]�҉h�át]�;���������o�}�8�~��Y�G�7���}��;ď��>�d�hזg����9@e��a9y�����i�^�'E=X9{|����l?}���i=Yx�VK����;a`�>�r��<���}R��)0�D�6�[d�cwI i��^$P;]��m�e����{y��
ή�0'F՗u��e�L�;��_c��r�M<�+X��u��Heo=�Pt7���;H�9]���vY�|2�k㙤�m�ӮJS��SÛ>ġ}����+T�=Rx�A���v��%���倧o��~���R�;��%ޗ�
 U3 u�ݘ����{�e�3�V���^�xxX���
9U��U�����Z�������{��)����wm �ԣ�Lj��,�n��fP�g�)S��j��ׂ�#��^m=�J{�`����{܊E���O"����JN�ϒ�gT�DG:6�|��!���Cj{C�Li4�Cw[d3�H��|�Q�P�h#B��S��+.t�Kg��bOk3������ǋݻ䑭�,�}pb3e��Վ�_ ޖCFaiK�\�N�-;�!��$lrվ�����r t>�������v���Xkn��A$�f����}r��Tiy)A5�Zw�{w|��
�{����}0�ۨ r-�R�q��,{������b��ɍV�Q�i���ף���"�vU2ts�����	�\{�5��%]��]E��+��.���T��S:Q��훒�4'��g�BY[�B�.!�(F[�
i��j��O��1x�r�hۏ�"����f,�U-��`�E/�ԫ���,x,������;�3%�f6�J�qW�OB��o4�`%��c5�.�M}�7D�x��۰U�����������$C�;��A�K�j#)�^Q�&�t|�N��i��6m�{W�vq��36]UVn�J�ؘ�}�e����m�W���`�ބxS�ƅw��#+������w���N:����o�gg:��n�L-{�d�1k#�Ɵ���P��dA׭�@)O�NJ���O�ySw�煀'V��Z�F8�Z?:���.��/XUεy�O�����CIK�?nۣ7yd`.դ���
��V:�%`��V18X�Vu���֡�VEj%1�s6�P2�(�K$����R�C-�a�����zsƅQm�ʍ�^��� �Uʋ$�[M7���� &�sDG׮���HW����	u�`��-u�;X�?�^-��朲v�މτ��� v�lwd[�tp)4�v����(���q�kܵ�����)������&#[R��3�,զ,���PB�¸nCaJ�����l��y���jx^�ײ�z�8��c�^h����*��U>�!��}��/3�=�H:f������ѐxf�s�y�v����{״�v�����@����i{Oi!����y�����6�&���9�C�2�N�^��۸�/X�-/ݘ���]��mlF��N���]n�]�m��>T�ï�E+��B9�	���v�N�j]r�~Sc����Rj��vRq.�ͥ�X̷�:mL�F���VMq�c�,9k	�)P�V����xs�M���N�ܬe�P��Z�����H�t��,���ҕA�����z�u��&wm���6�����mL<�ljr�^:U�L4'��)���:Β)*W}�R�Y�;��19���@m��f�Ԓ�A�1V�;�_,̽�R��S�՘3*+	Q�n�2o<+R��M�ѽ�ܠ
��z�TY�C�����)���Zξ�N�欷�a�'i���|�	;��+J�ѵ"�F��j�Ү�
��$k��w%�զ�<�f�x�����6�[�ի7�H:6*lw8�
��f��^�>�g���d�-����w��th��;�i��p)�*QȺG�񝼱������I�F�E��o+/�X�<�7��ik�=��@.��_-��tG)[�f�R��L�9eJ�
��7�-��	��]��5���>Q��L�t;w��j�%�mn�ŭ�Xhգ�a�g3}�����É-��Sµ���軎A�l=�5:1|��Mi�|�]�덅/8�C���wf�����˞=��jѪd�*����n�Kp]P�['L',���Wt��k7.5����wݙ�<n�pJ�n����=����52�u5)���<4q�6N藰&�:�>-��@�je9w(����*��%S�4)��.��c@��*��#FJ8������T߇�]��d���G:�V�j�ݛ��Z��\\��~=p�s��K7�(	V�yG�� �ĵ��eO7z,Z]�$y	<�,!;b�����:�u���գ���4���M��S�Y�o���*�J��b}k�WԎ}/�փ�����"��-H��5t���e\[�C��:8����W(:t(^�;
 �D/��腣�w*]�� �u��N`d}m��܂���Y_P�b��l��V�M>e�D�f�
�	%5.�<�(r���(�J�m�n�먍ՌTNXףi��zGu�Di�ۇT#7�2�!si"5��)㩹@��pBWm�����ϛZ�pX��;-;2m�Q
t��9�n��8(Ñ�e���0҆��.x�Z[�Rڅ^.��������.�<�;�h�V�4��/�s���г�Ue����uP��k��tS#�Pn@�f
Λ`��^O�Wf:A,�r�.�wd%0N�j�Z.8=�(�Æ>=&�w=+����m��kBX	�4rd�&9��;:o:��mB�n��M�rf��5�5M�v�>��A��u����t�̫E�v�+
s�Z�`c&�����*\5Χ�P�������l��%��Q3��s���Wz��pg�|8�m��;Z)�����cF��W�gFj4i�t8�*&;��X��műZ#X �3gZ��#Sض�R�Q�;i6uQF��L@S=:�:�ؓl�
�mh�lUUci��(�+l�D[Vb�b.��5L�1Q��SLbδQDT�EU%f�*���ղD��E%��Q���Q�٧U[v�ճ����hլD�D�Z�L�X�Qi�U$�1EAE�zꪪ"��T艠�*���;�s���:��+F�m��T��k8��(��Q�0EE���*M�QPSF�V�5M4F�QU�6��55�f�@`����]�PU���347e��*��kUD��[�F��j��ã�h�I�Ӫ�4�|y��߿wr�Qݧ�t��a.�60�x���IبG4f�s��t�WRF�7�z��v^Υݹ*#{}ݙ�DRNn��;�磌��H���������q��X���S�)�zK�]o��-*��\7ؘ�:M�L��I�izy[����6n��5����0p�&Ϊ��2�O������WAzz��~ѱ�9�+��{��_+[3�Bm���װ�/JX�t`�U�G�i w'�4t�)��*�z�}h7+�7�ڝ�	~��xb���[���=�u��{�UZ�bs����>����>^W��8�|�7+�U��on�u�\O�����U���L��`��@xt�G,J�O�R5yx�I�&�h��*���-�T�j�=>��l��B{���|v���ִ�ԬƟnBĢ��ݚ�C�&�����L�����,��a��u�A���9ttk¼J��;DX�W?���w8����S�����[��(JZǵO�n����?mT��tt2x�ǌުwj��2��)1C6>̄�( �٨����X�ٮc�-ay��H�>GŦ�[�F��"��E�1S��3'�0� ����x����P8�)��zNf�ވe�M�r��]��C�=N������P8\�ceb�H�3t��gw%�y�.�ie��?ʛ�~V}��^�R�2:e:�eh`��ze���,U�ݬ}�,]9#���9���>�2F'���S>�ݕ�:�f�|*�6CՉ�ߙ��{͖��[���+�aq<Z���6����^5P�j�����-���K�ST�A�t�_���i�V��O�>*���ҭ@�֑I����aBv�����%��j��j�c�$46'�@i�v7����L;��Ƈ�Uk��n��𥴰ɦ��&VŊ�lPe�͋���;�U��~�v��+_�����B���.�\Jqh��Eä�/����"nǉ�RU�O�O�Q����0>��9q5���y��0���L�M�쁖Sk�N�g�^b|������ν��º� ��'\���^���7�M�Ѽ����f�7�,��3�m٩�ޡ^�����u����Lz8E���$6{�j���g��"�aR�Yv������d	-��;�8K6.�k6nB�L0U�.�"J�g�J��Ǽ�ج~����J���:��u��cf7�l]Q�=�JO~�0����o��5e�tӢjr6�ƻ2E۔Y֛,pm�\��5��f�P9�R_X��Ur1+���li�����/0-B
�
�;�:���U�8���Y�l��E�R����k��z���>�9�ۂ�=�<�J�.��w�cŜ6[�Ǣ<x���r�]�rZp��ב�n8�s�Aآ�5mq?<���9�V���y��f`��Gsah�:B�}�������p�5O|��YH��-�F�UI�+�@���$�� �V���or9Y}��:e<a����k� f���ڥ;vk3��~�8��7ƒ�M"
�av /;��y|c˙�|��1�����Ӯz�������kk�6N�K�@b�Wk~?$�#�*�yL�U{��W��҆�iʼcMj����X36.X��>�ܫguP�fvj��^�.ԍ�P�F��ԶQ 
s�׶�|�s}�w�mN[����uſW��	v�8Oy���_�oP�\95�jQ�G�%R�{���޸��2�y��,1��z]�e�����<��4��u�Ot��IB�����>/ō�y�{��k�T�Y�s��1��tD�Lq_I�w=�p^�R��+��~S�ޕ^�^�/���5��՜:9��tj�/y�}i���Ұ�����.�����4n��)�`ƨ�u���NͭB'ZM�Uo�
�{�{�jzH�h�35�n�]^������ӊ�i�r�3��&�����Ҹ�܂�s�&o9ۗ%�Ϯ��ڒ���iT�<��w�)���[]Z��|k��%�����X�Ni�/Z��}UUU^J{�\l?xj���ެ{S��g�g��g����k�7���D�:+������ct}G�q�|���V;�cU��[���G�쎳kt�myVi�Ȅ��1{��5�g�����qB����li�Y�t�V'�ڷ���yï�^^��N���?Z6떕G����[ʡ��j�j��X�P��S��ɒ��5��SHF#9�U�k]��q�©1�M6 �5��N5��/df{�^�V��K����>$��K��J}�uީ��8v����S^���y�=gǈ�L�w� m�'�f�G�٪��}��+�=;�W5e�Z{�n�z��^Ko�K?��-r�����$���gK�=^�z������C�N���	6�5��6یu)Ye��L�U'��i�B�1�l�.�!�^��iDL5��R*Sҝ5�^Z�Q���MUhy�ofЬ4��2蔙@�ey^�ջ�b�� �{��p��'.iG�Ec:ej7��vХf��}���S���h1�vg*[h�c���u>��3�^�gY\�Ӂu�a��rۓ �];���@|���w,�9�t�h=g�]!�vL���(5�ȌQ7���y��U-6�%c���m�+m҆�:�h���w���h����o�s�U�;u����E�]�+��o*L�&��}�ŭo�jN~~���j�[I�F��q׽#��}�yeq���W-gW��]�SZ��j��h���*Xc��B��c��ʈ�po��������Vv��j��6�����T�-����������^V�������(���$?/^w�U�5�śD9�G��,�[�%���zo����R{���Z��Œv�P}����2���i,uZx�F1�� ��=!���}1w��[q�*R�Gg[ul��
�jŎ��;{�����E=�l��}y[��D����>�7��^�-�3�p��q��dias{g��=�p~g��&=���|�J����*�ʤ��T����TZ��ɖ�Q�Ylz�^ܳ�)Q�w*�����*
`m�5��V�Z;q�C[�W`������V�(\�'_4�F��BM��+k�c*a�&LP f�tƣ��)��K ('��+̝��d#�̹���Σ�_wi�֌W�����5z�bLP�.c��hͣ�<����cܧxxj������32��G&J�Oq������@��}7§��k	�{��Az�%O���P�e��fX8�}]ܪ�z��w��>�4��g�ΞU�nF�ϱ�����C��R.�;�r92�)��7վz���R�t�.�m{]�b|T�5L�̤���}{���khՍY�j`�JZ!}u�S�F��od��=-��u8@qyb[Gym.����*�{��Y\�=�w��kss��R�C<��{����{�6=��A]Ŵ����>����&Mt�4P��1.�Cwg~�/�Y�o^e�.�������e1[>���R���_ygg����ռK�'W��>5S����=��|��Į�����yZ��]�C2?8�����&Uzp����*|���U�vIp�yT���ו�9�[�"�����WeV�~W$��rzv���zeϾ��v��\ �O�=p4�B�g�ȷ������V������e�\:~��:u$.��[x�K7ɿz�ޘ�[S]Jt!��0�ܸ�]�ݷ���}��y�i�D�N�b��G���$�Q�o�eq��a�o9�ʎ�fgW1����O�E��|@���e�Ĕ��t������������~S��y������;<��:�5��J�X7�\@��uGg�(x��[[���3ޜ<M��nI�3ƶ��{���S����B��s�y�xե=�,�����q	�EI�%s���.��;L�n����b�*=|�6�R��2�^�٣J>�b�#����'��,�g���lYwZr�TUw{����R����B�5lyUv���؂آ֬޷7Ӽ �ݝ��V�j���{�W:fF��YG)��0ې�e��m�Ye����-��z�Ag}^��)	sw@�ۚ�Y����&���(de���B��f(��8�NY���?%�{[�I��|2�{&_d���^kM����#J�Sy����;� 6���zo�	��>{T��zF�*��08�qF�H�LהT-u�O-ڧ�`{��>	v�N��`q^���M�v����R�VӱXr��I=�ϐ�WHA����S�G)F*��)�bt��/���f�p��Ӕ�� ]<g�3/��]H�㻤S��joc�Us4H�[�G��q�K�7�\Ν�]8WL�9�s�v�ԹK���L�1��z^n��U8a�y>]�������a�d�$rۛ^]��SKj
Ta�;=��?Om�!���3a{�v&��%�|��Dm���f�t�������>4�Xߗ�{^�m�i�,����!�%���.={���HSW��Hx��rx�.�>��ɁQ�뷽;���>�q�n[&��ӕ��4��G�;�)�k$��4�mɶ#������B���?*T����u����T=����s�뽜{!�+Ҙ��6��E���|{��Um���D�C4�x֓=�{�!�5[����y�{t`��NP"S�w��%�O�q�W���(<;��k�;
�R�{�O�dr�fCM�Wvٶ�|�S��JQ�d+�i
����[
�2E�}����z�i�ϴ���<m�u{�t�T��<=�e��y=�)���k<y׺���^~вm_z�z��Y&�av�孲9�(L�64�2�:����N��<�;�6!.)C'��e�Q��Eh K;>��d����l�)��W����f���r�ޝ�@��5�7��.�΃U}�y��Bj��أ�w!p%.�:�' �[�iJ�!��K̂�N�a������y���o���b�X���6-,�SnC27씬Z�:�s��?Vxr��3����0���RK���0WPN������W+� ��W�����k彾kq���_Z��5jof���l{��,� Ŭ��u&�K�%�U�|��ן�Y?yvX�ziڲeK	��Eg�=$%��I�ܻ�sYk���s{���4��=��x��j��cn�a�hf�ECRz)L,�jw]�A�����v�ݓ����Ib�MJ�X�Y�&���Z�̲Xe��\�׹����e�V$��35��R��>I��[O�T��CW�ِ�o�Z�3��H!�~+k���y+���J��Y�.9��}S��q]�Y��^]Ɗټ�53f��8�Jݸ���U����מ��LTD�͕�RM~9�~0zq8竄��s��Ѫ��m�ץ������\�EJ�
�Z�Z�b�vS�=W�:�gV�K�p�qŻ�]��g���(�KF2�l�[e[{r|����V�^�@��[�:�M��U�X�w�ܲu&�ak��i��op�
g�teЕ(�����.L)��c=-t�Z��y;����'4���It�V�O����Y�{c��Ƕ��~�;�^�m>�Wz3]޷�y{�����{i�ǐ�f���Z�Z��W)Q��kj��G�i��q�)���T%P�M �`�}�T�/2�DF��"˶���x��$��4���o��������p��IPl�C�D�����ڡݼ9U׻�}����kz]�6��VC9
�H��m�0T27Sl2�;']�����*y�e�	��]�ڀj=�_����V��<�����Zc6F�b��eu{�׏�����X���Un�����NM�{+�knX)|p�>�ذ�W�Y��e|e���pi>z(��I^�{�L��j,�5*ڵ;c�|!;F�BW���V�hc��r���FOy&J��]�1Սj�z�>�J=�km"��`e�Fn��C����G�l�Cm�g��})Z��oϪ����ͻ��^g��n]&�ʾ��^&0v��vI�����H�\�uI.ɭTEv���խ��W��/�{�uYh�ﮢ�Z�Ў�nea�����BO^��'X� %k���X�G
��t��|8dʎ�� �k}���`F���F-�X�.d����
���������R��Y���8@(�Ǭ��L�ڴ!ݍ�Ti�x;ybZc��WO����%eA8
�UJڌ�wMf4.��u.͆&mlGJ5��ϲCw�;E��,R�j�
!^����թ��ޢc�1 u�79�v��W�X����9�c}J+�n+�U��Xv�6Y!���	Y��[�F`xk�-��dU�l���`��v�����/2��������ybI�Oؙl�i�����e��La�g�Kn���&!:H�^���+x!��T�Ρ�ep[��i:��ħ,Z��!��^+^�������<���m�����Ɉ����Jh��y�� BS���i�P���t!}��}�8�7������Fs[};"�F��i��kJӼ�������+�
R�E�]۸ufk��l��9Jy���-8��7.�+0jwXǹ���^E�r���L٧V�NS	TX������b�8{]��:�J���:�(�]��Y�o,ã�������}��N
�:��(|5��09�Q���]m�&���T��'�V������^ʟJw#+{���YJJ�2f��oP���Aj�ϛ�V��)�f�ڰ-WBp��c
�OغC�s�C�B�}9.^������G��|��>+�a�N=r�B�"����GW��Р�K')��XXS�S�&��c!�o�l<U�캖47��Pzܒ]Ǒ̼U��C��&��
�{�Xq�)މ�����%��4U��bOә���^^����iB��1�J͕Չ r*>�e�[�p�qut��3��H�
�Ƶ����c��ӈ׳�z���|k���x%n���7�K���>���*�1�'o6<�-�z�뎯 {��2������MXy�U��h��6��Z��4 ��
�`Ú�Z1P4u*�J'�.	��r�Q��蓦�f_�R"xJ PZ̐���T�Vc����Q��4U��S�T������g���V</Z��t�i0�,����H��pr��և<��7�U�X8�����1\��Nd�E�f���Mشٯv��鞎P�#a�R��U��ϯ4����t�J�э�(TX��˧R��"WV���fet��um�����{���-0��({|�p�8c�0���\�����s{:j��6�]�E8�q���b ���t��@�\��z�D�,�JiWuv���u��]���8�Wlh駩��L�U����Qxc�Q�fu�xu��V��_��1�|0�}�`�η�v4THi�kADv��:�E�( ��(�椭�R&��������D�Pm�(�TV�QQu��SSZ�Fƪ����b��:�SD3U5��l��lRUTDM[i�����Z+GI�A��������c�b��Fi"�5�b�c�u����K%T4�ED�h��.��8��֊�����h:1kEEE�EkQ%DTS��S<Z�"#F)�muE[h*�"	�&���U��=�WI�i���5Zzu��N��* �gT�����k�����Ut�"b.�N��*���֊�u�U1L�US���p` f��,:����x��6З�P�n�}��]�o�I��q��)g���� =-��/qY��i�kw�^ӈ���"�Z�.�����f�0�RK�CWsߔ�`ז�{��G���Gg~�-|i)�K�z���9��:B�f���J~M�S���N5<X^!����~�+<ů�<:ιS�wꄓ�u��=��x�T�c��*�ӆ�����y�/�M��_q�Įh�k-#y9{����6�;��MdI�R�wm=N,�zh��;��,%�{��y��}Q���9��>~�s�T��Ɨ5��7����T�p�4jw9�U�zz��.���>�mp�%��f��eG޿g[�]Yc<h��t{���	�9u�=�l'EWy�_�ͽ��;�Up��u:xuy����q�J�S-�s��8Қ�'v�ѻQ��ϕ�R������k��o^U/+���q��Yۯ��es�2X�V6)k��C%�BP�bc�p��(6�:Cpk���g������ �^�^[�3�fB��hQ�a�Lk��f�E�W�Ǟ�=�>���h-/3ގt�� o�5C�����8W@H��Ka�s���3�lصh� MZ������yS.�zŕ����,�C�̜�!)�4$���d�/�<sE5��E�e��;w�V^y�埃���ޛ,�3^���B�p�b�����y������5���b���[��;�Q�6j��|߰J�T������2y�|䈇�ܴ�'C�W�E*�o�7�䗢LeR��ߟ�Ơ�{˓6����m���[M2�$�-e�,�
���jU�^�.թ�?�wm�W��X��"ܙe�(GT6����krmL1���R��k��o��Y�j��w_��LC�](S|Q�SG����4cUL-�n�7�{2�)����;R��A's����W�v�O�O�ś&��{Z��VI!�u�`�gWWW��O������m�,x��5z�kO�N���Ǽ����f���$���>��CT9+���ˎ\�NwɿnT�ü��褿�1����3U�J�[[u�Y{�lu�TjF��cq阉�Dt������U�s�������řv��T8���ۖ�a����KR>5�Ϋ�/U(����W`��C�Rf�@���:e��N�=�j�G�:)���h�kw��ځ�R�s#�9(����6���O~��u��⺨���>��͉��k�c�B3!�\�:�(��4{t:O1�6wD���ά�Gݳ����J10w�VA����jy5^���DЪ�y����������5=-���m��k��k՗*�ኔ�`��l/V�C����h/ݻ=�}{ɩ+���J܏4��6,�j�[*�?�����mȧ~�SB�Ʒ���]��]B�]����"l�G�jSB�ޗƩ/v����Ľܷ�osb�dJ���2�5YHy�d�;n�w�fg���w��Ś��z�����g�<1c�O�w�ʇ&U������ZϨ�Y���6j��O_����]BF�&m��kb1	jP�5�YS�E��)�>K���PT�{�c�@�G�^�Ry�^�E��lW��h�4̵���d�Hv<�ܦ=~l\�q/�<�b�ы)�/�Z����LT{SҖзЀ��͞W�I��<ƥ%�c��'�ɩz������PُZ�֩E'��!���>�u�=咗����}�|�����~�bߗR���:����>~�J;7����h@߫)\T:�,���(����tG.D��u�`���=��AV����P���]/��Z�G��η��������݋�̥3Vvp�0��Es�;Y�b��ٛ;�q'ous{����7�:%U�¡����J���k����m��-~E�]K���&��K��K�����T�!�2����ҽYz�"_�F�Į>�u�K+�߈^�>��2*���l0��I8�X��wr�2������������mv�}��q����+�K#��䭩��=�:9��3�tq�Yڸ��P��us��u�v�o�g9޷�9������^�˔��6�n>�
�E;�{C��j��s�c��Գ�d-N�'E����՝�~yƷ�g����\���uۛ�=�{4�v=-��/��P�3���Q���q&�A��"n����p6�.����!����>�k�)�(��j-�r�OP�L�nL���NeV-�0&�$Ԧ�P�oS��Ӷ2u6���Ӧ��t޷JRu�Z�)fe�7%$���[R˶�O��ڴ�:l��*��>�WM��~"�� �F�a(*�n�U�N��=�ԡf�|z6ਖ਼'�Ns�tn⊺��j[������l��n�\�$I�18)ݭK���W�:��gq嗷��B����Z~�(�g��V#�wթC�^���\jv^��)KK�Jb���Sn�K@�z�I�8��ٽiy&I�E��Oi�έO;��着��g9�~F���E��+m�#r�w�blS㩃�1ԥ�K����DxT�>|2Nt��(�s~?)����j�6[Nژ'�t����<�[�F�7HY�sb�_˙mϝ�Y�%�H�o�å�)�.���]=�ޮ۾�t���G�`�y��y����h?��|���1���֎�>�ےM��"CEr�'��K���v��P�U�6������yk���W��3J��<Q��$�q���*{|6w�����k��r*��m�����n��5��7����W�*v��O�*�N����}�ȍ�Y1�����AV�lus!:�vU���i�i����Sæ��P�-8����c击Z^�mA�^�t�=1eu�L�#��=��}�{�
t�V�a��Oe�89���~g�~�����U��Ro���v��Ǹ֎c�V`ɞYj/L����pj�3}��U�[�kC�v𖪤2�^�5aV�Q��; ڈr`��0˞��G���97x�;Vl�����:�&
u� �:iu���u�ܧ �77�nhS��B#���u�HD�P}�q���Ҕ�^���e9�Ϫ�����+�wI0����=�=���m�;���z��j���9;OEP����jT��:��q6���ij�*]��!�F�����x�x�F�U����h�\�j"�S	J�kS�]襶��a�I>\i9� �^�0˙9'��/וn�KE����WkyC��g�V�i�{���T��.]�z1`�Ͷϥ##໲��s�\^�.�`�:$��{��UY�y�N�%F�	l�Xp�W�ڙ��z�쫕�v^��Rc)r�mS��6��t7k�,v��Rn<���*��ρ��q g�����+�O�|�D���EL�X���a�w�d[?�"�N�-��`e{�-�?#A%�&h���r�Ӌ���I��U3�ߣ��4/x�{Z�t&�}^C����}�9��w[�/�}��R�/k�S��o�jw�������ڒ�r�+���߳�wo�nW�ۍ\�_�M�#�e⹭�\����j�+:����+}�/Ng� J�0j���C���S,붤ɐx��Ӟ�a�����z;��S��v��k#':�=xQ��KmI�Jֵ����7����#-��u���h�S��v:�Q\����U�x`>��zr��^����}�^iں�m1�'���N����}%h�������D�I0�����������ʮ\s~!v��Ŏ{O����q��>g�y��������e}���>��)�O�s���{}7d�㾛ZT��U�p��'s��^0��
I1��{�W���N�݊��޿iO���|C�p�;��5��>|�x������o�W8k��vZ9�m��x�}�E=�ﾮ�߉~G��u=&���v��gv߰�{�Y�iq�Hwb���q�=Ne?x^�y�MY�6�<�ԥ�o�y���~�!X�K��S��Ad����j-{r͊׏����J��/u��컳9;=Pt֚�ה��-��P��(�:�}�u�C'�b��l��s�V�mn;��sv�H�S�yVo
ڡ+�@��}�w�%c]{��ޭ�i�Q�Dw
{��;�ii�����%�7�.�����y.n���1'�#�岶nd�a��ju4�+�H6�����A�>��Q�ś-�F.��a��ո�A]�k:�q3��着<0j��}�fk�6�>8�lAݛSb�lwJY��;jT��k, �B#D-�l�x���}Ȉ��*��v�X�̈́'m��CjzR�V����ҏa�����V?oS�jz��3:�ƭcn�6Cδ�j	�)�ٛ�R����ܼ��UN�r���P-���-]K��>��ά�����*d>A��[>��0Ua�X��mИ�-�w>N&�[`J��3O:Ӵ����-b�Y���nr����7��ϗ������ܕ�kؕÝK*�q�k�+��g%�2��Sǟp�����v�N��/�y��O�"@���fQL��BD%!^��������ҝ���FԍŖwb�n[�c���o���7GgV��K�<�y)Qz�ʲ��&x�w�tY�g�w���y]<�N6y	�߷�p%�z����W3���Gg�=��*q�Q��z��vv��jI�wi��j���[:#�-[��i�[���ubYщ�Sk4)�XU3�s'u�bZ���)j�����/536uq��;(���|�K,mY�
S��[��V^�y�Ʌ�Mn���2#Юq)�u^�9�ɥ���eŖ+@.�6��s$]f�����
��ѻ�R��y߫�.��z��d^V�t���.{��N��BjMփ����B�诼��T*��ciQ����e�E�lњd�fXN�P2��&*�����J��Zm�PƵ@T/56����:Y���Z��Х7�mvK� �ަ���w���\8�~ɗ=:�ǘ�mX���1�ݺ��6�cG�f ���ѝFNq&�*n������h�&��L�C���ʨV��k�y��=Y�&�����E�\�b�g�h�^�_z���3�ބz��Ey�;o̺=�bOR
���`��_����X��#��Vֱ�I���
1�Z+7kD����2���a��츶����#�Wy�~��eׯ�9�}���}�%{��(ר�/j������{��4	[]�������ݬ�V���]����)�R��S��jw�Oj��{ܭ��J掫=�;.U�^�u��U�g��/�iv�=ʔ��e��AU�,:�0�S0n�np�
�PW$�7n׳��Y%�w]���2"Qo�[nH� �:���\!����v��QL���9�T��`��BJ:��;��$�|w2�t�r�Z.���;*w��W�_,Z���>�˯OkB��=)�'�UJp�N����]��Q˼̦�����Mһӵ[��d�~X�W�bp�8}�0�:�5��{T�}�[�����z��]�/
��Խy��a�EKӥ?��uo�c�u����՝�d����]w������)��o���k$�{kvxO�t���
YG��Dx`[������՗,�S��JXe����+�>=E��&���6�fb�i%x�w ��ݵ7j<U�m��V)K����ۮҲ����{w W3����Hd}�=^��|&u�W�UO3��1������O�
���l���,���G��<���AM\��S���K,�����
9L5iқU*P� �sl�,�f՚�%�-,���{U,�-�gi�'Uܰ��6}i�B�^�^~��t�Fz�.�b������5�<}��W���c佭����{6��{�	�9
M�N�R��M�U֚s�%��ۤ�uصp9s� ���@�̞Z���έ�b�',IV��b`Kv��P`#E�s�˕;�`����z�"ؽ��GPfX�%�'k��y�ܥ>pY�N�9A%�xˮu��E�-Kэ `�p#+������\��`�:� Y|kn``m�2��:D���t�����ךּq!qP<�0/ef[o�ͮ��%r��̋��n- j�B/�엲� 2��Ư�K�xx��.�5֎f,����mn^`�L��{�s��I�V��ގX\��w͝o�%�Z�f�Xn��k�b���ZQoO--�&2�WY��,��*�ac���}�����S�牔��$�G�q���v^�Z�#ʽ��0{��[7��<�k��eOx��4��[��G�V)�)������J���}����u����_<x`T+A�ȗ\��:�vO.��3��zJ߂�.�=�5��IU��k��[Q�}xڽP�4��S
绷*��6B�xCǯ#qS;DR�&�98}A/q��&����Gڈ@]ȑ�v.��X�>�<F��9���éM��7��"�b��N��r]eb���Ǵy�o[�3�`]������,Wdh����76P�ݓ��r[�k�yV!��_e����.-*�g��5%yD����gX�.Ff%wOR�$}��-1I���O���}�0�<�:���"�2��;�N�%�N�¦wcM���ʖ������gL�I��͇������kj}��n��rq�NVt+��J��2> ;�Ro{���9�Hu���Q7]�����o+qt�Z/$�ҷH�y+�t����A��Xn�=�/Sv��Bv� w�+S�O�������ڻ��o{�����el�n�ʳ���v`��u:`���;��/+�;�u���6�!{`A��#�K듙Ү�9Van�s�8��բ�YO��66�̠��g��u�"��p�kC]i	�n�d�fڕ�3�� ��Lan.U����x�Fs�v�]hj�%�[x۴�Z��2�"�[�`�a�� �-�p�K:LxvԛNi�i�8�]��zMt(�����K��r�s��c��.��Z.���΁�+"p�������c	����`��Þ�r�MAL=*t��z�*W�c���n��Rޜ�an�Sp�<p{=㣱�:59vx�2��@��L,%U+��m>&�Ήl>���9�*��������V�|�ie]#,�in�\��@`�3{�jL�u-6�]܇
)vQ�H���y5�{�6����3�a.*ެ��vm�����s�4Rb�o��;[l�ج� ��B�}���+��R��a��vK��p��� �-)��T�����c�B��|��{�lGS��+��!,өܷS�-���m0����۲��չ�u�O¸��L?��2�}���ث�#[�t���`z�f^�1��������{��o�>��63�ܓ�b&���].��h�T��������4�Eh�m��4�%$IHW]�Z*�����Ѩ���
(�-��J�9�ц+�4�=��f*H�"�h��J(�ؚ5���Q1QD�;cmAEEPL]�S=��66�5T�䋻T�L�h�SI1DշO%EQ6�0���&(��ͣ;jm�l�jh��(�Yh���+������GTb���(����TS;�s���M&��CI�TST]�TES-���h���i���[9��m�;��3UWlEOl�8f�ZJћX��d�f8��{uB]�l[C�=�8���"k�Mj&�� +�EQ=�1:�E�V���j�޷��w���k�y�F�Lk�С|y,0�#7�^t�:�lЍ^q9���*��Tx����;.^��&����)��UW�^�)������|щ��)F�g[$�e�����ĸ������j����˯�T�� �m��u8F��"��=)m5�j�/�*ڪ��4\�q��Y�q��bR��j�f�t��e46^��UfY�B�<��9��8����[�dk�_KU=CRjQz՗�L�3�5fͩ���!�%�����뗻|�/��W����E\���ں�;�T��N��3Dz�z�6����8!�}<��J�W�kؕ����W.9�.�=8���ݚ�y�Q+��N{��>�);���&�{��iu�oa��ʸ��"r�����(p�ŏ���̡l^īܬ��*qD�ޠy�J�r*����{�({��RN�ŝ�B��N�����Hg{�^��;�W�s�K�엿z��F��.�Z��W����U�e9;���u2s�n���=��<�j�� T��J��[�.�g9��gݛ�p���Ȟ���j�T�EF�Vfǌ&�T�cqby�S7&�y��ڇ��jz��V�3�+��5�u�&��>A3��}�<ʻ��Z�6EwՔ��S�ɋ�5�2U������j���2���(�w꯾��e����ݦdW]?!S���ڧ���=�y�iW5s�+�&1�]J�wq"j�+�7��6&,����7�+��V���Ț��%�����F"[6. �*N�dnf�&UE�];Cm�B���k(�Y���7�>勞d����
Se���7�b|}M�ʘ(D62�@b潮���vy4W�쐘�1���5�|p�wmM�Җm4��e��N�[���x�c8Ϥ�]�n=IqvjT֧�Dld9Pש��GTy'��wO�`{1
	(罸3w�������l���_x���^�3��g����o����؂�@^���L�LZ�n��ˋk����_%�iu/oϨL��v����=}$�jk�	��U{��җ����/t�]�s�-~5I=�]K��>ET;K��a�ݼ��vŷ!�꽜SP��>F�u�J��Y\������p+(���*ѣu-��a����!�������a�;��QK��d�K�j�C/
y�e
�'�uӮ�A��n�[�]���۳n�/m����_q��)�����Umԉqe��8Ռf#W<Y����:�
�(������2,�6�=����ݴ�-�~�Ӄ��Rآ�)+��a��Q�l͝܆�|1sl�'"��L�m��Ƙ��ۓӣ��u�����u�b>V���$�N�R^�*ʮ<kh����)�v�O�ߗ,�J�,�P��[ZƝ��ȜQ������/�ܮ[U�&��[D�=��*��ŉ��Q[�]�N��D~��Zʯv����r��f�ض�q5���U�k"ֲ@�������n�/7Ϫ���xn���Vk�졽������)ݜN�)9�n{���޾�M�н��m��Wm*���/�؂ܢحz�5��^�;Zb�q��*�`t��̰[U,�M���O�5i�tۊY��hŚ�1��
C!.�pj���T{�k�ײ� O/'|s�6�j�s*y�G��!绱Y����0ff���Dۀ�*�/T�vj��S�8��S��$uh���Z���X�V��94a)���u�>�.�*S��Gk��m�*���b�Y)�e�ʝkN*Ĳ�zv'���x���Z�Ջ+�V�:�c,�]����*��M��Y*�/���o��]w:���\؝��髪��B���noRΙ�oi�߾���C��p�P�0�mO��Y}N�rnۖw����E���k�:�u$���OW�5�ƹ�y��I�֮]�/r;T�l<��\^�����8�:�Px�߮d��1M����-c�����2��jSGT�yl���M5���cX=n{r����|�gz���Ի_�e7Ի|N�x���>�m\Վ#yʞ���W�!�f�{/}6�Q���B��S����:p���}*��� ��(|�g"��S^jճSZ��L��uL����~}�1ݴ��zwfV��� 	�e=�W$rwmo�>�K�}b9��ȫǶ�3���΁^t'��'��\���~Sܯ�΁_3޿n�p��r*ϙ�Q��T�_��cudiߖp��Y�bA���z-��|;���4w}9ׄ�qɈ��**������R����]�������w�kg̬R�צI�٢۳�C���h�&ޛ[*�j�<cͬdU��<�umj�qe��8C��4U�j�9��^T�w3��s��r��ͣo~R��`��_Co����������v����p������LKD���9��,�Z�z��,Q�#�j�f������@��r]S��"�ñ%e<�jv����P�me����s�*�o��w��gW:��!�a����	7�y��Y6��ÞQ�Pnz�����8i����U3�+D�M��3X�g���ߏy�|re��CD����m���Z�[�%�QI���P��͌����W���&/g}�=^�=��5�����⼿(�	`oVv�%�>�tW��%R����7��&g�~.�W���ӵ�+/L\��@�$��j�ECm��L�dL�;uVZʱ�b�i!1U�7пRX���a�*��o�V�����Cj��
�N����F0}��uK��p�x.Uv0v����Ŵ�����,�u�y�����
үz0��Y�B��-k�V	�)ܭ�|	P�l�rךB���]�ǔkX�T2Fbùbn)�kV�jJ}�R̵�k���o�W�+������!v��&%��d2kI�_Qa-�T�$4\|�k��(ԭǄ��'+�}�s�݀��q⬖��5Ǉ� ���_�[�^}V&v]wϵ�7�q7u^V�=�#f�����c����~T��ʺ�fnam+����W��>`�\R�&������U�P��%^��$��=��xoN��{��iu�mw�{�_v����a%,L�ɂ_����t?=�>�T|�5����<`W���;k����ԉ{��y�{}���\���y^��x��3��ty}�{��o��1����q�����z�{�򖧸:l�b�yƴ���=�Jk���<�y�Ӕ��T��C��Z�^���{��
�ߐ���qm<�M����h��o��{̫j)�}�]�;�?{xjU�5��Al5͹�ЧR�e��I_xt�h��'��,lV�o��бz��-�W?]��yS;]����bԝi[�sI��X���_���1�[�;e>@M�
l�-�(�1�YK����Q����=~�������^^��)���w�LTaKD4�l�X�+3#Bw�w�׷��� �����Tx�҅.��ޚ�h��Q��X�K�
�a�d��&�+F3I��b�W�|1����k�L�s,h���t,�D�����N`��
���uԕ��q�*)��rW�ጷ.��I�Wg�e�.�L�,��3�.�+t+ |J�G$���-��ҧ*r�j�J�s�t�������:�n�۱/�4���"Y얮�ٓ��Q��=�}IďRh�{�7I�����~�6�M�BG�e��c�!'�-�]K�O���<���_�ټ�=^�+S���X�7�����3��yk�6�"CO�PS�S]=�YY���9Q�V{|:w��]�vy&Q����\?gR��ξ�y,�˵��Ŭ�{�z���T��S��;�ƪy�4����;[y�5�-��K3�s;/{B�z���Q�,n�^�������aM�YUB<�:�pX�{��h���-�W��a\ĕ��L�wT��v�"u]�PBz���#w1�Ţ�~��n!����v�:�����q�&x9ݯ����qS�ڣp8�o�7۸�wSZˆN�yQ���ed��ӵ<�MY� n���"R���?{q�����]�b����ƻF�v���j-}��U�J3ǆ�W����bʹS�@�f`U�ve���tr^>K��)�JE8���P�ܙ09��˦y"=ϛ f�`� |STʬ�Nqm��[�!�g"Ǝ��+3��+�PQ�*�Ǫل�y��������4�;���Vv%�ju1>̆b�cyg���k���e�����U0��w{Ɩ�T.3S)��ӥ��M3ڰ!`�p��|�yф;���,&�$o�?_�,�U}���T���ʿv����r+2?�Yx�܍1��p�f	�6m+�/�q�h%[���t��4�ο3=���zG��5W{��T�,ez`�/k~E�K��]��Ymz$e�a�Q�U�3\�O厔��g_I��M�r���4�J}Ꞹf�`���7�2�g���{��Y�ſ[G��m��ǖ�ǭH6��mY�0��{���߮q���g��m�{�5�a�U3���)�/J��4cUL2�A4O���F�k��1��q�]�t�0��\Fc�z����}S���N��a��y,�K���"i����b��|�+��h�0���]S��-���N�y�mva�'s2�}���kO��,�w����q�J��\p��TG�c�~~��=x�]h����V�o)����1-�ƛZ�+�ap-����L��7Q�c���;�#�SeT����x_���7�k�x��2������!�`�:�g�둪������*Ǆ�]�Σ��"r{�nz�1b�����e�Y�M�޽,�����쉈�w�3{ªBƕa,{y~�w�q��ߡ���;��U�VUx񣳶���zkKӫ ���N}�}���s;S��gK7��z��ë��"��x��WF�Q��	aV��L�s�8'I�'�s/VR�:ڡ)Gv}E�P�T�,���gg�����Ǝ��t)�y.�9{���|�{ˏ�.��;^��̯IG��p�J��)���-��I�=]���׹�_����4�uk��^�/�{Ӣ�Z�dۡlz�^ܳХ*b�əa���3c���CK��(jǱ�1g���=38x���K{s�Z%wmxl�Ӣyf�Uڽ7&9�yY��1)�����=3��^���*	^�@c䪽����|��a�+v���;�ڪ�
�'�jb�Վ��Y\�^��g3|��i�2�����m��"v6��ڵ;dB�a��H�����m���~��=�w�$��W�*�%�h>������U�����N�V�'1Ƃ��=�9���o���m�g@��/N��� o	���W�"�mm�ֻ+ K�L#�dK����p�-S�Ò	{zܮ� �cNa{�B�Y�+"�e�yƛ}�{���J�}c�4\svNF�K�X�y�&{�/Q|���O2�f�A��{Ov��Uzy`����0|���e.����,�B{}\���ݺ4)��bR���������m��e���,x�!{iu.�<��_���cPC�ź�>�>b���ƽ�OErU";�y{�:ӵ��8o���r,�J�{z�s8�[^}��ON�1Z{�M�ם�v��9z���2G-��ǎz���h��/{�f�sS�~�>Sƭ�-��������PO�v���}��JXcd�I���4vy����v�����|�����!�꣖�0�Mڕ�	B:�rϏLv�'�4�M,����?u��n�7�ަOu��^�Og4G6�Rm3����]�ew��:j��oǞV�!m�s��"�P�����X͠�Ix�ӌ�ܢ٬�حex�g�Y�W���.+���gl6#�{S
�'m5ycH���cO^���f;�Xw.��c�x^B�0(��R���	A���=ѧQ]x�b�>�,�X��.�rK�*!�|v����p/d��m�$�v5�9��<��g�F����H�V������E��������L92�}��ͪ��WL3�J�)y��m.<M�I��75x����І�6�}z�s�����y�ͩ\�DZ쾙Xf���A;I\3��pRᇲu��	,5[ز{tݽ�O�7ȩ�����]���G! �3����I�o6�U�
�EG���S�Gvld������V)�W�ùW~��|�@@�h/vw-�i�1�{�R�/gv��nyӸ���ު�sc��&�{m�y0	�[��S!����i�r�]s�M$�sm}��5���h]�E�^u&�3H&�Dt���X3��[,[ś,grIz7�X��}}V����K��9�l�%ټ����k9h�Zl�d�Y���D� ;�У7�S��#X���T�n���i�K{u����k�f�&�YYΤn
I�]V�CX1�ID�ni�n��G�ފЇx� ^�ѵ/[݀.ݛ �!�u-6�P�N�^����qc+
�Оn�)PeqG��Ą�2�_f!3,Su8b�
}�m��k��9���釡��qV��X�|u6�J9���È��i_m:5�0����	P�qSmUgڗMqi{X��`�֘�=4�\���o+S�˫WC�ń��pA�vm(�F���Y�V�e��,�B�{�o�:���\��U�v��T�&t�}���S4�蔾�����J�y��*f���]#�����ލ��*o�+�c�,�f��7�t��[�6g��e���36�.j���*$v$(���72�>����C����%��y��|-
���Vͩ��7�(���'V�W���aZ�K�{H;�-J�eo-���қt��/S|6�v����d�ŕ9�N䫦6�L��;ݧ@V�Z�-�P,�Mb�D�Իsn��>�G� �8��s�q��	�m)�Ž쥋w�Z�d쇹M���wF����^U�ȍ�E����O�jz��L#�(��X3zN�[,9'6Yǖ��ͫ���R������\���H�iN�)�r���:��F�H�dշ{�[ԠqPgU3�ҡ� �t��]��I�yt�w�%X�����5&� \�V�@a�ψp�M�U�sgE
�+�K9S�������ܺXw�M���in:�4
1��%ןe�=���S��&����%��.��v�B��d��s�ٻ���2�#�g�td�w���;=����nFrf��qQ��Q�X[�n�<or�	�-�1����U��=S��ޕz�r��;z�`�)�E�I��`��4:*�	�N����A4E5C�kl�E5lj��5�lj�l�J�V]4Z��*�b���S�;j�T�'ZH�
J�4�6�T4i�l������[�E�Zh��"C���)��Zh�.�qh��b���X�4tV��*fh�j�O\K4C]	�F����i��&&kmRQ�E$��JS����j^�Cl]4�a()ih))���(i"hj���������
������t�f��(��bb����=�֩�AE��&�-���N���UDM&�3�դĕZ�t��bZB��J�*��`��
��.��4�4��ڎ�]}WW���,��	Jkb�돴�8߹��t;���ڜ\����ے��=x�C����'V^3��x�*�SV�^ƒ���������)����R]d�熡y��Qm�Ye��&5���*�;	>���5���s=^�l����N�O�b�t����(��Y�5�[W,�_b��]�$�
o��}���{ϭV��|}��B}�\v�V����0O���ӎ& ����&�K��uK��]���r�G@��ϳ�n\�6�!���;σ�W�ݧ;���c�+�H��ޱ����{x�9���/zsP�^��Ok�-�2��qo���i'�mR�^�b[r�����ԯk�Gs�	+NM��;���نWBam�DN[l	uQj^�m��6�b���V-k���j�W��>���]'�ߗ�{�\f�ؕ��g�kw���>j������=���t�>�/l�i�	5����E���}���)f�+�_j������a�9(��o�a�u��V�{qwz��vs:��fa��q��g;k%G��Q����f�xK��K��wn�M�uZ��;,=�X����,��n�H^�dЯk��9�����^��Oc|�'�#��7Ԇw�����o�F��p�q{���g7r�gJOz�"1S��ڂV�6.\��{�p��n�՛�Q�ہd+g����bU�ƴ��Gw�wJ��X|3<2��{;`��;���@g�>z'z������:�����q�&xi���'[�T��(���Jj���;Y�{}�q{8�ݴ��f�ؘ�����m�<ɣ�D���nnC���dzjWo�P��	�B�4��"��HWs>����u�����\��?c{�gj��_{}�{�����W:��eWEʮ�^	e3S�o�n{��<�@��1a?_y#|r���#ѵ����Z��mp�UA�9��R��j���^U$%o_�|:-C�x*w촭�{h\!����F�I�4�-�M>2�'%^������Ȼ����)h�e�s/އXD�L6��W�8cܹ�ܱ��K��3of�����5+A|�L�A[-���~�EF��[SjA���/��L紗�����,��gq�}B+�O�@k@��k�:MW�?X���k��)'f�ST]�gq0A�2��owh�7ì�z����+oJ���$�&�2��ǋR�x��=�"6Q�n�?8���"�8���Iu�?c��Z��N��2��nh�=�V��9e;c������{��㝻߸��S�m?P�gS�&�9zT�4��V��S��w��;�%���ߑ[���y)��|����3��w�I���v;|��5�O��s�jQNM���X�Wcg��S���V�>�O�*t�-���'Օ��/J�8!�~��O�7ݵ��;�X�q�������pn�ѳfEc����ۛ���;9S�,�R���e�)���4�lhZ�@�*��Wd��'\�vɵO�sF�s����es�~&�rܓ�n�^s'��w�<f#^�|4�M;�$�ޏ�ΧZ�Qݠۯ�,6*iw!De�LF�R���g�oݐ��=�MK����s���Y㽛m]xE`��r�Rp��:�O5'mYL��\dv�
&���z���e,���`��۾�ش��y�ٱR��D�2�����玄����SE�]6*��5D&�{!���udfL,�x���H�G]��F���֧�p3	�h���')|T�q.Xk���d�|��W��)Z�l4�.��ۻz��۞���{ݠ�d��MMm�T	��&RF����,��Uˑ���R����4�q����U}�
��������Q�?yl􀩺��2���'ϰ��x�FAT�������:3�sTsC�d���Xlڭ����le�_�������Kq�����@:Ǵ�;�XW~n��=[z3e��Ҕ������	ʲ��l��J�㡡�8�ym���L��ʉ���{vλ�h��辛~eZ^�����a�8�\!�6f8N�C�&߬���Ƽ��B|9�I�gݸ�/�tv�����u_�=����טX�5�S{�g�W|t ����͹?���� ��\"Ĵ��i�J�:��ͽF�7D�eFC����n�k��6Ϟ^�;�g��-i�p9��\^uL�e�ٱ���d�7�/�}��������L�P�'M;�;M��:���Ι�Y9�Ԏwd0Gw���~��˲岛�$�+{%#^踰v�d��W
�K���n�����;7ds��w�V�G	�aݘ(�%Y,�l-�ԄF����)�Iی9(b�z�K/g@�͋�i�4�(ok6D��#���iP�K�N��aKcǰ�u)���
z��=17��Ԃ�@,�q�e�זX��o���uwANcz�!����(�#���5���`���Si�;�r��A+r���ں�G^0��|Jri�u}N���z��Q�@1�֩�p����`��Kux���p�6�zqv�}UUW촳ϯn�N|u?�@�=L/��@��}Fi���%�)�J��L����	���A��ۗ̉�]b9��_
�o<{����5�\�*�.��5;%�-YP�}��+9Td��:��NHM���ܝ@��R�
c�SYp3nϨ�7L@��Sb��GCϩ���Yϕ�4����3%d�2���g]����⡸�L	N��	�����EI��C��%��غ���9�SB+����������>)��Χ���3�yS�A|�δ�;>�͐ﻚ�3�{5{7={�@Kj"z���xTk�<#m�L���O�)or�ۧ�̰���-��f9�#�Q���'�؉�Ÿ�d�D�[�����>�BƸ(o�8ӯ;�l��_cf�Ke򱍋Ffk���䤉����˗��i��YU�s�����\2�3O����>��nc��nrӚ�\�l�F����3�_��Hܧp��	;e>?�T\�UoQo-eq.c�P��H8�'�}��U�j�9�A� sf(tf�"��w\Оڇs�k�>����X������E��6�����z�+~�R<Q�΁�͔5>ǐ��z���q���Ft8�YA��{��Q��M�4��gF�v��15�:���州o����[��ޕ����۴Q�e��v1�Ws��R��9��=y�vQ��4D��tfZ4ppO&?��ꦲ�'71#W��k��t��a����Y�ag>t�n������ng5F�����%=K�t(�i�g����#�J��&m8��!�\�B j����v[�B�c2��CL�|�LX�=�\���=8L��y��L
&ў bM���Ή���O�z[yJ&9����'��ڞP�n�1����`*[-E�jw�k����/y��Ő��N)���tA|���c��M�m삎�d	@+|hװ!��S	�=jyf��5�+��S�[5�`Z��/�~���ߠ�y�����<��k���Es�s�S��4���@߬6����2��/�?�s{r�Q��lP���-[p���0�z[��v9��nΑ���eGL�3\��9�y�l�t�uQ�ƶz<�ͽ��߰���|:��܎��MWG<��������,yeDE�U���ٟ����,�����$[~�wl�c�'c#��q�r=�x-�t�8�;��M��ig�m]Uv=\읷�
��+~h���*�0��ݱe&����x�%?��yyB*���Y�;K��eJQ����]��]̣z�gm	��1���+���g���3��|:����.�}�=bHZ}�ᕐ��I$,``J����`���
��}9����euAS)B[�����H��7���|�[CV�Sn|�L�ui՛�q�9�_[�]95��?������m��� ϼ��rT8\q���7�^L��U.�B��sĪ0ղ!��ڶ�c�y�w���P����py�[p�>��r�r��.���ޚ踰�՗�B˹2��(x֦�ٹ�S7@v�$�y�g<a�Dp��7 ?~9F���6��2~n�G��6 �;�:��e(�����2�2��^.�·`�a-����\�-�̆�Πb��t9F�n�Cr��^�Z2*�[f�2�O�E�z7�O�r���Q�O�!9�k�neu����?g��|f�T㋆;����l4�e��%���d� Wg�8pي@�g�ǷT�=��DB9�Y�\�su���ji�W6I�]��g_��Vԧ)�Z���+�w�Կ���5gs�rh���Q�9�1\�Q~�t`�4�اFu;��#wKРq�(ej��Z��;M;�����S�}�1�%�f�v�f̉Z������=�մ�l�px�����5�A<�΁�D5���Àn:컼������Ld���6<�S�$E%gQVu�V�*m7�f\#��u ,����w���U������Z��OI�R<�]��-��('e�x��f�W7mu��čJ����w:��33L����])=��[�m�y�O�p�����8!P��5��6�zz�j���%�T7����0Π١���ʽ�x�Ǽ
�]x���d�i�jqwx7|׾�>��� T���yT�9Z�7uG#�ς�����%��:�Wy��P�z�ro����;���,C6Gl�5N����[5��	g��:�]pE�/�Z�]?��7���q] w$%�l�I���ŏ]/�:�14��)�q��di�z�Ko���s8k	.�w�/r���9�ué�\ŉ�wND3�I㢋��T�Li�4J��'��ا��c?SV}d��<ϑ@�S�e l��̪#��g�i�s�o�FAT���t�]�s�S]��9����R���k�n�Ϯ�ǜo<�?0���!�.�� N��0��df��U%^c�T�ɯ���0��c�[#�p��J�㡗��Ͱ�;���5tZ���Z�J ���1�_xbzw�m�kx�-��u�|��ͳ1�a������]���v^�gEr:�V:�~���~�ޗG)����\����3�+�<�! c���k�q�R�����W�]�W8y=��s)\P�Ta��tAf|�!�Ku�Su[�[Ϭ��aZ�M���e��y��Ƹ�y��YdU��.���r�&�oiTBfp����"�u������۔�.�D���i�cz�N-�$gN*�!_��{��'�^bc���:��t�8q��Kn�7���t��ڽE܊J}:M����m�̥��ܔ1n�����9\�k�=�n�"�\N�S����oY���L���v�^h������m�`�������.[+ݹ'L���R<���L�x��%�*l�7-W�7+,��i'p�f�p��հ�ϡF�>|��l�,���^�"y��ɓ�~��*�'��0�������F�;�%�Ȑ���'�֛�Q�gΪ4p�i�W�P�̸��iC�˪��L	���(1�,��+ϲ����@���g���Y/�O�F�b~��ѵ��h��s/;F�����)<��� ��5�\�B�a4�������f���5S��M3�ݓ�Z���_<mw�<��4:aB��^��$M<����ݷ3ڬ��/�N>�fn/�w�<�w��q�e���Y[�*[����P��,x?#>�g����x�K������Um[��1=A5��n�:�#N�dô����d1�/	g�t�ʎ�q��L._�����z2vm����BeTD�V���Ш��xCm�iF�������0/�n��yt�Wp�NV�sZ�gE�e�S�|M]���F0�a��!���:�"�v߼z���eAR������x_Ө�U�Z���������t�De&ڦ2�M,Iø+ �Xzn1��Ś�]�;Q1��g��!���I��I�l̄�ǻ/)ξ�����$�1�۷�f�T�\���?�~����)&�g��闧:�U��f�B�^Ȅ'�j5���a�8��g��ۋ',N�Mm�ѷ|��׸=������8䳗��i�]�*k��1eY/nˍ�� e����|%�� Ktok�0{6��<�,r�/ݶa��(V�FG��������e.�m�����h�9B�����a�&�K�3��|gֺg׺�GoTD����\�td�k{��!Vl�!� 2�u���gg�e�DV�{��,0���Yϝ.��u&Kkr���ѽ��|���<ۉ~9M�7���O7(�:.�A� W,�s��z�x=j���`M�_]>�w3�u�#�&�f�g�y�f7	V�Va���M���V9U�tH�[<�Ѵ@5���yW/�;yv�\���l��O>P�4�7D���]4O���2���x�;���D����D7k�T���z��|�ۏ��͵�����pWk�r}}��1t���}�U0���O@���ad��.��DX�m4ܣ5ma�����2�w����e��t��,r�P�f��>�S@g��t^�:��Z�<���m�ݾ��~ֲe-�\��=WZA�Ȣ�5�6cN�
oe�PW5��f_vf��V7uM���n��\�U׃K��wscR�soiO�G�f��m[��mT�˷Ӫofk��.r{�Vۦ��,��2�� �m���w�8�}V/�Z��m�T�R�x���-��}[�8��o���sԻ��w�S�a�t[0�jU�#"+6`d�^����Ɲ��i�蘥��JW�n�w(�1ڱ�c#�[D_&N�H�(т�6��o6k�TYpRh�D�ē"h}���C����-z�|<:�����-�n�K��o�:�T*\�j+0L8=�1�\���~�)�	QI�κ,�����=�ݖ�mc�s�f[.��F%��[���|��붜����i�B>��U|�	����a&�D�9^{+U��t�)}�� q �u�y�euB1�ԕ�L�e��T����hƀ�"����@����v:�N�ػ���Ƞ�9�"�i�������l�h���.��ŵ4�CvA9_�����\�=Z��h^h���Pԗ�!J�C$��Z���o_A��Нw[W��tZ���*�F�ѨS���g,��`Sn��>��[�*T�C�8|��ćNo'���q���v���x��%��'л<���GAǩ�!������S)�yW�s�5��izT�Mfp3-��܇J������Z�!ѝ�vE�k��� �;��<�#�y�����;ݖ���-��u�L7o҉����;w�/���2�d_d"\t��'��¨MXd @�F��K1є�ge,�@4��M]*:*�(#;��e�=-Ewt(�s`'���v]ǚݻ=.^l}D��e�W{e�C��30�hK�|;��]�5�����P	�H��맬�v-xRN��U��t�\*n+K�V�u��~Y�lpB��E�qw�,���Z�ŗ�O(���:�gn"$��姲'hтw0�J���Z��s�S��U�y��U��MkĔ+2����9Y��%f+�DT-�aa=���9�Z��C�)��oNyݔ�O�I"�JM����[��d����q�ִ�}� �����5��yT'p��鲹�2�^�1-���OgA���41���	t���N#��4�=�p���x��n���n�o�Zf�F�B]���sM�y�)�ɰ���e
ǞNp�ɥa�$s7�k~�Dּ札5
��Ӯ�k;;�:�
��tV(}}7o#�QJ>�VX��s6[<=��Ë{T��u[���d�'$|��J[������,���J�i��3*ᓳQ!�nP<��X�:�_��]��qw���3��.����)Xދ��h����o�X� :��pV����� hd�HgJj��ݾ�M�6JV�Y�W;ʙ�t,�ؼV����2o�:�̯^Z�2�6��p�%�Lt�]-*��}�����ԭ�����)�C��%����-��c��/548y��×zNi�v�)[��I��N�7��r������G�5	E�&���%(�J͡�4!A5Pt�*����&�Y��
i�F���TдR�RR�D-��5Eh:N��H�""���
JF��bfbV���������)�I�)�����j"!zBSDPT�RP4S@Q]�G]ڒ��Jh��"��&�ihi	�h*�(
i�����JR�d����


�Jii*�(iJV��ICJ�	ESQR��@����A%h�U)ICACKJPPѠiT��SkCBD�4% QHR����-.�AT�M+Qlbh)J
��(�
�*�`�
�{��z�.픣�KFqz;b��������K��o�z>�F�"I��j�!9�v63[����o�A������с�ٱ�ZorX��.���=% �#�Ф�Y�:�P��m�z5V^k���t��f5�������
Y߰��8u����
Z����y���jF����c6�����>��\��,�
��3u�������d`@��q���9:��O=�e�i��A���]>���p9���~�<��:�b��G���Qq�b�N�8?��bv7��C��$N���Qq��s� :{�@�iU��p��03������iV{1*�X��{�Ǎ��@�]����� ���#���B; G��G9y���D��b7}98:�ox]\�t��[�ǂ�556�����7����lc��:��r���3�8��v#p7~T:.'�g��v� ނh"�i?�F,����{/�Ns'��g؟xk���i	�c+�~ye�1��CFv�����;��|�=���o�T�\��Y���x��m��@�<ӧ=\�)ͼ�{��'���qMU��QO�1H}��h�>C<���e�q�fӁ}>���b�ڞx���-Og�q)�cL�Y��4Pihu�>{��GT�!uɕ�U��tLn�5���Y��jwZX3s�l�zg��|��ur���l �����M� �\%8"�#����)��][X����xvg���6�s��[XqZ�r�R�2��M\�\���:��Y��N��R`d�sD=�ؼUܻ������U㙵f0r��/�,Y׮�"��3ϩ��嬦��;�0�&�����nTt޶�o^]��Gw��mdn�C�h�V��p�g�w%L��Ń�62�T�4�i�nY�ql����+�9럙���>�2!����4ҝq*v���q��!��QQ�=F́~�/F�Wh�/��ֱN�*#��	�u��BO�����l�,}�,���}����L�GI��rs_�-U�5Ns0���6�����eQ�@���/4����j��-��NSvA����F��D�iYx��t��],��湗qq���ʍ�%�H%iy</U����1�u9;N��v���R}Ω9|Df������t�Qp�����x>��M-{��e�s��ٜ��<r����[U�ti�<��p[�R�TBr'z%����h�"ẺlU0=���n4+��}y5��G�.��"�.)�y)�u9ٔ�"�|��d�gd>*�<v\�򩽺��YQ]P`s-~Ô
��>�#9�a��Kq���:X������Έ}�~���B��m�&X`�Ӻ.d�4E��f�&���_�{��uk=�۴lt��6�)T����[՛}:�%[��(� #��̫D��^�/d���j7��ޥ�lo5'��v�|�Q�{�Z'��C}�-������3;�s
�{�<֞�D�G�x%����t��\�,��]��j:��;w*+3�I�����3�2��<]�W/�q�>�p�m��IDZ��<r�=@���E���z�b=�{����ᒃ��2[����X�qe��8����F��w��~�~��dfu�u��Ds�ƗT[�nב����r��+2�!�O��)���-���պ�o��m�� ��uu��:�g7���y�'�����7�g�#0׺н�%SŘ{���1��Sv�T�tw��c�ys�זl.6�:X>��wП�=.��l��F��)����}},���T��Y���V=I���zf�֞�B���"5l �
5g��k��N�����b������O����j=쇤q�E �Ԙ���S���2؞Ev:�p�GV���{d��Ҥi)����#�S)�����9��>�k�WT�5O��S�Md�8�t�<5l=N�i�=�,.SN�nW=�]0K���Gn�JO����^hׁs���O��s�K]4��hjU�4C�^Cw���k�rtԩ~da��B���o��,�:<�a��.]\*J�;gk;�{v9��1Fب�LL�X��m�%��k��n��տ^[���¹�wz�ltk�Y��>���.��4�������ՆdVw{ ��z�9@�3�y:�\����ۓͽ���e�q�Oq�4:aF�z㠪��$f���qx�4N?LwL'������N>��(����i���g�Xg�{	�*��SҢ�x?#6��]4��]���{Ν�l�K-FqܔءLƲ��������q��⟎>�~�ܵ§��FuSx1,�vM\�U�����,��"�Um�A�R~�P���'��}0y���p�<��,��պp'�3 ��O0sڐ��k�3�CZ�x�[����ŕg�r�І�s+�KU�*�Os^�Ws��I� �=�@���ug۹eMw�,�%������ԌJ�~{��1u��F=�l��>�݈|3i��etE��n$O�lÇ�P8�5��)�.l*����� &���i�ͮA˿{���q�ݠ� +�~5����愶K�����[��p����к[����'y�Ћ3|���ڶU0�~�vٰ�=6NW��Ѡ���{ o`���چ�/\�������<l��GH��F]�I��ԶC��l� }S'�+}�/���vX5'�Y�w�,���.-���)����_��U�g��6s��֜�C�vɶQ�uա.S�*.��~#�J� �wg�ל�s�+8b�0qo ���Ƭ��k�][�M0.��S;up�ێ��5��aY��x�Ŋ�kV���C^�Úyz�_^��Pug�Cݓ���1i���s��[!�9�"=��P~r����CKVH������v���X��ٮūw:%�fV��&��4O��=�;(��ܞ����k���C�g�ٱ�nQ��!"�o��`GR�a4���6C�W���&'�_��P���K����4�,�#��������w8
7>�	Tl��=�r���1�Ʌ
¬OO=@ss�Z�#���6lf�܅����]ʹ�Bkvt����s�Ψ�/�7OWX�+x
��q\̢6�)�>S�;X����~�:�8��]M!<e��=���=S��S���l�o{���4Ŋ'�00OGTЯu��������(K��2Ǟ��	�@��U�q�_^v��{΀3�u�8�ڄ��u�l�7�ށjƪWQF����;*0͜��;v������`�������������EG '�z�\!�~x��w=<�˹�*�a�d0�}��}=O[]�f:h�(ݘ��2�x϶: �%�z�L�l:'��������ؾk��Qf��FLPN�1[�t��3jM�U�c���Q\�U!�Pp�7om@�a��O{�y>�%��g�s�^$s�/��m�x��-��W{�ݳ�x�·ON��s�SB����Q�,j���'�o0�=�Pgr���r���;�0br�v�{��J�^^�M�����5���'�婞|r ��^�q>��
9�I&��̱1��TM-���荲���l��^�^�GKp�p��+�~ye�^y\�g5���a,��U���^��4��e,����Om��.����Bsϑ�bYBh����)h�36�@�:��v��;����,�g�]9,�_`��r8p͊ u��M�̖��d���W��e��Fa�O"�����)\9^�u�	t�)�i����a���{��U�l}�}����͙ Z�~.�
G��`�γ:��KY?N_�,K%�j��S)���Y{q���^���n���ׯap��tȆ�ڟ`ԧ\e�V�]7vI�}B2�*Nϣ3=[Y�cc�5��M�N��>܋�%����~��`%������,�6u�l2�i�(�H��m\�sallȘ�{�Շ�8}
l�R@�U>�y�H���F���G��,�.��{	�i�Y!�^�˫���m��gCa�}e�O���hفb[!T�-T�K��}Q�P�~|�Y�\6�G��B��X�ʥ�K��y��	"��4�z�z�C����!W�;Ɋ�
�GV�S����v�|�EA�)H��j����9}6�.���.�Q��Z3���GS�U���R����EZ�Yueb{"exZ��ޗ�`�Op��}@@��fnj���U2㟶��^�@�U*`Otq�VI���ՏM��/�� ���=�~
��/������Yqn�&�j���:l�RG-�R��D'#y�7����T\q��b��\�m<�Qֺ � );��;��%qNe�t�̺��2���%� Zg�cx��W���j=1u95�x���:Y
�~Ô
[:�����\!���Q�@�=���A�5
�wRȌ��h�E��v{Y��c�f�{�����#�㡡s��m���BxE͕�w4�������� ����7U�,�]Ga�����!�fc�뻢3nk؇'u#�Oo�<�oq�S��`;Zg!i8f�E�+4��+���+�?�p�1��T���[{�8�s'z�'2to���u<��.�i7D�g�2W\d�o����9�W�!�{���d5k�+�o7���GE��m�8�l�<}���ˮsM3*r2̷1W�k�"�+�˭��½ck(D���w�n�tɎd�|�-z��ϰ���/]o;�G�>.˖�nܓ�U����욡�K��{��J*��:N��nm�R�]G�Q<V=����r��k�z�����{-Q53���D��\��1�j�e���#{�<`[R���*Ie�Jӯ��s�u��]���D���ócT&	\Y8B�+� x֜ܬ؝�������N@�����_����!��~��J�c�Y9$Ej�A��t�)�����yW�Ꞙ8�i]q��޵�gM3�E<�t���N���S�Ց!#����Xn�߳d���MY��ѷ�����PᦇC^.�(tð����� KU>�D���K�N�\�����&&B���Μ=�ݍ����\�1��L"����:S���XI���s���8�m���9�i�k��T7J��3ea�{��R�	���*l�	kv|G*: ^��1���.�mV�^Z����҃�:�7p�>{��}ǰ�3��P�����c���p����z`�9ssw͛m�"�6H��(�Fٻf�̌M��_�~8������x�m���XG�KVU�D�U�������֙d��;)�.H�T�"�~��Ш��xG��4Ϗ8�rC�a '�q8��y�^t��ˮ���ۙa-����&[{q�,�蝋seY�l�,G��3��X��S�뤰L�C-*���i�����3'��t�y���9xF��w,���9�zʲ^�foX��to.�һj�`���mڈk��Յm>(j@�Թ?��Q����XӢl`x��my������ �y����R��%uodb��N=&�ڒ�tZk��x����"*v��l�y+E8�����/a��OW�4�{I�Yۍ_G<�[�H8���wk���^�y�\χ�f(M�C�w8��t;�=����IXkϏ�)�("��m4]�"������AY4�lVn���dtqw�Y�#��t�"�w��Y��hd|z��E����$�O=�X�=ɡ3��mI�/�E�����|Es�@c�ag�;{�Y�}.���{F�DV7]��c;��U]�=�捧Pڸ�<)��$�Zp-NC��t �SY��µ��_n����y ���׋}��Y�{����s�읦�,,�S-����5[��_<x�gE3�1z���ԇ���=L�Ӕ���}\���̍8�%�ej�Z��3�w�wl]�׭57 3�X��w��m�4'N��R��U�b��
;^�!K'�Ǧ�{:�S�H� ���"�+z�s*��~��_ �Zاh͕�p�2��%OG��B�<� Yus[=Қ���C�vɯ���}�����ׅg#�o!f�aj;p�紊.˧���\(<6oX�bm��Yǣ���1e7f�d� v?C��~�#M(��O��d`S�~Âw���{�Or�'gʎ S�
%NE��;5an�6��*J%��?U�O�[Vp:�he�����\ڞo+��,��O�+v߻m�����)v��5�c��7�(k����M>����=G-�'�jr�3�	�ᗙAZR�}�"�õ9Z���s����߼[t��?#>�g���P����F�i���t{0�;����I�^���4ve���u��:A�@�[,C��ya-������Ǩ��p�T����V0vTA�F�ǆ��X��U��e���㠞[^8�� ��].��w���n��附�v7�f�i��2z�;6���g��_�dCwsW� ?m΀:}Ơg���B���;�j6������:�7x�B�1��:Er���n��xk(tle�y�3�0آ8u#p7~T:.Ѽ�<�u��Ǵ��4����[�Q�2:ζs�/n���n�T0Mo��>d�$c���j�F�ض���u�7gm������-�e�
t�fm?y�@it@Η�2H�wS\�-n���t���g��P�3�OU��+�¯ہk�b�ͯu5�C��#�U�b���[�UE���W�b��/M����Vq�{tS*s��e)��h\z��3ϩ���44rr�4-��K37��̝�\� ;6��.��R9��S�3��޺���Ń��3@&fD��=����)��~�zn��cOZ7]cZ��WfH�k�2'w�U`�x'sD:c9Z��|���̘s������m��"�;;B�V-rm�����C�
jW��x�t7�=[K��2Yw��L�x;�@x��	�����7+\�ڢ�$�-8��1h�C���r�T���a��;��N�Y3Uld漓N�%9k��B��f�ٻ��
�ً�����,m)���+r�k���e�1��5�ZU�2Eoۚlf��w(�}�@r�B���ʉ�z����PE˂\O�s
���*��yRWm�Q�Z �+�ĩI�Vf�p����f\�/�z(�3]*��Ik�,grŀD������<o/g�*����=���P��㭼�7@�_i��K���ob���I�{�R��دv��:nQo28*����Q��;�;E+F#��(��X[ٙio��ݷi�9��^��)ź	��/����J#Y/��*}� �B'w�z�%ͥ
���̼� �7چ��J�K�������Q{��z|9���Vč��.qm���6�V^�r�)�w&�b���/�2�V��]su��Dg8��i�k�ն�m��*mLp=l�^�i�Z�,���H�dp�==�s�"�Y�)O�2Pgp�ښh
H���cDKWϥ̶��	��a���j�%�C}h�"W�@�����wa��p��M��s��j�`�V<�E�*��)*T�$s[��X��ӗ;M���/v��K�eM�� B�5J�$�)�w�����=a�|�lV�Ryt�$#� 2�4���=$�*p�ygWKk����}Z���)Dݫ�}L=g�ڼB���]�tn��FB �sY阂g��!u��f��ak�Am����s���-�vBl�v�b6��Ԑ�;�,��hޭ�V���/� {f	�{�����.ȲOJC�ծ����lt���:.�C��Y�2��h�$�7�b���߽�+���Xy�f�T�aw8#�*SP4f����E�M��I��d7�zs�z�zv�3�&� ]ǛH]�#��.���'�8� �@.�n���M�A�T�W�����8h��y�V��ܫ�$�:���U��0��`T5�J�	�'�`(-g��d�v�h	ŝz�U��Z��ĻE?��eu����,wk�\��ML= <B-��\"�<��6��X!@_R�a&T�(Y|��:#ʊ���°�:�Cݠ�3$�C|�ݵT�V�gb���֚,4�a��+��^�}�*��VU��b7	=��a��@1ty�b,
¤���)*zz*9r�m�G9����)�2�e�#{2	�����G+.�.Oo.ݹ��:U� Ž�d��:�R�����Ïr��1���+#�9˕a��]6����p@D�S�="�+s���Pr�:�,��,W��Q�!Y�-/rǁ��i�t8Q��i��%}9{�5[�lі�v��� >�τR��HRP�S�M%UCCKZLAE �41S�IK��TE��$

((��Bj�$֚R���*"���hJ�(4U!S-4�DM%PŤt:R�IT�ES+�j��(�(
P��Z����N��)h�(	�()��
hZ)(q	����F	�Z���*��)
���R�-$E4� ��SUBQA�"h

���M$UAT'�� ����)�E6��P����"CAн!v4PSE!���U=&�������F�:t��ӥ:4�_g�}�aY�-�&�S�k�\�g&�W����Ñ#�g�L�<�c[�[�ڃ���oU���M����c8B/�E�lt6(�\���Ǘ�o�{1�v�w[�M��R��#Gj}����-��x��È�^��6����Ǩ���x�/�5�:x�RE����u������BE$�G5:�.�e�v��%c��}3sg�fg�-�ݢ:L��� ��(fʅD
��_)�;F#���6�RhM̺,�d��ͿCs��]7L��uL�1H�TBa�m��6B�Z�֗�S�[O�P��e���@t��#Ve�I�I�r�(gT��-�e�Yp�� j��.+[#��Q4��"9-�ാ��8T�Zj9����m�g��2�y��6�#����S�E��I�x��n}e�YQf������]�ڨ���F����od7w�d�)̲��6Yuˈ򨎂 =����<�V�.�5�����^ҽ8�Ⱦj���Z�F`����Xy��O8�t�y�G�26�v�Ź��ft<bYs�����t˼F�n��Mocŧ��9.^	B5�CB��U���� U�T������w�ܰ�K��I�k�4D�uռ]�U��2�؟x�C��q;���k�g����]x`���]Ekr�CX�,by�63ʝJ�;���{�T�Y�f�Y>�&�>r�J驇Aɵ���S�E�!�
��U��g5��YKs����(u+
��Lê���r��>���;�"fIM��y��ɋڍH���-�Ob���������7=-�*�m���X5L{�j����_��tv>�� svM͊bk�W���E��]qB[�|7]F�O��o�r�������6����j�5���<���*�z �1�V���uF���|<�����c:?����#%�v�G��雷ӼD�(�1-�w�v�_8�y�s�X;m��w�zӮ��Xݹ'N[u�esQ���=3������{b���"��I�$�+���U6;��� _�l �УQ�H��q�Zm�C�m��;s�)�{��m���s:S�GM�
�Q�4��;���#��Q@�6��DI���TN��6m8�]���h�:���2�0�T:e3>�[��'�O��S�J�P6��ˬ���.v'w�a�͙��~���0��i�j'u�;�;�qV͐��k.��Fch6��Un����By�~Nݺ�꼹n���1N��i����zxSt禋���zݝ#�%���~��|�終{���P5���Xrn�^�a��N�V犞���ӝw9�'�Qe��Y�v�ݸ�<8��I�|�R�#g1��WF�dДb�874��1�?g=.r��{D�Zf� /"Y�b��<8��>'�5��S��oN.=����̲g�}���D�?�{g=<�ڋ<A�꫱��"�J��pl6���m$��J�/��g��M$\{�M�iFٻq��|u��6�S�خn�k��os3��,�͇�-���@��;ǋ��rE�j�six
����x�Yǻ6�FE(���6PT��@t�u��\e	K���|�u�̯�i5�]�E�a��d!b�y7M�:�^bZ����s��\�'���.��%�t8w]�`㤕U�5�s�̭�/7P}gq�{gyA/�n��1홎ͮ�|�?]c���m�f<r��aw��kP�i���}i�����
BR�G����� ��-�ͥ�%��=�";z� ���b�aS�X����œ�'��e�k��*�oB,�_8�yl(u'�����,�U?-��Vnp�ZG�8w��)'��ql[��j��{�h��t�Q<*��L� 3�Z�}��ޏ�U�X�O��it����L��MJ�����}�-Сa)ݢ��1i���W8�!�4�<�����u����Q���nk�~h��=^m�4SgY�|���2����7D���T�H:�>k#���ϱ&fe����/gg��nM٨� ��g1�����v�����9uͅ��aS�0猼��{�-
�z��nlܶ5u<�1���e?V�ƣ���ƺ�=�h����S���.��q���;���-'���p��9v��o��� �qc6_|�m��nd���~c8��\:Uo��-Gr٥J%��f�׳�#��� J�����}{f��2CU٘���Ν��Û�3��	s�KqNі������%OGc��R�!I��k�@����a�"�q��&j�l������l�gO�jt��S�Q���-��
Öc˧���ZKf@��zݱeU�f\?d����u vlC��dB�B�ҍ4���>����~�;ZЫ����H�CC7��?wH����t�'ڡ<��,��۳�Y^��'��hQ�[ov���s
�7���u*��T��΄y�=���UpMw-b<��	��O>�p7��õ�R�� .5Q������'�nFe`T���N��_���~ nw\��\#��/#8���4�]�u*��p20�D�>E�;��o��z��-՝{y��3��!.r��.�㎂o�$^1Z�u"�/�?f
�ox^�Y.m���!������N�;<���N�j��|���{����y.>�g�9M��-�(v[���>�p���nBv�9��CU�%*��Z����a:u`փjд�*��i�du��O��s��k�<����-����q�7�Z�t��ΰI�G�W)�Be�0�﹬�ۘ������`�CM���)��G���gV��#����������wQ��T�l�ށ���uA�d�8�Λ��n�f��5�řkO�[! �q(�U�f�mv��v�X[B��UU7���*���<��*�k���(�g�-]9,���dͧ�6F,�D�)����61X*�lǞ/;��U6�P�3}f0JWW�"ŝzn�"��3�!����QړC'�Dm'�#w2x�?2<�#-��\�@��Qz�dp�k�ا�bs���J�TX�t/4p^:��$4_����D�o�Y����n�l.Έ�{S�f����l��vI�g�s�b��)˿]��^f�p�3dTpǦ��<�4��	�u���BS(P��(�j��*/'&��S@�T32f�*���gKu73��}��ٰ#*'�O�^Y��;>����j�цg�K.�U4_K��KQ�i���磜���=M�m���I��ï#f�l�R�S�/4��N�L�ǡ�m�\P0�t��s��ͣ��9_@;�zd[s���/k�V���6r:�7D�t�x����;�����;��a�2K=�#><�Kj�8)f�q��,��x�-nϨ�p~����^Moqq��ǆ7�Y�-(��.�(L�%4^��}u���`��e�MX�*&�e��Vsq�6���bʼ����TyS��z��q��5vvp  ��#��m^����U�;�:��Y+\���#�`�1,N Q���JV��؍��o�9�|�g���~�v���j�x����n6黎\S���>nPC���0E�7P-�m�qM5�r�p�;�^���vv	��?a��*��,���5�X���~a���H�5���8Nf(���B$~gZe�"»n��=V�1ͣc�28^�%
�/ݓ2��|��'�/��bF���`!�mq��_)�a��Ƣ첦��È�/��\��M]��q+��թ�O;t��sdm�r�t@�4̞�D�X��g�O�e~�t�2W���oz~10��a3�V_�j�6��0 �����m�?k�s,��;��M�y��ٟ(�{RC0V~�v=���`��OI���6�3�<����.T ��<F��h�K�u}r�yS��z77���Ȫ�,$��(�̅�;EM�<�q8bi���o�Zyl/��0{�O��Q�O+��e���Z�P�ke]�����㧻���)���Z�.£Z��jw�*��,���#V��3C$WW��a��QG��[-t�ڲN���zE=z:lN���w�f��ަ�D����IF��i�~�gq����wU�>w�9��甽Yb��K��D\EN�������Gn��f��1r������FhS�����#D�����g*��Mno	�ݚ􅜳����E�@M����Θ{�&\o[�%%]Or��܍��\����ݬ�*�z��BgoB�"q�����G���w���7Th�:��R�0�|��)�Z�GWT�5O��\��������&T�����*�F�'�1i�fR����p�g�(�k.~'@V��ׁjz��Ze�d�i�˸繄ö�qyf�n�yjʆR�Ѻf����7`{��*P�n{�r��e�H�8�A������W3����E7*8��+�F�
�H�yju�n�z2{Mxv�S�;,���.�}=�ٹ���1ט�{�Z^����v~F�
ޠ����B�(�7`�ُ����5�J~8�:�*�t�ӕPZZ��;��t��ˮ���O	��?i��g��QrE��R��2ԟ��&�c��R��X[	]��ة�0�S�O�@�n�Uq��k��ت��8Kt�UE��k*�CBE�ꖠ�u�5�:�X�n��#1�\�oKk��I� xn]$L�H.:My��Yu�~j�-l����{QYh�c��#�K�\7#3Kn�?�p/��DXu�۶�8xnP8�2vn�g��u5WO͵5z:0��Qscjޢ�l�%̈́dt�KizD	�~�-}a��$c3C�4�Ղ;3;;|}��s!��8�[��2�Jx^#�&S�da�qd�oI�m]ۑEi�HGX�.���Y��x���BWYS�=E:T�3�˼'�w�#٦� �QZF��Ns�n�4<���]%m]*/oa�n���ny��ڭ�j�4̽e�+�F8����R.�?��c�~�(]5�^�zfm8�y�l)aLzy�FnJ\��`����$�eυ]�6m����ʃ��C�;��	���®�$� Ṙs��i5蓒�}�y7��Tf��.Z����s����,,Ǖ��M�Ʈp5d��X��6*��b��q`Ѽّ"<�vx=z���\��6�}5�/:��4���#���D���굕Pv�j�.;vGnN���~
qD�m��w.T��_�f�y��
;M}B���X�s{8��/��B�	=�ͪ�Q���QtW�K�R͊v��c�+M������^bܒ�d(�&
�3���ok��<�� Z�D8��\l�'�����H�<���Zore�E�6�#�lB��O7SvmM�F=sd�|s�Z����e��c"]�-���b���69���u�b�~?]��?A���#~랦�M��O�]��׋=C���4���:/(�9�sS���j�ޭ(s�����Q�o7]�8�J�e����S�j��V?���n�AW
(�T�|��&?��]ɲ�9֞�u��u*o�2����j2��a��u�Y˛��X/�����
	�{���R�Br����N���[X*�v��\d�Bh3;B��ֵڑk��暜*r��3\N�nWE,m"fF���or>��+����=��|S�O-� �e� D�Y�HGq��F��[3p���2�걹�=ڪؼ{��'��K����{
M�e��x��@(��9˧�w��2�Ve�N3�Zץ���P�w��n�ӓ�U��x�B˼z����I<�L�����ú�`1Z��s)Kr�~�Θ%�8�Ǩ�=V�>Üp˄�#��N�N��=�uJz/׆�b�هL_���_����J�C^u��5}-�F��Mv�f��on���-��f[��v�ʭ .�� �G9\`K��b�)�s���,�e��+�Yo�0wz�@���?���ݯ�i�#;�p� �c��j�·�E��_Y���Õ�,��*��Q��Ҫx���v�4,/�lkGq߅�t ��Qy�(�h��S�����pBM;�Y}�Y��;%�b�F<�3@GZ�h�S��i�~���]9�4�>��N��3�l����q��A穙��fﴽq�}� F���'�ٰ#�P��jz҄Ӻ������$RO�bh~묋^�N��*���B�ˊbۮ���7A~�2�b�yW��|��Љ�Mu�{�y��s��b�D#��g����~˭�Eoo��M�����V��K����A|��|.j��(ľ����Ϩ-��Cz�k��}E�r�E���gY���Y";CSNf87�o;p�?R��dn�\#��u ,�F́P��5O�^Z�#�o#��W�2 r�%sK����C2w,��܋�@�B�Y�n���'�wL;)�f�u0�S�._S>NGU�s�={r�b���Y:89�S��LݒE�f�0we@����X���.�=�1��\��kf_TEO �����Nd2����>�|e��t�Т���
����օr��=1��/�ۮM�9̫��0ZfH
N�d7K�F�%qNeG@+�\v��u�{M�j�v23-�{+MjPG?@L�y�㏎Ę�06���P����>�F?@~yV����*�ӽ��������!������Y�#B�n��=^���b���dp�ׂP��~����^]��N������_<�C�]L��ʉ���k�z"e���]�Uw�[�.�����Zjj0Jٜ�/�z���n��֢����=+�dc�F���=i��FKu�{��I��cۈM�gɦ�'f���d�C�Q�w�<�h����[]눝�A��Kӛn�ʌ>��6������zhe��9��pf����y��*��m˹2��+��kz�Q�Ť�������pj�	nLn��[:��0�Ԭ�E7\���hܡV9	RG�w#����BnF�ۏ%���+:h>g\�X]_�(�X5;�����GG� ��b5c���tR�jȑW�u^��g�Z &}+F��']�p�.O�\9�ұde����E�o%Jz6�Y9w��౤V��p�1*F�H����wu@��
����H�f��qE��q�T�m�b��t�ZD1�-�ơ��}��L@W�D�uN!�G;`��B����W�lCWtIn�˞� �w��G�`�DN�����E&���]��ު��$x�4sim�C5�h�;!�v�\����Ks�i��7�&��n,�vm�c��oo�J���
�� �pv��9�����AYtЌ�{�.�ٷI sY����jy�s�=֌�i�'�v[C�NwH����p���xR�ݫ��9CFU�����8��1~)�p��lL=���7R�b	Qպ��Q��w��3�.��^�M����h�K�!�\p��� �لK��m;�Kṃf��ۋU{�&�G�.�ns��sq�Ve�9�gt�g��)�pbg%J
��)5����'ON�*�!Ưs^�oU"K��6xƌ�X]�m|�npY�2z�kV��Æ��{4�K�vMyt��]�P)}���R�����>�9z,X��jN�g3�fM��E��������I������$0`rjY:��}��X�'�rYT9��wcQ����]*_e+��C��(�++Ņ��c�O�*��L8,��7�#�������|V�%��;�>�m���Z�yW�N�K(mee�F�2��e��%Հ�����'��i��CE衋���m�@�8��a�y?Q������wq��6M��ք8oA[V3_b�m[�C�)�����֮�9N��\�s_ǃo�Ψ_J:9�é�!Iwd}��d@�3��:κ�Ɣ��a�����)��:M��2�#r��5:T�h��˴���H@��Tb�p��nƾ�W5RJ�/wpuu���T��N>������i=cw���j%��C�$�E����c����s{�:A��I�"Ӱ�_RTaݫ+�κ��_F��W����t\�c�AazɶCc@�5���Va��+�'���]�m=�w{$I�xk���훈����	���kh8j{������-�N� ��ZsF�]G_j����zh�S;S[��ٙu�k!H��O@���@0���f�w%����]WW���F���9���^?��Ƒ	rm����|���jN�z��'R#r]�Y�*��p0�5yu�����o[�:��(� �)�)�)H�(���h��h�):T�E�: ��@
hhhi���MC��(zt��RP4"b(����::������kl���(*�4i
�@��IK��U@U)II%B����H��4EITąQJ�j������%�����'l�-Ĵ4�$�Z�%)I@LJQM���WB�F�Z4	M-�4�P�QUZA���#�M4���i�6J4&�I���R��X�zE�V�iM� i������:MHRSIA�ACT��(4Tv�-ST!�(��U��q�X�)�殨"3X�:�u��r�Ꭿ$�s�GjsY�U���)X�5et�YMb�Գ,ʃT��qb�FI}�e����r���{¸�L+��o����7�3d�k�cM�g�[u�\WF��|m���!A�͓5[4E��eq8b��v�N-<�aq�,إ���q0��=�[�����+�؎0��3ԟ��?~x��������Q��(T\O��Ѣ{J�B��$V�@�>L���w��vo�>B�G�^�e-�����;�2�y�t��N����c�4��3�@��v���d��yՙ�#�qM��+^�e�a<�t�f}���]R� ��N+�̞ͺx�'�y;��9��t�b~������t����$��P����ڝ��.(����ˍ����O�#��;����s�ӷ-yjʆ[Ϻh+=���؎�R�7=�9S�����ꮩg�y��u�����E��|���#��SH�y�Xf��q���N�V犻�0�k臣��OU��k%��]���>S�8LT���]6(W�(�7`�љ:]�5�^FV�m�h���oq*m⦯��:L�w?��wL�㠁/��O::�.H�J� Ϛ��̫�Zh]<B�+x���fQT<�4'���Xb����9|CI�����j\�8�r�eSඍ��Xk�i����wTB�>ŵ+P.OU�zJ|ke
���>����3]r颍yY�%�w����97����E��(�S�Kjȝ� H�]�T��6R�&�|Xg��E���f�M�������}[�t����f�4�'�s�l.T�J�0����艖���Ktcӝɾ�������|�U,�ڶΈ;	�P��G�9������w4�sr���� ��=�s!�L�P�Gk�I^�U��VS�D�z�m��']��������o;pÇ�`-�v�uA�=eg5=��v�y�6ʸ�����-嬡��&�Y���Q��?����xZ���آFX]���/�9���Y�t�i�8U;՞�[Ћ6��|l(u'���e������mn~��~ިky�����ܬFa��4oi�H��]�I�N�r:���9�ˇ�ظ7Q9�i 9UT�z�XT�E7�/���}��j��hR��2�SZ��=`�Ȟ��.,����Uךx��X�d�D6�����cod��i����f�	�C�ӵ�k*9T�6�y������u��N���7�3N�olwANb���V���C���ŉl낊���!5\�.lP1�؋�F�j������#ʕS	jz�yj.笗d�اh͕�pח?a*z8m�_����Y{�
9�O\{ bݮg�P���Yu0�W݄<0�>�(�����(� ����"S<5l���
ᑋ���!#=w3��Aԧcy/�c|uht��bl��M��� ȸ�\���3t�򱴨*L�K9H�^��T�]l�sM'�7;S�+�a5I���؛����~|7��P{�� YMɯ���j��
Z��L�cӖ���Ȱ�w2��\O<Y%�����FTT6�}s��p�GL�dB�B�iF����vk#Rܛ|��dw�����\�u啹�*���Z޲���[��YQs���:��u��V����gMSC�D��'��/��#�Q��e��9��T�r���i����v�E�ku������̾����;����p~�od���[^8��� C4��p%�;��P �F�y�n���b��z�����6�g���Ƕ��r�s��[y��\� M�Un��U\<8�W�Q+3M��~�,�N	c��t���f��/�Yw���F��Q�睡s9�sͭ��rv�ݺ�C&|W��.�p}.踶�g�����ey�.�S[��q�^�����1�5GV�Z��^�_u�M_)��<Ö���\\S�ِѝ�^ry�#|�Ռn/
E�ݧᏀ˭��*X,�:�ن���r���s�}-��u�	�B2�92j�d�Ѯ��]ڼ426�o�z�7�ʀ���K=�n0?VвC�<�hB���%�����*��r:n�)�;��Wa~u��v�JW~���X�}ܱ��}Y}�v섽.ޖ�>H�H巪C�U�r����M��b�g]��T��<˜���ǳ�mO<^}�;
�>���;�q�H6){�e)˳��by  ����{���'��r�(��Ƴ�7��;��Q�]y�GF��N��s��K���0{p]=<��S�Ţ7x�X�z��h�WM��i�iߵ={����#Gj}����cCN4T0G��q�3.T����;9� J4���F΁�
��S֔%��i�ly	NB	|vqv��GK��O��m��Ui���3�U��E9E�=���QN��l��P��Rw��S�vd-<F9�ӊ_`��bq�WfB���/c����nvʖT�\$���L;n!ňl��� _�K`eQ�Y��Vk�nݓ����[5���>a�mO��dC=�*`w?e@����X��+\�q�s׷հ�����L�&��:��vX�q���r|٪����1b%D' ҽ�h��<�w�i[zsjx�C�]�8�4\q�6*��{���w���6J��(�y�3��i'Q�d�!g3b��p;z���-�1�r�d5R��i?a�`P�f��1�5خ�c��6~���Ө*f7R��u�G�}�)�K���<~�_`й)�Z-H�u��:R��+�v]z���x�;\��+��pr�u�*�8����[�Ә�3z	4���k���y�I��;ri�=���|�۴F�{4���b���u�mU��A��!Ъu+_�.߫�YO�!K^6FӾ�{�Q�6~
��t>��dj ��Q�@�}g�2���t�a�41�z��蜎o|-)��bV<Ķ����&nA�n�����7�%�W'��艖�qvYU�v� ���h�L��&�Q���(�cb��Q����q\q=ĉl����sђ�f�呷*SgNsD�f]�Ff��?23gx��G �秅z눜�@��2�ℳr��߬���}��w����6/��<�*[�r�Y���5����S��So<���������0��ھU5�i��H��#p�"�:d����I���lR���o;���;x�4AǾ8��5�^�򟳮庳`鎧D�k���ڎ�.�*.'��h�=�n;����0�yZ�	z����!̵B0��=y��WvI��L��!fP�zh�!�B�i�Q��[M@c28��da�ٞ���0�F(�=���,�z�C��ޞ�U�<2��;LB�0��mk��^)ǩ@wS�4JN�8�t�'�9^�0K�t�;p課�''s����ԋZ�w�ԣ�*���Θ��t��UL��	\��J�D�^�Դ��F�eQ��Wj\i��������F��j��$�x^��gu�sO�<�yw
�:ju�ΙK�	����8�g(�;Ǔ��̖�l��~뾙�k���J��K�杒ז��e-��Z��G�H��C,F&LnR�����Q	9]��0Gi��#���e�Ц���ݎ�2O���i�'M�䳎LB��u���_3��0�*!9ЋGZݟB�h�"㫦�)��c�Fd`��z�w9��k�W���ݯх=��R����L1�G:!�Gm�a�ed���3+;�JF��{�D>+�OJ:v>�2�8�q�����,��v,r]ڶ��p���"�L��~��]��&r��c�G8�c�~��y���׈�p7�~��I�!2����u��v՘jdܥ�o8�N��/�z�Y/�e�6f��s�_8�s��F�E5�,\���K��g/m��^(��J+y�2ʸ���e���� �t�h2��ǝX7��/,,̼u��w\О�r�w�������t�q��ބY�N/�����(�	��ѕ���:�F���Z��a��Fg>t�S�_]=�A��7C�7�Ф
�u���tr5��8��Ȧgg�cr�c(+�/��T���ţ���y1I�+5�ۙA��F��ޙ�u3��ߝ�H�4�6�ߵ#�j���ޝ��;�>3)T�I�.�r;|�e��ӽI�ɋ^��}�u4lE]���r��7d��5+:�n�a5EZw�m�	=8b�4�R���7cQ�i�ss�S�6~�����{������Ί3�_Ko�؅����0�m�fZ��LBƅ�#{r��ay�C����G���!�9�"5l �
:�o\!�s�ƍ�gtw��;���a�8m��E]�]d��h��wME֙�t7�6;���H���w.uQ'�bĶv�G{��%;�{s�{8���ׄcף���J�����<�����ӕ�yFɏQ\so?a�-�68j#3K�Rj��Ǚ�9Y�'������:�+�فr�
h	��<Z�#�O#�Tn�ȍ�� u/�1ʲFƝl�Շ�s�<���m�AB���3o�ʎ�>ȅF�Q�柑�����D����-(Y=auDf)�î��6�vZ�G<��Ǒ�v}+�sķGT�嗼�\�OVce�݈烫���9�{~FO=��ڧ�]u,��*����p7��f]]ֹ�e�͗ȵ���]j0sG3w+��L��7t��z��p���`�����%WK�[S��2t������|����1���3�����Q�=�'\[�6�e�: 갵�t_͘��0)���.���!�S�Z��wq�k�Q��է1K�u4����m҉#����Ne:�Ǻ�ꚬ��I0i��/���VM��.�>Ӱ�Q�d>�o�����/l�R���Q�iu;ޝ}�Ѩ�䝌���߽��~p��w��n�rpuz��z�.��P�m��v!��R5Ş70�\�VF�Se�h�w������t\O���8��g��=Moc�3��۠*��1��լ��i���m�t��{���Π_ 󓆹����^+�of$T���m�-e�{��_ 츝 OS�����sȫ9��%�m�<���Q��G]^�Pñ]\����9�r"9�2��2������6(�<�}O�V�Es>���8n��M;CC�XC�P���e\�2���_\d�I5�C�b+�����ڍE���-��b�
���eԆ�n��ާ#�����ؠw�4ej�Z��;KS�j|%}����4�M��I��7�ǘ}W��y��e���d�v� FYEB	�6l�T*"|���	jwZ{�k)�b��4�n��h����9��	�v�P�[S�Ґ5;��'x�jj'Os)疀�9����d�3���q?i��.<�z���	�kYp��:ï=0,g��c�1�/�ݚN�]�;�=�Y|.]����	��q�%����؅���ʷ���zg�.�<��1�y�K+��9��Y���h�O:�gk95�ͮ;� V,{��i���nG�/YH��S$��E.s��Ly�ǡ�<`�^�lz;Y;����3�u:��O�l�f%����|��i�	n���M��MK�Z�|��e,�f6ff�m�o�R����Mq��5C.3|챞㑟1�ruI\É�X�۱�\t�SV�'Eoc�ݐQBm����"㫦�W��׻7�U�v��=�i�`��6ՑG����w7���^]r��<�ý3�w!�ǙS�`KR~Õ�P����.��qM����w�Ԣ5�3q����Kq��G9|���e��0+���=^���a�=����4���}�]�vwtM�Ћq��ܜo<�<�F僘��������uɨ�,�l�9�p�*���0i��+��qÄl�p�mw(�W祗D�<l���8:��g����C�ݧ�Ȳ����ܶ��E���q�! c���qϹ(?�.o�b��3�����մ��]�*醴�y*�/�4W[�^�uVx��[�`*�)�'��k���8ջ���4\q;��o�?2�9g�=�~t�p�ӽ��qi尸�R��g'�+��gb��]Qs236����=�=#�}\3��{�^�����I�uٯ���^��:�X}�2b�􇑔�F<�3�$S�/+%�wn��w�T{�ӏ`aҝx�g4r�r�S�y������#S=w�ٮ���])����Q{MwS��k2��}������t����|�씍7EŃ��[R�E�ӽ�-�w�)J��/�pK;CEsr�9�7{T衺x>B�\��{-���'Kmz�D#,����6*�F=n���]Zf/����߂�ȑ��'���N_�T!���+���S.�(tʵ��6c�v�2%����9+p�{��`�}Fi߂�M9Q�W���3-�p�~��)�\>��3�-�n1\�0�3Q�k/���w�3�	�\�B�a>����Y-y�vYϘy�����B�p$ǔi���5B���FldW`�浪�E���t@�l�4*�#�������쵲2{Mc����	ە�g�ݱ�L��֕^S;G�	�
�g�6X�W�$\y��lP�Q�m�9֡D�(�V4�6����ءl�	&ޝ��?y���Kuܳ§��]K�g�K��B0;�dl�U�k�޿ODe��e�fԕw�:J4�e��?@~|G�Z:���W�C:h�2����SζGqǮ[uF�0���Z�]9�����B�3lCx�4��ޖ׈Ɠ�������ڬ�����
��'"��T
�|����\�`�mU.�3�M7'ud}SGj��Ð�f�*��zN��}ڕ����r��w&܀vs��!c\G7<���)��^���KM�$�;o����C[7���4z����iR�w���Ǫ-��P�Wm̮l�*-j��C����;`u�V�H�E*�Tf�n�=vHohp�V��]X��n�ވ+�;�!�j��M=��]��c�d���r�����u*�ZjT������*Z?J	�x��^n�W��R�ҧ�w.���ç�3�u�<��F�󥜙�9h����Q���hz���"��D�fmm��Zb�I���f����g������aޠ��pi�(7ۧ(�B'�̑���@ �V}GdX�|ja��PTU!�;8V��9&�����ބ�vk\�ˢ�=�����ӫ=<)�,Ab���tVOg���-���;-fR뮠1f�fxj%D�+N=�9˞��1<�`�3��ƹ��b�!]DV��*%$���x���d-�ݝ������[:p��2��ŎK�M^4.�#�L�[w�\�ِ���n��Wڸ5#.�� �B(OGR��퇛�J��IMy����V�WՋ���pU���;X�C�[�����7!A�؃pZD��vӗe�zdA)��XI����o�Vh�s�W���|+ �7�'@��ni��`�<;_Q������н8��1�So{�g=�ӥi9wc�
��,���D�cnƼ�˪���_m-�建�vwQʽt���I�}�
�hvK)Usq��8gۚd�|�g]�:�h��0n��uo{8�a�3����y�	x����䭗�%7e�%L�Eͻ}өL���X����y�#�gx�4'��ƍ:��x���}.W�����qb���|���a�VA~�7j6��]o�3ݝ�9�%�S&u��n�R$ڷwh"���_>͂�L�И+���L��]*��Q)̧6�X�� Su�A�����G�MϢMN�C���`�l�{�1��Z�b����"�Pf�S�:�a5e�_q�·.����ej���Z.��f�Zf*DB�r�n�;�tbSA�S���t�>�������kW,@���Ck���;���i��wj�k8�b�ӹ���WT\0eCE��d��^�Sss_�����-j�x���"i7u(�#��
�����=�oF�F9Z8�M+����0Q����:V��c �H��l���xl�WXU'�8*X��ȔN�:��޷ίwh�`����q�Zx�����Y���s���F�$�u���=aq�{:�b+�]�CY�2�3��oM8Q׏;u22 �7���7C�Zq7���|��p����ۭI*��g�EǃVP�x�푌yh���T	��ٝH*�z\����}**��åW�Q��lؽ�<��v4�W�ag;sG������E�|)������������I�i4�$������<��mBtZC�v-!��B�5v:��4h�HR��TiB"��֩��::M	H�H%)��)��A��(.�Bh��+I���HI�=%��S݊(�(�*J�)*�(�`4���i
����t�JP5A�D44�IMRWJ�j��
 ���(M���:�:(6�@h(��U�ON Jj�
B�I�)��M��BtiN������Mk@ga4����q���T�])�WNئ��CE#�=�N��4����.�t�,F�E5M:SNf�(
����O�Cud�x�[�V��3b���z��*
�|�����T�!�.�	/uiB����Y�2�R�I�)�ώ�aGVek�`�n��p��r�-[ߢ.��Ӝk*�x�e�=�0���C�p/��wL�u�!�%��sV�- ks0���}�H��8��f"��=E4��e.��P�ե����b�e��$�`��za�Q�ͽaҨ�m�P_�7@}=<.��"��[Ћ3�N/�Sk=k>�T#����w�r���aM�����g]=�*�g���V�*=���]�I��1(Jhw�Wݑ�8�P�nv4��钎©���egE�+�^y��q�9o�V�J�U��f~��+���ٺ�M#�Ԝ�l�\�D�m[<�b��ֻg��� �6z�L뛞mj���cк�h��N4�3��W�M�/��;��5��)�#y�˕(p��ٱlzN?l���=8�a殓�4z�sr�#e< =F���J���=jy�	s�K�S�v���l��k��Ę܋������T
m��G-���� jֈqp�
p	jz���#���;�-&�����`�w�W1{q�:$����]��n:
���:�+~���
�
�w^Cp��h�5a�0MۗgӹZ	�Ƌ����9�Aqzr�̫ԍN�:̝�U�*���~�pI�?a��n��y��Rޮ3)�q��{�-�LZ5et}[��5����Rq=mg;����ftm��52k��/!�-�?:!���ђx�}������T�Kx��T-�������_�=�]�!זV�t7T�ha>]�M˴r4Ŏ�00t[uqצ��P�f�䪼3:�*{u��áя�P�{~F[Ǟ���<���q)ц���=oF�5�f\�Ft���4pv��먣^'Q�b�M��of�G��� �e�@��\���͵M^P���}��s?@GeCč��t5Vӹ�������vQ�6�k�Q��ʊ!U�"v��Ơ�H���Ǆ�����f��U��'X�0�����6�����m�ӽ��&�X�UdB	����l:.>�?#{���oT{���g9��Ц6z���"���k��:�n��x�Cn�����[z�Nu�z���n�7�	b�Hެ��e��v�#v���B߼���q3�8	f܄���B��.��>�vg0���������� �E��?�����{����l��v6G . ���2~§:([�k�1�U҅ѝwM\z���-�(ͻУ��\�W-�N��-�)�����t��/m
8Z/��9�+W�=X��R��{F�Ua���9'u��Rj;j6D�\�;8cj��V��[ʝi	�\Yw��Ij�SK�<���x�L!�P�*�m�AL�Y�w��l
�r��R�z>mU;� �8E��5K��ܐũS�35�E��iٝ�˥c��
=t�$Рq{�hj��I���ڞ��J[3��[�	��"Zk��e�:���t�y��\���v����Sv@��(�A=F́�T*"��C)�i��'�tde�ą���O3d`��ӸW����e���[+�����o�@\�� ��{7��o���W�{ �2~Ӳ�qA#L��CQ�r�A==L�x��n�,�L�0��n��Cd������YYY�}�F��d�/���Tf%�����ʛ�H��*`O����峪�yЂb���_k��p�~N�gc�t��U2,�Z����c�����<,�O.8,�@�{�j�r�si�������峮D�xG������.:�lUx�{�d�1}��m�M���2�6��6�^qٛy[�%9�tt��r�S�Aϰ�>��9lѐFU(�0%sضLٮZ�:�m�i�ݎg��ȷi���[O0��z�%S�!�8d��W]9X:��c���c��/�Me㭜~���E�E��Z㡡s���.;���`9I.��n���[4Ș��F�nT���eG��ѼSq1�����+>}'=	�҃U=6DW:ys����,��F����N�g]3ӼXI�Ŷh��@�v�b{_n�>���bK�n&<���zJ��U�=|T�Y����LPp��?A�ںm�^�V���C�'�gM�"��=���X�{��3%�ܢ-ds����V����&�]*��[J��ckxV<�VM�C*�z9eqǖ�@��G	�z�'r~7���)�FwA�-l`���Y7��v]@�%�M'r2�td8��\�7S[�[�@W>6��8���4>�a�m���sffk���c�p=wd�fT���/A'z)�˪w�v�N->:�K_�ͺe�Sp7j&�o����{�w�R|e�r�^nܓ�Y[�)n��j:@�jP����{E�:�����b50+kS�us�̟dh����ϡG.zgW��5�#Kng�u��O>����mM�2�Fn�2g]��g%e����}N�oVD��#���P�K�N��aKe.�	��ջ ��]&� �O���mH�O�f��Zk%�,O�u�Tp[m���g���5�͝Ҥ��(��\���tC��]�\w<�=�k��YL%��s�K_k*N�n�k+#���Z��r�����>Oo�:G��M�iӕ���$e�����r�
hU3H�yj~�yj̆O��ۖ�cf1�Y�R�4�ːp�X~L֊ғ�GE�٨W���`����tr����Cvӈ�x��u5�$1 M����s���W91<�<�m�S�'V#�e��P��[CWp�{ي��e��4�\O���mR_���6��ޒ��e�ӝ�K]���N��ݼϢȌa:e,���s"TBs�����gв�.H��WM�S�g�ph�}J�m\#Fn���~v�ǽO�)n��v�*�r3>��3�σ��.H�������[�ӭ59�3�H�mTT�A�v��(M��<#�od���<�]0��0�}����L%�懆�N�M��3k'��9�D�,�^�ݕg�[!����x7���k�㦜�7F���Qo�9���|��\a�g/��"�Y\�9���ۆ\v!Яk��
� ~'��8*��-�bM�mgν=�!O�lÇ�d�qXi�28a���]��8�Ŕ�.z���;>i)���7��Oe�/1�=n�-uD�Ψ.r�8:+��S�Y�f��fӋ������{�=}�;@늖�{�v�#�����}}t�Z|ܬFa�t9�{L�H�f���(�lh����5�/t���u8��ta���9W���U<�
;
\�+�ٲt�2�!a���'C���S��O��]��$�������{�-\�oc��g<���Y�GY���CEga|:p�����B4��_�<�]��E��U�����z��u\&��� %~���,�	Ǌ�;�#�s/V!Y�:1\L0�Or�I��jV�[�3W�'n�\)��*��[�2��ʷ��_U�ٷFj��:1k���Ѩuv�R-z�zƓG��'��g��W��gKX�j��Z��3N�7�{�RيhKq�v�d��XmZ��	�#�"�6�^�j�J׽*�y�ƀ�����S	j��e��K���.�O�N�5��q���v��5,��5Sv�k�è�<�xi�(�3,���P�f��9
h
3���S�wr���uGb�;�9�.�����g���ҥ�0�NxML4-!�t��l�Th=N���]S��ٷ�����?q٬�Oa����u��܎�-�����,��۳�Y:��#*��o��̾{�;�jhQ��ov���s
�����`:��[���9��_8�pDa���NO>5R�qW	O� ZOpŭ�gr���VeF8?�x�,S�O����Ui�b���_\I��8��{݂?@��^Fqˌ�3�����g��1*��,���	����
m��Y����p��?9x��$����7NN�X_-Ւ�ʿ�"��7��-����(��c�H�^/G4sk��h�g:a��8u27 w�����9M�����͎�k{a�<Қ"� �$���,҉G�ueK��}���[�x;�*]m������C��T~��cƃ!�dK����$�՘z�0�ӑ�k��۝3���C����"�m����C6����}hJ�9`��?�e����]`�N�C�]�N4C�����/w{���~�E���+\(`����˞��z�K6way�4���d�^�B��@έ�ڧ�܋��ڨ钇3u�Y�<-�͑�>�"6uG,ې����P�+��r�1vjqQm��W[����=\S�8�~d��?y�k����4�e��~ U�+S��d�eKgE�H�m�� �u�YX� �]pQ��S�W-N��,�SF}��.[: }O���gt�Rc���k��o9�����ж���u�U:��L�
�KD�I�=OѨ�	?����c�r��Y��i��N�3�[}��odʊ��l��P��3�����O��Vl�F�y��@v��üz���e8\ikI�A�� ,�4l��2�%�t�s0c���)��u>"�R;��9Z�7؟��vA�:[�1�*YW��I��T�|.�N��z�����S\�fsGL�RIZ^O��0�-�Ѻk���=rE�U;0.�f��q�ַ/'3�F�m����5������l���LM-{��e�L�^?x_�?̉�fuM��Ǒ���ŃZ%�v���.
C6)�Ȗ5�A��=b�l�m��4O[��� ο
�ugoJ��;��Yp���t��e�$�+g^՞�L�9��y�+����m.�2�X���6�=��ڢ��P�:�����S�.�U���e�sœ�d��V_Iܑ�?��ߑ��*!9ڠ�BZݟQʋ�.:�lUx�{�lJ�|!���۬�*2�,:f�!����v���jp6��.!�Dt.��}�1�r� ��U)�0&��H�M���.�B��rD����tt����o����y���6���5 <{�q Cy���ϝ�,+���<��0�:v�ⷲ�0��e�c�L��1�,~��Jͻ������:x���`t�#ܜv�t%v��U]ʨ|���g_�W1QvYS]��-��ۡ��f8O�ܢ!\s�����{�v��p�w�Ifؼ�fG8~�P�ʌ�Vi���[���,�\m�! nzxS\D6nJƧX ��4�v{&�0��u���ݷ����m���&ۮr���"�����
aq� v榽�nl�`�����d���bѵ/a�ݗ'�+�3t�{�M��N�o��֜Zq�WZn���;宼�Ӽِ��\n�=i���n�s�Y�\q=��ށَ�6��.zf3���W1�5ӕ��d���y��"�����"5l �У�=:���e�/����B2��O3l�g�T­X���"���F�w���u���V��$��M��P�I�<�=����ڨ��x}y�J/�J��Y-f���xr�w���IK{�{:P�bX���jᛮ��<�'�ox��]��@�T�9Z�$�U�*��]W�!�7�X��ӓ&)5np��2��J����)�i�;w���6l]�w�3N�oc�H�<�f��N-t;��8N�Y�d�8��h�\3n��m�=s��w{<1?l(�3��l:{ 	���(n͒���-��nSvJ72���y~��q}y5jvuh�uOX!'�w�=F��S,.��S�Z�Օ��Ѻw'�BL\F�lg!�����c�\��y��j���,R9,��e�Ъf���OݯE�Sa��/&9�L�=H���W��Y͜������nx��q*!9�\�����>���rE�utءmK���t�ɩsWV��Pz4�gfF&�]���>���n��xe]`�:�i�膍��ܳp�1G�1{����7-�2�ΰ�£��O��oǜo<�?�̺透J�2��7�I�u������֮�N�5Qnb�Y蜄,k��o9���ޖmx��b5=�N��Rm���׻�ln�31=� �ܔ�/�	:���;�T2WQ�a��%�q���4��r֥Jl�Y��Kҳ9�x�̺"ơO��f<r��a�����QAO��1嬮%�Y@[y�m�G�s������(WJȎ)6��뮏�vAOt|�s»h�c�Yr�d��+������}b]�H��,��Q���d��C�nb�H�a8��S�������5�a�A2֤�m��i�#��\��3P�@�-kl[�ʛ�wq��Y��q4v�����G����/�˛���>�����v�:�����Z��Ɂ˼�*oB�� �ll�����a;����:����������4�hި�&ᄺ���V���9��2P��3|�Z��x�m�c��%��w�����B°
��k���5�1Ff�Yzl���&z:XY�u��N��qV�C�.�F-t!G#���(h�U!��}�Hp̺��7��P�]5�C�Gi�Z�V�Z-�E�J<7����Q#x�;} <)㊦�)u��y�,s�)�L���r"�ۦ�{=�T�i�S�(�:ӕ��r��OB��^���<�r��Zz�>ʞ��NSvA
L�c�8O�*�����z<�Q��<�v�&t�wiB;��gO�t�,��]�l�����;�,R4m�W�0-E=����i�ڽ�M����E��A��;���
[";N��8�#���.�2�VY�w�^z�'�Ma��5g�t������m_b��lƝi������BӬS�7�>������_�(*"��D_��*"�AQ�

���PTE򠨊����+��DW�j
����_�(*"�T\����_�PTE�+��
����_𠨊����+�AQ���
�2��o��`�*�������>�����	�������*-��T�B�Z+5�W7f��"�YEH�9a��a�+U�j�f��v��ۛe��
���٫�v�vl�w`+]����裻 K��ӻ���55�nó�,ڪֶ��Jp�elmkkV�[
�t�jհ�գB��e'e��թ�l�wqJf�iFV�f�n.�f��m	M
�     jy�EI       S�0��J       �bdɣ	�bi�L#0O��T@  h    i��&�&	��0`��$�@���a	�F���bh�)��{�=���Ƿ�D I¡�� 	 z��ID&!!!	=!$$�r�@HHן�?����O�Q���ghF0&@�R	�jB�<0�A�R`@������Ɉ�?����>��$$Q9�*�R���N4ϱ>?-�*QB/üז>a�	�i(��w�����i���u(�:B2�аU�j%��׊�ʕ�	�>�L�ːMu��vp֗�\H
���V�U4�ԊX�O7Z���r ٫��֝���ìw�0����7v�C+ �zHe����]�Y3#3pe�Q*L�O+3�!�;t���� $IJ;�p�c�n�Ʊ�A����nG�%���Y`�{��ݣ-�%4=�B��D��g�)]�k	`���ݻ9w�L[j���w0�]�e A�A.^��K�X��� ucF�i�4?�ןX�L[B����Kpy����_
6�+akm�bk{O&�pL4�ʚƆ�r���tl�U�)�-�)�b���k+Vc�A�wZB�.m6>��&�h��{jZ�*%�6^�#0cR5f�҄�@�TP�gZ8f����9�%n�m:r�GkpY3eM/1)si��ܑ�B���wXԌ��f$��Z1bK.�1M�KjV^؆!+"%�5��v�0�Sy���<�ѭa�t����f엲�L���w��ki����bb�؋uxZ�)�]���+ z��7"sb���N���j�yoC9�E·q��Е�EI��sR�,h,ZFa&�
��;nP�&Z]���[kkAM5)����k)� ���{��� *�N��,i�v�H���7�˱�Y�ì���� ��n�?,E�O$�Qڭ)A6÷h�l�f�f�!����/M�AY8TF�J���[B����޻N�b�`u����_$�k:���ʵNO�L,ب�H�/Xy�c�E��Û�B�	36�K{�I��:8��d��Z�������6��� ��)PV�v��ɥ�ħ��3[H�ۍ��P��s\15���Q�m��åkȭR_f�Y�VkkS��^+�Q�"�혀��p�Zq�Q�y�0U,�4$2����z�B�5��# [V�*4NǠ��T&���ӆ���1���J9�����RcYt�̬݀ �ܧa"SX#ؓ�wq��,�j��Z$��1����$>/�^��lq-�8Rw��6��݌�t����2�7,O�� ��-��T(�N]n�����v��+����U<?3����M	�Z��H��%e�.z��l���W�7P۳�UY�����t\hw'm�9(��v�:�	F�9n�yk����ڧ��$w/�sG�M���*tc���$�"$�/�x�J]�k��w����� ���c�ck巻u�θ����2;*R�
m	���%�'��ju�g$�ܧ�m�/&ˌd�G�U�EJ�V�Sj��As3��[�{c�N�_���;L �����׭�w�,��1-�\52R�X�n<q%jd�SF�q�֥X�^fN=`r�����=g�E�.����wi�G�2���-���}�@wÑ٘%Y�j��}�Y�ؤ.=F ��:&�nv��l�ϒV\ňT]w[�ZtA�k盢�3���@u��cn��y����ə���&�^494���}a�K�BXס%d�dhǅ]��rr˽CgIX8i��.�j�9���s�P�4YYf#oD1�/-�r���hl��;36��bX�`������u���ʖc��:�d�n��w)�P�Z)2��F�L;JSwl��ew=u���Rv"7.����P̮����Z{roiN�^�ܮV��s�wu��j��-�B������_A�*J���V�fl���MaW"�d��"��� �"�J�
��ϯ�;�μ+M\��i;f����)�b �D3U�e�v\M�i'�4\�w�=�`=f��1+c�)�V�r�e#���IX��H0=��v���ٻ�Y���#x$�3/���>ǜ����b�L�k<3�d8�h�%�I<�s�Q=�"^��z,���y�񙗕ҡ
ƾ�(�F�S<"E.�bwj��#h|Hs�!�ȥ�Ԑ��mm8s���J�t0�L���n)Sx�͉Um�Ɋ'-F�d���V�7����Էu���]S�ʽpޓ��ix�؇Q&���X��bcPm�ܻ}V;��o$Ȭu����&W��18���lo53d@�۷�Y�٭':�3���e��ij�b"U��+�7ev���#E�o#��q�e�K���`�9ku�P�SRF��n�rc*�侖ld���;uA�!5�\�q�]�7�h��X���Qp��������B� w��:��n(��ԙ��:�gUg9����ֵ����ϟ���~^=Y1�I! y��7́ <������	$$q������}ޯZzc|����9�d�k�ѾӁlaZM�Ě�1��J�8M�a>O�*ai�2nAn�@��h�R����g��b:�f������K���r���8�m��a^|���[�4)���X�#
n;��[���1�Fl�[9��(x)��6�� b;��Xb1B���'X���ܔ�t��Ŷ-,"�^��-Y�K]��G(SyX�}���{�r��u�8�a�[$�+�T�n�
=ْ�Y� ����'�(<˄,kZ`+_NՅ&lqh�ݽ���K�ʺ�رH�u��P��]�c�mݥev�ܘ�w	g�h��y����W\���@�`m`Sʽ�L";��U��$tY}i��cޫP�,�����\Lǜ�1dA)�~(�BYN�܈�?%�i>��/����W(��7�!O�^�˛�P�K�X�^��i33�@��J��b�V��_4�ۡF�䓲TR�1���';�lbf�k��`��T\�(�w��/fv��л�Ȩ�<$�	�w8�F�	Ԯ�f�q	4��̒�j/��*�gx��qN{�M�Sk�[�9��=ꕝ[Eɝm�����=��]��|�,��Lk�ޟ+�����⯜z�F���x�^��*��i�"�.���N����e��y�t`9)��l�C+������u��Cv�� ���* 9�<�;w�4�ƓC��ӱ��3+��k����X1l���rD��m`�G_6��Uu*��I�Ei������&�R���C���2����ӂջ������+�6��,A��0eY	�|����ةZ�@����)4/�ݚof�]شh��^�l���qᆕh[��Z���R��)QN���e_�Ы*�ȃS_[U}��z�<�Z���am�ٴ�3)��xc��:�b����k�qkېn�
�G�V�>Dt��8ӫ�Ei&::����F�ޥ���嫏i'�JaR�� �h�dZ�vc�Δ�-څA+��U�`Qv�M�V�v]fc���aR��5^�`��������G@�������i�]Wu:*��i���A^�r�h�r��i�z�'�	!  ���<�r���^)	�g~3�x�ўju��y��;P�څ�Z��t��;��7(�{F�r����]|gIH]-kz���(��=&��Vq��u���(Gʸ���(��������x5[\��Q'^�'�+�)۬YϺ�u]r�پk���c(dVT��nRJAd�*U�.�qm��i��)B4�H�E)���XS@E��2|w�x9�>:�t��ɜ���g�� �"���J���&Kϑ$I�=����b�:���(�8�0OW����.��_@CzK�� r���_������f5aS]�'˽x��&am�|´�GC9Zc�`���7�.q����LC����3��>T$�b1g�7u������n{]" 準��H����K�|�l�fs:�go����,�[�w�EQ]�䍟��n՗��ð׶e G��z*�-U�빑Vb;C����U���]1��["�9Қ�w=sDpp?A�s���(Di6�
��\#��VǞSz<8`��)�Q��ʬߤL�\�j�3,�{����U��38�s�V�=�z�վ���v���%��@U�K��hio;�;�b�9�Cҥ��T����=u3�j��͞;w�����EFZ�3���g���w�&��<BRTtlי�گrS�]�i����[�;���:�s{�>.!�<�"��ʲ`�[׍�`��­�ԩ������!Sx�y�L����^b<V�b��ˬ&���x�s�V����;��2��kq������h�u�#b:�C8L�Y<����܃Wg��%Hǧ[NBa:;kv�r�$�����tuV��L��ļ��K"�[���ܚ�{,4bwYt� |��Uz(ν�ի�^�hs�EP�-�N5 ��X���}���1���~j��V�_�р�y��7~�4=�/����2��wn6���!� 	>�S��*�&qu���r�"���?q�x��o��:��kOX~f���(�z�7<���|5�[�e����L�6�x�f�c��4�b�9�n��<x�db;SVb����q�Α��G+����OP�z��5�k5��]�`k��in:�Q[Q������������9�T^�L���+{�f7��k��t�"n��m�1���5��h��Ӽ��,�VZ���w�q߯�͛ӹ嘬>�
��[�udR��d�Ѯ-.%X�m�oDbL[a�������R����S��X�㕂˘KY���M�t1H��a�	�"YNS���)*!  ϖa�D�H�5�t�qa�˻N��R*I�u/!R�u-�.Z2�L�.��f O2�f���xӲ�^ӟU���a9T,��,H*�L�,V(ILY)�oc=U���f(FFW�nJb]d�B�U�zs��S��9����q��0y5��~lt׍-$�ʘ���*k�PӞ��5�#<��p]Y0��M�"ӌuAV�]�`��Dӫ�xVz1O�X�>���ur~wX_5@�==�1�;�Jg!�I;�a��+w~v��PX<��筛�=�bUL)�Em#��{��N��r[�Ό��q_�yz�v����4��W�2C(0�hRBm �H1�	�gW�L$2��$-wD���,�ZI}��BCli N�!���2�a$��5���C�D�����v��m��z���L2� E!<0!L������o�C��N!$�I: ��R�Cy��ˢB��VjCHN! ����:��Y �)��M$�Y�!�$8� �Q�ϙ��ܪ��釵�۞��|��n��_d"�)$����;�Hm	9�VĐ�2ABa&����!��U ��C|� a����I�HM�Ӝ䐬ԁz�]���F��;Ӻ0��ڣ_�TZG�쩌�k}�|OR�1n�$5n�9'����Ct-�����t?�w��K��'qO�C����VV{Z��[J]X�a5�����ෑP��.����r����-v˜�-eX4��5�׆:��S��)N���W��?�==��s��ss�×��d=\F�"X!T��y�Z�}]j9�O���9�T�.�^��x��,���W���WVB�y�krDˠG��)[�U8�SݝG:���v��ր~��&�c��d��f�׽�ς��<����2�>dy�������i���#��i��u@
� �^��+��ʷ���F5�u�='D�v���멩VoG6�yώ�	X	Oی�t�Q,^>T�nS���ܫd���+��eY�w(��&	j<%F���/4p�'զ��л����鲖\I�dCY#����#�qg8���&�ی͞1w�ﱜ��e����tǞ��=�]��&�n).�y^٫�];���S$���O�n>�ߏ쮴Bm�ʆ�[;��.ݛ������[�^�Y��DVx>�� �~���Y�zg��-`�ٷZ���<bJ�g�}S�����{��y�k���i�D*�0��w§��|�n�Z].r֡��g��|��)���*u�	m��%���� ^�gu�Y�+�`�k6��I�;�j�\(����l�}*��[mq�����߲� <?m�j���ڼU���n�n����Qw���U��i:"�5��0LX#��)�.�0��L&�T"�d�R���j���b��(�24�(;����vQ��3m�kC
�WJ���UR�Sb�b��S)"�CHUQL$R)"�>�D 	���韕O�߸��kۭ�)|��?<f��w��e�_:��W饬N�֔=�]�P�/VL�J>�}��}Qd�g,V���|ѫ�;��+m}.��*�ɍ���+!�m��ݔ`�)�$�VLk��Q�'��\[4Fx�{�9½[�'�c^D�3�ُǥ���<�'O~�u{��Ӫ#|#ՎcvW[=!hN5�5����Q�ݤ�[��]#�a�c�����
S-):e$�wzJL��t��e8f���XN�L��Jx�b��q��oi�)0�'i�w��j[{e%�\�[fx�X	�N�wF�)-�vQ-�{�s�e�L&j��=Pi!�Q������r�֥+�LMJ٘����7���m���
��5�J �T�4G��I�)��ktctR�n���J~t?{��.���Y���"���`�+U4�p�JB����2�:m2�wFuA�iˤ�;�-1�&f&�W�V
C���0���ц��ZC��k����K�qZ!V�
<|� AS���3�WM��{'uq�"蹮>���ã��L3�wgL/:��3(a1�YWE榙����ʛI�)S8�	�ޓU�k%!He-6�a�&�r�B�Rm-��skί7�1�a
gL�ιW+U7�<z�M����ᔔ��f�&�a�m�p�{p�	�l1���>"��j�APW
�j������ ]����3��S�%�trN�_UQ�T�E�JN�Sl����:vop�a�<%�eb�&^�t�n�oN��Jf��1w0�śL���V���I�����VR��4o�_l��m&�Ax5e�;�%ޞ�Z�Rö�w݇}r��F�m��ғ�f�x�t�wu�)����}r��E�x0�x��E���ǆ7Շ��0�������5}�ʟ5� c7T��tL;�O5D�����|6�1en��>7~1��Kfɨ)���,;�j�?�Z��|�1X˽Ѷ(a0��&7}�;���	�Q0�i�)�Jm�-��V��|�Z�	��C]f�{��GU0�!o��M޽� �,�JDF���
p�m^܋ � m�.��G6g2k�<�<&/[a�Hm��KL�L6ڳ�	�UQ��8�%n�0��6���cu4���h�4�4�M'#��z�޷��t�
��S�(ۄﾞ��)���\�Ѻ�L�U6��hb뷭u�ٌ��zN'*�hR��{ѷ���Vkӄ�x�T4�-�Hw�2�L�^��&��!j�O��UU#��W��u��&Ä�sx-��YChc5<3�[��3g�Y
���HyW>MbZe6�l��0ՔK�8v��J�xѳ]�!�UuƘ�ː�Q�G�F�u�4zV����<�R����gx�Z�-��hZJ����g{��ZN�GB&YM��E��Wsv��׀b�M(�B˃��P��D��@��gz����v�f�Zc�0ͺM=�Y���a7���aѺ�)0�L�x��Z���in��&P�1�1���I��5��fY�i�Ӈ�S����j.��R�E_UxB��m�L��cJ��#�٥���������
���[���w��e�6�Rv��y�������������w2!��ֺ�f6	Z;x
%&�c�=���͵�d��G��*q���`��*��.���3I���0�[SU�H|d�������y�+n�:$�{�T����RJYR�1�X[�;�,���g�aW��W��;b	�X�v�-eq6�a�d����xqL�VfZ�P���T�$���Y��ü���xS��7H'�[�E�N��!����ۮ*��HSM2A���Qe"�TT��
a)�* P��H-%" ��b�����%�BȜq����]c�o-�� �c}'nɼ�Z]P�����F3��/L��2�)�ќ^v�h�N8�˄�L!W��d�{c�9�(�i�2��(���8�8ЭU�H�m����B�{f.��N���+]�RZt%�ي����
2��))]r�+Y����;�,P������31��®�'1FG�AU�x�qGV�qO-��ˉ̓fD^?JC�795����'"���_U}Vo9n�I��Ǫ�zfsE%��Q�i�f�(�:�f��6������0�N�n�ĭPt�t�o4JC��
a��aުZ^h-��뼛v�ͦ�2�N&ay�w�x��R�}�sX���J�,�(P�@UP"��"qf����Q�U!ز�d �#Ȣ.*^�`ҋ���S�'{�T�U���=b���؞*�ݥ���D���M&ܲ���o7E0���He��aj���.��&9S���2гZ��5tC�m��#�6�dȚB��v�t�-���7��i2��u�`�В��n�%3�Gi���zφ�")B>c����s� �/eC
�'m(���V����z����G�%P�xt���6o������J�c�9[���4�5�������Nbv�0���xr}��&�wz徵�,1J�ܶ}s.�fׯ"�GX����G}/�t2?��U}�4/ߨOΩ�O����#i)/�v� j��+H��\�cf��;��V6�vn,�x2�,�J����Z��=y��՜���W��	HF�v�m��(�R��m�3�]m��w��U}_R����� m;�uG6*�Є�Y��@�M��j���K�f�"�H��}�*�M�"7��,hy�0�Sn�9;F+j�1�-���HIEk��ww�q�sͼ[W�����V+�_^4&�ao�/J�P�5m�b���ל�����������x���!����=Q�ۡ�|����調.=��A���9f��IeU��&���ᙋydO�x��Mw1ƯJv+M���m�}�P��(��#�SyظJ�غ�l���wf���n�)������fO̙H��dڗY���~p~�ݖf���X3��pn�	�/-���]�S��
���.�}���aO5��-enГ�U����4q[�VCocZ���� �~%z�EDP�5�^P�D�p�tv>���V��J7ѕh�Y�М�h��]�������g�	mcu��ٴQ����d4.f�As�E���G	V`��=ZM"_B>2�o�ԭ����#c�C�=�tA�&�iԈ��O'����[t��2��)ux�����ޗ�r��1o1B���S��˹޽���.�L��:��zQ�{�>w����{��g�;�
�	��ugck�n���z0RBɝ��K�!}��>΃�;mɫ��!��"yi��uv�dc��T^c����k}���;��i�nZ������� ���a �,*R�b���Ql��n�����Ʈ�*,E�Z�AUQm�U ����[Qb�R7P�b
T"1Ee!TҊ��QUZawV�ܪ���E���Ȩ���$B! IG�5.���̜m����wxs'�E1=�jr��>�����,~ǂ����!e�wL�J�u����hھx�	�,�|�Y��|�|�����*�,5$�|c+�CS��}IV��n~�ǓC|S��k�JF٫�Sʵ��^�V�״��T���w�G5mc�y��Qvw.3�T��U����9�Ɍ�x���{N�Wy��盕���(ϣ���X;)R��{J�\u�3H�Zɉ]�@b����]l�;l;��*�{��؊�Q��I�S�����z�3u��φʒ��Q���e�ֶv^*�@Q�S;0�X�\f�����l��g���v�&ǶL�?sEx��ࠫ7#x��]�a���Z�u^7Cw~x]uŘ?��M�*�'���fC�ט�/���&�,=�J�1�u]r�l��Ū�wM��ԣ�*���Vlq4�*�Q��n��3��o���s�}UT�x*1_��=?M�H{K�G��䆂F��5���]95����ةN�k��D�6��,l���sٵ���S=��uUK�P����(:.�	����9���_!C�Ֆ�÷��.	R�ÕG����Z.�m/yf�J<���o|�#a����+D�fout3�	�wTvq�y�-u
\�a�S��U\����e�g.ũ��|>�[��.Hk���"�i�')���g�XV���y�<��r��Q�alK�`�E���<����фM۞|�����:5'~������m�8���!^n	��f��Q���܉Ht:��5���P��B��WbS^�¢�7��j�H���S��R����+3T�����V��u���#����U��n�������{9�P�ݼ�y���6��ց��q��k��3Rg�q�*T�d��=�F;m��Y�w��fXU�M��8 ީ���0��ڦm{$ә�2�B�v{6�Πs�����8�i��C�V��%^j�m'�ۖ��Gt��Hu���7��zsw�R��*ӝ�S'�e��fNv���3�"�����KG���a���u�{]��*9�K�s��qŸ�M���X¬�3�y�G&1��W�ټ���4G���FR�Y�8i^�Y����
gWr�spc̒gnէQi�}1�>���?^u�rø�u���cx���\5M#4�U�EE��mj�b�(#IQ�T%!QTQ�
En�	iM[E��J)J1KhUJ�B�Jl�5*�K���K�e�l��F���j�E�uB��EFU��STK��J��K��)�j���B%"|��BH��ʳvw�?5�������6�N�C��Z:��O��?:W�m�� 6+d��7~n���_���"����K��	��|2�v쩖��7��)N�U{��m�y,-���Ĳ��#���O�1�OҵcK�f=4uW�˘ ��j�yV�d�ڀA�~M
x
��Y������؎&�3p�<ܮ�ȧ1��9��{�a�N�(d�)G���� ��%S�O?��B�{M=�tJ���dm�1/o@��(���Y;2�#zk�h{���)��{+8_:C)�pm�R�BFц3+�*,Ύ�]ث�յ� =�~#گ����4��ls����`�.z 4��WN����e}��dw(���t|���Y��3�|�)��T���Q����gV8���o9q	T��<$�w�:rf�8�]�^`i��_�P��l軇��G�(���Ex��U��tn�x�Jz)W��mܼB�����(�)�Y�yӎ��w�:������ 0H��|�L�Io�˭��m�e����̟,^נ�Z�BN�a��Am3!��w��C}�q�͔�1P�ʢ����ME��U.����wVN��l�O/&�_< �'���E���B�,S!�Į��[����&��ׯi��R��짇l���(ة�b�ڠC��l��+����.���j��������Xe�v�~.�h�(Bt'C�ދ���1{�T���v�S��<�V�h��9��'cV��uuX7�U�:k���g�9��Rn>	���K�'V�l9e]#�L>u�-&=e�Z2��뺎��xF�Sn�R�[>oonXb�ޜiݏ7���A����;P���K%�{�{����3S��]l����N�(孹㶳��)��R�C�g{v����*���#��� �ȃt�3t'=�/=�V�g(�%�_������V�w���&�2''Ky7�æ�EV�v}i��<�����]�l�M�\�p՝�bQ��7;�T]��r��4�%NgV�tP�`�H��v���`�8 K�������~Y�����U��n�Ia�Ř����P�Ԛ&�'���-9b�#/$��ĊH�"�V(��F�rP���AP�B٠�2A���v�F�&|�K2c�QS˺F���ۧg.bO�#$janPFFl�0�x���9�K"��c@�
P4.�i,E�����R����
e4�t˫�*-���%��D���jī.کH�Yv�T����K��Z�n"U�5mYH�֪��Z%ݩ���9���#�T����t��:��-n((�����OƇ����X�O_E����ٲ���䧏��]�hr�c��^�3��꽛�u���#��v���Y�wʯٔ4ݑ*�E6���\o�����fj����� �0����7f�F`���YZȞ���%��۳�^�"�˪�Y��&�vۡ��70��-���c��F�&�h��%���ϴ����i�@�F/o]��7� �0�]���F��h����z�o$��N��I�撰/e��]b�Ԭ�-ض�dQu�jj(<�/<5}�Vv������m�n�{v�^'�^�Ԉ�֛VK�6I�l.�*�v��ok)�)����9�a�ipm>��e�Km�O�:W0O%������.�Q́�O.�4�;O�(P�>v���_���`�������t���}5!׹�F�+P�w�s�Yw�%ziq9��\�+Ə�#�����(/'��ѕ
b��/%^V[^�-��*�;,^M�ͩ^�Er�s� o=�I ޺zP5!�=�D:�5�u����֛a��,��f��? �"{�_�g�i@l�� ^8�f��{�׭������i�v���~�4���^( �[t9����u�D��u��h�)�ɣ�E��B�E��TfDa�ǙJ��o4OG��δj�O�}Gcg�1ެ1���w.��g����Z����{e���\n}�j�+D3w�/���x/�}�]�_���uY�=s�"�Ä<ژ]f_��10�f������Z��<�MW�	��Â��3E��q`��p�B`�SI	��	dzfo���?kZ�b�}~��OW��u%��$F��Y/2c��f��T�?���������ray{R�
�iLY=�n���0Ǳ���aMa7"�Ii��wv��:s�s7!��0�s�$v��i\���ts�X�G�h`�Xx�"K���>V>wz9�`��{�j�:��R���F��n�A4`����T��3,��Ԅ��+�ra�C�yf�TZ�+q&+���9\�0%�<��eѦQ���d5�[�wdf;h<�7+�![o��g.*5h ܥ+~���,��M2����
Zj#M�*�DF��EJe
�
JF�j���3�{����s��-�Ni�g�T��dA���R��מ�@�JŰ*g��ؿ��#)�W�z�6�������{=X�����f������%��"�΍v���
�8x:U1��*����]B��TY�k@-U�7�(~��ݬ����`��B�<�Y�G5�D�ǈ���Ӓ�)�2.���b���*q�J���ٯbr:��Z�'¶��i�v|�[r:�#F*6&�o�lF�cd�G@_s�v�v(}1�LL��Σ+����
2g��N���O�k���3��L�YʛF��<#gsˬM��ق�{�6��!����Aw-�<���q��)vk��9�V��㖩 ���K�O��ך���~�����!�;~ų���~��&�i�RI�x�':{[�/=s�����Y�!5�
��3@4}j,��{\t�H���I���|Vh�s[��͘�Y+��^%xRZ��?�J��܃��O_;�56gra���������N=�i���Sm�}v�w�:�^X��gx"簓�i4c�:�OI�.���Vz�xcn����{&c�a�y[ZNu+׵�g�;䡳�2�-U;Uγ݄��^Ԛ�o4GR:k2I����vk�5���:�1��f�)�`��x��z�X�j�1t�B����� -D�H�[��c�9��*���agPN�"��Kc+,�y���%/o��9�a����p>5��f�{9�����gum�0S4�����gsɥr5�r�B��}������㕆x�3�Y4�-˽�����<X�w�V��D��<�Γ��y���]��wٞ�ú�Dg���V,���݌�4Ք�^*��sj$�fJ#�GN��x̅�t������-�eCʰg��y[�b�HM��V�y�h��qw����	C5t�ڑ�}��d�.q˻nӻ�U�#"�V�p���n�cak��tP�R;��2\�Ɨi5�wR�t����z�X�\h��a��stv��CEH���$Z1+Z:|��3�i���α��*DҹvPʗ�1���V%2��9�]eڼc%Ll���d�a#e�1��
�	�e�		�*K�v!�������wy�DDUr�U(JDTJ�R�T�H�R4Д�MPTAV�(J�4ʍT����AZ��BE$� ���jk{���o6]�*��6kF�X�1v}l��w^�]� ;���N)t��� ������+��<܈:)^�Ŷm�m�5�,�h�>��r��&�uw;�]Ci�����L�OmT{�	��z�v�??26p����C}�s
���N��ͲK����M"������3Efbna�7�h�G���'׵j/�ܨ�����f>:Ҙg)��Q����±����˞c0_����R�ۭ&PE����o0J�{<�}�h������R����@n�����z���q���^�_��q�f�����Y���2��F�����~h�"�����{�U '�¯8jHW*sT�@;qF�E<��n�)y��ZW���[U��0�FǸ&��݅-���;BܿzŴm�<Ϸ.�Yq.㾳I�5d/��+}3@�����j�K��p�)�W9G����S��U꣊�m�4�W$Q���=֜�KA��>�\�k��͹�a~�"�	}(�5���2�2c
a�پ�ӃS1^dT��y,�4�U���Ym�"�叠:��ot��ykX�K���r�yu��'=��i����Hg�y�l���W6��B�s������n�N5����(Hi� �OE
��_gp��s�ieE�:1��r�k�^����[��x��>S9��Y�1�0「Ue�~ï
+,����	_]A�LB.��ib�748�~�Pu�w��=��҈�=�{�v)���JC���w_������s��#��l�%w	kJXyJ'�c/�b�� �g�u�w��;�}�D���=��@&��i֓�-=~�l�s�Rs7��HkQ�6 �M��] �CKst��+�9P�58^�bO�K���U�<k�*�"��=^��H�[��Ĵh��Ɖ�3����b�n�Z�ѥ7�e�t6s�Òaߺkv���.�yҐ짰�~f(dK{)֖����7�K����c���ͥ`�"ʥJ���}.49�x�<�$^�Y�O�˂�l�fwuE
Uղ�i���9�\m�|�΢�7�e�`�*J�<�eΓC{5K��Y��P��;A�yw8C���vb�òb d�Kkv-'��uئ��*��g��G��aź���Me��Ƚ3R�y!<�y1>I �QB�"ȋ(���L�� �"�b��*�,�RR�+"��"�ILmv�t���55 %t]�ݡ�������?���i��l{߿r�����T8�0u|�>�Kٔ<"�3��xD���|4��/a5�Rt�:Ey�]�	�y9o��9��R$�I��uQ�6w��+���n�b�C��mx�Aid�<=�Y��3Y����{�VS��8�$�ir�ՙwԀ��n����m)���^kӃ�;+͊J��2+�W`�4<3�. ,Ԅ�+d�*���l�⎻�O�cDvY^��A�]�H�罝�˃/+ݢS[Ji�L�@$����dss݋+�/��̵���Ա��V)藾&��3���T�VM����_�[=l�6`�3ۊ[L����U勊�����q��̭��2�lL��{���E��v����i�r�d�76��5u��h�1�"kOH�xyz^���D��(@�Mwn"�^q��~���q��՞�i�p	��}�k�+U����48�;/�}hQ>^ǸePo��l9���Y��*�0kW��`�(d��<�o�7��-�#��mW�B�\^����s�|�����;�w���� Р�է��~q%&��x�xw~���\�C^���L[�d�[�m����Y��2:}&��v�<��X����`x�
ɨ�н'Sjͯg������,ӛ�kjc���ez8�(G�"�}16���}��cEX��5��S�.�w������x$z|㫎�������L�۵2����Ϭw��~�5_3�\D5��N�gjY���&b��}d1��i@h�Gڴ���z4���l����,�H�}/����IWj������x	z޿dB�F۞ʂ�N�����v�����^��@�ؙb�j!�S�׋p�w���}Ǹ���
��)�UU��UHH���P$���}��	! x���E������R�^\(Ɵ�Ճ����;���!�	(H�O�ufv]�-
��8CɁ�Χ�1�;��fT����-HHp�|ݡ��}9�<�o��/��s���g>���x��C�Z�A�W�%����7�#���ff��HH��q���ǿ�� ���� �?�=��
�Ϭ���H{h=���?�A>�~�(�>W�������3>�9�4|>�B@����s���Rx�/�8Kg�,CS�(��z	��+�~��i%�0_�g��>�}��E�|����MU�ğ��4\$�!��	$���wu���	! b}����Y�J,�z�l�w���6�0�����$$)��B�ƾ�zL�a�)������:�������:<�$�����>��	G������_�G���B@��T�rz뇞�����W��F(���kҮw%Sa?g�_O��k��sI2�O�z�����}~?_�~sg���$$T������ȳ�~�a�L�X���hϪ��!H�ϔ	! ~���?[�Ԟ�Lp{����
x2O�����$�U��I��叮��G	��IHɒ��bI�=���1��_}���IPO�쁙�.�G��P�frc��0BHHK���oD��{@������� ���������?��C��v{��D�>_�<�Q����>{�}s��a�C� }Ǯ�=�F���JHH��=3�=H~�U$������$$
���k�K?�������g����yO@�y���wf�K����!r[𯟚L�����:��C>�����_�r�λC>�$����G��u�����7�_��v'����sܞ��To��{8d0IA��$��H0�B@���~DO\	�)�~G�o��y�I	�'��C�4��{��ML�:�'wK�;������	�e|�yBx����rE8P��C�