BZh91AY&SYk�HT��_�py����߰����a3^>�   t   ��   t4 
  ` t � +@��   A}�� "�!m��QVڈ�*�T����(�  ���!$R��s��C��j��6c�p�]��N�v;j�����tu�+ۃ}�������֝�zЗ�!�"kO}�P<�U�*킑ݽzTKv{���Ծ�}�pʷv����q+pSGN  '�E���^�MF�$lą���=z�s݂�ws��wv���b��
�n��L�hwg@l:4�k;���k��{v�Zr��v���t� �S5=G�=��]���A�m��S�P�z;Բ���\p� ��r��9�]��gm��u���=uz5�v��{+˸b� � �UbjP8��ܬ���wc��ǣ�]�֛���gA��wFv5]\(
�·l�����MV���;n̗s���Pw
� �I�A��7���k��ӻb�>�wy�/}ý����'��u[���c:�t݃���]ۧ���f��q��
�˯O��N�>� �     
�B@ 

  ���AA�h
���`                 xJ��g�R�P� 	��    �%0��UMQ�  �h�`   i�R�iP@  �2d   $�RBM�@=C#@ ���  "*B ���=z��G葧��� TH�IT�Ѡ�0�F#!��1�&����и���"��t�0������,�>PTQ�I ��H������A?*?��������%C���EE��T��/��?�G��G���ڟ����,�V�?�*M�$H�Q������m��6D$���Z���K @5U�ߍ�%�@@u�C�_��������߰�Iݤ���f:Q�c��D���Æ31����Ȟ�����=0�'�aofN�p��צ �=1��i��}1�<u"8t�D��"I�|�1����c&9�
D��Y�J(�"�,��	���D~D�&�1��@�s��b>Ɏ�<���rb	���%�3И@�f:Q� �	�	~������&N�L'�{s	�&��Ӕ�|�>����!ӥ�xo�����'
9RM��0��.Y�H�|�"p{ɄDVa0N�&(A3�	�$/���x�^LaG�f0����|�1S	G�D&OQ�<>�DN�L<'2T��a�f$���a�0}���%.�p�A��27�X��%�X���<GD�#أ�7d�o���$K!���ӵ���"sЙ4O��ė�`�ag2�?C��Ɉ��"9	��O�aҸ�ϒ�,�$�Y�_��H:1�?c�ɘ�Yד"\���}0��"X����!:vQ:���y�xK�c�pN	��b�<��C%��ǩ%<�X�^3��`��='�Aӑ8 �Ĕ�$�Y(�U�.4e�9�8p�vqżˊ��bc������"cُ#1���'������\��ވ�%s�	�}eT"_�0�5	�#�#�DL˘������E�2"���+���BYC˘O	G���aBTGDF�a��ơ'����"p�A�>�D��@�33��"#1���.LaBz�������.;0��=�B"��,���J'}1D�ʙK9���D��#�̉�̉�FTŉ�=",x�By���/������@�~HIy���&�%ʸN?cFp��:tD�)�w!$��F�'� B~zI?BN��G��֢Q0Ly�ad�܊(~X�P�t��N��/!(L�� N@�$9�,�b",Fa0��_G�?5���$��@�#p�gN�#q�������BX��Jt��H<KQ(��,Hb1��	¾�P��q(�ǉ,~DN	Y1�P?gD���":q!<�J`�����Δ3�?!}�&I)���%���E��	↮'��'�z8Ju�JY�/Q8#	>C=��?�Nƞ$�\ƚo��1x�����F�"R`�������@��=8p��'DOG"R��=:/Љf|�������7�ֱ�y��f�K4���<5ɇ�g-Lt��E	Q	�x'G��F�afS
�/ݘD�Dn<����`Fa��c�0�g"�(���F���D� � b>~}2z8"B���'o�3Q�
�fR�H�r%0�oИ����w2�"(�m�p�s.q����'�rⳖW|��:�ꞝ�����4vI=�zvjS�`C�>�d���E	�8��L:'g�rbz#Q�Ǟ��K�a���z"<#qN3�o"S���O��ĢU�>({��)�Ѣ��Dj1���?"O�D�9	%�E��$��D~NL#���>�D�d���?"B���:�M��gc�0G��Ʉ�E	E1�<pN,M"[Q(�,�ɔ���rb�	"S��Qț���`��)�;�'�q��C�H�Í��O�6'�12"3"&je(��������H�!)bdD��J=��'�!�0�LJu�J>��D&7¦ ~< ��>fl���Ba�`�pN	c��:py���@�L�I�9?1�xK)���,HO?"$����т&:K�D���#�Ȟ�i%3�Ja��t���G�I�Dg���p�=LǊ9�N�q�I[3$��r!8#~�O.La�Ȅ�2�����!�V�tHOf'�x�$�gR#���c�q�̉��yp�I6c�ds��TM'��oI�|�>���`���RH{�R���8[�R�Q���Ӥ���T�o"x'N52I�����)����r<'�ȣ���K32Y>������8�g�y�RDp����"�$f>D��9�b|p�r&B��C32�$�%�W9:`�2�Ì	s��s:LΔ����	���lDG#	>�DN�73)�a~��P����ɔ���ǹ38p�}p}�X��P����~��N�a<#�$�%�(OL"=�r&��bzpG��~����?<�Dn/����F?G��D���'�8%��O<ȟ�~�B'��D���舉"a^Ģy�J`��&ı̉�1<,����H' A����&؟8q��u�J_#�ŉ���,o�=�Ȉ�$g��&�ĹH�f�vrN��3 ���]B'{#p�s�#�q10��<91�L;$4Wj���Ӑ�rN����><}ߙ�I^D؜:'��'���%�ĥ�����1�8��ȖM�"w�{�FY���G��x��8TQ�N�ӧ�����Y=8I_"u ��;TB&"p��tf�>#�	����$��O3��/�G[����:M	0QP�P�Q�_�N>��܋9�<t�p�3w��ZH��b�`� Ç�$�T �|�D��&:�I(�D#��8D&z:IĈ������H�9	�و,O<�0N6L�P�@��$���X��#GJ��tN�GD�1"#0��a�f(��$�1d�$"G�
Y'�$���P���Y�ncM+�1��4��i��S�	D>&Ix�ID��H�Ӆ�}1'��VL�w0��>D�0N���-%$�>"�;�!873	"eׄ�D%�I��� �L|��+�8_��;i)Ҝ'�3�|L�*���a }P�� ��\rc�^�G�0��S��Mb��f�%�ƃf*������F��A�����#��	?_��.�?;?g�,:P�a�9%G򛉉�4^rk+���dc��>�k�g=�묰��7E�#�̱a�zh���k��l��%Ep�:�~��s�6��=�!��8��rq�����g�Y�E1b;�ō�z���d�>�=3x9�����}z}�m��ˍ#|�ZO�ďQ߳aʇ�/����E�M�ya�}�=��y�Q;��O��)7�}C�I��/w>��9���\C�?A�g�DN��v⇊]C��	���>X����i�&�����j��mdX�ygz;��6�vL;F��G՛�����Ѵ1j�S�LX�G���{Ѕ�����4B)�\G�4��!�K~�N5i��.��Ld��CJ�^8� CL8CJQb�eDB�ݘ!���vv�#�]��Q�����taB��p�]2��R/����H3EB� �b���dD!V�O)��!��(�!8d�"�Go��F"b�I����A�B�/!��
3�cPt�AB�>�F�ӣ:"�
.��b>��ƍPAҌ�4XwY��.p�M�B���Dc���NC�"��ј#M��j4��h�A�~�iU�b��xmUN��m�U)H0���g�ѐO�d�A\QM�� |���f1�)���? 胆�@���8iHSFi���HB����DCO�3M4���ьF��Y�1�Lt|�Nw��T�팷1D"�^!�2<Q�SR��Ae(��S�)h�m<����0�3����X�1���H�w�Dh�c�FC�)�&��Ҍb4���d!A�!���#H"�4�<���A�,��4�)H2�i��(�0d[E)FBebH(�R�HM�u��!� �<��"�j2b)� �����3J0���vB��2�!0�y�4�DBbdFBE�d�@e)�J��Aã�cKH)�8pa�a��4f�`ͪќ>A�zg���D!ph�e(���ot�4e:"������E:A�c�OƐ�8"����#L�*�S�i�EmӨ�Ψ��M��l�lK9��~X�g�1|v����ͿG��3�{�±}v^h��l�(�	�=Q<�{���<�=F�$:�,���r�POK�Ou�8.t�Ґb�B������q��ȟ"���%��7�%���$Y�̈�f�M���#Y6��Q��/�Ae���w�i=�r���q���Q릤6��F��V�,���B��4޲]'�w�čh<u0bk�9��҈F��L��&{E�ϴo�K:��}C���xz��Q�{�e�q�ߢ��7��g$}�����{�r"8_��Y��7�p��C�s�w���V_L��������3�S��!!8Ũ�7"��rQ�:��ѽ(��z���/��q�č �՜��Qޢ���z��k��6!�Ny�}x�2�ә�S;�0�f�M��������G��Q�gh���=-e�>��q�?�y�w������N%�b��[�z�{M�rѮ�,ΐ��/wt�����8���}�r.�tmiy
�+�9�=I�pY߉��ihrQl&��P��~g[=�%F�s�b9qN�,�7zN��y86�q}�ʂ��FԖ>�"�O��q<�|��~�?R�?��b��t\�ɜY�7�&G�}��M�<��D�\CA��
���r�ȉ��{��#Ϥ�O����̻D<�6�^q��v�Q�%Nv��-f�EJ��C�{�U&���Qu����}C�	�\�>�c��UE��i\=������p�w9�z��K����y;I����5i����d$9
�}�P�ϸ?��>6�>&�H:*������]��I|}�)Ӎ��_�?�>\��?s�Y?p�e���u�8�矸_2�7!s��m]X����g�U�<���8�G܇~gϻ�D��<Ϲ�|�W;�s�����y���s��r�����p|C}?JN�B������q��:ˆ��č��+��Tw�,��9�M�׉���<�ZO2���O"�����u�\����٧��#yӚ�3R�0BL�r��G��6����EG!`���=��w�YQ"��B�,��<��k8������y�g���	ٟL��}s�{ȩ�1�:�4}�q|5�u�_�UVý��gu��p�j!}B"Q�=�C�e�g��|�ř��r��?p|Ӎ
�Բ!ss�*Y�Ig����v�3��I�!��~�}s�:�#;�'G�2���8w��F�f����&��k���:���>f���G�3�Ĳ,u��뤽Yq�JZ��?B�R$��L�=8{fr�G�%�g�u��yg:kd�������ӝ�ݛ�����N�I���X��������+YQ�I������x�Pl~F��/�g4�|{/$5�����Ʃ�\K'YE�y�C<�����BX6����̌��2�
C�t�t�gw~�.d�~hv΅�Q�g&�_>��a~y�ԍ�����NJO,�_�=�K��h��������>����g�:C�;�F��Ѫ-D](�=n6<>d�]Y�7�{��p~�'�Y�(�t^�u��&(����#ч=��;Üү�<��-���>�-�ϔ�����1f��������N��'�~�?<��~��<G���s��_|��R?��xO�~�a4~'������o���ܨϫ��w#����Z���ڗ�jf�``���'�{��;+���y ��FEwћo�N��~�n�߭�^�v�O�S~��w��7Kϟ8oz��}����oI�s���{���O��&��k;ӻ�ߑ��F���Iy���y�[o.c�X���MR�s�9'������^����^o8��MM)"=��>qvO[�g}�����o�g�������v���ߣ�������AX���!��l���sb�1�ߤU����i>��:����J~���rj�F����g����x�����[����y�=��\��Uת�7��_rsWu��:����}�o���=6�^�󕵰[�-�qz�_��z$�x��7ˍn�e>c��^Q�l��-r�O�'�q�^C盧��g���3*{�*���ߣ������Ǽ{r"�9��x�=�vo���=W1�Ț���O��}T7<��ˉ��~�|��7�y��w�~�9��>|��X����#������ډ�8�h����U����7��]�g�˲!�˜����pr7��qO�6���j����4�ݛ�_��_}�{T�M����wM�ߟ�������6R����x��}�s�S�q����g��ik��E�i�?�T���r�{��%âeqr.N��}��9�ݷ��]��*-٢�k�n^�y�r�ls���o>�$❝^���_;���W�G}Ne����׽�Ȯ����iM���|�n�˿?��u+WԆ��C�{ϝh�k�y۬��q���J�Xx���x�EW����!��;�X�c���;u�at/.�ܡw�����g>oY��[=좞���$s�%�|�y�)M�#y�&����%�TSQ�Iz��/�D_�_]��w�{K�ŽW�%�55���h�΋��������͞���7l��ywRǟU�Onyw'�ʾv�7\�q�b��tɞ�X�'��?�B��a	���O�	�i��G������2AT��MJl��&�Y1�p[5���r�ɸe�D�!���D�Ш4IB�[K[���ctΛ5C<����1�h8�&兮o-��R�5��n� d�%�U���z"eoGU�۫'ɋu!�bfԗtj�:�	�l����xT����E�G��ǌM����"��M� ��'*�Z��o&q��LՕ,Y����/6%�;�٧xkg�qqU�����bF�&�5Ƌc����gD�E�	Y[[�
E#p{�wcF��(dmXⰢ'��syq��ź�D���!b�"5(��~�H�ۤt�Pm�&�r%`��$��A�Bl�Q�g1��R�̅B�}u/>C�]@�:{�{3EKpϖ�Cp�$'�Q�ww�	$s3��50�q�����0K!���]8�XwsP�e��i�QV���M!d=x�Y�����=V'R�E�cA�|W����,����������&؀��e��S�^��!-���ݩ�1�^��j5�lѸ��<�%��UuR�um_}r_����HD:�'d��xq1m�V%]���Y�T+t��mpo�3��9�q�gd�J[bq��u��%�@y;��P�����̨E�r��U^C��������܁s�j�5%8���j�v[��q�J<8��x^����y�ޏ>���{p��:�X]�(�<��W�==���46i֝�u�|�b��n�	�����Q��RŬ4�{M�Y��Sńb���R��-����n�TV̒|�K��-q�/t�8O��S�<�r���g���У�XU�ϋ"������g˓���1�P�J����r8�F������#��A4���eL�."7�����&�	^����*�
;]�m0���t�Mѵ[,5j7T�
��Zܶ�f;ņ��IL�?]��;e,rT�`Ą�l��n ݓ��D�,,��즇DU�Y�͸	�Y�\>�����!�<�=�@����ىdGY�U�L�z�o��x�F���Psd@�MgPu4@yub��ƃ:��ė�A���\�q�Y��u��0M���s�7����?��H��5$?v�ZTTQ�?О�~_��J��?W(�D����?�_�:��?����
�����K�o�������^*�VUU�eU[EUUEU[�.��WUUq�U[YUx��YUV�UUQUUQUV�EU[YU[Ͼ��DdUB@I ����{�vo��U|�*�Ux��U겪��*��wswj����������ZUx��YUVՕUmaUWUUQU�����>���>� "���>�^qEUUEUWUU��*�|�*�Ux��W33.�j�U�U򲪭�*��*��iUz��W��UiU|�w��{�����Z�H��ȉ�C���n���ª�"���������ͬ���ffe�V�W��Ux��YUV�UU�UmeU_+J��^*�Uz���}�B*��#�(�$C?w�~��۫[[YM$I���}�߯���}��q$�_�5�O翉�?������د�8Ҹ�I ���:'�N,L(D��ab`�%���OxO$�%���D�D�(D��K�'Ȑ$�8q�Ett�U�ÇW�!"H�B""&$`�I""$�Bp�:"y#�&&&	babX�'K �0�bxL,��:t�8$��8"t��"a�xI N$�$ �_J�8'K�Ib&	�&%�<t��vD��r��[e���Oi��n�V"�N�X*$+jI�dD�XZQA�6([r	(�|2�1�,gU��l����r�"Q�Cő+de�%b�z�pcy6��7*DMQ7Q6��y-����4CO�
���Q͸ª�E*�! у�2����(�8!��B���E(�["���R0Tjc)%x�JB�B1�B A��|l6��4MįFR���7!�D1���i��U:��!�X*�"��M��9X�B&�&2	DQ�e)J18�I��$��X�
2�dPE�bJd+L�Q�D&1b� �eH*� ����R���dX2f���D+ ʮ�Ӛ��2�D)G(B�У� Cld$��a[-H�!F�B1��ԴeE)!"I�ٛ L1��9�׬�vEn!Q$`1!�L$a���6fY� U"Ǜ	�K,a��#�1!\�_��c��Q�$TW)-��f���41l�m��Ȃu�R��	{L��83�a�L0��E��[hƦL�R�L�!����v�Y�,�����X�HǞ$̡aō�]-�M4�a�ÆB`��(�R�
8\C��JYit2de�eVFvK�a����k4�W�JH�a�t�r��1Rc%��))`�	IIGD�� �)F<p����4׋F�>{�+��L�Jǘ�`�ex��&Q�QA��U.�KN͖	��M5�v���� N&�0�Fef�C��d ��8����75�b�II��Q�R�H'
�����7K����Є3q+=�nN�:^��ǘn����K�b��9ݘs/�ͣ����K,c���1�f�Oh��ګnBH�fL�X�9�fq����YM���4�%#n�wG�+h���'MU��R7lݶ����f��M6����M5�7[R4�#�HWt]Yh�l�14q�!�B&��5�1�ԍ���Z��l:`�û6�i���ĩR�k�4�V�)�%�]Ρ^�V�fib�:�Pu[kE`7�1�E�
HVT���CW�]�x��ee�l���@�If��F���4ڹ�E=�Vx����ۖ��;YX1��� M���y���[e	{Zz��zZS�Qq�`��b3uV�v�HW2��ZESB�������,U��p[����h�N�ʻL�w�p]ېc(�C��'e�J��D��XGH5!]�HUͪ��������e`���,׵`�fm6�0�&��	���2���V4��0�Y�i�a�Ӿ��o�������t���wwwr����GO������˻������wwwr����x�E,V�<l��g�:l���%a������y�W��LA����4	e�g�����"�	D(�Ҍ�(�H<p�LDDX��	�d�162R,��İ�B������+�K���(�!��)�oD�KSD�cLYFQ�̬Gl����(:n$�Ɔ	�)�Y�J�H��sw)���FG$�^*(�g��e"�y�����Ud�H�GT�u���*Q֩!ȭ2���<�{�%�a����,��8kmy#e�����Ԟ`ύ���'"4C$%u[SEI*Uރ31�����n�����ҝ�c�t�|���{3�N�����:p��{��[�d�9.�G<��u��������a*���鳣��m#��g@��E�d�͸6lb|��E˶3C�s,f�A�����w��='hA<>۱2d�!��Q���:,�CM�C���8d�х�!���U�T��0�Hip��̖0Ö��T�l�6�$4�~�g��4p����"@�BQ�0Ox��ȳ��>�\BrE��h`# �0�)�%�]�d�c�B�7)q�|x��LT6n�O�,H�e�O����dAa��9�o;2�!�Öt��F!���'#Yf4���;�2x̍�2B�T��!�Ƹ[0��鴕�_��>9s�:Xzd�(�Y�"Y�DH(J0æ	�$}}s��Ǆ&?m�������l�-�b�����x�ɡ3�/�Μ�ca��l�4;o��bu밽�,xbb8&�nA�����h���s&pu9T�������!�>�̣���k#C��ʎä�.jax`�6&�$��SU�&�hގUV�tq�MD���8x���"@�BQ�0Ox��Sm`�P)��M��sLτ�L=�B�(�S�ŕ	�쭥���Hh�0�ۆ�#eQI4x9pn1����4ds�����c�C��u��.���J��	�s|imi�ޓgS���:[[�=�HB�If�O�I�;6�2d���<'� D�(��'�<Q�g�")����#���c��:2i4L�
�M(�UL�M�#C]�>�!1Bq��u&:�yR��	�lvLP��WZ`�jh�Op����Dυ�"7����:RPݾ�Q�%�7�鼝�y�Wvi䗼�=���9eGs�L�ם�wi�-��~�;��p���fZc���z,��8���Ja{�mӨ���t<�g|���a���R$)�#E��
Xu�Z`�-�s-v��7��3���idf��D�����j>cϚM&@H��E	v�4;h���(t&ݙ,ᣆ'��$�%a�� 嬁'���,���^NI��Ǳ�$#������4��;iш?f�x�tA�-�2�Y^FY]�w�Ω���l����u�.�	��0���`R�N�p\$�c���v=����C>!E)H��DȜVȩm��p*�K��>8�!��mPۦ��kI���� ̵�'�Q㦝4D� D���8t��D+|����� �ÇA��=�T5�_ �$c 2ȵjU����>�M��U�̫��%p��M揱�̕��Zf�2֓RGd7�'�,&is�s����2�l�T�g\hȆ\͸��hԛz�I�N���w��CS\��lzS�����;#N��<af�i�<@�%	Ft�<'AN1�M53u+e�jI��b@lpF�Q�-V�)��)��!��3�0�TZF[����c��I(�g���49�5�x:mvhr�͵���e�mxy%;0錖O7���vܺ:�o�ݴ���.MɧYzUhz�=��r	(p,pp��&K�����-z_����Ϸ<a�&�:h"@�N4�맮;qڻq��ڬc��I�@����B��f��Å��Q�.4R���2�Y1/(�������L)�)8#��j>����}�
-��E���զ�t+����(� �b�of~Hx�uY���Hi�k]*Ma�sm{��!{�*9�l�R�x]���o��N{z���;�/w���y[���|3Ə��6ݯjF,��;�b��wd�+9,�BU��2��Rn�Ӊ���R��K�1��wR��I&�4�W�v�/A��xl�r���z68:�c�E� n98ʽJ6�V��BZ�BX�)�
BJ��F���d�f��x����Tʏ�Hoֆ���2p�5_m���}�pD�ƚi���"@�BQ�0O	�>��D�F~��Ii��ƥ43���r��g��<��T�ʑ<Đ�gG%9cs �g3~�����)�I� x�C�]*��Th����6BBf=E$R͹x:@�ƍ<�A�
H8IP�٦�Y��*!Kx�b�2D�c��94��u��NUs�Ҳo|MIĦ�|��M�<τCqrgQ�86����h��9Q�$hA��0�4(�4�M�O�'L'H��$�i:E��$ᤤ$��i�a$�:N�⨍ ����M��t�t�,Ҥ�t�N��f4'H��sN���j,ڍg�>k��[|g������b�_��q;����w�����<ܴ�t�g�(�t��'HӤ�l�i'��ŗE���	�x�,��O���^��G��+�`�&���i	���tI0�R4�#�L+HN�O��4�:$�E����IY:x�:mG���d�\Ɠ�h�Y>#K&b7�c~����1�L���>b��~c?/O�+��h���t�ǌ+�d�$�L)0JK%#L&�4��#��œ��๤���bhw�����B�=㓪_�fn����v��}�}	��}~�����Sc��O��}�s��S-=dN�o���YzKGT��^uD(h�����Mp�{s�{��o~��>AW����r{��<}��1r9}�"b{��L��{|�Qt�9�\���-$;���U�7����ɺ3�x�畿|{o[������n�������e��������7w33.�tt�wwwۙ����:}�4�MO4M$�J4���k�������]3-��m�J�Ĭco�.T/dr�4aB�?5JS��ٓ�0�ZM�:��hL��}�'R��0��U�rL5!��G/Z�S������#	��M'v�O02A�ƚhNE
alT�ǫ!J\�,��*\��O���<X�i�tM���L���H�U)5Q�bR�r���2z���OK��I��&�'Th����7�`�6�I�:X���r+�S��T���Û[bK�J`!	n�C�s �^ꃬFhS ��6ɔ���~��sqzLI⪵
>,�K7I��t�$U�����70�������>~v��>I��iӂ'��Ό�>.;؃��>��ͺ��'�m�UQ�ae?RjQ�(}��*��20C#��*4�b
L���փđOS�M,�\����JMK4��Z<!������~��oa�t��u(LVt�c%I[`�*�G�t�Fҧ��t�K�m���2C ��)rǌF��o �31o�[����Ś��:�]䚵�fW,�Ŋ�m���K���ɹ�_i�N��,q�=�L�� ��d!jo���tV�*�1;��m+�~�I�Xi���b����x�nc��JmUSG���5V�,d��3
�M���W����b�P�d�x��'�Y��l)
j���R[TBi(�Z�����%gOM����'��'�����4�M(ӭ��<|��j���V�1�M�������HCt�DB���F��c���D)�.���DVl���2L����j\O�cq�% )���`�CW:�c+�z\��f;Ya�(�I$�F�Rt�� �h�\K�8t�9�?6�ΖD�=���]�>�����D�����E;��yw��x"2z�yf���|c���
.UN?x&ח��sI�4�sE��>����>:ƕVc$[�$����,���#�US��6� "YId!�(h`�/c�6ꄼ�Ul��#��H��Pm��1URfL����[����ISc��Q�-BD�A�i�EU�F&X��1m��P�UN�xx����)�+�4B��:�X�6�<i24�l[%�1��&�-iUFjhj�Tbɞ�#?7������'��RY}�}=$��@с���/���;ݚF'�-��"�/�0����N�Ӊ��3���������$4/�-��	��Lj�̑�c+�����UvE[��`��0��cAc �&L�j)��O��`��������4�M(ӧO	��x���]]�R�y�	$��nnm&�ɖ̛�:�7��ܱ�SR��A���f�V. �T���̜1zI�����,4{P�Uw���i%8t���j�#DVX��e̋55F�iUdU2YK�MM��%%X�q����������Y��Y;�i�Yl��L��;Qe�V��S(aS�Ji`��Ua1M���Q��5S�R���l|�F�X|~gDLd��U�:�,�%��n��ɺ��j[��;�i���Y
i��1�Kmޥ.(�˒9(����ꪡR�IS�T�bY�^2�Ø�GLB�QV�B��������� ��d�{��&�p�Uk Չ�ǚ*�����m��0����M�6(�^�ۍ<z�����DM$�J4���if�����d����I!C�C�oZ���6��<�y(ҖĪ�a�J�g�pac�Ƌxd��:b��w;Uu���LT[-\1(�f#Pd`�K�)vR$!8��vE*b$0����c#�)��V���@�����\��7[ۤ�c�WDbB�'��D�L'�Q88q5�2E��#:2Cj�_�^/�ʔh���7��p����  �R5e-0�F�(j;)*a�Jҫ���<�z��ש��1�bh��0nX�6�<56��c%L*L�*��=m��1�M$Յ�*�2b'���ևU�u2N�[�v�,v��\7�#�4Kvd))��x�>�[45SJ��6��J��)�V��0�*L�<�Z[k	�,pP�Y|���@<e�ȿ6R��lP��))���rH�����~��4x������ѓ���$�J4���if�,�s�MF�E�����!�~�y$�B��"4�#��q��2t���X�-%�zf���Z�\�lTS����$��$M�)N1�Y,�0�KR�׶���1Hl�Q�?�?!�*�6^k|��7.���H`"E��"�-d�)��e;�SR��=+�n2,`�5GF&�%���h�*+J���i7g�Cّ=�Et���:�ឱos����2ʬ���)���׍�4�y�\�q�V�T;��
>b��I&^�+,h!�Q!�C.UѺ�V$y;�~q�t鹇J�JR1D\�W""�-պ���J H��cMZ���f�/�tW�:�Mv�nc��Jzk�K�t��d��|�ǎ???;t�M4�M(ӧO	��xڋ�#��A�@���)`��2��Rı�G��6m(� ������*���0�(�1�Ո�״Q'���ij&9c#H�ȝl��&xl���6ʶM(!5F�)�I$�!?ߏ��77�i�E$b8<��Ү�n��n���a'���ݟ$g�xkʖ}��y'1Dy���>��_%�a��?������ﭽG���5�&�3��>�d��bV1*hє��x���&��f��D23����>�<���t�k������L�.�o[@�3�򿭄����1 ����Z�R��i�
x�ra��0qG�.ʓG<:2k�.��ˌ��4���JmS��ګI(~a��Da��a��>�R��"���Z3���5�Q�Y�Ɏ���b1�z��j��j[�{���˒^r�e/Ƀ�w�^'F&��eg�1���1댦=!��,�\��⻱F��Ip��Krf��^��}��>+T�*UL��Gnޫ3/[0����N��~,�񧎘	��M4�N�<&�?�'�k̨H�&�E%��u$�A=
5ێ7�>6m��Bi��Ń� B�-�dh���^F�!P�Ja���a����K=)�S���fk[N�7+�[���Gq�i����3�*tܵ�ӡ�I�x�n4��7a˖I�ݟ�x�S���'ZO�.r��#�fiù��!�`���D7Qd8g���Y�chq=�b)�aij��կ�����+Jh9��6�>����EG2"��^�95�яx�O��=R�Q�o�d�A�|�:;�l24l��}������~<t�Oƒi�iO�����_�n&���d�N䙒I B��ь����>�B��~�^��w`�V�4��ɽ���'⛕��Zq��4�*j+�b�Ru��~y:U��<O<��A1�d@�c2df�?�4�>�0��N��-1\DdPnK-��2e/rI&��<�D˕6jX�Z�Wjt��ыXrcr������U���ۀ��P�a�[q�|m�VظU_�G];[�i⥞[�\qn�ʛ~�J�醥i��2X�mC���8b��		ܲ�`BCH[�If h�T��,-��x�5��s杸���?;t����M4�N�<&�i�C���AI�I�RI$�3����S�����l0��O�����E����a#1 ���qi>nk1�!��p��$�+]8b>6YԄ5
0m��L6�_��!M+����}Q��:|Ɲ&8mm�j���LT��ѵmXR�}��t��1��S��U-X��`���9�}%��{_e�c��хZt0<d�$�ܨd29i�6v�bW�)s%�Ͱ��M��irM�rgy*�ٶ�M^M�d�4C�GNM�G��b���i��Ѥ�D٤��t�t��	)���?��4 �i)����N�N�di�%��:F�&D�$�8N�I�I�I�	���Iӄ�َN�i&��4�'���I�M+HJ�М'I$�HO����F�4��(�Ѣ4�6cf$�(�4�	'J&M&M'HӳmF��i���$i�	�ٍ'�Y^&�8x��'�||t�����N��I�t�(�IH�&2cI0Ѩ�8i>#'��$�s�:i0F�N�1�L9�<i:a>,ڈ�6!&�؋g����>���+3��������A�I�'B:i:tҼa:Y�a��o!4�N���di���/H�?"n�����}4�t����[��=K�geD�C�X@f���=�!�?���G�`�uf����(Zh��&���3HpA�i2�*!D2 f1� "�R�G[#(��83F"��:Q�
���b�T�4D�4D �e�ejz�Yd"9%�	�ety{�7��qؾ��:i��=ɓ��vC�8�8.��Bpg�T"N)a��g�1��&$h�o5���ן3�j^�8�>��->�>͚3���uĄ�l"�vg:�����w����5��|�TM8#q�p�}ڏ�|��5�Κϐ�OM-�2h4!��������8"u��k+Ǌ�`���T�����7��_�w����l�w;������J|����V��]~\��f������29ü9-O�{j
E��>����p��ff{����^�����D}LO c�%.���K�D#��7u��mof-�B*QYM'�������\d�c�`�w��G��2�z\x��ah�6�f�rhӛS�F�ur���E��{9RU���9��.͵� �%#7^�H�d�^�T�l����7�MX���q�%^�e�ÖO_jy�p~������_�����ª��fffn����fffn�*�������@��&	�i��iF�tD�������\b�0� �q��J�n��c24�BW1���e�.�ь�Uc4�a����kLBn`%	��hi̲�# ��홴��XM�zٺ�k���1���t����G�KH,� ���q#�����Ya,#n���Cu�-�鬤�1�C�Q�'�
X+r�.j���X0��V��j����  ����6��k�ƫ,�M %t,���3$m��[Ѳ
d�8���ƒIb
v����� N��?&aot�Y�1�ѹ�a�d1��.�!�:SGy����T����k�����go����UI���1�i����{��u30��y,�p��ږ��۷J
O�|��$�6���#��t#���~�!T���ӂ�������InpA����H�LKr���L����3�֚�qho�ŗ-���aܙ��ܡ��!ǚ_����܁!���J<�?��R\������@{'c��N�e*���ny,D�Ag:Aℳ���'�M4�<&�i���yG�:G�"">����2�N���%��AR��S�P�zI��Z�4dJD@�4�]��CB�~`,�{��(�����h:I[f��il�go�p2=%��8m��:�p����^}�d{zQ�؎�#n��I����3�t��3�V1t5f�e�
��4��y|u�*[�;����u�h�m�@�KT3K�8x�*T��l-�XvD�t�i���LOĚi�J:"p��t�p����N	Sx���6�g�i�6�a#�~�<���$��x%�����͙��c�ra��i�N2<
�lv�l�l*m��G��.����!�n���0�>*߽<:rxŢp!�F�?�Q�����4�6�=����%�,�3�gވ���*��%!gad�>6@�Y��M��[w��%��N�r<ɠ�nK	�f��.���:����ֲd4푆��l��J-��FC�u���3�������gN8Y��i�$�4�<&�iÜO����VD��ğRI,@�4��ܐ��0���Թ�^6e�2w.4{����:cJݚn�������9 �#S��g�yL�6I�ܿ��Y�ی���m84�|�(���\��k{L9h�"dxW�$���F66�{�UF������6k$�
p��:�f�I�2��]�]]޸ljǍ⎾kI����]m��;m���6�0pW�N�r�Z`'OI���Ma�8`���N>:h选�M8iGO	��t��?Lυ��%ǅ?�A�h�1�X�Ȇ,�8�=B.V!�$C!Ş]��q���(L�Ô�=8C��;�X�5Q��UM��w^����x���KK#%�\M�QN�J��oYBm1ua��:|}����9�� �Ev]{��%N����I���Y��yxtBWj\8��~Z֐�/�I�Z���dJ<.,RN�G�#+��,6`tކ�lz8L�ۓ��>,�TQ��f���I��A�t��0�~>�R�oFM��]_��O!��S��V<��I^�7�f��ʏ�%H��t����ݰp�R�N��ƙ���e��)��'w�oI�3��e��Gi �	,�:��J+VR��BD���u���v�����(�s��Q���̥����NS2K$��'��:`"A��p҄�>??Ut_��LB��o��	&�*�U$�0;I��:��D8I����;(�1��TS��#-��*ڬ�b�`B�`�a�9l��͌�O�//>��R�On�B�gO��UU��4t�Jp�(2�0pI��n��?g�g�:媪�M[eHU,���x{�Q�S���e:(��s�<4;M�XHi����h��z4�(��-������v�\���p���o�m6�Ǐ���:`"A��p҄�K4��	�=ڔm5$��
c�~�X�d�s͕�w��1�C�	c��}$����۠ۓ$��Ym٣e�p`��|�>�������I�O1�J��������*��T���������1��I��g�eͽ�3�*��ʟ��f=y;a�7�ƞ.x�6w�������3�(1���p��������ɝ�AXx��u�Y�s���dnRM�2Y��~�LH?i�J�xM:~�|���I�9�H�G���ޖ�|wwj�T����#3��>�kC���c���&��L��Bx16Bc�!2\a̻��i��� �|:��RGݲ��fe�Á��}��_=x8!����O���3�M1�P���7roO���4=x@�P<v4�|:L45���풴�=4�n��'�4�!�Jl�LY���ǎ�2p �M8iBtO	��Y8Q_O��������R��76�B���?����i��t�E���B�lN��Ȧ�mQ�;K���Yej�e]���vtK}35��^�I!�6U;�EN$��B�t�w�E^X�7O+��>Y9՝K�8ƽ�>�z����.�#�<��٫�y�^���_}��ޝ~ō,i��!u���ߙ�L4�F�
����<�Ul놝�4�s�;p���x�Y�Ph&��-�^Վ����x��M���l�zʄ�ɠ�9~t�?K����G!
"�m�Ǹ'��Y���L(�eل�� �shx�b:o��)z������9��1D0��0�5bIS)�� )�dz�\\5&�1��^�q��0 M4��K7쭟��}ϫ�dY���)�̃ �XʱA��q�vI$��8I�&��,�`��<S%t|l����CŴ=����F/	�����'#_�����ᲃc��0x��V�nZ ��@ܧJ28e��t�j��;������U��.m����A׮�ox���L[���Y�x�N�jp��-i�)0/rh̪�kr��<3���`;�2����Z_4e/�m���U�|���1�<}ջ��>b|F�N���&�&��Ip���3�����_?3���?<c��gkҨ�L1�:lƞ+n#J�4����$ӅpӅI��1���J�f<DƓ��+M'HJ6���i:I�QDѤ�nY���zZ銻��-|Ϙϊ���&�'J$҉�4�6c��9�i���,�(�H��:N��QrcN�sOLi��p�$�#���ڏ��tJ�0�]Di)Bx���t�~�M*��*M%.b��6c�4ٌ4�O醕���J؍%"�6�&`�J�4#U��k�ұ�1q�~Z���3D�H馜9�I�*�''DғM+I% �	�4�?{��Ȉ��Fw���Fi�h�C�}�{{�?z%��oN�����Ͻb\n^���MDz���9�(ٙ�G��o��k���9>�6g�^vc���&ս����3��1�s��_6�s��G�l2�(zV��Uŝ����j�m}cm{�utE�gse��W�81߉����j�{�=]�:���y���������۰��^�ffn�ʪ�nfff�쪮f�ffn��J4�L4�D���NpN�㧍�,&��H@�<j�US�����6�a�H�0h}50�wf�i��t|��<e�\pFH0�y�Lpa�h �'��X�%l��ݬ������۶S��L4|F�@�с�kE�x���x٠Дӟcs"� YM1���e����0���[�|�6q�����h4��e�s�u4���>x�篝�xq�	��4�D�Y�}�ϧ����t�5��\��I$���é���D����8L����_�@�>(����)jn�e���
�qR����8탣x�[��B�R@�l�SN��2u�UD�d��iA�n��I����$M��.B�M=l)�I��������\<d�6�c�A��m��&8��LF�tzI~4�64@�����6l�;>�V��Q2h�gN�, M4�:'���(�oW$!DPB)�Q�DR�<�)���s��8D.\)("挼�A�-��Y�e%EC�<Eϕ^Fr2�Q'�l~�L���iq�hh�N�6]m&�F5�U����O|�I!3��_O�ѯƜ���!F��.L�þl��s��h�w����x"k���.�?H�$9x1�q�`��͎4h����l�V=&B�q�ӧM�I�q0���^��m����~�y��G�yÌ*E�r<�J9}���.�N�a9�BJ��\�_c�CjA�rmˆ�(&L�xi�ɈE�%Cy���R����61��Oq���l000X�'�IYq?>G�E4x���2l:q\|��;t�<|�bu*گqxܒIc���p�h��g%�
��8�Ac��UCㄜm�C�>x4�
�3�^���#A"�����?"~�0���~!�.H���3��:t@��QG��ZTZ�*��*K!D�����$�Ǐ���D,>�4̏�r�j�բ�*s'��M���-��l�Ǔ-�a�t��o�>q��O, M4�:'���'�@�D�ǿ��1�t�I$���/RDr�~��0m�TQS���, C��܍�zQA����LT��[��$����=�XA���K�u}�!)[U�_eʈ��F�	nf�Ҟq�g�a��N���`�ʽ���}X|ӗ�;fO�7
�&����T��8r6<����!���%N.�e���T
$�S�i�����Nθ��~z�����n�qi�8h�<&�i���c�DD��ej���]�߶�mS�Y=x$<�˳HY���y��.��]��2l�V�,�ߋ��fn�i�`�WfK�b��2��b�G����2I�D�EϰzK!P�c�˞��
X�~1������>~<I��NL%V��H|Ǵl���$�S!�i� a��\M��6�i�!�B&h����6�h�%}Ϩ��<t�4����$	��4�����O�T��y1�d+)B�!��8ǃ��sj�p�&�zV����Kȶ�!�� ���)�Z&�c��Zd�n#�I�[*r$���Y 竖=+��I!��#�SJDQQB$���p�bZs[�p|�LC_Ӥ䝉���_Y�Q����Nr�#Y��Sl��n���fp��$_���b�{��G��؇��ݸ( ����O~zӰ��nD@@ya��+�ȯ�3�n��_�ٜ�&��ém�<�;ڔ>�����ޝg�800�>�>�$C`|u�#�	�����$�Jz[E��hv��!��1�W�ӯ��	5��:x�"�-��k��c��F+�8%���e>bP`s��9C�Ǌ-�*����I:x�,�a��, M4�>8p��t�sWYTq3�-�]r)�&��ŔF�wVE2k�I$ G�6=i��X�~�Z6l�6�i�Ax��/�7��W�~;12x�ȱON�I�?v��b����c�ѣ�ePp���<��v,:~)�6Q�x�X�ٕ�"�.Q��ù$�Ȟh;�&qnaA�)��}��р��v�`ㄱ��}_a��Ǐ"a��, Dӆ�4N�K4]7��5\��ì%�)C�����dl�~���>�b��t��~8nx��#'ﰖ�r�$�HJ���T�>
!aÓqӳ;��>MY�C�h�*�¦�������gȀ\�4:vL�@�Y�8u����F�OVX:py��a��G��V��~�����J�K�r��f1�]�۱��fN쓡�a'^��ҋ;�8�u�Q���N������h��>?�:X"@��p�:xM,�"�C��FF�~�A,t��I$���jR��IE�C�6��ÃF��?��aC���N!`�iA�}JK��	Wa�a�f�cF��Z��ㄟ��#�p|�4�/�;0����A�K԰�,�+��O�R {O2m�n�4�:��"�Ӂ��a��Ȕ<Iu'�>��ه��6�Y��#�[_Όt������8҇�п����|�Y�JӦ�Iⴲt�#�'b
H4�(�I&���1��Y:xϞ3���6��������������'�$t�#J8W�hi:I:i<4�:iPi:i&�iZ3F�I�G�g�B���G��jX�Z�c���A��$�D�Se���i���ii=6bɓI�f>�`���iٙ�Zt�Z{j'O�?	?��F�1��W��)Y�&�fLi"F��&�x�+rx�H�7<v���4L���'Hb4�TGM6�L �4�#HH�<�*�g�}�/�������1q�H6b �v"$�i�j#N�����,摆�Ri)�V�$i���#$���Ng����♧Zr�Fl�*Ȋ Y���7M�2"CHB�c�C7r �B�c)�(���Ae�BFB&P�!Ac �iDZI3n=4�c!2e!DS�e[iD6,�������e��R�Cϐ����D�d)���p��6�q�6�;s���8���3��ѱkq8�#�鋽&�莑}s����.���T��N���'�u.��4.dۨӮdx��=���|Ξ�w]��g&��hw�)��ҝ�E9�L�#=�}Np��>l��P�2BqҗD�:5�4r1�d>?�����~3��yqשBͽ���W΃<� J�r�����|��{�u����h��bq�݅��c�Â���������ɼ�r}d�ok�=�w�N{��k�g�}�.��?*�icjTJkJ�o�m�h�Be˱t�qV&���ץ���7T�qR�JU��k\��C��h��}l[�m#�
W[+����a���-���=����d�6XғV'��XT��ؘ�j���9�\�C�c��B�׶�i�:o�S��"+���	�U������333��ʪ�^�ff��꫙{�����J�fnffn�H4��K0K:X"@��?�|i�������Ώ>e&m�e��fl�HZR�%�ƅZk*v����������%!r�d�(��d)!R�&hba&\��IKh��4�`c�����h�&�ɮ����ًHUFB)2��V��f��%c״�alx�TN{m>��Mj�v�� ��[�Yb��maz���1Ilvv���|D��K.�g"��V��.�S[h�r�c��X�M�x�I!��}����ɥ<�"�Bw�~Zt�ID����P��[����dǩ��^W{&�����}�Sدs��/}G#�9��
�t6�d,n���>ӷ{��Ńn�Q@�3>���:/N��O]M����f��l�a��	7�'I���
䁽Ҧ\���z�1����������ǋ��)a���kv���sx��&?�2����u��ݬ�%�v�� ��xHZ�ReA�Ϻw�}t�u��x� a��64:��eO�U����<|`����a����$��p�<xM,�]�n�TK��ԒI\p�>4�P��XIL� P�dԕ�>_ۿf��f�I���D�x`��tv�ci�g��h2�1K[m�,li�J`���C�ŴX�L?��X��p���EZ�c�+q��C�<�c���C�OIe�֎�#�C�GO����h,�>!!�le� k�����G�M�(م�<'�ŝ, Dӆ�4O	�����#'G���D�Cy�I=l���@0a���x��J��42:,��Ǫ���Kt<�� �ۗcM���3�H;B�@���$�y��m�L*9WS*�b^%?B7D�&��,�C�p�)�m9��l�*��$L>5�:�F�hz|�s�`ɷ�6�|�B�c��$��9M	����$��.G��ɉ-�v"��2u��"i�	�3�	�Θ>0t����Ζ�"Q��4O	�K4c�2�+2I$ d<�y��HP�p����_�����ɑT��qV�F�%aVF�e\�*L]�%�C^dcя�tva����;����|��֪S��D���������`�����8IE˙/����Em��㡒B�cDm�u�o�G�ʪӗ>,:SC�h���K.�6G#�Lc��O4��O�[>���I�a�N��~,�`�->|������ι�����Y�+�t�)�E{�FSS�߼Ȱ�k�N��);&y^j~i��n.��	oU-Oa��`�l��^��ڜ�s�I7ߎ��Ͼ��N��S�hzpI_�}����w�?��tkQ��t�����F^�"q��uq�r���N���.���������Z:���-3��
cXh��`0�ǺBUa�.��D|�������c�m�FB0gI�D|��M:�n�{����lh�ƞ�/\���KP�#3i����XiƜF�q��d=���U�A�yD�-�TyD1cM���F�Č~�d
,>��Iک$��J�Dl4>t�y�8�Xk�IC��,��D��gKH(�N&��<l�S�}Dm���-̒Ia�ia&�95���X懑8:����@�|��<>zd$6䁚�P�2I�9�x4X}�#0��r�!�D�W�Z`��(���lm���7����p\!EJQ	T�!�������/�:bæci�������Y�ߍ'�Q̔կM�1$EAs�����LA�#��ӗ͘��aƞe��>>4L?t�D��4�xOY���<���Ȭ3.,ʈ��h
�n�~�m�Jx�'�ۚ��f=�3�Ք6���׿6�m$|�a�U*����;xY��m������3sD=�$�����=��F�L�;�����p��S��l��ж�n�V�N����'�T�ť�f���Q���$�D�� X|FA$-��g=}7�l2d���vd�f�8|p�ٓ`�%	��t������#��+�H��S�$�/g�2zpm���ϋ1����M=(�d�=!X�1<�r�{�mHZ���������,#�9<`0|]��c�LO���������K�0�:`�Z�4��h6th�¼r���Q�J#�/xrl����i�:����u<�;O�[1��44��I�cC��|Ӳ�Qt�x&'�i�<i��,�`�%	��t��'տS�(��|�)��cQ�`��)�!I��UBi]�
>SMc���M�)�M�_ӷ��&(��Dk4ɰ�bř�4��ԤΖ�J6Q�n��$�HA���)����Ht�Ic����1��t����׫�痯<�'c�w����g0c� A!�GG�=`�t�ɡ˗M|��T��ys6�~w�����S#筚wFvz��*^ꡨS��]1���4�M��OƏ�&��*m����nw|Y�l)�S$�i*H@ñ��q�m8�n�=��N��P� ����i	�hb�1��U�)��ۈ����4�mcM��욨�Khr����N�Zxb`��Y.cS���:ǉ����n>q��t�D��ӆ��:if�^��m��H��J$��n���jw9$�B	Fݍ�k���̥��\�jTÃMPX�h���˖�������d���Lq�$
BР(�������Mg�5mPe�Pi) i��r��C��^̐��c�R�dg�X���/�f~�Z�<��OfL+eB�l~-��S�E�T��oV�=罼:F'�M�o4�UJ�i�.3��4�C�t�EI��'(L�"xD�0L,�$L8&X���<t�<t��DDJ<X�iE�4҉(�CCM D�����"%��p,HH$A���j��p��c�8��ǄD�:@�"%�'���&�i�&�i�Y`�,L�bY��0:pA��BxKH��L,��L D��N$ �'�:'O	��x�,D���,���ܫ�%K��wS[��[�D���.��J�Aƻ�w~әy�{�?w�o�}Z��a��^A�i �<��)�E�<�6I;��>���楢W��'��>�/_m��I9�Dߗ?>����l]z���{��g��\�����	�L�}׺T!oy.� ����oWw���ϯw�|?{xMD}�a��V&�:���_o۫7�������Q�ݱt�ؗ�T�z�c�����J�fnffn��*��{������\�����ސi㆖h�%�, \i�;qێ�<|�ũ�uն�T��x�2Y�tQ� /��21�p�ۍ�a"`~S��8N���5�ꋳ�+GCޅm�M�Jm��9d�d|�n���{4Svc�R�\�2ޏ�hxh
x�B�����d%UJ�����8�?>zrJ�p��ƀ���`E�`e8<<��2��A�Ь�O�Ƥ7�u,��<~04�Ä7��l(,�j�h�.>��O���	��4�,��D��ӆ��:if����	�$���"�LxU��[ԒILB
#�#��������6)i�H�|e>�����R:���֛R�:�X�f��i��8$�n3>"q�>`�#c2비B��vM}��48(0�ϛ7�tY��S:���^����|��MU�e��������϶y_�f��k�4&��Tc��-<�O8'DL0�Y���%	�n>v���/��6�cLcLh�Md)$C����"���aw�ˏ�;M���h�!�)n�L�Zj�$���ʵ�2H6�6����lmY2(�6˯M�I$�����,8(w)J|BSKG�7:�crw��o��hĻ�AouM�o.����n��˽BŽcy�-p��I7=�����e�::j�
)���Co�*ɷl��G��O3	��tzJ2�<�7:ȓ��Y]�94�cN?8�YWtK!�Wa�8���M�8ѐ�6X��G�]8�|䐠�%�T:V}�)�p<|S�C�?�Զ4�</<���L�QR��h#?	� ܧ�u�e6` ��h#!֗)��>�&�:xD��ӆ��4���h�7��$"�I$�=��:߉�b@�M2bUq�uU*N��,���wZ!�v�UL�:�[�i���UHI
�xr9���@�4�}�2<f<0jy���f������nL4�ɶ+)��(��X�eu�(i���F]�����%����OM�u:�>WbТ�y��'��!��P�i<Ii����#"}c�����P�bY�?�4�������p�<q󷏜�-}3.���fX\0n�e\��$�B��A���4^�p:Ӌ�;�a�\��Ĵa�_4��g�m]]�WA�E�|M_���IT�u�O��>1����d-!X*��S��8�n����N���C�&�!�
�.;�����e�O���(�#9%TÓfY�ӓa���ITV\�.��ǂ���f����G���9
�g�0l��,��J�ƈ�ig�;l��v�5!$���gRI$ p�2�}���79�J�
��k�T}���f��[q�����GlS�?1���K�KrG ���Z;��p����tQ��$	A���v�|x�Ti烧��0�1�)���pJ��%���~����&�^:�~����`h2���ӏp�d�Rq�Ι���J8h�?tKDJ�4D�K<i&ɤ���Y�k���hE(Q���Q?�'r����YD$n��S��i�)��i�F�a��'}%R9��hv5B�m���q5s.�әn$�5V��V.���$�B�y��+ä�S��pm�c�L�Z�_�y��;߷_}�����s�ύ:!��~3��'��j@�Q�+d����S�M�LO��=���[ǆ�1���a����v��̼(�t`��/<�B����N���%}����rE�ٓ'�WW.Z3��G��y�ȡ��F�����:RFD9+��&7���\�̺���'�q���
2~��}����i&�X����gD�$N�t���N�<l����S#%�V	kc{ĒI?%�$���p\�>�Neu�g��\p�*w��ђB(�gC����|ѷ�d����v�G�5��cg�ճ��l,z::�������$�}�z5�(0�zY�ܙ|��a6���GOM��#�S�'���F	�,�M0K:%�"%	Bh�f�i�:t#`�6�&jb�]�DBB1����pJs�8����e�9h�W�������o>f[w��u�����l�|�������b�	��	B*�p��w
fcwWU�P�}�R���u�8d5���[J�s�y�vVf�N��1�O^ۍ&1�D��q��;w?v�
F�|�M>��m�sߏ��GM:t����ΉbH�BQ���������&��C���I7*��I$��s�~I��g�C�4�̹�-?�\���<|T}�!TI�ʒ�;������P�����]��tzS�Gca���ɹ,�YE�>p�:r=�9�ն<8!�&)��֘`�J������,�A����D������A�3��D�bvt<����EP���&Æ6`�� ����%���%��&$	��(�(K���#�t���"""%�"Q�I"��A��x�N�h����$�!B	��t�"@�@� IDDD�"H� AK�t���L4�M4�,�K,L	bX�%��%p��DN����Y〆	�H�p��b!=Q	B`���'��(L�,�����.�N@�}���8]�
1
!l�ꨢ81d ˈ����q���"
S�SH�(3X�h�1��R������S�TFQ>���B8"�D)�#Dt�j�b�^0b�S�!���19!�3CƔzB�Pa�����{̇C��~��|��I�$��6j�V�2����t�0�_(i��d�E���xn�-g�:P�'�[GݺE�DmHuO>8��HQ�����ˆ�1���Ga{�K�DZ&I�>�[��SPE���i�xx��1=�3yv*��\f��k4o�}�7~'4/ЛtR��p������ǟ�Ȕ���ߞr�[�ޮoz����Y̧��S_ws����f�G����N�T�݃Q}�mk<��z�Ҩ�!�3�����e������X�Du�Υ�ln�ڥ����*H�R�����ͨgɝ�K�a35����f�>���m��k���F�+u�2Z�y�zjd�j"��q>'����Yi�.j��@�p�����s�&�O�^�)�����
�,�ҳ.q!+[B���AX'��ӆ���;-����{���n���W33s37wwx���������U�̽�����M,��i��tKDJ���,��d��/�O�s�!���]�)	Q
Z:1�P�X�BA��df7�J<\�3F]!��e��:K�R	p�Qbd-Bx�F�[��d���(ٴ��F�A��B^�f��[>ebı1-^�pG�)�� ��4I1���(�1�:�TXKq��q-��Ĕ�h�Ę�5��	��&�	�W���֓ÓԳD�j�)dj�)����N.1��&v+��.WM	s M1r�g]�bc+��,c�MR�,�Q�i�iַe�  BA��œ�ʔ��t҄��=�D�x�Z!h�bɛ�����Qv��w���J���;���Ac�ia�81�X}�����6I��.(>e�{�ã!{��Gr�x�b�=zX�C#g�W�ƍ��A��H��>.M&'�d:3Bˋ2>mzfD�����Q�r&,n��ǴQ��d���q��Q��t~4u�8M;l�2Q�d8a�L?a��bH�Q�i��i���FkY~nōSE��M�m��0��u�Z������U!T\�p|2ߜ�
�I%��=�*S,��������Hd�J�[<��'�M����ٵ;NLbv�ٙ�d ��{�e���pptPcE��C���e�J$�q)�ʱb��?쉍(+��rǭ�x����#����p༳%*�L2;vPA�����9(+ޕfSq�&�ۜ��9��q�Ǐ\4��bX�&aFa��Y�zH�H�r��җ:�I!�%�?�t>�����2�<tP�e��U|(c��,��q�y�d���X~!iQ|;
��P�hR	)��9mE5��#�x�1���l�����2SM�a#6d)�
(v1�d�E�P��[�����ӓ�˙����X�:�5�t���b&X�"Q�p�L4��g��f%�H��UL@$��K��"ܬQ���Ixt��8s7.�&�hh��	�#D�!�g���(�&䐩��W�F��g�r�MHb�92@�GC�٢Oa$tƇ�e,�~C���V0�T�C~-��Bhr}��$�р�����Dr@��G�Ml��{~��g��G�x}�%�u��~�N+�ㅖYf�a����(Æa�O�O���S�#��JHZi�l�)12e ��7M4���n1��+)(�#����8j��Ѐ���d��Ҭ��u�ɮ��5.>W	��Z!�[��I$���#�����qf�=�-�ͮ-}ҥ�Ǽv�ތ\��sC��?�W��>(;L�n��/3�[0ь>&(B��U��r>ۦ�Pl�;1Nʪ�(p%��
�uЎ�.O���(Ɋl��+2���r{��Ǟ;Hx7{,(~�{9�ӌ���������Z�!2�������$�v8}Á�5m�l8p飆�?ibxD�
0ᅚif�iLr~��?'����7�1Ǧ�ϒI$ �g�֦�g]6��a�ڪ�94�<[{hr~���	��uˣ�$$���oS�:�׬�K?�;=����K-*U1t�e���z�ٓ?A�(�#቉��e�e,)u��p������c�q������ݸ,'Ėp�R��4�t.'?B�[N���c�>q����4�<"Q�p��4�K4�d?O�5�&҉�T�RI$ ����(l�eJ!a�9��t=w�o�,>��ǉ8�C�0�4��K|d�a�JYi0�dv���G��4��x���e��%�X�)�|̍�)���!��Ò���8]U�$��ψ��'�S���T��~�fβbQ���~53����?8���dJ0�Y��if�13<�����SrI$ `q�ǭ˱˞01�;�i%�i�׍�O���H|B��Y$�eB�����ܙ��3�����ab����r��Y%����.�v`��FI#��o��|:욧���^i�����!�m�0������2�0��^|�i���G.U������!S�sB�m��;~~z���:qƘQ�,�K4�O���I�	"��(G�҈8�у1�#IN������1�rK�t��8)��Y�#�;���k^�����E)ꜵ���e���E��ۛ����ӑ��%�I$�ȍ%�\"
���.|Ѽ|=��c5�J��,��"���{����>�Sg{��m$�t���HHA٧D����|�v�����Ͷ�b�4�r�[a��t�L�6=�AoF���?8h=��D$29��np��}t#�G��aa���a�45�MUh�E�D1h�w\���B�3�!sL�~d�lɇ��T}�i�,��D��:"Q�p�g�<l�G��i��u�S��I���=t�(6����w}t4��ۗ�p}M��)�`�����Y��C��R�~X�HZ@�~3p��L�U(̝B�; iѡ���p�D���D��]�]��P���zӦ��ܙ ��	�&����Y��=�V�;d��i0�FǽřB���A�-�0J�|@���5�roo^;>m��q��+���"P����%��"`�&%�̈�,K�<tN�$ DDDL0Hy�Q"'���B'DDK��p��p�_1_6��6�ٷ�W	 N�$�"""%��@� AH(J:@����DM4�D��4����,K����g	:p~HD��'D���'��<@�%�I"It�D O%�0O'�LA0K ��+��s�qQ�ϩ�~�Y�Y8x��_o�y��"p�3����]�U{���ݑ��-��V�L�WOgH�}7w�>v����<�#���k��߿M����V�����.��U^d�_;�g�D�}�����HS�_�c�����7ɷ1f}��Ttɲ�z�}P�>�<�>�\�蟗u������\�	�_q�Ͻ�3ݎOyF�������s3wwwz�ffnfn黻�s33s3wwwz�ffnfn��Ɩi��h�Y�Eƞ����>x���%��m�Tѡ�AL���v�����O�U�t�)��O�X�N4ٮ��V|�ת����;�ҹDoA�:A��LU���u#$�H�F���}"���:��(��]��t�"۷��������������v@�7Q�(��m��~|jC,2�aFƜ��>ھ㧊<xK0�4�N��aF���������{�sP�V��DF�H�5�$�(�C�����ö���Y����8���ݞ8o��c�!�G���	i�v�(��k%���]�>������,��5�2d6|���#�Hv�HIC�:a�0`!�Pㆶۇ$:>"Ɔ؞TS�1�w)Ӈƹ%��Hp4��?9p���GF��0�5N�s��i���L�u�'4d���f�(8af�Y��l�~����B"8��JR�DHR)(Ɉv��0�.~�1j"c��!��]�Q
:����nEP��P��1�B��Nú]{��7N$�H@��9����-5ޜɔ�#ə7ɐ/sQ��kU���o���-���^�Jp�\����;�J}3�_�߮�o��t�����N3nǛ4zi��C�����!��gp:������c�	�L4�M�HB���7�C�E��~��"�BD�LU2Z�nG�<����gC���Q�᷶���q��M4||xD��:"Q�p��4�K4��?l�L�6�ԄaPг��N�$��Ccx�p���v4d�D��UT�-�hpC!c���5>,�nM#,����6CcN��B�>a�O^�g�̐�:6H[��%�S�8	��HB�#�t�F�m1	1n��9�ܔǟ�#���i�|d$4�7��|4�ل���MF����g� k�q�A��I�x�4�N��aF0����<c��Kg�Ic7WWEg:�H�2O�Q,>;����J��pY�46�1�.�-�Q$~ ��N�o9ps�ɂ2٭p�a*���I�K�Qm����pa��,�*�;�OJ�WV'�n�R|z�6i�7&̐��K#
z�)64�[K&�|�k�;�T��ܫ�|xJ�4���8&Y�&�i��O?�������6��(����ICK҇����dɂ6Ø~1vϫ:@�yX��uEH�)�٣�Ƅ�Y��f��;� �F�i�C��۩\6�!��^=R���0ٲ�`8�;ϳ�(�.��|�<�!C��Y������b��W߷:�1_~j�㷋������V+������a�if�(J0ᅚif�i�~82����CSdF Tє��B4�ES��!S�,�kÐ������pp��e�!F����iP�*���$V�cd�M�bg���n�$��!�|�xvO�莒����|?�3�\���2sǺs�w�[����^������V�#yFpM�g��<f�L�?�?�|9���y�TR����>�Zh��F?ܥ���c�c��K{�f	8S�Ҫ��`v���o�2C�|�>��`�ӱ������v��U6÷ƛky۱4�|$��:�f��?��]3�!�m�t�h�w���a4`��&�"if�4J�8af�Y���QNt��Q>��I%�BG��0�@b;RGќ�vF�r��"�=�IѷA^ǠJ���
h(|������o���!�ӗ/#���~�_-}T�Q,�10�!C��[I�3̥�U ����3�̏���#]4��	R��4C�����V��r����&�^&:x�EUW~~����}�(�a�&�i�D�(Æi��Y������>��+���ѕ��=�I%�G3��e�Tk
�.0Իb��jY4��qn�ocKk/�g�j�1ݷ�i�<���.2�Ȅ6!<P�����༔ǇHah�#�I���&@�m����ΈB��sUQ��Y��$2�$�A�V�a�L7�z3&؝�+�sF�^�d��f��h��4�P�a�4��,�/ߓ�؍J+MW�$�!Ŝ?*��x�v�HCe�'�!��Q���cݰ�u�--�a��d�(-��ry�
�o�"�)�d)��n�g�N�i��L�`�8�Ւ'M&f����J!K��`UJ�l�杸S8fH2B/��M82C jS��y�vK�U��xT��r����m�N1P`hX��"P�=��<'�0DD��ı0K,�,K,��:Q �$������H�@��X�'D���'H0E8q\b�q�q󳳷J����ip�$D��J AH(J�GȞ,M0�4�ML,��
����	�҄H,���<"&x�D�	�$I N�%"@�(J:`�����`�&%�xOh���2U�J�W�'	(�����#�-�mh� z!�2�?>��#�,1ALGI�C2H}���1Q��xAc1��� _���M!
H<�(�P�"���h�3�E9��g$d @��d(F\E<�C��(wN�E!@�.�CQҔ�Z$�߹�I��7��͂��A��"��4�E\ޟi��B�VD��tx�v���c߮s�d�x�'�g�L�LA�>�ё��};J$��R��Ji�|pߦ��p��7t����������pjk�"wK���0IQ��w%;�CQ9ќ6b�Ď��Ã�'i�h�
X�DBp�QM���DHdB�8�߾�3�"ȯ�g��#�E��:�<����+�׻�5II�gy��{���G���.�C+n�Tj�WS��|�|s��n�FO���.��S ��|��LrD-���G�x���4m���j�k�B���p���!�8���`�Xz�\�MfkmQ��kFk�76[��R�+R�h����r�{du�8�n<����ƢP���ȵYj�u�2&�")[cG@iZd��jm����6��O_m��.����N]_^t�D5^'�b�Ɋ�U���˻����l����www���������������7ww{{��M,�MDM,ӆ�BQ�޼q���?�m����dc�B�&Y!B!�(�H"���6�F�K"M/f;t��PpxR�![7F�� �$�tx"��i��7E8�3Y��X̢��F��b�K#�r��s�},4K,̭�[��tS��T�HL�z�0Y%�]47I��:���bZò�n��h�C�5�y�Zʺމ-�ں٪�kI{jEKfM4��V���T�QtL�)�k��31f�[UZMqv[nn���.R-A�ִ\)������$�X�0Ҿ����1����NU�i1�7���3f.��rri�.K��6�Mv'���T�>]������!�r�y�:N�� �lS�4�4�T�����Q�U��a��>p�D�@&h���˓�Gl/0$�m���$�`���<���\?��t��d?��i5�����6�&'�����J�s�l�B��iہ�-�L�s#M��F!R�2+��I�N�gh��F1-3�sw>�M������ļ�<��ƛv�֚&�i�D�(Æ&�if�QqW��-�w[��{����;�!-ᑡ��K<�~��tÇ�#.U\��v�����������ɲ��80jB9xr>�����M��ۜ-nrxnjv�1U�h����<�LE� �b2���#��_줟pX�Jit�B��ȣ���FWFJ*������Ja��64�3�8�#�(�����gO�'�<x�M4�4�N%	F0�4x�Ƭ�T���vэI$�!���׭�����MR����p�ތ����N;h6C�����̆nF�����<`�d�ʚ)�B��T�b0:g�"d�LC�r~X�c8!��1��!!\S�}ta�1��(�-��p��d���49t�T��(��K4D�8h�%p������8t�m�%��O]��By�Uk�I#xaftz84C�Щî/Ssט���j�>b�X�j-��V�ͱ�UE�ji�����!G�d�]�:�h�F�!N,�+���[W�̞�:�ڿ&��'M~w/kk{n}:�UI�4�W��ҹU�-�ݞ���}��j��FǄ6p��g�:x����%a���iӲ%Ç�A' �|i
Q1e4`�(�B:�B���g�78�pl� �2��\�h*,e!��IN�ox��g�0Mn��!���c��;%��r�n�H��$�!��1�MC�����&%�΋�ӝ�5	>��sϱ:�y}����x�=gz�|��Fp��K�� �G#��WW�dp;ke��|qz�xC���[��	!�����ia��W�=rnN�Xxtt��0fH�|h�*U��l��z`��ӱ��ۣ8:r�܏���tC�?�Ǐ' �&w(��6~,����cx�'��4l����4J�0�bx�K4~�G+2��p��@ ����{O6q�}M��(��w�OMwɶ��*��5+�q�N��ګM��M�XB���*o!
#���""�� t�,��j�j"5
k��!g3��<8#�b@�Y�M~����	�d3��S��K�pD`��Q�y��C��L��fM�<i��&�i�D�(��'�4�Mx�vm��ll�Kҽ�Q}�$jH(�{�@��8h��LP)�ߣΆ��t ��єO�!�%V#��!�)Ե# �h||1	����A������UJ1��GŎ8|l>㰄�F��'�r��zn�&�gF*�i�Ǝ�*�Q�[�h�8#�b�����0�*LCǞ;py�N6h�ӇM0ӆ�BQ�,Oif��"#�㗱�NE�I:k�6����o]2ӆ_5��[���`�o�d���P�d��N��Wmě�n ���E�-?;�MC���4>۷�:v���`���,����%�!��d�nܦ��m��L�bm��>ވ��L<�p�i��F'�3���~t8o�Q�lٳƟ���?i�M(J0å��M,�����f�!
2e�1?"f���.1�/ۜ:�q�F��D��.�
s4��]��ޚ�f�si�Z���.��H�6�;�V�vE�����*iqK �lz�q�w��u���$�!��G�)�������~9&�8$����+�ͯ��Ǿ�q/�ǧD�t\��y[�z��.��פo��ܕ�]�u�>6t�8c�D��2�D�����C����C��TQ��|�:���{46�B<S&)�C��1�'k%<i�K�D��^��9�t<��㧡	w.�`�6�Iold;Վ!NG�J#�,�c������7[E}��� Cj���7:g�ʞ=�9��OU�Uc&��ò�;��i�Ξ���4ᦔ%a�Κ<x��\!%ƓrIF5$�0����GO�!d:�m�O2V�������ӇJS$-ĒL:�rx陔�j�������oڛi��*u���:h(��lh�ǚ$4p:�!����{(�Q�[r.���#q�Uwm�x��u�ڨ~¯����w�_͋`�@|��L�,�2l�UR_H̏�;K�e��m�6ۍ?1_�~8�cq�X��	�,L�L L,K�3�%��<'N	�5����DI$J$�䄑0H8`��"X� A>D� �DN�;;;v����ھ>�.��q�""&	��@��"P�'D��"a�4M4�L4K4�J0�0�0L0�,L,�:t��H<pD釄D����@ � I H A"@�(D��,O%��&��Y��p�].�*��}�2}�V����Q����s�8�={5�="���^O
�W��g�+�.�I���}��O��_ON����	���2������5$��r�{�\�����k���6�m��_w�=ݫ�Vq.%��\,��*��,�̚ƵY7�%ޜ�r�|����w��Equ4s�����W9��>�'9��Tt��:^7�7��Y~{Ng8D��<;����r2�{�F^�����wwwwv����wwwwwn����wwwwv����ww��Y�&��a�,�g6t����&���fI$a�x(�%aw�A�F�٣��3��W�M=[��n���P��*�^�,6B�1��!Ҹ|Y��V�-�U+j��0cm6���\a��CÓ"�|�0xd�l*�49!�E�i���D:�LQZ4�3E01���K�Qr�r�Zm)�n��!�R�K�O�!���~��|t�M<i��K4ҍ4�(��'�<l���gxU��rI#X����dl>6�;\昴7�[��������b8!V�����*����.�5��fj�G�+Սzmo%ʕѽ�!�;r�RX`��D61٣��m�hlx���Z�ДUI[i�4�Uz�0�!�����6�!iM����fBI�z>泭N8$�h�Cea�П�p��4�L4�M(�J�0�;|����t���c���oOU�����BE(�A��̣�(4���sY�QB�ɏ�F�1��2$�;�,��J�eB*iѶU�ucA��H�u��2!H|�Ib%�<y11	|Δ��ɟ�1�j��Aw4��P�Ÿ����.����>ѿ��Ɯ.(Q7m�<�b�C��Q�f6`c���j1cj��ro잛5:1��Z��!�F]�$����`���v���O��/8xCm���#̻���=hxC��f��j�e�{x�a�"J5$�l|��C,����cjn�Yu��6�f����v�J"�)xC�6��r��0hك'��`�i�iBQ�0Oif��Wi(�y��R��q$��#�m��d#>�A�5L��``q�$חU����K�X���O��2,�$�$\=�cƌ��F������!�Rt��!<79%W%и�°	��M=z�N���Ne}�B
#��~88Q9ݍ��0�ZC����
�ك�M,�L4�M(�J4�:`�4�������$�X�{9���ԑ$�;\<:<���C2
j�ې�{�n�l�U�y��M6"i��),�是�F&~�|m��+�{)W�Q��f+�1KH����%����l���������8�t;4�a=(�Zr�d(|4���9F�e�:��zlm6B�b�hܔd�NX��L��{ơ	TW�d��]���i4`26��d��4x��M(�J4�:`�4��ȕ�`�I��$H�����$�!tI]�={lǉ�i��+�m<c(Ү�~��g����nlqiF	����= �!��.�>�(�
��hߩ�S�Kq>�����\h��7r�u��1pCnY<�c�)ɡ��W�B����&���ӥ�Q�.�>`蠐�m�:����+�k5��:�x�4��Y��iF�Q�a��?�?��4DG�R�c?�FB��(�U�L�bN<cn	�t*ơ��m�[�B6O-p�Yp�#�j��)6A�n�6��I%�C:�x�A��Ÿ�x�f�&:&��i٣s�&�T+���8p���>���;��x�~��h��RϾ����;s���b�qA<��ӥ!�|1/�7�B��Uw.�I�2o�%J2�=%/�g!��q���x����,(2C�4G�Ql���D��A$6�іh,41�/����A�)�.���(JISn�$����V ���6��K6iۑ���<p���,�J4ҍ(��i�M,�����Jy�\%�9��@5���ݒaiz`�DzB����j�I�۱��8
�.txћ��!��������2>L��i���GA~~�iN�h] ���!��'2�k(���e�%܁��c3�AG�>(9��i���i��88���<TĐ}㦔x�4�M(�J4���<h��g�ˢNZ��1��D�LAd�+R�u$�XH���[~<��|g�?�$�v:�lp?f���O��$l�
2%�NΞ6��ɣ֟0�T��+����N�G�Q!	`�Y%��n��Ó�r�����rBd���_9#���|@���>x���}�(�����j�>vFlf���a�X�i�iF�&0��i��Mt�ugJ�Q#����B��`x���2��$�1�h#C�iƭ��}�gM��v�֛ck�2���ȵY��ƍ�,t�'����t�aK�U�#����eQ:�9Gxӿ����f���$��*����I�4ĠٖG8��|�B����¥e��u�4?� ��W�E�4|��
�����!������O�J��������%�4ѺQPS$�&Ff����6[x]D�$ƃz�`IK)�5)�%)JR���)R�S)eE4��ef���K))JiK*+,�����VSJYZR��SJjSYK)���%2�)e*R�T�)R�)R����Җ�e6�Ԭ�K)eMJYM)�M�5+6��4���M�*SR�)��JVRҔ��ȥ%,R%�T2�R�m)R����JY*RQJ��Rȥ6��)����SR��jSR�R�5)��������ԥJVSJjR��V[)R��ҖQ%(��XR�K
QJԦ��jL��%��Y%ۛ\�MI�$�KK&��i,�Y*M%-*K$�M&M%�M-$�6�K)%�&V�2Y6K&ɒ�̕���Id�d�e��,�K)d�ee�RYL�&��VM-5&J��d�RZMKKId�ԖJKI��J��jMI&�dԒT�-,�Jɔ��,���\��&�l�MIIi*J��%I�Y$�2jK%�SRY,���dԔ�K--%%dԙ6L��ɲ�%�d�,���Y2jZd�L�L�M�ɲYiY*MIY,�+&�d�iY5&��jM�RRjMKK%d�l�KI�5%��Jɲ�L�K%��-,�L�I$�i*Zm&�RIRm%&��)]-����d�5%��5&�m��&��K%&�jMI��KJ��jJ��VJ��l���&��M��[&���Me���+%��5&�Y6���i)6�RT��ɩ+&��ɩ,���RT����i�,�&�Y6M��m%-,��&ɓI�T��ii��%�jM�ԛId�MJ�۷VܛI�6�RT�ɩ5Ie��m%d�KII���&��&�i4�%&�i*J��%���J�RVM%�jZi5(�e�u�U̙[)Vd��eY*�T�JM(b�**%�L���Բ�J�e�J�J�Q2(���*%JIel��Ke���ԥ���Vܲ�Kl��d��VJ�)KY+fZ�m�mq,���e���R��-KX�R�o1�mL]Q�4R�KJe6SJR���s)e6S)��R�e2�\U�+�+���YR�l��t��S)e2�J�Ԧ�aJ)�2��(�K)dR��)QL��*���jSiM)��)f�Z唩IK)e*RRқJi\�rʙK*YK)�M)���RSiK)JZSiM)YIY�M���K)e2���jk9͸���R�YK)JYMJe6VR���l��2�)���Vl�SR�Se2�MJe6��K)�JSR����SR�VjSR���2�S)e6R��)e5���e2���m)�����2�SR��T�ҕ)��R����SJT�R��R��iM���Ku5r�R��jR��)��0T��R�S5��FҖR�L���R��6Ve)L�e%%,��YY�*R�4�ҕ)��JZSYYe5�����m)�MJYMJ�)ZS)%,)e(�JX)aIB�R�T���jSe,�Ҳ�YK)�Ԧ�4�����Se,��,��T��T���)�*SJm)���ҙJ��J���)�,����R�tڹ�,�)�L���YIMJ�e2�SJYL�eSe4��ҖS)R��Ve-)�,�R�J)�,�ԥJiK*)�M�QM*YQJ���4���R�iK)�5)�,���S)e%,���%2�VYIL�ۖܥ�ҖS)e4���R�iK)R��QJkXk�&E�QR���R�JQJ����Ԭ�[)iJ���SR�SR���)R�)���ԦSe2�J͔�VR�YJ��,�)R�e6�YJR�l��4��5+)K)��Se5)e)K)�Ve5)�K)e,�e5)��VYJR�6SR�SR���MJ�)�M)�M�b�����cu�K)J�Ԧ��SR�����E(�JQK
�SiJ����M��l�Se5+6Se2�)�����*SefRқ)��K)JYKJee���iL�R�iJSJ�))��YMJR�����)b��)E,)E,)E%JQJ��P�,�+,�)e)K(JYJR�T���jQR�il����jVl���JSJYMJYK)��Se)L�e)JS)�,�����S)�L�))ed�SR�S)JJYIK+2�SJl�����SR�e6RS)���JRVe%*S)R�R�e)M+,��)M)e2���ԦVYKe2��JYL�)�,��e*SJYL�)��K(Y���(�
6�Қ������5��M)�KJT���e6���[)�Me-��MJT���VZSiM�*SiMJl��M�*V[
)aJRĥ�J)dQZSYY��J[)��T��J����YK)e2�SJVSJYY�,��L��2�)����YL���YL�����3$S��1�O��2~X�|д�����_�?����H���  !$���>�~I���¿�5�Ú�=��~����SJ�~�!g��������r�DW�������8�`g�?`���wY��?�?���?O�G�~��|9����=0~M:�mk�������kI�%������`x��E�O����?����@����	�� �,rI��P�A���EX��J�?�ԏ��?��'�?�����u*�.ⶁ�Q���"�O����?��f0���a�*'�6�QF�����D� �2��K� ��Y�S��E+�g���>	EH���)ީ��II�T���@���߭p�w�)���~_�~�)���$d�����!�����dX@%n�tI�I���"~�QG�QP*��G�D����Hy6u��Lb`���ڂ"��G`5���?����?�NA�/�DW�����?A��C��@���I;R�U$�aK(�&RL�c		%�R ��+,����a�+�����W��7�Q����������p`������6�`QI��|d�?�	Ԃ"�����v����DQEO�46�����46������ � ���������w�|�~�?���������4��SC�"@?�$��`?��+�C���4��g���?�QG���������������t��oG������p�ժ AQ�2�J����G���_�9���)��J/�X����p���.��4?�`����ҔӔk�$H�'���Ȱ
[���HRX���c�	�N��б�x�262��'����x�`�EQ_)�9���#q0Z?�v�G��By���	�ꨢ�h��!$����	�}�W� �(�G��I����?�8��_ͺ�������?��������c��~���R�������O�?�O�hO�?�?���?��H�_ܖ��E�?�?�?��GÀQE̡�)�j@���������(؍c��,X��(���TF��1�E��F�"*(�F�#EEQDh�#E����4Q4Q"��(���4E�#DQh�Dh�4h�#E������DF���"�آ6"�؍��F��آ"4DF�#DX�b"�Q�E"(�E�(�h�"Ɗ1F��1����1llh��664Q�4lllF(����1EcF�"#�����Dh��DDTDTDh��4Q"��h���b5��Q����DF�E��EDF"�6(�Dh��F�Q���cDF���"4Dh��Dh�F#Dh��F���F�"1"#�"�"4DF"#�"(�"#DDb"1�"�DF���DF"#DDh���DF""4DF�Q������+Z55�1�F�����Q�"1Db�"�(�1F1�"1Db�#DF,E�#Q�#Q�(��1�QF(�1Eb#QQ�"�E�1E�(�(�(�Q����"�DDb"�DF"4Q���"1F(��F(���Db��E�(ъ"�"���(�#E���QDb��1E�(�QDb���QDQ�"�c�h�Eb�V,[�h���QDb�1DQ�"�QF,X�Db,lh��(�c1E,b�*6�Ʊ����E���Dcb1����6#h�Q�(�Q�DF4Q�,ch��,Q�E�E�E1F�1�(Ŋ1Q�"4F�E�"*(�Q�1Db���Q�b��F(��F(��b���b��F1DDb"#�#Db���b�Q�Ѣ�(��#F�DF"1F(��h�1cE�"#F�(�Q"�X�F4Q��1�#�b���Q�FƋ,E��1Eb�Q,E�b�"1DE�ň�QF"�1���E���lE�"�Dlb�-��"Ɗ�4X�cE�F����DXōhŌQ�1F1cE�Eŋ�E6#hƣhō(�E1c1F�#E�ъ�TX�ŌQ��4b�1���4h�h�TQb1(�TX�4E�F��E�"1������F"�F4Q��F,F(��F,Db1DF#(�Q�(�b��Q(��Q���1Db1Db�1E��QF(�1E��QF(�F�QF(�Q�(�b��1��DcF"1���F(�Db"1��F(�6��1�ŌE��"�QF,E��Qb�1E��F"1�1lTh�E�Q��E�Ƣ1�b1����F#*(ƈѱ�4Q�F��-�6�EF��(ƈ�#DF�#Db(��F#h�b6""4DQ�F�"#DQF�E(�"��QF�QDh�#b"��E��#DQDlQ�"#DX�Q(�DDh�(�F�Q"��DQ��#Dh�DF���6#F�6#Dh���#Dh��^����:�����C��A_�Es���_�O�?Rq�����K������!�?^�8�,v��C��V��� D���,�0���[
?�A��C	���u_����A `<d�J��g�06d-���4iQF���� �3	D�_�?��������Z�\��X�����������~B��(TI?.l�:�u�������/��_��d�" ��G�M��K*p���?���? �A�O�L!A��?�R��:��@���� ������n�IjPRF� ��]��BA��!P