BZh91AY&SY�q�)� ߀@q����� ����bD�|    ���-�Y
��ik6��6mZKa��ڴ�iTl
ii�f��H�`�Z� �hQ �ְ3k3m���M�٪l�4�U��T.جi������35�3aY� 5�h�VMD�f�[ZZ�Rڲ�f �M�dL���ز�d`Hj�f���mM�2i���Km��lɵ[3Ej�6iF�m66��m�L��Fl�ʆf�ʍk�d����
���&Q6fBٚ�6���DA�Vڪ-�CV�TͥչwFZ��4���   �'Ʒ��k�Q]w:4���eN�j�Z�NƊ���ܬuل����î�:n�t-���6t�u�]ڎ���Я���d�($-i��@�i�mm��  ���  ��l]9��� N  d� T���p �@tp PGL ����  u�� :�u=MYV���Ռ��m���  �yA@ ��8 �ڹ���B�� o`z�}� ����}��  ���u�P ��^�tQ�=8����������y�Cmm��kM6�le!CM�  ���� �M��}� ������} ϯ=�( �p@�x��( M�{�� ���| ���p N�p��}�ꌍ4M�dT���,�� wo�����  w���Ѡ�N\  ���� :��  �/8�J�L ��P�6�:�  {�zfh��U�m6�1���4� ۷Δ ne�b@ �V� :����  st h�:$tĶ�t����tk�ݶ�� tgC@ }�{ZU�m3Z��X٥��  n��C] ���5w�@4�����t  �� a� ��:�u  9�q� :����cF�4�Z�m��i"ٕ�   6� j�+�� n�.Pn�� nW �P $� �� ���  NLP >�xR����kJ��
֫J��    �� (=�N  �Q���� Gn�A��]�w@���� WwQ�4j��  ��=L�6�X�(6V��   > ��w Ar@FL(U0` +������8 @�Zݰࢁ�����   ��B�*R�#   �� ��ъR�� 0�h�  4���1	J��� �L�� �~%*� d    R4Dh�hM'�'�'��OD�L�	I�THҞʞj50�H C�ڍ:�u��ܵ���~�ڬּ5������n���Y���;(R�Mxy�RI$��H` ? DW����fUUE �	�_��>?��|�5UTV�j��� ^�|��a@DW�����z �C���0���=0��"~�)�0��2�X��T�(��:�el!����!��(u�:��C���P�|�'YC���C��X�	��u�:ȝeO�D�+0��:�`N�'YC�	�P�(u�:�d�G�)�� ��z�Y^�X��!�� u�:ȝ`N��YC�	�S��*u�:���ez���:�ez�=`>�@G�@��0���� ��(���(#�G���� X 	�A�*�US�*�X�(=`PzȈ|0��EG��YA@��=d zʪu�� ��@G� d�"Y^�*�U� ��AP�dTzȢ��:�(�����E ���_�EW0�Y �(/XT� ����E�( u�:�"u��!��d�XN2��:�a��XC�!�@�a�'Y�`z�aN�'Y���P�(|��XC��e�u�zʝd��YS���S�/XS0'YS�)�@�u�:�<����}|�c������e���&�$Jfh��eH/v����JYz2��Kd�4Uͬ�967)�ʓ�\[��R���ؔQV6������O�DʃJ������[�L6�1A���ȫ̕��8"�"-�*ޡt���W��Z�L]g"=.iך͒&�'4ս�E��6����*�K7VN��d:QR�N]�f�'Yxn�4%��e�ۘ3u�u�5�"-�6����� �F�Z�oJ(W;�uh�jwG�V�x&A���R�	�1;�Q-�,-T��$i�m��Z��n�b�0�-"o*jd�I�E�˕�G�h	x!جnZ*������ٵ� k���w4( ��V�,�Z�q��Z��X��-o_M��)u5܎>u>@�_�C�n��7�Y�{D������,�V�R�ڭ�e��h����Y�-e��2�N��1E���shXX�/�eIFZ��08B=�s�e�U�����hT�а�{�T1a�U�{+'8ȬĖ�9P�ذ�D336R?m����m��m+hJ��M
K`M��yn���"�w�-j�RIlV����܂��$ʃ\�7�&@���ͽ��n�T2��947t:�n��Pb���i�4���4(iͭ�q�������q��������;\9����ODE-����x��(�nm����Ty��eeAx����ӫa�&����q�m�
��&���ZV���+Q��v�r�,a:�,M�vJp�ʴJ�P��pfQ�$Ǒd�N1f�(�Nj0Q�4�R��j�3] 4��KHݣٹ+72�B�,�M,l�@�y�T��enB�Sstr�*ԇǭ��-��\���es[��:��X�,t-l�s �+W��C�ی<��H��Ԙ��;;S1Vk���
{�2�3��A�6�T��e�t�����x�B\!��k��tGY�Cj1y�aTv��3���<�1�UȢ��	�AI��wX2�ow.Ag!1<�F��+&��9�'��dt6S�m�Z��$�Ȳ�ɛ�������&�-����n��:��+D��W��eZ�x�f-�(b���l-�$ U��*��+�Ҽ)8�T׻j�2���B��r�إk)ڬ�H�V:�/n�E��v�o�0�B���0���b��sey�����'V���9�q��Ļ�
��=l7�v^(\	�"�$�.|��f��b��b�dv�{�}���T�ԃ6�ւ�]�+�����,�T�2��m	�W��o*�+�ި0�P�ǉ��B,�/`Jf]�W18��+鄖�KE詷�/V�X+�̪ǔ��NↃ�u�
��0����Z띯��#)����N�)ieA�,PLx��3(�� ��'��`U��m�T�NP���orım�dL*<2�֮4Lg����(Va}�,�I�Uy���i��B6���H3����r6c�fMo*�4��R�V��)��]�I���s\���DxUe9qAWVnf��/��l/CW�^�(����j��Y��*��C�W��8%ifl[����)�hfM�IlJ�?�-���3lCn�+��n�!lʷ�O6���X�m�ER�� P���on�׮�n�{7t����"l�cz�� E�`h�)��}��wM}�1ٔ([yc�SA�Z��m�8-9>[l�'�U�US�����Sr��\�E���,,Rjy�T���-����(�oҐ��7F�ALVh�����L�S�,ǶkbJC&<��KF}ni�w@fEm!����[�Z��n�˖�ܑ��!q�����v��i�&�D젆�5P	ݛx�w+�tb��Lj�(�~BѲf1�V�8O0�9��]-�u[�Z��w�)dkZ���uv���R�u]!"�[+r�n!&9BXU�`Ċok[��e��LJ��B0U�ۙPZBU�jYSFhX��I�DgWr]���ۤ��G�Z���t��ʶ���h	Q9Gr^Ac�e�����t�a��¯n��XE�h%�*�uPU!>��A�l��+q���&�[�M��܇0��z2e�� ��5��z�?]
��u3[�0YƢҐ��H|�a�Rʲ]�1ٗyZ�����](N�	�o(�ɦ��-޺�"�`���E6۳��) �7K��9m,n�k&cٗtM�\KŸ�M��Wd�7V�-� �=<Q�tݰA���+e�i�i�O2��ˢ�q�dKZF�Q�"�S(@�ב��U��y���Rg\ʛk!��)���QO�+c�էQ�d=�8n���� ��IۗJ��Z�M��z��l�+�k �X(�� �Jƅ٫)���>"��t�}�[�$��[�sb[+p^fb�3sB7=�aA�Lׯ���̇MM�F6ђR�P�f�^�W���"Sȵ��ڨ�F�`K�5D�eʦ�ݥ��,�ȿ,�7�#n���2�*��Hk�v��1j��xRr�ra���|�b�ȉ��(�KI��;U:5���Pf�����vͳoP��f�+s#��L*MÖ�Q2!U4fA��1yzx�SmGz��.P�B���'�>
��,��hkEև��p6%�������7��")cp��5:�MeeH�ac�T-�m�7ie�x�G�r'xXp�ʬ-ˍJݼ��D���&������,�ıx������3w.^�u�d�\����ě{z2,��̡�V{�	L�m�����0!�}��Չ�I�>��]��>�{N�n�,k�K�J��Y�K8�J=��6��N3	��P��'.���H�hu��J���� cb;q=���EYa*>6��hd����&���^]����-9��l�28nm�r8�=�1સ��LT���wX�hX��F�ă1� ���w{w�Ɏk˹w[�S��}�.�ߞ���C������}�̊@�\�Km= MV� �z�,�+n��b3��«����7��ϱ��rf�Z��/p++6�1F�Q�]�4���]%2-��=_=��;%�A��t��ś�e�W
̀�3>M,�XZ��7V�.�U�n3�r�e��m����Y�O�j�>��  �j�2��!rRMÇF��O2tn�D?v�&�@���&X;B��N�-nq�ʽm��fh�+ߡ*Y����2��-��WS�3Z�m�Y�M��@.0��oIط�˹�9.��Nfl�Qc/��Y��u|p��j�pO�Ou�GQG&�qiC~Н^ VRKCn�w-a�*�g�W�zE���)!�rAh��&[�J��A�ɇe��
���pĬ�� ݑC��ʚ��.�]���a �x�dbRZ+fpC�Wj�`�ǆ-[""�'L���6����^��%eV�����.]k9���Y� G�y�,����l鹗y$Ź�`nP�ܦK2�k(���K��n�HAv�;R�{�©�KP�C�YB�
�u���`�Pݽ)�E�v
���^j#u�E�.���mZTo@0Ql�1L�36�Y�2�Kq���'�w.�.�D���� �h|��!��W�б�3�y��ʎ�T����K �r�k����ES�<�o3oj��
P�r�b����\� ��C�a��Yj���l�r��,�QBɭ�U�fC���6S�+�7P�g�j7/���ـ�R+���,6�n=^<X��SM	�O�{Q�e*�\n<��0����������Vff�,;������f��4�9��xrT�Z��,��n�˓-�8�E�CP˨�,ڴ��h`
�R�5��Ӫ=�2c��.��JT�5����;ט���a�gp�u�m�Q	h
��P���9�T�{���K��d�M�bm����C�U)�st��eV:%��Yڍ�r�z��ej7�ǲ����e��O4��3#��b��6.[,a�p9	@Ą�/0��A�{��j�0$��e^����9Q�����!z��
�w���-�4���7Kx*]k�3)�	�+R�)*��`Q�;���LAX�U��e�7I��zK:�w[X�7��m��>zl�Ÿ/�J�ZR;��ݡ�d6��Չ`nl�E��4"����XfS9���b�F��g��4fP�M�����p܅�e$�Ѥ[���#n�ul�m �fj$�D�փB�8jƊ�aɵ2UX�Mc7��d;�5����݅����	�\��AQQF���U�4h�M��X�����˃Y����qk�B�<��)2Z�d:����z+1,qm!)3	G�Y�w��Yd9��sM�y��`-Տa-�E�D�EȖbBEic9��+6&�Z%*Z��XF��,�"�7 �Aj��F��E`���շ�u�:��PԻ�`�/�r�����3��3xP�O.#�墁�W�ܘ�Ze�2e�zS�7����6�(K;V���a8P��L�Ǒ|���b�˘��J�*m1��S.\Bڌe8ޱ�,QX[B�̩	!�Q����de����Eeج��G7E�����*���٬[�:�P�)cgmT�`�"j��J�aZ��س5�[��OqKϢ� ��B�S�DXP��"K�Rb��^[{���� S#-B�,e+N����UZ�:5ն�C���1��֌y�[ݥ�6��5����FЁC�қ&��7un��N������F���u�,[	�[�2�n�EZRn�&�U6n�6�^�(k� G7q<%�O��7�%T�Y�՟� u���)��v&	�XE��nEKF$��H���ͥM�b)]���m���aSjb�d�{z���*eIL[44������gމqb�y�m�[��a�ɍ2I��SU3L��J�ۍ�ML�C��p�Y����[�dGe1�����K�i�7KXh��	I��&�T��M�NK��3I�b\�U༱R�(-I��,6f����n���WO��w��q�2fDuP��֭��ő��*=�WM n�%[:)Rfƽ�fX�,J�j��*��u��֕�v�%�k�\q��Z6�'�텔GZ48*	��NQ��� ��8�[WI��v;�ʦ8��y� 4U{W��pm� �un��G[FC�^�Ȗ�"���5GJ�{@��	Rʒ�a�ɨ�B�����ȍ��˘n�M�o7��f3�0�U�
�ڨmSÄ��v������:
j���j���FL���
����YH Ai�wF
7lL�ƖX&�k��v#:��f^P;KQ�2���`�.V�tRto+,�llYMǦ-k)�8���f9Si�n@u�9E	[wH�10nfm�)����z��)ހH�E5\��56Õ��G4j��z�k=��Pn��f�_q\�nd�bZ�g i�Z��Uu5EaX-���L�
#V���	������Xj����3sv�F�H1*%��1�%�v�L����I像���m���ô��Wӛ[C"��|wX�|�X`]}�D�@�73,"�xvdA�ۼse���f��g���i>���%��q�۝A2��Yf���ػܟOr�[��ҷ"�Ê ��n�	��X�B���%��:�/n��r͐t�<v���%����-�[,1��	�[Z�5݉;C�ud,z��Eq�tPxޮ�/+M�w2�U�R9ܸ��E�1��Yh�� ��V�yt'�iS�tDB=�{o�
�ج9����@��뭡�9Z�������A[������t�i��{΍k�1�)0����^;XBS{�c�ZI�5+���k�ylK�7�kv��YSK����ɱ%kB�q0�B�Y-����h!�0���ɥ����7�+t(��d������l-\�V�/�T��,30ɄI��)�8b�f�ߎo��7���%�t���#�!-�-�E�m�+
.��łw0Y�Y��XhТ�l��d�/1V��p)�V��S��aG�7e�̸��� Qn��`�H%��v�áj��Mؗ����w���C+1��^�ֱ}{�-;�9��e+D��DB��E�j�u�#��OWҳ`��RIL���pX6�Y�,�����B����d�mX�A)�ōL%�5�S[)d͘bÀ흦L�,)���X2�l2�w��~V�#}\�E;�k�iX�}H���Tv
q�A����2�!Dkr1v�t�/pX�F�4%A�}dx'��.�/1��,�wI�zq��yH�{KN��fWؓdx�����/vC��6�y7�P܋R�4�w�Z�m�p\�.�'v���,n�S/�^#sk,�b�iZv
���"Qm�q۬��h`��@9HV��1m��0]�$�ǉ��;q��5�WB�Y�+Օ��b�X��l�����^عV.��"���/K8�;��Պkx�S��b��,5u���LT��e�Md�28�VQפ/��\��N�Sz7��y���z�^r}��?�YB�e3a��ml+Z,X�֬7P�iV��N0�66d�ei�l�Z�,�-Hi���y�:���k�"�/���]G��{pS�s�4VՔ��Z[�h�*����C2e=��TF��iiP�!*��5�YTa�!��T.a-Xݷ���*�ƴR����JV�sq��,�R��w3�m�o(1��'�<ˬ��ky��O!�l>�Vv�hұ�ɺ��MHU]�n��Q�
.^��55��d��"���f״���q.9�g W����X!Dg*˕��{�mՃH��{9ubB����I��M�p%0[6�:��g��wNYSa��@β�)PaX!�q�qAoYS�k<� j/Qi	�70�Zj�-��5ݔ�0:zͺQ������Q9�����z��lR��y%��oMZ��]HH���-�6�g�oh��+E����fH�^�Ǩ�å�6z�lޔ�y\l<J�������;��芜>369ռ�	K!�^Z��g:�sx��#3�]�U�p��K��y��T��U����j����5����A�)ƛ
%��y�3n�Q���IB'��&YJ�S�+�dEslv����Ί���6S�q�m�j��ڍd{�7�U�-���Ry(U{2v��\�r�U5�R�����ͥ���0�R,v�yB�v���(Dv|.�]K")iR�3i�l2ms�3&�����N����Ɲ��y�i�5*{�;����:N��@M"(���tҘ�R��<&$��k��;��jfu�xuB�˰ef,��F�99+��[�N�a݂��):�?���Wh�v8�3pE�l�V:�ͬ�Aq�����Lo*m�B�ʵ��.ӗ�\�4)�X�{Ec��q�<5#��l�K{{���ݽX-a7���T��ͦ3��^V��b$}e�t��aA�|E)��Z/`}���0���'�tٔ�R駙�W�F����FCz��&�(��Z�Q:a��y#��YwA�OOr�[�v��lj�5H�v��E'���ںӁ�8�Yu|b�m�e�Kb��OxX��c��+v�S��1B����]bhp�OQ���'�8N��홦�����Oż7�3�
Q�0��$m��R��޽�ӛ)�L�#�����s��,�i"񻗍&w6���7���&�Ҝْ����lwL�s���XZ�n-�^�Z��X%��נ�6/zrv1	ǝ�R9X-������G����Ns�-[���	�ؐ�6Hu.9����_j���)JO�����&��U�#�ZYk��'p*;�%\�}6�G�/�^泑�ESqs�K�t�2֛�j��nE۱�!h�%
�,ڣ�:��MԆ�9�%�G]�e2wF�Ռ?-ַsl�k�h�/���hM+]V�eh�bͦU5�N����+�!o)L)�#�}Ǡ�J�ޏ�Gu�I$���1r;�tus�˔)^������C�����q�E����)��s �
��[�e�z��e�W�P��nkm�Q�Qh�L������n#)yuyxz�V`����U
Q�\�޾�2N6Xc2v�$gy��A�!Y�`�E��quk��*���_�X^�
�>VG	�p�An�D܇ۄ,��wv�> �09�y/`����Ȯ<���'S�}{��8��r�%�G����g�T�lA�����C4�����+���>�fk����ؽg"�q�f����K�(+om�/���|1-���3��Q���U�m���ܫ���;_NбV��+E%7�5�]��q�iS� f�|vY�޸����

�JMQ���3�	��H�İ��{s��kq]��qLW>�t\�e@�eS��i:�:^7S%V�pq��QZC�Tr}.�c�L�/'K�����U������B��r���Z#��j�u��E��7#�]�K=�Պ0m^̃�K�C.*�+`h-�Ԃ��@��8><ZP�!�n(s�7�p��՝w-�p�/�a�� ���V�M�ez���E�ڨ>Tv�Č$p�J �:]��N�>�*�}{;(�MMM#1
��Mb������[�]�ܼ��T6˾״H�l�Ԋf3����6"eN��LrR�h\�^����z�4�6e�����;��7�)�:7g����o���r�0��K�&Y�'����\X���G��3��'�R8��C���wr��1VW��J	p>�Nx ���_tX[Y�{)Q�\ShREvQ�"8GR�Y}��ʱ�\&̭ZWRX���&*Ȳ��́n&�0 OV���L��\9��W��cu]Z�����7��z{���{2���H���0��)�J��i�x=Ɨv3nʓRz{��>2A�Z�t6�a� �'r2[�F`#�9fVu��Җ
Uc�a	������&�VloR�2h��W�:d2��֝�KpjO���Hh+n�݄wC�\�;�{,�]�6S�2�Bm@�l빝�L�ִ��{�`|�-��u���L�{/��y&�����V�.����Ў�yy�r�ΝQؔ]{w4n�T�B�ꘘH�+H8����iW	}�u�d��V�iL�@R��+�u�ᇣd�r��c���V7��Z@�Qw���楏3 ;��e��4�{���oC�5�Mރ������*�r0����\1���1Y!��\��)Mh�����	I�鏖�<J��o��w;#�$���Z9zd0Ԓ3�0#H������|�+�0]�]7�@v���+��Xk r<ײ'��W�d���r���]��>�Y���� Z�nd�K}9�v4
+{�>H��ђPWX�� 3L�ұ!�����?�K���S�S|vP���b����'"��tYۑc��E�u�+�ԟ���P�r������b���,�H���פI����ioa(αO��x$�Z�38ZV���A'(�ksk.�]�E����X����9쐨io�]���^�^�2�r���}e���m^N�GC�}�:[+F���a(�P�%�ڏd�7�����i��!K�46���l�ڜ7�'PJn56����t�ѓy*�""��3e�j�4��坼��n���
M͚���L$�+�!�����]"�u�4z�M��1�N�g1w�����'bx]���fqw�n�d"�u��i}:���Z�H9Ռi���TB�N1+vF]Y]a�N��(�˭<����_q��:��9\t{fY��wL8�Y�(�~�WߕӏPY�7Ue��
���LDK��%���)v�|t������CQ��+|��CzPo�$7u�a���P뎰l�]�y�d́��읻��֞$����+ per�ފ��K\&��-�ͷ|�NA*��d������·Dzv���f��Hp&2[��S��z!g+�|U��h�K
vs��P�� �\(Ӕ_d3��w[ƭ��-�T�m��7F����9�n�����ow)�Z��BB��k��r��67�Fք�g�ʭ�:��L���Ö徾��	'{*�Q8��ך�e�!�4J�v���M�����<�]s:�u���J�FO,p���k�� ���X���)��&�sq[]��	O,�6�quqEv˘�'�oA\�oe�Z��=yzx]m�2��gP�,V(��謉A��q��
��]h1�9� Z�۬�#"��|�(bQ��Tהt��y��"��R�ە�t�̿�<��X��;�>�^Ty�[j�iw33��#D=$ɂ����q�)5�/嫇��:hK��v T�L��|��&�j��P��ے��_�T;KnJ�7F؝Y�c�t��k�*���9�6�q��T9�P���,4X{E.73�v�"'\�����]�u[��=K�vVFt�X.�V;�H��)tpY��,��\�n9|�Q�1Mh�u�D�t ����D�#l򢫅�a���,h\˰M԰��v3����������DZF������lmP:�蘠�����f�*{}/���7������J����7iPD�üu��1V�\	ō�6�fԼ�m}�:��q+�{����r�/$j'��]�C^�ӡ����K�
h�Ms��RH��HAS՜)�q3�sZ 9�n�}���"�;k:Ը�)uq�u,�gI��Uُ33Uw4��B����o�s6	}"�e�u�cf�,"��{Ќgfn�̶sb��x��4:�Ul��RqK�L/���r
Vw-m�v���A��_sw˛����.ÇZK��J����/�͝���4�e���!�Y�/�N�$�"r�sNS�d,e��Km��xa�L�B���CF�7�u���6��=�<�4�aX{�[�;>�R����E���]i][x��FC,����V��@\��v����R�K��9�X�.�2��w_T�Yo�u�<�xۘ�}H�,%R�s��6��m*W���D��*]�	Vc�nM��β�?�R�N!ǖ�T6��WMp�@{.�EgQ&�ΐ�<�o�hw/w	ZY��T'�ԧ^q�Ӝ$1o �WlS������d�#�v��g�*W8G���|*�۱��ְ%8Κ`!l��.���5ᬆ�)��-]rI^[�jP�ՑLb�E.u���b������i0�.��h�vށĎ���ܺ��e���{����8���b]��\ő2�An92a[[�b<.�𦨆��ju��r��[r�����	U� T�����2�!eދW'�1w���LS.p!H�a��Hlvm�R���͍���+��Ү�����-|5��+e۱�tF���b����X�5��(RhnY���*e���b�J,��mη�M�>��b���S�V����J��k�@�D*<$�OI�=��K���.xJ�/ZRCO)̸P��}����Q<����{k��
R�S���S��2����1nr���#���f�=�(�f5�\}�^Vm�KA�,'sY�%²�e�]n�ǵ�]%W4�z2�Z+�`�3�g-�Iz6��R�$�+�� ��E����(W G�v�����W:j�V���E!����E�M8G0k�rs0�-���Wβ�����r��݈l����Or��F$�]A�BSSOQɷZխ���5�1�	�ժڐP�'ŻF�<�P��v��f�����^N��������wW6;�x� ��kҔ�:�-��e��%�	����jP��/���I�e�ڻ���]4�[�}p^�Lo0j	�Dͨ��f�����[�Օ1|���6b�p:����ƀu�Wiع$�N��h�B�厬�t��L[�tRݫ<s�1A�cYc���sKw��u(5�#|_+f(jm��ھ[#�k��¹Wu+3��Rd��n�޹��$Ƴ�n1�D.wZ���)�.�M�Ak+K"sHespʸ���vݒ�jd�N3���.m�sL:w'v��[� �t؉��iܐ�;��J�h��&��;�jz/�T3��r�Z��@q����c�l[�t�C]��*��k*[)��R�&`���/�޺t���-���#�ĝ8vԦ&�����*��jF��8*�Ӝ����S-��etr�f����x7�X؅Y��
"����O �UU
�B�$�Z7��!u�;��r�ۨ8�s~\�]���-0�F�d�9m\O�X
�gX|�t�"�nZJ\ɄX��U��b��N��ZkE{,�R���v.�Lz�q��<���X��/:���K�vB׷�����v��%>�EKSfh�^�p�G���mR�� ����2 �ҮBZ�T�=�{���f�ndDĲ�NR�N��i=g��
�M�B���0į�ۇ.$�a�YL�ijsI��דa-�CJ�g`��]�`2�箙e܀wXi�HGu�����yܒS��u����k �jK������!YB��:����b�]�;BU�V�_\ǘُ�-([d7��"�����|ant���[3yA�&�C@�ss��.�k�x�nýn_q�y�^>��8��ȼ�;|e?�mٻ�{.����q���Ӗ2�(�C9[J��<]-q��UQy�k>��I����Y��2w�Ľm�#�ܛҨ��+0�x%e���]��-Ekb�y��@������<��p�r�̔��;l]|�m+��������{K����&�,�;�t��S�o~U�Y�7��峭���;#���q�������n�ͪj�u���i5��u�����ُC�{]h4�ӳD�����i�9P�p͇j\I����x{`K`*�L(,ם�z��{d����881եZ�ԭ�˝w�M����}d"�:��)�_��w3P�0�Ss��1�x�ۇ(�r��V��S���'�������������%sY�5+*h���0kb���Ti�Z�Y�&�cB錇��L�ݣn�#(�����NV�U�k�u�Rc��H;w�^������
t���ߣ�R�TE;�܉�#!�eesl���$�U��(X.ɷz.k�2t~�Q����a- �uW�5�.g���wwY�z�B�J��|c�қu}�����;q*����v�K��6O���)Ѥv�-�ԫ��Yl5��Y��J��9Yͅ-�o���%lUC[*�]t�f��H)���w����G��.��oZ��n���Fij޹������+p���=H�oS���,���%��^]O�5.-�������n�
[�z��@���2�I�&���|�z�4��YDT]�o;z(�5�4�2:�.�A�D�e��GA:-)�Y�C��.�����{r%��{P�ጻm��1fc�Pm�ҭZ�b��w>d��껗��b��x2!HB��A�}d�s���p�����W׼6A��+�΁���G>z�y�Wp4���g��2���G2u(���{�!�����|�^ech���[Ѽ�A�V^����X���:�Gy\�	�=��4�h�&@0��w'��eGz�m�I3���d�������
�*w:q�SrY�����ʘ;j��R.�ܦ�A+ Ɔ��j���vDL���-�6��wL��w��hZ֧m���[;wf����`���偻0�@�EreY˕�gX��!0z��L�(����Zn�P�
p1�2��<�j]u��6w+�౶,��a{ςk�m�F�<���7x)"��=�L��2I�r(��'+w���J�R�������fX�X`&~L �a� S&Q��B���ee2(^�6Vպ�X�ML4� �au�-+F��R�Wά�Q��,?�\ls������B�2�O��I���m�+��IP�D�
���0æ�� د6�S�v�	�(�pE��TaH���PD�,�l,�2����#�$�����BIq]Y7^���y�� _���Kw�嗃c/���Ɵ�0�/����CE����4���Q�;[VA#;ǅ�v�Z�c��rMF���ZO ���z�#U�^�7�q����e���)�Jq�:�5��T�!}�r�^*���+�XI�0�S������}�Zɨ�{+�1�W�-+��#�@tz���Ă�����ɗo�KŔ�v�a�����S#V�yᣦ�U#q�ɂY����ӯ�X�;F5��YM_"�u9�����U���Y���i�ӂ�8\�Z�f�sBr�s���G�r&!�R�����ܘ�[�cq��%RSn����٣B'0�}R�;j<��d+Ao.�l(/邭����[����U�a rL�5��z��Y�9۸�H�/7*�2&i�QĞH��[EO����(۲(���dom^Nm�����n�&�K�A%ٖ72@��ş��.v
"%4�z��:@����m��"ML��!��kZpvQ!]�;\Uƌ�oOp'T��ń	a�y:�֝]W5{���� �\J��͵�Wn������Z���eLk�Z���L�s�������EWxE���kq�s)VP��=[H\�]�H��w��,n��$�m�V��N�(��Ŵ��,�z�Q�Ѷ�c������-i���
l6�4�U�;^�8��A�g;sr,�Ce�����Q\9MVV��r��v�۠�t��ر��f-Ja��Z����2�%8�ѽ���eF����R���q���A^�^w<��ၥ�r�D���f���)Cu��r �E�:�������9X.�i�j�'�P=�%�X�+�c�uc�_X�{��S�)w!aW^�,�2�	Gn�y�������ug5�	���pi����ϡ*�)�3*kTVby�Z.:umg
��,'&T\�_ע��'2P;���^07v;Mn���IWE3�{2[3-�����Vʗ�q�V��vjB�=��U�R��n@\Z��e�AY�0�%�X��c~F�B�h�%�V��lW&�G&U��G/�G�{yR�w�a�R�ک����ybJօ"�Y��D-��t��e7�tS�.�P&�&^�[s* �a:̎�U����V����7}Zب2�q�w��Y(l
�5Y����!�fS��OpC�,\��]��L}ʖ��LTr��sE�
��y�ԫz6��ݴ�Tڬ�B��nkhh�V�X���2ַ�WKhZ�mM���5)Rc,U�q�D���j|����ŵ����w.�;Ժ�,.�{M4���2�Y�e�a�+50�����Y��7�*j�k[����S\�R�}u+��Tb�^��]��T�mYE�#;t��ew��� z�{�]��40�k��顊PnR�km�5����%�[��3��]/o�Xz�um�ýT�Ϝ :&t�[$v6B~�Ȕ�3fGY,���.��%|{{����������9��j�n��b��7��j��f��jDv�F�H�J�YfFN�5��Q�y�w	Jb53Ng�#�x)�u�m���"�.�aq�7���6�A�KGU����]�eT��\�i^�1��l�J1�7(��\�X�����h@6��v����� ��]!�',Cj���yMi�g�a��&+��lJ�*�����FE���jj��o����2����Z������H�����eVx��7�}�EO�����`�:9��s�Qc�E��H��啸�"�J%`
<�w���˝�e��wMĥ�v*E$$(]�w�K#U1�h�j���򻬻V����%vQ�)ޣ���C!���oTJ�lѸā_wA��b�(w,�q�#+M@��R�O:5W��OYK9n��o]����qx�Y�6ܿ�j�$-c����t*�6$: {+��I��T��<�f'��ċ�G,��a�a�w)^u�`nv3�
9�n���{���3@bق�TY�ut��aTh��A�mXw���9Sڃ��R��N���n���݉q�IM`+G
b�͋����k��Ռ3�v��օ���	��j�\E�V�b�ptN��ٝ����Ċy����k�`_<�q�R�
ʗ����z�m+X�R�0Vc�Se�=֜�,��NL1'�x�ssM�fc.\�2��������w�`yY��UB���%aQ͊V+O`��v���hP����e�d���l���Ep[�7b^�bW ������(���*��Ǧ�9�1}I=��h��p�I;�.{���Xb��4��lek]("A����zdo&횺/����n�B�z���+$����U6r"e�d��%a�r��f�rnGR��O�=���
�Mٟr(�KMe�ĈW�\4;3�Qj���;yi낡�vN�r�X��qes�Dl3Fmwk��$���#ٚ���9�>jM}Ĭ��]'��%|�n�i[&�V5P�{��c���FS>S]�=L�И�%tA���3�OD+Ax.�`2N�9��i�@�*��(�%�����@*�N�]�4�d��P�r��ksm<]YE]�o>u,l?=�s�;�-��������l-����blQ��p�Υ�N�
�d
@��f+M╛{��:ckE��.��]�nn7�)����s�  �jް�S�;m=d��it6u*�/pm��&��Puk=A�x�Ǎ���:�nY!],�]펼ڸ�3Y�H�պj��Sk��� �_ʂa�!�]�B�(a	���/:��	�6�V�� 5�r�EK-T۳H\�n�Yj�㐴�v�;��:O��[��`T�B9NVJ�ȰȚ�y�e)����<������+���q�u����oro�h؀�;׆R�w�,=W-py��{Yp+��71\:�O�8�#�-f�s��T�+��kO-�yLLa*M��/��'j��C�U��WЗ;�u�c �#w�I<�ҩO*�p7A�K���Z���FnmFɮ1�e#+X�V1��iuP�vX�����ݮ}����՜���q���`���̓5�-$�˨V.�]MP��떓b�v���,�����Ɗ�1�d�{�1u�=ֹ��r8& ��:�Y�y�)�L��]NSB��g9'^R5F�|�mjb��R?A��q 2��o�oS .�5l�0���ut9G I����DeS� �r|����yz)�VE}N�Om#������]h�����Z6�Z9��A�q�Rv��&��ɡ�}MZ�; /�g7��Q����5�h�Qj7i,Ύ�jb]���M�(�U����w;32�I�f�wu��xƆ��x8�����MJ�ь�TkD��ϻ�ܼP,[\�&#�Ůu��u3D�;��E_Z�T�{6j��ǻ�m	`�E��:�F���w��*\����豴/����x����X��ˡ��%��v_�hh�H��6�nd&q�+�*��J@}���Qu�Q1�)Q�ۨh�v+2� l�U�yx�V^b�be[��i^񯺶}D��88',�6�XOc�q��.��ā.�'6N�V���
�6�f.	�*�6������ܾ�g42��):[0�.aA�6�[K]C��%��&�ui�5W%�>�\�rPE������Z��hALt-)5��ʾ�[IL}�K���*eT�#v�)AըѷX�L9��[\v�_,*�ZP
�DT#���0���w)g1𳒍>��/:���Q��;�lET�mD&۽�!��M{H@��Cl+�:�т��wF�5qGY��`�7Y�=�JfʸT�"��zԇ��$#�Sq3���hTD��w� �W$0[�N�>Ð�%A�@��lܩ�:6�ǩ� ��ϙ��t�y���jmD��E}|��n����r���	�/�#t���$�_n����س�ޑ�Î_����1�K%�U5��:�9��ޗ�0hB[y1�G9әJ��!7�-���(�d���d�!��mhY4Q��nV�Y��b��L���N�ń
3�+B��&Dvum�]�)j���γ�M��(J2eY��^�n	��݊���Ҹ�@܈a��j-g�m�ά�p+/*�&�3
�ֲ�wNԷ'ep�=Ħ2C���R��%)�k��A��vT�p����䆩y�������H#�f��{����gXy�:�С��VnoV�A�+tV�׃�t@�m%.R)�L�Z�������F�]�X�7�Uwl#�h;B����?n����\�'�
`��;�+I�T�W�ԟ3:޺]��(�j�F#���ǼE�h�)n��Δg`?C������������Y3`wYJ*�{yP���+�!]#S�I���^@5qc:�Z�Z�{����ۤ��b�5����I��� ��njN�hP�bvv3*�	��9eh[�a�[daW��%v������x�=v�f��B����0���7�E��	��io��F�/J�e��S��Y&��H�`"l=�[��:����s���n�Fl�K}���ke���!�n��Hq.��RD]�|�+FY�zƵ"X4��s��&]%h-37�Ϥ9�s��ER���sb+0dA6�.G3e١��{B����U��RX+c�A4y�2RϱgL��g"�<�I%�4�Ӷ_;�{��WR��U�����0sC��<�.�429��xt��Fc�6kC��Z���iAƷ\'4�F�$!�up��8ag��Ȯ��+��(;I��Ϧ�1h�[����q��8џh�����h�KLl0Eݫ[���S�+���-1��k�u�����&-ɴ�#�T��|jk,�"7H�$JT��zF&�½��y'r�]��PPs�-���v���5��xn$�-�X�g.,K���t��dmiu�F=[��2��z`J�s�q�[�ɫ#����Nn�ջc�ᬪ��g3�`'X;E�P�s*6�`Rfͭu�Q�v3G�r�p4/lJ�8�B2
����_J���n�/��T�
� o�s&��Pz�2����n��]�|<�E�)Ƭ�j�P[����}-;�]���IH�}O��
�\�cu�w�6�:�l����9[5	V�������'v�����T'�I���-jV۠0fl<�/��*����J.����wv�=y%���3��l�(�£[���p@���w�'gsr�M��,�r1�4NCA�Y�����H�PNū~��2���S8��pd܂l[������;��!ZC�ٯp������j���Sx�ډ��YLc��q���w;��@�v�c�+� ��i���9c( �k'�r�3tޞ6D�{2�lG�=	�x%���w�:�ͪ!�����wЫ$$�'��=X��Z��b|n�u���ax���Y|ɻM�ϟM�"��y7��=��w#܌&�&���\���P;<֎˘j����6�0v>��ZC���ۦ�d�Jh�t�X5WuM!���Ʒ4,U�-����â3f��@���1c4��lzi��3d�Nm:r��H˾�o脻P?Z�td��8q�y�rv��-t�e�ʝ�7C6�a�uY�]]�w
j\��Ptvp�еX	a�\��\�K�8@A ��δ�CK�,X:��=�.,{�dy,�S�t�]!�$��']�e��7���7�O]�ua
���f	T���\%,�,���:��I���7"G�@�
�ա����mL�[�]#C ���2��+9t��UՇ�<Me�F�ˬ)Q�>��	7"
:�6����8�1���\���׋�p��]��uჷskr؃[B_I�.ܻ����vl�����(~��rჱh��6�f��+3�;��F lP�s�g;{-`�`����'Q�������ѥ�gJhV>J\-��!�G#˷;l6 �Yj>����l�|�7b��4�}�X�̩l�߅�isAq�e�������;�
�M�yr��x��4Q��4���*���׼����m�tkl��X\7�����rI*Oq�#r��S�B�WX��hh}2��4/7�;���Qd��|Ƣ(�aN��
���F���fVm�)���3S �ܔ�D����� c*N�M��f1���Z�̶�x%��h����'�:�.^T�Yq"�[+V�F�������W#M�77sU)!��+��ެWԻ&*̬g8��
E*2~ޕ��y�VN8��&m�v-�Q���sLXJgmm�m�F���@h3�/-�'i�{����Q��\�NFU��7��)M���Ʀ��P�.�k�)�%C�f
�W�Υ�u�D<�	}W��!���4U��d��{�Q1UĖ:G�*�p��Mt�ܔ�pr����ƹ��m��"/W"/�ZX	QL#�`�Y��-V�@*���g}4���P4��)��ws6���Wy}�$��:�w� ���SL);���<����U�_e�Թ��8.պXV�ݴ���!�ݸ��Kzn��^Δ���+�]�[����З�$�C��Q�i�z��9}/��M��[[9��W1�Zb�Eʳ��/F���^8:�B�Z�s��/K3����R�UG4e�1eې}�g≯���gG]���km��Cw5�B��:e7�XN��m��@T��.v{�^���5}����M��%&�*|S���㽜�_Hbx��OL��{f �չK]ӫ��n
����e�ǽE��S[��5�a�:�]Ma� �#\uw����.��غ��i��5�9\S�sU����.���U`�E�s!X��.K��`k�Z6iʇ�7�X�st�x���P�1�6�l!��wK.���R�Fo^eLQ$\X-lE>�����z]1�����}��E�S�M�6��s�`�ShC�kp��1A�͇c�nZ�\��V
m��N�{��ƾދ�   ;�e�|������ø^���x���A�I$�I$��>��[m�M�/��T�­��$�&��ξ��q{7'f{�p�X��{��t�]u �(���S�wL!jM:x0d���*cfJ����%�:�Q�WD-��ru��5����[w��:F�v(�}�ZR��J���X�K-�`ӊbT4]��eÀ��X�n�V�j�F5��S���Q�d�
#
���f�,^�|�8�-��:gr֭9P"܄��D%��e��G2E�S��ռ�����$��gB{�*pee\v��2��'�1�T�pA�Q+����-YR��0<[��o+p�t��X��f���mȐ�Xzvk�}}��Ķ��^��|����[�I�z"�$�9*쮭�wq��p�MXX\�a�٦��g�'[���&��A�n�Y:�9iO�
7��K8���T��7*�ʀ�����o+0]-���QE�3���h��8�[����AkvN8�kQu��29`�{J&ۧ�\s]�.��Qv�}�<���]a1w�-p�fMj�ɐ�y���|/��Y��0R��!ż&	��urGI�a��__�'�e#�x
�nN���Q���z�d!H��i^�q��:�e��뻩8Q���Q��L;�!'@�=�:t˃~��r��Ez.�΁EW��Ko�`��œ39�s��i&9I3-���Ld�6��������ţ�5�� \Gi���S�]���r���Ud�6T� ��=��c�e����_L��N�"��((����bbj��Q�DE�9�����Z�Z4F�t�Y�*�������"֨��#cU��'c1TELk��Q�DIE�Q��DAP�U[j9�6(�A�#j�E��kDM3�`��cZ�6��iѶNp��U�UQLS��4�[A�UIDZ�EFkh""(Ѣ�����"�&`�T�QEUTA��X"�h���cHREQ5Z��ө��M�\*�(�g55T�M2�ƨ]�5Dm�f�����Mh�δ[55�p��Il�j�b)j�A���f�5m�hi�lFɢ�4�i���mF �S�k�*Z��*")����RPQ�[) ���h֪����[�U<�EUR�b'Y(�""��X������9��"�����x���Q�{�"])΁�V����TQ/���K����Bq�CZ���fm=��(`����]�͠]f#X {���;(=����v���+��7n��6F��������/~�;)�n#bh'B�t�sٻ�����Y.�{�9y`k_��<L�2jev��i�V��������i󥏸 �"����c��^�Ƹ�ǋzn{m��3]��6{���l���6=,��+/�fh����7�px&����ưn��YqqG��=\�ֵ��4�ʕ�=�qʇ��^s���\��z'&e����?|ٞ�S&��t�]W��כ�~���9`��J���d��\����<�4v��;ϲ�ce�\o���?7٧�G�N��M=���^����:v�9�7�͚̇�k��i��J>:�� �3/��o����=�`{�#7#M'U??-��sO��)I�,�P���q�Y�n�H�h�����YY�h?��V����vh9f؞nq�X�^�8�	E͉�\xm4��)|�e�JQ��kN�ڗԥ��2��W�����������]{Z/SέJ��y�*�`KC��"wO�vC��a������Ӿ��t%��-0^�25��t^�2�rv6FfR<_Dz��O�F�������^f�RC��N���̕t�Z�M���W��Z����tz��r{����&:�]�s3�c5s�X�T���l{ގ���Vs�_��ν��6+�� �O�q"x����x�_mڼŃsǁ�����>�3=wѭh[�Hs~/�Q|h�ñ������i4F��;G��v)�T1͞��9����7OƎ�6�q��٬�����|A���Q'Zso_<[���FN���
I�Gr1�z��T�h���&l�Ɍ��i �0t�ͧ�'y_���5-���,����g��|:G�A�H���1rv��1w������{ �������5�/w��/`�k;��R8�V���]�gZܬ,�4/̱��z�co��^����������ϼ2şP�T��N�:����+w��g�{d�P������0�7�|~�yz����1¶�g��Yz�#���u���c�Jfe��V�����w]hڬR�խ�KzgN�G/pxoS���N��jw�w6RLt7��,�w�	��;ܫˢ�KXL\��ُ�2�ظ��[x1m��'o-W�pY�s�AկD�N��ԫ�(��G�z*��C���qojM�m����������l�y�en���\�NOyż��2I���L�(vW������k\�cs��I��u}4D�]�M���T����˳��]�X���U�w^s��e�rD��{ɛ׸��Y�e�{���o'�s�P�r����e|��O��Х�q�G��W��ϑ�����/_���7V�����l��&3�S5o�T�ؕ��#5�_0��[�/�Y�u4���d�c���d?y��ͫLX�S�����KI�>Ljq�+�ߪ���9�)�rF2*�^h��{�-��|����j�6�s����ӻ3��<j:�n����whCޞ��U�ݛ�x��5����Ӽ�����z��w�;��:^�,^^�=��^]��7e�EU=�>�X�Ζ=�{r��&�^�>f��z��x����^$ߟ{%�x��K��\7�+x
�X���2w�No�B�����t�~��UO�O�_�9�p�b�vy�S��0d6�7= ��TO.��07��?�?��ٺ9���Г�CA�؂�����WY����P"�+UIY@��E�K��]����ro�sw��h%Ǧ��*')n���vC�5f���������^�ug����l��2�iy�y���l!��	^[������|=1ywty|�c�,��ʁ`�K��պ�c#�p9m�+ON�&�<�&�t�O��.Y����tũ{g9�!��K({Ք��Z8V�^t�o��y��tъ��D���t�.$��U��]�����b��F���dW�]$�i��En�\f�k����z���c;�<�g�S�k���ۗ3������3�Y4��~�^��K�s(���}�}���S����W���-
�u�~s����]���Iɞ4��eOu�q���Q��9 �������I�]'�b�g�4�{d�"�Wb
C|hӓ{^�.8�]�@��ll������S�Z�S��cfL�<�~�����F�������g����ű|��3j+��c�+�����1�cqO!�zK�ד����ջ	,�z`=��\&��lgs�dP}{[R�TV��c~;h�Y�ݣӯ]ٻ��)�r)yS��A�93���Pb,��}Sp:%�n]��׻	�=4f�,�i��+C˼:�P��8�����T�X{��0������t���孕w����7�H�߷��}F3o���S1WL�4��|��l��2��m!��z���}���/�z}��!�6<_�O{~ý�cڡ�YD�~�tn��mls<wA��#�!�{�k���[=��.2��Q�=��׶������_�+k�w���^��q��V�>��!�m���ז�(E�^������>U� u�yt�2cg_����&��Wm���я7]'Oh=�NE�>� �"	��oV�� �����KL��'ľ��q��i�;�ux워���K�Y���p���L��P�鞤;[q��n����2�e��|�Ns/��'gѼ:}r����wf��X��k��'/�Q�d>��?y0�Fa�B��z��<��Z�۾x���zS�r�f��}5�M�)��A.�۞����r7�=&Ժ�Az��HP
;<�c1$w}F{$��S���͚���߂�;����[Y-e��K����0\��ЭX�s#n ;������7q��Uه���Y�u��0n�t��%��y����K&�y���u=!��~�]����YA��`��N�n;�o+4��w�\��׸�C�nM�&���72U7�-Tt�2�8e��tw�Y�zLT=����t�1s"6wzKGN�����0뛓��Nv�P{��ә�r�3�>M�|���V����q������<ДB�!��z�3ޞ^D��s3�ؚ5ڹ�*�Ե^����q_��UV�W�g��fү,�|<btz}Ld�%�dȨ췵q� ����h4q�3(�u7l�����] �q�7X���I8�kǻF<��e��Q�z^qk��f�}Z���ڼ�x=�s7;����$V�Ϭ�E]�VR/4e.�u`Ҥ���E��L�H*�ø���5G�S����ݹ=�c�����)1��t�z���Lخ��=�q�3d�Ɉ�P�Aoe��_cn@50yS��+�o�+�d�
v&姙S�-o��LT2��⚒�U��*����[��ص|ݯ�����B��3o�"�U����� F	�o�Y���n툅�u#�Y���xN2c���w[�d��m.�Yff���}:��i�J��*���K��Α{��`��3�l��nD6�냦��vn�3N>G?�7�M8�dנ��s��g��XK�r\���M��&�O;��>�k{m���x=C���5^�p�֏�uIJ��ط�ķ�sE����A���+�G���������٪����[�����9���j�l���,��6E�I�|Z���;���E�o��(�`ǻi������9䜙��T*��Wj>�_^ӭl�[��>�(u]��n�O��M�k|�>�߅�}b�I��M�8~�f�g��$*e3���6�-n�����7���G���;����S�/CU���ɻ���oz����%5���CW�k��P�����n��߇ݢ���V�p�"����e���/]��0@�boK�q��ǋvH� ��b��h��eK��P~�o��j2���_S>W�ܕ�L�2�s�V�Z�͍"̙��YD�}gu�}��W^�ԓ��n�)��9�y�#:c��w]�vҺ鰬{|��m�phR|�Ƕ+�p�x�(2�5ٜ *֖u�We 6}�<}; ��vѨV�<���~tݏs�ĜN���8er�Wv�]�9�����P��{3=',�P����}�Kُ��q�����ٸ\��Bc�o�P���(\�����9}�������i��f{=��f�]./�0�r$��c=�⪧Fn��3t�6X�������=�]^���f�ݨ7�.G��)��^���j�T}ǎ�w�]_���T/�ԫ��{fo���o����A�d��A�r�F�9�l���϶Ms}��*>�=P��Η\�Z�,{ޖ='��'§��\��I0��[W�����wN,��,p��,�'����W�r��>������C�A3fU8߳nH�o>�mi���[p:�ë\�\Zt��}���_�g{�{��Q�ߕ��Gh�Y�ݼ�������3�4��W�NC'����]�IXD�

�K�L��J:U:�v���/��m��aNU�{xӡ�;���s,�rWEΟU���)xw�T��,P��.��ۤ�	l�.}�%�O*M�Be�#W��Fm�pi��]��g+AQ�ѵ|5��]�V��o����#�̛�h�H.� � &��5�IR�iM�V��ͩ�z!�x]���q���=/��uR�;3y��p߄���1��q3�$��u�C�Nfy*��i�}�Xϫ��S�r����V�>^}�;����G�{�h97�9C�uQ�����Wyӫ��T�`�]l]}���v`�Fq\\������k��2c��۞�|�^�ƻ��K�=�y2ǪZ���b��zf���W����/�����B����Ĕ����>J���߳��#+�st����[މ�c^���0� m�pm2����<�����~���p`���T̯V�����6���BR�Ge�Kԣ���N3�)�ó�'��zJ��>/4x�7gA��
~;���_��;��ذ-E�˞���;<<��ߟA��K6Xv�3c��_hoݑE��2�+�ϥdπu��&�Ll�_��Ě�����1��uC[��*8�m\�	�S&������ή����t�a�Q��.id�:@�����/cVVɗw��mg,�(��Ѵ�M�/��s���hN�@�B�)m��L�J�ν㛲�Lm��|�P�IM�v7����e��F�y͞���3ڙ��߯�!~�gϥf�3Lz�6��;1�~��!������缮�5z_�*�C2NU�G쿽\~�+�]J�qv�[�Nʱ�Lt���M�y���zx��otx+��+���ޮV-y^��%Do��i�{r��=�s�t-���=�`�^L8�/���a.Afvr7p��3�}v*��Jq���;<��o��g�>�3�QZ����޵���'�fXù}x���s�ҩ�@w���6�ݭ��6����w2�������[�V�Ƌ�`\0���l�����T������8�3;c�z�i�G+�9���36�:�Ӽ���}B�}�;����'�>��@W�,�~
���=�8צ3Ԇ�uJ�R�ʽ2�.��v^^�j2-��I:�7{W�<u-�&EF3WS�������~�}>߸��eI$�I'�*��h\'T�c*		o_��4��7����M&AKJ)������y;S㝭�X���ި*_T��8ivw�!��DP��Z���|��EN��CZ�\��=&蛲�{6<�[��ʘC�DH::u�P�����F��y�\��Oq<]s���V^��ۙf�k�Ш/�tzq6+r�N�nYso1��١�� Q�����d�'J\D-�K�m��0����y'i�:f�wW�s1֚��+m��~��5�я1�V��2.��R����7�%nWg/[rT��E�NWv,¥uŒ��b��v��NP9-��T��F�vb���#�������H#EekV֒:�Q�JǄ>�FɄ��	�Q�YO��V&b� U���mԮv����,j�ήu��TN�5kDɏM;x\ln�f:HՃ����+����+>�,6چ
٘����R5�p�+s7���]�������.����`�ݝ2�y��7�����!��C��O*>�s�9t�}�ev��V��V�څl�16�ƮS1��u�dn�Р��
�����5]�2�ܵY^K�f�tkr���Ke�|֍�d#؆�q�|i���e��=9X�k�p���v�h�d�:ɦU�`D�G.�<����\ne�t���%_Q;�Ǽ���w�ِh�|$�5��]!y�>�Hp�OD���N�d���q�Urf^��B�Vu�N�� �%����ך')#��AKR�Ywyi�D��7Y�Z*�a�`�`���D�h�{US�R
Y˝Ժ����{u���ʸvsf���V��#n
�\��t� h�:�L��`3��)k!�klSU��v3_����P�����0�;J��_r�KY����x�U�R؉�^�̚��v�82�9[u)���`ǯ�xh+�lН���2EA*�aL	�\xc]�eZ)9��oj�N���<
�Ssl�LJ�}s����u㛯(U����ws!�k�e�ZZ�������<�c�=��ڢ�Hi���Nnt�EZ��k��qr���riC��"��%*B2���݋�T�)y�7�����ENGnX�����.0j����s'Uŷ��w������b:���
��Ո���3��:|��7�lޑy����My��Z�����Eo�&�ZY���@�Wr�!����]�v�v ���-�L(.,Eu����w��]�*����]d
ȋ�r�o
V5�5N'`������}ko�Z4#�{�re1[�������򽤸 v:F�p�ol�r�G��Hn���J�a�t&����ҙ��a��v�P�vP,e �X��C�wPv!�S�^��XO��n��"$:6�aqX��;�9�����/Oj�5����S4p����1�f)�/e`(����m��NN^,ww�v���t�st�!�W׫{CUw���(�w.�8V����:2c���R��O��C�(
iӈ&�X����" ��lj=���EIj���"N���V��SU���!��*(��b*��i�=F�+�D�K���MREEQ4m�������[cQU��j�"�5�Ѧi	��EDRUkETEKPT�"�-V�j��ӭc`�˗"�J)���1��6o,Q�F!��S�A��4QUs("^X�m�͍��b���D�j"�*�4QE���/*9Q�c�N�b��*9ry�QlQN�"i6�-���Z�h�[N�8�kX�y#���y��^���b1r\gN��P\�LX����ի�kۜ8sADQ��#����9�r)2V5l�Mm�jسU� �ryp���I[\��vN<LDA���1Sȸr8�w-A�.r���9�����Uƈ��h)�jn�5PV٩��Isj��DHr4r&L\�9gXqL�t�Pk��46�1#�p�孱�PW��}�w�������?[9�Ȏj�b3vm���Q��	���'NY����1�ջ�c����eΑ��'�V,茬�yx�fc���:A�9�1f����bt��h9���
^�BA覀��z���_D?i*�A�����[��ٟ��h���՗����"ŗ�L=�/^�x�Z���H��L�W�Xu%t�dÇ�y6�ӔI��v�#e�j�'�:��r�p!�<��~hj�
Lde9��G>^��W�G�vn�2�*Y6�����~<�ga�������ooE���S����o�K��-�Xt\	��O
UX�+ڊ�;�Rjo4��4t1g]y�ѺԻ�`52�4^���
���p-���[��0D�YBd${6A�BY��z�cDn�n�,��p�	�%�{)M2�%Mw����Ο)��= ���]���=�G:��5�]`�7��!fIz��(I��%9��E1����Ϸ�"����v{d���3ڧS�����a�n�2�0�ٔ�'�iRN]�9K�E[\Ø�����݌�.z�aN��2]x��I�[W�A�t �W��Cu���¥�@�	��(����A.�R����L������o���
@-�a�?y���k��s�׆\�=r7X�U�e�x#��������*b���!W�A�������w^G.��=+�c��bE���\�Q_.vV��i|�
�	ݑ�Yt���40���E2�
�e��fD�ͤ3C��xw`u��
ٯQ���q㬸�-���%!���{����B�ff�牎7�D�à/asׂ��.b��1S�L�Oi��l���#���8n�<_=�]{,�l�z���y��������U
����n�pz�؋ՙu�wo��^�뮓[�ޑE�9�z�{�O�o�b����t�v��w���Лv!���1f�����!햽	P������I86��0VSH;@��ԟ�z�5���k�#��Ս���js|��p�ghkLL,u~�����P~|/���d
.��]�H&:���z`c��he��aGeΰP��6���w���C@ێi0S���}ھ2�}�������WD��?)�h̾X�{Nϼ��^����^m�+�d2l`����L����>}3m�kv~mU��3X�u�{��p��p8^��*�.�g9��� [:~`%��qy�y��z`��b� �鞗J;p�V�@�QX��zO�g`�YX�]Z�@�c�d�C�p͞A@������]|��Y���z���x.����桓���2ױ�):Z�J2��������������G��P���6iY���C7BVZ�w�	�����3���:.v��̧aq�x/^<X��O
у�Ms��B2nŎ���y�wHuلlxZ��7nq��A�kWhF���GPŘ�-wk�Y57M5�Z̰bJc<�kU��`Yǈ�����3t#��t8B���>��RrI����i���!7���k�	x�v��v�}�s�	�~w���T-X�Ew�c{���v�ֲ��us����qm
��z$!�H�H8�F��eg<3\1ch˷RYp����!���/vI���΍���ׁ�8^��[�	;��PB�kL>�@OH �a�,�zʠ��]����o�q��u_a:�}�6Ɯ��̾��Hk����	��(�(���Y���}����e��ΐɞ|GN�y=z�0���U2����O7⤰��B��v#��85У�p��K��}�R)FT����-j�S�I՚N2�7�R�Ŕd�>���f�V���A��sۇ��0o���,�e��n���m"�Ƅ�m��BՇR��[.��Vz	{b�q^��<�/f�)]y-m
c0��-~�T�����G��NZ�>4'e�nt��0�@��~N�a�S�+����0t۴�<WN�f�l����=�rw�\>�C�m�7�r�u{���0����e��>��������Q��p��虘f�m��l��\	w��`L�����Tm�2/��2Y3��S��T�T@�E
���m�ۼ�~���t��-�<��\��P����[�zF�[ܽq�y�l���*�V�v��]s	:-�B�8��L(��/�n7ٯ]�.���n��+���:�^��R�M9�u�dbni����a�/���i�ϼ<>��ŏ�=ڮ��>����C�A!�p��r�v��-�����������]��F�u"&�[{u��f�M®t&���g??�����H<��C���B�&���.�L[zW�E3��&ւkt4&-����ڮ�;�o���fMk߄�cV߲�[����]ȞIP�>�[xj�w�Y�]�l�i�k�Fp]���S<�?5�#��l�����so���a	���'��
fd�)��Y��UqXw��	�׬z������`�q�������G7:��ӷųbWUDmn��C�zo ;c�&�B*��E�z0k�<'�����<�t��3����CyD��� ���+�O7?N������ٓ�Ş5�u#�)�y#I�k�8jSB}��$fɈL8r�|`UW�)
�gN��ܯ��Ug}f��'���0��<Sx
��1�噃kؘLZXL�ĳvD(Rwz��ݜ���X��mI�HY�ZrD��I�U{�+0�oI��~n;���p�5E�?%��:�b�o+�:�$�>y��[a�U;4]\���a�qv8�0�-Gs��!�@���Uk���?��r�Uױ/.��f�N���i	7ڷG4��[ [*���������6Stq]{���j䏅�4k��E���9c�O6i��+�\���'WyD�i'D�݋�z��1n��y��bqG{�"W�J�^���m���x�a���u�����W�D��S���Ds!�G�í~��mQ�Z�93l(�2��V��4�u�ת�97����]
�,na�y��{�0n�����ͮ��v�}�6ɽ����Uq�Sp�9ڱ� �
�,�����3�@�vS2Oa��p��(�x!�:�\�{ܞ�xf��6�[��O�W��;)d����!��@�LW��� �Pwc�"]� ��!C~uy�u�[[7����8B'f�ؕ�ONmc/\� �
h�BB=P�_E���a��w;z���+��;�Y�3�ZX���!�z��^=���3p�4�Aa��#;z'�����)ƨ�F�Eu�k &�a����6 ������!yxϠM���8Թ*f��(2oI�+5�W�,���6z�L��AV{>�`�y�x^
_�܃w�-��Xt^}��U�3�Km��8�`��f*��j�C�x-kC6x2e�%_�mq�����!�@����_`�Ad@H84R�/����[gH��yh�ɭj����"�
SL�J4��Dn>5{gO"����o?���R��w�z��=��M$9�Y(Qބe����0����Q�ӝ91��ү11�)�ղ��l��th��� �7i/�������[8���T/TTTB+2���J���u���w*E��C��buaR��r�UΊ������T��]��{�zM�ℵ���f����U� ��Qz)�|"S��S	Ml��������`�$q�}a�O=F�u�_=�/p�f�^���P��ư�0SfS��4�7�`1���F����-�%{p;��i����{\��졲�������-��G���&������6�^�0�v�0���Z�C'�t�=<Xn�}��I�2sd�!���Jj�`#�%��1���G4�z����i���U���	�9,�f�S�V2ڌ�!W#�C�c��'�q����ь�!ʗ�B@p_�=�f����������v�!�'�nQƭ��<�J~b5)V�u���@Uf�MV�ۡG���=��ך����C�Q�����M�:�NçT0��Ba��5�8-���b��m�uv��`�Y�ǉ4�{S�����x��}jd!���;Ϲ�Dw4��a��`��4��TQ`)?t�:���ݘ�:���5���øB^��q�� ��bac����k%`oP~ys�Mq�.��]� D��2_oV����;��g��Å�-���y��CdK�CF��i0���P����R���F��v��6$YWJ�����-Л{��n���2�	�ܬ��CԲ��[�E�p��U�K.�B`�tZy�*U��4��i��k]�F��:ŷ�Z��s˼��5F�X67k���Z���R�=��=#y�K_;)��D���ހ2�l_s�쫾��C���=��/m�$w'ȍ����X�o�d��8�v����y6�ͼ�.�/1�T�a{�e�P=<�SV^5�9gB�a��-�òg�yS+0HqB�_�w�{+&�W�3���8ɽYށ�	�i�w�h�#D$�v�ӌ�y��������WLN�:�����Ђ~c��r���V���c��*.��3 l7PG�6gkꋞ�DZ�\�ėit�&�d��tB��ܢ���D�%QaM^[�����%F�U�*;q�����ǵ����Ƴ���P���'lܗn/�1j�'�b%9��O��긖hwsU�h���1�)F�0�zhXN7�HB1�C�>��_K17�]�M*[�M��=S���߆=�
~�g� kL��4�Y}�[�	���!�!�O�= ��dS&�nP��1�!��6:!kvo'e]Ry䘦E���k!��F������ 4(u������r
������O'�w�;
-�N�
Vv�
��tKw�d��c�狛U�%<;�@�ǐ��ڙ�C��E3M����-��5;�cn��'V��f���|\*,ӎ�cZ)W0���>�jp�g��g�Q�y\�M�jI໫��i��P��T� ��F%Za��D� ��!�[�r�9�	NX�ky�\}J��W�J�U�{o����t�s�x����,�8<���u���n�T:�N�2m=o#�Cz�#��G�8r�ܩ/gY:<��ƳS|< ����k���r�����������
*�9���hZ��▾�����{*	{kU�mҖ%�]\�c�v�I��p����}�(��2�� >'4'e�mgQaͅ)6�ۀ��A\��7y��
sw��ʼ�mj�t/^/a�ɑ.��ƈL <F��D��j�Iѳ.ŽD��0P*#n��
��0^�%ځ2����f�sl�tg/:��  `L���S�xNP͸�����v���J�7�.�ȴt�$? �G.�i[*ohlg��`K{�gů֯���z�օ:�esĽc�^����(<�0�z*�!A^i��t�:b��yg��5�g�jc+[��G�:���xE0�ȹ�E�U>MF5u��R�ǔ��� ʂ̡Fң������raT����|��o���LT:�b���:m��Ҷq��mT�5t)�ѐ�7����L�[Y�s|��n��;�-�o�B�Vte�S�;@ Ŵ�8�*`$'��CH�S�u�.�u�K־s�#����!�]%	�:�}BН����x��-��$8X��|�pBp#�G�U1����������ҵ�oAw�J����}��%�6�yg7�1.}:律X�j�(�D-�zmK��:�b��(�m�q��I�u3���TU�K����hn�'b:;�VMT���L��s��f��u�����C9�W:�q��;j�ɚEx|> |?W��{Kӥ3<,�A{�ƽ#�d�E�K�)��&��)��׵��f��a}<*)�G���V��ק!XD;f��يN�_*�]g<S����c��S�mp& Y����m,g������Н���!L��&6jD�N�ʮ���Z~k�x%��;��{�"��k���S�^���, �����sLP�n��N��0,F�.��0�-Gs�,��i�}YZ�T^�-���y(_Z�=��~`}��p�_�vi�\��:Sm᧻��nQ-v�M�;��o+/x瞥שG4��f���?OH`�à<#�ȇa�4c�n8�)�cnNl��˞�,W��L�̣���O��G6��,ƌXgc �f�\>�E�ټؙ��{���7k�8OC�Y��۹�q��^=$=qh����zb�Aݎ�;�R_-�B�1�f��X.��bT�<k޿ƃ��mc/C�$�)�!>G�A}��+��;��n�y��]}
��q,�9hjC!4�{d���^=�����4�4/����WA����a~3�h����b���P�c�^�ժ񡢳Vܝ!#�W^�O�y�iޕ��N�*�����Nѻ���������H˻���:�=1{��َ2�3���Ҁs���}i���d��Kf�������99��7M�-ԜC�FnQ��FDc��������oVR:S3��]�a����z/6�ӯ,���- /	�ё�����y�{ӵ��Ee3sz�vA2�H��!�Vr�ֆd����͋O�ǫxTH�x����E��q��AUc����v�݁EU��ьQY�ا#���yY"u�ɔ2���t�
���z�o�[� �f��3ה�6�=3�S_^>�YC����d�sWD �qxd_�SL�J4��#q���ȧ�p7(�_�[[��3��P��.�k��O0�A}$�tD�I��"S�P%�$i5����MQ}�z9�ʲ��z�βW�=r��3cX����	��ʀ�,�H�)�i�)? b)9Y�y_�Ćl|/�}�������-�1��ϸ�-�?�9�h	�����~;Y�̇~_�#U����/I�𩒯=ǩ�q��ڋH�]4�$����C��s��,��%��w�C:Y�-l��~�YcN����[BO)H��z��%�T8؀hyD��}ga^6H`��0쟌]Lc��,e�rЌ~@NȦUյ��)?6#�eG��[
����罫��E���J~_����~�����}��o����=�4\�;��OQ�h��sz���/�-Q�#�'C�^�6l�]% ��J
�G��u�G*(�����_]�]�܏b��"u��7u�J��-���X)�!Ҿ��f���fj��S-��]�P�7&n��[\ܖ+��u%�1��F��Pru��ن)T+F�c�Q�v�ϰ����U�e&�A� |tm�}So�P2�?�3�E�:�%�5�ud��;����I)hc�#h�������1�C�8�uE�PX �P0j`��9�R1�H�:D]j�h��w7���%�͡{Y�J�f��*q�� !��:[�0ޜZ`PV�u}�":t9���Ϋ�+��Bv���rR\D�C����T��ذ�[�_Gvk X������8`�Lخ�sr�M	覜K:�h�v�]=;RWt�д��3ʪ�mn��d�T���rw��W�qSd��H]n;�M��j��� 8[��.����m*q_C�ܣ�U%:�nw��"E�]�ғ���+���7�n�DQ�J��7gfX��450MLR �\��Mv�;{�*�o3���:��^F���`�V���ɪb grk���]�����q���]f��9<�XA���I�,����Ҭꈝ�Tp]�ݢE'v�6������⼠f�x�䥪���vĒU���25r�lX7Q���[�v$�{�t˘y7t|��`���װ�m$�8G��p��ZC-�b:͑��9u�9�_��Kxͭ����R�S���n\�I��2�7�����EGp^�)݋�W���Ф
�N�r�����ņ��@)�p��|�u��Z�����Kw����KN�hTe,Z:�t�&m!P�E���{z�ʉU���e(x�Xr�L>�3��|���Eɩt��uL�[e-9�1r�*�m�u�{,	䮝X+'W;
�ִ  �(Z�3�����7h-�꽜���c�}�T褒����L��<��pU�R����']vc��5�ٕ�����=���0A�n�:@S�M3_�5үNsZř��'!<霂��s��x%*cm���-*gm/�,J���r����W4��l��vn��{1I���įWE5������Ą����s5<��D�˚de� �G�[���v��d����ڰ �9��1��y�VJ]2��W�u.�4�a9��B��������=,.WS��V��Ī�iЦ�
�m���.S�И^�y]�� ��:�̬��}vfGΧaHgVL�Ⱥ@��r�]������Q�=���j��]w��1P���F[��Jm���Ś%r���l��xߋ�kz]�ƥ�!֤Fep��T1���J���GF䭺�#c.Xʢ�e�1�����*=��ya���%3�n�K_m��+x����A��CUX��$0g<7f��s`�gaWO�X��xY8��y�n̙� �6���j�c��|�Ce��9�}�r��uց\�.�g*�,���f�<�\l����D(Eq� �@��"D�4�ל/�Ϯ0DADHp�_P��X�F�Wȶ�í1PVڂ�(�tnpxF٦*�j�" M�QV��T�R�ܴ�"�j6ڋc5��93D���7"������U�
��:��K���&�&��	ֈ�*	"�-h*#l�UALDT�ܗ�ͦA�F��V����PU��Z"��u���"j�M���b�sj�h(����ٵ��cW!��i�����*���	*��(�����y5HU%1%LDTQM%Nڦ�51AL'y���O1cQPTT��BRSIDT���QT�����G��&�J
Z���*����^>��i�ӧ�N�9��6))���5TSEj�CL�\�I�ş���oQ��ߏ�恊���ׅŚ8��m5r��i���Y�҄��o�&��ͱ@���
ݪ�[��M/���'�s�K�~x{�����ӕ�z��+��v�Z�;�hg�R�p/���r��ؽo����@���i�����̘����-��4Ali�:l �Pj�r�[Ƅi'�#4�YM �O%��T�+8���(�i���K�.{��<
By��'-b&9����z��ϰ�P��4]��#����m�6d��O������켲�Ŏ*�Ơ���uz$sH���GE�ӞޟM�EveK��ڙ�_O'jJq�j�N���o��x;]��2��!�-�}�:���~poKf�᝽��u�j�;,�X��BFu��g?��l�瞝����W�b����*�l�Ы�ai邹����]sz��0�?5���YX�]Z�@�c�VT\9*��?��2�
쎋����8�x�d�u�PɅ�^�k���XZ�R�%��v�"6�S�P�Jw2���ot�3tJ�Qp�B��H�ހ�K5ׄ�$��4_Jb��'�)���Y�����f����m�_V��iu+���6q����г�8ށ �ƟC�Ll?K��:��"|>{:/W:����6?d���x�(#X�uq���bfh��4�� �n�:��i����3�by��G�{w����w �:�w��h�$�q�/�FS�`!'*�[]��͊��k����Ytsh[��5%Ciƭk��K���˨kԲĬ��2:��):�W�}^���{���ɦ�K�HU}|���s�,��y^��~��/^w�xa#F@A�v!?t��ΒԺ�a��o&���Bء|i��`����X^4�摴vk�����8{h8Z�[�nuPX�ۀ�=�����f��t'"��MУ`�&�0����O6T�4��0�û4vC������΂���[�t(l�cZ�@LKО��0jq�Ù8�½k��̩�hOtZ�`�3/	v:��Ӫ�:��?2����7�)LnzG6�q�j�J�a�Jײ���{���ya��uJ�:"�qw*��y���ƃ�a��̆�5���zv]��΢Ú��@���~�/�>f��Zȇ�b�ټ��nô�U-�@�/^�3� ȗx�h��#m����d�����ݳw)A�p{S�TM&LIv�q�?c�fa���cB��W��c����^x딉�;'\�t{{�M�0}�,J�� ^E��!�(6z�D�O��\�OplgƗ:���+F��p�
B	q Fd��&���f���t��Qt9���5��t�<#��u�8K�Ύ�5~��4��������sӡ�:�'n_)b�N��v���ݷ�f��,X�v�&�s� �7EI�qH��0�M��qg;H.�y�2L���0�D�Y��(W>a!T�/I��в݂'v��*�H�x���s8hn@ F���u����x�/P��(�x�,,2...�ؚ�j�ʩle��㰃*Y�(�<9M�zᚲ6*Y�8n��r-�`��sk�b��t�׃=RZ�#��t�.���殂%6�à�]�o�}t��w�����=�B�0��V��^eA=B��vc��}��-��6i��VS]{�ۼy���n��)��LT"�[�]�}Ǆ�-��$8X��|p��S�23��X������`�B�@S�&�:fRtY�u��<�$�&���=��}meB!Ll=���4N��l=I�װ���w�1I�R"�s�1�]N�_��]��:µ��we�h]��5:�<0f�t�g��8jD�i;��YU�����PX�jQ[bK��k���{�+zts��Iĸx;�XG� ��kH���;4]_��c�7P���Va�E�F��6�������5Yޙ��-,C�z�������#�n�C�Z�Bvi�_�KS#	�	���N������O�7��3�{	A/�{��B��m�g9�!�8 �x�S�;k��7�P�f���&.^DU1߯GA;�-@�5z�P5t`�����|���u1��=�[�	�!���=���x�1c�Ó��>p|����z�
�s���is���׮�mP�C�9��J$��]Ѡ���p�:��d�2��u�3��G<cy��2�����ڢ+�I$�,	$'��o	}W֝��g�W	Rc~eO�9O��G6��,Ƽb}a��8-9^!��v��5n�%��n��T:~̀�6辒_��zHzZm��uv=���͚ɝ�!�<����C�����Z��E'���t��9����^)� �L5���p�*�b4���@�����az9��!�Za�z
���|[Ɓi�n*f��L:X��~dC9J_��z��Grt���[d�8��Ca�����pa׫��gɯ��o?���Iw�����[�Y݉��l�eK&��;K�zv��=[��5E�����X�mk�WLvf�U��l,��H<D���(2j��4�F0�ј��z���>á..���l�O�}�s��Շ��� �����C%W7;��h�Ƚ��4�ģI��7�=���P�w����J���\���N��]�*^W�|�_I/C�%:O��Js`j�Lh$i5�G�	�j�+,�]o��m��\:�����!)f����p�0SfS�y�M�X�b)9U��p2��Z������V �ټ�?U͝�f��*�.�ɼ�EX�̳A}�kF���:yHnmftI�ڋ���T8�ʽ���D�҇�Ҡ�0�����&@e���oVE���v<;��v���vB�mk$[���Y{���B�Y�Tx�.1Z�f�b�NK�c�[L���)U�P( �T�To{�x�{E�8����2�g�s|z0�y�<�,"�@!<�G������Λj/~¥٤�F ��_+�z���ê��u�]�	s�E�u.�a�?`a��a~S�P�S�׆\�H������m�r�訓׫�*��"�mH�0�
��M��Ļ��ga !��n�w>�-��E��6������ۉ��c$Ir�H�.L�V�I��#&�eG�S,ٯN�ۃa�H���Ȧх��Ыt(a���ً�:���Yʅ�u)�Pc��t��Vؓ�@��TWv�w��)61�[ݽq����'lB�pmg��ŤC�W�Ŋ�t�C4Ў��I����0K���b���-�V'n�7EtowJ� `�tɨ;�gg�����<:����md�ݴ�p�W��	��5�g!�8�0�ݪ1��v,K�8�e�m����8��o�q0��Ӎ��t�g!�+ɽ����Uڼ���i�wI�j	N2\��!T�_��A�c���v�e�	d4V�NǯWM�j�Bj�՗����:� Ũ���3���l� [:ya>�|?�ڣ�o�]{��{n�|P ��j��{)�8��*� ��U�,�k����z�V�U�2bcF�mįQ�%*�9��r�e��Bk�'z��"�b�Ωj�����"k�p����V����0�i�%Z����B��5��CEѧ��Z����=��f4�K�.���҈�"4��H?>}�������|�HW���ُ,M�'���������d	cA.�g����)���;�ʈU�&���7P��;�@���29�tc&���}2�.|���Z�R��1�aKz��W�#yK
ds'�Eê��3Ĉ-�Pe��^v�nK��L{���$��\���rll���:Gj4����-X������a#�-�W�q� �Ƹt���!�_K1L�Mo
����voe[F��<^b��I}	t��78^���`Ѱ!#a�'��G�S*��/ul!����1BɧijRy��m�u��̷���s�s?;��z��`�.t�;/vwC^�d;]���s�s�I�N�a<,�熵P��Q���a!<;�7�F"6:	�x�N�~��@>:��`����|���W&�Yb}-n+x�,-ts"�k}9���2��IZ�q�3q��zd^�9`����C��BcBzG6��4-[�X��X�e��9�w�F¬�U�l��h��'���w2`0p�3:����-��E�1�z��]��{�/�&�W����5�/e��M�&<Ct��
�Fr:
1�S�o���w���x�Weva���`u:��sK8�ge��ه9r�����σ¯��M�E��g+�Xz%�!W�q%��#gfΒ7.w���������B��E�{�Uk0����m
�s��{ô�j[��z�����zU���"�f4$����v>c񟍧J)����t�,9%��.��]��D6 tE�����҉���ڤG:�?;(��n�J�:k�8�&!\�w`ާa�d<״�$:Nm�.�i ��e]ob�6;�l⥴�����g�,q"3$�Ľc�flz�l$Z��@��B���6ئ���W�i�G]�iyr��b�׾c�Ѽ�/���!r'� N�LmV5.R=��� �`-��ȣ�]�J���v!��*<���ӌ&�*V�3�BcH&O��s��l�%~کngܜ���U��Ra�k]�o�w�5�
O�E���V��Ol�Ʉ���4v��г�oGm1��x�U�u��p%1��)͂�0MB*�o�����C��;d�F��Ġ�v�;�}�,=�8 ��� �ʽ:fRu�/Ⱥ�s�1����_8���On��*�ݬE�'ko��︻ A�K�W����װ���i;ȳ�Иg+��s�)�]Nݞ:��?���Ц9RHcPAgB�4͘����p�k�Z�7R�����(��C�:\Y]�g>0ٱ6f�_�٨�`��l<�K#��+��³)CD˶{���6�m��%�(\�QXX�g1[��O'>�r��q5�qv�����i#�gtE�G\%��Z+,p��ԏ� () h
AY�����f��0�7��v�GS�OO-���kǜ=00͍"��1ц�Q���z UYU����8��.��S5L��{�ou<de���Z��ɇ�\K���|���M��[�	٢�ę����U��R�r�쓳E]8R�i�{��#����s*�砲��{p����/3�Xtz<�ֿFĶ�)���\�x��>���=ة��kQ=+^ʂ^��u~��>�/�
G�o<x�+\^��w|�7��gn&��S '��[ׯ����1��:�,r�N=3<�v��1a��p�W!i	Խ_T�^aM��u�'��//~Lж~�}��3��8���x�zb��z�c�j~K/6����'n��~l�|.&%M��{�H��2mc/C�$�p��TK�y3�w׌���1���ޅ����EC�<3߈����2L=�O��G}�C�7�M�9):�k�Ƙ��7Gg*auu>%�7�~9\]�������~_�Ì�=5>�{�}!7
�a,�ֵf�����XM�7X�(2��l$rC�͜O�4��"��`qmâ�{�1�sm��Q1o�Aet�N�:�c��xb{ݘzj��.:��9eAHr���2f��s��%K6�V����{���ڃiM��� 6o@*�܁�l}�)�͵$��NO3�!曀Λ��豚�KhvU�R����R�����S�6�@��{+y����ܟ#cMR�����B�

�� �z�V�?aպ�{H�mRa��ڊ��%6�)A�R�4�F0:�o�q�^��;�k�]��&]�����4D�F�2}��d��tB	�Q,��Ji�#)��-�e︉��]�	�N{���}w�$!D�f�^W�A�}$�;�t��D�7�E1�й㥛�����O7ټ뚙��ȸu^�����!)fڝ��2��Y��'��,��SOnݪ��û\�rk�殧�Ɓ<��0�z0�c��E����r!6ҮqD1�3�Hc{�78�`�&�_����/�l��^&-?,O �����]�0��>��W���/�p���O�«@ke5�拺��u9�L�;�Z�b�^(ZF������'�q�c�!��^xa!��Z{%�Q��9\6��wf�+I�IՉ2)��4զ}k=O+���T�e�wf��-��0��or��]����hs�0윧��~}�3�V�S�ƲǱ˧շ&+�'%t)W3˄�Hz�������?���;l�`�73��`����'a��gՆ�pB1,y�#mu�&��RK��h#�7�nZ̠��Z�q8q�3r�7jY�̙�Y�A[�� t��^�FcChh]���b����pψI{ٴ-���4��Y�.]�xJ�ͷ�Mj7�4�����e�p���K�m��Fo}�5y�����y�}wz����)�H+@�!J ̄�&L!��n���3���m�~�9։ǫ����U����_��M~�c`k$w�?>Q�0�Z$�.��q�_u�5�<�L��	���^��6�v;�!�[�\L$虮|9ն�W4�v��m/y��/-S4׆�<�IN2�٭��g��pߴVП1`��F�Ԃ�=�T�X���s[}�K�1��MG�޼�j�(8�Y���Hj�Fu��l�,qL�˭�e�F]�L��}7����K�q�	<��=06��m�W�5oA	���a����%լ�����SYt���c���/uE�8f���vzv蘒�}ɷ&=�A��'����5]�,�p��u�'T�c�Ks�]�����~^��x��A�k�xIچ�p��Ls��=�*b"FOKn��t�-��"$��$�Z�*�qo�l3�-�q��{}BDw��] �c��jU�Y;՘)|�=��#�|�C|+��H�k�X^b���"��\h��.͔���dA>�}���\���uN(����k���'���N�,Ԥ�~�6Ⱥ��9��y�m.)�x�1m��	d��A��	,��(�����{���#W��m+��RM"�+Ovg�����=�U��SQ�!#�[]' �>��� /����"�Pc�#'7Wزs�5�k&\z�H=��;��3�+��q��w6�=��ٍ��:�T�/j�G�L���n��B�c�eb�O:�_M\���+ӄ���g�5n:Qʌgd��[��`�V1H�v1�7�Y�T� Ɔ-��m��>�>�;��v[�S2O����|��/�/�cxlp��-}n�2���a�����TK
����s�S�;D~����H(���dAX��mM�b��v7U=�W�a����:����̝7�MoDVb�{g�h�Y�'_�}��f��2���d`�;f�Ժ��[li�v�_5/�����N���`[���L������.bnS�Ի7����X�S����U ��N)A5�*��^j�[ΐ����:��\�1��h��Nvn��u3����D�jK }�J�d;�MD�
'-�jȡ1��5'lW
y�-uJ�;a�j�V�\Ôl]�s�t���2�B�@R7��Q�NsQU��s7���_��V�`����2���f���̀���\���f�.�J����O6p��Јs2�,�M���m�ѽZ:-@4����_B5m$��|�CKa�F\�6�)�$
V�5({�C��'��De�ul��]�h3��N0���qz/�f>�:c2�����:��g�����y�R��.��0��A,Rŝ�6��#���V�O"z�٩J��g���\`��Q��XJ��K��(X�X'u���_jR�b`WC�G�^�ײ�S�ܕ�����yl:�����F��X����#^�}�S���w]�Q��6�b�[��-M.,�I`��z"��Lb�,�-⮼�vl��.B���м���Y�&� +�qZjd���&\C��<�/���1��KA��uR�֏q!jeݛ�kD�C	fJ'zRuu���mA�ne�2�8n�7H�')�u˂Pͺ��]�NGM�Pͥ�5 w:��M�!�kS��uϣ#�}W<�Ð��QGfn{.��F	�j���Wyt�)�h+�$̐��`�����|l�ٙ�Y)'�A;a�u�&Ƭ��Bm����'�[P��6ڝn���S=��(��89r�r���L�9����Ĭ>��
�daܣf�M�Jߥ-�#�FY毂#��Ӳ�c1V�|&|H˒6ٜ(7)�v�'뺸��m�x���$3�n�
@��R����U�xEc�N����We�{��{�_��h�����M_=�=]r%kU�X�\i���&.�h�*�s�T��������r��4��0^��4�+�7��H�����2c��<�v�%Mh����C����j23��`�7y����&WT]db�y�K����R��)9�p�uW�1B����B>-,@}l�D�U^��XӶ
�9)H�u�5�M�Z&�j����Q%�NO&�cEED��堤�͒��rm���$��l�M�Q��QA���s�r�&X���L�$KMD�&��i(v5yo1���b�<���������N"��m�DǑ��Z����J&*�f�(����<�'�!���<و��@j)�<�QIT�-LUU�TST��ITMEQEA��R�P�����g��(�*h��٪)6�y�sESMͱ���

����[�j��/ �y��j��j -H���jC��˨�����3y���~=Yɫ�he}Ͻ���3Z���R�y,�d�޲�nʫ�]4�:�t�Mѵ`��n��;��{�$����^|\�<>���!�"�E�h fHf@�0�&L�s1�7[�5�f�o�Ӎטt'�����
6�aT�\��j�'��RX�:��a�����6v���=}��ʝٔ�><�}e�-�qx�u�Q.d㋰8�,-ts�쎙�&�l��:��+��`���I����?�}`:X>�4�0�ק��9���hZ��+p\�!�U(ڋԡ��{w��^̈́^��A.X�m/a��0?�G��!��"��A�[.�K�s3�)/�F���=�#��\3�,aL��AZ~�ǿr�i�&������Pg8dK��t�b�!�JU9w���Y�K�vv:�z^��d���>��k��S����":Ξ�����Jǥtg/:���S#���T�^o&��m�b��^D<��s�VoS��^E��!�(4�].�pE�~JV����7ݭ��6h�_)���.3�,Ȥ����I�j/����5�-�a�T!�k;Mix�[g3���=м�A�-Fb��>�F�_�A_�.D�`N�@1�YO��B����˱�J�Z2X�v�hfe
7�4y����	���:��hBli�0w�3O�����G��o'I?�G=�j�םE��8t|1�s�!�,���|����COnBBp��<WNȩ����4�HEl�� �%>�O�˘��?j�S5�n�<v�K������[��m��N�N�e,��t��r5|����S9�Z$�|�J���e�3#&�9��Wz��j"z Ir�0�2�0SH�@�I�P��߯^��?k�i�]��o�pD�m�!2X�J�a+�����|ioSCX��gh���I����P�0g)��1޴0�˯�	��a	Ll�NJ��6�s"���ǡ��𞅾;�,��4)��:��5�3��.�|����k�ך�k�8̢��"�s�1H�a��/�^���(T)�vk������ƾ62��1	��=1��H�Abql�e�:a�r�E�x�#���z�Sh�{�Ï5�o��]���p���� ��Dp��^���װ�
8e;��,��v���+�7���U���@f�e^]&���K���d0�t�Zc�ktlIu��6��F��B�l��3��m=�������J���s2�w?,�|���l�`g�:=í~��l&!��+�����-KaBz�[+�%X¹t�r������Ѫ�c�P<��(Q:���W��n.j�T�Z�G[���NY0���Ͳ�-�I�������>�~1 so�ۖc@ņv73����'��@͚��A�8u�;�'��;_�f�v��E��x���Šv��/�|���E��Qf�1��bZ"�3O7��sk��[��9�not�#>��3J�f[�p*���>�nu��Və��,r���x�f�暆�匱2(�+tW�w������Ŏ���/{�S�����Sz{��ʙV%Y-�VH�mh�ݏ2�����c�i�a�<��!	�@�
D�� �=���Ν�z��q��6�wm�a�A����Y|���K �A��6���S�(H<�y~�ª���Rv����ܨi���H؊�U�,�D���Ai��I�OE��ޑ�.2Ol�X���vwYf�;'�$�B��4]U�ǂ���_].?��~�!�U2O�꣍�noe��_Fv�/t3�q�@T��aD,�`Z��ڦ�����z��@t�w��ŵV��+^=�j̋��
K� ǥ
�a�e���D���)A�0?g��`_�mq��Lߋ;�|^/���VR�7��|�߁pU&�)�2 _l�(d���'�%�{�Ji�#)���Ay�{�T�^��O'��\�Ξi��Aq��;5�&
���'��K��N��"S�r��N�"�Y��\�V�Z�1�-XL��^��-O�p�<�@0�l�C6����a�`�Y��:���8�ȫ����:P�ʴ]E��yh-�a�^=]����"� ���tۢvx7d�ƒ�*���$���6C
�i��M������M ���R�>=!�Z1��0Q�~��4hRoeH�d�9�Ȋ���Z�_��]�$��j�u��3�� �Ѫ@}͇~/k3�4��n/\�|M��S�t"�L�p���ǬWWP�-�ߎ�u�Qر�.��{�.N�Ä�A�'��TFE���V�n^Z�/���:�n>�R�Y���t�ϟ9��~�O�	� 
*��)
E	�F	�h ���;�|�[,�oK�&曳��W{��BӭFW�.��a5�^L���*Q��H�ّ3�����ϫu��C�y�d�О�\�ęƠ���0��Z��yJ�Ъ��;/��LE�^d�
yV�9��Ӫ�ٱT0g�����6�/�ϗ�E$Ja�Ʋ������"������D���+ٙ���=t~t�B��(�:
�"��!��������K��t�ї~v�Ǿkփ��Xnc@8��-I�c���w��#Ds;@�����X��dk%eGn��2�u�U�v����T$������1��N����y��.�0v�o̞\�Qm�Z�]e�����eo�7�є��kL�v���F]�[�Zz�m��ȧv���C�\5R5.��H~`���sߦ�}�3bq�d$U�A�QW$1F1�Fl� ��mnU���ԉz���gz3��r�=;��`d���"1邿Me���jzO�`� ����
��Y�YS�	M�goB�t���Pʋ�4=p���X�.2���.�d����_��ƒ�|���}i���#'�8�hZ���u�&9��%g�to��8#�<l5�+wJ�.��w���oOB0i_m�{�GB;�"}"�h�7��f��\�}ΰ�)�暷w�_6��Pv2T�T~��slC���T�����k(�nN]����] �$�DдKIH�@ĥ{�������_oW��Q���z�(RXKjܜn��u��D�Y��v��.��$�5s6���l?N�n���\G7sو���R�j��E8���a>�hTN7���!�o3�M
lu�v3�]&�ݭk�{!`n^��dɇl�J�,/1V9�QzK�qӅ���o'�2�c鬪�3�tO]�6M-�e�^��_�L��`K*ʧi����yE2.�x��e��u^�ϓ��n
��wAy��s���!F�?�`��`` ���7s��E��'A�L*��熫W)<�RX��Y�%Q�ǫ���kn�Mw:����!��(@}e�LlD�=OEs����e�q[�*�7���E�2i%]�|Z�g�6�5J�������<{\0gA��X>�4�0��@��ƅ����L5NRe����{�R�V�NK�PK�]�y�Pw8�<̆�5�93�R�I��t,���|��.�P΢�6$���5�|��v�5-�^=���pȗx����{�5�M�ݛ)���X����~�.ȹ��v�r�
bK�qdv�mm=�������?*�gԽ� *}.6:��[����;a��>4sg��5�<�p�\[��4��i��.�:�efԍ��X������*6�ɥ=폻N��JcMr�9�]��&O���T4p��[�i{��������o`JTՎ�v���w�ں��.�L�	�lCW��}�X�(V$h�J)}���3 � '{��+wY��8l	��ݡ>0�F���z����9�A!��7�y���f�&F�E�����������%����t	A����ؚ�Ƕ�3as�̈́��P�٬v9F���s�(_�"����l���Z*��7,������+��%ȟ�	�S�1���P�F<�Y��B��6�gGT�(Q��󇡽8�E�U�`حa,΃�Ʊ�cZD8�vY�����
�g��YY't�U�Z�=s0��"So(	��"K�%v� �-����u(���W�=����1:�]�U��&BNW�k��:���ħ%B`��*��d�=}Ǆ����7ʹ��.���5�T�pm��B^��@"o�zF�����YY�x�4F��uq�z:n��W���'˘O@s�HN͎����!�{�*�f���1I���R��̦�"�4^e�v�-K٦���w�pw����vll�����7�7b���(�QQ�$+��Y��y��_q�u�ز�%��a��p��}����6����S�E�y��4p�22�]�+b��y����*�O�b�`=Å��W��� ��Ky�t
B�p�n�{E}� �h�mg�%��Y�kr��o�k+��:�Ն�XBG3uW#���������R��F��;-�Lt��Nna���6k@ݹ����aHɁ��5ww� �)�H�iF%9�߶����ɕ���6��F���s7J�s���@��@G02ã�\��\��!�o0��sہd��;4�X�I���J��]+^�PKܽ�Q�*�Y��-��@`�VF��1]vY[��t4F�ϡ�9i���mǡ����T�ߙdк~?6����w��N��C��b�W�p�W+튠3?�d�!�Cξ��t�C6C�Ⱦ�_��IC�@���J�f,D³W�͕���|�l���v<��ˎ�Se�N�k��C����
^Q��շ���f�M�U�^�hO�=PŴS���T?VD��BH!��!�z�x�r�+P[�L�Nu�"�f�P��ݖi^�����B�L8{Ȥ�9��F��ǬG4��&��ٕ�^k�.��H��Yv6t�Z�~SS�ǡ{3�@.J���A�yd����3g�C��WH�~���Ǻ���F��w��`�S!�����)Uc��Q^��D��P�&VbK�]:Fc�J�?�����]��t��,(}w��@�"X,�mPH==#E{%W5tB	�'�E�=�/����#o��ɠ������4��ׯ��U)�d�j/��zj�L�i�8}y�;9C)�}�8���=v���I�Lw�r�x�"x(GCՓ��u�����]]q��\{Y30���ᰨ��k0�8�s�\0��0���Ɑb��*��ifqȄ�a ɂ�I�T�B����]�����{�{������毄�|>r�Οm���'�]�*^B�H"E����	�u���mn���e��l��F���L�i5����S�\:�ty��a��D%,�Bvx2��Y�Ps�Y�a�T� �v��E�*�5��1���F��0�х����� �� r!6�i��]77T�**nnÑk{a`n^��e�g�&]��&�z���'�K��ZG.����z��[2�r͋�W7	V�K������O�ĲObz曬gֻe��kz*;�6;��b]�Vr�e����V�ޗ5x���.������yG@�u�dS�Vצ}b16�����S��/P���B{�<��/�|�
�wf�@P��!�a#��^a�]�$����BՀ�S��5�9H>�.�ҳh�5��;Y�+�Qo8��A��� �|����W��P��G��Q�vgz�p�{g�+n��t7e���8���
���s�n[K�w��4G3�
<:�$B
d_!Q�4��Wv����#��uO"�ޱWFh�P�.Ť$e�m��ȗx�A�6�������P�*�����&�Q�yf�
=QIX�u�vB5���}����j��g;g��)ټ%`���&�q�6�;GJvI^��\;�e.�M������9�2,�t�7]V:S��e�]o��@7�ٍ�2�<i�O�~�T7l�|7�f.�nj��>ʞ ~���`< f 3{���f  �����7�D���&1>ܩ��~��>�yf�����d���F]�
������1��1�l��U�n�9	wD<!0���%�j==�͊֯��ǚ��Z����
3��!T�]�ʕp�&�>i���e,P0-�9iw�^������¼"[� �QV�s��[���Ǡ��V�ˬ�Wy�[JVֳю�ƯeEê��fA8�"K����i]:ɲs����l��CT��TC�pe8�ۯ���PZ�R�TX_���:�uW�!��J�]	xI�z��q�ٻ1�$����o�
�-�^��=��NJR)TS�����M:q� H5�g�4��g4k!Y��Ö(�� ʽfY�k�ٽJ�,�x	��y].2	Ӆٲ�V�΄�h:zm9�v�t_k �F4à�G@ ��a�,�*���JO<��H�e��5��ݠòre9�J�k�}~h���GJ��*��G�ݐn��=��n��0�es�U���v<6��X�#�Lѽ�������vsB�	 m�K
4pk%_�x�OEs��t,ۙ8��X�y+�i���e����!�vv��7w����(	P���C��Bț�c�15Z��9����%�K�FN�{0|��$	G00':���X�Լe����ΝH)["�}�N�&���ܬR�(��D̳/�H���v�
c�S
&���/��������h((�@)Ws���}����;���������6K)�R�`��>�{p���O�}n���>�a1�'�smF�Ҝ\�=+�l���Y�A�N86ǥk׊�^ت�	�'Z�=�~�("����s�zM��nӗ���En�z��i�zv]�ΔÛ��@��6��P�9@���<���/a���2k'�-3���;��u��!��FC��'z]�}�(���$�W�˷c߬5P��/ʥAJ]���\�F<�ɼ�_>�x��M�e���/<W�R|aB6�ާa�,��0	�@A�غ�eph���&�����.��D[�Os`3`."@B,����ؚ�Ƕ�3cY2��Ul�~�Ų�F=�]o���te�#�e�y��)�P鋇T:)�0Aa��8��ue�ME�p]@��y�X�wH�� �����L�糰�%�"N�G�8�¡���M�8&n�5hMj��M2�Xt�]���e�6�[��M�/��	����<Ԟ�vM=�x�o4���귦b�r��Z)[-q(9�0��/��W����x���R�m�g|oJ19����d��$��eYE�������}����T �]���y���v�"���a	W'|�=bӫX�ۢoj��e�fj�5 a��oC6�n�J�ݩ{;��`c9]�W�>Kq۵8S�D��R����j$s���wY7+ahD�_VC�9Hqx�iPݷ�/�%���U�X�!2�k�/���_D�h�3�j�fEσ�Zw�.�rj������-�]�"�Ww�[�2bnV�f�wYG��,��6K5�z*�2�P��j_v�1ɳv���Ώ���n�,W-a�Y:A���.[��C��p�]��H��[�t]�8O�M��Ի�.�
��H�ɖ��іj�4k)�"�pF֜�w��.�Ż��U�)Ϯ��H�#��4����3��ۖ-�"��w���N[��6ͺ��c
ފk�,���`83�E�6��i��ݬrӒ�SX��&���^�Tq�94򽲸�
�B��xf����5��2�W\��^=�ڷ)��<u�b�3]'A8]tM�#l٨.�Tؼ�bQ��Sv�=3s
���.B��f�so�Ow����;#l���h��bv:�,��
yF�\� n�)fn*���Jn�{ݰ��i������~B��=��u{|N*{Y�N�u^�}֬������l�i�ܭ�7��c%q�W���]>\��e�5���Mt�B6@��8�*r�)��ϴ*�:�6�)"Q�;��,�K�ڳ�K�v�p�Jɐͭ�ƀ!�d�"d�SL/���׆�N��h�0XM>1�$�-񽤠�um-��lRt~F�1�^n�3��cx+-U%�	����<�1��Σ��>�.�+�w8���5�u�����&�'z��ܶS�hu�l(�{p<�4{�ٙǬL��ԯ��s�77jXn�ϳ�@W)uΩc}�
��|JD�����k��t��˺v�M2-���l]�k��ӷFb|�EQ�|��^b�4A��qBw���ztT)�ܡ{�\����h�a�}}��g�!T�܁��d��?��'\�];r�A'G�W1H���&=咢�w&��U�u,nlwի}u�.1���Iݗ�˽	�2:bT�/o*���m�U�ġ�e��:V�*�����V�qv�)擶vQ=�oP.[[[�>h��VB�d���8�6��JZڥ���8��wj%1��+��C|j5�m��*�`L�5+w���f$�Nt ����|n��`�n�>���%`Yk�	y���m'X�;L��Ot�[܌��k���>�ie�h�槼ut��7g$�jV�4�8dF�J�]�.�u���/b�쳘X�汑Z�����< �׻��.�}x ;h$���_h�H�2���1a[y���۔�
��/7���ř�ԛ�]s2����E5��%b��^�
��N�]���Wj�t��o���=Z�`���� �,�<�49�*��(��]lŕoc&����۠�J�Kۯ�SIBD�5?�$"��LUO,ACUKBQ$@P�L_6��6SI�����TD�d)*H
F��@fJR�B-hZ4�bh������'T�4MU4Mù��\�G1�����$|���	����\Ψ
v��4�m�cUK��(�43@U�JPQA�bv�;��+��Ѡ��D<�4�4D�Vq�
]�4DD֝5E	@h4��Dh4Ě�PA43<�PE��ҵˑ�d�W,�79p�&آ��A��s���j������1$N�"|��r�D�5A�Ss:@��/���(��C�'���2hsv3X�M�ߟ-�����Z�
� Z����5�d�U܉����i�%+�N!�����4�5"�Ht
��5_W� ����0��x:�U��\��Ŀ���!��d����!=�pEq�i�I��d]g<S,��O��.疭����ι�sָOw0��z�CH.͖B`��9��p���'y����5�3e�uR�§;�n����*L�B:}���BhiF���li���zBcXn���ɚX�Pk�w;�2Vӝ�]ů_0��1j���T4�L?5y8�u���=�d��#[��WM�S�����~��1o�vm�j	�c��V���ߩP�u�9���a�$H!��ּ��ɸnѶ{��I�}#�/8{O��3L���&�W	V0�r�Z�
�^��R��=�,�C��?SR�	�y��ڥ�����^|с�z���#D7c��3lo�ʓ�����<L��yz����?���SG|�X�ͫb�;t�������y��|/f�v�ҋ���zHvј��ǧM,܃s{��L�دn��-��C��.������^1�-��Ad�rf��ŕ��,�s�%�_x:��'��
n�T?P�Y��Aii��C�$��������jڻ�|DT�`f"�K`���*�3ݵkn,��.��#(�n�čJ�yc�]��*Ku��}�v��`�s��ˇo��\��x�*�$U')�yY�f��Yx�쌩ǗY��%@�w|C=G_`�>ƪ��#oxq��,,�3��b_0�헻5W:²j5\�9d�F�ŐԆ-��|�>�C�|3p�4о�é+��0a����z�o����Y��]�Ȇ�u�f��ҵ�g/�����K��[.*Y�a�PY6����z͜OC��+���Ee��K!��	w@��2/qq��^UX�+ڊ���7��əc�.����a�ٲݬ6̚��)���1�u�z���6��v^�gDK�+�A
y��A8�Q,��֬��i��Һ7bk��O?^��jBV�k���Ʈ{g/Mn��J�.͕�/	��_	H�K�t֤�f:̷l#�����%��LR2���nO5y�.W�<��kgJ�'g�.;�3C��S����Vg���L×���� �I��NVyV�0���/O���a�<��2�tq"�]�;�`�L\�a�j��P��a7C�(���@%��Ժi��4u���P]�hv�39uq���	�g��:	��6%�=�\�u��Z�c��V�kzGs�O�㻞l�s��P���o�.�����������v�n�����D;'�;�uޚ�Lk�M[^�I��#&�k���&��;;���'.����$��]�_2�ڹz���Ӯ��8�q�.���򦔛��~���x��u�Jat�u{()Zoj�]r2�G�00w -�hɈv��K%KN�!���]S.�t]������V��Pu����"3r��Q���5tɥ�-��0&d�qd'�9K�{�jY��a�!�ga���@A���nt�D�r�C
�jéL94>T�=r��J'/!�;�Ij/xcӈI���a��۹�6�������v>�nr_����^A���v�Ph�
��8��^y���c���w����*���Ư�g�k�����z���_��?<�Ρ48�j�v- �ԸF'��o
�D���97���W\	�}�m�ݷ�����	e��	9�#�m��{��f�d����U�a�r2�m�I��<�/]��R9�}|f�9�&�=a/��.W�bq|�Vi��?�l$U�A�PCi샓\�k(m���
��Jm�8�t��zw�NI�1���&���B�!?2������?U�q
X���,�~��Xu�+K��#�*��
͈�q���i�Y3jf�v
q�۴V*�ڽh��]��WCv���Z�B��TXSW���W�����g�L]�A�kƼ�jE�[���V�S���n����%�	�%�P��=�b%9��Z�%8�K^
uج/��������}�%���,W�ǳ z#��묪�^�Eߗ>��n?s���������J����2�.� f�;J�u�@7B�:���I��7��.�(�f�ΉG����jdGP��Qo�"������	��j[�,��Q���z���C�x` 15�*s3�$�C����xf!�/���i�I�g�C�E���78]�B�ͅ��k"��Cwu�x`���"1�C���	��0��T,�v�5)<߹M�.���a�8��$�Uzu�g����M�~g�=�����)��@�r(��L*���w�,�t�Y5�]�Q�gj�y��܂;P�Bxwf��|yd0t�" &��=ήMг\gFt0W���n��Wyo8Ŝ�0�k��͊U�'�=�}j�����9�����>&+6f�1	��tA͑�:Mm��P�4-X�N)c��W+^�PK�B~a�m	�����?�G��0S@R�9\$/s�Z�B�}��tgRa�C
T��v��i�Է5�0� ^�9�g��EN������u����p����V������ۧ����7���3��6F��*�.���c���s��l���t���u=C�>0�ۜdw��p�d<�� ������cYO��W���3/H��.Ӹ"۫�m����B,��̔��5�mc65�޿?�BO�ff��ǈ���Nx+�ћ�WX�934V�G8U���sޤ���;�Z��⦗���S󉡡�0͹��]�V�eB��V��a�K6�b��IWA�lb�f�'ėt;&uG�t��#�} �D�Xp�}(g:}EE]��v�Ȧ�&��w7p��e��o<|>ox���[7B
F��M�f�	�T;��M�S�������,:N&.拹�_����d}�0�s�[Cj����!p�o҃"�hVZTy��ޜap���ĳǐ��ֶ��X��uwko"���!!;H�8گj����%0|�&T�P��$Q��~�=[�Wk���h��T�l�=�b��4���	�����>�S�΄&<x���R�&�!B׽z�[�<����i���l�(�#�1ᩭ���!�ļ�z�p�[���t�.p�nc�jHbɟ9���������>�-+�U&��+�w0�����H0͓�.z��%ˌ"D��I�9oT,�;�[ug1�5_-��wS����1��d~�.��
lў���@�b8Bn�OHLWOu�n�������zF0�w^����='��U�K0a��8�`>��CM�v\��w��{T��z��`�j��N�J�`Z���w�Q��j;�͊T;��Y�|Ӈ����^&x�ڡ;�밹�С���c�7;4��Қ�%�r�Z�9DO)��]w��??ޘ��~�o#�4��Ճ���CTx�= �K���R��&�fvr/�f���5��78̧�5�%�"�μ�[s gJ��go((wZ�b2_vS�3�;R��nBAz�����7�����8Gm�r��,c�2��34b����QY�ej�D�eb0r���#Wr��R���L>�H`ϣ�<yIݛ]5�C��׬oM��*�eO��r�N>��b�L�6��7ݍ}Y�ҭ�&�R��d������ξ�Nç��l�m�}(�te��c=[i��&�����vo<�lZ��;�xA�����f[�l��;����m&s+j�l��din���A���,!�wB!�@"|	ꆐ_E���a���Aid1�S���X��e�oZ휷�zޡО�Ok4����,�+�O����W��E��z�xi�έ]�3f�v���t�x"ŗ�0�}���~����Έ��䩛��eT�m�d�H}͜OFz�q1㙽���F�w8�6�z���ŴxXt^D\zxR��	Xڊ��)��)A�R�4�{/.+$ �jb^gj�J�z�CzT�D�cз�x/V��$,.b!�v�"��+��t��T�Jح����?o-�c�ݨ�S���L�J4��Dn>753��{w� ��Q%ٲ���A��ʖ��9d�����Y��\D��>�NoڤSH�kc��i�h���4�������������U��$u�y�׶.�M��wM#����k��~2!r��f@7K�K{��Xz�	��N]��U?������OW}�m��n�
Ή!͂��CR��Qp%��M+w �"m���	ۚ�_VT[�۫Ӯ���2�su�p�;&���������T���v�������g�f��4�.��PR��F�W0�z0�a���>0����q
��L����S�v�!��	2�*ΛjOxT�Yt���>��A��� �Fi�ǹEK6���z��R�N^R��c�5�q"6%�=��n�S�Vas���Q����E��7����:�%W'w��w���@�6B����vOƧ�W:�I�LhA5mza'��n�t�ͱh����.��͕�l_X��V06�5Z�۠�C���6�/ﯜq�j���
{�V։�u�;9s	E�S-|�F}[o�'���JDwBm��tg���ާ��5V����OnW��T1U�(*�a���;(��n�r1���;��E�ip!j�����'������Z����
�'���}�:���4]��eش���q'DYz�m��Ů)�-kDR�m߳��t=��4
1�&s�N{z}�i�kL�v��� ܌;<�X���4��먣{����h����tO��|`���ϣ}Qs���Z��H8�fi/�oM�;�3�3V�в��Jh��v6��ƒgTm�׿b��C�+�l+�ޮ�ɓ%�z�u�;%�ZT2cџ����;���9lva�W�+/+a�+#׋���tǫYD�%�n���=pہn�L����U�w�����]0�ٚ!�f��}�^�<��S��������&z��?�,#$�!��<\n^m�nt'U�en�'59�\"5�ێ	�d	cA.�g�c���Qp��3 �V�b$���<�tƂg�z�\��J��ݮ3���z �Z�9E+�,R�R�TXSP[��C�.[�>H��CK�[��75�n.NF��ʤ͐�K� �"�S�tBd������T-\�E8���;�L�l-�"���!��W}[�}ƫ�<�"%���#`�4/��w�]��iRe�/1V9�QzK��)����_RZ$��͕T�;�0����0�'��i�0%�YT��fe'��)�E�N�L�۽:#<��w��#����JOc;�,@Eh!�בCw<s�s�MУ`�&eQ��Oq.�^�k����U����.˝O7䤱�v����vh���`���M��6��y�^z�����ʞ��$�9��.�����c6)V���.��_=�~��rѡ��]���ʹ>�c�l=�-Kj�*�ĨZe
�w2��-r������~���=�P����w��'Eư{��1T�7�'��ۧ�^T<� ��bZ�f�&�ѹ=�Lk׷�s|"�񱖶�Ri��%�<�U�䦹�v"{�kC�Ӭ6{^j��e d��.�b�+-�5/lnf=�Kʾ����9T�v�a�HΛ�y�ëuق�zd :/�'e۷:SnR�m�Mc���r�5-�@�/}uxy�Ι�c���z?j~�}�
9��&ǸdA�
x����쓭�v���Ë�v��]��(���J�]ƭ�P���e@��r�.���:��>0�s������!�/XiAU݇P�h0{P�� �����-�<S���fp0(E��̔�%���x�1Fkm[fknJ��:��嗯��z+��&|�댁P���X� ��a�q�� ���oZgj��Z��U��ӈeT�5 �H\�]G�2�������;>Ҩ�!����?
or��8�h��Hh�-0��i[8��کnj�6��!2��Ty�=��g�1�"�b詺k�ѹ�KNh���������Ŵ���L��W�i�y�t!)���Js~*Sx&ь�'D�~��-��7U��v�>�HGNc�s�yOx��C�d���|��o��N���n-ٚ���yEb�x&���Ok��L��I�k�8ǻ�O���3d���s�9l���谸f��g,o!7-���WYm��������	��d�|��*:ś��2]fKe�[�9�[�@�"���*F\��c�Ֆ�b��h�����"��e�J⮒��7r:�2L9ٻV��s��Y�f2N�-&T��PY��{L[�8LYۇf�嵣���Ldw��?}�7�]w��X9���v�1��p��=2	ٲ��V~��wN���@�������&�{t)X�E�U*������
�.]r���?�7�u
�Jױg0���?l,=[�/��53�rּ$�'Pb��0��v8�0��Q��o砲4������k��ʐ�ң<i��F�4=��dz�Z�������N���ҵ�%�^�G6=0���1���e��[�Ι��`�*C��/"��O�!�q�׽6��LB~���������7�����yze�dεvܳ�������y���v?P͐��EeGC�s)��Us���7˭�7G���Zex��L[ ��y��
,#C�q>�Se�E��iD�=�������ƕV3d:�6��4�C�����>/���툨~ǆ{-,�7e�		2*^���ʬ:%k(|e�R���oP�3p�4���@%t�#&<�M���6�մɷ�ۢ2#w�{m߲����ZZD��3�争�G>���P\�3vA�&�H��(0l��(��$��(��
��񦦸)g����,Yl_�i�d�*l��e��ѷz����U�﷪���ӓ��̹�7��d���w�"5%k^\��V#�
���X��TQ 'O�JO#��&\{M�+&$NgJ];[��̒����6/jgV��cC;��H��c�:�U��"S��4����S:ؚ*v(FI��5��e;����hN�n�=B�!%�L�������֙�D4�ɝ��<��kTV�BP�mV��N���C]T��%�ɨ]m\��1�ۢ��.Z����ޓ�zx����M\vU�uc�}��J\�tp"I5!Ǒ\����lp�t�%�Y��\�!j����뻑O�$̼��k�m��]kޙX�Z,��mbd�W�b���~��/�wed0E�Iڻ�@Wk�7G&����W3w���ui�8k��Җ��횪���C�e�r��%)L\2�LcTI��ݴ�%��j�W1]�*�3��å�R)��y6)r�g8�:�Kw���/��9 &�5�\�]����� �fʷ�kTՅ�k�TD�g7��&e
/k��o��cQt�{�]17.�ajO����ش��Һ�J��@���f{�Mr�d�n�SW6�u����	�V`W��}�-ZKN=�{�Q#)����ɴ�;ӇP�4'	�1��w���c��	qKWv�������7�Š�vQ	2����IX���A���ȸI���VWt,eg�y˳b�k�|i�gi17k�H����G�{�]���Z]�u��t� ߡ���-*^��b�OOL�G���C��P�ק7�NT��"]
��e'W3 �E��b�o!D5.�F��'[���m��y�pX���4)u|w\�݊�)���� $m�����躹+���3^sC6	��<�(�҃����.�}��\�����Y�.J��g:Xٸ!�m�3%��6䋿�9Od���v�j�+�_]Л�EP^(�~��jͫ��\p���<����l9@��a��=�u5\�h*�7��h4ܽ��tv.�ةJi�5��n���S!�][>qɦ��@�4!xFV��L�����-zr�Q#�)��iEs��/��}]\�;�9����HF�:�[L���|Wg^�͌nu˚᭦������������s�N�5��i:�7Q��2}Ku�����C���w�w46���o;<��,��Ekٵ�Ꭰ�ɜ/0^��Ө�^����]��틖i\i��rY�5V���/W�u{䬶��x�k_:�Q��-0V���jTCht1�%�G�j��gd����q����Q�7��tB�@V�r�� CCA0t���Ȋiu��V�	%,:j?�p��8�ei�E��	ͭwX�fT�p|�5zވV��Hi�W�&I!��,�vӻ�຾�������P��W���^Xo���6
�YЮl]��1�VoJ����\pk�(���Awc�ڝ�8m����<�i��5��
9-�9���A���4i�-r�I����T��P�E4�P�����-Pr����E�I�伌I��� )��kZSF��I���%�kI�SA��''�E��m��>K�Q��4U�Ʈp��gF���6����-�Q���%W �\6M4��9H��M�N��N�&J�EAlء4��ƚP��4@PZ���h��LN�(�����l�ɥ)��f�^l�퓕�D�
C�:���)���V�(�)���l�E>O�Q�o��i<Cx�=��J�z�ķ��I�5l��V5���a�cRٵ7�l%�3��^�H5e�َ���W�.g.��]��K:3�(���B��A�y�dzp)��8K���#x�M�9J�Nvٲ�K3��G3w���Gfu��R�m�����.&��?X�0Z�	��.�W�UsS�jچ�:�WS�s�٨�p�y�=���+��I���|j�(�+�a6��b�x�c�#�~nC�e|����zY�t�~w��?x�JscT�cIMl�qͯ�p�G��kf����;^rp����;*�4��A�f�'p}��$�b)9Y�"���9�#:�������;���M�f,S}�;"=�&U;<�gM�'��K�ۦ�����)���@��t4sӦR��y5�Q���T�Uǃ���[,kL:�@��e�Q-��q��2��zԍcX7�vKr�˅�n�������i׋�pd(�v�:1��6y���;'�Bz�s�dS�k��j੡o�2F�g��{�����������H�ɪ�^�@�z��z��h�?�e>G���?p�͑BQ���Ė̓�(INe��T�.�Vܘ�j/��!ݺ����C�9��y����P�.�	�p矼F��E\����K�ɼ��d a*\�I�HL�+�]����^d}w�[d�ش\���tq��̲�e�&�cJ���d�
��J�Z�S�!7by����;#��N8��ЮV��<�������t�(���P��0t��73���g�s	/]��kT�ޝ�N��ʄu{$��bXqgd��j/��x��q��ގy�UD�[nsB�vC�G4�		�Y�s�Nm
�F{�����Y��`�^u��Fͅ9�7����\�Swػ���9�.�0v���i���GE�Ӝ��z��3N�<�[в��s�&�6D���	�'ֲ�^m��	w�ϐ�a��E�j==��ZԶ.v�c����[��Vr���2䆢L�=ٶU�l���޽`���IݳX\M�&;�2�)u5;�z@�팎��L�f����YX�K�Y��/lk^�d:�����,D��R��w�핹��o��f���l�&�~���2׾QI��"T��VX[W�̜n��u��►���<>aj�u�yFft�V��l)f5/��!؍��ŨtBd��1��J��RS����49��K�>J�k��մb8ޏHB1��.6eW��CM�iiRdY�b�<�.�۝X�pF��[����y�Pg�e<0kܑ!�B~������eS�٩I�|�b�5��rW�&M�6��l�0m��Nie��W	;I1ҫ�9]�?LĈ c�N3��teY��A1dLӺz�QT��Õl��,rM]��B!����	�����Y+�Esk����ތi�N.�k'm���p����j��X�2�ĳ��+yS�cF���m��Ɵs��Tgi����]l���O"��F���������엺pbǈt�u�欅շ܋���VnRy�T�(��	�ݚd>;��`�bn/pJ�bj&�k���uc��l(��ʑE�:߼֌�,-t70s0�'�<��C��<k��>�f�j[�-jd���Wk_`8��@��fʓ!6�q�j�J�B��eI/��������A߳t�DЉQ���=u�0CDx��=�cZ=�~�;.ǳ����)P6˦��;N0���V�O�W�d��Q��B5׹�3�"]� `<�C�m�FC�N����sCV�`S�vSїιX����Fx���xG��'-�~�������>#�<���ۜdsz��̱�A>ҍ�yW�o���B�G��drA'��8���p=2Ή��5���2�Yp����j-B�ܵZ1o����¾|e]׏�<�s��BW!
Dך@���BkꌇTb���#X>ZqD���ǅY[s}gB��B٭{��j7�R����ȊX��E):��oLc���T9�?�
���W��J���Qʂ(3�#��<�������lL#J�T{k6���-غ�i?�������Nܽ�BמC���oR��e�1�۔�+R������@%7{K���m0c������m:vZ��Ŗ6S)�3��N���Co�!��~X=��l>�g�M$L�C��ig+��KsWA�o��ʖ*�d��MS/	0٨nj��+Y�۷:v9�b��B��{kN%�p����"�O7:��x��=�"�eD��K�+2:�i�o+�8���E(՘_���	��"�<~�hx~�YN�x�U�+2����_����JG_V�K�<S�F�׮q�w0����H0͓��sО�%�_6��q��B�z�/�<���/�������E��b}�ӱ��5y�6�y��@AC66Z�g�L�%B��j	3���+iS�*n�2��'��]i�?7qN%2��0�ԜK��v��s����m[����ԣN��EЏ�J`���"�&4'f��1Ln�/��}j;�͊T;����}�۲��o[a���ʜ:����a��@p�_�vi�X��[d%Z|ỡc�A/r���H��K%Y��{����R��[�!�8���.���2����W�*��G���A����Q�+6}8���v嘿��l3��n������ߣ̻��˦rv��kT��l�v��4���&��`v���^��y,�em17���PqM��Մq������j0.��h!�'NL�x���3nQ��^=X�M ̎�X&��2ĳ�D�����o��[&j���wǱcٹ�t���;Ϗ��yw�Q�:���e��)��Ϩ��Yh�	����b���GD��Ņh|.;8�7�rgx(=�����5�+�h9��X�F�$=xqhH�;�<tC�۷g���'�ePv��2�ҷm�"Ő �gkd_'���`��(sNnf��,
U �2a����|�愍�n>J��7ϙ�m�<����҂��##)͎���O����n�'ԃ=,�`Z멊O��k�w�9=1[���l�A)F��{����)���E�Eǧ���	pڊ��%6�+(6�*��D���6�j���ٛ4^F0�ј��o�|w��`�as	!v�#{vTT��W5��6v���d. �pK�"�
SL�ҍ&���|j�ΞE=������>�I���_hT��ݛ�ԁ޸X��+2K׺"S��D�7�E1H�jn�nO3c�:Ώ0��s�����ٌZ(�C=�3je40�0SfS��*R~"����F��0�х�k+ak,ٱ�u�*����l#��G�0BSttǆ����J]���=r�O�s^𿾬�}�O�F��+9�iݲ�4��[��~�-�<�V���gp_�E��(��|��e?o)NN�
�aZ��v����{B I�N�xf^��/%Έw��I��!�rq<�<ЙYb�B�kE��8�	:�m�B^�M�`�O���g�Es��w��������L'Ǡ?K�
X(�v!���\�'�i��r�k��W5[nI�U���Lo^j�3����k��#�x�"�}��W1G�ݙ?�Ό��.o��t�j�9ڸ�#3�ߜob楝)?6#��\� UR͔6-ݛga���A�ݛ]���̱f�*��}�|:Ϧ��ۛޑE:�é�k,{�.�Vܘ�jXF�P��.�@L���K�{	��ݟi��xw�Ԓ����ژ�*>��U-=i'�#4qi���i~娽���OdI�\c���#M��b�N��U�nyui߶�3A�]�s;f^8E�5�
y*V��mut�%�\�E�y������F��i&
usӍ��z=WFY���<�z�V]�y�53��K��_i��/�ʜ_�T7��b����yB̹_���ϫ�6+Zwo\§�fSó����^�����H��z͛e^�Ξy��,��|1����ǻj7K�_u��ʊƢ@��Y�A��Lu.�g/���2������A@���FsQ���d� e�� ?�J�^����������
{H]�dH'=���\�Ov���%���R[\����$1e{�g�!���|�֝��r�&f�;^��b��xMe�u��{0��M2�sd؎��1�5���KNS��;��u_]l�V	�|�-���s꿿o����[��L.z�k�(��֪�J���a?n<��z×8
�w]M����r�t�ރY��/��r]�_Ab��	�r�	��Z�%8����(�P���y�A�}e���T�oG��#a�\�Y�},�4��.�4Ҥ�x	����,�ۛ:��\��/���Y��78^���n8��i�'��ц��YT�V��%�2�1�l�b-W؎���6�:��9����f������!��B��>�.���_�����7�p�=פa^;I�U�\��j�'�Ib��0���� vC�Ϝ>6��tfb����l�-���r�ƭxǒ�J�l9��.�E�Z��3t�X&�o3����<k�a��5��l�Hun�i��[L�t���T-_�J�a�JװT��*9����CpL�_�佧\#����ܫ�y���sBv]���XsV��&�}��;����ٱfj�ki��]8{�5����3�D�Ǹ!5y�d�<��/��;�e������Sw�ɕW��(�ukɓ���~��*�l�{e�ey�2no6��h]\���w��u0m[��+&���5�3�.����=:�M�ʫ\$Yڷ����D�
�Q�U�����N/mN-]�����"�Y�0T�ٴ�(�ni*t��%�bF;�˜���ݴ��c�����W&G���.����M	9U���K%W���h�/"S�?��nq��PT��(�6���}]��!]��t�C�Pi�]��Y�463��B,��i�݄cgh���U��ٽ�p��ME����:5��2-W�E{���PZk�"�)�WL\:�tS:b��"إ��GU��hE���B�� N�ϱ�YO�w���{mT�(QJN�~zq��ݛ��Z���6Ôb��Ä&Ɯ�G;H[8�_��[���u�Rn�2+
N�LS�W�s����lv�{yg��0�p��~���H|��>!��kk�	�3�/�8��[�%VF+��ߪB��^�T.�'1�k�<'�|w�Hqm	��%����| r����9���u�7����<���K"�9��F�׮q���׵��A�lwL=�y�)��D��D_ol,�_	��w�Y�N�_*�]g����v�1���?D�p�nA�����mWU�t=��i�����&Be��I�a��*ʞ��Qi������`��)+��Q�?�~��Y�>vD��!�M�RX���P7/��*�����Z�o�S�(I��
ްv��E�/0����7YO�̊Uuڢ<�z�����̣�g���u�`�f,+���Xۇ�l��+��h����N5e��1�W9h,�mX�[ɗ��!{ϭ���w��|����cH�#YT��ubL���'(]��Q����O;��J�s��o�5���H浞��5̅2/N; 8�Dk!�G�8u��'f�U�Qkd�c]]���g��^
rk3M��7�V��9o�isT(O��Q�G�o�F���ۏ@^��*��֙BO}k[����Սi�>X&}8���g��ܳ1a������!�y���z6��]�����۔9�۔=�!�H�$�Xc��Šv��:"ص��y�a� �P��m�(#h�lU�hY��rW=ʌ�'��'6���-Z`��ᅠ ��b�)�{P���8EJS��3kM��q�t8Aib�d=�/S�x�s��9�73M�,:���B���p�./-��]d>]W%F�5��E��y�,F����4���s~����ٜj�����&Pe�[3��u+�F�6�yk
e��������M<-�N��a�w��p�U��y��=l��&���T�o�k6x2e�%?J��z3��[�z��;ǐP3�w��7�/W�fb�%¿,���Ʌ_弟%DIǙ|������e*�&��׬fl�'��C�:P�r�3��	jY�;2p�}6��]j�Y؟)Aq�(r�k
��f8�W#���+���C8s����tw[���jz'_ok�$D�̿�d�ֵx���Y�R�er�&�[����t�On����t�	ŝcڻ�������vv~�@���*�$7ҋ�_��'��D�7�O����Mmq�<�"������o:��yWv*'���{��l��!��1jY��d�8a�-�)�N�T�ሤ�`�F���eԹ�߿0-�ڛ�'.}(�O=������[A�:�cc�v�M��aR�l�S�(������hȅ�;Yo'��N�qi@��	=��l�Q�0�s���e�Q-��q�(�r�iE�*�ō��oQ��{ ����Gs��븹�wn|gaA���y쟍OP�u�����w�G4eI�"�q�k��S�b0i䫟/Hj�f��Ż�l�0g?0��_#���z�M�f�uF���M�:�Ӱ��{
�j��S��6���G�8zLW5x����c��X��I�$��C!]�v^��е�p�ki�M����|�F�4���a�Ze�^/���q�b�~OG]��\�;�ggC�[;B
O�ac����A���s�Mq�.��]�w���$��&͔QD�QEl��	�ޚ�o�c��O8maW���x�_7s���<@�5.�13y�щ��Β�l�m��(49n���˖PXsT��*�SFa*�+{V\MɌ4��Y���U�B�X2�1`ԉ	������gc )��s1BhcR�l���Z�x�A��!���;d�����S2��Rc�veF9u�M��*��6��R["��q{Ԣ�uw��s����	�o��@佱|�6+D����.	���0eE����Br5�f�p�N�H�{�fZ�^^@r�xh=<�f�J��SĒ�Uj��X��us.���VPZ5;�Q4�(��ՠ-3\�׵�G4��'a^YX���,��1�%2�Q�$���7�,Q�8:wL%r,��s�Z�R��T�2�ڍ�.��'[��y\��/bh���Y��u1��9l����h��۝҂7-N���#/(�̾�ˆ�hf�R%���u�Ҥ�=U�Ҩ$ڸ���ua�����!ޑ!�g+�1d-pJn�]�r}�q�&[]V���v^q��x^��y+8}�$Z��b�U�Ϭ0wK�C�kwXLY�%RX6�b8P�M���\��u
B"�`���k�0���=��9��2��J+\V��H����ۮ�Y��Uͦ��[��� n��K0WRy�u����Bㅞ-RT4�ż��@6Z�s��:�a{��e$h�o�A�m
�m����^ҩrVB*g	�������^, uB�Y��h`��WӃ�� j�~�j�a�^H%\L��j��k���b�`h۾��0�	Xu`[Û�ִ�NC{����דp�q�0��3kr�Co!����\�!2v�x��9]N�۔��^�W%Lt-��Q�`���_I�k����h����!73�K���o�ZBfk�d	ѝ��UU��h�j�c�<�q��@��Fkv�nK��N-*�f>E=ǝZ#9�cv�"l���Y��n���5�2��U�WԿ��z�ٮ~���v����'��5b���W�z��9T�2o�]v8�o{sO=�B*4:�El)�
��'���+�'����}�����u�u����ݻ��k�jt��q��%n���4�S��������ۭ*eɒ�ʥ�ǝ����.�5�ٽ!N�yZ7�����D������홫�r�MD�}yoj��m7� �c���K��d���f�B�):��l�6k�,S�Y:����Mc�3�g�������;��p�4$Y��n��V'q�u��S��-.Ǆ��!���U�ΆЬ[o�fM�De�I�&�+y���ik��tZ�ח�i�����h�H�嗖�.��Z�k����)���������ԃ�������Dgb��Is��r�HX#��������;`Ǻ��1͓gCE�&�V��h��rW�C8=�{�,�E��ނ�/+2yw��d�Ղۻ7��L� 
R�Z(c2KJ�p���y<����z<�ʽN�tmb�I�(��L�I�j�T��j#cj�����<��٤��,dtDDb�CQ4G2k�[S�[Xk\�Y�\��6��&M�m�&��Dղ�id�l���-!M��I�tP�D����$�j]�ih�Ѩ�j�Z(��í�&���[Ri�:k&�iӴ�.��l4�F�h
�)�C��-��ִ�ATV�h4f��Ӊ��Yڵ�Q�F�TQ�DkN�@m�IAgQlj�5[b�cA���m�Vu j��6�l�4j�&��K�1;h�sͥ���	��Ŷ
u��UE:�ш�&"�c���HE�*��M`��a�C�+N�h��V#^y��R�����2�k�T���T6���.Ԕl�Z����:l�-���=�Ur̩9J��5aD,���2������V6�J����	����&���*����+�� �G�g�I�	���s����2�5w��B��
��_��V쀼�b��JVpg�>\)+ҵ�%VhΤ�ԴT ��=�5s�-��fyx�1/Q)�vL�o*d�$=3z� Ŋ�!�gY�fͲ�dgO#������z�O�xN�7"�1�ag�w���]�֡�xȺv�Ђ~k�� ���������v>5{*.ۆmF���-�y���Kꋓ���㐘��!t�y�Xʅώ�2���):��P�bUԷ'�-��	X���s4{�����E=	ԥ����v�I�}^���}�%���$�����5�L����8%�ؼ;�{ ��U����ƅ@��HB1�C�\�X/����|e�tҤȑq�fV�(v�W��*I��%��N�x�6#��e<5y�� ��;�T��q���a�P�Q,D�]R�2#u�`�p���/6�E�g�5�a;5�^w�����az�Cw;���CK��<0���Qo�N�
W�XUY��i�L��%�;1q�O.�v#dP�����#�k����_�yZmyu������M�k���Î�JUx�`P���'�=��I��{�m�ř��zקX��י���y9-ծ��o��Ui��v���[b�.�g-��v�l�����5ӽ������*���w֛\.�<�I�����t	�N��V7C~x<�ͼ�}��5�����I�N�Mв���⨰�k�����k�!����9s۝E�{t��U�w�0d4=6�k0����,�9���4-_�J�`2�Z�9/LeG0����y����w9�!ns8T���'�AC��G��29��s^��e���,n�@�нY��B�F#,����3ӛ���U�KkP�Pg8�w�ƈL�m��%�'V7�ۗsV֍��c���c��-�ܱ��?=�Ga���~�V=9U���K'�x���_D<��\��*��;v����ީZ���;��1��! ��Pn]�p+�'eJ���
����5�ғ�m~9����ɫ�]���Y�0���+��'�K_9��"g;��t�P��ܻ���N\��w��,�x����q E��{Q�]yU-�^y ��ǡUٔ(�Ty��i�Z�mN6�~��τ�e���}��C�^1L�65�	���9�lc%�j���t)��HL�'z%ѓ2\�Z���ٝ�!^�u?{����B�-���L!ݘ����CM�e��xy�؈'��^>�D�M w�^:v/�a�V���4��)J�h��h�:k���θ���<G�DX'��hL.kP��s������n󄹆�Q<�ի�Zc�:9%�ǽ���˽im�OW
9$}w��{\y��s�����q+Slb�Jo��i�mܑ���P��c�f9�?5����s���	�"���}m���-��Cj�L!�|�*�K�-�I\���]�{,B�5��d�E�Z���Tq&e���!�����j�C�U���/��e�?+ٝ�ح�ˡ92��H�@Y��"�RtÔ�.�<S����u9jw�^�YG�7�J�Mt���(�Н���BeS��t(��'�����Z�O�`� �L?1OJ(^I��G�uWkur����#�-�0�kuN�'o+����a9BB�w9�I�����P�v�mE�Woi׉���f��Ti}���8���"����ۃ[�-l��a	��xb��ު��:���e׳`��{�sJ��m��q���d�#��;k��ێ�[q�Tͮ����e��,_�K)��X�ӏ\fy��nY��ɀ�����ꫮ�:�r7e�����{��vn(תu;�f�v��K���=$=-���a�����\�'_u�-?�SR
]���~�-�Ĉ�7�`N�k��ƃ�6��4�L�~b��D�����o�ݛ]x]��N[z�C�8lڧrs�@˽��T�[�+']X�}������ʈ��N��WJ��x�fl��-<�2AMΟ����k�j|K��+��	�;�j�[��]j�(�j���!�	��su�4������b��Z���ݳ��h�_G���ถr�5!��fXE�Obz3^�oP摛����$���YA���W6�e�pm����0���0���ZX*��~���9Tq�c����+%L�Mp����.��<[!�z$6r�әÙ'h=����O ��[E�E�Eǧ�*�`�HvJ���8��KU���7�!v���ͤ���SI�O�[A�u���\8M��b�j���D䦎S����o�ZC�l=\��'9D�/`�4��Mw����l���� ����:z̳��3��lJvcR�u_	H��^�"S��b%9��E1��&����O5�[$��E�5m�U�䵥׮�P���0�m"�m���a�`��w��$��S��<�Q*��1s޺����*\cG��/O���=�� �y�t�sd^�5�aR�6a7C���X�/��_#Bs�<�3��S֡�!'�j-#�.�a'�?Ha��`�Za�\i�L~�>�G�-�t�Z�~�߼3v�;{�l���-`ct:*;��|w&%ݠ�gf�G����{�d�o����i�E�CV���a;SX�^��]���	���aыͅF:�q��6����4�LaX$.�9"�K�C��f�[���9��'�dV�A_B�a1*|dr�R5f�"/J�.���z+[�'_L4�!�r<��u��P٥�kĽn�ٛ�M=X�r:$�_	ǯ�����_�M[]锟��O$+�@�wL�~�@��P=G�_0O�n~��q��ǽ'?Nֳ�f:�n��I�O���BՇR�uy�k,{����LW5����0݆�������d�v����h����t�^�a���AzM�NF%�q�|LW7sCk�xL��O��.k�X��C�!�a�@/�?3�LL,ss�5���A��u	�]�0���r���}I��:_r33��297C�>sͼ-��!�[�X���GE�Ӝ��J�,U�n+fZv�;�3J��NԔ� ��˴��Z~h���"���	�!���w��ׇ&��X����3��W���#�PqB� ŨrCP(γ�l�,qL��sӼX02��ys�vV���M�ٳ�Iuu�鬡�6���s��[��	�,�,k�po��A�֬��t��s���gm��܎���
�DIq�&']�F�k�Z��
|ε�ܢ��U/5�ʢ^�B��A=��Xwr��{���2�T\:�\c<�-�B�k�xI�r�m��-C�$�b%9�?�r�m駕�2[��\ONL۳m39hz&�]pR�^��0`���e�Ņ<�cHg�,� ^���ѧM@]He��yJ�(���B��b��[��Hl�(���l9:9�GIwg+W�ΩMX@�1c6Y���dBѻyu�p�_`�j���@�l/{��k���k�%QN.�l�0q��аt�z �Dc;$\lʯ����0���;��\�/Q�귪4t�W.m�q�J�(�%Ɓ�����[�	܁!�!�O��.���v�n]�L����噚��vж+�Ɲ���%<�)�Taq�Ao<��vk������c�
���8�c��^��]����X���Ru�IӴ�U�\�Ԫy@%�#�%<;�v;�ܒ��t�������u����c�LK����7&�Yc�V�TXP���f�V����>�*/���i�s*��5���N�p�\0g���@`�O�(LhOH��ƅ�u+p]�PK�vQmL���0)�x�tE���/A�:�^ÿO@`��fp��4�|Nca�n�:�j�����i�g�X�u������:;���͇i��R�ǜYr��D���D&�o�'%�'S���M;%�b��\���UI�]���v=q����-�tg/>חt���\�v�V�̍����t�����)�����a9��kL�C���A��K����e]ok��<��YE���S7Dpm��+4��T����)K�٘).�TU���[�ZW\D��c`b������[48��*���s�{=�{���z�\	��v�8�_#z�X�Z�
�Y����ND�|l 5��
�n�y��]?���V�<v�U�&��{P#-�=w@���|#2Q{��Ƕ�fƴ��-B��%rDϛ@��t�D��e߲��-�f1z�((�~XU�EĈ��/sQ�]�0�ԹH\��C]
58 �#mX��Y���+{x�8t��8hy�:�ϞBcH�0Y�?;P[8%cj���q�g��ӭy���f���jԳ6���"��c�ǫxjkgk���K�z`$'��C-��z��)Ж��x��؈ݥ�|[�\p�n��)̀T�	�EP�ː��w�,C��BS����ޜ�>We��e\7VB��	��^��e'XĲ.�s�1�%^6�6�󆪈Oݞ�f��]��_�q�j�)u����^���׎r�8=]%ߚ�����Lk6FχF�5��f�Lm)�����P����^p��#X1�lj� �P�n���P�ʮ���^Q�S�ql����=���o)��,!�����������5�6$������/��]�ZBf4Y^K���9?n�%��!R�~(eW D�:C�0e��'f�Tt��U��ژ��܇���$x!u��E|N�Ǘ0��Wtn���4������i��x̘6I�^��~q���O����)���[.s
�H�*��1\�ٛ&��G�Ό���U�p��z���K��9�3� j7���8칼OI@�j���_�u����c���	{��Q̮a�pt[���?����G}���{ʴr`����v������E1rd� �:�,r�N={��5�f%�3����぀�aﱶ�3	��XE�s�f)�<ӭxN����!�f�Iz�c�C׸��&+����^�D;�!sZ���w������GZ�DJ�Obv3],�6Э�a:IX�'\2ǋ�{/wӄY6pQ�����y�$TG9�p�Dy0�ҡyF���ӛ�GaG����m�ue��g��'Y�/���g��{�a��D���Q==W��ӵf�:�n�C�>s6V���(��A�F�:ӛj�]l5[a{��͡��b���636z1v�U���70��y �yY�岜�m������E[:
�#���e��&����B�$ N�[�^��V%J4
R�и�˽T볐gzwe ɪ�׽�kޖC�����s�~F��"/���	��I�ҩQEP�vm����D��)�f����C����4w���e�K�ө�#�{�;Ax�N�:��zVe��b|�oz�5��|�纯���Kr��Si�X��s�Eʡ�	X:J�o�qLe���M}5�>kh���e-�J�����gyE\��Y�_	p9���:�b�dT�net6��o�� �Ndr���Cv7���T�M�Z9�g��<pf�v{�o[�ѽ�E�.�{�c찷!p���]\�v?K��Q��)�2�X� ��9ٵ��O�8��|ʐy�0-�#zDl�3�%3�����Գ�<���7�*��`z&��gs���0�� !���0�����Ww'�cj�8}$Ђ��NM�)m]��UC6Xm��ǻ��9�����滽 ��t��/�����j��\��˺�Ę�hl�
�^b��n�a{ӯ�ƃ��}���<�p��e�|^5����-[�P*�g-�1��{��WFwt���z���3�,�F�uf�u-��o�5���V׼�����1�ه����m�A<��3�Ng!�4_@xITu���E�te�=�9�{��ԫ{�H�<%+#O6z�Z�9���#�Yo7�K��]+�Ƽ��w��ڍMإ(`��kݻ��.I{{}^��J���w-��,T:�QG�=Ϛ��Q�gtU�#f(4��l,�����K���R�ʋR��0u��S��#���Us���-�������^�X��,tC���d}�%.�D:���nn���q:�k���ll�HP2
�$�ư2Vzպ��ѩ�e�n�V�x�83ja�3T����ʌ�L2��6��K��Ǯ��HHs?�����{^��jdB� ۹ۈ��]>�Aer�N:��5Z���l���qxw�Om�D�Ul��PE�:BF�w�V��) ��NW5OBh��"tnoI�F�5O��v[��ȐFC�.G�HW��幂2��O��ȭ����Uc}>�{�@J\{���rޱ���-��x-\�3W~���-X�8O��x���"qAVK@�4�)�V��:�[ϳ��[c�+��K�f�e7oj��{��e �ȃ)9���UesҔ�|Wt���;
�S��^q�ٙ+a��KYaY�d:\�T'��zQ�箨o.U�]�;һ�:u�ޞe������~N�`���8IH�Gk9RNʷYj���o����z���o������}��/du?e
�kdU�K=ó�t������h{���lm��.��]Q,V'd].�q�"֐[v��(�mt@��I����:��;�Q�Q�u��^ʊ���NS���۪�E���T�D�,��*��`�3�8�ɣ6��ȝ�!��gvp �:����l�7��F���J�o6�	#�܃д��r*�$T5��a2��7�E�`�;��X�WW ��Ʈc�z��|��@�>_Iה�}���5F��]��m�ooK��GS��eW��=J�obm֨w;B�	in��aa�6���w�����3R���z�B���jB�m�K�\��4�Cz@D�e�M5!�e��+����52><khU�"F���w\ard�&W��\�Z�Z��3νV�Υ���ƶ�����q�ܢ0�*����h�k�l[�9Go2�"-u���+G+��Cv��*���/tB���B6�eʫc��%��b���żd�7�&cBWe$6�,�{���k�SP�Z�fg��#��E����W��:K�{1��\��«a^��]b�?���}}%�]i2�(TėLM�͙�����2��r�oq���!lwrS~�jݤip��<;�mgu��̩�ҙY�ĸԎhV�Ut�{��ځc
��lQ��sv���^v1�R篬qy���	4M[b���6���>kjP����V�V�+�4r�s>[/]!���5kN�S���K
=x��)��t��pv�v44g*�-K&��jS/�eּ8�Y�aI�@��K�sPV����X�<��_%UP� s.����V�̡.E���Wqї��Q����Q�RUU�k�B�n���x(�Va�v���SQ��X������zޫ���.���Ls
/)f=�*r�e�v�T���X;�$B���j}hS0��7C!��w`��B"w5D��"�L쾊�=;v�w܇[�ڜ7nn��)�ŵ�ƯK�+o*)���}�b6�&�F�G.*��jb�k�Aq�/ ���m��)�p�e
;��^
8[�-�0R�x1]f��e���u��`��U4L Qx����-Z̽h�{q��F���z�'K��u<�ԞB���m�lҾ�w��fO���;��ۉج���+�Ԑ�we��mW0�qȀ��wx{r����դJ���d��̔��1p��F���Y�;t�d�̗�1ɛ*d�Ȼ��Z�4�l�X>�7��0aV�.��Met�v�#]\�e�'H��/+M2����\�m�%��J�&p	��\`ն�)v�]�;QћW��mX ��X�&@�6���n駢Lٸ"��(^v�d�����L�u�[6���vu��F��bۉ���]L�uʃ%�'>׈|r5u}����6|�m��V:ըe�Đՙ�P�Y:��2�e��eh}���@݃�����}��@��J��T�=�F�ПW}O.�w��$=�M�ri�r���������P� �ICX�1���UPE6�8�)li��lZ1�i�4�<�.nr�[T-m���-�&ڴ%l�h��:)�.Qb �э��h��s�����F�1�F���Z�i�P�Ӵcjձm��L�DE[&��*"5��5T�f���lV�E��F��FJ(�c:��AE�j�E�AAAU��Tj��-�Ul����Am�����QmX�mZ4V�3i(�Piք�4b"b���kF�
�4�4����1Ú5�%LPi-�m�AE�h5���E:X��UQնj�tQ��� 5�EkQ���))4�j���f3���m�m��TkI[�¦�N*Z�&�gM;"�KT��SEQQMU�H���#��cAk(�N�Cg�����m5����-(�ֵ���0ElU�UT��X�j��:����Qc ��.��Y��=(`����fK��)�\ǿQFnU
�:���4�.J���\���ɖ�Ų�%Y*Σ;�;�f���$����~��4᫜�����o@q��c,�zOIO��<3�bbSTz�V�v߳�䶙��sE�ڰ׍�0a�p7���x����&,3D�z�7�vu5��/Xǯ��q�'��������C�4����mcu�D�^EU]*��tN3�%�W�����ȉI�˚
RE9�ʋuStN���Ƴm߳�!��!��P������x���#e �&G"*b㕙�=���º�����)������:�%~{�4"nz�b�j+�aAo��Bʬ�|6�*�Q�;7C9�N�֜�SsN�e��+�����n&:�J;6�7��A�ު��NGf�ʫZW� |��eQ�ˉsb���Y$e	��J[�\�f�μD/W�r�x]\J��U���|3-��@���?e-���9}�u�"��>�#µy4�2�
�xEkGh'�`�"?�Ϸ�ݙdmUUXGߧG����T9@_\��������n5X�	�m5s��ڗd}v*%e^�N���a:��	���S�΄��v2��Lc��%s�S-nT���9��Wd�tA�q�.�ݪ��]�Ԧ�"m��Y�$a�Ffmi�[�7�t:��	�%�� Ϭ�R=E4z�IVJ�*���~L7���Z��ok���f>d�)�dy�;>��kɯO3Ek�:�j|�O&��ӷ�����+��~�r�������b6J�D����No�?І� ���s�#թOfy�k���cC{�����#gV=���mmה�8e�vLi��Z'�ܪ^V���i����K�O__�� �V�|�C�st�������d���+�����Q{�:A�|h7@�Ė
e3��S��B�ьtm@x1z�"�>ϯ��c�E{�vI1��9���4�4q^�WGWPm3ㅨC<+5x��7E嘑��<X���j������zog���8)OE<xsd3�Y�6�G^Q�ͼ�"��Hi��t���	/�;�P��>$�B����s#e��E�� ��hD�'���*�7�Hb�����̹��O5ɪvFޕ�����^��h߭�D�6}C�[>ەzUj�Vҭ4�@|�Z���׳)�Ā�8&^Aҹ�;�2�`�7��o�4v�ϴ�}��2q-�o+���8���V�2+8���!l�$�D��c,�y}A2U�]�ۯ>O\�;�v��؞E���"����W��Y�`���fӲ�z�קջ�J��ӫ&6w�[��̚5N�qX5�74歓�#�e9���m;Q�*���A��	�����r�J0}�~���6۩��3�e;E3�
�G[��V���@6���%P����3�	u���*KA3�	9�ݲf�K�E��}�o$5ә� ���?�gӼ��*������~���pr��sN9���Sd��<óWP=�Cf>�Ab���}]�<��,D�X�1#�>N���sy�l M.V��qsl����t`0[F�1�߫r����@~�<��->ڮ�U|y�
+L��v?aC���,8e0���6���m��qF���MG*4��PR����P4�H��a������5d�e�-����%F���T;"��1+����r&:=~��9&4N�ߑ6�z�bνY얕9���C��A�\ŧ�x*a9�cph��6K�+���)�����EZ�>nԧӎ��ۚ�;�[�NS �_Q��P��/&���W��I{S+AkE��k�V�x���1��,鸢��ns8(����9�a���d_���z���i�EEJO����g����79�&�ϷE���2���9���:�~�:��y�fp�בݹ�p����[<'��H'�<tQ��s#!�/�⼒K����[3v�=E�o���^�j��#I�|��#O4K-sӜ��=�y�m9s�,eL]M_O\Ѿ�	8��j�߳cdbo�����/)H��:ۯ"�D�S=���p�}}�z8w*�h�=Z��xړIv�:�����hk��Ӳ�{#���f��Rg+�X�r"8@[��J��,�R�1X���9��˩={4g��:�O��;�>���L�9�A"��[I楺���-[a�u�;�c�T���x�],ܷS�̉ :B�4���ʹ�KBi�z�����h�a��Z@�n�#|�"��L��d�s����_�	�\�u�.��)��;D�%�f����Q!�(!\�Z���*3��9N;y�\r��贼��q��.(��G���l�k}�{%4�����db*|�<8I˺�F��M�1�{�,u�"�5�0%�Q/��̀�j�A��il��vSֺ��V5�5����ÿ}�I��EK=b5?��i�<��y�a�U�<�����Ov��u�hc�v�t��dY���bUVW<�jJ�]��ur'J�;Tm���55�����[���-p��;#ΝoDl��Nz�]P�\�Z�0��2�EcU'�̴2��+�� Mt�Ln0t7��5��#;U�J�+|}h�����F�͌'a���uq���P�V���Sto�h�q$oHq*�["�/aWN��Μ3�:�{�QB�J�t�Qs�=�x�c7�0"����SJ��WvU�dQ��k�q�d�5��l�V�*�"G����1�p�t�[�6o��~�C��:7c�zM��ܯ֊��.1"m'	
��T;��X��-e3EQӛ4c/��i3�b��)�m]vnm�"+��F�|���z.��"w3���L�� �<�z�J<�rk�1��Y+Q\}㞯)�K��72V����o��m�^ZV��/�#f�@#�=��q z��Z�gm=���>���Ғ���%���#F�v¿j���jO'����g6��z��wE.Lݽ�Z�ae�(@�dLNٲ*0H�ޱ�a1E�d��WV\��F8��K���v���b�(�w]���t�\ӝ��)�#��|��W~�T5��D����Q�s#����*��)�^x�܊�s5l���V$-�#9c�N���C�����\�)��q)T"���e��3⛁�ϳ*�&t�N���|�d!�O�IJ�/��7�d��ۦ�Uؤ�8�cj�^�{��0q 9I��'x)B����$�R�\�md�h�̫�Z�n��Q��ɶ<y7�њ���rh�z+^���%��}m��^�I��T��)�[�������[��|��6��$f"����찎����m��/"�s���k������
�oPp����Q{��e�.�FĜ��{�>~�ZR��D�P��`^J}��9ΧB�]�f�6�v�e� ,�E�A���v��Nq~�v���>�E��=���Ha�z�?g��%K�Uʘ�m�k�)�R_u:
vYz1�o�5�T$m���خ��{;E`�+��mJ��$\E�=6;��=���8�9�ýR��p�W	�Wd6���-�9��q;
�v�!�z����*�A�	[R���dL�n��77\}�.v1Sh~$*��e�O!�$^��mG#�Ǥ׸�a/�k;�3)��y�[���>��/!�c1�f�n%@f�ǯ���'����p���S}܏����r;-��J}�N��j �t+�?$���63�W-�jֈ��sK�p9ݢn�\��a# D���S�O^Y-xG�B�*���예�x�[��;{E�td�P�C��"���fڑl:��zݚy�:6o�b˛�#�~R�uf��ɍ��B��R�:I�T{2E�9鶖���	q�3jr�K���!\�� .�7u�+G)D���^��Kcѻ9c{���9Ul���T�tU^��|��t�s��۠Ύl<���l��أ7��<f��nGe:�p8\y��{���Jo�gL�*ʵv�n�火����C^z|	��{�ُ N�kA�!t��8�?�Ӱð9f)WK��B*�󾵨�T*�ŐÑ�"��qx�ZB��J�ͪJ ��4n�T��c`�=����c�!K/n%YCi�4Ct�Yjdʖ[��YZ��c������" o��r-��4��y��9ܔ�i��
��ZO3u6⽉�^�4
�|��旎ۮ V�Ej*()Zh�E�l����� �	�f.��v�"j�kb�ؤ��Lr�S\��
)(+���c�v�]�.V��XN♧պ��C�a��s�o`�Tiɺ�iJE-ފ��U#$=��C㤬�Q���`Dy�j�F$f;������j���Tz��)-j���e�DY�����AO����|����#Q��[Bx�(�>��~i���8sr�m�D��)��&y8��6du<�:9���E�Kt����./'�͹����\��:`nƌְ
�=du1��p���}�^;[�[�9�0>�݈�=�^��Ȍ�#���p�E�h?���������9���w�G({��"j��jԁ�(*���E\�����I�����g*r���p.(.�=T�D��1r%�� ړ��C�8W	U��*+c;�Y�h��퉝�h���Y�tE\�g.(Gٌ.�b�+(��Hr�aޣy�٫x|���T�
�_A"�8-��o��{�R	v�Vr6#��3><v��2�3v�������� rw�⚧Z���6��^��KB��:-֊����+��gۄE���~�Y�,�td���B΢�5��/or����ׂ.�z���T�H駉� y�	ȹ���7orȺni�m�{L<v���>�]�Y�⒟9�T�N庑ّ��C%fR�"4�s]`Zr�r�
'��s�U��K����j�3��X�'"1n����w\�2��bO�{g���U)���CT�7����ӱ����ɾ��~��j�t����^�a�C�L9�5=C�*����%Ewح�'d��۝��wH(`�8��>`r�ި�*�2,����I��A�k5�7|��^l��_�Ϻ�?�?��k�+�;V��&���+T�F�m�z~�ͻ9�d�Jo��ޖ�vo�s@#y�-�s��j��{<φ�ڸ��KD�˦�=gtl�i٣a��Hop-^�m!|$�H�2���S;�G��T��bȁ�}�b�^
z8a�lQK/i��Sp�����E;ʙ�THo��+�U�k0uL�|��L�Z��B[�f��fۣ�\�^y�:��]�7�}]lm:;eK�C[*��˝��
>=�8�~߶�	��ȼl�Ӥ�#x�d�;t��s���3��*�'1Ww��b4c� �J�/	�n��{I"|�Bys�y��.�w�v-���2s�(��"�·Dy0��J�m�u���DH�q�wfȵT���������A�M>��oO���a��t{KJ_2Uz&�E�ݰ���sn,E���}z�ټ����+�񔺚�D�ݖB�����GE^E�S�yf�U�]v����oJDق�vHn�%͊�@��e,�f�,�0�8�Wo^*�B�y�E���AH���I�U��2�3+m��e�6������^����^�������Eo��IX/��=$�W^�G4���;yK7��C]9�`���)m{Ӽ��QE4{:IWʑE�y�c]G4����h���w��l���M�-�5�8�l�3�Vuʠ'[���x��|���I$I%�4�U��\K6�Yy�]<B�Ӷ]�����f�fV���T?n�y�W�ʂ�m�}w�7��j$4��1�M.�JNV�=�nu�'U��}ȉ��:��j}*i<����ڮR���gz�౗�/�����TcE._Z���=or��n=\ƾ��nJq-�Su�ۻ鼬�L�6xj����@�]ޮ���4���;���]��$��׀V[��V����Dh��ʆ2��I�љS�15�LΤ��kej�m���;�ew2�8�%�IU� �\�wѧ��u��r5Q��{.�.��ك�o\̉��S�+���NϹv�m򛃪0KKW["�Q���)�z:��B�0X�`�{��j�t;�A���H�~W{]�5@��O_�2�m�r�����=KR婟��
���G���Y����l���)�h�����A�fV;�(lÄ3j��w��8�)�j�k.dyv�*H����PE��x7-��s�!J��Sh��-�;��5�B�oz�Q-ז��ڂ�j�E���<��z�Ίum+���%�B��q�x�1N�O�J୤�fթ�t�ʾ���I%2jի�3�����e��i(�#G*��X7������c��%�&���H��}����t�;.ھ��!tFp���Sq���s��tzgm�����N��n9�6��k%�aW��Cs�G JTM��T�ͻTu�)��Kz�j�Ow�R�SAź%��r��b�����
�*�!&;oZdJ�uu8�W����D��pX��Ȋ�(Z.��}0���b�8YTU;z��Zcnft���� 	�j���z��=���nE���ݥ[:��!ˊ��6��9R����e9E�΋�^�q�v*͒|e&�u�%��(η{�`��2�r�SP۱�
�8�H���;���IӴ�}qE�d��}�jN{��HB�h	ٴl���]�n�4K�YÚ�iʜ���7z-+d�1]���g�R҆��B�7���I�c������� ��XMC�N�*G�oٺ�/f`��M[jH{xd]���uz�.nڨ�)\ጺ��1T�ʝZ��q^0%Ԭڽ�N�)`_mI�k_bWz�ٴ� �]�-��n��C��9�6#H���:9%�+M	�o[T�[xDcn�N:��¦J�3+�����N=��D:Ny����7�Y�b����(<�3f��wN1�P�/���"�c�M���bd�c�3���]�wEWK
M,�g�U�u#�;#i�t����β^L�{
����5��ͭ�����!7�(\{�u��ΕJ¥W�h�2Z���%hӂ⻈�8NEv��)��ٸ;�&d�9^ɢ\��S�sK�2�3-��Wԩ=����݀a|�	ٸIO�ڧ���^��R�%�U�5��������V�r
�<�-��"U��oe�F��Y��c�*ŞY��+)�QAܷ��vef�<W`����_�Y�zP�ql�]h���1�[c~��,� X,! Q4��˜�\ޱÛ៯Eb�[:)լ3�����֑�E�5�MM��ږ��vq�5�m�F�F���Vm��Fu��`�6��6��I���Q��IN�Q1DV���k�j�m�%��&���4iѱ�ѭ��g4�j��TVڊb�mTD��Q�QT�h��m�m�4�Q��F��3Q2��b�Zt֚t�EI�l�$��P���:6�5AE!�v��i�Z�kV��0��-�EDF1cQm����V�65Z��:m����%�TE���֢��Z��(���l��lQ�U�������F�E`��&��֤��bحSlj$��*)�h����$�*������A�Ӊ���"6�2Vڣd�S�o���)���5��ch4�I��\�ĭ��b�����iأ%4D��SVƈ$&65�i�lS�Έ��X��h� ����6���;`�mm�[m8����"�F(ӊ�Z�*&�����b���%�M���Ѣ��F��DcV������b(�j���gw�p�����cZ)��n�@��^zw���WЬ�	�� e��_Z����4K��艙�o�U �H՜�]�k��f� �ѡ�����������$��EK�y\RD�E�Q���[}}a��~��eh8��35C]馹���H���ȡeeR(��Y��wA��i����ަ�*�`�u����s�����@��\�`~�T���&��0.r��]S������e�|n�>�����ܑz�׃����{J���:|v��tte����n;���CY��8c?�F<�f@�e���E�<A�{�vtOS�;x�n_m����)x�jM}vt;�3�*��J�����p���r�੤ی�vlКm=���U��&���g;���OՒKI/�����~������⛬-��~��!(��WK^]�le3�c�
Dӳ�\tFA�jV����ٽ����u�E�^�H�䄊�:x�41������t�5=1���x�
Pѽw=^U��ɍ���ue�@wAZ�:z��va��c��{U�]��K�J�ú��~:�o�6E�1C �r*���=ԭe;����YծƼ*�{_<T�j��~ҥ��]��sze�z�V���1�b�8���<��k��͏�C��	P͙Դ�KbbYo��5"	y$��}]�����5�+~�k�H�[��[�Q��*v�����>wO=�ۍW}���DV�E[<��vEm�����H�8��s)�f�S?f\6���2w"��}��S��Aΐ��B���oZ�iГB�C�;[�y��s�<hk�I:�����=pB`9`�9���Kf]h�/��X�����j�o*\�'����so�|�9�Ȉ�3Ug�����z�A���;��W-y����˱�Q�*����gLޫ냛];��u�:\3�0�e��gUG4��)J�b9o�uX��]&�u������;��F�F�#>���I�]̵a�&���33���:�:U!Ӻj������� ����o��^���3�ި����n���nHm2��[�� ����=!��t3��*�*�������_��|�G�i;ǜ9���3�Oq���w�5�1�j2BwD�z���p`׫&�_]CH���+-�(kiaz����7]nF7vI�B����-}���
r�G�&:u�RѸ�V��st�2�'��#u}]����ur�l���ёO��P�p�Σ��X�f�F���tq�tQ�cc �t:-N��e&J������5=ztN�2���j��"4���[�S�tS��L�J��<l�������s�:#�
�=�特�xvN�YBDHr�t��E�|;$�]�9��}Z��V�GK=��@`SUG<Q�1r�-��A����片�Տט{����+�����Ǫ%������,�$,�k%t[Cl�u�.��殥��9�ݛ�(��I�`�;��/SL��s�H<�x臘�ըMۙ��o7�q��q,��IHsƨ=��~�|�~[���m�$���4�5�͌�	F ��A+�gB&��*�<���l���rk��ni��ɼ!�Aܼ���>���9&cxt��*���(�T5J�`k�+y�]�gh{ֈi�L���:�&=e�����=1��p�k{�r<��$��?'Z��PJNN)�,�����Sl+bt��p�;k��s3�˧�/UF���B�P�p�O����U㧟6�*M�J\�P��͋1TV�_I��#�[np�b`�W�O�P��Z|�9�I5dd��\μ5҇P�y�����!�E��������R�սB6J���=t�Ewʍyka��so�7�zR�TW�nʺ��a��Hހ�\0+�3�d�%�;Iڍu�fI��u�=��i�w�ԬJ�7��=�G3��o�U�b%����^�wK[w
ҍ)e�u�.B$	�V*
�("WC@�ּf�7p�|ьtj�<+4#�5�d|�h$H[�A1�'��a�mzc����oʡ��B�<*4#/������$�$�Rq�3P��W�P�٭��'F��ȴ�A��`=%1�u٠f��Dܔ�KmC�<5flH�a�Nr�Z�e�I-���=�6�u �Q结B&:ީU�hi��@ȼ���by�d�oI���c

@WF@K��������8B���˄+�G���u1ý*�U��!�9��$�B�B�v�ji�[G��ׯ�� ]B�`��$�6fE�]pE�'vS�a~}z�V��<W�Z(Jӈ����>�7v9`� ؜�N�db4�m76����:��N�0}.`���x�rʎ�8v�3���I:��7.�S���ְ�2]�Ѹ3x+j�غ���n�J��4M�M��͎7�K0js�Q�DG��	˹�X4��JT"����Aȇ�"D�t��u^�wS]�
�C0C�\�[�L$�:�1��.�)�}f-�*���\�o>��o�˫��\y�]A�d(�ѝ$��fb�<�n��W���wY�}
l��0��{2m���>g�>�\���&"a�#\t��w9��y�H�[���y�m���l?ɝ8�4�`�3ۍ���7�IP�r��QyB�9��k�����p��"��Zڂi�`��V���i8�sR�#��t�)bQ
������/o�v�p�I9���Ԩ�U|+ܦ5�&���[�n�zT^��S:�b��gVM��c7D��v�!�׀���_fz����<AS�
"�t�R�W�볲-M�sDW
wE����Gw�xVhF�T3W��^\����n	d׉�T������M���W�P��Jo{�+D������uۋp�'�.�=�>+��'�I��*�z��b�-D�;7)k�u���V%�!9D_>���![L1���AN�W���%�8A������V�͑��4��7�G/"�8��	�T�C�N���c�z����v
:��c!�p�t�dD�c3LC˳��W���#5�舜�]Ib/���S��k�0��{�ƛ3FM�m�|�g+�%I�{�.(���J������˦U�,�+���li��p�}|8#���Sw��t�������KM��Ǳ5�.���ls=��~�A�1�,�O]�E��d
���m���'�5>\zoH�_�/�$CC�V� NEO��Uz8@�Kʧ�vemب�l���ݗL����EU>�\��/�\:B<��[�����*U��vXS�WŠrR�uǹ�H�'WQ�2ُE����E��F���F^Gj��7b��}>9�x�rJ9J����;%w7{���&o
���Q��ˊ�B&OTuOP�3>�K�-RQEw.���	:0Pt�/ʩ��Um�3�����)ae���!�h}�]2�M�0}��� �9 :S���X䮝��^~B���}�l�_tgi�����H/�V�	v���b�����V�ѪN�� ��L�@�V�Ҿ!��eg�xf�b�8m�p�b/�����n����W��<댈��Qƍ97Tqp�E-޹�X���7A{�~�0��0q�#6Pޏ8(�wd���bWA.��sE�]���U��}����|�=����Pn�N����؍z5��j�u=����ڹ=�ƻ��;*��ݒLt��du1���gDF2��P�1Kh�?WoH��p��������s�q�'y��xjy�A�'-��N�3�Lg�v��W��h}g%>Օy����$Di֎Yj�6+�Z���{�7ї�O��p�E(
3�D�Uճڐ6_�p�u�o�q����i��wt��T�t���>�aDyꧨ�=C&.@\�Ɯ���5lГ6�GKl�k�o�G�co�\
�s# ���0�B�E����_^�)�]�Ɵ��w8%�l�s�t�gD�M3�B�,���Ri�}x��*`loLNgfe�m̋9�龉���J�w���iwj�&ܚ����t�����V6ěR1�h��c`5��S9�a��z�]cVR��/����M
�2wv\��&�]�ӕǵoC�-��Tޛg7a�{ǫu������:�NHwEmξ<�ݐ5�F�xF�I�ǻR7.�
�rL��}i���+�V����r�"
>�Eq�tN�U�E��eoyI����k�<��^�>�^g��]�dy���t�U�)��Z�o����S��Y�jU�oC��%�K'��t��dY���*�+��'U8�-�9�ST��eu�lɼ='yԨ`����`��V��*�ѵ�Ɏ��,�;N據��Og{6��%U��+=�>W[�½�����`W^�n;u�U˧�ǡ��mo��L�&��Y^��J�+�-��-�7�9�]�_�����u�h�!��79˖��]7^�=Ѳ;A�G9���V�Q����аc8��<�צq��2�"�q&�qh��?dS�����%7�-�C��p������6,�j�y����זbt��?{�����!
>*`�v�QGՊ]cd\,t|.��;�n�cl��b��@B��7\w��[*T�WR�:n�]w96����,̲-P�4�siJ��!��m��GwZ�^h�Ɩc�J�^YM-U�'by��O{�(�������nVi��[	F��yu�o2�^]H�g �ZR�ں��oNy���c�a��+�9�b��L��=ɯ%s���PowPA(�|�2�{9�Y��jsW�y���ge�΂�\�r]xPS�td%�ה��϶YТ�[7z���vh�>�	���Y1�!aH���&���>[w54�V?>��sR&!�VI�4���;�)YP���0_.�t�L.�%*����s�j��i�m������>�󦀮�C'��H�Ei�>�Ip/ōl�Y�_	ؚn�Ʈ9q�_{���w$s�5ө%�.��{S��!E�q�8�4i�B?\M!�׽:?͙�~���o���Ŷ
A	n&3Ww��M��52|����a	lW�Zֱ5�+�����2��ǘ_C�-ڦ�l�5���˱R��;����di<�q>�;���i���o_�I��#sYKi�����eö
���cӅ���Θt%�o�j�-P�S2$Fqd'�{/C��OMMl���,�s�u�<���l��R�Ǜ�S�fܧ*��X5ܗ,�Z���P�يS꺼��qA ��3��*h����<���q��t]W=����i�|�~��ꎓ/�F���
&��qp��0�r�z�ښ����L6S�������$��#[rE�Rb�u�:T���d�Q���h�U��5� ����GHv��}�>�e�/K�|�WE��3�d���\��$Y3�ΐծ����/��<��
����A꾞���P�r#�����Fu�C!� ��P����*3�l�f;;�
����J�t�gq��X���.�ԧb��5�-��j6:��i�x<;���j��"T�^�J䄊�:x�)mʹ2���N�5C2��3�wi����Wam���������-��>
〭k3۵	��&L���ĉ̑sNdP`���pxB�S녳��D������A����`����g�?ywj�U��)���EP�<G����z��^>D�I$�l�͓m4찙��x֝^�\)�ê��yضX�^��'^��d�� h|Lr�}l�Y˱vW
���ȅl��c]�>�v�s��L����7����[�s8JV�ke�@�q�T�x��kz��LR�<<������Se�ZܾN��n	cvv�� �v.�Uk/��a��-����ψ/ec��ZR|%/�]�'>s:�X���g��r��!�&P��PGw5�^UF�f�4a!.�$Xҫu��Ϧ�l����|:>����T�S����nZ�5�E*�Cn��[�5f�^*TX���v�#m��A�pm�^�|M���U�۰�����MLmfaN$YƷ�NϯD��N�	�y�l��][S;��Tv4RsC�Z�[�4G�]�ZQ $_nz�,|�l0#�kN۾����|�Y'���zd���݈��cPuב�4sl	��Z�OYw\vޔ�͂��汽�I5��J�1��.-���|���c��ʁ������f5
�Z�u�Ep��j���md燡��L�j�c�,q4$����4;���elpuk��\aXkZ�@cv�<μ�3���� �H�rD	�J�I˶fk��u��5W;yٻO,vl��u��r@�h��`�B]��Q�-��iB0�kZfԢ����3U7iI�V�7�(�3���_v������uÛl�հjWK:)���*�N�#Bؤ����/i�6�]! �\C��!�u�;��Mzp�^��_o�����V��z�"��Q�|�3z��I�	��j�cJ:�+;�Y��\3^hg:C�r}�e�}�C��t��1��gY�u\�u�jQ���]��gV[ɭ5S/���H��sG�-v�e�M�G�	|�{f�ؒs<W7eO���W6ry<im��9�}�F�5PΦ]lB�����p��i�ň>R"Q�x��쫋4�.���E�z:���z�A���ݺ�DԆ^Ә�-����U=v�w6��]3uWE�6�Z� �hT��	��c蚋��}�[�hq�8\�z�v,70c��Y�3��⋢�N���q��E�A�Ʊ����Ff�Uôa%E�GSBV6�R��./D}Ƚ��:#�t5����=�	6Ԫ���r��a�w]��B[2��ӧ}���X����3�l��N��;
,��	���_!�����)f'w�{��sfJ�z�{�z7:wU9��A�X�ܩ�d�:�q?�{d�����]�%l�8��]�e�91,Fa]{��ŗV�d�q�M��f'�9	���=tb=4>ԑceh@^NUzm�� ���v;Õi��VͧK��˗WH��4Emc8�(m�*B�N�����+��%��4a�IB)�<�寊�c9�}�ؘ��9(ғ�|�;�i4�s^��v�j7���U������3�8e��%ƛw6�DT(H�B�|���.8���*�Ui��UDZ,[TD�Q[`�d��j5�j���#�k5����Dl�vsTQNv�*���#c1PLE�s��UE�6�56�Tӱ��-��PEk5DEM5U-QV�Ѣ���&hv5G68lPSE�H�)H�d��F*��"u�"J��"�SPTNژ�bj������&���gT�q5��mm��ӊ�6�h�V�6(˶�9��V��tD�Ƶj+b4੃QTN��kN�QETS55ST�SEEQV�lX��֊��i*(��EEDlꠞmKAMQ15A'5�UZ�6�&8�$�[5������TS4�T�D�CMDm�Z-�Z��V���"���CPMM�U50h�KMZ3l������h��*h�"����\�������F&&�5��A�j�T�͵h��&���j��	��"
�m��kZ�|>(W߾�/�o�������c1�͹G�rG>�=������^�nǱ�8��շ++JS���3��;�jD^�F�-ނY���hm��\~�A"���p]:�9�L�ΐ������l��k�NE�5�)�Z�IX�\k���N��{�{.+FSݧ��hɫ�]�n�-�	y��()Ц� �\���r���\�>���kE䨖ǵW��N^SYax;�Z#d�GT�v)�\���RQIwQu�ۑU[��:�w��\��v��b�0=~�<f:y9�:��W�����s�cY[��N�
��y�3N.������3�̈́7���;�oM'i&�[9�̌.��z�vs��v�A��OuW��I�>����.�����s�Cٴy��>u��j��������ݒ	�;G=���mƄ+e�6���S��Y����<YڋH�y�=�r'Lu�-�z�[�So�	�e�Z�:�ȸ�[�����GyL��ũ}�&�i�^Y:O	H�ӭ�^l���h{C�)�k�[؊Y����m��D�Kޗͅ~ԇT�^�6��A=�1_�vE'��muwL
 �5et�r�U[ǭ�㾪pfl�L{�mr�}[5w,���(Em�rm��ޫ�RZ��-��Een�;�E����g��� q]{��JQnd��D{�ي��5u^�;+R��f&��g�w\�u,}�θ�Wz�����������g�&-�a�p�y����9�����e�M�5�ZO\Q.p����0a�념����.k�sv��W%rg�^.B��E)Vd�K�a�ݯ6�4���q�t�fz옓J/��v�ɡg�H�p���:\o��))z8v�n[�:��k�P�5J:�o�y�zR��!r#\�|�W���.9�*��&W��繟�K�u��[T\��j���Z���t����*�i0��+��c�~`R�C�u!���s	����K�VH~�9�S�|�.�k�H5;��n�k������׉�|�����a���d>�ꍒ�:���&�-q���2g���q��x�]�*V쫭�a��ޏ0���,��NT��,&�&qp:��e����0M��G�l\s:�m���Kܸ�AVMº��9��`ͼ?J��y�&��K�\�A�p�#Un����ц�j���)f�3)�uN]�#�P�nыY�N��1��[@^�*[/3����o-�R'Ժ�(��9��Az��=�v�}b��+bD$b�`��#X���έYC�u+��-��:�����]+�ó�_�_�Й�j�a��V.8R!lV��;��kn}%nK�Yu�l�WPk Hm��
�����J�۷��x�"x�cz������1ɰ���v�7����<�ב�����:�q���7u���f���b#�:ѱݳ@բ$q�88+Z��9�� =%>�u��r;w��§Zݕ���4I����D��r���a�wPA"O�W�0���_f��F����>��qy�J[�PR���.ƑyjE�9�6ZN�ED��{��u�^���`̀���9��B�)"�*�vI۷C��m��=շ��xw7��N�c>�k!^4$:��˧�#L.�8��/;�m�n�v�{d�����n��>�eVKq��<p�0�W0
�3�RM��Y��]���?A�l��W��\��\���
���yM^:o;��}��ǣA��	�ͯ���z]{٤�V6�6�o���{�8U&9�1
�T�9��0��h�e�0���B�h�veoh<e��T�x���h�Z5f���)߹����ݜ�IlMK��a�M��6�?�#�����57�\?���󤶧x+!<��\#���n+���w��Oj�qoR*���Y��]��l���*&;UE>V�W<C`���Y���/����MVQ3�E�@F^<n���f����W�sr�'퉐��\|6�y�	�#ivq��(�,��M�2©t7xaD�U�4�%��X�>pb<�j�:�:@R��t��Q5�Cy��F��q��܍8�o�����G?��1�m�p�~u������O���"}��ܦP̍��C�6��g9��x>ِ1_��������n��M��d�1:=?�T��g�:(Ϻ�9��&4a�< ��ٺ��M�3c��"g�#O�*����4�7�������E9�������+)�2�U]Y�'�[B�u�?�舜�<���D�Uҝ�s�om���Z��V�K�H��rM����@8us����,�+"b���U�\��%:f��7W�)1)������E���'!tM���U�N|)Ս��k�oK��d{/�M�*�����Kn��'���WF7�:�0���Ȯ�8�_�3)ׅ�ɵ��e^�H<���:x�5䎲z�,�ee,m�B<K�s��kG�1��{/P���mbU�>�!mrAF�Du�\J1�s=u�]q�םPp�#�x.i��y� �,A�D_v��[z���0݂a�%̘��C���IJ�]3�r5[��[<�����F1�THf�Wz�=����+�@�H���*4�UA���t�t��q�V�z'�6�EgkgeP>{ Ȯ��m0��t���O#C{��x�Pg,�MJ�Y����Ǉ}>�!Lo��Rrh�(�9R�`'���b^�h9�ά�s��h�utJUm����鍕�S�;ȮZ�E%s,��J�f��C�2��wI�^�q�� ��.�\dFΪƍP��c�ߴq�4��4���9Bw��Q�R3e���oC���vW����꽲�e�:�6��%�jT"�.���%j���p�7W�7@���*��מ\�36��&wbYp���:`�W1Ҟ.m�h'�
�����2�fԮ���Y��Y�f���G�C�XQ70�Y�lX�)l�:7i2c����VW.����:�vw����3����6�[�vO��ŵ(F�R/�͔z��\�=�@ol�6C�<f�8U�[+wqF6�a�@ѯ�s[B-oy�,�w�q�'�[�x��:'�~B'�q<��w����r��7�]_�,��2�V���"0Ǆ��ii~f�v㛼Z6�o���ew=�� 0B`=�5WU�ò�	�g9�i���@匆�Y�*�t�*�������/A&���g��4�F^>d^[��c�dwoI���� ɵ%.��z�\�	�~���=�s����'-�O���G>�+9rC'�@�Ab(��%��;�>4�M,9�cS�}��ٷRη,�t�i�Il f�,V��r���%$�zKݨ�6��x���cU��秵�G�!s���"x�t"o��|�w��H4Ж���HJ���b�V	ȍ8@�&EN�w����F�>����C�FJ����U�1�U�D/4X5��m�	�tj��ʆ�M.��-�Ԯv�EO4�{6���J|:��(Λ�0J��c������llQZjó�}6p�N�KAC.�X� [:��3��I�Y?Y���N�q���s�x�faYM��j-��j�pݧHʚ&�kl�td�>�;=,1�K�VH~���5~��Y'}o�Y`�m��䱀�%�Q�h��yԨc�:�a�;��zFG�;�w�N�֘�69�T��<��r�[��;é��0#{�.8z�Z�MmgJ��}�ϘI��񔃥s�Z���P�dl�����~����Ѯ|gr�ʿXu�p�=���ƽ�#^e�u�.{�v�<��Fs/����e�e�Xn�C �g�Y���`62Sx���=�#" ��4^���s{��º#ق��[��q`��f�����{�ʩ�k�oQ�5=�u���W����H�R�9�45��o��11礲^eWN78����}��}���r[�/9�9��{�Hl2��x�g��y�q(A(U,�3-��!�)��k�h�%P
Ac�ƖVz3�{��G��ݗ��@�F�����O�
�4�������^(�����w�$u�.�	�.6��TM̳���!�Y�&H,�	�˗`�Oh����S����E�y�8H���O(��Nc�"{;E���a������ˬaAJ�2�i��q.cmD���:��ǝ��9o����4��8H[�W�b=�B�)")T!ve�{8w�w:g#�o]�wls=��N����Y'(BB:���w2K���zǚlhν鮝��R�q��r�t4��Dd������b{��=B��6�c�3+��Ïi��P'����ǖ�u#Y�tVקx*���ݫ�o���O>�S�Qr�+�����������` ��
f
b�f�E�fF�>�����P����~c=rh�w���h򴉑��HF^�؄E>IV�]򮦟q+&��\v����A@|��#k�����s��6�Z�b^Ri�ʭc���=,KX��,V��Z��)a]�l<��j��y���r�{5Ş�� o��q���5�$ޥA��j�yF��aT[�e���/�(l�NJ�Ηud���O��Шv��z��#�r�@�!b�C���?�tb �Rc�z37t.^-�k|F��Vʝӆ�9�9B}�"pg]���<�'��`����*�M�orVAF��y��'@��	M�n)��k�U���2�8�3���[��W��T5o�N��W�`}���5��XOs��46�Iߝ}�%zO���|tQ��Ϯ��;���3וwF���7al�oS�ɍ$׳[`_Z�I"x����`�;�>�l�ٷN�����'�m������8#���9�����䬄9cG����z�9�Y.ռz�Kɞ�%[Wߴؔ�B���������	�C��i�O��ӽ��BbXWx����E1 �3t��>�g��g�iV%Y1��B���`���Sw���������5�ӹg^��U�r ��ڲ��MT��qwuzЧh��~��D����>9w>�n����r(�w����z|�ϝϗz7z���!��1%#���x=\U	M�c��k���X�"-��3ϳ�(:|!���V�o�f�H�ax���\z{��}���,��v�+�~2z����/�֙J���m�A���qa����T�\9�Ѿ�t(�C Kp^�Wd#_m�=�Á�	lךG#�-SC��Y'P96��Ԗ��Y8c����d���/n`�%vA����#�&�"V��m悵32�)g���O��C�y�r���ɢ�%9R�a>�bƑ�`���Pܷ��~�i��ڃ � r7�6WP��6�/����ϸ\�#앀eq�60���4����=�f}(M�!�lC�/��#�a��髣�^�0���"��;�t�
�d��3�f���U��X��k�m�Ok��P־"���rW���uQ��;cdu��7����N�Mӕ�s�����&["�m�{�9�E1�(�l��_6�?Ꮖ���m�z�b3����-�o7Y�:�5��{�Y���J�� ��g~0u�n>�YM�:�B�/�����i��"'Ǐ�����9���rl��\홗���ŕ�:-��E����ѡ~�����=4� ɥo�͓���GoA�Mp�ia>���X�s�y�8�5��Oo����`Gd�@
��ADT_��c��Ȣ*-��8ol����2�ʳ �0,ʳ� L�+0,�� *̣2�2,�3*�̋2���
�+0,³"��0����̫2,�3"� C�0,ȳ̃0�����(�*̋0,ʳ"̫2,ʳ̫ L�0'�d�f�Faġ�adY�fA�Fd�fA�a�f�a�fA�d�fE�F`�A�Fd�fA�aY�fP}瞇�S� 0 �J�� �0��� &P �a@	� '��@&@@�TeD	�P& �`P	� & �>O &  �@` 	� &�UW2 Ȫ� 2���0 ª̪�ª� 2�� L��ʪ�
���� dUfD �UY�U� eUfPY�fU�U�VdY�fU�F`dY�	�y�Of�V`Y�f &U�`Y�gN�`Y�f�eY�f�@�W���=|A�w���QPi �UTU0��i,p}�;�N�O.�����T~/�׵/����J�7��^b�??���G~�  ���z^����U� _L������X����2�����������( �}~Ի���k"d�>���	������|���x~a��W�� �� �  P  ʪҪ���  B@�B Ȫ�B H ª�ª�� 2 �  H2������� *����� ��� 
�H?�H��A G��E���?��'�UDTZQ� � ���o��W�_����|{9I$�@Kل�}Y��Or��P����K+�^����2�v']�� ���P��<ȟ2� ������҇�!����%W�p���� }��Aa/���P�I��a&K�KF��Zcc��x�������?��~*�����3$��/�/%�v]��Z]�z$�I�����%(�  �����?��*������~_x�����Ӈ���?��~��t>@�z ��	9��UUE}'�~>�2���A�����O���"���#���F��H@a�ߑ�h��$�%�/�b��L��:�S:�5� � ���fO� �w��/�J�JU!B�W�VU4�D�����J��1E(*40[4$R@�T[dV�UU[6�l��[jU	EJV�I���m2�m���Vkomv�ҍj֤ҭ�#HZm���f�i�icSF�2��Ml�fj֚F�l�m�d��ƊŌd�kf0f����{s�Y6+CM4��ڲZ����ֶ�r鬘D������Z���+jTj�VƵUTԶ��j��i�#f�l[4���	U�ڶj���6��;���5���  M;[ﶗOT�p���W�{��j�O=�u���{�vݯ{{oFȦנ�^����D�wn�=n��/
��Z�oO^���oo�[���8����54�zzײ��.��;]u�j��6٤�� ,=
��v(P�=����hP��>�C�}�xP�@C��o^<��=
������ziw]�ݵ��w��zzj��5V4����{ڽ�{ץ+�{��'���v��{:��5�m��{h=/{ZZ��+K6i�6�k ����Z��]�g��U5��w^��^���v�p.�V�Ҟ�s�ޮ�ٯm]�g�{��r���ջ�{U��i����k����cv�L��v�+v�{ݳ���v�w7gz*�͈�h�B63i�ZCA� )�aCOjYv�;�m��J�J;�������wR�������6����y�OS��v�]�{��פ�zݭ��S�㵡AG:㎴s�B���e�fիjTTV�j�ֲ�G� .{�T
>����;v�t:�@*���\�뺌��DUs�q�iFc�U���'��n�� 9܋Y�K[n��h�3R���l�� ��wkGs]`+�lvr���EN��(鵃��O�*�uj���Zs��:�-+��F�Ӫ�(n�����.�j٬�J�5&i�bKL؏� ��i�(� 4���j@�滜jD9�5��hu� �V��7�[�p�ך����(��ǡ�)��Si���Q��,b��k|  ��С�:�� z�p�
�{����M�����p�(4y�j� M֍��^����@�z� :�1�Sl����jCL�m�V���  ;� } �{;�P��4A� zP n:q�@�z �н�y�@ �x�  6ݻ��xz�@@�=�6��j�����wnl�ئ�  >�C@
��� �=�� 
��p��z�h�@u��4 ��z =E� ��`= ���  ��Oh�*��h�B)�b��H��4i����JU=T`  "��4��@  M�h
UA�� 
DLj�  ���?��~���Џų�3����uMv�+��m}+���؋Ar�O��U}��_W�|�K���APE|QTS�PT_�PE�
�+��)�ߟ���k_����迂��o"����B)sSJ��'փ���/Z�i<I��P�̔���[��m�'�ʢì� ��Y[��1�/H�e]��(nz0���b�U#��V�l��,�K[f�U��7F���41m�.���]#��2�5�ce��;Z�H���43hayA�XI��M.�-\ !f",�0 �xfHՒ��8n�)�E7Jn����ܵI��w��Qѕa_�<���ۖ��愫)F��D�V��GH�i�k�6���F
LԽW�Q�CZ���Y�aD�a
jf	e��(hIk�w$څ�B�f���1����fR6!2e�p/�滘�kVN����P��>���4�h��YIZ9
�BAl"�h$�	-P�ln�D+v�L�=��bM���Ҧ)^��f:M������c��݆��GV���,���)zJ��TT���``����A[����������Hkh�͢V�Gr�rdQ�!,���3��q:�On!i��4��8E\`�T{�k)5-O� U,#eڻF7��N�h��	�
Ґz�˚.����<Q�+u��l�Eֺח�(�_j�SJKN%%�1|�6e�K�S� ңN΂ �\W(A��V�[Z��fm5�WG2�w*8���bt&�]�2D��r��{y�KUj`%����Su�D�JɌ���Vj�d�&�GU�@��Elu�,hil�%�?ab��\�Z`ۥ��m=��$��gUbV��2H�m�@�f������n��m�1A擔�2-=����R�O)Yt���N�Bq#���n�[+KSIǴ��x��s�0P#T�G���-����7 +U�ii�{��
��+jG�@��̱�n���IA-��q3�4�u�a���f�j�=�{Qaa��3������3Mݚ�QR���͊�q��qYJ�Y�݇�R�4n,J�$:�uk���ݽ��e�c~Dn+(;ov�Zu�� �� ����H�.�t��LML;z��j���Gj˼�u���hS6Y�J�c*G/N��dj�CS(U���1�m`�se�@��pi��I�\�I�v��^�@��!Em�
�^���ܬ�yKKݫkZd
�K�k#�R��T�j�`�{��S,^�[n����KV��w��'�*�:�tF�&6�n�(-V�XnZ�ӹ2��)a��֕��K���#9���-�(T�*�B��F�2ЄN��f�6�M���{0XIA�x��Nw�E��8�^R�J�3N��h}�`E��b�d�։d���b�1l�.��b�82[��OV?fkE�v�4dט�mh7�������J��^a��@�B�F9 �E��U�P�K�O+�2nԠ�f�-���gi]�M6�}��[En[���� ��-j35+�$94=q�����1 �J�{+R�K*\��zU���A��6���u���`���ʅnc[B���ZJ��Lv�M-:�]y��5��(j�RF�R�����W-B�"�
�%$��j͵*&���\�&��;���	�����Яv(���I�YI<��Yw����
�K\�v�nR���|]��HYdV�ܐ) �ʵ���Mi�r�r+a�Z�en�{�C��5F��V�1뿰�#7L������ͭ�i�M�1���+�K6��O)��yL�/f���Y��0�d�*�
R�b��/`[��\!k��B�n���%�T~�ɢ��m���&(���"�-��jA�����h����U�u�^�E��Ut*B�Cwo��:�,n� ��.�:�֨�������E�ٰB��f�],��VF�'v�5�>jeӧ �t�����$˻�V5���u�2nAu����;�&.Դ2�:�ۙ����@ObZ.�I�̭ӫ6��@�n�
�.�����ƙ����K0�����;r�Ӫ��-f�Ä�/�.Sz�+P�p^iʙQ���j��x�b�YY�K���G��+چ�����^^����i�J$����q��J^�2山�(,x�n����U�VowU�f�f%���V4 ��t.5��c	����B��ii��g���W�i�k����%|-b����q�gi���=���RZ�bp��d��b,�Mѫ��[{(�j�ʻ	��r��=��j���Ђɩh���*�ˬmf:ݻ+J��i�J�vM�Fu�2��m�ܺwnG������^-v�:��)˩B�T��uE`��u�M�@���	�6��C�W�nZ����
f�:�u
ܱ��{��*WQ�>�Œ��e�{(���\��)�"��64:�Z2Y i��swm��[�H��ė�-[�N&��S����&�J$,8���Ԥ���̻q�HQ3u�M��,k�}��t �X��b�WWT.	-����K�6e\�b�Ec�2�ͺ¨wa���	��qn�jHރ�/j<��3c���EY�L̸�խ��q�iJH�y4���^%j+b*��q�0�/�w5XjJEۗ�1-1F�4"��D���ˇ2��W�nEA�׏%$M���y)�1��9��3��b�EC��J�͈�\5t�@(Jj3O.Л�{eU�WM%d4�g-A�
�@�͊��e,;+N�w-�*Zik�V)Z�'a��pe���%�.��k1Kzop�&يF �JV�ǚ��En[ʉK�	�,�l�[2�DC�$��=bޝ���)�^��d��vӱ�T`l1ܩr�!�'[f��b:C�Đ��g���f���WJ�7Cm ��P,РVR��ϝY(n,�x��<�E��;��Q�:ri;5f�n���Xa?AZlI-umdInY��J�U�ْ��i�/��
�l5tƃ�k���H�0��V.�M�3Lx+�I�*��GQI�~q ��{���Fi�ܚi� ���f�������eGv�{X�N���`�����C�t)�ki-��;�����a��i3j�d�N9���Ų�S[��-�*�V�(��7e��q�e�z=[�Zڶ	
�t�sv�� !�m�od�O2�a���,Z��0&�*���Nܘ0R�V��R��X��j��j��\�Y�)"��Z�Gr���K�w��%��UZ�e���F(���dq:��h�M18؃c��쟴
	�o,�G`�Zr�q*vv)yE3ݳq�u���^g�+
vi"��YZ�X�7j�E5m�0^5�Q#k��e�VSMK�0���c;�^�F]#�j��*Q-���r��ф�ͫ��\�@�+kA����2���
��ءY��Fʉ�!y'������я�Ǩ�Ǵ��Z72؋N����Rɀ��#R�V��� �2��l5aZ��صU6�vH�hڸI�����n�Zjäj��������enP�b �I�+����6U���cAɤhᨄ�;wx�<a���7����5@*;��ͬ <ݦ���j
��qB�i� (��Q��u�K�m'���f�01R�!B.��.��j�w�l=Z�c%Mx"打X�j�-��T_���J�S<����E{��@��!ٕs`j�N�J�Ɇ��*KJM��0x��2Lr�YvT��aة��KC*CmPY��,�i�+�!�TsM"kr&J�O)�Z�Ō�HN�����)&R�"�4EB�Fei�k"�$��T���MT�[��z�Q&L�-7��.�a�N�Faj�'qE��Sr�+ (h0 ��q�f�eR�[���e<5(c7p]�J��ut��g0�i,�(Z��-�y�L�i��V��o�^ȭJk(l����n��u����a�,�8�(B��0�6�v4�0�Q�a�t�Xc0v��1�-��V�Y;�k�X��\�V޺�Le,m=C�P����6L��d��C�ncJc.�m
vǁw�L�[dRC1�Y)��ze�Y9��;r�M���6�L�F��#�51(%�wvՆT�d[cz�
r�A���X��,t�����V�Z-ވ�3��E��릞hzN�:�w^��Z#�L�q��+kXn��m�R�[�J�Y���;3>q#JW�tGZ�8W.�H�`XK)M�Hةh��ө�i���u�$\��б�5 ��9,�aՈ���ml֕��)U��-S4��@��B9[&9Iޕ�zUFوݻRբ�.ح,^���C(��v���ٳ���ә�7��;�[�%��i�LHԆ5@J�i���KO�*���9v� 	�B4�YF��|N�z�(��O�v�}�2w@٪�GJ�Rݖ��ic�2���@x�����j��˫��o(��SA�4�d�N��^1��	+qZ,,՗2�h��5�\�&�F��a@�i^m��t*�]+V��r3�m�+E7�����r�7��[���߃Y�4$) � �!�z�e�j+��MM[��J�.�TZ���\��[[w+.��<۳��%Z�d,�J0ZA�%{cn�/q���:�0X��m���R#QR�ɔM����7wnޖe��o�H��#Y�[�p�Җ�V�˽:Ôފ�LV�]F�T6+��r��Ъ�Q���X%�#�H#�hU���&�ڷD�V^�;��[CS�Xu��0�ݕ�t���<Q��LY��T�X���J�)������0�P[�N`Z�ZzH�����-%!�#w�e�pX��J�RvHx��&���F����5} *F�����ɩ�z��B�^,z��+^U��pdZ \���?c�c5q0�-:)�b���q:��3p�d	m�8�0��/���Q���Y�Qa�1�,
����Dum7[J4�9����&�Z5.��f;�A�#�vZ���
���uҮ,����.��A%�R'7\�z��y�.��F��:h����ƪ<Gq�
5��} �u��r-�0��b<ML���n���{�r�HR|]⥛L������"�a�d5N�2��Vm5�HbV�3t�e�\�o@Y�17u�I`� �;KNt�;V4#X^*WRU�E$���^e'�"K2�-�r�q
ؕ6�S�61SLǡ#km�M��Kפ�fGC���f�Kq�mި�h�h�Hq�y;o�Է)��c[4�Դ��M]3S,��ּձ�W����P*�FI�d�J�(e�z� ��SI�P��p`2]$���N��m+�KIҳ�
���F�V��5�W�R����nd<�՛cy�hU�Uu[вڻ�(�6���U�P�-���.Yq]H(�!�Q�*�<���c ֔��2;�p�<�	�+��4�M`L����M��֓��f�\��ǂM6sU���u���$��"�nM�:a�ۗ3d���hZ����.����M�VY��l�!ݛ��ffHi2�N�������$�bhܡ���Ee1���ғf�Wh��lI@-u�5 uVH�Z�b�U�e�Y�.�����ZN;H���E!WR�����M�W�B�	�µ�S)"�Z��Ɔv�`��!Oq�n�TV�ڋNT@|�}V5�K�
eQt�y�ؾ��� ��N[���b-���i+p1A���u�����ի[vtփ�O>n�����X�#+,�KA֢v)���$���9_XZe�}����'s)�BjcZV?�t��8`�n`�vۑ�5�J��5�h�[�`Ն�iZn�i�P�Hܭ8E��ͅ�Zh"����mT�M�{j����J�'T�cQLJ�:���U;��KN�7v�ۺ�J�4��%1˾��a��+vi���Ӷ�Z�oFd4U�D�����m�qe�a�/+*�:����VIa)�h¾MCy�j��:^m@���6��h�E��S�A�D˃(*/-�H�7 �A� Y[OF�L��6���J�0"e6�'je�k�H�Z���t�r�+!a,5��N��P;�39��2hB�c��SۖC�i��\���4� �����STm�4��)b��?a�1V\�Z��]���3�4&J��t�����f��L�* Ŭr�n�j*wh�z>6n��37~�)�w�����t����wY�N��vB*�D;�)U�3qA4�S�h�2]ȖQ1�iiP�,]M����0=�h��EF�
�Z��V-��,X�M�z�˳��f���(;č�$��lC0[���kB����;�tK,j�s>�ӍM�7��aɡK���Umm4�����B�dX%�,�t0��l��a��V�3!�Q\[��
d*^��:H�Z���f�����V�$6ƅ�ՄiV����{�,:��ځ�n�cOm�N'�H9H$�7(aZX�Y-h�uXq�^8���Dz�`l�� ���|��e�O��i�Hn�1�F����ij�ְ�V�\���ʒ��F�_ �b#�\�^2
�U�ۗ�%��VIG[�v�)V����!34���n�8����d]�KK
(�Y�K5�fm�M��z��[a'���BcP�6�>��PGn���"��ʁ���%�eK�J�����`�Dfm
��#�HXP�u�ql�J"��uu������b����ښ-����hj��+��gVkf�hJ�뤆2��rۭ�H��ս�VH�۳���.%ݳ&��G��v�u�5��F�D�Dh�2����(�Z�ȓzp��0���̬7f�){X�j�-HUӘ����XK6p.Ak����M��	�v�ZI�݌Z�,l�QJ��F�yyjmG�-GJ�P�r�8O�X�G�(�O�v���|��ۺ�FKU<)nec���vm�Nʪf�@�;jJ,�� ,52��{�^��AooI�%���YQˢ�q���VB��,�S;�"�T[�\�����J;]��9�J.��/o��Dj�2ZYx+]�k����i6�X=N����u����@��)�濢�ݹ�wQ�Ʋͥ�Gen.�-��U�mgEl�;�����$��Ս�����k6�[\�A�W����{Իk"��c���-��P��L�A��J�fRn>uz�!`va��qE��m�|���x_�݈uzr�!^�L��t%�cCb��@"F�w
�ͣ�r�L���*���G1�����CfxG�~:q�K<NϬGt%��WQ�LE�������v���ηC	콲��Z�nᓹ��j���]+
��y���6cƂ[�ͼ��įJ�/ZO���ء�X�6��PX�9x¡s��ߘ�;�ƒ�w[�5U�{op��Z��C[e=:�)s���u�O:s�{���:�U��͸ЉM�yZ�m��.�"�k��FlXُ��*õe��/��u���Y�53H���N���ݭpN���5�=FRgb�o5�-o�V��GGr#FmCŐ
�Ǒ;	Ø7���7'^VB � )�p5����+�GU��vm��٦�\�\����ؑ��Xn\�]c���u�i%�Yu���O���d�ZX�*e^&��}l<7�嘴�ք@�mB�pY��ʜ�Z,�Ѷ���TF���0�=~�^�>ҀW�B�y�_.��/%�v/��.kX�htՍq��e��[����;NZ�U�
wSh�Q�V���fh�p��ne�,�HOP��-�|]ѕo��I�Q�J�z�4�b��x�(�ӕfU�"ʥ��-թ)l.tM]������eG��+on��j��V4�e7����;+�aK3����4r�(�5ܥf*Җ�S�uWۚ7Y�k���By���\�k�*o1�㾈@�e!�<+-<���e�Yߡ�'̠�D���Z�I�ož�ʁe�\�ɒQ�QJВ�j8�2o��Q5��#�xM�ɂ��9�B{(�d9���e�ڑ)�%}�̼�ٶ�����`�ڦ��b�ޖZ��ʤK���T��9J�����)��U���6�˗Un!�N�¤��V�M���Fڽ��}ma֩k/]+��qYW�����ڈ����r}���)Qj]lq5g�Ѡ:���6�7����9��-��-������=��z���}�hZډ]�����.���60G�b��6�7@��vu�J�l2�C.4١��Dz��(����;{*�G1Q�N�oK�L<��$*kr�]B�\6���Vwbj�#W��܍ƶ����k���IR����4+pQ����]+\�B��@�c�U5X���t��^H*V�m굵�g9%gk)�z���· �;�P�s���-D�]Ε��p	o$���κChY%�ЫJ�P뒯��ά۠b!�c0����e�:eX=�����O������T>��d�㘖V\�\��e����+[��n�j�yٱ��-We�s����3��dݨ扪�(l �ڬfNd���꩓��ѵ�(R���n�3d�����9��a�up�d��f�e= ���\�!��xGh�t�"j�,q�3.2�)���j4� �@�6�1M�cwt�gQۺ�X���kr�1u�x�7vok������G~�Qo;��h`��щm��u;�V��lW(bNYGl��v�(��e:f�t�)0pg���R�v�g%j˷շ�{�����O0{:�����biC�VS69��6D�{�d���>�sq����\qL�]r�Y�A�p����r�yJ�������Zfkh�c ���dx82�v�K�th��,\��QW)w��֫	��!!r�Y�Y������ڡ�bj�p@�]$��@Aʼ��Cv=����p��)׼*��p����	�å����Nϛ�&���xD��'�B���M5�� [j;϶Vj `)��E������;Y�9^��h`r�=��"��5"��)l�
�� ��]�1�d$B�[YJ��ghO�`��� C�Yi�)Xy� v$W"�R��dwX�yY{�ye��� ZC�����7����c�d���ݺ�B�U�j��Vu�l��N�T�@z��%�zmτ���XDȮ��[]��͸��]�����qk�}neҭK(���*+�G3�a��p�H����(֕ȼ�3MW�M���Lhik�>H����@���d��f��{dS�n�}X�*rT5ʹ6�}�4�
>Ә> ��� ��K��wW;�#��JW���G,4)H�:�wR�縻	�:�T�I����A]��0��8CP��w8��ڜ0fe��������Γ�:j쮹Ҧ�6�y���V�>�&̇�/(�[�d 1�M�bJj�α�:�˶�MP�Αw 5�D�ajY���٥�5Ε'��t.��N�]�Pm"�9�2k/�d5y��P:0��B%+��A鼾$j�+T�ǽ��N��!n@�fe���6��v���8ԯu�i�����ut��w�@'R��><�f�t�c#H(B�k/5ш�R�	��-cE��F�9&��P�I���0[�y;,$[�R�Ԧ��@����t��#Ga�.k\��,=C�}+:��Z��j��GwAM��*�,<���V)ո�hZX} U{��;��L�M�UfL��Ktp��$����v2v�,�t��	�4������z�/� ҁ��A�r������i4��|6�,i�+1�{�(N��9�6�6�q �y�������n����ז����� v�e!�e�'>co6�B���Vr:��8�iy�>][Dr
a�f>�B���_ko̾��F<֛�wx��5�� 
�����X�\��nI. ��9n�A�)Vc���Ve:a��՜�c*����Ԭ�F�U�����-响� 7n,�AQ�(��a�D�w�h��j�(�{cd�E���ʻzWS[3xS̀s�55���j&���w8`XOS��f�I��e<��3��Us��M��kJ�uΝZ�U�s��XM���.;u�q>��@HM���է�����t��Un>��l�}�d�TE얤�XЎQ�;7!2��gs%�v�2�h&K�%+Yr��V!|-{3_P��f*h��]�c���p��K��{��v�D�b��U.���5d���Վ1���U�G�Q��=�,m���,�Ul��2�>����|�l�e:3��sZ����G����HB��K��Z���Γ���^�M�SgZT"��}�!��V��42ú=D-�U���m�1r{;.�L���7���4��]�%�����o��`�8yfc;�C�f^�7�-��;�a��&�Ƅɧ�f>���IV�7�]�.Ʉi
��������,V���ܼ�_4��B�ʻtV�r��*�[�]>����2��r�#���Z���でw����}��F�bƹ��f�1�N�|���K�5euh�yJ��ޱ}�T�)�ţ8,^a�	|��6
]it��'j��n�%�W�8LA��x����d��uy�� ��
ۥ+Pp��K���ׯ�� 1�㄂�������<����hRN��r�S�9�e#��u ʤH����3S�CzT���a]s
ٲQ��)�<��ë����=�5m�,�Ơ���h=�9�Pn\kh�aU�Y/�]�7i*b��Ş�v�vֱ�q6��{]�,Di��Z�rX�`捖�oP��7K�I�6%*X��x���Ю�I�u��5��Ut/� ���[[��
S(�"���
�H�m���p��)>`��6�-nI��lс��S&�\pt�7���@,�֖���lUul�56e=:ʼ|*:
,�%6�C@W'����2(У���+��\��<�ty%JˌbN=�����'c����@l\�ܼӉ���D$�í��P�f^�Ԋ�h,���+ԡF�g�D��X`�N3���ԣҰ平/t٠+� �V	�q��Q���n2�r"TZ�8L�P��u��`�;���rD#鰲/�t4خ��!9(�1�Ů�u:v�κ���M��y�YF�}S�뎵nuT�;WR�m>�%��î��h�j�SA��D�r�ځ��{E���r�ͼ�I&�lׁ�d�}-�t1��	��WT:�S���V(Ռ�u��:pA�;����3,���틹����؂Z��ޮ���.����GMX��6�RiI���V�2X�[�T6�r�/Y�,:�\c�N�N��r���d��:��.�昩E2�5x�'{b��n�6�Wm����N6HΦy����;�uΰ���(�j�&+}
pd��5��|&6���[״9�c�q�yvJ�aq�n��=�;�%�\ҵ�;�cd��->ק/�`��m�[�����+Z邮���ѻ�u&��ʙ�FV�z�r�7U�GrHW�~��nQ	�5��%�6�z�$���U����f�3/q���u�X(Ƣ�M�V�\��T-n�4V�Ib�٢��HюnXz�m�fl�d�;o�e�~\UpZ��F�-MΜ�n	QÓ>s���`L���5�VP;�z�#Y�Y�A-ᖞ�
����X�H^��0ۤՌN�d��k�J���Y����,tJ���6P܋X��B�����3:��
yJ;E�9d�c��-7�2���C��75kT�w��Ռ�z�-W
�ʵը��֘�'J��P.q���4�M���ָ��pL�׽Hk�h"Y��@�����ڛ}�gCY�ġ��қY��ŷ�%�m�Dġ�ט��3��{��j�)��jf�Jyy:GLa�q���U��+4LI@h�腜>��o`+v(V7s(b�u���LWY@��3�P���<���kb��K��Yu&���wZ1^n�ӑ�T�H6����IF��@ܨyھ%w6�'��y���:��x��!�����;���Sl��}�+:���OA�Ȝ�2�\�0��\�WvC&i@�D��E��6�a��z[�>���u�<�SGp�&RJ��ąa+�HƉP��ܬ�H:���k�Mc�M����w�#�S�«�������6CH-U�!�T�q,
4�qY�w���.\$r!����lFn|�O�,��G2�_e7�կ�Ci��=)Ѣ�,��ŉ������Z�d���Ӗ�����P�fAV�Z���	 ]݅hˍ� �t�d�(7��yw��h��-1Ì�3 �Omo�鍣��	��PQPP�9m�j�{vz���4�qɔށ�j
 o�c@���4�`��z���t���#��9��K{��p�L������m��4�ʶ����S8���d����պ��,+ZV��.]�{���������^\���k[�Xn�U�Q�]�}5+B�u��@_^�mT9�ܷxƑ�VwU�%3z�t2�g�\3@{6�s�r���ǂɬ�����K ]�O���ho�r��s��{k���3�s�1�Y�K;�yr�k�*����4��B�hnR��LbW�)��|��c}���Z3+9r�c{h�xrN��p��N+g-�YCR�x�۵�,��u�)n��C4J*��sm|����W+u��1�����}�'��%�]J�4��vYm��T��[���k�ұ8���"J�}B.����:9o��(qʚ��e����Ⱥ��[%���h�S ���%���RH� ���K-Ǩ�����s,,5ٜ�T���=]k5���W30�P��VV5�2}�R+�|X�̤fހ�q
5+��Cz�.�s�:�m�v6����Nu��Fk�Z�8����Ƙ��G[n4�
�A��6�:��ɠS�o�;n�t�q֞��V�q��_[���hʹV*:�:�<�.O��*�X��p��T{U�X�a|�Akt���u�+@�0t\�r�6)o�bO�D�XZd�m�x)�xik�2�I�.N�Q\�Y������p2����-ӻ�}ά�S�U�� 
�Y��`�ϴE������ۏ��OI]�NL���r*Y�=�K���z�s���+n��$�]��M�O�$�j�:����#��d\��w�)�(�1Z�=))�vGr2��GNa�#!.��[kz���7��M���S\W9��wWu�>=��N_\�iY��V9���ƃ���Xf�
���o�����c��ݝ�B %�;���y��A�FD���W���`Ô�'�ݖ��W{��Ç�=����u�ޜ�0v�M�u��c*��ʚ��sV��`���z�906e�=*d�1�A	ʬV�I�����r�|���S8S s�J�'���i�o�Hs;xE�,��V�@�N �䔳0S�Ԑ��!���2$��ULQ�ƽFP#�Yi�f"�dn�<%���tj�a��,؃4�q͗�4>��]��]
R
x�v�}�օ츯�d�%%��kF�M����őb<}���K�Ķ�ɻz���Bי�"��Ӫ*�t���v���!Z�Vw@S�^�B!��HΖK��I��#��s�=/6T�:�a@�+����`W�:�;d�I��6�q��[n����-ۮΊeL<�4��]��LM��Qu��P��]tk�$�w0���0>��QZ�{&͛$��Ml`�N�Z�d��MM��2j:����q��kb�ڭee	<:v����L]��kt�!�s��E��iflN�Z@Q���$1V��d�7����y7#�AJ��䇼�o��׶Hsr���y��*├��f����)�o�5��wiEnϮ�4����6nl�}7{w�8���7��zm:y5�r;F�嵗.IV�A7�11�QQi;����Z�G KM^�II�z��E?�A��{��}�[η�;nL��e����ٓU��qQ׊�8����h��k�e���ۃnX�	И��A����z�4B�z�A]��:��T���`=��o��h�qJ=���\6^�Xim��[�K��!�	��=:��}�S���ۣMe7Ƅc�$~�̺���-ۋ��W9��=��-�`I�c���$� �v��{����Ǖ���h�Fd
���bdW������H���-;�u�t�ĩf�����!nK�)O�*��v�la�e!�ց�e�P�*�v\ٴ�1[�ҤΥL�Ǐ7M[.��r�j�f�ʙyF���İ^�/~�Pa�Qk���z�
�b"������o�W\����*h�\5P�]Ѡ:�5[K��:��,CJI�w�&���ze]t��ȮЖ	ժ�>���Nl�[0|��4��Y�n��9Mm�S\��K��u}1�7d�$��(���>�S8�)�;ҏ`�h���:lg�67Zss�iYS{��s0d7]S-��Ք{�/#h�'(�Y[�
/�q���������YV���i{h�.Ґ�1�{���N�:_	VO'�i幱�޸E��[�]vNlc�:���`�|����h�oVִ��^�v�&C��Hj�>�R�r��%��6,Z@��+ Q�����wM�/�7^v̆�|�z��kE>��+-na�}Vz�e�d�UMJ��ڃ�H�6��31Ԙ٬7:���AT�k%ۮX]��>c�W Sp�Ʉ�3"5�$�i�f��f���(q�{&�'<��9�ۂ�huX�uR�pΔ�1�n�ɺT(h�h�]��7u�[��ΒYݷXv����#�7�M���h��lN`vbh��9���!��(S�lôiD�{0ޚ={("��:�Kw�������xo�P��:d��T@A����,:W�\�o`�,�<��T�a�{0k��V��<�`�!ކ��ou;g,�ݬ�I��c�zŐm�����NѺ�$���#�:�mʰ!S���V��J1]w٥� T�MWf`˜7E��J
�\wN%mL�UeːP�y$���UJ����}���j��g�'�0�c���/m��c�,ޥ�o#8'����[)V���`�2�u��S	+����Լ]���X[�媲ħ˘���B�4`�x�霫u}u��c4��&$��ұ�]Ov����fx@��T�y���+UvP34�KQ�2M'ݓ"�d��鈢�@�����a���
>��ID c����bd��k�|��bm&���='jl-k�Ֆ�#�g`<��ob�[F��u�{V� m�W��=���gh���g*�@S���7��i������$��Up}¶�L�I�-ѭ��eV�du�i�u�Y�*��j��6�_^S��j��v�e
A�p�(�� ǧ@$�e���zz�p�r:����ee���t����ϻ-w�.�����G�l��Pzt!)���y�\V� 
�иp����4nrR��%ܭ�*��{N��m#�;����I���dӎ�Q�+�l嬗P�o��
 ��{;T��l��U���ű�A�0�'������b:���Yi����֎+��X�N6���')��i�Ty��ir{�#�t8����2�$6Jך��g7���J�P�g0��Yz��ⵕ(V-\���h��zgQ�+Tޅ��Ví�.K�AT�5t���Ҵ���jƺ��eՙE���\K1�NФ�\�v�{�C����'�js,B�>��,퇻�c�^���R;��ÈCk�!s�Ep��v� )�'��.V����˩Ge���].��*�^�ûϗZա۽�P�j�&���^�
_99���e+|���.-�x{��4iUnQ6q��WX4���d����m�Ne����Va�w�77(���kx�'��z�DȺ��nZ�m��ę���:�r�B�
�6ga�$Q6�cْ��G�en�Ҳ�r��c9ݶ%֟�H�C`�uG��J[�j���9������)}�&�c�f��zL��%	$�ųf�#�[��b�k�� ����VU<f���j��$�v�u���^�ʟr*-��lP�7Uw;IU�}���V򋈼��ĉm)�=��#���X�F��3�Y�觯��7�'���n=�r�18]������uh�i�F�؋%Y���Yշ�$;Px�e`�����pH�����
/: 9iCq�c��T)�ƕُ+�*(m���ȫ!.{�$�f�Ϋ���D���;����V�`PY��z�+:��n�-#��e�ɼn�]�RgY:��b��qW�u��u>Jξ�n�:�X�͜�1ht �";���F�ksx=퇎a��� F�H�K+6��X"�"@�u�rn�����n���+�ӌ�I���	jx뮧����6�g�sCq���'Lf�S:��H{5A[w�qV�)����O�_<��C5�����Vv���w�Q�ʡW���m���\*-���Ի�8m�괾�jM���t#Ku��u��q1zVD�#air��c�U�:s��R�\:���:e12;���X�!6k�6[S��(}�B���uKr�Y-�ʃ�r��V��Ȇ�\s��hA��8��"0c-�M�[�v��;gVbJ��V�V�d����6�ᾊ�Q��dT��ݷ��9Z�,Zi�X�X�o��O�8����֗�̎Ǵ����V�ict]��P���57�mv���`U�v9�gl�H�%����x�Զ�l�w����y8䃪��n'ES`��]���$��Vܵ{u���6&�]�W�`=* �u�{��(_J�P�ڸ䇅;�dĮ
�eD�s[� �R�;�;|���0)����rAw+��2ã����h-:hY�f�����
0}ʑߑ�rM���^8Խ](r��G�XU�·s�д��ë��]c�n�=҄���H]o2d��h�����nD��6i	����*�j)���Ԋ'_�INN\�os%쾵�P��cK��wKo�~ãIĽ�U���y���3s��9���CPí	��ZV���7�V���a��}�+'�m���\l�إ���&!¦(��|�@u�p33�i���zﲃlv�� ��i�iv3��hM�Bٽ]��[E�z�+�>q��+v��$[�m�/:'���jZ�B�ls�O8���Tf�P=.��z��.Z�1��3��%K���j�{��f�u6���T��39pukFS��D�o�n+ɕ7�l���j�LM� 4n"%����pdx�
��Gvv�=9e�d㙷;{j<�B��G����5(��5��ʽ��։��5�]��.np�V-�Cr�`������G�s2'��@Pг/b<�mi��F�,�]7�:ޛܸ�����7؋d��f�-އP`�l�$b��2�t�u�����5}U�-�V2-]��\3vA���5�7��ӭ���y@V�Ѹ�;��&�B��D� s�v��l�
]&�`Χ��U�57�PB��Pe�yft�j["�x��o�)8���aV���ǧ������Ɗ��4)�x�R���i>߁JBL��[A�X�i�C����8�t���uFk�9���0�O��A�S5���}��P��i��)Z����\g~u��Ju54::�zJ�SO��:�E]�:j= �HrH�G׍��ef��x�۔��v�n�����u�$�me��W��J����C0�7#d�d `*�1lӐ�T�n�wn�~�5^�(خ
K�-cip����YJ��i>�n�E	�R��ttFN-�Z���=�����ly�}�L}��Sz3�#iN�V^��;��!�Ϯ�%��B_T,��|�$.�F�-(�����n]
9�푻�e>g��n���MJW��ݻT�Z9���XWIW�����J�[NC����ǭ�Gqm�&��/bY];�@.���U�rY#j ��i�t`=4R�@P]����y�μ��V��B5}�2�Z��3+cN�,Φ�	Y}7Q���*����%�C���j�	�,��i�����pE�%��$�u&g��c��`2��9;&�x4���/�����B�t�]e�(m�lɅ^Qu��)Nm�x�QN���L� �r1�͏�G>bvc��uZT�sU����Co�=}���碋�4u��z�P�zkc��`rۧ�뙭�,ou1���.*빆����j�á�^]i4�$F�ǘ��%�g-��Z����ŽqűY��|s�9;
��l���s�t��d���v_e�L�:��Xf3)�d�ͧ���\�y���b1�W9ca�Ze�u.��h��ȳu�8�:��TKF=ɓ1 Sf�H�;�2��@���\�
m��+m�ס��[so���S-�՚�;�{M�mTe�붺�	��\����+�������^}����^���vk�JlR䷞v>�Q��R4����U6�5'8�-��%C��]a=V�uǈ��ޡ6�̼�"9�6�xD&��Bsy�'���G��Z�8�\+���=8i���Xv�to�"B_�q�/tD���I�Ո�Vf��Wv%&���gT��r��6�h'(�D�d	�neQe,�u��6
%�Ŏ\�>��-���ή5reR���6���#�Y1Q���*sn+L	�'��µ��nZ�4��������xu �� �����L�՝�u45���FP��nث�{��fj���=�8GH������I�ybV�xTю�#W-�tk7�=\�ժ�Y���a�XgM��R]�X7Y��S�軧ò�z�0U���4n�aP}}G��e�{��؜u�p��^#9�R���G��|�k(���y�l��o�]0�W\��
V��\k�Ԥƫ6X��S�ԓsD!6g_Mia�<C��#	��K�N���S��M@�eN}6'�w5`�/�u����N�'.G*���Q�&�l��|3��w�J�v��9YP��c��y��]������X���S8�us�Y��Y��{$��ʉRA�,ȒŜ��/����nQ-Ɇ��M�o�\���JA�5�L�40�L������9��V�*�`m�ŭN�Ng<���J����
p����G 0�ڧ�ֱ����F���#lWEX��H˻�Q�)H�Z����}Ԓ�����u.�^����n�dE�|Y���/Ulѝҳ���]�Z,ӡ�V"mku�eZ�DR6�t�W3Fp���gyv�!�K��݆���lۣVS_m۽��Ű���4&n�%�]��/�4�c�H��Q��u�Y��\Um���+Rs-7����b���R9|d��$>�� ��]��`T��8�ck9+Ō_J��m9�q�׻(d����v����:dM��]��7w�����u��y6�`���NB��9�ǃ8��!x6�03I���H������PfV���[H#B����k��
zWp�&�O�!p��3>u{#�m��#>ۋ9�]�(>��3E��FTM��m_��jY���8���F�I��G�s���퓥2�]�e�V)�U�+J'�⾊^>ёH1v�K�ۚp��z���k<Vr��C���K�s�P����W
��v�C�'i�U��q*�d	P���5v
`�x;(���YZuS�w]ZA�9M�۽�J���N�o1���X�����g%Gr]�C��:�SU�so��9XY,3+���o�-P
m�ebY�1�]n�z(n����v�fdu���9�(6^^��뼫����_#����U*l����F2��2�}P��pT�](7D�kz��hZ{Y��V����P�8:�'dWp� ��Iݣ9�e���[Z��܉>W�w�C(�j��+q�"#�n�� ��Qx�a`K�:.�L�H܋(��%w ��gw�Z*� z���D/K���P�߬u��}�lUۚ����9��½Hkj�I�N�J���d�z�M��ρ1��AS']*:��t�M��U�n���Ɔ��T٧� ;7�ޠ�A�ki����#��zMs`l�]C1��,Qo3p�
��*����F����hm�����k�W�T�ڭ��(�/이Z��\�'�h�/�2
@��Kt⳹V5`��7��6{���/zK��G�QJ���k��(,�XL��@=�ҡ�c���ZxT $�.��D]p'�]��d�����
5�[�,w(��c��%*Vh��'�����Q���-�!���k�ɢ^��+)�&�����㗹��i�ݗ��,���!+�ÙX���iHz�à�X���&����T��JS
JaQ7b�Jf�����e�cik&�^�%��$ĭJxb[�&����ٽ����/-\\��)`*@�5}ɚR���ݍ{kF�oz}ڰr��MVY�.F�*�)���1w�cV��}YP�XGW0�}[!��'MڻΛF�=u���Wv�JYV4X�C�ŉ�z0覞\���%	�-��^'�_<���<ݤM��x*�v��|���}��T����f�S^����yʔF;`O��ic�`el5f��lLj���v
��}��2��q�+�Ud�=i�.��j0"!��:�F<�4fNUp�`�L�9�K���*��;��&�&*�f��gO`|�ލ���KJj��"����=�P׀Ez)��"yL-۔�Z{4dS@x���wo�9Tx�\��V�8#/$�B��˨��Pi*���6����{�Ǣw��I����{�f��QJ�y7P��-ɵR�]j��H��pk(!��9�ޒM�rṂ۸�WHn0�r�j��1>�7�&*�`/�8�ʆ���o{��o{���I��Ԫc�������8��7+g
ar��o!8��m21��gM���c������Ds���*�n�IY���ġ`�)�[��ۛ-�z̛���Q9>�#�&	Y�/��6(3�j�:2���f�p��3�˒!P�`����n���¯�[Xkz��4Z#��-��^mû%��Ɛz�IK+��]�%&^.0�=)�e��`�-�PQ��+c�tu�`r
j�ZxZ��(w[/a��B9��f_�li���-�GN!D^��,K)�ӱe����ݓ��`����h&��k���9]��k��W|����V��y� *V�ޓ|�����-��ݱ�O��(�lh��.盓��秵Jƍmw&?��Ŷ�3�|�ֳ��F��۴��ٯ%g'xަQ&�GG�\��j:%h�O��'�������QV�bL�^v1����.���#�L���m��Ai��/R�8j��&�:�	���r��\�c���$ l��*��*եb����J��Lu�p7Y.L8
���ڐ��k7�V��*
���&·��gP�P[Jb��'5w��q�i,f�t靴$����m	�X�E�yP�K�f�:r�����z`�0��+��r�����J��kM�G��k"�p�W��v��ɘ�b/W�2��c}7pm|u���{�=�u�Y�xF�*ZJ�r ))���
�!b2�\�"�����2��ZZh
B�������
���Ji��")("�i�i*(�(�����������iB��� j��
��"! ��h����(R�*�hh����"JB 
 ������Z���� �je�JR���H�"
h�hZZ�)
�jjj�!�H�)��bZj����()�����
��((�(V%�)
T�
 "�X�hJ�Z�B��;�<�n��	]g)ǫ�و�k���Tt�
O��E-��9Wk�/���D���.!]q=��4K���
ar̷�ݕ������k�*O�5�������a����AY���*�0�� pSGv}��/�MOB��vA�ٷH���<ګD��t��M���}�x�O��|�S���W�;���ֻxE=�~ٜ���}�i��_�<#���*��� ������l�� �3u$���,�!�!���n����Lf��Y���O��jTk���8��B����7�z�g�P�����ka˪Wa;�`�w�N��ʧ痥W��˿U�N�;�~O�;���I�ە��
��*�L��k�N�,T���Ӑ���/��+�=���O7'u�T���/���6�xg���a�S��qخe-��'숝n��b�����	��Gf�
T����H���ܕ9�?�m�2�BN�'y}��W��\ߎ���$�|'�x�Ǜ��̄7�'���j���k:$�	�N��C��g�.Ї;*��`�(�onhV��׼R�A�p����UK��9����uD�=t��Q�Q<�E<U�T^�{�3+�>&���;���v]���"�_u,��%��3�!�����xQ��%l��K*kl@s��V:�˗jB..�C[*�RX�s/'9��e�} 3��L}$;��|1
�Y�ɑ?�-��n�de�um�(��p@�C����p��]��yn�1:�0�%�\�!���9���B�Qd�R�e�ɨ�v�O�Z���m��	 "�O�Q��N̙�mg�s��0��>y�&���5��<��]��h����&w�i����ʃ/�����N�$�)߃v���s��ʜ[��,5fce�h�g�1?J�s>Y�b����&.6��S6Ln��W����T��^����Ӳvޅ۱xA��i�X�Ux� ��� ��E:���P#�D?]ׁ�'�3�"�KTP���
��nc�T��x~pɸc���۩�p��\5d�QW�����,y~�Y]����|�J�4ͱҸ\C9�a'�M=���s���uUw���3l�h	t�3׷+mq��#P�*r����3LAE��)�M*{~UGp��vz:u��8�g�����;9�k
����\n��j����Y�zᜪ�m�Þ����2c9�9�)�b��bus�(G6��8X|H�c���������eNG��+U����̠��:zЕ֫�'ȔR w7B� �K���oosX���YW9:�׋i���ȰM�f��:r�(�.�V��lf�MfFΦ3�U��<k�=j���[k8,��o;u�H��D�����Wٛj󕁯�Ѳ������g�teJ&��ʚ�0L\��P1S->3*u�L�o|d�/=wOB�Eg`����2pыi�g��,�W��=rU�{��YT_o@)m�����������3�()�Ӱ@c�g�����\���y�CT�h�j/��Ї�꿌s�"\�'{z7����\����݌����.�s��Tی���Lڣw��ۤ2-T\��E㟲�jwC�c�W�?�1Puc��x�V�
�g�F,����2K�X�tHBk���t�o��]����{��>N�����?_x�����~�8ڿ�̡�.��Ȓ��5���r)Ӹ2B�dt§-��-I�D��w����Q3�n�� �Ơ���{��u�t>�DV�곡������R��3��V�8��Ut����\��N��.�6��,(�$��ś�GO�tݼs1�Y���g�Hd��3��'Pf�u���fn_$��44��U=b<E걏��FԶ�`٩��Z!�4�gȻ����w��Y����_SR��I ���Jst��;�\}��p�ssʥk枨�vD�4eԢ�坱�G`뭃`��f�,󽙡u��4�:OC�W�rjcZ}{�;*�;9j�s{��ϲ;��I5c��ә����5;�Y	�*`�{k�M�}�������6X��KΫ��;�j??��\�S�=~�=|�>S��̹�Ī��9�-�������2�I��:Z���Tԋ�{����UTW½��Bg�4�ﮌ^��׮��f{,��f���E�ϸ��m
u����6'����{���LS
m����/mg�ݸη��љ���("+MS�43���nW�~TE����=eQ��u���g���mL޵w��U��Q78�=���pS:z��g�-�V&v��8$�%��NKk#��nw"�*^n sC�-\�S�̨ڇ0�*�F���߅����YL�Yυp�A�$O�K�Ģڇ;���M�X�%� ��<���7:�;�f�C�1��&Ż2̌"%#MJ�j
��g���ֆ<VX�+������m�]���w0c�����滙}Ղ���z��:����ѣ�,*�KȜ��� \*>dB�촂F�)�a���R��]{�z����$��]�AK�]�,#"_J�� �^G�C�xS��5�z���]h���pQ��*А��]Ȼ88�6��ǐZIm�n�$地^�ћJCX�,�^2u*�X��[��ki��$��E�.�R}\q��58\�N�д��w(���Ɋ��:Qw�& ŽE��B�nm����4i��a��rt��=\Z�.;+|3���
���'S1��	�)
�T����Ƽ�=��}�[��������/W.|�fƑ�����I�b6Fu$4:jv[ܘ��%�:؃v$Q�P4�,~j��ܾ�čU�0	t7�\�w
{a
r�2>넎9R�V��@.��EX�8�qȪsw:�v�	D΀9��F�M='���̤DVA6��2�K��f��0�b��s�Q��#��rQ�J���U��W=]n�����C�l�:t�=ӽ�z����S��;	�����KV��&�U��*�3*\=������]x�G/9�x���f\��F��kn�t�Y׏@|��6�nl�q�g]���(}��y�C�vѯ
��*�D}7������c����r���q`8&��}�*�z#>���wp�g���<M1\=��4< J6_�z�oOob▉�??��	������Ý���s�:�䓱���׷HG��g�/w�o��.^Uٖ+����^2��v������O�z�K�ru��N��$2��3i�c$�t�M��V��{��]ѩYldW[~w��,қg(���f��S��G��6x���\��YvV���M����v)��0b�^wP�ռW�p��c��>��iJ�e��RA��vKkS]�r�AN���=b�\�BP��p.;b��sx�9�97J��2|CЌ� 4W-������'�/������<���ᮎq�|������%�+
S	�z<7)c�kHfU�t�g�+�ε��T�KlP����x��K���N�ô����+r5�&#>v����bFGN��*�\���^;�gv*�xɎl���Dn
��R�#x|���Kk��g�K�/60����K���Ĥ"���%�T�DS�X�!u�1����n����+�$8��>�s�ۨS
�<oYU��.��i��]@��
�|�U&���1z��3��ϱ�৷yf_&�.,��I���M���� �T4!`y��hι��u����_}��OM��5�t7h�zq��I�"�^�0�2=�ޝ�h��-��ʬP����y���6�#�Z���:f��5�)7p)��K�.�H��A�nBsNfzMq�}��)����w������,:�h�o����D�A����j�I��I�Cw2^ľ̓1`�P�����8�Re�3�|�{��Rx4<fIO�s���&ŨNJ���\�\ �[4���W��ΨN�����;�����k��i��MR�$��_l`��,b��\�S��pb7˥�X�l��ri�e;߮��Ve&��c*��b��q���#Ut��tña�N\NF��Tf�u�-�Ź5-��ޙ���}�w���y�0zʳ�>iV��^HJ��2�������+[T+�:���
<�#�P�S�����k�o���X�u��L�
]Oc}�i�sk��u�
��ʡ�T7X�^���\뻩�M�>�8�+b��vLd*��P�ٖ��K�Pl�?yE����ȕu��]1b�0�B��:�ږY��ogjyI*/1r���ya�&��L⽢��S�x���+]H��;-U{��O&�#���0���x�>T��rP��<�}ϲvw���鸘)ր50c�fx�u�#1.F��wTW�]]�3��>u�3�܌e��0�+�>��E�:`��A�Z�_���\�l���(h��n�?���j��"���!�v�v�c��ו����������l&�I�d�ˤ=tBNHO�U�o��t��������Ѝ��N�x�냂'jqD��a�w�=}��:����WEEW �p"Kv���ڙȬ���3I����V�Z�[hV�ng�f��VG� e�zI����m���G��Ji^�j�+NYg��'g'g�N�S����xNr���%��m��gu0V��NW)&7Z�g&�����Ž3�=4��Ҡ�t�-T��#�9�#�/d�Nsdʒ�]��ۓ�f�O!�}��k���rZ�lS`��{���V��ǒ�I�{ƃ�<i�����JH��|����نĽ���y�8�&*��!�"%0f7/�m�)f/��Y�u�T�)�Rc#�:�#��'Pf/��Ux��$QJ������sx�A��{�~��,U���&����]	iћ��Iࡑ	�G<�W}O ��I�T���.�	&9t�\N/���4�GX1y{�\3#A���)1*���9�"��&o4T���V��fsz���.�q1��^�wOڼ�Ե��A8�#E�rUS��r�\�����$�&��b�a	t,�(w.��hRr_8�.�l�R�'�jyˍ�#.���s�d3��=���a�.j��U]�ݦr�&���Y�0��Pɟ��y�ۨMW��(��z�:Z�������z�C�We��α��ώ����%��6>�S��4�O�QQj�/�*��j�`S�7-T�s)}=p�/⨰�o�-0f���Y�ѣ$hu&c����Ay���b�c�G#T��~��fR-��d�mn��͠_#�R��`/������L�	��U����KP�W�u�g��,��:����۶�Bd���n>�w�_�:�gQkC�Jec�j-a�R�Q��5��Y�}[7���8R{�+��+N�D�\��7��e����y�Ra1�"ݙg,����J���ڔ�yd��t�If����ۤ��^}r�.��̞���s�Zo����;�{^;�n���/wVK�gz�}�[� �W���D+��H-G2)���ƺi�s�"���v��E �۫��o�w����g�#n����Ɏ �uH�Ƽ*��q�_�e���E[A}i��9Ϲo�gK56C8VE�	C��13m؜n�� E)DC�"��@�%�	3�ܾQ�~�W0fƐu2v"���lHΤ��u1p��꘩�UA*��1z��(�U�	JMϮ4	�U�8�����d}��G�a�L� �A�,u��5V%,~Š� @�}y��|"�t����ω�/>e`�9��֒��ָᒲ�일���I.���:dV �:"��;�@��G�V|�=ӕ�P�7�Ţ���Fء�B`Z�N;��E,Wt0�eͷNg��:�a��w�N{l^*%�Yr�'�1�v��W:~cIL��V���9�*f�Q�I�
����878�1�\i<��fb3)GwvpS�5���>Kf*�Ǝ���;�r�Wݵ�c��v�q30	��}�Y`��>4p�j��aX�ؐ�T,�,�E����N��T��!i��}2��w���"�9(�Q�R����gy-/��g^�=�4����xTNKu��fEB*3���2�*����`�Ɠ�}���茈I�aw;L�q�
9U����[�o}I�U�x�����Cm��-��(_K_}7<-��s��d9�w\�ߛ��t�26������U��'��Pk�}�@f2�*C�1^2/����.�>S����_����rF��s؁Me��r�k[�������� ���Hhg����?,�{�Q�wė�?dN�Bh�R#ۙ�\��t�Q=9w���T�^pxn,Miϭq'KD�!W��P�\p�!�K�i�@���t�Q���r9�6�GL9x��&#�s�T���6M*��'Z\z*�l�ww�ZŦ�����3�6՚�޵FC�XV��F�Tdo���9
pAD܂6%<,	e/k�<t�V'�/�6���a��>]w�;u�NL�����:�����w�T�����\�������!R5�Hu�Or�E_yl��mg�o=��������Y�8w
�֐^�)��Ę�Y�<黋d�ɻSX�bGu�2�N���fS僨A/ HY��u���h�f��4�^�9�Z�riP�ʆ��cx�N
oU��ZU�z*�|�ܜ���A��Y��;��8�1"�.]�W�hR�B众O1��Z3�S0B饓�Ve"�����{�.6v䳲�*�q�X�����N�-����Xt��>�1`�\v�7���d�v��v�V�P¹�[݆�6���^�ZY}z���"�6���'&�.�PwU��u���Vpf6�#i@��M7v9vW՗f���*<M�)��|,�r_A�Xj��;���T��dҀ�T�����qE�[8��s3n;�	Ly�-6Ѱ�^�#����w��X�����V����B�6��ͨ�\^w�oAt��Z`��0�� f��sR�s�M������S�{�=1�*b�N�+w��Մ�F���u�^��4��o�<{]yLi,������XQ�u'*�"s
I6��$�Ѭu s:�5G�p:���UcK�+���ǢV)**_3î�}}
=U����ծ�4E�)b��pؿ�d��_
��H�@�)\�E�l� yL.��2���]��MVU��4B�'.Ε	�.��5w,C�V�ڨ�S(ϭU��7b�miS�q���,@�f��y���,���c��@H);���b[��e���:p�G�����KZsAR}z��G�"�h��R�?���h�4�gg}��]]blN�,������������%@�a�qc�/�cV�A�:�醤t�r�撫��24���"&@)�u�3�=Z�����j�g�v=� *=�:�[��+��N�B�N!9i����c�U=���v��L�b�١�;��M��[���|��vN4`�]3X��c�A���t��H�����(N;KĨ�p�2DB���VKN���sw��|&;�j�K�q�o�S2�`mvi9��|����"���&u���:�ac�X^�d�Nr\+C��WO$1��4��.w��q�K��Q�Cv�Z��)
�	yxd�0H�Rw�����7�q�_:�v��S����9O�KZ%��y�K��Y���H�:|�l�8���;heK�J}�S��e#��u��9	�q��c�t6r��L=���i�|�� FK�t	%������)��3����^���&P��
��K@��i��z3�?�H:ڱ�غ�{��9'�g[�ڽ=��6�G"�
k�V��ț�f�T�jw-�*j��Z5$N��-��#š6Ѵ_0;8����B��ݢ;� �,�Y1�X+��*Vr�}Ǻ�,Y�f�U8lj�`7�u�2]Y	!��.�R]��L�z��jX{�D�dn�Pط����q*7m����m68��f�7�����5�e�����(��)��

��
((j �h)����(��������Z�$�h)��&�i�)H���
 �F�i
V�(hih
�Ji
R�)�Y�j�"�Z)
Z �hj��i�
R����()�JB�%��(*aJi��
B &h�����JhJJ �)��)Z�(JF�)J���i)P�ZF�)�@}�����s:�Wf���_do�&㼍R�G!����X���V[�nwbj�Y�}�B�R�)Ђ,��s���fb-u�r�o{�k?���}HV�5w�*���������~�k0L����W��5	]���b��Pj�{���s�>~�4B^a��}֩Թ�2<>��_���r{�s�T�,yxu�.3�ܯ=b2r~��*fc�FsNC�y.�^�͉��.f<����%;���k���d�0�HP�������X&N����:�C�j��A��>�Q�O��p�O!����Z;�U�sy��SK�}�T�\��<"=�L�5.�����u>˚ǐ�3p���<̽>ր��FN��������>��Z��ݎ��~�F��a웩
M�ϣ����X}�{�?a�U�ℭ�69��G�*�|�W
����Hn}�����4���J���}��A�'k`�F�˫����:�$���s��=A���:��u�S���%�j_cq�k?K��	7������Y���_��?�;y?ޓ�{_�R��}�.���My���>Z���{��;���?}�6w'w�j�>s{Z(9�S��4�����}����v��6{H}g�o[�C��Gիv�ej�C�4�9#>��30'��@f#p��y%��.@{�=����.G^����%�j����p�\�����;�2y.v>��K���	O��K��������4T�y��w���u��V-��θh�2~���D}}�9�����?�Pv{���5&��<�BU?I�3W�?A�K�;:�p�#�ufѓ�\�=���4��d��~s��(yG٭/-w��5;�����zz�U�v�W$���f"6\��?z<�.~�\���5��I䛩
vw���u���{�s�5:��<�֍�S��WF���P�OF������oA��y�W�����2L���͟�'�W~{��<;H{����ʘ�� LG��w\��5���4%�9/���y��z��0����w>K�tw�A�ػ�T�u���ujA�������jz��#�J}�zÑԝ]A���z��߻c���{��~��@UxV������~��?]��lr亍K���w>�\��|��w	Tr\���j����T�.K��j:�v������nԺ�ToX���2�#��;�S�_k:̬��n��ND��N����CE&�U¯�L�p�2��+��2��1t�]1)}��q\�
��ش�]�y�Hq���%$�F�z�sO�r �!�[�o2joJ]g>��W�$1j�{nZჵ�[��H�e�\]ɣ�8��^7��(�/��w�	�����u�˨�%v�ޏ��0wji���mz���������\�NG$�rѫ���7?G$�}���J��k�<�R=�y��֣�u�]��{�٣��z��k���8;�%��>�!�:�~�?A�����p�/~w����=o���|�K����L�������F�:�?}�1��aw��n�W��i)y�����P�s0:�!���u�A���:�;��2L�fkG����;�#����K�jNϼ�pu	o9/g\������Ϻ�ד��\��y���g��9��>��Ϣ{�x��������|g�+�>��}0��G�Sݫ��O��%?]�q�5}���
�G��f�/�L��ϯ���]F��'�b���_���J}��G?d|�#f>��
,�}��{�*5J����~���z��\�=Ǹ�}/����������Q��К� ˸��N���L��C����������`�jk�a�r�A�>���\�~kD\���1鏌�<`>�E�j(OfE�w�߼���Д�=�Qן��p�=�����K��������Y��7=˚�Ϲ�K�>A���5�	��?a�ܺ���j�ܺ������EO�3�j l����]�ι���Ru&H~�j��������ZCs�9:���{��j� �>�ݽ�'pjC����� ��`��j5r=3�'P�$��u��v���7�q��v���K����zjO���w�ٺ�<��c�u?��}��}��˗�����/����t�����=�{͇Z�2ya������j�>�G�r;�V��sPP~�W����<٬Y�5�QT�'Wz��W�0}��Q����X�����n� ��u�pj�l�^�K����'��r_-OQ��zJ���z<����P�^��/Q��L�L��]f/��pڻ��o=�a��)YR�.~3�����=����K�������ܹ�!��5&��=3?F�)�=��ޏ �BQӼ9��~�Rv{ޓ`d5��O}èFO�s��u�����d�5�Z�~/~�XQ7�" j`���l�\��)�n�6��K�
�[�L�e��u"o:����&�������,xt�2�{5�d��6���.�Cv�m���-v_�"��4*�X�L��X�%�pæ��%MLh'W��Z���}U�䳙I�k�}���D�}��E�	~����o�2{� 5yj���ːy��rnL�;���~�F��'Ff��2}�����A�u	O�a�?������]i�I���~����v�6��
����)"��#�11���~��#$����Q��<������%\��5߼��P���w'q���!ߘr6K���O#P�k��~5�5�ݨ:���L����翹����]׶<Ո�%Ͼ��3��#Օs��}�W �~5��KE�sg�w	s��Zz�nC���5��Й?���0��}p�G�߸�������K��������j_֧��;��t��r����'[V����}�'g虊�U!C���Z��^�^`�f��]�/�Ѹ>ך�%����3ζ��r�=�5����\��@u?G$�{?�u���%>G������B^]vk�o���W�w����.�����9jO ����d5�}�&�=����0���]C�w�hܺ�d�=u��:���_`�sA��\���s[����.�ģ�ܟI�<����r5��7����]ֵ=�W�̔�,�Ղ>�?9�ُP���=�BQ������y���U&A��oXЗ�<�[u�w���d�yގ��=����Π�%_b���uPd%�}��k��|�'��u�����z��g.��^~�����Gľ�Os��h:� �q|���k�����j�x�A�0L�n��rj}�K��:���jM_OZ��U-h�9��K�N�;�u?_C��}�{;��|��x__�p��>ޘ�evI��IQ�d�T��33w���s���`kXr]T���a�����j��h�^��y=�`uT��6���k�C��79.f//cq��O��`l�>�4�\�z�k?/нj�gyO����g�5V>������wЙ>G�j?}�6?Gp���|�j=��5޾Ѻ�C��y���`d5�=�ͯp����5�~�P�<>�s�sY���JFK�p3�z;3�Ck�ψ�C���?T����b��))�z�Z�<�cR}&U�`?�����ݏ^��>��7�6� �j�Z��N���Fs �I�'��A�KX=�Ѹ�����fk<��N=u�����FY�,=:2TY[&�<S�$�qc)�]��'c���K�&o0�u��o�r�'VF��G*��N4�o���K���r�Y���hQ��B5���fu�t��ׂK�Y�ř�"����yG�%(��[�z]������Cy���着z���_{��I���>۟��=A�J����9�Pd���ϥ�7=K�o��~��y9>_�ևp��.s�:�
�����y}�d~9�r����5'�kIO�9�W׽�wq�_o��:��s����P�KE��A���-�ט��mC��:3��)��N�0߸?��%u�h�\����wޗa캩����>��K��~�s�rA�fsݿX� ��
�k�=8����~�!�S���}w�u��Úӹ�\�_o��Z�BS�\�6}�˩�R�A�q5����Fc���?G�k�֎C�:���h�N��<�R~�&�y^I��F�}�@��g/����o�Y�Y�u�|;��c'�}��w.��>�d��d9�nA���k��b~�sԹ�����))�6{���j5'�u�����<�GZ��;���;�JPUAV>���J��PN	�����������Χ��������2z��?����߹��;��P���Τ�29u���kI�	W��������}�9�˸��T#	|��K,}�
�¨��W5�T}Ε�mn蟹�|�|�
ڏ-���	�{�o��jMO����S�9����A�%R�������B]��:���:��y��;��_cߘ~��@ta�
c����$��o�^�UK(��9��=��~�uS��X4q����?��~��f����
:��9�O�T�p�GΟ<�J���s�:��^��u4I���RS�G,��������W����xl�`x^��:�_}����[;�ǳ.e���kB�q�y� j��{\�q������5g�pmR3n��~&�,呤�K��]2ޘr��.1�n�C�s>�pxnR��m��q'KFx������(�nx"u��L�[��F���DZCMP�G������)8���b+�Ja�M���f���{{��Zei�6������������F�7�{�hb�s���wЊ�K�T�f��S����+~3�O��f���W��B��S�섮���
����TV$�������Nd.���^漄�dC�~�+z%��K�xu�Ip�<�p@=ݣ"��aB�"��9v�V 0e�sW�dl5A�GO�t���)π�I.a����w�}S!�޷�m;��K�K��Y(��|���x��t����]O����M9ֲc�r�v�|^'�L�z*x4t��(�9��BF�H���r���N̙t����7�����MŹ���c��]���U��dQAx���*;���FyFr�Z�=�Ҋm�Ź��zޜ�o���f�ʗ�1p4�<�m�V�˓E����l���o�=�r1�u��¸�7iif�r�K�$\v'p��mِ�ә����r\����~T�b��ׇ^��.i!Q�N�0����a�L����5bo&�L�R�2Lŀ4� j��fm�֣��eZ��N}�د|4[U��vyo�]q��<juI�X��u��ґ���w��u�(�:p2s�t�7���@u�W]�;y�2.�&�ϩKΫ��9[;�.�P���Ӎ�����!��eoM�Uy��m��M�7�w�g�)ՂE����l�d1��.�-���>b�m�s�;���-!�+Nζ��� �x���h�|�S�]��-�9m��x`;��3�úv�خ��JFf7�:�;xv�It�8>'n�Rн��}�&�"�KJ�K�M�J(�Ъ�#�U�7Y��`�����^P\��������3Ԧ�
4��i��G�r���aڼIN�p��#�O����ƅVu�)���YRlB@!�-��j����V#N��|2��.��u;G��4곪9q`vʈ�0u9Y!�Ң�//�%Dwc�3Q�YCg# #83DJ��W�
q��o�� ����2]FW4"�;�dO;r2 9���`�o>���ӝ4��v��+YS[0,z����p
���:����q�ʘ�s��tg2�g,��.�:�ïu�\��K����Pc��$�W �GU$H�qN��5%]9َ ,ؚ�Kr�{5(q�4a"s����-Z��A�y�ݐCk���Y��6��^Ǌ��m磻s97է���k����jY����w~�8!9�@^��	�G��@iP��(I��
I�|��4֤���q�ެ�Ƣ/넝�5�t�b^�H��t�:�EUrD�7E��ꙃ1ZA���]G�Ee;�ߔ+�x>�Ư�G99E�\[{"��3�����n�XT
���B�w�M=cFu�"�lq����!���f�F#ɑ�����ٔԨ�@�Q�s��^�� �WTHhX/f�u�#k�j�k!�R�;����λ#.�+US���>����UV�ș��1�;�Sc>�@���:	�2�DX�{��ٛ�U���G������ �����P��Uyc��ʠBǄ�[.�.ļtf�E�Iࡐ�Dsʴ'eFX��m���=���:��*�� o��!��Y��7�YR֨O��S ��U��Q���N��a%�%�r]g '�S����h>&o�t��{����q_
�H�4G/�)�����;�l��ѓ��L7��!����E[�hS�������<~��%�/��S�����ђ��ǩ��fܯ��=u[	�����m����Ԥh��`�{��R�u�6�m!Vd��vD�H����5U� Mα��ώ|kx\�F��s�/=%_��V&7���vQ��Nj�]Tlt�W-V��s*:��9�!���}�b��Gۇap��q��r������\�3;[�bf#�W��5���52�ɉ� ��®н��;��ix�ߢ��pO}�e��,R��rTM���(��kJ?(.��˛��%�Oh��v!D����H���v<kD�ҽ�R}v_���N,ꨞ��걆�7.��hqǘq�Uu�f��<�������u{�c��n�;�1��Ƶ�kչыr�CI�ֺ܋hD��6�k@���%2��YUx�8.�7�����Ϋ=۾B.IB�d�U_}U�^A�����It�
s�k����y��W]''(�6�b<����+t��|�{�Z���d�"�4|�;z6��vF��zn�ё�\���Lu�:G�;d3�.��XiOT��!������ȁL2�rxl'S1����ϝZ��3���ĜC7����v�&�TlHN����S
�"�2v���l��Hl@u6��|�3MN�p�_�ۜ��m���R=����D*FtL_�ÞR�|>���*v5�����V{ak��e���j�jg��ebMT �����_ٔ���&Լ�V	���R�LG�m�z�Z���ϥ��dhgy��wΦC�;�C���BӐ�a������!ԎW�b�ó��;�{N��v�P�-[�u�yC#C��-�O��t=��/���Y�b.���|ww'r�ߥYHy���T�J���S�й�ʳN>��Z{�8Cڭȁ`˅��x�f-�]��kj��5��5L�`1�Ry<��?��^�G�=��/���
�C ����}��.8+�$��jU�.�ŀh�����j����.�G�g�T�l ٝ�U�=c!�:���Tx8�w���[�K�1�a�%�gI�Vx�v_fc����z�:�0i����+�9�K�DE��^��9e�;tK�j��$�`����꯫����7��������1ҿN��Ⱥ�\��֦o����p���)���k��͝��cP�n9�7��j���m�_q��*�xZ6���`	��.�,T�8s8HJ���^R[�K��p.��~H��{˷4DЌ�ݡP��������Վ��׀���|�zv�Y?9�t&�1Qn�C�s")ٗ=�[Q�P�,���3�հ�{�ʭ]��s9��n�EPhC����̅�D�o��=0��F����Κ��9# �!H��f���c���՜��rP������bT!�SZ��F�A�F����|�K��'��MyuL��`��ڍ$�{�Hv�x�	s��7�~�~%㿪�ӓ;8W<H'GA��٩�Y�Q8a榍🩺3
������'��*���C�J{��W<�8 ϼ����!>S
/�q�3�ܭ�g��� d>yJ��~_q��T wQ�h�(̖�n|��.�yh�ZQ����<Z�����<s-���`_ɻ震�"�%�1?.0�!U.��}㖫���^�\��wt��Gw�8�cj��%xu���f��<���g1$�m�ݵ��!1x�UB�0�_V�[�*��HH��z�Mڷ-ݜ��a8�"�8�t�%]�ᶫ+tc�y�7\Vs�]4�uK�Y
�Fvu�=��ﾯ���%˴d���ZЯ�3�9�F�WMِ�"]���c�����S�����r'kٻշ=m�y�߽�+e�m�����Ry�&�M������/e�d��f��)0`CN�O{W@�^���LxX��e^j]sΨ��7���Jƭ=��Фv��n�6��U�aC[��6;EhP��+�EB��5�X�פ�g��o'%�AV�ØD��$3)��q�%C���ؼ��K�Y����Y�w,G�������l��^/Eu<4��saĹ�-�0e����+a�,FW=�b;��f��2�r�6Ў��蘧��6��OS�޵Z��3�`<�����D=e�N��l�_k�Ȃՙ�9]7�[B., ��ob�d�UG8�h��U	�qfXϖTCBx9FC��E�z��NDwd;�5�ue��*�����w-�
~�s��Mz�������������#N�����9��Xz2��ض��Ɇ�X�u�Q*{*�/y�s1v0��Ҡ
��\�ܷ�.��*`���������Mǻn��v�2�3�֏u�������Z]��d{�6H��/���S��i�������;V��M��1����;��!b��&, ����蚄���IHsl��y2T�f����-v�H���R�ܮ��)��T�tlX9�J
Ԯ���4���#�N���B��a���'�l���ww}F��۩����N-���37������+��*
�L��h��saKw�
��DV��Z�M>�'M����.��H�s#o��5���M�]����;l��)u�'�K��7xm�Xsu91�l�u�EKb�k��L�ة/� .��+���;��c���Z�Yu�qa���Pa�4vL���<�F����v��VGj�A��RNL�}���v�&6�f�=W\� i��T͙H�(�3+�dAJ\4��f�rV0Un>�A�f�I� ɉA���Z�6Q�m��.�����do}Y��lj8�t�B�^�ىvV� h;���\r�[��DKNo>/*P<4�:X���Yh'�ˆ�ն姢L�+x�ɜ-���s�C��+H#U�h5��ݶ�˰��ڍr�P+�s.�d����b�Z�U��%f����[[��B�t�oV;b)ϞH�WG���*U(e�ݸ�4q��L˕��*��8���ۂ�SgtS{^c� ���Ş��n־���F�樕+�p��Q�H�I��qŪ]�6�@p��F,��.ތ�J���Y&:���Fk��M�P�)�	%f(6�}n�WPj����z�_re�WT�2��t#$��}y���٢ �
�^^�%�K�6�K�Ր��84�Ƀ.���A(�sbl6i��!��̗�aޫ۔�F�R�̦�:VPI���qƵ�m#ӻm�ܗ�N���\�;���,�ڴ�|3H�*�����\�!�G�K;�$}rK�vZ�צ�p�;�wIޮ��5 �S%.\Л���{c^�+ᆊ���j�y;s�B}�S���efr��[K<7pX�)�{�6���\�e)�j2�;UjiMX�gv���£un�e͚NJ�q�n����{t��^W2��:al���6R��k�*n}1�\X�Hl�����޼��G�W!�#�ϓ�1��l]M1����ʸt<��V_����Siq��P8�E�j{���&�*��!&�Lsxٮˎh�|���QeJc�c��.�u�*@��v]!�bC���Y��;ՙ}�0�����W�V[�u���
-��|������2�S:�1�DRm=ɝ�=躦�}|�p]&;g�P��e�$47�o:�ls` �ip첀�bJ��{�s-���q���f�3y�Ϣ{-[���c
�#�K�םebD��0��3�����֛wx�LV��CZ/���Xi�S=����ƫ �R�%�_J��<ֵs��웮�_'L�Ҙ��C�(:�[H$�v3�d�5�{߾�_�ȥ������������"���$�������(("����(ZR�((h��������

ZA�h*�J��*����JD�@�$(i"��
R����2�h���(
�(�2�r2
�I�2Ȫ�Jk%ɤ(��������
j32")ZhJ�J
J�E�
�(*��Z(
P��b@(
ih
JR�j��' ,�(�iTȢ �����4>��r��lwu��M�$�O�k�g/�(���i��\��켚�������.�u9�S����e���h	����꯾�:�s����C���t�Ϩ1P(|I������>5P�]u�[zf�E�0���.�3��u�#b9�����ЩT.����|Ί�4�"D����3�Kym�Kf����"�![�3�m�;�����yP���<� 4����i�Nȝ%G����U�a@�Ղ�z���'iu]0���d&�fK����Ds)��v5��K-.�� ��V�w[Or0�/���i-��=�f��f%^̰N�:�ފ�Β��IT40�)T�Ec*�B�	�����v%�f�BEءe@!���5KV�R���m�d��ɥ{c$�M�'�����+r=���7�oRʖ��'�gOm�X(��)�R�J�Ρ.��n��������x��b��An��/,�r�
�k�H���\�R�fE���Hl�h^�8��s���~Ts˖s����P�O�4�Ic>�O7:�otW$	{%�5W����1���1�oa�12������yp7>���| M�#D/b�Tb�jR+7��mX��n�J���y�:�*=����-��7V�P��۝m0�u��ف�]��j�����݉lg:�'�&��e�z>%VR�8"w��Nr�8i�gz��Y���d�����'�Et�Y��gL���꯾���=����K���k��"��|.�QY�e]�s�v6��kx=Aձ*!�)T�;<�{��f��J+�z|.��뵃�`Z�j�u9���`�Xr�L��[���ia[*�v7zD\h�X������h�S�|�φ���7��N,�������^�u��+T�d;�TVCO��q������(��^�q�Sg��W��Ǝm!����z�G����w#]̾ϓϟMh�Bх�<I�W�G���b�˖ud��y;����븢=c�>AS��5GƷ<��Y�������"e� �Jx�q��p�5
�s.'����Y����5cY!�A
�����u�֬5��8߂:d�.�B�({Ry�0	��O	Ȧ���I�1��q��2�z���z��Q��=��`$�e�I������Q~�oJ$}�#�`�B��f�r+�=�S����\$qʞ:�u&�nj�Ng-��j�087�Y*��\�҇��	T��S4ty���i]G���Ug�����^�\�%5D�s���_7(���Pq҆"�CM��[fR�Uw7O$��f�����>�G�RTmĉ��	����w�����8w�璋Ry�9�����QCbj9��v��B+;�yHK��VieT��	d�NҵTb�[��������<䨦�v�I��/���-[�g�H����P�;@�Ӈ�����:�AD=���s�MШ�4�d�^[����h�w�]���uy�Լ���x������TPE<��{���X,�<���#��l�u7��Ϩ1�/�6�P����	V��k(�0�4��K�ϖ��]�gc����3�
��@�� *�Loc'�n�ؗ�冚�Zw.H��jCs�y�)�|�������2���xzﲼ(3�Z�=���ۊO�U[��W�N��"/^�J���ҫ��x7iΉ��
�;���]�TS�=���2�\߯�{vx.�~H1n���Y>i4;d�K��jk�u�E=���3���Z�O^��w��&�ȝn��b��{n`�;2�W�{.�s#@�|�6����aɴ]Y��륞� �s%���.���/s^BbK�%,z%�6M	�|�a�5CA�;�u�ې8�35-�����VT!�SZ��C@1��|�n1vA���ױަ�m�3��V��N�&��:����������ff. g�P��<�en��'��,�r=�0ƫ��9��¨���}��YĠ���a�黆N�I�
�m�
�Qd|�[V�^��Ծ�bE_��]p.���m�����;2��U�������>�f�v�jAg�A��~����5�#8�k#t��m+⼻���ɝ���"��C�m
��g���3ڼ>�QW
�<\��ȋ����&���\�t�']='c"؜��9��2��Im��q�m� c�Dg�L}HD�U��I���f�Z�=������$���5��6�\Yzr���5�v �Z,���	��[��OKB�9��h,t���� ��i�����5�o�/�h\vAWMِ�%ۙ��,��)��r6��-k�u��*�[r41���[7�.Zc �DbO��M\	��R`P��̗��2PD�!NIGd�\�g���V�}��q��()�,;����iu���p�sr�O0��f�t"�(e�SU�9�m)�#���0��+�h	u�|.���יc*.�&�ܗ�2��q���3����/<�E�W�����^�^{MJ]:�u(�Y�лs�Ә!P��eNHƁFW?�'��Z��g4����oMÜ�)�b�;,FAus�7�|��л���ۢ���r��Z��C/���6�J��J��K��]�м�GV�?up�r��M/���L"����̈́n�(e^dg�&��3ʖ�AnMl[;��6�pY:�nS{]�u�v:}crc���Z�ꗯ`g�< U֡��Á����t�mN�}wV~F��~�#���)-d�Ɖs;>\@{P�d�/*Jʆ��_k�Ȟ�]KZ^�F�3��b_d�!�����x3������N�(����?3�RNVDHr������=Ϝ���uJ�*��%j������I!:��� ^����A-֗����#O�����!̰�?���|$t�I���܋+�b�xi�=Ż%�9i��xs���5����LƸ�ϕ0_O_�Ѿ�b����}y#�jV��s$u����DT���&�X2y!u��u�n���|6�p�Wz�q�6��\Կ�ӝ�K��ΧB�[�B��j8 ����T�j �KܕE���8����!���^;yr�dwBvd���&u�)� TH��# ��p$rY�tj#'�z̃!��L��K��֓�����llײ17��y���"�7}�w��A�M��ŭ�
ꇸ�N�]�ڨWxޘMk�G��Ü���n�>��P���N��~Ꝺ��8�M+�wX���jo�
O�ip�]�l��,&�}k�ƻ�Z���P�7tJZ����;;W-}zmF�c��pP<	����4�n�3B�c�3\/�nxڡJK�6��X9�٠c��jج�fDEN�&�ZIZ�]�� p�|�<��qsLN����ˇ���TiF����DD}�;J�F�Wk�P����>}M*㤀M��'����cq5<���oRʖ��~D���_���K����mP���O�yx]O,:�c@���ea��s�T��d*�{$���a�ۋ�#��?�c����犻s��3��`�u�H*�[B��x��bx��U�GL�f��E���S��>��U��_ǩ���q�ȗ����^\����p}<��2'�}WP��z�_S�7ȼtS��ʒ���1��hl��n�Գ���7���8�v%e:ϓ~��1��]�~�5�ټ��1��=o�tg���:��Ȟ�sU���;S�z��]{�9���c]�*����(N��؈�<��[}c�S���:�Os�8R���a[�[�ˈ���Bt�;n̳ �J���	wK��=�i׾��t�v��} ��%p���2c�%7�;|���-����>ޟu��o0`��50����5��L�-�%r�b9��i��̴q(�<������8k����Mv!�c>�ƀ��C�V����/u�͉jھ�t�"����5���=k�4H8'F��\ѷ���M㥽�Y���Sh.w�����N�ԭ}������.�"��Z�[W׻ܦ��������D�V�^�+i��ʗq�V�Vm fz�n�� �~�#��"!����ܻ����]ׅ+��O~�M�:C[!�A����'S1�]��t]V6r�H�_.���t�`X��P� �,���1Gq�ٓ��6#dgRC"|�:���n�״;�z/Y����Q�To�\��VZ���BFz&._:��✼��˙���&�#�V�N�GM�K�E�bf1��K���+��H���/>
a���"��t4�h�*�S���SoWzyJq�eJ��f��I[�g��"��{(�����v�G�)�2&����l�� Or��V}���ynS5t2T̩7Ng���s��}5i�N��&�MF��{)bs�~�V1yn�CC�J���fN�AE�˵[�'��2i��O���_2���qe��1\>�vU��j,�L/e��qr�^"��(r��������6geq:sh���p5&_��}��cߏZ�����F��㻽P�R�4�2��{ �>����䓦���׷\ċ�*�}�xe;O\����%Dx�Z���6��#O	���7�We�+DGOד5����]����hh8���W_�^�8�A�&w�䩹��X�o,�q�6MlЊv�0\,�Y��M�X�FئH�T�٩�L+=J����^���D2�wp��h����`�� WV�{����>�4�.ͷɕ
gٛ����x�f��<T;�@�+ڮ]��"�F|o WSq�u�>�җhH��>J;QT���ߢK̟�u�q��u6��<**�d����Ֆ�|I�n��RAz�	zw.#�&��M�X6��b��s���L9{���SV����%#[���F�ugsx��P�#d �s9��p�]�ue@b�[5q�dl5A�F���4�V�})t��gV.H�̎��]`�T�O �E<U֕�|��X����93�F�֍P�!�\�/��
7F�Ć]O����b��/c���!�m�{��#��u�-̥խE��}���ҫ���4�	� >�P^?p���;�ZM*S�3Spˣ�X�n�49Œ��/+��CB��$�)��
\�-7}3���U����$L��W�C��H�sl�"]a�`�hu�K>ssB��	�25�����.��8�@X�����{��<ؘ��1����O�Z'27BO���@��0(dCn�K��N71t{�S͝�vr�\M�yZ,��zM���H��7ي��^��ݞ�AV��uk�{2��3���1��5��qۗE�w ����\v�J�}�>���T���Om��{�����7�,ev�B��ͰD�`�J�1�v�&�˄�)��й�F��}��bu�o�f�Y%j�b|+(xX�ML?b��s=]Uλ��?[Y��M���r�֔)|�8���;���C�Z3�"d�W]�c��^e���I�Oo��I-�I�U�3��y�;;8�vC��r�.u��x���ʭ<N�?z�F�k.����ea���q���Z��U��w{�^�s�!Lk��� �S�7G���s �P����gO=�x��gl��R�}5
fh�/jueC`d:�_V�
�tc*�=׹�W �?d�J�=���8�,d����r���,�,3�s�'";�\b]]z��h=iu��=V}�՟�d�Õ��Uۺ�j��r�,�v�d2��*%K慎�=�{=B5�VH'����:�WBOȃ���>�ַ-�˴��|���ɕc��d���:���?5���Q��Z��n��:vǏa�b#]��T骄�Z\�
�l��(<�o#AE'k�MN;�;9��#y�����ЩT.���|��*�E��2<x�޻����4� �*	��B8�er��f����wZa�Z�!�X�Ї�H���P�ޱe�R��V�{'�Lr��2W] w��X�h#SX���0Bp[�m0�-]iq�we���Q�N�=�d3Yۑb/7��N_eh�G���C$a8����D�����Y�o �@[l����#]D��;|�+w�KYG[����� a���nO��î�k�m�&��StGL64>���	�隮�pj��lЋ�]����樀�'�X�~�.�#����}��it2�3n=K��ڪW�n*EH�91�BW�����|hiE*���k�x!c��[R%�v%���7ky�Ш��T9���T#��[�A;��}>}MI�:H͆�/=G����k��X��K`�����ᮥ�Nwo\ce8;��N$�*rSꭺ�p�%�Wԡ���6�]��ڵ�XV����[�҇l>�+�g�L�>��]�c�̥�`�~4����)քӘ�욊�P��O�����%p�/m!��6cd�Lf�[�%���択YGW�kG�1�~�

g�E��?^N��}�r�A�&2)�U%d�3�Jb� �7���f�X�|ox�]���6z���Zev;�8u�\��7]����R�:4�c܆����^��\g�J'C���Y�v��w��k����!y�V]�1�U�u��1����Ϋ��=�*J���\+ۡ�3Q��G�_c}����c�.O��ع��wxp��S�mGRNg2#��$���8�D+Ut�r���g���aŧ��jnX̭ A�WXkm��P��]]��Lۊ�/x�2�9��kAX ;\p����mV��� �	Y8ڷ��:���Lͽp�#�s��U����{'�|@4��!V�HI��Z&o0P]��;)jۄ&8nۮ��T�dT(�;*q��ǁO�kks�^��X2�k�@axJ`��ƀE��Ӷ��v�
��K.�7��G,mv�X9�BvU�v�[���u
�,hf<B@y�I}�KO
�f�C��Uz]r��8�2ȥ�c^��U��>�.X͝7�{#вJbnKTB�:�: k`��z�7��e �k���Q :�PWIٛҢP��O7p�;�L;���)*���J+��҈���C{˶���W���ċol��Ѻs��)�tF�Ki�2�oZ�u�%�˵v���$��1�O����K5.�����U�1��j��E��C�]��*C��J���!!�T��{�l��஡��PV]9d馛�vo�2��jIoNK5�G/R�0�u����j��Z���Z\��l��ݭt��f�(O����_uod�KVa������5��T�Hv�z�K�݁�g5#F�S��:�H�����AU��f�W��
7����吭ȫp�E�+�&�s�!�eѲ�_c���^]�en���YQ�-�.��֌��f�m�HK�~{��g?�Q�S薾7yR�L�y�·���W�R�+f�v)p�i����N�-*�f�4����hJ���ZR�����cJ�ۜ0;�7y�{�D�������
��l����Z�<�Z���*-�h'�k��a��h-�I5h�7���ڻ��Q�(a񇖼�V�Y�\�gÆ@pv*9�_�6b��u�l��pƺ��.w�p��&ث�w�4۲����W\y���@t�W�����V�f���3�y+�M�9�����)�\�W�ţ}�Q{t��Ц��cJP	�ŽVxT�j��v�'H��t�ڙk/�����䚈K�q��ٕiHi��5��L{��1���rQ��ؾ�����iu�*��)�`*����ln�:*���:��O�s%xi\�$�ڹ�J�j����lmѫ���Մ���n���m�Eu���%�����u�BŻ���(��[�ޡC'q�.E,-��3�U2wqR�� �]whS�=���[�n�i�Q

���]���Li�^�5��d D�@���;&^�	���WWS�mȑ7�Coӆ���ڜ{l�W���9�Pp��&�� ��n���(>���CJ8m���u�.��H�A�CRvw��OW�ۃ���:�"�8krWR�fEf3Ɇ�O;����9Y���C졐NK�M.C��D�J4J��E	��$�CACAT1�DKJUQM9%&B4"e�MSBP�P�� PR�CBR�  PP�3D�J�@�A�Y-CT��@R�ҔQBP��@��B�!KIe�KMdRS@ӓ�RUR!CIJ��B�FI@dd�dPR�@�C��KABД�Te��Jddę S�LJe�Y	M4�EU�o8��!KGL�&p;��ٳ;ik=݇P�݆W󮅸�:�%�y�r�M���G%lb��6%�����7ȿ�����>{�^�� �v�c��[�\�xl/�\+��\-�
���4|)־c�*ŻN�l9y��K��I��I7��(t�Bt�;n̳#�Q�����YT>��ǲ�9�Ӊ����E�B)��e]����N`���̘[%����w5���O>|2��LXi ����6N_F��N�p�k�MUG���[!o��E1�a���+z6��vkۿ {�E����>jU��:�I/>~���5?��
�yW�?��q��s�+j�Ц	�9:
u3U�n��͇��]���udU��`I*���=!0�B�\j6d�'���fͅr��f�z��jܺ���Q��&�]y�8�ܶ�_s�j!#=/�xn!N]Zr�{���ڇ={7�]�>���˝�M`c@�`,�w�TB�qW�sU�8#~�.��7�	�(�\"�>�/9��s�,�|��rʞ�u�s�B���m����࡚����[�f��oZ�� ���{!LZ/q�j����e���9�~�ד�/�9H�V^��g����׍�f�r���4�!*�3V����mu1��1 ۼ�[��w�hݻ��+�{Kc��Z�v�X�!#Y��8K��F!�_wC�=囬9#�AN^"=s(�Z-�{7gPj5���� B���u3�DG�C�x�Iz�2�k$ѮѶBJ���:�a��^��zP�F��J������i��;�+�x�}㸖_ƸT�k����,�:n���4��Ӌ>�UD
�����!x���y���R^a���&�4���irD�h5&_����eE#ə�5���;y�ҳӄ�
7�v�u/ۙʸS�e�~�!#���?<�+� �|n�_½�x�%x��[��~�r��C7fT��f����N�����v��Y~�%�b�5](�ZM�b=.�Z�d������+�E�\�0��7B��kbK̟����M���t{��S�.{ko�(�_&�B��<7{T��nM�.��z��ɚ�7An���m�|��7��^�k�LFE5ny�.ȳ��f�|�o�46�Hp$�t|:er��8ӝ������\"���>����Z.m�)��.O\��?EP*'8��@�TO �S�^��~��o|W��4/9�ĭc�'���\�9����E� _T�e����p�a��PA�D�k���R��ޢi��gMU�J�`D<����=˗��ާěCSi��wE�BGp�R�
�;-���K	�M,�#vU̡�ۘ/�µ��莗Y;���X�t��«eɸW.Ñ���z���w>Ub�L�f��k�9�s2��h�K�S����쁍+�ʼy��ꨈ�r�qO8���^��4���7���N�<��L|�%�&R���!��,Qx�����\r�j��ʖ�A����'�&�L�DK���&�]����#�ʺ�Yw��!*�E�߳��&��62R@�W�и�vA�� 4/���~:������xIǚH�W,'��/�õ`yTX�:��y5'��zetfO��Rw�]V�9o�i�I�Y7d����T��,#´x!ٗ�v�ttv�����QH�Uy��`X�v��V"oDjr>�.{��}�a����Z��`�B��8���;{�1��h�7ݯ�H�����K�.��Eԑ]};�sR�ۭ(�3#tB��»��'2m�m<iV�Q1��l���̜�p�!
cX��=~�2���,���O 	c�O�N��ڋ��=�]N����r���fHb����y�|���W���=�(�B}�4�19hZ�'d~���n�4���1pыj���,�W�!g�U���(��|�>rw����znNcv
��0A{�r�g�\�KR�#Oo�׽S+�^-ޅ�}��z����٩Ԁ��8*�<�;Zm_%jXg���nd�1�L$ �n���7%��� ����4��\����}K6Ԇ删��ݞ6�G���VL�m~����3����*�Fߡ�t�gVP���@D�΂Z:��o�UԾau���X�?���B�}}o57��3<� �-��ۣW�C��.�"��@�W��-���k��.>U�+N�1��gr�PC���eҜ�2���C;�c뉹�4C�Ep
�<�Us�^�w����X݉��-�X�^�=�4�:�}^���GK�Z"���ޮ���(d�´E����ˑ'�jk�&3�y߮�����y�	��ʀ���ಷ~I�]w�y%�C��㻻�������2���1�_ț�'I����}{"ͽ��=�ƽ7g�dpBAۿ�L7A �i,�����Q�[ݶ�KX@��H�ȸ����q�l4�jH�uX�<|�I���'� � ���7�A^�����Т�D3�OnJ�VM>�mWt�mob��t ��P)�G8U��d8��W���i�����**�[�8�4k�UU�[5z�ϔ��<ʙ}��!3wG;�l��&��5�E��3ϱ�Fq���Z�({�a����L��}�Һ5	�>|�vd��oivPv�}�3�*�F/���1@ڱn��ﭦ���f�_U�+���Ms|�7o�+\X�v�ɇ,ޮt���V)Rۥ��,]J̜8�I{�VǊwEmr�"���Ƹ�D>�M\�>�*Z2;)L#��zsE�s�Uۘ���;�$pss�yu0���n�m�R��{��/��n�I�;��b����S�1�����[���yp:*�#5��h:���N���MϾ~��h���cղ�j�t���Y�z����"�g	�Î���|Ҭ�A6N|p���X�S����.�	}��:2��cܲ�+=w=3D��F�����^���9��[�S��mU�/Q.Q�v��,��C,�W�A�eF{�>��['�_od����y+~�w���(v�3��0vݙg`V����&c���`��p�Ga]~�p\����w�wf��G�d��]%���qP�s�w2�ϟ���0�	ƪǹi��
�#;&��\G�����e��E1���+z6��vDk���Y�:�lAUB���Z_1|�������Dp9W�=5�z�]������1�UO��Q��Ͱ��&�� ����'�:��k̄���֕�<++�l/:8'��D'�Y��=θ�}���.JX��)eq�oԯ ƫ�3�����<�痝M��L�z�;`���j�X�Bc��Y����432^�g#ɳI}%N��j�7�N�I�o<���驵��T�]#{0o�/�y��7,w���C�IG��}���P�8Mե�`�D�tP�#&97p2�����=��_s����3�1r�ׇ(��t�l�b�����R�D}ɛr��Fx���|<��\��qq:�	T��6���_`�[��f ���r���i�Q�eK��Y���V�{S�/bo홨N��P�:��bDx�ݯ-k��glAij��I�p�ʅ=Y��B�E�)�����z��?�n �r��;Ҁ�x w��[�F�~���z�ED�J�vZ71�W�a����(t~ۿl�[Cst�k����.������e��P*6�E�w�~	�YИ^��N._,m{י�\g�����`��VvX]̱��Ub��.H��jCk�3�S��E!�����ٮʂ��Y�Қ\�\-Ka˪WaC���7y$�� ��n�b4c*�!^���י榮��=�~�B�V�ū�S�F�s5^*v'�N;���!4+\�qD@=�>�8b�	I4�[�	�ϪX
c8)���R���#�.1Qn�C�s:2�LV��a.;j���r����.�vU�ј���ڨ��RsV�Q�롉7���k�o��n��� �m��Tخ����ٳr������N�[J��c�����|�O!�ֺ��n�:n=�f�<`����	�r-P����nR����$�<4e�꥕\3�D}��[N��Ҙ|����j�kP�k\�B�bK��c��^���U������R���M/G���՝��l+���\���������Q�c�,']; �Tlq���m��D4>3��� ڠl]T��'�T"�*��9 �����Y9��4��vg'&��2T��.x��.��ͧ?m��L+���PM>d*F�I��qg��Ӵ��HG8�����Q����ɗM_�^�)��;��~��c�"P�	l���<���K~'c�~����S����̼��o��Żb;n:G\:"Ȝ�vh�M8Hθ�2�Q�v�A)�4:�(�p�2��n5�;�i'�s���fJ�#@zg�$5����-P�א�����:��;{z���].���B�/h�N[�U���ݵ]�{W(��bb�p)��lgo9��sN��o�:�jz�۸�.9ɨ��nwU�S�	S�RZY�e��}�C:?���=Vח.���r���l�1��*Ŋ���]�(��맇>���{��KI��R�\��nm!Q��p���+"�9	B��º�Q}�JT0�m��'��8����$Vռ�Y�,-��DU�+K�ݟ��N�z�����ݷ�������g��5�ZS�m��Fz�'��:�-dV���C���[;��TE�/S���~��RE*> �&I��h�4���S�MN&3+�|�++n"i�1�8�,dB���|Z�ܺ�-}vfݼ�������ȑǩ�lu�k'�+�nn
-��gB����n�<	qXJ��ƒ>�����`~���d�:=Ӯ�c:��B��kz�^8kq4�SO� g�iL�%�}ti��T��y^b�-l�h��3(?���̵���}q	��ڊ��\ɠ�'=�+�V� ֔�2�V�����;��Z���k�Gz�;*�I�W����8vI�k/��J}=)�S��\�[�NJ�{S���bb�q۳�*D�q���%��4'����Sa.����C���<�I0���z���a��OUpW~�f�D-���j�h]B�P�L?\��vU�Δ]:N����XU��`�5��[c&Sn�m*7+�3��H��\|�%�eA�\2Gg����s��X�����J!���r\�����ɜ���X)�5�����Rz��t��V�>�W��>$N��i��g����b�	F撎�����h�i	�#_G"��ƺOoFT$�T��Pqy��z�¸�H
���������[�bX+��S�ƻ��I���[�<�6.NE���p�7����eY����alu�D���ss�ҍ�P�Em=���7�>)����N����z&���VI��ݨ{�U4�5�67u�=�O�%��^��ҹã��y؞;	MҞ�����#��G?�l�N'N긬f�l�N���]Ց?�v魾Ty5iV�?����v�<�����+o��1�:���ܽ��%��&D�ߖ�9�<ψ��'�9a5��AC2]s��;b�2�ݵŔ��湸(�8�>�V{�a���Z�e^H�W��v�Yk�7���Ȼ����O;Y���(oSO�S/����S<�盠��x'"7��V�B�J�͔Z�ٮ!k]�\�)î=q�ͨT��G�_K甩��g��WI�ޓl\���<|'7�}޸_I)�&di�l�)O�&N"ƞfM���8oq)�lձ�=���E���tk��ec���Ao�Pd�7��#=q��+�CP����\��'���Z��90+V�Aok��#\>���hjj��:]�N�ސ�o/�^�?�]A$�Ya���U¤��kTk��Í-�hf��b\���m�QR��ʅ)9�	,�u��l��铛�$�Է��xn��j�h�ڣ5b� �VA��@K�\�2�\��-�v�o͞�4�W�>o!��"_l�nv�1P��q4��H����Ӛ�ީƎF�����C	�#z-g�3/!�r��j�(�:�ז�j�Pԧ�)M�.��3�\e�Մ�q�٪�N^|Îy���Nĭw�p��œ���9|�fyČ뗔n��]Yˮ!�!5b�8b�q��Lk��]�̰^*�N:��O�tw=\�J[���U�{U���ɧ�V�糧��Ƌ�ՑK�'J�}����I۴�Aߗ�����X}��+F�OJ��4�_�_��7�d͸�'��@�8<��ŝk<>5����Z�i�֑3Wu��m�v�4B�49�#L�����գD�[[�:�#]c+9�wYWO�T�W�-��rSK�Ӻ�%�6�N��	�Ѭ&�+z�.���J��ʐ�����"��ؤx����xY�ڗM����������݇ԶƁ��nNF�7k+2n�:�co��[�^�%�.�֝+9X��}��]y�J��pͼ�\�N�����.���y�^��+Q�;6d"�<���@&�X�73l�������ġ��v�;K�ƴ�
��`Y� ��I�w�V�eA��8����
a��/9�|X�P��eq��v怴�����򳔭ܗ ��5�/�9C9�.g!f�\����dS�mfՑev4~YI7�csv�ӯ�w���r�<�6s����M;���^b8��29PKwzJW(�7�n^+���f����`���)[��gvvX�g�i��Bq;Ud[Fڽg�d��׉�`�h��E�x���p��Kl��B��JcOs���K~�pD&8��B�	J�ң�ȦsI�W	ɖ4HX�U��^>5�aܬ�y��ر��y�l�Q�%��In�{�doE��)�Ʃ��Mͼ��7�f�8�����e�C�hH��,��+�y��1��L/V�_���#B,R����,���}kk��K����[S"ގ����[Y�p�f!�*k�����iz�J7�v����oNx���]c����JScZ��v�t.��P���i�j$��u�o3���cj�]�]\��Ʈ|�V����C#($�ǳ�Y1>�a�\rr�]���Av�{����>�r�j󜘐[9[Ъ�ɲ=FޡM\�ξ���I��°֚ʖ�ɹ��Eӻ�㔵�˥�Е���Gk%�lۍV�sj7���\�d�	�]�P��F=��:Ju�HY��>��.=�̓�|z�o�d������n��Lb�l.�� �P�o3s�|����W���O3�M`�ˆ�iZ��%�폍�q���k����Ng��%�	��\ցy�'�o����D�E��'h��9,$vÚ-0ga=����ܽ�^h�;�^��!fm	y��:ۘ�-�e�
��\H�bd괻(;5�����!?�h��@���܍�g8ƫ������Gi�)7����Ŏ��JJU{wZ(�4&Q2mv7�6���{�K�S[�0�ծX.��9���y��o\��I��B��W�L<ܹ�{�a�J���W���h��=�m�������[���pp�:��E���WPZy��B��Ru1��2ɡ��6:+4�֞X��<�f�!�!�.i5g����W�f�Pe�E�Y)�V�Y�Y]Z�C6nB��[��0ٝ��u@x���z9;�6���QAle]���F1����m�B��2�^��u�x�-�%]l�OZk�N��
9w�:1�j���֥ʾ��L�+�߶{羙��R�-P��9 VK���K�b�9	�!CBd����JY���9�HQB��I6NIT&B�M,M d9%&DC�de�e�A@�T��NYR吙%�dd�C��af)NIV`ae%Q�5Bd���!K�e@�e��%Y	����AJ4�M��	�9!A�C�C�Y��%���@d�5�19!��R�% dR�&K�f`d�T���H�d��F�[������2��;b�Iutt*[)fմ�制wJN=�{s�5�ml���*P�lE�[�{.'l᥋�Dw�ʎgf��T�!7����i��Ȭ����U�wB�ά�t�8�N��_d�yED^��Qn}����ԍ"��wS��s^0æ���\M�Z��&��Q�Qc����kJj��aM�ӹ~�W{��xHar�s��#�Q�޵	d�N�7�"�o�9L��QO��*�:��-mۇ�Ź���}
��u}j�\�g���k��opq�w2�����Y�'ZWd�' ���,����j�3Mغ��㮇(uB2��҂�Υ�t�ٮ�>q�m�yܭ���7�$�f�{�v�FE�j9�͊#w��L�|W4y�i�nv�%qr���2�i����������FzJ�lq��2XiC�:�O�WW���f���U��*VK!����J�a���&D���ڇ+�Du�M(~��<�3��^����iciYgC�^ɣ�7��C��9=te��V�q���:�L�H�E�"���wt���W׾r�VT�e*`'d/6�$����1y�Z�	t6�q���H)��4T�^�m0��7ܚ����\���^�X��"������B���y0��;
j�gh`��R���d{�����b
,Zl˴1:tr��jt�C��%.�WQ����E	S�W�������=�j�\��ݺ8��N��M+h���:����s�[|�N�Rcl�@�n��\�
״sb�=��Kt�|uvU���}��:Ƣw�=�v/c���q�Ս�����E]���1���bs�|�y;�μyS�\ർ�z�r���s4m��nոu}^ͮ�ң��>�|�IU����^�����U=ca��Aw���˓���uS��H�{���.'(s��vU�I.�+n&����*��B���}dD�c*z�O8Ê��7"/0���[.v�r��k=��T5����s��gv�a��F�g�k�W�!�לs�m)��]D�W�N�:�1�ō�<�Yf�iG�9��P��&�=��{��3�|�.�V�V�O��?���Sg6&�շ�Ջ��cf����O��@>}Z�۞0����W{��6���e*38��.��2a��ш�Sa�K��B�
�����mΙ�k�p�̓����L̾�q�g[�ʍ���2�%G�I�)���<��V_%0�� O���TJ�QWb�7�:���_ȷ�̵���}q	��ڿ�nMAs'���2��6��A�P�t�pC+Xw�΂���3Lc3��./"x49�W7���>GJ[7;�g8K]7���!�s4a�&z>�c4=9�s|���2/�zo����U�|����:L.3��M-��3����am���V����K훈-�[�)	F�i+��3F���Lw�8u}��Iٛ�18K]�9n��f^}/<=�U\��S��g�	j���<�j-9h�e�5;w�&ktӅˮr�6-$�&�Y�V�s�5�S���Ŀ���w��	hf��㹶OVo>�F�g�;�1m��/+�	�@M|F<�����ʝq8z�t��O�w=Yׯ"
�عã��'��a��,\�g�e�m$l[�;S�\��Kgr'�E�UOXq�e<�R���U �N|��(���8�V�7VkNQ�kW+��m�oZ�v\�C��)��]Gs�\�tG#^���=�j�n%��g/7>j=���Št���EnE��P�Il\����y��P�H�ip5+N����w5�x��Ahh����)�e�S/�0�y�k�B���\�ǳjC�3`<���Ý�����Y2�N�0��/b�uOF�&�~�|�|�'�c���s�*�x�[�ݱʥ�dT�ˇ;�Y���ak��:��I��v�d+=ذ�v�R̫Ә\=w$2y��Sh�7N�ن��(���%�L�^��G����Ut_���h�2���C��K>9�\+V�$����J+U�p�ts�Ҥ��� s5z�nMF��*.%��FXn�WB��>��Fm��#����@��^�ˁ���ΐ�Mɨ?3_Rsq�%��37����|��]X��W57b����k�8�z�s�)	U���s)t�r�򸫪�׶SնN5u�3�T�����%��lg:b��`%�OM�N^�2'[��y�z�7^~��L,Y�w��Yi��e��dKب�HQv��: �$�u�(�/N@e1-)�b�.���͜P0���Ԭ�4K�u�����;��-������X�>m�l��5^u��q�N=n.��Dm��G%vv<������byw���t^�s!���ι�`E�]v�A��yF��K��	��)ims�
��:�ow7X���(��Z=XJw�w�������"V�v�o��{b�`Һ��mxK��e����w�_��Ql~�OL�S�NkY�	\�����Y�z.�f{�ȼ�yf-�����ݑyr�
�q�_������-��D�lXL�1���c�e�o�_��g:W�G�5���[ʽ/x]�EO6T����~nR��M���Óx7�)GM�Uws����(���ֹ܇�*/Yy��s�C�e:m��aS���a�hfg`���{;y�>wY[qFϴ8����B���;O���}y�+�.�`:�Ra�qIL�qnS�r��ϩ�lu�K'�����5��f�U�~����7�o�N����y�Dvֻ���,�[(M�&���m�󜲜��Zh��q�4�}M>��n&��ǀ�������sG���yy��0j��Y��{LKC�v����κʤ��puME_os][���*P��=;�(1۝]S@�+��}LJ�Ial𵦵[�OSܝV�{Rj��أ�Jvھ�ӷ*V�7ۇ[��m����t�4y���#�k�	��*8����:%3z�)I1�t�|�z#]�}���EMɨ?3A|K�e�yTK�X:w5�od�*�0��_��a����8޸��n!�W�ܪ?s}/kV���'%E���*\�6B+u:���9iO�^���6N��
�O:QYy\PH�����Q.@K�������M,�̸v�:�%(��y{[��sە�ҷCW£��y_�="�U�G��=�/@�~i=u-
!i�/!H�0��x*�~�Փ NZ��l���h����q��^p��]->�%*�K�&��4�\6�D��v'b
�S��%�qEVuu�5{�\7�u��S<�ټY����^5��o<|���3��
]��.�z.M=�v�j�����*�b�����\nU���ˎ�C�o=��$��,������-���|Z�z�*���e�.��m�퍬Yq�J{xU�UY���x��T�c��{���w=����Zz��`B�t�!ڌk��6��sS�w�Ҡ�'$�%��O�>�Be�%�\�	��J�J{�+��^��伽{,<@�sw��c�����ܧ�x�ke�*�e��cN��У��=<AJɹ�������z��)�lV����&ˢx�2k��^4U��d������n^�@Y_H�q�5��V�OYU6���@/�ԼI�׉���u���7�j3��Zח��Kǹ��V�xGn�7����k>�nn1�z�|���3�`7�z��"��T�۝�
&v(Z.�SVv��g0+�)+��̵��Zi�@��nLP=�U�T�s2h��glT�M��Z�Ғ0����T��������sw&��{��{�o�E��/�]�%
�� �;�⹚?:d�g�ҭ����U��Y&��_���j���9��z8"�N��N�d�+zˣ�}'�d�����5��e7��ؤ%�����3W�{����L^X�d���O�`�̼��\+�T�*{bAw��2Z��]J��L��dӢ�C�t�4��݉�6Vm�4!�S`=j���b�������v�[�z��(U���Ag�l���or$)@GW+��+�I�M��G6�qMJu(vkZ��`�����<�@� [zմ���%iN���X�[����P�<�������E��-3C�I9��y+c�	*w8��}��Gl���;����5�e|�Ͷ��7�#V�
v18a�����|,L�;0M��j�bt#��6������GR{s��ׅS8�â�Zp�2�Y����i �{�WsQX�;��`o���|�S{ض�46��U�d͂�5�8D��]�z�O��.wo��}�`ݚ>���A����q����ZIC��%�-˭|[R*�W����lv v+"��{������I(�F�����no�r�=0��?B�;v_�.��>+��C09�b��HJ�7]]F?O;Y:��b��4��z{n�쵱[		������ֆ2��ʡʾ�U�ѧ�0+V�Aok��\=��˻����5�,���N*^2j������[�øv���I�; ��i��EcT���@�Q�^�t���;��]����{�le�H巪��I]���y'oVܬ?PTBa���y�N�8n8���gX�+j*�nw��`9}���J��]��&�Ԃ:�D���U�}5�g��gv:뗯rV���f��JnWk�Ҕ��G��	^�y��}'��C������؜1=��q��5ۗMV���5b�t�D!*���r],Aܺ��z��6�2���f�ZS��Y'4��K~��6�p�BQ���8Q���SjS���e�Y,o�l����GZE������+�H+���<��v��Q�쀽c����"���a����l�$��8榐�������@Te�uiGD5�'L��}q+%v��՛ˑx�j�	��lX�n�)jUFoz9dJ۸�h�58�6��Ov��[��gmM
���g�Ӥ��F�{��=��|�ã��z�۸��e�958����>��މX)��ޯi�HY��M�S�*���_s�7����/������Wd��8�:Q[HW��&����/Yhj\;�S�ݽ�x7R��#�2pw[p�Z��uey8�]������m#i��Fj��0��=�^��&\t��C�EU�����:��b�&�u��}p�)��\�[�w �J��`�<�١!C�A�sosu�Ս�G)�(�b�-�K�M��ܴ�.^^'�̯�򸬭��P�F�QaQj_��>TwBV7�����33V�9�+���w���i����nj�R�c߬�zZ�)�j<�1�����'���=XבgϰmŹ���$}t���P��Z��K�j����$."�
�uv?�\5��2{7�~��_3�@�YWt������9M��nr
D� .+�Œ�g8k�5��ei��ɯ���_$�7�"��+Z��Ƃ�B��٫�t��\���׍ΰ�Dܣ!&6���w#/w���Ϫ؉��n8&�P㩞.�Y/yv�}���Ӛ�M����Y�Xo�ȓ[�q�p
꾴_)Ջ��I��ٗ6$4�F�b��o��n�3^{�x=�&ڰ:4�����3�;����n8�/
D�q����k�[ 2
��	ܛG���^�Q^aB�L����J��=�n��-3c��m��l�/�0
A�Hg�c�+���[�K��0!�N@�y���ږ�X�N*=�.J�mH$إ�s"�{/M��m�D�7�V�0���-�)�3+��N�����w��#5��1��o����v����E�\�w���8b�Ԫ��ֈ^S��rT�8n�c;�	nPvkLF�P|�C��4��魘T:�w)��c��Xt�Z܎����o� ��[b�j�8Z�����K�
I��Z�֫M��%>Y��*��S-ٛi&aWh�Oxp5��|款Q�4_n�)um�Z��������K���+q^-bU�8��&Ӽ	c�^���&J%�`��Jmѻ�+���p�iX�
iٕΘZ�4u�\��G(�^�"�c�JeX*�l�t�,-䘲�-)�$�7ZGL�]��y]:��S01���/Q4�t�;+{kmk�Y�r�*�}yי�~�q��o�h�\1�U�F޹��i]e���6�.�*�7CԹVQ��b�j��
h��w�fؼ��jm{5`��f�`秹0��ȣbZ�t�dC{�i�d������rH��ꪔ�\#a]���#���|�љw����w9@P�c���]�CM�l��T���c�Wn5����Ǐ��a��۳�������#�>���Eeո����+��s��	��pU�n�@�d��q5sZ8���'��-K���Xs5�TV�ܘV��8�Tˮd�;]7-]<y������Y����N�9|�Ƹ$�,T�=�����,^%�ٟD˭*hk's*(�:�]>�qm-ʾ���hYL�ٷњC+�[���`Ws(�MwvPU>'7`U!��n��-e�;��,��5>��=�,ֶ' s7w�側��W��
f>�W;�uq�cJ� S��Z`S�L��N���X���m�ܼgAtJV�5�v�mcy,�Ge
�,�e ��n�R��u��VާOb�MR�s�'�,G�H�y��,#�{��Ցf�ŕ���7@���y��G#��G^mȎc�� (���
����C�b[�G++�;%��`]�����c�u�t�۝5-]I�F��`ܭ54��.��-<Y�YZ+���]���Q].��t�pն ��K]H���[�@jX�g�1�Y�k�V�9SI�1�i}��w`4/V�N]u�����+���x�f�k�W7@�b��J�����Zvi&s��;nL=C%ͺ�x�Nyw�!'!L�)�*�S]ci0�k4\v�85�y{�`�\SNъ�yp��Yg2�$Q,�	�9uH�f۩K"�W�W���.�`���$ʽ�b�5�ܹ�gw��wa�9g;���T:���}[I�ӧnT���Y!8&�z�T���%�������	5���Us��Ոθu��K0u+t�oXVi���n��<�o���҉�;%����gbX�q���
�mG ��F�� ��\�R�\��S"��JrL�!r)���ɬ�3'3�2J\���ɤ2�!2������ ��2K0��h���!�(�L����20��J�I�' L���) (
!
2hr
(J�)Ȣ��\��ɪ�ʰ���(Z�r�0�h��"��2)�̆�S �����$r�,�� �22��B�""̦�
JB�����Ȭ�2ip�jB����"������!���3!���"�
������,�Ȧ�02(\�L�*\�"b��j�33�������%#$�"`�����!b
���������|��9��rJ��j~�'ꗺEX�FQ!vMm��4W.{4�cT�d�&��*�_uY�x���q�)���ro��n��D��W��9�j�$�6�S��U�MG)����q�]O�Gʵ�H��{v��q���F�$�L.p����On��˭��w��?�C7�yQ�\:w</����=����O���yE�^s��q�{�{�4_�;[�y��-��%�=��V>�������z�@<`�Z[�;Sʭ��n����v�Ib��q]a��T��Ǖ�Nʵo��c�c�;�9� x��<�b2��v���r6_,(�ݗ���vj�Z��/�ď���V��7�䢟Ӛ��(��<L�ݏg`�Sk��UXP��/!�|xj*V&恘�Pժ�����7������Q��3���w�m�c�H�ރ�=��Uꡳ���90+��Z-�C2���}i��-�ˣ�Ҍ�7�"�-��pvg���I3Q	8U�t�T��\���}|"xw��87c3��:Yk�[#*e��6提Z�旛��)���a��|I�{ �1Y�
c� ��o^
�����٩�՛
E�0��NN�E1=�sVh8kq#{��Ik=�9��+�TíTݾ:sy��C��b\��X�"���l��G&ЛY`��̓�K�4rmb�8?#A@��o�kT�Z���N���Q�˯q����w�W|���ۇHW�J���TK�K�8"�a8�)��Ⱥ��޷�����!�7�o7�K훈M�[�+�%�i(��	��.�s���e�FE��;��Z4�ca;�GZE�ٖ�%뗟JȥJh�ꈐ]\d%[<B�W����N�cw�
��[X[�ar��͋I9�n9��+b�؛��!��߷�!��{<w� ��C�J��i�H�,)ظ��m��x�p�ˍ�Ǳ&����I��Q�����7Ot��ėݵ��
�s>�����_]Sn�s��L>�6��SF��}�_���Z�υ�o{ÔI8-���\zy�Vq�Oe=\y\������2�.wnʉ������ �����>�g��ӱ��- [���ms�1��.wo�ul��V���o�����]�����i%�����9w���&�>�ʌ˶/)�!��D��O1�3";�`�ȗ����G!l�Y[n�=��.bWYQ'�S㺖ǌ�	��x������&�fǜP�3orN	��p.�Uhȧw�X޻��E(��3d�����Y������Mˤ��=���g`٘��+ܦ4���d������չ2�:�%���N�7���4�S/�:�N[�Ȳ���`��mnNg�U ���5}v	�G�����o_dW2g:N�X�t�W�K�5���7rj�2��Y�֣wi�e��P�*!T���k��U�:��\�t�ٮ\c3�
���~d�P"RspIF�g-?ƌa��E�wp��Ҝo\=cm���?A�\5��s��J1��~����P'�6s�M'9�(��7��銄%^��jrY˧2�փH�\t�]]G����GZE���e��1�VK��pFM
�����_w�LZ��;j�Z9B/f��a)�!6���I�#�v7��Rc(��鳱�8�Gj�-��U���񸸜~�u�-����{�.
c��8�}�K9��@���uҕ��{��+���з��!��<�\��w��θ�V��c�Z����%�ߐ�=���n7�%��aQ�R2�K����솋="=S�R��wϭ�,�֯�
�̮ٙ�		��n[ss&�J%�p���:�H����8m�<�[w��rjqu���7�̌��yL'�ꐭ�k�O㷜S�?.p������r���)5��{��I�!@�*x�_u\�R�*J���N���΢�|���N[�M�m�/�������`ዺ��`������V�M#;��^��Ըw��w���H�"ǻS=�o|�Ph߻�1�j�����M(g>����X�V[�v��m�_��v�N{��{:��[�l,����Œ�v��,�8zyL��/�)5��/Om��Sl�|���s�k����@�����w}�v�3�֗��7�Zg"�}�3��Mɨ*g�(�˱���B��I�'Iwc0��X7Iؿ�O��5���2��J������F��sf�Q�7
�I
���!����;f��:V�˜o\cs�����}C��x��A�O}]w9t��S���p�7�l�?,y؞��|jD�Q�yĺ��1�*�sE8���ڐP�ڂ�����`��u5J��]�k��Z���~j�bva�ߐ�~O*�9�x�:樫p!76���B��NCui��6��	�G�|\�$�����;����M����t����M(y�L'�6#�[�AW����2���OH�_U���aW��I���cU�:�Q�۽�GR�Y��ܽ�-�t;b�Ą���s�6�V���U��m�c�t��ѭ�16̼aƼ�Y\x��6��:���Y�,os�rluf�Y���p�ןBj��NE��DL��{E�k�����=���Y-�Z_�]�:��x�}����oBN�>\���cQ=i��<.
�u�Z�Lծ�Jw�ܾ�Zkj��|{�Z<���>4�yNq��ށ2���n�p��-P�R��T�xI]Ӿ�巓���J��?����Y���E��J|����k����.wl,�V�V�NNJ�T'�	��{�.�w���q��9}$l�XQ�lc��7=�~�P�Wg�4�fO&���o��-`���R#P�l�̲����{j�HL�݃//��V��\�����0����_�T�N�a80�K�4�VU��,ʷ��tZ{���fw9e�Om;x�vXtm2���]�����R��{5��J�D�肧�y%[�f��΂��nn
-���3��s���6��l��p��R�-֔Sh�
��q��������4�}M>�O�=	�{2{+���w[��^���e�1�'�A�박%b�E�ϙ��K��4�	�k�dʜ|ˑ��k��5�e�_;$�t���p�=ƹ��aTV��L�
��H�&�b������G�j��M����q��s4>�5HD'�u�o�ou7�g��5�N��,�~��3&��'4۰2eg&7W:�(�j�oO�s���_l�&�.�P��M%q=!���quՑV�5�@O�Wv��Ʋ:�,[l�ȗ�\+�T��
�7J.>��1;�ͥ�Z�w(j��g� �֋�p��p�rq����:��B�+R��ut�;z��bX闘�ڏ(����T�m����g;x@9\�hR���&痢5��e�>Έ�4oe2�VM�8s��h���}���U�b��]��Ƀj���0�;,��њ�&�aH�_J�\��]/%�𓫂����?
�y}|��(v.��-��_R\�)S��x���LF\z�r-U���v�G����y��t�Sݳk��__ݷ�&�3���w{d��I�k���::�u�1�_ڧl)�o��^�B��Ǵ/�(V���KϛG�{e�JZyr��^�has��P��������Z��Zz�\��7�i��N�����U�a�2��'{���,	t����;��)�ﾰ���5dф�487�͔��v�d+=���X����BĴ�xt���[랷���]:���%�O;Y:���2�Y�c&����]m4JKVZɾp��S=P�=u�D��Tq����WCC�$�&��z�#G8�d)�'s���i�@��-�r���y·$��<˨����h��s��J���5�s���Oь���7��y���>�>����;2R�����%��s}|r�"�2rV��	����6������H��u�=�p��b�F��X�j�Zȅq��kC@��9ԝ��y��8�O�=	!��M��/O�x�M��v$���/q�Z��<8�p�m��_D
ۗc�N���>��>�v�!G�����,���yl�]�I�B^ae��͙���ck�j3h��7����8��N|���9�{��cm�,��̬Yp(�h����p�z�\��F��/�n����E�a�y��r��cW��[s|-gN�j�t�����\������Cf��T�!k/zy�Tc��(vu�}૥CS�-�9j�#W�qq��圧l:3*<�>3�ޝ�6����M�n0ێyC���Y
xEB�]��^��a���y��������j�޿+z���vuZ�)�1z��}���:� �)o*�`U굻GR���Mg>��������g��y��,ª{�8-o;�{�]�V�r��4'���E�s�N9��}�j�P�x57���Qnw�|�'}��n��̚�c_F��&^d�����7f�3��+㨱�+-��B�!�k��So{��Z�0��wV���C�վ�߷:��۞�ӈ�(,��ÚL[y���P�E}�Q�op[�o_k)�%Wg2_����>��mͤ�.�:MIoka�K��Av�+L������M[�w#��Y���s�T�vl�)K5sp���R!ZZIY����FWj�K.��	#}/o�&r)��of����5�T�yC��ъ6��:���{���3���{���9��f�?�p����~g(W��H��(X�Y�	sYa�E7b��9�]���#�9��6�m�tܼ3�g�)�d&H)���SZ��R[Z۶j��:V��9��78vgbjT��&���M����F��N�ߊ���ϸ�P�z�9�K�\Zf3&z�W+tv�D��x�z����.c�L�c���j����@��a(��l��ݨ���YH�[�9�ȗ�o�M�\;b�����W:4�ѣ����Ӿ|�n�-�G�xH�L�i�-ˌfV�|�EOT���9W�ō3VXU��E�i�Ր��E��MXĜ�ێy���v&��򓀷��]����V��%��lm�{����o.�oN����1���OluQ"��AP.{�,m1���K.5!6��0;v+vӧ�IX�nc7�t�GK������5��Z��q�����Ӱ�V#:�|��5�p����v)۶u^ר�N,��g��Y&v2��]��WTL���0������ٝ��]�Zsc���UDN#��������ɬ�ǐU>�\�]V�]Lh�7�{ŚJvm��=�>��u���n�/�j��]c������^lJw��.9��1�~��y��{)��<�zv}j�P������cN$�ab��1V�&R���H)J�:�)6j�XQ��nj���2�alE�*G� Uu��ynz
-����C�ݐ��Fv�S<����㧯+{��r�u�u�
�s��<��8oSO�SO��z=iûC���h���>�1��z�E�*㮍3vJ��[�fZ���'�f�+��P��o���8��.�nQS'B����I��;��Z��7��j�FTM����4�On�G�8�q��ڤ�nU|~f�
J]7����fn��bsD��1�]ۗMֵ�+Y����ۈt��Y~J�� %��f`�u�����<_Gt��Wq[�@e�ֈ8̣faAmj�9D�B������6�3Ί�U���&�7*��w5Vp\���d��mG
נʜ���w`��G9�z�t��eGY[���+��u=��lj��v(�5��8o��>����К9�غ��ϹvNWϪ�e�Y�kw*�+E�W�oBЭT#�7r��9˵ͪ[]1Cn�E�L�O�:cmޖ0'�3�:�ڮ�T��́C�Iwk��\Z8Vmd�m�h_8��W]�;�����_cJ��O�@Tժ����vX	^�z>�fm���5�w�B����*[H�	
;�n+�N���H��OZ�U�M���J#M *܎l�_A�;�����)F��sx	P�_<�pWY���]�P��@�\�
�=v�R|X�%��7����x5#5�|�S���2�Yb
��Ύ�wnA} �)�"�Y�f�{�	�C	V��,R��"�z޴k�+��^h��;ѐn�kp�x�y�l.�PA�EkQ�f�f�S�Y����)	�m6Eo\TȬ�@��H��푒���0I�����`H(�^`��F?/gTC�)��S�;xR�f� d��5^�{�AyX����{�pl��k^�bQ�˾w�EӳyB�sfɺ��ך�±7`0I�f��1��J�զ!��#�<l(N��f�oە�-�Eƣ����ڻ��*Ӣ�����Q�觝�,�5Sצ<����E87���-���ieh�YJRm����Ŝh��^6](�kj��[W�d鐫��;�cv�BWU��xT���qm�yLJ��Bm�n�:��i؍�yَfeY�si�צ�YV���r�[�F�NH��y�q	��z�j��罠9М���7/��ܢ��I� x�wr��oN]�8fA:s]me4M�h>�6�on7�y�D��h���RZ�b�kMޑR��`�7i<4� ;�ٙf�|��Ϛ���5�\Ɛ�RF�U�"x�W��vR�n��(H4��h�eSJF��4��M��y"�v��i�;bmɝ6Hxi'�qjg�N���yvʵ4Rs�����L�7�V>������w��۩MА{;�:V�AKc�YN��	�A��%<���^Zn��*ۻt��z�ԧ3�uһ{|�D�����;*l�V�X�j� &T���a����Rm>-�rV�U�˘��]�ѥM�o��5���6H�Ym�Y]�M�X1�v�n0�M6i�1wj��L��B���������o��I��㬋8�u�wRv�rh�^��9eԳ��t9�����7`8��rd�x�;��x�A�ve�fZ,|۾O3&)��O;�:���kt8u��"�;�3ʭ�_��[�3������خ{V:�t*���X�f����3'jT�-
�V�f�z#�"�:���h����; :w(m�F��|Ŏ�yW�R
vh)�U�j|�[��٭y���}�멉<�"iJi*�*'&����� ���h�2ʇ',�\�
���̤222����H���� ��`���("�����,b�����,����i����30�+!�̘��H���������" 31*�����J�ɠ�K2�
*���2,�2��%��
�������22S,�h��$2�&,Ű%ȩ����0r�(l̩&J�
� � �2ii
H��Ȋ�������� �����"������2�#(��3�l0) ��&��#,ji+,����*��"2�L�B����#)����&����f(H�2(j&�(��"i(��ʒ����i����C�(9[�5!�{�r���2V��M�ʳM�*9����c�ḽN�7dY�Ɓ���C\�?�I��?����3`p+M8%ֶ�Q���^،����cy��}�p�طl)�vi%h�V�9Xk%�kM�Z#%��W��v�Cw�����/>��\+�T�S�Rz����rړ� 7��:�T{buV�6��֋�i��r.qΎ��a���}z��H�X��=_N>�YA��O���-����?`>�ː�mu�a��kR�P�{�=em�s�<��N.��a���v	}?�yB�</��\��M���o�t���k��y\�^�Μ.7W}X���ۮ����d���L�y�Y�U=�K��S��%�����1tz#\ק{s8���B�qF���FNN�:�0��s����q;��oכqq��w2�SM�j//,�P�ʰ��ר�^J�5Z�nl���C�����9z��Q[����K�)]�[��K=eH��u(ED�N�7��4�y��b�F�PY}c�'����2�v�U��Wi��eN�u3R��7�]I�n���Ε��:��f�Yس+*n�v�>Փ�A�Uᙝ��̝�Y�m�{� vpߎh�]��З	.�za�lu܊S��P+��G3��Q���'�f���qH[��X�D���k��s�j'���<}G����o!�u��*�mz����O���I?2j�,����WJ�i��) ��-SzԵ�\>��gmRWMɨ?3*�X�YY����3�W-��W铑+Y��z�ۇHT!)ՌÑ���]��g��鿸&�P⸞?*ic�lK훆���4k+��ښ��E�X3�6���� �Wmڃz�ބ�NY�3�N�w�J�{�O�'���p����\u�ή2���S���Z��TM���eⓆ-�er5ZԷ.Q���YS�/>r�X�o����v��+/o��Ko'1q6�)���mP8�16�}+n���.Lb�¶�MQi*����޸ߥZ^[=|���V�i�}��ë�s���r�����3�4V<T6�}�8�^�Zcr�|sr�ED��`�t-��p���^��8���qw��
��3�d���+�6wu�	��v��JZ�i)zo�f��%!ʘl���;�|ď�=՚a{�}*��Jv��=w��r��=VJ(D�W����R�ru�'d^�����+F��΢�Ъ���\�M����V<�����w��;齃oz�7�n��NoVk-�K�|���`up�Mh���|qV�C�x�������mr����$3�:��,s节�q鬞�<
�Kz^����+(�;j�_��5aM���ղ���{����n�׸*8��U_t��-O!��u|{ݩ��]D���Ǚ'c4ͽ���W2�
����O7��Q�3��쁜nnIS<��W�;��n:�#Ml�C�-Pe�e�SvOO���m��Ҽuf�F)�����-��q��qq$�q�$���l����|�\�R��á[^��^2�&mf���C���g�vJK��kw�8�jd�:i��VA���:�-3ܳ���Zy����q���?%_D�_f�-�˪)g7GG����r��yD)��~ƧP�BX�I׫\b,�r���%��7~M�N����X����c��g.&�u<'+�@�uO}�=��ո�=u�\8vnxX���� cX3T/
!�L�019f�7���wt,�:��1�P9���7����.�]A�4�ר���$B����0̼��n{�A�HJ�Λ�2��j�P�ec3�Z��ϓ��hu�XM�i��V�B�=Q!9�� �2FX�����'F�.��3�^Y=Y�E�)��9��J�t&�*N�땲�>8����@��P�WmWo����-�=0��F/W�h�U�&�n�ŵ�*հܭ�M���&1���A��Z?r�Ҵ���yd-	Nn�
�nY[�(��tj����U�.#T��.7P������<�q���ؗX��.���NH��q-��3��}<������.Y<!��;� +ԧ�n3呾�-Z�Y������#oR������R�Wt���>I�V��j��Va���
�[���}�8��;=�5��x�yX����m���&zW9�t��:�q������L�4���1�Ue �eǣQ(^�.앀!̄��N�)�5��@&�o_<T�Y���2a�Rb�6}".�R�f��gK�z����2m)��f�I\��l�$uN�a��� �Ƀ����i����(9kV�K��ӝȬ�r�����GFnP��{�`�����:K��^��W�F�����h���X��ܧ�ç���%��y�2{ ZQRs��M$���I�.��Z�A�in�u+P��:U��y��h�8ӌ�r��nQ��_%������I��%��ջoN.:���oS�S'"V�ڟt�F7;n��BUA�*����d�"h�����oS�j��q�\g�i&7��}�p�ظ�l)�y�vZJ��1N�
ʞ��ܸ�`�Vm�!=doD$Xm�p�Jr��Ӵ>�5x�c�1�lէ]���NƳ	]h�v���r>���XZ���ӝ:��iv��v�^�%bh��]q/(#��i�d}���F�:��*5�V�Q��-����.q=e��=Q�MDN.��wM�ݳk����rf���X�Szx�u8�W�ɳ��ã��y�ι��.0���N��g��-Ö{i���
��Wt޶�R>��mK|�m�]��x�L�]��>T��싑a��a�o,��op�=�����u�jQ�B�}�'���r�D�^>�(_�z��`U���"�'6�l�:�K&�3\�Y5oL;5��-¤��vw���G�E��U=�K��W=~ͯ�-����d=�􊀦)_Mն[���۷�VV�D�3g\Te�-˭|a��ˉ"��b�yu_;jf�cNwn��W֯�(h�qQ[��������������GVɾ�}{c.Ԟ�*GTm'W�Z���#:��������+���z��/�G)��3�X
g4Q8�uӮ�.�Xw+������7��&�Ʃt>���}����}�/��ɨ*fω<��;z;;x�ah�ݓ����[���E=ƥ��Lc;q�nMA��h)��s�W9�ɶE}�\p|OV�I�:f��y8�?cs���b����S��=�jFjq��˙k���9�o_�Y8���ƨ~�]~մ�8�=b�/v��{���cU������D��_�h��bᤷ��Oכ����u��[$W��*9gb!׽�r�s,9٘#wz$���d�5���)9c@�9��ٸZ�����rC��bOr�zz��8u�:^�����J,�Y�+���Y�E)�Y����	���l՞�X�-sN[���䙗��34MI���ͻq/zn
ȨT�AtIq�+�\G�"	O���s):����).�#�I9nTbr�)T��;Q ���v���u;l(��-�G{_���l\F��?z�ʇ<Ϸȋ�[Y>�H���ч/[�wT��;�x�竪����^8�����V���{�G�W,J.�C�|��gֺ�]X�kح�Om�px�=O�yɍR]@���˞+˽����s/ �A����:
xe�ޥO==u�{�j��ǵa����G{6D��՘�0ӌ������)о�
T5�sA���\�=��8㹐���5*(���~ʹ�V4�m��B�qZ��Rre�"M���vl-q:�q��<�o�9�3��6�ݩ���"a�7b/���� i�����j9��8o14�}M>��F��'׸���:*]j�/䱯�]j�Q�\+�c�,���u�e;X�hu�0i���kE:��vqE���It�7��o��xi�/n�o������]B��Ğǋ��p]�TqԇrML���h++4d�sZ��]j�X�˕���](�b��ى��Y+Z�'jv���~�ߣ���7a]%b�%���\F8{p�];򼸘1X�S=�AF��ܺ�a�
I,_��f!��I�Z�^�ofݜ��K�|���\e}�M�7'�g`L4�zKXP�z���%WB���	rt�$��ĭg�ݗ�c�R>"MDw��K�!z��h{��"��]���J���5pr�67�F}��~���Ι�VxUê ͊���4O7��~�
�����=�{u�t��xdGy����P�~� <6=U�o���<W�C��ě��V�������5���OVMүs���dZT�&�q���e�m���W�O�%�Teu ����|=�ǹ\�oey�@9@/N�#�KD\E���W�ߣ��-]�-�23_�}U��bRp�[�u�%+J|fF{������L~o�r��$*:�ڐ5+���.}:o/ӑ��雭����k�9ݘ��R���WBr���ߩCԵ��8��Mҩ}��Q�OO�_���MW��
&�9ǻ��$��㬚�EL��/u�N{R��R\��Ѽ֥p���a[`)��0���B)�*]n�;}����IՉ�S�Q>A�fmJѨ�������jo���i�J��H��%��@*��[q]u)!v�1v��;�H94�B����I#�>�kY��w~�U{�ʏ���+g�V���S�Àx4z��/��Q����ך+���}�z�@xluW�Wy\�Ra��򹃰��KU�0������l��{M�u��/ڋ����}5Nw;-��6�[��锢{����Nǲ��ׇ ��z�ب���=�x�)$=�Fy�wߑ�'#�[%/�-����gג�^�*5ǯ���o�fL����s��^ܽ�%�Z\���±�v�xd`@b��P<���W�Y��[{�{�Ӽ��R��]y�y�od-��C}�C�O}<�a^����a�b���}��I�ّ^���9����<w�5G/�J�ކ�C����Bt�;�.&�33>4b���J�#!���������{�7�ױ����\�����Hl]���~����`��U�V�1j�����ޡ�<�ʫ�:F"-��q�#� 眎A2�C~��oޮ9�:��޸���<*kgLxF�M�5��پ�SnZ&o�M��D����7��g�����YRs��zc=�,����J��s>�s(�^]�1�f=JW�A��뵘
�$̋kNp�vX��?vq\4gN�[�q'�Iu_b�2�]���WZ�q��4*L��.Z�98őjb@8�e�[�7}�����b�%���$ZjN��}�*�����x�H����
�q�>�vn/���75P�Mv��f�c#r�
�&Լ��`�N?,ʛ���}���{|6��O��xљ/b^GL�]ԍQ���n�x�S&��vU�o�+��������c=[FoK]��S�%yC}��(���$d/u��uԋ�U���dgê�n�[����� U $_N�qč��8&=׈Ϗgdg�z��>��Y��ۀ}�A�(����(���؟��|�����w!�@x��չ�t��5�6�<��u~��;���C�V��L���7Y�V�@��s��Ӡ�꬞��u��.��N��]Nf�ylzuݯo�t{,�-��	�Y�_>�}�r/��5y���~��C"@w`�ʉ!N|sׄlw3��^�+���9	�g�{�lQ�*��vm׬�����E����ꆉ�QD�O��hDbe~�Xώ;�n����m�m����E5���}��1�������H�2�*���X��s!��a|�ޝk����x-��u�5Φ_@Cۧ2Ŀ_�oz��ݿw�<F?;����+"$`
�9 T �O�=��1W�
�fd�ci1�E��.��3S(�v�Vm���"S�����q��ťS7�
J���i@	�K7B+�JXV'���A�V�QwQ�6�T�ԯ�����P�Լ�]�i��'f^����er�#�ip5�����׆�%=E�I�Ț�]"`g�d{n�TtJWd%���r�%jG��$�J�.]�1j]Ԃ�����ǒ�8��\��u⹖���67��圫ʚÑ�PT�Y��%�:f��6dޘ��N�(����M��Օ�����>��pv������ǌ����,��.�@�v��ࢃ�7���b̴v�2����*zs���)�:�BhFiɆTE�8nmdj�Jl6n�����q!X�5��K�F�oh�����|GLW��t��99U'1c;2*$�[�wnV��שB�J@���u}�f�oq�˨Z030����^5W]�����ýQ�]nC}�.����s#�Mf&�SDD��u�ۡ��^ ���o����Yn�N�@�CD�n�w���5ʎe=���v��[n?���wJ�t����\�6+[�,��Ž�bu�'l�,ܛ���S1䅷���-V�7P� )�]Y/z��.8u�o�2�5�R�{`��.g<�}���U�[׽�JT"�F��ҍ��W�`�������"�L�*���ޮC��l�<��
P���x	��j8�M�i��1��4�eZ�ti���W^�\�аpĘ��&V�d�6>��m��T�p��ơ2\'>eS��e>�7h�Y�AK71%�\Cg��Vَ�bj��Ƙ�R��<5����	IQ��V�	�d�a�p�_T�������ڷ'=.�%9�}w�PwҤF�9MӁqB��gd�ت��m:�G�*�.���l�G�7�����o����x���l֨j�G.vA�����7�\����*е!/�\�@fb����7\E�Rn�*Ԩ-(�����|���i���+����*r(ծ4����Q�,��5�dX���{*��K��õ
6�_ݷ��]ML�%���*9�Q���`p�w� օK�v_i�G�wBJo-���ջZ�lFzS0���(R��r�X브"��c(��`�<���Ywi�$�1�
X�U�vi�Ks����ۧ��%�ۜ��Ju��K�ь��б�}��a�Čx�z8E
��]����fjH�'�k*<�c�!�r�%֢�yX��Y�z�+��eJe]�zQ�x޺ˉ��c+�+��J�8�|�&V�����Z�c�9F���!����w�y��Y)��;$rf������T�9r7���9X���G�jm:MKm��]]���Pވ8�SOLH^�T��N��bˉLǝ�w�ޝ���X|CU��h���H$tÔb��V�5p��uZ�/ay\�s��fK�sk8�9N<��)-�Uӣ�^�M-�Di3�kyO�`��|4�T ���"jj�230p�&
��B��(����
��&�X,�32
������r\`����$�&*������jZ��0(�&"`"
*"�J)�"��"��"�b��"��"�&*���d�ɂ
����(j���j�"(�(�("a*�r� �*b�)����i�����*�"�*i�"&�� ��*����2""
�!�����0)(�������l̨�b���"*(�)��ɚ"��&���2��0�"&�h��,����*�(�&&�"�h�''�������X�*���0�*�d�)�"b)� �2b��3�30��"(�ʙ,��$��� �
$���]���� Ot��V��[.�)�ʒwC�|��cx���H�.��sK��@��{'VHV��x���_븪�Iԩ���S����ޥ=r��>�z�\4��7·�#{�>#|�9�a����lS�s��)�mZ�t�b)���q{�F�M�+>)w�f���S�}�D?	��}�����w��Q�Fd��t�>���-ˡ94'>5^Cw�+��/b�:��龜9�(Ϻ��r8F���{�����=�N��B��n�����NLv�e�p�Yʞ�u�ޡ;�+c�s��e#��}
�������[3p��U��TrEJ�Ȁj*7�
�C�;�s��}�=�X�I6���}������n�#��� ��{4]�T�'@'�[`Bj#�F���뜻=ޢ��G]?��׈�kݑ�~y�3�u��{�3�R�2p�mPB$�{�N�c��0}��z�������9u�=~7�_q��"��{�~�"6�_�do�'�{7 �Ez�����(�9�y�H{Àq�`�]E׼:r!c��N|��G�!;�l7��Yw��=�}��Ʒ���^��{0��X��	�������Gj8�f�Ҡ��*��|i�K��f_��c5�R1|;{z�{��oGsy�g@���x2�Rw���;dT���N7��ya\����k^`�2TZ'�ćo'�&�J���uf\��;/��
B���!���n1��j,b��/L��!�'J. �CrК�PRV��#�s��=��$o�h��*�~A������YU��קɥՎ��=���QWק����/*}��^���M�����|����"������H������3USg=�N�\v��v=)ğ��\N�`��	��,���ٛ��6� ����*|�j��]Cܖ�s�U
����u��TQw��O�ӛ�h��~b/�#�bi������7�5�C���eO�E�A4$z�S���$��Y�WuL��ɬK��3�G��o�|8l}Vkj�n_�F��(��C�D/D�-	���Nf�B^���Tۭ�r�����f��gH���i���p�s���G���<F��t[�p�'(!pD��X���4�/�\&��N����}G�����C�L���']<�޺��]��Ty?�r���5˗���*ӗ)�����B�Dx\���o���U��x���O���m�~����tDn��紷��ûT�h�b}���� ga*��Gy���������zw�"]���?$�����U��I�(J�q��٤6�eo�5b�8WX,�r�	ua��3���u�P�OIAY�;��&u��Q�4��ۃ6��)�6K��Y��es����8�%��zQ�#�)%{2�d�b�[�7�ؒ��/y:�}��殮��<L_��Z����:�.v�O��J�׮=�+������G��e�?>{ q$��
�N�x���v�v�{��q�'!�͗:߳ �F璨��ӵ�GQ�3䴪��u^�u�rޜ�>۩�<��MwY~�ᐲ�|v8�Nm ��_�g����++�w�:�x���oz�G��W+֐���x��]���^׏�/��z�GQ��Vn���g@cЍ9��,��C��w��#޸^u��pr;o�ϫhjF�ꧠ+��nd8�i���B��Q��4 ��J&�yd`�,����B[
�рl�w�钳�_�ln��󲦼4 �Ҽr�Ϡ۹��镟O{=#����e?�<9�΋�s�W[*�k[�u�8�f~����;���|���a�9)|�]R��}y/g�~�9�=~���
;��'�����w��n�v
�g�����P�V�]��,ʊf�ܘ���
%:��ɽ"�*Y���35���>9��9��.��A� <*M+���Ug����l��5=�@�]��wU��Y#˥s5�'S7��8>��ͭ+�@�ds��\���1�K�:,S���H;QC�mm����_qS(b��m��:E�Q�²�!o8�;�)"����Gr��y��kA�)N��LHe�vs+��J4=����������w�g�do���wn^DH�(��񫠦Du쮙�m��-��L4g��G��~|n
�d^z������]'}���7U!����Z���-q�~�MBj���g�)xz{��(dC*��lG���=�x�~�G{Pr9܊�w��[�S���u���QA�Sg��!N}�w�T��mg�3�{��],�ԃ���)��{'���2'�m�)����&�Dk�;r�
�&Զ�b}4�͗9�co�R�x�ƽS��������?K[�n�f[�n�JeL�p���o�ء�Qy��]ȩ�r�s�����7����3����<��_��u"�W�W#e��:�v�>�
^�#�Eif	>1>${��	W�={p�'���L��?��p{ݹ9���^�������욻���[~s��U)Y���[ �i�diő�B����� ,�{×�k���"�;�8�ˉ�`�=p��S����E������r4�Vw�ǧ]���GG�ςY�vW���ܩ���u��:]Χ]�m,�$b���s�m:=}\oᘥb̏KT@�kA�2x4�	�nc�+�]"�// X��+�R�Cӭ�`�ygZ��6��[Ւf��x��9|9dQoN6^GaR�ՑA+�k�G8�
l��Mo�;ܑ�oWa�d��=|�jʮ0;�Cۚ�ru�-�ϟMzd��b���x�J�U���]w����נ����L�yjIh���n�f�@�z$��=�c;�o1�4N��W�Ŏ��\W���I�	��Kޣ��s�~�>���6�({���0^�~1��f�>۟L_�I��oH�U��X��+�Dx��w��=�z��ݱ��[�~�.���(T� O��w]-������XmW�f8�?D,��=r��"��ɦ������,v3p�±��5[��C�wwF�Ζ�}�0z	�2=3���LVA�s��
��M/�~�=;�g���>��u�	.�X�0ӼŞ��)���v�<���()\bD�hN���]�Q���إN����.��{q�k�����8�]�w�'����Z,��ɡq	�w�L����b'&.j9�-٬�S�������ݞ�3�O�ӿz�hlO���?z�d�=�W��RȑRؒ�����p��
�|�N:ٯ>���2��8��X��Z�����y��7�S��`QKߋZ+R.����?;}�+/��N�Vuh�P!\-+@����Qs�
�W|��Ҥ+]�ke�.m��s	�h���	]���S�V%�Mk.ֶ�c;RsQ�lK(�x�ڧ�T�&۬�r�]t�܉tc��s�ܷX�gH�\�z�).��6�s����Zvh���?X�K#���$:�J��^�k�̡�F�~����/��d�ڡ�U)�w4�e�L�����#>�:���''ղ�"�p��������f�6�w�3�X��9�0s����_a�xÝ�X<C\N�yd������s�뼟O�;�؝��O�^V�X�G����H�O*�G�䅑׮�oR�&��~b�n�K�$\�˭����� ����������~k7�t�H�{ּ��I#`����N�B�v|*��u�Z(8�Sж�B��a���c<�Ff}������){�7��\w�o~�p��<�¬��������w�[R�dj�{��pBס�{2�<��7��/'�~!:^>ˇ�_��O�ԟ����Q�}\�����D�]6��NU�R��r��FA�sN��佉>�HϷ�>���ߞG���|tz�F�d�Kw��x�d���#E�9��5��Ӟ[%l��ګ�2"ۼ�k���G��s���u���'���s�D�>��p{�
�!�NPAO�
C�1!/UI�K�r����x�Jw��ͽ�{�ZnKSO/�ڋ�bK���:Q�ͻ��y*�]H���<qS�`�ͪ������v1tn���S{Wۛ�k����p<b��T���y�u&j�ź¨��%s�u)n�m��/tL�ڊޱ��8���ӻo�J]ILg:���d�x���9������0��x�):��'(0�b|�C�� a�^�:3�9k��"�.8��/�w+�T��}~@�WO �޺��]��uA��2�X�	;��u�2���퉿ozYQ�� ����(sB��C~�ǀ�=�Ǎ��^̘�g�\:�~s}%��ǲrFTڛ���n��'��'jm]4:x��2;�\��z������|�%�L��˧j�ޛ���a<���:6���U��E:>9�����1�X�g��,F6����N��{"�&�����o��Ig){����_Ζ
��4C=5�t�gN�;�Ɯ�6\���Q�D�;8W�V�^����>�~�c�zrr��E��
�j��!��a��Lu�B�W^8w{�)���ϳsӱ�~#Y�υ��f�#�*O��p�GS��+�>��`���g����sJ��}�&��4z�ᑧzv���U�{����~YF/��S��-K�:u����Oޛ���R�=�z���D��Cc��.������y�M\�W�W�/��%ޚ�?�yuY������K��Gk5��Ԋo��bW��n��}S3vm`�ٰ�e.`%28Z��ڹU�����Z�޹{I��gB�1�y�32���{m����a����i�z5A)2LT�j�K���U���ԋ��d�A!��!�)D�ÎK��s����۪Jt��R߬�����YTuzeGz�!:>G�=��-�����`
�W�����W����q�n�d``5�)���(�8r�������{=��盫:w��Q�����F9��[al_�O���k��ŏ���~.���r���gݘ�>�N1�^o`��s�I򲼦w��q^c��3�_?c�,Fr�� )�py\=#���Kf�{�w�N�����<s"�ȷ�X��o��>tw�s>#|��=���@�{��\ˈ�VH���f���Dz�}$ߤ)�������{"=~Ą���~��s���Ogޫb�Ϛ��sv|����*�Z�K�<�I�bG����CP�I֐�z��c�����taG�ؗ�%e��0~�~�ݑAČ.��_��k ���q�9\|<�<r���9r/W�9#Ќz(�Iԑ������������.M	�813�6�>z: 3^�ѹM��Ϯ�YPK}�Aگ9ފmoo����̩�^w�=��^�>ߥ�t���eHA�zEK"}�L�pݏ���~�2:U�;K*h�]����S�&�J,W�^�n��S\�1��]�gU�ʍ��N6Z�UuηzI����4��q���;:��"2�ML��ӓ>���F�u��X3j�8�m��+M� Z]�ѡc)�?i�j;�n��:�jz��U���W�r׻=/ή��~��V{��=�u���]HC�.�,�y�iW���ߴ��]���j���D/�����~�!|Ϯg֫c�� �ۗ*}�X5��Z+����%���=�U�c�I7���[ �q���ǝ
���7�^��2����T򻏭`�#��K�����+FB�WdU~�\D�t����ӟW��m��gylzuݯo�U��j�dU���\�B��/G�䓱�^��k�V�Cu/<}�<�ͩN�|���evU�+�S陫���J�۞,T�����e���Ԓ&4�����υC�p(�<9��+��U�uBR6�y,�c}�闾��0�'���/z���>[~�>��Em���۩��`.(/������Q`�>�SW�^��n�B�SLg̼�p}^л�>�����~���ed�+�3^S#�8z��uER���@�U��z���.߫��r��"��ɬ���#���z�����L{�(
U�����{�z�d���L�\@�3R�xVM�,�w��z��G�ا�>��&�}�����5���cf��Í�*���i��|;s�;��
��2
�p�@U���],.��KtM4zU�e��W%��j�'Q���s�B	w4�4�Eu�6����"96�0�h�܎XOx�+�Ś9r�*��m:�b�9m7�#.�̄,�D:z��{�?\���dϡ]�"r��L�>�9A�BrR��(�Ȏ~�*N�*1�*Z�*/=�;I-�d������3��ឿ\U��/�&[��WԽf�A�hx�����F٥��9��GjL��n\z�hlO���c���s��`z�t���Bx�.��Z���/�R�X�ݕ���K#�1pq�����R<�/�3އ[3���
�T�2����*߼Q}�`k�
�+-u��N��}K��y�~`�ߒ�F5����<�������z�O��}�<8�{&NO��ή�Qݩ�V�٪�T0�t)=�g���;�M�ddCY�[�a��/�$j��Qk�ݚn뫷/J|�g�7������ �v����g�p��K�	��fx~N$��=�y
w^�	�]~h��z9��z��\�Q׳sp��TKY�w>!���ct�_a,.V����U���gEZ������ږzv߳�+��׃�;�$N�n�r0;�C��+�1�ꊕ>Q�jח.4K��48��=~����^ڝyKޡ��u�hs��A�[������s���s�fE^�/ն�:s.� �k(��]�w"��Ĳ���ιю��^�jK���6@W
��;V;tN����P�$Hi�D��4��X�Q�:#���ȅ��/Y��8	�ō������gU�';���s]u�>ܖ����=B觚,������H�Xi��8jg2#ٶl��_���q�6(9�;����i@��[�Jw�=ۋ6X��h��2Cxݢ.<�7�0��-b={ISUlY�`Z`U�(�q]�8�������n� �h���V�F�9�wۘ{��f'��فe�56VBʙ�9��uy}[��W �m��]�3��݌ǲT�{2�"��or(�9��,�Q�f����f]�ػ�҃��^��e<7����IXx��2U�+U�Y�q�dV����Υ��n��Ep�m#j�t;�Gf�=�F�t��xLț��nU�M�Ax�����'�����NzT���N;��u�T�aLv��IH�|nn>�A�q޺\9��(��t/��b����J�&�V
k:<�N���of:�vKEǸ)��G4�g��v;z��&�0X��]%�QҝBGS��B�r�å�b4�|7�m`$':��Q��c.V@�z�%�:�l���r_c(���uv_8�$��|�3"�+8����Sxf�km�E��:7[�vr"_6�y���셰�V ^;/9(���������@ʴ���XjCό�Z���Ob{G{�v����2��'oz�� f�7 �7W��v2q�)1��Ģ�Y!���:�+#����]��WGj�R�=qhָ���<%u�{Pjğ4�s8;C������.k{�̬)�Qnv�C�����6M��r�o�)�'�i����mY-��͜A��1D2��hhW>���EݹJR�P�um]���`-��*S��X�����J�RG�;+�`P����;�b�"���dq�gxvM^�Ѹ�nW���]KJ��b�Q�q�P��[�wS�R�]�5x�����sB����҂�^'��0qb�Ip�+B�{�ܐV�#�WK��z�{�^�^�ϘcY$�I��2��QoNCw����U�6ݺ�K�JL��4��nZ�]&'ٗ�k���;�f�V�"����A�P�d���,�Sc+ʄ���o�M焀�SMq��5�HV/�:{]5���w�QPν����ں��k�@�:�o=�,<J��nݺo��=���ذܩaӼͰ��8^	:�h���ŵ��^��L�D����*���u�v�+�,��ǗQ8�-V�`�e,y�y҅[4oe:�����2�&|����p�8N�5��X�kidt���@�j��'H:�5�����\5�`O�(2N�����9�7�tm�x/g58k��ɖ�KW�W(c���|�b�Z�;J�Rڈ�m�v'����.�J�AvL��o�:�@
+��SET1dUEVfTPDTAE9EADMT��f$faUbeQM1f`RQ5,�4S1�95LCfSU%@TMAe�de�TQD�YET�UU5AUESTDMAQ,�4�-Y�KA��UF``PQUASFXQTQQe�NT�4�TE1PST�b5TQ%T�TUD��UDERENFQP�T�MS���Df`��E-%$PQFIY&9���Hd�Efe��d�U8ANFMTTRe�Fa�PUQAVYD�cT�ET�`�FFCE&Nf54AT�%�d5QQ4T4%D�CAfe�T�ETA�NS��13Eu8̢��;��V��쮳5���d��j��h���.E"�u�[�N�)�sJݽ�;d��Sq���d��h���(��B�l(�/"{��2����܇���	��b��y�71U��qcȉ�e>�@]Q�\��D���dA�sN��^K�>�Hϣ}s����n��l���UQ��K�Eq��=�
�/��`H=
s5<��9k/�fU0~�n�k�zL�-�E�(g<m{f��^S�>�@�;�t����r�x ��Nf�%� 6�C9q^je�@���<[ţ�웕Z�g�ٿ0�3��d��\�yrndV����!���wY�U3V�����^׷B�C~W���w����~��G��S��5pꃥ32�Y�TZ~ڎvz���-�V�"3�F��+�>�b࡟sB��~�ǀ�=�>����gL�ެ�o�"�ώt=9,������`�����$yқ�Ym'�
~�B��Ck=C���V�+�����Ü��gzJ��L�]US� j�P�*��t|.sq�"ҧ�5��yfX���J���ɯwz���].b��=�bK�Q�����A�nv���k�"�Ν��߈��nH��^���Ep�(ݻ�,�e%�L�f�!���7���"yے����H^3��^�-���I�C:�KLA��ä�h�J�)��w�E����c%iעƐ z,�54�v��`7W;�o4wy:��'�b�*�e�/u@��/��˸եM%۞�S��s��\��=���2�u[�ϳ�P�l��W���'�cl����`�|(uT��27��ۧ؎{�'膳�g4��~N��l3�[�w�d�'�U9���F��1�:�>�7�I����l��]>��5�6������\/:^��ۗ�`�������е�0\���5�NQ�3DU	��ߥRVK��Q&�w�G�ݿ�{+��<�����-�OA��~����z��9Ĩp�����Xr�����s�[��L���g�bv�=#wxP�i�u�e*���+��s%�)�U�*�Qd�N�H�s|Q ��r�ؓ��|���[B�큻}�*�w�_�׺D�}�=���������#��)F�����\󒖯��ym�B�H��f:��j�W ◯{r`�J���{�^c�;�3���|F�YFVNPAK .'B�W�M	��'ܤ_��-�-g2+�>�x�VC���'ι�w�g�o�	���ȑ�'�@�n^M���G�-w~������~�# �~a��(k�,��_�!,o����x���OS��i�Nye�<�)!���t�����_1�v��-YT	�,�Ԟe��bs-��	���$��"�.[R�<%+�FW�V�J0���'n��l�"�S�F��4{�$Q��]MAؓe�F�ZZgާ�gks"K�B�V�Q��Ֆ��*�m�HB�7�?��?ø�bj�� �~u1Ej���?cb<0�a���*��M��L�����Hj�o�߅MêTІ�$ؚ�ʮr;^��O���ʓ�}7�Q�C��5q{�O��w�9$s���z��=����ۿ:O����%]��
a�K��f�׺'�G��"��wn�l]�������A�T�+������L�C�ٗ뺐�S �H�d`��z����jo<rr�j� 3��vS�7�r<C^���*����d{��=�u�mT�<2��z��è����8������{>�_p���C��Fi��z��g�3�4㽷 �ےo���xg�
�l�}�/��/z�C�ңF�7���Yl�G��Yt+� ��^�K"�"߶�븣iV���׾��~]�U��OWK˭�ӂ����2�;�c�J�<�^�=�*����R�N�H��>_�$�7�E��ۮ��Cۚ�s�xF��s>q�������]Ǯoo�y%�3����S�<~�H��[�:�Ԓ6ћӷ\.XG�P�_�\����Z"c�T����g��T����_�2�u%*����w5.�@?#���i{A�c�8�mn�)ݣ,�έO��Z��J�p
u�n��]Iw�F�Վ��޻S�Д\�K�x��Vo	R�zR�OA*��A;��zwq�}j�5�L�������^;/�����շӑ?�ɷS<�D�fL8�zĭt��=�>U�S��gG�5|�Ę[��?D�e-끫�;�����
Wأ`�SL?�y��$���{�>�����~��YfW�Μ�����b�i7ӗ4=��,x������˶���r�½깮i���GxO�j�^�8�@7�w�o�(��C�@�a��2C
�V)��D�^�Sa�7]���SY��)�ǂ-�bPǸ��=��Ia,(�;ȏA�O���@�]�'(1j�W�$Kf��Ʃy�9(+�ݎ�ϟ{s�sJ]ݾ�3�Y�zw����<�w�+����1A��Be���TR���ݿ�5��Mte{xo��>}�p}��mI���������=��������{"��z�g�*[�f\ �/���}M�/�}�a�c>9^@�W�q��!������R=���C���ݺ,�����CSk��\e��� ́�%��S7�y����cR�FD5������(g���
��d��2QQ�����&�i���1ڑqWL��%�?,��N��������s�r���!o���7>�⮮��=wb��B��0��cr����,n��ؒ#\Lӹ�B�5�֣�h.s�X�N�D0�R���
�s�ɓy/��y���Թv{�`�"�ѫ'f;΅T�$�(mԾǮ�;ա��i���q��	��w,R�bS0�wB]��;��N܉���{G��do;D�� � �v�����yu�8�� �s��ԩy�}�/L3��}���ߎ�Ǐ�W��A�䃟u���/j�'�g���ߘ��R�����t��w�w��i�W�Y,_{d?|�9�����N�;�gxW?Z�{�y$�;Fw�U9���*����q�XQ�v������sօ�B�Z�"h43��f�5��yKޡ���ߡyڕ�l��i����}��F�c0���VT���^�*���Q�xqfX�9N'�l^��Oz�'K�Ǿ��?�_�A<��>�@�������d��j����1��y�JF��? ����^���F}�p�c#8�^�߫�egy��NB;�"�@�3=BA�Nf'�97J��|�n�ϭ�ɨf��DZ~R2V�f]fuyɟs�_����>��{�_�'��< V)�Ԅ�U9�m�Xh3��{���w��Ǣ��5>�~�t�������7֤p�n��D��O�
�=fӥQ�g�hW�%��GW��T�tx\3��Edz��N���?Y���'Lz��0��,��Lϝ���im�����ol!6�U�u��ڇ\�����+��՜io�U�ثӚL�d]5�Y���l�Xpl˖H��V��ͬ�w>[��զ��n�jQQ��NV���[X�0ͼ@���>'��O,����boV�:��
o䳺n�����mZ=��DBj+޳#�����(dG4.}�~��Ǫ��xp񾑏�ΙUj����Y�>yr�׉V{(W�@}��7�|d��Z�Tv����;�|��.6��1�����T��wA!��*�c͌�|��H����Uj����5
�^�Y;N���F�E�O���b}���>>�냷+���T�V���\���?W�O�%�u��`�-��M{D��{��~"���NE{|2��O�'S�q��K��͓)���Dk�Ϫ�=���9�9'�U#�׀Q�����m|�{x?1�uJG�������g4��S��Ϭ~9���Ƀ
���O��->%�M���9Ş��\uU����_	=P}��0]>�!�?���N���z����l/e����ۼ��\�}���n˫*'=��9e�Du	���RVK0o���TG4�B�<�k�~c�]�j�h`���~��7�Ivރ����[Uӟ/P��Nv���+_��n�Χ��R�{���H��뇠�^߻���[!H�e��q�b��Y2p}��s�r0���1t?�9�W�էUh���4 �)bYx�1t�2���d��`˭��P+�6�M��V�k2���͔Z��v;1���]L����ϗqy��E��Ѥ$��s�7TQe�e�Y|�ŝ�Ƙ�}ڪ��b�60;C�!�wض ���J�����'NI����M�D�������~�_�O������(�ZN�n�LF�u����G�#�y��U�yn�ݸ��~���ؕ�gN�z+�v��g��ψ߫(�ϧ( ��w�I�79�	���5^���5в���s"�2��Y�{���O��\ψ��+����>��U}����
��>$�Ke��L�����;�!��7�PמY��bCC��D?	�ފ�>�����5�ф�KxxM��dU���J
❉�ň"����(��sV�lS�6"if��L��{j�[�r����d/{ vz�¦����7�&��E�W8���=���푱����2i	����u����'�{�z}>V<�w�{>�؛�n�0�T/dMt������ٕӫcڣѧHҍy���6��O�}�wrگ ��^�>ؗ��7ٕ"�0Ċ�EE���r\n駲�����z+M��I{r׻=;��F�\ϫ=����:�r��Eډ�M��4��d�Z�3��H�D`��Yj��X�!|�224�d=�?fϪg�i�{n؞�W��Or/�گ��nk�d%�n�H�7OL*����#��eV���M�$��s-���9���b�YK����ɣ�g�Xs���j��95��کa�>��-��qY"�e`�ܒ�"5����̘��zkɎ	��f���/)]m����w�Nݿ�xwUnDr���dOWK����,�@#x���j���_�E�L����ط�߹*��n�՚�+�Cë������y[c���j6�vJ����f�����#\��v�<R=��޼�v�{�ु�����אr����+GK�������K/�+����3>�w�xT�~�Hq��u�$k�3zv�F��x���H�gS�r�q�W)��~Y���\ϞğfL=���NDk��Q��۟-�b�I߫lͣ�S��(疪�b��~�h����б^�9*�c>����e�Cؓ���T�{�;�ʷ��;���F��kԧ�6;�Ɂ�ײO�F �z@��L�D�p���u��u�~���N��T�2Ed�3n����̜mI8X>�����X�ȑ��P&|��Nf�R���l9f�+ޣ4��.�ѹ-��X�fv}���<F����]�'(0�fR�P�A�BHη\�#p�`"'�7���_�{�N9R��ܿWr{��D�{"�g��p�/�&[�� F��A�-z6%F�P�G��^@zM�A�s�6ȶ1v>Im<W7�|iޠ~������WZ�2�����QV��]ܖt%׵ֶ���փ��'kV[�Z7z�f>[R%>w�&�r�(`�3��u���<X�H���{<��[}�;�lv�n�ν���O%?� {�1p^}�mI���σ����|C���r#�슸u^�Tb�lW��&�n_�Z�wD�
�c�)�V��=�*8�6��=�R���~���}3쎡ر������\��Y�^u�t�
��(d�����nZ�66�FC^�kW~����{����:9q�y��s������'[T-T0��NLxd���ç;�M�d5yp�[{��}�V+q��pb�X�ע=��PϷ�����G�V�#�(�t����б� 6���>>ͻo�y$�����3gӿ|���W�>O�G_��.dڧN��R�'�s���������cX�^������l1�+�kJ'��ki��G�zfs����z�'E���$��h���w0;�sM�7k)�X��=^���w���w��|&�`#�O_�f�s^ڗa{�=u����JYF_�K��oB��(�����2g�]5��֮�oe(�9�ʿ�u� �Lv���0t��J0�z򲽜�IW~��lϾұ|�1��0�����? ����c�?/�߿aS�w�q�״��Z�(��g��T��?U�Y�WvΝ�:?Z�ɺ�(h�u�F�I����Õƅݼ�[Y��;"�u�w!���C*��<��6t�� b;�y�����d�l��.c=�K�+[ް��i�:4�r�����]q�ݛ���Q�@�HZ=��6��y;�"�4F����G;���=6J�_�T���=��@i��뗹��TW���=>.=n{{�>�G���y��- �)�Ԅ�U4�ǚ]����}�S��]߷Uz<r�?a�����^���\�9��#��P�ӔS1>X�<ʛzU��5sC3w��#�s������.
��"�=~Z�^א��d�������ۚ��e:�6c�Vߚ�z}c+�L�*�9�7fFMw1pP�G����{����c���Q���_���`�s?�af�!�.�1�К�����|��O!O�#����mg�fOJ��5��^�#��`�ު��[2�:��0j�T/g�U:���OK�lX۫����~L���z��Ä��xJ�x�X����z$�F�`�-���g>������Ιy�=饖��z}�����_��I����s�7�˜��Ug�^��6nz��E��
�j9�G�F^���P�Oh�W�B/�j��e2肳�gM��S��|Ϯ|/��L#a����ڪC��惟��5�w~�6����/<��b���E61p`6������y|�PV$�su^���_"ﱎS9����(�39{+�ŋ��Ͱ~�Z��sC�(S��l�n�9��IcF������TL<����&T̆6���1�#yϻnC�V�R�ge�B7{��/q��t�2��6H�թ��2q�Wͬ�8а���@�� c�Sp^m�dk<����M�U�x��umX��tЉ�>� u(��ή�.�Ju-c s�}uZb���;B�EՍ'6��̐���]��Ǽ#���Wn�I'�;����O1f(u>�X�ڭ�*ɹu����	g��af��d3��ۃR�^(6H��]��_����N=�}x2oO��Z�<Bf�卨�sv�t��jJ����5j�ۨQ::��K��wW����1���@��r�abn��/N�dQpC&�n��+T�U	���x��T���ͺc��b�����Ďu.���&Ď+kIG���ԅ�ME+b� �N��ҋR���c�]�Ҡ���J*PRa*4w1ɾ[��Y��O
��f�VЇ��������@�T;җxQ��׈�Pۛ�n^��+��4�h�gf�+��n.�B�m;�ƕ8�bT��jG��y��86��sĝ�4��fm�/,�c��[ϜŊ�<*�3�����r��:zjnQ�xJT���c
nj#z/���Eu�����έ�)\tm7�ro*J���``JnR��(�����̭4�PV��������\k��8�U�Amc���k\gwE�Iö1Ir��VR̃���ڴ�ۘ����pApε�����e,K;������ -�7�L(�سNR�_9V����7�+�6��X�U�C$�%�e;l��<ֲ�P׫/;��Jۗ�b�b)�h�왧74ٙ1^급#yQx3#��B"��f�rG�e�I,/�S�-�����7�$���Tr`R��&�[�����68۳Zn�&�Β\%ea�2"{���mhT�V;d�S�'�Cz��oUµ.k60��GU�=��ں��C�,L���뼢�;�Lo&��=����p�ξk�1l�Y]�k�0&���7vˠX�A�bq�U�UV{R��5��ek��)E�n���h��ؚ=w�a�6u�1+��OT�M�t�DX=?6���h�\VK�h%���IM�nѕ�(eW�^���&�+�o#�i`Ӽ/O^)�(��<h��B�}s4f�cwu]2$�uf��y3�4k��$_���9�.�۸M;ޕ�.S��WPU�0�-�f��s��j���s�>�
[��J��^B���"�>��]�Z��/N��3u���j�+�b.�t�{;_+�N�ʂ�����j��io+j�SRm�&�WR	��*�j�U��u9|F��n���K9��S��j����A��h� �ZJulmuؾpM��EECL��j��$����
fk,��� �� ��"
���"B��32�L�j���"���%ʚs1*��b(��&d��22(���)��ȢJ	�)���	�hH�����R�Z1\���b
�"I�r
i+,��+
*�
���B�"Z)"��"!)b
j�ii"������(�����f�)���*���������(�K,
i��!�*��ɤ�����$�	����f �
)))���������)��)")JJK1r(���r�*��h*��f��"�)JJ*�����Ȭ�%�"(k2Mp�z6����R�
n̻���Q ��m�#
9�3�h�	���ì��[ø��uI���m1��(�3 }q[�K���a�0h%���� �t��?Ӌ=.����~�-W�{.�}\������^n"�A������n�*
��r˖:�c��eIa"��4luS���Y�wo��*�3�P�u~���a�bI^{~>Y	j�"�Cڮ��9�xc	A�U-��Q~c������m�cD���J]��#���zF�{-��� �w�F����R�Ȣ�˿X�����3�����o��k��,o��w��"{���������߂����5�R�'�'��7|]O��I���UCx=�0�)���vkan�Sȋora�J���{�^c�;�3�?c��VQ����}p��\�Zh��=`�
���:��-0�!�ȯ���Eg��{���S�G{�3�27���w�nھ��'�c&�W�W�`�ꙗ�f�%��!��3y%��E�z����������z�O1���k������	�)��T�/�PW��#~"����b��sV�d3�Y���w��K�<�c���і�},\��!�D�"��3�=AyUʷKòg�kn��ػa^h��Q�3i��TYn7;�j@�sy��h�X[�D�\3�#>v�뢶V���#�6�벥	j�ڰ`i�8���_�Z9�k9ڮ��eҹ3(ڲ8M���s���T��G!s��3�X�*jEVZ1ٚ(��qn_���/��._����Wx�덉�n�!S ��5P��M{�=���=��:�ivQ�=�=�ew�^�W��Dy<�Ͻ�s����
������~̩��]g7���}�����'�Wz��xv�\R����������kݞ����P����d}�g�H󝫛�z"�S6��m5��u!��r{��V�������C�J�s��'���L��V�-���tnVu���f�������8r�[���>�.�9�U�?]��lq���ǌ�@�������I�q,���B.׃>��Vhl~b�g�xuvEW���OWKȺ�8-_�8Yrߪ�4v�p�Vo7�I��|u-�K�^�HG�ς���$�ZD��pϐ`wg¡��אs�ϸ��{�{�KI�\ϵ@�s+���3p�ؼ*u��zG���'���M��)E��8>�z]]�uФϋ�j��]�6ǅ;��8�,g�̷�I�dÎ��J�]/z�D{mϖ���N�m����K���䅌�ERʝ�R����+�d���9Ni���y��O��7��O��{�ʳ��^�)umUX�YG"��`4�������א.�?Ka�S�͑0�[���y�2<y{		��:�������wkz�TkL哞�mp|�ʹ9&]rmd��;&s��G=�\��	;�3��s�u�	�
����<wy�BT4!�$�7ٲHTI�nwՖ��# �§ uNf��ᛪn�)�]xW�W4ӿp��>�t=�ϽG�g�J6�o��G�^�@��d3�+q7!P&|�9��K°�l9�g,������}����dם�zz[�[!��O�o��;=v�<��Ũ)O�N}A�BV���n�����	�F	�V�f��#����J��_�9�Wrz�3�����Es�Be�\m�c'd}�M>��U��==\mX�Y^A�5����pߞ9�W��WO�ȇ�_L���dW�����bnN�PZ&}�T�*t���_S6�+�n�����ڿX^��H���3=�c'x蟼�Y\��%aM������n��� ���U�0*ٸ�o���xu�	S!�mǔ?<���,b��������U怡�q���_fN��Up6����l���v3��߸�"��Q3j ��m�7�F�~�k�7й����z/�27����}��/��
�v������^��[*Y�*�OLY�̟n��>����#Nfϥ:�d&}r�O��$�ٹ��{n�t�7{�U߱���ߓ՚B��̰w��M`yKg׶�бS!��j�4R��aY��������Ί|˭�Pr/v�c�v�[����Cʱ��go�3��\�f�C��زr�zRlop»�s�"znf*�w)	�e��(i5��Q|�Ż+�[&WE%Ž��l��F�Q�H�H:"/�E�d`�}#��q���yg�]߳�)���~w�H�;Fo}�S����d[�LO���\��O�~�|j^��������\׶�~yKޡ�ˎ�^v�F%0�na�g�m��������[AfQ��{��p��̰l8�0��������^>ȏ\����y�u����|V�Ba���'�jO�kht�g� @S��j��9w�6�i�gגΥ�-̍��}�3#���a����c��X^�Di-=���w�>ӟj_��|�fҎ��w���J z���^Mb^�I�>�[���\������X)�Hs*=;�Q���`*��"��f�}T�����(�{L��;~Ν��~aw��<o�H���3����{��:���V�鉼�3/�@؃T�s~W���>������2@ȍ��O^�Y����b�ٺ���~ɤ ��A3�U�t&���#�����(dsB��7�lx#���78��}�|'�q6�q���<�}�pa�(�%��᣾Z�}��L|�)�w���~CE-#�}�|yBٳ���d�!��Ш6w1�>g�U�wc���])��-F��|����
���\t��9���{���ݏ�WQ�KZ����Qr�HUf�R�s�{�!rt�װr�I����r��Cv����j����X�����ꤢ�s��v�R��]F�>����Y2�:��,�����<yOŌ~]����C�y:����'�oO���ħ�wbo�(d?W�O�%�u��`�.`��g"&�����X=�ĥ w�|q߈��~���l�ߛ�e�}�r��z�2}�9'�U#�x#ڟ���Z�Γ���������_��b��I_��:��>�;�������{6Aڹ^9���Ƿª=�^�Q�����T�:�:�F���Y^!��pD?�zu�߻�O�ʳ�¤
�3���3mQ䕥Z�_����j���r�~��)��%���~+����܏y ��y<^�
��)RkAݕ�Sy	o����ڮ���;"*���Q��d��Ǧ'������گ4��$�m�h�9���g�d'k��=t�9ٸ�U�C�N�p������bA]�ęZ�<�MEq*������ؓ��{����'5ǯ���o�o��S�#��Gn�� bkۤ�W�E{t#7�vz;��Ӑ��ڭ[���ܘ{��{:{�=᯽s>/���eU��W�S�!mZ��&ҋ�=.K�ͮN�1Z�����F��ImQ+�� �C�hr}��b�S���tL��9�خY�-�֣b��#�e*�4u��ANt!�)pt�'������ZU�Ǘs�ԢH���!�)�dF�����Ԥ�2i,�N_�+��p��^=p ب�M@J����ߙ̊����Ed;y��>tw������E�n��y��c���h�[<�����ۗ�0*���⃙�n�# �l=�o$��<�/��HW��j��,�����n�8g��G�>��s���Og�ثuR�PW^�5ݙC�s��(�#}%�u}��Od撏v�����xG�l1�<������r׽��#�ra�ޘ�FW�����w�W�/s�)ϳ��ʓ���K�+��؟\lM÷qV��`^�*ڼ����=Q{�}�o/F"=�#զ݌ܯ#W�%~�g��>�y]ܶ��7!��������ʐ���|7:*휑g+�lr���D�	yPV��ey�{�!��5��N���(f�\ϫ>�{=2G�����	��o���gW���}�R,�\H��:�VD_��ge2<�BT��9�S�a��@u"�צK�UQs.��e@�|�nJ�eVt�,m9Y=]/>��O+�@�x��>�W"�c5>�e���w}�}��W��޵���2�YØ��hϑ�um�_���5h��5����������R'&���Db�����'��JSA��@d\�g�x+�����[Z�s^�O�^��s/(Ê�q7�%�LxRpW# g�Jc��7%���XT�����.e��ٰ�����B��l<�}\���d��غd�s�����:�l�YԎ�O��m��gylzw�v�����>b=��'~7�E��n�d ��υC�:Z�?Got�
��k:C'��^���Y,��]4�V�>>x������~1�g	�2�yzZ��$U'\��T����G�H5b,�q��p}w0��=�`�a{���m��߯ا�k}�z���7�i0|����}�R�2>�w�jn�d��͓���t�v������|=׫�N�{s,e��(Ĭ�Cn�q[��Ee�Y�\B�H �S���+���n�=r��"/޼�SYU�q�;�oǽ*�{<����|ީ�9��d3�+y􌐅�>W��D�^�Sa�T{�LeU�����F��fǭDY6��߱ON�}�>��r7���!��\()O�M:C�;�;;5��C6�O�U?*��+9���y۟�Sވ~�@��{"�g޿\U�A��>_g��0�3��e��a�����&�_W�f����C�5�&q�<s��Z�>���޾���jC��kzʭ���ڮϤT�2>��k���Y7��|����z�{�|�7#=c��.��{����I]<V�o:��{�C�y���Z�Q"�C}�&�����>P�+7�8��?��YB���wb�ŮX��V�L�v�s��9�:,�MS+f�!l�G3�v,�z�񖱱F�F6vp�h6���Yd�|���t�{�w_	�e���"�?�/�~/@u����`e/~7����o����^���2��{�О��|{��T�K����{�P~�L���̜�=�AaW�''ղ�.���o�n�ǕQ-��I����ٹS�a��^�����~���{Eh�#�+��k'�����Kx }����}��~ �s�ә���N�v6���3���R���FGw���z��{��n��Hp��K��/l����F�3+;�=;����ּ�y�I#Nњ텾�l��E�.�vʉ�u'�:����	\z���|.��[=nfn5��yKޡ��uw�ǲ�~����͵��v4)�߶�M魡�^� �l@�p����r�O���.;��<���7}�{tz;��Xō�.��O�ԝ5�:s�t 7T��5F^���dw4�ʞ]>l�3>4i �؛G��亂��s������{�°���C1Аn9�� ���j(nD��%E�/\�*�_��{v茋~��Ϛ�zL�����޹�8��<w�Y�"r�
| H�ϛ�ţ���?#}X�#��OP��Xt kn42����:�����ާ<��sFb�j"�>ʱ��Mq�QÇd.;��U�:�A�w�k��a�a��{l��㊒���ص��`�vL�&�Xuњ(-��r��RM6��r���q�8���f;BW:�<y ��1:]T�W���r�^��.߳�~^7�\�9��#��Pׯ����I]��It߇|�ĕb��>t@�T�9��?,��_�������2@}��x!U�f�R��X�[��o��5j�z���:��QMّ�SC��\2#��6';�q݊yK����5��O�n{,=>�nO�����D�B��'�X���M�,���Ѕ? 
����U�e��&ך���>�9��y�>�<����C�uU6�� UB�DJ������;�Ƈ�9��F6o����-u.�����}�,��Co�(g��^�>ؗq�����4C5��)�3շQ�(��7��+:w�Z"�>�~��Ay�.u�f\��K�Q�zd�ޜ����M�U_���Z�f5�>`w��#�]�DZ�ᐲ�G�%��9s�ө���}S�e�w�d^��)�����[�;�Kk�Zʩ�A�L�?q>.�t�����GXY�w������߻�W}U혔�q�}��ԭ�*���׼r�vv�M�[CrzG��TWOO�RXO��ia���ˮߖ93UEm�������KN^;Z,�B�d|^V��|K]DЉ����o:�t���3+��Y�1��>�>��aD��5n�*L�����jn^��rV�Q�0�:¬�%�S����:����ܜ�c�k5v���ؖ�R��I��᥊��R�[����ܯ�ew����B[����Ut���8pr 2��`3�G��V/֦����3}/��@�S.;����xzF�{-�x�	�w�EƝ�ᑁ��
s�ԽR����lpF��P9O��&ꝏB�s��$��^�z�"s\z�=���������#��C3G�.���R=�\+%F����	�:r���V��<��ra�{:v;�^���L��?c���E�k�<���EH��I�NPC��H�>5��+!sȯ���9���l/T��^,����W�GyY6P.e��=�
��ȑ�$&gʺ�����4�l=���(;�K:���<��n����=�U�":��s���OxS���P%=Br��#����)@���3��\n�M�~�=M�A���Zq�>���d�W�O:��`���"M��D�cxp��ι(j�\�hb�>ϻ�*NCk=.v=^X<7��� �'�q��\*rj"F���1G��Ϋ5��g�a�^"+k��5�$y�&׮X%�Cwu)*`5S�9
�f}��+�H*�� *����"�����PW� �"�򂠊�PW��T_�APE�A��*��*� �"��*��APE�
�+��T_肠��TW� T_�*������)���h���9,����������0��ǕU(P�R�U!@QQQR�R����@
�uT!AD�*��J(��P�P%@�2��"(��B���*H�R��R���P)J	�T���p�P����Sf�kSXٔ��1��ࠕ�'��ZD�! ��  ww   ��  gp� ��JUR�p�+c
������S`T�i��0���
E�PR�;��l���� 5���k4Y��d��F�aEB($����4� 4�@���� m�A� [ � AB�'  ](4�*�5@d�@͍ m��*��d `VU�Ep�@�� %@��@c �� ���HR4R�� �̬�Ul�5���KZ6�%�I6�V��C���6
�i�cFZa���%4�h���f(j�BA��9�*��j�L�F&��l,�<��$ T�DL*U(       ��
R�T b  @ �12dф�14�&���@��$ �	�0#M4�M0�T�dyFA�i��d��hf�$i"h)T�4���j20�h2h �q뮷[���ٖX��yV=���´[,��DH������pDH�/Β�0� B:�$��a���R�DH��V�~ߥ>��g����
���QQ#�*,���VDH�6TE��(��0�"Dʑ�ϗl��Oۗ.�7/��B$M])5�i|�r��Ҍ�����q?b�~��C{
�H���s�ɣ?��9C��P�6��x��X1�K	�դwY33�[4n�U0�ї���6�6۬�i�kU�nT@���H���@��Vr���ugf
7��"�����QXHoY�hQ�9����7Y	a9fɆ����ݙ�mhw*L��f�<I\�8V���������W �m��62���@�U�X�.�M!�ä�˯yg�3@���·_|�/�6�-���[�j�7`ܘD�d:��4�u���;.�`�L������ǫs`r��ڣ��N,
���Xq2�8��A�qJ��H��%��woNR��K�o2�3���'�>KvU&㙻OE�v5X����%[�͗n�5�<Z�X.C�h����S�XK9�wj�����"hf e�ndŝI�K�QA�ʬ�5�����&� ���w�*��&�s9�V��%��[r�IiF��0�ٔ+4�]ޭ�9lƬ+��A]Vf�AYr	��uv�Vmi�ьF�؍w������C�t�K7N�ӹy�xK�n�&��E4QJ���]\����M�4�7����g����ִ���K�����tl�;y�-Rì�4����R�-��7�;PY���`Gk�[����E6t�⧘a2֗�1�t�{pZ8N�@��[�ڭY�1K ڭ�K���.�a�b��.�儵���`�v����3���m�:�	vt�8�bn�[Z"$,v�Эhb�e٠Q�\��$����EK[b+'{�X�Q�,Zo���$�66� �(P��L*�~��9cd1��^�j���]X;E$�2��40�����v�@���O:��]Z�B��sG��C��6�:3�m�L�E	�*$B�e�Ӕղ(���F��'���l��U���4Q�I�k���l��Ά5I�ڼ�;�~o�I�;�M�դ����5��;\eZ�/6�Z�T�vb4���������q�Y���1���]�%]C3���˾��,h�`R�@��Eck7�'t�jl9.�5Gd���+�v`�|�-���4V(�c;[mr��m�wm,��(�{�ThS(^�D8�L�Y.�
��HV4�f����S�ya��n�gN����C�����f�T��*��BLNoƊù��E�"�V����w$�.���hJ��i"Yb�e�rf<�2�TZ�"��sU�kv�(mKb�����h�l�[�n�Q�FH�׃7>�kL�V8$`QE�Lm�K;�ʼ�(֤�e_�K�˭a�X�U�,H��H,ƀ�/��
�"������c�A�e�����MR�~��S#�SB[4�U���a.;.��F�--��0L�YuQQ�*U�n�9���v�Z�H�뮞��0v�������A&�8���ܺ�s#ku���l�j�l�-��tYZ��n^-��C�ܳc+���X�VZ4�$f ��p�c���x�H�փL��Y@+�c���������ڔD��ǵ.cAӽv����KJ$(#f�ZªH`�����s��A�p8���jG{w��FXsu���B1�Uj��&�@�&<�U�ʼ��MނN
���1uhe��z��-�-���]o;Wd���^���{UD���a-��ȵ���3~g�
C,rvU�r�ϑ ��L�*�nP�75
���*�V�:���V�+kҮZY,�Fn��-��ۢ/1��U�"��,3����i�78Ϩ]��)rKx�F������2���ܺ��bwg7"R��轿���-�ܺ�]��zް��� M���	ڧO���;h��c
:�L�"�N�h�љ���u��۪zY}L�ԍ+Wh�%�mE�w+[3�ܱ�,DɃخ�V�e�p8��캋TЕ�P$o(�4V�8�Rc�Fm˵mYEf�T0]n4wfG��n����IV�F6��eܓK�bSV���sD1֠��MY�l��7��C:H[���Vj����q����#���c���h��v����Y�
�m��
#TV�����E��&��ۈ�
��1�ʷlҮ���`b�pn=G��h��p��8��ww�7~�DXT9�ı0-Rf�R5�:�F��ٛ��HЁTѱ]�QQ�K�R,l���j�LJ�w{ciZz��C5L�:�ܖn��m<�vdP�c*��SJL���N��!,�gX=���e6M��i��,��9����4.�8�׷�elö�u����VI�RĳW�����R��E+ul9W�IG����f�C����k ���F��*CM[�V�қXf}k4�[��[�ތ�sv������R�Y��ݕ��2�]�Gy��M��Q��M>���ٴY�L��u0������P1��lY:-��aͰ��H�b�a��˛�"b}���*�*�3]�[���Ų�r�m��H����p5^S��1��ʅZԴ�a��E��=��0I{
���hd�I�xA���ˆD�T��(�ɺ^�T��;���nBj!�aabf0[YNٳ�,L�k���V'�B�s:�ކv������<�= [5�1��I]]�5�
��Z]��i�o����e��6S{L���Է)R1�4[y�ړ*�l�� �]�yc��bQ'��W��q^O���he���mʠ6/�o�W�o��+-%Z�W�b`d�U�n�t	�'�x퉚LƑ�(Ǐ^m�6��r˺_"V˒fп�5GV=�K7"ɔ�E=7Z��Fd��S	�znL�R���ke|)W�WwHѬTEmU�Hă]�Wy$�B����8Ϊ51�qIyLR�	�3*�����(QtK�y����pm�R�T�o.%��f��f�<L�`��]�'!ó3*#�Zv�f�ܕE�R	��G^��X�ҫ�	gE2dp^��[�,�¬iYARWYE�e( 8c�܅�P�<B��1ܹc~�pBV��4p֗�^ 4Zg��ј�����F�8B_-.�u��W[�u���{�E:#A�r
��#[���f\�w[�E��u5ua^��֍&2�fj�U�����J�a��Ƈ�nMDo�{�ɆAj]�Gv���q���Ne�!��/i�Oْ�~4f��P��jД��#��Q��,V&�6��bG[3��/_|C��������A�����S�H���7�o���P�v�n�ϡ�&Zgmlq[5�#����.�@\@���ԅI��U՚~�������w��v�б�k��$�ۚ˷��YLGb�f[t�hQ��V��k�^˒��ԗ3`s�6���	��]]1���x�ă�"�U�G��]����4�7��q�he�T=r�-���f��-�*;)�5nnƵ}z������N.,5�$���(OM�%�3M0+C+-oG$��(p�%�k�O�T�n ��NNq�����m:�ps����G�+��2�#WoqB������4/S+���3=uy�8`��\�ň��c�V6���T���ܫ�f閡�x�i 5��@��Gb��4��%}�R��Y2�hX�u�Q�]�{D�p�����D~1R���.��6�W%8k��D�҄�>��I���n<V��� �BQ��������/�y�}��&�#&�X�o��+[���rK�.�:����,\FlpT�7��ɋ[ј7����U��v��:�ٓ�Ff��wN)��eu��G�!�o���g�"���K��!=����U��LO���`�����pS�s �T͚�;{1���f��ϳ�%_6
�y��ܚr�-B��c3�v�1o S�1�݆�	e;,"���$��>@�X�>�r�]c�\f��U��5X<~s�����Xf���+n͆��;�fvv�1A�vu˜$�t��3{1���W%���D��.�%��RӜ7�Y��n������&ɼ�.��	C���]�WP�40l%j*��Fmc�Ǌ�L�OMZ����`ӝo9�rNmuK:$��%�M��u0�^��
�d��T�b���V��ś�]�����|{'H�k�N��w��@F��q̘i�f\\���o�u��/'�3r	�`틞�C��v�
��B�2��\ ���׽r虡������t�j��R,��VbRձYK�=��X)e��(�BK�])lj4��׉h�Em���앢��JdaJ�����*W`��2�̶�wg�M]]��e2��@���j��L���kF��!����u��x���{0+@�Z�#!xۓ�����83�z���X3+':�s~�����*wB���1�̵ٹ�V)([������.�B=t��P�oW���'��}Yo!Z�:#�����La���HAs1����v]��yY\L,���o�q5�����6���DO'+�g�s���QB�g�2��}(��i��R�Q�Z����F��UՋVM����GR�\/5�4�~��J零��<t���LH0�AU�y��n�}�a62=3�������2o+�f���cɗd ��/u;��X�{=r��2�2%
լ�s�c�ӊY��	�386���V;��]���6Yw��]�ˍ�v&��M;���v`��� ��:�̕L�
N�OY��4^V�Ĕߞh�_f�OgOWg+���;�7�\�������&2-gL�v7�h]�ǦS*����}��Z�:���uö7|(�J�x�D<���L��s���n��P+-�嵨��U�wb����R ̳�봫��OFz̃��N�Is���\tcyh+�3Z���J�w],��v�<ҕѸ]ط.e�	��g^ܷq�]$h9c�D/083{:��o ^i���&^��K���hÔ�ͳ׀��a=5B�S�73�/�ӡ���ke5�(�9ӛ]���:�4����R���|(��2o
])5�p�=XD�Y���>WYx�2�KX��sNܝ�2v�C����',�L����X�r�6����\��.�����
���Q7 ��Y���c}��^n�cn�N�����}�]uqW��tNr�m��]Pa�M�Gu��*5���zer��.J����v��M��u�6���^U�i39���RwU`�A:CV�m'#��h��T&އ6.�4���p�4��c��F��쳝LkJ�ft��$���3��h�{�O[����O\N+P���f1��S�+{̈́�$,)
y�)Z�ȃ����t�h�����6�rzi��R}���K%�V<ĩ,(d}d�whi�sWsjV�aF����vlQ�/����9DKBk4cW}W�f����T�-�[��u����굕I�n�CB�+7�s��6��n��D8rm)�W�\�{d��Yp�7����}5at��A��V���j���{V&{x��q�u�Vl�j�KH��1$2e�a���R���ҚE$Bز�,�,uND�;Wg�kV�h��<�v����L��R�w���6c
��U����7�y z��Qؐ�m��J�%iއ��M��4�,Z��K;��z�Rx�N��EY��h�.(8�(,�/�fL����f�Nvd�i�t���x�՚�2��ɏMU�X3�"�u�^d[�]��H�`کFt�'��*��b�ЮH�����!�rf�lB���6�VQ�W� ,8��1E
���@��-	�:�<�Z��e�i�x����y�{w���$y�:c��t��(s���:���`�^���dEo�E͸���B��o!�)5,��(�rz��s(���ɑ�kFw��ź;���mr r�Q)�� +�.V-�!ȑg"��p�Ne�q��c�x�;J^L�N��Ҽ����N-���AR�J3c�I#NI$�I$�I$�I$�K̝2G,�k\r�!W��A�TS �Op��8�����&7��[4��7+3� �s�uIܞ�7V��@�B�['M��k/�շ|�l$�u�3��1��SDL��Xj��c��y�b(Mda[���?�M��5��k3�;4��w׏k��s0�b�����#�I|iK�֖�9f�i�(X�Mc�Ԅ=�76Y%u�o.�
��s�moE{B�r�!A౩b�y@eNN��@5�p���׭U/8k]�(��s3�7w�Ts��ˣ�!����۱cHX��pRδz�)�5�|T{�֯���³�ؕ��+E��jMXw�=cL�D�^$xj���kΛ��G��MXa�Z�3�w�5jէ�?~sM{w^���߆�����/�)�7Պ"I"n�U�D�F�[*��<��"u�U5:��}����ۖ�8e�1��ܬ�̧�0J�Z��ï�KꥻQ�hٹK��̅���)�'h�~
��&6� ^�W_q����[wFF��;�u��C\��tq:����Y(r�Ȑ�b;�O�ed.[�(nM�ǁ� 5w.�ZкߞZ�Z!��̫W
��o��՛�ຓ����os��.�ڒ, -���JV�"�S4yv����W�Ի�{us����5H���f�NQ�u���������r[�.�I6����(õ��Bxi�rOu;<�V���n�9Zb��H8�0@��UrZ�bS�6�;�\�t���xr+ԋ����W*�T=2�0�q;�$b\����V�{]����-A��S+w�=
�;�wV�j����\;١4�]M�fV�Z�7UV�#��کYՄ�,aݒ��t1`���[���FwU�x�HMB�򨶐0�1��krţ��F����^s)��-��d�ﳦ���"JJ�R�/���/¡��=��m���ܸB���l��٠�0�3Ռy�3��}b��k-1��¸���`-	
�Mlη,w+Agv��1$ �R�32�̰g�N[�0m(��Skk@��x�@n��N4J�[���#��j�)lt�EwZ)u5E\ę��Ԇ���1_�.��dv3Z�JS�tM/�Z4�dV��y�����Y�8ܖ�����H���fj�����j�{���\WrK��o�-�z��Y��Yw/)jT)d���r�1[;1�"���_%��`k.�T�J�@:�P�EtJ�sI���)�@s�쥲9�@�a���NI���3qk�p�#Џ��uU�? eS�<��I8�Q;��mLb͞���i���1;�I��[�nF�[/>͇[�!�]ep�D���p$��K$�C���7n�<���k]��]$^�:e]h�ߦ#�v�$�Cn�̼�Q�d^u�׉H��oi(n4+ѣ�#V�y��+;�r��˅K�9|�XV�t�Qj�f�dQ�l��̛�99J�m��@P��:�^ ¨-�κ�ee�j슃Q�T̊-����fj�]�h�Ѻ�K7�v�i/�G�1�wK������ǣ�W�g1�©P��6@�Q֝�ˤ�����W&��ca���#mZ��}nh#�$����9���ْ���퍱�.�P^Aj��_��"����je`�X� wq����z��y}h�Op����Fv<7����B��kX]���r��;c�<]�cu�ͱW�
'������Z����њ_56�e�����$���]�p�;ͻ�FԺ&���`�e�4�G�u4�=/F`�5R�p��t�-7��.�^LP.zst�\3fe���U�Ħ2��uݯ��γ�m��ǟ1�͞Xi��n^�Uظ^�"��7�_MUi���૖�}�(l��uጕ2�T�fpw�=z�u`Fu��[�`Q:�v�Q�74W"2�ؠ���y�f[�����E��V�U
m�Q�}`�-mL����6u�r[����Yg��bo�,��}x��Rq �ٙq#�Ka��$�w��˝ݘ8�:���F�s)�FWJ�툋A\lG{��]�K7lJʒ�jr'Z��z���W$�QրrD���b\վ�ѹ����b��4��s��g��t�+2��舽2�]��{-�AX��!qj]hɏ0v%gۅ3�U�`�Ύ��\E���!�UWΖ�ě�;�]�-�6��kP����붦��n\�Vp�hu��<ފ%Ga�η�gi��2��4ޮ{�&u=����F�B�O���\��R��%�r1Wu�ۺוd�9�^�N����J2�b\C<#�V�dL:�1�KC�1w9{Aa��rr�㹚jSc�w"�C�7u>�6���-!��c"ӊ�랝Qo�ז'R�}ݴ�u�g	�]ƺ���jA�\�P�4Y{��Pc��u֊�ھ//�"���
�yx��-��16]�cv�fa�Ubw�u�����]�NPv�;`k�Mk�͑3p�ݼ�3e�:24�ͽ�4Κr�Y��F/��f�����A
�"a�WNj�;;��Y�w�w�]Ī���8,f�u��	ڸ�9+:/��@�k��B��yM��X�4�b�ޡM,�u�7�+��;BI��	42�8M'|��_`�:�UCz� �!�UF�qx9#�iҭ���[��$κe �y���]�SI;X�,<�η��VB6`m$Pw�����f��a��1��9��';<�O�:�g,�q]��b��g+�:`�2fw`�gOWc�;NYЛ��ƨ�6$2`���-3�Wp|�Pئ"Ǐ��0,��xWWE�`����P��#7��F�8��C�\���/��m�$ʿ��˗��O�Sa���f⸚γL\�a5�Yh��j����Z��e�,q�>�W�t�������e\��b�q.�u_P��)�d:�C�G��W�N��o` ��B��A8��צ0�S����bPٷ���_m+�A���*��qR�v�
�W�Y����%�9�{�wY� @ͬܶt:�R{��+� k0��^�bM�{�b]�R1T���7f�������������讳�>\����m��8bw��-�uu����ݗ�ͺ�V+j���J�8��Q�
ħ����f�c$�s\m���e
j80�{�L%��|*����o$Y����A��X���{yk�eD���nK˰YF�憜�VQOE%-����9RC�[���=����m�"^c��V|0ڙr� �Q�ol�kRQ��-��ł��]����%�e��Ν	t`��s|ugb��N��|te3�M�����B^�K3�N�3��F��K�:�Qv�͂+s훃,��ב�XE��5��ɓ�F*Cs��̈B��tD����&g��*�+����7��N�P7e�	�Є���8�O�G��������ަ���^�^��6����e#N�k�'(��l�:���)�5�M��6�;7N,�n��{LQ�I�,e��{��%(��v��c6ު,�����UC���=�;aK�7	��o2Mb��Ҩ���u%�ev�M��B$J)U��t)Q]�?��8��?|w�����)��|�9��7
�ąnm�Z˺�z��J��¦u�"����P#1YWr\Z��mvu���tG�  ���v��j>�f@a��2*��S��m�K�K�p'A���٢�h�7f��[�ժ�:#O.V�<5�d�ǚS/�29bD�Y��Ef-�\��J�D,����q�
3G�c��hś����\�W!yn�$��5�e#i[��f�ʧ��E`x�]^Q6�3W®w.d�y��C��x���+e�������k�#���S2�fF�RT˥EZ�xf������	M�ԯ!����ن_-����qҠ��c1��PYj,R����B�bF�M��E��Hb��1dUQB���d�@�UTe��ł�RVT�Ad6�#���,Y""�dY"�J��b�1%aU,b�X,ea4��X��+`�LdY��m�H�U����3�έ�Xa�}�W�*}|��;W����ӓ%�ܰE��f���i�Ag�߫�
�����DhT�e	���rq4�]J �o��j����(��Z����\�w�*�<wZ�!:�Y؎Cƫj��%�5 |���˅Q���@�Y�)������S�t��c�i��wW���=�S��E% >,��0<�@ɳ{l��5l�����+�Uxu�L�������bDS�c[�]���7H�\�N�Y>�qB�����0�κ�\{�s��#�Iq���8�����J�ª��s(�x{4���s��c���>Yu�O�4��$��9�/�7����x����a�X���5����3L��2���S��0:s��S�Э�03�M�2Y�D��Nm�ۋ�^H��c8�r��n�1Qs����M(ك���G��O;Wl'�(�wDއ�Wf7o\�EI@C��S������l1�u�wC������x�a����P�{j����)Yq�򣪎u"�#��/l2���"mM�}m���vn'u"���w��]>�.���E��f�%���S��dO��BN+X{�nŽ�TNG4�Z}X��uP���4�P�N�b{	k���uJg.m�sBHsG.���Y=u��X�JB�0�dRT��C� ,���zM���V����ނ)�!�4�*�ի׸,�F
���u��"w�&��NQ!�����Ģ|z��M�1��|��k�h��hp�`���R���׸��^��=�B�j��{B�{/iZ<nĭ��:�on9J���ab+�7�n$�E��2�;	�Z��qo˫��X�!����?O	R�M�	w�Hc��C7�טؔO�"q�jٰ�l�fͦ.
�I�ڷ�N��0�E�v��E��Gl�Ꮤ��:Ӥ:r�)ew�|�4I�IvnK+xE>�I�s�R[8�m�gV�o1�	s{�GOF��hf��cr3+�ץj!�81�5�̬���~�%̒���ρcD�3�a�u�ٝ���a��e�ڌ�<�t�l�Z-�&m:�!�H��E=q38Zط|��ǬeL�eA�ۨ±"�v��f���#��j�=�>�������S@�<"�������*y�;��[qը'L��:�fr���gkgn6�鰺�p𹃷���y�7�;O��<��H.ƹ��-ƘHU�,�nY2v�^�rҢ�:�P3���Qv����>�.�kp�@"��Ծ
u�{�j�I��̬E̅����1�GU�k����ձ�u�X�NH4�L�չ��)_:�G��Z�.i�Aj`dk�v`��TN>�k�A
վ�T�/��o�;e��aƍ+֞Yբ^jH�`��1	�����]&W��v���ro�g����Պ�b�� �
/x�u��\4r�Wm��.,6[��;��^LvƜ��Y�:"���\FR�$nFv]le���N��H�K��#.�-��&�Z�	k�;�Ȏ����e��~�ދ��>�cıd�����I�x��^�������Ä�Oz�vqT��u���6�H�* �2C�7��N�c�O;4�$={Ι�s���u�"wkD�Qc<Ts�7ـ��M0t�E��u�D^�a��_5�93����dw=5eѵ�qb��Ў���<���mwuU�y��e=n�69�\�O�X}fn��\�!j�)DuS���������zް-����q�Ý�o�o��.�C(:��"� �
��%��ڀ�L��Œd̠�����}^���yf����%���w �ܵt*����'R��W�zrǼ�{�Kg�TW�C=�y
X��b�ڔ�i�g��aM����[j�،�UR��C:��J�a>K�~9ţ��Klƀr�|[5<E�7<㊁	;��5�<&���9S��c���_V�y{���w6��r5�u��!x)���d'x��@���h�H�@s�"ӧfD��絰��PM�Oi����Vh��E���d"V��������,jkV�\���X�����lH��2vѨY2��I�4׹�ٴ�љW2�����S참6Fs�u�q�sk/�bm�l-��9,da~��x�j43l�������f��"�k��n!�����oN$C��ҭ#�2%�２���ٸ�A��*,4��I�UԻ�����2��|��`�z��^wY�)�*��ji�u(�<e�ْM����x�N+�_��Ou�ܶ׎X�!g���3�*8��D`����%�GX�՗�t�R�p��7r���N"�Ut0�g��GJ[4�{q�'�Eb�.i\sbc���?dLfh�ŝ~O!��*����2,��|��SN7�j��<��Ȃ`p�� F/X�߳S�N�a���|�q�[x�x�����Z�@;D�v�^b�����Y�uOv��:ѿt��MՊ�C��5�d5���I��:�D%�!8�;w>~N�mf�{���^�ϲ8�����^���~��a��������}m��%-��l\y���њB�~��]���`R�G!��T�g�ڠHʎ��+U����.�
���.e�c��QAZ6�(:᧗��6�S��\bu���X]=2�<F�m���]F'B� k������`�U�HR��gN�2��}�uAV�F,�6�,��H��h��}�S0X5ao�(S�B9w�;��&�M�zr�*�����;]-�-�v�$d�EfK3u��E1���Y�u/-�0-�]�������� �Nv�V���Z�$詶�9!�8<�k{�,���c�Ek�O�u��]و�Y%�{�����-=�^��`#]�e��9��]|�&t�.�<�J�E�7X�~ﲉ������ש�<ZM�{�@�n��Rڜ���������Wty��4�D�q*�a�H���Cv��J�d,��h+:	���� ��8��h����WU���)(�.�̼�b9Y�����U�<F�q��xDV�gm�l�f����m��Gc��y(Sg&^�grs��n��<bw+�5q�8�[�e��j٧֩fafi�QĪ��E�(VJ�yrQm��OV:��Y���5�����b����ƾ��İaA�ܻ�RP�Xc�u܌)�l3#q'.����"�,;<o�G�Q���+��z��39�>��C]2z���XTuf1Bb
�AB�X�P���!P���(�F�RV@DFJ�@�[�d`�Ʋ)i*LJł�T]2��ք1 QY"��@1T��*Af�1���
��E V����m�P,�!Y6GY���{��|vu�����r2�e*���l$��Sm��r�N��3�4�V�3��d��֟����;�l,k�5�����M\�r��������y�\�.+��7At�<���N8艫a�UTI�\�)��{7oD�`��m{Q%�eC �8�u����M�S����B�!&Grz�S���h<\g53�G/���1�cS�-5��XՅm�0�V�mͻ@壭�����t�W2��pj��O�v���^�#S��D�ٰ��#�,�k
S�[������0�:���m�Z�*��կ�g���ٶ@����������8{�T�2�qw{!��3
�1o�k絽W*�yJz��R�w�5{�r��lR��%3
9�O�ڱH��2ض����#��U�.�9���A�'�1C�1��Mbq<8�k�����LQb1c���K�N�j��{�T�א�eo��C��4�7N��/�mԶxd������W]��hc���XD�-`�z+`m��o#o�j+�xh
�꺎�/���7k�����HMMv����}��A�J�⣁�18���3�\���KSO"CjSX^z��g��O�h�r�{$`̿1E/a��8n�;�z�k $�m�w�6��9����VFD��Oς�:��9�lEa�z�WGa��wk�*4{R��aHl�룞�@2K�.�2�������w�y=O�ݼs(l��a���Y�ݞ����?g�>�?�b�����
�m�|�;{�T�����뻐A̛�!$�}K9"��q�����W[��z�R'.�|0�#f���=#"F��%U�M-�Hq�=��DA�8A6�su�B9Áv�����L^s�;��-��v���M�s�2�����]��Yq^P��Dj{r�5Q;�	�zm��������!���;�}g7޺��d=d>7}H
���O��>a<;��0��'}H?Y����g~s���	wa�Ğ04�����>I� �T��>f$�C�I��s8}�[׽y	��d�3��!��x�:d;d;{�$�!�l���l	��c<d�ߏv�Q�u���ڜ��iS��.��*�ΦjS�S���;�����f�NL���F����Z�2SΚ�q��R�_����d�	�bI����'��C�'Z�ā�ɴ;Bu�@������;�ߞ�s��d턝$�2O^�'�'��H
|����z�������߿s�o�x������!��:@��)�B:�$+&��d�J��l!�q��� o��׺￹�<I�O���x�8æHu��v�$�$�ud�CL鄞0�$����w�~�y��7C���P��j�t��Y� u�C�5� 퐛M���$1��{�~�Ϻ�p+a�L��q�v�wd=d��B��'6���	���La�@�n��u����|}$<g�i��$�0)i'I;Myd�!�����j�^ݰ�`v���}�^�����N�I��!�@� �($�T��!�7�$=`v�Hq���{�\�1������C��q�0� �hx�<C�t�Y6{I=`al'<N�,�1�����Y���<��9��Hl6��i��}`bI�C�<I'l�m��uI;d���|?�����E��l�-g?�I�ڷT�E�ѓ�������ȸ�j�[	�i������M0������u���s�P�$��ud�Ci�7�d�gVb킇���� �'l�;a&�;@>뿎]u�]s�4�{�$8�� |��!֯l��a�Hm�$;H|��$�AI�OP��u͞{ּ������Co�H=P��'�N�C���L���@��x�*m=B0;`,/�z<��>�=��ߠ'l�.�2LI4�����z�
�ON$�,�2j�iXz�K�Eٍ�{｝�Chc$��d�������������<M�8�c
�7�hz�w{��u߹�\��y v����!����I�&���$����d�J�d�<8�{�f��;��ć�d;B}���CS��3�x�{zd!Ƥ�d�@62g��Gy���-׿w����$���$n�v�Y��� t�}S��M}@:a:@8�/]�߻o\�z'�&��IX
��GԐ�`,Rq��Mn�<C'�z�:`z�g,��ě���ڼ����{$>Bi ,	�t���� z��:q���C�� �̏��]3���|�:`�߿P�
Tjz⾽;�ʷH������l&\T��CS/k�����e��Q�Ip�N9����>�I&�Y?x�6��HQ�i���&�t�2Tr�� g�;d5������u����!��ē�1��I���t�Y4�vC���8�o�	�)a�!�>���]o;��}�4�Y�zj��I���!��8�0�8�V��!�ɶ�~�t����xt_u�7�}�'�X)���$��
����O>�1��P���!� x�w���}�^s�$� �Մ�L�	��Hq ��� x�>�x�:����<Hx�w@<dϹ�z�y�s�`���t�|����!��I�>d<Bi�,��!����!ߦ����ϼ�
a=� ����NRC�,�@��!���C�CL=H=�4�!6��<�ts��_w���
bq�<��������w���|8���@�r�<��$6a����͐�+�,n�GS����t���)�Ȝ���5�@�fN`��9ֵ�V��]�$��|��V$�6�3�aα�t`�QM�y$jD�U��}_P,���T/��j�쇊6숂������7��yV�:;/x?�V�t?eП�]�M�g;w�J��1Q��X�N���{K�IzW���P9E�x]�M��i�k���:*�C���.�3�
|�+�r@�):(W �0�*c�C�ΟVi��N�
z���{�F�㏚e��Vi�Wž��Պ�m%���i#a��:�����R���X��)\?[W��{~��AN0��^�/^�Z)a��K��B���_}U��R���g�EW�*~)�t����ygr�^�FI��Rkh�1��zb;S���N��e���9�/h��΁��/�eV'ƛ��B��h]i�w���}�%��IqQ���}F��>R]#�)n�PY/|1f�_U���z�̡�Uq��E������
,�-T�,���+��꿯]aL�@^U��7��]��Bg�`�5\^CF�y��U>�cMUʼ�9U���Z�g�)o����h?n�������4ru+f�ө/f��s���U��#�@?���F|�3r.�̉�h���s��{�C��=�������j�O�Mؘj������Ъ�w��wcq�ns��ݽy�7�v�x�mP�o��p삎�.n�8
n������t5B�G9��@���B6z��q�W�V���\'��k�Л;���;���R��S_#�Ѻl��v����׋]z_�;^f3��\��ҥ~�
ݱ'lVz�Ya��F�z�}{��������{EE9ҭ����ۤJ԰���Z�nu��Gy���v�)�!�z�#;�_-R�94���Q,�OϏi��6�Y�I����ڷʳu��`����Wε'��{5��t�ВT0`������p�6k������h��`c�W�4)}��밡�ϥ8�D��1b+Y��OyU�4��[S�q�{y9R�VD��m�1��p7�>O��ݏ^)u�s-�2����A�!sG[��_Ӵ����_Mw��X�V�r�b�����P��P�]Hin��&��cb9�WP5�غk�-AW���0�/sӕw)����/r��b��kU��,�`m��W��e����S����k�X�K�}#۠O2
1vqY)�ca�nf���a�\wʽF"~U�e���u¯����Θev���z�hu�xB�[���������6G�L�)�z�tf�����f�	c�����Z
���0C[ܤ@�m+�V�����t��բ7;��DA�t�x~���,e�P]a����}u,嫺[2�R����V�D
��Y)ݢ�N�%�g����kx�h=�Gs��;�uZ@^���a�'3e:n�Y;i�1�i�1�'��$X�����2�f6�na�>��a�-�v�*�g�:�t�S1��~��"�_�?'�������Pv��+R�i�!�CV¤r�|����P�
���5�AH���Xm�7j�PY1��i��Yc%m�LDf;t�����Mf�X"�
Ɉ��
$�B��R�6ɶJ��X��H�f�]�"�[Z�M�@�I�� ��H��ID�οk��o�z�q8�kzj���N��b]R�;�Q|C��������BE~��?����әC�s��͛���}�c��mX�O�p��̣/|%�5��-�éV�'nw54;�w��ڱL��|���h�v��쪘ͯ(��V����s�iG}�"�B�~P9�"�M�⌯E�I�T�WK� v�p�\��~5xq�,F��7#�s ����+�EdBl��2`���{((jЯ}�=��\s	+�ZG ��
����3q��N�D�{�����J���b6s5F(�{`�����2{�������J�z��k*����+�U���˖�k ���ݤ#�DpQ����[f;���d�]�|�%
P�mV󝰩D��x;�qyk�buq�+�WLB����		�9/���Xj��.�3���W��[R��������;ɯxx(�i�}���5c)昙}�\7/�v=|���V�&65+���˶�h�U�d�[��ǂ�b��h=��o/,�O��|��]��ַ�֯��yeaۣ�֮x{��<B�g򵳹��	;������R�	�?���{��_���o鯄,�˔L�DwYYĸ>;��Ζv���J�rw��=��R��A�W����Q��n�brr�=-��g[���3�<�.���I���h�8[E�V�b	$reǚ`>���^��'W�ӷ8�}�$���4&�he�x�a����C��؛y�T1�L.أ��k���4yx�o�Cܥ����U��q�vSz��S]��m�qU{�z�U~YmJ�Nn�L�a�b�2��{�K�jX�
�z=����7��EU��=��R�mc,�1��C3&6}{�D��*@<������J`���_{�������FSV/6;!	ѣ�zd5�93��Ǖ�1����p0�W��χ�5���IOf�J��NA4f6%(�[����٠���9
�����C�T�p*0��� ��ӄm�X�2���y?u<%M�pc|� �j��R*d�%�ˀ�s ݫ&�v�+D]{�GW%�H�-�Qc�������2\�q�%�諭��姊R����@k"�ҿ��|c���l����\i�X��N=����ɬ����2���vp�ĥҸ&�&Q�7�%пc�E����ǜ�̠���a����E�r�ɋکkϼ0E�ᕞ�+Ա4q�u���\v��	F7��=E_bQ��c>3�7����q��3e7b��:�s�Ƽ�(�jX�����ZOkX���E��,��GO+f��.woḃ"��	_G����RGz 0g2�O�%}�{�����@Q֨?�*��ț�bh�u%X����q4)��Qrx����&_S=k��g"F�V����b1v��/!����ģ[ga�����E�}�zkTQ���g
�'�핆 ����v�7K��\�l[�O��>Y�8��9��`�8
� ecq6/&�Z�z*:�0�+���9ڧ��\U��	�̖��] ��<�������ֶ�/)j�
��0���SbnӜ���OY��Vt�Ϟ˝�1��W��٫�S���V|<��cq=ń���s��ݾ�f�-c����q� �_#�gp~�X,����OV��a\�I	����KHwzZ
�K��,�r�c.Q�X':q`��\q*�|�f�=ek�s�O,�wqcXG�r��[���P���e���K�<�O%4�� |+��Tʮ'����������J���
��{4/'#o^�	ۺ��U��4���T�
����Cc颯�3=�f�3��%\��+g���~���ֹ�yٕ��O�e�̈�N�I�����)D����l�`�b��ֵ@�1s�޼�7�r-NEϹ��D(ʻݦ]�G��z�rS�H�y>U�;Qy�o.FaOq��O�A�P]� ˚��S�	�5��V��xF�~�8�������X7or�q��<����W���4<�`M�|I>sZ�1�TN�;t��!g"v�:g}���{���р�z������O�Ԯ���K��R��{�7]HH�p���%�?W�UW�	L�c�b~��!���\�ƛO�bi"��~u\��C�xw��l�IX�����0b�e���[*���.��̫��vrHGka��O��R����$�8�ΰ��CdhN���w�c�3�M�WK�-mۼ����{[�G���`a���eߺ������EP�
Vfz}k(�5NU��"S�P��C.���Y��7�-<"�b�V1�u� 87Z���t�a�h8'o'J�EqD����N����}��D����_]o�^��.XY{G5	���/�"�:/�����K����%G�8=���!Ӯ��J~"���p���VP�*��~�nr�������9�O:9��`a��c��F�O.��r�Ox��Y$��}f�{ϼ�i=�Х��yF�c��U|^�[�ـ� �m�yD	�P~�vȳ���M}��/�����Z���3�a��N�A�(ig(>yt4��E��cr�ܾ���@(��Q��-�M����b;tE
2[8o.�r+� t\�_-h��K�nõi@�!	���pw�ҬܳGM�*�\�f^ɗ��m�KL�k��m�ۖ�0v�qV_'Ғ+:\i��cq�{1]�R���/���'�p�Z�UO�,��ի��+���*sQ��}w�+��-�³�X]�\%/�^vNx�K5V�<��oh�!�A[���u�ero����=��4��*ҕԺv,�]T�cDp�؇]�(*��4wIh�Ǖ�қs��b�_:Y��F����m4
S%3hu,�p�(�+g�1x!��"Wن��	��Чā&�iS��A�kyo����	q.f�J�!/�CRn�a�W63m�.��޼���u֒n�_h�;/����A�{D��YUogd�Q�VN<��4���7s�� 4f��R2��f�(��!C5���p1�BY����`u#v�:�T{�s8:jŵ��� JIv�*>�U�z��-2L�b�}̂1N4�pxNܭ�&��+�;̹gR�g�Km_4^X0X9������K6���o�T�pj6{�H����u�`K��+�Υ�!��!a�i�Ӎ�;,T�9�VbR�Ϣv����ٽ����9�Uq����>6(�Ԙ��fR
8�((��;f�2�)���dQ�*E\b�#QaX)YZ�M�
��U*�DBc1U-*UR��Q̸�m��ʒ�e�ea�7�K�f��Ҧ0����jTT�2�bL0�X
VʘɌ�m���Ƞ��dP�b6�m*�*��X�TT*Ks+1��P��:́�VM�R,FBbV��R�IXJ��Y�:}�-~�iK��8�uj���v�X\�z�l��U��|wHJx/�4o1�5ʾ���Y��k-�M��j����h�����7V���/�B���u�ׇx�5�Y>K�Z�N�YJ����+�=�E�K�r;���R}G��!��q�N���{�.��)	X3]eE�
Ꮗ`
��ޗx�rc6ª��=�Yڇ����<J�t~��슷5�㮻3��M����ۥ��]�G�)�����i� ��Gy>��OB�����8���g�m��ȨbUn�7s���1:;���M)$�UU�#�?i���s��͜�;��w.ٞ�����= ��IZ��1k�v�w���
K����޾����v��7��+��D	��إ���1T3Q��T��'���Q8�Ea�c-t�V�c���A� ��(��S�
hN��[�B��o�`k��dIG��-�\g;���oEԀ����oN�UOc�hzТ;$��TU�0���L2�13&���6��㼾�����=;M��e E6�{��E�_un�Ѳ�v7����ԆS�"��ޏ{,��r���'~U�]�:�v�:z��� �����'Mι�ɼ�֒�}�4��"8g8Ф��ةoU�J]ά�v�Sb�QڶFW��R/�/M�f��C7|�Vp����X����\.s�P"�3��������YB	���Tک��qދ�~/�A�+��W�f7j�{w�٧H�}�+psA���c���
��Q̹��,[� �ȱ��^a�wr�@����� q\���5�Z�J�u�Uм5�*;��Fё�����JP��V���eMl�F����Vm�l�˾x��\��bQr�Kx���sni��y�c�NC�p*v�/�F�Į�]��wX�A���6�fuX����_�|E�ʯ�������ݎ�2q��V��(�e���+{T��U�2�ǻC��7���I^�lx�1Ql�NT_"�t��SO-�tA��D�T�9ƏM(��i�j�ڮ�����gWʉ���e>�����g���/!��$9�(�!'Ϭ��b.T4[������ȩ߾��=�MWS���3S�SZ�[�oN˫�8]8����p:�j9#��ڊ���;��(�qщ��B�h!Ť!ӗf���r�#�n1;����:�Gj�0Ӻ���ى��{���ًw��ɫ�KKA�����Q�n6.�.k�{h��bu�x/�b�u�t�0NYA秨{��%8�n�,�U>^�g���l�JW��r��C ZMSB�f1p���,�`C|��f�"B@3{8�`���j�$iD��DFww?M�u�b��c�B�V�̃����S2��Gנ�@�G��'݂��cؕYg.�o����-X�.����aqC��ay`}wB��݊&9�+��Ŭ�5 �]ok�R@����8:�k7u9iu�%��5�6FB�g��2B�m��b�aWZ�=Cy���S��[�jt�p�[����"FcB��Ĥ�/ub����w��һ��3v Bn�^D�����oXەˆ��-R�-�r�4
5�q!̛�8�?UUQ���d�~yX��\K�ģ{LS�^�^�V�+���b�z���QX��ǐ�aN=t^�8)p+BoN��������3rW!���*Z
���lz��W>M)����Hf��<ٳ�Ǐi��v�����sx�$��Y$���8���A��u>c.*T�u�"_��Q��5u���Ag�D'�C��#���|�CKե�@�W���u�t6>��P�ç�Vό�e��{=�-�y�n�xȝ�G�q�!uHw��BY�t��v�Z�`��Y�+�t��yȱ�36�W�54���5�����a䲆�x�8RC�?Z�q><i!��^��v�!!���b�=�h���B<^$V�u[I_U�h�Gǉ;���0����g�U�am̾Y��^X�8rfv�3xW�fv]��5�c�)S0��}V�}�F��"2��}���n$HӸ���c��cK�!�,��ȫ�%�e���▸T���8�Vw
�m�#�ڼ���?^&���Ť]-%��U���S��h����e�eb�R�EE����N�XH;׷�\a������D���Dq�z��[�\8�~<�<�p���<(��������s�1��V��}�>˵!�v���<䗺��)?}���ED:��=�S�AR�\F�0�_Q���6{���q��$��i��ܩ��^�Ukϸ7�s�T*��3�0&-	a��C��i�w%�{��G�<h��ޒGj%0�-h&On�wm]�,8�t�#�Hz֔�?V#����0U��bC6
#��{ֆ1HKW�>0����	{BV�}��k�U-��B��i��k�[J���E�p�C����	�@�1�R���Bqw���:E7�����D2���\��)�x���J��^�����#�Y�)�9�=~b���L׼;oEQ&<4�<�i��W���J�!�ݩ�q�@W-�%'wf��қ���u�)��UR�Sή�Q�]R��؏t\�=#iH��mm��ؘU/j!m^�r�����ƕp7��o��'�;9���j\�$��ڎ���T��	�s�J!����XwQ����-xg�=Y�,�!��Dx�lϼ���@%y/y�}�{��6|՝-!��$��]�Q�����s�:�yM@����h ��GN�H ���Y��W]�G�����3�aE<�THk�N��&ﯨ2*�1���YE���"̓�H��{��(��f�5~s��wT��2��jg>U���5�T��`b���G���J ց+����ȑ��:��6�����,:�+ӂ�flX{� K��8�6�^�YM�'���Z�SE��7[�D=�7�#G]M��I$�&q٠֚�7βr�H��r�-=`����H���Ch��C��\{N����+1�H��c��Edi��R���8�w+�e5N��@Ԏ0pv�R���HY�B�s�wr��3��JD�S��w�D�x�i�1�.X�m d��C+:�.|�bW��/a�Awf4�9�Cq'|Z1�E�46)G�����R�2�b�\����
W8�k��G���ӂ=05��3�1u
]u��y9M'���T�j�w�޺�l&������rY�`w:P�,W��h��͵�|��1�@f�3�u���l]�CA���1�M驽����q����]p��J�dx�-V�[�+[+�!�u���������:�mӵG�7��f��������ܵ��[���Z:SԾ��3^ o^�P����:�]l�X�roht�Y�X�\LT����=�����Ǒ#c��k1˧6F�kB��Ή1��s�2����Q�]K��6�J��+���oD�\�6R@*�C}ܡ���q���=0n�Wz�Ž�>���Ws�Ł���c,�7�]s�2����x\AIY*)U*KmKj֥dQE ,wd+1�����m��[HQ��Ub�XJª*ʅT��d�km[I+��UP�5�YD�ʁU����kej�xH*�uTQH�QKaJ;L�QH����IPE���h�,+*T*��R�XcDQb̶6�uj~�����z��;���>q� V��'�$
mJ�$�E?���ᨷ>�Vw?���2���]\���E!5XF�eM/�{��C＂8p��/gA��.k'H2��g2VwU�a�_{���Ⱦ'��D�R{{OD7*�w_�p�\~i�+
��@|��g#\���x�[����<�cP���S\I�i���w��+�ZC�MP�y"͊�.<~�N���j8/�v�6�KQ^�p�K��r���FC��t\֗:ʪ��ΘQ$m�,�ج�2��.}LM�\�<���h|�p�n�4�O�5Gks6�K�z�����T��j�$9bC���0?yM�\��#QYg+����A��heC&VF������G�9�A���1޵�wn�<�K\��}_!����ە,I�NŜK�"��H������u�������_wS���f��e���`��#ƈ��jEa~�+�^�>w�{%�V�H"�hB5��9q����{/���w�Г���ZR_�|��r�Hcvx&��ə�*�����EC��B<k5��ܴV�l�.:I�Ej�"�<"���W;ޟtOT?W���U���z�\��ֲC���W��L���Z'�i�4�	��^{3{���H�>��$8�2�1���*�*�Ǹ���u娅�l�m+�������^�a�EY�'m{��m��6`�\��Ut{�͎a��p����v����U~�H~ ��"�B�
kMcƍ�-�zN�y�qBSZG��<x\��(�:_�7�*�>dV�w�O+,�X����(����N������e�>�1���h'o5P#����cup�v�j"�"t�<p�ZFD���F�0�(����{w�\P�Đ|����1�&���Mj�:�88���
���$��ϐ�����e�X�o7�|d\YG��A�D���H�D�@a�JA�������C~7s\��3��q�f���s��w���<aDi�Ƒ�AHqÞ��r:��Ǹ�۫�8I�f��s��EU�ʈJ���1�S�эͫ�3���9�)]����{�� ^`w���ٳ�k�1?;�ĩ2bT��*����^�v�N�L��t��!~S�W0Nk�I�e���~͛�qG�x��*����#چ�1�3�v��\_x�Z��C��ħ��)�pW��E�ٻ�����?���mQ ~{G��굁��g����c[.�Kھ����F�-m/��^��p'A�Ij��������;��E¯=m��$�FU0���Hi�-8F���y���3}���I�GhrB�;��3fj�YJ�ݎ��k}�v/��+:ZC<�$b�@��ι��Vg��:�>��v�z���2uݍ�:	����{�� ��	A�x��2�.� 0�s�v��T.�����]��|le`�2�����4���ӯu��;�f���^��FdQ7�������{r�u��#�I�:t�(�3�!fρ�罍�C0�%�����CǏ��|��V=5�i$�0��1�=�yW!D1�꬞�ы���y]�#䰺_Q��g�X���wP:F;��)�sݸ�*#I��&I�J�^ʧ=8��nǜ�|���#�q~�_M_A�Y�8����T�Ü#Ðs�f�t�N���|i
�2�9ίn���=#�6�Ȼ��5�x���'5,� Y��oLP<Wg/P��X��Z�wY�;5|-붰��0T0����k*��
� ;:���k;���n޾��	i%�A<c^ _*�s��C�[��T���aơe�=�<Y��ä
�ƞ�y�́���)|t��ݞh#���W�ی���vv�;��C���j�$X7����d/[��Y��@���0�k9�#H�O��<jV�o?wy}S�Ɩ�ݱ�tߕ��8R�ΩV8�#����1�_y���?X�Q����������/��C�>��,�0yg��G%Uw���^ �&͑g�$,�j�������E�&�NUF��t�2�:��dN3p.�y�@a�����Ȅ��տ/��[�%�}@�j��������(3gCbJ����8���6�t��N��'g-��?PđR���^,�����$�"�}�r�=��3w7H�_-O��o�+�x�4�U��ݷ�:�L��u*>����&aU��<֟��t����^Y�$i��F��2��c�F����u趽3<��dk�&�+�#����Q�6���f׷`��@�n��yD��xf.!;"��n���x���*��4w�g�S�
$��M,�L�k��e�;0�9��7�{EGK	Z�Vrw�I�∧�Y�Ȱ�D9rp��xt߃����0��
8I�,";*a����w5��#(]Y=o$�8"�;�+вԗyЈ[Q�{��&Sھ�Nٵp�����Y���j��D�[�8F˓��H(��|l�ڰ�i��0��HfⲫGt��߳�7K(��5k��>�đ������7EuOoek�hg�"�iPZ��BΔ��æ<�u�����Ȯa���q�0�"�2r�Q׻wK,�||~���:#	"�������Ej�!Ӆ�yO)\�8A��F/��^�����x��k�yP��n$E�~��D�g����!�ŐH��Hs�fRf�~���V�o��D*ok����Ϗ���ă��ry�����gƭa�2�0��n/��dC<�rn�~�H�(���{�M�*9t74�!e��V�}��|�YuZ�ƕ�,p��Cr��ԥ%l��o]�����>�\��ݜBKn&b>�H�쾒�ܩI���p_�7���*�^��I
!�y���P�>准!�<{+�y7o�,����g�X�lTV�B4t�*z���%�nb�`0�_�ngđ�H�@{jK��W]�(��|C�SPIv�f��G9
\��y��fH&���_/!�����(��yx�����Vq����Ay��^^:a��hcX�x�Ut�o�ج����0��k����?.<F��=U�����?q�F�RC�K�'�1i��~�Y�Di�K����~"��>c��z�¹\�����옹��=�}�U�-��	1���޸���i���r̲c�y=��g#;J˱���ޮ��>��/:��bK�~'�F-:~����=(}и�h�1N�BvTµ��?\_x�������h��:����p����5��(ts"Sޙ��HY�Hq�&&E�"��4r��|�.Z"�f�[5�<�K�Px� W-�r��;��*��G����Q���Qi�����&g������*��] ��8Р�{���ͮ�y{��0��E�a�Z�	oQ"��D�n��Y����:z�E��`iӅ%�e@��߷ޤ|C��>'�3�ڂ5� � @X��1�����=;³dõ����"��i���9�D�λ٤)��-�(nf�\ca����XUi�1O)���g�7v�*�r�#�I,[h����Ӈ��Z�eǸ@[����$�\��F���7�3��]�3:�Y���BuK@J�ñuj���m�\���X�75�0Wj�P}�xf ���x�l�k���zd8z冨䮚�
pJN��)Uo����u��n����S�X�XE�M��.L{G�tRgS�7���4�����L� ��w�L��%��+Aq�ZU`u��&"����f�7[��Et����ƭ�vY�0���8���W(k^>�y7M�GSż;��%�2H�r��"��;c�_�yt���!�d��78u����d��+r���㾡�d����Yȸu�RR���9�o1ZAGx&�Y�b4�K�`2�!b�h�-�t�mD�Yߔ�=7�͹$�;��<�@gw	��mf�y���[����U4�P�U,�_I|B��1��2M`�T+.�а�=6�7�/0C��jK(��3XK�\��#v������L��w[�nA(��]���9k��d��/��J�ʐ��q��#���rF���=s4r�KZnv��:�P��	+��߇5v�����[��N�X"t�Khz�,1A"�-���1��-QB�9,�p*E��B�&�#s2ULJ�f8�TQ+P�bTQI��8�s2(*�
��ҁm��KhcˍLLI���K-�T�`����r�)+�\޲cU��Z����c�fҺA5l�1`���][2��+)X�[Gp�4�Mƍ,Yc2�Z,r�M%̸��Y����޹��}u����;��e�q���m�LιJ�������e������|F��c��B����k���J:U�t��/���E�`Ag,>3�^�s����3
4F��ډBՐ�iM���ճ��v��U罯�QĄ�$iæ��_:X{P�A{j__�әs;��I�u-8`���'�~Ȅ��{�]�C��z�귥�<t��hPD�d�eqU�<���xl��	�ƭ��i*���u�}��G�*��4l��r�2S_!*���o=��#iCFD6��3�N1�|sP��C+;��������dU�
Va�>D�bä������!�fl�M����Gi���=����h��c7����.Lj�T�	��	����2?�Z����u��;�ϻ�PVX6p�)Y�y���/v�\��'!�3�ڄ��t�_X5�3#���a�4~�8�Щ�+��ii���F�Z��W^��a��g�l(Q�H��~Yj6caf��=)����a�s+�H��CKA}�0��a!��	����li�.,��W���IՕؾ��Ĉ����"��a����;��n�w0��6.#ևe28��Ƒ�hB�e^���G-����������Ӡ�WOTOAӽu֡������]u�W���)�\�8A�]�n>�=wI+tV]�{z����ܦ��;l߫�L֥����/)�qo"ot͛�"Je��&˕ l'精!)[w{r�V'�zxӘ���S���gID�P1��<�<PZ~�H{��*:�U���<G�^ �o���]�~MQ��%�P����֧:�߅�߶�)m�^da�B���.H�P.�&,&+=���j\���y�}��q�7Pff��s�9��^p�w���]-HC�B�����X��?i����
�����V��Vww�3�v��?��Vx��>l�}�]o�}�m�9F6�|�V�I}����G�߸N��߽�c�������_Sg�"��k�ݗ��V_{�rR��	&+�L2�����nX&BƝ���(s!�r�l#Ҍ[�iuY��bX���E`�ѷ�ͼ��l���������?b'�"���:p�e�1�"�]�S���E�4��S�d�����CǏW]9�{�ݽ���}	(��m"=*;��ىu�����-h]S�f���6@��l�������=�������D�B�"c�Ey��'+�`ey��V�3y �]8h��㶸���ƁK�
j{�ړ���� �"jl�({<�_f�^�	�_d��䡿_�px��Bt��l	ʢ�ن
�����{���뼀aT�����,j�\�@�VG���Z��V��������FbCqag��Vp�lg|�	=1�{�h���L���,���)���PBaŲ�ǭ�Y���pT�^��ć2os!���e�, W��)H#���A��ڳ��ұi���ma'�|��pw@Ȣ�>έ����t��1��H9����Z��������+6�a'�u�7�*}�zu!�=>~Zh-b���GN_��5}�aW�v���,��N|G�C%��M	���	��Wqf�L)���L۰u�a�|p��^��_�f搅�>�>#�V:��dKZSl#���֗h<zv�_��t�W��<Ip��-c�R��X���{\��
O��i~H�!<x�'A~���7���}:x��rz��ZQ��<t�_!�z׫p�����Y�B�N�J�+���m�ѵ��;.��`
�E�����b{��0��4�7�ѝ�BPj՞I%��0`!ʺ��I�zk�מ(�Br���[%L�}W�˺?x�ր�D��f����}�Ѯ����!^XE�8Y���I��GrZ�|��5��v�S6����@�
VG˕$<Zy�M��=v�E&�x����6l��R�C�Y����$�m?��K�z`�5�?� �^/�����ݶx#�����(���qӱi�v&�κ���h��k�8F��
7!,a��B
C���+Nə�O�X�j�b��a�i�������yt��^`��a�,�ƾ���P�D��|I��gu_��/�h�k��܈�5�w���{�OթYAaQ�4'��)F����X�ӝ�^�{�Sl#'���P]��K�$G�k9�0�5��%	u^�{r�\�֑�i�
d?-;�m��ι�{ٻ�B�>���?X�y��N����%���ay#�楧��E�X_=�{�m]������QD*���i�70�HU���A�w0����as�,��]���r�\���H��d�g�l�N���2^�wq�b`*�u{���g���{~r0�>��ֆ�FRz�j�A�a��y��+3���y1\�����8�ܩN��T٬�h�r<��3�E�؅!5z�!��='<=Q�Ȳ�/m���`���c*x�a7 ����.��!}�R1�u��N�}�BIkbx��d�y@��\�ӟ����!����`����Da-�>w�ݮ��ZT��@_�LA�6՟FNl��]:��l� B��8�, �㶃���4D!�����-�a�>$�p�9�����G�,�*�QS��Ab䆱�N��E
��e�FLƆ���$�#yP/�	�9є�{a׶�U�4����ɹ����f@QQ�Q��B�x��nL���=X"C�/�M�#���������^�۽�MD���x�'U|F:~��f�mv���7F��"FUʍ�n���<�Ǌ#?��۪p���㬉�Z	Tf��Q�����&�s�u��Q�\Q��*6�h�3aӃ�uE6V�Q�����߆g������-Z��_^"p�N%�Jv�oL�����vCH�"���c�����<l���+��ě$אO�5q�h��W�~����a�CO�k�h��#qYȸ��.7)�{k����c�(�@t�:M�=�x{����xR�%�_ �N�C������ �^�Εs�=
D�D���a��S	�e�lH�U>���_��{0���F�D�,X|��˶��5�$�?Q:V��vb�����,(�7�|F\�8�Eaf�+7rI{����g��,j�+�E�c5	�KA�*z����!�&�դ#<���͛�9p�3
��v���6�D�,�m]l�[2X�!ܖ:��_}�Ǚy�gM��=3�g�VA�V��-iI	��{���}~��j��M[a�$iç�*Xob�wU��u��YO)�t�./Q<�����S����hxZy�˓��iG+���I�V꒞ev�����Ĵ���kØ��>@�`�Uw}y�O}qфaC�DbW��h�i0�ٙޏ.��>�!��ss}�^s���Y�e�ķ�}lq�g/_0ȫA���>^W熽<���+E>.c�(�-}�H���+,OH�_�ɖ�E�K������b�X�9#��?d+Y�����*z�͕�R�y{:���[b�Ŭ
�9��(�k�,p�n�뒦E�HP�l�k�7����N�u	�l��(������S���՚)��ɷ���k��}��]c��w���p�S����L�rj�;*���	�C"���S�:�AƆ�r�|	oU��&[��4���J��BNX��j�;�R�diR�|5�6+b@H��۷� ^����8�+�5�2q*�i#s����{�XbG.�M�+�N�ǫcVJT+Y�[�\��x��i�:=��а��������^ne���-꺴�L��.Cd��NM���f��m�,�`5��*�۳�W�0Ȯ�])��05�aY�:T�c����`K��{+_T,\W\:l+�5�e��x�Mt��ձF�e���4�.g8��z�{۩��w�t���"���H^��nb�`��f2���_0�5���`�̛��Uw�Y@ڋYY��y\�V�;E��.��$��6`�wQ}��/e�{�Uc�}�� �0�ы���X�Vv����uh����r�N��m��)T2�M���Ll���6�]IN[o���L�B��đ0���b �sE�sE<���.���:T�K܋����D�7'ub�݋)��+q`�94@mnd�Z]���0���Y�S�cҔ��q����G*2���-:r`�7W7�q++DX��n
��B۫�,��ME[���i�˫���b�kijJZ�`��c����cD��A-��(m�R����b���s�e�b���,���-���9r���\֌Q�ܸ�)E�C-��F�V��t��Y��5�RWN��Z�2 �D�B C�7�OwK]�����K�ZS�ΣE����u%��n(}��/ �$��E=c���OHb!��n߷&��-z���G�6G��$Z�喅,��Է}[�=;&|��L��V�{)����bqF�"E@e�Y����yq���u}	>�����ڞ{��/�S%�,��#�C<��Hz���7��*�7�x᤬��C��qe��~Zvc�L��[3{o�xx ��O��L>?2`���A3��W�����I��V+"������ JD��7�7}p��S�71=B|�HT=�/���0��OS��׈��t���q~_q��Őh���J�Q�c�z�OM2���{��)�̖��=T�V�U����;wx�I�H����q�N�3[���Ӈ�G{�Q]�I���A)����8F��~��/P�� R���<k�:�]`q����񬷦��H� :�j�S���gu�g��m@�{�q��9����d�rǳ�_�r�Ў$�HY�?��oU�oMt���6��TY��e���b��H�hJ��`�:*�1jR��}1
��:i!�pά�}~�|�k5_��)�oV��v��r[�U��	 ��A8I�3��g$t��m����!ԫȑ�̝.!�2�0���Q6��խ��Di�{FZ�1{W�?N�:�	�WYc�7�N�ޮ�_$]a�9䳊�^����^�ι�C��*R�r�f�a:dj��m�d�#N>��jC3���T|G����H�֑�^3w�C�����R��wv-��Z����9)����[�{�����1��!��.!�:�t��C2�a���!v�&�D�#5a�\G��h?cYB�nq��c�H�P��)C�/�5�����n]���a�H~����ɑw��o·.��Og�éQ���[l3�M�t�1�O��uW��b�A]�>�,��a�,�=1�}�wݸxRà��Jb� �QĺA�koݹz�h#������ ��?K�g��k��8tl�Nu{U�9M�յ�Yf]�N�l��ó.'��'538���ŏt��\���Y�W�b�Ȅ���{�qT�򾪃c�f����腴,�͂�PK:�S�o��K�x��$+������B������Mzg�����d_i�,�(��a�C��qV�W^�R!��WyF�:t�6Jc�;7��^�V_Oa�dW����F��IV��:W�G����j��x��B/���a�$ix��E�`tT0T����G���+*ǘ��2%ʞ52��z�H��
x���9:a�<�(~��5�V{β�+�پ����E�� 0�G��:�
,�ʺ��Y��}�+D�����dbWɄ�6ZCԳ�=�~ԝ_ӆQk�R����id���b=�vfZ�%"ْř|�u��4xnŮQ���諭��Je�z���!�G�� � �_x�L����wmf���!��Y����-!5g�^�߼�<횗��ٞ\E��b�}�*�b<��:.���p�p��ϊ$��,D߱�?��E�}BXOו�޿E���d�͐����B�1C�N����J�����Ԧ��,4[A6G(ݤBX��J��Z�
Ad����r���<F�A}�'r\�s�":�$!qq}�>YˍD�j��m�Ol���eC䇱�o�#;��$F#5W7W�w�/�#�i�:~�Z����B����t�FŊY' E�2����+���ُo��8U���O���s`b˜�v!�Θ�rC;�L�FS�v����R���~��殺R�o`�`�hY�N��}���^_!>~�A0_����v}AQ�2�8@�b�(��ߘ�U循k�)~���]����O�tޡ�iq+q����ΧQ	J����~c��$q�ZYmF�v__���*�Kp�C�:=�&-o!���=�z޳o3��/�X�Q�Ը�i�LZ�PlG�T��P����5�k^`����9߭ݡ��Ϣ��Fi(�=r��`���RbP$,��������پxV���z�����F�(�W���q���H�m��t�Om$�,V�`�c�1��V|g�m����y���9��Vv.M'�m,[y�TF�]jE��}�kF�;�Ծ(N�mU�YZ�: �8f���앻߾ |r�3�\H���_�� )!qf���H$�9|r_r�L�:�ðy�|x�A�#b�b�w]��w���B�庈#լ�0��2��^\x�&]=��ίk0�4���a�x��6�hA����P{];���l��q������gZ���3���~��ɐq{<ö��|�c�K���a��^�I�A�b��$�A,j��q0���i�����#��x�ㆾ�p�x��o��\;~t}�Sjg�wy�q5���Xl��N��}���ۉ����}��t�7���˘DHB'��c:��fI�_�XAٯV�ԗ�o��;r�uc׼^��5��xc�x)��'*#J.��N;�T���u�L�s*wo~�� ��^t����5~<Y�lx�e�CPx�������x�د->�0��il�<������F�i�KO)x�uoy	jȣ�ug�j`�u|=�����jL�4��7�1��^4���F"x�V�D�գM����'U�.�v��n�i	4�m�,��i�����`�ZlZ�:�WK]��ˢr���9�6��.,��HU\�1�z��8��iT�=T�* 9 �T�c��'��t�	7�;��}o�P�GFlg[�X��rA�Z���y4(��l3��G[
��i�/���d�����a�w��1v�rj��[��;��}�*o��Qv���^���P�5�K�f�XeoN����v�:��lp�6�d)\K��08W�3��\��m�5"�5�����f��3��9u����IƝl��������Xzr��[%||#��Z^�x�ҎH�T�gۘ=Fv�Q��j�JQ��w�HX'Ƭy�$���]���*ddK�
'pnP2tO���ҫv��o�b>OjU�:�c�ь�����t���%6Z2~��� ����f�^vE�zDp�՛�I!�-;.�*�/k�ˡp;m(3�r������ � �e3��
���ywE����a���2���7���gdYC��������mg���8u���b�p	��cL�@4�03$�`aM�6r�޷�҄<�Vw���{&)�1{z�^�*���VYD�<w�]��7�o9������-�ن��Ձ��lQ�쑙uh���3P�i��Xv���n��&��aN��Ej��+{��w�aE<�.�ٺ��
ͼxNS����	'�vq��
�k�74f=p�6�QT?��dp!
ԕ_M�/8��$�<�xs�g��i�8ꩥ�{�;�1�X)�X��t?���X���q�A��"Wu��3`�F��j^��nk��WGآBgJR��b��έ>+JҴ5/�1Ŧl�:"�E���1}pWV�w+�6bma�pk�m�-�g��K8U�Z��6�'fZ�N�d��w��ƺPm4i[��T�6��n���a�mN���Ko�8(q�y'�*�Y�u��&�8��2��A��Ě��A�Le�v�Y�Y��W����w�5D��um�]Y$���rw�'ܱ��ɶ���o���	�w3B�֙�V��6d32�lB��-����v�8�0Z�YSAp|-غ����Sn���T���;;��i���S����`�����T��x��f�5�J�7%+�X㝝Î�J3��Y�Ǯ�۠���`�& *i�&��퍄��[KxJ:%n�Ŭ��B-�ty�'w_9@1�P�!�,s�7���Drq��$nl�W��3���Τv�VG۪�ڪE��\,|�f��D�$y������WM0E��b3�W�-�c�DV�Z�+KR���][���t٤u�*�bܸ��Fն���.�T\�X�-X([D�bb���#mm�+U�DmDm�8�SL�m����J"-kim����mի6�b���y4jت*r���Ef��2ʋR�Y�6ł�"(�aX��m���V�TM��+���*�"�V:˚�X���}�|�r���Y��Z�K1q�N˥��@#�;�%�_�L=�L�Y�Q��8��+ݝUW�)u'�3��Ь�Z��!p.��aQ�>����c�Ge1mf��� �r;y{�0lw�)���8�W<�����=��Ŧ'��w����v�,1s�k�Ǔ��c'�������V�=�]N;�"�iP$��Q��1N�뻢Pl/Ew�m'5Ց���5�5"����s�E��u��ma��T���*~���B.�B�� �ftz;��滕�k�璥�;�՞2"�H�Э콱�)�o"o�j��ʝ�f��wy�k�S���f�K�*��Cb�����:0R�Zn�56��6{g�ү2�p,1o./�w8��Rm
�7`��q4�u�@S�� ��u��$C|���VP��,[�>�bϷ�{�6'L���֡��;�h/9��♗β�)��<�nYN�]_�2�w\�ѻ�oyiwS��΂����TP��s;�rI���	�F�9�iz<b�/�X�^��>�|�V��껙���q��5`Z���n��ZaX�[!̚BHq�Z9�8s���]��$e��n�s59��^1�����D��Y��=Ճ/���2`�B�\�i�q}3��@�������:�e_���ֹM�a�w��MO��Qg!T�~�5��ZT�)��`���� M�⡺ ߮b{�)�aFBvy3uݺ��k�1�v����ܥH����tc�pagh�S���bz��,9����}P�OQ�I.m	cw����U�����C��3�py�OF��K��&����eF�@�ׅf�HIO:l3��rD���F���{����`��K��,e�ך_<��6u�Op�m�*&��Xb�!��YW�w�k���Iַ�]_Yu��[��?���SNu�zo�fF�����:��$�&)��Qb�u���Y����4�NR��#��6��Zձ�c�EjވwN���e�e�ʌ�WK;Ǘ���`Ε���Τ�W�z�t��qiW��[��b��h�Y���b/챰C��@l�r	dǺ��_3Ѹ���Ic��ނ��gw����H ���
���`��wݻ�1=��#8�o��v�{�e�� )���:�*6o��mmp�{y������Lqߩ�{�f��W1�<�0@�f�Y�WS�og�������.ޱ�}�L����}��|�C�f��G*9��7�{�[�u�N�9�K����/B���#Z�	���]�ɐo����E�LI�-G�fCdͳc�"��	$��+ΐ�T�!rr���1Ê���h�i�M����:�odD��-u�R�6���Ԩ����q0+/%d����s���ݨ�-d�]"Z�E�bc��j����x��j�	ud�LӘ�-�!�9�e�^.��y=�����qV�e�3Y�K����V�vuT]�"�Ӌza��J�&�{s5nn@�G�֔p5�c���u8ʘ�e�g�z��Y�}�Z��LWV;�{���.ĖG�p��xj�h�Օ>���*P�MY�j�n��U;#.�𔨛z5�(nw�tV�i$F�M���Y�-�����F��:���Ն�Y� �'��i�ry�m�M�Q1�^��:v�=}\2���יjGg�ͳ�x�Q�b��r��7b&��Vŷٳ#�c�'���UWa�bt*�Q�:��1�̓�r�ɮ=���;�U1M`I5�e��xK���^�h��F
-�|O�j_���/ �۸��b��[!n��KծmWk��ۙ9�Z���m҂k7�;sipFD������G�� $ɝЉ ��u]1�E��D�x�'x��$��{ʝ��V�=�Y�W���w���'W�8�M)1KB�O4�|��dS篽���=FqJ�N=��	���K3ʗ�ǜ�@�8��?>k4���Ѐ�4�% �/}�r�_V_�%�����������)uҰp��Ѫ޵��Pnf��=:&k���:�+0�aWe]#f���.칙��f.�~(P���-�o�,���(f�Iw��7g����04i��ի("WN�wk��d���A�sY0��3x��	�p]O;���a͓63���U���c�J�|�tW:@f���������'�����8b1J��_h���p�t��Y�u:1��^��	{�XpꥫX����5��÷��WHE+ʖ1�Fvu��^ �`�G��A�c�t ��Zx���m�ʘs�͍�*/6hF[��N" c�w�z�r��O���w�\����$} ���y��vᕊ�w=?G�ܒ�\���'K형{��8"���h&6�{ێ�{D��V��}�;�V^��x7y���w���a�Gpݮ(U��n��a�� gI�W���ه��E[��:�5ҷ^�D��>ؔ��%w�����Y�Ԓ�8�Ut漴�<#�x�R�yRe�Tރ\0'(�%Q/�klL��1�xo���s�����z���+��c�PA��8���Ǹ��S�<ʌ6�M�`�)
O;`!��{�}]��$oz����5=�D|��&Йl�cD���+xl�=�}>��/�)��8�ph��R�F�PR��p'B�9���9���
}�x:Qb ���p��X&�"�9o��P���e���q��٠燽�Yt��Il��Ǫ���wƀ5w;��Q�W'xjW���9�qe�l���N�F��yVo��-pY���e\���kT����/�|�E��һ�s0@[`>���/YUq� �F8����N��"Q�=LVω�6�b��w1m>�o�Cҷ@���nR�)2�7[+b[)*{�2+�B࣯
�6j��M6vc���E��m�R�E�6�3ɓ��Qˎ5]��%qޑ�7�x4T�V�tf�yP�~��U7�y���-ΎM��jQ�/-���]��R�h��m�[�t���e�磲��Em�h�N�j���1K��%Mu0*�ם����E�v���d����SK���S:�\9��}h��ZN9�_�a��3�j6��ef�-�Dm�s�k��Y�F�夂����̙�/����j���%�XÃ�����乷K ��Z=�*xQ�Kw��{]ApP�w�/��
�AUY�S��[`�cl�����B�ӈ�X�&-�[j���5�J�B�Z�AVZ��L�uK#ĨT��J*(*�S-� ���E�U:�K�#V*�q��j�
*��DKJ��D�&P���R��KE��l���0Ċ�,UF*�c(��F�
�����mTQb�(�m�(V���f����{�4���1NBu�Ǜ��m���N�Ak��;^��n�ם�o)v9��H/P&�����2�����`X9m���Tr5��N;z�޿O��l3���N�0��䙫�ʲ��p�|6o�JS�����5�jI�n��Qt��+kj�������'.�욌�s��\�yo��r۶s��=68v �uIo6#��qu]�[�߆z���g��;�}
�{;�����7�����Z���]���Ň����`�/+�^z)��S��!�eJ�$R8�A	:����^j��nW�J9���`����,�i�٭����j�A�aNDe.�5�]d0oMs����𭼄�����xE<�_�xa���p�^S��dl���G�4����}��q�B`m���C&��À�>��ֹ�i����-WV�#��tu������9���|Fe���bR���B��amQ��{|�D}�G�~����cx��u~N3u7��;!N���ڙ��1��R�ղ��5��F�OQ�G���d�S��9�����5sq$\ ��ಟ�ѽ]�;+s؆Œ�Y^��ӂ�Aޱ21��FU���d�U���jy��#P5�.VY�r(Iw�&4&s	E"&\��e>#��=#�%��Ka��.���3�1,|v�
��=��a�}iU������y���������c`�]�{��������`�xi{�,t�s[锞^���nݪ}�.�3���=J��f��Y�����`���\�s���nJX�IO��4�9h9Y�h�T�4���K��E�ù���K��"���Y�)y����puz������<9�qUK6Nnw"e^�,����:2	65�r�d�|�8vj7����cP�1��E��ތ�X�ݸe��c8��K�5��������(x)�rTwƃ�+&��q��������^����rL>r"pv��ȺA�lGv����<kf��:Νm�rI0ga��uY��ǳ�e1�}��5ˋyi���kf�_��n����zo*�෡�
��Fnʎ9�J�����㢮��b%�}E=����H���M�zEOa���[2������UvՉ�s�-���;\�wp��Um��4��˭!%a�`O
��N�5��l�C���p��5ܡ��=�A�h3���u�#Ur7>��rѸ�|�<�4�Y��N-��y-�k���ʬ+�Vb
)1��.����T_9l����׳}j��	FRk>��5Su�c.U����}��a|]=m	�X�U�i->�:�C�k��y�[��0�s0�%���~�(:*�֬le3�����w��6���a���B�ʄbZ0�^�s�w���#u�D)ʾ'<��f^]^��t�85\2o�=a��
�뮻�|�.��gT�W��7v{{�k�$L��p���99G80Jh����ps#�:�W��/����2�8͇uណNldrl�r�#���5��HT�1Ҝ��:p2	�)�M�bd��v�cҲZtY��q����q�������R��`$+{�a�I0-A{;,��tk�+���A{��f�{;�cܕ���y9r:K�Z�o��+>b$`�j0��t��-n����Cg�m>�@��M���{T��Ti1p�R`��S�OT��ⷭcD���\J�8e[��W�����!g��u�0�(�'�Ș�j���D�76�˳�����C�|�l;�܄m�|�tS-�Z�+Ϭú�إy�my��n`�4�PS���P8�[`�:����\��,BM�㗛/��r�''-��':�]OWs�#*�=s~u�A��^w7����A�����;�����,��3���!���
]���25;y܋=�\�����>�{0<�:�Z����sk6�����֭��5�2=^s=X�Wg0�«9�k8��o)�)!F�3�zk>"-�j���st��7x5cڦ�j��"����@n��w[�p�!,�8|,���ӛ�[Z������7͗7Z�͌R[K���N�N�Kx�W*�{�M�H}��,��~*��3���$W+��	�|��>�9p��q|Ot���R<�I�M�	%��HS�]WA��u���{��2�̘,6�:�n��{��S����<&y�xmGi��^b0*ds����3K`ζFBp�3MY6Ƿ��^`�y�ˠi���w�>��$�6b��<�d��S�r�I���˒ٱ2����yC���h+�xe%l��o]���ϓ���8��������N���˯9�RyZq���Ǽ�e�[�Eo�/�;��E�a���Kf_\�%��,oU^o�h��ƛ�ф0U��X��Ƹ��)4��>�C�6�lG�@�׈�:=��)c��o�:.=Z���"�]s�41���o�wi��c�}{.�\H�Vx��"�V�.w�����=��d��z��
(~�^j�~��U��V���6i͘�l�{�+r��ؔzFl�;q��g���ޗ}��
�O^���i�}�ag۬TY��s{�r��]z��d�dnH�l�=��Ә�u�;�m�=7*GWWo�xZ_*�E�����wп�Z�,��nL�D��͡;AIP��GR�tS��
��ӻ��v�MR���*n*�G�g/���u�C�J��wk����Ҙ�م����y7V�����ǟ8��6%]��݀ɻ�e��,]Uʀ��#�q9R���F�n�0\+��#-=���#�2���'��őhрon���6���t��H�Y�T߈odr�j)';���v�B]9��z)=̀��苡���V��Ȼ��CP��1L%i%�Up��Rq�-9�1�W:�;ñ�fjU��f�yD��K�KS���ۮais3����˺���r̼�{z4(>̃r����@Zu�	��u��6p��W����0�"�8�=���jw��<E�!|5=�o�XL�k\�et�:��d��M!Ƚ��%qWYRg �`�V��v�Pu,���L�-�����6��)�ܻI��������t7��i�����ȕ�9��I����I2)05#p�*e�Z�|)a��i�c8���]��E�����9�ώ�D�b��U�(��[�
���+\VQ�*'Ir�$�R/-b;J:h,tՀ��V
�����Ӎt8�p�t�.\����w�!�w1w���lRTee32cH%�!�*�(�l����.�LV�"�iPU]�d�H��*�PQT1+"������n\�� �5���Z��{y�7��[��pF�HoX�0>�M%.i"	'fW��צQ��_x�f�a��M���4&1�A�Q���;�nf��K1�GF+�"�W�S���L�h�".�;��[y�]u�|�*�Gr/.�u�h��RM�hp�JYɷ�;����[�\PKk+f�N���(b ��w���d5Zk�&7�fu�\c���t��ޛ�S��ƞ��W���Y�����_u��5��r�#~]�Qe�#"JM}�������}�����H*]���#��;�N��i��.�d.�t�d�2]痲�S�qF�q���tG��Q�?Knj��({��(P��*���|o�&�����N�����k�@���t�,p��@կ 4�(��٩Wu'q1pR;T ��O��2)��f�F���r.�:�b9���G�ն]Ek��D����erW��OV<���MeGm��)�w�	�\��`��`N�;�&�/�f�c�ض��'��Kf�6��L`��:y�ʍ�#��7{��ќ欤4y�ª�9���������#�#Y��Yڴ���[��}��с�sW+�R�I�#�et#ZS������7��2Ƕ�W�n,����#k0���LΆ�w���b%��9/���b���i���%��m\�kL�I��:`
�gb��@��E���&9:9����0 ��q1mU�=4jp�u+ta��o;�+VҏLW�����Plf�$�0�$�ņ��8&>z��.T0��n���S��N2:]]�^�3q˹���N����{m۹'�K|��TD��b���D�]�<�����c﬜6N����I�{zy���cU��̴�B:���sGOi�̫L��1L��3�M8�5ʳYӝ}�\s�A�o
�	Y�B���A�	�6�	�ez�)�\��O'9f�dm��2ˮ�mVz՗��9$]��
y�H�Z5]�y٘3L�Lũ�%t6z�ܳ��\� 
�ᛍ��o$o����ے�alW0FvX�����\�K7��L��:ѧ��<�&��¼�ΝV��S�Cʡub�O���\��=��g�I�x���ϔ�[y��'�U��<)�ç@�����M��@�#�T=+���_��<^x�bk��~�S/N�4c ob�3����)�̭�v�bI��|"�}��sz3d���P�jx,�@^�����Vl�;b�V�~�Ne�f��{2��:��+d'S鶈�0ԧȑ�<��ݽć2os��Q���=KվY@S�4(�^�yd��Y��6֜�;�tp�X�>G��U��\�le�de��S|�9jr���[�x��wU���u���ܪ���R�c�x�B���>��eT"[!rn.�,��ht�RĎ�|rI�����!�W�Ro�F[�P��;NRX��"��I@*�UD��f��#�EO�H��������S��֊�pU�c�ܐ��#��q+[�)���oXq�����d���<��l�ckgg5N�f��(5j���W`-��F�Uڸn��k4ԬZ��j�B�%.����s���iy��W{1������	�_z�Za����&���[��=��75�"I<s�}"�>Pc)���=�AgA�@�y���ܦ&L�G�C��pk٩p��g���D��5s���(�
��"�����{���"LA���N�q}a/ElFy�ݭ!���R��V@������GcOQ���j�)f#�LqM�Y���}I�7i��|����E��;����ڳ��Z!��'F4HK��uⱝ5���E&*oQ�{���cA���ݔ\�K��a;M��4���C� �.�Dk�ZPھY�e����oz13y���s�<*E>Vho.��nuuy�\V�,��y�����Q��{,tp�ݺ2���T��w.��4�Vr.�A�Vv=U��D�.�TVW� l�KN�㬕X�;͸/ ~b�F���,��-ܓt<J��ٸ�&;�4-M��i<� i����K\�1�z�8|��Mj��O{�{�|K�|���iqn���q[�+��ҟRcʞ�=�;qV�OW��������	�^��0�uR�˘c;,T=7ԷBTO1簅E�q9}��,(��K��<���"^2�����pf�Y��;�fuX��Cy!��ox=��΃�3%t��Ut�	���Cǈ�\~�`�vP�b�{̹�\a�a��K�DW�	�Ńyy�Ԭ��Ub����짣fl�d��Ȣ�W9��n���J���,FG�tD�><�J��J�jٮP�
�U]��>�E�C{��a�Y���'��8��*ck-E��R�)��i�a�Z�Xɋqn�wƄ���B�@��x�,<@�^��gCR�m���\��[�JΕu���t�ix�֢t=���26.����!�#�s��,#��8J@X<���{��:W�T����_�~��O��?�?�J�EX���A� BBcO��"z|Qd�D���������`\�{���v���++{M���kQ�%�XI ����VBB@+I0��f�k7Ú�u���ꅆ�)�"�l���6ʘe-[�!�c��-�轄"D�RUn�蚫}p�����l���Y�YJ^e&,N�^t��ౣf|�g��3ȼ���X�O>[�9���8`}�6�&���@�������~��5[�$���RHD���&bDH��:b*��]�?��捫'�'�=�b���sO�v?y�bv�D�go��C�#�o�Σ�IJPٌ����H�H���S#9rY��]�1EjG�f+�E�,0�[�|��c��Ύ�E
ζ�y\�dS)kҹ)?,V�"B'g��g�&�ˆ�����HM��]$��t�@�d�
`[�1��i�pe��`���"n�"d�UT�qdr�cŽ��ox=�c�*W��i�17�ڎ3t�v'D������s{��g��g�2�Y��*X��Ii*k^O)�;��#��7��Ɂg�M�\,�k��X̏or�~�l����U�p�}�q�A�7�$�2�;�Oi���B$M�RQZt��Ҋ='��ѡ��u)��f����#ȉ%��"D�ϩ=�SQX��'*���8�0��%��$�Ȧ�bč�C�7^�$'A����������"|Z&�U�"D�h�1ZLS1I]!ԛ_���O�u��(���!�N��~�	1%�<�{4w0����\��u9<:duD�X��I��Q�r�r������mk�ڏ�5�1����$s�d���_���]\���wM|�=q�D��tH���4�>߹a�:��z+�J�J-e�r���W�B$KI��˼�%�#���p6Y�׭7�l�%ۑ���Z3�h�8*^)��f
���v��ܡ���9�jm�#79�x�����>旌�SY���;��D�~��t�(ú3�銹�ݹb��OFe��j7p&��Q�QeVgٕ���Ac֘�w쎊%$�H��*I�/<�Ǐj�GUyO'	����HH�𤄒I�'[̜b�4��e��L�q��RN�|����3gR�!�`��<�Q6q���.�p�!I�r�