BZh91AY&SY�yG#��߀`q����� ����bCY�    ��D�BT)B��R�D�R��JAI
)TJ�JTD(��)H���TB���H�UT*��	$U/�JT�H$@�%R��)AHU�H���AD$
�� �*�����@���)P" �P\y�%*� PU(TURUH�A	PR!*��*T����*�*�% �D��J����T��J�**�R�IT�����K@�  f[겶�ڔ[)66�ST	DU��(SC��V�̚k6�띶R�QTQ�%%��5UR��PP�ն��:%%%P�2�DJ��   3�IM������%K���rZ�I-G붩tҕs�uХ5Wf�t�$R�wb�T���,u�Ʃf�t�)Ϋ8�R��i�xUH �)ITEUT��   L��*�.�B�!�JJ+�;]wn�j�7rU:���/s�mT�lj�稪�JW�窔�Dz�=�#�*V�M�o{TRz�-���D)갗�=$�IA*�"���  g{�+�V�a�_w���]n��-ʮݲ�`E*ίy�W{"�F�o/^�R�K�_y���XJU�nUu��K��J�ضn:}�ER=�<�J�׻)���QJ�JU*R�UD�|   1��ǭv�Z�f�{�z���Cr^�R�6�����|�{kmH�Z���u{h��V�����H��ܗ����:p+f1ø]j��%Ϋ�E�'�x�P�)$J��� ��  g����J���P����n)�[�Y�C-��[�X]�Kj)n�u�U۹��8�J����*JT��qT�*��]�I]wj�}ޕT@�ITTD(J�  �|���ګt9F���v�-G�V�	���j�U�-ʥJ��s��R�n��(T�N:;���E��.Kt��֍.P%U JJJ�D�J�  wu������\: V�w*���q�PUc��Q�Kk�8�Р7C���n#��2���!*���T�  �P=ve�8:q��($�wUhj��E�UA֌�c�R��� ::'+t��3] n�R�t�*@��*B���  ���-v��P
n֛� .4��ꚹP+\cN��c�.�u�P�Å:
ɀt}�  �"
�*R�0#  CLL S�0���@��	�10L&�a�$�i?$�х3Hɡ��Ɉi��JUOT @    "��	ꪧ�       ���z��'�y#�� ##~;#x�6�oy�*oJf���Nҹ�ι�s|�7�g�݋�'"�#6�+�" ��zu�
��*0� ��@]�`��?Ӯʟ� ��DA�`����J�� �"������>3 �u�de�ʟ����X�2,�	���+��,��������������=dXC�@��=a}a>�}e}e}`_X��W� �������=aY� �`Y�W�W�OX� ��=dY_X���=`3/����+��+��+�+�����z����������������=d}i�=`Y_YC�W�@����=dY��D�(��'������ '�(�������� z�(zʨz�"z�(z�z�(z�zʈz£����(�a=d=e =aT=`=dD=dD=d=d@>�OYTYd=`=eE=aT=dT=aD=`=` �e����P��P�������D����P��_�XOX OXOXUO�@��A��A��9�D��A����Q������A��S�_�A ̂�����Ȣ�ʂ���0(����"/� /� '��!�	���=`OYC�T��=`OX�aX�T��>���=`�D��}`��d�eLȟ�)�������	�ȟ���(���
zʞ����/������~z7��|7°[��T��H�,;B�n�L޽r����d0:�%�z��a���D�T�`[ƯVR�IO�v��^(��Qݗn�ET�%������,�Z-]%.�l����ɹ	ƭb�ݼ�f��9S^;N�t���ɿ_�-h�cQ�7�{.W2F�T��,�=kvV�M)P�e�ܫ�>��o.�ۻYL�n�}i�\zpB�y,\��v��w%�>hق�d{L�Sݧ�2:fн���=IH�����e�W�Ĺ�KA�p��w,��U����ed�E�#���U�U"�.�œ��if�\v�"i�sX�Ʀ�l�h���$��-Ͷ��� �Bkd�Wun ����EC�{zvS�2���	�i��������i�[��/��h�#�V�i��`J��̬еR�o�ub���b�Ah,;cA�]eB��N��,ڑ�N�!���]���X�ݻ�b�T�a:�4�=b�i4l:���їhd̺w�Xz%�Mѡ��̲���-����Yhd�l��SJ����-���;���q�҅Z&�(]�#q�Ѣ��t�)ugb7�Y�[�y�t>!�ٔ����TR��8N2��b�	�Q�	�[ya�B�tѱX�1�L�Sܳ�e���M����
փ۵VP�bLׯ�M�ͺ�eL2ؐ�դiP��2=���(��ي�\i�e4��-�MM��f0 6�ݫ0M��\123i՝�U=���U�[VR$�g�NĤ�kl�'(�Shw�A6���L��/6�RŧY�e�ͭ��BHB��Sɯ�,��&��6���ݙSQ5�����E$�ْ��y	�>�S�I�/��H}r�<jcN+4��4K�+"K`X��Îѣ5Z�˄)BkZ�Al�"'0�wD�SL��tPN��	嘪���fj�����k&�!֯\����M��aU���,��@��������n�n1l[�`�� i�5�ʼ:R�����9̨ �Bi"�^V�i3�.��p�sa8"�Cj%l���Sړ�a�k_����1���u7��iA�ڷw6%L�J��.���i�	�ǐȔ�$t�7bbh)�4��ܴŝ�4�qӌ�e7��c�ʐ�f�M��E���e��5!��1VS�Ƌ�")f��I��قa�@L����*d��Q�Ɍ^]�5����ZN�i��@��Z���5�v� 1�7!�7�K�u�@Bڭ�iA/f����7,��D�jMt��q�F� ����oV�����z�Y���Wh]�KwYfe�/�@p��Ec�h[#4��PIi[Q����e�G�'�U���M&���ճ���V=V�6��*�D���m%$7q,����˘)�H&�hU�8�VC)=�Zi���dU������R���eA%��z�I*���/oi4����Dk��U��̘�q�l:���2E�p��t����n[�5I|�t��g�a`�W`���&�o�p���ˊQOq��t(���M/n��٣.�V1��Ĝ��0DXƕɓFH���w1f�[o/�Em\�[z�*#e�����l� J4��#��U����7SWX�~����hS��3P���R��Rb6��a�-1a�-ɲ���tQލ����1P�OThK|��2�i���Ka��pPd�MRB�(1
ͻB��`mU��׎�N�������h%L�wuwyQ�x�օ$ӡ�]��wl��:͗�,��	�V�oU�+ص֧+)좂�������y���&V�U���+�˕���H<CjV��ǲ��6�dj�V��Ů�t�� y�24콲�$%�[�RH��e:l(�j�.�Ӻ�.��]tp�`Tk(]D�պ���Ml2Y��-��΢T�6]�gX~פcI�i�A164�4$hƈ�w�KކֲS�A�(	��<�F]�*�D�cn9u5�����q�*�k�����U�l�Z���vJ(�5��D��m��"�f�S��)�HF�V�<�.�P0r�F��iCLG�5���.aYxDQ]r�ك^f��N0��WI��c��	z�$���H�xLH�)Iy�ڼ���iT��l��lz��9�Vbmm���q��+��b��յ�e ���0���-6��F֨ݚ�&GZd]�)�Ih-9yH:0�n�g0[T��X��|$��o�4���[�#���V`���8���nD�i��s-ڼ4H0꣊�f깬�M5dS'"h�����2�ɵ�ʦ��7�؟Wh"ɛ*����XV��o95�H��Kq
�+a��b�oj&�	a}���t]�6��� ����VAv7)U��Jɋ*�\�oo�rYkw�Q�!"�c�`^���-�XB)5���KU�J��n�MwlhOZ�=��N�Ќ� ��D�P+JYA�db��=X�ݳ�jGHҼJ�IFV2���aT3)k��"f^��mD��fe���i��uVڬ�#n��Uz3�]��1�-�����*i�3-�V�B;s44\�)�*�y��L���z-Q�`B��!^����T�k�l�M���R��ڳdխ���VDpMb@��-��w*%/0�B�,�s#���+6�V<�#-f6�1 �ɰ�w��!�)��CU����h �
��#xP�(���XO/b�Z�+2V!�yB7��	�Lz@�2�6i���(	�%]�CZ�_�ӻ�j�J��x����t);4�Om�m�"Tע��˟QPZm��ڪ�Ȇ*����ve���C	T��ϓ�2n��>נ,L�vF�H�����DC�:�=�r���㗏�AdcR#N��.��E�6��1�eVg°e @'WP��7]<�y/�n��v�kmJZUh��؛�aTУ��ZP�Z&�Z�!� �q8�r싲�ۚ�8���Uv������n؍I$�y�IrQY6#�Z�n<ԙ
��ە�$��v��x�\���1cna�a*��t�u��]���w)MQ�s,`)�������iG�p�tں��%"�lT���iP]ѹH��Sc��oeh4r��ݭ'Me h��Y�W�ZB��X4X&#n]cX�u�b��A�4�
����KM�[Ku�DfQ��θ�7��jSz]�EzΪ���-Cy2�Gl]YL�c�K��IZ��B����<{�P�q����,G����wJ���k-�@6�6��ݍ�z�c7x���$?�B����a�h��2�'3���J�� =�vJ����V���Y�J�M!���t�2^�m�H�����M����*�b^"N^���Z�U�%EX@G2�d��,�h=�J�Ů:c3M�S[H�k�ؼ���Q�J����!���;��/)�hbj�U�S2�Z�54ѡ����h=t�[M�qϧ�/M�շ���^�q�1�mZ\/.��<n�ԥ?{|]�`��ح�������2���Y
uzY7��OT�P#CM�]�b�X����2!ٚ�:��$�B�w�WVP���\�ՌɘHˆh˵"?;P\�KC:��wFˀ]Ёޜ��\t�������Թ����[��[@e�S5�����j����$7��6��p�V5^#�|8�]}A�V��ݲM�rkL�t��˩KBz��"��@�WYK]H��@ݜ Ne=�W���v�oʻxF��eG#M����O/3(ŋc����c9�&���q4Тi`��Ŝt/+ �X����mL�ք@Q��Vu��#n�v��WqQ�|�{�r��3�ڳ����,c��@�X�wZ>y�\ �e
:Ȭ����ز̰��KAêQn �[�U�d
�7�5��P�Ф�aL��#+M��,��ҁ	�����3^ѐÚ��)�W��W�%�He�{����
���3MJz�{Vc��ۍ�����sX��9Y�XT�J�ĤQ��ě�n���36T{1�����wr�dhb�;�O� Cf�_�Q���jkE��ݵs(-a*�p�V4���3��+pk����I�̣ ���<�����0!Lr�^Ga��G1��P����Fn+:��W�N0�ɚ�ӣ!�eL&e��/]ֈ�����ѧM�H�A����4G�Jv��h\�y�MkU�+��g���⩚헂-`�,eܷ���.K��#ZV� sb�&⭽Sv=�W������[�������h�&7S�Y��l�O1@��:skj�%�m&kh`H��j���aK�ks^����Z-C��*��%:ѨIL���?Y��9P-�(c+r�H�ͬ[m��Da�AfV��4]�u)�׍D�0^ȯ�w�W�dY�����ҮE35<w�Ň���CL;���)�U�(Dv�P4�9�4����[*Y����ӆ�S)l@�*�H(5O"vrҭ,���sf��׏`�8i5kZ�Ф���$Z�5n^U�+�krf�q�ӷ���J=ղV�2�m��q݌z�&�8�`jKyYi��z�-!XP�٫{Q��p	.��Ɍ)v
�Qş<v�Z�1�f8n:�.2�u�*�vn�ڠ�4�!Ǩ�&AZ`�F�H�Ժ�)X�M�Vi*�lI�ћXSƾ/�x�6R-l����t��VZ���I����r(�^M*a�f���fikC���Ϸe0f)r�� Sn˸���C��n��U��^K�ƫQ��P/c��2
��� H�Kko �w#�}`��Y�rL�!ԅ��:�S,*��ј�mų.]䣰t��>B���z(%� ��x�	v3*l9�V`�z*%-7�854%Y��+"TAn�m<�#���	ڲ�9�cr�iӻR���}���n<�[rdc�r+����f�Y��@ܣC%�*�%�]$4�D8IO%�%ь݁���7u��x�Ij�To�`WX��x��i��vQ��)����Pk$U���B���Tֲ������
�÷g畗mb�el9"�U�M5�ZЎ� ���ѭ�u��@j"�G\N۹wx��):��f�o`��co�ͧ
.��&^�
����64n��Դ6ll/TՌmZ��Y�J�B]�۴�����M�Vmf��U�� _��Z[��X!��>���sR�I;s`{�5�ɶȫn�&J�t�!h�k)�A0��
�1L�̔�*�
S��4ӥ�n��O��Kp�yv�j���Tv�e�P�Z�DM�J�e��N�f�J�6l�R�10�iGE�C�r��J.嚩p�&Js�����!���	1���IR]n=l:�^���
��Gu�&m�p�w�ik*\�]��[�^�X�ѓE�$:%��[l����Mi�I�+di3��G/�^Ix���Y�nJܹ+Z�6���R�X�0J�K*��75���	�V������u���U�'/R����3T�cJ�����a�wZ~)U���v��`e��I�BPՌ���<Be\��Ԋi���&n�Z�ZE*�����B��z�bKLJ�;j�Pk-X�ђir(e�@B/5�j�rʘ�x���8�h��m!�(���'��)50��R]+�:��ٌ�:����*Zge�Ė~��V��X��k�*�)�PDM�L�j�C>����n݅����4[���� ����]��f�K*��R4]��ؤp��#�/�N��z��k3n��8Z0?��)^��&��5;������N�w�ZeHs#�&*%a���������K�WAyʑ�f�$��r����k(�.�É;���a�]=ѹ)����r�YX��F&v%���#@;�34Z*�:9�����v�'3STN�ñ�{zU�Lb�@������^֨H�/�+�`.؃j���o[Ķ=��߳n���P�l��J1S�,�l��ʊ���P�usB��R�q��`�%c5G.�Z�u��q:��i޴1|�钡�0bݤ󫲜�,�J�[;TO+ɺ]*TXW>�LܗiѺ��Y�ʻ�A���5�E�����&3�;�),6*=ϵ�˗��vUa
PcV]唬�#]'�{t7o)��=�֩1e�6���^�׳)�ʼF�
��b�@��
���J	L�˼��!xaj��SM,�R��Cr��8l�%�X�&r�,�+`���f)�r�v%%*8�^*��d�� �Op0�5��J�,`�J�Ę�^������[�e2�ɖ��#ZT�ɁmX����V�26h�`��o"B��*�j��v\�������QW����J�	n����Wv�X�	�kgE�(�v����[�j]���M:�5��l�fŚEjM;��՗�KZN�(0pU���Jیh۶�3��Ҷ-�����X2�32��ɭh8 �Ѣ4Pu��"�luvd� �y2-X�2���y��x�XresNnn��,���%ɩ[մ^��,ӒM�m�B��/��C4�t�mK-lX��)���H���3-(���+P���v�w��^
M�
^��i�䫿�n(˩��b�N�߁6�k)�^�7ڕ�d������#NE	��z[�Pj'�]� ;P�㬡LZ�],1Z�'�n�v�k4�ۦX���V�wt\��Et��v�\!�#u!�pP��ЕgC�@y���<3��@"�!�K��i�l�˩��.G��*%è��<f�DY6\"�qD�yi���08#� ;�4��Z� n#�l�U�#Hdf��`�``�h��2� 5|�p k��T*�Ⱜ=e�hr=�و�;i�:
���e_h,8n���ţe�5��zy�#xy��3l�	������<Eu������в���`w#XW�;�� :��$ #ģ��:JEq��t�7A�J7� Z&�������y�G����ɯ}�D���m?��c�8�%Uw�ĝ���͍���j�����W��|Q4�Sn��%ArǗ�ع��meh@}��W#�$�ܕfq��t��,���\�nee�&��2�1�y�킬&�NiK*�	A���,�"��Ϧ���2��6��d��T��O>���0Q���;����}��8��;�:5���ʻ��cg ���4
�� .\����\��W=�ݞN0���d�jcv���{N��ʽq�jg;۷��)be��śʧd9���ٗ�wf,u�4�B�ݺ/�I���	��o:�:J��k��WGJ�X�����G��F��V:,��v�Y9�CK $2u������M�une�iK��/�l�Lmu�!���7Y��{i��m��;vX�.waEä�����o��ʈ�Z�bfY%�ZЎ���n�3�&��2#x�1�h3NOZ=Np����WXݪ�M�!)c�Y��p]k�%�W�6���(��y+���1jR�,��	�2���Z�V��,���2�1� ���0V��]�O��������ܷiY`uD+z�S_m�H��p����4)=Ӑ��N!,�i�P^�=Oj�"�9���8���ǋv޾���hu�7��1F���W�;+j��@n��v�@'���}��
�np��U�v������u��V���P궉%Nؠ�Ghr��]J���b�*���IwV'n���1>1�(����
��w|)���mblt; �ѶcR�u������"I��^qŒSB���p��ݥ�.����a�LE1.8flFKV��u:w��C������H�٢\ͭ�Z�8�u���*�h>狫���ƷAьv>��\���P��'�]^	���oW��T�ם��6țǉ�m���7�M�J�a�^�v�*<�<�l���ǼM����:�rA��8&u����(�U��� ͠��D:$��O��|5�r���h5�֣�^��Y�B&�]ۜ�_v\�:owy÷�l�˶�B�n�;"[�|CUMc�)�u�����(v���fҥ�C���+�Lr�+�J/���i�)����xt�u�i�gCn�	��ꂤ.�5Y�w�A�c{�Y�j�nd� �+����f+8���̝Q��o#VUrGE_.�Dxp�H�Vn�\3�p�n��}�r>�O3v�ϲ�ns�#7�5�E�Lsk&jϸ�iX(��qc���Ť��'w�աu8k%�r��jڡ�^�N�^-:-R��+s�=�VoQ���N�S�r�ẟc���1��,%��^����.�4�&��ƥ"k��`t{3�����P��y��$��j�9��6��;�bh9���š1�=9Bn�vn2��_d(o	2C�J����E�r�Ь+���/pgN�*P�У�t�Nnc�:؍��.��uϢܓ�p��^8�;���&P�Ί��,S���b�젱VҮ�������^S�ݫ8Ǒ���V�A{��{��w� ��[���RǁA. ���a�.V�c��1�Uz�V��v)ֳu�'J��h��Kw���n>b��B�	�"��f�t)�ǻ��۴�t@ޘƀ��� �*�?�{ט�KO�p4�jR�Z��g%D��=N�S=K�	`ܢ��r�R��6pa�\&0.�Ӡ�kVBm6k��S"E���;���	�̾*���̔�J�`Y�#�[��j̰�n����
m�y��1��MᚗY��Ԛ7�,�Ứ�%$��9ȹ�4�P��<�;.��8+DWK]d����&���PQ��i�GN��#c�F�¤	#1�.���5vt��80��B���n��r�])�{�mwub[�U��"��ؐ��L\kqt+yMT��^Sux���p��J/������+-A2u�i�4*@��z+)V^�B����p���9���ccdWפ왼��wψ &�h���W��=V��5�6>\2Q�Y�CY�Ou�v姮��wEw����rˢ���\�V���%�x����i�\���vc�+Z�;���L�O.^��y)�䤹7��xvv��Oe�v���3���H��Ŕ\�c��$)����t$��+)�uۜ9/�v�|I���*(�ɽ-�^<$x����7�gk�+7ٯ&wr�5�G��Gl�ybJ�����um�n�_D�6�Z�X{Nl+��&mZ=N��*�,��gJ����ۋj�+7J_�_��쀓{-��N����~G�d��*j�7����#ZE�+���Үj���n��ب�X���5�+pۗ6�����w�ҍ�����I{��lZȢ	Z�X�
'��7y�yt��XbڻǢ�*��Ï�Բ^�D�Ӆ�u4�z�v���k���H�4��Gp�ʝ���u�nVgwX�ky���SLs�+�gu�ϻ1�H-h��W�.d�|�h���Y��Ԏ����۶9Isr��};8\ucW˫�¹(X�b��6���F�6�gXi�|Pux5�d�9ʲ��j�O�NZ���L�v�0����xػ۫��(�ݥY�]�A[��8S�5���_��y>kmb���ǽ�F���O�W7a�JCQ��s]e��&��wQ�<0q�{���q���4�3o�ݫK���dzl^R�5���|�I�md���ԅ�\�W5�:P��k��-�)�1�;����S��dd�c���v��7׉�y  �p�G:�3X,}uau73���2c���I��hW3�2dׂ�I�0��u�61��0��X�`�������ZQt�0*�����6�N�]�4�N9��ʴ��8���4:b��TB��ugrʼ��0�#W��8�:~��Hho���{��U�Oz]�Yv�R�Ȼ���E��M#������ofhB�̙]��"���(n�,�ĠTwGr��.`\t]�W�+�Gjf.�7��Q��F�+�:� �p����)uL�����Ր	}YۑTu�i�Qa�G{���H$X���kԝ�x��׊��[�^�=��ʱ��F�Go\.bu&�n\�ǵ��9,＀���E�k��In��׮����F���i�Z�Р��;�kz�c��oC�Gnl�Z\���HGc�Z�s�΄q��dάǀ���y��6Q&Ƥm���	�J�O5�qlk���p����/��,�^`$�`��Ռ��Գ�7'&[�],�Cځ�	;^���uf����qY Q�VzP�s���|:A�f�]�~� �ڎ�7��F���p�9w!XV�s�Ә��lY��V-w>�Tg"�����"�G��[ۥ1�I|�R:d賮ݾk�`�M�
^�cA;`p��}9�F��W��
�ᙜ�ѷYD�3D�9%sT��հb�DZ����Ut ��T�y�X�:��P�-܍/�����r�I��K��L�ŷZG!�2_+�.�ʕb�ͻ�ҵ�%Rl[C�Em�}����V�FX�h�f�::� d��B�;9�]䎳(t#gk2J��l-����D�������Z�e��˰���u���J���Kͺ����Oq�vlI	��B⻆�\bjy(�x[�s��ew,����Jۘk�>q[�;��}� ���:�vB�K0m6z���h��t	;����\��'쬶o�^��C��8�,��ò%{t8�d��b�:�h]#�H�w�ve���ǧ������H��+�L�����\���s` Ү�f#ݐ,�a���qW�z�U���1;����	;yGC�/����0����C����)b��ۘ��VZ|�5���G�:f��t �S%�e��Jk=�f�FPr��=�mHG4]1�����\���Y�X�ْ����Xf!{i_+,��[v�6���p:�U��������2E'��:�w|M�Ʃ�; ī�����3�w�ڧ`����ޅ/�kzn7 �Wr�*oU�u�eܶ�e�}K���NY1�μYb�וv���`aU��/����}8Kl��8�b���1�EAR�o+��T��1�Sn��qԕZ�F*�.t�E�Ђ��P�e1I�]�+N�Y�q���cW*7XYh!\�oK��Iݩ�Ry��Y<�<�3Gh��ӝ���8',|oH�i�
���r�ӱeS�׹uۛ{L��ciT��C��}g���m!��v_ϐ<����h%B��'�9�6a�h}w���v�h)�v��6�r��#�9��M�E:7y4nqt��N������ωެ�+M"��`�m�eC�.�Z��M�$��E������t�Iof=�ة�����|ln��i�4x^#�[V2���5)��a��03D�.����])G������k�U�r��"V:��5:��d����Z/DX4�sR���mt��v[7��$�M�]�X�]����h��Η_:�c���z��;G�6���+6�h�aj﶑L��G�n���}�"��v�i=&�)�C�n��O�f���G�-��G��F4���WgS���h�`�w8����)�u��!���CE�7a��S��FJ�l�8��r#�ʶw��C]�QY��OlU�~�ۣGޕ��W^�}�Ԓe��3n�\�����Z�0f	sT�����Z�gZ�]�G�^o�Z?i��Y���m��ݗvƅ�34�ۛ�!��'9�[���vx��V^LMEa+ǽ��;�����p��s�@Z�Z�g#P�C�� 
l�B�B�Ytje#*���=�#ˮ$�x��%�4b�2�Ѐ3J�8O�#����Z�W�u�
�WV0���Y��@����w�2����M�4X�W5w9`x���Sz"�b�z�]����k�K�6v���u�����}SC�mwoZ��Iv ��w\�}� n��_Sj�m6#�C;;���o5V�W0\�&�]�p�v�� �Y;z^[��P�������ܙ]7-��A�@eEq<��"�!�x�ʵ:�[������=/���+�8��b�%c(�*�0U֊Ɠ�V�1"r6�a�9y�N�5���N�$n"3��c8/6�#%4�����5������gP���
���Ԯ�v1t¬��7k��/`՗ʐ��*�軔�B}7j�W;gR4te�;� m�;�s���ֆq]�.�voε�ι���dCFUƢ�ɛ�]����p�Ԧi�̓��U���P��|�!̓�L��zd�J2^�yKzs4>c��X�V:�2�.Jld�>��}�{T7b�:+C
mp�ĖS���>U�N�#����[���q�ޫ��t|��f�\Չ�cA�����[���m�j�3�;4=Ùd.�"�I�Je�kF�m���v�"�j�Q-�UqA��(6�s�x�Ћ�wj�wVU�4�
CV��W�\�3� �����N��X(5-��-��Q#
���`�\1JWK%��5��uin���S;2u��4�'��.�r��1C�[g�.K^����]f�ڝ:���Aq�n��y�ʔ-�9� �\hZ��oΖ]e⩙��Z�LT9���O.�:�8j�'�[.냫��׶�ٯx��f��{r�4��� ��1\�{�f�D�.93h�\�tAc#s	���v7AU�&�ubHsJ+\��gwf�,Fa�5��Z��wd�-����q�����:�	�]�{��*�g:O`S*�6�%`�-s9r6�9��F%�7�tP�]���]���[d^��7Pt��ɚ��+kL32��A�a�n;-�{2�<�mu3q�.��b�\X7:�ޗ��W�ƗLg2�����Ý�}�5�e��	6m�ٖ��>��n�e6��
��\(ct/�Qj���̖5й���+�C�-���^;������]�`=B�)RKΘ%JV�kx�%�u�Qڌ	�Y��\�fm���T�9���(lS��.�p��cK�b�w��@��.�3��o��j�'��]H�K�bU�]Y(b��X��"�EV��)	�Բ&X�s�u���w� ��~'WG\�k�oc�xk9wW~ܱ�`����z���Y�t3���B�h1~5�T��b��/�Vn��7ɷ�el]]�;}rK(QBS�@��,k�ɳ�����l�}\N�f,c����r�m�TUbM�hn)�B�5�Gyt=��3�WZ�m7z�<;|wZ���;�̀�r���-um��J+Ψd��Ji�B�Զ>����5؜�7{�ӫY�n�8����M����v���ʧL��39^m���M��Zl��Š�P�bp]�/E&�f�����'u%�u�+z��}!��qj�#Թ��r;(Ǎ�s9*WZ�wIuʦU���:{�\�[�]�7����w{���.���5�5�sI6oYݜ���t��Y��!���\�HX�W�O��8��C���kWv��T0v��9c��xU�@,V�����y�5�1_u�I)�ڱ\h>�M-���\�;b�>�K��(�k5�[�)@���$��q�g��8=g��,�Ktd��l
�v%㝶yws�<�]`�\xk�w���<��׼݈�6������� �i����B��$��]�L��3%�gH�s�}�H��@ّ�����橒���2�9P:,f��D[�8Y���P��/���O*Q�;A�8m݌Hĥ᜺�_j��r��ѓ�r7��R�t*=v��fܜΡ�
jQ���(�1lͼ��j�m�N��b��w\��Q=�u׽��g��v�k㝏_u�s��C��úi� 8��ݙ����)Λ�wuW�^����{�~BR:g���e:w����� S�Z)K��C����|��!I�|��GJ�p|��	�'�'�!HGЊ*(�.�ӵD^Z��'��PTQ}q�~C��'�7�׷L�r�w�U����r��HQ��^,�G]�ǻh8���rp:�Uz|qui�v�_.�ф=�V�������o1N9��nV����@�C�Gu+G�m<�
:�"�B��7qP_T���G,%M�hiq��W.�GWWkH�B�x�
���Yqy���D��ڹF���&�^}�Y���Ϭ֮}F�,[��ʾ�n��7:?���u�\�5�rJc���T٦	o:VP����ps]���9��NTۧ��t5y-s�S�/E�0�0 Ä޾���a��r3�_M<��2�-q�Iҩ�ꌡ�`�ೖb�t���LWGt�&8�F���Q�����V�̂6m�s�����}�V�Nv�]�W[#D�Tv�:�������*���H�����r��%��h]gv�ۅ��X���9.���'>���Ք:�nr�(Yv��.�Uٱ |��+Mb
�E}L�A0��+Of���cmGtT�ϭҤ�8����c�Έ�a�umؐ�5�`��۬m��¯�f_R�F���[�|:o+�{�ȩ;�;v�*V�B� �Ƹ�S,mX��z��57��E��7y��ڳMжz�4-�=��ڱt��P�y�L�K�@�}�~Y�-Z�`������wU�@҃����1�Z)p<OkJ�wqs�+�LM����{��4�z�f�lt����z�ps���'79�2����|���aw]��,f�:ZB��d� �y�f=�Z�%-��7W��򹫊��<�
2�P�wxp
�����cg������-��a1[��4
�v�s�Q|6�w)�hT�&�
�'�w���Z����6����c"�Ru��/�W!2(�	�4�vL��Ar���!lӴ� �B����
"��t�R�`���Pׅ�\���'��u<SF2ٺe���V�]������m���]���qZS�^�-b��*�!ۼq7Md
�s��<\�e�9�%�n��T�-]3�1�@��Dƍ�9{}�t�`�&.Ë��x��e&A�ܱ�:mN`h����O� �|1�LvSIJ�^�B�d[t�4]6�g�O(��]Ϥ�z���;h)+�ؖ�;w�"�S�h�!�<j�'�ڛ�ݫ֕ɳWm�] �	"\�/S�L�f ���.>5}���  ާGlCǞosi��٦���|X�k���7�*.����0k����I�k��
�nȬ���w��՚�t�N��<�U���V_V���.�Mo_+���?TH��� ���釫3;�G���ĖݫS�|1��Q��"�{|��^�}لK,�T�pP�F�N�'[���]���*S��P��T��;���."�@�Lqݮ��$��گ��F��Of>+ ��[om�.��[ҵ�op�yk�B��!��Rz�g����﹌��w�������P�#Nv�^e��5ú�Z�������%
��(Δ7�`-��ʒ��f*�s�W;K�yێ��}[�ι�
z�\'M5�Ԫ���fiZ�ÏZ�a�^�@���[�u��2�آ�s�*�Z�BQQVP�n�7R�DOC2��h�d7��`h��V.ι`B-Z�D�PD����[��f]�}�0�`��B� �:�p��Ne�,�)e��W�<;c8�sn�1j�[��
v�Uw�NQ�)Y(򮍞e0kX8��A!���U%��!2�WV�]إ���5����EݑL�.�HQ]�q�1�~��Ղ���]BL�[t��bV�M�
WY�\�#�8T�Rw,��M)D�.�6��0����T�kE��9�%��Gj�m��n� �ZYD=�,�A�@�;P�X6�f�)Hzg\�_&c,�Q�V9n�|�vI�c�ǳ�Y����{�r�s}�z�}��9O�t>
�0��c5�h��q�������C�\�?&5�赘x�-��h��\�� �Y�K��̏�@m�X���Y
��c;����vwlȮ��켋�]��BZ����pֲ�
���üH�2��e��Bw}>���w`Jt�s�ҽ\��L|�hQ�Z��PE��Jncd�6�l�оt�ܛ��JV���|L���6�2��W�d��^r�[Z�m�#�Cw#�z�;�A]�c˚�\y<=��=��ٮ���l�6m��W�Y��������W����8ᩢU��r`����� �����Uyy�VGqlU���)�cD�8O���Qyb�� daֽ`��|��U��P�3�����$t(�0�cG.�Y��d�j��t�?��a�j��T�J_$>�2��9�m}��[#yɣ����|t�L�xӠ��(��e���yQT۬p���T��A�e,�]طj�$4�)B�'��t6��s�h*��2цM�e���@�*�CB^��j7ݶ+z��*�3�W|:������k���d�4�\y/��[�;��Z�����b�0m�Q�|b�����bt�a�f6mCrV�qt,�e�ºF~�wB"��y8s�@���韀b�����Y�����酨��\��ma$��	��\�gl.*�����n]s��Ĕ��z���o��_gWl��j+���>���^�1;��*�i���Ș��jr.^�|�%��9Y��n�i̢P8�Χ!���w�(Gr��jǂ�jy�yM��1����f�d���Ư�%�WE!v�#���o]v��Gyp��3���X��zDK�];R�ûs �u&M�;;�(���j��'wO��Ѯ6��� \�p4t�ܺ�U8o�o6�gl��=��)3m�W{�5�}Y_Fu�;P�WB�GF�#���3���ߋ�����ܼ+B��֖�K��8���ݎJ+u���='�yY�Yu��7|8�B�*&
V��;%���}*d�l�[ط�k�w+>9�&�2�×/$<�������Ȍھ�t>bs���<�2�[{48�G���Ӌ-��3]�m�D�����M�g�U��K5�./yo
����M�R܂�:�gu�j�|�D��_R���'G�kopY{W���0b�r)�]�A�kV�S�C�}�{]�R��9V&��rj��	Ͼ�ӕSi���:Y�m�G]�p����7I0iJھz��>�Ź��]n���r\;�s�ڷ63���e0g������n����;J�N�+q����8��|2N�����:3�+�V�j��R�%�r�顐�!{\����x�+Q���&��$�c�S^�"ѻ�:X�K:�R��],��<V�A�����*&1$�av:T	ԟθ������P��8���XәNh��i�|��C����=�0\����!V��ܓ9���e�;Jº�*�u�J�����Nչ���Ρ�(��n$��it}wdW�>ی��ի-��g\�Q;��u��E�)e%r�9��:�l���¯a�흥��n}�vS��rf�F�t��]L�Ӯ젠V����;E+�ˡ�X����A�CQ\:�*�(�t�)ɓ�����/�Y¤���pd�-�C2)li\�0��՛U�c�Q�V��ga��l1в�o����WLu������C{�D��������m�y֧XlP�^�΀wTs�1�R씴�GBj���1J܇*hZ!�8ʲ���ي�I1��E!�"����F��7���!Sj�kY�aǷ�,`���,npw�A��Q�㔲��c�*򜶎��ݼ�`_.���:YS��@�/ky�@
����������;%��la��a� �
��Ň��;�
돓����4���\��z��c�b�?���b�Y�ݙ�;���%^f�㚺Rx��3*I��'t'��h��3���8*��{z�<�G5T��;� 
���<$��]h����X2�E]�n�b�Nq�ç:��ɡ�XN�DZ��;�ۓ:�Olf�ތ�\�Wv`�[j]c��C�����=J̽�b�˥��A�}��f
�4O\M��%��>R�5�*<��ެ�E�������H�0��7PA_qwt9�Be@x�2�`�]w)ve�<����I��U���d���>��żۡr]
������P���Mp8�c�;�u<:u%���rjsr�
|����򷲺��7KdJ�ֆ�P�f�V�5�v�Q��6c�kU���Z�r�$k�.�Xi@�;���x���n�u���"�2��T{�+�o3(�5��x�fin��wI�FWR��&a�n�%E�Z��ϒ0�We<�IZ�=
�kM�Z�n�˲:�wAQ���7��j�Y�0�DM)�����E6� m&gn�Z2]\�Y ���r��k�V2j�B�N�ZʸV1S�$k��2憭w�!��
j�6��I
��r9}���c���3����s�	�s{��>JJ�[��)pynRg�.V�4���C�ق`5cs�:��f��Y�*��+hW)	����F�}����S�����=�hG�^q�l�Ɗ�#b��MY=6��ZG;=\�>�h:4_�ԝ1�4���R�nj���̭fܠ)�bԤ��]�+u���w�;,tthb���ָ�:�"��i2%�Eʙ=I��1��]���2�;�$ۭ2�������ʆjN�ӽX��U�hת���q��#�WL�ev��R���mK��<�W��+�
���|r�
B��[j>�F@�bif<��K�e+�Yj9��yJ�1Nk��yt���0�����Ѝ]�)���^L�����**�gZ�U�d�ގ�@�2��p�}��Ա��\D�=������N��E����Y�PD�j���b���S����E�C�z��@)� ݰ*������g����(�H[o$\��ule,�j��`9�b��R���l���x�]Y�X�K����e_�x4֚��&�$6�C��h�V%h�"��]5���s�Nq[��7jڹI��p�*�OR�Tq��ˎ�	����+pުŽO�����ԳK��o;Os�N���)���\6G���w�&[|1[����oP��w�����u�-����VKǭ�A���\����F����$�7�o
u��k"ۓ�<��n����������K�V7!'�\z�yVY�z0�Tb�ʖ���~����Ky����3�k�����[GWj/i����)��a��N�Y��!�ʘް\D�+@�j1�4:�޺+�]J2�I�}m�h�uƫ��s6����.
�u�r4��t�;M���<YWo����{ef8x�9��n��\�M�xT�[q��jP�.��ǣ9��C��¯�u��i�7B�6r��g�k���Wv<��3i���Aq]iWJVj���Y�Pn3�
��ɋ���P�o]a��WL��#G%(�J��8u�E*��˵�+;X��*͇��^C��W[�%���TP��8�t�%c#�j�s��TSZ�����F@����w�q��bf�/j_o�kW�]�V�\0E�c;�;�������nsic�]3h��W+v��a����-<�1tu�*ݵ\���ᮮ�t"A��ݺ�һ+0���ܑ�C�&Pvm��"l3tô�e���N哃i��m�ܶ5]�cܬQ�^ֵ(�K����٠�y}��s]m͏36�u� ���{���),ٵ5]g_4�d���JV��]�WP�YA&5]�\��	:s{�W*�ޝ�kl-�i�rf��D�G魗`�Չs��z�]�\����͗������U�DMַ@o���H��]P�j�*�m�>:��qX������6����;O���m����VW�҃v���R�+�֠�Zl=�W9��{�:���JVv��V:�t�R�ǯ��R��T鿺+�؜k��ⵕ8��2��DN\�Ԯ����;��Č�q�s!mP��}�d�f0��Pz�#L{1�&�]ٍbo(6�,nV�j�r�p��'�e�euqJ��cV�t�����wG�<���"��m;Ub��#y���r�;����l�j�/M,y�i)����:&Ur�����Ya��n�K�oAy�qW������듵���=	�c:�h	3[rv�ޝ�Y��+�{\���G�3yo��.�1�Gu�TSV��r[��9G7�Z�������+v�Pަ��@[ʻ�����gT	Aut^u�4Ri.�F����+��)��(}-Q��u�.��SfM�vÀbaᢳ��)�I�s��	�>�Z��ܶ��p є�4%�=y��W�t���<4^�'$B�=׋��d#�_R$�:_@��(`��ѬλTD=V�4�`J:~�*�Sʴ���ʓz�G`h=Wm�N���͋vcw%�V41f���Lo)�:Wgi֒�m�����^�/n��C͋2�R[B�Y�n���ޚ�˳�����V��J�3��1��/�#١),Jlڵ�jC�u�66+;���jW;��'P�Lm�R�9%}ѻz����폣�W���o��J��k;K�#�Ӥ�ӕ`����G �\�왲!�p��!qwc����i�<�Ǭ��:��B�w3��լ4�YŘU\�kUw;�lԌ��M	oP�OA.�Jȕ�=��1���l]8�%��5ٸP�}Q+�lZ�2��n��]�Hj����Υ}��ww;U�@F�;5<�����n�m�j�Z�grE3)˜-!��f}6�j2뙬��Wq�8�n�'|���x![���b�D�Թi�غeD��K��I� ���d$���v�ͣ�a헪��P�����~4rt�%��:[ڍ��*�Q��^���ۙQ̖uE </0\U�蜭�c�v.vƖZvM���5'�oh��fmֱI�p����"�H���f:�(m&���\�j�P(�:"r�5�2*�:"e��^Rp���=��:�8����b��EYnn>#���.��U��v�N*���;D��r/�31G�֪%#a�`�i�WċVV�m�W���� |A�?~���޽��<�n�7��F�<��S����)�}�um���v5�xg�kR��N� *�m*����~u����m�;th��;�����ұR��V�|�4i�I&Y��`J/���	~Ũ��h��ПI[%�m�H�E�ĭh�g7o��'%�`�fX��5dC#�L7v��¦U��r&�+Oͥ+��dd�&��U�n�w���)�z$]&gz���Z��i<�5hv�pW�`p�V��Ԇ�m�u�o^� N�ֶ�gw϶�!��(�R�"�B���[��wf�,a��bg{;�}�T�.�Դ��q�6�.����uIY��3[�?����v��sy-�y;t�qT==�s�\Y|壢b�/�˫�[�Љ�M��`Žt"Ǚw:��P-��UO۝C(��q.5�۬�)BS�4�őY��[˙w��v��֥��:\�p���k�a�l�jp@l�hP�f�4 ����t �L�Y����*�r:�eɩ_B+�` D���(��1-AV���q��7t��ә��Dx�6ob��$=�]��M.�˝�oσǖa��ѷG���ٙ�j�w%j���嬼��g�ܮGIxvF���GK�I�;�\\�Y�'W[�B�ٶ輆��s^��r+`j��3%e���m� �j�v�۰�8�Bu����n1�7�p�rC�%v�+���4����e����aה@�R����'7����_K��KY���`B�����ڙz��27��w_]�-�w���ρwQ���x[#A��e�/�i1D WȀ�a�I�h%E��! �_0�&�(�ӯ��D&���hJ����@�B�� U�(��,�@I�a���.2��iA晤 n��� )�'�L�)6R��)�����ѪL
-�J�$��y��γ����AGX�j

�������QAAIZ5F�M�TM��V�趈�F�J����C��i6�D�PS�]5��gv�Q��[6�j����٧Q�ѹ,��Pv�X��P��JQ��QMk��G�;*͘��X�Kj��XM:Q�N�
*�h1^ZK�#mmZh(�ֈ��������0�%:��łں4q4ch��
��'�1Ѻ�V��w�"*5��+N����T��V��)(�g��U�f15��,Ol�cmTi���4;Z�6�ZM'Z��:0��k��mgi�5Qю�m�����T�TD5��l0��Km�V�͎;���K�TQT���"�A��c�h:-�����A5�Pk��ӣb�n�h;Q�����j�v�f��AE4;5�֪�ti���'ZR��b5��y�'w<�:�͠�A�M%jڍ���:������b)�>�|��~�닾,�
�DQ �A��c��z�ھ�����k������THԽy��L|��}ƞ�n�M��/��E,�Νuwn�7����_K����v�yn�����Z��bז5�^]��_G��v�7ݙ�Tg\�aڧ��w�\ʡ�Ơ��6s6{R^�r1xLI�^t� /H/'p駛;o2[?C^��y��r���>�{\߾+j=�+���� ���k��3 ]S=�n�n���}����!6`�۩U=�}n��/WW��;j����o����/,%�Z���K{�l�W�E�6�=鴺����j��:��8ǫo�f�Y�Y=�}�b���E]�7˜=��g~�z#Aټ3��c6b�s{���M�;��A����i�o}�<��+πT5�xb�b��J�@M~�=���ݞ�=y�_va���C^����G�q�;�V�ϳoK��;ZN鮆��p�$�y�rv�1��z�	��1�wNXs�dSfeE�Pm}b�~�(G�	�?O�C��Ig�%�3]���?u��,��Ỉ)xo�o�t��ݼ�.K�~�[�A�:�Y1{]G,7����4�W72�2��5cCyD�k��]��q@�(V�wr<V`i���|/^�wx��U�ۄw��r�:���0�o��&h@�+W(�ׇ�����s��	��Y�I9���Η����v>�ז��U�jg�#ʁ��xI���&Y���$�v`ƹ��t9ﳠ8�y��= �H��%�y��^$�;�DJI�{�=�+�/k��[^��v՚c�ƅ1g�}�]���������a�z��`�	�f��6�v��B ��Yߩ�̷�XRWz��m��鬄���ے�0Wp�o!���-�X����i��w=���>��g1'Nނn��w3��D�lЮ�����f��0����sGL=�ۜs���Y�w@q	�n��GF߮3�{h�\������}�^�]��g�!S�ޮ�ʾ��S�Y��>�:f��H�տ�v��T|�����y��E�Đ�~^k�����v���q���<�1��7��GK�3uk�l%�i�K�.�䮻�}�̝ʬz3�x��<���I�wr�j�G+��a���kS%��}��f��)m��WWб9K:�k�MKØ�]Y��uZ7*A����0�_Sv#s�]���fgY���a}�k��v_1�f<p��YȫS2tᔩ����G�B�fu�&e�6;�W�̬��ۧɥ�|�-����#��.�n9�ώ��=sDVj�'�s�4^Kz����Ɨ��ۇ��#���ӂ�����ϡ��p�cBsY�Viw�<{����H�Pgv>;�y����7��V+��O�]I�=;wP���.�����{!�G��׼$�+�����P�FV�֮ݿ�*���ݙ��qx���Ɠ<Zc�v!I;�*�}���������K�^UO���|�����gҩq�s#Y�6v��w"#�C�v�q9�zr�ۘ1�M3���an5�:��w�O`�Lsf��@}�ev��S��߸v����C�P��W8[���g|���ek,N��WV߃�{»yҥ�����ҧ.���w�B����(�h͝G���S��g��^:��*׀�?3�� ���ަ�\`SN�mbVWoӘ�Q�S�DR�ʊ�'C}�T�?������֊� <_��5����9�-��؄�A�
�n���==�{/EX���=m�&�q���V�̠/t�r�]�3�虱A��ڳ�����0&���9���?�L��7{�|�)ݝ�Gv\T�{X-jӮ��]�W���R�:ћLf9s�Sb���Am����#������>�Z�g�V���Vy	�-uԫ�
����,G	���� o�{<NNQ왓�-��^�}�f/�Nx�����p]"^��VX�#o��,�ߨL�?9�O<�K�_y��5e\����/S�fN]M��m���Xc��x7A�'�����r��{�4�~���WXp{�{I޵�ad����Os�K�n�Վk��ت/�O_Vn��#Ʀ�RUa_z,�i=����}�M�Y�ơ�ٍ����'_�o����=`>�O�9!λCd���{ه�ڬ��Y`{7���߫���{��G��{���=[k���Z��mF�⛉{<�S�c=�՗��$�{�#Wv�z�#<����]����Y�~�=��S��1M	��>�N�Y�ǚ��O���䯓��[���V�ÖP'����-�b���������x�a;0�@�+]�t�^�]ٞ�{���䎔�K�z��o�JmT��Kե�.��3Ϭ�]�u_���a�Gg#��ېV��'��k�7Ϟ�{37]�iq�B@u�L_K�T(r��̎�ёw���  �.Y�����b��ۓ�k�tk�yy��}��0"�(Ww�X�iS�~ڷ�����{��\>�4r�k��r�wWN�Zyou*G7��\��z��'](yUn{藶�g�d=���>.�M2F`�ڼ�0ISO������!����/�Ѓ��}��e�#�]�w��9ۧ��=�����7}�ng ��$��"*p�4��[~���3�O�̈Cۛ�sݤ�X<���X��>�b�x&�H<r�n��3��g'$.Ѿ���M��������C_�ȣ�G����l��W�I�7b�^Y�������w�>�-'j{��˪����:�]�^^��&u�Ӈ��2�^R.���Z^���V#��I����K��{�}O�܈'o��cf�%���[�f3/tA�q9�1���f9շ��5o=S�D�e�r�|�/P)w�/D�K�	��Y�0������S���9l�h�tΡ���vC���I_o���i`��D��z.���ofvJ܅�걝I-@U��Ѿ#^껗�yV&��i�š�J���C>���L=݂�3.;;*�Iy��aCNg}������� ^���<�6�e��	9�����=�=�M����x�粼��j�u������w�ޞ��zw����.�c!��پt��4W׺xe�:�k�h�٘����Ċ8ĝ�lt�ۊ���F]M�w�@"��inޑ��n�����q!���{�q�������+��^�ׯtA��o{��Ԉ�|)�Է�#�q��>�|n%^��֊��{�^�zZ�������ϰS��_A�N��`<�{w֛�W����Wa���Ǭ�a��W����X<�8��X>�	jU~�~R�m��7�0n��9��F��h��Sa��/+���6���.��L����k5x��v+�ӝcޤ�z�>~7w����w�-1.���0d,���+����{�W�_��V�Q���<�� �8�޼��D=戗׼��a#�r�u�����Һ6�����M�u�k�Ǩ{o0zdw�N��|fpZ��`�d��gE�}X��v�K�+oj.;�:�����gL��K�>w1q{Ζ����z�zޙ��>��g)�[���f��n@W���	e_x��Gxz�okɾi��ԕ���i1/�h��
��NePn�Q�L�'>�+D�;^� ��Ɵb�=���~X\�^tqÑ�E����&�4�Ɵe�k�»#y4��
l{;����	!��bw�H��c	��rsA���+6�� �=S{�^j��S�O+hث��;��6�P���I�q�����&��<�b."��(Z��w����b��m��ƮC=�~��cǧ5�fi��q�mU��}�r��Of��<fs>
vg��:�n)�s@�fHn�v��t�LlxE�&�p�U�J����7���y�v�\���Ko�,�7wm�臧mf?q݊�̻� ��KSӞ=}�#��-�>wܱ� =;7��7ٰö�ǟI]���:�q��}���r��qM{��{f׼j����H[���p�)�ڰ���v�����L\h[_ᕵV�qWE'U��8�������D{"٩;q�Zzfg$f�bQz����}��\��N��չ�Ì�(�N���V�[����>�7�`���]1���6*�k����tZ�TYu�>��b��s�1�yy�[t#���`=O�z���W_�]����]lv��<��t9�TދGe�����A����HU�<xWw�ʗdnE�'�˯k��mf���|��x3w$߰xzu���`�y/X�y*�%����mޞ>�n�3�h^at���j�w��}�n|4q���cʳ�q{Γ�==�XL�U�M��\��|}]�V�����o�~�#�����_B'��/Q���i���w��t4#~���#Q�{'�簛���'%��6X���ڄ9��r�-Uf���G[3?v�z[�-������C^{�~^e�y�}�ϱ�+��o�4��^ۥ�w�Q�Y<����<������s_w���RSU�*�5���������{ɍ��r�τ�C�Ю�K�9�uA�{Ξ���Qgb�F3ݗ���S&��V��ٹ�N�pݟ\�o3`�A;7�j��fyi��kYɕB�T�z��I֓��F�l6:�ۦ���T�+J��ZD\���6���h}|�k�󴲬q�׺�����t]�=����ƕuG�7ygX����Ɔ;c��uid�\ְL;v���s�R ��C���E����u�h�� �#C���=�9����}��&ۋ��NO��w��zvZ����e�y�S��g�5�ʯ^��u�Ǐ�=��3�S���̬�i/�VnCJw�o�T��	4'��Mo��u�Eۢo��[l���f(�ԑ]����Opo��{B�󷹒q�[z���=u'H38�g1�0F�<����le�0�!��9����ϭ�*�36���'����ә��.�q��w,���7UU�'ѳr$1х��y�2�D�F�ʤ��f��xVע�c�N��kQ�����i��H�$t�7�Η�k�7��mu���x�q�0�H��D��^bFN�C����v�d5���k�z��;Wq�Qyuݾª�->t����@���GH�l�;��l5�8,a�ٜ����w�z�N��k=�[�{S��ׯ���w=�X����^�6
"���j��e�/!���y�����R�ݨ/k��i`��u5^WQz�VX��Ъ�T�����M]��ֽ|b�ֱ��/,G�Ӛ�%��
�ɤ܆]�&���;{��a�(AV{��KLi;M�cz����9G����3WBA�s7S%Nz��a��Ǉ�CW9��>�1��Ϙ����y�=������"t�����jJ�tn}"DƬg�\��g޳˨i����=h߸���m엻��?q�zc�&m�����������E����y~f�Ou���;���P��Ϸn�鮫�ټ�7Ѡb��͌��Z�.Z�{K�w�v8���j���=8�p��zG��8~�"��ܔ����[kkTݬ�>� 9����Z���]�z{k�OD:=��\��׺� oi���\�JB��"yf��/���Dc ������LI����OsQ�%��J�J��� �T�Ӟ~�jF���Xs�<���z����[�ﷳ��yoݹQv����<x�ʘ��?wL���\�7�m�Wk\�L{�Ct��t=�$�l�,5jÖ���hѣGA��||�8�y�3�,0�1��A����d���2����z4()�����i�]u�e� �����z�mX���x����1:ƮT�evv��7�+����K5��cWWsV'֑ ���[<�l�4]���X�{�+���ݢl�	�&�Tv
y϶��,ܓ`�T=��z��_Gf�d��$b��-���z��B�Kgn�ɴ�,��9�)��ڳ�E�[�Pz����)��8y�Q:vt]4��)مe��:e]�Z�wX�W}��5�X���ut�0*����)G{�8s
��8Qp��j_�`��߸���Wʳ�A3��ظu�Y�]��xk�[���.<��CzK��1fi�8�R�g_s:�^����fN�ۇ� ��}��M�-�M��(U���B��yk��)�w�iT�>�x6΍��0Y�޺��8�\R���"X(̒Ž���F춲�u�� ���	z������YT����MڊeM��K�o�CFR�d.#��D�ȩ��]�;�~�E]_0���nS��L��3�7nV�;{�.ݣc)cunm��DoW�h�;@f�5��:rI�[7�PCr�NKG��d�*bˣ��e�僴�Z*>�;%qŶ8f*���r|�mAYIN�^ʗm�� Zh�G�ZB�{5vt��k�OvU��{t�C�ne�:����ilՏL�`E�J��oV�n*1�V���A�0:�=Xx�'ƙ�3y�Kyv�7�Sm�<�k�8L���"�f�����!�l�u��k�Hj��(uR;x�N)6 �h��<�b���K�SY�'g:�ax��{3w1@6����\جdΗ�X�K��E�<Ѭe.��=&����9s�d���H�a��S�Z���1a냚¥"^�!q���:�v٘@�1(��U��@�t��"�:��s���y�X��	���;���{��4M��8�^�\�h����m�������{7��[�
�W��c6���|��O2�f�ᠱYG���V#o���9�A�Z�����yK<�7"��!y�qK�\�-��첂�(<���s):�3�^�o���B��d�wJjJ,cH�5�r5;:�:���o&	���BĆ��;��G�hꗵ�3��3lK?����y���M*��nvD�aЫ������e��b������c�u+�1�$zRP�[IXL૧�u9}	6zm��R�WMu��1���7jwn��ޠ���vN����o9���4�![�����n���}K�E�@F�sZȶ�-�E��-��|0���l�^丈�z�Mhol�G��[�wR�^�;7Y��n���s�d�򬤍t�Թa�:E�36�h"�ז��m�&(�*8�Z'N�vި4���05�Y��9\�S��ٴ�e�֔A+��up�} W��6��z�С�o��>o<���;��g�"�����tkM4y؈j�m�WF�`�V�:�)��=v�Wm5�*�)*�1i���*�`�2UkTV�UZ�muN���b���F���Og1������F����
jݵ�mF�v6�q8�w�=�F&��Ƃ6;c��趨���wv^�`���;[�����v�$��݃qv֞�<�w�m�w��Ń��9#F&���n�����ww'�v�k_�j1N;�<��"�ٻp`�����f7j�&#�۪;�~#yyآ-�kUۮ��u�y�D]t<Th>#����]��������bKEѣl]c15���O��>u��#ˮI�T�E�A���|Xm�>V�Gj.�;��ʎ����pQtmh�<��X��������m��"��;�n���Ƶ4n�=�U���AW]�c[i�b�b;<�*�V�E�<F+qtW�o<N��-8班�A���l�-�FԖ���b���&�V*�]�z�U�������&#b�v{��Yѩ��\ch���-Ѫ9�Z�)�[��A�QET��������[%:����UG_n���;�}����g�0��6NOFB��� ;�&P@n$�;�[�g6�p�63vJ<׃^o3xT��<|��v3[�D���9��C��������E)MRf/A�v��FuA@`���_�7>�;��Dj-���40�1l�gs(;wq�v�����8��6�=7@:z�Y0��I�u^tL�]��%��aB`���W�"={�O��UDH��I��k��-����.����Cg�D�2�WQ��I�ߊ��'P�k����}�V��uF75�vzC2#�8_q�	�)ط�z�_�?��=�hS�j���M��sC�>^��`��R
y5 ��J�l��L�ګ�]���ɫ�v�1mY׾K(����xi}�Ƚy�$2�Q�#�>�v%�gK�\k]I�>bcg�+��o*e�ϟ*g���9�178N�fò���<��:i������IYT�K�p/Z#,���<#�O�:<���)����UՓl5������^@P��I6���(3ư�Z|����6q�s������57��I�p������E��?f��=���[uuLkQ}P��|rO�p�(11[�H��t��q�] <��%[�h�������Ƙ��JOYaѤ�X�%p!;ʽǙ������NlO�ϋ�[��#B�5[�KW��Y���Qf�v�6��녨��@��~U�Rju����ݼ�)I�� '��Z�����͗y� �*Щ�:���j�v��wjL����z� k��3[Ǹi}�P�v�m�9^���w�����[ �?s伧�~>�#�Uc��%��.1��宝�u4��Ћ�z �W�����|}C/�i��ly�3��7��/:��9]O=.p�N�ev�q��3{{��h�&`b������>��,�:�����i�d^z���f�{�$�G�1h�3b��q�՞s��8�ȶ�Kd?T��z�1m�w-F=`ŵ�:h�T� �C��^����
�C�n|+��]{#|��������N��g�eA�'�%/L���e��=�ؕ�6|7�
��(!}���ǝVP=Q��������&�ON�A��3��5E�������x!�`�Y;�OK9�I�?�E:�Վ�q��]�U ����G��uZ�7����������+Τ�q�m\�ԣ#�o��y��5�-�N�7s�u���Y¸p~�13oB�g�9,1���bG���&a�l�'�sP��p�H�:��OZ�'�9."^z˾�D�xd�S�ڛaW�+���e�G"���%��[a�˺wb���ǧcǻ����ν�M鸧#N.��(�s����J�Z���*ذK�7��rSŽ'�`���T�(��G�T��)�e���VԿy^���?lE���Hc�>�l+.�뮈Œ�쫾��Q���ld�����N�H��ȯ��"vŪTm�ɼ�lҺ���y��ꮵ��~QZ����x�Ƈ�z|��ќS.u�)�|0�?���`;�.��4Da[{w4����m)dC�|���V>[����(x[8<<�k��'�m���j��My����P-�dW�:Ҭ�׷}���Ȇb���`\E�!�F��I��a�:�̝86�bwsV��{̨?q���W�/�V�G|��<2�)`ϣL:5|>��a�{�܌���oʽ��LD�K�rT�q�LS���2�~�9����gB&�*����>N��`�a����B�N:���T/�qBͪ�,�� �5���@�g�;�Y�Hv.�1�6��M^o*艉�R֥,<*ex|Ǯ�ܾ�Y���A��m��>5�q�mx}E�ӋH���0A�{��»^��I`^@��%�3HA�wn�8*)��m�ĭ��⤽�Q�qۇ5:�}��pBf$}��`:j8�>����/(451
��R���j޿���O>.�s=U�����-��GՏA���?	TzS#�yP��;k�ё%�p��vO�&��#~��T�t�Ho���5g��ٽ�(z{tL�k"%j�v�vd����:�.0����ض;����A{Bt���T�$,�j�7���ν�&_����#�O��\nN�F��j����0Ν;U:
�z����J���T�sS���ǈ�N�ڙ�>Ym���觏�_�1>�q��{�qL�
�MNnY�R�g�4"=��,"eN���[�9T�zsuV�ݣ|�v��-�,��b!F��N�~�m�8�$ [F)�>�}u>����{U��)���/6�o�-8���C��(��{���s��BE�c��6���hr&�M����v�5���.��{��l�y�R.�е�!ٯ��
��u����[=�Bh�YA4�Y^���f_�뭋���\c���(ύ�`�$�����Uc�f<���?oK��Y9��Át�@4��cs{A��G��N˯��4h�͑�P`O���� m^�]��������
;e�"�4�L]ffGc�����<Í��wf̱���SlR̬�j�FE�.��}h�ϥC	���m�v��Q���z:;����=!���%ؼ7��-݁*����u��M��W�ŉ���|#�m��'r*�2{dc)�`��u��ZF*��7�ڇT��"��^����R���R�=�I�DU@5�.}��+�/0W�?B�Y�M!��Տ,��?���/B(�\];�돝H��@�G�֥�5\
�<�������h�>����8��n$�������Kc�.��~i�F��κ䋬L��<�gk6�UJ�sy�=�;��]Gn%�J�cUs{kRs��!��T��Z�̷ʹ�)d��9�n��
�՛\�ȱr=�G8fn�ũ�|wp\o�냾��a DB`7��[df�[�ƣKI�_�
�����%Cfl! - a.�C�3oHC7r�(~]�*�c���X��[�,�Xs���
#k�l����Y�h2RY�����ގU8��3�v�71�9��!�6�/��l/x�̇Qn��m��\��*�u��#Z�F�:��=�� Q�k����~�`��4�~HT?/
��'����L��׸�Z�����BF������|t�4Q�����w���cG���^�"��h.�z�I[E�~���?1��2��y2j����F�����9.��k�"E�*@����AְJ��u��V%3��$��%�l�KM��Q=��sFe�ܵ�vԡ�(,�5<�Y�s;��V��F��;������x�Z�S��Nό-�E�.K�u_�&�m�Mzw*3�Q|�3p����s�X�/�Xk�p���/���1ͮ�-��{��8�S\?��F��z��ݟ�0�\�N������%�bY2٩O�����	Bj#r`4�`9�1�|>�ΠFRy}��n!�˯���ڽzȭ�WE�5�{q��wx�i�ʝoR�S��$��l��Yk#Ž�&z)YW���7���5��&�q�]ς�30]5ς�L3�h��e\˛�����_r͒e�������m����p�s�s�m����꫑л@g�@��>��Nes���{�_:���I�ǱH��Nc݄�FF��F���K�?m���6�����wւ��w#�E�ou��bUr������,�a�{)N��D4B��i�e̟q���!`��x��go�\�I_su�~J�d�7���,��1�.�U(E��P6j��q\��<�zz$�1u�$��r���,�\�-�z�:�osR�?��(�F6W�[`���w�3�i�ρ���П�z�Os8i�om���}�1��ڳr�C��ɫ��	���<3��E�TNWڰ�6@�C@u�aG�x�2��t�/֢��n�]k�+"�ЎR*�T�m�S�~�j=�&k�����v���,� *��-�z�n���ꒆ����B\,QX��B��<�N�(ȶ"�H|�UZ�	���p:�)ʗgR��Z�o�K< J�o���ϧ�������倗�F܎�1�zd��K��§-�F��7YV�2�$�d�ꂠiG�P�_��Ǟ 0{{v����:]|=7���$��¶l�.�J;��F��'�7v��5U���]�\U+���s�u��G%ⳆP���ʁU<�#!��1���o�<w��ϕr�b��X�û�WbG:�*�r��ݽ.�B���k#�X����ۂ��ky���W�*����0lf��w�Z�l#��1l��s�;�*'L���Mh��J���e��s�L����@y�^�S�dw�^#�����wDj�y��L9��A�1�S��s=��/l������km#;_GM��I���E��f�9�O�2�ۼ4�C㚈���@�G�ጻ�Ů����+��˥�g�B�/�A\Qsim
�gKhn^xk��C��Mwk���-�l���- ���L�5�g%h��X�o&��v���;�9/�ȼ���Lt��:Z��%T���!�"=�����௢O�11|ު�-�c���d�T���fr-�Қ���4��։�x�r��9[C���@��;'�b�@��L�8���ؖx��X$�ԩ|���Φx��'�c���l�Y�`�����r�oO�0�˞��w�ǅq�ܤ[C��x`c"�Cώw[~�Ǚ���~.8��װÄ�������[Шf�|���Gh��OÛ����Ys�Az�s��\�qf���4Y��jgƭ0���2*�_�{��#����`��ױ��t��^{�L?@Ql�C�]Dn?�t�6}ipQ$�+c�`Wt�յn�7Ֆ����-M}]Ҷ���n����G��x��މ����˸��,�;H,
�I��ۆ�û�K0NTBf���O_$֝�Y��59e�u�����vx��Z��Y�j��^�����\�_݃�}�
Y�����1��-),.b����sb�EN�Mq�=/3�ҍ��߃�-�S+Y�Ҡ���,|��)�����t���f��+ǽ��l{��ޒ���}���+�����Pt_W�4�D��D�E�'����s��w.��xࣝ��~X�H�!��G��ʀ�H�(���z�� �X-�B/t:��OEf�ݖz��UsQ�C���s=q�l�
�MA��;��M�Ǚ���M�"��H�Wϸy�0��u��#L(�̔&#us'����\D�T��f����ok+�Mp/��%n�fn��g.TH�dC�|��5�/��jZE��{Jn�&m�j�w��('yF�Y� d��憩<fY��"�
��ˉ�1}f~�(�T������K
���jZ�3�I��Z�~�)�q��7�b��QF~�	���;���U�α?�ռ�cZ�0����tP�p ��Ӛ��[4_��G�_7�qw�=�(��_���&�&xf=﫾�x�$�u�f����������CD4����)>��1T�̉�����{��4D�����˰��>���;y�R��׹��|0��8�q�3u�pvq���̑Eݧ��%v}S�����C���n��=���\�NrA�Z�R�hs���:#���U2�8yV1ʊ`S��O�y<�[4}��T4�7���qЃ�k�r{;�<��H���%:aa.�,N���pm�GT�d=x��y�!�2q_���kY�Q]"�Јnw(�PX�1���c{��c�\��IW5���m;:+o�����^m�e��\Ёvt�]y�<g�ϭ^����ʽ���z���	�+���8����Ҙ�y5�-�9�=�7���iq�L��#Lo��c����	,odEL���^/��H�؉����J��$�dq�@�B�	��d(->�.\l�@o[BQ�tX���2����@u��:���7$�YS9*Y.�E9��[r���5r���-r�h`���k7����e�,n�\߭$�2[�{�Y`�.��w�[w�m>_��=xY2(I���(��t$�4�����uW5��u�w"[�`�5p�;/^�lp��l05��ˈ%߼k���\Nz�����^�ј��vr���{�����?�Z��%d��Tn;6���݆������ ��g��-�n�*�Yx$�%Ws(��]ĝ�p���I�c4��u��fWj�����ҾХ�V�{�+7K�]H�p��l=�G�{�ٺ믫��	� ֯�-S�;h�R6��mt�K#�6�XK�$&��n㺍�J�#�W��^�h�[����j�U��B�|z�.���6Hg���$�W躸�;`m׹�ٓ0&#s{�B�7"���Y�9�dqn@��~�]&k���*'L����K6#�s���2�UX�|��n��r�S���\��k�+&�/˶���j���&�jz�t�9�<�E?Y�:��v9�m��k%��*��2L���r�=����n��љ��P�0)&��M6do{3#����ŸI�"��l����V!��߬��>�����櫍d&���}H�O�F�w��X�W��y��j��S�H�="��p���S�׊�O�P��
=
�9m�U���{��j~b�?{��fn���P+5��� ���2"�z�"����a���R5t۩U�o�f���\v��6�ya�@���X��rj�����n���kG�����g^��%�S���I �(���&mΨdB.�{F�61���F8�D`��c�%w�,�����ɉ��i���Ε"�����=��О���r�E��/e�ݶ}��� ����0��fNZ�nٳV���^�rR�})����k�f,hmp�bV6��7���^-����\�Rf��y��ґ�(q� �i݌�GY��X�R���Y�Xz���������R�[}pn��i=`6�C8�# �j���AEf�n
����G[�Y�5W<>�P mЮXW���޵1����l1���v�����v�q̽���T���NN�Aµ	׉m��k>WC8wʹT��f�k8�n6�'c�(�yޛ���z��,l�6��4����n��y\�N(cC��mo1�H�����f����f�K�=�I�Z׺�R�4��th�J�bׇ��E�/Ǘ�ZG&`ko'K����3Z,u�6eǘ%c�/��ʖ=iY3����g���T�6�3~�G�Lsh��������C���6�;3��_ �-^�{k`��n��룆�4Y��*uw8{���WsWR��eA��$ka�,-����y����[�9Ez��	m��M�8,�J�-�2�=�;w;ķl�}��N���EN���Ё�c��p�FV98��D�ˈt\�]W�
���^�Y|�k��+��c<n�M���KOT�R�r��wۇ��ݽ�E��7P�ѝ�ګ�A$�Ң�X�pn�L� �����f��NW�m=�dQ!	�v�m�K�Ub'��6)ny��SqR`�����V���uۙ�]���t�'H���y���]��a^KMw;:���*�'e�lt��z_�iw������C��ݵ�޻�w����h��w$��%����q�X��ԫ�W��߁���Yi���.�����7;��@�c���q�2SeU�d�PP���ڏ悷p�
<��Q�w��,����PU��wv��!e��0AE���r�ؗV�[�`'Ɔu��}�w���(���S̻,I&�V�4ȶ�u[ ҝoG{M�:Wm�a��K�[�uo
��=j�M�6��:��s1D��p�2�o8�bC���-�]ܒ�����Q}]�]��]ƍx�Է�mv�K��+`�wr�i�b�����*�X3��B08���Y����i��&]��Zʷ�n�"�w�����0.�R���N�F}| rT��ګ����^,s�ǩ��v%F�o_y��U��]|�
�Z9��ލ��S�̃��e��_��>����~�j���������!a�[o
�Q��0��ٜ��n�D������M2��s�b��mK���Xi*�k4ȹ��n�N+fHW�#6�����Q�ʷS)[�R"��s��+G!u��[o{�sF�3j`�wR0��Y�i��1TK�E���6���9e�yY�c�&5��g��ٔ
�C��b�@70RRi�������JX�+�G}�iW�Fq��uZˣjۢ��V�̎y�����̨6�q�)�Y��;���Y�KNpwRV�`T��Wǡ�z�$w����+4J[E\�i���2k�=���28XT�n���n\�^��Iܺy0�	��%ۺY��+6���O� Z赋�wW~�ޡ��@������ݖ-�^q�uv��E]ۢ�ŷmWX�ET݃T�AE�E�Uѳ��b��&��v������ԕN؈;m����Q]v��u�����c5Ѫ:0E���D���j�7X��mt`�8��4�w��z"�ƌEb��9����vַ�Qh��j��������طv�Vu����Bq�uD����8����ͺ��RQTxX�\u�"M'[�Z+��lUkS���l�9�TͬST�E�tV��֊���:iֵ��4��Zpi-�#�آ�3E��Q�����RPSM�2TIUZ�m��:�qk�TP��Un�ɢ��R�Q��-�j)h�5��]h�X��DAV�S�!l�d��棻5v눤յc�h��Z\Ѷ�(�M�Ch�v�l�(���M��IM�iW�Yg��h|�l�)�'N��3���g�S_�C&.�� G�e�][�������r�U�5ܥ�CY}+D곝��Q裼�̬���޴�b���4�.�Zd�H��%�L2YI������?hT~|�+6o��&���߿�p�A����BPI�~Ϗ�$Λ�t��=<w�1����m��y�=yfϢ�5�Xa�����_�ˮ@gf�c{�q��/�1J����t!�[i�]ި�3���(�Ƶ��UV�C����q�&�W�s\��&]@6_̈A�B^C�퀹l��G���V:<����cl��V���UWQz-�G����]5��"�q�u�P4���j�5�:��ݻ?~�PDxp�q)�y�mfc�}7��;����A�YqD��N�����k�\[r}�:ɥ]�&�^^�Fb�8^�&&v� ⒄ͦ��+~� �s�E�/��B�Po��;�ίاzd��������3��f�K�
|׆*Z�{2�������dKr5͒g��P�'�ȣ�!W���b�v4�reR*�@Y,
���s�Gj��~΄C��/�Ȝ��c
j�;9��~��!���=ؑ�jO����8F��ݟ��扻�L����1b�yw̿��S:���s�c���V�wD���)ǭ�[�.��DE�#ݿc����&q�嚵N�m�t�-�L�4-0%�͌��ê���2��9]ϐ�:�PC�*�y�{:x��Lbpher�T��Y�Ǝ�)5'
���oY�hEX3e��AȔ���e��M.)�Α�Z��uf�`��������Ҳ��\�47��8PHa�7��C����Շ�|< 6�Gf�A���>]>D���^YyCQ��{lw��0�|xb���15솓 �Ƙ��tZ��E ̽��*{鄝XOǟ��g+9coƦ�"�?�PR�0�����0I=��NS��K0/KfY��{=LGzSe�^�yׇ_�=10�����8���ʯ�yت=�8O�P��m�0"��σ�TP��<�ڮae,�y��N�ϭ���fB����j�>�@8�:��KP�2��������qT�L�7o�]:���H}���*k�[A���T�Z�Ӑ kߊ��A��52��]l�t�|m�4z��Ńa�LS^e��n�̥��:��Kʪ�Z�Ƃ�<]�qg�A��3S*����e�u�k1^!K{}f��
|'4�_�֋/���؟T�Q4%��z���v��:2"|'g��y�f���z�0��~��Ng��=��(�]���1G� �_r�G�=I}����ˑo2��fg��W,���?��t�Md�}�}q�2-�_��?l!���$9�_��g~��l+s�g�+�B
�8�	���7�W1�Vl#�����|(��(=T�SB�*=x�؃�X��cU��5�ꥇE-3����q���a������v�z��a�*(
����k��S�Wr�W
�/�$Ǝv�p�2�RޣG���X$�y`�y�L���������Y$��W��DKd�Ɗh��*�+�+Ȱt��ŉW��<������"K�`�k��y�=W�C���;=���2L�(��*FO����K�j�UV��USsX�!6�ŕ�QT��\�P�ߩ[�O��©Օ�d7���)uyW�Z��`]g��wq-�t*��k$����ıʾ���y�qr�60��`��1б(�����e�� uT]�DC�`�[�6y�tAevUSw9�Sm�.m�r�� [�ajiпv��#���!o�a��{�V0�:˨?B�_�ħ,
�-�Ò�n��q����0�Ey�e�Ъg�-�v!�'Od��|;qC
/�&���DR��E>��P[�7���⢄kwX�eʊJ_Q�p�F�t�7�|����s��M�Û�.ޯY%�EUr}�S�V�Pj��jlk�5����^��*<x��j���^��}+�)I��Hnn*-l�-Aڒ�2��3�8&��j�%ƿ/x��bp��qrF�7����C��	���<X�ꪯ"t��y�yLleJ*�*j�f�}��.?�z�{�TU��-�~:���T��&�ŰyT�ɸk�yQv��c�yPYP��ɭ-r]��-V��Q���}�qƺɋ_|b�r
3�¨s�靀�������L(�=���&^ef�`�3����{� ;W.r�R��d[����}�*���%��ֵ H'~�9�|*�4 p��Q�|{�N���L�>��uϨ�������4��Gt�j����1�m���=̙�0���C���2�8�\���Y�:��wF��Ƹ�����b���<��.��%̷����;�="������Kj�M�>�0�"/(�2<XB���Z��AS6���v��r���t۶0d�B'�Yյ�7M!L�8x���+�'C��1�|Po���*�X=�2}��U��<.��P����f�֩��d&�}j;�X��ؘ2�tY�4N�aibF+\�M/��p��Vc�F�'�W�F5���|�eO��i��o���z��<h��K�h��d��R��޺�;73�<���Z1^hE�Luw'Z/�8TC�#�.�]�ǳ�����-�r��I�"���1OM_Z�r�A�%���Fl�M�<�m�_�|��ƢE���F�=�^���W��ůd���ȏ]��*&�}-�_dpe#�u�/
w\����5�u�$���䢷��&��d� Z�f[m�*��:F̡^£����轻2�����v]�W��@���,ȇ���;{��F�ʅ���6T�|=�~�\�73sS!�\�Éff\�Z�:�功>�ղ^wqa�������ֳ�|w���������� C��
1� ����S��eЋ�������y]c�TE�x�eW��9M�A�gj/'��ΚL}}����+�n�ٖ��\�v#W=��J"�����KP�R��ܪ�U�ץ2�q���VP�!�3qL��~�c=�D���!���
�$��ǹt?>��GlR9�����p�/�6��◮�O�2]�;��6��L��z�H��7tж�����О�F|�O�-¢sNF��;Ez�;Q�s.�^u;��,��熂辁G�u�h�x]�����)�t��3g�t	����l~�{;QIs�k;��j�D�G3�(,Zv�zO>��C��+\j��)��-���"R��:�UU�㚸Mq8 L��*��(�1}���ՁڼM��/�s�����������4��Ǣ�}��٩�H���P��GM����_��ǝFHG�~Y�Ѩ��׫��w�ܫ���ּN��&������Y��;ꂢt��s�,��8ܾ5�=���8rR��������hh�����|F��ۺ �T��Ο3���N��#V�P�ݍIw6z�y븬dr{��]=#)k�`uxe�WSg��P9ê�{�$�ŵԳ��n��nJ�U%�S�xb���>���k��; C7�>ީ���ڝ�j]4�rv^���q\�;m��o�o��߇�~y|ߟ?��H�B R����f����oz'h���znN�K�8��w�^)e�_������K^�d�~�%͍���w��_{�G�7*ۗ.��ǤS���xG[��S	:�k�\��*���br�ʐ��[ �X�h���"�u"��6�ME��2~���|��J�ԹK.7������u�S��n��SL�9\���[�.��a>��mtU�����-���]h�O�*@uU
�8�m�fei�c���*|���������F�\�60����ba����Tf��;v^:"mT�A�%Hf���c�_�T=Ǳ��e߲�}*����(�K������e�j�B_C.xǒ��)�|�@v�L(S�S��L��5��+O�P����ݿ9�%H�Y;�:�璜d��ez\BcNqy��#�<��0X_�ӌqV�(�e�Ѭ��h��xِ�>�O�bA��g(��壑:x`�hI͊��H�4*��R�x��><�wa�Q[�����>US��,$\�(� w�
��x@�x�L�g����u�
Zn5��K�
�r.��L&aRj�mZ˭3^-�а�ܹjP5и	���D�gZ�\pjФ:m��WJ�����վ����f�����q�;Eͷbw9�u��:�;!*�d�.����a�w@���+��߻|<�
�qp�,�|-����*;�$=h�UU ~�"�PR!H�J��7�q�w��_��R�"�G3�yUEG�ZGƂ�6���mx�C�f��¤l��z<0U��Ó#a��/.߇	Oj���f�q~i}k�!�L�f2!��� o���Ҡ�L.��;:�g3O�kGT[�K��a X{ezg[@�u���`go֤��`�Xȃ�>!�)O���5�MP��y�޼T����
bk��*��x�}{j�f��%ߟ@w!�G#�QL���97�k�V�z��x��ɨ�B�%��>��tab.��W�J����ݪik�,a��B�5Sg�g�|֓�3(���zn/q�w$�;/5P�O�!����޽.9�|*f���)]���V�a��N]��y<7f�M	\�Ȼ��8�L�W�r"�<$�ر'�� t��pT���Q�d�s�����LԽ��r�q���<R=����6�.-��Gb����p��^���6�l�Q�έ>��M�83L�W�W�O��,=��s��6�K2��S,����e�c�.�:��G5N�M���Բ&�ۨL˞�9���ҩ`^�Lsn��E�ǖ?i�_3_��'V�\��մ��݅r��J���tE�b.����f�n��=[���p�*�+`�BZ�:������͇C���_p�^�=��!ލK�nr�!�&�g�.Co�w�]�-�x�w��ں+�×Hl�9��:�j�NH�&�A{;?�����(	�P(�
(~�_�Ͽ�����]	G�C1b��	X��$hB>�u�M޾-!���mC��%=��(�3F�]��\½�u�����g�-���1�8���
��	&tW�<����#ү���{�B�=����^K����]+6�F���p��Nq�荂���5cEw�$鍈�5�T��O�I~�!���cY���=Љgz��X��$�i@�Q��f[��&�$c��6���1F�G�`����-x������[�Cڌ�I��,�V���Ig˩�4ߵUkR-r�h2�����u[�0U��s����kJ��X�^DwH֮��O��3����󀜚����w,�zR�TJ\2�+�澖Ɇ<q�,���&!�B�}��a}7��Mx3�9�=��w��,)����]ӹ����}�ӏ�?��"�v6��1�zW��x!�������#�TDS?]��٧u�zm���"�Lߌ���N���o�	��M,������y��t���|6%_e�#��$&8����SiV���O#���W�$T>�o���Oȃ�#dc	�|Үx�\}\-��Qu�7� w;QP�b)�̥����-
���������Y{kskse����$:�.�ҏ�mJ�7����,yc��d�0�@>w��:O��޺���qs�m;͙��L�X3�^e� � <��B� �"�  �H��}�Sg���'e�9��_jD�KĆ�a�ݙ�/o�M�S��z��y�偦���he��izj�L��4M��'�~%қ:w5�"4���^�"��`g��Q��<=��b�)p�����]���P]MVe���v�]^D�����I�^N	��Z`�$V�P·��\����RuϞ��OݪE6^�E����C$���׹���8;�b/���to�|~x��;�F�l�	�k�Lr�b�K���q��{�7L�=r�۶�<���Ei��Ǫ._���e ��D���j�πu��Gz=o�+ԝa��<8�	���.�x�؊/����>V��٫���psf����c>��$s��~�˒���"�2ť�E�j�$�L��P_�q�9 ��nv�}a�!��2Yv��N��Q��fݡ�5�R��H����"��|g��_�XL�~������*'4�8��㖀C}5����"=����\��\��ؾz�q�T<�0�c��Y���9��^o���ne����@��5�@~�g�,L��x\Q��*�4�<dp&-8��oy��{�Ur��\'lJ�hr��0Wk}c6A����rW�Su��w�̓6p����V$I�{�2�]�U�"��E4�7i2�j�g�Y ����ۜ���aV<����D�tRBi�k��Rb�6�EYƘ�rJU����ߟ?�_�
A�@�0���7�����F�]M��_	�j��p5� pD���$k�&����7���T�m��ѧ6�M�j1�n��0�f��sB\�s˾���mvN�^��	��ݴ'r�	1tC�޳b�Bx�}ݎ@��'��"�O�w,W�|�gɫ�$��
��'6a[�i�#�FON�ui�E�hAFF��������	�ܟ0a��p�	� �9�]r�j�U�3�%��mI��!�s��E�'�b$��Q}�L5Y�(���F���|�$^��	=��QiٗSٺ�͇�J�Dl줏®�ʤ�J�j���&̈z��=��їj�}�g��rW�����Ÿ��Y�����{m�_DG�PX2A���L�^f~̩�֊c�]�0wQ,L<�Ʒ�ͦ#�6c�M�;�&�%X\]��aX�˩�Ӎ��:�%�3��,�#zxQ,��n�%�b�&�w0[��es��S�M�����Y�^h�l�:L*&� {C��W������͉'�	�P�M`�?�=/���"��s�O�Y����b,C�>>�&Ɇ��7f��ջf�Z���5�W�W�n�]�h9��=I醰-�]
��x��3Q��U�<X�I�r�ك��j��n�2Zm��*��A���ާ�M��Ҿ�l\_��T���e�Tj���[��ƦGO��u ��==x�|�ؔ%�_jW/U�n���bUi�6���|���[{&ݡ�P��)*�m�{Ĝ@g��]�*&kz���L�C�YPo;(����v{E�N��T�����4�j��Q��\���X�����2���)�%�_,�sWZ�`-�8���C��'m"7
�����R�5����pU�2�7:ヵkxjշ9V���ZS<;^�u��u�〜��M�k���ul�V�Մ��������U������k�9�eJ�(%�^gC�r����{mJ�
���p����y��ꊝw8�.��4F ���Y4_Q*��ʛ�oM��Wѽ�ӝ�Me���q�I�f�X�^�M�}2@�qs��N�u�Sr�w<=}f�zV�
���WG�d� ����t{�4��.���y2�{��Wv];���)2����\�e��5G� ��B���٠�3x�|̬��1�y����r죊�X�gV�dPʺ��q���h=�X<�4n�!BhԂ��`�=�A��:��Ţ��;&�uj'u��}�ӓBݥ�����8��K�����i.�Fԇf�:9��q'��`\�{��u���lBwuGB�zwjr�k��Fnw�K�K���p�Z �f��G�[�]{�wL�^�����`���s˨�&��>���}���+6�j��"}Q�7�;�� �}N�x���f� !p͒j�Ӌ9
"�k7l�'��r�H�z�u���wxYψog3@@�;�F�ʔ�T��ɪ�������u���uzTp�Y�Lz���-m�r�y {�1*�����*F�=˲6�%[*�0þ���\Y5��35��k�(��ku����u���Iʙ��=;�5I�{��e;�[X�^�ٗ-�6t�7��'t���օk������tG�I[7kn�Y��D��v,�6���S�b�\�����Q�{$��M��YA_� D��VN��5�H���"��bD����+5Ԕ6�:�.!��/��H�I̸������;���:h�i�8v�k���h2���x��d�lcB�v�\��$����'�������cq�:���ykNQu'4�.��y]nPB�ͫ��P�b��;�c@)�"
�Y���'}ٜܗ�z�%ًͫA��M#e�N��u\�w�V
��/%l6��y�,�0������;u�]��`���dڧϮ�-��h�Ә������}���w9�Mݨ�k�{i]�v}ʰ+Ů���g.��6�)7���)�rk��Ѱ���y8oQj�c]�5M�Gn����/xu_�Ԯ|��D��[�wn��SC6��j�@�g��SI@ݵIAK�S���""�%�SE�I�Dm��I��Ѡ�����n������
#X�����u�h�mj�jK�f���+��DKkQkDkE���'����f�z4m�+���ET�v�E&�j��(�F�);a��j�QUv8��:��Y���9�֤�cEEh:�{"#b�]��OQt�:�؈����"(&Z��ѩ����(��4[:j��튫�mQAш�k��&���"��kj�8�A֪��8��j
J���V��Ebz�v4�cU�l�5MQT���d����5���&&��)(&ֶ�`�*���(�������c�'E�Dک��3`��i�����������������Λ�(%S�{|;�Y\��Je�=���O�+��pu؝�p�q�u�4{����l<N�(?�UQ�(��B��
ji�<�#\�8�T��*���=c�{��=ن���O0X�~�^r�ğ_�_�)ws7��Y$�K-U�����,v}�üp.9=��UE�4aŚS�(��nR���'!����㹠��y�m�`�Q����� �д/���E����گ��w�4cH��4�&Hr4�e�m�>:[�0�,9k[N����x@��L�g�d7
��矝�Ic��������� ��ў-��cpi��8�Jf[��4�h�;0IQ��F�b'4֍�3٬�P�k�0�]űzJ�j�7�,q��|{*���]K]D��� o�OWs[%�5y�1�=����.���Uѱ��ַ;������~.)�
�MA��;�S����a'����W�T�t����T*k����:�߯2P�>�x�z�q,NdS.�͆'0�0�*X2M�����Z:})&6��U�#���3~��ps���xy��tiw�����?y=��~�ڥ?w�E׽p�|��E1����`�^L��p{ƾΠ��y����ťc�u���OfJ*C��ε8�_R�XXZͩO��*8b�g2���VY�����PJ�:���Cn�6�vT��m����|+?�c��ɜ�!_�nM����r��B���n���3�J����2��)�S.�J��4�f;��_;�A�� D) R�ox���ݼ��6ʱ��KD���|�jD>�1T�(�>4N	�`�+�2��~�@���֮\'P��Wؐ<�%P�Y��W���~��i�_�V����ڤ�FFl� ��w�_u-T��}�᙮-!����n�a�__�a�0Xf��e��^v�8���Y��(9Sy0�2�[,2DN-��ӱq���ߛU�3"T1��~�^�9�3�Nܛ�2�@R[�Um�Pa�0o��Z����m?l>�PZ?��}����F�}K��4�/�Hy�4���TS����I�a��}<Ffg��Zt?w������x� ������[�pq��~�o�!q��׽��{���=�մ����$��1�^
 �]�u#��ڣ��_����-ppD��	,o>эX^1廻�V��<E�n�X��o�H���KT����CAx:��l����UmG��U���s)]q,�O��衭qq&t���ѐ���ov&S��ܵ>f��*�jZ�ؿ���6mk/S�O��fߖ��t4�^mO�D��}�Ui�\�FG.�gs������:9���C�����"���?[Wr���lr�[��Bj�΅���^��j_\��A�Ry���G���s�ѻ��\�T�48>բ�����i�/�L1��Txqp��f\��{��>c���5�ܘy8�wo-m���#�.rmű�j�Ê�՛���dsnH����������xxzF��o�~�e7�� �$}6�!� *M�N�Â,���C��>'w�*a�ׯc���o+�����;��&��2��r܃M�+��U֦�~���OR#<c��
��c�3Y��dDg�Wl���4	�O����9�[#39;����QQ橘>^�,�D��P���Z�2�X=��g�,�P����|�{�����2L�P��V�	�l��Y�i��i�Ig������3��;��杫[�R�׻(�E-nK�_e�)���������g69π�P�Ma}���8eU���f-�3�LF��v3�=�Yu1��hEԨ|mJ���M>9��XNԎ~�����R3x�{��f�rkv�!d�%D�9�ms�ۑ�"�*��,פ&U��1}4q�s�u���O�S�-u�,Ai��Y�f��-d���('��ϰ1��_��6&|䍯�t�x@柌z]a�^��y�j:8��30�W�i��F�u��i�7&^���]x�4�˲}�q�`܃-�]cw=��T.�7��b�P|�(�nY�<�VH'��;O��1�P�<~_��%١��N%Gc5�"6ѷɮ���.�ۃ_�i�{�6�O6�Y��4��n+t�>QQ7����i�b}�Yb5|9��{9�]ȅ;�;��Ą]]wɛhq&r��~�5e �h3���Z8N,H��@�=��
@@�IJ� ,��f��<<wjr�\	����O�j�K��3�nQt���`�F�PH�~�IP����mwYn��[��+O��b����"y�	l�2a��&��Q�����n���]�5��Js5�ٲJ�J~$�&�;AxD���./Ƣ�i�t��f�0��^��Af��X����T����R\��,��������<�6�w�^].�\���k�)��I�Y$3�������ޯ�ʍ���y\��@�H��$O�!υD����/���3�P������8=N�wO���u�­�9�C�#�3��>*��������w����7��'���f�C�d����ۯ��,'v�g�}�d]�r�+����Q:U<��M[�%S�����Cy^Sl'�&-�����%	�\��~^Ms�`yԐ_��^@�@��Ew}��䏾�!Qj)�K�Bq�5����w/~���&(!�T9H��1f�V����Ѯz�ܺ$�~�%	���õ�׿L�'2�^R�3r�C֞�NG�l<��Я+%�uC�ה}v�ųMT�\r��]up�ˡ���:�vd�)Z�s�HNڹB�[�0j�b�0q�������<�ٚۻ�u��Ք���=�ڋ6v>��1R���
#��]we�<h֍��G-v���W�j�W�m�� �5<')5[t����}G����!��(EJ
?o�a�B�ʶG�����yN��������x���d��?I] S����B�j��4r��!=��o�<��>�k�糱I���h^�9�+|e;�v]����V����^��x#^�����K}V����nj�h���\��ҕy���&~m���d@i�m�YEV�fiI�s�W8՝����{t�[Y�i���*T�:a'I�X��y)��
�XۯGx�=s���{�/��;���r���w��K�*z� ��z�}|ZCϻ&ƥ1O��*S.����p�)ЃuN�j�y���i�_R���g�i��z��C��_q矷TH�d���U��m	Φ��ʢ�r7�t�|��X�j��� �V�GJii�)������&,\�<����2ݡ��b�{݂Q����6��5���{�f7>�R:r���� ����)gǄ�S{���ݽuŔt�w����7�ϲ�����3��/��;�T* ��
m�=b����d6ph|0�@zdh�neBs��;�8��>5�>��3<�T"=��0�����;>7bw2�s�3%vk��ȅ���ҫA�s�����kx���,��Q�ԁ������u����n�!a��_��8���>�bLo�g������s�U�\�]����u&�e�����j��g�d�IK���3�_UM` T�"����*�t
O�{�>�����S|or�����?S��	�l�URh	���:�ud�}��V%0N��lㄾ��H�Q��	������� ���j��ވ�=V�)^]���Ea�3<����d%��s������H��P+�~���W�WU�f�a���X��uM�=��n�sd:]6� F[U��ь����O�c���p����w�4��˘~X�=9L�k��-���"SM<�cjʊ��
�ߞ�f/����'��ypO{<��u����N�xW�/z}X;���>:��:>�o2��!�QFl�:ʃ�f�����q��~����9�w�ƟC:�k� ��Z�����2�ny*�\�TS/sY�����F�N������Q��s*=���ԴDM0����={���h?B�]��~`�
�-�uVݵ������;�dh�Y�h%[�ߪl��&C�*�\Bw$X��Lu������H�����<����Ļ��鬮}e����\6�n^Lx���N�
�ΑC��+�����X{�F���aGe��K�3��q���n�����1D6��M�������b�^�B�x�Iqs�7�J<�S��8g�K�a�ǅ>@�S�W_N�݇͒��q��a���I5�"�Њޣ�:�Q�{�Rø�C��8�w	���l��q��.����W��~0�����0�f� ,��R~F�pj�"*�,!����5
��w�����K��=�_G㤕����ǪJ�UfqMK�9h4��6�����j��ʦU�2�cs"��-6�z��MxN8�#k�m��he21�(��;$��O�]B�q��>,TI�����Ϸ��=��|U_���ߤ�;���FŎ���y����tm1�?���3��8�a�@|����*��q�u�՞���
sl���qż���w��5+Ȫ�w�ۃ���Ͱ�a"p��!F�ls�Z^�Qs#[�����%����"��0�1��^L\?�3^4|�?jDgQ@bx!2�|�
Ʌ�3Q~<�b]6�m�Llڤ�����0���H�TRp�j]�$蘂P���k���y��hޜ��{�^�]�?x,̪B��}�!\7;y�"�k�0g���G']�����_�j���&G8�l��&�^��a��_�Ì2x�T�d��i���"a겖�ܻ�v5b�j���p�J����wH梯�-�r.jc���i��v��
"X�_���3kUmv�VX!��~׿�w���ر%�};<�G��1q��4Guryj�
"���tK�-jzvHh �J���S��%��Յ[/Jw�՛A�-�;��8��6FZ�K��V����
2����{��tι�Ѹ:�y؊?H�q*V������o ����*U�*Z�&q��1�0ظv�/争_5(�fc�W��o*e��`�Zhl��!���]X��q�Tq��hg������~J˟���*&�D� mb�fs��#w����4з.�	ڎ���� �z��OI������F�z��������%y��W�gln�N�3�eCė0�ܕN��38���f�>Q_t�\��(u�WN����1�9%��<�퍧��tg���,���K��)��q�\��ǹl}kH��R�Ѻ�w̔|�ȿ0��2�q�%�"y��T-����7 &��8���p��������s��]���^i<�F�m�֒C������xԙ��n����������-F��7L�|N#1a��˸��_SE�a��Np�w�ͯ�����T��1C�Ȏ�C��V�%%^6m�t�e<��u*�L��]M3�W@���8*$_�Hts��:u�h�0�~ot��M�5�ͮ���f�s�;�8�w��K�3E�9�.^��J�lĒ�A|�ތ�e�j�c�6U�n�Д�H�Ŷ��)Sϩ�x|��8k��8���Wd���u�jm��ƫP�Z7K��*�)p6�h��{b.���l���X��e����SQYf�=�%d�9R�6A���|<��{@�%;;���cs�a��\f��>�H4P Ѝ"ҭ"�#�D�rT�v����m��K62�۵�������~��b�)��zm�=�y&�Q������\�Ѽ��M�鉞R!��X~9��x�	���*QM�E������3��^M��ٵg�� v�)�<��[S�ʤo���%E�blȗ�w�[]8��a���{��Jm�c���n��i�Y��O}8I�TJH�t�և��RW�T0��6����^���>6&���N9Ǒ��J0_@�.*gl�+o�ַ�5ym����e�э����q�I���2�j�{�6�WT����z7CkW�D�ƾ�,�ּ��WX�
2�'a�QxH~Ь|�}j ���!�8���oo�iMxXt���0&/gG�.�Qkҩ6��K=�+U����l>6��
ynQ�髱۶���~xdv��h�C4�)E�9�E�n�c��B��_����ha����9˼�s����/�/��'�;NY�Tfw�+���S	jS�b�k�+������,����p�SB��0��r<@�����n�K�n�z`&��1矱<	��F~�=����Y��ʇ�ݛ3����̵���,ǯ����Pދ fw�-�6�oj��%�a�3�����: ���+�r�46j`f)�n�-w6w�q&{_>�Ҧr˚�%��j:�fi7[4�'��%��'���w��S�m���{�5_=������U�T( ��>9�t�A�x��|��2,c�v(kg֢�A_hꔴ�^g���s W��{,,YT�.�^s��L�(��ˎތf��1m������� gt�� LAkxћ)���	���3��*2Ơႚ|��/�%�����T�ȡj9��̍�x��*���u��L�u`�u�]�����T[	�Mj�i��zw��b�7�W��=�E�^����P�P~sȜ��e���J�Ki����E��(I�gbH���d^��\�g�����ew�XA���W~��{ܒK�?4Ԃr�;����K�j���������,V���{����2w)�K&Y�Y�2�����D@����&m�5Ҏ�Jq�L#������Z��8+�:K�Ġ��r�����cc��\���Uc�tj]���v�O/��6+��{<��}�t��_ޚ1��v0gz	چ����i����9\a8b�Mg?/�߫%�ʰAϊXÇ�zC ofD��:�n�r�N���\Fη�*4���O.����ޏ_��6���6j�����ɓS1M+Y�1��9K��-$J=�ס��A��m�z��96	+짥Z4V-�ld���qb^�7���7�Y��X��Tϧd=\���[��X�vmL�]��[��K���n@V��]���-1hv������%�c��&fL�&E6��2(e྅�9ː��7Ȟ��44�q�95\��Lr툵K[�wr����j�$t���Χ�������sgPt܋�=.p6�F��	��T��x���Y��7y�`|�i��:�w;��cS;)j���v?fr�>������t7ʹn�/�"��6���*��v%PS�F���HEs[�v�N�6qS{fuZR?_W]��p�z0�iԎ8VV�q�Oh.ͺ{۫kA�ou�����o�b��^�b���ғRe2Y�ʋ��vX۵e_�j�䟱v�����W���q[C�T����Y.4���Ž)5�f;N���|��;z�u��b�<<�}tB�k���Ԛ(t���������Y������fYެY���5��@�҇a$4���iP�����.������H���wF��a���=�����B�
��x��l�\:�J�fݴ��E�(���N3F̘��o�λVb%]��sy��ܡ��r�����eCQn<�݂��D׼��R˽S���Q��%�a�%��01k�{�B������oNo���N�)��}v����G�����E(���NT(nIP�p�w�QV���_@�1�N��j9�]vG.�9�/��\�7]u�\rm��+(�с=D���Ȼ�-�H�`#��5��u����h�V�s�R:^��:�m�F�ݽ�
�X5.Ԭu*�Rr��8�{�:������ڳ�߅�:Մ���n�"W���N�2�Y�r�,W\�]S)r7��\ϸ])��T�Ȼ��"ƍ7�)�L�ήx����H]�l��ʳw��Mq�̹68�s��Wk�����|lbV��3Kw]���''5E+l������,
���؞9�:=�leJ�W�9��p�o�"��N�Z���6�By|�8��!2��(Pw����ȧ��D�P��:=X�t�&,(=�ëX�Ue,Ž��0v�;0""�e^7A��4�v*s�Fր����z��I�^��k��iv����U�=W���^�6�o#9;S��*u���i�}�"�Wj=W��VA���vm�f���:#������j�%��_Ub��Nc���>\��C�
]��KpO(_w���N����qtKp^��5m9�����K=����<�$7+P&�uF9`��=�����{�$i��qrSX2��#��_vl�+�hF�����R�Z��ֆkY3U�&{h���óWo�'��v@���˫����fk�`(��I4 ɍE�C>�M����&�+�su�E�09Wi�$�����9ۺ|llJC%�{����ܢ��Z�+��Х�:_gǟw��~o���|�QM4�ccEUG�4�33Rv5b1Z�kTD��TUl�(*���V��ш���Ak��0AMk654Q���J*J*����2a��*��=E[`�b�4�a�#Y��"`�u��(������Z�T̔QlDEm��t�L�E1D�QZ5ET�DTSAUlj�����`�*)�
	�����EV�;:�(�'���"��**)�J����*ja�����4D��v�*if*(��`����
i���*�lTS�Ӣ*"�***(��Y�RA�V�DRTE4�QSEL�TMSP�UMEUU-35�Z��US1]m�:��kl�E�LEDR�b��k�MU�UHU4V%����1PL%QLQkE�����wq�я
���V�Uտ;�Oxfy�C�V��Kl��V��챝��CO�c���[���i銦m՘97ԅ��b�-��5:���Cv��AG��)�4�.�:�cy�y���mъ��v���+@���!IH��h������%r2VP&�<$�L�ᦪ��(����[O����8!�����x,'ze28���\���,��/Tg\�,�&*�"7�\�qx�Z�poZ#2T0��@U}�6���S<#��Q�sceS�ĿJ��q~�p���^>.�U��M��=	���(��	��<��^��]�+Ф���m#�y�)��o������n�x�'�WT���	&tG�i���7���Y�hO�g�Ԗ��?oK��oz(B|��ۨ�}X�CT`�[�	6`�hi�Nಹ.`�qo�_T�P�z")��L�n)-M�M�R� ��KM��^MxN8�#x��oG"n�S��^12z�!�.z���-BL����q�u�ϵρ�s����3��1��;�͟�x'K��z��A�#<D�l�	�Pv��<k30��b[������>�|�d��R3�s7��`�I� ���8��z0N��F�Β��	��HQ��c�9��C��Ud�i9�����
۴��2P�I��bw'�.<����\"~Ԉ���x�'�1~k���R�SDTD��mEm�æ-����x�E��4��ۗ]~��1Y�5�͔E�-���Gϥ*������n��t�݁�wxox]��)���7�|�gT��ZP��ƞ�)�;�}4\��勪���3��i�y�|�����l|�c���U�	
& `�0������i�gI���8i����C��bJ�N�K��yw�fvf�������٢�/{����Y�˯ME���O��feO�X�t*v�Hҁ��B,O��L~�,�q�u����R����,=�(_8	�3�|����M�~����{=!����08�(^C��Q����py���1n�^!��p���=��c�6�ەް���_�~c�pvPb���k�Z�=��t��T���l�w�xJ({���u��$K�4[ Ў�8���+g��L�sC���!��\>T�cQ"��s�Ŭ�1x�w_@_w�ay�3sg�j�Z�E��T"��%Wܠ�O:��jX�:�/d�ײ�ӓ�]B��U�֯s��_�X��}4��}����<��DS��M>s'���$1'\4�Q{�A��;�J�_�E��*�/x�GW���� ������e�+��|(��b\��U�e1i{�N��g)֮7(�o'r�1ѭ�;`�,�ٚ����U���!�J!�3���
��s�A~:*D���R)��&���М��0��ƍ�p!��A�E1솃bu�JX�ɕ�7,�� m��Z�g�a�yB������
��N���F�+�V�-�}�7���L����s�U�b6�K�W`���S]�!傐r��,Vֶ��ۺ���]}O���k)�E�#����1 R�-4A L `�x3oo4�����[6��ywzE���
\ �����5�˽1U�yZa��'D��g���쫺�h��������_g��~��#OJX����Q��X%���.,���d�y�^�f���ʤ�\ghcE���R���@��
8�2��"Q����3'���Ǆ����g�ͮ���1�gټpb��uP��&w�
����4=)�,��*�����?��^~�RzS�1�!�A���ԭ�_L�2�����Gw��gFs�xŵ��
�MC�b�aC��L<����LAt's�����I~Z*�V;����
�{�>�a�:W8\ǧ�TO��aU���WB���_�ͣ�~��/�{i׾���++V����}�u��GK��&�tu���yV��1H��g�I�w��뗇-��H��yV3��X��9��+�./ի�K��y�O����E�,�9�ְ������\����'�}g��Ў�&��3uC8.�pW�9e�Imxl�ɮ��8��j���o�ҋߌ����Eԓ��aw�Wm~|K�3�8���wl�. ̡��$�Y��0]�L.J'���^T��5�5��it]Jv�v:�>�1����I�G�+��(yoމ�d6���C��W��hb��ڏft�en��en����oU�z�G7/Fﵝ�)ڸ���+���fњ�3�W⎤)	���$HR0_����׬Jt[�+o���q6�=\kY5�:ͳ�[̫}�>D�İf��d���Q���e��m��_n�4^?��
�ocT�����f��(��3(��� ǟ��f7i�jي��0F$%�f᭮`�3a�@���տ��I���I��@|dzq���3~�3�Sa\jS���q�� kT���sw�[59�5��Ʀ�"F��$�uD��X�ʆ=����_���1�=��EdZ��Vo�����]�e�յ���G����6���1�(�B����W�����"m���s(��w�}kQV/W���l��[]��k�'���z~*7�� �2������z���Ʀ*���@Lŧ�yc����z��+�T��M��g���4s�.����66�ቚ��+�������ŇL/��֮%�u�g����a���>n��-�?	ҥ�ʩB�wM��XJ�j �3�(�"$N��.������b�i��q�lr��>���x��Q�zy���.([�0J;lҹ0t����ʒ��ƽNc�7����J>�vVh��TBGV�S��,(�����ͻ�F��X�{��-j���G�7=��2��S̓�$ݗgWc��L.�(�܏0�W\��1�{՛7Й��w�\6�^r�7��Ч&�7֥�} �
��T����JŤ胥�՘�5A��|y�B�No,5��_��Z�E�L�1y��ka��7U�H�f���gimp���r~(H�)M�iͳ��w�Z"%����4wߕG�#/{����������7C�ԡq�ik��P��P�$M��0�?�ޠ[�M�#��0}��̌�wQs�D��8�R��K���1���]U���T��;P��Ad��H��z�۲*�܅�~�|=x�O��c�'{&�m_G���[ Dwfo=p|�9�>-��|����s}�L��1V����e�#��r�#�<�I��Q���<9 �;�K��P!�'ӧ���]CX��+�:�����T�ݱVz[�����[��M]�"֒����/"�w�=���*T0��f�@��L�nJs�I8���m�i�k�;��T��f�(���yg��j51b�%bV�#EOBc�0��4�1l�,�ѷ�F�?S]2��R&/�*u�q�L迣Z�����%<�G�WP+�JI�&��-��]D�)�l��.XBk}�Hn�oV#�"�;ι�ϼ^��t獍4�ƨ؇ӏ�����K�5�Ϳ�je�Q���V)�I/��u26_i�lD`ϟc�Ɩ���}���p�.]����փ2���u���w[N-�՝A��'�rcn�!�6<���]�^ w��s�)�p������6����A�R���N�Խ8�td�����RIN�6�:��{*n(�{ȝ�e��ω�w/+�e��Q�#���[ʷ9>�}͐�Czng9�<���&Gt|>o333a��|�m8�������7�KЗ�t�%嵟w��{R�n���V���!��YSZ����j��T��#k����	F�{�b��_Is�Ua���W�)�?�b�+�z~�j�w���z���!�O�x��w=���(j�H�yED�Y�an90�'Iyу2��l��R��A��!6���W����YS��G�+�E:ԈΟp�TK��{9�8��\��8�.�<�$��Qݰ����Ϥse��#�6���5���'�rI�7�f�U^�NP��x��Pq4��I�י?1��0ۼ���R�m{��i\���7 :x*�H�.|wf�!�N�Ò��˘�n��MG���2kuiS^�p�'�*Xi��sh�z���n2�z��9M
��)~���\eY�}�k/�U���X��H­k��Pd�+)�7���ۧᢜkڡ��{�Z-�P�"�p�����t�&�[ κ��"�ʘ6����웯v�گ��؆�3��H���s�785�C��ƪ��I6/��D`����=�ū����ne#ҠI&���lu�Ť����KCc�ɭ��;w��N�8sH첡���{�Z�<@w)k��A�;��v9�M���"�ru�5�c�{"y�X����3�D-���ՂK�sxZ�n�g �NT3&M�=J���y�����`���c�]r�)Xc�%�������]Wk�J-?u�*�kP��= v=�A�1�P��.v}W��d��S��d������:-f "��E��@�W#�+�m�r�����.'���!"6@�����!����Uo4�H	WUFI�&��~��xmF{��&Ly��e�tUT�qh�X>�~>ُT��PL������W�@��~��/��7X{m��^�~�Cz��cൕ�$�r�H�v.Y�^y�{��y���B�+�5��B-n񍖭-�+�Q1���͟E�&�W�bL6���F�� F�<X�B:��<7�2A�q
Eܒ�H��J�>��g\e�ҬK�αJ~�O�e�"�� e�F�l�8��Y3��]��@iߞP��Vǳg9X���c�w����56\S�r��靈��P������1v�8X��}0x{՛Dm�^��v������eۃO��M�n����-b���l8��r�̓�_�~8�Ĺ��c��p�b�*�W۫�6X~�׳T["���9ci%=�V�p5¹���.��ޮ�zw��#6�8%8���Ȝ3/z��}�\�~�ЀY��T���~�Μ�<��N�Yp3�K����ܗ�D�>�$Q�2Ew�W!:h��y�Fe�h�7�)S+���Gt�
���"��u�G	�vk����~�����<���p�$�;�Ņl�WN�#��p�C�Ϳ�L7�W*�?~(<5��>�y�z�#��������z�pk�^Y2��K]{T�ϑ�w���\>9�D{ 1sI_Z����oFc��޵��Ud��^�w� �&������^�ѧ��v�ڊ�~�A�"�GR!�@X2����^YK_���jFy/"i�c;����0Tw&�Yތ{Q{m�鋷�DD��#[ޕz���Α����K�k�_��-e�t��7��f�S�Y���e�*|����xi�eF�r���04��J��������T�;�8e3��c�P�0����*s����Ly�,sm�Ln�Uq������������#������I��_a�e_g��}�b�ٽ����çFc�M���oì�j�}�p��n^�.PE|�6R��%1���c�k�n]ܲ���e�wI�̣�9J�(ڭa|L�E�sN�όK볢c A�Q)iᲆ�yMNO����xCj�}B��+s���J�ke�Ϩ�댴d����_^��p�Ӳ0�)��!�N�?M�j�ܥ[�R�>��
3�,���uy]v���;Y; WV�/�+O���)[H�vx�}���K�]n�|�9L�u"�/�/�8VRhՍ�[�N.��ܛ$���#�ח�q圯���)����2�e�Ie���\H:3�u}Ӱ+���k���������.g3��{6�R�*�
|  Nq��L�o�*)�������cs�I|��S��aUScWƂ���q���vmѼ@����'���L�2��}����1�'�O;�k_֧�ƹ�NuY���Z�'��%3Y���2�$�����B&�Ǖ7�<_̏�:�69�~�'%^�{�gYS$GM�ɋ�|'���,	�����wX:%���n#�m3�5Jw�P[%��4У�nW{oj1{Oyj�5�vِ����_�f���`�6���-�?C���3ANB��<��M4(��υ�jm6pt���BE}z�<�Ci���z�Ƀ��DD��3�H��C��[����߻��f8H�|`�K��f�G���J�����M4�Bm�%�+��yKr���%}�7N��mnkN=O	�Łz2:��8+2'ŧ�eV5�)d�lK-�8>�]`4�#};=x׸U�2H�2�{�E���3(gЏ2n��z���j:$���2�h���s���&�f��������St�w\Qy0(^2�H�����Hʕ>8=��0D|r&�)�_p��ޅ%ʖ�Yo��<}2�խ@�+�Gǆ�
�Tw.�̉����wd��������XD�r}-���9�#K��u�݋.[�M�D9}Cy1���gP	��fR@gu���v��:m<Hƺ$F�ە-t�� [T]��ٳ}�6MѪ�����r��W]'T�l�\�}����z ���l�"4d}=	�����y4����gt��bY\������⁊U���"��^���ӳÝ(�'�WP+�W��IW}���|7/8ud��j�=�|菦��5
��뙲׼_���64p�OM�iq��y��Ԟ]�]0�́	���B^A%�鹑���
��[�n�q��gɯ
��du�z���gP�Ȧ��J���>��+���lܙ�a8_˷�v�7��y�f�,���y]@1
�C��V��%uTW��q���_g�����	F��]�W���8獉d��ƌ��[9��B>��}��3R���G���=!�O�R��pv�2+�-�!�ɋ	�=�R����p�wQf�ޑ�6��S�����3�9��g;���0Q��.ǽs�����r�ě�nivL������շ�\Y�3]�~�A�v��n��l�8I�o|�E�9N�'�r�b���,A�����ܯX��~ZM,�2~�9�n���QϠm}�@��L�if0ݫ���9jջf�^�ч@���h�۪�j�W$%�}�VƂ{�$il��M�:P�ɷh�:�w�x��[(F.!Sk��g^CB�=�7%�F]��k[�����7)��:�9S�,2"����S�Mj��8s��Ƒt�\�ԟK*����Ŝ��N�̓x1S<V�L�XkN�(���� �kFѮ�
EoF��ۙ���9�_���溒�A34bǋ`r��od��!Q`�X�1�b�;�[��N�2��=����hm;2���N�鬛K:��[|��h�mvt�;IG1ܨ�n◖�u��.��nͫ���;��Ww'Erq������׫��}eo�R��� ��׉���1�%D�U�u��Kc�:xP0*ۄJ©sE�`���F���>��v=�+�N͝���R�u��''�{�����9Y}K;���y�K!T1A�6�m.��^�@��(��i���L��Z���MX��z��[��˃�s#�>%[;f�Z�|�	}w�oRT��u�N��K2���ͥ��|T�b�J��X]K��Z@Y������8�gGÚ�����]&�q��Ȇp�g��:o&�j[�}[F�b��Sݼr��/��y]�b� �䎤���ht�k._��ڭ��c岈Ӵ���L7����0�Ļ^l�s9k�����[�����P�˃7DHu���(�lbI�X�г:�.���嶳6�a��<��jj��H:�tmV��(�q~�O��8����۔���V��v����o�Kв��TꕗJ��.Q�/���T�[�y��T���#����(]"��{��PU�R�]e�ެT��V=�1��4�Kc�%�8��Ia�V�.5yGFѴ�n,SF�Jլ��ox��Q@��1u�ifP�W��7����B��t��Gag��� �oM��gD�����k1��W�nm�%�j�]t�I�X�XԵ�m��J�}��r ;�5�b�)��έ]�JN������CV���y�3�=�W�æ�R��"�+;b�0�K9;�k��S�ն#��Z˖�unҡI�ڧm�f����I`�BX�[X�wrF��i����^5P�s�[�=&]�V�u����
��\�'��)oE���|R�����L���YOM��2�c\_�c��7��[�t��vᱯ��N���[i���yr�L�i���0,X,,|�/��z�=}�\��9�*�gھ��M'AS�꾬a��hT�M7v�<?u�%�Y��7'���~��!�&����5�e���7x��V�N&�L��k��7��3J���@�4��Wr�Ow/eQ&ʙn�2{DrXn�͊�;�i��3`�@��C�a|�-5!�]��XنewXKS/��=��h�����a�ݮT��P>QQ151!E��55}Al�AT3]j��HUDEj��i�$PUV�4�kT4i5lj�QTM%֨�")���TI0�55SU0ALm�zt�ғ3T�Ww=�=��A@tb�"(Ѣ"*��"JJ���b5���$������"�UDv�%P�AT:�֊�-��j�(�J�֤����M�EPQSRAQAKQR�QEQA:1QOF��huMMD�i��/��*�\ILG�c0�QP�U[�b�JY�a�������**��j������i���'�T���Y((#mU%h:�-�Ul�QV�v�QADQR��DQ4UT�L���ux��Tz��ܠήu�/�mҥK/h��@�w9sfN{���t��3�ձ�g�v��_M��{�9�9���b�~ƆV��}j��zs�V��vBz��������s�2nxר�r,�ڜ�_!�'��{�HG��K��L�9�\�Q�)��^x^mU�7�xZ�}5�P�KS2&x^c��@��~٠ƼH^�y^'Մ�B)�&����a=$��j8]��F-Y�����3V�����yW�g*g�9���[�1���#Ր��D�7���H��Y]m�Q"3�BpӀ���z_�\��4Σ��/ie[xkP�'+i�FǟV�b�S���3j��ׂ�����Z��S��+x�-��TPO\���P%�,YQ�Dq*!��5��w�
�>�j/(%������P���������{��u蟋��Wۭ-�wX�����{�Ӳ8�7�.�6����;���vC��e�?��=�E5z�ɇ!�T�ӏ�Ty��o�Yq�s���ߌ��-¢r��F�%��D�ɮ�<_�Ѯ;�»���S��UPI��ǚ�)J���xi����ޚ��&��:��`�9���{І��q�MѼ�*�:��n0���ta�H����ՙw{�����\=���u�,����^8bH^���t�����-IJ|`[���̔���ʈ�\E�fͣ�N�W��FzBUu��*r.�74F11Ds�gs{���f��X>��$��k��1�zO"7��&q8��F�5����T֏x��� h�$�"Ǝ���;�^r����=��T�X�ط���5x�����6����3E�9�._�fb�8�s�u h�#����������͌w�v�=�i���aw�8˵�1�������}W��5UR�?�V�$뢢t�j˝*U�f��?r�̚�_n��1T�}�&5�:�U���>K��`Lw��>�^}˾y����'%��/X⚅�V'l��[*��E��#k�����］x��͒f��Aע8}��~u%%~�Y|he���T>��o	����%�ٱ�����fY���V��h�nJ3����h��ŗPٙ�:��S^��q�Xk���jI�����+C��X�qɇ���z�ǵ���q�ι"2�Hӹ�����.��;����bpTI����dc����X0�킧ț�b���g@v8���QS�MUD P++e�]�4���0��.C.��C@�C4�yJ/a��.�z������ee��ἂi�r��]�0� �zjn�v�QN� ^-�}ڀ{9���r��-bPj��J��Y1���r�8�W��=�e��<�3"����:�~U0H�hNv}}7�ʱ�|��v,nӍ*]EW	��X�K+�]hHH�-�^sW������|����^�RW���\:k�m��7�_!:z}�{�厹��n`'�DcL:e�R�7q�����
�����i,�嵸k�ڔ�C���U,>�ck�a��"�ST颖�)��P�x�����}E�Y��̐��֢�*��Q��6��`��=<"q�`��A1� ֎��P�18�q�W�u�!�0�	gζ~�ƅWV��`ޝO^��2���Bֶ�V������r�G��,���5c���L���x��s/,�vK{{�P�Q������uT4^湖�rs*�\��HV}� gLJ�s`jb%A�}_\�&1���1Z��5����u�9����?�t��Ge2?J�@o���A~�S�N�xԐΈ��B��������j�<�}=͋�.s�g+]H��`��h�Ω�=r%&�jA��z��T�s�b��J{޵1�	�s�u{����z��)�
LcH����_� Ct��x��(͂�}Ҏ�IH��#�ʂ��)K��Ә"�0�_dd���ͪlld��� 6w�t�}��E���)�FB��L���1Q&�Y����%d�G�r�b�~����&��E;�>`q�.��W�JZ�Z|��[dx���it��O�e�;���âN�"��7z���T��f��T��S�Յ�nP�7G1}'T�9W;]�j�;o~��[���K�5�!��� �}ݠ�6�[pc/m�mN�K��"�i������Ht��$ҮDۮǁ'�;�8=sې�Ǜ��E2��h���`�:��_�y����}���2�Y4�skM�,C��ٱ�Y��$�z�$h�h���v���6�_x��h!���<=�X<��u�ΨYt����\��X��\�	*/�^C����n�&Z�1�b����Ri��nu(&�����%J�{�u�XYU%��%XO����*�)AyF�0�XP�Dhf�=q��WQ�N�n�#󱭨a}y�a��Ƒp^T��(�O�~���c�X�r�,m�卻�_�~�袑��<DX����2vP�}|菧��x�.*y9��]��w=Q�͊����SJ��&s�e��Apy}e1 ���/�xX���R*ڍ-Sk�cW���I�^"�4ފ�l�V.]�x�a��U��tX�����FX��n��u��Y��twM۩R�^O�w�f��y��_�I�}����(p�B=�E��E��<�^�='�CGq�e���X��c��ZT�*�Ҥ�^�x�+��)�2�ਗ��7��y�J5�be`���1�Q�/�:d��^�N�i�Vy��Q+'�烐F�t���r��S��LTt�;��hx�+Gub��ogXm�:�7�cn�h�/��wWײ6#c�O���w�;��z�ρo�Ц���:�v3��rjk|�gr�,;k��d�`9���>�׵�Z���lp�E?�l?����.dckX~�.�8�������ZI�����mo�V�bvwvx�#}���V�I��*�{�h;gq�v�c ��"ĕ6�=zӧ�Ʉ��Ƕـ� �'����=�	�i��8=y����h^�����4P9�)���W�r��{�sz�f4�Q&��?����W�'}*����QB~V����_uթ����~��ee�c���g&���w�a�_��k��(S�ڬ���~9H��=�}W)c��5]���]��g�*\H��'�:�Ԯ�IL��A����u�{Z.�}8Jf��1��e������?�0�7p�������-S�n7�2���L�㘡�s�nۜ'Fi!΅�G����ݟEe=@�/I����F殁��p�=��8��+^�TZrs˨^д�l5�������N+ջS4�x���������|�;V�{�A�ׅ����f���
�K��y�C�,Т�V��,�jŶ兊p�30T�Y֯�����Y_`�]R+'�X�)�&��`bۚ��K�+�:��J����@��[���]�67�z�[���#ݏt�������m��w�.j�)��\��n��S'g[/X�N�ܗ�Ӆ�6���� *��c]��zP�5!��ߚ#*���R}Q����
"������}��5��#������z�xm�/n�(0�)#�^�j����Z�U�ewT��{�>3��(T]Q�Pg��^�h���%���q���d��g�-�|�ю��1�D�iw��<_�V�o��7�L�C���IT.�q�óc��Y���͟\x�҈?O�i�p
�j�}�Y??l=�R��&���0�н�E��ث&q8�(�Ƶ��*�ׯ�V�`���C7�9)il����٧�YH}�4/�Ϋ;n�}���ɾ碲W7-C��01���(�6t�3�������5�6��-WƢ`��Q�	�����;�I��~&�Z��֣�EY�.{;"��qH��j����]�1X��Oj	��@~�N0�ܟ{��&����U�m�]t�'	�ힸk9�/.�ͯ\D[4����Q�%��k[Ι�~�����5&�ōzk�-M�u�Yq�8z`�"9�H��z��E��~;�G�[VI��P���J>��#�N��������!W�{U��;kJ���l�biWa�a�g��j�a�����*�/_��m˚����p5���s����U��oB�f�V�6������Qˬ��O<t�M��Z���Щl�r����>�N�YM�ft��w�q�G>_��2��z ��@wo|�g£-�\�K��d��:�L��"��+o�ְ�Z�s�]��.�l܋�]W{;6vi����nA�[���4� ���Ʒ)�ܘ|n�g��^�7[�/��D��SS�U�v'�%2#}ȅ���8>��	�
��s뇅B��x_�}2��%>D�-��; ���Ց�f8L��!���A_�ʍz��%�=�·��NC#C$hh��ͼ�䛃�]{��푘���׏}
�z�Qײ�,u��{u��jo�<2��K�C�Q_@�8<aǩD��yk��9��EE=��r�
�R���j���A~�����MhD�U���"Jc���}~��k}'�N�I�a�Wƌ8{4��M�c���Ŵ(> �c S�q�S�W���ut��PԄ�[�P����G�<;8ؾ*T8��]N��Gs����1��a�b��D�ټV���ږ	�yB X�3��A/�\��.�޲ްJ�
qޖ���H�.�آ�L��^�xz�TӑA����ί���CH�*0j�)ң��U�?.��o��骧��/A�eS�I���+n�\Wߥx��T�Z�?wC���1��Od�?d}��]�=�{�f�fy��b�
��L]}�GL3�ם��{��sּ��y0�L�-x[�����;92�Mǚ.��'����TЕs#-|D�Gϱ��\�㫣2遪�0���v*����َ����]�?��}g��L�J�T��F�Ty�o^x�d~:*�>25��f�-sre<�5������c��Q��|����꘣�K���K��DL����$u���ǉ��.8]ê��b�fd�N�rw��m��H��T ?*������/R�油�D	~(sÌ%����"^�����3v���<���T9	t5V;��#t�8�tND鱱��K����?[#��*FH'�ڄd+z@q�U-�0����"I&�o*+W��'"|�/s�Y�8�E*�^�(��(��Ɖ�?b�mP���i�Z3f�Z�B�j�R��Zč���# �GA���l��<�#ψZ�om%�b�=�(�Y�u�G0�B����E�9�@Qod�����R�<Y���i��e���kv2�_����2����`W��fE�:9�#2"Tp|kC��#�����3>�T�M
�n�]�/)�
*��v%V�P�}���T�8+�,L�J�����7��9���EV�P�
�Fp����c�E�&���Qp^T�y1όB~l����7s���#x64��ַ��&g�B&��T��u�޿"y*O@�m�Y]:E��2�`j#~S�4:�����Aؤق��G	Y�MN}�B�!�F�\���o�J/���^�;�S{Gp�پ���+�PE}Գ��b3�Əig��N��O~\V�=��,X�A��=�"!>�K��k�<2ȾV���y#��/a�{}D�=��;v�fM3�ۺ�{z�j�����5Ʋ��5���M%�o]F���E���0Ņ���\u���A�l����,�?A�h�����l����εР{�<2�/R�}К�<�3��F�aJ�gg&j����Z_PY�E*�5���l�b]�sZ��]�.��^�t�#��&}F��a1��ƶ;33�`�uR5�2q�{i��� �W�r��8C;��ĳ�Xl�6�7Ad�.u�p*|f�[��C�����c�w�ӣU���~�]@����gS�y�����ή�xS�Z���6的��c�$�m�h�)ہq͚8��y�I���y$���\ܻ�=t���&��%!M�̉�[38�{/'��2��w�;E��Ux#�h��l�5��w˰ҵl��������N�aVI����{��q6éj��-��9T�i�!������Yzřp�Xj<�he�>؅?�j���	��at~�b�-��w��d^�ȏ��C%`/̘:�Lc�W��=o߷j�bl����X|�sCT�FE��wOh�1���+N?C޺@k �bX)TE{ᛞY�L�N�Q��'̀60�����;��N����+&Tt#E�Au�\qINԹ��Lz�����g\�}�:\;/�����o#C��FnGgu;��j����0;(p�Ϯ�c��T�p�,@~YM����`Ի�i��w6l���0��\@^�~x6����&m9�l	k�*��f8�豱N�GZR�n��)s�Y�I��!�X3e�r%�Z�f�4_�������ҧ��&����`�=�:�z����pTP�s%�/��X"bxO��3�k�Q���Zsk�����\b�zO�Ѷ4�̀V�m��b"���t��f��a�����>K���b�xI��
�_y�]��\��*X�����vtke��6&;�3�i�k�c�=�w����r~;�(b�riz�B-�J^���=�d��s>�B!;ㄑ�ImxP�
t�.�Q��"�ȴ}�`=�'�GB��.(�:�Ȭ%Ra��y�=yfϢ�5�Ga���i�p<�i��P��n�_:��,gT��K��+��^}�lc�e�ҰO��:9=$�+�Y@�������<��nU{�K�t��b � �&���Hs�k��>�V;���P�cN��K�
8h�WG.��4hѳW�цn44��<1!�]��a���YEDY�ʺ�Ue�	]���	jU�)�_K�Ԥ7������&�G',y�p�p�bF�k�7�u��6�f脾D/5���u\��E����E /��O)��q�ͭɍL��#��9bng�<��y������L������oL+�]:��G�'-��R��ڣW�6�#���w��.y�-3��ulD�O9>��Y,3L�8�6V����+��C�ᓥX�������P[3n�hYC5O���H�˒����[���҇�d�mL��#]\Yʓ��Z�j�4q޺<��v��x���
O:d�]؆EٰE�w�1�Z��݊���<޶nb�����o6jjdɢ�|NZ�+�2u\�x�=%^$
tS��j�L����3o	=��ɵ[F�#�Xr����1 C��ss�P����_*(�S�����5�e$����[�^����z�4i2��Z�W�.�.�T**͢����R.��e-���>�4�tvrݺ�c�J���c+fR��� =ԕ֚U#yu�Ws���g�.�v@k�moZ�zh�E���Q��i���u��&5�f�d<�̏�7]��FY|x28111��&-"����d�\XTN7���+��B�n�g�����qH���kre�e �'qP��S�����R'i�'�9-�Vݼ�.]q�'q�_J-i��WMT{�m3j��Wz:v%be�Zru����u�(�ɬ:<���*Ҕ`��2F�Hީ�Jl�w���n��7�R��@5��t��9�]	�[\+�����y�W�9'P�-�\��aؚ����i�9+�t.;�eX�P�=�3�嵭n�gf���kwA9S����
�y�� 
�V'h2�N�J�ǐ��Κ[���x�I�����2+f������)?Jوuav�϶B�3����s|�a5FDm�i"%p�����д.<v�[�w�7U��{\��|##^�XE��!��>=����-hK3:�ΥՂUm���d���a�����rm:]9(M1[�v��	X��]��f�O�Yշ�8:�5²��.�WPӏz5.ҕ���塡����k&�&}�:���Vo�����}�r�3�{I�\)<�c�r�R۝]���fV���"ևl�R
��fK���g-@tr�1|��U�wt]o�T�iA���0 .s�ة�;Wl�[�I�r�6�ھ�.pQi�*���.SR��V{��X���nh<�4�;�=�}J��ǗKYB��̬�w:�]gt�n�9���dަ�Y�W��\pMN�u
+�̡&�7��B�ϪoC"��{�-�3y(Q�M &��F�Wk�u���ؘB���+4KJ�s�5�{N�1���\�	�ݜ��f�o��=5���il �@�Ԋ������x�"+����Y#�=�z���ځ�	4سDT(P�.�$DTD�����h��v��b(�Y�������2ES�4j�Z)�q!V�*B*(ћ�5�h*��&����	���&������������*"(j!��"����5T�%1TCM墈�%F�)j&��M���(�h�LSElkgy�,AME� � �4�v��@jF.��UQMt���F)������:<ڊ
�������@m�UP�DTDRCMA�ZJJ*��	����������]�PLSM�i�*�k�5Q5DESTQ�h�t꒢J$�*�	�+Fں��Y5TU�F�6
H�(*���ۭXˍ�5M$��Q�:)��A������*�6���a�|>q�wq�U�F��������&��:E��R5j.U:5v�5�cUyw�9_������ރ��Nc�\�-o|z��쫺��TJrJCH
H0dw���&l�g#	�����6k������Aj_-������hnϣ�Mk�C��4�8����6��Ś�K��	�-AʰY��2N�ZnzaLK�0�X�n2��ag��l넌���g����x������&��;��^}��G~2�OfE���i��rT%��6f��h�4�Hn�v,1�*��@�-���9�K]S��(ͻ�t�㜈��Zt�� [嚫\͆�J��p2_i�Z���0�����A�9�/��'(#X.�y}P</���ծ�O�빓�j܉���?I�$�|ϙ�ʝh�0w>z���ǵ�@��?���Ʒo�}�eK�q���a7��z�E��i��j�)�H�	�u�Öϫ��s���F����c�1z��0��J�}�N4P��٨��Z���C��|*_��!�W�A�C1����x{r�b3A�u�5�هⴘ�\<GV5�k�O�B��6������|)`!��$�q��<}f�7FU>�/N�M!��Ra��&)��EI�X��j#�^���%'5Z3
��&}V�LNce��7q��6�M��/Q�F��p�W�rߺ�FL����@ ��כ�t�c*=�k��4Fcғq����ԫ{Ҙ�]{{;]ŜU�fC��ٜ5cPu���/��w��҅�Ꚗ3�3�vu��(˟ó���A^�`��5�.����e���+�3|9���<�W{�w�g�
���D������Zf�s��c�����fA�9��=2����+s~��Ggc��6�Qf���p��B�/zO�OIs�5����a3e�"9;0!4 c�w��}Nj��?l��{���VЮK�0��_{��i9�_>®��i�UP�]�f�D�5�:GyA���E�E�<���(z�;v���k:g2�q`?�E���81�?	���G��㴈���([<v��
�Eσ�m03�Y����Uks���1���^�ي�M���%�)O��nzaR=�S�sn�����f�W:�Ƒ�31{��<l��8�
T����:p(t���M��:]��Z�����3�^q�#_�ɨ�qX�٧�6���^�cA%(7X�M�]Y�8j;үOHk��N����}E1���/Y��e�;+�*;=���&�g+���{)�M���.lß�����k�d`������m�zu3�{�ND���zUc{�Me�
�s��Y�u�÷�J�Z���N���s�d��=��
�����Ҹ��¹K�lRt����L���0Wf'Χ}�TZb��E�����dbRNPr[������EKΓ����>ˉ���X�7R���\�X��>{4_��G�Q��Fm#�b��ʢs�`��U�7?*���z��N~ke^��pL�Ӎ-s^��;�n�K>�sc�e`�3W*2�h�D\*�ZIΣ�"l�15���z*K�+K�����I�^ǜħ,,����9+���8�[��q:���j`iEȭ��3=-6q��.]�W�xBn��fqi�q�\�=��y*gE�\5�����|법��|F�\q�|���_9������#c�dK+�.ޮ%�A��On����wj}a9�j���&�z�m`��8��b`i� xE��޸����	q�������ܑx��!pL�v����+7�{����$m}� ޘ*6��L��x�I�,TI��S�o�W��S����*�2��~� {"�y���j[%�׌0nb�5���C�t^9XŇ�}0M���w�O�,��fVo�9�DR{�3��猃�A��P�庼�a�|��Z�f�������� �1ȰP�{���%�򁤹���a�y��H�&f��b���01�-�p�
�o���p�S��C�����V�K�ʹM�/>v�ˤ"7QՀ�T���7V:P�'-h�!��^ݩ�����{��Qwm��/��8ވ�}f?=������˔U��>�Yh�n�IV��ϵ�����x�y�I�ξ3;w������v9���#Z@��Z�����{d[gwi�c�g�}�H�EeGEk7|b��|�x�US�0\'tp�D� Zv�^���~�8��|���Kd�S��u��w���n�˫�uw�c��@�L
���%D��d���O�8��V�zQ�l	m9]�jʱ�c/��m�{��;Q�x5��M�}��L=VRu�~2��#ߕC�������y���ϟ{2�<Ε@���-|�2i
�G����m�絢��=XL��Қ6/&�s������㐴B�v�~��=*�g��2���L��:�qe��%8�#��,Z�r���N�C�b�w���.�C#�E�o���bUr�����E̩���[+`�)Γ��ޔ�,�W9/Q�>ɧ� �h�fGn)p
/g��χG���Eei>�^W4f�*�����֝��i<yQ����r�ʂ���C�8w�PbkxI����u�}w���q
��� ��Y���-M�n<�q'>Dh���z����@hO�Ǌ�֔
��n�����󚛋L� [/�fL�����ڒ2q9�E��*�bC3te�`�%�o�5��b1�r�]Y �rA}�ζ'��o�XJ�u6���+:Vn������n�'���v�͊.U�]�/o#��w�d�o�+���%BQ���qn�>���,w���/���V
�T(D4?��`�����dSU�&�BhO��?m�TNTr@�K`/�\"��tE�N���]�wZ1�x��6_�\ys���L6�O3��l�.�f���a���F�����.��=9���C�*t��v�zO";Mŧ�ѡ�k����q���x�K׼d,�����$_�yx(Ϻ3e�(�u���cm�*)k���#Mv�16�S�����G']|T!� �|1TK61�v�zE,�]\��kĽ�-z��3;�F'z&]�1U	��#��f��������3��ÝQ�̷�M����gV���b$/R���^� �S^�ph���/�d��_��B�QfE�<�g���c���m�8S�2�Kո��.�)�3R�{2��%6׹H��j�9�d�1Ԏ��n+L4�{���K��~��H�LU�QzW�خN���eR�>h	e
6�k
k:�>���׎�%x���,0��KRMTyy�1�GO˔�b�����S=u�������Z+7�����Y��)\͢��1
���n�Lg��%B���ث�Μ���L�+ڦ����?x�^�ƶ������K��+��:����jɗ|��*=�VԦm*��9J0�\���]�ԸB�mk�P�b��=c�;uԪ��N�W��̙I9_�/|�R����C������m8��3��Y�֧X��p�6?��.��C�W4����ϒ7�=b��*̡��r_q��P�6�g��(z����-����'wjyql)c�	v�\��)�?6��w�ۏT�%_q�h��$J,>(�4^��k��֎�6l�4�z)=xn�5�2�H�R���1R�vy�y��n^���HӴMӼ��n�,��V���F��W��k�2/��/�H�ƌ8�6��YFK#���	�l���������˛އo����	�@�̡ܹh�	����b�q�j\v{zu=ydw>1ɶ{QT�F�*̓zH4�sN����.K-��1�� ����53��E2�"�����T3'\>�e�9P�g�^9B����:zfF�aqq�F���i_� |;�Ʀ ��{�sA��E�iqvEX3W���l�-�C֫�7��9_�82�����ҙ�r�7Ţ4��0�"vsǢ�ǰ�P�c�I�ʭ�Pq�	�dC�6~�c�+�0�����qL�L�.nY�W�f�!��6 {j.?N �ƈ��"�b��kCXK�V�ƞV���ޣ�3z����=���P����?w^��V�h�r��V�m"��c�/[�wb�\�hV��kd��-Ө�1km1���yd4!|5wG4e�C�qw�_��0Fv��Z.�|�r[�;�(�
�^e��xzw�fn+����
������8ug����[J�y)�(�3�~��"�m8�/GvxuvRI?~���CV�#��Q�~�xpt��SKP��~s/iB�
&˜�P��v�k��D����ۺ"&��2h�80z��&8T���n�h��D�5��Y=އ�M���2�jCЬ{�Ȫ;�Q�4N	&ŉ����j<��NN�Kq���Ө_�U�6
�y�p�2�h{�h�j̸��%�8K�V�#@;�����q����'�`.�FLoK
f�2�n��s�QM��+y�V�ᱚ��D���퉊���¡�6'j"`[z�5����d���f�Y7-�g��k���d۸]�jo�+%��Q�aď8	h��Y�8z�h4���\q�TS�Q�Z�G6�-Q
�zhKrY�ٱ��Be��r�R�&SQ]P
��I��i��#��9�������W'�ͮ�
�骝�O6�����xf1�*#��1�6(�1풸E���]L���LX��,�ށ9j���x#¨/h�τ�{V�q�3a���.�����]��i����A�vgyCQd�ޯ �F�nA��^R�g��A�Ѻ8�{�����`f^&���ֵIu_l[���t/N��۪��.��;ڟK�5d�O��B�y*<[��b�!IYϷ�[l`�i�{_�=^��位l����G��r��th�-�L��Ӷ�@f%�pj>�#˼jL�a%=;��4�wY^����"ضx��qY�-kT�*r_pqkb}��vqf&Om������4�0�lف'�1�Vw?Z�{��6Y��&���i"�Pqu�[�Fov��\�Ů��ϯ����;abw����+�o�CQ�9���*�*��c�wVlA¨`��=�q��q;�ً��e��i�Z����x�[��#a����(����M��/ܷwh�hXb��y./'mNek99���U3Z4ˡ�3�5�{��uk�Ν��#T�lS��3N���!D��Ī*��J�g���d���V�]�I,��4���A��P����Y#n*�����RY�^[l�)6�tK�⅓}������K�
�F֜�o:�;'k�Ue�,z�z�6Y�47�_�ژ�����e�>�����9j�	IL++5[�;�\�I� i��5��Jlmv&�
������j�ŽPs�8̊_:�gY�\�[����^w�r�V����R��hQE���ܱ�S���0����I�7�O���4���k��,K^� <�݋W��/�]���Jn&��y�O��z��
m�/���3��I��줨�^�ͻ�Ǐo]��먂i"���ʦ|b��["�<�sO�.���܋a�ѣcf���;H#���B�yC�Zz�nf��D�7������;p�ث޽|t����ޯo_ϯ�ے9� ���e�a��rꁺ�W�*p����h�my�~!��X�_��<wU��%��|����ܬ��|s7i�9��ogL�F��G�4��Ej�Jn��ǫ��[gW�T��skEJCV41����M�tWdq�uk��=��1\8h���Owj�x:l6����`����Y�YÜ�����BfXOr�ۊ�ĺ�G���li� �A������঺C*g��\c��w�뀊�&-=����������ɿ%�)���4�����	�+u��}9�/��,�xA�c���ۮ�d�ʧ�����*��x�/k���:{��剮X���_o���;��u�\�O�5�]ܩNъ�f� 5�������Z南o'I������#�rQ{vK��%sk�7K70��ܮIքt�-���OI�<D]��ϑt{7f'7�u���*� �}A��ƹ�+yoxRQ>�����w��xqݤEvO�m]]��SY���FN�7Z���~5�.�A�����?+2�wx�_�uk��N�{���p̵�o5^�q��>V w��W��Ņ
�&����]�*���>E@�Η��,���ލ�8$k�EE\�w����۫�>�x����Yo�[bk��m���Ej�eR}/�-Q�}M5�wY���{/�y"�l�U�^�yxƅװ��[,�@:��RW~8���ť1Θ�[y߅�rc��J�%oyY͠f��ۙ��Q;}=���{ណ��=��Cvz��`/V�\e�8�����^����>����'S5+7�Gh�w�f{�px�v:�W������W+Uܕ��v�3'bo�Yߎn߹�H>��	��������$�zO@��U�'���b@|�^oo������}>�_��<�|�1�N�ED̗�w�����FSdJ�X`�n˫�sb���իcB�^�Z�ѫ�j�˕@��y�볡�Y�;���-B�#L��R�Rm!�'H#��������M���f��s�ѡ�"�dH����=A�̌�x��C�Z��_�U�|C�����Uk)>��O�hܹ�n22u��D�H�4��j�e��d����h
vc:7����Tj�2��2f�s��s8ѕ�Z}f���r���y�u�q�����5�*ܒ]f�7#�����wV�X�$�:{�nW�r�����N;�ږ�|La�	9q�ZɀY�>=n���������`�9h�����Bl�-�D�}�1�ycT�#�Q�����
,����g�~ή�i��V�Z+4���:��f�:%��H]oGB�m^�Р3N���SΡv�X��%�6��o�6�N��z�)۫̢�A��6�5;<I��]���;3�kH.;`����<����A�pI�}�8k,R]wV���Јћ�Q�zfY��䌵ڱ�!�_`R���T2DV�t؏�RN��oFw#���kv^�	�[�g)ip�*_��Vft�;� �w.�z�!��֭���W�m:;-r(#��t�nM�.�Y��wL��wt�_v활"L��9s�]���)Ov5ge�6lq
�tY��8.�5��t���jL��l�#�1�
30J�^�G ���^f���b��P�-2���}Ҷ�\,�73{>�^�u���vu��m�,�F���M�qg�����7�q[f�n���c?��$'D;�O��켘�����n������tw:e�fM�m[��.c�&��V+U۾��@s�4�]N��]����iK���vj�+���e])���H�P�
���<*�Jgl�S��r�W}N�:�5��ն�������j��vts/;��:t�vMb�RH<� ̴� rZ�e��Fj�ɔJ�bEܝ��gX:���i��n��T5u�D�/u�u��8v�!Ƒu.�k�qʲ��ō���4M]s˷1�js�.�=�sh+}����7��gE��Pʏu7�X~�{$��t��K�ݣ���=L�ʣ�"
�����yw�7)⯝���*�<�)H�,-N�[I�\�ی�z��o�W��u���}���L��1Jep���2��V���ڹ�(�;�)g�FܤX˱t��{�j̮G����`���/���P%=���K#�D򬹊���u Į����C��Z�+P�w�NC�:��!#2���*�ƺ
2�tlV�U`u$�oZ��:o�k���"�����������N�*QC�nr�¢�v�=��2�-t��T��l{g�P4*:���s�
@nM���9^d�\;\qeJ�TwTW���EΚU���.�=Ք�<uhHE9�ٹԺ��{�u3]WW�@��6庻�w���KXi�
�1���Q�M�<�m�t�ٔg|��|�L�����j��|G�@ (��GN �)�����J
65�3QCN�=;X�3V�
:�qg15�� �)"+A���l�X]m���5[�E;UU'lth�J
j����Y��MvM���IMGF��EU�3v�DQQ%$ET�Qu������@���T�Q��

h�i)*��Hh~;u��1Aj�풊����Mf;.!:7NH��RMD�UM&� �E,Q1-h�.�4D�v���E%S[c�b��N�m��4���\mv�*%��QE#����i1lf8�*wDTRRQ�h���33 ��w���&Nu�}�ޛ�7S���*�M��ܺd�S��=Ԓ��(��3z��z�;�t{VIGZt6&��p���0�9ߏ�����%��;٭�[y�2ޑ��&��g3ai�b�Q��Ι���s\��^{�S��;�h��8��qhlI��[�˦i~T{��nƪ}R��᧞{��g��C{]�CD2�7O���5�n�6�����OTs��j�Hw}y"+5�$a���:�,��;��Xƃ)�l*/�����h�|��p��jDM�CON`q�ź�c�'H��l������^K�|/r��mI���W��eb��g��;���.���bR!?E�M>������Z�cT\P�ݧbu2��إ� *�=����٭Q�+*s-�Ʋ�mvy#��^��b]~Y!u���ё6d=� ܪC�S]R̺I��¾gMZo��o1�x���%K$�xYŴ�eP[l�V�|/�����)�ﲥx�ż�w)#?����2ft��U��U��*�(>[�t;����5y_�� b���_��1�,��ҵM��tej0(H���M�{�Sz�0!b�c��k���f�U���X�׋¹?*�m!������|wWbe��כN�b�P�����#�r�F�7�yÝu�(�WWl3=v#zL�}�����ٲ9����<�͎6D!�-r#�V�Ǜn��R*�)N*����4��3^�O�" m�CQ�r��3�~-.AɭQ��f��Hߙq��֣��*�#�d���-��t��ۭ͔ћN¹x2�8mK��M���D�R<��ĸx]^��>���vO�ǻ(9;�
ΐy��g��bzbmLmGK�d�2�Eo������2�������g�~Ya������5�<����匉Up�3ɯ4�hK�e@��T�YgX��!�-M~�f��I���_jڸ������y�N!}"��[C��k8�oz�_�(I�&C���k��������ݹJ@�f����kÞp�7ͼzޟ�&..�_[�n��GHe��Pq���xg��Ȫ�0;2;N6��hdea�}}����4זq}�U���=#��P�eW;�O��Fu��[$�y?}���;��
Z�1hW�'D�R�r�[�w����?�p��t�ʛ��x�y���"�)LV��G5�=}��vG��Z���R!o{[�t��{)�/���YM��Z����R�T�����yz��3F,��n�Qn)O�����)E�G&��uJ�\���6�aI�	.������eW?�ʶh�)�L�>j4��y���9{���n�軸W�ʯ'z:GZ
$��J*V۩F��̀�V�vQv%�C[�-}1G[���t��WBs��ajYCq�A�	d�s{U�,��n�7s�܆��,.��mCl4�\cַ��ee�Kd�l���0 �L�s���5S51Gǭ�U�l�}4�0SEg�Ejۯ>�K:7V�n֙�z�.�4��I�ʺ[<o�Aݡ�n
k�-�|�x-ax�38����l�F����l�uet�y�u���y�ق4�`KC�f���;B:Y��{z˰�ݹ)��@l��Y�9��Ss��S;b�z�DHf��`�8Di�ӳ�*g��LW�R��M���)���pR_)59+�o��x;孭})?z��m慎r+lb�R�� Nu�>a���cD�a�>�CjT�n�y�f�4������p�V���\t��!�3����RJy���Ӓ�p?��fN�f���z�:��`�����G�ʜJ��,I���K,g��3�pv�N����yuŨ蓹��l_e�սԌ�!�����vA؞~�tF2���]֮��ʶ)�s��uY9�����֓�;�Npw�@q�7�ч]5�Ӝ����e�P�;��{���2�H�vڽڮ|f������?��}��AH�0�&��U��|QS���"k� ���q���<
�a�۪�=p�k�䄩I����Z�m� ��<N��Y7{�Soy"3H�~Ԗ
 �^�%�Cq�B�<�2�Fwv*��7옚UB�t����'$#�'J��X���ݭ�����߷�P��c�Bh����R�Lt�	�����HWن[��	���*o.����V�1��������3)�qǛ��O���Wbm����y�qu�euz�ݠ��A�e>��C]�,�)�l�x�mMN�=97x_Q��W��`�X��Y!]�򫆫cx�6:�"�Kw�ha�k�q��a$�r���7L��~�\X�^�%��^[Cl���,�o���L���P�<$�dT�͟+�
v��zFy_�ʹ}V��yՂV_r������v�C5!��]��/i09�_u���Ϫ[~e�skli"qC��~i�(�E��V���3V��5m?LuCei&����N�)�P����,ћ�P�H�O'(���@1�2@�K�������A�#��9��[��]�0���=ҵpQ��i�6ho���	�u����8���s�����
 v�}�ڣq����̘�n�����q�g��ye�`b�#�l�ᷘ!�o�BuMV�sw��z���*��gb�Zz*�\o?�o�ť�*���2�Uv��ū��O���3���m�=�C�[O��(����q����Y�}�˴7Y5s�H�f����<�h��$�Rƃ.���;8��pÎg�g=p��_�?�Sn�X�c�י��H���48����ã3���]��be���Q�	Sf�_8�����& z������W�4�;��l �.<��rm���Ãf���2jUik�zZ���/0����k7)�`�9������ΫC3�,������J_I^�����]��r��y�ùVNR���V6h������(^�:�tF��x��.�@p��1(��N� EG���w;-�Á��zFDwL�W6H���vƚ3����q ����f��M.Ǐ,�x�j2��KܛB��Z:hEn�M��p렄vy�.��)
㰛X�ܟ-�x���w��ˣ4՚v���h���������F*�6����ЖP*R�Z��q�TU�=��I�5vދ=w�7�pz�`}�*��t�~��v�]��Q3٨%Z�ZyK�I��h��D�[��=@�W�]Hg����7�+T{3y�}��:�5Y��߉޽r6�1"V�I_R��wU��e�k�ٯ9��e�{U
uR��I�MsVn�u߹����v��\�D���8n�e��BO7�_�������g,mlc�gn�������s7�x�u��]ւ�BZ�6n���eҞ8�>Z��u
����jm�1UI�����*�7Mr��\#="�[G������e����L�E?ܘܮ�b�PM��p��uv
G=YI�;�W(�#�����[�$�F��6��J���̬�Nv$�vn���ꏐŨ�o:)ԳM�h�"��������v�RJ��>W�r�̾���,�܇���;=��C�S6*��
���Rv9W�mշ�Cx�p�6�Lu�+$E�yz�o�1�=�������K��֘Oan�����1*Db3a�9�{����z���]��gG��7�ݼ\�aU0ܒ}9����t�G"�`��v�zѼ�olϷx��Ffkqb��!b
����ؤ�_�j
�|�FI���{�����U-F^{y���ϊ��<�S�@�j��`�W�f��a�p��yR�-O�L��H(����m�F���-eS�*�@���Z�����cF��fCܫ�+b�@�Բ���TI��Y9Id�4�D��^��WQ�۝Ǭ!d�}�y�e+F4%�NoC�*����ʦ�5�^��9{���&j�E��L�3�;F�I�^�c��S纒�W
�:�Q#Ge��w7��2���۲Ӽrk���+ȓ�S�̇I��� ��~�T�0*b*�:d<����_
�w{[tOs��j3j�V*������6�lڝ��I'��^��I0�"�o��\0�U������t�B����x��Y	�3,���:W�`��1+��mV��Κ�Sr���]�]���|�^�d/�K�S]t�^�H�	���,�ٹ٢��|ϐ-)��+m�@����\���+x�B�ZW@>� ���� l���R:"&�ϭ/]x8!:��4��@���*����(�U⫸�<�2�-f���1�grr38�X�(0+��D�AF���4�"���&�j�h��	�`�	��uq<4�������hv+�;Q������OJ����NFG]FDm`��-wl�Mh���|fvG~���q�y�:0릯�c���Ge�wٛ�j�ЍZ��e�v�Z і2ϸa��2O�� �	əZ[v�f�����h�w��us`!���Nka��Q���8eH��Α��n�a��&���ެ���Q����W!BT .�D�抖�af��r�xwU�:bY�6c^y������u���2t���Is�B!��f�~ؖőn���'�5a�LγP4�-z�ܚzh�V��[��G[���Jʶif�C�*P�'󛼌��
;��Ĥ��w��}BΣ���b��H�c�Z��:��\��ov�����S���_r�Ӿ��(J\��[�}��b�t�"����B�7�MMm6����
q�l=���_�����}]��5�Q�N��R�J詇澵ѱ�N� l�0�j�v�ላ����<Q\��We+��;��f�t����6oW`��*�[�k^��L������P�;�JH߱o�ifd�T�5lfZĜ��!5��\i��N�u1:�DQ�"洦���\{g�y.���W�����ׇ�Tn��5��/�z�Rʎ�i�5śy-�K�h7�-�F��]����;�H��5�����. wY>�[Րc�\�}#��t-WL�r	��M��Swd?��Nj�7�>ù]�hɃ�S��<n!N�G	�����'[���,�N!-���ޗm��������\&�w2;���㝉�M����*�(���K@=;� �`�cG�z��yt��U\�=��ՉjW��1��An�J���)�#b	�C{�Z�� ��T�bsj�e
ɝ����0��{R1^�tY�'>��u:�fls����]]s�'׹{�Ep���^o
\�4��~[�V9E��A�C{���S�ज�����+yg/����GG��q�0zv������2�*k�u���ɑ�d��jE�&Fv�?Y��kI=bGq��=1��ή[|��u����{>�O�p�QR,_G7���_�s])��C�b�
������.�nU�Gd��v}_t��Q���ț7}�w1IM�ڄ�lǪ=�#�d ���B�v���v[���Bk��I���y�U�x�)�t�Wf�|Ov�[6�1W쀪�'��C�D4ܯ�����	�X���ί�����8����Y-[CV|і����Q�.����Y�YV�tEωzXd>�+zR���K��k�u����6��_lJ��,�����5!�:Z�[Y�@�/�O<VT��{u�@[n�;|��u{��M���=��ߋy<�?�+��f�wgü�>o/w�������}>>�p���{=c�m�:`�P���R��N�~}Σ�e��z/\�7sudk�֋J]�����j3Wʂ�٪�ҕb;\ۀ�\�rU��]ڇ4P��6�c�ܾ&�7��
�o;'�7x)��ap���&�vD��r��n9�Y)IS{U�+���F�Hi��pKIyʒǩ��hR�Җ�Y89��R��*A[ܫ>�7MNU���`�E�P���Mޢ{��Vi´Y�[B�a�����^�^������*�������9Բ���5}�C.�De�GEt�BL��W��+�b�NJs�7E@I�SY�u��`��%X�<�����f7����@����5���*ZϧU�W1V�έ�Ӡ�3�.of9?�tj�i5V�:�6�#!*��=�l��+�f�q�LP�l�@SO��qά�O^o1Q�;P������p��md�R�*�ɍN�ܢ]�B즻 �̜�iq��b�q�ӣ���}V6�W^�z�ݗQ��x�^��܎`)�Z������e��
P�[J�39.�L>��A�XWΥ�"p�Ịtd^��7	:���uMDXA�":D�h7b�e8���>Os������J>\rS�Դ3�޽�Sy���e9"�y/~�6Z���HI��i���R���!�������*�e��]t���!Z�p�;n��1�X�`���ҍiLmK{�g���Y�^�<�����[+Ps�KX�y��A��z�A��ßm�+�e5Q������.��G�����i���adT绩gt��4v�5C�`�wu9�&`��0P�OMO��P&7kq�׺{�V�8�]{��#No-���}����զ���f6�M���}3V���w(�5ua5z�B�S�/�d۾	�\����醔�ƙS�KC��y ��Izs��w3Zx�
,�E�8ǶRC_l�߹t�g�UM� Y�b13R�/3p�8"Z�}�F�/C�ǽC���n�/vCQc�(+�Epx�(num�cx��a�2�-o"<����0��2dM�W˳2��q�i쮱WS Di9��s�CdҩRڗ�(�v�;[�t��r��;\;l]�w`��6[��I
��}��40j���;w���ձ�${��([AFM�V��ׁ�R��׋C|�����2V����a�F.�0ň1m3}�Is���NX#��T6���{=��R�r�k\�9���:�C6�;�~t,t������
��̻;��IO^_ꔚd"x�+R��V�y��>�1>޽|:'I�_t�e�5	Y������4��P���YS>#i�x��ҵs��&v�VM�r����S7�޹��5F/��AI �5`̬���M�u��ׯs�of�u�|4ܝ�݌��e��ss3�ζ@�w�K�Hn�[�b���������ϊ���m���m��*"<�MuF�햆�X)�h����K��E�v!�h��&�	ѭ�lX�b�i���j�!Ѧ�-������������N�#Z�Ҕ���h^�Ev�[�%n�S@M�6^إ�lb�
+�7a�t�{(���t9�4�m�LSTATRV�m���c�BvƂ��wf���4�:���m�]��&�O����]:���U���K`֖�k���T��);Y�4�cG]WF���I�4�-�U4h�i�ڴ�Q���h�m�]�AE�Q](:M�:6Ν9ՓQ5�5ݎ�A֎�؍�lm��8{��ZT�٢*t֞�����;`�*���F��z:M��F�ݻlhѪ����(z�hi郰����ٜd<0�*����7�4�N����~��+e�k����.���n�gw9224�L��́O��N����.�x�h`�n��GfU�7�{��@T�r�i��ךT��xܩJ��~�4H�HѢ�0j�J����V(�E��kgܜR��(Q]�3�koI�h�[۟�%|��:��f8l
�<j��n���^�-�a�+���KvVVq�l�a�zv; o^�ז��~_���cK�S^Y|�m�)�:���[���φ&͐�2u���c�wK3�l�Ɏ��U靋�޻�h�uri&3���L�(dV��n���s�
�6��2Iͬ�0t�{��e�����7�p q{����b�jPl���-���>�FD�}y�F-�}�F2����P�����~G�^G^d�)���{���2g���Ȫ2M!ҫ��E9�>��mﾜz٪���k�J�y�|������Q	�Etxw~��;����N"��5|�����1��zt�r
�h��X��]M¯�G5�n��(#&j�b�9"&�iU�:���˽L�{E�����[�9D��j�3J���� ��1�'+L�aC�ٲ�`GoX�����4����/7�ve3�����σ��-_����
�_9�[oK|�"c�>Kko-.C]0�uʑ�w�<2t�Oj�{"�8Yý��]͇����5�Nsp3m܃ۀݓ>z�����䳀�7�\�$"�4u����O��udi�Ǔ���q�5��!r���Op��9#;'.�SVX�2n���U�Dg*�'2�(V���u%��k�	
�S�:���|&�J�޻墍�fv_i�>��8x�7+uǟڟ6d)�}-E3�ыݏ��!��x�g�����2EW��=<��d<Y�U�3��I׆�Yq��y�87{9�l��"0"�V�k�o)Ҹ�.���x��@s��)�k�=E�y��m�nl�V���W��0Kr�9m*��0�F�+�yrf�X�s�orMe,���!��mx�_�h��tH���5^�Em��A�S�Pl|m9El�k������,2u��{�͂Chv��.�ޕ����X:�j����d�ܜ�{]ܭz�6H
gx����q�5ۚߏu|���?7V-�����JLzE�0Y}��rѶl�5���-讜�XflU� � ��.��xZ�ia��7{k�4�(3�ةa�ե�.q[����a]��W�*͒XCgZ6u!�A܅��pW�>ΧGs�і�5�45��V�u==(,cV>���Ruxn�]S�{Y�ñ�j	ܭ^V���)�{r����ph����l�^9��2xa�c�ϖ�G���儤p���(馢����e�����d?)2�����ñL�<挍!l���CM�z(��=�2j���[��I!��4!*�B�.����Y�Tؕ��D1�0V���m�)�����ᇉ�^@D�O�|3��̚�Ȧ~���+uⱚ<M4t5�s��T���GLLN�ķ
�]�+���f��CՌ}��8�� wW��?Cm4���7CM+�C��vnz�ض��i��Of��\���-��{,9����x1�{����*���q���$7�p~�Z"�G>�Y�p���:�h�x�bj�Lz2�"���\��;+��Y'��f	��{ɳ�2�P]+v�\��垖b�=�g��S<���g����.�Z�,՛�WEXO'8{40���j����l�3�l�7*ݵ() #���>���͸�*����sk.���u'��[�y��e��&�y�+-��\ٕ���-�]���*�s��]a���;�S�m���%>�	^	t��)R3P��֏����wx���9�P�V��Cw��>�s�mwڶ��K�Z��W����Qs25_l�G����M�Z^4�a�t��:��l�e�F������U�]�&��U�]��+&�E8��,��o4q��N��Hǆ!M�����6N�M�r&L���M�DDW���me W5ϩ	����7�5���h����� R0��	�gm�>T�@V���Փ���i�n �����x�،v���D���ZSN)���.��V����������~�it�M�;�%���}ɋH�ʪ�#�q���L�������ͽ������u�2��7�;&�"��Rc,��IPt���M�S~����T �:�f��f+6O,�@�6G!Kw�b;#<Pr�5�1���.<�r��:]]#l����@Zd��qy�����8|�XU��K����[�m��wGeWfo�w����u��Zc�"���2T��etg+=[�hTF�=��vS�m�)�h��@V��w���\!�r�X2S�w���m�� U�� ����_Z��8y�2��E�V�P��r��| ���b��0[ˮ���1�n� �^�{��6��ТI0/� BAd}=>��}]�_Z�N�y]�õ�CI����-��6-K凮�f��y���}����	���zN���k
����GcUw�wpx�<D�$	�3����os��5���+��m�	޲��gzh[�Rޭ����U������>`t<�{��A�۫Q�#zYlg������ɵ`�ԕv�%�����fX-�pԭ�k;��*�jj�]���S��.�8�T�l�n˟���v,/�Oq��3���i�f�BQ��:ٝ��<S����nT�5���o�͖q^xy ���Z�+�^��`;!������]�_nu��I�k�-�a���=��{:�[�2=�}t�<	5��)�SyFC����Y~��֭��,~��!���{����i�IeO�h2�����1��d@Xf����<�N�;�u��?�,�_��+�[��X�ߵ��sLQ��WS�Cr���E[8�Wǜ��v�J�*���y�
=�{�%�e����ʡЬM�cemN�t<����T�(k��r���}	�|��P�f��H��%e����o��ԔI!���W���W?"����i�gF:�zV�x�	�nkNǬ���ƴ��,�l6)x��_=C(�OG$��Z	�O���(��S����3��1>H��Lڀ�K�1;+�ʑ1;��t��;}����B���D��I�m?@��P(d!m��x%N���.��=<�<3�e�$���|�j��KTJ�n�*��8��<E�q�E��O��]Q1tGvL����S����er�kz|{e�3�z&n�1s�ڮ��\��y�^J� �e��ƚk�4
�^a�i�~���Q��*"�'I*a(��9W �-���1�ڑ��>g�o'Dwn�j��7_"@�@���4O��K���~d*��3�u��9K^[�w��?p��/Y7� ���Ϥh����\xEu����>�Uq�V*i��ѤU��6��Eѕ�V��e�K�҅��h<�^���\����C��KkOMW�aN�\��RX�](�h���^�u�`<2VF�F!	�Y��YQ^�V�q��	�d���s����ɺ��	�nl�/:\�C�<���%�Ħ��W����5���a�+�|dC��\f�`������KJ��ǵ��vDdN�gO�Zn�n>��5Ό��;����ʮ��5���շ��h���#�]i�n����E��Y���ϻX7@6�����(���s;���������n�7\ue<�*gg��O{L��2c^��C�Ξ\�;��"x�9%8u4�Y:n�w�� �c��1���͈�vUVvJ�͸����M\�1��Y=�[���=�Δ��w,߲�t+q�~!Ku����^bmLM�`ʻ1{���$��!@����5�ѝܵ�i���}�Z�q ��`�*��]�z��H�%�ї~�3�NH��UϞu���KK�ߝ��3@&�CY�8
��ܙ�^/5�<���f`��l��x�ҳ�TU�wP[l���jzE����>��ge�̈�K����9�_r=�(^m�.V�t]���P
�6��P����yut��Y��=�� <v�{�:<q���gh���ۦZY}Z��7{3CU1��i���T�t��v�7�vC�$r��-����,7��v`�	K�wh�ͦ����b��mP�I��]V�����e>�������ao�h�,U|1��J��g�u��A�i�^~���IK��WU~�W1P������N��a���jf�w �ռ[JG��(�fn���&��7��/$��l-Yy|f���Sg��v���� Y���J��(!b�*i��ڰ�[pk�n���<M� �f�ݩ��a����/N�0?�J���m㾨�Q[����;�O��M����0C-����r�]���zwy�c�o�i�z�w�+�R�2	ݵi����^�A������[�Mgq�T�VL���s5�Y�(�ϩ	�cy\�geAp��S�"q��Q9Z����6=j�-*�c�|�D䶓���c6�qj��'V�vx��D٬6�L>٘
�ؾ�z�x?a���>=X)��p���0������m���E���g���.���xϝ�*l���%�le�Mfخ���s���H��[PJ��]]}P�_i�{�wӃ�t�E���Y�"��-���}ַӥ�3�.��gI��p�����F��*.h�Zݥr��<[g����׶b�h���Ϊ�j��j�����ߘ��f\��r�!a�T�ћ��^�ive���W�Ż��#�&F�g�����m{�Y��^:�=��'S#Z��I�{=�����3���y$6G)�T�}E�l�邱|�"�VV4���{�]�aeM\���6�49-R�gm��O����g����MQ��)cNij�A�$��г��(.#���e��]tY�TI�v��{Ml���xg ��j�����i-W�J/^��K��R��]C��ks63y�����I�U�m�E��G��Z�0�s��5˻�"�'�'uf�gT_�um�E�Vm����5U_oU�w�T��{�i���,�՞'�6�N��|�@����5�Q�o�w�߽�.>~c�0oΩ����ؖ�Q������0� �0oYP�oq��t�eW���#�έ,����˰ڔS4���d�F��ep�a��H�+E/�^T%��iPSk@�[���I��wrg���ES�ya.����I�L]�]U1Y��YJdn��O�oI�w������w�ܙ�G5��յʑo��5��F��=l��z�d��{�9�����n���L;;�d�v��\�h����Na&���m̆�]8�S�N_������ܸ�<+"���hLe�&�Y�D��Y靁���7qYgX��D�&�D��ݞs��V� j���֦7�n�L�9�_l�ʇ�;�ԮA�Vl�Ыk��rgLL>y��j�gd�dw��v]���@Xg�m��ӫo���ݵ}ӼU��?m��5�NOlϪk�1������4]�[&�yi�,^f'�ی�Ξ� ��Ӎ���N�"��H�6|��#��ώ,��D�ٳ�x�����.�Y�/#w�JDd�!YT�|���^TMNZ�Xe��!�q�*�s�wSJ�N��!<���	El]LGC��<���7.�S:-{!��<�P{����Q1�f�m2���̨J���Ҽ�sE�l�����W�KYM������d���� L�������yz}>�O�������G��5�$�k�1���"u����1i;[|�4Jm��E�.������V'i#ͻ�&��i��[�yZ��@�KȺ�K��r���z�@ۀ�A�6���Sѽ6�<6mn;��Z�Vh����t�7e,��P VMBFe��6lFV��h���d�!��C^1���#0X�</�,&��ܭ�m�ɰ_��cj�ݩe��H�n� y[Ư�vuN��ڇ5�5E�T+:T�k�hb��6z��2���w�.M�U���hַ�Ӿ��SYAI�,�V��Ës�Y[+w�.�����n�v:-�5�|Vv��(b�=�5p���u7���٭�i�m�y�H��7{�+RZ¿��Z�BR�쎭����F�-��K9I���'���0�	]^_Y��RX�`y݂E�O-�q�:��G*b�����۬\�ܖJAۚ�C_ljd�IK ��G3�f5ټ��C5'TB������7M�%]՚��jZ�)����	�̎�hGΓ+	M�G=uoz�k�K�,"m�:�Ue�Ӫd�wR���S��5v�@��j��C��$@��Yǯ��x]acy�ZP\�����PT8W(v�������M[w I��t=,i�}���]kٜ;VL�C�`<� �<�lwI;�����T+0+��1�ͳHJO�+R����3�첳kM�s�c�xo���x���̓'>��S�h��g���YBA��j��0l|�Q�OS7�;`a��j�䮸��`G���b{�3��ۧ�>�]F�����&8(d�؆�uf�ǲ�� :��y�v8�H�+z%���m�ŕ����y��Iukt��L���R�LoL9$麴h�2�+D����U�
]�,�}��/f��я6���o���Mf.}�:��k�Y�
H�T���:�oQV�Vr�f'R0��u�SЛ�AX�������
x��VeGt���Y�n	M����k�ek��H��Jvs��h�J�Z�#�v$+���E�oVŻ�ۦĎ֭�J�wo"��fCҒ�ڷs-g)t��/�_RH�Vpx8Z�sM���=���$���_M5ɻ�:�+mc��;­^�L��{@cy��b�Z�w<���꽾˚��i,f���;!�̽�tm[��7)�1��ŀ:5��*_e�坕�ҩ6WJ.��x��Q�7P�݊jb��K�6��/�ݻ��5vȡ��h"z�2^�fe����b<.�z���Ȥ�v*�Uի/1�rݣux��ubc%�x^����{z��e*u�5��39�6��	m������;,���ti�}i��=�#j��※�7�|�"���*#��&uy�K��ֶ-䶆�������b�`U�����Jй�p�{�TB�/5�!�҆I;��9�;���c�D��̱�PhE�h���hu<bd>Ev'f��Ύ ��l� �rRn����y׃����������&�W�,�zWV����@
 H6�AMT���i�m�������5�ִ���Dkl*gI��k����k�V�Ŷ�b�Ţ��ѭ�b-�;mQ[gkn�J�Mb13/F����q�$ձlH�tb�kQ�!ƵEF�4M�Pn�AWmNű�S�4X؍[��5M���IBc:�m��A�v^.6��N���ŰUh�M4��QE�Z�n,[c����&��+E[kU�Gls�T[&���j���l��3W`�fۮ���G�����bJ���hE-����n*���f�

4c���A���5�1kq�c���:JI�S�ѣT��:��(ŧѤ��F��UG[Z�4Uw`�����*Z��"ZɭkX�:��S[j5�Z��)���E����F�X�-lb�F0lgh��ڭ�gl����W��I;��o���$̤N�kj_U��_g���ܙ�K�4p��4��;#z��&����厥����N�$DŶt��N���}?��+꤭����N�ty[c�iaU{���7Xg7,ĝ��j38�:�'@c��]�Uɺ[Al�wf[1��'��;W*����J����!�ۃ[г]���o�-��l#���+æ��\�qJ��$��ݴ{m���CQgdGR/%_Km_.�\h�%`?nSԋ]���i̬�ƪ%��e�; ��8dC��\g��v�ʾ%��i!P�]��Mf�F�&ލ�3�2�T{�1� EU��t�o4��O8��7ƾ��������Q�R:�&�n�Nt�km�����+�Gj<�Z
��lnm�-��G��i}=:I̿q�v�ι[?w�����0��!p�T��Ҷ�(f1�"l��8��ܽ����MA�!��3�=]ܻ`��(몇}�Yjl�<'{��x]w��U)��U��Ozw{��p5͞Ё�J��a���X�Yj(_�c\�WRڴ��)̰����Y�+.c���С�������Z+��a��`VnhFE�W�۝�Ju������F�p�N���_�N�̛��%\ �7v�}���[��mmq�O���:�b���鼯�O�6l���i����T0c����ܑ�]����v���}=t�ژ��{jl�Φ�>���u"&����F�w[E���UN�t�mq��q>ւkxo'�����k2�y��f����#e2�m����^���)q; _A
Z3�;��!��eLt����r���;p��Ҷ[�!�H6b�v@ێ��U咶����1�ʽ�n�/Ռ�J4%]7�;unF$g:D$2E�zզ��I�s��%.W�U���i�Ҹ���OCӽD��Z��8�H��|,��o��H�:2��t�M��U���(u"jiZGp��kƦw�VLp]"���f���#o� o`�f�t��̮�掲8�mx�S�Y��x7Q/&���7�˼U�۸�(Z���,����up��]ة� :���@o{l{�M��bI�Ƙ�������ոv�f��pU�iZ��@� "/�,�1�h��?���GF�ddN��p�C��c��5\�b"ކ���S{*�g�u���[a���|0G�����z�]6�a�!�kOs)�j�]O�ϝ��ݘS*Din�X��E�K� V6K�Cq���:��D�)��wY�W]9�'�,c>'ue�c����5|r3rr�D{cei���^*Q�}1LGC�wW��-(�u!:c,o+���zv���;r\:}�C�ӷ1�ѷ�ʇ՝�~W\rX�����hw�C��a�8��]\ǏHh>�ژmy���fDfE��[��{K�W�]�ءǅP��š��H@�2�4�|ݗ�E�а���.yMM�FśJ&�<�s��UM��ov���)�#l��� g�]������jd��f9��v�2Ml�x�D���uB��4ө�l21,�]�\2�5�\=t��/]s�[T�{R�؆��Kh%�������ћ��b٦"o�'$;~M�7e=�]"����J��T��N-gle�m1��b3�D�Y��x�l��UrS\�����q��)n7���E�7u>�n����@�1|���n_�|�~�����a������vT�k(�rd8FL��	�=�,��kǹ�x�$۳|:1mu����"v���I��ʓn>��_]�_T��],��B��G�y`J�M��r�E>畺u�׏�Pw܊�)/����]����GWe[w^�X�JW�>�iR��i�DR[Y���D�;oa�mO����`1;*�&���*�]����8��g� ������@��)Y�qbs*�V�2�"��o#^��j�픕��W���υ�c�r�qZ�ox͑�oc�\uU����B|&��E������ fc2�g���љ�f�杹�9R"�Ll�26�D��%ܭ�u��6�-�U�^9!��Y^��Ǡ9�1�L�2q}����|pWa�%k{O��W:!�)1I"6��M����}�p{�fc�ȹM�w+�y�R����f苽��\����A��h7H��j�X]�#^ʇ�!y[��`���Ƚ��5c��Yή��Esq:@s&@n��v9�{/̛��lq�Q�5F�W}���H���}�������j �Q�c��Yo�%�{�&i���`���ᕍ�K2꣰H��&�l�'���}�GTrrN��ԉ3]>c�sF���Ws��V�"�m_�Pb��_�s��a���Ա_u֮7�f��7�^�-+ĳ��=��u�������ޗ����\�9�C>�T��v:�g��3�>φg��Uo��̖�-�h��|�*U�X�WQB��D�}:�V��R�j����Q��.��WX�H	�.]Ի�ٌ���r�1N��wYs��`���?���Pk��wʔ�������lA7��v���v)��J���W��<H�w�5�%s���"_�gh��ٽ�p};�$�8�A�����eVRY�I[@��Q��稳e�.VavջoK��w���x��G,{�Mg���F���֧�����}��uU?�A�L �o�o
�p�)��z��v+��{�t5�w[U3�tW���A��i��3`��/�_{��z�͐�W�j���0����|�r]6��d�Θu�.3q�6�0Wc;�en���<��c�Z�����r���M������pmL!�>r�����򸳿$�lٰ��r��S��W�>�3z@ݍ�WO�|^+�Y�,	��T�v�aq+V8*��Q��]LӔ|�m���3Fj��WNC-]OoqT]2�!\�w^K��l�H����#���4A�n\�Y5/Od��7%̛�M��;�ૻ�g��c1W�Hﱉֶ���ga��,W)kmS] e��m)��u�O�=��e���k�$3��߻�p|c9��pw���ni�u��'@��m��`R�5���^�(i�i�Ӕ і2��5D�^:��)�����KZwVl@�B����#���ƃ�n�m�x������=��1UU:9S޻aA���<�B� D�*��vb���oJI#vxN�tS����E���㩵3�C��<MR+ܼ�{��qB�I����z'��FG��&�c4ynv�nr��=��*D������n�;2��ʎ�Y�!:��V���o���`�cU	'�y�p��y-��hi�~O�
�g(�P2�)��R4IU�Y����2�j�����K����.1��lQ�ų,��M?A��]���jrǯ���}��LKE�fS��w��<<T֑H�ЛH������g'4�%�k�2c����; �:�o_Ě*�R$'���c�n�57�5}=9���p�ʜbh�~{~��v��.9���7,��|Jf[]��Nmh���	t�S���k���]G��%:v���Q?��f�W�Tv�
}�ɂ�l�{ū��c��l�Fn�P��ا̬ը�ͣ5o=�ܖ���qf���ʙ�ȦF��oA|�Ԃ5��3�{����Nx��و�/%k���]���f��X����X�[���S⻊�]ة�͘#�e�n�|�]����d��1G��;��];h��I�J���幈ǆ!M���?�{$j�����͎7������ۄ����s��|.~�D���Y�ʥ��;��ޠp�J����@j�$�/�\��Ocv��q�k��և�Ȗ1i���w=��EE��Ss fHc ^�u;��\+9b�/V�۴G:UU����Y��h^8��5bi�=bx��cA�����x��b��m��Ց|�Ci�9�<�b����;y�=���SX�c�=.�톰g��I�8Jj��x�nx� �&�γ~q"�e�\g6�D.kԪ�|��/�����-Ok��][�̤<��g˳_N���'ݍ��ul���-����~�,��W`���#�KW��v�\�-��k��hQv�Ǫ���E�
ח�5�DE�R7C7�붸��y���w��"���bFbJ(���b�m2�2ק�Q�{��Y���N���p/=�%4�{Tm��8��VNP]��a�rUl��]�9�{,�,z���B��|��SE�0���J߬�Έy���u�j�d�뛕e,ʠv��P��P��>��*X[_���/�rm����i�p����>&N׬���v���^2��Y����l�9�.z*�����D�q��yZTw�ܕ�]G�{��x�Hg�r�#$߯ 9�X�O�N$����P]�~ผy�K�vG�W�g�Hn���f�h�R�tN�Zӄse8j&�LV1�}̙�PYv��Q�U�q4(>V����N��C�0�-\]��w�Ll�Uk�x�)+�v*�az�d1]n�gNA*rh�D���}]���k�<n#i0V*�F�Wsx��>�' -L��Z�Qә���{Ȏ���������KI�~��B�J��u'�~�r��ŝu{�$�C��u/�!��y�y�ϳz�Ay�&����{ñ�ɛ����C�|]i��/W^�df�v���N��E�}�=L�)}��0.w,9^�t��Po���,�Vۛ�����E�w�a�#ͼ���:�����ʘ�5��|L�d��q%�Vȣ��v@&���k����YU����;~�o��.�ើ+ _�~�x��=r=��U���|�0�,�4��B��_�/L�b*�BZk�0ǆ������q�^$X�JX�'b�4�p�����ڲ�� bM�V��&�\�/ܳ2L���!"2t�bGm'��lɸ��ĸC�C1�4�>��x�jS�7�br����J:��Pf�3י�z-1ވx�ʼl��u��m�:Z̽8b�^���'L\I���pp�V�Y/q�w�@'AT�	8���	d��(��v�G�BOU���M��l67���aH׶cv{,Ke\�Bʬ��*�%�7�{!�a����C;a��t5g9l��`�E�8qXtL���
=�A�X��B `�W��2��msf�M�q}gTN�VG��
?�q�U�_� o��j\}~���#�6w:��� �������/��H$EB�yOMӾΈZ�#��z�oR�t��i�Շ#/2f�H�SS�W݇�D�"��k\>s��f�sT.
�>��=����r�{y�j�"�gG�s\���[��.�ܗ/'v��]
o�����8�?-�/���y��|d���N�sY���H�[����v�>���=�$��c��ۋ���H�� ��x^S��v\뎋��m�WWY�a�Ֆʻ�7i���\���;���!-|;���dBޑQw������gu��{'x�Ⰵ�UfV����X���r�g�~�2� v&�{�-r&4� *G �q#OZ�ya�[F�M�����y/�t���ԬU��5$p�c�q�dRIW���\�״�6᭎�lG���Psb5�����Y��CY�ddq�D��L���tW.����3��*U�*���W�XJ�����;�iןl��؉�U���ަ����+�5K�FEU�G2t�dP�c��K�r��W:M�k�y��?����@]�h
�/������e �<**���q���|����AL��� L�! ̫2�0,ȈC(C"(C(|���fbEì �{�Uì��{� 0�|�'���a `�P\0�0�00�2eEpȠ� �� D@P @ �E �T@�P�A�D � @�  � �UV�P �
� *�0 2��Ȁ���*� 
�  *�2��� ʪ�0�0,���+�2,�0��2,0,2�0,0,0,0��"��*����0����|���|�������"�
�L�*�L�Z>͸_���=�3�Ο���}ϐ8~P�">1����8�O� U�ߧ�v(�"��`V ?��P� ���)���b�8���
�����4&���<~	p����B}��_��?�b��r �+�)(��H H � � �  � ª�J 	( A*�� @  ʪ� JB �   H?�%pʪ���"�0��
"�c��b�������TTQih
�q�����~�A�����Q~�j� *�:���`���{BN�}l����N� �C�"sў�xE � U���������"����	 U�?����|C�x/�?��	�>'���<�V8����� zB���;���
]�!�;��!?ꇀ\d� *�`�� �
�@֡���D&�}�F�D��� �6�d`K�T U�Z��$����&[��ϫ���"��0~��D]��:�����?��e5��� cb]� ?�s2}p$%�.z�-�hV���*B�J���i!��D*%!4h�-f�U)IT��%@�@�����[eDET�U�Q��$"�U4��iV�R
DIM�٪����	V�QZЪ%J*$��T����2��PP��J��%A_YQo\�T��{2)U�h����$RU(�U
��iEeP�5JQ%TR�$J������h�����al�T*T�Q��ڐ��
/  1C�R�;��ڙ�WJ��*���ݲp��+mt�Mڮ�����;k�uv5;:�F1[M����IQU��Y�n�]MA��*�v�u�+L�
�RJ�M@�� 6B�P�v(\���(h�
�S�B���
(^�.�С�CQ�@-^�n9�ݥZ�֓�uZ��r����l��c�*e�Y(J�+��n�R��H��P��T�EE*����  7w�4�)*;�ܖu�-�ڻ�y�WJa�N�q݋7[g)m�Mj7N��n�U3���Z�u�;۶��j�ӭ�����˂T���\�T���ڽ Ė�J��   ���m��ۭ����-�۪�ؕK�
ۥ�iƫ��.\Դ�G��Ҟ��f�����[l֧u�9��O2��Uں���I�ISc	T���v|   N�ݯ�u�We7m�Y�U�V�[Y��7��zk��ڇl�F�U+l��]�K*�:��7]Gf[���V�NJ�Zk�׍�
�ljR�jJ$V�G�  ��� �q�)Թ����]rjkM�M�5u�R�$�M��:z�-�bmk^ѳnv�ح�!�������L�4�ݗ9U�f]�*�%QD�UR"�� c�T���u���Uuk]��ݚ�Gp��ӹ�t�m3�k������U���ֳ�7Vn�(]��6�jB��Uw$T.u�Hm���D�R_  >��J������
 �YE���c��P���}�/M{b�`lP��nR�AK�T��4͞�<=	t�;�\�Pt��nuCYz�f���Z2��[|  1�袂����EN�:wR�"�:���(S{� w��W�"P�9� i���*;9�����g���*m�$��"��  a��-m�]��B�9��T%:�� 'v�h���Kt�JA�4�T�B����A�6:��(�Tg'uER�C��@d�J&@ �{FRR��@�M�*�oE<� )� ���@ j��J�  &�Bx��h �����������Y@oֶ�䧠��'��|]�]y�z�{t��od��@�$�fr���IOd!	$$?��!$�p$�	'�!$IBI	;��k��|��Ux�ᯜ�6w"�ű����e�ҡ1��	�P�U!�V�|~u#��NԼ�
��YW�J��2�Y[�J˔	ۆhj��H�Ԡ����Im`y{$�G��s3����Kr�E��^�� ��LQ�lQ4�y5��L?��Q0��Y1�0��Æ,����;��ے"�^�e�da;¨����([t�^սYz"�Di�Z,�X�o�
X�;2�,��cn��.�ؠ��MX�+vn����D�N�&�	� K �%�*ɦ�u�A��iU��j���hn҄U�X�I�惨D�l6[��,ޛGlٔ��њ�L���6�����B�56��(]��v�mZ6��b�IT���	�2D���\t��m4I9�M��K���f��@&�ǚ�4�.�?��b�Ѫ�e��M�2S͍��1��]ajU�,jc n�N}��P�"Oe�H�`��������Ki"��f�L�˦ue���ڧPV-�Z�%!R�^�Bw�Z�@5s*�6�!�&�
��[��7V+e����/Iw�c4�ӕ�oN
єj�M�4�-��d%I�@���e��O�������Z��r�K3k!�%�{��u7���(0Ģb��Gn���W�u��"��ۏlؕz�����r^�[� rH�h�!&�y��W�j;̛O-ǥG�f�v�^��Ő�a����6���Ș�M6]ǐ�/n;M^+�m8��j�B�=7`M�Q
��ܙ�v�b�)��TSop��ש�
#b�7nB��%	!d��*�wY3H9��Rùk-�Cp�nص�SXX��p���l����oknd�Ro)�Z���]ņͶ*�n��ۗ��ͩ~���U6�ܰ)6��;j���U�����+Ǵ��Œ�۴�w���#/n�5S�?�я:��@E�iE� �JD�v)2��A�
۬Xn��C�i(n�B�7s���D(Ę��%��Y4�s�$�Zh��(�pl���z�أ˧%���`���#I֊�	�T*e�+#&����˶�K��`b�kZ�����Ϥ$U�P���կi�w��ά���Ŗ\�ڈ4jm�b�̦/��I36�,d٘�PJc_H�{��
T[OGB�RÎR����7��w4�qǷM%���U����[U��eFZ1��е�̅�5�w���)����@M[�Y.�Ԏ�7�l]��(�a����n�t?S�lw�1�+bL��]5e��VX�ɿ��Лh�ɹIah���bɨ^LE�b��L��LG(H�Y��z��r�O+%zb��b<cVf�.Ŷ6�B�輦)]�)��ǆ�c���Ҹ�Jݬ�4ci����w�/R�6-���C/{��ה�ZcӒ��+���2��)�F��N�ܩ��Y��@���c�Q��y��&�@jf�:�-�^��)�.�����V6]�vnRv�8�S,7�l���?�4@&� �Z����]������pO��#c��kɒT��Ί�4�bQp��\ek9�v����2��wkVco(�JZw"WrB�u��R� ��v�HRT>e��N���{6%٫H۷)M�mG %Y.e��ݛ�m�
�n��Ԓ�Z�ԣU�,+���R�.]��Q��Wt��VX�]&/-9�K4���5�:�T��3i�(����"8��m�r��Znrb�PC�njc)븤*�Z��t2��Y[WB��wn�#t��uD[|����ݚD�
 IlcvB���,����!��N����&��<����橮�D�L��F�Pt��E/j�$��N�æ�1#x�:2�ef�4�:��Z2��ӡ"��L+�E�Qyq �,ݖA�ׯ1-�btjIYS &��wr���q��xw"�ڼ��e��� S&�4���F<�p�v�"a������F�c�6�ן<�w��iC��Y4��̺��J�)D�B
Ԏ�1BA�.��Ht�u�Cfـ�BX��7P�.��0R����3hR5>v)Z"���%f|7/Nd���XT�0-ŵ.���ٺ*�'U(Ӻ4`��=����QLB��8�nb1���P��Jn[�$7a�c@׋U�x	e-�����.�)YN��8f����ׅ��+jC�(�2=�)P�ѤՅ�c�G �Z���D�Bh+Tj�8�x��]b*WD
"��.�ȦٔY�� ۛ��flM��SS	j5늕�]8J�S�Uܕq�����t�3R�r,2�H˺{Y#�Q��l�lt�,�Z�'V�3[��zBz�]�fQ'Th��˗yT#-|i�VwHv����J���(]2[ke�	|�1|̽�� X��i��fV];�^��P��|Bݮ���K.z���WD�Ř�
Vj���֩�����7e�b��UI�K���[�D���,j;Q�C,וU��/n0����%6]kH�f�,%bPͥ2���/B kݥVWAR*+_Bj�*Ã7�v����H��V��)������<��d�@	�w��j7�᱗��KTYV����*�@=Н@N��V-���E��[Ν�߷��+vV �D.�F�y�(�Y�[�}���=�S3V]�2ʉ嵙��:��%�"��M�pbtm�k2��X��mI;5
����ܣN��k�F�"�i�{�e���,4Ð�\u�t�{��ZKKWY����-[�ԫ�N�:���ӎ�0G.�U,5��]`����w&|7r�\���"�aIM&�M00�˽�e�̿��)l���=�N8�q�2�)�!�se�'b䈰���4��I�MD/����á`�z-F���f*�d45ս�0ݩ�?��4����2~�q;J�u�,�7(���tۃ/^�@�Oh�q�j�QU��e�X���Xkq��-A���43)�Ҧ�����V�]C-	Wb��7Jm���ޖMn_�tKt�v�6����fޓ���e�c�CV�M�J�s,�3.��$��	b�T+a��]�-j���e���-��"Ù,�����偋@j���C�7C��&��I�I���r�����*�N�Q(����[��
>���Ʌ��k*-v�yGU9��B���
�ܷ���a�j��V��(dK�MGq,$���*6�LԶ���^Uѭ��.+�/l
����������QU�t�N�s`,@V4j�U�X{�i�U. `�*6��8��6�[�{��I,Q�4�Z��4`�UZE8�f�(�m3�pKz��B-YJ£���\t!֬]I�y���*%ke�8��(�虸�e�{t�e�p��ۛ���F�T��WV`�F�"�9"!2�Z��)�mc�q��'N�M�n�����I���o!��:l�T�4�.�����ۼ��#�wI�^�3�^�.sM��Jk��ц�$bM ܢ�ZV���5����r����͋5�n��b����5�XWP�
���6hQK�ݦ�BX�R�A��p*��n����i:F�*n����T��H�A�β(J(lʺ��Ā7��65vW^)Z(��� Ĕ��C[���˒#搐uU�Eߌ'N�Л��N]$2�)��%�J��_�	!lM��!�BVK'F\�`X/-�N��H'D��y���Ԟͭ�[�<��xnIlv�L*3b\��<��C	�ݒF�`m@mAke�XHec����݉ch���PO3]��۶�R��V���6� ��Uq+':n�0&2��Y,�mJ��p#{�f�e�#F��U���;Sa��t>T,^&VOM=:!wI�}�=�"�$��6Qy�+��E+1���T.����7s-�n���/JڈԠ5nҙ�wVu�N�1�)�b�+��
��܎i�D�d�8�.Jɏ[Z����՚��N�Si%�.�ԭ���*�S�^�,&)�lB����u���V\9S`��j��*jM�F��Z�WN�ڡ�k����&jp��!���n��J��ͺub�T�U�8u٭�t%%sLkw�6��^Fԭǥ�/x^=����5�L�3%��RR�n�5�Q�"�%���q[(�5�P:¡KhV�U4l'[�(B�-�6�����`��3d"i)0`�SB݋%hv>�6�f��n��٫p;R��p�-˼w�ExP��:�8��.	S%���.�v�Z[u��&��� RH`U�����n��(�3`����Y�tk�0:Ŷ/$Ҭ���`��n�[׃q^.�r�ˑx�-�֬7VО�Ì�*�8 $c�RN�*Uӏw�@��Da��cR��Jސ�c�����.��U��)4܈�5],G4"��z4 �r	j���-�4YŰ��yhD��K�hG��;�,�b�Y�"ֻ�A-Q�)e<z��Ú7#;���>*�X�8ΉR��R��Q�"\,$���zN\���2N�����j�m�n��e�y�`�RdKiZ�V��M5��L[%i!��o]���"]���2 �h���E�X��:B��;�x�.a�n��j6�&0��2��]`2�7T!�&���ӅjB��İ"X�%���q&��v��6�@v�`�@�"�U��飱K�ح��P]4��!�
Y�73��b܁��)Z�?"�^V�÷,]5fq(��;ICt�0D��Ų�P�&CUwn�F�͋D�ʲ0�����;0�-��=�y� ��E�д�,P	`�¾x���M�<���_3�nt�Az楛*f%��v��[�u'6֤�ƃuh�T(6һ���ڙ��5 k˥���+(T�.޻4!/hlbq�n��u�X٨Z�޸�m���J��4|�v� ���� U��3A��:	�r�Cb��=�0��fʓ/�3ɱP�p,Շ.�5V�T�I6�;��ne;��n<�b��ue��Z�,k�o.��V�^�u*��iJ�6�X։x�8�M����}n��:T�����<U�������]h�*ҙM�0����ir�F���ݳ���`�boRN��l�(T�*����sf�^��+5��-��N^jaM��U�2	����Z�%���y$Un�?��N�+�[Hw�e�v@�'B�:��mc����,\W���w�&^�ɭ�0Wn �ꌕ/A�f�)�-�T��X�-@N*cJ�%6h�<�ɂ^ g�s
X
_L	��>�g4���X�����)j���O�Q��j��}p0�B����'#��E��u��r�,y�Q�ĄHi�In��݂X�&���4b���B�b��&^��n��f��z�%���))��t�f��Ee˦�h?�j:T�QU�*�/�WX��]���{Eb�d����MEh�R٥n��78Q�MScrE*�W[�K���ʼ	iF�V��h�DM�2y4d�t�8�Cqn7HLx2I,1�Z��jJԷ��Wq÷�м�gu)jV��L9B���o1�����g]AN�T�K�x��%�b�/5�T��F�U�1������Ա�5�Z�*����5�_Pٙ2��M����٬��v]�ʽ�w�r�8�p;��hH�}q:@��Ţi�јT�bE���E�;"ؿ��-tL�ϒT�^�p�(c7AB�P��弛J^�h�N��+�]hdK�п����*f�P�����)eXc(������ٴZ`����fNF�mX�]�銷XFX���u#u��fҬ�1���
�ڻ�eY��aW�恭۷IS�t):�r�9��+&,V2�J�)X �e�)��h��ca��8+*�{�"�`9�(Z2��GJ�j4Z�Y��f6�dM빂L��ԕ�u�Pi�u�5^�u��A#۳W���b����ĻY�%Ðkct��1��!��E遭חR��ʤ���c�"��ʼ0$�wA��icZ��OM�`�����M�cY-u�κ�ybsF���
�[����Y�jJ�M=�4^�Rb|�H"IM�2T7m����Y�5�,L�i\ĥ�v��J'{'Ѻ5x�F�a&0	u���3����CX����"���lƻGF����0Ҹ���ޒ]��z�3l�<�υ�Lt�Y�jf	B+�,*�yS����F�?1�bܠ�����5�G�`�@�����+7�߉mش���G��H@�5TD��*�=#2m�܀�L�ePĂ� �;q�sޤ��݆ídV�/�/�;�t ۗ�ػm�����-�+a�bB݉z��"Em��� �(�K7��i�� :N�8β�YK>�x��$,�V��TZt�x�CJ�x&� �.�M� �֥\&�m���,���x��Z�k�m=:j�mm��HfiX�Tr�� 
q7WaR�-�@Y����y�RTj!��ˑ"泐��7ʰC6�v!s%b��T����k^����yB���!��%��B�:4��!��I�ܢ�*�a���z�)
uf�n��a_�ӁJ5{�[V$ܸ@�4��f�e=&j�]+j˽(7�pP.��6񊱐i��0����x^�u	�]$��+p,�mb*�jұ9�s_�F�d3Tʷ��m�Kpn|��H���`���ݻ���x���b]If;��=Z���(�b&1v*�}@ʂfSo1�֋�7��|�U_��sK�W�b� 쑄b�-�P�o%֥��:(�x۔��$d�� �֪���F���a��՚��l:8���j����u��^YGqh,I�q3��^"��ʟ,Dn�l"�i��h�2ܽ�e�n�a�.I����.��YT\�Q��Q;g
I��'�wW%<v5�6�&	�����bH6J��/0Q@��G�p
�i��j�d�=D
Q��q���cB��G��pa�L��w�m�Q.k����;|�h�w�i�gecDs�$:�T��īku+�o�W�DyYG.�l���3T踁��/���=鎵r��Ua���(�1N����J�L��c<�=X)���M�-��!ej8G+��R�?�r�s��b00X�*�A'hr�6M�K�`�K*�$B��{G%�����c.:WK���*�h�Ď4�0̬���I�X�-�v�v㖟:Ô���Џ�t�!$�T��p����PZ-`kBOsT�����`�{�V�ќoZ���8S��deTFʘWe��U˧p�s"��F��E�u|�]�4Y9:��iu˖qX�5w7ZF�_]]9�v��m<�=�L�VSo]��{R����g �3���$\���WI�f�$�뻩�\�L������R�@�MՌ}�wv@y�3\
�k�P�K8h��O�Kk�������Ћ�u��v�#i��������.�u���љ\���\
)5�D�;������V���N=��G�ʛ��U6��m�2˒Ҭ��S��
h�v�10���Y29ցЫ@��h�R��b�59۵ϑ�c��M�ò�]4kC�]t`�)0D��f"	���&���a�o�E�S��avǮf�����^���<��BV��\x��³�i��B�_O-q��b[������z�eb�Z��lK%��C�swn�}�B�o��2����;��/�"0u�������2@�yn�
=H�kR�q<�����+!UlϡI��ˮcԜ�ɕi�%>gp��S�S���+�t2�W�c��[��H���Zw,�miE���y9݅���7z�/v�Ȣ}�zoJ��Ry��{�ĝ���zQ��[֙�km��-�-��!l7x��)5��m^(�l�{+Z�1�r�v�^�N\���4��xf�mf�t�Y��nq�hG;{c�Z�)���}՝���x+��:����-u'�(�L�v�A���2h��Y
 _v��UZSU�CE�1d� UĎ�z��_Q��<
�;�����3�%�3x؝����ja�sek�9��7t�Ǌ�s޹�xwp��1� 3��u}�Hժ�HuH�H
�ӝC�v�	�YH�=�ܱX}��K����u܆28��T&��;D��r76��л����vt�=l��uڭ^�y�9P],U��-��	P�.2��9��&�x�t��p|��=�N!������_n���R=��O��w���"��MLi][��&�O��(TKi ��2��ݨQ�7C�ow�$���8�Q�83Y��H�*�_f�]Nb����=�	4pok�S�s��7��s{$_Y�i' ɷ6l��9�^�W��W�z�@(�n��e��\�Z��c������\X�M׃nV�tu3��V7��jh�<7�K�Rk��d�
��9�Kt�n�Ɛ�nL�/^���NI��zx�.L�0��P�cJ+P��{��2P�ON�m��I*[\��-���u�e�}��cٶ誜�;\ݵ*�j��Oj�ě\��+��up;�/�x��;�,+3u�7�%�M�t�\�n��H%zWu��],����9���ds.�ig_�0�VD�
e��-�!���h�LK�r.ǻ��$v�WP��NA�<N�Y���^�����B�H���f
�)pE:°s�j�Z��e�{"7a����-���]�yv��6y-�8�	ռo/b7�%��X�n(��6=�m�ѣ~��fh��j�Ң)��5��h�sH�2��AJC��Ԓ���,�T���^t�cwtL��A��٘�I#U�]gލ�j�ky�^��v��_Xu�x%F[E��vl���L
t�^q}��a�J��rV��2\G*-�6���� �B�:f	@��^ѷ��Y�<z�.=�!N�v���#����A�&�7%�"�,k[}
�r�ު\��rdE�э�ꐬO>��8hz����k&��g$�l���u��5��%wy�;ʒJ�9$�A�jklM{��b�K�p�a%�Åuh��U6�-���4��.^^�/�Md:�]b[:�\��u���>}y��M�Pí2T4�C "����u�B��S��h΍@f!�~�'d���@e_K�8:Ѫm*�Թc��<��]�7�3��t�����Â�C��Z����jS���yz��)��ʡ��,ҽ	PE��K+��9O�9j�g�j�I��:�A3�U�f�(h����]�)-�;��(#��jV�'t�'Mq}eg*��1��1����ݴ�t�眛��r��2�����5���	���ev�d�!��e$��T�mm;a�$v��w͙���G5�����L�I��C ���� z��۝�U:r���
�&�P%Y�����W΋w��AU�OT�bU�-��;6õ�g��x����r��d��F7���<{�����Ү�Rn"��W�\��yA嚃*T�&�M��݋v ��m<h����Z�P̹6����M��`���s�����(c�X&Z�/�EJm3^NL$�;���K/��G��n.oޖ�Oi�	�4�'�Mu�`p��͝��l����>μ�"XEٻ�u��GhO��k�w2~^iR���l
H�l[�>����])s��`t���qi�*�&�4�WE�J�޺��n�42�~�q��8�i�k��ľ�9(I��|8N�] �RQ=z��{y��i�z��\�O�%���;���m5]�y33Z�{w-��J� e5Z�w%�.9|sj]��G�S�,�k2���[��%��nۻ�}���Uꡆ.���9��C܆-1i�C`0;��
�$�E^�	Ǣ��[]m.ۡƌ5F�6�n�4a�.��
�-�ʝ�������h:fx���=# K��
���V�]M���b:��Q\<���{�FP�KU��۶���M���&P��c0h�Rb�l��v��&#�#���O��*_f�l��A�7�-�
���_:Wv�T[��G�����R�C)F�bn���LAص����
<���鞭���Mlӗi�\��[��76��[P�v!�:r�_=��[�j��O5n\�w�RB��D���p^��`��V��u�W1jAj[B�uiܸ��\a�kVK4k��\j8㙂�\\���JەbIB��*�Cզ�S1R�:�^R���gs��-lqvc�S*�m�̊ O��U�����*T(a�E|,�=�Ů����J4\��n�Ogp�'n`�77�p$ξ��B2�h�+r���^��Mz\Ñ���YṆu:��F���lՋ�#UOa��Y���ǭ���k�eΔ��V���г���$[z���Yy�RT�	Ǆ{����n��wB����-����i|]jz4j�kI�c��A�.��uҶPOn�m�r�t+�Ƕe��1`�O�j<���S�B��Oq�i��,1]��f���[ǻ텞9t�����=�;�5�R37t�rc�̺ۤڰ��rGu�N���Z��z�ӫ\fsZu��H%+w���:lY��6����L�XK���HuR��}s��j�tZ����v\Ǚ�ᯭ���������f���b9j��v��G�Q��Z�WW�wWhrPIca�5ӕ�9����l�)P5��M�NYge^i�R��G���lyV�#���'a:��z���T=۷]�%D��H�>�'C:ɲ75C -���,�m�ȻP�v7�Q��w��Y�u##�����k2�}�8wn�ưS^��t�e:U���ާ[6�x�R
�լU�f��:��Ae
)������N��]�6��Xˬ�v�_�bǭȣD,Y,'�m�.guna���ը�kx�v�zn#V�ܵ$��L��erF�Ä́E�ȁ����׋�b�U�9ko9�x֮��͡�q���4)f0f����I���o�	F�p��muWs{���w�h$��+������r�ȫ2 � �����{��s��: �s�jZPj�J���q�]���`���f�Qi�tm-�j�V�Jun��Wf�vwf�]���(��
�lvR�|����[X��to��������>�4���q�B��t��̐�����cT�w�ڜ�^����YK�1}����Gfh�J g�u��(�{๥���K'[T/P���$�[�m��0����s��!t��zl �.<�%λ�g6�CL�[Y��xչ�{n
g�K\����3)���e���P�н���ū<쫺Y����:e���]���:�=}�z؅��!���T��r!Ӯ�V'ʍ�:�I����\�aؔ��p��� Ѥ���:`�z�,���4)���>��kim�����v�eҕ%eLn��H��AL�7{fP����^[�qj}��mU� 8��]�fw9F�khci�#��m��L�DQ�!g8%8lv#����;�����&9��]�&�.v�	�a78Qb<�M%����{�d����b�<x����mf���U���*��K�T\f����8������"�m���]�����*5�W�ɗF��۹����� ��6�ǫ+�6���r�4n�m������M�r�?1!�9h���W�˱�˨)^�e��l�/�WPu���6��L9�ᬒ��Ä۫&�r��`.C�����d�����s3]>�1wYmM����n����.��RV-�.2�5ߏ���~��Ů�.#�ap��9���7W�t�E�մ��v�,X����/����if�Q�.�͠�L��l�H��:�t��3R	Rêf���^�8WF�*��`͝/v9:���G����ǣI�ͦ�lW���j�D�g0���gF(��&������-���m��.�
����a����ҷ&ouh%%�w/��s�z�:���Dr�,D����b���uiLgm��	d+�lv5�=�S�+��+;J�4)�f2,]l������}۽��ʆS��E�R�Z�
��f����o����(��ݢ��Ԛ޳)�zx���h����-�v�5����E=s+[�������&����Y����E-L�CF��To�p��r�dl��	�Zf�k��z�1���oR*.A��Ý\[p�c��3�v䭾dm�����+�i���A�1*	ۣ��rZLM�#!x
�|i]��upX����kX�,WE��ᗋN�{f�k���F]��I���K ���2��7���"u�j,y�5v�V���}m��e�ѩ��"������;��T�Rv��§�]vJ�q�=�8cI+Q�vQ�R�7�K[�q��h�&��#��w�C���W,Θ�*�&rkP���U��\�ŃU��}y�dP�]=��.���Wvm�=Ƃ�A�k�u���
�� �Z�����V�C�CT����E��IZ��<�!�w]vN����=e��-�; ��$Ss�W��Y�ż*#W��ɜ\mK�;6�Ӱ��9`#������A;5���N.ve����h��-{-�W�_(����\�`6�õfP��K�Tz�)yCq6���#>����s;�[�Ŋ����MM:��t���8ڋ�oluQ8 ��ݗ'gi��o;�zl����\��9|��@+_R?�nZ�L�-w�t��K���)�l��b�<v�q�{f�}Ԛu{9ju.Y���U�����>z����A���Qn�`
�Gӆ��	4���"��a��;	o�қA�@��Y���|����r��wAy �N�t���a�O��)X�\�m�i_VSF�c�n�JW�'q����S%[����嚮�;��ynKae�N�n�\�D�:b�t[���������Sq��ӫ��f�L���f[J�-�u��Y���1tt��&�Y��(F�.���iЇ�9�q�q^P&9�f�ën�ig7�Z���Y��0-C��F��M���Վۉ#]Ƣ�D72ݫ��5��iAP-��gZ��la(�8֝3y��w<�����c�I	6A��j᭺Ѽr^���LāsnU�cC���K~�L�]��%� �)B��ȩY �<Wu�X�8�h�w�SY�\��+2��K]D��v�g���0�̍W ��J�v:=ni�/�m�TIm衅��T�V�h4u�.�M�S�nu�B�n�ߊ'(��`��b�Rz���Cq����䤗E�s�@�\u�OIYC�n��c�������+��+��f.����6�O��b�B·(�W®��w�x���X�o)S��r���nc��d��ovJ��ۺ�;����Nunr8N<�k��mXYp�Y���I�[�֓�\���{J	G+E. p�c]�n�6��6�o������lw*B�
��.�h^�q�Aj�����v���rm�j�-�-pIr̾|5<�۹�d>����ok��\���,�.�+��P�a(ms�*���]&��r����U���#ك6�LR%�U�on�K�h��YL�Y±b��q㇥��4��b�k2�-�^q�q�w�@s�)�FP&}H�B�]2�0\Jۡٳ{���e�ow3��]ڌ&����Qκ�`�����n<��ا��<"��.W�Q��;*n�,ǃ�2z�>9�!�m�n�E�:չC����4`הHO�R-"���r(f��:��$U$��L[��J�e�g��l`�n�*��6�1qU���d�'Jj����/�;��c6>�Q�����|wל���V��\��kjsﺟ�ɝ[c;�����
fIǘ��-�ݲo	��S�ñh<�n�{AumMZ��>]��u��muX�HQ��'O���s�:_M�.����\�M���/��%u�8 �4������+��х������Ƚ�l�*����#�
������|���5��~�@����� ����N}FUޤ1h��t���H~y����ز$2�ǲ���r��%�WՓzsbf�%;��kR��C)�o1Nw[��p̧�V^f���7���"�������Sb��y���˸r���h)�u�L��٫�����;�O��r��J�V"8̎���)�m�j��v��Yƭ�Uz{B�2�˄H �s.E6L�Z{P��� v�6��{3!�:�Ws�4���՝���ܶ�4��Y��N�YEe_�2�@�"q�!Wݑ:�o}f��"�Y)t�x��X����c��ü��YѵgS���*��\m�\�g;HJ*T5�riMR��r�1�p^�Py� ��jDQ#0�v��������Hv�u��"�\���n�Bֻ�F`+/u�ۖMm��|MUo>���q��K�]�8� u�|4h5u��n��8����re�F�YSF[�q���3C��a�s�1MX�̣�2h��:�_Nۼ7o3�9xã��S�/�}b�#��X�M����ښo5f>�ZkT����m��ࣱ[��W�3�����#����mt��Tɥ����5��lT�>�7n�� ���٠r��=�`9��y�P�N�^�L*U)DάC�&V��b�K��kr"�ȹ�c+�����&���W�(�i^�� ���S0e���hѤ��V�r+9�]�y�I�Ł�YRe�i��un��&��k��[�Y�%�*�Ŵbq�����Ϣ9X��D�H�.�����kۥd(���ǁ�A��{��6vʣ�	�]��!"�VV�꣪0T�!�r��s�t���)����D���
��m�&��:����EX�8�P�76�w��6� �|d���#�5�Ca�|��3sy۾�J�0R�!��R��-����Vi	�'���AN�+WP�����t֌�\3/��!�sct��mKm�9�eo�R�D��^-؏&�3���Ʋ������9����]�H��, ����s(#�����j9�1;��M�]���:�\ �&H�P�0�{u;�tf�8r�c�
�����UX4��#|nWw4�%S���۳��6��d�����{m`�C�T�u`.�K��hlVb��I'tG�	z5r-ꕗ��ʳk�s4��Yvm*�<�:�2Dt�+���U&!�0h��S�p�[;�^�YMQ�!][\��9�ݷ�F&V>T��t�1z�7ۙN
ˊK��x�(M�&L�UA�$�ޗ����R8�l�uX��b`�:7������W9�6�$m�c=`J�w������,5:���l򑺶4��7,�T�B5�gJ���C�q&WN��մ*���ӆ�D�j�(+�G�6�_
J�V.�3պ$�|��Y�,��;y�͘	�ƻ���y��}i��A>Fo"}*Ƞ1H�@L�f�MYۚ*	���-ؾ��"vA-�d^�(A]��.���4,]��S:4w#k^��u5��e7�V��3\�<�W�mN���K$����^N�z�5[����݋��-�����P�ϖ�a�u}��A��-�o �K�{ ��1UջxC�Q�*��궍�y�*+ښ�9j�I!�W8)G`��b�@�&�I-օi�#��˩���-�r�q�O���5�9�+��i�8l}8ܡ���d��x�5��V��k�(I�^^⇷��Z��C����7�n��� <]o��D�o;Bն�5����i]K]�ګ{X��4K��)�│<�կ�mb�m��"=�K������ۍ|��zs4n�����Bb��Wٵ� Y[�Qű@�G�"�v�Ǔ�t��Q|��J��\+Z���b�=��gD�$�dGfq���]�Kh�MvJ�EԼg�yt;�cU��U��jUX�a����7�P���m���8�R��z��JI��NgzMY�v��lc��A[;�з��@�u6�N ��Z{C��@ٶ�ugGw]G0[�oL�Á����R����bGW<�ͱ�2��*�]E}p:�y@c�7HQ�mä-[�6�~Ǉ&n��[�<�p�5ג�V�B�zly�L����H_irp�o�=;ך9l�k��3FM��� mJ�IT�\m��B��[�}ј��[�4ⱜdfW!btw�
QhpPtM���V�
�k�i�{"X�D�gS �C�.������\���w�r�l��2�GZT!��5�@;�娡åMxw�(����٦������l}yS�e��o+^Kh�1�,ǒŸJ=K$mE��˗j]��{&mZe�z��|�����6�2���9G�gN�0�ߠH�����z�^�L*Ȯ��i�Yi]���؆K�����K|��Q�T�[�)Ǯ��-�6�"X$��]X�wG��[9���`�5���n���w9sv�Y��`BI\pD�-U�|*���z]���qX��7�\��35���f�ǄO����@�e���G�s\ب��'ByWF���!b^R̉���e��A3�_^F��M�*�Ob��5�N�֐��t[Q��NU�wkuƻ�iΧ{cH�㾸(�1`��9b�eW^o0�+�-�5,+Nu��n��h(��6L�+R��#=�����Q��vṹ�N匳�@���b��pr�9K��%�Ǝ貕o>��r��']k��b�����=���%��EiBWQ�P��N��n� ��'j��GVj-�׏�TL���(Rɶ��������XՋ����qo��A�������Hd�R�c�|�162�{��R�e�_J*���H�͡�IoYC��Mt�hor%�f�&0t�0ۭ*�q��xXvx\K���KW`���)���ُ[�4Ӏ���rP��q֮�9���"5��#����* �#��l�LA4#�i�\�'f�&rJWf�1mm_-1\�u!�3w�0�HEus��f�yBe^���ĦT��%f[��o�w��hm.���&������{�S��*hv�uV��&�|��0A�e��9wy�3��h�za�iF�r5u]�gs;���{QV�ۡ�Y"��Չ!9�6ė���3��o��ݵZ�g+ѕ�]�>:u�t�t�RR7.����p:�Yy���`ڐ�8�҈�� �5��P���X�3ot��]���	)�zP���z�L�9Ǉj�ݽm�[.�A0h;��0Y�h]ioMe�h�S�r��V������X�z+�EִϬ�{�þ5�f��E>�}��b��L�zyV����Y�A�Wwל��^�_;�RG�{���ZuC�誼f��ۚyrt�V��� �:�"Ad\�l��x��]]=�]����&�yF�N�'�Alѝ4Uުl�{]{үhb���K���Iy7)�:�n�j��� �ړ6�^9����4&�*'�7��2�r�S���9d;E-y�e�v��}��h;1���.:�ꑖJ�i�qM�pR�p��x!T�	�l�f|��A����q쾙;�2�J��)�Q!�{9����]�z�&�ZZ�i���9�$��%��QwM���'b��.�c̈́�a^ִ�E�o��6�eͮ��F%b/e��A'v8n��4Ï5f61 ����/h��Q��X�:�_.�c���\t�K��}˾X�hu�wVLh.Z:#e�1�]�0VF��,fE�vd������֧�1e��;8�]L%�������D��������+�$;q���>z���t)�K�اnoovC7��o�zF��n��or���*hq��B8�h��!�/�"���!|�RT�R��N��b�WsluEG��ͼ�"l�G�Z�تṊ
/�[�*�u4���G/����XՍ�Ž;������x�B���5d��V#ʵ����BC�Mm��b���njW��7�]K�4Z"���=���\c�N�)���GA�$-�Y���_4�!k�E:���0*���{ml�͇y��ʶ�k��Ow9Kh7�FN�{�-y���y�%'�#'v):�1�#E�ǹYt6s����+� ��h�M.Rv!Ӽ�ovZښ�f����>���Z��'v�5ڎ[{�k0�a6Q���kev �v��mY5�2�Nwql���m��^�`֞�x�yJE�����\�/\/���ˬ8��g2�p�r��Ƿr@(m U ���gႌC""�h�{���U��t>��#�1JvMf�3�~յ�����Le�.�e)��¶��L��L�a��M&t�jA��L�y�H-�]���Nnpsޠ�_F�(�>���n���`/#̂�M�_+��k6�NgZ�=�{J�wv� As��x �b�6�;`���&7�;;x��,3-�Wq����V-N���ܳw6��OS�6��W)��2��4(S�]ZwuQͻ�q��f������OU�Ӷ��Q��G�k�P�hv�bPK�c��(�ۛ.��M]	1s{�,3�>i��(�&͵��vL�����9>��F�곰ƠT/:��U�x���]s��Հ�+=�o�}��r�pP���ۥ�P�|���*ﻇ_a�c;��eH1��I�R3OF��!a@Bt�
�Tn�m(���)|��Hq�
[D�"�h<�e<�4&-.RWX�3[��P\A�f�JL=�H�>S9/��dLN��%��!��/8��yj��K)�CU)Zpɜ.k"yR)ȇ��(.��:����2�gv��ua��meH�KQ���蔇@�m9j�w�ʺH|ѰVi�u7ʦR���p/��e��q�Cϔ�Lr�n��c���|D;�2�۳gFJ�܊��q�-�
���ɑ�F��+4}���hȒ�p,�bm ��`�]#^��6��c{�Y֙�zh^���7�δ)%�,hw��;q�����
�a�C �u(�� mb�{��
\�N����t��C����SAf���T*�f�Q�fz�n)�
h502��<��]�TZ�v��4��70ZVQ�G�iiXUcH͛��쇬�u���<D�`�Uz�� f�Ӗ����C�jD������-@�b*�������r���,��� W�s6��5�N#~��Rr����ف�H���p^t�]�b��N�x틧����Qt�O'9�D�F�[���.$�ƌ�� �X��)\��Kz��16����ݝ�z��>l=�1�uG�,��ewCo�]X�Z�R�o!��:4�g��
sN9h��ͮq[����n��L��G�bb˂����V(:�_W;���9]VQN�˛�S�I��P�r��2�!���q}ۘ7�a�$�� ��ժ��{.��c�_���t�h�;3u�$�G1���QV�P�1P�L�0�V'I.��,Iذa��@t�:����[(�s��mf�$���ᷯ�f#�%�6����Z�zyQ�}L�B��:n5SC9�`��ň]���v�Haj�i�z
<�:+�Tŝwk"��b�v����إaf�Ƕz)�U֑�]q�]��F�X�қ���*�)\v(2A��'f4��Ny���S�(7���F�uڴ��
�L���r�<٫�����D�X��WR�Bf���l�Et�����>+�`t��n�u�M��qbU��X�ʵ�ttŤ0P����9]�K��̫EL#ݻ��1S�ojvZ���s�Z.)��a#Q��z�qW�b�+�%t�"w�#䐜�\r��p��oMd$ʔ�"gnIn���9d����u��o\OrD�'	"��r'��r�K ܼC��T����tq�ڙ��|�z��,Ŷi���5پ��b�ړ������y�]�C�[����u��u�Fܙ�*��ԟ2�*u̫ܦn��ѕ;CM	Wκ�w�Z�X2bKѕݴ!�	o"a�A�yխ�]�}FQ�K:W�y]d�x�B��{��0�Q�d�D���!G	<�ł�R!��l��B�>m���R٭-�-R�u�l�h�]A�"7�FC���f��[��.����h2�pe�:q�벸�{π�i[{���V�.I�;��nE��nAєn��֜o9�δ_'V�ԡ=v�Z��4�rw��3>wp��ﶚl^b�W���BQ���}�K
eu�(��go2뷻U0Tg���MI�-Ժ�r���o��f�j��LI��U�=yfۃ|�G�)�\��0��
Q�&&Q}y�	4P7{�g'�rs��x%}ۙ��m�3"tn�m-�y��9�S�[�}��c��`��&>R��j�c�N�6�Lm���<ŷ}�ؗf�86�^\�plA��8%�x����(<�8���lgs(�|����Պ �� ���b� �&�uk+�ӏnK-�PUt7�j�.����x�����sfA��E�٬X�Dp��Ґ(d��&�A�� �u��w��>sy��=K{P����c>�H#1���,$�/��8�(q��aP�r�J�R��Bxn ˦����g��ej3"hV��e�fh��l����覷���K��ZYb�iەi8n��Z,U�aHNܗ��h��8P�i��p���HCX��ϚT/M.LK�W�r[ e;+x��A�[4���w���빲+�U�;��ed�3@��C:�,�j�mڋ5�yO�����vҸw9B�iK]6�̔Nkۅ*�뚒�1C�خp�|[���mk:��櫶���T�N氐���_-�+�R{9�N��Qq�t�>���"�)RLwd�^*W��{w�؆�sH�O�lR���a�7�T2e��~��B9&�],"Ӈw�k�Y�j-�ᱮ��]�u��+kilޜ�ݎZCn��c��a�Q�{�%��r\0�󊥌�C�<����e�����cK�}9&��=�z#��z�T/:u�tL��+��/T�r�}���x�G$z6M<e-�$�36��"�tDq�T��^�m�wZ�q�)�����Ԡ�ב�{A8�
 ^��Α5�9���A�iCP�u�B��2�-���ٚ:A�@`�\�����J�d����+���j�9̌K"�5v*��
	��ҫ���3I�htIN^��z���&�39��.�bcFT,��p�N���}��Y�u������dgusT6�u�{�o����,H&)�\�����iU�2���aٗ�&Q��X�-0J��n�;��S32���m���*�j�e��A�'r�*����]R��_\�	�Q�Mt9Z�P�X�;�I?�x��Y|�j�[�O�f�gqW��x��ٳ'��p��N�S�L��t@i�3v�-�Tp�v��Yk0v�0���RH�6�]�����-�UD��IK�T�Rf*�9��p�3u#���n0ۦ���Ļ�ewV�S�ϟƅ��*٦�105ս1�����͕�뷶�m���mD�q�n�Ql=ٺ�̖�J�;5F�s��{p��Ю�wA ��y��i�$e�<fl슳n:���j\1cL��9pŖcV�Cu�Hs�-^U��7��6xt��L�:T�9��|��N��'j�Z��ZL��*���}�m�=��(0)*30�$o7V��X���o&���C\�,ḝ�Ś��/�7���y�M���ږ*����b�4T kX�m�VR�F���V�$QV(��R�[b(5QdQeE�ZV-�LKh"[`�AA*6���DJ��6��m��b9,�U-��U�
1Eb�Պ�ch�*TW-LD�KkkmIZ[����ƴ[eXVT���0CUar�D��X.eS�.f5���`T+DBұB��KZ��AcZQ���fX��am��Rf2�A���Z�ˌ�e��帕
�m�*������b�VT�2Ҳ)Q���c*婌�#mj4�4��eE**�m�*D��\eI��LE� ��չB���PYY�(�+)m�m
�2���̵K�c���!F,QDeQ�T��(QZ�hQX���(`��(�b��6���-����ܝ���S��{���. -wX��k�Q���Taٹ}NI�\�u�>J�k�XNR�g�}�A��'9���M�pPR�ޟ�$����V��f�fAn�U�Y]k���
�F:����Ե���l	wg���,�"(
��/>�����a�>fWr��-�v�QY�ۖ (E�ϞQ�q��P�3���7�������Y^��8l��dW�ָaH�g#k����i%ZvggA�%�~�%i�����q[U�r�i��P��8�B�w�x�*@���nIǴ!^����U�/vu�u���5�-R���yK�f7CM�Fc���*.e�M�N��X�|����Z�pHs�<L����4����+5���Xv���G�����������U������}&�+#�S��P��}_g;���-*��z�HS����F^d��z{�.�=�v��Dt���𳊥iw�?]!mOї,��Vo:z�SE4�˻��^�U@���g!���gM�Z��F�K��M�:ir�dk�Y��yn�5�{eK�ɓO��-�A�滓�0�)�/��.	�R# ���k�|������*�m����	<����-fVw�-��y��a���k69�t[q���g�o�]�&g�>��+A�b��
��܆��f8"�5�z\w#6���C��*�����i�J�-��fh`��iY}��LG\�)73�^ݬ���`u�o�m��x˥ė|4B��J�\�9O[�����f�,r�T-DڏV�1v�-D��|�&ѵ��7�ԝ9�CP�N��=�>ۺ��a��k}_cm^� ����a�m�|����#�>,mk������d�W�ΤH���d�`�g:�X�8��#�r2��C_X���K��C�x5�f$D�Kρ�V,Fe���Q4�LХ���`6�MR���j)�渿�wL S��29j1.(P���і����Q�T�5Hd�Aa';��k�k�Xs�́���M�p�E�;!�������P;U��"���k�	�������ۭj��g<@�oC������]�))���V!��Y�]8����r����'C��N����aH,�B�qu�4�4\�-��B_nW������`���n�����U���y��g��
������:ɟ�a�htE�B�q�`�_T���+�%����Χ����8qW��#�p,ȵ�dWٕę��J���W��w�ӵt�]]x�v���9�F���$�Ayu	XvJ�uf��9�9K�B!kG;��q�k	�F�i�
�R_-"��aV� R��7E����P�'&�p˻���\�__oF8G6��x�*�f�J,�K�A���S�K5r'���NT8�����zֺHȩw�n��2)H���=o���E>�8�뼀��b6i��x�<&}o%CK=���=lL&�����'�U��ꋚ���|�,9����&�N���#t�:,�0��k�,p�8�V"v�D�3�J� ������ΙT�mn��b���}@=�Z��7V袲��J�5<5[(2��'����݋籥�̉=����6!��3ڤݑm���P�y�����a~��qx�mD0&h��a�Ԭ�{k��;�ɝK�\�Q���`�j�}y��V);����v?].Wz�i�5YΗ�.��Z�e���22��w�p4���9�r���%��|�{ó��#��U��qyÓw!��C1#\]Aв��i�"A�a���C����ڎ
�w�dp{�Y�{�ꧧD;�R�؍�	��#�کͣ�dr{�M�w�x�T4W�m���"�S�Ԕt�H�t�V�Ǥ�y<=b�w�q{6�O*��]hPh3{�x�s��ZTu�&��n�)�R��aѴ_L��Ѷ��#6)Ef�E�� ,.|ҁқc5��H��f8_P~�x� [+�Of?%[ ��j�u�c�M|��ܱU��3n�qϺU�Y�fGaWHFL
����J�V�)%Y�]��!ڋ+t�囼~�T�k쬳�֔���W�H�#{][XrV��K�΁?oF�Ry��vy��[��yuH=S�즕�ȣ��o0��,E�Y�^N�g��0Ξ�8�}$����
��y��z^ޚu7��!x�$��\r�ࢎ�yp;@����B�9�LiynS�N�=�� �:�vL��/~�"kO9V�{�8�}�Z��k�K����Lϴ��=ǋ�1��^�d��U�(�;�g-I�V�+#��U���dt[V�\�LV�QuO;^��^�=�˺y�T>⎘��΃�6rY;}!�K�ťs�ſ՝b�Y�BF�n����C59�m����[�=s�;թ�ؖ�pt-�o�9��A=�/�VoyZv�O3�+�sgFW��z����e�#Ղ��4�<]g��_]<��X�1W*�z�V�a��,��q� ����s5�}��r���������Vy�C[��ʦ(Y�k��	Ջk�"�W����H��z�gM5~x�0r��o�z��� ��XyFx��^��=9SNY�d#t�OP�m#xf�k록���}e��8U��Y�wE�h����'һ;1ⵙ���i�ۡ2\�}J�-5�( �o����O��N�!\;�:�3�:p����
�	���fQxPtNw<�5�Z����w rZ��0N�:m���#t7�nQ��d�4F��ݢKE�aZ[Sh2���]���]��,�ۘ���8�D����L������D����#�Yb����zy��]�^�ӭ"�.8��]K���Aw-5��u�ux�qW/k�m��c�("
��f��Y�}?-L�-49���z�8�]J��r5��o��@ld�ަ}�#<�@��S����R]�]�g����A��A��eg�	����K|��բ�s{��ʈ�֊�=����.x*O��g2��#��7��4=�k����9�����u2',��̒u���##��Ƞ+�e�_p�-���爼=����b�N-+�o����6̻���p��~��'�l$�����e��X��忺+j6�no3�Jsڼ:3��6aD<�gk�����;؋\yT�]ʵ_j�7A[�Y���c�M�>(�s�"wF	li�-�T`!��o9�7CH�����f�=�Cjz�0U<�rOqԧx>fw��	:��� R�Lѳ���$9˞&B�\��x�Z�P{��������J�&��,�30�ՠ�mu)SE��G8��k�����U"ޚE����8\�D[�{���O��؅w���oD	��h�w��#�w)VW��}����&��Ձ¯���Pl��X\mq�ׇ>%;��|hj�9S��0\�����K�:��:Ũ�﷋��p��a{	�i��U�3�S�+ѐ]��eH��ڔy�Cw'�C��+N���~�W��^pﯭ�M��\��,����_�Qxo���))�鲱v_U��w��!ѡ׎dE03`qܰ!���k�8h=�Z���&��Y�جt:���A�Q<�v�]�:o
���	�5o'V P:1\6���,֫����1�b$4��7<��~��8ىK�x��6l`�}9�= |��>Tt9f*��=T:m�(q�yH��5��w��v��$bQR���4������[��{����N��`���Z1DtFf����d��ݩ+33�W��5	aީ��%k��a!��vP[?u��c���7���:[��Y��Y7�����s�C��C$r�PivK�yܷs�1��t����z��|���
��y'R}����ｨ�r�m.)�<<���b��C0��/�&Z�H�	�keU51]Ꮨod3A8�N��v��H�AY�ڮ�T�N�qz6�z�/�A⫺"�B-��M�:� ����0Qȭ*�3ǥ����8���-1��N��_;�`��s��wu$;����g=��,���3ݬ)�4'#��#\��%*n6�;��QIc����l,�z.��}��Aoe�o��ǣ��D��U�Wq��1r�Qf�J�O5�w�W�/�0>���C��I�s�.*|�|�P��캛J�&�Z�CN�.���A�����ơ\�H��3�����0/c�މI���^� �g��ޮh���ʌ��d[���T.q"i�k��Wf�-W����O� j���$z��8�x!����P�&[�w�,G0X̳?Kp�U}�eF:�2�����V���>̜ ����tU�^�]�jN��S�e><��^�����;)Z�.8��H�Of;�@[X�,��ޒؓyֿKY�7}�8�Hu�{>w=:���Â���j�u���P�B{g�d���Y�e_����Y
}u�*��Y)ў�ف*/�dGШ+t��(a���L"e���r���X,:�^�]<�G_��1����$�h�K(hh��emB3���/b5��]��؇D����G��j�Zz���z9�hlG/
v��p�%����8�T�b�S��g�a�y4�f�1��LhcP9q��x���Y
X���~Y��]෱�
3���t�\>;!�����l60_� ��|,-���_<���]�J��X�{�e���q�"��7:�Q�������л���s�m���stko��7]B(�x�6��۷S�:z�����\
� ���['\�E�~���{�гU
|z���:k��;����>��x��<�I��U���gS�y��E�����x�]�׬+t؄��n��� wb�*<: q��;K5�
���<4��ǐ�1��c5;mЊy��8F��F�K���m�<M�Z1ҥ[���8�{�Y�GE[�ޛ�v����[hV����9�3��Rw=��̅�s�x��뵆Z�5�����K�({�(��x��}�������d�����i�	���BK��U�� �vؾ;��>��/��%�r|��l��~s��\C��e�;�a��`3uU��q������v�i9ϣ*��8A/�Z� ��
(�T/2GP��P�0�r9�x���ZG���h]א�0_.���׏+�d-��c�/y4�;I�3^R}Eo���n[�'-���`X���S�}n����rT��^����.�M!f�r�Žj<�y�+�c����L�R�X���a�ۋ���t�
s�i�o���|kMPh+~�� �ͮ��d/E�c�Z��6���^��^K�Z��֚׈C�W�v��c�M+:�H�[��^a�+}�!+6�̬��4�

�������_3K��_A�������rÚv��+i���-�q1ݹ7gZ�24ؒ�'�9t߫)��'gD�J�?���gz��Ҽ(_.��gd�/K6oo��b)Һ7��On��]�PwfU�!DbA�6��!FL��d1��VU�T��Cᔐ4 w���EFo���_<;�S�{.*u��9rc'����6�k&X�Lem{q�E_o�2�SY��ɩN�erc���z���@-tV�R��>u�N��:.�b�[�<�K2��5t�`柍u�rڰ1|�b��8�)�3b6W.�H�@f�~�)4�q!
��}՞�@����H/��rt��o9�A�c�Z��0�����8\H=˻�˝��us
"�FKn{}��ȟ t�'�9,��_D�s��瓫������8������Y��k�o���f��7"��%av�.�.��C�����"Kťiwf�Yf�9�ؾ�`Y�����")t#OV$Ob�f��J�A��
�VV���kɎ���Վu%ޭ\b�-�$[3D����3\�Hge�_p�-����#����Vr�� �]���dx�#wY��SQ��ċ*E�n�-
L�(�{�2���]GB�9r͑Yƻ��p7Xy݌U��������'�2QaZ��$W]r���pKh�N�'Xk79�.�]ko��2��Wu�a�Mt�]󁳭��yf;ֶ�c}�b�3:�4'�h��;Z��Mʹ9k�s:�N��빓��V���}��m[�%��}G��`k��t�j����[�M��>X}��S�	<�͑��"YlTU����4�3),��[6ei����QSI�.��e��VSQ���zf��Y�kf�̑?^�*&�q07i�f��P�tF-�L7��	��ә=��#C�X�c��#�i�-�+u��;���|��f.����A����䃵g&S9C���s�8n�?��]�v%u��H�{���,W\S�*w{8eH��i��;�I�ʕ�co˿Vs�O�94`�f?�}":n%��̹~.'�"��#�82}j�7��_��w�s��j��_l�+#OS�Gb���{l=u��A�� �zW!���(������ʞĶ���ʣ\ӫ`6
�U�k�:��#k�Ʃ2	��|�.Ī3~����}�N�Gi,tn�*�+�x%󿝃�ڳ`���\]��s�)#;#Nh�8�ړq�9��pOm	�*Ru*:�^��D��s�}��}C�ŗ�M�����O+N�����a[5� 8R9۳'�c��\�nܬX�q�J���;M�%�� ��r�D��tⶅ]����#�+��kz���|:}���f�Ã�鰪_o-r���1@Y,`x�������;���h���NAt�0f�ZVq�L���36��Jb�Kt�5]psw9'Aј���P��oT�c���5�2���Ws�(�[eb8��q���4
�[����Dwu��0�\��0 �{{9�P��9�T�]��kY��XI�wnT	o�+8<$,2Lڋ����*�U�m���)�셕����g�K�.f�J����6�c.���z#�r���?,}]�e^��� �FWr؛Y�$�H�YyVwd���3n�h�z9d8��(>xb�,��뾼3l��j���KA��׈�C�w;4>% {�U��jyZ���/�AR�i"��}ϫ� 5զp�v������0�w
�m�y�ͱ��F�x`{��f�"on�{$��,�`��ug�z}��N���40L����2��sW���c�/�Wܥ�Ww�������s��ٮ+7��GN�vu��u����J��}/M>&�GX6�����^�SH����#ow>0D�V�
d��6j�.ޣj�ŋam^`�(va嘻q���(�y��I����]܉�4q̮���R��K��';k3gn=�	���vn�9GP1���<Wkn&+�i����e�"=sJb�Y}��Ti�kZ��]�2r���G���*v��Y�kȄS�@h=r���d�y�e�z���/�Z�Y�Z2��9yf�ΜNl`*�
�s����������7i��Z23����\a���� �C��6�{��]Mi�|-qOZǵ��ה�-��e�R�Q�u�q��R���]bՊ4�6��v��N�5[�qЛ�n�n隋�Ӓ뺰v��� �P�XV/���y�h6y�ʕ����ǖdн��>�X�E�����b�A�fn93ۻg6�]ӨT�q.�9�=|�hx�ں�N��}X����g}�FQ�+KuM���˥U��ز�CE��۴�s5��lW�rs:�T�˼�>�̞FE5�u�eT�5t��@b����-j�E��ӨJK�*����\���u�e�g0��JH��
�f�f��z����nۢ��\:�)|&����06��K��s�A]J!o�u.�ա}&_���u+6�=ꎠ���e�&jF3�S:j��)s���^��z�MG"9�U�@Wv�5૫���ĳ�n�۽޶[w�80�n0p\�g&���b<��]b���]���7bV(���s���Χ
6ڂ�B����/QZ;�,X��{���Q ���`T�1�Y%Q�cBA�|樭��zطMVv�yJ�Tv�>}��sK��}��ݪ�$ob8�ܛۦ���-��y��^ۀZľt�B)�3օv�K>��QgOG��h*> ��b¥�c��TAAf2�̤n%�Z�Db0e�X��ű--j4�`�Z�X�-�Dj���Z*��(,E�B�kb�j�Yl�+QA�9eʨV��1X�\��kDQT#���b1Qb�-�Ld�ZPQT`�Q.d�)1++"�����PQb�apjV*�B�(1T�Aj��+[-�V�Qq�̱
�V�Q+Ke+DQ��ELL�m����EYJ�"!KTD��R�\lUDUr�Qb��Tm�Q���#hPcQAVڲ���f4��h��DE�,�VV��j1DYZ��D�ɌDB�.��5w�~י��^�+���=�pm��.�_
9OT���}8�)�7t�=b�p�]��6�qa�Ձ��ΗӢ�4��4�<��c�������$z����kz&�g�S�dD�x�I����
����a�bA|2�gP�8��b�����=�����߷�g�IS?o���m��Ӈ��{��<�gy:�٢��T�2�8�A$|u}Rz�g����[`x�2Vy���u��AgaR��b��?QV����A�����̼C�xì�1%B��q����7��
��+�[��V�U����7>���E,����`Q�x�/o�������w�ğ!YY*�s�I1
�w2ެ��Hc;5f�8��%G�ȲbN!{eM���Xc�3���c�'{�Oxw�y����=���|��iĞ�����>q��ܝ�<H*����i'P��u���!��o�'�񒲳��s����2zv�VT�����Ax�g��A���@�A?yn����NA�ݵ�����������Rz�,S���V��	�4�èc�>�I�8����9��LH,���Mv�O��Aw��I�l�zk�&�X����11���I��� A��!tx��y�D+��~���xʇ�*q;�x����߬�Y�J��<=��W�i�C�T>Ir�>�y$��'��h�n01���+�Ԃ�N�$�T4���?{h$�#�"e�ͬn��;�����sG9�w�G�}�}TE��
�a�z��MRc8�و~OC_�<H*�������1 �~CY߬���~���O�T�Hg�T�B��/߷�=@�:�O{̞0��,��Hc���`&�8�nG��>� D"��xz�B�*M!w�IY�`,�~��k(~I��=�!�q'����<H,�O�}�Xwt<H*�=��i'�T�}C0���Hz~���q+%eL<����*�_�����8�3D}�@���#�Vq%�&?�OR��L�`~I�%OsZ���2Vn���>qY<2���W�N�>�� i$���~���fϨk��}f�u��w�^��whyh�vQ�q��y~ �>Ӈ�>��;@Z��N�GP��a�����|͡����s��AT6§�����A|C�;�����+'�賓1%~O�3�k	�4��.Z�MY1&Я�!}���C�5ϧV���nnU�kh	�j��5�X(����s�.؋G�k���sʹ�Y���V[wu���~����`���=���$2r=�1-]}v�tSxD+HǟrT�4hwj��ky3�йN�䈖9��\�,���{��hD�uh�����%gW�W�~`b!��֨x� ����O��b���H)>�|����XW=;�<C�u16�i���kPm��~èx�Y6~�M!��1��j�aPY�i1	������2s^���~���������J�N�>`(a��M���$��N0�_g�'�m�@�i���6�y�d8�6ϙ��rC�?>�z&_���z�9��h�����h�'L�o���|�$�YĜB���/Y6�ͦ���<@�VJ�y����Ǭ1Og�C�/,=�����h��:�<K�VN5��Vw�*F���}倗Sԙ�Hd�t���xx���'s��n��x��_rMv�H,��9AM$��1%B�'���ST�q����Rc6Ρ����k�J�Xm�ל�� Y|c+M�}�g����}V��=���U�IX}��1��������*�_!���u
�Lߺ��sbO�CXq�&S�J�3�ՇP�ACV�N&0�
�h��O�.��nk�a�nQYs���*��}H,�=f'~���<H(y����z��c'��1� ��ę�����|�O=��'�4�eNv�I�'r�V�,�&�MX��%x��ii����﮲~Ѭ>����~��~�s8�d���O���|�}���@�0�}�u:�$i������s���Rm
��d�1;�w�C�J�ϵ�L��:I�\�ͮ�<w���YSQ�h�\�2㼡�Av�M���1& t<���d�Y�%k!��O\f�I�+�o�u=x���L���O;M$���&n����:j�Rm�{�OR�ͨ�ǻD�w�f��w����=nͮx�3���5@�m�Cl����Aa�<��r�ă�3�m���$�����:��M���i'�|��5��!Rq
�7�:�緬g������s��ov'�֐��*�_p��[��Y�J�X��RT*A{��8��0�
�=Ri!����_SĂ�!�{�����Ă���1ɤ1��1�
���CÛ���G�@W�9Q��#���Mcܢm�Y[����������q� <�kv���17�=x8=��޵>O�Tv�to�r��^�����v��r�ix4�gf�̾9Ab��v�[�W�vƍ�KNu�<p[�duÛ���+�H\�q5a��d�O������k��ޣٝ<a���R}��4°��Y.s���*��rM"��P�y�CYd�1XT*N!Y=O�.�X���}C�~O8����C7�1'ﴄG�@���h��P�E#[���]qy��<ΐ_X|�'y�>~a�R����4��Rc��kxT������}��Az�^}�T��T�E�mg�?j�I�*m��f� )8�l�B�"��DAb�9����潓nϵ��'�P�UDs1r�����f�!�����n����+����<H/R~�p��N!��L�p�3�G�0>CIP�=�i1P���C�_R����->�g�}�������s�m&��q?!������f�.��}N2e�|����i�d�P�����N�U��4���c�+�ݠi�q1�w�M��?QDnO�@�4�|���������~�v��IYP�>C�Y3������X(J���14�ɉ:�~���i^�Vx_�qaXW�X{���|��*߹���%E���N���v�����y�&�~B��>}���_��������u��"y���"�vE��Ȅ������Nr�0�Y<J�����A���F��b����<a�4�&=C���<H*�!��X<��H/ޟ~�Y>�d�y���~<���p߻������{8�2��;;�ĝB��=5��X
OP��;������P���	��kt�'���K�N:Ou|H*�D�P���$�{2�5��q��?{�Ԃ�3�f��xs{��}�=�ף�Ԯυ8��|	$xna�8��bOg����8��C����R��%}�h�'�8�C���O�����2�]]�y2��++�]'��g*T��8�'P"H���d��l���gt��#�"H����0*C�bw���6��u>N�Hq8� }s
�:ʇ����tCMaPY���|���IP��l����ed����!��w��ovи��OS>s�hx"�Gȉܧ��l�T�On�~B�ì1_C��$�.�^Y�c��P�?�}I��bA�o��N>$�hb}`Y>J�S��� �d{�C��1��sў�W��&��Y�G����1"NF�н�H�#t,�/��8\��F�vLҙn7���X5dVr���9خ"�]�������F'C<�Nwa���۔_d�ӚG-���N\4rQܮ�w@��rs�{�2��W-�G��Yڃ���KVe)&Y��=�n�E�g�Ԙ�1��U�'|���x� xe1�q�7C��e���Y:�z���Ou
�a�����`)<g�ܮ�:��S��q&��g)/����K�_������j���U�0v�{��}��Y{�'�3Ă�=-"�M������4�Y�u<=���1H.�3�
�C�1��dǈm�+>Oaw��%C�=�sǉ�LI�+���5����/=���S[|3�`��,2���D}ؾ��ea����_$c%O��Y�f�*��e�$�m1���Vi�
�����C�����9Cl���1����*N���?'��<H/T�h'��uZ��ط���g�G�@B?{=�N!�|��~��*�2x�I�*T
���>�LOPĕNP�i�J�*��B�ɴ�˥`)8��O=��<�B����|I�4�ɋ30��6��h�1�;��Nާ�o]h��h����Vy��P�A~a�7�S�i=a���4x�YY׉1�]�P�R
����2�Ě7�=M2g(~a�ˤ�E��Qt�Rq
�L��ߨkP�����~}B���o�������>&� m.����4�J�5M'��c8�{a������ �'���BLz�H=��q|C���3s�ޡ�z�Y�=�0<LC�1��
�XT�@��P;P�˭�����=����3�M m*Or�������{�ң�C&�z�7�r���,Z˚3t&�Y�g#)��o�r��Bm\lRx�ѳ�_A!��\L�����/�J�7:�_	6t�We��FR�l�]�l,�*��>����-W?��C)��Ɵ��#g��+�q�'ꀙ�a@zݨ_{�]o��i����Y�h<?h���q?��j��M���jqA��-���n�ڒ�� Mbuκ9".��(CZӧ7�U �j��JΏ-O4�k�ٔ�^���-����AJ�@����D��9����wT���$����զIs:u�P�f�.�>��Б���&,�p��jɹ��wro���x��j�1��wC���ӟ�����W��ӷ�Q<4�7�@��޾Vˇuun��W�X،CMv@�*5M:�b��(3�����^;�8C_,��<�zb:�oQ�ܺa���m1�D�}���K"�!��|�j��͂��n�]���_L!5A9�q8�U�]�Ǚ�v#���l���잩3�C�� ]Ƶ۱�h�s����b7n�|qy��XȘ4�I O?��,q�l�z�Ĉ��M3L솟Rl;���c��߹����ѣGy�qC����,{�2YE�6t�FG9qC�- w.u0��?Y�{�c<c�TSU�N?y���Y<ϰviU8���;��)�D}ʸ�.�ᢝ<<���ZU��l�+c��(�L���:�>%<�X���࢈P/�n]����|�hݪ�tD�p��X{]S3�d1��;�p���{;�6W��^C�	��V�I2�z]�8|��x�{�3��`�3���uI�ݖ��8�1�Å�׫�މI���;~o���K节GtW�4����w�B�"\��?���f�]�z�2����+�wƘTI��	Gjk��{-!����|3�&R36��}\q�QJ4on;�nk�)�U���k�[ؕ��V�����kvN�F�҉h��@��{\�{6��r}�F������ �̤{N_{*+�:�ōaQ�G�1y��9(��5,��v�ӌFNG�o25�yR?��γ�&�:~ǵ�^�������y�����ˏ&��wL�ؚ�.?YL�U��m8��V��PX�l�څhJ]g��bδ��G&#�f^�1�B|��j��ե�X74�\q��o���6S�pV^�l؟.V�l����28_=*�G���ʸ����2�u��_<����Hf)n������F;]G�﷊Q�z���\*CF�kG�%}�t�=wIP9�)W��E��pDF�L�3Q8�*��>����柮���Wa��o�_5�|L�5ç7]�+�xz�.*Ƣ��:�k�+;��ڃa����<lG�e}�zbB@c���|#�u*��vX�?i���K�C��w��a@�w=�*z{<k֩��9�	����f�US�Q�x�A5�}}�X�F\��:]�Q{.!���кI�����s��a�$g*xb�9郀sn��@�݊|���Xt�5�9}��D�Âywi���Ύx9v�+�1�lN�C��ګ������1],n�9]3S!˔�pUJ�PM�U���	`���m�\a}إ�LO-Z���խ�AA��]��F���36�H(]�y9��:�y����.�kN����@��ŝ�0MN��>d=��Μ�E>	�b-=��!�"�u��0��'�%��/�q��Q�ڜ�>Q���X�b
���;�����u��s�lC�� �:�4C�5��X���X�؆M�O ����@D`��%4�	�@��s/�[\t�E�sL�x5�!zϽ�ճ�t���|,�����)'�p��s���q���,��x`��Q�1�h��ǒ~���v�i�"�_��I{k���L�K�*���nx&��R{��$&Ĳ���6�[W����^��-: !����n����\�Ti.;I�E�����Q_K~Nɖ����=~��<6��v9��.Kp�O�+#���kO��j��M[*�=Aɢx�n{=�\���x(n���<nt�
s|�/T�����U̘6_E���G���i6k�e�8+�R�g��F�&�	��u'7�Y˷/wo.!��g�&1\]�ou�����g��9��%#Pc�J���5�%}�t�?�r5���n�>߹���I�i�����.]Jor����w�݅�9��I��X"	z{y�(��۫���*�޽���3.Ct#H:쐺�$�luh�֖_"��W�[h�`Oe!DX�=݀s���| �ޭE.���4�4Ν/6�1c�ȣ�d�y�f�#����St9�L��]?z���a������H��R����#�;ˣn�F�����nNt�*�B�����@�˵B�kCn\���M�q�:Qȕ�Q8�eq6�9�*)RՊ۷S*#�Q�A��d�0�J\h���_'-�?3v�<�!�S�;J9h$�*�\2����etU�c�RLcMԙ#H3P��+��]�f�K��-���"�K�T[�g���[ltv{fUτ`a�^��yP��a�����m[�,�y��xb����#:� ��M#�6����bk��.�%څ����_:�Z\ε��ξۋ��N�]M��Zⶃ�'��waI�db]�"@vS�R}��a��/����'=�:UJS���Wx��O�����p7f��\�d �ܨ��U�;���: ����"L��� �d_�������U͋Ze�¢={� �y(Pc-�{��"�;��TN��ð�+��8{j<STZ7 �-��1Ww�CY�1��yT��U��1BՒV�wPFOT�� �wW�*j�Ʃ��|#E�Ss�K���Yۓ�cf��+=\n.V]'�VX���+��C���y#�S7̜��1�|����eM�����t8s ܩٙǱ1]a��s+<�#H�Q���/�prV�u$�Z�<'� -V�ݛ��\���^�Mk��f�ME�"�2��&Fm��F�ϴ@�L���¬�H���ۼ���-x�6cqP�4܈�f���YT�_A!��������6g�`/!R�W{K��({��g�?��A�afH��u��5hu�Nr�<I�Fb��p��TT�sn�o\vJ��͆��|�5ΐ���gFᏓ�tܤ�Y�����h��� �ܘ�]�j#�EBq���V9�u���z�9n>�Lk�8i��ո�@�8U���ݶ�Xι#�Cpg�i/shmɞA�����4z�K��C�Ik�`�q���>�G�W��d�泒�gf���� ���yX�-5��ʵ��NH�g���O���͖9f.i���t�ј�
P�;�R�/}��V?�K̳h�ߙ�i7P�5��B��;6������e�25�oz��Ƽ�,Fr��NO];�֧����z�t��f��wϬ�Z=%vJ:�a�sl���������0��c�7�'�4��%�D�.(u�Z? ;�|�0;�����J�CQA����oy��`�Lk4�6�ut����74z�����^VFsޝ-��C�m�\I��yn-�	3c=N�rv�:q;9M���6sMv�Frik1��2��bj�f�Cf	��_���a������ʷe#ԴWU��T��}U�W�%��)�p�g��>זE%m�	fgm�/L S����Z�K��uF�V�k�U���%��?�PH�fpH���Չ��g����8V#�I������p�����'��ga��i{�T��(�)��6�D>�^���A�����N>ŕa��)���`�j�oS�0&����G�'���mэ7^�n�s�/E�Uz�zV��O���@n���CgVou���pF�E�z�� �U����G��X��7vU���X
(8P�s��ӻ�D��Ժ��3fc����~T����8a=��c��/��KV%�t����K��]̇W��Ę�-4� �-�,L�(=Ț;�
�hg��δ����1�����7M?T{�*����=V̞> �J�x�/j�9L�>[N�h��E��6�K�ճƤ��ֹ�-�݋�`v��j �*c�B�e��c��*��|�+�����wR+Lm^*0i��v�����P�/(F�QW�Q+�%�h��鎔.�$����˚IO=����'u��le�8o]�[@h�m:7�	'�+�4D�Vr�ku���ij
�s.@��r\�=x�����F��	 I��*\J�owK����1{+�V��lP�����'E�Smm��Dtm��Ps2��]ݎ���r��+5y4ܿ�c�Zl,�K�87�Gg��Z
��:;�V�U�����Rv$��5�-.���O�GB^.�Ӽc���_wgv梻w�(�p�3��Z-��',�����4b8�{D�`���"��������9������d딞�.j�- _WM�[C4��1�Ɇj��H;v_���x�FE�v@��Z��"�e(���^�����fs= Hb�u��xu��ߴ��[�ٮK��5��ц�nv�m�*�/������c�1:{���g/�Ф�d��Y����ӻQ�-\�#��8�)Y���j�g4չ!eK�h��)�)��i�ԭ؍u).�X�ڠj�Vm-r�V�O��k�EV>��[�#]ݩѶpdqQ�̎,���,u+iC�&�<�y�1�F���Hgsӳ�(O	c���:��	r��Kb瓟�����?y�"�RL����`�����x�u�	�B���&Ky&WHJ�"�k�A|�ŋ�S=�1\��{�ͽ��
]s�Y34ܩ e�"
&ҳ�d��A�a��'�P�ER�h9�^sҤ��>@	�e�	�󝑸����R��F��V���C�b�雒�d-���]�=���gPvc�=i$�g9"�$S^2��L�s/.
:n$���y��L@�M�t�-p�yV/�^W[)ֈ�pl�E�J��b%V��]B�m Z:.�4���9�,�5c�Y��O)G2H�c�;zHm�f���;c3&�;p��d}F��P�n�/�V�މ��da������٬����+9<��,&�պ���"<����sso��݀�1����m8�d��)7��Vq�b �MΗZ�0\ê��dt	9)$���Ȋ��S��Q���ʁiT�͵�ˍ���:M��5K���c�������:^�M�;Y��8�b���#�:��B�L"���&(f�6�Ҿ�Y4���U�W�6+E	L��y5P��6�����a2�2�U%`]V�-�,�kb�>���a�;�
7u�T[kG5f�I���E8a�(��� ��P�9��u=]t�y)�G9^U�Xƹ��Q�ǶI[+�l�6���wik�	.ɏLݩ4nm��,)gJ�o��v��NB��A�}�y�N}y�%Nq�P��V����3���7f���T�ޙ��;�jXn�^��N�Am��p:��pF$�T-uᵤ��Z�ê�4w��2t���9�Z�����޹�e�K���˥��2�s�]S��k7�z������6��9��PU��Xo��e�I@FV��٦�0><ט�sɋ�����Wxv�}Ht��\7&.��j2�62���a��l=o�;�R�:ҍP�~� �
�*PPDV�m��H����PT��+K
	"/樉���T���UX6�E#�"��6�DbV����(�[V�F�,�P�j��YQ����iJ5DTA�,���Vʖ ��,̪�"�1�EEUm�̸��l(��-��V
0DQkET��5*��U"����DjV��[��R�jX*��lX�E*PU�V
�VV-���2�TQV�[J´�6�EP��*R������Q��ơU��*���J�F6ʨ��%J"�j�R��**Q�h((�[h��&Z����"��ڢ%h�+EдjZ�EEH��Akb#[aPDXХDDE��
ڶE
��U�2���ŨQQ
�R*ʅ�#
�m��D`�֩QA[kTQ-������ޥ��jon��9Ź݌��K7���W�<�蹊�#��{9s�:��]��N�st�z�<-��ׯV5���3EKiZ�S&�y�>x����0�������l[L�xi�Ѐ�bF��K~1(���xG�fn�����鹫4XǓڅ������;��$lG�wF�v�Ǳ�x@�<�5ީF$rI=˨-�.��W�Co��ƭ��a�#����dl�]@����H�^+�؎/L�ׯ��؇�(͖�%�������Y(��(ݻ��{��(7�A=�v�#"ә�uZ.���ZwPE���(�v�V��Um�_Da�8F�iR�tG'�ySM8x��"�_mLm�I�� 75��O@f�'hPէ�Vs�;_8�p)tYq:Іn�(S��-��IV��S�T�G	�#�=c�/K���|��.��+�1V��T]F��B\���-(��w��C�� ������K�r(�U���X��<+�ퟸ�ڷ"�mV�û�g���{�A�˳F�J�aj�ʰ���yp;��q�v���*����hS�3'��4� M�֫��f�nf䀣�Plj��^�!9�"8���+`;���fgvX�)6j�K���A{ ]�W�-X;J!H鋌2�4j�=�i�GZLM�獗�ޠ,ѩR��
��Ȃ1vua�Ծ�J[]�WTn��e��QJ�������>]�ͮ��P3q��Gc�b_]9�|]�ŵ��W�P�c:�֌�e{*(�+��bֶ��t����h�3��^��Y+�c4]=��Oi��%@�qӯtqH�c�ǅ�o�_vE�ٗ�g���\�Ε�Ny���c=g��]�pޓޝhrBXWi4'�&�#�=��ED��B�2�A9׮��vK ��p9F=�W���i�M핽��
�^���./��z�N���&
7L
�
�:�Q�\<����x�j�]T�n��R.�/6�U��֌���ᒫ�Ϭ{�-�����ܢR�*�2yw��}/�D�gAE�n�Bs(ϫ͊����iR����r����� �<���R����'m����*d{I�\�"E&רt	+T�����k�ݭyCR�m�r���M�;t2.�:l�E���S�&S� �G�P�vWj���gN�g�/gVX3P/V��=��J�"`�\.- ��f����6Ð��NJsKz'�>�"�˭�Y�8i��j.$\f�s��4@��oǵ^5��<��X]�Oi��5p�-|(�>�s��yo�0�]F1y
]k%L�92�������yL�el A-g$���~���;�mf�L���x�4֪��j�s�9MĦ��.r���7���2Ik{^7q��4�	eGt�T�a�w��:X�Z�k�E�5�Ul�7�vw�{��ꯡ�q�{��,I�u��ygX����}A��H'�ZD��e�{f�z厜n���r��軛n��꠫�5�,��MXM�#$���2+���ەq� Dm�CK�f%wv���VH�V��\N��t��5V��X��u�� s�#���N��$������b�{�����g�{%���ڴ1fX�cy,�d�1���!�8d���HBң	��� ��<��Gu
㋠��騳$_&Te��cv��lk���L����u�eg7Z蠑�껷���p��0g�kE��[��<\hf-_"C��%<�X�:"�8����c+\ŭ��X}��5�G����e�b}]af�=g�t��Ab��Cg^^���mƊ
�p5,�$��L��<���s��zn;W�O�o�@���:�xeiu����첲3;��&>b�jih:�Ѕ���o��3�_[�ک�6dy�D��-/U�v����������L�1M�u��r�dj�\�d�Դs�֛u�S�\���ab���k�D�gV��<7F��dMmq��(���6k]MΩz.���%��	�9�`r�YN���N��'vRS7��O75���g�l��]A��ޥ�/�?��Ky&��ݎ�t��R{�:O��ʡ������
�꯾����G�����f��o��0��Hv"8��c5¡q���[�H�ξt
z��/���v£Ck$��ƹd�k��lU��q�Dq��(�'7>��	8����ft#�Y��S3²��e�D!C��x9�T׉a�-(g{�%J�=���$`�M	����Y�CK��A����S�q���V�:�2hG9�O�x�#f@s��͵C�Z(� Nğ��v&�T�4g2�xP�r^)ˬM-՘�|���!�拘·[�$��R�z6\p�#�j*�N���n���GZ~B22�ߜi���͉bSϊ&Y9`�Ј�{���_��B[ٝ`��z�y�@3�*���Q���G3[g����+�J<��o?(�{��ipr�I�u�����^*Ϫ��A�9	X*[����g�3���<^�JL��IS�����-zm�}V��W�=��]�'��!}����G�䥏�?��5ҭW���,RM�ޭ����;'� �LX�p��'!�`��3�ㅊ��W�� W��hx^����*���E{-4Ф�
����v��tmՃ��ɵ�	�k�ȍЩI+@A�[켊���q9���
��w��fvI;�Z��w���#\Ŝu�D7)t ���ώ��C5S��d�qz�ҡk��,Q�"*[Z�&�������ey��UT��/�h�8�Q̞ @����`�+��G���A{�N���ו��(|�Z�Z�����&2>�C���F)��:9[��T�z�9��^�H�	�a����+�����V����>������"m:��ptCr�u��Vᵸ���P6[<�V,�[�y�ӿ?���k�#t���tU��į���G��[�:�G�F*�F�N1�6�:�"���nV�'`_;�k��=[&x�Y��*\ߢ&�U���)�X�D\ٙ8�P;cb8١o���a�k�cOd������:_u�������3r)��.>��#���q�lG�{Hៃu!��˴���y|�>�s�"fr�]���j��V`v6���WCC���H>��wU���M�5��N�DɁ!�uFob����d����9{ӳ�@���
��;j�6y��Ԍ8y�N���8V�)ѻ{x!ѓ�*x��|`.�K����*ދI�|���>[f���s��؇=NncJ��X��@ѹ���=��ۨ7-#���y���A>����޼��~v��
F9BF��&e��T+4�f�v�cm�����9�c<90�;��P��E��ݡ1V�^�1�l�c����κ��a|����X��3Bx�Y-A:`'g4>�7�o7��o32�X7M�Rӯ�Ѱ�g�U1}i��&��{�ϔc������A����и\�潊����V�p���!=E��B�r\�~���ҫ臫**Gl�������;�O`��1�N�Dy3|eAfS8hs�,�Hqo`��u�l%D���XK�]u�N�wO,��Ͳ�Ŗ���Cc����Ha7t� �5�A�{��T�~8o$���k���vp���+`�$E�b�l���Ȧ��lE{r��t����|��DlCb�cl}�� ^]e)�����x���h�n��-1Z��vE�嵫�����"@�鶴���zO!"�"��d�~_�=�J�]�D̬��z�����gʸE��ɯ�_/�w��O4��
Z[���iA@z�w�a��K�9A��;z򣐡vc�"$��9��g�&��L�����u��'����De��OU��кtθ���c�ô1��ȯ�w����y��u޹��[���G1m}�T9�/��,�[~]ƶ���`�s��/��Ь��� W���L]����{,{%\�u��X王���.g9���N![tu��\"���W�������l��mg�:��X���^&�x���]7+!bmk�3W��6�6)��OI�;p^Πu��K�U%�S���T�-�:��@�ɶ�gQŻL�'[�Ӛ����}�������Q3��ZLN��'�[˫�IZ���c�2ڼ��&x�eJӉ����s*�'S�56l-x+�@gGцyp��.�]���=�{ޝƯ��s��Ns�!Jm!�ۚ�Dq`:�#���\mܥ�G�(�ki`��݌�zC����'I�;�(��u�b�2M�#T���ȝ�g�li�b$��1ІP!w,���䄗~!P+�3��>��;ό�g�q�m3��>�"�.����a=V��&~T��%.�t"	�R3j;��8�ZO��,����<�u�|�׮����=-_�s�FR�VI�j���3��P�^��+H���K��`���m�u-Nr�����A"���QI��^���W"I�'�~��z���6qcu��aY�s�QmD�q�D�����f|�<��|&9h��3���0����g�,�R}�+�y�hO�>Ы���
�|
�u�n�J���[/ՉM%�s����뮤�y�7��d1G�f7Bm\2]�:��|��3�l�Wh�ݺwN�V�<���k��g�/q�.��t(d��+�K�r��y�k��{GuG|�,ss
uNvm<W�%�0�!g*�Q��
:�01����6��ɚ�۰�O��܃OD\�EP��<�&K�L;�[r»����6����<8�\��]��7��y�m�rZ�*�ۿx[�J�N.�����g�?�,;����>����UPخ~	3ب?z��o�&�9nF|4z��F>y|���4��<���`����q.q��^���7�p>F�_z2~�)A�s�s���ܤjw��_=���dn��ᗛ+V��F���b]מ�W4�`�;)� �l��U������Z�]P⠠H�p��4J��JNdk�rdORX���k�@--b��|�o����l������v�|���<i���+[/M����Y�V���\]�}6*�Y:�2� 3g͡$4�RZ�ft�*x�����윛�Su:d��_Pag+��j���[n+�?w(K��@뎤�0�ұ"Űi9��ڥq��S14�ϕ�k��;����č���#����Qhd�bBA���|�ɫ�VO;��2l_�If_ܧ�f��P��#�.c
���D.2qCW"srgwy߽˰G��S��!��������-]�Sk1YG�H�e�����x�>GW[rdk�*5v6�JM6�ϼ����:��ٵ�@н��炏;���i����@H9J��zJ�ʉ�:"��4��wi�M]�l�h�*�9Wmi}73�-IWtIS�+�f�{����;ŷq��{���அ��w����
��v���T�G�_]B>�v���kGm��s��eq�:i7lv_L�1��n��Y��b6,#璒֜.��ӊ v�
=��5��W���Z�K'�ϗM��w�<&q*"��}&����@�J(��Ȁ��:ǿ{h�B���1�s��<�v��s��+�oN /O䯹�������=v�y�p�{M��]f����Z�s��a���ť���XY�S2p��q��{<:bC���F�uy�X�|�}�$����o� V���G?�;�0�M`Ά�-.,�,���c���ئv���ok��Nދ{�r�U�}"#��\��G�:���V�yTY�y
�!�׼��%���3dE�����[�Vq�ٗ��l邠���(F�QW�v��+ƴv�Hvg�x%�:��皊)47�ф}�������;$�G��x�*�ք+�u%�F�HV����$
�<oh�k���k��o���6�3f�[hh�9C��OJ���G�- 1���PQ_3'W����խ�ţe�_�v�ܝ�B<8r^�F+\nҀp���΃.��Uus]s�z0��G�-μӫH���3�#�uM|��;MO��r�޺[ �M��=�`yB�iap]}��5��2�q8��0A��mw&�ch�����7����X�R�_7���zY��R��֚�{�!���xo�u=*��·tmjJL�+��a:�����.*j���.�W��;��n	ʞ�4�
���Z�J7�¥}�p�� �(�y3�P ��z�|G�U���T-�hEFO5_'Ӆ=�6�
u��������Ǎ�r���2�Z1�U�G��5��-�S��\-�zp�K���zb�^�5�����T{�*�̅c�%�ԑ�Y�?���iU>�H_�ɉ�׌r��&��cgZ��o"O�g��[XAy!%�r	�3:UD=YQR;h���uP2��7~��9�#�<+��l�V��Їo����,�TA0Z��[>��PN5|��\��o������^��0�7�Xnf4��f=۵Ʈ=M��]��.-]P߿��~��^��F����zZǋ	���5Gc�2�#��aU'%�=�	�E�+��}$F}^<MXc��t��i��L�+�q���w�C"~ ��*�0&:�U���X���}Ʋ�.�����Sg]kt�Zm��]w׶�nr�DM�t�I��7oaT���U�
Z��I^�ٔ�U�ռZk��B�&X���NF�Z��m��+��6�����ㅻ��ݽmjZNIBuv��yrJݡGpVU�k����	�	D��*�Κ�6��޺l�T���	ju&���8P�� 3��{=�2�6��Ysiͽ)���K�(�$ss���m6�L��hQ�ogP�U���yc�!����xW�&!������$��@	����F#�7:7�_fu���or�g\T��C;�of�3�;5.�4pl�F�5���(tu�N'�Ѧn�ۦ��q�_H�T��;��$�"���o��hF�1Z
����SB��8���R=�;v��ʽ�BD�+�`��]��dN��-�/�zfo4�me�$��l�Ȧ�]=��t�Z����J�y[t�͹�%	]M1'�Rٵ��ȡK��SP`�����E����5[�gX�[�v#�ܴky��ote��U��kAEGa����5�6��Ӹ�=`ʹ�܆V>��n��%�SY��M:��eGVzo���B�F�xn�Ո�����.����w:��� ��۝!4zlR��]�Nw����3�R&�u�.:�=����nV�C}:��R�+\.�*�F��R��������Fif�ո���Zk���nc���n�7����3j�ٳʒ���cz}��ڹz��8oEu�>�2�B�lVv#���R���mʵY݃��A�����%�S�AG�:��]�`:��-��,Xf�Ĵ��%�//)��k�f�5�f�h�t/!qc�|�b�.w���������;�i���*�V��ۺ_Y�&u�kՒJ�>���rdhZe�V��&�Eݣi!R�h�S�o5�Yp[���(����ڌ
���à�����+kh[�މ�>v:�^,Jn�]�r˾ꂹ�ag�#�ՙw\�a�A{}��6��^�9��P.���#j��,\�]]��5V�L�}�bˣa��PۖT7�eLl�M�t����Z��;3C-�L͐m��������&�ev�m�X3���W^|
��'=Ř7�
�b ��2���_p�5�9=�|v�3V�ե�T��m��Q�9K2;If�O���\*�\��ć�ozBj1��!�=�B��s����Ȟ�`�*�)���/0�3�`�*��SR�*;���G�42�����fN��fS�c�;�N�jާ٦�F���j4��4��
�]�N���h�� Ҁ�����7�wc�nV�T*�Ș�M�w�����"�*R�+4Qecʾ��k�s�ˈ��H2T�[;� {��tPU��Y`U�,R*.������0߹���u�r(�FF"�X�����f5"ƴQAE�VF���Um\�1�����(�dU��**��"��#V�R���)eX�PřJ!���E��V" �UX��(��*PZ�,�b*
��AD�Pm�ŅjJ����DTQ�1!X\�0�+QjQ
�""�b��ET[K�&9��c�(���U�P�1**�""�YXK�b��0E ���*���\�dUb����R*ȥh�X�mV" #РȢ��"��*,`���X� �"�0Ym�X�eb�J�PU�TR(�[T�"*���Ve�Uq*��@QH���X���b����# �E�b����F%�D��ZJ�2Jڔ�1Db�FزШ (-j(�Z2Ԣ�DQ�UQH"(���*[,Q`�D�/vП_@2��VQ�)�v^��i;γ����Y�l���T�A�h��3�1xaE�^�i��b{�S}wD�v�l������U%�LAe�Q���Mpq|��
��]�7]z�+���u�+��p�]�ۓ$X��_��ע�ץc���<��d"�sB���SyZv���]��e|�AXҮ�t5��.����,�.�uu��@Y�?,�h�iN��c�F��.YΊ���n���"5L�Ĵ�`v,�F�VY*3̷*[k�9!Qʦ(Y�k����lء �m0�9���v�����]��a�W�9d��2s"&��!�4��W@��H�{A�������ב�ddԝ�̝���y�Sá�&:����\�H�
����?F.����85�{N��;�A�qj3��E�E;(?X���	�c�6�:F���XZyO�/�Fʔ���`�'�9)Ζs��v�Is	��3��7�o'WE�����@�]n @�����*���v�m*ha��7�'Nmj�2�s~�&�2ؗ���Wo:�]Z�h��"B]�k�{gHűE�p.���v�Ѧ�)��q̭R���{4�n	��v~n����up*�8���S��ץ��rW)�v����RV��'pAK\*�5���ef��ᘸ�2�����8��,�T�`QS�����k�׋2f�Ū׸)GS���m���(lΗݱ҂�̽T�5zJ��U!�;NɱNj�v��w��Tn�h� �Bvl��+r�wӛۃ�/���| �|:6��ߵ0��7�Q�=5r�������W��0�·���;�E'��� a�|ٮ"r3i<s�Ry��"��l.�F�����ݑ_�u��Ru��z}޻���Q�I��@�h�^v�������̒����f���G�ӣk���<�+S�^:�u�oU�U��t9����%�dq��wjn����z�Ն�!Bz�0kK[X���������=���QKpryS8��4
�f���=�D��x��(��_A��,͚l�bG�>�o�!��5n z�~�=�y�M��V��eV g����d���/�c�x+�ܖ�����Z�@�b/�o�o����nNYJӳ����
B�T�;�~1��J����'ܿ)�`�P_��FVCK9���h=���&$Ε���������(���,'6$�H:P���K�k���%,_Eb�l쪴��X���Jk7�ʵ��:�ؿ�x��kg���Ԟ�g'� ڻa#�{��ߧ��y]K�tq�A|EK`mxOu�s9�h���c܎��3�Nu��D��ƌ[�b?^)��L�)��u ���R���1�������Q``}�b%�z�a�#G�F�ڛӮ��	�@��<���I�Sh���e��{�/d|�-��'4j���}`u�;ak��UW�U�����JI��������7#qe����r�5�w+�%`�P;(@�}�C{Hm�P�\�&v�H[�t4���u7q�!2\�A��\P��D�9��lM��:��(���3�fM�`��D�<��i���B�74�< R��dz�Cb�a{^���,�&�кh�O�,�Ai�-?G,�W�H�Y��]j~�f~�9�KS�����2VH�ZU��w��1am�lv\��#H5�2�|*x�¶��_�^��%`��̮��(�;9��{F�#���v��l`�RR5ÅؑmDȪ�18X#��,wǡ}ywԵ���%ƺ��8�t�L�V@�ۓK�z��z��1Ӓ�?��]��aB�]��ڝ���N9G����� f�,��L�d&�7��`��3�4�N΁��P�6���S��<=Q��P�i�xi��w�b�vgeu�j�҃o���� �7gj�t��'�Ξ�CӬ�^��vZ�jY�p�K�_g���O i
P6��~�~�n�9)�z����8�[p�7`6`�"b���'ǫI�\9������uG�_A9t3D�ZNt�1��v��.�7���g�%����ٞПL^��4_vP����"�S3���y��\}�B�gi�Eʈ�$tv��� 3�x��f�u�?��^�DEً���GG��;=3�Xa�i�B�]3fiƅ1��pD%V_ ��ڰB=
�=��������r�(%�3^6�W�V�=�@�(3yO��S1t�Q1X������(Z,����l
�yP��a?=[3����D��;����I;���D/N��r�<:�.%^��S� �K4O��u�i U�Vƪ4��m��D�Dy��{ke�hX�?i���Pw�'#�[�2��Gs>y����'U�ѓ�1)4�'֒h=�&;�`G���&��XvXhc���w*h�ܤ'fl�=G4+7<*c�n3�\�u�������=�.��W�q�UCry���t"�Fh���^k��N��jx-���6�M}tM��@�Z/*�8���W��|��h�ˀ��n�彏�;�gA�K�O*��|���U���RR�W���=>Q���M*}��G��F"��me�'���o�GI�j�r��$Y��暿��/b��(�~��Δ��y�T��c;���G7���[�٭���V��5��"��=�ݝ[R%�]+��YtIE-�
+�ք���E@���gZ�X�9ó�ק���3J[���#l����G[d$�6�ꋭ5؍�ݕ}��r�V�0Ki�gh�q�4t7�Ȩ&[���YNmo&��]܀b��G5e�k$5��W��<�ӈ�,�h��1�%� �(�l����FY�vf@o:�}��U4p�_t��=�W�Jx<�Vı}�*�B�$m��T5!Z�uT�úf5G��I]`by���
��s�v��\}���^�Nlny��uB��[~؊��f��Rʊ��RV�!y�!n�YF8���]'?��]���V+�D�V�]�u�=z�]����λ�̣1y�.�ƈ���)Jfpܣu��@�*�k����Y(哆�i쿑�^��TN�	��L�.f��>��%��9�n���bY����(OE����yQ�Uَ�U������(�)���� ���%�,dF�"�~up6P�����=p0�K�l�v��^�<��x_�M�Z3׋����nz�~�U��P�<;���t���beڷ�yk��ӻ\Q����s�����w��g��V�U+������7�XB�������k�ݥ45��?9�8y�p�WAb��Y�kǬ+�8��^h_Ǘ
.�S����p,�O���SWeVݠ�,�;A�al��lgYܨ�o�����J47�Ƒ��0@����T��C��&��N�Ad�w]>s�:��_Bq��n��57��Wٵ�M�[lP
G�#�q�N�r�oR���ofHU�j��ýd)�����8��L]Q��Zk�J�WWn��]�%�-��G�.�_q����W^��7��j�z�<G��i���R����eJZ�ڰ�5xC��1����-��/2u�0�=ha��N��{�.h�:�@�.Օ���)����qt'=<��ׁw�x�*.8�n{����G�+�����9�p4�K�ch�K���Ǔ8����g����1�lW[f��뭩��e�{��4����'e�4��©ͥ�|��8�۸k���D�"Q됣�9"�Q��s�pv3�ʰ=�[��E����5�2&Kr�'J	�a����  tv��V)�-��ׂϭp���ҧy��;�W-���v{��e��7���xLb}�r�P��=I�,+�.��]5d��ʎ�<�q�y�U�7�mĊ%���[���=K��3�r��rϩ�o�n�8}���[��<�r�\g5�rkzIC!�t�8F�i�.�����'�:�
]�f:v,��Cp��\=��Tw��'�,L��Y8Ez��:|v�ֻxU}j��.���e�_?1����v���	�grNd��!�y"34�V^F�V�����|�g'BX~ȸKA̴-'Q����a�o��m�,VnM7S�2Ti���:Z�K�L���ʕ:]��,9��#���;�񌕆�W����#�kDv�##\��t��_������i�C�,��j��a���+K�}U�m`���z�e���걈qwn~�A8`�B6��%��TL<�}u���d8A��\����iq�	ث�ek�[x���ܝyt7(N��gA��ʗ�=4t4�Kt�:���rwǶ��v�l�����Z��U�b�������SM�;x�D�	|wp�U�gn�c-�p��M��y������%*��g�JT�J�kbJɸZ������ʜ)�6{����2��I��d����}~_ː�p�mTӮ͍S�2!�7���k��:Ы�Cs�A�����S�y΁u�i����6q��[�؇������V�݉Ҁ�˺��j����²�d��N(3;j�ʩi;�xj��5B>�t�]�!N�g��;j ������:� ���3`>/��������Qe��i��̻Ƥ6��nK	;>��O�E�\WNGQ{6�2!wu�� do}��;/pվ1��^�z�2k�կ���黜���O�a�ݡAt�G���Ɂ��y���;Jڥm�O��ʳ�_[��|������v�-UΎ�&Wn�p��&A��ꪪ���[o�×�`�ǳ\�N��o ����&0v��f����*�S�j6��=���f��ݹ c£� f�tB��h�^�k���ɾ��}9d-��=�)O4���r*��[x��mp��1��G�mn>�M{G?B�NWǝQw!et��Q{"���s��N�w��6Qom̹�w���'{旳W �KG����Ë��0��1�>��X#M��V�x��5������Tkk��A��A�u<�_���L�7A��k��E
��Qq8���
|��d�ܵK$tN�6h���Rpz��q���tt���ªp��1����8z�w_[�A���5�_mGeD��gP �GQre��4S�:��ֱ�؝+b�
&�c��ٸ���\V�l�kj�n�v#�S#|�C��L�k��b{u���ꏶ�>�vTz�c�����%�E.��H�5��n�;�atֹ�
�o��f5�;b��̩[�w��ܱ��EFrk�͏�o �j]��l|����VK�n�� 5P��]��owf
�b
�,�qL��Uy���ù�w�f���n�Njc�8y�jtK7r��Wv3]ʞ�;� �7;�~�U��k�{���׺�a��Ԟ�tᲽ]�.�|:�`wm�C\N�#����@ɾ\Kޠr�m�����i��ZН6ϒ�h4���;r$����ek���b�E
Ȅ��c9�2�wJ��,,��;��t��=���5��LHK.�/���b��#w3h�7j���Pu^y�˩d`�,s0��w��P�KhD�3��kf�`*vc���sV�s����̬�i���+4�������)a�wS�T�x�0�ojm�]j}Wg�]�ۦ���"�v���#�U��o4����m�����7?k9e���Q{ S���n(�L��kU��/��!Wz�����;�^]�G�f�}]--���������H�"�v�_�<xi웖���k��̀��Y��n�(c���Qݐ���%@)�>U��F�GA�#1�>�z{*
���#kr�#wx�9u�$�뻫��N!�[��:wG l-W�<����Fe�Zw��t��5sl#:�U�w����^�+@a�MsM��$��Gb�)���u%A��^�Ɠ�%�^�T�K}�37�c)9%:�����մ�	�C�K&�Jw3�K�i��hM�����|�B��'&��R�M��R &�Fi������,)�WMh��J�$Øt����T*A���^ML!��)����-�A)�I6f��S�lCs:��a��zw`a	+�.]^��Cs�]�uf����ݢw�o`�,*����L������+�Яt��ۆ�cܨ'�(4��ǝ���ڶn�B��Z���j&�q��0�f�i)��e#�icٖ�Nh���R��|l���2-�}�@�[�}�A=�E֝�����:1�4�ѐ�4�v]^jh�p��<�4v\[wx5u��g'��;���l�홸���tN.r���`.%��}{�^y��o�<}��ꝶ��ՊXՍ�Y�����<��Q��y���;dtz7��R���\�G�Ͼ��񤴮R�8pa��@��'v�J��I��7�Q��
�Ii�H^��V��[g���%����Un�L�@e�<ﯫ� (���.��g���CV4C��^g7㗝�zw!&�+��K��M�x����w�v,�`���RP��F�r[�	��Eu7��zs�=Ԩ;���Үduf�S�O��
�޻5�D��ј6��n�+˕˶�!�=0�(9��X���X�8�S�V��s�k.���*Z�4�u�֒���(�Z��/:�37AOyӫ�0��:(�&�tu�fc�E�-|�3�`��Puʸ�-.�bn��R�w
Rk��~�֦�|I���O7f�X�Z�X=�0��ʼ����g�ԃe�zdܭ�XAI���(���hWҏ��J��4vmq81�I	kq�_���(�u�ލ6wC���O�)nq�H�K��c��q��S幥�v�=�ۻ"���DQ�9y8"�N^�,�Y<�����Y6���Eem��87Fޘ�w	Y}]|�r=�[��\o`��<5��8�]t�U���w���揰���r�d����v����
��G���e�k�\����G`9�vt������D�W�5$���>B�.Ε��eL�!��ƪ��ac��҆��s���
h.�j:���לB��1�5�$���ܮ%l
�U:��_3��[,ڮ�F�"Q��mkY���l�Wv���̡���zaò̕:�r�0�1��+CV�Wu�|7���`��v������S{j:5�[{�5�f���AE��A�[k{�]W���ަ=�.`�9r��Vqs�Z,t�bv�V�9�z�C�c�w��wb��U*I��I*|��73.C(XwH�vu��͘9�t5&�g�s�=�sC���L��Gj�Mu󬙑5���`�z�۾R����s\h5�r�J�_.��jS����[!0�5�X�)�@2�Cs����k=�tt���{w���v�1K��r��<xd���G�[[A�Pi~�r`��Ր��=��oX0�]c<{{�*.�X�tv�K��:�s�Z]�5��]����=���qo�
��V8-��kKj�b=MZ�vF!�/@���X�y�gfgԝ	tXu焬yKs�i}���l���N�O�-�)�C]�\ʾy��f.T�]l�X*�;[țx�z�;�:X"�]�KT�=I(4K�U�(�`܂�h���p�[s7���)A�R��꾘^F�=yX`��T�b:QaB��>�0.��$�¶:}��.ꪃ9ˍZ];�e�N�vk�i��LVnv��s�ZEj���U���^,��GB�J�iή�K��m n��խ�z�5�R{�Vp�u�|���[I�r�w^���u��Z�Wu��@/I�uǽQ�t�N�f���wͪlN��oq�!��X�K��U�U�(^XE��U_�3�}���|��y|���q��E��ō�v�a�����cQT,DY--KZ"�ƵF�(��+*��Db*���Q�KlX,F#
�J�T(�YRTETDDh"��j(���fY�ĔUQQDU�X��R)#"EX�`��F",��eJ�KB��*(,-dX�$bDq�VDQ��V(�,X(1��
(�cJ�"LeU�!X�-�)iATm�dREX-���)QH��dU����cQF2��V

�ʤF��Ab""��J�b2J�"��´�B�+DV��UQ��[(T
¥ʪ����#ڠ��)LKhX�E�
+���
�H��Z��4��ZŐU��*�V*2*��RT��eUUAU�*�*1D`�FVQ-��&W0�
���D�-�`VQU�m�D��QB�"����e��"���
� �����h�u��.@��Zp�`��DX�Խ����w�(+I��Gtl]#�d��
Ӣ��p��F,�wb��� �6{�oP���װ��ih��R�s�S��jX�S�},�y/����/�I�oV�R�O0/����O��c�1!�78�\��l�M<�iv?)5#ݔ/حۿLW�)K��]YF��ǝ��'��oT6��+����7����C�x�u.�yڍ7�{D��Ӻo��:$n�a��8M�����Gll��1��S_:��'�tyڍN�������y��{f�U�'��7�o��e�"�\���ΡZ�e�iTrJ��*�'U
F �r��n��j�G���{�Uٮ�t*�φs�pQ����2�1A�ܪ{��Zi������A������;8r�l9�2��E{���]����.Gܼ��+�D��v�fac>ҍ�;i#�g����u-2�,�,
5'�WwM�֪�}�[� ��d�\�Ǹ�$l��E�����g��U��c9��E����p����EAZ�@C���
�̺X����j�7 �^��s�w]Em����8hk�Iؗ����E�����V�74�t���=B��+>�m�a�Ψ�e�Ǡ�
(�{�g�>�U�<��7�v��&4��sEw��a�V|{P=�t5o:���<�?�O[©�����qp�{(��;�%���*uǠ��9Wu�ܒ�^� ��I��[��wq��;���l�C��8�V������1r��+r+��M�ը��C�j����9@o32�7)�
~$��xE~��)p�t�ꛨ�nV�=8���;�*-��.u���+�����&13�H9x�+�Rՠh�m�ݔb�m�KU��Î.�^mrPb����T�h'6�zF���흫��M]Pߴ^��w���я��ſ.�T�VQ��g�v�zX�i	��8N��w��hs>�ҵ�WKD=k�Q�4�n���g�g��j���h{h�T���F9f�E������b���Z[C�������!{h.���6��£���.��z^�X��Iν����I�˙�W4��hq���C_�n�z�0�Mл��-f�~L��!(�����J�IN*�M�s�H/�6W\i����½7zx>wUV���9=���n��|��n���E};Q,�W(پ�y'a��&í�P��.��t��b\6���T��@�i\��lp��06�tx�ƿ������t��`ٚ��F��*�ѭ�I�K$���ʭm��3�6Z�.����Q8��R��{۶��J�mΪP����ж71�|�7�Q��0a���oaˊ�K"�p�\��L�Z���òV-&W쳙L��77�*�U�,��%uL=��~!�� �i�]��v������V
���ki�nϷ��k�(4�NK&v!�ڦs�U��X[L+�����ţ��nyK�^K����7��bt��ʕי�{���so:��i��S3V�Wsש�ֵI���6o8�Y����t��凼@ACy�ۃ^���v&��k��G�T�E��0�a�1&3����{E���뮾�+�R�}Wy5�!�Z�c����]KFRL��灂��K� ��7��:nP�5s|Z6qG�^z���������	Y��3����5	P��S�o+"��t����W�Ii�0��9�]f?e��v�*�qX�Ҭ��?�t�o����eN�y�hA*(���]S;�u�����V���4���N�ؾ�s���ߩ!����.�+����H�圼��N���f1(�J�4<9쪜�T��&�m�}]jj���0�W��+V.��7r�"*{C���N7�oM�Ώ�VD�f�g.S�7�*�Z�AJ&onMQ7�#\r����΁^Q�������ڮj����8��+}�''Ry�tDoq��w=N`�Խ������</.����nm�ɪ;���l�O5�ڽ�%�qh����o>>��!{hq	�ҝ�ן��y�a��{-���U�zB+T���2��\c���{�pX��$�E�j�J����.v[]��N�ӋkK۔r�i��Ia��������ϭ�}��\|k�l6�Iy��f�̥�%E$� �v&<�ٳ
!�זj(ޘ�XD��iI������gv+�4�wIvnC�p[[�oAѻӳ9�:0�ȫee�B�q����2�eY1!a��������|o8�d5uџ���q1� Ía�^{��3n�%Ĉ>\��wҕ{�{�O@�]�un'ؕc�+E��蓚|�<��H��u�,��s'e��m,OJ]�䮆������h=.U�ͼ�1�vAn�`IXi|��Vr>��*<����}_}K;�hD�w����&�����Ez4���=O�@�7�W*��9T��7H��`ݾWQz�z��K�ك��Zuޒ��_�*ڧ��
�����$-�]�<%�趷�����Es���e����-����q�!�w�}�B�~�{��W+�S���R��b}���~P�TEg��7�'�v����w[�6�lt{mѾT��^��^������x檩�\�����6��׋��{�{��^)?[/��r��*;�s|�5�p/Kn�w���+�R���f���1�W�?M���]��\j���F��P_�Y^����9���|�~]K������\bS���[i̠���;�r��R�{I����or{�6���N4���w�Uy��ΣS�{R���z�&d�G)m��z�k�|���q��W�I@d�h�����R��KÔ's!��Q��c:��:Y�n`�/�1�O"C7Qƨ{t\^H�@��=�>Ń)�������})����8�Mc��0¢!��K�����\�u��:���iR�W"hm���YWVy1h����z��g���J$�Z�`j�Ȯf��t�e�l�2�$]�	����P�=x]���`]d�^j����qy)-Z�֬s�@sy=�|5Q�8tA��qj�å	ɷ�YT�j��-.������V��������u�oѶ��ӵ��kA����"�KΛ0L��1�;�t��W?sݐ���Ҏ7�f�=Q�:74nC�WZVb�wY���@=�����6���D��c�c����?d���>���i�7lt�^�QѦ���9Ƒș}�������0��\�,~w�*na2(9��䩣Ɛ�s��o)���H�qn��f��Y-���Q�v����L��==!�=$����{y���ag&aY���~�����;Μ�~=ѝA��t9����=Sq�Qr��%8�'y������&�{�u��[��]p��n��]���G�������=�[Z���WCel���.چ�p�������i��8*E�\�'���f��O
~5ȋ�j_���%5��[��-Q��r��L��.췡G�6yۊ}��e@�^�:�I�d�m|���n�4q��I7���S)�����¯s���q����ޜ�zX��۫/=V���|�h�Z�y������O�Ki�y���Q�C��xoޖr���q���h����?g1��� ��Pz�M��(���'+ܦm/ ��m-�q���Og�oԭ����$qNO	���HM����[3]��:}��u�uy5Gv@]G$G	�(:]�fG��Q=�z����ų�睼}a��ܹK����[�H���T`+hᨳF�2�aZ'�Ƥ�Oy���t��t��gh�I���La
��8j�m���Aj�A:�Z����������z����:��5j8��1����vb�1�ӱ0���(�'^~K�����oH�-�S���[���X�k/Xʬ��(����Gtj�y�U�F����>yPI��f#׭�z��xߋ�k�k��9�*{+eӅj��1Zѝ�j�8p{E	��
~��J�t���Z��M�O��o_mi^zP�tP�V]d�s�p��vc�hn��a��h��8��*���A6�d�0�u��V��V�����F�vP��Q�!���͕�:]ü�����&"�!�X�Sg{��*��)��
Ⱦrn鼆��(셒��RB�j�5�&��B^�:H���7�\*M�/��>Y��z�ٌ닾y���w�܍�.�|R�K�c��k������z�Ȝ4Z���U�G3Y��'զ�W�s	k%��G���I�or�N�t��P��e�	�WG=V�p�i����Mڌ�4�kn/)-j�i�k�Sv�nr���������Z��SB���-���j�Ah�9�]�'�*��Ǽut��z��(��6T���=��qOa���}Dm�������G�z>����y=��A��p�Z:��hdS̀`�ڙ�hnK �P\��Y-B��jVTYk):���ƎꝼkZ6T�%�\#��hGq:��H]:m�oi�5�S�)��y��U��÷<J�����z�~s�mo��:��Be8%��f��r
>�Z��%z嵢��Y��2(Z��Gr9Hj��.���6�)��3�l{��MA"��֬�Fmo�b<��X��&o�%���.Y�}��CXO��c��iQV�%5�:7����1�[׹�t��!ъ6@�j��^ȇ��i�?y��UN�Y{�7�K%��>�6)��SϪwmr�$�'�����הo�Ԣ��m��f��S-�VrTQU����f|l�h�_�s�h�~U�9�����g��ؕ�4�m6^��q�RK)Pw���;w[�V:C��8Ǣ�;z��o6��U،��-�IO8�|��R�j6c��/����̛b���`�o{�Ek��GʺZR�D㭄�q�VƮh�f#Zo'7f3�\C\���r�dK1�qu|�l��e�s��xi����4.���3�\͌��HzK����c������E���ӏ`D09oTqY�8N<�Mz�9�YB;=�}�y=����tE.ڢ�!��{$.����mK�s|��������O�#(�h��r��U�K��n|,��ۊiZA�B�w�zx8���I�W�c>G՟IMָ��>;�L7F�c9u�l��R�v�F\�=��=ޜR<����GEX�B�vQEr���ƀ�R��bW��}��h>�]K���	���$�.�B6dɛ�_'���'i;/�}&��.�[}m'n���nά@n�nb�L��Τl��G^��G9Vh�h���Kp(k�U}ZR\�g	�6~gk����[VZ�喏Vm��R�-�cV���)��in�=�֡e!�f\�a����2�2��>S]�xĖEN��rY��==��P;ş7�HMſ{�Oe���Rm;�f�ð�GR�W��f��6��EJ�>�������ך�*�[_gV�r"�6$��,BD�Z�]&SE�U��+��b��R��ʂ�\���؁h�<��y�K�b��{瓵�Y~��3�֕�p-�e��+ħ�t��㜖�c��f�.�QT�]��Ԝ&Y��X)�e�t�8��%`�H�M�z��(J)��p��jXm�v�x��c�~�T2�Ζ�T����c��h�4�n�y#�U5�d�Mf��H��ۘ���0k����1;����葃��w���p�Z�t�J�*� �(TD�'���b����S�5�v䀇8�(Ge����8�g4kD��\e��eC6�`N�����PfsI�[4��i�H��5u��V�=�.���Q�q���F���]3��'m�����{xD8�ӊ��ڝ\�n���D5�-5�)��ki_6�h��"6R0��dރ�ȼ�BBÆwSe���r�H>͈eήȭV$����tk�'{mtU��������p5�I��Vn�tt���\���b^ey��o�}b%� ~�{$��1ZFWbؓ�C�WA0㗛�0�=y���%2z�r*�l���P��3Zk;�+9�Vδs�u��L�3'o&�j�t=�� ���MW>��9�0M��H�B��M�	C��MP�v*���p�p�S�j]�(�˜�p�t��Y5k�G�1�,l�8)p�w�*�om(�@<���t�;��'��\^�פSEWoYbfi��L�B�ⷳu��ո���%s\.�����)�w��pܘ�U��9�E�ӎ�u'^�����*.����F�w/oH�ڕ��$H��e�Y�FP�f��a�1�k�Z���/�Oz�%N�=� �\}M}��'D뜉�ر��.����v��->̫�<a (ʵ���퀪悃��]��rV��/�y��oSy�e�[o�ب^�`�݌�q:v��ř9�V/b[�Ρ��L�W�܅�N�gҦI���˾z�։��uۊ�m�U^��̠��;��'�yh!:�*�_g=5�4;o�,�Fqgr�fp�o9�7�	�u��wVF�� �y)�A���$�$��j�o9.x�����g��%ݒ�v���Jk���-s�X�oө�sh)@��+0��l��-f��*C]����8�@�Σ�n�n80�hWP��:��Tvݝ���m�ݬ���9��t���]�jvv���8�S���v>�㕺4A�w��3_!���v�T�6.��8J�h)�L���Ӗ+�
!B�{QI|85Zվ�<�z��I�g�:o������Ea�WX��A�%j6q�m�͍췎�ҳ��L�]\{��r�r�p�m7*�0��Nhcw)�.�XuۛY8�MaPJs�R�N	ٮ�5�)Ѿ��-꭭�;L�����@��k���ʮ`�5�X�ovl��1�d�����jW
�pj�+kw*�K�ZX9S�<���U��m��]�<�Jv�F�a��G;���*�W��+�**�f�tBv������4�AL�i�pXDݽW�L2Q��T7t ��}5��^�ZW��:�_Sh��;�J�����꺘]�f��ը3�ΫB���`���[K����sj�=S�t���q��(�1�@�5%�%��G,y��Cil�č�gp��#v�Ƀ�YL�=Bј���u�39@�:ټ/����O4���}>�V����1Cxn�Y�(�cn�V��R?5����'2U�y�r��X�s�k;9`���ً%b*r&CXc3��Rд�޽�H\г�����E�jP�G��rYA�q���+C[��̯߳O�h(�)��h�
"��"�QQb�bT��Q1�XbT��

������R�Zʂ"0KiX���V
""��Rڈ#�TPPR,EEV �D`�T�ȵ��T*+Z+"�l���0(֢�H(#"°��VE��U�(*�-��R�
�Km�%�ň�(�Eb*(���TDQ��X娌PT�ш�"�*�Y�PX)�AYiEUDPUKaEDE��EPX�X
"F ��U"�H�,P�
��"+#R,Df%R�h1�ɉ
�Z
��j,PX�"�E��Kj
��


��`�H�TDF�*0QTX��(EEU�%A`�(�)��0�UTPT��Q`�)TE�"�D*H���߾��RVt� �3at����Kt�u���ָ�,�dv�l�z���X����)�64r�y��r;?���lZJ�dD���fk�M+g������n�����S�4�R��%-��`oeS>̥��dM!�*:r�r�e�t�2����A�&5��_'�E�)̷7���*eJ�5n���c���;o���w�3�wA�$ƫ��H����l�9�N�+�"��~�y#�|l�z`���3s�P�.��6)Z������)��L(�����趂�ϴ�Z��k]FoRכxi�\^7J��$oNg�x���嬥���6�������qM>�����ع>�~�t3u�cFʕ�w�p�{�z����mW�L���EP�lO#��y]����2�sp��1�]=O=����k��mo7�{˙~Bmrm6�����E���LY{n�h^!q�[ ɷ�l�-H��R"3m+u�Gկ6�nUwr�y߮��M��}��?,�O7]m��8z�Z-�̦�*��1�a[ז.��'G�]����=�p"Sqv��.L��TR�IM��u��������2����x���Y����-��X��Q@e'��U��++~�X7�Q�Ǘ�A��շ��t+�;r��e�"Ӯ�w7��:����r�*����}C���&�>�l6bd-�L��ޣ�ٛ%b��$��ԃ�>�^kTb\�^��*�6�s��m0όL�(�ru��w�;�s>�;W-=N��[l���}�m±�%I�B��o;V��!4�Ƙ5�������&��+
*��Eϖ�<پt���ݻ!}y;K��z�^K�*
���LQ6�j�B�Ҏ�[.��j�����i'�f���l�Ǝ�)O?���\P�ۉ�e}��wM>iQY�+a�Ũ��Kޯ�m�*_�t�v�ܿ	�)M>c>\��U��gm�}�:�c���6`7ŏCݐ�b��|jctL`�H]�*u��e[��J�w�q;�jR'�w�X����t	��P��dF�I�����z�i�ܰ�S]jh�WW�Ww=�~��s���؇�<���_i��NCtkF��)�ʾ�^ɜU=��/�k���ˬR�^r�N�tܽ��L�t�Λ��#��y�s�:���4�)�ɨv>p䮰%(xP��f�eňD(6�w�&(��a�'P��!@�g�`�3�N���na�h���Иu�7����ɓ��}O{U�U�)�H`�Yt�b��ɲ+N�k�[�5����r����4����1\�qr�z֫�Z�l����
���dO���%�N�	C�cKޙ�����ﱜ�)_�]��r��fC��:n�7[���F�_$�[vk��o�d�V��<�&m�g��f���q��{O�mywy��}-�v����=[���.���!�P���%��h�i��c�Ul-Yne�N���^�n��|�����f�5p�g�L�L��'�
.P�,b�N���.4N^f�h)+�Y��XrTRQL5��6��jkaʼ����fg^�w:�M�]p�l��,}�I�Q'ne�q*Ie*����i��C�\ҝ�ط��@T����N�Ux�2�ɉ�jX]^e�jT��&c(��ti��;kIJ��D�lY!��ң��]��y��z�ˠ]i��A��JZ�C:�S�(��y��G����+9��]��A�~�޷���X,#c����h����يG�B�^��zP��C9O����]�^����#�xr���1�DR����=v&s��Cqڊ܈O���\̲���w�Jb=�RE�{�d-���H�@��}���|�S1u^ �c��4��!�>nD��U�ǥX���!{���4.<�����ᦆ����c��UBI�/
\˼jCn��;5vinL�z}H�& ɦ�ݸ�,զe�}���w,t��`�H]�E�nq�td=j�v��f�3U�ާ%�ӻm�8���:TĆ�ެI	�O�Z3L��^����^��B�>ߊŴ���/�V�3M�i}W'!0�NpxA�S�g2D]�z��c���UO]��r6�נ�3T_i��WR�}�Z}ד�G@]5���~�U[��#����mN�W�gnC�������)[�1�x��\Ò�{��v�|�gz���y�Ѫ�緓�W!�B`�r~���ݔ��$҈��8�KŪ%޺=C\;/��k�Gc��k�����.�i�/!t�T�n�4�o�{��]%���/�C�ٕ����M��Ei�{iz�<	��z��T����zm�g���h�B���F��s��]I�L��o"�>�k{*�>�*Z��[[�f)AA��kb���L�spx��%����sju%�;�!1��]l�V��]լ���]Y<��ǵ}���S,���|�/�'_��$e7�����H��M�|�q֣Zq�<�Jئ�o��Ȭj.gZ���r�}�euD0��}lL�lC>��:�Y�>��؟�Lᙳ;�e{��c7Mۜ1�i��p%�)�
��L4�C9�T�v��
���MW���.�Í'�@N'�G���/��_x��J��h/,��1S�U%�9�<LY�Q��
�3X�\�O��U;�j�P��X�kL�ە=�LU�s�O�n=<�{�|&ҽ�8�Q�ʾ9;o��yL��p}i�0;	Z��O5\�\E�twCm���5uA���UlV�}eE�=0�1agj��w���"�	�w��m�|�)v����/���m{�w_5�I'�f
�|ϑ�U[T��߇E������Wy�k�d�q���y1cP�,�h��׸���,M�چ��}�P\v�)�}4}]Dx�=t�_���{��CD���=(_(����]'Hܑ��/{* ;O]
��K<�4��;�k��*�"��]��<YZ���q��+��;6e�&_H�5�@ٲ����(T<��$ܥ�^6
��=�1^�uc���*��y�ZZ������V�j���lϷu�X�l�ζ�<��bE�Y m�]G'���X���2]Mr��y�i��cV�e�VB��iI�Y�&�*7����S�h��Y�Ջ��=+���*[�*o����.w����i��l=����i���̷>}��f{�C��Ρ�VQ.B.7�8y�y���3��B��u<��dŜqW���ex����pZ	׿T�#�������}=k^O}6E�\X�n���6{�z;��r��T�Yٗ#�'�<
�RT�S�e��&^z��%n��gV=ǥI% e؛�L�1@DU����sKDd���]Q¦�"B�a�߇3}"���/{r�J�7�p;�ԺL�u'��b�r5}�����/��R�Z.F�n����û��'v�v!+n)�Ւ�NMn%���m��e�y��������D
�-;�U�7�����^I�֕Xm>R�������̠�Ю��2�t;�4ȫ��lc%���-]*뭶�mnX�m�jʷD��f�sn�O�vֶ=m�Ca��JTOWc�Ne�>\+��:qAI��PueZaoL=�2���0!�]vj�k�>�����u�Չ�7����J��Õ��Ff=l}�!p�RL|焽�~�h�6����ٽ<���~n���K�8γb[� ���N�Ut깵�^c����[���w�_��`9�w c:�ɑwOFf�fm��T�7��VT���=|���F兪�j�F5��n�m`�LmU��#NM�����T�/�u�yA��g*��+��ZٞJ��n����&1���U1Or�d�s2��擯E3���P���[OP��D~y����/V��UT-K��Z��SvQt�K����q�����5j�_3&:��[��ܛT<m�w���!v���MG�;�aM[[t�0Z��'"�הV�%o�^���;���f��r
yA�"�Z��&�cwYlQY��AY���%7�Mah}�ΥP��:�gw��r��Ö����p�!]���KU{B&�2̯,9,�)*g�]�w`83A�4<`��4jeʑ��l��-��Oj�me�s%��]�X�R�t��u��te��c�9���E��im�2bco�X��<Kn4[ѾPm:�y����&+�/�Hun�����U��j^�0<RJ�Wm�7�������������y�IU�w���mI[эm(�fĜ�l�@�uJ6��%&�c1R�
]b٬C]z�p'Gi��ӈʲbBéV�+͌�l1�:�q�n����EP�nR`�g^�+�9۶�(���X�a�M���c1Wmr�c����cN�𗣤��+}c9�]���.3;��ў�-�'-��z���hq�����C��m���O�N"��n��O7	å0��������@oCtC��Lmm�����
Ӳ�p�����Q�Xٷ�Ӣ��Cn�ecj�3兆K%r�����>ћ��bw$��ȅ���ym0^7R.�v}Wjj��֓���hm��5<ut��z��)���� 5*a��ũC�q�>�!j�aڸ�k-j}�[=�?{˥ߎ�r�)�o�W�ٝ�h�7�����8�������y��=I=a�S�[�&K�����vP�����+���"����g�R@� ��� ���+z���ָA��n���]�m%H����,����Nr)de�:��5�v�;jT��p��������!h�Z3���������3�b�ͨڪ�y�^صz	��W�mUf�M|����(h��(�S����T#����������2~�]�h�m����ZX]zT�w�J�uyF�	�DӐQ�R��a�)-�eKg����;l4Q��ik�[��*g�ѥ�����C.��(���7^Lv��,�%N0��.d�U�*��
����u3>�O��T���Q����%`ԉ,؛s�C9�����!-��8�Ò���]tu;����C]=���\�g�pZ����c�N�NtT�y����B�%��
��O�:(����H�]�CX�����c�Z��s�t7c��<��˶�s�ԋųj7Qڵ�U!Y�K2���a(�R�(W�[Z�P�ri�Fw��ڂ�����ͮ����6ˉv�۽=\7�܍�[���Pr�$ը�&�o\s��Z�-�2xg&�z�m�Qs�pgTُ)%*-�����9`q���Cw���⮗��r��)�I
v�`L3���]��n��`�ft���;b�-�̚ȹ`|��/���7ؤ�����v_+���e	J��כ}y�WN&��h�e�i���سk+\u�J�k����Z�[W��a`�oz@{v�=g��l٫��O��[\�oIr9V�z؍�:�����irx\���4�߽��kB�(�ߝ��V8}���*���
���"���=~�)�x�o�Z~���E��h����~]�/�����	�4`����飽d��G�u��Z�(;oUGi_o���8��|���������i웞�JQ�ԝG�^�(��9�^�1x�ᴯ�ڽ�A!K+�%��(�_{�z.�u���!��͚l;�����X-�Ǉ+s#�X�޾� ��F;˩���Bʦ��8k�2In)V�j�ʸRR���
c�v���3�H���utf���6��7�����Qbj�����[E�f M��I�ђ��My��K0ű[Aa�֣F�#kTP"&��0ꠡJ�n�8F�c���9�űٔ���LҨWr�ew5�v�W�\'+ǖ!{ �Km<Qޙ�5�(v�6��]Bͼ��qΌjgD��;��Y��%պ�G�\��M\�P�n[����U����Z@����]Ο�-�(���Ђ�_h�O����q�N�3�`�u|ƶ���Yۖ��N���z�����R� <�nh��8��ې�%V��Ki��sT�3�3�������q��c�ۭV< ��b��v�����2�-j�WvJ���q�7�zܲ�¥-ں!\�ZK��a'�%����n��4]�o	z[�����t�iԝ[�(;��6���r
{�,n[��{C��m���j�1��&"f05ȳ���z��0
O;��L��_J��>���2v��\��֔��w)��R-E�+����Ȍ1G�g,�[�D�Q�_\N�3�Q�+6�m?�eb�R�&Һ�h���w8�x�ove ����L�w
K7�x��:��|Eg5-Ab#�;�v�{�.+^�ǳ�;��Jq�o3[�-���17��6�8L盽�+��@�����13:�ۮ�;�p��K:�]���l�u$;f<�����ە��6dj	I�=Pq�f$�̩ٵa��.���������Ǒ=���Y������m['�|��N�i.��U(��ϋ`-� ��H�^��i5N֏Pn�h9[�d�@��8IS ����s�.�ԟu\[i����z��NL�..=J�vge���;<Ai�Z�H|��9�&vD�L�z�--H�<<��=8;�mt�L����v�>�Ń����D��9P��c��w�������s񼘮�&X�Ԏ�y�'q]\�H���7���ѧ�e�W�@�)��O뉤�|�S��o6�eK]�S��^�wK�*i�q���.��2�N�&�+!5�x��R�5+���>�Dք�`2�Nmv�lͣ.�e���/�@]�����=9��g\&�����s�Q�b��y�i��1t��{�a�����6�i�ج:��)���B]p�ٷ��F��2��讧��s��Ol+x�}�+m�։��ԕ����f�f�(/f�Y.W��=��7w+1r:`�pT�wA��ኙ�I�c���$ <T�]wA���9��|�g)��g����p�\*��nG��'.�Q�8�(�\[:(�^cGr�X��͛�v��-�
¹Muќ�q1|d(1s^���5�j�����e9E��!;�:�_cCv����"9^PD��8�X8eD�1W]2AN�5p���;�߆ܝ�\��,v�ȵm��)���Xo�'䙥=����+PߴmI����̮�1I��X��QO
���M��Y�J�|�t���I�:`
���Җ�0�r��O���o�T# z���̰�I����[P���PIH=�z,|�wmn���cV��m���8�R�ءv0m�|����fT�ڀ�YQ�8Ҹ'L��5�3�!�7���6���nL5
����YE�.u]ξA'����#�Y�:�se�g�3��*+��0Z56Zj�����.��u�!Bvg�y��D��PU�b1V`�
D`,FR*�-h*�))�����V"�PYXT�DH�0P��A����H�+R)F�QdR*��ł���E�J,UAb ���70��1
�#�beh,�6)�R,4��X��(��� �H��DdF+#mT���XE��E"�X
B�,X.��
���5.�b(�`#dPTV�+
�GT��U(��+"�����XLaDEE�!T�QF��D�ɉ�Eb��1�"�E9JȢ�EA`��*"��1ch
A`�b�2

��EUYP���b��� �`TY�d��eV"��E�b��U�
QxyF ������h.�f�n����N�)aC:��kD��R�$V���V��).�׵�\�}�+��x*��r�����zw ��lV�>��(��Rl%[�Ѥ��n�#���=�4���gl���3���p�V�R�H�>
�U��SٚT恆C�1�����K���1Q�*���:Tn�[wM��������h��a*t,K�Ե��9�����i8h;i�}��3y�{�~����]��M��fө�8/�YCd�&5��B{r�R3|���ٽ<�_��$�9f��������r�2ϋ�;ϫӾ=���'��ߨsZ6{~)v�^lvD�������GM.U7%1�c�S��a1!�}S��O_"kX#ojbr`S+��n���9�0ֽl/e��61��G�i*fJ,��/��l�uw?g.g���֙�鉷�f�S�P�:q{~3��������^�������w��z��W`� �ʰ3�����D�-�3���s㋍�:�q�����l����Og��7�6L�8ɛ���9Z��BV�t�r���e5��H��@��{���`5�SN�U�hX�g�	q��{wg��V=��l=�k�%��vL��N������|�`CTV_��8i8%��D�8%�����nѾ�=�k�lZ;;�Sg���M�n�>�˼�k�/�7���w�s�#�������C�F��ڤRG.R�19��+��HQ�~�����s��nz�VU�iV��*�0��^l	]�9�R��f��%�ޡ-S�Ϋ�y�=�Fjs9��9�;����V�����1b�a��t5u8�4�\������2�쨏>n��$n�����n��ۅc�zT������l)Y��=,�>�Xu�1�;�*m�.Y�N��I�Ė��h����J'i⚑�V�=�=���s򮄿��mw��ًI��ut�d눚�s��c�S�P�I��1������+1�9�����t	֧r�uc���7)�A�(t��B}n��r��RZ����b�}����8O���4�����e��2���a��NVu���#�/rtc6�J
�bl�մ�J�5���x����?{#��k�6��5���a/$�?N��]W��v�u�w�eג%�>7�ʶ��l��<U@��DV�,m'��Y�L��{\��}�r��d..Ru;m���\���2�+U{g���Ͱ�_C��;V�)�YY��&�oGSRL�
����ȫ��W"��]p��M���l>;�������}�U�1#g�{���>|P*�/�;=ed&�8�M��N���eS�]-��}��]v����<��Ms���_�O �5�=�j�zX^Y�)����mw9��3W�sn8����9я.�>���-#ԷU(��0��#�
o|R�T��5�>o{O5䡩P�oZٓ7j���r���sT4?�r�R�#nw�dt�Z}t6�����9u��]�L���57Isq�Q�XU,fve�>�`њ^kI��)��#k�g2�Yb6a���Mj�,L��m�a� lc�nᗯ���<�F�ݶv#2c�PR�����3���n�n�;Kd���q ���s�v�\�MQA��+�*N��cW��<5ޡ@��L�k_��b��u�M�ׇ3nGǨ�D���Ok9[ǭ�L����UeSXM��@��)V��mN<�p��9�.�RԒ̜�NN���<�8G1F�X:V���E�'Jqq�9�0;��y�|�� ʘ"g�G>Z�9ҵ�f.f��%W�pҤ��P��j�v'�B����=�-.�4��cӝl'ՙx�ouH]��.��劣ꎍ4nO�9�(��`�b�N[}J��`��օd����IC|�U�� ��&�/I��>X���hε/'��e*|�5gft�p���跳�6�Ƒ4�qS��[��:�����yi21��b���c�܎�m�Ɲf���'e[�<B��}�������[;���/ٝ�g���*���Z�VMЊ$���v�@�	�_{�J�A����o���E���b�y��i�� ��JϏmT�����ō��V�R7�ʂ����2�kۢ"��e�b�&1����Noxd���ir�{ޛT�{���6�g�奊U�7���9�H�o�V7�P��Wo˽����6�/���������]\,F�C�7�W�51R�h����)�iAN��(9DwD��{�7�w/F+�)e���ɞ�ј؎��z��r��W�}݋�����t��:�ǵ76V���ڇ(.���1�8ڼ;ύ���S�D����Ɛ9ъ���a���;�`m��9���O=Ρ��W�t��\����i���ݕt5�lO�I���-��Y����Y(}�ٮM�-�k����=GX��-S엏�5�-��͏��;�{|�P�{rVI�Tg���r�^+�jk���OX����������y�:j'c�����N-����������m�ñ����v��A�q�U(>&�)���c���0����F��ˬ5�QjD�a�JS�Sn�4���qm�㚼k��<�"X*�l��zu�� �T��\�>����N�B�D��,@s4�y�c�O��uGF�OrWdK(츑W�v��3Y�z��]�!�:�]���a�b�u����1�b�`O�Ϗ/eO���vC��N{5��]�'��I�k��h.�t�&5��]�*u����Z�!V=PN攗V�h���37��q�0�q��2�?����j�%�� ���g��)վh�J�s\����M�b�*+3GX��Hb^��n��c�@�����F&�)W�Q�����Q62�I�E��������v|�9��Z���p�ǺGD�Bv�S�'��a���MMQ���{�#�3U�>F�,{�f���T��7^P�e��Q�Y{�l�D�|��d
������췀7�W��zW�l���Q���>k�;���^�	�k��<
]K�T�VU;�N��)f��eGk���gLeQu�d臙�!ώ-���q}�ew�g�Jw=�o�+�Z�����yF�D�Ṃ�n~�qY;"��Y�WZA��`J�r�zh~:��qz��~�}�>����rT$.���z����S���r�[3i�n�j��mQ�6����F}`����ڥ�bw�W_�m�Nad�=X��LΧ�G���'�W�#4���2U%,���(�ԙ;�2�0��L�����G���Z�f�����7�\���s"�b�Ī���Z��r�]S,���=�&vV�RNl݉�(뷡�0'�:��XĈnd�/�D���@��1TZ�=t���>��4�eM���2b��v!I$(�a����}ø�nZ�4XO)�N�%vQ@��j�"u�M���
J���][|s�S�֬���r�]:��^
�\�ڼ���S�R�Kg4>�7�i�^v��9ʎ�lf��.Lk������q���ɾ�����lt�r��������i���F:�a��ܹC\K*ZXg����zv	�X�\���' ��zP�n�����ʅb⬒:�HB��.y�}�ҽ��1E퓖�)����گ�`�;;�w-�&b`a�=�G%ڒS��{���4�\���6��
��C�d��2W*�ļ2Q5/���M��7J�9C���n���j�����x+��n��K��Ҩ��o/%�[u��Q-��-
Y�6�j��m�W,�ej�Fׂx���sޥ+�٪�R.��O�7��wX��]��Ôjk���>��xvV��-�Ƨ��0e%������$�:����]��.y�G*�f�_)�n�h�"�b�b�JR�,�5�,��nCRj�D�(��ށEWXJӉe ;���Q�yb��-4����,��{vF��GU\���&��h]���&�u6�����ж�����q�Y�cgM�{KL�����5��ѝy��K���Ԅ�{0���ܤC%s�h�:��f�bW*-�\5�i�+�jئ^�L�Jv�M3d4ِ�[-Kj
��5�P���/�k�4����SN�4�w���8
�PUj���O�{��ݯF��� !��\��ډ��Xt:웦OL�����A� k��z'�Lh}���m"iv�uL����t�3g��Z޸�z�Y�w|=էMz}>4\��1>Ɋ��w=��Qk*5�=�nܩnnK4�;�E�X���i��E�tq֬{La��:�h?O�0I�Wq��/עޠ-��m�/���";$c=����+���)l��?
�4.�~Ǩ��Q
��=q���v"�)�V�t�nm�1`M�E���Y��
�l��k��u��=P���� ��z�	�z-�E��N+c�O�{�%R��g���OU��~���+J�^�tKϻ��t9l�;Tw�{n���ꃇE/�"0L2�k��ƚ�v=�Fa���U<����L�w��s&�)�����.�L�꟞ó(������(�5w!�ד�Z^���?d�{�Z�5�Æ�y(�`����snJ��f���i0(������L鷼&c������f�B��VSj�\�#�{`*�*&���RV	s��s�Ы3�ͷ�X׳l�6�Ƅ�'vQ�Ox3%��S#��_6r��.��ooG9�	��S�׵��j��Pѝ,�!��SW+y��o@"�g�+L�ߤ?M��3{n�d�>T�q��[[���iS+F Y%�ײ���2��6��G䢽��֐��rO��ۼ�:�1�੮���=�VN�GU�����z/�l�O��E�i����1y53ޭ.�{�Tu��:}"�ps�\Fp��T�_))��Ҟ#r�����z���sw~"yJ�󁳀��[S]��U֖�n����ƺ�*��ؕA��t�X��wQ|HQ�:�̨/��Q|~�^Km���F�%��N�4��x�S]��n�y2�Gw�/7��6M��\�����3f��\���XNz+�\L�O�M�1
_��T:����&�`�ݴ�ht�3���lcϻ������;�C|6�.l\u�����j�Xi�~@��s�1C�-����Ґd�ћZF �#�ԩ�uʑ����Ib�pGP�騲�`�46�OJ�㴫�ѭ]��,����0����s�Ů�����˧�ܦ虆�`}�ח�0�[���C�t�1�����;h�u;D��J���{�%���0�����K�����i�fV���w����ꫦ8�T[���J{	��C�!�E������� ��w����C4r��9�w�+�U��������9�`.a�Y�D��e| @�?T�B%���F�e�⣈�-�\��֦$�9�/��ɩ�<\w��;�2���D��	 =X+�	{9*�?-��"ʸ��]5>s�躼[��izov'���}��$�K�{f=�
h�s�����%�td
5@�Op0��"s�����"�v<E����c�hq�xъ�[��� � �jD'��/�;u �u��c^�e��sq���2R_�F��I]�u���(j큂}��[9�)��X!�����?��c8X�HT�掝}�����pSgG8�˔��[s�]9�\a�Aq�h]Ͳ'�]�Dd�J	����e�$^4d�K5B�ƅ�'c�sے���~H�~��Hv�Zn�^4d!}?v�Ǳ�~��2�yze����Q��@Bv�6��j� X~��pN=S�+��e�B��m]vaa�[��{uJs�˫\�����u��p� ��E4��7�Lj�3�o�'���6�\]�S�5`흪k=Ұ.��r������ �A1�3�_�� >�o}�d^�m,*��TM�0}�<��*<o�qV�ɹO7��	�R��@���p�b v�eN���aɰ5H䣀S<_.�����`VRDu���u����,x��7�����z����J���۲���Hz��
�kH�Q�q)��Y�i�[�N
X���2X�5V����-�)�Ee�V�#�k�j�odO~�=7���s���%��언��q�Ӵ�s����Oo�Y��Y\>[]n�99��X��׃��+�g �,j�v*Ɋ��aU�6�܈��9ˡ��x�>�����vU�4wmQ)$:��'���l�/��7r��,&ܮ�I�|f��y�gX�:����ƨ���,��8h�ș�t��˶��b`�,��`5���^֋A r���T��^��ŕ2C�1��z�==�׻亚�]�l;0�.:/d87�!G�˙�<��Ց�tL,'�ս8A
j#;wY��S[�|��\���,��@�q��/�䋳��c:��t�u���-=9�@s�lu���V4�o��g�z� QTF�`�v�����2�wr��#��*��![��u`���uv��3U���zE��e�ܸY�9�yY9:���>ɻ}�JYe%M�٠�q�,�}X�ʝA#k|��듙ݤN�<*��im�S�ΪC�x�;0v�u��Z�ƾ�ɑ;)�*��Z5�2�;�lv��bC����@ɭ�caR�	����Pܰ�`�Ҟ`z������+�����-�+*v��N�8_`�Y�ի��oq�E��]r*��d�����r�(�u( �i���*m��=��y�Bc�:Vo��Ȅ�O��Z��@�-��7ܞ5�mqW���a����f��)��{
|���:!7�ժf���&N�Qۃ{u�+���fJ�*2�X<~=��3�y������WtN���t����2�=Vk�R����'h�#�2*�ԨJ�͟q��5sC���]jh�nLc���:Y&�f�D:ՋoTc�����/��6��k��h�wgCM�����w��n�.�ll[�1 �1����1.�^J�[(L�f���ܓ�`f�)ªT�����-��������݅8�t���\'7�fv'@W�,���8��u����!�,;w��O[���U�@�*��ˣ2���?��\��&+�OU����rM���zbV��E��s%jjML1���`���o�6G��9�tT�"����4"47�	�_eխ��7��腰�fM��y�S�m�-;YW_e�p�9�`si�ש�v�*����1�O2��ř�*y��������ν4�=s^$��Y����m[:k2=��8>Ipr��)�˜i�{x��NO/�&+xʺ��^q��{A W9}�cY���ժ����ܮ�Xr��k���c�����P�A	�VGĠ�,X
�DX((,a2�UE[a�jU$
Ȉ�EX�,��A����R(���f3E`��V@DX",��,X�T"�Q1��,X���I�J�Ab�j��(�
�`�Z�T`�(���H�#��X�H(������*"�0(�����0r���Me�0��*�ꅌR)��cV�"* ("�(�(.��EL`\�QB,D@Tb$b���Q�
*�E�YEQBT+"��TTT,���j��& `�V,���T�MP%@P&!X*�"�QK��I��X(
H����M[i`6ʩ�0�k���5�Ω`_lN�Z�al�y[�V)rS�\HF^�i�mPT������h��u:��l����3�K-������YD�� ����t8Y�n��T��Lr������։Z�����f�<�=ӓ��1�[���]���{���4�.����G �|�s��Z)�������i)=���*<#"��-��2�z5���}�i�wH3�9����D��\`��D#�����7���u��Xf�N�PvBmHH7!�J���,G]��2�I���h��-�����='\�������O�(���J2z\P,�`炣+c�g�DfO(R4uK�6T���F�,�e�ۢ�T��K�
�+�{��.�R�σ�Z���;j�.>��Ҍ=�����f?B��ǰz�(�<��G`Hff���<6j�U��B~�A=�T��w����Acs�:^Q��z��x��g$��=n��$?K5G`�����a>W���£�a����h���$��2%$�!� $_hJg�@=��-�W6]\x���\�Q[,�~�4|k\�P�P��w��L�U����--����(���T!=X�z��q�T1Ǌ�t�=���s�ٕ�ND��Qj���b��F��gk�p��{k�������R�����[�<J���nKt�����}�f��J��A�m����k��z���e]�l���κ즙:��B�)����5v�)��}q����˜⬘±�)�����ـ���w����ր�c�eĬگ��?`���
�[^A~�\Vb���#(2"�u����zI��Φ���,,gm�K��y�4ƈO|��s���7��C帛��홫��jc���7�>o��p�фn�wSi��4�geF�cp0c�)�ٮͻ��K��H�m��Q����c�@FzO8��M����[v�p:2�>�L��P"nl�Z$��FGY�O .�4d[�M3���!=\F.�iʒ��US�f��=�t���fC$�T>H��;��D���3{#Co{ ������GY�PW�,������+�T숵�bzF�ͧ���L��X����>�.��ź�V����wި�O)A,-��&'y���V7n�M�l�NgT��n>�#��Пv�h><�����0Ӳ�q)i-�yA-��;0"����ɰ��<���p�"��I#ވZ��x�>��a�N�Kn(@L�17oٔP�d\�G��f}��/Cj���]���p�䩠v���+ ��=�޾�FC��+������/E'���0nj��#k��.|$���0s&�3$�N�U���R��WV�P�gZbf�{E��VD	$��{Lf)���[���|��f8��S��r�X�V�-Q�'ѝ꼝���n�Y+�%`��n�Xc{%�p�K�tfE[1U�Q�н�U�T�Q=���2ȅ����u���Q\��B��wV�\�sW�e�l��:�0歓M��Rݷg��أ�t�'��49] ��U��ٜ�h��Ns�hȷr�29���8����[L�9��_N��M6���0p<z�K����n8�p5k��^�T����5����PzU ��4B}��z�%�5���\���� �(8ݍ����9�v������S0��ަ}��T�ʠP��X	́a=M�E�1�[K�E�[���Ǯ/�vg������g��<zs���e�#"���0=�y=�.�ש�U����N'�|=�ׅ����gc���܆N�ݮ�U�����sG2�a�詢�
s�ƴh�;yyThnk���P�m�S݈��=q£�Ⱬ��q�w ���W�����$���R��_�������寅�8�h
����.�f�=�����K~m�T	읢걬����љ�1�C�T�7>�ώ�j��{��:&=Р2b~��ëH���2�q���<�c:�J��z�lޱ"�U��k4?_�Ү���J�_�3.�*�(F��tNR����T��fƄ�����β�2�z�4U܄r���&��SR����O0�t�C`�qa�ǳ��o-с��&-��꺼?u*�����}`��$7��f�����ǟOWh�	��]\�4�S3c�K[_8&:B�'})��}}>ヾ1;V�抌t���PHTݓOQ\i�؎��pt3`8M�s�]s;(����\lG�v
���a��);����^|5�?!��]����x�Ԑkm\ʏm�k�S,-�x'o�sfۜ'u�YS"����hnR�j^@<�
��z��x�hS��{�$�#yt�F��p��ݡ��.��G�.�#�rb��8�6���MI�V�`���b!?W�J@��O0�q��qRPu�j}��\���V�B̀�}�X�|���%��K��U��n��*�=b||1���{Zfg�h�I�{�'��w�m��2�z>W�
�G9���=y!�3�S.�O�&��A<��@���)�ah��岑���]���e�]\�����J����ȼ�%c��NU�p��X	��O�ݷwL�CSb�B�����\���0����޶���/��h��h����'�cŋC�u)�v��?1��e�( F����]�>L���s�:[,�X�<qv3b��(<���&6^�Ƙ�\�=�إ���lX2bR�u;�e�"�ޔ�*���=J����z�V�:���L�F]`sX�32�Iռ�X�������N��K|.���G�7)�qۼj-���۹Cw8��ʌ�Wq�Ո�����nS&o����oӊ`���׮�LF����K�{g�h�㦾{�p�Y��P��u�2�������%�	�0��vܤZ{u�+���6P��ܫ\������J�G�JK�ΩL��|�yY��Ko�&��#sr�L���A�.�oL�Q]]�ۉ����:)�b�{� �MpLl����u>55=�s8���>'�wm6X	G9[R��/Űt�ˡp$u�{6m.�s������@�?�L1����$�;�>&��@\qmPyS�ͼ��ՙ�C�`���"�7m�y���c�vn�k�g���àc�}53�'�$��̶��j]Z��}�L����e�Ovr��!c�����������D�gra��4ɐ�I�`":���Dͤ{Zr/_U	p�d��%¿t�����뗾�%��?(T"	mMtI�����ܛ��p�cǻ��u��R3y�D��]�SE4v��l:�\�uc�����yes*L ���?j$�����;$X�u�������'�qZ����+R�ZC��&����]�t��0�^���ݿn��uN��W�Ab�-bs.�.-}�`�xW���U����-"�]��e,���ޝdj�vfӬ�K�����s+��*1enp���u��~�����-��uyq��l;g���� C�f/DL4u�R��F�m��(��}�RϪyl��dB�^*�[+�OECW���S�f1X�k�z+�5�R.C�g�h< ���M,��XT9�lQ� �R~>Q s��uM�p7B�a�=Ig��׺e�8Qݽ�nq�d㇣O�zє#$w�\� ��}�|���2�e�[�#��[%�`/&��L�F���y4<���Z���|�dK�d;ȋXp�md�6��<�xh�:�lw.�;�:��hh�,��z�X�h���	�h0����!���<n`k5�͝��T)�w΍C�5��p���7{��G�iM�� �`�� �4�fn�3�ر���}���lP���.T[l���]<�{���n���}ܕ6����ڦ;��=.x`�@p���N�����2fF@.�˕�;�=�����i1�9�Pj��F�:�v��O��d�P����u���.�e���U�n([����#�R��s������,zgaҫ
X�1���WǪ)&&��_U��j+IgN�[\8��qQ�.�8�{�Rd�bX��[���rюƫ}��M.�V���a��L�����+�_[�Ob�#���]D�'S��聽[�=�'!��3,k
݅0���ò.gQ�嘿���j�oԎӹ��}ѥ���s�;�h�O�JHްx,6�T^�F�n6��g���M2n�|�ϻ}�Yuux͈�M:(��[��D�9QW�*<"߮���	 �K�F�v�%��M!t�wC��v����0�˦zBgwK#.�j09��Yce������ɓ ,��ێs����G����5�+��E7t>W�A�κ��a��@��eژ�=2( ��w�����xCx[�	�|WRs~��]c�ODt1k��b)Q��F�ӧ<,/q7���)w.%@B�,S�\�!_NJƽ�7�3�s�KI�Q��xה芌�˅�ޘ�����Y�Ĺ ��8y=�S���2�,���01����>lM���3����_9;��Q����🛺f�w)w�l�?=�o!�0VD'�q.xe�K*)��$�]�ӹ����΄�#�X�*��%U<©���Bh=�jF�+I�����n>"�a�u�݁l�p��1��5q��M����	�N_[u����v	�u�4W,���7Ws1+���j[%*��	9u{Z�ax�]<�o,�jy�5��nvv�|sr�G����3��s*w&���X��v�4ռ*���v���oj�H
޽�����ŕ;8qd��\���.�X.���`zx����S\�#Z卙Z��"ވ+p�32���o$����8Y("+i���n�q�*�� � ����Z+5�5K=z���-��5����U���h.(��!�o�����z~���~8-��jʋA���0Tc�̧�k�����3�z1K�-]R�}�{�yY�/��\g�C�FKB�S�o5l��u�|��!��o�h	�g�,�KY�OB�1�X���sM݇5�S�/��,u=�sf���8���Q�Һ�˧�u������,��!�����@��~��*%X�z򩸋��M�Ͻ=��:��㇃��f�.S[`8&8�'}+�ϣ.�}㼲���k&�vd�:�%��+�7Y�HVwH���; ބ����2���mTEo���ѡ�&�x/A=�%ԙ^��P�g�e�rOH�զ9�[A��v����U
o�o�ԗ���c��%n1S哰���t��-j��ogK.���ss��(��P%&uQ�}�n�����͂���!,Y�Z�����Ҷ{��̲%?�LP����Ik��0��sЉbL�����V��v��}�\C�A/T�+�}/g%O�_7i��T�{;�M���F�-e����'cf�$;�9����0y��;"����7.�ɊuY��8X�k[TS:Ņ��c�����]���,��0wY3-<A:)�9��W(������f��n8gu�k��6op*�Ǘ
/~n1<)�r�~��Sn�k�ރ���G9�N�n���hc#*+{�M���zl����&�8:E3E1T��H�E
�R��[B���U =a��M.�CR%"c��nO����6ׄTi����q�D�'�t.UKw{�UJ��P0w)��~�yxʀ�Tk��UD�s|7G�/�M??�q�:�1�3b��D�.��5����ӊˁ����ðv�O#�;F<��w4f��K�V��O�Wђ��>��ȜU�	�nK%�؟]y����>�֮L�8�@~m9(�g���۲K�vy^6�<��̯qez/�f���8ԇg�����w���R����j/��7*�4ܲ���X������������0I���i�K���{� �,'<2�Z�]]�۶;���l�c��:� ߲��C?�n��v�茩�W�=Z�o���zg딲ˈ=�f OM<�6.��~�-����Ѧ��nOz��=���%�l�s�`�wsFþ�Bw��=��LC���/��#�Ǻ���bF��g�ZW�;�m�33s%��Ҙ%��nF�Gi�*´5U��w5��Ϯ��];'-�t}�v�sj�p'D��]A�z�3�(�o�C]��]3Tm�xv�lL��c6vS�ң����l��êX�V( ��3��31\���Jۃ�$\W`>���Y;17�l�Ez�ٽ��sCl1T��N�}3�D��*=����~���/v���NL�Í�nƚ������z������<mm���KpN�6`��莥c��k�Ј�"*�؋��_6f�<�z;��mݒ\.�o�]J�ހ~����eDڑ]}ӎ�;��Ǒ��M�}8Fg<2นh�2���,��[�㻪�
�T� �T�����������i��������pe���` +�<��.5\/�:-�p�]�{��  ε�������͏ڍ��V���̏?��(?�Fp��	�zm��^�]Nhl'#mg	��=�ȗ�������z �T��.s�q㰤c�*$v�>��i/)�GQ3��U�/\�٪\lP~ɣ�.�w����Օ#�B�1I�����3@R�2���&���k��C�����'��#���:�=�v�����x�脆�T2�e�Xi��Rsq�.DE^�_T�Ї1���wֳj��tb_*a�{oj^�ǜzcp0eD'� �f
Q�)���n���$uOc��q��nE�1�w줊[g" ��6J����uϝEv��#��=4���*�i��N��4|���y}S7;�����ʾ��ziZdr�%�/z��k>"A�2�Rd��Q���p��Z�\��{tX�"����v�w't,��"N��=����.6�nqn�A�)+�D8$G�d|f�-s�\.�i�l�B�?sQ��8Ы��͞7�a�A�a����Su7�6`Z(���Z�O7���A��w,&�JPܘ��}���0Ո�<f�4���>t����CK���]�nyf�lg5p�\5T�E�b#��{V
:h­C ��#���yy��os9-[ ;Y*AM1&>����L "��f���p�k���w\o݈A��U�zg(�����W`���:�iY �k�-wZ��׊� �����r���"Y�NȓI����-�[������G�9�K��
A%��m�&��|���#��ͻ��Y �j��j����ͱ��sj9k��]����2���Bni���q�Xx��U�T��bm��We�W���Gm�s�t_Z���6S�5h��G]���C�$Bb�+���:�|fst�BLf��m�A-�3q��ԭ�a�,0���w��E��bf��-��&�Ŗ��Q�>��	�ۺz�9���䇪���#�����.a�I�v*��}�0#��N*����*-8i;��zz�X�&$ �6T��+FuΡ�)^*y�@��2���6�tݾ����s�M�	�@��n���o0���]��5�aTw�j9��m���r����=f���K'G|����<j!��"��i�b)Z�Ce����^}�T���$���M|Z�h���ԓ����s������o,a��S�5[�]��;�	B�*��nb�&�m5�����;ov�C��d�t�Eqt��\�ō�ʻ�r7}Ɲ�o��v�ǝ;â�t1;���k9]g+:h83����ٮ��\��d�k{�3��c�
�����墊�$�Uv�TmV* �N���TTN=M=�Ը�HQ��EXK��V��}���Gid[�p��,4(�R9x�B�4�&�V�;�m]e<'0ǚh���p?��"���)�*̏�<,�{+��f�z�u��=oB��)GV(���F�Y������,j�n���l�{�]D]�K��.�j���n>���+t
�2�r�Vn7N���6��Y�qG����̺��� �.p���[��^L�)���C����w�#G�5��#���Z��멛y���ްxUB��`=��V�PG�1}�)ښ�i��!T| �T��a-�;���$PU+
�X,4�UE"��U��BH*��2E*9d�)q���*#� �B�QC��F)J1`((m��m%+ŊAIT*��U"���L��\J�a,�dƱYb�PF����Z,m��������"�("�eQ"*� �D���aP*@Y2��֕��
b@RL`VIi��+��,���U�#"����� �XVIQ`(Jʘ²�f!RP��
�AI`���T�mjB�e���"��2�DIUaRJ�aR�F[I�+$D̕��R(��*R�X�P���J�����˽��=�l:�+�� �+��̋�iY�V�0�[Yd�WB�6�̊s���ќ:�Pa:���{��hD�v-���1;�q�����z��5�5�9�8S6���c�\_)�	�]LP����geF���J�Y��#�ss;�B��#x��)�gO�F/`�Q�\�����b���7d�эJ7GD�d���o9�92MU9��CKI�˘�P�V,EGE��i��Q�׮#Da�E����b�5����ජ<Y�"�#�o<�$gwe�֩���G5m�Z b�S�4Ƒ�U����T˻\��1�ᮻw2�tN���1�ͰUc��81t,^ssś��m�้KI�P�ķ<�ӭ�+8c=nʓg����'y�i��{����HSg4';}�{��������:Q k�Q�ZǴ�љ�=��J�]��]o�GYf[L�L�k4.�E���C�ž�R�u�!M>�8:[2���1~�0g���v�=��f�d�N+gNlV��¯���h�6�`�K� �������Kj��x;�)�
h��hb�ңxc���/�B|+�>���]9��ל.�ݻ����L����b:[���l%��@ D^EK-�\����(�ݲ%>4�������9	� 颀}/iyT��1��ny,}�WM���޹H�}��6Ne'���������A��)��ǹ� p/���x�V6��\��VT�5�ߞ 3.�Kp<��;V��X�W�\����Ҩ!�.@�ł��bج4�S�f�?��,B��*��.�{>\V�d���g@���!c�S�����!Ö=�K���0L2ܹ�o�`��I�M�T#w����[@�&'�EWy�����y��31»���
꟝�<�� ����{�oo%����y���m�#'E6��"k)�
�Wu�|�al�����m�B�f�.�82ʙ3�7mќ�*B��::5�N?S\d�V~؊h�@���{ʵr^ԭ[���*��C��mP��1-e:���4d��k��lsŌlP�Ѹ�o���}8F�\^:[am���/��tء��Φ�W1��u��U�'k�L�v�8.#<�F9'���}�}�n�Q��Zckz���ġ���u8{�o�����ʄ'im	����f�=��vq�r)^��c��^2�g5�5N�y�KE�����ϴ��H��eç؂���|7�N�n��<dc�9�{W�Ւ��i�gP[ˁS�L��eW`�=(�l��.	�}1rH;�ó&�S���c3�D�J�/��"��L�낂�,�x �2ܼGJB����텢�����.jS�a�uL[8�����X�|��Zw��3����9�e�	w^ ��8�TΌ6�X���(<}:83x9�V��K���ٍu����h�g�H��˰��~C����u�W^3'g:�x{�F�k��������;e�x�o ��|ܾo��Ǖ��T�I���j��ތW�D���:��8d	�8�Tۆ���H5�l��2��)�'��U�֊-5��]A�N=�� �K*L� �6��U|�<fe���$��gI�H�1�a?19(8��u���#!ܸ��
|�� w���hi[=��Fex0��Ƴ(�����gM'/���q�n�s��L�W
Ҫ!��"	z��`,hu��*��U�
��"��G6��	n�Esν.3\,s�}��$�{�i�ߦ9*���P+M����`z7}u3�/nr��{�zEEO-�̉���pE%2�L�ݔ M}`��<8͊2��p��-s���景'���'�	�DI�O��]����3}�s�V��4�Ɂ;Ukͬ۶��A����r,W�|��eFO?�2�P���������n~�X���]u��U���51��d��l
���	��ew�=X�;�?m�y�9<��V���
�c��V�˲Q �c�mΙ<�=Ee���t@t�뜐��%�����?�<Jkbhá=��n���y��1v7�V�N�
�5�r��h�7�۹#%�u�Vq�s7,F�����t��-6f/�q��gi����)Vk�����&ƻ��8�Գ_�!W������D\Dk[��wd���[�#�&]��ޮ�ی�x
�Dvk7*�5Ҳ���u䗯]���B{:z7&���9ޣ�`�E����q�B.<y�m�T�euv���w+��E1�U�|rA^.`Ӝ��D����5�s�S�t���K�V�eWTs��\������R�θf�p�T�r˷Nʹ�[=�SĚ�3�:=>��� 7ѿ ����ʵ��1eL?Sr�/��#���9x��S����b�"Z���c�(���g70�m��!�;�ƙ�� @��x,����B6룆���%!$�����U'�煫^�b�������/�����L��OA�[�-�z)����e>�j��"�)m3�D�z��H���.�����WR�z���V��m4C�@#}�����w�՛���;_��V,#0�7p+�����\�5�>�׮��͕6�eI�]�a�{�<��q��A�� &v~�(���-�p�Xj�5�ٞ¸tf�r�|+2��}@v7f�N�0/���#�C"2�<�W�MA�8�8m��(s�C9Ǣ`K��^mn���7sef	��z�7w\Z�wp)\��(��<
�X|���I5���ZkP�)VL4i^��y��u6=�HU�q�n��wJI��x]�r�v���=29�:j�3��q�t�1"o�c��[�[�
��ړ�����M�V:n�m �4��z�d�����,-n��S�>(��"���H ��ƴ#k�R��\�c�`Z�7%?k�m�G
�o�3o�^��5�K��t=�ۍy4}`r�3�:�OVP�;�.sw��\��=�W%�p���_���ͭ$�w��9�f��=�T���X�^ށ��Q��¾�h��.zc�*71��P����~C#[r���U���`wC��Ǳ���On5��شk#���쀆�T\��F���;�Ej�}�;��W������9Q��Ɣ��R2%�{���=�(����Z����,����M��^�K�1]\�ٴ�';�,�0]��m�v!�j����� �}K�&���2ɁQ�L���s�<]��T��ŶƟ=�ʅսKdf�����(���TѦ�]��4A�1^�N�1�p�
z	�]�ѻ4@��|a+Om�ʱ���f�W9�O27�T��P\Ā�����(�U̼���O
�j� �HF�Y�,-K����$��������]\��nal�҃��iM���Z�D�vR�/��M/j�#�6'��2���K�]�����Ӭ�����|��g���6=Bܶ��x��I���si���9�[6��"wu�ת�1@���v��֩l���t%���S�w���z�)�u���8�e�����A���	�	Ȓy�+��[L�D�E4j�HctF�g0��}�vʷ2��'��՞���k#�s���t8��	����U�T�;ep,:/@ 5�k��%cWZ�W�kڝ�����ԇ5�4��h`ǳ�$iQ�1��'F��,WQ~G"3�]'Ë�+��t���\���1���U=@�	��T�ڹ�%��>eU��GV��ct����ݚ��Mp�R��m
-ߩ��8yc�$����2����e�7!SD��ݸhD����hSM������ܦ`�n�~/�Ƛ�^R4�\��ܞ�0�^+�����9��'">/<>Y��W�'�W�-+%��Wu�|�a/z��O�����\�q�d��z'f��7�B�~�0'��8�Mq��X��[�|������4
n0���c�;�5�9h��s�;3(`�&��q�C5���\x�*�碷!��;]���W�9lW_��+�����{u���܋��=��'�j:�f*��72����=z�3�4b�|[5:1t<�Tc�vo	B>z�_U�ޛ]��BFz�m����{�vӷmG���i�:m[d5x�t)�T#�*�kO;ɛ���hp�=�9E�qr9���q���.��li�(��bf�Y5k�NR^m𮨇2Y��+�;�s7Fw�̛�R뽻% �k�x�B�;���f�ʂ��	�
��i�\&�?=z�[u�\���~�u��L�J��
C]�+v����ϴ��=��I�"9L&{��{�c���������k�1ܦ��,���e���X�΄�9�}p����z1����R�*#�;��>�U�x�؃�lO�x�ҦX��P�\i���	}�tZ��
8�3[�s&�[f.�x5���d�����'z=0Zp�*���1�=4���?KhVA=~���>�׹�^_@��t�;�b����; ��ҙ ��u=*R<�
�[<�l���OA����i��W}o<Ф���A
+�M}t��\����Y� w������bI��1jJ`�Ӓ�fg����:滥 ^٣��r\n��uW�lU�E�ڈwZ#��q��ySѳ�F�S��<�dS6��݂�
��yMp��]�W��w2�ރ�.���F�l0�{�6-���u�k�S󚼐�4g c�����T�5�=QB����
꛺.���DЁꌏ�E�5ل��a�e-���d֎��k�)#Qѽ[�Z����?�e�nH�r�ɨ�n���W*T
y��u�tov�Y���5�i
|�Ŷ��܏i�v��wǓD�o_P:Fe�a�}w\���0��ݥQ���
��O,(�ڪ*���и�(��,ꈯ�3���z�n�}����b����Th����(f��O{����X����������|�'.��̾��[]��)�Fd'�\��L��9H"}�4g޹V������n2C��ڙ�Qaa|'ff(�ˮn�9�P~w;�a���خ�[�
���7辽��ǯx�X�s,�f��0��)��th���,S�v���R�m���m���*�-ln�sM�辽�`���p����-w�au���nGk����7�L��3��㜡{*��ب��Gp9�-�I]����t�2w��¾bci��9�x����S�V�2�\AQ�l��p�=4�m��`\�G�Y�*�N~�J���$��+���i�k�G*8����8̧x���3 �B�[�{�Q~핻>*�sN�G]
~�Q+�=����Q�h;��r�-�w�=
�I��Y�'sb�N�3i�hɇ�Y�v���]�ͭxzf��I�y����l����J]��E����Bg� w�{޺��xEi�N�|�~K�����Ce�TV�ek�,W#�{��#�2��._u�N��Y-����컹1O���"������΢�D�>�߀�F,�Y%p����b���!B��Ĩ)p�磑�v����9�b�d��uf#�p��.����N��8r��?��n�U�+�E���$_vIp��z��鯫��8K&w�
�n_j{��R�)���{h֨�W��^��I��.ե�w@j��
=-����p{����_]*m �8U���a�L��A~�Ӭ�!�Tng\.�XM�s��3�C�GX�I�Y�;��7���H�En#)��>�@u ؇-�3���(�zl2��1�|"S픆u�K�;����|`p��uR �= �@�6�*Y��`u�ǎ1�f:w� �u��/�k۳Ix�{�.ŏ8+bG��>�w����7?nH�P9�1�5j�\�2u\�utw��g��ŅG�]x�#��s�)�F����yz�8�ͽE�B#�а�'�v���&؆ن�kɜ��m�N�-f�p���}��G�b|����Hsc����M�A��+X�b�i\ϗl�b�Zѩ������=�W�SSت�	���&�F�I���*8W��>`�GE�ڙ/���S\Ft5F)r��zi����tw���f��<K?k���T�.�5�ނ���WV����YB�n����k�,+%b�(��k����.�#�a��;�aT��
M����.�͙pʱ�xM�E�b�9m�K9���`��v{�A�E�t+;}%��wXtq����a�]pu�t��-�y՝�����5��Sf�>�"�b�$T(���o��1t[NT�Xs4�=���`j���y9F?wG!��+Ex�l�weG8��8�2��i�{֊�^^]��5u����68@�f̪n7�<G>�Sn{^�����<Yދ.��b��-'|r5Ib�H�Л�{�L0�ut�Ui�췴��۳�t���/��]��uus���;a�s��sC$����,e>\p�&%�).)���ki�H�h�]D��#P�׌}��΁U�1�[�5�{��]n	𽝅�(�<�.k�L��"�':3=��Mq4�
5�W3E�tj���%Nl���@��*���T��uL��~����41�f� D���à��"�Q�B[h�7m��Z6�j�Χ��4���DGE���u�	es��,��l��9!iX��U@���$ɡ/{�'�ooM�K�xS�Oǣ����:�	��Gj*Ym�]��W9��k7j�6����[�Ӫy�����zf�3W����uO�a[�y������1��	�xx�h��D�جF��
�����KR����-#.���D^�a`O*��6`�T9 ���FFn$ف8�쵍��4�	�/cwb�o+��\F�CWwVR��ES���1�xj|��
�U���4f^9���`n�����Xk2%�\Fu����M`x��-*jcd5�� �f��Z��vo�ڄ��mv�v�������������<4m�m2��b�ō]W+k����@�����j�hu��j����>�(�zk�İ�}�h7�}x�&Y�#>�*8H�
��l>�����wԯ��!�YbY�\]��ϊ�:�� 3m!6����u2r�pf��ɋy.�Ʋ�v�����0bf�YiMŌ�(Ⱥۻ�F�s|�掅kk���`�AJ��Q�(o<b�tz֍S-�OYf��+-�fGc����>�e�B���j�� 9���Kl���L:�ӷaҚ׬V4���s'P�/�f��a󝷮�>m��e=Z���	^^��Kxҵ���v2\M��[9��z�����W#���	}����H]>� n�_4��i��6�ɀVL��j)��]7v��&��ɦ
������U{�fVd�LP��V̾\�pU%id�lpz��ZBq���t`������rP3Vƥa��+4T/6A��m�yi�]��
9�g%��M����h��F�W.�Y���rۻv�nx��e�r�:�Ѻ�껨�9d.�m��'&q��*��at��Y�z�XyB��J�	���wU�[$�Y�e�/�vv�P���Ш�����/twu[�"ՁK<m1}]t��D����5m"�Wa-Mb�n���P�7a�r�t����P���}{�|�,ΐ-��ӷY�;��;�rn����J���>ahY<p��@8�+2&;)F�˻k�����ؼ|Uu�z�{���i(u+椆n^�6��d�(@�!!ט�)Ia�.�v˷[nR	c��u��t!K7�>�6g��8,e�4�b�N�R-��u0N|�@殾)���}|3�Vr��j�Y�`�,����e`ѓ"ھ�ō�\㝐%YE��.�'1����V����5+2ޡ�-�%n=�K�e0�+=g�Rzr�͵VN��t�KD����8��}e�b&�c��X�$Y��؍���}��L{n��8t�4�}+gQZ5kc��!P-�;Iw=7�J(�B�@��aI��؛	�z9�n�56�V�s�s9h�M!���*��c3�gQY��ѽh�W���!�}.|�/��'U��lI{h���x�=qN�mvu��wW3��f=������E:� �:,������}*=I�N�W�%ܳ���Kf�cu�PgL��QYd��@v�wa8t��ūZ�de<�8z��',��!�� pm
��ڨ�˲%�s��+��yZN4ƫ{�k��!ΎAO�v�)�tD+��.S8V�\�3�ͭ�|�A�͹���6�z./DE���ң�AcJ�\�q��Nn�a��ϖ��bvͭ���z�{S�VVjyJt>�{����䶱�
J�C*E�&3Z⹙���!�V��IX")%nXV����eL���(��e�ZZ�aR
��*[@˘1��E-�+K��ʸ¡�+"��kb��T�J�T
���1�&%DTU�b!mX8Xfť�A`V�J�3�+V��YY+R��
����IX(�b�Vc���HQPY���eH��1�0�# �-�I����jF�VXJ�"�%J[+r�,Q`�q+r�,P�*�bŪ!U�
�%��B�X�k�KE��A�E�LʉU�V�
��Z �j�4�Yb$�Ѷ�Pm���\Ic-��*e�j � ���YJ��ԕ���QK���m+1�10W��5+XU���Qq&e�cP���DZQB�J�m�a�u�޵��g�D���9�:�e�K�[}]��G�p*OUÌ�����۹�)�Nܝ`E�x�ٮ��ej�"ހ�J��G7b�\�շ��{�a��7�'����f�ip�K2����1����4�e�Rv��Ӎ'8�G���~������M�n��;�	�b+r����n�Ө)�V��!��r�d�#/շ����&�W{M�E��2-�t�h�Ot����<���ې����<�T�V^��MAT�9V�\g�N�ZL��,����o�:��Ze=،	�#8q9ʹ��T�收.��퐄��wv��{�{������u�|ι�n�	���2ˆ�ˊ_���d����p�l	ÿ}���m�!��R�}�x��Wu;�����๯5���Y�� ��m�$S�mQwZ�1�-n��Ƙ�<e�L�(�-͝
�gBA��}zfSf��B[@ޫ��g�m�����c��'})�Ku��tM<I.V�lzR��~DU,���f�V&̓�HqЇXn^��'���#����)���|�^9'�
}Za��:m�_���"#�����o��tg/{ab�K��\�S6�mm@�܁Rd;����'�v��Q��zz�5���qp:p���Ru<���/}����g�|e��L���ƶK�D���q��H��W/���q������s�b}x�y�m7G[b����)Aw��ڸHj�`�e=�����\��zW,�Zn�������o�^	�{ɗ�N+�d"��� p;jGQO�W� �T�[�@�S�v�c���Sa�0]�p��K� ^�8�p~�.	�uc���>W=\[D"713�_B]�� �c�ls�h�6��CN�����^Xҹ�^�q��c�S�a��[�� 6G/���晻�C󧟍��+�EA�g��C��9�- ��KO,���E
�R��Z�R��9�̡�����PLKy��.RR<�ОZ��B*��������AП��]�wep�U�qu����UuE�f��[�vݏQv)� �[@�2�<�X��q�8+أ�f�MuQ�ٓW/͵J�;��d��i8�q��G�ۚ2�r��Yk�'�*2C�>�ʗ�����[j�'�h�P�%��ە���oЍ����.�a��2h=�8h��`�@V8�?p;�p�֜j�%�ӿ0C��K*�;B�:]�^����z��hft�5:�����u.���fgf���IBƁoAD>:�T�W���ʪl+��.��q���Fw�����t���+z��7������<�d켤�x����J0�=j�>O�f]��h��=3WG��L���� �pN�ԁ��2�gU���$��s��'>�uA���R���]�e;r�'�e������l��V�6��5�j��u'Mt֚��k&]��{e�Ŝ&������x2#���i����e�Ts�l��Q�4��®��Bg�E�3x�7�[Ez	��f]�<D�[�l��&Y0&7�
�8��,���l��6O��g9i�8E������x9�V�ڨ9�P�������H�w�^��wt��޷5̿t��չQF���޸u^��/�}�S�gK�����u�[s��%�ΐ��U�& ����8N��fM�H�[,
���I"��K�m���5Ԫ�t�S,�aѦ�\���O;���6ϊ�iV�+bL�;*Ű��b%�
b���/�&�G!�w�VX]�xF���H��H{�����"|+g!�K�Z�x�Et��qe��f!`K�5��Ӷm<s�c���;��7�.��ȍ�ލ�wT��*��ШD��;��E�Gb�#O���	��\+�-�b��!%����(�n��,뮠
d8b��5,�5�c�������b�V�h���_K��ͮsK����TԹK��W����g|u���e��v��J��JY&.5䪸�Q�t�SGu]9v�㕉���wz�!��W$u�������|��m<�QV��t���Mڥe�>�Yd��#vEa#`	\�X&oss8�;y�7���T��������cjkY��MY�rvLL2��켌*]M���v���;ܳp;�;�7'E{c�\Md�ǉ��{Ff8��*���0s�,��+�Kӵ8\t��ǣ��.�E����b��l�S^L�`��I��ͪ�/�ш|����ٗ��yem����s�)��e��'�0zC=	r��\q��	�:)�T�������z�ѽ�v3�ۓ��^k���6���^�1�:-���~���
�Ά�F)r�c�^��])QINm��)36S\
�5Q��6R��7E{�6��EX�	�Qn6�e;Ǫ7�{@�A	��z�X����7t�x�ǽ��uٱ<��7tv�����h�d���4A���N�_#���iy�j�:M�:�PA�j�S.�(�#��9V=�k�Ѷ�y����{1n�m�.c�ԟv����yO�1>��&u@�ӦH�
�.�n�C�!y���N6�><�WW<{&rt�D,�v�g���h�p�Xw�y�JK�̔Gn6�iH�h�]D�n�r5	�i�R9a�͕�;��v�)q��uA��˔�[ء2�WL�N=��{���B���j��~x=��\7�0	6�ڑԢT�xа]�z��Գ���G��V����b≇��=s}Q��X��]�[FBr�¹uw=Wz`{;([E{�Fs*�wL+"p�˶mN��|3lӤ{��O\qt)ej�����ovf�C��@��e�ۃ �.;��� ���v9�Ő���ו6�eH [@Dm@�ޑS�@���^�œ
n'�	��Ί��쭈�/ۣ���4�=L:�"���w]��+��@�h��=s�0ںs�	�w�F�w�D��29�B}�����9�%��?MyZ���������	.+�FL�\��Q7�B��Y&Z��#y�w������	l����s�Օo\���1�;�PWT���m�8��1��:�P�6�R��D[�P�u�2[��{E6��Ed���T��r���oS>�&��m2��S��6�[A�k�3�ȱM�9����Ot��#F`O�[����w;�$?K�e�Ww�xf�j�B;7e��ȱ�p�����W�%=���5�y�X��v5��ɪ�Y:��ɩ���t\*���i8�_N�E������jE]���u̳r.''���#B�%��Gb,��H���=R�L�{�zkZ��;Ju�7vQ~�2i�x$W�+[%�5���'9��74��1o�qz-�*X�ؕA��R�m���n0�O�ӛ�8l{�g�.�#ӛ ^3�o������
b�T��Ge�4����I·u�yl�o�S��>�(wU�'F�鎊�#8��z��v�3�F�~^X�K��r��fF4��:�u؇:��jm��[�6L������tӻy�+����n�;��}�`s�>��謚J�3F�tx�G��g�*$x�ސ����-�e�ʮVձ��9�.���Ǩ��v�N�tngG	3���(ō��F�(Jdķ^*���ȓ���=|:R��R�]?]Y��f$�K\�>�Gf�h�)��{`na��Ѱ連z���B W�����O�[t�	���18�㼹+��0֡���4�_[vy���� ����+�L��]kD��/�����;k9���B͍s޾T�+�ӭq��y8�=���밋�q#�z����[}^t߳�F(273^Kr���ne�VVF3��7�I#��8�p��L���d��PFO���.��p{=�x�OI��O� �r���%����-������yץ�k��r�~�`�����|0NSnJʚ�n�7-�?m�
h��(E?>��3]9[��)�DZ���zb@�Zw��h�|����|C��.�c3��L�9#Z*���㪸�9	E���×�,��h��C߭�=�?`4��e�De�#weSs*�C��a@�2�2y����~�\c����`{K�b��O�qM;�l����,���w˃l.�o���������v��N�%t�]�u��hԐ��{hl1�ۮ�>�,���[=�AÕ�s`�P�1=g+Y��[4Um[}4 ��wPs��-	|.�1�{�b�Z�ӯ��`b�8�l��y������k�n2��m���e,B��7/������<u�
��WjmY~���Ȝ͆�)�"�m����X�N��\���Y�*�,��
7m�D�Ⱥ<�e�i��뜖U�3�+ъ]�^����z������u�M��ɢc'�#VNQ~v��(��]�k(�mlAe��Pt3&c��c��M���-�uv��lw�/&3a��}7;�UWrbxp>׆�mi��vJ �C�3��؄�m[���*9�ڕ��M?Q�l��������������]m�(3�$��^"j7��O�a�z��&V��`��ڗ>s8v�U��x�����:h�g�)���wA��
���t���b����>��kn<p�ٝ��BX$#x,����V�=�I�����������E2���e�^�K\:X��&"�7�Xw�:�KJդ)�JB���]���uA�r�0]zi,�������6�!߸KQ�yg�X���ˁ\�4P��k�:W:y�#-F�5��f�R��Hc�g�AУ���'�Kx��;2���D�����nPyO�'���^,�;�T�m�~t�9��#��T�])��Dъ
�)����sX�w.�乗A�x��of�"	΢�p;�E�f�\��Y1]C�Ⱦ��oۗH�w3�Ю#ǵP���t�J�����@V-.ym�1�������Z��}��0p1hD!��.� +Ȍ�EJ}����y��[y�.ꇾp���7�u`�ݧ��Jz*�ܥ��~e0 <:�>��m4T�5s��vB��t�Z��}6�P��;^ ,1�#��_������S���j���h� �QG|
�W	�ŷ�0Pw|SA(x���su�,�8��N�>bo���L�0-��}���8����m^�6��m��( 
.P泲��"�{�^a�I��ڮ�YSw+h�u�zWU�MR��vYĦr,=V��������Z�q�~� �	�:5|9��T�si�i�f����m����n>��������i���a��l��^7� B�lA~7�W�#:��ʇ�X_V:7���Q;��>��=�te"yv+n5 �C@$)���w�����i�4W��5��E���7��:MO:��G�#�Ƕ���7�{E)�M��*81�h�R!{�C��6�<h�c��Y�w
����
Y]�be�q}/�>�FtCl�h3ss9�ԣyRp�9��k�It˪6�J��b�u�����*�̺���3�Ђ]u��+8f�;}��x���8�������-7.`�e4����	���sOk;��Ҹ�Ή�j��/�n�5�w��0�-���a�S(�О�auc��F�oO>�A����]�|{�Ίx�+�T4���G\����s��D�x�R@���[L���M����	�{d=�̦�x����a��t���V���y� ��p��@�t���^BR\XDu�-VЅY2�P���o!����Z֛{�h�Ьs�u�����~��'_Kn*e��&Bq�W`��������7H������[��-\��GF�,t^�B�,*��̩h����*7�>�������ѽ��W�4�o�����@����)��U05@怈�h�e�\��؛jj��ҳQ�@733�+~"9�-��~��b�E��?U>=�K���;s����7n��,�5�`cMfv��4��>�O<��F�P�P�Ƽ�~{m�B���j��v�.>G�VM]Diܥy������j�ZkVS.��۔� F��£���Kʷ.����^�����j���t"�T#!��E�5;1?-�Cr+�	��ǫ��v��H�{!h��t�nҎhAa��-g@��/����t{�5�+�WՕ����v��&����
����g���<�IT��XAǶ�ر�����7�
�WU����ғp;�ܚ�=�r�������͜�n=��N10�1ǣ��,�^l��ٛ��5c��Z%�(�p\m\3Z.gUǌ�J�z,��]���"M@�ݎb�K,��֧8k�������A�R�+��b�!;^�f݇CR�m eML�A��9`��%��)���^��}[�:nΞѸԧ_k�ݖ_s�t����GC,�/�^2�1Żt;q-����h\Fyz�����]!���ќU�ϴf�=6�q�t*(�G^�q���2z$B��!�N���p\�Rˁ�4�m���^t$	g�Vk�����,gs"S,���o(������c��N�*S&%��Uq�:y4c�	K��NJӭ��w��'�>�7�W�V�b���R�x�ۘ��(�ԅ�N���K�P����K���B��驕{��T�pz�^mk�y���~�c:�h���t��Й ����Ji����O���I|ו9h��<�f�:�2^6
��>yvJ21���ΩQM��>/3I��yڄ�@��-ѣ5ߛwb�e�2p[ ��/��$k�(�Lk��J�ty�<+�@�$��H�ā$I?��!$�$�	'��$I?�	 BI�0$�	'��$I?���!$��@����IO�BH�r�!$�$�	'��!$��$�	'�� ��H@�����$�؄�!$�p$�	'�@����PVI��E6U� >�7��@���y�d���1/��*�J�IJ�T�*�"H�o��R6b��Fڵ�P�j+mSM�)R���Ot�l��fP�����T������R0�*)N6��!�+jMh[5��V[@�Ԕ�%���@�{� ��V��R����� �:;bk(�4ڵ
�4hєQT5[SpnL���Yj�M�[u7imn��'s�jmJ��[l��[AwqvV�kl;��K��mW]��妷[����Vݺ�k�����wJѹ��b�6�cZ���a�ݪkY��nrNr%�d@��.m��՚D�M����EAa� ��+R��`���UAF6"Sm���K�wi���j���QU+T-��+4�R�[�	ӚV)
T��%��J
�����h  ����!��  ���x�%*�       `20110�L�L���T�F�i���4d����h�QF C#)�L�=56����3&�ڐJzH�Jz���z�0 ɦ=�����i~�:��&���P>P�9� o?H� �+�T@�}@@��9���c�?ԟ�C�!� �6A �`1� � �B4H��	XQ@���9Z�X�����@&G4&�,�4q�����^Yd��xt�H��L4����z֦�Li8^�lky���1<��
	rΐ��C{�3iӏt�P[s�RM7Nf�;��Դ�b[��zQ���4���$�7rK(�l[W�Qot�2a�wR
�"e5��ԓ0<*�Kf��&�<i����D��F�.��uz)���D�Vܓv�7{��'3M���Z�
Ԯ&�so �	G�JV��
������j�y, !l�V`$�1aAK��F7s
���ɍ@���5�%3l�ݘ��b�.�2P�j�;��c�]��n���:�ߥ��'N�J�D�3&�S����r���ɚe�⹋��G{��(�+Y�Yp��C5%����t
׺��F��hw��{I��%��OZ���xU
:���0�W��[N�B�b@Q� Sj��/*�Yu��[J,Y7��⫂�4�EL/b���;��������Ko4+�)@i�Њڗ1Mخ"E�(�Kw�c�NUM�oF�U{���n�b�kt]���5؆��J����Que1y$�w���{H�H��AX�w�+���[Z�1����d�j�B��`Z��FYa��R*�3hR����9�$�ܕ*k:��V�w��Y�X5Ѷn�I6�J���bU��YT�#�P'�dAGKi�q�4m��[,S�m^YR�r�$IS�XiGXQ{x5��X�6���*4�
�����N�ͼ�t��/��3��
r�E�1�*����mDfm]^ꥒi.%2��J�M�6�sc��d8V`�Kũ'�n��r�ݣ=�pN�U7h�]A �Z�ԝ�YR�M�n�f%� j{t��M,�n�W@�W��c��A�[���[M��Ј]�3�F�H�Y��XEd���l�#)K���ܺ��Զ�L� �O4m-��m��(b6q���kl��]8N��k0eIbYK-�W�V�,�7��LIn�dkԃoA��T�m7Wzj9"��t$��C�u.��Q�s*`��Gzm� y1�Y��^�%፡Cv��D�K-԰4�I��
�n�۵
�˦]c��ˑ�C�k!%�
��2� 1 ���eVBܳ�sN�7�����r|�	ں���M����B�9)�զ1�۠�Օn|��7AXU�ȋ���S���I*)�  ����H�M˷� /40�¥[��kl�ܽh�����]W4�E���&�Ұ�������4лZ-ðR�BD��7�k�"	oh�c�;R� �0w�2ζq@�RzU\� C`�7F-�M,�"+Pt�ұ��$�K�<��V�q��	f�vQ
i-�df�'r��ӄH㗑�{����R*X����4����-��њ��S0\E����kT�I�I��3)�ݡ�h��)b�B�M����ۄ6ov�n����ة�/�5Xi�ʌ�Su��H�.�������U�lh��J�)�A.��rݔ�;X ��"j=���A�e�X1T
ҫ[��P
%�%�T�8��:�K���Q�Ihң�����c33s�J��!����b�]LڴbN��u
�����n�t]im��Z��DA8`zb��Uc
VX7�У�ih�R�������
]6����<�hͧ�e3Q��{Q����k,#�X�x(,�&LIZB�wsb�+R���U�Ҹ�5��p���nc۔��u�qX�m	�Z�3@0̬�w(R�R�[$��&��1$iZ"�ө�kAd*嫭�y-4��^��Th[�C�V]���4\�T��qصz^S���JێH�M�<xÊ��B��u:�6@D@QOn�ڼ7b�B���v������Ŵ�h�h��R���&ea��3r�[�� ��o-+3n��c��@�p=*�Q-0��aR����÷a�M���D��+*f؅��� ���*�4efh�ei6۶�8T�'F�F���dB�+0�zA�y]�����i��ޝWj�n�e\��nF�r;X�F��)��XaOKR�]��c)���2@�kVn�tD�	���t(��ZuO�cq�V�2�RE
��^�h���F裠��5�f��Jtӹ��U�6SAK7��]G���@b��D�Ht�ܱ��͚CE�(M�Z���Ej���X�jܕu,�YVF:�5%��-e�Wf��j�{��6$���O��-�UwfV6��/`�GPc�lbD��NНɫpgw	�f���{�0L�+m ��Z��RԦ6�^4�r����4�^�c�/�0��',�z��q�U8��^�R�H~O�2Y��_�����Ί����u��§�LI���m뀘�Iq�2�㸎Xr�x�8R�;{�0���݄@)��Y�MH(�l�]�W_]��}3f�
��w�^D2
̺0h���2{]��.�r�ԓD�vغr���P��su4ѭJ�����ѩ�k�A/���� Uk��*-�[[��:n�U\�̈́k��h���1V����sjԪ�2 	��p�"���[U��U�e�9Y��7�71X�Ks��֫H��`{�|@7G��A]��(�݄��4,L��g���R�]��:�迹�,6�%r��d.��6%�g�㷠M}˲�����c=�k;�v��v�x�UטO>�q}�Y� �Y��D�����%mu��D�?�nƘ����$��%���ȯb���넓X��x�4h��*�RtĆ�z6^N�;��JR��bWX�훊؅���ok���#E�d]�c�X5.���'��f�˖�\�u��̜�i�7���i��Y!QT�!��7��j3)��6q�D}�n�edS�Ԯ�f�xV2��&@'��ﱘ*O��]��K��L=o�<7X�j��r]�¡���#9���L.��ѣ������]�GR��v�jE�T&e</0F�B�� �r���bbQ3��}wu+.�'j�#��u�Z�6P�\{2���U��b�7T6�W�����JTX����#@�C^��ژ��}F����;7*��� �����zf�V%��h�H���r�f#�J��Co���]E�1Ɓ����g��a�>�a�
���E^X����R��{g+
�>������{\%#V��7���C�V��U���@�w6�;k�k�雖�k����賻|���c,�7���3+�+��̳����G|����N� Yo��6���"�,뛕.�\��56�`���)���c{�����e�� #\�wz�,�[.^C�iL�gV7������	�K��u�K�yV�'	�*�	_+���5m�h�������1R�!�7�ڰ]m�5]���Q�.�+i�6���dA�eD����뻬�Z�K	CGi-��wݝS�p��ܺ�N�u�+�:�SxJ6K�Wj�Q9�^�tཱུv�:�g],��$f�8�r�7�]���ך�}Hl�l��ZWA�Wn�V�:q�VJ�j�X;2���a%J-�rrd�ڷ���Oy����$D웯Ujrdں��E�W��d��
�h�ն�[/1�/k�y��r�9��%�/�e�'؆HfRJ�P�U�S*��QY�)�'�E�k8ԑ5g��Cb�D���9@8�A�պ�PTA�\�P�N��B�7�:&0
��V0v�vFn�s������4EZ)�m���r���`��	�xx�����]w&j�[�y�̓IV��_r���=�an�@�X34����tf;���1<W�vY"�<"�Ӄ!~{�ث�j��yv�)�f����\�Y�|��yW:[���6��͘�5#���M���"l�2нÑ��P0�q���z���5����u,Flk�����q�֎�0	��(y�]�յ���LqS��z���XwZY�4��vw&�o�3&�W�$a�d�m�O��:�d�	.�քc`��%����È�5wp���w6�)D�u4�ZOd��*��nԤ��7�Y��7wʍĠ�h���M̭��6�<��{������Rԉ��@�[�����k�vV>�ʯ���P}�V�7�RcW�F�E�G�X�f�R�a��Oki�nX�D�tە�b�k75nv��Tᣄe[�L���_luaLIc�B�^r��D�T�",�����Tynd���k��TcR���L12r�@v��M�.ݼ� ̿����
�/jX
.४1�ԫ��wV)�!y�nT]��Tw1�/[�=�8
HVW��_^�ka���I{{�Sn�źkp�J�E4�f-�4��9��V4�B86����ڼ��`1[Б�vp��4��fjT�Z��蜡�D�|�oj�}o�Ϲ��5oGL�=|�>q$���x^�0�;�X��C*R�\N��]�i�躩�dE�����i���.u6�m��@��$��M��HZ�f2�c16	)KI$�	$�%�Ii$�a$�:Z��I�IZ0VAa9�P'�gt�Sة�݉��n���a"�%�I��g ��;v���XF�{*�F�td��ήÁ����p'Q���qCV{	�l���S��Gq��N8�o�p�՘�:�n��s��di����}�� $jH1�4��&w%:���@:�A�v�f���m�)1�-�4-�qX*�:�׷W]�,�ES��k���W�Q��+��J��JBD����:�g4n�!��Yc:Ҷ+�0�=�pc�tA� �o^���,�~�/����`h}��iXagiJ��,V;[i���=�)k9,_�*B�⻳ؕ��DγH��Ջ2�M]Λ������yCy���1�����+#qp�9{�sqP�M��Q��f\�l��n���&��ì�Uո�@��au�.�x�UxZ�3�`�N0���%j��s�����[t+&�-��s��Cpos8�&����ge�+4�9ϳ[[j1�!�������@��d
Ŝ!4UҴ_T�gp��!��,{�;�꼶G^:��I�\�r�;fv[�F�����[!�^a�R����dk�l)+
��)�"���׺���X�F���*6s��������$����Ut�D�X�I_�6G"	�#�	�̼(K�Wg������Y2���[ѹد�짻9.�J�CK��E�ʭ�ǒ�6٨��v�!3z`�$��75��t^�m�4C��R��v-#k�<��V���_lk/OR���[Y����t�+D���$�6�>�k�n����tܻ-@I(Y�XR$�f�7�� H���X[�J����k��#f�h�\m,ʵ���Uy)���7��e������E�i�h�3Ptp�����yׇ;i�
z'�-J�	��Ĩ�.��/DB��j�Snu�R�Mu�:ɌM$v`+1��)��]*�.w��oZ���I���a���v�D��{�K�Q��f̵]�/$nN���k)�o$�ip���s����7��[�Ʈ�Ճ�69�E1�t4���d�C�M��*�ρ��
9k������YzAPl޵��v�Ϸ�ࠅ�8�V�4膺�OV�V��Q�d��hr�k���on�;wj'��$h|��\���@��F�p�9>�0%v�E�l�d�r�U+-��O�9��J��F���q�/b���P#��NG��d�1����v
�j����7]�.�d1u9��n�Sq�\�^k�oQ�Z�V���V�S]N�ƞ�-or�U�"���kB�o>�1y��[s��m���E�2���>��w�R��PYQjA�[A����$��h��e��]tP	;2�Tڲ.�w���(�-��\�¹�5jյd�Ɛ�	*��m]r�LS�h�	����P`��(�g�;5�.S&���f���њ���ΠI���f*�koP�Ќ���ה8�Yt�n��vr�Ia7j�m��Ȃ3U�\j��EV@�lf�4�FzU�G�4!�`G>ȕ`1LJ�q<�z��̙���a��6 �)p�8��Sm�9R�ն7��.��o��P�|/m5^R5�[Lg����W7o�oX�sYu�B�����zn��ԥG�^��f�
΅ܬ��[�����C���3��2�{��؜��Ӣ�pnHNr�rԢ1r��=�����(�ϭЮ�m��v<7�f�YQ��CU��S��]\i��,�Xh��e�,7@�R�LTc1�0��u.����E]���z�yf�`�LK�,ym4�R�n@�_�86�8+�r�;53]]]/&R�5�ZB�U�B��BA^uI����́��3b��f�L�+S���ҩ�!������x�]G����k*�gpgC�����ZUm!��IB�.n:�ܥs��Csaڻ6v�b��i7ׂ8u�H����v V>v%# ֖Z\�(H��S�d�UvyR�V�7܅ꖳEo`�D=�3���{3s1�Ж씶�T� ,I0,1�ƃj���T2�wY�P5�g����q_[T��@����´�cy־�h��iWA�W)�����(:+����qVRp��g.G����sn�F�t;��ĺ,�ϡʹ�l-�X�[6�0�ϝ�����,*��!�y��,�O8Vs�Kf�@�w*�%���&�J�d����T���̧���lJA�����b,�V�0؛dOW״t{(r�*c"���/{��Z�dN�κ�(�.��qV�@�|�V��v���p��k*��N�@�M�v9Q	mwZ��w*�L��KT�k�s�Z㵫2��u �,iQ�y`c��}!2]�5A{ڥ����>�+)�ީ �R��Ժg0�+�w��%����.�4k��oP;�v�3�F�ޚge�ɀR�F9�;�JY73��(����+>4�xo(~~�  �B����KD����
U�K�������F��M&�F\Y��n�v	�,�,���0�
33W7��1���j�8 ���$��Д�������Kp�s�d�ͮ̚Ϲp�3�D����f�Ѫ�:�
��棢���L�[�J7֝I-�Uڪ�����)a�5�X���m����`s���sb���@��X�ؒ[n@"6>"�A��%��i�v�u�3D��ү���6�pG|�<"���(������bҼw�޾�H��S��w.��۝˟v����s�������bt��wcґ�)$�Ak�[V�I	"����Pk9�э�	iKJR��P�PܢP�*���M�U���TbR�����$@�H��&�8��T�vư�E�ZZ$�R��x��rTp+L�K��-��m�[B�b(�D-�#W�]a2"��e*H�D��F��r�J�X���\4��^I�(TV+��e&&�B�@�]��Z�>7�Y��b+7p�'������嶓�k�۩�xP��#v��|����)Y=z��A�[]"�ۈ�o��tO*+8W���O���Ԯ���ck(�v'�y�G��}+����|%�Ý�*8~qB��rX�����/V�q��W˼y�\T��W����7kp�i/<��-�_��o���I;`p�:���t�k����+Pr���NGb+�Q�k[M�D0�y�&|���@�k�ךB�W���C���ywZ�tRhc�����d
��Z��^W����D9���".;s<���ކN{@��b
~^�#�{�';�P�>�~-[���&�����A�����YU˝e���xf$&�:���w�U��+�\�0��%7�9�g)
X"�=s��Įޅ�����ov���ebQ�j\�s��|;������+3��z�b�H�<���X�ц�����V�[��MsGv�3�+s}�v�=O��ܚ�u��7r5��=��S�\Z�s�d������M�ıZ'�Ɏ6�-������&�a��0*ղL�/�v�|gT@mċ�sw!Ȧ3EX�����i
�O9G<���y�o�u;VG4�@�ފ�Z7��
Hx�]�=~>P��E�Z�p{����݀�1]6�rW��޺�� ���u�/�ڙ���L�+������xW.q=|us�|_lsƒ�����p\f��T0�ȵլ*�p�_otU�9�QC,�U�wB"R�V���T��Oddu��e���S�<�};��:����U|�� uN?zQ:vK����y!��(i���z^����z���
�^�����4m����k��^�����ƓV��_�&,�{ƽ���g�����7 k�T{����s�({��;u�^n��!h>�"�z�sk�.^���
nFYi�(��M4��jJm�{&�Z�h
�q�P��w���w �[֌ׇ,���!T_���iZ4_4�7T����格i;��1pϷ�q�A_��9����d���V����7�n��ȣ`�^U^�e��:���L���G�.O�s�}d�˗����l��"帯gE���υ����iM1�d{�V!<q$��V�.��q�m�cZ{�:�z�#.�uI�y�+xɺ�!��˳���U	���A�^bY52o:��]�h�x/cTX�����y��z��gi	����~权���a�O�*��� �z�x��Fj���A����-�1#��:
Zb:ѾX}�tA��T�b�;��wԺ��+�i��mgE]ۏ�(�2���ԽF���ʧXil�1GT�(���Sn%���չ�M$?1��vṼiy�r:�-�to�����ا+�u�t/)��e��ȃ�54v��_�i΋�V�Ҙ���O�������)L���m(�[��X3!�"��@�4�tz6��bj݌�U��ڌ�Z�<����d�+��p.�'Y��m��V�����QZ�b�乍�{L���I:f��6�)����"h�]]��d����8X,itE�ynlL��)<����w�b�rT��ӭl��H�/j���5�9Jx_{�m�ײ��*��"~��%aC�����!rr��^uĴ����ne Y����C�ngJZY�}9m���q�Rh[!�Lt�x��
�.!��c�;����{	.58!U깢�F��=��,�g��yQFs{��xຏ*3��*>�K\N�t���j%<��0FmT�ؕ�tf.)iu���L���v�`UvtY���T!m���Mft��^�K���o
�X�]�ot��t�xۜ�m�nZ���.M[DX�����xuyR�����Ǣ~�8��W�K	 P��-C|~��dˁX<��ݾ]����f[���|e�"ƺj�rU,�Fm©|;�-��m�Ĉ��
q�8sP:چe�2U3wz��0b��۫P�n����y��4�MI�XR�й��Z�2�5 f�'-�w4����P���j��ٽ��eޤ{��nHUҍJJ��6�{Y�z3K�;m���l�ΈJ���¨��R�}w�T�mG�73<�����͠jKٸHT�y׫��^���=�6��q�����-J�Ȩ�-\y��)���.�2�0���*��urҕ�]e3F[n��!��+�d���r��]�D]��5�8 VR-,MP��:b7�����tbI�na��"W�w��Vɧ�P���tB�	�l��JeK���:���)�@e)�1�#!�V�
�X]; ��j���&��%ґ����7_�Kt��8[�S���N�e�^Yξ�YU{�t����>J��Z�n�PP�QuR�j����H܌��TA��R�J�HK�7r�fn\�,Ea"��[z�E�`mP��jB+hKd�.�Yye��H7*�Tn1�[M�j�D�i��V�+X�LQk!h-2\�n�d%���R�0�%��x�EH�ܡI	K6�,R�V-�YmK�E)ԗJ�\�F��4�WPF��AHHD ��2}xlɫ�_�u(|^e���**�V��b�J�VM.�2P�YE��RX�"�(×0�P���?L���۪���}"�#<ޕ��G�c?A��y��\&��ĥ�tJ�h��5W�VE���Ƶr��'-�W�Hi��f��U#=�죶lևUci�2�7+��5[u��(��\�������R����I�ժ�W�iwgKu[6.�h�"����ࡍ�NZ����T7��Ʊ�"�Q`�z�"D7k1�7X����{������]d��^��ב��βռ��
����0u��_Y8s�9�c�{@)��O�	���
�#�K� /&�w��RG�����B���낭	�|;�X�g�[�'t��|&گ'��&7]r�B��37z'����r�)G;T���⎙;���R��>>����S��t`�\�-�z�Nrn�<yѫ�%�2��,���1�d�5�ep��T�T���)�����7�8%<�]�=�����XQ�ۭ�S֮�Ĳ	��=�N��%,4��ʛN�xd�q��ޘǯ�t��jc��aߕ{�����ř�1Y� 3A�|�dL��ؓ���wN�'@�^{č�����/5�+�:��rZ�u�7HQOS�WV��|���H�������2W ;k:'ho(���Î��'���ǲ��{���5DJ4d�6����J�R�Z����ޟMg:*�%�@�Z�9�q�8�|�u�5�Tu��Dh+HQ���!F����vU�
(�e<�����|�UƩC�ڪ6�y*����^΂�-QF�IU��z�R���UGZ8�-Q�r�(����xuо՟l��9�Wdf�ہ�R�N�_5�g�`>QK�!Y��3��v�DS�Q鵖�eKk�����ǽ�%h(;p%y������jrQ䠛֤�s۪-+HUtj�i+�UBڠZ*��a��+�Q�J+V��u��~���Tw�����(�Uj��PC�U_4B� �s�n��׽⫭R��
2�E�֪�jUQ�5EBҫ�UJ���K��Uj����Xh0zkMu��Tks)Te���(�A����߽���mZ�¨��h�%m��Tl�]UVҫMUJ�@s����[8��h�(�-�*8�^+��Z/��*���u�1���h�҂��i
-*�MVd*��Q���*�%h�o��g]�U̪�5G�ڬ5Aĭ�U[T�Q抭�e�cy�����TB����G� |�
�Ҩ�U�>j���U�*���
��q�w��_�X�]����ch���̷"yL��#_Ȍ��S�w֍!�x���s�������B����	Uֈ�j��k܅��Aƫ�[A���]���9�Ua���!���5Tq �j%Q��:�q���:�j�
!u�V���u���h�=�U
��-(P�A�J(�^��(�y
1�ƩC}0�AƍfYJ�TQ����QiZ�QV�e��+����t��������h(j� @�Ej�i����-
�T@'eփ;�5�n�4�j�C���P|�u�>h(,j��PD��>j����.;���Q��WZ+�Z(�cR�J!֨3�a
:�A���(V�U߻�UQmUJ�mQ��L�@��z�TO�y+�ϡTi��5Tl��}XǾ���5� W����#U�x�i�\M!ƨ9^�D4�-�S����$(���~�����w��SJ�O��-�������&*�c�ff�8�ж�j�%��߀A�����ٔ2���n�%���T�9׳z"���5ݮ��	}���Y��kj5�7؏.��G��O/B>j���a��IR}M��Qۂ��9+�^v!7�l^��|Mwn��}̅|��ͣ���'�-��h��]#�r��V쁊Y����uwwƼ�B�R��b[ru8��ݗ�{i7�{� C�ڟ�������tA�̏5�֡��Bd����]J��u�6���Er����*���<2�?eykw�+��0Fl(
2��K�j%>m�K5���=Wo1��Xj�/�Q�JFՅn�l��y����D��TB{,}]U�5��F�ӥ�{�6�F�ʺ��^�ENM�m5;4	���������������_��5��=�ݑk�X���ZQC6F�ve��<�N�M����Ub�n:M.�Fek�u:�S�t\����z^k
�P���̗�2��o��&� ����;�S���B{�O�_�F��CYi�~7*����өOD��Eã��4�ox�'إ�Ǘj�N����r\.�뜧x�3��q�Ř�{�xx%]���W� �==�~�g�2�"p�C1�*�>﷗�7�%��#�/�uq���WI-��o!=<�S홅�����-�� �c�[�g�e�8�so�m�@��z9`����tϨ���۱Rpލ��f�A���O^sӝz9i#������ݗK�Tx��m��$�ml��E�r^���ˇ� �z���N<�:���6;��.F��˗]&&[t�T�
���Ng��b@��S��KR�2tN��)D���y@2��(;m;Z�"�u�F����|JZt[�g�lu�]���ۗs�<�-�j�	c1[�N����k�p�yv8Fw�):H����s��F����k��*sMm[c�u�]�2��Hl�J��W��٘lV#�J�����sy�u���~z�ޯ�?"d��X��Rec��L��Xh,�G[���wF��N�+�cEغ��]���qZUrH��9yqVGP�`�B 8�H�Je�%a�x0`��u-�#���ʄ��p��3�^Eh�u.P�i�P��"�rL�ʺ�ET���a��[��Sp0�ϮIx�6��L��tpU��d��*B2�	�uwe% r���H����90+�Ǘ��iyٽosǿ`��y (��<�AU�"��M��JihED�2DE�D#�!m(�#����"
B(�Z����)$�-ܢ1����dZP�B�J*�F�E���X�H�S)���V��Z�B�MQ���$H���DYJ"��dSa�P�UswVIPH�0�TQh��x{��\��&�|��1��"i��m��s[|?a�xx��}+>��ّ����/=�B+����Vk����3Y(K�S�Hu���s
��=Nw��wZ���+;>�6�-=�ُ�m`]���w"9�.l�1�JI&�Ř��qhl��Q=lX���v�,:�=��D�K�|=k��%]<2M[/0�֋œ�j��c c�p����=āJz�H��s��n��o�{�{Í*s}]�:4�̊��$���BQ�v�P�5P%��{o#�	�8)oY�[�<��P��#�ozn��^�yfO),�f!�⫌�5�.��e�5����V�;CO�>�ݪq�Y��C�~OZ`߃ ��t �-ru*�1�L�t��P �7B$���E��R;;���9���Һ���6�n�g ��iIj�>����cz�F;j��L�}���u��C왰��y�㘽���7�Bo�k�S}z[]^tH�~{�g���lR�j]`��6UC<�zl��U��g������sB�<�z"g4F[p)g]`T��/u���2�LӢ]��f�:�o�ЅF<�z���g�LV�k�����%�D��u����M�-��:����3Y���{��s|��ߖ�f�_7	�:!�5V,�Qw���L!
�"��Zwq2����C^��Z�5���&WB�xxŭ;��'w}�3D�5~�S/[�sZTH�[,Z�[s���[��}��7N��AD^�}���Vb{L�"�������,PY�ի^���Իt60. ��I��i����6��^j*nN�9i6� xxJwͨ�g]\Pl�ژ��y�=��|4��>�u.`�f������.�rf�.���OCV7Lm�/O4w�zVT�ǳ�ch�{�)�n;�60�	\��i��hww����8m9����P��ۨd�Ֆ����,0S�K�{�6	�YI�t��*
�5��ײk(�*� X+�w]��}����ך�+f�Zp�q�w�7��=�{wo| �Ol���~5�/w{w�v	�3�T�V!e�y��F�:��g_Z5�,��~�I�'�`�b�9��w�.�>��%�U�Y1�EN�ngtC�ꌙ�!���������d�-2T��h�KY�"WB�������ޗ��Ĩ�����2u�3Z.����x�;c
�w�cu�فe� ��b�������N���M���=��)�	�VoM��3_^�\TTs���W\֬��v���D����{��L�$f<j,Qf�>O��"�8����^g�����4Y�x�Rtu=���pfL=�q�5�+���8�+C.�KV��;�;>ح����l���Q��S��@�n�M�wkg�y�L9<��(�w�OeN�ݹ"�uS��1�R4�47��kN�͖��'#h=J2b�r���s����Ϲ�}#���B�V����{1E���F{ƕ{�8�ڽ�u��!S�}��1�T�9�S�Z#t��7%55���gmfm�s����{o���1�"8w2!�.����=3��8߆c��$��V�u"R���KPn3R����ԯ�}p8S��kx{��&���s(=���������ݫLq-h�r"w,:���Y�FK�=���g�����y'�����r�l�#��]�����2��/̈́�g&h6�P1D��׃n�:i#�yG��u���{�����"�G���Xy���;�[�e��{�N��ٳ�k6`����e�^�mf>}�'4�c��!#�im��� ����p����$���o�~K~�{�d�l2���#�ΣH[c(ՠ;Ag�+
��$6]O�ٸ�����[qh���2df�v��� ,��QV�fSzR�'�Y�&p�z���ܹ�K��k�4g�yt����&�p�
Q�>w�g��L1��?m�7�#Ձ���x*�mԑ3��z�w���@LvVP诖3Xm�bK�3J^"�P�f��v�7�tZ�WS���;9�S7��T��۱d'gЩ
w4��sp]�{@�>X�ju����-h��K�ݪqj�e�1r�^�rƝ�h6Lx3�U�gw���(�U�zB�������t���6~�;,X`���t�M���z�؅W	�3�j|����qi2��.8��sB`�Ɉ��޿�]f$'`��O ��f���&]��� &����B�1t����ș֕���H�d2Y�QE&�iP� ��Ѓ��Gk,dm]]&�&#�c�E۬6gʰ;��9�UZ kO�h2��B�8�ʏ27�o;Ɋlڢ��P��;*�9N�ѫ�$�2�۔�Q$�I�I$�Fi����\z� Zn+%BJUV���KKRKI��
�ӈ�Ѝ���V&!�%��7#T[�*$cQRȩ)��*�!j �Ba��ĘfX������V2!l�$"�J[��QDB�&H�6��[�*q(��&aip�"�
���cr*�7MK����ݍ�c��Z\�a:nV$�����z��׾�H���?J�Q���'���2Mwu�q�G xTWO�V<ݍ��[��S�����y�}Xq�8�uPlh�{�V�s:���cæP���܋>C}�J��,�e��>�k5����ɣ�1,03lL����p��I�q���΅m���KJ��^��jeJ��bIC�L�J��V�V���� �٧pm�v�3%\�_{��������@����,�t'�O`ك���Ӄ���ullU*���� �<9�X8�����;�*�Gq{�����2��%��wf����7u-t#6z�Y�T�)I�s0����v���"�fLW�Z+�/��1{ۄ����9�Թ��J1��.��_����4WXG���������ۖ3���bL=��q���Wen���yy�V:M��`䵈�σ�ҤR��<�������^Z__�1�rҙF��On�sGK���uh�]�kmQ���,���W/����`P�F'*��J���
��7���Wv�pj9������
�R�=��Q����b&�q��a�m�<����}DuR4�F];��-m�
B��ә>���6��ˇ�Gj�����x��>13B�`(f,�ø5b�x^\@�R�KM���9B{W���3ں�a�q���M�������)4�ע
��<�-	�>�n�����޹"��eq�/k�\A�;�8s@�;xh�R�B�9bM��{��R�-����.2���{�(Fb\�j�ak�4�ۏ�����WS�,�,�$��J����N�5f{�}���||��%'9�f��R�6�����vi��bk�OU�=�����"�=���-ӏ��Oa,��}uo�T��������R��i�#F)�l����C�}��Y�\�`��Y;H����k�8�F�;r�O�����X����g�?mcT����f眏�*��#~�J��z�]���]��pm?c2��S:�f��ݽ�ם��t]VP�d�W̫��Lf=%dGS�8��q�w����Ŵ� �+��EHl疭�u���7������s��M>�5tz�@�ױ�(�Oj�T����8Q���(�Q^��)�{C�)w5'���OHR�Z�Zo�������}Yf�X�MT��ͦ�����48���6�R��2<��*�6~���~�GㆲZ�9Fe��oޮ8I�LKE,q�h��[�&&���/]��Fw�0�m7bv���.q*��;������L�ٺ��� v%a܉��dd5�d(P'(��ǋ�
;���e=ɷ�z���sRI~�����j����7(qM)��ʬeTi�*��K�{ѥ��l�m��C&b�:�����g>�ש�C��i�P�e:�y��������o��ZM�e��"OMa��9o��&S��i��]�Y�ӧN�z�u���v��CR��h�z�x���w���|��W]�U5t+Em
w�O���EW�	�9�У.)^�<�F�i� tlx^�cp���0�f�pc����/nbG���Ɲ��(nF�p:�Q���R?5�Y�	G��-���.9:��uL�\卹1���2JUmYW-�s[{�����bԎ���<�P����M�P��Fw�㞲`�����4ChѢ�ͅƬVa�i߻.m�p�� ���I$�4�A�[/�ŏ'�*�ٞk�Ў��3��;�kЎZ�a��Mf멧(e�_ONN��N�\R�n���Z��ƛ��:m�3�K���m�[�6��w����/}6�p^&��I���m�'s��^7�4a�R31U�k|jf���������*�ԅ�
�8�Y�t�fm+&��	x�u{/I@�X2�C��CN:܉�<7�[0��Ji�u��Q��o�<<�&ֈ9�0��c­W�	�p���kV�����N�vc�6؈�������y���nTR��{^�@j|2$z��l8�d���@��xi�8��C��ҁc�A��Q�5l�dfH�}�[g�v�UP�δg^�KϽ�`4��A����4R0&h���.{U_�GI��VۍJ�i�u�f�6�X��y�I�Y�/x��b簈�Y淮X�Q�`�b"������l�
3�U������Pb_Z�E2��5}�K�Nb�!��x��:����1ً�����;v6��fo+tY�g��u*7xg�#�j��w�8��tnj&� ���[f���>T�VKMJ�j�]`޾��ٸh�	B�V�`��a �a7$/v�F���v�A;㽛�v�'�f��ոf�a�ȃ���̃���[Hi�p�ht�h]�i4󕺁��/�3�ͫ�ɑI7��Z�Ł���'ymj�!�K��t��r��3s�<�6�&��T��
1���^ z�!���l�Q�|<���K#�����K�)kw���_0���56��Ǥ�G�i�2���V�����@��ܛ�B��-BԵ@��}S@	��+9�ct�*���U!�B
�ͱ�YT�Tv�;[D��zf>e9�!����Ǻڕ8�'bꓮ��4:��*2I�ff�D1�tX�����m��M��e1/L�m��&$L��ba��2��$�Z��7v,n��.�"�B��S7(�R(�1t�2G�7v�U�
]�۔�8`�U�U��ZjIDT\�˅0��3�&$a!(̖����,���*�?4iRB3�k�T�4Q(�*�Ez"izA��a��OJuS�����i��� 5�{��d��d	2>�,tɮ�H�5��~��b���(h՟vH�#�c������'z	�Ӫfjh�b�I:�9�}�w��<M�ǅ��~4��2{�Gq����k��r������|E����Ay�kӯZ6�9���\��)�$�7�_f�Mr��1�[�u�Qo����3��sgR�o�ow�J䇑y�[��ִ�K��ۯc��q���^&�-����
���|��������v�"�uw��V �hp�@zv�}��>2����L��m|�	��8;��|:�)�7	�l��5�_tm�渓��Y�,�B�:�.��-����9�Ekɇq�L�99�[{�Ǻ���]�wXT��#V��É��i��+��`ȕ7�8'ꂀ�X�cu�r�Ǉ�7ܸ}�wZM�e:�|����l]l��<|��w�2֜5�)�������K��p�]^��f��}0�$��]�b��Ѡ�(d2��4;z�x֦���]CC�1��]ey�����P]bi�5�:�s�6� U9`s�G�I�f�}�.:�e['Mb�zr�o�{�S�'��z*:FF@Q�A���}����}[EClC�ǥq2�-��<��}�k5���kE{�>A�
g���������V>����L����1�k��=�{�=�vF�ËL��F����KYQp8}��h�49���ѳYe������&�����e&'����s��ֻn�1�s���ӎ�ne���o5���B3R�se�Mf|�B�w/.���a�;k�yt�������^F�)��.l�ajL=կq�ʹ�{-pvMt�<J�3���%�pj�Jo��+=��=~C�̺��ñ�Z܍��l�پN��#��g�b�7��m�۶Lo[�ta�E�DK�#}���|�˹���d=٦�12�D�ש�Z;A��gG�6 VɊ1����}?p�/��0�+����l}N���Uhy�fk��s~��2ٹ����z��<�~�S}S�;#ꂰ1�h�����AI�}������F� }��2�Zk�[���q�����*�����u�ā�J��Z��Q�u�b#�4�s�G�C�7eY��;7�0�vL�Ŝ#��t�]�m��x{��~�>�~�Ϸ'�3ё�
�?=�\��\��>��T��ڶ�~%g�ξy��t�þ�.V�:��e5�Xk��{c[w�A�5�Y5�#������7����]���\�m�5���㾙�p��p���,1U�(G��ru�XtT6���Fڱ1 �X�w�9��g���^=�T�Ƽ
f�I�^5=#�J�����4���szލzi��� 숃��P�ׅ��:;k���	Xmy���:�T��ڍ�":�.�1B0�"m3E��<��t��"6�h�A
�/������U	x�q�g�Վ���m���7�[���]oؓ�4��IF�WS�Ε��=t��w�`���Z]bZ-cr�zw�9}���t�P�]1�4����N���ｳ{=t�N�vj��,_���B�Q7WQh�H����x1K���g�xցݰ푐Ѡ�&��j�*��µ}=^5�~�V,}����\'9!���p��U�~l��Y�V��d"���v��on�t�T���W1g%�wra�Vp�Mf6� .a�Lw 2.����ǩ����p������{ܭ.ᡀq���-r���*���P���Vhâ����NG��T�+���?S������2o�Ч:;cKn�q�tQ�x�O7�Ʌd\(�ؘ��L�GA����}�vqZ�u�a����ճ{�s�+�����os��ӷ�+����<>���Ί���,O��n�Ӂ^c��k8C�hN&.eۏH��p/�X�K��!7S����;'/��<缕Y�E��Z������>�1� �7J��'r�o�{ބ�;��|�J�CY�]I����1��r�=+Wڨ�*V�}��w����*/*C��f����<*�N���Ϯ�F�����`��**���n��#Ϥa��"�É��j���֢��dy/y��zv�W���t/÷��� �B�ǖ���M�]++kaDt�eE�6�s��t]�u�`��M�=WY ����Cד=�牣��8�;{�|���`"���:�T{�ƅ�����b8�� f<H{����v�gV��'P�8V8ݻě��������GFA�kӫ�q���:�T%������R�\k�N�m�e5�{u���h�[Xr�M:6�L�ά���ν=+�/�z�}A��d��p��z\�}I��L���-�_���D���ܨ��%��	��1��!Q�>Wk�U�b���"9fne�;N�6i���ן;w����}�ҠDS�p,9
)�
uA�ugR�A���Ѡń*��l4.\�"oq���d�J�}Lf$�E0�=�<�p����Ft��L�bv´��5z�{�w��}�y����K�MCvJ0����{�Et(;N(t����� 3!�װ��5Hh��,�c�:�|E[}:���Dn>�D]w*��x�%n��"m$�lN`���I�Y����2��������� �b��ي�m�]��\���kJ�y�#�sY�m/;��ZZ[j�*k����^���>�*B�>OU�b��C��	s�4T��֪���\(�'�U��}�g�F!�+�^8���'e2WXu�s4D��G�� ֬���L��Dul�H��@M��fd�h�	�B�vˋ��j�*���7Z�vu�|1�
Bab����p�f^�cR9�e��ǁ�-+
�)
#�h�Ċ&��a�:��6�b�1��|��pg_q��J�c����Bw.t�#���WK8!�m��z�%���B�c�.jS��d���bT%p���8�������T%R��d�/sI��9�&��K��R�//��HY�4�kE#�7f>X�)!W��[4�T�[��7�ӧ�mj��l^����@BO������.��̩Vj�����s0Q}ga+���v�"��,H�i7���$1X��õӡ�w�!�2�]z�6�������N��pL��|��7t��O��L
�;4��õ��Q�N]�����	6�vwN����O��t2s�3i�0���a��u�[�� k+7*��Efm��J��۽��ҹ�zۧ��L�:�qs�Χ�І���5�"�ZZ�֢*!i)3	rP��K�f�$�Y��Ȫ
�)��H����e�)H�KRT)DC̢*bR�a���\�T0,�H�2wX-�0e�l�rSp��J\�!��#Z�2�UiK�*� �.Z]�R�U�z������Um����j}���sK�/��e�o�G��"}�1H����8ޝU6l�g����"*G��1p1s����q�ݖ�=���i���Qr��At����Á��	�T2f�OO<�o��8�˲�t����YYM8\���;˥8�f�ס��Zs;u�����p7��ٓh�ۇ�G�I��4M����Lg_4q���.�+9��j����Iu�ER*�@�CDMV�Kn��kSCc�:nxldn}]>k���+��V��� d��n1�$�I�6��0��5LSaBs �G����'�f���U�zw��g��j�6Gr~R7XZ��F���kp��X4D�^G�=3�gh{����3X�v�;�m���2����~O=�B8z�k!`�bc'O
�5�]�5f�>�k2�{�s�Φ��{6���7*�+�i�B�f�a@2H�Q�;^�s]_N{<��1<�p�.��`�q��_��ɞ�>k�Z��;+ݕ��Ms�����}�m���ZjVg^����g�()n]a��s�up#�|}��7��ͻ��c��2\.c����m�@���EV��#��r��:���-ZMr�������G�0�y�j��m@���3�7�#M.8U���8~1l�_y�u�gp��jq��w�b�]������*ڨ� d%5�����[���'�CH`ЇC����5�\��>��6'�8�P��emѩ����}�o~�6�S�O30�Z\�w&9�.g˟Y��]^a���/\��-/8˝�i�+b
m�!o�)�P�~V]]4�*qW̚/ʩ���ݓٷ:�},��;�Ut��Y4�mx�)u�cy߭���2�%�:�9��=CW0���̲3[]�X�ɗ��I�_eN����Ob8C���s3�9M��~�A���q��GO�t��Fǅ�q�'�d�6��5�¸O�E;5��B��
cxW/6%E�e�G@�,G)��9��SZ�-<�_c7^�\���%y��o�2���u�Noߡ��7�NoZ�\;=E"[.�/S#Z#1n�쎯�p����Dpb�����N�J䔣�M�mʤ���׃E�qd��9��C�r㿦�>�Bmwn(�������:��_�>��}r*Df��D��fN Ue��j��ƃY�L��C�ǹ�^�՚c��=F}��-���ז�G�� ה
6qFur����zֹ��\����&^6���^e��]���N�7+p�ain��=�9����5<�7	F>ђ�W�D���4VP`|�/�p7�o{����<���}�gg��D�)�0D8�Qn�T8-+��� u6�k+�x���n�;��������4�#�*��R�$��x������̲�N���(��:�e����U��}�}^���0���߂�}���%���h��Y`��Ʊ�[��	w~����s��hhӦ���\s�_��<�p��9���hS�qK*8Ԓ�hTt
�����a)d�i.a�cu����^j�w�ˤ�9t-���l�̯$7� EG�xǤ\��|�7�q�ƹ�l��[7��{��>0��M��n���
�+ƬR���5��>˪�pX�\pX�G
�?!Lx|,���Uו�k�u�vGP�n�VЫ=p�����Ρe���T1pt����{��6Gp��O���-2\',�k�gcσ�#�/��=~���:�VZ�gǵ�L�i0F���G�����Ӝ�345n�=jܱ,T�Z�ʼh�qo+��5�rC�A3B���=��h��;��I�
yA�*L�p��j	s�Zr�����n��^�}*(B��T�[�]5��f��AǯU�u4�tfmޱ��� �/S�S{3H�7>7"�J'�#�����������[͌s�"d
�")ႬK,;�Ԓ�c�ɾS�`���&�,�{G`y������\>�B3�Z��a9+C��Ύ_���ˤ��9��!��@�P| lDj��:�q�cL��k� �j��Lh���걸~���HR��C�DS�y�p�]���\7�춬��h���缽�Ӯ�T(
������֫��$8xb��iP�{2�LHi6���s����99�n�"m�fݵn��&S��u�k��3�8poL�����:*���x�P��0����Z:�����/l�wr�J�.��f�J�o2�1��ײTݮI;�1i�u�!�xS����{wZ����|�qL�__���ś��˛��>ώ͝6g�em�s���ś헔�np�/��*I�M!X��N��=���Q�����O�`C�B����p��1�ه��J�nq|�.7�َ��v�1(�9g��E=���?+5�6tf��~xj�AL^-�7��W�N�Vi�/�V���R�{gD�}�п�q�#(.��oX-�m4��"ˎ�WF��3Q��'t�P��Y(I�u8��7Ojh�^��m���7O�|�?�\�mI��QP�%@ۋ�&���W�jz�ni�������V	I�t��Z�{J����:���{BJ;Z=⺦Ry,�d��ͼ��4�{�����̒�0���`[�=	��W�a����yJ��S�6I�<��ʁӾ�\����ݡRe�R�I�S׮K��8�K;��}�]*t���/������S�.���t�Dۭ�2b�v1�2䌗�Kriи%+�PK��������.Qdۛ�&�6 b�3�7 BexM#�X��:��޶mf��}6͔���E���v[���g�u�筊#(��A��[(1�\@�u��ƹ��RWy��0���9�[}$N�̾�}�W
8cN �m�P�S�0�{�-�a�mЮs�.VlGS�M�יv𼃈��@t0�:��
Ê�+��4�HS�08Pie��vc��3���˅Q-H���eY>
�5*�V3��L�+ a���L�u�M������4�"��q�B�J˫�0@� ԅ���+2P(�Z�*���H��)�*�fӊ��	CHT�8"��U�ϳ)���qF�D2F�X�d�T	�&]��DB�J�"�F�.�h ��+�iYt鴑/�x�A��ֲ�y����Wu{ytw~���!iH��L� ܉��--")i��Eԅ�K��9��m�F�K�ʱi��*�
�&�.)3	�4�%jJBH�J�\��Y.����125	v��%������M�����Hb����ͷ��nVs�r`��;b�,;lM�e(a��HWS�IĒ�KC�g-�UY����~�gdA�^@t$`�j�]u�B�ٵ�k`�>��|>�ԥ��J#�
=���X��~ĉ����l_:,�'��6�8 J�le�%��S5�x�گ*x��p�ԮP�N�K�Мf�H�NV����H�ɳo��L���|�c|���v��)>�TZ�^�+���0d��c�Y��Z��_�ڏ�.�v����1p*'swcA�K9:%�;ʠEl��ڴ�������( ӛ7�����*��o룙\<k2�綖�'�|��gpx�&��^�L,�
9\sF�z�[{�X�ɦ�>DDr�u���0;~/������J�~�3
^�^FP�U��<�oz���9E��n�R�Gc[��p����m�xt���><�0�ܸJ5ӭ|uMA�ɾ�2)Z֟b	��ɥ�23gfU+0CL�3��BMc���{n	`��X��r����v8t5a�T���5�k�wr���R�^��}�;�gϏ�$T�WS$^�Uұh��]�&־�jc��&%��9OƟ�+���ۑ5X��9d7Ѵ�'E���2��UR� �3Q��� 5�{}�Y]H�:,���t��b0-1��5,��[� ���h�Sɼ���oEb�Z�v�er���A]��F��F�q:,��.X�D�O��YF6��+�������N�윫iW�����u��Zұ�0���\Gi���Kv�yi"�}��W�v����Q N��7\�V���7e����H\����m�=;k�~�(�32����g��=�ضO5[t
��
��t�����3o�{�C����`��Q`묦��'�z�KZ'�%ۧ�ؽ���u]5�w�W��6w���<֛=1��ۗ<v�+A�#CYB�#�i&/q�L��xAv<ϖy��=�+�,%"��ی��8�8�K�y	�[�}��C���):��v�D�߾���_h�߶�*����)���L����d�z�7��U>ܿs�I+,�"ٱFޮd I�򖹻{z���z))�F+WM��ȝ^��ܞRf���U�O���V��d
�Tz��G�־.Q^\�\��Nk��;"�d�4>����<j����������iQ����O�~{$�D+��K׭����Tt룈nQ:���ޔ���<+�{a��IF���{+dO�qMY��uw��.��;�/o��:qf�
vgbi�^4b�&�Y��,��׭Rݦ���D���5�ub�tv��fm���Id�^i�;�= 0d.�Ml�ת�5���nv���<6�v�<~o]�黼<D2��@M��+<M�r\�zB�ۣ&�c��r��=���t�U�m�J�c�y��j
�WH���Z����gE�����Wf���Eq�}�KFt���J�M��ҧۆ��g�Ek�ޒ�{Z�4�.��FOx��]fx4�irb��kf�z�	{Ժ.fDj�����^Y%�^ƽ17ѭy`y;�����yo>xa1/O�^;�r�a�P����>[dM�9�Y�L*�5Ʀ[xn����,�b_�u�����o�М����ʱ݁�i��R������ro(���yskAJgk��5s����퍿m��$j���9�h�����4&�*I;�����w�r�C��4�i6����K�/r��W�[F�]�m��ýi�y":��������\�V�}lO�ؚ����y4�r٣����)���uLSa��9������j�b���7�#jF���Β�o"�B�h����[ڳ}�������V�=��;u�S���[Y՜�ٮPKk���ז��gp~�ڸz��GJ'{B�J{�G��O��cѾ#o]e\��R����܆3`4�U�Ҝ��*�؎Y��ie�L���|n��&�b��|﯌ACD���7�B��c��PYQjK�ǉӺM	/6؇Z%��1�J}dϴ�C��F�f�Ef���ړ�.�%M�I���(Q
=�
Ɠ�xUI5Zhw8+Dd�k�q_b]�ˮ�8��[���z�igMk!�r`�nZĨ��qp�Mlu&+�5,V���ǂoż��mk��Xr�3w���x���륒Z#���W{���B�ГvB���^�v�a��X�
Ymm�sAv���R��K�Po���0��4��yBR�q���D\$6��t�se���U�R`3#�)9v�Lf���Ԇ��h��QU�f��R�(�F�S�x�qt.�6�4��U��V52�]b��̉X
R$�2�
t��YtrPVAD<xbˊ�Lqՠ%\W��4j�����Lj�x~�N�$l���4գ@%1���S�ǘ^4������<e���Czç��z�&�(�Q ��X��ы��="�Il���Ip�b[F�1���յc]ˡ��X� �fB+���Њ4)PKHY�k)�������f0�$���1��X�V�\ j]�$�]f0���]ݶ��*X�KW	=��#[���#�	��ܗrױ	9�{�K�6�Q�U�)��[[/Bη�c��h^�=6��;���I�7J��Z^.nr{s������BFNIro�x�j�nG��U�w�D�l	�[�����y�>t:�����V���=�KZ�~�+]d���E�ԉ���\/�����pkw���٬�;�k�nK�����§kpY��0�f�o����w3�gշ�08�ұ3b
���	PIo��u�;���-����q�y�\o�E�n����֑qL��Ƅki�&�f�!�5���T#���D�C���+��0���L��/��Cx"�$2�m�@��ǹ�\{G��ls]<|J����<u���EB�Vq�sM�>� y�Ͷ���Ղ�c��i���:�hwqp�{'#ץww~����s�8O~% ��aφj(P��cs6vEw�=����3za�m%�!80eX���a��S^P�A.y��{��a�,hS�h�o��oC	��5�*���-�;�C���zH\m�.y���ou��E$'n�����n����������T���N�w���N�ٳt��K�g�xw"�D[�pg%�v�{�
_s��b�}{[��c���ڕ�Y�5�YzX�EJ9����[��˵���\�#䖄ʏ \��x;��6�T��Aײ���a�[���a��34�p疒oL|܎mxC*r9��$V|�w�Y�]{��t�-��c�䌞���n�WL�t��k�����n���a[��]�o=�״gi�-�\�ч1��<=���߾_�CEf�t#HfUKU�������l�ʙ�廡�Hv���P�ۺ�܍,�����弙|9t��}���{�s��xT��/��<�"�\��+f��ݷ��{�K&yD��#q̖�-��:Q��j+ʎ�S�;Ρ�l��V�޷��x8��%e�8���e�PZ��h�I�9��P�x!����{�7��R�'U��W�w"Ҹ?�c��m�Bb�$�\�b��췺�F��;�H{#]RH[&�__M�gKj�!�<�*�ҥKqIۛ�p�E�;��	G��;W���D���c\���֌X��ս�����{ݏ�-���\��Nۼ��Ң�)�#���PS�(d�V�,��]=��&p8%7����nl=��I��8�C�]-[YCߏ�#�����V�O��Yk�5&`M��y�q81��v�����ŷ2X\#���=�x�߮�p�}�aи[�Tፋ:�ؕ�ea���w�S�C�ܬ��Mݿw���hQ?q��`{��9$��w��0�E)�C�| 4��׾>��,�L=��%bɀጥ��]�7�*�,#���D.M�e�_t��&�Vf\�.T��:|�|���,|L�^z�EyxϭT�e:�}S�(�s{�rn�v+��k������n�J���W��FW��51����>�v��yM�������}ޔ!��Ǯ����gϧ~�~˴�qt���� �&K���E{����O:�i�D�,��Hà�Qu��z�N�{�R�B��������i�XlB�Y�R�Ƽ\����F������y����xk�y��Wٕ��"x�#b��������P�0N��ڄJ��YH��\%6�v���@�{үa�7�f���\��}�{����@��M.}W�墽0�ڱ���Һ�>�#}h{�&P��w0�4�n�����&����As[{{���s_`��>3u3�曕�V�\�=�_%����N�c�񠶵.$�<��'�0toum�X+o�X�	
r��g��<^�W;����.C������ޠ�3�����o�2蠭������Iݪp\M�y���;!����[*����mu��%]9w�^�`A��6�󗫺�Qs)'�vVQ�jum��8D�����i�A�䣌V䆲�!Ã�n��wRv�|�m2^����V.R�(�C��r`��Z�WX���1��[B�=ZrJ�!,�B��n�n݈(a�����VT�ĝ�u��S��u����/M�vTΊ�N,Cst��ၜ��e�{:
�ڏAU�%�p7�۽��)M��@��ef�7Ρ�vd8���v�RH�˗k�d���#��{@TG9��%ڭ6	b����!6EJ	R\�g.]�V$�s@�#R�a�7K��L�2Lvp@H��,�3���.�	%YV1��F�_8n��E��伦��hnv�V�5�Uh�!�0N�&�L��̤f �WWN���vQ9��@���7F<IB2R�PUlCi��è���f��ޤ�m��m�N�i��AF�����բ�jL]��.��ڍ�j��7�,#�����IWa���L�u� �\�nT���eU����wh����\bJq"ˋWp�ִ�D�iY"�1w$UX�v2)���,���$E�� ��F�S2��V0E.Ed��؈��iŒ����A���*�d-�KVԦ&�,�?�ֹ�L>̫��J��QN�8.1��m�{�Ro?�?��4/����ꚻf7@�9���m���6��+�oc���ؽ��=k�.���xǢ|�>g3-X~�8�9���z�[.�r��ŷ������X�0����.k��V��0kk�V �k01��3�)'X�����!&W`k��1����,}��wpƘ��ƪ9*�e:������r�3��:��Q0%�3���;��M�����y�b��`�=�zW���8��B���}9�V�u���V^�@��yG,$��o�.�W[t�a����۫�Uws�]+n��v��CB�1zF��C�c0�_'����F:���)���V!"�.S�W�8푯��f�wo�`\����i㜹���Ӄ��t�9�w
���v�ǳ�X߇��sE�h
���m+�}��\���c�>^~���n��ʯ%�2q�;�|��sP�%���J�v2�5�sK��i�q��]�t��+^.�M6Ө;�cct</W�oO<�ݸל^u���1痍� A����Qy;&wk;�����4�:x�˹�2�1iv��)ʝ�~�)�>��򃠀!DyUǞ�,Q߄�D����qQ��L�N�Nt�6m_�b���5JiX�9��Sz͎xF�Tڙx}�<iY����[�Lq��*B�ҳy�lZ�ӛN�0��1ܧ�ƽ�H~D=�I���[�K�'�vG\g�4������$+�W�3�p��B/t�i�Nr��=b�)���d�:J냕�`��+9Z��եY5&Sp�*�\Q�+4�6��ޔݦ�u�坉C^�1.��|�_?<O./,��5c���Y����N;�Y�t^|�lRJ��ZUr�_S���t�=����Ř�Z�ogFʵmH!�m�����W�y��lqH�8X�;�="qP��R.�i�K��T�z����$����.AS.iHfwg	X���ćf⃉#,�m��ۓu�nUQ���;�����3���
��1u���MgP�W]���R�[i�r��	��Q�`u|+�7@��!���C����׻&��՝���$����̡�'&.:�G4y�5�B���o:^�w'Y��~��b�������ylk�Db�1TJ�R���~u�N|+8��cS�����9�a&L]|��A��B���W�ˎ�{ksY��x���K1� ߫e�|	Ox�f����S�x��7,�w��l7�����O_�<7f��B�-Wr�k\FV��Bf�v���F$��
8���U��2��Y��Jd�1������xȗ`�bB��J�6�w�y]k�
 �7��Ek��2W,|ۇ�)q缵�M��4ۇ�k1��O��ng�#��M�ю���c��Iq�3:�<�A������w�<�$�5�G:wQ�]-��9ү�@kVd�ohh@��O$���샷N­�����혖��OH���I<�*��:]-iz8:
!nR>�.Sxy�0IE|�{2��=��xZ�8���b], ȍ��l�"�k+'[PT�����%s���"p���$uʽ��0�W��4/���ݵ�G��)0��#�:�[�&��@�VVu:�]Sx�:�ɸ������Og�~�0�*}ni�@�j��6*g����'8F�滝1����W�LO��[)߳:�vk�3dTH\�����یi�G^�`kc7v]�5$;�jt�=�舖�Q��2��h�h�y@չ��6�+43f�t۪[E�*�f%���bM��p��K-XE��V�I�D-ip�i,X���\Xo\�G��l
��`G�Bڿ}�Y���w<~}�5��N������/B�������>��o�Qy3��%�˹éJn��!���R�_-yX���ӝ��;D+��#-��{E�暤E*E]�V5%g��ܰ\l�n��a੷���G����!Ɣ��u?*}X+mf����vѻ.�boOB��V���]���素�y�"k�*\�(������fS��(�����*)�ZGd0�r�ь�t���
�)��:-zۡɔI��ۦ�
�w��4����N.�U��צ��&���TD3kh�Dn7Ǭ����������P��x���WJ��e.����krj��q+=}XjnA�v�FVH��ʃ�ٖ�8n�3#:�K��2�P�ۇ�ã(�B�q��iQ�}������C;U6��=��w4Z�5a8bP��������Q)U�����4���V7Q����w���ú�+HZ@��.K��W9�ZOt��p��;�\��(�e�����)Q��6�se��9v�Y��p)xq�z�eF.�v�d׎����cؔ��'n�&f�M��e��i�E�]�]�$'��\��Jڊ,VR�)n��Q�%ŬKE�Zc�	X�iDDi\4Ķ���v�)D�q"��
��j@4��șdH��*�-+%LIH��+Q*"��2��r�12�V�ÈI%�偗��#�e�K\��"4(�f.�\%+h�Nd�IZ�r�JP��hR�U�D��)hZD���K�\�4-"��fg�VH���B4c��.椅�r�K���
�v��jm�I��]ueϰL�tf��/��o]D���w�P��KH�#w]v=y|3& {+�����Bo�/�Un�����!!5�ݲ�ơ&�[����X��f�q���ha�{��H%�v����:d�Z:"�h#�}-��[L�v��7��SՂ�ޯ{�=���.�r�9�ך�^9�&�"�WT4��]n�B�6t�F]���7�����[�x�x����<��Ou[#���(ò�we��Q�U�j�9���{#~U~����ק9I.D��b{��/�;�m���;ۢ4��[�Ε!�[���wc�B�t
�Mʬ�v�[�#8���j�:�^7cB�WK�}�;���keν�d8қ�]Ut��/Yc�pэbe�j����0�6ΧM�4_
�Z�8��4^�US+��^ǹ\�y�7�H{
-8[ Z��Ǻ@���)4w�.�؆=K�xw�H�����v9z�y��>Z�0�A�2����j�_%7��C�=u�3#�)�P�=�ۨ:.�C��>~8���'�n�-�t��u�%�ŷ2�yE�H� �*T|��#'r��B�u�1["�R��#�r���g�h�ݾ��nȠ�'\�-?A3X�λ�6��U�\7B��S7.�hH���z��*���n���R�cf)�zA��C�����h{/kw�Vf�M�"峓߽�K��sgh�ھG�q�ӓ�gQS���_6�(�s��{F%:�&�Y�,�Fl�.��D��>��^�p��^��p�m`���bż[|hTz�����y�֭97����#x@�fw)z��u�Uyd�Y�ʂ�-{���Ύ���9w�EA��O�u��U�<ss+�;���QH�|͞�f��	�8{Q(��[՗J��c����*j=��^��[^m�C���[�rS�E>�����)�̊6�-+]3rq'���[mAMf��Wt�	�y]�34����]�+��n��jE���b�g���rx'�r��s�ʴ=6{�!�+-�l��Ԍ\������K�;s�q��v��`F��-�;r�z"ݫ�瓄)j�u�i����V%�9�_K=k��!�}[�kd�
8+�6omgc��aܻ֡�B�,S��9Xʨ��U�ƛ&bS���ٸ{b�fݱ!����t*C�%��m���q8.��볋Y�-���ɷ�Gp�շ:�z��O	�t!�9�\%�l���&QU�Y��S���N��ӻ��ۙU=`��V���0�r�xd�)�N�z�m^�	]�VoxE�{7��n*ҫu�ݕl�D����b4�Uv�:Q�k|{�����K�	���V���/G�x�P��vS�&�|<����^+8���3�za||�qs��8�T�n6���u�ˈ���q��-w�Q:�����xk��^�)�ˮ	/��%Oڛ�Y��88uN��ص�q���.�� �9��YQͼA�Smqxbm��,m�Q��Jo`���et
r��ۗ[�t
ꖠ���DUz"�v�=F���w\� ��NOQ�U�0�����vp!-Е�����޻KyЊ���@3OvD'�<��W��>�{j�ZQ�Z�W������w��.4�=O��9:���פ��و8ٜ��������8��=)��^�3wZ�z�X��R�N���&5�p���Uzn'���	�5��x�J��$���f�8b*=1�[鴞��.�z��|��&u��?��ɋK`�jP�m�^�u�Z%�A��_�IH�9�m=q���<gq!��J�m��*���g��������T�ЌUU_�D� [��"� �Ԓ� ɬ�pD]�&Xf���9�I[ǖʞU-r��1� J�Ѐ�G
يZC0��gy^\᭴�62��Cܛb�� 	� b3��5Fߴ��}�����9j|�[�H��a�eƨ����v~^�����'ތ�3��� O�k��g^�,}�P O�@�A ��$�F_�+�8Hp�����O;|�?���t,�h�@�8��c��~�z�C���&#@Kqh@]�d����%�5'��R�Ƶ	��]m�y��wF#Ҽ��]��Nd��A H՗��>���O���sA@F+�6Pv�DD)��Jm'\,Ҟ�;�ɦA����" 	�p/<�Mͷ����������\R������i�_��������_羑���L� �k.�b��=�����q��j+'���:�@� }���g2�]�"ɹl����=ZS4:���{�4 M�ac�ìb���Ɏ-�hD�$�t�!�� �Q� ���`�+��bWu������`X$"��\��A@�\�H��`ѡd#�b:F B5Y!Y6%W�?H4+����\bJ�;(3^��5�~�5mQݙɎX@�Q ��;x�~�w� H����Fǻ`!<φc�dk�f��o�w%9���X�p@P���˓ݔBz��!�6�>[�0
�P@:���m7F���%^~�pb��A ��_��Zǚy��dG���ؙ����w�u���Z$���T�
-#����Ͽ-Ak�Q��#�����լ7ӵ��  ���W Ç�i<j]1 ��$�f�M�kz��C��v^w�X*,��X^܃l	
� ���PwǓ��68p��T �w�Sj@\+�ï�F���\HB�S�t���� ��"E��4r����w$S�	
	�Xp