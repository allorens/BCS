BZh91AY&SY���"��_�`q����� ����b(                                            4P     ����B��� ( ,�h �6   `  
A@
� �((   	(     ����(�%R�  R� ���]�UTR�R��D�!%R�BI!QD�(
-}���z� ֔�$�R"PU�� |}h{��9�G*S��R����*���"<��{�O`�zމ��UD{�꼉n�"�ށO;: q�� �G�J(�{7����m��������lh�|���3l[���t87�pu���=	�{ ���D���s���� �ݏ@=���� 
 =��E;` �I
��$�D��ʔ� �|���u�� y�<�  ��h� -c������70�G>� ����!<@}�r���B�  ��}�� x�����ү��}It��l||�=� {���w� {�׾�Q� 7c��ްzx�� d�X � 
	>��� �
*�D�(�@��ā| 6���{�Ϙ> v=� �}�PO a���y��9�� ���������} � P  =��(}(�;��}�{� >Ǣ���<� �����+���Ϻ�R��!�������}����   }/m��JH �R�IE
RT��m���>@�p=���B}�}� ��Ap�s���z��9�>��zG��P���a� ` P )��E��  =� |��!��z���@��n������ v�;���� p   �y�Ҋ  މB�J��R*�
"��} ����� 	 tL�� ��:�C����$n� oyB��n� {��� PP�$�����`�g*zcxf= =��Ԁ�`G; �yEQ� r@7�@݀9��        S�J��e7�da1 aS�M%%U h�� � O�*�O�i�d���1�6J�aIRF�4� FL	OD�%*���	�0&`�0�"D#�JD�&����5CCM 6��|��~���n���ue�USA�n�jt�l��w3��EEt)w� ����T�Q_Ԫ
��'�4	��W��=?C��?�?>���E`*�I'� �������!�Qz�?��l�1E?c B��� 6�� %��(�6�F؈�[`�lPm�����bS[`�lm���Q�(��B�� [b�b���(��F�
��-��lEm��l@K`
[R�*F"��F�"�[`+lEb+lm��� �*F(�-�lm�-�A�(��V���*4�b[�6���-�`��-�`��-��#ؖĶ�m�lKdb[�6Ŷ�m�lcLm�L`��6Ķ�-�li��i�l[b����2ؑ�lK`�ضĶ-�#-�l�6Ķ%�m�l[cl#ضŶ-�m�[���%�m�l`[�6ŶF%�m�lb[�6��%�m�lb[��6Ŷ-�m�[��
e�)�lb[ض��6�0`�ضĶ�,`�ض���i��)�clb��6���c-�lb� �l��lb� �	lR�[��-�l`�
al
b[ؖĶ%�-�laLm�Lb[�Ķ�m�alKb[ض���-�lKa���-�l`���K`SؖĶ�-�lb[
alJb[�Ķ%�m�le0-�LKb[mb[�6Ķ%��[�6���-�lK`[0�l[`�ؖĶ�)���6Ķ%�-�lK`[��C�ؖ���-�lKb[mb�ؖ���-�l�m�l`[�Ķ�-�l�b[ؖĶ�-�lKalc����-�lKb[�l���-�lK`[��`[���%�-���Ķ1��-�lK`[�6�-�M��Ķ�-�lK`[�Ħ�J`[����-�le1�%0-�l`[�Ķ%�m�l#b[�6Ķ%�-�lK`[2����m��-�lK`�#ض��
SKb	���6�� �bl`"[b�[`�l m��T�6�R؃L�4�R؀�`lDm���T�
��R�� b�lPm����6��
�F��Rب�bl m���� 6�R؈FlPm����(6�Fؠ�K`l@-��*��R؀�`�lE-��T�"��b`�l@m����"��ت[K`lT-��%�T�(6��*[`	l m��-�$`lE-�%�� 6��*[Kb)l� ���
��؀�`l-���� �K`�l-������؊S-�0D�"��Rآ[K`)l m�%��[c [b�lm�%�D�(6�؊�
b[ `�l-��� 6�ؠ�K`��B؊S`lTm���E�-1A` S -�%O���Y�����p��ri�d7��0E�V��B��v�-;xL�׵����x-���p	�5��i���n<{:�rE�"�Ċ�xE�l뎊1V�z��1|1�g��ɧJ�C�oL�f����e��z�Q1:�p�	\��Pl�:e�	����W]��j��u�wb-��S���k\��Ń���}Ov����Z^����VE�>$�cM��ۛ����$s�ֳ������?��l�j�+P֗B ��;%i��������'9�Y�f���*H�bŪl�)��l���ywIí$�]�7f=qՄ���C���a/��m�餕9⣓�E4��-9�a�$�b�Z��.���o9r$�N�䜣˻���l7��%�x{�ۤ�	vG��o~z}.��_�[���t���OG�6U��g'�(�]R��)�t0�qǇn^�b�D��#x�w��7&Hɝ��e}y�e�=�T��Ėv��AܪU�4E�9��-]{`��FC�$<��D�����U%~x&��;!�t�C�-�f���w��s����q�3��A�������5l@�`�`.QСy{^���I ��ߤ$L�7���Ue��M�\0���7�d��k	+CJ�i�s��:q��Qh��h�vY';O.��&��,[�{&I�7�#��F
�X��R�.ʹ�l�+���vv�ȼͯ��U��ְT:���9tAP��b�"u�M�I�F0Г:��pɹ.���m�G[��;qiͷ3�0I�v=�9�AYq`1�ǃ��
햡@Na\���-Ǆj��^G7{^���#�	�|l�ByϤXwM�x�Z*���1R�h�xy��h/ܟ;"ܰ�:f�7�жLD�l���]=N�p��^��[1][�C��s�`p^� .�Q��u����T�.�o��%vb+�U狨�r�T��/�PԋH`��q& ���6bn��u^���9���gk��٧P�t�&�6:�r(#��u��r�=�(�u.;t�wH���(��R|��{@�Y�6ٓ��A��:�5V��-���\�sj�����=�''�;��f�[>;%��0��+�%��a�Ǜ{F���rg��G���6,
Oj��c9�h��=n���i�;Ga�8{
+^��S_&� �F\��$��2�2��|�*7yF�d��ku�"����	������u�;y������db�K����Y7���gf�V����Yͱ)�ҷ]oq,��o0�ƵwB�CGf=èS�)�ŔeKp�֌3�����Sx��ˈ�T�rg-�`�w-T��߬�9o8a� �,W�a�͓e�9��m�I���	@ԷUfڌ=��Wz�ټ��֋1ع��\�&&x���%����A�p}#��e�Ԉ���o	`1� ������H��4f�l<1k���2�Ʋ����Sq��1�]\(b�S�9��a�4�a��=r�p����8�$�m����b=�N�qn��s�p�4ҧ�d��f1��W��;�7zo

�� \I��Ik��ޘn�b��mۍ�N�# ֳ��'nS-o9�b��W�A���Ź�*�j=Ӡ�p{�<ʝ�V���I
�xY�n�u��D����O��W<mo�o�ו�Ň��o9�3�����L\{Qk�
t3� a�]��P>�쯐�<eN�U�]�&ƴ�쵖�Wh ҷ�a�o�i����Dbu��
a�&�[7;X>��X�㗧l�,��S�;u`h�suN����tMy1�9Mw��pD髎
� �;$Y��%77_bỤ�4%��X�P�����X�����O]�vs���ݻ��e��<I$��w��렻�x��:i��}��-K����;AI4���r=�o0(�ٳ;��Ƿ���l�sh�	˼��f�$}��/u���fUWo*'2x�m�d�]{�A�s��O&����Ӈ��|ۀ\�jˀ�Y��]��Ι�w������^�	�
л�-0��p{5��s�K�c��H��%j��:���P��4nno>j�޽3�JFN8� ~�P�1����3��{�*���{p���r�u��r��/��GJ'�Z���p�7eY�a�:������bɋ������j�^���Eݸ�u�ٳ��s���/#��'P�����d�'"�l4J�I���xd�y:�㳌���e���O�]�R�bW�u�a`����,Kf��I�[F|J��i�&�_^��yȓú� �s����9bp��,���!��"hTh�����\��/^�eS�m&u٧5�.;ڡk�{y�d��n�C��&�|x��R�]�H�؎j�i�䓻v挸�ɺI��N&�����.�+�s����NovK7���[np3Ҡ�c��C�u^`$s�4v�9���|�̫2�:���H5)��*ۂb�K]�m,�@e44Q;��t���9��M����7�@`]DpѨ+iSB�&���vi{��IpZ�_w(�z���՝��$��;`���=-`Ue�.�e$b�<��4p�n,���]ڞ��-��v��r�&��x���+�c������ԭ���s���$��E���s=�ҽW�^��_k�wk�'T�5��=���Ǥ����P�1����9��NZ_n)�CU�:2|X�l!�榰a�G+��\mM��=�;�l�\؇
0c�`r,O�*�m;3�fkS\I��$�c]�W0�aH�p��]��]Yj�����ќd�}���4��"՚O ��Ǡ#��ن�LGV�2���%X(�;\L�g��귙��o�I���.*0��s]8��v�f���X�9�wXy�v����M��⥻t�:�T��D�캜z��wf2M�e�j�r]0�f(��s��^�=쫀���Jo��m��u^X�Q�nwf�ʈrڔTf����'�'�{(�w:�H��f��sxqꪼ����[�mt�:U�˹b�d�{�>C�8�����ǁ�vk{�I��u�U�����ʮJ���#&4�KtlG,Yc	`�PNsv��a|�	���Q�'��ɦ2�ܲ�Yf.lS������k��2��S�ߵ܀�h�j�3{w.�껁�B��Nk��ȅ5l1+�p�΂�h+��7�\p�}]dwol�\-���oe�jiW���x�t�����$��c��Կ��!I�C��]��+5J�Θ;u����3��t��ckF��K�/ӽ�^^�G��g8����n�[�/V��u��,v�<��P2�6�}��T5^:Dq���V-��@�jȾ�D��]f�&]tl��!�J�C5t{,3^)�f�x�݇��������܍�r���ւ�}�c�x�i��p��:�a�`�Э㭑��`�\�r�,͖N��\ܷ��
��q��.�v� ��c-9�]�^��9c��y\��[{:�x�ː�p�`ǹ�c�������	�܉�q��Ȫ喳ʾ�hfEy�8�����t�6:;:���8�G)��E���c3R�vd�9���7؃���k=��,j	H��㷄˕��ŝd�OR�s�h��5�3OD]��]n�f�/+��zp��ç�nUP�\��V>���[�IK�E��su���\��4����woLx�odA�j����/q�E���6l��j�ɚ77l[�>������#;�t�:Ny{{8&�j�!�^\�9�]��B��r�+z�K�����=t��R%�Ev�r'���*�.;�_>�9�x�n 2� ����;�G���@��j���F�������bɓ5�5*��q��L|l��{v�s:�'s�%�h�M�lp̓r88Gr�MŧA�f�l-�3J&�����{z�ܦ�Υ5�o^L=�4�s��W<�z^�9��ksu��'�Kb� �pW�1U��h���棬h��;��e�������t7�c�j\�q��J�q�V�^;כ\�F�2�R:E���x��|���ǂ�Q�B#o�<�vMY��9Q�N���u�d��lN&�]Ǆ�;C���r6q��8�r����8冻fw1H
b��w�:J�Z��x�0`�E�n�v�-���/�p��b�e2\דCٺe;�mۈQn�G.ç��e�W��o-����p:[����ڲ����
/oF�z�{'���/|՗^����ݼUF�e����O�m'I�5F���(ܹ��}Irc���w��2u[L{���[�Z^�4���P;�dF�ξ�G�(��[�5Hty�����cӌ�3lG��QXJ�h�ȇ:MX^hAr��a/e��8..�L��ú���Dg���m�g.�hS��N��٣��n�7��5t�ҧ��������:A4}����uc�&L',ݕ�N:�9���S���<&�k\[�Wp�������9��ak(4��r�.0�z7B3���3�"�{F�<V[�l����.%����&n­;� :����/h�Q�ꩾI 㳕}�T�
[�_kl;�_h��[�5�ql��e!��m�3�����[�n�^s�u�9�̳�GOJ���#y���V;{��-V�/uV Ӿ�{��S5�����"ݷQ�wrNݻ�+���3�g-�U|�xTQ�<����f����5���S��붬�nf�C�A��#Ż��v�STg�l�ZY���o�G�=�9E�]���z̡�d|�m�c� ���Y�3��+7x�դ�m�l�w4a3	�7P�n�fEy�7����ϧ�s6��\�V���v(CNWyp�B�ɐ��7r�n	k�@hmle�p�sJT�F=B�4^=EU��w-x�8�`�$wV���:��v���Q��x�s�N��b���9�^����Q�o]֥��U��C.Ѽ�LLئ۷X�k� �p]>�C���t�G8ȶ�������[8�*�
�!X/܏Ξ�@��m~Y��8e	���20n���sN��"�.������|7���v9Nf��6"�m�!NOD7۴٧�ŀh���B��p>��)�}�c�Z��C�7x%h�嘱��d�b���ʒ��=�x����޻w�acW�w��U��F����FC��9K~�m\��S�3^,�94(Z5!ӆ�����U��� S��*5�D	�뽼�w!�D&�#!$�|5�>�B�@ ف|&��	��3	}�
���"�1�C�|
�@8�t���&T����T���g#AB[��T-.�K��+)^<za�ʥx��Y��f�p\CAYˉc�l��Rn]�k<��n'rv-A�r��E��!M���;/!�ɡ�+~���:� |;�s�ь�4L[�͌��1˯q8���D�1-�[{a�ז]�HX�ί�oagy�7sԱ�P�n"�ն-
j��E��Z��u�'"s�n���O�ҩ��3���3uu����=��ͨnj��E�vл㮱�=1vn��]�\w�փ�)0�su*�*\��76]�υ!+�mqy�4���8.GoY�!�K >���]>�ҟ!V�L�#O�f�[�7T��˹@C���ƳI[�w��_v��"�I�1����˖)`�ά�w&�����kٍN��#D�M�'`�6k��ݢ��މv���͛�5�Tϫ�@�N�7��d$z7�k��
p�1���>\#����nC5N� �h��s�l#[Ȇl�O'��80�׽c��0�a' c��S�BZԐ�Q��_���wn�t�Z"���v҉-�:������N.#\]��z�PH����<���H)mZ̆M�M�$g�S�L�ɼ�xoR݌5�����É����!gS`e)8�{soK!!�mJU�H��(�x��Z?{|=sX�t�_|�bs�0���❠���|3�K=3���]��}�7���Fm/������H�>�ӭm��A#j��jD>5�*n�$�K4��Ƣyo��|i����Gޗ�y�qыw7w��0ݨ?!����i=�ĚJT3�)�y���5�T��a��N��^������"�xY�E��c���mӛ����w��
ΓF��G���t��9�����S~潕�/g����9��	��xbҜលFUV��	� �3O��,�0���~<#��}ôc.�e>:�{ۏ�{����
<�I�"����a���ͪ��쯋��XL8{9dRo�}y�S�-8�^��׆���ݼ}6{=7~-���N����x�ccH��
x������[�P�d�^v�ֳu]~{&0�f�2j���y�#�f���r���Fg�|;�;{�}21
\{#��O_������/����h;�M_A�u��}nޜ������x_|7�Z٭i|�Skƽ�(�No{�j�Q�r�b�z,$���	���xv�
���=� �}{<��4`J9w���Țrq��e7w6��(�OCдҊ�>��s���'�"@y�se]��G���`������y'ꁼ�j���S���� ��ӈcP� �e]o2��(�x!`,�K*zdW�ǰ-��y�M��N2�#�?���;�/�3��y}C�fʘs&���o�sl��>�<��c4j!7���������8Y�U��l:�f�P1 3�����^G��׽r>��������|�+�]X#���H�� ,� ��-DQ�E	 $@* P$j"�U�*) (*�J�! �@�U�VF���	$	�$@AI�)P$BD
�5AREU	 @��IF@	RE$ABD�@ U$D�Q	I$DBDAV@	�E$@�	@�YA�* �PT���� (� !PFD�RD �AY�Q$ B�"�D�H(5  �VAdQD@�ET�P�**�PD@�VD@d��U�K���UM,޼/��-<�M1��W���3���.��g4���aJpӚ���������mX���a?�����Jb �� �m����&i�Y���	n��݉
��}}9�l�%��j^YĮ�ͻ���'�@�m5-���)=O6��::�����&O��</�?"e�xwl�̨2���<s-O ����c�Jѡ�-Lf����~�Y�1/��,�<.���|�(ߗ��$ϵ�/a��.�%v0�%��x}_Ɨ~�[�$7���|�N&�I͈`XJ�~ePY�b�B�u��ر���~8���8��[�7�O GI?�	i�͛�@~)��IoB����S6h�R_��a�E&`��ڛI�k6|)8�~m��@Qi��'u�!�
�8��0�sP�8�'2�
<W�4>Lc��9
Ð�{�����Ji��7��5���c��E���4���+BI Qt�g�>yV+|�+F���0�KA1�@�X�a���O�-'��u��e��Tj�u�/���@��?���QTD3ߐ�.lS�~��G�g�����~�������G�f
0���A4�8_����� ����⦍�6��u������#!�׷��~�1���|�� �7�t�w/�A�/�T;��)+�9��v0���>�xi�ݻ�[��=+�k�y����l������ �BA6�>V�B�j����i��]N����g���L���3�J��^��㬙������ߎ+�9N���=8c���~�����잃\�1���p�;r�L�ۦc���G	���h���_O4q=tp���
��D{[ɼ��yυ�0yog���R0:uKɅ�5^�61�Q��0k:vgG�^����x4[2�ݚ�ɠZ���jY�ڂ�X��ނs�K�I�rk�=�ln9g�}W�)u�H�	�ďfXǶwV�ֱ���"��\����<�����d�`��3�V�S���s�}h��x��cR=�<�'���r�G�>D ���o�9ګ��������Ur��*����l���k���`�w����G�XW�g`=����N�#<%�7'gy���'ĻY��;���^#��a��<� -��m��A�m�A�l��@���3)���^�V��Fl�s����!5R��Q
�\<�d�d�G�/�=�O�������8�q�q�c�8�8��q�m���ݽ�����q�qێ1�q�{q�nݺt��8�8�q��q�qێ8�q��q�q�8ӎ8�8���8�8�=��q�qǷ�c�8�n1�q�q��q�q�n8㎜q�t�8�q��q�q��z�:���Yz���g�5#�=�iڹ����{c���)��[7�PM�^���<Dk��>{�>ΏD��԰r��O���[`����]�^�v�mk͍��H�i����7w�}gCӒWϟs��~~[g�0=�H�1��G�&<V=��`~����/e7}�Z�!ba=�<%�{��Jʭ�,��yj���]���L�L�eP��*ab��su2��b19d�x+�ca��ѣ�x�W��r+ޔg+}����v	���agK���d�Ϫ^^9���`���o�l��{���r�V��ǫ�<��wa�y�!��t�┬���:����<�:�v�� T�i�w��"�iv�Z��{5��T����6�f�X繵$�#̿-������C:�{�Ǆ�D� oH$cه�i�9�)��ܖ�=<��fu�,A�z��ǻ���I��� ݰ
b�ۋ:3��5�a9��lC��������EAIĚi�7��sW.��3&���x��9�;@��3��{�9hk5�XK32q��O�+K;�yd󹲯f���n�z���1���n��d��/��ÔB�n�ptY�b�R�{�8X�}�o��Om.[ݶ����\�}kP�r���㧶:t���q�8�8��q�n8�8�=��q�{x�������ێ<q�q�8��8�=;v�ۧn8�q�qǷq�q��c�8�8��m�q�N8�;q�m�q�8�q�q��q�m�q�8�q�q��q�q�{q�8�8�N8ӎ8�8��g�z'1R�Cl����	�,�)NU���ݾ�?�d���ų2�#zn�qIG���}�Xp<�V{�;tgi���jz��䅞��+P�g5����μ��y�\;�$�B���NuO�q<fXlߊ�O��M.zW��/u��p_l,��)�Ut��� ~���%O�(���;�:���nw��RQ��w����_���.�ny�8��}�w��f}�z�b��>�7�������o}��,ؙ^�g�^�#W���`����_zzz���'����	(c�{�F+9�]�]����S�m�%;4����͠+�勆m�C��<��3�RLl{^]��m�d	;�����}��G}9��>Y����مX3���������?w9��453��;����f�G��foO>���z`�em���>w�����g̛�$c��ko����7��:�|]Q���7�s�#���8��6L�ϣ3b�{�rۛ�m��{�gc�a�>A�R������~���)��-�^�ǹ�d�]��2ׯ����J0���*:"����mʁ���#پ�ӯ�~�X�n XT?v��r6���Ɋ{���C���=�����z�����еq������L�g�Z���m���`�k�X��罞��*�)S������]�$���:�i���n=���zq8�8��q�q��q�q�1�qǷ���������q��8�8�q�n�v���N8�:q�qێ8Ӄ�8�=88�8�8ノ8�8�ӎ4�8��q�8�8�q�N8�8�q�N8�:q�qێ8ӎ8�8��q�q�{pq�q�=��_��,�FpkH���f{�B�XX[�҂Z(���h\N�+�j�=�Kh:�OM�x<�Obk�ȹ�sǊf��>�Iψ峢5�� ��{��d�Ґ���� Y�>��LP3�}a7`f�n��}�����f�}:�e���Q���a����\��V�z�G� �Ո|s��x�}{�G�'x�0���糕��{ݓ-|�����q��oe:{�uS��H��2���d3�4e{V�mR�,5���9�pc^�s������J1�h\�m��d��3ޫn�5��3^��X�r�S��o<�qZ��P������N-D��ok�[`���X~^��4��%ܷW��\���L���z������^�(��z��כ�l�̾��{mL���z1��]�s�>��s5HB;�}�f�M�5N>�6��9����b0�l9P^^�b�Ȕ����l�����YHף.'��l�=�������`�gC�6p[�Q����y<����w%�v TC�U�������E:t���&)�vj�8#��6Z gE�,��}�׻lM���/�93o+GG�����6',<��f��D�]4L2�����+p�+#�.����GV�7eҹ�kQ/�>�|%����}]}�znFw�gm�z���u�z~�4�(�a�{��{ҬLg9Κ>ϵp�vwj]��X+��f�C�q�ڰ���ٙ�.9盫��yj�z�O�����%U��w���fY��YjC��3�#1�F�!�G��[��sq����� �U�ʚYB��Y�Un��1��������}�w����j�}d��<�/�fO��DK��g�^G��yn��q�F(c.L���oG�u�߮�߳1XT�Z.{qB��@{7��: ����}�;�
�h�� 4�`�i�0=E����*��'-� h{(�O���S�s�P��gU:N$e\/�l#�h���"bx���7π�\ɳl9�6z��L��\(��ٗ��)Y.�{�;=�#�{p�?-۶!;t���˙���� �ۑ�m��>����nM�̔����\ruo.Y��	�x��s�ӧ�͏�;T�Ԑ�7$�ȁ0��)� @�~Kj��i�>���{�z�<�U�y�O�t�9Wٖ���ǯ��x����rV�.Ss�i��yW��x��G�ȉ"\��@e$�RW��Q��|��'r�;����OI����|�{��g�π���fVȊN�8<�F3��?u���:o�����X嗀�k���{�~���ԥ@s<�S��<��aZ��DJxˣ7��rE}�����cg������s���*5���T3�y�f�|�U��؆�!({}�}��g��~��/�l��hZ���� ӀV�k�����X��;x|�`���m'����\�2x�pɁ���
��I���s�H�����x�Oo,�;y���[}�����(��>C=���.	�xQ�������*vI9�:|��t󮞤����9�!g,�pyn�>���-��r��j<�E�OX��u�[V�W�o�t�7��]��_yg��n���*����p�}��{��zh����ܖh�{ݺ֋τٓ=�3]�r�n�3Kg˚)f��}|��&�f�˰xN��O"��'� x��#���t,����3V�Q�;s[�5�O7�9ʹ}�{�X����7tW�=|��w���S��t���>�I�y���U��K� ���'�8Q�?�M�� ��>*��}f��O�p���!��;^f��ܭ+_�q����� ������ΤǾ?b��Ё�J�A�����`�~�|h�S�6�y�#�\z{ǆq6}���ʘ����Ӡ̨�.2s,�o���� ���^��Vf�l���h��F���}�}�m�Uc�ȏW��F}���p:��G=���ރ˱�x���,X�t�sv�r�E�㣷</bD�yB�^���ڳp�4Q��-��⤣��Q�����A�9��T陧���l�y,���ÉIx�|b��폃�EY�zg��p��̗�}�������*�.X�ב�&v�U1�����o��F=�^Jvz�׀��<�\�=��>`��/�z����D�4�B�c�$�&���CS^c�7zn���u��?s8�٘���sŧ��tH4ެC�^F;�Y�Ez�GEֹ�퓐��;�@�i��L�5�׽N9�,�����۳���R��D��tj���O��K=�ˣڻ^Kf��W�ݹ�>�[�e��8�Z��2q7��޹�J���n���筂pЈi�q��C���`��ux���K�����C��F�B�����_j��f�v�2��|{;�>w�mx󖐱�� ��ʨe���*���Z��𛞋_�J�r��g���_z{�D�~��mP!#��`���4,;�z���l��yݭ\ܚ��:9�{�:.}�S=�h�Pt��=�8vw�z4/s�z`b5�嚎�V�p7�X'����n�2�]~��yyHY���1ӊ��re���7�w}�1��gK�t�!�^G���.֯,��O>���貀|ﲚy{*��5?�|w,��"y�^yᮄxG����݋����>�~K�"�aő.k���)�����Gڶ;��b��O�?��̶,�w�ȓz��҇Ȅ�7��fh����{�x�<0����=�-kgg�$�73q�����{��"�$<��1�2o�Qh��g�+��{����e���Z��MB���7d(j�n�Of*��(R������͔�E��u1�o{ކ;�u��u��^�/��9�bӇ}�kc|�O�Y�Q��C����{�����g�ʣ�Ҙ�?& �Q}o�V�^��3�D�o3�3�ӿT�,ocѾ��8���s�_{ⳁ����/,��w�������%�G�p��&�P
�׸�'x7�fթo����ls��������pj^��Y�msV=�`�Ͼ�^�ğ�S)��_: �����1዇�����֟dU�]%�Oђ��v!V���d�[���^�]:IލO�3�պ�z_��ER��Ȉ�%�=�J�ꭆ��&�l`��kˤNBJ�ɼdDH���]�.7;y@�1}�L�`��������_ס+�}�U>����/����`�af��m��q�i�!��8��X3��۞T�4n��
��}���z�o�OO���5I�o���(����~���ɋN�o����;�sr�:^�����G�X��D�l�G�C�3�3s&s�s��Yeov�F�x�.��O�����e�����P/��焷e�e��U���[��o#^d�K�e��N�]�7�|e�<=(����������������	 �1�;��\M$�kޞ<l-y⽷w�;��E�<�k{�n��I��x�s���E����G�9L��ط�x^�g����y�@ٵl7�7&Hƻˑ�ݳ�9�w���Z���O�</�%�ܓG���ǣx���9ĵI�W���;��C�z:�~�A��(�#W��e��,�|=�!(��_F<�j�ܠb^���{���_=w{,�^�n\~Իpt���e��;:��{�3�p�?1��ޞ���Ƽ�ސ���/*��e�+�W���-��y]��{q�����{=��)����t�����t��轕�q���mc�>�z�%;��f�y��^���eEv��od��&�e��_�����&�I] �B{#���2��'�Hza�޺ٛ�+�f����9�`��Qs��v �p�Jp�
Ǧ, �o���3�*��v��=�Q\d���a�]f�ڀ�=ǽ2z�Y�^�,����������7A�r��[^�fԥ�,�r�sx�n߀֬���Ys^�~|zu�-��0�%�	�����j���
ɼ�2.~��{��;�b^�����H�t���Ov�C��<�l��yzN^�cž�����M
��xW�>�E`���_Lo��6Z������7��c>���d�J���&�\絼� �����9`�R��˫��='og�O5�P��s� ����;n�s�%�?ݯl�M�5g�<�w�ᗐB�*���n�K�+��f��w���<������^];�7#��DZԧ�qau�����O������u��~@ٻ��w���}�Z��q�.�/PqN�|�n�{m3|�x#��}��T<>���&�ݷ�.k=����йչH�*�v��b`�(.!���r =/�St�P �g�/vO��p���q�1�/U^�d�A>&r/���o����$��燸�O�� �؞�}�go���=^o/m���ۜu������_l��9�i*�8�W&�f���h�6��W��1�m�^�*��6�F}�6��xW�ݘz�A睾bl�r]�"����wg����>�9���s�۪zT+�q�k�v[f�xx��W��η�� ��m�^���$�p��wI�^ƺh�m<�������|�ޡ%��{�i�0p���q�t�R?eg�����a8��|k����z��f�5��}�*��Sl���ū��{�n1�g�����p���뫕U��{�[�u���������P����~�_�ҿQE�O�~�D�����Zo����MroX0��m�6���ȿ����h$�Y���N�^�	,���A��?9����e�7��umgJvlx6���g'n7S�6�xg���7e�@�q\u�1V��- �))�l�`���!����2[�`SQ!+�u�b�Τ�U�u<����$�m#6ҕY�4��2�	��4=O`gn8�U�z�8;zl�jՌ�����!��]q���Smc̈́W�۞��v,�:6·�]cy宴V�m��,�/f4���Es�Z���!�;=s�O�v��V�\�GR���`�v���M�o��m�Vz]����g8���l>}&L/7Mqt1n۹{'��I8d��ۭ1R�hbm.��3��XWLk��s��3��C7:�c�<KcJT��->-�tJJ�V�$lr�a"h5+	�zR[,{fYz��ffi�؀��"^���OVB����)�X뗝�ڰ��宓.���ƠK����V�:HKu��]���/��yf�G�٬a-a���Ke� �)�GKjn(!i�3g.&I/V�֐�Ɗ�����f�W[�8���^Tx������ӣ��d�4�� ��.gDe��;\l5��z�nɮ#=��=z�yCkF�W��c"h:-��c�Ț�v&�^֧E.14 5�3��1���x�bI�,1�$�O<���x��w=�L��%f���[�Xq�����4J�	��l��i �vy�h���lgG;�(B�\L&F�,��u�FT���ފԛ#�7�fHÒ��c\�z����hxK��-����$&�f��c2�MٷoK�{8��V��ܴQa���at$��jGcH(�0���Ϟq��9�\�ru&�L��{uf�k��:�䍆�@� &��]h�:�ֹ�м�Ap��A�:��tb�KM.�aĲ�Ktc�s&�n��tη���ԒT�6/�t��{p�*��j��u��W�!`$�e�Xa���N%���L�Yt��K!P.�	��M.�"&1���t)���ɷ���㋱�x����|N��w4ڻ�&�������g�`����Yi�bC$J*��!uR:��K��T�Gn;K�����v�u���66�!����`�ť8�1]�����tl��ٲP�j�6�A\Wi������<����j�\	V;�9/0��,�0&��a�޸��r�C�xɇ����T��뜴�e��Ap���#v��#���Z���w��_`@���k���(y6�ՎǶ#�g�UZ��&�a6�@c�poZ�n��!>�N)���}��q�\4Ί݌�*c���W!���1���
[bs�[c9�����Z=q�Y�C�q8�K�q�A�c���Z���]uκ5���J�r��c.R���ѕ��ά��狞�0mQ�M�2�
����VYl���b -�Ic����Q'�ƺ��rV�����qI�L��sՎj���FĎ�P��I)�C�GI��h�oU�^H���yW�S�.�6�|n��Lݢ�:γ�ڟ]�"i�p�645�Ε�-�6v�;x�m%�40u�����㮶��69��e���[�7`�۵R�v*���W`�]n��p�v!��s�K��϶�qC�n�E'q���
�����g�qq����=e�n����mM%���pj:ڋ�u�<��E/���v,N.[m,M)��QRX�2�MN9��b��㵹b�08S�]�9]�g�����#����FӮ��a�b�*H�q�`��ZksƝ�Uq�^y���Fa�\{u�1�В�(�,*e��W2�s������ �j87b6-���z�X���=��[n�n�n�9��Aщ�s�u>zqm�I� ���Xɲ�v��0��5V.0^fW
��L4f˻KBl�f[f[����J�F���j�n�k�p[ Z�\�@���� ��JkViR�(�錹�o].�2�V4gL 'Q�;f�N�],�66���H���I#�DF�TT�$��a.���e��  �JW�U��Ҭ�e�'�������ȕ�s���÷�����{v�&Ɏ���=L���0�gZH�k�
�;m�g��lVU���BW�-*�儻�R�) ����E�;-��C�bz��g���u���jLY\�,�%�����x�`�=V;FKڑ�`����\3-� �>x#���v�nȉ�$Z2���Wd̍�vڎ��3��r��3v��i�GZ������;X�V��Lunq��=�\c�qN��ACg\c-�jhլp0��Y��
䉘6��2h��񌕛��z'T�"�����zy�<oP��:1��1����Wø]�"鉆���u32��)m��pԜ<V{g�n��n,j+*�4UvF���n�]rgǒ�a���ր�e�Z��\+�=Ѐs78�ڴ(�$���\�(�`Ybd��xN�R�x��m.7llvk]4��9.�+�e܉4(�t��Ż%� C�2`Mti)�&.;�S32��c������`��𝮯C�|��O[���+gH��e��G�L46�P�R��k�!VnE�3�p�[Kvܰ���!��r{0�Y����0\�+u\w\Mu�f
Ĥw!i.-�5��^:QL׫�nǎ�nnc�Gu����B�VZ͉JC]C��wl�F;&9��GYaMۀ��^�9�9�Јہ̻4�1%�Rn�i�ڼ���]f-N:��U���v�h��p���2\��Z�w\�mn�OoF�ᖄ���CZĨ���$��C�^P�;C�:�u֠���-�.h�gAk�g���I��.-@��x.�U�$��v��I�G���7\�H��'X6R��A�a�#�R�I����k��"A�k;Z�۸�m�<bh�l"-��c[���.��=�㮉�����\&��:����t��Zq��3�yr�K]ua�>1Z�q���h�[[[���!��V���[
�&%m��&`A���%�^�;�
��4�8hn�
ۓsh�^p��0!�-!l&���!�ڱ����Li3.,�f�FfmEFSH<[ �5��,ŷ��pW:[�B�T�d��=�sO)���0�:�ش�]���I\.�a{F�F��6�Mi&�Wi���N&&;ZWi�.0.�@�e��Y��HF���E(�4�fz��qG9�J�6v�����w=���.�>����vQŊ��Js���-ܔ�P���Xgr
�b[�f�:��/B�S��9=ua+`T�$:���M��ҭ��c#\c[��z6%�2�4Fc��� �[���)5�]t���bɳ� �-��Qc�����{8�є��"ڸ�h�hL�r[�_/1�]B�Ξ:msxNkjv�('Avu�'�뮜l<\���7���n�۰r��e��i�g�@��Wm2�;#sd�	E��nv��M��bn�W6�gL�=��uly�N/u�;T+�"g�S�8a�t�g�7mԗn�<pY�h8�� �`��E�Tc*i����6ו��W���9(�m‭��y�v�db��lM0Eb۬h�Y�L��ݝ�8�6FQ���^�.(1)M*c9�s��p�ӜT`��P��6/p��� l�[����bR�l�س	��q��8�(DR�]n�W:f]Dԩ.�Ism�Fm"��3�h�����R��HJ.{\q�\q��k�4�jN�:������+��fDAH��*��,qA.{Z.S\�5f�}��ڛ�vk{OO�ܶn���@�d����mZ�7Q��^ӳ��g[�ۆ�k�b��ƌ��w��N��!8&�ܻ���4���D��]cm��4�!D����1�ц�P�[��Ε	aIE%��u�m˭���,�U�um����k���W��7��r��R\�%�r,%f�A���ī4�d��'s �9�C�v���fz��<r�u��CA�axH�Z��㡫�,�w�o��{��R8ǑVN�O�ơ�pq]�����ˊ�b�:�����'�䣒����P��hB]�,��1�kG��M;n��4A�Ѭc)�����e��kq�=��S���,I� .�]�V�ř+W\�gm�[�pF]]Z��h=Gc��	�����v�b�৑[��7lzf��eV�ēl<n��H']�&y�Qۍ{V6:4�97�e,�5�.oj�����G*�U�Ӳm��Mu�WD0n�i�\�dn��sZkc/Zӫ:KĻmt�4Iۜ5g�mu�u=AW�q\�غ4sy�����C����$�.v���ݹ�.R��{O��$o9��k��ԙ���`Xyqۘ<�������Ұ��M�A��������/I�q���L�t\��oL�@�ڸ��A5�����������@VR+�eȲ��j��i�ҧ]]4�~y�C��~>Mi�IVVx���Wm2�j<���[1�iM�L���".�9a0Tq�X���Bɶ�PrAs ��)$�r�� �6G��q���J���\{{c������n�:t飒�X��R���I�V�XLʘGqQAe�\�"�@�ĩKuWQ&N8�4<xǏOn;t�ӧG9\V ��Ȯ*X��Uyl�9	Y0G�Lr̄
+.W8#��aL�	!ΰ�/���i�ޘ�㏎�:t�\��s��`��q�Er�".K��aq�\+��Q������q���v�J7�grCA#��fde�$���tl!�8�!;���:H��H�S� ����(��L�AΦfkUG S"ff�kp@�̒���[o(W0̘�"�!v��n�j�e��-*�Y$�M^���s�7e�Ms�n�X�%`dH�@���l��St��Ŝ��	���(9�,͛LY �i!pDLX��"�Ե�3%nK����U˯� 1�۰
�����/aq�1s�8���+ۘh���V+�+��-��[N��1�ы��$��c��
L����+zY`+IU�㣚m9�ݑ.�qoBVX#z<<:��8� �� �R$:5㮪(��B!$�	�F[H�$�^��&�HrVm��H�u�wtswK��U���%��f1���P��ɲe��L\q\D�"K*-�\5#��^hz��
<ZоL�g\���1d�r%��!�5"�8@��d{��X��R>	��37��u�dRJ�w��U���l�o=L�v8��i��:i�H2�M�����^8m��t&��2-��Y��VWS[����fa�tf���8�e(��([[�'rTCHBP�Z+nH�z6!!������s�a�v��x4�X}���u�eew��Z�D�u��J�p*C15��ҷO'��n�cq�� �Xĺ6�8pD��k���ZM�}���ә�ݹ܆9�Z��z�)�٤ ��4$;B͛�b%�MV��e����,3��M�rm۪0{Wλ\p�P�jY����Lņ���Ze ��qE�ֈ���`t`;���أ<�[m�)w��X�fF�Ic���+O]�R��Pg�������Z.ehpH�@.eq@�B;!4��%*��5��u���:�C�f�\�����0c�MS�x��i��^M�R73ɂ���]���iG![`��B�T���2�L�wcB F�kD�p	�m,�%@֥v1H!Cg��@_��5��W���;�����:�x��!��k���4�BSM��M�SA��&��NM�|��'e8[��\�I�㨡�wi壌�z�S�m�T�@��v�#��g���2�:����/K\�s��{S!3��u֘�ˠB� V�-'����+&x��]���ƅ�+���P�Z����;5�bY�x&�L$jB��N��/�
�[f�����;�����;7�Sb��������v����pnf��]�%�-��;,x)aRc5�ڙ!Ɋ�`�'K��1)��4Jԃ+���ƹ�Ҝ�g�r;l&���4qK���rl��\v��fħEW.���]!��^�fݜ�g%�m	�\s�V72�F�c��Y���L [��N��Ϟyі��`�0�,���z�e�h�E��R��*BB0��,	X+N��ee�դ 0�ƬiAW���[
[Q`ŋޭi/^����l-��4"JpR�ZR���؁��$�V6��F�$���^-9�Y+%ak��VZ#�Z��J4�,x傷�KeKKT-T�%�篋~�mv�k?�n���z⍣�;�8���ෟŪ�͔*�@����A	}�����I:vu�᪁�Q5�q~.%��崂A$��j �|H�l� �_q�M1�J_w~�|9�/���bE��Hp;���:̀��o�n�惩��vp*����pT�߾�y�ys��ZMݶ,(k;m>�)�Ds�n�`��e���I��][��F��[�ɲ���t/6�D� ����*��ԧ���jf�v/<A�z�x����֕������b�~0�vK�.����IG�!&[� h!	[n���2%�Kɛۧp�d�-vv�iSx�c�]^Cw�"
�g�g���.��H�k� ����^)��f
ɋ�������Fh�NE'ʳ<���~G�J^�\�<�����������Y�ͨ��O�Oe\����%��^���2�v�u� y�1Ƕ��Tx��y���y�@�c�HؘzqZ]$]úE�H�O+G�K/�l�|}��Y�����$M�n���6���P�"A,��,��TT8�f���P�/���?�>u� o��ϲ��w�0{���"m �h;�My /ʶ]�1uc �侾�U���|k5��7_"����a2`������r%Y:Þ���zy�����khe݀��푠r]�S[a:==|�_��m7>�g����G��Y��/�WR.ciF���z�J_��ɛ'�=q뵖-��k<��ן�fw�v���YM���5����8��$6E͙�U�8ē�bl9)��v��+�$l�L���7�ɇ�}6n��(� ��^��OEj;ve�3�V���-c��)Ӵ<�ˆuP�֏�?i�^˄*\�=�F"�M���3͠��F?��{d�}�̐Ba�P
��Ej���	�A�^^Zs���@�d�/$	��+Se���i�,�qZ.}M+yKЁ�Q�轝�4ѧ�؃�@e���A��q���4�7-��Y�8��A �2��'o$�䋥�\d(���7�:��k���I��K�+1FVg��^��r��X^��B�"of?��Y�TRC��7/��MO��E�Pl��!��v<̕l�l+��d�j2bP�3��b �F�f�7XCE���gt��kFl�7���V�>$�,�	
[+a�J� �Q�(������S��2�&�)��ĝŠ1�Փ �[Q@'!��I����(�m`pk�H��4��**4�w�m�w�Վ�L���=s���w�OF6N���}8�%զ�8��ɛ�-aV�n$�߰{�I����/��H ��������f�I���Z��>��yظ{��}��{ �����6�O��[i�ȁ1��|q$B�^G��{/�-��P/4v����qM5*�.6e���LM5�f�w\�$<����[v�R���ɼf�1 ��V�ro�b��Y��~���`���~��vyCM��6���_�0`ԟh)^m�8�u�f ?E���#�]?�L��F�QOQ�<��3�ea��;o�x���W�M�>B�T4�L77�O6(&-7�z@D%����o�_��ہ{�[2�����|���'�IV�9$����i�C�V{�sÀڿi�/�:��,&�-�[�	#j�I����5d�t٪	,��-��y�'sj"�T��di�Ch�ͶeFAȳ&ĈP՞i�Y��\ ���M�up��6��18�N��ģ�~+�}�ur_3p���!�盨���y�;wiu-�wL�n����k)vQc��d�X�,c�+�V�9���f�z�r��K���@��N�b�r�/b�^�s�ط6�]�
xJո�Y���9�j�1f�8AN�u��P�������^�:iK�#�7)�X�p͙n�J�!��W�VST���4!�͸�,��n ��l6�@MwM����Qök�b���tnΣ���ѹl�ܴ��][��|�h��f�A�ݑg�b�<�-�H��x*ܽ)�b���l
��A$m�y��{q�L �#�㠩dD�d���ml�O�-�Ăq؈o��.*uXˁ���� �,0�̟ɝ��*�c��:ɝ|<�n��׿s�Ǭ��}Vv7�cy�,�%����#ga�F@4�1c���;
-�ٱ��S^�$��`��N��A�9Y4�om��a~^���H"�E��,ʘ��yfS���k��j�jM��j����w"�BQ��7"�ߞI_�<�7�_`1ݎ[O�ݶ8z�������p;���{nu�*��������6p�Zz�����XM�_�NO  ~�'0�Z`��u�S��Ѭ�6�"�zl�;⥽!nKT:1)܆��,�SͣK�(��o�~C�
Az��ܗ�'�r-�������q���F=�xp�]M��%�g��hs.=�hj�6�"	�#c_Lx�o)5Dl�Z�mޚ�P�P�.��3��h��RD�m�I����0Ҫ�]XlBv]����F���g0A�� �Eٝ0Bk����n�칠^j�	 �SY�ٸ��[roĞe��^{�=N�����`Ǘ�x��AjƖ���UNH��؀|E>��$��^[�-C ��~�@�X>�4�:R�:�a.k�v�)q��m��9�5S�J�&�|���d�*�[ϒ�O�dc\ ��Z�	��^"A�9w.��=�����~~3~��p�,&�`ѭ@��7�)�D����;���|"��r�J ee���=�S�Dz|��*��0%;;2�X/�]�Q��Ø��>�_r��ݮ�J[K��nG���V	 h�Ϣ�}�J�v���\�#fn���g)�ک����4:��p@hl^y:mݬ�½��@'lsF`�AvY�$s�������v|���j�"H �c��9 ϐ[{Yf߲��ۭT��2$+bȻ3�@��S�sƫjD%0�2���d�͆�^�-��}��7�I��}YR�V�g^�x��7���P��ح�e��ԻK�k�IH�`)L���O���܆���y�*���|�t�(�و k:�u��-g�����	�x�	�&#�
#�b����<.�e���	�K2ؑ��^�3 �͔�&=��������9�,�)���x� ���x �0��n�3�$3�[�>�#��@��������?�~�.�{B�Y��D߱u՗� �sn�	V����w�����x��9Ek����\�'�O�]�'��p��F�z�C��}�tE&{<=U3ޔ��n�����D�jl!��ЀAN\�0H��{����X�gn��[>jӑ���$�l���۪'�ƬA�6*�o�$�U��,���Kx���xuӆ,to<A��YM-�Y\�,������I�ق�x`��^��>']�TE=�c؍h�f��g��UOQb��F���6�zw��r�w�M=��.$���Ё횼 {�h9y�ݶ�N����j�������<�A(�O�-d�u�@$c�j�2^���e��M�s0t���f�������_�2/��5/q�`��A�]a�O��P!��UwM�g!3:>J�xݨ��K<���J+�P{�ȀI6�'5��s�Cst]�M�� �S��(z�։���m!���x�����{?(�\3x�M��'��𓲓uk�*.^�;3�͓���sB�7:�=J�I��u�]3V^�u"B���y�ۮ�o�=�t��F� O���������+n;�h�	���}G[y��$q�9:&eȕ1�X���`69�Uie� $�mnw8A�5��ո���0�� �qN1�}8:�`�^ś7�{7nv���7[uѺ�� .�F���7X��`����K���#�R�7όy�ύB�<�k�l���+X��{���(�W1�G������s�6x�of�ssR�HKu���'�zz$N��b��z ��L�͆�sY�ޓ�D9ʱ�T� ���?f�6刀�H![a��F^Sd>����:���	��o�֩�1ymscKE�d"�C7�v<-�@$7���M��ɫ��U2N�l,��Q>$�k���1Dd̃h2n��X�l�:��UPLy�k�rA'v�S8ji����y[��"�쟈e������g|�u�A��SU�������/kg$㻓�9�(�M*p�9ER�kNȢ��RT��d{F�F�]�@hݦ�I���l�Iz�h�����7H��I���|����m>��]���@!�]숉m��ϒ&��"}x.Ă�v�@a��8��>]�^��+4r~�c���{n\`�t~]*��QOB�<L�\������:�4�*��h�'M�|YX�18�-�9��eYfȄ=d !�M*Ŵ�
���O�nD|���-��CV��>�H3�j���wv`�_�̳��䁜؁�"<$�NUekA�O�9���	���O�����X�f��<Z%�Y�N&�ǝ��$];8$��I#LXl��.�⨓�Y�s� �x�I��
�-��mp�=3�L�h��UC�~;�N�FK&Ӟ.Ӂ������@�=��꘤�k��lX�]u-���.��b�ݦ��Ez��_���w��,䶗�g$��P�	� ��_Lcc6񦴆3�ӱL� ��x�Vܶy�"�\��܆��E�S62���a>$������H5����T]2��Cϻߎ����v{��ZƂ�4~��o'w�6@H��|7<˙מy:���^�jq�H!L&��u7SYsB�eb/���w����;F0ּ�^L?vw������e��u�������׃^���@�������<�g[��e�a>�&l~CU����|	l�>3vC��9�@|8P�դ������
��8w���.k�u���q\�7v��� rT��_)�g�"���c�2m�����q�چ�_N�3�Zuק\�f5F�u���-w=�x���yN����d+_���`%��f���9zz�x����>��+��u��^j@1��k|���2E����D���6w(6�t�Gb���=�'w�<ݡc�S���K�����9O�,u��w�JQ��]�rqZ�����,hg*�Ո��L�{O�P��6v�nK��8�/D�w���i[�V^.{�����w��d�GT����_\�<V\���]�w�d�=-���=y7x��C�h�%��{�%�J4Lm��v��z_z� 3&�ݼVS�.�i',�=�v�;q����!G}��ٻ�y��&x�'����Cb�Z��^:1O|�%�qw�>����~�ʲ�$��gh�0�w���={�ɝ�k��!?�3ػ7�Սx��w=v��i��_W�\��3N��j�ž�&��S��c��� �8%��̕nL��!�Z@ʠ�R�Ϋ�}��i��ay²+�=�y��|�x���?M�<�#��3 ��&O$�eU�������'�a�y��Ne�=E�s�:��u{'�{�9{ϦȨĀ��+H
V�"�&.Q�@Ec�� J�G%����<ϳ��#m�OOM=���ۧN�jMV�.�Ƴ\+!3d�$d�W�"�ݦ���!dqql�\�1�

�$�*x>=>4���ǧ�M=���9����L�!�I�ň�Ӯl��2.`"(*�H�
-�LR*G�Y���p�g�㏍1��M���n�:j�Sr�a$�V^n"!���@[$�Z�<Ʀ32
�(#�F�sbᩕ��I'����D�2$bG�X��Ԫ-���W�����b�G#$H�"��ɮE9�3>�)�X��������4�޴�;��[�1P#�$�#�)�
�L�D� �Gq#+�I(��:�E�b�Y\R5
�LS2m���b �\l����r[F!��#-����H��5�ɓ\6�H�����2�,sP�U"�Z4�+[`K���E"AțH��I�L�l�
Cʸb��		`�dDQʬe�L�5�x��bF1�D��W�=%A)���/��$��=��c��� v{�L���ݰ�}�� �%��D���{bgh���
�Pߞ_��NN�@�-D�D�:���`�D�5����֢�{���g|��5�@7�Y
�Z��/�0������*Cok�.�o���0���$0|����0����>�گP�T+���QC�
�x���3�w͍E$�L[�D�%��u����f�6��Y�
H���xrd2�Mb%���^˓0��RUk]AKikn�j
�4�C�'~d�.]�e�C^P}�P�yy�^A���鏵�fޘ�B�T&J[�A(�|�z�nTnu�35�����L��U�����L�pJ���ߛ2'I��ʗ=�9��m��6���`q;`�=֠�;�T������{`�{�W�<b�$Z��j%�{߼��<"T{ߺ�]���cq�;��y����� D�6�g�q�[|�M��Us�'D��y�fƠ��RA'�����@��HM���s�2o�3�M����2�.)"g~�{�ȵdB&O�������<����m��%#ȏH>�7Ka��m�yT�v;E<��}eŸ<�{��n) �	;��j����Vҗt{��p�(�|�N����P #�;̫�`SU�5���
��[*��,�~0����7NȮD��|�xI-�^łW4w���uֵ:=i�c1�H ��#�Źdk7�ơȅC��}u+.���:�����W����@��E�s�o�p��C���2����`Af��J`��1�9]ښ`0���/��� �끙}f9�V�DY(%󤟥�y ��0�w [�Ͷ��=W=%�ۻ@�"ҳ�����i��$�������.�c���cQI�$���2�.\�G�"l=�$H>�cp��|R�uW��T�'^w�v5ЋP(�P*���L�ë�:-�m~\��g�7�א9 �Z#�$���o�����l󇀕 �k^��7����oPM��b\��[vy��q�QlB���wV)�H�� y�G���[of�ݺ��jw�����0�`���w�9�OYQ.A�5[���&���{I���5�I��oQr@<vӨ�!A
����^�8�:��~��엒�# �|���fy*�����߯�r)ƩI�{�M�J��D*׹���H�Ph!�oݍE�Y\ߚ���� {���W���Q<|��xUV�R�ʮ�������.D�Z�QI�zכ�{���u�e�^{���PM;�z�l��İ����^_Q�$D��kݍE$%w��v������e���M��l�v��R��~�2��͏c�ck	W�~T�#J�`^��G�hє�
���)���9�kɽ��-��h#�VN38�d�ig�9^�]t
Iʖ��0���du�]�6����㋎8�P���Z������k�����z��6���%���(x��Y�`]��`��q��Y��.�P-(]c0M��̓�%z2�������I��bט�l#N�2m-!��0svقke�&��p;��2���g�q�u�M�"�Lʖf��"ք����жZ�`���Xh�qv`h2��xfK�wa��͂����9}�y�nxP�͎4C��2ˈ�7m�+�e&�3g�����Q�f�������? G �PYy��1ye0	�,����DzO�#��ҷy�`k���y�\ ���`����ä"r8H�}����a�·�N����XCok���p�뽍E8B�:�^k�^��$���E$��,�}�}F�;�"�Th�ޮ�'��"W��Q���� j�wp�L������l�>�s|3���k̼����zĲŨ��Б0��0�>�/�ty7ủY��]�w�ܨ�J�UQβ��n)"��ߺ����dIs�v~-��wn�^�� ����s��;��1���3�㣪��y���G�TN�5����pd*�Q*-0k��Z�����w}�f"[7���D7��	'y�ߡ�7��j��&J��s7��NU) >Oo<��J�~�y�ws4���C���]�9�@*5y��Ȥ�H�������TOu��5�ח�%�B�}��ʷm2�7-ж-��`h�JF�FX���ta��b���RD��ߏ�IwK,g�P}bT/\��p�ȵ���c�^���2�t�*) �����	�PL�W~Q5ɫ��]+��������	�*|�Gz��8b�8!�{��o�*۶��xg�O��������({<�����3��OH�OH��؋�s"�O�Rj�Q����zɻ�o����Ҽ�3��_��q7���pi�O�Q=c0c1^0j�y�
b�J'Q.'|׻��<c�\B�T��5qv*Q����|�{���^Ӿ�^&t�O?*)���U���XCW܂vv���^�{NJ�QT-BwY�)&���D*������Z5��=���qI���9��9��"�q���[�W��[�r�첽�4�t���q��(tݏ �"z�x�fd�H.}hD���%<ѫ^b] ����L���M��ݓ�2�g4@����B��l���S�>��O��2fL�$�=��k�O����Fe&�FBFێ�A�g�a���~�]v�ekU�n;sC�Ov�-��L�혭n�\':�j��>�9�6����?E{8�HA#w�,K$�_�2�zms@��c���jH$�
�$/�RL�Y2*ZR�i��fs]�Å�y�<<>����0	��A]�D��=�Ҁ�J).�����n�҃���
ę����{���)ט�����rs$�SuO�RH$�eS�l����5J��,���os��M�c��o���͕m�ԭ�r�ޠf���U���h�R��I�=��b"�(���l��W���>>+=��f�8��U����oA#l��A׏ԲR�4Z�XtS����	���g���wP30x8$c9�W��|��%��@L���]<�+v9�VyUery��<��\��c}�2�3G�:D5��#�֢BI-�l��.��y+3hm?7�OxA��3ǒA#��(	��"[+��O���.[����PL�X,��)��0E����q
�ʂ7�n�t�Y)�,`6�c-<���}ɸ;�wv0���VN4�k��zA���Q9Z�
|�WJ}h[&N�_��ĭ倈E�Sϒ��)y{3����t��y(v�T��F����i�i}H��.�]�b[�*��S>	 �Hm[��	 �lg���������aU����$�3�Q�.%v�iԲ6 ����TNp��ke����=��x�0���E^JP	�|�Md#���'`C	��i�i�/[�i�@,�W=�
RI �տJ���H��g����0�=�M�{�i�����kn~�p ��?z���ޝ�+�:i'��v��t��N�uB"NN�1���ݹߧIpD�Ų8��*~�bc�	����{�sǏJ�
tS����M8�7���H��D.y��be�|�@$":(̄�Huk䀧�/$��f�֘\�]�����~��%��������id5�/X�葎�c�-�GY�]Yj���nt���}��S顒I�x��=ʒR[X��)$�[�����h��L'-�@���''���+�,�~�@23�V81f���������@ �̽�!�]�d�60���R�H$���T���(�ƀ!�ne�3�l������@����˦�7���"��{-s�eI/$��sI	�3�Ŋ:S��X��h:L����R����K�!/^��H�'E��i�\�66Ytx<yy�ZYp�����:A$���D���*����,�@|�*|�ٙAR�f,Y��� U�=M�H%Z�2O���됾��XI�z��>d@),�`�` 7�L�;f�q�Ҝ����X�4n-��z!����X���ogjl\�i��3������a]4+�Y�RjM�o��ڟ�
�\s��%:?O�L?�9�6O�C
%��hF-�H��9�d�'+��&;��|oŸm���h)�66�Tc����n�'�v%#�F�����,�yU)M�*�&m�P�-5q
���1T�Ӌ�˲v���;W\���W"s�;V9<���s��  ��mv[	BK�g7��J�K1��#�F�i�VPa)e�u�� e�1�-n74Y������������z�ﺠ�Є����i��!Ml։�t���l�ي�k�3$���<�A9a�&�גd'f�~�&��rL����L��P�C�S�qz=�^MĚ�d'����f�I�*EäZ��ֺ�|��OFN�S���>ވ�'<�H��9>�{Y���S(�����·`w7�S�_߶�6����L{0�z��X	7��e�8��m�nVAԗ�A ���Ч����b@@%ڒ��Őfp�BQ��}6���*M	[r�	 r-�O��W��$5�(� ϒ^�މ5�����lğAQ���o3/D�ٿ$�2.��o~K��%JH��{�%-�O�bse��l $s��I�ד2�ɀLd�<J#���n&1	�ă�ٵ�A* �y�D��Y������e�K�a]0��J�h���O�lv!	��_[�͟��@ 7���J���̗WLI �-���I?sD"��Y�f@@�%9�N��a�w�e%�a����N�RMp���~�\�y��N�4>�G���On�U˽-89�'��p��'_.��.t$� H,eS,����[�.J��� x�N\�I��3y-�y�)�~dY�z$ϣ���Pys�g:/&��$&�u�LY`v)�hw���P|����u,x��H��ښ�=��٩��Ҍ��~G���pnw�%�?b1<!��2�L9����ۡc$�	7C܄��I\�D�������[�Z�@����m��g�w,p1,S�r���-r���y�̳�ץ��l��� ��}~5I/$���҉$�J��S陪��-���ﮝc�$Wz=ԛV[�w`�����#h�-��x���$M)����T��G�߳׿�$ɉp�TI=[6�*PO�^b��u���J��! !�z���H�uf�w��Ř&R>���R��ğ�
�;1�Bf�)�B ��r>&�+"����7��1'��](�H��� ��8�T�`�L^�>��B�#\$��K�%�z�d�H�_4@$�Gj�mg�0�������f�F�L��!P�*���3;8�-ͼm�܊θ}��4��d[,)'${�x-K@Ƣ���?�>���?'�"����@R�$�;��I�E,����C�N�hK]�K^�M��PIf�U�G�W�@$���H���An�9��e��TZ�bY~���[C
L�*�����)>n� ]�H NtW11�Իg��ͽ,�PH5�rsy�I |���H��;q��-��=� D����[�ս�'p��v���o5fDXH����X��t��b���� �}��f$�l\���H������ޏH�w�iH��ݼ��G��GM�%�t��u}����T�_׬���vr���k���,�4F3˷�|&QI7�_]7eoO�$���iJ ���وv �H4K��$����K{U]�C5������A$�K;�$����7�%QH�p�p��M*�S��(��&�����̉�Ɓ~�d�U}��3��]��<2�r�9��&v��!A�dŧ�id���'��`�"��F	����Ո�n�/=��������i�==O��`G�?��1LL��d���N|�!/^��d�a�vI�k�Y��'iG����UzA����>^)yTs@y�27�0'��d��[zX�<6�'��y��0��:�eA��k��6��s�70�ƒ1e	t����UC��W}�����Щاu��	5[9�A,���@$��]�ґ�Hʁ�)�R���3��IfvO��)-�P+wls�	�]�3��Z�eْ��ɗ�h��g�� D��el�������RIl�(��}Ȏ�o\1����(�1.�����|e�G�:�����Gs=��\�������2�Iy{�c�O��d�J��,�`�
�,�t�y9�XY��'�����C�_eJG�����<z�u_iԐ
�#H%!^n�E q�&.� �T�:�3�I$ ��D.��,6.�W��=Dq������s5��UUU]���a[[TA2���lI�r��g&ň6�����������̓��^���o<�����ۋ������a��%k�o,q�]`�ZM�<#ʻNśzlg��G�5�z�Uz�/*��M�珙�����rg%��#��nq�6V�=���}�U��|>W�z��C�Ta[������v�ƶ�V'�G��V�>�o��g5;.KC�U�"�zd&�W{�q;%"C�oz׸ޖ,�O�7�y�|�)2�2��=�A�wOh��ϗ��{�Z�o����f�]��v<W���������Q{{hc+���6_y=����HNdٻ��)�{ڰ�����v������d��727A�p_oz�.<i���Յn���y�u:��ۛ��j3�ό��:���+�����f��+�[��/���%]}�r�5�0*z�6?*�xɮA�@���}[;����]��`{��7��u�8��/�EM�u�#+3)갷g1��[�ٕ�=��o�������0�<��
X�vT�{7%9<��N�/:s�,~�������A%�^Փ��DtT��w
�[�o������v+$��א�������o8��}�5�`3�kÌo����[�:�����q���<G/b��Lv��}� W�lTA5b+���v�;�yk�n���cq;��0������}d�&����z��w`ෞx�>"h[��� ��O�������.D�q7���%y�x����wviJv�SI@f�����:���D'��kNB��̣ʪт=ن�+��jk&"\�ı#�^�n�E��QJ���с�9��z����k����5����1?�H��ns\�q��'�<���{ˤ�Ry�F���dv��͑��Zu;){�2�<̑��5�V�i�4n��I���_�8�Kɇġ(	Ɠ��O�Kc��T�~�*�XH�c>���n8���qq#l_qٮ,Y3�.)	��.g�:ϳ�L�>1����n�}x��M��T��J#�F�	 �FE�AQ�1TNYd�H�r"��dƷ,g�	d�8��H����24�ǧ��q���ǎݺuʅQU*��y��Ԏ�r8N��I1dQũ�S(�����X�B)Љ.>N��;�q�:�<{{m�ǧ�;v�\��*�/z�u ���Eb�%����(�H��LrB
1���$�$̎*�D������G$#m���)!1���e�ED�0�zIHA]I-��f+ ��E��
�5�5̈�a�QFTH�A�	��Ȇ�l���E*�k��OraZ+�)�ĐW�lrB�8G�(�qGY�M��H�!0\XHE�E��Y���*Rb�@L\�cm��Qa"�
#���Л�IX���Qd�R%��8��L����&
E�J�&v�RNO�a�G�%T�&#��y`)�a��Է#\�Td\VB*��1e*�_aj@UNl7ln(�&�ʮx��L�Fﱾ**�;��U���e;���;i�x8�Q�]�2om���,LSL��he�[����vK��6㜄�1q�6�Bn6k��B���y뫮8�1�en���S�-R�����:2�k6�x��{(�x�n3�u(bn:%%5�M�»���L��::Փ=`굦1[z����&������`�X�	�uv^A����'�ܥ���gcΰ�6͓�8ƼhL�^�����pkW��R��R��e2��bn|����d���"�`,g��.Fs��<�]��4и4 n�7��76�FP�k�sD�B���M.K�=�]��<��A۩��8}���DOm�y���Q����-#���3zĎ�&q4���4��F�M60a`1Rݵ�7SH̓&��`�E(���6�J3@�vۣ��y�;�è���Z�і�thi�1�fm�԰������rsn"X
$�smvA�h�����l��n��׉����є����l�t��6�o�d¼�j<�$�t���k�b�^	�k�MՀ5׎C�a�����O���)n�j�Eqj"�M�7��̪�H5- ɶ��We棜�Ա$�Fa-�2<��^�aQ:��7k�����Ը�XU��� �u�����t�X@w7����v��QΝ���%���p����^�x�\u�/��KT͕�x!�q����宨�8:np��h��u뗹�[���ŝ��Ŋ@����Ҵ�2ĚcS���f
H:":�!Dt�,] 1�,a���iu؂De����'C`��m�ه;�^n���d� a�M/r�Ե��=�'N�]t �9c)�U-͡�C4�j�&��K�@\���h9�d�tC75��2v��7.7>[�!z���)����b%@�s1L1C33C��oJ�H�k�l�5A�]�����5�&�'c78�=�4\��%��b��`� �4,hH9�U��Z���
s�(]�m��g�huɜq�������q�³PhH]t(L�:�aY�#�WVw��v.��[��Zv5�a��6ԝ�pr]�Èji31�hbX0���!�7��s'*���W14��yz��v�n��Z��+Su`�������R�9d���%�(5��N<F2%$o���/n��a����n�݊����2�}~�)T֘;�'I:xy)�h�����9�.�s�J{��'ȢP���R��Hy �9�A(禩B��W4��m���Y$8t���x�n�k�n�0d�E�!/y+�\�w	��&)��Hk3�y��^I����o^�$"�ĸf*��MS>���+b��`�O�S�t"M���f��<�|��x�X����w�ݏ+ow�.��R36�ī1r��P�	GK@�I ���=/3��7n�0{���5k�$ͭA%�-��2��w�h�&�w]�E;��"��^M�sK����k��({�����fp��%�����h�gI�'�k��J<��g$�@$9�9���9`��ހ�*]�+̽e/$�Y���H^��fA4铖k�@'���4�+�N�9���oy�5Y�Z��=Cl��eu����C������w�vnx>$�L�2�sͬe���YbqՌ@�!#;��˓�� �b0`Ȍ�"	�F���L|$�	 ��y�I%�<|�J(�I��Ɲ����JH7�kL���(�%ޞ�K��! �H�n�|��	y&ک�34>+	$���D��9H��״3\$d��v��k��}3kT_��A#}M�JIgDY��I$2y�U�ξP�����D�$����뱓��Y���SW��ǩ�������}���K(��j��KJWu�Q�� @H���(���f:�*RvŻ�����X�`SC�f۬ڡͤv��,�ڔ�ێ��"G��Z�A�����鋲0a�;��m�g���H%Yҥ%��Z�ޠ����褡Vt��,�����>��2�����ᙋ:*y�����e���,b�'������M�[m�� ��=�����d|��Ф$��N��c�k'/�� ��L�w�2r�����B�	��N6EH$���zw�(����or6n�ROI�c�����z�V�>�&��k�
P���;�̼�2���p�陠"���|ޥn���/���� w�#PI�%���U%W~�~@���d�O���@*���݃0t�4���^����8��{���2�$I�־B���^K{Y���w�����R�}�8��C"L�햩D�	5�2�'rr���H6�T�I$�W?J>����bw���v���s$JHAX嘻�N����竃h���:t[��톊l+�WfR��3Y}�����f%�1\ĭǞ
I V7D�K�ȯ$]��Kv^."��.�� $��J�eyT�;'L_�T�])�˼�{*��Y@>�hW[�N�\��'<�T�w4zA(斆��ҳ&<����m�H�N��p`*�(�m�@��f�#��}�v@$�׸cmˣs�>^���R�	��S5(�$��L�*� �-�蛍3>�3�l����I%�[��Hm��~;�Q�i����gq4����y����-��^��y�{EVZ�u�� ������'��^�c��z	>(�'�� �b�$U@��*�yR��0��3��HKk��	 ����"L�Dc�_D���o��p��j�A%�[��xI������>3+7��^7�d�D5v��d��.��4--ǌdL)շt��c�sZ1�1Vy��'M��f!���z��!\ٙ}��i�d@w�K���h�%���Qr&|�S�[eu���"���R�y���i�|��,t�!f�"��.|�)B}����`�Y���C%�H-�h �`$�y�e�L�
K�SXn�Zϙw�E��]ꤗ�۴�:vL�,/�ɨ��	$�>��yW�����LXǝgfuSڻ���	Vk@�W��K�:W��R����49'	��pHIy柣{��������H�L�@	f%�d� dl���k��}�qf� �w4B^���̷Ι�;UPI�� �+ʼ�˲�a!a1�4��=)�H�s9$�n.D3^oG���[�a�t��W\�M��yL���jzO��=kn�C\�U�5Y�w5������gd��q�$���a�]�u��vcn���0�@��27D�d���s
��i|��cn5��$����`��D9�'8Yխ��2����|��r�fC#3맸'�ۣc������5�/[�7p��^��u�e�]i�2Z�x�cМ��ꇂ����`�����E0�d����b���]�Vr'km�3�����m�z�qUL �4��BcŔ�:�c#���UN�<����;F��; �/W��I�C��e�[�D����jͰ��4�,e��߿~߱�-����S��� �$�2$�@"Vm?J&CN\t�'ȩ�g�x��^Yѳ�2�d��%"؇`j�F�D��/��Պ�1��ܣL3���q�&BD}�OХ$���4�U]���$�A&�d�!33��V��T����u7D�Ag�n��i��Y$⾍�	�i�,�~�>@%�Au3�d΋�R[2�<24ұ
3/�"�މ�RY��YQ��$I;���`d�����A|t�M\����CN��jN1䚿'�k�d��H]��aZ�lj�s�z	3Y)$����R�����ٔ�N�jje0H�)�,����aͮ��;�/��gѣp]�na�֭�{0S���k��?=}�c�칙���	7�&��%�-���K�Z	&����p���m�O��D���1���\W`����J�*��iM8m��x7x����]�f�1uӆ{����i\q�z��?!�&��<��_5�@��)�]��.M�L&�����<�u�$��) � �"���*z�<"�A$/���! �'��p�#�64#�3w4��W�/��B����Al�\�)+�0��$+���fb�r��������2:��
D	�p�I��I�z}�m�t����z�[�.62&w!��;�����H}yOЌ��H+�h<���w@5q��2�+�%�~~�5�`3�(�t���ddI�x��h��2L�� �7N�_u�=0�A$i�T���9������2����[����>��:6�-ј�V3Af��p�6��8鸍�	6^u�Rj±��_��}��@{k|���%�}�f�H�F��0�	!�"d ����y����Q2>D���?�W4Y�r��;T߂O�tIRY��h�7�ٖ׍�-�.J Y��U�.�	�#L�Wy"�������,�=
��y���e_�]�wb��%���RI%���x$�
2��Ǥ�=(��>�ڷ=G�p.��&���%g�����G�u��c0���x����ȻH&e�W8���Zq��E�"'���A������NO������l4D��Dqe ��_9���f=U��Ms�+5���=�Ƞ����K� ��3��3!?��/lk���;x�%��Y*�g0+�c#%�1g����a�|���U�n�x��A$��<�D���S1�2@/c���'�p�s&'�	���,A����h��A�͡��,��#��u�Zm�b��?}C�fr\�[�<�L4z-�H%\�R$��6�*G��/u]mٞ;���pU|�!G�,�|���m6���8,�;�U��n��@S.ɰ�A׶sh�WOҧ}^l�u����]�5d��s9����w�$S36��;j��O��-) �]8��I$���D5L�T�J欎�	Ey :m��� �G�+��w.Y˳&zr_��"�}�5�$|��i��JS�fG�������IokN�HXIkL"�D�۪���"g��qX�ڗ��o��[|�E�a����vᯝ�	C+-RpYUe��!�^`X�¦�}�o]l���b0 ��-A��*�UD��𪢾{�>V�;קq�^N��0U��~h��ה��^mn����M�w&�I��;�~�g�ߵ�P)*��M�,@2�.�h
�F�ڼ��l0��a	s�--�X:h-�K�[��1W!�J�Xղ��y︖�����s�3�y�҂H$}R���|A$���^������vw��mO���eL�� �Z�Z|	VH[L��3�傡U�醈H%������ޅd�j��(.�3$6�6ZR�/7� ��3�H�qU���i޵'�)�f!ؘ
yD�ٿ:����nƈH ,"��wbO���o$@+%�e�����[}
}W"�������;URO�X}��o"���t-�#��������R�ƈ�32@%�<�T�7=O�I�t1 �O:,�N����ZY:�	��L�h� �;�Be�zZK���c=CLy+�h��@I%���C�gϽR��|���5���� �����$D[\dP�E;��D='k������8�������ٯ�|_L��o���[Ნ����0i��[����IFF�t7+���2
�1j
�l��S��Z1�3<s�Ўn;;�U����K�:ʛV�kRhl���������sc��z��i=K�9�u�͎ �HF:��	�-ə���B^���\&�Kf�5؇�-���Ώ2..��݋@�н��h�d�м[F��;As�W���s�n�ڬg�v�a�����o$�݆�.�T;s���*5[,��&��6�� (]�#��(�iKՖ�/���߸-�r�)�>Zf�%��b�ƘD����)��1,	��3R��P
����o��Kݢ޼C0b��%->H��](���^sSD�� e��}�J�� �1�� $��x�2�Ƀ ��]r�v?�����re��,7-��������h�� Q4er;wYuխ^H���^4B) �x�B����pȇb`*�� �/u�3Nkp	%��]��	 �I%�׌RiH� ����F�{�,O#1�l�y��2	���m`Ag��a-�=�`%*�#���<^��Iv�D�f�K)�)!˺	ߝt�?}��mz��nM����Ku�D���e�Bf�aL3]�Uie��ϟ�=}9���?9&�h�I9mJ*�3{t1#[o5��YÇ�Ȧ�hI/�v��})��Ȑ�˲`��q�� @K2�l�<����oj�\`����ID.K�p���<������yKrh�ܦr��`�؅��&�N����\��*�%�Z����"���Ɔ	@A�I��Q�G����y ��_sƩ�$�H_} 4y%��Y��h����^���A��RR��k�$� ��I$|��n�I��.f>��$Z͙�&RZ���/�x�`�L?�����ل��l^kf��A(�~�)$	z�d4 ����|�Sv4���;]T�C�" �����y�d	��f5׋�D;d��{t)#լ�`ɷ&ԥ@3z|��ud����I$���?��B4lS���d�"��!��2�#�s�q�ٞΡ�'S�<p]�c��m�c�����$��A�O$�O���Q�fA 8�@ �	 f��<!�C?S����<�f8ȔR+]�В껍(�16]��?���{��w,K�_��fcƅ'Ȥ��� �@%]��(������Ǝ�9)^NN�	ܻ&
�����L�%�u�z<�,��7���<F[yn�
T�p�j6�2z4�6i��N2w^���e�"MVP�wU@��[k����'�>����{�lo�6�9<h��
zk]��ۉ?S֩�r\�4:��|�	�|�K���-<��&q^����\��=��;��fVN1W26՛0�F_�A�Ci�V�
�g�������g.st���B2����S�:��Q��0�O���9gw��g3���!r�s�ݎ3sð/b�8�����H���x�۰��S�������Z>������3}���.eyA�BIX�:g&g5�hx��HȌ�=�孵�O8"7�y'+� ��'��="��؊]�p�ӞvL�)���φ�zY�g�*J��Oq���TY����uӣ��H�&C<�Ѿӹb�u��k��Ȼ�.��uM���Ml[��r��j��vO4�We�@�P3+�>�^>OV�~�:v��4�T���/`6�w�k��F�j���P�3���E��W�<�ϥ�u���'n��n���4�(�-�琩9[CC���.~�C=!>���:�'�}�J����z/pc{�ϲ���6�j�=�9UB�g�0����i�ڊw���m��׻��b���x:=q1���}����=2�������z}`�N��=ݗ��O�S(�Vz4X4%K	��%8����LS��3������*SI��>y�̐��2C�ĳٙ��c&f���'+�S,Pw^� �}��,�Rs��Oa�+�X���XJS�;�fk6,$�K��jt*�l�u���w��w���M>���ۍ������n�&�#D"�H�F1���䘍 �LQ$��Mu�,#�b�%�!�{�>4�O�{zz|q�㷧��:�g*t��$0I ���|c-,��1	e@�P��P�k!R��t�||c�L|cǏon:|v����n�m�U$�[��UD�S#Kj}29�"�`�D��*[�E��$��U*V���X*�A_Fb*M�U#klbE�QW8�����U��$�ET�
��Icq�	#&UB9,�����.t�nn^<AEA�I�d�E%�jW5����bELX�Q�!��1� VH�Y$W�c܍�Eqrtȑ,`Ȧ.A�$Dc��uI��6�R�E��&(����q$�0U���,���1J+q�$C"�H
�VL\U�π���A�N��H�  � �=����>PU��}��d$�_��	y���+�b��d��.|z�pL�ζ�|������Z��@/$gu��@��Q����!��X�zs��2Aݶ Q�_]��ӦvtĶH3�E�a$&)vP"���.T��AP����$JK;"�IgLq�M{�e�5�$
�"��ر��y�u�ў7j�QN�����*f$�U�k�R|�}ߓ���dC�'�����y�W�D��")#��/fw�Mhjt����>�B>��d� �o0!m�$��D�w(:�5j����!I�,Ǧ��c0�Z��2AV�@�H�O@�M�5ch��<WbԚi$���ҋ�,��Op�U,�<�K�r$$��)����(�wP�4ӊ$�,�i�"��7"D���I��˲`�OB��K��UrggH%�yD"^]�o^TH�I ����6���[��קl�z�qw7P�-y"m���2gn�*����=��^�Qɷ��)�r �l�/!����n���N�F����N��^X8����Hy7���|���1R�� #C�""VUQ��]��n�~uH�ߍg��r�`H7L�$�U�^&莝��U���I�[v���	%�7"	��st(�3GlPn��_A��;��p4���؛۩�Ol]Yt&�a;[��v0J6��Y�g�ٱs���g�
�@��A)��e�f��n� $��oV�2��T�	�\�p(��̜� J0j��-�bLHOˢ}.���h��anД��gU>�d�K�ڙ)$����BI-&e
���覈U��yi,=��w(:o]�J.2$�H�Ŏ�0%4��<Hi��֪Ȧ�	���dA2����t(��7��`k'ɜ;����fͦZ� ��|¼�ɼܪ�A2C��f 	m�[�01�(�v��̗�v���Y����EM��ۇ��$�I�w����s@�K]�6�gO�����R&BI$)^C	 �_4OqL��9\[�;u�c��4?�o&3�_� �б׎���m6rJ�{�$e�]�+�\X�Y�2�Y4��)�q��j�Oo,�&J���㞤��"X�6M�ܨ*�CY�:ۼ9���M�P�%lEl�����h�]��UikvSgف����0LD � �
����������X*a�K���%]-Im�5n]�z�;�kp�^kupr˩(]	�d��B��\����y2{'C�d�8�UA�/nط;x	�`yD�K7CKBYm�6SBn1��PFY1f/����.��Mj��^��E#�7c�n�`�q5�[�$]�$n��ͬ����H������tیrQ�n��C
�38�X:ʁ��l ڔ�Vly�o,vԷ6W=Wlvo|w�$�ኁ���7m�ђW�Ü��32^[���3��vʏaܕ��5oH�(���z<�{v���]�dZ�*҇��H#��V�r��v�"0�I$�_C~JBZ���Ly���6v�1��8JS�s����Io;v�4؇K|��H��G�$�J|�.Oi/-8(�	.W�ē	ns@��f)+�|��P(�O=Ѯ[[k�>��D��32�xt��I,�c�$��#�j:�5�A��4z����s'D;8vr��݆�By"[�s@���mp�����L$�U\���e�=� ����즭�	�j�ٖ���C�=G�ma�����1�c��X�-p;��f!�׬�X�w.��w�	�y�� O���@=04oN�Ȧ����`g�`A�7^H3$�TeK� �:�_c��-���ޜ�_�&��㱯��w�xp^�z�'�gǽ�㯺{�u����G�����kRm~WJ��0n���~�"��|�PE�����E����揘����ܐ'�|�D���-�����_P&=�"B�gEܖt��V�"�]7?Nz<�(�[���[Me����0	"__��cP���o;,�� 7]�
2䨌��L��6Q$��p���y9%�Ӏג��x}�ȡ]��w(:����H 3�U�#*%��g��Ɂ �9��ǉ/���aQS+Nt��Ws�3���r�Nn���p�C�^��9���Q��v,��u���܃���~i��M���{���#��g������nYoٻ�3�̸����D���61YܺfJ�wMDkDV�'����$z3��D�+;�<�����Yr�°/"�A��u�A�9S'���	3]� ~T��+�ih��:Ⱥ79bp�t�f4a��芸�tB�b��������ly��M�Yj����sSpíދ�h�� |���� ��� $Qu���BG��� ǐG��@��w%�1r�D�Q�F��f��5�&�	 ��ym�B}7�:t19�� ���#9!��L��\@ ��[��kSS�F�{h��#Ē/�`w�_�c��Mԧ}�M��m�C�t;��o�Iwf�DD����t�����!b�ӊ��h �n�6��o�9ړ/�-� ��}� ?��z�;��f\�s�|�8���,���'�8g!g�tc����齍!�ol�cω� ���^���s���/3����$��9���1b���2S;ힹ���@��y�ܫ�̤c�Tk�[��^Ё�vl@�~I��㽻�/�y7�܅Bm���!��)���T_@�[�^�d�}�V�0K��!D��m55o3C�����[i��b�=7?�n���rȼ�W-v��zկC[�|O��q{E�r��iAv�1WvΌ�! b��i$��U>�@����TQd@dA�|��w���~=f�7��f.SP�n>�I9����t������'�"'�#ě/{�"<V�/T?G�D>f�<�z��GȄT��;R`nlM�*�]ͷ�L[Mk�1� �t1n7����u����rC,��鈀H�+g�W� ͽ<{�Y�1�{�D[��� �ݝ�����Pu!ts߈,w�r�S�۰� ���	=�� �r4I��:|c����)!����3��A��$�r��	=��$�pi��UאI%���;��Cy+���fL�]3%�t�E_v�2ޭ�*�Cy|_ʲzD@n�N{v�i����y����x�oq��^M�w!P��|�>$�^�Ή�����AgMlM�tA �V� Fn�x��)�3%�e�{nrE�f4*Fr��X��4�̶PA��@�!C��ݎK�l8j�8t#ۊ�ؼ-�"�A�	��̱�F� �H'�"<Gwu�S��ӫ۸6W�u��4���r����PRB� 0eAX@EU�L˭闧]t���i��!��q�`OU<�������Ճ�t�+�
��C����YݜAÎ<u����1��b'ƷgtlqM�}[���5��#��n�4	�[qkP#���8Y5Jͫ�ls��x�4�<��{%����L�N�S����WnR�\Qe��Uls�gzӝF��nJ'\�0px�\�LJ�*
r��PmcNx�r�d*��u��,�X1'�~>�_�VWYü�=�~HJ��q$u�8�����=)�˪}2	7������`�`�R��Ϡ��r���3]>�$��� �Gݯ� Ǝ��lY*����Pk� �r���-�� �	���	#r/߫B��� �O��!�w�I����M���t�9P.����m�#���*�=�	�;ϯ �'��	$����!�U2`�z{ G��]��33;��̪�:���$�;Ԣ�^h�y���H��'�ݐ#����}A-�p!gT�*l�z�g%^(�;�籧tg�C�s���p�"�Z��-r�Ҷ��߇w�X1O��8� ��ǁ3��0�$���M_s��[N�Ί�y#���U�'�6�%1r�����A�g���z?�����w/�u�A�- a�-3{X��}~[��Bu��=9���.'8��]b�͜gS���\6�(T�'�|��>��_�j 0�!C � $��w�_�
�O�3\A>-���A�0��utdf'Q����Kᑿ/]���͵u�Q�&n�<��u�;䏺�`@��~��4��(�!ܰu2w5	���u�N�$��~A���A>��5�5O�ϴ�AuV�y̅�!�w ��^uު3�1 �F�a��zﯣr6]ܙ��kǀ	� ��D?� �ާ���I�Ȅ����}7�\2���M]-��'PG�!��໣��]L���st���5icee�>~������Ywz�*#ĒZk�<A����;��*^e�K<��|�������x���#�#�A��f��/Od��=�D�C;�o��DI�cIZ_+�e�ω�z�(PD�%1r�� \�@��Ƨ��HPz��y����@���YR�vCUEV	)�׸�f�`�sv�i��n42�{¨�X�1o� m�Y�4@�`���w��^r����{��bJ�> "�*�b��$ Y 	��E�w����ݻ#���=�_+���$��.gt�F=|üE��M/�X;�7%y��	y�T~�c��Ä��s���NTD5���Y��X:�-�n�O_c�ػi���B!��Ĵ_DI�h� ���@"�oj"�B�+���U7�#!r�[lu��W��P��7<iAx�4���fdB$9r޺��'%���������n�L�$�������Vrw�|p�]�|dq4s@�%��kD$��vf����E뱻����c�=ƣ��۽�@7wr��2���7H@��9~(�����g�ܵzB��#Ę�s%�py;^򆋯 ��&9�� ��A5�E [����Mr��蓻�o�QЁ�W�.Oy+����0G���6g~f����8I�������l��66V�S��Ȇ�
2�lJ�mS�\݆�9�d�F^Mf�db��*/\eUk��j�ݘ��Z浩�;�X��}���$��Z�!"�"����kk�S���왃�IL�����������]h$��<|Nvl@$���;�8�B��|�=�5���JzO�jm����������]]����mv.�����O���>�w,@�!��=�^8�Am��8��^ԃ1��=]�70i��v.�W�Ę���*��{�37B����o/"V��$�]0$������'+)�	�����BLΉwfk�|�MdA�3��8�3 �׻���${�c�	�������@�0$����ڹ�c�˱�Q���	-�� |wc�q�mcޟd�}۳�H.�)�\��i��}>x�<��&l�n�i� ��\��/'��"������f��y�s���E4G��\�9�׾��K����<��4��=��iɝ�bJ��}- R�{����p8;������,���^a{W�h�ٴn{��zY�%;.�3�����_w�q����o	��FD���n��.�.\��/f��*��*�bZ��_+�j~ۓ��'��^ʼ��+~^�����s��!Ɏ-��g��l�/�{��ϦK����(
Z�d�vh�ˎ��W��V�=��!�����t�xt�M����^����<sQ3��Er��GJe[��C|Ua�0�<ĝ��;u1�^��myw,��bY��>}Ԛ��j�����
˝�{���N�@u��۰+�x�]���jYp]���^��B��$eL�D�#&֔�
k{���1?Yp��G�g���T�j+�n��w��5=뉛�-�!�9�������t>a�W��.����c޼
�����{g�p��d��ԛ�o��õoY>�������q�ȴ7<@{�kh�J�rq6��"X��0��Xw��j�i�=�b�c�jh�<�=�}�����<�� w�tY�@(v��5���&ۨȥM/{z_��19�!w�����cc�n���si���Ded��=5�юP�%���ȃ���9�pBl9����W[2בuIV&��?{��q�t!�qȓ���p�<)"�,,8�_ۧS������ ��l!��}�t9W���3��D&?�� $�AH��#ڇ�?��;Ci��Dcc#���w���.���2��M�S�����	s�
�
��rn��M���<����0_[�A�'�����1��c��}���:���APu��������_�uu�AV�$\G#�������#��˪��UJ�<c�L}cǧ�t�����:�g[���x沓v�Eaj�\EA+#%��n��)RI*�1�>1���ۏ�ݽ<x�:�ǩ$#r��2)�3Xl)fW��Ip�XI ]Qr���>4��;x������s;γ��9����[$ȑ��H��q$2*
��d�rɈ�s���,�;rآ��HclZ��F��#R8Gd�2@��D�u�UT�(�+�Lr�o6@(��{[e"�Ę�㋈�X���f5��%�V���(�!1:��l�A���Դ��d����!	3�@qK3�
(.(�B3,�"�
��"�d��s��0 Ͳ�$I�2(��YPD�EqQ1,��q����qTX䶩���H�$��2)"�
=%���jI{oV1�lf�@��k��͚WwA�rN�b���n�;=��!�8�Iݶ�ٗ��Y�mf��49F	) ��$,�մ���kU�s	�]�� E�&�i��m�#`G@a�W%h�,�7j��Xv��mk��<7.!{V<l~���Gf�፡��y�ۈ��T̮)�����\�!A����n�.u6��Ct$)���zN�ޘuv9e��y�WH;]n-�!����	�4���<�5x:ݻO�rk�|�hgΉ����Ф�Il��9�P�`���.�� �3U��0�aF�`�d՚n]TnLҪi�bHk���6�A�s����P�mpS�]��vU�iYP�ݵҸ������e�:���V�I�i��5���e�2�ƃu���T�B�mQrk�m��Y۷g5JR#C\j�hM�X���u��,�ܾ��m9&8r`�'�k��<�'�8�����Ut#����m�v,6��0�e��pK��lP�/kai�Gf�]4�vL� 6��/kHa[O]�k���;����Cv�ō�Z4��Ga���R�����sy.@h˦�2�Me`d�f�l���b�L���T\�+�̜:���6�4Th^-	S+��k���xװ�A���9�ݷEO.�i����kX�YRk�:�Z�4�T�*�7M�պ�s��<!]�ƱؤJα�r�� �ȶ�s�6�(�����[�n 1�����,��o":�F���:lZ,lr�=�c��-�VΡ:���S��Q]��5	���M�����kc�!�6��fy�n;Q�h8���BЭ�K�C��[/�D��c��C�x�;u8�Ta��z���ﳹ��nwlE���6�8�];%U��N�k�gis��d�dl��a��y�y��k4��2�auI/��a��1�%R�CD���	 &��?f����`Mn������-�q��@9�w/v!��4�iu��z�Nz|����q�i�x�n�G���+XJ0�й�c�i�
�鉥�֐�T
�X˲1.8w/����&2ϊ��k8�����u�\<�N]F5�<����S���]�:�n�v�P�kh� ���=\Y�d��sժ�j ��������ٰu̝CX��j��۵�)?>_��&o�,��.����	�� _�	 �ys�?�o�f�V�δG-��H-;��g�"�х3yذuTX��&��)��g���F��{�$H���;���b�$A��+Dl\��n�u�>&�N3N���َ����ۖ��4�֘�"%�����}^(3��<��$��[� �9.��U�ɨ#u��Sa��̛��O������#�˦�y���߲?�X�C�_�3��[�qG�M]��;�m4Ph�������� �׽Z�
k���@�y�"���3����s��H��+��K��u⻮��1e+�Y�߾�ԋ#�r7y����6�$�:��x�I�g]������i�`D�sٗ9,�Q.��$_��
�ݼ�*��G_���;+��"���Đm���SŇOG(4ę5��Վ����[���l[���lI�5�ŵ7����aM���0@��"���`�ȀH�-e��h��_>n��C�[}���y�EX�u�)��ɏC����N)��Ń��Es�/%ۘ��M��s���s���Lϱ��	>t �	{�#������à�U���#k�fO�H$�n" �+� I잦�;+r�.x�բA>j��8䃓�����]'I�j%��&�z�"j�v����p�u�&� un� H#�z"�%��bu��#�l�Ye�}���[�\�[�uUGt؛u݁�8��`�k�-�hl�e�ؑ���_��������y���܄A^J��I"�z ��8�]�C"%��1o3��� ��	�lAI�V�'!�H�\��o5�e:�]��g:����ǋ�^$i�I�61�e/�ۜ�ā�25�p.âꪽ}"|H=Sq���	�[vs���h��NC�m\�q�'�o��v��%��B}�2M�>�HʂD�g.'�t��w��owν�K�3U#���
`<�0B��UB�"�|߳ĐN}�A�>x�RO)��8N�|Z9�}u�']�Ǳ�><ՏE�d �r9��ʋ��n�q^|�6���gp�"�(oUw���Ս�ܝ
�� UoC��.n"�Q#�_��MP�w)��|���s���m���,��������5����qiSFf%���qp��>z�}�`v�߾���H$�FG����X6�<� ��jm�Iv&"�;"��f>`Y�%��'�� Iy���n�7=�^��_�{�_�x/'�*��Y��N퀪3V�yd�L��%nr4�񆭏A�1���E�f써�]ށ6���#_�F������w.����֌�5e�4�f�A=�1 ��{>��؊�&�U�CV��\�j�%*u��we8�k�'&z�.KN/��g;�B h���?-������Y�ȉz����f��b Fx������
Ah` �EI�^��}�����<4�o��@��M����Wz�[�nK/���@�1I=�`���.ؒ�Ag6��Ld�*ԃ�ƺ��7or���0���G�VB{W<����Φ�n;m��� Kc�n�b�&vr�e�\�dz��a���؃R�-�a���^��F5�>&}�\�HK�᝘��v�z ��Ywם)���^DH�@��Y�� ��Յfz�x-��;6R^�7�0,���|�sa�Ǎy*އ� �id�/׬Ʀi�P k�lx�M�>� �7�{&I��)2K�$�:i5u9yB���G�w��Z��O�Y� �H=�����UU^x�Za��/d��d_:N;�)́u�ܩ�s�u�O�^^��aN��E���y0w�o{b	����n�����s˦V�x�;1[,�qc��=�O�l��ё��Z9-� %�����W���Ҳ�u�5i�������4���hc>�0a!/�G83�N�uclN�d�hƳ��L��
�&��u��Լ�Rݎ�X�v��$(�2��4�]���W��9�W�<�lP�p1�b��-��5��sV��P��[��v~�v��(�{.�꬗�AL[���X�a�8�jǭ�Q��#�P;�a*�N�nuq�u�#��ݖ�]�pg"5�b��c�n�S��[��wxzz�WT�hŮ�[��U���6u�����y)��i�@�ΌQpG��0�GC�lg�=�V���+et���<a[���'�k�<H$�n?B���v��P^{��q �}}��@��I�q��\���Z�x�U@L���������w��0U����@ �{_�D��[�Eh���Fz�����}Z�τ��F�3=	5�{�g�����A�Ɵ@@�����U]�xC��_�3�vm��N�j��K�A�xq �{#�z=�d	�~�gLb�m��r\s�;�!&I[���M>���@ �o<z��ȶfT��;7�@�'v:?��#��+;���A����E�[$��0I�0�f.5MJe�kGvV���N-��p�l���q��K��{�g�݊s���2uL@>'�z'�wf�[���ӓӃe^��'c^��.��q ��eMٚ�x'��g.�`�ֵ�Ux]�p��fY�[\{�Z��gq�#���ۺ�羏�:�=�@D���R����O��K�K���
�]I�Gр0`=P�	BE��s_-���5�d�$}��q=�S�[��upӒ	�6���%�ݜ�%�P;3pB�I`��̋�Qڑ�m��ދ��#<����@>�s�Kz�V���*��5�l�"/Mh"jn,M��%C�5 �����f_��E�1U����0}��L�dK�W�䵘����c�[:��,E�pO�^LG�$[�����gt�/�:ݱ�+���_����LZ��a�f�J��ln��V�D�Κf��B5� S8��)�dmH�z��Q�k���M�u�=6�������=LTX��[Gf�7�N��y�ǁ3$��f�3'�2sW\�!z<�:Eت&�zs�H8��`^�3cwDx�ޣ���Y <h�$X�X�N���k�ُ��$��R�O�k�v�NUe;�iyHE��v��T� �u����FiG����n��.?s�9�{7�O�]W2�����w�ߕ�su«���`PҢTg;�t�m�f���az��{d�{ݕ�̖��,	h��T*w/Ywv|lUm�	$m�<H$�ѳ���I��R�cį\r�!�d�ú
��_�O[Żѻ�t5��hm���7��`ϗ��k� ��y��u��V/@��)��p�aج%�lVV�]���E.P� 4U^�攉��8)9,�
�'��`����Q�A�nkϯ��y*7d���j�,�m��;Y� w�b�LR�E.��o�e�����ZPC�Z7��q�dI7�� �I��`�&2{~5�	�����3�p�Ϳ\>�-M� Y���#;�G��z�Hm�xp$Tz�,�;:FQ��}�=��.� ���A$��x���
qy�m�U����Az�K\1qy�IR7�#�{�eX=��)�-Ր m7&r����}�^��/I޳���N����Q(�|V'����1J�������o��ka�!���ŗ����-�����{����i�sd�N6�//� 	6�g���q7Yc�?9��Ė!��$��K��u;����è��d���l��3�S�g6`����]k4�D�'�)�\S��x��{�x��� 0�7����a^n��$�M�s$��0I�r�y��R�	\0�`k�>�^�K�$�@�ۈ8Y��x��>`�銲U������*$`�:(9t�'Ǯ� �%��'���ܮ�S��x���n��jȇ�^�%ѽ���	6#��fp�3�Ϋ#ra�0����£�m�kˑ$�b_r}>'7�!�Ѱ�Vo����~�L�X��x�;vFh�ǀ	3�ߞ�t�\�1�k�O���<I#��F�K4�.�؃��q�0$,��\אv���v�FyL~}����ڥ5$�_B������4�e�cUܗU���3j� .���x��<�q}�y_{�7��o*��ȩ[I��A��mlˬ��`ʖ���3REoTU�ϊ|���2Yӡ�?eW�A�K��V��.�s=��787&�:`�0�d�d���r/�uq!�F�<q��w��8�q�щrIM��C�5��Yu�f��L��7:JZ@�b<��J�l6�0[�`�.t�$�+U;Pī���̭ɣ<<�gVmiY�rv&�:�ej�4�c<�`j��g��s�T��N�Z���X$|�tld��U�J���'�q�V
��)]٪[�wa~�z��?n��ϋ�5���o �wdG���Cv�>�3�{s���^(x�͹�>�����tz��� �|�QMU�Vj*��b����$ov�Wv�u"��-�a�z�����	3�%�����A�9��V����{"� ���A��d	`AB{zb	�{6h`�:(9t�(��Np��8	��x'�x�<�W�˛�e��p�u�|H��� �l�	3��ܲs2c�b	 �e�c�j�W&.��T�A$���A[�"���g�߬9�a��ki��4�����1՞&��M���:SI4v�iTl]����}>�N��=��u������>C�'����n؀vf�y�)���xߕ��n}��>^��������,���w^=Y*r�$@��Fz��`L32�m���7�	�A���gb��e���Rݨ}�[�Z��Pbĳ<6R`�"�� �x�G��A�5�����_'�$>{����� Gz<��M'�kg֙{O�c�,,]!@����I<���<�����rl{��#����؃>A�=�Nߘ$��(<�ɇYW��;���<� H l[�&��ހi�j!�Ò.�-��7�����E.�D�k���H	UQ�&��X�wD�L� Cx޷8�z;�A8]8������ ���&,']��-�k��[}�(�۶(��=u�NK�:.�xn|��@h���L䳻�3��z��$/$z�b
�D����c1���B�Ay��M@H�$w'���Af��|���ӓ~1]� �GnW��r+�ZZ�A$�ET\D�#խ�<O��)�k-ۚ	�dHT�J�N�*�v'�	 ��Y�M��LM��������U��7?hWҬ��ph����������"��=J���a��gNc�wf>�Q�4�
����� ����w�R�]�g�ʥ�N��|O�l��}��oby��z=���wz�����.H<���R������j*�W_���g�U�/e�w`��9=	�}��9�q��M�-��ʼ����]�I�䧧��=��o���6��n*^ei1�4�\f<��Mh��	�^���O�^�~��9�E6�(��=���4��_��=Io�����>�����Iwf{}zz-�V�	�����W�ul��לW<F�#���7��'���_�c�v�6vw�n"��w���bg�7dQ���ϻ.���3�����7��b�b9���˗�����.?���E甪�O��6�����q,.���)S�Y2��)a�P�]��_|��YJ�s���U������>��;�K����УX��C<;*��薐�KڇG(I����L��`��-zX��k����c���{���?-�v��p��7�'~��o�-K�"��\�d=�b%h�rf�1�I3k���!=��ܬ�=�U�=�g)%�˓���<T�j >��w֪6KJ��fܠ4g�bS}��%��.B�:qF��8oh羝��/W����̍niu9W�&W��y8�=uy&�ٜ�[��?B�r#���K@d������"&��o�M����<�l\�:�oNk�t�Y�ޘ�hl�P���d+,�ed(^�	���_���x�wtոy��)"!G
�Y�� ��"T���\�Ի��������==���۷��:��q�jF��!�RB0���YQ�,�S�eE5J�t�|������۷oO<xr�
���B`�O�K"�V#ƵE�Z�	�EUi��pϳ�r>>1���|v�۷���!ʢrT1�2c&l�*��`�L��dF��ESZ��&��W8�EG�!0�1+��X&8�-Ɉ$b
�"2��]ff�Ÿ�9���l�0�HQ��&�$�$UI
�r��)�,�&�L	c�R3/#{=BԖ�olf/��`����>�Q����u��1�_&A��l����m��Y"N0�d���q5c ��\pEB�-��eĖW,�㊖���WUWA�ԁ�ܢ��JNI�]��"�
�DB29Id\E�0�� �1P�;���?(��׼vI���0O��9X���!ӯ'�?k��1�+��;s��-��Ê��^o��u�+��E��y��&Zf^A=^dS��y��~DA��x񮸍���"Rۑ�M�m�G�vtAʋR��]��%��~��F�v�����T[��s�u��ȸ齧"�e��d�PuY�0�΋.��x�ڈ7�`R�����]�3�h3�1��]��O��x� ����p�h���� ��*�<��wa]9}n�	-���PI��� �1��ڂ�;r��wS�>�4 �y��NL�yY��$u�<~Y��jU]��� �5^2�˖s�$ln�f)�o�$�dἂ��X���<9���D�n�d0 �6��x����{���x��a�A����&�<�õ�������T7&<��x>�����Q<���� po7<9���\�]v��TC��H0Jx �x�	��P	a�\,�)�t�ʨ}q �|~���|�q�ɘ>�e�e��Q�|Hܼ��O>���1��T��<�/���p�j�q4�@cx3�{7��=�W�m��Ŧ�K��5[i�/��۵)��a�U-�A�$���Ă5� ;�ڎ9���w-��H�́x�
f�Ν×OEs�z7ro��[y�ֺ� �ݚ��|���u@$��p�� $ ��@A���i�w����b<H$7���I^��9��YN|E��o4xN�t�"�s��"Kw�ܻ�`{�"Ss��/W�ܱ8�>dC�tn<��(���'�����T$9����}���+f��\�U]	'�]��m�]�u~U��"do��]����4�9�,Ü�k����.�[��[��u}�׹��ǱU����Z�h�q��}���5o]���ȟ�^����<s���=p|b��$1OGf�ݙ��<������f��"�-�*����'���8��v�^���5e���u����+�X�.�ϲm��C�Q/9�7`�4&;�o���� ��ӂ''Кx�up	�����[�[�i�L�Ís\@�q�����N2�5O7��c��й��Ϻ�iJ�0�{gmjA�F飭�Y�t2ӓ6�r��^��η-y�� :�6z��y����֚���q�.&���:�Z�h�{CMeʔkj�	���0���d�j;1������+(ٌq����sq$
�@ƽ�B&��m���H-X��ah����0[�,ē�@��"]��`����EG�m��i�"�/����H���K��'�a ��+}h0��O�ră�4M�:w]=� f�D/��h��=�����^�y�_�"	 ��.�O�p�J�]�`�'p�0;�E,����DJ����ޏA'ČQ��Ws�Zz��ӎ	-�#�����wN�����mc������ ꑙȶq����P�ނI����H�s�?>���#�=}��s��k- d*�Ea�#��h�.Қf�����O�~��XK��.�Y����p��y,~�J�����=%�w<;+�A#��0���C�L�����<C�'z��������hvWAq^����9�/'��Ў�<-�� /�R=g�w�_{O9l���x���SZ.�3�h޻�rh۳]��a=$ @I�~�O������}F3�W����s���C�'[��@$���E��x-~����
O��H'3z/�g͒g˜'Nዧ�@�=t����6�.14��G���D��~��f�����A!�u��Z"���N�33L�;�D� Tg/;s�kf��A�,�Y����=��=�/w��N0�����[C�m7�;A��!/�+���u�,ɷ;v�bf�U�����*?��L���_?~�c�|s�!��D���6������3!t&�U�G��H���҃"�Ip��D���g��朘SK[Zx���Uv<x��zy�M�s���B=z;[ͫ�b]���T���KƱ� ��l�]��g��֍s幐�!�Ol�7�\3�=��$##W��0��e3]=AW��[�C1��m�E9�eM/m���K�ʹ;�&�Y>�$`?�zڿ6��ǉ#>���W�(�$]3�=�h���υ���C� H���O�'��$z�ynj��y��4��z."�!q�:w]<�m�z'�eoCMUw=Q.�'�t�z'v��@Smb\�r�r��b��,�Ӥ!;$��m�..��m�
��j�CjZ�d��ﯲ��:gb����3�q��	'�����`1�%�Z��Ah��.4��EzQ��Y>�;��]�m�n8r}�6؅�EU��<�A>'"����D�-ܣ�z����.U3�UM�%u@,�3e\��ȳ�\-�vg` �Ү�1G��X+!�y�p��x�$�呝 Ex����<H�5��$�,���޻�]�rU���y �tDA��Q�I��X�ztǁ�-0.�d�۴�<tbvs��{9W�f��<_og���{��"s&�J���������xV��Ã1�`2%|d��<�^l�8UM]腃�z��ҏ__�;��R��*b$���A��u����K�G���?���MK$�xn:�l-���3�$]�jYEТ��,&qT�a��e>�tnOÊ��H���D�Owt@1vn�rZv��|�s� ����D� ��p7�3�fMv�`G����h׮˘H�ƾ�H'�{���}Տ�)�7?��_��I%������Pxƫ^�q �r��-����� ���H9��<��n�W��"��U՞H�,�3�6z1ow\����no(� ���A �W_?��y�ol���tCy ݯ�#|�;lhȲ.����#|���n��t���t�4��`]��$��΀!�`�dZ�p��w����b_l��h(��{$�L��_��s���v��B��ˠ�ٻ��Q�t]"��_`�_���i��*���̮�[��\��ɝ�tFq����5|�5��h]�����1����.C�;�{�䬺��f�][RP��Lb��}�b�㷊�st-v�s�bε��S�M����E�rs6�]�sr�'�☤��!��1\j�AAhuF�v�bH�ݶ����u/;n]�fZ�rP㸸9��`�94!�7˭�3S�v܁�=�f �ZcX�n3���q�9��c��t�ŧRɜ���׌u��s�r稗FU��s���>an�ѕ��t��I���ܿϼ������CT"I3�� ����fɈu����x���v���۴�:d�1t��Ɯ�w�(�;͐�mcm/	�݈7�y���L-�<z�Ή��d戽�yٜ&b�*���	�$Sm�����z2��{��{��|}���}>��TAf�3���h`�seq�"�"��$��<�H�N�	:�=�VzT�x
�����A7\Q,��$�U���@�+��l�Ǩ�.�#�b �H8�q����y�..�bl���A/Q��rPٓ��=ۢ�qi���>�4�BoMb��b8�%NU�9E�fd�]ӗQ%y"�w��[�`z�Μ��<-��f̈�$=�<�ܰ{<PN�	A��@瘨�w�2�䱳��*�`swD�Gq�P&wP��?`��ѻ���j|o�?r�sk`% �F�,X7�픇H����c �+��|1�d$cﵽ|�P'�j�@�̍��_8v�u�p$O�l�;�t��9t�FR͋�3䁨Y��Vn���~���I/���vr�b�'�V��ȇfp��@>�gR�|��ޣ�D��5 G��x�R׊
�A>`��5������Duȣ��F�/�kbۆd�͞ggwA��J�^�@$��<$^}��P6-^����j� � ��;�纕t�{��BgɃ)H;8Ğ}�l�F�"y��n׭���M�4*�؛��-����d'p�8]�3���|_!��+ݽ � ע�Ί{���M�V($Lmpt�f,��1�/~��a!�u/;6"�A�!���\�	�f�|�n����u+��۳�"'��g�	��(<��U*�W�vf�W�E^)��׍UZ�#�,M��n�3�{8e;ᩒ Y�T�2�CS�{=7˻P���@��&׼��Yx����"Cɷ����������  +;��{�3Ҷ
���_הg]��`����P5�S�s�
u^��@�.��1�b����%�,���!%qr0I=�t���t�`���I��9�� $�1����T���� ��F������H&��u�A�ju�X�뿦�'	>�4���E�`����Y�q�	�W�W��+wV�GTl]�ŝ���6�ˬ��7p�]�����%�I�΍��\.٨M �����x7����[)��.��WDs���2=�+rX��I�3{w������� ��^%y�Z��.r�I;3��L̙�!L�w� �	=q���,��:�ߜ���B�m�x�v3�`��@�x����ݞ�S��'g��!5c� �1����m��]�E��'��P�n����D�2�=͸ ��=�Λ���!u��� ����p���z����I�k�Y���
��Wַ�\R�1 �%[5�|���<�Γ�w-"�c���d�¡}�y��>�NK����؂|I��q �v�PK*ޤ��j�s"���S���c���걣�g��{I>���]M��L��-������`�K��Ȁc�n؂$������,24�ߧ�}*<F�d�f ���2wwA�<,��}>`ji�T������9�b']w(+�Cr1�*���/�J�L��1p�^/���%���r�����̉����������n�+�9\�.�3�!Md�D��#�Cji�P�W�x�F��$�P݊ '�䯟�@���K�����tLC�Fl��wrJb�PI��x ���|�]x���0���-���R	3��=�+N�B!�_�H���½��	=�
��3�׼l�ݨo����.x�w&�j{�CݨN~���oqy�{)qwW��Ɵ�q�a��ٸV��D��-��z��-�7�,E������ܼ8���x>�z����۾��%�q����}xcr�zo3�Z���n{ϳĪw`���h�]�!�p�������4��:��,�z#膞��3V,���>�'�pfwq�g����S4Ѡ���o`�#^�\�<ݧ9J��w���t�������2�`�>������9�¯����4��qi{��j0nƁ���i0���p85⼯��u�ٞ�8�n�O<���ù��[�.���#A"���f{J��3q�a��d���{�kv��Ij�n�.=Ob1;�.�1��~D��bӽ�s�۾.VL��yQ�oK9ć���jF�`��~b:|sڒ\Rօ��{�T�ܛ!������&o��h�^�=�j;��>(��ݎޚ�P^Lќǻ��5��u;&�{�srvÂb�r	 �$�w�z#�I>С�.���~��k��)n��ɹ1C�QNW��X���z��9���{���{O-���x{�xf�8Ǎ�(W�G�R����<���TX���,�V7h�b(w�ݎ,Μ��>���/>�x�;(|l���w�����%{Z��w	!v������=�㻋���r��0tO�Pd洿��q 3Hc��f����p���` C[>M��.�$����F�JVU�Y;|묯S��Q�H�1GS�*"w}�.%����w��4'����<4�4�va�(�\�6MM|Np�ʜ��u�r��b>����n��{��x��f��Ɏw��	?\���6����1����ʄcf�<N���<���J~�`o���[r�.8��Yd��ϼf�d�yiP�{��YV���"�	YR(�U5:H��#0����;�r1���O�q�۷nޞ<w�Jj:��"=$��(���[)�L��&��I��v!�&��D�%kT��x��>>1�ǧ�:t��s>3������W� ���ؚG�ri�����m��h"%A���Q(�]�]Ysr��Ƿ�<x�㎝:t���Bn�bs��ZJ5Ta$�l�i#R+��� �0��DVr[�[�0H�cY�D+�.�pqERH �qȩd�**Db�b*��V:R9#6��&��+dŌ�b�"F"*�̌`��F�$�V؛mU9-�1�VHsnAJ���J��sw@A�HjZ�u%��ݵ"E4b6O�Z���2�����"�����5�f�
�`�Eq!�H$f8�`�D�G*A}p��"��Eu
*��!k�*��@�qb��gRm���F �r���&!�k!�j#rޣ�zJ�=V,u���E�1�������M��)f#0I�f�hk3Ay�,;j�[]llb�x�̓3y{���GL��u���.�Ƈ�¬��`E��m�x�^���;�`9���=l�g���+�ݘP�ò � ,���%1����*n�8��Cln;��dmؗ4��a#���A3��,Wfo<<̡�3�+���3Ԩ�8��a���
�cb=me4�Z�fїpPL2J؍�l��dy��}��C��%,�=�h�
���kt�]��&)R�JD� �hU{M.#��m�6���$�XٙUې��G:��8h,NWY[P��Q����kq�V�nK��\m�X���W�
�%�4�1e�E��l�$]LMept����i)e.��JF�hnמ^\�=�\Z0�r��c��؞�n4nŹ'��x���;7f��5��X<�a��:1�m��2��'f�xI�y6�Svң�;
���t⸉51\��r��t\ݹL�n�6�<����>��q�$ez����&΀���lЃt��������ΦM��9��d::�ZsjN�0sh��S1D5o@�k��9N)�*z��#�����c�m�X��N�J��,�cp͵�-�	G��q�Y�f:ɕ	i���ޱ�*�!��2�3�+���e�б��F�K])1�%)�"�/8���:�J�3�ܯ8��h�(L�C��jPT�X@&�mccv�jDM)H��T�r�3-u��\�{[��ڑ�Y���1���tt��Y��6#^֠J:��
@�Kɰ�Q��mmЎ��c��[���,7���뎔xx�vE��]g/U�����u6��0R�芳G��#Em������1̗x�WT�j�l򮸹��Ȗ0X�
�I��JF�Y�7���
�u�/�v�����4�o]1��%ǝ<e�R]u�G��4nU�=63�X�Z2�\&H�Hŭ0/�2��JX�4��K�Ї2�J��;���.��P�����4g`���Ό�n(�ݘǊ|�$�q�8]ݍL���8�=�;{���͍��6�1,���Ό4��j̮�a�1�	��½�;3��_�ž� �گD��jVr�A���ʺ]�p����\��Gz�I�v0UA��D�m�{{$�d{u۷ ��I�k�!����G��������4g�z͠[\�N��<
*�>Ag>?��t١-���i���HBC��^=�`9���f���6�)1p�%�z]p�vEޅ����I9]� �ONwK�_;�v;\�쬼]E���je�|Myu5��	>�X��$�8ݪ=�,�؂H��p"Ii�>T�������S֭�5����g.�t8`��n�7Izۜ�������
)�jXh�O����|Pvw$�~㖢�1Vn8��Cg�`7Uw��#�ͺˡA>$���#�3��_�Š_�쨈Wn׍�=O.�>F�^�����}���tYX���;;��{f{j��ըS�vN���(�OV�����b̫��q���������t<P�u^}� �^G���/�� �O�#�1���!����r�DH�3��.�Æ
Wz\g�/~@�� ��%�7�ƒN3]����$��#ĀI�ہ]�2Kr!çr}B%sƝ�;:�v�ӏ��@��� �7r--ـ/���i)��$���}�g��@�+�Q�r�ˏy�T�W��L�������x�{
�P	���1�tm�9� �v�ir�#��g*F�IMV$Ql�����0ir�a��K-�V���Q���*Oߍ���9���NCw(�q�_��dL�|I��A�z'��;;:.�U]�n@b>�`-R�Æ�n�Ky gv���[yA"<�G�T����g}X*��,���ZEiׂL�� �GG+����p���a����є%yP�n��^�ɗ�������ɓ��Yu_t���81��n��w�*��N���H0R��[�H$�o�B�_C}�o.ek�9w%���>���/?,m�$�_DA9x��y��Vb�Yʼ6I��xܒD�t��N�<����ا�-̗��y�	������=H'�|��g;�<i�YK��׿�A�bz׶���MM�E�)u�RS��^.:�I����Z+�s�����>�+�9c��b���g�<˥\�$���׳��]�-�� L��� �0�	��\���&"���=��y���[;����q֮�Z�}$�f�W�D���Nzg��9N�˷ ��w���-��~�vb.�<�+GtKͻUEz�i!d(�$�E�tA7�']7�r�LZD�ʊff۸���Ag]P��fo<�v{j�dD�m��L�x���J�&�҉2�	����O&��)֝&�k��t�|�ny�Цq^!���<�/`�}�G��(ݟ��-`�0tM�\���ɯ9�b�9g���޹�	���CК��Rϭ*����R�����>��A�'����!�_��\_�t)��in��w�r�~q�ܷut[�|��/f�U�g����>��c9�{ॕ�11�U��>��qɶ�Vt�¡��#�6�I�kR���]Ӳ�Gc�B��U�1=}�֛RO�#�2 �A�ΏGx�c�sR�� ��u~&3��I�3?�S#��]2	!3w" >$��m�f݇���<�x�v�:�Hٮ�ANߒr�]ݓL�9S�5�Vdm�����\?��K����{�o5���vC8�����Ȩ�	�7a�"���v�GZ�#�cz<�,���>�w��s�A ��Y�N��h6;c�s�n��g��Y���ٔ�ɐ�f\����sw��_I������?4�Up�߀<��~��|��������jg�!�ɴ`k��*��S����t�}���Xl3od�,��'��w��,d1�&��낳�(	Qs�t�ª��1�z�X�C���6!�3K��32,&�	���J�Z�7����y��ɈVmcnP�!j�3��5n�݋c��Vx�rq��v��x穏e����\c�z\�X�Wq�F�����mNꌠ�Mq�2�bۮ\�d9�e�7<�M{9,��9�f5!��
������ϾNɊr��|۵M1 ���(�^<Z���f�ȇ�#�t���� �����$F]�.�C̀�L�0�lc�������H� �U�z�W4N@��͑:z�f�Ԕ�\�N]�3�X���@�{��B	��˃!uLz#ǸW����O��cA>���~�������ȫ�Q䏏�߰�u��dI���D_?AF�v%�W�h�k�6Og�r���٨I���Mwc���#,@��4fDA(����^�1���{ܵo���J���C3��cs���GF%[l�bi����z��[`ю��ZB��;��v�A�C�7u�-�I&�z �os�3:�����:�Ɉ�^��I�3�ݙ�t�W^}�&'2����`Ʃ�ϧ�%y�T$ӑ:�m�N<�]��6́�6��R�2�wZ`�xܻއ���c����W��7�wRM�>� Ȍϝo\~6��(�$����%�Y�ت[���ؗg!�L�ݏ1 ��|�I'j�,2v���;flr<[a�TIW� _�M�	<䳰v�/���_R��k�I�x'���<��4�����D3�Ea$�ns�A;38pB�穹��@�UM�fҙ˫2˱@$�D�t@5��+n��5mna6C�ζr�̰9l[��fY��W���*:�]�t��<u�`���d�aw�����N�ӷq�U0�׸�H� ���������`vv���c=(5�����r�;��i
쨂i:/Ú6��+�-���
|�[=�M�7]�K[�cJ�cӦ0Ӳd]��`�����!O��txA$��х��#��:�Ҫ�mX�$D�_)F��=۬G�p�L��&0��I����!��0��]��br������30���x�!"��u�!'���̈́	;��7]�g��g!�MT���X�NW��v�x$Iی�!��_ysLEWv��ٺ}��PuHH���S �Nߧ�O���W��jo[" ����r;��ޥ�8�-|�����8Τ����6��)������n ��+�M�Kٹ4��stbQbzk��38pB����]}>H�������~5<˛�=I���$�Iɱ�<��ӧt�K�bz�13���/|�]3n$�z��	�y �rrM��n�N��=��9)"����(����v�<Z�ϠA� ܪ�{�����:;�+#���6[�G�U�N�"���5���謊j�{n�A�'%v�!vtc����M�\���cCޯ�{�o�W��Wg�/�+�ĿM�ߛiM��_�+��L,(��ڡ}��;84��gm)?���\L@G��UƼ~ܰL�!ӂ��=����bH5w���'x�Ҍ޿<3�$�<DҪ�Gn�@5�I����	PI*ԼT�4�ue� �pGM�dl����ʰ�<�XRlFϿm���|��lC���� A�rU�0��"��#��{����Sb}�>d�ʮP	鮴�HN��8!��SU� �k;+a��d���g��%��N�tA,��t���|��zf���w�;�j�wRж�>#5�-J��=vKy"rZ�A �������4][�HA�]�P=�P3�pR�"H��vWZ�	�q�_�<���H"��C�p�~��S�B=���i<X&��Y>Etz'{2wz���n�aG������Q�m��1G"�\@��BE�fz�X2i���^n��2�m�vؽ���r��T�#�f��)��� ���y���C�-��w�Z%LA�T��t�N�e�XݛI����A1�1��۾����Wi���l�ugK2JƑ�N�^�,��4�9�[uq�ϒ�!�FSL�q��ۊ�����0�I�s<�泮�ێ�R-�*�`�q6ݪ����dp�N��[`'`���F��h��������Oc�����s��C�0읻Ƕ�CY��;f�z�>��l��ڈ���K����mt�����5�(�M�1{hT�솮�&�k�.f�]-�v��{�.�g!��2�a����xn;�������c��@@ �:� �+D.vg	Ó#e����!D��CM�[X��}=������8�TKmO'�I�I1�m�B���f��a!;�;9%����@�$	)�נA�*� �[w��<D�eZ�A3�� ��Ky� [�L�߻x��Oe2ͣ��X����"��"'�|Sθ�D���.Kyl6�q�Yu⹲byn��A;�KәWTA^KG�z韤5��p���k�&�/#�:����D��eN�`����_s���z���4����^ ר6�{m�틤k��ؖ�J�B�����/��%f�{�\T@$y�c�I t�qh�j�;��&:�z D͙f��20NK���"9�>/"��,[�Q�և�y0�W,�+�X#-����X�*�F����!�㫋���#]�:)�|��Oj�s�WU�6�DT�sa�_|<H��$}�߶>$�9���$쯟�$��zv�����to�˳��A��2T��#� "�Pѹ��u��J�`G�:�� �vu��;I�y;�;9%��^�ލk���7����uO���Ϥ@�{y�f�ຶ������u�_�ܻ:gN�]�e|H�1�ܸ0r^�7/[
�^W�Aݾi<�n~��.O|��/���JK~�ң�[�ͩe��e��5�]���Ջ�����^��G[n���uޠE�M�Ά%x�����<�'Zju୅8N=�Cx��ը]:;B3�&7�\n�������uT�εo��A>�k� ��oD]�ݥ{gj�2�����(i.\�g!����_�U}�#Ĕ<����<��e|%��
c�(mƱ�C}V!݉��
]�d�����;׶��%X�X}��^z=6o�y���\�nK�P�������]<HY���� ��D�����=ޞ]������y�O��Q��&���o� ��8��뛄N\�r�Q�Lyq�إ#)���;��N���y�<t�i�N-�;_���_邗���/E�E��^{����U�{�wm�O1�{GM/gWn���Ŋd���ξ\7r�v8{d/Cf���L��.�G��;@��ٽ����㣛ĉ~��3�]�'�5���G��]�,���B~�:nѽ�v/Bi<�	�>o�_�=�ބ�ɘ��OU:��՚��ҝ��H�C?P,�dL"�X<�o��yq�{�3�4��4�A��q������ܻ�6G�7��a��8'��� ��ː��<��̽�|:&��ǝJ���R��������tI��������%JvM#��`�G�yg_f�>�\4ػKg��V�m%�g�'��c���s�9�?j�.:$ |���!�Q)᏷wV{�j]��;=�{6 pr�wH}��x}I۷�E���-���ދG��C(v�FC���ؼ}0���y���0�[b������?~�iU��/�^���o�C4(���bY毹��y�x��罞��@�b�
iQ���!�iZ6)�8�8�@�8�}�i�F�c9dG|Zdx�l
�Y�orm�?G��
��^���?�!s��Ltg9�^u��=$H�W*�-YY�82J�K��~n"�
��E_���$�N��Ƕ1����:t���z6T��㓈Aa A�IGv������H�r,�!�1Z�-�w�պ��.�|c��:t���s��OIV�S#�+���`sa���X"��b����:����V%�WAT~Ό��q�zz{||t�ӧO��#��{�r"�Ԁ���.D�c��XՄq�'��U�8�1D�B��<�R�!� �v��N��-*��&kQU�` �kAW-�DE�����Y$��9�"b*��"V������B���m���!�6m$����p/M��������hHĶ��-��q1�(�ۑ��$�\��`�Ԃ.(��$l���㈎��>��GTEDJ��d ��#��E� �#l0Ԃ�습��*�$Q�W+dk��#�� ��E1qq�L]C���\Q�R#����D�*�b8�rE\UDc�PqnĤAܨ\)��I5p~A�`�y�~Q��TOv��}�0x�L�3j��wK�9�[V�t'�Kk�$�n<��K6hͰ�H+�F-�!���7ɝ���*�b� In�yzz��s,��%��
���	�}Έ{nk���C�K�M.�7TT݁훬l��M���b�/�id�ָZ.�8	�v�-bܻ:gN�w�)�<n���Dn�=x��2#�XZ�;Y��j<H'՝������	6����g��Y��9�z6��0 ������#�vΘ����m��ul�(8t�ę��UWG���@�6��E�5,1���Cvc�����?��>���vr�vj��38��Y�ߎ�S�-�~,7�>ק�b�ƬE���%�6]�c�Ieut��G�o
�ż̙;Bk4<���A�������D4^Hw��T�c%WR�.�B�Qa����x'\�[�91t�2e�b$|k��\	ї*�-�>H��DIk��}n0c.�_nLn��dŁfPS2wwJ��B�uV�mmi��S�ê�g�nxf@L��ny��a�fwN�Ah�b� ��20�Іy�����/t�["�z#Đ�x�=�\��wr���;N��j�A��+5��_��F O��xߢ=H��~0	���.��Q�1�&��� �8&�;_��z�+$cq��	 ���-Me��$�~��嫚RA\����;f{��+�1�f�,	17q �zk1�|H��3q���AF�{�;PH�[��-2�����!���x�:;�'aXٕ�Dl@���v]���t@*N��͂��1���d�\�t\�-XiS��Z.�'�s0f�w9m12�,�ŭ	��t�����s ��<���2
pd����0
2�� ��"�w��,����#�BN�����0�,�%�q�w+Xo�2�>q�Xǈ��q)71�]v����.�uq%͐N83ۮs�� /lڮݞ{�E��v-�Z`�YC�� ��aWb$�u��7Y-͌p:��A��4��X	c���γ:�qlY�Wj�K�!�Ї�o7Y���֎�d#�V�c\u��m���ؽsvQn������uU�w�A�,]=�'�x��T)fnP\�������_��H<��,H��ɪ�c���ހ�;s�<`3�:�e�lS�@ �{~0	oL������-4D>tj�4�y"u�⺷�ۓ0$S��Gns���f-ڞ������A�p �^�2r��3�We��/R�$�ǀA=���[2dU�&ߛ�x�?���5�� �i��B3�mC����8���"1{� �o!�y"	�Έ'�ϐcxNW����^,L;�$Em��N]&w]Ƿ���%�bN�[����@C���HD�lȂA'[:s�o��}��H�m�c1u 8'�!o���u�\��p��������m����u�35~���\"{�U�<y"�9��U���YTQ�ݺ*���$��؋�>�0�$���$M5�k���l$�ѕ"꿻�R<�v=��T���ܖS�&-M����ա�yt*�pd9�e�H��u��%mti��������f}�4p[�l�Y�fވ �|� Н�۸DW�[,�L)TҦ��靐-y�	$�ݼx���yy�q��Wi�I7�� :�� �N�2r��;�i�kݒ�ٱq�T ��[�E�<)�y��Ǣ"/���0��sLZ�S��x��Uo� �8&T<��X �H�n�O��l�뮡�	ܩ��|I挏@'#���oמ�y��?N/,����YrZ�k��-ǣ�>؜�QMWJ�2�3,���_�;l���lT$���J� g�^E��V%����TK�x_�"VGB���Wd�#��%�9h`�styo�I��f��X�p�	$�:�Ϣ	'�<�`�y�����e(����P��\�D�8bDS��j���)��f�:]<����q&�"�rn�����>3cx��nã��L[0�#RL�R4`<W���f"�U�z�����l\<���>#�6x��~"Ϊa�I����}�gN��x��r�^���$x��}"<lE�"��lC�}>�7��8wtΝKz�\�@D��ǃ�F���C�����y7��xo���{0I��x�-U�f��U�#�76�up-�p���;�����6g��n�Շ��`,�81�ApO(v�n;ҁ �;i�{w��Ѯ�����{����dH����F�nP5�:wI����}u5�fFSB)P�]�����*i��$�ovDo���J�k���jjD�$�`4	�!�N���g���w�H"6�_�{~��>9�rq��I]�z\� ��8bEU�c�5�E���<O�m5��s/� +���'�����_C>��w �xxy{��B�2{�}Wx�"�����V���t<��Ԭ��2��=��>θ߽m���{�e�4<�3�S,(�ˑ�����x�KA��S�wdE����������u�B�{ @ �fD�dt	����9�:��	t��Ń m��M��{I']�����fx�a�]4�R2��5�Ͽ}�����Åp�v�� ��9��w#��u�v���S��>39��D]�D O�lط!�2��|y���_˩�0imfن]}��[�	�͏Aꎈ����(�qXz+t�1UP40�wL�3�w��gc�	 Q=��3���G�� I܎��l�@�r���@�5N�x�X���E�k�Vv=�$����I�]jvN��֍�gN�O���2���:��o@����y��5�ڌ��v�w	$}����Æ)���1̮�b飶c�79yn�^�ű���c ��Eݼ�wy{�p��}qG����|1@�v���R�B@�`�/i0-�,7@�<�UF�S�XAѶ�p_�H�|��Wd��T5�y��R�u�M1b\���6�R0�`$��j)��l��t;�ju�9�����nk$Rcu�{� a{l�ہ�NS37��e��v�݋��l��{Q�%ħ4��^Ż=1�O]�ƭ�ۂ{e�-���%=��[uf���TQq�t`ˋm����4�l�7h]��T
��m��i�v�����Z�x�wg�s�I6]��j�c}���?ۦ���~���I<�p �<�'����3u�03]�y��J��A�q$�[c2��݃5P5�*i.�;�ӭ�7$o�$s�D����u�n/5�\WL�W��A��c�Pp�҇{;oK������7���ݷk��m���O��x�#%����4�N�&r�{�c7"R�va�����k�,��^�uv�fI�e�v��<Q��>����I!��R.�x�-��`�>`�7��&�7��O;v���b)��G��5F�H ��nY�mx�1�1(9�v,���Jk(��5RlG￠�I��C{����'e�	��l@���^%L������|NCg(<���S��wtL��O��Ǣu����w��<��@��f��i-��p�e�� :����Λp4�a%��r�%�4]�p�)�T��2��BS�TrAE�UM�@����~��H�*� ��ؓ'@��j�]�fC;�ou��2��݃5��lA]� �YwNJ���,�� uX���� �0-�%!(w���,jڌ��g7<h�-���vs��/A��#���O!�_���ǙR9Pqr��س���I&������Ѯ�^Ya��QU�A"��'�I7��������֔����x݆���F�A:̮6c���0�fY�H�V��G��~�_٬��?~*��>$�ǀ��}���q��b1�	��@$�s�L^#�o/L�i؃�d��A���7oV�0&=��	$���F��ca[�U�(%��V�a��w.�j}�|&ǒ7����n[en�(���ǉ�s�pnS��9��7�o�!���{ʸ�o]�=����N�-{v�~�X*y��=��]�}�¹4�$2� x���wVRInN�2	݊wd�b�˜h�̮�ˋ�~3���A5�м`��K#�8��>A�|x=�������.(v�tg�<X孕�vx�n�U�7=>3�>@.y����n�flB�	�� ���O�`���[C([R��)�-�5�����f]n�j^E:���N���;v�Q� Aꍈ �һ����q|��ש��=t� H'�r4��`I��Lm�t��5ٙU���&��T��u�x�M�tG���+mO)���f�c:���y�d$7�1[�-z���by#̷�e�,��[]z��A �_�A ��O����cE˹vt@��S�4qY��N�K�nnǠ�J�^����Ls�]Qu)�����^�i���U3�s�,��G�-�5��2jX[��~�k��}|�1��~.���JE�政C��W	���$9l@��<8+��{��uFbK�)ݐf��EC|go�<n�:C��g�6�ٓ�GR�B��蓎�T��V	��A�)N)IBYA��i�!|��
Qde��T�уn�u�����mi��z��#�\�;q[�ꕻ��=�� ynd�va~���}Y�$�|PM�A\���vt]�f:: w� �295��W�=�'f��x�۝'�Qq��z�]+�m��7�^)V�7x�Eݛ0��q�2�	�{0F�u3��LL]��#�H��{q䚘	�v$�"dj�ܔ�Lm+�J!���Q�Wn�/����n�Ѡ�U-$G��Z��"�;:%��v�$�],u�b����o��7ޅ�|��H���@8t[�!ٟz��E�¨t���n绉ɽuC��jCc>�/��8�&�u��w��;��,Ƹ�2���ӽ���������/�^��s�N���{�V��f�|x����;��ؖ2�k��{<��ܕ38ɡ���{n���O��U�S1 *����O^
L�ּ�g��V��;����5��Nm]��w���t�Ӛ1���R��Ÿ�Aw�s�q�Kɫ�F�Gq�/���i��M�����/w�y�C=��Wt�;���nxqR�C��.����N��f,�G�t�7�}�ǆ�oS�|X�{	��G�ޣi���w7��a��C9��Oۆ���k��)n�֮/h6��{v�>Lf�������]gh!�����)���<[o��;���;}���S�:��h�����'��~�V}��������X��<����pU7��P�;w��� �qԂ�u⺭X<
�����/7�
��������ۻkX0��N5�yzHwȅ�K68�q�����?]��,O=�iD�:��:7s@8�2;�U���	�v� ���}����s���[�3�o�M�5�����{)�~���{Wnn��>�3���m���Rh\}���������������{�Zy;o��8�����|�gOT�<y22��;��R��^Ns��x�"�"M�?';v����K�-�P��1��^1q�~����qFr���{8��Cq�?}���E�;{�	Fp}lP�=( !�aK��P�$���7�� �@x�>��,f��q��ǋ�	aa߶ȅ�)��O��o
O$��8
��tUߒ�x���Tݸ���X��O���M���o ��#�4�WR�t5l�ۅ��u�e�k�y����z���8���)$q�Oq�#1I26A\�,"����6EEq�6�棩q�G��1��������ӧY�K��l��!��E�qp�T[0XERBUm�1�j�(�������m�z{{q�Ӭ��ܹ��(���Z*�⪪�	
�#,��MaU��\W
�Uvb�O���������:t��z	uZ���1E�feqUH�\(��jE  �@\\UQ�Z�m1_f]��Ŋ���l��v��,H�r8��&�6`E��+*�#��jK+D�U5\s"bG+1���"��IDqyAH�Q98�͋2�m�qE�D+Q���8�o&�u��fL5�)�q����$�LUlp�h�#�XL��X�r	$���U	&�.گ�����(�9jrm�����$�a�C\Ɉ�k���eB�����T�"�c$1WFH�⬓Eu�$J�bAl���X�*#��.b�&E[��H��ӒhcGc���FYMid�>�vE3���R��)%&��6��G2#��]���Q] �z��#�o8/7	����u�0�d3�Xw%л����d�pǷk�.+��}��D���Y�R�R��\���b	n�ݨ�"&g�����ZG]֡�Y�\�8���������ݢ-a�4��_<<q��v�(f�<�}N�޺x�f`��`�h�� ��"��Y�$�s�vq�,�ֶ�O^.��ä{�����3ݸ���7R�N���=�I�ⱗ-㮣nEϛq�S�8D9�ö���P�&�t�-KtNc/]�#�öl�e(*�]v�4k���m��&4[����l�[x�m)�6��c�6(]s������e�x��a�=�C�닱6��@Fmq逖�S@"D�T��@�m�\vng��5�k',�,�tpqڛ�.܊�H�v��A,V�۳ �v�Bh�Ѓ�43��C��,��ɧ
��p����{�s��)y.������	]yf���m3�Hq��n5�C�����V6Q�cMc��%���G<���܉ �=n.���%rs��/̘ �Y��˝A�n'/V\W�iN��<s�8&l��5�q��(�wh��ֶ��ZLa�5&�GF\��b B]�1�M�6�����H�l�;\i��K��`�xq�7Y�ڲY�q�cX�����*���j�=� 2�܁�H
��Iu�2nфe6�-^ ��c���LP��׮ۓ�Lj���h;��K�֛��>=A��n`3�K]Md�7�5�l��c�u���q���3������\���.�8Un�%[<-�e��q[c��p\08mt<�7k�J�u���eGk��-�\h�Mi��Kl ��11��.���<�'ť�b����Y<��݉�1s�;�R���������\�]T�-z����͊7f��X���b��]�ٺ�Ñ�'A��Z��j͕$��XS�X�;�8�8&��	a���X;1ԛA���!�C4BA�o˱�C-�#Q-\b'q������f|���pk�7f�</�,���݇V����`�,�sc�l�Q��ab��X�»Gs]�N�7�i?�_�m_?�x�gc�f�ܼ�t��c�v_>��9���p7��9�oY�׉��<=ݿʉ��o7�G��:#���g!@�;!��/�@��Oe�\��ft]��d�Dx����m� ���Y��v>gy
:���%lt@�����K���T�7,Ӆ�����?m8�?��%�[f��ۡ��ѵ2=��BB���IЉml$�э��	Sv,�$v�DI����7�:8Ɍ{�Z�=I1V��gs��:�]�;���M�/IXm�86ɺ��=]r�B�L��kӸ�'.����:+i�׊ ?�!�$��kq���O+K�����[r 4,����U��b���3@��*3c7u>��"rhu����p^�_Kѵݹ�]f@��<�Z^x+6����LňyF�Ζ�2��s<�D���6�Z�xDc�9}1|W�[�@$��
�a���@��^� ]�uHC� i���$�wG����G�Kԍ{�9��v�\@>o��������;;��賴�a��.2�۸͎'I�|�5�$��ת<I#�2/� \��]�<w�.�Ȃ��X��K�vi�fVl1On8WFt#�g��-��	$d5b�A�� �U�!G�������1fA�9wr����w8ݕ�<ڬn��LR]F�b�h��"RZ���V�Sf):]p�@$����|�>�|�:����j^�]�H�j�$,<rL��,޷fr�ظ-�[}2��ʎ��Z��	=z��~K{� ���Rr���h�>�$���Avb��j���z�	"a쭜�����.37Qm��r$m��[;�F��v�����_� �f�j���߽�~͐8w~�_�qW<1]���d�7���	�����-�$�wv��yZ���%�v�y��cl1�	�U��Gn�@7䆳�YQ��#�d����m�\��L仴�7�t�O����4�lk�Ϻ	�k����Z �7����7[��.���d� Ks���/K�Kw룋ۮ���^���!pZ0��%�҈MD�������Ap����ee�A������O��,Q��A[E(��/"#�ݳ$�wEg���I�L���=�Ej�[u�۴��� �ǂ���%�	׌�f�i*��L�������;��EtA ���/�"y���~���v�$o���@;��P+YL��1k�P<�j������Wӱ�|f���D�l��O����T�f�e�l��w�-��=P�6!6��v������C�j���L���>�ۼd��FF���$]�B�b䝲�Ή��G��{�}Q �C�w�<�����jޠ>䁦[���ΕԳ�#컘�O��݈;w!�5��}}|��j�A�b�1RK�A�ؖ��&q����5�M
��.v�b]2���6�;����gn��L@$�e��	$�r�*�'�=I{`O�6^d9�ǘq �BS�m�-��]˺�3+��c�b��u��Suc��|���"	�%P��%�l)9�B��n{��^�"��f8Ίv(.���B��0��s4
��;[yg�����(���n���4��;�N��g�Ϧ{b��w����$r� o�L{J�P_��{�G;_lr��/�W9>���nw�ƐI��)����'���g��S(��$�H�rD�TA ���PȠ��� ����,�9��H�f��9rkI6�*+<�j�*��=ވ��E醛�v���>�
�n�l>���0g�?r��Q��q�;��Y[�a.E�a�A����hn4ױ6Fl�"������O\n���Y�LT��uG@!�f��������)I���]r]��[KC�r�v�$�NB�4a���Y�����-��6ݫͳ��PK*B��1&틨3jQ���fW��w�[�w�V���l�|V5V�z�7ZAN\cgbS��[���<h;7���'jm�^3'���ssh�Sn*�Ӷ����]	��~�w1�����ƺ��P�T�FolA68U��͙N�lΈm���b�n�����w��k��R$�s29�L�M���A�YhA#;�#�U�ϐ���+h�VLz�Ga���Iw.��]|g�]�����:�y��dH*Z�Ao;�b<H��E[����*�V�7v���n�����mVSo��'�/� ��J��$s�Q��%��C��.� G��Ĵ���N��j���<`����r7�c.�!c^o�I]���O��C��_	�z���P����6�2�c����5y�4y[&��̛C:\���g�ϓ�ԙj�;�mUCz���D�=5�m�+�A �}�/+��`]�\I�c��,��;˓A)�q��4�-N��,�E�!��"�D�閙��L�j7a��+`�-8!���r�s!�[e�&Ue���3;��ެk�U��}���bm�1�$���>D�����Ͷ�`�	�]r���2�;����wU������Fy"e���iɖ�w�a�?�5^k��yy^�>�q`_� ��ѺS�Z�d.�Bz׏I��@�zyV�-Vgn�5DǴG���	�l�+X��س0� ���A�,�Av�[�����cw<@� �_L�RR/�d"�����龶��-qs]P�������c�� �Mq�:�vı�����e�������˲Nwz�)�<��k�	��y[�m!��x �ODxג'of"�"��9f)�Ӱi�z�U�C���G�p���� ��A'x���,��Ǖ%܄;M�#)���o��W^[�����!��Q��A�O��	$۴����9j�!����wc����w\ ���=O.`꺹��=�ol�u?\�cJ��O���v*n�ެ`�0ܓ�����[�$�l@�A=-ܠ�	7TuZwg);�Nn�GLOd�u���w��	�� ��9Oc�����z�$�������{{(��]����y�������v<�yD��F<�^�ƂA"=?���=���DbD���(�L��X1�a N�8h`�<C�Ի������jKM�~z�S�c.;��ø�w���� �{�"<]�t�e��a��`F;	�$��x���xt�� nu�C���9Ż�	�#x�D�v���}{�����5���ܧg����uP�W�{������Z���R����#��l�����N������0�>0�u��������6q�<�ג#��x���ȓ�����FRa��3��y,�&2dy��/�Ú�燱q��;W���'г��z��Ju�=�Vi��#�}<�)x��>o��fkA7�:�:w	;�Loױ��H$2��{���������M �=���D���}x��\�;Q,
U��v��Bb�iy�����n�yp��d���҈9�H�!�U��o�=��nώ<���p�Mk�ǉ��zb��
�?t�J��!M[A�s/^I�tU�N�p��d�=Ǡ��_^^��7ŷ�d���tE�ɿ$��	��lp�(�\�v�K��#ݜ�b੟w���x�EWD>$˖���kަ�I�΀79��^5�:w)�ði�x�S�71����n�x�OnCǈ����y�<*����x��ܫ�!�w�٤l��އ��Q���f�C�t	�����1��l:�JsHq�29�s�16Y��BjC��1��B�uMi����ܿ<�S�w��Q_���X׆女u�C�*;)�b�$��y/���	gTzË,���m�V�+��ޝ|�<|6*�ڗh���MŹ����[s��v�{s���:.�8"��1,�z�,a ����4)�Nsd�	h[*��uv
��Vn.��E��&��#fF��Scv\��`�i�88�������6����n.���^%�k.��h�^����v�8K�ǝ�.t��+�Fѫ�0qgx��םqM�87Vs<�Hk�H�r�Y����6΄"�8��%��g�$��~��~�Lm���"�	��;[1�'�8}z�܂]ȹ빀}�툃��I�ӌ�pή�`�\ �VT�T��=i�m���~A�ٛS'��{�H3�Q�a��<U�H5��>a�\;0�V�ݓg��lGz^H�/
�N�n�D���'S�4|�����&.
�������[70�c�Ǟ����z+�$��^�舋���w���x��D��^:gN�'p\�P:r��^��g�7(�׉ǰ�C�S�����$G���A�q�[�<�Z̟�7�۰��H���V���\/q&h�0�Zn�T�2�+Hl���F#j�,͠lp����� �؀]�3���v�����؀O�hu��N��Y	�k��
����>Ƥ��8�r/��-��4=�c5��қΰ��[2�{�ȝLM��ʍ5�S������{9/QY&.j��
� b<�xxKC��KyS6�A���DH+��ބYT-��8�e�y�L�%�QpΪ�`�kG���v�)'�7��P���%s�� ���h'����)LMM$�1��feg\v�ޙ�u�-�x#�� ��	=��$�w:*oF^3�mlx��%��V�vbD�~���7�숏_��y���8�X�3��I��}��Fs�ɧ*{���3�	ښ ���� C ��H<n��5X����is�.���t)�ﯾ�K��z�&V� ��&ȇ�I^�@��	f�]i�a';������D8R��J��<����L �|NwlA �M�DDx�X�F�K����fZ�MtR�;��:e�3ѳH$���hB�L����:��~佈�w�=^�8�x��uNI|��GR̗ۤc{��oi��o��.�H�y�$�{���n��������V�<y'��]��y���U�c�P�g1l2}����t>"_Y�{����g<���:G�P�S�����D_5��}+1��w8�6��v�v�xu�Xw�d�Nm?9�)�9�-b�?0�|=/�O�{7w/v!�b�����g���%�w� ֬���q2���E����v��{r�.�������#��w���6��7v�n,�n��Y��3����/[��Η���]�K�ޢ�zxd�	�G�)S�X����J��(�f	�|�C�\:r���6����xu�۽�;#�X�*y�'<���i�y���c�7�ż���D�E�#'�dG�x�~���-��Һa�ݗ6��=vEC��8��g��7;��˂�Ċ]�Fx�e���
���0�!��ty��ҍs}yN�^�_�@Ȗ����)��,�Kً��$�$��ۉ���:8��`>{��'�e�ؖ��������\�Z{�06e�G��W��&�ú���ˆн��[�6;�#sP���qM�����b �*��3:���u�3b�]����1S��;�{������\/�����x`�｝��̼��3۹��۸��^xGe$�a��K�!�ɀ���
�Ԍ�]V��8�T�/n�:9�ZuF���ٝ��˗����8���� �x����Z��Pˤ�3{&u+49��Q�������<<�����&I�X�D���K�BH�*EVH�"��#���8�'Y�;i�c��ǏOo���:t�0�Tǔ��3�ER�D�AB��Ԁ����A�#�vx�����Ƿ��:t�ӫ��.�36ER$�b���9`��UU�ɉ���
2�K	!22W��m4�>:|zc�ۏ��:t�Ө�"���$a��1Y�
��X)�rHkpU�^�����"��8$��\�19�1qG�kU�b����b��;��a
"����z������DTMu��*�ڸ�6LlU�(��i0�����nb�I �$�U����rLR$���R��^��zӛZȤAs�aȫ�(� ԈBE�󚂜帠��1*�
��QK&[0l�"�t�U��8�""�ʢD��ޓd�&.%f]�j3"�b�"�	&b��8���u����6E2l����� ,�R(�r��.��l&XAW�Œ�+%��Qd��$��>��i6�|xofD�H�ޘ�f|�M���Τ<.���S���S�>$���I)��O;4K)�V\DF4$�1	��&@8�q ���%y 3�cWC8����k��h�6y���܈oOKU�O���d���0�'p��"z[���86�MIqa�B�h6j�S-��k����O�;1	����WT��S��}T��w:�v#�����y"�DEcκvN�ɜ�M{T&��������j����x�ws	K=���A��D�u�����w�={(��*N�K����+��=M-0�ԥ����%6P��]��2[�@$g���$��vt�G���꩗�V����м�55-أ��o��g�@a�4�D�ɸ?r��.�V4�1l�[��q>�/{��p��8'߶�jyxKS�ݝ�.��6Ecm����Á5Q6.�Ȟ	';@�(�[t�`Mws�ٹNd;Qפ�5�[� �e��Iݾ�,��D�� q��I�.�Ƣ�2W]ɜ-<�h�����p�J���n����%<[aBK��:��C�v��.~�>�� j��$��v<xϳM���yC�iv�s��S�� ��q��rgf!p�P���wNb��[���I�Kf(H��"��Gz�1���Ν��b�æ�ڦ[��$ev<'�S
�>�s2�� /$zVڀA��}x:���rT�f��r�����ޗ�:	��_7L��$���@[ �� �E��&�NG��=��u���ץ��%&Qə����@ ��M��Z�3�w�W����v�&���vD�W���U�ۜ��vol��b���_y�Zu"rs)�D��g^�p�������jz�\� �����1�X����1�Y�g����V�M��L��N���59u�f$�4n!+ְ����wK<�G˲����Ɩ�靺p�F�[�BK�0�����*�n��7P���=7���˭���0,�6�!Gq�)@��v뇲Lm��f��].��%�٨b5�$���[�\褣��6$HCnڣi��JD��4�ݘH�6�3ckH�1)l�b��Z7G]�y�[�c�:Osז�M�wm�:��E������g^�>�M4qZɸ�p��0\�D�5�j��=�e��1ћy����+��5�����<@��Å��c��\w�v�P	���,aBa�û	�� ��Ü	�;-HʜL�(1�'s��$M�K�<A���Ъ�P7����e���B�#�~�|�y 	�x�
ӳ�x�nF- ��ȂI7�1O�"��t��8t�G�Mn]5%>���}���}���A�m�UOb�w=kۤ�zj �mJr�gf��o>"�wg��C�6K�:9����*�ȏ|D�������Ә�zl�|,��D��6ͦ5v�#��PF�d#�wDm���6I��[M�='߫��;3E��0���['o�{%o#�<���hY�~� �r�;�Fl���.��A�[�������<�vxO�=�ך?-_�\S%����wX�na��1RC���4�q=o#7%�(���r���[�6%[�z�f$���/���k&��5�y:��&cʹ�4R�K4�Ss�3�&Q��&;���k�ϯҫ�x��d ��y�h{F��.��$�_@�I��*��,�N�B�*ؾ��-؞��X$1�+Ă{m��$��;Cɏ]��,g;���t��8v�
���p���x�w��$��M0�`�����ȂI������`����߄�������6k�,�5[�{veչ�x�u7�oU�[��sJ�u$I߇ߟ�f�~�������n�㙽@}K�W7d��@�A"������1ԝ3"���0�m���R���#9뭞s��_�I�Z�o�Ȏ�>�b�F����	�`� Jv��4�U�� �|a������v���C���ٶ�0�o�f��t�G�w)���$�5�6�hi��b�ޖ���W��69��$��kM!ds�@�-�~���	�-�n��;��br��P���;&�j.�DC����jk�s/"}"�Lk�W���i��R�P	o\`��S�!p�z��8�g��q�]Y*�/�`���Q�I��x ��k�'�o��卒%YZ�8u��e���Q�qx���"�H-����эu�֡=����-��]��O�� _*�b��x���׏h�x��x�{��p2�t� ���x'M�B`�Rgg��u�NU2� ��[Y��~f� �#�*�e�v��c_%fgN��a3�3�>$�>��	��'F�ƍV��{�9�X$�^8�x��A[�Kx�RN�E�wN��[�Ϩ�[5�|W���"|��:�#��0�1+'���N�(��2WZ騡w$�Ԥ9�ׇu곰��ӷg��p��N��ʉ��o����~nc~��z���Xw���=\�O�����L1˻0��&�x�I���<\��ܜ��h$�g���I �v8��X��BN�<&���6���Ã�ˌ)o�:�]�n<u��[�z3f���9��e�ߟ'����j~��~Aǚ�=�I�7?1���a$)����W@�;4܁wp���'��떘�nV� IE����"y~�1�]�
���'�v���(q�X���fvz�� ג)�����T$�U���O���G�@����ޱsZ�33�N�0������n��H$���A>֧� �{{c����U���� ������rJڣԡ���@D�׃}[��ٓ�w�H��Bx�y��+��+�-�Wf��%�Tg,���-�2�C+<O�Ç�8������-͘����c����4�}���ga�]��b�	X��]�C���z.y�[��l��V:g�N���R��M0+,���!�!�u�yѫp��u5 �N!�\�c#�/ul��<Te�1qCL�E$t֨��.=�q��9�:�ѩ9�mu��� 7Vz�����H��2��ۃ`;.��n�� �3�]�-�`j7^�'B�Dy��c��뱂��� �k[ �mm��:�%i��n-ǎ�q'={W6�`68�Q������m��ǈ���f��Gp\��v��l[uʜï��RS�wm9����7�Ƕ��>$�׃8�#Lr�3s���qos�%��у�$���V�8�k�n$�.{���2���!��>����R<�Dwv�ܖ;������7f��.�Y����Od�� �{�	$�Un�M2n���kx1�N�k�>�^
p�-F���c�n7T1�%ۚ� Fy��^�"	���>B�n��U���x1~S�a�G�&wN��0�Z��e��'Vf&���7�{n"��ߌ�:��}�'XK��f`P]n�?�10�q�����<����d���ɵ�X�F�-a3�>����Q@�w󭰉�$�=�	�9�����Nb�h�cf�)��s1�S
��k�va1�	��6T� �uհ��v�p�LWMFFs`3!�7Q�4�=!����jR1���C޼<�>
mA���|G�+\x=�v��8�o�Q3{�İ��l��dH������� �-s� r�77��уIoth�ΊvA9t�>�>KyWEȂI�y�Y��	�ɒAk~�O������/c�;6i���;yؼ	��e�ސ���ǐ�Ky��A�>Lω3��[�7Z`3�U��٘�������b�a�N�@��x�T�<�#d��y	pH���$����K���%)������2�?h�bFh��^�.�7XÌt��#.Z��a*b8��H�{�����`guz��@$7�����z7�@7̲q��4[�]q��A�|^vù��$Iv� X1Z��lĽ�T�FZ�F��y0%�:=�_� Ba�ƽl[�S��������L��'d U�] A ���$ff�5�jQ1i9S�[)�.�F3��zF79Y=L��8�{{�y�U��Vnk/ȡ�9����eǚ�l�Ŀ��zi���I�~����w(&�S��9)�"��UPwC\���a��7�������	�7j���ok���m&A�"��=S\�$��΋ă��a�ǘ.l��L�/W�Q�[��"�ʉ-��ĂF�l@5��^;C��b��A%�D<c)3�&��б�+1F�1�U�W1�G7=�/�q�+�XÄ�ׂ]g�s^������y,�ǃ�i��푮�u�D���@$�7b�#�&�e.E�˳�$������M8f���������A�Yj=ݱ���f�K�VWaǊD�r4/6�H�3��f�^ ��634����U�>o$O������Ey!��	�.,3&dy�9c3�5�Y�D
��B�;b	'���2	'ǚ��Fh�Ep���HM]m2�W�]\A�\}���#w����֝i�:� �i�ѝ�N��o�mSiH�����o�A���?�xK_�vH��*��_$��W[��E�FN��i?)��pK��)� Y�]�̉}�@� �z��,v��Քjֲ�\]Ɣ�����}S<ꃩ�`|\�ٻ��'vgo:-�b�PIμx �O�˝���y��._�m��h�$��� ޜ4�!��E��d��ݑ���m��||��Ȏ���/ �)7n4	/1�ߦ��Dz�F�fL�ْaY�+�Kwtx	��r�����W(��: Ǌ:��"C�6��$v�л�ڛ���'�v[�$u��$ s��Qg��� ��<�b�2fG��� �u�ex�ܬܡ���|W�U��L��jl����?��/�G�
���( (������뀠��~vY��Ñ᪀���AX! �`�X2V��U��0@1 0`�! �1#V1�  �# �EU�D  �@A�EP�@���B��@5�Z"�J �݈Z"����-H! �@!T�!�UH!�P!��DA
b "P�EX!VA�`�X!VD�E`!VD�E`�EX!V@  �X!Vn�V� ��B ��� ��
�B"��+ �� �+ *��!b+  B(��+@`*���B"�A�+"*�l[�B�VD�U`�X!V@ "�Ebc �U�E`!VEU�U`�EX!V �  2QX �U�U`�XDU�U`�EX1��U�U`�X2  �U`�TX0��U�\�􁾠Q�>��ED�@H�Qc��+����_����J������j���?��_�,=����0��U�J���_�����=��(*+�������_�v�PTV����a�3�@�:?4���?��?��
���C>�����B���S�����	ހ����l�J�M ��Qb@U�TX�E�TXDU�V$EXEX�Q`E``��VUX�E``EE�D�Q`X$AX�QYV#VX�X�Q`�E`�E`1b�#"���"A`! �`$�A�+"$�@��B#"0B)$D�"�a �D��XAB�EAET$DdV@U�Y�T�EY�Y�a�UdEX@U�E`@ #V$QX�U�X��bA�VaV?�R
�EE�EZ/�����?m�r�( � *$��� "*�'�}�������߰$/�4G�~'�_O쀠������ѯ��gò�v'��?������������>�PTV��C�O�����@EE~�PTW�����8x}����j�
.���c~@EEp'��%�iv6�]�((?�+�����&���E�,��y�?�O�����AQ_�<O�T]�#�>����k��?�'�hXt4�
����H:?�

���o�������.�����?��}��`x��:�v

��9#���)���z�a��v�����ϋ��((�	��E������O���O�����)�Ң%r Ł��0(���1�� �@QCZH�V� &�P �
*@ ���P�� ��(@�5T((E ���$Hn� �J*����D�A@DIB��( �"�J��D�QQPBT�J%H�����)H�TH�H	�T�w�   � 
 �                    P
   @�  h   
  �V�����{y��
j�
uZ��um���+E���й�t.wuc�q���w�u-���TJ"*H�N�  q��O��ks������[Y��8��0�`=��k�4 P�< x����� {� o=�y��ע��R�BU�  |    �   �
��`�� �`z�  ;�9� {� � n��X�= ���[�̀ �� �甽�P�k7]�

�RJ���  [��ڠ޷��ʥ7 ܶ�[�ݳ�ԫ�R�{�K��ڳ=۷�]���p 8�ե9ju�Zsnͣs��V�nq�j��$$UD�|  �  � 
 @ 7�Iͻ�ӛ�.5�;W-j6��mM�@�-T�������Թ�[oy�H�6˖�k����r��4�n�ʁD�JB��  ��}]���a�����m�t�g��y���j˖鵵^۽n�+c. u)֜ۦ�MKu�j鼘���;�W�3(�
��_   �  z @   >�|�ս;�S�55����)�7J�ԫ���6ٱ-��Nl.��s������Y� ��+S��6`�;)sUE�*�+|   ����:*mm�u�j�� ���nv�m��Z�4�ӫ��Z�u��l� :�v�s��M�[����l%�9���V	$���W� �   P     .�m���;i�������B�w6�%à������V��H��v�7��Z$���[8�]�v�J��J�J��  M���
��E�n ��Pם�9St����{o[�^v(W �����v���Z�ckk�ukQ��n�c���)J� 4hb)��JTh  ��UJ�
J� ��=)P  ��IP�4 bd HQ�b�Q��2O�������?�kQ���h�续_�>h����S?��� �$��k?�	!K`! ���$ I B��I	LH		���'�����ޞ~��l�۷�[v�bg(j�e@�Sj�i��͗����e���?� Z�n�Ů��<b�jܫ)^"�iv�=����2�G���pǢ���vu���}�,�����u�+��i��-P
�w[XvDH
�@��^�Qc\�*�ح�3-54-i"���qV�432����i*y.=�M֯�����V3[�h�V���M�JG0k��ڍ	��*���ّ6UfB�[7&���95���6A��S�˜k�7-�J'7��-�-�P�1��o0�7L��ի���U����E�wM:���8�ӹos0�S=����C%m,�ɅU�.���`�ɰn45�ǒ�aB�&����2�'{���f��V�n���C.`��ں��ܰ�
{�j����e-y6�"���6�F�S���.�P�ti��w*TOeE�M��fbK^�Vk��n�F�dbg5�V*�!h�S&kFh9zr���+k[V+jn�ܑf�+��諸�Ck.cN�����g�4]e�X���%����;j��I���P]k.�ԫ�������5xM�Eb�mF�Z6���^�bjy��@Q���G^\�{�qe[���VE&�����
�M�O6��R�ք̼����Wt�^�r�"�e��a�0��7$�3,\���o[7N�eeV.;�2ŭ��+A�ԑ�ɺ�����G����{���M�-�(�K0T
��я6��ͽ�QQ�T�Df,��a��)0��ӳa�o�in+2�8�9�"����u���G��ɊXNs����򖖺]�?j'�K/7�:p�:��U��j�����K��;,c.'y������k���G6��e��L�Hk�l��z��];M���K�n��r\֍`��r=+�����U3��b�ZC��Xg�t♢�Uhe�'���ua���ռ���G󧜞�%Ѻ�p�a@���%>�c@p�I�;y3�.�7��%�ͱR��2�:��a�EF��UJJ�QkZ��7�L�Zv:Ú`�j�ʁ�湲�V�Շk
�v��7���0��IDazi�����q�hM�0G�EmK݁<*�/5j��b��I� �Kf8y���9�o�3S�
 �j��m,�jwz�t-Ǵ=�_r����$)%կKR�M���M��:{1^�W�۹`�c*m[�(���lI�xSRμE[��V�嗊�nJw�z�ӂ���С��	�nD켰4V�y�; v�q�V�U�͗v�c[���(�Vk��o
UҢ	 �f�fKR+��P]��5l�,�T��w��mq�U�n�uH�5t��Pb������Ղ�e�PN���v�Ė�d�i�B�:Rf�[kv �$�\�U�ڬB���6bⵐ�$FB>a�WV���^�775G�8����]�y�u͌���R�ZL��V�3+�ڕ
Ϭm�^t��)�:�ju����V]Gxp]�re�T\�YxK��A��<�*�Z�F��Z��p���z��\���B��-ּ�.��]\��f%��aa�M�O�X[/�=�/us���|��ȴ��.j�|�V�s��ڻ���[����N��V��ML�N�T�͗BD�sc�D�AVՖ"�+7r]��1��j����
��p1���V�2��dT��^D�:�8U�S �t�fcsifU��X?]:����/aǖ�h��Xa9���NR�n�,7vN�u�!��~X��B�U��g���@�m�Gq�R�edR�q^:�շw6�%�*�*{ZQ�02\�aǃ3M�`��ۓaR��ݿ�D���5��\�-o�=����ʝU/�άc�3ѹn�V�ͭjf
vZ��jӁ��R,�,��r[��f��`����~W`ڂ�ʱz^	6mklw���w*1`� ��HG��0�uq0Y�.�ν�n��gfn����'�[`�)�@��]�BT��ײ �A�l9��3QúH ���[x�X�Z�O-�a�ɏJʴ��sN$h�6�d��
w�l�\i؛�"&��uՍ���ۼJ�Ƃ�Y�z�5�ɉв�n����PЫN9Hn^Up��}���{��]�H��\�cm���O�p]ujLP�,.vœt{�Ȋ�6V��8���ۻ{��n�L��R�ދ�ӵ��j��eָ�h+���.K7y�T��|�,�Pۏ1�de����Xn^�-��9%����~�CcH�[�-mcH��|t�Y]��/R��ى��T��x�N��18�$�"��J͈�e����Zv��V,	�:Ag+b-L�L��c<�d<A�t��s0�۷V��vb%�Ee��Gt3n�D'��t(Pv3*!1��UƯY!o1�� �+u�'p�F�Yt�2a��Qta܊���'l�IW��Xtu.m�!X)Xe̴#�����T�&%Yͫ�F�Ù�+m��^�aXC�(�ؘoiV={��2sl���(*���˨�;ܴ�mO���'�2�J�t���)^,D^���k\5eGM
f$-�F��`[[O :��ZP��Y�੗��Iś���kr�Z�����<��GV��	hՄ�*�bAv�NJ�=7b�vw,;κ�YF��UuM�{�P�T�����gr�Ch���V�eeR�����u]u�i��)iN�����1+�39B�6�-�t�;in���Em���]#@M3ZfR[�����[�oH �,1Y��5����"l%�1�M6h�A�3B��.�v�i�=���7�r��CKlvUt��tz�^��}c��+�����5ws�\ѥ��������eCFf��$��cHbs/f�Iv�慙��ڶ���C2eB<Ò
'S�L4�[�@�5w�c���;��H�v�%w�������n*I1��tnU�8�V�w®s�u:�����j��X�&]��ɭYNݚ��d�Q�{I�re^:֣Vdmd�M贴n���y�,��u��k�Y��kvj��f�C 5��X���!c\�wd�r�<�xv�ۙP��yr����kkV]'�e\W�[6[u���Y�&�Uz%���"����`W�	#[��w��^���:�j���{b����ot�v؛�b�ĸUec�	�(�ɘ�l��k��&�N}i�I�wX�ޅ#�*+"�õ�N��:-�V��,`��њ	;�H�/�(�P^;����n�G����6͇EnG[�}n�����c̥v��P����T���%�-����51�
�>Gj�pvB
�;z�h���6��[����-�!rK	-$��j��D�r�M<���6�QJ7�u�M+ս���͘�v�v��c�+]�Usy@r���t��Ajr�e��0���a�w/{��M�sv	4V.2�.��`ekPVZ��u��N�hA/C"ud�i������9�G��N�x�����]|+���1*��-���1��Yn�����!�:�j���Ue���Q)��>�ؘorM%i�@�V(�S�^��:p�؛�i�.� j��f,VL��IlÚp�F$m\�OݩI�`��#H�����;/l��SCۥ���ؖ1�=%ݪY�t��e���i�n��v��z9�����Y�PIdM�Q��:N�ןR�in�tb��cY�Gj�1���M����5b�Q���;M��HF�2�Ve�kE֜��;z����l�ؖh��e�P*�� �9�yx/5��j	6Q�G��dB�#S�Q�.��O<^1��`XZ�R����؂`����q�wY[����헹�%m���Wr^�̧������W8nnL���)ճ�v�;���b���Bý�Z�V�"ֆ[���-��>�ne�"���c�uk	�(�%�Y�ÕfݣN	EYݶM�
��t��Z%e��ۼPi�K����o1��J�*S�k-Z�.�!Vj��r���ha�-x���t9t�p��r�^S��em����!a�R%b�6�����gEԓ),�L�n�����B���bЮd,u�ֵk	���P]�uw�q1bf*���j���P�����%�kh����;����#z��ٱ���;^����Dn'o`�M4�N��i�f����s^���&�7�n�e�ᨯn�+��^[I�lS��mIk3#,ᗷt6V�Ĭf��#��O5�gP�I���5�lx��$�;#RɈM^�äهE�p,��ލ9t��� [[Oq�Gt	t�I�Ԫi�J��=� ���#\M�)v��ͪ�bxNBY�"�_��,\���6�g�;{w2�K�p��a�-\wl.�*s^j�2�uv�J�U�w-k�+
��Th8�S�dC��ZH7��f�y���j@�K�����#J���2l�U�j/�H�ӌ��j[tN���0�sQV���������q��
;I�.�ϥ 6] �ZĐ՗gV��A�p��Ƀ^80cKh�K�ۅj��:�tP(�[mV��K�m�9HV<����� *�L����Y��)C[1n�z��=�QB�w@�������5&�̷�ζ��쵭�v`�	w�TNݝ�/,��mⳒ҇�.5�Y.�>9�3,�F$";���6^��� ��Ɩ	X�w�g�0�+��.���W�YE�.�&���Qz\:�1���D�Q�����U�{W���jQ�!��t(큙�:��ʴ5&S�4��Z�c9[�/	��b�n7�5�:!v��d1n�n0/.��^fM�B��RF��
;,5��2M�Ķ����0%yz�.�n�������Б���n�[��h��F�9����[�1�-�;$iZ7`l%B����WPm"�Y43(����Gr�:U�VE�m������N�L)�V������n�paޣ�X-�'A�h,���)!k�tj�S7R������ו6d��p���Fu+���$=� �GQvܕ*<	T�n�wNا�Y�P��Q�yNMv��Ȁ˗yr�D��nֆ��--z!%^n�K��}`(��/\[�Eѽ������f<��xFiV.��ax���(�l����ۊ���V+�� -9R���إ{Q0�RP"]fC���1؊�蚯p�n/qX)�|ۮ�o�i��Zu��M1l7ݴ����2��0���\�@%��C[�������؄8^���a8�դ\����;�,�n��֝�?��wKY6�5R��J9s+kP���-�f��g� ���Lf^�Y��2�j�	�H�{S���۹T��A���s00Jqg�.4᧴2�˖u@��7z!%F;������7k2�!T����P@��y�,9��v�x�h����o���n��D@�����T1k:� �pf�0�ɬ�IP�Q�y�̤i��� ��ᗳb�[�R��j�����
�V���M�l�M�����~�7^�e
�/ ̖�e�!�nn������F�Z�mh�����6�qc�ed�r����w9�����|T�8����[Z�C����:RهX�2�;(<���o,g�c�l7{�^:P�$�,��`�*�Fpb��1ű��l�F��+(��(jQ��j�4�R�n`�Y�o)+�-֏ r�]wU�F�u=��ax�z���ãbV�E�0:�����*�U�hৣ�kv������q��.N��oɪJf��3muw�P[rҔ�-"P9"�iV��4�	��$�^a�1����5�걣~"�� 37��]�b��]��-�&ڡ�Qe�����8��F0֒�kb�w��fN��f`��Omk �\%]�f]fh�TW��Xu:Cy	��p�Y�
ek�[�v�3w��RW�����n%��CoC�K�Ǚ��j-�cVTdǀu��pn������}w�h�և�%tԪ������B���YtwM+
�%��x�S��I�8/]I36�{u���U�J�i��mސ�u�,�ec�^#���4�M�Y�Wu�n*''��x�j��M��i��kJ�dE'� �F�N�"��n�K�*���%�f�� ,�>�[�wt��.��oR"�^H�R��n'd٬�o�@�@�5
Ƭ֦�͂���3�W���� [�uXo&M��7�-A,�Xw�P�f�Ov�gam��	Rf��1��,4��p�NfI�I�h�V��uv^{����5���]8B��/5Q�O�x��{e�8�Z̼X��:��2�4��أ�ՙ�n��2�n�&赔����ϠR�ѐ7.��T����^M!�F�d��q�@w���ܪ{|Ylv��we��yL���.^��т�l��Ujj˛%:x�CXc�-|c��u�SU���bffmI�bA��ʛt��	��*����'�%�jRR\�M�u�v�<���u˙6�$n��
�v��l�jL��0"&��E�r��A�iaGu[��# ���o	���t�n8�R�.=�oC�X�],&m_W��b�*$v�����4�.V�[�ZAs>�f�
E�xfon�V�un�K6�z+U�B�l��\߇؉����i�^:�yED�^B�σ4��Beٸ��Y�Cp)w �N��!�E�ъ��i���N�V�c5EOia�.RYz1�o%+כ�m-��E<�r�䀠�9m*�Ê$6�r���u�^YY0ʲ�S^ُ-!H��WUla�i��Xe!ku�2���KL�j��V�#��:��N���{7�Cw�be��/B�n�-�"�F���V@^`;.9L+�}W�t��_gfbE6j��;��ͬ���a�n���7u���Uk�j\j�p<��f}�f:�̎;��)7�ԲHE+��.�rf*5�f���b�Z�	0ъK�ܵ0��) b6	6$�6$��	����:�.����:����븺��뺣��.���m$�6	&�B_ͤ��4�� ��BDbDimww�uwY��wq]�]�q]�Y��E���ԝuQ�]�Yu�Q]wq�U�d��BI 6$�4$�H�4�"0J4 �$��.�+��뺳������.:���㻮;������˪�Ϋ�:����.�ꋺ��;�����.λ���*�;������ꋮ���볫:�쫎뻎�:�컺����븪�뺬�����.���겺�뮎뫎�:������IF�B?���@�HH����	.o��u~���ܭ^~��5��f��_��h�#��X�����t��ܜ�.�vyʯ�T����D�\���J:���kt+&
�}W�HsU=ߧ>Ra�\���^�K���G%��W
�ٶ���(+��F�Q�چ���/��㠻��yl%Y��is���U���\1I4K��O��W_"�s��־�pJl���m�o��e����=A�ȇӶ�+9���m�����*�LYi����<�:%j��"����o�[p�]S���7f�ώ����GSRV\2��X�R��2�H��U���r.�m؋n7�j[���T�6[6�!
���Ӯ�c+xt���;s�S������l����;�ٸ;9�� W@��eɈ�/�Z�սŦ^�r�ʷ3F]�rҙvv��\�b-��e�����$�L�ql#��S����F�S�]����k)��@dN�
��ئc���9rpۭ�����
7K�eo*�g{���ړ�s�i�����.�L�3f���Yu�r�m�LW2�X�({�Z��y厤�z��jU�T�SҶ�W+��.�YB�D5�tx�&�˯x�E�+]���wp,�eSN��k"��2�#�n�낒�:�g4m.���+L�^�yT6�N:����:�E�R����nh�2�n;Q�w	��������ݐ�[�f�����nD
6%��0��r��)�.N�C����{�hz�W&R��sY�r�f��AcK9�<��lW�e����&���uҽK`�&>�S(ۘ��nMR�CF��BF��AmK�Lst> ���wv6�C��S7`|D͵�.Nm̩h1��P�{ůi�{��;,�XN
���k%���"�!�����1.���#��ZY[�WRA�VZ�z�6�P7D�K�ڣ���Y��$K�/u�A��͔�q."�sy��]8Qj�C���.A!��}g]%u�V�]�SR�`��ެ��2S.��Ux�p&�4���#���d�E��ʕrΦ�e��R�^�*�+U��Vd�[.�yM��N�(`K�<���i�o�-�S0���zR�5'E]	�*Y�k���W���]���׭"�yɎ��%fԜ!�����w��YH���K��ɉ��Ӯp�Gj�gq��S�]�w�hۏwWL5�a�-b����Y�N�{�8`RU%�Z����UՊ�><��!���'y��l�b�)�d}{I�s[@��+b��N���ש��jO�M�u{��y�R�(op�ѳ����V��AΏS�Y���ڽ���{D�b¼��´���+4,���1ne<��]VOi��F �줲��d������A���Oz<��^��J�uM��ۺ�J�}�5wU�d��v�.�
��*Yv�=��EWL��������Г�1�"Z�!��m�[�o�a��]:�%m��Z�|��<G.�u�A�[E{�*��뾤�ƫ6�*<v�U���n5�,߰\��q���)N_���j��Z�o@�7,�\�7��YSA<��!R^.q�$��9lM�{�M�˽��*X߲�ɴ��δk�c ÷q�<�s�=��u�$ڸ��y���d�\'_S�i�:�'����vgm��^o*͓��̫�"�H2tb��'d�X�Fl�X�sjۏ*�{^32�g<ݥ9�w�k�j�1�Q���d7Yӻb�ѰU�jp�	x�geӝt�P���b�pv��z��)�Te��C�41D�3��b'�8��/wǄ�0ɟk���I`���*�c1[v�#h�Q`��f�;R�8F0��&\�p��me�͸�us���D]�N��5l]?���U���8>r	�BW����C���M�Ǫ�싞Lg�z f��Pr��,̶n�į�ud�]pb�f�ѷ}����ƝTֲ^t��aq�h��/��Yُ��m��8ծ��;�`�vJ5f�7����hzΖ���{���6/����.��i�t�a�0ur=r0��Zڪ�3^�_M�[bUV�f����fw���b�p��Wx���(+�/�|��J�����Ӽ^�7�C%(B+�ފ�ɮooj��i��+��kI];W¡���كU᤮�c�V����c貳p;�%��r��H��F��aJ�v[%У9^SJ4�e`�lE{�Tݐ��U�E�!�Tv����L,ؤ�sʭ���*t��m��O�`�]\�Ji�Ϟ��6)�ֺ-Z_f>���T���(���Y�7bw�̕�c�7w�I:�sWX0u���*=�]pF��we����	(�8��[C&q�-�����J6��86M��	힫$>�m[]5��Ir�J�/�����4i�̜��K1u�&�]�u�61@�Ü{�`�Q��*�k,���c!�ڼYi����3���2����-�Ń��+.$;+����|��m�T��I�*rͳF�F�oob C��f�%{܋XG���ǈ�E�Ž��7�']J���j䶶����G$"��ݝQb3˙��m�Fﺢ�tu�r��<厦�K?��ѡ���� �n�4��&�(f'5͠�w9;��ԑ��c$w�e:��`�Fw.���Kk%Qٝ����*���gK���V��׬7�L��w	��l��(N�f�Sˬك^�����l��M�[&bZ�D�e��`�ʋ��ɕ�ÔIYt�"��mB�`��p%h��d���-�!ы��o5���=��aD�����ʳ`�"V_ek#s�XJ��m��Flo.��{2\���y�;}ldd>�Xf�iᚱc_d�N\5��h�|�̓��ZP�����f>H.	��(��K�v#ϊՂ�4��Y|��Rn�2�wS�ma�7 �M�����w`��`3D�K�W�'Uj��ֱ ��P�j]]�n��t�-�(��Ҡ���Tc+,<�@d鳎nkԓ7����ǐ��7���GA�L̬�l�.��'v�]���s8!v:y��r>=�.�:��Y�}&�ٲ��q��鷍];P�e�R��tf�ܝ|�))�Xٴ�J��(0v]k��d��7�@�V��Sa�ܡ#4��=�5%�	���"C���>��*s]hm�)Z�(e�5)�9����.����[��ׅ�5l�f���f�R�)�Q�#��R����M��C�W�ܶ�n�z�_,�Wv���:D�nܮ��gY�u�\4]�P����Ȫ��3�QBJ��WM�W��L/j��u�n��t����b�V�76
̒�ay�e��Xxg�j�TU��=rI���9�l��i$t��j�rhl��V������ێ�-��s�]Mܡ�T��=oRIFGu��5!݂1 �|0���خ�!>�Jng&q`G�����'O��m����|'#Y6at��]V�X��Bb2���q�+��<����>��6�meZ�ه-���3ef81��\ea/w�-�9t=��_^�fB&�q�'���_\�t,��J˾�\`�t��vYY��,u!�_-uvv渫6]cop5x!�7���t�}:�T�㌛��r��K)�Ù��F/�Tˌ�(3~v+��́����7i�����f�%T�L����V���X��z3��+�h�sj���]^�.�=��f�N�EJ�&�֕�R�a}��݉���ճB�W�!�u�#de[o[�v��=yVvdm�*�Z-0u�'d8(��9�ͮ�����\�[v4�P�%؎q{�-u۶�Sn���6]c�ڠ��b�=��0��b����:+O52�j1C���]���ⳋ�|������V�̵PI�%J�u�©�c�:����/�m��z�W5=W9u��ZF=��{S4P���fdu�il��w�S�&�it�)=rb޺oDՇ0'�����Ǚ�e�y�cǖs.��3M�����͆��N�V؆%k�����4F#��jC��r�Ӈ;���@�(�v5n+�'s�ս�֙К�}k�
�pȎ�i��9��p�c��D�MZeps;]�9�M,�I�;���t峽:��ҙ&�"��t9Ө�.nKaK�:��[��/%+[Ow%8DAU#w@�J �tiݺ��ec��M��C7KN���h.��G�����e�(�r�r>��6�L�ɰ�{AV��ZM����c'u)��f�SV�\^@���3��O�̓�&�	��;�V���AAQ�D�%U80��Ε�
���	�ٛI�p��E֨x�����#W�;N5�ְ��hS���Ѕ�3q���Y��0�Y�r��i�c7�m��61�P�JVn�w�3Z�V�/	�l��)����:ʺG���5o.gMvo���Μ��S76�����r�gX6Uk��2�kn�8�m��_1p�)SԮ�R��i<�4-!pb՜23DO�Lb��"��R-��[�����r�@�Z�N�� �1�V��&Ά�z�S��>���ݷ�|(��kQ��}�őv��&����f'�F�ͺ�,D���Ӽ����*(��f��VKBe����{�ѦN�jw�0c_YT��T��Y�۰�9˅����C�p$)Һ���PE]���^h/1��I���2͡��iq!�9�*�_L.�'Ф8wvK:m���%��OHU
�)��#R�&.�a��7����P�y�5���L�g��Z�Pۊ��Rw�xm�ԗ�����!�b$k`���`���֧���Ω�ge3+�m'��(�������=�N��
j�CNdCzNDe��º��I�E�v^���p3c�*�l-�eJ�7��]�l��v�=�^`�/[�m��;ޗW��������dv�M�)�W!�
@]�h%m�,����vj��O��;����|^�X"i�e�JFw�L����[c.�U�cn�G���2nq0�\��s�y[.Ku��[o�)��T��v݉�\JYTp��S�P�P���RF,���Se3�+{�X]��ŗ�6��ӡ�!��(2���Ɍ��i��j:B]�I1K�ۺ��[A�9:�(&�h��lg6�ḡba����!�vo�M7W���Z�Xտ��ow
��-,f�m�Sv�X�n|����;B��29��7��z�N����2��3cx�{�NZR��aE�ԉ�YVa4�\�Ԏ�VEjl��r��R�Z�^Z臫�E��e�sv_/���^E]��'rvBT'���rN�ܴ���b���y�h���4��[|R�P�E����{f��؝�V�%�n�d����96�hJv�P�M�����YV	�Vl�6�eс�/հ4E�دWE�-j��`}Վ������B_:s����_+T��X�UҺ������4����%��7(+M=����⎒�0�7�v��Ni��P]�^c��NܮD�S��e����&����;b�Kۇ�z������O��A[���f�ո9 ���`1��Ms�]�;�[O%��v乷�t ��\vv�G�K!���� t�L�%B{7��=��˨je�4���r�Y�R@�1���I�-ն���uZ�=<�i5Ʈ�ۼ�B���햋���j,�E5�6��/�	��5���+P5��/0�|:Q�vS��rN8l��v�t�����1����n_J��HM:.�.|��)��Z��3%թ|&ޜf�σ7b�X5����F��i���
)v����9�d�R��\r���n5h:������l
`�7�Ŕ��Қ�=j�XW����U���l�b��I�E3�NJ�sM�|Mv:L���ڢ��L����}�#��#p�L�JE��%K>q���"����ֹ�Ö�D��f+���A�Q[fΊ{)�}e��eCR�9�g+���`���TяIҔ��,]����.�V�0A'b<D�Vj��;j1#il����*U�3�l�:��T�DN��fu`�u���+��.���`As+4^]*6)7��jv��TTͫ���2�Vp��=1:y���xShD^�!p���Zy�4�Sz(�	�T2v��mj�UK$��"��Fm���v�#��nUf��}q�G�9;2�]nd���b q�80��Ŕ,���I��{�#]���Q���YRq�˕��CS8e�a�a��=g����x4��*��B쪨��j�+�	�X�N�X��%w:j�s,u9�ȝu�'r�nF39\2U���6�g_L����{��&���+{���7�k8������F��c�^��ͧ��m4/z�ݳ�.�\np�,t�9�U$�]���o!�g0Qo]��BA&��l:1��^c0���(�M
�e]p����]yC��,X�ŃA��9{�\�c:^�����R9f���4��:>�ݚg����)��"�Z��@t#.��Zu�b��!9&5x�P�v3eɽ���щ���mL�;��em��ox^��F��/2U�Q][��V�6�ګ�����3���7�R
�<�m]�$�Z�bJԎ�ќ��Z۳���9|�8/�nXo@t�����ʻի��������8
�G)#�W�����Ν�ܕ{�[.�KĚ�;r���Juy�es�bV�*3x�\D[)�d��pm(���
(ْ�t�|�ۦ&Е��Xx;���B���[kb.U,˽�����[]��[�.4fc>�ۼ���1ҷ�)syβZ�2��MĮ_VS�-w��mJΜ��i�'�.��K��eb啗�;/
�Q̭O��1���V_GW����:_��˽Q��X�C�2e��⾏e\��-�r���ժ��+����BhLU�2(��K�J�Uy	˲�ݵ�]۳�������ܺ�ά�f6o0^^ćX������h�؏�r���6ж�z��S.�=�����7Sx�d�\��¦W�6�����L���5�M���N>5��m��������}5������ $�	&������
֮��z�3]�qqd��@n�>������@��nۇ�ٶ��ԥ�X3/n=�8\���P��^[�N]6��ػY2>���y�ҕ�����>�z4IpݺKJs϶�խ.�Quu��ٜ(c�;f�-��&�I��gF+�m]m� �g]z��kh���nn^]vz�;.s�d-�Nݻ������ ���kh�͞���yyI/i1���v�4g�E�<L�s�v��v+t�V����jv��wmr�׹D�2���㷊v�;��9��Z6��e}pKrIƮq(lV�i�X9ɛ��G��ۚ�U�Ew	n7%suk�����ȝ���Mxn���s�p�
��v�\z�븮�f�6Or]�9���ℸ���<Z�z��=-��3��ny�Z7:�ޮq�bU�7+s��$�82��i�s�ɺ���9]�݀yca-G`7]+�]�k�ݸ�;��3��>n0[i}�{�[;=g��
��.l�bz=v��w�����0�G[n�ܘ���[���v�v7a3'��j	����wc�V��a)��F�=�����1DV�Ȉ�I#��f%�.����nɛ��@�����a�yp{mI���#\�h�w4�x�m�ݺ�b�u�j.�e���{opv����Ru/V�����xg����4�Q0��\�öcB\���3뭘I�r����q����<��ۨ��;S�g��ih!���u�ֺѶq��qK�/az����[�:R��L��Q���/���:�;�v�;���<;Yzw\^W'����yCr�s��]��������=Y��tr�yR��n�7\/g^_Y�v�ѝt��,\:�=��81���Oc�ʜɮ�<䮝��=��\������&�x��|�p��&U`�j�T*�М�h8� +��q�z��p�>�pۍ��Y�;��:��������콶y6ۧ�s�q���^��K�;� �x`��ݗ��6�W-�W��9���q��Dm�
x�(��FMٜ�x�<�2I�<<���b]�w+�;l���׮�c��η����
v���%�P�t��q��/���=�u͚����pm㗏V�ݕ�x�:��X�]oK�U�-�rU��mL'�{.�(�3�Y����N� �x��g��{v�H�*ㄚ1V �2 E,,��ثQj6%B�iq��^nz���ؓ����ͺ����%�\ۑ�;mǍ��n;�����s��3Rg,Ֆ��lg�u6��k����B����!��n�<��l.Ҿ]��Ё���.�ݘƳ��6���n�y.�r�����去��q��vwoGM��T���`xM�޺���e��[g��m0�l]�����e�wFF���%�[;���!�3�$�l[g���h��8c��c��v���{\g���Jv����Ƈ�F��q�� /n��=����d�2s�w>%N�=ч���ڥ;�gVx���f��fkQ���Pp���t���w;u�I���\L	yCl�n��m2Z�hې�T�ck��9��(H�����"�<܊rA�g�Yb���-�[����=��M�=��Tv�<��.��9.;Vz���{n8�m����9y�+�����\u!�0<I��r�`��7b�����ud͵aR�Lm;�KD���bs��:��n���|m''�w��1��e¼0��7.��/nr0sc�x;p��>jؔ����F;�+ie�>.M�grn�%/`����:W'F��Ls��2�4�QJ�mw6/v���.��n�rέ���'E]�E��u���%ν�<m��K��M�;�2]Y^Z�`s�Ӻs��.5{,�[���gv�C��+�5p�LbȐ:K�;�Y��m�q� �\�x�wu��\Y�cvkP��nK������M����y��c��u-�y�z�[up:�d=� ��㵭�8��;k�/2"g.ܓe���q�(����/F.�g������lt�7ha�+�^'6���[���=�����9�;W�e]����v4m��ga����6��<�m��:x<<۞{<�Vϡ�i���-ʥ�΂��-��WZ�2㓶�k�]�ݍ����Q�Ͷ��TE���2Q�{�m���^�x��+g�dA�i��:�ra��9�l��5�l;�g�Wh�1��ZG�ssg����3����3nynή��.	��ټ��n��7=�xg�,��n9� �Mu�Iݭ���ګ6y�=�v��������={l6�Nx�;k^Z_\���ܶz�I��)uݵd��'���t�kt۷93�j�Y�;�ۯ]��z`���r��7m:� {m�	�k��4��c>��u�e6@*��l����Zx��ԡ�j\�jQ8�{e�ôm�G�P�t���s��d�'`�s��5]�;�ד�\F2m�U�OZ��s�+�u��8Wюn��Oiqq���8�Nx፭c^j7��Nc[Ɛ��'E�{$����sjබώ�k�t+�ͮ�v ���w<4ts��h���"3u���q�-n�w3�N�cۣ��I��+�h
TDR � [�z�����	v����u*�>���Q9��.�|gx�]/n�l�q�z��X-��ob�r�v�n���)ӷ7gG\�`���m3t��c/��=���1y6�S%�m�p�۷T�ѷY�M�[�1��\W�a�yu������@;m�9�I{Y�m�Ʊ;�	��e�&��v�[3v}��Ng;v탬���W`{h�9OvJ���n1��ė��hʹ8��P��{w;�q�H�c��c����\;����XG�p�:�ù���Art�z�z��gH8]�]�Wm�	�a�P�;ݸ���"g�m��A�]\-�;�m�)sY�6�-�*SsR<j�8,h0��Ox�c���! f�6����睧�N|��(cT[/ckb#]#��s�m;����K����ny��\�8�=
��5�[��rg���[�Ss�W92oi�Z$+��Z�E�c7[ ��N�]���ڄOg'%ι�c]��OK�-�Y�z��d���,����M�eW�ד����c4��xN�n^{�݆�v�f�X�km�M�G��˹��ݔ�>����v��=�]n��1�R�z��yՇ[�X�A�ۚ��e��c��x�@"�8Mv�L��6밆��s�n�܊��86�k&p���=]��p;��m6�y���w:�wZ��t��e��y�;l�zN m�$��8˱�q�y�	��Y���u�Hp7vw�:��y��:r�%�Fk��</bָqƴ=��]St������#ʝ�=�[�%�۞�Տllu���'�ckhk��E8tl�լm͝[���0NG-g8�������ZI�ld]NE�&{��K#@��kr=��x�e�ַ8;3��n{4ckvݼn.�X��W]�Ɖ2-\u��[i��7n.�!��.�z�V�QZۮ��q��6NU���l8ֵh�{Z�8OK�<ݷXkZ6���P�:{\��&�73n��-��H��g�7<n�+��N:���;z홞^�ۮ���Q���ؓ�����8t�5��y�ܺ�U�knf�jgd�c�uz@�J���!�:��:wF.n7>�z��`+\����o�K�h�8���y:�/&a�E�w�6���֞ێ��p�:^�6��B�vSvl�	�ѽ{8xٸ{r�:�����ݚ�Vq�3k�I7}�t�r-��M��m�HNT�I���s�
]#��;�����ƽ[�s����W�s�����b»��m����r)��N� �i�`��T\�6q�wi˺M��� u�����a���:�Gjv��ja:�g�ۅ���;����V�6_9ywu�^���^5�*����G��m1��6��;�74�V��n�m��r̽����Ϻ���b��y��n}Ymn��7�;��t�	�F��ux���e�tn���}��p�mr��a���xL4�������\<�U���1��;f��k�ъӜ���[:k�%���Tr�O!PJ�*��UD�Q��r�ܓ�0q�n���R �ܳ���T�,�;P�ܥ::���dcMu�	�#�yb�s'nGNۈn���u���hڄ�ʚQùz��݇��7�:�j��1��l��j�v3�(l'n]�f4D8&���UQ�q��X�bb�#t�LT������Mtt]�a6�<�wn,=Y�f.�z�k�y{v�n�l�[k�a���p"�8��̀����L<�5�ݵ�3�v�|
�6�6�{��N.H�<��3��ݗ.6��vgt�=3�ZL�<;�luq����Z�a��&�qC��b�eɃ6���ywN��:nR��Mǒ�9�60vs{�{��Sp��;�c<�U��v�tq!��Ws��nѳ� �ӥ;U�n��n8f8ꉮ-�f2��L�5�,��#\2���Ťٕ�kOcm�=�_]��a�u��z	y ����V�Z�ɳ�qz�����v����l����3�`����v�v��WVې��<���nj�l^NPl<gn��g�\]��OA�pt����c�(�t�rp֍jc�a+��/,!���eW�]�����u�G�M5�s뵹�K��v���h�nX��� V/d�x���9{<lu��ݹ @�ump��^킳)��8Lp���z�0��x�=�ك��ݝa�c��vȯm���U�b4
��\�V��*��Y������w
t��n�X6:�\�u��ٛ��So��U{m�n,l=VX��*z�{�Xܶ�mm{q��I��]�}l㚊��"�loc�㡰�v��d�zK���մ�3��뷒�8���˹�x�Ÿw{]z�5���U���ֽ�K&�ӫ7lݵbn��f�sӷ��_�� ��n;��;�쳳��s����w:�m�܁�݇rtqE�q\k��_�]��ZAqqE�$t]�dYYda%G�qR��d�6��2�m�v6҈�"��mݜQebGr�a�[�8qe�u�ی�#���N���]��Q����`t��k;�;����E�d��	�n�ˆݗܜqQ���p���KJ����]�yݝ��rt8TqD]���]�n����J�(*�;�#��;���q��qEGrl��PsjK'm�v��wyg�f�pu	mj8����ϯǽ�һ�Y۴��>�e�Ӛ�*��<���g����N;�*��՞��� :����Gwhx��#��gp�kk��Џ�ks��d �m��"��m�r%�$�7���|;|볶�$qg�WAշn���g���l:�W[���m�K��q�h��"`����" 4;�j"�hr[7o[*F�;K�=������,���X���'����1�q�3���gg��
�1��^چ�p�^O��xf�v�8^��n�v9'�v��j���6Wa��,i�]^�/�g�'u{9�Etb��D&�9�p��7Ds�u�pv�0�J�ٴ�p2���\o<�q����uhy^�\r܎ȼ��l��8�c!جI�6s�lM,pq�n��i��.%�ӫ��z�[�=٥L�2l��"6�N�<��Ҝ8U]p�w��7k�8�n�y��d�:�� k�L�T�U�R6�A��)<�&2YR��zj��v�O�:d���>��\{5���6h��H��,�Gیx�K���n�.���s���:N����[k\��}�[Iύ�燆Ӽdت�;6]�@n�7�<�D�g�N��ꍶ�;m�{u�U�n-m��u���%W�㍺�����xט��k��M���Z�6ٱΝáG�GlG�C��f�cu��X��ï����:��<܌���m��S]�̚���t�� ���FQ��/�=��k��s�������T�%�u�ؑ��X��m:���a�c�������I��p��]6���Լ&�{r:�qg)�ٺW��ѹ�޴�v��c��算��� \���<z6��wmuK�]�¦�u�z웱����{�q���ݴ�|M��vih��l:7ssǆ��h᱓����;la������a֍�:�Z�֞^b�tm������lp��gv��[(O	�=&���q��.'���J��B�������0|�xں��b[��{ƺ�D�m��Qx6�_`8޼�Om�����j�Ӛћy�(�p�yϲ.C�o�ݎ9���]��/c�s�x��ݸ�'��z�y�gv1��<�c=�+�S���v��s��w.L���{{ �;��aϽM���lrZ�zl��Ʒ��e=�ݑ�W�ۜ�AƂ1�܉ ����D�G80�y�=�v��ceP�<\?�� Q�ټ/z���Ǜ�@�� U��(]x/���p���8h�<��A�d�Ay\-����yUɽ��llo����chy��2��s��kJ���2�x{đ�f��^7��n�� 햑� +��:����t	-�{t=��+��u�*Ք*��T�R�.}�Y�,����@$���Tzw5��np������]y�֖�H�uճ`,��%��qQ+�7��R�Pʒ�Me�n�I=��$�{�߮����}b)�R4�	
�l'Kl��\ĺ��JrF��J�Y$%n�(�ZC�[����R��T}5�O��Y����0%ڕ����� �-">�*.9`�� ������Ll;+/k��FR��c���t2]eP��2��l{�:�����|�Y�M���K�D���kj�l�ҝT���C��sk��sz��Y�<I ���À�	�I�H=��e�Oݿ��MZoM�RJo�� Ӿ�9e��͗�{�B��J���Ҫ?
��st/Wu ��`��y��6'K=�����m���'���4��t�u�D+�������6E�H�O��@j\��>"�[���(����� y.oᥖ$��oգ�yx�g�v��w^7^y���783�mс������c*<��x�7
F�}�&����~�?hA$��7tػ�Vv^�cb=�Qo��t�Y�c2����M��9��@v��o�׀���a|G�9�?���wA �8�F�W�R��Y�C��Z��(eg�11���'�5L
!�݀yi�!�Z�w)�{؀)w��/���a��0N�l3��w�b?m��XX���~�ڍ�����x��y��5�7���I��ѿ'�n�ő?5Y�4HTI���K3�ξ������S�P���`
{�c��G~K��ޥ����%o�=�(��nz\��i�<�&}�~����\�ǒ7@P���B��ڢ7�Ga�;�T�5���E"-�v��5\S�yNb��k���CNr�*��vY�o��3��N:���ݎ�<��@S�c��V+���&콋��ۙ˾Ι:��b�Y�e��p/�b���b�UǞŬ��%��P}hR�n�q���>�εn��y�N=�O��ARU�f��4ޚ�z}�m��Ŀ��z��@=ع��(=��G�O_�h�Ϭccۛ�X��1�x�dG���	�H�KÄ�fy���䃭Gu��رSl�jlV:A�-�sN�tƮ�7E�v�%Y��C[�L����K��I�ܭQ\���
|���ԿM�9�s1&�.��	��
A�Z����wu6pc��g�=��9�� �n ~��3A,D<��*d�l���8�kr]v�q��^��g�{r��d�+�b�n�[	��ys����Ky�_sy���{��/o:0l~!T�#������*�m�����B�a�!~��- ��uӸ��{��	����L�I�H"wޏ���:D�fQ��رe����`>���h%>�>޽�q�	=ޛ�OM�����k8��>�,���G��v���S׸�� ���Р+����
�I��ϟp����6uT5d�����*�������tZ3���f˂��5n��C|��Cɗ~�<CׯH-nk��(�6����5,\��\P����/��M��Ѓ̂�]�}g���
q�eC{�C1���"���ٖ۶6JjͶLv�/\�{NC�2�R+d�LU�N �"Q��=ֺ읃r<�:�Ͷ�u��z�u�cu���@��.�.���s�OF�[��<��m�;���GS��v���gl].Etcme�s���m��m %����V�w p�Z{WNk����x�m�7N�qəᗘ:���awnF93d��!r��4mF�b�!�y��LG<F5�o]tXy�l�=\�OR�"ł2���BoA������{�=&�'�� ���M�i��F̪?�u0$��K>罘��^��P#�������(!�+s�V���i �w��>���t�E��,������֙-��*5ida��w�ō57�g�4���>���� ��B
{�ءW���^ʅk��5uDU�u���V�8%��	�͏�> �y�@Cˮ_�hn���\F3��=���	XmY�9�����������}s��^�߬
yӛ� +���	��؍P�o&���E��ۺǮx�WްfC�՝��Ak=����3�A�W�!f��uAC/�7�:���ߦ��oҙ����c�o޿w�I%߽���p]�>�428���ֳ��Ic���nu5ͺǈvr d@�˳�<+``��?_0��߻���3x�U��W�e�Wuֻ�47��q�0�O|4�I!����I'=)�@V.�j���������A�7��r�1���� 
u�4F���i��;�٤�H�d� �?�=?���sc���������ǻ��\i�f�$}���|I?}������Y��e��zv�.�%��"EU�"��ޮ�����vk���!�NzY S���	9<������D��OY��4T'*�����`!��x��-��8�6��u���=="�󾾻���k1�Ū>�n��<�A�_�7HT������KE{���I�O6)�HK�B�+>���no�S������L�%ވBI�v�A?K���$ŋ��5�7�}:Г�ʌ� ���߄���w1�2w653*{�GPΪM�=�5=�U0M���{��f��h\�/�̂���q9n��˥9��s�����Â�*a�ީVJ<�_T�?s��픐����I':S#	��M�E�I���TK$�3=��{�7�^6OH�{��k��<���T����0Q�_A{��Oك	%|��c�W5y15MS��s��� �~�
�����|��7AN �`V��(Gq��]�A�%SD�ۦ����	�|������o\� ˬ_�}�����:l��~���	��i$��=�M>�g���1,���\T~y�����k0�벫#ϧ=���7/�������zo����@��t�	����adW�6��+�y �kN*��������i6��fh$o�e;%7���!�I��0h&�?n�Z� �l/�R`5��#K,gƷ�{��	$Uy�?��|�1�rܵ�G�d���C�+����"^[�����qg.:VLz�
u,�ۓ^kC�GauI٠߳�5׊YT��f{Z��.柷՛/��%9�tY��c�n�Ń�w��z5� �mY�XT��󾎨���\���>�{�>�w��~߸�$}Vz�U��M9k��rTM�Ϧێ��]c�Q��h�]5��$�53~����E٤��9X��I7]=�W�a`�匐^��ڮ�Ѡ�G���qS �Y�*�h=Ҹ�S���W/ۡU7%��$�w���
�2��v��g��m�x��k1�r�BW%VG�3;���n����Ĝ�'�$ڄ?nA��v�ѿ~��]Ev��vO�x���ֻ}��'��k��+���?��=����d��T��~�ѭBʩ�׶�@ <���t/o�Ҡ�O&�*�[��gw���m���7n�+tB̉�}�1Gw5Og�2£�z��`ɏ.�J���/��K>=wGұwPʣ�{{�}�/Ui���|�W,�Q��l�O�;���j�ggGA��y�5ç���c�2�˶:���\����ƺݮ��܋�Nk�6�6N�дa7w� n׮��3��]�`v�G-�uî��:�M�nX�r�mٻg���a�{]]�n�:�ԣ�j5���3J <ܽ��S��+���v�]���7=����G:�Ì�q+r��qvwl���q>L^���-����6)�6J�{����,����L4�.!�Mƿ?{����U%����}��16ۛ�ύ=z����M�>�ز^�@ �˭�!A���7f�K���Э��%�wY=���ޜ'�G�On�I����N�b�f�	�4�A�Yj����@�����r��pNL#~}@P&�h�+ϻ́�b��8ټyYv[��Lg���� o2�" ���Iq�ze��>��-У�y�p�F��h]���	<�}��7~sP�ݭ�C�v�H�=�	����Z�2������y�܇%t��P��s`׵pNwe�q�m��ok*��HB;��B^G�SD�b���c�s��C3�ɏ5,;��3�>}�l�c�����Y˻'-���� ���bWej�-�G�M;�a�qkH�F)��c��1݌�5t�[�p�\^ej�2h6�E4(�ڕ�s8�2e8�@���YR�&�&>����Y~��H'�?{��@P����� ^�����t��>i�8��Q��}ߵ&s�u6ۙ�o���c�=��I�H&林o�h:��	���U�ѻ�i���Vz��罤	��4h"����9�V]�8���cS�da,�����}ōN{/���q�'�$7}7t�@����?��<�3�Ⱦ��k��}�!�$1�g.�s������m��ZE�3��=�e�-O9��9Z:�����i*R�d�w�/�n��wޙ�A��0�xOfA7�6WP��`dշ7@$'���B�@�5�w��+m�ٗo/�4�E\��$����[���m�w�6������6I9m�= �j=�$�g��ǹv���u��`����x�G��Z�M][��ǚ�P�b��)�
+}�ԙ�8�Hۧ4����u�ge�t����q��Lbj�\q�s���rr�N=�W�ه�k�}`�f���E[j�4�(�m�k�B�����VE`�W����"!�bZu��ǣ.��}��MP�>�M�;�oOW����+�e�ܗ57G�S�0�b��i���eF�7.����1��]J�K F�k��1e�ʎeE\�������U�t���۳r�q(u]ه�����*o�NU0�8UK�䳌M���)�LM����^���R�enN�kn��2ڻ��3�����Ĩ�y�J5�k�fI�ٸ{�X/{:���LcWjep�Was��R�ͻW�Jr�m��Ꮽ����,�DYVv�2I7��,�U�u�O�,pM�:n3ָM7�b��Qm��"e�7��]ҡ�r�*�9�9ux���ǭùt�Y\�T��]�
�D���	a����6�n)�w��SG!k�-
U%Gr��jljvgL�}�L9�����s�v�`p��NӴ��Y�������V��=��>�mo`k�Z�]N�ts��V�PxN����'$s�ڐ*�Ɲ�a�sgS�nnH�֊.XN�w�}����mBs>��YnV�N�X���a��:�s��ZUV�	���e%r�5F�T�D�g����N�-M��q�v�N\��1un�z�C���6��-��ϛͬս��q�bƸ���/\��X�=|��8�J.���3���i�U���q�m�8.+��6ʋ���8�ΰ��$�8;��βҸQ�VgQ%ZU�TRty{�#�䣎�m�qv��β�����$�|;��.8��g/k��;_k��ˬ$�D#�3:+.�y����n����:H;�2+�vrE�qǦpy�oj�8��b"]��{ڻ�"�(��m\Y�m�i�G�Ŷ�:|�VVR]��t��:��Օ�/k�n��wKm�iQӇ%ݕ�w>��.�tD�˳��>ugs����J+.�^�'v{l�.�.����:�W��n�{4���6�}�T�!X�RB��?l�P�֦|O�>o4��צ��A���k/��ED�'�ѿ��ڃ{ѶkZw`�;��m�]햨��>{wo��4��������	�;����w�9'7���i��\B�6[/���7j٥��3�mT(�,P���,֐�nk���K*�K���3M���r��oM��ẅ́��{3v��n���*�p�i;�h]�����������K�}z2Cs%����?�5�n$�L��$^fI���+�]���D�%h�%T�
c� P��6%%��Y��пsϐv��t=Wݣ�#*��NZq{c��ՌYQmK�P��@| 8�͊k��,��I�g��>Vn2�ԍ>W�L�+%S���L]�P�n�孺��Z�ҭۭ=��r�>���Un*�q'be����_&��v��V7�8�Q����5���
�7��;�S�y}�������7��tk#��y��v|�4~ң��wXq˧F3��L�W4\G���S�pB�����7f��>{O��/�M����L )go�����9ea�|���M����16�_G܂e�;�-��:a�]�==z��~�t(S��t���w�K���U�Kn�0l�S���Y���˩�(,����t�]���3S���٦~'��n��oۿ�q"G"�]��Ea��5��ǔ3%�7d�A?2������V�%�:r��>o����ח/��G#��2o��cm�[Tr7R�� ��6�R��'����k�]S[�m`Cu���:�ӧ0�u������w��*����(���7��Q]5�׸�x7�&xo�_`ѓ%��WC��*�ot�����(}sl�9��θ7�n�E	TPK8�� �2B���j˶���{=�X�]yz��B�X�[���4�yc�3�1�����xڗv���l����>:x��v1��]�.^K�J�V����W;'<�c@�˞����n�hg�E�7j2|���K���k�pb��]nk����\�k[k<�ω9yr%�E�p��Ŋ�m��E�o<���������s˝]��;�qWO0�Qª�M[w���U���?�_� Y7Ɋ@W�c��h�A:um��Lz4���%x�/o�HV~��[��^� o�����I��T��n&��~'3ޛ��G�V�@��<�ꐫ�=�[�X��l�)b,�s9���i��ƈ� r#v$=�՗���(%�y?�M��3��:���T��nc����tJ��р���ٿ	����ω'�'��bnT�1^i$��7��A�+��AB�ޯ��>;|鹏|�~����2��K��f����&$~��{L�3�\[����UA��D�b�����pUe��m'�v�.���v��$�D�������6�i��}�H"�ո$�[��w[�����ԝ��$�q��G�#�P����wE$���Ѥׇ:��LX2��c��S�r�Y�D�1<�e�����u�A��*�5h�o�v��V�Z���&�4��8�r�%^���aP�]��o�*�z{Ѫ9��`Ԕy��
8>˲������ۤ�u/s��ꬿz;��?r�>_%������ˇ�"���[sz��2��\��}��7�v�|�`ҍF�z��h�����1F���ݴcF4F���f���œ�J���kr}�cK�JG���%i�`Cۿ75ǽ��7�ٽٌF����x�G��~�v��O<�}U��{}�o��#������H#-0# ��Fz���4��D»���h�s|Ｓ�r����1Q��hrN��+���ڸ��t��YS���n��~\}�rHA���i�ɢ=�7�A��b�#FW��15�(F+��Y�L���w���NU��An<߷�A��;"2��R1��G���z�[����V���~��Q��j(�el��|��q*{�ߩa�(�1F�W��"�14F�4Fw��-�ҍF�y|�}>���ە{�%��0'���5ŷ����r�0,dh��=H�!����z���Cq����=�����Gw�|},�����Fm��X��`�ybp���)y}6��Z��Due��,CBI��4;�:��A|rN9��T*7ݹճ|�3�1���{��cXҍA��g����D��϶�d6���cF4GϽ�P_ML���9�b���h�w�Q�cJ&�&FEw��1�����4q߽����g���o�w��D�~�Ԍxp��|�A��m��nKAi�����f0#Q��J<�w� �5n�{V*a�b��ߩэ�&��۾��b���(�y�o)+��7��w�oZ�S.�d�<�ٜmŶ6(궧�sz��7m;��mUXQewN
��?u�;m��֛��ƴ���>��y�A�H���-�lCx����R����o�5��p�����ٔ�kQ�Ҍ#���1�&�=!~�}9]v12�iF�������l[���������;���D׳�E����C`E�_=f1���w�o)�PC�{���5�U"��G���Gõ���rm�f�oZ��b��Ϩ�c5�j4������KL �A�4wۮ��r��r{W��|�h�Dh�D`o�稶,aQ�ҍG~�w���F�?)��=��H�Q��44^�����S�Ԏn�޺�s悄�$��r���A�n��� �����C;\�����f|۬ޜ|�7�X̎���� �S��%�,#����#抆,�8����G�뉮�W{̑���d>�+ynbX<���(tn�Q����]k�Ҍ#�}�1�1F���{X����h�cF4G���(-�LQ�b�#G��v�Ɩ���=�����Y�1���q���syH,��=���ݧ'��~_O�~_+Hک�T�V0L)؇����cf��;v7� t�=���F��~���U�1I��b�s����Q�Ҏ���4��&(�6���֌hƈ�5���>F1A��}�1�҃Q�=�z��k�$/\:t�X�V�ݸ���#G�粑m8�{Uߦ���r�w���y�/��A��G
��-e��6�3�����`ҌCa��9��ϵZ�u��W�.�1���;s_-�SC����!�r���F��F(��;|��1�l����s���W�w��[F�4q׻����Gy}�#��w�־�ss{4kz� �u���>���|��o'Mt�(�7���E���Q�b��/޴cF4F!�7}稶'wk�XSKMZ�������5H\Sx��ۮ�)�Ldh��z�m�D����-�eg���N�M�w������Wme����D�z��F5�(�iF0��=F0�(��[��rt�o[��oW����fX�Ø0�����c�[�̭ �ӷ�^`�U�Ն����km�?@�Ľ��iΰ�+78T`�7���y�꯳����\Q�\v�6�Lk�.�rn��=k�8�Ƣ���j1��/Ĺ{��m�x��N�8�3�|���b֍����]�m����q�X��(vW���m�n��8Fr!W]�O,��Bڶ㣫�I�t:��{t�S�\D=��V<���@*��%�㍇[mk�����ɩ�j�7&1ʺ�rg;�g��մr�n(��D�1����Nu�8Qi������<�om��:ޱVY+�X�m�v��~�zڮ��K���>��Ai�LCb��4{��h��iA��6���-����������syH/PC�Dhϯ��[��G+۾�no{m�orZ�b�+����4�_^���:��s�Ը��n��KL#a(�����1�4A�1D��s�c�X5U߭���V��v���{yIX�0=��wC��6m�M�l;����h1�"~�v��A��(�%�+���5����/� �d2&j�{�R1�iF�Ҍ�s�,im5����rI�i`ܰ�(��4G���A��<����֯����q�#a/}�(Ʊ��20%�߽f0124q������H7�]}��~~���6!�F�v��Cy��Bۜ$���޵h1��gr�b��J>�7� �7�l�9Z>�^��Q�1F���ݴcF4F�4F(���Ō#JF|	���}��D�zODhe����Ȫ��l<Y�����Mqv���qĆv{r'�g���4�J�S��'QA�U#<�I~hzW��bx�A�!�/���/��#�p�z���l�~��ͽ�[πƼ3���#Ɣj(�0�w�ь1�4CG�'5�P��oR�hƈ��o��4��Y��O�T�!�Ϫ�;����^_�c���mQ��x��:�#+&֣W�c�T6Y�M�����/j�c�WLn�܂�ԡ[��r(�a����[��_f߃揷��Ɣj0 �����f01���Ƃ!�����!�(!�Y��UvMeC��M�>.�b8���U��m�{6=�ܔ�0>�Wh�!�Ɣj4��{Q`���F(���g��w����G#أ/���c؆������Ԃ0/���hއ��orn�bG�ݺ	{�w}5��h,q��@9��QxADb�^�}h#-����z�me��I�g�m�F�>��a��4Bq<֞m��F�7-��#߳|����1D�4gy�����W��՝559ޮ�6���s�Ql�A{���Z�؇"=���4�u~�K��s��'�2���c�����2�%��[I��Z����-����ѝE���d���_�ż羣�5Q�4���������0��4Ow��F4`�3��d�}G~F1[/y�Q�X�F�MF!�����kj4���rtv�R��K��_��`��};�Ϸ�����Q}PDb�+ܯ�e�d`F��w��F5�(�iFz���*�����3ηY~
��(�b�G�'5�P��ze�14G���AcF���F�{��0kP�203e���_�g�Z����+F|A����
r��q�W��6zx];�V�I�E�1i{�[�>ڽ�(�,��yVj�ę��V���<��h#�����jqA�sԌx�GU��z����ܖ�2�/���1��y�5�3z鿀�\Q�o\��E�-0�a�D�{=hƌh�4F(2�ϽF1:��o�g����MF�j=U��+L���u�m���5�����;��1���W��h��%��X�����R�L�0#Q��ԌbX�Q�T�� q#�[?O�6]�[������N<�㚋X��������Sp�q��;�"ۃ��p8�W���<[�O�C������|�h�F(�4g��Q�X҃Q��稶#AY����ԯnaδN:��ADh繝�[�=$3�u�>��[3Im��_��>[f1��{���9�X��n��KL"b�#h���R-�#D#es9�1�m,�-gx���U�^G�]w��+Z��i!yLY'Gh�-U��IcCһ�v��A� s�^Db�s��}��g^jo�޳ﺂ3��0#Q�s��F5�(�iF0��=F1�y�>k�oN=閌hƈ������=��o���Z�N��y0�Ch����cX�6!�*���l��G���A�}��^��2����e|n��/�f��6��:k����i��ԩ�Y�L��y�t�'��sF��Q��$�X"�}�{&�x��eFOh̺�_P�DH�=���F<�,�;��okf�nKAj��-�`F!��~��(���n��������ZbF�Ք�h��#Db���;F1`�4���(�~��)+f���f���#5��z:]�ݔ�1��������EWi��
������孏d��o}-��F�s��4q��W�z��"H"1�_k-#A "=��M�o��?{�.>��kQ�l"aW�v�a�Q�C�Od�,T�3HkI��/~K�J5�I��\�ٕ[��h���H���Fd`B����`bdh �߯��Az� ����<�j���s���|�q�A���8�;$V�l�%��������餣ڃJ?���-��1Fb����ۭa��w��Q�#Dh�Q�}�h�,aQ�҃Q�����f��XN�W]�U�Q����f{�H;�ӡ_5���|�|�@9��(�PD�Dph#���Z�LȘ��;��cO|�}o�i�g�m�F�w�c(��?�;�H�ӄڴcF4G�wPZh�C�F�{��0kWG��	�����&��#�{�1����AƂ����jp�$";��񠍤����׍O��V��S4����,����A��k(\�H����tj�>�n�}uËY�K�:��R�=ϑ��bN	�R��Hq�����r��w+��5�*<KM?��`l���حZ¬�.��%N�Tt�̬����R�1�BU�J���5]��H&���Xnʽ��&f��������훷���8uuy�Жt��Շ�D̤��B�lQŨ�	b�����Q��K�-��PC��qj5ɗǻ��,��*4%5�+ʶ�ս�)�[3��{J5�+Y8Ek�I�iز���l�f~���;�����砙x��9��}��\��tQ��"��G1��L��P�$w͌�A�����Z/��-��d#�Ou��i-+��U�|=�F)���ed���lwm��*�p7^��wE?5��H��|=��\�lwj�v���j�o]��!�Lk�m�D\���7�F�V��}�H�8�.E��XȻ���]��,쎲��|t�پ6��1�O�Խ�(KWsW�2�h��u�(�H��Ѿ�����䫁NӖ���3=�Ư�l[��)T�T�:�xeóH�������<�S�@`"��9<\k��n \���?'��fvb�����e�����V�p�Ĵ���O�V�s�KP�W�7$����4�	�4zD"�bә���\��͛wT32�'}y4�9Tb�(�\����*�ҫ� W��J��Y��+|'Υz�ᵹy�����4=��J�;�cao2pUV
�J�oXࠇV��Je�,5h7%�����ˬ;��Y��l��+�N���;���H�k����(���8�y�I��v�dt����{T]ynq�QבW޷�>���uw�Iwy�yڕgVw{jN��:����}��:��gY�ܝ������grD���M��㮎�����Nzh���^�IYg�]���eg��(γ�p��{��:#�����[���R\����:;:+�9.̋���Y�fVt�fm�mt�\=�8:";lT��mn6�ze���=�{s��Nyם=�kq�u��Y��q�Yyvsm:̽�w�N�ᵝD��4���mf���Q�u�<��'VdW����杳�=q�ӷ=JuMsW]۠N;q�y���,u�]�T[{=�o�ZM��N��]g]�*�H\q.;6Lv�+g��3�s��/C���{v��#�5�s�gמ_n��{z���qn�^xC	u�n`n�x����әUϗ*�^9�F�]kF�K�f�t���e�j�;���h;m��v�A0�z�M�z���vW:�<G:�ۤ�shwktJE�B����Lr����gv+���)
m���;�X۪iz�Z��=!�C�_1mۇ�)��{60I̒��/�G�pƹ6q��N��b��SWV�j��],��d��0ܼ�{�����O/3���2h랈6��96ܡ���ӷ��z0��Jm�݋�8EiS:ݗ��X�������Ok���o=�b!,��<�D3��[�ic�]mí�1�0��u�I�k;��\J�=�8�]<�-��y�8�[j��hݵ��{uۨ�{vF��G�&�h۩ۜ�v9�z��Y|��m�g��jӋͳ��ʯS��M�h�7M�;i9���t�N���n��8��te݌����r��L��N�!���n��䧢iFɝ������{��"���\lh��!�x3�s�L;$v�c�(#����[K��3�\)�N�q�iΌ@>;0;=:f�s�ՎWs;��]�*vk)� $	�X	4� Gc�(4�z�'n�l���m�s�(m*s\捋��;c��Kջi�ègҭ�u��v��������<��9s��rW97��n�Ŷ����R�p��;��r�v�'�r3ƣy�8�:%y�����u�#�N���ۢ�͞E�u��˹,Ym=u�W��&��x��Ƶ��n�����t�c;���{��\�/Snr��y�I�9�
p��\���'I��;nl71���,'h�1y�=6��6第��mpm�@��[
�2�����H5����wE�n���x�<݊�2Ū�Nm�����h�9G=)�9^�3�̂�ڙ륝pd���7:�]�7d�;S�m��2Iv�齜�=�dD�&���������9Ί{�5���]���9\f�QC�^9�n�=Ǫ�����ۇ����7wEZ8�r{ �s���K*d�qn�x^�)�U�yn��Q�M{\��O=��|k�=�nշEzu�&��d��S�f�w  e!�Z0�ʥj㰈;�n2���Z�]��B|����g�<�"̹�'\��y�T��!��3������������ݷUZ�4���5����1���DҍA������!��=h�!�o]�h���9�}E�[7�}�1��6���j��0+۾}��r9����{����}۠���#/o������N�ծ�{�ܢ�HA�o���e�6�=���4��sw#�w�1�i��;�Ϩ�ޗP��7�;K�L��'�?nv���F!�_��R-�lC`>nz����u��`c#A�CsW��AD�G���#���}�ё�kF����[:1r�Ϩ�z���}��w�}�i��iG�ݔ���D�>�3��h�h�4F_y�-�Gך��s��Z�p4���iF��k6���as\ܛd�ѷ�4����}���c��@�?`�C�yg�T���6np/�:��G5��AL���D��3ԌbXҌ"a^�z�a�Q��tx��,����>Uǡʉ\���;$��kc��9ڲX��M\3���إ��*������gz&zp�^G<�}��SF������v�kQ��6�g=f1�柦����|�cA�s\�
��=�g)�4�-��zm�{[7�rZ�LZ���1���Ci���t�������X?�n'r���po�{)B���3�s��lo�
}׫m�]_�1�:���7~��g}j����i��vs�-�YZ���[׵ݠ�?���D���~Z1�#D#L�g?(�,aQ���������x~Q�ڽ��j�����曓km�`|�=��Pbx�A�"^�z�bAƂ?}�>�����K��gS2��;��cXҌCa����"�z7�ֹ�BnG��h�4G��6�Ͻ��_���F(0���cX҉���d`J�w�c#A��u{A��k�wc�m�|!��{��"ߚ�<z��r=�kOs{ޭ3����c10#PiF�iG�u{(Za�����o��bG���"�:�#Db��g=F1`�4��iA���^Ҧi���o���_?e�5����u�t��L���㝶_g���.�5���@�9kVSVޭ�p������K�Q����x�A�") �������#��G=�� ��g%e��4�=��6�Y^�z��cJ5�aW3��`�5�m�d�=�M�E�bh�;���@�1kyF���/�]�[�H���Q�F+����!��߻��
��'�t�6��G��r�Ǎs/���ǽ�h���h#,�_{�c1��ҍDҏ��즖�A�0�Q���x9��j�eܯL���Uk��S_(�hr���4���F��`����$�iԘ���9`�gpv�����4>��0"����q��V*wW)��������h��0+��QlX�F��(5�oIP�`C������G4ܛ[ovcF�g��S��Vk�r��h ��v����!�G��oh)���g��z��4���f��u���[��%Z�]%m!�8��cӆ��W�hC������n�ϵ�����k��d`{���l�A~��*��$���=HǍ|����t{^oZ{eԢ1�Z!�^U�7��v�a�+ێ{\q�ۗ!�۶x�=�I��%��ރ��njh������<��_>��5Q��Q������F(ў�z�m�>����-�W�Q�X0�(5Q����T���	s]oN=j=�Y�!�v��H�!����L�M�_��N�.��AA�h#�ܽ��!����z��cJ5J0��q�>޻�>bG|�܃��nG�h�!��h>h�(�1F�����4��bx�?��a��=��֪��c���A��^�QPC�3��R-�4˿C4����{7%���Ū������c�*��n��m�iF�iG�}��Ҧb�"b���zэ�"h�Q2��=F1?k��Vx��I����y�G.�:�zlZ���b��l������s���F�S=RY8%�}��~ݷ��:�¯}����+;Z��� �4��(5٫�T�0'ۿO��{�z�[ovc�+���u<h �	 ������%�W���e�8";h#���H#(`F!�3���(�iF0��=F0�(��}��w/�����~�l����t'k6Ǆ�
����Z�v�X����B��MByg�4FN����?iK�M�5�&�1A�b�#E���15�(�`@d`J���cn��Y�#�>�4q��sh)jqA(����F1�u�z�M޷�h1����>���&�j���4��W�Gw�l�ii�b�#h�}��0h��0*��QlX0�(�iW�>�z�(�ON*�ӗZ���$r>��� 똣Ic#E�3��lD$��z�bDb�5�H��{�������g��v��cJ5Q�~��1F�h�I9�$��mZ1�n���}꩛�nu���|G�0�Q0���(��iD�bU��ٌCh0q��������o���"4{/=H��s/���7��h���h#}]��6!�Ɣ~�e-0��f��k�F�D5��֌bر2����6�F!�wW����V��L���������2<�����A:;P����؎�v^����T�f����<{��}q^֪�&=��鱘� �z��ﾯ��Rs�&y�u�����**��Ol�ˍr7r6���ssg�{pY�^m<�[n�c]�ыe�,u�������L>�s�1�lo:�۠�=A��x;�4/T��z��nɰ&�Ɏ79'/Y9zq�j�n6������y�a'q�/Om
���K����\v�f���fn�]1�|�Ǉv{%R2�y.�l�5�ŷ.���"�H���t[.R���<��7�\U\�f�9�.SF��n����,>m}}���٠�mz����?#Gs��x�G� �����$�#�~�h#)��َ{�9���}�"��ҍA�F���1F�w�2i�pܚ�noT��`��\�Rh�a�3}�2��gټ�m��;�u�iA���#��v�`c#Ah 8��^�R��&�wU��G��σ#�O��(.�U�����x�����c؆�4������Za(�Q���f|ϸ�UwZ��U󨶌#Dh�Q���h�!��j4�5���T�����]m���Ց�i�����{g5N����Z8�6}��-�yG�8��� ���j3�s=Hƫ�^ٙ��^���gk_O%�������6��'sC��٣jэ4G���)4i�0�Ch�~�уX�|��k�HLX������r�``��G��{A�D"����R1��G߸B^}]�{�����Z#���q�{�
�ܻm�P��LoN��d�%d�ӵ�f{𸼣{��7����#<�]�v�f&j&�j&�~�e4��&(�1F��g�уDh�r�ŗ��#lZL�{�Q�X���(�����`Q��'�ֶ9����{����}ܠǍq���O��~]��y���T���t+e�U�S�I��n��n�8Y�3n��3[�]=�/ ���4γV�R�yĐ��|�y�/���4��n�e0# 0#Pf~s?)�(�CJ0�˸�r���Q���C���9���޷�oT��cD~�sh#&�0���R-��F!�=̛���}SnO����X&F�4q��^�F!�F��3ԋx4���,��7��n*���8�?_��4��+�okڿs�p�ZiF�Ҏ�U����A�0�Q��{=H��h�C`z�ثO%�+>>
i|�b�j��&i�=��ٮ1隑�Ց�m\�P|<h#�C`}y�QyNo�>�o�w=t���7�w~����Cj3;��#�ҌC`v��`�.��&��i�]��{�/����n��5طY���m�O����8{m��>�lN���9����5�6�Flѵ�u�n���y4i�0�Q�h�~��-��Fd`z��24�_�o|�r���X��Z��|jp�$"9�3Ԍx4��C#vW�P�$4����5ԚHkI�l����!��.={]�cKL �F(���=h�!�cDb�����!��j4��_�vV��^>\z�ݥ��}������l6n�``���}ܠǍq�l^{�^D�Dq������Y_�?m��M���9���:��KC�7~�Ho���j�0%WaF���3y�s���fkw[��n���5U����I%����g���?>�z�m`ҍF�`~^s�a�h�;��M_�z���h����3�k�wW��r��S#a+��Q�XҍFz���A�oh3vf��ՈqADn��R1��G{�Y��5�ǽ�h1��������A��J?�oe-�߽�z�ʖ&h��;yhƌ#DM�����b��iF�ߧoiRf���wk��v}�U[�l
\s��">M�ń���%��ݶ�=���1<9�)%����j.���|�I~hzY~��cƂ8�6ם����#�=�� �)0#>9��=��;�}�t5�;���F5�J5�a�s�cb��~���C��Fգ0h�'oaI�lPa��Yw���=�{�>kQ520=y�Ql�b�����D*�g	>ǿ_8�v��#�{�af�ލ�=�ܖ�2�o�v�f�6!�N��[a�0�Q����}�ֳ}ץ��G�Dh�Db�˾{�c!�iA�҉��;{J�����=�lݘ�����s�A�re��=�6��1R�e�E�A�n&�9�r��C20�����|8�tC�m��L��F]>2c՜�v�Y%�V����t*�!��~+�8��	��&z�i�����I���u�}�	�ZDo��E���~� $��u��Ҍ#���Q�Ch|��4�'�%�iK�H����ҭhL#F����"�Y����`Rd`Ng����dh �A��h4�:�$��{��c��Gﳮ���k����w;~�}c<�^(Ǟ�͹6���x;i�5{s6v9�a�U\R+m]�u�!��\�����>�-�L�Q�o���M-��Q�b��{��cF&��T>s�b>b�2��ޣ�aQ�҃Q����C4���|A�=3P�n���F��ߨ1<h#�D��g~毌�ٜW߽E���4�����LȘ�3��z��`4�Q4�}�����5���|�6�o����oDf�T�h��{W���LQ�b���}��������^g��Xs�������N1��}��tAD{��R1����C
6�ލ���r�i���2�F2�^�;��}ܼ��u��Q��Q�j��1�1F�g���cF&��#L�����-f}�~4o���F�F�j;�ˤ�e07��ƶ�ލ��f�24s��R-�lFHw�z���g�ML��莽�p�۴e�Ș�3��Ԍk�j!��s��[�Z��^"ԝU~s��#��
g�o׎�z���#P�wVF��H���;�P��R���r���3d	�^ᝃ뫰�>^FnBav]I�g�Vo���%��s$l6F+[M�-��BY��-��ۡ�h��#� ք�m���Ө���%��g[-���Z�&��r��97<f�.H�V�::�;���z���mz�d��۶:��1�ݬ�����5����j�at�� Z��m�g�����g�b\��b�c�lf�c��R�w>|M�.���e���L��lc�� �.jdz��6�!�	�"�Ǯ��%���]��%�wk�Ga�9Ϭ��cpb{;	9�ü6l%�����=��oZ޿H����3ޠ����a�џ{�Ʊ����#W���c
�_y�ʽ��=�r���$G�Ͼ�c�s�Yji�[��jKA��ż�~���6g1����R߾���X?zD� 2t�b��x_I�Y�χ��б� ��.�H,��� m��i���ʔ�׶���:�݃Iӽ��!i�j� �&ɡh�7�[���p�����Р���� �&#���@�;���$l�4`�mW֮���t������˫�0�s�=�c)�;ٱ� -~�@���E.����m��B@JLRE�r�!����\]u����{�a�4i�U2GUt����Y�u_���y���y1@
��V)pٖ��_�<��n���3M�����T�K�?N_`��O�u�A��Mq��t��T�����"�[y�48���z_!guŘ����޼�g�9�yA�;Ar��7Q��*vc��`�w�����W��o_ﴒK͟�I��T#>7mHi>����wW�/�m��`�)�^���$r�A&����������^t�I�0"�6�>4���F��]���%g�6B�m���i���}z�M��{�ۧ,��n	�σ����'i_6F|��m�Nq��1�Ѽ������r���������~]�����7$&��l�F�K@�(;׊������	Ş�u���Hc��l^]U:MR��y{�߷�}�T�~ �M�Ʊ�=E�`w?GLT���ܢY���������i��w;[�,�*~ǜ��\8zM����-6�A�W���}�

�ZDҺ�D��0(��=��B�1��i;�i��ò�͗yS�l�TV�<�ӯe��w�椩��r8�9W�Z��bN�&kD�7)t�Ϙ��n;���%s6��/#I��s��P�<�Tg&!��[]n��5r�4:���*uD4��}��o�t��v0�X��`ż��a�����F�bפ������� �*�k]һg��Ƨ�z9̰���7sn�'���H�̷X"�3g�`ކf*��\h\0晛\�������15̭ݺ���A����ok1[!=v���L���� �W.�ZI6O}��=G;*�����ͺ�6�LYr�4/�I�Ró&]+��i�v���B���69��Wo���c�J�&��(WW^����A�:���.Qw�m�r�2�WF`.ڪ��VW�Ȝ����*�tĲ�_����^e�e��s�H%���DFak�q�&'ì�yU���m�l�'\��������>.X�ܣK�T��햻fs�46]v��Q_r��W�D��
ĳd3�3ya��jU1��V�˝P���֫��mQ:��{
Fv���8L�ښ�TF��Ӝ��d�ei̢�E���Y�e_l=�n�.P��쎡쾫C�Xewrw�n]���fȒ�!#S��1��7��(�\��嗻�Og�G1�r�IX�:��2���w���᷏���B�|ߥj�
U����ɷQ��eXۡFt�e�{�������1Zr�﹛y��RIk8�!Y�	��b^q��,��D<���9�m�a�֒cQ�C1�1�vX�^���h��9��E�Y�v-����Ҵ�=+<����^S�ŷdVV��l��;���{h�I������y��zTx]�ז�ί)����owyY���t���v�Ͱ�{��n�VY�Ͷ۳�� ����{S�$zM���yd� [4[m,�ݝ�ն͋w�級ۉ��vck",�!/.�ف��{��y�Q�g�筶�3�ݽ��u�I�Y�L��Z9�/(�p)#����L���g����ye�c������m���G�j���y����-���ۅ��ٷ1��6M�k[-ݬ��J�s��`rm��p$ۭ���5y�l�퓖k�,��H��AkZ�Z���sM��(��5�6��߄  �.�� �E邁$~�{w�[���Յ@�/�9�:�n���[�a�P�Ry��OĈ�����*i��嬘(q��b�B��z���ϻٿM�=p�=~2 (��U �q���\�c�՟yY����X��Q�G�@��Eo�PT�
��6�2�ZiYe��+k��ڨ�V_u�����9��6cUb�W��0�΢gz=�7�P?:{{t�çF�j�S��Vs��m�='8�x�6�m{�����}�߈H<y���LV���W��5dv	���/g��u�6����$�*�z�{����"=&��_�{F���;(�Jգ��]�_A��3��~~�� �E��w�>.q�{Nx�UV��@�sp�T��"�oSc/Ww�;��̗����<��״M�Q�;��-j�cy�kw'y�Vo/JN^��=i�!$������������	���`�-��q�A�.#�T�̝�Է�h�o��� ���e����x_D@>��|;��<a�u��̇M����S�q��lm�V��kakRD��\���!5+������f�1�g��P��j�k��U�E
��Y�ɀ3ޞN�
6<6^B�9vN|�a�X�b)�=w%��ܞ��+7�7T¼7�e1��Cr�we@�~ȼυ=,U�RX�?n�'��y`�_N~����G�{Á�}3~'�O������V��V��==ϛ����\�2{f}��q��G�7��ʏ�wmWĦ�6 ���op,e��W�=��>{{u���7(����	��t� �?<�@'ޛ۠�7.�leZk�m�8A�G�~�3�<�&�7r��}�l9�M�7h8hec.���}�Y�(��2vr��̅���N��C��ʛ+��  >�F1�j
��Te��Դ՚��^z�2Z��#9M�gv:�=�T��R8�qoJ�(�瞥n:�����g�����u���퇗v�e)������f����z��c	��ݝ�{gr�&:H7)&ے���`�9��m����꺞���������@����s����g]��/�=���\d6�^¯[j�;\7g��%rge��ٶ�,����u��fXۢܝ���<�W8��6;v]�`0��8�8��Ў8�y�>�'�
�����8���o�!B���8�¼�'.���s���������=qx�_v��r��F���[��*!�)y�ɾx�?~�ۈ
�8��_��K��u=�Y�x�ܽ\D|}ܠ��XˬƳ;�k�i��{w�U;y�M�ܻ�Ay�H���M�Tt� .茼 ����<��<�W
��Fm�=�����h�W�G��Ur�d�H�劳���k��>�A ��{��f�N�^��(
�b Mq� ��}��车���7�"*���AHRڢj��cvٍu��ohʥ��\h&v(+�s������=o��&_���H��^��_$��<ө�
�f[W�?������$��zܢOw�����S ���_��A�s���R�vQ�˻��TŢΕ3@o�Y���59�$�D�]����K�����7}�୷טm=�LW_����$ ={��׹$$��������~��@��3�]y��<o�����h�:�jE��ﻜ[�A��/�@:�]𞽇g���$��$�U��d� �{�0~|ܠ��TA�ۭ�+*���jϥ��5>'gjA�H�1H��.G��ux<�@�y��{@.s[����I[�L'wۘ��O�g�̗���k,9��KzHH��\�f�G�o��o����H�ʜ5uc��4��Պ)s'X��h�펈�v��'���_��s�[n�⮩������� ��12I'�M{o�ۢQ�|�)���TqN��h����wTm�u��b���;�l�#��`���<��I5�ML:�M~>���a y�*|�A�j�yOx�j����� �=���y�4j<�I�Z�T���]��&���Xт�@�7��QN+�y0vI�O=WA�6_�N���D�~��W����R7˪��'�W3T^�si�ɇ&� @����� �}���?p�3�/{��MH�4g���}�gs��� =��愒I$�^{D�^�����c+x�s�@#��\��+�,p���n�۶�H%�q�|9a?�C�<��<3>I���BD����h�I��>������|�}�X4�OU�4
A*�/��/��n�j�s�mr��8����� Ƨ�����~�j�n�Fs�����{ә�����xܢF�wI��ó�S$Mon7�&���6ݨi�]S&#��w��4�H;&�����ĒMk��0��c���J�E��ؐ��K�q��*�X�v*a�=�z������f=��~�Փ����5<� I��s�^�	0���{ހ�u_�c��q�a�sx��{qZȔ�s�a�I�ݍ�D�����	$�>]1�
7�iBd��g�GW���v��UO1���j��`�=�7�b��jݻ[��_*up��q�yw��&��.��UQ���C��גH�?�@�v��s�?����R,]���/�@$�u楐��侒>u������D���I}1:�ws�g���m'��kŭ�kZ��.��on���/wϋ��Sa��§@W���~�Wn:�����ŀ�}��7���Hgw�|}u�s�y���
���N���{���4�܁\��&#/{s4 9S����ov�����/v�>$�O��l��K�!|ރe����Դ��M�U�2a�w���� �ٞ�b  ��2{�o�F�k}��pI$��w|�	n��	C�
 �t�6n��Z����9��T(B����ā|��UBI�� �$�^jnލ�jE۫-%��ǽ��/x�'��أ�{���i ���K0^�c�.��ܯoĞ��I	$�>]1� uG�z7�ɲ�٭Ub��3�f_��ۼ�ׂ��8"-6��m�s���g,r�o��j���œT�a�u�q׽v&iZqg���| �������������]%�a]�ou��R���ϣ����x��y�u�tuȼ�L�]�]��Ǹ�:ܴ��.���u�)C�M���'m�nd��ۑ��kA�/���v+�v���>?6Ҿ>a�u�m���ּ�s�kj��(�l]\n��L�{\����R-�^Z7
썺-p.3�:q�㰺�D��Ӯp�U�#����ն���Ô$z�凷;&�׶�[��0��֍�y\s�(�u9.�=��~��'Gh��s��>���=�sٻ��ܝ�LA�z��.,�;��߽�_�����P�ӱ��f-���Rݜr�{�q;M���Ǩ�S�٤�	 �\{�b(%W�'�P�y�s׼ߐ�Ӝ\#rGG��;ܹ�"W�x��F�I �u���ロ�m�� �sw0ϝ��桉�i�:	�fU�g��"�i��!���/5�H
{ؚ ��}0 =�;��.�n���~@h�9s�g��$V�O�H;�<��@�}��}<�9=�w��gA��g��< ��e���7���/>����l�/�ld�HꊕF�[�	�6�M��9ròM(Č�"�M��߳�C�1��4�1���~�6�{��������	��q�{�Aĸw{ش�I���PG_�v�*�܋0Ͼ�w�l4�щS5���!K�y�|��������ΣKq�f�d(��^(ę	NW#��rb1�2>��eԤ>��7��u�Gh���Y�1�T-�_������_�b~��rb 5��w��� 9ӽ^��A˳��Πwg�-BwN���	r� ~'˻\��D���k�/}��]���;�K�/�,��/c�w�Iy�A��R�j��KkT�oD|�؉��?�D��,�ݲBI'����lL�����}��_�'٧��'uj�p�{��	��?��'��0�SI5H�y��Q��ID�$j��蛿 YU7�o�[���_G.�1+�`��z�v졧g��]`��R�K%"��wݞ�ܝ�N��w�5D�c�k��$�:�1��^�GtWuK*�ܢI�l���8��6<�����>�.`����o�S��Q ����o{@ �}鍒�D�>�E������=9��p@BR�D��+=5�D����4�I&�c7n?f���oy^xp��^�zof�����K\�>���.Q-Z3F�R�W�c�YƖ��)�'~���$I����l��~�����\�=������T��fh;�{�9�>�؀A～��������ݜ�~b��ŇXD��RI(�i&�^��WYu�,�g{^0 oz���܆����'��	4I+}�� �N�[�˗�=g\�o1��a %'�"�tr(=�u�1v����jLw&�嵍6:�'Z�������ؑb���~��9/�Id�ߒ%|�~�����Z��+J�|�]~��$$E{�s4~�t7&G���<�g};����`4��ߡ4H�ݩ��'�F�Q�D���W��H�מ��O����`�9��~� �{˘���c�X~��\D��8�I�7}��ğ�����.&�YmM;b=w�ns7�yf�oq ��]�ɆH���&ݟ��0���7NgYd`GB�e`������Uf�n�x����W2!t�����75Q�!�:T׌�{H�.,���;L�*^'�G;��c�_}_W�|�o���G�u��n��Eu3ｻ��I$��9�Gw���ȟ�̞�'��v�^�t�����$M�|�ת��=�Gt������vQ�n˷m���zy�^���y�-c��I��{�����Eb�ó�=�.`6 �v{� ��}��{o���q���>��@�9���P5�Qv6���J7b��-���y/o��/7���/�Jo�j'R��M�	 ��7�Ժ���9��hNL�7]�ߞi�����{�Ms�I$�yl�>ʞ�W�8BI$�+ډВ����	c	eUڴ�G]QǾ���ɮ� Q3�GO	&����}��D���{B�e�^�m�$�mw3|��lղ�ӵf���K`|��;�	y���K8�K�t�ԉ_99�rI$�;�	W�J����^[�������=�u&$�C��9�>�5fPِd$:�v%�0�-t���j55�e�O��_k~2�s39�V��2nk������8��4�	wǹ�˸�����|Å�{\nn�l���˫�3pV���i'�Oj�eB�v[Z���hHn�E�p_UVM5U�i,����Z�u{ò�����U�g\ˆ���&�������ۡp�}���e y
h��ә&��'��a`S����vX}3N�Ψ�yy˓����5���9t<Ye�4)T�#�#2Lk��$��i�*"�i�i����=�r�S]R�z.2�X'�u�}֓ӣ�+�ʈ.�T���+6�݅�����Y"��f��u\�ׂlmX�L'�@���ܙ[Fwc�b3��Z\5�)4�Y���fj�(ؓ����Uc'd�+/9��/n���Vv=�.��
��j��X��}õ�\)*8�\Y+6��B0�]�ֽ�,jM�Lo1W�������`֬�z*�Yx˲����u-s�˙Eޕ�7����l���	�5���+�mr��i�X��f���eLU
��*���;.ob�֖s����
K�+��]����[��fS�����of�.�x	��q���2�V�'r�˳-��^�V:�N�1]3I?'v�����pM�8:�ICwG�Z@U��{�3����k4H2P�قƺ�39ݎ���v����ʕX�P{���r���	�(��W��ɱ}ȊH�O���\8�BhF�5�� �mm����e,��H���[��z��Gc��Xyy��G;�6me�ۛ�-�{g���0�i͛H�V�.R-���[b�R���j!ٽ�^f�-kck,���cQe����6V�Ѥ�&�z����6�n�f'�h�llN�lryy��#�mq�{�Ŗgm���������-��m���Z�,-�{{�8m3�kjɰ���R6m{�򃀤��9�I�mk$��N�c2D�̭l/m�6�r�{ޒ�4֎i��Öm���ڶʹ�o7��n��v̀&�]�mݎ��'I�n{��/I;�w%Ȕ�v�3k[�	m���Ύ��rf�m��L�yY�YgC���-��!�ݷZ~/�~g���o�����Jva�x=���\<����nd�Qv��m#/mzO����5Ŗ�9e����u�p�/W��Z�8V�ŝ�f7n���,�����Y�W�Xk"�nS�]�:�v��g��
ܹ�<Inp<��ݻ�6Z6����n\ŝj���9H����s�벗Bk���ЏM�v@�0��A;w��?4˯so&t�k9���5��ۍ�p=X@9���9ػjϞ�{탗Ş^xƸ麁n�vɷ<ɭ1:<�v�ƶ����ce�V�it�u�������f�q���X�+�D��=�p�܊68:SO�4vݸ�Fuٌ��m�n���K�>���ۦz��JG]n7ܸ�ӝ�\n�c�{G;�#ST�	:H�,�B�X`�YG���B�=�N7!mzi�<�����v��)�B�63t�ޚIC����;;4k9���s�����ْ9��#�3f�����
�t3s�Mֺ�KUiܣŝ�=��u"M;\e�x�CMu�ۇ��2A��t�6n�-<|��g�s��n���Ji;�#-��vJ�m�]�չ:u�uc�w	Nۥ�솏b$2�Ls��''d�Cֶtp�i�F�֠�#T�n����D�7@��ۗq�o9nȳ��:��-�����>x����22�IU
"����1��7C��\��ksl��uú�����kw4�o��;z]iْq��'x�ϱc��޺����q�uU�y���ވXwn��SY8Dn���'�p<��]ݠ[n"��X:��{b��#�Ӯ&�q�xw7%Z�R:��OC<ki�Wu�d۞�z�|�Q
P��l�*M�N����]V�9U5�q+ &�b��uy�O,w,퉻2��võohcs���������c���=vK��1�s��tYy[�Js]��q���-��M�P�(� Um�'�:�H&+U6���-���]hP�CJ�
��鹕��k����wV|�l���^�Q֮��{���������8�Z���Wj���H�{mV�dqc�p�t��8�|밇�/�ї)u��'c�s��o\I ��]p��p���ڶy�dzx�1����䓕�wk�1��D��`�պ�6�7m�vXq�C��p�;m G��'N�b�A]'%���ۧ����gv�5�5ϻ�k9�ʂ=vN�p�c�wt��.�$��n#5�u�����U��g�������Ton�I�$�~�~���������Gb� ���К$�%��0�.,8J�G�7_"	'}�d���m�Ëv1��3G=̹��Ǵ��>~�'�5sۈ$�I99�p	 �l��A�}Y��$�u$��E���hÀX����}$ %���M@V�)Em���H�y�d�I4_zcd�B��Vm����2d=���ی�
���hD���B~$�i�D�$�R�׵�w���K�<x$��ӻ�L��J�H]Я}/I'BSd�0^l{�#˧W��I�ޞ�J$�I�/ޘ� 2���Ŝ΅�Ҫo�u`�gԸN�Ph;Y�97cE�<�6�-���ӝ�G9=i���}wv�&�?�<�� �-�v� T�b� �~Թ{��p|b)�w{� g�˘=�E���Q��J�u�Ԓ��|���ʻ�I�=�sz��v5q�;�����ٮ����t��AóV���g�Pm��s.�E�m���������>���{}�$�Kg�u$�X�K�N����^�｜�>Q�������݌n�c�LG=̹��A�=�q��[��yBd��<���H.�ޒt$�O}/t%��u��%�yz����R�hm��F�@'���ؙ$�D����J�g�wvI��sll��$����%�?V�d��n���}q`��w{�ςycE7�b�kIoo�I:K���{�"�[�N��S_t�8b�z��.;"��g��sĎj����A�^Sq�f��m���둩��o�eP+���x�Hӱ� ^�I'đ]]a�?go$�h��.b ��~��$.sˍ1WmCjU��﹜[ �[�mN�X��D�k�<�d�$���I>�O��z��[����9�ۻ� �9$��N+����f�k{��o`�A��k���b�y�1��77vs�4�7\�n��f��^����;r|��ޅq�rv��m�q��k�T6�X�S3��v�()���� �o4�	/�/���� ����{�="qn�6Wc�LG#��[�K�Y.�L_��T�^�I$I�{�$��B�L^���fO0< z�k��&�}E���@�����%B�Wzb�wm��W&2�M0��F��I+}1������A�`����m]��>n�͸�vCf�%�v��@��=��竆m��z�h��V�!~~oݹ��=�ϡ5D�%o� �����3�;/�e&o�x�����q(��bڱb�7G�$
������Ύv!�$�����H��^jD�Ula�"���l�<�Yv"�n��l��r%%�LL�I'� j�'fON�6�$���������\Āѿr.H�r��1���<���z��_��]�ʨI&�@[ٚIВ
z;�v}]��K���t�eFE�R�e�B���R�[��n�ٽ��:"ߓ�J�x*�o��ْA��C�έ6�f(h+�$�]<�s�I����	?����'��;T*�*��G�]߸�A���Ň�����Ǉ�0.�~����H�}�� ���ߒ�����(�%Q)��:���^�;A����^�[g��e�苴9n��|�}8�RB�9]��#��w���H �~��?j�5��L����,Q��{d� �뙠+dj�i�g�/	$_O�-���	$�o���I|�w�+���}�*[}�~�$.���X:ب���=s4A�w�0 �-4}C|�����R{�_��w�1[���U��q��#~�w�C7�Ēq��d��$����jD�~��t�H3ܘ�M�	 �y˙���rJFتr��bf��3D�%�����y Z��<N�=���H���ؠ����w���+�����{�3f]Ȗ0���� �E�z/Mg�ܵoڒ�y���x��ɪ}y�ѐ�e]���x��QT2��{�������|S[�\�&�y�͆:]�B�x�st�:�����.[n�u����� � #i4�1�'n㌦�vsku�Gi�f�Ny����}�2<����C8�\<W���G$�J���sN�8����^9:�.���'�]��c^�x�$�E���$�ݶ9b��6�t� �/kpYnɤ�����`���c��	�vRX��>3�:���ӗ�˱�1�ۛ2.ބ�F'$v�e�Ee���Б~.�[n�Q����I'{�d�O�}��7�;��u�{]=�� f��C��g�#�HRG+�p�}��k`�Ӿy_L�,ʩלA"Sr�V��_k��w �Ht���1x߲�ܒ�Y�Z ��u�H\x�N�� �{����U�ݗ|� ߉4H~����$����q|�U�Q�?�;>���Q>�@�^�v�J���$�{�lP�S'�����@F{��<з��m���U��^�'ВM�v'�>n[]{xw�t�$��Y̺�I*wk`BIO}����qƓ��F�%�;@b
��s�qvǧ�����Kf��Ev�rp��
��?��۞7\9@_~%�\n�&�[��!4I$���0蔮Q�s�s�mZ<g�zݐI?/{�H�һ���h��LH��.f��2���J�{�뗦��
~��9� ��d	mu�К�~��]#�f=�#En���6r��	���]��OV�@����o��BK�3�xIHQoctH4N�~��k	���R�/X;lr�����`��fw�����y���*~��y$��l�w ��s�0	���ۛi�B�o�{�h��v�S�{=�Q$���ʄIk�0 ����O]�M9�_������Ck�l�i�������  �3�5��5��~/<���s}��H$�g��D�D�����5��)-�X*�6�Ӭ�Vl��
q�m'a����7@n8z졒�-hs�伭���W=����{�I�݉�~$�'���<�����՚����o�z� ����&*����O���6Q��y�v��Zq��I$�[ɆI$r��?��O�j�9���M��@)��Yb��L9{ˍ�I�{ׇR_%��L�q=ž�-�{�����|�jh��u�l�t�+��yH{n�	ژ�v�0���s�`��xWs��.*�y��.�Dmt�V��w�����_ﾪ�����$�h���!��?g�`���p�N�\���e�}-y�C��$���D?�$��ɀ�I�{���R����k~I-�n�I|�S⭷6�'l�ǈ3��Ł���7�}	kv��) �{� {�1�Cs���f"Hj_z<��ن�|ն�֪Z����6]�R؎���!�WmBj|�b�0�����u��Ex���7�wx�D�O)�H��?Tܝ��^�ݖ ���w0-��u[kU85Vb=�ݒ�4M�����V͞�yma$��;���I�O)�H%#u��Bw��i��b���U(��A��w� ����{4����}���$ 绻��w�����	U����6+c�r��z�moE7h�wh�D�'�� �yM��h ��s��"�x����.��<�P��תR���n�W��N�e�s�j2(f8�/�����X]�Ȳ)�-g]�	�[|fR�����p��U_kWo�h��ܹ�k}�1�%��~��߿l���%�]i�ʹ;B�g0v�_6J�iВ%��?wI�O���HI��>_#i�֢�EY*���:877�Gi������g��ZHo;c	~���~�~s��I~~隣d=��{ vs�0$zy^�G������C���^�����O�O�֮�(�zoي�
�����{f��V��&�ޛ��@?��֊H���1J�}�k[�S�H�`:�U���_u#���{[����PI|�Y����zNL$�~nn�H����+<y��E�VQ�-��	�S�/(�eL�h����BI$�/�v�$�I��z����j^v���+f��"����r��+c�����6kA��mӼ�&;+�^[���?W��I4d>�� v��vk=���R�k�7�59����TL�s����uf$Jz&��m�[b�07�>�8�1�R��u4�ti���d����|'�(~@�\]���-��6DЛg��F�9�z�A۔�r�k��]��d�E�&v�a��z<�{vz\�:'��c��z�;f�ӷk��G�o�7����{�8z�-�u��v{$@�x�f�kv� �mz櫝��VJ���ȄFB��Q3M��v�n�v���(�lX��t��p�f;<�<����s�5Z�U'L��n��ed�}�2�rt�۹K���v������q���F��-���r"�~o�� ����U�_�����=��u��~'��*ݩe�ꁬ���I!'�M���j�� ir��"�D���d�Y�_H� �yZ�-��[ ��}� #���d�|��%];�{=��^Q���r�WUx�L��J�A��o4�6 ����E��;��6#xw��� ��zo1@�g�T�F�_W�7B��{��;r����I�v�$��de�I5ӽ�5�7��=k}O�S���_t��$VQ�-�'����$��l;���:�\��I�;���@�{��HR���'~�>J�H�	�/��Q]:�m�N!r.�&q�y��r8�H�,qXhhv�qx}�lm��vz�$����_$��=7I�	���������A��}�\o�'��5�_̣yyG1����` +9�0&�]�sRU��o��&�?�qE0�Y���hG��p��0��me�Ӵ*'/c"���K�S7�i��m��=�k<`d~ɛK�"�UW�Oy����$���# :$���$�I*s�`M��eS�`�~����q�*��#��U.<A��LZ&w�7O�Y�s�,k�<���׵D�%vh�I	�Ӹ���Eb]���e!���_����N�]o��#�cd� O{��I$�Ϲ��b���{y�`?��_�@h^�zNʇX�j�e/OIP��$�w��l�-#�*�?g���TI��{�ID�J������u�r}�Zq�Q�Z������5�h���
�z�8%�-t�f�nI����~oõ$V:���s{��� �=��[ �P���ms���{{ŧr���ZH4I�>�x`�C�H ��Kk@N�M��I߭���?=�K�2I?iｲO� .�bT`h�Y6��Й��� Ո�/��U�^Q�v��wI! �����I�o�N�����f���[ɪeX$�4+������]��ծ,��WY9LqfG6�,��L{�wK��n���:�dtq����@���>���������2��HPٟ���E�l�8-�ėh��M���^&����o�)m�]*�kyi����ˮ��Ur��ԝ�-�Æ��?�3��杲����>�g/�
0*�]��K�hP?b6h�Hd5�o�KE���}�DŻ��^d)`p3{Qǒ5[Yq?��QX�/�«�
^;�=vƕ�c(Iq�y�|�dܖ�_��2v����18)}�{F�E���RD�v��l��J��lү]I���s��l���1�T�ǖ�;k��k�����Q���QI,��vBsr�F槖�m�*���~�b�-�֥��:�g��Mu��`�R��Z-A���X����Ñ�ʱ���{rl]IfYt$�6��Ү��E��N��2{,zx�]�ܑU�%�����mt�.C�Z@F���&_e̬��|��Rηg�q�u��_Lu�ҝ�*�]�ե���U}�85vY�nc�,��j��.W�b���]H����T�t��Qf#��M���@Ɋ���Z�8!PΚ�Y�^k��[�0Ntw�X�x6�7�4�](7�"��y!�%�x9�{�5��pK2^���F����re1��Xݩ�U]�̢����rc�o%��>�;3[pf*���Or�+���m�k�Ή;}�έ�L�p�BEY��Pv��5Z�n��j��d�cd�'4�槵dH�'Z{[���;ڷQ-������-��ei�d�;^Y�[�KlQu��"���m��3L��gZ��lqֹ�tIGFE��'m��C�:δ'�6�Y5��
L�ˉ:A;-J!��pmj�,�:�QD'�[��$��P�{�Q�nBsn���&��*�J��rڳ��:-,gu���g��3HCo,����Eܞ��Ύ��´��9(��mT�ذ���kH^ٍ�n����fts�m�V�앭ͮI$�K�;;,���Zt�W�;:�-�L�rv֍i�)n�D��9��m��螽�[-�X\Eek7M�����RPmj
r��4�j1y$�~��m�H_9߳�I7S�s����ԵKQq�����g�G�<�������{y�����rbB_)鷮��^]St���������G��WQy��=̏=����Oa��%��)���$�I+���h��O�nf���\�=��n�m�AƁ�}������mlۮ�s��^��!�Ě���M�Y�[��|�~�Hz��Q�W�s��� ��ب ?~��L2k�Y��g�+��G�J$�.��}����h�Ec��34���&����))����M�ЀI�}��I�	�m�'R{���d��(�/�}�G��%"ч�9Os1P@��:$�>�xTˬ�|��I$��wٔb �=����>�h��l�K�����c��Ԫ�)I����	��I��tI$���t�������r\����˸0�6�,7��x�Z��f�u���9G#RUA�8�u�z��0���r�&��盯���ߕ��By�Eڶ�kU{�op w��!�'}��4J��X 3���$����'7�����L��y���("i��sx��٣i��琐cn���m�Pll�s��I�.m����[5t"�/w=� {��u$�Iz?N�J��n׾�՗�]�)L~��	$=��JX��l�՛��i'�j�)���) �IG��$�K��wpI���6����7*� �����mY �� L���ŀ�A�s��m��!�o��rOo�< �������绽�����@�ں-d|�����=9��P	6��jA$Q�;�$����Y�~��I�ws|�q:���KP_�绽�l~�؃���=�e=g�L�$�6� Uӻd�h��}�1��C��c��*�.�������똓���t��+xnP{j�RYY#�g:zKt�X&2���n�WKFkE��M��ڭ7_Y���z�!�'v�ۛ۞� {i;fp\e�-�]��6c��ڸ��3��,�Y�J��8d�n�c�mD4
F�ꄶ��PV(���v�� ����\᳹t/G�j�y���o�j�#Vz���yx^�vᴵ��7k�]�KUs���^#��Nv�p�;g<t��6�������\8ۭǂ�4�V���a�L�&�P��@Z:����]{�Ya�wm��,Oc�6��n�u'n�\Ö��/7��rjԮ"V�L��#��P�7`����z��@ ���f�� �{�x�a�ǣ��|��PK�y��H:"!�uR����w�\���߮w����}=��I$�s�I(��!-� &�Z��k2k�,���� �}�EK_$E@�^����v I��U��Ǿ��n�A>$�i��$�Q&�%-�0=��V�+(��\�����nK�Ή愐	m����%��ӡ$3�/1V]^=JԱ���F��H���@���&#�ܹ� �z�s>�B��
�M��I(�HK����4wϱ��^_L�߭�9yߚ��D?(ۑ�%h��F^�A	Tۨ��2�D*�EB��m�b~�~RX]��O#�緽�����ؠ 	�>L2gX�Ϻ������HH�w�<�}E�5e�rFLx�v��yrI��������������)��_�j��굺кST��-���q�\�!!��U�C�ok��ߺ�����٬�ʹ���@��y�����$U�߮ZI$���w�	�0�u<qȐ��,�;� ��dwB �Ϸ=� ���.` ]�K]}���}�� #�d�b�4�{�3@��`v���h1���I��ԛ�!$��ߓ��($���i߂I%��ޝނ��^jG���ؠ��t䮸*T��w7��4O����>��:eo��!=��,�D�3��n��������+�����[���'�y8۫^TO\�=��;]�{=�@��u�d-��ɝj]4Ge�m��@�% ����9��$A'<�u$�I{�ӻ�EyϷre�J�޷d$��zcժ�UwYy�ˢqۣ龒Bj��P�����\D ��$s�N�J����A-�o�K�/�r{ؔ&�Q7
)]n�����{��I$���$�Mצ:B�ƭc�ܘ�ރy�k����.����[ӭ�YV���n�Y���آ^�^Ӫ{��_�tr_V8D�Kj�tލ�or}�|>O���"R�?u��+������$��:/��q�t"�1{�ά����Nh�e$�J��xIԓ�>�y$���ӱ�����#3ݹ�z�<�+AQ�9�T  �v'D�h��T�|((�~S��d�L��Q'�Ik}�9�c�>X�'��G)�5�ں�ۋ�]��~!�v�kn����vG����zpT�$'$����A�s��m���ɇTN�^Y�[�V٣x�6H4_?H���'�)-@��U��SNc�߉?أ����q�䟞!�D�g{��%�b :�|��(;[x��m'�O�Gmiؙp�=��{��@��_�ԗ�/x�O�磌�a&��>�I|���s�}E�`��+#&<�g�ق�g�����w��I+�G! :y0�D����̯w�N��Ve�Cy�0n�U�0��&0扽����3x��3��3���.
��i��k�+�a�=�8jWtd��-���}����7�T����3�0�x��+Nqksjqݥz�^�I$��;�.���=A{�$�t��?h͞� 7ݸ�W��)������JV"Q�H�W+a��n�GY�8�o>1�sl�v�*�7	U��;�z����
��x���!?j�����I ���0����i�Cȧ�}'w$Jt�{���2��VՕ	�$�e��]�f����[�no1�ߖ��}�	 s���т�}:�f־��[����"�Ue"��iQ$�'u�D�I+��t��#w���0%'��:$ N���``"���+�sޛ��zo����7� H�M���~$�I��&I=�v��7�����w|�� �w,U�d*��K}�6�I%����,F�3;]'�$���ԒI7+�i�ޏ����]��k�z�k���;Q��Q3]�X���]3��D�2)zgU��<����Q��JDѕ8z��z�쓸YMn�Sz��M��"�k���?��|ϑ�x��vl]v�sغ��R84��������\�k�8�u��:�r.��y�^]�v���ۘ�\@ipx��4\oM�y�9v�8��ȻS���{uYɭ��=h��7(�ޥ���YMV6���W&����6��=��������;�na��8�C��K�g�@���t�{����N�=�t�m�j�{k�۱�Δ��J3�͜\s�- r�u�Ǚ��p]J��z�;;�#�������_�~���K�y�=��s @I���]���d�D߇�r�ݫ�/;gi������h�}7��#������ݚ�t[��'I�'�F;O�׽�C��[�� ��� �{c}�&��ZW���N��4�>|�&⭉ڜ!3�oh��v�� &ɬ����l�<ĒMǣa o�����T�W���RB�Ud����w�H����H��|��OĚ��쐒HS}���������?�;����
b|���%�9.^���BI4J��@n��U��ğ�����v쒉$�*o��'ia�J��������A��3�y��(�>�7la�4s��Z�T�c�=�\qW�����>�xI����$�&��&
�a{ۃ��mn,���&?7��$�bI?�e�(��S��&�U�S\1��<�rywwh�ձ�`x �W��k�k�z{���m�gD��F���s�r�*n�����x�kT�r���W�(���X�'���ܢI'��� d̤S������/�_�Ao���(�\C�����%��N��D���q�'�K���H{�d|Ho}��I��=F�� ���*�Kfm�>�9>���F%����!$�[��.�?j���4�K����
I{�����c�УF�Ud��S���$�K�}z5M���mf%�ӛ��$7���� ?Q�������-����@i�r�S*�Y���۵��$��sm���R�Q��V�����h��2�x�>�I	�M�_���I$���L?�.n���:���z��v�H-�Sv�	�jV�ɏ{|�İ;�xܓ�7��\�I�$�]�� 3�}��0_x�������5�n4�bh�L����I&���tI�o]��`�'������Vwb�lġS T�l4�X��l�悤����j3X�YÛWe���	�}*L����r��."���	��<߁�����4?s;s G����tغ�tX���5�fTI���b�$]�2��$Rw����}��4�Ú;�"�Iޝ��JH�h�3(�l�	D�}�9�i�4��LM� ���˘H�f���\=�q^��~~����6|�}�מ�;E�-O;�;:�N��������j�ݮ.���H]I[g���� =�r�� ���~�����t���Z|��v6H?Q&��n7�%��$w�E�����.��'�^�C��<���}ؙ&�?k}�L2I&��=$�H��������=��w@)��o�P�vFLx߽q`��oُ` ��������u$K���{��>������]��#n;Eb3�z��|S�7��f-� �s�>$�ܞ�~�v�
�=ٙ	�٣/$�sU���-	��F�ͤ�6m�y��Z�
�+'e7�nj���ʨ�iM�Q��ܗ��&]S��o��כ�$�u���=��
h-7�k�H�q�o�VH0�W�n/$���:�	!����A;���e.w��N1*��z�U��8ٝ�v���0��@�<�m�������~����?��p�M��<�9�q` �����ؐ	ߞiԧzo�&iP���B|����I!����� ����.���&#��\�$�S�;ړ��5$�H=�;�$�I|w��5����x:E�^լ�`G���Q�=ϻ��l �v��� I�U^'{1�F����$�c~���	���f��}Y'յk��1�{~��I��S��{��`h߽�<� 엮���P5�X	/���w$�5�%�It�Gvz�).�^��G�{��y���=nh���]� �4}���*�T�!U�ڷ�� ��p�m��]��1�Ys��Fe�;%��KP��l��s:J���V��т��^ɠ�gQ��@a����c��LF_׎e=��ґd���f�V�K�x퓻s�̲�*���sj�v����s�)>��^fZ�1��Ⱥ����H�ڧ��L�(Ğ�v#7��tu,�몙*��2�D���
���@��,��.;���5(R˕+FSt+�r�M��pSwkr�n�?�}����xeF���u�}������;b
�j��4��#���`�ިŝ+rT�ޙV잒+d�|P��}oe	,'�̕۷y�Ù��r�D[V)�9ga�\�7u���p�y6I���w�uh�y�iJ�����\�o9)#�o2��6�bg(n�R^#u���9â���Y�����'9xk7dJ�R�	dmX���zw���$*Mg��m�n�/��bc�)]�]Z��//x��-QAJ_ea$�;�:��ʑ#���B����	�:Ԝ����e1����(��d'wn�����~�2���rjȔ���H�[I���gm)���|�����I|O�.����"}��
�Y~�=���L�h�\�gh�V�����6��^Yy7'f���:'$ᖃ���dr�k�#���Y�xi�wRڮI������y%X�+�+���^I��+��[�^7}�X��Yْo�g`�X�:V�4����uj��e��ŝx�P�]Y��VT�b�����P�6�����m�QtjQՇR�����ɮ��3��}�~����d�D��的ㄵ�ft���sʲ�mdt{a,�O:���,m	I/;M�{T�Y�k��vt��.�+�'�tQ��^w���tmo{Y�r��c;��W��/w�Sm���^gHQ���+H�{D��g���ru�[l�ݽ�6���u�y�^�.8���'#�����(�����̡�7���N���Km�ֲz��=��yŤ��=�����3����ҥ�� �g�Vi�c���ge%YnBFa�ٷg�ݒ+N	i����89m؅\�;jʒ;ʰI/1�X�v�����ۂ��""r���m�̰%����t]�6����vQD2$%��� ���"$<��ne���D��c9FYH�:���Z$��۬�2���?�_��om��.���h8���N���z��yŻX6n�9�c�v�])��nttGfz�n�ˇ6�sjݤ����1m�6�����7`2�c�;����x�Kث��� 5/V�ܘ9C�G�4��<��)g+���5��ŏ����n�J�� �4c�qҐ4`�]����0�m�^ �j�ݯl��:��m��D�wPN<��V��]�vLF�q�y��$���]A{=n_\q�ܱ�e �0��0�Nx�6^���ܝ�� #�>c�|g���x��i�E��z�l;@�������d�]���l�y��s��Qv�֘�9��צ.I7=:�ڶ�6�����7��84�7l�Ir�=;شk=:�������{N��N��'ѕ��<��M�UQ��|��x��/�a�-j�q��p40r6�Z'	KdB%h(�^r��ۇ�;��pS���ݒT^&��Z;v��'u��67�=��ڬm�-�;��xN�6̎}=�>)���j����no��/�S��<[�F��냑۱��E�m͍v�=��2ۭI�Z�2A�=�n�QtNXv��5������\{j���8�����ll[9���ٗu{l�ۓJ�h���F��-m�ݘ�m���c��*m��y`��󣋬9.�c���[��xɻ`Z��f9�{��v-����F�k�AZ�8\���s�*(�٧A'DD�ZeA�B+("�1�y<G[iW��mt潞���n̓��p]zx"&�)����{X��귆��:�c���p���A0�@��͛{'��������]n��U˹�&�N��뮐0TF71���Ǉx���/n�#-Ʉ1�0���V8h�����&���^ܸ�@���t��ǲ�=�R���(�t9�;q88n���8��2ώ��:۷11��fw8��v��[@b�-y����'y-�R�x��^�{^5��\;��ܕ������
����+�;����u�C��&�W����O�u��\��v�n��s��h-��g\snM��{m.�`9��<�Q�h6ڞm�j	��F�{&r���v1m��n��7��`�ƕ�e�j�������Ʉh�%pS/a�;/�/�y��-P<�-�WA�v(]���ܶ��cp���ݵ�z����J=T�Y�.�ezb4��%e��\1t=��!1��1��o�j3�˸�w`ַܔ�C�U;Z�"m{yzy��u��ݸ��OZ����{�q�6�O�D��w1d�7ڮn�D�I/�$�:�R�Coz��S�7_w�	ϻs+��WE������dd�6k�-zw��s|�Bh�I�>L2Oğ����w�I�izx�3ބʕ9U5��`��o�r� 4�����iG��A^�6ޒ �}� �$o�o٠5�y�RҨ��=�gw���b��M=݈I$�=�L2MQ>�<��gKc�sa'5�璯5]�!X�n�6���~��/�M|NΞl	�S&�F6�K#�iԉ/Ҟ"t$�ӽ�K�/����<���>�&������:y�kf�H]��[Y�ӌn�S��Gc�r5!z����mKR��.w�0s���6ٯo���Mo¹�܂to�������FzSݤ��,$P�Bͅ��7Ӵ�H�N�R�q^-�_�!DL���эόAm���w��{���|T�Z��Z���z��&뽆�a{��y��L��>[��Mh���f��$�ӽ�B@1pɪl�W��Ai(�H���"�V�'��t��h�Ov��r���a��qs.1�D�F��S�� ����!&�M�|��R�&$s�r�Xՙ���ޙ�!�߽����ϫ��<��}�q���ffC�����Y��>�t��I'9�&�[���������z�,�k��%h�������|�{Ʊ��y �*AJ��1M�%فv������-T�S ��R;SP�����蜍�O�����,�9��3k`��a�+�W0�f�T�����R�� �g���i��W�!�+jQ�=˻�I|�a���7=�ݦ�D������H+~��	�Ji�����U�����<i�6�VE����N� I';�'�~$��c�l泌���IW/+,Tb��V���Yޫl��g6�|9d�x��WC7��d\VUйB=�1ܒ�8��[|��vs��}Uݜ��~�߹�� H�����4c[߫�拀U�[tK���'�4����rM�I!~��t$I��x��GǶV�4�������,��ʊ�.�TfL9�f7D�@�kyY���5���+=9�JI|���R($����<%o%fﲹ�|�;������䤴+�h�qpj;\����;e���:�2���|�`�*���wI>	\�В"W�Q�j^S�5�TQ/7�~$��n7D����0D��UiԽ��+BB�]<ߗ)E��9��������=���h+"7���]��}��\_aSP��G�$\��b��H7�ŕ�AW��>�}w�o� {�� ���b����;�a}b��u^o��Y�10Ǟ�´�@�WȆHv�;d�$�o������g[�v^�yi�2U����f�X��Ȩ7�8��+�67f�V��.�
���sn���K]
���#mW	�^,��v��$���ݓ�A��`��`.��%���$�+��ʄp���<�X����.f^� 9���(3@}�����o*�ܤD�����H���Ο;k��(��;gћ.&9=��ۑn��L����򦫗N*3��{ə�@߻��K O��6g�i늄1;��� �I��{s�<��^}�+J�����gu�A,[������s>���4�����y���H�s��J��~k-t�k8u�n�&�A1�gy=� �}���! 佫7#���n�&4V{�ȟ��=��� ����o@qu���QM9F�`
����ͣ��]�/&$��I;��vh�6o�r�4H��׹�:{;���7i ���j�� Ցan�����~'�LL��}�2mv��'ʲ�[�J���$SӤ��D���$1W�=�91��������6;�Y�3~��a���m&�Q"��bq3V�W_;�opuͭ�uos�刉x�F:ô;-�����~��f�ͮy�ل��]����|��;@�[�����66�����M�t��>v󶮺h�on��Xոs�z�ɺ5���Glt�ܼQ�8%�9�+���F9�O������S��:Z�O!V9yt��yG�=m4ssy�x0��7�5��Np��i���m�8x�`�����냷C�l�܆۴�����g�=U��������3:q�u�A=t����xj��<av�Qv_�α|ܶ󎲜j) �mۛk���\�kru��o����:9P�$���d��{�.Ϗ=�dI�_�$�eF<��J�T-�d�%���=�՗8�*Jvh�TI羒J$�#[� 'XR�ޮw���i�����_.�BV2:�����gv  �g�؀@h3��7��2��m@�	/�g���K����*� `b��@=�!��ҸK��"�o�gsk`{3�c��'p��Ꙧ�w��'�Ɔ�PB�4��r+��H%Ӫb�A�M�W���$��N�Q ��6H4I���ٺ����-��2"�(�"#)!�#*j��AA4�a$(W�1�EPGk,��gyҲz��YG|qzzHI$��|��I$�ӓ 4Y��?ԫ^��>$�I��ߛ���k7�깢����g��İ���9w��l�v��k+$7��P�=���Ue!���N�{�r�M�j��N��T��h�NO�X�0U�PKl�$���Z+���Ky�fӗWs3do�B�W;�Y'�I��c 2T��S���\-4��4�S�?]���a��e�F���\���|�~/s} }��P`��ۍ����e	Z��z3��y'�:����H���$�kzr`I^^�����2���N3uA.|���6������A��{5��w��i�i,�o|-�����$�h�K��� +�}$'6ϳ�{���O���l�8�g�݄�8w7���՗%�f�$�mru�n���[����?F7V��.���I?=/��I��T���J'�ˊ9|�`X|��Q$Η��=8�Y���5�i�qI���2���6M��� ��s,�J��7>$�Ddr��3/���T>5��W4J���f�;��d,�ٺI�	��/�WC~QJ�1nV���yJ�]�v�L���=����I^{��T~�1X=�@�l��׎�4���B��L�\@�L�=��3@/��o{�Y��|�ԅ���8�w�d���W���J��tm$�K��nUI���Tf�<�1ФA�B��N��h�G.�g��ʻe���$ ���g�|	�W���{����Y$�K����MNo�7VMp�I^�"b��߽�)C��ʌ
If��X���6��u;���;k�*����������ڪ(����g� �>�}�޶��]�9ov9Bn��R�ϋ��n�$������@N)
�V��Ә<�y-�|>�������3V<�PI���	 �WһQ:M�;ڗ�����vEwT�'/,}����3��d��I���D�6g���)/f���h��� �V��uVQ�O��� n͠�9�=�Y�Ē�o6'ĒM/vF@tI���u`�ؕlЫЮ%N�\�.<_SzI�s&�*z�Ps�G9��=�S�'Y��>8���K�[:5���Ռ߮���4���7���i��ɩ�*3&�&f(��=�y�xG$����u���'��zw$J�ݤW� ���vӧ��Q����s���q���eݢu؜m��S�`�z渹{V�;�'^xz���|����Ҍv�sh���I*H�q�I��s��>�J�{�cc�'w�H�]�)<��ҢuEV�Ϳa��(���.�.����[ o�vo�@��fQ��&�9"
����5�b ЪVRNC���b���3(A�W�}�{�N��$�H,~���"�_/E��BM���fʴ�^�7۲��'����D���� =}����[�/�,W��m0��w�\o���ޫ�R�$&b����<���o�s�ɻ_a#6�t�RJ�y�R%�G�h������H�����c�����iA���O(�خs�PN�<�v�ۂ���Y��²k#u����G9�W:fem���F��2��G�.�Ĝ9[�ZPz�	;�.�'Kiepi6:�$u�-�v�u�;�m�yu��Noc��v-�N��NGS��]=��rW����GF�x8��m����9����tzt�'��I\��nx�u�ڼ�=�ix�#Hvx{�jݜ�� �(>K�>e�\�3�n�fE�D��^� �K��y7]7C�Ϥ*ݻ�úm�@���v��n7g��q:�:�(AvL�lL�81�&5]C�����~���!PⱩG�e�?�A/E�h�I{}w%�c6s�y�r��Ln� ���n��O�+�f�!T���s1�nNu׫���\�q� �{=̙� ׽��{�I$�NH,�v^aZ#wy�/���GLN��en����w� ;����zȻ�������47Ӽ̣����<!�G~4(Ք������=�����i�{���e s��7���3���hUh��r���>��|I=⵼$���7#���*�f������ 4�;�߰'����y�z=���$�����&�5�;d�� ��'��N��Y�y� �߀o\��v-�.^kg�Y�NB9�^;G)��˫���kQٵ��y=W��HNx3��2� ��߹�� �K9���zN?o�WO[j���'~	/��ϻ�Iv����*V3#�w������<[a�_���<���ŋ��0T�O!v~T��{%(b�vb�vܵw���������T�^~��F^�+�>���3u���Q �����3����0'��y�9�_����q>Y�A��r�a�}7�0�_zbd�I6�sUWf�{�<�`'����	{鍒yv@,�`�ê'�����fB�|I%�qʄ�$���a�h�}�s�M�hTI���	��W��n�fQ5�6q�ޒI=��٤/�S����I_�{��$�{鍒 '�g;�~�eMa׻�?>e��w��,����Ok1�R��ζl����8��UG,�/9���"���*������$�~$�>�|�'jp*��2��{���@4^���i	� V"�U$&b��x�}ׇ�R.����yű�T&�4I���`D��̀�e_��k(�@=��ٙ$�C�D�B˪:@ɇ;̹� {��ő�����}�����{|�<r�������F��&��:v��h�T��De�[�Sqss��͈v���v� dYcuWKf�z��$�������OB\:�':�}�u�x���P��}�(v�[���Oioca
;��7�V��㔑k��`���# ��V%\:k-er����`ʹ���1b��/T��ON�	���<7���N��L�r��x����gD�粦۪ns�N�'o�|iu&���&@���>���N�5Oo&B�t�]��!��6d�.c���خ���ޤ���C��}%,�=�ո��c�*͍DUFoJ�pZ��%X�6��^�b�\�՛u4�ܚ�j�(�e��6�o`���4n+����d����\�$3�9V&,�5�e\�4͒��շΝ����N��V�d+��Q����,�x�VZj�m㝽�	���Uw��G�#ff��t�8z`�kw�{.�NΣ,H(���'�t��l���u�疷�aI��+U�Ѕ������)�pi��Z5�n=��_f����F�P?)Q:1ժ��٫��n��.[Ҋ啍Z'm>y�
��at�ֳU�VHu��.�*bN�^�B�/Rp^Y��vˊ�5���Fe+8d�V�_Tv�Uެ�{Tx.��'�{%V�Ų�ۢ)��S��]5*͎�*c2��̕kjh�Z(1 l�����>}G�qXy�̋c�*�.p�v@�3�P�Kokj���[d��d"Ee�q���d�˼M�^�]��ww+K�)�,n.���uzѢ9����_�9~�Y��2����&����	��u�����Z��8�4�s������Y��řGm�$���;�k���wee߷�@p�Dq�e���s�6�E�dE�a��tڬ�s�jYg&Z��3�ô���-�%$S���;Y�r�:C���8�8�]d��gZud֒J:.(��ZY���Q�-�.Va�ٝ�DD�vv��򽷞y۔]�YYM��IJ�9���v\V]�gam�.m����������fӹ.����ζ1gE��u�frG$���%ۻ;����m[�QFVDqqЙvVڂ���;���.)̳�՛��䀈������n�J�VQ��ug[h�8 �f��J�\FgKn+���m����� �ќ�\�m�����:mՒ�Df(���މ��%s���{��7�٭�w�f�H�)�����h�E��6I��XX������ܞ��$���~��ff�|ks�I�ğ��&ğ�'�/��}�ӻ�P:^ε��૆.;t�
H�Ս�����GI6�\��E�E��{�2�Q��������(�@�|s���� ���s��/�H$���;�䞚�yd���$��]̀��Π�׫h���>�7��o�[��ok����_�o��n��{�t��D���|�ܱ�q�S�Y�D/�;ƛ�ET�L����d4 {�o���	��6XߖnI���1��=��fA�{�o���/3puGH
��׎L��>���I&Ӹݚ$��}�fl�9츚�s/ox�ʰ�T��_m��{޻[���g�O�y�g�hhR��<��ݞ˷]��:�}�Z���}������eAT�M��UW[�����dq7ˈj赆���w{�	 ��m���G�eE�jC뻹1�K�O�^�ˢI;�9�I$��x�X{f��G��s�CL�8qUX諂�Nx��µ#��8���P\C�����9�����߹�=��������� ���co`-��0蛫y�{�X�e��d '�Ѿ��'�-R��HQ:k=/I!L���ak=�N� ���I4f�c�x�����{�(x}��eV�KET��v�D��IךA"|�����e̋RI!Q��w� Ak�^�K�0���`�*�,�o�_K�{V\���w=Qˠw��s�g3�c�l��n{*���>�Ҏ���{�Sʿ]�;]nC&h߾���|��Y'�ū� ����W�t�h�W?c  ���nҦ��{�;~b�4bp�֥k�1(n�<5e>
�s5�5nP11����)��su���
��.�\�Ho��WXk0-��sw�$bRpL������:��n�C�=E�c���ڗf8���A�n�����7 p/l�Ѵ]��]�S�f���Ov�ܖ�ݹ�Phy�KM��I�x+�`�uE��t�q�j�����32q'����3vB�pQd��ݮء7[�-��ҵ��a�a�N�l�vR��rD�϶#Ta։���^�M��;u��Ѯl���b�c��񚗡v�ps���sK
Z�;���W�-��Q��cP( UW�2��M�@3WE�><����}	��4J��L�I�L��2[)�1�Yׇ����BI&���o�O�f��KS�*�6�=܍��(�~����o^�h�D�\�0 �=/̀�(��n�=�޹'���"e]QB��x�x�I$L}Sv�H%��Z�v���$}���@�7��fjy�QU�V�@�"�_���3�'��D�و�&�5��� ����ov����� ����5���7���34�����h��9Xy�f�U��K�y�BK䒝/��j���m�-[���΁�<s6܅���r� {
n���^�3�n���s���y��3�;5�]U!��w�r�  ��7`O���J&�pBgy�{�tuf�`1 ���G��������-a��_��<֜����ܙ>Ywg�W�wn��/�r�;�X8�5�;�7�t]L��]�0c�g�r
d�WT����ν����H$�J:�N��s�$$yf<�`��;�$�M^��E�m��F�<H>��f�� �ﻛ�٠��Ǫmc��G�ϒ%�N��޹���$$pS$uE
'w��{��ތ�m���H%���m��^�&�$�F�z�K�0ne_�N[��ב���x>��4-2��d�D�%t�L�=^˙�^K7���'=���w��@ ���sK��L��sꅾ��qs���=e�a�h�ی��Ŀ�|��ڞb�y��g@W��|���5[��}�3�� 4�{��BI ��� �H;o};�.����{�́wEm.�!�����~���Ʒ[جS����H%�'n�Ih���d�D�����S2�oY����`�*��~�w3�cbA��/؁��㩝�g.����z����0ذ�6���G�U]`���ƅ���Q�o͍�]���� Ք]���:�;����Xv��V��'wz6��_=����1tUlF�'~x��rzfd�ݡ�۳�M�'��D���	�K�"E�
;��~������FJ�IV��D��<t�K�꛴�Lh�_9��$�?G�O��Wb'~I'���A����9���Lq2AR6�;z�<o1Ź��p��m���)]L"�teh����^q��uJ��[h�珽��������f� ��E�: w>ہb2��$�M�{� h_<ߴ:��B�ǘ��� �w�L�0�S'o���눲@�}��"���<�嚥��ĳ�޸X�᭠��D2a��fd s۞�d �~��͍��ٽ�v'�D�~/���H��1P��O�� �MQ����fe��s�����Ͻ-�	p��e  ׽7�n�$�{�H�>ݵ���Qk�N]]25�,}�F��������v��9��p�#�eV:���m��.k��tҞ�!#8��Ƹ �_(����eV�i� ��=�)�4���~���^�z�k%�;d��'�3ٔb{��f��1��"��{����P�7���E0�E�θ�u�{1�Lc]1��v�J��3˯Ͷu�ՒE�_���� ��d���'wp	v��_�+�i`�~�V��o�f�z=�>���V�'+ۻ%Bh�w���I}ۺs��MD�MN��`:'�[��Mr�I��sOiI��`�*��X����27���>ռ�BI ��vGV����\H�|o���}��{@Sc�d�U�Є�v���Bf�P$��/v���I?f�s�OĊ��m��iT,�݀w��O�i��R�?�;����`�;ۘy�}�:����<��$��\թ$�W�o��I��6{���7Td|��$�os��������˩Ac�.s�9�WT���Y��p� �	W��2�f'�;S�m�[�G��e����U��"��������;��H]cn�[���ۗ6�E�]�����0kx�`����v�]j��;Er��-n�w
mώ��.�]�*v�٬�xxG�ջs�����$����v�u�S����#��ձ>���[��8��� i������m��\[q���;��qy�:���d��l��N;:�b^�{Y+�ms7��ύtp�����g�ˮy�
@�5�T�������eEq�N�ƞ77H�]��]�/��|�]�؍2"����v{@}�;������g�����BDg��3@�/��s��R�S$uUB��C}�p�H�*�o�fv��sR�$��9��$�!��h�RA��$
��ҟfݲc�ٯbгuv��՞m�K�		M�D�M�G�������O���I6�=���`>9�F�mD+x�s3;ՂE����I�'y��B~$�$o�4�5D�=����Y*�>�ѸMM����UXG��{}�Ł�s��C	����l���k���BI"��S�@�;s�}�����Ȇ��Zs�kM�/Q�.Plf]�e�u�;�ë�nN'��� �HHHQ4l]Gw���HOs�d�I�}�؀��z������@'�׽�}�ĸa�=��Q�#.<H=��Ѩ��6�D��ݛ�*oϭJ����X�7e�$OnC��_��#R��y����)�7#=�^_׀$b�c�����`�c[F`�Wi}k;�,e<z�ÒI����I��y+��s�X�d�&w���>4гT#�o3Ezn�L��$Ν��I&���<\t��,`�ղ� W��t�4H�N��?zǣ򪢵l�Nf{7��ʱ|�>�@
��'L��ޞL2MQ'�I���y�~@���ـ�>8��UMD+x��o F��4Ee��o�2�4-�� M��$PK϶n�	c��b����Ѳ�?t����u؂f]���p��7�6�}Y�����x�k�$�����ݼ��	~�z��H$��l�����炽ـ��0�@!�����=���� ࿊Ъ(���Z��+���}�j�ym2h�I���a����(�pf1����{���ϳ;��;�ݵv2���w؃�@�G�T'�I8�Ty�ʽ�o�S�B���ގ�@��s�Wu�4ywUF2�]^!�����e�a�!��Η%�3�5�ujj�v��9$�|�H�w�7�	/�;gw% v�!q"ʢ�Q9�{�����E���"}��`h�w����l�����e��v>{�}@�������ꨭZ�DO���v1>$�Ml�3qzZ�L�6�(�h�t�n4�Ѻ�|q�7*V�Ͼ�]���1�a��ƌ����3�y��]�v�9s���U]s��;��ꚈV8����w��$�>��؄�~�����YG��$ ~�:I	!:�&�B��Xx��[���<�>C�w9f�&��:7*� T�D�I�r�f�fd�ْ Ϛ�w��Q��P���w3�`� ��o��@$/���c~˛8��t�$��D�57Ѡ��طdfe+(��ߒ����t����$���l�$��ѠQ$���F��v��,�K�8�<v�b<S���R�����R:�O�L-��^^eY�\D�vh��pA|/F e��I�4á`�ڽZ��B�z�v��5��_uɲJ$��X8��mV(D7��}��f� �s����a���>��m$'���	 ���n�)$�Tݥ�d���3t���uP�~"��m�.ͺk��ۙ-�����C��ӽ����n�:���c߼ʪ�!DN{Gs7��a�4~���|�	!��5hH���[��w �;�ľf�uMD+ �;.:�`uƆ�v��X�;����4C@o��ɀ�w;�j��L�^�}��2x�BB�$���4�ބ�{�,�$�>�~n�$ոU⒦�yg���$F�wy�� �w;�ŋ��/SPQ��P��{��}w=�޵�('���BI$��3����$vQ�v/+C] ������Xݵ���;��n�h�{�9?L�ݗ���xwU��H/>��)Bz>����_��d���iSa��QƸL�)��w�q1���V���Yʠ��I�$�XƗ��-hw�����ʒ���T��ʻ���U2s�co����_9nă��9*p)V.����Gyd���w]��gp#jSB�pazWr}G�n��&|�U�;U.��*�̈́�]r��k�լo�%%5�UÚF����L�/�P�K�1�ƻV��d�ļ�l�KE�:�h������W{)��<{��8a����%|C��+�v�`���8۶N��z�3\�[hh�r�YQ�Ø��ԍ�H1i9tvJ{���s�)�H�f�%�<���	��e@�f�m�U��-U�����f������V��M�u���*y1�o(M�FM�^�9{j�ذ��F����RJ��d���aoqNnu��'�8��m�8�<6��ղPl�m�ְs�hT6�ٰp�Ǜ�轌,�lW`�j��N��͍kw�J�fܳG:�1^�G�Y�����.:�DE�ܸ�0 �gd���BƓ��:�t۾P���7�W��Q����[iΣ[��Gpa��Nd<����;���o^�sz�,�ˎ����)WE�g�=-V�-�znu���}�r��t����[���I&�8򜥢�7��wy�n�x��Y�[�O��܃[�$\��ʪ��\���6=NtM�B��a�i:s���h����,�r��a�e�t�y��;��q�*��s�-�骵H��ӎp�9�8���� nN��8l?[��y��ۓ���p�mm݇m��2+mqEed[k8���q]�v��89.+w[d��:��"3(��.�9"��m�w�rT�AEyy�wl���J:�������f��Q�Bgm����)�8cZ:���.�ά�8�sj8�ܮ�GaݒvdR\Q]��RQ��]V݃++�:�mVq6�ӊ��/+�����<���:�s��+�;"6�ԉ�sh���J���q�GEݶ�����\%qm�mVu�D]"gVY�G\v]gG��gti����m�>|��*��8��ʽu��q�n{K��_;��k�&��<��h�N�f�q�'kr�ls<��V{v�Ay�%{�m�n��6{c�ٶ#��g���=^��v*�4�x��$24ဇ�a�S�D�N1o#/Q�=l��C[��N�kcv�q��w�u����01�w�GSí�)g��;��'��s�l��N^�>�	��Jv�v�;�<�'+5���t��c1{�������ܩ�rf��99]aYn���8�[XG��M�mQ��ۦ=��ƴ��{�L��Y}�������-Pp��Ƌqu��$����#�6�b�ڭ��5�c������Ó�ذ��{���Y��źL�m�׳��hY1ٴ�s�:8��mn�[�P������4���u���<od,L=�fy��T�F�oa���h�n�`��h�s.J����q!h�0OX�����U�ddQ��)��؋u��9+�v�Oc9��q�݂]�����`�N,�M��7z�α�k���Ȳ�j�Z\� ���ӌ��JwuŮηc#:/vⳭ���2�m��6����c��m��{k۱Q�z6}�^N���c�T1pOe�Oe�u��l����t���ph�_8x�-�N���#�k�����-��;WKŪ��í��	��	s�Mt�n�R�q��#��Ș@���|S���[q�x��ÎڷU�����lfͭ�wl�Tg�k�۞��l�v�Ӌs�t�g��n�l\���˞ڌqkn�,�U�έvx�rnݻri�^���y��-��ӌ���[�w&�-��u�z9��C'���=�x�:�<4�ڎ�c�!�^cs��=��7a�^wA���x}�x���qmǰ��#ui]��l;�=۟q���om��ġ�T���	+;d���m���7Gg�ᚚ�p��ar:m�9��Z��P��lK\�\�sڭ��x.{t��3>5ٞ�n	��b�v���O���������[qk�6���q���;��	u����G'vۯ\�vr6������&�rxl�	7W�u�-!�����1��v�j�N��l)3�8����ݤ�)={�q�ib��vu �7oFu�;l㗎�N�n{N���,��F\�S���۰v�[��Ɲ�f�պ����7']�|���t��u����IV�7'��;k3�*X;gy��:r��Q���Fx�C�Y{rXVz�����cx�c�ń���K�]}ηZ#&���z{1@@����$�����=�p��p/:O�Sr@#�߮b@z>w�����J"c��&�P�k�f�X�[�_�� �O&j�5]��$$�(4�S���RȦϾ�*��5�f���� g�c���I�u�.����Q$�M��Б$����{�o@����.#�����:�����J}D��~�L�I>��H��f�����e�߽8�YJG,�$�o�bX�"�8�D9c2?���w`�D��� �u��ܴ��D����;�lnQ$�f���'��k�1y$|(
4�1������답:��F���<� ؒ��Ȓ��7���7mCu�_��s=ۚ����>�lrD�O�}��& �{�b\܈�=˘A�������FEM������ [w�ًɠ���A��/�"��/n\�������M:�J6nv��CO���U�x��X����my^�����!F�%2i$����������PI��e�}�]�/���Ǹ�u,$�&bG���{� �{~�  _��^Σ�[�A�{��o{�=��hc�%�E5솛%�����Ya�3�I1l�BI$��Lө ��y�����
�I�e9e����w������P��\G=̹�i$��z���5V��ǪjH����$K���RGϽy�.�
����Ae�����b��E�WP�Z��nCGV�������nn6ú�!��.�#�NQ�ϣ�w��k` o��� i ����x�{�z�{����4�H$����5��i�w�������cd�+b�+����~�k��@��y�6�{���@��9��s�Y=�$�(��������ߖo�{� A�o��y��M��wg,�����:�7�)�ip���B��ݑ�j�b����D�d��+F)�	BJ��Ԭbܲ�*,}��56����'7��ӯ <�{t�j3b�j�UZw����\n��su� �ͱ��d�M�A T}��Q�2�ΠH1��	��4
�����U_[̙��s��V�s}O�~}��������ϱ�;���پX��mB�\tNe�q��uu�Mӎ�Fvv�)ө���G"����|�x�	+6��2<��v��4�Q��p���J���(
�}��t������X���=����R������m�5����}��%;M��/ٕ��n���I�J�G��2k��7�	�o����3������n�A"���$	x�k믑_P�y�g��0��I��&���������*��Lw���"4����d]l�êe�]Q�c���S��	���>'���ȤM���ʛ餒�T����3m�a���]&�����}t&��W��f��F� .ي��ܗ��t��/H�A��^�v��ޣ�@"�*#6ð�]M���;m�������ν=񫘸Gs�=d㳫nޮ>.�?��"�����4ޙ����=2�������<�?����t�t����a$.͢No��yxH<rU�^oܮ'��n�%G�}�'6[_l�����Nw�ծyH!�B�eQ[��  [�� ��"�w�u����~'��� �����m1���`�o����1p#�4a��پ_:�e*�(�����z��'B_���z
$�E����}C���:��w�̊4t{k��H�c�fn��2>� �����W�FڵJ=vz�)>7�W�&d3�	���lS\K�N&Q.:=h��{$#/�v�#��m����V�V2�-8^�D�!��I�{��S6WΎ;Pm��5�ƺ={W�ئ��GG1�X��6x[y��;��/]�g��1�۟XAPCHB� "&�%�M
��V��Ӈ�}�,rs�m��t�:�%Bc��>�l����m�����ݷZ�Ƅ���p1#˜�g���p3}�r��wA�?���ܸ��`6��k�7�q��|���;rh��#���+Ok�紛��KR�z���[k%�s��.˛6���[1�\��|Uk
�cu���o{�M�֚��@PW������w��v���%.������O�ޟ43NMɭ�_��*�~��.�l[�^ފ|튕 �����5��
K���P�h1����Y�~����zO���� P�wS�,��Y��N��P�w��boY�V��r�>G��s�W��׍�Kω�5��A?(��2��Gñ#G�������HfA��*�t�7���ʘ>�jc��n2�z\c�:�|A�st�Q��UB�o���/v����1n��#mV&Z��h��C��n��׌��(MK�UE	��m>3�6�A���1��H;��ߴ����X������A��M�|�֬X6,�tM�����\�Z��w���j]y���۽�*夹��Z-a�����T�O��p&���S_`Hu�w�[���v�Q%�י�W�؜�f��g�  �����}܆۩�yN��o)|C@�)ZUC>8�ۣH$���I$���+E��W��V�H$t�{t)��O]�������_bO���䄫����m?}{��H$T�O�k�Z��֗vo�O����bo>u�uG!%�
o���m��!��ެ�]�l���	Gɀm�sY���ʼ�������<��R��kc��]��0���XC]vvyv5�j�mm���OT���f��ś�������{����)P)�m�������0*[�ѢJ$�Zh�l�����;G�(��<��>i��}�&�$u�o؟��/���`�����Bȥ`�[�[��uA���P9�P6ƫ�z[�[����!S�}�hS҅f^z�]�ٳ<���k/D�P��;.���'N_<�]�9��^�ݫ/�2��_e�ВCמ���u�a�ȍ�I+*�aɞ�򍧬�j�,X7}�� ����`�H'�}�U�7�����$��ۤ���)6Uj�7K�/�:{~����!K�����f�A'_��~�=7A[[�{��|q��@$�;A��`�YT�a���;ٹ���u���mV*�����s�I��r^P6}Jw6� (9�� P���MhAV�q��1=�������xO q�5D�&�*�{~�gH�ջ]R���m�k3�R��|�*�c����Nk2��$�I!���H(�9r^Iݞ����f���ȩ�}�
���I��{;��7�q�{���9QY��fg0���I�4���yr�I#�$����kbEf,^֙��i�[�.9Aj���!i�-=jgn���@��pt�"Y-,�3S�U�P��56��jX���OL7P_��{x	Y��S��,������Q�>}tz���(ցTT�HP^�����?��R���}#>�7ˬ�M D7l��PD��5��t�W��%V6�{x����:�����ܽ�]���T(O�x�Oh�I��t��^�2���xA'='�@$f�6��*��g()o���wuL~]z�z`�J�( )o{��n�7N����\�7�a}���7}��e�D��.b|��?��~i�@P����=�3{�N(�o�t{���D��c6BQ8z�N�is��O�^\�|�����O^��a��ʛ\؜m�^�t�c ��^��j���ު'<����`,^��A#��wA$�;��P�î9��>�j��k+��vG��{=�|�Y����8���C�v�pM+"�^٦�����ӆ�FH�^^�br�tV¨U�(�zj�.tQ̛��pH��]j�YD+5]>6ڃs����pP����K6��;�j�K�.������5���1�n"�wg���ix�RM�;<��C�2�9�V��������3ө9����g��	K��T��H�RoV�����"ʏlpj9�� ��7����:��5��x�[g��9�簸lU�z���[p�ܓ������wV^��._u���a�wm+\��I<�����3������t}w������i%f���c{�sə?L�[8X6�{dg��� ���~�EP�a%UthP�>�� �t��7�<���w�{��&���@#�F�7*���;3X�`�l8��¦R����6�{ߧ>n_�՗"�1A�: I��ni$�;��w]��dTc����|W>����D�k_�4�I>�l�$��N����L�u�yOǅ�l��X9r�"͞����b��N˧��w>� �I}�x?�I顀:��H������+�A%̍���()TӮ�c�e��8��n.^,Vm��sתV�6�U�4��yy7I��g.�H"�Aݑ1]ĩo�I$��<D�<G�J6����:���}z6/d29��"b*Vx�9�4j�ގ-���J��wz߫<�u_z�\�/0QƼ��x�ٍ���9�˨o"&�x��znh@ ���U�=ٙ���S#�XT8�I*�(P�>��?���߾#w�:����$��20���w�pi��*ɰl��M�W^^��Rh*�[�A#<���H�����~sx��'m��jg5�*�*2��>{�{1������NV��!΅C�տ{}�
�w{�ϖ�6kFfz���߇EA�4hѺF�%uIf>�]p�oh�\z����@ݍ0R��$ ��&ޏ� �!D��T��?��H"c�&"��%~� �ZG�Z��l
�oIv�V�T��K�9���|�\/�:�%N�O��n�L�~��~�ٞ+V��s'��U�c� &W$_i?�=���A����I&�oU{N������kٻ#�5����yE���	��������&��{�G\ˮw�C�ʼ3[n˛��xv�w��/u�Y+���kq#ӕ��W,T}-K���J�?]n㡘dfS��]9;c����F֬�.�j��ۗw�r˒8"��4T�/F��/�����AC岠�wf틧wl�[
�v��Ц�c��wB�k�r��QtmK�|��h$�_+ڜ��*,���yؐL��H�e�w���Z�5�T����ZO9�j��ӹpgE�ڳ):yҍv�t�^�,w9���"�-6���$
��:�H[;�Zu��8WV ���_ogcjZ�S�nӱe��t�۽Z��m���*�$���EU%Nj�-e&�%K�6�A�VG5g�j�Z(�̢os,�_���;׈��D��3-N��ʊ��N$WBe�gJ2��YVz�i��/�E8ZS*�_tux�S)7h뢳j��wvV��W����H�/o����Z,\�ﱌ��9նq�)�D��·uJ�5��n�kf�e���V��]�&uvQ���I·VlO6d�1�&��f�L�kE�wܫ�s3n������T�Z�I7x��A^X�������1�Ն�fꡑsf]�/����a�eJ�����Jy��E,9+#ޓPS
6[9�h�ҍ��5�(L�e�W!1�AmX��hl��Ù�@C}±I�\w��왨�#�V;������Ǒ������iu����\l�{g��ge��kU&tbe��u��37gC��д��*K�2�fe�����5�	�ʤ�z� �&���mY�wQ$��ݝe����tGg�e���ڬ.*.��m���\t{^{�(㮎$�ʤ��N"���wNTA����I�����9,������m�A��w9%�eYvQE�uQ�e�YY�9VYp�Ol�.*(N�9y�8����v�:�6��QPwgYI�\Y�q�S�$�v�h袢���AEA�hw!�RP� ��\Y�e�c��8⋢����dw%�wGr�w����-NX�gTu�N�QvDt{j�f8��:���N����.⎞n��H.;��m�B8��{����/�H��7I$	X��	��l$�X�(n�g+��2�l�Sw���~$Y�� P��t5sJ��q�T��kt,v�F��*e)���&�O{�σ7-��~�t	}��������ո��|���.�����m��"��2���ŭ����l�=�OWZ%�����]Q�V�&{���E��2͛�U:f����^�� ��Q�c�L���ɷ��٠�Hu���%|@-�- BH��>AgW��xׇ�����	u����A}�����z����^������DX���VV�����	��δ� �L�ν���X��H��է "�ZDF�Y�����o���e��Æ��T �\�(l��Hs~�_��+6�%�U��Q��.��d@�����=��x2�~�~:S�V#�\l��AS��q��免}�r���W�r�#jF������n��Ǌ���	T_b~�'��f��K!�e�o�߁!W���I}+� I��{t�0�S�^��4�-�eR��y�����n��m��gm`���iv���`��*e=���߉���x�c�{t1�m��(����I �t�")Ɩ��Z7J��7T=9y� ���l�I�j�� m�@}@{���𻭖�^�Y��/Y|����|@8��(G_� ���Ae���T���M�sH��n��溢,U�(ث+}��#�^^ߦ��e�F������S��n�P݋��~�g�G��?&ݜ���S��5�� �H�k˛`�M�i�	��N�{Y�_	&F��7�̆�ϙ��@�w��e��%�O�^4G����vU��A>��}��:��(=���b�Pa�fW_y��;��&��#'b�Y[�#�Ǳ�v�	�m�����6�muN��]�f��hgqC}��wK���X�`�7�ڏ��3�5�����ݜs�糷]luPv��uO��q۞��"W�|���'[[��4\/>�p�;k3����;cR�M�qܲ���:��=�c=�i��3:�Kǎ`�4c���-���3�Rp�,���]qFx�NxHGK��r�h�N\`���.�Ӳ�� vn���E�'8��%�.7[__���M{$�[ӆ��<�j�#Cc�s��i��g�t=�6Q@��*�@	��6ƥ��!S)���=���d��c�r�|$���o�}�� �$g_����z�ޙja
QH乚~��coO����H7�:k�
*^^�����$��{w~<aa�H���p粦�^�ZЋ�w���:n�$�:|�ޝ�{�M��I<�"�Y"�*��G�u�G÷oQn�=ؘ�)mJ�l��i�� ��<[^�Y��Q�1�ϡ&�*EfK�wg[��v]���sMs����o��ڀxvz�O�ft���7�W$_���3��=��@$��y�8Z���k=I�w���H$s�wA>��h��]$hn�gJ�D��7�U*v�x���B��(\���Wu+Z����Yd��a�([�W{x5խ����e8W̫�}d�'�9�Gc��{��[��i$�G�4y��	������ǐ[�L��U
�J�XU.���
��ު40��o�2�8�龍�(=�������egY��^����ޫe?m��_�Z��?w�2�W���N�@��cu��`��n��!
 �vB��ir�r ���n�����2�+@J�>� ���O �z9��+[�Ӟ����w���1
MW"
�d&l��j��l�4��$dJ�����>��Ԏ�[	d痷����k����M�z9��s{���{�=}���G��ϑ �d��O}t����z��	�g_�=쭴�f@~-��G��n�E�I�K�o����ܻX��>2-�J�#��iB��|��1�������y��,ڬ*���o:7b0WJ�/d�:ؤ�^�j�˖�Jە��`@����YL枺�L���Y��cĂ���O��I�H���ZB��R�`�X3������Լ��'����I?vG��� ���vh�d�d:y��H4�{��T6�&��T*���d���	>y��x�ҵT�_6e��	���t�_��V=��j�.����8F᭰��M��<Plm���yx:��;+
�]8��4X�UP�3���{�I�֯��c�r@o��ƹC�G6p���3kH�^I��}���!EF�Il���s��&q�{��\$��������ʝPW�<�aP�=i�����V�I�5��־��k5��X66��CsO��$�Z osb�ߗ6y!�E0lD�I��z�O�߼s����?y�ti���y7A$z:�]�m\7��9߬��K��7&��v��zJ����vϊy��,���W]���u��u�u�׊�ik��ӎ�X7�m0�-ϻV5�?�Y�wF͜�p�~��@n�TM>�P�dMY9+ �;�~�d�$�GY�!G��bʾu�xw��������62���=�E{��E콍ɄKcW[�#%��j����}��R;��7{�DS�f��?���!��
,S/~~Ǻ	�^ٺKB$~<ͤ	H�H{.��*;̚�Â�[�4�O�׶f�A?GY� ~7�3���UW�}�0H����e��~Ԣ�N�H��X�ym�ێ����t�#�l����u��#�J�"���PÔ��=F��V��Us��P����(
��^$��	�~����F��aT6�(*�UT�@;%f|#��ۣ����{~�~��$�n�� ���������X��3���)��367�o@��d/�e��jk�SNUH�Aʝ>�ԋ0k�~dc7LՒ�����D�=�tY��&���
��+�]6�Lvg���:�gq�L�usMf ܮ��ayޥ78�Í��.�n�n�����ڛ^b�6ݢ�lK�nA\���u����u[��G�����g|خr"��f��N᫹�Z:ٸx�tn��@���f�v��g�طL�[��]oڴ+�[�q�8��w�l��odͷhyv4�mk`y��vi��j�y7`��2�R�ڳ�qv������A��a�vh����@�ڳ%"#�����==r"��S��߉#��$�1�۠�$M��s��� �[u����$��B��ߏ��k%���V,��@| ��a| ��`.{�ec�*�s_|H�4��1t�(�I�O� ���4$� ��׵^t�f�$d{y���w��s��8Q�k,e�cu�݌¢*8w��|=�v` �9���$�������#��N�}��~m5�ّ>�j�RM^z��zn�Y�N��vqb̬����O۾l 	ݿn�������	����W$*5]�(70�sj��e8�]F;����:vm�_�^k�^pEd�����zM�w��k?��~������}��+��ގn�X�I>�8�%���K&sٍ�c�8�iG���ѺG�f�]��':��W�廳Ր�����|�Nؑ���g3G)�Y��b�:���̔U��u�m_� ��q��IM�F�2�V}7~�����2���@���}�cm<�{����]��m��]u/V��P�z9�I?]7���D�ڸ]/��Xs�Oά��$?��{�� ��s4�Oǳռ֭���B�$����!$1F�F���~���߈&����	Aǈ��F���/������y��=��-��?��v5m����-	�+�wK=XHvA��To*����Ujusi�������j︽L 2�y?��O[
���vr�}��wX�}׭��]�س��5��M�-��qK�;b���:�����i���@m]�q��\�d�Z�}]�b��������i�����6�>ｕ�HD�$�LL����'��J�[o��ӡr�E&��s7()Νɐ�C|��ug�V����R06|�'�A�q��\%�Ύ�S��O�[�� �o����6�y����t��g=�7���vVA�|��${���MǷ�@���kׇ<o#K�PMi�CZH���Q�DܻM4���qb�_�W���,���P��P�=�N���w��~�n�=�[u��Eh�ɹ��W��s��I��ٶ�B)\������Ttj�e���� S�P }�s�a��=��X��[�� �~��O�g�K	�/��
����¸T�p[����ȥ P�ޜ$��{}���}e�^#�%�����`�)b�zg46߻��,i�
2e��=��Uph������	3�~n�[�6VY̻ ^a
�?.}���(\Q��G�=}^#/������E�Y�>YH��x�l��J.��Kt]�����n��e��ha�����N��+e����e�5�e����o�����w
lv�������F��ܙ��͛yN��{��>��́@{�sg��;h�`ʎ���k:�IQ�]Lu���ӐD�n�Bv��8:�Ӓq�m6���j1��y�d��o=������6(e���Y�@!ح���}���#<�mtn��v�������y�Ym��#��w�� �%��	���3��q[���ӞM�k�=Ki
�.T��d�'�A~��w��H�����'o��O�d����%
�E ie�%����5~s��*��w& NK͏���S�i�^�����?s�T�A�e�˳C36k�Θ�-*=Tp��f�7�r�w�_U�6<�j�O �$��HH@���HH@���B�I	_�$$ I����%��BB��I	_��$��$$ I�HH@�� $�	.���	(�$�I	_�$$ I�B��$ I����%�RBB��$$ IbHH@����e5��^����!�?���}����u�# � (�P	Qp�(("@����     �$  �vf��)K��:b[��{��.��9�k{�HP@��E৪K��*�;��Fx>����ϵ)�h�å�  �{�U ��:Q�Wl����v��)nwUT:  ��EvaŠ3��@�;/x䣼�)RUC@.9���+�Ð(4nL�`��ʨ����*T4nw;X
{c�    ���Jh       E?F)T�       ��T��*��dɐ�ɉ�LL��h`��ȩBI�       ��@�UM@ �0�� "I2hDh��@��#�z��4�#O������Z'J�y� Pbw},�<�TA�?��P�(���������������]!�Gxb�A�@�?���F� �"2	�P:�qU����{��/ר��5C��ͥ����ʏ��F�l�E�s�����P���J�T�k%[j!N�M�e{�D�ʕ(aM[�y�!����~����V�P��I^3B���%�F��nfn��vNS�]��aTV��\���i�<��8��5�H�8�PC�[z�&:�]2v�[[3@�͗q�KLї�@eAqAm@Đ�/*u�KI�K.'i��w��^^ءr+�ņl�cM�I a��L̛.��g*ٽZy��$9-̬k>{{��n�G���SR�U���/j�kN�rJA�O�Ē�b�X����he�?K^d��6�&b`�%\96SH=�Wf���<�-fC�����6���ƞ�n�ZԲ��#��3N�9��b6�&X�*AL5x��z�,�AY����v�'���WJ�2�N#�mo9W��کx�e�����%6� ~�n�ѵ%�T���R�Xyw����8�S�u��b�S5��V5��
L��˷�졟
Ͷ���v��Ñ`uA�R����Z�b�g�[o�swhڱ����`��f�x)"�5^Zє�I��N��n_����x����[�:V�N63tV`����ofL��Z�75��@h(7�,�4�Vo.b ��nc�p,lP�����5�j�B¡f�r�mC�Ĳ�b��[�m����8m�n��D�i{9���Z�x��+���ᙊ�$��T�b����ͫ˨����ּ֒�/J�[�yn�Ř��u�t.����ᔖm�;�r�5���m6]b�XǦ���h껁��3���{�!�Zp�&���{�f��{[r��[�j���t13�r��k4TmA��th�Ȃ�y����{PHE�C	̷�e�u;P��;(j��sa��nQ�k��WY��R,�,Sm1����7V��E�g��%nTa`�6p��nչI�`�.a�@����	sY�|�.���P�d�/E��v�JˋJ����*Y�0ܫ�������)l�{(�,�s��kv4n���\"��jȽl�5��p]�:o)n��7t�in�a�� ��N�Ҫ�n�QQ�w���	�|���V���n�ˣz��M2���.�,��)ET��T�*^,q�e
��mCt~��Dim9���^���!��7f���iрV]��Cy�2�Kp�Ŗ�ٵX��n�gCʱB�պUe�N�[X�]@N��맥`�hF�
ǃ>���B�I���/p����"��()�%5`�%�j��;�u�hX��B�͚1S���{4���+Ro���l� �;Ӑ�a�J�ˤ�w�$��M^*yC�"'=	䱆f
b�(�UX���^�J�A�or�aY"�:ݵK0e<��DCk
ÛXĦ.	�J/���r���u{�[�zm�S��9�A��n�����[f��m��$جmHE�y*�6)����/P � ��5Lԇ��u3�걇I��LX�_pi���;��k�0��6�H3J��.hXN�E}�Aj(� (��� ��UI**� � ,������
T **2((2(H
���"���xpylm�������TQ�Hm{kqy`�@�MOQ��A�=duq��4/��kq�Wxr?�����]��!�C���iˮ�LE�u�� 7:-�<o�n�Ѷ������b�V�VU*��#��A!`GF��u-iyp��6��͹BaIw|cX��;�����WR"B��SE���$�\s��|=&V��=��t�f�:�u�UI'vo^��f˓��6��]9׋��Ǚ��1ȳA3 �p�������99�6r�� �ĮWd66��CPo'+�% �
�j�lڐ�N�Ӝ��T(>.!�����C�Rj+~�R+sj��q��� ����p=#�UE`E\U؍)ub�;��_e(G;�v��4뷕Ǵ����n���Fm��AX�/)�ac���h�5fң�ާ�oZ(�Fwb�j̹.`��&�sS����D]H���)ȳ�VH�Ji0Y��F�r��nj\�ّo4��B�H;:��Ԑ頩��ݫض�R.6�N�K��o3s+3�Z�uc��)a�/�4wWH��e���坧����j�!�`��ō��"�&��_b��c�4D8��҂��R�3`ը�P�~��\�hI���x+��D���j���V1X���p��4���x��;�P����IK���6s���6��#�W:�X7��#�bn��'��%�CV9i<����P�P�y�D�������3�4j,j��WGv���+�̊N��4�V]e5�hRˋ�Cwx�5m�e�;}ݚ%ʕu���;3�W]o`Zшλ�:N�����[��܅��:�m%��l�m5�!\�g,�Q�i	,�.���#7��,�ͦ��ۡ.�F}v 9��wV�����7Z4��U��]��`�K2�rU��a���]�&���p�]���̂�r��:����fY*ZPK72˅�B�-d�>u��M%��"��(WUÃ�{*��n�Ŵ4&ܑc��VZy��G��;�e�`ZB
�['@�ݞy6�k���`�O0�hȳu�=�w`[𕉭}����j��ݠ�tq꼎����]�V ��s�5K�S�`F���ҹ�|3��2��Ӱr�� �m��0��i^KqE�N;N�J�_8M�kథ��Q� F��H^H�r�5oL�[n}Gk�f>�ct^�b�(��Ķ�]�wx;��Ǯ�+��ޝ��8Zt�Kb��fZ{\���x&��p����ZN�&s|�a��W,����JJއ#�ZXZ(����+��i�s�͌����L�N���ti^]Yʷ�\�Χy
��:��w)s�&�)��n�\��V^�;�W�r��ʺ�-�V#���X�?EG���0���1�����Br���1n��#qδxP��l���/vƮ�{�K
�:YM���;�������n]Ѿ�,  6�wlN�R��[�*N��������cx+��Z�p�NȅV)Pd>J���tKݷ��j��\S�c]-�l⶛X�!�@Q$I>�5�K�DG����> �_M�	�m�٩�n�K�j&]tPb���au�d��ve�n����J���r���c��h�t�`k{Z�MWjZ�l�M�f�ݦZ`����q]]�q�q1���ݬ��e�j�t����٨�b'Y�&Ʀ6km��M��m�)m��[�nc����K����\�VŶf���YI��Li����-�V��么t�Ղ\�]+s�m#�-�b�GQ��xn��b��n�2�էl�%�S[��m�u���Z��a-��4	�����lkVi�ɪ�u#kf]j릺��ʁva����l��l��
��ڡ�l:���[��Cuc0�\��8�7]��nة6�Cj0v`e.���m���i�d��\l�7�+�6%6.l�f�GK������aM��ٙ�i3]�ڴ�.���ЮLؑ�m�J��-��jhR�.t ��(jVfG,��H]��x�u�-�[is6��gdMTF�!\:�fiB��G��X����J�S=�2�%3�%��Qֶ�2�(����Ccrn�:�j�N�a�
�1).�����t���î��)-�٭���ؚ6 ��ƚ�h�#W[lΙh�IW��;K\�ʍ��%#ɋA�Dճ[.u�\+Z�3��`#��I�Lh꣭���JgF����۵]sҧ:�0Z����&�kp�Z�[,bSif3��kt:��ʫ#��jjЫ�..�]v�aKZ]���43���+F��,���.��3��%���C#]e�-`�Xccpإ�%�e3����ˋ3�Vڶ,����	.��k��\�݌kK-�e�4��0b�e��v�,۱�K#�h�*q65`�;�n����t���ʚ:Y�ť]I��ib:\��k���c�A�.�۶avui�s�ɮ�iP�c��,�:�E��L�Q�`5K!+��)j�0V�����m*��-��ۙ�ce�e!n�%�u��6���l[�b� 8��䪊��EhҰM
Z�R)I@    �8   %�5�v�#u���Z�.���Pԅ��:�R��p:-��۴���]���([6�k��������N��H,	崀/N b+�WJ�y��ũR*�+��6�AA`��9�ʐ/	#�c@d��̡ J���A"�*(F3Ŕ��t��Px�N0����Y�]����!��V�.�]��k6��U�lJ��
M+��Y�c��6�!�������ip�����yHm%�qk�VWȔf���8�ɳ��6&-�4n��&�T�IE3��m3qfHZ�a-i!ce����#f��R��:�f�*����H:R���(��L1�J��[AܡT�e�P���eI�7Z$x�������5��*��n�v���5�:m����	��\c�A��[i%PFR�j%ib�U���F�-���ƅ��j�}���߉�ܩ:���J�I@����,�����D��(DnJ�*�����{7��G<-4g/=��Ɯ�g�*B��(Hyw�z{�e�m	E!3���6�Ќ�%�cG�1�'�	;��i��?	"�N@��=٢�B�>8@����mN�s�c��%"�yq�p��, D{T���"��إ�h(z���(�	�����N��l�p'}�col~L�
@J9Gkw��l;1&��4Q�A�׍��/�Տ�D����q4��JP/�Ww�]�zx�²z��6Ur�����{�ew��DLHCe(l(��<t�<rm�L>�ǀ�~�0Ze��ǩ㽫ʱ��{�<�ł�w-?w��h,J׫&E��f�O4�g#cQ*᜸x�{���7w~�]��b�������z�*Y��T8����Z�o�$�
J{��F��)>�lz`�����	#p6r$Pq����ir <&/t��۩t@��u\)�l圱��<�]���z�Y3��$�	��A�Hs�����hR��VRJ[�A�h�:]mJ�6��v$��m6��v��$��#��@efU�(ۀK�W�o�݊Zb�A�)9$�;��9x�D&Q���`�t[mR�hE�+&�^u�b%L(�.f�L��b�3X���Gw��uHݱ}�E��t�ܼ,Nn�g<(:P��ʢ��BZ̉��/b��a+(^�V��j�m)'��q�Z���f�,���w4bg��S����]��c�*>���� a�蹤��
3��٥����/Tȍl�9P�s���}|���P6��W�6*ΌTl]J� ��#Rr�>�v@�	sy�y"�ȹz�J튽{�Ab��b�1�&�Դ�Q�BPr姞ݻ��&G�sŋQ��ݸ�s68.ȴ���j��tYn߲��Dp���Y��9�����	�6[+�;V
<D�iDE�t�G�p&j0?E��B�1�V���s�/#�S,�7b�p���N>P��fp�#MŠG��I2[�RT��j<�O�v6�����O6�,�H@���Kؕ%5�0�e�59��	`\%:���n�`�Kkm�h&\_f���� �Q��t}���b��G:(B�3=j���b�����,�ow��ב�	3�X�+�%�|�Zg;o�� I��q7ȉN���B��g{�����hk�8E�]����E��x�mXk;]��J��Q��D:qǪ	e��<�
o��w*J9,Q�ٰ2Z��Qqq�|��������b6+#�}�D`GGa'sy�L���45�-5%����(��:"�/]����*$���i���<N�C��v>��"r�^�w�M��e�>5�v�dk#�9��G=��� E��	t-�絯E�v��|�����O{_*�\9�6�ʸq�ґ�'�o_����ՌA_'�;*�tH���0^�\��X��'tצ�pn���e9
g�iZ��Z�#ء*-�bE��ǡ��X"#3�zX@�
�E�C�D��$ ���"��E#c���x��r���a ���Y�R���q��!DTP B ��VC����9P�$AC�AQR�'@ P`�b >���������r�9P���#[,|�V��=�$+/iA�0��ɽ��"�Bgϙ��$�m)���)kuܴĬ�	E���wgj��1x�|ߵ���xg<"3���q�`�C/֮�ǁ����&��FhDu��T8��c+he�>'�G*�9�`�e���L	o�/y;9E����1�ُ	x���Z��}��>t�Iɖ�w�u�D�Be���	�O;l�m���%���m��KUu:fW�8J
�(�I&'1#�d��/4���҃cu5:�D��:�iq����[�2A(����h�<,mQ�(��X��Y�r�D��T�3�����tK��@KL���6��,X1I�Q�{v�:��<�{+���`.�y����K"x�aBf�{X�F�^�}$VmW*pL��̛�F"z����9�>�K h��=p�j0H��^��7�Ҽ�}��Ku�rk{��dV������kn�d(W�Euj¥)g��R����R�޼m�Nް��k�+�J�^-���P��v0*��Ѥ1V����������ϝ���ҷ���k��)��eVNK�֙��r�t�*y��6F������rqwDA�H�2"Mɓ�uU�4RFf#PNL8,�f���8�hn�!���T{nl�\���.�;j/�^����J����~�~e�ޔG�S��o�]~��x��$�'�Q;n^�n,���[���8�KK+�����0���M�
�7��ޱB�E�Y�a�/��*�Z�i]�%0�%w{$��o&+$����V��`�ʭ���C�ʉK]�$���tc:TCDYk���=���5�w��ͥ����ko��2�e��΀���:��n[�����̀�l��e���<}�B��+��p���zu	mӬʟ����8gp�}��{�_~���&?Y�t4͒#W�w&�˃&rqe�Cfe�4�w���B���T���YRߖ�Y�Ձ�{]LI������TD�RH�b��������'r�$��X1��m���4�I����o�8�Q�tE��ʣm��9�nj� ߣ;�NjyP���!OD&G+��CȲ2`I���ʑG��uDS��]*���4
*K�S�#���Y���Y���lL�T�����Sp#f��\���<˴�]���GjkP��v�7�
	�r�̾jundxs���R|���^v�{w���2��mڜokz�\T2�]�J���W�Fgi��5N�Ļ��}�5��Oꯆ6�� H� B�C�9�:��0�/D8�=T�a�c H�*H�� �V���f6B B"��� "Da��H�sHE'#b� C �&b�/�f�lQ����l],m��^ˆuԱ��Qw�R�����Zd[��p�%��-ŗC:j�j8��WM 	��v��	e�l���r��42�]��؂�67B��J�m�15n%&�����ͽ,��θ�]���<�̺Ų�,�k� E�lպl��tv����pRh��Ne����o\Ku-���r��q��X���(��` ����b��ۦ�7����y=%��ZƖc1��*G�6g.-���Y�,�m�7��y�3�`[D�AHL�3���&������w7V{����iL	4����Uв*�)��}���r^�gC�F>�U�*!*\V�X, ��a����='�,�Mw`��f�F���="#��%�7��<< ���}��dS~x2��n���]�@��rc�싚��KB���]�N�hFT'�����qj��2��I�$Y�L����$f٭p��EHQR"���_����������2�uq/�J���"�/)����p�Â��a�f�;��b�]#T{���b�)+��pf��}D2���~��W���W�h�w���̿���������߿e,��û0n���P�C�m�����k�Coמ����㿑@w?f�f��=��O��5�����PI��0�*�**$5c�{�*n^92�gJ��f3��!�-iw:ܭ�f�l�q�M)a�J6c.ؤ(�D:��o;�_8]{޾j]�����<�AP�e��fs��w}����ICK�zh��=ɛdvuqk�&�"ӈ�c3��=�ݻ���t)j/y�I��L���������U�+�f.�eL�>��v��ҕ*QήX��v'*�^NA��PXjb���/���H�zT��2������k�U���S��q��%7�xx_��9u�;�ꪌ����\����$+[�BY�4/(�$f�w�g���	��t%�8l�K��O�`v��dT��.3&!�C��8�l��=#W���_�����r�m��]j*�8PI��*�{;f+�)��O&ſnZn&�����m�)g�(�%�`�1�g�{p���a$����z���A��Z�rdܽπ��J�BeC/cL"j�[{���݈�Y��(�d�@,s�%�c[I��P< J ;il�;�z��Fu���ykƖlЁ��#�E��+�/�]1 � b�] ���$�H���5A�ԉ"�h�hc�u��9�PN3�mt	RA�H���ĴS0J����L� 9ef�S0�b��?}�w����B��"qzD�q�Gh�m-��� �O�	c2�dk������V��E8C1 �@6ڑs���]3 9Vymt���@�y_7����i�] �׌f�@��k"�T�gk"Z#�Z�:���3p��h�"��Y�k��$�D�sHZ	"��%{d��V�����ϟ>g�&��ύxH��m�S0D���L�Av�[Z0"%��-/e��D
���f�H6�foq[EKba��O£(�̓i¨�ꪚj+��LP�eBԨ=;�!!���m�;;l^���a�t��E��-�@*Q���D�J����L��n�]�/���y��oV�%F�������u���v�m�}uw�˺�݋/R�c���+�!�1q�U�ב��w�D��F� ^G[cM�hi�ʄ�� z�#8�A���0�A�-��*$�0R�F2
� N!�$^cՉ@k3f��5��[��aV�l%Z$!��� ��D��J��G�����2�(�
5�r����� �[~WSX9��Fk�.�B�L�L�',m���.��
�,��@� @o�����Z��� �_^6���,!Ÿ�m�}�p���Z��<χ��	QM��Z҆��㍮�"��%�,mF� �R��h&��H���p&"�@3,A7��-�p i ԂH�bu�7�f�m-dL��54��������X��ec�>f�3^��nP͜���� �<?{�@+Kq��� �Q@8���� �x3�v�4$���,�f#+�~_x��E����Z	�)KB��p�ۿnl���Es:���x��i����J���+��f�>�7Q����W�z�f�u�������jJ��lC���3[l�`�9LЮ�1U�Ř���K��i�*Kհ��)d�pDt�J+(�����kڵ�it|����0�
�K���:16�z�:��ng��v��y9�Q�S!��n�Ҏ��:z��VTN�@�Nͫ��s��=� ~Y��^T�����徭mF0z;��h~�u'��Jy �W`��S؍ ���bE��Zf�V3�ݼ�Έ=z�9=ay��f��]������?S�{��
/�wNevV��6-�P�e�0�ngp�ܯ�Wt�
�(c£�q߼y|;�V�Nd��Mp��qM�(B����d�=� ����}�kVNs�Q�X�8�����X�Ҧ�e-��:/j���:�dc�ي��A@�0� ����g�"J!�r{)N����VP�뿀�F|���	�z��y��(eۭ��ݠ�J�hZʊQ!8�iڢ+)BZ���;����u�f�D!e��[;�%�ϙ���-��p�o*G�B�5n#C���p�뻻v=Q��z9˪��*���Of�+=��{���,S۔�U����Η�B
R_|��˩T̤�X��?6�M��I�ٽċUwt��==�.�+��̨]ΪO�鑯���+��+ifݛ��}�WϷ�������E)p�9�	cg�QLқ�
flCpa�Nwh�ݚ��I�+A�K���FȊ�+
�t���J.�\O'�����v�����\�}�W��[3����C	0�8b���G<R[���:b`�C.c/N1=/D�L&8�uT�!nu3-ۺ(��u��0:-K�Z�W�1�Ri"�q˰��t�9u�*�����>�V;]蛵f۷���Q``Sr���v� �2�4���ǚ���Ӹ%�Gv ��V�(l�{��]����q���eg���4e�tu(85*�۷c�5`�j�[���1�k\��0��;Xݬ��P���	����A�@�yz=τ�B!a�8G�,TR �"�$ �c!))P�^yXp Na'0	12�����e��ZJ�1`�w�۴)�W!�3XԺ�t�v��Q��Y�Ws5�4��6��V��U�f�]�.t`�pk�K.v�1GDmԺĦ��T�l�c�.m4��D�fmqf%�mR���F�2�K���ح2i��Z��ޱ� 8B�X�!��4�&	����<�Ֆ��G���)�d m��a�X�f��05��5e���`��Q����Ism������`�S�_!Y  �:��)c��cl��wt/�Ĳ�&[]5�u��=��K������a{V�Dơ-� A�lf���j-�Xb�pa��o�~��Ҵ�z�hT�wִT�:�x��@-À�{�Q*�n*��N��W��d�Ƅ�pS�L��=�O܊��s��ͱ=��@���+X���� 
��3I5�\�$h��/˿F.Ժ�����R�(R�ޝ��d8P�D&6s/�x]*�;�y0���ݚ7	�����b'Q���ڎ�
	\��B��{��Oے2I��uQCﾽ���f�Vhi�$Æ�O^����*��������7c�{�}P`�Q���B�k�'�آ��[�F����_��&;NO�0�Y
[pb�}�w�a��T,��gpK��,�.OgM��ⷝ�{�u�דWi^�DԾ[��$�>vAj]�]��{���e��ūK�T��-*8G$u���l���3c�֪Ki�ƏUDVR�hW(7=���$w4�z���h"�s�)���1���װ݌6E��Xz���ۛ�Pf��GEc�
K��w:��JK��.>f4�)�+cq�N��+2����ϼ��7�}b�����·[.�]�#c:��{r�R�ͅ,�6bmCK����������\"���3=(���H��Dj�/vޱ7:�����퍫ۓ�!��OGʨ�G6*��i@A'CM8���p�L&�k���k]I���=�B̗'WU���F��2{���9sj����:�>�O�1'c3\��CI��M�Q��w,��ٮ1U�>�5��V3v�5/Ř�՝�-�G1�Z>|�k� n�]�7Y~V�~w�NM���&0���ۦ^���ﯽa\���X6���ir�A6�Ű���n4�u�]U�Ԟ�l�5V��VX���hʅ	;����͘,	o�3I27���ucbK�d��|�Qsх�"�
��봮�!���֋ �+	K3��,G#�	����%jy�\����Ó���\�I��\��_V�����x�Ps���'9��vkl���۬�������x��{�N����L�*�Y�6$YU���h��p<����nS2ҌQ�LDh�c�d����s��1��WƵt����56�;$�yo�o&�p����4�xT��� ��niF�YI���w�#�o=���ۺdkH	N����L[�L�,QV��ܟ*�)��}j�p�]`���I"������}n&b�%�9)HZ^/k)��׉IUP�lUx�d�ه�uN��Q@��i�I 1d�m+���L����$��
��[T#� G�b?��o~wޛQU7u/�2z>�5Y"�X�#!��L�0�Qչ�9ג���bKk�[]9%��&c������V��|��8�.v�`�.'�~��iO~g��Z��FfY�D��Gջ���>e�DF�\��!�נ�;���S��q���tT�\�����^��;�3URh��=嶟���^��5���Ζ֑�R٦�B�[CD�.t1l�����7�%�K%Q�k�"��,�;	bb��|����m�ݻ]�u�5cT߯�Ȫ"���,�Z�rS�%�x+���g��n�K���s;����#�srNM�;ne�e���6����}�|�(䠓�E�?���'�rO�(�\�[{���ܨe����3��f���q�*��1)�j	�k���k9�E:�a�]:�>�|#"�f���o����X��N�f�ʲEa�.���b�YOWu�B�܉��]ه!��g�J�b,U�"��hZ3��B�9�Qۢ#o��F����p!T�F�A�4Y�l4�_W���t��RM=}w*/2�8���`��ඎ�]�6�W�-#R�|�

�YCv�2!C�:��~6�{����LnFz譳�*��VȥuۍK��%��	L�X�ٖ�W����85���i�h5�!��wgvgި�@��έU����􌉢�'=�NͰf��R���2eu*��i�m��M������4��y��ch�﯎�&��f\�x��=px��������zl�"��͔�ejz�����&í.�$��Xb:���Gj�)�K0娰���
����\$�\������{O�T�ṥ,���>��U�e6�f� ]dj!��)�h���x��8e���3d�:h�ʮܙ���r�8��B�āMR��.w����w�q�N?;�������s��N�'}G�tT�*W ����`��FE�k�集C,��'�]����bGE��sm��bw �j@���^���}���j�<us�ݽ���`Gh3oRUvV'�5yQd�O9ۘ���^����/�q�gc�9���㨍�U��4��UQ��b��%�%�0�ܡ��d6��_%#o+y��ٰ���/��\U���y�y��|䒡��ն����,)rȐ���V����D,]P:�y=�HQ"�	�H�p�'RB�(H@H�jR0�0Mm�Z��(�ZJ��z��-RJ$ *Eb"a6�HX�kF#�*[j� J@����I����v�t-��2�b���kNf�Q6&ڳ!lsm�*�ѭ4��qs]oi��XYW62�S4��fvQ�J���:#p3\���mIt�3��23P����S�c5�^��h[����.���В�)0�M�f��i�n�	h�sjQ��-͆���љ�k�;(�;\��Ҵ����olG�,��hQ;!s���w;R�Ff�K��)@� P���0b�n�Yf��)�ҵ�ѡJ�Zݦ��e�m6�bZ3Mi��v��Z������R�..��L��߾y�΢�E��}�l�ϑ��F����Q͵�O҇�-��׵D�m��`Ď�����2���/Y�r��:e�|�vJ�Ss�}�}�M5�O>�eŘ\�������GF�{n�N]Ø1o�g)B��f!6�j7�4o�f^���r�ڎx-�f{w�S��?R���`q�����۝�{/�?{��आ��{��}���V1B�9��A|�a�މ^�PS=IK��c��v� V��y��Pl��
�ַ-���Ln�d���}���ӽ\�����]����a�4Jf:�ߏ��#[��+ב�]>�X[x�292���H��@ʇ,�s�oS��t�-�z`��}@���=�f���YE��U�a�k�w�jLM;Fgh�v4�X�e��[\�K��.j!]��|��j;2�#�����-�>�N%��y�hj�u9yh�vh�$LH�Eal8)���I���υ:[s�j�kF�qfczjd�v�v�W����#�?}[�"歊4~�:�B�&}��&E��	�`=Cv��#��i����6�(��Ξ͋�ܡK�/����%��i9��  ��Q�yCYqd��G쟰m^�!3 �'sL8L��!6�7�MD�����Y���xz�ݐd&����l(Wn�]�n�Ϗ��b�����OWע8�����L�6І����݆ԑ;]l���˵�e(�ܡ�:����NjT�o�V�ݶ`ۀ�*�0=��/�|< ��1sP�yA-͋E�kW9�R2�K6��;4�nG]��cU�Xk����X[)���;�|㛘{}w�M�Cw+M�%*�kA0�Y������4R(�	�墌Ķ�B�`v#$�Q�So2������f��,�M�:��q�9�1��S̼�E�Yb�0�^e\�hHm�B��lb�AG�٥�b����vw{��5��R��3{vB�k�=԰W���oǺ�~����4"���A�R��˝u��v���<�=;o������6q�P�,}�6o��c�=ǂ��CF���F�[{	ul�+��f��*�B���i��%^��\��O#��!1�,]h��A���+�����[�q��6M��֥z�EQ#�+���E�Q�ԛ2�sjKт$JIRJ U��XIH$"([)
%:��q NN&KJޠ�9�tK���B 6�����g��+��פRj*������*��O2�Al��!����{�DY�#�T�\�&(>1��ٮ��Ε>�T5�&�=����{&W^�r�A���/)a�.�6T�P��!&�6����pF�y���Pj�>oN�;��zӝ��7�C��C"n7�c �z�!�^��� ��wd
SZʙׇZ\l]���o���ذ�����V�%.-6�%F��m͕R02���S)H��-�")/}�;�)���7����R��}ֽzR�GK���||S�!�Iղ~^�K00�T���r�H()G;��W��2IN��s�P�̬r���L̵���=pD%G0ն2yh����e��j�T	Ә�i뗔@H�癘�E�hᄧ7{:NPm�EYqGN�	�����}�U�5�tT�+�6|F�1֣�`� d�=~��l5�h��Wg$����+�PV���hT[���Lmud��}ū
TgvXŜ�<������=�g]�X��|���U<�T�1[h[�P�$_�M8���ᦝ��t��3��+���}��2F�P�5�C��@�0��m_]݅[	Okv�F��m�C���9��v�;o�Wi*��p���­h�]cmmV�`a����`h�36:�6�kc���m�������ښ���vaX%�>/!q-��9t�*g�϶�+pR̾b�و)8n������Vj�O��,�S�Q��V�11}�wn�x� o��zP`��q�{� �P��d�	���ʇ	 �M.�����;�bV��oD�\�I"��v��;�W	�E� �C �h�y�r��4TR��\�2hQ�K"�0�jj!�����,�[�&z�K�2I�=��@p�0-	�ێ��z-oY���=,|l��2��g	K2���"�ړ��ܦRPiÈ)����L֖k;�Y��c��'�W���IY��������2J��O������i�&�.!�)��,���
+������j���'��0�I"(��ڥ�+3�cd=�K�Y�/BYf`����`y�zE.�2\�D��b�qD����)�G�����ACg�-�E��������\�]w\�^$sk�$��Z��/�X������{�R:�{�Kb�`�	X��f�T��x�F,%��[��J�bU薂�pLy�t�B �qFgi��b��`1�a$ebD~���'T���MH� ������&�m%Ѷ�v�jW��ɵ5ى��֌�]�������5r۠k��q�MSXic�.p�.���f��X�F�r��f�u6��ڗ0n��汚We���%��;K���j��3�t�Vvu٪��"�f7e�%��F^i��jW��PRi��j84����nv�3�����n�������� ��@��Tk�H��b��]��`�]��*�Z,�"���RD�ԫ��.�Q�U
P�(�mAd�;���oZܱ<V󜬶1nJ��������
5B&�O.�u�Q3n��!��nmF�gp;�{1�����p��
;�U��^xQZ�tߟ��ׂ�Ɨވ��I����^k��\6�]�m	H�s����_�\xh�u��^��9wM�9YZ��x���B���8δ��vyu,Vq�6�s��ۛK��$�����,X"1���%��?o{�-7�؛��6���޴�.�N[�S�ƃ�X{��z���5��S$��!f�����i��vX����@X�q�%��S*�3'b�"�ȱ	��C��[Y�K� �j�q�,/mE��`@�[���Y��݌�NB6��s�i�^�ۡǶU9BWj�����d=�`�Y�I6TU��0���/3�zg��y�b�e�(�*%�LDH�plz�3y��p�4��kZL�W|�6D**�*�R�(@`9,�9�9����V��(LV.۳�mw�}��I�%0^�cM*�yS�k#*z��w=@�!�:���,��@���NH�����ebj�9g,� 0S�$����Mg_ua�05x�(�	�F��=�*#\hI�yr��yQ�0h�d9���=Yí��-�R�M��mM�r�"�N:~��,���� �H;�l�C��r��G.d�DL�����`������9�ݏmf�E�Om�`�B`{���V`�C97�وO��c�2�~�KR����0��t�ud��d� ϙ�(��{oǎt��<�2.�l�&\��9o��n&s��4]볖X-؞�[���t���) ��ھ��p�"%�0Ӎ��ϣ�X��Q��"�:��ӌQ���4���.�
o-�Vr��2�͑���Ѱ-�s�y$~Y<��rT���]��x�{���r���k�h(9�nO,ØA�;��;�>���`����V[|�o�ܮ�"�0�kz{�T���VC	��5�eCG�0���X����Yq�e����T�z�]Sb��K.��nj؆0����9��+��0 ����.B>���J�B R�Q��E��D���b�Ɩ�\�i�Z��8*�����P��}��!LB�|tҠ˾q�b�����y�c��N��KN"X�+b�Pz�'1>���<�n��lP����u]����S`R  b����E��iG����`x�u4H�lOZ)���p��Y� ˗y�2C�b��=����E�2��vf�R!�O0ElQb�Q� Qn�ؽ�X.�pU����;L�P�����c9�=�����ҩ��\����.�i��<D��ea�YdބwBM�b�u���把���8����Cis�Y4��'��0���VFAF�W,�v6�.�sq���Nj�1�8�n����J�h�dKFM�;�mj͔.�E��8���F���{��DZ��C(�p)��f�y�DXÙl�Ѕ{B��h�Њ
��e֒�p��(��ex"f���pR	$$:RZH@$b!���A�Փ����P �����2�G��)A�G]:W�����p4��tAA��m��Q�y�	�ty�6�3%oNU���0�R�^�"��Y�e-R$8��#������2	0����Z�f��p����[RٹQ�6�C'e�>��h���M��j��A���9�� �s��D��(A"iS��n��K�%���(iH��E�/erK9ӘdB�=���`I@��,T[�(i"��a*�3���m�gw�,��Ж�~9%�D�X���z�-3Y�:�\��0�k����˶�P��-	N�q0����-�µ�J�Aھ�
���>��̢3)�Y �a�,˅"�4X�Ƿ��:�">�Q]��6��Q�(]I�(PP��nS�$�P���s3K��������H�/�� ��ı��V9�O�>4�����xb��A=��ݒ0<&)��$݉�����Ty������D.<�>qli[�a�?D&
L�ok�j|�1X�Q�fwia�AP�u��pp��TI�A�y��虓M���\[�%D������UnPU��@���Œ��Y��1H�"���V)r�P�-���oU�ĝ"	�{��I��+eQ�{�*��SL�p��~۳��PŶ�g�9�0[�-���P�%�^a]u�Q�^����h�*����}��xc�umxV��^�޿XPd(�/��dM���kZ�ț~���շk��������k�Ԧw���2��TF���>X�g6�[Jz��1SI��l�X�HO;T����WIʞI��g�9����O�^��`�l�1��Ջ�p�D%r�Nغo<������j�@�u�u���a21��36����%�L��m�lN4L�`�%��p$����tK�g ���&ZT!�ʢ۷�,�Ϩ���>��l�2Y�4�}�?b��v<@�$��s��<�F��zb�^�t�Dtmy���\Fʹ��ߩ�ic�*j[�h�s�\Pbe��gk��x��}���ӭ���P�Z���r-��C�^��9Q#p�H�7w��|��y�1�����;=)��圂EM��gw}�d�9��mw�:���F
���n��C9g$�@OH����}i���-�0�	d��U�zPm�(&TVns�td���I(T@��ܬ:/K������,̌(�@;�H���i:���:�,���'�z|������+����@}ê���6}duZ��l�.!"�����NP�7e�P��X�]	Y�C�f{^'��V��*���9$^����'�:��\þ�ݴ�B�B�\�p4�=ǰ�=A��$�m*I$�OrU(�iG�� ��ܔ� ��}�&����)���u56}Ϗ+�J�S��/��ڬ@�S[��A�z�L@��ʞQ����-oA�:�Z (�� ��:�i�:f�����N��^7~�l�ۡ,v�m�9�5�����e����!�@��,n]���k���?�o�>[r���ϼ��TQ�8Q��j2%-�A��M<����?�� ���r�ϕ��l�SȻ���@�w��A��ƿ{>oDd����#`K�� a�h��6�7I�}�^�Z��4
�M��o��y@�y�39��g�1V� ���A�^oM�]z`����""�l�TD� ���I��E��:�-Zޯ��C��s�>��y8k�ǒto�vr}����xS��9��8M�}���>/��F��������pF�A���ze��|��;��������8uc�Y�h
u��W�w��7��$�t[�����{yےF>�q�u:�z��f{}�q����WL廛�o�����
�g�AD�� �3O�'�)zXt�7�|\��
����A�`괒��6']��9�(0�r�����O�ŷ�&-R�Il�B��d1�=aD�M�/sL�(?C��wt1�{7�<�
 �>G���o�Ph�c�rÃ~� >��`>�����-)�C�'C�|�z$O�|=�Z[����4�?�H
 ��'��Γ����)_g�2�� �/��K2�����6�����Ԝ�����f鋦�p-����-�}x�p����/�6#��{$��~flj�t/��󸂈>�㴸m�{{R[�w�a2CרQ��} ��C��*5��vd�h-�./���EE���:�{'��|N�^��j� �aޝi�,��C��f\��o+>6��'2�}
ÎH�����w$S�		$
J�