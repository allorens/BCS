BZh91AY&SY�w`G��߀`q���#� ����bC��           tUJU��B����)T�DUE) ��T�(��P
�@� ��"AUTP��� )T�Q)**JQz4
T���4���(�R��IH��)QQPT��J@�UD���UP���
�$!)UP*��(V�����%UR, f�U
�`h!BUDw .�(�Q*"�k%QT��l�1!TP*�UM��I%"��B�B�z�P�J��Ҕ:A��֟ P�Gpr G4�QiX���;�G�
;�Ք�@�1�J��w�on��� Y�%TTJE!T�E/���l ��ʕDS��l�J���n�T�*J�_{׬�R����QTR��Y��R������T��}�J��Kޗ���([��ג�)*����$���AJ�7�JH ;_)RR��[��^�U�eއ�j�U/k��WmT*<9y��J�w���*�������R�<��סQt4�^�ԪP�������U*�=%�
UTR��>}$� ;���JS֥g��sݴ�T�J�^UH�Tw���^�z���{)TUU��w�C�����
����=T���U��R�Cr�r��P�ؐ)J�T�-���IS��ʔ <�ʪk-�n���Rs�]�*�T�F�QT��7K�����gNr�R���u*Qn�E(�K�Xꔅ
����*Q*��!�
��!P�Y��J@wִ�m�7�wSf�U��:��kJ�93�P*�w܄�U!`ƩSmJWv���T(RJ�����nے�����P�ʑP�PHU��w�J�����@$R�7@su@�m5�
�Q�s��������9�(�,�r��@��UE"*.���@<wk� Uf�� ;�ܠ;`��  �gq Pq�`l�K p�:;`���cAE�UT��*P$�5U)H!��P ��g� )�X�wn u@u��r���ÊM�N: �w� �c@��� ��Pg�QR"*'YI)QM���J��_@�w ΓuU(w;�lܘ 8�EQF�9� h�.� S�Wr� w:.P_>  *� �@ S �JT�a2`#C #�"yJJJ�C�4�!�b11�<RUHm      ��jz�J� h     ��)���0M0	��2h`�#L�D��I#LI���i�'�d�����O�����f�F]����Rb[�מKyK��y;�|��;�9��@^�؀ *� ��P� ��_� �
�q�$<?����Y��������*��A `�I'��� U�KЊ��������޿1?&��Mb�X����u��`�X���u��X���.�u�kXk1u��]`��5��]b� �.�X����`��u��1��C&�`�5�k�\X�5�k�)�X&�u�b��5�k�!�X��cb�5�k�5�k�$`��	�SX&�b��1u�k�	�CX��a�M`��5���.�#X&�`��!�CX�q���]b�5��]`�5���!�X��5�k ��]`��.�X��5�k �.�b� ��]c�`�5��CX��1��q�k0��X��b���Y�X�5�k ��X��5��CX�u�k��]b�`��5�k��X8�X1u�k�	�X��X1�kX�`������u��X��u��X��1M`���u��b�X�0`�X�u�k �$f�`��.�:�5�kc����]`�X�����$b� �&�u��X�0u��Mb�X:��.�u��]c�u��SX��5�kX��5����b�X��u��]b�0�!�X:���u�kX��b�5�k ��bkX�15��MbkX���&�5��bkX���5��bkX���&�u��`k���u��M`�X:���u��u�bkX:����`�X:��.�u��q��.0u�k �.�u��b� �k1u��]b����]`� ���]`� ��b���k�.�u�k�)�]`��3X1b��!�X���b�5���5��:�q�k�	�F�X��]��q��1�k�)�X�f�M`:�u��5��X�b��5�k05�k�)�SX�Ma&�X����u�kY�b���]b�cX�]`�k1A� �U���X��WX��]`��bc]`�cX(�@�
��E5�.�D�(� ��E� ��5���D5���Uu��0X��WX��P���5�!�Uu��P`���b k X��T���T5�!�b.�D�D` kX �X�`#�Qu���A��u�.1A�":�X�`+�Pu����*:�X� 5��1U�"��X"� ]` k ]b+�u���1X�]b+�Au�.�� ��(��WX*�` k X�k�u���Pb kSX*�@���WX.�U�Uu�!� ` k]bk]`�k`��D1���`�kX��WX��� ���`�X����X���.�u�bk �.�u��X���8��.1`�5��X:��1��M`��.�u��]bkX��5�!0u��X�b�5��X���&3X8���u��b�X���.�u��]a�X�u��`�X���c�]`�5�kX:����$b���]b�X���5�k ��b�X:��.�u���1��X��5�kX����u��1��q��`kc����5��M`�Y���.�5��M`�X:��&�u�1�.15��`�X:��&���L�}w�c g���<��3���y�a�Iٙ�&����JQ��,̭�+b/(L��&V�6&�i�E4B�d�����u�!dJ�!y.l�-*.����<:e��KF�-QG,��y�3n�U@Ŋ��J��V�[Cu�+h��0X�Y%�pֽ�
�l�3pm�8(/2bݨ���fPi�r�5�R*��S����^���\ש�^�47U��Dt���U*�^^IA�E] n�mq:�[��H����q���VI��]Y���.�ڂ����oZO�7<��Ȱf�UNK��+t'�m�7X!���-T�.���.[��Q2��^^�Q#UD����4��M��4 du��wKi�7/������kT#L���lPU��T�F�ǎ@@-�"�JTւ:T��F�0v����y����x%�YoR�G�;�(�V0V�0ժt*Ґt�Ov/)ZX��6e3��,�C~p孔��c�5h��@��$*���^��ٲ�j,�%�ƕn�X��]Y����j�5�R�>++mq�U�(�l�{m��j��sTyͲs��Q�u-�V��������Q�I�٭�M7��K4�3<
�p�/tbZ�����oM��i�F%'t�;�KV������*��UJmG�(IV㛻X�	���LZ�D]D���wCH�.��{F��X��PA����oUɱ�xM��)�YkXͦM"���/s �A�7����
�Y";MdF��ջ��jT��ܘ�1w"�黺yP�l�L�U �\z �ɒ*���C/����Z�t�����M[�D)n�\l3V�M�ST�B�z�<k4֊ ;-��v��mܼ��y-y�޼�Uj����Z��//b�������P�����\�c��R�Ygm��fJ��4��:@�g0@ۊ�ą�"�;h���r�bl-%�7s+kr�Z��$F6*�F�32���3T�M�y��D���7R�P�vrMr�2�%���և 8SM���>�����Î�GOZ��V-����sh.�4��˛�Wn֌J�(*52�2��"a�g!o/v��eU���B�P����v�@kZ^�#2�ۣus`��]Q��j4bYi���*!dF-<(���%u���Lb�Q��7̎�.�Mu`ưL�Kպ"LQ��ͺ�aF��y)͸��i<��ބ��N��suѨ�@iu�W�����M-�n�OKK${�"W�;���fQ��&�96T�j+�a��Mm
�h\�wL�╚o-n1aei#jf7�z�n�����&Z̧t���n����^�e�OMխ�S{3���"����!�i*eLw�uNT�I�nedVv��^�O��'9�kL*��j-7����'� g2[�A�4K�ډ��́(�`�4:�cٚV���5lw���<8���b��g֌�lXĪ\�Ñ33nČ�HM���x_����K�x ���Kn\*�-�LTa!V]X��nK��u�-�ۑe�`dRGJ�Y�E�K��į/ ����d�5n��[J�t��L�Ŗ�����)m��I�B\̽��BT+���[J�U̹/2�z�p;q�e`B�]�n(}�2����e�ݬ�B0֑�n�2-�� �Rʖ���+1�a	�)j�c+v���9�ȣI�Xh����Im��Y$�s��Z�� 6��̚���L�PX�r���y�,�e�F*#��b�Wx�:�^8ߝ���6.e$�j�Vԁ躶�=�����2���s"�^չ��.CQ�ݡ�ᰴ��"�!4�ѽ2EP��ۤ��M���ujnQ� LSzK�U�G@;�r��١�4���)�6�;5^��45���qn���e�"W�Ӽq�dڦ�;*��`DP��I�%(��Qܹ���U;��Y�&hwZ��n11Ȫ)�Axʎ:ż�rG,�a�:�1�x�h�/e"�iӘ���RO�t2�*m�iѰ���[[/ ��m�WW�&�!b6�wk1i�r�K�P9���;sBwLTa��yA�4�� ��19
�F�ݢ4xԲ/ݧ��lSUw{)jD�А\�S��X4���%��ٕ)�ݪ[� w�dc�t.F܊�#6��WN�@��-�C���VGB��P�R��j0��6k�-����!a)�A�GHӼ��n�.�B��X��*E���;��; -���K,�,�z���wkh��F2��f[A#�n,����q�,�5/}���'��sUe�b9��\��|��m�+��)L!k�-��6P��I��؜�C4�'�m�%ԩ4�K@̹x��%�7^@�*
 d��(&N�usCsq��[-;y��ЇLW~*��vS�ɭX�Q��ضn���a���T�8d���:��h	�"֙Gwݱ�"MS�����{%Ҭ@�l��sB#n��(剬YVw$9&G1���c{2���49yq;�(���W�D^1��(&4��\��,WtFԱ���n��4�f	u�պ{f�����{pѹu�(���݅:[B����t��^E�=�˥n��o7@�Tѽ׎1g1⨡���� ���<���9F�w5T�ב+�4�����
��sX�ҥ:"�,�c��$�w��BD����$�6�J�Hb{.�$ŬjV�&A�j�m[B�T�d��2-�,v��j��GL1V�IL��Y)	\Y3&�t8ٻEny��͢���:T2b�sq�zU3L6�X�Ż��ژT��̰�����	z�8V�y	�N�(�
2l�k^V�1�ȱ1 6ιZ*�5��U=VD��jN��5��4�K�+{W�Txt�A<�={���%w�V=��J��Em���WJ*�7z�	�������a)2 �7V]��d�p�F8tنZ�E1V�CH�U�k��Q��We��Rd���B�ڹ� b¡��{NP-*���X��֫V���x��4Bz]��C�"Č��P��)�E-7��f[m=Ra�ecm�ؗM�YG&��຺�̀ ����ZIS1�fP{��������\̹x�m�X�!�M#V�Ub��w4�nG�[kr���.IG8�il�:AyFSS�-�J]�������Ǌ,ųn�(-��
�V����L�kp�!T\0��Y��\p�m^Q�;�hF��aX2F���cj[�(�1��Ӛv��6/^Ը���&� 64]T��BQ�BF"^���RQ7�m�EZ��V�$,�)D-�ͣ�ØU���QeV�M�1'������1f݉�8��4�Ft��x����&��C�J��A<6kRD�PtB�E�ܙ�����'rJ��f�/&�z��S��C�I��ۢ�x�hn\���ŕ&:�(���CO)n�yjJ,A�ݚ>�@�-;��9�n�7Z�C��Z�x��N�L֖�B�'��',ɳ�6&��5�(J'cۦ���ة�Y���bR׌'�(E7�wf��~�ʍ��Ƿu�6�D���f����Z�yɲ��;�]*IP�`�B� �xV�V	��S汵�����e%oe�,�EF^F��WI6�ܡ �R6v��6a"���
�������a�*��!(�ݴ��dK���.`�����P�f�@�n,-9��ù�5<�Ln�`�V���W1��ۦv�N��˽p5���uj4Bȱ;���m�3 T�`'�Zt�b�mK��,XDP���WB���U��@K�ZmT����Rm1��)Zb�@v=ױdG0C��7UJZ�tr�j�hTZ��9��=xF�{{i�@IX6'J�M�ǔ�[9��S�Q���f=4���$�(����+3ט��Z�����4ս�z�X� �J5v�oB�+r7	��v걨\gX�bݓwq�f	01RJSul��%	��mM�ou�+*�s&+&�t)41��;*]���(��@)��z�#���]�Q��ct�5�j#���a	f8pa��9yM��6�;�Ӭ���x���f�Ck*��.Syq�b��6J�ؙ��ݧhm��e;U�p˥qh���
�D䷊�k�����j��L�Ôr�<DV�խ0����
�!�yJ�Տk�n�׀L��nVԺm6-Y[��S��Gf d��qT�P�:�ed���B|ű��9�zwDYKqʲ���d�I��۩yv�͵tZ�D�$1z��l�ql�k	��B���2d�W-hՖYw�*<.RS�Ӳ�(f����\tCݤV�z�X٢�pX�f#)lǛaҽی���eZ������@�	#[��<
4��f�@c�0��.~�!m�12-2�����^B@%Emg��92�[Ӻ�S2��̻�3R�[5�jJ�m�d��Y3�3E`��M������f*	*ٺJ�(����T�o����ASԕٙN��)$��w�,�<�o%d���#��ژ��v76�b$����Xɂ+-�*jh�770H��2 ����3ܲ� 8��,c"D�II�@��d��o%��Y�zN˲2F�56w�S`v[x��r���lf�!��+i�����A:���%W[L�X�{GV750ဌ��h=��1��)	�D��II��uS��ɹSD܈q\�J�OI�
^�4��O͔��̹bb;t��e��䨥�ʺ�F`[hz��/q��n��o��Ʊ�5�-�wgv��l�)�G� ������-�h�Kb�W.�Q�T��LX��n7NЏ �5e�n(0c�m�o���RT���
�/c{�+k�޺;��M��^'����Y&nPF@��Un������o���qe����KK&�;�%��w�[����L�N�O*L(�z� o30�$�s"�չ�-
�x�Aiv�&ݰ���%��ܐ�VVT�Ѱ2�@ժ�to"b��jVG�Ưi2{d:[q��@�]�� C��b��ҫ�����cyp�r:�J��5��-wG�X���Z�d�j���7O#���j��.kW��y�馒 j�D�q- %h�<58�U�G
�j��Sn޽�"�] t!�/o.��N�M���ㄩV;8*�h¼�M�偗�"�zK�́&j%�ک%`�^Փ/*k��M$�(���mтm��ܡ�KI�m8��8��	�[��Oa&%]��[4�![�6յ��d/�kq����� ����UtK�n�6��y���3&q#:M�<�!�\ʸ��3�a�{3�hE�hI��ǖmK���n7(a��<ؘ���J{�Yz��Uskf1N��3pH1&pKR�)�`s[6�t]�`�
mh�����R�l5�.�A�t un3�a�t�^��Cv��Z
KM�X�9�n�H�I�m�Sҝ��d�;a�t��v"7jeb�J[�\��´b�@���B�H5��\L�k.-�t,L2�ʻء�Ɯ/�#{*�ô���K��k�Iv�ՇQU�N�l��╶��<
﫧a��K����݂K�AZ˙u�N�*�=�1K��k#Z��%j!�@ċWIzK�8	/-9�U��r
,:ԕ]�Z�ȫl��ٹy�a�n64�a���A������l�(�k,���BZ΢�juw6���n۠�<ݬ9�K3��sP�m��f�n�m�s���$S��:;�z�`r��C�ص�N���be���mZbH��4ӇLbV���vģB�/T[�-����V2�P���-@^�.�޼�,e�(�@%wwI�c��Qd5�^�A3\�;W.��5[.`��OD�A�f���/C�O�*s7%� �,ծָ�9Lݠ��L�wZ�!:��L�[<�ڍI�e��/\ ���ZU�0�4�!�m�cH�-�c��풉0�k��^��2�R��Y��*rs%k�
0�b�[<�Y<{��+�ڴk]<Ǖ��2�2�<;ǎ<�Ї�j�m��2B�D�#�k \���z�{��ݐľwCt)���70�f��2�:J��'Z9@aT4�gl��\������$���
1���-��j�8��d���K�l��s�eP��Yy9f��.w�$<K���V�Ʊ���T�q���,嚂�EV>��B*pܜ'dˆqA�d�+���&��cu����J�����t+X%�����$�5F����l�5ba(�&b��0�ee��t��ZͿ`���yU�&��1���zoMX4(@Y��B2at+�S�o���
�tX������ևAYd�\��X(,��V�[�v�C��W�N�;�AYkf�;��6��"'f�o}�i�9�0��J VΦ:��t��剝a�$�rq`��l�'h����L�,
b��Cn��*ěv�&ɖy�c�6cH�vvؗX���6�g0�u�[�T�����,7����Fi�S;A�љ�*��%�*�KJ����6�Ag��OT	��
`C��hʈ���I]�q�
�v�ι����Pm�U��+G� ��F^D��I��]+�t#u��DI�d��t�g!���D��$�7�_:�CHQ �C��L5�V.�d�T{�c:~�ʺ\p=)4]��	�-f��v�)��J۽��a�4�F��h�*�j�3��j�Q+����һoY�-�	r���� ���S9��I�˭�4��ڑ�8c`]|�����u������ ��Y����p��9���C	�i�X-F�#��xJ<�����\��<�1	�q�B��	d�PE�C7.,9e^ZusB��8�$È��>u�3#�e�]�0ve$�`����ˠ�ɲt�=�镏]�=��ku璚6�����{0Q�!<KǄ�*�CO83/E�����i�R�[D4C�L*a�s�CD���¬�.��Gג����ggG&%ų@2wC+�*!�����wY�{#�{��,�7�� �/��������ߢk�~o�f�Ӻg3Y�owM�{dY�t�R��<F�;����7s�=��BT��n뱐�X�fE��.�w��s�D�l�}�'y�9	K���4��v���ܭ��I����O��@ѳ�ۍf��/%�f��j11��O����㱂�+�뻳�p�8%u��k���\�32��rc��C���آ9�t�8�6ڨ͚i�X�Kw)�  .�V�m_r6��uy�+w��'[޾���֤�ƹ��u�pb4��R��Y㵽Z��Z���Ҁm�
�6gr�
ll�u��,��F�,�=L�{ak��L��{��GE�ǯX�7��Y��R�imt��.�;�F+N��ۄAQ�k�0��v�(kdS�YTWr��ޢ�i�F�Y��p��e��+�.df��U�'!�h�o��j"؄�@2l|lP��k1Ø'6��s2����/v�(����T7���)�1���ml�]y���)FAظq_6�p�������<D����aְ�QKYu�6
�\�Q+�w�uNv�{^S�-Pu�/Z�K�H͓P���^�9e=1ڶ�w\MSܭ�I��P֙��po����;[a�X䟈���H,�ƺ0��b��b�Tzԋ����=�MW�QF�p!��ȵWr5:��{�j�[�X,��@���ηENU��e�J*��%	���O�{��Al��ڮ�RW���R�
��X��l7Z�7k2w$�Ǉv=g%�g3;�N�9G�ps�)��������v�`� �sU�\�ɾ����YY�P.��!/7�V�]�H4Vwd��Ԝ��Y��}��ZC���o�7]k�N�uLu�T��'+z�oc��Jby8^��`fJW�Lr��x�rz�ow*S�XY��w9{n4x���Q��aژ��Ar�B��;gfx`�3�G%0z�C�eCO��ǳ�&])sZ����r��9o[�&4�M�`��V7��"���3TU��.�l�Lǅ�}�2Ⱦ3��*�Y_J�*Nh������.��ۛ�l�t��`�M��fݺ=H�ʊB�۪���TJ�[d� �ɫ��J��*�����c�OBg/��m6#9��ĚyX�Ӯt��X�`�M�}7���I�;wՅ*,!e��`EZ�:b)ևG�xZ�Ĳ��>E��RR��rW�.���:3J4�Sf�c�L5\,sK�:��|y�2/s3t,k�T���ӱ^,�je�kX�	c����Y�U���G]��r4T5kd쮊�Nhi��J�[�yYu1����ޢ�7���w`Na���݈G6!w]��z�X�Ԡ2�gmN�eF3���p6/+jR�(Aj�^q{5���h���ITN���݇`9���]r�p���ӢD�Y-���s��g����;%N�	GyG���s�%���]<I�X̓�"�;]���to��r�fZ�Uk�v��.z���G ; )���� [�<��:��	*��>�W%�Ul�n �)�V��]�U�F9���D����(25�+o���=���o]A��<��wY2�񫡬�Ƨl���o���lG^�b�b]���yf�҆���Y2�M���Cn5�]�ev��)�zՄF^#bV����s����"�E\���Ѭ�_43��hǫo& ^e>:os*��~[J��̺d���V���m�S�F��v�omf�%Z�6����%�����b�vPz�ԗs
ɩXb���>��F���]ظ��Λ�HR�d�y�3(s�Xc�y�Z�
�t���nf����N��k%�-��s��U,!ەWZ�mf�-�,۾͠��-�t:؜�P�x��wApǪdK�ժ�3sp�: ��Yfݱ[�� ���«5{��ڱ|���l��N�h"��Wy��|�j��=��\2B���qu*�ө[99�\�m㠥qam��M����x���	�n�/�ֹ6h�mG�KgU�h3u�z�|OfJ��A��31S��u�Ў��R�#6\�w�
vr�y�4�7�^�S���]<8��Ĕ҄��b���y�o�ob�om}n��F|S�z�n%���abKt#Y��� V`J�':�5o�TC
����l�w�KH��p�DG��í��ق	k�2ys��L�)`�&(s�U�NO�e�S�Y��\!nN�"ͽq�TX[��`R��jwT���o���s��ɔ��Kʾ�uˬc.�W���ZL���cQLB�tr�����j���Y�}�t?}o��bh����gCvBKu�����o�vV�)���Y+��w@k��̸l0���ɴ��Lu)�փާ���b���ck�{�:�!�c�I�sOt��}��qQ�2��k���]"7H��q�¶F��K�2�s{����3aZ���#t9W�{-��Qqq�֯`����(�V�{��[�1w9dSv:Y�E.f��[�W�|0�x�}xyU�C�n���ws�m��X6�f���F���mM���}�]!u1�.���˼w��,��LY.�Y	SV4n�ȡ�f	�AN�;S+��l2�.�u�e�=���H91.���x]�C�Y��ӣ�rY�=���(Jػ���N�ы���6��;�[��
ô�l<��+_�Y��΃����.�+���e�>�c����%t��4�őƚ�7�3��͜e�sr�G6
f�n�dΣ�����s
Ȭ���Q\$��,->�]vdF���ѢWC:�-�=qa���[}|	��{u�;�aVGZ�n�q�f�-ۚ�@��bq	S���on��ڠ��r�vܖ�tH�i�F��W*� ��&e7�Ԉ�2�%/h
���ۚW,�ŀct�[ �B༔����jD�鋬%p�,%��lwK��.j����n�t*=;:�R
3d�K*�ۨA��E;J�$�|�/:u�F�p��ɲ�3��c(N�7˭K}{�Bu��9�'�r.��y���aU�I|7���S��yH���JKsz>�������V�.m�zXz;�A���]8��_��]N��=�]�]��<�e�_*q��_l�d��/�[�a��X�������.�Vzv��7���ߝ�$��&s4^rR�n-�*�J|C��)H�]�����]�y�/�r�8�mSW��`����:�oGVyţ^+
Z#�/q[����}0�w�Ԝ�1Vp^բq�;���e���'���|�2��7u��)����)��kgme-/ʳ�Q@�V�W��sT�6>�h�/Vi��I��'7�y�8��ܬ�f���Xir#��+�uY�xF��c�s���Ӯ嶦q���ӎ�o	��R����]5.]�}�N�k��f��|�e&q���y���W΂�A].Y�:��l5r�Y���Ғ����;�.�k�߆H>���z3x,m�(�!���yǦ:����ې��M<�-��^xu��,���	���U-*�x��yJ7���'*�r��b�7J鍳yJ�|��|���.��D��k�dewl�|��6�J#�C��ڇ:��r��F͙$�q��s��r�ڑ��B(.��pg9X�*���1c˙AJS���H�`צ�5(ڭ���z>�ƪ\E�+��p���B<
�ڱY�ߎ���.֠���5��g O8vs{}}����Z��kr�5��Z���:�PU+�RP9��zje��=�r?��ۗ��ӏ2�eO� %�q��^�ܜ�G��l��]ƕ��8�M�b��|�w%
���+��j��V�}���5�(�nN��/`�Yo���uu,��oK�=��];��i��Ft��Ke�����W������G'�G.4g��6�	h��oo[�ת[�]��V��A��E�o:�
U7]a��.��ۧҙ�+��W\��jV���*�Vӏ��HnuL{�n_,�a�� ��>{�Ǌ�"���]u]�G����T�>�*���b��u�JS�\����]����������V��
�1�E�9�}�-�//��W%�{_A0���,�VV�Lr����\����L{���Ex��V�C�E�sr����_��w���|�:��1�۔�4���1��x�սR���"��Y��Y�T���_Tm�N�Z��Y�ChOz�]ֻ@o;�!�V�]'��u�4���[�j 	��9$�F���������4���w;תvP�����79 �4�e)˫z����mP�ї.�Q\�U�3�	ڷ��Ԡ�8h�me�����߭��I�e���_NU����v*�Uس+h�4e�}tKB�M&d�sud��뾺�.ٙw!L�c%-�a�6����"f�x�j��N���f,F��Z�{&��,�ź5�j�Uu��y�k\ld��=�o�j��M�\`��\�=�E��8�J��4T���V��3Z_�H�g�+��\M�yj1�ĝ�����7N�̈́T��'qaD3cS��:�~�C�2�m�9�u�H���w��M�ι�:],U�fm��}E#k� �Έ�vu.�Ρ�6����;4Ғ�d��a���Q�
�}���\B�gԄ�§΃��aޏNЊ����s�R�̼����>�|1MF���M�Z��]�F�6�-��K�̪r\���WN���C,�u���� �G�U�w��ݚ:ceL[����mf󾙏9�u���V�֩�̧���s��nr7���i�L:�}]��R�]ۣpX:��t��З��0��R��:[�8�U��K5)�U�K���ݝ�:�U�M�ih�e�,���:7XK&Ֆ����k�y�|�Æ�wf̥��:]�;xvM�mN��d���r�n�N8*�����>�84Y�r�����{�y��t�]��%�'r�O�ՙ���%�O�'N�^>sk0�����Eg/d�z�+���e�WX
YWY7�K�g���{�:r��l�X̷ϸ�z���ҒU���y�f�k̘ΎK�R��Q8_@��S�����u���N��XQ+�m��Ar�K)�F{���I� �yU�s��Չ�Ki�ÊllQ#�5��}�ӭ ޘ)�7:���_�y�<�IOd�.�a+�:B%���]��b������YsFuGy|6 ;��
]�d0�©�����]��3[�x�u"8�ōq V5q�T��ɷ���V
���{S��o�Fpc��^5��g*�B�*v*�
[�e�u���f�w ���L٬ƪ\Ib9d�3WjG�s��QT���u.�no&�׹|�z-5��i�]L��U؊�Wa5��Z9`νy*�x�ak}o�̙��W:��&R<�����>�ɓ{0)|3{Y���������+h���Wk�D0��ݮ��pu���}�i����d�D�����5� \�i�gm�"F_@��uoz��q�y/9�h�+w�Z�X�@;;v]Xp�Co�j}0N��K�7V��Գ2��t��L�R\/�x$76��*�v�Z�"���[1]�d����vL�L��2�juZ�!���x����4ي��[�5ݛw/_bNۂ,<���rp�A^����)Rڇ��g�����a�ӷ[K��,��]�p�	u҉/��:M�)w>��L*]���1�f�Lr�9I*�Gk�K��;���s��d�����ֲ,	�c����=V;FV��c
�l�))��}��V�К�]�ݳ�����)���4P��U���I�,`�=������:�FZ�	����w��z�N�tq��H�Nչ3%+�슾�i�*ͦ����fE3��Gt�J6�.�p)y���m�#igk�:��pZwh�kT�l�:�ꔷ:*A�N��v8%�yq��V�W�4	3�1N��>�c{�&��f�L������I$�A��s���>t��''Q|�Y<��������999ϫw$Rrs�5Z;2���
e��YsH��(�h���x�c@S
��/�0�9�[ˠ %�K�"Ac���0�E�J�W�,�v,��%���]Ւ<,$J!�{M9(#F�����$���)R�BCAT�
�HRʕ"�L&R-��\JpB������*>M�����l[I3:BjR�L�h��
�lT �����h�APf���X5o�4���u<��#�U�Xh���M��UD �
���4��:��!��,T�r�4��R��Mi=��2�[3M ϱ��
�Th-��d�(YM!c�����YH � ���/1:�1�4Ѵ�<j���&�W$6
�e�L�6ͻ6h*��E��!�\�8�(����,0�H�̳N�@��	H Ph�ƚ���e�I�)E(��Rc�^N4&QS^��ai�*�A0֐� �m�)����4A{��hYƱ�L��P��4�Eexєˣ��D�i��y�t�����&�2�C`##��R�n�0 ץ���i��|, �0L�vhc�m$�i� � 2���mi1L�e h
)tSTA�)�T �T��(�,ف$UQ 2йq�i(h�@h ��S-mK�Xu��¦�$�3E�(u�di�xCU �7B��WY��� ��D^
-�E���L%I�T|�Q�u@���%�g�n�)r��� ��o���� ��|u������?����D������U����'��?��g�Sy�v�a��A{kI&��V�s���Em�!X���VcǢ�%��[��+s���`����˿;�1��+��W�D�v���-K��%uֽF��ì��qzp��ml��b�kY�B�%wJ��z���O��'&����xu���-J�
"%.�U�]��ȴ�шs	4"��o�- �I��f���ʪ��*�u������a��Θ��Li�:j3h^Z���Y�p��ٯ��$_�L���j�g>\E)��:l�Q�������U4C��ld3�&�⬏:�=KE+�ߣ�+��\��j��v��)�6sw�)�mk�}�r���O���fW$i�0k&Mu3M]k���EJ���ޙ,�:v�Y�JTn^�,Q�n�v���ΦR�;<;�H<�����(8�+�J�1���L.&�������򲖎�j���()6Ha$��,�&f���9�N䤉]�S�6KN�P�f�̹�.��ԝ�jGwg�p��w��9�9���2��x�4���J��u`Ƹ�8����Q�p/ib����)q����>�K�-uPcFzVN�/�3t��Y|&c�X����ޮ�R;�;Rۣ�^^�p�����Zצ��kZֵ�kֵ�kZז��kZֵ��kֵ�kZ�5�kZ�ֵ�kZ�Z�ֵ�mzcZֵ�k�F��kZֵ�Zֵ�kZֵƵ�kZ�ֱ�kZֵ�cZֵֺ�k^�ֱ�mk�kZּ��k�Zֵ�-kZ�ֵ�kZ�ּ���<<��kZֵ�|hֵ�kZֵ�q�kZֽ�kZֵ�k�X�5�kZ׷�/3�w��l�b��U�=��ے�UU)���@�m��Z��c�m��F�j��к�%�x��]v]��w#x��ܧ���2�R�劋�l5���߳'�(G�b�=�]��<h�%W̵C+3Vc�'u*˗�� �|%ڣ)����˖+����|�WO�����+���Ve>�:��<i��/\�A�D���Q�wk�q �s����^�RrY���ʪ�	��3[���k�	E�rm��"�i�z�d��g;��7\��Ctjm�I��k��+q=�W]�3[bE��j�a�֠�Mr���1�H�m�z) ::S���S���*����-���/fk�bZ���Bɺ�;�<%9W�@�7���X����͊�J�7n�1��*b�eoUÓ*�hnKZ��2�U��
�����W�GI;�VB��Qs��c���Bѷc��{+$�58�"߲�n=�ۮ�^!�]t���e�#�\�9�:��;+��p+�\�����\��6l��i��N�!n*�1��]���YZTN�T�B	�:�w�e87h���&�:��I*w�t���nL��t*�vO��d��^�䡭]1V��2c�C�J	w_f�9z����X�Y�(-��(<m﮳���ז���><���xkZ�Zֵ�c�F��k_�ֵֺ�xkZּ��k�kZֽ4kZֵ�{k\kZֵ�k^ֵ�kZז��u�kZצ��u�kZ��kZז��xkZּ5�k^Z5�k^ֵ�-�1�hֵ�kZ�Ʊ�kZֵ�hֵ�kZּ5�����kZז��xkZ�Zֵ�zkZֵ�k^ֵֵ�k^�ֵ���{����#�FdC|���G���kX�=���j4u�E�m�.n�(�ܦ��=�@�<z�]��MS�u���Iҟ{2��m��:]��&
d�"����LI�E�t}|%�ht�T�TOL��N-�붒~��).�4&�m�]��wj��t��iΥ0�z�;���b�adʫo�w#=����)�ڳ���7P%:+�
F���.�]|�d�G5fA����;�{$.��\���H�<�-W[�>��9ۼm�2-c.,w�r�Ƨn�z@��
��.Zn�:�<��F�%��Q\�I6G@����7�� �*�o<7�"*����G'4
.h����Qi��s�R�Û�����i��W�ܨ����]�t]+�B��Sv]:��K�uT@c�,�17�b��v�[y`V{0S~H�l3�M�f�Y�r���t�w�ΰ��pu�S�X�Eֲ�`��P�z��ܕ:���tg�J\�l�,Vh�wh����Gbg	�ë�.�^u8+$k6,��"�u�z �.�E�h8�ew=r�Cgr�WUm�oD]B�α)��pV`�JK�7�W�v�u���As�n�1;B��.طU
��Ֆ �+ Z���W[�u��7R���s���V1Ǡ w�J��kҽ��b����Q�^Vn��r��c��lݻR������FG�ccѰcb��k�Zּ5�q�kZֵ�kZֵ�|kZֵ�zkZ�Z�ֵ�k�F��kZ־5�kZֵ�mk�kZּ��k�Zֵ�k�Z�Zֵ�k_Ƶ�kZ�ֵֵ�Ƶ�yk�Z�Zָ�kZ�ֵ�k�ZƵ�kZ�Ƶ�u�kZק�������kZֵ�q�kZֵ�q�kZֵ�q�kZֵ�q���������6E�S�g}r2l�[�UU�$"!��(�����w4��	="9b�l���8�8�����9>��t�qX���P-�c!�c���L�S�b���	�:��K���0���v�e�N�������B�řo�L����}4���w+���&�P��CS�8�ev�,���>�s��{k�<�H�����ѕ]�t��94�ye+�n���EܰU{�y���+��bl甶"���;+�������ڏ]n�:୬��<jT�y(u�6�38���T_[�&T�������\}�vđĊ��@������Ý̋= ��7j��t�*-�W���N����+�PgZ��N�ڬ-;�fX�-�Ob��[���z�bR����Kl̚�2%N[z �WlV�$b���<O�"͢l�FHԵ�n�l�s8ДUa:��n���BZT���tǍY�N՗�M�[���0��r��U��e*�c�j=�.��zM���jR���y��]��0����U�xIw��#��yU�@闤��[��h�I7ͧs*�uāp���lO�ǭl�5[�WRH��K7��KJ]m`�:�̫�����]m[詮3���y�D`�O״���O�^�6B1�X��3�@�ې��=k�@u=3V�S��	�Ա'C*�8�i�Q�[0fh��HVF�1�;�wKyz;V;�*Q&�Xc�(>��T�#�����J%�a%��$�}L��!m<��C�;�c�{�@S�j]F:�7A���)gVik![�m�j���Ǆ�һ���>M���xun�ݭ��;.����ibUn[�Զ�E�y]�	4UY"��,�(�q���y�Kq<ۻ,D�D���\2��_;]q�u
L
�7X�Zo�u�L΍6Ea۬aWj�9�c=��_�������)ٻ��J1n���F�j�&��k)���3�̇1r�bkS�jz�E5{��u�8e��w���r�1'u(�&��[Ā��,g�5فqB��H���Wf^ܗ�e�.��;�v�[U��E�	�����oQs9&��y���N�2����O�^\��<fX�m��䙾���wV�XD��R]RfP��Wꠋ}J̔z�i��:�EΫ���O���>��q0���/pUk˷�ă���5�^9���Fc�F�(nwv�!����%��Kr�;�@��r�vÖx�T^*�u|��-kD�ޫo]�s:��/t���x�;1�*�(�C�2��&�N]<4G��9�c���0��i
��Ǯ����'��Z��ޯ�ٜ���F����-ܽ�r�:c���6��A�Lg'�p̫�q3�zb|�|{-�E.����[T�:v�$z���Y��f��ty���.��V��Cez�
\�ԩ�b��l�\S�)k$N���x۫���C��c�zV_*�!Sv:��L�M�Jm�t%�O[��!�}}=���@x�V�QΔWXA�n�i�֘�=d�l�� H㙃.�G�ĺJ"lU���AF�7�ar%��r�@�v�幁e�� ���=UZ���4۬�1���GŎwN]w���Iv��Ӊ�ܹm,�
*�e!@�[8M��z�7����-*��U�.�](�*��R&�[�3y4}�tַn�{��޵t���&$OR��qPE�gS��� ;�Ī�\M܆�������5X0�Wq�b����Y8j���5��BbB�Ci`�C������މx$� �|�Y�i�vq�maV�op蘢�u�v-��c�U�o�W�x��+�R�a�G��f��&��vp� y��� ]�f���� ��Ύ�U�iQW)k}1\#2��Z�39�����~�C=�=�X�E��� 6��ji��۽h�fM�wf�S�1�ܴ�s5 V�:�@��ӝ�z�/�w�G1Ἔ_,�l�y��ں�{=^��u���JWV�L�N��Is�3[}�,�ı�T$ى/�/�����=e�+���zؠz�Ջp��2�[ϸ�ip�)�~�{��ۣ�eK�1��S�4�rv>7��]�꽕:�uˤ̄�����f�*紱��J��I�+[Wu|�я�t��[���B��n5���[glN]��X<tq�Vا�);KTp:�m:�"Z��K�%���v�m��:��e��)uZk-��f��6=U챊L�4�W�>|�<�r]x�������-�4{]�/K�!�Ќ��9��_c��gM��$�Т:��z�A6�7�J7����㫎u6,�4;�rW��>�K�P�f_X���K;0J�w�f*N�=d�s��K}1����S�� Vm�]��r�;���(�{�� ZӢ��NL�]��cf�R�v��^��W��F٢+�=j{�)�}�����Ρm���dj��f�쀢������oL������O����`����3;2�P�a���S��ӽm��`>����^��K���Evц����V p�닼z���U���DZ�*�k�ƻ��8��A^�崝���.�9�3�\��ǻs$N ]��\	�p�'��n�q]v��"廮�V:l���{B��_ޞ�L�8���cjp5.�Δ+�=4���3we�K׎��mI��꺽8B��A��Psq�w.M�[J�s͐��|P�7YMkݮӴ9eF���h�ïx��V�XK�*�$6��T�ɛޠU�(Ԭ�o6���6��9c�	����4��]*^y�_Yh
8dҵi��ȫ���rfc�����b��.#��1@��(�zM��ˢ�Ƌx�S''>�=�kO��wvh��m�M�tv�X���E��3e��8Xwľ�:��_�]k��,���MKű�+��YM�p�x��	C�ɘ����5�I#�y�>Gx̝4k�
iʯ+���ޤ�.�c/rj�=Y��9�����Wvj[����Sxe)p�[I��V�MN�;x���N��@c�]|0���,gSZ��}�1G:�N\�����<��v�3j�@۬�F٬�,B4��K���V㽻�`�;b�.�^G\�~L��O�46q��ά��Q퇫�����t��m�M�s���;�YM��3)aqf�)���!�Gv��wLH��v�B����Wv1�!Sv�M�ڵ�w3J��=�O���]B6�W��.���n��
�k�ʶ`��dTս���t%��^ї]`�
Q��mLg	�[p���3C�u�)g��Ur�0�x�׆���|hJ�u*zC���뗠�c!b��32P��(z�7�-o651aV�`�*�z�	���W�y�+�>b;�x(�+���������s�6	�X՞�;��F��)�u�586��i0զ�3�� /(aw�ݵ�􌱝K�h�S�p7WTb��6�;H���wR����f�F��}�kNvf�7�kb��Z��-�Vj�`9����r�$�}��i���|`��iaoz���\,V�N��ټ7�wyi�-)v���o�fX�C6�FU�ui�:��a|�k���W'tՎ
BOv�9D���:��{2�����N�s��%s#]qv*�j�uf�n�4��S�D�v�)gJ��bV�D�1�θJG��k�4�C��nU`��:o����{��j�O5rձA��۵����G����>�=�w���=���l-���u7C z�rt��B�&�2�q�Z�e`�Ms�5Ҋ7jf1/�u�Y.uk�6�[;(��j�j�ά���\�K��K���l^����x� {��n���1���:��C}�s���WҮ�9]\��ȷ7�՞�;rAg���K; �V��sr��ᒓ�&Dz��oc�]a�;���U�W�R�)�H`���j�E��	��	�
�tc� 2�U�-Cɹ��L]�eWi`��404�f �F�6����,jn즮ix�LQ�w���0���f
s]��oBx8�Dd�)9IE���O�kא�o8�U��w��[}|�<t1�T}z{�e@���B�"��X\��=��jU�;!oT�X��ţӋ� �炠�1����(���VѦ��A��L��+�Z����6��j��9��u7�3*c;/<��y���ٗ��X�]5X�Z�j�L>�ࡘ�0���"j�"�8"��ee�bpS����Ria���*���V뫸=w����o$��j�cܬ���C
xm�ה��D�w��[o^ۺ��\��,�o(+�P4l��x�/����O�];
��Uyv�t���xK�ʇlb�>����!B�u;/gv&�7#�0X��;,��[�􇮞��n<��$:�ǃ��|j���;n�!H�ό3�ܻ�\�6�+����� -�^�� WՎw��t���t��%%�[���]}WƫּS'�<�&������Ed��V�v���	���3DYȽ�΢Io��Kݼ�JR�ur��uν̨�E�2oN��WNc�Y`�>�N�s��Cw��ϴ U�Y���w�}���r�C�?�I��\�?��E#�k�H�A��?�۞�
t�c�6 !���r�n�z?���P�R�Tj����h��/S�����ψ���#ѻv�K�gV�E��V���Ed�ʙWÆ*T�oISdUpۗPM�-�w��t�)P�,�K�|�-,���CdheM�|�MVN���2C�5�s4wX8u*W�#��%��iߗtU��5sg4=������2:o�\���ǵ�{(�حd[9�Ѽ���9�n% 7+���b��^���P�Q��7�1������f�"���;�L��<����\Ʒ�V��z�S���]�j��p8��1���W�W���t�9X�pqi5v��]n�M�f�MsШ�u���^��y�۝��E�G3�ALR����ׯ�7-��C������K/�{F�1v�P����/���'Z�����V ^VA�Ɲ�kf�627��r}=�j�Y2od��k��w��k��e[5�{g�e����l��)U=xf2���Ht2�$�WSv/wk<�Pz{�� 4�����0*n�&m �rV���2�m�{�+�	y�-�z��K3h>��#�o�h������*�۵Pd"���Ѱw�$��f�y�T���:j�5��'�ۣ��g]�K��8�iӥ'h �E>��_wou�J����Q��@i�и��9m^h�=WxJ���@�I��(dt�T�* h��	: �N��v�"�~p*�<�x�^"A��u4�EBTSd�"`� �Y,�([-��(5h4��U�(ZHy��=�Ƞ�۴i- ���y����~o��ֵ�k_���˥�"�W�s�\�ndn�N\��Z��^O<�}޵zk_��ֵ�kZ����ח�^__���]��߿+���v���z^b/]��k���"HI8�$ޘֵ��폍kZֵ���~o[���{��z�{��ݿ�Wd�\d�忟n�*f1�o;ו�ᐦL~�I~wy"�qr���@�$��Ѐ�i7"�0
)8���кw#��.k;�|w�p=��ج<�K�=y�ζ|�ؔ�[��r�n�^^kEx�t][w����/��W�wv�.;��wu��Ӥ��4I]�;kuΝ��w;���\�˹�wj̝���ޛӷ]�koݎ��23!�8�a���g<��']��w��;��pu֧I���x]�צ��.���B�'x�x�wH���uݺ^޼�㧞=��z���r���O"x����r�۸��s���Yyiq�I�&B0�	�B�B��]㼷uמ]^qΞ;1��c`�`Q�1-C��
	���n��������\;�@(0�(HI����9�S���������GP�V���,`Nm���y���Pvs�'�3�j�eK!�*��fR���v=[�m+ֺ���1ߖR�%�v�B7vİ��@p`���N�����p:e���{&uvΜ껺ü�Q3���r��Yf�ϳ��9�I�@��f>bO��*̧F��n榝U4V+�F<�"�6cΐ�JB�*ᬍ��J�EO�Ik]�6�{��*◪�ϓ��"�$�����Sኄz�c�pk�R��4K���vn1V%�� �l���T�F0pi��O���j�'NG�B��e�W�m^N�ٚ�/j�(l-��u����z��0�n�ᣍ��Xk�!g_l�f�[B�(�:�n��z�kpUe��Z�|ۛ>�G[�I���Բ��N�L0��n n���
X�B[��`ߩ� mre��Zc+���N3��x�P��DLdfQ4R�1v�6NZ������|������H�wY���Kn�P&v��@�Np���(1B;8>��k�����6��&�}n;�
���f��\�x�	F|�v^]�Ҡ=:.��4�OҕF�-�ۗ����%1Y)�aP�vQ$�ֵt��%q�|�R�r�7p�ʗr�n	ѭ=x��m�0F�BrV�2���� e�y��7or>���Hj�0󠢟,Ȁ�(@�z��t˻�N�E�-�6����"�E��[;B<��A�A�Q�����3��1#J�����ϳuH��cIh8(�v)�;AN���3ĩ�5%3	���8&�̲�;�V$���ϫ{GT���\쪬AP/j<�Ӭ���g�ǽ�꺄I�)�m0��o���U,	i�����.�N+�`6bˍ�4�hk"���x�#"�
��
s��Y)�>��4A0L3�jZ)��ff�T�7P�iԁA�*�P����e\{��Z�|Lգ��M�;;heyC�YU��%��;�9S�X���+��u�u�gU�5iܔ\���U&BE7��q�N�Y���I�g%X��ld�T�`t����[l3�除|��ࡰp�d�2[8ʴ�S�6�����Y�5+���&�hcG��Խ;a�.�=c�%�+��r뛭�dE�;3%wn�y����7|X_TH_AfM�+r�ǯ�M��t�Z��B"N���zgu�l]g) ��i�; xG�:����ngi�����������P�FJ�y���~�U���(ux������m�I4�[�kf%��&E1�R+��b�'��ùɍ��e���[
�z%�Q�^����*�[ٔ��v�`��s�aNWmy|����V��|s�9h�4'eN��m,'}��z ک�V0���!��l��GU�� 'melO��pZ�2��w7z�O��$
x�;���;c ��P2Cd�`3�B�{G'!�-N2����Д��t�����$�V���K�CМa�B�V)�7��EjX��i��Z3b�mҝ�;�b�<Hq�'g'����˭����sYL��а�;��is累H��f}�����f��0ɍ��k1I��Y
�bШ�8*��!B���3(�g�6l���;V�f�H��t�knR���0g��B��v�����m��&o,&%7���Ҿ��k��
�SJ�w5����̫Š��%ܾ���įz�s�j�o�ĵQ��X�Ӱ��=�B�����vM_1�+X[Y���>��k���u��1SQGSu���Gz�G��|�*���xUP�/�_	�s�O�b@�ȿe%8�{rE�9�nz�X�ޥU,I��;�ɼ7����9�t]V ����4��Ϟes���f�uY��(O�6�?MX2-�~m��R`�XE�А�52�}�!{�����?�EU=�{.�d;*e�MW[w��I�(�qE@{�}[Bk��<���{Hl�m�d��mC[,���꺸�Ɲ��CB�t��8�6G��� |L���c�m�󤞢6�vV��G�&H�Bo�Bم�F7mC�oJw�k�[v�I܉t���K�voG��츨�|�� �I�cQfi	}��'7n��:�ZYًxx:)�QAVB��i�0"���w��gmeX0d���Ƀ��z��V+�.v�K�g�6*��yJ�k�^�9�,/XO��Ub��gF%���´���#�£�F�vR��sj;(�}�΋��-���T����FuN��'[N��:vj��9��箅 +��n����I(���i��p��I�.Iq�]Ó��sn��P�����������M�<ͳ�.մ��Ǖ��%�ʓMRY$�L����ib�~ݟ�I'l��"ŗ�Q���R~�������<g_X�p�}NqXcUSć�
�o`FԵ�� ��v����W>�t*N��#t+~�z��ڒ����li�F�F<�ؤBa��7�"&�/!L�uv��؛t/������J)��+)Hا���5���ٺ���el¼l��>D�/Mf�4hω6�yq���\�,����*8���Z'iáBq�O�V��d�Vu"�T!�v�UP���$ثy���Wy�i���
��zn�ܛ��R9��fH�	P��lyPVZ�����D�#Rq�����4�}qW�>G��0�$Aq���.vǯtҰ��9U�WW7�T�}�c�dڂ��H�lC�E��W���u��
Ӻ]�6�\Y�uע�
�%P*kȬi�>Xt�8!�6@ht��M�a�I��~���;�i��Xt��ê
"�[�2�mn>;aW��r��լ<(�dM�EZ��C��x��/eL���d��-��<���ȶ�ͮ��s�}5�Ja|Ƶ���ه���Mɧ1�Yx�X:�������5��Q�p���o0���f�	92�j嗁�v#Ӧ��E��,�q���a߇Y�@�ڈӍWG^��j�tA��gf6������X�A����16��۫Xcw4�+�g��;�f`��Z��#6F�mxME ��3@ǧ�V��j�O�8���0�N���~��շQ{|t���~Gzt�lVο�=�B;�(J�q�Ǟ�W�H{�B� ��$�v�-);9�1������@l����8CN�<M�m/��p6'@�m�.{/\�J[��2�W}�u����5�j�vS��a
����_s��:���fNi87ш;�������/�R^F�V��2�!�)4Q�/.�&�gzX�Y��q�{A����U}�L���l�%ZH�.}�g\E}>>���-��Smf�����,�������T��i�'`�t$�뮩���]yC^Q��y�K7�q6�K� 6�7;�E�ܵ�<�6G��S7�����lJ��������|���0����Xs��k[E�.��*�kGL��W�oE��;Y8�[mm�-�⫵�Y��n�t|�rHy���1/I�n=Em}Sm[��A��HL�b�Nb��-Ǽ3&u�i�8l[yZ���(Ҩ�3�{,�M3�.�u�ٺj�.�O�!�> HmD�x�^�}��_}���>xZ��n�l^Z֞���=�v=�)/E&��¼�2����l�JQۦ�K��N��3�21�[0F@�Q+c/k�h�E[���,!���5�k��RI��u5^}}����wY-�����l�eZ1I,����eDٻcB�l�6m ���.�������9Q�Dfa�:ot�>�n�V[�%��$Ūpfov���F>���U>`��f��j4��Lv_�}U,�o�	mN����ͧ�/�jz»$˗.��e^��\ҍ�^&�`8�}�X�òd��V�����O����^4��½��]���uhy>�	�����#�ʺU��_uMv^��>�s�^�U-�-u��V֙�`I�U�>!]tX��ԅ�SU�p����F���"���}�� ��뻃T�=�sxu�h�~M���1͍�f	�2)��+��H��9Y;�dibH�m��ڐ�iV�d�{�0�7�a�1����#V|��y�p�He5	]��h�`��������s�\���o ����C�(z�����u��^c�`FS�/�ĤZ�����-j�-�^���]V�}+���FF����["�;)c]�M7�VO�B������}��z�<�'1mE��f�%oX�U7���W[��/�P�	˹�VO�ٟ׮n�P�^,Ep�܋�*��*�nּ%A"�:��-��y�ﱔaV^*0.a䷭8�H!E蜻t�k���PlҨՙS���yRj�|�G�.�������Z��P����[ߺűQ7�:ȱz����	Gﶉ�4�@���o>߲C��0H��؋}|"��F2%�M0��]�b��H�^�`�S���`�����oI(������Ӭ�nN��@���	�S�,��G�v���yݞ3��j�q��ݒ�;�l�&�
l�3��u�L�B�942S/�i�[�0a�|�� �m����z^OPK��u����ffA����2�
�{lm�M0��H�;�N���j&V�L�2���ma֖q���^
�(72�%m*�����N`K���2v�=a�����(�)����AÛ�*(ɝ�2	մQ5AN��>��G���l����S�kbQ�"<��������(󋨜02���r��1� ��"����&ꡞW���̝�f�@l��Y`Q�{��P��tn�2�E�f�Xc*����.�K0F��c d2��C�h�L,."��UL������X�ȓ�N�l,0U��OSa�0���Nd2�����$��[2��V�~�4<h�@�O^����<n�������]�u�UP�L 97Y;�v�� �"�?�m�	x�5}O���S�wt�8pzףs˛�̋R<�w�ڣ���6
�u��ʻ��g��fhSGR�fU��nPܔq���W����f`v�� �mSX��kZ�w�7�9;?)}�N��( S/+���a�-�e�LVZ�}��Lw��,�w�/���^+��y�]��R���_";gQ��kKG#�xp�q��f]ͦ���y�UoF�i�ܪR��Y6����ɓ:L(0`��t�7	7"UM<	�q`���U�r6sa"ئ���L@6�Xk`���A�eF�8m��an@�j�Q�F-�^�9X���f;{�-ϟ,M�W����)$����ji7
���
�!ݛ3虠��{z"!N1�4�A�Xm�_�E[d�Xt�3����Mr�Ӓ��Y�i��J�09Qjkz6h��n8-��	�<y��M��;�ޚ���5�;z$��¶���X��U�8(�Z��+�6U�A�xV�TBjLn�I�zg`�쀫g^C�w6b-LB�ͽԶ�%�M1�+t��giR���Xd�eL\��x�CM�3&�3Q�m��e�T�Y�4���rfPJ2R�m���zϨ=�6[(�q�.�ܙ���� ����� ^�m��<N|�I��/�Ǵ_AT��P�Z���y��Ӗ`f3��!jm=�1Z��l���W�h�x��2nf��b)�Y\[��Ь/�u��9�fҙ���S��f?��mp/��%��]�!pٌ���T���]BP�@�ٻ��w��F�;b�n���`�*f�� ��<�S���`���[�Ԇ�"����*�����nF�(3"2�������� 1!�o/8w���L����,��iN��i�U�LS��Ya�q?a(+��#
��/'[���������n���gj����qho�k�/�}����R�Nn�t��X�ʴ�G6{g`��y�.Vc�q�Nq�E�d��l�*�&YJ�z8ݬ�=���3�kXKL�C�Xh�`��y�.���M3x�y���1й�\��=�
��-�x��,;��bК��BDuú��!����k���/_�<����{�}g`6ˡbf�m'K�w�j��T�)�%���M��5=Ѣ�R�Q�h�8e�����Ky���=��Y��a �]�j�\�����i�N-έo��p4]Dk�Y�vt��bIӠ��8�E�"�v�n�O����FZ-�ݞxK\s�Eo{���޺C���OSmc�8;�zo������ኬ⽥ϮRb��kb��NV�v��.Ş)t��sY�J�-�ir��}�(�ȼi�x9b�B7E��뇍�^D�6i����ᣱ�b@Lux��w��^Oo���W+��
��t1e[`Sg������MϪ��M�n�Vj�3��:���+���^[.L=k�T�T
U�rc�/2��z��+۵��Rn�2�i򱒜�:���{R�=v�4���S�������JB��T�IŘ�Tӆ&���PyR�E�w���6��c:*��#zJ�r��)l����,���4H���
A���n�T\��;N�����ddŦS{Gx�'z�O@���� ��f����p���v��W7A�h윺ܥ�uL�1�-a��4Y���.ͣ{9�|�3+�2Ecu)(\�L��ai$��!���kS����d�w�>ƺ��nuְ��w����������]�R۫�r���Z��B��n02�ˠ���k!��ɰ	{��;�՗��,�Hw���h��R��0V�ݪ��GJ�fD�X�T+S�ƳK��׀��kX#�
��t�U���߂�O��*��|v�9M#�m���Q:�WyMT5p�Oz���vZ+ax6���w�:�D����F(`��3��ԤjEK����J��Qw|��ļ����^�yv,n���E��%�Vn�����7C�C`y�N7+B��_K�����m��ZSJ�r����%riɐ=�¦mK��x���(P�hP�GC;�+�a��:�˸�7�:�^�02M�	�����5��>��k_��__^���G��FI�7�n����,}�LJ;���&��]�I0I&d8>����׷��___Z��Ƿ���ק���x#�w.�n��1d�����DJ	�4�H$�L������mz{|k���������oo���OO��󻁔���7��l���ޜ� ��;�}�c&0�`L�&^����ܑ�!�+��}�}�׷��&wv�N���Q4��[�D'��h�/;�f��WF{�� #}����:|��N�<����"�Q��i	�"�u14��) ��v3'v�\����HH]u��ȁ^�@E!�E�\�\%�q2���NI1��/o]�$���رI2�=�������^R���!�_^���:jL�i��K.vG$�z�(�&3�cO���Yv/x��Z�|�R��(P�(
� N�}��5�/<���V7��r��ۮ��J<�����}~`��q�P�ĳ�^��A��W���@�A��
zQ���f���pCWF�#v�RoW�Aw/"�ʲݻ�����[�����g) ̖V��W�0�<��
�ȉ�LR��;��V��� ]8Ú��][�[]��b�����Q�w1�d���y�����b��=�*#��@�V[Mx�9���%M�)�j����!�ê$�%�E�;�c��=[���Fy���1���8���i��iovCZ]�xצ�9�Ɇ��\�H�b{�W9�dcR��X�OE �)!Q�����{�ٜ�+ǔ�~�ٟ�<Dw����#�Gk�OWvt����}\h�S���� Ǻ$��W�,���͵��	� ���D��p���z�Sp��Q���6(�e������Ԕbp2�s#���u�߳>���B�|GX��\��>p"���m��iG3ǧ�\Y�~�d��.�P�c��~�̲��N\�� "����ap�xۋ�m�F`9l+����KL����*��B�k�ODD��Ji�Q^���]���?d��-�;Σ�ݶ�wK:�GH�uB%؛ï��M�p���[v�-R�u��у)۝J��]x'A�V�p���{3�H���.�����l�֒�^ͪx�hs�|���W��>p�!��y���gV�^ ���ιkw���YD1�Ǧ@v�g���6��X���qk�y�!��7|��{>_�P�G��S�(qc]H�$P� ���HyHh���5�w��>sB�M+3۠���y`�&x�c�|���Q��6qZ?j����|��.yz�V�"5�U�	�y���rw�9������D�������k���ᕹ+�QNf�W!�ᄎ7��i�M̚C����Sܳ�Lά���4�1I��?|5L_��zc8Mא+ϑ��*� ��
�d�;0��*���7˳N��#p)�Z��x��+��֐�~���7����.�h:��'��v��ǃM�T�t�%���N,1G�,��ѯO�P����	F���솭��ͱ S��~�v��j�*�w�;�@{̟izc�r�)�[�~��>�6}Zŕ�H�����L �ڒ.���e��Tؖs˕͝c��
�3ma5�^���w`��L�R�g��㋇�uz���8Lv�z�1c�N���8�{Z7�R��ū8TM�,,|֮7`eWʅu�z�
j
��u�Z���5×��o��P}p���b�������>�S��^� dɗQ�^wۥj�xoV/=_aW}�8}|��Lo� (v�@��E M0[���ɪ���.�i@��x_��u�g���˫Yy-��\�Jgv[:�:���Q��閴a1��p��&������]  �K��IGiAR���a��	&&R�����~�A� ��)4w^�w�}�ؠ� �g��sz��˘Iן�M����X�㺵'˶;�����F��9�ƺ��x�ɽ�s����	/M�@���6W���u&R���܁	OR�?bx	���(9ܛ~��ĵ���ZM�����V�Y�89�/@;ݸ�q�q��C\}0��cǈG��ZV
���9�"7s0�RO�x5o��yغӨ8>\'�)��5��@�9d0(�pBK���l�\�qK��;�|X�S�%F�2�9p�N�<-Rk�]��^��B��W�����28��cX����.>�[����U�]���@{XkF�Kͺ�&|�����.�fi�����o���N�Ӱ7S�ܖDMOek�����=��ʦ2���c;�Z�O�q|��M�kk�	o}L��맚��0�9�y��~�(��!�C�A3ß8y�;0���>�t�I�ֽ�w0Ѳz����E����/f�
?@sU�UL�a�>�?����|5@S�?W�TTn9�f\�h�f��ڤ�Dv�Z��ٝ����.�E�_�C6�׻�����[q ��)I�0�|����E:��?*4�v�2Zgݯ9�Y�ʣW�O�������^�/T�7�r��dh��jj��]�E��Wt'O9G6GM2r��gZf�\�G(k��!R���8_V�\��ZO;���v�2v�9�}Z��li�7c����Q�u\��ё�dc��y��y��D�C���Y�3�p}��|Ń1�}(�}�	�>N�;X�7�<"Ӎ��&eGMjiӨxn�$�ړ@(�~��E�"t��e=��WU�oe�9P�5F�'H8K�Q���[�O��j�!��j�(>��L�"څ��2�j�<��<��o3�͐1�:V��v̳sq�uF�1���΁�!f�(��P�'T��ެ��G5#�����+�6u�,f�yb�A#\�O���ʩ�7Ȝ{`&��=�-q����P(��c잘�+�!��ԭ�ζ}X��S�}�.��	���u���Y~xQ�mbR�ǹ_���<�{ ��.x5e�c0�|]VN��,2��w׀+�<ۏ ,}L�ȿ{z)��O7��;��|�`y������;u�G�݁�i������xg�&[��y�1���f,���)��ck8d�E(V����@hx�=nZ=m�`�u�n�J� �?���Bl��X"ԉW�o�) ˁ^J/���Be�:��� �f<�j�����vｷ�#Ԃ���r�,>+൰C�~���l��Z3��Ժ�����F�����H��g�O�9�Yv��x��U�1�9�'i����ʢ3g?�^io����}S~��ܕysȲ:�|ӎܽz�/�3�;�a�.vsO2�`G�ot�JTjM�Y|�@���7~�\�,ţgڏ�N�A`�0`�������n���t�CM%/�����q����$.�L�g;&D�1/�2K
�=<^{��z��5�R��J�ʥ�[mT���UĂ�:$kpVc�!���Z'-V��?}K7ۯ�����n�Ѯ� ��\�{��@�c�;�ܡQ�@G��HE�0��/3b�0%��>s=��(������
��	�X������:�T)�
���2D��;90�5C�OSI��i1??��J��E�].��7w/t�j@��L�{��15���rm����!
J�h�����Lن|/���L��%o�U{�c�^Z��8v�ư�t�.z��zW�	ݡ0ul��?=�#�@�N�G`��ג���M�w�����I��@ILX~2dp����%��4�-O�#��\N4���L5K�qo,��n�^q�7}��
�H��E|6�EizB�e��,��&��ޡs����ts^nϴ�r���SooO7c�:�1���������T-�sb@�#d$�ڗ�6׍���f����`h�.%���_ߤ
=b{�W-�g�VQ�tR�������x�;��<
��[��t����A���66_7\��@�9o�ͺ��#�d��#��h�Q����\�f��rL���[���-���vr���iK����z�ևx!Sw:���)�S�O��5�����`�@	���7��I��*~��W��{�_�d�Q~1��.�MԹW0��ۚ�Q��~ݤ���u۟a�U�F�i�����1�c��"Z�@�i���{�H��Ws��\��0)S�Q`[HǸ��Z���4�O�w^� �ꣂ���!�����:=Ѐ9��0C��4��t���.��}]˩��~�۽�La�N��
�i�T[C{vh��_}!|�BXf�X_ϒx|� "�`������
*�^���Nw<�t��,7���)��.��}��F��M&1YDv(��G���L�������N�*\�����;p2���wOr�Q}�����l]���)!cȂ�������y�Z�	WW�+!w��ly��%픋���Y�,x�Z��3\Li7'5e��DPh�|� �od���m�饲����+�C�Ny�	�=��K��F��86�M7���r�>Z~;Y+�ϥ��MV,�Wv�e��2�+(��k���3ؾ�%�9�2A��r�xP&%9N��]�)t���6��=c��t� 	Pu��Y^�����0[Қ���F���p��A�����cG�y��4��9�_A����u�@zM��H+6�\͇EE����s�ʒ��8{�}�{�~���^���a�%n��^E,"!t(j:
K�:����K{�-�}
�8A?f��.�8�O�Y�:���E$���[���Ш���slW=7��%Z���ESҥ$[�2�DU�p���6$AP`�EB�D#�(}��{���nB�z ?J�~�����L��T+�z�*�{0	����pxC��Q�W�𝛳H?WWmz�}��n;��HP�z*ݓ��|���l�Eޘ ��~T�����]Ⱥ��{99��߾������à��p5�'қ������D35éS����oCL:�ʵ�m�v<�U]�Y}����	�a�>BCQ���&��Y��cO~;	�z�O�������涱�g[�eGOp꯴Ѳs��\�a�8U����`]/�lV0� 8�X���w����GlP�ۙG=~�l���[�q�ޜo	�Mcd�d˹~�x� z/Xcޞ�?:��M��N��
��ux�[ HP'_�"�S���P].�Ӻ���0t��rސ��b���������i�%��J����n�'�}��۹�Ǉ7jx��ԩ�|�H
/�86g���4�����bhT�c�Ѽ��~vk��Բ��*�O013�8�{��@	�*�����?cX�.����nwQ��.�fye^\���Lp��З��Ci���<����ԛ��<d�U��Ú����V��Ǳ}R��T���^^Z�S:���A[�uqB}l���W=���+y��Xy5Z��[����"��Ê�^�i�2A���{���̾�yP�.Cȴ���cP�=9�\=�1%�b����\��Ut�7(*��<<ݪn��6�ٻW,�j*,0":s>�73���@A�pV@1rC��Bdކ�J����(�o�C�.��zn�ok�e�)�9ɴ�Q��\==j�ȯ_��6������XZcL��뚝"��G���(��m_���(V�Kn��"����N6�������N���|���`�>axK�l���"]�>30-\7�[�+���=� эa���f8���ȸ���>xk˼
���<������}����'@Uū�F�0[���#�U�TL����+D[v��2�����CS-�?x_�''I^C���?	z����ߓ�e�� �H].���~�:S{ڶb��KjY.ٍ�����>h��@
HD��VCG�1Oa�{�d
�M{�[P��Z��Y��xcy(e��>>�i�TyV�~Eo��x���¥�M~��
*�I4qc��!j���(�([�	�c�B�G0�����U�=��\.���'�K� =����Ҳ�p�ٙ��tp��~��nx�ږ�qg2��sWxVj>�?*�������q\��?Nb�<�� �!�I`��9��/G�*G��ge��:��x��2o��kfM��ރW���FIp!u/tQM ���K�v|���K�/��e�t�ýN|�`�b�	 '�:�-P�u��24�h��8{�]�ݧC<�zVݱ/�,f�*Z`찶�*�}�k9E2a��o}sO�?/q\P�#"� ���ߞ���{��7��/��ٞN�� 2籽�C�W7�y�,��=܁�ŅzD���[�vP���^S$Τ�w�E��lw��5N��2.9;��~a�`.��~����Gc�Pw��y���S�{W�ue��l���8ZTǁm�Y�=q��4���{�,{�6yX�<֐+��^����� �9�j�;o�!�;=�\k�B�����e�c��&����T.�K�/Wѭй���q�"E�� �&��|­7v��PӰ~K�|��ƣ⭭� >ZGѪ5�ʄĶp��;E��5ʌM����6炙���~Гܽ������eG���m@ـA� ��U򖏌 8Ȫ�l�|/���{�����4�s���0T��({*}:�>�i[s� �v3�͠�����eð�i�ə��h��-�V�C5:�3Hvɛ�\X2�K$�C�Њb���0xm`ݡ[A\�W`n�L���,�݅��KC�BGMua�7S�]� ��f>�������1N73XŤ[����� b�"R�e������1Q�w��4\�3��5��w=Kս+�qwF�V��U!�о����;F����5�����~��
�li��K9�[�;��Є}�0���]X90̕�(&\jt�Ә#H>1�m�� x���&j��u��E�[Z}}.�О��M��W�\�x���-������wa�Jv��G�߲ꪏ�5sk^�?���!@B��+}��ץ����{���|��Sa3���%O(��:`K�g>_���4������vR\o^n�TQ=�19�N7���(>l_>�{ .��)+Z�Qaw�Js�>��N����k�8V���5{�HIz XB�P�l��Pd�� O=�:�栌f=p+p�?,$�p.l9 ��kjF}]9�;�]Gx`����æ��!� ��,��Q-��+���>��֡���סcR<Nwq��ug�܇�^�}��	@�^�����D���Ɵ?G2O`�Jp:�H�������sP-[�A�gڝ̎ν�o�JmI��1�Y@}�%�z
�0��������ρDs.�3�KK���x�8�e5�n��^[�y�7����^p�dP��~��X�-��&&8鱾xzW����.K���d�W�I��lHP/v%����{!�XX��j��yZ��U��n��	ٸ���m�t���	D�������:���+�$>))���H?�p9�뤣��J�pݞ��nhK�0�p*���ݲ�5��»cS���}�N��s��@��<�L�*�JԺ�����oǔ�~�(�I��ք��n���}�6^J�D��J�xim䝸��mB���F�C���Y�1c�L
2��@̇8�_]�����u��ڼ���ԉ��62Fq��tŞ�h�����5���}�gmENn6
��P�chY��e
������X����WMX��3��g`.��W��.�6.�6D3a�h�jż^;�ܼ�Z�{:���L��Eu#�%�&�V��CS�[��è>N�*�� : sz.7���{���K�K �p]
�K\�j�㼱�&o޴[������p�4:j�e;�8�(>�\õד��e=y6�1����q���9��u���9�v���hWK�YNF��]�l��Z��5���\�1Q����ǀ��}HudX��Cƚ�ۙ7[K�ֻ���/)�\��h(ᾡO�؛�m�f!$�d�=��N�'��";�D#Q�'vc'L�]k�5��-��=r��*���y��ǆ��}��&� �I(U��Q鳙Xg��u��-��N��eΛ
��=$$wT,�ޭ�;N��|zf��@e��^{:O�Gh�[���.�b��©{kU��˓Qꚦ��Z��渨�/k�9���L����3"ʇ)Ԃl��aw���@_\*�[R�l���5*
���
�Z4ޗd�l��~)����$�(�73�D[X/D� ��dK]��ʿ:���ǑP|�()Ol� �'���O�w4�������*䉼砩���yHYT�J�hk�[��j�\���t��j9�]�e�G�#��g
���J���*��tw�{Xv�3��Y��7ݹK�-���#���T�YW0��#����՝��
�Yml�:f<UݥjM���������l��	�գ�.���Xh.�1�`���49����573�`<��#�,���a=�%�ԋ]u;<z��gF�ͽM��Y�ް�+��hl\���چ�;q�X����٩3J��Y�j�"ㄱS"�p]Y{
V6�*��b��yx �/�]��L���oIih3���If��=K��+zJ�S6�^�,���_tj���W��Db[/̼�r�ɶ��(�z��Rr��`�1����io&��i��q�8�%ᅠxNX����xj�+��5��v���U�/L�]d>)V^e����������K�,ڗ�n��8#�BKj�[t�PF��4��V��E����-�-o3&���ǧ1f����M����ik�!(޻�yJF���C3$�oU��^ї�V7ӕZ�}{}cibƪ1��-
Z����}��E�F�M-n��sx�I���#��v���~�AXRF�4�I0 V�j����F��>�2�d(S��D�� ��OɗM��B���2�,D��J���QLdڈ�^*A�M,@xb�F��n���� �)&��c�
I4@4��耼���"|� ��	�� �@@���F;�A�빼��I d�$����/�oO�Omk�������_������������FM�x�Rj���wh��`�(_ο��|�w�Ooo�u�}}}}kZ������������FI���|��x�'��5��b�I$!:|}|{|xz{|k�kZ��ֵ�������̈́�w	�d���7����
F[κ]�D��(L��� �+��C"/!	�;�v�������ؒx��:���\ō��s0�F�WP�4��`��X10���"�v����lgu\#�]��Ddb&I	�fFfS21����$H��z����e����"$��%��J�5��!����%X+�SU)3{ul�w��k�tV�n�Dh!�ޞQ�sl�3o�WiH2�y�0f�%�noK8�u�Ҥ�d�L�A�2HO��H�1�v�ԩ��u��u���-��LD��Av�W��=�� �T����ƽz]6Z�	XIa��[��Ҍ���gX�O���zP&����g>�7{�=��<>A���5��K�y6H�#$nO'3�����hh@jڳZ�R�����90o�l`I��(�ơ�;0R�Yr�|{�$2�ĭˡ@ Ju'8�޼�]j��;���$p�s&���,+�ف)8��8-nB&��+���6�@���x��L�P�x�Wɶ�vOx�e��1B��@��
R�)�u�
+*���n�Iz9
�� �0������/�s=3ԨU�*�r��x/����� �z�ɗ\ �j0���ux����K�
�W�k�Or�gO� x.k@�0{ݹ�����{  ������k=(8�.b�����⩔�%��l� `&��yN�^��8�o�����<kO��H�}:D�	۹��f4J>�L�y���T�!?�1��S���F0�x���������E/6��uc[��Ì�4-��(���b����\�o��p=�=O�]ß�_��:X]����(O�>��0��ސ,�>���5'��fNO�f��mb�X_�w~ݟ{����L�ʁf콙@ uKy�Q���>⛙d�U����KpC؏	�/�\�'�a��sC���˛�#�9vܼz�=�qIZ�MOg�k���_��S�����"c�� �@c��.88Ϟ�{��>;���=�~�����
��o�5k�D�&�q��!����2/tʩkQ�S��G.��)���ZB\�Oa(�]���23�)�\�&�L�pP,��a����^6�{z�;C	�_�̉4r�xU��/-j���=ЙqS4	��
P���rp�y�)�rw2�B��C�fdsu��='>먟98�u|EE��zo��G9R��i<:�����o�|��p������@����O2�05��	ov��Q�}�~O�?�������aыs�M�Ó�����1����xyi�rDz��{;�l���5@�y��.��]��`�$�Q	$���e��^�`����D	�P+�0O��,���G:���	db�ðm�}Ġ@6�]����f-��ãK��9��C2.��g��ʬ�����&�$bG�?�C�}|�'_���7��5���8�se���⛽v�s�&|�|��F���n�c�O���q�����Sb�2�;ڹ��iĈ� �<̳�b�����U�}�:�����η��|}�ɵ�w���67�2��gLd@��Ggf�2��h����UҔ�c��@�y�Y�7���G���s3���|�.���N�߳�-�����uL�֝���9
�A�Ok��`z�Q�K.i�٫�r�T8D��!D@Appr �� ���^��/�w}V�������ܠ+�2i��Ӂ';�����~��`|gަ]��zK����Ͻh.�R"E˦������ŗc��CF�<�-wX0����w��<U��ճ)�ؼ�D���Q�^���6H��i�]uO��Ǽ��T��7gN�h-|������W�֖�Ss��b�v$�XJy����.�ws�^���V��,�.�f{何3��*t�W>J#$Q���1^c�Z�@�2�}�����\��wuqʵ�w1�Z�L���;9�^�ypk��Gǁ�0�v!���R7%'��V8���������� �����-ִ�V�n���o����qb��ބlK���{9殰2y8Y^�4�INs�3�2�q��:.*�-�44M$��iJ5�M��Z�%2W�*T�B��/��Q\��{p��n��7��.�/�v���E�hk�큧���C�ؠi�ʒ� ����*4�?k�54��2%��QrԤ���7;[�:X��bP���ЭFS�d�J-��X �cX`|�D�qhb梾����:�4���޺��TfYE!�hX�R�0Η��0�P�;�2���-Iݝ��Ϸ�x��+�]��}C[ӺxR���fL�����
;��q'ck�:�]كp5�<�����[�L�;�gk-�U�\���`� �0 � G"1��E�Q�"��
�F�:;���_���������֟T&�8��Jz�g`3>��fn�7<p�%Ҝ���he���Ä�r��@zθ�#t1�Q�Q�
Hn6�F~n�.���A���&�����=��2�K�H�\>}`?j�����^7�H8�*�Af���ʇ�#��xD1��t��cU�F��A��IK_bel|g���C@q�#�V UL�����,��o�mI�+��Ғ�0��3Jj�/��.�w�w��/4�ӊJv�?B·|��b����ٽ�"��;�ʢ�������a�ﲂ�ˏR�@b��X�а��0,>M���º/�����m�~V��2�|�~��aw�$=��P<j;0'�w�ȿ��1h�X�*�df�I�8|��o\���&��~y��>Dg@nr�C��B��9<c�`}�M��\�ն����I컚"E�OU�'ӗ��O��Ǔ�.�XCb�#��԰/���D�������SS-�L�K�{��R�;)���Qp�@��7��=�'��7S��[����g�ʈ�72���tOߢ0e`FQ�{t��P�u�s�3�n2�.U�@5P���C(+�w�;�m���%��G	�'�ȟ�zi{�ǵ�#�@6�I�v]kO������ F��|��}�`�%�֨���c5�b��]�\�я�C�R��Ku}���풘U��*@QH�aQ�&@�7$��� ��P�W 2" w���m�~>>9���
*�!�����*>���ߜ'�5@���k����\��yWi�4+r��V��~�5+���#9���#~�}�)�?_�>�`Hc��oD�0>�Bӂ�|۵�S��'uJ�VdL��ނ�p�DȞ%jԎn���%��/�I�VQ��A�'�����{̌�r����cA ��z��Տp�X�2&����/��y��>U02�-�@�`��� ���yŕ����ol����ý��S]�@J�ɿ�WV��=�x�/��U3�9^2���z�KwB�}y��>�m!��TFD�y�
�\e�|�<��Z�>�ܮ�i��[���xǷ��eαK�F�7���p�;�gg����0��[r����ܿ� ���/mD;Q�t�D����wln��@��x�[��%..����/�8�.��fa�C#�O���jpW��t"����w1��o}(���5J�(�?y�r��L���D�k��{G4���S��x��'JE:5�܆_��ƣ��h{Gs`�h���5�+�����×y�ڟ���1XR�GFZ�g��C���^>eJ��+Ú��wv`Uef�N�6lfٙI#t��w�*�>�Ugw/l���q-ٽiˀ�Y{%M|�,��ŵ0I���쮡`U�_�f��u�~��o���""68B����@�G  �ٽ�~7�}��Z��RB��w��.7��������%8Ϡ(8��=s�n��=W}w;��{isk8�&p��%�@E�q�csckc��o~;	��
�<�p���@���-��Y�}DY����T�����|GA+�+%����&|����I��ǇҚE�˻���ƞ��\h}A���Z�0{�ճ��e���b�.�G7�`b�j�T(���Ξ[�^��r���gJ�e��e��Es��k�COpS��L�����S+���>�|q�8��k���n�ٹRy��J(���c���R:6�꿕B@�&��a{o*�_�=v�s!�w`�8Sp���^��)�I�r��*�J/-^�`Os�t&U�T0�9�����u�����o%:~w�-��,$3jz������NIN,����ph�WT�S�!�ڟM�Kxug�������tٔ�!Ђc�������Z&m��*�bo�����vvL��ߌ(���ٽzk��oc�Q����V}I�$hPK����4neEΑ�a�J_Q���S�%9Q9Q/`����u5;J����|�+�צ698��>�Y[]�pխ*�Q��i�,_JY�6��˪�8��,�����5v@�jvɢ���iA�j�xV��c���vO� Y� b ��.88�88*��]y�s�qݾ��5�k�N�TJ�	�'�Χd��
skS_R�n<��y��F��Nu���+9�e홒�)���r^��a�%�)��Т�˹���	�s���Yg�9
�m$htS��柘P��nW�`���g��#��Pi)K��`�i^)���OfIC���0��kf�	�`y	v��J�Tlѱv�S7����"A�Ϛk[��P��Gr�wf�Wv
K%2�.e��{�3�����Q���Br�k�q(=�m
dzzE�^��i�\9=c�T4nڭ�wi-��Y�g`ؕMOG��1�F��=,��������w��UÏ`ya}:M6���C����=#��qW�s؞[A{����2)YE��ِ9	7-����){D����k�/HlN[��`���ޛ��.���8�=��f?O����j��T���V�앧�<��W�-�T���,Vߤh�f}zg��y<Ku:ފn��\�YqOv��F�N�{5�]�k8w&M�S���txH&GM�O$�'�9T�~��������^Z������#��TBF��X:>f-�YRX���ԩ�xr�m��$K���EZ�b�p�j� ���͵M-����@`[P����[�݂���簬�e�p�%$�s��ܰ�f����L�%3l�u��L���z�Yɓ:n�� DC��pqq��QG;��^<���>;�'�@�0���<���;���H����àP[ҥ�,�j�C�)�J�d鯘��>��:֚�	/|�/L�\p�������>�w�-z�5�T�R!���աgj�$�yWT��t;�n��cL��RO��|�F�����6g��R$ň�e�u�u۰e0I?��}��ʾ���`eF^y6
�b!�и1N��B����uv0ۛ�ǖvf��+��V�P�/�l���ג��܉/A���i�̞���5]������ߔ������[�Ǯ{�+��ݣ[;��ʻiA«�DV��/�z���!�$.�>��<�q�_b	�Y��Td���d#b�u2k�}A����X{��=��Ւ�>��o��#"�8�ɛk�=�����@kǹT��_^O�=ۊ6%��k�]��� ��ζ�ꞃ�t��q�`>Y�Đi�L���/�>�q�$,�/�	��*W�'��^NVS�O���ΫreCvi4(��At�>J�}�t��*��������ars+��]=��B'"��ׇU������}��/�;ҟ�?�vTE���y�}R[Ͷ�?����Z6t��&}�=z�4I�L��Txثf��.�p�+�n��o[�VI�҆v|����*�l���U����t�s+8 vbr2����Ic��h�>���g!�ɠCV�f�8�q�q�>@W_��1��P2�" 7)n�?=��=֮uyK! ���!)]�k�Ї��c~��Տ�x5���q�u�"�;�x���-ٶ��]-�$�+9���m���r��ަ�����=�SM�=�*�A���\5.V�W6ʛ�=�����'�y���y�|C^cFE��<���R.�r���y6��k�S�ۯH���py�=����T��Y��"CZM?�.x��5���SV��(��f�X�;CJ� �P%x��a�K�~��y���=ò&&���DlW�U���Y�d|Y?&�����[��ӽk;4'~����'y��/�(G���y��O���~��H�M�pr��\DV��w=7LԴ�)��z%����(��B-8��ү����H�ǅ��]o_�?��V#��a��L�	�)������k��?r/�w��8��T��&��/��_�~�9��μ�6��"IH� r��8�������ώW�Oh�:G�S��{	�m���W\���9�s�{*We�e(뿉���(h@��$5��U g����)>9=���4���a��?R��Be�)}I���)��jՊ�h:{�wFf/������]T�Pm�V���o۽��^�$T��,��-�f�i�D2��6l���s�	����t�Fh�LtŅ�/1:��4��GT�LN�n�:�g����e#܈�{�`���g\7����� �8(8�⠹ ������J1]ݲ���<��dҞ�A�2��9�}kn@c�݌X�������&|�;h�l����:�
�?|��N�+}��g��V&�s��~<���Y˺�iz~���3���-T�����$n�ׄP&{�s���2�'�8/����&d�&���ʜ���zg��~���]�c��*���C�t\u�k����~>�|�w���l�kW*r�زX�d]�Oo�z}�7�@�V�¢�q��h���{'�$S+%Z�y��%��y�7�_ýSՐ	��.�>��_+���T-aaS�?[�;	��#r������f�_s7�\�0I]����t�>��=��e>�w�U���n��ln٨j��g���[h6���l��tD���Cz窹�ߣgH�wP��|��xb�/)w!!�EEe�48h���� �f���3���;���Ĕ>=�5N�Vr�ﲅ�Z��L��8'�����\��Ow�3������1�6�Al�%=�ܟ��i��m#40W�@ D@�ҿ8�z��eP��[��W�Q�V3�-��i�Ҡ&�uӌ>,�e��gN�ś�)��b	U����@F�9���k���|�u�ɻo%WL����hb�)s����n�m�c��LPܜ�Cm]��-���8m:�]�k3ك��J�*;p�\؍pz/��r�ά���#{w�=K��m�5���B���m�b��.���r�b����.�s�;թ�]SCd^Fqq�Yý#�W�m�c&fMZz�a�d�ܻ讶��X�"w�Ǟ:`��a����u���q��,3�\ew$��뭭�]��ҹ���^�:�-	ӯ$�f����o�{��h��W�%Sb�	j�[ys^k��"�}��g:�Gf��U�c�Q��
��\{s�e��g`Ơ�z��wگ��]<�͛�_��V�"j���3z�xy��"f���[�Z/�\KnX���㽧�Dmigsg�\�����\h)gt9��˂��H��0%)C�v���,6�(ok�Kk�ue�t���v��1��yK�M[|�px��u�V�M)���h��򄇕2W[���
����:����֎�wC�����M�W��9��-��Z�i�f�FL�W<����d��K����!�0��)yP�μ�A�<��X�b�b�Z�Y利t�XZ����[���{�_���Y���y"�U#"����t�y�t�U�xt$���g�����H���&�b��pnu�'�B�L�X*N��77��ġ�`�L�����՚{�y1�9��m������KEr%�n�lb�[�̸�w�sV��Cm�+������u�ӈ!o�Y�[k.N��H��s6Y�A���)=����GB�%�b{m)	lcn�&Û9`�y��S�M�]�g�NB���a�b��֧�77�J��:z]����l�sS�.u��vaů���.��Ц�S�is��R���N���oCx�Q���4)r#�@���T\�+�]�*���4[�R�Zv�K��"ʽA������t��*�ӓe:1ہ�S"��=��]lڒ��m-#�Cp��5{�op3����م"��K���m��g��]ڎ�Rr�uP����.��i�=z��*X��3cӪ=��M��X9��ùic�+n��0����L�ᵅ�}����׽"I
���漶��%U�ԁ�4w^�d���e�}2�rR9���+�� 0�R!Y�����t���Oa�u�2�qt��t��1�S�X�����ٕ�=Z����c�Ӹ��0WI��,Oj~4������Hf(�O��ԔI�	���ֺ����׆��}kZׇ��|�7��H�6�O�����Z1�(�-��Ӷ���!�>�>��:��ֵ�k_Zֺ�����I �����H��Q�E%��]�}n� W�<�2��wO��n�=�5�kZ��ֵ��ק����~���0\�_���_�Y��^-	F(&X�@I�.�
";��=uJH�#
#O��7���٣DX������A��-������&��ͽ�w{^d�[hF�ȑd��咒Io�D�}����:C�,A���(l$F4Y�v�j1�J��\�Q&�,��%�;�c	�Ch(� 1��Z$�Ѡ�&��f�F(��Ъ��ԫWL����:n�u�W&^_=�$�w�����}�F�0"�[�A@��Cd]�&^.���^�W�?#��� &88�����$�nX���!�h���^1���	@��nʣ��~���������t��U��1wB��{m�Hp�{�F�!||�si|���@uuAl�qv��0�_-ҽ+KK����'�Kq���67kӾ3�@ȑ�ɆJN��# B������]{IN"��oa�:��~+r:��wBOm~��V�ǵ輱�`0!�0�yi@�����OcS
�x����U3}s��f�4��aM�W�bq�q���\&�����;օ��#��Ĥ�ɬ���WY���^�����Y9��7cmRa^$�i=ʆe�^������+��n��l��{�P�x��7R{f�ḭl/Gz�Vќ]"�6*yEc�n��+u�����ذE�Jlz�
�OV7B_mvZgizt��*�<�	�r��V�ս�ۀ��`��Ǧ��B���3^�=ٻw��wk��e[ZY\,>!��C�������D$��n=�"�֞�����l��Z*(��Cg�Cit�p��8�n]5�y�Lpbˋ�2�z�ۅ����6YPՏ�L��lO�ʂ ���3��E\wJBp�(�e�*����2���� Mt�Ty-�(s ���+|����!�I�	�H���D�H$.������ٺ"�X�DC�����+WJ�fㇺ�(k��3%���Y�0��Ǖlv�����wz��l�=2��|?#�.88*c��H�)���q��Ǽ�^�pu��:�QiX͑��v}J*�p*�@��>�v�0c�Lͬ(�;3�I��ȕ2�{��<�N=�y���0ޕc�Sj�_�����4��J%��eL9��;1{y��r��?Y�嶰
�,�l�������,��z)��O0>^w�e=u�x�3�ٝ�;ms�܂�b��0�^��;>��S2�y2�}�W>0�U<��yn�+�>z�S1S�8�����_�O���如@��">d<�\9{@~Z�ƶ�"U\�pqA�wǝ��f�g��Y�I�-�.��^��ޮw-����0�%ưB�a�~(��X��xêj�"��6a��[|�����*�"]_?u�Oګ�cL��&=�'��Ϙ�8~�'����S6H���Tv �]2%���I�����I�W�;#�:�F��6~��c�E&��o�8��4\rO�������Ҋc@�p�O����mz�����3��{��ŤkN�旾���|�vܦ�&O�2�3\������2A­�J�'z8e�z"�br]�L�_�7Qe�[�q����X���Z�Ӗ��[ѭ#2�X�W(�[\��k���?���R�j�̔�ܒ��ن�����⫊�rs�mi�����5;1
}P���SVhn�;C�M�f��L��g�,��uS|A�W�N���T��l��2f%�Z�� G���  (A�"�<������{�o�](��OH���e���OB�0g�("�w�z�5��0v>݀99Q�����s!��$pġ��>
p�i1P��J80��-�G�ܲUZ��&6g���zҭ�7��;zy���V�.���>��94<���2>�V�Wۨn�n3�6��Uޔ���x��1�br80��|w�Ag����RWNȤ�����e�z��V����/(}n���.aw	�v��C�'��}ʋ
�Q���[Ƽt�>N\K��i���F��nkz��(;,$��:}q���pu�9\���{�V����ܕ����n���%UB�J��)Z@H�(��'"��<�Q<Dـ��Aa�A�9�{ȉOÂfסz�OCc��9s��s�֦}�r/=0���A,a�}������#�[�G�e�qRA� i�D
2���W��A�FQ8��0�x��ˬ1�]]��.Y��Qi���cϣ.A��X��;r�D����,���@�xuR�k�qxL�{�kO��L���R�W:��v����a$�r�¸>5=�Dh����j�k3�&�E��z�����)o�w��؂���PI�Vm}�w!��|�G��ӛK���H6�r����A�1�!Z��%r�㏵�κ��ԭ��m=�؆#31oXގF�C#c8��%ݷ2�nxv"�/�⁎ 8��
 �N��ι�a�K�gk��xl�pЪ9=�h_�8�t�OuW,H?�I�VQve���z����jo��K�gA
�K�|{�&D��bO�� i���=�U���s�UR0�eT9��5x����3�|`�$����̾�Z�<��KmL�ؼ;��.2 y�-o��WK��E�A���ixkUd^�AО�6 U~d^�6Er.s%'�9n�*��̞�/����Çs@ݠ��(�bɵ �(��.0s.���u}Sfi�[]w4��I���+z|�_���L���WB���߾@R�8�6=t�_��	�rZ���r:���aK:���R,�ĐHz���/b���:��zT}��c��֏��r�Si�^���v󪪸�}Z�3����jϹ`�q\��.�0^��������dz"0�F%�_I�fsC��r�ߏ���%14�N��R�TEȹ�=��r�f�|��K(��
�M��TY��cu�V��=�PnU5�����u	=R9X~�u�,�T>G�_�'��#���<�!�ð�[|Md3��L�9���w��)�19&���s�+�C��v�ॲ��o֫�;:�r�U�:
�c�ՠβ���m�E�D$6q�ԦQ\4�\D��Sh�8Խ�R���u������m�!/������
��	?�W����q���({�������q�-��hV���L)����j.E=��'���tT��L'��[�%������BU��|w����R`�_D���T:��s�^vF{��6g�&���.���������>u�HP΀�ǽ8�8i��vMs,j.�Bn집\�B����/n��ȟy�s�F��u���Ν��2o�`�y�8�SFKHܩ<��nQ��c�z���bK�Z���ן?^����r���/ЗTy_/֪W���N��qCrQykU�Gt&[��܄m<ԷF��#P������j��\}-�>�R��T�@9%8��St��9�)�v�:z�5�g	�c<�a���;�}�?�>6�`��(�0��ي���)v����&��3 쫻�:��w�T�����]'�	=��a>F�Z�^��0�f�!�J9nVzKߪA��z��k�fxd�w50�	KǋV���N�T7�{d&О�+�Ąn4|��G�;��/w����;��{�L3g<�ݚ�mW0�LR���s�3������+�}?o��U�_F|F��FͰ���A	?,o��Ԏ��1� ��Y3�ӻ�6����1 �a�T)G�S����z��k��:^7�*XC���ǟqm������VU���el�ó+4�=�&���0j[C��/�p\pqG \;�^�>/_�:���1��_jFeQ�Q78fm�4]�3ϳ'��<'6��کYg���w��GI!^�짦zxc��`0'��x*n{�Ī�F�՚���Lߗ�6���j�m�hx5��i�F0�
��S�/��7R�����>��w5�A��H��7o�C��3���8�5�z81�_]�+p��l*a��"��0'�t&�q��3^`:��Sw���e��kީ�(Jk�xdsu�^�bye
F3Ê��b/�|�/���bWs����\������lgHɏ�^g	��O��L9�9_�י��n������,ҥ=�Δ�q҇� �=n����pEџO�W'Y�˞��s�4�u��@s*��ξ�%ob�g����pƢ1�#�����5��e�e�O$�'��9?u�_i)��
�#nM����lw�m�J>����l�fx|ᅁ��Q#��6D����w;�'[�����c)[b���H=mp���1����������p���B�C��f.����#��r�I�Vv'p�R��]��JY�[�T_5���O;(��u��iHKk�˔鲹;���h`=�׻V*UѲi%H���,HML" "3oy3b����>�a6���q{����r�Q��MG����*͕�_F���kXtù���J��\�jR�St�3Q���(H�A�R��Y�&���  P�(��@@�2m/w��n{Ǔ8�(zG\�%��ꋼ����r���΀�v1�Gʒc��s����)+������ۃ�d���G���;;E����.�����q^iWr0��^�`S��X�2�K�M��o78���a@|e�r��kȵ�&z����Y��b@ǫ)-H܊��r�TC�قO#= ��
`��b
G�)��s�J<�b�&�\���uę���ߥ�菟���s<Y�f��#�����Ǧ0K>)'8;9zI	$]��BC���r��P��T�����jƏc�~赸�ڻQޭr��?2|lJ�JZ�Y)�pa����Gǹ34���S*F�r۩!��ݰ���K		T�*58�#��/6�ӏާ���/�3��+��:e�b�;��N�cѯM-[�z���u.��9��e�gyP�@�E\6�ׇ�Ӣ�����
W���O�p{Pr�L��p�`�����ό[5s���'�}��x75vD�׻��^���/�-��:���W�UtCƿ'f|�X�an����g-xE���p�1-��ܦ����RŚ$���=4eE�>2��nȓϗ�J\W�����Yi�����4ӏx����w \W^#�t���(�QK��nt��,�ї���+w�#j�(�q���%�x�[�4b\N\G�f	sK�,����K�7>D<~G1��O/G]��_���<3�s�Xj<��@:V�����C��Ƹ��4S��.8_b������[�;�q�4�<H�U��`/�����+�=�M{�P��Y��!��@������&����N8�U����̻�ȥ]���_|��K&<�\A�~��XmU#��ht[�t�4�0#���`܂�/^*/����ϥ��۪f�I0�Y�9ܩ긓w�F��}�r=|�|�'�=N7�[I�B�g���n�>�^�>;�O�%�ʋ��q/7ׇt�*W����$p��M���5Lkײ��{3۵˘��N��=L#/*���5�[����Ş�ۭd,I"h�"��i��c���kй�����ٮt�����B���l]5H\n��{�b���Q z�G�d�� 
�:Q����/P˓7t�z���h�2�U�t�o�\.�~�`��,Е��|d$0��ҋ��4�Z�&r}��Rw�@ ��y���i�d7<Gc��7fyW�h�n(��`=�ukƊ�0ч�%�9?��يW7v�TS��f���w]/��]���v� ԫV�w(���EN�6�����EoZ�Ԋ�/=��7^ͯ����P=��ݺ�:�۸����mrz���MWp�p�N�u��3]�+�qb��$�Sh
�w���
�
� ���nwmשʯ|C����݌�=�*[���w@���.���|�T�L���k��NT�Uf>��;Y��G�*������y}�ڇ*N
���^�����P�Rǟ/�ڣ��6o����9�lY\�e �X����Sܑ�ya���m�S2�ze���C|�#�Hn[;<˿]a��7hko.��y0Zr鯫�G�!wa��Hi�Vx�������K��9�V>L0��-���(jRe����ԇx��Ϗ_}"{D�|E�r\b�R�Ҳ���0�?�_EԾy�:�5El�]�Kf5A9н�$vG2i}�Ľ�<�ܤ7���:�q�g�k�1��1���趥i�����ak5_o�g=8v�˪5�4�j�t�-�x	���\���P�آ��E��2�|W������`���+<&Hz|����;q��U���I簔Sr~�-�ݩ�m}��9t׫g�۷U����a*,x!e��dx�����@�n@��ь!�^���z��S���N]�m&��Qq>/.�7!���o�6ע6��/)��H' �%jBڮ`�g�|f�g1\��Wj��b�jx�ث��V.��;�\L�P���	��ʾ��Q�u[���[/tQ���rU@+��h@�� ҳH* 0	>�(�VG�N��&�nf7:���|J��o�q��r����C0��%�h/*u���Wfz��I�0?���
��B	�J!�����w�>��~Z�������όꤘ�|6�����+�*F�vբ��vzX̛�[lv8ׂ�p�3��.��э�qDO޹ƵY��CC�B_Rf�w9�(���]5Y+E���g��1�����q͵9�ð-���;��ս�)���	�HgW���׵�@j��-}k����;!�o�]r��VH����>ֈ&��Ob�3-t�b��q����s̤�έݮV��)<���,���A��`}���7v-����9@A��%�0^:�<�����n��<>��ZC	ʓ�a��N�~�k�dJ�Tlѱv�xm�[�8�����bkx�kv�qt4Z��{k���S�%;H|rji=ˈ-[���+ދ�Ͳ�����S�۳cŅ����B��*JV8z��'�1P�^��C3O	�,t&ξѺ��!��.����5�q���B9�xe��=c��V~=Y�������)�͍�1ǵPܵr��5�n�y��K_�y��Ɨ�$�0���Ja�^�]B�ѳ���q<�r[c��%�r������&�[�3/V�@��;wI%z�q��P��Z� g�����[�7�o�V�fcDxr��#��R����oi*Sz�*�ol�ū��ɵ��	���рδ�j���7��n"���9HԒt[�z#��C۱���ۻ��9;7����yj����L�;��n'��ā�(\K�<�oT��M��L�]Xka��|.W����v�7�Zm��^���Ӊ�Y�����ﯔ보RgT���l��o;[[�:���Y�O�}O�P��1�US��#�j��R�h���1n�U�����ݣ���Q��<A3�˂:��䢱.��H���ݺۭꙙ����+:�"�!���]˯�Ƣ�X�JR#̹Is�n�~��Gw�3�-�Rs�b�a�.��՛"�[��q4Ei�����{]��3M8���_ch�e9�Mv7˦f�����k-λr@%^�Ǌ�[b�+�v�`E���e���-��L>��3٠��l�Oh0��d�N�&Z�~���;0�%�zЮ����~#.$*v�[}u��S-E�yJy�2�-l�ͭ��L�-��M���eҢʗtGTUmw!�k�J͵�����)���ܽ�j�o`��q�����|��>Y�WE
����܂{��R�8LV�,+�(/*L�#�=$y�IGA(A�8�&�N���̷^4U��Fp�n��`0���`�Ƒ+Ұ�-?Z]o����;V[�j�ہ�/.� 	�C��*�4�J�8KhDkFKU�Ɠ.OEݝdVtu�=Tnqw�� -�f���nQ �3���_:
}x:��ۘ�v��]��ڡ�Y]i��ћuWm"K�r"��z�.1�!j��v���R>/�+�ӛEM~��;k4D�pu����qc��B�I�A�Ca�����U��L��9*��܃bN-��w�"�KCj7O �"�"��1*��T�A����o�٤�7��"�a�#kjt�{y� !pWXWt{qvt�ذ([[7TW�4��Nǭwm�!=�R�^�+/��F /�agb�F�P�]=��F�Xk^%+]Jr��u+��{;�}[.+��0D��[��Μ8�NsŎ`�u�%U�:-u�Lk�OQ:�` �α�@����݆G&ʼ��;3�Q,�����b�wQ�&��=b���)wK�x�]G/�9վ�/ҹc�S�@�d2��P�W}�o�v�(j<�9��W�r�^�y{j����u)��كb�P�\�1 ���J�Y��������Y̷ٵ�"�[�<�,Mn(�Y,�6�ʱ֧Wgv`��`�Q�ou.��WyV�a��ظ�:��7�[���{��T�u^�r���mf��9�nwv���0��>��R��hq�4�D�����>�	� A�f��D�LAd�X,��R$�2D�'�T�AUa�L��$ JKn� BD�L�!A M�i[q�TD��$�(y���A�L`���s����կ�~4X�I�.FM�-��]��!$Y������ק�Ƶ�-k_���������2:HB$I6)1�-�;��>����������Zז����k]}k�����F�A�_}uy��F/ƹ��6�O���w���Ƿ�Ƶ�-k_Z�Z����x#F��~-�b�ō	�zW,ZI(�K�vŢ,�ur'�4Qh�>6��x��O��l�MF��}\,G�u*+~/�x�&��h���a�6��g�k��F��r6(�V���m%X�
5%�l^����nyk�Q�MW/��Ω�n��m�k�^�,X��QRh�أԮ��6�UhC�&����z�K6x��U��]|�1�݅Kb��ڷ3'l~.�l����}u�5D%�^8�u�'�i[p7��*(*L���F(�$��28BB�B (9�V�z����l��|i&����e,qq^cEk�#:_|���9;�������ݧ�huo��)ݩ��*�8+�|���c�}#)����v}<����BM瑆%?0�����<����V�ݤ�N=���� �(]�kw�:�Vf,s��q���{"~�ߧ�~V.��A䥽~����9/C�8p�Ns��|�?Tv�5��!'|����`�´/��ґ~�8�C��O]���*y���@����I�]5r���=���>���&6�@x�Ba�[tLmN�rcV�ۓX���R�	�-�.v�qiL�{�Ĥ�O�q�n�������`����L��Y��x��8�4u	�a�=�v��jH�}*�_ΏV�Ӄ������ʽ kQ�	�Y�ɉ�l��Tl�p�OA��'F��p}�s�R�,�`��}������E�[��'��ᡨ��ۘ�wmd,��i�W��Q�'M���cI�Z�0?'�i�K�wP��Z�b�wQ�֮�2v��v�����,������T���E�A1�e�嵲��_QQ�H*fK�����+��N��)�� +�V�=����~4Ŷ790.#�HTr�HLd��Һ����l[�J���A\*��k'��*�륍�g9t�WP���W]B]��]��LDl�`G:ŭ>%�ŀo:)���l쭚z�<~��!B�vs�zwp��Y�g���[��H�R�R]��E�-�ׇTx]P2>�q�D�W���?�i�X @��4�ػ�|��ON0�w,��^��9���K�6Ymy��m��f�u��ՑQ!��a㉞vF����!�p�7q������<����g��5Dt��y�x�{:iu���P�HØ��������H���ߣ`�pK�-~S��̓79�f����I�
sB���Ơ^��вƌd
!�!m]q`�c�m��AA�U�g卣/���n�=�{ˤQ�響�W;Q�5�k��c�,����=C���N��w�V7�*�?�� �۸n�]'9Q��N�˸1��R�gu���o��������L�ȇd���-���$VAK({�Uȝz�r�_O��ofy�d�0#a�\P��#u��Ov�ݙF��ieL;��C�;;-}�O���^�j{H��Tw=�C�$/��l��GKY=�}V��?���/�W�a��d���:^="c�*��^j`K���V=�/�y�9>�ء"��֚�W�H��-��vk-�Asj�f�]W-Rw��,w���K��1���ⴈ�n^� N˦ck/J���fX�#[�m��(*�*�g��m�e`:����N���ҹ�YRa������	�o�#��B��B!
 ͥ�]�v�G�*1�A� ��XCཪZ?.�o���P��Կ.�B���.c���_���j������_�:f�S������
�����j�� (	G�_�,�,�[=��p���V�V��0��^e���Ĩ�?8S�a �2�-(�����kw���Q}X��z`cr��n��LJzC�i(fo4E�{g3�%߫����uFvI�;p*���}�wx�`����!��*���������u�I�w@�ǔ;`O�q�s��%��4m�c�}��)=�.A&4s�	�Xa��%�,!�렧�ɨyu�źw_@C�И�������7���}y�`���Ρ��DS�>��͟r��]x�R���]�
zD����l�Es`�"�}�z��]Z�:9�~BCOUz�D73�����t��~�n}���}<b�X��O!_�������v�Ҳ�s Л���T69�� k[�o�s��6vP�������w�-��D��� ��O܅�;##�쾨��,�}��Ĉ���WW�}m��z/�!q䩻��K�,$�'L*i��s���.�B9n���9�S.^�*��+�(!��~@�}><S��ͽ{2��[D�+l��Q����U�un8��؄���0Ql�Y%D����ƹ�8.���"�!����:�.o��IĈt��Y <�X�@&r��E�&��^Es���[�5��Ow���{y��n{���d}�vxd5�n,
�C^yᙺEd��ʓ�iE7'�`sV�p��lY
Rm���z���	�-s�{ni=;�/ޛ�d�0g��^�ځ���aB�J/-���s4�����f�Kt�Y~5uCu�*�������>�Hc- B"I�C��2�9���#i���[�fܴRXΤ��ˍ��W0��&5t�O��Ǝ�'�
�?	��p���p9����2�l��\E�a�	i�"��$�BFx���R�����mύn�¤k��z&7z;����/�vզ�T�o&�|�ͷ5)�i���1��)�bJ�i�7�Bj�z�f����n��I���? �<`����laُ>�v�=ϯ[�0��%>�36y*f���V1j͵hN�Y�6l)e��������|��H/�"�Y��ﱒ0]�*Fd�^]���U�`�Ol6��x`n�2�#p;7N���	�8s8���*�Uj�h�P���{lқ���qQ ��a:δ4�렙QDR�C\SEō/w �Hj̴TE�u ��9W`�[���/`YmY��^�"�fV`*2�"�x��X�:�X�mn퐕��X&۷�-��5�3_y�	'\��K'�c�e#��[� (\�H��X���~b�#��"b�7�����J� �Z��yv}�>)���m<�^���r�57����i�W������SČX ݮ..擙2����C�J�1���l	���>T-�v87Z�i*[P�?7d`�t~�eX����]�S{�/�]���*�u�s�z��&�|��	�FGw��v*��B׻soV��2!Cw:3Qd�c����2o̍���Etk>|�%��s��q��Ew��O9ʪJ�7���Vl���P|;���_+F�vW�HM��˜/ɢn��+���,��J�Q�M�ݴi�زᮢ�@P-ߘc;h`����p�����1A���Uy=�����ڞn���a�ИA���$>�n��v_p����LĎ>{�ce�Kڙ��N2<:V���L�%�Or����<֚�$��0�%Ʋ5U�x��|�;�ϔ�5�̀
���0��CO��4�����u}*���u^� ���r��J��%P��x&��٩&��p�=O�p�Ϊb[L�n݃~pOGk��I�^�\S&i��ߟ����������*�6�X�m:���Y��!t-�b���v�?���� ���:�i��xB��3s*:��,��R�sn������˅b����N��&�)J�WY4]��gטE�K�� �J�����~�y�G߅�ACG�A��ܥ�K�$��^�g����^7�l�ӯO�S:z�=�9� �&��w�ʹa���}�{3��c�Lh}�C^9�ye�M�>O�}[D�K]M��½-�p��^�{����	�_�P����a2'�{�k�m�(��U���Yf�107����T.{� #JY���S�0ju$M�ۏ9�Nc���꿾���1��}dM��;[�z����n�J`�_A�p��Rs��|]&o��߳�|N�t���v�lv�=�l5n���|����G!��sP�YA�ٳ�����{[
�����ӕI6l����NA��$!e�an��O+#�s�F�F�͜�y��ND��ݿ~��l�h�L������b�4��-�sa2.��>�W{"`ec��cѨd�o�ش#��v��j�uH�S~\��_����U�q���Ѵ����B�	|EbY*��c�έ,էV��u	�{P}4���{�l�ܫ��� �9��p/65OT���*��~�[�j�˄`^�ܧT�Z�xMM.���[9z)���i,2�)f,�o��!�vn�����qNʴ{"�<-=y�ϙ��h�f>X�˛zķ�+�$Û�+�ln�Ad�%u,ǼV<�������<+�¼�M���18`#_X.�IƙS��Q˭��]�X)F%m�zh(�q�}*��u�����D����
2�H;	���{t�ٽt#4�pE����2~��_fgnxz�'��"��ǃ{���>z_���X�a�Vc���#��Ws�Nhv�?�WO�u��Hty4�Z�D8�c�]�Z�Tȟ.�aįW�զ�Q���f��軜�Í����z򀗵w�O}s�^v�q���/��y�;'��%��XZ�]�EJfi;��(��(���<�V���>�S:�_m�#�.���T��h|t�j�˵mAm4�7_>v�	O4��\������s4¼S@Z��М�>z�{�5�C�v�e��9�'"�r���^犚����`���3b�����z����}�$=��#]���������]�n{��iv�2%!��|��7��p��mCvRz��xf��|�'����u.�3��� Xx	1Oy��W#y�q鲙���l�PѮ����῕��D�Z���ϩ
���-d��:�{w�Z���32>�r���d��.�{rq�nQVc�7�'L��O�����}��㷏.Ċ�s�c�huP?!<<(>27\ֹfp��XO�2�!�fv�\�WD�}�u���k�����{倣�q	�jm3���xt����^���f<��~�F~�{��7����Bʵ�����r�4[:)ۺ���:�3�럆�@�~�cs=�������YRJ���qp���7EPO�>i������Q��SWu��N�X��;�bXqb�%�:�[�������H����Y#��@�\<��<p���:�Xbn���J�~i���;1:$]Q� ,|wV��#�|3ݍ��M�8�ȶ��ݜh�a=\O[���G9 ����c.p����1Z������Q�.G���8n���{�P}�Og�����{*��Q������vcO+Xy�y�'��!���W�΁{��W�r���QM���`� 5<4�A��*F��x�rǙd��j�H&Tj'����|�U����+�`�ճ�Nuk��6�W`�>��M)=�sڀ���?Wo�ȞM ��b���!q��je������Q=o}�Դ
��ͳ��Y
�?�p=ԘM�%���@H�����?���!���Θ��w��}�F:�����E�TbJqA#<^�BOm}PXO���W����|Oc�ܪ�O��[{&�߅�amf���!ܝ����c���Z�����nE}L����h����+R����Jw|�G�

9YP%�0�C|n���3Fr����=Y���Q]0cPX4匽����Ö:A{�>�1�d��T�/�;=ٽ�ܔ�F�ƈ@Ph2�R���Ѥ�	���k����D͛�z�랝����VЙ,���1���'ԢO�|v=���dR٭r�F%)�8[3ch���zl���9���ﶹ���O� �/��M孹d��c
�Cf���9�%�t\��㜼�[�ݝ��d);� b��)I��>R��(:v@�$���ݕ�?}8��1|��GxV�{�;�CP���U�=�*S;h����U����X��3JM˟�ʋE�F�r��ն{o��jf�i�U!
�k�7`:j3���:����pi��1㶱����x�Ncb�����&nE�����dm]^JV=48͜�8���~�>x4NHx���!�_Gi��"Z��A�j��� L��������b�\���)�y���sN��������:%�>��{k��1	OHvA�SxtcC�Z������e�ͱH8|�l�d�2���f��w�Ә�j��H�iH"�|��6+�h�F}����_�����o&��V9[�Sa]��}�W�����]���,/��R�t�e�����{���x��3���Ʒ�3������$Ӻ{�Q6֝�>�}9c宛g#5���Ye)8eY2���l�0�A"�D!�3E������҄Q%�Z�}������*��%tк¬�٪rC%J�k���>;[
�Xy6cfӭ�M�w�J3,��g�7��o0MR���-Z��lR~a}�;Wa�J�<F��?�m"�>Dўb�t�<6q�q8��M]�"z�V��qI�I뜱�ˌt9b9Ĵ����gE���:��]Yz�q��3�MM$Agg�<��0-Cs��z��_F�E	�q`��a�-�=�����0�v�y<ʈ��5�A}��L�6�O�H���Et$�/~�ț�9���GF��gj�#+���#dk��q}�
3�>(�\p4O�LW΋���{S�^������xCg5�mX��z��	���Nxł�ֽ��c_�+�}�P�yd�lo�;��ş�g�ﺶF'�۫�j������ �{t;4kl4\㔧��G�?'�i��b1\�^�=�bK_�K>�d7�>�o[��LDl}�I
J�hՂ�`	K^���3t|�3�nO�f.�cq#��ۡ鸽Kսu����*�4����.�!t>=��Ro��b Si�Y����= {��8�v߷9���L�� 5��ޮj����y�u
���<wN�C�e{:�-v
�����;���v�E�j���d�eYY�t���7]N�Uӭ�>z��C]u��'�C2�WGn�陕t����zs��V�}�ͽ�΄1���V���:�(:]��<��-ּ�!43J�$v_p�⡥o��~��)��x��ּ)�Gg)�sc�ws��lv��������IZ�� P֒�7%��[z�x��
�u+l;U�v r�˶(3.�3���w������>�)8f�\ 8_�K�v��:'�9���]Z���'j	�gf��+���Za�|�g:�l�M��N�Zc{�R���پd*W���K9�)�̍m�q��ɳ8r��9�bmJ�]B^�#��ڄfk�VPX4EV+�;l�����a�� HsmQQ���wWvt��Ǯb�t�ޠ����
�Q�
���Xtδcf���oz�K;q��Wq�mi;+�"a���-Xڑ7..+K�"�6�A� U{�]oHU�\2�UvJ"�;WpӨ�1���_Uqhn��hi�̵�^����1f��r���h�b�!a^=�y���,��r���Y���j��Ďg,�� Qtר�Ꝏ��t���T��O{V޻[|7���k��C��W@����W��R��v��/uɎH-
���U��y܁Y�ҍʹ�^sX���R�,WJ���e��]Al�ʍ9c�ժLY���4M���SQϡ�W�}F���E�J�I��ܘ��]�k�;V_"�/����)q�p|�\��$wR97�N��S���3J1[��ص�w\˖�vYG ����<�oW�B]�R��9��a܊b��Z-rb!���P՞V8���n.�,v��ڭ��"�,�g�i�\�o2'��*�V>���[b�ή�%�E�"�)�A��b�9z6�E����N+�����\��WL*E�w�hl��:s����t/Sum.��7��d��1�=�K�k9d��S�7��+^�R��J�|��T�ʴ���U��9������!:�\����+7i>s'h��eѵ�jOͣj"o@�J��g �w�%��~�N�Or������諫�tB���g^t�E��S�vS�Ov�PZ;���������Y�oe�Y)wwWged�p��9%�r�n��/5@�8�ci��${�C��Y@�J�|>kn+�U��w=��t��Y�ś0�ާ�*��{+�\:<k+�a{��38q���u:P[D$�SZic�"�{6�Y��{˄�5��Yi��0d/��� �\ �=���F��$�YE��;r�j|��)Nޒ_f�6uϥ���݃�M���u�K�]�I����I �*4P�v�F�0�22�><��==�>��zk_Z�_�����)�U��m͍d�鶼W�c\C��BO_^���z{|kZצ�����q�����̈́dHA8�D��CF�[�m�clXԄ�F3�o/���=>>5�k�Z�����>�===:�ؤ��$�9Q��.PjƬcE�Z1F��V��TlF*��YnT[D[_�v��0�[EDm��ƾ��[��
�W���������騣IXB��WMM�Z����^�]���^�z�u������r�-����;U䨫�W+I�b���ơ~v��;m��b�׊�
�(͙�+�z�]�{����mAst�j�wC7*��۷�y�W��%�6[���!���"gLl| �a��/pgj�{*q�=ol�;"��0��o�a0����d}�_�P��	�ј}T��̾�w�g�G1NW�$�H{�lT�]j�?�D����	#|��ȸƗn�7�l�YC�F�X�;�4��A�[����f�\�P��-�g5a\��L|�S�R��O=�֓�]���9vo?��{c���$��:�c�E7w)�}��f��c!迮��[Jl��7H:^�U��]���`��`=4􍴴�c�]<����u��s�k�i�b=�1=y�<�i�=�Vݥ��
:�w����G6àۗ9�=�rܜ��r�2�[�����ѷ�Bz`�F,s��_�U֫��.�/!�Q�\5	i��<^w�B��{S�jG7C����ؖ�R�YX�宍�83E�<ܢ��3�	�ֆA��;�T@�~�۱�Z��O8��}LUS�+w<w:i�F	y�򩁖6-�@�`��B5� �^| =.!��{���ӏ����E�s&f��';<	��Oʶ$g�AL����C�1�p�48wd#��w�]�Ӷ�O���1E�&5%�K�%��n5K=�V����N��ƻR[:��9�s�h�H�[�-�J��
\�<v�y�s���h���i�S�͞�v1
"�n�!o	~���>��k��Q�'���Ӣ�Vg����φ @�A�"��^z�����᚝r��dΪ��]?��QM�YiU��O�c�N�̇%��#ٍ�ɬ���:o��t�C��
ߡ� ��d�6<��P&%=ɧ�C43 pE>ό�\����^��`�{�}��H�ĉ
R32Ħ����3��B5�=��&�e66�Q�.�����;���^H��O3joC�8M� ����zf��� �t��Y�a\͞�d��3QM�Г�!��13��6��&����s��k���݁@�t�ެ(X]�Z�n�������{e�dN�W�>�E�����-mY�İ��ʒU��q>���Zᛇ8�	�1���J�j��^%oY�E?r��o� >B��]2Wʅu�Raޫ��-��`�.}Ol�!EKk@�t35��n������T6�+��!u�͏�K鈞~�cr��)s�gX7�+m�ڕu]��C�f坮��h���݅,//r��R��kPѾ�� ,�&��\�Q!�����^L���;u���L��.><(�|������%�nT�z���t�lK
�h�{�Țu��@���>s<G�/��N��`R��:�`�\ή�_qG�0��z��x5�h�j&P��9�[�1�YAr��X2�Ar���-�x);�B��S�tQ}��>t�k��V-�Mz�j5�ƇVp�n�;k Hd&L��$% �`�d������ũ�9p�u���s׸���Fh���6�J��Yc��ڨJ�[Q'�B�[V���
`imV��$�X=*z)����w?�ݿK08�l0=�ҘHy���a�ͥ�ӎ�Ŏ~A��23�OP�.9=�.������ j긮�~AræG�$��}j�|ٖ�!r�Jq�&-嫤��jz�}���?r�]s���/�8p�Z�����q��C[�5Gv��9���'�>2���4N�=##���
c��S���	X��>��}�iΖ�Y�;&�pM�S�g26C2	��~�uyq�Y`}�� (�>��>:��tn�s�F�nf�t�w�DS0-�<���nUP��ϔ�<���xk�,�)����+j�;=��=��Pi �/�zZ#E<S�~��	����hN �������|%�4EW�O[j��u�{��[��G�����u;�uH��Iz�~w+ŕ"��ܱ���qZ*9K�����4}��p���{���5�m���{28�]J
�6pS��?U8D1iB��v�|q����ɻ�E��p�s�U�:��.�*������]��Y�����T�9����`���e
����uk���ݓ��ԍ�VʾK��������Ni�z;7+/�c5��W+oWT�ƾ�Dn����?�y����[������7��@M�9k����ܟ>��h���بW=�-��Z��U>���}��g8�}*�3@(��Q�!&�6;�q�3�ɿ�ӻ�ys���y����|ûq�����u�"�"��j��SJ�r��]��]��'r��@��������-��a��|��E.�m��靖���(+�|�B	�;��-��~��l=':u��c���w���/ ��~a`�����S*�4
un�]י����8\{#4#�Q�v�a�l��˄�����j�'�8���Q|�]�� #��9j���J�и&����&�4�������;��]�D/ K�� �O_�^�!�C��P���U�Qsѭ�C��/C���}\�esmz���>i9Aw���EG�>�Թ9��ٷxw{�`5�(=<^��I�]����FaG=k��o����ȶ l	�5��o�	h��!�V[����=Cb�w�*X.Ux�Wl��T�úG�^�w �OیU������暙��8�>��~���á���XW����Tvs][79�|����hq(�}ŀA
·�W�8�K�|:�����:ϼ�[ޞt��J�}�@�
����{��+�\���pt�'L�arOL�\2J���WZ�Zl�؃�:��w�p�y���<.r�j�_���=�=]�cT3�PX��n�g��Z\n�	fG�Kz$���r�V�O½b���۲kz�;5�_�d�Ól'�����Z )K0�K�0���s@lK<��*�n���'��!��*H�LS�M�zV��thEn��������"m;��F��	���F��?}����=JZk��G��5o#9���SjmQ~����{WN0�G_zs�����8���lYs�A�L�eg(&��q�e{]�j�lN��<ӣ�+��?���k�ޗ���QF��y&�d�!�N�.3��kF#v1���Q'#�� jÒ.[j���	ũí�i;9�a��t�>��1,y�r�=��]�-D?�t}G/�qy)��Z��Ѳ�N��3�8a�j	I��&�������X9��]�O�=p;�������]�׮v,K�Z®�r�²���!���
ܗ�6{�mWs�e�`I�k��	jJ1>#۪"m�+]�E�U��L�y���@��H�5L���c�<���s~t�������F#���2.p�q�Q�	��rUj~�h�
���И�����ޗ�L�7:�I�R!K����3��˂(�=���ͬ��ag�1��,�����P��n�l-����������@�ݍ/�(zȃx����}^���~d��x==j�|M0���h^�8>�2(;��z�>�m��F;^/Qd�Oc9��k�m��N��la������|�Lb���c�B�R���ȟ.�b[M�;u<�Y}�Sx��:������q}�yOS���FT;Ha ��x���R!�?c��ӳ6j��2�;h�é��H���)���s�ꏞ˩1�*gZWs�3��_�k�~�*�%n\Ɯ,�~�Y��qd���߽.��6��7!s������{4wW����uC ��&�'e�����>���5���=t�p�ڡem������Dp~�D/�˂��58�Ì�:��ҟ�ol�"j|A�,[��T��$d�/�0�!���!X�&q>*�68�����f��eN������%�Xh��������ľ�a[��a\s��t-�*�|���w�rfҊ��Q=�㳣��랆z�Hi�zl��Er�T����]͆��~���J�bo���������|�͓�~�e^���2В�g����C*-���k�[��_}���R*��a1�YB����X�;�;�^6�]��1���wv�!ۘ�-��[7:�v���T�%�����1M]K�s��`��i/��q��-��ܓGuʹ(��b�B�j��6�k�۽���D1��+f>�匤ƴ]��3kh8x�I�aP,U'��vi����6{X`��q-zZ�Q�_"!��^���q4_[Y51�>Am��s*�T+�z�
dn-���gɻ=SR�_2mmdEQ5�U�g�#Lys�9��ڦ1)�pϦ|�5��͈�~�8���TZ�8	����g��MO��r�������6pÉ
��.���-������fCD���u8&��t3��;v�_
��v��&=�O.�`���Z����@�F�[�Bc5D���UV֌5{;ײ���z)�?c���|���٭[	�7�B�x����O�}���#{�Z�+�5aů�*����Lo��������2\UC	�q^��.�G�my��hL��2۪�ܳ8�ͭ:���07IN.�R�;C��ψ�wӧ��u�8���)z& |DzA!3���^jx��mL:[9��d����R/dWQ�)�y#<^�BOm���z��ٙw��瘋o��e����3��h�͑�@���<�(�v~4­R!ٺ�T��L�s����k^����:�bܙ��c�sۂ6��#|w�\�<�t�u�\'��OC�^ �3���e�"ݚ�l�`�D+z�D�ƁJ.��������-hG2��;�i*�j��K]�u�u�H,�����	�y(��_bt�<K�lDMW�U�*�Ʋm8��p��f� 퉆MK�֭zZX˾%.�O,��+[�b�ǣ���n��;![����^�w�Ri=��>>�{�'-ws�	�R~�,Y/����C�������r�qⲨ���S#��v+�+K����q#0�[O����n��4;є�m�6I�OT��qf,O�^�c���o}�,��ZAU9�A�|�.6�X�~5#^Y�2LGK���y�{�Z�"8`U�K����]��V���#��o3����%+=לa7czu�
ٻN"b��ޚe��)<hC෦Dv�Dȯ��΄sX���h���بW>a�PH�z�r�G-O���I��9�fi3b��_���$܆��� �+�_�^��5�x�c�i�wr�{��gQh��GO��w�H���K���W)�'!/�|������"V�L�~�c2]e�qLԖ�{���]η�%�V�������^w�.���1�Pnb_���<_�S߯v����y�	�x#����)?0=1����2��h��6���f�9���Tí�p��C��	����-H�B瓉8��=>�O��r�ʸʇ-C�K�/���O�O�[�IX9��av��U��\�=���p�6(�������K��x��ō�"s)P��,g�id�d����Wo{sp[X���l���������9Ӟ1�u��VQ�M�˲�����VxN�Wl�Ґ�A� ��]����o)_4z�Ŷ��֑����,5�n�vWR����l�Wt�@|]D�=`����[�ۺ�\4�*I��	��GF����t?�)��h3�~��zx���У��ї�5���
� *�f-����}bCW�{ǘv��͖�(�2����W���Yۚ�rh�ǳ����;��l�u�(-!m�-!���f���xG'�1>/���yMj���aP�#S�]��KF�3��9��@'��ϵ{JD���Cջ��齰�F<;�ņF��.��Ȍ���Gr��a[���W�Cd�`�;�����!QR�m�_�3�3r�m��7��m�k�p�_Vu��h~�&|5����)��}y0�tf���a^��j��!V�s�
߲����]�W�AY���F�UH*�^U0�ɑØj������"���(n?��rm-�ǹ��*����8��v������t���ej�l�z�1�"q���ϡ�;�U9��ٌsy�-�7����c�]�<#��y���V�ʭ5r�1VM}ǓeO��U�����2zvZ�ņR�f��ƽ%�9�y�z,�z��+.�wJ�h��귪_�����x�g�3%����H%B@%^�	0 �B��Y!���D�C6�����;C�;�P���5��=aIP�Y,�뮠��m�bM�&۫v�um~�
����#q:�B�lsC�&7�>&*߱�.����\��g>VV��&��5s�k�sی�v��'9��.'0u K�r�����r�� n�9����.Ο��}�n��BH$��v��"5gJ8:sUޖ�3��� _��P�g�7���ɴ��r�ys`Dw�9��o}vC�l=0xO�O-*����t���[��T�����9��1��p��6���r�����8�s-5�R�v�n�ؗ�%��`e���^vsm}��ÌEO�3�8<m��0�Ȼ����o\���������5��@W[9L�<ù� �x͸8�z��gS]���:��!�J����m$M(��m���۠C5��Ut������}�>���]A��Aj�PYG;v���5�%#T�	ڜ�rN���>��ÔI���v�M�g�5wW�soH�X�<<�G=�48���o�e���a[W6��YY|�è��Ǣ�0���ygF��ip�SF�lj+�
���;����n���p&Wty�]L�Y5��a�Ө���T��H�aG�S;�v�H�!�V�<z���b(.���vk���חc�!W���R<u'�X�q��8[���LX�2-�i��6��o\���:
ֹ��*Ak�%��溉��9�q\�i\�#%mm�v�rFԾt�yǶ�j���@no5�x��4s���ԙ�
�[69� �KR�gpu��U�>�6�h�ͧ��a[b-q`�W�Ƹ��*l�!}�Ӫ��I>qݝ��1ٛy��m����H&K�#���T{� æ1�j�G\�s&\��YP[��I�We�;�S�!����aN�����X�f�C�����y؂�xb��:��E-��@C�P����G�����%�2����ݪ&�W2{J��4�7M.�T�����U��7��=�s�=��-�7J�e]�=��|��;R:*���wu.���3�u��m
�k����\KeD�Y�ڑ��Vwd\��v���f���}�q ���k1��ɏW(�/�h6�/nV�O7�ms1���*�)�N��k�8l���l�3Vw�5�~j@���i�o$��r�ԩ؃Ef]ca����Ly՛�eِ�:TE�cF�MS�ձ[�D�ʓRRC�RB@�`S�"��.�5i��Ѥ���Tο1@L����$�	�~DV����{MP�B���0aXe2���n�+�}:aT��W*�nq��u�uyc���Y�Q�*u��3����&͠�Z��ܵ;�32$�i�X�R���S��q�@�Ks�jᲵ"��n���:�c����є�0�M���q���ݲ����KO3�׫�՗8[ZT6]"��ȥ�҄�o���%ާ5��n5]�'˵�G���3��� s�t�52m�)�i����>�8#,a�t�b���=MB^ַ�g% V3��g7,Vk~�t1���͹i=�&��)�
\�Β:��w��sOF�@L(�;��xhotMsx�a�ʾ�;���JٖK�2WCK���l)x7|qo拕����1��V�P�v�%.�M��\��3���)�2��'i��j���L�X��(��?t���6��ziqoN���Eg��˼f�l�=u�5��Ԯs����ow+�Z�4�q�9�M,�z:.���&X�+�\+
������G�o�\;I2��Tzj{�-���=`Z-�s���2��=�a���r��3`�Zx��\N��8��/\}}|y��XĘ{�����@mT��)��o�&��!ane`�M2:B�<��saΡ!�rw`�N}�U�s��C��p�@*6��L�$�4���H9*��<@A�t�B�@��� )5@�0�S�:�D�q ���R ƙH�k`&T��L�-�	�6��I�[��I$��$�C��RrU2$S)1s2B�@&ۚܨ�ޚ屭|s_K\E��ח��==��k^������}{����y�|�m��\��j��Tl�/���KnlXƿw�OOo�z{kZֵ����������������ֹ��[_�T�".����O�z{kZֵ��������ˣ�"w���&�0Q�mJ�{ך�wv��X+��Fۺ�r�Ѩ�r�h��^1nj�i5�~7*�*�����sr�^H��Lll^5t�h��ƮW*�TW���ڹ��Ώ���sl��5��6����o}�V�\Ѣ���r��5�m�x���Z����E���x��Wwm�jw����r��K)���l�����&�	2�gn�����V4�̠U�c�m����N3��/�@�mM̼*.��;U��o@	�!)�s%.Z@�[?D("{�lSU�gZ�a��cD�	s��MNSla��L��'��ʭg��7�-;#X��13�U��A�LVw����?�-��-��FV;�u������S輯�J��jk����W��"���Es.�k	4���޷�ae�|��ʕ��f����l���Mc�f�T6��*U$�<��G��\K����]��cW|�ߥn#��
�~�R��x��3�
�#�k�MyA��u�fm<5��'*�l�wtqݬ.�tv`��y놳Ė~�ܹnnS>9�;�P��|F��Uve��,��݀L y��)hݎ%��[���4bsE�[,Oa=�yE.3@j�\(Ⱦ!�T;���Q��BK�A�oT�Q6K��߬q�qRyS- Hwg>��(�&�E[ot���(ɐ���8�<����VԳn+&=4\����iъ�]<��
��]����m����5�_�|��o��
�_�[�{Į�3s/ys��Ua��\�)�Svܟ^�iJ���\VJ?Eս:�h9��e,�����@{�˻��I2�j�h�*���H�-���+^�*�5���?��s���ݲ}�MP&؜d6���ۛ���?���"�՟{����_���B!�8����/�_�������m�Я�r�#�P˼���Ϯ3���U��(a��!nȵ t��R�x��[�y{���ő�]Yx�i�eR�i�U_�w�t;���:`�F��{�|l'5A7c�ʛq-ٚ��
�nt��=�2�4hP�8��X���
�Q��{T,��i��'g3����AZV�&|���l3��r-G�:�Ŝ���[�<�m��=�3�V�n�fY����*~I	)4y`�\���=��(:⺪�s�Jv��W�^�Ò�M��Q{9���r�|������M{X�S�u��ON�w����-�-�k��12�8�hx{=E	�)-�[�hq|��c핤n>�
��m��(
Bh���-�_{�Z�#٣�
���y��9@c�v�+M�7w��r�*����g�p;&�:]h_��t�T�S�k���t��ŵ>.��tg^�����W���\u۷�+�L���J��V���E�%I�o׈ⳃ����̿��ݒ�J�mhl���/�u�m$Ipʽ��9�� 1�R��wR��/rgp������`���a�Y�f��P��?s�t�}����i�\�W�G3Ɣ�#LŶ]�k��x�"x�w{�m]˲�l��J�����;��rDive2mB)��р����Q�^�݇���S���ٖN����>�T�γ�2mAzS���,���ٳ"�@�ka�>�]�}�O�Y��c�G����y�	�מ��{`�:�&a}!�|d0܇�Q�GuA7��u.Q]��մ婪�.+!�M�&�ŐW���7���Xi���S�=�	�T3e�9SNd���~�#rj�͘�Nfo'�u��
a�lCxx6[:P6Sʛ��	����ֽ�����[1�!�ϵ��kC��W�ʃ� i�эB�a�\
�]>{�Gt��_���G`f`(<c�
�z��NY��p�G`��<+��-�輁����5�s��l�F�^<�ed��=�x�4�P��&�����j����	����V6X�u�1�G{D���*s�F�}ԮW!��k��Z�lBо|1��mD(�j=�N�,�[0���|�P/;��� ����VW�Җŵm5N�� T�A���}�/�}�r���^E85�û�=sy]^ʩ硙�e*A2�Fn_fO��9�#��)g�ݻ;2�]�4��A	���`Ȫ��G��f�N��� �cT�O��lm�_�Ϝ�9Ӕ�a��X>yɿvb홰��A� �rE���Vh��a#��vM�儋9�sN���t��9��_�!����՝6��y�+�b�\v<a:1�m܍�~��w�x���	a}ZJ'2�sqF��7O�H�R��n�hk���]]C�uW�|r�_���蘳ѸoU+�u, ܁Q�B�'\�F�����d¯h,��0�w�6ى���`r��{�p��\���#"�D��[x�����aNc������ ��}�g�Г�2�MO�=�`�\���$=��_��2 2>��R���@N�����;�V���q�;L0� ��U�f/�#����PZ��N���>ݺ�*G�>��*ى����G��EJ�/�o��W�'��A��}aC-
�"�`���H�����O��ѝ��˹s������%j�R҉���NM���Qyo-��5�ڲ�u�p�#�GM�E�-�fXr%�
Yi�%L�2���?�2=V%��v� �f��� k]����(�����\c�~��(dcǹ��m]��]M۩<��⏖��у{�E����x�oR��v�F�m��M4�p��z����D;����Q��a�,^�{����vQL�-�~��Mc�[�
����<�W�J�LJ}wA��Ր1t��axy����"��Ę�N�-%��;���I���[/j%��.��&�vv��,�N���F1V&[�����~�{�.��O���-�,���i�96�{*�/�b��ɲ귫��T>ڽAj���D��%�ɉ2��=1�	��7ᴧ&�X�P����OT^��>�EW��4T�%�(�TK��h��xw`u��WM^W��U�қM2���.�4>�0R��h��;�ϐnRkЌuMM��81��vn<(ܩaH][��/F��0����O\5�1�`��'yOs*����
%����%]_��������P�/���FrT�
���yYw��1�nx��"���n�K k:�H�������"�]-mC���ެ�wC�p�܃K���M{۹���	U9�|��UX���N/�6��]׳�/�&E�����үQȑu��r!�e�
�o&؃L�W.l@�[l�m6�,77i<s]����1����r}&�vd���TzC�*��x{$�6^�W�����7)#R��Gjs�IR�ת�ݘG�v;\Ŭ�u�w��f*-Eln�y4��bE*��%�V�����Ժ�hF6foxN�������B�D֩>x�_������9�f8#���_�����j�vB9���q�D�ΛS���k�Q5���9;SÓ?^۽�f�%��fђ	D^�L{虿Lz��>�%���(>��u;�k�NN���7X�5�ߨ��Gfd��� �B`���լ4@�ϖlG��1�vC_�R��LN�C4�Q=�d��	9�&u[��g;�Fs�G��my��[Y�i���E_m��g&��2HH)4,��sL᙭xL7������)������x�!���p��	HSԶ�{u���\����@��+;�w���o���Bn���8	���T��LSF�A�X�ނ�YӸ�z]Jѵ�IJ��Ц&m��w��tk��x�ѐNsk'n5�of"�h�6�1���w���� ��1H���w�>+j$5�N��љs�S�:wkD�sSf�.b��ؼ���s�| v�"5S(:�E�?���G��睌E��#��פ)�I�d����&k��F�Z?O�i�Cw
z��	�&{;��AMPڝ�ؕ�f�7H�T�q�v7��H[wQ.�����Dɹx�]]�	��XDt�m�����Y;2��3�t�27b
p������뻊��g�A��uvw��!�:T��ȝ8��hD�f���vt-	G��e��s�Q?bg �J�T7��j.�����{�Z`I5��Ԩ�J�<����rs/��C0�[[�;U8�e����2���"7�l®Xmli��=�CF����o�Ʊ�4a��3�=��W{�
�]"	���T\��<<`oxS{��ik5����CQ�i�}%��K���1���^�ΟDq�*��9�2�j�*�bsZ-���06��G��_N �N�.��'�Vز�պ�*���=)�:��v�]Ai.a�[�p[�{�-ڠ�e���KV��f�]�Q߸fi�σe������^ͦm\�㾾>w������o7��ŘW(�\	q���q�ܕE��¨������t�3�F�o\�ёH^����F�
e�K��m�|Y@i��H�[@A�� f�5v;ǧ�V��b��ޟ{��5-����iq\�o���,�~-$�x�d4�j�O����k��l3	��vµ^ E��F}�RL51�2s9�h/lU9%����r���NWuE\���/9��̇�=9V@���[&��/CM����ݛ]����M�]�\�O+�j��W�J���lZ��i�Kԫ�{�_��nt��� �=g�Ú���4-y�<��Ȭ��̪g~�����h�n�I�G2nk=
�7��ecƴ��zz��'!g	P,??���=��t;�b��&�*]���B۹���=�2`Lëy�w�o�������a�zD_l7W�7/�.���MF�y����p�s������lu`�8g.��b#����@R�}�]�6�g־�������{l\�W���vQK�0@H��e���4��"�f��/;z�9�F�e:�Yec������VD���3Yp�~��S�4b�X+�߱��JD�KmYprKq2Xs-!- ��0`��
j���ٛ���vu �Z����V��PN��`�^��t:$ߒ�UL�u�⤶ݬ�kݰf�-i�U8��T��w�>���u0��7�B⟠Nn�v����$�*�	7�5=�\zۛ���^���X�[�����	���m�OY�茺k�-ޙ�Jg�,p)�]�{�㏁;8mqٞ�a�o��)�33�p�3���:�t��i�S���T)�ꬑ@y�R}@��A���ͬ�{�6�|�z{��[�n%��mմ
&�Q���a�^Ju�/������F�4x���y�!�f���vͬ�}�ߧ�i�k��/&�H��s���V�u�3�G3���+��w�.��ԫH�s1�z��z+Y��T�0&����xY�&v�����y�u��� _)���P��{Ue6���%�i=�����+�G�d�����>n`X1c��
_m}��^t��.�6�$�i���~����e֪��M� j%�Iv	y�4����)��<�lj�{����O�� �4�a��Y%�a��.����Z!5
�aO�ٛ-2��ˉA�n�1�=�/��N6�j�[��b�B�〓]�iyx��7svpϋ�5�gF�)~�>q��<�f��q�q���~_L���Om��
���W�E�����YqmX��*l]}��3�'�R�.L��8����.�����
�(��jIcJ �����3�38�z�%V�T���݁G���/�|�4i4u)�2�Jj�U:4�g�w6��i|>7=>��5u��=�)�WB;�y	���x��Vp�ʌ�g<V�3���X��.���۔��ȑ|���@�!�rw|x��v�!d�`z+qz��_�u��\V����U:�fW��������	7\�o���,��%4��p�+��B�d��3�[ot�xv��ɟ0�izw׾�j[Yy;��d#�u �z
�Q��ʨ@�='��D���OCO�F5C>߼���;�t�Oy���{Z�fWP� ��9��_�Әق�����5���cxT���Ά�;��ΛS�9K��;�>���4�+E7�N�A���v&�����L+���Gd~q�p���xT<�����휝A�Ove�寓=�Ƭ��Y&�Z)�|`;hVr沕�91vw9����T]�8��e�u��g6�eJ�.��
}w�7�9�$6FcПodG1�qZ�ΝyD��er��j�h��we��{���+0�oN�1��#mOn�4��#$��_Ğ��t\��Ar͹-�����y	3���i��(@�	W�����s����o�Tױ`]ŀ�w�Gyxo&V;i�3ժY����L�j+n>�6H8�b{Yԧ*�F�ۓ��g`��:幸�V�]a\]&\� .�9f����S*,�`&h����XBԵJm{s����&	+7u#G��P�7wkq��Z�u&m12�,kv��}R�N_]#E��kYG-[ylֳ[G�loR�lÉ�싧b)��ܹR��-�.j.�f`�r�C�Fӕ��q�G���8��1������b���Re�f���FS�k��� �3U#��V⇪�ՖH�i�ڦ�u���J>�v�^dCʇf�\b<�್jܥb��-rȯu���E��R��:s��E�t�t��q���r,"^��r�S�m4�)��V�\��:Ty{s<㗌�&��&:�WǤ�%Ҡ����N]�c����=ў\�Ys|u�̿�EJV�Cȍ���>9��Z/�\s����~�V�)�xo����[�`r�V�n��Vs�nT�ۊ�E����sڵ:
�m7��f�]m�z��N:Or�)I��y��G]�:�G�,�2ķ�r{hot�im$�|0�]5^�r��u��[[���Â�:�{�a�m+���o�B$�A�J����N@��Ƴ�݉���8�����u�B�u
oh�9e�r̲������v��tmu�0�����E`�����y���M�T���nk�p�T�qa9W�1�v�R-�kyTM�0uƒƞ�ed8��ܲU�ԛoo3���B���Oo����a� �nks;2�eҲ�.�م4�_슅��f��n�����*��UՔ�N�e����/7n��1�t�c��-h-gE�3��Vv�G�t,��Z��!�6%u�5�q��5H ��s���:W��I�`T�H��v!�u�bl��V��ˑu�]��;e���H�*��x���r5������ug"��^ް��L��mhl_T��v,�\��d��*����R��zxu[ځ�\9Һ]����d5����$��ǹ�]�����=JZ�Ҕ�VF"��$��g�R��ٮRur�8jtλr_Jq�]�a�*�����6f�C���D|H1 �mʹ���ە�/}w��s�f����������ֵ�{k����������x�&@3�٤IF/ݕ͠���ܹ���(	#��������ֵ�k�_Gק���G�2y ��r2)�Uة�x"�z�����==��kZ������������ �L�u`��_��j�sj�m͹��>;cET�U��O{[�ם�m��W5��zIh�Z*�߶���6��W-�gv�k�yjn�Fѭ�n�b�^�t���b�׋W��7�.�6"ł��Qk��sh��5I���o��׶�!�&�d�6��5�W-�iߛ;mm�99��n�0k���b�n���4�y�W^̙Q����[ԏ
�sr�S�O(o��U��:�c�+�8�@1z���>='W�~ �o{�WG���4`o�����0�/�0:��&�z��G�Wyth��(����$��9)w�B�<��fY���~rn	�|
��`PT�W��HΆ�x���/�+z���g�(-�*KU�^�j�(�<�|�^��O�8�X��W�M�������^�}��y�ʪ��;�c��ӊ�Sor�E�o��_���W=��~Ԡq�du�ژ��Ur�,gp�=��0�p�����.WB�9pY�f�3��uY�V����5]w\ӝ�B�C�49z��ӑ��q�V�F����j���mb�U������Uh7��gq�6�/z{jh������F%�<9���6����m����wh��1\^XNq��e�4_A�V։����^������;����+m��4��ƨ��Ǌٵt�q����#��u����o_)VWM��J�A�U��y�9����N��h�P��@(��R�v�k�^�G""Y�r���kx�]�+�t�r��og-���IMy��}ln�y��������� �BP�� ENgb���9���ϲD``��_tQ�z��W.����EH����NX��~/���_��x,��3{
Er���3��m����Rś����rg7?N�D���(R@v$E��'�l�ޗ�>`�Gf�#��i�uI5��eDFF�);g�*Ò�n�A7��[����L��㏋{M8�3�4+j��m����"�v��]]�Ƽ�*��pfo����|��O׽{@��'�L�6.;�R�]*F�d���җ�؄am@2p�N:�6Tfmb�l7��>~"�է
皳/��`�C�:��ʇ!��Qj��DVG�i� �_������Z���whՓs� �]���40��f��r�
>�'��,��T
�I"bg��~���oU%镆�����U���A�N]�Ղc~����:[#$��A")��D7!�;j��Ӭ��Q�v(�����l��J��!���<��z�4A�[|D������ҙx�Z��@��'B�A�U�u%���Z6���$Iؗ1i�>[W�w>�y׊S7�{u��Y��S¨p����⍡�e��JV�{�8=/Q��*e�J̖��sL�'KF'���|�o0��ۥFt�#��
��mnޅ���w}~ñ���zJ�>0b�w�|��5k���5�����n�'�j�i�;;�:�t�»!0��fs��nH4�>,�p�z�B��%��C�:���W^k#M����a-���`��:ԬѲs��G�*7�H�*}Wb��z��^�{��׃ԗW��n����21v��Rq��Q��\:ޱ���c|GO��M�T���ש�J&&�un��1w��Kf>���ס�v��ʯ(Bz��7wnƷ�n�����`r�J۶<{\(��Fz<�,�b�N����~�PT��t��Ӿu0ʪP� e��Zv=(�tW�r2��v|��<6�6�t*R����5m{zf	f��1���DAS'Ƽd�P���]���t{��v��[U�*o�W�@!=G�s�8��Q�Ѳ�ͪ}���ƁHT�{9�Fgm� ��5g+[l
�6�x-�v���A���˩AV���.'Z�#n7�*`nN+�wW+�	cE!N&{r��^,�>u9�ov�M���,�ubP��r���K�A=ޠ�݆jF��l�J(�'ƧU��"!wF�����_p���`}|9@p�`��d
Wo�x�#U���:�"�[Y�wKy�I9���"��pr+�j߻�{�c')j����gt�Y�icҐ#�6�P�����z#�t���髬����՛����ϗE��S܄j,{)��+!��?��A�D<LWC�ٹ����3���a���-�s"���ݵ�����|��������8�CS@z{G��q�\^�^�֪�9뎁t�����3EJ��7r�4���_CJ�B�j��n�B�����T��u����$�z�_}1y�LK����Q�smu*3��דӪ9��^�[�GsKĵ{�1�s�=D<��6�� �[*9��f����^_s�ˋ���l�vݼ�+2$Z9�2]�ϛ��?����~��ǟz��.����◩���ZVy����zR�_=ϭT�T�3��un�j��7S�`���8/ �wJ\�L+h�*Lf+�l�8��]
t)�9�˝r��};��-C��N�7^u83#n�	y{v�7�{ى���f�a�Ed+Az:��B�1{6]���
0`���VN{~'Ƃ���p�0nJPF����v����P݆n,�[C�ɣ]LKR�����|M��h�14��������eES���	�[�ڮ�c�X������fLr�{է�?��=ds��7�|6��6���W�6Y����$p���D�Y�E�ǵ.=Q���2��V��vz�q7d��t���-�����㫻Gm&�P��r�;<�KRcz�FTk�>:�F�E5�`�q~��YUܔn�Q�V�U-O�OV�I[+���gU��V��y����QB��]�1ޅ�vu�]{�$hwM�dHH)2�)�^�?e��&l���D��}B���~᜞�MJ���/{V��)��Ќ����d��N����*�ϭ�}v�<g���|���_�e�b��A�v=�UMLr��"v�CUk ���#�Ըb�b�o竵/�v�?U��t^�SPeGowN-I�^2ı��Hmy:7ϳEq��y����DJd*�wt��N���c�������q==D�%�w���.P5p�t���#}j�tz  '>��
u�۞0o���i����u��\.,o�2}�ٝR.��\���=�jsF�^���ޜ~W�����u5l��d��!������=��J�h�/$���Fw:���wFwϾ���E/T����bh�|�o¤�j���:�Ƒu�N����/��jEu�,�@�N�84�9���üm2�=I_�3d�Y����	G�@kx�=9t��6`���e�Ѿ���vO��Q��:}X��؂��`�%i�֣�+{�����rޞQ�� ���ѩ	0I ?���
7�Ųor����QQ4�<��ug#T�7���6����Z�f+^k�8��S��OQ+�z��p�]X����n��Z�!}��3bu^�Ζ���w�I��YZ��@EaV%��-�-�21Ywk�t�������Ǚ�Q�]�s�r��Վ)��@��g*�5�5��(f��MH��wu!�j�w�B@�b���hH�z,	V3[��ņWtW�kA�,rQ�C�5�E��9KhP�c�ˮN�I,[Z�ڼ5��Q��To�պ.��hPtA!� ���L�E��
�ޞ��F�Y:Ҩ�Di`����in��D�˶���3��$�Nb/s�bߝpt[a�f������ލ�b{:�gmzE�t^sɁgH*i3�9�]I�E�#���WH��X�^��Q��wW��U[���g�g��֭;������{�B�>@�lt�nzn�q��MT�v�U-�B�K(�ݜ��P��o�|:AW�C��3��<ψ1%���桓�����s��*���N���5Vg
��H��:����/|�d��tB�ۼ�����{�ͭ�<��C�#��d,�b��`줹G?-��k���S{�wn%W[����@N9�O��Vh�Y���*�u�F�3k?o��\&8�}��1�@�52(~��^꠶�ۥ�=���2[���=�,���e�� ��n���.U]$��d�i+S�ُX�	�c�������NlK���9@?��G�޸l9�g�����ܱ�i�[\f;ȜP�k��o
�;o#��F}��w�]�����@y��>m�B�T���ƶ��hi�C��m�C�6�5��[wv��7�����o7�S�V��+"������#���+ǽ힒X�[����CM����bw�-Tz�?(�2U3�_����U�^�wA���>�!��q��eڈ|0f¾�i���i�4g��ILF)������t��^��(+"<���a��h�bfj;��d3�>Vg��n��O�ܤF�
S�/gQ�[�N�(��q��ul��5��0�a7�U�2�(��`��a���+�6���ef׬i�}���fy&�Ix����!�=���	��j����&�O�1�]���yG�xbD2�]�Q��u�ǉ��>�c��c��������B����]�r���O8L$����i�[�q�Aq��x�<�O�f�F�V��a��K���RH�ـ�����q++�;Qw���u�k�v�JO����%��4W���c��WS��q9ݓG��Ս��@J��@ĵj��v�
n��x��6Gp�]J�����b����|���������ͼ�%�>������ a:��e���(݃y:%�]ʇώ������U�p��V�[b�*(�ZD)�� �øA��+63#=@s�.�������ۇu�pjŇ2���=q.o���_zpL@w0����ff�P���1��g���u�̓�ioNԣ�i��i�s���X�����/z�*zB�oI��Z,�Vܦ�J=���K���s�O��7-�|s"E�p����1�f/X��c�Cu������������6V�	�0�O�}�;�d��o��ٳ�i�,4\ʙhJA�SZG�����ܾ�+u�nOMk� ���(�٧�OUOg�n-9cPe#�EË�Y�8��Q5�z��&���[r¦�9F������K`�a����B�`ު�^��<�ê�k{,��uXk�[���4zA>�>rVY�ǦH�}�/3�_��H���B�rl�N�;bKs�9�C�F��4`k�}���>q�"�C����"w�Klf� �n���s��r���	��q)T�IE7."�Ui����ةν�� �bi��9��7����kW$�n���
�n�]��׍f���T�h�庝�U�ń60��8��!G�n�ʾ�o%q�;pU�ڝ�xж��+���Y��Y��v�F��Ff��y����lͬ�9ぁ������3L$q�@w�)]�#�<�9+�2� �R�G�
2=��2n�!�l���9j��l�і7)��P��U��a2$
@4"�ɇ��X���;�>IF "z)J����	5�#���^n-H�]��ڵƳ�]Ŷ�\�Z���F�>����E��y}v�ǟYgw`��O�=P� ���Fv67��Q��+���{�x��:�����ĺ�l�����=�QT,�y�wǹ�,�gw.�/5�<͡�������wv�tq�Ǯ�%��fu�g�]qk�������ƛ`��p�����;ԑ�GwU7�v�۲ރ3�敢)L��Շ<��vF�d��?5i$�S�X/	��ҷ�o��;����W�y99�][y♍.@և�BP9lWs�O�Ҿ���n���1v�Q:6a�'aUNq�D��d5?p���=��0�W.�!竣�wݏUʠc��([������N���t�e���L�s�����=��mַ�q�'���t5��m_NԶ�ٲ�f�ڻi�Y�l�1�w�`v��F_�9�-}T�[de�۱xގ�����;XГQ�˞�x�"���wܜ�S�4(�����E�߲iu7��p"Z��^�&[2�KS*��A�����f�o��R�emt�18�V)�`��_t��� �b��ͣ]�l���ۧL��|�ڂ��o^K$ǖm��F�q��`�ifb�\ ��gz�R��Y��p�����;c���X�Ӹ���X��5͕�7�F��+���
3���VEl܏�ڊQ�LK�{['R\��7|3;&ۦE���&WSaK�֝�r]f�U��Z'/y��,A���Pн��^���73}m�\^ix��Z�n!��0���t�UK1�Κ�k8��^��A��4Q��A[O����u�.LOhow�$�2<]p�IT�ہ�:uŹ�R����ǜ�NB��^�ye��|4��q%Ӧ�V���e��И�.��#�9ٕ�rhv�чpX⧘d��;+����P"�̮qw+��G����3��h9\z�v����i*��Ġ�;z¥*�\�5&Y���Ïu����n�;"��)�DIɱ�9}5��髋GBSZeF �"�\�S��xݚ!��X* �F6�kZ��,�&���x��W:��WyXҭV��,	D�l�@wu��@�c�G�I�)Dz�e����6�}j+[�+!�W�9�{��*+�N��R�,�;�A_@9x�Сx;u�]�W^�ܮ�O�u�.�n��2����L�]Ӕ�/i�v-Ю��3��4��ΝJz�e�娍@�q4Ʈ�|ao'e�(�XR���[S�L��#����i8e�WV�����(�s`x2��w³Z�騶�	Cd|r:U%��
��u sZ�wS$Φ4�(�� kY۵y[KV�Nl悳�Q�px���n�.���(��WmA��#��)@�H��6���{D�ԜЫ�1��o:�h-M�6�
��`�N͠��)F����SueC�y��u�8��E�����r����\� �]��d�􇎥��M��oU�գ�E�:�.��'���m��Pvݽ��Sۦk5���Y��F9D h��L6��Geft۔��X]� �j_ �#v|�]��@��n�Ƕ�V�ܳ�M6�X� S�j�7E�N�Ӑ�"���V_9�f.xĆ�U�2��X�< ��@-\��ɏm]�n�(����2�;Ν��Y=�/.�J;\ ��N��e�є�̑vm���`�l����X��c��զ&6���M�&:�;��e.�U���:5�Sާ��'yN������u^�Vl�A�9�0�2УE���&(��(�I� �%*,y!H�N�40��$%����-�6��>)$�e;���%�����D�`&�Aw\�*WMӠx�Q�ƺHq˓8�8�ن:p�9O��1$�!���/�Cȉ�C�����z{kZֵ������^^]y"�%���Q�.W4V+�z�����==��kZ�������<�����fA:���O!�D�9lj�j�n[�5����r��==��kZ�������<��������k�oE���\��r�oO�zj��˷+���y��^-�zj5�:n�湣D�b�(��<Z湻'��7��o]�w]�b����s���_�orB�\���I��k��T�c*�]ݠ����\܍����Qi(��1��F�`�wV-�ţA�A\�ю�S��`J	n�@ �l0\���,�c ���i:I��[�pɩU��$����œ�2��M)ЮRT��fJ��n�s�-��RE�/�	YESM%��$�"fC�F[d0d$�L�R�2��d0`� 	uh`+dVݺJFc�� ǯ'�i�=J�� vņ:�-F�F�w�Ã<�}Ȯ3U����I�~��`1.�\��}]���fϕ�3�:�V�ⴆ�ECA�bc�Q7����(��@��^\�Eu9����'�Kp�iW�۳qY=]��@���dЖ�g�č�1�c�F�vV�;Io��m��T����.o�c5p�O3����O��\Rk�2�mA�� xy�Rȼ0�-S�"���m�<"�c3�@�	3���[�n6�@�B�e���39�nպN�G�$�P4#�ٞ��Ca����I��ȟU҆][[a��l���AY��Oo*Bu�WJv)�z��0C��=]��zkr��B5e�����������#��
�����:W_wr�o+�.�y�+k's+4�}�ٻS�s�[{��W�GO��o/�G�Msz�s����EL��u���z����'h\}�������|vw[�5U��4Q����]h:�vQ拎���D�Z׋&#��vf�Ym
p�"��,�N����nF������ڽ���ޒƀ3��$�,�ݺ�DZ��gCr6�{��ٖ�_aW�2��"U�0LΫ��F���\����/�U���=MMVK�76k�wϚ��Y=y��7UBU�%^�E������F�'fr�[��3����r�4n_�j@W y�����:��c�1��uD�zՃt���N���&A[ƂV�6c�ێp�O���H�n�Vx9���!k��ɟe���\������Gn�ñĶ�;�]DԄn74�oy��zb
�
}:�����ע�B�v`�	�y�լ�+s���7O���W�&�<K6��Ɇ|��� �;;kOt�o��\d'lv�}�����v��>���A�|���q���7�L�hh��A�����"ߍ'����FכvXo�P�rd{��r��������V�*o-e���(1S�7%ṫy}�F<����1�d`�WV�����3�������ۃ���ԣ�� �s�8��ڠ'bE�ݙI�����"!�&�fH�7{��y�ȸ`:V��V=ȷ�ۦ��E�Gk��p�}6�ڽ6�N2�����[����:<��fͻ���_�� ލ�-Yz�3�����A��-) ��9;Lc �p��0�o���^3fKNe�q�����#W�.�<��]�\�3j�'��=^SnV����e:W���hмFzf}���DnoP�N�ٷy��v�8����#Ol�"&�bpג0�����L{b���w5U;0*o푔���V c��rS��fk�k$sR�z����4�����}n(�����p�v��ur�xV
a0v$s��}����ͱV�#!Y�P�Rۼ3O4����%�ˮ�(��75Oj-8��-��r�`�ww 8�r�.;q�w��r$fv�4�/X�T���i�wN��I�dwd���zz_���M���n���W��^����7+�*�>�y�d.��Q+�r�]]����Z�: ~�ǆ5�}�+���%���G��Ǝ���E���8��������O?y����^��t@�ƌ�&g;�s�@ә��T��WR[:���������|�u�V��ט�}����+g�]�}�%}��Jՙ�ػ7�r�(���}ǳ;�r�ܒFi[rjVx�o���y:�K�N5�7���&۫ը/o���P`��ya���i�����q�e�ٷ�7�-���M�^)�.�X��u�n�M�Ow��Q]^�_�{%e��q� ��p�f�:�͒haބ�������~��΀	��J;.U#�J�]�xq���V`��c�&�Wd��]V.S�Q*�ʣ9	��{Td�N�Ĥ*��C����j�����|e8������qݔ(��-0��
�$pA�+rf�#Zv�	}�|�a�8b��T�*�ܜf�h�a2����a+F��F��9X4-�n� Z��|P����Ϝ+�5;NȻ_j��t/��?%�oW��E�
���omO��x�	C�}�3)P����hokŬ}�H�m�R�^o]nh��x_b��8>l�=���ni��*g�oc������ɴ����|o������U]}~�S���Gz�b��LU�7�'�W#��T�N+*~�U�m�oE�k\mc4���n���a9k�vf�a�i]h�+�Slz�C�p��� k"6{,�tF��`)�E!�!@ %
�wY2S���)�v��T��0���U�[�1pU5y�+����ڻ�����&wL�+�����'��~dPA���1?:�@yPT�9!%S tL0`���f%U��f�~ݴ,�L��dC���Q����1]����OwE�l� ���y]��m[(��g�3�}{D�Y���-�{���C�߃�DR��<������L݆���+^I�=�=�O>[��p�,�Р=�f��/�}��ܷM��0Pэ&<ჱ6�6OؘV�JGLeD��1�Q?WgEDR���9��:��n:aT���C�p�S[E	�s��|���xiq9�Ӗ0�R�*�u����"�N��|eSw�-rWA���8�d�Ɩ���ϢLCx���4J�ArU7�3}���i�����'�ީ;�<�Y�	v@܏Rq��6�7������N׊2M�_���th�v�N�^��0 B�/5T����&C��R u��&��[���:Y�oFo5'�<b���.���;��������=����u�ݗ����<NE=�)�*o;�i��b'u�p��� ���e�3{��e�t��������ڡ���dW�;f�|q/!T33TI��,�7���J��y։�}�i���0��[���j/�rBX��M������t�͗P�3�&�y�xxxx{1`Vm)[8���{�AM���+_ld3��
=��{�Ѧ���%c�ٛ[#3"!�;���Z�֩E�UҝETN���Nќ�U��DDӿ����!x5��G�~��;ht�*�����r�nn�םh�me��Y�|,1�;c0�s*�H�q��]x/s[��G9ė�Be�v?OkGnk܉�uB�*�E0i�F;8�}�<ҁ����*�3n�8��N��W�$��U�3*D�����Ɓs�u@Lr��)dP�J#*"��A��Ӹ�e�ٻ�������U<Q�����uS��n�����Yܽ007�!���k:Q�j���u9�P>⫻�?.��$��v�;0�3v�:��j���'�9B5E�M��l�*i*��kn��a|;��'U;���,�+#�)�iV��"���W��D�V�E�"���v��h�O�h��KW���'.}Z0�x�d��T�sqsg`ȩ���&��n�4D���z�l�	�C*��T�5��x�c}��!A+%$�K/Tpk�`s���s�w��A���p[ԭ<�lR�۬)��|sZtx��#�Û�Y�ߧ��O�猟:{�A��F�w��)2���S����G"��j�)K�vhm�}���	����S�8�7�͎š��>���=;��(�9Z�z��n�Νș�$z��`�d��dO�|�q� d�������쭄;Z�Ў��{`��g�e{�I�`2���Z}���j!lq;�TvP��!�E��?Z=�V�:� ��O�@����C/d]�Q���>���w��;ExZ�QW~�x\fQyR�C=��zS���_t%����)��WO���;��t��^���UWr��%��D4VM�q���ʷ89�q���Y��a��8��Q�O��L����g54�<s�����{C-]:�[���������p=bs\�L�
��m���{��F8��p�{�G?j�幆%�M3�G�^�����+�g��.�8�yu@��ً^�WCB��@X7{x����ɬV/�����/�'L�U��8�wR�k�=ϲ��!5m�]ڸ��}wg=7��<ѳ0��ޡu��7O�T�B8�9�+�x��ԣԫ����� xFJ��2U5y�A�.��𺻖�2�\�ѹo�wٺy��h~��;�����_
�"��2�wYy��Kel�L@�ԋEă����w+�b�+��;�OW���v�r1'��%nOPFx�m��p]�T�w:�r��3z`���6�=���";T�;7,��:MW��� �-ay	뷷ku3Z't�n�(-/^�+�-��A���}�5��!o���<�1�
�Y�R'b=���cy ���v���q���kz��q�};v����i����o�gS��MO��Y�h�сz���ԡ����n���a4\iN)C��<sqs��	�fj��n5-���qˊ�ծ�=���Қיs��}���31�,_z�u3�䂹H��/&&�Un�6 �W[��>��^��0����bc߾�{Vߌ����Z��g�����]�jb@ǒ�������N�8�����ut�7��ⷚ{'��l�� ���z�(�8hC,רS!Q)w�������x�
�P��s�pF����jv�i���ܥ��՘ؾg�p��Iy8`5��k�_�Pl�BtS�Z
�0����'b�U;��g=�&=�Rm$���]��|)�����(p�q��j���I��
�_���gf��c���l,:�r�\y)"F潥�'�Xw�/�)�>|^��O*�^.�N��:Ơ��+U���ԭ$i���zn���W
����P���0+��V���4��������'<��ٕP�Om��ӥ�՝5j��u�t�7��d���tk�}�$_l6��lr��?����%GP������v�)SS�4�:�^ڞQB/�T��Y�	�ǂ3��ʾ�Ed\�	n��2�N�Y¨�e��Рq褍5È�'���,R�2�ɚ��RQ�����i�
-Hmm<9y��s[�Iq�ޞ=���5��n似<@��wh�gbF�ޢ��-.f>�X�0kr �g��/�7��"��{9e������㒣<big<����\�-��t��q\��S��D[ktb�� C�I�#k����h�.!A��6���ϑ��;#bC��6�<��72C�8��O7!$�!"�i��%%0�[�y��{u��5Ҷ)f�9Y�£��9�{��f�}�[V���VA�ص\�jqu1]���'_U
����I���;L������Dj����W�`ܫ�*�Fb��V��^y��LV�;~�*�+,��}��y/@�ks��z���<c��%�cɉn㉨�͎��g�T\�03�m	�p��j���,���gN�'r��,��kI��Qޞ�d�l tQ�PW��5���h�x�U�#b�x��YM�ݚm��i�'��8�8'�b���o���ed�&)���p�';qp��˱U=���R���r���r[�����'ޫmm6rH������=�x~��T�}~�U��{ht�����sl���h�� m*N֌��밍�=��_)l2��>��	�u��7i�9ږ-w)��m�n���Y�q.�_� ܈FgV�'�����ܸg&.::{S������ɯ\��T�e��~��q��Tr��||)�Ͱgjp��6p�d}}�ӷ��t�Cu��2�	��i[��I9�8�����5:��f��M'��6�5q�Yi^(Ie>��yhճ�_E�+w"b{�%gd�%�lm�w�E��o�ЖI:�m�"����H�-ۑ]��F��0Wq�3Z �W��]�v_f +�U�s�MK8��q�v�ۊ�Sc��`�଩��s"���>��s�b��h����5
�}���h3WJ7���
��5�X	9
f�s��/�'�d�h�������x7e��s㦺��
�	�����+��waL/M*�e|yT�em��\��97[��Ku�6ڵ	��PTڛΕXe�]�6���:bRK^�I�*eXt�Z�S���%YO�V����5g7mG`�2:*�����[̜� 76����5ӱ�ް c��:=��ݝ�=�\�w2�;:��8(��	���(��s;�j��|d�R��n�r�U�:	A��ǝpN�L�i�%�y׆+��B-JWa�N��D���=���p�I�J�3�v����]=1GE:�l�
��-ɮ�Nn��<W����w��hꛨ+󒉕,���xwu��ת�ݧ�+�4s�d���J��B0�8�<l���d̝ה���b��b8	e�*����(-V:��b��asM�f��}J��n����@<�]l�`]
��ղ��l�����oL�VӢ�e�O%n�����f�u�c��Ջ��d흕�B\�z漥��fl�*c��4��,�d���%�k��4��z��7P�I�9Q����|-*�0{�D]�p�i拪l��etxE(xؗDE�7�����H[��dҮ�w�H�����U(����^L)I��i�W��$iBY�^�I5����D������
���Rk�:Ū��	G\�c�|��u;Y���Sю1q�P�@��� �m�W箚(�k�%5��k��� �9�'e��f�[�zu��h�I�����3pJzU�{j�H�N�]��.q��:���oo	-�����B�!h�����]�u���V�649<��Ec9����j���V⹕�}l���*:Z{S]2���|z[���4��y�� �ҭ��t�Jٺ�ܭF�^
9��VsR/n�b�����	@�����Z�)�:t�˦�ݮ&�v�q��Sm:��9���xK��ept�uҭR^�v�U�匼:��x7�l:�F�`���B��Wo`ǣ8��,��(���t&�9��������U�� ��_'���9�.��;�b��Իy/�)G�YPV�(C��ٔ���l��ϣqU����m�h)5N_ft����ʭH��=j1٘�i��jUQ�ˢ�#��ӂڷ�J�oq��\�[�Gk�<�Z"�M\e��p-83$JW��V�1A����9C�&2�^6���Ȇ���.
р��G/.[8:�.�J�'.\:t�d��I�^�y�E_h�Ĥ��V�q��I��C:�&:��ӫ�����9���h��e�a;�ڙ-�`ȩғ��w���Eo�N��d:��gp;�~���>|�X�#_x���M$���Lyyzk���ֵ�k_�ח^^^y<V!a�IB�Ͻ��6���wv�����������ֵ�k__^\y�����U}zm{W�5���4dش���ƿ��E��޷�����ֵ�k�����ˏ///�1��܍{V�(���݉� MD�"��|�=������I��v'����טM�k;��������r��i9�nX��Y.�1��v�:�F��}����מ���JJ��O:�ܽ��S2��f�((�Q�`��;��sA��A;�d�&������!N5��ڃ��"���@�Δ1��Ĳn�ܯZ��A ��A$�"	�7���c��}w׵0Wȼ9;���c�MN�9��5Czk��h݈M�\�o7]�ǈ��wX�W������i����"��f���n�|�It�\��ɩy�n��`��?v���_�a�7H��@�J�]�_���$��BV������8�=S@�C��!�4qK z|�6�A��!�l�Q='ɧ������w��-��������̦�fc] zC�v�(��Rok�\���[SWY��̘�����ա�A���~����f�_j�"3��*���׫4�-7owv����9a�6�{��@5Y�՞n�Æ{I�!uL,���6fh�K��J옣H���/ݴ�����=��{*�>c����#C1��VNn�q}�.�B0"ҁ��
)�r� 3������D�Aj��|�7�ϐ�da�y���Gn�0�u���K>Hk�>�1�s5>e�>3������GD`9�)y�T����7R�܄j-��mE�������[�$<���S�K�
�Z������e�lt�g��]�\;%���ۈ.�G�%u���b�������S��*u�q�gd3�t�^M�W8m�L���2t�$�0�Uǧ#<J�b[^c��D��A�'J��߂�W9��tX/)W�ߖ������H׬�7΃�L0�	�E\b�4��=�{VR��x�j�vy�dЄ`
�Q3�^����$��n�F���'��G�}Q}["�)	+e�u�Ci��=P�bj㛶�p��YĶ7�����Q�R;�eT#��L6�L�\O�����d�)�NVQ�����1��y`aG!��V��܀�󢪟/�����88-�}�n�K���pB� ]^��.ȣC2:G�u��u��սMT)�H�\B�~�X��~�}
9t
&�z���QeӈL�^ˠl·���*V�oY>T<d��A���O�,�C��F�G�p�Z�#Y��oR��=���}�)^���T�"O�������d�O���� ;�D+�~0f���eT5#��y�3B�ݑװ�峏�y�=��Sʚ�7��(RUHV��`T5)ln�Ս�Vܣ>r�옞Rљo��ʽ���|���'67�4p��V-���:��D`���ԅ+4�����gh�3�=7�',����3�hi"+.�*�%n�m_]�8������\�ęN�;ngJZ����GP�L�J�
	P�˫f��0`� 0`�g�����V�*��%=�]q��;��4�*W��q�3�l�����>y���ߧ'�~a� ���r�Q$��n���`�;/Tl��8�o��`�k�ݽ��@��H#�\tMK[����^J�t�{�!�%�&jj/9��з��nڏ�	�
�HZϡk�:'��4�/��ږ�m/�1��ޗ#����mɫFz�^��n3�w��F�O���K>N�����u�i[%�^y����&H�I����)��@�;���E)ڽ͘��� /C�ze���-�
yu�u�wa�W����3kṩ}o\�� ��8 �gG)����q��*E ��#�������PnY>[wy���P��Ϫ�os�g�	 \a��pu8����~�>ot��c!Hau�vo�of��@����u��s��[���_*/:戔w��en��R���mYyٶ.��Kݴ4��$�rDNk��xe�%X�0�0w\��_K�vuv��'WJ�2�Rґ	���xN�]
��1՚��Mtt��W��2+&�>.��Թ�۔�x4�l{h��%X��F�*#�}>a�{#U�jPV�߀JL�V��ݒ��W��BGlL����A�;�z����?����� ���������S���� �@d�6��_���[�2od��@e-�6����;�z����v��(6`�`�Ш4K��f�]k��>.�7��`��tg��q��<�� Za�Cԭ����;>k����޿d�J�����}��Ց���0�]'����[�$�ʄ��U��_UW@�2�᥇q�q�3�K������z=�JӃ5ubE����M��Ya"�;z��=�� ���Ba�YL��+٨���ff�g6��a�H�; ��ε�?�^3�M��aA�3�s���b7U?O�ٜ��ؐ��)�2�;0�M�;�VX��ӹ�bF��{�] �
����T����1����(��饷�N4��=���YZ�hd�ri�s�c7�;��w+�1��9a}�w��鼥�i���Mw!�t�i���ź:�F�:��H��PS�x�������ٙ���k�4��������΅��=�
[�oRС�zJ���e�^A?�վC¨y�2�j��ux>�bƉ�Y3�1U�j㶆'����3�y�r�4wP$�^�{1|*���;б/C��z�ڷ�����jL���[լ7H��b+s����U���T�`: �_U�\t����>&Ѥ��b����[���$nɧ�M3���UQ~�o��νYnƚ���ɸ�ͅ���GPl'k^�%�u�ࡁÔ��@��*��2t���;�4 �	�ٵ>���W��Y���ޔh�]�X��e�VMWQF���+����n�~�팲z���r{n��a|ѱg0f�����3������뻻5�-��2#���77:f�s���B]݌��;z�CH]u�]CN�����)ٷ�5����߱�3�Ò���lYe���ܱ��v�I��'wc�tudnS��o!��x�`��cT���~ 7�?&����s��/�ļ�6�7��P먠����#q�K��M�	��مIu�~Ah
�9ݤp�w~�7���H8u�t�ډ��0�@z�9�g�tŘ���P�/�*�E�Q��y�wt#O�aZ�W"�0�����o7�� ��7}i[��ɜ�_y$v�i�S�VHڟ>Ϸ;`Ge{'8�;�Y�cg/	�/����t����#Ce�BEb���"���wC���x��R�Pb�?@i`�V��vϰdz)#�=KjAnE����lnз�j��RO��vX;}d@x��\��0bs-�p�#�~d�Ɛց8O�ۼZ�=��0�T>��!q���Ú��Q]���9��Z��v&�8���Uؒ��+)O�ӏ2�j;�US���u���EU�i�7�ze��g,K��:W~z�[�q.�Z�Uz�r��b7f��� ٭�U�c������:��%C��P�zB۹٤���;�w5*MT�y��������~��i�5��;�7.��꣆{l�MoS�3��Ѧg^Y�B���>�=��fyY~�[�����Q�kv��#�h�����Ş�;�������$�� �C2p=*�T�'�qR��Pn�%�vm���vE�S`
�Ml��� �A����J��$���\�H�P�Õ��-*�/_`�Z��*��o`D�����Ơ����LSh6�A�"[
Cr��8� � ������yO�h$�A�V�vォ���k{��f���C���<L��<�m��t��Ya�[`����]ҵj4s�1�҄�$������ۂ�y�+��9�E�m��;����Zc�Wu�d-/�Ѹ�6�u��l0��Yd�7�Ǧ�P�(� ��w����W��#�w���2�2���OV&��'Esc��$�o0-�I��r�s��qvqD�_R��w��AÓq]h̓��G8��;���]X�l���Z�$��x��j	(X�D^fl�5��6��̍(~`y���]�8��kL���O���i�N��E�I�vw��c�#&~���n|�y��r��jgu*B񽃻�_r�IXH���M������<�V�9����Qn;,���e[%{3�¨���B8�u=0�)�p���[S�ԕFf0�r��9���C�ml���JC�ܓ�\�NL�wo�Te��V	�I��t�X���.��y(��v��-}���{뒢l�q�j�e�9��Vn6H�M�oa:���ۡwor�I�,�.�S�.��]f��t80`�`��^��~��_��T�Tf����+��)��X+6V^|ۜ��&��/.vf7'��V�q�<����U�7���:����˜˸�����E�o5�nD�T�O��`U�n�z�ݣ1�͂N�v�.����ͥ��{xGl����e�1�x�\Ou�'�%�Um��4�.���m�Wf��T�xZ���}���}�z�G(}`�6Fa���y��W�[���T�ǹvy��ڼR^�۴�l2*{gg�1;>�Qw(�i�>�wgi�.P���}�66�D�k��w�����y�mf�t,�L_h�X�w�އ�k�*eUz	��3�q���B���[�
��7�����^-�oU�����^�8#y��Գ���y���Ѐ�H�uu3�M�N{�������77]~���T��\�vR��x�k�>Q����}\"=]y������V3�n��X�-l�f�d`O_m� ��[bh��x��L�66$�����jf�5�U�� ��%=;grI�䦰Q��<#e�w1��3�m͹��=��V�-ѡw�4�yf\���I���`��`��{=i}��ə1�}�#��nV{d6��h�4��} E���)U��W8����ɭ�_.?/�vu�2H9����^�i���;7 �?{ӥc�M��&̷Z��ǣ�+*{�P
Jh������l`l2���L��ᘫL=����J�������g����g潱��r�Ԫx�	�A�T�7N�و���m�����y1��	$n����>��|���Z_uS]wkLU�7��x��Ǚ�ն�a�Q��D0���Fj���׷d��wY�U��6�Ч���#Q��^9#2m�{�U8���z���縀��$���:,k�0�.��탕[���k=�/G�.�=�����J��O�Eq�~D�ywr����?N��t�0x&��7��{K�L�Fq�g5�,�\��eo�FO{������(���A���hn��_$C>/6�_S+R�]�&�ɺ�N>���w���t��'�|En����Y�T����Z��$���$��-&h��� |3��7��dN�u"mu�T�*M�fpD���4�u�+����,��m�N�Ό�rxs�+V�z�y�P0@0@uy���7�/�����w��cG�ߢx�isz�����dln�k3+5�7!B5+E����`?�?��#��\V��>����ԫ+)�����Mi�h�5�vi�L{��]=��Y�-��}�!�L��η�nª�\�޳��r,�+��T)��Y�k�yC_��O��i�k�T�zDB*N9��mMR�99ci�=�m��>�9��9Q,qQqz[�p��vg9B�e���}�E-���e[�O*�am�����gZ�܆��,����������u����y̕,̊�l�u{b$�v�*��,��W�k�z陃k]6a6�6�!�ɖW�J���m���{.cʗ� ��p�p���-®�:j*�菫�N���Yd:������@rĶR�%hy�S�V�<�#PJ��N��������9_3��@\�a@G�_�����@�P3���H���{ow����4��[�Z��kKZ�1���L�T����f���V�2��J���Yj,���Lfښ���3j��Y��jd�kR�j�m���KQ���jbͪjki�+SR�,f�����m��T��6�������J�ԵMM�jm���MJ�Զ����MJ�ԵMM�jkSSZ��������55Sk-SRښ���j���ԵMKjjm�R�55���TԭMM�jZ��ښ�T�զ��jj���6�ښ���V����֦��55��V��TԫM��MKjjU���jj�R�55SSV��TԭM�֦��55��V��i�����5*H�D"뮇�S�B!	�V����֦��55���MM�5-�����Ubq���!A �^�I�[�M�T�-���V��D �C@ �mU-M�T�+j���U-M�T�*�KSV�Z��B"�n�!� B(�-JکjZ�KR�T�*�KS[U-KZ�jmj�b�Z��Z�֪X�����Z�jZ�KS[U-KZ�d������T�5h! wD4 �T ���֖+6Ե-�2��SkKj�,����5-kέ��5+i�5i��f���3Z��i�,��R�1���y���V�KVc�MM[5+Y�m�mK-�c5l��Zfٌ���k�j�fe�,�̶�SkS�m2Yj�Lf֖3Z��Ͷ��m������^������� $T#T1?������w�����>�ݧ�ٜ����.��٧��>�����?��~޾�~��?W���~o����TE��H��*�����9?4�"���}Ї� ����~����H���*v��a��y������I�G��
��MT�SU5���-R�)j�٭JkSVkQ�M�Z�6���f٭M*���)Z�ڦԪ��E�m��ڤ֦��5S5R�j�Yj��-�U��Ij��[V֋[j�6�P�""ސP��F ��QkU3m��5j��TҭTU���T��6V��T��*kS*��j-SSkSMjT�KKTٵKf�,�M5R[SSV����֥SV�T�5�ZkSl֦j�VZ��֦U���Ml֥M�Z�֖ٵ��ZZ�ZZkS+� �T9��&����O�?�E�QQ$�R@@I���@���~������}��4�w����
�����8�s��S{�p�� ��Xr~��''�~P@Z��>�~��"�
�  ���A��~ӳ�PD^~��т�������|/#��00?�3������p ��?a���C���>�W�
�������>��?/����(}�����������W��R��A ~�q�p}�!�H�j���`�����?��ǀz�x;��A yN��`v�}���p����v��	}_�(�����UAD]����7��xbj��d�Me��4|�If�A@��̟\����EU%H���P�%*�I%!(*��QH�)$)R�ERPJ*�*RAP���*UIT��IHD��� T�@�$I�
�UUD�R�H$*��
�$��W�QUJ�HE%JU!EH* H%J���B�;b�I)*I ��IB�B�QTR� (U*%��*�UH�T�J*�"�QD�J�B�IB$RHDIT�  �v�#J�-Z+Mmj��`����e��t��e[TԨRcCSR��&��*lR�ڶ�����J�L��J����e�%�P�T(�R����  k����v-�5��U(]�WG�D�m��[T١x{�F�uB�СS^j4���m����fٚ�jYSJ�m�3J*ڌ��Z�Jl�Z�f�*�e2�E��1J�*I�J%�   6�զ�mi���T�F�-J�[f[kk)��Ul�-Z����m�[R�l��u֦�֣U�Զҩ�������
ړ*Ƭ5B�Z�HB�R�AD�)*   3.�b��UCLёh�
 ���56�)��q���L�kR��j���-R��E٥q��کR�H"*ER�(���   �pڴJ�e���ڦ�`��,�ƀh���AjȲ#U�R� �0�*�SE��,�Җ�SZ6���J�*JEB�  ��4�V�kUUR��C$[#���j^�):*��Cl֦���Jj��[��+�5SJ���H%�"��"�*�T�H�x  �=P���X:��n�:�UJ��nJ��Ӻ���U�WT�T�qԐ�4�9wEQ�R�l�w
�.�BQ;��Z���T�"��!'� ��WC(7P�T���`*1՜�"B�8�p�(UX��QQ@�Ҙ�J�h�g#A-��%E
�:�U��f��D�H���V�  6�y)EUT�U�*�	3��"�(M�n�A��wJ��)D\twQlAͻD-��p;��m�[��t����wUT���uDN��*"ERI���  ���R�w"�����֔�q�P�(�;�Uv�k�-�
I��tW:;���m��\�U	�nU�
)R5���R�$h 4dOh�JJ��@h*x&P@ �JR�  )�@��U	� ��$�JDM�U2  3R�VD�H��VOW�������x�
]K��)ş%԰�2��>�������ޞ��絵�m�uZ�����[Z�����Z����[Z�ٵj��_?�����_򔥏�Dc��%z���A5g+&Ь�[Xr�w���5�u%eaU)f�%��s9�4���R��tv�y�25�sB�m l�kn��c˶�7�j[՘��ecı�e���%����W"q�
�6b�76����6쇢�ٍ�N��"���m�OR1wn'�[�sv��Q�jU�b�v�jVʏ��k�F����|�FƽM)Rj�۳a�JD_�L��6�h��\��ʴ���O�o^�����	�f� 7rLǐ-o\w[)��f���/e�&���!��O"S$��r���\6µOVenGx��$��M'@�+&|u��e��t��v^��GD�Y�K+$���شwuu�Hq�`ͫ�	�H4]c�ie1�7	j�[x�#o41f��+.���Wb���,CJ�F���[�v�m<012J��V,��El�b�
�!oSZ̘Nn�N��'� �I��^�
nFs*����ܨ�<��[X�lX'#�l�An:������
O�F�h�[�#[wB�4*�DflZ��L�w��)��'Ъ���<e��O>;���ٓK��q�Yuy)e�R�Rג��D1�6���Z~9���Wr2pkB��z�3~�c�7����e�r��i��]��I�U,����.�-�	m�F���/*4��V�HVY��(SY����OZ���#I�s��M] ���rdb��At$&Z�-J8�<���Zo��eӁPT�2�q24��w&]�OF6����JyCTh��7+M�v�Í�a�5��'+iR��
�ݦ"glX֍��P�t\�Xv��P`7pLɸۺ�����v��t�I�Alv�.2r����f�1CSN�5!W[�⩀%[D6�\Pf�P^l˦%�P�[c;
B�T`!� 2����!�s+I�X�.�RDi��v5*jL&����q�;Р�|����!u�3 gF
D�n�I٭̥���fE��WVF�z��.�%Mb[�u�j�毱K�Ta�քtд��R*5oE�0E���#���'sEu���A���s,@��+or�ʘ�R��5������Г�Z�ሐ؁���A�%@0��c���2�����L�	.e�޻�������-�(�h6su�LثB�?i����C��U�{�e)F��C�֝��X� YH�Q^�oX�EN(^dj��2o^�7kt�J��V���d��OZ�U8�B3W�4�|����@R	�m��fe�t��7Lh/9C���IAk	�xM��l�`I��pk�u�'W�F��7B�������5�3+U�-X�Q���P�*<�Y�o+"U��n�3Y5W�h�B�s1X��Yhj(L��0�QR>�di����)�|� ws
u�*��)�ݤ��GT8l�\La��+����\J��Sfܽ�qU���5�-�7�ŀ�*���i�V`��0�"�6�4/+V�t�k�d���z��l�I[�J/���",,��Kd��ɪh\��Z$V�, ���Ѹ����X����Ի�������(tU(:éwIެR��BJ�m��a#��#5��;E	��d��sn����45fPf�tJ�3A�mK�%����!j���-l=�c-����@c_�u�<�X��)��]�|��G	[��U躈���u:�g-)e[m�F���3*�T�͜�H�c�����+��ĨX�4!�a��J�r&*�X��IYb�5��W{��
�V����l2�
�e��#LJ��R��7��:�J���KPCf�N��Lw������Ibi(�K{���Ʊ�B��7N:T�W�+�e)[�)Q�����%�5��L��'*K���w���(Xc����R����\��X4[����J�2]j6�M,� U'��x���F�n��SY����b�ȏH�z�[����R@Y�N³1���,�c+%Z{dV!KF�b���|�ܡY[��HRf�32���;I�

zIk���Dm���U�ɇ^5��o&,�(ʬ��:.]�J��u�sB
2ڀf\;42�Y@�
�*;'�/_Gz1`&ԥʁ���nL��-�c���^�� f:e`����m�'!�T�P��I$�7v��K�Bl�J�Z�kj��EM�Qs ̫�]m�Ә��F��NRo��3Uҕw��`45��tԔ��B�����%S*�!�e�j�ֈ�ܡ@1>f��,ԣ5����c��}3ATK9Qt�t�m'��id����X��I�`mMWx�iNw��wim�p��*�֨:g>p�UԅK'�0n�4an6�n�c��d�R5��͹��=;m*��A�f憬]f�Բ���rP1b�8�"
7[&hxV�+H'��Y��f�*�T��L�V����$�PӔ�¤I�`U�����[���4 �IZΊ�-��A�1��M���u�Y��j�FV=͒�#&2���ɭ:�h�wlcQ�5��WF
L!2��OE+˖*��qR�(����m��hf�f�e�u��v��D̛�J�4�X�m��{�l�ʰ��z��1A�S��Yc4M�kD�
])����ݓ�M�E6&4�wDq�.�ʈ����D�ޭ��rn@e�����Xؘ�h��Kwr4������u�&���KM�su@�0�f�\T/PP44fJ�RYn!Fn�t�96�ͻA�[��f�n�o�(̈́�zΊ�ҽ��>�T�n�L���C�4DiWpGE0��Rkr핫MO����TM	�ģ%\շ�e���Rn�Av&�Y��٪!��AM�����劰�[i��#aa;j��4j��Y" �9C31m���R.2�-�%5@0��ekt3j]
�B�V�C@�*n9���R-��֢Xk���s0��PQ�Z�m���;&n�H�%����Y���e�\�2[Dވt�ѭ���ݩ1=���7���V&L[&�;Zj��Y`@Q��z؊�(��oF�qrV]�W*ͺ�J��7�HVF)M���q9V3a���ֆ�X�b�y�� ����F�5,B����h�ǉI2�N��ж�M{n�Z�hmT��7f�j�הB�Q��HF+��5������n�j��ulܧ���(�F�{����pշ�1��i��yJG5ժף ���8L�*m�aU�n��˩@$^�m�xY�DK;n��M�%���n�($L�@�J�cՠ\vjh�n�f��Aͤvi�woi�ֲ�6�t]�k�So#����4B�c	k��;T���[6%rn(��qf�J��*[Tnt]�����9j�1cE��h�9�]� F�y�D�H�JFVY�������­�ae��k@E(���̠N4(�,�E=xe����E)&�BpH��ЭkF	�)�Z#�4̌Xl��kwcZ.k�e*xr�J9J��]��3R�Sc3Qh`���4>Q���Q��5��W��YN�dxu��s	�=)�YR��+3,N�OYY>��E��L��
`d���-��MZ��ҺlB�f�a;V��Vh��a���V"����c3n�NA��Z"�v�>ö�LەJ`�.ť��XYAШ��H��Q�f�Z��L��^mȩ�Í�������	�(�x0n[�5����R��+u�YTç��"ESK��(��X�Ov<9@�f�A��v�8�W��YH7�77mƭ�.�,^0������+��$'�k2���,^��0��6X�C�޽�YD�\����t��)�khZۖ�����`�3#�ۦħJ�n+�C�
,��X$xn��;y����%�6�Ռ�����)�RJj��^f�X�˫	����k���n�����,�4kl�ׁ�vEЩ�2�Pj!?I����'E�7/d�v�M��n��<`�가
��B��u�Q�0V沭k!�Wz�jX����u{"�~�n���G����kJ*�!1h�,�Sz_f䱲\ya���T�f"�L`x��q�6ٛ5F)X��Ts(6��]M�;¯^軀��Ò�AS�-�H[�)ޫb�  �so��vVb�:�`$駂ͽ*L�{��Mcu(�T@�)bN�iצY����Pܭ���.<��.�De��,�kkl��==c�k5��홻5Z���h�i�#y@��B$������w��[(<����E��6TP�S2�mZ�2@Xs.�����n8�v=ڑ�\��|�m��Igv�D�Ô^A�%���又�> �z�ņ�Za8i)X%�5wz��S���uj�E�.�ʶ+���(�����[�J[�[Ld*VF�Lh�� M�P7B;gpn^Q��(̢����d!�`LC@��f��Q0���_�5Y�(S�Xr�:���KP"eX�A�Эۄ�f����0�&DNde��œc3-�l��L7YH^�/&݊ʈ'A��m��u� 6��L��ޅi�*�J��wH�-]�&����6�*0 ��m��
�Y�fb$�J�U邆�^a�����o5�uF�vV��,�4�V��Mg֮^6im�i�1���G�wN��K����yDf�k娣�T�Z�ct�h
�傄�C�%�q�*w�b�1D��`�l$��x�2f�a/
�*�
�ѫ�X���-
N��!�+K7����� ���)�5��pXa���;�K�&\ĕɬ*�%5z�AJ����F �Kp�X7�쌔�.��k^�rY�/"ɶ����6��2T��C[.��!fY�#EMN����e��.��Z�Z̅!�)��f��YBԤ��c�G�}׼&�0_m2��0�;y n����`��do\á�Xed�v֝��MXoi+��Z�Й[Y��P	[��A��d3.,�Xp��,}���J[Z큫�l��OS��.f� �y��֢^�K����
�z,Z��n�̆U*L��+�i�2��������K���M��wB�r�?^�!)Z&�WtsX{� 0���$l�K-�.�ǃ+ �*dZZ�e�y *��Ö�;?L�u�ai#E���;��1j����- ��F8���&KY��M�Е�Bu:`$\�2��X�YeR�b�bp��X�"ք�I�Y�X��x�j:K��4Yd]�.|AL]�pȨ�H����+�Y�\��v2Z"m]e#n6qO��-�x+iP�ʉ��j�U.���("u��ZB�7ZU(2ڽ�J��lc��4Y� Me���R6.&"�����b�*,Vn]���0J�Eޫ9��mI��I�n^=�L5����0�@�V�,�K�q*}bGS d�Th���b7R�n��!ݬqr�8
��Wl�PJ��N7t]�j�t�7�=���������n&r����R����+-�wEe%v�0Ǵ�A��Qx-̙��q�pb&�̖�ec�5�6�%Y�9�nQ�ٶ66��[a�El�uZv�e�jn��W��6�Dlj�֯�������l^��f��Ku�yk*QWa]mç0TwA�3M:z��RS(����*i�h�)�L1 Z�V��*G(�����U���Y��ӊj9Ooc�V�w�U�q�yi�HE�Fԙ�/N���aŴ)"�:ZPu��iݰo+XD^�^�]˔X�Y�T��ښ*^ƍ��M�JYE
�N�����o(��l3�{M�MbW�40�&Z`�SZKK�ێ��Cu]"�Xin���wx%*\j���&��b�ƥ���ӈX&ƷY��i<�1�eX��%�5�qڌ���VO�<W�Y�>#i�J�0fIa*�or��m�������] �8�.E��Ѵ%�W����e2CB�,)	�ZҤ���8�����(��f��ӭ@<�4�1��.-���7������B��b`��a,8f�Z]�=����v��*%F�mM�XxF��(�� �$�lSܫ8�"�֒�ݒ�dX���JX?���#R/r�v31����,�	��k�a�k0QE�G�E����ҧ�Z��ʺ��<��i��
M#H�L��-���ݥ�$�9[{.�4ƫ3f�F�v�55�Em����L<E�E
�J�d2jݚċ7��)�a[�y�bE�6�{���w+h�D���w���F{I�x5��wQ�Z��ʽ[��b��)��ˇ.�KE�+�����u�<B�����]�v0���"d$�wL�FVciQtL�S6Ln�,�Q�0L���yp��f�u�Rb �aF7rb���fĆVUڲ���v���(�܂8�ڽ��T�{Q�f�V^d�& � 6vJR���l�Ն M�feS	TB�4�m�j��Z�PF�5�I8wb�I���`���#��Zg30ǚ���tb�G[��Ayan=4̓[nz('���`!�iN�a�QZ)'�&� ��T�2�&o5���y�q^�x58
� ���Ҵ4>��%R�Q��tj����*7D�n��u�mh�*h��z��NYժ�D�����+Q�uh��E�|�����du+2��#�^��V7��na	Xj<{xι,]ܽh9beb�9h3Z�V+)<̬ʻPI*K���f[.��܌3R�]�����S�l䢵ښ��b V�
)���8�a�V��@���Xw%m���d�ZyN�ĕm��"�Xٷu�n-uaDſ)Q���dwxT�V�4'~��x%��n�x c�K��\wiгY��V��8��ڽ��z^��h�b@ �+%�'`�<��X���]�m37Qe��.�k�s��r^R�#e�6@v8n"͖�`��(�7�#U, A���f
�й6��!K�{�1&�^V�8�C9���*8�E֪8^�ӛ���8�S�5��i��*r�V����WVf�ບ�4���nn�K4:��Q=Ӳ�$�6Gt�p�U&�W���&�0�:�-)B��W�����V.��R��N������+��W�.���9	�`]c����PCW}��d�E-�+���꾓]��}.��������S�b�ꁅr��C:��VR��s�V���r�����+%蚍�{�Ћ8K-�pŦ��u��Wb�q����@ɇ���6UD3_e��ĂwGrSpt4��U]����h�
¤�@ǯ\��
|���Y�v��]I�.tWH�S��u��lͫ�%��o-$;	}��v����#�n�Cr�6p�5�B&;k�4D�ݑ��sa�he�Qٻ��6<�q�Di͝)���B�=fGQ�ڴ�ԮC+P���8��b�X�}��%������m�i���Uv�;ƶpa Ռ���K�6;bL�Rov͉\֎-�˾���y�MM�6�N�aJM�X���D���Da��	�ٗ�4�U��o�7��9����De��-.��@�ĭϳ7�>�q)[؜slZbu����7sd�5F�&q0e���i�Y�u�/����5Ӊ󦶑H�Gu�؈���A��}E�D�.��mk���d��\B\�����P
�<&��^A'%��Kw��t��؞mΒ�፧�i�Ś�kG�AAWJ����O�y�k:ۮ�h@.A��%�|;o/2�s���t{[���aacN���9^٬Gr��ܚ�=WM�{�(�K�,�7�wZ|��eb���N����*VFU<ݗ��]�r�x����m���&iq_N�2��%�	�cj�N������ulΥ�`+2-�ϴ�lm�f7�ң�����ʚ/�o+���P���0�G�oZ��Xl�ɪ�n�jڙ��
�:����!4��N���AF�*jS;���6��f��[ͫ{��G*l�'Zٛ��]q�л����,X˚o%M=tj.��-��sɲ�)p]@b���x�J�ڪ_hdM�[��V���k�}�Xkԓ����m�A�P���M�h�yr�LO���9FN?��SiF7��Irogo�� j_��E\��7�'c����l5���"ov:�����`Nt��+��������<{�-S�3�e��[}��w�1�]2�
ᗖ�$�
d�n���5����x!�n��s\ra�l�ԇ�]��q��`�kn��m`��"����R�t��A�R����C!n�wI���d��۬�s��QdCzoI9]W؂�|s2������Ux[���Rr��M}QQ����?v�x+�->���u�<�}&�D3;�W:��픯�¬T������ �w�ä�,s,RP�|se�1�t#���9y�ԛ��\�>�]�5���j�X{w�z�O4�b1e�{�Fy�Z�Չ��r뭽˩��{]��b��>�Yˁ��Mm�N���D_XX4��$�����U8u��*ZQ湻td�ƕ;�o\�u�l9�&;���K��xp�g,��3L�t�"f1��0V�4��#�]�DR$ۇZ�a�`t�o��aë��6ٓ�W1B��S��Uk��B�WV��w�cq���+�z�s��˨?��q����կ)��}ڊˍЊ9��C3�K�0�;�Q���zK���]����({�b�����ܨ��� ւ�I�����wh��|`�7/I�g#�ӭ!ם�mhֶRʥfe�m�5���lf	���3�ˡ{#s�v��e#`T��Hz�X���ݡӉE�ۗ��nJ�����_-�Z�t.��b��(�r}٣@ׇ��ͥJ#-��	y_wE�)s����.�6�ݮup<�}���\�\V] 8"���C{�
��f�a�9C�`][���S@��������n�.}0l�g>��Bu�ó�ą��'.=/jX�=�0u^�d^N��Hy3oZǷָ
�%��<9�

u*�nw7��Mb����*_,�4��_g�������X�2wN�9o�.uo��2����uՃvA�s��ݚ��ˏ����Z�g��b5�R%�*��ؾ���M����3`�����1��unM�Y�EW+��N�»��ջ��s�jL4i�ˆ޽�[����@�b�xal�CAP��Jȕ����fГ2<�)���~ E�س;(�,��o9�ŇD:�۔�A9�e��<���G�kL�:�����'�z���ѩ�լ�]0�u�-V��<�]��\}s³�#T8�f�gCP��ZbL�p�5e�N�O�d"��tl`�Z��(]���`�\����J���mm{ԧ��A� �ѥG5
J��|���w�����z���siP���r�64�S�;��'�������ܵ3�靴�Ҷ½�(>��xB�m61��u\�ãY7��#�*��Q�T�MgB.�sx�����*,�/�09O/���d��u�9�\��]��\��˴+���uYLj�e���v���b��"+�ee�trX�
�}�\�%t���{�n��!�^K<�y`��%�/��\���YF��U�u����Z�+�w�8<�*��$53X���v�5l9/�PSv�V�wŞ4��n�[c`�ÖJ�:�tMCW���e2��k��&u���ڍ:գr�%mvV��$v��4�CS*u����"6�e�u�w.u$�2������w��.�^Sn�S<�,��Z��4���,�°�S7r�-�G��Mf�n�*�Δ�sT���D�|4���C\�t�٪Vrݮ8������ݿX��]�us6��V���C���Q�v�}�[O�Gl����`��Y�r Gf:8����¥�὇^��D0�u6��t�M	���c��tJo"�d"�q�b��Q�h�����v.c/��k�doL�Q��WƓ�H�mq�Y崺����)�@�\L�r�bc��Eq�#yY4���h�n�3�x����T��ö�)K�ާ��Mw���{ ��U�6�O���Ć�VG�hu�c�7]m����WD�@7��1�7��6SёΊ�h�ޞO2_Q:�$җ�,B�V"�/�[ڶ��I���I@�Z��V[�j�q��d�I���.�{j�w�W%�B���F�9FW7�h�|:I;7�h�T�=���ݼ�}�a�W��N<���x*)c6�M�Z����m��e�� �݂+��͢��@2�=���+g����:(�9�(*�Wי�Z����6����
�oJY�7v^l���i�KVŤu�r�M6ւ���;��c�=���+��u��H�L�|��^OyP�v����t��f�W+=ʑ�>yy�s���s�&7z����;� ��[��Ou�F��t]��j2E´�%ǡ��q87`��k&�o������}���c�uܴ�9ThV�t���eՃIwmf��F
�2��c�3LW"/f����۶(E�IV)���,���^�u	�StcV��A<Y��hC߅�˶x���ލT��ڞ�:����@��J���#���O���ӑH�Z�JV�Wh�X���d�D]f�Q��p���4f�`��71o5��v���t:�*�`H��xl�Ç���i���hY���Z¯MӤ,e��M�ꉭmK���ρ�*�vӄ��
������W��@>�ث�Z�]�\%�8�<�GB������.�i:.��e�5�H.M53��T����-w9ۑ���>Yo�����$�5a��d.���"���������\jഓ�^S�;���y׌�.h{�)֒�p����-A��눨��6�Kt<ݨ�gD��V�Re�R0�{�n��u��2�ħ���M�̭���k':�nf��k5�#մ��:7+�5�b�&�Y�>���DG��+M�Ng�����k��]a3��T���^�7ut��|�7���Q�����y��Q�����4%�(��֥r���:OG��@�)�P�]���;��,�*�>�c�Pyk��[���������
�+��©���[� ��u�\���(�|b�V-�w]�!�l���ʷ��,����b�rN!ǘt>���	R��f�K̬�`�h<���\k��~Z����e��C�v����l]�4���$h}�'}Z(�<�-r'Q��q�#l��P눶˼1$��=���}�x�{f+���!��T�"o+�G ����J�5QZ%<�,��D����W����s���9�n^f%j�N�ƙb���dbZ���K�(�Y;}�|x���Hq��xM��\�,��yK��5��%��4�Y�n���]��c��4)um������e'��bfmu/�YZ��u�P�&,�R��;PQ�}D5�Qte՜�MC@� ޘo�� ֩���V�����	�`捭�}��p]��U�|\)��W�b��%��Ybj�6��[�t��}t{�
�:
٫�W���s�0��U/n
���`���ꄭѽ��}L>�u��T�r��Ν�R׽�� ��r����k�-��>
�!�X�ub���J��52�+���Su��j��M�7K��AK0me�J��YE>}�� �*Z�H��;Ei�E��B&P0XrӫÃ�<=�cJe���G��u��X��Q�[�H��w�vbWK=i�����Y���/mre��$�������T�_+��T��2�_^i�9Hk4���(��c�����hU�+tW.(!�$�N�R��m�aA%��{���/�IX�8+�o��rݤy\�0�6�N�(Q�c�D΀X6��X���kk+���I�¸��i�w��k�̑h� �����J�ך���q��A�ˤ�k�Dκ%���BԜ��ـ����N�\wn���Wm)��������De��"��k�Gj�ņ{�x�������ĝ��ˏM�y��VLZ�2�;�y��d;��߮��S�j�L:xN�Y��|@k9P�����UrN��X�Kv|�ˀ�e�*�<�e�)���iA�OVs��;]�mQ�6�
weVi�=�z��^��s��z!�A�7�@&���G�	������nPIf�!|ge�&w,��֗V�`��R��,oH�[zk�6�k����a�[��&�6n`���|�朹�ϻ=J͎��jjv��\n]ˮ�ǻb���q4���XM�w�W��l#�7:3�;ie�:I�g;�9\���=���t���Kxf
�v���9u�/����c�)=D��3Q��e�8��Y�s�U��%m.�u��qN8S�}յ�%��˳0���ä���Z�Dg8��Q�ڟ(vRVmbG���qƮ+w+{��pW}Q�&�K�A��t��oCQ.TR:Pܤ�n��ڎ�[��eN�2E�0f�=w�@nJP*�h��#�N��W..�0�t$N#�/9�}:�f�X4Թ_{R�]�W�x<�+|��o)����nh�4%���fcƱ=��1-h;�j��W̩W���l�xۭGd{ٌ����Z���t����k�/��yϴ�4l������8@_E*�F��0򃻄����`R���.�r�ABPw�^���N{�����H�1f�vT��cf3h���mBu��ۚ��������9��&1\�a�j�؃ۯU���@���b"�E�u�k�eZV�ӆL��2�n��k��|��Mƣ�v��&�j=�|{6٬c�8�qӺgS nu%L�t�ѥv{V+};���i�Ҧە�{��rnYh�1��]lO���09^��t]B�f�7��&�:TD]�Ԩf�P�۵}jn��Q�A���訴78�4igzmѡ��T�Y�ǻ'$��}�j7�M6&�JY�D��,��:�{���t+uK��	\��.ʎ��q���۳�)fZ1cq,������w�{Ʈ92�tٛ��5+�>uº�q`}3lf^���p�B_,/Mw9n�r"���B���R��,�O�U�:E�mTOy����O;6�����+ﺭVC�6�r��ne7S����ٱ��玔�+Xkx�k*Ty2�r���x���#w�7�k�U�\P�z�IڲLH�c��`^�66)򣔆ܕ8��Zy�J����Y��UIɋ�CLU����\�]���;�焁yM'n��wα��AP�}:�7�/��}{jmu�9y�x�Y��Y���#K.q{Sm����J�)�\��1@X�k���kz��euN���B6��|c���c���כ��y;N�:�mnp�v�.�CSݺ�>��h[R)'%4��j�N��T|�L���C�O�L]>�%�Е���-m5wrG���%���N�$���v;��陬n^D9(ِw١����7����.�췝��1�21YWR��	務� �ku�i��/��(����ܤ��E�601#����)�77|��t�����fr7\햣x�K���Wn�i��[7I����f�yb��g(� ��>�YH��/�`V�{�gu���h�ϊ��f�F��yJ1�x��z�Q*��e?���]���>��+���8!n��*�&owÅ7W��T��c�(,���6T<��(v4L��#��FK��a��ud��(l�[٫ /"+�o�4�D�O%�s&�[���%
��"4��.�m'}X��ְ��Y9"k	�����7Z����)"+��}�%5���ʺ��&N�緻,�=�q�h��2��N�E-�k�;����)D�47z�Ԇ����f1'G9��"�d�M��ٷ]��rW�Dxnk���/�u��q���g54�哶����M:X���55����K�܆r�iҨ��U�k.���@�]�+J:�N��7P�靝�(��m�]�p�*�6������S�8��(��w��������-Z��������������|��>��0���NbrĆ���.�0�ciQT7..�����3�j<�:Qu��Y�� ��3e��ScYA��G�X�`gx��p�9-p��f%
-`R�M�=��Ӂ�ʙ0NA��ݴ*!�!�.�,��Y�m��ÍG�<�(�S�z�
ӡ��Ks{~�3��25-^v��ݬ�j�1��6HT�aLt\��uCݡ]��rP�Upl� �|��r��e�W �s�GC�-�K��SZOWVw1��K˨Z�i�W  xY��U3���V�&j�7R��ʳ���]	��I=Y9{�X�WkOiGnͩ@$h�4�g:��C�(��̑六�($j��ݕu����i���{,'e:��Vd���h7.�˝��	��؛&u�{Vb�@��%��۰@z.}�w�v�)��L(��+*�jxj��%V��=qt�D�tؑ��wr�1s7��[���e���ȍ˹Іd������z��"l�6��(�F��3soZ� -�r�y.�೚��2�`،����[���T�V��^U�t1Վ�*�@�joa&��9���.�<u��.F;�i\�p!]I���wN��:l��dW>-���wI�QP��k��\ʅm*T,�wRL���o�(�w1'�ZY��=@^��9��֙2���QN�*t\�f�e��mїy ��}3{���u ;���'���o�p`�Kز���Y�q�)>��q� �T��R��N��AL��K� *_70r;e��^1u��P(C�뾼�^����|Wk�RP�ˡ[9�`=}���N wt��\�}إ�m[����V-%�����vb�F�ɓw'#�1�F�]�jq_�G4�)�aX��+�z눢���m���ҵ�^�"ꝯ�:�ӛ��� {�v�Ѕt�!�sy��=�Ѳ���Oq�ec|����/%�� �PF�%��n��V�`�]�	7y��*5zXޮ[.����s-�N���2��:C��v��2�QVНl_;)m����>�����Q}Ӭ�7��ئZ�ib��6ؓu��m�x2�Wtwř��=���Cq)��h�[���':� J�Q�{mQד��,ۮKom��	�s�K�\�}Ok�&VVuH6��+e�P���u���)uN����(i��AC3]ս ����Ŋ��	�d�����X��qT�Q�����[�R�j�V��Q|�[wwR-���au���p�N1.������ż9�+����9v�w���� u���?v��{s1tC k�����"a�O����Ml�9��U��7ЪJ���1n� Ք�E"�|7����2���0����Ֆsh\�c�t���n�M�/l��6 L�,�PM]�q8���WCW�x#&���[��us\:�q[Ń����[��qN��wM�����ыk2��vj�ݝc����=��|�&��J��A�s��p��:�iqٲ��"p�s��!�V����ef�q�M���6��+�&p"�Tr�Y���W���j��-�y��̙l�Ω	X�S=�J����/a��a\��pn��!Z�lS�9��L�(m�m�i���A{]��a��η���w��N�Ӎ�.�I[���IP� s�h֊h�w�n+3��L\vR���Ԧ /�����M.�\.�ltЩ	��|\G��FxR���������۪�q�u�!����ǂ&j���U��A+��oljV0�n�Nd�6�t�m��c�C���Gb���or���{z��E�x��p�������z�"�˻]t͆u��ea��Tz��}�_rռ��b�������GDSn��y���9�]�5��v_.<�j��qCiT�E�5��A���W9r�i�E��y���=g4+�ZEƶz����+8$�����m�B�:�8��T9S(����JC��p����N��7��K��<����5�Q�ъ��P��识v�a�T:�ؙN6Y�/F��b��e�:k�;H��)Dm�������Avq�eJ뭴둭kt�ޥ:��ܱ��=��I�|`��]v�a����7���ru_�8R0m��%�϶枑:`�.�h��&[v]�J������V�m]�=�pr.�D���v�Z�jThm�,4!	p��rd��F�<y�>�R�kμ�N�b$�Y�1@�՝����'Q� (���G��Վ�
���iyX��3
�c��������Pi�1�Z�bn
�hl�Kl%L���$M״*�K� �뱯�E�dC����B�,*W�a��m%I����MT���_g)
t�
u��cQ�k&������Y8oZ}�.b�NR7�9�'�V�%n�n�������+�7]\�����ی�V��,t<�YfbZuj����IJd:ޟK���M�7J��>�h��=��0�\��h���4d��/������]G���.��n��[u��*p.�Pn*�5ݹZ#���"7����J0��݁�.�8ޕ�]�����ڳ�L�EE��Q-K�NJxj����ؕ�cσ���������(z�,�=O]�G{�3Z�.�jά8$���WC{��5�w��A�>� jg"�hHqr�j��Vp�Ksi%A]��f���}zI�F�:��z�	�������z�ЭY�y�B�+x�:a�%B��K8YϳUY[h��@���l�i%�K�L�FɝR����廊A7h-Ov���Y�����bc��F=ݷ@
ȴc�4���SjRvH9E7&V���v�a��ӪC�hu����z*�3�I�L���\��t��hXJR�Rd�-p՗ص�j���i���k
��������-�hE���I2��ӵ6�y6�����,�:��4Ymfp���GD�,���7Guv�h01�D�Xͮ�ͽ��CtJEA
Ը�[n�T*�8g^��!��5�Zf�!Aԃ�\�8e�m�Q5$ݖ�C{�Es��K���Y����F�;8�ڦQ��+�}��Y���� �[�	��(÷ٰ����T��݃-}��r��Ľhm��lh��ڲ��䁂�t�:�X�w%��"�'F�'s�&�� 3(K�j�7���i�� �N��ު�2v�M�H_C��)C�s�[�S����_1f����(,�Lo7K.X^m��	h͏��8J:�����tf�J��s-5���|�^՝�D���-\���*�|�2�L�N�%�k�m��3�-;���x�3yX��Xy�]v��ݺ-r7�fc���1+�|H�� �^�f�-��ɻN��2�R�ɬU�+�giB �Vu��Mwi��ǋ��s�e*��_VN٪Sшۀkk9a��.J�+=׹��N�
ʻM�����$ e�m��^Q{�)��i@�����&����Ɲ�ؾ���!�V�8�&_]�)W9_[���e.�2�b�K$�Q�]��\A���̑�tn�6�a�d����ŲUt�w3(��я�h�@^	�������M�j���u��z��)V���=+�ʂ0�&V_[8���+���Ѥf�f��Ko.��6��/�g�r���*jg�p���Sv�Z�+M�)P`[}��!�C�O��J]Y�e6u�ȥV�EX��v�^)Μ"��Em��R%��@\�0�Rގ�yA��6�u!g�m!}�-�L�"R��G��H�㖶G>��Q������d���n ���G/q�E�PӴ�\ݾ/�-=}�^�2n
[�:K��^uu �1і�v��Ƭ�����L�]�ce��6�
>�;����J�w�o*5R���,�ë%oJ��:�$�:�M�-�ĭ������I�m��ar��u֧6�G��'\kX��V��G��1v��v1���ߦ�UgQ�kD��k;7�����,^D� st�o<�&��O�չb��F�����|�{� in���tFYCWəZA�8�ˣoo^���|�6����8L��JO*��I�K'5[��F�lh�jM���/u^A�i��gB�ww�"U���2w��i;OE$E���XH���R`8QK]��;��]�=;B��w��j����32��a}ҥ<r��[O��vͶ_�\\� +��]��E���͠��z�2�Ê#d>�z�,�u���Y-��ԙ�K������v32P�v�u��,�l�ԱJwX��
�ʧ�%�ף2������uF^���c��<$U�t��v�w�L���6 ��IZ�½��3/nF�%C�-W4����`Oc٧5�
��<��ӥ[�Չq;���Y)'J4pe��]���	�n�1v,,6�4�p�2�/>�m��-�z؂��!	=�U��� �Xee]�;ړ|��J��ݡ
��ҹMWT��8w�$�3s�nPصӐ��˒$w�s��Ƨ<��c�15Y6Mu'׻�:��K�חn;�ld$_k�R��Mj
q��%%�ڽD�Z4%<��} Y��[��VL7�O_A��ˢi�wy(��(g^��F��w!o��a>�kz��.��w,����"۲+�5d����8�\#�i�y�����S]��2��#�@��v7��T�0��WY&Nr�4��ם�m���-��0��;z�ZIB���e;�VJ���;�I�����.^���IB��m����x��3N�=�9����0�J�A>"벘w0���.��M$��z�sK���]�����BM�Xɬ���YV�r�ډ`ɭ1]���r5F��Yk�i�l����J����.7��c�Q�lT��g7{��J�f��Co)�(;�[�!�j�lL83v�N+|o�|&���4��:�t����6RX�'�/-�KiM���������aû%;|��c��gvHU�P���/�V>�}zc�ھ�D��і{~�6Nm�s4�����sㇷ~��u��2X/;�Ř:vZ�>�o����0G
F΋�]9l��vn������9p��g]�GJ�{j����-�챵�gn1�[��t�Z�\���kP�hKQu�;m��f����N�Y��U�@B�\r.ۺ|����]5p����RPX�jUʚ�vwC�:�lv��X�`�Jdld��5���z��}{V��āt!��[�/�o��I����k\�V.��w�Oht�V�Uw%��c���]n��\�X�-�~�k$����7���W6vC�����`a���t������{�Z��eҺ�Z�<�t_'�^C۶�:�RV]T5����vpQ�]����o�r��\�n_��g�(89� -n'��̮�A�7M�hi�BR���剁�_Y��ބ`�`�@������ҕ��
���3���N��wu÷"H�N%��=�,�m;`�	 g'
��Q5n�8[�]ذݷk�Yg�ojƧ���0�J�{Yn���'�҆j��E�uȸƖ�a�͆�7'i|��^�V�kP]o���y�Io�$�z�n���gu,�8�G���!��;�S�7t�R'�=���	=c%Α	'��ˤ�Ӌ�@\��(�eعq��m�JyL5�[�6j=�Etwn���{��)TSb�T� 8����=�d�c(\Ovk�z����{�G\��v�{Z�X�/�to�hѺE����[�O+e�M>1�w�F��Ӽ�v)������]cRe�䢫��K=2��]x)�[|��Uj�e�sy$�b�9�r�moX�W���v��3�pQ�QF��7���3�+SU����K�������S���#���g7tRg�ud�{$��@q.���<��{�Xz�����ы#e����N�8:��@fQ溺u�:!��iYk�y.�2�2�JnRs�X�)�>ˬ��e�b�w������W	���{v�:HCR�&�e�x�gI�nT�oT��e����:�+e�6ږ���W�W�S:gWG#<�⤺�r�a�ă��l���-�-Ԧ��n�Q3��5 ��ܴe�K��F�+ubp<3[�����a��h8o+*g!y��i��G{��:+15��k�\�q�,�;��kn��t���Uv>��c5F�>Z��+���]�/{P��gvjdq5�H�-�}�G3��u�{t���ΎSs���!�5�a�0�u�7�La��GsSV�j�C`_-��Mc.���>`�u��fڥ]W��P�
�h^�N�����%b���V4�9�M��d��2��1I2����i���3��e�ʱ[��pM�Ƴ����v���L�1X��j��&�n�1[���-�Ǜ��
C�<Tm���fn����]fWA��X㙶��hΧ�:��V(���iRnbc���t:�鎍ڴq�$�*W
S&�W���w�vl�OU]��^�3�u�1�VS���o�p�q�ʙ¬8�k}��l�S.��<�ki]��Vg���LQ��B����}8��[Ʒ*��hϜ��l��È��O���T�,�3�ذ���r�i�pEʆF�2�m��{�̮��sq���oa�l����L,��fq���-�!�4���:�|�t��_.@KGw:�|#�ϖY�.�T���}�0e��a�0�җ7ͧ׈�WAKX���koK�nT{)Gc�2�	�gO1�c�����ڍ+���@j]����tRS���J�=x��A�8��.�]�����``���W+�6؜%�}ip4�]�/�^�:x��iU3���X�8�zʦRaޚ�V-F1��]�ˬnᔭ�i�I��'D2��Ky}��=hq��C*�֞���,m���]� 1n5[&8���:"�T�5a}u;�8i�u�.�)uj���[G_'vs�«&�P{ۼa��%�Cz!N�\����=��ϝG��r|V]E�oogfr�g�%���a�{�`s,��b�\��.��c�⨨K�9]ܴ�#��u}s��:��N�`f��քN��:k���_/f�
���c�j��?ʫﾯ�����f�vr{�=ݙq-	�1|��-�k�o,�ծ�1E@��Rۇ�.�3��ɵ{��������ʙ!�F����ΰ��X���Ao	��R�NZ�;��W�ty��h�M4�qSa`���ɩov�Y��]��r�M�<pb�Mx;�5�9�tsNb��� ,ަ����nQ�3	�J�KN����63�jD�W�n�[Ӻe�w�+����(3�h�s6E:.yɋˀ�]\e�.P�a��"�oD�3gF�$��Y�9g&n�V��A��q�'A�\<�i�ͱh�pIL�gQw��]ôL�0 ���pWf�!���h^�g������j�𵢶/i>��Eՙ>���ٜ� �j�4��i�Ci_.�񋏫fP��#6'}��;�'A�5�\�cG5�U�b��脠s�ϐ-C��~�u�F�in�N���S�2S.�^���>��7���L�#:�����Ҧg3-�u�}[Vrf��zؤ����眈�G�'ǭC�Ԉ��H�f�L�jRB��?�쮈�Y���r7zW$�<��e]-��m�ڗ�jq�N��;��O"��ޒs�X�a�n�8z���1�S�skPG���d��4Q�+�Q�W�BU��0a.��jdz;�O��y�!�h]GH�7����;�:�r�B��ֽ��fM�VAŽ���gj��T�U���Eψ7�v�ks�Ko�F��>�@� �F ��ݱRnm�\�wZ��b*E1�Dh� wk��v�(����`$��$`�$��d1�ED�#�l�2\�b4��R�v(�ݤ����LR��&l"H�2Q�K���Ln뀜��E��\��0�Wwh�u��;�#F��s��h��t�5�3wv�h�J4��Lwnwn53I�(Lc�u#X�!6�JCd�Ts6 ���664�Ib$ۛr�P�Wv��$�(1DW9�\�"��P2K�r3��`��I��HCF��@wu̉)���n����҂wraL�E2
~m�y��~~����5x�TF���e%ԕ0R����7�8�R�)��=v:��7��;�P���A�a�u&:铩��|�+����t}���hÕG�l�\"�ڗYI�4d��m�X�%�nb�M��%R=Xp\Y�<��`����Jz�����f�zX���}�u:��7w�B1ݞ��0<��_+�ع�y�JC^�}F.���/;�'y�l �B�_�^��g��s����N+��tĬ���)�X�u�EB�r�W���N ��곽��ل��m��UZ>�I�3��i�Zխ1zsΊ�tC��n]<�B�Q��=B���ٔ�p!�g�M砌�_��V��O�^�� ?O=��xrw(���u�{�� <Zǈ@F~��߇^A�>@{ec��pf��y7��YMN�Оw�w�.��'���>_vF6�-$�#�YZ�#^��u
r��Xy�9��7�/&�*�K�\�VP?h�p���Q{��]v=���5�I�p
���i���5н�y<��Gr���v�F_ͻzR%���4BP��`#L�Ұ3�B' T5h3i�Rm�U�v�p���f�A��`�T|:ERh� uY��Gmd��t���"�Wx@O���8i-��R�[�vWL����F���+��q��&�G:��e%�-p�z�v��M�dC���#p޴%A2��5u����jT8�|dݴo�b}}{��]��*�J��{����k��20����T'P�8ۙgaA�hC���]��{s;�iZP}@Հ�䦰"�Ή)u�a[��	�q8���{��h+8��Z�h��S�{��9&�@݂�܁�����θ!
��V�w<�/��MW<�o%����Ht�V�(�!��� 7S����_^}����_N��<�o'{�R�kuJh��u��S�`�sw�P"�H���=���k�q������ϔ�S��Z�*�(����D�e2d�ɺ�|h~�9�[<nX�.�;"60���P��dK��O�݀#�)�zk�W�!'wF.1�Ț�����ь�o��(T-Wb����`�'����<:�m�]s¤
��N���c��m��w�?Z�%{Ҟ�o�%a��m'Gz/�C|_U� ��\��@ݚ��v�<,[������8�T��s�x�Sd�R*gF�ݾ�OC����.1w�y�;�EWY��RcI�O\L �}lb��`d
4�qzj�[��'�X�.i�`��Z�au��B4���\��d!-��-m��S�֪��(��O5w4�X��\F�4X\�ʃ�6���1��wQ�N��h�Z�Eڵ��t���j�a3�t8��;�w�<�-�!�s6�-�q�m�S���e��y�>����^�5S����Ho��;��h��TW{*-'г�.O@1S%����"�˧x������f3n�B���¬�0�gB�_L,�):�y�*Ӊ��L�3:�
�yˣp��V}M_�3�|ܡ���Q�;U	{u�fP��߰_R�B
�Ԕz%6�y]��
��鏯�p�f8�T-X�ק :ĔȜ�vY�Z�SXT�$ߨ�~<%4����������������5/�q���@Z��γ&)����%r�ñ�0}[�k(3��g˸ʦ���zR���h������%��^�&{8�P4��n`��4���͢ ���:��]�]��nϕ4�u8spj�Nz�坊P�+�བ��{Ѝ�������ִ{T$
#��%ic%�z�W§@���\�sl��������1��s6�P� ��9���ͺA�Dv���������rI�7
t�/�n����o�M���Rb�$�Ɉ��FE'B��<�E�y/s�̥�*h���.	�j�)kǉضh��<r8��y;��S=�����ȇ{���h�I;Ձv�Z�0(�vܾd:�o�E�;���uq��� }��/���LVR�ܩlb�34@2�]yn��
�S��c�S&�'1���ݩ�[j�g�z���ފq;�.T�4!��w�	*��2����S�	׽���㷥w"�M��������^4>�Z:�̽�WE5���󂯼���]xr"\�f�����P�"k8�^��[B�g�']����վ`֊WJ����g�gk[���#������9���ڠ!�K�vὼ������jdX�/Anx�:v�x�3x���.օn��h�bBo.;>u5ȁ�%�F۪�ok7�b�Ɖ�c8r�����[`wg-xS�;ٞ��.��d��zP����뙀��b{p�6~�����;�Ѻ�;L�'����� vrD��QBpȇ�#��d�}�T���b1ܶ{>�\d��Y�J�xvl���=#8���]�?v�TV�	M/i��έ!�eY�K�k��c�6,O(g_r��ōȵTo���1��85�<I�?A�>0���n*e�G"̏�"���%Tq��W���Ŷ�g �)�˶��]7�*��?y� s�����x	�C	�<S$K����I�|;��F��M��|�M�WKnD6�7�te��6O�M^6�2g�7������s��������8Q]��JV�c䈄ǵ�}�6e�Ƴ�l"����=m҇�٬rTXe_P뫬��;�/8���M��3�B1C#������+}ԽIp�3�U��s�
�x�F[��T3�D(J_L�����Td��%b��#�+;!�XF�W!�b��y�f0�Ҵ�71�*-�������
��]B�g����!�>Mz'�7�X:�{�kvh]9�2�������-�,�-����uSY[�o��V�'���g	"��F���P�4��;ݹ\@\���7\K�e��FZQY�:���k8wwuYZ�Vy���Y�ZQ=�Q����g�N��
Uy�.���}��Ք\�55�Lʁ�	
&2}��CAo�y����(=)��2��.���|��p��qĔ)�.�F?�W|u��p1#j�q��L�Ø8(tY�6-OW+���J�T�e4	&I��Ʒ//�ޘ\c��V��_���U�3�V�׆���W���ĆF7W��.�l��T��%N�������b��_Г�g#\�<�������[=}�3S��Cuݽ����QU�
�<8����F}g���A���V�۴�E�o��,��|+b�a8�D=Xy�] ���2���_Dv�SEwRfS��]QNu��_C/�ѹ�wyQ�AG}"�"c,nA��V��IXެYfV��������W}�e�v]`V��ѽB��>X��Jç�.�U��[�v�l�r�l�,�ZLM��r�ց���"u$�"9��ӫ_��|���_@����-.� =��c����͗�<����I�2�
g�/��;�dcn�-$�#�YZ�t�{K�]Cx�>���`��XQ��]�W�U ?p�m�6b�Z�7%d�*���5>gA'ZX�{]r$h�_��88u�]��2��T:�J3X��9�RYzph�6�WYSl�G�JH!�%�Q#[��=/;'��/�X:�bI�gi*��H����i���(��-�mz�ƭ���m7�nǱ����k�v�k �{S�xR���W��ḝwx��ҕ���aJl����{ly�D����.��� 0*)PL`j������ա�^W3��1�_��3��yJ��{yX�:�ϒ�8h�;N|H¾=��{Ne�2nK��4��~׎�nw87"�.K��y``�B����6�����"���קs�=cx�5s�:�ε��dMQ'ƾ�k�$T%)�&�7@s��@z�`*�8<�_�/
t0@�� 3k��[��.�O��N׳��;Ja����\b�k���6���e����5���3 ٬=�OU �;o;G���שu�r�ٟr���JI�7;8��IS�\5�Sݧ�Wp<���Cxn-��*�_� ��2���3��u�k����r��oR����5^���4�s��H�J�/���^��W�1�|ŐѦ��0��ߜs��~�k�����@�~W�Sv����~۫�;��W�ޔ����w!�g��w����X��N?�O�@�ra�І�H1_n]Bpv������<޽���)�)����`����ϟiݳ��$�^!����R���<9]w`�C����ڠ�1����R��PC{�!=�p����ע����Hm{P���`֊�AQ��9���J�*>Nx�8�x����T��t�f�wV5[G�E�4��K)է��xn -���;�2���C�uFP*"YtS-����z�Z�k�κ�`�|�27<�e���P�Ǜ]���&+�?�����sMT=������0q��p1RDS��q�X�t�F�pt�Ѿ��,�"�K.!�-��!�F�!c�5t2z�#bՌ��j*��<�S��(/��0��(��Z�zR�.�Z+|�ٜ�3r��Bm�	H�8v����1�B)��K~����,���:NNr����[i4����4cx�i��}2�գ����<�٬�}�Z�y1$	ׁ�H�t��)���[3��������B8ސ��oox=�-�ĈUz�p�蝄;�I��v�iA���ݸ�3�&8'�w�^\ ���A�]�®���xn�2�];T=^S�޳�*��ԙ�.pBG"�`6��:��X��<<kG�J$��EXWiv�2�frSo>R��Čhm�}V���r�h�c�0ɮ'�N�iUD���}=��P�yr�5r�B;~��N�TTal�guHV��I�䝖q��c��2+��Y�\\3E��7e-�nkd��}�}���i��V"���>5�'9��ZJ��!L�r��[,�����㔃`/�8N.�Wѫ,��p,���vc<+�+�qp�������Fg{Wj�z4�W�1�x�YU��hVx�w(=�|st���#X��̷�1��8��y(F��KC%��c�bw���4?\ċ�� �C��f�];o�wJ7����Rd�p�A��ێ�3Ȁ��Ƣ���jq�W�(S����0�������������ޭ������%��\Gj�<����3;l��������:'��-���M�뺫�KWʴZ��)o���^`PU}+iK��n޷��=�h���3x�z�u��f.�~
/ALߩ�)jG���D��$�t|���֭��Cﲊy��U��������.C��ylmJ��;p'3�k߻_kݨ��q+��Ƿ�"�S"��eB��U��Y�)�b�.C�ϭ1�zP�,FD;��dS������Y3��8���Z9J�5�v֟C@V����+_����\�!�e�t�gR���3�+��]�<Ʀ�Lĝn��M˺�8��g�!�QFR7�L���#��'R���GΧc���ji�{�� :��-Խs�`0��� �M��$Cl�r��ʎ�}����)"��Y[��e��q�a��!���ԋm>;�����Β�o��8�ܿi���vd=,E�zo��}ݶc	�+N71�*ۨ;n�١p��Qԍ>�����}�M�GPL6~��1{ ��{O˓�_Ֆph�M��I���NdV�>��i�=��Z��f�G�ā��&���Y(:�;�Bs��y ��:FyX!jλ��;�%���A�`.������Q>��Mv�fS5�Y�k����=t|B�����n�����FWe0p#�@aOআ��ŘΡ��c�A��٭���c�/�е���-A ;js�o�}
����k�We�'v���z\��q��u6�-�{�Y�5Λ(����o��z*%gFtl�W��9���Rgf[�
X���e�x���h��2��WٴiI`N��w1b�f��#:1��I4A�q��T�vo!]��#B1�W|u9�c��y�r��ZRyP�Q���k�r�ol ��{ޭ�0��[�Y���������]�����@���W�:�wn��s�xZ���'�	��`N[�1UV��'\�k�g��kLM\m�b��Q�y�,7RjL��L�
����Ӊ�\|ʳ�M砍�O�}��|!o�8���ۚ�˽سӹǚ���Q����]t�|,a+l�� �ഷ�n/ +,����b��J��g_W�u�R��-�^z,e׻g���۪�I:Z=��Z�uH״�]Cxݳ*/��m�O�	��#\"�
������1KT��Ҷ�_ڕt��<	<�����;f�$��;�o�{�`�DXH��!,�Dbv��K/!MT1�M��L�(�RAm�ʕ�d�����N`l�k�u9�&9�J~*
E�k���9U�O���b���\��+4�N��*Qj��00��}5�
1|�D��W��V��']ď���M�\����o��^���Y����8r�Ǭ��뀅�G*7`l�]H�E�D1wW�d̮�Ҭ��(���wP+y$��:�Jf��F�zX *��]��Ő%J�P=u�`oes��iNA8
�NEƲ41˦h嶫���ڶ.? �T�P���-�=�V=�t���5�P�]b�S��\������2��ٚ��h
�-M,�S�6��س��&[�&�p°T�s��C�����yH����#{��в<s�E�<Uݎ�/jYp��ݠ�͕C��o|�n��ZtKn�i�X�0�dڍ����#/wE�
��p����j�Z]�ڢE� Uz����2�:�#$�9;�)h6(Mw�JY%qVm�c�Ȯ���װqeR[��Y�;W�%e7��Ҝls��`�:�l���q�X�0�af��o^,�B���! �ڥ���}��K\P/�m���[�C�[��	�phĳU�l�������L��詪(��w(b� ����x�Fޑ�W`�����ӻ�]��6Un����h'����/�{e>ǎA�PZ�z�����3����WXw6�vYs(�t�%����Q����	���aq��`.ٳ���º��ƞ�N��k����r��y��M̵kࣕ�DՋ\6C��W<������.t�}H,���b����l�J4Z�y�ν]w����%����[ث�Wd�j8�9с&�t�q2�������ھ�3q�x&��]�t���p��c��6㕕c{q=xpv�H��O��|٩�1u;"V�qY8�J����x�j¤�#B��[t��9C%pS� Z[o���{۰u�@��8B���>�/7�Q٫XwON�� Bv��|+*�4H��G�l͐�^���k٘"�����{N�lD1����ؙ���!�� �J���[� ��|)��y�q��ʃ#q@%�u�n�۝z7tm�t2�F+�q�m�4n,T�nU�����+�PM��8�iklf$s�6���ݎ!�R�n���-�E ���wEoj��K,��u�L
&
��Ƹ4��)K�Ѯ�]�� �=�����^=�f��;$	�.��l�42�c`���9����Ñ��1I>��L�F�ۦ4��y��v9��"Y�������h�1ncO(Nk����^�<��[������Գ��EQ��*�BWY}gBv�`����wn�yc�G��(p�gX-G�V�T�꡺�;�ٴ�F�Bͼ���w2�+��F��G�]z�9��Y%np�6���ioT�IX�۱��R�F�O��2E.q��<�{j�̏p�z��E�gh��F�.?��a��p�]s���R���U�7"�Ԫ�����'Q�8�l=�ڱ��]��ko�א�[���a�;	b�����"����Ti	��5� x��������;t*��}�	����cF'���-t��]H���Ŕ3@D[�����N��w.��s�d�`$�wn8[�b�˜J�W7�#L3�rn��AdĠF�AH`�0$)�d���&%&ff\݈�#��QJ��&Ċ Ƒ��6)�Q@a��$f�#�Q;�wt�4�1��21��!B(���
fb\�I��21���"�D1�3#	D�f�$�n��!$�b`nn�1JL#M�J3"fi0bh��I�pS�IB��-�62B�$ws"i�3&& Ѵ��c0��I.rL"R
���k��2P�C�BLDe ���h�ܻ#&��!d�I�J$�����5�R��[�N��v����z�ZR�]y�����x�G���7v,�Һ|#��CN�.YA�WLIV �N�U��-\���� �G�b'�ߚ�߫��^���5�����������^��J�so�sם|��{U˕�η��m�z�?^��:�6�F��>���DCD\B~��c�}�,�Ŀ��B��/5J���"D!� [��<ſU���/=�>���ͻ�}����~-��z�枻n|\���^
��|����yڼ���xޫϞ_Z�����[��W��5��-�~���o�s�_�sT]��w���I���"#}�Cn�}3�?|g全�*~���G�c��3S�����;��|�[�\��o�|���޵��>{�{_�}{zZ~;xۆ�?���:�5�j5��/����w���˸�YrS���߫}�r�`���PUX�g�!��_'_D��@ }�U�oJ�wϞz�����M�~_>����k������oj�˕���a�r���{ҽ��{�o���������r�0��S�{V>����`���}�}�xS���>@���_h��
�Q����;-�x׻����~�ţ|k��Ͼ�ƿ��h��~����x����ͽ}����_���+�W�Ϳ����ۿ{or�]�q��`_=�]m���jT�>�����j��������z��*�/~]6�x߭�{���W��o��U���B��#�Lqѳ_Qx}��>���_�F�|��޻�狖�}��
�9|�Fi��k��c�n��d>2*%�L}��{x�����5�����W�η��Ƽ_���������}�?Z�W�O�~^����6�^�����[w��U����_7�������Qo�����׭�<�u�H��┋��Y-���#�D��o���W���/M����������5�Ͼo����n��}����zo�W���h�U��>^u�k������z[�\������x�-��qW�}}G���H�6L�x�sP���~�W���߫{>��[���|ܯ�><X��"�ޯ�}���B�󟣇�>Cnk�����/���x6��׋~���W~���ڽ7�߯ߝzo���o������E��D��*l��;����j4�PO���K�^>5w�lno��|�or�޿��=om����W<�ޖ�����������������+�o��������m��6���ʿW������������0D���rX{93�1����XX�u�W����|�`f�}���b�Y�fr��o�5��jo�w�U˻���f!Յ�Lɼv��������<g>�>��NI�m��t8	]n��p�������{�cE���#��8f
�O���O�]���%]���/k���HY@�9�o:����_P���}�ׯ]���zZ=/���۟˛�~��5|r�߯�W��v��?�z�_Z�}[���|��M�}k��~���|_�E��Ϟn~������篝\�����տ2:��n�]�#*�f��I��?@����\�����;�����;?�o<�_�?�����^�o���6���oϞh�-���~_:�_ͿW����m�_������ҝ�y��W��>��X����_�忕�����u�W���{���W�s\Ӻ��m⯋�ﾽ-��D�"��>}��F��}�BE9������}�dG��Ex��H��i�!<eRu�|V�s�G�|Ĉ�z'��k�ſ^=���~7���o��W��צ��[������_ם�i�����>-�W.W7��|�m��ޗ��}��}k�h��@��]��B����}�BnEW�� p��>�D�~�#����5��~�{U˟�����߾�z[�������{]�szo>�^��ޟW�_76���s�����W�ξ|���	��Q?hc�
�>�+�}��T��n7�w�	@�z#��C����E����|������~�>��~�r���҈����'�~e��\�A��L_�����rޗ��ץ鷏>u�/M�^,�>#���� �/�GSXn�r�ë�E��M!�`�����2�}��R\+�	��}W�x�{�����x�o����zߍ���Ư�Ͼz[�\��r��U羷�x�|_۾��j�˚������~>��U�T�}TG�Q�U��V�1�����%!��""D|l�������"+޽��M����n{��|]��~����ﾑ1�����R���A1c�D}>�x�{��y|k��k���W��ז�������G�0�����R��Sç�h<Z<��W�|E�DDG���h�����!�_��+�*���T'妾��
��~u�m�o��ߞ�_�������7�������~�}�~-��~o�>z��~{�\����I��(E�G���T`�y�q=H����[wv����<��j�s����?:��;���k��^��4{^-��4�տ�E�믫z~����������W����׵_7�n�=y���AW�my=��`����KoEt\�>�)���zS�w�}�Ka��]u��P�)�q���8�,�,X�k�չC��)�(q����y]q��w�ޕb%�����z��Ԁ㲞��"Rt]��c��UP����ۈ_k��ӎp�I��]�G�gM�Vv'�A[�������߿~z�k�|y�������/�z����7��7������^��w���n^/�׾�?:�7�7��ο��/kF�������ֿ��ߞ��3?FL@��& ,ю-���������;L}b"Dy�+��`�� ��L��"�m�����W�r�}�]���ս�ھ�޻�~����~�������ͽ77�_��\�����=�y�ž���r�Q:c�#�>��~}D]�q5�߭��@����ƿ[����o���x�����u^����_�{Z}����z����or�������x���z^����5���G�1b"�0,FO���g��EAH}��>��;YK�jy_�����w����o�?�}����5���]�������s�����?��~�����تxA� Dt�hG��D��1�~m���Wּ_�{���\�o��/���p�����W��!�4-�uا�z[���+��ݳ�?W����W���׽w^z��m⯋���_[z���o{�o����ǟ�o���齶��o���y�h�۟�<�o�޼k�\7����#�$D!��^x�i#w��Ϝ�����o�~����+�_W�E��|W�{oM/�ߝ��\����i�U&�1��
#놘���Ç�!�\��zW-�����^���W���ߗ�}o��h��>���J�LW!'e����2��}��߭���~�����m����cQo�������W��������/�v��x׍��A�}_��i�����zo��x��߯/M����3�Ӟ�uޯ��|)$��q�9oj�}��ﭽ��~�ſo��W�:�����~~�����/����������_?����+�~E��W���O��/>v���wv�ϋ��޺���wW��x�DG� �ؘ�ಲ��򡹅�#��^-}��Z�7��׋���-����_U:��#�"2��h甑Q����SH�tH�PG ��o�;,�=�5�iZ@O|%��<*P�¾��ֽ�ٌ��Ҵ�71�ۘ9��٠��/�������un�h=r�G.%~�G���_^�3=�ʹ���G��Xw�>^E1�]��z�쓰�W���nr���TI�}�3G;����⨼�ҙ�N\����.���_|^nW ۂq[��K�ς@��M��++��J�+v�V������bU@�ؘ��0�\@(u|{Oʾ��3�ڲ�'rޒ_�r�;�|{�:��9}^�O�=Ek9��G�P@h�C���\<��nBs��+>�u[٭M�Jh�'�3<��W��L}_B��F㌒�������h�Zͥ��Dbt��p���-�qWS�ɺ�7��`a}���f���u�zU����-Yd�Ԫƫʾ�"���|������?g]B�UXo� 9�@��w�*��ZRyP�C�k-�ex�f��4�g�3��Rע�չ��=��;�2�]������}u���]�V:*Kj���9�;��k��&�T�j�ʦ����r� ��d!�
��}p��gY�w�����j���	T����]���U����U�g��
�<8���xc�{���례�1b˽aBK��N��	���������Ƙ����㊵��Z]>@{ec�1�b������+S��3�] ��rS[��u��]W�����%`�T2oۂ���m���oxwkJ-V���囫�'h�Ue:��ۈ;�X.�
���dC���>r���Fe,�<)ps��w�BC�R�$�6y+��V�Lt���z3:�#\fԊ����	��21���Zvw.R�;���p�xuƕ@TaBs'pً�Z�5Vs2��ق��`	����['/{�'�]��`�Cԡu=T�(��(p\S���-���!���T�/A�Q�Pz�^0i(����+��ׁ`�)����f�*���R,`�k]�w��*�K�OQ�r��|d�^]^6ht�}ma��@��O�� *8�ڝ��<�h��Q>���垻�%԰��Ӹ:be�ɘ,�D�H$�@Q�~��҆���GH�+�KϺ���J!�>��5�PBs���<箜��(ӔHy�1�ә]X�$���S��p'c���>5᪇&�u���0E���`�ʫL_��\h���1[��r�0zڸyd��n���������[��ԗT�JS&M�n��p���ϧ�߶b��Ϭ5t�*X~M�w�z�A!`��?dKu��%i���.N��[?q/����j�g9�IVf�G8�.x��"[4E���fJ
�y������e� ᚽ����!ۖ2d|�Tt�\����"W|˙�1j?pta̚7S��������;r��8g�vj�*e�t-CR�<�`v��I($��/F�S�/�3�y�y�6V4�>6�)�l�5n���$�*F1�����7Y5�˱����[�}ݮ�J��9�����*Dŉ�}���G<۬<�&�Z�X7f�SU�.��[���.:���ryz�Un=lN`��`����s�sWB����Gm)�$_�!���Ê���?;�E�:��qZ�������WZ��@\AA�]8��k'�c��58 �����1yK�hQ^��,4�W$��s�ё�lt�7�s#>�LC�ٌ�n�
ƫh�'�5�3���܏�v���bz�^^�S����ªA�K.�e�ʚ���Ǉ%Yf]Sq���DR�����A�V�t
�N����Ɋ�����9B�A`#�M����ۭ��'kq)�1�A�q�ՆǇ$�QX�}��iW�Ѿ}�������bW�-����]��
�$f�	��P�p�N���F����*�����hgl��Ź�����+}���Ҽ!�~ә]�i�~T�&8'�myJ� ���:����{ibqz'({!�#}W�������TAs�8�+�M�q��'ʑ<�{UvӦ��S���4_L��5�ge���(|m�oa|���x��b��)�LP�{a#��Ǣ�[�riև � ���Vb�t�+_',�#�"|P���Ʈ�����S6���ck�{oe{��F<�W.���0ngE�Դ����$�[G��W�v{�S=�l�8 ����Xt�U��!���s6�YցIճCF�R���kH�_!����-`��=��E�bbꧦ�P�1�3��R&9'E��b1���&�j�gl.\��.&k����2�"+X8�:]��E��\5�'9��_�+�Z.ܺ�;.5���\����Y2۝ ;�9�k���̞�0��N����9����i&���Q�,��"����uS����^7A��s�dF��2�F�	�l>�WJվc�e�"^3�:��8纔�"E���Q�{|3�2V���^:�'��௓ʉ|�� |M^Ƀ�A���a��ukg�k�c.x�U��#�k� �1�P�q���b�ÿ����7��OH�z�Nw�3	��.���IFlG�{V*�����=�u
��V�M��<��,��gf]v��^Vr�P׽�q���¼#�V��R�#�4\iW b<�yAua�K�)�mt����o�t��3�)��<s�0L��=H_�2��ԤXH�ͻ�����5׫s�^�Z��ȃ�=��-�0=-���m�}m=�0�yo�L�	;pZ�kޔ�Y<�^�r�:j�;��{�[����ݙ�cdc�n�>Ø�K7s�t��q`��Z5��ʫ����sT&σ�&p������]�v��v��+�~�����6V�cb�EU�'e�d;����u�`8
5�'��*�
AHá'r/xd�of��
VfB�˲��c����R]���W��<�ـWa��Fwǽ�}x֯Qq�,{ex�9��M����L0���"6�x�F[�<9W��w�O�"�Oewy�g�Zq2H}P(�xD-;δ<�[�� ����yV���� ���Z������7B֖=͵�V�� w�1q�ˀP��~U���Ֆx�W��Y�i�n^��SI�{�>�\�Js�~f}��B'�l�N�^�A箫"vm��jy�f.pnEU��!=�Kϙ�����:c��Mӣ�����O����xZ��u{�}�r~�맳��}(CO��g�*�880Ce�GQ��C����h8��ܳQ�a��y��m�ah�H=�)^W��2x��0<��|@��$%瘴��Z3$�4µ�������=T5}�k�q��p�'��E��^��z��w��y�@/zd�;�~��yk��<��շ��9S�	��m��c�QX�r�d4/(�����1U⮿-&�K��>�ܨ͈wz��u��wǶmn��{��s��)���Vn�q�J�� �nn)6�Ji�:��T
�r������u3AY���Cf)p��'L�I(�>�>�#�{]f���t��|A5?��T-X�����K����H�*���W���� ���j��qn�������(%�x�~a!�{(�Ux!W��q;1��"�M頄+9�c��ŻEt���c���_��v�w���{,��C��@s?���4xO�R�U���o�F�>vf�d ���9��t�uˮ7���ۡ��E��/�{���u\ļ����h��\�b,E�l�L�ץPP��'pً���ϥm�J�LH�I�%��f�v�v�e��荮�=T3β|�)��x�����Ƥ��ƈC95p�F�}��3�}���xK�z��
 a�b ��8��Atw*�4�|e>��pR,`���Gc��*�EV���(��Z�l�z�;�c弬Vxe��WQy��* i��P��u�E�]-c��@S~S��^��8�1`��O���(�S�|��e�����b
T���������+��kf�����T!���癅�1�	M����U�Ą*8���0���dSmqK/��#n���HS�ފ�b��R�o:r�1u���ME)nhڒ&m�G�X�9Hd��� j{×q��u�"���nP���nh��:�f�����Ќ����>�K�������|���1�ۑ]�ܝ��p�\�Z�jp�ެ?�����ܓ�Ӈ
읳[��	��P�#�C�P���u��!
�`ڪ�S���t=�`�����N]�~��[X�}[���w�f~IuH���ɓ&�xh?P��q�fvo�٘���o�q�Z�z�\)�%�l���9k��볻�3R��ȚN\	�ц�U�ͅx�S�\Ц� P�0GT
�{0-�	G�$(1ó_��O�P׺��͵��W / #��'zS�+}y����_k�n�t���X�`���o�����.��P����e�ӧ�y��K�~��v��{f	,W�uA��~Ø2st���:d��`sx	Sd� _.�1UT0/��r����ǵ�jp@+@/����RTS_ri7�烩^mO=oL������d�f��¼6ϡ��U�J������ۚ�-��V���ƽDؔM���]�����o�U@��"Ytm�l����uY3����̱�~�� Q�{�2����ᮨ+��-z#k���rb����W����}�z�W�:��io��1�%FSTN���Ӹ�0aM�m
1�0��}��WfS�pi�X�It�i�s-���v:��(-��M��j�R��F���t+XP�&�,�� �FbgW@���:)�Ov���e����NII��jm1��n��v�5X9-�-Y�S�S��8�;����^�����ݱ�{�����xu���WV���^f��4_��xxR��ey������i㗮��)�+���3�_h�g&���#a�
z~](�o��8.�"���E}-���X��հ�t��-ǈ[�u+�2�+Tb��U�.����w~Y���Q��sd�W^�s�=[J��&p3�yR�(<��QjU��U��s0��#4(X ����o��ÇCMC^ы�p��.�eb'i�ʚwԪv`v���H���(�6/]Cw+�w$�k���F��d�0��yZ�}8��ޚ�����f�,&�!j ;��1��0�wN�v=�s�q�RR��!��ʸ*�b���U�\fV�X��F���V����]i#:�]����|�tU9h`,�����ͤSg��J÷����&�2.��9�9���ѱX�\'-�Z��r���mfs])��8��#w�д7rr(.���V�^.��U����,6�+��,N�W�S�������
��������<��a��;�0���umǋ�4�ќ-iޝ�M��f�+m*��hX�WVW>����Jo@7�6����e����������Xmч�X���x�K��R�M.-_rC2��c�Mwfq�2LU�X�[�r�ﶩikriɵ؆N]MU���yw�O;f_uG�����E�Vޗ��m]YMѠ_=��u�y���Y1�:��Η}r�����
��(DgJ�u�U���^�C�s�wu�e��uɀ� p���w��}�Q�+6Z�n� NT�,�p�{��b��.�v4´`U��ɋJ K���@y�(��{f$t>�����fm1��;�q�[7���|vf�fk�gE'A�>��4�����g#�dP�7���Ėpx�r*��@��7��;�q1���H�͝\:�ֶȸ���S����հ[����V�=7XPm5�tv�{^Rݵo	p�:��P���M�+�o#A�S[
T+h���Ɲ�7�p�:�틃4�,�+ ��l�kǍhե����q��:��T�`���{M������g�W!�(:�
޷Z y.��=���x����ٖ`��7����>��ΏPA���� ��;�B�
�M�T��_�� -��G�V dw���O�J�&��u�-im���.����Cz(�ײa���V���7�)f���V����]R��(^��z6i ��tZb�J��U	�e�N�YK���v'�9�ks5p�a���!���e`�`R�9�$�`��� �Eצo;C*�B��S*�<)�Ln9�gf.�\�v��U�g�JQ)�&i��]�H
!��	%͹�`b�d��vM	4��$d	)�"BbH)�H�$�3bH"H�ΔD�BJf�)�CE�Lw)I��f�hM2�,���a#4L�I���F��Ғewt�����`�I�̢3�*�i*A%$&�hD�2%&��FS
N��YH�BA�@s�)&`�]�A��wrTb����I�ȹ�E$�̓0Jd�I!���"nt�
N�.�&I%�����) Rb$X�JG9d��Q�2�@��%���,�:d��n�`�ݸ�	@h˺�%$��bb$A��@
�(|\�W�+��J�R�ӏ��z{���h0F�/�j�N�6�s�[a���.��p����+n��{�Ǹ��������&p��̩�~on6�ݧ �P8�/��\�-��x�tV����I[����EՎ�-�B9�X�p�v���k�V�(/�s���<F�ҧ��Sh�)�鞐\�B�7[~�Dk��G�����03L��-�1�:�6��q 
���51�&<ι&���4��6wOV|&�]���N�9�s�8�*��y�����"xa<�gsz4/a��[��8F�JQ%�c2|k�:L*����.c�19�D���(K�ď������\X��ۤ0�hڰY�$`C��aL�t�]��I���#��x]m�q�7Ƶwv	�%j�]�ή��2���\����i��Vvy"��)���/E�n�P����@�X�?�4GL�X�?`��U{SȌ�WGx��k=����]J�������Lk�r��~�i�f�;M����x�^T�,^�B���[B�g�'X2��7���יO�g�-�~�'��m��#a�5�{l`!�I���b{�ʹ�;Pf�!�	 3��-V�_\�{�پؑ�"��s!ø"�kÛ�g�	��W��6k���^6w� <�����y@:�Y3�<g�:����+LCO�ИznWH�s�F<z�:ew;����<4b�tT8;m	���sk7M�P����9 �t&�z����e��_W���Wr��D�o C�x�Ɲ���l�V��G�ڊ� r>�SuLGdk��v�(�&M��i��u$4jǾ��p��\-���4�6'ϐ���?b�WK�f�M��袧8UaV��N��
b��w�i��r����n��P8x]?&)��8�L{ea�@n��+&ޙ�Ƨ��
VH2���9H�E:��A��1P�۞9f ����?�B4��>@WP�{~��va����ҰƴZ����0���M�*��F��OT�|a)R1���/�w��Z�窰��p6s�!�J��If6����2������Ͻ>¬�� �IL��1k����ZpU��,w�����7S�%(��+yW�i�j"����^�q�>^�v@!�+�*��z��2e�ӫ�:�d��@���xE�Zg��ZKvٌ�oJӐ�ƈ�U!�noj�H�/ޒx�>���D
���&#�2������G'h!�����u=L�.R՛��/�E�5;�)�;���'�t�;��B�py;(xy��m��v��x>���\�B�S�}��u9һ�t��o��˫���Yt}}�Y"�nղ�V���!
��uќj�������HKW�ɋ�i͕$ѳ�A����a� �շ��0m���z�˫�ޛk7���9�r6�w%sY����$�WY�q���}�������a��g*NR�C���!�\K`�1��`$鏩MӢ`�=���|dfu�^Β�@)&Z�����ĕ]�<"�nX^46ำ�Ò� ��֞v��b�yޏ/��V�A�L�,��x+e}��	W���e U�����5,�Q�Z���EM� BJc'��[��`�1<6�(�i̯AG�ޭ��w׽u�=���[}r-u:5�]t��X��Յ��	�tk�՛5~?:\���k�Us�u�����e��^tW�ts:v������f��ǘ��AY�� ̿��#8�6gR��(�Z�ks6��t376�Q�=���B��u�'��6$��o��xuU�@s����u4�-!s4M4������n�ܟP0��> D�@�<��9B5ˮ7>k��kN�� J��"�/6ܽ�;�g>�@6\���&1��C���X�
@�(BgzW�jR�?=oF�ܱ��И�vӎ�vߺQ��&���:�i��a	Fk�Nޖ�f�X���\!�(�%��W��zP�t��)ֻ�1`p��,8�Q�ew��ns���u��u�u���t�����]%p��s$���:�x�dq
�����rd�\/i��N�{w���M�z���o�A3k�Z�xi�:M�!���tJ�=�fɲ�ge�ﾪ���Sǘ��� �����Z$��L�Jcjf9��)*����K�����"�Y�h�u�A�4q��G�\��cr������*� �-��t
S|� ��1}��3ng����
 �ϼ=<�e��]��cwM��?Rs��D@j���Os�U��w[�*z�Jݭ��E{]�RMZ��0�f0a)��Ӹ��!�����.�w�ф{�ӓ$s1z.4�z=Z$����>1��3���k��x``����0���Uc��}�ka@�����iYha*ˈ;?����k��2�����}��]˼J=� 5���@��nT�>���������s�tb�L`�.[g��P<��a�q�gw�f��}��5��[d���M�����%�O��gy@����U���׬�t�_�`�2�1޽���s#�b��A�Yw�@O&�n�p�<��Oe���}*��r��Z��ޅ���,/6z-cA��0Hi�F�
8�U��U=�t ^Y��Gm*�قD2����
����GE�����B�ǹ�/��F�&I\zO*�=],�~�.׭�C9U�+*�t�[��ޘ,\���8 ���90�d��q�27�w]��c�f���M�n%��-��פmۧ���T���8���ξ��-��u���_ff8��Q��U}UUY�������܄=%a=q0��u�����eo�/��{.�����ע�N���Ij;H����{����v}Ek�G��3���\�%'��\��T�1�ٌ�^���14mΆh}y��6@�:=-4��K�SKکqFY�Y�9ˣ�ܶUNٸ�S��hz��-|�N(�߭�P�R(Ag��H=Pe��dW_%�D�׷��LWJ�>~U�{o�kb�]o�����Z1�`q�m\>ª��0خ��'�X�}��iWN���`���D˾Y��{}��j�!�^H`�F��#��c�:��(��w`�uyC�n��Ҍ5j�30�������v|ұZ#޹J.�Z5�7��`o�0S�M'U.n 7ag3n+��G��vrp�a�k*�ʬ�b�I.pBG>s���&쎷ub%�*V�hZ|�o7�����Nl�Xl�������_a�ar�h��8C�ɏ):T&@2����Τ�����,Mm��H�mb`�+�C]XS5�R&6u�A^Yb�5�{�Jo��{�t�
�,�͸�V��gG��cuX�yp��}�����׮`��z|�m_˙֨NX�[X�8�ks��]^��LV�tNڋJ���P;�ø3��g���	u
W)���v'Y�X2������ӡ����]�r���DDEe-m�S@�Q����c�*�u�b�ߙ���1��X��^�e�I�1ie��y�/�QWS����p!L�X�S�
�qu�ё����Ƈ۞Ć�g��[።gU��K�Jj��qp��o8*U_y�>�9b��b�o���<�:�=�mt��ۥ;x���]
z{���Z9������tc�b{?{�E��TH�'5�Rہjʽ��j���x���6�r���3��Ua����Z{��|3���oµ���)�d>Ż��<{]�Վ=�>>�T#��>�0e�>�S��D�%�{J��:]s0 �<.�. I�H�Hl6�L��H㩱�	��g��b;�B��gJ�9��ld�|�=o,�
n�W�uU����Yø?o��Xf3�Sknx�8|��҆�L�!��=\�����}ݔ��RX?y!�l%V:5D�q��}���zo�W\��� hϩX|�L=װM�g����</,��au2�#�fBQ�Sß>��n<��"�޸�<��?1�Fr�si?�0lV�ѳM�z��6����q�6�ܭƯrWpbh�i��a9;~~�cw�<�y���Z���"M;��]�B�վ�f��/:�$�X�us���M`���}�,��gN�e�+)�Y�ϓ3/"��d�[�@j�oӸsV��ho�U}�UUB�����;@]�9�$��(}?9�f�ʉS(v�S���]ҕ�㖷��1������J���,S�h�>i�w:+|tV]sTg�ߖ{����0�mӴ3���2%��2����kEv�~�''��\g�D
�� b}��O�x\��;��ʍ*�{��2 �+��F!����g h��7EG�i�U��to�HJ� 4��ϙ�4��*�]����;w�OE��ɫ����~��q/"���w��ιG�eiD�L;#~T���e��>���OG�S��+�I>G���TW�x0Ce���@SCC�03�C���s:}+��o=�_?��nPt�x�~c�#�)L7\jO�}��W|@��$#��Po�k���.M�W�򫺗���Y�����X9��bxo�~.ez
?.�l�9��H�f���c�I踅��:Co�XP��տ�xj���\EN3�D��r��@N[��C�7;uٵ�M��Q����&8=��o��^��ja�*��*#2QU�����P���F�J��<��~�:t�q;���';2@�&;�����X\���`n��öc۱SꊚT�䩘�Et��i*"�0t��O+��!t��Wk9]�]B�U��B�p�v��.WM�\��h��	[��"j��.���CrQ�]O&�+[6�P
g�着��������77 rU��+���Ϊ5ϛ����sעg�c�t �{!_@��Z�v����kcZ[oV�u������H ӝ���t}���=�յ����nܟ��<aE��ӷ���iZ.�����P9ɖ:�4���N�-St�&���������>i\hש��N�c���T��1��%��������\0���K�����{�s�1V�)�lb����' T5h,w*�ҭ�O��Gq����&�����W��8*蓕�\'#J����RuC��,΢�+@Tp[�N�c�b���d�'�.���aI<��-}y~��x�q۞��э�6*��I�i������r�{�s��n�
��}_b�!��MZ^W3�&�u�J�s��M�oKVA`�N��� �m����������m9)��Z��\@B�N��b7Q&����F���E�l,{��I�>τ{�Ϛ��fa�/7��������%��=�+��W=[V����r۠kZ>��J��W��A�k���+YS�ӥ�{�gW�fy�]�oh�Y������e���E}��ӕ�k,܀Ów�ѣI�*��0�Օ�D1��mm�+37�zA����~L���R�{y{1=��{%�hN���6a�6�ہ��S���ꪪ��÷�z��9��_0_85�
un͎�g{U���s�F�wx����s��3�.d����nv��wC'��,���DkWe��k�l?�+��J���w2�ԣ���uD]
t����` �j�,��Jxg�����վ@�t-}���5�״�Z5����N�h���CX��(p����p�Q�R��\G9���=����������-��o��z03ի�A�̯Q��?vd���{��^�5y,l���K�Y��Χ�s2��܃��zp�}j7�����/⟽x���O�����;�M�a���e]X�.��C�od���*&/�nM�W�����-Ϥ̍�q-.�/9���p%��*���Q2�J)uNL�ݥ��I�!{"���e����qFq��}�t���N8;��/�������>��
��]drV�n8Y��br�|7
��)��l �N!�,�>�ULc�<E��h�}��8����R�:򮤟'ܖ;(nԙ��o&�x����zk<v/
�a�	e]!ٗԝۚ��R�ώ�Brڲ�����7�+v��i*#��͡L^��W�g}��.��S�Y�t�4n_5͵�������}���|�T�D��{ᯈog��.�
�jqyM�S=<�Hwn�T�c��M,}�o�~�����жo�U�M+��R�g0T&�����@������`T����u�v������=r��M�ιsW�5n+%�Ck��9�xK��kGz�]-���/'ZGk��5G����Q��w8/i͉f��m��W-=a�̸�pD��TLs�<��mI[�r�Mk��|���-m���(��p�g\CJ������k�
r���:�-t.w	��v;võ�W��^��S-�fkp�t�=�w�ë�{�{�=Hn�U����c�;�tȞM>��ڛ�"�^}���V����w�Y���ǲ�j3�������52��v�/�f#g2y��Pn���:g�YOWH�M�$�����^�]:���>��{N7�;l���V�W��_Q��U)��z�:��!I�~夆���t�B~}W�}��@X[1ǝg5��Oؾ�w([�a����h�2���C����[���DA))��X�;m����y%�V����"Qs%Mnt��z��@Ea鋍�����e��hS��+��a��_2+�a�5e���Œ����:��eqT��)H�[+^8jwYڛ�LR�A\ٳqX�i�3-�\���5�K4�nC;-�6��qKZ���ՙȵA�h�Jݽ��"C��6��s�,ŵ�5��^��#7�5�d�3�m��%�Yt;n�c���� V�A��&�!g^+�=j� Z��5�u�`��Yk4�*Gcp6}N�w0��(h�Wˉ����ڍY0�l��Z��#k(�͂�>�ZY6��4	K$����4�[{�b�I:)ŭ�2�z!����$�I�Գ���m�M��ƺu�\���ۮe��Qm,w��nf�о�#�z��"R�D��h��'�dQ��k�KՇ��KK�[�^�#{jr��;�qb�[���e��V��3@w�wlO��gPp;��2�L{D�oS}�Xw�6�x���U.�f�w�u�D��pI}���-�f�\��Q�Tg��z��%�=�tj�9��*��$�kv�r�x������R�(J�n�[x��p� 3"��й6��vws��4Sk��ֺ�����jG@˘�t�Y��\6����q�(![[�*s�"�h��>�p�=���x{��R$]E`p�|�٩]Yim��/F�0x�q%�}Y��q]VZW����wΦ�3�Fʫ�X���:�,0��e�E[��>����ˋ��c�#8��w�'1����\N�i���ՙ+B��,L�n�*`�(3�s�,V;_L�l3QN��We���5/�0�WҞu2n���C�󭔷�	Tp˫��N��:�����Ҟ|����&�º�L�Cc|�<����x]��<tṬ}��
����gz�L�d��+Uы�fLW��>XQ�Hϧ*\�d�/5*Jڮ��+��ؙ�%��dY���9H2�eno�Sz�f4���uh�O^K[dV�}I�v9��ÌBm��7��P��*��Lژ����{έ��ҏ{�03���
� U�(�$J ,N�])�&��M��+t�Ե�������rZU}ˢ��^V6���
���|$6�$���sfd�sS��2�!�uk�IR�v�y}�6Kt�J�XfoW�;��s)MrԎ恎]��:Zys�WYQjJ�4�%���OL[7b��J�z��}R����Iϰ_'�V�*������������ve�p�΋��R��Suxtӈ��2K�����P �Ch%nI�KW��d�(���Ƿ��w�˰��c�6��Wmj��$3u�����w�nJ�Ĳ��GT���K�9;����J�R���D��\"mj��ـ��2�*��mf�Ը$��}�/��O�������w����1���	M:9�
$ecf�$\�DFJ$P�	�v31�2
0Rl��L�0I��$$Ph��(����P�!����HRc&&J)�(%�iD&ȘJE!��F�	1� �hF*#E̍��i# L@2� B$�$�l$͍�!#�I3!bM��LJHbL��0�0���4�F�1AA�L�@hДĆ�H	 &�	����M�M3e(�	
2�X�4JXBM"4��	RQLč0�L�JXdL�JQ�(��CI{߿߷��H������j�ڇ�WRl汖�&.j��B�qPYi`�:�:�C5�f�.5t�5ev��fC���W�}��U�h��{s���u��gwE�-��E���G�����K���x���wJ� ������������6��������s���e����R�M����wr\��=���Nn�/��)]���|�<�8�5m��w/s����n�-���\���W�S����)F�yp�5�����Q���ˬ��$�v8n�ۄv�"���v�U'�����K��9{����07eĖ��hI�O��.y^r�᝘UB'����/����L�y7��}��疶r%��f�� Ffz���͇T�L�]��~�J�{w
�&�J��p;{�C.NQ������!�����9�S.k�!u��Z�eQr���hPN,Mѝ�\��W6r%�={��\�M�vˌp�1:b�Snk�}r��,:t�ZI�}dܸ=�5�N��w���J��s����̉�7Vu���]�7:c-��d��[D-��6/_k��[:s҃E�3J:���j�0)kk�BHQ�.�>��W;	���,'3�.��`Or�O��[ׅ4��P=��:.�	�A�ک>�mk`�vC�����7��%��ꯪ��,}M6��I9=�.�}_OfTK�5�,ΚYκ��ᚇ��L�3�M�g0�' �
\%ip��b/,�|�e��ή�
�;y�	Ͻ�q����{�2��{U�+	�괴zR\���VR�;'e��qv199\4Z�\+�ϗO����X���4<iNXq6r�~������֬hs{�p��W8�-�U�)�K��v���:�Fl��{�̨��q;.�\>�Q�\F���)��Y蟹t�{�B��Wf��F�ο�3y ⨒��G,�(﯐No����Z{S�ٌNgWk�	S��e�{���*�=�/�Ҕq7oC�9©d:w'�sNx�j.d���ա�q�R��8e?��T=������e50�o)u�qW"����vk��|19o��t��0v�~���a�֩-u�	qѓ����'�"z��5&n.�+��x�䙕~�ޗ�)Mҭ	@����W�3˝u���W~a�x�ڙ�~�)6�.��rmq8�6���=�kX5��[}�X�/-p���#�� qx3�a�#,wũ/ayĪ`����}U�}�|'=+Q����h��O��=�m�ߝR��NK�_5?�XD�|lg)�<��]�ՙ�W����|��;g{����yW�W����پ͡�|u�0�&�ONE�{��.����s2k��c���S|���
�ͮ�Tf���|��G��NX�4}�N��Ӿ�y����sI&	�x*R�gE��1K;�)g�r%8��%8��v�>�sWf\Jy5�&#:�Fr��8�<�-i��Y/��A��z�����ez&��:K�y-���fSW�kT��b���Ed���_�[�\9��R���k���끑o�ᘐ
�}��1��+�KD���k�Y��|���39�w������Ⱦ�X������3�KC���t��G{�q.5�3�Ϋ�'���������40��9�y�~��w���h��#��P'>����b���(�*'y��
m�DE������<wN��O�]���.b�/d��s��nùtyo�ٿr�u��1�&<��ڴI�>����q�>�k]�\M����(,]�p%�봘
�k�hv��D�V��蕼�7��4� 'H΍>A�Zr;ѽܲ��kFi�;10NLq��]��������gv�dn�����{�C����,>���:�5�����2'.�+�s����2�����OBVu|�������_I�%������6�Ӝo��Sy:��[��e���i�|�4�U�.�����Y�	T�{�znCE�}U�!�Bomt����������V���W�9���͗n.�N~��b�^��*�����x�C�CU|}7���3�eJS�sM(��!�B��F�s ���)��z��zes��Wý!�:�3�/=�QVW����N� �B�SU3l��>u=0r�~1���ݏ;�ޔ.�Ți��j͉�����"b�5
e�}Bꁵ%k���12���[�6W5�%
l����SM��2���0�TO��� �`mI[�Y�Rއ��V�6�R.�Z̘�Չ%3֜#M��fz�n����7���:n)Z_�b��um��j�!nD@w�e�Nu�W��vF��Ct*���T�i��(��!u0[cNQ�ZV�����b7��;�׎�]̀�˄��J�c���VVH���nW$�Yn0���*�<.s��XE���o�8I�I���ﾯ���~�v_��q��A�N�,�t��]x�3_<�;p��s�5�C���<�,�O��ݝ�
��^��i0|Ug��S��]j��{i8�x��w'en�d��2���!..�	m�M�0>���M��%�Q����RަI{����ھ��\��l���͟U/%���;l��9VU*b��zw��AҦ8���H?��Q9m�D��o;�1������PU�:�%�v�x��KD����4�L��9�0����79M����낳�Zz����b���Q�M�m懢\Nrm��*9W�{�0�w����_Γ�*�\N�ʊ�a�{E���eMց��n�O:�K�(���<�����p���-�EDɠ�>#�C�\o�:� �Y�>}r\��D�N�,4R�X�u���[s/,�MY],��E��#��6�SW�x]B���5��wپՔ;&�=���+ZH�Y�1���t�N:-��졡������*�/�|q5��o;��jЅ��\���K*Ĵp�W����$Wb����^�t\��;g-#��s��Yd���z�Nёl���\�ĥ.�*s�	�9�;���G�G�*^���ރFR�q>�ڞ`�ƹ�9)���]0#O�9�ԭy�YiB���U,�c��ua���	hM�B�{˜S.k�]B4����²�R���.55���/s� �����2�+���r�vtV�&�t�<�#>�;���sp6�s�f�YI��J��s���)ˤ��jk��c����kohQ{1��M�gۑ!���rRig����s�������s�s�.�jr��qf���t���3D�°^g9˫P���"t�o�f�m��YnQ;�{�S�sWU���Z]��=�V�b�n2j���ʞR_�W�ܙ�ٜ��������W�Z��#]�#Ɣ�[;s=wٻ:��{՜�m.�gKٞ���g�E�)�K�����o3v�Q�
�\~�QOO �f/U��Ǐ~ή�I�N˛���כj!uv�)���AT<f�q�V�ï[==�"	��v�N�ӎ��c�Yۘ�Sk����p�D.�ok�]Mpɇ}�z�/nU�{�*�V��l�����{,n&T��)&#,+c�/��1�^�Y��jpل�K��:M�o_+@��A��1��>�>��E���v+fw��9���u��"Tr�/�(ȾA9�M�jDi�u�;˧�e�����^�R1��`t>�D�ꉗ���R�bogbއZv�JwF�RVQ#r�&;i���n6�ߡp
N���!��{�L\���7��cO�4�T�R/����Q�3���:n�nP��?�(�*��2�ݜ�+=�vn���|�����ۉlc�J�����惢O�Y�O^���~9h������c��*��҇ZچsBok�=���&������ � �閞����V��u�{{\��|�l7@��隆[g�=Y�v)vK�L37�/Ҟ�ٹ�ir��;{���T�`&�y�+��25�JJ�'0�1?�<��qQΜ�O��gD�x�\���~ݕ�ҭqxj���sdeV8��M}m�)�9�NTk���UW���K���+���u�O[�R���~S��������.
+��B�i�ɶ�|�.nS���ds���<���5�ԅ��]]]5�s�6��9s��7��^sX2�{f>}��]���Q�:�x��h��fZj˚y
x����g{�Hb�ّ6D���S��U_}[����Iʛ����]_\oJ�Z��C��~�N����Vk|��S�L����A�	Ĝ�u}+V71�Z��V���;�g�+�ox�Y�7���m\}�����!,�z�E��J+k����o�%��T;Ϣ�������L+Rşm4��Vhy������`ꈗ9Q*V(��՛��!-�f���^q)��ڊCwg�x�{ϵ{�Lۑ�9���X=7:�o�=�u�.E��T��)r�}�P�ւ�M�/���M�.����+�܍���(˾��O���t���J���w��ᬸ�SO8��zp*��)��d���ݗ3+�r��6佩/��+{�h5����	�wp�5_wL�+Z՝/����!�H\�$���+���u�V�S���3�
�����Wljg����Yꝁ��{1}�>������G��^y�����Qw!�Z0�D��'>�I���:rh�Q7�2t�蹸�����zjf����B�0���t�Yh�p�|^������M�8{��ʲ����(3h�ܨ�qӵ�1�d v۴�9B�k8uIp.Y���g�z�`z��ó�d6��������N^A�%�����o��i�B�����=s��Sp��9�k�z�}[=��1�\�6)㜩je�q�N�s��1���{G�U�O��%�w������;�\c�!8��N{�}CkTg .�yw{�ٝ�o}�,�^Jq���ߏ8E��Z��y�=8fffP�-=��ޘs����Y��_,�<~s�
�W�ז�3^�0|��u-�����<��wE �U�Y�ڴ��a���=�#��L��	8�nsO��d�[	R�P�Ώ��>�雴���hڃ�m_Eo�9[�%���ZewOF���w��*�H�����v١�Jr�8�W��f<��U͌�Ackܘi<W(����ſyI��<��ܛ��a�/ƺ����׻�.�GQ��5���3����}q/�\����\.QT��UTm�%ͷ�g�o��|��ze#�ٹ��ʊ%Efү}���U)���h�����7@{h��L�.8�5��@�v$��i�����ú��/9:�׍�|+^;��d�t��Dw��Ont�[�9�t�ڷ�����SΒљ��8�-����rO{�si�g�Vڕ�v9}��6���{pU�ռ��1v�f,\�R��)��
`����Q%�R�DbO.�,��N����sљ�/uj��f�x�XW��wӲ��C�O��Ry9JΔ�&�Ȟt6V�bz�T	��Qx����|꒸���-�	E@�}7h����gc�`�>z.g)P[��z����5̹�2W|��gn;Z�-}�8	U�����/c�J��3hT&�*ӚS.k�!to���dׁͭ���.%<��k;�؄��&�;�\c�"a:a�s����qztSt ���ګ{�9����䟏l$�ms��!���t��6%�ө�v�վ�J�=9t�?k�d�[v�]~O�����=��3�r�;��[ރݦ�,ʐ24���;Q�WѮ.�!�?@լ]��z���Ż�z��ǐ_�8��{ix]:2zt�H�0.\�e�j��:��ema�DΡ�{��j{r�9Mv|�������:L�����Ќ"S4P�{e�Gn�I����۩ҫ�r�T��M��4�h�j���:J[���llܖ�G�e�҄�Ӛ$i�b�T��S�Wz4ꨬLd�Pvk�-�&N�ﭪN����wi�Cϋ
���BD�W�*,[GZ�o6s}[�G�\_Y�R�?�xgy���}Eހ�;�Q�C���ᨦ����;<����{�f��>42�� �v`��� �:�o���X��U}�s�rk�� tv�^�2t� ��`�+v]gM$W!�5����4�u�\�jOWL��VD�g^�+�r��yZ�X�J�wu��T�-����_�t#��M*ꋇ7�ayw�v=h�Pv��{��n�{�M$�
gva��F�c���0�''q�o-�J�a�MK}X��հk���W"�0�F���,Es�qg6�؆��=�h�ZY�m��A>��8�̓�b��C����+{�>�Z&�# :����Zd)����*C�^Ԧ�mc/�k|o�4�����ck]F�9�T-�=PP4��3�c�֞�Wz@}O�(��ݗ�Vը��2C�m�I����7�]]e<O�K�{�o_Ɩ�u�I�J���j�fqY�5 �Z���Q��9{ݴ녈�Yu���@&2b��v�CS�N������|.��-�um[��m���]pR�٩4�� q\l����ܭ�c3������P�!���}���.��7:���3z0p|y���*�+��que��<��1��s7�q� $/6Nx�h��/Ws�m��z��V�r���&�8��6h<Ƴ ΁�cwU>l�1�F�`��^�:��b���k���Ѩf�	����`�V�	��6��=��1ಭ�7��!͎׻͂�]�%�WzWJ�*��yZ�cu����{@ޙ>&������&Z�6o;:V���v��켶��f$!(��a��4[�拊�G5�`�f�����k�n��g"+;Q�Dkw�Ї91�7���ᛦ�m��ᏺs�3M�G}�Y�Y8WlaI�j��۳i��Io-���RoH[�`�8�IEK"��δ�u�I�犒�oV��w�����V*��r�Q�E!=�W:�^N�S�(B�MV�r�A<�Ewܫ^��m����N� ���q�t�]�OZ��k�jΡ�H@w3�أ�P�HN��D��`���C*�S�2H���8;���A���݋	�fghL��I��{�!�`
�oOwm���i��)W�
�^�Yz�����uې\Y-q��t��}�X��\|�I�qʹ��?�MEu�0ko� ��)�#�Y��l�t	M�����l��sUs�G��{XIO{�����Gٳ�`˗1lѹ-9:��/�x��N�"��2� �ξN�;t/�O��?�O�����@��E�14E&�DѣId&b�$
QBd%L1!(�)D�4@X4F	$1�1���a"0j)0fhH��S&CE"&`�3hƓ4d3"�̋D1$��"H3@�0A!D�Dl���0��A�BE"�&X,cDL��Ɔh�����M"TJF!�*RHD(1%JH�24ԈhL�$Ț1���M�a���R(�J,�Fhفc�b"Re�d��X�$Ib$�c4hQZF$�(�
`�
� ����+�C7*�����s����5��mU�'X}R���D�Js�y��|��e�ص�N[ޚ- ����������r^����&Dn*��׍�7���c���&�5�̨/� fv�5��|��\3:z�]�@�}�yУ�ᙜ���Ó�ޑj�X�y���ʂ�]����03�S>������R�:\�����}^�yC豜W�i�{r��׻����	�Z������V�¢w�3r�۔�f)��F9����e�W���G�j��P9Ωk][��>��aQ7�'#����eZ��{N�|�	�������]�[.�B�Ӆȳ+�(ƈ�r2(�v�1b����u|�e�ж�M=����T.I߻���Z�')0�v�9�)PPz��SXk�F����)�}-o{}�mmwӰ?�I���l6MK���h{��6��k��K��+}�	le|����f�4�^e���lwZn����:�����v/��M$�x�`�M�v;�ն�@]y�Y{]�Y�ݡ��r�Q�O0�c�(L�\�7��f�T��(�&6��v/.�hE��D:��X�sk�?7�=�w���u�4э�U����:�+P�5�)-����ti�Nnl �]I�d\�nvDB�p��rzWW.����[��OI��T��e}�}�騕���Ҷ9s�M�l.yU���kj�r���Q��pu�y:�;]j�g���_Z���_q�eNt;���r.�\7��7� ,�~���>ɞ����!�8��4q�C�G���WcN*�.�u{o�MZp�Bn�S��>}d�J��'[�y�HK!5��ՠ�}X�f�X��8<�?W�j������X��KRg�]�f�	�2=�/9�@@�mM�>�Y���?������w��?g�4�׽a�o��HɋV����e���Ù(�!w�����k��57��Jg��:�����)���.�5T�6���g;l�rÛ�ŵ�^���RZ���I�ٱ1&4�R�A���)%�.�5�>^�V��G���ut�R���cc���.7q�bnru��b/PN[oTD�}qg6�����/�r��!7%���]b)��3\a9Ǎb��kP��X�̭{w*a$��s+���Y휉Hu*��O[�:��0��I�*�,��q{:�>����u9��v+�qM��\�o���-��]���iq@�e�(�T��S�!(��<���eE�>�����"���1zg�Z�-�8j�8[_&��\�NK�C��E�(ޖ���3�p�,!<��ʠ;�\e�쥢�t�I��β7s�(�d�oٳw梾*��n+��)wB�؜�Ĥ7��H�r���{�n���;����U�|����>1�4;��^[z,��1Ӝ��*�oy��ci�9�2Ut��4���Q+^_�/��*lQ�p��x�rr���;��l�
�ȟ�:�u�y?���Agg����}��o�ᾉR2�_gNwIuO$�_2�+���yۚ�[�#9�-���U��]dܸ=��]��<�v�U5�#M��8�[\�[�}���^8���7 �+"�����K~�/2�g���N{a]������'M�s����t% �/�TF�0-k|���]b�^�}q�MKؖ�@��ѿ"٥m\M�@cש�L*�qň�y^b��ke9���[�.�8�T�Ҋ��);�AR�%�x�[.���8VwW9���Y��̷�ma� v R.f��	O��	��w{g�;�:��k�z�mI�������;KooVdfV��j��Mܪ�2/}	���=s��9w�etf#F�'�2�cSU�E�;N�'���2�73�/�-���/H�����v١㖧�4s2u��Ղf'�=����Qҹ��d�ݸoz�1�����U�hM�����OW���S��R��Dd��*&�ss�So�%�낳����9�6��:�U��m�jjP*���\r���X]T_G7x��t��Y*�ӗ�vG;�g����������}%�(�$���ky�(B��<&�,��u%�����>�y���
���#����T,]��H���QW"���ƻ>��ʇT��_/��	D���qn�_:B��=)�)���ϵYM+�n7�*߆y/+�H���
ɰI�蝳y�ʳ!�bMn3��.��*�94�7���ew�����>K�W�� �E��L�Ɍ�"�á��@�e�������O:�m�ON�M����~5��D/i/q�]�g\Y�+�-�O�RE�Y����]�y�ݖ��7�+xu���$z7��gEVީ�o+o�SC1�w�npx0o)l���e�� �K�7WH줆.��?ޒ�������=	���Ȱ���i,�}	��rrn(��X����]�N��U篻�-�����E[��O�9g�r%0���tډ}�6�OfTJ�5�s���ҾE���"�.�(ee�mB/ߓ��q{��w2��JK�y-��k��x�\�r�������N���Χƫ�vC��{]�j�@̢��ja��.���bulZj�\!��P�;���g�������-�y,]�ҹ�������n^�/,�}�Ëj�u��TgKߦzz�ݞ}���9����!��/u�[��j ,��U�A5n�uzm/Tϐ�Ϝ��j��ޜ�)���ĹP���i��X��_ՠj���9�>�K�z��P�b^˦����z3�L�P27%��]r�Я�i�O@є��#t�od��.�l��|�Q�II���K����Q٠�������~�}%�U���H}���\W��2m$�=�|�#].݊�-�;��{*���e�>zٶ�I�nU�ٛ�
�^,0�Bx{�	��S��ݧ�@/+��^V��%v����J�Es�T�컻�Ė�����o.�ޅ���SLn�26 w	1p�mK_�CH<"�Ol�6�wy�/t~�����W{}���=���}g��^�`-n{��,5겾S��������F������S�S(�}۔a���^�'��Q��d�}������-؋�+�I|�l]�fvFn�Y3��)z�B�
��_&uj���C���컟��n{������N2�g���\М�Ыa\.��|���ۃ���׶Ӿ�;U�{<�gj��҅q�q�j��`�n5���YF�x�6o��9C�\��·�繞�7]КH˙5��k�L�֜"�����}d�@��H�	�7��m�Փ�]�R��==�H��/�>�t�s=?W�k�{��ǳ�a>����qy���nt��H}�S�I�a���Α��V������<#&��Qo)WM��R��KZ1^��l��+��1@�Np�(ؤ7����`0]�:���B�Gw���˰�N��sܒ��p���p
)<3r�5��o4��T��'\Ӹf��q*�r�� ƛ�Y4�';s�93�Ⱥ)�;\�m�9ov�ZTEp3���5�^�-��x�E���U��Q[[���3}��r[ꏆO�W]t�ތ:s�-���L���iy,s���9a��=�uz5�$��qg�j��=^Yڝ����g�g�}����r:=���$z��z��EM�2�]�1<��*&/�n[oT�}qgWͭ.�����IWr��x��1�%�ٷ��U2�\E)J�Kwxᬼp��OB�]�@.�7���Z�Y���7Z��`cU��U{��{���[�u�]��fͱ�1��7uD��'7��k�s��?�~*���n+�)w\o�w�$����u��=���/�������K_ouQ���P���;&�w���9��v��c)$�nE���;|��	��ꜢJ���4�}5��g���=�7s �t�O�����v͠��d'NQ.r8_M����P���m1�h��.�4L�7�F�ԭ����ߞ9J�X�Tۤ��O��I^o:V;�,����կ˸d�?YE0�g�Z�R�����_a�>k+�N\X��v�vf��Y�#�;)�q^�V*u&�VG#�w������$�s{�\v�ƹ�K{�3�٩�ܗ��X��qit��L;�\c������nb��������Xqj �p:��e�)d�bɌ��IT�Zp�6�]�9f�%��u����ev5�������G۞Hr�t�#���l+�L��g� ��������9�sZ�8�5��;>�V�ma���V���R:���f�C�
�v1�z�0ee�Ѽ��=~��K���eA�Fbț�����Q��H��Mrp�90w��θs<�৪ۗ����^K��v��UZ���<�ۧ��{�Z����Nnb�壣���Ko��O�si{�C���Ӄ�R�Vs����Rg&n'���J�Ւ�������}M�O9C�G=��)��r/9�;N������W@�I}Q��a���9�Ifg��pz�ł�#�<����Nl�~=o�NK��;�Q%"-�(�N��.�ۮ�I��4gIӋ�d���k��,(�ֲ��r0#����-ܤ6�>Վ�;�h�{W׶C����^O�2���=�%�㲷�0F��<V��v��6Jwuhb�m�b��x�hj+��Gm[Ʉ�B�:�z'c[�\��[O�^�G�{��M�i��ܴ��CJ�O'Րl�*�Oa}�V��T�R.K��k�ڇ��K`<.���)�`%r-�-g6�6ډ}Vvn��{1|��Ұ�V��;�lmC�r�+�Zm]��&�UŬK^-t�d��6YM+��o���҆�5�6�Bob�ӞA�#R禷[����Q�`<�Ai��L\}���K���{;ށ�\cQ�n��B��0�����5W k՞|0�W������Mw�_K�x�%R,1Hm�\�L����@����p�F���v�X��m��eJƝ��2����2��{��ȶ�{VN���.����_���uV�R\�<��^fͼ��p� ���L�0����w�}=��o���'~�'���y���o�jr�o6��B�'���eb�OU���k�������%�p�Ue����e�5״E�dX�yr���}�l�Z�����֎X�u���>������B����SFpڙٳoN��*���i��D�|t�e�i��|��s {ʢ���#u�ٝ���n��@rR�%[ڟJ��F��tg
�9�����qSV�v�J=�ߨ^sQ[�����p��_8�)����ޗ2#�L�7@��E�˫����|�|	�mg���P��t�Q1���Q=��ĸn��YU;�e����Wy��s�ke��3��$����>ӕ�ʲ-�z��p��;K�Ǟ���j���G)��1�.��:0*�Oq=� 
ZH��/�w�2��U�✣�����zt&��m�@�*�h�U�f�������y������RXj
O/汮ϵ�u[�	�j���xa<}:s��Zi������C�afV�j
]�[�ϓ�m��g*�F����rx
�n\r���_f�J$j�6�_i\�J�m�X�*���۩sE�%������G]j��Y]�S�]�Wyьu�މ6��y�9�,��G�;�w\Jt�4�[�6���}k�.=�`��-��sN%ҾU�H��}B�[�"��*��xoP���Z2��q�J��n�c�������7e�������s
dPw3��²)��]�h[�]rr��.*���\�
ץ��r��)0鮍n	_/���9Vq�Z�@�Z�wwg]j���Sv'a�h_#Nl��q���v�N ���L�:�Y�c�ZAS��>Օ�����^�
Q��X�F]�x������6Z�Ɲ�ʑ�6��rYr����`�z�� |�j�O{��,���N�λ"ל�[U<�My�q�!�iu-s���ꦷ5#�/�EG�|��u
��7%}G�WR�CW�ɺ���?��'g��x��O�y���\Lk]3<�wg�n蛳�O��Yyq0+'M�Q[�L�k*���]Rn��c&�]��,��.Q��%>���fA�� .��^����!ţU��چ홹bb���[g&�U�����d)�ȕ�s�w����O��5�q`�b%��]}!w��5vbz�mD��#�o:Z��=��3Z ���HnWn�R��{s{E<�kS�)�V��m�	'��^��lѴ��
S�yۆ�5VQgkB�|��>��	Լ�uj��l�RWt�:I0�6Ղ=�ZN�S]��Ga���'=x�ڰ/���G���z��:6����;��x큓9Sō5y�u��o:ٮD|��\��;W7es��ivR��ӭ����v������|���G%=	]��Ҋ�JY5��c7r(g�_r���%����Q�]de�)W���j��P�g;z��f�|OAu*N�UY�H����y�t͇bCX���Tʗ�.�V�8�R*�Ս��|J�p���N/΋8jn���k73,��jL`
J�=��dݸ�A��)�QFn]!��k�[���u7�S3�39��}+[�Ӝ��o.����:F�K�0*)�$=����C���^�d�ՠ5Y/�o
����Ҭ�2A���G�ى:�LTz��ٽK-��+���ܶ�pt�i�q�][;#۰�p��쾵k�hz�<��5U��G�"X�s�eo.��W�(]�XJ�N>�U�Ho�]ۅ����k4��:��2�cL.�V��	���+.�U�p���� ej���<��5���Wc�^������jZ5��WjqM�����X�V�%��z��v/�݌���R0�۸m7�������r��-�{(�9�����;h�udEB�C�u��ݻU��������p����P�}�����M��3���;7���M��og-�	��܏uJ�����lv>��,]X^��'R�1Zo�J����)�t��W=Q�o�xi*'u.�8-S���{Ћj�P=��ʊق )��jaL�sI-ə[,YLu^���{�K�`d7s��n����o���;hY�g��)R�]����妎`�����u�����jP`�ޏ��N��@�f�z�3�R�������&�A�MLmHY*#X�ƈ�a �6��4c& �PA�S	��34I�Œ��EbLHQB��&$C&
�M�"���J����,0
"Ch�0���lQwqb�Xō\����\�*,2�A0ƋG-��v�h�4X9�ơ#ccF5�heB[�ѻ�6-�	���TX��9th�L؃�r�b�11�.b�Jh�����MrwFf���Ž߿��ߟ�d�XE�y%g	��t5h�B
�sWpUz��M�X4��TCەd2
�M�%q��w24.9Ae0'M;�bج��Et\�ӯ�k�jL�c�q�g>^�_����B�r�9�4w��y���}�,ߔX��5'�4�������{�?S��l'i?Lb-ߝ���� {���u�-�/3O�#��9���^�������}�y:��<^nwA��s���EV����e|�؎�?L�v~������mн�9s��{��o��k~�+��4<r�M�c�1E��2D�r�i垉��}=����P�p�x��z/%��9�f�9Ua���uz`�U_�����yw��2c_ȸ���Qp����u�]�l��X风X}���TH|�<����8�{wW�+�
���A�m�R��W����}�P&|�����4�9�v�#��er�R�-��8k1�΄��*�f�ٛq��3tn�z��H��^�t�v�`��x�U	=��s4�\�LR�!4{ں���
��`���,Z�0��w���������7C��suJ]�bU�x��j7�o ,�.�j�Q9�tiNaѨ5��=Kp�^��������ci�Ѿ�,sWP��b����b�ˎ���� �r9i	��2�.���(Ŕ	i�v�~_r�J��ݸ'3U��m�,f�S��b��5
n���'��uJj��ܶmw|��%�y�M\����^�z{�Ū���v�Y�3�*ck�T�L�Q�:m]:����5�βB�Y��%�q!�lf���\��o�b�s��&�(�9o��;rײ���~��M���ѝ�W�uO$�Pˌw�Y	��#!;���|����g�����χ4�g��kLFs�q	*�����k�&C�Y}38�p��`)i���z���hy�r�?>YH��N{`ו샳�=���L��oeHR��q	��8�U�r���?�����.��k�<|���e
��&�(SD],D��S����\�S�q�eA�H�Us��7�z�s�lw%`����������U�g�U��%����#������r�D��]�O�toqwo����N��	V�ZV4�8�6��v�?v�O���j9�>4���b�t
;�.�q�1d���4z1�XQ��o;S�p�S���[���,��\Z�ƭ�R��+&�T_��+8��,d��i��j��:�����D�ed}JVubd �Y�ұA�\+��-�ϥ���7�X��
R��4磛Xd�I�˘�qT��J��_laQ1|���ި�ϣ�J��swÚ��v$�ot����y�%G,��U��s#���]SS���ٸ{�^ec�����<g�W�U��`zq��_)E�]b,T���}m(��u|�n8Y��ht�}���ܧ�Gp��w�z��gb��Ι;�' ��V�!�z#9{�~�����q�!��e
ns��]��M�c�HQ�ϱb����]�[Jj����m��T�L��ŘK��{ڴ�h�����zC���o����҆�5����,SvC�-9�JJ�w�c�����թjxGk�Y^�)T�-:����J���&�=��;#�V���+��)0�&�)M��!�@�rs�O'�ٯ9d#�Œ���S���cȥ����W��8�)��b�BͻR��Z��9R���ue=�!����gx�d�U�;",�0Z������\��j�G�{�N����H��fɩD��&���Z��{T�e��;���ef>���Z�\'u	f���[X����-�Mu^�gN�.�ʋW���ur��&�]�9_}��K�����~�C'�Զ�'^sK�H�Ƙ��u�k�]x�3P�Aڄ�k��K�O����{�n/�~�h-dv���9�Ng�]�>y솗�����5��ˡ�p�낌'^�V�la{��k"�����+}ޞ??g�^�Og��o��}8�;�s;Ϙl��;j��*%1أ/�
�|�৫�8JV�<�[-�Q���y�Ug��Z�l��mV~�:���3�C�x��ӗh>�v��d�+K�ݷ�m�Z��kg�+��{W��:�}��V����d����~7�,S��qz�sЛ}r�Я�n�����Be�ftdOq��֛����qi:R�&������{pU�Y�]�w�q����^gw�"V�xZ1:�/��%�$�}�5�uD[ᔛ��+C\%bYs�UK�^y��u��;Gzg]"�抄�Z�=�X��=[��n��L�9�XN��ޭo�����K��ɷ]�
M��v�a�;*�)'b��G�
�3Gz����uhjQ?;��y�p@::T�Z����$pC�{O��ɒc��3v;ë�4�wA��ܠoY�{�w��`���g>&��E.������go�
++�e	��Ǩ�B[���J؅�R#a/�k���~�Ҫ>��wL򚌵6�W��Z]�I��M�.z��بsNh�
��.�B}5+s/�	����.���\Z�P�jH�I�2��5�o�����p�������'`�s�����|Y�yP�>y�
E��[��V�]SP�`�n5��dN���Ns��+\�fV��p��x_2��5���,��:�_s��N����*5��w�jqj'e�i�*hJb�����"[�^e��t�s=s�{7�{��pԕ�k��J~��j�$ӛ�}V��V�5=��X�}�;>�K�do��,4	{)=�8����~���p��4<r���8�'�o˩h�F��H�}������̞�=���)��ڼ�3S�����g�����^٢�z�]H4�xw���0�&���`fӮI�y{}t�!Y�P��G^�F�?_���!{�uu���ŵ�f�F�;e����z�/n�vC
�̥���D�4-<\��K��޻����kS��&� 멎���S�D}�˥Aڠ��呯
����.��>�{�ު�i�?i�6����r'� ��^���\>��]�F_ ܶީ|��Φ֗&Y�����X ��m��(�z���I|K崥+���юˈ�jOf�"f�*�Uf0 �������*��I�w�I�n�����qK|�--7s:�7�+�����?C��p�����8�sw���WL���;r�����m�7��^��#(wD��]<��hC�:��d�`ϹYM+�,�sBlm:�(��:BꫦġC��iv���<������{����R��C|��A\����2�<��V��s;2� G��f��m;�,�*�.��I�l��adl���.��\*z��w�z� �ׯӓ�#u�Əe��w�:��{�����Ws�Z����r"u��{�^n��y(8Vl %����,��YZz�p�v��ǳ2umty�+¨v )\���(=�:�ٸ����]�q�p��νup{�!jͶA{xC�J�|�v"���t�����k{�c %j�W3;-$	�t_&�k��s=+;xJ�Y߾�ų�k>������ꗮ�R��L븟z��h~�r��V�l������9���s�5O�r�����r�A�)VH�X�6�[���s�o�Z��k��,���??S�q�e|}���W(�
����f����5�&W����̝G��ƫ��8��%�q����L���pp�fw^yh�U��q*V8?_./�Z��dK�ۆ��Am�{Z�M�e�;3�*�:���U}.z�T.��ՅD����"�|:3F�QYPW.���I�;l�t����t�] �/�%G*��_au!������z�2����p�]:On
�W�������}W������ƫ[��e�Q.T�6���SyE�m��.m�8[Qo�����i�}��N���aC{��~����;m�V�?l�6�tFr�E��f��r��%��_r�����*L,�Z�>��3�<��o��=O֌X��z�6(�<[y���=��$7���ׯ"\�kd�n���EZ��x�p[DE猭 F��<�o�Hx,G�cT�8��,Έ��+�^�фq�i��c{%oR��s�)�'RӋg̒4Z;��!�(���Yjwesؾz추:Ս�
Hb�S��Kp}�9kq�6I;�f1�+����*�4��C6�L䩭�f^F�[���j_'Z���{]P�#�ɮ�N���O:���Z���˫9NG��Of�m��{���+�N��Snj#�}6V��ҞM}�-�I�MɆ�uqwuz���S�f���{��+�S�����A�_�'�ܷ��1�/-b� ��͍�� z�p�f�WTn���/��C�i9ʈ�O��ŻQL�9�מbk����@��g���{����z]����������SֽI��d��߻�禐*��'��߰���+[��wύL�v{�<_��6�;*�6[}>��Rڱ����?0�r��BY޹�����zz��6����J��j�ޘ3-�}�N��d�U�4	ʰ��g�mgW���Q5���ki�߬Gݖm���᫁G#�'!����7O�=���",�6i4}��SڻSuv��<m��~2�%Wc}���m�,7i类�����`�9�uՍmZ{Q���,8�V�c��:�ś��Μv,ݴfcTb�ٚA8�_,�N��۔�Z����_��t��5\D�������������L���0���A9�M�-<
�b�*xߎ��� ��Y,*�iq*&͸�}S+��JQ����>e�jOB��,��r����ɵιaSu�X�b`.U'��Ԗ�)<���~�������`OW���߶���x٢sXXv���'`��`o3PLV�h��
�e@��Z苇'e�Ʀ\N�x6�ʈUNi9-|ֈ�K�Z�پҔ��+r�{0��uE�jq7"��-N���^OɞC������)v]��54t�t72کP�8�������=����*�N��Snx�kRɲ.��>�Z�79��Mg�5��R|=��77�I0Sq�������,@�����ǎu��������o˖|����=�#P����S����J��fr���6�dk��st���X�[�Tf���La��P����V��Ӭ+�QFN�w��%V��j�T�3-��7G|�gM2ew!�m
f^ێ�-�|�bw�Z�z�b�Of������n��ח͓Z��]�j�ݱf0Bv�V�-����CD�s����^�@{W��^u�V�_�gZ��f�f�g���
Z\����<�2h���S��-M�2�F�;�r|����Q���n_[LFO:�����6�&��^�'��0�Ϲ�����ɯ��b|��ѶK�82}�
��g�$��t#��B�#__��c���ۅ��L���\�}�eF�5|�F3�����sj$��OG����ٻ�9�ܾ�Ǣ�CSzX
�K�
7�s7N���F��u�X���)�;�6�]�5FK���SnAc&�*g�o�rW4<�K���ǯ³ޯx��k������F?E��ᩩ[Yπ]H�f y�w�<��"{�}	ϭ�q����Ǿ�,�6:�p>̽��JE���d��;�v����.��t�0��2ٺ�Ax�[ʃR����<e���e�3p�|ૢ|{g��;O��6�~���G�]�� ��I�$7Q0Ǽ3�h"��v6�e��#{;�4M�p\��,3lv��3�i�9P�W�[�P��"�d���@Ȉ�Yk�vė��w��rےkPSW"�i��3$�ې��]fڷ"� cW���G��̚����u�imv�J,�u�!��+tv)�gX��v(9�dO�@��i�VY�;�up�H&u�"%�(���Kn�FT�7�>bb�v_2G.\g�{e�����n;+:��mU�][�o���\�04�<4�R�4����v��� ce����Hu��gt����ܜ$���QǊ�Ɂ�]z�2��x])�u�mpN�	ZtéN�H֜�e�b[Y̓f����$ë�$��A�)�ȴ�����X���T��B�[�7��:[�k=�:s�l�wv�r�G��z��N�Cv���i�K����S�{Vb��Rk.�u�xj�e*�HiW% Ep-m�90R��VX�[�@<��2�A��ӱ�++�>
��ۭ�j��j���6Û�P �{m�[�x%=��� �}�r[�������1�=1�{rr�0���M��|%��B��,sV��ey���yu�j�mC��R��3�^smf��ioC��6��� ee�A�bRp��s�hk6���}Bo�;gR�ӚΫM���[�����+2���,�ئ�y팎Q޷��S ��.�b�$�Os&�|4�
�S�n�/x ����cJ���p�H��O͡Ϝ���	�v,5"�4r������˫m`;��� ��j	v��v�΁ML��l�ү�Ri�_�fR�*f?���VF]��`q�@Rt�ޗ]4���CJ�:s>��N���õ6��ku�g;<6f�X�N+{�':iL�q�λ�	�K�>]����}\n�t�����$�xƒZ�7L�����X#�[:�F�L�mѹ;/i��i-�Pdq�]4 �����2���^�܎&r�ιf������8�a�L���r��g'��/*h��\(�u|��݀T��z���V��e�j���]�f�q�n���n�6��[��.�ը�z�Ή�#����V�P�U�s��_�0޲��E'|�j�m�u���+Q-CʑBu��w�V_�1]���k���RGX��)X�;I۰j��V�#2s�fݭ���̕ǯ�b��8G[��Y!6��S�d���!j=�,�+jO���/b��8�U�s{#\`Z�7n�[V�a��p��4>��;)����ܶ�����@&zN��5���g:f���:��h@}����ko�rY�&�s���rrX�Oz��5O,t�mqH����,��׸]&`�ͺ��4�[DU��hW+S�";tX�kT���A-��7{M����v}�+���9n>�,��|x^Q<vl���*֨Sͣʰt�|�5�CZ�/�'ס��4;���}ǞM[n�����O1N�]u�/��v�9�07�/��GFvT݁���K�_nQ,ټYO� [Ռf��ը��J�)F�Vk�r.��x�����b�B`�F�b�cbJf
"���5#ˮA	�1F���7u���1���d��Wwbɱs\��**�X��Dj9�h�c.u$�ʮDd�����j�5wv��A��iwj�ė5N�EN�D���ˋ��$����D��Q����Hl.QE�`����rWwQ�ݮjB�$��l���X�㻅ni�E��W4cQnn�0�Rk�ʍ��������E�Uңr���J��-��k��M]��{�����1�p�9>���.�}�&='i/�Қ���E��Z�����՛4i��>�NZvP����q�)�e�X�%OX�ݳb��j1�p�~��3��l���z�p{�U�C]UK6�Hj-�e�VH����t�g^5�l�3o�0���>gp_b�����1�}�g�=3��\����#�{(��Eo�K���Gh��S$oX�?r�td5�XX�ԮC��	��>��� �6����:ם�j0΁�=�z.�TF��F�FIh��/�p�~9Kj�����]R��i{cg�:&�3��Y3��YS��.|�XfT
��a����2�i����YD�W�����t2��N1�����6�Y���n��G58MTkS#��\�`���Nr���NUd��J�W�v_��D��x�kr��d*�|c�R���U9=���ax8��p�ݷ��F�PO5W���r���n!Cf�Ta�ɺ}��|���/���{�^<����n�q�/g�?��y���υ�%���;ō���t�+�`N'hj���2W��[���z�-�}4��W���R3``���霋8J@Ǭ��q�n)�l��]���/zjGRur}F*bա�*��5z��&^�<��}E,5��V�����^��R�����kQ�SW�f]�&*Ę9��A'�����G�@R�z��e���u�Z��iL�6�m����PB�z:�u;F�t1G�����J6��B��d������d�ˤ̏!�.�C��=�!Q�O%�PeT;���g�fPS�Ę>zN���znS�wy��^�U�=�^��\{�s��ò%��8Β��IU<�*�T�s��R7���%�g��U>���Ξ|C�x��m[�m��u�>�pz�3�?z'�W��ɺK�<}SRHǦ)���{�$����&���׸f�89�Pm��#�/b��]Q�g{E���� tq��SSY �ؽ\<��;`z����wy�\=Q�kϺ��7�`QU �Rfp�{� p��u"�K��&�]����7��5���׷M�����^S�8~u�\:��W�T���-�G�/��n��U��gp1��۷7��2���9�ި[���U좞��Ƽ �dZ?]�uY꘸S'�G�ஊ��Se���t�[}�>�����?-�Y����+�������P��;�0�����s�.z��7-�<����i�롘��Rm�
��vU���Ϋ��sKDvy�dS�蓵��)�֦�MC� ���{-�{(��F��(�:ָZ�l�C���Ysb�$��Yw{�5���Tv*��k�G�c�m�CK���,N-�����{܃p��t|-M������淭��n�,uwA�![&l��.�ab��D@;2��������:�e]Nk)Kܮ�=�s��]^���<���q�9<���K� ��K�J�ӑ��\\Fy��s�t׍,�\W]�_�<�����7Th���2e@0�D�������H�>���1U;�q���3�\xk��7���������N;���<֑�q ò5L=���L��W}����&#VD�`����o�W[b�ψ��c����{��󮢱�i,vD�a�=P�+�H���N����+׼k�{ѝ��3s逼Ϩ
�s���:��g��q��������AZ�J��	�N�F�Ņ����<]�WE���Ve�QQ��&��x4;����ϫ��ݐ]j7�q�r-I]�*�$xx�j]{��.�_�3�M"��%�=nh9���<4yK풎���q��>V�>7�����[[}ݞ��Hf��8�'��$\A��d���o4H��:ɸ��Oó�֧^�ؑ�S7y]����z?_\,�,�̈	ј�[��:=7��D�Kk�T1~��^��_g9�JHw�_�kg@��4'*!���3>��@r �p[����A��Զ�Ys~5�.W'Փ��~�ɝ���5w�4/�Lm�`��>�
�?r-��ŧ2�'0�żmb���Z�Z(4"�@�6�>�k�`�ْ������������� rFţ�fR�cΛR�t2�.h�'>v�Jq<n�鬄�Z*�=�q�pؘ1���e�j��y��(�A�p�W���7���3��������U_�\��X�RZ����?R;Js��flyB�/�����L��j�F��|���>��>�6�׉�W�ڙ!��`̒<��\��u�~��=�I��,��(�hϫ��"���Ey���|�!DkSBd���ubx'��u���H��AǨǺ���!A�ed�e�U,m}�����\c�2�|����E��P}32�ێfB�q�yŨ��$t!rN`�Rk0T!�n5zrTe�צ��U�s����4k/�l��R�eLs�?�U:��y�;\�-M޵ b�r�Q�u����)�a8f~?���9�!nBr�G�������i'�_�s�\kI��Ƿ�Q�kˎkd����'�
�����G*-�O���_ewL�;��86:&�C���K�s9�Toduo�c�cZ.��Ν���q�a�W�Y'^~��TN>ꞣ���jn4�}��
���x������Ҍ�n��+�~�\/t@�Q��VR��h���o�te@3�	%�,�{�s�K��1��z��+ԇ���}ۉ!�4f׷t]�ƜDE�N�E4��G�Mb���@�R�r��}	�_�o,Ƥ��w�u�ѯ^��o�_*�/��[-�}�:ݭ�V[��h.0�����N �Pbŝ�U�l�5jB���lW@ [\�.�zy����f�Sza/r���m; ���u�������?f�ov����$��0�K2��>	����ϸ�׃#}�v�/f6�6�ȋW�6{yX���
��_�'�H<�;E�eX1�. �T;�2ْP^=o*{ױ�f@x˅�N���Fi;����㷍L�7�TF�UxyG�]Ðs_I�$7P*���͹�~�g����#��=�jˊ}��:�<m�ўfpmC�Fq��y�%��	���꫰<���P�2������QS]��we
�/�b���_���W�=��*<�@֒aO�'�6��P��מ�Ƒ�<EߠH ��к�����]��C���1�}�g�#�8�y�򌉑�b���S��+sޛE@�aQ��2CV&�Lw��F����_�,z�+���ڻ�i��>�w�� ��z�ρR�E�@��*!�.�T/e���#$��1p}�0_�y�U�=�g<�8�\35G�,z�y�H������:M���>Ȁ�k�Q9Ղz�T�E7>��5�����%����X����r���م:���y:��je�O)zV�Ct�k��&����`��+:y� L�5�rs"jȞ��l��h�G�=�V��3;:���ջMD�(�!� [��'p˫U��R��1-5"�q���%�#%���s�)�ru���Td�ɽ��7@�f�5��s�]ի�V*ќ�f��FL\(]�L���S��_h�1�]E���GwT�g�l��,<�F]mC��S��8\�2\�����S�i���d9�ߗ�磡�y�ڪ��ۉ�r�C&��09���vC���/�����Mx����N�p#ȸyAX�{���"k��3��u.+&��9�e����\*�;���M�׻�c��E���+>p{lϬ]��xz5��G,�)\����T;��R7�9�ڡ��.�Y���}1���켇Ǭ�/ۅ?�������=q�п��}rE�$�RZ5UC�3�d8	�ʔs��������`���A��8���Ǽ�=n�;%��8Β��(UDL��0�\r�r��i/��u��N���l\W�k�����1��f|6����}Y���:7	���Vy�e����"��}�M�s.p�B��b�D�9�n�Mķhho=O���Hү�o�'n=wl�=���Qк�s;�z�K�z �2H>��J��tb�����������{ӺN=
}K��&�������zT�+�B��f�ʠH$�T�����	��1vHa?:`�B��S�j��	�D~]7�6�+��F�v�����Xe�a��t�/��OF���w�}�UI�O��ܤ����w ���H�!f �9n�lU+_ ٻ9��#���v%^`�;���;6@��J�MT��,�K:��I��=�P��)�9���cy������I�`�7:C�[3P�;��KG8=¾�'A�Ф=�b�1ב������|揅��8o��T6�Hv=^ o�:�)���۪�T��)��6zlQ������ ��4U�����.�$C=�]�=�����&����σ�}�E/VS��s�}�6���W��3����wFI�>��}�9R�g�Ϋ�g�G������9Z�ة̱�����I)S@�K��6�t���Nt���C��x�>�~��^�f�.Wv�58���9��p=
�W�V}�A;��Z'tø��q�s���0_���S��"#�2{�C�3@K�Xy�8�����㘫��/$v�{��!���Y�v(��P$��Q�`����z�2�!�O"=���}�<���9�)��94�Zip���w�����c[�����R>�
���9:^3��=�O����c�y΢�Z�J���ǩ�Qo՘���}8�D�1I��5�|V�07�Ϩ���>�Y�y�{��F�ǴZΰEŲh �D铩/Lr��z���VޞAȜ���/��Q�gZ�����V(�`�Yf�ݛ.�T�+�; N������qb�ѻ�OUX�x�!����%�yY�)*�ú��d+|vp+�/�I��W`޵�eiŖ�%eM�x��g@�sH��_$_x���Ƴ����k��9���?:�n�~�r�dFZ�~.�S@N��y2�I~�<�)+��l�T��m����ё��W��)���h{w	��m�����:�q;��2 'Fc�In���J�������5����M�xDK(W���h�T�g�}��\8��z�ۏ]�q�S�@r �e��_T���v �Υ��5c�d�{�Co��7���;Z�z��U�����|'4}�|H)p��7�?��+��g�+FM^=��r�8��>�����_ Ųm��|�ey�`M}�i����ڨ�M>��G�6%���*FХ�{��zk��T�q��0��)�}��Q�d`�op�fd�1r�W�;��2��2�ּ�Fю�;b�ed�ala��rV�K�t/�9���lT	�3^��cϳ`��^L���qF'>}tH��hǡ�lW�o�l�y��T�[�h��]|��D��86�u89c+ۅ5!��ڰ��eN�s��7o��._
�=J��kG�&�[�f�X��/ñ/�Tb�U�E���y���vj��9����I�q4��눵�DQ�^�o++���\љ�n�i7XE�U4�x�j��c:oQ�]�f�:�:�ۄh�,��l�=,C	��j�n�7h��ݾe��"�w�K�!��R�9��;�o���e?^��US�r!��^9ޤ����o&���!��l���O������=w��}G=�`*0z$�{�Ǒ\�����[�mڌ�Ռ+�x��{��j��9�\T䗵��<'ցjq�(z���h�r��O�U��^��:��;!;�ݸn��}> ϜWۓr^g���[.��"���,e@3���g��!��G�F�pF&=~��W�TN�~\�����5�d���[����VQ%Q��5eS2��>	ө'�޼����ؿ+��'�=��������m|�1�9�y�h�q�K�1�'��Po�Ax�%�H2/Ϯ��Wy-�ӂZ��н'�{} =+<������=��/�r NjO?���o���.$����:o[�wՇ�g�ȴ��n[��m�ўfpm<tg+�y�%�}���W��3�VQO�]�jW�9></j~�*ңW��m��>ζ�ǦwI���\�Ux���Y�DC���8��}<}
���H>��x��uH}	�s鿃}A��M�;dxg��-qa���5��,x�f7j"x5�e��&]�!���q���[��l"��+כֵ݄Xp (�;����/;"W&헙�u���%1CH/c7Xcuq��*a.��՞�s^���.
sVqS���os$\鯮5� �V�]��C|����>frD~��LR�k��g݉��e�V�r��Wt���.�z-���a��_r<T�x?�;3���d���*�W;��}���N�ڳ�c}���C�����Qh�'�� ���7�_�������ˁ�73*����TBk0#���<P�Y�/�찬�����/rwh�P�~ۦ+�޺k�p��jdp_.z���S_"�vz3��~�?�.��^���Yu���S��'�^���V�G�M�׈�\ןa�wv~ܐyN��i���p���C$�����M�ۏM�]뉳�[�p�Lo(T3,x"�=D_V����{&n�/� ���0�D���VV
��2��w�S����
�0e�e��`P��3�Js����r����>�G"��1���&�
�^3>�&\�7��������ڂ8E׀槒����<�ԇ�){h_���,��D�jKF���Q�"}e�Ƿ�O�7:&Tz'���xv4=�G�#C|K�s�ֶ{$X�z@���舾�lBv"m�3so�����氵͙-e���TV��gn����֊���nΙ���1s�wqweId�
]Y�)) �'~��UT���:���;q$�4�ʲ�I��*��o�H��(��X�x��3�lי�}@g�]��L��?q�I``�/N���3�*�ܹ�6_K|dv�az�m���r祁mo]��s�:e����^�#�Awm�o�
V�Bq��s9E�T���С)[�@�K'*�.F®��ʖ���gMn'u��:{�����;/i֖0�F�9ӵ�G��=r�v�r�œ�=��N��:�=O*qY���}h�)�N�]��:V�3GN�2�kv�q�6�
���;ܠ\�Y�}y{}�Ѕ����c�7�9f�d��hqCE�����I���D�S{�ܵ���\qUڄY����+�Z�=j��qZD�����r���S:*� ӑv+0#�0���	e`����N͞��`J��)WJ_c"������oa��b1I!tpX��{��3*�>-XΨ���y.p�W"�ٚ��έ���ѥ)d��[��ٻ}e�3�h��1�#{
�/4���T�*�/I�1k��i4�JN9m�<=�o���d�����ԝtr!Ə�������3FS�76�w
�9��H��7��'�������<;J7C�Zƪ����u�We���AM�2�rE��̸NTR9}�n#�d9[ȻU���\➬���n�]��԰�L����;y�b��0�h'mRyl�u\=qQA�;T�=�}/��[�4�-�ɲ���δ��'�ԫ�7��L�3�c�j���}}��壙��n둏_G�8�nګ��]t����z��4�ھT����x��캜u�dB<F�!�5zt��s	w-
��l�Io{T��'4�Gs��	d����Djn���Zy�:E��kVS�v��6�R�,�6��⻃�C����=��aem�Q�ef1���8`�]��m�֜r�kJW6z�l����*͊�uer�
�"�b�.���g�*�GK�r��q5g��s��hj�����݁F�'�P
�M�M���a����J�f1ԉ�/����w�^VU��a�Ut�H�][u��d���tl�˭R�ˡ���y���O������K,5W)��hO��k���7Q��$���:(��Af����K|��tw9��])g�I��w�����وٚ"�/����1Qu
F���{戲U�[6ͩқ1ps�G+��4�L���po$wX��^�3�(uBe���EVپ��x)�4ž"��f�����zŷ��R�;�Ť�k�9l�k���.��WNb5��V�&.JG�k2L:��	:G�.�5:���!{�A�DQ��Ep���P�"y�`�e�	������&B�vq� �D�s)H�^�gsf���:p�'#D1P��Ose:��Cj*w�^I�m\�x���%>�!��Wҿݭ��ۙ�G8&9�]6�vCsk�.[���P[�+qݷ]�1ȹ�h�u����l�(�(���mQ���(9���`*�76�%�sFJ�k���6(��\�5w%Q�lmsEww.U�+�rJ�&ۛ��-'5#����79���+r��C��bы�76�7wh��WH�-��8\��sc�\�9Ȩ�n��6�[��W)ݫ�ܥ�λ��.n[��ngv�둥�t��]ݮ�r��wnb�&ܹt���͹0�����u��E��\�Dnr���
4�Я�����^��E[W�ԇA3K�/`�H���)��v�XI�}1�U�EV[�Z����od|��/��E؝v�\�)1������R��p�1P�]�q^+��{��[����f|6��+��}Y���:)G��c�ͭy;�M[8�&<�8���i�]L���n�Mķhh�������G����p����ǳqC�P}:c��OP@^�[ +�k����^�>�2������;F�]g�������g�oΠh�^���SR͢ 5P$z����k;b��?-�k��OcN�<��1�x����<g&߽\���n��Sh�-$q���F�;Id���*́=�G�?#Q��W�7ޤ����X?]�3~���L�)�=6�6s�=�z3]kH]��DnB���f�*������3�<LߣZ��Ե�M��
��=��j�D�&�z 9��*V�O�_a��u���W���x=s|�Ng��/�;�ۏ�4������@�t�uN,�P���P�p�=-F]UϦ��O�.3�O2o6��>�հ�\x�V8�P�s�J�F� fT���6�i^6�c�U��<0���-��Ra�Y�!D���'Xk�^����ƶ����� ��-�|3�� �]/��6o5����>�`;��]�c��O��XY�W��Ԧ�P] N\�uj
V�}�˰�ܽ��z]ԁ��s��;t�_7�v�i��Ma����F���o!9b�=���:i�x�����%Y5�2���洍��v�6NC��v�Ѐp]�Ff���@���d_��dg��Ú��=�"<�и�:�+V��vA��7ޢn�3����(���#裐7\Q�����P������b�κ����F@��U�X����S���%��L��."���A�]]@�N�>��}��"��=�֢��zS�cC��W� )]O����^���$��ԪB�|�幠���<4w���{d���Y��U�V��-���mT��u�7�:7&Q�̢K�<��"���qS(/Sw�AoՃ���׳9F<T:���v��:��q�_�H��t���,_̈	ј���=+�n��ʿKhmSW�X��4M�p\޷6��s�l�7�{�F߮�~��OC 9�G-�	����ћ�7���8�'��|��
w�{��7�������fi�L!�IaI/�c���Y�;��ta>=��U�R�tn@>f�q�w�j�Fߧȟ�ͰϖL���0$�sq�b�\�leb�+�p^WV<o;$k�Mu`�˟[B��o]-�]w�t� e��W��F�T�����Wv�O����i�sk �S�N��/y�#�Ĺ����	�s��7iE�d�|1 ��$�R�*��	���h�����	�ྲ���Π��Cs�{b�	����H��C\�O3B��J�W/N��Co���m�̛�2�u���S~.ܝ��듓>�1����]{�[f�Խ�0[����c1UXa%�S�D��>���m��RGDӜ%�vd�7p�Tk�Q*]:��{k�9�=_&��`y��9;��E�K�q��P�͆��K�.<����R¯�*�--�9��-M�>@R._	�1��Z|7����;� U�dc� 1@X����[]7�/h�'<��I��yW;v��rN�%ؽ5"#p���Ϳn \+~�kUq�+ģz\	��ǲ$�x�r�y�z�/7�uk�3�����>O���u㱾גA�W�pe|&t9*N��#�oKV�p*9z׌�ׯ�+k�qܶ`�c���VO�ZT�N��я{��LвR��3ŋ���7�9�١������U#둧D�R��O���W��fG�7�SN#�ڟYD�y2��%#2|qn�9�����Q={�V�Ux�}5�R����3���[���%ܠ�q�,�(���t	��C���gEz���;�`���uu�F��7��x�N����.�pxxY������֕Z5#QVu��(���E�hB�U�ؕ�:�����Vr�kb�اZ���/�j�6n��C��	e�x)�ʾ!�yr,��]1�$�^��
ms��nL^�q*�^�JR�΃=

����_���J���9>s����|n>�*#o��g�]�@	�|F̯\��[�n�����,��K�d0�l}\�yw6�h�386�:3���i�dO��CxQ4�����o�𣞉�:~�@�ޔ*�kgC+ԑ�A�u{�9�Ty����������[��\�*�zQ��uU:zIp�:jhe9����]r������+>#��A�n{��ϯ���^�lW���u���wn��F�L����<��FCY5��Ǫ5+��]d�f+�q��(Z����e*j_���`��w���&TG�UD��tЮ m(Gڳ�1i+�:d���y�>���_G���\=n���?Po޿�����e��:əW���;8����Ϋ��֤�<�g0n;Z���U��3�L�)�/J�n��}�NU�L�=����x��VV��29��:rz�Zs�� ���o�u��E=�8:ǣNeg�ׁ,�0�9�f�Oz��I#uG�F���d���#hd�.,��>�7~�1U'�2"_���`����6���Z�ۂ���+7��{���|D��Y�={W���c�=�5�Ŝ�ܷ[]k���㋪�_��Rms��{fE�ç������2��
�������A�3:��.��@(پ�7�R:H��JX<���������%nlr��/,]��؇�2���΁�p;tq����)���c�
�Ӂ�2�3D�uG���#� �����Ś����R��H�%+�0���q^�F��!E���n��X����z�Q��?Ml_���}Hxr����Ǽ��,��IF��AS��Sb������˜�x8�.%�XK���S�|g�x�7���xv}/m�gIwP$����^���W{�����@�Q�S/�}+ǭ�37����}�φվ�����a��h.f�/�޶-.�l�>�l����&�ۘ��Oӑm։����{�h�s3��-[�vk���*뷮yX�pSuU�:L����� u�-�+�Ҽ���X�����}>�ʞU� ��Ξ~�*�����{��M����z��p�jY�D@j���`�T��/O�@�i!�gν���}������M�R��S�����87�������~ȧ3>�@���4����4I�^p�c��GRl$�Fp�H�z�W�6��@�>� 7�`�~��i��q!���M?�T���l����"�L���Zu�@�]o}��1h̘(�ơ�&x���e_-�-�r�T�y��x|,V�H#�y.�i�^����S�k%�]o�D��.G��.��)�7ӆ���S=*c��j<�rk}ǲN�:U!]k��G
��9$1#\�M���lG���Z?1���ʇ�ۻ�x�x�>����m�ޡ�L7&���=Z�gs{�#�qq@����t��#�2i<NVXȌ꺏_s���p���蓪��x�Sy6�d�Q��� ���y��b�jI*�Ly_�kC������^a�j2�};��G�Osc���O5�ȉ�7��W����cX�.��/���B��R��Q�3:�^	=�e_��Qqϲ�������ު���O����/x�Ϲd�<�S�kH��1�5��PKW|�w�=װx	��+����&��.W�.|5t����ϭ�󭢳畤��3�^5����b�W���#�oSZ��%�������x�E:��e?\og�c�u�P�ϺQ��X�詥5u����J&�A8;�T�S�'7���W��
����/��<��=��A񾻡2�<�U작>�>����9jH(E��T��UO���sA��k�xhϻ��cr^R
:�&��,foT�e��b���b��>��Fx	��}-�������"�����G����P�lzh{ݬT�o��s�]1�'��\���(+�n�N^����R�h���b��ˮ5�Q�O�y�����{�FZyu�'�W���򙽭�xɚ�.�ni���#�B����mP4*�Ϊ<�.��;�E�v�I26�ZS�x*vq���u:�oLܦ�.ui�;~A���{��*�ԁ�p�~��@��D�����-�METo��xO�V�9�#�d���&�W� ϑ��Ѥ;m	�uU�U�f��f_��'F�Q�T�M��xs��z�L�g�z t�Ya��c��y׼.7���3�$Ty�ٚ��0�����	���wt�,��bY˟Gt�Y�K�r~5��CMW��ĳ�3�'�� �w~;v,^cǔ{}�6����'Aƒ%�iSpY��;ll�5���UTc���2e���>��f��^��y��|�!Dy��2��i����߂�4�{�`�����1�Ic�tuߺ����uk����t=�:
f���O����>�$uDяmDI����[�C���)n&4ٞ����{?^Z��SGz��_��:�ȏzhu��nP��N�@8<��ڇ�U�b�/<��j�灞�,<��i��K��u�s�U�+#}٢߲����p�<�9~u�.5>�׷U�%��J��Q�%������&{�����eF�|�����7���Iw�1u�bB�[�����o���lc���P���ʣ/��(Gٯ/xCT�����V�"�	\0�|�b]�-�C���4��Y:��2��i^́��yd=�;����}VF�{���*�U�}��y���V��wݜ�h������:L�Z:S^g~C�,�K��/Z񁎽~�Wj�5���j�m�*��8�����1{��H��p���� �.�|��]4<�:�/1���_��Oh��Y@��h�G�M���C�9�c���>9�Y@ c���U1u2��>	��!:��j�[�\�}��\0�W7��n}��\C���9/)��h�q�K:�*���qY�IK9�\�me�����p6s�YPjR�x真9��P����^Q�t�n@	�mgD��ϻ�s9>�"�`FG�Q�_����H���x��g�hʹW��+�%-,����׽�0m̞:��L��f&'|�J���l�N_������L�Nf��q&�ߟ����k@����,jI$�e3�3 ���:�jB߹+a���RBM��Q��r����&����6C��✙�S$5bhD�>�Q�-l֖=���/�nH^�Ý��NF��UG���0\�;�TdϜ%s�hW��N�^טRz?+*T���Ʌ(�*ȧv���¹*IT��0�)ܼOfE'�*�l���qTV��q=0��UI�įnq������#as����V���5��!�u�k�3�Ԭ{O��W������<�X��Pw���*=m�R{�Ϻ]A԰��WN�����������7�@9�z�d|���\]D�$�D��hP%GE��/���e���qV�7�\h��WQ��uh�k��7ۦ+��z�u����;����([��J�%�Y��p6tu�Zs�� �_`�F]mG��E=~��_��r{3å��@�f���c���������''?L�*�����:%����vC�O p��1ꁑ�`�{��N�'�~ep��}]�+e-�v��W�u'�@�-�(��늇>59YH����&��C^�\M��m�����oWN?b\;�`wT��Tz�K�l�����^�g�t�2��HpW���/zk~�W��W������#=�x����h�A��>�0�aſ�l�Oxo�OOV�j���1�7Ŀ9�}����A�<h{{6�����o6���q��@���3�C s1����2��u�>��O��������Ч�ɫnw���̆pk`�
�@��b���.*e?NE�Z&�CF7���S~��5>E�LR�9'V,ṣS�ܖ�[�����,�G7���������5�[��{]6��L�c�_�yDyul֪`�2>Ie�T�u��k�����6�T���ڭչa�U��;E&k�+��|w��eū��.P}��hS�JǛ(6ް�b�ok��L��M�N*�f������:2L��J��X�^��T�n�ɿ,����~�FR��÷];�6�@����Uz��MK6���	��^�^�����:H�=\zGtNC�_=�>�o����|�g&�~�p��E[��V���q�g^xzI?H��Ⴓ^��Q�;W�f�#P�~�qޤ�z� �`u�S�߁�U���Yl���^���W���C��AS`�N����8�eB�|ۻ�x�x�7���@uCey%�辌����Q�B�$�}��:�ύ���/�'�\��>����=}Ϋ�^y�di[�
�uL���363Ը�\IN<����0ؿ����L5p6�;������lu���*�e��l}��V��'�+�W^�ߔ���)�׎�h���)X��f@̯���3x�x�Ⱦ�/8o�<���	bA�� z���U;�q����k*^�}��e)��ZF�t0g(��}=1Ғ�E�Y���8�8������@���P�ԼF}.�9��{k��>�/|���@z��Q.�]^]7]Ld%��KJ��|�K�D���pž�v�C�R���p��	vхլ.���c�A�h���7�.��� le[�P8x�S4�Y�*JO�9��gRx�*v$J���;���H
�BR�"�M�Y�Y��[�/o��pu�/�ga�AE�uuz��s�kgu�6t]�{����^��W��x/&O�+:��\��[v5l��/{��ǅ���%�h�.�zZǛh��	d�f��Au��gp9�o�-��[0�׀�jԎvEQ'��E��99L��S����w
D���}'k��,�^Kc��N�3H� ъ�Uf�-|-ɩ�(�����6��-n�V�����_ڲH^�fm� BĮ��0a�X��:��9ٻ<�+s�v��F��l�3:��R�c�^�W�2�̮x��H�V���ߵ��OI����嶷��a��=2��޾0�[��]:�����t�9����+��Rh�����,Uv��[j����y}In�k�]��Fݻ��ʣ�+����1i��:���F�yܡ�GJܷ۹N�t�tf,�tw� �gL��r�*��]Q��5��rD�e����HE**���;)2'ur�g�3t��-wf�RݴT�L��s���j�1u�~�0���u{��)ڇ����ɖ�RdJ;�1�閵�'ѝ��L^Wc��a�vѶG�a�Q�E��4r]�2�m�Ι�>7�t��l�A*�ė������*����EC���v�.�ç����9�H����N�d����m(�p�M���ڎ%̌Ev��35��5�姫}�,u�B,��>�Ru��aA�gS+�ss-nkv�`�:L�ʖN��r�w;.�hܫ4sb̜9�6I�:�T�uEg��w{�_2r��r�f��؆bsp>E�!�Y�[]B>�Y:�	��.D3��'p�.$im�ٷ����(m
͡�`�ΰ�8�v���(Rz��:75\	[���o��a�$��>��p�����b���a�|\g�w`��{E��m]ËZ�>뇳6�W%a&f8��7e�(eEg�ma����`��Ii4(Л'5j�X��u�S
e�T���&4����^�x�$����Wc�&���I']�yy��{J�pJ�������;(�n���<r�]��Mv<���滼=�Qɋ:�M[�EIm����ӱ���J䷊9��k:v�
`<ȹ���m�V�d���˜���	+3�%]�G
;ŕ#s.�	E���p� Pq�7���e�s�Aè$\u�G��)ZX�$�ɶ���,�H� �1��K4�S6�3��duqd�).�͎P��qe�N��7��j.H�e��U�Z4Wr��Ϸ��������Мi��1j�<�Ó���x���EO����fl�-�zz{eQ���[��gJ����\��hw�Y[���c��v��N���e��A;'.�9L������sW;����wYܓnb�9�wi��5��6�Zwk����.vku�
���Us�u�����b��ݫ��I���sr8mr�s��˜�ΐ���,nvZ�����j����ۚ$��]2vvn�'v�5ݣWf9]�:s�6��.��2���\ۘ��E�\�N[��r�c�'(�w&�˗(.�0R@�F��;�����Q&�ݤ9�b�Qr�r�,QQ�5˕���\2��˗76��h�-.�;��"�Q���m�r
wK�Qk�r���W9\�&����A��x�_J������x
�]'8]]N;�l�	ם�/��V���:J�cmcGr��\�d���f�y
���&�Fk�s��Y����\WUq����Ѹ��
�K�+���2�:���7�<�N ۞�W��F��PکX�.+���v]"_�^3�5���>19���x4<�c\�٘���y}��m�8�����.���T�3㖤���?�X��T��U>Ni�z5�<4trDC��̼�n��^w֤F<���=��7��ɖ\2�.��
D���[7S(/V�
�z�FnP�~o@F����VM����jpuE��0{��!�S�l�	ј�[�N�{�����ܵ����þ�3�c��E��&��mb�y�����{�F��������q�3/ŧ�t�yU�ex�9W��l1��oj���>=��C�O���>���b���7[3M*a�NR�?[��JZ��'�O*��7H	��/��\H�
�B�W{��^e�\2m��`�}~&*���g;Q2����U�E¬�F����'UH���&{���������1���lֿ ����tT�9�2[9���q�M	��;MBl�����O���zo>Kӑb�7O2l%2uY���y(M��[u���t�NP���S��3y��].�/3���qʙ�ƺ���,��n��Yk��Y�2s��WR�ڠڗt����\t��`��G{b��R��!apO;��Aj�Y� p����N�	��\�����<�T���S�j.dmC����(��Ϯ�QF=�3{SY������/�`��z$I����t��ʩ���<i��S奰g7�w������$\�mU����*���y-I�q�t��a��}�}ld*�|N|�x/��W����f�n�!��P~�r�ÑyӺ���>Pp/EeV����ap'�^w�SK��5�ڌ�ר�+oĚ�,{r=����gCl�#�~�4m�77 l���ɥ�/�`��d�D�o:�"b<¡�4�89Yr�9���m;�ݿ:���~�\�)q�2��Tϑ�rW�� �=7�>�S{;��^�=�a��?W�VW� ������>9�YD�FcȂ��%#n��޷p�d�~n��z%����Ԅ�i��%�;����1�*^R8�o�Q%�':0�;�搷^�g��V}��H�<�׭@G���?�Ʀ}����uN]�8���t�;"鹙�y�X9h����N�#�P(9L�E��^ۉ��[��f�V��#O{}R1�4�����ḫ�����yQ�Za��Eܳ��wAg=Ы:2��|��V�.�*E�����u�H^�}2������u�'��)��i��k�Q�����%e�wY����ahZMa=��2���PR�ћ���QU��T�6폨�6�jW�������b�A��d��
�~�+ ƣW�K��c���yv�V*�ߑ�mnԝX����>�KN��ݳB��T����	�$s⦗���.z��Tt�#�
���xo!�{���w;,=t�d߀��-F�����qNL��!��4"c�W��k&�[��&���͇u[c@OG�R}R8zWts�|��|�F �P;�^���@|*ҍQ�� :Y�>��|���m}E#��ú�߆Cn���?Pn=��x�qJ%�N��L�^GP2�\�p�/����-Y��x��G�Wۗ�9z��~�=&�=�LWd{�C��5���D��*&�x����	 䓎5���},�ꈉÒ��8G���̮�}�k�c�R�Sg��}>i�{����G�ri���r����$Y�'��`��|���K��2��d�=��ϣ�q�]�k�}ҝM.�;�h~e1����Ec̥��:�u�s������x̾������1���3s��{޽zZw����Ez�w������r,�)_�aᯆM�'��չP���Ӱ4~�h�5+������p�q�±6�_^�wAyx�h.���}�^N�Ĕ��^]s�t�ﷰ�F��s���R��iR���ǫ�kX;�`�#�y������W�%v��
>x_���1I��=�kC[}yQzw�x��:�z�.�:����Ud���Pa^�@Tbt����{�z��Gֺ[�Fw�x�V?�6��Ym�"l���*�n��7E�L��2��>��G�{�yN}�^����q�1�����\J�K V�8'fL�(t���/�Rg>�4��kw�9�'����Ig���>Yeg+m�B�DS����נ�,��	��& )@��sS)�i��=-�9�*��v�v��tI�o���{���=wl��ڟ ��0d
=+�k>�^���~����wܴ\�Sb�|���iNwI��G��qV�k�Uq=�@�(��u�^e=.���Ugۆ��cʱ�H�O����}�l"}ޮ�W슸�U雄d��� �y��W��~^I`}��a�Ǻ����{Q�k�H�;��~�p��@��<7��s�:� UA�;�4�nr�^�l�Ω�}
d�d\J�b���(�x{{��wE��L�y��P�!��n4t����>�B��6)X��`��aE/'+�_*Q����L$���Q���f;��:��X��k5��]��8�u4�rf�g��8r9h��m#���[�*)5�,��+G5}���tzL�ū���!SG<�͆V�#k]��X��������Z�C�s�|���S����*�J�f!�����-�V���;5�É�3Q�!��ؓ��)�fhC� މ�ډœ�E�ɨB���K�+�W�C��ɜ����u7.#�{�/�mK���uEDy�R�q���M؏/FEW�Q~�ʬ���Ā�E���徴2S�>n��9�w����l�)N_��7lv5U<���[�{݀B���X)���g"��Q\Z�&ϓ��o�\?mt��͑��6����v�^oNǒXdD��9��3����P�.��p;��J�+��x�K�l�E?\ox���y�QSK7d������{!��ETL�('�ʙ򘿩�f����U��V|}G��'Q6hn��w1�t����?�Q�,֌�x���u�H�i��1u*����sL�t�r6�����/wؘ��U�'P�}��?:�j.�C���w�x���,#ųOI{����j	q��v�S�䙨>n�m���Ƨê-����ΝC��FW	��Q �D�y�w�>��h�-̱��B=�}[Π�D����l?To������wlU�6�!yGݚ��y�V.�K��/F�j̼T$\A���[�,�X5����d�����n|;�ǹAH�U�%t���N���ݩ�W�IG�t�X\{�yݘ��&��hn�.k� �,���c�&�q��{�v(�[n���Nw4���z�q�l�q�� ^d��u�x7za�07ٛ���l9�A� N��R��j�Ǵ�b�p����Ӝ[;��kA��\v�h�^z�$�5I����%��>H�ڒ��C<&�V�ρ~5�.5�5~��O��{p��X��l�愨���"_��zi��s��(��U��s�)3��y���ȢZ�����Ϫr���(�'hC��К�.']��FG��&n9�hTp��"NЅ}�Y'��Fn��7k"�xw3�qW��D?+��>�wt.1�������u��qZo�P*�̕SF=�'&=	��Y��w����"�����]99j�\f��_�֥�P�T�i�l�ڎyFj����Δ��_%�ݶ�W���8',Ƶi���X+�����K���s�^4���Ƿ�+�9�H:�֚y��$Hy�P0e�/��T+KM�^$O�\	��+���d�K�s&s}~��^Ł^����p������5����t���E�Z:S_��>~C�)ZX�����
�}����)�;[��C�m��^ˎ��޾Q�[u�,�=�Pʀg�T�|�Ӑ����r��W1?=�k�'
/E`j�w�c���P�XN��6�f�r�;�]r�-�y�	��Z�	ffVZ�85.ooA��X밞nr[���%;�f����9r��V4�����a�9ҵ2P�/8��֬(�֫�2t�vQ��1ugV���]��YX��zZ�E.�7�=���3�+9��z��҇�Z�_��!�N���iek�'�CR�>�u~�y�v%F�x8���1sՃޫ���1����l{�D��q�,�2�6���枚�R��]���&ˋ���dw��K�b��&��a��53����ӗ�"��r}�f�ל�{(�@�3x\I�&��n(��k�q7ݡi�x�/�a�􍧫2^�c���k}�`��/H�G��M�:6��]D�!���xN�
ӝ��Կ[f/E�޿3�����*�"�ˆ�`�@͇UL)�$��L�v�����O���[�]�4�~�rr�"��+c�{ʏ���3��~���~��u5�7�Hj��>�Q�~�)��1n��A�/-�����3�\��������@~���/e����s�1�6Z� ���=���w���{F����m�ѿ�σ��z�`sCo�p;cׅ{
�7]�ܗ��Y*K tI��6*q���|�����
/�.}��h���@zO��:1�G�r?/uY6:�G��=�.���'�7�b�m�/9{}�V�O��9�%��?tp�i������^�9�����R���4��o��6_jT�R�:`���S5�T�_�ݠ�>6�p'�*ǣ�R��z��|��]X����R��	ɤd�����r��[����?��I�>�0�j�7<|\�D#�O1�t����ODk��&.5�d�/q�ty!7�?4�O\~�P_�L\w�#Q?����_�N%?��,��=5xK]�FH�N4{��N�|��������봥�p��+�O	���^OkW�ɖ�{?e��>�Kޮq;@��M{ c��=�M���l�q�}t�E�%P0�����'�j�.�e���_����� y\mC
���:^��߫��"�hG_������%��k�y���]eVV��pE���x����z'xV�P���n�Ρ�6��J�:�op�l���%l�H'�=�N�ӗO4�=μ��W�_�񺜟3�<��=;���&��T������#����\>�>�����̀�A�`q�/�1��`��2�ӊ��9���*�U{yﭣ��U�?U3����p@L�[ WǥyM�b�]�`
�ﴏz4�>^V�\�hdAy�c������z��]�J�g~D@j���""��.�͉�+�hd�תA��+ɃW��#Y�4�,�̙��>�J���{\X%r�>��ۨ�{�a14��ѹ��l�.[�7�[�e:&_f��}3��Õe���;����4�3�y_��J�a��M�z�+�>�K��ۘ���Yٖ�C����.��Π1���;ߠL>���!���0�{��3��oޮ�W�.d����\v�g�
H��',���Ou*2���~5q�w�j�E�ҁ���|`/H�EPWn����6���Q���X�b�O;4�b����4�5����z��d���]�cY{fYc ۙ]�j1}榄����8n|����Â�z�+Kñ����������Z��um�(e{Dz#�p��ǢNo�)�֦�(|@�{j'O�x.qc:�{m�d����>�ا�.�y���*k#>��7��i����+���U���yP�����y�	��،U��kq5X������=9�]vӛ���h-ϻ��4<�G���n��~�����\]=�ZS���n�Jp,1���V*�j19�1Ϫ+�\��A�s������	v�t�E��ܔg�y�K�*����������ΰ+y�g%�6{�Ņ��_��S��|�J�U��/vx^�]E�!S,('�ʙ򘿢��p߰�����W7a�zoif]��QY>o�S�w�+�H�p9��n���N����z,�;S�كC�1�j3����I:� ��-���_���嚎�9Q�[3��[��\[���ɘ�*�A����,�ԙ�4+�Y��p���Ve�٪5m�X�M��=jA�4b�ϼ:�Q�*��ǜ�2�DZ�
���@�,IR��_x�'3x��߰ս��F��O��Nnr5ǩ���Qg��ǻ>.�C�9EG��fL��7�ޒ��=�܆]�@�����.%�^�3�u�2�=H6�N���#+���sɄ7=s��9����s9.2 ��G�EZj/�뉹mb�_�5���Br�UzR�N������0m�������
 6�T��V|&�]P���r�8�wӵ����+|�B����U��_��ꭚ��TK
I����:`zxM}R��n|�\j������n��vi}B��0�M����@~��n}E)������Vy��sL�#��H�sF�n�z=
�+�7���\/?Y���s��"Ts�Ш��}'hB>ܬ��^�XD_��V�G$
��(�1w��!�wt.1��&�.gj�
���Ts�uDяo�jTvǯ��U���� �k��lR��j���Qq���~֥�_<U>Zm��k�Q�ߢ1�P`Xg��� 3��4��`ǧH�o�z,�';qq�@sJQ�d���2�G��.<���u��P,�ҷ팼��̭���Z:�X����M�ю��5�l�j�j�1A��+:��-Y�@����c�β��v�<�y2f↞�F9kn��g�mL��ivkk8%�U\�V�[�M��.]��Aoi�2�J�G��\�[�1,�%�qO���F��,XN�5�sםc���+9�(S��YZ�)@L�x��Ģ��|�ٰ���Vmx6�V�uG���D�R�/h�L/��U;����N���ᝊI��J4`��{��i�s�g�-`V�s0�5��7��ggX���֖n�S	B����]�r�����'�ҵ4�'|i��n�-�����N�Ԋع^r'j�ƶa�u��֢8�7A��mg ��-R��>��2���''�Gv�\ʔ�+���Y�q��Z��2�9��fN�˫	u�a�������s18������J��K�Z�f��v����9*᪎�]��j�uζ�ĸfՋ��8�ܭR����	��N�H�� ��-�f�v>��!�3O.B��[�w"no]l{�<1,9�Ct�2�u�Ŷ��N��V�ϊ��q�=�P�{L�N�n�}��Rw�&�fsO��7M�؏*Uۖ ��W^�]I�>���5ۦ���a8���J�ilN�|��\���G5{[A7Ian�Z��R�c{\+"�wq��j�0��&oZ�9(���F�d�8�vv�JP�?l����h���~F��s�h�T���~I����r���L�Y�B��i�1u�I=[��_]���JJ�l޽��tCżl%��7>�%�TXk(}���+T���uЖ6�^4B�����Z�:�;r�|���Aɼ-jy��@���K��6��N��R=��b�ˡ�����M�l�1+����y�v�N���������[|o�X��s�k�
���u���Sg�s� r��7�7X4�<���2�&2	���lm��t��ޱ���'m�F�Z�{�v�=t.�Zg��8�N�����l��;��&ʇ�ɕ���}BVV��ҥ����ΰ�\vA��)���������E'ZE�i��_[=�-�e.�VwBh�7ˠ:3���8�+�G��/�_gv�u�H���h�W�Wu��5��;�Z�|�Y�:�&���|�fv���6�ZV�;E����O/�:���n�V�����o�ՇΘs�e��;�G�a�n�F�i��t�ʙT�vӭ�y�h@ib��+�����+�M��LW���w�i�$�=�E��Vޡ+3�<���<5�����B�7`�����}cz�ki�{j�qU&.[;5�U��Nܭ��\��1ƚ�����WeoP$�5ge�}����)G8%�n3Y6']�s��d�L���TYZZ4����C(o����d��rB���6E|s�L@rn�o�.c���Y}T/��gqd+��\���D�$&-S��)����li"��4c%�m�;�˗3"�U˗(��ˮ�,"���]1��Pk.vB�ܢM\��;�Ys���9��,A�C"���Q�+�h���F���@Y$����DP��r�����4Zd�ͺuq\�3&Sr�(���Q�sW7*$�Rs�!� nW��E�"�Z!�B�@1P��!���C`�2H��m�Q#)76�"����h��4r�d�wuA����3EH}Dw2o�bV�����թ�[5��M'�}��\��ڽ�.S]�c�e�\9�}���k�����,o.ɏ�w�ﲋ�wgi�� ���rA��Jӕ;�E�aF]mt�%�����b�NO{��I���l�E���Kn�!�郇�·u�\n(�*#�1}�y��9[ �i�YQ����O#}����j�61��vm�Pѷ�E���}GE�S��7��}Zm��	k�G1z�.����02=^�x��+�qݞ�����Z6���PM��tB���V����;#;=��n���҃3�E{�C�Ɨpb~�	������!��.��y�Ⱥ<I���>�lgs7��c|��>�=��h���w�!�άv��������1�*^R>�Y��C�r�^����'��@���wFy���ax�[�������3�[�����GN���3:'ѰO�s	^��zjO1L	��H�<W�Z��In���<W�c='E�s��T�i7R3���n=��|o�"�d��
�{Ǆ�Zo�:���so��cg(��T�{�����ӺM�z��Ǯ�ƅ���n!� t��x��o���!C�ce~���Q�Ezٺ7^��V�|��fnk�Z�z�����t۾
x�=���c:)zk����~u�,����3pG�]��g8ëդ��k�ws� ڵR���3��b�%�s8Ʈ}M��Q�}��T�7
�ڨ�7�R��\v/zzC����C~������L�&��ꍁP�~���S^�q
d�����e�������j��!�*��gr3��{�)��k�w���(���p<i4�Ov7'|�)"��w�=C��XpN�0�xe^�=5��2uto�>�x>�de��D���P���e
��zV9��a#g��"�n�O��xV�ˇ�z�����_�[�Z�d5ބ����^N��sS��F�28M�OdN�ro� ��;�ڦ�5�u�{_��^��x�q��.����t��Ɠ����)Q��H�zO������#����/�q�,K��^ˇ����= y��B�����G��c{!�v��y��[g@ݸ=�u/}y 9��Ѻ��+��}��)΂�i�?bv����"W�����BG!{��>�F���֗x��r}3�>������˅a�>P�����Ϻ�+�Q]\�/zko����CGg�}lK��{��3�����juT�-N����-zc�g���\Γ�4���}�����S^���_,��
��x/9�hICOc���Vp�l�Xq����2>�m�ޤx��|U�:�%48������Ե�	19�n[*�����`�V0��p���{����*����;0'K��vn�r�����¢��n�æ�������뾧��7ݖeE[�~���q�WI�	+�x	U��{�W�5��Fy��wC,t�u;M9�~�րcF`qdpچ�P�|i��'Af�jH.��(��\T�^�[m��������B[|�T�W��}�ll�y�p�fpuE��^uLC��E��� N�������x�3�>W��U��e�z����.[V�w�CTC�n�V�@�P�P��,lxLK����S��5�[��grO���5�A/ż�L>���!����ew���ti7ޮ��_�[��i����L����`����d�!9Td>9�&�}��C������Hw�ː�F�uDM�n2���o\��r��v��UX�b�L�)��b����R|�Q�����CmUQ���yj�5Is�9Hy���3���֦��5-q��8*\�:2��E\l�.tx�k�G�W��6FUz55UF=��S�q����)�֦�ʇ��pǶ�qd����D_W��`�k�Bh�~�9�>[�x���5,�������-���l�k+�>��*մ��E>�
��5�x�[��l���B��[��r�U�d�9W�[һN�Z���V�un,N>og0�̏l
�)�����A�m��R	zz�T�WΤ�.]v���d�7n�(���ӡ�n�m���[xڷ�p/m.�yڥI^)�D+^�7�.�D�E\;B�>�a�)RF�΃����Q���}�z�G�^��eK<^�߼�)N{</qX5*��;��h�\��f;AݨwYK|�`vL�}|��ߒ\���s���pW�{i#�uI?Y�l[oQ�`��x�[k@��&�/��I��Ϣ_��C�29z���͗+�����ȭ���9Ug!��fG��߾�z�{!���󝢂��(��e��3��>S�9M�i�+c ]Gy	��f%/��^����*�D6[i�C�Y>�X��$r��s�L���R����%;��}��=
%:�/�eO�ht���5��������FIE�(��� ���]!�.�����"��pI/O�*g�z��:%�^��<�����z�=H7��������Pglf-<���ўٰ�'-�1�'��L���3qS0��W{�[V�w>㾇�x�{�F��@����3Z6�5��*�Er��� s�#����� L>5��~�˃��-���2�.yݏl�'{5:�[>@���G_��٢�IcaT�����HU�T�>����Q�}������+�{��[�g��#Sx��b�㸕
m�鵙��jٳ����a��"j�p��J_i���]'HF��yh�mM��WYV��:�FW	"�^�&�P0����t/:.���7�I�MVw9�aJ]vL��>V0ZS�^[���7��#H��@���8��d߀�ĵ�+�5L)��I�_)��V=�Ci��M��������^�k�
+��G�ʤ+�5wF-��>9�@�`u�,�K�^���.�=�3�3��y�jv<�o�Q������k�����~��}���
�p�;ѕz��R�=��\Z�五�}$�C�@��-Y���������{�W��,*��î��zhs��g�G�.s�w��0\��kRDܾva�+O|��<��e�[
���!�P���{�MT��>ˣ{��@N���*��;X�_520eD��X=��}L��pʬ>��~�^1���e|��v���]�[b�ψ��n�����k��#�m�6��6�'O��2O��:��|�\`Em%sw��>3/�yp}.�0ν~�[^ˎ��޾F7�j�_E�%+2�P3Ņ������n=h���{�!�l�kC�c^�
߽����C֣݅�>�G>��+����ި��O��{V�T���+�	M/i���Ƈq���f������?]��9/)Q�{+�����δjjfhAE��w���Q�{a��m� l�X����أ�����4�y*���\y��_��ʽw��[w�]�9X	k1�YEqU�����j*U��l�t�mS����u�,� g*�R�X8Hܧ;&wGM4Us���\1a�ٜX+y����G�g��%���0R��і��S>	��U_u6-��o���+&i�J��!6�;s������}����:K�r Nk�<�J��Kf⌢�r>���n[��t�ʪ�Lk�Ԃ�m�W@�p�?H����#n=ul�������:�/J��;Y��F���Tq漰\�W����0�->�������_��ƅ���n� t�+�4KUL�D�V{����e�>
�1���~�p}�g��7�*<�F��5N�W�M
���n+ �j|s_�;i��.�|{{���^ɭ��_jW!��׮��z�>ϣ�|�<��sΝ���1��^#������nj@�8�@�
�m(_A��@�b՘���e0�uto�j��{��8��q��
�ƚ��:�; ��]@�z�ԼǑ�n]B�+�C���gU�{����ɭ�x�_^��챻���3�6�L��Fo5��j��8M�OgӇ'�&�p�`2#0z��܅�I��Q��lqBi'��|"�\���''�~Fw���	���da�?Od���B7�l�_�-�S�_;3�{�ҫ݇~��nLn�)J��j@�%%o�7�p�I>���{:�n�:�l���%v��mGU��E�we�G�k�Ko{���\[�{'S��K���^�:b���8�*�@�өڸqq��K��%��wu����g-��O����zx��tB�}�q�_1�3^���y��60̀a�	�b����Ay����J�K��ub����U�쁎���o��hH���H^���&��H���j�cC���Ԗ.�k�cp��v��*�n"��������������W¢�(roTe_s��Iؒ�y���<�D�k�>F��T;�3�d8	����Z�h�}���u��R�t�=�{$�.7��OW�l����j�KϮP$���G�C��Jb���&r*y?���~�[��+�+r�fL�����}�'����Ig��G�Au�>�3��mI��g��
P5 ����}-z3��+�X�[� ���}��։�����瞧���iY�Ps���c��3��	ў�����^.���(ז�<z}ޚ�ê1;� ����;_����=냧�N������({�c�?-������<}�A/K�}ы�C�����]������W�[2����^�{�8��zUQ��D�@r�J��|wpL?šG���Я6�C�	q�#R���`c�Eɷ�n�t�׋�q�V������#�`Zv�e	cU�F��6�
�	�L}���S~Kt{��R�'Z=]ُ�Ĩ�x{������8/Z��k!��l�O:F�9�z�c�j�;��^a���F^��HM���d�fٲd6�G����Q]c�/�`�L�U����${�5*�9U�/�!X=�Fk
<�����2,�Y]��6f����� K���9�z��_/VR����+�ӂ���;�~�z��~����&���J�D>[�}�)��o���ы��%���G�c&�b��r$�a�n|1��9?o����-���)8�~�8=���3�.�xg�����y�d�<5൵�b��5E�OT���Q5��ʙ��@���i�s����ǅF���������.;�CǍ�Փ�z�b�S��k~��E���|�ۢ���sz;og�ҫ�
�y_�|�x��u��H�Ջ���7�Yҧ������������z�N�0�U���W�7E��7��U���Z���^Z\��e�#�.�#��Tf�{݌_��]E
�Q]���y�Tϔ��9Mr��gbܵz�g����m�>����п��c��:�p�l�Aap�P
,������){Us��=�Q���^*_�������N\=C�|������v�,"K��h�6Yʏ'(G�1�\\�?Cס���TW��l�,�����9"����r?Hj27��l ���A�-�f.���a����guw!�:`��.���=Jr�����vGM��GI��)�	�$����ĳ9jy�%��d෣��H�ۗ�ݔM�s/��@��s��޼�5߯F}�'��o�3��@���Ǫ�a���=y��+2}6}�x�΀����u3L��Q=��0��#������/���>�����Ez=wz*��K�� '$6[������b�e��:�	#��#%w\���*���ȳ���<�du���h��X�U%��$�ԅ]K��<����F���
����=	��W�����d߀��V��5�Ca�W��B�!�V*\��
��Β|�,�,��n�fݠ�^���ϭ�wF/�߬���@�/���~�D��!\L>7�>7��*�$��z'��v�3۵�-/���3��s�rJk��%�\λ�T,�-D�O�=HЖў0����o}��(��q4c�(F�/,�H<�����ylr�����<�
�J��3��2�y�c����)(ʑ^�@�߬+�o+ҵo��04�~M}k�OD����x::0vn{��Bm�ގ�;'^=���;X�_520e@|'��\n(�����A�󹽼,7��]/�+H�z����.�e��V&�Q�����ci��k�nd��u��V�ŉV�	���ր`ʸ�����]M}�~�.n!i�cw:�"U��i)�|MN����m�^R�`sV��*���y�w��_Gr�� �!�P�uqUZ^tp"ms�m���-��m(��,c�1��vm�CF�.r4��ܜ��6ݷ��b�z�>��<�&��������u��Ͻ��c|��p��b���5�U�x���6'L���l�j���15���{+�++ԇ�9�c��}r�f�^|=x��0a�u��\Q~ s�b� Zs_"_�H	�Ԅ���_�������]��>���@��Y�u1ΥoG�> �P^ڔnD�Fc�����.|9꠯�����㹞-����X[6C�/��n`xg�{�LvO��=��/�����BS�z[7FQ~9m������
s����4Rw��8�p�fpmC�Fr�ղ�ztO�Âu t�n�P<�(U{��[̫�è{�F���s���^�����;�[jk����|3�Hj���4���Ǖo��&t��Ě�v�WO#� ���]r��a����ώzg7޸��z��n��+�Zlg!Xk��Z$������y4*�k��r�IԄ��-3,��F�����>����Z����kkZ�ᵵ�m��ֵ�����km�]��km��m�km�[Z����km��m�km���ֵ����ֵ��[kZ�um�km�mmk[o�mmk[o���ֶ����ֶ����ֶ�񵵭m�絵�m�v������(+$�k:M�#��+0
 ��d��I|w�U@PR�(��(�TED�I%U*�$(�+�T�*���J���@QJJ�$�UJ*�(JQJ*��UTJ��_X��e*TK����dK�b�TZ�[2�ɶ�h�V�:=kұR���1(��A%l�e����%)*@�J6dø:�;bfh�ZR����R*��Y5�)P��j�Zh�"h�	B�	m�f�Y�:d�D�h�*���@T(�J%m�e-�iU�[� �>����T���jۼ�p�Wo{ǰ�A�ކv�=�j���1봣����Q�{���y�ު��X�^b�xx�ƀ�s��UM^��J
TT�X1o�  �y��}�uw��Ӵ�a;����:O�Gۯ;� �F�:�|<Q�P ���Ǣ�(�(�����@Q�F�=������@<�x ���^[�G�@6v��z�%c�p�E�"ɓ�  ����Z�[ޯxh���m����z=�׼Z�wT����G��������{��O6��U��n�q��7�Z��^�U��Wc��^.���U�s���^�iF��h$j�   �쯵���+ە]���]�ӽ�\�����U�tu����ve���uwomƮx�u�@�g���x�Ovu��ov޹^����{m�G�n���uU��Û��C�k9ꠢ�/`�T)@a   ���3�ݽ����r������kj��랕��CW�kջ���ޮ��k���l�=�%��݂��׽��n������٧�Zz�vq��]�]=]�C�Ukۺ�u�h��%E�-1#]nh��P��   ^W�O���w-{k����7�εͧ�����{����j����^���월V�uݯ%]w����m�������׽ԍ^ɽگ����Ƿ�!��e�Z�{��kU�\�)PU=j4¶�UF�   ���������z���Ӡ���=w��ގ�6�j�w����W{=�5����)�'\�z�U
���z��w]�[����W����Uy׍ޜ�n��5�y^�{W��wo6�5U�B(���5��  xWٷ�뷆�����2C]]]i뽴��6��M=��ט3�۷F���׻3�z׫���u��vw{�Ӯ��yѯw�j��v�y���T���F{ez=:s(�4��[j(��h��  ﭼ���N�{�[��w=��6�k��M���^�������V�Y�Z��S���OSvV�{�u�{�M;�O:��:�m���nj�y�]y6��n�*o4��Δ�귳�%RB�u��v�v5B��/|  w��ݞoS��{��Ӫ�g�:�����j�u{�����8��l��\v���ݽ��i9$����y��ީ׻�֏z�޽-U���j����| �?!3*� � Oh�JR��  E=6#*���d�JUC@` T��钪  ���1�R  '���/��e�� ���o컗���,[^��}~������Z׿xy��AQw��AQt� (��AQ�D��* �" (����l~�����F���N��aՁղe &�[2m�6��Eݵ��n�k��@�+#��[t�#��7���:,���-@-� �v��&�p�5&�����&ڻl@%X�"��F骽wul�6S�t�Z��&R���+`��F��.�Kb=�.5{��^J��2lt�]!�l���J�s��+L45�n^�9je�{B�[B�>���d�X���,�e-h6 ͌��<���1!?�AWv�"��+�Pw�N�{�\Je��ʛ���X� �.� �m*�y+,���o+wn��)<���qh����q�.X�k�Pǹ���X��!��%K�lfݱ�����lG7h��J1mGa�%�n���(��b�M�4����b%ڕj]�gqH�ATU۽���G�i�jB�V��uaf�i�(,��Scc���*gu�91����2�</34�%!�e&h���p���(З�ȱY¬�W&�9&��I+r� �ȁ��U	�0T{y�DbZ��4
������`[���p&�8�l��]�3(�؂{��V=pDr���~7�
 �%�q�F�n�)�&�5��mj�(:�7jhX�Wm-Z(Pt.�K��c�hR��d?��C���h��B��|�ef�%���d�y�e*������	�{��zn�,i�p���z
�%��``��V��Y#%������q��od�����6ވ���xd�U���t�V��T�c�:#Z�3���5�ҍ�`h�hRp�݀��[�ku���a[+u�r���cK�6<�/\e]�)v��3즢�)����^�IA6Т��7"��ˎ��8cX���,n�XJ$й-w�OJy���,@.h�i��mܖ�7	6$b�h:���/S��mˤͮ��#Eۄ\��2�W~Շ-6���O%����!C��m��2�fiH��j�=ń݁�S�T.�3`���jX�[�?+�aj �%�+���l]����r���ܛ���z���ۆ�퉦�5�-y6�L�R��Ӻ%�$�-�ýwg.eX�m���dm)���+�2��Ց2�Z�7�ؠ��וg1��I�r�V4s-PQ��S׷�'ڭIc��!V����[����(R
ݵK͆��
��Z�9
�Nkq���N[�څ	���Ma�+F|)��oPcqᵒ�,Qn�[����Pr����ٳ5�r�T��ChE�v0,�Qu=����R�2��3JOPl���6�)pd�E�A��k����6��(Q�b�O�Y[��r��E�I=��f:S\����m�N��&�Ҩ��u�$�����y�n�?Z� �
(\J]L����%-�v�?,�.r�B�B�neۤK�f��I �u,�O�Lgt�ݸb����ۦ/&��
kᔯn=�tEcX
��W#x+j�!�L��)7��Z"�RbvV��g�q%lIJ�`A\wJ��ER���MQ.�pH��1H��kE���ړ6�P��q�oc��G��bq�.��9dY�)��[.fG0D��l���{)dϞ�Bƕq�/(�fʖ���*<�H-WA����˳�m̍����M�BN+Ϟ�H���E�L��N�ъ����EJUɲ���t�L�J(,��#�̤�>���J��ɛf^ܗzE*ٸC��v-7n�ט��@:���u$-���2v��ݫ�݅���N�aV���X���Q7��ɹ�J^���35*�:Q��R�͵[$�;�����6�廃!��F��؎�E8#֕��I��k*�;eȚ�S�^h���͛a��S$h�L	REX�l�-�:��v�� �F藦���5JJFn�J��E�v2�[�]Ѥ���P��&���/]X����Se$~X�JZ�c�zUǑӫ�*�7P7q52�׫&�j�»�f��m�W�'�k���w,U�����`ɛ ulA8eC���2<��V�4q=wd\r��.ԭ�Ҋ��y-�z��#���[lfnRx�U�t��̫l���7.Z4u��<$nJ��A+�WJ[��M�k�l,0�ӵh���Ҽ�7�]�)W���r��xʷ4��yw����)�Sܦ,�[-�Kj���sL)�\�j�u��9�f���	v�a��n�,@�YXةeM�<a��D#t�mef�]�qݗ$����D,{�42��՛��gwi���8��P���]Ȧ܂�ш 0��`�2��M%R��Z�P;�9-�Z��H�WwX�9VFM��&���6�梳K�u!v	af{;6��6�ޱ�/emɡ�c�L�R�C7�����ך�#< �7qTXt`r����^�̐��b)�;��6�X�a:���H^}1he	t�+74Sw��M��O�g��m
u{��w2�e5��q����mJ�B`�n=7D����:@��,S�sm�6��c�)�)��ۻÈ���j��*ӽc[Z�ږ�;�$��MnЀn�3.�f �WVi\����]e�sZ�R҅Kt�Y��͙.�GCi`:5˄��I�Z`�zuc��dz�8n0���ƽ�a7H�25���4mc�9y4[�ni�eYn�	�,RV�۲���P��duh�h��@Ik��9FQۻց�jz%"i�ko-�A�wz��B2I��qQ�Y��S�Q��Z��!�4���Nⷧشn$[�b�Uu0bue��=te�ҕ�����S�U�}vj��WW���1+�G
�i��p�UI[�]����JV˖VLM����jRl(hv���f7P*��0��b�o�`z�at�w�ʹC����QW!��Q�h
�2���1�Z�L���T@���:�Q����Xe�i#�-4(��w��
G4`����D]m*X���I�r5��5���/v��n��V�(�EG(ӚZͷ,2�Y˙6��N'/�Yz1]m���DN��&0�޹�˷�
�EJaP����b�U�Eܬh	/`n���7u(�M�Vj��V�P�D-�nQ�\�ʔ4È��!�5�$�(L��Ȱ۽m�?rTuv8�*��P�2I����^K:@'%��fd!�M�B̵��*���dT�X&Tl����l%.���M֓��d6�����Sl��q�P���d/(��-D��V�I[�0M�z)K���.	�wX
��	=ɲ�eE��Q�w3!T���u��ؙvUIMlx�4��.ƨ�?��9��֤(5�5\لAyY����N�e]KtP%U�
��v-a^Q������e�U�O�nn��N��MheʥWBbN���.X���"K�n��I�)�v� ��㛸�y�kٔ��2��J8�SZ��R�SDK/kR���B��b�(�%��J�v�Z�h�A��7#ɡj"��͛�ɒ���b��&fP�m�T��ޥ,�c,!�cZ�����])oq�N�fZZ�4I�.���nc�Ce!%�[�mnޭa9��D���7V+[������CZ���v�Q'oGm�C�����N�̽��:n���d�񺽧A�j�����H���t݇o[�ˤ�Ŭ�P͘�YQ�(V���=��V�2���]5��&��6���mLv���谖�+�5'��)U��!8THֺ՗6��Z���������5񗎶9yn�wcD'1D��6��n5F�ugj�fb�C+>�"f<�]�t�u�AM�WXv�3b���&,��9+�Yo)�Tֱ0���p1�(NA�)2�d�&�ʅ7��h��[C,�=:�܏&T�e��X���l�2_��:ճiK�eбq�י3����1���v�g\Ս2��H����sV�O�}�(Y�K@�8�W�bV Q�Z�A�]��e�Щ�T�IQ3�e��O�1��s)V�3CyY�;�L˳)��,�i��NE��C�S��DT��cE��jL�w�!Ki%�n3W�� L�4]�M=��j�NCt�s4:հ�(����2F��K@�m޳�'
B�.aek{�Ɲ�D���w%�n�W`i�J+�m��#Vm-(V�CDM9-ϝG3uD��.8�.Pd܈�0�A����
{��S)��!P�p&�Pnl�IXc�z�{K��h!��3h�r�b��ɵ��<1fVi5���f҆@�l7�	i�rH�Xpk��f��r��A��%����;�ૉ��w��U��c*�w��a5���d�3o
%���x�9O�kU�wg!&]1��'��[n�݋�����1�0P6�࠯f��*�*ul_��ܬѕ)J�-CEkN�Ne9�)̫��IZM��8�n�xe�*m�)
��a�@a�SQ��+ +qї�O��p	��$!�ү�x���օ/ok
Eb"&9� ���	 `d@�0˦)e�i8�FT�:�Q�Ӹ0b�EHb4vV=+L�OU��2���#sd�v�� ��T���`yG�"��2u������ycEY��1�U��KF�ui���x�m2��4Uּ�f̊�������vV�5��Ӂ�5U�W7*V*U3XՂ3!W�i8M�n���ֶ�ɬA�u5�_]`��Hp����jn��A$�)}o*���2<����N��턔s%Z��FcUګ��N�,;Wi�l�
j���	2�>?G�wb����*�����,�ll�V�v�����)p-��.���`:�50��.�R�e^U�@�K6P��0�m�O�W�Sy�jeX��sfr[���>ݔ;��� /
J��ʋB���L� ��(��@HX�Y�\�.+W
36�*��b����[��w�h�ʰ��V	��I`31*X��8�uWť��Ut��y��,�0d��j7��9��蝀��EGd��ٵz���P�^T�e� 5�fi��ڒ�RxS^8�/d4Y[��d�OJ��'VP�j��j�Z��ˊ��l=�[u+/���;BS��Bq\OB��^G�6����· ��xh�]�b
��R���jP*�4P�*�;77L�"�y�Ku���̋X.�fP���c�Ӎ�(c���X�b�5�T̚p�@A�3G��X0vY1
��Stϓ�cnI{ v㕮-��%^=����he��A�p� R=ө���A�t^����;4��hT��X�H��c^+h�9h�u��(�ʐ5�,��q҇1�"���%��!��������j���oN[۳1�S�T�����0�C3PɣH�t�fJv���T¯	�N,�ͧc]�J\�Q�!�N��M��}C(އ���t���L:0�%HnE��Rm�x�����fa���jŝB�q�Ye� �gZ��j�W�0Qi<
�$C�["�;�� �Ǻ喥�DI�	��I-f½����k�����v����DQ��5���~b�Z-Gf3��35���J�uY�!����pU��z��4�k�(e<�U��Z����t��E�#8#���R��ނS�l��Cv�*�]�Ʃ	a&�4 ��Y�J�U�*��L������Z�.��Ҡ����B�U��nh �p�DbƝM�.�K:@�)ť��q�[xbXi��&
���!��V���¡sL��e����E��ցm��gr�P� ��>�ǈ�͐oQ��nш��%l5{HT�NXv� "���T�۹�����2�	���8u�B���*
���U��	��r氡��;z�4$���Dn���:x���͙{�x/i`w7�9sh��w&j�0"��1�C]�W	eŐ����T�q��=5f%(ԓ)��6���W�ܬF�o�Վ=���a�769-J2�B�֚6.�zF�l�347R��V��H���eḰ��ur��V����:�v|J����Xl̙N�e3${WQ�tN�J7�eTY2]���j&E%��+B��;!v��@�Wy�d�"��vf8"t"`�,�m��ʧ�Z�c%��n�"�������]�i�vșvN�ռWQ)��FDE8,+��Ef�(�ҁ��嵰���Dͭ�{�aB@̀�I���tt�XrK�����<�N�D��U�囕����Oq�M�O`-l��)���vV����*+6m(��1�Nd�tƊ��{s)]�4���mJ6�]Y��ݠ��`&i��3C��V�l`��wT�\X�<O4mf[҅MV����5ʈ�v����BḺ��J_�V�n&jP �X�"i�4El%l�sB2v��^Z-��U�SLi�d�i�nJw*":CY��]�Z�<��.%tS�D8�d\��5Z��p���Q�TX����tB���bH�e@r]^ItK�@���j�oN�Nd���{eJ�����cm͸RWg^���#u���ueaٶ����l��B�»vt@���kBd����f��TE[�u�4�X�iĲr��.�%�\чX����e���X���2��H�ޘ�&�*�ˬ&��"��d�-8�֝��'�5�[�&cѴY�n;��kzҳN�aܿ��u�qӣm�2�u
j�J��7�� 
�q�n���0�7�Uf�����4b�"��Ї�6L��a)i���J�VbSF:f���Qz�٣2PsFs+B�m�N�!R�^]��X��c��+#�CE�6)GJ�B�)#�/%꧘�0$-j�5T)���Gv�խ�u�����C��9RȲ:��UM�`S���F���|�VGI,��X�ThM_=SD6���p�J��E�bV+n
h��IX�	��2ۃV&�u�l�G��9��t���E:cE.�F�k����8Z���[�M�1,�-�g�-���jAЙQeY��N������n�82�U�g�SB��b�5��:	��
��I�-��"�]2�O��J�]Jg�Z��,M�UT�6����'E^{�Ap8�]3�]p����2b�"�t�e�6�7�{M`�R�e�����E42��{�3.�s\������x-�2���7�]b�44a�r�e⮮���j���,+rԤ�Q�.M�ӑ���0�i�mԼ��L9wܫ]c麱�K�>�ZB�\��`j�UM��RŽ�n�p����{��Zj�˙H�+�RX�<V��w�S*��Z[�=��iIN�U��<�\b�6z�,�w�ɗWѧT7kh�Ή��D2,Z���I[�z�'�|�[Ӣ�W&m�|,�V�!NV��h�Z�Ou�__Ԫ�+�0N�:{C��x��+	�W�6��1�;nQ/�a��V���I�̜6S� �����4􊈞�(�.5��ٚj�;�d��g�de�lk��r�Hn���7�p����&1�S9}Ks��pǲ�	��l������e䳴b�16=:FޢJ�5ɣ�a���zEYc1����>X��	5Pcf=cf���P��8�`T�`�j��7A�{O���/c��3x/qޕ��0L���kOW�_j�M��%Z��s����:ݙN鹻�O�� ��k�W�hG.��W(YW�(vqU9u���/1ɣ���pl�A���a�7�r�U��B�c
됛��`8������M��T�*�!��2ِXׅ�����uSF�8*�:�T�]����-��8!���F���wNt����Fqm)�nͬ�u!��
c��7����hM|��Ό"�|�����WQVɆ>bw�6�/���.�Ǵ����(�������N���g�jp�p�$.δb�����D:UyG��PS�u����4�t.�cXj3�>�.GE_�d� �Q���X�V=5p�9Ν��)K����ۼ�tunNKYc.�ky��-e�c�}v���ci1U�c�pV��rgK����a�t�e��u��eD�o�h�Vrfu���.*���v��q�b>��v�9�T���[6�a���=z/N���٣�Ʋ[��-��r��II���m�"�4���/DC��u�U��%NI�ۋk��T{�ʱ��6�,��-#h:ꅞ$�b�ҵu����_.�Rnmx�M��oh+-��S�8�5@A^��2��V<�5h�vc�Fخ�ژ-���&PR��Sg�����`뚞���!�����)[ݼ𦻺��\�t��vŧ(q�b8w;�a�41c�l��h����b)��l��w�y��o'!WE����sy��ȊF����V�f�^հZre�k�G���DlL���2p:�N�	��z�
�ʺL퇌ͩ%�Oat����W[�};{�ؒ�E8���D�#�1�[Vޘ�ec9m2	�����<"�cͨ�:%`������c��:o4�Z]���#R��N��	^�N+a�>�o=�jD3֢����)Y@fa�0�we���w�z���t�����돗+L�gi�P�]e��Ѧ���.�jk*)ʹn��e�x��E�X�=0^Tz��aO��k,]�N��
ẜp92�|��3gc�X���1Z���$JZ�mg1�fBDJ�#��+��Xz� N�9vN;�.+�E;W�L��A�:Z��F͌�٘�v���t�:�":�M��h���l,ӻh��?���%.���֔��J�����̦���F����"��֤��4m��iH6!6nr�n�*(��L��*��[�3j�2@�����*��IW���j7e��)��
�E�7n�.Vƻ	Wb��Lͨv-u�wK�	�x�:p9PС,v;}]��������T~���5�n.`�;��Qޙ�x
��6��GٷW�v#�5	�����Ŋ�$L�T�n��9fubw4�l�/_h�-L�[[�T��\�ʺ��
�W{�ȔN����� ^m�y�WK�
�E�5�2���ȧ\-�%(�����.%6�B�d��M)hu�i�t�)c��+6ItnK���*�4e�!^9#b�ʚ}%8]#ꡗ�s"d�q����,k��5�KAd��j#n�`�P��mt���@���Ҙ�^m�7�sUeh�:�$�vT���ށ���[@�Ш[��}��
�a�ȞV	@.��d�x�gt�d���'O/�/��X�@�
��u�R��Z��z�^������S�oP�lh 뎐�t��^�g���h늻 Dm)J�{rr؞��YG�
�{��Z��g6��5�-�3�1Cz����a�x�Y�(;	�2��6�wVsY
�~%�-��h�D�8GA��\�:��ls�. i<:�OE��M�lu.��[�j�6�-Z�����u�*���4p"�3�U]��';~�1U����G,-�|��Ť�Z
�FQ%V�n��>�c���vM����*�e�A�D�,�v��{M�(�!]e��s��^���+�~��ͧ����X�����Y�gZ��8�o3��q��hEh2��ٗ����2����;�:+_2��:��SY�X�1m����L�׼q��7��ޫˊn��S�HíM���D�]mA�'�܊`N��`����{&�8��*:��wE\����H�ڌ�̓�O����sh�9h[��^*�"7-ଽ�u��4�;���G3�2ZTOe��X�:�ж5,:)d�herx��t=I��T_4�Nل�X�z)ռܾHPdVG]�H<���&E.�c��i���W�;,pv��F�Uκ']��*҄.��^�W]���J��ܺ�M�Ε��i $�Fk[���8J@��������MBCg/G^�E���՘r����=-����ԸeD� �f��u���b۔�5N��T�K �P�4���fe��������ӫ�C�:�ո�bHz1ꐙF^"��yNU��^"�\L��(V��=h⡵����s�v왧q(b�{���u#;�voe����x�EN=d��/��Om�h�غ1�Y������u�S�a+�n�e�;zy�ӝ�|o�`�Үpa�|�9�fm�
j}��d�V=�o���1@�k.^�On|������ɳE����5L���f�(e�z:����������|K#*��x�a�5���u��Q�`��Ϸ44&��[�qwZȦ�Pڨє���#�������꧗#���V��٧y�4����Mf�"��rmfV��U�,K;�����>U��L9g��R��w��.ټ�c+.Wr2����)Ko.�X!CP<��~%�us3b���q�0�cn��Ьa�qG��!����rkˢ�*�Be��l���Ԧ�*��u+�LLO{mu�����M��:N��a�"�+z�b��#���i��7+O��,�u�E��P3K:�T>��9��=�;n��۳�n�H��v�쩃�d�����b0s����|��'�<л��r}�0QJ����ެ)V��K�i���*ފ��̝0%Dm2hw5`u�X�dYKY<����3zc����t�&S���0djG�ɴVe���zf��<g4�^��aR�WuI����8�N�cv�֤x&������.}B������c:�eX�E�Ox6�t�
�ǂ�U;����a���;�z�k���Lݘ�]�^��d�Y�|�	h����*��-��.���J��E{p�mT�*���4ZְSA�bV�ٗ�J_�:�M2�Ѥ���׼�T�_N��o�y�Јn�4|��ݸ�j��[�R�ْ�F�n�w�Ю��-����3�*`��JC_V�),��A�w�.xhH��Tj�gr=��u�C�Ї7�(!����XT�C��5�'���a�\�j�]d�R��� �yY�r`Wr�kj�ґ�u�Dn�,���Vp�6�g66kt�'�z�k�Ki����;�!�9��l��8�&刳�_���'x��&�4��t2��2�F�j�Y�.^�Z���rY��.f���Gxw�[N�&�s��U7ھt�tѿ��U@��,�.ZJ�y7�� h.�(�V�fd�2��_�%^���_�{S<�N�nu[��qÚĒ���<�Y�`�A�r�!�֭.�fp���{D�(U��
ث1_Юђ"×l���:�wچd͂�l�Ē�S�A�W��g1q�ʦN�I����=u��@�Ijh�z��C����ܴ�b���Q+����嘑Z��>���ئb-̴끮�b
�2���#.����5yx�[����y;ZM��(q���]%�Sz��r��κ̫��%�����Ks4�V@uЭ�P�v��@��u����`�P�3�A�`�����{*z1��|F�Җ��A֐*WI�vv2&]�7�4��{���]�ݣ[�N;$b��b��q�<v٥hԙ��R�s��mB����F�
�I�1�F���NB����}gl*c�<(u4ӝ�7%�bF�yA�{�.J�7n������y�u�/dɩU�E�{E���c$�;��L>��E���&��d+�݈7����n�˃�&<5ڬb4J	�{���޽`�CVi�1��u'3l�mg	��m���f���D�@����,*X�E�w�,�ã{�<ݕ[I��+�31�K]��:��A8��'c�v��&޻�ه��t��Ϟ�I\�(������{�����E�2�T��^q�W�R�����k�BG�}{��r�W��Q#��`�܍�;3���´��=�Z � ��_�m����M�|z�%+���/Eu�5>�q:id�]��l|�j�K���cZP���usr���ܯ0v�Fd��9�����U�\����{��:K��@�����u"��$�H��a.�V�b�8f�e��khs�X�"+{�˛\��&]�����7��Q��kAm��g����J}HwvS
��0l�n�K���`�oqT|��,4o��b�l�g/u�o��U��Y%-���˧s`櫸p�(e�bS���0�{k�V�-!���8��+i�HI��ج���V/�� ��,P
K5�(t�t+L�ʸ����F:��5��!�c�άƃ̢��wg#6V2�}Y���g�=s{2�1,�օ7��}ϢQ��#�9X[��9jŵ�uLONN"��T}��p.�Ilط^��C��;Ne]Cm���'E�.WhѴfb��Q�ឧB(��A���e�����8���F�bc��m�(T&��{1�o �ђ
�\|gc#a��om��m��Y�u�:a<�Zj�9�RM3x9�ofbNs�F	�d􇴽,Ӧ�G�x���i�Bi���������n�X� �O��>�p�����ښa%}v�U�6�1�k4d�NE\KwEvt�Ԩ��د�j�ʊ���pbƅÉ:�gLp��zg\���9��Sm�|�V����2��8��1;<��RY���B`�^4�+xӵ�e)�O������֊�/(�ƻ\���9���������,����1!Ki���ɝ��6�[wgLD��鼨�	٫��UэP���XqMłW�X�y�)j'�Q])���8sL��K\]ԇr���F�'V�Rm(6h4�pN73�e������k�)V��i[፨�zR%_v�\@���nq���]������9������n�z���Wej�%9+w��=>�6�a�ط��=���m�N�z0^'ݓ�ObG��uӜ6����p'@	��wu��Hr�q�ިD���+ٕv�yO��c_NL�Jf���юܓo��ۊu �a���%5+G&S�|�T�R�n�l<pݗ}�n�]�@���mm�-}�����H	�|(0D3t*���崺��H�7�Ctݣ:�a�c���/���-H���/�p�}&�9}P6�t�O�鬒�koKg��SPJ�蹴u9:���R��w+����8�|�e���V��ίyb�#fK6dEa(n��V�����n���9��%Yu^��l	=��z�>Z�gq��:� ��
�6:VjV��'ʹ�w6�D�4��Q^�;��mf�,V�+����I�o_.e�{��@�/�M��{�R4�,��Avr�B뮻��T��wz=�#������th��l9P���6�T��;p�+�.���v�(u���Ž��$���j�-Lu�X�;���L��3�hCz���vk���]�f���uG���AZv�K���m*S�s�(�ݒ�_t�MvC[�1��q��Yrs�e�Lm��b����5����O���kǌ�#e���v� ��(����!m�����dB�E��Y�ŹH��꛵���O�2�[�9���^��g���n��a�~�!�{Z�*�\ڽ[�%p���b��a5+��D"fmA�h/Nwew�n
�[t��/��Ă���zD�͍��if���b�(Mc�v��d��(��Jm�8AR�қh<�is�_Y��I�Ӝ:j��ܢJ�����JX9]�ְ,"�{�!w��t���
/.���N�:�J�)�z+m(c@9:.�����j�V��$wҤ�s�d���9v ��q���v1�<��l]v_P��G]�d9��O*l���)�k廼�1H�D�M�ϔ���1��^m�C�͍�R<;�t��(��9��#jX�`�X/��M/٢ˑI��M��Z�H���m܋d�c��������>���}���3o�k��E��g��/p}�V<Z)
*�u�t�+;�J\ɋ!��������c�q��"�r������D�+���YO,;ט[������)VC��f��Y�Ô�#�аd/gJ@-��vpGjCfP�+8�Jf6���h.�mmȯg.��"pq�����f� �@iy��\�"�"R��䱙�;����S��� ۨ�<Vf�������v�R�1E����]
 X��kyN,��;#c�a��ܫ��8`���*����a
�@�k���Wp\60�}a��M�U^�B�4�]^]7V ʳi����e������2:���c
��;4˶Fj��॔6����	l
Ӛ��[fV�wIyA��97���F�ݑ/y����/Eƈ���*B,,�̼f�\��kq6��<͙ ��CX�YݝС�pif�~"�ZG
�gU�Ú�s�1�Q"�/;��q�l6�-�kۗ�{of�=�،�Ɋ������o�-�l����j�b�T���f�����W+Or�׍>܎�46��(�اܪ�DQl��͇�t�y/�|,:b{n�T��W��K����r�w�+]�[��ei��M�h3�Q̘�v)�-�2&�{�����9{�a�R�̉��*����,Q]M��u�6��ܵAp��f��V�@Ӧ���}�^�`�d��K�P�[B�a#�=gW]�Go�����ܡ/JWD�(�h&퍋��N���Ob}�/;oF��9J�i���5
2�75��o`�A�6;8��,�'X���L����3�;��.�o�F0S̡�����2��W�iGI�B��9ܢ�V�>��|�j�S��i�;����xC�����Z�t���e�� ��),���=p;���97ь�Ovj�t�R�M�#aX�t���k8 ɳ�ϵ��1(3E,�k�=��
vV��PhҞ`�\�ωݝ���e<�|#��)a�g[���)e��%gs1�uki���ڛ��y�6�tؕIX&^
�ʍ
���c&[��6�L_���I��
,�J�,��v�l'1'I�b�ohdу�M qV,���;{%��`��4�YZ��ū{�j�Y�Ӧ������/��0R��.#.}z�Sد��7nY}�.���xQ�����UG��T�hgEt�*(_ �5�"	y�GLνA�)�2QH#��6�o�hgo��3��d=u��;:�Ⱦ�2��E\ ��P)r��d�ݙH,ʰ���&o�t�&�TtK�k[D^��^ʞ��+�VI�*@��MJI�E3^�Q�(jWyκ!�cY2Quz�#����be��[���U\�^�k��qAN���o/��u`�O"(���T��� �O\�b�'v�BsT�ҡ"�0+)X#q��ɮ��y.iK��}ۄ2�oӕ���猩"��]j�p��sN��6f�J��g$�Ǡ�o��ُ-l��2�� �[��h"�K6a��Z�Nb��5��MM�=�X�� FgwQCr��t��R�dZZ�T�ޣը�n�T��_3�c�����6�q�|�3g���S�����uYF�����C��
�׈������!��n���u�IV+M�+��n�Jv�zWn|y��Nڥ�w��j�E�&F��@dMN���؞�֖��j�V�csE\������g���<���8��}#��_�,�q��Ӻb�wJt]h�7*d���;M�����G��v��������b�]b��	�v%�nM��%lb� ��t�i�Ff:�/M�ґ��)a�mi�]e�Y0�/(�x�U��]�k��ڦ��x7sp7B��D�[O���f���m2;��vsW3F�[kH',�}��r3�^�
�����6�2S]zVR
u�S;9ĳf���B�V���l#S���d�ᱼ���e6wgKε����m�"	�z�gb����3m�x��4�hR�Ɓ;��|QJVB��}����ie��Ï�4�噋}�K�^��F�4���b�ByLo�>�3Z4�H+�;���rʚ.J̳��`gj�b�M����ڐ�љ�2�](XV�Q��z�1h���_ln��'Y�iv��hc��u���SS.h��y�4koo��@v��5jνU��vMPMbK�,}ty�_���z"�p�$E1zƕLm�(��864�Q���}�2�	ogY�1C�����̎0���q<�l���*�76�E@��ET�M�HH�Ԙm+�E�j���E[�wR�+��xܜs�c��D3��a��:���,��^˶x��Ny��������oU�72��i�]�m��4�w����\0�%����8��Qw\]�A�s����|vA��d��A6�W���U�� [W"',���6h��n�t#���Kiq���Kn:���-�#��X�Ȥ��N#�������]R�X7�f<)����)�F��>[�j�:&>F��6���{����u�#��^ 8�M��	�F�7ts�[yc`�8�ms���h���O�]�s����]��MI���$���$��׻G�@���ƚ�M���L��f�[Xڄ��I搫R��ڮ���j�us��L4 �I�N�o!� ��*�Qs�������αz9.���w���ŀ��ۆF�J��֭�&w�n���7�o�m�}Hh5��[y�y<���r��:�'����Nr�*�)	���#<�*У�/Y��S<�=��K{[���j��=��^��o���6c��|8v�F_`M�+��i�X��嵚c�f�X�l�'Z�F�Ꝍ����]�
�al�r�����Mf�wи{Q�Z�0nV�S�}��!/X\��"���'A�iH��(���ϟ�˯�b���vݛ���S[���
��7���+
�I�Yv�+S�F�3�/"�b1n�����I�ٜ�Y�cMfV��Ű�9tDj���v��^�8��(������F��/	.�����WWcc
ȕ�(]�x�l��~�G��6�y]&npN%[p�pޜ�Fz�>��y�
���E�;;��l�7�L�Bwv��C��K� �yD�˨�1W%��
�"zw�$[[{�э�u�X���e0;�u�x��)C�����,Z[�ȫ2r��m�� c���@MSVj���N��9m��9�u�Pwe�YG\r�ð�[#��g^��j�[��[�1���,���l��L1��@ �{�tI+��u�s�}��G
�*��ʈ� c��unof��4kx�L,lY���7H���4
Ztԭفe�l@��z��rd�K���h �l�>�����R���'��lo/X�෉�j�	nʫ$p���A�g7��S�u��Dyژ�*��TnR�9C�N�+}�3۴ .���-���f�[b�n�E�� ��)�F��R��}aL��v�7`65�
M�f��^���fJځ��uj�3����=�L5������ejWd=�ܭ4ӆ��}�9��Y�����9I, ��W���pWc�2��x��yǠSU��5$�j��7d:�"��(�fұh�k%D���k �#|w2ns�ʵK�{:0�kS��3�I��`җI��`��4�d@�My�&)Xwӯ���Ա�T�0���S�>�W>�Z ��2��&�`�_M�s.��wRn���!��"���X#=P�+���t�5z�-�R���+A0��&)`43���+ٖ��r���eq؄�2#�˔LL�����n�&��7z�Eun�M}kT�C��ʓ�����XsQ�E\ޣV�Lh��N5�d|r���'��a@�>]�E$�����f�v�;V��y�������!��V������u@�t���n��7����c=���grۤ�Q��Y��6�⻍uޤ�-��Ґ$W\�TU�Y۷�:���m�:C4b��l��к�:f��;���\�T���Nh�Qeh������+����Y�H��3�n���Uj^C��E�t������2ur���r�4(���Bv;r�f����E�nѮ��7{6��[ao#
9���ȷ蝜���LyO����ۭH�v��k�b����Hf*u������ge-p�c0������ds�=�N�����D\.	�6�ӝA�o�LF_S�%�&ǔ,�G����.�Vu����ޮ���0�M��&ʚh��<;g�7��,6(C5
Ɋ�n%f�Z0�v+��6\�:�5��Wݖ�źmt[K,}�\��#�Ob"�ݴ�Ze]u��.+/�$_W�5=gn8���b��ץ
�ȇ����k"�f�
 ދ�����Q�������>d�R��</p!�n��9�9t���\��s�.����РҗR�y��O+��<5�n�+���(����eĘ��#
�r:�(�/x�����,;��mrǧ�lj�X��k/Bth���:z�c��{[ef}Ԙ�pL�9�̭-\��vt�#��v�������,�,U�g%�	X���r��hX�qf��,����̵�^%�I�P��BLDTF_��t��y�����Ӛ򱫷�՟�W��F�aX]tFK�{suƋ�0:��G3��{���ͷ��M���<u�j�$���5��8V5-������Gv$�Uu$c���r�|��U:*ݶ^,���KK�@���2#{��c]�P�]�}|0�n��	��i�cgjTq�c/A�I9�Ig�A�����w8���y��j\���.��:C\R�շd7&�)D�!�c�grI�C�2�����RU�'���X
�Hvt�A��2ރ��6�T��uBY��|��[��hn9��x̔ssd�5�y\j3��oX4�%���P�;�J�k�p��\��肨�TU,u�w��[��&�3E���,O�Q�W�� w��0X	e�L��էy�M�F��`m臲�C9V�]ܪ��Z�W-����b��U���:JĊ�g1 3��5�+;^�yO��Y���]J'o�Ǧf�d3�J�odS7�"���2��At9��K��5ЕU5�m�\��.]�� �h�)"m��u2K��vܳX���aŷ�TV�Mp ���78wfF�:�.f�\M$B��f}�٬v�9`��kr�Z컬V��i��ɱux��ad �g5�c1VC�����w�/.�e�CrY�e�l�V��y
��iY���E�S�1��Z�u^��vp�ΐ�;��u&;wE�$�t5��:ޜ����9-�bp�YwV+9)\��ol�'��|٤Jv�f��������I��
Y�n�r/�y�,�H������gi[�O��p\����2�����=� 2���M[�J��y�g��q���nWw1�`�^�>ם4/c��o�9��[�T�λ����7&�mi�B��y	�bG���JdΝN�es��%�8��(u��QK]ּi�,���B����ԼA�to����#�a4��tb�i�� .@�ۘ2J�1�T.���`��iW�b�2�Ovb�o:�&���2�Be�9��G��ܳ�o�u�������T��t�|i;���(�T2D�F�+���r�N�Ϭ���N�+#�\��%���C6(G`@w*$�.�"�{¹e�b���b(d��,͍�unMf�'];�Y���b�i�D�'������4�|��hgǊ{<8�ӵ�SQV�vTVp�bwATn��cj�ݾN#0�V\�f��-U� r��eb�r�p�b��{���a���"�ص��M1Ќ��6������Qu,�|8Nn<�M��v-�;U�)�60vi�)�"	�/i]��RE	|��k�u��m����s���Mur�������3�4s�8��cI��1Y�u�������^bR��U��d=�֒��8 ]4��Uu��Q�� ��؝���-A1�����!�\��b�����vP�l�Ÿ�-�ۼ������ū���5{���	�{��h�RN�i�P��8�Jy�x�x��e�.�0��G8��W����:���6WǑ镏K�w��]�&@h��@��G1���Ű$͆�G_�2��y'VM�E[�m�eÚ3S+�������N�F6�rrj�b���ԯ5��^�;���LK�C[F,���Y}�V�ζ�P�-`���N�c�֧����u�r�ͥm �;�8�L��想�H��L�컧��A�MG�]��h��7܂'���Ca^:w�fRTws��bR��=G�KT��	|ɀE�`=�x��f./u3\V�M���@f�`=���&>�m.��� 6���F��͊����A�Y�-AX�����ܵ���o�Q�|+���r���Oi�#ʙ�#�*#��j+8E���݁v����\N�F��N� �c��m��_X�W��b�or�.鰖͆=����uʭ׵��V��Q�[\��w5۟*�	�r*4uI+�]�d�=ٝ{H�����b*�7n�-Aq���ʗ��
j*#��=f�!�d��;y[���{ܭh9���S��+�����2��ҴshTu���O�T:�vQ�4�Ƀ_H9���B�-�ڽ��歾"��H��S�`�=���W
�!��
Pn�#��h,�����C'�uk��M�Mw}[e�\w-�/3)�ۆSG(��܍T��业㝛6�n�32h���*�����_lI�}�6�`�`]��)@�w��iZB'��R�l�y�n�N舢lg}���d�f2=�ۡ��qPD���3:6�]�:��H���M2�����U��W�_}�W�:R벤C6Ҽ���@o���}ڒu}������-����d1������mج��1G&�	C=C��P��<�ͱ�D���;��֥9�X�:~��-�l��U���{���ʃ*f>�4���qr����ˁ����֘�[��h*GŢVT6��<��sE��ق����Wo$O,�W�gf8r^:Ӊt�Ic΂��v�x�F��;f��R���]�(mY���T��Fp���ʔ�'p�/�V4��̏"���2��.�kP�ENP���z
��%Ŋ���0A7u�$|�k'j*�4��Hl<�2�sV0r7M�+Ʌ��E�� �O��y�U�A�!�B��$�U�+I�\��1���9�z5yڣ�`�z:ǭ7�Nͪ4�!W�b�e���+�(K�Є��q�<]K;:��t��{�:֘�.ۗ�����B���`oV�ʕ�- �Y
�m��C�I!�L�����;�s��.h��󾄫�K���Zڻ7�#Ʌ�I�����҇]�:\������Cwqۄ�Zy�ܗ�u�����X�qwJ�i��ݬb��t�����B��X��œ�ޭ<mÏ��Q �<�w�'^L��`ߊ�L���Z���J���$;�� %���e�ۂ�:�IXt��1�"��|��T�Y�)v���J<��S���s�g��6���l9誖_��/߯���}�{��E��9cETIYم��a�eX�����fdQe�fff5DDRfVe�e�U�a�A���Da���ff9Sa�U0QFYe�0SFfU&XQ�Td�AVMfVcYcTd����UUDe����1SYQ1daEVa�fQYcLLQYQe��VQYSU�fX%��S50MLAYDTI�fdY����9a�Le�DŖVY�aPCAE�eSf51P�QVfXETSNYS�QQd9PQMEE�VC�TL�RFfQe�f�MPQY9Q3�4�e9DEY�E��ז����ֻ���}����H���b�Od��q�:�s�QvM�M�%7���U��^��gRvYz��%1sW�_��������5�n�ƻ��}t*'u8�p#|�q������t=Sy�5��\�gѻс�ج?����ϧ��ͅ��%�i��Ս�z�7(��֕nˁ�m��T�b�"�=�������ʳO�؋��r0</,7�NTBb��$��zLA�j�6�ݷ�
�Z�l�I�f����L|eC��Q�s E���e��V���:�;5)�Q�y֨3��輡�;�o�8�U�k�:1`/���3�o!��om^nÅ힋EN]�5僫�M�'M�uº^���9�{��`Ub0k�N;04���\�5����C��]46��Q9B�e�=��hϹ�}n�T�+;�Sq�QǨE�c���?-�Vn�	��+� �o�þ�/��� ��{9�a�J�z?d�k}@����P�*ZdXj5���hg�.��q�F�_�Lc}N�k������N����P��=˶lZ����h�)n����Ń��Xr�ͧ���n�O(Y���v*[<Gk����U����T�X�ϸº�Τ)�^:y��wmt	W9�w'y��y�Զ���.g�0�k��sf���tM\c\��B�yuu�i3X8vGqqrA�}��_�S'_�J�O���GOV����n�W^���Ϥ�<9�O�h�������y|K��p��m����8��o�H���Xɬ��ּ�L���d')�����crXZ�����i��LW��ލry�9��	0��ASW��%3���1���^������!�__CR[�'�­��ѱ�����`�'Y�l����׍t�ufk�����,t���{�S���I[����we�/�M�5�]�7�Ղ3h����{+E>��F^����	7�*gƹ���o*[�9��C��ˌ�3xvW�=�.��ߦ���M��V�����kV�U�>bNt��:R�p�t>3~�ӕ��U�8�f֮9�uԙJ�'ay�]��+���g�EF�w���$�;K�j��N�{����4�ghmpfm�GV|�ަ%u�d�H!�)��E�Yzg5�kgB�	>���ڻF�9�8$n:)���W��T(�[���1f-�(n�uq�q�\����������ztud�loJ���W�+qC�\זK8y��3
2	����*�I�r����t1�Q�N;04��7�7+�^3���y�u�.��}.�uW����.{^�	����)���o<�Z�I�SP5�i��Zw�QZ�j�:�Vlt(�,V.y4e�'��#>���~�}s�$�jM�y��a�<�_[���=�\���wL���vxl�>�ϼN���i�䘸�����N��]��Uuw��K���Sj��{ z]���.s�4�v	�]`IfY��3R�9����،�1G��<�O��b�K�>5�>�z_oy:���}bn-�ϳqfvS�����l�*�Tׄ9b����|��>����X��Yul�ĕ���P��`�}���<t?}�y��t�k��u/7�}�=R�^�ET���#%��R�w��T�3��;!���04@��c*���4�V'�ظ�*襔���u=�M��s-}c:�+�-$U���{C�C���ɒ�6�R���AX�Wfӛ9�Xeo9��B;υJ�ĺD��%��Ǹ��f�>��8�Сn�k�o��@��xh,�(J���<:4��]=�_����E)�kos��s|�7'����u��U7 �_	S�%`��9���WOnD4'n��ձrӜ�i:��?s�¥���T�&�\ޮ!lɗ�,�q4G=�0�!h�`Iݞ����S��������@�t$.o�����\�{����3��(�9@B�%�}�6�o:�.:��w��ȕ���}�I�sT�ٞ��T��U�(�az=�,t;T[Җ]fh"g&4�}ѽ~�����9=~Pm.[�:��jn5Ac�T�X��j���k������'{�'j�5�[[7������K49���3+ا={�t�uJm���t�`����z�v�i
g|��'gY�Vg�����q�w��GxAM�3�6���L��\؆w=��d�O-:{c�3/A�.D��S���YY%d�^����d�yPg^ݷ�٨u�tӀ��L��Kz'I��F�o��;�![�wJੜ��m8h�@�K�\�3�oy==��e\]��`�o��4Vv�=��	�r�6��k��M����s��ƴ#�l���Ru��u!�%`����>��O�R��j�ڙ���n?y6�Z��ؽe�f�	k�R��>����q�8m"a=Ǐw��|�����
j������Oz�����3'#�=�PHiU��T��C���	��y}:]��v�B�3¾/z�C���.����#�皯[I���_K���&��vnv;��vʅ���_�k��!�@�z�Y�ׯZ�6Zφ���鼩��5��m�X�<��9�8��:j��hZ�^'�f�Wʄ����|g��Oυ��N��S]h�W\U�$����Q�r��M�1�����'w�oI����v��+RWm��'v��Z'яW��\v<&�W���81�,��v]����rT�{�}���g��A|��΃}.�LS����;e�\i_��:�$xG��սx��ij�n���ۤ4"�Ɩs|ɥ7�K�T�_
f�����{5  {���̮��ަT7e��[�ˏ��㡀鰌����%UL��~-K����{]��������y^P�����v�f��5��mh8��1�n�cklw�'��U�N��w���-�j�l���~��{z@�y13�F�rc��r@ד�ո�m|�ڊ�u�o%�M����3(d�����G���χu���d�T�>��U{�%���(��B-ؔ5d֞�ԯЕ{��?8��X�h;�z�B�1c9�����=���D��{��WN�#�(�(I�k"A��,�il���Z�3�/�L<{��t��;wk��S�����`rC-O�|b~��VL�^}yx:ᚳ�{0̨~C9J��v�'��Sɵq�s�f�Ŭ9jX{e��:���{��י�;9Q=�=�1�uoyXw7��:s��m!��7���EK�}��gf�q^�>ͷ�{�mr���� ��U�\�E�P�9�ޜ��g���.�쫼�܆��~s�$��[ϨjC|���x[��cB�VF�֮���]�J�`iD���v����}���.�&EZW+,�å�n��u� aK��2Q�oo �������W������H�"8WS�[ՠJ$��ûdc�eur�:Gr�'"�Ƚ绗aɝj3a�.���d)7�<1���Mٓ^���g﹣W�ꦻW6Ǻ�����ٻ��L&ⴣ�j}Ok���a�" ����W8�������ޑ�>�e��W�7I�1mͽ�j�6��8?	��9��f�ð��x
���o(g^?s��WM�b���U)*���NS��z�s-X<�3��,N����M�wԁ�^�;���>��bb�vͱ�*�͹�Nt�z���p}�کֻ����Xf�ygP�zO�0,���C��JA8�U^�����=��Ⱦ嚖�|�����r��]E��<>t��V.c�o�+Y�6�W�����s�{s�-�o���X�O�y[�1��J�\�VͲ6P9vqo"����^�����N�5P��̔��9.u��+����.o����MwX���t5nE6��W{͎#��.-:����Ffy{�E���)^._��l��n�����hfo�o�j��,�2Н��7L,��;�
��Z��u�=��In�G0&,>qO�R�mwq�Շe+��s��	r�:�͖�oQ]$�;�uu.[1����t)b�c�~���H���.�S�j��:�����}nl�\�K�N��%��vw���O�b݃v��w��n��XO�c��K�oyXw7����K��R�ۈIS"k{"fp��/��b���C�1����̍!��8]��W6kx�� B��i����	P�9�ASA���ׄ>������=;%<� u�=o�1�ّp�>|⋏��k�����[�vj��b������_d��`���.v�c3�4Ԑu�m�+���t���*R���,��)�����{7=+���;{�;b���:S��XrlWQ�Fn�#Z��O.��j�O�dxB��w{��<�:r����9��i�����c1�s���6��:�s�X�|-Mݛb��Yq�3;��:��>v���*:ܪzw��4��\����,t;T�ƽ�e�`��#�*���(nq�$��^��^�b�\Ú���Ў� �̓�f+�;]���]BOP���<�PLӠ�fo����t�tsH�}�pb"��-��Ѕކ]�u���#�����B������1���k'�d��/�w6�1���/�Mwl5��'�Ovk���b�
Mn`���j*���X����-�^��;S����~��d��5���vof��j��"Z�wsSk919\l:��S��:�f�t�3�=T$�8���+�j�؎�w	�!�^�Y�0_+z���_ΧL���kz�MN���4�[�-vtU'iP9/�J�
���y��v2u_���T��>�Nq���7Jʃ�͜�����o��_�b�t�5��¥u��y�K;�O�Q�����~��S�[UPN�3����[���<(��s�]�c[Z�n��ۚ�My>�Fc�t�=�8n�S��/1SG�+��eU�뮄Ș�R����Ǥ$��Av��N�=�6��C�P�*�Eu�/�ƭK�ȼwV�H�2��{|Gvm;��]�`��)��lm��&x��z�[yyn�٩з��|��m��˵%�^Nl������-g�tc3x���D��Գ��T��B�:ֻ�M��q�M��dS�w�c��\�����4��9� F�}-]��j��z��]a�fQ�L3.k��Vz㼠��bh���w�R&>�OI��~s6����KT�����\���@ڵ1�� �[�2_��:�^9p����ΙGWm~Ժ�Ӟ�e�����E��h\�5'TT+�,��_��=\m�^s�E��YH�٦�e7��<�k|��~��w*�����~�[���=Gr�뗀�bLV��uZ�}�V�j�M�'���p���M;�I�,�Vv�ܼ �����Nk�;6W�f�KrW�j���q����T{â��u�����`^��m'�.�>tx���t���RP��{�%��Ҏ=բ�T^8�v,�	l��8v�+N�#^Y��^^���|y���O �Rk}^�_�7:f����t�	7r�����YN�[.�B��y͙(��b�kD�ބ�R���fV�N5n4f�.����,;�R����WA������<�Գm�nDUl͑��n�9^J������ky��K��4�%�88��*�G��v���
�	�ge-x�����U��+��Co����y׶��D2��$���r89��d�����y2��Ilɐ�U�f�E�'��x܁e�Ǣ�N�7m��d�zm�:5n�)��[�K�=|2��Ӄ�Y)��6��ܧ���Ò��e2X&ݵ,]�����#4-��a췼���}�Es��M���k@2�z@�L���	�������9b����ur e*%e�C���#0�ii��NK���j�N!�|�Yυ��@�
��p]��J�"�L2�;=�o9i���k)p�# �帹pFW�4�������t�����ۃv4�R�G�*�@d^��j{�Դ���
��CWa
��������j���>-�.�hp]Ř�fj̗\�[{�V╨ݕ��'���Od�s���J�z=8wTf�1gn�Qj���&��*�0���+��������7^fo�>��L��t�oRǛPV;�r���'e��6��q`\]4fj�QT�+�O^R�Oj�R��;�g��*�]��;iKF6�m�o�?n�͌5[MV��ޚ���y.n��.i���
��ڎ��N�^�]�áZm�U���K�Ip�sb6��7�$���4򳾌ռ
>�h��u�C�S2]w��B�	����)^��V���p��}v�mCX^k˼o,���
�׽�P+�]�P�1Zw���^�kG����z�Nb�W��T�-��QC7K���'
��v��p�w*=1��B�}at��`ώ��4�D�'l���Η����A�����* �w&u%�()���0���oڂ��4�fwV�v�9��q��*N��NT>����̬���w������8榪��m�ϲ5������+K��]��d
ܥ�N�YI���a:;�Fp�g"�0�U�]���ZǠ0��U�h�1*��2'Bcj��4_w2��ͦ�o��Q�S)\�G�kWH74b�9WOf.y6H;����֏ح��G�_��n9Q�ǜ�����(>�bІ����wv�x�k�n��������A���X��N��ര��տ�K�P�����M�+9f*�*�1���l�RG���.fl�7c6��!-�L�q�fj�����+�Ӏܝ�zQr�*��I�p�}J�4�w;X�4+��ZWT'�ër�<��L��f���Mv˹mͧ��k�����|�k�����C7^0Xz���_aܶ�.F���!Y"��WGNuN*� ������l�o������y�G +�N:�R��C����G]ƮO��y��]�p	�^��[v����7���Y�IW���6Ӹ�&�&2O�[G������U}E=f5c�T��cb�FT�Dd��S��MDf.YUHa91YVfPC3��EMVXYeLP�MPUfeAPY��USEE�Y�3UD�9FA���eX�54SUU�TTTQSDUK5IQUAPUQ%QUadUEfVVX�1U�Q��faUUEEYcSY8��TIESQRDL�fAUM%Uf!�5QETL�EENF�IEE���EQEe�DT3	2EPHA5QTT�DUUY�UD�A5SU��f3�aDT3AMRU5LLe�X�5S33�4AVN@f`�514$Tљ�Cfd��PEAkϱ���뙗F�`띺h�uv�b;����1+�i�j]��w�:����2�G"m&�t�Kn�~ّ�5����/^�\��Q���7�9�ξ\jr�����e_l[I���v�K��c_�v��*S<��tǥ����ofs�}��E[�]�ߗ�{�|�8G����|!�o��,-�|��x:�a�jĹ5�y������P���M�є�!A�Ľ� ��|]�K�������4{����S���Jn�t�B��4�NF����X3]���R�:[�Wp���U�b�8����o�������X496+�b5����S�~}ٚ�0US�}�Eԟ�sF��j�G�=]p`�C���s>k����e'������%��f{0�խ�-���۱�q5�`�q������=A̵t����i�*�2�;s>�,Nt���'�g�)�~�=����6�=8:^�Z��.Ś����❲!=]Ee��9���ܘꕈ�҉s�}����e��
�J�@��E������Q-S)k����C�ˡ�_U��ɧ���2�s=�׍@,m�Қf������\���l3Eb�E�n�yXh)}|�=W-#w����ԶO��Y��s�(�=.a4�̣c]tӏAc��杁���	�7su��݂N�Ĥ���׾�9�S�J-�E�(G�:Tu����SU��}�=�<��,�N�Ϸ�7����+�+�+϶V>�>F�A��R^��uz���7��o����ԛ���_���=:�
dAѤ�HM��]�>����@�Κ{ݎM����Ǽ�u��?_��g���m�"sϪ�(%GOϢ�R�v�����މwb4�����S-���:J�鋧&\�}ou~��ڗ�|�x{�+��v������o�{hW��
=���__czq��>���i��m).H���Eg�@��t
�T����}v��z�e��Cb�@�G�s��T�췊v?>R�jϢ�P��� ��������'�WO__�����8���sIz�Ϧ���u�����+D��8X�k:rk��@�i[�5���]2��8n��w�-qX+�m2�CVj�S�V�]����R�ј҂�e!{J�DI}nr��e��Z뻥�-��y������[�[5A2�+o*�
�a���|����8�m���z�v�~={����N귎���&���N�ັ�h��n����l�0����{ϳ%���4�E9l_��Q�[ec�Sz���i�Il���e�Xrs�c�,*i,�vm��WF�/]`���c��qsV.�)�f����N�輣����
9���܈ﺳ�W�=�B�}6��v��\݊0��N-�w�&�0WQY�[P}Zgg���6����T�o�V#k���d��5��]�f�a�ű{��*z"2s����m��(%��]՟Zr��B>��sS;��\H�\R�j���(��OC>:�Zޡ�ޭrV	��K����r�6U��ͫQkQ[x�r-~+�p�M`*�_u}�7_}��v���)���7'$?I�;�q���ҙ.���z9}+�?k�=�5ώhx�V<���;?9������}��r"����_����Gsٮ~�u'!)=���)<3�ù�%}�q��'#�_����~����仿O�{���T��{�jǄ�'Y;�zE��p�-�/���*m觨7{�e ;G)d�D-�Y_n��6̗([�,�|��D8v���*�6��K(���\�φ�9�:�i��鷒���VcM��+mε�u�J�%�A^i>o|<�o���" ������?}�����nG�ϵ�;���翺B�=���]I���%�
O�>��xF
�g��@dQ���'`��x���K�����m2_��?f��/��9�������4}nGR����|��x�Gqܽ��:H���}.��z~�pd�AI�`��~���^���w��w�{߻��߼�ڻ����,��:��~��09.��}'��H{!�;�4}n!����:��;��~�?Op��t� ��t�����g�<��o^��}�_xw���;�!�r�9�w��G�}���>�W���'���O���!��M��G�zy/ry����;��)�o��=���o�s]������g䜼o� O�}�Ӷ���D}�<�!�r_5��}�뫾��{~�����C���{���rN����>�G�3�(Y��~@S�u3=W�5�}��k�%R�;��%��~��W�~޼�u׹�r_�b��w/�����܇���$w'p~�.K��Jo=}��-J�g�K��&����~��Q��z;��R��%��
{>愡�^�����O������W�������5��~���~�܁���ä}�>�}���W�~���~~M����#�|���ײ�9O�h��GF����
C��A�����愡�^�9���K�?iu~��ش=�_ O���0�w��ܷ�U�ރ?}�y���Jq����'��=�<������_ ����AJ�t~ގK�����>NA��4���/g�����_!������a�p��ߗ}��	��|�������-w��H�O>���z��z��rϘ��Ի������߻���W����r]�@��=ù|�ӛ������ֹ�Z̿}���V��B�Af��
�k�����%��G��i6<2x�c��������ʿa6���r�E=�����5�[��y�"� �Oz>U������[�����ŗ�er����H]��T�z�ܑ� �y�L퇾ة�.Ys(�������΅V�✣�/����_��6�����ش?���;5��|����9�{��R�
_ؾA�yk��w��Ӹ�W��7��w�>���^wC�t����K����/���1_~�>�<��}��4/�����j��:�|���vk��9w��)]u�
^��?C�y9���;��c�^Ku_�d��7ݾڟ�_�����?�P�痒?�|��y���iy�>ߞ��B�!ۼ�%�O�d��Ի�XjW�9���)]={�ܼ����~��P'ޔ}?>=U���}�}�ȏæ��}�����м����wy#���C�|������#9ޗP��0=���<��X� �]�FJ����}}�v���~�~_s�#��wX�����;��y���2]��{���C�7���nG�s�H}���9��&�~����\����<�%�
L�����f��7�fa��:��[�~���)
?�y��ԯ,�r�w)�`n_�����ҙ.���z��R�9��������w��>�ԯ��Z��{�\�_��o�z�����x���Rt�ra�����Ox�GR;��`{//ҟf��?���}hO`9'a�k�p���`�y/rw~�\����{�o�������w��{/~��R���{�C�(���/ђ�����F#�yw��������/%;=֍�����ˡ�����lV~������;}ןy�_~͝K�?@s���=��߷�@����_�
Wpvo�t�����I��/N���u��w/��~��;���O���N�מ���}������_o��=����N�G�9+Øj^C��撃�|����Jre��_�
G���_�]FB�{��%��٬]���ޱ���{�����4}ׁݿ�`�WO
���*W�VoP>�C���<x`̾訫�J���)�c�x��t)w�Qe,�2v��t��;U<p�V�t�.���Ֆ�ˆ���'�o�;F������|!�r����5d��*��nF{͆�>�2�{�wPv�a���|y<��5��X<���>_Ϻ����&��p�'~y�J�d�}�rrW��z�pP��撃r�=���z�?t��o^t������?3� ���(��+n��?_�{��q���}�۸�X�������;?b���g�k��'�a�)\�����Bw�i(7/��vsBP�[�����?}b	z�GP*��7ߋڷ�߾�W�������$�C�{�F�~���G%�����z��v{�H�I߿h��G_����2S�|�+��}.��X|���o�=�i�?�i59���>����ڽK��y���G���Zגf�?C��jN�܏���u/!�>K��pZ��{��l��8@'�����Tnݝ���b֯��ݽz��éFJp���n_oa�x���/�����Խ�����������=�a�w+�du�'$܏Gxy=C�	 g��i���@;���Z���َ�y�;�{ս���G�|��ޏ'�_�{��q��sF��^������������mB�;?b�O����w�}�"/�	}�q�{�>�U�{��K�����?A@q�.�ܿFO}y�~��vk���w'��G%����5�C��|�^H}���B�!ټ�K�?��X���^F���1�]�{�_�������<�n�uO��B�n��d����仌����A���ϱ^I�7����G��m!�>_C�b�A�}�����?~�{|$�XjXqL��������d����'�5.�#!w�X����M��d���~������ҙ.��x��W�[Ð�}�+�x�~�[#+�r�2�n^����J�8~�}.I�'!�
O�>��w#�;�:����٬M��d��7/�����ҙ.���z�¾�
�Ejs�����#[������
��W9�hLB����,V�����Z�STy���}*v��a3�z������>�0�X�xk��0�y`�s�͙�stM�\��cz�������q-�u�__'�K�n��٘-�v� #��n�L��aa�}������{w��R��{���PP=c�2���1��^Gf�W�ww���#��9/�p�f�7��3����vQ�Q��ݍ9�����Ҹ�.��}�y��=߹�H�=���i5#�=������wK�d�k ܞ��w��G]�}���w�W>����γ\����~���l2_��?f;��װs�id<�����K�@x���w/��s��u/���AB���:]A@�}��%�2\�ܞ��ծ���^���j�y�Q�*?ڿ?�����.�W��}����a��O}��C��o����<�K�=���hy=���9ށ���οt�!�޿t:����]�߻���y�y�=��~���Ò�/5��_��u�X�����!~����/`z<ѹ�A����NJ�����w	پi(7�S���y���{�����Y��֦~Js�����߽�k쿄���KK���X;��.����C���!w��C�r^����n' ���<��:���Gr�
�5���*�䊫�U��yOw������<ޔ��]�ގ�y�.��y��Z_��:�܇�����b������{�p�����y�rG�2��Z�
�[���+?BJL�g퟾WUw_|,��=�pP���p�/��q����z9��^��y���W���������NH}����p�G��<���G�L�����͛�ۯ/��U����y>�����_ �N��G �|��ޞC��N������d�������<��]Kߛ������ג��>�����[���y+ۆw�~{��$�G��qԿAK��=��W�^h_�nOw�#�_������Jv�����_�a�� =��|�}���������Q����4��;'�9��yV��.��`��Wg?~��ժ��%)=XU{�z���h��pgbK�t�j����}�2��rK:����%.l�j�S��M���v��Ge@�(�� v"��ǵ~�ǔܑܻ�b��+��r���9U�M�Tޡ|���﹬��<�߿[��)��^��:��.�#��O��G���u/ �������^i�ܝ����O�i����4n^K��|�^H}�~���y՞����;�ۮ��~��=��!��>ڗ�<���O#�}���~�#��9���r^A@~��w.�#���w'$��Z9}?}��<�����_��!���٢=7��z�~����K�ۗ��K������C�w	队FK��AޱO'�w=�5+��I�)�;��<������;�q�ٿ4�K�5�����f�k�~�������5��kg�]�{���nG��Y�|���ϴ����럺]I�N�1=���):3�ù�Y�_`�w�'!g�g)|!3�?���(��9������ܽߧ��ҙ�?h��G�{w���r?�}���}/|��C�_g�~���O�;sA��'F`�Eh��¢���p��>��s}�u��%�I{��[�ҽ\�&���)ٽh7.����H}!�;��[�Խ���|��x��w/|�·R;�����@$�� #�̀O³g���W~7����`u��ъ�&���%~���=��b��kA�w��xo�!� �0��?���~��;��;��?i��{7�:
W�a���>5�g8u�y�?�{�5�}���r
����s��k �>��vh�w/��x�Wqܞ×��>��p���<�ZC��-����7���_ �6s��~�_k�����g�y�����{��AJ�;�ΗQ��}��!�r^�X<��~�������,��N���9y)׾�܎C��dt<G߈��o�ܿ�r����ޝ��~�{����'���R���o@�e��ԯ$�z��d/���~��5��}��WgX�>��`wy#��� 4���~������*N�û��
�r��$~���.�lT��wN<�0��YJ�|�M�8����]�7�d�Z���bC�qY����m�謝����G��޳����^�r0E<&��.ջ�Zj;��o3|U`�q:M��������#����}��O}�6���G�D#��G:G��>�3{�ܻ���|�Pn_ ���hJ%��?tw+�?o_�]_�y��-/߱�`�_��y���r5��<��7ϳ]u��5�����C�?C��GR���%rr_>��)\��K�)w��w��~~愡�^�9���K�����?}���{!���[�o#5����s�����O�>����)즺��ܽ��}�yK�+�p_�r>ÐR����q�=����g �sHy/���<��]@]�����{��~��Z��3��������Q�x�?��u����O~�w z{���^I�|��5.௺�B��pv{�<��|�Ǜ��w�~���_}��y�{���g�s��,it�"��R����߽�}W���S�k�;��C��^�c�_#'��C����:�pR���9/ �ï4����R��u��hצ���:��{ߝw�7�|:���9�K�w���Hy/��~9�z��h}�p�?�`>GR�;5��|�����J�t�pR���w'#������z�}���:��߳�/�o����'���w#쟳��w�?��G%�>ۗ�b��|��~t/����r^��z�?GR�22_�������O�}�s�#Nh��Y�;ʟ�����k�������������9ߚS%�?sG/�y'�ޞC��{bC��_��/$y럺]C�N���r_d����qg߽����k�}�o���p�WPu�qԯ�n�=�����?C�w��~�L�rtw����<�<��r;�֐�/��ߴ���C�e��#��|8<���9���j����~�y׿y� �|����~�����a���;���W�X������^w��t�K�:�z��R�o����>�>�����B0��J޺jy���;0`��0�-�֞Z.f��9��î����1[me{|�B��%�v�:��&k�yZ��
uk�s�;6$��Gz��(�:�j�}p�x\�l�W��y������wlZ�$���	�;4ը���8���4�C���yz�u�?UU��}O��P�lk_V_�}/��ևPP?�1�/�RP��y>:0_��t���u#������)����p�}��y�7���R���!�O�H<Q��O��_���_�o�~YK��^�ߝ+�9����|����/N���?Of�Gr�:��!w='x����o�ѹC���s�]����{����O��C��C�������ܾ���� �^�u���w��K����d��K�p�/�a��#�}��r���|����W���J�jo���.�/��_�R/d�:��NJ��sGR�`?9���_ ��|Ҝ��{�_�
G��o_�]FB�nL�۸�r�/:��.��]�}�����3�>�h�]O���/ �'���=I��}+��}��7'%vsC�(Ow�%��
{w�	C�=o��{��?��:]FH����������ߞ�}���y��߸4�_@p�/�C��~:�y��{�������{��<�%r2N�>Ѹ)\�>ޞC�(N��%��2N߹�(|�\�_�}���C�d_���������G�}���Z�����ѬNH}���u��S��9/P�O>�<����{�H�I߿P�@'�DX�������ZUV��3����j~�5߫�O>�^mT�6QY��>9��{�S��{��V�l��]톄��c���qnþj-�����LnH<�� �Ҷ�{%^�������M�b�s�Pkt��+N��5r����>���x��څ>��K��_p���P`�y��@ԂAE�]�kt���hJi�3�B�́�K��[�Ϡ:9��:�m�J�}΋v�)�M !��!�rQ�1���k��Ѡ�Cf�P�K�=�XPF�Z�l�2S._Tj��C.��m��=Z؃F�-�,Ӹ��NRZ���H�Ø�3�gڦ��鰁�n� �+747�m����j�qP��49-oBD��$�]���(eZ���1�n�)N�JP�0�+4Sn靰�VsbWƮ;Ti�:
͛ݽz�24�nt��ou��%�@�%K���p���oܠ��P�t���V�u}��].�i��TG'M ��_as3*A�G�8�9�&�:��>'X�h@�3�	�T�C��jv_
��
^>����ƛٞ�qJ�7s���Z��4F��l���-��ʻT��^'���� "�5r�Qm`�tR��΍*ʉ�0�����R�K��'-�@s|'ˮ�kק��ڭ��$<}ԟWX��g�Ljoh���Y����sx٢�q�L
��u2�ֽX�)�U����D��ZVȖ�m7�����V9iG�Nt�}�+�{�⍫9{�kc�6����Z>�#�h4�yC�Žr\�Zk�,VX���J��BD�.��76K��&	OO͔1=;�d���ECB�v��̖,�D�RWu�i��)��j̠�3�b�A~�����&�;-n,�nƵQ��X�d����aX[\��lT����*�=�Zދ��ZY�*�'q�)��ma=Z�]������)+�]���i%���yZV��Ԯ��F°�ܭM��0f�*ƺ2�(����n*O�,�x9�t�ͦ�#C>qUQ����=����&\N�v�j�Q% �.��*��m�Z���8P�'-f��yY��C�}{�����'�G��|��H]G���F���`^�06�J���F��γ�.�`}.'��`X3/���N`�-@Lt�kN+^���;���R��Ɩ��7�5��=\��B�Q��+֍Yv=��2�*����yW"hPih�ۀ��.�͟�+���fPǀ-��Wɦ+�'�Λl�L�lq���=���:�7+��]�I��]Է��"v���d��W-}Ǯ����vVs�{��{l����k�S�,R��ִ�����5;'�E��H,�q���Ȯ��Xɧ#|�Op���sx�>��.�d�����%Y�3+(v�]���k
���59X��q`Ӣ�Xz�fU�I�\f$w��)I���r�d���GXLC�.�D�B�$�G�е\��f2���b�Od�c5=F��A5����.�^]���j�'r�N�vU� ><}%��GV\3���Y^�������R���M
��ǻ���u�Ն>��ۛú�;�[���|j�v/���s��rwI��n��>�;^��c���xA ���&�(f��rbH��̲�����b
����jI����%�����(�����l���������*��X���""&d�02�	��"H��a��rr`�!����)��*��H$�h��ª2�Zb�f�&�*�����Ȉ* �����!&��H�"���(���,�hjd�J"�����*�����2���j&"&�2���&�s�j���K0rj(���*(���fJh"�&�3����(�����!�������B�����̂�������*�*��"���l�����j��(��)���) �*&�(2Ȫh*�"����Ɉ���(�"�)�����&"���&.v7)�k���m�ʑi�|)蜕`�F�,�Y�1������ռ�!��3���%xج�p�{3��As��<~������"�Y�Eu����
�b�1U�a���qǨI��Jn�����:���Wo�{[q6j�B�������/�z�r�����5�^9�\Ф�]o�e�J�w0��k#���&����}S�mrVJ�RP��{�g���z�>����E:=���xu~���d��x��Q�)ᏚSnkAH9�ޛ�o����xx��9���fu�S�U�*����"���)�b����@��9my謝r�s�*x�զ�߱P~�]��nܭ��?s\�j�.U�%�a�9�(t<e���CY8[ȓ/ss%d�v�(u�ݓy|��j��l��>��~��)׷b��Q�y����6�*�7��U�}F^��;����1`8����������l��.���M'g�ݳ�U��=5`��&D�]ާ�QM*�N��ռ�aj>�:X�8��/i����������:�t��1��@뫚+qP�B���Pݔ�^���έ�@��PIpG�[��`G6��u�����9mot��ֿu`��/*���X�\���U���O���C�_}_W�W��_M
DI��N��W:Y!��񇫎Uy�G�j�ȵմ/��[F{�=V֤�d�C�r���7A���t�Ϧ���yCN��U�(����ؽ���Aq9�O�:߹�>ޔ�qأ�.-x&�3�-5)l�*g%�q�5ّ��fТ�� ��.����v�+\]�Cv�<;�Z
>�s�Зz&�0�V2v3zu0-9�v����/w��3G�z��I��N���~E[Ϗ:�2/{������{�	8/}<�ݍ��z�+:�k�ژ���t�#;���:�䩜�ǯ����R��Ϡ�7�o�s�M/ݓ������v�`T�������u��o#ٴ뾑5��X�{rs�s��MŶ��0�l�qT�ʭE�5�7ٝ��������,r�zv�2sV%�g�q���w6Ѓ��F��Z��;�gf�����`��+��ǼNL�im=�Lڷmy��(#'b�a��Ĥ���V���.�#��.�Y���wL]}P��;��U�ܦ�s�3n��{:���pB�q�;q(���e�Um���m��5�+>ov1}����du:�������l�%(��Z��W�lu��؅Wy�ʩ��Ns\�4����3Ccb>�o���5u�_]���{�%��k5Ŧ������X�4�QB�}�{����8�9}r��0s�q�����u���p�S���й�J�}�O�αPrh��B/8l�'K�}󃞀�b��TLj��z����*�Ɂ��S���R�2�6�p���=#�dS{�]va�\���
?%�n��.ux�t*�/l��ϩB<+���y0�:��	�w��/I�Y1v5�
�PV��.;��?t[�(�I�27�p����{���y��kZ����"�k��p��2L`d�1� L���>�{«�����F��X��B��+˝x��;r�jfv�oV���Y���9��"�1��i��^A{�\�{��豴�UJ�+�b�*�͝�ںN=�vR���J.� B�ۈQ9o���p��K��X�S���i�{�7��l���C؈WR����W�tO�y|��7VQz@���u���������}����R�b��N��41�/LR������j>|^����:�0�~�$ք���iׄx�د���6�M�vm-1 ��WQk�_K5s:N��h���Ʃ�zA{z��5��T��/����?>�u���>43����[��G'�.(j��=޲&:��5����|z^�K��]]aN���z]��	��z[yZN��:�nZ]M[[��{�H����9L*��r�;���3"j�l]s���#��/AQ	\����v.�L����ڈ��Vf�"u�u,<����$���5q����q�uoX._�7{y��w+s�CƓޤ��	��: OU�pި�ln�V�짽�=�>�ʛ�
��ە�Xk�gJ��Vܒ�M�i�"M3�ʢע���&��b&7���ˆ�Go�㳘j�or9yAM�`���<�I.�����9�d�I�3��2æ�W]߲�i��YsЋ��P��b���B���bݨ���vT��G�z]rޜ��B=t"�'=0�"�"�W|��6;Sڻk�DDZǄ=�F��r�NE�N�jl��e��)ec�}��Jz8>Y���k((�\��{���]�g���꯮>j��$��S��toԚ�S�����d�j���ϵ� L]]�˃ȍ�t�z��Ri��|q}�V[&(,���X+��	�,�_qO��=�߸kа'%{�%�v���dR�sWQ@y����y��o{!�g�]��#`���}���t��Nz�E��۹��Oym�,>�U�G���96��ֱ��˺��@\��}��_M\.$�ګ�iW���ַ%����vΧ�����p�se��u:g���{�١�
b��m���b��Z�ר���w*��*�o����=.��6+�|��f[�M��2;��>^�R����/��\�]�|hc��j�eH:��:���x{�&r�j����뛋m�ҟ�s��1�cƬ����4wQ�ޜ�����t^o�����BC�s^����:�f��B��j{3�3\���[Ț�g�����-�3�`�w��]���2�w�A��(ةO/����C�X^&�	EaU��L����V��-�Ѕ��x���[�s�&N��L͍_vc�<�j�ҭR
�͝[������[���U�}�=߮���PN�~F6�3"p�k��gZ�;ݜpE�� Z��$u�\sJ���3|���)�gn|z����o*xc72i����Z�n�RE2�g�1� �3�J>�E�M)��
{����v��̰�'`����`��*y�kzL����c��0�{��統�Mo�w�O7�� gi��2���\�O<d�V�+�3{UҖHD/���6�%���B��5P�s��Ŝ�[9i�϶���.:ڧ�5ҷ&�·�k��W8�|e���B��6E�{�>o7JY(v�>ޔ����/l���g>Qmنf�Z&���>���F�����JE�p"�v(�;V�r�����vos5*����t��x[V�gñ�N_��^�	��ꅵg�)WQ����$^�
<ePo����<�~>P�<-��l�9��=sm�=~
�&�n�Һ�]��Փ���u����<��댞� l�����x/��sk^�i����I�l�=LaV�v?tvh6=�ߵYA���8�折5:i�VMXo>�;Va�S�o�U\�!�HK�)G,J�۲���^�?_}��}�U/f�Ȧ��w�_s^�l�w=���)�X
���`�N�����yp57N��K�m�v`���:as�M/݃��ژ��t��_�Z�_-����$��z�ͫ�����mI絿79��__�qm������>�}|���^W�V��^r��d�3�~�̜�7��3u��8����U��(��d�ftuwӻ������hs�/���g�rmry��gz4m)��|/E,�Lܜ��íxN�DXr�_�k�5gTͥ�r�]�Y��N�׼v�ož(�Qg!�tx�SEL4Ë����.�ǸU�	k�l�=�6c�w<T��p�'����#Z�e���S���.���HL�Rk7�eLĺ��ι���#��L��5�'����kk�ʾ�xϽ��4n���F#絻.�s�����΃hze�Z]�&^���2�ټ�Ӑ��s|�;c��ּ�L��g�z�]hcjS�����Qe'�Q�����5]�m<;P�Z�;�6	�%�v�6f���V�C}V������W�X��6V]����3n8֋��4��Fξ��q����s����������_�9?��e\��X�f�c��j��zU�q�p��/=��u�p�i��KT��^��	�� c��M�~=�-�
ȶv!�׳C��oG�돴�znrryF_���Fm�[�__S�tmS��s왇{�:[�<�[��rP�tǺ+N�#^Y{��WL��LyGrC=�����U�K����!��ѧ$֪����i
}xG�)�~���w�_�黪�0����tv���t6�So��9 �>������1����&��⯳�Ov���ǟE�Լ��>��xs��ywM���Ӿ�u͉���z�1b�ʧ.�p=�S�x��M�|�#:,橝;Вݙ�4_m��r��S{r��r��3"w��<Py����=ҭ�2.٬��;��f��9�K��+��I�篋(�G�G*�����,S!u��Q��h;Q��N9Hy��F�WJ���T��][��'TF��/��kb����}+{NW
�K=v�[b���*֦J��kU`�S��-�%̗׮qr����݄ǽ�tIQWQ�8һ%:���ͨ��E3O�꯾���qKSR�_w��ӗ*��>�p#3 �a�>��X}N�k�F�w�^W�f�{ػp��pm�[�u�xc?\ɦJ�Aɳ¢���=�]�hK�'�e�C���)o�
���!1�$��f�c��5O�N��w�;�jF1��O����/=(�L1D�)){��߃ʏ�j̻;�P���+_���i��Q��Z�5���N���<�����5�^�3�)L�m�q�ԗ�sۛ����Q��b9���z��H���,��rS�&,��~��?�7\�K�{0�\�ͧ*�_�b��yF�>7�-��_���ϗ�|���ysP�R%���G��|`i�s�/ӷeY�/P�K���-+���������ޡ�M�y�>2�ޢ<�ש�Hge�>�L��c�h_S��i���\^
�x�pM��sܼ̃������mx�/�E�^�΁��ϰ��﯅_�ȑ��R%�nn�`�ԛC���>�dӓ[ܭ�.��G�Z�wD�OwoM�G��4�.:��=��{�f� hn,��7o��H��vX��w����	&��d�	b��i��֊���3�+��Q���6����wS�y�3AW��e�'`�ء�_4�5g@�4`�Ʒ��N\2/?W�UUW�O�Z���I�n�}�v�e45q��du't�lϮ�<o4�y�3|'b1����/��"��OO:�}���
,���C�ƞ���n��*�0�\k����a"9�.�'\��(��=6�������9���kC�j��L�;�G� ��a�M)�$ŷ���G[��c��b�g��}�ґ?'��P��tx	�˗cms�d�ܤ��Lt�C�Ud�6yMy�k>TpRxk5���/�Y\֌�WgO.��,��,�9��*�Y߶V�n3��m��+5���u3ٝMT�u�x�ڙ���*%S; P�ZW�|f�����ry�w^�5��p
סi-r��*���ja�,�¾��G�r��@S9K<�9WL���/o�
�N5�>�.�Z�hM+���O��|�x�2�͊qw�5��X'�j�����W,	@;�Z���`�
z��|����0ץji��o���m��0�Wq��pc������m03y�
��Ȱ��:a:gg]���!�0G�"��/]��gp2��v�c7Ԯ�˕	3v���9%+��!5a�Wot�0��t���8dU�bD�,�Wnj��<ۮ.!y�>�w[Ө��d�\v]lW�����@�"��}��فu�ǖ�.n�s�Dq;�|Ցo*`�m��H�yD�v�ԧR���`��r�d�xm#��@u�ȢtI��[�{W\;q��T�tH�����X���5�c��;�GdT2���e
���������vo�赿@�i��Dsw��ĕI�^���K�X7�y}cN��[X�}���m(+G`�hŵ��;9���/��;��5�T5ѣ��cC�"��A��ھ�_vXۅ�rr�o�sV�ʱԏpx[ɠNt��i�hX�VpW�goS��:[�<�}yܡ�ɉ�Xy���Z��n+F�]d�ȞL��8b�����,�f��f�#*�&4!%�a�iut�1Ϋuy��z¤�4x��xl*+i�܀vp:�X� �~W�7)���;IY	pg=�_6xl� ��r�y�jHs C��M��R�+�QɁm��U�cqf�+*��I<�sK����۩ڱo_^��Ĺ�ĜmG�nAPe`��#�:ޤ�B���,�o7��nh ttr�],_hH�R5��m<�W	�=NII$B$1g޳x����i.+���/�+�P�Ee��C
D�!�^����v�v�(#}[g��4E�PQ5+%�J�@h,�9*!X-��OC�Lr�8!�Y�.[?o�I��R������WE9J7o���ޫ�V1v��S�Ӻ�i�yA�w}7wr'{d��ݸ�9Y,^ߵ<E��	b���6�Zn��ך����6�w+�c�s�%sq� ���>]�h̰��Q���N��r��-�CwΠ��Z�Ԯ r���,X���&�2b�)m�ե��9���3rU���v���¡f�fQ�P��q���L��:u{����a�Y&͎��`m�QDs,�t�N�"�j<��E�q�OR��M�Y�2@�f3o:K����R���uح���U����B��ٰ9�}��{���/����mU�4�;�'u�\�,�W[�Rq����G��l�
�fe�4ˡZ#`� �SN�$�@s\w�x:M��a�qUX!Y6-�Ce.i�(�6r�q^�b�⮺R�n��\�+�g[���+�%ī������u�RrŨ��,ΏF+�:���T̞�Z�l�'`�n�-���<Ԑ��x��^���V�~ؠ�Y�-՜}�U�3�Z�lpO&��ݧtd�D��?�Ep�Sv��Fnn&BԦ��қ�7��lfL�@��P7{@�\+�Lu6���H�0�H�4�9r�rw\9�e��z�H�&kqG
�e�X�OhE)���H�5B��cL�)+&wE��Q������Z��_9��VR���IPB�ޏ�+���r�7�������������b( <�����ɉ*�i&b&� �(�$�*����&��)�Ɋa��
(�f�����&�)�&��*Z�"&H�Z��)��
	�X���3)�#&'1�i����)�f)���e�
���$�i������* �3((*��"�h����!���
 �b��H**�b�
� ��,(�f
����I����f*���jji���0ƪ��(�2r,̒*(��"b
*�$�3b�"���f	��Zh���+3$�bR��("J"�b*" ����"�**��&i*&�(����j���jL�*�J��i��̌�2L"&���
,�k'(�1���J�
���(h���h��3)��)��Ɔ"�(��"�!�,��
##	�"���
��"*"**h�,���
��*����!���b����*��{&���kR��M)Hd�u"�d�D�u�h�k�#��������t��*1�w՛���wmS�
�k���鼑��� >��F����t��c���u�[�=*�y]n��H�p�xҘ� 
��[�~P�һ~�|A�Z�ӱ�4����<2��p������V;����\= �E1����7]n����k��:E�p\��=�6��v��y]H�3����J���)���iy���7Z�\]CG84�Q�T�>�nJ��O`񙪯�R�t9_�!}[�¼�ʅew��z�?4Xײ�*[v���<pMv�=.�7�a��3�m�6�,2����]R\i�WG{TTy(�yj�ۈ���|��N+�ޝ���*�WR�o�苴}��[�����;�z�AuDu��⬇���i������N4��V7���b��=�W�]��7o����
��YA2��y�P�B�u���Іd為e�:�-0�.C1%3Yƥ(�۝�z-4/�^��m4���P�e������x��v׻Xpק<W��d��vC��u�I���w�S��a(t5�_Ԟ�T:���01'��8幾34�M��R�Jn����S���q}ȷdtdwՊ�$�[�����tʻ�@u�GMǗ�I{1N�)p^��z�M6h+��Ѽ/!sh�����Έ)������-�36�J��A�����!#��|_�l�Z�|>��ժOt�uމ�tr���Cz�<�vVY,����-)�SW^]��Ǵ�2g�8){��׉o���`��0���|�����B�y�a�V��D#~�������9{����3����gޭ]Y��$��u�f0q�-h��``cѯ	�ڳ�;��}�%�r��[-����]Ժ��\�ʾ_<z=f����pXRP`��V5�xt��^;i^?x�MT���d×�����1~?;�\+^���'�J8,y����^�E��vN�m���&�ld�]�^�#�僞��f�j����V��N?|}�=Է�44+s;�q!
]�����1����u����*�s�@��𜂷��wY�����u-ߔڽ���lg,��Vӵ��z��=t�}����Pi����`;&j���NoWR[rE~ݧ9�VO�X���s2ҟ�2(u�&C��4U�}�Q�����wԐ:���=�%��rɫ�d�<[+�Ҋ���L�z�8�:׌�K��0Af�,�{ƶ��)f��^VV�TcC�f�n���SAWVd�v���� ���Y[d߲sB1E�B:�9����{vj�'5r�:�c��n�];}K���i�����2�͕B�Y4�v�Ak���P���.`�W��| �=���g�t{�r��I�`��/*��\�/*�H��t�|�.�9�jeNyYK=���w #7��%�O���H��u(�iv������exq{:���|���;�>))^}@^[�V�L�<*�!�Ƨ�;��_$�L�v2��9]S�".$[����c�{��>�^�%_�9�%�,����u�L6�+&��$���������U*���u3�y֣���oVJw��U��~Y<[�.2�T2/"j�}e��n[�TE�3Q\�VP�=U.e�L|s��/n^������jL��G�N�P��|҇�m�V��o�u�}��#��^Z):K�Yb�?��k�i+=/�`�H�"���#�G���kf���cވ����8	�]J����"�_�"̥�)�f� ��sV�]�.��ی��\��Bd��NG=x+>�Z���WR���7�O.7Zm���=��6�L���f��n��נ��n��1=K:Y"��f��Na����O.����>���]c�V{����7ׯ&��4���Ɉ�ci��M�����Tq�H�3 �%6�!iZ\�N�ð\]����(VX�\��qD �v�X_C�2�*Wa���9;�'	�L{ռP���T�^r�ø�Ox�����7�J)�o�c�{b���t�ب��q�������ٯ�����m-N���c�g�@|ly�i�rZ�r��X�^L���e��w�&�9��w�e�o��D���P�pW��
�=�P��:�uv=�=ভ���G	��_!��%2=K��~1r�]N`*���"� 5Z��o9]t\��� �z�� ����e�Y��v�-��L�p��c=),	����H�Φ�Ƿ�{a�W���*�̹5��z�.�h>+5@�gҞe45q���$�Cg��M+�g����)�gz�1��3z'h��g>Nv3�ƞ��{t^}*�0�\k����$s^�v9��!|a[5�Vf�����5Ћ��N�=2���3��e8��a�M��x�-hμ�&�v�/����y���ϋHd�����Q��v�X9��eB2�L������>��@��x����n��T��D��R��,B�:��F�3֘USq�3;�@���V٪����d����Y��G��F�Q�Fr�~�`�����p��P%к�o�L��u�`˸y������N�FISk̋�ߢ���f`�;+;��v�D��QRk�WQ�}���� �o�v�B���
}k{�:&�%����Ԗ2�T]��`PY�eI�ٛaL����-OR���䐼���dhu�{�B캉g��G�q�7�u�ET:�"��sb��}�U}_{nl]p�[�>ڿ�q��B�~AN���]R��7ᮭL<'�ha_]�F3�^jR��=���v�����\D�1OQ�;r��Z�hO�WyX��h? �X�tKpL��`u0z�B�kK�y�n��ް��d��i�8)�X:Y��(��k��Cm?�᷉��yb7�C�9����T��Z��`�:����fx۽��lN\E��Ԯo��:rV������C�vL�}ZrX����g�_>ͺ҅#I���򘧹/E�:����Aq�힏;wh���.|j��|�zVG��1>"UZ����_t��w�n���բ.IKzg�ɧ�/Y��Uh��xr�:��ئ�������x�O)�O^��<
E^��<�v�6*o�G���d��M�ӂ{��R�B�t9]B�\^Aug5��ږ������>S�e��w9C����Mv�=.�7�a,�}�Zϥ"�E9�l	�� 3}��6
t����E�qm���9|ק�ݟN�xO���	��t��s��}���;��͙�P�a#�S����˩�{�=ˑ�;�-Jl�dA�������H��ލe����_\����#��nF���z�U(N��Z�����:��Q�&�[M%r�w�ET=:��ዳ ]|��O!z2@��us��{!$���.w꯫���1�!�=��@��]Q��|U�C��c�MX~}�p�ÝX�3��l;�{Gwq�4ʍ�}�ȴ��y���fX�v^U��C���K��9��P�皼S��t����T碝[�Q�]�߮��(�Z���3/즔���x�t�w;�3ٙq��zp�
Ce��#���\OYM�>x!/�"�C\�/Wo�)����P�Υ�w]�-��9=�]�h���O��*����O�f�.�/�K8�$P�K��Jj�˰�C��}/r�{=A�t��7w��4�gZ\��a}Y�|]�����B�wf �U�e���� w�8\�\c�ї�{.my�|���K7�	�v��>�����Ne�m9�j�����J� 6K�k};;���[o{���:$a��R�]��6��9�t���±%����U�S�5o:�C��%���5��3����= Q����
ϙ�{������(�ň���sd��k���b�UP�ysJ���ygMx+6nV�,աJt�^��R�{U3,�" ��D��i��.P]�<ti�.�Q�պS2%B�o���;�w�A��l��dYj�$�1����`�2�Sd��N�	�VS2�n�m�����`�%�V)}�r�Z�$�n�G�u��\I�5F�!��V�} HnB�m��_W��}y���"�?���mY�;�����l{��$֫����O	����tg���d�ߒ�;��)��]�	��h���P�b>�r��~��tx��3��@]�����O)^�Xi���XO �c%��]Y�V�fC��ޡ"���L��9ȫw������}��O��}���Ϫ��,��	6.-��=���@�w�Ҹ���\~��F�2�/s������]�n��8���y1������'�5�K��}���xė?=>k٣��5�
�����ޫ�"�(�a.�0}J��N�:*S��)��[x��z�l2���ˋ]����'j �?�z��N̠E���h$�L�C�S�*��=��eWU�E����!F\��ٷ�s��5P����Y4�]ܱSW����"M�؏!��nOzN�ٛ�w���v�Ù��3�ug�N�נJ�!��P�(ӵ�yp�u���y$G�mӥ),�nX�7��d�/
�]
ъ��]��V�)��4�fR��L��F�;�����f���qu��A,����t.-�L�Q�T��=��M�Z���^ՈX|,,�BM�*��'��f�iВWE5|����>���g��Y���M2�5$��[�2;˥��Ϸ6����Y&�H��W=���p'wb����mݝ������>D��QKΏ�Vνt��H�������V|^��xm������~��D����������VQ#A|�/�k�`�km�>�=e���^%P���w~d_���jõ�L�<��d�ߥvWO]�b�&�Q>���7+P�b��D�n��φ������͓��Y ��ydu�J�뀣c�<DKO�h�d���4�Y��5�Yx��K�u^}Wj�Ȟ����c�M��ӟym�3���5�@|}:�-r�M�մ��tk>\��X<�����'���w�����K��.�t	V~^ۧB�
��YКK�߼c� g�˓+��~�eS];��L��=��q�c!�V�y���x�W�r��,�g��:s"���@��Q�b\�GϻM"!=�.*�e����֠-R�R���)�|�H�u"X&�"��o����$�v�+��8T��as��-D!��oަ�Ƈ��ԝ�)Pق����I�%.+��=t���sӦ"�%�0�	��}8��^�n��VQ���\'Es�Eo�V�xݕ)��U����h�˃ZH<�w�����f ��-턑.T:���{BS.��bq��Ա�V��ږ(f�ee;�W�n]�����^T�Yѹ4����O;{/#v�Fm#��׌{.�[������%c�v4��ji�gP2>�ﾪ���u%6z+;C��x'�檜}r���	�7�8i��;�G��TN�)4{<��ԔV:�{S]<�OY�4�[H;Ｓ�m=Z{�99��g\#��3bϜ�l��%��m4�ѵ<zG*�f�UJQ+���������^�hw\wt^�1KBΛ�5�xk�[��fJ\����f���ď�@��RK^Z9�o�]��ZM�Xx{5r������z=*f��k�����'Q�E�����Z��+���]$5��&��wp��Vjg<��=ULգ�ザ>��#z���][D��
z��h�DCX���v-���T�+|��3	�=�WkJy���;�-�����~���৩g�,��+�p:��LG�U��"���Y����'�}�%�s���f<�Z}H{҇��Ņ~s 9ueO�{^��=�8s2���]�Np��C�#����q�mz�۸f�R������ǵN�'�u�,�3�D�_�w~1s`�&���wYq�ѤU2��p����Vm��#B�~�Ҭ�:߮�r l�u�� ��wQ�"K.<��Ȟg=+n��o%4��-=d旦��=ķ4��g��IS�lP�V)ʉU#ܶ��W�Yĺyjm���|�������>*q'����r�f87|�\M#ư)>�^��},%��9�y���|>��|�og�*"=�p���|&��{�ĺ:)�¬���y�e���q,l'=W^�_n�}�[[{*��m*�b����G٦d��MU��3�҅��*ʱpw�t����� XFM>]W>}�߽��uSw������z2\/�.o�Á3L�[JL���-�E
wwQ�\5�ݡD.z|��U�.��{��mNP����'�ݓ��r�����a�PD�n�zOb}���5���VE�UT3��T��8��؏�_lbU��3����$�ܹ�-���w��,��5�X���PL��v^U�]2��2s𫔨9	p�م;�X�Y���?{���fZ��~��@�ܚ\�\^}B���Ҙ��(;�~}� T��޻�ԏr�>�j�ԯ=�W֩�OYUg�늽PM꺯��Rz��hʉB��I���:y�]�NU�O;>���6*_x�.2�M`yp쬲Y#bZS�5u�;N<}����Uv�ע�zt��(�{|>�c�,�x����;ʜ��~�R�`�兑�����쭦ԲUyR���M���"7w��1ܝ^�v�-��3LK��8�j����nt"�Cz�C�R���X��z][�e8n_vG-��|��e�h��=Hђ�xfm96�("�.,'�%�n\�}��j�y ��5#o#qne9�e�uhʰ �o�D��&t�擮��k��Q=�N��;�Z����:6f�]�=�m�j�]Υ����jV6����7�i��7�����u 5�o: �**�D��mȀ���X�r����0u4lP�]�����ߢ�ir�r�yO���0��Y%O2��+���¨���2p�U���mB���)G3 3��K�[�t��e����s@��:Ĝ}���z{hk��]��Uۗ�I������`?�S��S
���)#�q8�*e��2���F2�d�eU�$ض+d�]���wc���#؜���9d�J��'d�-βKH�n8өٷ;�T��2�J�hBwH��M�����53�z:��5G���]�V��Q���� _u �P��ֳ7#�ff��kv�c��U�ׇ&���m�u h��3�N�0��]���E�n-LP�8��S�755�iW�ks��;L�VV��� �Y�,)�6kw�h�Y�A�]��Y�b��/l�)�5�S��H��q>��M��L���Z�^��@'t�t�"�j���K���z&���(Į��jE݇�7�eFc�f�Pf��d�O��*+���p�1bk�b�p*-팁e����]>������jN[�=�?m9L_S�o6�-�K���4-�<��2�e��x�>���ʬ�����"���λ,kv��hk��b���ȩ�v���y�Uԍ>��sb����_d7��n��\tq܆!Sx=R�u���f&=�Iݐ�7}GS�X�+[��2k@�ԋ����^C�kKܸu7}dxvYα5f6�L�Tՠw��x��i�B���N���+�=�e������v�
��`��V��գ[oqƠz��VҐ����5��v��Q�$�9tC��M�,C���u{ظ冝U��+����I>A΂�X�@'��-���u�����}�o���FV;����\Z5���} T��B���!��ӎ+uۥ���-bs\)n�Εe:�*v2����w:���ؽ�^Y&��Q.=S� ;�CwDM�]��۫�ݴ��`��K��Tkt�rk��ᱰ�\�;sf�b۾��nw/VQ��v͌_�[rm�)�bR��d/;�2H�=n���Jl�~�{��&�
AҨ�9�{Ar��F���U�����e=;Af�-'�:�ҏ
�=��h�nR��p���.�=�}�^4TZ���*ek�w��%�o6��p��(��0i�.�V������Q�}x�frM�s�����F�|m��jj�s
 -��w.tgC�!�ZV�+#��Ww�_�,}4-UMT�cA�UTMU�SP�ESK1A1��Uf6aEUM1ST����MT4UEMEUQ9@MaL�DVA�E9%�QEM�f8͆Q55DUTMU0�CDM�EL@L�T�Y�R�X@0��U14DDCEES��5��MMEAVND%DD�TVf%QfeddADD�Y�Q��$C$�ESEMU�LSIEUAQMPMY$�$PMMPEE4D��AE�KL�IQQE5�aAMTE$�,�SER�T�D�4�T,TR�Ց�TTUS�IULSADLYaUD5T4L�#RDQQdcRT���UDIRMT�NSSDIQS�y���־/=(�Kx��*R��\���m[::�>ԻN����:���k�����u#i�Q%7�*^��������G���-�L+�ۆ�z�׵汏a{,$��B)˶���a�'J(�1�g�?oy��>�n�L[�>D�:Y�^��߳7<_���P�t���*��
ut�J��A��3X+���˦�\�Q�cg�(�k�yL�'ڋ__�c)Z�</����TpX�~��Y�8��g�{}��*Gl�/�[Һ/j��Of�j��/j���8)[VG�H���wj�eü�v��m��Pa_�b՚N3�P�%��<���Z����P>��=0#��\��Cj�'���ZgmC�`uY�[�C��[5��s�y�ĺ�Cڭ���e���M�YJ���?b�ӡ�e��_���L�W�p�|�ع���9�	{^��\���e��:����$�wv3�/���;�E�����|����W�	7�.-���(���&-��Kh�����^�X��`�6ߥ��Dt|@�v����R+GJ~lt�/q"����MMV��ۗ� ���e��k�u�RP�(`�k���=V}*Ȅ��п��>���ҩ�g�^]d�o�L\��sM]?Wb%d�u8�z/�{�i��R"{��P��j-��Mqi�x������C��� ���o}�l�R��9Cۻ�Dk,Я3du���If��9�+�D.D���q���ى�3�+� ���E����8������{�a�N}l���z�nq��<����(;S����̠E�GI=^��V�7o�\�E��]�x��	Y3��<�^�����Ns9g��TCD�r���e��D W���g3�6h��$W�i�ם{�>���|t��-��-ɗ���p�,+������>� /�P��72]Lu�������m��3��:���~�,yU�u�����;c���)X+��]$�y�O��X�e��/PO�9�i�ꋽ�)g�:�M�I'y��
j,��0GD��^sقx��(q���/-��7S.�
c�ð�#�_���[��բ�v�*�Pm8)�lt˴>�5����T_:�^��̖nM`���{S�=�*��.��I�TC?:�J�뀣����ORΖH�L�L��3-<��Ǥ�Y�lƯ�e䏆t�g_%+~�t
�W�zQR�wày�i`���ݵ�7�J⏟L2��s۫h[��d��pB�yi�5��R�u�۸}�1W�sK���u@��������X��v�Y�vՊv*�G����K�r�T4�����\��ΗVOr����K�qyHZ�4�)�Z�LU���VL�[���[�7ۏL���~X�Xo4��y~�U��I5�����V��8s�w�I�x�kh����_6�:�[`�P��1å�>�����ק�E�6�W��)�7��y`3�O�GZ��V�t���v"��וǣI��]�S���|������(A�H�>��Aqu���$O���QҒz���p���H��cg���h{�ƞ���ws�~�40�ԝ�67�38S�&j����ɳi2z;���я%�0�s��}8��^�n��*�0��\��=�٥�[��88�{��@�����a����2�vᮮ��(o,��L�};�G�ج�U'	^���g�f�7M�� b�UaZ�*\�H?T��Ϻ������(��:��Bk���k/���0.mo��;.��)4��k(&E�A����U�w�5�̷[�o�d]o�rT��̡8$�4���y��B̙Ou�Xx���E���qw�p���.��%�`jfoSNuPw���7Uc}��맙����p��fZ�pL�E�+��U$=��%t댺�||��Ѳ��^Us��jZ������,�T�.�E�a��ȇ/X�z���y��mn	h����l�v�x��L��j���E���Ȅ��Ԫ,A ��fve�y��p�:�S��ћxz/wٽq<�ҥ �d���ʎ���WV��U4�b<��!���*��V,��{ �'L��W0ķ���M\S�G?��U<'�߷{�PC.��X*L͔K����y��)�X:Y;r�ه�X�Y����Ş༼}�Оf��nə��w��6�n���,+��"�ά���k������O@�k[�ܮ��G�C�ګL�ͻ�{�ϟV���ǽ;3��+�m5�<XX(̵��{J�f����O�f�"�����YU1>"U���ǻS�M��N��ƷΤ���}�mg��̡���\^�j�cf�Z����L�*�Ğ�[�=C�YV���$G=.o%f��;�WW��a�t�z;��FJ��"4�b��_V{G�W�Wx��f��%�$&ۊ���-c��'�sƫ6����P�9c�&�z�����0�f�lT���=�n�n^EYy�Nk�s��c�����1,<�Z�fڜ�.W4��W�~�*Q�j�]J��ѻ�\����֛1JQ*�Uq�>��:��'���f�?e	��z=�,9�ۊe�s�>�dob���e5��,X)����1ݗ�C�N�z��D�uwr��[&�t669];�7!�^)o��-�;r�`q�L�ܩ.��ǚ�Ṿ� s��Z�]��Y�d`u�v
�9��@]���=j��۽~���+�d��d���1;Q���F�+�t�^1�z�w}7b�����ȡ�_UW�zt�=��C��o���bu"����M.���
fbiM\G���\��&��y�����7� �gӞ+�QBzʨ�>?U�^�����+�Rz��;��A�y�c�a�C�I�y�u���A���1[�]LZ}7���}�_��D�H�J�W^T�u+���j+�nZ9�bC�-���c����Ǝ|�z �e����:0J�������4��]�t����=���b��������Rft�K�s�3�ʏ��m�Mu=1-s#sJŘ�=�@T���k�����({�ZJ���}�3�1A%;�Z_5��5|��@8-�|���?pV��@^����J���C���5��+�˫Շ�ni��i�9>ۄ��[$�~:�)�p�ư�?3�m�����W,����[ �e���ɄT�Xb|++���3�<G��n�}i�5��UӞe��Η˙V��1賹ass�����P�v��=~�/+���'���w��㺣��n�x��˕On�/ۚ�!H��FS�Õ��XI�<�]���ox��:[�l"yK�Wʠ.s�]�I���r��Ǡ)Yp��X3�5�����]���Yn�����kbn��1�vs��w�k(��Y��K���u��Af��c���9�"�+zB��?�����7)�����}��j%��
�8y��;��lBe���=�I�k�Q�4��
^-ܘS�ܤ������4�����3%���ɡ}P���es�QY��OLgMQ����}^���헕Y��C�xȴʔ9TN��b��DV�����I{�ƺ�j.ˀ�S�����~�����X]	Ά	ƻz��*"%�m.�\^�t�2'xIg�T7��*�6��r��#3��F_��8�Ǔ��� �?�z���idp4��9�~�gm�oݛ�{�h����x�N��R�׿J�?[��Y���TC����劚�.�[�}꬇��ŏ�е8�5U��|E�g�ЙվZ:�ïD���(f��J���#�6���%���`�O�GD߫�R�du/���l;��gK;��S
k�m���f��з<-��E���yF։���\1eR];��^Z):K��ŎuQx�Vg2L�m��|z�3/\�S�>���˪��]��[t�8�~V*Wo��j��m�N��B����vH���'e��mo��}��hτO�l���Y��}�h���u;8,"Fs2�Bi�:�AːY.&8i{�f�z*��Cyv����9غ��m�N�����Q�:�(ol�%���N�&)B�J��{3jL�Ǚ��W�w�����W�V��9�*����B4M��I�:Q>�����o�H��r��-/W���lT�c�ۘ}-l��с��<�jrg�o��F���p��X:Y"��n
<��b�k	�R5�S����8L@`�}�sMLJ��#�`�c�v����.Y)�յ�mU��+k:3����/ۏ�n�F7���1<��a.yxLK�2�
�t���КJ�K~���阌'���1�y͖;���F��b�Y>fgW,�`/��x�V�x խ(z�ܿ�=�>{�\ױ��w5B]�q֝�[��)�"��U/=�]AS��$:R��3�[g��=Uv���":��x����W6Z�����D���¬��̳c{�׽��#Fμ�$�i���Գ�綋�CŘ����ƞ���n��VQ���\D�����1N�Z~�-��DdV.]��S�K�3=6х��ٓ(o,p�=���x��N��cHޚ�g5��>�D��&�,���!��˩u/��uSi��{�99����f�
�]�|�G�׶�[s������c�ݎ]�0o���`f���kY�����^�P���%o��<��J;�ٷ�&�"����u٦�De*���k�K}����@u����u�9�F�쳻�B#��s�#��Yu���{��Z�|�UÓ���M+����A2/���Z�=���u�a����p��{�3�홧�z��L�ʘ�_���nP6�ZJ..��{��rXgU\��L�ý�W?c-�%0�����z\ڳP�S
��]$,k5�&��۸{���I��\�6t�5o{�v}N�3�'������4o�=D��K�"�G
�"��F+���F�j"Mg�\����KsH��V=�"��Z`��Z:Y;J�f3%��W�=��wt��{ܼ�@赛�\O2��'�x*a���m0���9�agT�G[����)浏��7�������f�zW!P�ً)���M\U��Ҭ�ͺ҅ V<(o�������Y�W�.�[���C�_=�\5R��c�Y1>"U��Q�a�\���N���g{�'�[r��PzI������E�Zpl��Vpx."�#���C�WY;�Moj��<�e��{�rU���9�}���g����d�z*�5N�`�A���k��c��
�Ur�n��q5v�j�P���m����x��Ǵr�٘��V��v{��\�o8���h�n��b�x��D�y���}��5�8��X>�����&�<��j6�`���]��bS22S;���������lK��I_-��ol���j�7N�?�P"��+˪�V�e�w9C����]�Or\/���<�	��Y~S6��^	a�Zh���(u�bU�.i�{��mNR����:���h3P��}*�����l�^�eo����.F�*�*���uD<���
�Fi0���R�}�;Kuw:Z����y�����N��72���"ŀS=PL��vZC� �t�PYP��$~��C��,ƙ����|��av��Ԉv&�P<Z\�\^P���x����W"f�Z2%9�u/Ա�^�\?zs�}j�(OYQ|n ���"�C\��OWghŚ�/�]U�;퓭�y:�{���ꓷ�e��.�->3z����%�3ȑ���ٛ��?0��-����iݩ�f���R�wK�G>n�~]�^
����V�;�Ku��5r*�ϙ��t����j�o��WJ�TY��ٸz�J��K��S�|�ʻ�O��i���Rr�P=�3�+��gר
�P��k���,vG�kw̓G��#�V&^�w�1vN;���90��me�؅T��R��h,�W��h�Z�n�ח���S#�
r���@(Cava|���9^���em�J��g}p0a�tc}#`[2�+�wS5���Φz_^�n;���m��x:�9���n�����X֥�yX�r!*��6}+P��_K�*����A�w���Of'q�o6��R�������$[�oJ�J�Y�^
͛���|�&7��W,fô�^�����ǹ�����^&?R�f�,O��Ћ�Uv=�[�|�Z���km�c{0���є�;�c�����J�t�� �[9����q=Y����~;�����=�M��nvnc0�/�c;>K��R�z��c5;���]ë��X�m��{<�#w<ϼ�<��P7ݽ�/}�E_@00�I-1�rɡ}P�c�z�^)��e˞]�É��a̮�\��.��u�"��V�%�Y�uYy�*��������W}O�(��^��j���=�͋��G��w�d�9��'�����U���\��j�J���v3x��F}�'<��b�ו�*Wy��m�ז��U��L�<'!�Ƨ�t-�p/��uu������zg?z�\�v2��+�šԸu�|~�9�d����1׉0��d�vI�Go<V���!��V_W&�}Y�� �� aU��$v0~�$����E1s/�vQ.���n�CW������j.
��rfT�����sYI�æwb������o'�N�fXYs����wiJ��=����c����}�pg4n��P���Ĥ�m�����.���mзVA���'&K�I���ϻ��T�.^44V�]%3K�]w�~F�0�o��g*P�W%�o����ҖqpXrƋõJ�筻�㾮��B�Y���R�/���S��n�£��VNW�9��]N�Ӣp����M*KLX�z��A`�w����j�2�f�(��¡bv�q�1��i�7K�ă�ЙJ�8�j���ox9N��sM%t��Y������o��xL�=gpd��W��V�uho��\��D4`�*�L֐``2�qGD����K.���K(�!��zVL��s��@)�����!����zoYj�-EH�ͽ� �x*��ޚ�oc>B�j��W�WNe����`�Gka3qm*��̎�n�@��Z��8�����(�[wH���U���{r:�qY�Π�5�6��[5�Yl70����3�,����^оws]�cj�D����'GC/5J�Q7ݎ�x@z�ϱn�x���i��r�kH�1��2�[��'g+���,��?q]m���j�V����t��M<�;畊�d��d��4[�n݋u��f��u�o/�pbNǲ�����.��`0�1.��t9�������t������6�;[n���V�T!m�si�v��nc��8�I"($>�p��զU6]e.�i�/��q�M�z�F=�kT�M��ԩtr�E��c���!���ݎ���`6�v�N`=���K��uy�!z�1�"�T�tL]�k&��B�s�1��(�caǧ���o�!�~"�C췆��2�]�C�N��W�`��D�J��%p�����Q�-"��=CF�ޭ�4�Į�ܭ�@Վv����O;�K��7��V��
�+Z�:+�Xkm��n�{�v��5�竺0+Ș�wu��%�v.i�
��J��ԇ��]�V�;�j,�ҷy�D;���烴=+1�U{����*r�����*���*q�~�n'�$M�Z�[X
|�Ow
�3G]�hTK�=#0�ꆛ���m��i%lØ�k��*ܫ,X�����.��f�r�8u��*I���-6{�6��n^��-�bK5��o�{����6��7���x	4�6N�N�l��q\˻��p�\��ppg�ة�v�kkQ���`�uu�����l�]��q37������Ǘ�&���GS[���S�1����8�h�}���՛��O����.���8�4���R��Ì0��/>ͽn�oU_Q؁���a��z���i�Toj ��O��W�1t�������ghB�v�?{��4TE%QQ�SQD�T���AMDQES1ETA�R�155L�SUESUL�4�E,�D�QQfcSE1QAT�RQ@E%AQ5ETM$E!5UQ%1�LNa�EKESQ`DEPTQTTUQ4�TTQDY&DE�D�Q$U�faL�5TLUATFYRDUTT���S3�PTADQQ0ME$�DUS�Y�U4�13UUQTU5QQMATUASMӑ��ALD�0CUTSSSUDTTAQ5S�D�)DELQTT�N`eEUTAE1RCTP�-�UDETQ,TEEQQ��ETQ4DL�IERQUQDUIMTM1AQ�ddPQS��EU$IDIPE1UE51T�MQD�1RIYd��CbEDTY8�DQ4LKS�SUT���ELIUPT�A����ܖ$�6�_K���9�F����vWN-1&���*���q�d<n#�>� ��pX���j�0�����=�\O�)k�!�!BEg�u`�w�����(f��J�r���=x�cț��q�x��ݪ���#�.K©�Ԭ��Ca���w��vbaCNO/N�܂���O.W�Z3���%�\9+�I_JG��B��O>9J�����N]:d���W7���RP�e��ݰp9D�nQ�=�'�ۤ���~J.9�v�c2��!V�yN�ŗ{�5=Be�w�A�앮�h�d���a�^
Λ��GGax�ѣG{g[����ؖ=Shd^9JoT:U�\���Z:]�e/k/6�#Y�wi��s��9�J����]�����@�e{G�R�/ҭXN�Q}ׂj���v��'���~���/~Q3���ZxOٞ�<�gs%^�mӡ�W?�M%���8�%���G�9dk%�<y츾a���a>u��U.X���{�KX< v~�On�kPc��e��K��TӜ�;Gx;�˚�"'��$�=O���d;3�m�J^z�.�_�Z�E�Y�����.�ܔG���S�]#/% �an*�L�x _��{Թm�.�4�D.eH�H9sͧ`ܪKn��P	ṭ�vol��{\������1��2�GS��[����14�k��)Nj��z]��ַt�C��x^���_�rPM�CS�N ��hx	���\GV��G��
�Pvf���j�L,ИŊ�G��}���O��P�8�8�3�N�e��4É��|'z��=��f��q3�V�躖���6���8���n�v
w�_�37ӱn{�Y�ޱ��u\�u��iD
�K�rƚ�:�̛�ɑ&���A,�A����uSi��ܡ�2s�1�߳�]P���K�t��t$�u�Bj���w8fU��N]�8H�B���=Q;9�[�e6.��vj���w��P���eu�k~��a��nP6�ZV*Wyw_���>?+�(y����r�	f��y����%�K��Vj�C醅CO�`�����/ڙ�(�֮=�*=��j����G��՘{��h�
z�;b]��#bRCf]A�<��է���)�}R�{s�iT3F��'�$Tpi�n
z�J'޷��$>�}�/�d]!��o�3�eś�\O֙��ɞ�O��vXԷ���9��!���/7̺Ck*�lk�X�7x+�թ�61���wDL7�bVV��Ҭ�ot��m�wW�k'qP��3�Y����&�R-�િ[�,��+24mJVAE	���-=��h�//]��f�W�-æ�Z����bIuM�͜�h��)Ƶ=y�"�9o`
�k���9գgT�	�o��g>3�x�tqh0�mm�3c6��Ԡ<������&�Ы���Z�5�%6�������S���T���u�e�ƪYlz�#��'�n���ݹӠ)�����g�
����S�=$���V�9x�z�՞��q&B>�VJ�~���.������ig���V~[�=�4;�&��1O}F�Q��7�2[�&��1w��:���8r]7���{��^B|��P�B�p�L����/���(K�0���{��}��nF��w��ػgty�.�k�f=~���P!Ř��k�z���S�8r����u*���7و�8��]��s����u!��1%��搭'�!���=��Iʽ7j�ܮ��k��l�ӳrqN+�!��V;��h��S=PL�uE�P�B�=��^n�=��4�st��8�J��"T���3��n^����\�D9�t�&�'\^}B��]��Z,oX����I�6����\{��\?zs�}p�6�TA��*�K�M����%k�'�o$O��잽��z�k(T �>���7|t�-��*��l�Η���l�1�<��Y�T�&R���'k��]��ܑ��`7K�A�	���H5�&Z:Ă�J�2���S�K<��(ȯo�����+�4z�y[�)<�K��B��[;��C,.\α��+=~�9 �ߨ�Z��}������b�5�x<�w%���]�!��S33n��~Jx2zH.��R/�n�9_��6JZ��_8�D��������l��yeȓ��oeA��b6Q+ah��5*���J�K�ߍ 6vz�<�e5��_�h�Z�.M�W*<��2�^��s��gר
�ϩ�u��,u��}^����\K�O9Ft����KhX<��q[^K@�G���̣�x�)���i�/�"%^ZE�z�NNv�MI��zY��_#�O���0�~w	"�s-�^�o,�l�ו�a{U;���Dir���|㉗Y]��g�K��n�?�qT�w׶���k�) ����ʥ�nc�V�;-�RK�k�`�*�Z�&��o�.�� ���JzP��[?g|���^3����+:�<rB�����H�#��6Y����襁�ʨu+�6y��w�Ի�0������t���Ϸ]�w�^SƠ/�:�2d?nS�x��Z�^4֊KG����x �����h�m����A��v�y��wu��wG���������f����J�]�h�m�"�W����;��z����u�zc��b��g�t^1�̵ʘP���j��f��ٿ!թh��0m�pj�m�"H:����Y�]J��UY��j"��KY�L7]�!j��M�T�"ץ(=��=M���S���i�k����<�b�/)W���b��=toT��
�z�.F�!x��5�=9�~��έ�:j��U�	1.�v��:]�
%t��;�S>��q�WS��)����v1�q��<����I�;�G�	ٔ��{&����o�r���W�=�,X��ԡ�]S�>u.{*���;��d��l��T1�J؆Yذ�i�tww����d���D����W�q��:�W'P������e��Kzu�u�d^ir�s�d�{!Î�.y$k+L��`�v��l;\��㥝�O�a��'.��<��j������<�6|��ӟ7F֌X��_�Ò�t����yeJ�)&bj���'1��奧k�O�c�N�/�2타9D�a�>Neؚ�ݓ������Z�gI��i��]�w��#M4�ڿ{�cy�)�'C�����2��@�tC�V�fz a��C��Pz�+\������g��J�뀣`yǈ�i�-�d�����u3k��K���ڻ�J�DF��TՔa�CzļaL��i�%.���F���R��fr�y}�y�q�(E*\�=םoT�elq���o��a���'Z��zݟ��=�W�H�L��u�)�pξ�N�A8άϦ��X�SF��g8�l��_��Ò��/�|.�S���7\'�g�!
S��Y��8���^���W�X��r���A������~��zD����J��P�m@|t�P֣w��%?^���V�p�=���s�3����q��SV��5)��mh�ZU�1�4�H���^��<�,L�d�f��e:gs��x�˚�.�y%��{�s�6������q�WI���3�Ԗ=��\ی�P�&��/��{��9�͖����E��uaW�W�^�N�)=��+,f��+Ȫ��]C������h�=�G������E0�wG��r�rΜ[kWMy��޲�ˁ���#���]��:fo����0/�����#�+8�=��Bm��{(��ج�Rh�)�6�]���~+�w!�C����j"�l�<�T��Gi� �e�xu�,
��s|��{T�&��C�g�"������}4�C7��51Gs�Q��n����������*b������9H��T�.��]�+r�=t�ַVW�̽�.�(��9�csm;����p�y���*���O>�ۦ
�4��PuL��CmhN�n��]�ײ�-])X�����7�m���)]���rY-�:):�nf��S��-��o�0M0����r�&W��_o,P+A��`�Aso��W}�^��/��]�a~2��P�ZL�E�X,Lk�Id@�w� 3M�W�����;9�+���s՚���_{�ј�=����p'�X=][���:�2����+�D؅�k~�FS�k�=;��tK?-ͺ&�Y	X�䊎i�a�OR>�~���nU���wy���o��&$a�J�6�G�'�GZ;�>
�
m�i��VP{��(��ű�{��j���\����o@6���,���W<��~��qP8���mPu~_4�6��t����ñ��^����>u�,��V�?<�Q^ڲ���x��̗'�y�����=�G�3�s��m��Ю�]"���EI1�߆J�X"�-8;�g>�\E��R�
D˺�YIe��On�=8=�/���-�=�4;��p�J1O}F�b>ͣ*�7�L:K���/#G�e��3i��]�P
]hZt9]B�\=��YZY����rǎ}5���:�({uD<�[���yȣ��d�t꺌�J�8R��_��,ļ1sM=�Y�(vdč��F���X����X�j��4:���L{p�ѥ��U�_uc�R�)Fϫ��=�Y��p���6�s�Dԇ��a���b�n/#���~��������룧>�̓��3��N�.c�kD�������R>�������7IbU��#c�gs�fzߑ��׳�p���	��t���Ė�F���C��i��2�jX�DOns��q�|wu�Pp�=�:�R�?�e�y#���E�PL���w���yt�`���l��˚�B%vN!��ܴ�j��H�ss(���o���r����Y(MEK��v�������t�}�^�`u�U������UD��M��/2��F�!u]4Y^����|�p�Qq>j8^�ٷ�������&oQǗ�b�����S3y���N���x�#؉�\U�SW]P|�{M;������5M➦����o���hl'��v��ن���U2���I�wU�!���xg��3�]\�]*�"~oƀ�4^���f"�Xϻ�����`9΋Z09d�Z��]yOu0���k��I��t������z׹%��V��O�0��`�~�IB����~D��!�.�v|U�]+���f�-��F꘴�ڸ������	W���H�2ޕ�tׂ�z����k6��R�mn�;V�h-l
�]��|��hnj�@�4�dN]���K�����\[�����{��qEո"H��<eD��uo7�<p�ub�u���h�QZ���e�b"�S5��p������+��=�ǲ�=�|���_sɛ��W�c�G�s8�<��s�X��b���`ۥ��	����U�ū)�}g���G�{�|�ʶaoh�t]�����%,�𜂷��wX8Vj�OJ�k83�j��=��=u�KT�7�:�ҔW��T��;ܯ��mD�Է삅}}A�c5��k�B}��ޥڶ�+���3���������E��X|e$�zU?Y5��BO����m�=�������5��`�� r��	ƙּdZf}r�ㄲZ%���Y�R{�ه3�K�2����]V�5�X�}6�L��g҄�Bq]�U���\�x�P�V�m��op�VW�������21�"��������R��ty8��~.�3s�=|��u'�����9�u&v���R�ײ����pL�<�O*rkrq��9\�N�u��ywGc�a����JD�3�`!A�c8�vu��w��������nF��9����b��OOi�nl|�)p�	&��+�du+3�Ca������7F�wB�S�j�0��;�����N����D!��GW^݀fڶ�� #� .�%�w7z�1���v���6��n�.�l�����_��!�(�U�$��]a�nڭ�$�[�:h�}yEy�+���\�*6p#����wh9Ί�g��zrS
k���T�c�F�;ƠT�<bD��-�\7j��Jh�կ�1�ٳ�Q��SN��ݖ���B��.�."F�Q�=�#>�Jb����z���k��s�.�u�j͛������y�*��6�6:Q>s*�J��~۩C��F�w)sp=�y�� ��g7~p��mk>����uC�^��Q�8�3ԭ�U���R���w������Z�4/�y
]��{�Ҋ��mPg|��/�=�>8�Uf�U]�����ڳ�[�#ηr焱my3f��kgRܕmTG���`\�9�o&��+�Q�顊��I��v�`dwrяo�yMZt�JnW���N��mM��h׎����4�w�|�I��q��s���sW�'��9��� ��;2��|�{�*{&������ٱ�S��iu"Y�ۄ5:��u&���O]xD!��~�5�գj� ��m-Κ�h\��Y�>��T�.�<q����3gZ1��4ß';��)����[oR�-}�5����bnb��x �>RQ��������Vh����pC::J����&��.����5%�����)�ɛ���Ew&ÙԲc�-��
R^E�A�����3L���>a��d�Joj 7YYi �����>�:��dx�w$��{
���	f�t�
�'���=ԣ��Y�nnqUr�e�T��
�E1aF7z۵rY����p�!�S9��⼝{nC��]��� ��1h�݊L�M�wF����V��)z��7nH|�]I%R�W��J;�=4ݥ���t@����Ƕ�f˵�^r��c�o�� V�V�qe�.n�=.�̅�*Qղ����u��S��s��%����C��(Ӌ�z���Wj�m9�0:6�˾��:=�Au`�fL{ի��Kgo]�~4�|z2Q��]����\Y.�Ԫ�we��A�3�q�9,%U���(�*� į�1�hj���t"�U�r��K ��@XPX�{t��v��ʼoX÷Qt�m�Ls��2�)R`9Px;eL�U���8'h&b�� D�0�
�д�t���P[:����SUsX��ب�;� 5�)t�e��/EG�o3-���:[��X�'��IS�*�c���B��H�yf̈́��I���]�X~�!���ڱ��dV/엤/,zD9��ʶ+|0u2u��i�L�1�j��G �F���"[WZE�VŊ0�L�c��pٮ�{�]�>��>���4����ж�3xmA�I�Ss��Hg3�iMv���$��O��
"��1�����y��&|C��:"�<��H�T��3^���cYZ��YcCL]�1Cԣ#m�� y�o�USy������K�,@�H��m>����r��e��.��8�� ���$�����7W�d��*.^��'��Y����e$�Z5ػc��]z�/�e�k3Vɡ��a5t����+��˜�S1靜^�N��e��Z�7���L˘�# ���9��d��`�%m�]�U�Q䏬A�Z��'JU�i.��x
瘷(�ǻ�;���m�Sd��[��e�t�#�y�R[�^���d���K�`U�ɑD�}Lu�7zt���n�&h��-�I��P�c�V$"�u��t�Rs���"89S.��4K�/;,a5���Ǉ��pF����Z$����TJj+O���(�Xi��[a\ؗve�h��c����5�ӢM�wLD����%�X�W��v�I�.��-����m"���:Rm�rI,e[v�3Y*-f�BPM���l�{�ׂ�qچ�Ǥͦ�|���w{6SםО��+��ie;јol^H��w�v���LK������4v.8�ۜ�Or�������iYqV�'^�ndd�x�j�KrV��eN�M�2(�B���ǽ{�B�O3�*�zVe<�V��.�8�y�����k���~��}�0EUD�TQTELU3�TU$�DQATDUUUdeEUE%ADEUL�QE��KT԰DQ�MEMUEDT�A`EMUQM5DQ���U4ETCMUEDUT�QMP2TQMPD�UQQT�NNQ3V`U4T�ACde4EMQUQTCQAAIDA0���Q%TDPD�-�3ddM2U1,PPMU��MUd�DDFf�MMU-H�D�Q5EA�٘NC��U@�ԘQAjr��"��������h�������VM�f����i���f��59Z����2�(�)��������sf�`�(�bJ��jid����������̍a�D��1L����*���2(�I�L�KQUPTU%��)"�(����&���f�j�("�����(*bjJe��(	�������)"j�Y��QS2S1E1SSSS]����~�F�v�jý��2Z�ݑHrX��S��|�a�8��gs����9�7*ٝ����Vҵ���t��@��}���k�ӻ�ѥ_��lV]	�A�w.�'\��:fo��F��ˬǆ������L���{�u�\�w.\�U��M3��qw��Aة}僪�b��<�T|t�|�Q�� �xt
�-s�g��ET&���9���2��zOV��(c�'������>���z��Sw�+������}-�L�W�"�}2�)X(7=tR-+�T�.��F���3>�w��>|o=2��n0�f�:ʅ�.�� ����eB,J�bxB�����N�uQ��ҷ��*i>�͎��l.��C�"=����9>$��=�PóƵ-�p���q5��N�0�y��[I���.ن��mß{kH��a.�䊎-0|�5�T�4�gӢ~��VjR;'m�0�Ω`��qf���-kh�ੇ������*���w��B��-�v�ޣXYՃ������8g�����K帨v�.b+'�:_y f>�ӻ��^������B|Z��C���m�bVv=e�U,��ǖd�Ы.���7��&<�|6�q�����wx�5�%$�L �2��MV�Mh����V8/v�޲�Y$!d��-m�q��<��`�'��;���So�b���M��'���M�kW)���gH�;���!v	�f&+2ɅnwhV�K����\ׇ������k�������]"���EI�	��yw��l���%Qfi�x\c��>~e�^r�t.&CW]���f��q*�fp�3���QQ��4̖�+g�̋�	���m�3��W���CWP�-��u2�ZY����NX�y�����3���fܷ����8����m��e��(�\2%�L�C��b�b^�����ge{�V���ӑ�<���絔��.�qzq���'c,�O+��\�0�Z*��˪#���_^)�n�x,�=4zyM�sW�ZZ��쳀58�,�'yX웙\/���V:灬���R�4mA�"W8%��T7<�ehhC'���e�:�-���dМ�,Sf�sN�=��w����������i�2�'�#Ǔ���0:�����P����3ꆽR��l��u��suy�{�m��#�[
g�*!��01'��'ݚ����xu�<��:^�R�=�}�sĭ���Y���y��:�u�]�\O#����V{�xWx�� �<f�\�@����VQΚEFim���qY��w �%K&�97l�ҝ��6�TM��c��Q+M�� V쬃���r�M�1r`�&Y�;�T����ۧ�Gws��h�Ӈ�^�=��ݹk"1�`7�m�����ފ�"��3à���C�/3-yR:Y�v]Qgx{7)������#sm��BI�������ȫ�0q�-hϜ�t�Yj�u�<:�h�ؽI��G�ĺ{ϳ�+s������mq��-%�
D�7������ˁ����!�S.���Z&Gܒ;��&�xB��sǩ=��X�{�	^u	#C�oJ��[˧��=WZ���b�y���W���mʳ�oL�qX#ԤY�,V���>>q�-D+wӮN��y�l�3z,�l���q��\��~Yi�9o�N�>��:�t��
u��pg��ΤY}W:�-�wW?i�`�󮗷ڭ���e��6�x�UC�X�(U��梽'݇�X��+t�;�����v�����^u����G���Ĭ>$���[���}녤7<��]ܳm؈�����{�ƙּ�Lυ�
+K��ɛ}��>v���������eܹv^UsHߝ�=�]��Y(Nt2�/#��C+��f�z�d$��ǃ���գ�5�5�Nf�5�-���U%$��8ZJ�Z��ѕ��xu��	�[�w�F��L@�tP9�ñ�%X.)P�e�m^nV�|��WR�a�Ec�4��Y ����|�˯%ɞ�0��R	�{�+F���<��:g^�.u�q���msJU��Ӵ�T��bd^����{�h�y9�O�Pv��h�T�v����l~ݢ����G���2�w�֙�]S�K�^�W��s�Q�LS�}�h:�(^������K�wp��|���H�_��8���u��;�հ,��9c�^��n˶�˕�\���Rײe�f	~}�G�\������nuX��x5�*~qf�n�S��%�0��z_��ƜQ���WK�bʤ�$w�H��=�f�66�ud����f횊�2�V��9�֒�y�^v���G����a�f	�ۤ��������؋Zg!���ժQΡV���cޖ�����Ѝa�]ws�����x�p�\�'��b�i5f��Kl�1�b��}f���^U�뀣��1]��˫h�y�=�s;۽*ҽJ}��س�:j����h�h��g�|t
vi{G�R�׎�y�Pl��kݩj��®�v�<Y)��0h�g���Ú��.K�yx:���)[��;�^<���:<ݑ�.p⬆`��[K��0�x��q��[D��'�zg�ڙ����_/C`7k��Y����oRL�"&�� �)Y����B�;�-7�����
J��vw@��w��`"��Y��q��&�0�tT�&=~w����3�-����9�v����e����;�b�ӊ���v��1�������WOL����Ğ�\^}\��˚�.�y%��{�s�p�/�5�L'�X����Ww�ۯ,��yL���H��sn:��x��hzq����t#�wʡޯQzG�1�ڶGV`����͍�fp�l}��V<���d���[9�L�j<���3��7��'�h�f`�]T�K�]	���й��
\���k<�L'�>܌����M�5���f2�� ��=�w��֨�r�G>�)�C���>�Ƌ�픡�XW�'k����w��yأ9��	t��b��fu��Ri]T<�PL����#�'f�c��M�Y8r�u\^�k��t^�離be�kD��]�G��h����{"�ǵZn��2Ǩ���%��w��˸{�C-h'�r]O
ʆ��:>"�+��z�����rR./�w_ެ�� uW��v��Xa�.��p8)�6��Q�=���H��"�._�6!�h�u�x�I��p���|㕻L�X�]W}*��fC�!�rv��Ơ��lJ�l�娊�β��Pټh�[�\�U��p˧�]8��f���m!�WN��ƴ�-����U�F|���+��b��T��y�����b�J�d:���H��uL��nj���V=�"�۪���>X|q�9��==��'
��:'�0��rF��Cm:G��+g���<r��Wx����G����ǒ�7�����ή�O���ݔD�0�ud=���*ӝ{��u����t��yuRn����+�s���7���I�^�� ��[���C�_=�4Ъ(|��M���x(͔�gv�YOvY����ٵ|�z�ȍma�*���q�3�I1��	��w8���W�}5��>R#j�&E�dyW�n+Ϋ,��N%[L��a�����wW�Ur'�ՅL���Rs�-w�cT���`z+h{*!
�p�S--,�ws�#��t��A�t�ZZ��O���~�t�1�%������9�f��[j`�qLP�	��\�H^+�>�o�1M�>�5��ˢ���8�����pT�qu.Dz-�UW������������gR�T3{�6%�]r��ퟯ��Ő�yX��ne5�'H��E}]���'k�h������t:�*��d�f�N���B��
�)�0V5C���`*m�.D�8:��qS]�i�t����3�'�� �HTq���+邖]�Rt��q���U��r���rf��fFm�I�,WaۍZ�V7�"�����ڏv^E�oAv�8��L��zgE���T\k&f�b^�w����Iʶ�e��"T��z�I�Ix��2�2�e4���#���>��wޜ�_Z��=eD��)��b9�{u���~o�!�=��5�]'��L����63�j��/��|���jXW�Ի<h5�����.���޶jm�8A� R�#���:��.���ß7���Q�3�9���;�]j��=H���8*Ό�;r�0��j�l�;��~����v�Gwr�ZW�d�z׋��:N�}Ӱ$������|��c��3�>�V՟^�*C��}�ՈV3�$Di�a���i�-f���b��p69�rԙ>X��XQ}�����!Y�����Py�+�1d)�ڶ� ���ޘJ��p�-̷�{����1�c>u�8�Fr�'��ܡ,���cA���}�/Q���i�=j�x�ͭ��J���j�6��֫���X�YxNA]�E;��5t��
u��E��ȇ�+8�*�r�L�ڳj�E>�t�!�d��~����i]Zu��H(�aͼWj��u����i�47����p�ku��r�3�8�t&�+|�}�Cd{�[a�+-��������i���M���;f�,���������ۑ;��:~�1C5n�j�W}RҺ_PPgb���_�W�R�S�T:����_P`�M�+��.�n������/)���n�d>��^2(u�d�~ܧ������%�MmUq�Fc���7޽���=��613Ь{J+2u	��z���L�BE��
�h�W�0?�{�����\Sg
U�g�.��UF��?,{H��xV}2�<�:�G���i^��S�׺}�o͑�%`��=O �\^];L�J�2��
���ΧdЇ?oK��F��$��&�=��㕈Hs-z��28$�L�C����W)�C�p늴��T�j�KF��>�W-���r��������I����d�:D�!��B��<���<�"��\��R���5�u-Is��쩃�m��e�!���FY�P*�^I�r^�du+!�}����_d-V�G�xM����ཾ�ى�5�WcN}%Z09br����^�J�R=�G����K�/
V�Qh��Y�����er�Ãu�J�=,J�������rW�:KO����Y����̗��fY��̮��?��]F>�{��cг��;u�ç�r���t����\E��A[Z*B��ڷ�M+�n@;:%�e]�=M��Wd���WK�Ėv���WA�5�EF�y�3��h�8sB/������Q[��5B�qܚ��9\#���-C3�eZ2�z�ՏzZ*��xJ��F��2N:��Ý����+\�R�Ėɩ]�؁�����an%�����͡�`�����+z�(��MH�go<���9߲�{�ꝷu�e��3�f���O4���O��]o���{ĥ�� ��l�Jsh�M/F#����	�\�Sg�Vӯ��A�ysP�RU%�	u<�;W�r�I�3&�|�^�e[�t��bڞ��`���ZV2;��n=�=�5i�CR�=j���I��x��&�56�Ѻ<�F��h�ޭ0�b�\^
�x��5xD��/�������ӣ�mMQ���idv)K�L�|U�0o���ɷ��v���i��o�{$˾���M��4�W�+�@���ԝ�J��p61�J�������%�0��ðГ:�^����l���#55�~�-�VQ��\�\C���ܻ���Wj�y8EF��T�-��CJ�	5���7��3�;�G� ��`9I��C�ѭ��5�XY��vBr��:�I�{[��bf�S7��2M�"N����멷6ǑJ�7���"ZO��G;�^�m�	�
T�u���0�󖸳�LO 3β;+m��:�*>����(���W����i��3�;�#d��n�ޭq��-�:ջc6u^�7Y2E3[乡z��w��!��Ks9f��.�U	�>?9��N#(�r�J��&�{�&�d��N�P��~����Y�3���ے�쟂�yg���C��L�末��Di0�@�r��v4E��ih����֓a����Օ`˸{�kAɕ���Ͳ}ެ��:�:>�b=��B�5�\\g������,��|�������SB�����w������F�;c��qב��1��w��o���^W����Q/V�-����9j��K�#u¦�1�D�Xlß|�!9��Hnz��=���;�Q�X��9�)��-���ZF��>�Aa7.�agV}�	ӳ)E��e����xk��s]rc��z��oEb�t|�sG�Y��m���P�\�"u�Y+���柲�>ٹuj��� V��kr<x&ۛT�{���GX��'���rz�
ᮀ]#I��ԣ�^��}yEn��z�s�H�K|�(�ۍcѷ<�A21P��^mY�}�D�i���a]�"!��_�:סj��rV���=B�f�����:�ϙB��pG+nȌ�����b�e����Q��`�0l�#�u�Ǔ�,��t ��9:���f�*�2S�k]��O(h��v�-u���5����kr�2�AՄkd�gfe�v�}u{R ��V��V�]0+���y]���s[�Tb�G}y����T��Z�5S��ޗ,��U��h����{+�o[y�3��n2ض�͇#�
63H���A:`�@��{n%��Z7!Ֆ��f�'�1��8�\��״�_g*Al]�d�A*�da6j��x6Z�n�篍<�e*+���f�P���j.��=��EF�|@B7��k�Ŗ$:n��&�����s��gVB~�U�*$��&��>#�-N���`�g.�es��h�/C�Z�-;�֡۳��P�x��B3��0Jޘ�x��+�\j3��;N�2�Mu�^\Y�rPW��c�)��Ԩo�}t$ס��:`���Uu9K��h`��ʺ�E��N���f���G��崠Ƀ0ݦ�kU���ڥU�\ܭ�T���N��;iv�s��K��^��5\��}3�*����&t�;uGX*��j��
�\�A�q<��(�Pg�]C�I[��݆5:���EQǅ�6Fq�Z���f��3-��7�[���Lӌ��{��і4�X9�!��qKl><-��k2;���.��kэ-:v���#�HO.٬���J]*!�a�m�g9���p�x�rU���=�s�J<8��哶ka�Jmv^�rW8ݕ�#a�A�L��S�3�P�]����MHb9��捸m�^���ӴÜF"��+�ʄ����J�Mⴻ�s�o ��#P�����.t�IIe���O��s���Cm�I:E�qꙴ��ڏ���Zr��L�x�&��iu����7h���}ò�M��Y�.�_kM2������v�d#��ŵ�ľQ֎�t��U�K޹�U�3@k�T�ޚL�����ugzΈd�-��U�sʖ:�e�hU� ��m��=�W\u*q:GZ�چ��L_%w�h�n��w�NVBL�g&��$��17��Z�j��)Y�Ck3Ky�񾻬�yu�L7��r�!�U�|�盻oiVa �o.��Kg ޶�s�����4Gu�'��:��8'�R�P~xU=D����D�/b��7�%(Զ�]�qj[�2�,6��p�m��\��d/�/c�N=ٓ?H��8������UZ�of�y�3�Nf^�16N�,�S6����J�mx�ۘpN�Sf�t�kObc'��m��ht��}xl�q�#�myJ�s��7#ȴʞASv�ٛ��cb��v�ŅR��YJ���P��@I[���7���c9bDD-ҳ��J>x�8v�[hm`�N�����y�fʻt��#�z�.�;i��J�=jptu�&�tU��P���uwCPQRA14SU5$E$QTUP�5CT��UUTQQ%D�1SMDUT$DQ�PD�ILT�ِ@DDPHACU44PP�Ea�ET�LAA4��DIIE1��&0�̕1T��Q5�DDTD5QIT�5TEVFD��CD�`UU9��UA-QSTc�UT��d�YeT͐`Q�dM3DT�%A��ՙ�I�R�Xa�e�VU�EP�M�َEMfd�UTMaAUMSDfffL15���S���dE553��EESUUAE�4ٕ�T�MMM9��ADL�Y�S0ec�DQf8՘�fa�cQ4M$S�DY�4FcM����VXA2fbPDEfc%e�e�Y�Xf1DQ��w��{���~@��u7��u�F��w��F��aRu��0���_Ʋ�i����>��`���u��{�cIǽ]�+�6��%w�������&�i��W��Km�8�W�0sW�ifgv�z<ghI���|}��mt�o�v0�m���%�������u-�6�"��(Qf$�n�ڗ�L=~p����5�}��a��	�fi__��e��T�O%�R��ʪ�7�ŰC ��t\��՛�+1��]m��^\���,�54�??Z��̦�'H�ګ2L�+{:����;c�<��\�a��2�+P�.{Z2��H��g��A���������W���(�%��q�(S2�S2�7�S��������Ѩd=fU�U֍f�x�f89ow��=Z��`�0t��G|,[���|2���|���O��Q#�ء1ˆ.Y�^��c|Y�z~��u��tGAu�61%[���ps��*[~'3�%��*dF�"�˹��AVtd���9+Ì(��p���<3�Fk��K�1h�n�5��.�{���I}BJ��(���'��u�3�E�������2.�3�p�V1=w�^L��NV���%��.���+��n�=C_S��ײb��>gɡ컰z��.���E�k:�V�f�JV�M�7ц���BH�ɬ�f�����q��/�t�@�G�u`��dLF��F���3�������5m4vs�ll^.�7<s��3���Z࠷�,0\LY9�C��ȇ�F�ӕ�P��i�7A�=� 8*���"�Z�:/q?0X�o�/���k�f߈���0̻��|d~�+ܭVp0����	Mh#)F������f��MA�qZq=~}��r�l*����������:��cU�E�`�dLv�m�uVw���.aΖ֟.���i����u��Z���ʬ��Q(|��(cz,y�I�Q��u\���|)��xpd�}��������ϖܱ7Qf�V�K2��S/��t��b!f�=O�  ��+��6d� .\��ƙּ�M�N�p-Q�]���J��t�{�xG����J����it�=�]��	΄ҟ��bv�Y[����e�ǽ�\�LV�D��9ggȬ>k��)ypuW�¤�ds�vMxԡ����ٻ��.�xȄjvU�ٔ̎�x���쭥�E17R�mۢh������N�C(�n��T�b�������e0Hv���
��A+��y�=]��!�>�o,J0���~HYIhMZ,��(j��\,�!ܩ����Ô:�v���/K��X^d���U�L�,��6��� w2�i`was�}��~e��^��?3^*!�K�u,T����@p�k�Z��K���Xr��\��zV����^٧2��ԙ
ܙp��/��Ϣ�B�R��GR9=#�9h'��D�{�B���ώKW�k�Y,7�ӂJ���',�K�b9�`x���.��22���ܵ�w��EX�Ӧ��{*-�87h�`�P�]�e̻�V)�VW�n�2倄�-ǫ��[�E�Iq��Qqԙ����2׼�����F�XI��&���7Z�ӗ�}U]�K�Q��/�,�G@g���ު��-�7Jj��Oti0��kV봙l��X�Ut�4o���ۺ�2�h��9*V�12xm��Nx�ī�5�V��M�{[�}���k��X����hO����=jݿb�.L��i�9��)u3��L��y�9�w�G�q����H���Xf�}3���GP���ס���Y>�?`N��s�FE��gd�؆C�.r�z��KX< j֎�]�nT�b �z��_�ȕ�4X�d��27:�87n����N���.�@5�=��`��`���Ĳ�4z�h���(�ve�t;P�������I��VX)µ��s�̓�z�ޜ��QΩ���WK-����\��Ʉ�ZN�VT�ܔ�$lk�s���:�9ؖh:��st9R��y�ݻ��)��$4�mx�L��H�}�R%�N�E���x��r�%�5sV=|ޠ�l`�o%OT�ڙ���6E�ԨzU0t�(���_��z/Ŗ�ϣ��g�<�<5����>�i��A�^(�x��%�7�"�%���&V\j�WL�yZ�=��S�}��鈳by����p�w��e8b�)4l�!ž�QK���eך��Ǹ�q��ȯñ�j�3�MC�B�s�93��`�X�g�ĚƤ��0(&���^��O)�z�����mXx�W�݆�ݕ\�+���!�5�L5�>y5R/<}��r?I[�;��0?R1+�ʨz�.֥�ᩙ�^�c����P�Z��7�� �ji;�����cT�(o�u:�/.��-,�؁��:Fk�0�SڏB�TC^���}�=��	8T�q3��ȇ>u�lh;i���a�E��y��|S�6 �5mw������٭Q�]��)��҉جчΨ�^�jh��j�CǶ��2{	]g.�y��n�e)�Oӥ$������s��y�u�Ha���­rKk���&�{��+f���F������5=V�Y���J\m�:T�bh]5ua�y,g�[W}��AV���ٹ�}�����#�ϖ��`�}�[�<����m�cvX'�����,,���	�cg�3�0��M�nb �\���E�~��X�-�"��P�k�Ӯ��k�%*��sO���rЙ���͟^�H���sB���x@�GMˆ�ͫk���{~3�Q�3��^���W��2�+9�j�Rt�K�
�O��g�C�]w}�sj��{jEZ��˳��u��fA:Sс=�̀��H�G�'�WI����`��[h_��4�!^����1l5YE�pn�Rُ��-�O��N�΅�q���%�������#4��VڙJ�t�S5~��~
��ֆ�/.wpp,1��(s��4���_,T�qu.V�=a��[C0fn̎G�O7ۻ�rZB��%�᰿����������*�^u�*i�.�՚��^#���{���祣�8Ԥ˱�켪�XN����?K���	��/Q��mY��pi���Pu��|�;���*���z��3~�f_�\F�v��~w|f)μ(Q�MK�g�
�m�����	�S��f�������]���
�������eҵim�1`��z��m�ׇ�ex�������}ya���J�:z_u�	�j��I{�b��|�����M·^X�*q-�����+�/��D�G4�_vnV�s�v��O���r	똳�<�&�@���ԑ�-��+��ޖ(�m����~��=�I�3��L�|]n-,�^\���_��p<����G ��o`zqu\�[���	j^$罣�����-Pc��ϣ��? e�� T|"�	y��R>����;.���ВR���<.j���m;W.��ׁ%a��Xr��-xpr��҅��3"튓�[�]��]���Ď0��O�.�f珎5}�-%�
d����3�tG�3�g���'=�|:gw�=��V��J�@`?))W��t_m\CN�za+Ρ$qU%��6z�����W�����t�/k=]�q�8^�b����2�k>ڳ����u�����Nh����+o�Ok�R^�3o�WMk�[7��4���k ��"��ۻ�]GF= �S'/o=��{ӆr�-�=�W\����g#�Fw���ux9�D�����O���UZ�.a51��W��Pc�n����>p��'�)t|��=-�K��U���%��U��&e���3�/��ђT�Kc3-_���]yy{�}�ť姒��S7�{9 �Ǝ�����0��� �J��9r:�K(:{��;å��c��a[ۖ��܆=�4h����ο��R���)��P�Ǽ�Y�9L��-R���D��� +`���Vu췅7y[��l$h��d��2M�\[)�I�.\��%�[����N�%%�&8C�Wd�6<	��K7SE�u=��g޾��,?'���xg�	΅�U�h�~1��\�����^ǵ�ʃj�f$N�N��VG���^\�p�;2��L�ItH�FD�.|�ͼ�x��v�»���_��]
�u�wj����Dh�YξDQl���n��#�ŵ��w)9{_O��pL�<����0:���+'�D�����
�eK��)�LX'{c:J�&|-��>lJ�:p(f��IS�ˆ�/��ȼ����)�N��yڳ���;LCŅ7�Y��^�yYlUh�6S����i�%Yџ9br�~	cZ�/f̮�ŭ�̚�Y<VjV�B�����������ݣ��B��.��������Z.XV����37�<���iƉ��z�^Z2|�
L�xA�	1���k�؅]��u��D�1�����Dz��y���hH���^���4�T�}����b�Q�E��7��Q��i�Y����cBgۗH\�����r��Nge��2�9V�����:��}_vQ�3���LdU��D�"U�[�\�b���,<�]�Z�SVtÄ�k���˸�����Q����᳷|ܧkqJ
ܻا:u���6Tݽ�o��X:Y"����ٞa�5��\^_f�
�˙'}��o�gJ����gF�Ѥ:,����*w�|M�.�|,`y個鍇�j�X�^[�v�\�\��'D�3�̖(����W�3o�`���ZV2;��hǷ�~���y<e���&�ϻJ��g��p�b倿�:_=^�� ��P�]�9�t�zq�{Y���R������=Or`� �B��ϗ��-����:�,�`:��[[�ᦰٕ3�nc�yw�BGS]x�=��)��q��d"�Ll9�%�:��T�����\�zp����s�A�19�Ͼ�i����^(�aq���$3�Wf#�K�G��52o��L�T���7�A�=��Zu���G��T5�ȃ�h����"�����u�7�	J���yf�NOV����e�}w�9��c��ٜFU�*���x���ϼ<�*��K��B�Վ�F��;��۲�����|�1��,hy�5x��4�>��3"@��qN�{��� ���{�@�K�J���b:`wV�
�®� e��Ƭ��:YJ_��\���<���G~;� �G\N�h˹���>���ܬP�i�Ζ�EF}PC�oЦ{�}�9�6\v���{;�Z۱�b2\R=.�}b�	�jx��w��@t�a�����*��w����X��Oqy�v^Šɔȵb��T���\�gG�S~�����hY_e�#ڔQ�}�긌\(�����ݓ��]�;�!�bG���wdB�#C��K�K˶a�����Ȗi��=:��K����4��2������v����8�!2eśX)���)���,О�1SC�z�u��)�m��߹�
ۙȰ��:a:ve#�13r�d>X���m���V2�s�C�vL�V���S}~a`�\��i7��x崜Y��x�ʶ�7���Z�|�t\��e��a�LW����W�'��
ᮀ]#�b;�n��x���LՑp�%n�g/J�7L�zpO����.���<*�~�0��"��cq��ɉJ%j��[���.�lT�0Gq�o�(v��;=��W�-�@����&���������Utn���c����8㷩��.޹��,�3�*���)P�'w��Vj0�Z�Y�^�z�y==צ�}φ����7:A6͸]�U�w�[�:��!����KMX=���K��I�pt2��_Z��E���z�_|�r�v��+������J��}2gl��:N6��QS�X��V�F��ehވ){����0@YԨZz��Y�.S=4�ٮ[,�S��ς�\����:���I�W���J�I;S�]��q����Q`�j/C�o�'��俷�26��:���s:��M�����(�`��沓3QzP�B�N�z���y��n�sć����$�hf����ܼc��.����4�ˌA3L�\FN��s�J�g�(uI^Y:�MkE�'�6g���Xg���@pZ�R�-��_�*%r�u5Il�l�;�������z:�=������ypyP�}�8A� R�|��ѱ��[�g�p*X=���}�oIvu��}9���D��s��gF}(C���>����J���52�^Xxg\��l���}���g�����0$���a˶|��c�N�e�_4Cݠ�n�rq��Z��h�"Eϭd�����E줓��bKS:����^�;�S3������[��D埩�aAv����I���b�}־��<~��poCw���ܩJtIx�7��b��-a.2�+ǭ��]f�[o	븧t���4�!X��29�}{���a !� ��X5pl�Z�	����܆�����b�=��K��Έud#���5
�͒å]lh�ݸ�c����Ŕ5���Ñ��3*C�d%#�-U��m�4��fv�b�%�ZA�0��|�=e>���b��m"m��'�@�n(�l���,P���l;OZW�)i�x�a�9�d��j*�]%+�^�[�����9��+��Y���ű��υ���GգuʻNC�KF�����x���-��:����y��⽵���\�>O]�Z��2��Y�a���Ҥ7[صl�6�Έ�w�����*Bb��i{B1\�u�jE{�i�3��W��׋`[�d'N���tsVA�kT�ډ;���^PW�FR���b���N8K[s%l}1[Uu�xw�s��(^P���WM=�:_WBo6�%�j*ŵu� �x�,���3iL6 =˪�]���)*"��; r��ז6��ҫ�3�k����g�_���W��)�����fq�b!;!�1S�,GEJV�V�Tʻ��P�l�#m����ʾtx�~1F�{���w��3�)��}G��.��:�;4�@V�L�_}ݷ6��/9wr9�?�veh��C�`k/C���l�������`�#��"�v�|�j��H�SY�&���(H�Y��n��,�-Vha�}���y�vr=|!�̷w�O54vsA-��4��qA�����~�\�X<h�����߸�&�1��dùRU�VnF���X38"�ɨ ���]��]]�MY��'*�C�����'R����b�#(X�}�J�9u���`���vs
�y}��^s����i3)|rX�3��}z;K���w�چYO>�Z̾�(�TN�E%w���W;:|��P��zr���h�ӫ��F��y�g���MC:���ru�Õ�8�{�,��
��)�ם�_G�tV�J��x蕵-rW(.����j�hm���Ĩ;s�΍��/70#	q�YL�{��{�=5�:z���:�b=xvً�~ԯ��;+��6[��]�uܳE+�򐮙Ǘ\o��+���u^�:�]c��|�É�w���v��Z�F�vo�Ļ:�(-�Mvڋ�k��l��c�q�6#��[��n�T� ���դ��ֵW���[uq\l���hp��1P�+��k,c a�_#(�2�έ����*�}��J�����ʳ��B;�*��듞�A�k�^��4�?w7z����:o#�jF6�MR�����h���$r�N��̒iVJ;��k��N���������lp�v�J�I�.�a��Mܨ�!Z,꫁ue�sozv�#}K]��R�sh:�`v0�7:�v�	�槶HuԸQ�6�w(o�����1+�7��9�ܭ�pkR?rG1EE��\��p.��h �
 |�'��$��M�Fe�EKf&Y���T�RRETVAfPe�QE&�Y%9eFK��TFa���TY��fd�E�3dPS��哑�YaQTYD4Q�ff&�Qd�ff.FC���A�c��fC�L�9�dM�E�F`�UQ��fe4fff9��eYSHaa�Q�FQe��aQcLe�Qfe�9%aQS��fbU�e��fc�FfY�YY�cYY�dME9Y�U�RYYfPee�fdVM�FE�Te�F��Y�FY��Q�NYQf95X�NYV����Ffdadfa�ReVaY�eY&e��6a�FVA�NfM�Y.fd՘faFTd��XeT�4Q�������Ώ�p��﫱����z<��_�Հ�}T�;f�J(J�+���e��7��2�tȬ	�4-��.��mK��>����ʜD��y�6.5��Ұ��&>V(�|*#�2���л�g|���ܚ���E�}B1J���>�����ƺk_��h���U�ƫa��T���s.4�M/&g�q��h���+�b�&_��=�w㺕9ì�r�g�yo�v�<6�Ա� ҃\�o�a:��b�x�qσϜ.�[:�[��"��p����﯍�� �\��8���ϳ:����c�,�b��OT<d�r��3�OK^��bV^�S��$�&%�PC@��ڲ�\fܰ��G��C�E㝀�����vb�Ǭt��u������z�<�dCi��[��i��ZeDΏJdb��W+�b�7Zv_�L=�f���W\'�ŵ������]>y�(mB8K� �����O_[�!Om�r:!E�m��[�Kj1���_C^*�s���o�t�4C;��TG���;]�6d���fs4=y�ڳ��:�>.!~PIS秲2�T:"�A_�=w���"�X�n�^5t�5(� Y��}1��ˊe���;Frä����*I}\�>���f()c��t���.���Z���mrF��up�; Υ3�ξzy��Aeq����U����67�}&�e��Pɟ������9����*���G��Eeo��_[ى�5S�V����{F��9b�u�h�@L,��jk�:>�Xg+h��#F-�\0!cn/PL�<l�P�2탕������tY�v���F��a��قx5�IC�0�����p
�E.�e��2	�z=�cmN#Z�԰�4���z}�]=v9�;�]2�	4k��QS�k²c���	j���]K��Y���O�p/vKv�U�iǃ������&�س}��դ�z+粼|��ɘw�w��hO��p#u������X�d'�.Y)�ԫkbҎ�?nY���e4��Lk�;�d��:���
��^:g6��ZC^��뙃���-+�$�{��{|oP~��&�S��:���<�~��f�q[ @�:>�B��G=Za&��W�Ս˚�ZO+\�y$|���"�ݲ��y�u�𵔲��N����h_T�y�bu�)m�N��^YҖ�>|s��y<��WT�	:����Cۖ��hb�C��Z(zU0lo�W�!ga�B݈�ş����>��V
#G"XL������b�.�{�ym�D�c+V��W��4*�g2�Z�h����=FH�ĕ��-����}a�-eK�W�,���>�:走,���=C��ew�N�J#X��յ!��Q��M]��Gn��}��דh�����{�a���mux9��	ƞ���XQd�ZK�v!�ZE'm<�-�4�b��eV�&�6�����;��ѹ(o,p�=�N�Q���3��S|+@~�6�P�q��|�Z�,��e��(.�ũw'��r��s�8&u������*e�'���<wjV���:���uP0t�0�[�ȡn�Lo+ϝ�km�U�[���2�ūz��3��Ǔ�y�;r�*Tzr�ܤZJ.-(w�@�kR���f�y߮���)a�vs�&#2 չ�z=�g�r]
�hP��g�B��w�*��\���fԬ"�77�݇nM��s�NѬ��,5M��OQ�0��.�p:���G!h�9�|<6=ٌ�߃�u������>� �5�
�.z���:৫�'���6ai+Br;�M{�[޺ �.Қ�s�osա_i<W�km��7���
�s 8"�ή�O����/A�(�c�fV>�C�#����u��@�e�����V���kzP��p4���\���Y�x��Tj���']�+�]in�f��US��E��H2�W+�@F�ck+F�]�p��+R���� �;�+��:�X�����J�6��������+�Vn=p7Ұ��}5�5S'�\9�OE.���].�^����S
���y����<��o}�}���L�8Q�c�#��b~3�-2#���f}��t!����]�Wd��'�>�5X�{���]�p�P;/��՜ꠙ��^�g����}1��{�f�Vdm�l�K�b�����n}���x*�L紡gp��b��t�9���s��^�(�d)W� G���OJu�oSђ�}S�Dlf���3G����:Z+s��웻��R��
��Ԭ�\�v�,�S�%�g��_f����5�C}hl8%��#�s��`�I�Mij�x�,U�uDu���X"ş5e�s�W����΋��7\����W���}���C��*#,iL�H�7&eO]��0o������̍���+�4�);,���+9__�o��,̣���:��0P�e�;SW������o{�ou��m�����2R�5ګ8�&x秭�ό�BM���k�E��)�c)��rP~�zI������V6{�ϓC�6�����h�:�}�����u<��17�.Z��.�׵r�6� t����n�\��-�q�Z���w�-�,j#������\^�u¯lkb��5�����|�T�.7Pҥ��
Qg\�Õ�,�;��n!���}z�.�)<���m{yo�L���;.u��GSQl�� &�G��Sv��<�����/�V�t5�R��뎞�"�˹��
��fT�w,�<^����QI�j�c�[t�����:%ͤY�+<&��%���<2탟9E�Q>7�y���_��y�'�&�~�[�>u�����\e���ᵱa�
����v���ǽ�^��ɪ{�ί�.J}%.��"��g�Pe�_K����kг�ڸ��JǺ*�{��6b�v�{nzf�I}��#�I9�+��yX=����E��]F�>V,O�|_­q����0� 7�u�=ٱ�)ٯoj�~޻V���9I{i���]5��;7��5]��Y�6�߳ I�c�2�L{��"s��~��8_���똼|\M,��	��[�	�x4�z����8s�N�{�~ΆqZ�
�y+�g
�5]��X�y�����i���&C���]��t��a������c�ȳr����ˁrY4/�p�l�{N,�P�ʞY�۰V�i�վ����}C�82|��������JEh�~`t>�F}|���R�+�KwGx�V��saݫLm�C5��Edu�b5�	�5%�:Xݽ�.�Q��3�UnX�K�s��mJ�.�����Ϛ������/��,�q��/����B��y��r'i��r�`��ʶ�����*ڜܾ�%�L�%t�CO*V%��9��=��ܤ��Y�3m���z��(s�0M4���=VJ�!���	v�����)3�T���x�n^og�Y9��2-���h����w�m_ӽtzu��#A'|��C��	U,�����V��?$���O�����^A-��w�3��5x��Y/�x?���� ��֫�)����=3w˶h����f�g\Հ:���:�ˌR�/��}�De�0*�t8MX�~ccq����MW|�f�n���%�b�������ؘP�S�V٩2++h{����Օ]hl�~�d�߽���������%����Z��I�\1�cǱE�g�t�e��K�"yoR��8/qp�ɣ���TywJ�sɾ�@����IC�0��Ԯ;yvȡ���e'�v��k���<�����{������f�ж���I��I��=�^����~O������tsJ�&�w�f_����z��P�W�llyǄᘞ����+鹸,��pO:>��Ky�p��Z>$k:�)��P��,�����@س�������gW}P�齕��U�pg?���8�t}�ֆ%<���=�����,g�6��c�-�T�)<�[K�2���篶��]�/j�;dmA����Z	Z�|`km���<wu�Z���S��mf�
m���Қ�|`n�����d�mB�5dI8n�t��\�շ����a5�-����G@�j���b_�k�֯�%�x��-ۚ��bY�5�Ws�Gz�׷��U���X6��S��q^"��m��s�쮱�O(%��"������iÇH�,��S)��.��z���^�4��:'��<Sݵ�f�y�5y��ɿP��Ε�b�崮N��!AY���Y�S��vU����vl��J=�<��#���9�ϧz����<*�Q��\��SC:���i���=\��ݺ���0+�f�JǝC7ӱny�Y�%k �i��6�%g@�e��7E��qIj��'��V�18��z���uSjj�ܡ��򌾮#3�sŬ�y��.k�FI��w�oڝ�'e�2$�ҡ沂dW���dl��U2��]�5��vϧ�w�.[	\}B�T9�t��9V)�Ŀ����*^�����XM����S�9����e]�;ýͼ�É�t�@��P�P��P~sr���J�J��S~�a<�
�}���P+�X��g���	���o�����Q� u�=��/E\�Y���z��W,�-�f�ܢ*�d�ے�P4����u=�{�T6�"K�s���g<�8���2��u=�ų�e�](��u��H����#a��r�h46��ŧ�ΊZ������˽���놯�x3�^�a�����!�^F����y"�Kom�c3w,�z���j�5Q�>��"+3�%�wc��i�n
z��Nؕ��8R�%�
��Mr�Y^�OT�(��;�eRR�������ˎҲ7w�q8,+����:�t�t�쥓S1���븸�6Ly~��+g��u~�^?��63e��km@q�i���sAlo+���'��E=�aW��{U�C�=iYxj��G�c\2b~>�š���Ю8f��Y�5��\�vn�FM��E�r���y������3���Ǉ+�C*PE·��AQl*ȩ��:����7���#�e�.�IC��N��S%i�^�U,�Pi`[�LvR߷��tV���� ��w���11ZY��Z�~].��r	�z`��"9j��������u�;gfe��wm����C����@����k>{��mNP�N[��ƾ�9p�}���̩g73Ny�\��l��(�&j-��3.��I�^tO��M[�쳀5ﾉ�������]���f�����i�|�k����	�����f����!��pZ�{����-��8,���I�ԣ�˄vact�B�L�=�����B.�=��WcM��,]�E1��Rw�hpv{s[�z��}���#C;vc�e�F�_{���G<T9��j �"Ŕ�D���|���U�ӣ�}j��@qMM��u����{8%���G9���r�𝈎�72��M.Ӯ3
fbt��q^�U^a�J�9>��r�3Hw�ζ=9�f�&ʲ����M�+�u��d�4����ּ�p�>g��7[��I�6Wjϥ;���W��R׎�7��^<��Y��֑�+g���9�DW.��s8��S�+},���c<ZWl˹��H*Ό�!�Wd÷�`gH���x���B���8E1Zϑ��j3�]̕ҭx���J$����t�˶9E��1Wg\7�#�s�w%�`�ѱf$O{P��ܪkG����kbÃ�ZJ�兟mͯy��T�7�;�N����V�ek�x���j&�+E��K緜_��ˏ��r��-��|�7cTڬ�v�V>˃i��Ѕl�P���Gg+Z�|1����In�:U�/o�b荫]��qym6;�[�O>U�_��Z{-< {�`)6ɺ�-�n��fmk����jl���׹��ô�e63{�mZ��'v%ě�*�
�M�j����q��&��t�lq���Բ�#Q�3'�'���@����0ۑ�T&HϷU�ӗX���0z��1g�um<�gjAY���Q�fMݺ׾si�=0mŘ�z��|1c��o;�P�a9���&*�+��:Ixm
���5\�ጹ�Tk0UC�_�
�7��EU�5�u��|�[��dP��V��3����}�^v{�t}=T��Yȳq+��yp/�M_T$�.-��iņ�P�V��靫s&�ʬ�f�ּdZw-�M_�r;f-Lt�V�O���/q!��[��mҗ�=N��s۽��(Nt0M4������VD$�\��O)W�]KN�C�{}.�X<x����0E��{�i;mx�8���s��"[S����'*��V�ǖ���L�l��E;r>с�i��S��Ը^�|~c'<�/���-�Mv+�߼�۳IMbq����uw����^D�D8��(6�8Ѓ��o��%�ک��mǔw�P�>Ң=^�{ٰagm;�sjc�toG�\"�DӔ�+�du+3��Ca�嵠�foS����i]�[�㝢�y�_d���i�C�W��@k�V��{��\�३p�X�������|EP|+��h�v�ע� i�Yͩ�woV���5���/p��<��79흋Y��I��"X�wZ�Vu����] ����*(�g�H�.NofV�L^�����"��G��F����@�;E�U�$U�o.��KڛH��ú������ᾬ���Χ��j��]%f��W�N�`C��vU�G[�nX��n�-�E[2#aX3[�3[�w}A�1Y{y�n��RڮE���J�0Q%�/��{��Gǆ�}���M$t��ZK/ jq����nG�2�pG����T_L+���1YF�q��2w[N�q�;6'^]e6�4�w"�-�;��1��iV��ٺ*�nx8mX�3�:��|w:ĝVz�S����Fݑ�F�5� ����Cq�	a.��I���e����F�D���w����I�J�.R#�>���(%H�v�M����S���n�㇗<&�a�b5�U�<tR�u�k�wp)3uLTB��8�
�:u�sp^+���u�u�}0�Q��1���6�Ѱ��|0�¯YG�i�����g9{br���o9Eѫ�مԲvj�u5[�O�{�؁Kz!s=��MVUZ�p��v):s�H_�U.�
����K}c���n�'miV�r�o�x����M[f���C��NAg��N�
V�;̼G��Ӽ��ʥ[�%����U�U��tPZ���%f^��oT�"�g�ӈoDL���e�v%\��&�nf��
���Iy�p�Mv%GL�:�
\U:T�Y�u!�>�*0,ǀ!�Qp�eM�v�z�!J�*�W_e��_\�R�#1v���/J��g���eA�ӂ%3hg��LN��cPq�ŷ��v�|ff��-J���5�۷]}o�d�7.��f
�k�Ʊ���þ���[&P�����B��Ɩ��q|�让lFm'�j�&�V>��T5hh�u��J��+��E>꫸w^m���1�a�ʳ\��g�vz40=�ә$�6�r#n�cz��_w
�&tC�7|YO#��nL~��b���+J�/I䭱R��H��L�Y��p�rhާ�+z�����Ne���*z;/�����˓�ê�"�IG�\뼖{�ܑ�^�ͺs7�����Gwi��Ҡ��T�ϖ�غycsp��;!�����I��Z�K\��` X�m��n�^Z���;mF�u �Z�kom׸���i�Y֝�8����d"IAˬŜ7��s�x0�N��2�D3^�I�8.��n^Tp��U����xq�}ZnۊB¶R���L���𱃉��t�8�u�W��
�JQes��:q��+�R�T��Ț�E��������O7�}0gJ���]Ƣ@����]=Ӄ��;	;X�Ѐ��ad��[�u��{��J-	��� v�R��_0;��5k�)q�<1\����wAP�V�^�6-���Ǎw���9�af�|��~�H$AD)
�1r�3,�2h��̲�)¤�# �1����B���" ȣ$�2l,��#"�0�)�,	�"����̬��!�¨�(�3,̲(�2�k3��,��30�l̀�h��"�p̲� ��2���,"d̰�#"�3�ɪ�&
�ph2Ȭg2���&+3(�(b�2�*+,���
�"i+,�	�2�3,��'3,*2r��+0����b���0�L"��0*���
̌����!r2���!�ɣ0�����2$�bȳ̈��
���"�((� �&i�30��r"����h�� ʌ����	���0Ȋ( �
�#0Ƣ2iȦ����J*�,l̪�3'"�0������&ѕ�%��V0,���#�F��+�hX.�S���d�`���k�i__
ћ�����v��k8��)fM�p<^U���o�����0s�G�qO-�K�`�kn��O�E�n���b�&}��b���K�U�x7���u�~�9X��WL�BDD��/TN��
�϶θ��h��an���f�(g�yz����{���q�9񘞥Ү�f�4,�]7�jf%>x����<�};e{o�t�7����+�V<��2�����_y�3���mxX���͈h��^�z;c�i��n߮|��,����/g��(���mӡ�Q~:�4��_f�J��,:�`%>��%'��5_1�=�\f+uO�Si�p���t|�NO�KX< t�h���j����Onԋ��d����y\u�g��`���m�Z}Qu�����W�f��3��T�v���dXu;�ԛC�N�:U���erJX#ԝٱ�]���oe�y޾��kOD���뒱�Lłn#����'z�?_Wpj�ug���)���ą{���KSs���]l�
�� �x'����ϲ�IC�ϧg�N�Q��d��o�G���7��H�x�eЩ��%��͛�~��+-��e+�a���}��܉x��f��^uN}Yţjν�؆�,̡'��؛,V�=4����r��5z+#ۡ�U4���V<�jt�M�����0+ͺ���U��2�d��OO��qպ�z�5�Q��Qd=�����a܃׿N9~ْ蔹�*��ѻ��_���[�zȽ-#r�s��.$�ҡ��	�@_����~w,�w+��3��/�e��#��X���'��9���Y�,L��@۔�J�W�*�	~��R�v��������x�E�;���������P�����7)!c���Ԯ.���x?�����p��sy%f}�Oz��Y�G*����
�G0�˻"u�lk+�n�xW��+��v�D9����+�>GGY[H���<	w\��-0l8)�9����ن�R'�0�zY�G�ܱۛO���f�\Oh��Iex/�z)�e �,+���agUg�ҏ.���/x�bMw4.���dQ�9�C��ko)��Vg}���8V�czye�y�P�aj��v�(���{��Y2�H���85�֫ _��u�g�r��U���'G�;�3{y�]�n�Q�򣑼��<��]雧��=
gk�{q��?*
�o������B�-Y"Sh͡Y�q�6���t1d�{v%>�U`
$of���>��
��{���j�����j��[�C]��pm�ʾ�
[Ͻn�dǷ�<�W��գ���f����d��bs`�Ò&�1���0哝z�c6y��ڂ��e���,��e��ct�9���g4	,=C��t�}�����s��¬E]<�w��Udyy�Fzt�Z-!��M�=�KK1�KL�t0�t��d�_T�Q��o+�n��:��@}��ӐUm��R��b�֢^�4�=�a��(q9oW�^|�랿�jd[�7��'E����vZ\��UCqg�U�`TG$���?'�4�mٟ)R����n�{��켥x�њ�H��V;��|�"��S=}Ip�|��IV�L��Z�\l�W'Y�~�� e8��y�؟Wj�@���m�c�:�6����{��A34e;QݦW�"��]&V&��h:�̈�1�x9׍��g�zz�,3�	sl G2�/
OWl��fz�v:�\�vt����TK���_M�O����o�`��%�3ȟ�M�Ǹ��I���Y���NGC���v�|�����E�S�?w9{�Y����ԯL_��/:>�'ǖ*FF�P��L��f�~Qu_n�	+�!�T���6��5ܪ� ��
��[��ê���{���t�N_��r6�\���W.�����]*�Ŝ͊ɕh��B�84����	�.����JKѽ@&N�}�|r��jaD9�n�{��m�렁�˼r���.����u�&닏%��;3��kv��6�O�vN�喡���INDS�و��v�z�_��D��6R�&����73��}b|赩`�GU�z�BWϴ���._K�*�iZ�<4q`��h{�Ζ��y��
���0��P����Q�l�`�nV�8�&/�Y�pXk+ޑ`༚��6������!��Y����{~,�D��8����aw��3ϕe�)�[��a���h7�-�����b��]u�*��Jy�b�S��w��*q�����b�ҺB\�~2��ƣ��r>q��W(6���	>K��Rz��?��>2�����}'Z�t}�Sl�!8fО|i#�+�lz�}gc�t�g�J�񔼸<�_9���"_u�c��<kz�s��@R��7�ʠ�Ǻޯƙּ�N�	�K��,�����\eJ%ڍ#Lz/t�Ь��v'���k�z���(Nt2i��^�=V*Ȇ��{SEq~�y��ԚI'�����J�P��7L��h�����DK�s}tw>}�@�0�4uk����i,ob�x�:;Wh͙���tS�v��U�'^��CF�#���B�ѧF��!R�D7-���*� ]�3-J�c�.��:��Wo)U���f>
�y�N�u�w(��ّ9r�:ۿ{=%�Dȅߵ�b\ W�l�UJ3�������z��0�B���~���˔�d��9�׊0��k&g�f�,6��Wy;�q1�D�"���^q���뚱Ըu��>q��/	�1n���N�ٮ�wv��Vt�~8�>�K����J�!����w���`,��u��~ܳ�
�)�s�9^�_-��<�9`�.�뤯�#�]J�)&w�+>=c*-��\˱�(�ұAz�N�������T��u��rW���D�u�>^Z1��P�Nִ��P��Ѧ9�ѩI��������U���5��p.$��Q>�=x'�^j�{��!.�%��+3��k����ؕ�=R*�2��>���y�������Y����r(R~vq2�b����7��R���˷l��3�w2�j+l.-�����|�d�e��-�|��jo6kY���7M�3���7K��`�Zܻw���%�:�+�t�V!E�\���P���]�iЦ�rϼ��m�{,��Lv�*`�
މ������=f�m˻ޑT�v�������oh&����Yt[2j�����e	t�)�TN3�4�ň"N)��>��=K�� ' ��YҍREb��*�4E�Tǒҝ[j�R�5���9Q���d��5��↙�S���8ԕ�Զ'�;=���fF%\�徧<���:�Pzv͛ۧf#l���r���47c��w;َ�&N�����S�@Ԟ���s�n����G�uaV

̆ǯ:����:uKg��y��.�<lc���:�)����0�s��	ƞ�����U�jL�ǔ��m�S~�^|��d���v;>�|��:�l�F'�e�P��׎��%�����X3�rmve�,^2Z\���x�G�ԇ_�/��uSjj�ܡ��s�*�Ԩ�;fM�U�m^�癗�vO��1d�V�	�t�)4A�x�Ы�����p���b�Xxb�=��[P͕��)������[�����Ô�IE��P���K#_�y��X23��:fi^�	~C�T�����|.փ�<�E��a�뤇B�'R��ˁ#�Koט��{5Q�:�P� |�u�/>u��][Z\
��W���� ]K/�|��-8���n�긘�[z�����/ԋ�Z`]a=��Qό���=G��T�s\�k�0c�K�)T�)�֕��t�R�S���ϼaj��}w��w9[=E}ȶ{���^��BC4�`w\���#�wK�1���4t{	ܹ.���+ל�����䩏:��$��}��-TaH)}�o
�>��}�!Am�c��S����W;d]!��o�3�eł��x�u�Iex&���� �:�����	j��+2W��yգgT�	ӯ.艈a�:�-���mz�7��ƽJ�y�u����+�k�a�C�����/�
�l��ƑTP-i�ܶo�ڸ���%����gn[{�W����F�a���`�����D��:�
��٣lҠ��G]!{��r�Z�2!ɏy1�.U�<�u�_�c�ړ)�SQ�����NU�ǽ�{}�I%>-&���l���di�P7�p�f,�,�U-C�.�<\�<�����F��F���wc]�7�p��*�%l�EV�/R�C8����;!g���4��]omԿ)�_���꿛�̆���Áu.[�P�YU\f}uDu���X#�~X�M6�4��i䷪Wf���÷N��8�q�:F	�V;��)H�`�z,T��we��x��U[��s;].��ĮP�ۋ|*<���9�]bm������9��0������m�Զr���б^�3��C��i��uuu���7¦Wu����M��T:
׻�ǆi���]imiM,튪RÅZ3#�Vˌ����:)]�is!�&GM���V���V��Q��bn9�m4���+��)�;��l[l�z �-Is�ŗoD~�ry��~�B���jmMHs<q�[�g3��u����>�=����GnC���p(�!��<)��m#^Y���6ot[�����|�z��ze�:�Un�ة��ɧ�+>a��+e$̴'���Me<4�Ǭ�^�oY�{�Vބ�U��t�����#��q��y4��Oi��Ζ8D/ȏ=������*n�����<O�ѷ����7i�wp��b�M���Z���Wx1��c����j�t�1�ie�{wڗ=[��=�b��^Qq�p�����	S�Y����K�5������F��E�D��΅nJ��O�!I�`�M�'kϟ&]�����Ԧ15.M��P���^P��**:��t�qأ��7�h:�s��5N�����F���\W�����U���v0�s���؆���&f�W�]�ݳa#}�7�gs�ݺ	<n׸���J6�iiB��rv��ճ.�{(>Н�'��H�r�{�J�����j���9����r([���:=�k�ǅ��H�p�$�޸��tI��Dl���@�#S����ns���%r$�)_[�ϵ���Vt���\���x6k(g�k��󒧌
�������I�N\����$��M=����)�;�=�]L�����2Y�� �����{}|�3�ۙ�sa�y4�t�]�Y����kՎ�WX~usq��wn�J��3�=�=.���lM�T�O�S��X7��W�bcẟi��c�Cw��������=2@6�^�&��k��x�o���%:��X�R�o,g�hKՍ�]k���"�(�<�%�th���	;�0��Y�� ��=�/-�ɽ�ҞM֦����9O3�r������ؕ�Xb:Ο�U�Or����^���2˖�խ]��i���Tr��T��0�/�U*�sY�a]���l6�����=8H(�	uޮs��Տ�Rʐ�~~>3j�U7/�V����]�ټ���K���Ǵ��D��<�BF<�tc�Ac�����5�};�v���(�e�5����z�&G���T�$WX4���c�[�환s_B]�NH�;=S�}:��|�����*uv��rc�a�ň�-�G�^6�=���K9PYK �vm��ux\t*�ǝ����oJO3J˃E��k�O<�o�,����Gr�p0��X�ͭ�IN�)�����x�|�ęW�K}����W>|�x���[�:��j�<��Т�ո�)���o��M��M4g�d�z��>h���kf�`;�y����v�wcG���s��l�w)}��z�v��i���F��>�c���m{Ps�MD�|��{R��b����
r/�6!��|.#���]�����c��'�0�[�9�����:9�͂so�����Q�B�:,�\�M���*}6 N���GHzt^�mK�{rs���7{v��ۙ:�D�z��<w>���J=�r�ۮx�2r@s|�G�"�z��>�A7}�����t��D߹��:߅>ϵ����������
����
��� ���AQ�
�+�PTA_�AQ�
�+��* ��* �������D�
�+�* ��D��* ��AQ�
�+�PTA_삢
�4W�W��PVI��r
P̀�����X���y�d���jo�	���ʪ!�)J�fJ�$IKlI�T��*�ZTY��J*)
���5�%+MI^��{d�X6�[%e%�*��[-�٫`-b��+U��KV��6JcbkV�Զؚ���_F�3�����2ٴ�6m�1Y���S3[l�6���j�lM����l�-��i�֙eV�lҬ�Z��J�ibcv�t�&Y� >���R�]��Ԇ���q�R��Q���[j�;sn���������u��骔�q�k�U�wn�B��\�զ�keQ�[Z�� �j��
����Um�3�*�,]��PU[��ں��WW8�ʭu����
���Buզ���r��0���de[Xm��ml�m��� 	 � (�Gz�� 
E ����  @QC�� �� 
({�x�  �v�V�!UU�Y�һ�T�sJ�R��í6����ݵ�ѽtz���aZ�l����  {w��N�뺻��*�p�j�e]]n�B�Gn�Un۹�v��k]���u�5Qu�];�mR�9�
[t���k*Ҷ�jUV����  ��*�W�ܻ���Ea�榵N��r)jڹ��$J�v�В��p��m� w:�np�х(7]�aZ$ZSZ��  �����;��mv0�7]��X�d �	B��Gp��cE"�ZUKd�G�  �x{J����3��F����n
M���d�١�j��Ν\ mu�ѱf�H�mY[c� v{ �b7��n�����u�EV6 nv���"���X�vs@�M���m���< ;<h����ik ��48� t�*��ܶ����뜐b�@].S5bͦ�-5�i� wx�@s�p*��n�����0C�q��w.�U4�l�j��1��U< �H AEP��b��*i�`    M1�C��       E=�&��J0 L�  10 5O��IBd��#0��$�S$��j'��(�=C� P��M$��J#&���S��ѐ�4duiéយ��Z�R�j���8Bs�*Ӌŉ�I}�י�O?h��$!�i���0�PB���Jh � ��$!$!���	!�7����`�`��?��$��jHA*�$BHB��d"��! Iv��~��-�޺���f�aA��q�����K6v��	$8�7�;[lu�֏H�hE�W�apM8憬7m���92�y���Ջ�J��u�����ڔU橛ylX��V���U�n����X10a�\2�ɮ�҂�yXt�ϒV�����k��cգ~EK@�FU�V�+��l�����:�ق�mޭ��̲i�r�r�v�@�-��J���W�t�ǫZ���7��n+�R<ǡ2���J��*e� ��P�Z�[]���E�4�]�&�e0�M=���J���,�93�T�5����i������=N*-:t*(���r�pl��\{70P:�İ��Œ�mk�)�Q�N5��&�����m��z�]���P��'���T�3I�q���zޓb�Zn��(�2�f�����`ʱ���V��1��MQ�ʡ"�c!�⣚Rj��(���t��;ϲk��^25��/㔮��U�t�Eko^�9�s2�i1��/0:K����aU�-��O*n�t~wrԇ��&��n�76E�x�C��ҊX��2��I^h7L͆�rTce&���Ci�;m�����x��U݃���R�@cF볕[%`��R��#�+2�Vn��B藤�Jȁ�N�;{*P��K��J��;@�_e�ᷗl2�2�$'��!����m(n�0]�w�b�7�㚪�t��9a���0E'�#`5B��q�a+��X[2ޓL�q���T�� %!t�Xa�Op���pM�5S���/�ISYF��uB�4��$�Nf7K�ݹ�,�Df���U���P8���[_W�I+��݅>T��ڛ��v�4hM�[�H5H<5��s$ʽaTЬ�K0jp`�߱�b'&*�r�@�E����c+#n�XqnO��[���g�oI��0�2jX�Jb6����62&�kN���`�rF�EiV��M,�z�lYnEQRxZ����(f޻����]��a��-�v�^�`���z��6�����f�Ӭ
����d=��P\Y�0O��%Z�j�&-6Kd�p`w�!��+^��6�U�{�B?V��RE�Fv
V@�%�=U{�>�x*���fT�H�v��
aۗ�ed�Fd�Y��.�����7l]�l�,��z�h!V����[8��j���ڻ�a�К������,��ۚ��5f<�fd�*,�Ԩ�3E�uLn,!��n�� ��-�w�Y/I�x����/u/�]�:��Mʂb��.X����WOC�(��m�u�B9	ר�7���%�Ss/~ �âKfĥ�nJv�0^H6m��oD�iY:��2Z���24kjC2 "е�[����M�G��������[�aV����jlaI3�J�D\�2��M���#.൙Cr����c6�n�+߳Z��w�
�0]�-w���U��y�㷆ØK�Ĭ�sPb�.CZ�^�,a�S�)�6�5h���U��# �y����+-������4�7쳹+n�N��-�h�M(Y�m̦q�"��$�Z;8��T��Sd��j�M�T�S�oh^��*�n���U9��t�+U&��3n���Ň�Cm!-���՜�ȐW72T��9���2�#��05��G�CA8���r�Szo2���dnK��Yn����	���ux3\��N�=X��]Ȕ���ix�V'v���u֪\%4�a.V����n��ݽ���*IT�[��܁�p,H����!Yh�z%����6]KU�Pw��0�b�	j!	]���*60�2͜���]�V�\�0m��ڂ��ǔ5坛Uv6��xXۙE�!�ػ8���Xpjxq�:cSN��&�P��ϣ#M+T�s(�em@��k�Su�v^���T�ժ���j��A!�1髯���
�U�\�,�aZ)��JJjʷ�֗��P�K'F�M�y-T��
��Z9M��VXT��%��mm�('L����b��`��e|�#ٺ���H�͕10a�]1[u��$��(Y�����e�3/.U�ޓ�Egc��7il���`�F��ۅ���H�D��ĭ��ձ�"˵yxo���f葭{�O�^�4���6G��e�t� �Y��&�"� `�4�\�:�������$��d���WH���x�k(���5Vf�cvP+wi��㛪�P!S6��q��Z-[�2
�ҥZݢ�/*�	D�"�Y�a���77C��Ʒh�0'[�����e-�ƫV�YcF#%A�B3Y0���E��Z����U4cYO1۹*)��shD�a����ɭ�����0�����enXD����3��J3B�s#��.�u��P�2�B�	1y��Q&��1V���-M�5<�oH���f^]׌7������<��5�!��Z`���mh�bڶr�j,;rV&l�^H�^R�xh,:٭sP�z%ở6�`6"JF��fB����M��ªIl�[�pЕ����M�nÓ
��.tP�7h��R��ײ+�(��r�H�,�7&���lV�K���v��T�ͽ��8f;q��vwU���n���!�cʔskP����B��c�R�0��J�~೑C.݇YIjiY|/����Xƛ��M��ƨ^Gm<�Y�졵LLW���0�;y.Ҡw\�1L8sm�L�*�LX4�^�L8���b�*�-RUi�:��P�wEf��p�vjdn�M��j�M�)�1Z��G	$M��2�yEn�n=�#(TyV�#���P�gY�K�j��a�p�]ַ��jw��l�q�)IL�*�j�Z�Pرk�q�{�:l��E����ӻ݁�h�1���X���'B訾�R�Ȓ���x̭�V1ܱ��*�u��rT�U�ᕴ\9[M�X���@�X.�{�wXla��"]�S ��Ҏ��z�n��Wd4�
/�S�4�6���D�b���6����ɇoU�ڃo ����n;�m[� �7a�Xc������,�u7W8������ju����
z�&�}�2����َ��50+v�3���A\�"R�h4�ŌKt
���K[�
�03��v�U��iT����I�0ܱC\1UϦ�a��Oq�����v *�^ͺ��s P�b�a�kUnf�S;aR���[�\��z�4�w��P�J���p^J�	�R��ӭ��ShXq��!�t��ܽ��;j�&'Y.�:�3��](��Dd	��k+Q:gś�ia��a��n�.S�ɉ6oAH�Z�Wm�)C���Cf=seYƬ+wI�d�w/�GDJ鰘&�|w\�	�4�hO,"n����Lo*�n�ǴОI�~��=�p�f�FkdE�j��8�
i�����Ö-�b<&j��q�Ljſ%�r*)yM�T5�,�m���@F�8��ݭ�@�%���&5V\ݨ�ңrhW��*����.+���zu^�{�,�V	6|�m^f�-<&V|���I�3n!�X:w�qсڭ��C�a�Ya��Yc7f�E",�5�5�Vh���bn�iSV�nZb�J��vz/yo&�U��fm!��cuz�/JXм��h^����^\��t�`Ru4�H5JcCq�ͤޣ{�-��$�[���������b0dr�1�u�u�i�v4����7z�� �F�%�yv&5�1��%A��q��1a*����j�U�a���ҽ;�
�[���wz�#�R�0L��1;g�T�"�"̬�eUH�)�dj��Uy���e�{�c�]�iU�u���-%b�nY�/wA	�n������S��G|�c�*Q4��gl���U���{���c.��J5��[�U�Qd�u!%ݴrM�յ�tKqEw&��+,Pύ����=�6��$��Y�bm�M�Ӛ-����CD��yB��-6����gTm�R��E�TV��y��z�aE"nH�6���F���Z�Z��2�bv�S��Rv	dH)\?iѳP�Ot'cjF�!�Gt�<RC&��1�5J�d^��(]�+[��y�-�WukCIR%�mЬ�& ��kS.�4q[���J0;�aS:�a��aYV4-S7Kx�P�ʸ�U����)�:���o#z��Շf��5�-b5��J�x� ������w%� ���V5�
��fV&0�e��^�rk�y۵N�KvDs���Z֔�o[m���[�xeܘ���*P4�����+ߡ�h�*�cm�͙+sU�镘]�BVC�[&����GAR=��5w�-�6���J识��E��mF+��%�����)b�^ 1ͬ��a��Cl�6�����S�3��9�zС�m���r��z�m=�`$u��b���U�sP��i)i�MLR��ҙ��+b�11-.��x72�e�����RgB�DY��J�Lvr�Ml�)f�w3ht�:ۡr�R�d7�3�0��V�[/,Wz4���`Uu%G��ۓ�.(0�k0��n�CR���G�%uR=xrHM�h��+T�w% ������^��M�9�p�L��m�y�Um��pkI�J���<�M�e(b�lձJ�ce���1�b2���5vT)/�Rl{v)v����л��U�B�ȰX6�h�O3��[����qBT����B�f�yO���+*�	�X,b��.��L�r�5U����S(�[eJ�0�N<ݭĘ�-�r�h<�՝4��gh�v�`8KK�j&�ep(:gB��.�nݴ�dyXYyx�FZVZ�ǹ���f�.���e����=*��-��[Xr�R��
Z��&�0�跦�0B��*��ʹ7tŨ���MAl�����J�ئ��
;R�e��j
&�ٵ��Ħ��KM��Tq��s	E��Ux�x�q�s�n��{']�aYA�-P��`�,V��t�,,[����l�[�Է5KT4LOhJTy.�j��� �Qm���m�o�^�w?��3��Y��?�*v$O�~�ե����c�	�ceZ)ҵ+Vj4k
�q�^Q�z�Eo;���dT��y +�+�t1u-��a�t�K�;�R]�V��A=���]���ъ�� SG�9�ec;���E�\��G�:/��<��0���a��+����J��W~uisvFa�;��7���%ge].�{��b��Hjζ���)c�����V,8�d�X�Np���Ř6��h��wi�q�3(�����4N�Ѹ�Z4�e=�o�۔Ů� /{����?D�>����/��W>yW���t���*1�ܹ�`@a���'���/�����g�*�R׺������E�Xj��i��5*�����Jݽ9d,.�Ne�zQ�7D��#]�l���>��X��?$�u�ɻ�z����<�)[�j3�����+�������#:��a��%��ݑ��.Le�\�a_um����u�P�(6�=v���ԡ=t�;�]t
<X�o�{�"�S��u�K�0�7�Uly֯�����g1�i�!#���A�h>�� �lDvQj��S7��F��%�K#5MV�g\�l�B�4�2�ë��	���� M�y�i�H��X�85�����OB�M�bm�)K�to:�i�|1�n�����V�ﺙ�)r{�C�	�՘�΂�C��`;Y������hT���ֻܮC�GgLó�rK��������I��t�m�׳r��X�-���m�P�Ge�Wq!æQ�������>��Qk��+:�#^�3dkY���X���l���*t��[}�>�^D�o|)2�f����*��bV�Ooi���wU��G��Fuu�ͼ�3	���������;��]&�F�i
�Ӥh��;]��a�2//�z�U<��cl��'}���K�����y���(
c%��J?D&�w��ƜvT�%���1��u�F���N��.�>��%��e�QITȻjc���̼�N��jMʸ$�{']>���ApB��6N��A̘���a[c6͂^�m�Uh�S˰�[Z�BS��e�lߕyo�n�M�����s���6̼::_`gp�9�]�"�\t��j)nA���Dc`<)*[�է�U�R�1*xzV5�?�v_ �$S_}�yJ� �����f�NB���@�.C��Os��)%()�f�8_l�:�-m"\J����;�|������᥽9J=�DK�49��`�a�����,e_<To��G3y3�n` 7�M98E���1�k�#ӎ�(�<�t�z��8�a9\�4�opv�Nyo�7+���`�6���3�lZu�L˚3�][P���VwQ�;2f�x��SN���/+9��R��U�9^����Ai����?w:�ԫ� q�u9���N�q�����,kg*�9��0�M|м/6�ȚB�u��v��2��6��hw�Z��u���h۬���:��*�By�� �Y�.�,�G��A�X���Fʸ�w+2-���m`����,9t0MU0񻽵��Ԯ�\-.�J�s|{��s<�:�c4���՜�]$���]�����0*[�RKW���\�3&mn��VVMWC�h�R��[D#ȒB��Q�Le��,�(*��oj_۱>���������3{�3Tօ����ip�܎T�w��8X2��#�D����L�FϟA*�������]�@��}�)��|��i�G�<~|���(z��klY�檋0Dh'��2j����5Y��uŻo]�YX�P����VEr���K(�j��v�R�(R��#W�tgQ����D�V�331-A���,����Ӈ�ఱ����Z�M���id�x+� �)��0%b����7�,�n����\�f=�"���r��`:�	�c���f�ȷ�obWή�a�%c%t7��:(D��#mU�љ���Q�(u��1�?u5�-K�2Z� Ӝ��1� ꅧ����[j�ᒖp�����V�<(�j�i��o�N���X��87d0�S�Z��c�)p"<h�q9�@�� 0�M}YN��sy�	>��O�n�[����۠���Յ\���47�+7�L@ʽRj�kIBM�C*th`]k^�[!���4/9ל/�#�!K)��:�5d�b�9`��9�}��k���*'s 1�&^<�EQ����mv�g�M�ZTn�зR���;�ӔTݝ�q���%��u;4���
�]r5��8�E���R��)�{��ɪt�O��z�;FgE-�ט���g:��ڥ�΋Ύ�f�\�7[����ʣ�vo�R�i�Г��U�!��z�-���V~_m�{�L�u��So�ِ<友��{�V�ƈ�)�v�!���'��)]Y��e�HR�!�wPw�h=�;8��t<����e��f�JZ�NN49��{+2G'p7���]�N_-�dL5��}�*U�Dо�Z�˭]A�����ku$��i�3���WY�'��J[���h+���ņ;�.A��dYf�����p��(v�I0ԫW��6�C>�+&-�B𓕅��}B�[�qS�<�X4�t@��2Tۃ�ojTɑ;2���bu�0���g���OP8�77:lܡ�E9���O��d������i�����J���#�	r9
�e
j� r��*��x����}x�
U�wH�{gpΙ�{�w2��J�Uu15\���]�9ѥ/n�+t06��R��T>���㋒�v�4T����c/�g2%��OQ�ɜz���;Ȅ��Me�w�X���KUi�T:(�s�[��w{���;�e�WDz�95���b��ް�Q�Մ�	İ�OkJ^�!�9�!��Y5|���Xɪ�!㓜�鸳fQ3SV���ڟ#lM���S��Ι���*�V��5����Εf��*�\����sg�U��2m��ʳT�i�Y�v0bWw�7S��z�7(&���]R��]��S0Ei�ymܽ��,�npNS}l��*i��2�Lp��#qV]os��A*�p�V���{#��f}$ésө�`	�;7����=�>=6�h�m�t�AӀv�pG��.�=�Z֎H5j�Tk�����K5�\��EN�J��¤�6j�!B���ӻA<�+���d
�9po�+ɎX��4Pe��q<�g�D;#x���ʻ,n8��#�VA�Jq�ݙ%�=RdC��6Y�y,�����k:R�Q���5��_ڴHY�Q�eJf����I��3�T�v,)1es5��.yR����=U-9���驥F��	Z�{N��;V����> ��6N�w�+*�3�Fի�3c�a󕼺�A��v-�K8��t��^�}�eރt��c�9G�:��[�Ƅuk�Ž{��-��r�ڛ+5�MԓGw`�t�;�_D�f!U�&8F��U��9��ŕC�V�;�un��Ĳ����#*�����I4�>�
T�P;�]�^�d����q�do+b�r�iq��tx,���oI�		�m�²�Y�z�Jʈbc{�QU>�:��hA:$�Tm�6]
죝�<����+��|)LSk��*Sܫ��er/j	�D���U]}�X�3��ʺ�Q>(a+���k�\���F�`��Aݤ��i�,��?$p;�-���o;eյ|�i����)m�bJqN�u���̀�nu;[q�T�Es�a��C]�&0�nT5Z�������sݺ���X&�|��s"��Τj���ּ$�5�\�y�c��ٹ�9ʆ��.I�U��9؏�4L�9�r��Xq��NT;�p;;[��NjMںC��Ŏ��#����x�GV�-m������l�+��Ƕ�yR�{�D���aOՇ��)�R��eX}ռu��3�ة�]:ޮҝ����5��3���|#��V�f�?X�M�vV�(���7q�<�g6�=�B��[�a��r�D։�do��v�<�ܺi�4V7SK����ybd'-C�Ԥ�6��$Մ��S�ƊhN�/7;r�7�"N�b���
R���-([ܶ���#��P�.4��3D��E���ȄT�s�N�ܼ�L�=��"���4�_`5�����eH�B7h]{�lP�B��qRd̲�u�e�t`�z�,��5	䶬�F�ve@46��@�:؅�֨�Moe��t�"����:��י�q��G\u�&�Ȇh�;Y;��%%5eP���q���3J-"6��OX4�	ů���D�[Y�����1��ۙh��q�`�������8��̰��1Y�����yb%�}5��et(v�v*�M=����;��Z٣QV�["t��ָ�����ɢ,'.o8V�ӰB�����H��9}S����̺����UT�)��hgk;�%�8�&<�y*�C��pN\ڴ�����l�BT��͏�Y�s�YF�i��s�MS6)��p�7A�����y5�a�+�_lo���@ #WϾ9��i-2�U�F�%�\�`k���vސ�ĳb@�CK��i�퀻'�6��k��L���ڶMU���^X��-�4?r��e���ԝ�F����˘�]�l�U�>���oø���u������B'�k"�]�E���iq�LtP�ԍN�R!
,0�͋�3Zw�1P���P׉&P|��nM}v,����l�%�V�N���=�Y0��Y�*�݋�ބ�F2�%gc�T��,��3�sM��xnd�6á��Q���L��}�9I$�I$�I3sz'��/T��(7-������c����*��zf�[�묉4�gjA���rW2X$==��3.�=����f$4r#�;���Q�w;�h��wt��9�ua
�%Q���FI�"�l��q�8���Z�,eZ�i<2]���Lr���<�l�l��9�sbÓj(��nl�j�"��s���b��E�,w�u8�fd��)Y�t�e7{و����l读"� �)�u�uÎ��iH]���I ��b�Y��!$��㿰$�'���	 �W�iQ]s��(��ý����J֥�3��k��yU�X%�Y�w`-��fv�nl��2wt�Ĩ�O�nfA��G�͝���fm�o(q���YN�������:�k{R2-�1[�2�ue#e:���-��Q�9/�²r�>��u���H�
��NV����b���䒲Đ�g�N��շ���1	o�,&�Q�F㩻11�6i]�3B2e��u�G�;��
ɇ
��D�՝o�^�����n��`�W}S������\����bVj}f�(u�ǳ;7�X���&�9�O2�rҞ��a�b��u훮Qf�b���j��q���IMu�g@���8TE$���Z;�;#�6_]O
��1&r��TS�"�U��d�D��v���h���;�A}�V@�]�xʺ�I���Щ	�5����a�t��� Ů�0�����Mݢ6V^(x ���䶚��'z�r�8R5�sIVik���bX&��'�vj����F�A�p�r�=�.T/!+م�j��j���A�4=�o���Ł�U�e�8-��S]�ﴟ�˅���n0�V�)},��6�KJB���r7*!�\0 ɼ{w]L�u̟��vb5C1��"jb���B��v��Gu�E�����4�ʽ�s��)�E�\&�7v��s�v^�PX)�r�u���p��'�z)�D�X��W��O��#3�U��Q|�u"�J�{�[�"��.6��H�;��4��i���<��(l��^l�b����"���p�]�p�U�e��(��o�?%�Ul�]�W�T�EQB�d8�2�J}a��'1��`9|N�_�Z��c��"�P�V��5�Xi�m��w�Ņ�=�,��lm�"c`��QuŰX5.(�Y[&�V]��*�f���u�s�է�e�/#bn�|�\�PQ�k��P�++.������)�Y��)�ʐ�;�oi�9:����p���'�d�]�zqv��	��NV�(�fQ��L(�{^���Jp6��о�t
f놥��6�h�IVa��m�HȞ�x�f��+��qo<�V��ff�z�7M�X���I�@҂��`)b+e9�R�׮��[�Xz�uL�w3��|��*�b'�>�)��,l�X+hg$���eݭJ�&��91dcRG��t��76��$�l�e_l��&�� �EL����PwT�d0��$acI:�wC�8�@9��9P�H S����Ŋ۱����y�wP>&Q6��bs��*��V��ր�N�I��P�E��_mDD2���Cl�'BJlRH�vM{�Jd��/6����τ�++h���7�I�z4�)V:s��mʘ���@��'��8���kC9U��j�i{��l�Pc$^r�5/�oR���ɻ�<�5���m��v*45ƞ����7�O�T���R�ᇥa6�������79��@�6V�*[B��)�%=mnAp���}̵��dQq��D,��tJJ92��	

�C� �iw�]j���C]JѮ㡶[�r�X�.`՛�N��)|����{��7hV�h���f��O�*N��f�%֤]]�ajRWA�i��6�%�g���5��̻k��ET�Ub�v�D�Skmf41����i�z�	���2�pw<�z����jI����NFo38q����e�a�Z��$����:�]��lnnp,�VA!1S+>��c��ǛǍ�۬��)�}y���ɏ4��|�5�K���[H�=� �f�Mw^��)v�L�/{����b�wȫȎ�%'�����zV󲓵��1W �S�f��������]�v/�7�6�u����q�,껇/�Z.����:M�+�*��ut��ə|�÷�K�bC�:���PU�k����3*����gA�����Fq�:��CY��YB:��Q��rhD�N����:�xA�{1�#,l��G��m[xUm���oY郮��0�嫘���Hj���YN���^�]�dunKҢ���y[{k$�C57Pn��4��D�ȟL3�:���6�Q�P��er��J��!����EuS���6uıf��B%`ä9���v1g)�����w�e��)�R�۲�֐��(��=nK�<��r���q�lv��S9d�Q�y-8(�\(S���yd��X��uF.Ң�����Nx��=h]e���=R�=b�WN%vr���K^�6��1,��&4�ũ��+sT�C�X�u�i�
�ȭ]�1�;ܪ�їC�ϛ�c:`hmgu���'t�բ��X��h�֔n�[T��zvK�a���;��q�������㿻^ʷ�(r�Z��]и2����\�~fݫ��t��=E�*�lm��RU��-,�f{dEZpY,PE���G�Y\��$ o[v�]�;A��{D�R劏8�b��a����7���p���"���C������8٥z���ͦ��L��ĺ� -����ˋla^!ڈ*=ic8��ͽ��[{,	�$��P��Z�1���Qt�H�:5�5�n!z�|��غV� T��sCݑBGo>௓u[v������v���[��K���D�١$���G������{�e%jQ�.��-}M[�:�LmI�'
���e�}�q˘�Kl[Dӫ�9�G";0�H�<�*/���fAy�tr�m�t�"�w�����sj��L�@M_fZS�h�<՗�A�$���{�Qs=�{([�V2�3�)�3lDr]j]oN�挕w�)��b�A�w8�ͽ�Q�R���i��H��OQ:��ܴ�3)[N٘��ߕ���ܽΧ� ������l�� 'd.��dũU��O 33G/vۂ��̆�����R)��S3
�������ծ"�S��Tw�J
9:�`XU�l���a�5w3S��DX�U]3�(�K,��8&oW&�K��K�l�߱�rZח�6���+n=���ۓr�)���Kj܊�	AUV�b�P�;����P�ە�����XsS��������7e�7�F�{]t��jІ��m�pZ;���U�R�5�^�7
���;NE�D�z��p�T��Fp*n+u�XF�4�+�]I�$HP��%���2���J�wb��ƺ���j�%<�#�oN�<�/J�����>��8hֿ�kt�$�:��۠m�9R��q�amorf��f�OP�5�T9��d���{q�F@��]Y�lD�G7�ڬ�w�����C�7M2�d&�- 2�m]�pp`}�(U��5GHl+`�`��[87��F�F�/,��s���t�)u&�a���qٷ��Zr�k�CO�n�p��o(��Z�L^.���A���w"�ڍ<6\��˭J�r4�I{��{�*�٦,�VF�s	h�vbB���(�q�ˊ�-�9��{ov=��4cD��p��q�2��Z�|���۱�^�(��4n#Z*�k��!Kp���ˣ�vG��J�&%eJ.r{.�eЩG��+� ou����"s��T��7��FÖ-(	p#�Y�}��$[�����6@���院Ծʅ&�e,�E	6-�ە������s����u(�Y�o̂��a��噗���T�a�㽅����$�%�|wS�2�ɲ�)�SM�ЄR����wW��iɳ{3W�Q��\������e���Ĺ7�# aj�8��%n��v�v�Yس��O��h(�IG�}r��ǣ�
-�2z�.�ᶜ�؃�n�^f���XV�4!�nv�������ƎL�N��]�j��4r�hY���H�?E���}�s�qx�w�m�{Om���Ŗ�0�������UAݓvn���jY�G9�[�t�{�w�h����&�!u@�wL������&��{��W���>�Ze��V�8�4�A�<Xr�i|qjp1Q�*;�('�K��m��a�}ʻ�*��r2�{jиS�+���}W۱DF���5WO��i��&��Yfac���q��7��=�kp�D��'{gS6��<���=��Vx�T��+H��d�e	�X�Wʩi��醍:��(�3����q�wës�+�Ru�r󥖕ŧ�.��iEs,�3Ff���]ZY"�:͈�i�����))c#���+���I.��Sذ���S��]@�x�T�F�IP�C�zVh1�k���Pϯw)�r���U8��Ev��n
W���(\}#�Zu/��h��{t��`�J*�D��{w�i�M8]�����p�K�Ո�d:o��sۢ���$v�m��S�A<@��{�p��t��GV�%�h�:�A!e��z�bf��]Pk��+z�M���'�u9�,Syv�7�̑r4�R�4�%jןGՇ����8K��\N�yn0�@���Lm�ej'�������)�qd���ƵZ�$���˖�}�uJ��H�b����N�h|Ƃ�{f� ζ��LU�	��a6�-S�pM�>\��:f`��_�K,�%YDښ��ZK�I1�]��i��U��eӷ��e�	
�6YmNK+:Eחܔ���$SZkE�K�u��^P��}96�W/*�z��^�j�|�����c0���B�T�P���*��7,�u�9��!��<��˗sY�p<��.�1�@�������qx�C�4���Ў��R5���6ƾN��a'���fE�%e�w[z��uf�I$��M���|�B�O'E��0�{�%uG�L�a�|�-�ٮC3VC��^q�����\��jjCh(o�R��[��.���P:�ε�n�4�e�֮��Y\F��[�%E,�͊�-z�89`�rW��=޺t�F{֨�@�R�	�i���݋�����}�ud\�!���zb��Y���ʵ�}�|�$�VE��!�s0��d:�߄?Ak��p+��TI�����@�Ho�,L�C�E*wyQ)�!x�I�&`c0��ҶЄN�Y��m��7+-���md������ͽ��֔��Z�@w10���3��%�a]#�5l�I�Leܺ� �6��c{`v��q	mU�-;O�6]�+2W%�*�b����{�ȳq��P�"�S��+��r[|�V��W���6����t��7c�g�[�����r�D�� ����4���͹�6�b�� ʡҏ���]�+�ˍ86�������=*8t���I���2�[�t�L*��H}j�`�+]�[�٢�hs�Qe�&4�A�����`RLy3i5ڦ�c/��x��r#��U����E�9��T��yo�	�-��Kk6`O3L�	hݭU�7�Ӣ��|�05y��&���`�}���ti�_>p!��v�*Sǲt*�*��Ƶ���U$�}:���O�v�$[ɳi<����Rj�L��V\�FN���{���E`�����5[E(V��m	P�m�l�DEhF�U
�J���)F(c+Ub��uB�-�X���
��Pm
(ԕF�f	V,jYb�"����Ƃ�EU"DrؤQH�,EV(+��&55�TUu�q,cYUR
�� �F ����0X�QDcj$T
�*�Tb	\B�*��QX�D��ʵ%���\@���@c�j�X�,�����E-,b���Z�QU�!#�x��Ӵю�]��s"��m��)-fjf��Bs��a��X�Q�U�J���Li�<&w����h��,F0�Ǐ���W�������b�/���4Q]�p�^u��^p,������7�U�(\��A��A�J6���3+$�MA<�dX�P7.g��H3" ��6�y�����ۜ�����K�6��B�ާ�M\~�Gǁz͠�6��_9�^���;]���"� ���/��P���������a'M���X���N]�a-��R�H�֣�B�dB��	#����4͸��:��B�{{x��� �y�Lc⋗P?.����&3���6�[�7+��	�M� V.�Sb�P"�%�3��A^���s�b����s�*�߱]{}�:�w�o��C��-Q�^Q"�_��T���"!�����g$J�ў�E�!�r�v�K����%V��%\���C��'����|Sr~�i�9�i8��[�\��0����"�����G�$V�d�(+&*��55��:�/ʝ8ˌ��{���н���X�T�0�j(t�n�[30�vA�g#�>��g��hoA��������/t����"�F�T�����N�����z����yo�֯#�go�r��c�Tav��uk��54�$��9j�\t���c Cux��2 �túh&w1�y�@����B�h���!�<<G��,�/��8�.�m�����s`1ӦCr�"`�f\*�"�x��#��oo��=��ãm�I�8�;s��CR1H0��
�9���k�\�i^UjG�0��V~���:�]x�q����eP������:�7%��%���34�X�0	�.���>�T��!j�Z��� �\aM�[7������2�)ȿT�s-��T�XR1Y�Am�Q���h��ǡ���=��8��qAH���0�^cy���oe[�G��Xh�']0���ؗ
0u;{ʹP�w)�������$�3O9X�բ�1�Ee���nX���7��ZK)R$M�0��0���rm��I�}jNչ�S���[���WJ9P�_��J�?\�X����^H��2�ԣ�No�D1*g�f���=�L2��'ڬ{X��1;B%MP�)H��:��A�zS��/f���8|V���а��ј�T�B3�*�
�Q/�KW��!��^���=+ɞ?����M�t�T�e,���|�Ը�o�yA@���N��#Z�fiMZ6#{��G��;��e+�Q����6׬GfV��+� ��ҳ����O���k���u��^��xTBt�h3�;);2��Z�����xA �9�&#a��e����8�R�3F
��^M��N���:�G{[b�r��<챊�D8�S��SC��FS����-	���Ol;hW��h��#G+3]�G
І�$�I����7�u7ڭ=x��ժq���)���}�&Lɗ7�����q-|����$��*�xH�q�,��!-�V�����Y� "�h���M#N�쮭����v{M�i߼���}���AsnA��FE�R�L$\؈�x�I4�� ÇN�7��8��i�zzz׎}No�}��.�S��-E��f��~��|�K��O�>4zž9I�<!=YŔ���1^��,E)�W�#&�ȅ4�r��=�)�{)+�H�C՞�_���B�@c��c��0�_/��^i���=��M�嵚��=,О� �!9�mE�!E}a�����8<2 �I<�po���P5�=�5\��X�f[�#؍LN9z�{Dڝ��Г��>��k-�7�o��l8��nX�^�N|�����e�T���7�+�^�	�}�Q�Rb�q�B���~���F�Y���H�9y����!b�U�Ǣ�96��o�j{�J�]_o����b�N*�6�����qn�{b}k7_�n�
�sp��2����+�V�o\`�j8{4+)E�_&epS�Z��%Ih���xk��̢1Z@^)7�����&M�02�)�~5n}��wȊ�B}�7e��Xͱ���v�΍��_�W1�}�"�!�FVnu�*�"�c8�+c�qP�����۳Ŷڱ�o"C��)�B3���<61qӤYuc�@�;ư�ܺ��1�J���&<�ʀ�tg�V6�������ùe�4:�D׷��v��Q�<��v6<�������ny~��s���b���K�|���Jء'����	#}_'�8�<�?Q�S^(��Z�r���픤\
n���3"�Cq"��X��g�|��|-3�ܲO�9�+�������hv]�(v�b�iZ��b ���ߛC�C��=�v��Ƣt��/ �sܫ�$̩	�FK�Y}�z�a�xlWK�#����N����3���m�/qT"��L(f��v�[�i��6�zv���6j/9!���A�34�=0���Ě�r66��̈́�4�r��e4�@�9K{sn�U���.|^凅IR�+��6O9;�Gu���}�,��v��.0��~�b${P>T9��Uo��Q�ɵ;;>�_��)���<����%zN2��(*>?_v]��vs]o�~��r^���k�!�٬��xV������қ���;X�Y{���t�ϼ��V�!gl������Uk�rn�wW��w%{��hz��D���C�6Qx��Ҷ0v�;��ȃ��[i�e�!Ըf�C� nOxc���U^����zNn=^�6���C�xx7F>sU�����9��L=@`�V6�yu�f���ēVc"o�ΠO�k��A](gD�sȷ!��� �9*r&�\�&8S�Ȟ]� �cR����Vix�1��[��>�Z���1
e�&��뇙Cl!�ϝҟj�܇�p#���X	򀏛^���t+͘E��fߤiu0�[yM�~�B�4��=sf8N��J�.�$�V-M�KjfC�D��cf�5}M���`E��
�ۧ7!���; ��f�� G%|�MrNn���w�*�����>S*�R�f�TxVyV�.-��9�ݼҨ*]H���V�*\p]�ӊ|�[��Pj�&D�a���KW�
yª�PS�#)�������e�U1g�5I�*�����q����p|^/���ψbS��WH��=#�-*'�l@z�u$q��,�n_���0�[A����Μ�^^����IqUqe���N�TK��2�aV�(C�t����K����Ym
L�*�Έ5���➿���h�63%��>��jIT�9�/���>X�ɘ9|wƵ�_l���+�RC�f�M�~#���>���Ѐ�`N�b�Қ�rl�>�*����-D���W��"T�eJ�Ȯ�;�
�o���-z���w�K!ݙ���ufS���~���nR�M�$�;�����Rdç�{���ı�:O���-�`glɕg:��i����K)��I�թ�,��}�G13���8�s���bv�����q���K��m:�!��;���G�0[���ĝ3-��
K��2(��P�2aǹ	뜩�B,T�"F#&5�'K|UکLu ����f�YȆ��ڰ��������Z=�ݜ<���6�y��r7&��H���Y����A�D팕�+����Mb�`l?9���~���Tӛrd##qU�P&`�PB�����C�F�9m�憗�i��z�^5�)���T��t-B����Τ��j87^���1Y�yi���K�ָ�Y�؝�[�4���n�1F�������Z�X��@b4���څO>$��g`��V���fHŵz���h<@�όc��$t�ϬL|s�gPg�kRj�C1X����G�{�l��/��_l�4!�+|�ht���
m|�����T7L���4ዪOrۭb�c��\�;�)K���I��B����]�:2�G��.�<j�R�&Mp[����f�T�т0��ٽ���&�#��ʮ;ܓ3��7�n}�	N��MB$#��e�����QYv���6k�`�0��!L�c��z�C��nX3���艋T���Z�k��E�$/�-8FEa�R���Cv\x������(���J�b�	2(3B�Y��ڤ���X.�Qm�ܪ"4��Wj1�[c��������B h�]����.׼�HP骷d|��A��t���M�C�Ņ�h�Vnu�*S$[�q}Mt�՛�4l([��������Heg�w�! -���.:t�.��@�ߌ�v2�e�w���g�1�.7��päa~�O>�y~4�#7��:;�`�<u����aF� �k����=?O-7���6���!����5=�����w�
�}{~q����X%�}��1!��xD#!�uy����R%h�az���ޞ�v�Jz��y���AL����(ͫ�3Ik�5�o;˺fQ],���-� i�Z�3
m8��[ �\n9�^L5ܤl�7�~�S-�����o�펱�\���q���^������4^���q��l�p�V�ںW�����׾�G���C�R�CT��t�\|!\���qOt����1������+C�C��5�*
�PP3R��벬�|Z̈Pӡ��L�c�.�?�<���<^���數�Z�osjH�ec�b<�L��uC+iD��Ч-�؈�Yp��ǝ'9$�I3��W��*�B��uJ,�[��^<��G
Jɋ�\D7�&�2�Pi_���aZ�=��ℝ>T��Sc��ǩ;6j��z�:���HL{e%؇h_n���3�p�:���ͬ^5h1�D������k����)�/r����z�q�t�%�6�����{��
j�by�:|��w���n��dͽbZ}�
�/��ܿ�~���'G�;�H:17���8��˚gλt�7���SA�|�Ug�EF]�6z:�����0�QDJ���+h������F����Y�x��'����t�4�I�7d��Z��k�V�X��*�j�v��D�ɨݺ[��/�^!;%
0궕b壬��i�$t-�gw�	Lޞ�����9�\��q��B����f�:�_^^Y)J�<FA�E���n�}vE&a��d��Y�$��Y��R��$Np�m�]y�ON_lY�d�*��u��ÈT
�1�tn;���s]u�Q��ٶynbJ+�j�J�n^�|:K�;��b��UnN� wu;��^�r<7�cf"����[t"[}0j�}��V�$ڏZ��Nsq>u��*������ҸU��V����*>�.����ͺ�����r���lw*�\u�YB0#�#�仆�Z�c2�%��\�p�-���G�]{�\�T��^�"p��7����4N��3OlO��4h}�����2�E�V��F]QU����!��q�{YQ�qo�6r�Mю�T�u���}�/n�/\����>My��'fxl��j�
z�KA�f���st��V]�jҙ�.��o��X�Wj�q��n�,	J�ژ�a�؞u�Ju-���������@q�HZ��8�r��luU���Q��9�\�J�g�RXO�5e�hޛ�A'�RP�S�|k�(V�ʗ���k�~�i�q��ǂ���m�|GDȞ�ﴎR�RùZ�c����M[
��m��U��J;���,
9�� ��b2��p)0w:4���ǷF��X+1�?i�:'8-�d�CEJ3�H{���"���k:��v*
�����+��=(OnlBƑ�A���mP�t;���
p��tVx�A$o���V��Ah5��Xh��bKtc��!Mv��LA��zJ�%3.�b��%�ޤ��-�`4��|{Z�)���z��ۏ�l1�q��f��"7���Wu>�s�Z��/	�w�9`���9��듺W8�%I��O��sg!P��3��s1ŉ6`���8����d/^r|e,��`��~�]%�
��UAEQk+�(�����
*Œ#E���QV
���Qm*�*����"��Db �cH�Vb"�ȱ`*���F���0Tb��(*$Q������J��DUQES-�(�TQE�"��"�E�"�*(�E�+-�PPU,QH���*UDD`,Q��,.Z* �*[DTb#� �(�#X* ��F��YF*UQQ��E+PF-�,U[h8�c%��TTEFj�UQb����V�UlUG-�Ŷ��#X��0EkUQm�S�Z(�?+�����g�:$W^�������Ax@�S�Ea��B����>��넮w|8]�}�l���E����O����K�.y��!��B����$ {w�<�B{C;�v"��@��ZgBVEOߦ�������̬0��z�����mz�W�⃂��4�r��"x@�p�L���"N�h���H��ԧ���m�C]t�A�
��S�5(��d'+�mr�yR�qk7��l1�������u��q��r���>	QR��c0���s'e��U�JiȘ0�v�S�2��	����6A���PR�����W��+�T]ï��*D��;IX$�K�1�Ja�����t-6~���$��A���BR�M5���J�4�2�@rh0g��=ˇ��/�U-Hx����:sP�=m^��{}�z�e"U�}�O=`h<`�Oj�v� �U�P��U�}~}��\Hg8N�c��jX�[���X*��_
.�I�~Zrϧ�u�3�m*
s�y�d��3G�f/�}�n���+��khǗ;30�b�y	��j�8��Q�	 �rjI�r�o��Y��oʱ3�k%b�����,/q�&¼��KbB�N�Q��>����,فp��
���X3������ˋK%�D�~�t��쮟]!�U���a��@���=��"���l��̚c���ޔ~�Z~H�\�b����6wgv1�����\Y@9ο8�:#�F��4�=������K�=�*�ww��%����Ld(�d3/g��)��qtV���n��p�{�y8�(�I$[���[�}�1�c��@���ڰ����:���^��]����C#h__�^���+�oH�}���H�M�/�\s*��è�2�tOJ�c�?���y/�]�A\�.>�w�~qK�����,y�t������4��3��@�Z47�Ys��|ˡ��E�j�^�)�Q!�WgF����qS��w�<B�n%����{{)e��.�i��@q�~X5�MAS�vB���o:�]�P��u�'��r���ޔ�հ�rрg�j(w��͗9�Pń���/�2z�W��2(���t�-�2+�ܸ2�ݪ���NX��B(^^���3�3P�nr_T�SI�Y0�{"�P5)OEv� bT�Ԩ����,'B^��܌e��c�j@��}����v8��}������$��V,L�M�>�4�V��L! 2:��F[��r�8GEK-@�{<�$�`n��,�y���cŋS��W���R:�Z���p<���g ְH���Q��몜l��A��~^�k*4r��k�[/oc��'"�V.��r#�����,�ƺ��~t���-��V�[�5��>�e��5�+�����$'� n�rqk��5�����Nҋ�f�s����+��6F�wU���4��w�>�ߡ]�6�L	L�'
֛Y�r��3��3q����~�nx�K&zUb�ì!x���L�}b^�º�>��[$�ڸ�0l,%��tb٬�ش�5U����k�;�՞m7!W߁F(ψ�^����륺���d��q�06++�3V��Z-T��F��hS����O���K�k��Ai�R��?��^@�yq�������LZ�7�j:EH��ꠜ��91ߕcj���_v�|3�Q�1�H�!)����rV��Az}��0$7�aó�oTb�����۟t:t�o��XMH��`(��̿@�1�*d�-z��{������1�6(Ϟ�(�[�x�ǬR�@I���7ܵ��)rc�����L�.-c�UHnB�b��壍^mC��7�D#	4}�cg͟- �`P<�q\�	�b=�f�a<Э�ڈ��4��Ǉ�B�@اo�.]@��~��D��O��H�V!K�(PrL�5���|X"�6����
�|b��S��Ke\3���Wݘ^qJ?���+!�
vs�p>.���lc��Ų��e�?��ޖyq^��fG��-��o'���S=Z�s�w��CY��Hi�r�ѓ����Y��Y̡9��d�ty�G9�_�A��J?600�Q�q���^%������L{��or�+��ϑ�*B��F�W3��+W�w��l�����%�P�7��Kǁ���l��}q^�$�/a��媕�I^r�~u��5
��!�c"��C��Z��l�i��+��H2�}9ݛ��?^W�����nr����K�.y�#ux����,?Ue>��-���
�kE,}>A]$QЕ�`O<0y���;9;��n��"J!����3P��t�$N�ʄ"�A�'5̮i1����?;lWu
V�=�ڹ?��b����V�ɫ���}�4��R�}��[���۷����c>��K��A�X�t�}�����<̺�D�0�&��9�"�Lp]�]X��ꛟ������_ó�����o��GY��jT�/���S�"�]��%ǣ��_B,�y��Z؎��Z����on�T`�:�[���b�D��)���'��ן��k��;��3B���\����u+0yq���Ɗ1�4+�D��AX=Z޴��3�21r��$Q��� )t�P���ڜ�/�َ4��XȊ�{!��!g�S�5-Ϡ��5�fC��1�:���Ojx�_�]���*���,�w��f:?
@�J�&vG�8̗Y���AYb�b�{�n���^Q@��=3���9��E+0���/�����!����C����L�/��Ӵ���n�{�_�Ot�e��A�;)_�$8�]�L�֠�'���6p�'���7�(�>��$m����^�"������N�A����2�O�?)��!��*4'I����3�G_��B��Ә�o�W/Vny��}=��~�REޖ��*�e�xr����(>�����U�s6o6O3����a���&^t�B�O�`ͱt������{m1iU�����;d�֧�kו�d���oZ��s1l�E��:�n��E�s����O����ƙ�}i�r�@]c��c���;r��O^��y��E�\yܓj��d�`�����.� ���ckH��f�ry��H�5aM���$su�$yi�[>����<��=�/M����S�S�)�9S9|�s�jືm�������c]�dc��a�&��K�BR���a��=�P��~�^��=3� ���c���/��c/��z������x�����@�_`�&�<�zqȍ�\�V�~ͥȮ����F.�;C�1*Qf�EY1٨yI@���6Q��>����"*A2��)1��تLA�!":�Lv�:�Tg!�!<b�R���O�	������C�
���C4�����D�9�
2.
L�������-�-O/5��[�m�*�:��O���>U���_���u�����Ċ�cY��Ԯ���*��<W��; m�]�5q�p%^o����h�iq{9].J+&�L�ā��F�z������>��O�X�t��������5s�rg:��y��ɣˋ��2n2\g��V]*1D�F>P:���s�|�)�'C+�ĺ��4��?<�v��)^� �~��ކ�p��F�(���D=9'�ρ���P^?�ذ�CM�m��bn(�؜nt�oe��W�7Q������I�y})n�!v;9���vsi�Xz{{z�ͽ���b��ߏ�,,#�tZx����S׾P��M����b�O/�5O��q��v�Pt�ǭɍ����qr�w&{�J����v�����6"+���"pEL��۠5�	��Io{�Vߐ�p���^�m��JE���7Ne�1�/K��ĩ��.��"��zջ����c�Ļ��܋�N=b�(16^�7�N�f���K ��t!��t�ev�ұ^��M�������9��S��'��x�E7��E*ys�I\�N�c��g�'�ma�0����A�4U���6��R��v��<�x *��ڱ| �F���j#ڠ�ίO�C�AL�%�����w�5�5���#�-H��
�����^��E��r&��%�"<�DP2��8#�$"�F�;|Qr�>�����v��»w}�T���E
JspT�z�J*�õAOqr��[DTV��	|�V��nj����D��aj�V7X�C���0�Qܔ���0M�7=���)��M����`�cء�8�XB�l��j��&���pf�7y6�O�5O��t��ix���-�(���_؆��~�+3a��[>�z@^3���x(�s��Ր���(���w�7wO
���ꝲ7�Px��;S���r�V*'n|��T�0R��dCunhKiX�b��>*�W] kh?l����ux���L聻!�<#�!ztg�6l��"q���6ƒ��I���a�I +�O�{�xL��G��g���D;_Pp�v�(��ĩ���1\ss��T�jm���3����ۼ��+������ ��Y䓢&�k��8�7�d���C5K4k ������M����dĔ��Ot��G�:~�c5�B����\���J.��܏�{����$=�5��?@�~Xk�����:�]B%� �/}[v�z'$�NǨ}Sî��EC���B��k2� p�o���oS{��
�)�QQ�U[Ps�.}��n�������jg�����!�*=c��$>t�U�(��:�Cu7����y1�jO�=7v?&��oy���s����=0��{��N�Wg�~M+�d{� �:�	���d�+8ɬ�@�ۦ�f�7�������8�}f�R
|�E�jC_c�+���o�&$j�D
�@� v������;�Uv�l�OXm��^e��Y+s�|�I#���& /Ma�*s�y큌4��t}I��d����|���O�
���8�ߜ���7��}���9e!Xz�1�AHs��Ğ8��βɉ�'a�3 ���tÜ�Ă��+6�+:aQd�*q�H,���8Ɍ4¬��7�V�f�d��.����;��|�)D�'����gWj��v�mu�	o@i)�����}�[��MIڎ�ױ���x��XՋ�� �e-�SH�t��։����hH��tʦ�q�6�*2����+��_��Զ����`� �۰�ـ�6ʾf�X��+�mD)�[��)3p�rl얏u�9��m�������o��m|�[Wm�;_f��ĕ´�N��*L:�	�[�c����1-
��z��{C&�=�l�y�eo8�e�n��q�,�s3��X��]e�&R����%q�SIᗎ�%;5�s����@/ykSf#˥�F���L��h��P�����fP��4����e@�&�^T����A�Q,��m�j��w�0�Kh�hX�8�3�)^�Lw''���]3�����O���8=Ț:k��t�_V`�r�=��P��k��@�%[�0S5rj��\�}ףr]�]�r#��#��N�N��7���F:{XO1�v\���1�r&���i���-��`8��T8��m���R][�T��"���ya<2&ig����\R �RǢ���#0,l�gU�O6�������n��w^k*P���W���L]�J�6�|��Xj�����1\����P� �
B([��g����XcU�κ2�l2r���z�=o� N�t��M��O���Z�ތ'��!�΍�Mr�������n���M�s7_��O��8_O�/$d�#�,`z+���̹�h��+.R���ho�,�%�l�k�>7V �]<��FT��_7˷�+Q�s���ZqVA��[X�S�
�����a���ڼ]]H^XhğN�C��+�%ʙ����Ue��,��ZE��.>?-��0U�{�g&�,�̋�9��e������9�7/�AY����tm���8�(��ݳz�lݼ͢����9������)�TJ�g�����hы#`+��%ڳ��ʮAF�Y�y����g-�p�뜻W��x�l���f]ő��U��qi�
���X�ñ�S+_Wd��c�bl�����r.e�������!�߿Ӭ���@���U�=jDƱQF*1�QDH��%U����
3)UQ�3)12���l�EQQE�",����UE���,QƊE����%LLTF"��cR�������%b�Z��%�UQ2�E"#Q��ƲUUƢ"���X*#Qb��UX�[T(�X�"�TTTE��#cF+X�ֈ"E���T\�%J��A`,"�R((�*�,dS-�DAH�PQ`"(
�,TX��V�P*()�TFVTTT���Fe�B���"�(�łȣiD��N��y�<o��:�>��vq ��K$1[۬�������jS] �Ѱ�B�y�����U_U}V��w�=�}�������&�R����N��T���*����<a���&0���W����E ��w�$�*A��9��"��Y�q5�7δ�y��׼����Ay5vͰ� ��)3V0�z��$+�t��*�u����!֩1�2u��4�a�
�2u�a�2T��M,D���Y��W�k�wrg;����8����+��`�R=���Rz�La�1��
A��X�=�;a�AC�P�ά���T�Xi�Nn��W���L/�ך�緣]�~w���pXi�C�Rc���x�@Qv��S�
�����!X:��R
��3i<qG��h��l��ҰR���SL=��u�y�q9��k�s��\�JͪJ�jɈ�zʞ'Gy��Ad�ՙ�>d��� �O�����3���VM��h�B�=a^�4����L�����Qw�W�����}�r"�@��T��eH=�j���U
�d��g}o�MO��H/�����:���I��c>d����:�2 *X����u��V.�t| �t��{��°��f!�ݎ��2k�aRUT����"��Xq����6ξ��
At�����=ՓL6�I���~�Tߏv��禵���~9�<N�bAza��}d�6�E�0���7l�AaP��
��>@��
ϓ�XiE�&��|�R�u�ԅg\�L9� ����<��o�s<�N�@y�1 �����r�0R�;C��n�v�@Ĭڰ��ΐY+*h�E&$3�L�vɌ=N�f�
C9�>d��;-��*�)��<? &@c����_h&0��}d�3T�gl��1�5E ��q6ʁΩ��9�T+����+�(b�J�!�����G��S��~�[�˶} ��H)du_m��]H��G0�֍�!<�X��=�l��#]�*d��j��f��Kv��|�#Z�l�H���=rv��5]RrzQ�1��odB������xz8�.H��xDύ���wg�4�P�^�4ϙ+"���J��;�,�'Y�8��>aY��V�Y�
T�J��{�@�x�,�z܏	����5���9}��s�)�Ԭ�& (���񘇩*A�N���6�a��q'��vLN�"�aS���H,1=fr�a���Av��~>�7��ϟ<��y�7&�^��d:N T�G)t�~CL=� ��Vi'N$��b)+&ky���r񓉦�!ﴘ���ڲ�@Qd�'����9��:���o��)*AN�3�>d�l�Ăɇ�d�1��)�@��gg�LN�/����W�M�M$v�_;�IΨ������#��=0<Q����5W/�\�|2<2�6���� �M��1E�I��m�2to�H=Xb��H)��Rc6�Xk�1;I^��i�H,�']kz!Xv³:�:Ov�޻�g]�s<���Y�r{CI�J���)��`m���!P���'I"�������
i�3���i �S,X���d֬Ğ!Y��[Ʈ.��{mr���"<xL�|�$N����V3�)���u�OY4���:�ɤ���(oT�����0�RԽ�
ͤ�j@�� 8��퓯r���U��A`���u݆&�*%f�w�M (�h��N"��:�0���d����Xi �׶�Y*��|�S���C�����}����sӾ��s�y&�v¸Ó7�� �������QH.�� hd�*KH�Ho,6�hbA`i��8� (���'���0��H:��z�0��`xL�����D�ě��<�ޘ�����J��݇I����0�a�
��O5H,�,��IURT*z�X-H>R���i�AC��&3L=Ldd'���9��M��{�:��	�����>ǖQ�6'L��ԭc\�%����>��W�l�N��}h�'lS��X"mTT��k�.<+ER����juy*E��)l���i�������TTuf/�x =QZ�u��� ��N�
A�1g�ã�I�+:��fN�
�_k�4e�
�̰Ă�SL����X� Vu�{��uy�m�zL�s�=��#i�N��a�X�Ă�Rz����<��oL&��g��0��n�$
�=�U&$}E�����k,ă��d�	��w�~����}�!�@�C�'�>H|����\�$�'l��'���>d:g���ox�n����a|�{�}��3�������S�v����ua�̆�q�@�T8��l����<I^���Y�ͳ=��[����c4�̤��&'*��:3ݼ�N�׿}�>}�;O�*O�� �`p9t³�Ă����1��1��1 �=���f���w@ěB��ӾXt�Xi��)�P1 ���s=y�������g'��$�3(,�%@�+X>@���j�~��1�a�����YRa�󤂐SS�ɷL
$������]�����x]�)~P<" �u�J�X��*z�J�� �Ͱ��öaR
�q���J��T��P�AN�5���
�W]y�v�$i����ߝ���Ǆ����NىP(��măi���g$>��q�C:eH)�m�7�R���l+e�P�%f�kR.�@�g���&�t������s�2N��V=�CL��:��;d��J�G�%@�z�n$�t}f�m�&0:���AgL11h��dDz�xD{��!�8g>����m+ɼ�V,�x����+9:�z���î���}� x��0�Q@��P톒����%Iߴ1��2h��!�����`0�e|���_���P2e�7�(Øs1�7������Q�Us
�p�JwT���gXjί��;t�.|kn3CMt�eA�P�Y1�/��t>X�r,�ҷ�]��n��'N��Sav�U�(�����<=]WŦ���4�Y�?��E!�����8�`�@��8�����C
YLf�%@S�d�*m���T���f����TOi��2V�~���}���s�wy'h�h19��N�
T5�`u�!Xm\k&�
y��M>�s(��*x�FO:�M$i��j�H)���qa�*)6Ϙ�n�xWg������ xD�׷�c�L;aY��&!�J�Y��� (�P����^�1 ��dֻ��_i�2o);�g��6��w��� �}��xA�3wD��b��^��Ɏa�:Ld�vbAf�v�s�E ��Xz�$�a��V,�=f�N�
J�}�x?Y:@QgYE�'��1'Z��4��E��]0�H.��g���~�w����d{cޘ�d
���u�Hr�
�HV�yOP*Af���� (�zʛdی{��A��������H,4e�c<T�ۮϝ���^uߝ��y���&�Sh��&�H>Y��rN�m�I� �ԞN�S�
��$�:2����>Mr�>2v�������d�QN�� ��`��^��޳z�fo�;��~�6,� �d�厬6�T��0��Y�εa���:��I�����a�
�P�JϹd�;Oǧ�`}jͲk7�+�z�k������?r%t|����H?�zٶJ�é�UH)�7���R��T0�>La�Ն$i��1E!�30�1 ��VL��X�i�� xD8?�t�{�>�����(��Ɉ
/<��O�@�;-"�^QC[�L6°6ְ+6�S��(�0*|�5I���ɣ�f�
æK�h��S�Iۈ
,:Ξ����w�{��C��,��1 ��fXo�$m�&3����t�Y8ʜE�T��m�La�
�����Y�5��'M�T��x�W����?�_�»rI����KG��mdef��Sћr��mY��b���s���ީek��!Փ���;G����W�Z���s&��mR�ˡ�W�5=��������-���) ~�1��N�vc+%~d�S�y���Xq��~���sVT*[�$q�C9�H)_&��xDj|6<*<�Ύy�[;�q��ؐP�J��%@QC<��O���+>d�}�9��
³L��u�Y*q�>�J�>`��6ԇA�8B��>Lg[�$�AgI��>y�ٯz;�\�~w��s�r)�����f$�.���:��q�I'R��[�b�wq��T�(�{`c0���Ri�aY2{f;`VbM] (�`T�^��uo���\��sv���p��e!Xt�c�������O@QgFY1:d��̂�{�u�i�9a���LJͪJ�wa��q�8�t{CI��w�΍W^}�=��Ͳc0�=�1 ��r�H
)Xtw�N��T�����d*v{g�4���c�Xc<d�̝�X);@�'Rvzyd�VT*O~��Fs�z��s��Y��4�@QH/Ϭ���
�Rf�6�i��4�P�7��t�PS�(��N�1IY�&�y&��;aY�O;�Z ��J���|V�ҿEu?^{�x}	$�����v����?��]��!抂hN�h3��g?Y���Å&��1of�d8�^t����E^AG�'���2�_�3z�W�Fw����H�@�40�
LC�,�V/�<�;�	��ˣ뇆����"m�J?qY�����
傱��ސk��kUd�H�k|ثs
�,����|3��j�:�9Z��-q���u��^�b;m��u}�,�fF��A��j��9�q�����;��VbY���5�ilM��S�mD��� ��*<���q�_�t^��G
z׬�1��姫_�#�����]˨���O{=�-a�Cµ�*���c�K�gcx�3�ZΙ�WpuV�Jn�u-H��Tߺ}��v��j����#�2zd�4�OZk%G�dtR���1�=띇*��r���F���Fd`��/o8��n$�|�����<�g�zd~��^ %*/"#5UB��[E�Y�L��k��G�����S���G�}�61�A���TTKB7F�D�64G�N�Yx��JR��� ���,��|V�'�+y�8����wIL�؈�Fߛ��\k��v;_(V]��MV6R2M���^�.}JZ�йT"*���dԞ��O}�7m߾Y2�����ƱQb�`P�k.�8�|�����|��aw���9��w��=��fY�����:��]Va��:bQ��'���M�s6Az��`���I��v{y�P��o����"*R�=Rۄ�e�L7���E��$�� =�*��"ڎP��T_:�HF��Q^ޯ#7��j��!L���s�59Gm+��lW�Z�&Q�W�<�Ho����4�~ڏ,�8�b>O��s�?b��6���6��[~�.�L8���KuAh>�3���f���Zx�!f]n�0,8o�-�K��]z�^�L��3r��&�=&\��_;����=�O��|_�� A�n�����wNNvx�n{��~B�)a���c�F+�x�)IE�^�H"pDM�#/o���PI���q����A�J7��d�!d�
-�s3$�қ���՚��g����Q�	��h6u�\x�-�9^R:�Gc�r"UX�u��Q/�j���s�q6��͟0�"Gj���;�F�ئ��Y�����C�F�'Kll�ZAT����_��B�O��+�kznW�]ef_��{{��|P5�%�w=n�	
�[�ٗ�VT`��\%R���X\ �\�kF̴��P2�w�o������%�=wg�dȜ�����'I2*{�b�� (bSX�X��A����L[��d�9u�`�VK�o�J�C�L@5�B�7$@5~���������T�o���/(�T����b����Y�&5��7X�?&��=��W|�IX �@��^17j�c*���΃�:/�C�k�rG=��Q'z��3u2�T��zA���F)���O�x�0Z�6Q�D����Y���O��4�:�9�^3ac� ��~�C�\!!97=�z�V�����p���mώ�1
�tc�<�5����xeR�泛j�?	��Iΰ6�� �kE,�~�;�10C�x㱄�:�f��Idx]�0jvzY_��C�$��@:b�eo�m�^�{����%〢2��He/�k���0���\��q�Aah�֍��H�e�),q�f�7}9���Bi��rV�f�����`R�e���sL��t�J��y\+���w�$,��dէo����]���W��uؽM&b���! �:" =S�}B�\�w�Tu���1G��rC����'����5fp7N&<*�e�R*�uz�有��՚^�|�L���z}~uE���g"x�~��7e�.0y��ٌ��*�O��2,T�3-��T�Z�������v�����M7o\Z3P[�NLJ���ڝɈj\�AX��56�Ey
����}ښ2yJuC��Ǧ����躱����O���W����|�g�N(��T���vn�f�~��QG�VQ�Y8x�.���i������~��i}���Wk�򜾦"���E�pč��#6���rBC�&j'�+�|X눿�����5g`��\�"��]�/�Z\�ʱG�]zU�W'����(�,'�5quGf*<��P;����ڔ�c&���`�
 �n�ő[(%�/U���n�ө�^�7d��p蹆!.nΥ��b�)�<�ӶZ&+����ր��,�o�4�a{&f�9{�+bf.{��x���Mj�Q��h��ѳڰ�y��J�x��3DcAQ/z�+<ӐeK�ՙF�����W�
�6��PsL�.}��4ss��T~���J4�>hx�(E��������_��2`(���s���AXо����ρ��O?�-�(�S�-��QBj�س8���f:&��h�@^����f�S������)�����,���	\�*��("����&�.V�LAf�5��YA���B����vd�x��~��]$/BZZ�U�H�������ѱѐ�i�d��^����9b:����c��ei�E5ay��5�'�e�pD���Q�I��^?�K,�Lm_{��Q�����/�;�E��'�i�}�۷>�A���l����>�\�͸��ʹ_Ce��T����6�rK�iwݽ1K�ۤ��k��Nt"��e�a��]V�2�\.4���"\9����T|q�[��˲�R��2JԳ��ʍ�rN;�YR�ʻ��N`i�rN�:��v�n]�W�u�wU�	���qh\���+��F�U��|mz�/7Lf:�v����'��umE����3(-�{7SO�q29��Y��)V>��٣.a'�	è����}J#i�u��I=V.�I�	|�>�~ݨ�EwY����� 0���_�I%�4��h�b�e�3�I�~�if�f�f����#ƛ�l��WkgjMl��qe*�S;#ݕ�6J�z�ŉmXjƗ�����b��'�qc���ڻ�q��6ƞ�u�����(.+�{X���<+��1G&b')u���V0�ˌV����h:��;��&��v��aۚgآK.p��?��F>�ٔ2�3q�ҳ��B��JG�J�%}L���Y&(�_ny�\o�7i��ԖK�J�Q�z�x��w�䥯�yW�s�V�5��8�d�a�nޖ^�����{�Mإ����g�1�Ls\�G{��뇥�%Ս�]9e@6�7|c ��r�"�W�'j�yS��W!�j�k��l-���Вb`U�)]'�)�e�*1��d�7�t���3e�Y�z!�捾V�S�c�EF�ѫI�r{ڶc���L�����q�dd�]P���*����lD�,��}J�}_q >���n���`�q�r�xa�@9P[|5��ɓ{��qR�F&/K|+$���.�Jru�����GVN�c��_G`�3.�]+��XFrDWL	�oe&����hǹ[Z��7اV�z�N[x�X���+nT���Gݍ]9�D�|��k���pڴ�A-�gh�ƕ��,��76W�u�A[�n����{SR�t�9��u�t�۶������,uԭ�n�X��is��՚� F"��?���RhͰbý'N�04ԇY��V��h'Rg��:�۝{ù��;HX��@R��P�U*T�KJ���H���Um*��	�����5�`ĢPej1UPQEQb�m�DUDW�X�1`��b��)X�1�AEUU��V0U�U�1��C-��m��X��6Պ�Qb�2��l+mDTQYUU���U�X��,���*��,Q)PX* ��9��1AAdR�ciT��,�ks1AF�R�h��a�*" �K�Ub�R,-TKh���fQEU�++U�*��-j�EE�4�0�1U-�U����`�j��ZV�F4mV��Z�[��(�Q�m1��*U�R�$U�V*V�ƈ,[�[��'�{����U�B�NǙ���q����x��zI�vGrq��ԥf.�l���=� O6x�b�����-q{2�����	���X��'v�y˒��!��'<��G*�:X�Gg��Pu�f�4d�t{r�t��U�c((��}$���R���4"��$`<p�^�9M��V�����z�a�o�����|f*7�Ő�j*�AqK'�bU�R�\^�ߪ*قS~���b�}�V��U>m�v�㾌Δ��d��^V�H��-���R9���嗏�1a1�X�&�{�8|1i���b�E�����lq�9t(d]��B@˦����'��*�Nm���ۥn��@��4�CԬ��a���{��������}����:�c����Q�( ��nK>�3;����{��c�}C�ڿ���M��c�`3�R��@K���������3��~�|P�3��1�&j�G��`��iz�nM��kF��C/rQڹ+��wyȾ֑Vb.�퍕�7�L;ElV(�s!֯�$�}GIl��v����M�]؟����KM`(G�d3bk`U�qAH���wˍ�1x-�!)ie*�+k����֥������^>xg��-W^=��2Z��ղͦ���r�!I�x?>3���������$��`R贇Q�V2�Of��ד�zC���+lqQ:r��l��u>�=q���E���U��6sZ�T:��T8b��q����]T33ʲTc���%{�0���n��}1瘐a��E���R���Crq����]�4��꽐�h�v�U��b����Y�'��ڷPi�����M$���Р� #>qT��*���΃�1�x�e�"�7]6���{�%�7�6��^��ϬL�܊�B�F�/d�'KT��4��Ϯ(!�1��p�"�6��kVC�y����u+�%���Ī3�ά�qR�G`ok�e=g�1c�Z;�ª��o�A�ԕ��9q`����<��}L���	�-�f3�9���iK�Z͝����c��Yቂ�Gn�0&xp�kE^߽����r��9��ϻ���#�^Fj�n|_�P�tU��ma���,��*s9"�L=�S�E�3mX�ĺ��5w�����|���vLw�)��W�~����q~2�1���.���BR7�� Z�H�ۦ1Y\Z��@<�J͂��}6a��]?��������rr3!�������4�fB�������$~��dD�ag��}VB�d/&#�}�*Un[�}>
B��o�cDQ6����| [������K�	�:��%�,!�ǉ<w���a�/�T_Rݙئfr������U�􉁆v��n��P1�Tz$�1^����z_�g��{��ޏ���4�H������CSa��Aby�rƑJ�V�HY~�9W����K��O�k��}r��2���x�[�Y�1aԽ�L���s�}|'��ڗ���+)v���N�oJ�kv�d�+家��D�|)�CBe����I:�X�-�D�^���,��}����P����$K��f� �*ЉB������/&���t�+5�ͮ5��Ni4-D��c�v4d_Z�_O����?y(�5}�K��F��3޻�q�L��忊�/n�_�ѿ����5�����1��ف�"�|ٯ �LZV����@�/���l:���$�{������Z}{j�
���b;�U����"��I��Hj��^i4.{OY��H};�[���u�S������m��zy��6~��SL����Pg|�-���0�����="/
蜢�xV����c��5�����Q����P����
 n�u�Z�')h�^��A߈o�-Xz���@Ƈ����V϶��g�������O�j^s�A�����۾���Z���t��Gh�+7�@��(n��%�oN���\+n�4&��S��{I�Q�ˡ��C����.�o\�x�]��[�M۝��捗 Q�<d�l�����m�"������>8��k��2�E�n��� ���V�U�xA���)*�u���W�w��#�x7���>>>/ʏK|r�Eg�?��8�NP��e^����E�F�p�0ѤH>Sy�'�~��TP�� ~�fF��*uy��y�� �&I�dP����'�@�=�����G�}���
��WyyR^���	�!�H�D��f�h#���	t�Z��`/c��x� �^�Taޖ6j8_�=L@�-��	�U+�162�E�Z�2x��Z�{��[!F��r���(fOH�aX��Te� �'l���~�i�G��f��>?Yg�b����!P~�"\��ʸ�6�-��)Ϟ���:�L`��d�������S;f�m��Ȗp�������i>����ȋ��*���RO.\���g��\#s|���$F�*�Y�w����^��M��~mTI��T�t'|���ںY21��gm�����/m�pmE�t��	S��̖y���Eo-���w�>�Ź��� }�糝���Q��FyY��4��x�/��lq����Ra��_XuS����o��9q���0c|dl^�GPX.\��V�@6��ۭ�|��u�5�N�t��f\Z|����O���j�6�O�ڎ�BD��n���:��M@-�G���~rM9?H}7�厽�3�R�6"=��II9��>�6%��*܎�B��:(��m��JBf�;�vo�o���7����!��r���ƈ��}��Z����zJi[�X�k>���P�z� �F����!1;W�c�U�^Ufwb�PUY�U	�S,BR�
��z���wV$����S���VV���-P�L@��յ�<`F�SS��-^�^{��氢�0�1�!� =4!�1#�>5~�[ٱ�1V\ɵ��Qj�zѻ�$e�,�l�Yͼ\�d�)Ҍ.��ٟ;��A�����}���Zv�G* q�2�P=�kv�y:�ڌ��T��+[��r!vNĘ�kO/� =�*���ڱ�@����� ����s�b����k9��#;�.'`��Q\*e�q�(H���(��~��M�{f���nPVVA8�'�u�M�ą��%�y3�C�+�7g��)��uH@�p�@Z8t��fhp��[���
�_/�c���J;��+�����lھ�u���G�W��C�>*�Aױ���6�m mV:�.�A��3UW�N�Z��0�ϜU��p$����b�L���X��4��7/7}�_j�L؍�yᜇ��.�v �*y���U̾��[�G�F�K�<��->46y���:=�m��3�$�:�s���d�R3�A�C��;��T���@������'�N�S��m�^W<e���3J[��?T����1�t2��}�����S����a��n��l���u0�����;}oaCoP����u]Xf�R��x!�ғ��]2��{j�)��r��P8�NXb�!�Ԯ;nA#�]�۪X�V8-�:"���}�xA���S�ˑ0�b��.�s�2�� ���(`��gNM���Kk!E8��!��<d]H�2����)��$���,y�kҥg{�w�@�����pW�O�8D�9b5Hjr�6�,�h�X��r���pa��m6<F��'�����Krb!�
Ɋt+��^��V�1���I������?��||_!Ey`����2�F+F��o���}������ƌ��Wk������OyFN�;����ct$t�5��'���b�^V�h*��d�/w��H��i%��^�P7U!n��$kV,�5q�\�/�� 6 �p����^H;�|d�a����t��(y��j|�/����P�^����J��	ҍs� g��0��ya�cVg!�c#D7v����Or�qLߚK�O1���w��!��Yy6(�&0����wqn�&���9r�)2�p�V�Ѳ,P��ӛ��]�
�*��+y�U%� R��K}�{��9��{�}�vg�q��Y��`hx��b-����_kǋE�,,��ra܇sd�D�>�Y���`ht����/��e�k$�n��:h����Pu����Ѧ]D�!��Ʉ��M��u���������X�>�.��\B=����̃����ێC�J�z-�i*^LH�WPؾ�kք�/���*(��t����ێ�U���|ҏP~3
M�{���8�[���s�;
U{��9�5�͎c�g{]+�k��1O��ǵ�#�#�le�r�ы��*����E��<V��qv>����H�`b5A��.-L쉣�nmf���=�����⇋��g�/fAR���<����3.�=�X�R<��3� 9~=^��9&"t�TtZ�[��� ���inz�2�e�[qۣ��;��mF��!��P4���/5䊜��DgH_(
[�WfK�sD#7oL}(ej#0���qn�ќ�����to2�NN柇� GG�j�Bݡ�|����q�NX�^�N}JZ�dT��s�ݕs
Q�:��c*:�N�̵��wK�pٸQ�q�Q� �E�q���ډB�XN���)���U^���vU����~�e�E�%�#�EO������5�a
����L-ɯ[�#rArK���	w���|�ʇ ����YF&.�������_��A�.�r*^-��v�L=�G�oo�-�N��5{ʌ�r:A�����4#gmݷ����� d?�砂��/��O��v���n����N�����3{M`�#_���:��[����_O��>T1ߨ�)I6��7���Ͼ�����cЩ���<M'�){ �Q��6�X�4��{��k�3:F�yy,��-F�$7!C����dYzG��X'd��81qڢ���w�ѣ��'rh*����p銙��xŻ����=/�/�cR�Nսs~� \�.��ʬ�Bӣ� ���
x��z��XaJ�bnpT�F5�� �7H���1��yƻU^�&N��a>u|�ۥ�J�]�1��֋�
�9꿰^ ����}�cmRCX���4�8GJA��/0�5/*�|.�uvr�t�%��i�߭���k{��{�w`�F��l�6��VV���+Ulm&8�r��u̫2��H����	1�F��l�W,�$�3'k�w�����m�p�=������Ds_<�g��R.��ѕKvMvhG�Wr9�N�޳���C���[l[Xn`���)k)-%ܞ�^���|ܣ�A�Ոݩ�Sr(jeen=�HSc��\�I=W�k�σͮ-+wӖm^!�d�f�8���K�"h�w�L�a�2a7�&�nQ�ҟ3��ig{M$��K"���
̑��qSu�rލ��� MF���	�M;Q*��3Eь��<�|V�sf D��+�[��-��R���:��be�ū�T��n�M*�&�rm�����b�����![�o��/����d2�m���^�_<�#�GZ'���t�ʉ���r�-�7�5�T5+DT�N����CT��� ^ۯWZϡ�1y)���W�n7�Mo0Nܽ&�@�Z��cYy���ʭ��j��ؒ���0Y��4E���Fصԗ7�M�c������l��i�s&ٜl�oل�`%77�p�$M[�$a���s��ՙ8Wȵ�Q	�UH���)�a�r	�a�	�`EK��b@�/\��3��w���,s�%o��T\�c�
��1�I�=E4� ���"��O\�I(:��)o5F�_ě&�j��uv�J�ۯz3}]I���F�F�V��n�u��w��=�ţ���Mm\פ�Y�w:����S��9K��4��4ej���3�3/:N�'5O�s����G$���pr�<p��$�A$*���F�bņf��%G-A�V�����Ԩ2�V�1�ecF��cj�f9S���\�Y��m�
�T�0b����m���V�*���2�r�Rѡcm�ib�m��ʂU��0��VJ��E��QYkB��J��1���`�Q���QVVZж��kR��SĹ��h��-�V��ڶQZ,H�X�Z�jT`��*�E�J�dqJ�HV�ڔimR)nZcmK-0DJV���LnZ4KX[V�,eh���ѵ\�Ķ�-�b���YE���m���PZ2�̨f&aQb�-U���f`喥ʃmQ�1�أmE�(�TP�QVڂ(�(��Z��Z�R����т�J*1��2�bF	B�h�Tm�(�
*��Pe�\��&4�������|/�WA�Z����r`�a���$8/us\ȭ��}xp'����r�*�W� =*��S�����;Y�c8��|g9�8�H�y|�>adY���p�'�w͒$^��e}���������F���42����/���j���|R��,
:��)-Г��z���5�c�b<�-ؾ��#�1���PfF?=(�u���&"G���x!Z��-��Ւ���5��ا�
g����'V�|~����s	&��xc���R"�#�1�1DU��*�u��c�[���S~�L�2���Z��{��3�=�}⟞���J�4?�ݯ���Cr(]R#�1d)�mgX�1�!��ҋ��/�CJ{P�(�f �X�Hʝ�9�vTt<�n�t�.m�V+�\��r��&|���Z�:��~����«!���I�n*I�*\��F�,a�� ��΂Z�7+�@���:�1a���
f�z����<x�����/{�㮞��{]�i�Op�d�zHQ�:°\ݲu�e2��u�f�.q������V�G��!��̽ѕ�n�<��~�?x}&�O��[��3��5��w�,�/�޷�ֈ����;V��2�C�@̠do�+4�x�����/���O���p�n�$>d��QN�rm�Cr3�A����H�*}�dD�a�{�2�Z���l�|�Q����q��U*�Rܸ��O}���X��e�W��kg����:B5dg�A�c�_y/ya��>7��{`�&�%	A;��W�.:)��Q^���LS)P>uLE�!����՛�]���V��>��0*�Y�7��������S(��5|}��KRl���z�yz.������O�^�g�&%u��ެ���Gډ���b@4?�'hD���A��%'���u����[��%M���!�D�����а�ƌ�
���%5O/��� �5(�=�F�X��/�m����IsJ�Z\�+{�\��������Xi���F���7�|����C�N��9�s��3ҭ+�7B��w�\*�DX��Ѐ���]��S� �������w�~�\�|N��RtLab�&g/����|E��eq��xgh�q\����?n߶�PP7M!#�Ѱ5�Қ�lBUq�5	��EQӇIP�r�K�欻�0� *��
VwP���+�YB�O&�<|�S>�چX���M��P�\���)x�����çN&3������z�b���C��в$Q�m��3A���-����L�;yu��w��~�S���ƚ���4?����o��T����M]�m�5����R�t߱PRޑ���j趂G
cC�������Z���[Zz=~�u���ۑ��]�W'ˈG����O��Y�J�9]��L�<������������|�q�
������EM�u�����#J�o��-?0|t����)TVz3�N�b����'2�\���z$N�h�/Y���wna�yNg)��i��E�)-\jc��v�����;��R��[�}�|��S۰}�y��;�$7�+r�Q��٪�΃�R�댾ݗGs�x{�ԡ�i�66I���A��M y1�a�> Q[����6�ӛ��j,����V���>��������"�ڠ����.�b��9���#5�X�LAb�(�$(5�2f�ng���,�|JY~�/,	f���B <�?�yN��H�:k͐s�~���QJqF�Uq�hdZU��
͹czD'>�)jm2��M-�%�\"����(�� �S�F�1v�~��0�ᣛ�Ry�0jx����\�=��<�������1�j�㷏�cޭl�1�q����d��׶�1��J?Wpnv�^Mzܡg\�X
���Kh@��\�~Xp�0�W�4�@��g�+aǹJވ���R5�β�N���[����<p��,ˡ�_P�t��hwk��{*��������y"�m���tKY�uz�:��;m�Z>�:�]�|����5��'noyV2	,r4��3:eF{6n�"݁3}���=�;�'.���[��}+k8�����$�����%�8�{����G���O���;T�Y�~��������������i}f��g¨u�=B���{V��H};[����۸])g/��������}��
�$o�X�a�t��q��Zz���̼(r	��dX�P[t�m�A���zfߡWE�p����t��}��`��?b&��	�8thCq 4W/���)������DH�R���:|��s~�����42�ӗ��{���[�*�Sp!�X8�\���	�b p�5!�c�Ղp���K����`�Q�b�>(�.1^]�,�=�.�g�W�&`��dv.m����c�g��O7�^���j&��R>����U�{|:�w��(p���µDv�qD���c.U�G��o��:5�Ѣ����5��c#wa�C������z�K���rU���ɻ��>MT�[���tb��A9�i�Z�bi.&�spP����[!zy����쬊�14Aɛ�"'�gv}s8����e�T$`i���/����jρ����_B�)�@X޼��Qr*z��ʍ�8�j��?��W�fٔt1FJs`l�^�Uq�ʎ;^�.2E�S�#���9�6�$��U��(1q��u�A2�Iΰ6��03�I�N3��w��i}4z}
�"���<��;KN����9�1*Ӫ����}��;�����hT��!B�������\��6x!�c�[�>m��C��҃Vr�i�
������X���kӵ>��p;�w�>Lb@�3�{�������Q1��k�WS�x��`�^1.FT���X��e��Pj�(�P��V��+��>��Nυ?�� ����A�]z�Y�Ȥ�]nɳ}�6�l����L��T]FR!����(��M�%�~'�j����x!��	�5M�Mn��xgL}·4=IL��.�M�פ�#��bp;���wQ����k�~�TR���Pc��[�@�8yJ,�ۛ1	M��eL�[�܋�����&����M�nNW�98��XQl�N�t#d�Y��g�[QWI��J�\E���B������k���z*�fgE�F�mnkk�Z��^����NWB=pv0�ݼ�-�����/rVc@�N�εFT��M%y���6�U!9;Ջ2�g�&�|����8��� �'Ykg1��L^&�r��;띡os��8��:�G>˓��5��5�~EEQ��"�R��/�Դ��P�a��@��p�ȩّ�t�
�hIF���Shz���*=2���6�Hc�A��!Et�kl)���z�cD��q;��1g���ٶiy��.��[����R�!I�����e�MH��<�ޫr_�A6�'��������NŎ�²�uԲ�2t�rtr;O]�g϶<�D�+}] ^da>E�S�z�F8�H�.^J�b���Ė��IJ�����WE`��k�3�Ӭ�G@x�b۱X��T×ǻ-s�/
�M��b��`RA��
Y�j�Gmp�즫E�|�B{uL�&)%F��{9�$)�E�^J���&�uvd��%��`�B=�Q���\��Rk1���(�F�n�P!�1%�@��*�l�J����H��δ�j��Nj�.�Tv��cLrsA5ڳ�"�����j*c� �fZ�ruJ~���}�d����@�)�%߆P�xR�x�.�ud�y퇮���9��;�Wά ��4�<��!��*��7*K-9����lv�4c=Ӟ�79#�Lr�db߅P~��إ����(�Ö�NҺʶ������C�ք�ZV�]����(F֠�7~�5��z� �8Ԯ��=BK��7t���r��=�+���}�Ղ�9ey����=���c?p�º"�go�	���hj��[�56�ա;���F��ڻ����9��ug���)3m00��{�Y/>{X���2`��ý�0�w���H^2F	�u�N��XL,Uթ�ۖ�P��-��]�+m�?A���\^;sm
Z��=���o�{~�=o���رIR
H��x����)�j��B�Z�_T7�X��zJ� �JOf����C�ԝΡ�(�w����~w��
��[YC���#�rɬy�hK����y�.x-	���!��D;�w����ĉ=v,��ռK�^��G˴�[���|N&��bO�#%�zB�N3�5����¦�+����Tq��:�~��4�eM�ھ�x9��*�g�m(�|Z���i:�������B�*��Cm�����|�\��{��l�Ւ��v=�fM���lڑ�:�,���um܍�$�n(bU�Iݻ�B�t�+2��kIkU�h�0�=�i��S�cϺ����ݹ�wSIF%�S���ش�j6R��[]�.���b ���xNUu�֯'�v�4�����{Oj��o7�7e������2Dm���e�;��wa��T�p�����KN��p�X�dG/S��=�$�j���߿ D>�K|����]b�v#��Ob�4��
IFp-)�����+�r�錢�p�9�R�*�颞A���n��+�N�^ݵr�Z�O-�u���l���M@�׷c	M��-D.P�D`�3Iߛ��x�Z1
u��s!č��d݉Uf�$����H�@�����지��R���wfgF��]Ia��]J7�Љ�q]j͕K�T���NW�z��FU�U*�@F�����K��14u��<0>Wם�B��Q��4;�)A@�wT*�PX/Kr�Fm�ɰ8%0�z�c=K��-�v0�B�r@�$�$^룗�n�ά������͕�P}���oi3ε���0^N��ܙ���GbKU�F���V�8h�6���s3�����f�"��[��9��|5q61�i.[,�<�`�y}hҾ;�4�$V��'��̈������|%L�Cᤒ�/�p�:]2nw������9V/MY���eùť&��[�/�E��/i�X'*�}����W:���:�`+ã�t�ELGxN��B��"����+�D�ʌgr�o�_f�1)󶭭��Űmm�}\KW9�	쿍�R����sV.s����aF��WFi^JܲV���R�8�ʟGg�f�	�r��c $B����|��07�JQ��W�r�ĲR��)��%��`G��K~��垷�.��d�+�$��l̇tKn6ؚv��+D�8���P�Au�u3%I�$����<�R�[[31J�ʚ�J'�84nf[ƺ�F�$���N����b5W�,�U2���o�a�Uo���:�{�!5���Ӌ��ʸb�\�]Hr�s��Q�l���:��GD5*XQbLל^F�K2�{('ݍd�K����}X�օCL�_�Ӱ��s���t�sh��Je4�Z��^c��9fP�sN��]�ఢ��s��,ssR�4&�r͂�����[|UG]�5�*�ʎ��M��M}��9	]�p����"�Lۇ{���V�"Ԡ�)bZ�P��+AQdQ�S�"����)H�Ũ����X)l�jڊ��-�
�UKs
,TL����Z�m��0W)cD���-���J,eUh�
��)b��DL�r��X�Te�b��V��T�AKhԭiZ�"�mT�����1QX֢��2�j�V�(���1J�mik-��Q�[
"+-�QE�,V���(#F�3��"�����S+b�miU*�PU�(�F1F�,QUX*�/XVe��W�b&-�U)mLh��1���0���\eiV
-J*�X�ֵ��V�����j�h�p���(�WV����G�b�ʔ������4� �#�&0D��$UcEL���1,AAb�?�����O��gl�o�ɸ�t�v�wmA�[��]�	kz��bf,��ȃy�����V���mcT��I(1�)h�Bu<WX̪k�֦t������^��1R�i6㟔���4d]��փYY�kRj�s#r�ч�������%���5��ь�\���T��AX"�YW8�JT厣z����@�������
}�jB���^���>��6�Hg�5���i8Cbɗ>��p7J�j�f(��^�%zK�Y2j�>���UדQ�6�$�=�t�RY�T�ikt]]w�I�:MXU����c�4,�';KJ�{�|�C-�~�����b6���O��:t��Oi�':���/7Z��ָʔ���y�
n��2�c�]��v.ħk�1���iCCO�d`c9�i��5Ѝ�[͇�i�F�u<�Ԋ�[��iց1^������M��#ݍ��4qS��m�(��Q7��A�]AosMD��+V�^����������Fi6u��U:�sHB,u�4qDM�JZ*M\�[��_�>X��6�^�|W֋�엙���Q��;(	�*u+��NV�Jˇݼ[�)��b-���}�j�:h��hIW�wp�s-3��*r�������tCX���{�c��3�DF�4�F�{�,k�{�nj{��}�ݱ��2�dpoa�I��y^����plWT�V��vl�|G8&E������_��ڊ^��;,�B/���:7<S���}4���'m6.���@L�4��2�(!]��*�]�gW.�d6	=&X"6s�Br��Fn��HN�Pw^�L��^^=$�W�{��uM�KF�簻g5
�/9�A�2�n���O��hc1	zx�S/��#�l�̇Y|RA�U�hej��f^�R������E����z��QmX��:ۥcD�`��� �yD �w�o4Z���,Φ"��D�w4�w҅��������k㸛G�k'�&��[j�i�64���s#e�LD�Д,�=�����'��fY�r.�X�{z��S����UT.b]��L%F�����D�+�����+��*N��|[D��teo�(�#�С��Ԥ���Yӽ���wJ~��t£y\��M�֥��/G�%�yy���Z��2,��p��uvq��dT��Kt�jp-r���<���Hn�QןD���9	�o�Oy��}&)����l׿�T2��~Ț�>7X��~r�k4|Aۊ���JL봪+u�[�;Br<�eX2�n@	�d5�GR.�K�\aa�:\T,���2����]��D�Gv���=?��m~_?�W����(܈������%SŪ6����R���W�ak�m��3�OT�DY�nū�I7�X�������r�6$���5�G��4�'}T#���c+}U-ҖZ$��cDM����y���	 �mWV\�9��γv$:�C8�Fj���&�X���&��j�	d=j�� E���gSA}�n�U^!v�V�m�U`e=a!��A�!��z�����J4z��EW��sԦ�gX�\S���Rq6�q>�(�3�>��~nǞY�����v&.�T��Qm*���r�X{K�s�1��SAnM�Fy�v;eҙ�aj�<���g�Y��d��"�9'55�a�P ��O���.�yi'pn��[�I�7'pa�KV�V�fK��A,7Z:�+�fY��&�m���s��W��}3ץ$�%^}�ڷ�e��'Y�َ�g�wڑ75*����f�JR���g伞���ל���{��^�by�s�¡�D����'dS�e�+j�t9�;��O*y��{��z9Д�	3O�l��1!�-M(�~�ԷFr[Xy%�LPA!��&�ʜ6�+�W\�y%�϶j[�f�[]��R�iXm��u���^�v�)�Tĭ��}�8�Sֹ�}���9Z���9y�6��@�cz�;%U@"�YW8�R�.�[��|�˸]� �?r(_�� �a�HR�X�ɠ���*�bK{�fe9,ZiƄ#�ˑ�$
�4=��"�Y�fA�,�,'�gN��|b�����cid�Ф4%��r�
�[s�<�Xp]<b�YR��S�v�5�ծ��E+5l_d��"�xd��Ʈ$�յ�n�S�~�� @'1�^m�ς�9�Q��g�j*���ѣ�'���Ōfѫ�.�J�Q<��EW�U��[�ژX����{(V[c���c\rZ0Ь�9ڋU����̻�vV\�Ƃ� oZzZ�>�%����|�'jƊq��VU[ڶFߵH�%��i���<�~��e�8����v�X�'_˭Or�c%��8��^gTP�@�ʙ"�Iz�
ΥIn��~]���E��r)�y�N�"��2$&��ކJ��z�x։�v�k݋>p�a_�b^}�AJ�ΦQ�lʞ��гQ݂�3��������(�<���#�y�9y��f��K���i�f
Ңm��������V96���WGa��,.��q��rs�Y]Q��p D�#�J^�pe�#�c�2���bMK����Go6���ȗ� �T��\\���2T�mûQ�X�]��^IB��Ω��F�����ӕ�ȴ�es�aRͦŊBA}�$@R��g�"��U٭�%�F��]0Ɇ�$��#vs��,;s�g"�B0��^�l�s+!�o�q'����$�S4��(�74�wҁ9�-��ٛ��Z��j0Ȫc�qDۻ�MU�=�����KsJ�������Ѕ,^�s�8+��2�]������^�Aj1�M��wr�Pg��W[;J�YVߡ��;1�5�u�'�Ҭ���F�.��1�ܸ��".�O�dج�Lm�K����J�&9�Ű��}�Z+�抓:b��1���4t�KiTW��Nb2�wkV8^e�\e@s���흁l3�#��g=�9,����=R9�c9s��^����RXo<�<1@��oB6bv�]���T�P8���c�z�wʵ�}�-sE�z�Q��C�vu����+�7Ԭa��δ��#���w_N:�XΕ/���W,d���!wg|ʢ~�p��,R%x���ս�xЅT�ޔқ�`W:mvmcK�m�?@#:���uw-��Yk%��������u��N�c�*A1[��O.]�Z4���T9Bɱ������1�#m�WE�d��5��!�"&�8,$�s/P��.E(����fud�Q"��m_	q*��4�{��q�B�[�=HK�`�#(�Z��Y9��c//n�c���n�#�6�H�V��kt���Th�(d�W���"T7�j�_@n�NH��&���Z-Vmi���d�d�um=�Fj{>�-Q�p���E�TJ�:ULv�C1����8/�����3*b횲��ԗ���d땆.�\�4���_�*��[0�Ї�4��BLK��������}&p�3��������R�T��y�mU��hV'Y��0:���;d��횽d��/ܶ(<C���C���g���x6u`�.�Dj���u�Mk�+�F�L�^��Oi�a��.��q{���W���R��/��В�n�t�J���)�'�6W�I�9�<���� ��hv^�ce�-m�I0'���A�%�]��*V�ی4�f��{�U�놐���BB�Ez�7�^S��.�9�u!�r��'\���4�s���~�k����[�5h	�����9������W��6V�k����m�6f+F�Mw�@8�jIbo�2vA��mv�ӖN�������4��*1�_M`c� ���u��C�,Օv+����(�Ń�<ؔ<a�$)jk�7���9�0iu�����%*��k|ӄ,t�s�+���y�Z�QOj+��VWPf�x/S5p:��M zt�xt��+�f�y��,ӫ�n�҅x�Q�h#�D�u�&�)Xg��6��M� }�ؾ���#Ӻ�n���L�.$0�2�ӆ���/4kCS4��3n��E�3��hRcg��,O�۽�r��෴-����U#�U���ax�ՃO���@������śL*�_�_a��n�-�sF���!\H���_-7{Ch78�� :ڻ=�9�wGj�\��Vt@�)���'(3��
�FF�{�[�WU����q�}o����\ z�=�d�i���^)���c�)5Ҁ�b^b#+922�υ㩙�hjմ'�2��Ͳ4K�ik����Vk��f�^��Mv܆
�I�j/����{}�F-�*�v��*&�V���4fEe͐,ǹm��Ԛ4�V�ڝz�"S-8i�p�Ȟդ&_S}Dn��L��*�w�txr�ׇ:���Y��1���2���N��n}/e�������r ��p���ۦ�����3��2�[��6Lu{xH�*.��.�0n�ק/����t�!�Z:���A
vWƴ���u�.��Z��������0TB�*y�=6�)A�.�b�׼�V��[�FJ`��)U��k
k�v&�REI�Ʒi�4�J"�� �����z�\ҫ����0g��aK.y/&j��uc^�.��әeH�3�BT�����Ei�-_�dv�R���9Ћ��g��*Km[@M�x�=n<��"�kΌ��K�D>}C8���4���w{����I�ԟ�u�:��Ah�}�HIV��2�٭��x9X�(:���=�v~�Ո�C���O-�W��4�R�7�ʚ�kZ�oT��1M�y�����R��lYՌ�w�g�tr�v�����2K͝��j�f���r;�Y6�ӬXU��d�E��ʙD��_ٮw�����|b6��ghB�֮�B���v~Amn��.��Y��Ӭ_9l���h�:�Y�u��]{l+�Ν�~�ܲ.�+o��4��ىc�]�L�Psz;�uջ�ؾ*��	5^]�Z�G&�K����)�����l{���W��i w/
[s]��@)�n����U�X�$`�l�U��.�!u ��D��ŀ)��M�?-���v����W\D�pI��*B�9r�n�Ŧ͝z�)a�-r�i޾����^�}�"��2�V�E��UQUPQX��hUEYl+l�`�`��1��Ur�Յb���\J�*�T��PPW)F9h����T���*�DDDƑQEX��j�PTQVQe�V"�[`���h�mkEQX���4eQֱ�)Z��U�J��Z�V��֢-�b�Ҋ�lX��V$s2��ĕZ��""�T���.8�1�Ո�U�9�X�m�T*��ST������b�EQZ�EQ����C(�"cKj�#�h��""��ʉEU&���ʩ��b�D���H�+DAb
(�.Z�
(�9K�H��$Z�W-������EEb(�X�Q�)[`��ʪ�h �,b#��h��0G�#��1X�(ֈ�p^��z�����36E�*'M͘aؾ����vdg���o��$c�:���Ȳ�W!Ѷ�Z��ފsB�y�ު�r_:Y��w�Q�伣�9�
���CQ���$����t׼�3�o^�9D��W
��}BѬ�|�8����;Ѩi+�1Ws�
���g§��R�v�#��qeko����4V9�NvIpg��eauם��[����t��ua/!(^��:��U����D�X�w2훺�^���:�ؔ<8d�U��]�ʙ�-6�1y��ڼR��>@Cb�U%E�Y�����fR�m��bN��������4������zQ���Z.�}J�j�]�b���T��F=��2�����)֊� c�f7��ji�Z2j�s9��^#����q�G:+;齓m#�``�R��i�1ՙ,�,O�L2�J�A�qjv��鵛,���ؓ�^��?xe*��]�����Oi��̶�C���(1]�h٦�*��2=���74�:c�O�Ц�Xyy^w���"��*��jwFB7L�{�-T�xfv�g����Q80��tBu�8�{s�~��!~+�J�p����F����s\��9W�$�a١
��Z��H�B�}�5�~�sB������7gHT;_����*vim2�gH���DL���"�"ı[�۪z(���-����?oWB���wR�߷�T��ȶ�+�y%�H�2������n
�/��V�h�5�Qt^�`���J�l�}���[+�W��3��1[���TV�9����h��Ƅ� �ͪ�7�R`&;`��ӯ�!��KF��q�5.F;�.���\`-Pp��u&N�ÍѺ;+��B�qz��b�܅�P�������s���iU�<�=bv�i�m�a�wt���l߱Sע[P�>�����N��Y��V�$ �;$p&�pUB�Jܶ�)��8���F�e����7�z�r�h2)�]��|�	49��B4�P�dv��M99��f�d:�Ry�T�oE��9,<$�Up��e��̈́"�h�RN��s��c�g�8Ҧ�D������W�kU�i*��q��ګ���,�i��<�'����ID��ձC�YV�E�+��N�;P��"m�U����e:ҨafP���Y��._2mj�����z>C�3�h=�B0��]�m9(^ፀ6Tݻ�������GI+V0J	��7�Xy2�ѱ����
�iL���r2��;��7���1�`��JÙv�&ғo,��	�rb���T�>�\���|�P$.}=q�y�fVk�K�f֓v�Ex��۔�3A�S�=�ڵ�mi~�ʷ \�<󎽺#`�A��"g���kF�ͷ��]`Sg3Q����Jch�Y}�n��`g�@y��&�W�:q�u��J�o�Q�u �Y�T��:2٪�;4�uU�]��>l��QڣYM��'��K2)�M�#9�m�o����,�� �*0��땇�uTV�L�a��7+#�s��B8�uQNpC�u4g���dۙ�m�	G�W]�����T9u�h�����f�Ql�e��d��j��+�+�D�����o����|�I��Ε5��E�r�m�W=H�>X��c�K���aod��f��ʚw[{8�[��]C�4�^mX�u�Ŏ��ʃd�@D���&l�OX�kt���ɺ=����U��0VwXw������93A��f�T')NM9d[�8u�D���;�O9�)�KYre!�b�@���kIS�Ғo�Ӡ���޾E%��NvU�L����R{������4�Κj��Rkq.�;v����3������s'Y7
�,2��r���Q�<u�{�r��mqy3�R?a�Ϸ��ӥ�YHm��[N�q�[�S跳�}*�s�N����p�p�iE/@�G�qza5���y�������YW+z+��z^Prv �|2+7:���+��M�|}��ޮ�L�m�sc�.��1�zq/9պ�-��a�dgrUri���cFf+�䯗�_{3�����k�ӫM��A�|��=�N��I�����O���1R��e�l$���������4��2�����rFٌ�B�Utz"]�l���-��~��Y�[^��1"��ml>��*�g9��B�z��%S��fM�t{Cg�>��o����>�,��у�ݳ��ծ+o]�;�OJ���ygj�:&�����C��s�����=�}��r�v
��|�"��cW�;F�}h�(�J7�
���=X��=ͺy	�����rm3�Z39BX۩�v'Q����}�<�02����s޼5+uA��
�u��Jl���fWV��vB:�I�_k.�:��HZ_L"fO��\yV�c+9�ܫr�q����>��ԛ0��N�F��UۥNQ��;�{W"�1��p6��3Da��Yy�/*c���|�JWS�6B�K�;� `��3"�:�J7rG7[_��w���'GQ)H@�$A�u!X����)�י �v)�ofZI\qO���vUAWX�-Z�8�̈m:6�$:�9{m�x�w
MA,!�m�H*���)׮��O@�����g��A5nuH*��ংKf۩�	���.�̪����4���~�:�k-��'�`ڼ|ʋ�c��bJ��k���>���Ʃ�b�N�ZՌfѫGZ�9*<$�U��S"v�Z���۔@
Su�L�0��+���q��Y�R$�v�oJ;���5B��XJv��Z��<�f�;y�3��ʻ��:E�+[����]s��qP�X���(��Xz���_s�1D��V�2�ޕ'��Fꍣ�w�iu�2C̸�ET+�C���鮁��R�&V�d����R#�ʠ-�["�^1c_%b�����~�Y�y��;)֕Cξ���4&�q�!��u�����g��#o=2EN�$�5�]�E����x�:�����5��������ҁ.���ߠ��CA�rה��݆��ڌV7�^�Jqf2��hk��J>g5.�Wj겶s�5Я��	~2s����t��4���1˃�}��X�]䰒�8g\�3b�F'#�!g3��q��3fN�Q=P��Y�U�}�o��d��:�ݻ$�G���yV<�a����k��\���@ʽP��)�2��x���Qh�qƺ7�� �d��p���\@PY������{��Df���M��! �>��g�\�_,K������V֜N(�u�V�b9f�_\v�[��}W��e;:�R�C<�s��l��	˜}ǧ)�|�6p�x� �i��4�\��V�<�R���E���S�Bh�̫M^��lomC*�rS\��QlB��]A��{�.z��OoY*5������ꍚb)6��^����[K��D��X�]@�r3J�R�+���| ��j�q�/����IY��as��E!K{�����}n�g)W����I��\v�L�}c:FI������>��]�%��T���tH����gU����	�In��ë�p��mQj�V�:�U����.���M"Fv.�)wJ�(��3{_B��ƱP��<���PT�jʩ������!�#o��K�#\�2+ν��Z�^�Bǻ�?����b�+����7����Q��u��ժ�� ��紤k��G�f��.:ڔ�Xj�4��NLBzkyT E0�V�..n��6�}ٵ�i^VqA�΃�P��[�g��H��a�8-��]aӡi�t� ��+�aS�I}!z�K�(Y8�p}T%�
X���ة�S��9im)7���ԇ ���W�`m��}wcM�v�[h����(��Ee�ھ�PvgH9s�Y}��TD��CZ]P!Ob����P�J��K$�]Cvm��eV�A������{��R����l�U�g�GpVv�b��3/��:���n9��5��A0;A�ne���hozIu֏p�ɉ�V��0�x���/��#C��Ol��n%e!/�����&�,u[�5Y�v�<y�H�<K�T=0�j�|�~-�Z����nE�ؤWYu��v$ș�LBt�Z�����NQ�z��K&B���X�^nQ�<�]Y�n7��<E�)^J��x�b�7��w$u՝r. \��2�KHJ���]��h=u�k ��LQ�dv
�w�	��jط��"��s�p�zz�xs�첌")�X�c;Mdګ�
]M;�6��!,k�;�d�¹���p���. ˖a0-JO�K=Y��m�eٽË�+�y[Q�Sq��VY3uWc�3���[��U��Nf�TEn�׌5n���)վ�)��k-G1�չ j�5�A$�[\�PA>wM�����l����+u�ݽ��G^%uʊ���5���w)Z��s�U�Lz`���M^s�W��㙱L�(T��PÛI��	��pK'���xwg�q+��\}�0"�n���7
�E<��-���T��E^�}�'I���^k��)ƍ��r����k����Q!�/Dܝ�3jZ
�^�饽�Ay,�Ɩ�r��	-������|83|A�zwVV��js;��m�84�ss2��KN.�Z���[ŵv_w�ЖՕ�[� =W��ώ�A��/������e�=2�H�4�K@����Hdi�a�HX��
Y�}iC�� �;�����t����bR��"�>��#X,*�LϷC��6��z\]u��t=��	�Nn΋dy�E<���YG���	L�;Z���s�Uy%rg+A�l�EuH
W+�b�>W�բ&�t;㧶�ʷ�f�p�I�dy(�/�];n�Xn�1�^zw`���;��j(/j�-��>[l�L���r����49�z����i�N*�]n�Ot�6��w.W
�qL��sY2��Ҳ�7�a/������N��L-{c�C�٢���u+1H���){�*��'n�R�^�X�E�S6E�0͜�n<�;��\�c���ȋf?��7WWUuut��b#�;��$�J�F*��jTVDX��V�EJ�*[j,AUEQX���QJ�X�����eh�X�QQm
(�1��UAUQ"�������d*(��*"�j��*
֌ER���(#k(�Z �ڊ"��֤PTj*��Kb�",����KJZQD`����F(�����TE1*,�R�VVPb�mV$����Z֔jKKETU*��c��1Xy�n���[�4�z�
�Z�|� ��(ɱ���B"��76�\�[�i�۝�����1��8J�7�W8v<��NT�և�n�6֮mD$���p��>�U�W��4���iL-���:�D�!����]�O���ĹgLb������a�[9J��7잯[��\�*��,�J�z���愅`���6vi�,Қ��КU��mE���N>%�(����$2.��[Uϗ=Ii���H�bT�Ib��CA��x]�j:1c�I!��Ox����ܵ�����hg�&=K����|���|�&���ֻC��\AA��&1jK��oi��4'e��H��:�V�:�T��h�ֽj�'b|���,���Z%��e�۠z��5l8����P9��^�P̮oC;��<mI�a;�Ղe���\=s2YV��\�Y�Go�qY��Ri�սg�����>�mr�m��B��<:w:��)H�Dd����$kh�Os�P�zTӄ,tᇜ��m��]��k:������5��".���V��@����//�mQLf���|sO��Ju�-H��jκ����ˋV�l�fU���(VZzT����׉4�fv����-�y�С���,%24wj�Ф���Ei�Q�����Fn�U��M�Aά)+XX�q����֗C/G���tˠ�T�K��;ݬu�+W`i���Ȅޙ��kO�j�]c;:^�{�8�k�nT�U�}.�;���Q��ɲ>�z�=ib�����]
�,���u�Q����*�(��貰���J�u�\��<Fr,]��LXu�c� )�oK�E0��tgbt;NHB�Z���h��u|�8���F)ĕ�JG4[F*��4*�2��wL����#�WVq�w��h.���s9�^I�8�Ԭi�v�j�])=]C	v2P�ҥ��BrC5P�u.]���1o"����b�Է���lJ8� @C���cM�2ڵW�1�إ��U	f��I*J�*�ve��v��gQ��16Ny:V�n���B�洓�*Tv�͚8A~����#6�m�zP�F�X�;�믥՗��|��pr7N1�O�;�����{��&�tn�׮�;����Fn+�P-�b3���|Х3M�rua�*yq���� ŗ9�چ^��G�lˣS��r���W�m�[y�sZ�ճf�K4��s��q���R�Q��^�Vt�g]t�D�'ڭCHDu�z5`��úN�He��T�(X`�G���T���nf<�b{�Mj���t��lJ�ң��
�ʀ��8s�A�/Q/�Nwv�Yù�!�Z8�O�#Wy�����,�[<!�â�w�\h���{ͽ��,r;rFm	dP��\Ҹ��ܻ�Yϋ9|ۢc���6���T}���^��`3�'�'u����_�-��H^3�`��[Q"�aڭ��Zz��mrͼ�M��ۊ�gh�(f�ROi-U�������jGZ�/m6.��#u	���GN�i+	�������ϧ�����/}���ܫ��ȝ<@|^t]I�:U7�_0��m�ZD +�z�*���(m�t���%gt�_i��\��xk]M����訴n�:�,��Gk���Q�*SA��lS����G�f�g�ԹS�~
����VC��۳2�6�Fb��`�b0In�(��֨�Q7S���3+C�ު�o^�j��`�-&�[��ֺj�<FBuy(o_��ݛ��<ڪ~�U����AF�TQ����o���2x�K۽�#\%��p7k�,�N�i�c��Ҡi�;�Ϋj�X��#�˪�7]Fn\󨻒)�6��)��+V�H��z���U�+��I�������-�(7���6Y{ZiP�4����g���}�r{�0���\���
���=�	
�X+����}�2���NG���k�c��t�e����$���5C�����b,u�o���W��pT/��U�d&X'@�����؊va#����N�1d�Pm�A��M-q�r�L�̰v=M2�L�k��l#'����/{���ݶ��t��[����.��Z�Tj���XbP��P�)�khvR�Nr����Z|ڍ0ד��&�f7�:u�8�-k���|���av�d�MW�Di���U^�9"ڼN��+[��ngt���Q��𢐩"G�nuH2�V��X�y�ڑV�v���f��@&�q��7�l��0%��7sOE5wu�I~�*�9�0j��y���541���SɈ��M�u�)�(Q5G$z#6�W88Y�<�$���hC�G+{3+���B��T���;E����������*-�/1�u=���I�b�ѽ���ܣٱ��Nl�{;�<%�ƣ�����ئ�Mg�]�t� Eߕ��S%�r�PeV=��wpƺ�K\�Ⱥ���)���rT�Ǥ����I-ʖFm^�Q�����dlOg�����^�}�w��|�4��N��g)��<��/T���)�R���J���@�]�8x;P��̩%:5�Q{�L��窰�f���\'#I�g�j���:u��<Ұ�����R�Md��8���o1�A��많��/y����]H�<��m-&>�/I�;��ѷ��Xj�p�9�^	2+�O�(���[e���]�ܯ_�7y(PiR�pδk�4H�U-Mͥ|��r��Z�w���N�6%1ג7��VA�Q[�Qj�b���#)��>��j�IQ~a�{1�]X����t��=K+���ٸټu�X(m^k�_-m.�J9�fa�wA�k=�
�yj�������uf!�9P��u���)�F�H�E��Ɔ�&�۹�aH�wў|�v�y�0ed�iXҽَ`�	���u�����+5��Vo�3�j�55n汷c�
@��WL�5�?�A�"��;J��g�p�ӓ��W�MJ��a%��!��њM#1��x)�fY�Sv��ٺq!ųV[J��bm���v���i1��Іm0E�p���7�e�W��K�{���`�_J<��zSd�6��b��/ݴG��V�介�O�~�qH�G�x6��M�_JY|"	��qKm�����1���׻]���큛���}M*��'v�V�P�X�N�y��Z�rx�#��o���"����� ��px�壥t�~���F�S:��6�C��wy��p=[�Dr����u��Ssy�ul�w"I+���r璕>}�ns[E�����ES��vm���[��}���\kW���)��	X=��vf.l����n��i��-n�n$�&�p~��<j�ia<�6�J�f}�MV-���u��N�bsH ��)��Ũ%����
��R�1R��R٩��|c5$���*�pv�mh!��>ʸ�����E6єŐ��#��ʢ���������`Fv-M��،#�h5�����e�~���3�jnN���,�ig�Ҳ�])b�e�e�&�o�;t��kiL%�V���E^�2��Ҥ��n#�p�Q�U�m�{$,s�w8�ʸB�֩�y�#|�T�|P����Q��^�����41���"�]�w�#FY�#����W!�9,�:է�>��=<��Gi]v
�,
��pn���<.��%앉Y���"T�y�̚�-��[9���$'j�T��jvi�4'C5������-־lE�6t�P���}�y��V����O�Y�)�jө�`���&H����uv=�W~�ׯFW�|��-�F��l�<�*�mI��C�k)W�;X��Xy%�I�Zz�qw�дq�R���H����^�H�M{थo"���?)ZjQ�����z�h���"�"�NO+�J�RF��jlC�E�;7�''&���P��\��T1�!RG�΀R7W��,��Z����`ʡc��.��l&�p��ӆ<2�-�G>��蕖#S��}��Vzo�ӓd>�s=& �F���F��8䙡�V��૞V�>���3k14�-��,��1�}$l�t��+r���&nWHdzL��#6m�j��XF-�`U�8	e�el��GdWV9<���C��6�W����%�eBV��&C���<��f*�\l���`کw�pҼ�v�\J�_&��v���xuk��֨�#w�qv1Ր[S�QH]p�95Mޗ�d�YeRۣ]����,z#���5:]��פKx�1��[H���ّ����v��V�d�Y�t�̕B�Y���]��&NH�v�/��G�}#����4�����ۓK��8��5j®<(��ӈ����da-��p�Y�����Բ�-����=7�J���/V9\����+�_v	u+�3��*m >�V��q٩F�����GS���z�0�w�V`���t�K�{hеF�Ђ�����O/Lf;��Е���<�r�OA���Ыu���J���Sٕfutdn��0stөFh��=��"�)|k��{}9�r��������}*�M��u.�r���L�,�b8:��D�Qe�;�ɠ�dTT�Ԩ!Y�l_q,��8t��Q�"٠�0�ʶ��<%�
ÛwǗ7\W:�l}�S9֍�-;1�ӷ5�%�G ���)�3�μ-T'5���B�X��V��r�h��b��:� ͙F>�Q�M��I�
Ղhx*���xDz���¸�w`�4F6L�o5��q�&����)�񭥂�H�|�ԍfe�}2Nu�|kV�!�����oAz.���)��qa|��)ԫ�K<f䤭��LdL�U����J5���NS�#��7of��b��xu8���׶�����uC���v���w���#�UVSo�x��Xj���������}�yl�Y�V[�μ໥���Pלr��]h���r�{��/$�AV9�t�Գ�\:��g����a�qc1e�s�(�>1��Z{h*�B���7�Y��hہ|���cL3��',B1���)3��s�5*M}���_cJ��#kJ��+ie%R�ciX�)oXd�iR����j� �*��*�k�Z�X*����R�D�8ʘ#V��,kF�ZV6ʭcF��JZТ",ZԶ�*�lB��E"�(Z��1� �j��$�RTX#*�-5(�,U��)F
�R�D����� �F�U(1*9L�B���(��j(�ET+(��Ȱ�V���U{t�뾞�z��1�ۇ� Z���fڳ3+%��r��7�\���ww���\ծ��FaW�VL��*��D"�bh��L�t��KV/����n�R���t�F�䤉�uq��x��.*����V*��M� rЭnj��\e���)͎U��+�im����}X�fpd�}�euSD�S�D#KD�C�7��rfKC�i���{�(Rc\�4���ߍ*�8��&�NSWW�s�n�wYj�<�ow���δV��4�0o��ݍ�ڬ�s)PF"Ò�=�kB܇_�����S����^�L�,����O�ɡ���ʽ�u�1Sy<�|�;o�+s�D#GB�U5�*��q& �R���V������Tq������iێ��:��b����{�s�/=#���NG���tgERcF�49uubu6�:���%�v�(i�ܦtq]�Z�{e �Ԝ�=�g��|(T���ߴ1E:��FwPe>��t�ye�������3�pM�w4���n��I�T�:�Ρ�n�	K�Ӵ��R�w;����	����e�:O�D�	&��So�#q�9�$)��%�X!�fy�V��[֚������Z&��w8��C_T2�{�ծ9�{�Ҥ���5�8}�E����m�t�^��^��~���q`��\V�T[���
�:��I9:c���Q�gG�0|�ʐ�P��=���H��+t��\���7��rZ���]�:�UgG^��y��w������u�z�Y͛�)���p�w-6��Av�8�����8��Ҥ��/��Yo�"1n�Y�՛�Ti�f�u�f�u���N�Pp)G$�
��y�*��+S����n�JNL�8�:��N���*������Y���/Al��0�z�{җ���q����3rY�O��#�F�w:"�t��Ҵ��2���N�~�o%h��O��|��Qt���^�c3�IY�ʽw@"��"g�=��c�JTw��qY�6����\i����[�$U��{פNu�u;$�95`�hN�L��U�l�>�]n�]���ee��٭���Q�)#f37GF�*V�\�eސ�	��;q�����v�
�6�v:�Z�����5�E���\C�,�gVNN�j@x�B�^�=ͷ�l]z�l�˛0^�/e�I�_At(�u{�P�R���*�s�6����s�\�U�)��S8������:�q��[���/�rQɨ�}��*׷��[A�r�]����{2p��%��3�|k�ұ��)n=h�jΫ�]�ܫ�s3�j���f�e���d���n@Ҧ�LM�g��X��Z��e�9l���+onP�D�*��5����4~�3K��v���jvt[����9udD*���a~����f83�T!�]%!�W�d@)�x��'�&�ϳ�:{
���ʙ"�dK%TS\n>%,י�y�8i�x���eC���ʩ���6�!��������|w߶��J�b�O��;(�\02�bx�􆽑����V�zf�t�D���D���6l�]R��Ov[����P��WdP2��w�&X����jY^6���>��z��y!ܻ;j������ �/�YR\��)n�Q�trJ�+\e,�w8A�ܸ���4[q�~R���L��t�N"��L��L���֗Jcu�.��A��$i���P�B��nκ��[o5�B���n�i�-�R�$�c�nv	�d�!I�YMZ���U�Ӳ�lPMSN4(�iӂ�\ٝE�u����N��{��0hB���$.�ix)Nk��5��
]h�mw�Ҭ���
"=� Υ�������|��.ɛdfe��l�Yha�����/��-��7��:�R&���5�t�N�A��+q�Xcӹ��aND�kD���VSQ},����kT���ך�R���ik��it2,嵵{ʹk�	[�{�]k_mnl�j�/���P^��ɾz����;�v�c���B�ˮ8�jly���$�9ql��_j��Z2�s���
�ڬ=Q3$`���j�'m��b�~�~Q��X�֯��'��P+Wg��D�tv�NlU��$�6Dp��B�Y]c:Fu���<��I��ɋ�[�Ɠ����h`�4���Y*�������4q�B��ٰ�A���K�ʳ���cb�`m�ۗ�R���fFd�
��h~4�7c�|̙��^�yY^��tٽ8��C}!�_ʵB-�T�&��Ob&�-����BR�t��b� dF�y�#_-%�`��������x�[�d6�����K�o[f��☍��xE��ұ�[1�;����h�)0E8��J����^�G�b����h�m޼�j4E<�j�G`�7!Pw��s�V#�;x��gx�)�>Enh��5�ۭ$���-�3�u���?7\���g�����UƳU��}+:(*�ӎ����ّ9yë�:��!؀�H%�$�p87M�y����,�^mU\����'6�5��U@�q��*�����I
��D^s�疑O�A�^�
+��3��	<�T9u��L�1go#|ՙJrM�g�Kw��+R�����働�e���w8�v�����؉BO?q�X����J���Z�V�<��[P�*��V���I��S���iq��hGF�|�|{�Y���;�Y�.��	��#��n^uU:��TC�N�m-���m�kq��m����}9o���cZ�k��NH��S6+5�ٴ1%�u7)D���.��|6��y]tb÷
�9صBY��p���]�>�(�`��{7��eI������+�-�Q[69
qV��� ���۸ֳ"ᶛ�z�pٴ�6rF��*��i.t�K�~�z��$@�}�~���"Ȅ��p��8��rh.c�B�6`d�j�����T�gi�_i�	�H�''�pIQDӒ�6Ѵ�naT���U��֧�!EP!H5����ʨ��_u�8����\�V�\��m��!C�ƻ�t�۶���c��y֥V�-����AF�TGY�&�ce%=�a2����)�$VZ�mϴ��W(�g_"��Cn)5C�*���c�mйC,a���TM���.-=JL�k����N�=���ܕu��%�Jl]��O�]���7�p����QG���Z%Oe�qj�6���k
���s/㹬���n
ˇf�_����82�h��c��#��������)��vT��[�ji�31D���p,�O3�(wq���#����D��X�x��{dm�ӧ��*����1xp��+H}75��&�R�!�6g�w��ħ3w��4�Ԭ�����X'��l��;�M��x5'�W5?S���w<o�T��H�k[�=�sp*[��:߯��Sm��Ai�(�P����찉�����Q���˳�7��������Z�o���%ճƓ�,Z��7b�Cx�I!_�nv5Ȏ�-GW6�'}5Č��Z�>�g!��ҡ�,�K��s�8:)f��We)8!h:��\��Z��2���V>UA�=Z&�B�*�oaC�:2W�*��;��{P�B������iIм�{f[ݡ@eEz�V:�l�ņQug �g�͗���D�sA޳��nW���/�Ny�V�"Dz;�n��ۭ����_	�7*_��G�^��It�K{����N�>$��y����4�$.��3��̻����T4_�	4���� Ɣj��
sȉ�6�J����_uv{�����َ�|�޹�&�cΕ�4�o���lv��5���=���N�:��h,��:.z;6�v��N�����#MF"�:�N��k��K���y0{/���^ ����J��O��V�E[�%Us���X.��� ����U/bZ��r�j�5x_5:�vﱜr��\����.6�L��E�am��^gp�"-3�m��Z���I�s�E�'1l
:Mj�[8vٗQnv��ʧY�+�@*$VS$��&e���e�&�칝u2X�Oq�݃�db�
[�:[ltf���j��Gn.�iJj�Td��ժG�y%h�4!p�����%�Ek�'
4Ź.�Zuz�:w�*śڪ.�r9�(X�A(��|,��$�yjz���g
7t:�t�XGo<H�'ld,�B�l��s�J��&<��\��]�`ָ$��W��>�oTR��;{b�k)�Λɧ��� %�u2�i�
��'�G}�]�=�C|0�{��H8�eӳe:z{y|�P���i��w9�@���l[lV1�i�d��R44��5��6���N�nL5��鶉���f�%>װ�0[-G�c�d��d�����0��ܝ���:3��+MAc+6�6�Մ��٬s�r�;��װ�K̸0N��`�U-��x��ȭ�gw"%3{��
�Vno�u���^�$u�+�'m:��{a�8��u�7t����4vȕX�/�pUW�Hq��чͱm��U�uV��7 ��[�G�	��
�:q�$�g[�a�� .Л�A�`xn�83�va6Tr��:#k+E��作{�60(b�On���{]�r�vWP6��Sh_�� �R�� ��۷ܻf�������:�di���%m�k���U۠T��%�u�� z?48Cک�ᛷ��Z�́K��sZ��&��Si�����8EB�{���)r��䦸P��V��u�lU��nd��2��9;g����kj����|�%/�����v�Ò���iK�iYĔ���R�F��^�iEx����#Th�Fۺ��y���w���M���ZN{��Kקz'�� �h�@�3����㼠��y�k�3@����օ#u��y�	�M����(�Wj�7����0��U#݈����ձ��KR^�ʝ�N�C)XJ�]1���ӭ��G�lT;�V��Jv������L�r$��w%1ͫU/`�)���e+V[�ӵ�t�m�2%��Cv�*O[=�[��Eʈ��[U.�U��9Km��-h)m6�ı��EV-
5XVb�[V�+PYU��B��mb�iL��FTm��R�)X�*T�+[HVV�i�(������m(��dR��%E��j�ж
Ɩ�C2�cJFՕ
0���Ŗ�H��Ҕej5��RT+r�r�*Eb��(��ѵmD�@F���E-j���W.eF�����ڥ��@X*ƴU�hO����Ȣj'��4sΆ�$�fs�e�*q��ra��̱���;��Ҷ�Ge�C�3��.IǕ2���Ct*ŷu��t��bda��1W�V�.iA��H�ʺj�F�R};�f�����N;w�C�KQ^"6s�B��m��������+��H�vC�C8ʢ��WC��r�FR�͡3oy��q���9�;���pn���Gq��<SZ��4�������MPF���'����ڈKX��VDM���������7^�ȱSs�7ɭ�h=�9N�eYZ.H��>��o<ն*�}�/;�{9��1�Щ������e
;���Į�i��%��S�V=G�p����S����de'�"X���ۨ��vk����9��<�n�uP�iˬ0�L���^��AR���m'�t���=��d���b�x5ش	�+5���Y��&·ق��SY����h��|U�
7S[3w��z�Y�)���/�
k~�|:VP�)Ϸ�/?'ޤ��x���*tn�V]!u���PQ	;�$����j�U�YI��eX�t�o l��=zOJ��j}m�1�BUr���?zq[�d����L�5z�ħЯ�F)��{̈]M�Ŷr�Ŀ\O
�o�0t����b�*AH#fK4�s��i�h>�i�-'��uR�,W�U�*=��"
�XG&�&󯞍�_x����"�XkPm�~��ɴi1f+�o�\!�9�$��[��LX��뜭n�"ұl�l�\��S��(g�����׽t^T!���E����Z*�n7W461<zl:�΋)-���M��t߅3�D����Q�%ӡʵ��-���])x��/"�)��.�f�ǫz�t��^+�-Ǡ
xc���c�z�����k)��.�m�m$��n&�l7��%Kނ�,uÔf�N*����aj����_"y�tX����T�8'Ǭފ��K+j�o����
:�+U�Rtd]���c�ݕ�;���NSG�z޲ڽ6�ˡo��p�t�y�!X<�B"JkE*�X~�Op�o�g+��[�3X;�S�-:,ݐﴶjn}#�#���gL5��d��'���Ŷ�>,-}Ĭ�$0h��O�R�Q��>�\'Oa���IBLbU���J�qO�'3B2r8��\���a���o�>�M�!�*A�'tb�XqOEۣ��4d������yB�uJƉ�KW�Y{���X�(��t�ظ���ٛ�:�ǫ`��-C�����N=���BؑQ�=C�	扙Y�v�	\�C�O�����I�*q�Z�*�k�n���bP �+:J�σ�{�#)0$cS������K4!��6�R蜁S��E�9pܾ1u�S������0���.���I)��'T89�ڊ�mP�J��M��o,Z`�'�:����*B��v�]�N���2�>�i-���6z��#���g�bi��(|�Hړx�b��:�Z����Ƥ(lֵ�ʚDHF��&�7�t��JP�:u}����Y���v*�0��5U�2ڼ	�7
y�J�ܵ��_�ֻk �u��������ޔ��*��/��,�5�����C��ҽ��Yt�����I�H����ѣ�z���������Ҙâ�U" d�}KZ��9Wd!h1��}Wz#Rhs�3a�fh��\܁Dݢdu�P.�Pon�=����SO��'l]���M+V�f�K+J��wҤ�Z�xzp<��[�����z�<Ss� r3&�P�7���-��KZ)RQ��k�Լj�㝍��iG:��!OI��Q�B4'���	x�b۱X�.�L���b�K������.��SDd�R��Rt�ڝ܆�L�=�:F`C������ �m�n�c��;gYE�N�0�T9#^E�戫�jE&�ث)�Y�/ه���bAn���b����f���Y�V��)�I��z����@m�,�')�f
�w���5�:IW�9���Ǜ�KQ�-�o�7C�q�<1���N;�󯁔�ޝ�Y�o[V�Wk�"ϋ�4�flB����[�jķ��a�ݓ����>U�Ȭ�/Ҟr�H�� �.�V�����0�)�[9Jri��.���oC�������ڒ���ƂF4'=��*����˴Q~c���N�.�w�5�;�T�����)6�']�c�ך��)���;u�;{���ڐ����{k-���S�{�$�o��;�#���$��v���s�W�KX�;/z��Me:m{W��"۳���}6�;�j�{�&9�N��fp�[ٲ�>�B�cw1��(.�M�?3��z�fSj��l���T��5��])�=�N�M�KPRɁ���v�����6��mNk���A2�r�U�Q�:&v�ե®T���Ym��eu���#ɜM�@gVl��m�[�\�)\s,h;��4��������sM5g&c��L�v�{䳵9��χ��`��IQD���-��[V��A��Iٙ�lPMPi�A��r��I�,hI���:�vC1"��j�K�C�`��4�ai^]��I�z��Ͻ������'��?���3��@�v^gzѫ�}�x�&��'U/{>���t�r��FR�ϚI��ٸz��*����+n�w��㚥2�)�l�D���_a��"��kPھ�(��M?I:�X����t��s��e�i��C=���nE� �<5����l���ɼ��J��c�|�D��Jp-bCʙ�Bs`U��p�ޟ��T1c�<Guĝ�W�&��/î����JYj��{�b�z��vs��q3�f�˽�}�ދ�ӛ��.<k�r���.��W�ܜ�_Tp�;A�r�ʚq�fp�4��J��	�l�&���3���N����02�3WQ�̸B/� ۮ�����	�YO$��w��~���E�����
�4�8!σ�_���_l�\���{��6��ʹ�*5�{��9�T�FiO����)�wP��
�r��E����l^�dg�cr��{� !���"x����\�f�G{9���\tS�^��P/%�R5̷AL�Hp�(�p�*33���tǏ�@�zC���6�$�/dr�p鈉��3{��M�B�xϡ�Bz]-���t�5���K�j'�O(�O!����@�N'b��76	�d/��B҄1�����!G�Id�c��陻Ι��2W�����а�ƌ��Zlz�}�p(|�k���>A5ޞ,�>��}�!�F!����_�>,V�l���[�H�r.������d{��v]���/�M�q����-��{]�):���7��3W�&@꼪�f�����AWz�y�h�s6����NCs4�D�8�S��c��e��z72X!���\rwa�gȊ�K��꺮�����S��l�J U�K����{���b�/|ע�ٓ��k�v�]+$�U{��SC�8m均"ꦸ;Ɠ2��+Dc�Q{�=� ggԝ�K� ��N�X3ѹ}�>n�o4'�<��p0{��C��>)F��cCǨ���] %v�Dͯ��4����0u�/�eFU͂+�S�ҩ�R��8�]Bt��ִ<-<R����q��gں-���0hQ uHqP�F���x�kAg���O�i�x�0���W9ʾ���c�`�{�5�1j�D�|��W��#bi�p�ИY.*r��uv��L!]�\E]��Q�膽"\�Nت�A��9�W���j6���t1Cydl����ڸ��a4����|g��/eA�p����6b�x�����y�P;J��/�� �kۮ�j�`�Į�ٽ�S\�x�* �)>�WCV.
����[$�b�h�V[�S2֦�vG��V�,����}�JVJ�o�]ݨ���p����l|^�+��	XA��j=�.���]ə��Y�^?#y:>Ao��l�4!���	t�����ǛX����`Ma��MB >�"����T�����wn⓹���ԟ�S�5�\m���~įղo�m�h�ӗ�v�֗g�+����#Â��(�l{>��l��/��R��b�}�!N����l�[�F�m�w>�3�]����Fh�
+���q�*��Ƿ���	���Kݡ����^�e�>�t�/`}�`�<�� ]͙��Q�f���"�c8�a[0�����=fR=e�w��ݟ,���E.���Pbje׶�@��1le�����;9����,��$4F�/�(���c�����9�?�����ߵ?=+UUQr� �Ɵ��@$�?��$��	!�/a������<�Ο��}k�=����L��HCH� *('��� �~�g��M��~����P�	!��`��ğ?���z�u���NC��=���nî�6�܀���$��==�w�ǡ�q{ۂGG�͝O:�ן�I\������~�����~�$HC�'Đ	!��XE����ã�!��~p��K�(y��PF^� ���9��HE��w?��3l�
w Y�b ����`��k�p`�0~0�L�p�~[���tNP	��/�Q� Bȷ�5�_ɣ�2w�B$!$��C�f�!�Ҭ'��^����>tP9�����؁ �z���qME��`B���;w0̭�ڑR���K�.��ЁΞ^��b����@$�qL�t֋�O�K��P��c_&u`�	�w�E���TG����ԟ==~C��������P�/�9�����=���'��""��@��t?L���?�Q"~g�֓��,�� �����`������P?���d	HC���X�1�0P���zO�� �c'VN���v�O���uZ�'������'}��A�2��B$�c���H@$�l �5�� @$�G����-v���x܏q�"��}��rP��⭋���eeo���������M$##R;v�&n�_r:� B7�ЈK@j?�?�������?l��3��Iփ�:�8'�O�r#& (6��V�9R�
��X:��y�J95eCWG5$���H(�FↅϾr1��}C>�`a�c�|�IR�?� |��I B��'�g���������:��$�Iޖ�1m�0������,��:�,�����I?T�� �Ċ�&��H�
	S>�@