BZh91AY&SY|)�)�g߀@q���#� ����bG~�     }_f٤��j��ͤh �L�
i�QB� F�L��5�Պж5*+L���X©MU(
THT[-�i�S�٭[c�{�RTY���ikY�����m�֒J[m����V�hĨD�U��e�j�[+%*k-�����L�&���dZ�@�Z�`�P�;U��mQ���)�%jZ��0��"�H[*km�Q[bM��j�����3Y$����2�XU�LP��R�f�ѣZd"��M,�{���}���؆ �   �9���vc:ptD�X����Q����[P�;j��]�ڵj�N��r��.ӭ�vcn�Z�m;u�uJ�{w���H��L��[a��`�   �w�):���R�Jq`uB���u��� ]�b�ҀV�;�:
��ƨ �ݪ�
B��
��U�zʭkJ��l�k+[[   ������-9� T;9�Ҷ�A�]Խ�=P^�t�kmJ6�w���J{���AB�����B�T^�o;�+���� (y�^l D�iD*KF   w{�t��ޓ�t=�t�()A�y��mPQ칽�h
Pw���z� (�=�Ҵҝ4�z� )֍��h ]��;B���wl���m��Zd�ذh0O  ��� �;���t)��\�\�
 ]�� ;c�':���	�pu]��i�6�B��k�T�t��@6�4Uk6*�4���
�  u�� S[�k�  ����V��8)�N��p(
V8�@4m�3�٭PQt�MA�u��B���J=��Um�4����͚�d�� ���tU9�� �� �C�f��, �T���4	�j Q]�1�+@-]8 P�훎��<�{��V����[a�  � G^��]�u�p (�2� ��:��8UGuuk�E�7]㛀�;�ۂ��{ț%l��e�0�6��*�\   ���@Ҙ ��u  ��� 0w ��W@���(v:��m W�( �Z�حb� 5�@Dx   wx :.�  �  ���r� (7\p w���l�� Nvr��k;�ƀ�    �   50T�J44h4 � )�4b���2 ��  ѠO��IR�      j��@��*0      EOަ�P�S� h� �a	H��D�L��O��j42z��M�M�u�n���g���o�]��+S�ʌ���5eߣ�^[��������� {��O �*¨*~�����dW�?��?C�����?�������#�*}����
�?骪��t
 *��OȄ?T��QT�����wj��P��	��C�&�,!���?�xʞ2����"x��0'��<aO�"x�2'�)�"x�0'��0����`O�D�<dO�T�>��T�̧���*x0���� ��>2'�|a	�<aO��<d�D�>�<dO��� �ʞ2'��x���|aO���8ʞ0��)�xȞ0��)�*x�8S��82'�	�(xʞ0���(x��0'�	�v�0'���x�7l��x�0���� �`O��<`�<`OS��|d���>29��|`W�Q<e�D�e�|eOS�T�|a��;c�T�|eOG�T�ʞ0��)�/_S�A�|a�T�~�S�Y��<dS�T�<aOS��>3�"�A�|dP�^�U������ �� �ʠ���Ȩ�Ȉ�Ȉ����� �ʀ��!�� G�PG��QS��PS�S�AS�S��QS��DOQN0��0
�0
>2*>2*�0�>0��0
>0>2��d�̢���
�
�����������/�����"+�
 q�<dS��<`S��<eO�a|eOG�T�<`S��<`��Ȟ0���
x�>2'��*xʟ�D��2'�	�x������m�|�g�������=��ȣk�6�ze�hb��҂��X�m�')�cɷX���&�-ԋլr�2+Geeb�ۦ��W0�`�0��cw5^rT�ɾ�6���,�)9�F9�9��Bq �N �U��[�N���|���hʹl�ᶭ�r�9tMΝ��բ���'1�V%����o;fq���]�A�a6��1f�d}2Uu'ENS�D��� ��_ bZ�y�rj�Pn>�,Vܖ�@웓5��nUݹ���sK)��h�ݱoQ�������^�����u/:���:��ҳv�l�����˾�i��^ѡMFAЪ6�ZK�a����!���-r�Q�M��V�1�W�;���0���k�[���� d�����p��ܚz�z�3`��d9r����Zĳx�փ�0��v��hm<�5��M�y7��%Ql("ut�c�{H��
f���U8� ���'3�$�OS�K�NX=MuJH��oS�+t��g��Ӎ6��3?���9jkqB�eKg�c��\��wq\���hh,P��4�w��qn�i����{T6�V��f<&�w����1!��b��]�ڄ�ې�R�8h�����1ǁ7f�\ٖ�Ɉ����J
"l�
NX��
���r�&���߷+�w�]�xu%�՝�f�S.�(�꧘zM�D���a'h/t�,��=�J�E�ʧH��ɻ�Y�"�J|�ٗ�7�r=;lw��w	ؚW9�}����m�Cx�-�1�4�.�Cs�]
���"ɼ�0�׽T\�E�z�XV��:�$�]$-v��R�So\��)cP�u�aۚ3r��Xv��=;��=	��d�LS
n=n�r���E�ɳ���`
��+���y�m�����dm�sx��t���:J����5꼢l`6N*Zބ�e�zǶQX�꫃�!wn�A^�
Q���F2�V�iVmd��BP�?��C6 �6l.U̹ba�qJ�JO��*�Jw$��r�M؀!q��+�shwp!i��M�n8d�۰����5K7ᘔ��)�C�,*�Jƾg��1�x�hT�DǄ��F��(]���p��wiV;f�X�qo�V&�D��-���;��,�7�s�j"p�L�ܺ�Z��'���=zCd{����[��
rn�Ug:Kۅ_�D���@[��T�D���w�Bכ�=��dĴ����"Mp��s�3,�c�t�S.%�gv�JojZ�<�(rW(�!�¸򸷊yHWH
��V��j�!�^髺a1��l�M���	�.=��ޓJ#�׻���)� �ߵќ�sgj����r��B⭰x$��\QW��nU�v�'�W��sՐG������c�h8͊bl���tƗ3!!D,9�1B��qY�{���3\SwC�s�$��Xico<��FU��rTn�%�f݈l4biE�f����Cn���^ËPW���g.�r��'i3�i�]f�,�X��|ś� :��w�-�k�l搒+��G�6l�:'n��@��a��r\�k��j�v�N�6ɱ�[,��PPv�S�(blM�L,YQ�M6�̭�hS2�Ԅ����(�;U�N����ѿ���k(bM<�X$h�c�du�*�Ê��n�+��[���w���.�֓4����-��Mu�oZ����ҭ{�j�z�n�wq1��ڐ����*����}\�SM؀F������1�8�}���&����:�v���mf����3�Z<��IƏ��ޤ-�YJ|"�*�7��a�ۮu��Kĭ�$�Ei��'
��m�Y��d��PCN�X�uY������_!���b;�vk�n�eÕ�FZL���t�rӼ��1|o�&��wʮ�,x9��x�6�%eE4�u��hAۺ6�un���nj3Tp�)<_��&v.�.�*�jm�̄6��=Դ��vv�V�/ZUgP{��)9�xU�M�7LN�w����3�p��;5%ܥ�%��%{����]"��R�O�!��f�ʥ���O���ۥ�}�	Sav+(��=F3
w��f��f�*e�и�<��\\��!(����%['Λ>�y�]���(T�*��n]�T��j`��!�b/H�*V��f�!9y*��!AS2kڠp���UL�ĳ�+��.���H\�Dޥ�oa{8`��w��Z��',G�#�'/4�DO!<>P�;'�v��h��y7l�ܯB�}:�����:�Ό&�ȋ�C�Z��B$V)�q^U�Do]\�E���*�I0b�wy�e`�Ff�6��ɥ��W5��γ^�A.�'NwP���Q�v�݃^\4�tn>Np�=p���[���{dE4s6ŕ�M�q�����jpNn���>���q3��&��7u�Qf��m�2ܹÃռV�};�j�6<�2�X���M�枙��C^ ��P�H|z�򁋮�;�R�yK}�c5����t\�;T5�1�r�^s�:���h��ʲn׹w���RM8x��ġ�H@Ռ�in�y����q�rc�0^�z�6�\V췌�
v�6���I��͓qk��-��j��S����7�nA�AW:�!��74jKT@��k��2�	L��q�v����)�ӊ�.u�����\��V<�o+�,կwopZ�a6�X���Xy�v��y%�n!%����*��nHw�����J�*Y&�t�ز�ӹl�h�&79�R�i+t�[�U�u|���K\ՠo�5��n���j�v���1�K.Zt:=����C�ą6.,�{{��v�ƶ��,T�{�3�{5�vƃ�lXd�*컦M$M����ա��"L�Sgi:�6�T8�R2�ٻ$2]�p���C�t#����e���NG��������&޳�H`p'FHw*>e[�g r<�ᛍ�h.)�)أ\;�;nѥ��Y� "��N���oL8,�q�s��f^��B���;'�g�֢vՂ��?���ۇK��.�+��ur�e��V8M�"v�]��U݄�[����0�B�:"�A:�;w�4.��;R��Wc�*拶bǗ��w&�����҄E+;k+Q5E�v�74ղ̔� �wG�RM������ �|�66 {F]�n�&�֗qG�:��ar���{��F��׍�����7�ѝ�&Qh�.�5��/Zt�-� ��9��OS�s���Mmɹw��k��N^���h��4F��1v���|�s�G� v7�=q�%��ٙ]�&ݬW��,�X�mt�Ժ�C��Dix<��T�9E��>۟�4�1��0��0f�F�x�4�jwY�a�T��%�V)�3*�4����U�7����]И�餠.���VR8HR4�0>ai]	�ztp���ע�dҩ�ZP�a7&�3�g5Sczwip)������s��t�=	K�3,�+o&���/Q�F���R!��癉���춞Q�9��TT��:ԗP0�� ͳP�z+
�V�A�� � �:��'w~Qm������ٰ�9-�C�
a����n��m�v��r�^2�����#m��A*L}���(�m�/*�A��wU���Llg2ͭ䡤i��+��v>P��7N��J�q�m����P;-Jb�x ���餠�j�:�\�'f�rr�����+O�77����F��S� ���4�IӘ#u1�⣘bd����H�2���u�^h����#��SNְZ}D�����#\�)v�>��gX{6>'{Ғ����AŶ���f\�Hv�,�:"V�h�'�Z��a���̐e�.�2HBu��0�a��ur��epa��Ἰ����3z6Ά��#x�ʰ�E��#,X�)���˷���^�hpS�!<.�v�:���^���sm3��[jU�dˬ���p���n��Y�P�x�A Z��l�h§�1܎�UR.[7K��N8vB-x��q�3֪xh�� ��>'r���<��c����m+_��(������S&��vߙ�'f�����k
��X���q�����)�Zu}NŽ�|lT<g]�Rݷ8��AY�٤]�9Zr.�巰��u��m�G΅;]��ͬݩ�G$�1Q���Q��+�誼g0�{��0[t��G-���.��;�2��Q�o(�X����KN�He�doTY<�3�gY
�̇2�7����f�Bo�Ա2�k5���t��r�f���Lܸ�4gFg@E����M�y���`a,�M��r��� �nQ�6JJ�`��u���O&���"��X�@�c]/7(��S�zW:��c5ՙ��NQ$���ɷ�n�mk���Y��`��y�v��nƐ�ˁ+c[��KӘ��:��dL�[R�)��M��>�J�[U+)c��-"��6p��L;�`�ٔ�V�
���踝�:L6�*�!����Ĕ-����Z/yv����P�׏rK���O��0����2��e(�Ak�g�X�,��7y��\����r�h��g*�Fsw#6��fƠ�4s��i���Mc��f�����Yk�ܯ�Gm�H���^b��j�R�x�Q�2�y���ɿ�P�i,1��p��&�����N��.V%�@�K�Y�l��lJ�'u���ܤp�I��ՕwZ�?�{�v�h	o۪6n���5.��.�(&���w����m��T�}��j��v<Y)Ij�W�j�wH)��C黓p��9X��{�³�f�gD�:�i������PC�U� ��z� �^�0+n�6Ej"kE4C货L�a��[NNbBMK����o89%�4)5��(�����J�v��.A���L���hy �n�f�ܺ���ځĊ鶳��#��Ƈm׽Ҥ��U�o/�ުX��Bc<�7�+���]�yY��k���޼��m�
�*/.gq��m��v���Cvg7�ݼ�Jm,7J�E{���� N-��{�D�rp�ٴ�6n��~Ln �t�
%F���Z����خ㜱ί�,�p������x�ہ^]��z]� ь��qD��R��M-j���V5�e�@�Y�]�NR8M��Jk؆û�h˛��t�^����˧�`V��H�Z]];:L
�����m�y��� ͔u���tj���ùئM�7��t���3B�I�����0ڬ��X0(�/*���3+�Ѹx�E�Gb����9E�q���i���1Zy�Fk�~�dʱ<���%�&ڳ�hjV�t��WoݨAΞ���b���{5=b(n��.�X:�x.⺥�38�Pc��p����FK�� �C���xɺU��a7;��z{u�VE�Db,҃���[_�k��뛫���t�RX���H��R�d�pm�5���Le��q�ar��K�Ղv�����8t�H��c�EF,��Hk�;�H�ٱ|�[��;Ӯ�0\�X̵�+)�X��8�c��2fq�[d��G4:Z��b�U)�N2B&��`+.�]��.��~�}&���d[�^��1�'M�w�Ng'6��m�7q	qԔ 3�S}ǁ��2RU��ۃmy���5�/B<�#Z�4�1��6�pJ��ƙ��Qd$����g;]Y�3�ԅmi���sd,��z��YZ��f��\�'P-�� TX�w��Pb;�I0:2^r^��)�M4��A������c�ʎ�d�k�)�'�w�y7�����(of���2�of.��Ȁ��ٓb�0�7(�,����)m�ù�f�s��'Ne����G�{�5;߻�����,�q;�s�������8��T��F���$|��wv�i�����+"p9��9y��t{��X�Ť��n�v!a3*������$�&\�/5��.أ4Gj#��.��g-�E��i/���yɮ��Vh�{��mo�c�xM@>IՉ'�h�s�8)v���O��w���U�N�4tn�!����su,u��Y�*4��"���;��CM#�@N4�T�e�ڻņ��G��eܣ��f��=�C؜%��V	����x]�I[�/ASm!��s��T�+ �k,AWXpۉ�P�IA�<�x���W7��Vb�Z�,�Ot�h+Z|�0��m(�17�eD�K�h��]�n�-|��̓O��.�(jn��	�䱐�Ɠ��t�������wz�����;~+S���ç>����͹�.��� �x�_�Z��P�U��]��M-M��u��xȶ����'��=(FI��\��Ɲ����c{�Z1�׏�8���b]�B*�#T�It�V�ؔ��{b��U`^�Zo8/�op�s���Vؽh᭽�Gs(!����8�)�y|��W�}D5�U������GH�G)nM�(��ŰLɈ���B� P�F
��if��޳zJ\�������Ɗ��CjޅF3�azt(&
	�,�(I��Ȃ��#��(\�������֮��RDKbt��r���5@���ݽ �����a�P�xwݨi�����p y2�(1�RK9�]��A ��:���H�B5%��$*�p^��A��uX�J�4� �I��֖��048PT��{Y���*���D9�ع�m�NXÅ�@�m*��,%3�UA#B|ձ�u��C��x��X_ݣ�^N҉��į���+��RI�嚲ˢ���&�U�!�`�QWoJt8l�p,L�t(-��U{ͭ`'�Uط� �����<B3{`,X������~�����v�h���k��������7�����?B���?�J���?�s4��N<n�w��m�jn�[c��Ea�}���b���<�kD�&��,��\$!c�y��o11��u�Y8,jy/�����B�&�j�j)*��5v�;�#*\�F��'	|��5i�����)՗�kF�	ۤ3�	�ͨv��nͨ��&�����X��� �����V�|:����Yx���u���,�˸�*�|�d0�Є�#�CЃ�����>�C�}}/��/�-���d�\����Y}iN��XX�Nˍ�U�n�4*������ŭ �+�y����W\z�wW�͏�{��֬���>�7+��|��$���]'pk��G�\[:�vz�蛾��,�/���*{��ݞ4<��ºT�mK�»0ǫy����)9\O$/5 ��G�C�+�rIB^�Qn݇\[N���]W�=��bF���޳��D=�{�ҷ+z�v�fʥ�e�}E��]�5ݮ�	��wVs�������呩�p�Ym�l�?v+K��&��m���-5(H��t�>6�{ގ.���[�=2A��k�l%���9�yu�B����W�u�u=�d�{e��j�oy>ц"�}��]�T��u�GB�
f���m�}z��3�޺Ň<x�sy����1�pA��x���>��yϢQ�͆o��e�r��=�)�3�}Ok�S���#ç2&��t���N+�P��)�8�q��ǽ4����yb�;���+�8�x��Y���\��[{�Oj��us�1'�[�^#N�{�k΄���5�� 5d��%����x�*��l�k��>;��mlr��c�*�]w^����0ۖ滚ʦR���X���zw��!G��Ε���n�f��M��Xົ��H�9S;�7C��s�'�{����'�K�6�������)j$�����1��x8w+P�=NBh:PV蕔�sK̉:˪Y����*Ec��r����8ma�O^q}���;�0[������id:�V�So���,�^A|��2S+UȨۘ��IF��\[�G(Rv��I�N$�m��yU��^fK��«���7��W��=;i��V���i�훍)�Z�,�˺�]��84��?T���������ލ�g�ŏL�_$��$�%�6:�^�'��C�W��U�����7�ƽ��q��96�q�#��yW�,���2��"��4֭��3��K��!��v���o˳� ZT�C�G����qjXs���Ν,��3E��a��뫹��.ko�gm��U��d!s�;�nk�]z��
��&POV'E��{��YV�:�%[f9{y�w�t���'B����~��ɏ�sD<�m�G�G\{_E}���j��c�v�|�iMF��I�t��ܽ�@v٘�픗���;�s}�[���qC4Uf��ڄ�x��RoՐR^<�M�Z�[��.�����j��(��#����fUaO����%�<�5�i!�����N%B�����SuX�Mc5���v��`;�:l�u��sS��ҕ�	�V�@���]�-)��&e�m[Q�ڼ�)N݃�|u�?!r�y�p�r��`3�
�,��b��ͧ��w�#��O���P�5���t^=����^��;�`ջ�n�D'Yy��FgqiHss;�b�q���Zgb�P���w�eh��A	��钸)l�yv�nQ��ck�cd��Ɗ�x9�W�p'�%6Gۻ�BJ\��2S\s-�h'�����/t,�t����F��mA�\����Y��-����Ԭ(eN���%��=��W���6�Vc�&(h-ʮ%���Ko:΢��"��}Y�;��W>�pz�1�P���J�[J�+7�ľn%VU����x��*dr^�J���a*� 뵆�����e��	���k~4v�}����B�6�kB3�vtU�H�ϟCWy�zQ��Ƿ�+���E/YSA;�����,$f
oWn��Tx�m��zt��m���#'9"��z�u�p��/�$w�'����09�p[�>�f��B�����P[|�8#�˼�GV�W#Ae�b��=|��7:����4��U�l�#�O]�?>���,Q9�{��9�u=҅�!�]�QK�Yl�9�Z�c��Q���pz�ң�������T��WF��2����(Q�7�v���;�4:����QgP	Շ({kj�	��g�@L�k3�h��W�(���`���T8�9Am���9�J��S�Ձ#�{^�=*}��ԉ�|.*�z�enۨw�$2U>�}kt�gh�on�V�Rُ�e�J��+��
�<�B{6-�ɳ9=�˺��=sf�:��8���h�R|�x�-�ʗዽ�2�	����n�X�4�-!�v��</���r+�éR����b^�h��<C(2����A�49�g5�WVh�%�"ksrU�`��j,^���n�M|��oG�R5�/I�4��Q��D�k{5��/B��'�j,��s���(���೧p��}4�{�\���͕�������B�9�����g�es�FYR6���eG�C��eF��O'r�(*P���Y-r��-�q�Z����r�l�F��U��;;+��A�lt{y��ik�-jl�^Ėl���obzW����&��֊��+Ǘ�Ԝ��>)uk1�,��ޏ݊1�X��݅�o��x�5�E�:�f�,�/b�dc1v*M��yl�z��\�X��7%a�ۧA=��v�@��F�LΤ�_P�۹u��ؚj�r+�R��fª�K�yǕn��/9"E;��#���˕.�We�i��K엮�FY�{�&q��3rj����j�"��ֶ2'v�v�<�;M7*}|$f����������������#���*�o�{tҍ��6N��K��MQ
y��i��j��NH���J4kk(*鼸���lV���+�U��O�̩���������2����5]'en�z�cG��LvO����Eݯ�t=s˽���K�Kj�>��>���Q��pɡ���~d�{�Ý��{r�4d�֯%7�ok�\�\>���]��+E�O�/-����3R����Bn�SvӮ��S;���e�Vo��/e�=����g�4�.0u��,ݴ%��|�q|��i�]��p�f��!�M�6����c�p��M��R8��Qw�w�������6�'n�e���gON�-k��-b�o{=����I|��s����]/D]ݶ���m�A�a*����*�Ӽ���ifGq�+s���a1W�rV_O�V9>�v_!ɍ�y��^���t�������
�G��¢2s�����V'P���Y��h�#B-	��a'ϳ�+;gw�0���S\�l���G+2�LWų�gZwx�q�Al�â�+Rۏjk#����K1ʾ�N,�u���T�u����}� m����o<���u�]��j�A�A�j��k��ybLA#P[����� r�.l����{�Ř�i��Kh���}J��A� �QҘ�Z##��۽R�aO��y9�H�-�S����#4���r$��U��b��CI8���^�o���f�w|�Iv��V�fu����m-������XZ���y����Û���^a@�/��¯G/�L�29��\C6f�*��]��I
5�$n���gF#XWr�@g��Y)nq�[j@3�ůtΗ�X�Y�å��'�t���i�rfu,�"��&Ss�Z��#'s��Ի�C4�+l��SMuO[
y��o̪�}۠z�S��Z�*�JϖV\Z�v��2	��ޘ���[8f�\7��J������-�e+`B��D�3���V�.b��e��S�s�C�a;��*V���,8��=M�M��Z7홽��Vf��ے���^����!���V3�n�B�;ɗ�'T��Rb�4�C&hw@=M��9d7�]�����*�k6�b�S��4:h@��K|#��=�E�t�g^YP$Ѻ��od� �b�K;ݻoT�11�5Oq(ˍu@YTWI�^��"�{���v��1���}��0a�Gnӎ;D_;�g�Q�oR�n�Tv�֎ۣ)y�{p9�y	q�zpb�M�o	r�ӓU�ִ�+�IB������AE�n�rݗې��i�D}��nea�֌JMc�&
@����u��	�v�6��>$+��:+T��|�b�^�����m�������fM샻�xm��x���F⹣#Y$�d(���_7u	�_C���|g�XC]s���ٵ��^n�e��ذ�Jqf����3�����Mv;f^XVj���|��]>�<Ȟ�z��{l=e�z�ɳ�	�ږŌ�\�#%���������H�2� eҥ���{�ُ�=�)y�4������w*�|M�.�v)ә���Y�9g˵>�����nH:��/ ��E�%W�.*�g.m��^Ax���*��D�>�La"���-�*%�p���!H��t��g4����P�q}�����C^L\�,cϢ�taɑ�&n=SiX����i�ox�^��n�{jKL��"�ys��=��=�`oN�ѹ4:�.�ֆ62����T˝A^.J�3R�3W�=5{�,6.�,&��W�~���3�K�V���A�u9�3���O}��}�<w]�	�չ6&F��'/r��P����u;ɻ}�|&&'{���U�_��2{i�P��P֍`#�
�.��:���Q�7V��-��Z}�:�ގ���Q�n������SW/,��1��}	�KN8�"460��oN��R�k�C�t�J]x-���w��}W(�kť�;cy��g%���÷���i���pkz�_Z!��<��j�<,�Ē�HB���6�\�*�u���Ae+���6������@"�i&��jQWuڬ�۫��6��'�dy���u�k�g�LN�n����j�^���/p.�9�P����FN�0����nU������)Xî�{��C�>��'E�&��+�T��X�"x�%�i��e�z��Z/��K��:�2��}�Q���0���Β�:߼7bg1�!�R�x��Z��|¬�E�Aտ/�1��^)p���z��v�CLg_�Z���� 6�̽����YXj�븇��uosOd���l^��0vL���i�j	�Y��71�e��ν�Ӕ&���͝��eb�c��������z `���1yK87����D�.Q�LJ�l��m��q0w�O#�q����H���T1��L��[Ձ�,��\)/n�֊�|����q����˴&�7{#̳�<����N����J������Y=u�&̕���O���s%�c�8d�L�`�}OP��j:	�ڽ7�[�z%N�G���Q^qÖ��H]̻�z���{�w�D��T��S4�=N�$q͏�2�.�"7#��]�Zfݪ��[�u]9I���M�|S,PT7xC[p�Y[0v(��p��MN�`�mL6�s5kQ��\���J�" binބۜl��B+8;K�����OGW;$���pػZR�G��d����8h��{b-|v�
@I�\鱤c�*�����G�<�u���4)�JX�y��)9sA�� �6�w�O^�WŴ������~I�.��ޏ�=����?���A�7;����N�
=���.�J��zX)��:�l��L|d��bI��>ܨ6g^պ��<}�v�x�0ڋ.��C.�'M:��Lꎣ�Y���E�Z���^p4��=�{s���ڎm�嬝�n&zDK�k��yA�
��}����JnN�_u`��
����y�(�n,�;��ٷֹ�p�e��v�CnVKM5�g������Tչ5����� �����Re,�N��36��́=��s���	�V	蜃	S�q�:�mr�s��_=� S@�,+%�%��X@Ʒ  l*I��m�9J����)�67V�	[ԟo�z�n��|�����6���Y'�Ҡ]���W{(�ݲ(8.�<��(f�P`~Q������>I��LLwR�t�tz��`n�����p[�����&���ϥ��6�K|�3�/w�h�7�QK���z�\{q�`,r<0�L��Bsn�W+�0��gS�p���m�;�;*���J�[\���s�Q��4�ޤ�Y���̎�(�6��r"{z�K�VCJD,D��ԣVB� :������Է��A�`*��������\�X��������wq<]&c�ޥ�D�R�w�Vi�t�#������u*~\<dt�V��k��Bk{�-��U��3n�t��Uq��K	U��9Վ��^֗u�LԶ��*N��+�g{�.�I:�SW��N�B���%�ļe�$ȿ��R������L׷n��&��bf�FfI���l������� $�[�.hn�˾M������M���e�W\j�F�*��:��Ȕ�&iQ������ڼ�s7�}{ӟ�|�����������OUY��ٔ��ut鰧�[;�IW2乑0��Io-�iɀ!���d����GKq&Љ��m��ˢx4k���n>�l�RkY����2�l��K6Y�������݉Ē��B${ʗt0������$�I$�I$�I$�I$�I$�I>����P����w���/��~A�z�]�}qC����'q�'ԭ��;�����t	�G����9ԝHG�;��������}G#��~��������>p��4r ���9/�^������DD_����zUQP=������'�?�������o������}�>~��ߎ�}n���/�Y��wݭ|����Y��}Y�\i~�pr�^����#�.� ��7�Q\ջ��\�%���~�K]Ω`�^k��t=q֥cI]��UX�-6�]�v^��ӻ-S������
�m,�}���䭴�ޕ��_׾�<^X<MFY��R�W��G�r�\sMN��bY�*R}պѭ��Jm�vlZ7�I��ј�hV��[u+�$P2*k����_l�ľw1m,�%�<G4`�1�VoFE[���=�axy�u����ٱ�v���Ψ ;�����S�P�Ruh�-n&u��L\!��zn����k���9������؎z���㈧�|Z�eמ͵�����	���~�gW+�r޺͘��R��P����S�ZެYh��'�ʷ'B�z>U ����w��d��ѳ�I�%,�%�)�s����_���:�]wz>�ھ���m������x8�̧���ƠZ<�U�\�̈́�ݝD����2�;�ˣ��^�0��kh��L+�'��9��qe�{q�r2m���H5��NvM�2>�1�Q�)͢��eckg��rC��RǽNx��rcp��U۩g����2'���}������T���P����q̄��k�Q+�,��WF���F,��7;*�Y�r�X򻧭X,?N`Og�����_�Sv�;��O��M��W�q�Bu��E������1��y"[rm� ��Jv?_�ޤajFt]�0yx|�є����n����ٮH��-��xy5]�p�̾8;��+�j�6�I^IY4���(:Y�BJΎ��[���K<���?;�Ů�t��¶�ۢn��{���ӧOFefF�fFwI�m��2����ijA�k���I]��sD]Jf�iQ�/Q��̒�=��h��#�5��٢7� �����Pv���uo�����+�I;�VU���y���4���Ӱ�f��]q��ܮ��g�A�os��(���&3[w�:5&��V6�X�+������P���=&%�d�M�/`~�������`���Z��m&E�l�\��>g���Tt��"�Y�K�g{8�l��M��i-hM7�p���p9"4�ٓ1>��Tb�T�P��U�`g�b����iTX0C8sA�7	A��|�E�P��������өM6Z�U�W�WJ�|�3�0��>
*�?�pr������m�yQV���@���.��!V��7�ic�^_6Ӹ��:e�*��aS�9��KmT��2�u�*���'f��G�0�
<z��@D��e��Z�c�sn��6�t��o�5��C��2ϼ|������,���r�z�3wC�۹�-I%�R�d�*��h��8���7�b�u�28�[��\��r#�v��u�j�@r��ͰΜ�S�f�r�lQ�����h��4�5sBp
�3����{�9OmP���U���7ׯZ��ds/���9Gv�
���u��lTT0��o����Ρ�����
�Wb�w�ݖ�ow�jN������3h�u5�O�Ӷ��2�,�\q�.�V�F���=�6����g֯��ȝУkt�	���(��3���lZ�{��Yƾ�&��I�����9W����Xյ�.#��fn�y>#�/YLorB�S镘���|-�yI�x�iyj-�Y�VS�i�C+O&XKbA�7.�����K�
��8H�5�Qq���g[$u�癷�N�3��:A�s+4:�ii_:r�:̥��]�po����F)�yB�yf]\���weL�O��@��lR��{��> �v^���n
^ntF}��L��=��^X���P��zPK��}ݢ��NU��e���y����s��u�J��r7o��M��X��,� �g�=�r�O��3W<6c?u~��Iл�Rw�p��̼���)�u��M%ZF�5T�Q��\eAo�Xg�R���[N��Ӥs���'�;)`����޴<�=9�g�M�X�C}��+�@ܭ7�~;8 ��2��R2��+M���p5tJ�}����5ԫ 3��#���!�0u�VKW
�wfJ�޻c���仑cN(��1�/�����EfĿU��Ѯ�;6�m�s�M�!��sq�J���v�o���N�Ş��%jp;��,�B�.��:��<�Ǽ��a{�I41 �j����L$(S�d�֮�:��f����e�pĖh��]��2N4ܫV]�A|�'�J9:Y���/t�gg��v��j`���n�;������E�#�瑽�9_)�0�=�(����yз}��}���W�~mO^�ς��X���2�
t�[��7(�ޜp��l��d�4)�\ v=ַ������ݏ����
�2lP[œ��b�:��+:�k5g�lB��
���8l�+�[��[��:	X���ϻ�۾�Xh�l�ò隵��foAq��ޠ��̨���p	�qI�ҝreQ8��r���sQ��<�:v*.�3j���ݫ,jĆ�d��T�����0�+z-}Y��d��Z�����Ӵ��i�K�8fB""�P��M3�l�X<���ݧ�-T���������̰:�Ӈ�w�ݨE��<p���ۋ���3��/���u�2����'�b�e��gj�rΘ>��C������Y*�����3J�`��l�{�%@�VR$ʛ׷��M�):�"hon$���#r��:ub��l:��
�yB�㯷��1��hbuպ��}�S;>�dU�j[!P�"�H 	G,��$�s.I;`�ܱ^��-H4��*̾�sp�n��8>����)z<صd!
+�fKP�8-*י=��]��@JsͰBA�֛C���[P�:i�F<�K�߮i��z�8��/��ɽ���Uf�G�G�6V�@�k�+ɢl�����S{vh�,5�!m�_HԎ�i<�饹*�'Q���z�<�taoCz�>�Xo��z�>�a�#�=�ayMW�$�O+�~��}7u+�nDa��c]IR�,�jZne!Z���"���w�*3�)/Q�S�� �M��x��^iV���f�h��R��w����J��t��ue�\���D���i8
Bn���gOWBn��H`���7���"�m����L9��(i�c����ؽ��j��]ץ�y����j{rIn��[�X't��X8��M�:�P��clmnZF���Mnᗵ��n�FO�����Ʋn>�C�zys=U^�rL7܎�^f������ķ_}�����oi�X��|�����|$��;4��'N S�f��%K��Ѫ�z͑�I��'%a�+Mև�S��qhOD�g�Kvqo��(ּlfɽZ���@�#�Ĵ��u��
�@�'qM�����Y��X7 ������;
I��x�Q\�NS��nE��%^��T�=��^t3R���.&/X���wH����ƫ3.�X�tw���ྈ���q�*zIB�8��f�zN�&)_�������Wg����ͫw ���TF���(���>�t�[�ˠ�x�"�7�z���_�ڻ�t���
l�S��yq��/��ZS����%�`
^Ụ���.��'Y���eqj���R6kv ��U�o�'�6{}�]j�%��=��;��ާ�}3�x�x!���88�Z%5p3#�S��,f�T����,娺& ���_o:lms�:%�5�۹v۩��[[4U�o�C(ҬN���P鈻�����)n���0h��8gt+)�+��W�@��%�2�s�����DY[�q�]�c�t)��T��ׇ҄6��J�ʗ��2��(��	���e����#{u�m8�l�Ᾱ��uN�ý����7�mrjT�j��pT�+'���tf!�N��Yb�R��7p�g-�(���3�%0N_ݠ�ލ�U��s�Z.р��ЦW\ԙH';l�ޅ����7�
B;'����z��O��Y���{�G����yeI-w�4��fƷî+��$�B�p�`����!����
�U{�e�!�!��&l�����	 %�V+��w4;�X���[B�/�+�Ǆ�B�hhT6m���61��'Fu�0�}&nv�CJ7ٳ�R?f�8篡8O�6��7���$�A$�3�>����_K�[��X�3�u>w�'�u�[��<X������vwi��%5v�qTA�ۺ7���^���=�\�%N�|���M�D��:�7���3i�U�3
�t�����;�b9t�¶���Ǐ^��%_iWkT莌�>��dt�I1�j��53+M1HU�-�n�s8&QC�f¯�*�u�ۍ*�����÷5r]��95;�t����T*��:��02Y��%�	i`7A�וN��f��|G�6�a��7��i�+}�q��f�ɻ��`��i(I�=ݲ��S<vw�I��t�؊�8V�-qM-,�\.�Ra*�l����ϲ��^ذI�&����Áhgs( �[�+���X��WK°۱t�j*�5Њ�V�	�A�
ͶMKOe����t�8�O\�y@m�;p�-��1[��m��ЭSl-Z������k�2�s+�'l}A��ӑ�8	β1k�������V�b�����r��c�ޣ�x��9A��OM�'A�li8�W���Q/�N��ɡ{4"�.�	���zr��bt�S5%��B����+��K��8�4�1�,ÕkTC�B������/6���䓠o�� g]`�A�N����r�uZ�*䲱1v^m�ˡ�yĉ�L���7s�/�Z�����Z�X|#��2o�ΪW�]+eV"�H����U�y��YVoة.����N$�vx�۷nr����[K���efT�l݄������h�>-�^�^]Wb����w6�p)���B+�\����Ոl|v<�1%;T9������H�iX��jA�����VS��δmޘq^n�˲w��5P�)��̡\{�
B�pgxz����q>����"���+rv�Τ�o�/�|��hˠ�xi���A�Rwc{���Qm7ulŅN�fʸˬEC�mn��1o<���Jʼ�u8^�y�(�@�N�����X����_!L��խ���q�5���Y��]��j,P�O6�2�U��0�!;Xk]Ft�"�gʴfCε�~�Wm���ֺK�fEk�wfo)+��!�.��<eR�,>���h��3HS²$yYL�k�^$���uĖn��\^t�At�c��EN���0�=�(���o��n?���g��yl^��}����֒o/�ީOy6gQsw����%�&��b.HU��wG5Hnz+�֟8zs�ע��_��򗹹��s��������i��Q;����a���1,߰@�����E-/��H!��^�|�LI��G0_P�f�z9�A��ޜ層R�������N�3fnn�̾/�H�ֆ�\Bn)��P[/���۫��V�m��j����J��fp���/*�&q�����yr\�Z���͸�>((
��Î�Y�͌f�p��,m�m��x���$s�g���^���|��dD�.o����ǧ#����V�8��='1CG��.��|d���+IF���w.wI�0��1�'K۴�3�۫x��McҠ�2v;4J���˼w]hb�Wc3HO:ē��êM>�%��~��F�%����Z�m��b��t�/rrʵ8o��O�Bͱ�=�0���WEA+����Kތ��%�󷅻{���=�P=�]86�N���U�[�z�T���"N�֤l'�|�Zy���!���:�9�i4�d��v�bo����6�������TvV�2�]� w�:�|3+2ݒk��0�L���'WÍw��ιQv٫�(ׯ�l���)c�+m���k�;�vK5�T�4�qzӶh����IՖ�i<���uq����F���u3`�iW������a:'�sI������=|_��S�@Z�Ն�˺h���S�؞�(�ZV�WO���C7�U���6�w��E+�Pi,���?\>�is��w�;�ν ��B�=��y/����uh�$ ��{�i�N�M�;^��Lm��40�jAf;��7�n �1JU�(f%�~e�-_
I����b�,�!cJ�5t>�ߦm$�<$�E� G�vyo��GN����~�����w��DG^�X�P�8i��aoP�΃u�Z�[w	��n�]���n|8�`���S����5�������3 ^��rS�[+��Њ��$�sۤ��>�Ƽ�k�����ً�Ϥ�*[|L��_�F#�����x��g���*��Gh�cO��ؚ��W�#P��+g]��&�f�I�2�"� �ef��b��� �(jͺ]A:�B�V=�2�E<V5(5��R����e��RIVVQ�f�E�n��z�W������s��8��e�y�Ԥ�5�P"�+�X� ���]8Рx;���0"��vH�Z2c�Τ�Nh-��Ig��d|��	.e��?s_6y9O�ꂸ;S��-��3�,�Wb�������x���C;Ñ�Wy{���5\�!����j#�3�f|�9��\XTk)ǂwٚ�W7V1nQ�M8H��Y�U�B�{�m��+�\��j��S�&`��+.e�X�8$=7���Po2n�c]J�s	�W�H$Z)��b��7�c0�2NT��2wh݄&�m^�`�X����d�}�s`���b�g���sͲB��I�W��z�J�x��4)�1DwNZ>��}5ʹM�.�v���Ⱦou W7�7��u��M�&�KH�Wћcn��[�lhۧl������ �{���a������������O��o��O�����o��~�����~?�O������{�}����G~}>!���<8�`�I��$I�G�HH4�#%��%�fE$�$�r���#�J4�n)z�b�ih�8j�N��O�Ȁ�$��.F" �(OƄ�-��G�����5�d�δ/ݓ*��Vx��(�7|���\=��Lr#�+�g�Z>h�\u���`x=����2��ok�N}��S�]�̀���#��V�����cT��B&�XwV��t���"r|���S.�i�,�m�=��nJ*���������b˃w�W�Y�e#�[��0�׳�9b�k��kHaT�q���ըR�����Ϥ�j�]��<����gm��Zb؅-Gͦ�q�t�v���3�5C+9Ļ�X�������w*i�d>9wd`8S��}�@+�2���i2����>�dl6Ѷ(�o�����U�;��T�"a٭�\�d{z��G���v��s&q
�b�76E�3��X8���꜋��?��$=��9�&}
�^(�1:���M�yY�a��;4tR��6���������	��	JN���l�^�,!Q:<��<8����u����v��ZR�^������c{��og.�u���VV���������f�'�/
��/����3g��a���꾢/h^����i7Y�2��=bQ��|�]3�s���;�&=�f��	" ]nռ]�ts��q6X^�:����u�ۣOV"ړ�����m��z�R��p����B�v�{�޹.��[�..Z����t#���`�N.�Q�`@�-��Ȝ��!4TFџ���`�H��l2�(���(F�B�|��h��L�`�7r8Y!�͈��!?و�\���E(ل�'�8�, p"Xa)"�1	jR!A�&%� A%���E�H2�e�)�Tщ��q�A�!8ğ��B#$�~�7#�4KE��&B�%C-sc�u�u讣LkE:t�D4Q2TD��T�S�i�.F>�(b
��(�"650�uh�76
B&��Z�`��c�b"����Q�E�e�UDw�UL�3��Ţ�4h��4Q՚g���E�:�4U&��kT��Q�`�`��**��\���ւ���h��bna�6jyV��Y��Æ�(bt���-cgM5�rp���b�b�J�-�6�\(�TDEIU�tꨚ�*+���	щ��qLG-[f���傪"))����ڊ��"�MRwc�A1Z56�b*�lm��j�)��ۨ�Q1u[QE�qUAQZ�DKWQ���M�[��%A�mb����sb5��*�e�STQAm�"�*9��!�+Y�4�"�����.nsQQSEUMS�V΢���Ɗ�E�A�E1TU�/7w.�h�kVsST��j}!���i�i[d����D�RB��ү�����塖��N��F�˱��E��.@A��y] '��ϡ��ʂy�\�9eo��@e+8�3��]%���5m"�e��E��E�\�##`ġl�ʒ@b���l�S`�!����];��Q\�)����d�%�[�<�}�י;���������>Ϸ�/~�E��A�l�e�2�E�z1���q��y�� k�r�>�d�g�l}ʸ�>���,�3�>͕6Gn�q�"�G 6�@6����u��N��n6=��?Tl��V��^V���+�������9���?~��)h3;�u��~�/zz��?���T�T�����k��C߇SW��N�:^yO��S��f3>�%�[��;{���fFv^Y�+#wL5>iy�M���]�{�/��P�8���ee��9TU]�]��=��~�8���Nݓ�{��}���w|�TۡM]m%w�]I�J���;�Rj�S�����=F����p��5�:�gk�v�d�f�9S�h��X,�	�a��h�~'���n��σ��a��;�`�eA�[Wv�{�uֵ*�f×���6t�ҬM�1�AV&�c��H��I��R?���%=��M�y�N�`b¸
>4�:�ԗ���4_����Y�Y��> �����j�˷K4��)�4�q����O��R�-o
�����1�c��٥1e�Z���3�Rk�~��i�\�On���>[���+Z��V���>����/�ݎ�Ww�L���{W�B͏T]�s�Y=�֛;�l.:�a��7|(���$�\�NK�q�������`'غ^���r���d�j�Y�垬5�C=������}��F,��n���8=7�.�b0�{�ډ�5��ʍ$m����{�'c��Ȩs�y���)��>�1�S����� t���L@��r�z�w�>�&��[q�{����G�}]�ۄ.�n�	^쮬�W�����ǫ��|Ƹ�w��䝷:�b�gH�g��-�Z6��c��>���<).B�h.�U����&��x�;�d���M��m��5ә�*\���z[�cp�$�5��h�F�5��3g�����=#�ݳ�]�dP��X��]���_�a�uۺg�6+R��BV�u��������T�ٮ��Mp����.�)! Þ�t�=�E��Rݡ�N�{���6�{�q�{�ث����:�>��*�SB��8���KDp[b���R��MO#�,�[Z��݇���/zaBD(��R���bW��Hs���t>/�S�(Ή��q�|톉v\k����zٹ�E�#�# ��W��5�n��/}���r��6Y���|������9u�����8+��_��j��������up���8����в�̭�-�YK�O��
^�����MM�]�������my!��RuY�۝��^׎3V}�4~���;+�����?[Qί=N3���z ��w��]���7�)�5Z��6�1aS��ɔ�ߵ�NT�Nb����O��t�<5!�i˘丨�y�{����-*��N�}uGA��i�z����67�VG%?�{gޭ�/��__"m
�_�9#���M^���6>��eJ�W��S]n����y=�/�TCe;%��N�~z�ڥ���2�������]X��Wr�ޙZ���䤨����>�F9����y�lj�FW�J
��L�w��٩ߌ7��.G�0��r�
��eHp�oG�~����ɢ�����x����4H4Od�e�ߗ�l���f��j��pToC�*فb$M��*�n�2�a������u,���_.���sox�]��f�|����Bu{x��F:I�i�}f�g�b�'�����x�=�ݷ�H{��<�=���̀v�vR������oB�5E箥�{/���r��6�� Џ]���on�'q�ė�LxQ�L�}�t��M͊2�OoSU�N6OV����}M��[6	ὼCl�zIY��]���H���Enzތ��4p���u$t����+g�wI�5z	��5f׭M�^OZI����͗ӯ��a�m�`�Ӫ�к�����n>W��c;���9��_�5�W����ȼ`�>�Z��⫝̸���vĜk�w�!�.�1��cw��duP͖�\��p%^�p�I���(�u<��>�1/x?-�����y�{H��yT���f��*r���~�z�r�������-Fk��6�����j>���vM���{<|�;����A� ��?
^]N �K�*ˣ�X�_��W�T��mu�뉑������י�q�g:V������8?���[}��V�*�;��r^��lJ�|᱌\�UZ��+��%��F���G�j�H���f���q�)5�8Gyt�4���a3R?�	<�H(*��ƕ�����罿I*[��P�C�JRX�xq����i���{�*�Ы���C�>�rǻB����*�=��|@]!�8arG3����yT���Uw�nh��Wg���������q�߆�kJC잿�W�����+�t�h�<2���ӛ6>ꂶ���[�f�C*�|[o�jz��d���e��=zA�F���ӛqQ/Ƒ��5�w3���q�zr��(O՝��!�5���Ϩ�4 ��m�nW�Agj�^�oQ5/x�A���+i���Zv[H=M�z�<p��<��:ݕ�ݤ��G�2��܌�s>�h<H��p1���6	#�]B�^K����gd��Z�x}�xխf�}��ԅeAl/{`|5��A4�D��OL�x��R��<@6~����{����{�R�0�k�ExP�Z=�1�O�^{��#�T�C��*��Z�Ό���h����F�֒�6;���F��-�q�t���#2wr�
�W;/�2�R�荬P{�ζi6_q,iԙu+���ٲ���}U>ʐ�縦%8Ps�y��ֽ��z�m�:6gJn�9�2�ΠΨ��.H��hv�gbz��{��K�v70F��^�Dں��{�F������C��w�gCT���'��w�V�T}z��F:�Z/�؍/7�ݝ���i�L8^@3�:�':��Qbl�>'}/O�Z�����}Ă�-���;�I�s��Y���1�ˑY�i����7"��z�wK��{=G�A%�s!o���>G��VK��<>����5
�i��h<�g��v����SF���*�^�ڌ�柫�`/i��Q����F&q�����yo��H�n7��u��s�Ql���=^
g�Y:=:_{����������{��DH��8߬������箦h�����u&��lp�;l|GF��Mz&6@����F�MN��E{锲����s�b#z�����X����$��{��r�x�|���������;�@��M��=�u�����-�<-4�W��tk^�yIzO{�u����!�%��_�g���,~'�_w�[1�Z��ۥqY�x��I>���vU�LM���pVt&�\�U�����4���Qݝ*
���`�p\���אǊ�Yk��)s.+K�w<���~��Q��Ϯ(����o��_��mA:��R����׳���+�5�h�H�%͙�۹�n��xpc��9����F�XD�2k���-���d�m�W��H$���{ 5ә�8Q؇$�ӽý�ߔ�&#]��W����\���>�}=�l���gꓡ��DsZg=��{�A<��%�9 ���h���5|Zqא��_�>~[�Mz}?f��㾍��rR�-|��}�yڦj��=�t��~{��r�'�_a�����ɖ�G�z��|��I�U�y�8?*�an�l��*�r��v�FN8��(/��ݪ�h�y]�Rۤ�5)�s~�c���������l����#��{�x�'���T�Zϟʝ�J��l�l�l:-��I�k�BxFܞ���]=��)�Rc��/�ջ���*C<,x)�ұ��׽(ޕ�1�{}�^�r�oȑ~9���a� �|C�"��"�199�8����y��j��F뚆��DF�[��N]M���Q�p�7!X.���Nͥ�*���*5Mva՝�S7���ȀJ�����S&H��L/>�ۇ�S�z�r�N�I�T�<���Q�˙T伨��w��Qg���Y�#�����]N����z�d�+ѷ��7\
����x��dO`�f^���h�oQ�o+�_��lw]׉�F��S�/#$� ��#���w���q��5syC9X;�ڮ��;���P�KH���O'������4�"�~���~�W[���"�t�z�}�w7~���A?i�X��Q^��Q7�N��W����\vϵ��I5�&K�*�f�Ϫ��Z2�������Fr��x�/�dA�-�@Zv��4��&O$� �w��2���� Ro��~�7���ʕ�@��������>ޓdq�26r���O��z�{���<�.���
ͧ�{(��/�M��������g�}Dq�m�
�>�������_�>�b.����_�ȉM��3�0������������f�e7�cCP�����V�
��Q��'�&��J����=S�E�:Xçh�A�n�z5Q��es�͕i�в-�/�]�%plup���ת�U���i�R�jafץ�O��>z�=�w9T~Ӌ,6��>�O��u�bw��Ld��p��@����r���,9�\EI(TH��ξ�^�׺W��=؟�,�"�]yߜ�d��og�{|��.�{����= ��X}�n,y���?��`&�#�ٗ���}wޚ�z�Eu2��d�hӓ�E��{��������l:.��w�4�������[������G!���7�{jJ�jL{H)��Mj�p�j��zɦ5A�l3�Y��[_g_��龝�*��h��2����?{���̿ق����CÞ�O� Y����)��=^��z����������4��lH$�<��(�ا��ޱ�Esn����֬R�C���������J���g��O��{����!.{&LF�k���݌g�w5dQ��ˇ�Iھ ќ��ފ��ޭ�&�>N/g[Y��o�W}�b�*��v4F�h9D�Ll��9@&|(�.z���,�a��9�͕y[9�L��v�񏍯=W�[��l�(�2���<�<�p+"�'�t�=�	���kodμӎ�Bc�)|�ܟGa�f��n+`��Cr�.qp=��7{M��ǒ*Y�P�;|����zP7�������6{*�n��wB���69��Ef�#�4�2�"�	+x@�;-�M�y�����~>�u�;�D;u���q�*_ކ���~����~]G�d�Ux����̻��c"��5�=`j����f�x�2�vy������#�kD�Z^���٧�?�(�4�<lk�O�s�f|����W��.|�ĭ�y��R�߶<�0L2k���Y�듺	�/�a�5i��F�W���k�N��>=n��{�K�Y6�Nݩ=3��>)MU岸g���ww���]�>�w��0>��������5����	�~�3Ey�.����K�����e���a�Y��z<�=��U���=�UŽۚٷu����/&t{R���d�j>�Ƅ�t�Xu�ϗ��r��x;85�x���]����b{ᒌ�ѓ2����\�yb�T
�?��G�{}=?O���?g������||||{zzzg���{� ʻ��L��|�Z��F]�v�F��ڕw|��y{��P�z��˥ztc�{���g�*�0f5rt쀍������w��9�u�U��J���\��a���xݠ��6*�of.{%m����+��*��ĺ��rN���n���X%bt�Ɏ�!k1����1���\���|��"��siа��wL�ek���
I��=Hj6�}��e�m�&*=�i&�v�k�n]n� %ɺY�i۫�G����^i�6�i���V��� ����ܭ�)�i������K�חi�@Ә�T�P�wpi��.�c��׫fB�Tm]��6��ɛ��i��Zy��u��rb��x��n+���E��R�c��"3hSw}Ռ�����҃�:���`[G�{a�N���'v��*pU5&7�J��l��7b��ze��l$[`�p�ذ �z	�>��5�|6rhL[��Ǹdd9�͔��ڲ�y�-��Dǽ����G���U��n43{tK�����)�V�;��� i�,m��b�'����oWINj̹C� �)A��b�-�".�'�6����F�R������C�?Ĝ����Os�6z��{�d�cWn�E3|o���`�-�#��јR�g9 6z����AH��oEt��u����w���0JF6/��r�,���7ch@���,�J�u%s��仺G��c���b��:*�'�3��;�s�cM+rd�ڀ�KtV����8V琪y�f7����sk������1�Ƽ���~�.j�)�;���Ƨ����w�-����L�-%V��G]�4\��N"��79���ۺ��FH֑[}Ϙݗ|��X N���L#��ҁ	v��mj��ӫ8���_I��A��;09w|?ɷ�z�L�����)�Ç�-Ԗ�{k�x�~��r�JMx�c�Z��+ Yއ�u������^�S��f\[���h�U�V�dP�ד)����鄣�T�&<FBzOM�}��c[q�t۪��E���7�:���ã/;����k��[G �������T��t��(���<g!��t6�^yxN����y�����Ez<��x�t��>Qg����i�t��{���B��n��7�����`�&�<Sp��dv�����2��jʾ��Xa13��N[n�$:I�SI�3^5��A�}y����n�b��9�Li�ࣼC��;�0�L��+Grmk�ٚ���3#|4.���iF�L���,���X׍��cv�L�V��.�Jy;.�ǟ4�b��F&�Xy�$r�3���O��}Q�,K��35|�#$x�ˋ�Z��谉ۈe��v��Z��^���[��r�I�[�Ë��㬣�������l�m�~{��ܙ���439��.b���C եn쭹��T�mi�����!�\z�:���B�f�R�a��1N�vr�
��{p��۟g����F5�4b���U5I4m��5�Z�U4�EQ$�Pm��*��a�-�1�b����5y�TDIQ1<����ڢ���TASW'AUs�8l�&1:a�(�
+lI1�b&��g������5S�Tlk�tTT��FJ���i��*)*�uQf*JM�:��c�͚����Gww��:�(�뛚�j"������(��ZpMcjcmh�SM3�H�j���Q�4DPQ�l�բ��r�;�WFCv\�PUQDr�U�Ξ����f65U�EGh�� �,F���7(�+���m�7#�\�A�kf\[�5��b�h�b��F�1[f
�7�p�"=t�1A�ƹ����ָ;QV��EG|�r�5�X.O[�bzc1�8p�sd�\�*��-Q��F��b5�9��sf�XƩ3��X�<�u�sm��F���Y��`Ɲ��q�j��cz�9]G.PI�b	(/Ā[����u�a�ȥ�\Y�-���q"@t^�5Ů�Φ�=}[W��K��8.I���/T��˧�Ǹ��zق������{}�ڰ��1�q���	��skCrC���	�`�z���K��t�V8Q����v�ӂ��f�wOח[���od,kb1퐇�\������uCsf�i����WAP]�轛N�a݅-ޟGzń���-�g�Ԁ�= 0�|�p<yK��T�9U�˒�m�1o �-�`:���j�櫔5Ty��*/���M�����1z/M�$�!e�|�v����0��ȧ����>:.�[��&�����?�ޝH�?t����d���e#�~�~3�t���!����?6=�v���εuv;�reQ�9�O;]�LZ�^Q�$�ȿ��(JSW��Ưs� ����A��Ip���k�bc/�Ou�����93�=�<��]'c�NO�H�4J�[ ���k{�\:��mb�2aէټ��}Un8�Q�Y��c#�]��/���O���O��T�*[�Q��XsQ1���TQ��nC��m����z�n�i��,}R�a� ���L! �7Od���0�v�ft9/I�2�K�=я ["J3Zm�2�B�@�\?c�
C��r9Ĉؖ\�:�i��3�wy��0�������M�������Ɲe���Y5S�&��w.��_%sɗ��.�n}�+��iH[3�+���ӕ�]���P�z�܍�y�ɪg���-.Ny������nԩ�E@ Ծ�� %����Z̆�L	���~��!�M��9�xo�DKl��s��q�K�ՅC�t �܀����P�?P<��&E1��z8��u���m�n�Dc�1����ԥ럘�HJ��1����ipW�4ux���{�w��.���Τq<���h_Xe7�Qx�X�	���������:�G�2
и��.�[ɏCC�=+���N��- 0
{����=���4�a���%�� v���C˅�(yXK��"�f�F��y]����)h�����!F��H�Pny��Dש����C Z�Ż�\��J)��F�Nn�nͅEз�x�}���88e��|S_|�|쁔���Uר�C�w�>e>�V��R�=�&[C!�e�m���{������#V0y��XA�G�-�~��Sβ�C]��hg6�}�&�8Za�U�5y#:�^͜eY��Ϻ�"1�`|��P��l��l�����dEBfg���q��^A=Z�,h$k��;�T\9�\gAG����D:0�N�T�ʚ[�0k�"\j��� ��桓��D �^ъN��JĪM�M@+�iz.7���L��p��&(-��A�5N�U���^�����I�����-��4Yq{[��=b��N�`�p��l��i�]�������N�%Ք�EܻS��a�WVjV�P4v=�/�v�H}8�v�[W�%�4�Nc/�)ʔ��m�At��%X�p��������&O����S�M���(I���>���_zc����.������sWD&Iؼ'<��j�RN-�{M��cm`ncN��Q�<;6m[F-��l�z�#ا�0v!��˷�^��HޥI�y��?����Y��걍P�
����de���Ŧ��3������Ez�*�����0�o�)B]k�~�z�5�[��\4;�kk�	�em��3l��c���4�O>�ߊ�? ���U��r��q�Z!~۝Y��w���3I�Qo
�S���P9r�Մ����;P�Sû4nC�ˇ��`鹽9�S��S���r��'�L�-͌;oHk2�o%�uH�Nd㋰J�t���֑<���Ɛ@^�A�Q>�wf���cups�Tu�|����(OH���"�:��:�~������U�0j�X=�y��<nKDh���P�u֬;����g�`���s�-��,9�aJ��'�u^>����~�R��ҷ�ҳ��!�~�c5W+zA�0C��o�9.�:���t��-�иw.�c>���1v����N)���{� ���g�9�+�j�?�1'�<�<���ȿ���������dIm��g3����$D�<���r+���i�������a�׋���V�5.%��v^�[�^~�wBs4���,�v�ݠ��{�ߴnT슃D�mLі�#��\�U8���

^�Tq}�2љ��ffUT�t9c���i��wl�����ٟ��ήO\�}m���C��H$=�a�<tE��WK�ı����4>B1�vI�>�}Kh��w~�NX���
j-=����Z�&c�yk� �x���F��q����p�gomЊ2��=��)�-�;��m.e�s��cW_��[�q����aT-]
/�J��G��~K�D̮tx�����{��"s�G�Y_p`|p�k��#�a��ڨ@�C�����L�ҡI���X��O'�xE�!�vw_iᥩ��OM�?���S!"��C_w��b�S����6)>4U>VM#n�����~@j��pZ�R�v��V������k׭��$8��� �^�'�ƀC{	+Z�t,������|�]3��D�X<Li%I�k�8ǻ�OC_Z���.p'+w��X����4�'h���%���K��EL-�]`�LV��T>�b����
���~ũzی�rIjR��O]�e��U��
��U0ТvT8�jv]�O̓���+�C�XN%���3=6p��G-�Ij�A�#�1i���5;4]_�����NP��2�Gs����;����bz��iG�Y:.
�x9V�׽G�	��x���C&�7H3q��|b�����a����ہ3]�e'�'a[�� ����$�7�8$���/{yn��2Cj���]�g���9L]��T���{}M���(a*�ǝ�;������w�Cq�ݚȶ����>�Vty�-~�;4ڬuQk`�J��+���p*yص�;8��b�M��~����=w	����~�+�0�/~�mt��}Ǳ��l�׍���&O1�rn7ucL�bY̽�T�u����Q����+yhp�	��(; ��U�82m\4B����ĳ+;fZ5<�%��}fQ~���!�������b�AݎtK�z|�CxV�e9;s�5nkf2%� D��p,	��~X	��6q�6 y���8�'��i�[�v"���[m�����^*�k��l�--:ɵ�C�qz��ǳ��9�73M�,t�9Iw�rJsP��0it����vN��}jZ��Ň��y�cǔ�r����fq�.J�������v��m�<���#����p���CZ,e-�_��d�zxR��	l��
v��ݞ��c6ك"y�g�8k��C�Ji<#�I�ױ�X�^��x�
7�E�l{� �k<qk�4����7_}�P�c$��A8��d^�Q���ĥI����lj����[��01������iѓ�ƋE���F>�ø�ɋ���r����iª�7@�)kZh�j���33E�K)��*��N�T�̸F��/U^M��t�a�N��k�拷R�>[�:.�n�E&[}{��'��|�nͳ/���0��=Y�c�U�w�~�L��#��}�N���bS��S	*Fͽ�Ɩ;k���l���?�w}������|��f�~0��1����v
������%�Qv���h-�Ø��k.M�U��vwS9N��o>&l �z-��p���n�^��/`���?���=7J�d��A�y�c{�y��C���(��at!��|�Ƽ9�?k��M7X�U����1U�QL_$���e:�腒��	�\��~>;�/�[��q����`?��5s���Ȯɻ�vnܧ��}�}�pAb��[ZP���M�����z����H�����x.!��]� ݶ&���w�i5}��e=��x�r�x�j�Jo��잖�
� �W5���#�C�s�`1\���,���Ι��y����P鰸'a���M�2��|��0�H���瘶�r�n���|�OV݋��y�+�Xw����������؝������8s�I0�meذ4��U��3��koo�Z��"��j����`�7��tZ�����g)w��@��L�~O�i'�1|��ݝd�aa���|Z����!>��]��ʟ՝�Œ����?[���R��{���6Q�R#Ex��%*���`)��f;��E��w�4�K��۷��T3��۔�A����f���e�4�񽹇�뫞��-���ＲrlԂ��^nꋑ��"6��T�����.�f�C$a�m��={��N�kdS����A��V~��W?W/�SIa��Q����1�]��-k%��8�P�*��Б�g��0�C�e|�ĨX�����G�����%o.�إ����XʊƯ.��_����j�Hͳ��{k���8fߵ�d�X�FZ�y�]��f@�) �Jq��هp��|�&��^�B��#�^%B�ʤ��`�Ԑ|9��鷨�o*���~osD��&�
Y����m�v�_Jnj��&I��[�)̈́�o&�����&�-e��ڝ����j2q��E�*���zA�" �D9�n]�5����7�Rdޞ���\�אs��뎋��ۉ����I�lA�*�%���������uǇ(;#|�ɽ�/�haf|�0Iժ]�; ��y�'�S"�s�c��1�\��~oy��6h|�Tx��S9��|g�3�%ȨF\��hR�0�aT,��9P��y) ��ڀO�û4{r|��T�
��URCF�S�Z@���$�'7�7B���N8�T�� ��4�u��n�p����p��¼�z*�.ʃ�����vZ��z�B	�k�̐W'j��/�z���)ks��j�F�;���Mzli�/7��v��_[CLô�p���T����stW&�잋rs��{�x�P���Jp��
-��k��k�+d�nV,9������x{��oE��I(ME��<�>`��� (�5=#�kݦ��u+\rn����=2U�����w����6�@T�|-XK�`�<�W����ag��Z?od���χ$�5��&�|�;r�WE���x�p����Զ_��tO^/a�'�D��y��h����\ȏ�/�wBx�����ۮ]���5YD�LR,D�e��虗i��Ž^��^}�.�^�]��x!��Oc>�K0���O�b�[o$��@��!�zA/�j�Pi�z-��������(`����In�۲��c<�p��q��[c[_�cZo! ��/���
�W#^k}�M�1p�n��MWK��3g
5�5�5n�ЂXGE����=��Ʈ���ƣ�B籆`WB��G\;ztg����Ŝu��T�a��6)���c_�	���q�ޟ-�N2Y�R���Bl���7��#~����ֿ+[����c[]&$�	�=���'C�L���<C�S�a�I-��$\�}�1��/7D���NX&"T.�g1�}Ǆ�-���Н �S'�7���÷;��}L��=�}�靍b�k�W@�iw_6�mrի�K�yH���{���b����8Ȥg�����{;A~^����/|-��'�����h��*����k4��_)�")m�9�*�}9X��m���V�ڬo|��>�'��|<�;9�F�+�.�8g �y^���^s��x�))L8>��o]<'�}iٱ��#Ht�\&���5���9S�-aX�r�8�'���]��0�.���5(�������ڢA�n�~�~̞�q�q�dŦ�1�0wa�$�q=jv]x�Z~d��+�C���l0����~��;��ݝh[�@O@{����kLp�n�N�'W&m�P�r�߉Te�,��4�w�f�nz!�B�9k`�d��p���8,�zp������@k�zvi�X����	V��;{x�����F��e��Zc��t��q�>7rʹ9���s	��������Ǝぢ���.��:]]�%�i��n������N��y�ǲY��ɏg��ȉ���r��u�ݒ�s��О�N�f�vپ�_����C�"m?Ohv|k�5?/r�.���U7��K���e�mS{s��נTњObv3_�k���6��4��C��D�^WA?q��]<�F����⧪}g%��D���A	���s��9����9��4�7�X]���=E����h�2�]_��oF�~} w�ȉ��;`>�z2�~��O�[�V�>�^���7��Кi�h�[˧�1Ljَ���:��.���{�A�2�t�W<��rQDo+�Lm�(�/�kj��!T"3�(�����"7�'��yk�C� {�z�iG"r�
������p!���� ����3��ɩ��н�U;.JY������N��a�v�i���a�-�oj�������z��C�S�-��{GUX�	?��[�c�0�%'͎�zFN/��LŐ����1l4��_�U��V��E�>c "��&T�{����5b۽шI�]!
&��tA	�/��IM2�+p0e��݈<��5�<�۸�����x���Z��R�Ivc�� �������~�s���"���T�؈��V���u?Xkr�^���oK)��6= �5�zK6��3��v�R/���ޣI>y�Rr��E�[�Г�������+~�ي�h���yR��w߈xE�H�A�/���9#ry���*]�Y��,z&�u!��rꮚ�T������'����0�W�����Gόk�!L����J<��n���{�f��ˡ��s�</�P�ԽH����$Xׅ��Bsϡ�?�^*!m���W��p�v�x�p��?!="�9�*���2���Z`�Ҩ��Y���n��;��0�����{~?O���~ϧ�������������������Vمh<eX��N�{��3]���;��x�B"�̸�,pY�~[��X)%��PY�]�z�=����s�����2���t�)2�;��G	���WZ4�抡E�n�R�@��ۮ�w����X�4�>�Z����j���������%9����W*�IVl���\ ��dݛ|��:�T{��M�YD���{5-o*TWN�U�O�upm��:��+�D��4tqR^�n���)Մ].�� �֜�2$n�7Ox�Xf�lKNYoy��o,�d#'�Oqk���@L�G����L��J�F64Zˬ��jٹWL>����M&����I��t������K�Yoi�w�+�Ʋf�":���j
V�h���ӏK��1C�)l��
��$���/Qˏx��IJ�^.����yJ=�/ޱV���f)o/���%���&�����MG��ɩ[��	[�q3����[��K������k�7����9E7���1����/��)l��b�[���Y�=��L��n�+�n�Rr<Į�e�`�����KU�o�3��P���Y�4Ƒ���so!L�ƪu&p�b�̶��ٮq�Z=N{N@e�عN��_[�!�*��Ÿ4��]�k����T��j�S[�Y"!�϶fvE\O+dl��E_85׼�}2cp3�X��������}GK�l����@�>���8�)��V�ۮ]��B"�S�)OAy�=(�ie�ȵV�"��V�i�oj���ur*`��O�	z]���ٹ߻�M�9O֥x1O\��a��`����K.��Œ���%|���c����H��sc�ܵ�����=R�4��+FtֹVΠZ��[�׳4.jC'Pn��r�{���q�9w�bx�dv�hN��̕���%����]�U�[��9�wp+'�N�n���fn�O ��nO�n]��{v�Z�l�r����N)��X4z�h��5��^�(��j�����*`�{l'����M�O���H,ںG��6]�D�˻a���C3e_j�¯q�Y�n��v�q�N���z�U����eEܛ�x�=�J��Yz8(�C)�{9&�3m���~,�U��x1-\c�Y��@�%a
�[�Ժ���ǫs_a�h�ul0��]Y1&_k����]-پl7���oÄ3D�ǧl%]�
�%��C;,/Xu[Y(u�M��փ�&B��0��:�x��%A�ii��m����X}Y�b�6��2����2�;�_'QXg�<�&���u��W.��(a�ˊR�)* tؤ�Ŵ�w�8y�@�Й}��{6����26չ�2�kW�m�K"��_��є��sr�m��e�_NCaU�����T	�p@XK2f�AMvKAK��Ӻ������A��n����u�n����g=TX�PJE0MT��*��rS�;��_r��+����Yw���}4�.�Dp�4r�s��D<��;mm�e뜩�k���lQsf
7-���TQ��b�j��bpng�s��1Ѻ�j�ÅuѮF1uǨ�4u�,��n9�^��-�(��ڮ�
��sZ��As:�i(�n�i��5W.Iȋ��p���Ek����D\�A|� 麞F��M4M6���w�PMsr+�AպƎs���35�-�r�3�II�i�I��
"���q��1�Q��njb��-SZj�Z�^s6,j(h��[%k��r�����"���wQ�����9i�C�#���S�L˺܈�I���)������4���E�E%4]]�;����&�(�#l�T:Mk6�T�SMb��H]z�Qܚ6�EA��1T�k[�њփ��"��q%rq4>�\�CEEGV
���WYܭ�*:�]I��F,��j�X(���7v�Q7Y����%Vڨ��9r4:(�F��:N3�s���z�u�\�:��&�$6�jL��w��-��
��~%/Sub�{�2�2j�D��O�VM�3� �}k��0j(����������R%&�h'��5_��H��!$%~D*Bp������� ��~!�Ԩ5�!�y��3w��^��;s�z��hv��Bo�^5�=����5�^/��!ݹ��*��/�W+���s��U���QLǌi6'�;_{L�?pZ��i��
$@��+��6�g��Z����M�l�吵a!���E����b���iJ�&�W�^�4&���voD�F̽�ʢh1���D3�-�M���^h�O�/�������/����m�Pރ������ܿz��1z���ߢ���l�Q�̽J�32˞v�%6�5L�M����y��[$�y�?_�"�n��@Pw��h���c�����C]�v �+Z��A��^�1j*���g�f�2��l�瞝��ت�vA�g;�*�M��<��|�蛑���m���׆}('���F�z1���쨸r�赎��1f�-�1]�1�`x��1:�5�M�&=�2׿#�bR%B�^p��*K��_�/�m'm�?������c |G�<�	���#�_O��̓߃���n�Z��UL��_i{�@�*��]�N0��E4����	<͌�qa���t�C7�5�?/��ͣ�Ze�n���j�1��OUk�X{B��fW<�]�#��a2�m���ju������)ͅ�o�>��=3������{s�[��p�&E��z��%�C��$�<1���G92Y�/?ܦ��q{�z�V.cnpL��=�ЍΊ��r�:��~�  =�;�����f�����	�K�H��?��x���<0��}!�p�'�pG8�7�sn,E�iC@n=��F`��L�l��c�V��z+�ÿ1�`��qz�=
4����:�қ;N���8d�]K�{�J����I�Y����.Qz���4چ>��f��}p/�-U<�fo��B��	د0z���G�d��&(�\��e�qD��,��5~WZ�K݇� �4��dZ��{d/cVv�uֱ���錆�G�D�	�	��]���P��b~s?s���I�!�g"��'�};�8���T �s�w<��g#c�D���-�v�a�XR����ô���gff͹�lg�)����hR����0���d�����0��@sƏ������)���ȟMFfQ}�,�s'"w�E�ǍK7k�&Eߕ{��U�������A�١g�����9V���[�l�r�voS��ȴO@$?�a��zeà	��:�}ћ*�]�����7�)!�� #2W=�E��Xݍk�$<��� �s�g��O�ʺ���������)0��5�@_�����k���VKЙb��\���(��g�:ڭyƪL	��FqWwک����$z;%��2��3�㆏�9����/��$�:J׋�t�a;�??Ir�8);����>���vk�N�� ��5=����v_vӵBnN{�z{��_��=��x <�?^:zsՊ���y�O���������O(&����R�ԹH\�X�2�WB��m��ѽ*6�P�`���u}�j�M���'���K�lk���\m����.کnj�"So���@��oM"&�������w�8߾��L��顂#4Q~����P�y����>�?�7yN��K�NR�&-[)�'��c_	��/:�J�ߣg1�6ہ	��
m	����OP����/u��;��0��&��_��AN�1�d]?��tHǂJ�y_���_��%��<����~�����������t$�g��Ƒ*������t�Q�E�x�+L�wx�r�nn��;cY��f����i�%.�>�h0̘	���S �Oa�D�q<q]/G"��XJ��.ōk�c;]j��Dl_���Z���[���L�zz�f��1Lh�r��*���v��Oswfz�Ц���H:迱�4����k���k@n����6%�o�KS&��^ꋢ.�ឳ3M4��v?�q���z�����'hy���(��~/p�}>U�?k�T��n���egg-��٨nGGN95�YӀ�љw�x$wuo�sv��"�qO�Pwb�u�!E�	��V���V<�S�K;�a����k���'c��Ɓ���^����7�S5u��^ý�a���^�V:����vB	�u0�t�͑[����~�s��;>���EhED��xo <މ��orX�:]��f۬3�ɍ�������uɈ���,Ɓ��K�j�����gk=l���fpәCd#N��n�^���7d3l�J/ş�C�"m�:"ص{�C�oL޶�ަ����<u��pɡ�ۼ����ĩ�x���&�ͬa ����$_n�T�c\�;���ի[�V��7����ʱ���~05g����'���#73z|�^�������S��15�>Ȼ��q�4|�jAK�~T9KL��Y��#�Y�z22�~�>�Q{�:�1���x�=і�\S��Lڸ�h,�`Z���Y���/H�~��с��ǧ��ꨆ}h��9����*�.m¶�^}�Č�ɪҚOŰ�ѕ��5�z�q%�|w�o>�e�ky���A�\��A����k��!��M���0L��";��Ӂ��zT�T+z�GiEOK�d9���*`�=�`���])�v/	��"��IRk`*]���ۚ�J��7�fଵM��\�&9����'Z�~�h���y8��4�㘤�_���f�و�ۤ�l�`�l>ȝi���>��n?���~������[��ά˳<Eg8�Ž���g�w}غ���upa2�.�/w�*�j�̦�sg��g'���ݲ����^-�өs�����+etF8y�7��-+���u���xo�<��������g� �3�9��]���� ��"l?ݶ�sI{��@-o�Æ1f�i���eZ`����2����̤����u ��=�.��&�#��5���S)�B�޺5]q�إ��ܼ��k�b�^(,��e�%�^	��t��v���熣��T7B!U���-g�r�i=����oI��P��I�z���4 ���Г�-2m��ϠU,�@l[�6��`�>֬���H��Lfi=v��0H>c�0�]s�;�����:�è�k,rz=:e�X�eC�r��=p�z��nf��u������ � ( ~>05�~�;�|�C��lA��I86��0�D���7f���{O��T<�>^���U���PT�T����|�c��^zƟ�݀����u�b�mӜgm�_f+���<�˶��K�Bhw�_�KOհD��^�|`h~�I��m��u��������.��w^Ku<30#<��e�I�I�d�� �x˴��*���C`��y�X�u�̃�6�=V�m%y�����ϫoV�-���.��rC$c�f�2��-�<�ӹ�y��I��|���uv�-�ͱ�����r�N�0C�jL�
m��R���J�i�L��g�w C�,����[c?������OB��Ԫ��ŷ�s���J�YHN���D�c[�n��'������"���"˻84�Y������j�F7Xގ��fx����~`<<4 P
R��"P����~()��|+�B9<�|ǦM��~ʊ�o��vA=P%��c9~�����}}��T�z�﹂P>b�9���i�{Κ���b42״b���ĨR15��PFD�M��-���"�0�Y�9�{Qp�1�zE	��(2�p�;`ܗn})��A�$�22ݐN�bZ��s�n־��Խ��P�r�'��;����<k����G�.��;}��	��1wph��vrO��y��[t�/^	@��/��-ᄍ�B1��O��Q�9�%���N�(@�C�	eWƝ�_T��dͲ.�q̳��\�.+�AY�J��P�����ѿe!�0�C�mשy/���k�«�es�P9r��PX�v��gwfN��٪E�4�Ύ����|�|��������*��A�u̜qvJ�t��ַ�����G]��W��l������<c��!���[���Y1��ͺ;M�+�[�Mб�Î����f���ee�_E��~o�O�Ou���r��A��p�_|`a�9��v[]�XsG��L�-Η֙�i�(���]��ۈw+>ي�K�
Ҽ���ed��<��K�b�2�\�}}�Z���6������1��L_WR�Z���-�xT��g,�P#�x4>Άn�Rr�e<�=�{����6�rG{���'��������ϾJ @�T("EH�B}�SG�
�xqzA���ֽ��i�Է5{��*V
��.Ah_�&��ܚ�v��vݭ�0�]���7,YE�bK�0���L˴�lk�[9y��������WiZ�Ӯ :y�5ڻz��vl�7} ��TG#.�tE�>�5�M��~ǅ�n�啜ƺ��O�|<�ω�d�V�x���z���$<�z�/@���r5�o_7wZ�hr����x�?d�O���\:��L�0�S�����5��쪖�\�-~�A�{��rw�	��E^ŨՏUW!��\-�d`��*[_X��8��#�d�fX�Oj�&)��I/4� 8�Lk֕
O܊��ס�V��N�� b�S�!�1~d���vكf��c�\�k�$=�g�:]Қ����V�%9���5IP������𞅾;�alm�!/�lD��8V̚�.���xS�3	�5����1,���b�����\p{���N��X���ۥ�t�d�(d�f�����1���%P����dEL-�]g<SZj�����_�f�~��Wj���[�j\{N(����<��~���g]i��L�,`%n�|�3{����G^~�>t�'�>5d8	�E�@bφ�Ԛ�:7bKZ���4�w���=����>�=E�{xR����Yͣm�[fҰ� _lI6w����6�}�>�*(�
L��
�@@�H�D@��oU���vu����;��`��������	�Ga�D�q&��v�qi��^0(��0��kۦ��iJc��%��t�k���D�������J�==�l�u~��`Z���o;�W�mY]���gf�S�I��q��У�Հ��s� W�U���Ln���q������WT�GS���#'Vkm���OjرBV��
�Z�9/T�+�eu۝��zC��|DqpB�����l3+U_V��{M�,�d;$�-)�W�*��x�|�gӮK`q�vB}C��G�@�5��R����Q�}��{#Ht�f<��|/bv��n�f�m�E��^=$9!�f�b��(�b�]�k��M�������i�ꠝ���x�����ę��;��h1͜ay�>��oR�nv܆i������*�;v=�k�Ô6%��M-(dv�I>Uj�ú���&�c�s<k� ��Z���75��l5j�(��p���z�<������ߡ0��	_R��S��L���XI뗬捉D��Z�.�L�c�ʖM�-^H�����1���N��-�â����E+p�&P�{���`����ޱyϮ�s4}�o�,ng-�d!�r���)w���]�#S����fZa���c���p��Z��@mG�o��w���l�w�eP����A�=5o]���<Ý���\��]ֆ��#Q�c�(�c�Mu�O8��k����_qS�	 �"L#J�P� 4�A(P�@� ��>}��`����=W���n3�~��=�?K�)?!RX�H�g�v��uVD>�iO�$Jm���ɭ(��(�8���V�o��!UG&P��K�g=y���K���<�{d@d��:!�1,��IM2��Rk����c3rLx�c��ߺ�9�*�~��I�>h���� ���B�he��~w��?1)��ڤS��o���c���#�Jou���w�c��
�(�?�f��JY��82�vK�R/����i ��ȭT�O��u�rc�2 3y[�jr+��a����>G�d0�aA�"m	����%��rW\h�i�o3���v:��K�} ��u���u#4�A�Ӽ�V�6(-0�����}�*qtڎ�At6��+�U�v)E�H�2��w=��:|b]�6�8��@C`v6k�_I�8b�4!�)�0��o������,tA5mvJO�koƎ=��QaU,���ͽ���Ynn
�ҸM7��?0~�Q�Q����Nk��o�Z��S�^5�O���V�5Z��_'T�K���t�&�w�U�L�v���Dy��4��ω�N���v���4��瓙������gg0W�:e����O~_p�YX�/Q�5�ć@��S͊b
|������2��m���E������rq�޾�wEM�%w�u.nܞ^ι�2T��aTe�RH��;@��b�r�L�fJ�� ��f�F����%��Z��L�~|���	2%�)-(�0B�̨4IPJ"I*o�~yy�RZ�a��&(�s�ME�;��v�h~gh���ìs��5��wPn}��Ly��QDj..�SZ�\�ش��$�/\�o�D����B�AmQIז�-�w/"-_L>�nzr-���yIO�,�4װ�iڼT���d˴�}kO@sͼ�.��͵�O�"T׻�3B�����=>1�����6+Z��H8��1n\���}͜e�)�>��t�PV�����Sd�^WtWE�w^@�����c���߲���t�����P%�Fm�n��w���Y{�o.��V~N���[�à\�%�T����M�Ʌ�^�k�F):�)�tX�I������ʢ,�Nû&���xT����7_���g�%ۄ��M�pɕ�O!�s���}��íx��$hZ�)8�ض�ȶ�э��i�H8�C(�]���Wd�X���<�~v!���]�}�*L���X�(���o�g�ǣ-��B1��kd���2�vso�[3U7B�O�` �c�n�|i�o�Ky4�Ⱥ�Yyiy@��n��o��}������?�����s���{O����x����8N�}��3�x5�)����<��]3�⪝#Q�������a\���_W�u��^~���=}�_f��	�l%������'�I�K���y����3'i��6nb�K3�DK9���Q�ں݉]Y��c��=#�aƥ��I�9[����Ӥm������Mܰ�)�1lo=I�B�f����
��$L�Q��ӭdE������*��a>\N���۱4����:3���I[{R�,s�u�6p���oGc���_��M��8��I�HQ:�[�t��&��,�=�V�N�Q�{B�R�,T�Q�`�%�[��z��Ce�����p'��עuv�&ߟ�Qm��3�W^���)�tz�����x	��Y�Z�!�{3Esn����÷�)ę�>���v�V�qQ!e������*�j�Nɦ�]Â�ى&�ʏkw/.�A���8�F5���Q0Nqtg9�����j@o(�E)��	f�K��;T����[{QZ�L���;2��ə^	P�<)�;�>����8�vy��%�+�M�1_65���.�(�2��4a`�6�V(�x��t�[ż%�Β�'� Pb�AW�����Z�7����ݤ�����g��k`t�Q��֞�M�3�Mù:�f�I��[���.�ǚ-69̃�=�a��X��w��\�㝊F�(γJ�q�H�Ce��c*7�ڙ����L��q=��CPx�������C��u��6�K\�h�Ζl �[;ȯ�i�49䝷&�}i�.J�m���g��Q���F�E�vg��JǺV�ypo�z��n\q�ܠ�5g+n�t��O�R�"O:�P����E�(�SE�n#ʫ>��Nژ����| ̐y�l���{x��C�������O3��������K�jܳ���j���Q���d57=�O����ر�ğV��gE�M����p�eu���kʹjJ<��u[�1j����;UYغ����+��$�p34v�X,!��(1�#	����Ch��;]%[_]���~�e��*N�vN�{�]@����.��'n�U�ܒ�e�
\c*�N�ڹ��,�����R�Rv���Շ���u
Jo^]�"���F4�8��a�����B,�4v�T�o"��b��iW:�)��.An�+�kb��w7iRy5^	4�l���� nxA�r�r-|Sb�����˱L�r٣�r��b$�)i*O9k��ˎe'����jA	Pk���=�(�z쭠��L���'W��ǖZ�q1��j��*^����}��=�+��Ss��Z�����$��}��=V�<���v�X���b��!#�se�&,jC���WQ�`=���n[/���@�R'��$�v�{����"5����/s4KAud�vW
�u:ǘ#Q��SD	��Ms&���}%��45,Լ�Ǽܷ��Ӫ+��D�;ũ���[�xvu�As���r(�y����6����u��Ɔ�t�9��
�-so��si����E3���""��:��ry�QWq�lK���U�cF�A�����#�b�I��N6����5��F	y'#�h�F6��n�뚘����"�4U�UPw�\������5�[`س�STDS�m����wJ�1�Q�0CTD�	�8�6��t��Y1S�F�tkՈ=�\��y�-�zƚ.mP�%��1u!�����sb�$����mb���ˑA�d�)�i�fNlP���**j	N�������q��֩CF��(�Z
���R�P�PUI���=EPF����ij�����;����sEV�lh$��i(
�e�r]TMRU!U�|�r��cK:������}�w��W�<�|��o~�0��9�'ߓy��B��{�=��oQ3Ċ��g^����V*���}��Xo��k�2v���;�������f��7���2�J� A  R�(R(�P�(P�B3{��f�j�k�X����� �9���2�y/�&D��L*�.xn9r�Մ���v�������%]U������:��!ٕT_���&7��� ��"yķ:�7B͹��.�TX,��4*}���;�wL�S�5�Ź�Z
��~/�qZH ����}ni�a1���-��B���V���b�֪��q@�N���\NY�u�9=����{�M49XK�+���<5�,��;.�s����
�f���qW���5��ǫdr	�k�f��j[��=�V
��D����� Ї9���}x�F�Q���]Oq��K��3jr�
ėj�7k׉�%�|tE���l�����TR�yO=��f��j,e����K�
�e�6���"�,���	�@A�9{���Z)5.��<q��1�7y�g��<1^��8t/5R��Db�ӧ���{kݍk�$<��� �x�����3�E�c������d���C���>�P� ��a�q>S�V�%���ʩlj�r���Xn!D���D�;�Օx�6.Ֆ/�a��z-�z�*�ئxBc`�-bG;J��H�z#�D��˾S:�ם��ח��,u��^�C��e�X{�6����藤i�Cb�tvА�Y� �S��b�����=�P�%2J_�����xzE���ͫQ�B�R�t�u�c9,�{�pԢ_�}I]�{��cݔX��6�H���]���|�o�^�~�@P�4�J� L� $�P-�@	Q*s�]����Ѳ��ֶ�h�ڔw�2^�T)=�G(]�t�T1U�e+(�����2iB��qQԎ�7F!$ �z|�Փ<���%2�%:����dR�����𞀷�{��8����W��4N��%�d5����0/#��>�5��):��%�u��cI*L(>��*�;��m��/�z�|�}�V�2q/��,�����*����<�L7�Ԣ�9�����QQ.��4M7FR��{��@;�׏8zh@�63�tݓ7Oa�F�҇@⮗Q��ATԸX��M�WO��Bb�?7q��=�O�{��8O��xt��~?��f��ʃxR�u��Ԁk��M��x�Cx��u�����w:��Ӈ�n@p�A��[�C�Z��U��ʍ͌�Y�'�KV��51PUk
�ҵ�r^������]�v�;!t�a��S*z3��ެ�U��0F�z��?;���}�lo�U&)���Q�N�1���Y�z�]k�Ǉ��D�+�*�l���A/>����bv�P��E���e��^�"mx�������5
�9�^�dL���je���*ʰ�R�x��\q?,��ӟd���=̴�=|���W��*�4twyP��z�<��Wҥ�U�Q����.�Վ\d@n�okyd���nD��c�6e�\Z�4��_L�|��׺��[p����< `�H$���E
��D>o0��7��of������sem��[�ǜ���3%+�DO�>���=���|�x!���4��"��<k�ס"	��#6��4��C�|���>b�D['�hθ���_�[���¼k����t���f=��umtCA��E�SHݸ55�s�Ԧi@q�è%t�r����\]&lj�;�?��<��Z�1/ӑ�\���.0q쇵�Al�5{�T��0���&��$v��l�zǫx���X����ݝ�u:�I�����r�^��J�U�7���N��mA�ZQ)�Q�`y��=oV�]�.�����g��f4�t���� �ø<0�x<��VJ�j�D �R1,��Ji��)��O9K��=9MKOw>��zd-�^i���A�>D�'�L�0xO��ܫ��$�ħ5���ma��b��Ȯ�z�9��Z��nO3c�:���a��@���kޏ��ȗ�>��y!���&�Hw����M���fi^�s�~+��(��,9�񝇧���[�@�4�"uLXm5���%<ٜg�T^�iP��OC�-����R	z\�GR3L$�������_��������՘�s�����a���Z�'�M�wTlJU.��ը���Q�N~�TV`�]�L�xE߬?<(bC�2�O�vn���䨺+�QW]	ܴ�6\��JRd�y`��G�O���9�Y�϶r=��!�;�WN{���9�s��}�����}��S(��*��Ҥ� ��8�[o+��p��K����:���(�PY#Xˤ���>;����61��3=0ӆ)�ڹ\;�1z�1t�z�s�L�b��5g�JO�kL�z�w��i��ʩ��s�������֪3��Ba �Iݛ�K秡���MV�S���X�OO���{Z�vhz������a��Z�~�41V�1�����=h���T�xW�����w��'}�6�W��L��<�hO�ܱj��&U~���G�?�������+���]+s{�;�|�k���&�3Eڽ�]�gy�!=�ߕ~�-?V�z-�Jcy���3��@����I�eo�7��2��mӾ,�^M�C��i�Z���x46E;���x�[T��5'lR��a�-�<MG�{6q���qV�栕�I�z�l�'��F=��;k��iwyS��|9RZ1���߃Y���.l���2�!?5�������KIm��V����V����jV��ІL��d�C����(a��x�m]:ɫ�0���#���O�*����Q�=Cz'�8��jc;S.�f���<�x�Gm-DkJ�l*ͺ��_�mڲ9�hc^������tw�K�����|#e�i:R�q�LK�򲓷J,@���F�2i���X�i�E5F�t���/0���}:������|  H$~�eI��id)D�篯>|�)�D^8]o�L�?zz�
jvN5uEê��x ���f���Nӹ.�V�p��Sd#O�d��V��:�b��D��	�JN+�t�Ǧ���� �3�AƄ�荎g*��w�P��]�i�2�;�i2�b�t�.�2	gןh�f�%!}�ϭ"�9�ߑ޻C�,���` _��1�/�;O�g]��"���Z^�=5�֙��Q_/�*˰ld�	;����y/�:�
7��
�����R��JK�e�u���dٖYU�=�F�҆Sû6o�7�����0|n����ׄ���u���-X����L	�6�p�>Kf��'S��uʏW޺���v���h- �?|���ZxȀa1�OH�����
�Z�n9�hW�� m1p�sz�T˂�~��`�%�����Nr��A���+�_'!r]qL�d9n�g���y�𩯷&�s!����m�a�v��nj��^�{�|dK��Nнi�4b�p�� o>\�z��:��e���E�]��f�rb���tg/޿?�`�/���'�o��l1���kA�7����2�uu!�7�/A���}��Ofܧ���ܯ�o�LH\'��h�޵+�Xt��y�~���C��D������ٝ�����t|�9�=�{9o��W���x!�}�N�#�.�jle!EI!3�vTΡ���O���w��\��%̣@��U�e|��]*w��.�Z��)�F���ާa�e�zA!�4���h{��&������G��gB��뉷�����cG�����2}�qV*8���Z��_;9,P�^�q�ݺ͗���W�A���g�-���s������+�<�S�]c*��f�f5�_��\%�p�E��B��;1�R$�*���:k�5�L|��m��7u�L8҂[4�)򸈵MրUR����)����ʽiP���ȭ=;�X�o4����O�f	�%�V��lus�����HM����<����V�%9���MP��w9�^��xOv���,��moY{��`��sG���������7ƽ#ze'X�%�u��)�$�0���V�7U˨���#�f�˄��>��H0͓X*�E�����"U4]��(�a�mJ.��B訖�/r���f'��{�X�b�g�ϩx�HME�>dᏃ��~�|�=������n��s���oGDn���z.��r���T?2a�;`>��CM�"8F�FėU��zf�38CGt!��aiWp�^n���J�}�ְ��A���u���n��]�K��Z\H�91!d�<���]��OU��J�n`eQ�|�ɷŕ���#��n?b\���e���y�ڳ�}�u����� x|�����{&ܮ=Wi�2Vu^L�Ј�5mN3�Xky"��z#��XWC��di�zp��#Xw����0)˪���^�ô�Kʜ�d�����%Z×B����N���]�v�;!tϧN�O�}���5]@�y�y�b��q���عR������z1Ɉ�'�Y�M��l��i�֊����s�����0J7������mA���ߧa����m��E��x��$8재ߟ��<؉Ż�����v���-�F��q������\LJ�/s���12��Z�O�����]�f�ՠ'�������G��_��n���
�e��'�OE�ٗМD���3ff��M�[��0b�]�L�Vd�4
�P�%���/j|��)i��T)�|a�������<>��,Pm��D�ɼ]o�j}:�fg��Wn��ʖM�-A#�6->�7�~چ�$��P���>�Ρ������}O1q��3���^|@�Sm�(2j��4��(�0�ј���Ynϱ'�/�|�﷾�N}t�-<�v"�����?D���h�U�]�q^F%�t�u:/G��0g�P3C'm�3�zX:��x-��dS���e�T��x��C�7>�ne�K��\�l��A};$!u�����*[P�s����p҆Ա���X��U�s�v`�>�Cm4r���91��g����]ŀnĝՂ�{��}|�뗯��"(�T�Ϸ�w�ׯ~/�;������++�+I��]�*a0]� ����C�%:NH)��s. �ܹ�ݷ��=O˔�n��&���X���<��A��'Z�g�s��WHP��;3+X�N.�jxp�%�Չ�<�)7H��K��az|�>�h���D&�27^2D.��1x��Yv�P�)-I�
�k.������
.B��:���	�?Hh��Ϲ�G)͘=�������c�u�LKv�*��E�dc/�Gs�|w Ļ�69������<��y�NE(g`��K�;'�Bz�s��"�נ����(-��M�X
���n���{8���p�)�Ч��Y�1�]�:��'5�h�B�.���ƲǊ�6������#j�]��WL�"�a��۵�6h~g��&��v�x?��hJ�rl�ʑ��5��]a����������Q\�\-x��HX��z^��%O�{﷙LD�P��EELN�k�֣1��r�A��ŝBh4]�q�b�\��DYz�x46D��A�7���yV������3[�}��c�OF_�T�D�1��+P�J��CFB��7ػ���;��Nm�ܢL����j�;DOu�����[7�R����^������xq[lu�f�"sgg*r�[�
3����B|�6��of�eNH���s��� �c�m��N��jV?xx{��n�Y��`��3��|�J�m��z}��3M�Qwj*m�j�e��Z��E<�J-��=���k��Ҝ�U!�>�N�L����ϫ�6��� �qe�nnJ䆠��g7VL˱aKNaM������t��N�a@��;�c�&�yQX˜���0�	�/�ts]��ȯw�m���U��W�Ks�����A@��C�;h]:ɲs��٣�zMn�7�<oS�����~^ĨRo\�L-��8�uB��9oW�f�t��.�s�7Ͷgu������ �u�2t�?1)̈́�W*�qw8ñ�`�����+�b���u�eW:��K��}W.�E�K���L�1������QzH�����|���\3�j	Ī��o���A�?��#�{ K*��������Ͳ.�� �yryk0�I�Gܫ���#��Űp۠���8{n���n�yO�:�
7�4�U�?A�>����fv	?d�*~M�h&�30�瀣�~�m2'&�/q�P�/�H�	��	�x�bE�8����=�����w������c�j�+7u[������.�c�\���p;��S�B�O�D��ׄh�X�#{v�3��i�'�F�|���)�<ʥ��5�l�N�g!�St[��ڭ���!���<�O�\Nԧ�U�F�ښ�8kM����� =��3M2f30�=��1�S�7��i�V��3���Ѕ��u��|}�H�׷H��D[�b�/nx�� y3���~������ʣ�H=bu�s�w��0q�<��ls8��#cS	��ە�GS�y���;.ةm&�R�HO�X�/7��P�s�C��^��%k��qL��,��Б�9���2��	�v1������aDėj�7k׉�v��-���dg��MQ7���5=H[9yhwCF@�������X�8���;��Yy�zA!�3�����u��M�p��#t�s���P&�|ğ~B�x��zlݍi��C�6M�T�4��'3{ַ���X�X�F�L���7t�[	�}� �O�:N'�2=�I�_H�E�+���N��\Vo�����b�P��J��zzq���*��3ǐ���0Lɼbbu��dܖI�:��q��IvIO27�R���D��`&G֕
O~�r��ж�}U��Y�ڧa$�O9G�����L���꘿2"��"ʒ��D�V�%9J�T-�.�{��������^>�/W����z=��W�����x����'���lv���gB��!��,��D���U�]��et��=sۗ�Nxi�<'t++f\D���An�e&3�*sQ^�e7��r!t���J���� ���vaLȞ�7�x�k����Ԯ���o����lxo��3}�o��	�̓7Q�	�ԜE��H�T�u�b"��$�P.�6��Ü����Ńw���^c9��rvtg6��i��.�i��Gg��{E�8m"�a��4�&�)�3��1��en����;��1A�w-���x|Z�/Q�K�60��������-���뢣F����� ��0�#�ބ�����=d<SoQ�ٙl�I��(v�Lˠ���QǉgV;}y'�o v�w��ı������:�����Lsf{��'���^ɥ?!JG��;��O{��	aK�s*���#�k���~�r��7p����0��0�l��pl��jK�dǒ�l��]OO"Ù�Q���m��������f�z��q��m֙�cw��{�ΡF0�e�ʖI����|u������5`���� �v�{������h=|.o�`:Y$΀8��>����{�cL�w'�gW
��Q�w����⪓��²�Y㻫�1X��}�IS-H-�wnkVa�g�ZT��w�S/�[���,Tx�eD����!�%�ʸ���{�id�)S���u��b�X]ϵ�VǰI7L�1��!+Ր�:z4�UӢ�.E>��)'��}{��p���}�\�p|�>d��5m�Nl��u~�ڗ�̌j��1:2����H��y-Z��"&ש��-��0b��
D1���W2#��cm��J;�79`m*8�����쑻���\�Ȗ�_cli�����E�|I��Ivd<�.�`Ղ�m7�P�{�v����~M^D>ِY��=Ww��,�
k{E��	+���XA;�)S�2��9J�W���oh^~��Tq����D�k��|�H<6,J�kz4I�%���h��5v�g���O+��3�%�Z�'8G��rv鍲���#Z��k���ж^��b��&_w����{�%�a�A��Pu�pL�;ǝ���1�V���#�.�ᓢ�H����Kn���uդ.�u��z�+cE�w,�
�i�r�`ѓ�,9h�ܬ��k4,�*v�\9�1ʲ��r�"���h�d�O5���K#�T�]��3V���É.�N�2� �&����O���}w�f�wt�e]M.���%� ��Z����E�̺_<S'[����K���a�#;5�כ֘2ӽ�c|d�R���U�7�Iv��L��y.���]���m���iɩ�=�S��A�|���[r䛼o�O'	�]�B#������&������I��۾��/)wU�"���L?7���n��$d��TCr�7�������k���3b����2־2}\Rn\�p���s��MS�<�H�
��_u�pPhM�9C F6 (�
��Aʖ�:�����I��65�(֝�t$T�RC��AUX���@R�'6M.�X�G$)��i���I�r�UC�r��U%S�M��&I�F�^�Iɠ��lW9�X$).c���TII�T�)�I�F#M�h4̴i�%��lP��JM:�s�������'%�r�'�Ѥ�Z4�CI@U��R�m�U^�z:�ur�k[��͹S�.�i�:�\��T��Q��:�wsu��Z(J�'6�W\C͢4m�M<�Ӣ����STQ����~�oWG���FAE��A�ߩ��yo~����U;DHB���.�|ji�RL�WԸ=��JilP��xw���=κN��V���9E����u�P��0�W��cu�sus�ۧ��n���"?]z����u^ϫʓ�0*I���G�/�5y-�����By� ��5����N�1�d]`�c3p���E�٤k�2�O�|����Y�L�����}ʄ^���J��.�����n�B�	��``Q��ɋ�U��<Sq�0�_e����8zh�
�����	�Ga�F�N�ܷ8{5]m.�ewLB�q�r�2���pJt�~j	Ļ��}�0�t�Za�����讻�jkc;��oc�E�NP��`��²�߉Te�dw9�R;����Ӈ���!ú���6���A��8����愙�G�SS.��XW�t�{J	{��q�!]�6������])܇�S{��R��p�+�A���a1a��h���C����M��*��x�|�gӯ^&g��:LǄ�cU�BX�w����3qa�������:/p��Ӱ���d3l�J/�X/��L��U�����,m|�����ЎEx��E�m ؇e>1.�����\<(��'c5��A��;8k]P'�_o�V�xq���@"GN����EC�dK< ����Za�s���5`��q��k�(����VmO.����?ݦ��t�U+���`�0��zK�9�o7���a���ޛ�&+�呬l�k��PY5a��D�9	�Ŋ.�f��x�f��g^{l��hg��^�N�n;PZ(c�n���+Vr�n����0B��h�_U}W�&vO^�ƾ�c�}�Ui��L�^�X�B�R]���O�~�-3�S��	x{,z��u�_����
���œB�:~,o<��2䥛{�eK"�Б�C6q=cռ"B��[n�>Emꮊ�-�kG�:瘸����^}��"SmzѤ6-�M��(�0����S\���;\�;	�]3�j���U�E/�c0&F~̑�>�T�{�p�6U[P��F%�y�s�Y밎T&?�����h�~���ߧOR�:&x�^S�+I��2|�8��}�X��}=����T��-�t�d�׼u����H�o	+Ml�q͡�.s��f�t��pLpdA������Ny�,[�3:vQ��j�R��9zN�l	��5���/O����G��]]�e�L�+�Vٜk�0*lS2Y	�=��Λa����L���iR:�3L$�쥯5:��)���������u����+�Bp������M��u��.xo%�5��%�I��wV�6�z)��\��������������,|�[��aؿ hu7�W:��.\����E��Zd��y���ڇ�Jުvz�[|�}a}��N��צ�����������ӫ�S;
�n2MlL'�V���,k����'vz?�9Yd�卹�	-�zl�`���,w\�[<�v��Z�.��F��ۋ�)��m�vc㪥llҘ����磌�Z���g����N]������]X�P�n.����c�����ML�0����u��0�������Z������5\���a~��Ph��������mqϕMkϲ��.$�Dg�����Ӻ���s�`'3L( v���@�r��^ø�xg�,�KChN�ov���+q��:h�꼭3����ק�&F������P�&h��ވ����=�ߕ~�-?P�"W8߲9�)�}kN���)�C"���?g��m�oO�,�4�='����A�r����-~|(0�!�������3|��nQw^�%��Ľ���WXͭi��H8�0�sRW$5u��ޛ�%U�x��ɇؿ
+�T�ǘ���N\�rO���C��]r�n���nwf�e^+�{	m�'|oY˜|nQp�W���<���v��u����sk�O�.��n��V_n.�C3o�k�E��{��_�*�U&��j ��:����$BoG��]�=CZ�fg�3�2Gz��ba�����A�$�ħ6��j�*�qv#�H�hT8N7�����{"�y4��ݘ�WW5oQ��ir"͍�p���N]2!���Ӷ�{���+G�4�ݻ�����`��m���=w�`t��@,ן
�j��<:U�og ��0��j��j��zwCG�\F�	�W/Uˑu�=�g����Z�YڂLR,�'�_U}��)<�o
&v�>�A�v�ۃ^�;g���e�`&*�t�.�2	���k��"�]�%{7�Ʃϕ&Fb|<����mdE�i��)�ɛd]`bށ�4� h�L�:Q�ח���Ste:W���Y��8{h^}Cw=	y��У~�I�U�\���ʉ�E�T\��n�6b��k��)�#�;�5��C<���X:n������W:��{*��5W���3;��̸���`����WZ����g=���(x-=���ly�}�(v���<�AE��=�J�Z��%��,���;���{J	{kU�OX�j�ÿH��y��)�R�-m��q`�{0���  >�ڝ�e���,9�
T��5�`��;N�5-�G�az/a��V[���R�^��b�OCmJ�\�X3��V.���u�e���,4]���7k�&e�U�L�!=�4c0k�N�8��ASp-�}�.�0&tF�!�>0�ۜds���"�}6^��HzM�׬M��{Ҳ�'i�{#%:�?�����ϳX%bO��!?=���o�+��ܸO������v�O{���_�i׏�c<�7��y�3Ƹ]@Z�W�A�0=�)�����.����Er�P�˒���ˑ�B�Q�I���CH��.���u}o��4�`Cx5ZM��L�$�e��&�gEN7�<�&���{@b ���u	�E_ʪ���WXپ�'6�T@��>�M�Q��*���F��덷M]1p�)�=���8���.�-4�p�x^��Qct�E��n��U-��@Z�Yt7�V,�K�p�������U���fx!6��������n�f��t�%�8�L!��m홆��t!)�ѐ�ZR%?J9B�Ӻ��O�b�dnT��)y�Vɐ@�4�q)�0	���7�y�?!)���Nl%%�j��^�h�k׊�r�R�su�&�S�o��8i(d3�߰��{?������������a�~�a�VAO��k��w擙7�U�b�.����Yp�Q����a�$E�S��%�c �H�fS�>u`���b����2�V��q�L����T2�<�>��H:� ����8g��y���2���5l]t�謍Z����^J������^�ش�rĮ��IĻǻ`>��@`鵋�WO�}O��v5m�Ż��m�2$�^�6��b9B�>Le�dw9�R;���4�^�<n@qH#�n)�fKy���+j/Il~���^aq�p�:�٦޿uQkeiN��#ҵ���/tꟘ�C6G���#;k���A2e3!'�t���;�Aj�������1�̐\�h'ƕ�	��~�d�������'�,JŌ��e���"_���4���g�}���dfl�[��No����@_��O�~�W@����f���-c:1C�Ø��wll5"���U�Uj&y�Em�Z�R3�
�"wf�M~��mǽ�]Rci��џN�{��T��.�SXE濗2��f��E�v2g<�о�E�'�|���쾟yu�-���푻Oyw��j,;[����fww����lZ��<��<��Ņ�Y��)M����t��y�1lj�j��7|�a��Ș$=qhHM;�O�؊��vĳ�ZZP�M{w�TeO.��z���E�]	1i�WHּ�,�[ÉW������/e��R�3T*{3��_�>�r[���T�PX����##)��Ҟ�f@�<��o�Pe^Y6��$v��͜N������<d�oyj����S���I	o�@ȧx�-�X~�{GY��	^�W���Jm�O�v�Ji<W;�3����fyȃWjf�7j�]�۫z��z��x!@���� Wl�+%W5tB	��M��K}�n��#^�/5s��M1�)��5�G[�W��=5�܃�vl�L&
@�iv�9��]ծj����<+�J"q�vO	��ܒT���vO5>Eê�� f�t��_���6F.�/3#2]ل�e�VEcf�X��1�w�Y���tj�h�����YvW�u�j�+v-��́$޳R���Ӎ���v̗�\E���K�:7C��0v��:��'�ڮl��*�w9T��8�Xْ��ފ��X-��'t�����\O[f<�l-���A��R��N��T�㘤�`n�F��a�^&0�c��-�va>Eќ7��;-���ئn��-E�
�i��M��'^,YH%���%��,~�-�E;�j�F_b]+������|9�>�[](�w�Mvz �� �F�x�$�n��T�J��h����$/�N$qqDW������z�P�u�rf���JO�]��>�wK��@�˵z_��������H��ʒw����H�_y`������t�-�d�وP�i��,
�c����+�Ԝ�I��F���pb�^B-�O����W��/��no�S~��/���zRpJs4���x�sQ~���3�Έ�v�]ػ�P�-yj�G���(���rdkr��χ:D.�8˱i�.�|tE���6�L�c��7Y�z��9�g��]!n���X���lON6۝��z��3M���T� �9v��68������l��w�Od��b�Դ�X�X	�X>B��c�Q|W>��fִ���qe�nl���c)t4���xq#]Ӝ�+��iN���u4���!u�XL#44�l��N�i:���|�j��n珡����J4Sa�O0�A7�~g���k�8���b�%�vu�@��jڋ �Rl7Yk���Yͧ
2��x�,�W{������->��=���z	כ��7�ӳ���͌cY���{�
c&��~k1Q�=�)�%��/F���ς��s(�V3��L ^���Y\�՛���@�~�|��O�cO��K.������qj+-��M̂����e�a���(ʤ��j�T\:�q���$���v�xTsc.���}���Lڦv�jY�Od���L�ߜħI��I��t�Ǧ�֟8OtC��׹�'�cx�}d!�$C�c;r���z�oR��	�M�me�7 ���2�Fg��^b��;:m\��w6��s G#D9	����!�z�Ӵ�����Ͳ.�u�m�4�֩՜�ݎ37��W�Pm~�ʂ\W)�e�>ԏ����C�~���g4�a[���=��)�L�l���\nW=_��Ƽ��0�'�vh��lm�&�	��	�t����,��n�ǲn��1t�w]���Μ}W�֑�t���h'�W�!��!_�~fWL =;Nv���x��Ʃi��X����C(X����Oҵ�%���Ts�#NV�@��/�~6�5'4<�|O�(Ѫ�����<�=�����`�f�tn)}�96R^���$�{�� O��) SU4�r�b[��WaGM�i4^4gV�d� ��)R��"���z\�7�t�c�����}ǖ=/����gu��%>s� ���w?o��?w�O#��]N��Q�`�b��f�!�m"�9��v[^�Ú���o��f��O`fl�v����-P-������w���a��;��&��o�9.�:��.�#QaDėba��۩�B�JCіս���8VG�C,��@kW�j�|<��<�j|��na��K��z/2��QM�9�o�Vv��BpW�0��D`��g�N�>�����#�݄�f���Ѡ���Kue�4\e��㼹���Aϩ�d���\�(r5曍�M^鋇U�L��X@��8]S�
|�HI=6t�N�f��Bj9��*���q��� ʭ]
6�p��8�E�T9������	��z��v�uㄏ��A��i���N1W�R��:��~FBeiH��(��Ӻ�䋍���=)���{�:M�D���Z���8(���J|�0���>�S�܄&\�%9�bTX&�-�:��Ĥ�!Q挹C^����~Ȕ����[H>`�'����3�ޙI��e��t��/��u����\�Y�$�T�6�󆪈O��֐]�,��s������X������-��k�.^ܻʵ�}�%�#N��ϝ���g}n��"�k���Jɝ��`J�D�:����@��Uv�4�0���^����J�>nQl�L����s=�c�t��$^������8OQ��y�e��윮���k��:��V�y��p��{�A'p�v����>��%R���'G�>�S=Cϩx��*/��H���	�c���4�e]��~b���7"Ji;ߚ�*�^�r-?5��2�S\x|�I�s`!��鋪{ނ��'�r��Ѧ�;E��`�e%9���NP�%Q�X��h�]砲4����u��5�ɩ������t/��_��ֿT��i��E���8�����^��+�g�v�f�k�&�휵G[f���H\Y��A_�9����GW�\Ȏ�Ζ��L[֢:�'�#�Y�v"������>�u�d�u�2��όg��2F�Eݣ_��:~���m3���2^�c��������s�ǧ����������Xh��J��1�g�O�~]�Tʬj�3Lي���k��/�7�3kCrC�g��v�_E��w�7/�6%�=�#Z%Ύ�n!�k�]�a��O8�̄?2ǎzǥ�#[��*f��X]+��p���~h��̄�q�Y�7:���Xμ���4(���u�z؋m<�3u��ʖM�-A#�����yz|}^^�w�����{�ޟw�������||}�0M����txzC��D�v������R��E*�/��=b�m���hH�mӣ��E1��u�
�����n\���|cY����.J���hj;.B�\�}dT��]�e��gI���7�hy��}��E�����NHK�{���N��Dj�+,�"Z��놖�;j�]:�9��Vt�J��Cf.ۏ����r��KR�o���͞�2�wI�GEt�J�ҫ�;X�Is���`M�\�a+�f���;*=��C�2�Ac�t��	[���@u�B�3��9�Ȓ;��.,��n�j*^b���QȤÈd�4���(l�,t���ǐ�.	!��0���
%]��q�t�)*�����;���=w�QՍe� d&<��U��ʙٽ�����c�los��5��*"����'k�.�ӷ��Lh�s�u�8��//
ĆNNV��`����"
D�2��&�����P-��(���{��wO5x o�[U��P��x��]���:e°'�b3ygp�8��ͽ����5٧\�.2��&��j��9�EU�M�����4��O��OB�PFW��T|�j�zsا`�>�,�ot� X�V����y$��@�M���T[��[uV�B�E��ں�5t%i\��j�rݛ_%7�fΥc�;�r�Yl���7�-@��Xj>u}N��|�v�1ͣ�!v~��nQ�L�mi�*bzR+��sb�K6�m�3r�\ig�Yn���ݺ�<��	b������j�|�?G�6s4\|������:}����������w��Jre�1���ιP�%ڮ�r<��z��zgp+�J��:\�GP�/�o*��G���U���zr��*��&�,�x��*�JifY�x7�6��ϸ=!Gc�a>IY�����ᜤj����K��8{�vX���ϯ�:�Kc=��}ł*�d�RT�g!Rt�F����^I�6N	�7��7T�����L��a]fz��?J�����k��ؗ
*�onfjm�]`�/{/x��+�/�7��ޞT�eW��|�W���S�x���\�:yn��A^�;Y�;��-����	��u��(hklҼ|�M��V�s�o>���e�������������ԸqbW#YZBq	@������E9q�o%�eZYF�z�#�a�.��U&��MK�@�Zݹ$W���d���j��__����\�U�M�N�-ro3Ԛ��ni�ܼ��Y��k��mT]?h!%�ۯf]�,0^~�n>��|JL��; 9b�����]��f����Tv�iX1�۵����[Ӌ��Y܈��ȖLN��\V��ԕ����ny�r�{�m��Ѻ��EM�Ή����?r�;�fԕ}�j+~���?g+�o�QM��{l����X�=���Q��|T'
r`�s�h����mS{�y_7�w���5^������v�80�T�� �4���� �m��u=�s�v�Eh���12�\�6i4�g�y5��4�w�X������͞'K��O3�k�r��9&�)��F"�M'M)H�r�rccI������:�lb���=gG���5EX�tm%�r�P�s��8�.��5���1<6��:����DGpr����,4ncA��9:(�܆�C���F�9���9�nV� ��lss��sn\��IAf�!�����U�i�������U�F)4\�h���b�9��j�]�.l���&�ᶟQ�[�kN�֓N+�i�Ŷ�9ˮ�ʜj�P���Dj��լV��9'*nw�u��V�8���
��DC[s�J�Z�lh!��m&��r�E:1�m�6�9�[9����Q�~���
�SR�h\\ǘ;�l���M�J5�{��CZtt/�Ӻ\c����[bii�����<=�Zw����U���ޭ�W��A��`qm��]��aUc�mEz}�D�����/n��뽸���h*-�d�k�W��;#�瘫����Vq,��08E�"!�˶A����P�L�8��~�:���+��xc�I�bd�`)����t�On���(���S	�9-��A��IF�oZ,���הD�I��Jsk�SIRkg�m�.Pq �5��pk��Ucq�Q�^�LЦe!d����3z�$��)9X�Q���j��������g���0m%�Ӽ��J/!b=0�y
v6&n��%��
�n�9/I��Η��M|'��ȻZ�~޹V�z�CF@aä01�0�s���Z���M�3�s]�^(,��e�Xꭦ֭S�����l�U΅�;�>�E�xQ��k>A�ʚ4��'P�_X�"�Ђj��>��?q[Y�Jzzc��-=*ެs�S�cb�ٶF�p@�Y��Ov���@����@5<�v��h� �s<��x�X�OO���i����A��YA����/���������������=��brk��K�M��#ѽ3N�;Ñ����^�}��>R｀����*�m2�y�r[�Qr�ז�.��{��ӯP��K|��9�_?U6���S׹Nt�&q �-��%�MM;����UB���}�)�_��o��:uQ����4��i̢+����5��׍�a �2���W��v*Чr���ޛ���!�m"&:���lwPnys�M4]������`DYu	��P�ys7Z��W=�=��n��2D�ǈq\s=�a'[78�npoHo5�f���(�k�����#��q^;v��z;��E^'e�me�m�P"��'A��ȼMG��6��l$�m�j��l{�y{��xf��YQ��$εC{6q�dgO#���X03���o,2&�e�����Ok��+;�ŝdG��{���|�ۡ#Z�@��Ƭ��sn��X�.0�f�x�/mV�=��wX�/J�d�y�?A��#�g���J�RaMAvN5uEê��r��W��j8\�JmgZo+o�f�酮װ��;%75y�$��%:���g�=QI8�ӌ�0aA)�;��y�ʚX����g�yaG�5��ۈ�3��Df�*L��� �E'�:,ԭ��V����x�ӳG��2�{��N�o'�r>5���^�s�8�Y|i�E�IO3��{(o�|]�d��k��N�;����}��gSy���4��i�42�4v>/53�a��Ɠܐ�Sɸ��w|A�6qR�����1m*�`9Ξ�Y�t�dX];1�⭸.�z[�*��İ�uŗW�7(��[��p�ٰɵ����r����|kstX�F{L�d�)���Y�/ �0}�S��s���r
�>ԏ��Y S��=���/��/[�]�V��xR�PFx��\���'�m2 �4����h,;_���yU�s|�[���j:w6���F��(zj�Zc
�V�U:9������o�@sۇ��@���PM�|h�y4��Tn���m�-,�ls�}A7��\R�[�c�@A/mj��H=bu�9�`���Q���7vj33H��!�G��X1�"�uBv]��mՅ*�~�ǿ�4�T�5-�G7�PR�Vz��i	.��3��)�|���,Ba���:;���0�	�.�;dbm��{�ͱo6�`T}�1eyOڢO��&��Y���>�c#���4F�-5�'�äz8P�Y�+��o�Tmv��-����466�%��c2Rz�l�ӧ��\����^Y �Z���|o��������r�r5��t�P�^Y��,!�-������#������~��xxaӗ3l�)��A�Z�l%G\=��.b��{=�h�Tۥ�J�E�/�4;=��vs�Ѳ-�'��j
�f���0{�1�]��>6d�Whޒ��;�h��cM���'����;6?�o�=����sn1�w����(���.;+LS%�B�8�]������DE�\_H�9�Gv.�U�{It�5Ԩɘ�����u�i���_[?�BsO	�i�9�B��J��[��ذ��$Zk�R�	�f*�����w�@P����]�w��:f�z���)흴k����! _W�i�S�O�Jd�s	��t�N�4�!���������e!��C<6�'x����(L�c@"@�5��9ͬ�R�I�Ʌ����Y\�,x$�0��|�+��U�K�̜��Gܪ/���_��|��0�ᓛ�*o�sD�ǧ�ը���~FeX��i�n�`Ӗ�p��će�8|�E��7�:�Y:����\��b2�,T)X�I�Q�=/�"��$��C�&�~��6�k�u�]�r�6�6�����tۓ�\���6��a9B���F^�Gs��q���{�����iY��l��C��+p�v�!02(�8s��'f�WL��]	V���J״���r7� �'�Ux׉�1<v���B��?r��� ��9�����;��zm��*���}M1G)7�m�3��&#���1>1a��p�\�轀�㿊��/���tɽ?*|>��n::�ojg��uq7Z�7eq���c���5��^��t��ft�ը̖�meҨɋi���'�U��޷��fc�Q�՘�0���A�u�1�pՋ}w��R:/���53��BG �Y'� ^���QP$�ݳ�C?}���F��:�Q����;��Ǥ� v���D[�:�;�D���9aC�q����3���oVFf��Sщ��h1��X��.y��h�#��l�}���X���0������p�57�5�lcH��\�=���]#[�nf�����R�9Iw"�m?`n�d��r��F)_�y76����
P���$(-1���&=�/d	ƥ�S7X�(2Y��=k�q��x��yh:��T*����X��,�%k��Ua	^�W�����X|eʰ<:7�}�ro�@a�~{L��v�oV�^��N.��
w���5�<^�&�1�N+�6���p�Q,���YJ�]�u�753��On�$*$�6<�f�s�̈́b�4�?Db� SHB@�'���.��A�Ns�ȦT
T���y��.o�t�w+'ܮ�_�KI�g��U�i {�|��7T��;%��]��Q���'+�Q�-�Ø���2��O�U,�-u���"i���ǚ�wm�+�jb�]��P	v�����;c5�p�������׆'1�wv���'��F2�#z�fo�/�}�^V����ߏ�w��ԩ�`\G$Ym�Mww���/���d�jgB��f(�̶��b�ȫNn��J�%J�K��
wUͦ��̱\�����^(f��>�μ�� ם��k���S�;�ɦ4�~�l�Q�>�0�~e�[]4�~�U�w�Qx����Ѣy��4��M�U!-��r��^X��<�GVE~�k]�4~]��Nu�dS��44���������RS�Z�&ޭZ�zUܳo=�C7s�jA����6�/W��=(-���i��py���g$W7Aa�όm�=#��W1n���uv�v���k0L�)�.��hѧq�-�������v���4��>Nf�P$@�1\�~�����U�[�)sdd���0�`ygj��z&9��~o*�tf��v�s~ܹ{PK����@35^�	�4��vͅEռ��UzD���4dsLL$��m��{�yf���zO;?���IAp�h���n�ȹ2��b2֛�R��-��������[���όUM��?��U�>��ְ��ɎU�p�^�@��#Ϲ���dgO�.�`���	;�c�
�fFQ'{���v\>X����J����	��a�h�Lk��z1��Օj�3:
�g�ȓ�gܳ�ז�����%U��)r����VN�60�&�B����C�����5�:S6A߳n%��|��so�Wѭ��r���n���sV�qJ�Vk���m�WG��'f���CBU��n+�`�m�m�e�ӧ��0u���dq�ݯfk���Q��E�c�\o�bq�VβjɃ�A�e�~F):�dJ>�I�5�8����s;�66fsi_)让X�C�yl)f���s���7	2SsP��&I��Jua#B�)I�L+nl�QK�t����Jm������T�?���m{��k��6�<�/z#��_Ze��ښ���\��75ٱ:q����s�sǺo�;ռ0��B1��O��/�lyF�j��vQEތB�s����ee��E1�:��2���bK�3�V_�j��ܪ)�罯+�Sŉ����Ze���^J�
�R����V�O}��=��(�ð�=c��.��2���r��v޳�3L��IՉ7B͹��k�	TX,0X�WZ�|^���sۇ�p���qi����?PN�ml�:e�;�е`:��:���{	A/m`*�`z�kZ������,��cݬ��;u�����@��?ġÿz"���6�nIa�|��-�6���4�r����W�X�j��C2k�=�r`C���x�	�<F����vI��K�a�,���o�`�
���#�6�_m��/p��+���H(Q^='�{�׿����ƫ�TF{Uy��>�_r�m�T�tqn�eOpn�=@3���)Kt.�Ʈ�x<�t�[(�n�J����+
R�]��������`������^��K�6�Z��T�(��ً��O;~�,ۯ@��c��tg/#^]� `L���C�|aQ�8�Ӣ���B�6+�n{����e�% ��� ���j:"�P؛xc���	A츹[Q�v&�ț7���35_:j-=����>��<�}*�!��k�7n�����?o�3�C9?b�����<��$�r0@ ��L]�kߦ���T�o����`a�Z�R��}�8�c��Vm.Zk��^w*u+�k�zYPx:8`��n#���d��*[��A�m���*�����l��}�D]����cռ4����Qm)ė���y��5�E��j~BS)�	�z&;K�y�&�9���.��0Xs(IP�ػ}l���o��[Rt��HO=� ����;Y���lx|�D<J�[3��(�E��ƒU���!J�?�~զ"q/����[덈1XB�G9�)@nE4�J�}E���`���6�܂�n���p��=3��x�Z6����#Vч-�&he���B`��4(�N�⮗��O�iAcK�C�Rq.������3����"��Uܷ p�'+�o��j���.[�C��Z���r�ޑz��m�@��d33xcLb�Z��W�c:��	�����s.�\2p5i����'nfP�{ |��i���粖�7W14[]�5��:n]�#k��Kn�&_��?0�d����hN�W&m�j��.�%Q�����]��?I��B�k_�=�|6�iip�+�"���ֿF����Uml�)��w���r0u�ʝ�+f��E��~��[񞻄�s�N���s	���(:�0��{Ώӂ��̚����SΙ���1I�S������&g��=��h`���	\<�z�P55g��ݯ��D)�6��9���
)�j��f��~�^=%���1^�tE�j��y�ސr��S(�h~S���[�Fu�K�"zH�$�k�&Cɶ����$q4� ��N�T?t��ڸ1��Vs)�l����C��^��oui���j�K@���R]��=�̶^��'sQ8{'}X��-35B����������/9�z؋�:ԥ���v�eOsigH���Z�67��y�,5��$:�l�zǩ�ī"��-�����U���뀌�楠�uk��Mm�q��ZSI?��j�\-U��V�'�����$=�<�x��ۅ�m�^�Zx�����C�K�R��ח���V{.�zY�D�X�>�{+�����{�j��׳α�n[]x6Y�s�#t���`�IR����G���B�ɹ�����vФ&�}��iZ�(C)`�� ��lG_ʪ�
1p�=C��{���A8�bY��z���J�[�S�sS�}���^�D�,���.jM,�~�?4�L&
BƑ�}}'���:O�bS���)� ����Pm��h�p�۝�ӷ�nv����^A�mg&�Lpc>�`��.�w��O��Rr�@��h��}H��tTM��=Z���gp��r��<�>h����"m1��F��Q|(v�M��1i�.h��e.��m��bh�מ�3�����zQ{�]vG�#�5��H��\
��M7_��s\�9��v���ŕ�NvLl����Bn�H�~O��Ļ��(���ߏr֏˽S�W/����H�ٰ���^�,P���v�_��Zd�ի�G�T�f�;�n��?0��_-LSf��x����f�,����.���N��UV�S�^5�=����5\�����=5�S��%�{��ם�W@��!��!�az�����4�$�߂r�
���+���,���-oB�MqE��WR�����E���Bi���c`k%�!��ÝBk����\eطxz{}�=��O���<~?��������������~���`��B{G~�-�ܶ����<��έ�Mo8�NE]��5������z+s���LL\J�j\ʨ.�O�L..>�}�lN��A�z%&<k:�{��`Y��y�U��`ǽT���J�"����I�+ڙP㘶=�|�$qͭ��K��>�W��m�+��	p�q�k�ӣ��(7xQ��m��-�w��6n�N�ܽ��-�^m�h��0Zd��ؽ\^.f�mv�4o�Q�J����x����V�Κs�̋l�Rk�B�JEV�	h×}����}��4t�� ��R�w��e���픵������&x/�o�qخ�\32��.b��o~7��9��8V0{��y`��LG^|o�tz֮�d����P�$+;9�N̸��2RU=Db��R�$^+�������}9�<{ӹ��ali�|�x����#ê��
������l����)(�R:�BŜ�̌�I��k5by���v�����5*�G26/~�͝*�׳�<�
�+��-L�//�]�����Qn�s���z��V"�g���!��ꁾʅ�<��n���\��� �9���^MaL�N�b�\,F����C��ʍ[<��*{��6��k���S�y�uh�6q����&5eh9�Y@!�T{� ���f-pnΨ����GMmb۫Q[�<��s���"y�,A� ���fq�<�R��wVXon�h�B}��ٻ���<�@���Զ���Т�;��i_�6§�"b����p��Ͷ���
��+f��q�}!ݤ��F���;A�3RC�U��ie�uYYJ����n"�,��j�]ތ�ZyM;}Mjtq� ��;��P<vwͻ�nC�d9i6�b�<��9N��k7%�;�ݛ��ՖiX��o�7�	�LZW���9�_r���9ͽ��ڟ,���s��x�cf�*U�F��ԉ�<�q3�X�M�e��gt�rb��AD�x�bCz����xJoT���O���E�����m��=��e޳�а=����.U�d�D��r��6��.��Z���P��Q�ip.�D�0R��(Lw�}vi�X��v�2vJ�i��C���f�.�����z�<
����n�<+}�R|o���h��{GA�le�⮵LO�A���-d-E�%�z���:>4�kŻ��K^���C��pF��p��Y�a�Y*m��Pf��i"֊scxN�}�N䍅��^���Z[����Z��m"��H�*�f�����/��q{�?G�]mr�8.�=z�Q�d]V�J�I1+4��Tb��ɇ0\�N��낇ZDsQ���Y8������!�y.�[n#����{�｝^�,��MM�OI~}j:����a�lO�����MI�3c� d�}���6�$�@�!���3kuw-s�ӳ�9v��M��K���X0�@CK�'�'�'�F�t�c�<�
1	���\��"m��C��A����%�hӢ���N��z��'(��V-{r�N�hK��70�X��r��8m$\�$�9r֝-m�tm�j ��ʝ	�AG.�����M'7&���n[c�"�:ti�u#�*4��5�ܢ(kX؉�Asn��y4���ݖ�F�:�"!֨�u�IT\1�7,�޳��)�hѢ-*Ě���r��뮚�F�9�<����ÛCD@r9s`�r4kT<�8��E%��V��lYvƴQ�a�QZ���RR�%)M9�m-'�m���;��JC���`�Rŭ-`�V'Z�G ���;��oQ�Ll['pb��kOPjb��Kg?w�Ѳ� E# �QQ!�LMƆ��|�~8/� qR��8zJ�bCh��X��,��sV��2��=O�r�e�x��4�Yi�WG
 ����a��@�-�JG�n����D!)��a�/�2+����Uz�w^�͆v�|��J(c�hx�`��C��=�@yKO�l'�|f��W�']=8�npoO���3Mt��L;,��9�Iދ��|�M���e��Z���x;]�`0%��������W>����9���TZ2+t��yk �5\�����A#:�Y���dgO<���`d�����=�ͮ7�𢯺O9���!�_�������B~ka��P%�$uX�dA^��;�U޷}]ߜ�I!$�A���ahZ�4�LN�H=:Ųs�~�k�1I�W�Хr�0���'hMc�d�L�WX�[�M*��}g@H�ހ�K5�	;O�e����M�A�(�/)�["�n�"ڤ���;=�r�j��a>����� ��_|���Xq^�Gz}>?Pgݙ�?�?kW��m���qR/ױ~$�b�zw�xa;�!#~k���cÔ�b��9����A^�,N���vAuN�����Z�搴�C�+���S�
���ڠk��,�Z2x�i��ͭ���\#.P�4)X�I�P�+��\���+�a�gwfCrAã������A������s�����oo��[�^v�	l��:w��d�A$��	�g���IY��(q��[Y/r9�LO,gY�L��ɫ�Z��Y��6k�i��&�(��iQ�#�݊���t����
�n$4�h ]\����V��s1q��K7��ü�CdB�W�9���n�|Z?1��I�NlI�l2q�߉TXRΞcJ�Xh'ј�ŭ��,�獚O_VrqH0dC�\���sO�Ƅ�m�v��Υk����kߒ�^�K�-�$������k��K
���=�s!���4~k��췶Kk(�䟦��kf^ng�͜�R�ݏx��W�Աj�1= ^�90!߃x�|�	���~�NK�N�z]��S#���<Cf� Խ"����e��Ɉv�tE�W1eyMQ'��hy�S�>�;�����}zq�[YYϛ��������y��	E@A���c��tM�1��̀��j�,jd��v�����g� "���j/��݈�qy	��}*�!��_�=z#m�t=C�hd{Q���V�����X΂X@��L]�'�5�וR�ǔ�e�b�]
6���#{��O�7V����v�}'�a�LP�)�=�9��C��!�s���q�����t)�ѐ�s^�q���cQ�eս��HYt'�(]�M�X��2��|<��y^���^O�j������kޜq��9���r�����CX:����1?�[����n3�E/+���(&����s�ǩA�*���f��Dy0�vb����m ��xa����]�T������ ��T�l���f�x¢�q���[�d��uq��?�U�j�c���:�U�V���S����MP��v"�����o	���Hqm:A��!=Jt=�[O�C�glи��,k���ϸ��1�d]g���J�
�|��a=k�@�a�3�]\S��w[�ل��-aX�K��c@��_Qw�}]0E�,������P�@��-A�6��A;�%iɜ��ɱ�B�A�b�BcS �vw'qG���O�iAb�?3Ck6��"�ʊ$�v���h[�zߟ�A��֑#[�	٤�ę��a9@�09Te�dw9�����1S���a�F��x��zp��>��s�:�ꝚmV:����	V����K�����J�1�f�״�'�uO̪��;�;!w0A��c���_񣸽�Fdn\��L���]�%�i�r%��ٞOO��я���j=��h��ĸf�ƈEԤ�//2��U�(�k�;%�+�(81�`�#yWm�>�^�����	�����8Ū�C���.��o��r��6t�ԫ�m��� ��q>&m=�;��4�ͬay��Z�Ӵ��o��y�=�;��N�VW4:.���ogaJM��d�AK�P��|8��� �!�S�
��}��ޫ{.�/OI����'��|U��[�fGd�d�S���t�u9�y� �RT�W��}�ھ�#��\��4���җ���G��]S;^/���()6o?�����$�T�_�4�ϡ�����|!�z�x�s��4��i�_I`h�����n6q���.?ޞ={�������mw�.�f�S��a����1�[����,�a���m0K��`���l���|�1����s��ߧL3y��h?��<���(����EG�TͰ&ҬQ�t��ݏ=��ι�<2qx�[0�g^JPd�z�^�3�(�ǫz�����
͈���U3��}qm���3st�f���$�^K�*&��܄�|�K"�%��R�T���s�:y�����m��Ҽ���+{1� Y�ٵL&;�#���\��	�{s��R)� �����*��u7"��b?+��=F?���}��c̛0?���~v��*��0�zjQv�-�7H���!4����k�7F+ȧ��f�c����1�no����U�$����E�P�a�̻�4��l���ު�Q�}��G1��7OM0�p���[�\9�}��k����Ǭ�8f3Y�;V�<B�S���	��	I��:mw^�6-��!�6C�y�ߟ��&X�0ݲ�m�
�lK�B�	dltV�I�|8\O��r>�F�ͩ�e����wi���-�,���u ��!���23H4�R�={=dؔ��V�}��j�I�;��}}<��|ީ��];�M\�P����:Dғ�wLBg��ک�Ή��;�D�n^�LMM y��R)��4՞=)8��<^�G�ƪY���n��;��Ό�A��6㎬o^8F]C���I��m{�w��س���L��ܝ�I�֞}����X�f�1]*�ݓ;}�&�Ŧ��,X������9}��hu2��`'�Ny�tW�j�i�x�x)4Mn�M�*��/[�w��$Agh�`@x�o���	���χ:F�����J8j���F*z�|��bm�3�KkW-H}������D�����|��6'9����s��ay��6ɪLӽ]�Ri�e�|_Z�׹��l�g<ğd5n��_�ח�E���㧣)t5��/j�i��D8�r��Hd������Y_)ʒv<ę*�0�j��y���"]����@��y�:侲a��P%�Fm�|c�āsT���8Eށm���S�]Lv>A�����p���Al�&��\��C,}F+FD���,$S��d5��3VN��[�;�ϳ������+)����|���_|�� �;'ǻ�L�ۘ��}ޏ\�f-�n�z3�Ǽ�,pN�d(��>�lNŒ���{��;ܲ@[:$t{8\�뱏�s��W���ߔ�=��.��_�͹/w�h�ņ��ˎ�}�즵,�][�� ����1��y|�y�ܣ�&���uu*-�Nၡ\"�_>��l�z�D��Wþ渻��'ۑm��8ޘl� ���e����D����gU�fiƜ��O�4���	���"��L��:/��|ǆ7 @�DcL:O�0�Nn�֗%�p��ǡ�n=�셪���1L��n�Yix����;�ׇM  �cՆ�Ҳe�MYt��i�y\V�W�*U
YҘOx�yj9r�������{���ؚD�ƱB�I�e�,�Һ�
۬ S�� �O@N�s��ta��.�*�
gO1���^�YCv8�2o)Vn�u�qïK��æ>d��r�w�Mo�R��=+^҂^ج�SV��9�w\`�0Jbi#�s�#��K�ᯊ>K?^��\Gͅ)r\����\3��e�4�ӭP'hR���z�Y�4��������>G	�JT�<��άy�Ӷ��Z|��ėba��Ɉ�D[����x4>g`B�1+L+7F�VF-�
:�2��f/"�'�GpU�c����Fhvf�I��	���~��������`e\�!{��X��h#"9�ީY[���Bի��ԓ�յ)��HIu0��ͺ2ʳ�ƽ8ju����.��B����'�#T�u�Q��׀Kn������%�J�y8Y��>��gS�9{|SNf�_�ݖ��s&5W2au����#����&������v��@Nw���7��
�d�U��4���L�M��h��V�f���V+k���hxC�_y��y\�	����.R=�0�*Yt	T[h�1�	��ٻ"mm�t3'H����� ����#��l�%`mT��i�#���s]٢��e(9�Sj�j���rO]�4�5l�@׭<]����Mb�A�v2��x�4�������`��$�^�I�>�첹���A#���U�3�g�u�5����"w)ޒ��0�b�$�Ϸ��N�s�4��wv��V-wͦ7�����Dm�T��di'�|{�����c�ol�ZK��5��n������V��9�
�vH�푹Ҫ�h6�'����D�`T5q*s�f���f�ϲ�-�!�l>AT#k��rʯ{�4m�wf^��F���~UOwa���m�����7��q�#'� e�����M�����A��R{��dh��}D��D����\�E���V�e�n#�I�"��V�t��l���4_z{i@춵��le��C�;J�_!8E��OOb�4�"���Y�⬫X���
 ��3���vg�-�$�J���*;�A=ϧm@�ڤ��,ys�ۈ�߹r� �jhN:d\�z�uw�X�<�� 8�a.}�В�\��Oc<�E�s+k��p6G><�Q�	��� t���d4q�����������ٌA�ౣX���_������1IM����hn5\��>��]W��:�[�0-��>�@I����v���D�,t�]��4�؀遉�>���ʣ���+,:�l�~I?VI��⮈����q�(Ґ׻d;��qཱི�Y]�/�!_�s�j�j'���0`�e�1���t5�3���:h	�2|x��%�;��,��,����s[[�f���A���]�$�E"�t�z�&�.%���<���vn)���n��z���1��9k�;�pvu�*���I)T���z��cCd�-b�ݽ��6�ώELj��n˳]"9�o�Th$� ���:��`�Ɏsad���>~Z�
��m:sOp�t��њJ�3�=2�#g��[�f�QTw+4�h�~ёy��`��w���{��0��"�ގX/��)�Kf���{C��w��{I�%|�<��{��.�V�&��/_`ʞ���(�?TO�EgY�Nmu�Lؽ�o���^r�?�ڲ��7�%mˋ���Ɋ��7�v:�F^�u�D�ُn�Bَ��u3DZͮl�n����]Q�'Je��|�v�SOsw�Ba�#z|"̽��L���˃+:[��O_����p�H�%�>]�Y��-����T�o[�wy�;n�Nᵤ��&��rn�I^�O iA��³вy�f30�����*:�"7�i�U>�����x9+�>�����3���ԳzD�X�M]ni�ۮ�Q��^�� :�hF���;"�=@�ʯ;y�T��W�?h;�u�i?wj/j�g�,|�Z��3��In�6o�7]λ=�n��h�M�]Ƌ�ix��㢌��02�1���&ɤc5�T�[�7Os䃓Qǯ�%؄JG�Df�h�-��Nth�b<����ʩ�7�>�m�s��k�/�]��W���e��%oˮ�����{�����W��`�5F`��'��q�3��/�b�⒁����������f�t�=�=�b<=q}������O�]���O�{�zG;��<�b��|�`V��/�������Jrt�{�$��ÿ�Ә��� �$`K�UҝV�GKG'�����]�:z�E����\M����+h_��Z�4�Ɛ]��9��yj�թ]_w�U8,�$����@p��"���.�5��q
�"���&q뷢��#]��.A��kP�̝�y���9~��+xX�["JI�J�	�[6��6Y��|ַ����'�9&�)`ܷ]�����O�[���[����ƧhGx��'c4�b�W�y2�2�[!�
s>� F2\E,l�b�b�s��@q��}%a��WIG�q!�Z_gǧ����
�{���=�t3tb�p�5�����P�J���t�y.�:]O��5���l6Ձ�°�g��j�n���-/�Q��FE�����gq��w�����~5\��s��J�ai��1C�u�v*�ҧK$.Փ�[��z}>�O����������~=�������߾������#����X��g�e�`U�[�8�Oy3��c�/<������OcO:���_))�\+B��?{]}y������T*��B���(�k�n�����+�jl��`����Y���X�ǽ�����i�e�ރ��.�<�p�vs��޼:��;<�4�:�(�%���[{{��quf�\�(In@�N��l��'.�D�2��B�8��(���GZ��?w��t�r��T�{enp"F����ޑ��U~;G1��z	�dZn�Q|6�6��[ �[{·u)1�.����i����f��x:��6BnDyf~��Sׯ��u��9�n���b�;3��U�c{����w
�6���j������Gr1��� ܃AR�&�Op��^�s�ȅ�C]�pb�}r�Dڴ@�D�i��L[��J���ʇ���+�M�;TΫn:�k�C�Ƕ�{����1�$8ｻ�9F{=��53��L�O1�#�͝m��n%���i�*�j�J��.[yN���c۝�j�/� JI>�gx
�]���6��r�A�:4e��*��Y �s:n朒-�hK�8a�{����;D9�=���jucö�Ob�j�B��ۏ��-t(t
�E���'�y&C]�A�-1b�#0��ʶ�@���m�Mw��7E�y������
����}���.|K��0B�-&�y;�%x��W�S��׬�g�!�,�8@q�pn�C�V&=����$l+۱�o�-�74h�;U^r��{|���r]�giԮJ(�!�*ە4���wuhUͭy][j�ǃ�p�([��esY���EK(��/�"��J^��}r)�T�~��o� K�Е���N%f�]k�.�.�v���o����=�Mԇ�=`��yR}����*m�z����ن��+1؊kݭ�,JqD�c�:��[hZ�A�kq��;�{ha�.�*�}�b�nc�տޘ�� 5gi]y���>��xT�����b���΄F��]Yh}u�)�mh�Į��N4l.TE�)ϭ�O9�{e�6�<;H�����[�Oi��ƺS�b�àBT֝�y����x�/ޥW{]t,��-,BP)S�v1�J��hk�)��=/,��=X�h��$�mw]�*̣SVvh���Ty��zz}JQ�����'�+�{�a\)�Ny�L��o���ꯐӉH��s�μ�2��@l-�yv�	�i*Y��f̪�"��n��.�-�}@�z�-�z�wH`����)���呬��<�T\e��J�;fȴ���!�ٝ��EN8��-]c[����ec�doE�X_'%ѱHEg��C{^����{W�Nݪe�+m�R���P��%J�<�n1�]˩ bK���גnѢ�)1E���E�;���}wν{�����F�p;"�2Q�h�Szܓl�հ�sW)�8nbu��u'G+lQ�O�h�hګX�"*�[b�=�\�h�ӣ�s\��.F��7;�:��E�9��N�,Q��F#堹gMm��]�!l���9r9W%���9�W9�F�4�m������ːDscգl����$�&T���Q�3Q$5�kk�{��퍺�W!�:�
w3���ܜ��SMQjڤ,`*c��:���;[N�E�5͍�CNء�m�ېꗌh��S�4���(�4p�;��j���v�ѣF��X�usb;�ͣAI�SF+a�F����.���p���E:����m�A5k;h֮�9�Ѡ��e�ŭ��h�؞��*�Q�*�t�MU�(��4���UI��ړAI�-���::Ɲ.�u��U�������}|��^^�	:ܕ��.^�7[I�5�|5q��*
QA[�	O��̹fk��$ ��Q��ٗ���$���Z��B����{:�x�="=����9��q�=>��-G�;��'�ӿU�ݼ8[ӻ��nw{8<�J�s7\c'�7�Y�l1��g�^F^f��	U���66���t��E��'�d�G^ Lv	�4�0��T��*Ħ��U�x�,;K�j��Ļ�u���<IKa�Z���e�)���4��W3��: ��ly��n{7v�"'�Ǥr�'O&�����-�`�/w�N?d�优a���
�`���q1�+"��Q]xPBz�ᙬt
g]Ѻ"e?dqǚ�>�����SsN��,�B������Υ�5��1"މ�x�Zw�6�.�#r��K��gY~rG-���i�E�&�=���2��r�t�]�����C�܍�P&��u��n�L�ؑ8�C�q����f��/}����u���;e$���IT�}-t��zbnp�\�|��.|��ܩ�����,�c+7q��sh�L3wH:�;�y2��R�"�:���Fp[�?Nn���~u�o?{󠚧�Vq����r�"��OXn��m��:��3�:�<�޽�3�|��`�L���W:������&.|\�3�{w���4��f���m,�?���p=���/G�����"���@�[ݕ�."z&����"GgM�M~��}�eF���4Su,���:�Z�fݖzډ.��`~�)
��1/�;�������_�k�9\�Ǘ��dn,[NL�Fd��;�[���3�7���y�ޘ��ї3p��ڦ[�q�z�����q%�8J�Dܩ��X2����Y��S@��õ<U�=G;)�l$c%iJb�����;^&8�!��sS��V�oN�DMnSw�RW�:�[G�[���xBd��UF/�{��I�3�e^�]��2몁DП/pJ���K0em �"x��T#e�WKN���ͽ�x�]
Z���C �EsrK#�(�׶ހ".����CB�;��v�\��Պ�O�-���S�,�:#�'�7��������|��������f�-�<,�0gV���e�%8���{���*����}�ۏ�����x����U��:<���O�t�Y[���Z�8h�r�@��ÂF5+q</ww��|d��#Y�76
��¾�G�K���=��z-�p�)�U��m=�E�v��L��$�#�5�֑�jn�F�?��a�ػ՗��5En��x��;j���()�(��=k�̛�}�}�CNFU]��3��y��gдӗdt
F���JL�;VD��y���3����[g��D�z�g�	B	[����G�i�{�����x˸0,������@�8�$eә���E�w�B_��mX/��zRMΟr��S8~�s���`�t]�Yg$wr�'��}��B���6"*�r*��rH�4Mj�.���ބ�r,�s��ʞ��\�Ñ^�y�ж,9�#{+{��8TtvF�+�3\u��3�.���Y�8�kC��+~�s����ӧ���9�U�O?);�&��]�{�&S��T����݆f�\�w=�q5���j+Ǆ  X���;�F�NJ�	�e�U�g[���+y�{=K��׎���C�҈�άSwiEהz�w�]�\�<�à�]�lTy��R�4wt�
@^%�1/ޔ��'�����������,k��g��ޱQԦ���æﻣK-oBD��af����K�w!�|�Ϩ/m�;z��l3�3vOv���|*��́�~�j5ç��dYG�l'�����S���<�ƪY�26|���ɖK*��gU�|� wxk+C;�Ȕ�a�35�TW1�|xj�	-E�c�ҁ��}	'���M;��C��=/[Y��ydFx��Pi��[k����`���i�]�o�č������eD�����!�|���TD�*�	��Z����G4�l��y,���5�vĎ`;U*�mu��<��z�����bCIw�OYx�y�zĹ�L�:��w��ܕ��Y^�c36D�����深�����UC�2GM<	�pA��]�B+s�'�kf�F�EN�ۍԟ8�Db���Һ��L���Yt�2$[���Bh�fm;�[e�W-��;��2�݂��a��U�y2�3���j�23# �g����f��s*�ۚ*��9�|�G�m��v�AY.�%ca��u5j8u�Ó�{)���ݜ�ڔ��t���s&��{��oK���ܖUv�Z�,���m[���p��7������\�ڷ�8�0��]��0mn�-�s�c���� Kم�ǅH�黲����3��=�1� �o����+��и�6�!i}����Sˮ,b���Y3��q�C������3�/��A�GB]����"��$����{���>zi�5;����J�ѳ�9ܹW�wz��1�a-���Y��[�7%*�e��-��3c�����@Nv��4�:Y[/z*/jvEG��rsT��˩9�i)�3e�=�9����1`���bw{Yv��	ɨc������Ѹ�~��z2|;�dv�5�O�;�����¿��#�����ӿ���o�����Qg7J�I#�A1��4ۙ��;�m3��*6'4�]�}3{xT��e����ז���'�#�c�e��Y�\�b��[�����=0��"�?�lG��dE��ں�����"+�o*"����b\�n�ތ�9s¯eW/tS�����rhD�V=_����}>���š)���ڎql�-'|��4�A��|�w�!A�X���!�?P���Ǘ8�'{�^v�|V����e?�D�@�2b<�^�n�{h]�7gl�)�����,�{l���	���w�Iu"�	�ً�:�wے��-T�K�� #��e���)���i����6��o/�4�@�%����p��������r�-�"iS�s��\�9������F�Uh4�E[:�,�)�s"f��r��la	)	w�s�>]��IJ�ҦګL�M4�>S�,ٜۇ0�Zn�-@. �#lDV��I��)������V��D՚��;{i�ZZH�8T+�����Q\Z=�<�5�E �%�!�rC6&@���ܚ�������c�)�8n$F�Z��U��y���̭�YU�FҝjM�5S8�䌮O�����0��
=�6(,���������y�<��fb��ǌI��wd\@���ހ�z<�lD�6;���͚�?F�Q?8W���'�P���]��4�����#�oVO4�ݦ���w�����3�ʄ�-��\�n��x��)���c�6ϛ�鈸-
|��>ӏ��2�Y���[�#:��{�祥�{h3�~�e���
��珹z�ו�q���l`!u�u��~Q����L���7VS�<�{<c�'��a�&m���p��Iv7�3}t�����+�
Z�[տ3������nzs��L�]J�N>�o�c�S<|�!����-ʥ�H��0n�L`�k?}�OO��N�Oޓ�RSF��)�/�ߺ���e���"zd1.�Öo�
�F�U�6���'|�2'T[%u��}Lt�E��h��lS�!��WC�*����c���rʚW�(�����>MH��⺼�  ܋G�)Hا3�{N����X���+^&"�c�{]g�␮C�q�h���6��+�g��R�ڔn9�8�<���OE��=�AbE�j����{2}sN`l;��[�6bYY���$p�8!\��j�����E~�߈��d��{at��H�e�������h#�
�EH�n�a|�d��;@f�X����{k�&%�V~�=���[�t���A���e6���ޭfy��M�ț��]��K���V�ƃl��˨�21��B��Y��O���w�)=�l	�Ly������íf����2\HP �6�ݤ�ݽ_���-��g���[��h1g�QZ����Ю�Gv����E-��#�	�����-*����v�����1}M�,�I�m���>�&��,�Ge����P�Y��~�)�����O1�9��岧���>-RŞ:*��23�Oc��t��J2d���֑��]һ�e�ζ��^�sY�iNp8ݘ���a{�����F��uG��{�s?O��LӾ�����=���{�����Z��h ��8H�wfᕡ�]^O�(�N7sy�zƛ
Y���Ta��7p����6�t{}�p]~�F���;6Q�x�3;���	/F��~��/j�_�����`ih9�hA�� ����{t��$C��d�q{��[�2�������|$n��Ė�tQ��02�0_/{��;�4�4O��V$g�ȷ���ެ?8�{����;F�-���k�h*$��qީ��fg�j��F�M]VfDv�|A��'�.*�Nk|�j6�,�z��O��єS�O<]�p2b�%�/�3EI���A��?�.|�>�+ʱ��G7왢�J"���^�|"���ƎWh�P�_L�&�]�Yb�GI̙W��<I MEѝj��f��H�����dl\�M�S�M�AL���K-J�n�鳅�(�o�ݚ㛗��[2b���s��������t��h��ځQ/z��+���= ,�hd���B�F�vvJ����Oe�W?d^N=;B;�^=�#��&���("��'S��h�E�N3�/�/g�x<U�iW�P�Ew��T-N庐;2�p�wL�C[��6�\��.�x���+zlq#�)s�H�l���Ng2��Ts�F^���9����n8q|�r:�ԚŠWITzW�j2���==����^���Oq+�}�$�#���=W�Ux]n����c{� �>�lcn�9��\6m�L��g6S���oTl��N=u^�\��S�ﳩ�v����/���"ۧd�&�=���[f��.qڨ{��=ھW��-�,<��>�w�h��'�#�^W��W�] ��n�my���Eu3��y���ܽy�@T�Ы���M.͜]X{�+���y�>�8ha��i�{���)i\���ʚ������FxL�[ۻ�dz��C�J+�n^q-��dSk���W��.���:��<����ׇo�rd����m���Ҷ�%��N�k��Z�w�N���>Z��q]�4˾��"�[y ���ݽ��13�56ͻ��z���#�t��ȭ\hd����1��F�sU�R���5�j�ʌ�[��:�X�@x4�+	�׋��FF�&��j�:.�e[�鉹����ya������Ϡ�,�zJDm]u��r��l��̄)}�8���8�U.��/l�觏l5���rj'�-5�oS2��-�Q-�1�s�GM*��!]o����6�ni��W��ן��I�<$d>Dg����"�h���A�<��iJ�B7 �܁SNg�l�C�Dq��{����q�f����GGW:�A��|zG:
WB�JFUO�r6�\f[1�m�؎�����B�(f���]o�I�ƠI).�mR����s ��o͛�M��8�q�ܞ
[(�-6y$e{����M{4Z7���\A)?w�?I�����-��(F��Γ^Sh:<��>>?g���>3���~?�oooooo����L����G�44�vM�a���w�g��"��Okۅ������]�
�Ûû��4�%�ư-�(u��B�^�v��c��o>X�i��]�uÜ'�@7�ݚ�c�t��<z���<���J�cHxx��G.�e���r����`��a�e�v��. �k%����[E�	���K���ث��ܭv�@���U�Qs��DS�OrU�jF㖉o8a�E�*#F�������������vN�ȗc^�Dស+��=�61b][l�6���,^�����?���t��.��H�>���.j
9�چ\Z�a���^ػ��Ǽ��4��Ө�ͻ�þ��k1�)�t4�.L:�R��K����q�(@�$f�Ua|�xe>Fx��]�k��e��{|�����`�����w�#&�-9��~�W��`������H�w6i�n�^��:��'}�fz{��a6���/�T�X�3&��&�a���վXk%{C�͵0�og.��H_jЫ��*nP���#[�s�nffl���D]��g���'5����ͭ��nt3>�о!쭔̺X�YT�P�{Ow;���䟈��b�w�E�Tc�/��xl�r�����9�����j˛t��zfw�Kᢵ;�9�`�����	�n9<a�z�7H�c����򫰅��r�M�Z���s R�̕�9��=��u����u�� _�-C:;:E�2"D�Wm��F�&)�f^���	,P���Z�u
w��M����8�H�CS�{WE�-]3�e	\��� ��uv�ư>'�����a��z!�&~�o�X��>�j 1�zˑ��j�'V¼\u��q
~)vӌ��q�"OR�Rڢ��w^�S7�
��y������S|��XB\!�[3���#:��e���C�z��m��z»��2wYF<B^36�(�LK�b�6��b�/m���W�ե˵��]�}އx�U=+vu��<���0���P��V;j�:���o����6��ֳi�'Y7�t�ͤ�
 �՛F����"��s�n�SU�h���o�w�{3n����[g�m�{����WZ]�)��6��
��K�0)ѣ7��*��]��;f�j��)�&�ޗl���jEiՍh�rU�zJo,�̩�Uj��:Q}��Lݲh]�m��J]���TWj����\%Ts��-��7ǖ�Q��E�le<��Or������w5[�1b���s���FqR���D<���`��'�7]ޮ�'5���KE��!t����:�$܍a>�y�0/��#�n��Λ%��Azs��޶0V�[t��o��f���,�!�d��Fqx���*ܔ�6o]��X�l�5����ɩ�lV\e�q}SF������B\��p�F�zۘv��ni��j�L�uYoS���k��n*$�m R$GC��#�RSE%G
�U6���i*%��(�٤�r�ͶMumNd��N�kEU�֪�j(�)ֶ��6�h�Ss:����A�MPAE[m;��}`�l�Q����DT4܍1Sh��UZT�Q3QD�T��ԓQQVڈ�
� ��Um�(�6l�ƴ�D�D��y�US$ss����gk:��b*���4AA2L�����"�ZuL�L0S63O-����$����,�8��%�F��SUMQ5.�Vf�c��
"���:JH�0Qs<�I��j&Z�`�f�*""&"&�9�%�Q��Z"�52�0ͥ��0N1��mcI�Y����[gl)*�f+��(�1�Q��kPQED�ld�ѨӴ�$�&&�mSPQ�M���C% ��B�x@bE��2#q���rT��5e��a���
���]���z=��[�=�e�r>^��S2�D/4f<����-c�pT��Q�h�n0n�v��:�C�?�JQEc�6�4T�6���TA0¦�FAB�T0?�&���*>�"�����h��^2�<}'��A�3mUw+'�en+	>\����v��a]��6������"_a-���f��/#�T�0�:6�}���i��q�ޯ0ޅʻ�T�=؋�+�3����E�=��֨�[IS@*q�"�}J;�{�
��yWQ�KT��2�qO������`9] ��\c4���+ͱ��i��V��;u�Cȋ�0a\=�ߛ��N�m��x�FwƤE��1ګ��ޑ[���Ɛ6�>�8#�Y՗�K�F�Y�N�b8���Q�/go��t�����l��>8)N�?H�a/t.��%B:��=�٠���ۭszm�=�� �ȕHo"�YJv)�CX��S��|7>�۵]Ժ�0cxmk�{K�+���HׂG[6�K-e�FEʊ�5W�zt��
R���|f�P����-E����E�{���=�CR�"�g,�@k_��d�������*VW�qw�.����!=oj豵��ȭ��������F-�W���Y�b�5[�e�1��87�sW�;�3͸��cy{�%ñg\����g�h�ȓ&*o蚪;Ѫ�c�Qۘ`ه���9��t��un�PW";��X.ϵ�*�9�E*�=t��v.M�m�"��h�V}
�N�S��n7ˤt����sy�ݶ�x�[Hҫ�K�L� �R=��p�~)���S�C�gډ�k���hK��D�d^r��U��)��ُ�pB؅�Je����n,�݉���v��P�ky�V���\�e���=�����%'%��%$��_X�Ѧ��9c�>���3�/��rןu�f�]�c�v�c�%{ە5�xN�7��	.�0&(z��O�N�&�%>W��F���򵝍tU^�����&�������pQ��;�����θ5J��l]���_Eޮ���;A��6��\݈��e��v��{r^7>#l��As(�����N��Pjc���p-�H�]~�wY�wT%��8|�3��,���#d�Xn�֫}�_f.�ԄbbzE5z�#k� �+�v:��u�=���V��7R[{x�ܼD��x���8^��<������v��i�;� o،���h�B;�X���W���\tV'"��ꋦpj�d{$8��3X��'b������6���tQ��1��_���I@�Xn=?{S�]�<&��P/-�<$Di�崹�ʍIDT^my&��nM�s]T	������W��^�GU�)Q��N��de�[ټ��=Y,�
�K?�'�Uz@�=Q6z�b�r[W�@�;�dUL"��ǪU�i�<��.%��gA\b7	��F����C�K����m��<�B���=&�U@�d���� z��-���l�W"ڢ�SM�p{�p�)JO�0�$T�&����[���"�ݽ	o�E�ɼYѳ�ϒ� �m�ށ�	�rEX�g�2v�U9�Z;�L�Ŋxdn�4�d�f3�������p�jU_�+���q��ei}���!��*���;�s[�g]TzHa/�W�(?S�u��䧎.��p���w��;�0��F��O׀ށ,k�����efX
��<&T����we�κ����\�M���5���2�V"J������ҭ�k:Iba�UdӼ�a81%�_$mgJn�kШ���^X�RS��e��b+�Z%M�
�y��m��b�]�s]1��:k�Ԙ`������}[�^�����x{�;���e�r�d�^~0�G����vA��t�|�Flv����{�էd�%fL���q�DE������w���aWA� u7F��s8o[r�O{2�)-�_�]���e=��ؙ7>)\��'��}ϝ�p�p�� ��f���Ұ�f������Q�i���V��$�$vI1�Y���l�F��5�}���1ҩʨg9��Q�x���yo��$�׫���	�#{\*�ШǗ3�Y�A?Z����m�_H���)�,��v�kg����깬�"�`����见���ЂMw�"c�ʹ�S�Zr�m��wxl^��bAtd%�ה����:��=��&_�TB9�n61I	.F�c8�x��J�)T!+�w����=մz=�eL���E̎7����}�PӀ�XA�AK�x���(�Y�<f櫽���~���,�x�w5�iļ3}�c��.�3{�z�=u`S0��K���7T�6Y�%������:��0[Y���hV�K3u��	����W4������dy�d%��dɄ��֝d�����0�����;=����ؾ���<�]̂��R0��ګu׵.n�xw�'[�L4�1���*:؈��47�$��z. ��ͿS�ꮞ挹I��\��g)�[��@�gM���x͞K.��ΔN�����=s9e���v�M���:��j��'�ں��UX��|���i�]��@Ó�h��$L��?J2�y��t0���᭦1�k����N�Y��{T_O�J��eQ(��^tI;�mq�7��Un$tOv��h��Oٯ7wśNS�H8�2 �4#��~�4y-H��T�Eϲ��[�A���+��i��D�׈�C�S��ܑ{ԩ��l5��~��װv����_�}�s`�r�D�Ě��`>ّ�'p���<[���7=Iu������כoB����5��
�xF�T7F�}��7��g��c�zP��{��$�5���&���iY�a�H��
YW8師WD�_6;�؟懑�}���i+��ią���g�h᤮����(V��nA��c�'�s��w�{�5���hf�*�)�nn��՛��N*��>vk���>���n�&ƯM���{�
��&�3��%�j�/W{�������B7���	�XRח62Y�c�96$F�~��yñ��>j�t"T�x^�H\��\�q�u#�9���W��!��c�U�5�v�WE��!l��V��Tl�P�M�PR�:z�Z���o�_��\��)�ӄOW�W�B�x@]�n��@�a��R���N�A�7�k{*��n�ުs���@)���"��_.n�3U�Ul�����FNU��h��ISuuK�`t�~
ڢنݩ�	���W9˚��.D��T��7.8�=���	�3�6�.�:�����sm����z�����qռ�+QQD��a��,���{�T�7=殜��+We�H~�?�#�F�OU��^z�2�w.��Z��)I�w15[�'픠���U�\{�7�kI��a�{�v�jGdo���@�l0c���zx�=�T�d{}{](��:�\I �_�֤�m�޹���r�_/zm컾X$�;z62rrI�j���<o�ݛ�ڮL~�M�r�C9:��i�af�-X�=�&Ψa]�v�?Խ긥m]��Л���|c�>�<_cWG�rj�id��n�w�'�m���o��<�����h)��ǯ��3c�� �̜�wd�p�bWf�ڪ�/&nql��˩Yڪ�gc��N�m<��
�X!�vЍe��
_�ݧӊ��,��o���������2Lt��g�A�t2�Z�����`�x���\r�1�m[�$���j�|G	�p�>�:$��c�hi�e����y�#��陽��!��ϵ|lf��"Di�r�W����ҚK�%�y�4��OU���)X{�hD��{3+�*��BTA*�/�5�����ˮx.g=�r�&��z	7z�b�l�d���p�J��md��q��Oڷ9
]w�ߋ��=WQ.g:
�� �w�e�� �1}F!�b�b��me�9D���$�&���y�x�g���>�%C�w���6l�Zp,�]jo74��%k��uTe��RM䕥�&�*ݳ����yѝ��٭KS�K�LgfTY�U,R��SR��kZoqL����t59+VB�1}o�7}l]�s�b[y�gL����7�7�얛/;��28"H���mE+�J�)�2��Ů�KS���ma��M5�������hJ��b��f�DrE 	���D�f���޺��^��=�3}�����b�p��O����*��-�J�zW��n	���G��������1h~�(�t�a.B8�d.�u��䧼qt@��g5��P��5#8�[fl�EUN��ԅ7+�5�,m[���*��"�����2�\�k4�W�3:x�U���n�7�K�f��6��]A��U�d�T��b�"2�­Z��.�]��	�j�􍾦���G6� ����z�x8·�79|���~�6��NWtl��s�]�r5�`��j������@��Y�c�:�b1�M�ej㠙"@&�0h�t�/��A|����f;��^�l�;¾����,�£Q���p��{�op�;��&�8�j���y��U��	���Q 2p��*���g�P,�22ɰ[~���NY�c���zP��+po�A��vo�菏���:���W{y]9Z���etY�wafU����pV�p�nEG6�d:B.VV<�э��+�Z�������Sn>�T��	h�KC
���ex*5��o��!0�����{w_���5��j��jD���<�E���6�w@A&���]��-�W.���g�錎�!�h���oi�f���3�o-\K���:k��BgY]`��ͽn�3�;��@��7�d�Mrl��R2h=r��EM9i(nV�{Nk���o让�>#�T[wvw��aF|_�.��IJ�$��m�_^Ch��c�{��v&e��3��C+���Z�w�$���2E���x�G�͊7�W��s����]:�뀅��[^���:�g�=p`� �Ҿ�]1^6��;�
�h�gegl���f���ŸAb>�����vr�Jwu�=�ukG_lH���� �~�g����\�ŝ�{H���Kc�|
���{ro�j�'�oI;�<mt�`��޿�]������G���nH���=�nJ}	���]�TNb�'���*������'r����e�K�$/�I+˭xul렼��������ƕ��1����G\�\�5�{O��8��5ʱ����H܎ڴhf�ok����9��zn3l�oxٛ�鬜���~Ʌ|�&�}F��R��h�[A"jh*�z[���&�tC��$�ۮ�Os��8�f5�q�z�9[͆�(�c�#�x�j궻�g�S'w�0;�����x}�ߠx�$n���q��]I�yF��9�Q|.�����GPg��Gt{0�������N���1�p��]����$qcy�ðQ���u� A�
�Y����c:�x�񞽙����Պ��[^�5�=�MhO"�&�ּ�͖���I1f�u�ش��ت�e��עT���d�HO����H�G[6���0���K�{������/qz��m;,��]ow3�h�>b���Ap���=�Ĺ�|݌wn`��p���7t��3$\���`B��nx^.qʽ��M>��WL�n��l�<uX0����ً͝>�g�������M[@2���B*w�>��z�^^>^�p�{���w����z�^�w�����~r[�����'���f��ۡ:�F���b��e̫R=��Ai��rg�'��!��7�:T�,��ݽ�_���H8Ҿ^�bq_�+��.�7�}j ���[g9�����3^O-��dd9�|b|.�	F.��4�y�)j�\oB�w��Aێ��7:��z%�vyv�Ƚ����P�#��o�V�"x��)h4 �Y����q���aǠ�gx'3qp�L��@�੆��ι����*WHouj���`�Qd���v����N���,SV:N��)s���
�jps&1�Z�����Epܺ�]�wh�s��+�6�� ��o�(�]��"�F�L-h52n"�RÂu�W{���풌�+B�\��u9c�m�Vz��g	Ҭ
<�V���I#�Ν��z�㑜�e7Zz{5�{����
��bvM�,�9M�3���7Om�YG:D0��5���.s�zƞ��kw��L�je9�+��+e�
�އ�;)�]��C(T�ד6�K푿��e�>�8Q~sH�%%��Z=|d��w��e�W���Y�˺-6L_m^'}��������m�vپ�]����Iթ����·��bj����dUaJͳ�C��������s����Gc�pKt
�۹�uW&!ݷ>������4R�,��mVV9���Dm��T�:�su�n�A2ͪ#8��'��jrgdd3x�n��P�;���g��c�����`q�����
���[�j��K��w��I�w�	�A*�0�l�?Ӊh���V�]���ۊ�6'���5��Mr���i(9wd�9�j��c���G�����I��Y�q
%(�,^��=*C�;='7=;}�;&Y��=�U<}=/�c<�����F3��H��Pd�)�q� u��p��2��C:�T���U�o.ŝ�%����~:`W<��3//��%f-��&N�o�X�!�^n�i�FW����]gʦ�x��N^-�ۅ�<��$�վegۛ�ך��pL/��u�c�چxb�}�i��Mk~tnZskc�F�v�@�]ݹF�wh�H�=�T�/a��_F��ݪc���Qq(��o1� r��k+��6㷜C�:I�k�m5���k��d����\/o:)]�|ZWj����)|�N+��i�]�H[���SFs��R��T�՝��ofos��<��^g���!c�uu%�ya-�����U�wܻ�`�m���U�皷���KzǶ�f�.�t�n%J��Թq��B�귳B�����'��E�l���b���:u&�R���c̚ws�D�I��R�a�r�^�x�Gܳ�{|�+_���ïn��'��D������DI�A�dX�qݚ�Ʃ��tVO-��ϲ�|��b_e[Qѭ���d�Gg��f�Ӧa.K|X&*�ev��/7��Sv��X�����sc��+�)'U}�W#6�1E9�-�V�QPTZ��uUI��y[���Å\�+�� ���UMQ�QDQ\ƨ���	-�Q31<����*&��i��jֈ(���ٛM�sW#Mm�b�"��PZ1�LG6�*�(��劊��bi����������<�CUW,TQS�TkU1Dm�8�DTcf�

��D�5���4A\�)���LUW#Rm��w2pf�������Y�"k��T�IAL��$APsb"�Z4�X�qDDr3MLki�V�F�u�IDDQ	A5Ur�DQ\ê�5D�DUUL�Z�ws�qi��**�mE��&���L7#TTQ�TtF9i"i�d�G#14DN���NV�<�"u��a�G#�D̑�ELQQDr5S���rm���u��(�h���-�Q5�4��44m]q1s[�*��b���cRTĻj(��U�Z������Sm���Z�IF��L��mh�؈kK�&9h����IA �����{geOLNA�
��!6�3Z��:^��������-b�����˸'�Y�9&�b�w��c�7�y��p�+����7+
u\Ӽ9�{���%T�p:�֛��2���Wp�FBǽ���n;9���[�R�\Kl��WPG��x��[<��0�\Nj�l�#�	�l� V���S?�դ��il��|��E��6�kT;���X�K�K��xϠ�N�����}�UB��oQ���I�ʕ�ٯ���|6M:����)C��\dFΪ�4h97��<��۪��φ�#v6���N��ّk�L<���7���FDwf�u�i��v���b.;����(�,�Wu���h6�o���~�r�����LH�����u�׬�ϯ���|	�	���du1��8�{r����}��Z�+�4g^#-��)��f1.]è֐z8Op�$�:$�S�T��m�}�]r{�㮥��dy�t�Փ�j� <$Di��/H�7�SW��$���%�}k
��U�����h�xw-a�ӡ�;�'�jCg�S��J*A�l�,��ԩU�|~��Y��69s˩ƯR��F�r'AW;\:
�C�Dfg^��<w��cK��Df��B�I��Ϳ�f�Lwuǯ�	�j<�U���l��W�>X1B�=�5WTf@XH��
�����C³���W9��q�g`������F�c�J�z�g�����lּi�.�tt���t�*M�1꺉s8[},�Ns0��;�&D�3DL�c��J��nk�EΤ�R]��Q�`���}�h�gx�Qg\E5��a�Ndt*��`��#ս�RJ�c�	ę��kr�f(��d�*2n��>OU��H]��vۅ�ށ�a#a�"��L�L!Zn���6��ی�;6ޝ�
����p# 9]"�u�J��Z+$�и�n�f4|zg;��9|�{�r��}��=��\��_���f;�U횽"�4K��*x*&:#@ق7��{��K���,#��<���,�����H�`ע�8V�f��s�/M۾�{.�ĞTw&���{��q����a���V�Y*��UiͶ��xZi�nZ�N.8um\u��N����[{��oY1���JZ�c�qV���ed���-���L�T���X���[ܐbM�\���U�ay�/��kc-�Z{zK���\U7�aY�A�|]�x�\9{G���"���Ӳ�������S�Z06zgtTԵ4�c���k�U*�J�Y@�Jū��=MѾih�W|�y�gx������Z�ϗY��
F�~���2Gtl��3FC��M�����u�A��oX�}@x�����fV�4L�>$O�(��]a�D��눾���"�B�q=��/�c�
�z2���/-�&���57�z�n�)���>8�[�Q�/�|�1Yg�$�W=Q���r[,ʵ��}���w���ƈ���H��=���ЂP93�]FL�wmN����n�o6���H��;�o{

@WQ�R�j���4�a�4UE��&y�،�(A��@#Q��r��+�`<��f)N�g���H�[�_y��h�6�R��\�&��a|����ua)����������������˘j�߆Q�P��
#'Дu�[�w�$��#���y�5d��q��c��q�$״�7Am�օ�A�~������I�7��ěX������_��@�>�B�4z���5g��%���
��ò�����;nM�aE�>{Wm�I֧B�w`fǘ����&W�I@�}�P�ǋ���ڝ�͗[��Z|y�Y'	����;>$������[:�`�S�Em	��m�I�nJ8�)����L��|�'G��ŹJ)7I�,��}>b�)%�,9��W1z3��g��V�/���)�kbGuV�3���B3�����a@7�5V�+��n���B���k�.��J1�W�N�����&��=D��5%1���r)�p��Ô	��cM��R�� ǒ�H��,��E�^�����gz��a5MR}��`G8(.6���ܛީL�oZ�֍�(��[�o:/�4�U~{�H�!����z9��#���2��/������&�^;z��p/x�S(��r}�#�_O��8�g�C�c��Y�w~9-n�s���h�}��� b��$q^uȶ������u�b�V�sH�Y�:��8�.�eG^R�j���$�C�1��;�<�n-|/���4]M4;�h�^`Yߦ�s����T0A$�2�h���Pu��A�.��,��*h�y�D��{;�l��+��^ل|u�5]�s�cN⸕d�r�J��1��6��U����|f�=�iy����)�2��w\g�is��ez����,�A6nϐ���_���=������HMr�QK���F�A�P��h���N�gd�Y�c��(+�X��qAM�p��.!m{Ƞ��m���%��j�$�UN�ܹMݙ"�MAU���(���
�h�����ܶ���xٱIoJ��JUFd�Щ��d�9���m!|Z1d�h9�nS�`A�2\�9�h%QI)�?_]T(���j�����Vv�:�5ϒ�`�-��l��J�q���'�Q8g���lXm��z�uus��o��a@r/�8lm+SV��I���e���y=��N�Z�"L�w�?�v����[�a�ޑ�F����O)����Hǜ=U���Ǥǖ�=|ݯ��V�s�p6��Ͷ���Ϊ� Q�$�A��S�Ͷ����LfI���e�{�v�8#4����d��yi�֎�lǋh���?��
^�|��N1�O�>��pxR����+�{co��ߎ���u=���͊,�7����?��p��i�`XU~��Ϣ��m]<��ESԫf�p����݋��d�!O]�]ڌ깖 �ݷ۲@�m'��Մ�O��ch6ǵ�6���e�֢�gunvS�^5q��JBŲ�z���#�A1�h�A�{��V�<���3�{YU�U3�}nY�hǒ�����}�4ρ%�}��o�*2�B22�Z*z����("�����h��1ydD���Qq�.��5t��m�p��6��{��H�a<!E���WY��a#�N���Ze�n�Y'$����\�P�㕂{�|�Wfu[�Y�`��ꧫ�6zr�+fS8�2*�x6Ë��'\Y �Pu#�>=p*%��ǬA7��L�ߙ�z�{�7	:U�zG9�Ji)U�\���D����ƬU��+f:TV��=א)%:ah�V�[����ty"��5O���j�)8�O*�6�����^�q�ɂm�oG�`�~nH�h7��
fB��t�=�|�I��������?W�5.a���v_k�Oe����s�j���nG��j��Z(�b��>�U >��^!3�H�x�T�r\V/��R��=8f=�h����{��'�u�N�G��i����U��'j�7_T�ZʝgPFo_^��E�4�-)��M�N�1�#�r7@�2��OAHQvjQlո0Xɞ{�4jz.�s	u�ǌi��a��\Td��.��u��w�F[3]�{o�I���{��t�%�'K�P�q���+�V�0,��*v7ZW7��n(`Fk�}Rz~�����[~��y��lͼ�z���r6�b:o��;ךDrG�J`�+;�;�d�*�9��-�R�o_�iب�'ov4��75��3�=5�\�r�F��?VR1���*a1nxL�q��\k����v@M����u�^6N�'��5�z�9��c�Ц3[�7���͈�dj��3�\h�Ψ�e�6p�W��t�p�:7���yAr�7�qHP.Z
�k���3�Ba�)�zM�T�5����KOt���C�ǯ��Ǥr�$i�״��� �g;����zo�S�%��4_�"��-��`���*�w���Vt7��k��Yu
U�YDѭj��P��Uڎ<�Ѫ��-�P���;���te��Y{�GQNU�όuw�t�s�鉄�����<;���*WJsyS�]v��ݵ��j�_0�e�m�
�N���L��JN����q�|�n�c&�.|t��XPT�ĺ������+��>_��_�o{�����u%n#C&#8��y%BҕA�����V��u�~��]1ׅJ_AVtm�ɹH��D���΂��68ȩ_ov�k�=�uH�6�j�j<�b���"��%G���"=|L��э��I	z�WtFLeYm��0�H$�@>��V5�P����zxd��V`4I�3wb��i�����)\St�Y�#��C��
A�b��l�w8���sƉ�!$�B���[�upH���G���m��j����o��u�PE���3c�^�wg,� �bU�D�wd��+�l_6�ȇ�ٝ��6�Tz�8����Q�z@��T#�H�F�䶼�51�k4fy7s_=�T���Pdv׾$׊����t8ǆ�y�H�s�m�"�ҧ+c��j��Y���IVzoq�%e���hi����eg,���jK1�ܔve!��qm�|bs̉��>���3�'���M�d������W�Fd�����wv8����Wa��z�u�8F�*g9I�q��)M�OR4���0���a��6�[�c�|჊UW�1c������΂0l���:�e����Qq_RċO|����x�b�)�Rc1�C6�1b��&R��������?��COT��f�3���ڂi=^�}j0$O1᧚;���F�Ӗ���[�7�$�.�ιuz:������"'���U�\�VJv}����iq�*W�;�s_Z@�O����l|9�z��:�c%rBk��2�4]n�[�g�wι�Uw�o-�]��m��qA\XE��E��1qQ��*D��ǝ�މ=7yg`��H�/�Ӵ:z�ٗ���
�P����v��9����Ug>L��p9U��iL�i%*����܍Vꭜ�r+)7V2�Cy�=[�a�#J(�B/O��#���UI*���u>�SO&�Prd[~K�'x��V��r�z������R�ܸ�l�O.&���g���5/S�C�}7�;T�u�ᬱČ��v�V�iT{��S&�4v��c��w�ɣ�����|7�I�W������f=`�������9�����Ch�s�Awb{����7(��<(;�q%ۛs[�����#\�ܻ,�"�v󹮢@d��F�َn֦�ZJ��+�ܭ���Pl�ٞ3S���l֚m���\���-��oLB����/�b�Wb:�{�@Ezz��K�UNm!��ǀ]�[^z�؀�s.7:�G--�|������u������"����ޓ(̋Ѵ���|3`�y3MʰK^WDo[nv���,��WS�\�qc�{���v;hf�m��a�B���-��]��z��C,�Q̶{͔z�_eP$v�&:Nٞ��1�4��+��]�f���k��u�R�;�G���{��s;5�Xf��EΪ��{x��?lВX
��v�
#�/�<$�6�����"A���XM,��5���So�������]�G�X/
0�hЉ���fw��`MZyV�g�ڵ?FL�;�l�t8��8m̈j�<��}O�����K��#��
��������W��aA�TAQ7��p����st"�F`Y�	�f�@�`Y�f��`Y�	�fQ�dY�f�`Y�f�aY�	�fQ�`XdY�fE�V`Y�fE�F``XeY�f�`Y�fQ� �aY��`Y�f &�`Y�fU�E�FdY�f�dY�fQ�i�f�dY�fU�V`Y�fU�Q�a`Y�fU�FdY�fQ��@�`Y�fQ�V`Y�f =g�v0��E�F`Y�fA�d�f�i�f�dY�f�@�FaY�f��.`Y�fQ�V`Y�fE�`Y�`Y�fQ�@�`Y�fE�e��f &�aY�f�S�L�3�3�2&$�#0�3"̃0,�30�3̃2�3�#2�3L#0��3 ̋0��3 �#0³̨,Ȣ�L*�2 ��(  L(�2�� '��Q�  L���\�UVa 	� &Vd	�U� ` 	�U�UY� aUf �UY� &UVeUf �UY�U���
�0 ʪ̀2��  L�3̋0,�0,ʳ"�0,�3 "̣0/3��,��̫0,ȳ*�0,���̋0,��*̋2��3̀k�}����~�� ��B 
� '�������{�g��{~����4����3Cc������!�����l��o���~� ������QPW�I  
����p��02��'����p�O�C���
�~��<����q%�`��S�~����}t�?p~���W�eU! B�T(Q�VT@�
E@�U@�EV�U�d � !VD  	FV@�  H@@ �UY% �P�H  G�~���?w�?� E�AB����G� �������AA���t�?�{��pPW����������=���H����lvO�'g��~ ������������"�
�pW���H~�����g���
���~�ρ"�
� ������c��o�C}�N���i��vp��;� ��?����~��C���t� *���x�������ǳ������:���0? �����c�"A ~^?�~��8 U�@u�:>�i�AI���i���`�O��������>���{����
���}���2���������_���� *���z�}v�*
����|�;���������)���#�c)��8(���1#��|* R� J(T�*�	**%R*�J�(PJ���$��*�P!$� **T*H�)B�H"
z�ۻ�J���:rl�J�T�UVwqv�RB��$) ��Tɋf�A%�����6j�IV�k3kaK4��j ��MV�Q$V�Q`U)PBER�j�$I��dQUP��c�J�Y�iZҪ�FҰPIIP�l6���M[z�4��mV|  ���uӥwj�y^z���C��R����SN�*�]����X�v���v�:�KB���J�ŝ��S{���˦��v����P�!��UR��Щ�D��kP��6�  ;���(P�4(t9�a�zm���CF�xx���H�ё��D�{�p�(hhR;�o\>���:t��իVY�����e-[TV�Kݻݺi�v�k �eݭ�����םԫ�Lc@�BTT��`P�  s�𦚶U>���z��tC�7;m�UC{��ck�J���X��)���N�k½�Rm����3�P�N��ݽhQ��V=�����k�u�zh���s����E)T�P�  ���-���=wZi�.���:KF[m����os��vg$jkl��ݧ�҄A=u� �R�U�k�P�Ӝh�fٶ�NΪ��kD��Ҁ�RED�|  ��i@*�
V�^ۍ ����+
ي�jY@Udii;��F@fUE�P�Zd�S�&؂[%m���KY�   �
*���QT��զ�)m)@�8WF�H��P���Z�Y@Q�Lhf�c���-m��IS���M&���[�   v�*�C�ER��iq֔V�5�A�.�4 -I�U �kTY&}P :�up� 0{�P ���i��*��RB��   ��� ��� � �њ�]���� ;G. @=�� (v���  ;������  휽����J�����'Z��F�+�   ��  }�A� ��A��� zE��� =(<:` E�t W���� ۶�  �B= �	�4[V��0�U��J/�  3�}�Q��� �}�=  �*`( k6�  ;��{�AD��:���a@C��5�
^�
t > �~@e)R�h0�Oh�JJT�  ��<F��  E?�MC@ b�@  L�BaT� l�?�����~C�7�ݑ��.Mɯ��k��B�d��?Z��dy��y��� @���ן���cm�o{ccm���cm�o��m�o���6����cc�|�����W��q<�_�ͥI
W��%��9�Ȧe����*��GwU"����k�E�O����wծ�V�&.���H��	{{�V��w/XӉIE�7�;(8ԍ�}�nn�ـ��"�lnir�X�T��Ҹ%h۳KjFA �:������$��i`��X��rY���c�Zx!t^b C%��V��7o5at) Cn鿞����J�ީ��Y7�T�n�ą�EP��7q�t���5��f�[X>��z��bJ���a��o��-)�����I�I��v�e�6k�	�-`�U1��$�n�۶@v�(3/m�]<��E��ݡN��9S�|e�r1@<�j �%��[�G/�Sx��F��'���[W�!��b�QA�ҥh��g4E������ЅǏH�tJ��d��Zb����a֫	cٔ-ڦ�"�&VK҅��vQX�+6��˘�w�=4mJ����z�$���-�a�2`4wnc��P*�D���chًi�D͡�-9L �w/#a ڬ�r�3.���"����^0���a;�ʴh�i���;�����*�0����^��t�t��;b��R�b��Y�b
)�k��L(7�5��NT��
�j�ib�\)�Rأe�5�a4��b��*$E,߮�h�)���i��A{.�ݪ)�S
��&(�P���U�� �324�JD�e��r�ݴ�Z��
�҃j+@̔.�� "a��r�V�f�����X��� VM�a�Օ��V���姤��# �uv���������Xf�Q�4�(�d�qZU(� AQ'WXv�E��^Z��%ZT�j%'Y�V�y. �D�dmmQm�Ke(#LXd�N2�R�Yg\�*M��H3.�fުa�#�B�]M�õB�ǲEW �U)�nR��FtA�*��Wͭ��wB�ʲ�i-e'x �i�G���M���X�5#1j�-���&R��9p��g���-r��0t$��$��7mk9b�2Dһ;d�=W�w��`8�;��WX�66.���ѐ�+z����&�Zh�E6hnsZV  �Gtf(��o67+WWS��2E�����e��Y��R �7�n-hm��[Sn�vF �iEZY��hnd����,̬���`�W[pHQ�),Ȗ���y���N#Qf�����������;4�����	���#�74S�N��S���E�0��S/.*噴t���8�^:Pǡ�(8>[nmjz��Z��6��.�5f	jf�\�c3Y �I���}r�y��4�5�q;T��5�Mh����$��E�J�uЧw����PsZ�
X���]�μC��J�U�a�Q��,㽑��#z��<�����Z�(�dI�`!њX�)�K�bz��t^��4�z$6&:��"k�ذ�e�R�v�F2�FS��^:�� ,1�ٳ���I�9HP�&�TJ��:�[��U,����N
+f�w�"�bPM����
�2Q����IQ�.�'`iQ�z���s �52��M�Y�3*�,4�r���m��M��_M�*�����ʨ�����f�1!/(�l�U��Y�&�9�m�Z�6���{V۽���{*?^Y�7��[�w�VI�����~�1FڟZ�eR�w��
�b߉5���i[�tl����T֧�"�M-�`�U��ovԘ.s !%.Žדc7���I�IF���?�ٓ0��X�7
� �cvr6jlxTӮ���*�V��a����6ZI��C2�%ȱ��!�xUfC�� �SrS��RT��Jf��V��T$8|P�m݁̒��j��	�{�c!f�ڤ����hk�w.��$����JM�>U���5�H���[$�ll�������!�Q�)3�G&X.f��a��f�fI��Ϧ$�,"���+�J$.�L�D]��E���y@�i�w{�2,��i�&$"�.�bT�MgLf2���T�E姉]�K2�e^����S�
-:�ʍ����v��v��$N�}�^�Zj#�Hp�kM֪ZlhYt�=�`�B�H�{�z��g\x��0���J�	$�!yh��7u>k6Q��DAh��J��
�n8#�`E�j�퐆=��m�ڔ�遮�!�#;����}[�3vG H��OZ�V���9�H�^�h��`�фn&N;�r;�.��uy5m�#B^&���+X:�L���Kn��xĘ���Je��8��b��t��i7y�����J�=&ڢ���E����M����)�/P�J�Qb:�#���D���;*��q=�v�n
��]]�Xb�R���Z�[J��M�K
���VAb��@E��i�)��v����w��7@S�Skq��8�]5G�D��{dK�׻MV-ÕV��O5�2c�"/�����L�wO1:!��b��Ŏ�/t6[���sh9+v�"L+kke�5�>�uy��Lc����r�o4�%RPL0	Z+ WV�`;M��b�i7�w!�dY��p��$m9�Ј�CI�w��_��K48�0\F4^���5�FnT�XF�E��Q��Q���A��G>��Қ��ہ����ڸ�2��dնS�������I���P$4m�̣���6��G��#ԁ���C,�uxٖX@uN�G-҉�'1GD�{F���Z��FF(E�	5Q�u�@5��-�����x����1�E�˺�j�A�חn�bK
x�Zx6
�3nQ�z2�?����"�h; %f���$m��lBM��xZ�n!v���>�7`YOs�!V�����CwpS#�v9����`�����p�1��7	.�:�-���m^e����ѽ�J64��Ǹ�T꺈!1c{�&ib��KskM4��jK&ctpMp �#�� �ʂ�ӷ�ZH�}��!P�#�l(mAM��V���&�[�q�M��t����zj��\�y�L�1����N�ʓt��Lb�-YM��Х�a��'Z�E�V�6��F�KI��A ���ıXq��ַ��\�U��֦FЩoq�:1?���Х�t��E,�qlAQ��*�ܢ�f������E�Z6�k�{i�f��HIV��&ƹ�d)d4�6�4:B�H�N]=�5���6��ghĊ��{j݃����0_�e1�j�<b&C��,0(���CV�M�b$�s�����N����0����*�$�X�e�ph�C�a�eR�]��)�Պ$\�T���)i&qB���e J���t�F�ܭ�L�m���F�"���D���X�1�ن8D8��ʓ.�/RB3����zEdd�M���`�Ժ���ث`e�,TS/E-Ƈ��]oM�Ʃd�k��-�Q�@ �c콁+hz�wMJ��[E�~�`�m[D�DF;K)�1��T��H��uʔں1�2�(�aX^��F�L�bl��n�#[t����wu%;�%w�+aC�ӫ(��"����wD��Y�KN�=��](i�L�Ǩ�N:�(�Jh�wqMݫ9�6Q�)�B�b6��ǿ\9Nܻ%\lio�pV�]���؄�T.RܱO�j"�u,a��b�j�Ʌ����%lܫ.�n^:�xJ�DYu5c�6P��bY���#qLH$	�����n�~[z��Tn�DGSqiڳ���c�D�*Ģ¸�hU.��&'�&��9v�-�nU�V�wY*�ŴFd&d�)�oh`�a���{��E"/Z���mj��]�;a��ƮƯ1��Y����ibTӆ�h��B����[XqV�� �k�jh�͍^Z�hB8lw�n���TGi�A��y�fNӷSsd�5D��d�=׋4T�H1oz�틑�ÊQ���*Ӑ�<SY��v����X�јt��4�,�1`:�R�۬lm%y.���KpQrm3-4Vk����%д�y߱�i�����f�$��kl55��ĩXA�a�d�m��`�ۦ�"1K�&)�l��85�P7s1ꄍ�$p����4�!����\:��n��z��n�-ыq�d�[nE�M�ޠ��]Z�8����ز�A@*�m^�rҹo ���d�
�th�E�X�z���Cd�q,�"ҵ�fC�C+"���4���4$۫
�HT��ߠt�P�V�z��nF�Xpc��Ҹ�PIb�Y(ZYhk@�A2Np,7�dz/T
	5B��.aJ�iX��h��7��Y��D��sʻ�\��r�)�X���f�m�yV^k�!Q��ʼ��3�š�M���g3���'��f��wW�0I-��uꥻ�	L��vq�M�]DY�,�5\.�b<-����ه3&�d�^�M�WN�һ���N^�,�ҞClj�K�尷,���E`̶ޝ���
��1���l����,`%e�T&Bۤ��-��D1���7(��ѕdh�����0F�3hV��r�6ͬ
�'X[��QS2j�$�S��iQ���I��zF輔ʃ8�č�̳��*����<�0j�(�ݎ��]��c
��[@�4��`���cԲj��[���=��Cr0#�n�A[�k7>�a��xTt����s8�GL���L�+2��]���E/�,���ڟ0�SPh���75R=/-Zn9�X�ш���2"��uF=�;-9Q�w�X���b�]#�nƶĹN01m�6H��e��?j�U�� ׳�5��7t�T�]̲L��hB6�S'jn���9�r�Tq�Yt� ���#e�Y��l]=05���I��$Մ��-]
:&���'��9O)*�Tѯ ���L��V���F�A1�ˈ'�I�dj��a
V��K�!�3&զ���tL���U��,�09f��p��v�Ƃ�*ac,�Uzt�tPX����nP�Rmh���"۬5yu���2)e[a�#fl{Aa�n���5�5k.�2�(��h��&^�CYgA'7�E�sjm&�S,�IXU��Ʊ�CR\f���ɐ�IV��$�r�l@J�t�d:J�y+k/rc�����EGB{Z����hS�)\\���rj�j�T��!YX�n��bF��/
6íӸ�M�fK��66���������L�5�-"�mѥ�{�lԣr��k
�b@H�S)"��ڊ1�3o5j���$Ƭm��5w���t�&d���b���:�ZԱ&�T*1��ڵ$z$ZNP��4�Y!�:�R�e��wj�+h0�Y.k��SƝMYW�5�6�ܽoI�s�Q�
H���N��,8��y{j�(+�\�l����d�����%�t���6�L����bn�Jj#5��f� �:���a;��f���.V@��^�6^K���R�c�M�R8@S wY,JWo$�j���e���E���d'�t�:�m�V�qih�A`ɮ�2��kn*Ug4 �[6F�3t��8�H]ְ2���W�MR9u
�[,M�Z��4�����Z�5�y(��`jQ�ɍ;�`e�n�b�����:�dّ�;�G��P���R��c��Pb�K��[ج��J���	�BO*�@���v��/!R���)��-�����7F�8]��5,��5��7��&�`�
t� �Kͫ�+d�ƓW�ז]f��.���U,@�Q����wJ���wA�^ �^���U����ܰ�N� ��;�Ij��$�*9R�U�@�������aR�{"Eܽǁ�� U?��gp$���h�d}�1̅���1+׵�r���φ��4on�]fCɋu�P�:���ތE�ŸΏ�cU��4pӵ�HU��3+1��	��[7�o��GX���yz� 6ciP��������ÅGsf�K�B���1Y��U-��pֆ�b���bSn�bn�v��,!-��V��'S�5ysV��b�e�:�W�m=I+�z�3[��]���V���R�����A4�U'��	�X@cE����(�®�T��X�Bq�e�g3�V���ȅ�v�F��ݗA�����7�J�m�KXA�5�ǸcMޢo-F.��r�m8q�v�݂�K��S�!�u����������h	�#3*:ťQP��ۺ�ˣ�f�`ۚY �Y�(��ʉ�Gh%-�*%cD������Se�p�5k�����G)=����&���p-����J�Bܺڶ�6�ȅ��c�bhY�W��˱,��o�`M2X�Ȑ�Ǧ�M���˶��KM���(�< kҍZ�5�8�B��ЊS���aR��]j��za�u����V�Wr�i�*�^Y�0�/6���Ffހ�Lci(JN���v*�i��0վ&n$v�]���V��؝��Yu�_�f�M��UO�CU8���R�LSTO(�(Z�]��Ţ�2҇�$�u{a*�qe�ZDx�;�OCSpA*;�W�0кc(��U���X���U��*gK��U,�*���U��������O5\,�n���E�X����z��5аh�v�n�n�n����3����t�����LtՕ.'&�Ha�VM��0�[�-���s0�Eb`@��w���T�)���qV���ì����b�m�z�cS6�b��u�L�F�lj�GXc��J���VX��u�D��0�v��ɯ̉(�I����be���D�f�ksw���<��u.DbͻߤTn��L��)f���g�I�c6��/,���Kv���,B�ϬԱtQ���pL{�4��V�dK���X;u���k�I�֨.b(L-ݷAe�N�K"+�h���6�o�\��D���u�W%�)�rz�=�O3�RP��A �:	��X:�wkY��B�ѻ�X/]I|4�r؞�E�"���)+t��\��9��F/��㇒�����tKo���"
ؼ���.��$��s���Yj��h�;�9��)iK���nAє�=�o�jN�eZV�(��4"f-�t�Z����٬˽}�������yi��c��6Y�@�U ����� �K��N'Y����+A�N�wO1V�Q+M>��e�w/�M�^+e�ݙ,��NV��,T���*=c�p��� �'òQ�%���7Ł��ty�����,�fXJnkW����1��mlOo�����U��9�{����!�#x�x�]��)�٣5�Ӊ��T���D��)�������as��k2�e��8�I��}�N�p�Q��0�����j#�T9Iw�a[*���ڹ]�$͂=���uAwLh�ݓ_��B3١��,��h����1�}�F��_9Z�̩Itۡ�8W[X�G�F��v��ȄՙV��[��P�.4��<�7'���c2�Lr���������'��I�|�����8,Z��>�
�d��x^����9�
�R�H]	.�g\���|0���,�սHт�mD�	]Mm#���^D%�Tòc��wt���]ĵp7���%cs\�6Y㘩���e6D�V�#�9&3ݻ�1��c��h0>���G�:������vm�l"���ShpWfA�2vd.#��{��*�n�H��x;�}X[�9�����Kǚ�fP�
(f=���{d���v
BJ\����1�x�s��:���D��?#AZ8#1(�ᐬ�`)(�I��]r3h�ۻ2�9s��So�[�i؃�Ɠ;�,�n�o U+x�_D�)�}B���r�m�K��$y��������}s͗ޤ%�si��4��8�64(��`6+>�5.�/�����,�f�s]ӆm����z�**�����Ɏ�e��(�z$�\tX[/�3�#K�5��e��V�t��$�����Ӈ����	������w���&�&B��w�ؖ�j���jzk��G����:,�q���!���@E���_]�ҏa�Ҥ�s6�l���� K�i r�|�oW�����iц��o�M��^ �ˮ����j]s�"d�r��6"��#T�B��7�;K��S.�]��}:|s4�+�P��͸�\{v:vkeW[�����7�1b��"v���3�$x��&�k/X�(`w�Zӎ�g<�1�(8�L�&�⼘7�8[v�0V��SA�,�&J÷��/c[���Ц}n�[3>֭��R�7���R���w�qLW�=ܼuS�:,z(�Z�*:re��B�B���`I{[!��TG6�r�ޜ���m�Z̘�#t��ywVu&f�/nU��K-��}�X���c(��8�9K���aɴ�� ��C׉�ۀ%oq�v�&����BU���=��d-Uϱ
��X�[��ݽ<�JK� �L���i�٬�\Yn[\���*�뉹�;7i-�[�_Kz��
�r��+��7�/� ��~v��V�c�dæ3��%A�Ҥ�|8�nCM#�r�W
�dW�`u�S�x�8�uI�ea��&�lu��}�R���ҐY8�������n.Ꚛ����K	�Y�V`ď_��o`x�^Rkg���Z�)U�]����	���%o*j�^�ӯR�Nk[�u�����:��Z�q�8��^�[LQBr<��@˰�p�3&n掺4w��:�ݠ������H]Mt���S� r�s���2J�YZ��l� �z$���ԝ�)�3p	�dɜ�n��9CR�\��u��<b���(��H���Xˬ�P�]�n�Xv��k��"`�����LQ��pD|\��ν�[zi ���P�������C�k�j*�]�����{����!��Y�਴�3�l*93@�=��nV^v�ێe�Q�ͺ�e��Ǆ�\���J4e����Z����PT�m�Ֆ[��o[8nm 
��m���R�~�v��E����K��e���	��"w��D=+i����5f��5��`Q�I�Vd��J�Tܮ�nK�����u������|�a�Eng����O�w�:�4��>�>�s��P͂t9׫E��e�����5�'����}Rq�մ�(q��f�܊�׫2��V�"��9+h�'\�Z��LS}�3B��~	PٸU�7,�wqVۥ���Y[�ظ�Su�+i����X�"��j`�T8��/3o����܌�h�7�&����3�n��J��e�]VT]��5�
��`�ux��U�9��2�,�xFV��7��V�h���MNֵ�+M�;kw��.G��0��]1w���C9�a,=�Uw�^��I[}m0}Ee{{}�׺<f+��Hr,�4�n=�͸��^棖�a�C���ok�d����K��&G����]�{]-wƝ��]p6�౒�@Y��)c�^�N��Msu���N��W��%��2��}�&hF^	��͡Bi�k��&|��XKG�{L�Z�\Ά���Y5�̼B�R�E�Y���R;CCYl�1��2��o�܋7����+����j��V�*�7��Iæ��R���ᬗψ+�-t�Y�y���x��a"�i\�\����c�b	.o<��N8���ق�?N� ,ϋ�b%�1S
�eA��;����������ԾԲ=�:�4@�Mm�����Sc���8��*[�{�$��轭�"U�%����S�)��I�ww���XW��x]�3�P���+'Q�#����z�"Fx<��toP��.VJh�C���M&ج X�x$+z@h���a�c��<]�9A�gD��Mz�J=�tv־2\�P��co��Ġ�y��٥>B�������u�v���n�X�5$�}�{��I-ᕔk+�\ȇfK@��e���5K�RU����U֏PJ�쌼���-���5����Z��n)��j\]׌�	i��(^v+��"u�s����@U��h�1HV����Z�9Yv�uBU���i�Ng=�Gkfڬյ&�Y�
.'}r�2�"�ɼ�5� �vD�9W��!ΐTIк�,�9��,����چ:F��uv��Τ�����p�]1s�H�yk�)���Q�fj�Gf��JW�vn)(�����,Z�r��q17e�؄���>0�鼇D�51&�o@��c��Fd�I�;EǞe,�t��=�[F(,J��k��g:�7��+_��ַy1+{�kMt�E.W��[է��ijה�;��\�O-bƩ��7o��[���^-����te9��r��ݍ�}u����u|s��)���ԅ�9�^�k���y���r��r��cjM�V�5��:��<�R���P���6�\�U��^WL�������W�*�%�f�ݛ�����DGgh�ڷ.wR][]w��v�� .إ;�E�vi3 �x�u�h�LՎ�ӕ�ښ��pt� ��V.���m�1�	��|⮼ࢊ��2�N]m]�����n]���w9l�_Nqn����d�v�#z��S��+�ee�XU�<1���ÍMxNլ_=�z�]�zl��w[�Zhurڇ���x�y9n�ν*%���d�� [�o�@��҇c��W�gP+C�����ܾ̺!p-۸��I��iջ��i���L��d�q��%��I��"�OVo5���a���eؖ�ͼ�ZtҒ��eE.2���N+�}�zo��.;��Hv&�$��D��v�������=װ	�B�p�u�9���d芳Ե��8�r ��y�V��Z����%�fL��n��r����/��EM7[w�w���R�v�Y3�����ǆ.5�S��3C���Rb����)1�nQX�f��z(��ݡǐh�y�Zf�W�Okh�Fe����Q�[��^JW���>T�ٴH�ή}	s;rм���f��nV��L��
�vd��M�9��tV�p�փ5t��/���5EE3�m�=���9S-r��u���p�X)WY��M�T�c���p\bS�{��
���U��_k�Z��vM�y� ��fD��|(Y�0��7��#�:�E��\6N��m�tn^�XVtz��S��g^4���;�Y�J��}x&�N@�+�r�GF� ����^.�I]ema{����Z�/\U}ib�M	G�;)���̿V�K�Ai�QF.,f�z��L|��z��J����_��潮����wM���n�2�4�#X���Y.�vO��qֺz{'v���#bj��@޴7@ă�0�U)��n���V[x�JrwB�ܾpa8��/�1��Q@
����s���E�o�	M,�(��.�_^Iʣ�KC(ڃkq���owni�+�p���^�@�^�e��e��m��jZ��c)G��0Su�MH�qI��][ ��Vf#��8��f�fo*Gu;6u��r�PZ6�_w}����u7eK���>R���F���c���aC+ɴ�7k���U�0����q�݄*�a,��5z;���XUA���Wӄ���E[��I��
�2�Gg�\Z՘h�x�̛�h�%E	���=������߮�9����ir'z��O�v�C7�(ޡ�W^�6��!�������f�Ҿ�G/2�17d\=���lM��O�Ӟ���Zi��/���B�fAG(ܵW/6חK�zg_��Mn륨HWc
}�&̃j^��힎��(�'S�K�X��'9b��vr}�FwGt�v]ң�<��/%�Nk�֬�2�;����t��JN�^?y�0�s2L�=Z� ��c4�uv�Ԡ���P��u9,���	V�鳀-ښ�����ڠ�|C�f�&)�k�*����F+5�-�X2tu�i�BV
�#����]�eb��JU�/-Y'�}Us��=w*kH�qt��;	�ÂW���[娩J�q{ n�rݑ5 �Z���(���N�wl?wVW)��u�beq�VL�U��%u,�{�ڰ:�jS�K�n���wk<���~�.-��;�:]͋��MO��q <��^��!V���ni}�:�l)���kR�WYz_t�3sA���X[���G.�nw#�h��2Ŵފ����ݻv��(9m�;�Z��pL�](g[S�`E�8���[�:m�E������g$��d����K���yə��R���Ы�Y�s^Rf����*)R��Փm#�|',f�Xu�l�����`b�li/�{7��}��w����T����i�(쥘�G�E�7,Ģ�6.0%Ng���fANI��+��I֕A�B�u6�]�a`�Ojb��/�MC <�=��2Q
&��b�1�iը�45:���Y�:̮]V��#����s1��s��㡘�$dˍ+A�1�gM��a���3-�D���'ɮ��R�����'=̴;,n�?gP3]�x���b�G�C�Z���H�in�L�9��y�-_XyL�!�]oN�t(�&֋�͇vQ���=̃g`C�fR�W�����/���:���z���++R�����N9K��y���{&T�|F�v��O`��s&���-�Ѣ���I���x��=����(��pY��M��I<<�9|�2�ūN[s���αnV5�;���d+V��ڮ&�"�/��}Z駗N�����G�];�tJ |g� �u��R������a�tL����[��6D���]e:ٺ�T!��癝��y�4�+���)�$x��ɕ�eL��N5l�}ʉcifD����%gϩI��s�H�z��Xw�jXGԁF��kt��*�UJ" ��o{�eD0j�X@�X�S���e��*)vz�G���XR4%�F�
��7���g7�TВ7�x������H�rc������*Hսe�uv�&]qS�i����')�!���2.'-�A�+B���>K��I��(HtV?��[���Y8�#��X�(f�]�^�Ȉv��W�X�+{E3{)s����Y�� )���:X���F�}��3v�vRU�|�M\z��>�Zy�oLr����������}�}��ʵ}[�c;�:d���Y�)Ր��E���I�*�q`Л��L�\37�(���lel�o��׎�k�.T2�lr_=��5�`Qz����X^;��M�:�p��"�h�̠3Mu���R�S+�wv�f;�/�U�/�{2�wV]�Ch��aN;nJo�����aQך�7�2��䤩�/Q��Y'ou�.:4�.�\�*��<o�o�0˫�;)������+]��v'�s`���%C�0�Ζ�����f�f���OA��'�V�_9>9u/��^ͪ	=%�ڧ�i��3c�4�~���W;��^�m%�
���N�Db.s��9+��aeb�S�ycV��]�fQ�o�On��oK�AЊ�]6�5����U��3�j�gS�͡y��@+���(��޶�Whb��Z' ]��Y$�1_n��,�R�)e���Q��t"�Z���(��hJ��n��^ygY��JP�oV|Ӫ����u�~���SU��Q�O����.�5;���޶`��K7W	X7W\_*��U�3O���9��l}۳p%"�-'�/����m�ԾDK�\�{��lHL��M��h�֢��)WZ*��D�堥8n:P�|��%] �嚩�G�n�]�C�;�
���=�<�wzV��Q�qԫ��S�c��sr.w.+�������o8)�����n�ޭT�R����·bZ�}��w#�U��1��>Z\�_\n�4Ύ�v�:x�J:�`{����qu��{���u��ΫE��4���ܾ �7��KTq��5M��[�/\w�{���ϳջ�b D��?L�� DB���j~g�����,���-�2�7�M{F]����$�L�������z�u��:h�T�)Ks:�8]�y�/�����kze袏 ����4V�b��+��fa�d��;�؏h����q�b�K{��K��Osn� ���nAQCC�vՀr�[hl=)�
��º�#[I&M���6mT�m6u�{f��YKp�Gbc[���ʹ��"�r�����W���)fN�nu*�}�2oܫH,�/�qMB���GKÑ�Hu��J���el[ip�Be.��2��:�v�>�ĶS�uM{n|���ǌ�C�`502>ᜡQj�G[�!��Y��F�;)�3�Һ��^B���q᳴����]���Υ|�ˬ�,��8Sa;}�.���(�KML�*_"g1yt�FZU�vV���h�`�f��45
;j�1�`7���p����(��;�u�d�Q��R��l�ۮUb���u8�|�&v���wW�1�e����i�!fhE98y�m�,L���
i����{�f�Q��v9{�Տ��6��M[l]n���5v����*��{�����弳f�o����Y����z+)rUU�.d7ύڻ=����zv^Œ��]ֻ{�������Ԝ{Z���Z;V��L0I��V���Y4�[v���_��x��X6�T)z����`�֕����/�gˆ�É��7s�A�غe���P墕-������`o�����a̜�u�v!w�G�dγ���O2N�w=�[����1��R��s"���z����&�`��R�Z)G��������ш��P%�RtF�Y�A�]yV�ڥ^��l껝]	�Y��+NT����ӽ%,�uLT���/�3le�AY���tvpV��@D��cIft�:pa����][YH-m^����z�e`gBX�d�5����7��n�IȐ{���ѕ0�,7�zExN�郰��j��R�%��M���D��2��k�C��v��(,�:��X���0K�i�605�tj�c@�����+r4�݂�͞�\�WR�����ݣ�	�x��u]�`Z�d3zi��껳-5�% �5��+��C�m���*2����v���*�[A�#�}��nq�aw� ��[8t,Q��q���}x'VLW�B��c���'��[��p�z����U=@��]ؑ���J���3Cl+����8�гlgV�Ey\Z�]�t�m�X�����VT�16��ۖud�����̎C`�n�.Y�SQI�bgl��d��bF�	�C�gR�r�Crn���"����U���W1��&�9Zzó���h50+�m�΂���u�^��9�6�G3�i<fRmL�'^WdW�|�#*n��:F�]BjP7C���̝�G�Oh��"�:�˹)m*�z"�Y�lq�\����Q�h�WM����M�)�hj���sZ��{&	�ۺ�Jh���e�H��a��[V�a�ǖ�,"+�����f�]�Ok���i��ô�O�u*�2�'jk���S6�qܶ��2� ��T�����>��E�D��sv�7� `G^e���m�o��7���;]st�lH�>��u���]�[�����8���}HWv�m�8�:����fp�M�ݸ��#���1K�N��p��v����GY�`���EU�&���q7�����5$5����9V���m��E䠻
�����b�w����x묕��� -��r�2���b��@dn�a�ڗ[�n7ڀ��z�*31V�{3#{�4���<&����b�]��4ٻ�S���C�b᣺-�>��n�Zh̢9[)���m1�2�)��Z�s�����yz�E����Ǽ����0�-��΋2��g��-׻f]��rR8'%֙�Z���.�Җ�շ�Ut0"�.+*�Pn�t�]ѣ�J<�;`'⸟Iv9���lyJƷN+��om:-of���S:C��@�g*���uG�b���c��p�Ř��84M�u�����9V;��t��*諚���
�׸E��X{�h��:�(��Q8k��|K̟fv�,nXsr���A�2e8e�۽?�{�>5;Z	��w1�W��د%X�]k��S���r�X��y`*m�2��#�SL;»;��R��#CtS\�އ�n���x��d��_I�իa��p&��Ym��Q��^NӠ�3�����k�-�"��<�f����T�S�\�������R��U}Rʟ�ܧ$���}�@V;���V����+��c��aЅ.uy���1���>*�M-^I7�a����ETS�mf���XK����#Ǫ�Q�Dk%W<Nh�:+չ�W�������YjV�p����&&���b�+��F=<VՂ�Vl��8�2axc�A�²�%q�q��󍷷�9Ɍ��h��Ȯw��{[�V�p��j���!�ʖs�m��O���c��^9��,)t�JBq4&�±T;n��rh=\�����m� �o,��rZ�r6QI���ea�֤Y��[
��:0�w���K�+S�����J��떽ߠ�[闥*�m̮֕��V�N��/���C�sUD
\0'�)�K�4q��Em\�[�N��p�ӚT��*r�n̶��ik���	|4�F.`���{z�v���9����l�q/sp��De*q��wǻ!��`Bu��cW���,�;t_:P�>3P͙N�N���g��8�����6� ���¥���s�d�;+_ ��I�0��hm�'p����PsF�3��e�a�#d\@�8g+9e_#R��:{�����<J]׫W)k���$�	�W�����2d���pJ6bw����GιRͥ�
�K����t�c���4lx�4-��<y-�g����V���WV_-�%�Xɻs���*
�	�	��y�Ù/o<�h�௖�H��A��g���cRRX�����-����= ^��}7������>�Ef>���
��Q�.
ӻ]Z<(:�m����F�GrV�SoP̮�{ϕ��T�O-*�Tڮ����ҍ��K<U x:��|�Ց�Y���S����fS�0�aK�:ʖ)�-TyJ}��v�x��iNe� �Ã�}���%�������]ힾ�͍��6���)�Y<�'3fk����h�W���\�����f�>tR�Χlh�+H��Y�y��o��P�q�"�oU�#�z�����T;,��@+��oz/�T�ۮwCC+p,հH4�]n� �aw5�R��M��OB����d����O�L��x��GJ�s w$sh�:���½�4�t�=���Y�St���+ȋ�����l^_ax�Vx�S<8'��0EqX���6Q��5��w���+��b�0&��� R�؞�M̛�~����xnD�Ux�Tv�`�\���Yd!�JN샘�8�7��me.���wq Q�U���Wt!�<W�+^9k�6V�؏"�� U��DXyغCp�J`Rʒ�r�һ�ͧ[0u@���������9����kѐ�n���V�{�}syx��DTX��W��SE� 7�֤�����jCsZ��vW�v-r�-� �x��J��qv]]�vS��l��Q�%�/�B��іmb���SE�u���FUٷ��tl#,���X�.e�a֬�ԍ�c��@�ZX.V��c�PVa��cy�K��;R,�c'���o����gH�E���1R@t���KCr�|~v�[g!��W�we�H���t�v�۠���A�SJ
�uJ�ȉ�8��@�Ot �����{��!�*0n��J�`�jس4%��a�kpX� ��bJM�k:�J[z��j��:0��aWY����~l�rA�� �×��y��^@$ķ.�7�`Q�����9�����-s�\�Z.I�Ve˦>1���m�i*!��u���Ul�.G�{%iʗ�l��2/&j��V��5>V�ܱ��t*� ,Ez��5xE�Q��U˃=f��P��֬}�h�y��]�q��=HX��D��,�F��%ǪR,�iذ���3��s6��0��:�&�]�M�i������[8J���b]�KΛHL�6Lj�����I8�s}����df�I��F[����RAn��q`��Q�M��:����������ĝ"���#�	�eCJKDm�>j���֞�h�n�)B��f3���)�]���J�^��j!*sVe���0�4��_�_B��x��@�'�/���E@ݲ��%�o5���}Fе��q7]sk�^z�Ø7����:�CvkM��039��&�j��]����l��p�ܴ&��\��j���	�+>�ˊ��og97X�l�Abگy�;��[�jJ��R��e=M��!r V��
����pVt���RKlW��bWj�)�zkYOi�wk�MǺu��+X����O39��Y�`��3�T����G.����#Q��{�K��Y�U����R]i*U-�I�x�^��+.��q����W�%�IQx[�����򒺟�>���K��Ud��wX�4 �.���7\�� �J)�x�u-�x�3c��w�tXr�4�g,�73�~*��_7�����J���k��K9�ĈLAS*5����/�65�|y�sh��V���]ݧ�{. ���Wf��L7�:e�jD*��ȴ(�=��WEF��@v�9�k���2�2�F�"���Aԗ�	Q"6ӗα�z��f��ܧ��*�R��M����t;��ƀ���B/Dh���G�N���ݓ���xv����Iv,n2�����u4�f�ƱU��Z]F�V���ЌZA�+;f�v�v����+��<�>d�p�̖�U{)�zJ-��Y�RE�J�q]@ֻf���wWN���k6�vN@v��iЅt7�M�WRm7Y\R`�����ĺ#�t�̾��T��do2�G�U]]�pQ}�)��ՉH/���Fk�rMi>�]��@�],�s�����yg|�b�+uZ�/1�Fn�f��܈9��y_�Fh���ޣV4���M�WJ���9���]%t��q^Ы}w��P
��̪}��;�x�AU��a�\�U�*�� ��v�`�q�7ucg�8���r5Vw%ŗ�Y��w�>�8ฝ��榛�|ms7��~���p[f�t�d�Y1tEuH��X�co�t�̮�%�qֲ��C��%��y�.>�A��Y�򎳁W.�1�.��C�=*L�N��}�z���a�'�(���7f�(�P-[	 2e"D�j��Q�����ooNw�����Wc06mVEt<p���!���#�3��.�љnsj�/7�UjO^$����u�tV���=����M+��3�?�o�u�氊k�b�q�fjܘ.ٜ.�v���\ȟ�b���'�N݄�.W4 ��V�'kJ/�����u��)R��a@Q�'�:�2��a���vf�VA�6}��t���pY%����^�K�;<Ģr�Sy7*�{V��v*��1�i����$\�h�mP�6�wvy|�N�C��+�t�<��$lLDsb��v����7 �Պ:�vr��	T�X"��/���k]mj��w,mc���Xw��ǅ�m�C9�vL��ݏ�.�ͅ�D�E�V�v��=p�~�P�BkZ0U��Q�W���,)+����96MZjIً/�;|�>c� ����h���4H�"�����kLE	�,t�|����9k'f\�/���J�V�朮�[�.�g���-��m�E��GV��`0�f8�A^�|+��}F�����B�5��(�Lne8g��������r��p�}E�:p��$���c/�E�"�w�.*n���;�c���aG
����)��c�Q���:��͈J��V#�����p-���qK�,����;GK&�^:�#��+{u�l�`uN�}А�B'Ry	];��P���u�op���Ļ2T���t�.Y�>�6���ԙ�r�ۅ�P�B��5�ر»{�0�����ǒ�ʓ����B�ʀ�HC���`�:�ފŸ�1f�]�)�R��6 �|�,��I8�6+��׺�Q�N�	��j�2�@󡇸��﻾��ja�g
4���HĲ�,h���J�t�Yǽ	Ou����an C2��WvmL۝�\�S��}1��;jw~��x��VnWo��w��LHE�Tq}c�h���wB��gz�f	r�����È,�^�/\W"�� >�'���\�oG,��:��싞������4��U�xhL��o%c�{Qr8�3��X�LJ�z�:u�׃��XW�V�:oy$�gK�������e��X��R�-�*�me̳�t��+��z���cL2�_#�ǭ��K�����Sj^*��z���yn%�N���s��l�vjq=AK�������#���fmfc:I��m�o[2y�&X0BC�c�y��[�Y܉���%ͫ�c��t���\��50z��׫5�e.�l>w��m�C�&���"�K5������"����z�ɛ�t�3z��i�T����MӴF�j��%oe�5Xs���k��vo4.����5�x�)�,��6h�ť��@t���s#k4t7w����˺����ᆶB��EN�P����W}i^^X����a/tN
4/j�h���Z{�9uҊ�m��T%r[Z��V�Qh�R���Δ�-�	P��J��cMܴ�̫-�u��8���Z�0ޭӡ�囖���>o��N�}�`�y�r�<6��اu�]������b��2��xG����oE}}����e#w��B�3\���p=ų7鷑�O�WXx+)��}[Yr�N[uR.�U��" ��;�T���~W�9ͅ�V՞�M�]D7�'Z�eY���������L[�������:W ��xjX��I6ڸ��CB����.�B|D�d�y/*�.�"돖��H�:k���b�n�v6��w��ۊ��vG+��WKX�zZ�8�M���P��+�0G�`vq�P�n�:��c%����;��#�yX�ѷ��+�8�;�35�5��>ˡ��3��4*��zp��ؕQ[�G0�V��,��ו�vG�
��p����v��>�i�1yP��������t'Wr��*�؊ug�t�^;:c1�,m=��/5rZ��X��W�܆<�X��M���{^�����|c��r%ù]�s�cB<RPI1���;�G�h�A�gS��V�EmZ�WC�Zb��3)�u�����U�����j>EUڬ̷���]��(gw_�"���u�&���*1L+��Dv�i�}1�)��O^��V�,]$�pڰ^�-�5ܯ����E�=�:��N-b�AosW��E�-��4���(�c�}x'wr����[�R4P��C��DpƩ��O�[���Z�u��޵�()��=B����;�s�=���u_�Y�D�.��u[�^,T�f[}�;��۪Ք��p�V�7����eɇ�Ed�)^��O�ٸ�)�P��դ�qi��ԛgWl���� bӹ��3$�����YfgAA*:Z�4K�,��NimDA���9�r�"2H���D��&r�JX%���G �ʎ�T�V��%ID�")R�XZ$p�Ԃ��)P��"���B��dZ�E�*Y����R\��
*�U̒����B����PJ%+9uhh%T�Q]D��:)EUp�9D$�(��P��QI��Ȧr���*�4��8��.t�0�&U��҈����¢U$�UG#�U'�TDUY� �"�:TDUY&M-RH�J$Y�2���\���L��pʒdD��r�d��"#H��Z4**(�Tp��Tf$L�G9Ȩ*�"���(�U��t�"*�TTT9ύ�x����_+Ǐ~��Eu�%YG��m	r�0��oR�Od��J�9}�:^ø��b���.�t6��ƻ�K��L�|12��>� TE��Y�P#,�5c�6�p��]"s6�f�G)i'M�H"$���{q,o+���9�xd�a��qd��Aa�w��,�A�tl�ۦ��g���HñƲ����́]Z{���������� �֔�\+B1p�-}Δ~6>�x�������\����ѵ�_�Z��!ԇ�7�����+�/�u
*����c(�~8���\�܇S��)J�����g�ˈ[LԮ.z�:��{�nE<g
zs뫲}3Ǘ;�]{�+ӵ1	�&��ύ:��߻�23�I��̦w��}�S��zl�.L]�����R���[�G�@O�4B�,O� %�dDR�!vO%=���)�S�U�ٛ��K �1}���Y��%� 5������!���3js��P�:�ݻ��O "��������~90U��ZR^�ޒ;YS(�]0f^GC���*n�\�BX�̮�ڗ.�F��%Z�+�O-$b�MV��XK}yb�&��7�Vx[���vJ�7�P��v�(`�A�en��\у����8<k���u闓פ�ŴX�~[ܦs͈a��Ui��v�'��K~�z����Qʷ>��*�v�[N���<J����6�+}c�Sq���i�*.���ki��$�h��p�e����s{�sR�ϝV#����P��K����W��~���p�t<]m7]]�j�{��5M%�P�q��q�:��+���3�)k�25[9���n���z�'��g�`:�z����r�/�"�����-�Q���aLZ�W`����3�.�1l�O�]G��3�+��Fm���h9-C$��T��E��OJx�W�3j�h�e�d�SL��wZ��z��)�TN았_�><9%�δ�z�0U���&}�z�O�nx=�΂�������>�0�l��j���3���!۔ɕP;�IξS&q
Iy^v��:�a��ʫ�Od�m�7R_]�-���yp���F3�s�&�ˀv��7��7� �s������˚i(f{*24k�,8*6�i1f��Ѱ�R��y�5מu~� �����&8�l��<�$��`�Ra��) ׮���)s��|�s1|�i�ͭ�}R&���<�&�C Ϛi�XNd��l�=��J*���'l*�����KUwp�]	5��F�+��ˉ��� �L��s�姕{��NY����%򔫱lٛ��t�?4/u{�B�9f���>�L{�pn�r�sk0�Y��]���x������K�k �υ'�{���.K��:)�C(sx�N�;��+q�T�,K�%�-��&I�Մ�]�f��Yְz��b4��:.%�]�tꑿ��!�q�.:��.xY�p��"�{�Ȯw_1Ⱦ1��8m�ܛ�"M"ty�KF��U�<�j�X��v��wgG9�ʠ�I�ퟵ�t��0V�缶纣(!^O�X�N�W�'�hyg�r^@��p��Z������G"�(�q�(�s�>��HfC���:�m~?0�h�nfD*G�ݕɿ<�D�fx	"�;0��S�7�$\�aY�ܷ�)z`B�T���>㤖�1��O3�/��X�s�����"Frټ_����JW��h�r��9Z�aq��x8q�+K���N�	�S%MG"N���u���qw�"�d�S݇��y���bC�䵼)C�z𸎙�3W+tW�����ƶ�⠥�Hbg�T��:7rmK�Zn��L3�+*o���_'�����p�-��%�#X��8���U��C��fu��/��ۅ5W�Y$8E��wK�z�Ha�1��vd�s��F�"��xd���IW���ߖ�kU�Ws��5����ѯ���z��"E�v���l���:�F�vB���W�Օ���y|���9�	���#)�t9��S����R9-)�gq��e2{���zqA�.Z�:���`U��nK�q��M<���-��NI:�GZ�s���A��k�0U<��������H��9'�/ K���E!��$�si�N;.�h2��]���~(圮�!�o[#&�����"��̢R��EԾ��=�z� Agي�s�
ߐ�-����������7)]+?G����%��04NÚ���OՐ��_ي��R���xhm0�Lc�	�Ԙ�W�V�nO�p0��W��h��Z�ɛ�����d��e���3�������X{�lܤ�[��ۣ���=����Y�s֙(��V��}��뵢a��jS,wM��S�7o��Q��8��GwO75p��q����e��A�g�S<"��V}�Յ�]|B��l�v\�\��Ţ_;�]᯸R�w������,>��}�eQZ�#KtȁT~����z3�|&�{D=Q3K7"o8��h���ǧ�#���Ĕ|���2���,�Z~ߊT��㞪�r�I.r��M�OU�m�T�����d��Pڈ�%U�L`�=;����ߢ����0�v5��;�YƯ*Kb5�GV�F�{lǕ�u5����nDފ�.���mՊT�[4&œP�Q�{�\�2��ݗLNH����Ma��/�J�O+0V�Wp�I��.r��v@Q3pgVr�ֶ�r���[J]�����FIt�����s0�i��玤^ÚFj�": ����"~���t�a�#6�2ҹ�9��p�k�\;;l�@9���3"��Q;pꙑJd�P�~S���V�.])]K7�)Dp�!ĝ��wT1�����S]l!�9j�0�W3_D�Ui����6'�����y����![�ߤ�\�1W�H;�Z�[=G�IS%�3,��\SuG�D�gz'�@���)T�Xˌ_�R�:kak���?&k��;�:Ury�Fh�3Ϻw�>�`�N��moG/MԠ���d��mI����?S9�{��J�탘�:�3���ԩ��<!4��n@rlH��Yv/Jٜ�p�r�F����j%5v��Y�:�9�C���e�-���W�F��N+Y[��\mFiB(7�Pa0��&En�����ˌ��Q������E�Yg��\1.q��n�odw��E���M����6������Q��B~�X����%�la�b�fD�u�n�3�J��(���Â�#����G�X�=D�oT�<G�\#,���cܘU��3�H:��m���	�GX�B�3v�&��#3$��
������w!c-Ğ�L�O���Bb�ħnR�����6�Uě�+�KR�f+��Z~�_,�h��ΐ�Va������bږh"R�?X�'D*�ഺ���-��	܈u[k{��ܸgNj�d��g����t��]��s��7T�%�!��V����S�4�b�j��9}�'>Rj�K���Dݢ�p�c�L��Ȝ�`�1<P$�L�&�t��^��:��^��7ׯw����YP(����ϝ�-��#�7�p��8����<�l�`�z�k�օ��7��_������]9�{�,p�pֻH�5'J���?eC�B
��A�'!�~}|5��D�E t��!��<��D,s�C�M_��ic[��^:��r#~Y�4�KWu����!��ha�(n�XM*[��z�G�����t�0T$ա�]"~�婢3-J��)�9�"$�W��}A���*7T��{���t�z�9_�V�j2k��,'9S�m�0&,�۴�LK h�c �T��t�~��Bdq�-��hs;GZ}k*V)�sL�ٖ�#�+*�-r���MT V�䚡��Nu�8D���j�6���Ņ���ݲ�mq���U�X���R���:4�
w�q�*����P��Ւ����V����p��֭"�	��H���E��˴F�1�VE�ċʖ�uuvNK*��%H8f�`ã���K���y1�9a}��:`�a��k���d��� �y��f�mcO��b-P}ﳽ���c_k�N�<)?g̚�.�n���zg�q�:'F��*]Zw��#':ҍ��A��;	�:Llf�l�lCT�#5:agѮ�_c�"��,Q���;;=��B��p��E�����p
�C�%���W��$�V��,)s��Cu���&�mqf�'���Nˉ����]_Te]H���N��fG��j*��)w��5��ol!��*sHUaMw{��9��FEi. ��ݛ��詾Ǣ^�F��ω�q.��u����3b����ƅڱ���^>ՒIC=���D�s���u��/�n�Σ��82r$�'G��r���yOyoL�S=W�8�a��P�ξW5���eb�;����Q��y01x��gZ+�}����[�Ov�嚩XEXic�76��qJb�\鏞�<-����j��|g�S��H�/#uU�vԪ,E�v�� �*�wj��o8H,�ca���_��l���k5(�S��Jf���"DiMp��5�`�&4��*��r۽Sf�����0��rj�V!c=�ҥp��o;IA1�Z�5�hj��U�}�Cf�zE������y@)�`�q=��$���z��C�:W!\�ݡzQ��n\�+�\�%�}��mܻ̈́����8����q��A�gO�y�tYQ�mGyx�(����`,p3���ۭ��@x{�φ��4E�y�	�k\�D�A�0�ݟP|�y+_<���k�Mř�3����q���|ߦʡ�Մ��d&���R�U$	@&xA3���&�e�Et�0�ts�[7�����ܛ����Ù�K�E��N$>40�)V�:�LMz���f���3�ͨ�՞�W��u�*A�%=�g�.�-��M`�`{�j�c˩4�vj`���c�d�6�rs��������9:[��O����\.���v��B�S5� �'�����MX�f�*��xv?u�5�S-�]W/��j����?T��7҄>Ϸ��2�X�j��[��W�u��ԙ�*=Ɛ�V���J�9ʗ�#jn{UB�,�9弍ҩ9A���ϻ�ˉ�k3+%�_.3::7?{/D����|5B��V:S���:�}�_����I����t��ʪc���ϢT�2��C��}�η��"��{��g�=��F�^�ܿ��/�%I������sfP
�MC�L�S�l�����#p$���хXi���ڤ��� ��ZM���lނ;<fF��[ϰ���mgz���g�����nE�x�o!B9p�Qhvo)�Sp��=�Pų�E0�!^ݤ&���ۈo@�V8�nN���:���m�d<���8\��D���܎I38��\�'��#�U��Ҡ������.��HE��g�>�R��6��"�܏6z���j�`��4�#�F�i��if/2�d�;�l�C�0�>wOv��{��S�-��(���To�t�r�5�qrKf؆Д���n����j��6�z���1�09k۞)����L)���|���n[5����Y:� =���/�*��q�{���FR��~�y�^��p��t�Ex�*��V;�#&:�����s�DLtǫ�t@�?����1��|�ul��#�P���kz�v|��f2͖�C��M���uLȥ2Q���OM��kqs%e�e/��$LD��4/�ul"�P_�����-Yf �J�k�f~hnp��۞։k,��ؗ��R]������А��&���z{G�i�49d���2[�*���*�y����X�"���uD�D�!i��WV�ȭ�ck6���-���Xn�5`Wo6��2]�Ѐ',/!����y��aX����g��O��u�p��,�f�Z3.��AK���j�/uv��.�bpK��v�S�Z:�*˛�n]C1�<�a��)h*�=��]�B���vKE79��/�
&��&�p��/C9�p��F�d!4��[cC���+.��
�έ��dj��U��t5�����۷���>9>9�N�:&ATm1�X�;�9��N	^%�b���ˈ0�h�����^X��Z�&�33=׺}T��-+�D�Ϸ�3q�j�ó�b�=<Mi�&7�k/r�;P��;����@_�+�~ai�nnR����2]+�#%�3��uc{�j0�!*x�c���\+�ڙ�����;�N'd.@xe���}7�}ޟ	��L���9�7,��|��W�|E|���ׅ�n5�C���TW�*'s>N>@w`H}�Ғ2+��g��h+�9����^+���]���V��i������ �����Q��F�z��aNM�����r��"�ae�;����蜭p&���ip{]qT����Z�a�9���w}�hƇN`#_f�֥o�Cֹv+�i��^P�L��ATV)��7�%���9��r�/��0��͍������N~��,p�pֻH�5'J������m�7r����1��q�3� �����El�5;��Z熎�M_��9��Ȇ븑GձLh*�������DnkY:�]
�{����	�J�0�l��x, ��W�.��ޜ����A�� �/W����s"���s�V��ҫ��`��K�t9}�V�Q��q�F�u���v���g^�w��L�z�\X��"��!r�l�]I��{�Z�]LK�'���̵�4�ç1��9O�����/j��4*��s�JJ���g3L�ℳy�e&� o����%�f��r��ސ�"��������ʛ@�C�4�{qf���5F<�
�����5�|�X�-5�
n�Ǎ���y-��R�ҡ\c�5غ�=h�#�L�Y��mn��d��[�d���´�F�|z�L���TS촃Q=Lwhno$�.R��û��XLmV� -gs�&��4X�D�$[��%W=$iyVr[�4EJ���v��0$���`t��l�Ǣ���ɭa�ŉ�.���=3GJv�Ss��/,�h�ŉ��Y�ϭ[�{nIѲ�v�'����vؼ
��5�6�;���G�������u�I��9Z��:��̭r������U�����������`}�AHA���U��uL�B�YaK����q�:E^+3B��(�i ��孳0����2k՝���l��sK��Ŵ2�М��%�M��{��Iw+9d����|\g�]��ԖȾ�rm�zL��P�Z�x�M\C��V�����^��Q���wx��#�
�R��U)]@��]i0L��V4t�k����%Џ�K�EΊt���%ZXm�͒�\싱d��7Qb�'sK'H@u`�z��,�TsA�s��o+
����&�z��:����Pk���el���	�	������e�����L!uۨ
É�u�0�\�bUX�>�O'���%��&�r �:���<�ѫ���j��t�+(钬��錵ע$NY�B��9)���﮺�7k�6�ƞ>ҩg\��l!��Y�e͙�b��5�(�9n�E%��!�Ջ�}J�Z�٭�SSt!X1�D��{9��'����V��c�Jj�,@9p�0��²��o��6s9Dٮ���`�)E��xYe�Y�2��Gz�r��'�ىb�]��Q������o�z�U�)(�\uc!��_&RZ�Q\��R��'2n� ]����ww�o3Gq��QT˗��dR��F���C�������q)X
46 ��
U�otB�����@��p�MX��%���+�\
���\NS�h��ƭ�'�myč�	^�~Y�-6���T���qs��6��g���Y�h�C0��<}kkZn�q�6�Yݹ�	�z�kF��T�a��Qx��!n�m4-i8^�� Ych���|̭�Gn%q%�����SJS-�sz�q�x��9� {�`әIS�ذ��Yl.�Q���]��:�KJK7�4�N�j�QWuӏF���LEj߸�*�g;��]�C݉"3�"�(�EU*\��s���2)0�Ŝ"��΂�QY���r�r3�r8��H�!jȈ�U��r(�,�Z�e'#�G�Q4��!2�"
�N��U&U\�.�(�N%G;)�*ʦ�ĹEÜ �B�s�sR�"�9E!��vQEp��*���\�UG*�*� ���jQQ ��U�r��9AE��U
���B�I,���A"����",��Z�g4*L3���"�Pp���� �*��E�r*���r*�(�:p�U�"�\�ѭ2���t�(����E�K���	%�t"��[C�jTQ�TED����jj�(*�#���MH�U�X�A\j��o���͌6Q�s�i�Tv��guK
����M=�⑩���o�>�^-�
:�X�{�z�^�ݯ���k�-�?��_P1�yN�c��L*��9$��&�|��eӿ?P�Q����Ʌ�#~Q�E�k$��!|�g�0(�������^s���$���m����F�/4�����n�b�G�>�DH ߿����	����~��Ǘ{v�z���=&xO;�=��]�ǐ������|�ݼtbw�x���~M�97�?8<;�}q��N��{�aW~M�t�����nBK�z�����""�|>`����_i��������]���~M��&�����O�M�	'|C���os�!�� }y���۝��S�s���
�\x:����ɯ0EMץ�{H)uQ��ޭwgl���B��C�s�>�����z�~���0��[���nBpy=}�c~C����߿vߓˉğ��~�7��P����r�������	������y��� !dV�H{\�K���`_m!��xv�zy������p>|x7�{}&���G�8�c��,�ΧE ��7�x=8��C���x����y������t�}��߸=>ݽ'8>3�[w�`����V��I��O<�sVDA'k��!�0���=Q�]�� |O;����󿝤������۷'*���<&���v��ߟz�N��z߾����&{����F��|w����ʸ ��1�Z��������#V.�Ѯ��}�O��xO	�'!����9�'�=��	�]�ǂ��q��&��92�On܇�����������{��7�'Nׯ�xp)�!'��~^��C�(���ٹ�(��bVڝ��t�^'�< |~��w�����&�����{�xW�������P������;����F�<&}C�����P�U�ǈ���I�����ߐ��G��H�F0���ʷ����d�3uR�	��F��N�O�#Hdn}���}_���_~��]��|HO��;þ;N>o��=�xw+��1ɿ;�M���x�xw���;����i�0����Q�G���7���k�4��w���6�W�I�$��~���	��w��w���ܜ��������~�������0�~v�Ǯ���L>�۽o�yW|v���i�=;xy��ף��v��O[ro�O�#�y���}��l��8�^S��
Sk�TY��"���Վ�\n�lK��jr�d�cn�j��n�pV:��ޔ�^Pa�$�!Vn�G��;�Wn
#d3�#u|�-�d�Fʈ8�o����2�YG��Z[�s��@X�K,V���	G����xﴫT���w��N�r�/�;��}B������<&�}���o4o9w��������O�<;�����O�9>��N}~��<;�~q��?���~C�aC�e�������pI���D��G��τ�z���ep�`#�xO�`��ⷤ��v��M��qYs�Bu�$��D�t�q 
�pI�7�ޝ�0����{����������v��з	�ў������@�(I��!��n�����z�?$�q��>?�7!'���x~;|Nq�~�ސ�z����������	z<~�~t��iޏ�{!����rn����ĝY[���������=�>��	��|���1;�<��yw��]��PzO9��&�@�(��>;���a�l�O}~���v��=wq�|�m�P�sqD@&4�/w�#HD([�zY{���y���i���>���}ꟴE�����{q���<����v�����&�'�=���<��N��w[s�< |�t�Q����G�i0�����.��&�XX��F����%}X��G=j�x���B.�NϰG��#�"1t�H��aC�����y~���;~�w�e������ ��]��tz���;zM�	�z�c��bM���xO�����O܀q��`h3 �F!?|}�ᦾ��8�;�鿅��0�>�H�#Hd#^�僝���?c�|���]����ߞ7�~w�9���ɾ!&���x�<F��'?���v<�{IĞq�����dC *� 2�F�<'�ٳyc���}߽w��_��90����V��]�� y�=��v�����z���/�������m�7�{y7������bw����<;�ra}�x���zqτ9_q� (��G�|�~�@���Et�{��oV�������۹�ܜ���9�:ۿX�W����Vﱽ!ɇϏ���U��ӽ����򟝽��I�{��S}B}���DDq�LE�r�b��蘭��#�q�\�_�e������.��Q���}����&��c��]���<���ߓ�r|q���]�>8�x����w�������q���Ǐ�I��|q��y@�����׎�}���TG�y�p>T��O�S�&�vY�y��b��߲�u^���`�v�{��RD�d��	�S�7}����D�5P-T�3[�5��q�)ýS�Z�>=3��6s�T	&n[��1E{�\�Y:�:诒t��\UȴVwH�Rf���`U��������OwTr���&"2�0"?7~�(�b8�B8�	��ޝ�}�����Å�]�<��='�J��	7���=8��ޣ�!�ܞ��h{O)��_G�;˿;�b,N$��Dx�����t��EW7}�Ҋ{[&�B�h�����>��;ǌI��v�ܞ��x�W�Hw�",�D@-x��x�1�!�zO�:w�C�xM�����X$G��C�����K7:~;Ou:��n�S��Y��q�
S1f��9��'���xWe<|��������۾�o��M��nN������۾G��}C�aT����ǟq�!����b&<bk |D��G�1��8�Ϲ���ɺyw�O?/P�#�� #��	"I07�y�/�����<������<!�{���������|eߝ�@�~��}�;������ߓ�O��<����Dc�/�qda��n�kڹ�9�^5�Y�l����1dB,��0LA�$��>��=��.?w�{v�ߐ�G�����8yǿ=���'o�}���x.�� }���\.N����bO���������o��9��G�r�m߷/:��ц��ن>�>��=&�!�90����?����q��c�Ą����)��o�w��<?��}Iޏ1�Ǆ��v��缡Ʌ~[y��DY ������1�!�o�����nm��vٲ~���b0�1�>�Sr�oi���\
o��y��Ǥ<{�N��+�9���:w��㟮�ׄ®�)����~���9���1HC�T`����林��^����ݹz�(�⟫�*��� (�/�#zC�~>�����ە��z��(�}v�����>;yM�	��xO
�S}�0s�ۓ�X<��:v�o���w�w�j�O�9w�iSw﷯?�y����'��y��j�OB"'ǌG�w�����o��0��}��c���G�xW~M?{C��߼��I��y?~�	;�ޱ�m�ۓxO;��bH��� ��iz��n}�5=ZP;WyW�O�ч��b�Jߏ���g�ɾ'���J�`da�ݛ"+P��i���Ő> |�������xw�}C����¸�Bq��������7���<��� xK����T_ӳ�҅d��IG'}s:X�s˾珊q]�T��h��i�oo�`lVLpY�v����+@X{Ƶ��׀��[%_7عMSʝ;�ԫu������e�P1��t7%���w�.H,��� N�!s���fMV���SW���y���
!�1���	�~�S�rnB@�x��~v����}�����;~t�o�_x�~B�m�|�\
o�y?}���o�_c~�ߓ}}8�~Nq�wbw���9����bQ#�k��J�w��#� �PxO�xL>-�	��o���!���<&~�c�G�������<wݯѼ!����}��ܮ��^�py@��~v���yw�i7�'�~�6��{���m�S�mf"���=D!c�D��ޏ��þ;U����{����j��~|9w;J���c�}�9�����bw���n��o��]�c�	��9ǽ��c»�i���z��I��e�Cs����Q�^Ugٲ�U&�b4�8�c�߽��6��ɿw�:v�R��&�����߯��v=��ޝ�=�����7�xM�99��<���S}Oi���7�Q���~w�=����0�y��2k�I�z�T������G��7����?ǃǴ'y=�v���7߿��y}�r������?>��wc�a_�y�~�'�ސ�z�}��xO�M��@�����x�;xM� ��/H�a���Y��s{.=���.7���_)��������~M������8���s�G��^>��2_c�c�?Eo��UAյ��F,7c2)D����z6�p���#'����|'�';e�z�C�\1����ũ�����أU3��SE�^��Mx�4�5�P�i�����/�+�uᗝ�߭uN��RJ�rOMެ4��ϒ���[�2G��#>7lW�5j�K���f�zi&����!�-�[���])y��˥o�[��r��N)g)	�Ć�b${4��\�	��z�G���T�����٭J`�6�+g,�S���mp7��GYa�p��<[�&�����汦��Q�u�Q��o,�2���,�uhV�s'�<���K�xdԮ�Z�]Au�vכ�nqoQ�����fg��ݽ	��UP�Dj��Ξ���YgP�Av�7����� �iIz[�D�'D�%���'z��J��+5�|�PF�F�֥o�5%���Cju�M�Ƭ^n�R�t>��d�u{w}�V��pO"�1�3�F*�g!ۯ��8Xkw�Rt�����)���W:�by���hٝ"�k�D��&J�C|��7�N�3�+�25\3�P���&6��r�wz�tF^�㓸�7Y�~F+�"�s�,&��|��OUh�_Wҳ�����h���
�4���:z�1p�`d�� ׎�h�f:���1�����2�fݼ�ܿbp1�9n�_��j2�:�M6�y� p�F0	�T��L@	�������@+�FM*9I���jor�xS4��}���BOo��5(�k�I���s��ɑ�RI�1�ϒ�<���':tN�pXb���{}��h}_N-�/���U�����ь�?2m� '��Yz���{t$�t^^���;@�� L\��xpO)�csepv��-�}�����V�m=�o�on5z�z�/s�W�+9Z#?t����f��Wv%L�[��-��K�#`n������Z�K���:[5��_�C�{%Ԯ�<7)m9��1kPoS�����Ƀӥޠ�㜖hg�J*9/8�y@sB�u��������x�%8�L���#����}A�@�z3o�W�( ���vU��q���@u��g�z�<1���VUʣv�tӍ�*�"�U���J�&/�{_��q�&�'0�n����V���^o�)U���y�g+t"��ɸ���0�<����.�tg��5Jc�[��KF�9*,����^���4�(���؄�T��<�U�Xd��Je���E��j��rtoײI����DsMn9�l���e��WLlu�c��t��s������ߟ�������
O���Q����=DtV ��^�׾7Sm�2���;c����`3�k2��#���W��4��#�u�8��(1?qd����$�E��-T�}�p�K�0����~S^k�Y�A]�0W�`B�eKN��ڃMj���Ƃw_���r۱�~��wv�	���@Vޑ����}]p�Ü��v�8����_:�&��S�����v-ͻ�/�}�2���=����y9"1�\kꄝ$r!��Վ~�*�wua5��Lkin"��!�72�C��S&���&F=7if�\���2h8�i0 �L1���9Ul'.�����}5aJ�=F���Q�6�y��	tI��C굪������/I=��*R�Ee`�|_n\���Y�䥝�\��K�±Z�=v.%k{?UW�}�V�w���x�@BF�z'�����t�oOMu�7�pa�l��ցP��!����uiݣY��yz�2����Uv�\t'���:����Ԙ���&Ә�uA��:��,��m;�U�ED��$�������f�˵Չ�~�/p�����x���#kmC�T26ܿ�7`_%�X/����[@�^']P�]�,���{fuף��V�P��Լ^� N��rg���b.1��ϥ�Kf��q�N��7B�Ø룷�'��Iq�]�6�ʡ�s0���V�$��&V����5Fg\���V.�:'��Nxh�<��;7�_ gr�+E8�UZD��G��Gc�Ҧ��N��[j��s�{�f0MH�&����X֥�Bח9;�[���t���+�ǵ]b\���1Je��[<���n��s�����O�������;�o� �xm]h��W�t
��U4�)�>c�^8:����X!t���\��ww'�R�dv#��pk"�]s(�fə3Ԃ't������ �žذ��0��U����u/���x��lN�OXg�(B�z�vY���S}�_����s-��4���[�yW��g'�&��"sh��ix���swk��\� �y��+&���ud`�9Su.���2]�.�@$��"���ʏ�pa^psW�>�>��T��a�*�$&ˇ��z��������4�)ũ-��#؆ȭ� W�8�b�K>[�ru���AѲ�3�A�O5%��{D-7�ީj���N�@j#�oٖ��N����i��0����cx��ڸ��,�S0�il����sH�B�B�'-�h��s�t�+x��Y�4^b{���L��Kz�vD*vٌ�se��f0Sn�u���S�/��*u]`5eU�p�k�$Dwژ���xe������*!��ȇ-Yg4�sa����z�����iR�>t�����%[�a��N�&��W���A�U!��^d�(��g\���k	�6~}�H��̰9�,���/IL� ��L=���Ϙ���.�;����Ջ�)+�nm�Urp0ܰ4��v�\��1���V>�4,7�h���{s���ئ<��-\�R;�cE}�u
�w|sS�������X{�\+Ffy@0\�*��Q9�ԮF�~ut�\u��x���<~#���ޭ~�x����T���n�P4Ƒ]d�FS�㣝�J@����8D0X���o�� PVwrY�����5�%�E���Է��Je�gܒ6/V��g����eƭ�;D�Ԭ��ݹ��T�ڜE����n�_��<΍ލ	]�Σ��f;�ۜ�������_U}�}Y���38a����5y!dq�ݝ�.�D�x���iz��
%Ҹb3�s���f855i,5�>��h�����1�s:u0B�>(TU�a�7�0���|̌�2ǗaK�E�~�n�	�ϒ��e�����g���=yӵ@$��ɽ�[�u����v�P����C�[ܷ>�[𮔼�xeҷ�܍����Y�Sك�)�k�"��w���X[0�k��w
9�¾!���c�\��|mS�삩!�JK�44�t����*��ݼ�yf�v�㬟4�k�S�CƠ$hM}�[�|Ԗ_!��p��h����oC3kS�m9�T0��P@��y�Ѳ����U����}5�8`�k]�v��em>�c��v���p-�Jy��,X	9��e�v<�v�j3�*1:��!�W���q����[��u�X'Bz�����t�@�~��	a ����NJ�8���+s�#��R7�:�zz�JQz�36p�/>&���Knp�㸑����5�� ��h���ڋ�y��u�P_U�M�rC�<Y�s��E�W���/+V��9mAUvJ\�ՠ�''`���m�ΫnEK�T��X�~�T�78K�y�w�oQ���WJ��+����"�P��I9O��L�I귔�o�/�N�F�֨^�q�������V^]7|�u�ó��U�}�(cr��n��Wx�ƴf/��%��lK h�c ��R�5�J'�������٣� ���Rȱ���`���\v���/��	=��5DU�L�7��3T*8Œri5.Z� _�
�����aQ�e��b*�
�{��m�ái�W�����ȗ��p�o���Du����a͵��_чt� ߅�>��f�W*�b�epv��.��m�'N�m\*űڭAdjz���]�X��J��(����0�*a�P�s�� "�#yz�V.�"l�Ȱ�˜�)γ
#���:�~�q�'ڸ��k������C���,%�.���绒kn+|NѬ {��DZ��lX���Fy�Jc�[��KG3��]W׼)9ڙĭ8HuO��t�Tb=2�+�JE2�|��a_������+:rN�톁V�&�췯��W�4I�Q,k����4�UM��4���3����g�nS*[���gGk�e��
o0b��Bk�,!yL���)�,�iKr�V\�OPeX���;N��$��%�P����4^3�X׷�k9s
L1�t�u,��G��i�;�9\��Ʋ���G��\� Ǽ˥�t����DI��B�V����]���ᝄ���1�we #cY\[�U
kPWj���ۓ].��]�ް��f��M�a�
{����a���lhh'T;i!\�/Y�p�����;Z��w+>���E�t�'w�yI�]����a��P��v�v60����t�>N�+nt��i�ي�crS��$`a4á+����y�j]^���^��m�[T�_ei��Wn���t�1D7�P3�Kf�y�PZU��x���/s�.[ǽ�y�R�(+�^��W���������|(䰕F@�S][.m�T�O��/���\S���j���k]fV��Y�Lᗕ.�	�ԳNv�St��-,T�O����Q�G�;�t
А��8;�⨧�����ϣ�n�v�5�+!��c��S�q����r��:;GK �n�����^�"p!,w��)^��O����5�	�slsC���{7�b�.��J��msx{"��x;p�wҊ���.j�e�CX|k;N�[̅E�$�Sm�D���Cl>�Ő�6[7���$;|��{�s��ӵ�ˏ��{9��{#b!��Qћ�k\_5�X��V�3w{�ʲ���x��,�w�[����N�t�nK��F��+YyN���#L�6VXk�$)&��Cs*�o$��EM�(ې��}$g����^��b
��FӡV�fKgdƸ�J�j���o8������Q#6W.��.�j�ΰ�JKة�KnD��1Jw-D^����z�ŧ1�f��K��Z���I��Y��=�߷;��[/eߏM�B:�-DN�Ojqu�3l�0�ή%�z�Ve�t����-:��=�s��Xyb��N쳵Y�,��'uvoT�i����7��1R�Y� ���i���f2P$�p�Rt�C�q[��\�x�¢Q`A���2����l]��[4�E�xNkT[|ڼ��_R�K�����F�l�q����U����wU���*�����<��(�ۘ }��b����鶎v�iť	ź�G!���g�śW�'3s�nT	��T���T�����Wˊ
�]Ρ�v��Jx�d�c�s���b�5s����m�ӣ�<�*:���M��_Zf��vs�w�^5��I��+�Np����7��B���ĳ��u<�ZAp�����4@��� �R�>I�p�R��W��mN8{���4 ��!��X��X;�?�`�7P1A�I�P�&��Sy��ݏN�'1u)X�}�}�U����+I����EN�����R�O�K�O��%(�`z���hNL�3e���]�a)�Ώ���-�1������=����.������oNƾ��j���^%zUꭜ社ӟ9�Ԣ�W0��ΝO��W�kn�a$I �$��H/ĐDTE\9�AG.DTAd�#P��2\�"��(�QUs���9VID+B)D"� ��E)�E�L�.���(̊H�\�.E9G9��[#R鰎Q�*�I�"��8U\�R����*�Qh����8Z�)��M�*�DAG4H�I�QR��+���U¨���R��Њ�E�UE�]�
"*+��r��*���")�=XG �8E�8GT �+�vr�	΄DʩD����Ear�+D���\��+�Q"B*�$**�Ur(�U\*�VTQ\��'%��9������h�T�s�D��kB# B�QI
�P^��� �.u��_��z6��ݩP�f��彲TF%�Fs�7��8�g6�\'V�魘7nV)C�\�Nv�I�7����MTʹ}�}_W�fso�w�к�7��e�	ޠhb�L'��VbF`/Lw�`���U�긪M�*O��&rf� �;��0��;�c��J�B�rQ��>���'	�ebF�}Ac��[y*��}a�r��T�8_�r���N%�A���Icш��3�+ڛ�f�����9�[+'��sJ�$Fq��ƾ��$q���|�k�m� ͈(�V�}ڞQG�Ǜ=�x�V�c�]�p�=/���ҙ�����u�7�s!�M�_#Z{�wII�3R��Ol���Gyɀ���fa�Y�kVyŶ�S���Rb�$�Ʌ'd��JV�o7o�#���,P�ϭ4�������+k:m+8�|�T���]	����\�lw�j��vd
���ٗ	� ��s��w2Dl�z�L.��~�s�n+�s�p,�J� �d����J�~��s֜��bt��K���(Tu]H�[V�o+��ϰ��c�6��C0�]N�ʼ+��S#��f�o����U�㪦�yz��.�X8a{��bD_j�=n�{EP˺{`����z���V���Cyu�;9_�4l�����V�۔|%㹫��o�IS(lJm�`��bFM�Q]w�>;�O$��.N	�A�}$>��(�G{rsC��]��;�r᫾�k�����b�OM�:�W��3��}U���n2W{�mf��;�Y�z���������C����xɾY^���� 3.��==���~�}\VV3P{m7>K�	}�乛�cڰ��0�8jS,wM�3;P��cY[
���2��͙���W�n�+�`Δ$�#>�TY�Յ�]|��Jq۷�\+�_&�Q�@���q��Y	�!1�r�P�	aF�+��b���7}Ht{Nnu��U���z^W]�zQ�WuGyS����LZ��N�qu�*4v6���Wv���}n�
7���R��h�c�!�{�#n9����ר�V�q������p����������cx�j��A�{��;N7$GT<w#-�#/f6���k�����Y�r�Ӳ�A��"��W�e2�`C8�з��b�m��6Z8�cYwɺ5�j֓N�"2ȵO���Nd�J��H��O>�\��
Xw�����8V7[>�++��ާ ���[C��{;!����-��/-	�py�ӕ��z���`s����,*e{�:i�G��OՀ/,�&�X���c]��c��[f������v�tX���1�]�4we��*�ʒL�<ֶ�a��潭���i����mc�V�E�(�hf�g*LHWT�+Gk�9;�.S�)0&s�+�9�?���h�!�_~�� _��f��U-�81d��7�y.���9�(�%����R��(vG���K���)��@,��T��s��h��O��P����� 1M�K�v�\��=,��姾�:��hS�W�a�R���;��1 ~G+��ͭ�hV��c�y�����u!,����{^u��g1��# ��8?uD�1��J�������N�z��s�&��ש��,,ˬ���0(�ꆠ0�<L`�Y���(�P'�'.;iW�d0Z�^ma�K[�U�E��]=E������m���wEW������E��}f���C�+���"[A+�C����-�&{>�_n�Ok��mO��](��TN
�|�F�<�X��o%5��U\ѪT@�䊎�䧵�1�h����h\�����;�7ԯ64-�j�8�C�J���\P9��J�Dt��@�,��p�����7:;�ɍ���x�|���5T��A&��1�<��a���`#	��[��,�_-r{R�+�s��[�-E=ʾ�o#i79{���n�϶�X�;�3��PG^�9r#����*H�f��pvTn��NT���ff���&�2�H��{�a-ꏖ*�0�RP ���&؇�u���Xgb�{I��,�Nf��/�V�y.:ggO�������9�8{��z��
���pD�iq,��N��G�UX�|���NX��v���3��K6���"�����!
$�z �d!i"�g���g�V'\8n��g�t�_/!��t7OުaA-����J��A��\jS�Aݒ��Y�%\̩~n�d�����sٜ�p�guV�|��+�V�|��&.>f02i�Z�Q;1����)ua�NMJ��]���.�//:��)��1QѨˎU���p/� �h� �T���S2���B�Un������4�3&�3C��7�+�����MTV�2d��lL�KU0��(֫N��oZ�{t�@�$���i�uF֊t8Aͭ��}��gcU��Ͼ��ь�?2@[�ب�uy���^���ez�r�'j�q��7t�f�Er�&/��A��6�S��8��NKo���N�>�C�-s����p��ڠ<�/z�q�
�CZ��KM�gdi!f�ƱO�rf������39���G���l'�mRӹf'C+�ڣ�:z�MrxS���R���fYS���Q\��4��L'���S��g��o��K�E���l�W^!s��wh��h����s5
�y�/��7/�vu5\~�i�t�������h��fËV>���S�J���I��S�܊������J�1�Ms9�����37k���5�	J|�}�$���D��������ws�S��=�V#M�O;����/9t�Z6�{�2���;�1��p��%"�z�_�+/�n�P����;����iF쓁ڒM�`K�KڪV�a�����~W�VnS*OTh�e�:��>�\�=�
��/�H�h�HOIpW�CZ���m��S�L����U�d���^!���^�t�㩪��q������Y0����H�^c1P�!r{I��<�����z�uOE�!�X�X�E�5ñ�YC�­N���4֡��-��*E`����W����ӑ:s[5���Ĺu�zq��M�ق6��!4�J�� F-e�9��ș��7[2����ޫ�t���<��}I:H�pCeC���m�npA�w*l���K�uv����D�"NqpL���\tn�:S7�����ܛ��8C�d�4��.��E�����:n�w���$W���	��ᵂ�L1"���b�S�DƤ���J����!�4�t�@�`6�q<�V�m:��+]r�fs�ۂ���x��)�R�hIV��l���/C�p�Vtߔ��
�s]�io-�v�}�\y.t�.�3n������$��x��d�󙢊앥�;��'9�
�x>:�&^ٖ^w꯾����v.���Q:�5�����X��֚S�,�m��"�:m+?b��S��|��a��a�*��R�����?�Wr,6C���Ms�Wѯ*A��d�a��'t�Q.s��N���{7RԺe�9eX���C�e\�q	U1��fVK�nb�u]H����S9��v:ݍ�+��C4�T��\��+�f��x�0����;�*�q�S�����3��?�\��M{�5�o'P:a�*�Á��YU��)y�j���c/��-O9r\��9����Mw]U\U5��7[\�n��C��]�ٸ��tO�)/��G���'�զ����2��auy��3+Rn����q��ۆ�Q�Ӏ�GuDB�҅�S,EFҠ��.�&P��чU�S\&��8��A���p��gW��iU�z7.^��#����y:hKy�!ѹ��:��(�7�t,�'r�F?�n�c�0�_�h����	��z��Q�S�����6�c�|��oL�t"5����ʠ�P��Q�_R��k�����3٭���J��2�����}(�z�g�O��{��n�lJv��z�Z�i���S,m70���@�v���x��^ǘF���r�|�"wsg"��q{�cU��a]Ͻr;粭�ˍ+��v��b�)����yt�	�]G�Ňe���퓞��������_U}_Wڑ����� 	�Ԏ�VkEJ��x��pf��m\U�g��a���ܑO��WGF����Sn�E����#.6d�˒.R��|6S(F3�ޞ�B�m���o"�vL�;�̨*0���5:��%�}�/���D/��jb|��xe�Rø/��'���WJ�B�u1Mi0'h��yԹX(�%�9LzìOZ�Hg�B*`w��:
�U�|5�^��O��(���7�k���[=G攲ZfX��"0���ڀd-6^T(�����n��[MNnV%�Q�Y�C��m��ԕX���v�\��=,�13�����ٛ�]<��Ǉa�z�?3+�GyLh�4!l$���F�@97h}�	e؀a����z�qۥ0���pz�!�<;�F�ހ@���S{~��)ά\#��ms��'�/�n |���%J�-H\�xZ��.�D��rWC=H֮7�$�e���jNU��+.:�ՓW���S�p��+q�\*�-���P�i�����/��t6��ܞp��_�2�w��oN�B����t]^�z��x��Dw�,4����͜\nȲ���z:����g�E��F��ugb�(*�\�:&o4őr�[y0�G8)ZS��'�0�T�����]r���G��4�Zs#+��]��9�"Qc=ng� @w�8��x��(}�ר��i���uI��U��Ok��ƴ�|Ot+�Q8+��X}oļē�~�"�W"�J�W�o��n�Q�Df���^��]>^z<2��o���h\�.$�/�[�Q6����t�!�/U���W�&7N�P
;�]�����!���0_J�r�v� ^&3"�l���6�Qt��XR[!�7斡�"z`#_�	�ԭ�Ƥ��ƈC7w�����YϽ���6��<y*��
��NK  *O366R?^*�g!ۯ��8X�n��%��j�J<� �r.9�ү�|��9�#dkT���L�!�HϦy��FxF�L��v6��+TA੾�a�W+��҆t7]���q<lK?J0�"Pt���u�y��r"�9���+e���p�F+�Wh��j�e�&ry)�>&������2J��[��"���=]��4f��[��qJR=y��+�h�g)�OD6�y�3L�
7k������Cۋ|W�8�������'v�U��}Ҹ�Oo���jS&M�n������Ռ�5��U�4[��WѬ�;yW�N��`;�u}�[:;Y10��_��?O`�����^�Uw{֞{��&�ww�wD��� �32c;�zAJGθ���e<��Y�Is���\�������n4�����Q��*��grUR:��k�:{��>���f�z꽷d��-
Ij��oH�<h���P�=���w�k�r��'�w�BN��+�m�B�?"oN@8�e��2���E]�*���^�a��ԫ����E
5(
v�3��vL��������T��\^�{j���f�|��
�a�������6�^�%Ҫ�ē6��z����38�s1|��ϵ�}�S"���faa䪴��r����ܨ˟���0Q�h���Gb�k&Wp���wv˩��)�G��q�!5�fhp�.�87e�ڇtꑿ��!�lˀ�a�IJe����V_ݻ�a���`�}�%�� �U5Z>b$�X9�U�l��|��q]0Y�ʳra'/1r����4G׊�	ݨʄ+�������|�
��-{��#�_*`���w�6�ƥY��3rE+?���3�gjW��HH����,�����H�!��
�*���Z�0���BC�T�P;n{P�J���­L���5�O��UEWP��JF6�%n省�'�4%J��݈�oH�g=��.jR��I�rGs�"
Rt�k�f�Ymn�dZ<{P]/V��g�Q���۝Q��ۨ�t�m��l��֦ͬޢ���C8�|!2�>/�j�Ѷ��͚c3&.�>������U��}��5ű���ە�\^g���1>��t�8\)�|u�ᤧ�mC�BiL�;��͜�.�ٸ�
���|/'��/��_[¾��'INl��`�m�8�r���-�*���9�wNt͚�$�����IF��)��^>�)��<Le5���Cs!�(��ފQ�5���H4�N8ց_C�D�F�R����åʼbq�5>�]�gy���Ir2y�샷:D���W�pW�{�I��`{�j�b|��JF-K&��]��]Q�◆�q�X�iv���e��Fw]������\�s4ܰ	�����cj�x	HWG��c�yW�1��]��8�o)a�(F�mp��U��~>��+�x@p�Ɛ�q�V8����-��]�Եk���=����վ�hnR�Vj<���֬_�����/����/��!1bY豔)U]�������**���R���ڛ���%�������J��Y;�3�)Xܜ=֯{:��[��f���3V.�|���%����]%�l#�{V�X���
?}��{��n��b�����n�o���nLW� �6��[����s�ޥ�q/u�vo�n�W/m��z)�6o�/����h��]_�-�L��wWir�CA'w�K��{�x{�΢Pea�{O��5�(�X+�=A���R19��fh�[ѕ�ƕ���p��,�1N���U����Æ�&�`��v�}I�w1Y�c%3����:�(���*PwXuZ��b���Ҁ�@�Gb��+\%�r�.�E&s{��SV�kA������g�aU/��}�^�˔�$���ǧN������6J[��"p����w6�=�)�_gX��]ujV�;����V�i�� �
9ի�[ns"�@i�V��*ʢ�Ev��հp�ʖ�Rd�\�NH<�'!O_G��Tn��,̩|�3U���R�c]R�`tz�̿Y�.�7t���im�#Q�TT����0��v�QA�h騑�V,���;uo"�M|�`�����ܜ�N,�^�:�V�����ܨ֍�չ����bv*�O4��b�r���OP9����ҙQl�O�dI*Ԭ�-�{��GA��:�]�Ws%�|��kol�f�d�.&�U�� �NA}���{��>T���g8=F�L�J�	΄�y]��j��9��o�d�fuu�o)��0f���a:�#v!���u+zd���>0d�7�(��,��W��oi�;Y������	���n�̡y�k��[��IN6
�k9^����f��r��E{|��<7$����[7'1(]+cx!�ؽ D�pd���{z�-Y�u��Q��0X���+�/��;5��թ����Ѕd8h��Eh^��,��k��@���7�0�c;G!�6�,G)Օ]����V(d8�}&r��r�֓���&}�D7�����*��9�����3�9!da[���4 �cv#�d5z.�^�S�V9*�֞kuCt!
�<����ܽ�I�(�uv�1��XV&���h���B��_%�I�lOf|��ݸ�O����c¸w�J��Ħ֞��Q0P�՛��Р�aj�`�$��,���6��s41Y5��͔����wan�)mj�et2})��yY��9 pol嶓�뢕�?A�Ã���CJ
�wVBN-D�h�����1�$1n��};��;%j��7`��3)�DU��L��\WjWԂZYL��ɡgU�3l"����e�R�@y���d�,T»#3z����b��'���٬�A�&���˕����+�c�q�.ܠ���ʵA׈6�WI@��r���ݾ���C��i;]�ڳ��-����bW��^@Ԡu��=	-(wfT��7en-U��X�+��"���]7j�Ӫ�c���C�D���EEEf�f'�����A5�����s�a�yE�L�F�MĠs.���QT�jG��G8��v._N̊�+77���U׶�.��"T"A� � �`�t�L��.QU�2r*�r�
�TL�$.�G
�e�3��"�.y%T�VTAQE��J�s&z$*:a�U:5֗;�1(��Wt�]Ԍɺ�"NW��h�.U�r�t9�Q�FA]Ԋ+���r�Gt.%r�*+�kJ��H�躙ʹ*�TD��A�0�H,8E�ZĊ*�:K*�EG"�1��R�����%ȹ�QWu.A��*"��G�es�PQ&�u˜���E�8G=]5(�����z��9��dNBr3V�'(���)P�(���@���G;P��ڎ�YTy��(�Q���t*(�̊��%N)M.y!����s�W8w2���<�s����OoI��G�gw0�tG�I�/�c뱴7��18��΋{nCm����U����+�=|n����jy	������>�����N��ۇ��
颲��n��oՆ����n��p���ixS�|�+��O�X�Wrݓ��w.��_K�"�l�}N�5����e�0h�3fz���z��VZ\����Z\
��TN�������a�{D=������8�8 ����Y��I/���Ϸf!p8�.@��NL����^�a�jK1�d���̌Q
��Ąc�I��iƬˮƤ��tM� 騉<�SE	p��oV��\A�{���a�ӐܑNM�x��Qc1�K�p2�]H�<���ke�8�a���\>{�H����9���xS'_~��.~.>� �fV%V)�{ΖO7���<]s�����C>�Ul"��ts�r9�|ѧS4~��|ϡ�VY�F2S�gʕD�*N�1�@��'C����t=99�wN����#�:a�kW!��g��M*d�\�N���(��d-5��U��FkmK�Ѫy"[�ӟV�!�{�B��&���a`,/��P����FӤ�����E�]m���آ�c*��t��%cM�0��U��Cb�)Iة�^�q;y�[��v����\�ָ�n:=R����{�{U�R��j���ܸ���9��z:���5\��f9WĎ;��ܨ�Jy�mK].���3OO�}U_}T���3}N�$��~�mA��<�>x�ţ���6#�uZz5:ɿ���6w�����[2�zwF�����^�Q��Rs��;�F�	�����ey
sn��eZ~>��9�z����^R5
*��-H\�4�6��K�Q ��F�޻�$�y7 /������ܽ��Tp�.q�nhf��W3�B0�*�}�<*8(��UfOu��{�ju��(p��;�ddRN�.�=����k��Yq�@H��>ۆ�}|����:9��"_ŉf�:� �q�E�nH�[)�퇔�+�]pcs蜯��۩\���u���u�6[$�Y^T�|j#L8J�t��@�,{P���1��b#3�	�����[
�b�Iy,&�;�5��q�`ꓺhM}�[�Ԗ_f�k(�f���m<g��(q��j�*��1���J8�3�e#���]9�p��vzw�Smu�+Р��*�+���Ҋ�cH�2֩���L�`��Hϛ��r�W�ؑ��b��KdwAl9�wZ�S k	��avI�U�Ё�v���w�+��ѨXi�fąp��8�w@,Cgu�ş��D�UkS�w۷�D��ň�<@L��gB������W#~��ɗ�ա���w:�r�)�9/�Z��1u����UU��}��t��n�{�]Hp�M_�^�1��%�w�?b0� %�'I�5up��oް�P��Y]E�9�q�W�j�#BMR	ˤL1;����؃���ۦ�@�����̯�T�3�J��t�z���֌�r�d�m��`��Ⱦ�]�ou�,�b+�T��_*>�a����7�+�O+��A��L�=���R;�\�m�Dq@�p�Pۇ1���zj��Ǆmm��+����/��r��D3��x�ק}!@>xk�ܾ�_����w�n8�3���.au����<63������-���积u5	��2�-�pz�����0���mՊ
�N��~}�9�Jy�p9N�K\�VU�./�lp9p����T1aK�fr�����voؾ߭Ƅ�j�s���M�'w���Œ�>=��QU�TR��&�u�<�'!���m�\#�O�ʼ�'r=�=}^�PD�V��i,���[>|�[W�ϱ/P�'>�������Ͼ��1��A��7g����5�V5X�X~����q����y#�YW�\��E9�%e!Y� �iv���L��Q�ڝL��"%v��f�E1�I�i�_R���w�kY&�τ&+a�:jYǗ}P�_(�6��SS. +�_)�g�#��E���{k���g7>" ���}�:�&P���CޫG�I�'G�K"}�����/��5��́N&�c�v� �`� I�\c�Z��=�W���)�h�HOId�WIk�����cۻ땷=�Mʫ��������t�c��6�d'|�L����HOI1"b'����U�-oZ�wX9M�x�vr��pSڻMoj#*�ak�[L�_v��{P��f�5e�I/y��Ze���\Z�F��_b}q7�q���9�C���TF?7�wk�����O(]��a�cV��S��@���h7��\^蟳�'I����9��a��W ��Գyw����/�t���'��>D�f]:i���L@)o��}��v%*�t{7$���x7���F�撲!��q|H���tR����åʼt'��[����z���Nw����iZг�'{z�Uy�E���։�(�����.�T���9ѻEq�T���ѝQ��;�Sm.��N�G@L�3_?/ K�+?���/��B�v��j�j?���^]s�>��U���%`ՙ�;k�*�<y6`9/	#�+Ĉg�%�Z�ڵ���K��ݠ��Bak�7F��:
a��;NN�Tv](�-=�Ml�����oZ)�A�A��vu��wˣ]!�i���LF�kRA�к��=�Z����_}��C����C�S~�ā���^���wK7Ԫ�����3+%�M71B���Fg�g_J�c�};�^�� /X6�-����h�Q����o+i�vK�T�4s���7$ڎ�b��t(�k�~8?\TDu�٠9�T|�tv�Z���1���䩮e�\Q] �ǘ���C<<}Ch\�}��~���p}�)Z�����t�_�y�湏j��.�����4/9B�H�d��������g�@�l������1zp?1�P����1l1���3:e�xry����8�UXY���,P�n[=��Ys�T.ʔn�>L�GӊҾp��4����lU!�RWbn�c�0�[�!��w��q7::(�1�Ok�
��<�n^n��� l}^��]�3�"�0�(�?R�O5%��{D=7z�h��L����gR���M���5�I`O��_	�hgO�)�e��jf�1�.Q���f����:H�"�H�g��l���,�Ҋ�ph=�X:o�ףd�S&�r�V.�}*���߽�01}	��K�
�8�2�A¤��Xݤ��Mk)��(o��Ox�`�Me��l��%V�v���Jo5�n������W/R
�����jn���㫎^�)Ǜ�o�X��;c�K��Sc9�iս32��	��� ���gK]d)��> �ך�!D{�Ζy/2��<_4Eua"#���yμ6��&��cZ�j�(��p�Z?eG>��-Yg�LOъ�D�Rv��s���RŜX8�2}����P��I+�3��{ԃ����ų�~��2^3,yDF1	�:�c���na�ݵ	_,-f�C�-��5��^W��l�]o��m��5W&���Sr���ɡ]K$�%���"���F�G��t�@��F��t�ի��Kkr���u�'љB�'[}�� �o��گ��u�Lr���g;N�>��^�wKj��Y�-�^:/r'Ԥ]����f�}d��z��	�+�����/$<;�a��G9_�\�c"^>�n�o�{�4s���*��\�K.�s}�����ʾ�z1\aq|������+�nެ�;T�r�o��V�j�e�j;\@/�''�6�5q�Z�إ���i����[����֢q��LZ�1V��^�߬����=z�����	�Y'�l����^�-hyz'��koGc���r�E��B���\��(��2��Ǻdή!���ʳ*�TV�;������.� �Gu������S۠�=���J�\��bxq�|DDd�g�4�_7J~�녘�Ω/��bR�kyoCX�=��Q�X���{]\��#���B��`hQQ�)9�bR��<�rT21om6��X0��F�y�l�U�O��邠��f�jJ�V8��\�0�:����vE�K��Yi�]�>���q��1�wI�BZ+�����[M8j��nk��Ub}�ZW���E<gYe ���+��R����S�~O)�v��ji_̾��+��æuLmYV&��A����!zÛUn���'E��N������6�6c�)�3�2l븩����;�^;�:[Ubv�89��;<���{�;����F�E}Y;I����l ��w�V�"b9���;u��eb��)���0O�����T��6pd�|�����nkyU�ֱ���3}.�K������Cv��`9��մ��Y}��6Z��ӼC��=�3%;���&Qmj�����Vc���#��$R�1%�­��ړ	W]�Sޡo�p�ls����Jo0�x�)�ἧ&�;�s�����:��gt	�Qk�_+�E3������G�}��K;u)�!a�B��{�ڷmKیN5��t:�Ǖ\��]��`������i�(��uܸ��+6�K��ڢk;�*^2�>\����������x�[����3�q����끊&;
�ϛ�[k�L! �gm7������.���]��Q.z�iCW��
�cb�$��Ug��8C�j��K����ۺ�.�õ�h9�:��/�iAX�����qH���M�E����;m�&�\���ʌ���v�u���'��y�Zצ��5]��~ʋ�>��P��m��5��=���6�
<��x����f,���APB�BY��Puޚ���k���Ψy�)JT(&*l:���LR��}U�־��*�wN{�ম��W��7�*!�;�̉)�->��e�zm�t�?�����������9oԚW�o�o���4zs�[�bsl1����������l���Y#�^{�30l�$ҷ2�Wx��g�^�r���Ջi�[�ͥ�z�
�e.�ﳲq�l�,[(4���0�_xJ�J�����	k�睉�ͳ_��6�~���+F�-Q<r��G���Y���Hg,�;e �
]@O�����F>9�:���5.�
��0&�����;G"~T��㎁�:Q��j{q�QC�y�/%e],z����$�5��w�#�:쉎Cb��wo�<:L�����SG7+:�J}����uZ����֜3Pہ��<�ׄLk
��x���/r3��k�3�y����ŹV�!)}bpʿ���o)k�6뵿	ٙ��\��8��Wp���1}��ev�_E�s���OZ���Z�*��6��()���Tz���������U79P'�:�b��|�td�/b����֟{H�^���5Hk���KH[=ih�V��+�ίB�*�Vv�VZ�������F����sM�-�}+����Q���4qʰ�+�ZZ_��^JWff,������lT,e���t�_V�:��^kV�^|^��>�F	����)i�oo��+n*�Y���[�i�җf$���L.
�l��)C�bl0�H�2-ޭs�0���b�!�^r[:4�[�]�s{�aMu��,uo[�ѷ�����v�̈F�)���QX�t�������ewg2��aeI�ٕ*R�Q[���k/=m<�7��<���Hl���n%� ���@����K�+�:�RҊw�4��uCeS��{�u(2��t�A����*���%�|��r��zP	u,ޜ�o+U6N����O�Qϑ����KE�SY�t��M�]K���A]��{;���k>gpT6β�"���>��i�#Y�[�{�X�oBJ֛p�4��ش9��*������<�(%�ta��+;4b�F��ˉ�����M>��a�\k��ȘNȼ���86gvU�=Si
�c)���y��[W���=i�=�2یc��.^dޜ*�g��>��� =Yd4�O������^e}8��}����0�{eD���9���6���>˰"�έ;p��;5�F��-�f-�yQԴm榾���hM`0����a�H�Vy�xC�>d��m�3���#���p��*ak0�K� �����/1}oU�wRyZZVv���Z��&@@�N���jV�[t�Jmș���N�y�:���)[C���	1M?�B2�Z��}�8k�M3Ě�w�Pt�a�-c@����<��ԙHv�Cz�e�����u/z��lB��D�a0@�s�����櫇y��C�W.�$�*���o �c�Kr���ѾO���kv �]{9�9F�����+T30LJe��k[Mm�w�>���:�{���&rVY�-���ڈ7&���Y�];־t����W'���&�j�0[�x�\v�e��4��R7�Ebw9������ȷl��`���vf�����q��qp&g��b���E�'��B��ȣ�Uy�٘�>\�^,l���@��9�5R�������tJ:�}��=��f�^WV\G2�9���c��k(����
9�nVҺ&j3y�%�*J�'dp���Д����L�sc�U��a�q�iB���wM�6S��w�<e,�;�I��(̲�m��}�Ь��]i�{ͅ�ed3C`Z@��͚���"d;0�\Q�G:'��Vob��p�k 2}���һ�XU������?m�"5Z��q�u{��u�K�R�v�֕3�E��)Ƭ�R?
�g>'�u����ZY�WB�S�E!���Sy!��m��g����,kY١�ak�a]�7�{�X���x76��u��SmR|�є�nRԑ¦\��C������} �z�vn�i�<ǆ�S�.Z�[c�0�ޮ�8�E�­�n[���nnV��{Ô{�v�b�F�����t��G�Ƕ���'yjB�{H��;w�G!Ӗ=�i��Ԩ��ޖޛ�+�'�1V���;.��!�\µ�e@k�r�5+[7�2g��v�X10�>�V���4�����?b�B���85Q��:��`���h���rP�U��YE7iR�8l�Җ!�J�����F�L�����>��N/��mdvd&Ծ��J��aW���]�>�fBl`iZ�����˕6�J*9]��1�e3�]�d�yYA�w}-A�v�N�m��p��_��bZl⠋ע��gV*������Q�ċ����}O^/��c��d�7].�#����U�,�JWC�kW4��n���U,��ڷ�t�ĕ>Ӽ��{��T�9���ܩ�(M���fB�{ZƵ�E�������*�-�wƤ��ͭ�bjP��9��Vq�_M�c��@�Օ!��&B�p)U��vα�%&j�r�eJ5���蹑pӔf�΅֛�81-fm�9Z�uc9��j���Kj�f�,V��Vy�d��͹�c�����N��j�s㯞t���_
&�tk5�:MS�*×J�]����q�5Y��AҞV\�ε�А�{!�A�W��WI�,.�ιj�������������^=yǖr%K�"9��"��<���.^�qj�J�E\�����+<�AB���#�3�\��.Q9��4C�msD��PDPI��"�"T($��QD\����H�EEzЂ��RK��r̓$§\�(��I,�%4Kj�Ý*G2�bT%(���Qr��s!����wt�L�QԈ��4$�9:���Zy᠊̝ݻ��NEr�US����
��+e����t�76���B�40��٥E�r�ChhD��� U�QP�TT3#7\pBTUi������'t�C�/V:���%wn��S�g.$�j�pԴ�$3KJ�$$��ܜ�eW�V���\=�R��gP�3(�dPs�8W("��q��g�Kb�)#��/�r�WJ���T��nӉfr�x�|���Zx4v_Wsz�K�*YWi=�R\����������#[��K�vL��;/.>MƵu�c_�s�<�v������|$^p�*���y��UG��P��]��ASͅ�yz{S~P�*u��8�-��ˋa�N��ܜ#;82�n�>��������JM��ޕ٩�tFv���/Z�U�g,^��j;��ԏZ>�NX\8G�K��e���B�����簦��9���uuV�-��j��V����yTI}[J
�J��o/硬�q����fVj�
p,��Or�{�(t�06J��);��
������m�9�շ�'ff��O�5��=jr�6�|(t�|�J�;���jI�4����K��.`rʣ���4��_�k]��u<g)�T()ﻧ�6�����jGO�u6s���8��+�O�ܴ��[����x���Y�B���^>�]�.ԝ�)��W�j_�3q�-�qb�>���ضyl��ʻ�Vٝb��9�f"r��8��Ө�q��.�YojX��S*�1�N���I�>3^��cM�_Z�0q5���:V��-���8>P��ۓ���s��[�����)M�����4��$x�����Vf��'��|n院��kz>}-���ꪯ�b1;��۪�ϣ.�ꁠ=ryvWGru�����6�1�9q����n������Qi��"]"f9�8꿊ܚ��qܶ�<j����ڪ;��5VfQq۬mƻ�g5������8��Od�t��]�>O&��N���,��l+�^[���V�5��tZ�Uf)��"��W"�ԻǞ�Vp���ڶ�y؜kZ�m���7�]���� �;s��̺�1���mm@��.;TV>|T�g!=j������~�۠9.��gJ��ޙ0w�+YP]�r4o Jc�ob�_|��u���@��z��;�ϫ4^����n�|;*
�z��=S����U1���Òg5.�����!h����g�f�ϵK8����9Α��}G�����7W��kMq}%�n].c��5��i��O���ݶz��T��<�mK
�)�,���_pԮ?m����_cl)l+F웢�.�N����)�%|	��4��z�h:]�e'�8hV�;�~v�u�i�C��d�hn�j�-%�6��o6G�3O'`.��CT��tÊuhp���O���<�_}�}9�ܒ/��o�)�U��P��������|�{fگ������$�V}XmU�U%f���#1�ȥAԷ��^F���=,�^P.��#�P�V·;��%�2���`�ފ�o5��v'Ǿ�/��GnD7�8퍞S��إ+Def^ΙDw|�1�-5s�W�xe$��8<�S��6������u����t�B!t�F��j'�n���ʪ��8rW�ҳ_:T.�hˈ��5�o�b�}#�*������@뒵��\��`�����vt]vS�%��}	��5�B9�ȞCb��)��k].�;Kk�B�[��e��[Y�9uZ���է�Cn�<��xFE�sՇ���6w[�K�P�^�]��қY�l�?E_9��۴���'�t1jVg*6�����cU@����&2`ZU1T��+�v����}/X��R���||�AI�����+]�:(�y�u{@���0x�҂){ju���I��"������n&���2JF�p}�����6iV�K��T�!;�7+2r�pv.w���D�F�c�:�H��4v�jg�;a`��p�N�0x8��ͧ,-g�}��}%\�>�0O+��_��Q����.�{M�T���uv�zab�e��S���ܽG�g��������FU���3* ���\��/1�U�ʹ�CkГ2':�4��<�����I6��%v�:������\�\y�W<MuJ��-���.��1��5|�}q/�Y���3<���460wn�r&iu�)����ė��NT�*1�qCY�t6��N�nMA:��^�ѽ�i�
?v��
��!.خ��ZBN��<�
�7[��܂���6�t�=�P���}0T	1_IZ�θT�u��t�k�BU��Ĩ�5V�N.����r��!LG}�0X%-55���	�M��ʞ�w��Z�����+����3�)�v��0�\B�V��X_�8�䞭+��xC3��g�=�ڈ���/��gV�D�*Fc����X�~Sao.�o+��'LM�3��mLK�3��.�#�C��4��s��S��ӕ�f���m�
f{rir� f8F�y˺VV@�R�x;K��U3Y�q�X��ZC�V�<���Z�o9f�NP@s�)T4���Vǝ������a9k��U_Q(��|<]fR����SQ6�j����Z.��4�a���.R�TFf%Y�뱠I����
��˜�q��S�К�i�<��
�[��!e��p�B��)Y�W�e�{h��%���9�ק�T%��V��́S���5��gn!����g��=��wΔ��}�UMb���������Ӽ޾?��Q�>}���'٣K�K~���& s{��M�s���8|1k��\�<�R���Y��z���r��E����4�����ꛜ�����D���o�I�r���Wf�'��v��<���խզ綨C �sմ�-����Z��v�� e�y��,��Gy��rx�U����h�@<�$���PU%*��A0�����V�bכ�; ���눖�
�߅���_>WRw�u��L
��91yV��D�ni���a�n�XI�Z��7S旜�w�s�쭃F)��r��pt��U�J��OAL�ׅNº���,G=QN��Isgw)X�i��s�϶�ehr�l-�:����b���`��J깂fI<�F9V�5�����tOr�}}빠�ܺ��}���|�z��[fҨ�C��z�Q����DOȏ�9�;��͙��S}Ҷ[��pֵ��uD<g+�)T
��e�$��֨m(��oX���B9؟oD9i1z����O�Y���yy=M�0���	�ڣE�N�x�����L>C8���\#��^�_+��FLz6єQ��4YZ槗m_ru���s!�6�vfVkg�&�R5���p�B�9��e(+rny��r�t��yQS��[k�8�5:�J�[Lmƻ��ׄr�-m@v���� '��{���U[Zө��E�]8I�Dj�\��F'շjʯ���X��Z�
DgI��3�A����2-�߳����m?yE�[����q�k����Uf�v�'7{!�@��B�;}D�V:�����O��/+[ګt�M��*6,ȹ��*��m�Y�uԔ�cK�+4͸lԺ!�.�Ma���b��h�i_^�V�3�6��Mz��lsd���iSź��_Y+]]��>�[��6�e�Mvg;�]�-$e�KJO!�c��?n���G7�����������)S��{v�:M�xU��s�%1�Ob�Py�a��T���)޾]&oV�I����ڷ��X��Ʃ�WM��\ՙ��i�/C3{���W/�o�kU}�v���<�D>���A5�:�ݪ
�l��kb������o{h�Rf
��Lf���m��p��)�m���{��6����yͧ��Gt��ym7�j?15�o�ٻ�.��	B�k�Pu-颓�k�|3�q���f�Ob�����
W3���!-7��/�1>4��!o�޵��cWy�(q�V���u�P�����j�:��h�r�@�����=~�kG�(�i�����v��!OJT4)����.��Gք=�`�x,1{��g���o��gh\d*C��χX��[ C{}W�+��=
��昄�ь}�ˤ���m������`.���T��J��f��9��Y�}�tPC0V�zh�b@w�^ޫ���.� �����Y,;ͧu�Z�^�:�Q��h��N�Q���I/�"d��Yk.��u*B;Vm4�r?�U}���{wLZ�~�ݮ��t�Q���q����vG!���<q\�|�j�a����a\��˜�f���j�:5�3M�\���9�T���^�.�hC�/�>����:V���nU���N鱐)������m�p�-����z.������߄�}���s�	ݹƹ���.n�.5�(
���R��Ck��j#u��]�b����=�Ӥ���|U�u��'�,õ�$���Oz�{WO{���j������7�����V��?N=L���b��q�S	&���|Wfl'�:��Sє蘜/�$���c�Tn�v������=_HW`]��}r���o_T�����ٍFԨ��rtet�:�=�2�oԕ(���k/=����4��j[@d��O�7��Ps�s��!򯤥���)i���ٚA]I	�{�������79�}�
��'f�� ���珸;��w�M#94q9�3�0{�/�P})����e{��$_��^N�2��ۑ��ku;D|�'��B���U�V�<�ʝ5=v�{�;ȶU�nΜLu˔��F&]��F��D�����D}v�j� V�B��q��:c�|W�&* jJ��t�cG,�U��T�]Խ��p�>�lgS�q�P���Z	t�'��g�S�WY�����N.�p%��Х�q�9�g��
m��,�"�HJ+8ʼ$^�����b�G��Ow=ςn�����������{��K��=-f��Vq��P6�k����W��}�P�Q�i0�̝J]N9����N�#��u�;�^�ȼ���\f�psH�z�(�����c�D�u��k��#�����?yO��Ƕ���[�.~��}xZ�ʗ	�uj�V�ɞM%]��*-�;u�=����UgҒ�˲�*����5.B˙B��5{<�.��8ֳ]�{�B�7Z�eָI�]��msIA�ˌ�q*r��2�TLV>wO62^>>����ZB��O'<�noU�K{����+)˔������>w��.Q����$�(��n��F2�au����L8��@d3���)P�s�r{y��Mc��B\wA�w|�A؂ۻpf:ަ�K,���"��fa�5{u��Z�k\����`�/�	����W�f��_�ַ�O�8�~Xqm�С�gKbN�9��t)9��[�w��s0��4X�}��Ep����d�\�L�cS{��=*�9\̕8:��3����2>d�=v�zX��=6��ߗv��VK��3�E�����YqS�i��ޡC��W��!'�������FV�|�T�2��+R��5�B���-�iT
=��*(.A�8��Ә�QT����X�[�N_cX֧�9�7��s��&���b��=�i�����5����f#�Q��2�L���EC�v)s�S�xN�;��9ﰰH�!o�����=��\��X��$Ҷ_�zvֈ*��ⵍ�*4�A�{٘E���k�˲�Sz���=��݅Dbά�������.;upˍv�D�Bb9�{�d_�Qo�z�u0U����5����i�2�.�&��)����+e*5x�A����G�Zu�h�n��e�q�����2W�zS���^Kx�6�
�艙��K�vV�塊d!�>�yu����� H�7jɚ��l����-p�����}Ɍ��cxv�Y����
i�0u�otu���Y�g��T��((mC����`�;�ױ}~���^ 
x]"F�,^��[���;�����6��������;��:C��h]�n:)Z�n�;��@kGy�=Bu�;v����*�s����|�u����F-}k)�L�X9�n��rFX]����{�k��V��k�H⺯�[��N/z{B�����\R=3\W��,��دqTw�ˬ$�O�,ӲI���R���J�7iefZ<�Aa�;�x n�=�E�o�1ݡm2J�%�FF;5�B����i:V�v:�:�fY�y��E��ή�U㊲�\�5aX ��v��e���߻{F1NX�-z�}�X���l*���h��c�6��2��i�_r.��KN���4��N��`J̈G��=�g&y$�����l�{;a�-�*�-�{���C	�w�v�1��\M%��U����i����"��p��q݅/��m.�e��������*| ǋ)��e�������e"��Ʈ��,�)HEb��M�(JԔ�e���bX���k.�=�eɝ�n���8�3���|��e巉c<��[!G8���[6�+ Y��+���I���$�3�M�*���z��Y��5P����c��k<[M�ޱ�T���Rw�W�LyY���'�|+a���������۰�To��<��-���ٵ>��L��/���)�K(��J���r��&���;�Y˩������������E���y��ft\�8˱�ֵ�щ�	��B�&vU������s~5���-��W�uF%�4!\Eq�sݤ̯�-D���l�˽+Uӭ�iN���!����w])��eAQ��*D�1GY�j��#֨�Y�o�s�F)L:���4%�72�f]�����4%J�`^�B�I>�:��m��ւZ�p� Y�ikH��M��/jm�ئ"�E�.��b�j��`
�4@�kV�����{��DOm�=�1.M'Mc�p��W4`�,���X�勴�ޞ4v3�F����T�ѓm�j�
��ALo���-qX̏�� �]y"��
~ �;]v�p��/T�(�"��G��U�	F���z�׿:�\�)\�f���l���*�'1i����ca6pQ@%�C7�Y=�寋��nE�Yg�"e;˛���.�)4F6�6�{.B�aV��bׇ�l䛘�&���tF����]�	A1Y�z�0%�ݜ��`Ĥ��6�ۃ�ޝ�X-��º�ƴ��^xUi�䮜�B=仺X$p|����bK_#�U���*�5�36�Y�f�IUR�9��C���
F�9�=��QsYI�W,P�"�GL�H�j�w9�R�H�\���2)$����2w
��!RDV"�㫸�9�y����UG")S�UQ{���rJ�;���Ow;��Dj9]��*!�;��,��Iw�8AK�p�⒡+D���9�e�4D)��{����]�ݎy')V�/'s';���*��$2�i{����,���W�,�ЂN��9���J-�ZG"�����,�`�sf��IQ$���է$5K�])�/J"�IM����,Ԭ5KBAs6��#�y	%��%ez,�]]�2ʋ�Hʭ9�'qR�����Q1i�/q�S�R&h�a��#�I���Bg�����9�B3U
���&��t�j$�pL��3K��BE)5��`��� ���ݪ�E��TF��7VU&���DVY�^\hp�Q�g�VN��1;}.�j��K����u&n[_)����s�=����b��&��Z�|ۍv��k�&#���9+6� j�m�[�m%�fga�O�յ���u׉�5��o*�Ẉ�9���vͭJ�/��z�P�~���߲%�7���;٦�x��N5��]���v�uEɊ:C���z����C2����m�	X2�TLV>wK��ֽnr�1�zi�e9e{�Y��>��iz�T8��~��s(Jc�(�\P\�k�ŷ9w�)"!z��MR{�3�(C�[7��U�7�s�:��0&.���׊6S�����7���܈v��}�mjγ��h�p�h�O�ws-�J��f-j��N�kc��k/��������������*Ş��&o.�v9����m`oj����4W&���އ���ڌ��7DuV��BP3�%�.��;�4�~���-5�I嵍v>�1��n�fon�ER'�Kj{���*����W1��Gv�Qe���@������({�
���ԟf�n���x��͓)������(���<�aA��W�[W2Sw!]�p+��fN�s]4�d�����Ж�b͢�(��.�Z;�n��QT��P.d#/��
�.
4%�~�=�UpSWz��� קk����l
�O�]��xβ�"�|��Z.-��U|���4�[��ݼIu3�H7�3y�9��3�+���;fQ
~�J��S�ͺ����gV4{�X�o0�����j|�B�B�&:���Ȱ8^�n]oy:q+�L�h�q�a����2��)&}	�օ�F�#v�"�[���b��@��[�m��D�/y�O�����tjӆk������bѲ'g;4����<���&?{C3�"^eGR�S�{Mi�p󢂖�޺�b���Jt�\}zź���p��.��:|�Ou	X2�9ox]�n��o9�mD�3����p�ֲ9����i�7]�E�{D���ȭ���bT������\�	�]|��y��b���G=�ʳ���AW�*�dQ6��Z�p^c��-��vnv�V�O	������:�p.�:��"Re�֫b�4+��O�\�Gu��f���K�w�ok�[}Y���(�#eM6UlAf�|���W���c6:�Rq��v���ۏ�vc�ZX	ig���ڕ�Tfo;ת)+�L��.\�	�}�GtaLRI�n��]�}��J ��ݣ���p��H�G�r�uD��*��=P-!_v�i��/�A�a��2߲����{��x*=��yTIr���c[ǡ���N��XXy���� ��n�3{�(t���v��f߷;��-L�On$�����R���v+�|{�F��L$�Ir���g6,�-Z*/	�q��Q}܎>����_<g)�3�!O}�& wJ� E4���[+80��d�K{��KJ�֘�����N�����0����ɵ{�ac��7:���}��S\ղ�;gL\�ی�\�7oS%Z��V\ae���F��z��mo&����4�a�M�Z��ھm�
G�ӎ9ݑ?r0
��ܼ��{Y�:5<��@����_R�.�ˢ+]̴���<5��`��T� ��7f�]S���x�]J��d��6�^�}ξI6�}�Ɋ�s�C������qc�kυr%��YZ���,�(�g���Mk���,����{6��� n��t�
λX�r��n9�}�gۮ8��D#3�cp_m����T����]y1m�Og�ΔS�^��ػ��NQĲuY��L}P3��ٚ�4�YwJz�kU�6�y�׵��x����'��}iX���\�Rc�z�;u�c��jnr�O!�ڢk;���/\7Y��{,HﶵEMg�w���qy4/TV��9rv�[y��PQ?_.{�����<ۊɻ^lR���{����wo�\W���	tF�j�62��*f����kW'0����ҹ|��7��s)�y�<�"K��PT+��8�y195�h�%en].c��ZǩꖟY��:~��*�S��ٺ���w}�+]:
��Ԟ�����B�y�n�_
�>�9��0�u��Q{�6ðL@���*�q-�e���k]��uC�m�w�[S}wWV�U*~t�VWl9�&˾ﺓ�ѨLr79��TS�+�q�mp|�cV�s�n�p������̧��`����sC��@���s���a��r��j��5ǯO2QU�Ɋ7c:�:"�ї�x��x���!��I�ɚs�����C/�}�s�1��衼�d#�Q��[������
L�:��qSKruR#(�2�Y@u��H�O=����qU�.:�J�
Y��K1�*���Ü*{�A��*��(s�	�k��p;B��fR��I���2���5�o��eƻ�r%R�l�=�2*=���NH����޽�!�^��Kj5<v��V��M�ց��xD�r���ɞ�\�-4�q�P�f2_�]�M�:��[Z��'4�qI@��yU������D��a�]Z�����ե"��槗4�R����ʍ�u�s�$&�ͭ�����}1�xZ�$�J{k�=�.;\�>abVu(r�s����0��QTw�����^je��g��Z�y��в�L���-���S�9DV?��43�X����sި�<�es�;Η����EV��I^�~+��V������xJ;����v���D��t�J�|a��)��ת���0KwM� VΝA�!)w�f�'-�CӹKb�G���S�dze:�74՚��o�F�,��n���Z\fu�2,�=����O
Q<����i6�t��}�ڢv���O!��87��k)�s���xe�)>����偬�������F�!�;�8�~ei���zi��-�D��dvOuW6���k.������Qq��I�w ��.��g�A��-.����KM�[MigoaV������ ef�{�F|���O^�n{�55w�8z����9�pz����0�}��ෲ
����f�>�|á���*����<pwa���G&��9�d3�*{P홈D)���h��Ev����O��z�k��Y�r'X��\����8¶r��Go32b��DXv>�<q���U|p'ٵ��nt}��}'RLT&�Z����tjf��\���n��K�\y�_n4�)�5����gz�Q���(�k��Ʈ���ܥ�cZ�b��;]�w^v�:���}i��LΡ1���*�sr�[���甄6�SG�6<Wm�r�{�z)�]p4j���L����-ucH��H���;���
S������%������SD��o�s�znf�\�{����ӳ�6]N��(�.ʦ�������gu{K_do'�֞�{W��:�bK��De���T���K��o w�)�m�)����u��d;�ja������O2�}&�_����ֳ]���k�H�}�w%z`{{h�2��M,������17¡c��ϊ�l*�����ߋ9��֗gEjX�g���R�;q��\D��	p��
���LRI��+s��<��"T�������cQ�V9���t7�J���P��}ػ-4���R;1���}�r�'h
�f�^ٟ���<� ����ebR����p��&x�Wd�@�x0{����On�P���x��]A��\��������L;�8o��������^Ql+J�P��c�;v���FB�\�\������}Ҷ_�_W�c�l^��r�ʕAO}�A��
0܇Q�'z(}q�,g����s�9�[�v�J�V��DFƯ'=���$�E�;׵���Z�t���w�1ծK����s��%�Synh֚Ӹ��=��թ+U}j���K���$1T8;#]����4��qv��]p�|JO+��D�	�يG���%!������:�c�vږ����������w�fƮ�%�yq�9R��Th���N�{	wִ�.m\2�;�s֘�t��q����^[���q�b�A/N@I������m^�u�嬉UT� �+�9�m`)��kb�>T��9ì�+p_;��[A�9��Ξ�n������IQ���mƻ��Dl^|+rvK̺&����w�;���͎���~��W�	z��8f���V�7Z�E���b���Ţ%�j|��ˌ�=v����n�[����N5�r6ݯ�Ѧ���a�ܦ�T~��˴�B{>����P����������*[�>��7<2�'.��U%��}Z�1�}�$�ó](��^�ʳԪohgw�WQǷ�UL����o�B1���y�Q��W�V���={+��ݩ��W'�9o��V�f��N�nQ]�ˑ��V�r6�&s��R K��;w�P҇k�h{`m�6S���Z&�M�w��/3:���vX2F����v�Z��
��U��Z(k�ڶ�v�*ڗ��q�9��7j>�qa��������E`"h?�y-�v��}��1V�6��7��yU쨱3G�	a57o�9�ʠ�ˍ]]n��j�OT����􎸎@l�fC�|�n��c�J±��Z�*��[��T<)��wR-U�]�Pk+Zٞ�&���~=[3�\5L7�\��ֵ��gS�bک�} ���Q���C������P�k1����}��[������=����"�=L�9��߻���<�j�|�ub㱌9S�ւ��E8z �[ҹ\C8�o#b�0����y����DK��Z��g��YWK�v�O���|
!R�lC+��ܓm���wx�sU}��/�Ovn;�֦��5	s����D\r��O'��2�uo��s��'﯎N��ҟ=��m��N�ӄk���o)�	�&`���B�կdկ��O�SK��%D0���JeoB7�|yw��a�C!k�2V�b�;���
p�JT�x��p]
��,�o7&WG�of�b�9��vΛBS��f���S���0��	O�]fq�N��tѮ���}�Y�:^b֝�;���z�;�}{|3:���{nju�V�}x�4���:|Q�>��^c�?}ym�8c��q��]��{P'�gk���ƌ���d�n����н޿8�/�m.Ojiu��E��"ԣ�Q��kھ���Fn{&n�����7͌u����|��챓�vTs�;�ʊ�Y5QsuI�y[y�̭�W��P��4���I�[����Q���H|����\|�E�Я{<:���@/�϶�:��_����[i��K{F����z� �ȮK�3.0f�����OuN���9�6�ކ��yuqip��_JZi4I�͹�g��~����+�:�����'�S�su��\'��=C���E-7���b�w5!/��ћȯv��8HA>l�����;_C�e�;�!�{�/��@���^8L]Bf	BP��*];J����\�6L���ә�iht�>����T]�Dt��p9�Eu훾��T���#A%�d�{�W�i�=�N��mv� Y���w#�vX�8켺�g�u���M���FVʅ1=�bF�����㮮�j뷦�*��D��R�f�F���������ψ��1 ���:�qj\6�X$J�Z��$ڏp�b���l7yg3X��٭d��#�(����	���t���
�+��GE.��t$�WG	�.�u������u�$���N�9���hWwEI����:�O#����׶������*^� &����g�b�
���j�to8!a�<�m]�ڪ�ݜ9ƍ�1[��CWdR���R�����,�����C�&��@k��Q�������;��aN��qx�h���܇8���A<ɎB�B/
��5�5ΰ
Uv4�8�A;Xv�K:'��"n[O�o�.m���*�4��u�O�SA�p�в]71M��M	!�'j虧q�����ASw��,�{�ok�w\�Ǻ����g��ה��T�U9:��U���xs5�iqugCJ���3�6��:�[�Ct�����]�֙i�[]����^:S<�.�E��Z�e �F;M��Wp����Sz��~�4a,�Gp�ک�;B#��k��%!Ft��YB���J V��b��io�y��A�ا�>K3s�*޻=,E]^95r�k�3E9�Nv\C�4"���tos��M��ю:�r��XM*V���hB���NZ����C�@v���)�Iڝh�������f� ��|�^#�o:{6��6�-�L�v+%n��H�s����Λe�P��6FV���!KJ�r5�-!�aw��,'Q��#V�=�oM����df⵹������}I�M٠lt��%��<��z6;�ܴ������q%�	b�}��	��_Wsn�J�S[ص��&�#�>��.u7���S1�)Vm9t5�ޡ2"&���%��k������-����%�7��nV:6�щ칸�YNn�zO&ì�s6eZaK�jL�w\U�*� NN��z���ř\��{�֕'P��V��o��E����b5��cv(�B�ŗ�P<;�A�t�}�>[x6��1+sNh�B��kH⋋�s�e	�	��mbU_SX/9S%�
�6�1�4+�&E֞Y�Ԇ�H�?�>7.�D�����ޫ��>�=޵�(��Q�B�D8:�F�E��	Ԉ��}uc���u#�b���\5+�2��Zj�Ug&�kqt����t��M��h8k�����.����c4Asƀ�bg5�/���n�-���f�޼��Ħ^��xؗ�5��{�'&֝s.��Y�ܽ��eH�K���Ofs�(�YUR�4"U�*a�xE�Zs��e���TJ�w]�(��QI!*I�����YS�U�L4AUZ�!ڴ��g*-
ʌ���T�dh\�
%pQeȢ$�a�I�B��Er*�p"4�5�\��K&�g<�!�*��J� �"�ցDR�AYi�ʂ(�E��t,T�
2�Q��*UT**���P���͑,�I�SL��D�4+�=2�P���mB�<�RL4��m�E�0�KK<�*"��#0�
Rl�(�-+��t")V��Q�QT�Yò�9U$�&�E�(+���&UvW3H�&��Q.U^Bz�9�7<�UW�e��-�)[��w�W��E]�=r/")Me��UI��:�C�p�Nk�^Iy�R�:�Q�t���U�f�����Sk�G<�gC-1.V)N���M330�KV����d����"��EL��]�,nwO��S�:��;B^̮�#�� �7<��I��uZ�P��sƽ8q��!�Y�'9��md/�.���ܮ����+�Ӌ����[ؓI��͝�M�t�B!OJR�qT�ᇙ��۷�c�F��3��psu�>9P�:��l�	��T��9X���k�2�i�4��m[9���8�����ޚ7�1P��t��M1��P8���ƮiWa�^�d^Io.<��ni�<��j?o8���By��������a����V�#�إ�z���Z�5c�CX)W,�*ہ��iˬ7&{wV�P��C),��7�b�E�ٷ��H�t�ҷ��Uq�2�4����eKˎOZ�#;�ͯ��7Q�w%{�^TQݡ9+ϓ�;��xہ-��zx���Z�����ߋkHY�߃[#���>,�nR�b�8�9B\>�*&�1I&źo���Wj���"p�D�Vf8��㨂�˪Ѻ@܂�V҄�L�ZCc�v%�0L�����P�g�P]|u���ݹ�u8��Տx"*�*��L�ڹ��ʳ9���L̫Տ�Z���O4uOJ>�Y������z�q]+���r��3��W�a��y�7z�K��Ar�����D�_N��I�|nn]ǂ@��<�:d:��<��G��/*23=v�xՇ6����eTbT�5=���W�=Vۊs�����Y��6�ٽ��P�@B��dI�מ�)�y�e�}ZZ�z����Y{�p�|�\4��jvR��P����P��7���kA`�7��8[X�S�r��,}��Χ��9JB��aM�[��%NV�ؾݺ�J^�oЛ��~��g��C9���M���D��tv���"����U!o+�L�v>�7O5��a�F�e�gfc�x>�Z�H.4�AƼ�T������ak��]�q��F�p����,P0uz��0*��F�����~?#�?* ����@w%nT�J�s�Z Z�l�Wd
��J��t�ƥ�i�5���6�]���k�62�nT};�3�pSkZ�w��#J/Vw�O����wz��8f��7�_k�u�T��� e�0U{G���o����c%�OmL�ժ�I[�箋֩Y1���sqZ �l�s�G=��:yi�����4R�LY���$� �3��CV��w��й���)�xt�w>�4Uwb�6����@����w��nW��k�ZgL9�{�V%�y�>����M5��:����N5��t;�G3g`�Zj$KO�!S�8t��h̯�遘)f	�3�GV>wKb�}��<���
��r���&A��s��p�𑞈{5��}��E��a��.�I�G�K����t��}��z����w�2��r�vzb(*�jv��2���<bzWN�ֿ�o!�7���_eD;����3���� �e=4���b��|!1.~��AU��\m�j�����񽞡���V��e:[.����I;*w�2�ʉ:����I����i<�m)I�k��qO���x�s��;mY���Q���P��E�,�mc�o�u���Y��r]�� ��_?��>�_	h�毡����}�E���yÍS̄�L�:�ѫ�S�v��1�t��wO���3A��_pQp�)��S=d_O��Z��m`A�7�L��)�:��K6sG̱2I�L[X;{o;͡7n��Ӡ������;�A����2���5�x{��ͺA�AH��̢c��`�4�j������w@���1� 9E��ޥ+���-e.��F&�[�֢�f̽��l�l[�د��0��� ��]��2w�ڹ�OQ�c�%�o�k�m�k�q�#�*���Cf�f�j1ә��<¬���t�,e��M].��yѩ�I�I0k��?
���-`���f�~U5D�b��@����=5BD�b�����ϴ��w�o�8F��f�jQksҦ�oU�w��K,���"~Lt�-�|3:��Z����nU������c�w!�iu��DF���6�ʨ�u�d��q��=�+\v�t�bz�!ȫ�n��+r&ɬ���x'�����-�^je��v�EC��Ep$�*�"C�j�Jf���P�퍵��T�a}^��}��O�[����;8�Q)
��XG�teˉs�z\aQ�11M&źO�Wn����*��ձ���M.�/��7rq�iBW�ҿ�����~����/�B�=��van��i�����o����Q�����(�������4�7Z6����%ZJ��w[�]����c;2��	w�|�$��gd���i��I峌��M���ݱ�P.���b�3|�le����1�k�|�y+il:,Z���:]��6t�_�ҩֱ�-ײ���z�1��nc�ѠH�yi�P0����m�މ��|�J]=!쥡U�v���X)з��������v�-�y�KE�d��5%�(j��;�[U��՝�/�/��}���x�S�e�;����}z�7U�����@{�0,���)i1z�gpSl�C�e���ҹ��r;k-�V,�K���X��r����a6���*!�j��_p�0�Ȟ�<��C�Y��<��	���(�����z��m_��ִ]B}F�L=;�R���yő�(���O������;�+s/��{Y�9s�;\	�d�T��:� U�8�n5�9U�������_TK̯�)k�c/6�}��h��Aв
)�UN��K�^<ž�yл�8j�N��'�ȫ=�����뺇RRv��l={�x�4B�ͫ�%C��{� �S~Je�Uf��J��	��{ޭߖ�q���c����y����rt�+�:���:���:�D��]pwrL����2��Ll����~�0��ܯ��o��N��^�:Aaͮk7 ��vv�d+��T�����eKˎN5��Cj=�ڇH�1v>��M~g�f�獬�v��8�N��>�O�GZ
mk��v��j�$��{��Ap�ǡz+K~r���-�ίE}LΞl[��;t�u���▴)D��������}LwW�\E�ݥ	\i���8��Th���5�Q�FV����r�����9�H�<� U_W�J
7�����SY��uuKc5[z��|Zy��� P�@l�����= i_�;�ū�y���N���yѨԞ�>mㅵ��Z)-:{�ыo)�inu�j��6�����n�M9}�	k\�^��r��W��OB��&�V�Ū;2}�����F�W�gR��nZV�k܆�E�=�S��+}�N�dY�,�":{�E{'W<�|�1q��&�� G&���9��/����%!u}�'`[Z5C��Ӕӓ�]]k2�>�w�姺�}��@��>�c"���O���r�b�S]��*Oh�Qѷ:�3��<��]I,]gS�9v��Ս�/�{`��x�{������^�]j`pf�v^p�L�y:*���p�m�T;e{J4�z'�m\o&�^D�d�2VB�K�� �R��.7w�Bo��\k�G!J&���N�q�k1]������ݯ��g"�ws��ڨ��j��i���vDơ�/�Ov�]p/$��hQgӒ���R���_ݢ�u�^��*#�����v�f�EzM�~��!�ߋ ���@�#�$�����?t	z+�;a?@�Ю��Щ����1�λ���{�5�F�S��X*Y�~¯Ld�`o��#�ˍ �1켩�l���3t'tú���ӭs����W�K�^���B�����W������#܎8SC4���i�4x�2���.���+K�6�J &�J�}*h)'����E�D�x�OJ�>����ۮ	{i�vO\EωCne�=P��U#���L{ܧ&�﵅5��|�R>�̠�o�Ķ_���.��-��W�z�óG� ��g_�� �����_�(��`~������ПN�M�w��߶��ӟ{��VW�ǖA��P�a��q����:NQ��U��p���gl�Uy�ٔ�[S�SU��eMOT]���l\�3y�vG�y��-�Mu��h��*V�c�:g�=rv��E��⺲�9�A#���Jv�<RrF�Qj�;+�΁���ג���]�u�{�R�2q]�'��E���/�\��,I��z-ee��;�����zX����=�:�h��\�x\Ӎ��09f/ƚ��/���n�f���/�+��=/Ճ�����ߤщ�+�^8<��yyW�6t�*��%.W����c�as�&�J�z��"�_�ī�]��L9��%��A��9=�|�Hq7�T���T�ә.ir<H����nKG���?k�uWt{O�{�O\�ۯEa�ѾF����m��}��=Z��z��s$�lԶG�*�хWwۣ�*�o/�W��G�hR�o|�F�����O�>>'<O�3Z9�H��g�u��3�u}�B2��[��/&�+���`���f�S���K����z��]ɋ���2m�}���F�����]��]��[^�4d�iD�0��.�tO�ތ��׸�F�1��1П��\c�3��x�v
���� �u��{jA�����N�>�ô����W���o/��n�1]�����ש�_�����^�̼���<n#�ڱj�e������Kޑ��ڋ]iZ}_1S��-
��N��꽳���y�A���WBA֥
����qx�(z��W<!^dA��{�D�|���<ӫ�*n��7��H�9RVCu��'�s�qhwT�f���'�N�)�y6i6kE,#;�����]]t������F63����E����3�ڄ	���R��6��Jձ�O����u��;�;z�8_ЮrN\t�t��2����s#|d�r�z���Yw�y��m_�>�S��r ��-j�������w�\��y�%���\΍��:w%\��(���yQz6��w�ς��v��>��=�,z]�9~>�-���M\wc��1Ѷ�:�p��چQ�/Ӈ�g	^�2�P3��I�;�[������O���z=LnG�^�Qq��j{��V�/r�I4���	ߐ����K�Y0��Z�ؖ�U�u�E%�!`��z:���!� �c���`�ǽʈ]q�Ǹ���QD�\��Lp.�#�	O�m���x�<��K�7�{�ΟM��7^���[ӟ?I��u�ߵT���S��U}���I`L���������0��'Ʈ�׫�Z����\M����Y9⴯�ޓ�_��#o�L�|�Af�PB+ц/:phB�=��x�lʎ�=��H�bu�ʐ��׭��޿3���}�TN�z��B��Ԫ�2cʃ��Y�W��r�ş*��c��=�42�����{|�Fw��<|�����;�_��myvg�M��؞޹P�;M�+�0�����9�R�����zV힋�9�y��z<��e�ۡc�4l����#9�RiĞ�"V,�}�̌�L:�\�8��u����K��rp��6�8���s�^�:(e�h�{պ���_Y���[���H���J��~t�W��vU���;dK����k���=}�r<.�܀[캐6���W�|�6tOp:�G�7|�� ҖO@!����պgJ��_f����tq���O;4��u��!K}��uro=��~��>�����ڐk�>%T�񳳁]z�O=:7O��������He�[9������v�\6�U�F�P�g���b���g/���|rXJM?"i^{{���kk7��=���u�o���7��7�u��g�c��Wx��]���?^�m�«���?�ޝΟ�֟�o'�����C�gG��(�����`+�,��%��xT�/�������|��G�{M[��V�w��L~����m�N�1�τ�E����f��i���񐾦�~�z}#`ǫԱuR��/��Ѻ}�H_ڶ��ş������C��U#����Tm������ItQ�&�G�;�7=�_��9�!��r�W˲�mI�W�A�P�"�nFD����ov�(�ܺp&������W��O�܍��򜈯:�윜;PU%���K&�tG�es�o�<X��m�gl�m���1��
�=EP�0@%��
us�:
��˳sf��jm&�D]�l>]����ګ<e�t)��,�|)�]���Wƕ�Z3g�7�9�%Z��On��J�64�2�4���rٕVW;�to5��ɬ�Y�Hs]:�H�6 ��gn�a�p���5�e,�ju��'���(�`�4�U�a����W�s�b��a�nwl��C�^=�Ã��0V�V_&�Yl�X��썎��>���������Lѕ��"8��>�����
Hj����W�q]-r2�a���4����֊T�	Ƒ�}B��7T;ϭ�*
�k����2O�ۭ7ʝ*u���,��6;�A�!/2'r�ܒ;�!���4hp��W������k*9�> �9V�E�\�a�,�x�8䣕���|a�:�.�:��WQD��̫��'��ðV��l��Ԟ�\������}��4��x i��r��)Y��.1]]��Cr�ZX�j�.���K[�H�qպ��T�kDc0����[�Q�( N� ۢ�..��E�Y�����2���,�T͊R<G&
�_��B��'p�Un9-����Vu� E@�%SvwB����x��B�P�I�;o.�wr�r������9�T���:��:��|��k6�Z�,�o#�f�\k���YSE>a<C�>�q���r�9;]�w�g<z�/��9���7]���
Ƭn8&aL�7��D�Z]��/
�mh=;c5ڈk�W���n�H�Ք�G7V��CK����bI[�+_+�su���pZ�w\X������|���(����+)�KSJ��ʵ[�r�95�=�Ke
��|��\��n,�bqі�;�ň�I��9[V{/m�.*���<�ˍN�˴j+��t!vӕC�5�
���+�C��A��4������r&�`�K�W,=5�fW7�hsQ;��m>���ph<J���wg3G���7bjԘgBJ�����{xnu�����̔�u��[���6�T�c��M�63{��L�Sk���C�}�|�x��f�^`_	�Em�#5�S���l�S)���5V�������0+�1e����X�|�U���@&�:�5*j
��a}�&d3�=��mq��I�b�\�OT�y�����s���w��j{<==N����ϊ�r\}˥K/�"�[C/FVU���k�Y��ٲ��gU�X��x�n���8-*�ɫh��g	�&���զ����;�X��}%X�tP8�-Ǳ��qWNmU���k���۵�ժop��t�IK�(V,=n<�$8U�[x�M�V��]f����̙3:����$\�&.n7�P[y���֎��3f��$2�u1�׹B.�L����w#�ٺ�T�vZ�U�TR&%;K�0�]�7r#��)����ّ@�_Q={wO;x���;�Iv�ѻ-�3	80AMU���BF�g#�>Q̉$�E��GD ����^{�F%U\�:h��Tm:\���I��DJA"�3�#"��&ʌ�h��dV�"�Cm��6UȢ�(�LM*BR�Eb�%%Үd�f:�NH�a\�J�6r��Yp��+
�-*�kH8qi�r�NZ&�)	3�)��URiadEB��Q���$�G���4�ԽJQ-9I"��IX�j�AVt3�Q��w(�"�D�g(��5D�wJ�B�jE��^bdT�jA̖8k��"��E*k4����&T�Q����Z�*bj���uU�"T�9Z�燚(�����YY��FfHQILR%=�ENd�.�Y:��U�3-l�R��'**�)���D����S:���V�T�D���ҫ�^y��T�ұ#�q9baUDt̬.]:�]P��e)`U���Y�E�Ǔ�ϟ?�{�fo%�����yJ��������k3�f�\��j=\zLVl��n���nL�cF>R�V>������s��
�?�~�*gvP�WE��n�M��߸生�7��j�z�3���Dw'�u{r���3�x�=UJ�#�U��(	���f�K�c]o�G�ԅ_�ֆ�o�m�):UǷ��^~K!Ď��6�}��cG���|.J5� w������8ٝ
���=>tǎm1��>�r"b�u�x���?V%�g}A�>��9��)�A���^���]-v�u�Z��"��hW�U�𤆘3^��e��:<O���:=����3�`�l��"b%�z��)h��eS���k|Q압6���y����~�{ޤ�<k��C5�S�rf��xQ�~6T��QK.���J����+<�y�{�Qħ�o������M��d�G�����߸�&MGL3Ӟ�c��V�nǒ97؞��s���Oi�qZ�ؼ��|o��yp�?]���.3���=��;�;��3쉪���9u��͙GȢ}Q&��ևqS�:-[�'���?���xcu��ϵ��z_�ф���y�wS(��7�X({�yS���wA��N�qY^�u��.� ������j�*�t�7��'S�F}��b$��lR�ww9�1S�
&�ҫ�z��elԅX���e9�ܹ��G�|�e�Θ��VL|	�p��b%���z�L�8�M���]�C;fؖ4�Κ����I`1y��ejٷ7]~δ�p^٧�yx'�!��ޕcp��6e)�W������R��T������&:ԅ��ꉹ�*
_|��_Z.-�eߍ���|Jzro� ���Eϧ���N�N6��^�CQ�=�s�Pۙxh�T"'��K�^�{��{{\<����Ҩ�G�3��o���r�}�������+����ӒtS$��b^�
u��JGxf�y��۩���_�O�����z�Ƕ��ӑ���W�ǐ7�gl�MOM�+�ϖ��=�gO�-I�A�Ah�\T�^9k(�t�X�k����zX��>=.���.�u;>>WۆW�(��(��;�M|�W�-+��V�FW���y�A�׽�$_ާ��8�'}�f�j���[�T�p����::UǶ��6��;+���A�e1�����X����)��f�qSO ��&D��A�
��D��Z�;�z��}��ުbY%�B 揤������a1�s7�4�˱�<����f�Z5m��9�����h>��@�p�Ih�-�?c�ٗ���x������4g�-͊�R��Ч�7�F�n<��Mǽ>D��w����6!ͲE�C]�āǠF>߃�Up�Yݨ�ʋ4���J;8?�ȶ��`��25Vgggk��8'�+� h��oV���/r_�Al�z/nS˥t�kסj}�8&:���T3���U�@�,=R��uŗ�<zT�7T�o�2R{��KM����:��ұ��9p�? ���fcU���3Cc/Ը�BT��s�H��+�1p���/��7�'�'i3}��t�e��T�B��\t�t-Wl��Y���0dV��Ϸ����w���?]�����&�ow[�`3�t��
�dt��Q�ɇ�wL.�V�_r�~�ʂ#n�wzVY�g�|�W���z����X8v�~���[B�ؼN:�~0�:����;{���6�w���\�o��T{.}L�)���_�K�����kSΦc�С\䜿�X:v��xoԗ9��2��.^`���{�J���5>�(��e���o�ǲL��'!���g��^�G\�
�S�+ήtU
o���u�i�+�82	��>��~��)�X	F�~�_��z��*Z�ݞt�9*��SS=䊛߶%�[d~P��ƿ*KRݠ�܂�.5-�����<��}VF�W�G���=�hٵ��-@�3���ph��*Q�>$�0�ARĒ�������U���pTLϹ=�
l�U�<��3��#�{�Ǹ�<��"�[0��Z�du	O�n`�S�gH��~Ǟe���ѽ�/>��U/t|��[%�k�N�m�������B��z�up+zBm.��sK�}����\�s�6��������]�˒B��1{x�����oe��],:��.���u�J�Vs��t]��P�
]���E�^tiF�Tapl�)/\I^�a�9>s���j�n���X��5X*s���#�z1��+g��DK��t��U?+��W�#��w�q߽�:W��#;�L�G�d_�_����f����{yoҨ����lt�7C�E�5:��c=;��w�L���z�tT&�h�Xt\�ޅ����YC�$t��U�(k!}H��LGޥ��χ��\�����1�z|��������H�����IP.4�[%����18��=p&az��b��z��K]7�S��s����`��2�a�v	�H��d�_���*��Y=���z�2_V���^=}�|��0罛�g�w^���=��ԕ������}��X�d�;��`|t��U��u>��;4+#}6�x��;x֟C��)E�q�yp���9����g���yt7�ٜ��
+qu�`ӻw��މ̮����=u��
��Oޗ�q�j��潦2�Wx��T_�^�^�߉��j�=��z�p�,��;:O��:���x������|�<3�{ߗ���_�ҿz"G�VM8|���$�3���w�u�� ;�u"]�����<+^+���%i`��{ʮ�)vΜ���򁞸�G�\��r��/�i�|��nmI��p����y��֤<c��ʋO��6	�$����#.�(&{دk�d�"��Z����s�uf�����N3���`����٘yȱ6g� {��i�Q����+�@���x����y��;�e���|���Ȋ�!�r���[S��ωJ��< ����R7n�oz:�Q���v���};w�!z '�"�l��/�ǞW���¾]�#n�xԕ�
�d:�|ج�k]��wٍ���\	f�5z�w��W��>/s}p��"+μ8��P(���I���,�G��vgo���c�vLg���)��WG�[�����G���#}!���ڮa�e�����S��=���C�* ��
W��å��>���_�
�W��z�>D��ݑ�%�k���)����ɜC����"we2T|���qo�q���>���G����^�[ۧ�ӽ׼�TՁs���q>�TN��W�&���z'���W���t�}��1��m{�v=�jf���l;qs3^�C�ܭ����>��&���p�\K'�+A�ٳ�D�/��MC�/_�zu՝�=~~��������zJ��Hdx׀�f�R��,�f_���r3����2l\<ɛ�����{E�k�N��|u ���D�(.��]p)����+�s��$32�kP<�)��#�.�w����m�����S�T1� D�)C��d�E������uy�y��j���R��6�
�޾ŉ���DX�`�O�Z+*Z;G��q���n=�?;�7�x�>���j�\�V6���·��W����a�a�P~8�JӢ��~�/J�yp���v�k�O������8s�F�b��R5۱��+��c0͟3�U��և'�pj�\OgѽLz��xd7^�Q�����X�z����pd����Ղ�Ղ�ü�á��/!;��Y^�f�h;���=�hQ�nn�d���}��7R+=�����g_��^/U���/o*F"���0���wYU�����	�}�f^��S5=�.�+� b�
<ܕ�:�]9�n�,�{��S�z��C7闄�s�F��o�{�êxe�+���r�y������=���z��W��vG�Ь��:�S��lѪ��[� �L��&~Jt�Қ^�Z����������7����{��T��{�mw�������ѥq��F�Y�>��W�PE��T�s�YE�nhK^���774j���YuY��G��%q��8�uMj���Kd'İV�FB���c������B�6�74�O����"����}�Mܺ.���{nFI��w����$fR
��^��S�z�y�r�6N�>���F�6�n��n�w�:q�g;�v�=`G����s���ئ�F>��7����,�ފ�X�du.���U��-z@���'��tql]%p	�j��7�p�^jXL��W���my��Tt��m!:m�H� �\�D�@Lp,.�Īǿ'�f[�)��U~���{�>��k�D�ז �O���{ԇ~�T����9��sP}$,��J|���{Ϲ�n�WJ� }���v��oZ57�l���������|�s�Y$�l����U�:=Pn�y�{Y����T�Y�R�#÷������5~�q�O�>9������>J0Hɮܼ��}�pz���(�j�%p:�T�{ƅ���q����~���w&/�߬�3��v��==9�ۜQCp1��eْ}�,����O��K[z2�׸�F�1���0���#m���V��S�2O�v�3����E���� ��+~0���W^��(�>��	>��~�ӷ{����6�`�+��~����P񗑾����V-^T���N�8��wj��*��&r���%N�ʼ�GƧ:_��_�s>�y:�jy���׹���s�r㥃�J�1�z�T��w�ڹ��ۏ>�����ZnJd��v\
��Wȓ=���w>�^��P�|�G�@tN1����X'-m�u)d@~���$ܴۡר��<�^��b�dv ���.�Ɩ(��f6�\�n��4n��u=�-��O;D�9��39}�lSl,1�N���bv�`iwfʎ�&��j�[���춀�oV���G�E�xk�3�c֯��V�^ؕ��Wb8r%������:S�����ߝ?��x�
���U��k�4Ez{��1z�����)_�X�x�u3�z��Z���4�����W�i+=Y�S�����KG�^�<���O��k��|�^�n��~��c�તΌ�V)�7��y�J�����z3�p�3��=����9��X�(�,��À<��ӭU��~I���fz��}~�����\M�-ߴ真9��Q��L��TÁD�R ��V��)��L�*��z�����X����U�G+�Q��z�,��ZT{�t�o�Ftzi���X-l�{����T:v}@��3�=DLO�\��~,n�:���R��m����_������7�җ�߻:�v��]_�k&x���d���DĞfA�<�"ì}r6�数�{�O��>W[��y
�9��y+�[��G�����O��-��,���F�Z�J�������&'ޙ�tU��k��}!$��?9�>G������\�JY= �����_V�1�,B�f:�����>��1�[ �,���&m�o��aGn9����5��\��
�;�OCr!�٧{x_7��Jp�I�[�����g�}��n�s�b��Ђ�%�ص=��:��|7�O(����}�Yײ�r�J�^v��׷ȵ������������m�c�x�@zn=��}��X��Ԃ��Z���f+��w�����z���n������R��u����w�5���������,py3g9x�c[��^��G1���Há�l�W���+����ޗ�gZ��DK����O�]��;�p{+��[�p�j��Ka�g.5�~�?��zg����>ѳ���9G@�?�ͅ����,��K��ef�n���Yu�J����y:�ݑ޾F6�gJ'1��'ȱqY5��4�,��LW,t3 W^��3����^�G��ⲝ!�_�PQ�jx�Y�)\���s�k����zdz�e��vs���+�R�3T#�{�E������������'+�B�\�O��s��zݘVO������2}�g<z��>=��wz��=�|^����NEyׇd�pW �+��mQ��
��x�"���MS��P$�<�g���>j�-�	�n��<���9��K=~�p��'�j�1�sy�ѓ�0zٿ`���J�-�3�}u�>�J���CC{�|v�_V����0��n�7���Y�/��ٹ9��=�pž�`NP�/�-.�=;Eݮ����s�O�Z�A�#���r�q?9��%8��|�`�/����ؙZ�%p�[�6���}�{k7/�&U뚮ww��J�]2�NU\������2����j��gl��<tߣ���}3�p��^�N��@|���P���;�΅o�h!\>]��>�V�r��W�{�U���R�o�������C2Y��D@n��1?J�u����:k�x��b�s�>9�ױ�ܳ�~��F�d������R'�����\���9�L�6v"������W��`'i���on^yQ�S��^Dr�~7�f�m5~�~���	�|��
�I����g���(�Ǚ��r�����v+߲Mw����&�ݞ����q��w&���2o�{�{!��le��P�g.Q�w���<�q���O�aM�:Ü�V�Z��/7���WP��W����3�q��#�������n�� 羄�l�{��>%W�&�Z�Y��}������	W��`��f3���O8�%��������b��N��ݳ0�t�ج�q�4�A��m����)G�w&o� ��=>�^�����/>^��#�ԅ��H�R�ݸ3A�}~�j�*t5�f4�~�rKs�����y����VE�*y�9�:�]8ۮ#�l�>�X�ȿ�U&��^>
\�j�]�͵�+�Kˬf�:[m�R!���<��,2�����[�B �Jݲ�X��.�bm]]FgM��)Ǝ%xn��O����tdt������յ�5w`� ��t��W��
.�f\+!om���̙NQ�6:���:֡�ٰ (�ua�6l����ǚn����_$��|f�"��BD��p���:�
#��5;�zh����w���9�$�h����f;�6�юݤZA{C۞�{���T���,n��|��3�h��%���r�9�}�:��6���ݭ�5Ñ�liSA��x��LwN�6Iu7t����*�X�>��w.."�f�E��Y[�.����Wg�4�'��2��_=|�J������Q��!�\sh�`��&^U�x���s���������5���X5���0���@M�t��,�C�A��דl�7�P�K��o�Yl����V��ծ�к�����OmMB��L��=��Un�m�o���*�e�.�q��R�he%+n��&)SB��Wz�w��R�$ou;�g�_�J4(�֊�CNq��C��.���0gd��qHÓtlZ��
o_}�򌝽M���@'&� �Q��Y��R�r��W��v�M�[F�V=����� ��[Y6=��;�Wu��T+x�޳��������Jb-��X�mc��9��2�K3pI�]��v�Ԙ�5�)vg��-z�����Ccr-\�T��ꤣD�U��ian_V_`�y}G\�����Uuҗ%E+(rY]�v��������N��]��\bk9R�x�b�6uǐ��r �u��F��/2w�N��x[�{ϋ�x��[��K+�wE26ei��c������T����Ze㒯zCg�*�8J��e��q��M�녚�/))�v�5��+f%�bݿn��C,�]R��z�^��qk�3���c�/�xQ����C�ͽ`?X��=��W	���}�с
�1f�4
���p�.˅��,���M�Z'}˺�Ks��u���k%\�o���N|�^,�ܧ)6�g26�^ˮ�w@b62p��2�#2�Ԭ�O�Q�y�Mbΰ�xx��ٝ�Һ�Ӿj+|��:ެ�,vP}��	�ۋ�Tf[��Ê`�'A�YڻREk��֫` n�y[��5bZ{|B�����u�	t���cѯF<���:�Z���&��Bp����ug\��]]��/к��Wv�X�c�->N�@(6f�清� Z]\�^�N���-Ֆ�����6�J¸�[uh�om]�YX��� 4!(+"v3f�*�C����II��@�v^u���E*n����ւ��B]�)��̂M˵��H]�)}����f] ��f]�:\�[�<�Ӭ(j԰k�r���ke<T��m+S5z�s���#��{7��b�$�2
$�J!@$��*�W�M�кf����*Pz�DQ��d�Ą**U��̺��&�r�U*��(�<�)%d�̩T�J�Ef("�C��8볢9G���u2�E0�\�=ۆ�E©4U"��(=�qdG4k(�g9p�*�TJ"�FE�E�*���.UC+Մz!+2,Ud�M9��0�g2MNEDr"���Q\�L-�eh*%
�i!N�Eăh�z!D鰸�$�ˑs���"�
��$��Z�J�9U���C� U���bi��*�0�iȳTT��*K�QAj*.EhYEE���"��f�Qbt-�TsՖ���9UiJ�D��ah��+�ZdU\����$�9F��j�򫅘b�H��EfE�F�G*焅�Z�e�S�U�j��(�^t*�=NAU*W#��Edy��r��W����p
4�U�{
�`,K�U7�vd�t^T��u�odY_�F��Wڻ;o����x貍NCD��dT����_t��mG���T+��F���<�GL����-�����&T���y\+��`��X�q�Ŝ�ڗ3�&�q$�xw��\EL�L\u�����<�ޯq����{��W?(w���.�M�4z:�g4׏a��I��A�,_�*��}k(�-�	�k���z5���<��vH�X0��oI㩪���3�0��F�GĔ�H�Ge%9�uѥg��럑s�y���vl߬H��;я�^eo�Tt�����:�b�_" y�n���^�rw�3����T%Uz3��{�5���O����ב�zxi+�o�G_��&�̗5� ��v�s1��]\�c�g#풣F��O*�l)H�X��TkF���[g��x�OV�~�����Ӟ3�0���ؙU�H��l���||jy���D�Jt�]*h��
_���j7�W��z|���L��i�|�M^�!T�{oR�s�G�Dd߉�= ���V
�\����K�bT��G?T�[�g0��5��^�؊䫱��6�;�`kbc#K�$�d�@ɇ�'�b�%������z����Z����+�k3�)��4(4Y���r8��S�P,�!����wz�6&Y��s9����4C��M\�	a�L6�ճr�]��_Hs���#/��r�5�#���/[��lm�и�Wv�&V̓��0����U+����m>AM�'sV�ʱre��J�G�ޠ�oޟ z�{4X��ԃQ>%Pɇ�wL)�����Oo�����k�r����1�ݷ��y�y��2�}x�{j�¼�{,���x�ψ)EȰ�K5z�\f�;��x��i:Wx��W��]W���:�jy�PQ��g�8�(��O�U�<��}��ܯ0t�D��GgG���M�K�(�.�:�g�d��;��y�%���1��稩�FҤ���Na��𿒓�n&|2��u>���])�ٖ�����y���1i_�Yg��z����碗\wg���1�m���Kv�|l��K�Y��yu�/�����^��}�����tQz Ϭ���܇�����!�s�.��v>��=Fa��A�L\T�D9!�Ξ�����W�*.�A��K��{>�~��|�?u�z����
��EI[a���g�7x.E9��U�;�z�>��3�V}j�7M�Ė��|�����|oڪF�Ω�`�*3�`��O{�-������T�s�
�����@�å2�U�G"����z�i�3�+��N_{}r5�d��{o"�t��w�5L�[��7��Ρ�HHYy��ud�%��xȫ�9�Df�-�Nv�f��B�*�8�-M���z�P��3�vT3�P���	��΋5�O�&��������������yqX}�N���3���R/�^�ݠEo�'-�J�3�{��Qzc3��@}�O���n���X�Σp�R��m��N���ݦ=z$���H�*0�Z'��q=��K*L7�:��+�h]'KǷ�����R1�n:�M��ՙs�GR��}�/l�_G�����G�����O������`��QU��M���x�+ۮmO��+%e]y��w��B��]ȸm׉�G���C7|�� ��Y=@�|G�`/����_�ܽ���4sr��>������q�k�~ήM�?P�z��/�ڱ}�ck��/���_��vx�
%T�������뮭�{r��v9K�q�yp�]�ϵ��������orƯs"F��I>���N4x����A��V6t;���ۈWO����o:�ǲ\״�B~���2�>�]U�i靖q@A�D~W����~3�����|?F�r��4��;���Q{��pDf�W��"_�&����p>�WZ�Ͻ�ݝ��cj�t�,�ۈ3*�.+&�٧@y[`�X�^֎�����n���ը��Ey��z��+>�Hw�3�gJ�>% a��=P���	��Hڕn֜Thg��5v)�Ifs;�hIί�����-�I��4B���	�B����<�f�qL��˜j�u��p�Nm�ڷ�c	xx��7���V.��'yhu�)��֛0���Qd�oa����A�#d��G�K������,�rЌq�]n�h�+�����޵@s�5BctG|�Ss��c�}\�D�p��R6�Y'�����(��B�Wٛ!!�0�A��ۣ=���Y��[����^��'�����:�순�
�Rۺ�����b��ʋ�o�J'@�j��Ks�֮�7MՉ�n��#�O���,��,������q�Q>�{���d�^��D�}p���X�+�o���a�Nx��<+������́��^�x��\�/��G9:W����f�rY�����IJ�@��r¼����w�}�m�݃�����lg�z�;b=�\U������<��1���%�A��NI�1�7�K�\�̮�c�y������k$h���J'��tx���\���9�L�6\��x!㫭�opΔFd{�z���)H��+�x�Gy�����Mǽ�@�#Ƽ �d3Z�re[�_l�_��Wۚ�qv}d��E/x�8�5��9q���n����n=���M�9^&Mǽ����{u;7W�{����<�����s���:ǧ����{^�ާǝ]C��v�8���Zo? 2�_��Y��k���T��/:�m>�ɬ��fu�����ոի5��3ͣ�.�ӭ�:G��䫟)%���Ɩ�����.+�1��
n����(~�.��%
�s=��������z� y���9��G[Msت��J,�g�� ���د���T����{f��L�>%PɆ�ևu>Ӣ�V��ަ=�=�@�i��n��w%>�vL������P�K��X+}X6��0�����������V��ڙ��m���R�����s>`߼� +��+�ȗ^��z���/U����B��e�d��V���>�t��<gr�/�^�Ui�S�Jφ� bj��S���u�s��pY�h\j��ܫ��S}�j͌y��Ю�-�t2n�90�^�F���<�GL����������#�p�^W��uY��\��s�[uݼh�����rX�E��z�g�����|�/�B\�k�Xqޟ��G��:�8��`�YY�8�Y�̑��'x����P��+%>%�_j�ҕ�ֲ�2�Й��6�ҭ���@�e��Vf���<��1�������3�0�5�u|��>%���>[��]Fdo�j���x�:�.�),�J��G�O���GJ���˘L\�P<��8y���a��\�3x8͹Y�O�>���|j5~U�=^X�9>G}����o�G\G����2\��G/I��iۮ3�*�?*^ߓUy<~�R��97��3N�K�ם���b�R_`��K8T�+yƴl޶q���]/��ڏ�x�졀'j,�h�nΩ]Ĕ%�WoI;��r9��W(ӹE%��i���;�:�E�����
�z����#S��㓫5��/�ֿQ�!R�|�çȽ�f�Q�h�s~�ˏL�x�ޞ�������%:λ��uX=xg�2O3pjR#���Rt��á����m����x��>�~�`�鋟)�6�5%`�4�[%�ޛd��zA0���D��NV�]/K���ݗ�7ʽU4�aJ��N�Ǘw�ɿz}���lq��'d�a��'�`���k]{���T��]�ý[>ۺ���+�1?]ȸ�~��oޟ z��E���ԃ_t��C&X��
`z�n�[��M~�˙�6��~��G��~�V����9�C�^��=�Ջ�yR2�Y;���bߪ����KS�˭>bx��G���������K�Υ^
%�{I�N�Z����חÛX�W�ګ��JVxw�K�)�t��ϰ�S��L�x�"ˀ���{"\���;���1�G����ݕDO�f�k>�2��߉�yT���::���	My�ܮ�&������ic�uzvU���9�{p�>�בY�qݏ���ƭ��q|J@�x�b�g��[��N���	p��5)3���Y���K�4�N�A�+�)��MM�����I�m����U}��xh��'�ۃ�1R��3��BdC�q��\Ǯڕ��yG٨0%�+�X�x��]�[��F���s"*o���+;�PT����K{p>}�Q�w.�Ⱥ�!�����z��҇�Bw�nSz�)rK$&;�V�3��`Ah�\��s��]W}���^���+��!`��z=���~�#�~���9��X�(�"�
ѝ��)�v�k�-1�������P[Q�F|������뉹n��"<���g��!������q���xL[O�}��\+���9 .��O0�p:[/"U�G>��q7��֑�s;��{�t�oށ������Z��"�"��\f�̂�(!S� �<|:_��/zxj�RF{Oh�x�sgJ��{7�R5`\����{I�{�ޙ��,��L7p:��+�hJr�v�x�ς�j_yC��׻Ԩ]TפW���c>��Y�Ͻ3�%�x�l
v�&��'��3���/��n���Qh�H��6a��cs���7�~�����w#��UH��x�g�3�;��h�� ��Y=P��]�����xih�T�|ƨT,e�=�V�-����m{o�"�\��~�=7��~��ڱ}����R�)j���v�x����C�������?pu;=�
5�^��`Q����g���B�Ă��VF{�2�������]c�B��H&��Z����V)k���ɘ`��gm�U=MR����J"=���[ޤ�[���:(��4`nVopW����!7H~ە��ğR]yw"��K���b��w>}O;F�%�H�ΏG���MD�c�+��?}�vg.�Fa������WO�㑽/�:�G���i��W�RK9��5u}Hv���cɜ�G;�=q���
fl�>;;s>�l�w9GE��_�܅��(gb ��:}���n�V8�vy�ߎ�Õ~���S�(��5��6FW��y.�kN���Ej�Fo�w��SFjo�W���iK}k�FE7��9�~+)����Փ<z,����<5��}���<���T���W��^*��棍P�c�-l��/�ǜ����9\\��0�Ñ��1^�g ��̓�gW�^�ϑ����%�n�o��^���F���NDW�xrw�Ƣ��
��=[ў�y�����x{b&P��ȩ��Ig���7�߸�yI�|I��P��=gk/�����~�=��/��QP ��2�����6:[,>����ԅzMdx���z�=�++׬1��[GȜ=��D��Lø�rYP K`�ž�.:ey��[^�f�{ƲMV�@�R����>V��:�3���_�o�K������7��D�K8���D	�c" ���zf]养�n	�����FoN��s�WN�8k	Y�P S�����'�}�ðd� `v�w�1w[R��T�g�uI��%��e*��s�q�u�+ vA:��R�N����+|��E�N��$�
M_8�����Ե��;{Rv� �����|�Yv���KtjTz�V~TW���hu�5�����<}(�8���o�{��_��Ng�*=�7�;��:��A{Y�����"buS�(�en������΄��M�{ޤ�<k��|�hy�ҬOi�*i�h)�X�>�3��c�e�pTਟuh�˥��R/J���CU^7�9^&H��$��ӟo���#H���j�x�&M}��(v�=8ԭ:.+__��oS�s��s>��\퇔=WUVz�w�+� S�1��/E97����훎>�8o��U&�����������Z7���ٞ�/olߴg�+��^쌍~�ޗޚ���X�yS�����0��sL8؞��u���Y�挤ߚ>�Y\�� E�W��׾3�{��/�����RyR2�K'uzx��yť�~�Y������pt��T+���pj_�X6�TG}�����1t�6���=
a��/S����΋�t@�n&tO�f:T���0��
�:d�R��wP�OVw��F��9}�Ή�+����4;�h���']R\?:	h�i~�S�З7��a��W�=���{c�=J�.�T��z��ܮe�:�'���f���璄�fH0�+��셹TlуɼD�l�2��y�P�<Xd^U�b��h�<��jP��۝�Fu�[Y8���F�DS}I<��=�c�)wv�mb��a���S�%u��=�@DN�3��g���q�)�W�ǐ7��(�rA����c*U/�YE���bs{7����tܪ��1>\�ÆyS��>YCﺇ�p���P�Mj�_$�S�X+u(S�o���v_n�J����vϗ����~���G�י[�GJ����:�p.K4�����ǣrngw��BuGG@��XM��h�u��F�_��߫�g'��z��}����&pc}�k(��pn�NϨ��" �4zH�����-n�5�����o���L�x���>�C*=�!���F��s���n����GN3,�R;j28�_�
���F�
_����5~���_d�Kt�Q�"l:'����>��)ͲB���^�Հ��47��t��%O����JҊ�op�E�L�C�$�����/����j6+��d��\�C���hK��x�^/�Oް�9U}��9Q��Eז�u����1�	��E��3~���٢��{jA�����#�|jϰ��k��F{*=�c��t�Et�>[��8_m��dG�W��~��/>�^���ڱj�f�B>��#��R�R�OL�e�F*sR�)���q6X�w]]]���d�m1�A�S�ʰPPR��w��!ڂ�bȯs��E�\��9&��"hvi�J���3�t1 ��U�I�h��MP�.ī7�Л�jac� q�7,�]�)�֚�Q�YXS�����'f�5��.`�u�C�
9+�%���m�)67�Y���a�um[x�����0g;U�a6on,;�� o9���`�:�X��\�\���V()��m�b.j��x����׆�)WQ�v^]�A������]}u�c�`;Tk�1W5�*^�d�L֓��.���pm�9���4
{h\���5nQ�_Z�J�Ժ�Qe���tZ��2Uen����-��d̹}��6o\z��܏L�j:jtt�w���$�ޥtw99�f
v�
�5��7g����� :���%�V\r��XV��'5���&%zJ�� �*��y�
$��mE�ONs�_;�}i_S���h��h���[*Xv+��Q:���ki����̎�a�%j���Yj�GS�����c��5HC�iH�����omϻ2��n�k f^������W+Ķ���c�Z����N�㵐��P�f�OX[�u�l��.���+��!�6Ry8ԓ��Q���.`�޶�����+특���Yx�{y��|C��u���ڵ `;;gXz�(9�#V��A��?iIw '�����u�úU�k4��A.�U&�T�l��^`�(�o1�f+��C�9��*��諠�)��֩������:����Y��W��c��8᡺�y�L�޸�M7����B�u��z��F�5�hE����Y�k��z�u���}2:J햕fp&sw�w�bݭ�뜷ŤL���M�e �����OuW(*tT(���mc��[�,e���p��Ml�'�����t.K#�!L{&)���n��p���J�Y<��{-�:K������;)ݧ��: ��f�t[�}<jKF��z���y]Į��\�4�o4���@�1���UkK�\�5p�<O^�4Y �G<�$�O����� 3F���gLq�{R�J.��]��.o+&b�SKC��l�`]r��Uø��4�w�Jt�<Jŭ֦{�V�*;�L!&p<�!+^ˉ��;�k)��Qf���4�hC�XVh�;>wI0�!�Z��ҳ#	7[n�{�D���2�*���xU��ַ��yݱ�,7�lv�-�R�{��(�hݍC^���Ƌ��<��
�z��V���X�������}�r;���[�طB*.�[4u\.�jS���%�:�]�t��CZ��Fe$0]��s{�S�,2��q:�d�-�|���>��1�*N�5j�����2��W��x7�=)�X3��1�9��F�9rзi���uӚ�qm���ӊ��m.EX��p���5������bӹ�՗�p
B��|*(�5-�QD�,���ɜ�d䲪��
rI�	-#Zh�r�r�
(�OQ
f-w!Z�䙐� ��PB� ��ZK�����$�r�šT\��DEt�-Rg"*"!0��΄qGq(��
���$Ei���(�J�5���p�K�r,#Dt"�9z$J"��t,�,��\$�(�\�j]Z�wKL�"s2���z�ZU�����N�I.S3�!rH����XBUh��Bs=

�����z�!"wr�U��RfBs�k(�.�*�Ԃ�4�VbБ
2,0�8MR�M���U��E�� ���(�Ds0����-SLȰ�D�W+0����r���iHYY�YPPs6i�t�#0�3��̡P#B�AˑD
��E�2�MR�	ii)�P�j�4H��0�(�()Xj�YV�Ҋ��jjs0���]$,�2�D�J%O�P�#��iSP�o(TmE�2	�X[ۋ3oBUs���Y\±��ՠ.�ۮ�Y�\Hx^�!]b]<����*�^��,M=��iO�]E����s�?څqY^F�K�t�.��y֯���a<�F�9��������!��v��;�P�=�9'�p�vx����ʮ6jW�Gˀ�ʣ��4�|K�_�C�ɫ�3k�M�&��3�����/_#zo&tZ��;q2�W�g���}GD�#�{fX��К��m�y
>�}`��"�u-����w՜�o�⨥�[�q�V.-/�!&�,^�e;��S[�AxQ^eU��}^[��csޯx��RYg8�B�F�OT�㱹y�'O
�Ƿ��ź2|Ǫg<n���"���{޽�|�?��G�ަ=���*�G��|���sh��n����_Ғ���H�S��V��=�q7��~��O��u�ߵT��Y�5�J�w�EQ��g�F
��l�dޝ��&u�o���o��"�����}INx����n�_x�5���<x���mG�y9�͕�cB:�|Ѩ}Ӆ]��h9�o�ʐ�WH�oG����'��K��xc�:�3���n=�\O_ު�Nd���{����Ȥ�x�gփ�3�N��,��we��on����.�dCȧ���(j����)�WD��������ă��ْ�k(h�t�]�&��}��d]���;��N�)�7�1yGa�X��%�������8_5�FA]#����=ϯ���[�*�Ҫ���vm����k���O��������Q�)ۨ��rz��/_�{*�{�N�L��Y��
��2�ʏ��]7��1����G��ͺ�>�������~ːiK'���f+".�?ݝN_兯��W�[�x3����k�^	��ɸ���q�_���v�W����^���7�](�+����U����ﵰ~g=�vz��C~�㑯��� #7jA�w=�v� ��;�,\2�g.:X(��i����6�]>'�oK�εq�lf@(�z*�sw}�8�P��q:��Gz�_�׼|)�������3��4�{�NQ�f�~'\�& �j�RA�'N���g)�d�����C��^����Y��V;��|�^�T�Y;��y_	�,a�C�>��O^��F��_�>4�z'�r�k�FDS~����)��!���[S�����^S�{��վ�}�j=����_յH�_�<�8�V1�"��n{~��1��C�d�p�gO�O�^�y$5g�xmK�~�~��Z�n������?�VS�_*�wU�s����I�{���~S,W�y�roΦ3��=#k�I8�'"a%%�ܶ����sTU���!��~�j�?"�@�-�yov���e�|��mӂ�d�,pĥ�}R��Q���3�z��v�XFS�;)����5	��SR����-S��ʾ�o"֠��ܸ�z���;7�Z����ĺ�H�|�e���5�k]��7��np?@6O�O�'�e�0<����tZ�,�sBw����}�Z���q��w�Zx0<ϣ��{ڪ�l� �(�( yW�X����a�Nx�ϱѴ����&�(~�^��cF?w���Rt�{����!�5�@Љݔ�C�ݍG"_�"�nz�ͬ^)]^���g��<����z�팈��_�o�K�����x�z�Q5�e��嘸��g;ӵ���Q��L�>�)v���k֮F��2=>�O��������\� m��y��oY�p�ɝ�F�H�J��E�������y�����O��@���^ w������l�����]v�eפ�C�O
3)����Q/�E^]/��K�p׶����J��B��]wT�G�&�n�����{�dp�̕0�M|rP��JӃ~�}~����:��w3�9\��ɞ�?Cn��z'�^z} ��׶x{��>%PɆ�mhwS�:&u��MU�r{b����ʐ��|ɴ����:��|�{�25��z^���W��-�Tῴ�wA��}5��Zq�-��Ы�q�=h��g�$�J�o/�'��h���C�x��Vu��sv���[��WQ�!�]��=������f� ������؎���S�Lm!f���K��J	����9����Ӝښ2�e���G��V����Wl�iQ�cuE;�cF�8*b��%��]l_^�_�s��Q�Wx�^�ǽ���ʑ�6�}S���!m�opGkr���+>;�����M���V|6��5dy�*�F.�����Цvbף����u{Vt�u}��b��눹D��3�5z�]z�������>��o���Cr�}����[�~�<�\K����jE��z��Ł�?�6�:�P9'�c��t%���Xn���Tii���oE��v�{��������=�s�#�ed��e� �.�R�7<Ë�}�K�U�ʌ�3�4'�w�~<�����g}��d�w䢇�+L�zGyu]<�͏.�� �>��-���{8H����ϼ����*:UǶ��.\��%�=�BohL�z�:��]�*�����q#��x���F��\Mǫ�g'��<4��dnk�:f���q���旴��ߘ�l�S� Jt�"e��lt�}��F����o���L�x���U�f�ub��FM�������2KF�ԶG2%����M�@R�o��5>�=�/m����M����S�(٥�e]�P��9���M�f���j�rR��J�CI��ڵ�H�VV�+�n�u�w�u��)��/^�3���X������$���ڪ12r�5�H-��pKً3F��O�A�u�N1+Mh�U�(��'S�A��ݸVo��ԁ%���	�I���K9��w��>f�
�ͲEB,�tR��*��yo�ī�}��������A���e䬫�=>��
��]ɋ��Ԛ���}|�xb��J�rY0��@�1NV�K��w��2���gf�`���K�����_;�gП��c�2�����E���ԃ_t��r�}�^wW�gۊ51���{�|�zT��>��r�v�_�}�U�s_�x����<o�{j���s]R��%
9䷎�8����哵 ��#va�ey�R��8�_��Z��U�'"�֧�2�w�n�l�_���P�o�wnxz�ɼ��:v��<t<���pjW�G"ˁK|�=�{�:��=8�3ۭ���E{p�>�s��y�w%��tU���^��Ib��qS�:$�S��d�eb�͛��2���Ӱ;�qV����~>"=u��SW������jxݟ�,^@3Ń>v�/�>��s�=���||����8��<�O������/����ȯRY�����ײ���#�����1�\}�3�n��
����,�?z�d{���Ͻ�G�ަ=�}9<.��zc4��ov(�V�vn��E2��jg��7�hne��Qc����+^�]{����Eڢ-M�>�z��]&���(��D�J6u�����7i�<�o����2��W(�5�v=�����^��u�8`��늾�MZ+oaX�ۮ�*��>�3^ty�q��l�*_Z�Ʉ�wX��>�+j��o�&�����=�{�������X�}^ȝ�s!zEyU!���) yMI`Hn���l���X�s�w�qW�ZG=9�6,�y�=j�����}�9:UǷ�#|e��24��Q��r�p6:_��:��Y�]���[��U��c	�����c�zw�����{�������E|�K4�a�DL��4.�L�����Et�1y�^�o�HΏ5~g��ώzg|K������B2������E��s�~��(��1���h�VJ]7��xz��G�����_ͺ�>���n4
~ː}�:Ƨ�$�}0�^���c/߁�5��&�2�|�^}����~urq�@���޿��R�46:��{,���ɐ}|J���t��W^��q�/������7�m���o�h���3"����~�` ���WPw�ˡ�Gl�_K9,+:��[5\w��g���C�s��`�X�ݽ�sn&ɜ�g�������Ew���]������7���8n��ۙ��CgC��r����ʓ�wW��ӓT���s� +}Fe�Z�©բ��jW �Rǁ�KT��P��O��[����bCb���P����.�Y�v-�p��n�׷�cF�ZN�`�f��p���u��y����_=�'cS��U=MG�;b�����Ŭ�3ۻ��k��|ɿG� *��#�%��xT�/��ݝ��b�o*t�"�ݿ���N�F}�&���������,�A�@yh�B�k�FDS~����)��"���[SǕ��#5���}�!�f_�;��1�j�C�uH�u���T!\nȸ������1��C�t��up���.����bʑ�Ė)}��R�ڪS�_*�uP�ޯi���yB"n]E�sZ�� �/-�ǧʟ�}R[#_�%�q4�#�T�s�J��-�	޹���!��wN���ff�׭�%'���ίj�}�A�e��Q�*2���x͎�� �7��a^���xWK�}�}+U�V�ֆ��o�m��N�q����Y���J	T�6W���W%c��\ul��)9�3<����z����_�o��.&����q��D�3%�g=���u}�W�
)^�1�ɉ��to���/���q�d��~v�z}H�dxΏ�zt	�8q�����8��9���K�_��q�Q	~���T��ל�������zJ��Hm7��&x�б4�Zx�{�Y9� C3士z�����{9wJ֛�M��͟��o������.�ͧ�CY��/�5�`��B��"eҜ��az��5ܳQ�����簌�����&;��b���4�[�[���g<=B]ȵ+��]`��<��ցQ�&j�xT����/�EeJ��=�R��^ۏ7�q�������j�����\�>��2o��P�f�p�̞0���:���ivk_��e�:dd�_����~׼��͇�u���1���7�g��{Քw�>�8o�>%T�j�ֆiN��{ۻ�'_o�����Y��{H��ޤ=�Ucá��dg��C�/{�`��}z,:��9Y;��Ӄ�Ts�Wݫ{�f]ipw�%�u��٧Z�� _^�_�}.�{�;�w�ϗ����l�P��pR�K|����E.��H~�:N������߫*�������6��5d\����:�]#�����t�]=���S�dW������d����P��e�=P��T���.���@v7��Fn��w�o���Na�=�u�+��m���Z8$�$뤸~a-�/ܫ_�^ROs"*�.{=W�N�n��rV��ט^	ׁ�{G���~��Σڌ�G��7�����X�W���]ݛ���1<���Qf�z�M����C���{�����u��;��i�SW�-����v�Tˢ�!#��S̺�J�m�^�i4�.�	�2�f��3���V�.���]+��5����ֵ5p�%Z��{��͗��ҜTC-���,c쏡�B����to�EE_b���p��Bڹ&uGw���B�aD�M�_�8R��*vh�Cʽ*�L$�n�LW�w��i"�ϗ����{8H��������+cʎ��'D:u�l��q�N_���)��\�������/��J�=�w��G�޿+��W�!��k���{ԇ�0w�h6�����{���E�ElΉD��" nj���끸-n�Q��kF����KvnQ3*��o-��F�e����|�zs�Y$�D��=$L�Rt��á�R�8��+�z�Vn����Roޟ"|s�;�}��hm�g�L�/X��R�h�4쌞�m-�|��Z��ٯ-4��>���G��]ɋm�̗��>�yH��M)��d�6�`�k�3X��{>�(QάǶ�z}���Ϸ������c>O�r/�~��oޟ z�^�/��ԃ1�[��*6r�����ĝ�@ه�;�ӭ�t��|�9_����9�C�^F��;Q�u��Q�[��7��P�]\ȿ|���gN�C���6j^��!t�ε~꽤�����x"��S�`���'uo}��Q�7���t��.���ǨM�⠥��j>\�qg�Fr��]^��E�ya\{�j���\��w4T�x#��r*����+m>1Nx���⃃u�ɴ����p��x>�M�ɡ�Hgv�} /�i��xT��ڭ�H�=�����!���
�71ୠv_p[N�ƕ�XC�*��ť����Cuq�v�$�H��g���^>��<��p�|�|�����t��L���஧�tt���J�D�lߦ�����K�!̠����Ο��ȏ]{�dE5qݑ���ƭ��Cĥ�e����Iv]g�ԒQ��n=S9�p���y�U��i�xq���cr#ޯx����Fs�TB�F�e�U���?nj)>��g�qtW��>i~�>{����,��z�g�O�܏u�z��9M���`��1�r�e���`>�~+�ubK����du)���A|�vTOKw�9�'�{�,�ޘ����0k`Lm��l ,�GY�鑞�S�H�H`Xn�ql��ƣ����j��o;9�+��^�>��q���N�z�c2���,҂U>�'�n����X�1Z��ɾ����}��KS~�>|���^��gޝ��;��n=�\O_��dT9��|�a�De�O�gx���[w�Ѝ���G�g���E{�x��>�*��}^z=>V|r=3�%�F��v�&��:�"�Gn�5�y�L��#�.�@�f*siQ����o>�*��T�:�"�IS%����'����`���x�`���&6�1���6�1���������6��lm����l��m�cm��m�cm��m�cm�|m�cm���`���l�X�`�����6�鍶m��6�1��Lm�cm���`����m�o��m�o�m�cm���
�2����0">� ���9�>�>��*�+ZU�	%6Ҷʪ�QH$I ����h��!M��`�*F�E%*��UB��kf��E*�	��DDSke��ͦ���j�F�-�6��j�Fվ�9i1������}ismmmMm�c���j�ce���ci&MT��S�S���&�P�geV6Z���}��l7�v�5$[,��������k�&UU��[6ƥ�յ��������6j*kSV�kRi4�Z��aMkF�b��֛6ڶ���"����m2�F��   ���.>\��ӷ�T��˽����^���U�W���Sln��{y�{�7�n��j]U╷G�[լ�����*�ks�n�h����yֶ�ͺ����kk)�I�ձcPe#�  ��Ԉ�7���ם5[Q��szf�5=��ި�|�(��Οx  �F�Gw{�x�  ����QѠ(��G�=�    �6��  � �t�}� � �y��+,{��>��T[V���π ـ�}�1�h�6��%�^��g�UW;��=gC���h=��#�x���F����vԪ;�������ǜ��'\�t��R����bAkjԚcm�i�-�Mi�  mz��MN�ﵘ
]��{���Q��{��׵b�����Ӧ�bz�/=Jvʞ笵��f�֊�mn^�<���η�U�z��vn�����z�cm+�=�{fQ��&�lMT!�,�  �/��+���칯T���ͮ�K�{�P��M�Ǟ�o{8�v����M���y;ݵ�/6�۔��	����{��9������7l�pʹ�57�j�Ӗ���s�S�٬�Un�����a�i��   ^��o�sN�ޙpOI�Ηl���GS{z�7�^���:z���k:��{��Pz���m�׻���k�mwu��z�-^��j��yo7-�v����컕�]�QJ�;��۹�����4�u�U�4��n�]�>   #z����یjΏm�aһWM���z��q����l�;�{��m�ܞU��M,;׽̽�y��׎�����ڷ�K��v��^Yw�K��7Om�+���N����cǲ�b�m�V�l���u6dƖ�   '_}ٓ��v[��w�v���r=*�]�U�{���k��Hdҕw�Wv׻�w�v�v�z��=�m9���wm�Sݵー��Q�󞺳�o4V�<ͽ�u�4��Ooc�#k%-emU�R�F��\o�  ��}��=4w��z�[mݥR���^,ֳ�JǞ�k�k��ڼ<���v��ޫ�/5km��5��=��W=�������N���s�r��{�lsg������=�{,�ֽ�黎^�[��h��   w��>wv"+ޭK��E�n�o]�;ֱ���l�zK۷��n���޻�mt�5k-۷�	u=�wjTcʴ���[on�:�R����ڽu�˞Hk�ǻE�V������S�i3*��  ��$�E 2 S�15*E'��O��T=F E?"f*�M h2 $Ҕ�aTR@������W��/���fin��]�u����U��v8{����<��?k[η��	!I��Є��$�$ ����$�BB���IFI�����Ǳ��?��X)s�@b��YӍBË(��d���.�;i���,� 2�F���4�s#�b��b-�Bw���̌j�ڴ#��Z�C���!�̂����{��Q�J����t��W�ia?^U��$\�Yۓn�L^DV��z�� �8%6mo�b�����(1Y٨m��4�����:
meZZ�u��і3P��he];$��T�CZ����M�#q��Q�i労��NS ��iWj�X�i
b�>Ƿ��8����޽��p�R�No�2�
��a�Q6F�mReZZ��h�T#(Y'scҥ;�kqT
��X�
=��l�b�(��*?&jKV�R�\��"5�ǴG�}���86��A�g/R�D��Gմ09�� ^�}}-҅���ڷ�C�tJ��C�+1M�h��G��!a�5�<���5�,F��{���m���=T2m+�an�"��]iO-i��Ӽ�1T'1m�1,3kx�غ��M��dX�짦�����	N��)1��p`�X��H1{F�ST�r�,��W�`�:�H�:����WCz�t4R��X;fM%�GQ*bBM�f�.f���X��8u���T�a
[�4�ղ��N���Gen�@TԬ����T�4ޣy��]�X��F��3_�U:�!R[KB�ۋVj��X�ee�jBñ�6�D�d�q�d��x*V�ՅƖ�
"o%@q�Wi�4qR������t��8�U�F���RK%�t
�ٔ����(��+#�$LX�;J٫��"5Y���5 0V^%yӒD���N��Lm�fj9E���ae(�f<LY�,��ViԼ2K�fb�S�`��u�-�b
����H�b�l���6�t.���]B�$��8���ݝ�z�̄�fUᕅ�B$kVV�z������Yy�w"��R{&�����h�(,�݊�,��P�)�u�9+"!әcQ�1��̔t:f�P*ͫ7��������)s@[x����׵�����wn��u�4���`Mu.�� �`��Ovaac��[d̓b�Oiۦ>��0�֍�-��� �JTEm�]<7Z6Z�Y�`�$��ωט������; ��!nh4/M@+Q�d�h��P�J�L�kZkk��.��iJ�՚�S���á�\�)n^	�xN7W����Ґՙ>���ܧWw`Ԓ1�hYX��WB�aI�h\3$��:��5�Ӻ���4���I�k�_c��g�H���jR�`�^�����.\G*h%m1��J<���L�s�*�mҵiQ��ӦD�A�z˄Y�9X��1mh��Kz�&�*{w�dʚ�Џ�i%A��f��cYz�0�kp(�0e��s�v���2����b~���¦�`h�oi{�{K�X�S8�9y�]B1J������bϖ�����c%�X7*�Ct���7Q��XTb�9w(¥����#�S��Q�ڻ����3	:��Wh�@����H3pF�0±w����۹��ڼ���[��^�m�@0- ZPVp�nF�%�+�S!Mm;�����LB���-C�aq�f�B嫰(���J��I!��r��C�a�{��\N�Z[��Im �ɶa˲tm!���"r��������̗4��I�֡Q�4<�uf��QVZ ��KJ��٘�Y�@���c&���F5�C/KY7*�cJ�k+��ǹN�
2�`���3,24��a4���@r���EJ�F;�P��3Q@j"4���iVm=u/e��*aO wA%3*�3�0���!Y�"O-f�aۿ�Ad���=���W�M[Z[,hd	�u����em�ȢZ����8b�R[��%Ep�ڕx`��+]b)/���H�+7&쁅�F���dra��w�U�hf+Y��'o�0gִ���hj�������r����%�t�.��ka��B��ǅㆡD�J.������5�����5��������G7E�D�7rD���0���g&Qں�5����q�r�&���1���*B�� �4+ ɣ�ّ���^hTҭ�KBEp�۹h0
i$��*9��屌�9�0����5��&D�RAu� �o%Դ%�[��������d�oV)�Aw/�z�K�c�3@b��d��ӂ���Nӣo�0�Κ�B��ғ�Z5�!'
M�/[X�k@�M�	�����ZP��V�O[�YF���?"��Ѧ��YsS)������DI�u-����7$�u݄r��8�^�b�ҝ�/.�6ZѦ�T��^M�f�[JUr�E"�Vs�e����=@Ԧ��	j��]�c#�L�J� ��r�Ce��`7�,���Y��Y�L��^��M�LA�6��tn�f���,�vPBkv��v��&.�)��g"�+Tr١����HL:/K�Y�X嬭�Q�H�^^%$hi2n��k(;&� �ld@<�Jx��um̔,�꽎M�4�%jd5%�j �f1�8K6r�V��8��<��q�"�m�E�cnV!�t�)1ˠ� l�5�6�+�̥�Bك���֔��h�GJu�%��`^i3qm誰"�Q!�[=3/�)���浓���
�<�O��>+�h���)�^V(�% ���	M���e�Y�QT����1�E�V�1Y����341�鑔�Z�!7�U���JJx��7Tr@�e��i&�{ʸb��f�os�h7W��@����Q�F����B�컍[(��Z�.�Y�m���fK�y�
���+f�IPv���U����?�)V�ii޺Ya<��^	�)Y'TM��
[�;`�]�à�m3A���qD�96��Q��5uc���Ùp+�8�Bm����l���DBE(v wv���L�����$���f-PJݺwI��8:e�y5��e�����)}�aI:���&�Y�M�������àڽ��L��əWm��w@�L��ڽ�$���p�/hĆ	n�fM��t�p��3���YƱ��'v�����7�K�`ҙ�'�2�(d(EЙ X��
�l�5�EZ���t�5VXH8C���0�n��`s&�0�
iJMʙE=Bdoo����J�Y�T,�pYn�<��f**�,@����)l`KuR��\@ �Ҕc���@(�
6�M���۟*���I�̱C㢃��F�A�&,������@�j�1�%ZWX�*ӕ0$�.�O"p�ZĲ`u&�r��Q�P�9�|�ܩx#l�.S�aW����j��s-Iq��.J�����I���mP�j	sZ�Y�Ŗ@e:��V�q˦U�Ц˫�f��c��ݵj�� j��m���Ⱦ�M�Z�v���U��M؞�*��lX��eSxj^b�(�C�2���xF�ijpf�D���-�t����Z�2���a:���N=
���@J;����J'�n.Y���^�s[�ǲ��Zv
OR�0�"aJ�J"�=����gIr�k#�D��J�ݬb�Bu�˭��v[6s<��2��;G(���khbz��w3O�cB���U���,*�4xb�N�Ŵv�ɐ�
�-�uk�Z�<���
`źa��J��v�aI@�	E���\̼a�ť)�O�L�dOH� p�f�ƒ5��J8.�G��L�WsJ��Dͨ����)����`���n��fJ2jT��u���4i���`V��r�j-DÐY�e���CNl��un!󚠫+��#X�ƫ�Ph�	���z2�b��Ø��m���l�ܔ8�׭T�f���1G�)+���S]M޷�Z����@TIڪIH}�T7!TM�6�v�T�%�����R���`�C��p�,�:�zیXr�W�K���e�ͬyt�ii��d��J:9Na+
�)(v���6PN+]�NXA���2��y5J2)��4I�� �Pm�Xa�E�pEKkr´2�!,ժ�D���A3F�k�xS�N�`otҊ�����()Ф�"c��s0VSI��c�ԩ��û�7]�0^���2��PZJm��ᦣu��$6�n�v�V��k0�h,Ȇ�O��a��2,65���Cl�Z��n:�VݝZ�Ui���]�3���;��GF޶�5����J�̠,�4@9���e[E�"��M9���D�Q�ғ 2{R0�p�cW��8E�2�2�G�6ź�3�,4��Q�;M�r���n�a��Z���լ��QI���,�4��aVZ��m��2:nMRYV'z�%Z{�SC*�^�%�*1'�.�[��ovV�w%J �ik�3���2���,l��అD�٩ʹ�2I�ϥ�� ���mI�s]�Xl�yH�j?��dǲSЉWHk@�,�^�3w0�W�n���8�#Gd���`�����Y�0ͺV�%k�z¬���1�@�鰼d嬥�`4V^3y�ʗB�ɶ�eH�2�kC�"Xkq�n�2��&��b�Cx8�y���[0���@*"4iKfJ�i05��;B�,3/4��,VT��d��9�M� �N���caݑ�lh*�Ǯ����E�X���RI�0���ɻxH���A5��6�[�n�#�7�c@ݦ�̦�.�6���Q�(���xA�r�[��+*X�S��T��-WZ�I�x�{I����,���I +��fe�A!�W�A�F�{V����v�"��g^&�8�0������X�c����"f
&���j�_l����ө��U�Hf��`K�p2�SFm(q�O`�a��Y("���[$P�o6�0��
�f=��,�)`v���kiW@^���=�˭wy�%a��)�^�YL�Ҷ�ڷ$l�,i���l�I�&�2!��e8��D�9�JDY�P:�q�,�U�2!Jm;ӓ0#�,e#�(�х������OA�ʼ��Θ�B&���Z� ��q���2��	$�8
Zq�����Ǎ*G�f�7@Fa���萞�6��ō�ln�Tf��&�a[�!��+����,/bZ���Ű�y��ئ7��%޻ܲ���J�6b�����N��{b�lh���lf˼l�I�&�ݥ�7C����Fڱu��I47Z.��s	1��f�܂�\��+є�O]K� ɩyb�Z(`�2�QMD6�%��V�ܺ�3PR1'�Sc(fW[@��ؼ�z�5$bd���e^	�F��L9/1�R�Hw_ŁMn��9�@[7lYM��M�tuЖь+�Y�o2���Ub�JB��b?A����M�i8tT3�X�w���V��e�k�i��.��LbJ�wJ�AV'�����L�E�'7%64M�.b��3wf���G�Lʋ�Rqԍ�i鬹GV�R��t��BPT`�I)k6�1[$Ut��{Y�@?lEc{�}�TQ	�ʼ�V���f5P͠�h=� Jo]�4eY�Rʵl���4��^F6�}��r���dJM��7񫴅Mg)Zٹ���(�j;7`9��nV���S���t��5$��Ƀ�Ҹ�]ɚ�M�r���d�C:(�]=8��U�vP��2���	��o5fj&%,3��r��	B��gؙw�ˬ�o�^�y�Z��jc.��u����u#�&��k��H���-
�G�J)݊�e�Utp p�-P`p�T��B��\p�dQ6����xS:B�͒hb�F`J�啑M*F��X��b����x���ȩ`X�-��E{��͔p�H��J�n�Ƭ��u���7SyT(g�V�&��O�V%)ܗI4Z�W�"u��よ���BЧ�e
�
����v1 �Fa��Se��$M��2�
�V��������w/PLH���̈S�/sத�ã�f���uw�b7����µW��ܚLŘ3����'JBm@仐���CV7A�p��Z��(�n�XX
}��,�]�лՠ����u`8����r^������V�Ĳk�0�ai�駄�[�Z&�j[�D�m��k+�
�VݙV��.U�l�Z��ZW�m��5�&8R��̌�B����ܻx��
LvUf�����ژ�$�滲�*��OKY�r�F��`�uef�*+��Z�|���w6S�5m-M��J��9�ph��GQ���w��qnXv�ی`�2mjs.�'�Z��1�2ߕ�ff$�R���1I�R1�-��lؕu�����\�4����`l�!���\����w�V,o[��M ̣���2�K��3w*�Պ�r�����͍�#t�ܖ��znd�{.Clb��F��K7��+��
;���i�y-�u7��8���[0:n����W,��f�y���h*�I��D�,����ڹyf��KcV�Ղ�����G&"N֙�\)]�a\�M���5��e2֡�ٴw���%l�q�`��6��f&bT��Eqn+f�-<#bɨB��Z���,�	]0Pa[�]�1
���36��JӚkVꢆ<��Yv]^�T��?iW���r
�LJ�r�m���2m��M�E�5���U�yqÈX�y�:�5;X�(ZѼ[������-�����0ۇmj��Hj��N��AA�*��8�K�8�5�TH;�=��V,�uz��Of`6��(�a���1$�rњ��D�M�RlH]�=M֫����3�T��Y��q;��iCt�������^�&8%f<��]h!S�	m��a�V]�ݲH���+�i����i9��-)k�~�K�o��4���՝����ж͘+
��S5����辵]Le�
�,f��L��uM�/�]�>��.��ipL)u���WB����FpZv�\H/��_��uՑS��u�n`U/�%��&Q�mD��nj'�j���h�y�M���|�J�:�.�I#�b�}\�h�s����q�"������I�Z��ӄPigu�6;�z9QLͬ��N<!B҈T���ۺ.*�e�H���mgpd	�r�Wd4�C�f��YY�����pJ�c4���,/��QgAv�Vͣ+���[���Cw��V�a�Ma�:���i}�v��:�+�Ror	���6�(�����P[.�e7��t��]"�۝;LLH�s��Uդ�O
��+p�G�ΌN�������e:�Β*]�XC=D^��׷�ią�os� wPr��A�oY�f��@Er����W��7m�zw�f!�DPz�f�'d��ޗV1�;G����gT&�-I��J��y��u��T��+t:�M9�[��YN�9�y�,`��>g�Q�V���A�t��ȇ��'v1�P�`2h���1I�Qԅ�[X/l�:�쒴���cd��Ot���#�F��/%�?��;w]:)4��es��ĐmL]��JKU7z�Sjue奐M���-�i�Ђ�������F��O#���<���"����.�wh��Ќ���ã�)W*u���gtk��m��fa+Z̵oG�r��A���C�w\�;&�Ě�I��t�Fu�jT���"��&�m��RX�F��.���J�Vf�z���H��z��2��nVq�Q+���nC��9Ѫl�PFf�0�6�4��v�λB�>ZuwJ~	�	��IɽJ>��{��h��X7	T�Jt��N'f�c3^��ev���ؖ�S�!���q�r���"��\ܘ�>�lZ�V���:��q��X;�#{~�QVV�Cqǥ�ȃ�sW����'`q+�ԅ�f��t샓�:��R�-��c,�R��Wh�A�k%`���.@-֞$VbԈo5�q	] ta�u��%Ո+%;̠_mڍ��KS[yS,9����3���ܧ�9 ��E����oh�ц��D.���Y��]�#�*K�	:Z��B��E�ݺ�
�$:�����<7!���eN	��S�lkt�P�m�*��,�x�j҃�Bb��eP�$�6�e���l�.�-�Sj1o.]�G^.2�������(wh���v���{\qX�s�tM8���Me��iǴ38C�����ҧڬΖ�"R|7$V�_(PɃl2��M8��;�u�e�+i�r�����Q�nn��}��>��7������"4p*��Լ��qQ��`�\��fAȲg�C��&�*��d���դ�ǯnL��]c ��S�!8���Aįd�;Q����!�n�����w|� �.�9O1��MXy0M9��]�]������2�nr�����]3-t���I%J;Fd|l��Lt{�,=4��c��J;�)��;��&p&��1x�О�����b�|��ɽ�kT�[��R{kE��4&d���g�t皸����D��J�M%]Z�V���:]u����I���6�ڑ�7�]vg���%�W�8�	3:loo�-�Ȱ�*�*��Nj�dé���u��,�P�ad�=΢����:˩�D�EC�m�WҰ��#�Y �E�ˤD��d���g-^�h����T8�T�S��H�ۻ�a���z'��Eqcf ��2���n�j����Pԏ}�U*�<�f���~iP��� �W[�d�.5�fvcx��I��e�	��q	���_:Ŝ��`��r��pH�t8^�9�5��ejЕ^&�:�*v�Ŋ � �+q��`�v��Ӳ_	����oֻy�"b��f���\�tGZ�!���Z�����k�D�cb��9�S���y�(
����RWK�t{�9����*����4����-n�&fήJ�3�V&�oq��(���9P��H[n�`Sq��mBP�rb�0�ox�Ws��:F���]�ɛ6-/�{mb'J��:<���G�U�Z"RN�eY\��W�%�ب���a�f�Ug �oe�ҟO�̜Է�Z��YRd1���"r���8%*�yy8�9�j�{Ma�,,$���h솻��1f6���xZ\�)���t'��h�����A�6Y�[+�l�������[ۑj���Ӫ�*�u�im`���"\��X{P��(�q: V�Egd��E>ѩ��Fz�j�B�srၭt����˟9k@�1G���|�u��������0'R]I!-�άG����3%��V1svN8;Q"H)����PT���|�����/ ���8r�F�Gg��"�lpIc�/Gd��K�i�Q���:�SMsƂrnAC��Z���i-��zY�e.ې#��ǃ��2 {v�'����]��-��,u;��H����۽�mI�z������a]l���pø�x�I2��ߵ���4���Uؾ�Q��r��NԄ���a7rM�Y��mv����R؁5z*�[ޣ�Y�fe(KW���;Mحl8�Ryd�{s�&n*E���]]ܨ�5��g3�ms��'�bJ��|��6�fml��[�8�|\<�ɐ
Ji�:�ȫ�;���i��s�ͮ��P0b*1����4{U�, ¶�Zr��uO�I^�Elr����&����K2j��sukb��
��FH��ݧ�E	>��-,F��S��;n��ތ\V�v���:Y�w0ăI��1��̰6�1;�^͕:�U��&�ôڃK[���כֿմ]�l>�؅�,�/� �Z��0��_#�/	���4��tݢU^ꥳ@�2����F[ŝ��(��m%���o�[2!��������s�\�a�v(�P�f!�F�[�;�f\H7$�����N��|.��l l8p+8Gk=b�]i)݁��k~sk��ʲ�Y�Z�D��H���\.=�!�Qs�ۚ�.����$���(�G3���5�Ć�ʸ#��1�U�]�����Ώ��q�Yv�i]������Jm2�\U-��C��e��3��r��f0\x�� q��W�E�7�j�A�aH��R�*���2��j��>]�%JV�-׎��eE����C� S<�;��:���aݥ˹b�ٓ~J�v���z�,���1�Em)B�=�ً���L��yC�)Fpo�ϥ�����]܂u���Dbam�K+f��m�wi���1ڔ9�Q��p�
ub��Y��]c��ڵnuڔ�غ�*Xm{��,�U��<�mG���i�$��2]���S2t�q��XU�}�h/qC��:��6������!��skJlZ�����EB�wt*'&��tV>r=%�Fi9ɭ
�82�vS�8�a�͘��;{L�zX��ލ[uf�T#�+xd"ӳxk�]j���W���}�"}W�ݎf��D�)m%
wW.�0��d\k*�ZЇD��-ԝ�9n���{ώ�4�x��z�/xL�08��H� 
GљK*>��}������KXY���c�:E�4����XT﷗w9������v���R(��7Aq[n�T�)f�IMw���u�m���4���ݥ�rhq�Y2@m�\�+�8Vi��le�2vK��/��Q���؛[[mTǁe��%�\�y]�p��+Z�b>�nLv�5Q�ͧ��l��7 >AJG��mvuЩ;Ed�7�PVo{S��U�+"rZ�jJ�f�S޲������0�\�6����r�ӛ��N;l9�?O^D�'����^�Q��n��楲n�ܺgP�r���O�R7�o=�meYzr�#��ۚ�rΖ��aμ��k��C�ۆj��V�+��C�u�^�}�m)���;ps�6k�m� z���NyYb*���`hdk&w*��Z����b��A�y�z\�M�����&�p�΅���Ȟ�T���qmo¦���ν�]��h��9w
�dI�h��v�h�X0aAe�K�1n�J�ٱ���ξT��r͉e��/�ӱkw)Ƌe���E�f��:���JM�l����㾐h� ya�{rs�U�'�E��F	��k��(�޺�a�Nl;��p����یTέz�͜�lhۗ�rt�g*'����u��_X�ܷb���5��S�:�ퟞ]�j�^gtu�6$�S�-�/~T����c��yC��c����-��T��,Z�Gd��_����7A(�_�-�ia+�Pӭt�ɀ݉E��ݎ�[�/�=����/^(j]�*:
P�֞�����{�;�Sb�0U���l�z�f�kp����I�k;u�m^ ��Sy�Ŵ#���]�ON�ni:��^�Ө�ܩ/��a��z�#��7��,�����6��x�(ws<�wӯ�ږ��ڌlyL<9��Ҩ)pCz��̴`SZ����2U˓,e�Wn[q��|:.�����v����4t����48��
�T���:k{�U��C�Ś�M�j��ڽM2��.aT�=��m�$��i��_T�&7Q��2��U��ʡn����a�d/���gK�(=�K��,����D{ �=�ԇ�g�E�qD`�����6��ܔ�C��ܵ�u;�B�ܬc9�1b�}�l�C��㴸�w[�yp���*��b���R�F.ٻ컒:Ӂlt�o$B2hæ�b�qH���d��:��ˁ�u���s�u:6�u�s����������#��XU���e�o*,K	
u2d{8�f���0t p֣�"�.��EMaT��{k������P)ҺU�ppve��]ڤH����r�L��2>��lwY�h�p��+������Ǖ�WCVZi���R�v�����OnlÑf·�*�w9���Y�y��}+��M ��K���r�evܹ]���g9�K�Rm���J���94���7���F���0]N}Յ���ME��m� G��Q�o�`���!�ނ\�SN��P���o*�D�H��v@�,��Qn�4;��[��@]uM}�wp�����ا-�Zc�/sR����(=��s�+�Cٍm�bS�u��N� ��T9��0�+h��ùX�5V��r�=A��J�=��8����+a<��Z ̬/���n�QF�\@�n|��i����݇�Y?�j������h56�v�&;E���,zxf��[��,�Ww�r��;\�(�p��C��	Nb蓻�V	œ��]]m䙵j�sv��/r]N����`�o��b8]@fi���BEZ�4=�ne^54��%ow�;'�u�S&݉�d�o�)q̼Xxb�z�8�r#���mK�@�������`��6�n�(7�:�Q���T.ʩ(����.�߄P���>�X�!�1u��緤oPV1a�^�����8��a�8Q�W�_p�Hj�
0��30��o;;�e��6��Z��÷�z����RR�Xʸ;tȻ�� �`��Q��c���yHJ&�����u}H,��%ٍ�9���~��7w�k��ĵ�a���Q+�%��V�nIy��7[��%�:^��b�Mu,�ܬ���P�a�1a��O��w1t쩸c��9\�J�2�8�h���<�x����+x�K�h֋��$T��h�]�z1$v�nP0���-"ީɝ��7LG�y7�%L�p�N��a�"�����/^�Ov��3v3i:�u�<С/)r�9�lJ��Ycd��S7�u҃y�25D���b�חq��\ð!]7����r>��A��p�൦l�l
"�ʗBM"�H�h�[0N�Z�<7&p��k�i�����jQdu:͢��\wl��xH"���������Qb�2v
�$�`��G{���um��̼�%��4�M��33A��i ������l��T�4��'����V>'ln5x�ن뢢�p.���^���S�k�tK��Ssc�-�$��J1���KǺ.4�L�,H�lZޔÏP�E|�wh�ot���79�����!hn&���Α�t�6[m�1���{1E�t�h]�qք������r�~C�A�m06���H�s]�\����rG����/��=R�L��MJ7��}�I��m?���Yj�gDz���g���Go�k��]~�!��19��j��2S�ٮ�pMCWm��v��sC��Iʴm��nn����7};�7�'��Y��[�W�դ�k#�T8����E�[�p
-j�e�<�(5[�6]�&
ɤkB����C��o����j�e&��Qޫ��:wm�iA��/S���l��"Y����㙽pV9>���s9�v��]���]���乵O���*���&DMk�r2%���<Tn��̤ask��� ���I�[��Cƣ[.d��!.���F�D#DE�s&s7z	��T�G��rC�Ξѻ�5��,���o7܀�1��Q��:4��P����r�;I�[�t%YzN� �锤�o�R�ie�bj뮺�K�h����t��v�L�;n�	W��ru-�枭�v� *���S��w`ri�;�9h�\"�֜��+y�\0�9<z\Yx�i�7P��$Tb|�\��g�9������ƚ1�bԭ�w;kkh�y
��i:ד�X.����2�#���]�fp� ��8c��r)��7ٽ�3'G�����ޮ|K ,	&��y�0���NWMm��+�͜�y��n?s\�g���7���! �����W�_}�%~�?h`g��鬬������g.-��F$��[�+Pcy�&��O,��e4	�Opq�,��x��0k���)�"�Օ���Ue�u�˲�F�}zfǖ�Q�З5_�#2u<�����X%=�\Sb���b�Oz��z���v��/1,"�j4�wIm�.ʬ�i10����ίldٳ�G�f���mL��6�]+��k0��*-Lu*�>2�L��5�63�d�T��O�YW�6۱f�:��Ѩ���±W,�M�b�x׃�h�"��{gm�y�6��-:Vl"'r��Yv���$�ݣWM[�~�h��_Z��`u<�ޞ�;��ϭl�;��Xس�a���9��C!�4PDc}Qi�Z��QR����ՠ�&�c�붝�te��Ί��\��E\��َgXm�ڵ6��b�@Өz�h=O9�T̬��2�i���b� ���k˺����<�G��͛>�pN\��|2��o����H�d7��#D;�<�ɕ��`�+c�ald>@���u���UԪċ[.��ꦵ9�{�T@�2����.U�d�/J;эT�Ӄ�^]��+uĭ�t��E�6vu�ǜ�݆�A� �TK ���eؘ�E��Zs�U��Z9��9rn�w�O	0�Se�3/AN%�vEԄS@Sh���3�5$�r��.��I�i��.��;FcWR��ZɂP�"O�t�T�W7��C��� F£5��QK6���[ @��-������=4�7sa�V0(ox���v���m��-����b��rpr�f�+7��2S�$�&m+�ɵ7�/��#r�cǋi��I�S�m�;�������e��@i���j�K[%�&�[��,�ՙ���n������A&�rF$�;.lY�v��d�Q
ԏ��Lhd�,�ӕ$f;GBX��݇�����XU[�[�nU���^� �ھp�P���\VD9\�J��/�q���E�����[5̅��ҷ�ȓџR�+]���
��tA�O�K<�R��,���(;6�,&ˊ�d�wlu��WCJ홸�PS�t���*��D���j�6�_I�X�� N���mE��֒��ٽѳO>��\8k�Ȳ���(� ��<a�B�H�0���c�Mi2`��c�I�+�T�y��VjM��ެM�bp�nr�ۍWe�f�c�e�}�����(N`.n��t�3'\�#��z����r�Za
籨�h�hgJvp�z,؝2�X��ʛOnD��u]D��+4�$�5>8)4k~����s2����rՊ���+�>��`>�L� v+l���j�\�x�:T,��K���[A�L�ul�#���!�Vf{�㥌L�8
Ω/"�e.؊�Rξ�M���JwJ�QlN�yY�M�K'�r,e�N�;�|Ѷ�
������]A�+�ʦ�#��&�,f��G;ݮ�\B^(���wL�7r�+�8rol���֨nZ��:.�c�8��I`U�jU�֙d��H�" ^kؔ��������X�ۓ:��pX����03��]nczW��.o
sU�[8)MK����f2��r�u�2&waP�������c��a��!�Iz�9��,�xW)+7�d˗��7K8
��->Y�ԭP��S;�����F6��2�$0�1��Rh�� �Pss�[�L?9���m�X�����P�P�Í���q��#���m��jR���/�1��-���:�$�`Ȟ�L5�x�B��V"��r�-�)�R��z�b�+N��F�ZR�cJ��X�gY����mZ�EX�+z��)�P�`߆�e�vm^9T7s�����uo,r�[��<� ݻB��+������ls{/�[;h�P�I�`7G�M�7K���)*b;�����%v�wR�WAa�a�ɦ\yY�Lצ�δ�����ߗю�Z6�v#���f�#�Բ�#�Wӕ�SclԴU�Fц��8#���|ؖ�9��,u���yWώ�Bd}���37�h�H^}�s��5S�--�Z�!���r҆Y��_@�rvR�Q,����[H�F��-�T#�*��N�PojS2;�z�r(7��Λ2QPf ���fM���	]�����_Q�h�C:6n6�$ ZT�ujź�v�kOR=�Z��<���,Y�z�`�Z����>���l�'u�3m�cr�'��\��ηVE[2*{�����K;[�k϶��n �֩�HK�8�d0[r\��G�e��!!v+{�a	�8�0�5�z�"�Lyj�
��m.k"�Ut��t��x����8:U�`��@���}���ug\L�b����˥9�:�w��-�p��]D.�՚��l��r�4��=!Ħ�l���O�Y[�ӡ\�gma��^mj����EwB�B4p=�3- ʜ�'s-X��{]��}Vw�a7I��2�M��T�LǪ��@�))����e��eM�	֤��sZ�m����6�^ؐ�n`��CMf�/�q�t6���\�[���f�M*:E�SNu�G5�s�>,�l hK�j⺶M�%X���|�-T��#��#���Κ�#��voL������و���ES{��~6��4mF[�.�O���ɣ)��s�kk#��$��'ΐ�Y�v�<��0d�4���F0���m>S��xE!6�t�&��.���]L7 ������[�����!���%�>4�C����G��y"���8�����H�+�����l�]��6�Af�t���֜4'e�
���/f�\:5jmY4�^����$)���+�ٓ]�22��[-.ܢu�b�f��{��6�XNVS1�Q��*]d��>1����<!jK)�lj5�BݱP�\ۊ.���1�ܹ��=��� ��Zva����m��˼�/c�t95�5�zN+��9�����xG Y�� 7S��}�M&7V[MĲj�Y��;e�|�����	�V6'h#��ޝ��Nq�w�l0���
(����^��6��bw5�F�=u\���˝�H�[n���Бb��f��� ۖ�E��`dQ���l�!�=	%rX֦�5��ձ
F�A3�ӓ��x	�5��s�̖4�C�La�+�҈�w;��߈�A�E����k$v�6Pj'�ެG�8
N��@G�*�X����˧
��9�^�µ��V����d�5|ߛ3��	A�N�1�ҥ�բ�-N+��s9�]�K���Rm[k��F�,�SӁiZ
��r��+�{QL�ᄬ�V�j <ܠ�1*��om1���יu-U��>�k1F$�{E���
���2��>��냫�9bY�Ʉx�Ș��Y�W�n��FP}@�Sr���P����>��:����a&k�!%P�G�ea�j�:��t�ڷ��V4Z�u+ӡLp 3�A�Z ���Y�����P���{�q]EQQs/J�.�%�F��Mӝc�˫����}"��k[q}g��NBMe�/�~v�j,X�}FXi:�ɹ\3c�R�;,Ż/HϞ��[*2��FX�ΗF�k7ڒ���A\#&�їϴ�c��7���N�%�4�p���Rx������)��F��&nul<�B*���Ǌ,.�fT'1N�T�fi���ҫ4cf����1[��@�0aUخ��}:;k2�Y
-;��ݺ��n����0�: �oy8�C���rK+Uޛ�)c/4ݜ�̾b-����0Һ0n�u����E�3�~�7-7ű�2nk�C0v��5*�P`AR[��EW��O}(e�\7�]��"��� �-q3k��F�����lq\���y̥�0û�Z�Sf۾fP4���U�+N��W�G4t�R��ĦQ5Р��kX�?Ǘb1�XenQ�t�B�&�|��mۖn�)i�)����ս�E��;<��C����tH՝�㵩��������l�څu=�0��K���s����&)�
:�E��o2+7bG�m����\,�j��Աs�m�a�]��k㹷��
���*=��"hd���P�e�L�U�I�@]��,F��Ҁ�׹&mGr��@:W�rW^pMo�9�悫��i^��`V(�:���͚˟;s/T9����h�<�E���$w�lr��S�2W	�TZ:�i�7�PW8�I�1z�^`Z��&�׭��~v[�
��R��q��B�Y���5��8�eoa ���9t1��uITx��K�bTo�c�K��'V�S��e�Z}|���u�� s�Uf�Kt�`aTnfI�z�#�Xb�$���ťt�	�IO#ť�r=�2�m���v�jL|���9���
��/6��{toC��H��*n��DQ،�9\��#��k@�Pq�]N��c���v�Kl��@L��I�1�L�`\I��h�)��'��۩�p��*z��xq��ʌm�C�aQw lO���Ĥ��왈�Ph$r��@P<��)	��#@�9RJ�P b�u4���ő ���2C�i,�*�|��3���>�ݞ+F�$�T��h�ՕaGw�Ыe����;K���[��n�=n�R�K�ҸNw�Q^�JE:�<7��j|'��%0_�u��R��ٯ��PƫC:�*;.L�i[�F�Vn�̳}�h�o��PY�A���(�T
�s��o�M�&c�W=\MӱJ��;)��#����H��+����xE��c��2�U)«XM�Co2�����u��Y��%�+�, zk|�Nۖ�}���i=���|���Td��2gۊ1��4�4ɉ
q�o=�8F,Q�'�@�JzX"��81�3͑�&�B�����E2q���zRv���».�$�J�h��o��,N�;�N�hn����U���ڲ�,��%�;��,�̛w��b�t�[D���
�j����%�n�[���U��X�/��*N�-�5]�n���й�]���O�SnV��4(mit,�.d�t!�E�:;�9����fdi*éIE�t��6���Rį��D��]���P����U͹4;ރ�����]��fbL2�SK֪�(����M�\��e3�2��-n�|���c�����;��Wl�����x�l\u��B𩵒�V�c5��.<�ϐ\�Q}g\�8( ˜���]� ]��E0�ff0w�����>�Rʷh�(Z*X�3#��ͣ�q�:6iՒ�,�z�R�w>�7R�z�-Gaé����Y��2��M*����
�U+�����Zپ�����Ԇ�q� n��b��$����L|v;ɋ�ӕ�,�B�&�3V-j��O�\x�%h���&��[h� 0�s��]�>6����������v�P���ӄ!s�n
ן7��D[�[w��ṳ́�b��&�
�8.��`�FQ����=��y]$�W+�5��ލ��
폆aGU���2Bʺ��nf��&wq�\Oz޺���]r9�(�����6��yV.�w1[CW
֦`m���xጒQl��A�F��4�m��:����k��b�e�dڍ�ӹ�*����+�s��v���nS��R��膌�f�ib�v�ذ,�M��;q����]�K���̨FМ�Շ];J\��4=��L�Am��.�h5&���Yx�#;]XD��n9�,H7N���vq�E��hBl\,����0��a���H���5:[�¤ն*���'etH3��*]q�].֢�p��%iKX&VS/������;��AgnϬ�O�:� �����4@��EGO4�P)_F�2��sv�#ա`�3����W(a�+NN̨=�q-�dhΔ���w�tnģI�l�ZYZo�XHoN����[�{/mJ'�ze��X�fgP�7|��Y
p�m
����+r��X�73��8���I����e�!�oÇZ�;��g���k ��Z1��ԦRՒ�7�d����ԛcf.�1}��-����O[2�b�c�I �3w9
��C�G�G+�����ic��t��-���H�����Wet���^K�A�2+���&*�w��2:}uyk��@�%����ݏ�D�L��y=�RU��S�u��T�[�WLR�h��^g^d��[t�������TH�B�T�|{q��ټ�Y�,*�d�H�S�����4��묄&X79�غz>�Ba�wHU�A�7�:�JxF��RDyS��PxE��T0�DVlz��;C{v]�rp�NJ*�Vq�[o\�0��A��K�{����w;mk�Nʘ7��Og`�����-��{�7%J�9����S��3˲W����lS���#I�P��\b�i�&3�����(0ivh�ڧ��Ɲ�����<fo�2��mAzi�H��Y�h={i���>��Cc����Ub�78�df�
����%�h�j��k6Ҽ�Q�kD���)�w�4b�u�����T��c�B+[��Mvoq�#v����h�a-�Tka���Wb����Ү�X>�s*=�z&R���筟���Qr��j�44c��Z�t�kn�3;F����c� �o	��U�	v5v�g�pvB��Xk Ietfp��gT�-](X�Z��֬B�0���Y\oO4�}8����0'wF
��Y��u���CԍE���j�E��ي7�u��yݠ�{k6'+Uw��5X����I���*cҳdy��g[Ŵi���;�`}$�)�Df��}t��bD���6A[a@��I|�p�H�[���2�m�m�R��t�4&�4��X��;;�T$�	'�S#����7�uy�y���h���mt�J9�H򹓓�Vv�h�).",�ŕ|$\&i�e�9*9f	�]�N�PV�7�ڝ�[��n������ݷDk��}aCVf= ��ن	����<��ԍ]9_m +Ah�,
�Y)m 5����q��3J� ���|��`���"��x�=���B�rťua���T�X�:.�u�,h��E����
����3���3P�#/v�����)p�������7T����-�ʗY�F/fκXr"�X0�����U����gxw-�m`�X)����N� �l����v�4�R��pWsv����c�?�Zn�wfr���z��G� �/��WJ>x#8\!<�k�ͭ�����Q�\�U�O$�"f�Lj���F�y��ɳ!^O�(+t�tN�`kX��a�3L�khf*�	.fW爉�Q^w<�I�b�`\���N���R7�t�g��ա�j����L=C:��{_ x#�.�`[(���P3h'���X�D\���w�R�ma���v�fA�\T���L�Onh�f�F���������\Yh�x\c�9�&`��$9'�`����[$�m˺bq�;bY�:v�H��Ʋ��a/�]�ە�1�9o^�S$u㨭��k�^p�o,;��71Yh�Kw'�4
�M�M*��ܹ}ϊ.�߿F?P����"�
""2"�*��Z*1�Jb����*[(֩J�ժ
�A�Tl(�(����Z��ŌEPXĖ��-h+ ��P
"1e��
1TX�[eb�����*"�R��(���R�*(��`"Z�Q`�iX�(��ʈֶ�0EV�ʊ��-���
��PPAX�cmF#Z��JT�UX�#Z�E*�*Ѣ��h��+Z� ���(�����iiQm�YR�F6�[DDQ"1EQe�m��+Kh�T��[m-1TUAPQ��*)X� �V�,DEX*#m����,EEE�A[lF)Z("���+X�D���AV��"[b��(�6ت5�5(�b,QF)mZQ����V�*֊*2*��F���UX�T��,�"+h�QR�X1b�H�DX��TQ���"[H�

#Ѣ�b�J��*TU)iUUF
+���,P_}�R�A�=e��N��p����-\����J�
:�X�m"���]�(�y+s�)>�\�)���qW�,�ؐ�Êۥ���C酛�]1̡uҕn�hL�@8m�\1�;��
���uĐ�WDzWX�P�_k�*��ԩgEA2���&���Og�7d:�ֽ�S������ht����Շ�����R� pd�*�#� �b��Hyz�i��o�H=���W�O����՟�#�9d=�v�f}�0Y�R��S���w��.�$���~Ĝc����&��K>�X�n@��pf��o�2���N��ڱ�,A�z���e���+�5C�;"~�Vxw��"mv�j��;[p2�>�:3a��9����#�y�o���u�J�f���
�/�V�Y{�f�]N��+sj�b4���@���y�c�����^�ju�ׇb�L%Cs�:#=���#�zpi�T&���.�F��6	Nݴ5�p������RT�e{L���u�W���#'[��N^��m F;"����Q��5�s�T���#,�!�	PϯDPVp�L��Pu��^��yz�]�Y�UL
G��]ch�������`��k�H�C�Ȣ(��[�N7tgq��ŕ#Ν]6T�5]x�f��P��m��y0`�N���r��Z��/_6!��dS�W��MJm��N��{]�K80d�wZ�]���5�d�m4�LipK]v��i�#�-�OY�B����a�a(=�8�5)}Nu��8�w�7=��c�}���J����3@�<�� (�Hs�꘮�rɺ8�\�>Y��^Φ���3�Y����g'U�C���GMq4ǅ��CT�Y���ę��F뗟�.�"�_-��C\.��{G����Õ&`�w �[:�̸���'M!�7�ʈg�Y.��l������ŃR�,����*��4
�S(P�v�b�O�}�Pr���r&Y�A���Y��b,��2�Ù��3s��`�D˃f��cA�ɳ���i2���
�%�ﬦVx$w��:����/!�B��,���ztڗ��v��Ʃ���v�ѱ�:�!U����i(X��P��0Y9V�9�.A�γ��U&P��-�}=�1�x����W��`EA����iI�&�5�
�=�=�W��m�5gM,{��VJ�\$A�@w����/��J�Fϥj���N�`��1�5�����|�����y��[离�? ���g���U�8�s���.f���wɩ(ɽ)Rz+��M�>lm�3(�e�<"����Z+x��9]�Gɇ��J��6��c��l)F���ШXܭ��5�AZ������JO5J�yj���o!��K<�ߕ։�\�9Z� +>s���KVT�v�ҡ[�Q�{l�gu#���v^��{P��o޴_i��P񫞽��6�RV���:�w��q'�q�i�'��O����ڇ���eq��Cݔ��հ��n'S-��k��zDoŕد���'�����Kս�!=aXuz>K�K�	sԩ|��uKl��ا�Oe�n]�lԥ�໏=�[SH���+C�JR���/��Ih�����{K��<���]�)ћq�����4��g��"-��es5l�&��'I����~�h2d���TqW��D��~��$J�]M>�f�Ӽ	cx�`j��V:���]�!�������DF��]g�����2���|�(zu����x�{�
}쩷��:�{:v[,g��/7Z��n�
�
������Ҟ�e�n� �R��6�s���K�qzgHrL�����Mw�w�;� 	T)ȋ3x�����w&~�KY�o:~�[�nb[�� S����i�;j���h��ܪ��wH��+u�"ԑI�6^,���ŻM�_t��u�l�<�aԆv��H��:&pu�������ҝEY|έ�%����Sw&�S���cx�W,��N�g]p�M;��Ӑ��[%rt�vȵ�+�+Y�]��	압���)�f��Y(�+Q��_�<et�cLc:v"F�'O��'�awA��Q��&�v=Z��:�4ﮗ��DI[�GY�K�E'Ip��^%�մ���/^=�s6��5L�f�VJ����rꆊp�<H<�Iu¡��xg��h����ss�0#�d��=M��kFi��gپh��|��j�p[����6#5`�^�4s���z�=�o���h�����B�C�op�p��}�AF����T�zN5�{O�Ǹ�c���r�p�{�^����S���V�L��Z�ԙ�P�C��S:�<}���~��oI�s�.���� ��<a+�ƒ�.=	�Zג���^�fx��a^l��}l��#���r�+�J�;�ǫ��*����<��债��}]O��:��6ף��c��� ��Oi��S���Ї��f9g��l�>F���[]"�MpK����z���P��ur�ِPqeD��[Q�[<=��:k5y��(;��Z��i�w�:�kw^�lb�*$ؽ{��T8�42:N	m���r��.7�r" �~����{Ik�yt��X���U팶��pC���Ӥ}�o7��l�k��8��jZ�T�z��K���s����fBp���d���6�Q��[�x����N�O�z���^oo�=�iYk�%��+���2'���U�X����l�o<�g(����A����W�]*��b� ��9�i;�Y���r?_.�bӜ��9 ��t1{_����^,$łg&��CF�J��>@җ���2���W,����F�pN��R��g�,�/�z���F��,��k�0K)#w�py!y'Ռz�AƗ޷j9G��9MS���wV9t7=O\s#lud����cxY}�84��b�L�6Á�hrl�;��[���o`�\����D����q���`ކ��9
�1Y����ؼɻ����݁uG���;+�2�k&�D�����6��޵&��3u��p߽`�z�R����3�y���;4��Z���:�3��x��C���q5��!��M�}���X�0��jg?�WB-�d_RbU����g��$�.�Mf��V;���$��ɹ!�JV��'�Hr�a=�\�]u�#N�]��nP8����O�<VP�
�&�ے�ڙ��� ���(��T[�=�a��#���Υz�sھ������hr����{��-����A���̯��1�_�~5g�[�c�G7|��qajW��֜�-�ůd��g`�ʰ�����C��V����G�68�rMў5p��=�On6�>�`ϲy��a��(�T��W�62��Q���R.������ǝ˞�R�|pu�ڍ}����;�X\�=�+��H���u���t��j)]�P�M�D5Kk��롡��:09�\�`_� .�Xٞ:�9{5��;�o�A�a�틄��>�MK��:��a���C�B�R(m�1�9;U��X�5~^�_W����>�S*_����AB�E���z����=�N����b*�ёg��d�=�2.X&rO�넷�H����N�kt"u�w C�ai��N���Y��s�"��s�n�/]vzi�{Yc�ྊR��a߈��}w���j��;h��A�r5��^�G�z;4RJ}�r���N�(��9*]5��·s�z��T�|��/X.D2eN���}pk�Y���a�?m�3�����6���Ǵt체>l+{�M��`������U�'Z��3tǁ�䆶f}'���gg���Coq�0l�K�W*;PG5L��V�����������v��K��'���hrt���1ۮr�V)[srv���x���w�Z������v^�>�j���7]�w���?}��P�����t`y\@vV5�=:�׾�z��y�����ɨ.��ۏ�n�0k�C\c�_9�k:{V��>V�F�s��5�M{��yt9䁚��-v�/z�jȾ�-�<㥓&�>[HO���ʹ��R�oJ��=�q�h�����)�����E�+��ܹ�Iղ��o�z}�#�=�&V^u[_\E��0E�w��oJ��1�I�|c�7��\/�ҋ��k�y�T��j����V�`ڃ���q�t���Kc�lN��ɢ]G��Ǫ!�O�8:�h�>*ٵ���g�2f�֭!�BPwD��E��2�n_.f�[F%()V2�V�w��s�X)�i+%���sJ�%Θ۱YP<AmN�z�pӓ�G4κU���nֈƯ�tf4%��ޝ�
��� ��N3P��α� 3ڳ�s�Wm�ׯ�������/oQ�)=�=�M�2m�����|"Ƀ���b�hw�\�H�<i�z.�zeZ������n�5��<��ii�ߦ�F�.���%Ʌ�T�hubI�i;�o)Z�O��;����j�e��_\)�G���o(cJ`���R�}A��/���'�a��̲U��K�r����qYި������Q��N�olf���i�=uk���=� W[�O��?}��z�P�#����짲Ǘ�w����O=ɾ��n��S7-���oB.9Ӄ�pz�V��OJ�|Y�w��2�΋��u���%�r�^�Bӎ����)J��U�W4�'�R�woI�DڧH���vg�W�_k{�<�s��,�!c.������o����9V���+"��E��~�g�~[Ɍ�zAށT8[ӛhI�	���]�֮'j�_�nA���wwTى�[w�M����n2�&���!V݋��ޛ�U�9+���k��l^��x!'<x�r�:p&k�l��Ĥ[[�n�_C�|�3k����\8%%��qg��R�<4�p�l�HE;�_B��u=ϼ1'<����A�o���3}3y��c�1S�u��Nk���	������W�����w�z6�t[�;0=d}rF��ŝ�^П��
{c��@��\�F���k��� �ʒ���BsV �'�(���'f��p����Rc<���n ��;�6�P����*�g��]��v����Qv��y�Kq63�u&���_�ӥ>]V�}��L�IG�o�Spm�cC���S0�V����mD&ZR�j�8����}��wb�7̒�/�����1�V��#����\~�u3������ȹ#�2���D�Ϫj~ɒf*�Y��ӱF�/�ύ)9m����O�j7'.~�vi�P�<~����Ί^��dHL�5�S�{yP읋 �#<�J�-�Ff��=�;��C}�K��MS{�Ö��/�<:�eڟN��=�ڳq�ְ�2�wAK4;�Mٱ�F��f.q\�8o}�g����l�pdڋ+j�u�ܫ���ڝ�;��0f�<��A�h�CW�]r����:8���޴�����&ދb�Į��\�ř1*����K��{�ó����i,a�:R�s�V�@���6�sc������2<�8�!�������:����s��euqj�k�/w�]1�]k��J{��w�������熽I�ckҔˇ���^8Z��&�D�v���:���T�����w���Z�u�e9��J��ً��fΣ3�by�Fv������D��ჽ�0Z�|�ޣO��z��=���N�~�U�j��X	�wAz� �N�zr��/XST�d���G�c����~ך}bR@���+7:ی�E��Z�n�q��Un��mIE�֣R���\
�M�x�7�Ӈ(p��F��*�|}|����x��/7)΋�<���٥秹T^�K��?a���@�Th�hv/��\�?T�4����;\�>3�Z/�c��"��YS�8:ƇV:09�T����h��,�;^�v_�t�A��Bo�%��3r�A������8
��� �:�7d�������92t�V�͉h�� �3�)���W6]��B��͌�5%^:�1}�]f|76���N>��[al�QF��OV7B���v��Y�A�R���vj��5��T{x�I�7�x���(�={�)P�{$�g @� ��Yv���SKG_P��]>��iH[�fX��y]\�m�Z��bY�i]������)�`�Z��ʻPLQ��Rg���νܓ4"�L��)�[���R�⡵�^E��U�Ίz(mS�j�:*�f)��b�5��O>k�47�;S%x�u��K�k.��a��L��/c�5��b]�2f�&]�0+�Ļ.�{-��Au}(�.×L��e>�r���,-Қ�8��������I�v�����YjTۄm�-[����m��0�D�&t��yВA�)�!k���3���A��Y�zZ�3&QΡy9��R �Ns�8���[��B)��T�z&�yjoB�k,���vH��c��.ڮж�.�CF+~K�{7t�0s~G�j����}HV+�)���fsg&N�$���J1vp�ĺQ�����v�f����pEs��bY���B�dQ�@7��yS�is�lc�0#���N7��=L��=L���5�ݦ9����i��	�9,�r�J�N<��Z�}����"ݢ����[�ʾ�[�l��]�f(�Y�pE���q,yig�/h���v9��|t�%�RZz�|v>�v���wkP����츫�2v��"���΂`���m�Cxs²��I�I�3�gS�FۖU�	��%�Sdj�r�1mV�eɹ�Y#S6i=�/i02�V�Q ��W��������#�
�ֻ锾/��������������ظ6��L��N�\V�
Ë�Y��.�wD�6��3)>�M�W`	B_iΰ��}�Tㆲ钚�jѨE��h05ᕨ`}(���-���n�d\�SҔ���N��S�fE���`��iA]n����[DE1�M6$�pʽ�(\�3J��52s�ءs���ܑ�y��lM��:�9��h">a+�xT
���̬*Azse �su��S�ݵnfQ7�gj&du}��U9�� +`�4]":ֆ��˝xo�Sˀ���)-m�X�&���X�*���=���]n�����w�E�gg6+�3Mq�L�_u��	���`�����;��IHI9f�eH��r0\|.�(�T
�Z,�W
%]j�����f]�T��*K��Br50���ف��)�wi��-��?����pF�p��(xVl�2�gGod'-5�^6*uh��6�
�ɋm]�	>pPh&7U@�7�rǭ����o�����-���K��״99n�d��2N|��4ۭu�֞�Z����Qh�9��G�>�����jE�"�P�m�A�JU*-�h�X�+J%E��
�1A�Rڠ�TFJ5�������TA*Qj,UQPQaEk%��`1J%UQU��j-�-�"�E�1XŊ�-��б`��#-�PX��b�,m�*�X"(�F11�$�+[E��-��UTX��EQ�ČQkDEb"(�
(��+b
ZQ*QE�"���QE�TdV# �R�H��
���)PX�(*-h�X�*J����X�[H�QQ#X+�V�E�UUF(���* �*�c"2��b��" � �ְF(1Q@D���b��ڡR���jax��+����^�b޷�#3�\���`�c��9�-��}]��2�1�.��(M5���g�ܻ��Г�fkL��O��T��yt�H��jX�v:� ��s��������O�Ŏ3�ת_O`��=���y&�$�y0M��)�]-��2�n�jTF��_؜G.�}�7?f�7tR�t�K���*�I���;js�:��Ȑ�0Ǩȅ>�΅�aF���y�Ľ��X���-�7<߻�UG��)���,��*��׻�o�^�`y0o#c�uf���̗�g:6�>�^��W�.'�G]v ^�@[?-^ǧ%J�r��آ�<�{�#��$L B����&�f��˚e����b���I��)Z==�^{]>P�Z��sς���緈2�xXiШ��~��/u������G�E�C1���8��z�Q��<c������u��a�hzt����A[�� �k�N��R{张��$r��pϩ��y~��-�V ��v<��іB�x�ӽ�y��+�����9o�:���`�ݬT����ݵC���"�]�kjTh�m�(�ol���/�L1��G�[)��LL%�j\f}��,�6*tC.�����<B�C��+}gPs��*���"�H�����|����;��U�e=����ć��=u.ċq��
zq�Ӥ_k��H����r��V��؇Ӳ�=�1>͹�z��Gv3�<����E��q�{��>8%��o��z0�s�=�'����w9��^n?$+ժ���C�R�~��CS����$}�~��a�dj�uk]�vZ]��p����̣Z#�=�o&�{˞�����b����}���	͝���ɋ�U�"xJ�V�e+���?9�}:�^�MNJ̾T�q)fdw�sTk�i�-����s�A8)=�sk����.U3�E�O����\g36��b�s^(���@��R��x��ƽ�yI����1	�t�c�S�,����E�&D�mU��U�ӭ[�[W�9�鹔�Lk���Sγѱ���g�Z�Q�hp^����%��Q�Egٙu)������Wv{>;�PK�X%m�&��/"�N��q�P_n�-�WN7[����/O�OFr��C�$ޠuh ���Ԟ�]h�\����݊]�a��dʜ�%�яM.���Y�Y�����s��r�\�m8��?� �f8 �]��w�[*/N�0���W� ��A��/���ջ�D�F��6פ�K����D��K=2�I�=IOr�*�('9Kl��ϯuy=�:@�*^��疍��#.j_��xŭ��y��=@gsw2�c1^C'�{�u�f�z���/E�X��򦢷k.6���*�0m�r�fI3e��sb��]�M}��,�{����Ϩ��\�}�%ߓY�J�՛��>�|�jsj�{Q��O5�g�ϒ�_��U��7���~Q��r�VRސz��p9o�(��8�~�ӽ���^En����[�ם�fȕ�cJ�Ay(�S�ʛ���ΙN?d��|����/9�?A���X�O>*��.R����u&�)�]�Ћ�2�5��w�����_�k5��Ɗ��<���[t�|�x2X�F,��؏!Oo��n�5L��gU	:�����Al��K���9�rˢ��Zﻨ�9O�Ozn\iY���w 80�����`�
��4���t���l�I�jƲ&��ɱq7ϰP)�&��<e�C�%}E�}�����tWf��&oc��LȬ�]pR{X����=ï�ɡ���"�=���OsK�I��H���b�rYM{I�s���>���}�ٻ�gٵ�&t��vk;�[�M;�`w�T8�^Mkr�������5��*��%�ݿ�x�����-G(��zd힮ȸ�	>��+Z��Η�� ����}���Y~���7~O��&G�Cl{Ӻ^v�,YX�j���û�vw8��e{������?��&�>9��<��C���Ӵ�d��s q�d����}��QW�w����g����	���a0��0e��,���:ɴ�3�`���O�����:�3�ĕ�$�M�E�ڰ*d��'~d�!��X�+���}���=�ML�������O����0�aPɾ��$���py��,��I:�l�sԂ��M�g��O2d9�I]2N瘄��'�8��}��\��m����+?'=_�?U1�h���~��e��<��z��Y:��7�m!���XM��i�N�Bs^��N��*;�@��l���6�y��|���>�¶�o�/�zWL�=Y��9k{�����+0�N3ڡ��Bg��?2y��}�6��<���	4���l�~d�3gw�̝J��k���7�O��@m}�W�x�)�~�����v�Y�3�5�ι<�^�f�4�x���okN�M�Z��ױ�����[�}!�{���f��E���h5Ĝ��mW*�W�Q��[�Y[-���3d:VZ�����}DǼj
���1�xkƝ\Σڥ�=�0Asp���l�km�7FNw�4?⾒G�����s��>��2����Ry�?2q2�gY2��d�%g�4<��L�a��,�Փ�:����	ĞC���e�|��2u���\��s�^{��Lk��w�~���x�&�7�'��I�I�gVL�?��R~I�g'���ɜY��*~���I��f̞Adι�):������'Ry�7�z���~�����o��������L<]��'�On�a4��m$���q%a�C�h|���C&,������S�hy3?P�	��g��y+�g�����緟��}���c����*M$�ʙ听�a����ē�5{��z��Oq�M;d��q'XN&f3�*M�>ed�����'R�d�C�s�����v����3\k��k\�����*e�m�>�|�Ĭ���i̞���'�~=�v�̙I���=I�M�N���=�B�M���ĕ&���B�u����Ly6����k�}����9�@�2e(�2������$�㟰d��!�{��������`|�rwX��M2e�]� �ԚI�G}�N�Y2{X�a<��^�o�޿�
Ʈ�z���3���ƀ���a��Y4����|�i8�जI����N���`8��l����&�����<��	��Ǟ�i��'���l2�=���To���t�����;���eR�<��o8%AB`��J�Ԭ��@�N��30XN�m?L�󄓬�߱��<�\�2M�Cس�&XN\��1�+ؿ{'jo��w~
��(}� �G�g�M�gP�C�N��8���T�&Ӭ+'�~Ru̜�L���d�kvp�̝C�Y�O�:w����]@1=��^��M�V��>��������L<�9���'Rm]� ���h,�wؐ�d�i�I�wX��I6��d�b��M�{�0�u	ٽ>�+�ó��v�6 �؆���q`��|D�mn,���:kl��}}����k��v/I�W�:���9[��>w���Ҏ�ݮym!6K/�Z2�7�96ax��.���7��m�u��
�c�ζ�),���Tƛ�@o��.��:���$��YL�� ��8v��·��2e��g���L���Ǚ&�����0�L�ؙI��}`��O�Y���'�?�'䓩3�bK�$봋'��}�z�����}����?o�~a:�O�������O̚a�o���e��jo��$�V����,����O$�
C=�&�u�iXk��&�~�8���������Y���o�'���\������$��"�.�:�1a�I���ՆY:�gT�<ɔ�a��6̲u��}�'�y�f���,���]��N%d3�`W�W�u_�w�o�����Ms{[��k�a��7�~�u�?kWI6��ы	��eC�&��٫��	��0m2��I�gx��e��:��&���G���]���n~���+�i��M�[���~d�VC���i�Y6�'ǻ�d�&y�������'�d���ɋ	��2̘�����6a���8��A@�5�I�<���}����{z��ce������c�]��O�{��e$��2wvG���O2u�O��@�����bJɤ��N5����Y���ɜY�I�T�fè)'��3}�>������}����0�((>�!Rm��Y����<�Lw���4�<���A�c�a����u�|�ĕ���(m+'�fqd>g�N��{�{�W��w>�?}���;���{�(~f�
I�����O%`g�`��Y:����!P<��wܲO0�{�̝~I�O��q$��L��u��3��J�l�K�&�{y�3�}�~�>�y��VL���b��̝L��O!�a�'�9�u��X��J�̞~C۲��{6{�	��ǻ�6�L��d�v���N�٬�~������w����Y'���+2�O�T�Aa��C��J���N�ߨq��N9��C̝��=��N�y��1!P��E�G�p��+�׸9j�~����� �Dm�����K��%�Q�|x'�����\{D̋&9q�{��<7u��:�}Jo�_g�aY۾��Zv��t�qzf�ew\T��ף�1��g�S�{���0l�1�mu���T]<YkWL����3�q����쬺�
r���#�?���������o���C���0퓌2������&Ok��i���IPP�g�:��P�N$�'�8,��:�C��	�}9��O?$4�6��N�j�~�&����~i���I<}�m�&�2�G��<�d�L�̈́�?2n�"�:���T&7g��J�P8ì�O�XN�y?w����W��]tl��E��J����z�h{��$����d�	�Gq�̙a��$�e��2����e�'��RN���q%J�bn�%d�VOؠp}_���q8�^���l~k�ҳ����Ogx�1a8�'���&P����d�|��~���d�׮̜a�����M��=�y�{4�>�pJ�_����^s�{��~�C�_|���I�O�<�L0�`h��~d�'�����&Xg�����~=�O0�$̝AHfw؂�Rm���)>d�_/������c\�������㬓i=>�	YXN~�$Y<����e��~��N�����4��>s8�d���$�*�b�*o��'Rb>2(g��v�w�{;��¨��t�<H,>d�{8?0�@�sX���;�x�d��O&a�ì�OɓT2��C�`��d���gx���'�h�q�hV�M^Rmg�{%����-���]U�IS��L�J��,�N2|����Xm���q�$�&y�Iua:����&S8��$��Ψe'XO�:��e��:�������,^ݐ5>�k��>���߲��i0�{�<��m�;�O$�+!�{�d��w�l�d�5��O2d���m��P�~d��bβO�S�z;�\�����n)K��Ѧ�D�|2�_��L�u�P�� �I�P�p�<�8�&Y'��;�O$�+!�{Y<��i>�p�a�]�VO���}���c�(�gR����Ykr�O)t6!��^�d�fY��
ΰ�V��4X��˞��7�	lU��7�*�+E�=��0���ӫ���[o`���$͗��x�O�s�+�H�=k�`�\$ə a���cM�X�v��7Z�|�k�aa�{���?<՟�����k��9޹���?������I<ʟ��m�$��f��Ad����O%N�8��0�;�ɖ�5y��N}a5�`�'�:�'�}�<�>w�����y�w�9���Ǵ��������>���VL0=�ed�ÈdŐ�?2q��a8�O�l:��`���O%Hd�1'Y:�3���<�8�<d�a����N�a?^��������9�=�g��{��$��O��?���q���C�l>J���3��?$�2b�m�d�a�����N��2}�AI�O}C۲��/u�i�{�j������>�w��̓L�6�i==�T��2�!Y&����%a���a�VN��RC�:���:�?Xy?2N9��C�:���'��w[�Ƿy�s��v�޹w�x:��L�g��H(C����d�&Y5�`�d�M�+	��&Og�&����IX��7N!Y:����6�Y<��,��:�a��~���7����}������^
�a4�O�b2o�!�_`>d�'�����N0�����&Y5�`�g�4�)���',��J�u���*
���Jɏ��u�.:���ߏ^����Ęd�{�i���46�I��sX�;� ��d�xÝ��,�a2s�<�&�q�ky2��MOka�����Y'P�����{���~ß���w퟽���s�T'�*L����i8������u�l���<�u2s�H.�<�w�N��z�G�`�2N���'mG}�<�d������6�.���y �PC���W���#��*I��ĕ'Y*O2m���'P>M��&��y��>;�^�eϷ��	���i'�N��n��d��׿��~����[�������)�`��O�Y���O!�Of�d�a��%J�y�9dY9��N�m���d�!���Ӵ�d��s q�d���d~Ÿ���Z5�}��7�U��ȯZ++Y��p}�or���}�b���M�dߏ�s~J�D�c�x�j=��4Ϯj˘�����m�&�3x�@�ܺ�3�|��!�T�g^<L𮢶M�d�;��9z`��%�� ��H�����m>x�;�o7���0����pm'�L&OwY:���}�(u�iXd�AI�'�w8?2N��l��$��ċ'�`~���I�I��d�!����ÿk�\s������\��c;�u��I4���b,�C[�<�m�C;� �J���d�!�`4��6ʇ=H)>d��~�$�&NkWL����&��<��9�Nw����߹�o}�RN�fP��L'��3,�aԟ� m2��[�	6���o�<��m��d�T&u�M$�M����>d�&M�I<��;�9�7�n;���s���;�����C.2���ń��&S&,<�|�fMP�O!?��,�b���bM��O �7�i!����e�m��<�ԨN��:��M���?uf��|���~��ޟ��C�}���_!�����>jO̜L��gY2�Şd�%g�I�'�aC�'PY3ϱ&��'��[�u'��;���$���=����s�~�>�|}�}�k�Y4��{|��O2wt�gؓ̓���VO�I�'Y�P�'�O&qgXN0�����L~ـ�'�Y35�IԝeL��Z��6n�ݿw^滜��M$���;�|�N�{O2u�	�oO�2h��Iē�q�IXm��Z2�y�P��ɆN�ئ&��a���N����۟~�qu��g�}η^2~J����T�I�TϾąd���<I<�W��aǬ�d��I>xɒ{8��'!��J�iš�+'X����d�g�ﷷ~�������9��3��(~L0�0�>ohm��X��Hd��}�bAd�j�v�̙I�{8�&�4{�!:�2g��(�g����k�����g�u[��s�hVO�,=l!�O%'�u>͇�$�~�u��̆��̝d��=�䓇u��d�&Y5;��4�"�ߕ}��A��߀����`�ߞ~�/i����Y�j{/&�/ޫ��3����-�+k�|^&�ڽ�M@�������n��D�� '�ht6�����*�n��Qu����^b�#��Se�{@rH�*[+TE:��W���[2�Wm��Y�uI�q��1������ �5����o���+	������1�>B�q���I�Q$�O'��I�w��q���^�>a4����O�L��zɦ`Z��s�y�����=��\�����2Ͳq�_5�N�Y2{X�y��	PP�7z��y+%@�N��(�u��ٝ�p�u��ì+�O0��`�$��9�tީ�?���?~����{�������a9��d�M�k��<̲q�4{8	�6ɓ��,��~;�IR��&����Y?LRu̜�L��'Y6�݆�$�'P�}ۿ�qۗ?~�~����޿}�]��M0����	�u�O{�y�w�0�ԟ l�̛Af{�Hy�g����y&{�IR��7z²q�LY:ɶO~�{��y���n�s��u��>��α2�L�C�s�a���̓	X~�py��L&g����AHg��:ɴsԂ�I6e��}�������}+�k�f�v�o��};׿}Ϲ�,�z��N0�z��Ì�d?gX�~d���,��'��c̓	X}�y�Wݳ�8����bi'Y6����Rm'���X�����w��~��s{��vu��'��ĕ�I�;�,4���ɋ2M?&ua�N���'�4��?n����:�����<�}��Y%L��d�VC߾�o�9����Y�~�9���9��Xi��Xo� |��z��'Y3>�$��m�ɣO�2̆(u��<�5a�a?g�6�d�O$�gx��e��;��L���}�;��5���o��s��ί�ό&�'P���N�d={�2m�O�w6��L���B|��ԟ5��'R��|��>1gY'�S�0�	��q�:���������n~�6����-������C�M �{?�8��^����i�w�;�	���O2q�'s�@������%d��q��a�>1d>g�O&qgY'�S��5�{�ӽcY�3.-LG����HֲT)G�Q;Нΰ0
s6��An݉8H�}@����ޛӝ�8d��G`Wc
ֱ�����N	�`<0Z����-����p�*ҘŪJ��^����ޙ��l�=�\�ك�S(܏I���CL�Mr�3EǑ�jh	uh*'�^>��I���&Q�������JИ�%g+:���8�l�4T�m���-����|�1Ĝ�����
CErR�5O��83�h�����Aס�L&cT\(j�to���F�o���g�lb�;���1��I�+��ʑ=�4��p�X���Kfk�.�=;T)|������X�ʝ$kw������
�q��L�ͤK�rU���-�+��ޗ��&qZ�S,�&�k@ȹ�Qb����LP��م&U�&���L ��]���/V�edN�E|f�UXE��顥i����6qT��j��j=�O)Y�,�A�1rQ�]�C7XR����ͪ�����E3����hb�::��d����0�?9�߱>�n�y���g��;ؗ�`�s��nMWW�+uV͋�g�d`A('4H��Ս
	CU�h�iĎ�:�â���z�?r���r�}v:��v��aM���ݫZ�p�<$����zqc-Ҁ^(:��4n�ڋ�G��H�}Ѥ�0:���Y�R0^��R���JVZvM*ͳ%� ��h��\�����}�e*�sSz
)\q)|��:��@�[g)��SYW嶍a�Z+�k��X�=�R>��\�m;�k�w+��	mD�u7��Z���j��}�`��=s���*L)P���F��ɕ�;c-��m+��06���9q�n�`EV�(�n��)����Y��N.�\��Pވ�,�A"�E.�������s��]u���G-|��o��]\�w{Y����Prf�N�r�]Mἷ��)��o����k5e��O5��CLЖ�ǋ&�6�V@��N[i�swCAͰaH����`ܝ:ėCG'�Տ��v8m�$u�ҹV�ð��Q�:��>�\9A|�np�hj�����GR�u �R������&��k�]t�sQAfn%���Q\����]L�bۤV��t��5���}nFq��duY�[6�)�:�jQWf�����F���L��×���xݕ۰Gu�{5�C�����"�?-�'p%�xm1�Z7dθ��ok�h��{��ƅp���i�-.�����Rەӎ>ح�Ȯ�	YR�m��{&���p�b��YutK��{&KwLU��,:�k+�'EVpw�#�bH~��(�=��`:0���p ��K����jR��
�������,�ܧn���,5��-I�Y{�'W+ɏ���(�]��j�ԇ�;.)&j�hAS��ܫF�nT��R̤�j�&���n��Ch#���l*�EVUXDjTQV*�$QX�2*�%�UU��V*�V"+Z"%��
(,F2�0Qc%J���*"1"�*�T��b�aUU�+h��
,j
F�IR��b*�F"�T�E���`�b���X�")�UY����PQTb�0D�,ÄE�EG�#UDT(�&�b"���X"(VV(("�&,���VAAE���
��%V"R���1`�PUE
���Tb�DDFE��	�U��b��W�
�QQ��m��V(��"��b��%lUQŕQ����3�K�k���qϱ���|l��T�:��6
Tz�:��3��tyF'.�$kc6��U��Mg<y�@T��%U@��5�}�}�ټ����u��?aPRO韰���A@��'�:���w:��f�3,'�h/0y���&��@��d��'Y&��8��y��9CiY?$�3�w<������o~��}�c;������O�鋆I�f�
I��xP�'R�2s���'R�'~�
��?OwܲO0��2u�'>��'�d�q'XN���y�����w��g�����}����x�4��I8��RC�'S!�a$�fO�<��'��!�N�`d��J�̞~CG��
��?�'�a?2{��d�&���{��]~�KV9z�}_���N�߷,|k����Vd�
��,4��d�T�'u>?P�?$�s9��'~�hi���t�s	����s��yu�?lr"yܟ��Y�����n��o>�r�'0�w��*y$�v>���7s5�#.�>�����b��^c���U�}A��RW���=���c�~�=�}7���<�	k;>f-r^�"�?|�Q�]u[j��m��~�>��n��22��o}��-G����Ohۿ[����'Y����͐=���TN���\!j���_{a��G����|�����}2�9��yI`^����s��Q�vUi(�x���]�s�	"}Z�8&<�p�H���t��7�m�u����I�\��Ʃ_�u�J�*�,yxS������l�^X��_�=w�%t7}������8k�O��B)�m\����8%����O�V�C$��&<
"���l"����Oz>�k�Bӗڳ\�/�UU}���<���oԻ~�TC~��2�x�5�>߲�veV����ݒm*�a��O�)�(Mj��؆S��z���ٵK��[��B���6����������se`Ց|#�^�\2y��9���ؽ�ؾ=�:�؏�i���oӴ�ڴ��y;%g��f�����Hds��'��~�����>�Yc}�L=��ũTV�QZ.�ѫ�n��mIT\���[M����D\��8r�j��r�A�md�gU�� ^�)g�n \��F�!��z���Z���/�<���W���vM�~��=]� t�{�Q�*���Ν'y�>��=�|���`�v:�hu`VƁ<���x�*����J7y3[+�SS��R�L�T�/y�Ա̊�AՎr��ե��bA^-�WH�V�Z����{����ip�&(��<�a��Y�JK�=w���l��w�=pz�)�2�'���z��G�q��F���f��u7�Gd��a��=�wwe��F��X�DmF���:>B.��o_\�mml]OwgöԒwRaT2om��}a�렭"
��+f�v9r�OrގPj��Ƶ�j�-�X�������Ȭ�G���������t���v��E�&E�&E={���S��^�=^��u�1�*:�_�N�osaz;�cs�;N���1��ެ*ґ�fvɈ�]5gmvT۰����nsϋ.���Lu/m��DT��������ҳ堪�GO���\A�T�ò�/}j���w�-��ད�,��}�|�@<�2[io��s\�`��+�q
�eX�p�s6���(8l������h�(O��1��R���ً�΂����S&'���u�`�ֳ�=^�;^ŮC�:Y1���oK��</�����EZFH�}���d;�y#='az�_^z1�jƛ��F8�D�|.ݜ�'��&����eb���}�Q�ؑ~�
E����)�s(���&�c|�-)"�M���}��m]Zޫh�� ����'��*D^��h]�����QJ�L�n���"��13��v�int�<���%��*�+����q��:j9�%�!Z�t�}cM�L�Y��V��>��Zݻ}�~6�oYd��3\���A"����6��X{���}ӫ(@���7ک�M�g��>�����17:�	S����L��|&��>��*��z�_[D�N��[̗lǫ���+�{���d�.8�8�qY1����C��� �`>�^�˸��G!-f�TczN��R�L�H�����*W���߷�I�M|��T ��=�J_حe+�|��Qu�r:jC�_��R�����I��"]WX�]��&��JbW����R��5�v3!���/8���A��:�\�L�x�C]J�ϐ!��[�[8~���'�j�7;����jk�{Oo�����꿋�k�{����T��Š����o�F��c1}&G���p^��P. �]r����&��٣���}f�_��w��/l5�dL8�A���³�!�X�����iNr|��_I,,�c�ܦ�jǜb8�p��=3+ҁ5b�����0^��SEm��EnF��f�ڹ�����H�q."k����R�
}C4���`{"�����Pm�A
�NAp�/�5�w�f3�/a�T;`����Zp�d�l����J���.�P��ǚ�����i�k��+��^��.���UU_W�?%��z!��Osڈ>�EM��[�ٕ�xŭ���b�q�,A���|�˔�XG�q�D޿4Ap�[�q�h��y�by���/��X�;�\�m���>^o�>�-jC ~�u���g�����d{^� ��c58���}�8�rn���א�4�s��3iGf?&�L�5r�V|�H3[�\ɂ�w��5�<�U@O-�]�ғ�����_���]��Dƅ�oC���Su�g����=/��vE�p&�8�-v��3�t�4�U�*T���־�|���|�I��%�N�Q��G7�9~^|1NW�uJ�Ϫ`�������IO-Z�q�\ٗ^��wTAs��Z�M�{u1���&>���em�t�1b���(���G}�j�,�9Z���Ȧnt�5	9��2LQu�]mJ���,*%�ÒPn��'i��bÀ�[�Q�pԤ���!�� ��=�yP��bXzܣ��ӽ�9�@�,�Y�%J���E�8M!�W�)�k[��f]Ar�����T���t3�&K��Ev��1:��=ӍT��:i���8�oջ���$�����.7�{�8�w��>��'�KY��1k��tȐ���~�ϊݼ����n1	�ǔ�d�/v�o��R�s�o��97fY�q��J��w^�銨��Oǵ����<:����#�m�<�mѹ�1l�{�.6=q\C����s�̣Y�ϴ�yT��Ӟ���Jlמy��	�[�U�.�T6���ިl�Ӥ}�
ӳ+J�8�P�Ew,�N=ɩ��|�g�{��S�0k�O)j���ƻ<���_[?'��f���#���p���SDpo�u�1��9���~ԃ�=��a��,9-���=Wҭs]����3��)�^�K#��	�w���z���rޝK-�9=\���_#����F{\��E��w�-Vt���w�퉾ZZ�l~f�9%�@��uZ`���g�7�w���}�ڽx�����S���`l��c�/����d��;Ē����6�hw[��[ �8��٦#u��~*WD]8��7�D����Ken�Q:��A4�)���wI��W\YE	�<�tc	�Ml����}�U}��o�>�<�H0��ۈם��6v���j��=n�a��su��#
�u�<�<���~�<%�|"Ϧ��c�huc��S����'c����b�y�:Vޡ�7�o�	bf�Y3{09O�����4Zb{~�S��s%Ǎ���f��m��NS��_n��x�݄E��&t2�� t��oJ���V�	Gy
Skw�������wI��r�Hd�C��2r��#-=]>^�}�� ��SW�[��^���n7-GB���uHܓy<=���Z�u��k��"���-�����^�/��c]J������z�%K������;!���rz#ʩÕ=�یpz���Y�R��a������CW�!��ߜit��ʓ��3�Y�z�'���(���rw ��,����O���h�8 ǵ���p�=�{r+�Z^�q��ڑf�u1��6jP��5ܳE;�/r�(���r�����"Ц���GN��@N�T>[;K����Ū��*��/�W9Y�ư�`jq�/�Au��o���";����)�;�0L%R���:l�yK�����.$��U_U}P=�WyG�@��*o��ﲫJ�EL��\~�n_y�K&=�:�
�����~���6��#9j���߇/i�϶=�8��F��o���Cr7=\�&>�~���yw�ߓ��i��ޫh�H�V��l!�s�&g=Y�f�NbF�zwv̖������G�'�*��U����_U�3O��s�J��9������P��ez9�:e8��{݂��[`W�4���3�;�H����/i_��H&��΁�|��^�"|����L�o���k#�M�k�B
�D	��� y�OrM�ʗ��鞑?z�+ں�U�W���<\7S��c�L/�hszi;�i����zv�7�g�`h3�l~��7N��T�R�BU�B��A���w��ڌ�돖�Rz�y�ޘ�8b���7&rA�n�k�Zy����$�FX�骍��z���N�#�!�m��NT���k"�QFLMlt��M���}��)/jk��ⳮ��P�d5��Fb��h�e�Y���o58�07�
��a��+0��C�����,�t���c�'���]u�:��%\<�Ω|7�{W����>{9��Β��{ߣ�y-gc1n|�\2)�`n��]V\���Y�#z����S��3Q�:��l̓������c������l 7�7�C�oC���cbm��[�������=����G!ߤL B�=^��8o.�Ͼ�gm'Fߗ�S{�w.og����2�k�/'�{���_�G��ܿ�[<�S�I�c�x��ߕ�T�����/�;����\^�V�b{��%'�<Cp�k|=6!�*2����+v�����ԙWw�7S҃���^G9��pAE[��t�OM�G����/z��v*~�ёNԨ���=��s��X����d��yq槼����gU�ԏ���	ũ�}��ٸTY�j��������2z�(��S�s��z�k^u����;�nN��9сe^�}|��_[����lc�/���8�e��콏�j��ډ�]l�L�J�d9�{��A��|������i�uu���*Шu�dL{�a��x-��Ĺ��.��ou�w�̫-Ln�b�L����SJL�|pt��캕�L��N�3��|���=u���}��7�'I�~o���j�����[@�f�<�y�3���jP�o��9��r�L��N�|�YS_��_�W�� OjլW��x���M����b�U��܄������{w0kv(��?����뚻�w����g�{��w��z{���Nx��(���;���r[�}��i-�&�*���������<�y-gc1n9,�dHLf^��LW"�^<�d��n�}�xJ��}u�����I�n5��z=2�.������ܷ��\����m�ޮXf�B�Z�'����j��к�7���㛺��`��zя;/#�i���Y�J1}]��+B�����ue��{��Pc�W�0�Ժ;3;+�셯xboj������{��D�q���[�??y�s�2��	�u�z�yz!�X�g���!�Rkɯ4�z���D�]tD�&F�t�B���EllY��+ANx�,�[�k�H�qj)}65�+{�B�9w�} 8؍]�S���T�h��xu�LW.���抶��p$\=VJYz�d�������Z���D�����I�X�ybNt��j+T1��Ӄ���˜v�q��t����`�FT�.z8�6㺻�^��U������T���x,�oh����4q�$�J�����J�dBJ���;�PKDe4�-�ݶ�N�-@�{2���vs�^�;���-�(�N��қ5|�9���Wd\K^�;����J�A]h+&�b�����*��GU҈Y$�,<唓Bp�ͭ��U`����e.=N*�՗�VdP���!ɂ�n���U�^��$ٽ-_L婼�Y�ws���]��N�:h*qux�v����oz��2F�Wg-¶���l|�nV|�te�{|�h��a��<c[� ���y}4��u��b�Ť���N���Dr����0�'�b���s@��6�D'��V��KAvO�s��`<�(���C[h.�0����z.2�h�ۏ9�@�@�)vJ�\�E9Gp���Z)öl���䮲�/C,V�a"��#�z��2��zZ1���+^��J�>�P���'����[�R���:hf�Ϡ囕-�Z�cb�r�m%.�:�/b
�ȭ�-N�<+8�6;b5\�/�n����j땎\=�yOt�K+C�-Cr�k�JvnJ���U���.��%��+-��X�}50��عX/�.�ʹw&���1��6V�PY�bm��t.��2:`V����
��[���ս[)T�p��S�����!���+0��ND)�pl���E�(��Cj周к��f�.+G;���X6�Zǩ�� U�ir���
]{R�C�ӝ�],W���*p0����G3e^(�V���;�I#�(�)�"x`�jŻ�w�����H �>�\���=Lݥ.����9JK���/D�q�jg�UhNXd��7�A%E]��V �ksI���Z���̾�
}F(�s[��C2����49�][W�GIOn'�:�]Q�R72�Ym�tr����sY�7V��۸��sjP*;uNu(k�(r���BY�3b��p�k2A�򃨰��	�4zh_)�o1R�+��9������u��K��}��DH�t��Z�ѫ{Pź�fvQ��m&����H��{yt��54�9.�,nϷ\"��G"��=R�T���lA��0��ˑCQ�GF�Xż�gv�Fi*�S������pH�u�GI�,ە�v������t�M������]�[ �wk�óX��V�0��nb��x�(��9�\:V�m�Mry�V��\�:��P"�ԓB���-*Ls���#*�p5�LKј�ߺ5-�ӏ��~��?o/7Ϸ�E"��DTB�1DX�DX�m�UR�X�l"��UVa�Q��V*��V0EE�`�,���,Ţ�"�EX
"*���V1�0qh�J�X
�@E��1�������B�
�k	
��-�q��*�DV
�PF6�jڢ,QR1`��X,�Ub���FdD���k"�Eb��iR,PB��Q���QQ��+YQdUV��H"�ł�,TAAX
�DXDE�p��ElPPX[b�+0ыV"
��qk"�bȢł2)iTX�*�b)T����m%m���ȪE�1EX�EDRd��~���)2h���&L3�tϊm8{a�{�ĜPV�wWB�CS�m���q�WV��0�ev�7�4O_}_}�|��b���5���Y�߂�Lf���槠>ؓ�}�q~Qz�1�X��{֜��Ũf�Z6�<]n������/�������h��7�|�X�)y>�'C|e}�6�t_eY�h�to�:�[��sZ�gn���q�ݧ3��n{g)\��T�h��/�갘7��Y���&�ݖ��jx��P���>���G�f�˚*���=mv;[��b�4bL�fb�nΛ�'~�6�̛3�{݁��*��c����Gΰ�؄��u���;��~�lvΝ��R|���ދ>����0uӱA� ��]*�z5Blk��CޙTj;�s+�q�ַZ�*j��x��=���s���~
I���L�=]V|�t���vt��vy��^ד���u�M}su��vr��R��@�����Y~߳ahw�ŭ�{�Qǖ7�ץ�Kn*]���S�Q+��C�ㇵW܄�_`���hWi�W蠯o��]��_lJ�NX�ǑyA8���;J{k��2ѽ�|��X�Ԥ��Bƚ4t�gI�Eo�Z�1�U�Z��R�Х5�s{��U>�,�ះ�}��H��rd��G;��op��E6!<�Q�]V�e�scN�w�m��Z���H]����#ϡ���_95L��yU,p�^����v֬�sCy�vQ�Z�>��7��r-���;/;+�{�FŻ��}�X. |�.������S��T�e�?Wz���v�i_�^�l��.k`�Vr��/��!���(�����^���5�-��]+t��Ķ{��r�P>)j�"��Օ�qx�_o=�w���蒇�$~�q{w��Gst�Ӯ|ە��{�~ִ����;��Ib�uچ{��-�"p^em6�{�	����>�lq��I�����zv�Qho��ɚ��>Ƽ��.�ڨ�>�u��q�@��{݂�*�z�l�Yǒ��ܤ�'�ٰ=ү�^'� SD��)��oj����OS-n��ײ�i��ؼU�l���'��)3/T�ǍJy=��]�j�d�m�]&��*ղj�Zj�+o܆��Բ���MB���yY'|
-��^�E�
�n���C�VA}/�7;/��3�.�Kێ�`s;.�Z\�!�0>��xri�;?}UU��ݏdg�&.�!�
m�u�{��t�{�o�	3�.�N�-����^}�Y$��-=������G;��\~Ν�s'U�i}���'�mwr��x�F��R��ި2�� ��S����]7ʳ�a�ҽ7evq��j�����;�L��]z�W1�Q����ݘ����mm�hMVrwmsΓ^KY��p9)���< �e�>6����ג�R5o���{y4��u��bdx!���MS.v�����I^���T]Y��֭�����D���W�Kc\A�,S�w���'OA'^��=�lͧ^7�3ޕ������P��(	�����O�:O{��0~���s�\A��m\(��>ֳ�$��54���(��il.�ZЬ����S��[��Vk�s��b| �rays
U��;"	�)l���>ъ1�%Ǩx��%�j��ꄍ��M�H1�w�WL�w����Ϟ��^E{w]�N�A�:F�]�\���o��:���2�(6!�"��/. $�q�CmGֳ˕��o�0��]Qdۇ/�0^c�8'�������]ޞ�_{�7י�-i��VE[�c���w�G��}�n�y��+s�B����},<Q���ް��3�@�8�q{#�pz8�}�K~�A��>��e0W{�L��������b����r�
-�s_|K�����nz �!.�2�<Pd߭c�zʣ�m&/����>bu,��9��c���#�;��v�fț@�ۯT���'Z�|���$���X�j,��}��&��=�B=�ǵ9}m���:��għ�j���Ƹ��0:}��&6�
q�s������<��>q�&Vؘ*�|%g�:{}��K�[	MJT��O�cL]}L�~~�sd�Q���x�"W��9��T�[k���
�෋A���<�KY��[�9,"o[�>�)��5�s���J�:�a��[�ͅ��Ԁ�s�����{YCQɦ��ۊ�'��� ��G�F�j�ͮ��9��
"k%] 2d�w��������3޽���1��l&J�u�����K��[[ǳ:�i�P�E���$�.P�%3o�����#5��&t��(oK\2cS�/�VU���k�ڱR���>
��w%2;�û��0K�5T@�]��^�?-^��H{a���9eJ�B�cy��݇:6=��5o���x�\e��N��kFP�=ג��}�t�}ޑ�V<��8��Xj���}��^�!ӽ��kp)y�	�g�?K���P{s�C����C���ʬ85<t0er�3��RC�m�}��.Y돂�Lf��G)�R��h������J�o�)N��z���[}��J�9���}���c�W� \Y�����^�:M~�|����f��H_��n�\Ceu�\����J�}�Ûy����}��El	=�>��U$ӷ3�����8
!���侻~��D���ɇAǾ���6�C�������qd�b��8���׺4)�,yJ����{>���q���u�1}�b:�A�P���JnYG+sۈZ�VWئr�0�hɛ�c=�.���*宨8���ͷ�N��ă�V��\D�-�|we��t�17	��r������D<�:�pqv�+��f��quǰd@8�Dz�Ҧnk.ǓDU��S�����5�}���qw��q�q_�9�������$��f�9Ox�O�9w�d����R�S_&*d���iK�V�ǾZ��\�<X&I�p^O
�7~�x�w����Οw��++��覲�)x���;��f�<����wH�P�ݑw��IgN�\��/���]V�־��l/>[]+�v]nd���`M�k%u�^��9/�\�S�*��s���-�i��k�Yn��i�Y�����N�x6i�7��$��?Rb����Įʞ�z��"a�x�5a�8SB�:�:+i�˕�lh�8RX��Nz������1�p�:{��Um)�J����`��oti޾\�:vV��PC����}���S����Ϸ��s�K+C���9;�m�n�{��57�:��V��_��Fϧ*�4��T�T�����kni�k������粬���~����5���שC��{�bTSkƚׂx*���߲�f�^�nP5�9F������8ǂ��.�e�	"x�c�Xn����^L}	���º7��Mܮ��+�7ZS�(;��hvŎ��U�$u͙���l.�n:��瓆��Ep%K�P��+X��km8�LM�$��Ri�!�\�@�9��ձ�=�<��<ǳ��  ]㽱���մ�P�n�G�"�/{i���\��v[�T��V�CJ��[�Ng!�Pf�o�z=�}���=��_[���B����¯�~~��),g�o�a'q����3�WY�L�g��PX��κe��8z����|+x�v$:�B�- �x�`�ڷnl�뵱�y�J�ጒe=
*��5*�|��IG&م�&
qs/Dt��2y���K��ً����|��'�N]��a2���6��LT�ڐ��;�M>�e�D'��+���Y~�F�l�1�K2�c��?�w�@��:�Ϭ_SYmX�i��2�UY*����ܷS�-x���sX��l�3՞�1S�"(X��Y<�g�,tC���ۓE]9͍y�����i�񚇟���Ǚ�2Z�/�O��T�<,�K �H4��eX)&�Q�S�;0y����O�!��k<C�6��˘xEr��*	�f�{�4�Co���6.kǄ�e�ЖW�6�7J�|�S9�:0���v=[�H��Bq}\����T0�5�/%\w[�19�I���=����.���`v����!{�������}7*y.QQf3*��}E�݇/[H�fgFgXü(,1������۩K�|F�V��u�Гo��1d�"S�\�lwx��Nu.;��W�U�N��{�&N���Z$�=���H��3p��1���W��r$�a�H��{:���9���ػ��P�_�w^+�$&w��u��0��5^qpφ�~37���v&��,�F��Q�{���|xj G�`R���u�QhB�ԬLx�{i3KO�m��=��1�&7�l�O	�����s=Bå=���Wn���V�/k���g��.�iG�ʮ۷�xXx�T�#�^!y�_���}���ϡ��g�bd��?ܥ�����h���Z�7�mI+us�����`ηK�a(+<�A��p幘7��=>��v�=c�m����������ɼ(�8����>2�;�},�W!�� U�؞�s=Sh9��ܹ�!Ks�y��w��(�V� �Vz!�x�(P�ɯYf���lU��#��\���a��]�:"���y=E+�[����_30�Y�H�+-�*��7�tJG���w.�N���Q���J�~!�ܮ2>ŧZɖk�H�R.�
_�%Uf�b��ǣ�V,��-�i��8��=��-��k]w<��Q�31&����Vj'�m��n������ʰ��өy��&�ێS��>�&�����v7��Wz��C����+�V���n��s��oY�1�j��M{\xP
��0�]i��꯾�'�5�ځ�ߔ���>���K�l�'E�/��I^�F��,���YظZ���[k8X������|]�:��Ͱ����g��3+��{V�h�4^��ڛld~�o���K>%w��"�-�d5��53١�q�9sưW	� �s�l�����;i�$cں�������f@�]׬¨$\>����W]��z���"��_T�M˗`*�Gr�@�爒5��%����L��"W�X~���޼��ȩrt��g�D�
|@��]�J���HW��vQ�7V_o�JB6���LU���ݣ���v��c0���ޘ,��Q��8X��ĩ`o @a���7nQ<�۫@շ<�08�v�o�z��{�N���E7.��r�����&4��hw� $��w�s1j@�蓩r��x/�s�K4�xiL�3����Vק�i��>����}Ri�y=�{�os�M�dh�\��V&���m���Sσ��'��x����y�P=�uՐ��p �Ag�>�-m�off�JH[�%&+U�m���[W`yk5��.4!�zR�E�;�"�L�"�r&T��Ao�c��갦��}���H���o�3Nw7goA��5��(Q7s��9�gS]r��;�(�r���b�?}_}�{؟�����EX���1�����	��CN���;A/��⭊����V�p�{����wˌ��c�u��q{�mt�לy��Y��#F6-�ϑ�i�|�KU�*��_&���}7���a1��!�nS-�F�����!�!�;c�b�<�&ߤ�]uTՈ��v�=�a!P��cPq��;�f���A^�p">QL�8s�h_c�1¥��9��3#���|D��I��V]�E[`��י�w�!Ϧ����&xmA@6�T�����h����A���<�c�f�B�T��u7U1�OM�km}L��W�S��j���l��t��<���^��`�����K��EXx�I���u�d����ŕ�^n�[EJ�#�6/g���1�)�	=3:���a�X(6E
k��PzS��k���v��=J��0yOo��4Ԩ�R{��z�x(`�D˃z���A� Q�vP$>3=<��Ʒ��[���3�Y��<�v;�s��t�����
LV8.WX��LJ�<�jp�m�&����e�Bv�C�&��^�c�N�[s,����YH��L�x0�~�1�؝�tWF��3w��Q�������p�[�ǂ���y ���YI��8M!oI{�V�]|Eu*K$ǛzP�郄�om�/k�yh�Ri��*uo#`��ɦA��(�k�\dVސX�mP@W=�������ǂ��U���`��8ɰOgNK�6��#�vZS�L"{8��܌h[CAwz�����e�c��Lfnfت�p�/�1��7WCV�b[�v08�ɬйH3�Wp_cͳ��[»�&�VU�kQ�eө	؂[�);Aodc��]��	��CI�U�T�\����
|��3r+q+Z�z��W7rՏX����WM�^dO,T�����*8�]Z�6�	]a}�_>�����0	;9'e��B�d�X��e���"����wQ1fq\�o9)�����<�3�!����غfgY�n���G~��A}�QR�u��_@^�v>s+�I��Ź�s��L����:����x�]L��9r�Kr��O�T�h��K�a Q
���I�Cz�I�n���݄>�촁�������9�凩!���Ϻ��7�3/��O<X��-qC�]�U
���\cXq�~��7��]�߶hc�.c\Q��3Lt1�z��ӈ:ü�H�.�Y�/�&��bC2Vy��9Vuj��7x�C�S�:���`�`�ݴ�3��^:Lv��pf<�t:���v�J��0��~��tSr����4�MN[�7%
PfQk;0�����V�u4p�0fQ��S]��wB��]�>7aY��d�� +b��Tiu�X�@ksr��]�m��s�:�U��"�hO.����5�l�����Q��^s޺�����]��RS��x�J���.�U�z]
e2F1:����Ww��lV��sTn��}���r����Ӓ�	23`���B:[���(g]�`�b��w[�ΰz��}�������#�xP�k���(	XX�vӳA��w�ؙt/����Ql��`�ݼS/orT-���dcTZ��L]V�U���O�]�ɚ��oR�'gp?@u�v�HL�P*�<��.pժ�T�Y�O��J���BC7&�k6�6��s
�t�]zn�Ч;�^�Le1U��6X���&���Jl�h��WAhkɵ�{|��u��A�2���6&�\�q"�n�[4�ɭ {9�.�f�WQ�Ft�PE�0�Ȟ�/3���*�����!���yK�Z<evJ�|v]4���O���ᇸ����d̸�C��'K�)WKJ<���clX�q��r���N�V��f�]�u>Ыyގ��8�o"�����jhw�)��!���^Tۼvܺ37[
h-��c]]�i#�+4Ǩ�:��.�0�1էqމ��)�m-i�׺բ�s������x�߳�5�,EPX+l��+E��T�1��)U
�+jA�������V[PX�YEb1b�QEU�Q�*F2"DAT����[jEEQ���
�#l�U-�Z�U(��b�mDQ��F
#Z����*TZ�*Q��F**������EL5Y*�V�"(�e�V�AE���T���[ke���6�VѴ"�*,)R����
��Ńl+bJ �%J��ڃj��YJ��0[++`�Q[eQ�KT�b6�V[EՖ�5hPQR,+QK[X��dQT���ЩTeH�iR��T��b������VQ*Q�H-TR��+Q�e�D�F@
"����A9I�-Z���ނ/z��Γ��ɶ��n���r��wti������]N�JXqԂ�+dD�n�%������}�%rk�T�~�z�+�����9S��|�%�(b�.��eV��}x{=�ǧN��Nk-\=�QXݧ�J^(G������0r��I��{���[R�FWQy�cS��ٯœ$��.R,��=� ]��TֱH]o{�3^�SjED�?m�H�Sù���� +*?c�o���;5W�"3Ǒ�d^u��ƌg�˪%eep,^�`>�ԧ}�6�Of������+�I_���E���:%�ϕY�1�I����{�*۝Y��3�-�+ay��L���S���F��
!��*��Z���_.A�������[��~�� �R��k�]LCK9n���r��O��8�v�Px����Q�dȒv�ɇS�gJ'��IA�ɀb0�-����0Dj/����hex�g�M�m�X�2�#P���'İ8��(7Y3���BG���i�l�&wV�t������ɉ3	�H6�'U�!X�����'� N�	�{��:�ݾ�0|7��Y��MP�)��d=S�����2��L����C�\d󱻡2��ef�����x�a��jصO=�;^��v�!c����k����岳8�vd�8`�-g^��WF�ev�{�:ͥ�(3h�Dj@��i������;$�Y]���K�� ��c*M=om��Ú={�+�~�=Yvze����,V�b���2Ŏ��qשt��w������7��C�w�v��7`�Fs���d򪔦Uк�@���OiƟ�L��MW��������`��k<C�E��0���	�0xx
�bo-QV�>�Ƒ��&]���^��9)��s:éJL��Hm`r�y��ٴ�-�o.y��}ִ:؉*��f|��R%F�Z2�j���������efϪ��)��<�TyZ��_��vZ�v�!�Tg���ue1�9��߇q���W���f�{ܵG|֫�Ճ�� G-�WCU�r��/ja{��!���͎�G��g�59�Q#�����ӛ�5OC`������Z�� ����N���I���yI�̍��WG� ���,j���2��{'��]�Z�ru��P�T���S��OѾ�4O]�9�]��r[�(+<�A�R�=��p1�z<�q�:H'^�x�{ϯ#��D�t�����0v����yP=���%[��a��v�^��N��
o9x6D��U���[��e�*�tT{2��l����љ�A�bQ�a�s�9|��>�9FAQ2w�\�ihx��Ȋ�1�ylx�W���W�V���׳5�}
��?T>-2`�1y`.�0ڹc�%U/����n,��Pں�ۮ{g���վ[�0qX�����Ch_g�̻ڈe�V�nX��Bs1�OA^
;�?FLF��.|j*=�:�_3��Y<k�t]1��5���
�b����/{7���,�Z��#��h!����q���ؑ���
�N�u�]�7/`��Ӈ�{=�a��`�rC�E�+o���N�B�o`Tѝ��[��M�ϦrKm���-���l��\��j
#*�"SGl���2i�.��^��aI�=��O\��$9�6/�V �ݘu�����T̲*Ƕ�%�Q��~7�(v��nx\R��}/V
p�5����Cg`��>��PV߸�#ƅs����NU��� Z�������E��t����1��Γ��=c�$��	�*T�]L��	5s�Qv�r��S�\/����>HnG��9r�Ed<�p@�/�/H�m��Le/t��<��}��ڋP[�4g�v���arלL�,Ÿ��k6��?)y5����l�X��t��`KV�>_	Xz��z�n�I|���u�Rۜ�U�0ٕ;�N�m
�:�.�f��Z�N�l]5&Weέ�dZ�j��.����U~+���!)~��Q���ۡ�7�(y�J�,RzNtUZ�Ut/M";UM��%E��a��>h[����Q����l�C����k�i85��_y�u)S��[W3;�gZ,��K��A9�M�+Eh���y��u�ԥG��AY��A�C}�y��<7L�a�ygMsZ����,{����JÄׇ�iZ0y�����j�~�[6��9ܽ�\�<�qu�<p�}��4r⪦�Ӛt���zP�7�u	J�뙹�*��Aޜ�`���[������8�}{������&�"���/�ބ��޽�o�����
"�ŵ��X����8��{i^xB?r���6��BGbrh5��|��)�o��,�!G�����s]�g�v:��4�������z�&��&[y(��|��z�0��'���$�ۻ�Wؐ>F��],C5�¨A����J��b�����i��@�j��f�vi���}`��T����Az��T�z��̡��RǨ�����[OL�g<�&�vD�[��ͽ?2�`�'=�8VS�f�%b��[&��s�3��Af����g��k-�p/�q���D��V����g��7{!7�Db�)gVֶ��u��icsZZ�AYSN�ӲbrMkgT=Q:���O��ܓyY��΃�_W"���DU��e z�2��l���
aO/k�Wl=�>PB:A5�=e������C�70eP��ҡGP�NR;��o�8i��@�����m�y�̨>n鐶4#��c7��2�+��d��)U �z�xG���z����{�e(�|Wޜ�>�t�`��]HT!��'Y��p�,J�1*���o"#�[�����{$	}b�z}����f�\�Δ�uܾ����Y�r�y�mI�9�w���0�1�SH��
�|)���R���g�F��>s�v�Ք/<���Q㕀�"�TyR��T��{���/�}>�W��wt���~��z��Pu.��<�{Gl�S��:�\ּj� �s٬�9|��܄ܳ]	��c����I�v�L}���G�f1(��x���`��l������ �E���h��<6�'��p�3�m���c|z�q���XP%g�հ��q:��Gմ�zsѩC|U�
�ԭ�t7�Z�!�xbO�+1�!X��̸���4]\�}��_fzZ����xpjX�D<o�>)�.��T�t��އ��X[�� �DM��^�W�"�Z��M.�!���[S4�v��7�ár�/�K�Tt�*��͒��KK�<ظE	��T5������\�a�K薀>�I�]:���0���p幐x��N���|����Ν��ev�V+��e_��\K�Z=>~`/�� �h��ev#�*q[����'���ڧT�;�!�"���.�i�O�t���f�S���Ԅ�UEu4ӞJ�iW��㨹{g���m�^U�`�а:�
��*����v�'a�w��[E�<�:퐍>P��%����z�*����nW/x�>�%}�U��`���������Zb�aVr�o�����ԧ��}�k�ƊUR'�[=23��n1�T�	��Ӎ��Щ����p�.5̀�Q������T}&~�x���b:����e��곪��9������ј	�Q$�����{Y�Z�ϼ���E|!Hm^�T�эN{��K3=�vN�۬< m�O\�&Y&�Y��/�Z����/�Z�r�oEd�/,�zV��ذvǞ��'*4���P�H9u��U׶�����>:&g�����&_��}�gfI��4�|��oQ���y̺�C�"�M�i͘�:m���!O/#�G�{�-�&1�醕���'۲��9��v�f���-���QU6�;�'�K� �+��@��KMv�A�"�:=u���.m����
��^vJ��o���V������C�y̰r�� p�������yQzψ{�ڊ��D��ygkݑ�v��=դL؆Cz|��]z��i8��
�^����Ǘ������v����j=���y��m�*����L��H:��ac�qC���A�L���S��[]@��
ǗQ�ms��r��u����S.�Ɣ�����}nf��#���m
�e�Oˤ1s���ӱ��Avl�㔹`.�0�^���V�b������q��):j�}6��������p�ϖ4=�^#
��/���a;Srث\-�i݃ɔ�kwqw����{0�����`��M�[��,�>�^������X��k<&,�^��)��kiqn9�h�~�p� ����L��£�\SB�>��!K�� �M*��_����xǚ����C4�̯*��j��_{����kA�|���sp�7���F���b�S_64��B���+I�����Yu�]6�s�a�����e��"4eاѧ��mQ{���|��h0�L����=���R�ue5е3�iץ+��u^K�������	m�JN��'�x�rΨ�U��/�� �8�u< ����}ATy�8\�ԻsgT�2y�2{~T��O�;vÂ� v���Ė��'��ҙ�]�/�#�U�π�{�y=��>���}r�+K0�v�3����α�n{�V��"��{�{$O�'�nkNvz�+L�}�*ɗ0��ڳ\ɦO|�xs�߆����"�E���D�I{���[���n�Σ�R���w��u��r�&�$��W�L�Ew+o�B+����w����W[D:|k���"CK�@�*��0Vۻ�|���3��.XhR{7i���8歮VT~d/�{s���ۡ�7�+�%+C�ޓ�tUZ�Ut.���5����b���]#`��|
�R9�^��S���rǉ�5��C�c���Zox`��pֻ\�~r�X=L��E��mס�e�C=������A[P��C{ʟ�ƴ����3�ſTY�R��KU�c��o�!�k��%�#��������!@	w��xS薙�Gi�;�U�0V�q�N�9�C�T�:ti7��w�.������M�|*a�#�zmf�]`��u�7���̨��!η�r�@����v��<{�\8��y��xg�(�V��w�O��֍b4g�������0��]ɾ�O'v�dDRT���Qluշ�t�	�]h�	�U��X���8f5��䬁:��N�:�E`ms6�`��|���e����G�Wxex4�p�Yr}۵yT-h1���q}-gB�[�Z?VR���j���n���:�ڜey�C�4�����!ö8=�f���ܜ�G;aF�.� ��uÑd���;�(9������]j�X��K"��lfN�Ǔ�BWx^�2�"�ME�݊���
�f��C&��G�V��� 'k��TǼ�h���Uc]٬޳L!G�ÀX.�ƕ.��gǼ�m�����C�9��Oo�ز��(��< ���≃(�a�,N��f��!x+9��c�n+��7!�WA�Z�ɏ�<������C�70UФ�
���rʅ
�y-ެ1)��.sޕy��y.��>�dt�<ܼ����z��ưz?��*R�اƕքF�̗^��2��=��qC���8�)�x.�^B�IӀ���ĭ������9���{�IҒ��%n�"�Y!yz�Hx朧��+0oLJ�����Ы�������/XX]����|E�Lc*��=��:��S X®(�.>�Zuvƺ��Zr�r�h"�g�ް,�M9���i-��%fdCp��M����œl�]�(�a�x!�.	�@����=yE��ޱe;C������)�旯����!���S�5yڛc]�����4���L����[�+hj���GxΓ���ܹM��U�"�;�T�RO��wלׄ��w�����]p��x�w ���;������5К^(��a��V\yhenT���?��u~ە�1ؽ_��Um=������LA�ہT��<����,n'%d)'�g���YR�Gk�k��PUC�Y�7��[Sׅ8^�ѩC|�*�����螗���:5������x.��n�����+�f�q�-�p�n)XD�}(H�{�'�s[��كu��SɇK��Gǥ%��-���W Kl���>��b�,l�MO'��vk�wcj�Z��b4��4�=����͠�]�]�H�sb��{�;g�S~�i���XŰ{e�g�����X�V �v�'<|N�.#6ф6��'�h!ߞ��*{뤽6��)o��3՞�1X�"���b�����^ꭧm��캺՞� ǯ'6����p��ݭ��������O��<�+�J�o�$������sp��.�6KM�z�l�S%
Z�z�|����?>�t{܎��B(�"VE��8�� ��;ߌ���m� ��E��X`����:d�o���~ޡ�X:����>Z�9S��X�ˋ�)�
�_�X/7z�ب-�i[	G�z�eh�S�a��]q�M�a���D]ss
Z�T�K���;�ǥ�&��(���r���_uY�:1;q Q�v���on��d���e]ome<o��$�q��^��x^U���AQ�;:��&��ːAmsάt6�c4I�{�m��[���Xnݶ�F4��F46�_�qá.ǧk�i�����"� ���v�8C�ʕ������p�)|���"v�6@�0-��Q�ł���E�r,<��s�l]���̶��Uۿn�x)��r}7q���M�\t �Θ���t`UvD±����5&-���Ü.ې�f��(m��������4P V쥛Z��b�ϲs��,*��B8$H̊GK��MKo0�ɡq}	8K�o�(���P��'��]��ɛ������q\��0����"�5��Z۫�R
K�2���-�ZK�y�3�/�Ep���en�ڴ_S����2�^�xҤ�z���
��$u�Q��������m�R�~i�ns���K&q�][��_=�f(0)3/��{Z���&�T�n����du�&�1��4���$O5@.c�n��̚�2Lg����9���D4U����4�Tn�v9:�[7�!�5�q�R,+��`G���P|Hmb��t:�N :�t�<�!����۩ ��ƥ�w׺o��w���J��u��-o9l�{w��P[��n�'� 2��n�4*�y�ΚH�߳o����;�oP%��Mc蒧�.pG�Q�_q�}**z��A�d�_Q	�GCdC[w��Y��Ԇq���%��6�'c�t�)v]����,�;qiţ�u��]����{��[F@�m�Î9�Sh�Hi(eoqK�7��
���s�9�j�ܮ��LW٭��tr��flW�s���/у��҅IW)j� `!@X:���s�MGVO��DA�V>/P����hB_wK$In7ҒŹ��;I:FIiu�[��ٟ\#%�����T|�Z��nokS'�������n�з.�e�`t�(y>Q�ͻ�4�4!t�A��r5�^��v�bc����#]p	(v�w�E�	�L��}>�G�Q9158IN���`�kd�d*�`�W�s`K��"ɠ��]+N`���%vZ�S�wP˔���Gx�܅�Ad?<,��oD�3W/z����e���Pw�IȋTT�Ln�@������l�l�KgCJ�г+t,&�np�'I��*�+L���r��RhY�뎜%l�]�\�(�`Q�iFoK�vl:�S�)Q�f�gX��7N�ǣO̶k�%�i���w����+e���pY/��b�ל�
0/߾��s?gH�h�J�m�T�(��,U
� Ѳ���R�6��*,RR��
m�)-����+V�H�i(�Ģ�U*��!PF,%�U�Pi`V�PY[J��b%ZZF�e�*�X[UB�+b�X�C0X6��� ���Ki*)J*��Ĭ���Deh�YD�QEmP��"�AJ�h[`�TjQ��FKd*��ږ��lU�V��Z�Q��4�b��P*�b��VT��-(�
"�"#(�[X������*,R�dm��Q��R��kP��G*�+
���R��U�
��ҡZ�dTh������Z�E*�mR�T����X��UQm��%j�Z
�m�V"2،R�`�`�*�R�G���QX�`6�T�Z1�b��J��b"��kh6�j(T
�5������������P��ͥ�L�
�R�3��7}1�L��lSd[�+ʘ�i=v�"����'G�3	-������oҌ����� �B�on��^�\(<>g�`�0k���!�N|��=p`Uٯ���?�Y'��vN�`a��=��-;,�~�|)�l>��X�4�
���3Lj�"���K�t������ؚxO\�&Y&�Y��/�Y!�Fx��s0=��]����y���v�n�����g�˪) �׊y�\~�E�ʿhUY얚ݮ����c���y��x���Sฦ}�e���8X�����k��O|��j�@��&l��ztɹ�O��A���!g�f�����s�@�����x�'�g�[���A�;���5Oz0�\���x/%xd��9��7$��l=W����_��]��wt��l�O��*I�������Ig)/%�/�䠬w� �H8K�O{|��u�{�zc]Mm��)������+�x��@eHr��1����k�Ī�4�nR�x2�o�oTL�ޥ-���N'�Ї�_�e�͟�Q�t���:��q��g0r�1����M ��r�Ɗw�ӺfZ[�-V���Z������f�x�Z�a�{�;��9B�{(w��$��~ !����ܙ#\5��U�wVn쥘1 
<��e>!��x��oD+�ؙ�*@&�����:�]�emwd{�b��v<�3�v~�߮9�'��rm��^��e�@�:B�a��Od�����U龧m�,b�-g���upNߪ/&�p���;�Uq�,�/�F��u��v�����s�b������КPM!�������ذ���X=S��oi�a�m$�|��9�\Q��?���`]oYdP�=F�;�
����!��u��ʞ��V�]X�2=36�O5��v�����o��Y�iل��g�����R�S�pk7K}�R�xm:-�t�n�J�p���pGsU�.a�<,4#V9٦J�S˸j� �m������G���i{
�ƗF}3�ڇ1��`��1˔�,D�E��@������F�n��q��$��K�QZ��k�	�'�L���2��h�Q���ئ1x���n.
a7;��{�Js�l����v��~��:v�f}�0Y�R�
R��y����I�{:�-ȏD�K)��_�Z�ׅ�\\K�7ڶ��N}�
��[��F��	˩�ʛ�>8m������|t�itN ���/������2r��-��SZ���!�K�8�c���+"]r��4��{[ړر�:��b�d���[]-
7�C����e�m�wQv���x[����:��b4� �9I4�"��~��Ʋ��2��>?^@�f��Y�JT`g%PVl�P������J�r�<Cp�:��eٖe��Zo̭�/׶C����,�E�D�+j٨� �,�0���oM������D�{QТ��=�&'�Xߐ@o�������`���i�Q*~�.E�7��*�1�����e`��x��ƣ�ѓ��1�Q^>i�D=vt�þ���ݾ��\����*Ɗ�ru��/Pu��
�̭�~�h;�=�JE�􌌓�go��ބ1�6��!�X)��X��0���3>��JB�ە�24q�]wx����m�xwM�HL��&�
]�L��]�ؐ>��3���
�3�U/~S9����bK&���QU�M#W�f�_Q�p�]Lwu�FH�p���/}����o��m8O���ߪn1�5����4/�&���b�F.��!��ga�G�a��k�hz��t���m�7�Y�x���L�u�lR�[��
��B�3�b���B�8l��b�<+1ȡ��<�;����`w��q)���L8,�P-uv�tv̮C���ҙ�]���0��l�H��2�gF�=�Y�4t&�-�fNáNヲv�����.#�WJ��H7S*w)���r�6}�o���t�C�;�<���a���l��n��'fV}6"�ϺD5��g���\k�+p�
~#y�Vq��1��-�P�r +ԝ��j3�R��r����L�}��R^B�IӀ��-����U����ݸ��E'�c�.�	]�Ȫ�$A�/�%��4�{ܥf�ɐ��D9�v���y�}X�Tx�_�����n��w�y`C�@�/�H5Y���.�,vQѬ�lG/):��������u��곴X0F�
N^q�o��]d^�gר�N�*��Ǐ�0Ov/f!Ҽ�yYjj�=\�K#i]p�\��w ���;N_#�ק�l�񔌳!;<��2�U����.s�mb�HOӔ �0{7�	J��ׁQ�{)+>��1q��d>���t 7���i�j`z;�f!��r(bBք�V
��f�u;�ja��z㲽7�B����s~|��9V#��������x �F�Q���1a���8r�̀n/Z%�&7*j؆�/x��ekV�T����^���'G��~`*z� m�;�<hN��X��L�29�f�	�Y\����1W���N �K�Pn][g�i��L���zD�����uv�I����/����Im��GBJkv��ћ˝��D���&9t!㣹S��LLD�E��øç��r�eX��V�k�N���F̭<�OPs[Q�G�1YWt8����� ��왁� ���{*�"��b]���^Pl��s��ؽ��L�z!|%�]�lV��x�C;�㡒�W���M��y��/:�e�=R����C'Ӑ���x�<�ed#�ϦY�I ĖT��
쏵�	��ň�غ�?;�5=r������"���t��{��ik���y�en�c�o`= @*� xvO�*�3��J6�TΓ�KY�����=��;/5�ݍ��!oR�>���g��������B���?:հ���*g0u�]A��a~	\W�+kC�jq>�0S�PnӼ�#�>q	�`2�e�zO��}BлuV��g;�Z��r�|�K�7#\��v���d�Pp��t9���S�Yu]��l����G�_Լ�^&%��;��>��d%���U3ם���*q�r�L�s��(��, ����ʞ�-WV�����;t=�[s�><2�P-C��L��=�c7���ôuܡa��l�qݞ��[���=�i;=�r�s����u�����5g	[�
��*��3�WV�O��IVq�>�!���!\�|���]�䬝Ք)N)����{��b�|�`fA��&��Y�@{�z\� �j��Z��ӛ\���GC�	6-�m~��y�j	�m��c[���XO������ꦂ�9VbvOٞ�i���S&�U�8ܤ����z���˼�̓v�R��ts�%"��YH;N�������]��W�.R�@=]��J��2� (Y�[#�j\ZR��NS�!9U���y� �㢴^�8��g*�,�`*����3e	�Bٵ�fg�)��ޏ '�-�s=S~c��C����0w��T:����#�}sN��$X^�>�}7xО�D� ��Brj����'�ܛn�GW�Ͻ�Ϣzi�p*�>�����F�>���פ=ݛ�I�,��w��!����[�c�,�|��U�s�j���Z�x�b�\��OW'�0J;{@)i"��H<��O8+|]M��Js��*ɘ�g�.I:!��/��w'H"�Xb|�X��FP(A�� �OO>;s����vSX!��~���L��>��ݸ}��Ts�I[�����>%�v�2E:[��ÛoI��=v��D:x(���ח�r��͹�X==s��ڲ+;4�V�SX���T<����J�6g`Ѳ��`���쫄Z���m/l��h�X)$���m�ר3}�q�WFC^�T4,��-r�Z3i�2�E�B�Y����@�G3�$�ﵢ��Sotk�Ս�}�q-��9`�קy��+6��OiҜD�.��g�DK/mC6U���=�`��>�UTf3�b��
N��TG�`�r��,D!ۻ�pg]�:R����i�b��Nv���˴:}�5c~e?^������L�8�\�Z��	HT/)
�X�s}+����2��\:��!?vzn������$7BYb���&�ݭW�..��3z69=�45����w N�9�E/��n�Ͻ���W9YG���Uz�
�e�[�V�K��d@��@A�/|(�סy�k��ʫ�����ɯa��&6�ĸ]Y�m]���¥lU�ڦ2^��t��d��>�X�t�?Ki�V=>����U��c���ĵ�p-6=�es5��}"T7���Ͻ��FK�8'�^�t�g�%~��lg�V�xDg�]I����%�(d�
�^�!87��;c�|kc���z,�m��_4fřK֒<��&�w��\��|��CMBD4^����t��u���w�NWᦋ��΀o��3�ev��i�#�V�`��ff�PVŎG����a��N�e���49rFR�Hkip�����G�0��J��H�kG�&ѯj�����`�:N�Y�0=�;�P�WEh�R��k'^�ފ��4�|҅��w�]s��,�N��Z�(�,�x���+^��18��>!9[¦i��1ۑR}�5���I�3�
��j�g�8h��Z�x�@����%����ܛ�`�\(�y�Fҕ��ۅ�7힘ϝY�����R���ԃ����GHD�[@����beW�`~�7�W,9{�u��/91a�f���۟C5?z��ys>���_CT%��cO fu�-ڹ�$f��)S�߫*� �^[0n-!�{P��dp^^'�U���L��(S"k��������:Ro��r&Y��/���ٕ�M��2��\�_��m3s��`�G���9���;�>�|��;�t�s xJ ��e�������w!�t�g�&�$��S�2;��#~~�gx�ǳǱ�Dm{�`�^��	�
�
�Z<3�Jx�oԁ`�/���%��T�t������Χf�aT��b�Gt�*���߇Ba�j�T81o���]��m�XS���~��f�o]׸����d���b�)��֖�R���g�q�ͺw2��ވ��pM�F�����f�R<%f�z`^��C�u�g9���
�<����{�>�r��D�XC
U%�ʣ&���&���w�aT����^��;��xj���s�]�Xe��VVŒ�����xX�pUc$�ǁ|���P�FU�]�]��Ċ���"�+^NP�-ᕼ�ٳ{�9�۾�j�uc���֞W�y�Y�&��e�תB�U��Rt����=��|uj2��*W�8�Um`c�=[;+��tp�{"��Az��G���]*�ҭS�.�cN����$�`հ��n'S-��k�S����'��(�A����7�)c��Y��ެǦeܭ%d/��������_�pu:�S���E>���Ќ��}��YAxM�Y�p.9T���T��{G��s%���aw�ryd�*3����&
q==�:CY�L�������O;QZ9\�B21;:�7�L����oD�ֱu،]CfX���WK �B�3��lW�Q.��p��M�}�q���iu�J�7�YV`�����~3��,M8��"�(������?b�Wz*V�[�Ε����ЩB
��wOGE}e�i����R��6�����f̚|hp[c��J`�Y�[~m�����T� �>^��=B�k>5t��r(:�=�Ƀ\6����f܆�n�y�Q�z�O��;�{%e`�)	�f�t��ʻb���S�j��ϰґ
��^�o(T���\�4/�vs`�E[st�Zj`�U{�qj ��X��þ��{�5����B���5f�G�O��Ў�FB��H��pB	9�f
���mZ���]�u�[J�Kǉ��Y�[�mu��x�IY�7�x�v6����3�ul�R�ޏ->5=y��������rx\�&Y&��f����-�L#�ac���Z/�M�s6�}u�Tފ�O�)1X�����^-]��� uʿ�Y�[�	���%\};zҧ���/=���+��9��C\ʢ�u�_8-�R��y��7��zg��i�:9�v.q�@�5A��E{�Za=�c>�m����(kPQ��<5���Ĝ�R�z{)��6z��]�k���bvn�>kO��{�k�7)|�������0�j��i��^�o�^rϞ��y��\�~��<k20Nc�'!��fA^ܾ�~Vt��6�Su�Ϭb2���L���n��{ZϪ�+6Z蕏C,r*��������^O����~"U%�0��؅�Bw��z|!��Ol�޼G�P���>��vq3]��~�kvgh��}P��j<�\��fAX\^���}ltb�����\?a�`��P��ٞ�s^RR������䘮��L�`ʞ�v�	�6�`��>}W��왕�.����B����m�˾��DY9�@�j��#4"9�*53Dn�WAݳ�o&��IJ:ޞ�0I!6E#!�l>�P=�Yb�є��.
�im�MK���h��jq��\���`.�]c�9!9�(I�fŻٚ����Ĺ�)�(+?.o���R�V.̺:]��t��n�V��t�P2���J�ɬk*t����U`��6��ow�Ƴ39���u�Н2NJ��e^}�:R
6�������vd��c�� �z��iƠ�R���"�׺�y3�	[�i�Mb��WX�AY(#�Ǯ�����Ol���@1�tk�Tu�P�rq���ij�8Iݭ�ˀܜ�V	���#�+"8�g̤��	�KQ�-I0�}�k^V��<Ɍ-��[9�r�#�����f�7��$��	�CXU�t�J �b�3SƅW�h�P:S�V���U��s�f��9�1�V+�bn�(�M�W�������o�b4���+a]uJ�'��l@�3k�v"�;�jv�×�[m�k/�	Y�s�H�o��û1m�n��$mY�
�۰�v�a�ю3�9	�v5ɚ�!�Zt��f�V�mC}��,��!{o��_#E�5׺R�t�>d+��i�M؆*
�&��|³����m`ѻ:&i��z���J�+�2q�|�ʖ�� �}ڙ�5���:�S�0u:m��H��2n�k���r>ee'��´N k-�q4�EJ����Q���;Y��V��B`�ú@��E�yݥ�S}ʷ���.��R�X]l�����,Y$F�!P��1ewe%�*��ɫBN�P��ʔ+)�d=��r�U��bp�3қ(�	��[��$�u��
�X���-[%,�c�����0ڵ�v����q�$��,P��Iu[����ik���<�i������hQ�=n���d�i�-�:��j�O�o�=��Ȟ���p����&�feʻ=�"�YQ�Ag2����|d�J��1'Ko�d:�$��,a��������[�4Fܲ��}4�<��&Y�a,;���:�`߄}V��{�o�!<w��75����䝀�r*]��u�f�N����g-����Q�����hM�ŕ(��ͳD����M警-ۅT���cJZ�s}�u6�m��Lޣ�:j��wB��y�����*��Or��K��z�V��Y��������2H�(�d�jBnkBH� �J�N.��
�>���䵗�\�=G�9C�osQXO����z���a��M,�f�=�î�$���u,o>�h=��L��v���k�;t&���s�r���n��g��\!ͺ�5�����ݻ���(��^֭�j��u�oɭ��O�>1�T�O�v�r�����(�۶����b���U�,[#6<�`o-�5�)ˀ4�����Wm�L���+�2��ho鵺
Κ:>ĭ���-c����~ߨ}.����	
ʢV%�E"Z6�kF*�kX��TB�Ek
�e�bE%B�1E��-�R"�XU"�qA�б1D�h�m��,Ph�5(�U�PQd����TQ��L2�0�1F�Qb���+ ���6�e�+�KDV�R#QV��+[mA�,P��Z�Q"#FU����E[m-U������iJ��UDc"Z��T�EUb$J�Q�DEQE��m��(��Z��Xk+H�Ķ��V
��b�F6���!Rł��Z�U1J,TIZ�DTRҫiEehȌ�+-*[jUb�+PX�%QU+Y"���T��e��[��,[R�J5�DUA��0X1��\!�m��Qm�+[U�1cR�����H�Ե��`���U*6Q[*2*�Q,R"�m�V0jW���Ѣ"�E`���QEm���#}�k"h��s�Z�Q�٣Z�u�������`�"gT�f���#��Ms�$��Q] �*�Mu�8�i�=�ts�.~��-^���"z�D��W�$; �񓕾.��F����[f�pb�בҷ��=!oq�P�#�������0 )�QVi��c��]�/Oy����5������=��3��0�.�M!��Qꁫ"�s�	%�glB��Aʲut�I_Gt$��4º>wҪ�!���=�=�n_���0�X˘f������2P��j�b�2���������t8�
l�r,R���[�Q�L�B D_C�wS���/r���s�	Y'(A�}��\oF��zk��j�և�yA��Ci��zj�J���Z�	�CÎ��Kb�J�t���!���2CY�ݞ�[�C3�����ЖX�nW��1��q�e߽4�����u5����p�3닄��<{N�]��XO_�~s���N�N��F���eY�7��� 1����*�!x�^x'g�r�쨎A�}[c��t��\�u�o��E6v��\ny�d���C��V��sT�öC��yZ���������uB��>�m��$�D�Xn�����́ں*�iG�E��#ܼD���V��=������ Z����Nk0�@-��FW��n,����v��P�/�j��F��LA:0��u��P;��vrJ��&��&w���ې�\9�Y�0�L�/-��x��]���棢=]���	�W� Ӥ�U鐙6�q������̛�
^���U7�P��AX+�\'>�N�}nfV�4���G׿d�+���1eow\m��9����%Zg,�"�}b
�\��_ݔ��y�i���7uA����Z�w���ލ�N���FF�p/Ғ�|A��[9��P{ff�R�+��9f����$����ؙ��!u��=�4JP-	�.������H����X�ܯr'�4�vT�y��+�`�}���\�`�A�Ʀ�ҁ�4���U�b^o(����V��&ν���z%3A��s)i�Q��u�CS�)�����P�R�a�u�('���6V_����4��>��>��^=�+��ZC����K��8/��O�n��M�i ���J5^�K��B�c�r�"�Uul/+�`�,�\�֩/�е��(l��p�����ڙ'W�sz���� Q���Y���ٔ��ԎHv��̟o�)^�5�%�*79ܲc-�|k;ڂ��Ⱥd0��$�c�,���ͦ&0r�^]����qn�XFr���&q����h��Í��di�p���Ͻ�����e�4��d��7��->�.�cO[_t�bEN��>�st>ջ�rt��R�9\�_��f���^��"�[�xg�XxeX,�Rm��<ORu�,�y{�c��ɞw(�b�5�GK��A1)X�Ι�VxXc�L��<Y�+�V�fz�����{��c�u�z+%k�%����8�7[�4���N�l�}��KA�fn��b�3#����c��nv���4��Qs*��R���ߨ�>ӹ�<	Y��#�U��Q(=�9�=~���9��@aP���d>����b�Jp��ϣ���]��Y�����t��hl�б����o��^u��\)�%���~�L�97�ث��O����J�ƥ5�U�2
^�����!�j�!���=w�F�Q�AW��a�M1ܓ��5b;}'E	���Udd��������b��֩J�&��.��8.�`QUy	�9"��L���r�2s��wUSe��G�0��3���8����g3O*�'I����ts(+z���m��3=�aܥ>\�v��k'U�㞖ɱk��8B�>�K�ᵹ�Ǎ7�ki*�uzG�|0�V}��ݓ��/w-�6��U�͸1ba����E����c5K���3[�IwgiKa�3�J�]S�Z���S�&>����ʌ��n���W�w[�
?uK�X뢺1� �ǚ7��{�NR�+3bJk�A��v5a��˝d��=�r�'t�˲�����j�삶+!S��#��?h�4�q���vC�&�g1ݼɮWdP��U�L�`�c��ȺϚji�3T�p�������X�m���5������O�Z��2@�Xj�Õ^�r����ͫ���gm����#��l-9�=��]<.R�Vj�K,�v�u��_� �\+��%���#
�i��W3�d��
Ck�GF|��	�r�$��t�O�._P�/Lr�_�vg��=��T���ލS9X7��P�����c�T4R]x����Iu[W�Z7Z������HD�|�-�V�F˺c�=~ݸ;���<��+�s���d�R�� .̫�|�464ic�3���ݝƢ8�ꕍ�e֟
)�o	��/�zط3�,:���X]�>��3�b�����.��@��jڀ�X��Zs.�zz�#@�n`u���C���1Z��������e�q��A��d �{�#�[�r����`c�20Ng[O���o�9zL�l����͋.���SB��[:��M{A#^s#�Pe^�ě]�XcVbR)��Jmc�����7"�Tc/&��Ŋ-��2�iҖb��*����B�'�c2�Q,��\h�Y*J�w���)q.Vc�\`A%�2��ݬ��	[��a��`djWq���h����e�&Ǚ�\���u��SdV]������r��=~z< �]N�	�N'���z|'�`�^#��P,�S�G6;�k�VT�����V�p����'e�J�./T���c���0!WmQ�����6�/&M��|.�B��гc^%u,.�+�\�����ܮx�ĉ�o��jЭ�R򑭶��f��"F��ڶ*��?hs((��]�˳A���W��𥡃.fL�竛{�>	nz�J�[{r�u=�!���0�2�A�f���M/|_�9�N2��3�0S}aOs�a�e�fÁ���Y|��W�n�9`����j��]5|��!�~� t�O)�o�╬�W�����}=sU��6�V9٦Nn�U�O^'��c�)�zǲf0�]���l�}3��):�}��X&\�"{��<Х��p����D��J�O���ܽ�0�-�,�!�P�2�ʶ�|�g�����ɹ��y�i"�
׷���ظ�\�D�Ёb���ΰ�x ���/�O�z�fn��t<�Dv�f1�ʚ�V����4A۽׽t
:��`p|���.o
<��6Y��_f	����ԐWgsV�f�;,�����u�B ~���\7�@ʛ���Y�u`JB�~��:�C3z`���Cb�E=Y2�l�2s�fŷ�+U�P��-�9��U]:C�aML������u�Ȳ�����T�}=nw�A�É�ka���JT��@�[Hn=�4�'^��W�	٤rDg.������4�;-dV��:�T�K�}��f�x���x@=fխY�c�\~�kט�@�?IU���rn�ض��_�jCO�z�}"T7<�tF}��>;����n1���Sz��o��O�\+O�Ɗ�m�6�B|/x�U��B�U��4���G�x����T+V�(��~��..<M�V-����H�U�(z"���p�L��+jq�=��� ���p���z�_���xq��BG��=w�g��!Eѥ�3	��a���hVb�ݾy����s�f�	��=�W�
�g��U(��G�!G�C�]�T���v�J�e:��d^:˜5��
0s	�/�kˡ�
��s9:�:�UcW�#��i�G�¾��b'������3VoK��M�Q�Z��{�� ��q(_ �����kQ�t�(��z�bݩ��Ү��şC7-S�l�M�\�NY�VT��%�0��}�w����
ju:�	��ǁ��XjZ$�Fku�5��8�����tC3 ��5]�sg9f�r���z�%[�$'��_��z!�ԧ�e,�b�>ÿ& ��L�@;����ѵ�����;�r���膌�l��q���r�{�����g+�dKk8O'�үvⱷ�������^�eСG�!l�$+~�n�g)fV}6"�Α~�=]�n`�ۃ7�֯���ġ�{��j��Ԫ��1� ~�e�\+=Y��ԍ�\V��I�C7�����7j'�R�_��)>>U�+�1*���f��˱��y0A0?&�,��9�nT���d~wu�'Ӟ%Ir�Rf1X��<08�������ό��T2�T�����t��Yi>�O���QG�p�h�ڼ�yԩ}ܫh:�SN�Xk3�a�}�[#j�ܽ�8'��ݻ"���W��'��v�f�����G>אYT��;J_#�x���oVo$L#���{�iz�� �XvT�F3Hu�
�ܳ�V�f�64uk��U���-�����˔}9TC�;�9n�M��C�X�b���&++�a�4��Mv{�քO�t
�;us�)j�+���]����]�^qG�b>gV�y�x��� �Oշ�9{&�r�ȼ�"�8�pd�:�����:�P�+9B�0+�e�+�f8��$[1"1��{p�7�,�H�nMw�[I�ұ6H��'gv�ҭ}G��8�����W?<Ky[ZR^�,RE�A]r���6�&8�G��^K��T�{J��Z��j���j�~�cM�'Qn��_P�U��*�[���t���-R������f;�3%�^	�CW+q&�~jՌ�> J{dF�Y�>�#S��|WTad[!�����v�ݩ�K���7e�~M���Ͱ�X�.�$*�]M>�`L���i3���������%��]���Ɋ�(�O�a1�6��[��QM>3T��	���^��y9ef��INF��rt�z�L凿=ۡ�(���Ŏhb�];w<x�R��6�t�>̗����qwnz�Y�Pw�?��u�U7 �*xX�v@ ֚�p��5��)w9��7��\�v�dk,��O�/C��s�	����"��x��
�~�-��Ͱ���(����u��ϤT�g�a�C�,������=^s*#=F	���R�zi.���-{�3|ԥI��UϮغ¶�<�r�謔)�)�)1X����5��eL���Ӂ{n��^6�v�����J#i;H�q�Z�/�*���\��W�-�{�-�Ύ�s������� ��E^���a���E���4V�U���4��w^���Ѻ:��_�P.2�c��/�I��ދ����H5�����K9��pJG����$.^��u���.Ct���Vw�(�>�*������yA}�Q=��L|�k~ڭ��B`�#�&p���&ii�)��x����>�U����#q��g��\��lxr���zh��mxAkf'd�@�ii���L��k��ǩ�A�R��y���94��l��������|�2�l񞪻\}�ZJ%��q�{��S�Rmf��
���1��p�3�K��C#R��v�`���6Z�ly����Y;�h������bW� ��V��x� z�-��q`������{f������!9�}ۡM���b�>G��8`�.�5������s�@�~�"QxeZ�[y᜽\�����y���/����
e�#g�����2t1r��v�O!�(�рt]�)s޽Ӛ���b�>��T�!��C	B�Q s)D�g'���]O{�uyn��H�pm�^1c��ԣ�����O��v�������0 �4i4��F�R�{�
�I���|_���ٴe)�b�����h�x&�k��R���S���G��(�����G=W���t"rġ0ur��GC"`���>�9�[�L�LC�WF�V��b��7	���`9V��r���M�+k��,ث.�P�RV]o-�<X{�ό�fq�]:��5�xO\�����[�VE_;0�]FP'yV���zh7��~�,R��7J�~������g�,^����O\�g�.a�{��E
��ה�����r�ϗ,��x��kv\S(_:�n߁��g>��*���2�<+>�r�Ds�������!샺��7�D�y��r�Bm��Vj4�D<�[�,Hp@�Cx�	{���^1������Wy��@K��ʫ�*����<��n���0Y4���ķY�dg�f��P�בּ���a3��01�a��+���c;�i����R�^�k�J�n׏�������"G�pk���1Y�>q��g\��5��7��e&/����ԯ�ez<(z��0y��7t;C���s>�!�eez��Y]��i�;��tR��ջ�i��O�)yZ��돃�p?��[�{�
ުב�[���^�Ȭ(_<���o)��kby׆}������b��	HVp�LVW��N�u�W����}��� ��u�rWp����wj���*ݣNb��E+�y����8�����'�+apW=�R��֧ �aZ�2{���Z@ד�6�;���4*)<,>�� �at0f����X=S`ީk��W����O!�(�YY�m,nJ�mm��v��"ݓIK�d��g��MF��x��;�=�U�n<��Jj�b��PT�'5���h�A��󽦑�#�+���߭X�:��lUȥ��Rf����,�3Zb��d�T����Jө9�\�oD��c3�LwV��8h;ymv�U�j�mt뗸����A*���(ڲ�Q-�e�&Qt䪻���n�%��[Baɀ��'J
i�SL��Wly����3{���QL���ϻ!S�%��w�V��ۓA���V���9F�9�w4t���qw�S��M�6�q�5*ZF_�L�dZx˥$��wZ�ͅ�@�zB.���h����ּj��i����GU�)���n��i
x�n��:Ė�<ޜ�җfR�U�_Ap��՝L
�����]��ՀJIL�:�Sz�᾽�Z����^B.�s.�u]�ҕdT^)�iF�����ʮ�'�$��	STr�h�hI(�D���:�r|�p�ޑnD�p�,`	��]9�5�K.)�m �-��u��g�VTs>�U��G<v�o��f��m�����)
zY��i�fW ����ѝ��|�'['�{q/FU���}n�e{C��vp��s/��-��:v��2�jT��e��������H�X�7���d��ә�*�\o�L���֎�2.�:�l�zm�Lɐ�r�y�0�>�Fr�qk�N���� �8�#��!�jަGP����:>V�u���]�Ւf<SD��Ij��7	ը��L#�mL�R��N�T��fnˬ3S�����M@�S�ӈ"��[���a���z�qTQ���z�k�Î���X�uǯ;�=�,�m\58�8̮�7�}��X�G;�|߿.�ɏ�j�Ѳ=KrT�'�%��õy%��Slf,8A�;�J��w#b��q�Xo�'gh��X`8�ղݪќ1|o
�Ļz��Q���ԛݶ�u��YS�Jv.�v������a�or�R��LF�^�+����]W�d���%�)�$t(��/�F5�كk,DjV>v¨�_tQL�b��Of��l�'^����dnb|���U�,+y���5%e\ke�%��H�����9ݢe�N�cbz�X4]��/��k��w�G��!+Hj�n;�x�m�oL�ҵ����`aR�8��V�����ѹ��0��ʸ�J㨦�ܙ�P�\��BRܗX�l�C��6�Q�gl��G���p��[C��k6�w�T� ��(9�7.��_+={)q�3�!��[���R�6L�0U��]��/PDA5Ѱ�H{�]��ز�N}����ʂ�UV6�`�֨���
)m�����jZ��R#QFШ��U1e�⒣jX�+j�R�a�Z�-�(���TDX��V��TERڢ*����֕+cm�S���V
�m0��ŔQAV�PIYTAZZ(����+Db�ֶֶ�*��ZQDD�Q�1�+Tm�E��V��b#(أX*���B����(����(��I[b�ֵ�����-(��A��2Ҷ�Qb",��V�X�X�U(6�+A�ZX���Z�kB��""�j��*�EQD(QhDDEJ�*Ukm��j�*��@���(�V��,�U�� �Z�V��X��[l��aZYj*(Ѭ�V�j(�R���*�+m��,EQcX���UV ����*�(Ң�T��j���(�F!m-�"��DX�(��[X��*�؁JР �#@�5�b�u1��Ę�	Ɯ�5>/6u��r[	��&��9>ќ�ic�b�3�O��:���6����rlMż�����ʱm�4=�P೨�]�+�a����{��g�vS/T�@b��v���$����ʠ�{5�����Ţ4Y��=),g�[Ab�#��M ��ĭ��U���5�HS�r�����:�{����Z��,��$$�&Ũ��|�Nɱ{�'�0WK����C8�t�Mk��J�s'R�U�_4����4��:�2��y�8�ݫ� �}\����Sv��?\[<��^��РW���m�@��j��zrӑn�^S_7Ƅ�߮���p�+ �w�Ql������ň=/C>�`�v�WmĜQoH����X(K�(7��*�3�]��Y��lE���C_���Wa'�6�Au��5;K�E�t��8p�"Odꛀ1� W2P>�˅g�̦�jG$;�}��w;eX����jR��X��~��	v�RcjyW�?FǄ��8V���^-�Y0z���	��ߙ�5���eS��g3z`�P����1����jw��~�>�j��g�yw��4���J�`��E��j�X�+���4w{��sX�f��{x����5�sH�m=X$K�Ӱ�;{G
����v���S/��+F�6�u	�o�hg!��D�_C�)h�|\��R_4t�У��l͛g(Vؕĳ�
`M��dPUt�;Wh�3W�kĝ�<V���0g�����]oK�{\,1[��:��r�ِ��p�o4�g���=���nߞ ���~�(�� ϫJ�+��{�3^�z����;�T�b{D��x��͙+L�&���vKg�����}�V}��գ
dum�}��*W�8�U��mV�L�^�<̚�SZ`�RC��cf��0L���oş*���
{Iu
�~�`#J|����)�M�pM^�=���z]lyv�Lѣ�E�ʭB�?Uޣ0]��VAcҼ�ׂ#Vj/<�ٰ-!S��L9r��s2W�D���2���:�V�����=),����zA�[P�|5o��V���S�- :�F���l¡�D�N'��GHk9I�л�GL�1%ώv�e������3��UOB�S�-�	�uX�>��L��Y�et�=��ߊ��=����f6�/#oOw:���t2�|K��^Y���[E�5��5J�Xy�r�z��=��m�7�Żo���*m�n�U5_u+ '���F.E�4���5Js`��%,ŷ�h���^��%�e��3��2L�J� ��XH�G=RZ�������:׃��ɏh����>�L�N�n�/��j���a�
��*�7�u���y�r	��ϖ#���_lkw:���a�Lv����g`�]I+u�oK��Y�N���] ��B뢊l�b�J8����eW��Myh��WUc����O�"Åf�A¾��Ŝ���=~rd�=-�W=�^{M8^��˞+���ڸ2xY�Y9v�u��4�Wb��w��M��b�с{�mw��L�u�]L�RX��:08��	�r��$�\o������=�*�z���e��W�]�c��3iL�r�d������˪)|�׌*����:!o�"R���Kj���K
��>:%�u�8�����>�Vo��z r�����R��7�5�7|��x>}u^Be��w����3�Qn�����x/��#�w���3	l� 8�nu��3(Xe����;���+>Z�� ��v]���o���2j�;����H��\i��2��V������$`��#��ݳ���}v�#7��wO�����\�f��+Q�?� �.$=�K��Y��tc���>��UVl�������73k��oF&�>�UK�p�;ڕT�[������\"z�|�k��������,r��M�n��}Ewh�)���j����ºHYY�3qW��Sp�|�UwoǢ�+2�uz
�i�;��Lw^k�z�2��uS�`�Ĳ�>�h��*e	A�d7�;+L7h[åt睮c�t���';5�5�};y��0z���iBϑ���u2ث\-�k<��N蠠�ʊ����Τv���z�̸�)�^����;.T�x��ՉHP�,�<�ԆL�<�ʛ�;LKՕx���m'�^ۛ&��Ս���\g�T���f�U( �=��I��t��?2f���υ�o�n{��Me;E���C���X&^�AJ����;0�_���_c�z�G�������W�K�Ե���ë��V�yN(�垺:k�����lc�4/���SC�(�lE�k絒�i�p�2���"9O��ζe���W�;��0O\�`�sOwC�S6ƶ���乶hOK#I(�� Y�(��p��1�L�@�c��Pے�^��:L�rk\�΄�=c܉"��Z'>�hL�ِ-W�i�Շ��Wb:���ދ�%�d�=x5t��8�ʋ�U���K���*�N���e�ՉHB�W���u7]��
��wѭW)]�0c͆�!T� ෤��V���Ү�n��X��.�#�F�YJ�j�)���
4[{Q��=�)��u�7�$�uV�k�V�}]�@���^]n�R]8��wzL��LTk+o2��i�f�t{�WXz;[�V,�j�t�qfLo��Z2VAS�JC�mӧ�o�\�k;��i���կ5�2���3�H��ɤN��q�霕��2�O��I���s��:ӟtʭ���PT����8g�Kגa�ܨw����C~�oig�2T���0W�K�k�ϼ�2p/b��*�V�Y{�v�b9~�Ol�8�s;�F�����yX�W�+X$4��d�P�;����v�t#H�0�"��x��T��dK�v���K	C�\��8Z�+>�ip��N�}nfWp"���ؖ=Ӝ�7���r���ܦF�T���VȰ��	�ϑ�i�yV���V:�z�)Y�� ��e�B9q=�P/.y��*�~�k�����#C���Lz��,���:����/��Q��b�̝&ɟl�ŜpԤ)ιY�qs5��^��0���-Ĳ(!!c��1?tW�x,���;�Y��S�Do�0S߮b���k��=��k��~&}�N��b�f��]�z��E1&�8���{���Q�z���O>i�0�s�8:���{jn&w�h@�ߺ/8�j`S�>�Q��t|wEY��C���WV��d�{�W����hL�|�8u���3w'�%SՃ��,o�<��)Hne�]߹�Wc+-�t*��T�.;2�V$pQ+(
��J�+�#��[���&�I��Σyo��B�4�E\D<y�k��_P�.��9��S�f�P�蛘�k��g�����[�[�ym°P���W	B�3�b�r�Y��b,�"�%>
��p>x������o��xC)q����T�J���g����y`	SG*�#�g��P��oM�;s�*�}#x.�*��|�\0K�H��a�
�Z<3����;��߰��c���u㕳��LoLJ��&c���70=����&�� T=9=�\��)��C�lg����A#+�VJ�@�a��/�|:]q��� �v���s���ޡ�'�JV�Gʥ�Lprס���;UX��@��
�+}�m�Ȕjo�7�����"b�\ZЄ�X{*[#xm\������M�~�3�*z5�5��⃈ �9<l��ݪ��8�.84���B��iX��.	1^Y����}�D�%���.�����|-��h8_��j
�ɚ4zh�U�^��&'�"�,����B�]a��C���_�Y�*B\JV��="3+�� �yT�v�e�(�w�V��e7�m (��0Tz�U!�-ۑ!%AbY|�c}��qs��!�V������0J�[V�w�]�mƟ<�!n�W������ԚtѾ��yr�E�������W��<���P�c5�<�F���.h�|�����l}o�ǥ>��Sy�k	�M�X���� �#�]�Ð�jS����W3���w��	�z�2�o������L�&:"�t�ɘ�䄏D.��}����ص�l�L�R?{�������Mm��m��ka�6�	��;4z��mX�SO�����ݶ�FĻ���:��'�'�#�;q8`�e�K���~��u͚����̱c��Ⱥƚ�H.�[�u�^���K�`�ה�H��!��}�	��̐�H4(Ӆ,�����/t���s����z�{K2!�����?Cai�.a옥*��r�*�X�e��ݏf-Ԏź���[��f}A�deu>|���t.,���!��9t���">�W��P*��������O|�7����a�����]j>�{��r�oEd��8e<����˪(zp3�
f��w���$㖇�ݦ~k@�P���	�T��K c��l��n�<@�s�Pl[�<; '���]�v�����	�v�FW�Z�?JƇ�o��+O�o�=ϖ��}k;42���뉏h�C�ɷNj��I��jr���G$�V���[}Չ5[C;SǑ�B8f=VR�E�:�C-�C��L19����x�pj��ݹ��1M����vuE�3w5 F�&g}3����Q��uk�\�ނo)	%u7׷�;C��ݗ��)H��W:r�u��3]�6�P���w�
X�� ��v]�́x��O�H����le	O�)^O�,����^q.�������8e>��ٶ�q�G �n��	\pX�I
�>A���h��q36���ِU��05 ��s0j��_ }��lJ<�\Tұ�xL��^b�}a��<��k��\2�债�`,Ur���X����x�چ�/�W<<*csp罣/�7W�l�b�R�F�{s9�t1Qp��k�	�̂��*uǵ�w<�����i��B&/��`J��Ϗ�0R��5�s%<d�T�^����T�x:kɸ����<�>��4.30��f�|x\��J�
�6��i��
~94���N��۹Bc��lA����M���A�8�C��,X��>���8�-T�l��`����ۋrC�]�/N������|'�PłfÀ?U�MYz@����jT��44 �����
�����g�,^����	�i���D��랧2�v�`���V|q������x*u5�ҿJ��CXͳ�F��Ǒ˖}�j�v�E@:�z$L�QY+6��7��sN�ё��dY����u5Qf[6"[��`��B��y	��;F��O:[��,):�������1N���tU�C'>�p<��v��|� �}�l�e�xO����{[;Y���n��a�	>/hX����/�u|J�}Qg�J��{�t��V�����a��{��A���iY
q�dUGV�0A�R�T�UX�a������/?vz�ȅ�Ԙ��=����<�z��4,Ͼ���B��NzN|:*�@��t����O^�-��mN���W�ɎD�������3z!���9�VC��N�U���� �"EG��Vl�Z��`}/�Ɛ��o����[�̂:[��P�RЬ�r��\�K�{
&�����h��k4�%�����=�G`?g��r�S�����78HF�/f��3w��`�v���U��fL�"O^�k=�L�+�}Su�2��/�#��<*���x͢�P�x{�̏��6�D��(��ڳ�n�z;�КFz5^�����#^�ըp}gQ�U�(/DPV���2}��c��Q��.낟[Ȍ˯��;ssGE��<N#�h��Z�w�ysUӳز�d]0<�@E �6d��2C�K9��^�A�wH'L:� X��xcI�Dw"��Ɖ�
�p��4��m��iWzÈn;r�����g_5N�e��:g8��;�w^;�ϩ������ �t�3������!�:��P'��D���]e;D0?s�>�� ��<\��D{�Oy����,D��\&?fH\����2�2�d`���3�B!sZ���g0N�X�Ny�pe����ok��y��Y�(��r�u1��֐~#{�u�0!�S��o�q3�7稤�&k�#o���Ը���M�"��	��=n�X�Q�LO����_�V�r���U��;po�Sތ�]ݶG^���
�A۱B���+�g���ź���R̬�lE��Wnb���]�n򮎝����i��(l0b#�=�w���1�  ��P��� ���c���ֱ�r�w��LVwH�r)=V2K�4�ƎӕxCPoT�`���Y�����/O�rNT��4f�{�Y�.���)�LJ\�W�f1NgG8�����Ε;Δ&����q�|��t���.�*�$R�٫)�ǫ����Y+\$A�N^3���Qfg�}�ȷ#n��U���߆Ba�j����r�1�S��e��Y�FҺ�9� Ͼ���j��ffZ�B�wV�N�`=�r�=��sul�u2�	�:
����\����V��=}EՈx�K�ަ�Z/��;J¥2��Ef9c0��q�����R���R`���W������c,�6����hR�d�k�(����İ�.t{h��kC7��]�$��ucO6jR���ڵg��ߣ��P��\ �%+�A債xE��\`m;՘&�n���K�b�r$W]������wDb����4�>� I5J �"�32/�r�$�)����k�Jti��.�Fs{ʲٟ>�n���u�^�W�<wK:��Ɍ;ԍC@#6�$D��(�7g���z�6-���h�h�`�6��0�q�2��R���2�ΫSKK�����1n�TsU�뮛 ���Z����\��9"����t�ysi�V��gS��Z��!��� ���)��ӕ��CB�d�c����ʊ��j���Ǻ�]^��X�!G��Fl
���������b���������0$*+��b�� kS�f�r�frCۛ�3�;����{�D+鮀��]��oWc�(uc�h���lt�er��j���9��]u�ܭ��:oJ5,�կd�J��Gx)ӾYl�KmA;a7��yJ�&�cL+f�PR���9�~w��R�sL�;o�|�X�H�Z&���� Ц�
�FVr"]�iU`��3h�]��u��V�ߖ���7I I3)B���Y���+H��#v�+���\����8E0_w	w�`n�����}d���Q�:��h����5��H9Vw�X��'t-Fvҫ�$Agik�y�.�� �AG�B�mr�F��&j�ZwcT��T�p��c���II�Hj<xÇ%,��hŮ#6U�ח���ե�cL��lYov�Z�_T��Ykv�C�ě��9u�v=�βG�9P\�h.�oh���3�+ojJQ�X�����;NI�FB
鮹N<)^��sBh-"S�C�����2���
�������3q�}�D
�in�G���d�����Uʶu��jL����%���x*�7dle9[ִ��;N�ӧ$9�f���%��5S����[sG�ȑ�y���S�&!p��n��R���{:e�%�J��U7i�/� ��7GJsGs�m!ś��w�$�p���EJ���7�����T���s`�H�Kp< ڶ%m匭r�J5ʖo:�k���Q���������F�;X �\IX:2�|��iV�����h�ݏ�e�[J�rM�^�;��WU��ۻK �_<���1
}� N�Jn]�n��gd�%�8���S��'�F4{�Y�`骷��D���c��p[����ɇ-e�/wb�|�!�t���B���֚vy��9u�m���4�g��k��|��e�Q����-*2����U����%�PV�Q
�jT��������U��QEPk�cm�)Z(�T[IR"�m�1m
�� ���PT)m��b((*��QX��-h��U�Um*��DAF**���UD��Z���"�%JZTTT1EmKQE�Z�R�j�A�؈�X�R�Pk*�mdB��UEb�����F,DDU���(�m���DU-imDZ�J�PUb��Q�1�T�+"��KU"�"5�J�Z�V��U����(�J�QTb�-�b6�Ң6�A��[c��j��#� �%�PDU*�F[EQc�����#
�k%Z�DE��mZ�Jň�Fj��j%@YJ�FڪőVE�l��E���,Q`�R�h�aR�ekcmP�����b��V(�U��UF[*���*�
��%b����DF�g��˳����[�
�`[�gr1}��E�s9XΘ;-�M�T�aHɨ,N��� {��!��O)!����퇚q5�ۻ��(w����3+ҚЄ�X�Y�{�¥��\�~�f9q��`\��8=w���6ݟ��k�) ��c�٭�)+񒗝a}p����Rv9�M�s��<`�+i�c7���6���^��O=���!�.��xe̚����ˋu�Yw���~Md"`�Ũ,AH}޳9n������|�P��Qڂ���7��.ݩ|�*��fy�M"��]�&I2����*��Kl���Ϭ�F�c�1���G�4=z�l|���l�;����0�}j����(�<��&���bx�ޖʛ���+z��b�s��Q҄�ί���V9|�ڰO�"v���<V�t�\��f�CǦ�u�����8������8���U����G�k�,WPb�y��,s_b�]'�6���儊הҎ;�6��j�ײ�����ڛ2i��7��nO2@�����CsAك�(`j(���Xaٞl�03�g�Lᵄ>�N|��=���YY<.R*�L��_�8��ڑ���b7A��6�A��Φ7�]w):
���2�ݾo�g7sn�Զ�z�{s���Cj�a[����$m�1�J�혻���gDw�u͜��u�Y������k��Sy�~b}<��~��e0L��nWnzd+�~�z��(����%�(mm��9��]2�����ht�!��]#�Bq�=�c�e���'�E=n����&��7��~8-�P�۫��C=�S9Y�����ҫž�b;<R�|1�ɟ���t;�0+h~��,�iW�m�x=��-yh���x��إ�a|�X-�AQ�+x�ֻY|&f>�W�^�\ {����ק��|C��3C۟yd!g�fӗ�[��;�+����|������xw(ϣ�O�z�a3|��Un�xM�oZW�D�z>*nZZ+X�K�܃Jx�{��L~&���r�3��~������yd���G����t���{V�e��������'k�Zz�>̂����v*��z�]����yG���A�����΂������ؘ�&r׮�?}n��Ȫ����5��uJ��5[����49���6]��m�؜Ž�k<{L�.���>*�P�P��f����*��n=��B}�l�+��d�~�f�y.~SBHڭ����F/��T���YF����:�Vll��ԆL���+R�6��쬏�5&�3��4�i��^�2�G+�ұ�R�<,��*�#��T�X<��1ם$(�V0�˃r �����;ˍ���9��I,�xD�4��x��\l�i4���_3��	z���3D�r��ܹL<�I}h_Z�*��7:�;nT`�8lM��c��{�s��/�k�H�Rj�	�|Me��\��R�!{yA��4oS�����/UE� Ϧ�����巴��!	`���+�Z)��Y*3tv���7���`P�Y�����ߋ�e��
+�������<(��5��C :Y;*Ν-�ҏ����T�gġw��"��Py������g�,^�ܵ���a
���/�w�d]�oq(�Oy#���^�BӳL�n�5��r�܁���*��)����V��c=+�x%;\<����w�aa�MBL"$^��%w�|���Y��MX~�܀j�Off���)K������ u|�[Dx�d�S�l��mV��g�(8{�oHld,��;'{��;�f�������Hn��p:�[�|��� 0��'�P�pEJu�}i���ve4`�[�3���:ݼ#7�Nk���1YS�8L����)�l䒯u�5Nk�͊ѳo�^r�������J��]�
��/�!���<�>���n��2dÝ��
y��_e���$-�W�غJ�o���R��`�+l/��|t6J�P5�tvJV�����,�㺭� �wfY\�[I����P�u�|,Q���Ω�
@�5�m�a���:��c�颞����!w�@nl�L봴>6�Q�$��#�k]A����;�O+u�a�L�/-�{���"T4X۔�]zcg�_k~��V+�{Ǡc�{���:J�,����iHs��b�o	���L̵ޤa�i�5��գ���<�ƽ��j��@��p����4�*��u
��y�y#�ٸ�� ��Wh;L��:�ڜexqT�k�����J243�xz|�3�0�{�7�Y�$���ZM`���]v�%�0¾�� ���F���^��0��P�v�v@�]Z�������>"�a�wn� ��r�M��u��;B�d�%s)�:�t;:���R:^c���ww:a�$|Q�5��!���wO@iW!G��{�=~�~.i��۴�� �ݒ9���u��BIvhpD���t�X�Q�LO���ϋ��ۓ��b�Ǟw�(�f5e!�x��&�yzy<9�`���b���Jy��b�s����P{�[�^����A�w�j0٩�k+����-f���Od��`
�'A��x�xFI�_�qQ�]5�6�����M�H@	۝�)<�-��-:>�S�\�^jm|p�eY�J���������c���8Qg��4�a/�(I��(*����3\�f0�n�k>�֤5�q�ݱ.ݵ0.����[h��0�|�!���^{��f}�es3�2�4.�����I��U�>ĭ��<�h���{���E�`�6����Ey��t�sNT?��%Ir�Rf1X��<09�p�ǟ���кl��6Е�gKD
�LX�S ���{Cu�r�d��	b��O����o;��{��3��=�a�do�WZ6}5xi�U.|�b�=�4���̍�u�;�"@����\��~<��Q�C�]-YS�ڏ�Bk4��C
e
��d#�<����x�b��}[�	1z�
��8Ѯ^[M�^�wE[�M�m��]g����"�����R�.��ڱ^��u�"�׾�c��tu�� �ܙ�G��iK;l{N�1�y�)�����p��{�e�K���s2W�����#0s�e1Z0Թ�ױ����Ðp�p�O�%��?0�ix �Ѧ���l¡�D[��o,��bV������HճZM0�%��W���6����\��D��^�~ zD)Y�J&T�E��qN�@R������3;���:d5�֡xb��T2u#��}���o&�
��"��O)�)�`^ޖ� �5�����{"鋩dk��[(�� *A�wn
�����M�\D[���H����-��\n$��5����D���1($�&Ͼ��l����x],6+��(�C(��P}Yo��5��B�ʜ�/w���օL�G8�;\��\��Dg$hT)�36��5��=��^.,����{Q�ѷ��e�>��³�=��2i���	=l�
�y B�����M��c�φ��v��FP���3�&~�Z��6�r�ɊR��*��}��%Ǻ�~K�D��Γ�hR���m��s���s:î�>�&�Hm8E��@�s�FG��z�G��SEz�d�﷑f/-�%�P�o�׾c��L�s���r;���vz'�u��ָT�����O �"K����h��n�*qK��>����q�a�xޥ��+�}�x��29V���6'�y��ϔC��P���a]M���Y4䦗y�Q#��x;M�(�{�*x�'ET/��J�ޯ-}Y�ٴ��y��V�7ЕBC&w2!9���S&�_k�7)|�������Q�d�����]ppC� |r32�me�`1��F*6���L�t�ˆom�4��'%Y��tSee�e�oh�-mo%[1�2-܄�2�̼/E3w�Q�*٦)�Bec�Sv`7����p>�B�� Bw����[�CzA���[��7m�Λ�>ԯT���7|��4�C:�7؆�!���`,�+%w�o�A��p�3�ܦJ��yEc���|��2�����N��
�=F�XVl��+�债��T��B=U����V�z��;kaDF���y��|��`�$/O�M�8�?uɬ���P�b�|�[��1rjWr�ڽ>�a�Dw��1Y돍D&y����]iVt��ڰ�
e�f��(+�z���Y�f`�9&b��ޚ�^���z�8'�ڕ��]���\g�!eL���� �����ޭ�}�+�WY��)KY	C��:,"5?V}=|�������L�1oO =d��'4T��^��
�ʀ�%4YS���Øus�+k�qD/,����j΄���{kdӛ�����ژZ%V�^�Y$ʌ��[��ߝ�6߅�+Y��+E7/8�ik�e� �_�9�dy���r>E�#�Y9٦J�r����Z��yKp��1�f�!��v��E�e����[��#g�.PS��x�5|Ţrݡ3ِ,�Y��
S����:�3��I�}B_;9��yLMOq|Ҿ��ޠ���G�7҆�\�Sw�k{~tCK�3�)����>���a�FC�v\ջ�s��p�gYU�ӣ� V�#9�`�U��>�L	䙵�")Wvp|'k�n������)��)G{��<<���#޹Q,����� :r��=����i�����.�i�;�����J�%s�P`�Rk��~��ވY�<�Cu�U1H8-�=�E�8="�=cP;W�uv��vǪ{�s�Lܴ_��J^+���!�;�'�(y�b�*u�2�j6���d��V􁥉�p�¼W_��Q�7�{-��nd��z���5����ɛ��	�/�ދ��(�]�Zm2�N�#^��m6=�P�|D�������r�gD��ݜ�n�ZxS��8���>;���λ�ߴ�*����_7�6�C�e\���"ìI�z$+/ϧS��g�T�s2��F��3Ѩ��')]�~F�I�Z�>������UuwGY<�ly�s�t(W�Ut&.S85Q[S��qT޼�^^�w��k2�[�uɻ�����e�4FЂ�X���t=�9��5)S�r������L�8J�)x��If�������ra��l�@�!�ݡ=Yv)e�n�}N���l��	��0��s8 Aɞ�x�7F���+[�d�9I�/U�����3��S�k(�a���`�&�P�b����%�Q�?\�ֽ{�=��?5��*E�ÖV$/1<g���	Y��z2r���J�E\u�s���/�gn6�ِU�Z���Q������gG43�u��³ao�,�ptEymX�(f�Tz�9`��cJ�|�
49oy����,κ����VP�	�Ǿ�X�z-����� *l�4/�(�C(�a������L{lV�s}�wH����\�M`��X�~�C����-~>��N�СG��I	�h�Ǣ���iU�3uP[�/�M��G�
}�Jz���a�12����0G��yn�3X|�绷�1#�{첔� ��N*C��L�t�.����!I��pZ�^�PvOf/˶��Ջ�I˚�o������R�����<\,<,vn��&t�d�e�L�+>r�{��>�������N��{�ǩ��p�`FP���.��{Cꢂ��L�s��*Z��}x�ץ�6?TyF��a��^�5��'�h����TyT���-�����c��x����?��Nj���)N z��{`�r�;5W\F 8t��̪qC}�����'�e��H��"R����Usס����^[MگLc�rぃ�c4C�b�������R��z�<ʴ�I��B<Ua��,���!T����[�=�X󻋎���'$\�)�b��Jm��Sv��\�vRm�8�Q�֯ט����f���aZf��M{����ʺɴ�4�s����A`����o΅�0M�:�!�X�@�:��N�mL;^�q���
R�}� j��!盉���Hם/G�n�*D��Awդ��X��Xb��l��اU��A�T��Dfzձ�0�:v*8T����+Uf�cT��O����Ih�~`/��/ 6���ݶaB�Ow�X�����(�O�ӵN���Uzƹ�T0�d��֦:|���(�<Ԅ�N��8i+��%�<_��ʝ<WY���qu�^ʜ�K��
��+'I��'<}>Eh��3�lY����\��N�}����=��_�Э}d*�РW����凳v�V*��f��DE���u��ń6�#�-���5Jײ���9��S%�8�	=l��@PF��W^Q�������{f��VDE��x��3�a�7-g�~�Z\1Ξ�Y]Yᆯp_��v���R��u�3"V�,���)YB����aΧ��S9�a�C�,��)�!}if�mv���K����a�>m�x\�2�=	�����Wn���3w�q�7�>�ԑY�Ř�9�mv`�;�ã��_6%���Es|^�*.ݾ76	�h�K��q�8񣸉g͝�LOc���Iz����%��l>퀍S��heؕwJ�Άf�L�0s'g�Cs6�d�y.>�g�4e���kY�{���ͬ�����i���\2S��Q�T���N�lX���A匜[���R&6j&�ʽe��c)�S��:�x�n������^�B��4X�t)�݇-e�u&��9&���(ѱ(u�X3��1�x�=���,=������v#������U������fΨ1�}FlQ�;�{k4PiT5�r��L�����ႧN��ٶ�R��K$��.fh�Ū��+'K�F��,_�� �i�P��Ԥ7Mf�[+z�Qb���4�6�=b�.������1J�Z��<�9,��5��1G���~*�Z*���7�0��Wz
�	ϱ��so8�K�"�3^ 5�D�t�7���Y0�ò�Me�����<!��<�n/����E#�����PY�jS�A��@�0m4/{*T��/,�mofk�0I�P���:�[R���JM����%$�ږ�3�0�3��Wͤ�wġݣ������h�,�A�ٟ��CfWa�/�P�e�6����r�xĹ��d⾽�C��Ee[����N�8��c^-���Y0.ctM4w5�7�]c�1;�V�1��B��ۢ2�đ�o��( �G)�p7m��:w�x~�*&9ҵ�01:f��5r���G���ư#�;�iS#���ϡɷ/f����@�|�j��Ņ�\��fޛA'���][��k"�%a��XV,=���I���G-�`�9pw��YQfoJ�v�̶��Ƽ�(���}�k+�xߓ���y��vol#뷚͙�Z���c�$B���S��dh̠���J]��E�;�wb��'(,�$���B�z����k�������x�)�s�Ss�+��{�q#]�)�ἾV��r�=��'L�Z�xlZ�Փ��7�xS�O^�Y(e>�,�s)�9���]L�LsR�,�"w�W[v]��^�r��`\f��b�n��
�[�WV��Վ �,ݗE�1giO�9�k*[ɻ�ˏ��Z���̹���$LT��n�woq��rI�!�����;
\P�(�Y��\\�R�����9����(T� E`��[叻&�eM��.d̫͕�9�%���l9��z����v�Dk�M�*ج5yh�7�*��\C�G ���\&7KrPNw=0���긫4�r�N0G<�w��i��f��g�����5[G-���\50��:�.	S�F�]��[G	Yy��Zz.b)�h��p�^�Q����ެ�;t�[6�Z���{0�J�]��8۹��uf�iFj��:���Z�A��e�˜��n��|3��,����Qb����l�+m
��RJʍ�`�R1R-j�lH��ڢ"1V6�E�T��A`�ciE�jUEDY
�J����¥A�#(����DDX(")X��DEDTKj*[DE��U"�cb���Ab���-j�«F#EkVKlP+Pm�b1E+*(��,Y�Ұm�
T(�PR�UJ�[J�TT����E�Ղ��P�J�#,UYP�i
�AE�[l����E�1V�V�����XT*���XV�EDQbŶ�i@U[*"�(���Qlb��0V%B��������1dX(1���*��-,X�+�,QUQEQ"��h�DX,mZ�Ōb��
��b#iV[T�X�E"!R��)R�(��Q*1EQeJ��UER1R+mJ�V#+
�*��(�U�lR�Z�`)DPb#����.�P�����J���K�WV�0gvS׃�z
>�B��W*{���@�k����L�݉z�]r���n�T�{����Z.��G`WPp��u�[l���Yk�E��7\�]�8fZR�%���yd�^��G�Z�U�Fj���Ut5Y疄��>!���!�����S�c^�ݯ1��&lC!�>E�p��֠�H=�	����T�յ�y�I[Wa&�|؞���N��f0���]iL��}�8ܥL�/Y���T�c'f�������b���k�I��{�`�_�ñ-�"\0�<�N�=U���5 ��nffS%��'����|�z�sX�>3ϱ�Eh��:r�:&�w��y���Gk� �v[�>���9�v;��$VV�	c�8V��M�;��|U�l�>F`���*�	��]���݇5�����70��:��`���Ƕ�c��re��G�Gj��e�k��|Ѽ��4���=�9�hp�iЉ�upNؼDʛ�� ��и��BꙄ!���Q3��k�����cr������)jBgܞ2pWibtXDj~���差a��{C+��b<���*(Ṵl��3�O
}���gx�%�l�u�@4}�{de z׼�0�c�GV�ej�&o;հ��/[��Zv��k��4 ��/�:�`�,P�E��,��"��we�ɖ��s�޳1���o:>�o���4��ɍzY�(0ƚ4�ʢ��ʥ�ψgYz_�Eu�S���M�(���7�1��{��'N��~��xoݶE_K0�ۨ��^�۰����)�^Ӫ�<w�o��)��s_�]RM�è�S�0���_<DU�L�n�5��}�(���7�soZ|�����5,	���;ylt���am&C��eL"x�"���%���)\v�wq=V�|��Fg>fռ4Ĩ�?_��X��^T��Ci��p[�X�+T��)�V"/�_t���Mm�Ǣ������^d/Ovy�ۡ��0Y@y��*��*����G�:���uMZ������(����,	g��	�G (�O���xFoD4��\�1��S�&��e������фސ8J�,��<+�b��~���h�O����~���c��i���wlb����� �,z�c��q�?Ki��c�����	�H/o))�Ż'l�d��`�4���Q^����8��`����]$��iH_��{�l����ez�
g#
z��(�!е�[)��u*^`��ݸiAoyhD�{Lu�����S��x
�JmLY{��5+]H�Z�gl��K���l�r��r �Y��ozɘ���|�vք%��ܩ��v�3m��x���N�l�`�XP~���܃�Y<Hk�����Ѩ��ە��5�A�Z�,�"���N7�4W���\^Q�Ϯ����
Ͻ��3�Pu��^w�d�^��ڷ�8v��J��3��'����ryX�@.��lJ
����_��;�A��pz������֪�c�n�~*�����y<�B_���2�"�J�إ�Z���c��;��9SZ����,�=�T�Rin���lZ��j
�h�����=f�B�S��u���A���\[<��=:$�P�ʔ}7�lYa�}Js��l�L�@�L�B��e=n�X�Q�Le0|Hy烞�1�C��9�U�b���c�S1�6l��.���BP�\�P��p^%�;�E�����mz�7�Ņ�y��z��0�JK�n���a��J�{ ���P`
���� 
�3.��^�8�}V{�,�!�P�)��]3��`�BK�C�Ф��8-Wĭ��w-T����/�r���%V�.�<s�,t���m�9�)��P�oLJ\�T���6���k�����k(��Gg*��1˗��i� �����Ǆ����1��$ӿ�e��^�����}s쌜�D#e5ot��L�d���3�sC-�:����o��_'O�/K�=F�����,�h>�$��3 ﭅
�I�p�g(w�`�����߄��FϦ�*
�����.c��eM�� ��S.�'˧	�-��g٨p��g���u�����|fu�^tyT��r߬�j�eC0�/fĲ�rj���q׃��*�� V9�}aT�8!�^Gë`��=�,�J��9^��ظqK�����ꈸ|3ye~�u_����f�w��+�i����������Gr�X��B�R��ޚ�8�Aб�IAY][7���ãh8_lyv�Lѡl/����Kս��o��P�%��K��R{J��R�,��)Ö� Rޜ������s�ݯ��wLBP��J_�(��k�ݡ=�L��W I���v��T5x�q��ou�����z�\W}��0>5Β��Q6O�e-Lt�V�^Hs�&��c1=�$[x_�ꐩ�0*ͿW+!e=�X�ˤχ���.�b�Y<K�;�f����rpe�}���M���;X���{����j���V{�a��Y�wdP�]A��(��9��^(h����e% {c"�֬pcB�h���w��?x�O�<��AUyn�oT>�N� 6�˙(��Ùqe�dQN�H����2YB����*��'�w��]l�h�x>��iT2��6B	�wz��e��[S���i�]���{��i�l��Vt���˨ji�������BN~�T�s��ֆJ��@�y��nZ��x����s`�2Y X�	
4��r9O�u��z���XC�l-8�����?L��.�g��=�zd����FX��,�.���:�͇:��|���:î�"ɁΙ[�evk�Zjt�q�c��u@5�#�#Bq���d��f��\��h]�ð�S>~�����駔��7d�O�W`��c�T4S����A��$��*3N\�7�2�ʞ*�Bn�n���:zx佛�i��>�ཧ<@8� e9V�����ߖ��OԪ��j�[��-��&'�rA���L����m�h�(���<5�T�zJ�v��A�+|�O.����֜���H�f'd�x(~Z}u�E2j�8ܥ�;K��z�����y�\�ASۅ��l��'��ĥ6ނ�Xc7l�~]��&V��.R�ِU��1�[�4�/7^!c6���zc]Mm�=J{}{�'cѶlU�f�]��e.X��({��s�~��e���j��-ة!��fB|ŭ���&9���{D�f�kb�63;{ԙR�l���l���Rv1��q����u���z2���r�8s����.��<��v�㭔���z*�R�����s,��vT�N��I�y�b�9����Ӆ,��=�-$7�;MD'�;U^�����x_��_P��|��qu,SȪC������b��v=��]���s�O
wۭ��8˕�x��ڰ��%�ձ{՞oj\y�c�gPC�Ok��v��&Tܮָ�z���Do�#Dӥp^(v�l �\��K����'E@Dv��RV�ibv���jyX���m�XO���E��̽�{�i�I��%V�.���( ƚ4�¬�ϖO>;�w̾=AEu5=&�x�ǳ����mt.km
���HxpOU�MY|��Iu߬B��(6iͶ�dʛ���̮˓�9n�j�mO��^q���!TF#�O|�\ɦN�[�{2��(��:!��d����eǑ��d�9U&Ba����b!��I���@[���n�ܘ�a�{��w�m���F������%Kʔ�m3T�/Mq�+P�t%5TD��eVn4
�Q)��J7�.ق�xŁ&���Y7n�f��e���B��ڞ�����DMe�3���vBկe�ݺLB-n�<�M�:���腻�Zŷ�6��睁��o��ų֞^�>�Ʈ���M���xz����ݭ�CQ�����7܍���-��9�7��Ġ:vqUcj������.ݼ��}NJ���׎*;'R�m����p�ނt��yc;�	٤r����ߛ��f�CI�p P��쬺�:�~Z�9�MHȠ"_�� 1����(���/�죐�|=>=�o�{���<�%������]��^��	��1�L���J?Ki��X���!ጊ�Vm����ڲc��;��O�/T�����Q���>;���Or�;\M�G
�TX�<�6��KV��S��mG�Y��j�P���{��.%^��zE����.�l��'�B�q��r9/=˙�"��,h�E���g�[�s����F󹕣�NY��7j�kd����~��7�x�V2RX��Uh����3	A�aϦ�J��N_2ᗷ7Ƿ7w�1l�=2Fwz�>@�3���@���'G��B��}��$3�������
��jM�s��J��m6ruXt8EV54���4����.��T���AБ��W���o�����)���xy}7;�P;**K�C�&P�*�~��b4<�?֐x�M7�
v6�zl�n�������f�e�E��d�;�s�t��Sع_��p�M��Gl��k
�1I�����,�C������h���2���g��9�l�g�lf��8
��[Y41����c��V�|�M`��Sz��T�:��)�>(���t�-6�E3k��uL�mg<��"�5��ڀ�1���2j=Kk�6S��rUպ�2'fV6"���!��^g��7<P�`�G�����<�ͿL���.�ly��n��	��(Y��Ą⇻���N�g:D.�)�ή�O0n�b��0ίE��S�'�c�/f=]�Ȱ�/�+b�m�9�)��T9�oLJ\�+K�G���b�[<��R�ݡ>�a���00y��}h���@��|�QI�|�T���)n���~�����Tβg�v�r�'��>Wr�������QW����R|:��n�u��i�ךtJ�Y�F�+�*�� s^Aw[]��)�pC2�)�O�0t.�2�8k�)���$ܩ~�5
�����Tv/T��V�yǆ�2ǼtG{]�j��*�=��WLx�Gy��c�)Ws�e�4�Aп�)&+ul0gۉ��ja�N��ǐWe����{�H�ɰ��!b@`�����3�/%�R�OiS��-��>�ا	s2�s|��k/��R7z�)ǳI��A�.�]֤iPcޤ
x���x��Ol�1�Vt�j�%@�ە�Z�N��B�f���R�I����3S�`3��z{ vU%'vr8��	��%SǸ�,��ET�{��ܖ��r�,���������J|����W�޿�j
[U�7�WY����d���*0�l��9�:A8o��9hԔ���fi�i������!���k�Zl�d'���7��(�6����~zy
O���K�����H��]=>�u�2lZǶ��g��H�x] Ep�(�@�ee�Y�{���?ks�@���Ț�|�({�NF��[�)�k+��S,֦����ƈ�M%j>�k�*|O���_Y���<`3T�p��s���K�q�'X6�����[��'�����0��N�UX�)�Xp���^g�c�0k��٥
�X�C��3��f�]nI�ϧD��f9�g���'޺^�!o��Z\+Qb�b�g��ݨq}��o��iWd�f�j�q�E�g4tRY�wH���pO���$�K4�p\��j���>�j�[��a
P@���Y������qY4��v�7,
��4����p�¡�{%�LD�� ��2f?Wq%{�]*XV���=S����\ʢ���Rp[���vW���-W*�ϟ?eL �������I���DD���$�i����"*��?*�cѴ�oB�1W��=nx${2\Ν��ʑ	C���6t>�5�Ut�PNt�y:b�-������!����n\�U�=ܦOV�mQT_/c��ú�)�Sa-u�Ý�'źo^��e@�w�24g�f���ôu�kC���
�/I�:*��OD���9�.�N{�ep�Akv]���d�YC=�����X{�z�
�{-�q3��C�ZI29��C4��-[�T8:��p�|���a.yx:��z��� cRǮ�o��7!���'���Z{���&z<�#�}�-:+E֝9l�g>��s�紽�9�ѲF�r�s���4ޏ $�Bz���=�c�8v�Og�i��b�R�Ѷ||��3�׉��5}����4%f��H�FBab�{��V�[�f��	�3O�OP��,xާH� �S1P��S%1r��v�O!�+ /Wq}F"笅��K�,�ض=T��O�`�t^��X��H��d̤��%P�,N؍���kG����m�+5xM�I���Ax)��8g���0�0Ѥ�����~:]�/N�]:ǀ�����������Œ�亹�2��ִh*��v�w8.���7�c~!$ I?�BH@�䄐�$�)	!I�rB�$�	&IO�!$ I?�BH@��B���$�	'�IO��$��BH@�t���$�$�	&�B���IO�BH@��	!I��$�	'�!$ I?�	!I􄐁$���
�2����0��������>����?��>����_f�P��X�Um�T����R�J(��M�)U��R�Y�P�6�w��ݻa;;�Z1�KF�[3Mj�[M���h��Fi��f��t��Ul��-Z�5�5V�*�-���s]�����ŕV������)V�k,,���R�[f��A5Zm���Z��fb�Xa�����a��㡱��{� �:Tֵ�!(OX�W@�1�u*��7E����lV��-�j:;s�U+f��ɺΩ����  ]tth��n͑���:յR�:�
��R�RZ�˵*��:]��h֯`�޹��m)3 Ѷ���Z�mf�j�6��  =��8 QB��� �� ��� ��`  ��Q}�x�P
 {��(���Q�����m�mF��5*P�\݆��Н��lZ��L��x�  ��6Ĝ hG��k�{t;A���6�nSM0���+�n�Tl��l��h�1(,TC����LN�I<  /{Ю����P*te(
&wt��u5���@ҝ���k!�u�T��+C3�;X�F��խ����
u���M�h  x�wN�U�h{��m�km��P�� ��՚���M�P�k ;��w7][,4%�f��  1�tL-m[wvk�� 0ѡܻ�
�!C���ph5�� 7l���h��VJ�f�  ;<�� �.� #X�*t�!�(�.X���рҺcV&��1&�C� �{TF�p ��� ��p$W3 ��� �vi@6`(햰��t�&�f(�V�f[H�x �Pv�����h��i���K�iC1��KL f]�@�T���P    50�)Tj`!�h` MM���* �4����h�E=�&��J0 L�  10 E?�T�� �    %!<!�heO'�bbh2zOA�	4��iU*0      ˲�|{0��ft�l�RC8T�1�&q���:VS
R7�*�V��`5=H��'��`� UT 8�
(�G�PD������?P,�q����HJ��	!!K2Y�
�(��í���s��ӳ~B�
$�R��O�iF����;cM.`
!&����6��m�
cC,���Z��`�5��3p|·p5�K�y�) �Sb)�y�,!n���cP�����L����$���� v�SڄÛ��������Z��1-�F��O�=��@!mT��%���Ƿ)lu�̱mqp��j�C{aбr��ƭ��S�䕠G���E�1�f/�+�t�dW�K�z2%��Ջ��#ٶ�T@�Ŧ�^a�M�*��M����HZ:u�rܣyb��r�)���0�@n�yc���!�LT���w$��7iG�5����ijݠ.�,n2�6�U�T���n��Qm�փ�\А5A<�[Y&۹N�R�
kε��E����A�Bj�+P�	�n��h�ٔ遢�׸�ڙV�����+�H$WEڒ;�l5�5��LV%DㅝCJ�D8����`T��1햰�A��i^X׺J��c(fT�W,�q��(���hڡn�3)j�5he �{����V8i�}�������Ĝ�CE��]��+p�6�|���)b�LF��ѽئ �����������[�%m�]-�X'���w,m�/!��޹��J�P���f����@��
�y�z�B�kKĦ*$Q�-�žWI��q������U��Toe8�ԳX����[x�)I�@�Q�r�5Acv�&�j���[n��Q:.�>ܬ���P��By>gq�vk��*k�j1V�+k*�ӫ�Փ5�f'��ʂ����S�p��Qt˿����m�C+s�H�u4�Dr���{j��;I졶K��V�&�ju�`{����Z���H�h��5��"��b�>C --�;yJ��t�Xt4=��Q�� �RNC�f���J�5Zᰦ9J��?)�b[DK5�	V��5+�B��F靤"�35��τxPr�Jb��9����Ue��Zz)�s7lիB
ǥ��f��0��z�+A!�L��{�⧈���8\Vu�AFS"�G�1Q�/�/ƨ1KM6.���3jʽ�Ne��x�[ ���U��4@��Ԏ&,	W�+�fm�߷uPt����Z�˓V:��+6A
ZĲo62ƻ�����֪�f n�lɢ�4�q�R��vb��`^8ѻ�pf���-�Z�hr�:�,B<�@���!��ZN��t��ctRf�V`���r�Z�b��Y����Pr���B[.�3m;
+��P�j3�D1j�AJ��|�<�1�` �E-�Q���M��J�N�an��{\�ޱ��c;"L��dѺKC����p�W�%1�X�Vk؈��N�
�M�^/V�y�����Ej��1�q}��j�� )-�# N�i-��΋,�6���[�[o07Dʂ��BҀ���=�݌�"d�ZIZٗ�F5#L���["��Iu`ޚ�«(L����+љtĻ��č�t�Kj����F|�ehJ{��*����i�d��Bt]n�SQ�DEk^\�P�R�$�l0nФ0훸)0�/f��-�4�h&�ն�\f�(��נ�6Xy�D�ñ[hT˶q*�M�vV�Ed���f� ����@�]�Yy�նvMgVQ��\�,�[���r�s*�fU��M욣��02�kh#IP�IV%�hA����ê��U/7r�!En4i�4���N3�Xu�4ڡR�%�t�6����{�vc9��nbR����ELa�b�8�4+)��a���En�f��1�ޜ��t�`KkvT��l�r-Pۭ�R�+�
�)�jˍ�p0v�0u����n]��4,����y^4I?+ͦ�ە%MO;�N
ܣ)�WsN@;!R�O#��D;9�ML���g�ڣJ����I�ze�D������5*i����,�֘�EA 0RT��ɧ�-�Bh��)�ۤUG�,�R��e�F����(^��4^<{X2��!߲� �Sj�y��6r�[��)y�Ӽ�Fm'���fmǡ����8�3+1B	ܑك-̋o�W��d�9+)�x�:Un���*��.�+@�V^�3>;oC�0B�HNW��"0�Yb�'e���԰��U鹖��!��kwX��AV��~L�]ux4�5R�>�mn��p^Ö�
X���-�a퀰�l�s2�vtZ����j�au�������oV�6�6��91�T��n�$�A�I�َ��Ң2�t5�L��2�T�� Y��̦�����3Ru��)���g+D�W.�<{�įv�P@��cZ&�:�A�K��]▨�b����(9`bhY��8���hTLQ��^��������0]�����b6���A����[,�ٗ�)P�l��^���݋U-]�T���]�#n���F)�%䆡L��b��3)��h��v�;Q��'A�dh��@R9��i`V�Af[ͫ8M*PY�b���4��
����T��M0�Ru���9Ed�Bր�=��-�n��eGh�f^4d�G��H�Nj���x�(md�a���m�(��y�a@�SwQ-b�#��kJ+ծ��,SA�k�n��FF�s!��Qɰ*�&��l,�L1�Y�DW�1��]G���,�j�����p�+`I��n�5�Ȱ�gRB���nEmcRhM\0��W�8��Úg�0��oe��ŀC�]匼:�Q��b�K���\�[�ѶJ01A7TTT� �B�.��x�ڋ��V(\2j�5��cN�D��3�";AH�t��1�9� dؽd3����Zx܉lU�]�+v�0mc(��ǹ+0&�ٔ�t���S�{��P-�7wo6�3�N�Pض�3���*@)�3LN�R��j<ڹkH��n�T���-Sy3c�v�J�E�H� V�EX�4�b^ܧx�Rt0�1��պ��A̋wu^n	X�����Ȓ��:v�:4c5�Х�.���7i��D`|.�Ca����	���3v�$�,t=������E�/,M��1d�U��ɖ���!z�ѻm[P�)�5%�1+��L"8�5m�Ac�{I^}z�o*Ώ�IK��Qv�Ǐ6#�Д[ӌ �R�`�&պ�Y�h�7%G����^;�)�736WV�T0!���in )��R��7�Иv�b ̄��X��MP��I�VІ�P��#� ��t �Cٵ.�dn[Ҫ��^�$Ѵ�����ۇ�[�"�:%J3m�xvRsaij��_'*F&+�]E2�]\[+6�F����֫�����j�X'a�r�ַ+R���<&�)Ӱ�Ӌ+Y�Nn�ˈ�u����JVK�J�%��e��ZNdRemL�Ȭ�i�v�����xv�ċ�h�]̈́���r��i�Kl�Uv�K`���k�vn�[����s�������h,���̣B�t
�	����s�2�4���QSÁ���;rR�����U��nƝ��e�1m#ĖS�\f���2�I5�Qѭ]\CNnS#+(|
V��5M���F�mi����k^
�̂�a�ۛ���j#v�B���Z\s7M6�WKإ[-� �+~̲��eG9����EC�ˡxA.���&��M�G@ǉc!%�[�zMr6�Z��h͊�9�x���l㲫��?q�C�X�WN��]���f�T�2�~��-ڸT���m=4�L�&Q��z&J�ym��J�������Ռ�q7.��x��ڠ�İ��	>u�Pk7�7��i`�x�cHU�z5��N-X�-����#�;3]��su��H�o-ZAP��^���l	y�	��0�qm-Ŗ2�aš3�Vыa�874c*��VbYn*7K݋5�����.'��P᐀�ؓ�ի!�6Ѝ,M]-�,�R�h���km���.�e%���t��yl�9y��W�d�Loiņ�bA�ԙ7wĀj�ʲ��%�V�Gu��U�����f$L#3�k&P�|��������V�Q�HV�PJn.�8撫
�:(l�oNj�-�nJ;d�4�yS���be!�J��
P�Wd�ɚ�_�>[�ۤ��T�ۥC�&��y"Å�����3q�Dݔ�(��CYfS��b���Yȴ|��߲�ō�ERR"�â�m#x�hbܰ�P�C��h��ث'ƈ7�S�i)T+�a׆3`]��n�אeӑ��ڬ�3�7Zi�j�<n������c0�Ӷ0��`/�VZ8K[iU�i�m_v}�wk6M���"�ͧ)��I/#�e�9]����oZ�떛�T�Qx* Э|�8��ل7-��Um������5x�Tѧ��:���)�nkB��3sp$bR�43N8�n�f-�M:�X��/�#��{a;'�0�V�c%�n(�b�:�A����ٖ�Jd�ov�n]�\@9�\^�8F@7t@d4Ѣ)ɌM^e�2�([!*��g���u�*��,T_ʊ�f��R��xa;t��Bs-w�¨	Q!d�u;���0��샅h���A)1f�;e�{E�l#aۥ���,^e� ;pY���a�y�$�aO�u���4��[r�F�g˙{��]KR�Tw|F,R�7���t��ۭ�����>�4R�u��Y{E+�I�[�\�t ȪB����Xtp�Z2�m9{6�<�{P�H
��
'-���dX
�LR���-��V�gđx#-�Ur���ݦ�!Un�@q*�A���!�M�J��L�$t�h�6pXfٓ0kؚ5���˳OUkWj�'3&8sN`Y�q	���\7+�#���U����n��Io*K���B��t��ݘ��t�=�ه2�e���4�2+)�1eʷ�it���ܷ(�d)���a\2��ҹe�������NU�.A�d�`"�C�?����7�;ѿ��^�I%�Я�]Nz��;ha�uӔM�]M�8.�����TYk�V�V�P��u�VVq�)�X�ʋb�w|��u�7�2�hQ�o�^ȩ7��ջ��*TU�9����E�R%���d�,�f_�#�������&��`|ƙL�k�����;u����Yc!{����ZX�ӧ�P�	�ƺmJxFQ� e�����R8i*삑�B�X�g��$��,�k�$�-��P�pxLu��e;KL��L�c����DZ%�fͬ�b�]��FF��S�gv��b��ؠbn��K%�Q��z2�����pv8�ӄ:�P��:p$i�HfP�2���U���)A:-_^R�Wz.�a���[�.��8t��^��5�iՙJ�J�xr
X���J�ԛ��Uݳ���&�C����4�׸���2�λ��G��uj���"$�N���TDJY�I>e�&ȓ.�V�kx�ҝ��+�Y�{����3d\Y����ʗ%6�
��wPҐ��\�8\gE}�ŧ�V�\m�WS�pQ-����r�ғ��e8�����1��t�l-��_(esT;L�(�c��)��m�n�%&U��WN�Z�Z�2���Ծ�y�u�^	S:M��|T����E�6�`3WG�=�Y�}b�D!�PЯ���%m�FH��}�3��sM��.�N���j�`6�I��.d"5�ՙ�D��n��u&���gg6p�9e@�#xj��7*�4t�z1B����̩Ƭ�;�:�JwNR���eciǗ�e��X�Wu�;��}y��rl�Ro���5���P�q���O�b�� ��~&���S履ؒ���ԝ���8����u�u��Ç:���Q}y2�kVSVx��Ɉ
iiuնs����'0X��{�WW}��^��(�y�U.M��,ࡸ�#�b��,K�b����'T��uaZlh.�Lr�k�(�4�B�����f�(��fu��{ݓ7'H��ݘVˡt ]��IYk�z���r�fVA�d?�� ���2��@dV6���ˌ�7YX؃9i�X��fN������a�Ot�+̵�\����2_gwf�v&�
�u8�E�mKDI�Q�Y3{:rgWJ������Y�΂�����ܕ��_o�Ν�!��!�^"j(�nn��i`4,2vnI�r%+1�k���f<K��v���!��<۾�iS6�̳�^��GV��Fn)
�v��-�vG�o]eI|F��-q�=��8l�[��&�����:�P�LOJ��74'R��&ͽʾ2��m�I��;X)��ma������$�e��%f�Ê^v�K�%��B[ת�dP�������+�湫ܣ���Hc�L��v;�Rw�X��y;b+���Q��u]�z�˳¬2^ȭ�ީ�j��e�؃'z.QF�]��$�g(k&fv�ۥI��Gp��z#�5Tͱ�\p�o�`(%��*_Hm��6e����%�r����¶�sC,,��/e���c0+�y�ZH=�O�E��p�&�[w�jw��[�HVh^侓vPn�oő�u��#z�M����
a���c6H�weg.�+��Pd�m^�	I9�ٛfd����{�uM
�"�׍tt��o3	2�L[��o��YpJ�������YMA��S�W�7dR�i�(�p�P҈/�DV�H��N��.�y
�kw�w@;$|�'(�8=��8�4^i[Ț��Sٛvz���Ž���d�G��L�3��m�$F�LǷ뽴����ޫѵtn)��NlF�^(��b�.jݢ��39���:��wP�Vr�ۅ���(����sQ5��M�,�(K7�7��x�ӏ)�E,=\����.��b������T:�,b:T� 99�H-Uʵukޝ3 /G�1�y�K��,GJ��9�y��J����0c:�eL�u#ZѨ��v�0�
,����e���
���ckx��ϧ�����mIع��.�S%
.C�����-���J0	ܸ���-��;�K��OXW�/�Wjc2�f:V.�JS�4��J�i�g+���=i�}}{��Z@X�)i�p��v��`L�@��z�彬�G�k���MfW=M(e��N;�H_hY��\�����VS��XZ�'Yx�*�%��J(%��\��F�	5�qdR����]t;�b�F��j�#���}��@�pp�R.jML�Y`�ʚf�Zq���w�]
�qR>�	��`ΛDAh=���gȹ�B��r�s5���[���s�_�S{Ԗ_<�v
�m�j���	%��+k0�e�n}�wd�{Y[1=��c/+n�Rq���3�bn�aK���aӱ�%cȕӭd@wN�7�×/;�<O���[! nR��>�ɽ6��l�de��j�ͺS 5���V���̾]���5�:�"v�M6R�!�KJp����WnWd�p��շ�6�f8�6�o� �F�$���2�3�]����WJ[3��73���1�:�u��@i�R������E=���Z�]s�`�\�d�]�2%����R؎���9���!�J��Y!��ګ�=��n�B�.�V����E�2��s.��/���woL,5Y�v�u-wrV�iǛ�^Fki5u.�+1Rw�jY�V�{ ��;O������F**�E.+Ȯ�����>� {�4	u����[p��H2)V�r<L�O�=���چ����*�i�a|9��m'{�{1u(o�kt��{��(���y[����4z�0U�I�m�R���"q>�� b�y�Eb��L��݋�{8��`&ؾ�E�T��ZJ1Ɋn����yJ' ����M�ՌX�ˉ|��"$Lu���&np�-�ۜ�F�+����v��p�����o�����P��sWAweB�S��������is]���0�!v�C1!��]R�7��v�Qb˔lrb֓l�o��)�V���P�K�U�p��g�>m��u{.�#w V�``]1%��I�uv�!a��w���G T�>�����6K�$�Ւ%Y��o�5�Sk�%��s��e:Z�S�m� �=�b(����f�rD�u�|��I��F�Dn�6M: �N�ZsU��.��܎�-a� T��Ψ{���@빷23:��ʳ�h԰ʷZ�N.��
:Ԉ��u���
���Q�c%�@㦙?rɬ�X{���z'յ�9�\�5���BԳ$}u�!�xd���,��e�k1ެ������8��M}­�B��V�c��m��{o����=�{KpF�4�zL ��A�vn�/���n�&�I`��ʭ
�����ZrD3D�ܣ]6�[�\Y1c�gO��0e��xrnT��ir��z����iu�wtw9��T�qU�#��������ݟ�H�œ;�w��j֞�'j
te���G&SV�H-�nD²r�cQ���l#)�]|��Ru���xLU���,;�Ө�&���<��y׮��2D#�����K�b;���ڴn��E��g�ik��U�V���
��R�qw'l��@�oY�� �X��'x����=M]ݲ�W���[��\���7���-��%�)�Vwk�蜔y_\3-m�9I��Z�X���������'P���%�8z#i@T���qyզ�ڀ���6�_x��$��[���"��*�#��v��OV�NA�ޠ���U��c��e'�D�xN�U���`�'Ph �x<�r�[O�hh�{%�aL�s��_-Nl�C��E�Ϙf��U%gpP���*v��<���q-��7�{��\�o7����"�AVyDv�h�\� H=E�T�d�"��,(��yO<�Z�e��~+b{ ��L���M,�3��(��s�s"��W��d鍽�̗����!Ǌ�ܦ�5ָ9q��!8��:i1�';D|��z�R��7X�\O`#FjH᪾D���������p�י��-ݪWï�HN\�\���j�iI,�p��	
�}�2GKj�E\���f��-��$7YZ��y):b�.9���sz=�
���B8��X)��{�I�<k�3��A��\M��w��ũv��˝�+@��묑01�jp|�.����Vw;�9g��Y�������\�wx�mq%k^����w@;:D����������[6�^1ݡW� ��	}�2p�T�^T'���S4�j�t�^X:0�"�/{�4�W8Od��J[j*zWY�W)'$e#�u�q���V���8��� m�)V����gGE���c3���A�霛��Z�B����B�Y�L�:�5�����-�����NIr؃�����GK}��r�Kw�d۴��R����&�r`YΤǒ��V�ل����+Ť�GQ�`���$��\n�p[J�@�)��O�g.{�=ơ��Q�q`JOm�z�wj�EH�35p��ď&J$�j�k�㇈��oRQʔ��Vu�y{dG����B��h��� �ڕd�VҔj�h�E,��Kcv�˫H�ЬYR�t�4v�z��h�}R���Q��-�;���t��Њmj����b'Q���%v��ӽ0�R-@��Uݍ��N�y�4(z���oM�S���$�`�7�u�tB=fM����������\ݔ5�,]r��<�Eޕ�w����M�ГS�s`�_6S��Ւ�J�^��[Xh��U��36u֍X�����/�!�v\�i3Cq'���jf�.[*������r����9���tR3�q	���е�o�w!M�x:S"��8{���	�F��fU�2R�o�Ind��[mqRboA��5���K����Y맷��T��Xr0b3!�7�w(��u�ZsA(D<�0���`��jgE9BeѮ��_8@��{�w���f��X�@�l�!����PTMwʠ��\���T E�1+��5�$��G�@����e��*�L�q���xQ6��j����eX������Y�u��dv̀�,]��:\�u��2e<ThG�>�Wo�N�u�óz,�����=#N��܄r�5#��-.y4i�E<��mM�_t��.��[.�����n��-��~��������/�K@٭K���"��#��ԭ!�We="N j5i埵`�^vҮ�q��h�$�.��]��3�s�b�d�f�C�-����YAf��{�j}j�<��j�pC)�VtT �;�J�j=$��%���YH�����3h�a��s i�3�7o�]y��7Nf[mXU����t\E���`�5�[��wf�Yo"��>q��n�@�n�<f��}|:T�ʅ���bĘ��Wzu�jr��<��:��1�E�@U��v`��՛Ϸ��[0˼U���۾X�L�ű}t�j�x&,��'X�4����֍��:T����X�J�#\�hq�sN��SN����o;md�t3�Zi͘f	�.�Y�Y���	��'�y[��CL��oyj`]p�I�Z��!��\��w��q���c�᳠w�X<+T����K�:�� ���X���{�o����AM�6��@�cU{(�UBN������>o�*��&�N��Ni{Y�a��*L��2k�7��2p��PݿjGi]nQ�:5�X��0�9��"�̼�k+u6�XEA��f�W�ե���2� 68�K��®�S+6�@�;	�z@��Ȍ��X)̮�9�Y��W!E*����mFS/�snu����P����`N��0�ɽH����z�uۄ�@��6d�X���-J_]gIg�xO|ZN,ށ3"\�V`�ulX�(FL-+K�C�����{��R���u`�4��ԩmu�nu���S���r��ewkG���iԣ"��e�H]*���}i�Y|�E+`e�k�e&e��&dV��Tǁɛxy��.Z*`���Ep6WӶ_�1Ɔ�@�+np�6e	���_\�Ai�Ec϶q
�=����tr��4�5}�-�=w��
� �\����0��N�e2�[{���)�OO��гԲ$���=�Dn���Pg���N�qڴ_���\+t�U�n�ҳ�`�q(m2	M�2���[]؇`&��+$��p��2n�6��.#q�%�ůIu��8��͡�hQ��b��.��/n֚���ԣ��+#),b�b'&�	�XL���<�i$�����U�4���h6; ���+:�w3��M4㹗�X��tzl��[a�\�����w�>��v!��.�b���x�[9�<��7�b��t���a�Vu�)Yh@z�j����,�Ӭ�Y���)WX4[[ۙ�Z�U��am
CXl�]�v���x��fS
���eA!�;\��=㶟�T8��u�E�ǔ6��HF���@�B7n��<�l��sD�y�v��j�*�3�vb{�9jt%d�5޺���V�b�,I�g]�Q\;x��]OU�G8��J���-}s�*]�Nl�NL:+�;���:�a�z�%�@�εH!���0gf�5'y�{a] �t\}[F�-�������Ԩ��1O�-��-	�g`/1A�vԑn��j�$;����4�q�a��$ ��f��'�>� W�3�~���<���ÎFF �i*�ǲe�D���Jܲ�c�ڠbMVmӆv�7��]f��@nZ"SM�he*6Ʊ��5�iF�\T����Y��붜5�"�N��\Й�a5�u,uCJ�N��b��P��w_q�§IwX�>�:��Y�-���|���oT���D�u�vX��;�fP�y��[�L|蓔����*[G�E������w��Z���f�\r�R99Ũj�~���',��G���H��d�˳*Ȓs�G�<$E�(�D�-e2]�2-�:�#J)��2#]�l��M��xs�a1�X�I�Z������=�����7�����k4-	���:R��M�E�3�� �YSywc*�S�6Y�q3��c$-�#e6��� �v�E�:�tѵx�nL����H�K�xs�L����l|N�u��}fH,���i%��oo2V[r�m%��#a�-	.��8��t&��D������#+U��$�&��O��^�W\�����w�̽Y��l�֮�,l�(��Ն>�or���Y[F�����`7�e�d�CF�a]v�%�[��r�����C����:~�p`��u �B�;k�5/���rc���}\�;ӚBʂ]VS����JJ��2�N�LƊ̾f��8i�൭+g,�V�#i�ت�Q�֒DG�`\��l�X3Y���Q�En+(JY���r0�&�j��U��Y��.�͎��B����!D�k��XUꂬ���]�OA���D6/
�����cS��k�H.�j;���%"	���%f
h����H�-�C�Xv�i�澉�W�ff���+���xfq��l�wpS���қ��>��A.��/�$J 5�ٳB�����k�4��]xj��ǜ���U@�]'��nJ��u �,��Ɖה]�r����Z\̄Q	d���nè��t��Zj8�4rR�>��T��N3�ݼ����u��;�A�h�̦���:h=fq�t��\'Z��z�_�D�8N��N$tJ�l��1�Ղ�x�k2r���3�М���:�+qY�8�p��وia�Ř;v��8m\뮆7�P}�ԶF�ú�Z�d�S�۹�2�p��M�r�(\��}�kcA])���#
���c��u��.�C7�$�%3/2��{�\W%/,����Sن��8
躼΅�괪7>ə.�D�RXy՝PVů����y0.�6CjF�H�m����u�)9y�L��BE�G��gaػ������s��7�T(�����^-����%:J�pF��uGWú�*5�3(-����QL��ɥSz��
U�%rK���|-�5ǥ�N��$��_iۮXZ6l�oN��2�� ���s�ifqQ�GSk�x�|�P5��;kTu*8�JiҲ����,�r��Ev�s5��ӂ�mp5�� ���B��ʳL��6��w$�(����<籡:T�/�6'l�p���9so���-T��9�r�!39e��5�m�P؎#�b�j9s\tr�eS5\J����9ˢ�6cnqS7Elg���/;T]W�d��U�o:��+6�uuZudG]����x��AG2̓n
�Ӳ]̐Rjvwwr/$ǚ�a��Y�����2�M�V�����1��J�p�%�1�=�}�$�U�\-ҁ��L�D�uy]}�7ٶ���P�:�[@�8:�Eva�[[�r�����Y�*"��H��M�n�ɡR���z�+*�o�2h�$ε�Hr����-Q���k��M$�֋qj��c�v����[]�ҡ+�Z(D1Ef�۔kt�Ši�7�C��V����P�B�7���м��J7wK��ϲ�+�����	[�{ ����Tip�4��݈Aܔ%���W���jKq0�F���&.�D��ou@8�	N���PJL�_WS�h�-^q�z#8��_�������$b��ܼq�xe�o�ʽnZb��]��((�@Ϋ�fu�(���JT*� v�\�4� 9o��M@]�[�c%����&q�+�JT(;D�w/�a���=Y��E���]�Y�'��
� ��v��I�T�d��n��46��'V1	�J*�X�������²�f�#��i�*;���0�n�p���5���Z깊V�#&^�=r���d\��L��C��gm	[G�C�o&7AT����7!Y��u�)����J�x�Kf��K6�1)�l�`3�Q�I��i��_�fj����t�m�QTʹ�v�z�:�"��sx�|+#a8$�X�qIl������֭�N&.�K���:�,+J�]s�ڢ����]N(�V��Mn�76�Y���=����&+䍂AonT\�2���b����?v[ɐ�͡�����zl��P�A�Z�2��T�򕿤����٠�[Kx��
��>�:h'�h��(�bV�U��S1���E�X���hY�tJ˹�9V�Բ�]�}!�s�u���Ƞ�}Y�ث��/T�j葫&=������Q�����s\� �gc���Xz�eM0��]�l5*���;�G�-7i�v��g�,���9MP{y�%�9ݦ|r��Χj�{gL�q�D���z�����9��-{/Wu�:��jf̤��2�{'`Wu�t�t���X9��Tq%[,X��ΰ��ݼ�����Z�����o��u
k)�(�KF�@�gk7Ŵ��h�t�IRذY����ce��8B)'h�2���l���3%��AOo��{��b�ꎤ���Ըl�l+�7x�}��}\�0[�2vQS �!ՙ���3w��)V���XRr�pP���(�L�pmՃ��4<g�J�7h��ܗqW_b}	�3�e6���[|��dX�V��L.:Z�r<�vðkq=[A��w8�[�ا��SU��ݸ�*vҫN�(lc0z�vk~x䬴��:��ie�Nc�1k�K��ȳ��������U�r�r!����k��r�*g^�.��;v�c�̻'���r�At00h��5�4���Ŋ��'2(\�	�uwZ��Va�E&�Z6��,��{Q��u�'F���!��݉i�Ζ`˳�5�3[�N�g5�K`9�T�h�m��K�y��s+�u�0��7E(K�-u�����W��K�h���r�+��bZյ�&Ի}�2R�@Q͕�@"�dS7��$7���VM��'>4k��=c�*��H�y��SLjTuA��uu�yz��H?�c�kI����7t�P��.�b�;��U�Ю`����[>�"F�oYy�X 
9J��U���;. U�t��>)LX�whGyAuñ��r��͝uݭ�܂!m��c�9Ek%�4ۡӴ�۬�Y>ck��n�8ޓSw��*���Q�I:E*��������AQ�Y����\Z]�/�r��J7 yDU2���<�G+�y�]���\��O	�L-�x�n�XBWP�+nj�[}��P�"k�Z�M��lδo3�Y�U��ݓ1�h��ڼ��cDA�TV���w;X��@3���X6���v�%>p�݃y_R�����PPeY�}$�+Y���7�(H�}�н��]���Cu�D��RsY�"%>��������J��r�Zz��EM�M[��kUѐ�K�F��.���5Y1�Ȧa��ْ�Gc1]�
lfd+����a
pP4�~S���s϶�E������*�)\@Ѡ����:��噀��zzfV�,+Yv�nY�@�#"�aYs2�����1��S1�
2҃l�f�uָ�ʚш�����-"�PZ��k�X�جb��Ɍ�i��QLJ������X\���`��W�Y�m`��0�Ƣ�U2�SmMI��C�v�nb������X�rܻ�E��ʵ
���q�f0Y�&Z5�F\�S-�Q�Sm���,Ƹn��*Ҡ;b7���[a��*��2�u�����L�+5�%��LT�]qn�E��wr���Ma�n�]������E�R�\0�Vcr�n&����X{籓�npcY�ʁE� �{�fu�	�am�F�rh����]	Eg{�[y� F�?�ٕ!5^�?Ғf^|�����hEPܜ�ݴQ"c���w�rU&�㧲��/Z������Ll��5�}���.��f�B�a�uj��gc�B��mG#n��=�4�!��6`)�=}%��U���b��;��G�$CLq�
3l�Y��n��c���G^9Dh���AU��-��J�*����Ⲵ�*�����2���'��!j)+M��1�;�6�(fe����v����h��j�>hw\�ҷ1#\��e�]��c�Ì��G&b��߭����<��*=^p�ueW�����\u��W����wѼ:���2���ܬ]Qn�y�jfU�̙Yi��?�#���P��ʙ�/��A<�����v��U),6r�r��c��;ͷב�y!��$�Q���zqv��}�'��&�h�½��$�~���]Y�VRJ��)��v2�h�v�^y�u:��{n�y���&R ����vr�Y������,0�ʑ�����J�z��^%Xɕu���b��i���b�8؞"ڗ/���M��=n��H���g�pb_�%���+���ּ_OV�ebڹ�;m4�խ�I��G:����Q)H>��5'S��|�fʭ�z�Bq�5��ְ[�o�%n�p#�����WO[e���wK��K�z�[��PhI��K���r(V�)eT� �MbW��`m�`�+������w���iX�"����9{1eL�nݥ�Qys4�W6oLj��g9��N��nf:�|�x!�4��!X�ZP]�\�9;1w	I��5K�w�x:av�ٜbۚ�46�pf',����7�y�!�$Y���ƃ����.�*�W��,�.79RDj��z#���pS����j�☎��{^�>�T6�J��zb��^C��+\Qd�sҵ�>	f�����S�Z<�Y����鼺��L�੆*a&r�mu"}e=G�`q����d�v�ֶ�{'�V2��w�Vh9蹳���^S���!e��G5�q7 7�H��Kh2ɞ��jM��oiX�Z-����]u�^�%��73y��D�0[=C)k=��Xl�W+�dp�r��^tC��d]�d�2cg�R�ޮ̻�.Eh��W��2oyWl{i��L����:��À�LVN�%�5�|m#-�4��f��\.֢�s$U�P��5�{�P�Y�������8���jI����k��@�}	d���N�-k-ɷ�S��z�ƛ�K,�R�hk'BvR���F5{��͈���k3YI��ͮ	@�#-쐞��nƍ�%�nj��Qa��c=��~С�>����صgj�$\lU6iX�/���#�i��t���/���'�sl�m�y��t�Ve�d�,)�� k9þ�� ���+e���B�4��L��{�:g�C&
H=Bs.�z��y�D�+�wcU�|t�/�lwSN�XB8�U��p!Q�ô�C�pw�5&���gNT��@EofQ�g�]��i=��-��9�V�[Ⱥ���Y�.0y�SZ��`,��u�gr���5jEc�ݚih�*�MDd����)��J�!N�f�I�|���E��.f��� �O�!G�e���Mz�:79�RN/��* ���´B(�5hp;�����2�gbUû�祡�"�H}+��]���*�X;��%VՀ������)�(c@tbzE�Cvi�G��#!7B��TOj�g��e��B��è�� ��U�G�Y�_��54������$�kt�?!�Z&���,�����t�/�сp8'��cO^o"�91M�ch"Ԉ`���I�r(��{U7C�h����^�!O=�����بҷU8C�%H�(�dW��)�nF��C}��wsA��tT�H��<�|l׆�Z�Pu���Z(� Dr���Q���M�b�aKP��q�r��o��K�
(j��L�se�ݏXj)a�휮�0۝s4/�.Y�����	�ڲ[�.��S��v�Rڜ{��7f	"��l���y�i�Cn	�ǘ'.<���㉍�a�jJ��m���^�� ��[k�4��]KU j��=��\KSqNh]��)�)0*Ƞ�d5K�$�U;σ���ab��}�ߊW��6�t7��X�e�)3^����c Q�W�]���q�]/R�k����HOj
��Nbd��YtxT�xW�1�L���6w�cd0�
�7d%�݅]��T�Q8����jԹ�w���2JR�������<�G�z�����'�����O�s�t�r��9�2�K�I�B�	I��A3["������M���4��V��Q�����9)}z�������x�)�������D�s��&��#J6` �2�m� DP7��dx�
ۛ���{����Է.�*v�y<�Fԋ��A�� �_n��R&�4���D���yB�Ss~�5��٭�ԗ!s�Yz����4K�!w;@wP�A�S2p��C�>�*Q�/�xmI��.ގ��R�=IK�]���X��%�_q��2r�\�Jl�B�-�v��6
W�3cޞb�TΏx���D*�\��a�O��j�yŴ:M���^�P��ˁk.ãX���p��
TG�!0c.��H%0�y�D)q�X!ҀFˁ��p�st݋*���x6z�[<���7WP�
<`Nؘ�t���]��Cs�}�\���z�!��p*gO��D�Q@(�{��6�&��Ѣ6˞�������U��pk������+~��k����ޅnw���0��D���O��*�_�aD�Хe/Fwe�������h�a�@̪� !��1cx���r�|�R����aA��M���*Y9S����X��2���r���ޑfE;�FS,�VD0�6}DME9O�m�F9: �rTߜ�# tz��[�
�(���DЦ�\����u'�aVQ�,�;�B).����S�#�kɻ������WƺBYT��4V���N�d�9dW�Q��;�Gm�� ���Ʈ�<x�+�u}�`W��
?*�Y@��&�e�*ï��l�eT���E("Ԩ�]]�35�{`e��ةEǯԫa+ja]��&jy�����5e�٘1����;G�B��ZKh	�,ճw�l�l��)��덅�.����_����pN��
g�M�S{kW�RJ/��s���y���7�P���ũ؝�3M c!V1�l�o�i�0*�ѯ��G�E������Y�B�0p���&�M^C�VZI��J�@�à8GE��&g�^�Ϫ�Ec��~ѧ��,"O�I��;���q"4ȍ��B�P2���+��**:��[�\g�9���=+V�yW:⾥e�����+�Ή���V�'7��iq��O��v���
�/W�}��Ѭ:�ޞ�}J�}�q^G�x�^޺�_1�%nKbh��'F,�������vEQx�}*��[��ҭ[�y�On�vd�t-Q��EE�ǃ�MB�\�L����t�o�V֙��Nr��/�'S���
N�7�Ն��Z�2z�7P�=��(n��0�T�c�S�u�N���������<�\������_foTwaq�O�W�Q��@�%���_�c�Tko���3=�1|��V(VW*����})��T��?����-����4�#ad�>��+y;,A��Q��Ѯ
�D}�)��w�x�愘�(�,eSlר�GL��8�۞J�Mb���ψmZ����δ�'Dz�X��@t�^OE{:���t0� �S�c����G��~�FZ�)P�@(�@�&ō�S��r���n�)R�P�՚�!<bS��I����#�C��G�Y�_Q�ji��C���/��	�71�|~M���-X��?\������q� ���rS��GH"��J��z��=���R�Z���<�q+�b�óx)��E[��~��]�3�Ă���ŏ3=�y�f�.�V��1��]:)��]JV�n0�}�����Q�_��:�{G:47��r�KZ�qvR��	�P F1]�f�#"��zd8�Sbw8�n6(nTs���P2�n;��N��Q�@�U��P�O2&���s3Ŏ�1�J�ʈ�.xl���7�!���B8ȝP����u�Ʌq�J���,ȓ{j=z�(؉���#� 6v�FE����J�<:�&b��O>?����׼ku^�9�����6�@АӢg�D�J�P��ܗ�I�y�x|o>�yL���`@��Wu-H�������7꜁gy��|��*�5�݆s�o�=��A8����^x�_xօ�=4�r�^U��8R������K��͐�x@��Uڬ�Ǹ�ĩʢ.(���\<c�&��Rr�[����ƅ:���l9�W�W@��c#G��#�~��v<7�D�=���Cߴ�Q�h�;x7&D����塌�o��c�6����sk����}E:�[1�0���{b��<�4�6i�\��գ�,Ŵc���!�l����0��o������R\��4^8�Y��
{Q��;$�NӶ�R���&b���侾}yB`�j0�Q�k��`��f(�mv�3eq	e��2��8�D�ћ�TP��l��ȪgM����ɝ��,l�@�9�>#)e�f4Mr*o˕�x�;��YGb|G,��xĂ.����e!}ܪurɳ0��ۺ�L9���-Q�ǝ��gD���i8�بT���M�YWɽ�v>��;2�˶~Jj�K/�V˧��-�SSy ]�>R��ڰ�<�N�5��㊵3MN�ַ�^S���s���#��Ź�A�v��%K���u�U��45�<ū�Bk�-oQ:�.��oQ�)'��ř��!ĉ��e�tR2�'6��i�A��U�qI���z����ܰr<�va�JD�?Or=T�=yy��]E�yq#�l�uK���q�uAw���Y9�����o[���7Z�o� �-,�����Z�t��]Ũ(܍;gr�X[J[<���^d9*�q� oX:�̳9'ılRUK.�_h�O��d�"�Z]�uT͗��!Rݱ�K�qfhX�ɨ�pveEkc�TԾ��i�Vڡ���Y�5��e+\�M"���d'���p�(Ʋ�nh4,��8ݒ)�N�tn�Ҏ>)��M�\7�aU����X���lg�aۨ�N�jE����R����B�F�4/���$F��N�x�aK��κ�d��þ��|�)1E}0�ʼ�sx,�\���)��So�k�
�[͂�"Wӗm��.o|�E�@����5������-	��!� AG|����f��0��mH3y�LLtf�g���L!�Z��ٶ��s�g^bͨH�M���u�y�h�sW�%��8v��!�Ȧ4�&V�A�7L�nbd8�Γ��Fpf4%����vM���x뎝!��|;x�j��!K������?�Dj������D��9��C-+�D���[,33�+j����0��wmɉ��K"!��Je�aUG��ㅆ"�S-�-\�Y�k1-�v�2ədęnb�3(�����3*�nm3sw&V�iSR�H������;b�w.��Z�e���n��cJ�nm��Z�)��D�Y�e�
�����.��m�:��na�(�p�R�m�2���EۢV8�L`��ֳr���mc���cALT�1�*ܫ���r�w3-���v�[�n`jaiq������Kq�-�+��������T]J��
��%h��+5�����S]Tܻl3(VV���GZ
���u��֌���������M@R"&<"bD��N~|?.����ʲ��!+�}S�������L�&�h���Gċ��r�Gs�F�����%�s���@@��pk�4U�Tk�βQ�ҮE+�����Gv�x�wQ�_�R�=�4Za�L���Zvr����7���㟮y?^����v;<O�F�ܿ5A�K�.��uM�:�L� 8����*M�+<�Q��a׵M����Gj���FT�!�|%_O���(��ޓո_���S�;	`w�3��a��&fQ�zF�^r,eA���E�Ԋ>���s��R"�38���p��Ngdb�1�8g��*��gm��p��<�&�u�M.�C�e��[�&�c��\��gФ����F)O�HA�/���]͍���RB����j���ב-��C"f��ƻ�
�{��e�����CxywӍ�C�3�l�=ңjL	"}���^�����m�{jN^�%HQ�
!�~��4�$E���ͷ�_!�LZ����"U1�1\�}Id�u�g
Ls3���%0lDn�ʣ	�[�c��Z�I5+��h┬��qEj�N���Of�nU����¿8e���S�.��vϝ�0!�꬗�N���b[��#���	����heځ`@�g�Q0�i��|U����v{��G�C����H�rs���N}�T>��T٫�y�*I3t�6��ݑMЉU}�1%ʩ�# g�J��+�9>Ɍ�1z�2�<�k=��lWO���W	�7e�t�7��78;/���
�o����*^6,X/�	���
��*�ET)��R���V1�n����Utnel��ןu�j˗�fmJ���+�̘y��r3d��7������R9ci)Ȩ�k*H��#y�*���A���`5���*��*��81�F���ĳp��tW=-�0J�y9Q��o��3'lN�����㏽�8�W���Rė����72�ޘ}��U��"G�/h�{2���6�w:��2��0ū��U���"��,bLnQ!\��m��m��r$b�Sb����<6�)9Z)GUnJ]�5���)�p+��*�yL\~��xK���N9X5^jY����V��u�9/�;]{
�"̨�^���
�
\(������ڍ�w/��^ʈNQ�ƻ����%��UңU�q��<A5�
�q�nC]�*��-�ÊRCو;*�]�;����wi�m�kW�M��e;aڷ��:�jB�[�m���[*&�ˣ�|��
�y�+z���ފ�.F�U۫w���PUN��
=;
��u��jUȲ�uϚtb�*5_p�(�*>JO>'��Y��A�3������9��NE��\k%���қ���l�'���崢���tP��f����W�7
e�HQP2���*N�g)����?`�z*�^��Ӂ}�WY��V�o-Ц4�+R=eW���q��^���U�1�i���զ�����A4e�v�[���^�f�S�r��g�.��(�N�<%]��_&H�.�O�+'{6 ��܆)F��8!���pۃ>�e��@Q�sA�s��衝B�P��UД��V�؞�n2�B��P8 6k�IU��|�]?��.�2ӻr5�j�-%�����x"�@����T�yW������]l����0��ןv�����:}|hLtuM2"�ޏR�2٣�A�`½�5i��Z���`��Gh�ȵ"I�ޑ&aȡ22%1je��(�	�PQѰԞ��w#aЧn; *�� J��	����;+���i��2"!K3���㘁Jll��kӲ�T�q�/����8�B�@Q�~���r'/mG�]�-�=,G�u�s��%}��q�ɡ�ן��s7�,G���������d�0bo�⛞��(a�s�|�
oiW*so�H�uS��1�Yץ{!{E`�R�Uo�TZ��de�v������0��W<��v ������%ҫ�Wt.N޾�K���p�?2�o%�O��vqM�<�H��K���sQ�9��������b15L~sp�)�d�S�EL�z�Ks`T�9^p!�5���J$�b��1vk�2���ƴ-��12Ue�U��zD�X���0B3Y����;sq�i��R��f��]�^���4n��]�)�Sw��7������%Rr0T�W46�}s�l9�WW@��c!7��E?]��z�X���  W\�5���;�A3�%EEӻ��k�B��tg�ĴQɮ�4��ʍMeO,��F-�P���oV��������ic��F@B���"�c�k�RV�ĩ1��vO�΅*:(��og�R.=�#i�'��M���-�U�|���h�l{�y���A�����LW���]ݹ�}6��|�ax(�#R3b�UB�P2��͗�]�g�*��@��3~�b�@}5AM@�X"ގpJ|�fY���c
�}�~D����_@��ѩF�Z�Kǲ��	mx��E�!�0˨��P�N��ݮH�II&ݐ�k�+d���7�lN��u�\����y|t��:�ggW��<�Z;e�skC�),���R�0���D�N�<z@rv���j3���Qκ��\�M5<b:�>�$e��!!�W�l �f����fױ��a��\�i�8�p��]����E{aCsШ$S���{��{�7�b��j<.⭧X���X$��Y7�n��ǚaP�3�T	�ˁ�T܎�>U�q[%ME��騹�IkK��ޥ^Z���3t��u<�L�
�""�{�{��<r��s\�c�t(�+�P5V��J(wǱ�ƴ`�Cxˮ�ő���u��\�r\z4��9���J���+�G��Y�����u�v�J/s���)�F��ڥet�
�ʡM��"?إc��'GZH�n)��>f�U�����h"�ӌQ����F��m�n�7�2�H�<3��a.�a�]Z*q�`<�#��G�gf��z[��e�������ҿx{�3�g�=���d��$a�+��36�GD�@�]g�Lh"��"�����.z:,dڑl���JE��1���J7
��{t�&�VB7���Fj��ίmӿL(I�q�fA�/�o֎��]^Է"�iS�3:8Z*�ʏċU����!�|=D� &���o� H�nz_�R�@�@p��3M��K� =��c.�(Ȇ�-(�l�n�N\�;�~*X�TH�/EzC����
a�HE����)�0t��{b�eD.>��#�\����%��Uҡ�H�.l��L�2(Ϙ�qA�b�E)Ѳ���za�@=C"�+��ص���^�0ś��#�p�h�9�x���(�.۞��EU��,!D���8���N�*_���Јi���yݺ��y���P���}��`�X�*�I�hhˬ�ޙ��Q�
_&���Bñ���5Nd"�8R6Z㡑(��{#�r	4/7%C�ЮP'|⶜[]i��V���"6��ptX��۝j��U�/i$��Pg߽��U���8!�ʑ�s9
�(�:�t	�l�u�ޒ�o Ñ�n�����L@��
+�^��8.K�,[1Yë/f�X�p����ω �G��U�M��2�z�;�]q��謻�M�ɨ�Mz��q��9M��V��E���`�92�F.�'t��c?L��YsB����2z(	���u�y,���o�K��TN��Ю���@́~R8M٥62}�-����y~�Rm��ʟrP�����=Z{��3�p��<�϶���|��s�ϋq�;6�-ϤZv&/��i��w����]P.�сPr]u=M��r��F�y����=��jD�d���tOl]���R��B�B��ca�#�t]��r��N� H
Dh�<|(� �O+��8�T���ӣc����i�����˙3s�Ԣj�CQ�Ò;���tXw&��=̍I�����!ݦ:��)hP[�/t;Iۜ;ƕ�ڊ}{}[z)KofY�ړ�UU���(�B��C�S0�ǬS����JvS�o�R�T�J�*"b��&��K�b�K��ȐҾ�TW�߇������*[5��w�+r������.��x`��Z,I������^�N�5�!ا�OE""Ȑ����>�4�]��\�=Ϳ�U"��S�s��_^{�%�m�Et�C�rT(�JL	�C��8K�"
Zר�������ެ��x�u6H�V��D6�t���+H��K۞�̳X�����9������5H�BT5��Vt�v{��9ʢ#���a��%1w�-��jb�`���eHW7� M�)�>i�Y7e��m�����y`[-�$
��pt�x8tRf���td@p(���H��лa�	�2�N�b"}Ck�!��)�@�Tc�݂q�]�����g�J��5�f
f��,sY����ٻmI{��^��������^�w�É�@�(��pot�D?��JˇKVr����E�_Bg�#�.��W��K�{Ê=�S��Q�sY>ؗ;����8���D���B��"��f��ʍw��!�E�o����糾r���O%)Q�>�5)fs/����L���z�u(�)�1�;	g��3��&���ceXq�oo)L0�6F�SٱR*�שˆ�a��T5�}H�����Qb��=BB���|>� ��B���=�^�υy��̧K��iNN���O�Z4�_����Lk��;bb��=A����VW��2�[��Rc�9
�B:L����W�l �k(}9-]���|�A_��f������\@�U�{�V��3iz���m��2���\��b㢜�P���U��	�A[���(��~^�|�vdkS���p4T���/.ې}С�C���
��/e�0�b���G���g:n��A��IwSa�2'n阱���:�t�8�A��i�A��3N��z+3�9�Y-F�fr���(8)�9��w��ڡd1Հ`���Q�'�L��a���Z��|U\hrE�F���%�	ak�4���b��]�7ēi�;ɱV���rk[touj�.�T��̮�.�����N�%j�We��k�B��խ���Y-�WK�r�P�Y�9L���!"�8e��hxw��cu>=W4i��5fu]vc?7!�{� ä=�y���B�穫�B���r�!���>I���"OM���wͽ�c�.Ɂpbx7YK��t�<�ӓMe���E�4p�8PtS��������pA�}n�:���~óu璘 �X]�Q;��R�2��5�����L��\B��;��lf���Bv+ `��Tl"h�w�<�Y�r-��j�,^�D�Ɂ}0�̼+~�e6xt�[�%�Z�U�TYe���/���u��D4XD��8v��
�W�T�v�usC)u%C?P�$��^����o:$�˥��WSq��dMT��Ɏm�[ʥ,�$c�/^_T��1a�@�s�Z�%�$�4��!FM�ł���BSCp#�<�ն!ʵ��e[�]ُc�w71��)����挥7�x�]�5a��KD�FK;YN���i�C~]̡��6���+Q�Agm�1�T��4�'���@A����2�^,LwgjV���Jd�O6
=:Nd򫥦�6>x񽷸��G���d����b��T�Ie9g��ĊK+/��\e_R�n�&wkw�i��Ĳ�VM�*�ǻ�i���p��]�9��9�0�T�1w�jl���aVs��p�K �A��th��;�!�����j�� �qj����,Ժ)�x�_a����Yzq�c��e�w˅4�#�We��@���ށ蛙ot%�d&㝱�Wc����&b���Z�k�۟7x����%�NG/y���cf�����	IJ�"�
�q\����{z�Z��[D,�1bV9�j��1��U&�)��p.�)*m�����e���T1֡�Qu�R�ʎ��e�+�����ҁ�jы3n%LTY���r�r�P��fep��q��*Ki��]7&�YZ�-J�)��
T���Z���e�i�c.��L���ܛ�DRL�Tę�b�em�q��Wr�[q*j��7l��b�svƹ��mq�e�ŕ&[v�i�q1dm�MM��ډZº0�WQ�c*
:�P�C6�w1���a��LF����ܵY����2�6�F�V.#u7(c%��ێcmMTm�ۭ�R�4�q-��ML�-e5�Y�f˩�Y][��C.9o�����������s�=mq�c@�B\囹��LoX=bf�X9RY�Tv]F�ໄ��
~�}�W��[x'��z%
YP�E��98*v��� f��"�x�5C$Y߫Vf��� ���P���m?)Eb��_�`S�tM�Ⱥ�w�x��ݗ�=�{�����aa��]*�Y@��&�c��:�M	蚆�a_���:f�v(DڥƑ���#}`eP������)����:T�����P��1'�VO|��La���R
~|d����۩'�=�S�N9�C�1�z½�jc?rɌ񒸆�s���>������>�QH(
)=VT���z�V}�<g�P�_�0�I��v���q��$;gLǉ�& /ܸ��+��S�=�>y�3�����x��&�2
Ì+'�m ��O��UH,�dRq�8�_i
��tu��
A&0�j�:�&2q�':��A��R>�����7�^��֣�# xD|���?3��bB��T��٩=B�7ۖ�a�
��?0+8�����J�AIP{� �HW�>����H������}���;���w��8��t�iR�~�>�R�?}���m�$��H,���R
i����*�&[>d��3
C��d�%@QO=������^l�;Om5Ȩ�~��@����}1 T�v���)�<a_�:L�B��J�1��E ���`jO�����R�*�큉��表
)3��ã�`xǷ��\�W}:��ߘ2����]l̑���L󐤝���+3t�c�ɖ9*שR ā��+2u��͝-
��F˻��B�GKG*�j�3c�ʺZEޝ{�F��\������={����@����
���N0�ܤ����E�W���Y�O��<@�0�>���Y���j��v�I���,t��dxLxTE�s��������_�� �q+1���
/��>eC�)�5 ��X�S���>B�yd�R(��*|ϼ�ԕ
��/(�V0��p�������s��.{�u���{���=@Qq��5 ����i
�wC��Rz�g[d�t��u�1�����k� ��:�~O�>����LH,�r�E��Q�ٿ|�f ���`|� �3��à��*Ad�,�q��)����4�:CS�O��ó����~d�jAgL��d�~��Y�%O8����=�t��{�E��~e��	���� �i�>CP��La�
�_�l1TY�
�SӪ)1�8Ɍ1�:I]I�ğ�&<���c��1�c�cǟ����|~��ӭ�~g��5U@�*AI�>q��:�*��8��
O׬
�a��������ă��b�OXc&ͳq
�ܲy�o]���gy�wώ��(��O�����V���(�V��tԂ�w�<d����R
L�޴9� �@��a��L<�O�W��gc�l��R
N^�׿~G�������辰_��^����1:���Y�Y��M��Cԕ'h~�p��2b~��XjAa��c<d�f`�;q �<V<��c�ȥ>�n6v��e��b߼b��0�)��0�r��Or�At�z��m�{�+]?f����Y���� V0�;������^Y�x¤;��>��z��>7z�~I_��Ϲ�E�W��$�
�a���V0�09���rɈ
�O��'�g�R��!�=MH(vwI��Ld���Pb�/�3��3�>�]���rȸ�Ȗ��БS�^zo��~���W����i�`�I�s���3x77f����i� �K�2_�YF�O�)(��w�r*'/^R�N�k��k������_��<��>	�Ad��]C��1 �N��!��:N0�}�I���[5 ��<�T
��+?yd�h�V~7!��&�Mg*At��@�xDz�'뛯���sI(~p���$����˩�I돌>C
�s!������_h��}���R
xyUI��Xb$�<��TS�ޡ��*cW�k�s�O|���$R�?0��!�ԝ2z��?RN�q�!�$��a�N2�Xx��I�uV��}o����s�ܜeg�bC附0����5 ��|��Y���b����&yHT<I]O2Ȥ�
ϙ�C��a
��u=��ZA�2V�}}z����y�]yό��$��.�l��
�S
T
����?}I��7욇����䕋58��tI����^�~H,5����������{�;��7���g��H.0�(,���v��
�]冡��A�Si5�a�Ry�H,ĝ���>B��ݓ�X/�~��e�jc��ĔG{19�v������}U�ҐY�ܒ��J÷�bA�f���~a� �l��Vx�S�N�I�T��O̝}��HV¿��$�?$"=q�f�9y|{�OѿT\{�G���}I'ʞ8�m!S�vz�jAa�ϙ�1���1 ��=�N!R��,1q�`�P���'{���
$�:>����]{������+>�쓟����(jC�`l<��̕�����Ă�S�q��v��k3��N\H,���y@Ă���T��
�{����lGPSӷ�/��{ݒ�gi��)'�Va���'���[���I�u�5 �E���1 ��^Y5�2T��}`V��jO�{����P5���=���߻����3gb�@W���X�o��ŁN��K����z	��Ly�����4��vEj����b���2���vP:�䛰�	}N��mI-<3���־yfj�B@�	#X�J��TR�3 q��*bꁩ�:��a�O��z�*�ZAC�+:���ԃ�gG�?0�@��Ă�̕�������s�����o�v�vɮ!ĕ'hT�>勿R�hz�Y51 �{dǌ�e1%H)8��dԃ�!F� �_���1���R���~0��޽��~����=B�����q�H����{�j$����@QB���`T���s�,�o0�CbC�I�T1��T�j�R
|������wwy�7�{��xE���1�����Y�>O�����2���a߻�߬��1<g��%B��VL@QgfQa��I���ԃ�K�n<xL��݊��7������WG��x�P��d���I�s,|�+a̧gT>CR8�r��>J�'�fE��X/�\�tLg��a��FXc=T�����~�:��>;�� ��J�NX|��Y�,���'�PĂ�Ri������'��y�7��a�w�5�����2W�M�)�@R=��Ɔ_��qKྈ���>��O�<>��T����3�1�a����5'�T��?Xq�"�XW����v��Nt}�~@QC��z`T�2�f=�{�U��YN��H�l�����LK
�ĆZO�1��VEUR
Cy�J�8�~� cY�c��5��b�C�d����1��dϬ��?'���䂓��6���O?k�9{����ӯ���Ɉ
/ǿ`~a�<@�z�CQC�r���
��\k��J�i_
���u�M�����?0�y�O��=T����#�wn�7F9��|Ӟ�£����I��ԃ��fX}�H,��Lgʒ��*)
���=B��;�ɬ=aP��LH,������ud��&�+���үz��`��i�K�u��v�Pos�ͣY]gv=��7U6�ͺ1Deq\4�n��m1,n�s��Ạ�o����eoKS��,@@m��u^�4���*d+C��?�����梜l}�\fH���a����;eed�>�y=� �����}�}��T*�S?3͞`�AfwE�$�
�Xrd�8�pװ��T�$�\����$:I_�xtɈ
(~��`T��uf���g2^�aXT�֜@�����,�T�ɇ��ԜgHty���l��z�R13;�����{������E�Y=eC���~�3�%bκ��5 ����yd��1�O�+��bA��y�&��+&yf>�+1&��~@Q}|��Ӫ�l���-�:� �����!X~O���'���;Iۉ=J�:�&08�~�� �@���?0��H*�Y꤬�¢�P�y���@ꅰ�]��Omw͎�:}�&0���$c�L@QJ��Rt���VOsܐ��l톼d�1�A���+�N������a8���?ud��'\{﯋߽_�������Y�58����_�����-#�a��^���
�;����Sz��`T4�t���O��'��0�:�t��Y*Zʴ,%_I]�#�_��""�G��O�I�;q������3��
Ae<��É��N���vʆ��ѴR,���E8�R
"�frɉ1*,1�O�/�s������=��p��$�
�z��f�8¡�������و
/�Ϸ)5r���gt�`��m'�{Lgx�MJ��C�Q{B��39��/:>~�3�{ﾝpS��a�jAg%~�d�R
�&$�
���g�|Ɍ=C�
AN���j�q�!�'�f���9�B����S~��=ϼ�]}��}'l钸���;E �e���eH?]�Xx�Vo�LH,��?}��E���0�I��u`g�Xb)��H(x��׈�ި DUr0�ب=^{���N�@�;�X��t���6Ի:�b}/쌯�/��{��9�0��O��p��e�Q<wq�
���B�d�+�=�Z�����S��-��x{�{X{�b��@5%|`T�P�gl��d:����}��Ag��spU �dRq�8�v�=�+Y��0��R���8��Y�l���T8���k-��~�;�ǟ$�T�Y�x��׹!��m��{Ca�*c=�Rz�`z�E��N�@��g��j��&��������w�w���q�#� ��d�L�'�$�^��bA`q��C����s���a�:�H,��=����S�RT�!P�%�_|�<�1�NWݥ|*�8]"�N98:�N\�;�~����*$ExȍS���<��D��b�D)jT
���{b�b�ƌW��Vׅl��FGzֻ4��I*�'�Ԩ��??����J��՟����#e�ۍ׫�9�TS��\��kҹR�5�*޿���y|��W
Q/xة\R�n�Z��NU��/+^�(�
ZD4!�;�Տ;�V'y}s�}k����/<�vp��1ck�!��D'�*d�����Z5t�a�r���]̦$�0a��u��'�!�����z��YU����Y�K'�rM�Ayyq�r�È����p^�F���+��Uc3u?���i� UKu8(�h}�����K7L�M�,���;7����q����|�dΕ|���1f�h�z��W�xx ��)�f3*�1]={n��>9R�3O(W�N��il��y9J�f�R��@�pK�ː�&�Y*6��9K2lwU�1�{�Rj����ޤ��o�Z�W+P��A����)�s쎍Ρgn���0D��x�b�a��:j��ߍtM]�@HrK��VM��7�K69�\eN�s�YEHMе.f�J^����";EPT�G��YY���(�&rhm�[���3|�Չؘ�d��ȯOz|��
�n�h֪f��P�X�p(\�Q��n�r�v���܋
D0bn�wh����12:)��79�:.č�T��aV��ޭ�vu��r"|�@$,ҢG��{�}�
\lx/f��3�{G�a��&:�dК��lD
U�;*�Ms�7��ۮ���A�u��ʓ�m�P Y��o\���ڞ�7����n�<��U�3��<�6:����"��"p��Օ;��������))�{�M�֚Vx�[��Ғ(U�2�u�K9}��{����s)�Tl��;G�P�௕D��B��]	G�� *:!��E��:hDN�B��)��I�Ȑ�}!��]M^DsiH�Bٸc[���㢠��P�	��� ���T���7���R�c�`�N��	y}�/�YC-��X�^5�aZj��'/�)�;�����lHtE&xW�f��Hm
b�mڬ�PMଟ_��ġ�6n���Q<$�t�H3����2�uӫ��@��hv��-��}�@n�jl���-��  ����/4U��@��u!�Ns;IQq�!t׶E7���g�i��p�����Z�>Mg٣���.0�o6;��A�crk���qPV�����$l��$t��R�R�<h��D&C��<4c�A���u�-h��Fg�(%���S�9X}%9S��x<Ƶ�W��;O"H�$'Oi��
�� ҕ���F�n�HF��(�XXIEК2��Z1�ųA2��ԧT���(�gW����sWǋb���_Q��Ê��}�ܝ^ߒ�Pfp��/�]�{������B�>
��<G�kKl�i!�����V|)�&�S7�,NfJ]ɠhSt�}c�ۄ�H�*AW4!�L�C^HkFiէ�^���o@nzt�St�����>�5葂�)��C�m싅vh�2���mۉtu� {�G��Y�WP�H�Jvו��T^�(a�"�B��.}{52[���iR�Z,hh�}�B9��y�z����_�px4X��Uc�q�
+kd��r�@�ˉ|�˯d31:+���n�
#���>~�+h~���Π���N{7���~(:�TV/��J�#����$X����\�x
����;hz����Q�T�-4�в4������ӿP��v��u��+y����5� �R�����R�3;��XB�%q�V�F�,�O5��Ԃ�t4�Ө)\P��$�:�/x
�!��L%�[\��td�CU���< ���1&,\(�
2OG��~�UlUϔ�*a@
�G,,��NT�����hε~��鼫Fˆ��(W #��r�`5�ɒ���J�u!��H�@�Sݵ�ί�L�)]Su�$���B�a
�p6d�� з~��.hȰPN����f�u��m܆t�#��"60p�ԫ�Rǃ��>;�~�.S
�=�8喢�tt7#q;ʓbt���.�yА5C�Z���c/8��c�F�'��@q�}��u<�@�h	$O�Þ�W���J5y�6�R��0�9y���r��;�R��!����p�|PB<�D@�-ɁnS��lU���4b��W�Ѭa,=2���dW�}��֚S�&9H����ˋRCޠ��j��!βn�2����� <�AV�g{g���]֧W�۷m�<TGt����$e�L��X��K5SJ�tηI�|��
'2�����Xj��ȝ�:��j]�A}����j���Z챦�s��0�N�-�w���MCs�Ƕ�6v��euf`kT��
��C�xF5��=�E�N����r슔�����QT`�
�E�`����u����͈e1=Y���,�^�6�Eo�8h�zP9	�`q���5���D*�l=���ﻬ��k�J�W���'V�,��eq�;3��v������}Y1Z�WM^d!oK�U��7�PfU��;��Ҹ�7#\��V�WR�!�w#�\;��g�k��-A�ء�x(Ȗk���X�NI;t�4M������6�W�`��*������|���d�]�]{Ʈ�N�Z0ܽ����٦%�Bt"�%���md�)�v��pK��-`�wsE��Y�#H��k�LJ��:<���_M�j|��e���=2��4�u��K�0T$���=�o�wo��LU�Q�tvBq����)�v�U�7���L��\�2�9ےrt��-�4�	��2h@d�C����\���̴a��[ُ�]�Lix�.ه"Ni�B��*΢uo���T�jn^Å귕2N��3T�E3Q�|�Ve��M] ��Ze"=��ɽ�+ ^��#�f�GY��T��yE.]iY���l7�;HL=\OJhw`+�f�e�>�I�����J&e�{ȊP�v�B+��<3'cS\���������hm�g5��ځ�5x�L�O�NƳn�t�;Y�>+�j����2�ԭ�Tn��ZA�)'�[���A(v[o�o�*"����n쾳��V�'Z���*���dBR+K�MpգHy�Gul�M����0���t������L�E<�A� ��;�]NW��J�����`�Z'V�[�4�U���N��b�C�Ԙ���Qۏw!��|2�#Ot���e
*m\�.����bR���/�Tᢴ�#���\��՛S5�t��U�e�+��r��PF���-���6�0-�ָ��MCV�Q�V�1lR2>,��LU0(��%��e��nn�Tۊaq�rnSLh��n幆��1�������p.�nij�]w\����[Ac�*�s�ۥ(�r6��ۗ6��
f�`�n��۴�(,�U-���6�C뙙+tsܺ�����V�(빎�r�ʷ.:�u�SWQ�b�n&74�\�\����3sm�f�2�8���S[�EUp����r��˗*#���n��n\w-�\(��������m]���v�pۍvَ���U��\̦[�D7+eR����F�бSpݮҍ���]�v���˥ʤLs�ۮf\[iX��ˮm-�drű��6���n镹q���9q�n�e����s5°K3
8Z�nmL3[
Zc1�r���K��6��c��o���u_��5�jMPȮ������9Eb>v�R�[��� �i�)��G&`t.�OH�h��[f�L^��W��n��q��xfkq��A�
�\g(�*0�]��+��;w{��G'>��e}!�ޡ�~U��`�O�*P�)��j�m�wi"����2����ѱq�FE�58ww��re1�JX�Qn���6��A�>�+4'����������{=G��>��S�P��W�xJ�k8��/�a��+`M5�j|_.�^Hm��󞉡#8uB�D8��h8.}�=z+��\��E����ttʄ��P؛4 ����t9�Tk��`���/g��5y��,'\>��(�+���^�+�@z�8��B�O���;;v��'�ǟ��C��M}/��f���/���'&�E{��c4����RS.���j��,]��V ���\�
��ݻzbPdS e���׌�*
��۷S9T��Yuo{:�.��2�1�\ Nh��	�����,^��U� ��޾���1��k`\���G�I�[��A��DK���T�K�3�FHs#"��GF9p��H��Μv�r(F4�0���^�2 �) u���Bf�s�ND��\[��5E��՝�Ғ�lHp���+E@z����TU;~br�9�ȧ[��K�=(@l
���#��,�����P�U�|���Ȩm���#�B�B"u
Ҕ��t�H�@ƺ�6]�5r��(8���^̡{���U`�����{�EO'�ҍps'v����G��{������%��YA}�v�^5��ȞΊ�x�{��&s���:ã8�o��w��)ѷ�5��gK��J(gn�x˱��N*�0P�t�L!�m{ƥ#EyU��� v��U;6��cB�j�.m��;S�;�Vu��a�ʎk�H�F�T��t�n��_�;Qu�>�r���F��Wvk�/���q�ӻ��ul��N�kkf���K����k)��l����}y9���-�o����pj׃�p.�K#0��K���t ��V$j�sY6��%�LK�^Uخ1C�"w�K ��7�R��U�(_Q�F��P��JoUa���p4)3�U7!n[U{�0���P�S!E#�֯�#ݹ^:6
9�	n��o��l��C��O� �r�؝d�=��{w,�u�r����H�~�bFr�t��4R�A٨�30z��8�V�Kl�iW�<<W�p�g�h��.;�5A>�3�J��)$ъ3����pb��<���k�M����
���K��@5葂�{���p-{����B�ی�.�b!0���JU��{HV����Ewr9$\c�ue{�q���x!�~vP���O�ഋU"��<ռ���CW��x0��i�)�WU�sz� 7g� ��Gr��͊o���+q
t����aK]Ķ�\�γ��.��#�h�q��aX���4J�m)!x�⎭��Kd�򪇽�9���غ�5*�}������U�t�x.4�C�٭X��'>m���M������w�DFl���J"7e��q�>��� ���Q��orpsԤ1���n����J4��㡨�,vT���ާ�t��~��AZ
��n�E+5��4C�QA�L��,^cf�;���G�p�I���i_�NE)�$*	�͎5��Qlh��0&����c������"&�(�M#5N��ps���Š=B���|H��)���\7�2�Q��׋~�@g�ɀ��~���'��gׂ��Ex(2D`rw뎁�按v�&��+Z���[t܋.�db��6"v+��s�pK��ј��]*�[�E��z���5����N�h�@駄
���������g�%&�wĕj�nQ�P��[F�]Õ�2:e��#+�ĭ�tp���NG11�j4�Wg�z��V�!��S���#v;]��i#���
���s������ bI�R?L�cᗶ�._J��81��^:�R O�<$X�'L.wy���I~����NqJή��Q��S�QT��eD��/Aڈ���̱:!!^�.*dFˇ-�s�=�T2�r̘�!ti�����_xt@���*<V���TSU�.σ��4�=�J����.N�˙�⽪�8j�V�~~;7S������w�*��Q�=r܆ 
&l�!G����H��&���J�P(�6Z�#a��~�vk�ܢ*�&�ޡX3>w@���ʳ;Ń�ƺ��k�#F��@1�7dt��y;4�"ʎTy)u<%�M!�EZb��j�^�u5US��t��B��M�L��#�����rdײe��6������5|u�|�5���[	ـk˗Y���Lq�N3��ܹjo^�n��qv�e�M����}g���DvT��ߛ�(�xr�s��R�3��J:���[��x 9��-��1��`f����OX���}BeǶD�r\�!96E�{������
���êp��UCbL�"r27��u�.GR������S���TO���QxW?s�q�y(Q�a�"3���s;*-�P�l*q�����&���Pflw����Y��G"��P�#�D��H/_����`�p*�tQ��@�'�l;;`���7���Ƹ=���<"�s������򙏸v�/r�;�n��n�4/z�洇M�[�V`X� (B�jh�����>�{���ֲz��e�GE^�
�LE�4&�{1V��P��В3�Fi-�Zq�5\~`i��^�>��8/��*����>5��k�ln䎗z�@�Օ�P��W�܍�
�SʻVRB@��t��պ��)"Cj����4�gP�p#QL��ļ���g/@#���N]�1to?c�S8�N�nz�Ԡ_w��H�eeѓ����{�kkL��r�	�faͦ%@;UQ6E
Է������{:���ax�O������\��U�����Vj���Nױb@c�w��yH�x��4:%�΋��z�\\�t���W
'`�;�X�7�
^��YF���8}d�,{Ƙځp
��W	jH�::ۼ��T_���%]-F����Ԥh�*����}��st��Ó�{>tW�oa���k��עf hЩE�Ӊ���5%V���V@aH�7$>�E>�0l�Qc�(��b"�ϲ劻yg_�,h��J��!�����Jlj��4��p.���p�\Y����-�B��"C�t[���O�'�gC�����KL��N��o^"?UЩ�]A[���Ҵ(9�#�ʄ�)����jl��J[�-�-����LA�f\ϦO�65{�8q!o������4�P}�gc�͸*���X���+��V�]x��
��r��I̝���d��j͝V�DhF4l�.�2���֩w�c;��nA��1	P�ö�b��OϾ�꯺����d�t(����9�UNR H4b��t ���FΡB��Y(#U)�p�p6��H��,G>�5��=���N�v$�}0&�V���!�߼6��¢��VtQ Sx�j��p���4$Hs] �P�j}{5�=QD_�@����q\ػ[ˈ����<5)?s���\j<.��ҋ6��6{=����T���� ���R�Dݟ
#����^�����0��i*8p��ΆPP��g��Muz'�R�h��������K�'(;?{�]t>�c��UO��X(�f�#O΁Ok�q�l98�V*:@��
2H�_�*�*<�J�dE�+|��Ĩ!���.��<���2�i��ܫʴ*�ب�T��i1ok\�O��� �ǵ!�f��h>��m8�:cv�B�K�\��㸖Xm�E�-Iղ��k�G�������2j��f��2��ZZ�It��:�K#W\W�Z��U��W�{����a���s�z%�R�>�T)�s� _O��a���̶�L����U0Z/N�~b�U����~_G=p�x�$E���FL셒EH���Qs'�v8@�>D�&��>��ev�6���0�ߦ5!F�2'yS�ED�4$t���r��}r�wEL��lq��>��:ո�].�C��m���R I�8d��i���Ի�`ja�]W�l��r��]'.zӿ. ���e��ĈaȉB�*v")0`R��z=�U���4cokqeX�lt���{Hρ�i֕��8L򢩪�g���㯙�n�_��b����vL�Q�}8:��F�p�͛�����X�j2(	hީΐ�	6T
���(� ��|+~�~�C5b�@�kCĎ����ъ��aXqǣv�UiJ|,X}�3��Ji�Lqt�|F[H�s�I�BK�Υ�a�+uh�O/h���X�S�<9H}ąɒ*�t6�Oʪ���+uqL�WPȳ��ˊ7X���
�W���*j�`v�������͂1u!Eت��dn�~�zA�ٸ�ѿdI�|5e³9�YB�D!?O�fa�*�L`�B�^{(�>�#"G�mc���1�T9��6n3eL׈�����5��_*���x�z�ʐW%�pؾ��*�5�b7���U�~��!V5S*��5	9}��{�����l(iy۫%BS�U�2# "�6%��@e��n�e3���l��cbL�yvR�����P�|Ո
�Eb\�(%=���"1�s�F=fG�Hʷ/���Ջ��sG�Q����ʥ�QlU��O���Mt�Р<�-O�a��h랭��e��B�Q��Ŏ��R(L��ET*�nzEFCtZ��0�QmA#��n�Mp�IK�.mK����1�gn�@8�x�u�aG�(�t�[J�^J����o�Mծ�);�ӭ{�m��U������[�,�е�+�g3�ʡj�}bp��kK�R��.a�b��L����ebR᜶K!�'��C�9�adt	c�f����5E�+�G���Վt[��3,6����)S�n���0=�}�fA/��(�2�"��]�a�s��m�O�E�skVs�l#p=3�7wwe7y{���QћVmL��/w�ZI���Q�����7k���{i�r�賮e�
K�ܹ��!���2��'6i
�8��>6V�p�6�MY6�&�`��-�����O���Y���3nI��kx=�Jdunp��J��	u� �mR�Gb\�kZ�Mʉ�lρM5yD��0rU�y4	Δ���w�aE0:�JXv������e���e[����A[�.F>�J��M�$��2�0u	�f���^9A�0���R>F@P�4���\8��ힵ���c.�fK$uJx�Y�teމ��h��<yI]aԛ�4��w���:T̃_o�4F�ޫJ��7�1���[�}}S�.��cN;u`�/�<W��g2%��g>�
�c؏��ѵ��̚�W��)�f�Q�n^䔩�H�'X���;mݕFR;K�B��Th�R��u�͚����`��hj�Zע��w��W�8������OavR[�^D�+z�Vތ"� wE=s�LX�bβo�}� w�<��ꔞ��s9��_>�3����͡	�h�r�esPa�V0ù7 K�q
RK�B4�$�UhT��<hZnE��%r�<Q��+�X���d��F��C��X'Z�� #�4�9�[r���lk����j� gG١V+���麗([��j
@�[��Y��̦�,���\��E���j��,�֙��j��c����w���̷�t�MW,�ŽΙR0ҩ:�-[��j4�Q���T;�q�=�o�KJ�ݕM��\��%�k�t��=m�\�Lvfa��R�"ٻ��V"�*��2�\2�e���j)E32�Tm,r�a�&fdʙ�\�ݖ�fe�e-)�f�.Vj�h�Db���L����̙b��V��Sw7kJ�U��0�8ѹ�,W0��ҫ-i�;����8婶��j�f��v��S6��b��-L�r��j��)lieݣ�p��bۅn5+�&+����c�%eE��#��4�̶am�nUV�7\QU��[Z�qȡZ���\T�sq��QK2ܴ�һ�aEYQ��ۗ����70�-l��P\(ڭ�M��eb�ZTE�.-��[��%�i�0�Z�B��܍�k��m,��ef%q�aD�У�r��3+h�X��Y��s���(S;���br��Q�<c��� y)HG�k�Զ�ۤS\��\�)�M#y��)f�q�<<<;)�%8>��n�8�p8@��Z�4�W������G=�����	Q�_��Z�~��T�H�!@؈1o��T9���^U�S���тXn�z�uz�aJf����0�P�;]�H����&nΞLMԄ�qQ�uJx���U}F�f.��P�����]-e�k�ء�B��������A�^RuY�!v��T1��)=]�8(2��W	q�g #���}v��2���Gm�U���2�:�S���(��nqDʺ5j�p�L��	ƽ�Z�P���&K�r�4�5cD7#_UTh��ji�B��h3B���g^\�|h�����,I�-� O�uJ�#�ߧ�,N��|5!ƖR\�q4�y�)���!�p*�����ʁ'�l��.0�b��'��Y�" 0�f�o״%̤D�����6�6��d����[��f�^��"�<}B3��d��gW�hp�M����D���t���P'�fd^\�w�(陼0�h��h.6���=�z/�������HB��U�`(=�b��6;�+,p%�lUe��۲�1�,�nC�C�d�+� �� ջ�d��+�e��I�TI�غ��e�����ԁ�������	���x���4�t�r�b�\J㕸������~tk<]e�E�ЇՇ�¸��t�$��+�e�"�l0��g�zuA�s��Wn�@��ъ3`�t��Js�I�ˆ���*�l���Eԍst݋*��
}Mz;�hf)<,���Q���P/5[��<�Cs`.��4��w�f��I
�f[�D�BB�rRU�P����i��{q��1s�"�_�@,C��sѕ7�*�
�ę`�*?s�<uP��ae{���jԻ���W�����_h��D*����aQ�]*��
'3�x�kFqG�v�[��k؊�[��>�]Y8��S��2%ۡ�t/�o�V�� �=��W��ܥ���r��C+��p̲7�}gY��������J9����hq��{��-�S���#��h��1�6��㸾R� ��a���lQW$�o�.����߲�� �mX�"����0����f͖��;ɋ����j��X/TQxxX�8>�}>�*qm��,_�!�4��EG*���ݗ~��],�BS��_P����d���=3�%��A��sA�sݴw��,��Pw=h�C5\�DGFT�3�4�l�����*�~��*7T�e&�q�7!�5�3�.�jE���)�3�&�v8@�>�B�r��|^wno��лަ���^=<���q����i	"E���
�f��}���c�|�:&���N�*˄.F��g�C�R�@�][��]̱P�%Ll�ϭʀɆ'���Z60x�}c�n���93�m= 	oE��V���A�d�^�v|s��'e��ҬU�-���w̻�+���zgQq���Y�$L3\�=NP�L�R֫3��
��+�)�h]�o� xU�=�1W]ؑ
^���^:)|�{��.uV�������ǽ����S
F(�Φ:NOO�f��BnCRv��u
{m�+���zc���F�� W	|�*�hYF�b�bћ*��3W��]��XIB:3ҕ/ٶ��5ԍP�=B�Z�3�>��D<��Q����r�G�yJ��~�=n�۔��n���A�V �9�9��L���W�G�-��U��e�b��F�04lg*�΍��!�M��\n�P&d�����R<F�A?yӇh[�\f/�
�r�{�:�<�s���V7�����2D{0���-΁rD� ����y[�{�޽�lD>�R
�fT �O�qXڑ�0��;N=�q�~��9qu���f~�<`�֪��\;��U`��X�וe}m��V��J���somQJ�5oE
u�1�Vv����|u%����&��(`�nE۬�����
縤�v4`EŲ�����Yo��a��B�ky-\�����$?�W����ۼJc�����`%X؞���+�Z����:��Y^�����^}+�x��r>�b6�S�{�F/��+V��f��W��}����5D�W{�ؙ�4�����\��)�
�R��C���ٝ|'	�{�o9&��B���,ˉ�
TP>�*aȩ�vn�UT:8nc����<L�#���m�F��j=�2b�H4D{!G�fA����i���0�sceŬ7�!�KT�2�����ܸ0F������9FK}BmWG�hu�0��V�8}C�4uf�Uow�͑�1Lz�����箆�u����~�NE��:4"$j;�)Z2�A1����^{���m�����
r�����0�T���6u�-qǧ.��U	a;&s�EL�zo�(�3��8��~ɖ� �	Vx���-�,3�D)ʪ�^��>�[��Y�1����2	�[�\|�<D�ӑ��g�e���h))�=�9��Vj�<@H�IreD��̛nB��UU��̧���"�B���`WML�MZ�^����L�Ǽk������]���qU�F����y�>�����E@���vB4,��smL��w�"=��GK�"M��+UtQ��L�m$�#3��4؛�d�����[B����6	|�K��Wz��ke����R'T�H�B�`Z��RF*�S�!B����z��%�wH�jB�L��8L��2�rz��d{�ex��r��<�.�nT(v]�\xZ4�X5�k�PTMw��~׊��Z�ܥ��4Ӌ�6*6j��k�<�u�Ӣ����\Oa5��7�3<����Ϯ'%EB�K��c�%T�yH���Sn�^:$��G�����n)�:��6�:�]H�2���J}T�ۢM��Җ3O=w�D�Q��ך��И�����<��'���DM�u����Nc�g��Z}A���8攷^��MW��o`j�48Z3�Ѷ^ɓM�F�M�B+���=���b�ت�!&{�����N	띈���؇#���{)���w�:L�>�Ed�(Cs��jpl����!�L�Eu1(�fo�x�©Vhhأt~��P�S�*ڿ8�"E��=@��*�|�C�ƽJ� k��g"Շ�"v4L�ˁ1nb6	7�
!R|���a�]#=���#�SPL�w�^�(�!~h��M/t��F�~���H �XV,ȥ"��@���/���ē������{к��s�W�Uu��`��W�to2�擏�B�.���Q��ʖ�\Z4��)��bY��ʃ��w���'�>�ش������K8�(UC�����	��2�x�+(��+��R��O��}���3S~3�4�mzC��TD8
z �
�����5h�����8�.Cy�/Y���!������׺�y�c�O"�d�&�N>�|Ľ��j�cu��9Pn�1K�
f�3��(m-����s\��ݣ+�i|<< �ӛ�91���2/&����5!�1jO�rd؉����ut��(>\�48d5.�P�w멥/H���O���"D±�avi|�;6�꼪C��*u�P�\Tr��vn�j��ng
��Ibh@n���f��X2c�dÍr�4`��z�%�w�ns�������(Q"7�H��_hY48�h����>����;��ǺҞ��%��t���i���14��1��>^�Ǽϫ��QNK7Y��rbԁ�A�3Ej�OI�p�W�SmV�IO��b�VϦ����۞���(@��JrzA����Ch۬��I0�C)�e�F�ݱ�~ğ���VX����o���>�
�ϼ�̷w�ީԉ�E{(��@�*��2��,��[�#����n����=�8PQ��1Pi��C�_��1F.Kz��f�#����{�M�C�"�p�2�
c\շ��k��;IT�$�MJq2fo!�����f�� k�q��?Ͼ����w$�u�(���S5�FП4*TZ˿T[t7$�ݐ��ӳe��������^�N �wh����*q��b�pʢ����W�z�_�¢	� �)%[f��Gl�*�L�8����¢�k�C�E�4+�t�!�����̨&R��������$6�E��҆:�'����f�r=+FZ����:��<s�����ۼ��+~�-
�
��R�:1�F/ߕ{V�}A���W�clN�ޜ�R����7=�OW���R�T�.'�T��rɏj��.����e�Sn�N
�,[�q�(A~wL���s)^����5Wl��⣺_���9^F��%N<��G U""6f{����<�d���=f 36ʋf�;!�K�Uk� h=�5M�(3��*���{R*n�4׮�]n����s�
�ٻ�A��u���W��v]�-�t���o�Qj�����7�!���]1�Z��wX�t�o�V֙����}��f�2��B�aO�P���סרdÖ���z��["�mvV'tx��M,�^����V��&5J���x@��cP���8=��Xz�\����1떯�(ׇ�=�cd�S�pp�XB�;�$H7����({��t 4�ٟ*�L�K��?�K�/�Ƴ"�_m_2\v�ú��)�q'(�����6��]g�th�^H����1�(;"�^9B��P�k�デ�:x�QN*�m�9z>��2��;�Ҝ�EW�Q��uQ�_���>����裃o�S�J4F���U�_��55�RX��C��1�#B��eQ#`�xu1et���`�|�P�(n+)+ϖ
��8��b�c�^��-������;���`��S(@��DS�hw�~��Z����?�:nxVe��̣X���b�됥�u걧9��Eػ�6�6P@�}�e�EL�s��/#�n;T�T���\�:�#5��IK��7Yyx��0�*[��qR�V)
;��0����M]d&pN�������XY�k�sA����4�u����\�`p��#���$�Kf^�����Q�_Z��.5!,0y��X�:e�m��s<�Ų�7�Bf�ͱ��Y��a�/P3_1�%˫HDmn����\�Ht�c)�C5�2�Y9�t�Ց��c��s���^��5����	�/|��x�9�2�}G_Y�f�`|U�R7ܑ��ƒwX:mǆN]��`(��d}�9���Z��N/�-�WΚ�Еd�^^���zsF����� 8Hu�J�])V����|nt��AB
9x��^9�u�(�	;�4�TT)sJ�"n�ww���~����+bd�F�a]�15��_�a��թL�W+�`�i�tC:�5��y���*�إ�vR'o/�Z�O]�R���@�]��\�>�Z�
�t9/0�gD�9(��t"Pt��D>��p-q�i�f�@H�}Y[F��ك	��Rm��!ۜ�T/Z�T}Gx�+��5ult3c�w	�J'�PU��m��2���@�x1Q��6����!�g2re�.����}ZW<�[�{0�Ot�@�-��tLYh� i�K��+� �,{�f%��!��ʇ�/��B�l��na�p>륖9Kz��xs��E�{�;���$c�X;\�؞p: �`Ui�++A��ov��u�@����T�	�0�z�m[�q���J���Д�%uO�����֗	�R�#�v1ZǨ
��mC֖�ۓ�0�Z͵���y I틨�)-o"N�����9[-O]���.��Q^lU
x:>�U�+�3i޼z��ј�*%�����A[Zѳ-�C\ԍm�gNCHz��	��vtʺ�j�<�2�(D���X�BJ�ve��t�B1��~
V*(��=�uAґ\��m�A��Uqh�-�+�6��2�3.��Y�⩎���C-ZW3�he�̷s2c�Pm��r��u��F��bV囷n���n�3&5Vգ(�Z�v��L�WS���]�2KL�7i5��U�1Ƣ�i��.\pb��1&��0ܸnѻ�w2�t�ɗ�ݺ��`��nWݸ).�(�S��Ě�+���2�券Z��FZ�+��J,�����X�jۮGv�70�Uݻ�Z�c��,�(ۻs76�6ܚe�c��9��1����Q��╫nm�-˻�]�b�mLI[n�m�\V6�cT�#F�[3)��۸]ZѦ&�iM�n&��fj-.�t���������/�ۋ��Y���mj*Z�q�6.��
���_��'~BV�@u@�����ǥ��";T��-1�_^g ���ua��"pEb��Y��q���=��L(����R.����HEL���S�Ọ��9K�_5$74dl`�pۯwX�(u5��2b�åӀ�<�g���%��s0%�W�%K�*UA�5�}~J���|h���j��-��DÏ8ڪQNL]�u�,��c\���[��S'�8x�G��h^��CQ�
|`���N	���Cs`���Q�8#����J��E�3��� ĩ�W=����{l��j^�﷼7 C� j���xD]VK)|~���JA]vT�Xa�ONa�}֮�-@�u{P���u��Xx7�Ұ��>�Ê<x��4�5�,9�P�|�"��vБ�T�X&�=>��F����K���7
TOI�u;{.\�"��P`{�h�Ɛo��O%̊����F�lVxߕf@��Y��L3E^�$)��LI;�w]���yO�6=�g�w�gr�l��]9�I�!-��'�}#������'�׮�<�����u�6�I_{��9��%�dGΣg�D��:�Ƭ)�X�j��B�`�w���w�
��L�2�����o'�
E�&�ߪECx.�k&�/�*:������7{�[-p��A�y��X�\p��<���B.<s�4#M�3��K��v�,�ɚ�~UF�/��䳏Y#��N�~�k�:����u'���]�.7ڒC�S}~�HQ�W!QQ�{���w�'`�*��s:k0���bC��{}u��W�{�uN���H	P��R.�>LQ
 F�L�'�T�a�_h��|�o�8�(M�FzV�I�܈=���Ϝ��dÍrɣ%���vg�ũ�kJ(�N��M�P�D(�Ex�lؙ�������d+]�t�����X�!(�3/p�������-}���bn���o��-���ѿY��$/�fU��r�@�
S; ��z�./�\�����]ϴD�T`7���\��U�Σ'GP�K�iQ!Z'Csd��� wnf�LWA�T���8#�	�P��"�*�_�B�5��#quu-�zh���(��6g�]@K�m�t�*@�%]"$
���t�#��V���8�i�<���,]�۫�_,�^��U�>k�wQ��ڋ{{*���'��]#P=�ה���W�X�V4ig:f8�ɹ��oM�"\�"�k���>Fh
���1�[v2��we'͖��l0ם�dPEX�Uy76T�'�@�����\�[Q����b���DU�6����,�d4�,�ame�P�ۆo"*�����m�G�:�C2\���.�.x��K�q�jy��n�&.�<��і����Ȥ���Y6�Jh�­�Ukqc(�`C�CCr�.�O�����^�_��3�͉�0���1����O#�"X�����d�ر
j�%�
Anݡ{]����.�F�>a����Ԕ���x�����/!BӲ7�h�@kh�h)�ЁJ:�rR��{���M|.��/�(p�l���zF����X�2���窟.s�K�I��'b#��l&=Z�Xk���L��i�KBCr�Z���}��8S	UB����];���)��
�������)��6�	^��`huXv`s���������D�Fh�*˭�-��ۚ�Վ��w�ٽ\��]͜��Jn�W����*�O{�[,�eA�?b���F��pC1��[�L�(�WB�o���a߾�]C�l����Y}]�^x:j���h���IH(�:>�(S��5�r�����,���\"���/��NP+�N[.��J�e@�bA}:�2gdhP9�TN�(m��֙���1�f�ĲL�W/��{N�61��3C3���ǌ�3�p�0�Q��X�KL�������w��,/�[��H��~�U;�=��s�W��"�a��+6�R�R��,Ҷ˅sy��2��f�\��6.������H܀���Kh2���%Q��e^�\���l4�-��쮂4!�I�>�3}'��G7X�j�=Z�[g�\#g�KB@��{�mά7�K�X}Q��[J�qŸ�͂`��٥W航I��z90&gѦ�7t��;Е��/ђ�3;Yw��1P�!������^뻭p�i��cMvwjHU�g J9oh�ެ�oF��op����֤\��]Bb��cB�d�V����"Z�����e8مZ�]]�-�ghԙO�v%��Fh�m�x
7.�>�ײ���joBsk�m������>�
̚fpΰF+d��(���KKN�0a�Oy��u��_�t��e8��Ah��GTi�SѺ;d���0+��0ky$F0�mX���(S�2��ȥ�S1�m�xql^~��?g,���O#+�����6��#}yJ��/K�6�̻�VV�-�"G]m�Xz�Q���KY{�L8A���)X+-��/;��9���ꔢ�8�6���:$.k�t�W\n��\5��Nb\[�%�u�=6�8����E��J+O�wMR�Tq2��-O�R�ܲ�Ru@�֭�<<�{l���zIK�W�p���{R�l�ȸ#����3ֱ���CkғTtT�X�J��ܻ�5y�,��i�Y��zo�"l�V�8m!N� b)��f%�wfdlUm����^%����hTY���7�������o�R��b��B|�̦��8�Z+�J�RI�]D���Җ�C��U}�ޛ��[Wއ��%A�:��h޾�W��(��Q �G��m��p�h-/
���ij9u��:�N�0l�xt�يj���q��)	�?|п<bVa;5�ӱ�Vv�w�r��kbh�t�h����ePՓ\w�i
���K��;yVX�٣��e*fPFN�Yxڂ^l�Qb��F���+ٙB�U�F�f��Q���X�~	�ncC�����2��f<�]����ܒPv��ƫ�(��D��2���E~��75zF�n�vw��~��%y�SgM��j������hwp@oaDK��x�+&�B��M)�[�R�ɋh�SK��	8Ф7z�B��W]�Y��@�Qj�$��/�u�Z��--|�ZŹ�gu���2�o�k�Y_z;/5�W�Um2�T��S!>7��_��l���OQ�X��uŶ���keP�В�)��gt��&�ӼM�a�r�:���U�>Փ���*��!�M֢Q���=�n�bG� ��o�f�%YO`�:�sW��~k��ĶK����,�~��l��0]OV�1t����:\�qjֿ_4���W��6�$}�hI�3��M��z�(C8���ְ[�}i4�%�D��uI�ec�%�����1�k���CxSTVΧ���v�,V���;�n�U��`��A2U�,�W����=��c��T��;^��/��AɈ�}	>V߹,�����쮲Q茉r���W%s��w��]H�^d#8e?C�ZW�S[���2"fd!��P��=�J=� :�ٮ�a�})�Ή��c:����?�<c�%7$|u���|D��3t���5T2��<S���0%��ltč5C���˨u�KA��'����{&���,�s�TPlŌ8q6��\��-��\�Y4��
�KG��y�]]���
#ڗ��S%
n/V�at5��Ob��5dl�,U���b���^����	pr�Y�N/Ux�,��#���8�#r���H��R�Y�3J��o�Q���W��E�rvWF�:}la�k;����|K���%��5�l�W%z6xsC�L<^���Ŏ:ĳgK��M[�8�:�0O�����x�Q7�`�ڢ�)��+�ȴP�[�[�|��=9YH;»�N�4mv���0���u�3Q�H�bvZ��fF
#Əe��-K����s! �UҐ�K> =�����o�R�3"7�����f������!u�ve՝i	�x��zu)w�cW��wZ� ��Z22�\�x��N��PJ0t�ꐞ��n�m2ɩEݻM�<6�f�,V�O��@�JÔ�ۘ����NQmsq�T٥�������/F (���fg���)?G�e7�Vi�K|9+TO�R�Q�Z�r^�=7gy0���t32�m�C@�A�8Iѳ=�щ}6N�/ީ*j	�vC�]�A8�~���%zRY�p�z�V�GgǗ:P�Z���˄z��W��:�p4��*��I
A�NSx(ȹ�=`�2�I�3h�
�x�M����o��Rm�]{w��u*�i���4E	��QLܭ\N|y%5n�]�*I}��M�) ,��񍫡j���D�]l��
�©fj�#��P���hVD���S>S�g[�3�q�J�@����5���B��@t]`8�'���/9��.
t-G4=u�|CEr��j6w7R�d�tn�[�T���%�^n��i�y�U�(�9�k*>�ݎk�%�fP;	��O[\�u��\�]�[��.�O�M?F��̨��Up=+�ü�atj<��Cٶ4{���^|"�e�J m��AoƏdV0���X�K�9D~�������r�x3K���"n?���G%K����P����G��f��_�͔CR=�;w9th_T�7��
dIPw	i:8�v�?c�0AW[ģǮږ8'��`�,faV&����:%Z�wm����8+�9���SS��핀�ga@�-q<Uˈ�؋�H�Au��t�S���+igf�gJ�,f�M5n���kh��ծ��oWW��0�I����ږ��J�O��F�o.B�Q�G���I�3$\h�(�f�i��G��7�L�d6��jKn"u�ִ�or�w��K:�<n�s'T�ܩݎ�g}0��P��@;����D�����p�[��v<W���lp;J�7��꿦$[L��bbx�u���Mb�A;�X�ddv�*�d�)eE��M�̡�y�[��sf3[��#}ĩ��#2�`٘T�'�ӹF�+v�;�1>M�w�-�|rJ�����WX�Vn����:�t��36mЭ2�C��"v��^,t���WJ����]����j�('G���N=�vȾ�3fx.����$ݍ�]�G�|��NA7����M,:�.�\�9gB��3B�.�e2�!��ܝ*��y+l���I+����X���AHv�d��V�$����p��5��{TU��Wx�����׳��q{k�7W��C����Ԣ'(��<�r���l+l5]��<��q�'!��[XQB���s$ɰ��/xZ�o�<�$G�DT���Sv�sp�̹r�c�cI��r���d\Ke\��`�����-�.c(�6ܲ�i�����c2���(��i�\[eƘ�a]f��w)��d�1Ů8f��Lnf�iEcF�l��cm��`�&V�EQm�����cs-�F�F���aYs��R�˖�(�R�8�P̡��X�+6�V�̦R�Uk.f`��Ur&�V:�E�&8e0Tm���5�5L�aP�n�KZ�3.2�l�m��Bb�b*�Z\V�0ŵ�r�X��)�aS2˔�RQ1��Pۙ�-��ܴ\�8хqpc��#i�Y�E3+n-�F(�J8��5.ٮ��Yb%���R�(�ɉW3*��U?yw|����N9zX��7��&�5h�+H�:��íQA9WѰ��;ͷב7�~���\�i�^�&~�����Ŏ+��R�P*�fk�z����.�Α�SRY��ՇH呹NOzg���9�n!��.��,���J�*�E���H$:e�B�Gv
���ukP$E%��3mU2�C.�V̐��!.�.�t��KZ�{ǷE��X1)c�T��M��+۟���b���6��-��jj.��mN%>��p�x�Y��3�xQ��AtJY�����N�x3fP�8��z"�tEZ�W��2�1!�f+�t�CgX�eW�d�9o)�&:��/�B�:�̶f�Ncn�	�5�NW��v.���Kvh�Y�Nؐ��S���{U����io�6���M�sy������� �:v�[t�	;�@���v	��`Hr����F�ໄ���/�����[u��Q�#c[W����Uz�i
U3S}�wnu�S�����7tv�ڻy͞	ĭ�v"�w:ː�9&��'����J�u��b �l�9%g�yWgx��Q���V�6�eJ�Z�鉗��:�s^�(��ޡ�B�Hk$���7ֳ�L`���dc3^��_;����6Uwut���:���O�$�,0>��}C�U�����%Y=}+�n�;!wal��N2�j.��p�Fؔ��?��Q4���۫��ѱ��z�X����W;�>hL�MF\u�z�P`�K{/[�>㝸[�	D�'�^�~9}�h�j^{��Ff�S�s,�#�(q}�f�q�Z.Nٝ���k�Hv�<���{|l��OZ��Q�Z�����LjŜ��R�t�V�"L�Z.֢�s$U�P��~������%1�������&���>����!*�:���w�����^�g�D�S�ԏs�H�{����ŁXՍ�6���vfDVV���c
�^�2�![#�����ci۸BË��}�q���lE�#w�+�3<0Д���f*]��S��Qq[L�,*��&�>/1W����H3��r��y�4�������s�P=�
���0���ޢ�Дq�8����V#yP�n����m\]��;KHXB�"�>[[mJ���^E����չ��B��|%P��z�s��VƻΧ'n齎;N��#hj�����iQ�`�z���+�� ,V�4��RS�s7$��VAV�)���kN͔쇴7fuRQ�Ž��_�3��
C"�L�A%��E�;��=��Y��pn�{;6Nqz"�Ѫ�`�1�瞎7��j�lW,y��w&�e�ٰ�����������:��TR�Ի�9id��8qWS;�M�g�̡�?�����m���Z1;�&��AXC��4ب^ƻ��	��n���rm�gb<W
y�*�I&.���^N�å�ju��!��{u�)A�pcG9�T�n^׏0\G�s��HR�^�ݢ��9�un�.0W!���F���7�E)Xr��r�F�P����{Ԭh\+P�:js�3���K\Y�KHE�6h_*�N�)��� j��_(Vz}a@�pl����>�r�D;���!Y��u'u�+U�y(a��3���fs4�!�2��ad.�Bm�64�����lꏂ7\U���`��(q�zI'wΎ!/��9�r��m}�<��;�co~aȌ����ʶ������MS\j��{O���^J�~CgU9�鬷��+�gqN����7���9�8,�a���m�p����*nβ�.~�y)��]rB�%T�7�D�[F�R�.qD�&$�0�P�O����kx��[
�H��;�aS�}�6��oX���ם#:�ww�Rt��Z�.ȯO\���	A�]D�,#9V���ŌU��̲��A291�-�����X�J���6�tf
���cj�5r\���O�Ipg��z�M���a)G.�bӠs�aNl/n��k�$�������hNƮT�k�fP��q�X�e����o"�TB�f%@�!�[7X��7n�g)>�]m�sd���-PpƸˮ��5;�ࣹ�����yW�x��Y3����6R{'��xƷu�b�[�S��K|SN;�f�{F�w��)�Z��}z6��k�x2L�^�8����Ts�a��/����KD7��0L#Y.�v�3�ŋ�*߈3��+2ښ�s������=�Xs�0h0�,�RH�S�Mf��-5Z����f!Si�(7��)tF�7�e�+��]s���͔�]������5�j��xnpJ�:#��t�ɖ:y��W�+��VO�Yc�^(ಝ^\i�G�iW$��k�o;w�M�S!^wu�%�_����z�ҝ�/>����^Cews��XU�۽F�������� ��m�9�v��ne��V����\kn��Z�1�hv�S�����Y=�Ѱ�ɩQ3�v�ܐ��ʺP�6�0L��u�DGs��3V����]B���9��qOϘ�/7*V���isK}�̋u�n��e�.ݶ�E��+���l+|h[*'HIsݓۛ�G��_>Ϟ�_e���;�A��w�
���gY�-���=�>Zd�%��s���d��ޭ#�x��z9?L�Í�}�k-�|�A8cc�Wr���x���C`�02[���k\�=U-�잒1�"��wZ\J董�0��Ma���K%�u�3^*gJ;���~�����B[-<�c��eF�ZC�;Z�rA�pJn��-��}�Ɉ���mX�;DP����Z/1T��y2��5�jW�C��q���Y� g���}�*�ܭ+p�� NU�����J�=�W3�ԍ��|�]���8fe��؄"!X�G��h:�'ܫ+L���,��"��-�)gx�Hq�C�2�(3r�,	�
����\!��U��VUZ�o-�͋�Y���e\�}Ŋ�ڦ�W�P�����K\�C���5�E/d��j4lm<%P�u{��t���N���Qd�.�v--��N!#r�7]m�f���,��):��.��}��rk�nNͮ�:���K30�rz�����\���PԺ��ĮP�h�ue�]�1��Q��w/�����n�]���v@�`�M��̡1�%{d$�WT�޷Mإ�e��\��z�Hl�2���g�H!����F5�1��g�uV���c�c#շa` a�(�gfFr�2�T��Q�)B��D֧�����H^��^_Z�Iq��m���h�]Gyl�g�t��;��3��.�b��F���qQ�۬t%��Ҡ��wHOT�EOwT�8��)��R,`M�נ�Cj'z'B��M#!Fur���a�M�{���GC�F��s���P!��bޤ��-�w7�/Mz�*�2��BA�;W	ع˹R�g����%%i>X�"��w�NR.z6����s5&;nJ�j�@����Ne؜V�n=�!n4��hNՖy8=J���5|#�V
5*��M��5E\�X�QdZ�7yلmaU��H!I�NSe�[��r����SRh��O&Zl=Iŏ�+��a���.k�cA�%���g;��Σ}�Ny%�׫�Sr����c�����*ᷲ��a\�[�wK����:�Z��42]���,V1s�U��f�������k�3@,E���d޳G���E�[ى�e���?\�;g�ƔW�e��O:D�����'!n�*Ժ��m)�d������r	�h�Du	m*;S�2�O���ͦ{�%�p���5&�G{e>�.��q��
Vȕ[����e��R��G;s�z3���r�q�8n�8���,���v���µԷ�
i�Cpb�D���5ܒ��$���+�ӳ�!�P���P�����☮�o9#�MbV�V4Kvc��D����w6*�儧��u,�7��jh[��m�!�e��f�#[x�����C�B}g]�P\�kg�U�feMU�`vf��g"㹺c,&�j���hS���g?M��F�K�N"��o�O�#�<4TE�CzR���0ʶ�W������^-S���s �u�j�D9��|�Nv��_�
�dUjHu��1utC����Dy����^��P(N��\$���f��"!<�Y�#����)�2�G@Q9g�-�iWZF��B+��T�P^]GwOf��wI�o),���x�a����i���]
�Z�*.��z��Լ��溹��b��Jc�N�=�5R��h<��\�=�ۗ�-���Cb<�O��t2
�6C����0n�-Xԙ���\�B�Y��M�f]D�Ґ�j�\��u�ɔq���޾H��;��]��2V�r���O��%�2��\��hQ�O+W�,$�e�i�47�u�.6;B$�\g�c8"T��D`�ù�i9q�O��� �]�Qt��d-��D��`�4[]cAA��4����gv�7q��'��NZ�Q@�z�+��EXn.���s5��ց���r���j-�XR
�KG^�+�s�U���rD��R@,��"�Xe�����v`����Ùqg1�&S���=j��n8�M<�Y�`-J���̸�/��ȁ	I�eU	���T�w��!
:�`-f��"3zmNޡD+%�2�W[�6�E�p4���a�X�n����R�Oj�4f(܏1GAN� 8V:�E��	��l��e�Ԃ��D'��%�zK���֙&'s���cYY�NV�2t^�B����e*�ʱ�^K-cr���-IQ�UA/�,�uK�AX{�l�Z��a�GV�q�c������M���Q�PJ��#�Y�aa����]h)+޵�+���hb#yu��Сd���m-ie@��6uw^�F���B:��.����Xh܎����/���#h�J��W�nܫڔ3� '�?�^�Sz�,���6!���/x^m'�����s�uI86܁��n��;��\T��h4WU�&�V�7�uŎȢ���bnNVd�#Ր�.ty>�t�M�Y���9ލ3��7�;���߯~yё*4�Ȣ�`�����3m�a(�c�H�,Y����i,�m(�B�5���m���8�)Jmj��QKh���ܵaFZfQ�U����E��ACl*�bԩUQ�@X")FVs2�&3Z��[5����ԅq�l���\q�,im�3�DLu�km�����Q%AkQMC6��ˎ,��"(,�°������Z�%AT77&�m.�f�Lq��"�(��P���YYYP��.%��m1+1��*+i�U
�Mf�nS&�b6�w2�K���cC���[sЮ�ƭn8�2�K�6Qc�]��UƸ�MaF�y�O]�3Cv�np=aX��P�dv����W��sr���K�%
�C����E�V��}Ad9�<��<Ֆ����m���\�ݺڡg���ȃ��V^+ʼPs^��rζJ�
��\^ɶw�S+�%�!��ۚ6�>~_���}:�D����WƮZ}d�%��3t�rb�'�=��D	�+hO	��SKwF�o4��sq���,'�E��lH� ��a񵷬�Ŗ�%:8�R`�˲^�K��ؾ��J�h���q��֢�u�s]�ii�֟w�X[��*�DK�������^l=�b0B�)��ܛ}~I�ܿln����-1;b��{(��N�ֹ|T^��귖��O*{YԊ<`ǂ�@�̤oqQ�Ckm}Ku:8������
�Jk9ܩ.1����nd��K�9���3{b�y��s�!;AO!���tb������R�\��{�HrĊƬhuv��iV�ɷ��nxm��@����GHT�N�*"ns/��o5,#��$G�	�_,�3�&�%dӤp8OY)0w��T��\ q��&�cLݪA���u���l�o/)��')m^�4p��J�5��Y��0�rA�q]�qU�h^W:E�����#<яԁsͯQ����m�{H���tgNF;�D�Ju��E�D���g*Be�}�eh;�u[��j,�wC�ݛK8�����#,������g>MŸ�"li�+r��nO.�9�Z�����݆��;�u1˳�P����$%D^fG�*Uk('Y ���L�T�	�]���q�؝�5a�\�Gy2�c�IV�cՃG����u��B���73QCH�%�w]�}�2��=@j\پ�K%30*[��+$�M�T�촕��C���-սs�#w7(]��]	��Kjd���:n�kS�d5=���_��q�+�	��3ޝjlC��5W��]�\X�����j���1E@�D`�{�lx뱄�o��R'K���x3b
�7�F�6lL\��m�2�ܦ,���V5����#P�5��Y���^���м"��s�7�-��J�[��I5@�ֲ)NtY��[u�`��#1�u�̯ZoPє�I�..��m)��M{��T`x�9����̓Z�=W���jV�~Q��b�z#7�ӊX�Oo"���駳�B��#Q�aw��������g�9�e��dbt�r�X��4��sw{��..��T�K�/���MΆ�%qQ�>m�M�9Jj���e�R�X�HF�)��E����ec���Y��ڼQ$)"UU����h���2.�ch9�9�D�A�8q?��ǽ����OjN�A���%vv��6;��$�h�]a�z�JC*̶�<<�:g�k}p��= L��q�6�UcL�@���eК\,�OuH%��μ�IiF��)�S�N�ɩ6"{e��.��S*p�nU�)��*N?Wku��s�sk�Oz�}��e�ŲZM*x�{�S��S��!3B�,S��{Z�XB`)x[OF��t���2����On����Mȼs}}6��u����{�o4�q�J\RÛ,��e��X�� t���ɔ��a�楉Om�R��e�ߵ���ؚI�{�z�[��'�k�*�RN�������J��IE���B�G�G��X�g�McW���o���i��ԋm�#Tiۗ�|���&�ڝ���m�.�Dɼ�$�2b=hn��9ASdb�ƬU�fa��.b��]�*3��^��z=[IH7��ߘ��n�9�t@������>-4;�m�fp�,m�p�W��R��w�MK,����Sr�U�x1��ӌ��WS�%�]\����!��(c/i\m�"E�{ݺr�P�,�m�uw��o��lM�	T�_����I����*�%�|\��t$��{g��@��rxH}K�X�J�>����79{/q�h��r�ĎFգ�=����G��U���9�u�Ӡ��:o���z6��!�d��_6�)k�Gg���:%K�1V���>�m�C*�v�܎Y��%y:Z�Ɗr��y���?�߾�__y,�;�b���z�n����s��ZhKN^�~}�uanR���5�h�m����nץ�L���k��k�o��F�y�W3�1���g '~�d1��,�Bdc]��3g�&����%%[��1@Th/�Hr��5}'��NȊ�=�����H��B��I@�2t�?K��8�N{�j�I��}C�)ЭҮo��Ф�N>�٧+�gڳٿw�u���N�l�fm��y'ϛ��a�>��򌋷�-��9J��J����'��������a�����Z^�7�2j/E�A�i�$l�Y�2.��DQƌ��x'����G^ڃ:л�=��,�w���{�6&��*����vK�"�o�Cx��z��Y�T��9Z�7ʶdr�:���%9�3u�nj�hYx(ck}["�V������N�jN/u����]��A�YP|�L�)�Y�ƫ���,WE0�Vr�94;gf��+��/D��xr����\����\kģzg.�����]:'"l�����!���2,Գ���H}�ve@�p���&��#�&&�$��BΤ�}݈���m=���09��.	>�ҕ��鱓1@dM%z��㑲���=a�saz<L�C9;-UVC�WI8ئ��{��V�e1�@"�t��'r20
�Y1��_��Mj�\�l����L2aq;�Cbd�Ƈzs��*����b8¢w��w-��/���)8�݊Ŏ�n5^�b��5��نM����N�)_2'byu2��.a�F5S�GIcۮ��� ofY��s��xȂ�JYNo����t�hs�5{-�}���a/�b��s$�f��V�U�7c����L�Ϗ������9M��1���3*�z��AE��D��i%��	�nh�4:�F#Q�Y8��׸�T\GC��YQ[k�t:�X�S\8+�jU-�Rj�W6�J�:-␴�,ڲ�+�A	�=�u���՝܆�Ӕ�
��y���M��8�x2+'����>��r�pT�|a}�R�Oqũ!�9z����H]�&el��GmJ�%��ɸX�y5kO^r*�i;�B��d�F�#�XiU��ҹ7��[�Qu=Y�ћ*�����-S�#g
��ϔ&^p�����PH��,�yS��+N4�t궧u9s8��m��M�Nu]��.������H�&��&(���u1Ss��4�����a�%G�+�ѭ�{�����߷�8=��zM�yI)��BԈ�ts�sk�	�m����*�o60`K���v�[���u��p6y���MOr�ġA����/mލ�z��="����S`�gq$�_D�btG��@y�&���J�Kr��{�$�NKh]/U�.�z^d�[S��o��Ϧ���Tmu�؞4�ԹG)^#c[W��M�<�����Ԏ�'��w$�A���O�B+�za\w��p���+���7�G��dùt=,Q�f�O"�| ���묪�����yi�fw�����f��]UY
V��M�1ycк�P灉�S3��oD��8}�`�����e��3���u�Ώ�g'1gc������IrĤ�q�j5u�o�R:J��I�W���yDT�&�h��#��5z������P��g��lP���N���|����+#o�R��n0�r�_WKk��`"F�=�����=ۏ���a������T�o�+��6`�5bF�ەm6��+����ZW�c�����W�a,�p��o����v���"B\���Zr�+}�s��;�)�\,\u&!Z�A:����!g[m�u#n�3�Yշ̲y1���x�iH���2Y���EFV#�5)�v:����QY,	j�`�*0��;3Ϙ6˛ä�تl�	����7�Z��8����T����f�
+�e�Õ���d��!�@U�<�8�ؾ˘�v`ۉ�`eq`�����i�χ4�VM���W���$���9����y����NZ�.dܢ�ڠ^���Ӻ	�h�u¹�����K�7a�*-QY����8r�M9��C;����c�e#���A�-��[)���9���(Q�Ǒ��˲�r�$x�E�k�۱o�V�n��V�wt�r95"c]��c�+^��K�����ej����M�F�:Q[�em\�hQ`ty`^�)��]�U�+:!���,���m0��:K/�0����Ϝ���c���	��������=��;�}����K:�����0����(kS�o��̚Vҹ�k���TQ��\6މ��v'	%�`���*�iO�gax�WO/s!,����B��vi�Q�֦<��+�/�c�qRb��͎Ƣ��L�	�����y�D饸��Z�H�Uel�� �7��}�Fy�ѳ�xƄ��J�dV;j�v��-�x�o��1,g���Ϧ4"��#��WEyF�Ȩ*���fZ���|�>��>5wS��I5��Wg1N�k�Yg�����d�� �Ȧ�ց|�֪ѷ�.��+�4OJ�/:'R
Wo�����[�b>m��*`[� ��y�����Z��~uwe�f���'xm ��9 ��S;*�凂��tϺ����(�����sc�:2�a��&� �+ff�9�*[�]#͊WX�w�Ǫm��z���{�@[�{
�̑P]o�4����r�6�3v���.\�N��1r���1J{�g��Eg2qp��0&��ժ�hR��B��b����6a�:��r#�.��֢�{��S4��E��ƴ\4't�\�8��o2l�W�c�pۭ��]-ti��� �ʼF8���r�q\�;V�c:�bv�����VV��fvD�L�S�]L%��|��h�+5���34�"˧p��.{핌�b9��٭t�V��77Vt�[��!��}�4?3v�b"!���2ص��WQ`��B��Q�j,*`��6��T�Vآ%��+�\B�Z(,Qd�`am�LEX�[b��1`�P�Y1��iD�b�b��+�c%Hc�J&���
�1Lj
L@�,�[&�X`���[U��Y1�Y��eUX�+,1&3Y�X�R9A`,��E-��TETLd���$*��Y�jfR�J6�EYXX�h����k-�1.�I�V6�bȫ"�����Pj
6�U��&*(�m�P�T���Lq��WRbֱ���r����^����:]f�z�;��,%�f�+`)U�Z��Y�.�Sʵu��E�*�t6�ï	)�fv�X?+��ү
uA5NL��˄��o$��T��k7����3k�C��WI�I�������&�Z.1�*��Y��H{��fj2�DZ��~L�Q8398�1Sf����82o3O����柣��L�M]�a�4��X+f�Q�Bɖo^s%E���%�i�'��x�TUp��t!y�<��^�P붤�=Ռ�9�#f��+��Hܗ�Z���B��ݯٰ4�V;��x�싉śk�z�)������T+�g�jY�Ϛ��PŜY�J���.�#�JO��o5�V�-;�=��p�Jو�.?`�ےwG�6RiP�Y�Q�cwy��a����s;jN#�E�N�)j���Wt�d���/�%Y�a�ۑΙcʍK�k'25�2"�]���flJJv=���sF�b��*z`� ��{�_q����}���Y�`� ���/@&G!���. �w�Q�{�e8GF3��ֺ��@�(����p����I�30��k��j�6�O���L夦�
g7�"���=�t�join�Z���ut�h>���]ܖZ���0Ƈ;E�e5��U����^4ũ��r��*t#Y�|�y�x��;�ʴ�+�:��n����1Y75�L�Ōp%��q;ٹQ��p����$��gkX��u��)Mp�Ě1\r|mkL�	�u�ghj��e�W�*��Rk�NV!����Zw���c��kl�VM쭶���ҠH���4-�u��s���l�D{�C0ۮ݊R�&��Č�1�Po#/�\��[ɵ����)�-�I-=��7�r�IV�=�ATf���T��=>鵱�Kj�M�n�4��e����d�	P�+N\�e�u���r�l�։������0�֭�7�5/��
E��2�^6\dm7����8�E��Fh��#�[I�p��5\o,���N�SiwkT1;�fODw��,��R�N�we:Ĺ��^������P���^'3gB��=��M��{S��j�i���w]��R�YON�l�yŶ'` �2�������c];���w";G�<Ý�q:!N��k;��L���!`��b~�G�I\�10����oeo����}�A����//c���Գ�L��-����\m����
=�l�6Cw�XBh������V�%�u���8���y[=�j�m�wol근К��o�$��D��)����?/S�2�2j�%Ux�T'u���'=M����o����i
�⦉J�3������"�!�{������შ�ۖ��5��$�],���0�dwC�Օm�2�n�Ӓ�۸R��,u֥WOp9�T�&�m��|�0�Ȭ�{�89L=��;�4�ߍI�����Z�ѹu�f����Ҍ���m�1]N��G���R֧t��//���m�Ÿ�C'����J�E�s��FĎ"���\k���\'�����U�����ۇ�id�gM��s77Kg��Փ��T.,
�/�&S�c �݊:-�On\��T�!g*���O�,aHD[��\xV)V���T�o�w�K�'ո��Z�
�*v=����<�ŉ��S�T·q��+�!$ж	�)�9����;''�3tL�.�۽}j��v���8�N�����p�pHu��f�'ٵ�x�k��qb���VUJtS
�*$h2�А�m�^��B:W&7�ih鰓G�6 �^ڍ�9=���|�Rck��s�.h^��kC>"5Է�N\� �V�Ԙ�~B�oj�1m�Uc�3�b�S����\Zu�LO�W.��vx��k�p���S�c�������u�b�%]^6�����ԁp,��e��یЭe4��,�^0NF��N��9�ֱ6Ę��O�U � �Y���s�U�C�$u��-\���.$�`b{ʍbq���gk��Df�;w|���9�I�� �Bu���S�vdH.&93i�K�+��+��k/���q��5v]��>�zd,Iӗq?��������#��@�{!N � ?㹸_7-r�BkdR��zp��ܚ-�;V�Xȭ�|�J�I!�f[q>C���Ԑ����Gm�팹�3o��غ�e���U�������酹��{�6N�\n֢�8�:�&$�>��jDRq�u/��-F�n��ktѷ֕���&G!�ȹ!΅��9X��ch�p����n��{-�ƕH���x�u�"��5�C�z�h����za�2���=�U7�ZB�7q$B�nW79{kh�!�*���@�
��(���-
��"�oo��d��Oo-�ie����(9D3a��f<�AJ6j�ӆN�˷L�Z69u�p��^;�I8�f|խ��L9WIN��۴o,u�<mdFCe(���[*c�r/�u�]^=m�{׼T�-/EX���]`X��EE���򘡺��&k�Q8�Ne�6��&&�-ҵ$:y���r%�|�Y��|&T�"�9��n�]z��f�L`I�T�0^�{H��9I��Y��ڪ�쎩ڤJL^B�اcw�r�^O���ZZ��b��;\��87]i�s>e�tL.��s��mAܶ&9.S�'�A�%�zHj���1��w�J���b�]b~�]�q
����g̎�V���)F��i1<e�Q�*�����X�����;ڪ;2�i��/�P��K�	���ݥ�e룝Cr���qq J���
Y��a3�$m�(���s/=�C�u7>�m��wCi����Ʃ�����2�i�V��7j�����.�e�A�3L�O�p�`�� q1�6w��ݩ�j�д���wuحu-�s<�;���5�LU�r���!��ݡ��ˎnb��/14�!�)b�ā�48���N4��9��(�q���"���Uj��J�x�i�r��{�b:2[w9�w!$F�#�+�J�b�ɚ�����]��hffUi^�>��8��c:�}�!i�viMGb	9̵��j�b���xm�E;r#��Ԫ��m�2�i��6�7R�NNz۫#+����g2�4�)9�6�Է�WE[H��x��;sz���U�'�g�SW���{\lVW��u�뫺�)Dp��=�hh��}A��"�tF]̾�� ��:�3bxe�W9�Q�E�{6�x켌6C�M��I�],}�@Ȩ���|�oS��M]=|ܠ��=˔,��Sd=۩'1_�|�g:�U�;)2�x�p��f1���S����c�?,�V��*��WR�b-��\�q6�:1�]��� ����'��G�[짷���߾���pڻ�S�[H�d�&��Tv
ޯ:ZkR{����cx��6e�]%Ƅ��k�v�B�۽��>�ze���n9.�����N]�HC��2Y�9�����j��bz�Y�Ke1�D��A|Sۊ���3��Lp��z�T0&���(W��=�(�
\<�J���+`��WX�+Q�v��Ӻ��&�m��,9��.��b�[�V1���P�1�T:EJ�if��\��N���vl��tT�}δ"U)vp���̤l��R�����3p��e���U��&kݨ��5�3��!&@�V�W�8���,�O7�X31T��<wgoczD�He�/
kN�NR��I�;��03�}8��H��i��n��V�X2�Տ�<�Jr��[�D�r�$�X{�9��ǉc�Yap�n���mf�z�D���8ɘnr�$�E�k��i�͟�����t~�{�����'%h~`�H�S�kf�בfƙ�J�ry�yͣek���r`�ٷ� ��Ch	"Y��}Քv&2�fU$��i��,�W%F��k�ܓB�r0�"�w2�Qj������&	 ��6�WLO[H�^�Lv���+]�Բܛ|�9��'�EW꼯_R�i_����4[�i��P�����V�^1Z�}iV1s{���L�"�k���>qT�B��k,f�搳���f̤v�gt�1�Au������0Z��Q-4T	�sM�
efn3qeѩϲw'�_u�r��ڧ��/�Q@�P��R���������YM��)s�
t]� ��fA #�����ʵ��[�q��1PI�ϖ=�++�S�TU��Hv]*�0��w�/fJzd��r�Qps�N��aCX�ܖ&˸�C�:�������|�^�C 6�r�u6Q�E���u}ֈ��.��^ȶ��`��+�҆���mW��+F[Xq�����ƭ�yb�R=���� !up�{���}�
���jP���B���S�X��Nj5��@4�%7gI�\j��PF+z��t�X9��2�y�x�k�{&kˢ�л�(i�oΚX��|�^j;&���=v�e�Gx�o��H�3K]��1�k�S��t|a*st"y%�/MaX�ͭ��J��R�i����mݰ�3:�u�܈�E�np� ��KP@���7��W�z-v�����+<�B�3p�	�iƭ��d<μV���)m(pH�oSGkxU��+Oհp����[��!i������v|�ք���K��/�L�7XM�M�XcU3%��
�@7�f�a��M]	w�zu�N�S,U6:�;\g%ڶ��6q�1q�DLʣ>5�!�Ƞ�R2�����F��jB�ˢ��PK�d����]�����Vw+"�S�k����Z�����}�A�̔�9|jtKH�K\�-�uZ�GK
�UԐӛ"Ml�`ǚs�Wu=;��r�W8j8t����B��.˻wc��l��d�<�^��9�w��uf��syV�t:��!�T�yu��Undf���;e��N�(��h�<�/�t2��9{Nf\�z8s��9g+��ӨN�yi&�^�[��!>���kY���F��a��xf��Am@z/~�}�޼�><<Y+9h��H)r�ڰb(��g,���JъC*��(��LerՋ�(%@QuMfeܦ4ef�J�J���M�ͤ�r�V*�1��,[�iE��K��B�w([aDR"
5�`����X�0*��S��*TU	��B��k�f���q����D��"��mQی1dX�۸@�Z���q��R�Db�h�R�+��E�XV���4J멉��j6�ҥf2��dTA�QR�\d5���ZUAkX�B�����E�(VfWl��T��XUG.&e�3IF6�\�\�+$@���w,���ksJ�+��Hi��Ү�)����^�X��vp�8M�E�Ո����������ϒ�یb[�����P/3Se�rl�A���/]z��:06�����/�̽\Jz:��+�I���e,rp'u�_�9��_���U=;�������&pt�:}���So�ul�k��FD�yU���y�E�����e��KO�������^�u1���'���\gq�(;��N�����g��Y㔪�.�95��J8*~b�J��Ygw��I�Y�}�.t�2�v4Ыݦ�v�-��\�-�D>(���A1d�[�*	��k��(d����&������T�5�p�Ȋ��{o���_��S���ܸV�S�<}F`���38w��%&��t-����=�1�Qr�NPU�eG:|���uݳ^�Z�� ���pn��i�L�|uИ�I���f9||�����sJ7$��#�g��k#4mh銾%�=���U˱�~l�ȸ5:6|��ةPtAR�I4�cL����T���5�N�A5&�W���k�֎�.]q���j����S��]�
��HO������f�i���w]�֠�7U;�ښ=M�����o�i7���S�+[֔�QX�g������!O8bzI=֊y�8تa�V4KG龨`��*ٵ�+�%�<*��V����j��m�! P�KG(*W���.�����	?J{uyY�i*�s�+)'rw�R=Hm��WY�\����e/a���I�K�⣴сr�~3�wޣ���%<��ʄum)���Zr�W_Z�[ɸ.Z�>����1��v�|�Q7��	�NB��.:�vJ{'2 t�%p�W��M_vA3&��<3���Nӝ���W��c��tj�D�8	�T�VU[vE�čhç�Z+Qj
���r?.+[��+)w��{Q;���x�%�W�'� ��S!?�ت:�u7�2/&+��P����f�c���Tƪ�)�,+4|�=�\~(i�,r��mnOU�+�4[qp�����x�%&*����OK�V�~K%��N��gE�� ]�F�$��wZ��1;�!!0]	��N���I��w4�JX�qR�jS���;P���k�2��]�=�4�=!'A8	_(w�̮��C��<XM�畳���M��~��Y��x��nݛBMF䛯.]`ܼ�br�z"�t�n��E�>x����F0�}�k���<�>�� �֣���
�:Z�;�9Q����5�eK;&[���TIQ���&�T�����r�X͍�n�{� ��ڂWM��\�Z(_4.]v��mM^�����@��foUl,�E�wXM����U�f*�V<�C܈k$7��snt6�ξ��'���;�w-����s
ޔKn;����74�����W�;4�yXɡ��bLk�ᕌj]H��pȪ�E���y�f00�e�Z级s^��6���M�A�6`q��d�Q��i#�)�-�	�=R��B�h��u��7�fo�\���)O)����
=u	X�s�OCN(8�X�7����n�b\xs��.`�0oY�Q\��ޡ��ebZ]�ř��]��/��9�U�/b4�I�2�5Jb���k$4BTZ�9vi�;kǋiGh�!J:��R�H�I��ޞo�#~�î�C`�e�n����ץ��#i���q{�T�&Ր�
��s����Y���ԘQ���K��bI���W,كu�u�c����A���������	[�^�ND1R�]��q9yȰ�0�ڔ̇�[Ku݊�R��5�w��[���+`6  V���U�w�j�6�|�tO�QS��m�,|iߞ�	#����k���Ǻ�G�ȗKb-Q����������u�gg��zFEm5Z��� j��K�h�D`�fb�g�ޔ���}�y��')Ҥ�I/��ҫk���_+J��<��Q���b���(��f`�����w%2�*�G�u��ػ����u��KԱ��1�s�)�&u��	ތ'웳)#�z9 ]m�u����V
qㄔP!&�q���ǺF*�\����rfS��Ǖ[]����DVԺV+$[��0�zM�iֺ9�̡�w�6^]r�ԡև�&�st��z���u�ٕ�ZnS{#f���WD��ԡ>�4.wj]���oy���os�������n���t���p����wz��$ׯ�"��(E�����3�+y���E�ryг5=�T������&d�wg�����c�Vz��ҿ>}��{����g9�m���JE�.���NGy��9,�B���;��F;)����j
���%�p�A"�3"�f��ei��e�=a���odB]��q�.�n�vu�E�k��m�<
X���u����vS��g��n:�X2��	Z��	��3�@���Ę3YbqP�ö�b��C���r��/yd֪=bV|]���Բ�
�'^�Es�خ�K�Ԭh��s���'���jc�ym�I�E9�VT׬���� Gj;R��6��c����Sz�{Bq������k�C�1�'/�F�SG9��ecsH��Ne���e�{�0{��w���D�c-�cz�%��D���.�Ř}�(�^r���sMqxkJ�Sg�?=�c�B+1Uց�8,�(bo}H:lE�U��6ޔ��މ���wOM����scE�	m�=�t�2�
���k~[\�7"t�!:��Y�_h6]V_Y|���^���.Ih=}+@ĩ�݈�	R��m{+6�E`�0��[�D�`̣ңSv1I���ְq��Z�Ozyv�<�Y�L����J�]$�O��˚;2�N��S]JE�c�@gi+�l���PɇD��ݒ�Ҡ�����(hl�R�.5l��^�>��絋�;��]V�6���W��k���oc��<{�"�r{�rq�Z�ӯ��R� �	;^�+�t�,]��S���Z�O[�r<m�O���$4�UEe��&:�O8Q2?1�r��CxST7�ƚ)����ob�aw��6��࠱K��p-����n�ҩ❦沤�\�#+nQʌ����,&M�rL_���W�����V:}��]d֔S���'���[��p��xQ<���4Y�잳e{΅,����(nX�H*������.�u>#juu]�����LM⯔��k��G �˯@,��~����y��cN_{�����)�դ�7/��]��|ޭ��/R��&GY����H .���d����p����<��_�"F�uϙ��5c��p��r☰�Yo=[7�ZD�e�c�t���W��u1��^�ܭ�C��S�B��\�'Մ�8md,�gx��$.����N17 7�D��-e���"�����֊.ݶ�[prytI0�ׄ�͊|��ZV��N.��Z�Ïk]͜��P�:CBa3p�ȱ�U��b��} T�SI�㊆'sdĂdqۉxu��ک�Z�li�$�#M�n�KZ�nM��%nl/'�����$��0d1�BvCuB�#��s�e�+6VꚎ-�P���@�� -���e�v4mV�Gz�h�c���t3�=L���a� �*�X��L���J�ոڷ����V��i��,�2�M/��Y3q澩q?)J5�v��������K:$@/�MuآL�����MK��'D)f75�����z:���⧽}�eO*����e����9�
zY����b:1��j�rUh�~R�3��?o"g�kޤ�!��ݚ���+�������/d�]�}gN�ፆ�s.�:����+�ܴzU&�񕪴��{��A��8R�VM���^�g^I���Ņ%8�kVU���"Td��n7L���C]G����nO�CaO�6+gʽ�(ak���#��l��+��w�	�,�I-pf	�%�÷tU�gW26�gսB�ʥ�J�*�9`g�V̬���y�Op{��)Hz(Q�����IB����$��<}�G1UXC�	.��(�F�LZ��=�0�\�(e(��Z����*=С�NA�w�����I�б�t�� O%M&0s�g�V��-J��\���*�-n� a*�?�Yco��K�K��03z�8�sUPQ>���{3ӗG��p8���b
���@D����%�i��a�N4!�P����?=U��T���K-aܡC��UAD���>Uۤ	 �5�ĀT�l+�Z�6��2_qK� �*�mn�/���7��c4ú�`��q��(*��L����*�f�[�,���z�P�&a-$��q�R�Ҙ�)Z���!�Yt����UADѸ�	M���s��WG�Z���H��y@ݭL͇�n�����@�������-9�h*��v�ʄֻ�ji�3�P�B�i�-(��q|y��:�|�1>��ٯv�Կ�Og�bn;�TM��0&^�C z�����A`ʤ�Hzn��AE�9�QU��>bÄ��Y@��fx�� �̋%vȾʊ�(�nn�����R@��2�DE1mE�� 8��`0���akRRa�.��ص[އ�#X��yb`[��*��YUAD�T;��|5 z�*����;T��7=v�����O�^� ���	��NQ���(�?q�:!�_c�\�OOY�+�p��?���*����a�j�����;�TNK�[�LJ���~f{u�@d:.�`5�������[҆a�Y��< �ݎ���p;���f4.�n-��Ȫ
'yWI�~��Ҝ�b&P�Hl�7	�� B�[���y`���K f�"�@D�/�|@��܀p���i���� E��9��%�w\�7X�
.DcZ=��á	�$>��S=���.�p� HKh