BZh91AY&SY8b�?ׄ߀@p���"� ����bF>�     ��R���P�Y�VͶک��(-���C` ��%U*P��m�V���R*�6��$EJ��Ɣ)VVl��� i'e�������Qa�6V�Uc[V�QZ��k2٫c&�ڣZ6Sb�k$4VQleQ����5ZR�f��6� �@�uR��eřkkj��mkR����hƶ�ڈ�[Z�Պ��f�)�a����Z����V%�T[kU��0M5[I[mkSZ͹ۥ5m��F�   mڇ����4��U�\�wX�n�ڸ�QB��u�֭R�Gf��#:7vѣ��i�GN�Z��ۣs�ڊ�vEHյVؠ�@Y�^   '���}��3t�{���e-�޲�R����k{����T�]�e��)�ї�x�yJ��Q�<�{h4�T���T�U�Nw�JJ��g=��]6�����6eUl�l�F� ����   ��E�v	O�z���%	V����{^ڲ����,95�z8V�{��Utem��}��=/����o�3ﾕ]��%-�}��ҥ}��kK���O�k���
S*��րE�l3(�V�V�� �|�֪������=�޲�+��=)O��T��W�>R��Z�N��<�T������U�M+}�X���=i����=����T���m%C^�mꞚ[V��檤"٦���em��l�і�  o���[Pm��W����OK���U��������FN��ޯ'zSӮU(�^;ҡEu�c����jW���.�ж�*���懥)By�^�B�Ռ��*�mm���ml���kZC{�  ����=���ew�s�F���.{�֋V4�y�:�h�k;��uOJ�U��n�w��rw<T֥�t��AT���O=J������W�jBS��b�U5j�l&�II�K>   nr��*���{ޏ�Ҵ�,�붊V�Gu���Uy�'���g�<;�T&�oW���v@�����p݀��� i�{�[� hܩIm��MV��U��Z��  s� ������Ɗ���� �` ����t���� �{�Ǫ#��@�(y��
{הj�(�ح22-I�k7�  �w�@i�ϼn \�� � �y�Mƕ@;��޴z��u��n�4豪 �v������G�<U�Ԭ�5�*J4֩�[�   >� }��AV�. �y�=:��w{ =��@h'��������A���AOz��� �     4   ��R�H�     "�Ѧ)IJ��     6RU5F�2    ���J���h� 2� O ��UU?T�   4 ���SDɈ���z�$��zL���G�~?/��O���~Uu�E���6�U[s�FFf���������{�<�>��_aW�@aT>�TW�?�$W������?�����*� U��5U_�q U�`�	S�Ȫ�����??���,	��!�?�"|2��?�"f�L���
u�zaN�'X厰�Y�)�U�*u�:eN��X��,���*q�:dN��X�	��"u��@�*u�8ȝdN�'XS�)��"u��a�XS�)�
u�:�=eN��Y��:dN�'Y�u�:`N�'Y���)�D�(u�=2�YC�	��(u�:ȝd��)��"xaN�'X�)��+퇬	�P�u�=0X��3u�:�a�|2�e�'X�P�u�:��`N��YS����"u�<aN�XS���A�"z`� ��z�=eN��T�
u�zn�YS����
u�:�?,��� f��XS�)��
u�zȝdO��	2�aN��Y�)�D�"u�:ȝdN�����#�E� ��z¯�G�"���ȁ����A�#�Q@� ��QG���X^��=`Dz����>Y�
=ex����T�(�S�(�XN���a:��u�~�T���� )����X� =az����*��@��3
��TG� �XQ��=dz¢���* u�@:ʣ�&���zʝeN�X���A� ��:�0YS��T�*u�:ʝaN�X��Y�:�=eN�YS���T� ��:�LdLaN���SO��|�|��{���w��^�Qt�rˍ��3�loj�AjXL�PE(��{�[pU]i	V��`V)�I2�JO3o�i��/.^�/4�F�حyR�Ez@��-z���{�|^4�եb�r�]u�V]�z���Ćz�e[�6ά�`�Y�!��kؓ��XG��n��^�"�u�Q����^h���.�tqk�0�;��l9-
a��Y�����kN�qbN���f$Տ�-Q�~8ҳ+wN�wy�B�7.+8��b�j�&�0�SB�a�@&�tJ*�]JP�[��O�n���d�L(V<�[Q�p�h�$Ysl�2�h引�ҫ0Q�4p����Eȣ���n�ج�y)�&�-�ݒeJ���HZ���ѺvM1:����q�u*Y��`wpm�[=�H�c�qZX\��dr�;��8�R���n5���fZ�\z�m1jOLSY(mh�6�Զ�N���G��71%����2�X�1*��tPGzו�Nl�v�X����i�״�2h��C+r��n�Fs3�F���-�ɪ�#qf6/=��9S^6��ȀĦ���4l���fֲȥT�p��X2�����Ű�;[!u�[�8l�T�D\۹)r�i������ͻɚX�hLJJ��n1�	���[�m�U�j�����iZ�a�^��o�U��-�z�lB\�u��Y�a_�85�jCc&��k}2��ѷ�6��H�̵q�n�V��L���ŧ=EB�m��M���!�SD���(=���$���Szi���3B��;-�V�GnTT6`F�9YY0I$��IV�f���l�.�y&0��0]k�(��F:��j��a�l������*�{v_u�/�Ya�oy�xPa"V���� �X��5+݂̬Cf�MܔR�GP��C,�͐�@f�r�Vf=pK�����Mv^=� E�2$������Z���#G�`��XuMї)�֚CstcaN%��X�8��7�	��N^j��#�Ub�36U,�E��r�P�l��:��v�i�&�I��@��{+�l �^^���)5{,֫ͽ.A��G�Ax5��*�f�r҅�	O�>F�����7}�]f#bA�^��̑yֱ��:,F�ss�ee^�ݭ%+�ͳd�V�+P܈�/K�t��{���},�K3��ջ*��
A�V6�Ͳ�Q���I�RYY5Ø�Ȓ��mؽ�,*.
� ���~�+pP���TmH�Zh�:>����$�W�6�r�7�iQ�t주B:��O�m��Jdmna	[�Y�hP�R�%)�ra`��{�Z��䔮�NP̼h�в�kM�iv��+���[��d���m�Yi蔎��5�gt�����iTq��OTc7��\���h�M%ն�7��f���fP�S*�Ki�P��Э�L��:�4՛��o`[4�l*��ÐҧwB¢�<��:����^���BU�R��z����fV�9me���X��3,M��U�#1��v�D���+�¹f7uop�:FSm�\��\� �v��x�ܩ:;xl���f�m�x-*�e:��H��L��Q՘�$�&w����45��o%�256:����[�T�9~x�"auOI���	TUW�I����t�f ��b��9�^F��r�6t�Vǖ��FL��Q�7yr*'k4p�r�㦕��̭�cٲ��Z�lQ�4�T�fٺkd��,���ٙ�F@u
�m��葶�@�v;�k
s[��7���L���s2�wi�+�����1���ɖ�T�r��EM�;Y���P��5��e ��<u�lUx�e�&k����A�M4�DH�����:T.e� p����{|�fCH��v�6*��$�	zS�V	�v�M�q��.�(�N�`s,���TC{{��[6U�tNV�5�F¶��/��LMI��՗V��с��xe�lH�m��W�D��X�`D8��d���9�n��ki��gW- iV�S6,�ik��͍u�gqA��siR���]n��7*���m3�S��[h����Q�暷-]�a>Y��nܩ�xsh��:[�ݡM=�)�DQզTӋZ�5f��Ye�W|�Zd��L�[dэL�G��"�SA�q�IZFm�ċ�ɋ�*�n��b1!�i5����q�_��e�F頌���3|�����̨R�u�ӏUe"Đb-�f����@�vpg��ར��.+ؑ0
5t旲��Il�Xs����{Z\�&駣h^�Kp�A�E�&ʼ�����&���˵�j��L@��d�c�d�s SX�V3#��Y�C��#�.Rv$U�Y[y�6A�kЪ�*����>7L=S8��Ǫ��h��rME�]�e�VT
m�%3��h�
l�i`@��q�%���-������+yk�פ��Sj%k%�-@Q�ɔ�����c&���e����-�l�*�dnKLyE�0�4)�>׊�=#5R�dLDK���n�����W�Icq<�3{�Hf�nh�o�爼��]b@����7=�)�Jf0�^V̑դ4*�;x�!"����������v�����T��܀�Jq�F���ͭ�B���%{qDsP�s*�S2��/*^�˙b\�F���&AYX��"����YN#�@�i��M��tP�&�t!�~��,��Jtb��V6��!)��$Y/%c˧�c۬����eֶ�A�xB�Y�p���T��᎐6�5	զJD�I�Y�e�"����)Tڻ.��(d6�Ɇh��1��RK�n��`"��6^��e����#�N�����K���F\ݨn��F`Эf
�t3ob�5V�nƪ�r=�1o�r�e�F�f��Rd-k��Y�HoW��Tot�l4��Y��~fc���l��{A�a)Kc(a�����CZ��Qb��� JK� ɑ��*ֺbdu�M{.���a�;Xn���.a��5qh�k�t��i�A����vYN��Cr�Ez��-�����7E+ɹKٯi������ո��7j����r0J̈�c2:z�Ŏ�&k ��-]�,��W[Z�(����^a�LvHtO��VtV�ı0e~��Fb��^T
ABԨ[:U-fh�Q�ۙ[�y�u��'l��	m���Y:��ͭ0��1,��[Yu6�b����R���E��2G���1[��չj��7f�P#�9��r�f�٧2�8�[����:��r��(*��q�R[ʙ�@Jø�J���]є�k)�R��$ [�`dV)�/���L�ـ�q��,�ecL=���&ڋ�H�'e���/i�\gn-�A/lx��
E�n�2��V�;��5�DL8����^kN���a%zc��p�����2`�y��B	�^��hnJA(N�����!f�jy��H�ô��ow�g(D!��s�`�+6+�d����Ҧ�4������������l�h��s=�x��KB�Q�D�l*H��J�r�n�
2����3n��}҇1T;bT�5}���������䩪�-��&#@�5��M�rS��"�.f��	u��{oY.��~(�ǀ��Aq\KD���B�jE��N��%Y��nɮ�ÆGJ��#��ii̦6e�EnMW2�7�ۚ�โU��
�kR���XL]3�5�{R�.�Cu��|	�I��y9����^�G)��w�'N�L;��;�5-�xv�� �,K�{�3J����ԁ3���ǐ�{j�B\LQ�,��y����J�fi?��.�`[e²�I`����o��կmi��3%͹��6�T㹪�A�7Or�F�5�r�ʸ�$J�N<��YY��]*^�F�.��A�(G��[�=ʤ�^�ñZi��K����ز���&��RO�=�u��M��ݸ�`ܹoX8�ճ��2s� �UGl�J���T �#Gѐ�v�]��df�E2j�OY�p��n���쳷Y2��s*k)�I�J�`�lP�t�\c0<:&�THї���^ʰ���A:�Wx� ��V!9P����آmE�w6���e�؍7zh�0�6Z71<5��&Q^�vJ�b	#\����4�dЕ�8c�2c��̙R\e@��n� m^��c� �bܛ�*��:�����*,)Xn�J�c!Yx�{#T���l�%��fnG��A��r��[2�b�� %��*�0��*��i�5�i��X9X�ʲ��2��c�:.]��Z���!��9�oK�X���6�;�?9��n٨L�)��eQ��s/kZ8m]�_rT�T\�{6�𭬔r�P�:�hn9XH�@�6���ON�A���]A����T%�֪@��yn23����dh��Y����P�&+.7���y�if��^��GzrAI����Y7e�Ѳk^ب0��T��dflW�T���	L�Ԭ��/�*u�Q7�]�{���b�����{���N%NZ���2Il͑�Bɖq�����N��UZ	�mZ���;�}��­���N�4�3��3,M�� �ӂ����F6�6ʅ��r4k��7S4P�)�.������Q�ƚ�gF�
#U]LҌ�.q�)��%��ˉh�af{${O5Gh�,�f���L��01�*����te�,+v�!m95����p�cLf���k5܁��I�L���/t���ɅT����[�+�SHtP'&&�`�8R�8�������ǈa�[Z�ݲ�
��ͲJ�ÏpF���)C5<���nc�����p��;f�6���fML��uW{X�Sm�N�0A��R$M�3-�-�����?QJ� mk�1ͦ��j�#z*b��r��fe, �I�ͦ�Y�x�j�*�^SaQ���kU��'QG��2�`WJ���YÉ���7�vmG���n�F�(���RsI��5�@�6��6�@�7,���	�Bm�Edڈ�H���m��r�Xv�ݳOho�lJ�q9ycuy^ʅ�{����v[4��vB6�����7	��MƬ?��gR�!�
hu	0e����[L`YA�A��:��6��6
1� Y6�{v]Yg.3�nѱR`Sv^�5�#M��.���㵯Րd�2+͗l�%��Qy��,^������y)�
�5�]2��i�n�i˶/��b8�v������Ħ$S̒7��Xyu�"�l$��)� u&C��� ʫ4onf��%�ԭ�]L۳�"�#�rZ̀�U����5f��PP�X�bxodgb�:{�r^���6�[Q�1[vv�'qm��D7h`i�X�Uj,��Ị!!���F<�%l�ر�8�v+�k��i��u�������M�=�b�K�0�fm!Kc�n����յ��k[v��|	]Ͳ�U�q9d��8�8�XR�HN�h����7wmH�^KN����*�����,1Z+<Cu� �=�����VL���]#��*ٖp��~�u�1e�ז唪E�M#R�`ܻ�$j6Μ�. vM���J�HQ����]⡯�����+n;�a�7sCOv�r�Z�Jj�εL��c�'t����*Q�ٽ.)0����Zŕh��L�YaG�cI��p�Dha꫹Y�D��SoCvH�P�NޭBQXV!�-8�i�Ͳ 8C݉7�ⲷpsQi&T��0�X�2�ƛ�,�W&�Xhe��I���(a;�PÖmx��D�n��c4��9jSyEeI'mM�^m�P^\�2^��6�բ�$f+ٛ�6��-Q��N�QO�`7�[����o.���Fޗ�\cp����T9���QVwB$b�2�5`&�{��p��+F��E�ǎ������7�rcpU�+E��U��E�B#N�	�w��-�׹Z�ֲ�;r�Osm00�[���Hiګ�Q�Q���,V�9)Q)Q;vF�.��$*�f\(:r;���QZ��Ӓ���8E����d�ݬ��F���:��E,�՚�v��[�b
%�q�ֲ0J�5J-�7:a��EЕ3�.�ڷA�Y{q�		��YmhY&�z��U�B����S��������[W��j�cK;Y��ȣu��ʁ�����]Yw%c"�������.X.KU�p��k�,�i�IbӯK{��b{I
�BT������4��G��i#H\�Dv,�����J��T����������{Y7/UA�-�Ս6������	Z}j�
�N#��j�mm����q��c�3dy��6���*�6�y/��r�'����mMHI.v���/^�͹�5Hm�YI�Xj0rnM��!�9P=7I�'uM̌يJ*�f��{Y�U��y�d�v�p����@�Ԥhe�;>{��Y�Bm���4@�O#،:ö��[* N�H��/��0]��a܂��Gf�֥E���g2fN�7ײm��U&B0�l�w2� \����!�=�#�C���w) ��ʕ���x � �	����3UM���"F0���B�'W�!�J,�+����ٴ�י���B�|KZ�VJ"2�2(dG5�ut���U�fL(��C�n��F]����t�![�A��cg`z���&*\��1+!NA�VoSES&�,L�`P�ѻ�@\�Md�fӑ Q����k��3"f�n�I��f�dE��/FV�lB�.]nj���Ag^BfJ02�ř�d˥s{y�8��y	Z�C��s�u��QM뎍�ڷ����S1e���ތ���7����N�cF�i.2��L��ɍ�����22��Df+���n�큰^ �:���U�����1˒�gX�ImZ;�p��OFi9�4]�NC�O_:����ZD��S3�D ����<��Y����)�P�F�b����^fZ����?�t������ ?��`���3����?B���]���̝� 1��.��\�l]�,�0�,��/�%�����co%$2d����Ea����=:tSML�Z��+�G	ɷf�����)=<�ŷ2ٲ.-5���aaJ��}��*�������BrN ��V互�R�G[ӹ3�tՋS�,]>6�����-�`��D��97,�T�;�����H��'Lv9+t���d���'_+�5�ݤt7:�D�Y����8��I�yU�c��3ow���\���K��J�ԵNiH\uf����5�a��tI���O��<j�d\<�C�����X�n�iQ����S���K Y#`��ݚ�J����a� ���u�Tt���;0N��x��)^enZ<�f�Ҙ�$���r;��SCZD�s1�"��9�Z��r��F�뷆���b�/��R���]�N�vs��U�y�S���1���B�i�.��U/v�0��]�O]N�FJ[B��0�!j��2����UM�@�������we��]�y�N�v��8��.X��xU�������#�"�w�`�BC����ej#p�Ά�!j��`�y2�HWV����*�;e;� z�d�a]�T8��R� ��Ë�K��ff+��E��:h��pm�.3"���H.}�똼%��R�3F�>խ�����{��Y�i)p�B%���
e[��Hpc�ݬ}@�������]�tc��>�/�;�?dg�}hG��唎��\X'K
�,��Lm���u�RmrS)rjwR]{�	Bdi���a̲jou�
�n��JCX{�Eo�!f��=u�J+��α���p�h�#�p55�b��e�V� ��̘����˾;�pjf�.�쀆b�;�s�s����N���o�G�2�%&r��<���8-^wP�rM�b���+5]]`L�s��Z�8/^e�bY${3W#7[�4��fÎ���]ڤ���w��W}�� �];�/iwӲ��\��zz��Ө]�
=Μx�9.�n��u{\|�A0Bm���7}��j��r��漼j8���c�<���lҙ��Y��'q�yA�}�9~~彽�!��\���&��5�8Ô�n0��Ӭ��Wv���P.�d*�>�SU]��4�\���]�.�k-��SD,-�>�w{�;u�E,toh�����&����qNw)���#����Z�y��s-6�fi9�����<�$��3o6�oK\Rl��7F���!	EI��^�e����->F���D,���BǓ�<s��\������[�V+S:'m��O�]�e��ݜ4�ڲ�Rȡ�wa����@k�x�I��4���8��傯�H]w!x�K�#��`�R;�hB�<P�C��Vc�lM_oj/�[�J�F�Ei7��9aҮ���,��V�ˑ�d���n�	¢C�3{�H��L���X`�ݏ�W:��[�>����D\3q�v����^ޢ��ڹU�U�#�e�r،�F�B����z���C~;T�_N�t�n
˖7ih��K�qrdv,�����I�;%���\�SW��=م����$���w9�x��Oc�L�B��U�ʜ	��s��P�IJ*d�6��nL<���@2���f�X��Z��wmٰ�3�t��J]Y�j�o��W��댨f8���#�
�m���Ҟ{$0w���Me�U�q�w�`�H�F�R;�����J�n_G�
Vj�rOJnP��c��f_4�p�'=x����ҏy��/Ѝ�^VD(���ӕ�\q�,⡢�g�'0��%g��Lb�Y�̹��aN�8����KR��W;���I|��Խ���ɏ^�(��a���F:ږ2�+݌�3+2z�2�:k�Qh�q�Q���c�;e�x5�F ��[�A���uݟ�K�ɚ�)o6�,���w{ixH\\@�5gk+
���
�Մ��s��,"svd���g3��Q�S�^��^���M�(�4��@�/�p��ae�\�%\��'�ْy�+RX���gk��+S1҂����[�����{3���ȒL[�'�uވ��{짥�C�J��v�	�҂L�%�uڪZ�{�����|T�V���[�[km��!WU�f��ӛ�qB�d��i_�[+������S�������`Oj���uGjqT���u�a$]�]�V��1��k���p�z;��.rpc��ZkufRB����]Ȼ����\�㾻��K�y�Z��]��YjIݹv5j�۽����,���N�P��;�.sJ�ӻ�:����<)���_sH�X>�V���U��PE��L;��M��[�9����Q�����I�6�d{�鈙y���f佢n����� (�W�����k"�۱8�N{��]ۯ�
�ؕA"�̫�Cw�M�D��H6kx�6�u�f%j�g��w �ٔ{�D������Ud��P=c�<�ک��l-�r5W�v��0��:�}���v3��>vU�#��\��k�4���+p�-�#w\7G5T�/���In%F�{�iM�K�5���ky��Q�eoe��sq":r\���#�:��	���9bwd˥�"��U�4�3:�t֡»wo��Wu�v
��fc����r����z�tG7ۃea�td�5�bX�Q��/���]����6)!�9��*!�ٷa�v;�@�rm��z�(��{\�쬠���B�F����7�9�[��I�T��v�Q����e��]\a��=����6�
�ܾ��V��)Ҧ<�big�L�Iغr�MKy�3wOЌY}�V,C{	�&Ѹ*�[�	�������Y��Ѳ�M�$~��m���P��};a�uKP�R��-f���5a�.���Mbнݬi�<���B/�x�M�oz�4���r�s�Է{ns0Aa�nr:B��{n�2�n� תpw-sJt�$���fƝ{N?�PAU�#n>F���rv�{�S�9#�9�ھf�g�Stڰr"���ۉ��9\����I9/��ռ��fg+8tM��*����#v�u~�\��6�s+N��,Ҟ:[}e����jq�3S��)�/���f�Dn��ūm�-��^�eW9֤j�Yx�,v����e��B��7)�FY�7�e)i�@c)�.����N��GZ��X����Z�Ǎur�1fM-�fb�����·��&�o]�q�X���`����]�v;��ٚ�d�����c���v�qa�H}~��xf3���n�sU��B�ۖX�ӥ�k��v���:��kw]\�%�l��R�:�|j��d�M�X��/#P��Cs���
��ݧ��2���:�4sg:�ݐ��K�o�,Ŏ�/�v�W} �ݍ��ʚ(�:����]?��e�Q� s��b�(\-��V����d�R�I�6��4�r��_�n��ᕈz�q��T�NUn�%�*��h�c��`�+1�<��ZtX�+��xZڼ��G�d��1v�\����!;�C��Ɣ��x���&^p;�1��&�`�k�V�5��j]j�n�x�J�R�p��K�8��
�R�,�]-��5]�W�dP�YI�e]\of	�L���o2E�)w�d�	�@��k%N������F������婨j�L��Fk��JĨޔ�mQ��˯\&��w5]u�gZ��7rI��yZ�rޣ��mMÒ�3a2%�2s���[p����X%��m�λ�p�������z����AN��*f��o�l��阙�'t���Hv5�8W���\�_Ν]bY]m�ui�G��Q/����RE�(ɯ5�6�Yf��Ն�A�*��q���M���]����RZ����8(��s�u���R胸pn�Q*F3F��6$kaہ��^�d��{)9�N&^U���z;���t�=��ʺ����;�s�Z�b�Ʃ�	����(�vrwR�b�G��\ظF���5�+�i.�`^�r������&�G.�+��A��<�Բ��Ɲcm7�R�� XX���&Y}J��'�r���5VN�A����m�n�2vr�3zu�"J�u��:%�o��V�by�S�R�����.�d�+ l���k�̥v^��(�+8�/Y��^u�[��u%=;7�� gt{ι*N.���Z���b��t�@p��%ɑ{��%[���ks8�Rp���P��h��VU��*�Tw�n�e�J���!�8��inL�<oib�x3�� ��];`�:��������V�Q��r2���;��;v��1ַ&-�6x�ɛp�DL��[b�ȟZW�"+�[�Ю��eDGKvB���z����r�t��U�c/�b���E�绷m��);�n�Dtҕ�hc�7N��.�s�bi(�7O^!¨'��'i�����N��`��m8��V;���!�S�)�}�G����pK@d0DP�k�O��C��*ouW�އ�6aY��}Z�e:�2�V���iؗ���K�J��|soN��򍱌2v6��[J}��(=��ަ�v+ ǣ�rYk�b�h>K���vU�Zʎ���}Z9jkAsk-�Q<��{�`����[5��~5�.d�V�p����<ͺ5��5���@��T���	�ͣ�mL8�SĨ9���'9z�aն��J�9��R�x$�5.�.Kq
ޒ�v�������-�iƆ��y��6"���vl�w}��ډ�tpʾ��z ���=�2�x>�.X�)m�����/��F�V���wt���N�b�W�mX�v�Ў��u.��8�9��N�9�de�
@AJ�/����ʲ����2��fԻb�K��L����u�Ri3���8b=J���wۦE������
�9�䧦�\�9Wc�'Nj��v���t@q�{%�ځa^���p��mSJ�ȳΩI�ثy&uډ�؍���(g-yڸ� {LȂZwo���t��Қ�A��Ozw~���p���g5�Z�{�x��ϋu��C��8� {pT͍�P>4�VD�1�9!0�}�c4n12�^��A�C+��+�m��J浅-<�,�N����rS�ݸ�̓����({���A*��wr����N��a���E�Nf\��՛��®������V�,���©o][�O�����V.>��cа=��yé���$v�F��탦Q�U#d���IuՑt��d���o� /o&E3Z��u�[0�|0aB�.P>��Vj���+�JCT���c�XsT��wmg��;�ɳZO����Y��,B���f�v��#J�b&>u0Ԯ�b6{]�	Jж0%ͨ��v�zs;�%5]E�f�7-�gp(�:M&i!p�Q�o��K�L-$L���aJ�P��vs���.ͫ����ٝ��1zQ>v�X��k�|n���ag*���ɇ�ȶ����Ѹ��c��y��V�N�l7���m�k�z��<����:��`�U��l�iHs�X��-���N��bѺ[�R�N�u�Y°��NU���u,l�4wi�[Pc�C��5;�R"��t8YǸ*�g��r�6�y���������o>79����-�otl��X��`�"�S\���"�{,U���c��A��ZK3)�L%�Yf��n�<F��]�pu������b�����BN�9�h��fZ;��p��7��Ұ�%l���H�RW'��jh�'-M�ܼW�8l�M��0��rs!+^��|l�V5�aTT��L>l��(�>�a�f����m)֏
�d�E%]�91���2�b��K>Y+�>�z��Ӗ�S�{�.�>]כS�Vӛ����M�M(����'8�&�].X@V][λ9�
	sC�<ugCx_8yo"�:$��L)�h�@�u�YS�@�h{P_����}/c�� ��>f�	^�En�&�bv�9�1
��9CR�w�Tv�{��������Ws]��r' ���5	ۼô��a�@(�F��D�.��۽j�<PZ,��B�7v�4X���M�,U��q���͡����/pLv�����1��u�r���ve���ӹ*��s��6].���Hg2TX�;ǉsBZN��N�U�toV+�6�AJ-ź7m���Qu��\���`�S�|���6�je\��v:`����l{�)����p>�u�s(��-��.nԔ��n�E�Xή�R�n����%N����|B˙Ȝ���Jd��>�8dްk�܋y�ԁ���	{ϊ���HA�(�6.�.�3![+�wm�5.GvZ��WZ�Į�I۵�bܾD��:i1�t�RH��luJܪ�N\���s�o:z��i6������㗴6Gx֪��{��g����4兼�=:�:&��:��Ըv8�F�ABQ�eXbQ�tʎN�ýzX=)N���ƚ�;�k6��F<����@-�� �so��P��;�
x!M�|6=:�b�1(��5��+�F<�e	�>�2�ť�{����sa�P��:Vf�������P�5��G Yxn�\�k&��f��_IWfit���)�Ɋ�k:96m�=$�'$�n�OgZr��4�$�
�IrI$�I$��$�s�I$�I;�������rWgBF�,/�~q�"D�مI�0�&f�5E	��"�+���\zt�B���%4h���
Hf!(�"�UForR�H��@i/K.��]�V��F� ]��f�0R��9��tq�0D��x��"�CH��m�L� �#;tZS$`���L��e0Y֎QL��w���H�NT��I��(�����D��d��XJWiHS��e��KH�KA�G.�d$Ah��M���\�?��sx����=T@E�~��?���*�}}�w��{�QD_�J~������c���O��0��6��ܩ��#�ב�v��(�i�u��fRK+�s쿸Sλ�����Z5Rvm���N'�r��+ �*R����ؑR���k���g`t�Հq��wV���s<�^���v�k��>��d�s�D�L�WJ_��+JS��������؍�㊛4�]����7}�:Q"X���x��0R��2�@�dJ�,`i�+o]Y}Y)Q���+5e�9%����l�s�=�-��DA���xڀ���p♼�g!.о�.JQ�mKL\iQ��ӽN��K�n�ǙQ.p����\�ڄ
n�"�_���ܧX�Ǜf����P	BUO��I�;l�X�F�g:��譏_M���/�[����s�&^C�l�T%KI��Ա�N���Aj��F�th	(V������O�o�bK���GR	Z��Q�� imu�ݥ��}�B���s��A���a���+l�y�n��<9�7����7���`�֪qAo>�}��/�>���v�nV�gCo�Qr�h��QKz`}�Ama;�PJ�<'�<2�j� �N��k�D�n�49���雋��2�3��,���ʎ�qd<�9���j�bB��o3*<y���vp6`�mK̡�hb�W�b�0&�0C���<����/:�مY�B֗�⮇:+�lG�
�o�:�ME�
�+�S4�"�l��S�\.�c�j;gEi�]��tb��僷c�2kcFr��k�1u`�[���J\0\�E9G���yV�3SK{ ��30Lڜ����\Y\��t�+E����z�m�Oz�-�aA�Jxoka4a�5�`&
�`�ty��z�d��\�0S�(pZ�m>�R���:����2i��N�Th
݅��凕5�q�WHᦛD�Ƕ�i�w:�Js 
�y8����u����u ���]S����Z�|�����e>cV��������<1f6�B���Ť�M��yMQA\���/p;Y��q�1�J�]�������W�ط��v��kN�2�i82�ve&����ˣ�)bl�=W�U�[���V��N�r���:���[�2~Tu�5��U�Ƴ1�Zy��G��.�I�e»J������Ҭ޾�k�3e>�Tg@�n�(\�AV��0Q�]c��pZZ�8:�����g872T`'bl����(���!q+B]N�6�VS�:��P5�ϋ���݁i��&eD�H��Ă�%w���8X9�H5��j� #ZӶe�����߇%i^�`��O5S˦��8ql��`Z��X{d�F���2`���*;G������ek�4;�b«��� 
�1C�)Qv`������Da�4��j��5�VL㢨1v򹝕��\hEHB��b��^�4f�(8c�����>iY7����Ү�,>���w�:㔹s' �[�L�Д�ɗ�.i�k�E�J2L#[W�L���9q�-hE
����,�c�ܴ;)��nb�y�*�ǅ�P_h+�e'�Du�]Ϭ�0oNwp�ʸ���4�L�"�k�f9R�b�����Oi:��BuZy]/B��t.���Ogk��:�V �9*�3���r*��l`��%���[��PX1��
*)|��ܻ����8�`�O������Cݴ��tm;���EՉ;�n"])�Jpmj����a�6�i�;~Tڸ(N��o*Ln�1��n���=V]&D"��T��o7B!��u��D[1'�9��^镜Q�s�����\�1ͥ���⫊�3"��o�;Ѣ�Vc]h��H/�Xu������{�p�p[�`͕�^=��E��Ȇ.�OF�`�h�9[�Dѱ�-T8��c�m7� �9Z�t����S��AI^�n��e��1��-/�յe�];\�Y�e�H���E�3�t:���f�TRT�i���yے����q�4P���y�2���Q�s)ք���H��2��;[�A=��Y�s��g��R�^�M����yx]͙�&����f4��ޅ��ܥ����Onu)]u�6�eT��ԗ3Mv]�s#mՂռ���)n2ԝ��2���ŨwVB��KI\��FP��{Ǆ���ӄ�'si1[��<���7WN= Kb4������ Ѷ7���+��jOs�Z(�z%L�wTxyUݳ7���z��}�Ц"���7����x^��F��r�%�+{ǳZoI\�Ry�����椩YW�iI(º޻\mڃꦪ���_v����X�/gN����}6�b��v�z�PTN��U��á��r���9�=*����4������R��q�HsB�}�����t�z�S��e�:RA`z�Ź%����;78�����X0�P]�+.��ѓl����7*x�lOŞ)YV�7���:&�+�uN���ܡ��Hq�N�	/�Vfl�t�ŵ99�ܾ�Z\��۾1ǛAiaǉ�;_I��z� �ލ��X;q�
Yz�̴��_�=�j%�n��U�9\����^͋[iۭ�gT�&m�����~7�L��>���͎m���� ���}����(I�<:N�5�(�s'VC�nE��$��0P�4����m�)�����:=�<��X�{��v\��afpgFv�O��H!ņ��[�w�̭Z����H�_��ri��P��x��F�^'���}�4q�嫘ۊq'����tз�so����f*{��g'Y��FӜ�{&�C��nQt�#�Mr�{P�#WV�ݨ�{C^��9���x���u� �'�[����Ǭ	䒆�!3%�ᙺA�Y��ՑA4Ư�F���9+m5.^����@���n`Mi�u����j�̤1�!���FgF��Lg��4r�lJO�î��4^�{��fwn_FwgS�b���0�� ��b�*	��-�����lq��l г����Y��Cg�c+K��L�|�u����C6���S%�������5��s��b	�yR��f�+ɍ"�� �s�-BE"�x�ǗN��+�%��N��*���"94�5��"4W�c',V��O�&�� �e�g;z���Z�l)�W9s�I�&��@���Jwn�=�	��r�9��X����],^۷��wP.k��n��V�-WMl���'k�u[dE�����b��N\��p�$D骜t��;&<Qy\�����]Aj�/m���-3J��/��ՋZ����(U�o.����D�k7j�y�L^�Rsh��T�b��Ԇ����v(��al��0!����-���ȋJr��֡�����
�٥�\�N ��!{�:ͷW�g�f�S�VxF��Fe\zǫ���Dh즴��!�w�fߊ'^�e�U�Vr�Kt�gs��PJ�)L��.��ޤ�WrB������;1U�E�/�>�g���RuӐ* �ʸ��%��#���'�ƶ��t+�IV��7���s�e�^j�T��[o8���c�\��u�q�{o�[3SiԻK�[�fT�x��[�r�uǔ�f�Y�:k���.I(2@W����W^�� OE8��6WM�&��tW*�;����Y�y�n��P#'��޺�9�)WS��'rSB�Q��@����I�2k+���X<-�ΘI�#$�1]�km�=�-�dX�E����vf��X����wt�_a�~}\9�U�63/4���o{��֦SL��t�h|�l�}a�+C��6��H|��|i�A���u��T;�tX��s����i�lL
������*|H�[EG3��mvp�A�o$�2��$V�Yz�c0EE=J�X�,��	@�Dq������V�jH	�+�Ջ��5�;a�
'F�����F�p��������u��&�nn�ՙR���U�F��/��˥y9��8����U�eh��j��[�{���&mcط\��72��H!�R�<M'N#�}ۥУ�� �rM��n�gc�z�JN�b�Q�f��w��/��K�<,j���tj�f�蕰0hu*�!9�0^�D�;����wÌ�nb�Zs*'�-�l���+]���n���VY`��C���,���31뛶ٻ	�Q<��`G�ycY����$i�A���80�wrJj�̽����h����Nj���8't.�2�?�#w\mW���IPb���X2�$w��[����Y�2N����C[]�H9	Z�xs@�y��X�+&A|$g\��^����$=u6�p�cb��]=|��˦6x�hǪP����ƺ�]����#�����k�w�+ZoѨn�#e�LP��{	D��Ӛ�+�e�^�l�=�R�/����S��d�^�v���p��sT�x;?#�W-0��	/Z�I�쩣�;X�x���'M��-���k#ഛ�&I��x�{eM:u*�gyضMFu{�(��7tCAYӽ1��ރ8��n�;BM����Ҟ�]�SB�D�/dĉ���v�vP�5��a�B�Z�j���}�]]9]S�v\���# �]��e�<:�1x��-�ג�����-
p�������')�OM�n�+{��%�rߍ���V�x��:�Ek���>7m�Քe�ᬳ��^�9�ۙ[�������#mծ为v�	�囤�'t�릱el�7�hP�G�Z�)�x�[� &]H���q<u�� ��o8t����Djf��u�n��,L�3	+&-+��XP�\LK=g`��zT�����H�̺�eݮ'��0J���ܪ�F����%���}ΌJN���F����Q3�/��lj�[I����]b�H�ʳ|����w5�Y,��`[N�?'n�nsb%=��G(h
�
��'w'���u%fU^g^�������$e���V-_%�jV�aHQ�jWm)����S�``�^@ES��o��f��	�%��e���(!Eٱ���:2��y���}�4�����m9�긭!�H=\��ӆ�O.5q^m��1G T���b������oW0����x��������+~��"r����f=��/Ccta�/5Cp]�w��̆�L;�,u�@�#[��J�ڷ�e1�lѭ����i0gr���ř��t�;<�A���Ѭ�4�5�b�;l����;�効�Q�˗}��n���ieDp����k����t�ŋ-T��j�K2,��<��������rk��w[�9�P���E�mn`�l��u*j	�Ƭ��b�{@h�e�����i��{��S�՜Wiv&]U�F�:�\O�=�(>��]t�޺�_w /�7k)x�ȶ;X��ʻ��ݧq������ꇮ�1Bb��RzSgf�A����X�-�ew�!(o�����0�F��&Q�Ǆ�3�lO�ի����39�fT�8�Q{�g6�/��{Xzkvn�%cO,�c*IL界��V'�2�������zgD���j�B�����7/����պ�ѷ��2=׉\K�>��WY�|Z���hJ�>�£�T�3}�vm�|��Y�Nt?mh/���d������;H��s���`�y�Sw2�Yg宄4�$; y�n��T���u�i^�G{2��:�A˙�tv�#��g]+���P�αJ�)3\��2�u�=R�{�kP��j4X�e�����v�%�6h=�Pt��]�2e�Z�t�� ��4ÔzS�:��=�p�H��n��pi8����^�`3R�l�_��[�*kj'�YE�]����ň�U�:��VV*���,%�5ņ���Vwvs�w���p�4����&�w����b������sZҦ>��B��1�#��V�Y"q`TיKG&<���ݓ��ƊW��N�op�evWeE���y������*;��:r���F��jD��n.'AXv;��y,�Oqͥ
-ʳ� 5J����!p��K������*^,�LV��I��{4�˼��ؘ P`�r3�y[k:��G0��wf��Xή��~[L���HFuV�w�k�Wt7:Z["�b�6�VB�L��;�X]J�$�0,���ؤrΣ��j/*�Ӻ�,Q�Ǻ���(h�3����ReVއG�� �+C�\��ث9�s�KX��Sb��N��Tl��Η2���E�xOE�zr�hb�p��ԝ��
��IƖU����p�c�2g@��p�}���d=�#q�me��c�u��毩[���ܱN��ރ��L"�on\����r���bБ��`�V�<3����Df���͙c_+̀Xd��f�.x������K�"���ap�������F�nC�6���+�ai'%��#A�8��M�.��N��=�{,�ޏZ�C���+^7�ּ���X̗�0�-!3$^=�c��ǫ��,� �*g�}/�b�n���3hr=l��(`lH�n�e��W�z�(�4X��rQ�.}�NIF)Wvj����o_��͆��x�a���;m�W��rg��c%���|e`�ߴ`2�M��S{�M�)��;��՛͚y3�`��ʊ� ��kP�{	͕HT��
V�	���Xwي��-Ԧ��x�EW՗P�����*����Xř���4��N�<FYע�M����Έ��VQ=`b%��W���@��A�Y�Uw�b.MԻy�Bc�o�\N��:9,�y\@��	�\Z���C8�w*gJ�������)�8Ŵ��W�dC��r�+��K8��'���Õ�L9��݉�6�@z�\��.?�%[�kE:���)�K����3���F�ł�.�q��Q�銩B�^[iQ���_r��P��}�|���? W��������w���O�����_��������?O��?O���?O�����}?O����?�}�r��3	��$�UB�)&�?SK�����>�f˞�ش�݂�MY�/U�a�J�^^=y���u���M��I+R=�a�R�->�V3Cّt�g_��3j�fLX��A[�Fvoχpw�,�v隘-�	��F\
��`�I�*9�%���$���l��8i������f��)\br�4+��t���8WP��Om��uo\��`�g�l�=��������9j�f�:0�%ul���8�LN��E�#2ľ�e�wh�¤��u�W�N�޷)$�R��i��YN�=QDnr�d�{]\�����q�����
�*�h�ܮ��97yC�8ީ�`��iL���Ų*4o:���g��U�,��ot�1���@幃��E�
,pD��)`�粌�Mkz���3��Z�u-FC9v�AP�|���G�Y�4���t�>��q�E�Ȥ7|]�����2���̰.=�lЗ������_Eٹ�{+mpS'2���1<���-�P��3u��$`�R�k�-û�Ԡ��K��:��xS�:�Ef�!uyT)�fG����9�������)�Ea^WDm4[��W��Y"]-�P�d�8�jNR�"����c�j�r�Z�c]�v��fuu�'�e������/r�I�N���g-dң�"&Tc�+Y �g���|��$����e�:"U8�M�W�`�!�) ������>sQ���y\��=��@i�F ���u�
���y�D�t�U9��|Ίbb(���<፳MAQ�)J�&
i�����j����4ŬG9�[h������v�p4�r�SAl�U��j(��t�Kb�A|�A\�E:�k5T��E2O�Uru���LU%M�*#mTţU���1�j*
(�'�s��UU�S[VI�N��Z&"��Qm������������ ւ(}`�弳EE1%Lm�$��%2�D��DԐV�QEATl⨦�f��J����(������mIZ$UU�\sM4�QRrެ1%,T��8��&���k��UBDE�KPT��P�:MUDֳA�QQl��f
��I����/~}A�s��of����`J��A��fr=�6;��D}��<��:逩�E��'ju5ns����C,���ǚ�#�l������N;����l`�x�g?IpX�Yz]9�5r�^�_T��:��.L�-Ƕ�^FO{h�o����>��B�t�nD�l,�y		r�pk��n�ϟ?�oy徨��d����{����$�t� ��#���	�nf��8�"��>�w�U��$�s�6�N�:�of��s�zH�ƃ�u$+*W`���Jo�{\���&�`ʏ4�����G���V����dٷHX�xx[G�~~�G�G�i�?)��=E��H��=U8������~R+YWL]ymH��Z���ʓ�=�54ͮ�Rzf׹���[�sɷC��Z]h��Z2��jo�V}���W���:�{����Ǵ��S@�Ǻ�c�1{����^�Y����=Q�`��L �y��sB�{����� ��}�~���=~'����r6%�ږ�~#}���g�j���&0pV�J�j���{�6u}��S�A������[j �1e5�t�����#.�ľK�:�8J�oY�cĳ[�P){o��.V\V���8�I��I�U�,��99HѮ�f�w�v��XB��˽��r_g��6�!zmG�U찌X��~��a~�w�o^�Ie��ӻ���U�~���̨�ͦj�Sexr/��u����Tɐ'�%v]�zz���=^PeI%l�+)�yQQW���,z�z�e?d��DV:~�>��]9D'�:|g}^k9t�.GS�մ�.��(�^�c*�C�W��yUN�w~��^������.-�s�H��뤞ƚ��J9��s���H��a��C�{l�t=F���k�& f�9]��d��k�ip8/"��/��w�{j����������~�Ü-΍<Ǵ\U���c��9'��LQ��7�}�h#��;tk��Ǫ#��eﺾ!��g؜���gy�M��}~�?�������#��J8=�^��⟪2fE��B��5�c�s��$��x��O��fZ��y�џ���oW�;�w����3l+|xS��'κH����]y-m��C�)����:��꺆kU[�s�� 6��ĵĄ;�K��W��θ�q����l�x��mL��pE��8f��V�j����~���#SC�ӵo��!=�j�I"�N���xѱ쾞�/�Eqב�GM����o��l՛0ӓ�3�_nn���˄���@`z<�l�;�1��ӵC��H7�N�94��=�~^�ڥz[���Т�z�����U��Omc��v\�c��{��t������ID��}	�5�H��?�P����t{�-omOC�ۼ#�s�:��r�Ǽs#�-GW�
�����w�;�'����o�J���!t;�h�ZsD/͘�=��(������b�Jk~�tb�j����kJ�cמ6�s�5q�O�>���Tk~4�<���d�RT_9/>��cD»]�mv��OO1���o�z���4���<+c���+6��8�y��Mz�b�ǳ��1�����袻g�Ʒ���5^����'��T�{P�m���}h_a�������M�j�MQ��a�C+�ݞ0���#�p��z�2Z�,���NVI%f4^��'Y�]WQ*^�b�U�t�����fv[�<�+Y¢޵�D�V��ѭ�lk��L�q�Khh��_a#��]�m�#%$���/,葴�=�ˣRz`��9I�������(pV�~>���;����$t�q�OcOm܁sO�(0 �궈�Wu��9]Y=��)��6A2�r������C�L�ڹ٨_�l�=v�DX�<�6iɹ�~��z�Kt3��.·[�!��^n��OQ�$�>��s�\��A�Z����s��W�ײ��n�������$߃q�6	9�m�4���cү~�'�������ޫ�4%y�Jo�����Ϸ;��ڄ�x/:|��N��Y��������͏o��0ܹ�D��7]�������;����2͝<}˚.�����������o��W��U]y�9����l�j^j\�2�wy��\d��{��|VT&�3u���Ryt�O��\{:�|���9��">�7���E���T��#h6���������V>�Ry=�V}��w`�8ĩ�>��������dǱ�??����º���6�^�h�fX�OS��廁���g���]��S[H�ov�.Ne�)S�P��|=��oE]����(�y'$m#��u�Q��� j�$�,���<d��v��y���s`���L,\�7�� .T��R�(�w'�ǉ��-_Y�n�-��	I
��U>���8*��t(,�ӵSh�\¹�r��6L��T�������BsV<}=���~��V�~ϖX�T�]9���[+ޟ7G��u��<u��9�;�8�>rw�~�G��������}���ĕ����yO$���W����*l���?J�(�������Ƙőm����pƉ��m�"g��l��z��&�����۪Y���9{�O�X�VX'T'��Md��8Eý�oNC��;���?���-�K�)�{>�s	mJ]S���Cd��s����gͤ�����
!\����c�t��2�^��7�O�V���vp06ۄ
ށ���6�#aǏ�Fi������R�V����8�!������@�q��'_���l��ʵ;M�|a1s�)�4��w��q���d�3����0�p��a�巘�����������ې:����d�ӻ���ZvS)���W+����][���Sn�V���H9.�:t�)$�V�w�f�WK@s�5���-afq��{��;dX�&���o�$��I�9�*"�z�g�<6�I�ř�/�����f�7�+Z���Kݝ�8����C^~��Z˦��;�;]س=^�S�=��=�d54���DԞ?M5��i�o}�&�/��{��^�y��	�]׫Ԏ}u�u>�y=�ƨ{�~�~D{¤��/qwl;���,|���va-���B�����7�دS���b��u.g�Ozz��#����82���Go�9��Rm\�.��)԰���~��+�*�囔�)3w�1�<{��eX�����A�1rm����/��zz4\�'_G��\���%�@s.2�|�ӣ��8@���Q��X��2��������4��mȸl��nvj��ށydD��H�DH��їg���0<�O�/>�J��K$�;��X{�ꉍ����$e���'���g��K�C��h�w�]�C<t�o+��z�li���>�d�=��+��|����oNt���rC%�{��k�P�V �lՉ��\�]���k���Ya3�pRO��5޶���b��í��y�P��T]L���!F�Y|x��c�>�x;+���]{wZ�@[��;�р�}�qLX�hr78m�5�BH{SoU6��AT9&�w8��w��7n��4歧�9"۸P�.4� �����]��8vz�ks��1�^��h%�q{]�i;k�Ý�T~�nA�g�ި�ܮ�����F��`�9�q�2j��[!��s:�`�������<i���a�����kvx��x�l������}���M��K�&���k�u��_��hU�p:H��3�mH|��y�1`��t4�dCO��rvz�_eџy�U���Ȯ-o����=�f�^WEo�~�jI�?j�Y��߄׻t+3���� ��O�zz�ٙ2��>vF,��'��B̏UTsvn}��-��_\�~ʔ�|)����Mz{'�{ގ=Mz���4�'�x��Sq���e=�x�T�W�ieg�w�S>�����o���{�ޞ���)���t��VX��<�,�	�W�t�Jn�Ǳ�}��6(��=�|I[�l�D�F/��DL}��ϩę���G���<���y��P�H�8NE�8b��'���8:�r$��u�����󩬩wۼ�U:����D�{�!IJ�(̙�;$�2����=��Oƫtk������9�q�������j�Ȝ��z�X�tJ>��x����M�<ef�rV�<}�����o�=7Z��wa�\�Ez�ڶ�WQ�.���<Lv��8��vܳ�����&�$�T�u�E|��ߝ=��W*�`�����%4��u�ގ{6D;�� �/�<����w74�4�QB:���u�}=��+۝0xN�Aov��;����h&d�^Ĺ���y���t������&"�3W�T߱��]y�ӻ�H�<N�$�>ֻk��l�X������U����~c�5���Q���7d�~�q�M�`�a�"g��3�Op���{s�=�O�]<�#���7x{����{F�6�8�o�X-Bݹ^�^��(���[��]W����7�%���"{�ܬ�`s"�[�PP�,ԝ~Ǿ��Hh�֭_C�k��.�j󺍹���D���Hs�+pzi�J��G�R;w�*Wg�kZ��p���
�t:rooz��SEn�2�g/i��9:�%="�v�Tc2���n�m�=O ���0fiԂ �  Q�Z�p���5�˓��{7�}4��o�^K���,��<��;ё�?hW�{ϑ��<r�v������9쪾="M���kc��R�tWޤ���^^�8o�J�kӤF� C�&}� n4���d���푗Lն��<WL����>�{�ڏ(W���$�}=��X}%b�1�n���z��x��u�6�VU�Ai�|�����~N�t�d�g��"�s�Ð�RǅK<�'���	�i>�|9X�|�����e�^�
�yR����oL^'�Y7+3l_��t$i�%�
~��y�`����j�vN�4[t�c1���%�b�wl�W�"Eo	�W"}g�
�26)�Ş�Sy�u7±���C=�g��w�����EQk��:�?c��|��s���T�/�4L<�w�,
����#���2-�#z=�2 w�l�1��绉U������G��
�)�iA>�߼�c!�x��4�|�⒆�'�np[m��;`�C�[��)�Z3#�3�8@w(�t&�����-��%���*[8�.�N��gv�r��J��eb <��'f�����t�'�	���sw��y���M<	�S�2��0H��z{[�Π����{3C5�<�%�*o���r#*�w�YLR������7���M��u{���̾{�#ꁹ�{�{�v�`�z~�A�}�xk�U�����'�L];�wE�ko%��h��6�$�;u�j銺��U����{@���Α�#q6c���L���=tw�����^ˡ�F۩^�*�\�{|n��Zpz���M3��U'�mW���Ž�p����i['���Ac�'V�i�#��vl���[=E����=�.O���:��5�$}�fq}���7��y)˥��E}K��ޑ�,8z�+Iڙ���<j'����mS��>������J��p�|¿:��Po/s�щ��,���*�/'�nH��+�h7@�gC�_h|ޟo����x��������������}>�w��#���^t3Ը����Y_S�ȴ��,ު̖�{�1�I4+��Vk�a)�����4�	�^�7�+l�d�����4BP����M�5�/�3{P�W
h �\�����o]��U�r�]b=:Jɯ%��f.sn,(A�"Kd�� ��{�z�vޣ�p�,M�K�o	`Ź���U���\Ʃ9�`K�k9\$�=&#Ͼ��G�u���&6Vj6��O]���������(m�҆	�V�ͳ|:IJ�E�,29R��^uX�$n<�C&M��m�����N�1�pQ��2J������P���t�6jݒZ���d:�T�҅��n�ie"k�.�%R�nÛ�<X�tj�X���v�tFmpd))D�m��ve��=W�t�-�luw-D�y��g�ڻ�����t�s�s��wB���^�qŕ%"���|{��R�^�2�s�3N�;�2��}�i�]ǌ�]w���
����1q;�r�:rI@Y;��agu���q�[o�FnQ��v)ʒ�b�����f�vJ��N��(�*�Z"76�\�lgI\l�l���L�ڱ2��瘨�wn�ٔq��w�V0�ܦc����ߑ�K1�X9���g�}�Y��oX�+��Y���s�r]�9�J�js'R9�����bJ������{����Ν�Tk��`��I������(l �u$��sd92k�G��}E<d���,P�)�W�
�A�r���՗�s���y:��V�p�mWQ�\�'*;�	 ��*�U�V-�
N�F��+��}��ŽxT8��羬ٯ�"g69�h1I9d�n�ܔ�p�[Ӳ �]"t�պ5�����tz#ku�u�控C8��G���zͩo�B.��\G�,�{������.�7��8�M$.��q��m^(9�i��6�Q��.;�t+zl�b��-p5f��(gS%lZn��]�t�!�qe�={Q��Xʋl&���ڔ��i�I
��E��T����X.��e��X:��s��fWZ�U�+5��"�z,�r�OM��U���-x�MS�|�a<���$���V�p�w�ʈք�4�]Y�U�ENcl!d �aɵ{kiE�++3yIo%vG�y����Eh�_=���s(W)Y��L訋��P�0�3N�)��[Ҁ�s��L$H����-�е]c��\�'6f����+���7]��u6�}q���	�2�f�/��eNlT��A|����F��֢�l�|��_uBÂm�y���a-��	|��T���ը�:�jowo6����e�#��6�:�$�D���ջj�>��zS�u�1N��,1����Cr���0�Y�o��\��f�yk�;NS�
�������cT�0b�K{9�<7;iX�iX�b�#]�N��0����	J����WK�Akwz�r\�_9:I$�������rD�ERQM4Pz�D�LD��b"{.*(�� �
�0QE3P�4�AUO̚
������<�A%!�tMT�U�j"NmPa�������)*j�����$��Ί��������	 %�("
f(�ǫMAAD��M6������O!�!�mDP�4�4�T3͙��	�5H�%QAM?����B�gHSL�ڝ�T$M4V�9&��9�m�k�1%'1�i�-��;o[�3O�֣����h��ִUA����s�z��BDm%tQM RQeyb�F�9Q��U�g�2�#��K��/M���c���ېČ�s:vǜ�c��kN��p���Ƶ��\�X��*4�v4�71���4h��干V��<<+D��9.���;s��&1�ɵ�ZLD&3���˗����]=��,��MR�//yg�롚L�Z.X$�5���ܽ�mU��-n�KQ�8�;MF�s�oe�o�w�<���I�3�6�Ϳ秣��׃�mci=�� <M;I}��6"���2%��q��Bz�X��ƫ�s�yϊ�,�C#��y�uE����P�њ�3VgI`k��C��}��N��{�<�b�Ļ��Yzx.���2�r�#)=��u�������3m�2�*���Tp��q��i~Uw��7�\/������H+�"��6�b.=:*]|Cv2��#x�M���e�U6h�O1��/;����5q!���']I20�ј�-��з�t>C0&Ec~�O���!�<��q/�"�z�K��b^]g���q��A��@�/�Ϧ���L��e���H�-g�|�	%@�͍�p��E���D����2����};�ꆛ[��-u��(��7I���9��ȸu^�3�F��lTs�bm�fV�ne�<~���OT!�>Ȉ��]�t�I�9�o&+�R��XsQ1�����܎��SeWpٹ��+�!0�����������S��|���-��1`�Z~Y��	p1U�筋3a��a��l���\1�٢3�[�",�g�ޝ4%H�$FD����h����ݎ��8 ����tV�v|��߮��
��8����LFl$��훢�i��+�.إ�F[�
Κ,ee��͕��F߅_i�q�}�6	�tw�����}��γ�*Wr��
���S���ܬ �GkE�5�6�3l��\e]�Q\"ٷj�P�|>�MbY݉6�N[%��ʹ|��Ϻ%#Dy���uH�[�;B�;R(� �6���N�Fw�ߐ�H�m�
�^�U�����ڽ�\1�W�>yF��'������y<$��p���4a�X�ǵ�{~],���^��˻cӛ����~�D
'�b���H���6��~e)�̛�b�̠��E/U��Օ������Đ��7(� q�k�r���մ�\QU��S��T�ZrSEb�F?(���62DwW�s���&h�P&Y�O�;/J�7S�)K���E����jmFW��
j@�/���`{����0�f��u�L�����ۺڮ���d�?)7[�����̓ݍ��7ʹK@?�`���`L��<�Ƚ�\���b��&�Ȕ�Nfs�n���[y��p�A�I\�CP_ziT3b��1�WˌJ�y�����7�zo�s[��}su�Ә�%�Ȳ�=m^*O�~�'���,h�k=��C)�^�?��>1g��.=<=3n㋝����c���=��N{��-�ǿ�^#B��U&�^�������}��K��{���q"f˶���]6�N�Y�`Lr
sΊ�q|�*v�&ܮ��*E�+�R���ֽ5/E�sX�H<o�:�u�.xQ�*�!�-�j]����>�&9Ӭ�ok��[7�5�b�	��ײ�N��f����|z`n�+�=�O�_e�9��e�T����ID|=��yE�v�몜k04����oF	�o#��}(轎:ql2ڰ�%���V��qm�r���|�q��t��r��ͧG���6~2�s�O��0G�a�����
���;�˖xjt����q���
�`�[����Tš��ݲ
�8^��ZdM������DcÖ��x_���8E�_�7�~d/��n'������(��Z�D���r�u�5��ҵO�VO�^�\�@KZ}9ע`����Dek^�װGӬ%����(��7<z�eA@DA G��_)/�O�L��U�ə3��L��n�1I�آ��]6�N8��,(� sU:�|���C������<���Q�Z����!���G�0iu;#Nh��_�2��8�Gc��^���0��'	�-��4a�û��4�)�J�@!{��;`����'e�m{��jR�o��kɆi��<�,�t�5�x�W,㯓�U�8^����W|:D�:��-��&D~�}cz#�=�� �������{��de�f"ƹ'1V��=�Q�B�~pG9��O�T	��0��yO�*6��{�����[>4���x7�[TY헑��٬�ؼ�
�|���P��+���� ���ˏ�{);Cm�2s�!�%�O=���l��$H�ނ��e��R�%��Ù��Fv��7w[ZH�H{5��.9ƻ��ѓ%e���zֶ��|���������ｘs�*U^��f�!慂h�j<��I���'I�f�J<�_��K��3r�s�=k)��=�[�~s��j-�6F�>^&Mj᫇;��{_W���-3Cf.P�v�sb|l��T�C���ӗV��,X�"�k��TcR��j������eУ~J�8z��� h��9��ލ9���q:��0������0ה��r2>s�>n��Rtז�p��t]hФ�Wp,��|��طE����CPΛ���Ҳ�;3�'�ʌ}��`�A��O5�%1oQ9�z$4��jqI�U5��K����)P�ȫ|����p*��D�,�M��	���ߌ��ʽ�Z!�^c=.֋���b;�e!�'>; Qttȥ�z���k�b�:	��B`��ǧ�M-�i�[����5��,��O�����y�N�XF�X�ʟ��WGR�@$((��>�ܼ�MSH���5�CS52(Bn�09�Ga�G�q=�U�{��O�~*��P�m"�+��mv޼���M�as��C-�"����+���
��&�b9^}κU?�uuXw�������\m�Y�o3@c��ɭ@Y3%�V�]ǔ�j�O�f�-�T�u.�]�@�p�X^g��n���7]#���2C�(�P�!���u�s����K���̭I�g^������ڕ�N2�u7��1o
�l��wvoY�bY*���k��Ep����a�G���^����-;��F���c��s��_�z�;4ںd�2�J��zV���j�y�)�n��tT���YI��۹'+b�Z�>�:5,F��D�3B9�g�6Y���Y��"'b/
�}�Z�>�|��|��;�t�G}$���'��p	\'�A�O�K�>�?/����s��_�NB���MG2�S���!�Z�_��(�R��a�������ƶ�#ӱ)C���G;C�D�1ؼ�י��8��h5������N�7��`&���oV���#	$8ὲ�r�k�2"�i�SgJ�����;�B���=��t��K`���!���{8;�kNn i�o��<WAP]�?�d�~ۄ��y���ox����i���b9��	�FFS�j}<��3�״]�9��gP}��r]S)��U����fb��N�}�ѠS�@����@�T���"�Ӣ���� 7*(z5֫ſp���Def�嫫������։}?]��ʼ-U��g�hY��p��(Da�Ź|�L�'���Rt�?��@�6U&�B	�bY(Ĳ!R��qk�{U��*��G�t^^�)<����@^I7�`;�p�E�ͺ��m���NI>Y����݋���=�*?���o5,���kf��&�X�Z�_K��7�}�i�yh+Bm;rm�9��6wlN���\ep���Y,8��&�o+zu�X|N�Q�&ԙ�W[�*y���}���{�F���6��h�vk�a0Rq�p��ϡ��i<'�0� ��ʊT�����b��{4��X:q����c<ev��۟$*�O���*��)����.���4�㨮r���)P[D� �޳�l�7�S��ٕ�H�Bu ~q�k�[�dha{��gѻ��T; �5�\�����.�;=!3���ظ�`3_(��Rv�#��E��q�ap��dIz��Q�4v���M�n�i��R�Iyٔ��/2l��}k��蔌d|Q�������Bz�s�����H������;{�����TfV5߻�ԯ�j�*ޯ�r=�Y��6ZD�k ��~���̶/頓�ng�U}�{����u&�W��B����#x�.�x���uEi��~���-O�d���i�����f˅͜���~}�2�$��s4���I��_�͎XШ���30�Q���T*
�b,��S7���0�c6��8s��k����@�f,Pp���@ZiY�t�vM"��^�y��["]��8x}��!�,���7Zݎ��Ϣ��]�����'�Ҿ8��8�2P��)��@oL�J��X���٬��Y�Y����Ӧ엽/rڍ�࠻��w��C�u��:0z?^��`V�R�fI�b�ܮ�eC��-�y�X�T������9A��I����
,9n��m�B�)�Ka C�}� ����^�+Q�Q<��d����==�֛��>2�?����yC����?y9O�������5�U�3�2�5��?^���a
���	+��@7y%6ϛݠdgO<���`d���X3٩��U�=���rvB
��nv*ڼ�O�xa�@�4��g�c��*.и�f$��0�n;*�~���E�DN9�V�l�Q��MC&g��\��f���xR�T�SP�q��y4�����rF]N����^xB�q� 㤛�L6���gЏ	����Ka�O~s��	���J&�e_	5Pj��C6v�\�����!��э�D|fa	���r��"�e�r�>��,bv2������<T�q�-�:�Ě������w G�B1���n��G<��ɽT���V�S\vR�z�ᛚ���f�z����!������حU䴭RVa�)��a��Z������uu�A��.�靑%b�¨䀹�T>U����*��"c>�L|� �8}�x����WM.Y�����)�I�s�s�Mгnd㋲Ut�*�t�N���_x�{c̹[�q$%��0%�=���M=9kW跕Mc�@s�U�/��FjѲ�[[�����^L�W;	�{�w{_f��ߎ��7`�r奛���}�_+�(�=�%���AȦ�m��z�E-P34RqE���/�Q�ݷ�)mL�%,���-^e^���������ޮ�ټ�N9�Z僦��4�zvF��Ρl�!��^+n8����o1�ouuxn=��u���X�@Z��="<Jc#L�z1�bv]�{d���aJ�L��p7x�y�F��(��a�76ɺ͙��^Ovr���[#�JQà,	�^Q}go�k�-���)��wז�38�b���#+2�:rw5k�'���=�2���{P��|1.���2���)��V�oCf��ś͋V�k�3ǲp�C�!0��}(ϻ�]lM�=Y ���}��Ͳ�Zr<���gKwf��G�%k��^=�7cZE�$Z��^�U�C��6�m��*Q0��S^s_)���_v֋���!7�:��K�Q�]0���y�x���n�D����j�^�9"y~)}_.۟��ֶ
��s�,��li�0�D }~s�7���:h�$s�,�j�֪���w�7w��&8��)��ث�V�� ,�:,Ϛ��A��>!��O0�S�ĭ������t��npzpr�X����nEh���W�g��-|�HB�4�_B�w�Wtu,�������~����lL;X���x4޻-*]�o�ω(�d>����#�պ80-KN��t�ѝ5�zfI�qWR<�C/��xA@.Z85���-a5��鋢�Μ�&��j��&����3��N�t��T�����xx}���u$ّ�A�G�����%�u�n�d��|��1�þT�~lm� 3cz	��K�i��}4��K	�R�2��"z�����.�XF�X� S%�a��rԐ8��w�:h+�^�17/���@v_��f֑#X�������N�x��TXc�\�]*�^�L��(%x��arw���1�*dG�	�3#P��.���Մ�x]�Uz���sO�~P7���ڏ5��vz�8�E��+\���Y�W�^;C�/i���'&�;U��M����t�j�������eG�&��umv��\���{��Mܓ��!ot���
��W�fc�G�`1�PnhO�wg5&n���\�F�6�6��t�qwDi�#~��S��Fxtx��ǃǴB.m�iض}|���\�Vj�Nz'C2A9"�{��C��g����zA�ū�C���.�wN*�ڝMj�(��ީ���>[�OxM*�x׽~]��ͬa ��"��\7�;P�c�6������:/n%,�Խ�p��q%hZ`����+-�Q+�ha�0�4��X*� ��>���-6���ب����5����$+C*���O������<:���1
�g��R�!�~\ƾȲ-��坋)vã�`Gw2H{���Q���B�c�`�`���M�ًa&�ù$d�7�N�X�r�m);�^��g���Ǻ��g� x{�\�����:�ؐ_�[/ʿj���ʧd�D��2 �s`MO�����5�S6�������̥�鞺��ZPf�sq7!�"Ӂ��}�(��})�5����U�\eܘ�i����MvM؍w�>^H�Mv4�2kJ%?J3�+ǣ1���o����(�ᅷ��ǵ¸S`�"�DO^��7��+C�d�B�z���N(ϕ��E�t雿Dm��@Y�C��H=P-�#'C��}��@��ĴK�&=� ��<��S�����]"��7e�5v嫷{>s�2�a�)aǖI���Gt����ߥ���$wQ��� �����2���mc]�;dnR{9�����&Y�	�߫s�oC�	��86�G4��aR�q�t�������Q����b�U��K���sz��#��+#�a�\5	��0�7/�Y�^U���Xm� ��nppUd�rS���!��Ĥc�Q0d��w�O�K�{�q�ޓ����~��~S���ƻ�'浦M�_�ϠuT���H���A\A _�������=�^^�w����{��>�_����������]��:����]�p��SsC$S�O�)��{t���YV��E��J+�+�����̦�\{����Hf`�M�D�Q݅��nJc׆�]L���J"c�=#/MdΤ�[�r�Z/�;ڴ��/*���/+���)��kPp�-ڙR���8���'I�gg]��E�\:�0�ӼKqPHJ�u�۰�U˖�i}(��@؄�:U�]��)P�ٽGs^%�h)�4�h�v9Ǆ�c%f�J�nl�N�V9��vgC'�^��!�JK��s��r��t,��s��b��\l��Yr^�C�cT<j�Łe�-l�z� �[0��kz��9��N����jj�<��+.�T��F
f�;�;��}x��l�&C�LV�N�^()�M�g�׫VE�FF^���l�Ggw-q�����T<5��g�S���
Z�}w}d#����4ȵ���u�(ڙYk^�RgS5w��ck��D�L����p�e��S�v�Xf�[b����GWT�A���a���9O��b*�vs[�:�<�U��`�\+����N+Ŏ���3O�ʒ��u�&��f���a���p`��,��c�剾�Q|��=�;Zm(ki\�iw4�e����R�9Ձ�ȳxP�5�F��+X[$��$��Xd��9SQ��QU��L�:�^jt,fδ]kWh��J�|7B�%0�n'n�Uû�6v�җ���T�
��FWT�EW:�)�MY��\LQ	���)�����
θl�.���r����cu�Ӷʡ���o:��o1Φ;�����B��wI뵧v�MWe5�e���/�D�PI��w��Sg��XozVm"=�ҵ���1u����5[wx��&!��l=��\�TW7j{����
����dQz_=q�uk�Z,6��*S6��`���osQq��E�weg�غ�u��K�7����ƫA�����@��10e�}#c��uG{n8�Wv^ &��ዡ��J��a����gN$�%�D��2�k.�N�w��+1w(�+v֪G��[�,Wg�L+g���t��yy]1=�f0��rh��Iip���2�G��KX(�AW�<����]���Q�Ĵ���P���)��d�6�I�v��ىuղ>�qF�=V��)ǎ�ұݴ�˼7N���V717�!��),��:Ц�>����U�]���]x�.��w{�*�k,V���5�f,@����޼�ʔ�ΈJ�ҕ���QS]d����!�E����	t��R�u,��r�dȩ�:+�Y�ծ=�Q����ޚ̮2�]8�������mݐ��ӄ6'� s7����[��H��b;u��,�����BfT}�ZW�1ݦ����¬`��(��
�-��Dѝ�aN]�{7y(?�����>T����}we❭������6��Np��kx���w�NrI�;�3�F��Q@�.�	�� n$M:�l�t�V
��LFc����Ja����&|���6j�z��G:Ճ�S�lX׫S�V(�X�pX�b���Lc-��snmD��cF��)�"�Z\ϑȎ&�1`�-�ny�0^[�cm11�����pܹM�,s�ႃ�0p!"ij�� �8vC��Y� ��&����d4Q��QMX��4L���5z΢b)�=��LT Lrt&�S�b�щ��*d��� �lPQE1,N�PD5˒�N@��4,R�h@��T<�UEQ'6�Z�(4�j*��)
5�AK[m5F�y�

/,�S�m���M5lj�M;`��Ś�"�{�AN�6h{أ�3%I�����.�I����������b8z��6�kI��T��d��J�F���4�����6KZSAAAT�TDѣTS�d�{[V�wy�5}����2��+=��9�+=�T��Z���{�:���ۊ�>�<�w�m.l\	��˛���@)�#5p��ux�qB���N_��~��yz��b9�uv`�z��C��ǯOC��v��呴9F����推�<v׉�èC�7��S�͂�6�V�u��׎�2�%G�F�3	���P�0�7zB�����<x�0�D�^y����GOh��m��k��F>����q�!3��0-"&9�Nφ�V7�?<�aΡ4L�D���J���O^g%¦�6XތH@=�p��ܥ���D��t�xۘI�L[m9��#��;v0&�Gd�ZJ^Pj)5��{���7��?{E�m�4�(�	J�! G�/+�/�R_UlK�T�9�#���:0�J�kP[f'�:b�nIN��͐1�dgO#���X01�����U�xŭ���鶞�����&#^�P��nr*ځ�!>���OAd	b�x�3��ơ�[݃U-���o"�-�t�`��2�|�У��p����Ka��X�4���)XUI�0��:*��etT]aռgn���S�����q�P�:}	�7	�s>�@�7�Κ[��tK\|�&2R���2J�{�K�������HyK��e���a���x@�|��?O�q/����+����}��Y"�7�([�|(cyL�|���"���+���h��^9�v!F�5\n��|H�BG��m��������{�o�^2Ο���*�r]���R�CsIn���%�#�Z�1Ox�qde��W}�B �Xq�\uKk�G�^���y�P߼=���{��x3��]V���f�8�g�e �V-��O~J�~�8_|��g�8��B0ϡpkhL_�@itE���ꗋ#OM�
�9��d��'�Ͳ.�1�^r��;f�W�ҵJ
� ��"�%Z��������/�oBѾzwR�]P4�Q�4�¨�yj ��/IAbE��KP�03�_ 3��Y�~�%z8)�g����~d*71�1�*v+WX�����q��%Q`����WZ�K݇�/s��V�^�EVۤAvk�^"fD_��q�=#���^�r��5��[qܬ�U�d�E,\0H׹�7o=��2ā����B�%(�_5Ѱ�Gm�0�@����f���+o;�wf6q����0�O�uRũ�E���%(:�ȏ(���������b�xl��-+�~���N�,5�(��F�t����e�,��+�>E���/
����=��>ow'�A�A��2Ij�)`v��
��u������C��ϫ��H�/�W�%�{e��Y~�u#����#2w����{v5�pU�X#`�s�V����3������~�'��Oׂ+�{T�^�'{'I4U�a�1�쬾�S�kE�mc����؞"@�p��s��51����h����':�R���1a��*����:�u��+<�����6���t���ݑa��K[ȔE9t�/����V�΀��"�n�'�%�tEt��{�{�7��� �5GrK�`�*k�:)�zE��!a���Ҟ+�f��mkT�-|=�A���Т�����sXo��sNV]���M}C1P��E�|@�x#���3��Fx�]�>;��ف��A�\��Q33�sa�	�S�(]�xa��a��xs���$n}���@�h�/&V�7uV��'BӃTi���)d3A�u7`O�_*��W����!1����*�����[f?0���Z"d�[`��u�1�`�[���̶�ǢK��;]�2(-��(=��}moy)�O��$6N�a�]ٔ93r�����{����EL,t�q�(�|��9O:����Ը��N΍��U�e��7,M�<,8'�����-�;
60�wGszZ�ȴ�YPX���;=VY̵Q�c.���m��z�����|GH��#�ǎ�a��E�{ME�-�p��J�.�N5ؘ�����y6t��T�Ύ@�-.� 8��a��c�O��G��5L�5�y��nei�j��~���,��Z�PJ�W�q�	�]�9[B���`.y\;k��O���]Į��os�R&���#��>�-'�Oz���Y�����8K���������9-���ׂ�գ�co2RѲ���(�1]���E��z�}n�ȴ;��!�;���l����*�	.7kaa����E��,���۳��s�rC��� ���$�����t�x��Y}ڵ���l���	���3�עfy��HĽv%�6�0����aTul��y��d-�L<�I�/۰�E���Y�9!���zN���Z�`��˟ۇ��օ�O_tV���D"�~a|DX[�LOy��5�Տ�M3�X�`��$@"|I�l�y�5�Lo1�ʖx�<e����5o�*"��*�g���?|��� /�;�i�f�i��,y	�6v��D[M�^:t&>LXc�q �דz�j�>Pg�i���ǔ����`ܓ_)Ivm4:�:����wc�^gjf��!�Sl$n|sg�ǫxT:E;��,:5A|���[��>K���A��f;{��/�Y�yE!)��A�ZSI�Q�a@�ǡoV�^��}((�����[���7:�V��������:��v�p���i��hW��K�~�}4]�tͥ��l�5YM ��2c8^��tVޭ��*~c$9ؖ�ʘ�6|7�#���j�-�i�2yC]�dQ|ܲ+u�N�ElLJ�K.'z�K'ظu^���HR͍"�9��;���HHݮ���tS~�^^H��Xυ��m���~�Ƈy��~E�\*:΍�C���:�=1���O������%]�x������T�L���A�����*<�7�b]a�p�Eũ<�q�y�3Aل��И�:c��#:-w�u�%����v޻=��|.�.}�#��-�Zcz��||�[�ss\��]EO�
�
	JP*�  ����|���R%�l������1����<� 0�o1<9~��G���\��r�d3[m����6ui�͛�[����Q�ܨ=jFמ�	퀶d"�#���!���y�s�bV��B���Vnvd�U}y7�Zo�)�?�a�M�խ|��}C�$X��c����q��~�WT�u�͆uEFH�\�ȣ�#��ݎ�mi�<��Un�z:�I��E�NH� �]e����r�=Փ�G"3τ^$K\�<$×��i�j�JaşY[�'���E{��_�8�N��ΕA̹MO�ә����A�oި �����i�0��ʄ�&��i��^�I8)�K����.�S)�$��g۟w{qԮ�OÖ�\x�HX�9¦DiF>=�B.��rF�6�՞�ȑ-�E=Dc�L�#/�9;;\�]����ގK�G`��Z��u�)0B8-s<:N��m�-��<�}]y��b��{_^����o6I���E�,�Q����<����)�e��7X�"0�������BƢ�j�նv+Z��,���U�I�z͜eY涄��z�>�?���Σy�9^�B��͸v���4��W��N���D�g~=q�E^�Y��g�4�Z�%u�i�xjXM���M��Cd�R���S4��*��ׅsjmd̔�c4��f�?��zpƣ�[�k|�`��{:�Gl>����e#s�͏����{����׷��� hh@��J=���*�F�����¦nG(ǚl��!>���qR���A38�@�����C7�ъ�>}�:��[]�_�+���\fxLN�H�:ɫ&=�A����P�jT+̓X6s��{7{���ke��𾹄�tײ�������	��G.Ѡ�%��V�-�j{�î�-)��6�K����
�'b:m�c�Cس�8G�D&�!p.F\���Ȼ|1Zܬ	O]�T�}���Ӭ���"��L���C�[�	܁#D9	����TF�"��+�%��!�^�<��# o�-��wM���b���C�+�<W,AY�Ӽ�~Qև��___۷�l�A���Ď|��-m�B�L$�-yd\��~JKGjHj$�.4`�Kpn�~��"jK\��rBgdD;ʧb�;�B���{�.�*�
Y��jº���:��e*sw�����³F�L|�0��:nC=^���+۝[���9�Cm���f8�6/��L�=�ظ\d������#[�	l���"��2����:��w(v׈������C��U���1�0%�K������o ��jٻx���VmM�����w�Vq%�Uý�`�v	GXU��=��/��!v_��x77�6�T�{69�b�BԻ�>��F�GBa��F�6�{K�xF[��d�m񥃻�m"!ˑ2�2��  ��(�
1
 ���zr���kp���3X�
�i� ����C��V
��H��r
��YF��z��t)�md\4��Ί���NկH��,Y%�����D�7k�3.�C��W)�5��:Em���������e�'.��i�e���NX/G\�j��L�/"�S^��s���}(�`�.��ڃ��3�Ea��\ M��~6�	��� `L؃�G���aӼVou����CW����s�P��$|pO���7Ѫ��[�7��x��Tm�kڡ_`���&��G�5�bj2���9R�˔��aM�����.ԚWw���(A*<����g��T.��)���p�1���Y��ʩ:�A��,<F�J��8m^*Bc@Z4)������l�**�E+(�c�̴$��p� ���Ӭ�>����鬭��ls�o��2�SW�!)��1)͂��f��B�G�`|�|���J�,��80�_�j����z���e>���H8�8_�tBNS�E�7E2IJa�E��!�;M����Y??��tXb��>G5^����ȗB��)ߢ�2/�Ԣ�tS*Zj����a�Fa�����d븪��D�V!��q�z�hw��]��[��Q��N%P���	X\r����%ɗ�����+���z`��4�r���&go�u�'[���p�&�p�֘�`ٮ*���{�`��g+ˣܓ�3�D9�o�ü�}�O��h�A)
%R�
�"ZA�|<ގ�<MR��%�wn���pP͌����&n��hQ�)�OU��r-?0W�l����(���-h.��MC��b<��,�pF�ק&�>�����o:��K���i�nF�Va޼�Ȱ���*�B��+��� ��ЅH(��C�a$_�|Ap�X��8��'s�\��;U�t!vs5ks#6��>�x���WI���PO��d-��+F�P8F�����T�l��{XݦuApaۓ�X�عR���9�M�	�N�1^�=�A=��Q��@$

���eX��o����/�1Ig�9X��.�~(�3e똼zHz�"m�D[37l�t�V��m�!���'lU�؜X�3e�v3],�c#6��4��C�"�Cz�"6���m��,��n��N���O���O�XC2X�q�Ь��mE�;�CN�^۽�����)g���D��3_��1�]�<�R/&ڭI �ړC��dϘp��}+���N���z���Evn�7�wڀ�;�Y��b�M�,�\�E��}返��Ȥ�b�z�����]���:�J�_�Ï���ε�z�b�R���3qJZ��[2��n3v7�ih���>vU`yt��j<7x��+����������m�V
Ws��	Ie֍l����6���<��\��>�[�A�UGZ��-;��n,�jw{8P+�p��N��)!5u�>+k�>���
��	A�DbhF�"E)�JR��Q�	B�b������\��Y�9ϣGޓE�헟`�ل��&Pd�k��ؔgQ��z��[�z��p:�'y���[6y�5VPd-x��1t<��P*��?B	��u`$f�XT�5ߢ:���Dl��F�˩T�N%�s���x���a��_Or��|�|s���,�:��ɢnTI�δl�a׷��:V����mz�?����N�̞ق�vK�S}'}:$�O$b�Xk�q<'�����QUʋ�1�F��,9�{�}Y ��#�1��ʘ�rs��\�]�Mj���й�歝�>�ƍ�ò��E��<�^1k�ȵ�,3Ǡ?O�x�Qc�;v�_}�ш���$�xo]z�f�����v�/+ kt�uד���$Xׅ���t�w�����1�����Wݔ[�v�J:D�:$Ȧ.L�Q�mao:z�_�ϣ������9���Gm	�Q_i1//:������XG��H������(nuvr���(��VvϫluEi�J���5��m���5���*�#�>��!�g��X~�S�����o�>�m��	����U��[+���]6~���J��wN��n,~)`��7��ro���qUj+���R�Z`-����Rtu�p|U]����*��\3i%����vkk%����JxX�����+�[K�£a���o�%��"�m���[[��Xh�d@���( &�ZZ ibT(�"�T��%J � �xG�ʭ��s�Qa���8�\1xו��TC�>~1��/\��^��={�bj�j)���{9;��J�)�v�"��ZG.�N������y66D�ǐq.9�&uD�vݚ���^�v�mQ�}Z��k���̳Otv����}�֛�p.��l�<�t�A�2�M���͖��� ���5s��݊֯v�A�Y�5rCRFu��W�J��Y_.ٕ� ���v�fl���|P���1�L܄lNE[P]'k�� ���ƀG�Y�Y��6�f?I���;.�^Z���u�Jc`Y�
Z>?T��8�9���Ka��X�i��Zz�X�SR�LY�F&$`aW����Q��s񭨸N�q�P$GC��n�G>�nЛX��rT��v*k6Y�����E�]:�-��H��j�'��=�Ы�8ސc��!�&�J���b��/�s�f�Uߍ�{�d�J�c��L�p���):D�����/@;�0�qa#�x5�tU�3�F�"%�	�Bu�!�/�;H�%=Y3l��\sr��6�Ms����[�x�9����~����>ߧ��~�?O���zzy���}Ｅ_����oGu����:(4k���N����:Ԃ����(�Ҍ�mJ��ڮ�f���t&�O��N]��T�M�9I1��_m��C���ov;]�TZ���,�!r�|�hg��ɛv\�f���7�5�uw$Y.�6s@��WR��4���(��I]�R����Lu�ͮ�ྺ�QKUeo:�[�,.x��.�`�Id'PGc����:٭��q>S �C�gX�(���V��k�C%g1�:�	3i���eb89-B��P����/�ӄ#Х37d�PX03	�&�<�V�_p��ﲷU-�r�j*w'S}��%;�(�7&�RtQ�:���Ju�o�R��P�F�L�5��E�������~��xx?W0��ΓO\ƍ�n˩�U��p��W�+X�(ޝ���N���0b�D�:v�N��Jͫ1��l34�����m�[��v��J#�:��U��<mٝ��2�m��Q�n��.1N���A���]�-�xZT%�7�$��P�xɍbLW�4�qW$K�#oEcu�шV�c܍sꫣ;�KDڣ�nȎ!Q�5���f�A�#hkZ�%
'���ɶ-��dS��~��m�Й��Eoܝ[�����1���  �&���E&q6Oq2Ò�E()7^�J�tGh��eZ��;t�l#���tk��&�4+D�x�5�N�I�q��ǰ�b�vz�^i�{�6$CE���iH�!�i�Řt�����T|�4ֻ��������"nt��]�<�qqĲ��t��ҝ`�[�dܬ�&��;.�7���@�!��
�YOfJYa�r�d�/���M	���}��5F�!�p.<�n�q35:b����oZ�٫u�}��"I�m���
��Pܩ��wWm1�ea+�w�"�"�	*��Ȥ��g\yl���i���n)Ǔ������ۜN���;�T2e���1aK�3� ���p�i���o�1l�74��Y�;ze�Ѐ��q��c:�%n�Is���I�
=]vQ}�*Mn�g5-�%�F]�#�M�+u��ZC�7��u#F�����z����)�U�5#��́�:d��n���Ia�#{�G��K�D��,�B��W&ⴍ>6':m�F��]v�*����	S�[�6��-�C�����2�i��������rj�=� ��fc������̐�U���J���rPW9�q�irT)7y�\%Y
BNGB������Oy*Ŗ�#�[�M��o�1��T��:��}����\Ud�l�R�nZaɡ<<���w.>�+/�ؕ��g0O�V}bg�wPM�r��[do�W�X7��N��6��\��iu.c��ǉ���X���ړ�zo6̭��:�zIf��xnѲT�	����չ9m�%K9ko.o��$�$���}V���Q�(�N�T�h��*����+�3�����Fۑs��ZuF��by�El�IA��SBA�\�3W.Ap�% ���Ӡ4�X�N�Z9�KD��T�ضZIMȠyyrQ�r����9�trk�R�v܎s��)kO$�r)6�P5��K��w��O9�NF�<�Z\�5F*j����W%4�CDJhy�O!�����yQA�B����G�`���@A���l�M [.�@�Xy�h-��a�i+Ks)�
�%1��Di��K�9S�8O"�M&&�JmM߅������{<���
��g�̹>V!x�Gp3ri��/�(�N��cp>��ɘwK���37d�(��k꾽[������^�|z�}��`��R��P��i ���a�)Y�
eZR B�I��#� �� ���\�R�{�0@�T����/%���
8e0� �yc��rRX�GjeN]�m�L�Ⱦ5��a�$K��h����Τ8�/�����z�Y�9��.�*�
:y�V_+}u�^�ce�GN^�9�X ��{p��x�c��Bå���~�Ρn���'��"�w%W�q��E��B��6�F�>�8hh
�[#`��<JᑦD���-W������(����M���&���(����jٯ���L� MKsP=׋�g2dK�ǆ�L/j�Dt��Y3�u�,���w��oK�O��	�.���w����	�v��"�P�W)�#����u��왊���UR �A�y�<ѵܳe�p�d<�= g���T<��L�{W�=�e-{�'ci�9H�zA�\|���'ܬJw�́���������U�A��c�O;C��|���^d*6ܚ��9�L�~"X_|��W��t����y���W��:g~�G/ӻ�m���;n�m�z�PU�?71P���fΌ�q�8� 7���ML����hl�~<�完.LO�kk���5rt��g�W	s��C1P��⠖kyH�F�����C�o v]eS�gb}��^g�'U�\3���[i�X��
���`ѷ��B.!�jS�lD-��zM��&>|�Z_��C�8C�?��!�J�	R������(hJ��J"�*X�)(B��w���|�Rɽ����)�	���B���pv�g�\�Xe&l
VQ=���W��Jʸ�Իߚ���b�1}^`ͽ�4�����RX&�)P�ȧ��{_q���`>�|�W臲n�~�6ǜ1<�x��vA>Xu�����W��{�!'Zz$�Lj����[�VV�+5+I��u�d�e�&�2'��C"��x7ncH�W�]�(�ahԢ�s�%����C��^�nM�W�Flu�(b�:�Y�6��zh��p��S7vta���k������iw�KNY������\�/�t˄�D ������´,;���'~�#���}��8��g]����[(j�/K#��*����ki�{>��#٤A����-\B�?�n=f֨Yl:5�U�l��a^G�b��]+���4 �I�TB߶Aà=֑q�11�_D�{64��].�ڝ3�n>يbDI��'���cя���j�Y�xņv#k:�5qq�Y1��'k��-���?Gr�R��Ě�̐NHҋ�g�$8�>&+����7��Q}*T]�0�~���rM̈X��{��'�q�	�WP_��K�D�ցc���X���~�����ls����xص��K����s1/h�
��.����'��'��n���r��A�lR��Aqn��bN=�q�du`n�_m�q͋��3�&��Œi/W����D�B�*�L)��7���f��.g�f��Wya��*b�m�v2b]��9a h|.&%M��N�k���c f�0���Hw"�cD�� >�e_=K�M�,n�(�b�kؔ�w�H@Aid1�g��~��z;�C[����kKf)��W�|���3q3M��wA��
o&���߱IP��&C
O�vvܪ��0�g��t/Y}؋d�l݃nPeV���$r��_����责+�"��9��o���RG�ޭ��;a�������7�j+Ӽ���&Pd�-)��(�0�|gu���
DB�X4���ٿU/D�c�*�[�y�A
y��N(bY���eaӦo-V�?O�c!�[ퟮs]ڢ��e|�+I��d�9�'.��Wi���<����>1)��i�\�L�e鸩���)�cN=�6lF�\��T.�����)�'>��\�҈w��W���[���R<�C���;��Cٍ��X�:�.X���qk���*�����a����ۘ��X���Kv��um�Z�ƞ�^�n.N�ǝ���蘴䦀K���uL�v�lW�mGy�4=^�G�Y�q���Z�pАTQ�&|��^��O0>�w���bhC,vƝR7΋��P#]GhZ�ǖ���=z����]-��� l�ʳ�
��x��ky�q�d֑n�U�2e�$6u��g/�Ar��Y�����Ɣ���������g�~��>�}��IB k�0a�<�z�Xc���D8���Ԧ��g泰��d�c/B<��M���K˲~(��A�N	������;D>`�V����;u
����G�GeY�=)?5�2m���} �K6�PQV��u����+2�$M� �>	�&�'���-Y[�B݄��Q�����>���c>ĝ�])[Kc"-cce�B��8��W���e��-�hv��3��@�ڶv�*]���Uf�en�v�`�!syN��-.49XHiEH#J1�q�DL,sY+g"�"i��{���ff+�9�؃�Aa�^&h�W��b�.�G�;���9�ٴ)&>3b�pf{�щ|l��3)d𵙼6#OK�n����7g�*�I�ݞ�hs�,���L��i�m��	w��[�F�ӤfM�ۢs��k�Y+�9��&�|�2~2;�l!^Xބ��Hd�cW��q�����4�W!��*9Sw}F���J�RT$���L*f�br*ڂ�!>��0�z K��l����nkqw�ۺ4��g�{e����X�	���|�Ts��o������C�a��g����~�.�\z��)�{:�yx6���K��{1j�����p⒛m��މi�U麛���KF��5!êi�0.�����V����b7b�|�9eN��GvE��qy&*�xI��%��r���"�d��7�g#���H%@�~ڊ�Ք�7b�P�� 0�� {¨�r䦪��q~ò'��I�5.���z�Y�g���t�u0�3�J:��R�M]�wՋ>�:XN|�P�k}Bݺ�л�l'�-�W�N7�H1��A�~ܒ��we:ۛ]�&Nr�ڰ˲>���#��&Y��1�&�:��$�pg׃�[�	܀_Ƈ��bl�����2����`^{ Ho��oeIOW�f�$�ܴ����\�2(�*��.�/V�ܴW"�, �"��_���g�O�>�L*�J�9P����5�X �g��t;{}?R��򾨏� �.|Bӓ�����&���I�X����E��w�u
�j�o�Lo#���=7����0�{��^�h, �,,;$,;S��	�z��hZԡ�b����{6�i�;�F����e���w+6�4����V��8?����i�h�넊���n��߯c��agV��e6�w�k�c�N׉�nj=���p��`:�ȭ*a�m��S�^_!��As���z]��^��t��,+�ėj�2���	�v��-�tg/޿?��n�L�vKeJ�v��~e���F��h��g�-����ᤍ��du�^Z��`ʂ��ʕqj{w�VqK��b��*v�Y��4�j����}h�wyF���j��j�0sA�)����g����A憴�Z���p��5�5aU�E��k|�5�z���>�Fe���(T�º��b�[�w�z�L���!�0�s�Ot�xp�e����� �9v���0���tYs�r�os�n�Vܮ&ݝ���bA�w� y�N�Y���/ ���}y��=����l��ey�bc�`�ٵ�������P�E`^"�X_|�wr��Xglʇu�q�|�����y���;j��ˡFң����E�mz��_�Á�����J2ۥ�A�j�]������Rɫΐ��L_}B��}����T>Uj�VQc����oEl	��Ts��'m/�L�NW�4����� �'<T�	�)J��}7�Ö��'���p�W[=�I�L&�~!��;/�z@�I�1,����m�U)���Õ�.9#ޯ�C���K|��߈������J�/��ϻ"���jQt�u���m�g>ogf�:؀$�2�`Ӗ����Atg��N��|z�P�X�I�U(��IY޼���F\/E���y�8ZY�v@Y ��{|�´-�p�����ᵫ���<3�ӕA�n(��0k��F�w(rE_殷��s/&.��~��}s�1��]Y)%�k���2Y�G�
��3���%�p�R!S#������T{\i�����;Od��4wEDio���ם�L2N�B��PS�o/K.7�Akz:3���6�88W9}�� D4�HP�xx3 <��G��
�����c��+�*��ydg��ک��� �8x܀�<�a��z��@�A����:�o@]
���<��7��V!��l?���]+]�y��%��t[�!�+��{��me��Ko��vH,-
�8E�+�c��R��Y�)�6� >�z&g���bz�8U�\r7,v�G)í'���v���HF0d�w��N/�_��&��3$�{/��(���o�4�SK��Y�IU����.k���m���gD��Ņ{C�q"%M����t�A���0���׽SW�%�n���ݪ�{���x�v��-~��5Վ����>�cV~�WS�W曆����f��d��ݛ�w���,:��5�$�S_{Tڃ#�ai�A	��{��p��/zoIw�+i�j}:�L�.JY�� ƌSd9A�7W�T~@���+@a����Tqo�ߴ�+0}d0�A^)���4�]|G;ʊ�]My>�&@A�U�O~�gP=�$0�����쭽Q�2�O[�9nwCB��0D����հܕ\�μ�&%�M�Ik��쟬��˫
d��^�Ď+�L�s���%
����z��#�K��
�:� ]���/��Y�������'x��Ak�m$�ȣ�9���J ���?%�(v�J�%u��o���Z��v�ڻ�K�Iq.��:�ޱ0ٓ�J�ɋ�ej��n���{���{�f����8����v��获�CU��)ZP|�_��'(G�N�����z��I�z�w9�A����14����T�cX��+M����Y��=1�:=�?�I���J!���3_[3TczOk����\�����QI�����a������}��l �@r!6�<��f��i��>��Z��r�ڬ�5'�aۼrt�x�� �A/K���]4�|z��[}'T�������{vu��E�T
���V���֛��/�ך�w����S}���?G1��y?SͿ�&ᢈa��s��0�-����Q�l\���Q2����zJ��^��e��3jQ���=�����Ӹ����A0���yH�q>U;VV�P�`',����}�	΃�D��Ïe�����~���3�l/H�Єv}�A�t��g�8k��Bk+s�-���G8��W񹓓��_5M���pW���G�����2�ǀգ�ƹXHiENҌ���*��0F�h�h�5��*�3`�m�Pt���N�L�v�L��q��'�DY���4@��V����Iþ��箿(��B�v��m�3���yA×�e���Æٸ�O����[��3��f�ۻb��yZ�:�$������u��zۮ��/e�s���b�j.�[� N�-��˫��S/X��������i�m9o�t+��Z�)�J�dp��� {�����U�޵L�8`�m��Le�t��?[�L�//i�{��n�se���Y0�W�~Q�}t��.̘"^m��pƤ�z�EP!�i|u���Ofeax�W&�n灠�N��oT���,%�f]���s��ث�l��^�����>|Ǧ&nA1�4�����a��e7f.ZK����k}��W��;����N��%�B�X��2�T�F���Yܱ�_$H�r�]��ޕMu n"������hR�)���vOƶ��:!q�y�I7Ba�~�T�fVgc�ܹܾ��Y��؅�S&�:��=��Nm#BՅT��[��v1�P3�������T�:��5uY��F�{� ���u�8�y����t�����-=%��s_���.Z�x��g�㓮�K���N�08jߐ����R2;*Jz&)�t9Ʊ�xs!�Bj���F�]�r�j_��˧r���`��0U���m�K�~�:�
7�4�Q�\��'QzV�7����ɎB���^�ȹQ�{K��RD��k,;���$>=���urn��s'_��G�-��ϔ��6˽�ō������m�X�>.�7�.�u��n�g��,\7dG��"��hya�Yj��L��!�o�l]j�����z����wPrf�O:eZ*9r�uGyEv
�6���\�H���k�[+'�����%aeK�L
�:U����� }���:�0�r2�ի�a>/v���h( �pXvHQ�Zk�:ꞑ������Zb1�vR����n!�>I�5�����w+6�4��8kU��v�gls����4�U�]�n��Á2��K��i0�aJ�M�6�L3N�0x��s�^V
��(W~���������m�-t�c��+~>��v����s�憭�½�$�Q2����;g����2_մ�]Vº���;�ŕ�`R��8����C�|`�Q��wS0�{3�l �C��n�n]�)�f(��N�\ִj£��_(5Y ����b/�_}�Z���L��
�t��2T�{>��˩�_z�h^�k�"�m�W�b�������|�����	Ot5����lH�ù�'�=�.kc� �0�%�"N�]�,ز*��Ȣ��{冽�����7n��
�ջ���3��vTd�홆�nBb�L�Z4)=�9B�ǧu��=���7ΛI�s]Yg��9�������e��S�px`��|�����ߘħ%A`��JT.����^������>�/w�����{�ޟw�������||}xbM�来�j�c����r�K3+NQִʽ{�h�i=��e����8lH�����h���22�Y63-�hiI���jp/��Io]��F�J�p���k޲i6�0�Hn���)�U�Q7�
-,t��%�Y�"�z��7.�-QfE�!|xÖDY`Q�+'Y4o!��L+*��P��oCU
�MӚ���3+�"p�u�*�v+
fF�{(k��NF�nk�mN=����K]{R���S�}��J����m��q�&Kk�K����gV�;+,�usnT��ï9z����H��I����:u3]���q���;\�:tu��WM�o�XE�_m.}x5rk�ڙofJ���Y��e6�^�U3��,��ԷN\pVmY�%�D3L�Ǟ^������wyҲssof�o,"Y}xk;�$�3�5�N�Vh�.�!�:	���تVnq����ݝgX��I���,��AH���f2� |H��u��{zp�0<v$�Fz%�p�����9S3�a�Fxe����#�v�bT��aTՈ�J�]:�B^���7
��c� ѣ�m�]��ԕ�@���Ňs�{UߋXa2D1�x�5au�Xf+�3ޮ����S	��I�� i�YCT�� ��yF��l��wJɏ��M��Mwv��������gzp�Tv�[E��4jt�v�n�e���i���+N�'ή������gf��3��6,��s������ț4�P�W�G�.�-�W��}b�1��f03vrO-�#ڼX-w$�ѻ'"�̸H�)G�/���4��"�����%�%�$[̝6f�����r�Աo��35�k��m��yק��4��N�A�;�j�v�^fݡ g����TNƞ��M;D���T�r�U�*�|޾f�A���L�w-��2��ڰ�nwQ�ՍWZF�klN@'�H���ŕ{չ)YUk0�[�-�HrE|�z	�cظ����v�V�\m,���W/�:�0ܳ[�_q��g$QA_�.긯7�o
�Ye`Ǵ�q��s���M�Nzl����
������������&]C�WKܝ@��ܻ�B�"��1`��N�l��q.6VNh���n2��:��55s���:7l�S<ح�b��wY�6*�j��BU�:٭���.��㸱��h6�skS��5�r��%ے�,��=��c���!J�0h/t��Щ�k�ȭ�m;��:��_��w��4	N� ͔r�b��>����ٶ&`Ť�g�e�zg"��V-��ͥ�����&-����	��nDyj�`كI{�K����f����M\��d=T��4o%��� �"�I��?J点]�W.��6i�ý�ǈ�悒�s�a�z����Z��5�q@�SWr7�؋0ε/[t%�nksd�	�Ȗ���1�pj+�S��e+T�`�&���M\����l���K2�q9;��!,�
���q��d��?�V�����@�5L�um��=w�<����@{��l�:4���)H���V�i��}\���cAM�4h-�	�F��	I��%"�%���R襢���Py#���<�9
]�t�:h)"���!��t�KEj�HPm�]hKa3��ihmI�M�L��Vڐ�bm��1SC��61�!Z �KZi�-��Ji)4��M��H[�zà�ih�(��i%&�h��Ҏ��+��JRkl`�4LkIVƵ�t.������ZBi�#CU�MUi(-�T�7��(���i�4>���,f�.�:)��ZӶ4Q�����>ϧ����b�{z	�#��W�]4�ɂ:k�n�<�H���Z�`�V�ݕu�Yc<=�������%�e�(#\wp2�bĂ|H(�����ET��do��S�QO�<����[@��ʘ'�;��^�ٖ���Lb�մQ�d�;}���y^�}�k�@�7�j�"r����T����%_Iw�Ȣ�,��!����-��'s�=�OI8���4t�7P0i�^HP���D�n4C;S�ߺD��<u��-�W�����{g��!�җ��ii�s�<�-:Д�ݐHG�	�0>O0Z��zJu��9�W�VWwi]�}'��mM�MC�d�2���t;�bwʐL���{�;._fg��i�졫���٦=~����*��L-r1A/t��9���Y��E�~�-���B��vnd�k����X�^a�?4�c���{}6��I�����`����3<��_�����׮���6�Rf�.,vF@%9~1CDO$c��(Ě����}��<���ݷݑu����8���w�Z8V�+h���zb�AݗtK� ���/����`&��7�ude��쎝�����Pt=B��dr�kؔ�����1dϘ�8�0����yz��\�F]�DL;���L�[���o��m������vV�ɯk?u����Uu���)�����D��T�7��U}B�v���P�V��j�(�'��C��CdPѱ΂�:��J�b��������y��x�{�(�m�3�N���}���������?��NH��ٸi�j�KE]+��s�ΜOEM�3�J�X�2s1��Cuai�F�d|�	��_�Ɉ���eT�U��=��m�2�*�6��F�>��'��V��q�_g��9��;k����8�=����z���	l��x�M�(2j����O�u����SI��5o�;?F����8"X\�Cέ�E{%Wg��'^`)�)x��أ�z�\��|y���7qk�@j��O�ZP$��d:`���}����v_���<�p�=�׳���c�D�6�E2)Jj+*0��.�����B�r��-_5�a��8t��x_B<�y�>�{���֧b��"��XsP&0�>G�C�
!��>4<����Y�djѡKb�!���~{/�J�i9	�\����E��9��{4D��O���b�;e�U 쏘\|Q�"�����Go�k�7}��M�=*�q�|��!��=�o�*����֥ݔ���"-�l�@0�ݘ���Ώ�H�5�5��I���4�^�\��C�?x�N���U��\S�%O���>�T e�+���a뷫]�b�9B6��1������n�50��O�M�8��`}�y�t�7�( �<���P�\�+�L� &ޓOw����\%\�������n�kwey\bu?���N�9k�x�f��̵�5zH�"G����P���+s�[.SعI}*�jk������[���g��W�-���;y�i\<lB��*v>��3�$EN
�����O�y����W��k�O�L	;4�E�c��a �2�.(���G����r�!�H�<�#A�B;�ͯ_�s��L���>��#]�O��rB{_*�6��%��1�c�=t�7�}���P�	���Gʊ�ر�O�-=������L��j;�l�k_J3�Xm�����o>�v�Tl������ ;PҞR7W���^};�T�Ь8�0��BWD7v
;͢*�����Z�WUZ�u{8�
�@�~~iw�`t�>c�
���&��U�.��Bd�����zj����t@���q��ҳ߲����l�1pXs�eG �w�5�^�������{j�f�s�
Piװ�Rux�
W*�
jvN5��uB��H�ޅY�eB��2;h�<I�W�_�(�"�t饰�j�D�����j�Q�.�����_����G���3�V9� #������'��n��붴�Ln>n�f,�;�(6�f76=IG��ߎ;Ѵ0�i���zk�o�;�1$���(N*l�έe�h�Lr�"�N�wg�7o�D�l�H�Q��D�7o0����?$��	���sޙ��W��zA�����v��/O�C5)�y��_��|Ԟ�D��g��P�c���-����6jT���B�0��s�d	eWƝ�&
z�f�@��;S��C��s3Y����Y���D��\V�AY<R.uP�����]c&@��~�ܼ1|*��L�V��Wb��פ��:�v��gwf��|r�'���T�|���9�Sr����s�@�b�.^*F'��s��7h�8�=$�����a�a��a�H, �����01���aKǺ�Mi�~~�z_f���Ѕ6�=B�(X�l,r_�闕G0��Mr��A��?��+�w܆��OgF��������أNǨ�sj
T�?Mc��њ	�nj,��^��g9�����Nm��ܕ6�K��Ո��6������۰�	�.�2����f]���8lj�����9��o���eb�R���N\�B��"�#.~/���U��zA!�u�f�UYkSv��/��`�cF���r�?P�	4�P�
ʣ��~30K��;o�S���d�|+S?���g=�l�b�	Ts�=&owÝ;8_��Y"���S�]mOn��מB:o3|���+��f�w�,5cIb^��ζ
%m�c����{�W.��	�פ/m"w��6��	Å���;0�.C(P�k0��P����"�7SG8�z����yo�q�U{��c_O�z�-3[1p�lQ_�P��8����2#ps��ф"��΂=��OT�5���Z�N�]
6����?p���IP�pսU��]�+��V�����(q�>c�'{�KsP|BSm�ޠ�X�4)<#r+|zw_iᠳ����֧����d�އ���_� X�����7+�4�*y���Jca�Js~*K��)P�����#���6�E�^�qf�����;Uþ�5��UV�oO�n̒���$�w;�d�[S�cFbޟ�����[�R���ޑ�O�"UJ�v@ߌ�t ��K,�iG�M��f���{μ2_�-U%��ı�~ڂ��u. R@� ���0编���TϤc�d�4��O3\�(%\������T��[�p��hJQ�d��p�۬J�re���L�읝Ѻ��hRҲ��Yu�V=L���+ITe�?�uu[���o i�T���@AȪ,v�������=D4F?Q��	�q�';6��.�s�y
}2�>]ʩpwduܛ������,;�g��S[zTt��o[x�g��Ć��/6�t��i��2Ҥe���F7&V'J��n�ڭ��Yǥ}NCL���ۺ��[��&S�rhƱxn����'dd?\Aҫ�Rʜ��EI)��+�[%���&�=(%y�oxDV<��t&qs޼���tW�a6�8���ϕg�6Z�,�y<u>�w;��G��ɞdfj\n����s7�e�8�ł��	���)�8��b�����fzZY=���v�n��4����^�u�B�g�W����	�lJP\D`_r"\�(�x�����4�A�k���_ � ��i�0Hz � �M;�O�P����K!�Y�\��WkDF���j��z/\��ӛ�����]+��p�/fگj�Pg����&#�W���7y�pkdFF��22��ǡ>ɜj<�S6�m����#���8��2�j�%���L.�#���]��#�\`K�[G�,ԭz6���7c*+�3xK9}��f����:T�v�U�]�{�ٵ�ti�cݺ�V���$Ǉ�d�� l{�M�`�d���A8�l�٦IM;L<F����UUZ���=�=aӦm-�g�VSS�J��.2��K�eza0S�ƐA��KF3�L�tJ��1㳑m��l���^�tD���E\�3emF�_E�z�bA6d1,��_���	�����R��DM�N�y��#P�]�Q5�SZysYyC�����gvm��\p�8.�j�P��3����9�Ů>׊o�F�K�Q��1�za��7�GebwԱ<����L�@:wkt��fZ�)�kr��1tp��v���{.��T�<����u�I%/{2'������6�,˰Q�S��T�v��P�)-���	�/A�y�h4ctpq�9�̮�|�Y}��t4 �!6И��;�Z��P�m�l��1i�by��>Of��p�	d�޷�f��\Ȅ�����80��>�4�N���XH�қ[���Ն	z� G+���ø�����d�c�E~d���M
.�T�cPMc]��������Mժ'5vw
���X�����W�n��I��
�H�v���q>T$×�MWf���=n�
�3{�f���F��^��V��5H����H��%��T8C,�+�����P�н�y�n&�̽�������RN
c���p��+MZ+�G6QZ��ob���g��8�W�wNN�p��ٸ	� �����~ys��h��1v�e����BG�_*��t�T��+���ز���$�A�T.���?�۱���}D���D}� ����9�D�n�EC!h�.>y���s;�򣞛�ǲ*}#@�b,�W_+���m���!�6�_B[}�nJ��:V��Q�=9�7:�ۂ�0ՍR:ɢ�Ϯ�,d�/N�vU$����6�1�4@��^�K�,0����8��mn֪��)��0U#X���o�#����ǚ�)VHw�Q��Okx�����s1�_��͜(�n��n	�a��� ��C:�gw�y���{�iY��h�,�)�r����3��,	t~��{�a�K�~�!Ե�����cj�|`��#�,�,i#Z�F;�v׫��I�����a�!��9�ǘ��N�"-�ꋹ�߯�Z��~م�N��Z�LRuc�J���n�T\�k�H�>,��ݮ�t��V�g/c��]���J+�&��頶|�tK]a��nêm�#fȝ�,�����d�����w������hA�ZH˔t��v�wR�� c1C�J}H���/���}�^g_�[�􈜤ȭ,}���3	���5m��t��~���t�e�W_?G�M]��\c�����1h[ r��w5��ҵHAY�Cď��J��9�dI�0�aT���8�^c�=ٮ�W��X�T��������*��$LoоR_�glDw�j�O	���e�ww��g8kCݝ�C�}��`�E�Ύn�wXA|��6��@�������۠�B�_E�4�\�ށ�������	��6��x�7�ͺ�#��a�r��r_��~�����״�@}uV��������֔��FR@�W\u�Uc;Bm�4�{;���n清kݚ������W�N;D�t˟�I�ti6=2�<��{���˻s8��*�6�cE����7���y����F�B�Q:�����ލ�D&w�Gr���hRR��J��B��}�|=Qp��ﲬ3������Ƙ��N˷mv�aͅ)6�ۢa�v��nj=�!�Q(KoW;�ߌ]�W�~�"X1^���omu�r]�uc7�T3���.�2����kK��r{5nɮOcβ[mlgO k˹�P�^D<���ۜds���^i�0��Kn����j�Z�ڞCt'�AS��`V_�)A�&�!�"ˉ��I��Qx��0��j"d�"s2z�S v	-W�Az\�(r5�q����\'[T|#��,&��l��&'Y��b���e#&�9�Yt&��u�ʖƠ�HZ��e^Yt(�'\?oN0���sCb�u��u�-g��VgW�6X�1�@��آۗ쁖Ű9�)�Ґ�W����r�������ȵR]��b�*ֺC.��-�(�â̴'��07��pW�9��	Lc�bS�I`��[Q��.�J�ܽ�3kE3�CP�����x/L��Œ�&	�v4$_�锝%Ľ%I�H�F��r�u⦍��<��E���"�ؽB���j��a�ȟ�D2����ȗ�O�����ҦVY7nf����D���R�O,|W{~��ύ��M"r����W�<7&m���7����!'�:��Z(�g�/&Rt�
�q�mt�T2�m�<	&��+O��.���i�4����WA7\��6kb1V�.��]�:�qS���4\�7��w���F�}��b��,9L"�x�E'y�htu.4�8�4g�8'�1�v���:�z�i��1�Y���:�w�vWZ���-:�/i��~hJQ��g�#�z�0ن�OU��\����령��C�1�<��Ù'hY*L��Y�jº�Adi��ή����xa�@��h�m㙷d/!��)�ǡÝ[S�G�j��w�^}��Xn;�ҿ+�eQ�'�L�ɭ"Q���}����z`�1�,j
_�o$N&n>�s�Y�͗b
���x�|2�\���5_�/Q�k�I��3��~�z�E�|�O@%h�|����|�u�w0�F��T����m���1G�{X��C�+���"��؄}9Ę�_��4��^%�*���cUt_�?���yft}��{�^M�����$@"x�v�Ia����yoCu�"Y�--��E�]�+U__Kwe�4�C�,{�B-*y�C���D�^����1Z�
E��T5M�=�~��5Pg��Z���iMM-#�i�����s�ܙƣ�S6�R�a�O\�q�}��O�����x�}��w��������ޞ~��{�O����^�����7Q�]E|'3ëex�BE=ƦL5>ଃ:죎����iЫ�/o�ޡ���f�X�ܭ�E	ͶOo�)�;军;Y]#F������%�n��n��K�u�_u�t$o���#/���1{u�4<8y-s���İWEv[�m�բ��룗5��lDu�/)}��И� ��:�V��}tˉժ��E�ۮ�%���᪪e��P��H4f� �J��AyV����2e�v>n�o�� �Wd;���亴M���Z�%<�7����<딳��QU}�.B�Ua��e.�x䅝{Ė�&c7H��;퇢E��J�����k­V�l;�[�̰U��7�E��93#�Yt���Z"V�/�8@>���A��s��v#�Z	�[B+㝷��H�H�]���I���ͩ1�Z'I��#b� �\S��E�[X�L�n��Pt鳡�QL��w{pɍ_gN�Jd�x�B)�ZJ���U���S�b{�jŷ�D7@(�Ħ`�Y��m�2�ԥ�L��Q�z{(ʖe�
�̻��==����l<Î���f�CW��ɇ�G�J�+�ջL��������hP�#�qѡ��uq
͓[��ieY�{�������7�Z\�A�n��GO',�n;�|	7L-}���ɏfh��Y�R:Vl!ufu�d�b-t�8�-9Sp��΀j��)ېV݉v5́���Ħ^<����C��I᮹uEYt��W*Ϋ��,A���s�Z��Ya���"�����5�V�+�R9�AK��X�.1p���5N
r��L�n��3�Fpf�w�����o"�9atq���V�e\%���&�ݍ��/�Q7+�Ne���cPMm"�LeK]Ϣ�vv�ŇV��V��2sv��XtcP&�r��ůKZ�e�u)���s]��'F\�0v�e�H�(��)�)`Κ1P�T���.-��g#���_�Xŧ���^�Gb�]��D��Ѯ` Qq,����gk띨�·�R:�פ��jOr�Ac�c����;F<h�0tT9-�(&Z3�i����f�>�N����tѣ�ش�KF�ն��R�(N68�FK��ش��5�/��=騰�:Y��]*��Ƥ��cN����c0�w+Ƨj[֩vYλ�4��H�w}|.��֜���T3@=�=��VhuҫN�e�{�E�c�vܧ6R��}��ˁ+�lϋ�`���f��c,{%��46OP`i;�C�7k����O&�Ʒi��h�(��n�ZT�]Cw<F����m�V
�# ��75���\q���&�z����Z�G8��3��)����Pq�v��Σ�.=|�
�D�X��t�#f;KN�5��[���q�{v#*L4o��������Wp�'<{gaJ��;Z�2���X��4��e�O{	�:Ѻ�nf��ۛ��j�m`0�n���,��x���C�.���C�jma�h���Kl�[٠�������%:�ڦBc4:v�Bh�d�ITQI�Y4h�i4V�/������l�
]&"�#lh4;jJMh-���Ks/.@ZΜME	��ոb&��2h�bZ*�.H5�]Ul��8��I�Į����4h����)td�kN�EN��D�A!�gڈ5�Mb�<)������Z�h(�j��h�'PѶ��ɧc1kUc��c��Q�͋�ԛg͹i���f�v�Š=ƨ�A��Z�'��F�N��lkUZ(6��bs�kE�:m�I����ت����Ŭl���3ӈ�����f]�,�a�����5MoG,����a]l��G���	��ڦ��\6��O^��)�[�o]�4��8��齘����{�qI������Uj�I@�!f,g�Z��==R��ci��7�'�l{��~=�����PYf7�^��U���~#u]�3J���#CH"H�����#�}.�ˉi|X;9�k3�Smn"9�D�紌�+T���Ŧ�ya_()ZLA�9�NP	�ۗka�r��{�Y7��Q-6�tK]~dQu��6oѷ:Oʡ=^C�4U��uv����4�8�0C)%����'��$����`n�N��5��h��߾5���B��Q}�f��vF�
�C���b��ϧK����L�ƻ�5��H�T��#v3^ӛxZ�Y�.'�oz%����0$dt�a�B�L( <U��Go�u��QyYXː�a����z�n���E��_-Hzg)�#c�X�]���d�ά6ⅳ�McY�Ւ�@�/�)�oe�}Z�Uᯥګw>�uT��*H�� ���i8-�"��X�+��a|�9�n��2&r&.�s7]�n�>I`k��Y|���>����<����H�� ��-*8G���������jp�X���[h�H��l[-�ORꏘ�˂]ֳ$��^��ü�;�k
����kM�(�\����K�vhi��w�����Fo2�����<�β��[�[��7���'GJ^��5p�eF�U� �H<#U��mM��0�w�7�.f�۱ww�}��x��\�/�a�����4���İ$8�$�sP�c�-A!����ٌ]�ޕ�G��/�0��l���P{yÝBk��j�2�Zx�w����>����/�u�5+v�|�*$Ƅ ��p̈�m=�����t�/,�4��]���A��w���<Wv�T�'c��lO^�x�"��`P&|�c��E�j��׻Z��A��
x�7�1SO-v��#��7S�Ck/i�����f�?bW�9RV<�{������TEzf�*m&�o���x��W�d�{��l�0B}k� ����H�3�1��kˌ�6���Iq�U���9-[J7;5����]t�f���T�`�W���dJ2�0���8�=�����-����'�5�����N�J�*��?s���Q�7�Κ[��(k����|�p>�O���a͔��C�L���HmT¦�@)���<���{�!����{��R��1����E'u]����K�d��B�1���N�o'r Dc/C��&��!�_v��RS��}��oD�Nϛ�1�vr�R�+���0'�Y?9V��Jl�f]����2>�v���_˒�B�sE�+h�hU�����l]wX��7�KU6�M^�G�sX���h��U�J#�K�d�,'7��\�ڂ]��u��5�H�����w��^��`D���`� (v�UW�,Ux�(�0����X���Lo��\�� ���$x���kvzD��r�����N��Q-ќu��s^����r����s�"CP�07�0���<Y� 6��@Q�Ks�oc	�����uY}+��	�kI��U���Յu�<�Kݭ4+Aa<��pV�N�(}������ݔ4�**vAm�ڨZ�a�b~ke��w+6�4���M���	l6�lé;�}�׮��<�s��v��v�aͅ)�'�{�4�R��,%�Fcu#�u��{��zj��{B�a��h�"FZ۟�Ӽ�G~杻�y�"��/��9aټ�}�_�K�n�lB/0E���>����EB�*�Y�5>XE=���wBC���C^�RWod)��=�6`v�E@A���i:"�s�<1̀̀��ˌ���I��oW'�Μ����sD��|eN�2Ƶ��-���9P�C�|pU�|��U	�(���X.o%;�Ӗ�:�%��5�sQ�]~��lj�2��0�*.�J�8}���V3��|}�[�--L�-�	;e�ۯ�e�f�%���� &-]�Y��2�|��cf���bՇ+�z���Q��Q�_�i��$W]��g�,�7Ue_8���8�Wֻ�}5>��v�Z��:�J�8C���g���j�W!
��P��_�}��ǲ#��������i�8&0��Zq�w쪓�����d&UhФ�%�}q������-h ���ϻ�.��wK����oц��Ɛ1ħ�p����7�y���ǘħ1�w���~֨����+s!ӛB���x�R��o�X�Y���Dc��c@"o�z�u�c"��n)c=)ά��k�ϡ���(;��;]�2��>]�5�NA�N@���T^�<x�~��g�]��GT���"����I��v:ӹΨ;C��q��8� ��	�˴S��=A���u�Х�0)X�Q�4��Q�]/^9���PXחJ��'�`>��ɠIsCŇ�V��Ux�(�~^4l�F�^�����Sdq�Ǭe�&\���5j�w=,���yF�m󚻦�QW�:A_���!�:A=���&�;U��M��`}��[qܮ�~��gd��JԳOU�\�[tP͸���
��'������x��U�s��Xgɓܔ��y7u��yw���y������/Ͼ�^��Qr8��%10�#��NBk@�/nҼ�h��;���U�mn-Q�QG�yK�m�u�_En�.�A�&��1�i�k`p]Oi�����3,�������}hW�5�������.�k��CTS�9y�i�8;��燔����1�eI��Q�5Y}�mWa!����$}�2�3/�2�Y'_���/����LW���㟺�GܚT?�x��g�.���a���2���̮̍�Un����&�ͬa#���x1���G�/ؔk�2���t	΢f�D���c$61�C�o=��{=�1���i�j�3�	U!�%�=�SO�V�5W���]���)IQ�>2k�-����75>�zܙƥ�S6��0���6���6c�«��%uwm�յ����W�z��}�OX��{`XM���OP�X�-��o&�Cԗ�F9���:L�$�ҭ��G��{]נ�
��րT����%��@$<�[ ��-�7�n�R������^�$'<�K.{	�V��7qk㦊k�V��C���M�����T�6i����otLOoa�HBEh��|mj��%�G�5�"|I�|ݳ�]P[��\:��5HY��������oQ������L3j��dvK�7�]�wQ��򖹳�)��)�Ǜ�j6}�z��j�^W�s�PhL `B=��O4T���4�W���g'�;����܈��_���W��LW�G4d�>�Ƥ��'Ō�e�1gꑏJ�Ѷ}��b��>��ot5��Վ�Nn�ګTv+�Z8ib#��1��$�q*���v3P4�\��p��S��ncq�Bo
K.u\/���Ӱ^�4)ך]w�D�;�?ρ�zI�O!�S���n��(O�];8�"#�ix�el��k�7c�Yy�u�zVY�����Y8�l�^&z/���蔎/�"��$-�>�Zީ����AG��m~�Έ3�۶�5v��CM4,RS�_��0Y�d�yl���nקD��� ����V!O��S���ҧ�{맹���~���c���9do���;�}[�:s�2w�z���N���Ƞ[�!��ff���n�<����˞���������C$��s4���=����ߝ�c��{xM^tl��\&JΜ�|��G�k�}��6 z�f��ޏk6��3.L���o�T�o�O�*�5�&__ݺ�>��0-M��## h�昘)��N6ۜ�E�f���]��;����2�g�#���P���gMr��ZP��iH<��,"�V���~N/>����O��ͳx%�IR�������_�k"�Hd�[>�f�2��l�AʒbǾ������wSo�B
�Saf���&�aS�V�T �Z��&�&8��Z������r�3:
�g�����_u~o����ՐyNwx�;yL�"O.���]�E�:�qw��%�ؑԹKF�� �����2��	���{mBʦR��e�+�J���:��E-�.��$�����nA���5���Rj>���WL+9u���QsF�F^l�gV]�(�l�!%A!Ha?�׶x�ۙ��@o8��.;�LM�O�αj0y�?B�������#^�K�E�ߧ㲪Q��^Kf��Wv�ڤ��a���z���7�ߡ��i^[���-s}"�:�и�_+�QIntPa��ͪ�S5��������r��.a	�.�˔t���~T8�˴�S��QE��A�ngdb��ELZ��� �3���-ᄏn@��i�!.���؃?`��#����l7=�R�x͛�G���7s��4��������X���HAY<�<��J��j�n&1j��N1��Q}{q@#\¨��I�w�/�_9���*e$M{~���<Y݌:�L���=hه[����c��b��7B͇2qŒ��!gN������a���Q�[��/��Ծ���|��l����3ƗS�4��OS��m��^+�r�`:�"}�bu��w��ے�2u<l�<���lְ%�`���%xy�,��M����^#�aJ������vhȭs�)�P;��b��|p���Zh��H��r
�C �����E��f�;�}<Gyyz�qzR~�!�AzceQk��Un�w��4yz"|v���v��.��yi��y%zj���5.P����"ի�p��M�_#���J��������9���0׳O
]0Ӗz���m�IVu�!vwD��g"Og��7K8%n
GVU-A�����Ҽ{�y���ؿ�~۶�����G��������|<ăC�(S�j1��스��<n�]�&�r�3�ޯE"d��<��I�ʽ�6�ƶ6�{.�Q�n�3�볣�SQi�lkH��C�U�^�W!F|�q����	꒥���ncr�+�XiWWU��&�,�z�軚/�Ҷr�����Z�]J�D�	Q�@oN0t5�- �Ƿ܅٨tT�~J �x����i�9�c%�U-�^~"Sm�d&UhФ�}FcH]�;e��p��۪�5{:w^�*�E+(�Y��&bF�^�d^��?!)��%�6x�����U4��=�#���V�o�X��P��P$8��� �^ �����&��N�nu���g[3W�*d�8�%�t9喆�2(-��)]�5X��:	�}�z�C)�����L���U�p6�4+֫�N��"�����o�����yä�p��=4���mػ��yG���]��L�#!q�04���B���iW���:�U�E���9��˅��	G���;0�U_�D�����=��h��e�⪍tţ���*����qJ��ޮ�#|7�����P�.�EN�(<�y����{H�m���9�I��o���삺s��$NS}93�$�����b��m�O��`+�`7�t;2�4��x�=��V&cN/S�7�C��u�T[�`��1�%�����NH�%Q�X��h�]�ᕂ��6��AD,3���lQb� �PB��9lx��ldI������*��,{�vp�LF�Gn��ª����O�8϶�I�B��� �@b4������#�/��l�b4��1���/t�>֝b����>�z��W�d�ܨ{�ttr
|0C�0�ܲ��<�L�\BӺt�ˊ���w�3}$�Yx���	;Iy��-�W��D9��wA�	=ת���ESe����9�S�"jV��z3_�A����ǜ��4�!	���G�E/�5�k�����}�Ù��X;:�V�¾����MY�.��W�wP֑������]+��p�:��6R�b_ef��������)3��J"����X0�}~��8&���C�g��J�������L�����jxjR۸�����^=�A�6s�i��������"%|��Yu��k/�#y����M�mL�yݴ�W�6�(1j��4���<�B�Z~Ukc��08E�=��~_��̿}�}�� �qu*�#^X��NfDHr�M6/�S]�h���l@�4�N�1T#�:�o�"��Ɋ��.���0��R��m�W4�Y���;�7��Ƒ���Jl*	��z�'�Li�ݍ����Յ�s��Qw(��f��sK�t�����s�'�����@��U&�B	�/����ղ�*T�ߢ:��ʇ++��Z���]�	���w��Vb�8Ӵ�ơ�!��ƐD�̮T�%��ˢZ�{"����6lF�頾�k��a�8���H������x�}��>�Y��?y-����D}�^�$$��mR�1�'���=���C�ٷv�ofVm9�����LY���x.�Tƃ�3��\��r��q��t[Z��T���a*�կ��[i��!׻����g�E��k���"��c+f����M��D�к���+�+4�^^�
�y�Rt��u3�CptJFG��!�[�a�jz�s���: �������V��9���;�͵!�%?5�i�oJ���U,�C"�H��dP��S�p3�k�3��v��9�͖uE'=S��зa9do���[��V�U���^�	̂��]:V\�<�¯�n����Y��&~�S���C��~�)8'���
��	��_�9j��xn=�f71����øB��xrd������-�m��"t���D�1n��=>�g��������{���w����z�^�_����F��}��Ԡ~�ʾ�FË�����|�ѽ�� ;�wuu�W{��S�M[}}n��absZ�f ��u��s�/b��#9d�i:��.9V+V����#�K8�S'(f����o��PF��O$���{>θ�!j�wim��z���Rs�����:%^Ct{v���&�~H�����N�tP�������]��T����vS�����}e�N͙t�K�q�r��H��2����5��-��i�x��/o*q�iZUc����R�aTG��Μ�5�	�O���lp�#B�?p*�N�p��n�5.�î�r��M��v`d���&J7i8�X�1�iեd|��D�"ἒ�JNj>P�S��p���vK�;y�Qwz�E�C�m�\n&~w�U�t�n{hv�~��[��S�Bc:u��kg恲ɿ��[���p;V�rTaA��2�X�'c�\�t�/Lv;�!KQ��C0�O\��<���p'n�NEX�#D���Kp�����m,��ۆ��m���D*��pבpX�������k']�C���������mMS���&�T߯lz��\�4]��3"*�<��n�wt=����[..]\)����1D%�]�o�@�4�@�oVUh�:���5'm݉��(i�9�-�8u=N��:l��\;w��7fb��t��R����2v�zg*9�c(m�L��F���܋2sR�
��lЃ�U��|A&l��&�m���e�%[×����_i��,Y3��E�lBj7`Ѱ_Jæ�~)�&$͸����w9C���tj�C�B)g�ٽYJ�(ok�V[Ra��M��jor�4��q�c�˕~��2/�2��w���^gc\ؐ�6ng0-�z�Kw�����dt��)����܆�ˑ1Ku1\!eJ]\t��K�yӓ�r��q�Ǻy$�C��׏�JWVX�5���Yr��wD��a�r`WyZ��]���y�ǖI�mdl�∞�wQ�1e�
�����E�� Im�s&�1��w.�nPʽ�2�YX����֛��<ORV�=��1�o�w$����ò
�g^D��V�����Dm_:�e�nAq��9ʵ�5`�2	2�m6�2..��jE�5�rr��7]��/ SR&-�}|JX�$W.�]$��X��C=)Dٌ�����G��Nu��)b��Գ��5�$WOE7�C�0nf�Ϩ㿈���P�00���� �}b\�z���HbSN��5�w�i���5��3;�����itb����]
���1�٫�
3��e���+5��Hq��aꝒ�M('ױi��9�m�x���]|�탦X�xŧ+^��7g*�x:%E�����э�87p6)䷅t�Sk�;$@���k`=<�,��������b��O`�;"uk%�a^Y��﬜W.Wv�&D���l�(A˂j����w��ѓd6*��*���{�x��d��fwoww:0�l	��i���dَ&A�AH���FK����ns{�/{��Ly8��Ψ��V��m�ESZh�A	C��RS�ٍ�l�ST�kSh����X���b(�l&��hhh���Z���QAI�f��ƍ��:KlHm��P�B�h�M�ѡ���mm�[�%���[�*��"b4��>0�.�&�"�5�&$�����6��%;`�l�Q��i�N��U�ӡ���*i��"&�`�$�:֭�+Eh��[U�DjZu��`��4�Ӣ�V���DTkcZ�^c�ʝ-&(���X�X�bH�
v�RDA��Ef��6T�ED��f�����kA%O�jg��U��E	Q�Um��:(�"��[U�nE������TE��i֭�b���-@DIQZ3LUm�֊"��!�6 �mUE1؊���9�^u�~Ss�w<3�5��S�(@�j���Ywbu^ɍ��D9*u�*iޫs��y�U�ԋ��[:����A�H������s����4��C����R����`h���/�V�zL�W.�ٶ�~9��
�14�lg�B���Q{�gA��dZ�mV��["��`����6E�/sW"<��d�l�չxel�����2v�� �!���x���5��~+�/>�e5>�IG�8!'1��i�\Ő�6TM�(�=����F�8�N8�5�Z0�>���,BEn��e�;�z��SW ��HםqO[s�_oUeB�8�bu�Tk�d��u0_� �i�ϗ�S�O�["ͽ�ó��c�Tɺ�T_]����]N����J�"8� q�M�m��J:&�Y�Al&I��Jsa#Bն�(�*�J�(�͝�w(c�l���g����Ӆ�VNܾ��6tö{��&W�D��SY���犚� ��dW={�4��/^w�xa;�#�!�!�O���|�%��pY��2�T��F��Un������Y�G�u<�X} Y|��4�y�FP��^Kw��� �L.����5���Z�s7������Ia<J�9P��<z��!��;�V�/�G��쑥��O�R��Q���&��&�d��=����Pbf���d��*r�G�U9o"_>�tB�3�)yߴ�x�Nr��Z �1r����gK늹q�VLbu-
c���,ں�KOJ���1��HL$9�y�?�le�@I�)���^��~��'/?�K7��κ���@�I�z(��R(���J���gO1�WZ����g=�s�u����M��q��3������"3`8��'di�ΑL�8ԟ�k�PK�Z���Np`�1x�:��xor���o��Lm��B�%y��3�溽9(��nW��>���[5�]���~�3jY>e��2�6����qTx��c|����M�Ac��OC���7�l#�VK�N���tՄ#�����ɜ�0�dnj�N�W)f�z ���<�,4MX�0�)�$���H4<�O��Ϛ�u�i2��E�͋V�k�3��/'�9��X�Ҍ��]{bmA� ��t	}&X3uME:�P�j��l�v\���p���<�3^��lkO�!���� ��C���n2�5�	���o&w�d�c�{B*�}J����d@�.�~5鋚�bj1��ӕ-�Cǔ����`.���挍!�E<��u|�rIϭ���?}��(�1lȟ�K4!�f��~M�5Rt�����V���۟������&"�rb{>�w�9��ʭA�e��f|В�B`$;'�6�<���鋖�]e[P�ϵJV
;@�p����� ���BD����uY�'d��^"���&����;6$�*����+P!��,���<�a�{��ʻ�Cѷ�!����ԯ�dw)�{�G3&wJ�)���M��]�+�B�",��x�WA���j2�"4�뤐��h��*����+��+�5g�s�!�Ȭ���Xr�5��_%C�hN�|�/T�!�'b�D�0�s�|�������s-�c�K�Ʃ-��W���!J�<U�Ky����^�7��a���q=�gJ,']	rO�4�꾢�#�ɑo�_'�أ�� ;@tu.4��B�emW�cը�UN����#�צn�2$�N�U��E�沠��ҡ�����A�rpd�x�;e�[ta�)?U@W ��x��hXw=յr���`[	���ˬ~�5�	���\��j�4h�=9�N:`�sӇ��8F���D�N	ɣ�������`s�l}b�^꯵m�mv��\���W��1���TB��(p����'7B9�bܤ\��j}��O]��b�/}:܂x��6_��N�1�Xmߩؓ��j �����Ւ������Neu\�oi�l��Եs�	����-�^=%� v׉��tE�j��g�]慎pb�����e�A��H�Se�N�k��	��	��!�Ǡ��"�&��n���������r�wK�S7y���ݍ�,�3�Z�nn��pb�<}pZ؋�XQ��N�x,h��	漠������W]��d�&�4�� [����fjTyٖ*շ}W,�&��t�F6ui�����B�끫��/�	�Z�Ü���s��3��.�����[�>�0xc��ɐ�����{Gul�2�5�Xw*�DZ��(h�-*��$���Kêٲ�5��"Z�<��"�ZA
H���3�q>�~ȌnEfu�vi�#J���m�8vM�V����LSdo��3g�=���H�x��=�#���FG�aM��\�eaa�4r/sW�DJm�eM^"Kג3�(�f=��J9}h�p.lD�pl����g�U?��7���8���� ����?B	�ϕ��� ��
�k�^�e5>�*`��-�mY�U�^�����j'��F�ό�/eꥰ�h򆹸y�t͕��G��5�4����ک�P�yّ�L���.Q�5!�ݧM�1K��)^:���bK�R ��G{H͞�V��њ�#�b� s��"ymz����;�U^�G~\\�~�xsM~m�[Z���*uQ|��- �yG��N��VE0�
<5�(/��:��$<��Wjg�Ls�j�IO4�Bc/I����:%#�c�3OT�gzxx�d
W@��K�ux��Z/���閮k��lP�W��h�F�^�6��8��K�O�7lh7I�/�KD-��]A�Ӂ[̜(ސ-PbU*fk׹�� Z����\�\��A5�:-tP����ʵ�+\�ԗ�H͵]gK��*k�ն/7v�2���c��I��*v����*vX�J�]>����E2�B5�vzRqK:x�*�a��l�6-"^"��;=�4��A}r����vP�D��mP��~[c��[�呴�a/��^1���8t�Az�P�qƂ(���L}�yo����/� P�tȄ�5BrY�dw2��a?M0�K��&+��+*��w�:�bi�;�5���'jB>PT1	�������2d�d>�s�Q.y�N������*_���y�B�ʵYNrD�� ���J�ڿ���mNI���k-S�DOc&�KU�nGNVf�f�1I�jHA�v�ִ�9��=�c��|�ջ?ynfن����\ɜX6g;�6-{P�c��8�r��N7�d2Uy���0-�^G=;��`=��Í(���8�op"]z��(o����k�6�BO�xa��%���g��qp�wi��	3F�^�.�*3|!? Ʊ���=F�a��T����	�zѡJ�*�
mM��8�N�;��7g.�j��J�Rh��#�Òn�G>���þ[�VD����z���ˍ���E[�Î<w	w��D���2B��.
gM��Ȉ�n�{ɉ|/ ��Ƨ��9/� KSq����5cV��b([T6��
f�m�k�iRԃ��Y7}+`�ޞ���\�W6cW3*���7��ر�9B�Y�36�����y�����7�:L�-k�0n;/�t�����/�@ׁ�m�����7[=¹)_S��3�/=?0\<��i��b�%v����"1��~�s�`��0�g+m�t^N��QJ��eJO`Ⱥ��2��7pv�z�$W� �Upi\�V��Cz��xnb�!B��a�«�%pyj.Q{J\�O�û6�9�69U����
�έ�����A�j1N�>�q@��']������0n�c��a>j�����C	�����EVۤ�(z���L��v������P�`'/��/����s),��2�����l�^���at#KU�����F�����s��)P<$K17�=V��/b[�������ޘmd���+zzW�a=�
Yk�dD�D,��:�qN����l�8y�s2�3�LIv�e��虑)p��:�Ӧ�r��������m�UQQ����cn8��N����,��е������H:"�|5�� 3/{}^�g�]s]���mfީ��+7�-ة^�32NO`T:a�&���ju�и�mk�a�R#KkTh�\��b�kr��'g2�U�P�T����,fZ]�<L;31t�9�]����}#��W�r"���(qQ�KLꭏFI5�ǠU�����_��Kạ�_��v�H�-�(8
.�Y�צ~�~�P�/yp���Z5�k-39a���)\��(�4¬z�H�x#@!�q".��F&\Gm�5���HZ��eAe�7�j�<�8.��z5�n~�{'���V]B@m�tS��߈"0`��?4#}0��j����2�%3\��X��x�����nvH�^NI빩��g@�,�bE�XD���e���k�=��m��7K���D)J�&�m2��p u�H����eL�6�V���h�s̝��|�E]В�%�`��y��o�-�o�f���c��d�ܻ۬�����P����n��h�F��x�n�>��ݛmȔ�C��*b޽mU�ʸ�����z���"}���ޕ^�M�Ď�:�$�#���1�^�5o��}O����)@`q�m>g�ߖ{�3�VN��a٢Ŏ��יY�ɶ�s��x���2���z-��Հt�^�w�|GG�S;b��95E���J[P�5L�c�t�5�[�TӺZh�#Z�ȪfiSR��rg-�wP�0w:i�3���X�*~כڲ�O^��S;���V�Ⱥ��]6=�L�xUwGP.d{n)�c��Sh���p��w�Q��GK�Xvה3�*f7Gw>!��>����(��T���[i�}�b'�G���x�T۵�=F��k���z�����=�{�����:��Vܴ�_G�VBq�wZ��}�72`�Y���d����{�yt��rw=���u'�EdX1Y��T[�D�7`<U�W�Fǯ���A#���!��!�44��j����ITS��3��0��@�ͣ`������;�N�:�d���n�V.���1����g���Rs鸞,l@�Ѫ~?fͅ�_�ݳ=�J��C���zz g%����hE�G6�K-��P7B�0�r���H옲1)�UM7�r_���f���%*㤞�G�2�Ȱ��[�s:�s|1��MEunt���X�h����q���y#*�95���j��Ζ�U���o1]�몞��o§ы�ۍ���mH�n��J�E%@/o��zz�p*��_���7u\q|je���CH2��yj�rf_� �4e>�2��v�hӄ!ϻO.B1��<�Cޏ�&�&��̛����������ܕ����_9E�f�f��KY�ˑ{�]\�oU-��U�T�+�������dg@^*�o�����M!����9s;ϡ��f�VK���� !p���Q�ڦ���Z��!��:*u��r�sxT�����p��]n8!p�-~{pd
��}�#�V�D��S�7�����+�s��*}��v��`9�"�GI�7vZ�tSڽ��{k�^c�#<�t�����e���.��7�;��DJ9����ד<L),M�j5��=&V j�N��ˍ���<��]��z�2^V@<�u/Ss�\�U�=�csݦ��<�����9~�g��5g���}){���OK�s^ϻ͚L_���Gm��.�-ف �mZ�܊��;��!���J�4
u��m�i�׷Va��b�u>�^���ܭfgl�@85H�J�m&�c�����焤lU��x_��X>tA���5w�˯xB<H����c�ڡ��rp`0�#ԛ������i�Qv����r�߮������_��R�u]�\�]���zy��sM�;r�g&���4=��,�0�R"��aH��~��bZR��Y�,��y��z��9��re�vi=������8e�yZ�b�ʐfΜ�R������D�����G��?z*��2�GP� ϼU!.���A=��;֘�k(�&3��rj���"���3�w�����xV_�7dRR8�jAS���TU�u��>׹2�в=�1}h�Nyu�Q(�zK�6��k�}k�xr�������kf�&��]
����Z�CiH��8���s�|f�k����;����[���E���)�u�-�.+Y���=#����ou��"��RD�mh�s~�p�ΗF�uו;���/8�A��Er�V���r�Ҹ�K���܌�a��B=u}L�v�o=�ߺq���ן�'{a��J�qti��Q�Wq��|�����LwGB]�wbj���������<�[��=uC�rY�d�V�إ�j*���wq����Ɉat�8T��vz�j3z��R��d�ڲ|/�������g�����{���w����z�^�/q:�u��Ͳ���l�u�Xn<s���	u�tWu��o	��WQ�+5=��s�:@:���{�{�.�D]�}�мn�K��Ms�\�DnEh-*<����C�e�QJ�w���ew����~�+A���$�|�;� M�ź���.o|��x�2� �.W�p�V����MdY�5�*�fJH�����̡��{���Z�̱�`�ա�>�e�*�RP���%��3�n�A�3w��j+�r�
�<�Ș�v]�wt1���3ju�p{�t,@�)"5�srη�vИf�DN�Č�7-�ǗȜ&��Z��J������ܺO	�Ԗ]�@�u(�j&�taa5�͕��T㲸�VJ��5V:u{Q�A�q��4�ַ�mFpI��Y�t�x��3�P�VG��[]��W�v��ZrDy˸ԫM��'t��v�2��kk+I��h�%n��F�Î�MV�N��)h:��huC݆_k"=v�".k��Ï��Ӄ��siHd�8��҈;\�e��}/-���k��=�D���q7Ү�t0��[ɼ�J�P�]\�&K}��QW%̮���5�f�3Lt�-�&#mr���^R��;%�plܛu�0R����7�Gm�W:	:�x�ݨ��^y���!Bxʍ���#ׂ�r�#}��k�`��t��I]�e��%����F���E�61��g���<�7�C����vv(� �K�b��#{b� ��䥻5C׊�z���Ss���1uV��G6�#+Vq�qPxE�S핌���EvV~���!SWǪ�evΗj������;'VG_l�����툦0<B<x����S���^�Oh�o1��]��Y�b�(�&	���w6�R|h�7�s�le��.5�be�}آ�����(��4�)f�OE�V�f�Kp������ǧ|���RY�{�k�Z(�̠�c�!ב8ar���gk�km>�VFK|�d$H;��*�3�n�i�*d8� 6�ͽ���'��䖵u|t�@4��Ԩp%pL�a)E���A�8�VW���<����e�M�����r2+��v+Xe��u�x��vI�4L���*��[j�K�� ��W�PO��8`|,y�ү��]���XQ4d��ٖ)L��of�ӆ���Sy�P�l��vL@��x��Y7is��(��e���"����_�0;f�k%��6q��DP���t��{Z#W�K�嫳�j���̷|�
���
�Eɇɻ��v�9�Z]���)v��/2���$��w�̏�����7�K������ʸ/��z��.ʎ0e9�3I���Ռ�([.��K�H���a����pg.)c�Vk�J0������v�;�����	���;W3/I|*�Hră�vwb���i��]��ai�{�Y�a�l[�6�7������- �"��|gvwwqH���~'�$��Ѡ�5��6ƪ&���\b*b��h*�"<��QT�DQT�S�Fƪ���SEQf��lQUQk1A5Q�A��EشhѢ'��1DD\��UELr5͙�͸Qynl�G,Wj�����������)�"��j�����-:g3Z������J��6<�O ��ɱ��"�*xF*)ѵ���9jh���*	�76�"�����
�5E4�EQAE^F���Aب��/��*u^lQ<�8�EE<�"���V�kTI2TArC����#X���.A��&J�(���"5�uF���[79�$�������"��s%�j������8���z��^y�Uh�1�W0STr�sb!��;�:d���m�� �������ccD�ATAsb����5:4m�6�3���i�ep�͵��ͯ8��W�BE���`I�G�P�K7�A�PfB�	!��_]�P���yY��Zu�"�O���9�T���/�Q��7�q����Y�N^�^���ȍ�Qo���c��q��}�ڰ�6�!�|Ǟ2��C=�K�W���k/a�p1G�Q2D�H�s��+�Ӝ��j�V	ꧪ�xm��l�)��.��� ��đ#�h��Q�/�>�
UmE�Y�nuv��^�t�N��`����>��������W�$`y6L�w@��U�p!�nv=�\EE<\3����plD�I��+���aAQ{#v�r���Ri6t��La��k�YsNv�"��1���8�*Ɉk�d�rד�n��[�np� qHե�OB��WSNd
� nM�!�f*m3��5}�8�ߑg%,�RzWJ��T*�m2�Oz�="n%����n�w��6�5k
�c}�@8� 
�����ad�$���������]d��z��U0�{ox���:��KĚ������ja�\mB	d`y� K��L���e<�6��aW3M#�zb��JU��$i��8#m�e�	�1���������G��=�P�ӕ>�7Vd�@Uj�w��(�W���/d����[~+�����M�hݞJ�W��gk^�<�$�������2��Y5�xS���>��Γ@YM�Ď�:��pb.��Ӯ����}�q�n=XDw>�):�l+�������*�k��r��]�����*�r�W^veoli;�t���#><�;��7���Q��T����a��j.�^hk������P<�ג&����2.r���|��r8���<������s�wP�K�[����ɝ��9���v�1ǨX����+V�v�X��#�V?s���f�w�v�{q��#q_�k�9LM�)���㮎/Ǉzʼ�s����D;?�R�G(x6j7�7F�Y���A*�h{�r��y[��u�s//^��0���;�[ ?$�+$�MI�$[0�ٛ���èq����VR��K��V6 0׍S�;;�^��j<R�v��ݿ��F򓸨��R$�S:Xe�ti9��n�ر#���8Z&�{�
>�N	|&���\s/K�"�A#L��s{�:T���F���{�e�ɭ�ޑ!�k2G����f���Ls^��s`�]�Ea�a��sR���V�A���VIZP��'B�ud�NsHg��@�"��$�ƒ8�9���P2Y��a���S]����Wj4Ofs&�'<��c'ː[D��q�*/��o�C�49��������1�Ľ��G�.}�z�Ϯ�m@��H�FR�&��e��cd����u*�����ŸMA*w�_.�ԍH~���U&i�?d�,���V��ؼ��M������e6����ILK����ï[g<T�wf�;;ܸ�"��m��B��["8lV���֊P�⫨�ceu�ͽb,�3@r���l ��'�Wsv ��y��oI�RA�����f���w{�����e��Vv:����x���<`�mp>��y�tKR|�>��no_u�CW��3=�Ң���ٻ���� ��`�[-�DFJM�7����:q�|F(���vN�Į�'Օ�{���y�^e��+)��B":����Xa�&ܬ�O�r�kw�K�T�X�	z�����v��g~�!ڳ _m��Z�G�i���\b2Eu�U��h���V|]�>��'h��m��BD���b�2nS'kg`(�Ӗ�;us��6>��׼������U��y���؎�[>�;e-��Os	�����Eċn�ᾆ����3+v��s+G0|�:���IX�ny���dױ���t��nW=���I- ������1l��	lN�1�mśκ��}��#yE�;�Q4�r�X:-́��yx��iE3�˚���=�5 �k(D��e��(u��TD��e)�պy�a|�B�'���b8���P���'�ʾ �Pu#��|�"�nL5N#s��s�A�^x���L�+�b:��h�J��g�h%&��"Q�R�2{w�b.��v*�ݙ�/SL� �yA��Z����7Tƶ��kj�����3O���je�"��	��X7-��d����'zƼOC�O��\�G�1w(��;�Rҥ"e��T��� F��v�Ӣ5t�-�:}i�!�D��2�˶�\}��#����S���Df����}�2y����#|j�<�_����r
����}f۩�S��ntO�Aj{�I�,ĭf��u�on^�%��o�'�C؄�MAl�Rea}o�����w��{�)��)�-xG�����\�@��6ڔ�/�!'p�Ͱ�/�)�j���%�7_x�8��L�.O�x��P�U]�t��t��r���h���vG5{����oW�l��NY�a�܊[��q>��TGL5��fY��IoG�X>�3`0�`�H���M*t��&�r���j.t�,���f�޾��KʺU���[t_��G6z~���VUF�v�q:��n"��Ɠ�������8h�a��>w1�.��ZV_>�l.�����6h���9����h
 �"A#���v
���nd��UL��N'k'aLoͣS"8T��J�e�������'�"|�M>\*1���E������n����M��{J}W]{����=���W�.��������#	�ר��S�3�(��$�Pr&:F\Z�Vg���\�W	�:���[L��2�=~���5��jG��E͉ѷ�ݸZ�0.��f�:V����^]���wE���(�::<�Y��m�v����)gwd]M
��{�ޚ����Ne4*��G����q8a���5�4 ��]37I3uU]���}��l���q.oe�!HP�>���F<ƜY�Br	�����[�4�osw�u��h�!���K��@Ҹ�qX��r�Eɛ��׈��g0��)	�zCr
@=��D)J�>U��e4�(i���9�`-��{����AjL)	��"��wJJ�ˉN���Z�i晫�����Vhɩ�S܆�V�ڞ
:�Eqh��X�*��(!MְT�9�xf�^�NU�ɶ aHpXVv�I�YM��u�wa�A�n��$����H��.O��
$�m����cp�|qdWYu��FZ'���3�_�ml�xăy�>'vM��Lq��a��s�^����	�؜jXغc����zw�%��54��d\��R��o�1�7�6��q���[�s�{���q%LknN��nj��}g\�r��G���DƎ��4��T��KK�����[�fn��
x�G1�Y�i���o��F�My�LV��iP�����9�G�slg=uVVu �����N�]cK����|�=Ld�3�r��dv�����vrhm�CX�E.��H��;��kXe�Zm���S�43����N7W���fqq������3'���e�7�B��_2�q��F�m�G��L��nH�U��Oi2O-5X��Zg��1����6�AF�3��s�O�n����,Ht�Т����UY��¦���0]�T6m��Z�C��3�4���=��yG��s4�y���}g�P*��[e-ys~�g���!H��;3���]�t�#:�)$W d�F�8����Xާ]4����ᶥ;c�����Ϋ���-%�V�&��;�fM�9��$e���/cu�&l�]T��T��=�L�����
�L�A#*���=	�|�q��9s�U$R�Ul�s�Щ�"�n7��ڑ�����G�����	���䤈��n1��T�ܮ�g/@�e�@��d�����F�8��%�9]�:��|ټ�ۏ9�4�ω��8Fc��>���b����{|s%ٴZ"��Y�o\	{c)UY�kJ.:+ND�/8 �sS�jq{����]���Z=~D��ު�vV5$;�⾐@~���=G!��V���j��K�N��u��N_���jx����-pD�#�"�4�;Y�Q��8,�k��Df�a����	�ܻo��1���V�s�z�R�S|�-�Al����݇w���g�5�wFHD=*z�|f@�[:��<�K�B�x.�,���^�d��:���稃o�!WOT�O�4k�NUJU���XP�;�򄨵���f^�g"�nH�G�|� �~���i1+�>��{�����,��D-�f(oV�v�(�����1��p=A���[=�f�==��2�p�ۚ<{+vs���r��:|v�ƇXc����vu]^��ʪ"����Le�g3;��A���;���Ko��d3�����º��g�5wf6����c78f(�]+��zV|�?-�S�]*^�'�@o�q�k�B/.ڇһ��9�-9��dv:���Q����o/�_�Ɋ��t̪}@g���Aꧪf���	�#�%n����jN�=>�n�x�5Zb��V�ɻ�}��Н���:i�sI�M��(L�ג^j=$ȫ�����y;իV���w����,N�b�r�z�Ȓ�����%�7����c�/v�)wI�cW���nwJ`gH���Ric���[�_+b���՘��Һ����O+e�v��\^(g��!\a߄zգ��@n!b��^���)�I&�ȼb�$���ߤ���g�J�*a!�*lL��N΍yG3[�V���R����R+�q�'�p9o��^��!�\��y�k
�2s�a�Dz��'[�*�t�H�m�.o1��z��p���G6���$z� �=�: �@I���pQ�[�6� <�l�R"K7��yݷ�2nw���נ�d;��z:��_G�z8�$�h�Ś�t̸m4_;�(�����
�K�����>���l�PhϬ���ʢ�b뷶r��[��VM�d��W^�0�a�f@#sُ��e=%#QZMU�S\�Wm��>��7��$ڼ��=Cz[�����g��byv��ƺ�6H���}��rr�r�X�4~��ѓ�=�x�bG���zf9��^V:S���T�=n�D���
�\�Z�&[�WPNF�ӻ&��dԭ�|/�w)��+#�F%���r��S��A8��goRU��q�]*{�f:b�.�雅7բ_f�SF��[�0%�Ρ̀�8���S}E,w(���k�\�Ѵ��߾x���Ә2=[�Lk�M
$fH��]#M���oc��R�春�� �C2<�ԨF^}ï-�v�	�"D�%�֫O)�EN^�����,��_$bg"��ڒ�ں�����+�L7��+6S7��{�{���/׼�l�}v�C�	5��Nzz�#s���
���9�;�N=ufr��]rq.ƛ�R.h�t�(�)P}lh��1>�V��1t�}M\x�]q1�� ���*�eP��۹�5mh���������ɬ�v��j���� w8_�܂<�<|�BS�|���WWP_���<e�˾n_7�����}��"+x�t��tyl��J��NK�yi��:r�w� \�,pEO������]o����|�<��1x��ٚEL^Y��=��6�aO�ppU�S��k�`������������>ow����{����������{��3J�u�l�Vk�/+V{�C���ݗv��#ց1��YOv��Q�:�60����%Z�m��3]v�P���Qq�vM�l�$�øLy����	��fl�ڼ!�2ww1��n�gL�]�:mG5��vb�ok����j�l�K�z+���1G�av�Xp�r�N�%O.���Ɋ��������|�;HK��g���#!Z5,����t&#���\vZ%��v�mnW.Zt;t�֪u���pçM�s%���]��-��q�tQ�s��ܕ� �{WYÊJ1Q>��)���{�c5�:kV���[G��$qoF�G��F!�R�ٵ��+���/�G�5�+�:΢�#����rl��L���nɷ}�n���k�[I6��)���Vr�l �*�8�Ƞ��;�R�Gm_Y�7!�;ƶ)e�!d�YP^֍2��r�����7��/4^Y]%	��
��JY������r��
�^e��>�:s	�ȯs��e�S͌��m��="�%��Dmѳ�����+�;����xy�<�z�1r�fw20�!��j��p�1���ڏ-��;�
C�=�`���
��Σ��eA)6��̬���Ӛ�eLobQ�^w�w&Y�f,��4�N3��Uүiq�cz`��[x�n$-��3�gl4 ��aE1u�(ٗS}�MܾNfe$�n;�]�XX\���,1%��˕I��z�;F��g��*"�e9�����<�fdڕ�$XÅ+�!bTr���Q棶ګŲd�J+���eҧ��t���ުx��yW&g�_���uq�Q���j��hV2�2}���rc2���MU[ϔ��Zr���4��,!�;s0H)�*�U�!�=�ߕy��Gς�V,���9b��҂<՘*��q�a����j��X�F�4E$+5�,��j��]�	�MW�(ӻ�Gis�8n 2���Q*��0�6]g2�+H�i8�=�cz���F��/�@M#�ү�~�oMFQ�P ;nuɒ��wu.�����ht�& ��]�gkF3��2ֈ����
s�]-eu@�3],R��ܹN���:W|� �X�0�^^0!�lC1-ob�t�M{HM<Q4�����ie�nfw�r�����oy��(���T�NQ)bi�	Ӭ�|�F���*�ovlF�S�KOJ������[�
�p٦�����K��9�����n�^�F���0����pP<��[��� qJ&�A`��[�S��wVu�X�v���ϑ�\��I�CAT\.�sn�;+���d�z㫨��Пf&�K��.���ۍ�Ƶ�X6�����&�ޅ(�mZ<7X�!�L[��Ȧ�tr�N�
��wi>��=�\R�W�;y�p�CS�����.Q�0���lmݜ��f��gR�r�w�'��X�m��n)����p��$w&��,���[yS�A��φ�����afLםFgt���mb��X�QD�.�L��4�
H�@�`A3Dɷ��oZ�s�co����i���76�"���9:	��s�k�nlUQE;h*j�*h�$���ji�+Z���f+�qUcj�5Cmm�-ESUU'5��s��\-E�آ�2�-��(�y���4�h�0a�����"������U:�Y���3�T>\��*��3T�A1UM��f��6ų�b"���Z
���
(��`�U�&b��G�p���j��)�M$LQEm���Y�5����cEI$SAL���5O6�����q�EPDEDl�h�#IPLDN�*��f��֢�B$Ѡ��m͚/1��l�Q>g,�Py;Z6��/Y�T��Ah�i��bj(��	�("+��gZE���f��뙢��j��Z�њi(�1:����[ornX��������@�TAzƈ堍Vv�'CĒ)��ǣ�p%���Lu$�G�r`u�b�;N���+��.a'�2X���"R߭).LU2��ؖ9�H;�de��7M�莐-�]J�V���oUf����ۣ��H\�����¹��5�Z���Mwٕ�Ô���/��W��[�U���D�wd��~�6>̉�z���x�����߆��Ǽ�g=\��KR&g�?�d\���>}q�D9�]lx�v���,DI�uH��;���ஒ���x��1�X����9f���76w����5Be��-�^�^���"����79Ē���.�stsM�T�%�/gh3�w:�Ӂ��̨�J�����������*Q���b�ɉW���9.*�����,�����f?$�t�Q��d?G>a:t�^W_�����V��E�VR�6)̌�{[ii?AD%�m�8.��;�.r�����!5��4�Ɵfڟ]2����w�e��;j���ʫޭ��ց��]_-1�x��J
U�H'�Q����zS?4f䘘s��Փ�r9�)�ͳ���'u�E�և��ĺY�^�:nB�x���˹N5�%�`U������Mgh��,�Z��3xj6VG$��;��)��l�"���i� %`smrK����qo���R������h��D��sv )�����&���(?�<#N����m@�&QHP'"	���φ��_>���ڹ1�W��8��s0h#0BY��e��R<*���*��v���u�v�iTk�%U�ꎺu iq ���B��[M��v���֛���P����;�~bx�kzL��]@���X�B�&�����-����'Z�o=�2u��ց���&�+��|�;eH���Д�����]=�Oxr�0�κ-�AS�����6�F�=(%ܻv
��T���E����Ή��f�O0�3������2xdn{Q5���i@�%Ya�u�O���f�
"��ߘ�P�� ��ٞ�4�9+�>�ˋ��Ǟz.v�p�ɭYѨn��A��������[�^���Wx���]WD��ޛ���[��n/'l�Pc�9��e]~�"���%����tI��6�b���6+D)DZ�07��{sK�k��Q,޲��}:��!�O0�d:�oU��T��T��Qzy�.���X�:lY��ٽf�Kz=��g}�6������+����Vpv@l���y�������I��O<Y������k�L���/'��wQ��+�u���:Z1�� �jo"��nc�cd��F_j�ݍ՛�F�$��9�{k��қw��$m��ʮD��6� �������WU�����_��%.Z�:��bnٟ�^��i��Ns�.��_P�z�3g�ёR%�/�/#����ȉv9�t�ưa���'u���]H��W �p�-Z42W"�VEA�����i�����@�z�A�<�����M:�� �("����5Vk���~W���&|�$m�z��E���d�����(���cs�n�d��Ù]�׳��m�cv#�(lD�l廳m�c��!�F&t�6w��P"��>�G��*�|Z<:�и�}p���	ʞ���)��sV���/�q�;	}	d����v_%U㋢|n�w���U�\>v��[2�F�z�W7�-cv�1X�;z�V'��]�8�V.����+���=K=��V��.�dN�ԥ�$��ի'cܔn��xT.����V�%a��f,ܶ�Eqͧ���n���d��@RR����x�:��n��2�9Ă~/��h�\_!�Fl�������Y{��u�oj�ǥ[��C������K��v�*z���:��� �Q;ףD��5�o'���a=Ҕ����|罣�g��g�eK]�ն�+t������6Q!?M�{��#��J�L�˱��@��վ=��]�j��|m�s�I&H�H�b=�+��nr�;�|w��Z��*I����F�p��{����3�2m~�/wku�sM	6��E�A<�,Ǟ��ں�u�����u��og�`�R�k�/S��ӓ��s��S
�g�7c�7
��R��٭9�C�-37�{�"ﶉ�KlaAJ�3�'p�E�)��26Y��8���`K�Uv�zۮ�;,�3�pTJ�Ɏ��$U�*����ϼ�8��-��������b_b��%���Fp�̩ԥ9�/�I��0zۧp��$.1j�Gg�X�ն�ܸn�fe�3/�K��uf�E:���e6C��,�f�H�L��[{
;Gc�M��a��&�ܩ��Ѻ8E55���{ݬ�Sov�wE�!{�.��*=��I�P��⮯c����տ��˕?h�j�&�t����WJ��*�ʾM��dy�m�����U2�@8� +��&
�u�[�}�) ][&K�=�}�ql�ů�?;z����2����m;�T��ນp�-��v�NV����\h��t��vvϻ���ɺ<���j �5MM�����߆��[Ά	��'z�ٰt��Q'˓�f��a]�l�]O�[��>;V���Zd��"=5����KQٲ���wg��H4���?��r�y��Xۧ7Q�7ݔ5/����&_��Kh$MMO�9I�E>���Ec�x�ݵْ�_ċ�z�Sے7:�9�.�o�+��v�1л�v��N�+�"s	�{���� �B��dF2���m�v2=E�kTE���zh'x=���Tة�t��,Ϻ�8�gwFa�Y��}[�@��nR�^W!�')|�4�k��-�Ò�L]�mKö&�͛������P��j�	Ѻ�\<sN?]%vm��:d��Um_��rx�Ajn�������x9,l���}�FVL�p;��i�I���udǔ�+����X�|3�lA�u+q��'0�o7�����{�|t�#���S��g;�]�����t�B);�kf�᭭��_�]�׫�;��T��E�����~����g�`��Ih�V}�����������➯nFH�(MtyD�4KsmM�.��۸��jܑm�lȝ��E�c�g�0�f���\B�'���"�،�u���fyy������Dw�H��OY�г�҈��E�l��
&��PC�Lc�O~���wܱ/n�����y�����EN�w���,� Z�e��Y��k'`7�$����f�s�C�u^[Q�N��\@"�:B28+��a�w��uw5�k"��X�Ikr�M�d˨�[1��� ��ͭW�wl����oG�	���Ѷ��er�|��S���wf*�C�m���;���"��Q���#�{'�_)�ֵ��x��|�8 T�\{d��(ݨ����\��-v�?OH�ɒƭ&�������/��}��wl�̈́	*��n���Um&)���D��'Uc�$K��z9��ǲ���7_N�8�8M���5�`W&V���wr�����dP��u��[}u)�΅��zԤ�����6��?���ߟ�>�x�Ƭ&�y���\&�{�"]��3�0���ӑ��P�L=�v�7�8HȎ��2����1,7ug*��ea�9[}�9ڥ��:���|�C�"��?o�� ��~P��乩�/8k�i�8nO��gݗ� ��`�0i�=D*Wb�I�۸S���`�"��9b7�������L�Ic�d���0�Agy�瘄��5�q�ͮ��Ad��ͳ|�ۥ��ȉ��ADF�g�[*�U��^�aܡ���әs!D-�T��Ov���dЉ��������UX�Y��w�֑��Y���[�2��A(z���͞|y��d�4㝉r�55�w������m��S���H=p*%̌��`|���#�s����mfh���5]�{�����_j�.(욃ʏ]�駏Mw���("ϯ��Y��N
n�܍X�q�[���ɕ�vys�u�%�f���{|=s%�sD������)��b	�٧���
�,M�wJ��H\�� ��s��s!�1��=���ū���>2_,��ե�b(�M�ꑢ
�{�
���;H�\��5K$�&b��|	5�8'x}�;���F��5䊐`���S�n�u�ܢ;z�T6a����]�0�$)�p��i�	�v
7�ܑV�*R&Y���Ev�b�
�8|ђ��Tt�?�+B���#v�Z`/�G��%W���6ڑW���M���U���9�O!�?�j���r_��,H�3�/�F;��9�b[���n�������R��㱧�a���z�d��-Mgso3��}��{��7h���Ǭ�K7��*ݓ{,2�O����<��ec�WR)�nz�qsTv_B���I��d�ڲ��aWG��=M�������T���u=�on��.$�6]�/��aH�~��z2{�gݧ�&�ߓ�O��o�zrz��c��<+U�N`��\k��	�	����i-ز�X�gp��)[��a�R;�xV�ѷ�o�ï-�ݽ����c��6V�,��
���ٽ�9�k�%5�S^ג��^��He��JZD9��m'4��!�a���i;����Q	������y빵"�6�KGF�0s��5Khڣ���a5�u8��u����nY�<M�ު��.��j(H���+�g@_곽�dJ���j�	�hHA<
$�c������U�h�c�{��)��|�A��`=%>�z����+�l"^��e���
)EY���{S�կ���s�#b��H��
��p��l��j~��S�b/��\@݋�q���te.Ɵ^Z����,�S��z�Vn�=ɝ���� v���z]��GtFP�h�5�B��WV�fp=jSK��W�[������Sm�,XE���$z�*
R�jk!���a��r�}�Rj���@Vy�BQ��Eo�Iw��/iꝉp������ҳ�䣽��Ͼ���ׅc�|�4=���J.��'�Wt���Fl�Gj^�D��	�����r��a����e_�%GI��&�]��ۑnc��]�B�>}o�!_��Ӝ������Q�Z$q����~��9�
8�����8�M.�q��]�'v|��L7�~Q#nv���b���,-�o��aۮ�t~�S�S���l�'��xZ�=h8h����5r�W,�fv�n��4�"�*�{Wx���ɚs����$���Zg/�,nŽ4�����Y��ڟK[;�(t�$�9v���ͩ�o�[�I�������M�Z'^���*��VT�Oa������)�������G��	R��d^�;[�UuN\��i"��=�^l	�b;ے7:�9[<�o�Fc��e�nEϢ�Y���1}���Ʀ�؄a���,�n}{�z�9��n�nY����n�-�.�_��:�>�!�@`F<��n%V��;2hF���;�v:s2�q7�$H�	4��O�2��sYΩ�j�|H	7��}$_^r��.�Q��WDD��&��9����r[*�j��)]���ֳ���H��%���,���+�$�:��ͥ!��a����g�w�ÝHsY����5N�����\B�J
|���{��a����͏sx��ۺ��/s$\�F�y��QB:��T�p�[P*�DNoS#{y�����{H����u!Բ�G'��� rp����n#���z�^^>^�p�{���w����y�������"��7�S�3��P���3�t���k�µ�6�w���ː��G�K�b���'������y���6�7#W/�+B���遵i��l���
��wK�쭆eΦ�q���.���z�����L̼��[[mNM[[�g!��[��A����5#y!Y���&^s�e��[���7Ri��+���[M��q�THM�T�v�;6u�]6,;��^DH<;7���9�0��:L�nN��Y١�-��L�*�w�C���� [��kl�Xi-�ۛ)�\Dԟ:��Y� �!s��"�&��Uٳ-P��lYSl����@��k�ԧP�E�v�ܽ��$�YP�A1��Y�*���[9�lCU/w^��`I.�[����&�.d�{��H{4{�y���꺉F$�5�	�ے�'�[�ю�uA��{]
z[���2L]MO��;r���1������-�Vr׍�g]��`&s3\�r؝@;5��u��8;�V�5�8F�	��m:!o%�w,���(���v�� ҡs���`��hs�zEd֗��sl��:����w��u�h1ɼm�$���
����u�����i�M�w���P�Avѡ�ojVf����3�2��&�4N���ilC%�U��~��&�;H����v��@3p���|�"�a�(�qk����=���ȕ� ^d V��n�ҧ���C;T{F_v-Yw�Gu7*��NL4#ͺ"����r���貙�}���Y�p~�ھ�Юu�!����I��������ޑ(��Pv���s1���=q#]�X�XT�c$^�,|����V�2��Z뭝,7�.ɒpoon��]�H�-�啉�Њ�����GU�q=f��z�5J����3��!ϸ��ʓ��`S����.��xCڲ��!���F�$ �{a���4�Yk�����ݾ[��;��l�l3j43xf�͉�X�D5G܈����$J�oj�;!��e�;���O9#M�w�=R��k�
�iۜ�_�;�Pf�̬#���[TM�v��a�\6��˛b�0w?f#�.��NǗ��+'�/A7��xV�f���{�<(�Ӟ�Ɋt��͆;��K?k�`Ru!-�[�D�K����#�7VGl�뢊�w�{Y���ۻ����ɳ^�Q�L�t�L[�H9t��3p�,��mt7%*i��d���(��<�]�;sD�چ�3j�)����4���E����Ǒ���dAi̆��5^��t���ٳ{�K>8巘�s�V�+9x{m7���K3�z&�J���3�b��p��Y�4�w�	d��tU͈j=,�jà��y|��WZ�5Z��3���"Բŀy��7\u�1p��@�$��������pCS/r���Ob�s���+��1�u	������2�!D�d%�|O�@� A U�IU��jb�4gN*��(�h&��V'Z����1�o1�`��:	��ƹ�;SEb��� ��\�>���ƨ���� ���*��i�EQ��LPTD�Ss�"���V���h*�ݨ��Q�2ETQT��כ��l���Xt��F�����QF��3�$�y�D2W �TѦ��q��5Q�h����$�QS�;��.F�G��y��Q4DDm�ƈ�kN�"(�*�+k9k��C�j
����j�1AADl�kQQ�M�V��*�M��gS)Q��(�����TDQN�5$E0SDQt�sX�U4T��\�1͈���y1QA����+�Zj�+�UV�n\��$(�hѯ2j��"��y���D�L��^\#A������SMQf�W&�(�4SO�Y�K���_��dWnT�.s���F��
[.������s��}~Hoy��3�ƕ�Y]Ih�#3�p�j�&Ӯ��ݽm��l������='��+�J�?T�u��^kgB��ҟ@��:ZfNu�"���k� �.4d�<��:1�m�5�q������;����\4$�Ȏ��u���J� �\�2�Yϒ;e]fR"X7D�v��(퓭7,��41�T����ʾ�)�A�Fx �w4���+#On,�ڋ돴n���Ru�-���P�<d��]&�\�~8�?�tx�e�>۶��O9����V�}]KjFw�u�q�b7��q��(1ݕ�o֏�7��K�aU�a�q�Z�ƛz���FnH����6�����>�]���j�y��k2�Zp�i��\E��ʢGi/�(��`�}�\*��]��UC�N�����CHg����ܯy�,�H����4�%�k�:���y����١�s��緖 �cv<�y�j��7ydA�F����͞^GS��S�����k�of�����P���������l���0�ۭ�TI�܍�K�a IWZ<p"-f1��6��vZ3���z�g2r����y�!л�oq��oH�r)�ml�f,#:��w��t��h:�OK<�(��w9Bt�d�ۼnwQ�OQ��L�GD(�v�D��fb�Go��:0^��M�0�y����z��0���s`�����s��,����	��8��*�~�;����mo6�`Pϝ_���@�#�Ri#� ��ÚY�
�9l��4k;�{g�n]_��v��S�H,�J3G��U@a�ک��j@纰wm�K�:Uٝ�y����i�����kI]H�	���n[���\{e�v�L�|^�(l0�aE��t`��̇ G$V7JH������̓��̾�D�Wh�@���6̪�-��$��[�W� �m�ܑ1q�vwq1j��u=����%�d�����_%5Z�|3"U�����y{5��}��׸�)烂ߒ��б��d��U_aT �M���q}�|NfUoK;���vM�l�����}�F_����:�-�E��V�9�n��r?�3�S3/�͍���f��bg]��&������AL��J��3��7���X����{F�SE�
����
E13�%��7��7-���g9|s5[ر��K��ȷ���q�����x/IR�Y8�S�$�=�=ܭv2�L���-ef�ޔ���{��J����YD�RS�df�������w��ޮ�h��3&&�T����nr���M�Xz2}�=�	V��g4�㬭���O/�T����+ݭ}q�I������Ɓ2D�;:�yy�ެ[�o�5ƬVH�n�؃��f�������9��9��7�d��v`;˄��hptT����؂�����f��I���)���5�5��3'�����D���ɺ"s�����b�{ ����Lŭ�O��Z��H��vy�|D�슸�J[�|��]m������sA���V1�e-�����Ւ(��n<���r���!^w$�ZR�9Uy�A�qK��I��2�v�d0�Mˢ5a��HnAH=��%�ϙ�ekUI��v{wS���kp^d���\�;��3��I���b,V�z�]�$C<u��o�/Lٔ��R,[�E���i��6�X�ׅ�v�x�w���|�i�R��iY�z�εW��o0śps�{��Z���T��@̛k��t�
�ĪB��ٓ^&��,�`�Ik-oݽ�-�����!մ��:e���F��I���/��gY��[@Ol�����1q�˦���[sXٝ���i�;.|�ܝ�� ��T�0�B�T�^�,����&�Z�o9f�Y�T�b��7k��>�z��}1�H'O����\�	%���ٽ��Cd�<���[4�����x�bB��wM��`��#����:ي�����r�<.x�|�C���ꮙZ����<S{R&g�k�a�����X��:ק�\
��;�C�GcY�j����Z�U���_�N�Bf�'��&���#����ͣ�A�ٱ�'��-�͈Ρ�=���VΨ�}��#L��ϸ;E�Hj��C�<0"ά�a6Ldd��͖���ñIftNJ��P,���x�c�ϴ�W��\��^����y���d����_Swe���V���V����N�UG���oiH�9����/ǆ�*)��G�R%�L+���6�o΅�]g�ɽ�E��/rq���+.�SS_m9Rw(��&�\�:KW
�ha½��"�����}puV��vvb�ݨ�r_k�&�ܵ$��]u�ю`�DhJ�An�fU���P��Պ�;ʃ���*�P�o��܌�HP�|�K���GZMR����@#7?v�{�}^n�8�S���W~�-_r����w0���(�j��"����=��U��ˉub�
�P��</V�u�ݡ��G�/]�a���������R����N�U�)ȩ��1��Uo��Yx������d1$�s�	T�Jy����庑��!f,��_�WqV�M�= �?-�[{͝Ғ��k���Q8d�}7|�ea��0�ʻ��v�xPMÍ�xnۛ�Lm���4������x6C��d̿u�T[#]�d��o\o�u���_)���=i�_��+����uf^������jcQm|3|u���l�~2t97Y�c#T��Ṇ�N�^`�� u��J<P�T���ސ����zs*�Tؕp�X5Q_���ٵ�/7=�a�&��m'쳏i3��
�s2�^�_u�Zˤ�Z�gw�����M.������fϮ�hJYk��'�8i���W�6�y��A��qn�x����!:���K0���l��u-r�hm�MB���ѷ1�z8u�f������ �V�0e��� ���{��!e]�O�y/Y�t�i�۫�_�JX��=�/��Ď��1�v���1��;m����<�ݘ1\��-���	@��[�w�v���7F��:$�9��{�[��_����3�Q"�9-�H�c��DI�D���沸�]Ϩ��=���sZ�R�5�n�CXP��G@�������2;_h.�V<nޙ쫩���F�G�+,��n�g�z	@����3���k���]�w�D�|Dx�6��H�O�]W�`���
�?l����	V���������^�=��Ot� ��xQ�4 �=�=4�L^�qma�=�դ�a��������p���py�.��R�j�)<�z����-�g�#�ک�x%{Y��q�Hɂm�+{u� �nH�a�%g��`+�[����:��]_�k�7�^;C��Ԝu�k^Q��:�Z�g	U˝7�q)�g]�~�T�#o�{=����{��,�d��뇥�h2��li�7��0��i�q7HR�܅���b�wAJy��2��	�@X�HA!�d���6�U�R�f �� :\�m�Wź��xV��ǔ�w���zz�"t�����0�^d��.���w�,��\�~WȜ��J�_��:���+��u�8�l��6��d�5Em�H�W�Ϋ/�oW�hȳ�~��)^�J
�M�t�e�#7Chx�S�Ca�R[cw�_vP���МG�f�L��]�	�Ut,9��Sp�}���ܧ����ve��!5X-Ƕ7>}�
D�~x��1
��O�	�`���Ǟ=�;�7]�A~�`�2�|An|�>�l�[�g�i�2h{h-ζ�sQa�2}��+uS��C8@��f£Q��<����0�4�B�DMW�#�j陆뿜���h�TG��և�9� a7礥�j�/x�=$�>�j@� �"/�o*"}��M�yz�g9�<�R��ޓ�VX]��us�~����/�������dv��aAt�\^4--�%�9u� �<9��u��5c�Ap���f7s�����p[$Q#��lm>�5�I�M!��`7uЎ
N�w��ݦ�`�ou��"��ƫ6�7�ׂ�>;v(�K�ڕ��9y;�O24�KF(��ܷ���
�]	v5�,��9T��p����Oo�xs���8O�bU���=�B��IW�)U�S헶�����m�vT�Tөl��Y7.H���]�7/'�s��T���6�^�������9�A�}��4� u�Fg�%����/c��D-�H��k�̎���I��28��d����!O�P�����of���j�{�^F�3y����E��>̬�9 �L1��W�ť��nS#gxok,�E�EJ�=VSQZ��GU���R��>W0u��m�C�I���T��І�z�� Wu{9mP%�+΂wt]:���lh�ӈ�u^o;?\01��2������5lB/�f�%�&��s�G������j�%�7�9����+��@�@�q����;�J�����;�w��"��_�������
u�E���[ ʹ��i���1�+���PY�DP�B���k��4����|��Q�����w=F�3���7��t������!�m+�h�^K�%�]�]��W Y}�^��qV@pJ۬�U���BE��M^omlm�l��N�c�Ǭ@ �{4��J������>̚��n������u?f_|��,;�n��pܞ���ky���3�ú�0""�a���h����nl��{tn����H:y�v
3�~��bN�z��7l����޲F�W�]7��ݮ*���W���ȴz��3(��Ӥ�������d�^�g��� �UQ==[���+����*��ət���[ur]}{"��>��0.�ѐC�e؉Õ>\B��%�採*K���U5]�7��TfH4�G�G[��H�$�me��;'s�{n�7O��*�R�$e(1�j�U��U��1��^6[��v	��i�;ֵ,�Y�ڑ��os����P[P6�<���ZP��	��K;�{�r�A��2�u�6�)_���d�]@�({}�q���"��Uv�?�G�2K��b��A\s����MW�bx�ٛ!N�������>Òݛ��9큅2�`���F1[�M
�ajP��c%�{�v`�eip�C�X&ə���.��=E�r�ƎMdinvՖI)�3NpS�1nL{�f����1�C�Z`�m�SZ���(�ҙk5�@��2�u����]O�Q�K�;`�L<��f��;;W�gm�T_�j�,g�f��-���ת6U�d�9f��hf�`��3:��Go���&'�a���ȳǌ�{�����T
�������>#z}0
-:���%���GN��쾉Ý�X�ɱZ'���v>���f��S��{���պ���W�C�3ݝ�hl�Tsv���Ox�V�;-����v�n�z'ᛗ�Q�J�%
 VV�o���v=}{>�+1�1���9;>�!�]��{�����2��/��O�jѽ� ^Y'���a"FL��c��{�\����mk+WE��,��v�������,q�?E�Gs;^��07�v�<kD���ܜ4�!�}`<;�o^������%��#��
���"/����i"(�����������szA�2�ȳ�0�0,��"̣+0,ʳ"̫2�ȳ"̣0,0,���*̣0���(� L�2��ʳ�2,³"�2���"�0,³
�2�2�ȳ̫2,��"̫0,����3 ̣2,���(� C"�+0,ȳ�0,ʳ �
̋0,�ȳ*�+2,ȳ
�̋0,ʳ�+0���� O�^��Q��r,�3̋2���̋2�ȳ�0,���̫2�³�>�.`Y�	�fU�`Y�f�beY�	�fE�`Y�fE�Ve�dY�f�`L9�fG9�fA�Ffd�f�F`�f�d�fB`�f�d�fA�Fd�fP�FdY�fA�a�fA�Fe�	�fTd	�aQ	�& @�d@	�@& �` 	�%U|���@eUf  � e 	�U�PdUf �UY�` 	�U�UY� &  �UY� &UVeUf �y<V` 	�U�UY�U� eA�dY�gA�f�`Y�fQ�S��`e�vy<E�`Y�f�`Y�f�t�Y�f�`Y�	�fQ�`�oq�=|A�w��@(Ҡ*)2 �Q����o������>>��������ۇ������Ҡ~�O��i�[��� � {���� ���G� *���Y U���>��O�_�O�o��� *����!�~g���$�������C��������دɐEY@QITdT�( B$A`	�U��U�$@@� %V aU`F  �!Ud UX	  �  �UX�P�H  G� ���w�� 
"� �BB@}�������������������_�� ���`�~����g��ρ?����?��|����� ��~Hb~�y�'�ߑ@X U�h~����PUw�?1��N ~ ����&����|�x�o����xz���=�z� �~(����H ����=����pg�~!��~���������8D U������� ����g�!�R~k���N����C��.���r|�����W�{��>>�2� �~ ���z������A^��>�0}�~ *�������߇����2��b��L��Զ�	1� � ���fO� Ċ���U"�Z&Z6�Pa%�2���4�j��ŕ[kX�5k6�mF�m[,i)
��KAC(���M�cUm�P��YjıVfY�%������2�EնZڭ�ҫ[l4��3F�bBQ���i*�2��&4Ue��F���J��ΦivuWj[4f����Lh�ub�+!6�K5Vl����c���ȴ[�ڳZcRڶ�֑	em�kScd�J�����ј�2ڪ�UB֨�Jf(�ҭ���6LZ�Z�Bf�LZ���m��bٰU7����D�)��  7�}T��K��j�N��y�/=^��N��t���Wc������n�ڍ���ڶ����UWjڭ�v���
�5;�in��ڠ�j�={�/[ݲ���l&mm��SJ�Jڨ�-�j�  ���P�B�
>�����(}
(ho����h @;���
(�����Σm�k�צ�������^��$J�������z���{<ӻ�mM�isO���O][mo^��J9�����ik[h�1S[k5-6����O�  g���UO����y��og��^�W<����z���]X=�zWJ��շ{z�v��kCO^��W�z�����mۼ�{����m�{wt{m�{ہUS�=�{z�㙊��{�����]z��m�u��[[m�����nʚ٪��  ��>��Nu�y{��Mvo6���=�M{{�Z��9Y������x��٫�j���ݩj��^��ڷ^��{m{t�^˼=5��z���J�gE�2�km�3kV��l�Z�� ��C�}����R��ޭ��]�������ק
H���^�ƽZ��o+=U��ݻ����^�Pov��zW���ZoZ7�-k�0�5j�lV)��  ۼ�W_[���V�{�[���U.z���Ƕ�끪��;����������Ҝ:�ݽ�z���κ����w���ooy{fjԭhڶZ!V�j�Yb>   t+��b�9N馍��:���F�����]k���mGE:���z[uC�ǽy���@廯x� P��ہ�z�����A�P��f�1ZZ�kb�a�mZ��  w|  v�;hC݁�UY� zPs�p ���=�j�� tҫ�+ �C����Vt ��G/{��%���L��@顼{oxPR��ճu�i��Rj�bKg��/�  �>�@:�v��P��a� ����]�
���@(
w��A���� =
����=hR��y� E�[�
( {�m�fVh��֔ͭ2�+E�   ��h
��n�P������(@o<��z� kޞ��M ������B��y=�: n��(z����Р��A�)_ "��1JT� S�d�)JQ�  �~&BR�   O�JT�  �@5IR��  	4�&�UM�  ��?�����W��*���9���?�����yu�j�2GeFZ�Ҳ2d��B���������{u��?�H�}$$$����I BI�В@����ID���BC��_�*�~���>aJI7O^i�da�Հ���#@H�.*5�V�2�X+U^�G($�Fi����$��ٽ�8����X�f<N�iK�����X��M��y��ʕ2%r�w��>,D	Us&��XYq7;wJ������mK�A�r�]0t��`�L�emP�����\zM�彶�6�l91B�{�/m�A�餍��ᢦAp�l�HL�k9/�r$��v]�ܾ�<���䩲<��Ū�Z�A�9b�sBi-�Y��T�J)�m��1՘EfA�J��I�ݷ`�[�nE�4s^(�����*�1]F���)!LfӥM����C��[�ɕ�́q7B}6�M�;2F�oQ�O[U{1AZ"���� �{��I�{�AB��5[X���۲f�y�VƩ,Z����1��me�M��Qmv.�fa�V���nM.��i3	�"y���aB�:�?e�Ʋ*#	%`
���2�[Ņg2)�f�[)�n�%�1[-Z{��tꫢ��Tm���(���Ԟ�ؕ�.���'TE�Ƃ�C�*�mkrV��rFoK�.k̸�Xr:V�*�g�P����s1Q2
���u��b�/Ż4$�{��JKr�"��l�J�ⶨ��ˌ,B)�9A��$i�#�re0�o"��dEy�^]c�YwzT�O�4�=��L:v�XX���V�S[c\���!%�.�c�Tգ[3t�X�VfS��t�Sh^� �ͣ�ȷz6�h�{
�b�x\0�+��K$n 8uK�g̛�� �����-��l�&��hr�ԥB�r�Y, r�L������L=Xk\��0i�D�F�K�:��U�3�S5����K
�tDy(�wN�*,�C5C��͓�04X-���\YXK�o4,z/C`P�bSu���q�`۶UJ�|I�m`��u�Y"�EiQ�Jy����#L�t�nV[�DXZM1K!�sU#nI-�l�eԫ�J�mc�d��X��J#���>` $
8��-P����]_f�)p4]�H�M����;6�r�'�Ӣ��X�+�l�7d���A��,;Qf%+`�x%�a�u���t�� �P34}2�H�yI�`&�BӒs3,<�N�̒Y���(�4J�����Y��H�U���&i�p�:kh��m+�A=4��(a!PA��jސ�f*��Pf!.i�˚%B�Z�$��m�Ȥŷ�Va��M��ֵ0�6���Q�]��rR���EG�>��QFi0��QD��v��MH��W[ �m��h��^ƒƬm��A6��E������	�����T���ac�`���q*s��W�ؓT�!VQ�$h�L�����rn�����O�L'*bS	�ou.��J�MxFL.6�T��l�R�F������Zնe�d;l�QDj 0�{/6�id۔-�y���ȧ�P��-I��V�J�m71�	l�F�W��7oj8e?�FV<o z�mIl2��"ك.l��
%-�u�b�"�
�)[5t���*�l�Ш�̲Œ�
�A� ��q�b��:И����F�������`p��n�p:xéYch6&f�X���cL�N|DHH�Rl��-i(��L��N�<���CXk8�l���q���Wl��p��d���Qh���)�sr�Lף�T��aG{č#[Q9�haSL�f��mF��R��2[�$�@��	((E�0��)L|n|0]��E�٩h�&^咤@�he��	ͭ*6�&�d
���: ���rfSp���{�ڃ�YV�7L=�A@��I���uH�c���;�ۅ^�C)�j2�����\ȳ�)IAnAAR�dH��������)��X*m����F8�V3NGwe��)T�t)�Q�96艠k��X�2�Ȭ�� SYIC���Ӽ��.�n��ب1�7146�^Ku-O��Pr���R���9�X�Cd5��4ð���q,w k��aT�Y�F�d^\�L,�M��Z�uX�j�f�3/ j���ڬ9���������el���{l���!�1�Du$���" n:�4���Ն�M ��$�kl0rj/V����~(P8q)��Kr@j�4E��B�+��)�maQ�p��Md�Zʻt��*P�쬕��M��-Kr�(8]���b\�bc"M4iv���=����`e2qϘ̭�m�`�5"U�N�C2:#p�B���@]���v�v�b#@��=nc2��J��!�����r�d�&��us���c&��N�e)�} �������X�:�AmI�l��C@�w��D�P3FaӔ'֙�!�ϰVi$bz`P�f��B��7�m�U�M3J��f!W{�*Tf6�Meh���к�op��K�ik1���u�V��$�[��Rde�ГEv��[���˴q�
�%mh��Kv��9�"��|��B�oF�(�����HI����\��/� Ҭ�j��ԩ 5�sܤ$Չ�(IQen*�ߖ�U��QѦ`�n�-e�2a�ר����;A�	5���8�.�^T;0�ַTE oVd��
���JLƮ�s@O"�́w�a���)�m<Y����*��h���O6,��$F�#�W��4��Q�n<�K&���$g=}�,�,ç���}�l���>�,�u֘�t�b�XA&mj�`16�P�b۷`�Fh�@U��n��@Uu�ފXM�ī%�ȇr���(2k~3S�J�8aFj2T�Y�u����ujq;���B�R��A�RDW8%.&�i޼Ϯh�5�Y4io+u�X�5dv����fla���f�qP��7"wj͵Q���#ǏE-}�aEjr=�yǻ%<�U�'��fÂ�7R`�cܺ��e�ct̰�Vڀb��;*Y��FPʖk�5��H�M�>���@�D1��LhsF�L,Bm�h���ٚvD�RY�3f\���z�5�vA�I��Յm�x� �*2QU���3��K�&D��	�Ͱ,w���\��kJ֩�q5�Yu��p�ZD$Gr^7��� YkJ�cC_�ڽ�,�v�]�4Qx+d�[(Ku���1 �N;�h#�a�2�������#N��
$�oXʚ��3C�VF�E�:5K:i�D2,���<eO�Ɗ�d��&�x��
�n��cWW����R�Je�K�є�^������4��n�i&ތ��^O�a��˓�v�I'W���r��C!b��eJV�)&)�`��x��A�ɐ�Kn^c	�[�#@I�h�_��L�d9Jd��a��l!��&��2��ݧ��gE�
����v�ɰ�خ�䴱�(�[�u��yf�U%������mG�nl9-mǦ(�6%�m+�V����7�ǚ��]F]����.��5��T�$h�ƞKA���������.�	�B�MTs�d��qP�O�z�aDm櫼��������W@�1Sh���Fk���n���_�ԛ�u����b h�W�,6:�^4��v�K,T�0fQ�WH�g�H;�>ȮfC��l��A��Mom;��@�e;��(�؃��Q�wYF9iZ����̡���nP��tʔ�oK����/���i��OE6%Ye�K4IV�L�	E-�s5�i�����T�m1%栙)��J�l;-�(^����]�[{R�=��'��5�z1�Q��ŐL�5��U�V�E���cP�Nٖa�ԀUa/i���h�J8(@r��YR���n%D*74�����(�(#HYy��Q����m8�d��H�n+B���3%iEVZ[�#�)B�Y�\�U/U��{��/D�ӿ*���ƒ�=�᭤Ae�4��&٣����4Tb�H+�][[��Ri�ɲ
t�[P	{i�x�6����C,��z�R2=+.��"WLk�u���[��� �U	V+X4���i�vf�3���u���+�Y�å�tiDcr��I��y�u���T`3�7��2 hX���ˬ�	9N���'�b�m�uu��e��e�q�i*��l5��4V0pV6��n���'�w�"hZ������e;e���Ue�L��+kUJ4��]��n�u�f�b�j�N5���(��XǑBN��ڽ����
�CM^�LTWz*B�V���,KV�M�M^��{),%ƫF�7[�S�u ��mP���V�X��̭�٪�䂝/�ײ%VS4�=�0B�]۪tZZ��jV�n��
�.Da�Q�wZ=kj�`@'�u�p��I�-�:� v��ƍCE5b�����	��x���RD�fS�tt�R&�����V,Q{)[�q�5)f�)C���٣v+��5�tvDB���Z*m���ȍ�x�L�Qӊ�ܶ§׌�j�5��Wf�P�K%Jq�������b����#t�aH9d����`lFd����r�K	�.�/4�7o[f�")��fѰ�ޱ)��2�c̛�����	�L����a���7stJ:�[5�.@�0��3�N�fT�wel�jcq1�2�bj7B��r̬�(�)�{��i;Q�Ef�y�%�;z�1�"v�q8���^�P�΅i�Z��uu�fc!�{�: h���Ǔ&�V���W�v�3@[ۧ�+�¦|b���6�9y�Pt-��4fL{6Rnh��=YWt*d��V+�b���7p�QTԮ�z�N���ҍjl�<5,���ҸH���u5яU��+5�P�Ҿ�b.%��Gy�j�טa��ݑi[E�YZ&l���1����2Gn����{y -1W
��f�Sհ�Pfݶ]M�%F�(�	I�f�lX�/2��w�S:�Z��x��g#����3��WXc�D4��C^h�&����0\ڴ�m喚LD)�#-,�*h�fe[���X�]��efBtj���n�fYC/ਲ਼S�0`��X���ȺȠK�EX��w\���X��$i���B4J����"�R��ҒۂU��t�7/b��¬sP��w�qb����hL��x�Q����h仢���v��]�u���c�7T�0(
���>�@b�� ��%�6��omK��)B�V<���V��%�tT1�źf����%�AP�&�%�͆�f�eLD$jҳ/Zxj4��MAJUl�#�v���l��QVQ[*Ƶ�mଫ�MI��V��4x��f�E֘!!��&mEL�m=�r��[,����i8KT H��\��F`�h ���>�y�{�Ыv��t�x��ʅ[l�abZ��6����0��+.�Yi���ň�q�f�j��H@�l�����]M5�EY�-ف�*�ٚ�Q��
�C&j:��������E9��73:��Z^؍�7���c6�BB��x�A�2���9Vd[jl�¢Hc���8k�h���:�ڍD�Ь_΍<�!�v��p��[)Xz����j�D
	ɓeA�1b#%��&��m�e����ӤkFШUc��K��X�<ښ]f�@���v �9�61���vZ�v�K8��"��'-C���`*a ��l�L7yKh�� V۲�7�hl�/Z�A�L�Ҏ����Y��j�����
tk9w����f�)9��je�o4��V�4i�����v��R*�I��
�Y_*b�ܛ.���7(��Ts6�Ϋr���u{�9K&6��ѹ�԰VJ��F�����N�8�Rl��Cn�^l²;R�F���ࡣ^	5��k	����)��$���	����63*��W�N���Q�oc	�JK

��V�v�Zr�Rͽ�f��֦��h�He׭=&�#4�Rf�l��섄
�*Q�rSgCt��]8�6SZfw[S4P�A��D��cZ�B4&e���F�J�ݠ�s�h�G���N���;GU�.JL�������{O+���е�B �b|I�Y(c���J+�Q̈́�3+m5��-��)A�2����l6�vL�	����5�VY�JV�S�Ӭ���;{*j?J�],�h�ã0�L�.*��Y:NS�n.j�0'�䀫�=C���O	���EYqYw���+��_B�@��0e5����,���V�L-qʙ�3
�i��7k�)���C��Fmf<(Ф�mк��I54lCVht̰G{�(\�_K����;7Q�Mk�P��lZ¡���i���%��H�^�R4%� ���i�I���VL1�5r�֫&�ߟ�̭��Y�*��6�YY#c#��	�m3�jĨݜ��kj��pJŷ1�'b,q��? �?�T��t]vj=�j��:r�Irˋl�A[A��%�ͧ@^�T.�l����2JAi���:2�c�r:gH����R-Hޫ*F�����N���JK� :��(�H��-��Ve�AYictﾗ��e!֩�1u��͔��MR�Ѭ6�*b�C��/Jl��Yڸkc�m�������jĬn��� ����r��f��Ak�6�K{ �L%#n�n���P�f�\�16�r�^��Di�Yb��2EGl��ݎ�ה�f�@Q��-��dwwˎ�ډ	D	J�k�ٯP��*��!���Ru��7�Zp����XD?m����]�%�J�'xn�SW�-����aЂ���4�� WFd��R�b�z���zGC;�f �3PHʲ�}+(��m����əXs1�6�U�>��O.�(��gj�s*Q����{�.	֊�2[z���E^�l�T@so#B�,�w��WMʿ�B�	�����Ӭ�4������� �]�-f�,W�j���&'��t��K��%7c�/m\�m̫��Y��_����2M�����fuZ'h�έpwu��(޼���9��Ү��C���L_Ro5�Ვ���:�����	���Lt=B+$�Y��r���U�B�x�ͩ��������`��{�􎥦rj\s�s{������­���WZS}Ng`��[<1�WBm�dg���<�v����pS��Q!��p5ծ�L�[z;,��h�B22�\߶�G���<WR�� X��޾�7�Z�Ȫu\�t��:�2�;Nd�����i�:s�Ty�!Ov��Z���j"�y���b�36i�ŋ�Ӽ��f������h��g,����d��R��I۔sw�[]Kw'0p�:����o����������چ�ʗw3�KWe�W�"t�R�Н��=ѕ�ӱW���K*�N���,�P������)[>Ghd��w�/2>�=��z�e�% �ں_���B������ӥ�X�D���ڔ ,�H�hky2����읜oe�(�B��M�y���\�1��v�*k�Ԕ�{��]�� �4��gBӏB�
���j�n+�k���9+�����f.�t�l��c��I��wq�i�8��#�3��,�6�s�����s�Gigj/�)��ߋ�V<و�g��Ƃ�}��[K]]S�Ŵ,�$�w+��@�m�Ύ�K⩼�+�tMb�U��� ��Q����+�x�FL䶲`�RJ�t�{�*{4
|�;{��J}�b�k���-��Ap��9KT���m$�d������#�X�GWj�}m�,�p��ӳ���Bp������5�T�Yە�vݖ�8b嗲�9"Z¥�H�H�*u��2���]��4\����*���\,ΠΧ�6G��rB�u����tWbl	��^p͝Z��\z1^�9�^�Ǎ:Uɴ���`��vp4)[����b��F�������t�y�'�k&��Ǎ<�"Ywي�f�d���s�ή�*r�m�1���W�%�GS�H�͔��
�;��aYFwB(`�t�����*^u�\��$�8.��_Rw��B���ʲ�����ǽn�hwH{s�����ᓫ6�+�*�E;�.,�4�W8$D�G�`X���P�l�ø^���$�,Uq�`��$k�ܻ�#s�]�Ur��jJ�=�@\VH�^�+kM��5�$�@ޤ�'�ὙDpc��ӛw����;�C(��Uۘ���h�g*�8j���8+p��`�[���-�F�8��)�A2�H�e���d]��j��\M�����չ�M���;9�r��bs&�6��P��W>@LʏΖ�8�X̛�ObU0��-9�J܆�1��o*��Xs$��U�r�u�b�&��sD�o)T2P��M�����kh:Ӧ��9�����k�z'�X	��He�Nsm�/��K��� ��j`����h�����Ol�%�HS<�k�֓�;�O���#�rk(�����敒M靽�I��"Ƶ�Hm�Z<YC�Nw5ˀ����s�/8]��Љ�r��Y�q�>�z�	c������n�A%&6���xu���^�Q�£�q603�A��{����P����b��C�Z�F��]z�΍��e cwwj(��gEۓw����nU�il�qd�.�ݳ+d8����#DX�e=̈T{NT*�ν��M�g6�RTt/��1
7" p��h-�u�Eų��M��(=!@�m3�v��y/{�c�R`P����tv.�wl�C��nw�C+�3"�8"��/�Lъ�y"v��5A\��8�o\o ��u����f���5���0��Q�]Ս;}]�Q�r�h�hŜQw�r�0%Y�e�����Y�C�J%9M]"s���΁�`�wĖ[�N��B�[�����V�S��o=R�.E�$4�U E�#����P�C{2;��/f�G��e��ZZ1��B�w\��U�|u�x��t{(uA�5��*�0nܡa*��X/H#�ct��S�S�ߔh5��f+��dŌ������7\)�c�o���e�3*��F�r�ӵ�,\�:��k�1򸮣�X������6�]g�JxMwk��da�}��u������o��"��"���V�Nr�C2W9�n�v!l�Gy���D��3��ۃq��g(���R�	��a�YyJk�9�:�-N���q��/NIX�R�=�����xU�Ֆ/2��׍���GYw ���G��4e_k�@`�����F+����4>���XE�ht��I�\�#\8�.�Û�je�cC|��t�����w�Im]�2��J[��N����6��f_�z㵺��p�R�N�
[�o:P-��(�ï�VJ��zݥf�pTY7U:SEi1�#B{r�:=�.��o$mɇ�j���A0�A/�uxoh�lM�eE��n��_rL��D��0�	��N忺��m�z��X	�]9��)��!q�@�N�^����srn��"\�X��OwS�F������ց�&se
�Rv�ol(�U�@"ݻc�m7���B�ѲT�%r[��VBU&=^�L��s���F.�&͡Ɩ�@�u�Nǖn�Z��L����gN���4�ۛ��]���u��HV���A�}��C�2a��aG
�dn=���C�4�{��
K8���yҦ�];}B���)R�4����ǓE+$Z��LNW�t.^-�ٛ�do!k-C�ИЫICM8v=�a>:2P��F̬�h�E�"�\ʃ�94�E��_m�Ҹ̧���ae�q����
Ԛ�tr�M����6+]RU�]m��l�=T8�ե^��4���6g�(�ܯi<��FT���������dU�{�7���Xn�!\���D�zy����e�]���Q��;���o��N�]��@s�حFM*�5�)���b�9�F`����"�d��'���*�.� �mq����S- �Zj��w|A/3O,�����)Z�ι�S!-ł���k2ʺ��4:�v*��j��n�+�}-Q#��'�j������C{�X�GXju���p�P"U�Qm�%���;i*��[�r�E^ert^�or*�����n�t�����ܘ)P5K�����n�f=u��������8-���H����H(%H�5C�]%��[�f۪wwm�N8d�FT�p�G@%d�B�օ��M��ZZ�r���+4�ڶWS�Y���^��<��N����㍉@ųC]��k�Tz�jZ���2�B��{�U^&5nfrr�A�] ��6��L���m^_�㛿:ET����'��q���G��ZQ�%�t�x̛\$�v��r��i7�9v��f��L�,�}հҵ�)
 ����M/��"�f��1)I�o*x��^�͵[�����Dw)�68)�FB�z�`뗍��Z��nZO����J�a�e���r�K�TV����z�9��t.F'��꡵�(��|ͬS��u}�f����i�-��1�a�ݝf��b�=*�aG��R���Xjm���N��&$\�p���4�}*i�27X�{Ww1`�N�\����'�f��J{\��t:���o]7�s���%Ӧ�� \��\�ܳ�:���ky�˹Q�4�"��B�]Z�m!�i�������B�R!�dL�y����c���o�q��T,X�ɤP|� �)�4��ۢ&H�^��R8at�G`� ��l�?r�\lnj4un��k�c��e�����(j�g��Eer�5Ϣ�b,�P	�`c.�07��� �[ils�Y�D�����6[[�x
Do;7�ƦB#'V@%6A���_w`�v�T��#���V��Q6k�b��:u���6�ҩ�y��)��hPr �I�p����:�]pD�K�N��'��^w�_������4�K��j:�T��;%���w!{73�l>MäS e�\���J�[��e^7�t�|�Ս9Y/c�|��{�t64R��f����9Aँ��z�*�qШ����8[޷�#��U��`{���×;��
]<�IB�]W��A�N�g2O:��-���)�I�B�cs>V���=��\:��u��t��a�^
��՛׍f6����`�}� }�VM3�:���W��h�z��n^4kv6�A']e� ��P��M�Ե���+��s��ir��������g�P�AY;����iFtr#G;�"4�<�{��̝@��P��]�+��Ս#ff�7ڹ=Ӥ�ك�D�]�Q�ᛢ˔�����iJ�)]�|9�&��!�K�o��a�a��v�\�J S�u�KHͳ�bJZ��A�CFM�3Uq��gM��4
��[оU��LX�眴�j!3���ѢR��8 yz�\�ŉ�J�h���d��U��{7d{��4N���ɜʳ�V�p�lr���&��*�C�@�l�K����]%*��N�]f��	��g���{n��E��h�V���RNu}����J���(A[�2�XS��T���>�**�:>]�L�n�ɎA+�*&mI��E���@�Y^�=/ ںXGt��ks�x�-�L��{y�ݵ�P(z�QJ�U�z�0��Pj��s�]N���J[��.e> �5f=˙�����6�&S0;쬥�-��(�z��cs3��m�:wA�2�;������1ߣOs��+u&GJ��i;�T�N��v��k� �!ج;����N}���*�9NU
�������Pq���f��n	ˈ��Q�r�86\|�˖���%w �U�3�o��TZ ,�6����Z���Z�5��K��u�b�us��$���͜$}:�G3j2+c��-��.�:M1����7��XV�ǪV�,.�&���^��؂k�jQ|��+keҖ�ٵk���$�kiM�=}K���]��H"�$@w-o�6�#&�b���3���Ә��+6�fv���9|:@���V���+q>�]�q�oO��s�g�)�C��mڭ��6];u��):�\���B�#bWvV ��.�;X��Z7���p��EP N�z2B�:��+
ٝ&f�#�,����Bf����n�#4ȋ]�{ [k�;V��}}ט���S��s�,���\,%*\�Md�꜈켒�S;��zrm�uv>�N�����]fA2�J!=���U��V+к��]Ε�.s�n��+]�I
�7W|�s`�C��p
x�cI.��%n� >��ʜ�m.����%zN]\\�@��qN��s	��'L}����⣊�b�t��=g�w���b	��H�Ԟ���Sn��,���/�m��Xp��*��Af����ooTBc��y{0��>r��S�4��R�@��2����z�[M�ؖ�4Va{���X�D�+fD��U�R���^��mɥ�ѡi{yX�t���y!��r֪��{Cu�m���I E�����u1��l�xNXz�g3�&Iǘ::�]��=G��.w=�?m-I���*�֦�ϖ=���.Р�3.9fҹ�+;+M)\1�o���bm-{��0��f��pvc�ǀ�7K�L&o>޽�ؚoe���
c�e�(��V���"Zԩd�=f���#�<̝��6�8� �������q�f���8���<�x�CB`��N�VD|�-�±
�F��p�y�O"삳e�Uܿ�"kAw�#�MvGG'O������ky�L�wΰ��YSh����4Ɉ�����da�����d-V���-^1������e+4��r�u5&G�	]B��-U�@/,Q��NZ]�^Z�!���
:P�m��WO��.���rKg8ܓ�k̾תݓ%`�8��Ѽh>�L\�V�:�����{�X��+�I�u:؅� ��;!�o&��ʃ;r�S'��J��ng#�)����Ƹj��.ݜ�1�#z�J��KrtN��0΀l`
0o��vh���:nwP59p*;���#�|��B���;��
JD�W${�}ĳ.5���,,vIu0�6�(S��O�Z���D��:�438���gz��L�oa���*� �Q�+��L̥ٙJ�S��vwc;q#�<���|t�y�N����N�����U�S����WT�2j<��7U�t�Z��j�7�j�f<���<(VԨ{�ҭӚ	��ө�'5�}j����; ڷ��{���dn���1C�5{�p�d��%N�Ƿ� 8.�$�Y{7����:��wQ<;��X,`\5[Ƣ�N��|��.���	
����r����Ml�/�\�rh�#|;��`6���1�c:)F���o��s�	����Wx�ok�P9V��!:���������.��@}u�Vm�yl�J�wyB*�1݇�$DJ���ohHt�o���8	˓���W5��/x^��y�y�+R�W{[�,��RBoq���/m�̇�pK��7���BtyV���pC� ��\��;��j�ږ�CG;Pc��t�$��v�M]�RT��#��+
��T�Id*s�F����B��낂�/����{�qz���b�4�b�����c�a��W�H����.���c��*�}��$ ����J2+L���5�'A�wo1w[��.�C�ӹp��("�����qs��ء"���o�3����؉e��f��}����;4�͍$ni�;����&��P��N�T�ӽ���ua�:��-]�.k�(�!�a/q��7���;s�����VK;mDfCٮ�;SD�����|���k��64h���u/�T��7Jtv���bu�C���!��s�ј.�1e�E�����Ȯ`�wSe��H�J��PH�DGzbuo!��/Jt)�U�x�ĨJ�w�	�
:�zmq����ݶs��1��'�t�R��H۾Rë�m=���r�Y�6���J9�OR���9����HHI!!��$����~~|ʚ�7�X�
��7z�n�;%�v2�q�㣝�E��������>�G�maUAz��t�͡Wz *�L҃�Q٫�f��4�%�ݼ�V)2��Goj�o!s\n�Z�J�����Ɏ�4�5��jI�I��@%��>�N�T)�V(.�|{1%N�ɔ�`��f$�,�# �cr���Щ8�mf7L5WwO���Z�V�,:�1�j�&�L[���XԷ�&�
�����0h���d�/%'�`�pp��������>��6��p�m�%YmɗI�4�'���۵��k<fŔ�"�u����u��#[�|����Oonu:[�Ec7@�vE$��7L"U�(��s�gÆ���nGOo������V2UH�0aG�Q�v�ҕt�b��L��غ�W��$���/J=2���<�I^��s���1ɥ��֎8���k>��,T��MN���wF���82�9l[�goWd�j�K*(��)�kM�¤��΄��j�n�Y�d�4��C�]�eN�u8�w��`�F(�sv�U�cj��L)o
���
iq�*�Υ.m��R��϶����	K�DOfR� gZ�{�+�)<͝��:AEig M6�̬�\4�q⥙��d95�U�MJ��PvH���[�YV�T��ȸ��{PhX�Γ:9��a�p�B��Pwn�i��d��gw"��-���+w��Q��|���*;z��b��g��:u&n��f�u��.���QYeWN�[�.}b���
�t
� ��f٫����V��l���4�^�qV��m�a1������W��\�s~�R�t��}0d��V�Ꭷgmk�\p�
zS�4pޅ<��ϭ�y��/i����ΩM$PZ�a�/m${�d�Z3Q]��khdCz�
hF���0�h&|Jϸ�Ҩ�}{YSu�sի,'�A�%{p���.1�ةWQe`�ڵXaz�����#n�V{A��Zt�7�[�����n���r�LxC�Q9E����;�Wk�+�=Ҫ
�r��}-)ф�.��2�r��"�m�K{�b�r�5�1�A2�B,�}&`�l=�e�N���O1�����P�!�5e��)�xά�z	���������I,�ǚ��SIvJX嫵Wj��!· �Z�	7��Ll�u��c�+�r(��wx�H�	1�2�΅'roQ�m����C���w�K�E��i� 0]�z��O�<L�>*l��*�+#��%�/�{"�@�8a�%Yp�(�lo���)+����+LJ�U�g�����ԤB }��M������LD�#�s�md{�-+̰+!�\���(a����Ԫ���F˳T�<(��|ݮu�u:���cf���5�d޽Ru�e����;3'&�&��B��`��+5p.�sj�L.�@9�{��r5�@j� �Va�u���E9���.�Z�ͱa1�P��8���gD>D�O�����}[k��5jG�'fN����Zņ�u����F��7����+0]s���2(*�ɊJ ��3_jz*8��ZK߭B���y��|7ve�����]z�Ȼ�1ک��eՍ����/���m˹@��M���銈7;�e0pi�M[n'�45�N5��.�I�e�Мw1��]@�ٙgByLm�iO7:������R..�5��,;X�b��G��:�z�]ϴkC��y[��딷y��Ļi�b̈��C:�S�q�A�!�ǔ���P`}˗��6��2>�T/��:��B�3�W*[��F"���C��E��:��5;�_u�dIIq v�6J̮}�b)�v�M��M9,�@��i��g8)x��`V)}�0���j:��:��lF�|�.��u��X3 �^b���su�U�'��N���8�e*�]
��^� l&�&ռ�|������@S J�J��sd���#�^f�ri��ED��vg[_t��E�B�I�����X��+�d�j]��յ�uk۬@FU�Y�\�F:S�ɱQ�WQ���.�c{w����V�Dc���Œr#nI��"����yα3�^�Pٓ�Y���CC]��9�˝������8Sq)K����B�GHT�8�9X��ghY[z�K��*�x�4�&��9�Ѻ�z�m���s�IC��d.���A�dY&����T��E�W�@�\�☁&��Gk5KC���-�|�S���kdϯ7IV�Rc��l-=�p��@KV�s��XZ�JU�o�v�٤M����pj^�ӝժ�~L֚���4�gj��/��ն*��9�1�����Eƒ땃�IӲ/����B�Hu��I\��W�)h�2vtP�:Ƀ�&��]��sj(Hέʚ�[hmo�c1*�Rif�\�,l87�6l\3+{�:�Z;�Q}�X��d{�xv�Se��1�V1�;W�uܓ{�n��8ma;��'�-<\�nQ��ݕ�V,]N��]���@oU[@*-�ܧi��2i��`�����O��\������(j��P�Ԗ���z6���ʭ�Z�2���;�M�j�T����{'=���CL�p��H�FVU�7�m�!�Mݴ�a�ɩ�����Ba��4�y�o-�t�Qof�o(r�h8{Uec��H�����^!�b��t=v!N�E]��o�fV^Cz�s���LJ�N�̗�v�w��tn��4te��-�MJ�%
B�9���ǂ�#���h˾�`㢒����#�:�\���-��Oͼ�Hޖ��O��89�&L�to�r�����=Z)�)�=m�a���	$�㊌�'T��ZR�e,�)f;)��+�Tu�ܥ+BR;�����ݻ���;V�Y!��$��	Z�VÐN۫�x����HW@�P���ysK-���l��Ef�+��fZs5uM4$�7�\�`��B�Ba٠��S -�y*E�m늺\f�3M�g
'.�S+n�T����^�u���K�+���[mn�n�ޫ�"�v���1)��&���3%����"�Ȇf��&k���Mi��eK!�.<kf3�������7��Hi��ƭax���Ѳ�Hg-�V�tԢ'j�{{U�{@�=�u��{���c7k�GbTPZ������t��u�|��
��2Xa��m���]ˊ,�6��J�B���҅Iڷ
�H�98�l��k&�Y�U��w|��;Ũ��hgb4O�ڧ�Ӟ�4
z��x݌�I�A]�7��wTӏ>����9}/��AuZ�
-���E�xڕŴ2��թm_LM4��3�GI�������t0վ�;]��}4��Ξ�E����D�M���V��7DZ�d�;(_ٹy:�hs�����*(;���1�Yo<ꃻq�e�p�ϓ|�"z�[����:	"�!��&��ns�5LeJ��U
jYX)�N�FN�}Ϩ:��+8G�J��˕fPZ��b��l��(_J9-3W�K�t��;�aމ��(3���8*�vG�1�%J��f�wm'���.��)�A�y:�V��M"��R�F�鷷&u��:�K����c����]�ue�ZgJwI��%��c�x;��*��ْ��ˤ�DsoM\r���G�9�֕��#+���,��C3����0p|�"vk�⯳�ǉG}�{v�5u�B,����NN��n�N��Ab�l�3�b|�P��M�71��f�Ӄnq�S�����1�wt�,�����O�tŰ�X����+>W�`���ق�{MwV��!\Nu�-n4iņ�u�� Z)�Ʀ����[�|5���i�߶�Gl&��j1�w�3rq�9�����p�����5ʛ�sm[×��e,&�h��RJ��]q�݃�ŧҷIf)ѥt5�*�g�^P��B��d��+*�49lG��g|�u�Zݡ|�+6Z�^[�[ug�Np@Sxֳ�+�b���෗�y$"s��7������X�ƣ�/e�qr�Q�;�x�(�V���6�]�ၰ�\X:�X���8�.�������0�`.�a��c݅VK8^�8�h2�UʇHгZ򹋭���'a@�m����{+;�8ѵӁ�ګ��eu97+f���l)�z*<6�M��C�a��+V�0J��@ѹ�G������q�Y�Yv�����~4�9�uǛ��p�gL�o�wy���צ��K>mІ�JHU�:#t��+�M���bz^Y�0�W_b�/8[Yq�s!$�����\�VG�6�H�6����pn7'rC�YM�+��:�Ss�4��z�5���/���U�\x2h��|r8V&�h�:SbO�w��Gg+�\�|vXr�<�U�ݽ�و��t�r�����wXEY�.�wy�ba���plN��$%w4pltP�̹(ww����zk �Z̧N�KB����c���̘Zy��drHeiv�;�]�W�up���������$ꝛ�4Y�A��^��ֺ|�8��4#PS+��Ԭa���3D�.��Ƭ�T��ȱ�����'�DM��3�������.T̢��t��c�H���+�JW���Zt-�ieu��A�+e�KD�|9*=���T2�^R���Ő6��W%�J��{��V��&h.�us&���\���pX2�oHO`n�:�C5i��g�UIS���b�˧���5+�4��'-<�B�s��.��m��i=B��	J��a�j��T��֎�.�)a�MQU����f�TLؒɚ�v����p�$*td���Q�Z2��$��"ZáP}&�@�Gu�v��o��(����Pl���d<ñv$X&
ī�eP��hCx��_n���Vs*5��]J�R\2�(>���$s�]��0�*��Lf8�5�-O�����N��K��iYi���PN$u�T�(�N���2@�wF&���=�j��D�NX�T�`�*�c�}� id��MmM-�r��|!�X�]Rm�k�����U���͊J����Q�f�]�D%�)GL�j7u������0"uٓ�!�'V 9�5�HC��u�	4��7�2D:vp�(F[
�E>��St���<���sg��7$��	����F�Crm]�ƪ���+8.�Ak��י(�[}�5b��E0#�1��,��t�Z�r��
����Q�.�z����S,�Wf%���V�G��n�n�w����$p�t�|��m\p�g��*а��ȻZ���b��)�y;����re�W[�[�ヾ�9��ć=Kl뤖�V�o�*J�[9����Y]�qU٠ڻ\
�7oZ�O�+4���#!�ZP-��$�I�SQ �N�v�v��V�`\��� �Y\C����)*;�3�J�\�>� �7���>Ma��Ge�Lކ�ޕ�V����t�ߖH]��į	�z����j_-��")����Q�d�WS�CVP���w�Z`�&���$'
Ǎ%�W��E��=�rM[7�4�����r�u�L�0={����S�)�
�}��e��n��a^����S�<��)�\�rN�
Α�#/*��U�{��sl��4	4���@���q@��XZ���9X�]5ݗC���T���{�T���6�I3c�^�Ǽ-�r�����<�s�/Cɏ�V���mNlwF6�uK��\"*̊���ƚ(�/���[�`֛��*E*ش���o�uJ��tx�i�������c�qtd+;Ud��]V����S}x��8;�N�I��n�n��ƚ7�%����A�!�qAX*٘*�����a�J�3pņ�-�C�:��ޫ�;�@���Sb��Y��y!�������oW��������б%[��F��:�׎r�Wxݸ�ԋ[��9BA�냤�㝹{;��4V�˶�.b��Y�6X}��fof��(#�-��7���˅;啋�-e�K
������I�M��Ƿ�x�ݎ�(e=à���l���=(����.$�SW�־kn��SY`u݄������*�LB�'i�`�o�+B�q�S�����V�]h}����䈛�
��c�&dg:S3:�p�v�u-�w�rWIRWCk%��aʚA�!�wd$����K{�5f�k�`'���,���IZ���*enMs�.w4� =4s�(��\t�m7�JF�Iaݜw4Sf=�_NT�ܣ"�y�:b��"sf�m4J�o)fw;���I�[��ݝE���0#�M��-��	�J�CB�[X�є�7��Y�%���K7X�{̳m6��;�L	�v���<U4�rm��Y]xx�J��\	�tF�NJ�q�J��R��fҡ�^�LP$�L�J�5�i�!�|�	�&ʛ45%o�s�:�;oi9�wm��<;Wt�4������y�)B�^�J�]֕�v@��p��a���Ԧ�.�J�ѭM��2>�}GSFD��k;�"����b����IV��_P1���!0�6U�*�%�	���P��|�4��V��3CŭK%�t��Ț��A�:eoAU`�BfB��i�g�\� c�|E#���۸�Cᘸ�ӆem5r���WpGTz�N��2ZR�ܳǞ�|��۠��Y���_HHu����*��0�x,��Z�7��s��j���j�M����X�g�G�"���/�f��[rN�����������r==��V�WV=��6��q(�GF��LV+[����&GG7^�Z1ԛ��P�2:��ʊ��p.5�*59�F�Y��S����(8�����U���D@��ۥ�֭�h��}�&`3��烜�HN��b
R��T�+2�2�����Fē�J���p�\F����^`�+��#{�DgWmﴵ���*�W㈓��J����e)]4����䆦��?�{�����սD�I�U��!\y��%$I��b���=�5d�n��;��&�C�HʇvHb�,��D�ӂ��3�fN��!�³���M%fb�����݉��J���R��#|���#�B�;I����m1�AYt�f��pqpa.��3����u�F<ʺ�����<0\ٍRN��fR����'�\ڣ�ҩ�Y�!�#�gXω��ku�K��d��μ��`�U݄��X%�@$~��6�nCG������f������NQ�������9���[;f �d&v�GE�p۲0�}	�|�K�7,�\
tG��W��[����n���vnRT���W����8���ܷ�.��m#�߃�r�x�]j
Hk']t�X��|������4�d�^L������(	��]� �B=&��)Ҷ �͠�ta�.5�=�'a[�>��v�wI3Ʋ���n�4�^.��F��O�{D.�ng�`���<8��];�I��+z��-S�gvPN�f�-�� Ddu�Kh�/�@:d��hSU�6���ɻ�8ңO���ܶ���QE��Y�Ié*fs7`u��C*��!Rq�������,�_vL>nq:z��|R�"�Ru�)��;�<����=����IW˱�.���k";pP�Gk���Csn�/��w]�;�	ɾ���n�.
�-��^��+�T����C쥌U�*Q����b�Eq(*2�_�V"�7-��1WT��J�em��%�ѤGMTEUPb9J#��q����*�Q-��Z��3*��T�������)R����***0UTQ��U[ljQA���5e��1�* ���\n%E��BҊ�c����ֵֶA5�[,X�M��R�`�c(���j.
ʙlEm1�iR�����h)b��Tt�V
j��X���bccPr�D�U1��T5m�Db���
����YQUF����*�*(�U�R)4�(�%B�2�,��(�J�D`�*����*꒎Z(�j�D�����A�lE��\c�X����MQĸ��D\�Q2,V�QЪ"�UT*Tj���Sb3V����R&��
����Ep�Q#"�1m�b1�,ib�Z�UEe�LU�]YA�	A̹[[��}���Q4~5p^�'�m�k��)�FGw���U0Z�*�JU�d���4�D�c�]Ϙ[M�w���ʽk6v=�㹼{��54E�Y��D�!�ڮ��5��2�
u'm�Ό�Vx�%>��9q���mΓ��m�Y�q�b�{�E�c�~�,���ߞ���
�:�KΚG8d��ͯN�z��z}��Ⱥ����6a�J?�p���t"��;��]���%�i��pG����y���Fmv�aϳ����-����t�H�R9
*����qp�ʧ7a�� �[6�a��C�5�������wXf�ˠȷ1mm���u��MDp�B&whAC	�Qu\]�䤑݋�!���թrO�&+z��1��ǡ�klOO�y:xB9�8U���:�]QOV2��,Y;ޢ����Ώ����s)lw1�	X9���t�{���L������YA!�<�������$�#8������:+��']v��}Y;ɺv�+��	ཙ��W������߮0�6��\RY"#��^�꘤!�E��COv��Ø���z/0����O�i�gg�:U˨�&@ 8
�|RQ�xr}��lW�;�.x��fkvqP@�[,n"�&cU��c��.3V�����!�渣<�Z� �=)D+sd�����;���xo'eI���H�q�Ց,���R�Z�枼<j4�n������-�P�gB$�D�_���ʲ��p��r)@�Il�#���X��aɜ���x��pYX�m�)�q7A0&I��aӃ"�4rs�4�o� �-iku��=D�9ӆܾ�W��L����J��B5P0ׯ�����e�;�zUGdq07�-&�R�8͸�nu�{�D`�թP��3�#e��l<̛3B�����Fn��m�>Ar �}�VB+���I��Y�T�n|U��M���}��{u+z��1��,4,��E8������uF/��x�'��{B��tؖ�_-=��I"sO�Wo�q�(TrN�bB�P ���"Ĺ�W������n���ydŕ�8��>�\.)����:q#����63D����WH�wҬά^)���'��a�̉�8���eזJ������O��_����m�U�Nhf���:�R9mY�v^��Wƾ��#�.��$͕t/k�22܆h�8�Q|�Z�$f�*���O�+�'�{� �Rݠ�r�sU����]&��)w��T����,��w��M��!�4o�&��S��VoV�rDx�w�7�@�]Zָ�pb7�,��6���弔z������+[6��z]A{"�=g�c�H\E�0Z��p��CX��Qtﬄ����jw>��M34:���J1H���QM�נ�Z��{�t�y�k��Q�#�K��W\uHQ�T�T!q&�d���rS���`2h�����Q���0+"�Y�WBH����zb�.�8�����*�h-��i_�9Ӑ]Ak�W��k���j�5aT��Ed��x]즱Oy�>΃oEA��9W.SQ�AW��S�獴W�����Q�}ssqw��� ��s�y��`�PɀU�FB�U>�	Ж�Ls��E�5��a�_yV��>=��ݙ�[���h�j)���
t�TQֻvU�f�3�Y�����F#cV�Pt32�3{��$��I���K�f'��$j$��ϐ�p�#�<��R/�u�n�z>�e��]�HQ��pV��d�Tۭ%�!vx�%ڨ)��IP����4���<`��۵j1���5�o�L_R~��#^ӄ�C<�-��r�&z+�3�E!�dQk��y�m=荣�,�]ݗЦ�Ė;�dr��v%�z��>�Jp:�X���BR5rR��V��ӴQw�=���]�L�r�؎�#G#7�N�GI_���[�+�f�aB�Zu��o���Q7�xr�Y�$�0��j�%��Ω�����]��$a̬R1Үv�%G�_<��hH���L���7כgvV٬[���y:�զ����kZ�u|Ez�������?�<���{�eN �]SàX��8��þi�0��*�`d�E[���K��i�^�������s�]����X����ѻ4���.��H}��;hVM����gu�,^�a
"���5C2���t"]��3�'+���j﷏���h5_��Z�-��(���~;UGIa����\X[K7�2��麈�ݸA
( Ս��n��^�B�4�Wz#��1܇�v��泻����s�����E��d����*��5д���94V��s�nk�	��X�"y	D��gbV�0���c�ˬbsG�s�f�s�St�;n̵�+H�qF���MM-�Y�Y�+����.�Re���%ة���������³UÌ����U,��c�24���b&0�P������	�z�A]�gfBk��ؽ>.�P�7�LLf�=�Q�!\����o�`�c���#�W�5�y��c4��T��M�E��� �z��ۏ�V�>���͏,��%E�Va�p`�mc���a�^ΕDNt��v>�s֪�ny�N���ݍ-K
�zaξ0jjv
������2�{�G,��<��[�Mˎ��)EY
���[�&���&������p�rJ�;lE͈j1kU��V�F�v��i�O�T�!�ȍ���z߲N��.]�ň�֭��ه���.2U;mW��Xqȟ6�F8���D.R��>PɂɗV̮寭]=K7Ap��I�����2�����}���Ji�m��S�="33�Q�עj�39�5��7
�16�m�"
}5�M����R,�kez_t����`ӣ����VW���l]�n *��LtE*� �Xˌ!�4~΅�ȯ^�mW]�kӰ����:O8��8D�י��g��V���Y4C��~�ih>�W�qGk�\�,�/���:Q�Gid�Њ���Wȴ�n�efp�n�]�?jYw;�uU�C��
���^슖lL����vUokhe�X�@`q��F�Y��wŸ�a9�ET�k�� �|+��M���$mf��}�%���3�ǉ��ɑX��7]E��kl74wlk��J�ӌo�z������S�.��Z��<Fjf)E��Y�ZL
ޭj�Os�ᵚ'�׊ٓ�TD���(�9&�]�^c\G�=����N�ʔ*�R��]r�D�m�Ч�´]wQ���<����4x�9`.��2�9�-Sv6�t�1dCK���%}��s�0WY5���o ���5�m���CH�o�
�K����%K��>gz�C�
+l�cɆ�R今��	a!3�Ӝ���[1}ȇ�b��A�hsB^��H2v�]�gU��l˒2���pnSIb�Z���ȇ��W.��Ӻ=�Oj�9ݙ�2���&���4*K;b.p��!W�LG��Ϯ�s�7��=J*7o��Nԧ6'��RbF7OS�x���w�8�J�uEj�hD�K��6WD�������z��q�������cm��\:rgM��>J��
��σ��t�����(y���/>��W��t�k��l$d��t!�s�=.�����kvH�z&N�	�]R',��')y���(H��i|�8͸�nu�u�tF���,:@C��[�=��C�U38��p��� �%{�O��FvK�D$;AY��Sq�S]e*����}�)���\2`�������R�:k��7ȧTx�~���;,Oev�L+�������,Fn���bj�L�G4�Pm�:و85
Ib�/��H�;�C��ٰ����.������&k�	���n�6]��N�L��^����6�h���SU��JW+���o
���	k���>�U�m����+�{\���\a��ro>��z��@�ȳ��NC�T�!���զ�'�:�X�̢�Q��}�/�H�(��Xv���g�z
9�Jy�F�y� S�
��R��E,�	ޒ�`��)Mj�z������b�������Ŝ�E����ru��|rm՚�[�O���6�fÃ�]F�l ;�WƊ�C�� K��t/k�2[���㐤���Q&*��f��jzwn�Yg\t�7�7�>�sS�a��A@�R�O��X=�f�8 ��K!�N��FS����Y���"1 �}��!5fc�3���l��2�.�����|m�U�(��"��M>��}�oF�D�Ҁ�.��:�=A=B��ӕ�P�Ю��'K��=W�%ɍ*̀q{��BwN��Uz��|��G���k�6�����`!X�h�S�Aݝ��&����;������"̈��j�nW*��	*Gk�}A�v�w�Q,u�k!��}p���N�,@���`SgĘ�`�HU!����u-ޘ4�6k��K�-�+ZI+�6��{�vN{B�(���t-X��"��=щX(�]vO�ϯ�ЇF�����<sR����Xoq5t� ��n����u�ե��f|f��8��^4�%SM�1\��:�PY�3�_`�1aB����G�]L�i���41��p��.�$0'R�X֦�����ʸvQ��x��7�N��L��B:�fD8c����C��3���&,0w�p�#x�x���D�$�Y�wN1q`}� �Joo�в����J��*�y����ҲM\QM�ZM8��I��!�L�`�k�8
8��6�y��#%G���6ᣎ�7Pf�1��B�6��'���.��,�R�^b�.�%��\S�٩����g�ipE�/��0���:P��-�Bӥ	W���]����	�@���,qHز�õ[凎H���3y2\D����3���u{��/=�n��1�r�u���_U���?:^Y��\+�Gჰ�>^��)8$V�N��F���7��V]�+N�{ʘq�B�q7A���X��Qj�VȻ��j�Vl"}���Ij+Q�t*_��Ȍ����>�9�!��x4�z��pvS��o����ldͬⓩ��hUDaj�(��ss��mgĺ�>�����N�S�z�g7�Ó�����0+�,ߦmS�d��˚eC��cH��s��(a��by��Z�µ���{�3�t�ؔ�u�*Ɖ��eIj���/4�Rxr�X�4�J�x��{�/]�[��+ۻX�)�97q�<�Z��r��K�M*�W�Z���y�73D���C3��[C;�;׺��	3=����K3���5�
�}6��~��Ѣ����D�t�]x��������&:2�˘{ݯ�m���dX�֖�(
�|~�T|-�!A�).�@ۛ<�����fZC�yZ�"��|���>���C )E�"ؤ��Q*�c�N[�5�(y�1������`�My�~aUyÖ�3�uVK��\L��w.��Z��c=�Wrx���gE��_�X)�F:�ry6��;u�8�Q#�
"4#�g���"6o;p�#^�����E"�ĩ�]�sz]6���!�,���s-A����TF�B��ľܥ���cг\I��!���]'��!��<m��MX(�K��O���*��huw���o�5�ֈb�t'@��1���
E�""�Җ�X%�|����J�3�ӌے��vN�'oe�6 ��2+ ]�DR���A�T�v�b�2�3�C2��_c�{�q��7��YQ ��vPd"N��p���M�.׎���^�Fԓ��e�"�NdK5��PV�U�n�J%B�{�U\��j����ƶ��xkk�>u�\)�6e�6=�ػc�k�N �k۽�{΅���{C's9	��\@�$A��T�+����0f����S�l��:��іl>��fï�˜���X��k{܋�otwa�_�b��Ϋ�9%¯Z�����%��3�g�/��=vM�W�����7��N��$�o��M&3N*�.��lE���B�2E�B��8�!x}g4ddF۾��+��#����P�V�*~��Ȭ}a��9t�-��ܫ�x�-�ΗnC�F���zN�ON���1�UpUB��������h�3XV*v�y��S��wxnV2{件�ɝf�W��N}Ǯ��`%#� �Q�P��t���}ȇy�_g��!�t������Z|���[��cH^�Z�N���es���:)D�p�܄T
oxZ��<�f%�)x��g��hp���؋�;@�H@�����%�W�Wc�wf�XR-ժ��'
�����D*ka��j�U��3��hq��]@�+T�B%�u�q�b��"n��9���%��(b��٪��]93���<HsT8)�>�j�W%FXQ���2يT�3��D�kq?PD�Q25ĉů����a;��n_W����XnwR#������b�JC��F��<��&���GT�km�\yE�a`I��Q�ɺ�v*���W�l�C�;�&��*�dH����5Ohu�Z�س6�2����6㷛��ĵrAӱ������D�(�
d7Oc�2^s"�n���s�o�,d�RQ������	E�v�@� 	3jY�: 
^2n�s��F�JXH�JX���L��d�Ū�hiX���o`P���݆��8b{�n�;����x{:63��b�������9M���퍺d��iN����=:�Zv�[��	F�oA9������N�z��w.�N�3w;t�;K8=��\3'`�����i법�fs��ֺ�m�Z�D8tJ�x������f�9N3#�m����O���ѭ����0e����6��b�
."$ꖱI	,�w@L8��Z��;�n�a�pV�����h�D���$�)�@�T�f%1Ö%���Ev�����H�5�#F���8�[Βobf`��jr�#�f'eV7��=�7�wH�����)��ʗ׶��#���R��=�vɜ9c�N�ty�gm&Qu�ѷ(�9�z`�sz�8{)k�}oa�Rt0 k�/�4�3{����{�.��ŀ�ַ�n�0�N?��N9���m�WjY��b)<h��t�אV*�WQ��Y �a;E��u�)��n]��:r�=�ʼΜ6bj+��K���!̮��Rӝ�LW�IQ�������!�GRĶC��^��;��2RYIs�+�=V�y��ӳ���5���KBR0�6�!�/$7גĻ�!���I�ZR��&n��U�FX�7���K���SOAF��-E��!��B�d��E����2�4���4P��q05����V�ҋyw(Vc�����v���Q���Z��Yoފ��@���+Ui��H��D<%_HH�Of��:�&���wz7�Qw�W`˰�������9�Mdg��+�����q�lf���R��%Z��t�nV���F6�0
nc����y�1���݅�Zݛ30��e�\�CsBz�
դ�UC�����:&g`�e�q�enӦjw>�F�e��j6�:��8`͈a���t�o2UʝA�:ᇫv�hQ��T߱	k�{�)nL�N�k���9�GBd��}��rmu����؀�ʮP�d%G#}�Xw�����r���$���;�]�x��71���^6o�]o1���jڹ�Qj�C0bu�֨wa�s�,�Z��b���K���[
�C�A�2K�^;�0'8V�s��#�Ao�fv���$|V�Ox3a%���|��b.۝�i�#�n_qj-c��7��9\�wh�H�Ӈ��Ꝼ���7���mzqvt቙k����E�tp�l�\�n,�\�ݥÆC;�>���0�Pcph/D��Gn��fme��Vi-���9����;�����ʃ�M�>���;ߞ�񱈕�Tb�F�Tb��G/�P�EEFAk(�bi�Ҳ"��Y�cEDE����kcVV�[���[TV��d��UV�J1�V11��b�IX����b��Z��X��*��e%��]d�ˌE��iQKl"��J"��FZ6ň�e[TJ5�V
-U�DF�ms1r�(%���J�V�mX�m���j(��YQ�ũZ�*�3 ��U�lEcF֨�b�K)X����YDU2�`��1�YQ��"�TQ�f\KQ�������х[ETEm-J�"���V�"DKj���`�Q�cr �fV�Q`��F �E�
��TPVF��J�6؈��)ib��j�Pe��"�`�P�q�b�l)Z���eJ 0EQ��k�a�cD\eA3���k+��������<@���H�nM����G�x��kl���rB�a\{�f�2I#ͺ�(�mkЯowWZ|�ꪦs�O�ϼ���|��4����6z�$N0��ShbOM��dYY׈yi��LLH.����<�'�b�o	�M�^�}�y��A�N2}�1f2TP�����3g��ȁ|����1���Ν��xmϬ���;>̊O�Wl����D4�̖�������J���q�6��i��Rs�1�)�&���Ѯa��<LI�y�3���Ag��,�I��y�[�|&:E�L���wo��\�Cԃ��}戻Ld�Nv�4Ͳ\��;n�q
��~��3 R~B�f�(x��M!��M٤8����*N'S��+a�	��Q� #;�S�qA���������o��k�͡�b��c���3�m��y��mR
���y��&!X��):�&:d�}�I��aSo_��'�<B�m�|�bbLg�뤃ˌ�D��z�@�LB����/����>����������R|��5�'�b�~�>gϩ:����k$Yԟ8�Û�S�z�Y��������Ă�>�"�LC�l��"��'�{���'���>�����_��%��<]�g���7���d�P�i ��a���*�D�'��%OǛ��?2bb���d4��W���a���d��'_�ԂΜ�u'��n1g���I��-Ck����6_no�U\��z�Y.�
��=O�<M$���Vu1�'�?|��������ă�i1"�?2bf`q+?2\���g�8�ed���|��=��ԝgP� A��������ˠ�=\��� �,���x�R|�&~����x�����4��_)6�3�c1�~��4�Y�?3)�q
��1'�*O٬r��bc���fT!|�n�{�� �n��Wu	����&!P��ɴĘ��dR�l�&���<@�Q=7܇��d�=�v���i���Su��M�_u`i�I��y��>O6�'SL4�
��}��f��k��ړ3��y���(��~Ce���,���s�%zɉ��N�&���3��g��=H*�d�������>g��<Vm��jߓI�&�g�K�N!�11SYdě@G��hS��g�Ef���N-+�E*(U�	�5b��vS���Y:ㅙ��9y[�N������֝�uw^S��h�r�����b���a��5�[���՞B�B��k{�$���/��9W)���;n�F�l32�}���|z�'H]��]�ZC\��q�>[ۻ��n~��|χ�R+��ɤ���q�V�N1g߹�I�AI�_���d�`zwX��Xbq'���� i�N���~�uR
g��/�>Co�*E��&"By���]��f��o�w��~�����0����2��"�g�hy��N?$�'�}�O[�4�T�o�jN �§m'��)�H��D��}�2��ٮD+�Ϟs\Ǻ����!�;-�?!P��L���Ǩy�i�XV�ݲbLB�����6�û�!����������%@�_N������ȏ�k�@���Ϡ�E��3o�o>�������Lf�I�w�����ğ�x����Agc�1&堠(���+��E�<�ǉ<~d��=����l��O���'��d�C�;�򘍘�&�Nx���i~�t�"��J�̕��g���'�3��I���;;��i&!_��4��!Y�~���Y1�i�t�VKi8�RӬ� ��)�P�2\�~���m�#�=����c^���%�����˭��n��H,�?0��������'�qd�Y��T���&s��'���r����ORm
ʞ�l5���159M&�1�Rm}�O4�ǎ3��a�'��ȏL���������]������Ɍ6°;��q>LC���w�4�!�b���bbAg�;���f����4�hT�B����ԝC�-��?%aS��4��dĘ��������A�s�s|��yWq���c/���;*H;����?2T&��C'YY�J�}�qݓ�c=�y&�q�8����A�R�I{��f��y�u=a���=�p�@QC���s3�G���1����1)T�����K������e�9a�[�$|���9I��|5�d�Y����~�q<N�|�=K��I�+��g7�R
N!_M���T�g�3���']L\���l����L����^�]�}s򟥴��w{�3�%H/���C�i��>��:��l<��i �����!��S�1���1�����
�z�a�����Y�%��'����}}I����3a�H6B��Pj�ά|���Ҫ��GK���c:�a������j����,g���y*X����I�^̘�&U��ϛ�s��ݹ��l]V60���֥�hpZ��9�⸝6��sz��E-SdmE��K�1Ԯ{[����\�U}�F�{y�v�
��;H�G��
!y��<����g���|;�0Y�%Cɺx���4«?PĜLLC�%��!Y�:�OfS�>O8韙�u�C.��a�'�_<��n�ly�����J�K���V�7��	��ELz�S'�J���Z�N�2bLON�
�ɴ�O��z��/��,?'�����t�42c+=a���I�.Y?3əq����N��ԅg�w^�z�����׽��lVh��x�3�"��P}�È��O�@�dQCϷ��� ��ٮkS�q�Lzɉ��B��,��zw�CԂ�����Cϩ6� {h�OY1Y������O\g�w������7���n����>I�+�-4�V����ӶO?R�<ì�['���k	�u��N>��5u����f�s�1�d�O�w �N���5�m*Ag��>��OS�8�$��?7���������{{�bJ��c;l��*E�u<2�HJ�XxZf���u
�<��5�X<��8��Y8�)?}��x�Y*��,VJ￲:�0�
���I8�LCl����^y��뺚��ۻ{��T������|!I�>LH)�v���gP��l1XT*O�b�yI�2��i�Y��&ݲcO3<B�ݓ7�<I� ��I��+7�x�����������ߵ�^�aSC'Y�;��$�.�'��z�'Y�0��!Y��a�ͦ2xn�gbcx�&]$dQE:�C,=��3�c�Oǻ�G���&N��|�O���j�:�Գ����I#�l����{�����k)�LV|ÿSH�:���}��x�HW�{�'��Rs����LL݁��Y-�u�i<5@�q��-8�:�U&o/�����u�����7���)=�g����4B��m�'|�tN'��Os]�16���gu���I]����D5�*E�xw�u'�J���v������I�r�f�.Z�]�1+&���=ַ���/]}�o�>�$����ޔ,�h�X,�?[�8�La�]��I�m19��O7HVmӞwS�:�S�2~C�i�g��;�J���{z���?'ݧ���L@�_گ��C�V�ŋ�8g�Fm�����{l�����J���3t1yo5A��n�2=	�v>ʵKtuJ��22��Ƃ~(c���f�����i�&���[^KY�JA�y4�z��N�����ƶ�Y��jR��\)��M�X���QnV��������*��D��?x#�dA��A�3HbA^Xai�i&!P5�go6�g�����ON����&$��Ngw���R~g��޽I�/)
����N>��u1���B���0ǋ����w�odS����u��G�Y������<H:����3��c��f�I�퇲�[���$��a�%�&��y�&�M�b��{��<@�T�'w���Ru
�I�b�:w\�ߺ�:f�o����>���2i�d�ɷ��3*Ag�Ki�P��c%T5�I̡��-��B����0�O��Ag��a�|��c���gRW�&��R(T����ه~�ʼ�㺍�,�̀����}��2bOO��ed������T�����3!�3�J�����*ݚI���Aj��O��S�I�<�~���@��޷��ޚ1w(���^���9�{O��Ϡ�����!�a���g�i ���wA�z�Ɉ���0�*u�&>��!� ��<�0?'�=B����r�ɤ�?$�*�ģ&�R��bN!wC{y�v��ER���E̻�~��$�G���C�D{�/�C��|��M�����ox�����y�,�g�"�8b�|'>]��PG:�x\!# ��	��n��oq�Kou��ɭ�E�֥���ĹSo�����3b��b��nh���Hs��4y{o�nP����5��/�%�\>��75j���͑���Z���:��Ľ����L���QŬo�?k�fZ�5�X�=Ҋ�£��xV����؁4�j���L�;�<��E;��~�
�z<4���v�t�p�;�/�5�wԺ߀V2�t�����ڬ{�樬Kx�"}��r��Det�{�
�Zʏ�u:nT�ĝh�[Z�̇r��}\Z�wf�mI��6��	�����{jk�0�M���O^�p�cqɼ�`~-���9������o6�pT�ۄ��RH�mn��G�UG�d����bH�����T�{��*��hT>�v���)<RW���`�±Ee��ݓ�c��"��֖����Z�_oS��&�&�����ÕXV �7)�c��=+������$�~I��F�{}}3�X��ɦt��c�叡b�mz�b��MQN�A��q��s�f��y�����-Wt��\��Nö��7����!t�&	⑕{���&�}΄j�c��(q�E��J����*�ۃ�g_���kU��_�
m��wb3���"�Ks��v�D���+��B�E.�cl�@��Z'[��U�/������3�w���d^�-�қ0�8tq�}��)�����!�ރ^m7;0^վM��{;j��F�|�������k�4�7�Ns��#P����"J��Ոu=d��m�}�����d��^V�Y��H����U�^8�Ji�c��Dc��-}�����YEq��h_���Pp�BĽ��i�.��^ذ3��C��^4De0�^��o�m�tj{���X�6ۥ3��}=��������%'�NS�,H)�X��}/��ZJuvk$�ݦ�+�a�;�'���}0j\��]5�����S3�c�᧴<�U3�i��ɝM:���ʔ֨ ���obe���}_ �y��8�'�k�ʳG��)^-K2�y�C\��{��&� #���mK�h�kNɕ��er����*wC��?��B��s6������Ε��]�K�.��IH6���*��iv��ӓS3���Yy�]�og�<]�eҩ�e��c��X`��j
�����ĵܣ��F 3S��)����i�
u�x�5y�Z'ת����i�~t^�&���B%�:�j�� �A�SBjw�ȉ�l��Z�U������A
�[C������\�}�`��(�)�\"��L�9 �b�PAE���h�s�3.�c�ȼ4����tňM��-¡,�F$�*�y��f���
8�n�ed�A�HN�-ޘ4�6C:խj^޼��S��g%K9*���@��O��P:&�	_�$��bU�e؋ՅSy�I��q7IlV_E3g!����맀P��qb�D.���O/3���+�]]+cG,��f����S�j��F�����ƭS��s��`8�!�n2l�m֓N,��'��-w~�2�nn4�Y�I͜)��V:�7m�7� (��G�D��U�Om԰�.צ�V�>ś�6�c�,�g�;�0)х%�j���t�ʬ�IQ$�9I���D�)����N�.��q�����#�dG����y�ף��"#N�I[�w�V	��VD��ma�a�C�.C�	�4���[I�)�dtW$swj퍴s�T<�r�rxn��3�l1Ur'od�%��/Z�p���}Δ.he�n'N�^�gi�"�al�}�0��/���4�tu��Y��lhᓥ��Jwu2u�CY�j�8/�̜ɞ�q1h߼��<���Wk�,����dY�0Γ�zmFE�T7X��.�����E��2ȡm�j:�+hA��� ֎MU�s��r:}��E+������3Y����P8�cv9�̭�QE�O���|�Wjvj,�h��(��o�t!U���o;�m��9F�C����c" �
���:'�ia�|��}^�.����l��.m-������#}e��X%����0O��X��X�Ά]9���0�l[� f3y���o���.��ZjŃ�AR:+��+O�!gA彉�����̣�]?joH��V��|x���()�Ӝ#@j?w�1p����c�dlTXq?bݶ83���]�4M�M��)]P;�������.�XZ�V����Sw�B�㜓3��d�3m����R�`��!q86.2�JvV)��G�l��G��z�5����Õf䫌mn-���8���]ʺ������x��r�*�~�� 	�f�|�֛�����מ2=����ϓZ%�FUy���k��H�{��fa�+���*7t,NV��.���y(�Tl����A.� z'�<U�3}���]i�m�j�qt)���	���x��MdQMn��g-0�"6|��j9F�(���i7����Ы]�ӂ�S�5\g�F(渋 ��RfΝ��M�~*�+ Y�ۑ�"i��*sI�ڵ5����p���:���HΉ�s�xn�.YgCG�a�l�!L��%5�=)�� =' _W��:N�\��J���6Б�3Qڄ׳g����NQ"F(�T�޹��RT/;̞K�L�}(�&9���K$�Rw"Dv�b���S��gb�R�Fl��Mm7pf���|�jZd�d7�N�,�!����{�HWw�Y��'N�<ܶ�v,;}ȇ��h$:!*����);��@r,!��tl:�ؔtk�h4b�|�ļ������u{����^mv%�1sO׵��]�؋kq̅��c���ڒ�I�UO� ��.�ډ�6��ꂑ�q��3�ӽ���7��ѥ�7����&4a���Y,65Չy��NT�V��7NQm6��&�%��\6�j �S[oMe��t)���oh��H�	���s�/"��~ζeʓn#/,��Lޏ�U�}C�!��})�ˌW-8���A��n,�W���WB�x����r�2/�b�ݜ�Z�%ٚ�H(�xl��J��XX�����$�����W�𺶮o�
�8��oV����y
l1z�I�=:J�1}.��:�4'�Ҹ��,���huB� ��W2��\�h��/��^q�������:�Ζv�>��hF�p�#�7Eu��a��=�x��v�:��`�Lb
�#�Ψu��^+8C=u�9�P�Y�s�h�! j���Y��S����70P��n�\�5; �'�I��oS�~}	����ˇ�!N�,z'��v��2)�*��K0�`��Wr���j�"�ɝ����C���]3��^��ά/�w�s�~^�EGA��@��(�Z�/A��$v9ӆ×�����C1˛ֳa,y�u��Y >w���!C��(w:I���f�U�:�&5��7sI��R�������hdQicnp�v�A���ܥd#;'�=K��7;�ߨ���-�i��.����˻bc��2�T��AbDА��̠�b�X����1�g�H HD�I{pl&,7g�ڟJ3=g��ݗ:�vr�1gr�{o��9K;��#A�Tb�&�%e�e[��z_��6Uɹ��%��$ɡ�mX\��r���x{�fs�<��«�]}���3�d]oHiH�ҝ��d�5�B�莅68���P��i�/.���-�]����Ⱥ�c�g�i�	3�d&�M����ܓ��S'H��dh�*��݋��7�:�r�+��pȐx�������-�3X��Q��[S�"69���t�G1��Zȁ3{2�����2r���mn(��'pP;B{<��f};Ӊ
�Ŝ�E���\�fL9"�GB���͗�Ҝk}�����P���诼���;U�7D���5� ȑvO�V�=����:KQX�e�I�\�l7e��������ZB��2e]�}����01'R�g�?c6Լ�o���c�s�"< O},�QWq7�/�j��pT�(%dZ�:e�g@X��{Hc���]���ʮ�Ի7#Z�#"�D43��J�r�h?��޾�AK_�W^��;&n�D�[8�{s����Ǆ��b:	h�M/EWR�L!"�Ϻ�8��-u-�5�-׷�����ri{��R��|(��Aˢ�
�Ҏx��g��T������A��=_R5��y�j�K�;2,[o����U��װ��F�\���0��ɳ�+�؄V�&�)��5�켻%���ϲ�ٵ:#�����T3���u��;�l���"�M���U�k��ކN�*���2�WN�����!*X5�',{Zn�=Ӣ�H�p(�oVZ�!5H�GS��c���ttç�Ь;���u������pZ�ʒnVp4 c����]�2�P�� ��r�h�(��y��e�M�3�v{�â�I5��ew\�n�h��)�Z��(�8�9p�]alR�i��n�5�M������tѢhPK�{9�B2q�����}B���*�<��k����;rE�hS[�%9ղ�x�NLR�5J����t�F�Yb�U�ڲ�|�]N@,R����7�un⭕(t ���k�Pruh��c͛:��FI&���� �֍�jf��v�W��:�9A�-U�2�f���X����t��xJ�}�#W�mU��E�N���Tw�
�8��c�\�<�h�*>��*�|��9�ggP��en��ו5�%N��x87q���@�+1��jF���R��Vi���#�a��RճKXZ��pEî���r��&d�L_9�ft��t�o�+�NuA��U���#\u7���']fe�X԰�n3`��Pp�:�S˷�o�|��G{p��9��C�(��T��fK�7HN5�m��9W� Yx�7���w�>�i=S�[Η�X�E�(��qRpР��^7`�q�ȭ5c����p�B��]2������cJ��D� ��X��:���d�h�ߕ��xi�f�E�3�[0�fl,�N��w]IQWM�#�=�����FU��%���q��*�q�̲���F���:I7;�4��P�2�VE�q��Ա��Xc�<,ԫ����8LylS�sq'S/�X��5"�8M��\�{�<��6Ĩ���n���.��jp��4��$U��g�M�=�S�u��\R�H\e\�)�,t�L�]GAw@=�f݉����#�o�����8yM����	{���_RU���Ƚ���:k�-����mK�ٹ֌��&	��[���z�#Λ�|B�j�$��ق���\�hY�K:��(p��ۏ�`�w��1'k$r���kE�h-��и����$��ط��_b��We���7't��Y�X7.�y�5J�f䩋�Y�3o������kCxaH���ƻ�ۑ��%�'ov.��9V;��A��Ds�ӻ��_k6�K�ҧ�=n����\�@l�Z������>�����dƃ��B��2Vu���� �X�����[�XP�]�J �=�z6◭l:��*�����ٲe8��R�T���يR����'B�ۆ�t�MM�*<�'n������^�	���*3y�śßm3��G������7n�m��нL"��;��q��6k�c�p[�C#G� ��U��eUH��*,D-���Z��=J��
%�-R�(V�Z���[B�"�*�EF
�[)V(�m+Rb��������Z��E,E�ƕUbȨ�cTLF�X0Ġ�h�+D�҈���B�J�)eQVE���(����b*��YE�*�Trܰ��@F*�*�jҔUKh��
��%R*�b�ZEcaYUKh�E��X���LU[k�\�`"(���k*)6�T�L�@X�*�QmƸ��T�V
���V�,QX(��F $EF*�b�j�UC���b"�����K��)X�EW��LG-`��B�s1AALB��QDTbV���ҍjG)b�
*e�&,1��AH啈�UG������^_����w]]�6++�lUQ|���t����tz�ruל13��rJG�n�}*�3���J���E^�����{ﺛ�PH<���r��
/����t��ڎ&<V�F@YuP}R��L1wͷ��ծL!ӵ*_.��k44uF��_H��\��=���������Pц'h�VJ���9_t���ȥN��m��^�~�Dk�|�� q�T<>���ϳ�y�ר�4�8�H��_^�ڧ���=ɥd6��M�ۜ'\Y�U@"k�ʱs8Fޥ��=�- J�2'Ѱ�a���c�._m8T�A�s�:�`=B�g3^SvT	]SćZuZE�R�D�&�À��n�4�d"�K�Ⱥp�x(\��I�l;P^���i��ʓZиصOE e i���j�v�@g/B�&���/_T�C@�Z�x��Ө)�'�{�x���%)�ϧ�>�il�nm�^�7FE�S֩�BFqa�r%�K����Jm3C\�"�����C4V&Ѓ~٩�.4 6�d�0w\-�5R����7)nݵ[���E���j�̭�l��&��A�Yp;"?>�8��N\r4G��T��ɉ���<�9܏vg1:��<�r.}*�g)����ԇV�$i�{ܰ��3D��v��^��'5al��Y���Z�ٽfX���zl�w�l:�ƛ[U�ۢu��F��it��2.�֙�hv���M�-/y��͎5w�P4j�V�6��qg��xx�}ϼ�vsk�>Pk��x]U��'���OZ�{����8����.��ķ3��=~=:���k�"0Ɩ�D��Dt�4����Ȏ'��$2'�9�U�s�'�=]K6#)[�♞���}�E^�K¤ep�@�<.�^��{19��qω�����4����\�$�q�uc�K�Qz��ۘ�B�$d/s&u�����EJ�GT��M���~�U<F0sz��z`q�%���y�R�M�Z0�x�̯���5�K�OEu������=��87�g��̀FE�p�O|�CB.և�0r�g�%��K؄<�+��c��g��l�=T1V
u��z�h櫞}B+��U��;�ۄF�zy�y_��W7�gf�'��^�D9���(�>����,��S�͝;~�t�
������\�v`ںw��5^�ɜ�3�+R.PB������bMN�r��e��Տ����%�Lk�����UVV�gn�������<:zDH�C^hH��M����|=����b�Ct�x���ˠr3��46��>'�H�C5�"M�z���﷫�VT]J�6w��tXq�C�4�{2c���z��b[?��U�<>�k=������_��r�V�n��+���8��1��yٟc�ʁ�������xxx[������2�ڶW��4�5�w(�&9�DF�K$;H��ʥ��2��:[��i�����ܘS��B��E�9MU�Z�e�ɴ��M�񍆖�+݋G�f�C��������@�vz�*�3>���حu']�����l!������[��X�-��w�*��h��G�f.X��9��}�)�i�D4�Li�����_0������K:�V�No^�ւ̉��}��,ޟR�5Õ��V���Q�Jd�5��:w`�׌m;Z�9����h�/}Ы�~�S�*kK�®�!@� ������F:	f��fnܼS���%d�k75�2�"򖊚�7��v�;O�٦���ىC,���+��Ώ���!�9��o},��S9������Ft[ܷ)��+����إ����p���L�G���[���귪�f$s3|�!x�4jE�U�u��`��}p��չ;[}'"Fy�����β�f_QI[�d��!�MpN�n�q��z��k܏� ��c���I�~�嘩�)�K�O�R��
��U�S�V�86�����k0��=h����4y��B�uC�K5T�*�.F�Sb����:G�x�Dm�G�?ɵ=���,=�I;�7�;B�7zR���d�d��gm�'QH�%�CJU�c�g5�U}_W�}���]JO��U�|�'L�#V��;��Uk-��0��OC\� T����E����;ρ�'V�`,k� 8����#B'vB�PČ��}���q����Mc�scu�R�ݒi"�gφ��,s�ԩ���^�*�=�bAo�(̩~kp]@�|y�ף�Ib
�����}<yÞHPhYiHm��Ȍ&����ad#*!���c���9�t���3:�r��}:�j�Ƽ�ҝ�,���&<:g�F�K�ؽ��+�/swrm]��{>ʡ��r�c8�#!&s�����I�Cw2^�2l��t��D�;���ǭ�LT\�<*P��#���~}���k��V��Dls��
��v��#���*�v:
����T9<Qj�v@�`Y�������९�X�s��'�Ҹ-a5Ow���=A��'P�q�-՚4:�T/�<Nc�+�P��KU�6O�49�q��:V��tЩ�zMØa֡F��xR��m�~�����ev�C���`��{��#�b	B����;Hut'
��Ԇ���+u�ɃΔ�IY�BWLj�"�		v�R������H �z��f�;�Y�Ѻ�x�t0����w�o{S�9٠Vv���b��1M��.�f�ɰk�Y ])�������Z��op� �����i��h�~Q�u�G�Us��j*�'��b���\��2�a�gom�xp�-=.(�\Í����\2!��
e�>��{��̬���k!Lm.Yc8�h�k�q�a֥��D�TO	D��SK�UԾajw���nC,,����j,뤢­�L[���3s�����R%�+
�k�28�Fεu�+�	�T���>��[���I*;' ����:���rתe\}Ϩ=�ק�Hӥ���Q��+u# uA#!��b+;�E,���Ǜ���"����f�<��[�V����Z�q�\������;���襒<.�˦�F��Y5�u������"��k�ܽY�7:u*yqb�D.���O!�7F��zqO];�����U�?*seP7������q��qCjÌ�*���gl�q�N���m�ۼkh[��A,���-�	Gr�(F�jØv9��!o�\&��8�8�i<F����H�J��0.6��tG!����E�^trlȎ��5�q�ִv�E�OT­��9�K>��r���(���:؆��盼5��Y����2v}��^Y��i��(��{J�i��߰�����++�eGΖ�Q�ʛR�ah��c��[B��z��{,J��"�+��ꂹ��C*�t��}�\v��&#o�v��&c,WF�U;�x  ��n�rxy�C,`�NeS��5�^{F/����(h��k�}/XXx�8��8�p/�f
�\�J��Ng�Z+2�!�2ꭺd�:�Ϥc����-�n�^M],ٌE�ۺ�6V{x2��|[��t��׶�M�i��"�/����2U�Ѓ�f�?��8���E`�zq��7�ێr�uBȣw�گ��f�/�O���w�eX�6C�,���R��|�+{���� DͿ*:K
�g�� G�_Pw�4����,���L���'�1��=������[5��܌1���%�t��pY|Ǣ�Ը�U�[�r�Ð�����qTR�ӔLb���6�W�7�1��� �F�jJ�\jbѬ|o�k*��/ݚ�k|�{�,�K�7DZ*q�ur���d4�5Ŋ���2�s$˸�Y��x��M����:}�F�Q`��҇��Qy^n����kD�L9�<I�E}My�k��x�`v�F{tAv+�+7p1ap�OКA��W�l���}�T���D^e<wyB2���N��_r�M&�,���*�g+�1ss�Ц>��-
����z�F�\�w[�3���~�G��j��9��]'��r��:Nۛݙ��aC�⵿8�s�J�;WV��=�d]K����e�����Z�޶�b��Ɋ�[Y6v7���xxz�f�y����ꡪ�����]g;
�s�P)�F:�rxl7B`�=yS�i��院�a��u�`���D>�s�r�����,��RfΝ��M�`�����W����bپ�Z0ݚwQ�Vo��|P�OG�D*Fz&�^/K���D��tWk��,�)-U4��y�5`m��ǇG@�+�XHcf&�5�߰�΂�^���^��}"^��w8�q���H�Ml�O�t���5�xȬ�������
�z�q���5��f��賦���ǹeKx�U�G���o��jZd�g��'�Y4hk�S �N���-]Go"�ô�������o�d_S!����ճ!'��~����\6>���V���8������;��
�PxmY��_�[�L9�4��8��B��_0����Ⅽ��sѳ��
�ba�ER�b��C�T"���g렴��5p��t��=HV�0r��r���W��d3���߷�xӬr�`��<*To�;P垭�� �EQ*z�;NJ�BK�/�<n3�7�4�ms�Ֆh*�؍HݑP�s`���3�Y^^��J��\%BA�iowr��2P���]�'s�4Ǭf"�H7A޼N��nC՜k�;����#��:<idr�#n����π����k3{�)�a�S>���T�[O>��v�;���x'�d��3,�W�5 tM(]z'(�ԍ	۽Z;J�@l�-����C��N�6��+��ף�e)*�v�mq'+�׷��m'("Q�tH���</��B�dv�u��0�z���A�},툹é���w��p���81��S)'"#	�%�3���=�LH�OU����0�l�cs�n��γ�A�I�X�U��D�.&�֢��;����8Չn|��:l�\+&�.dٞd�s��$�(?���dc�P�Pa�N�D�;8F���фl�}wY[�;V���[S�''�����{a�$*��B5W�5��-$�1��6Wi��D�9�`�y��֨�qGTb�p�����ZM��qۡMA���@+*�-�+�=)r�KR�� ���!��+>rʚ��*�m�2��� ���X%ȣH3.�cs<����oh��kk��ĉhX��OV�І��<i��9�|��x�0(cn�K{7G�P����m�!(K�o7�c�;������C����N�2S.��EgR�?lYмERߚ("r��ʖ��&N�R�V&3�2ެ"�8�ܝVP�Xɗ���/*�BwbôAŚ�ї��(h'ZL�Ĺ��-#��Y_��k\���� q���óh-��L���i�uF-c��Ga�R���6:�pF��w�<�"U��D���f�=�l���P3���tz�i�5���X9�k�p:s��W��zǻ's*�H{��2���s��+gc~�n�[�|v�ѓc��-a��pU�B`<Yu4�V:%u���oX�̕��7i�de��N/�s���s�Ϥ���&L*��E�`������k��R��.U�R����Dx ����]ĸU���������9k�B4�y�q�.�ֳ1�rx��t_º��Z�C>� >T2!��S-)}�ܧ^g������ڕ[��X�qE,S��ƅd$�$�O�F�1`W��L!"�Ϻ��.C,,ר�����j�l�ծ��[�����=�Z�����L�e(�\�x��LKi�F�Hw����Λ�>y��� ���mE��� U�1�\�	MHYmL��|R�_nַ�ԯ{����&H������>�|����m8U��OH�)r�|�8
����/��)FgH8_q�M��{~����k��+2Ƣj�m�r����[��	R�2�[�]Vc�cz����+���2�.�Ek�-����8�i���.���cw�G��u���'�]����P�̤����:��V�gz�IN���DG�}�ܐc^����H{���f���.��qr�f玥O #��3�>H�kqTO�[5�u�s޽�y>��:�,� �e�@�=]�cת�T{;��t'�6��2l��n���[,ԅ/�ml�wD)I*��U�(����lv�9��sU�Z���.�HfPnF}/���m?s$�f� �zH�BC]�3����m�ػ\"ܽngB��5�j���irЇy`�؈���X���BS�\��^��N���e_/a��}�_xڒ��N�}41���/y�A�L�-�%)�����sH�`J�]�c����M��'���١�4��27o۴��6��>�d_8-F�d}^���
��uo`/�<ǽpr}����3���C���`Yh^�5�fܩ����F}�.~{�j7�&n�fwwΡ�ˌ��1�eZt�ˢ˯	��T&#Z\��m���(�L6��F,�^�k�íjXh���\3|˪l��F�K��	}��!���V2#��$2 z����aԒil�D�2u�Us��B(�{�mDt����xѸm�����
YK��oV.|4-�1�]S7B��Q�
&�T}KV�@0Eq�p����	e�*y1V���i)x*+�����p��59���]\��A�[���a�_wAe�H0�bڕcz
��C6wd�6��j���-=
�ǔ}Qmk����+��������LC�R�4�<�hu_X�����Ob~���.��;*S|��^Q����Ӗe/�J vu=̣0���e���cl���W`�����Տ�>��Vqr]J���2ucm�<kO5{.�o��Ӥ�^��K^gf�27����Fu�X]Gs����-�Z]2�Ք�t�U�S	T]ʙ�ֳb����m�w�M�N��Lԓ\/6�BM�dn�1�\\ Ii��[@�-�GC�+�v��;ձ֠]��J�޺6���i�����n�hu��ou�l+z��j��Yb�Bz�/�Ƥq��*��Dk4s�gVf�E��Q8��GYXEU�+��b;qQг�9��n�p�R��=�I���Ɖ�7$��TW��L��%*WJ����!: �R,V����5;�����|kyWM��au�7}�A)_��e���o�0��]�R#c�廙�fAE�����;\TS�7a��0��`(F
�^`<v-�4�2���Z@ox[�=�X}�� ɇ#���Ŏ��ok,�_t�n=J<j�}ھ뚛\�J��pa��r����Og�+;Mp�f y!]����#$�tq�g%�Ɍ�2v�P��ww�l��4���s�u������~ܫd${hk�u��ץ�%��W@��e�z�r�9�bl���i1��bn�v�ȼ�XQ��0`��51ǆ�v�è��^e<rG����M���.�)[7B�q�9�������Y�;E<
���͡M��9x��i��ӯ Ý�CtS���Y�ϝ�]p��]w؜�+�Tn�\�"�ãS�ͣ�4�O�P��۶�.Mc�g�H<u)����p�@n�o@lv:�򦎠6�A�2�ݕ���ir��a�v�����)��73q���ړ���b��y�u�5kq����]�,�~�҆���$�U]����Tޫ{���y�&��d\�[*j� �����B(��ZǊ�k �%Cݪ�IE��Ź�)�gr�)��̹�{H��LS;�c�*�[�-�c�x���
�����ԅ�': ���p���+����3f¦�w��5D;r�hc3"�u��3���4��ˊbV\0��k3����H��V�OOp��#K{o�/I���m���ctr�}d_N��3li�ݥ��w�Wu�R]�WT=�WN�vttqD���B͔;�+����cw��T)���EY܌������c�S��Ӓ:�i�g���u�(H�D�P��j+>��Z��[[-��R6�Ĭ�,DJ(��q�2��"���`bE�*,b����A�1��+YR(��EZ��`�UR��c�+�(��,E�TUE$Y2�@Rc**���-J1V#"�`�E"
&RT�q11(�*��F�TX�*cF(���2��UJ2UZ,PY.S,8��cLkDTE ���*ň����*ŕ(��ʂ���TF��e�i(�(8�@�2")���EUR)�#K (��T���`+j��9h(�&Z��"31bȵ%�T��Q,�m(��a�J�[+$�*(����0H^D"^��tv#9[�nr�n؛���o������:���[�ye)����b��B� ]���S�oZ��6B�gGvQs�_}U�W�_F���:NE�+�����/(u��+���5%F.4&!�"3�����7-ҭ�,f�Ln�*	��\-�ja���~p{����Lk�՚�Q��QQ����n�z�rY�̔���C�?������z`q�y(����EF����.�����b͕V ��l�ǝ�>Ǳ����ڠ��ؽ���v��&�<�^��[U\O��{mUnaUu���t|��I*~�$�����p!ܺ���j���"����C� 3��7��D^��m��y�\�1��ҟ� E)DC.d*]������X8l.��	�ͱ`��#1UP�<7u�G�0�wKn�����#��5�:�T��L]9�3����0na)��7x�\;�3��EU�/�Rj�F�\�x_�zDN��Y�5P^M'�Ѕ�re�e�JIE��%�vx�{ԋ,�/`}��v�N��E��"#W%�
�ؚ�D���"��=���uݖ�8�9�����2�#��3c�MB�i�Ym2m=�h���UM���bZ�j8�I��>��{s�J�Kz:�C�},���8w��F`]�p��V�^_1��=���~O${ǲV�����S�;[9 ����:�Gs�h��yt͈�P�oFk%���Qs�i�ٱ�!��:Hi��\ö�rM����������������<0�H��:.{m_p��B�*����
�����y�}P��R�ɖ����_.���Yx�9�FD��5�Zk�X��?���o�0䋼r>Cʽ���M͍o��*���RW3� �Cy�u���|i����jY�_|"���g뉢����9�+�[��D�)\�Q�╜�1��X;�I%�!�ͺ�|h�TUpT+��n��h�hR]���H��ٝ��S7��
�i<�C��Rϖ��3-S���t��x?fV�j���Ծ���O�x-/籁�ʅ��}ȇاr�~~���ʦ�C+�����;z�Ų�;� �↑p)_�� �N!��R/��u�r�Xg���Ш},���1�W�it�`�Y�
�iW��N�J]vSK�x]8�qt;��\"���Pa�t��=2�%&��8���ג�\���"Y��&��)!�j��6ۿ��t�u@�	�]�L����ԩӪ��c�u
GO���:;����H�Z�-��q^/
�cu��7�&|�����˘��ӳ&]*f�ǐs6>�����OFh�ҋU���3:&]뛱�>��OT�K�o��{A�V��O�Rᇱk�pǄ�A	�Y�8t'�4��Wh�!aʔ�fwm+��L!u�%����}}��fgs���g�{�ڞ��mg��L�q���@�^��Q�D�W�
�Ԝ��[�^���{\]����+XΠ���s��aÞHSB�J[s��v�D����竵��ʫ�b����aК�6�dY��͈+>sl�"���Rs�;�jY'MB��Y�f݃����9.����~@����G�{7�]Ac�dq�FBL����b��Gv�D^�E��3��������F�p-%`r؟+�"|Y��m�_��)�oT.�nB1mѡ�,����ck��^ԝ8`���)P��E� ��r���=4Up(����YJ;��i��U�k����s��u��u��P����:+�*�d5���כx����X;	Q®���g/�3@�:�+a;,FW=�c���o.�@n�$�uv�o����Dba>�H��fTF���3����!��8���{�N�^/l�-T�\'Ƶd��ky�n֍ ��~��uT\����R��S-'˚y�S�3�=�a[~�Kj�k#�!��+��%k��ym얫()P�9�����[]ڕ:&�(�"5nT"\S�z�,���Ӽ�n���H�:g���bG�; ���J⥻�-hy.��TsWL��it��Ĵ���ШZF^\�����;�2���=Bq}���V\�y8
C��4Ƚ����d$�%��Xz{F�I�/�{��cH'Ճ<^���m�<C��#�\$�[�m!X��U�zY*8�Yj#gX1`���V��[���7Β��������<n��O��mE��2F���[*8� �ԉݦ����e^���]k=O-ъu���ut}_��@©ll���a9�}���̻��"�3�K�G�>���2/�Њr�i������I��9�1���2��=KޜΆ��|��Y CHh��s�c�!ꉯ���7�N�
WL66u�E���l�����}�o&qlϾU���&CtZ��
��:�C�v�]�p F�4q�4p��2�6�x�pU�u+D�e�E�M��s��P"��Z�<k���w:�]��N��Ѱ%���E��y)<'4Ic��p�x(bur�c�M�\��^�\��;dY��7 I�z��ӌ�b��_���}ַ�T��q�2R�qg�� ��il�v���3������wU=�+������E{A��{K���o�+�'��"[��D-Ժ~��h�E_f!6�T���i�ێ�e��9�SF�L����P�}�q	C�;t�Y����HV�:�9v�(�&n��.��I��N�h�FZ3�f2V�e��=�{����ˬ�̵���E�#��7i�6b�8L�+��KQ�!�+��Iؘ�+1yt;k>�����p�A��H�=r��٨*	��љ[L؅�U���|�k�fJ끊��m�q��'c��D>:5>'����ee��
 �uTE}Z�{J�0��,B��]f�WnZ�0�����:�{Чf�:�GZ\1�����8/�j�ުS+�Ze�:�v뵝W���2�#&4PR6ݦ����P��+�����q��
��-SM7��H�4�pka^J�u���tft���K�
/P�ۘ�^�	}�d��ȡ�Y��ߏ�^���~���* �]y	�#���6���o!x�y��uZ�?6�T��==�g�������0x k��+Z��A5^�ؽˡ�|�X��!��*�.1${m$�,GN�穕)\��q>�Ƀ���Z��H6�ȩ�_��dc�N�="��z���~)�$�(�c^d/�w?���<*P᰾���I�\9�mU)ȡp�dJILX1�e���NeПH��i1mΕho,3#k%`�[#�D8g(:���׷�^�5[Pf�''J�6�.�c[�|�]�x�2���SK|���$a*Ęru[T���:��iw_N��ei�+�������g���� M��H�E� Yr#)̵GD.S�����}�za�E�[Ֆ�!��V[�ܧ��ң�5�z�^�<m��MX(�K���ư����<�&��L����#|?7q��`��QN�*��/֫��}��w桓��dǹ�D@�,32���Y"a��oL0���%eC��}��3��#��ה�>��֙%�n8�y=Lܭ��� ������	�F�W3��t^t�:�l�vw{5w�	�����R���E�jɐE�'��ц��eU�J��X��';i���3�9�U��Ö3s��Kz�Y<�I|�z��\+���wn 'S����s��n�TV�6��KOMT8<y�|&��>0��sӕc	S�qeK)d�����}[ϐts�r�5��48��l�R;؟ӣ�-� V_JW�M��֦ĲQӱ$�����%��n[��o��YL��3��u�t�YACI�m^D5k�Q�$w+���'�\E�f�IQ"�!�j�j�C(�p�<��7���T�%��^���:pݻG(N���7ݥ�&.fN�펳��`��X�z��������������%l&8J:�T��X5��J\͓���ﾪ��� �Ӈ[T��ˠ�IyA��P�V������ɓVg�!���^Y�����d��NG�^�]Χd��.O�+��vPk7W)�s�f�q�r���]6�Dܓ�;�P>�X�	,�W��
���Z�h#�Z�i�����|�fs��5��"nU��J]:�)�s4o>(N;J7:˓�s:]4�����鷬u�b��P~K�n��e�GWf�T�R͖1�_�Z�핪�Q$�r̵[3��	�͑��v3�N8�����\��Y~�s�᠙���5����q��E��ٗ�8�����b��b��ҩj;�]z��*������KT{q5s��gu���	��q�Sf��+��.K�G�����S�э�W�v���]�����o?�452C{Ҥ�>�{)�w+G�ޜ�[a�l���:Sx��5� �^����z�5{�OYK�Z��W�Bvu��K;V�>������"���
����]�įm#e~S:�����M�L82�R&�pN>'9����y��V��1s��s����q�s���7㶷�l��DV5��T�x��#'�w|&M�7f*�o[ �:s^w*{}Ӕ������א�>�N9��rn7�MqA޽��w�q&���"~��{"q�GfO��f�^���.�����]�s�v�g`�mӱ7͜M���s��hf�*�l�\#ޭ�2��fÜ�u��4e;9��o���������D�7���j�p��J[j���z��]���R͈k[ݱ47�ݻ��k��7֠-N���D�]���eosQvg*Y2��i�����	��3�	e]^�9�ޝ�&�#�oaZ��_�:{�M�~���k>���}�1���P\ɠ�]d�=b�Q�r�F{v\O#�b�˺o��Or>k�:��zF ����U�	�e��)E-+������-d-�/��L�cY�l���8s|t���Iroc`�k��O֍��v�<P]�d�w`��[�i��r���@}���0���D�����I�A"goe�7�Lf����O5��ep��q�����>5obp7F�8V�^�i�ކ��n��y\gi�Wu�m�1Js	�)��"ˮ/X�ò����ن;��]	��	��ߢ[�i:o�뻈QK��������{�+��1;$���x%�(�l��� &hwz$�z��g)�/b�r�˯W_Q�ST�ܥd1�^!��NC�$��WX�X���m��G4�
�6��*�3b�i9	��!�\�IS�k]_��޶��������}�����ϭ�S�V�um����������%��OӔ�R<��+M�������ľ�Y6���k�ɶ�(U{Nh�WrtC2tu����q���qX��KgoJf�3ʇg��Oy���*�Rh���Z��>��o��ӻpTO�����1+t^8�v���MV)U����9�|oo�9�e}#�cviC9�&.r�!����oF�tn����i��s{��&o�GG�����^,~�jW���(�\�
��D�soe���*����B=v��ù�f?y������
Jm����[T�bV���"Y二>��IK1��}m	u��Cs+9ih9B^Tޠ9�ˬ^M�Ç&�.T�Bd��A��(B�82��`'��#��K�V����S퍳|�g]�}��6ͷ������&6���;4L^���A���G�
�"���G��Gm��T�tZV�'��}-nC�}m��3��As�����G��&_������	5/���*Oq�k�K�<���vUl��8�[�VbH����ˣ�5|�����ZOԙ�(U!'��-֞hj�.�:n��!�����2��%�Қ�+�e�����$�,%�9v�FwSW��5�[j��P9��� �H�[j��,�%W>�K��F�8��Uϟk�i�t�z�V �P5r� ���B�BQ�ov�r�bY��������8�l�w	��r����L���&�-w���b���)�;�Yr�E{�u���j�'m�3�vfө;���׳{��/}]������G�K�\V�g`��Շ�w�`��t,��l�cUR���1[o&uک��v���)܅��g{~�
'6Zr/y���w�Ӵh2�4:'�&LI��)1��S]�:�j�����ݹ��U��h�S����=�u��Vr�:ɒ�J��f66�!"��.挸<)c��#^Tn���W��.�'7��U�{N��;�G(���O82WVv]p=�4�8T
�qKPr�!v���X�M4��'f:;e���1J �c�cRW+��WRw��T�[��Xu��ʱQt|RZ;�w9�n�˫MR�ݴ�i��FS�D������*�ZVeb�5����j���w6�v%[��.�u}��{��K��-˗f��7�$]�S(��X�����qSL�#�M<Lv���h����ԛ�ed�n��R���<T�La�o00:���2�A��R�F����ޡf�Dv��qՉWf�Z�0��b<9-�r�K ��6YFsاD�%�!r��B�
Ru���c��9�.���� 86*s�$ϤW��)`��f�X�9�@Q�9�F�B���{���%��N�Ot�#�["8���e�I˺�8�*�U����\W�3,�5�-W�&ljl�ۤQj�	N,����k�K�P��×�}�x�Q���5jr>2�XQ
�9Y�[��w1V��8�ks��'��h[rp)P����+���ks��Ӳ����u�2���Ĳ�n�N���r_v�}��6��X��w�����xNI>���P��֔�Dk���Տh�=ṇ{��מ~w�1s����j��T���Za�*��6oI\֋�����*�1- �X+N�;��t��5���e�b�)v���s�g^63E��v�U�rIIf�T!��H��ki�&%8CQ�=z󴡤;glEA��{!�o6�sZ��O"�&�M��A�i���jD��Yѕ���8���� �tsvv��8	]�Ch���5�����a��l��olpְ�JN�,RkB}�a�}4�W�+��)���6-d�i5��u�<�M�A��D�&����hdM���O+�K�5��a`B۰�����˻v��<�x-"�Νb�M	��.'mKӖ!�І'�ɻa�s6���uJ0���.���+�^��	�����`��t�:�oE�:�upL���W&5��T�P��N���<4�4�L�L��l1-D�w�voX��gN���R=�s9����(@9��=��-���.�]u�0�6�o2ŝ;wn �M�xF:��;�ҿ騥�d�B>:33)b���{�J�v�&�Wr�Q*ʙ�o3�R��:��0;i�z
9��vx�*�]_R(�����7yt�)�o��L0��3���*sczQc��;s�o���m��W�Ge��y�5�S%GY�|��[�^�8]	̲\E���\�����Go��:em@9X�t�C�q�j����_S�ɼ��[z��qxJ�Iဌ�Y�T���uk6��X6�N�s��;��p���ß\֨z�uJ��j*�*,+TP��V��j(�Jnت"�Y1�AeaQDE��Cf[1��-���ł�D��@X)m�c-��TB�e�UU����FT�� ���(�FEYJWd�A�����K�LV�V���E�Ҳ�B�
������j@Y1�*\B�X�aXVŕY"�`���k%�QAJ�l�T��A��b�ԅJʓ�kKHUb�X�X����k�T�A�*Ub���-Xbm����a���Y-�UB[,��LJ2*��� �
V�m�V�R�4*��#�v�7t�W^�E�ty�f��yH��#����%@qA\7"Ѕ���]�8Pu_(te7��i�X���*W԰�X�{W菾����祥s�yt;�6�>��N[��;��w>\����V��p*�������e�gu�Sn	qz˔R�6ﻞ��J�ۀ���C�_L�r�WK][n�m�5��F��2)&�"�g"������tv͝�(����
Ry#��;N���?�;!�Wrcȝnn&�b�k"�f�U��Oث^b)�K�t��p���0����R�g�܇�֢�=.�Z�'�j��l��w;|oc�1��Q�zsG��N1�IX��n�Ia��������fv��GV����φ%srj��Ib�H�Tƀ��5e���Jv��J3�k<�s�!�%sr��ЇL�[�&��mC^����	{I\�c��|����d��:�t�B��I�3SW��WISiώ9rW\�핪���I�2����o�	m؜�B�3�:��c,lR`g\Ǭ���=���
�(Gv��E1��l0�����37�L����_!�j��c�A�.��*#�����ܼ����-C܎�����f= ��.vo�>B��p#:p�B�1�+x��ۘw�6Zte�Y������d�Wo��U�X!�HF���:���^G�9��Qb�fY��î�7"{�M��O��֯*���Cb�V�*{d'�.ڸ�<ʧ9��~P���W�3��Ѿۗ&%;��ͱ��E�;F �;�'��skW;;Q2*��N��kҒ��mc�F���;�N��u�{w�Fs�ӈ��;�3n�vf��h��^�#�g}��H�n��yW�c��'d[���J����mh&�m�ҖͭT9�K�u��h����^@T����vG>*�F]��|ȍ�VŊ����V�Z�\��n�'�,��vi99�EaFn ��w���7�uOY|�'Gh̅͝w��v���mq����Lt�m���,��Ҧ'N��ڳ˞�n5�3#���Ȧu�s�C%ݻ�V�U� �h>��n�<�4�1��o)p�Z܆�9SL����qjg�/�W^��]�1x2f��Yյ�E^ąwm�ה��i-�u����7��ӷ0[ơ����ˆ�Gz�a,A�6­p��@��hBs�ty;���D��� rf���Suċ����O��YM��{F���X'K��ZM�@����oFd�z�s*�c,ҥe����"�w�NH,��o׹*⓱p�}�̵��_\6�`ƮnM|\�� q�<n'�O_&ܮ�����Q���Iҩf���y�sGY�7��6�Q�MY�Bc)�砨{D�>��x��q[N'��d��k=���/���3k=��余`aZp��}݃��K�9�V��F�ГI�1�[Ȩ�k����ar�\�9�?@��{΍yxg���t4�z'�7pN�:���ܞ��]O1��z�y�CoKf�{��ς���y�%�����;N���ۻ�$�8市W\"��ɛ�r.q�Z�~B�[���'�����w]ߏ.���{�y��}hެ�)ظZ���6���{I��E�q�������k�ލZs���tR�����νyS�N+�n�_����=���u�F���U>������=��������At;7ԦM;=l�G��PPX7A=��b�'d[P����i�5�Ӆ�V�ǐ�ll��_h)���ѡ�`�����il����۞ZF�3GЍ�8J�1������ 7 ����ۚ93�2��9�,F�wv��]�N�p�VV��Gc&�����KU��D�S��j�/������W��O��hQ���.�������i�s�\E�؇z�6�/I��\�l�<r)֪��k3���7�o[gf�Q�u�I7*)�r��OQ�::���b6�u躮eQ`�iU�ėf�Cxq��������k[O����G��D����#zVg'�%"v�u�1)	g��K>��G7�!�����i�V�]�7��[�1�yq�,p7v��o	v�"���ܝ��).�=jZ�K;|�r1T�۳|��3*��Ʃ+���P~f��)9�	,�\Yރ���-�L�|�C���?1��:m�p�
�%Q��@K��&�	��#kc8i��:a2L��v*icW���8�X�V9�{��@���zt���oES���Ħ�����-1�V|��+@��|��u2lk���M����^��o�;}��i��b/���v�)R9�w�us�f�X;�]�!��|��Y](E��
�����xT��.5u���u���#�7Eʸ�f��h�Jf�3��9Z+�=�M�rٛ�֐(��9ZQ���G@Ïo&�@I�_�ﾱ#����j���y:]mc=|SPʗi��r��s�6'�l�R.�jJ����&�S�B��VP}���_VGr�E�MP8�0&�I�Y�J�\�К�^��1z�۸OD�F����z��=�k7�����؃w�ːXK�Sq6z��?�'c�7�o����MN3�[��gk量݅/0<-aF��m�e��v#�����;��+�׺hp�((}��d�����v��[k�jqW��
�r�n���ʱ��ݘ��7�olۛ��k��TR��G�Eel��VXϩ&�)�r������&C��,\UA��1Q��ƹb�L+sGY�9]:7������o�-����C���liΨ˫�]�,w{nz�N���
ҥ�'A���K�ݦ���s�QD��m�mC��Y��'w��p@���#����(�YV[~���^�@Le�@�!w�N�Yǆ�؋��d���\h *��%ܕ�
��\#'�J��wR/c��"�kEO�Ժ�S�dx�a����u�;�������.����rfU��K
l^ܛ�F#��%.Z��1.�bo���[��͜�.ws�w�>�n��R9���=�����>}/��zW`Į&��������ٵ�Er�ɥ�%���֗Rd[�w!�jgރ#�g�?.����L��h�۠�"(��z�F?���/�+��*sV�7�g��ƚy�2m�G^��A7jq= 5�uȾؕ�Q�4��e��k�}�+�Uun���I]�o&s#��7#����:�����ۂ�kg�oݛ��m��\p1��T�u��5V�{��O2�ou���3c��fVv��rH���b�Ɯ��k(V�;F����ӟFݰ�byFc;;��EY1ee�-qެ���jp��7���g��T�g`��+f��C�ۼ%��]���}�ϧ����:��T�S�eDs�7�n�W�/%��K�'����Ԏѝ`,��$E<�aٺ����<��=���w��1� wrd�jX���m&����ƕ�29M�"��0i����qp}��^.���@���U����[b+�VEw�h��C�ɠ>��E�p�L��1PX�C��{�����b��)��wM���.�DKf=H��!�:�VM�)�p��8)yM��S�M�O�{�w����swT|M*�5Vڊ޴Ժ�5�=O{@�o�Aj
��q��]��u�{��"��kf�~>���U�{!���s�W:�θ��)�J4�mk�Ns.r��%.��_S;�r��::��۹�a���b��D���>��A��(�l�9<�ㆰ�i�����Z�z���:�h +=�f����OKoK���.��m�C2���|�{6�|,j�C۞����697j����>=BuM}:�[������=Ϛ��3��� ��2#R�oA�!m(��ss���A��K����bW�ȷL��5�޹�<��ۺ�̎`ܓX�k%�Q�G���C����Y�磦��ɲ�d1��ܡݤf)�����̀��.����nw�w}�t�\<�G9�F��p�a[�ƖX?6̼��r��Jr�� �;N�K���y+m�ș&zŚXb*�n|;�U-an�u��Q�o�j�f,�����%v5���"�(mv�7D��N�d8[�q�;v����9�@�u�[���@谣=��|��9;#�\�7�h���Ĵ���(��7dl�&�f���+k���Rh������9%ܛ�u���ר�����r�3b�s*y�����9F��95`��/3�9g\ ���o��tj{f;�Z7��Ac�O��OY{w%wd��n���q���@��&�\N�s~����_gV>}(�RvB�B/)g]�j3��e��|���h���_�N/۔A&���^�Ҩ�=C"��,H��K����F"�-��z�{y��};�G�lEem�>�yT^���s�e��-y�t��w��6�/I����f��#��5�v%@�|�JC����5��e�3����nr)�r����i����%T�I�kz���H�D��\H[qAp�	�F������ɦr"�fo�Zpŝ��oJ2z0��֦\����]�Y��k"y���־�����l��]��Y	��h��.�1:voLT�S='���A#�f儸`��z��[�B!8���9�Fs�|�_9�axnXR*o�&>�xHI��i�.9nPǜ�F�����8��コ����j�*��o��෸,j�wHNʎk��s-+��h0iT��:ʄ]�V>*�����%I�>U��n�N����\}����m1|�Me���|�Qe8�x �+��뇤m¤������=<$���wU�����M' ^��ir*�;S�N:��cY�nt�=co�HR���W�.�حU}��K5����q8���������Nw'md�G���{�Q���칎��e�ǵV��~���#m��C�Ϙ�+!���hFÉΨY=u9m�gM
.'���Go��l�w	��I��s���n֗�V��	4�k��!��PL�} ����v��1ܺ�|�T>��:tI�����Dak��xf? �j�sXˎ����L�N��>X3g�Yt汜�}�jy�=�ʶ�T���� u��Z�7����v�Z�7�r=�t���S���<
���Y�S�5�\+���3bo�%<�N��4*�+���WEɆ�ޱ�m�.�l�����P�dKfox�K��1_�<�y=�Ay� �I�؁��4���]K�$��*���!�pܦ@��Ѝ�� %+��Q����E�:<�=6�Q��[e��pt��Ż�	�a�f-�ے_'�u_�kY#�E��|�N��S�x��5{y>�Cf�� զ�R�0�f����?�}�iw�R���Λ3�溜����iC;*;
3$�!��k��j��T)}�9rQ�����t���Z�w�/(�oW,�MdN�7��� -QQ5.��Xz�k�Ժ�6/d��'�F��뷂{,N5�������;�/v{ZXSe��o�uk���(�ɜ��φq��5L��(JLX����K�؞�kR���Dؿ��}�̵���Ҵ�1+��_���H�B�ڝ�G/o���~���-�ަΆ���Λ������]v+WZ� !���u����.ϰ1D���Z݉\W3��K>�7�7�&��.�z�<��<_u�����}�����/T�W����X�2�;r��⩥Fn�3}R�S�L�c���M@��ϊ�:�����5��OA�Î��;��'��x����^��q�NFµ%���cG�+�O}��'�a�>o�ql���Z�qI�jv��n(�]ET99�R����R�]za��xfiE"ZUңz��̀�E"OT�Ë�e ,�bf%����`�Gg,B��A0�=��C71����})%��z����MN)AcR�,܀�e�	8]�ܟ6���mT�}w�1n+̴�͹s�>@��e!H�*}��r��w֬vd$�aXwIu��=Z�v���΁b��Q	en��׍�"�-4�|Y�h���R=P)�GN� ��.�fSCó�&��"*���%��Q����!��(�_^i�ox<9���&Ǿ#*O�o1�!�5jV���5Z.\�t;50Yr�'�peꈜw��2;ï8�-�Q8(܏��G{�QR��I�����2��5cI2Ѹ�jm�s�b�[�l׎Շ\�[ކՑ��z��Oh��cE�
�;��rV���e^.\�C2�F�F����#�9��(��f5�P���h빠JSs�¹����i��L���7�'\��@HQ�����
=[�q�K�Q���>���}�%2ڵ�p��.�mfu��4r5˯M�1�--�2���o!c
0Ӵl�m���+d�W�c12&d\sm�i`�{���bM�0�~�Ӥ������]k���D�R�u��Ę������SY�F�s�M)�Wln�P:N27��}DŹ9���+q�'���7ǛK�Y� /_\ݚqp��hk9Jn
'T�*N�m:Wy�c6�am\�t����t�Z�/σCB��\
:wٟN��F��G(fm]6��S��/�ل @)M�]A� Usf�8�:䬫srW%���m��S�j%2���i�ɣRbo��Uݪ�B��X&�Lf�5eW^Gn<5s\4yWr��ئ73;/�G�g�{X��>n���c�++���s'�}�xD�֡e]�}\eəM.�<L|:�M�9�����\��}}q�*����*Ҵf]��v-n�������̱D���:�Z�Q��v�}�v�k	���(gL�.K�%<X��q��x�k�qU/�k��샨�Uv1�#z��	�ǭ��_��0����e�--����7$W��	5͝"eUmv�U+��j��0Rz���2�3˼��L�ݸU z�+���з�[�t��wr���bF�#m�ov�vq�Q��N�i�gH0�`J���T�5ۺ%�8^-��r��_:�͠��䓡[G<��AE��Y��)�]raދDy@:����Yr�v�K��C��#���4)A}R��:m�� �y\��u8�ĸ���ҩ�����5'P�-�`�#7��2����e�Br�MΏ:�%��q`�v�o8�O��R���&pe��w)��&%�D���ޗHE��)A<����.يw���Igp5m�Y�_C���L��czdݰ��8>]���2:))җ>�|���J�VUkٙ(T�e��1%Kh1��UJ7���PYY+j��1ص�R�օ�+��kV�"��*����ˋJ�����LJ��+Q[d[��pkZ��Jʅ`�aU��,U�Qd*-����iE1�,Z�B�6�[aP�Ҍ�2T�*�A`��Q
�*�����b�²�LL�6�JT������EX�A��Ym�R��Ш��(�eR�X�k+F�Z5K���3���b��hE�5�0Bو�\ƮJ�[mm,X�e\��Z�Y(	Z�ҵ9LE\`�e,ĸ��E�XTZRԊ�X�"5��*�9��Kkj����jR�DEkj�ѱ��b)QJ�-(��D-�K�cK.32�!mm��F�F�[~�����]}��C{���+tur\��8�B�)9�[������u�-4v�N�x�Y9�L�^���+}S��_Wڟ��I�Ħ��%�MP8��m��![��&�quļf�oP�8��L;E�w��m��E�y��ѽXS�ϵ8b������%���Y���Zw�����y��qGtӽܞuc��jq�ls�7�n���@�8�<l('k�'���f�wU�c�[;�A�e�O�>/Q�p�@���@uf�Ԓ�J�HZ��q-�u�_ǚ޺MB;�r���x[�D�]U�){�Vm8DMV)p�I�M����>��r��G�^��ou�N��u�J�"��܎sܦ�M�Ŵ�W��^��o���	��ف�r��k蒑QǝwD�N�kr��[��s�i��ޯ�ٍ�|��Z�����g����9]��êN�`���̵�����yAS�R�6x�N��j$���I�,ɞ��f�u$�"�˸��[��掳9&�R����3���M�mjz(1V�2���J���^[�W��D���kρ��9�k�63��1����|�yWo^��7�C'�����r��v�QrW�5���l��\%H�-�o5v�������X�����B*e�I����������c^�4��}EyW�8~F��)t����cS"�tɲf0Ž9�/4�Ŝ*��pQ鷬uä)	U~J�Ȁ�M��/vV�PhY0#��̐a-��N7y,cy�n�n�󦣑���t�(.{QK;����y��	�S�Y4X��ٗ�ƹx��+Riߤ���y7o���֘�X��q=��+9u�Za.G=�>}̮l[���{"��f�Q2A�H�s�Ti=Ӯq�����ȭo�#�u�z��b�Z���n'�
�ciU�Mk�z��u���h��vvH�f����/��5O�~tEOD��+�E�P4Ǫ�7���j�A�{�Z�[���f�il����w_a���;����-T��=�i�E����t����˸�.������b�}-����0%�z���i��Rnu޳��r�{x6�ݱ�殮yɻ����XT8�X�6�]�A��T{^�Z�-R�S�7hq�O#������M���_"�>��[�7w���I(����%r��W�����g�.^�Ôn�wrl\����};��Cu".�pu�,e���nk����ۮ\�|���K\�\'�v񫢵.��J����g481��BI�B=�#��<齵��tPD�fc��d�}5�~�Ʋ�8k��}]��s�J�G
i��Y�����ͮ�bM#N$[�1�7�=A����7�]�YiZȞoq�����$�Մ^,g�&M�կ�o蛒\��
K*����7,%Î�����I���F��p��R|��ǅ��U���'c�|����fqwpv��az���#;wϬ��L�8��xd~�yq\G/��/�fhW� M�YikNF�GR�E�Į6���T�ƯXk,�����{;���Z��f�_JSi�'�.����)��F�ϵ���A�g��dT�\�h�ڄL��������$#Oeή��)���Þʐ��y�S�1�W�R#/y�y�SD[�@��]�]˭�/��i�̙������{V����S���߲|��:�e�3�E&
���Ν�{	��w7F���^tr��������L�V����1H� �.�<�j�R��8be�����b�X��KyxV%/n���]N3�΍��}�ǆ�LR��k�R{](�q��)�ՇTpێy�W��MGxj�\�2������M�5.	h%G&�.�M*K��?��9�N�#S�1���/F\s�S���f��;���:Jz�t��\E-���.�:����|[�ky���7�i����c�.���4w���#��`�&1��{�=6��]ٰ�9�wݜ���1\����)����c;;�WҊ���
�B��)I�I�}D&+�m�w�$4�_�N���$��ε�K:��a^�'�� �@��fVIl�*�����!��9�*���� ]H*�=J��Q�ǳ��%iS�Q���'yn|�Z�|��i��=rh����D��"�bv�5u_�AZ��ۋۓt]�E>�e�}/^qٲTܓ�'n�5a��˶u&��W�vC��f�$��yM�n�ֵ�LΛ��k	)�Z �/��}��oJ�ֳ'rV��h:J������C��z��	���4�J�|�\�	ɒ�L���!"�S��Lf�]�� ޗ�e���y��$���c��s�;���^q���LG{(&��5���l��Ni���"�ɞ���St���6���t�Ϙ�}����� �w����x�·ftS�LT!&���D�_U�"�#�ۄ�N�'���t2U*��ռ7tnu��7	�����%-��\�"�=|S�M9T$�;)J�)��	�/c:x��8:9Q��qb�P;:�I�W��Qi(�Yo��E�MP8��pیt(���h��; �f�������g|r�ED�I��Ŭ+4s��V�;�zQ���\�R�'����ic�в��L�'ar=��q����[�����;νy�T�S�Tk��yT� ��qһ^s��Z���PG���{ʭ.8��M��<�/��G����}'�S�ەm]ٞu��N����^�����S�pCY��%�v�`g.���z��Y*�E�qx�:�Q��8_�ܝ�����Y^+6}�8;���a�����y]r8���j�㤈���Q�@5�������Ex�OQ�c1�W�յ1&����e�PrAbX�d|���Ɋ�2���d�jv��t�P��r�x�d��� �nfw|�
W҄vOX^��:�Ou��w4�J��gx���Ԙ:����q:��I��)�s�]���-8;�;� @*�s��rA��[ug1�ۥ��C�q��)���<�䩸�],�qn�mZM;���Z�ʹ/�}-b?�6[x_K[����i�F����j�w;ݪ��,0n����|�S���/%��v��]f3B�p"P���V���r:;����Zu�:�o�d� ���|ӱ����{K�z�ޏ��\�}Ѫ<ug�x�@,�2o;�+��Cm��+:��P�9|��;q�M,�7��;f�����ύ%-k��4���f�p9q9�8�:�b$�z�ۆ��ٗ�ƹYlR�Pmov�%v��O���V��N�yCK�����(�.]�l[I�n5�6�7Gjgyo9�Qn��hZ 	q�T.�Zn�V�בݵ�稧@����^��V�#�N�����-���M��eR�Լ�0/��|n^P�bs!�:�;bf"�@{�)_�����,�i
0�w	f�IX(vus/.�a��嫥c�m�vh�a4��9H|�gAԦ=��<��u�:N��iV����5�������H��� v+���wm.�&/�N��z&��Q8�4��u˙߉]�X�2���M̝�h�=O�%�t��-Tє���N�����M�W7Fy� Y��Q�q#7���y��޲�������1w��'ڧ�Pܝ���zڦkO.P�8�qԞ@T���ͽ�7�#䋚W9���x��1�N�JJ��݄K�5�N�q�NRM���g"�����J�7�w����.6�P�y%�YR:�6o��	g�(��Sp���Q�j�_�SN��l�n7��A�3k�����Q#��A��%ED�{Jp��x��!<�ٙ�oQ��83�T��z%@�_�K�7.S�r�h�r������^N��8NZ����Ӫ��'�v�%��$	 �:�]YP2�[8m���d+f��L�Z�o�Η�cԕ�`���#k� ��5HB�����˱�Ŵ]=��SS;�p֙sn{��ۋv0N-�G��ٽOI-������-⳱�,8n3�_w�J��0�ޜ���+�
*q^�3Nt3z���N���oV�<3vk���p����T:�rB'��G����T.k��t>�^:��md�h<�{4T�����=�N1#%�E����]��v��z] ��E^;w��Ġ�Y��s��[H�~�j=�VH)�8����G�8�2���u��v��ЗT��q�u+dݜ�5c���i�+\��G���WU���V(�fN�yK��s[;������SM� 6�:�1�1�ׁ���.�@�v��Q��N~����;�+=����Ӊ;���������Ui�ܾ�ۖ\`�����o=8���cÙ���%�}�[��99 [�Q^8mׄ��J移T��c�������M5;�TU�/��<|[��Qn�GSv^�-Ɲ׽U��Ȭ�f탕/��V�l�hQQ��R�7��om��P?*�[��>���3�w�5�F�~�:#^Z���^�v6
�^��p�#�����,WGr���6tçl��UbX��eP���>.6�:�!��S�.�q�v�̚j�ᣕj�n�� ��;A0Y�'F���[��-nU�t�nQ��t�o/h���'I�4�f�/����\Zyc�)�]�0NewL�vP�t���eZ��Q%.߭��:�{la���Iy@�f���I�"��/�i44���we��m3�M37Ƥ��z��їȬ���[8�����=Xf�j�B����]�r��U�&N�[�Rs�3��y�:���&�^7��=��\�7�@��=�ݝ�o�@�0�p��2E�0�z��p;��ɣ݆qk�͐;�0��c[�Х�U���եZ�ۓX�k$8(j;��p-y!gk�={>·ZfJyIMbN��r^�$%x&�}�l�o�MG#�
ݓe ���#{p����95w��J��ҽ�1�Ya�e��>4:8��987.��[����`�ku�{;*t_u�r]p�i�!%�����OmN'ū&���y���H�gw9y=��������.��w�'_�`�si��d�������]�>��B�hY2�6���P�ٵ��狤)1^Yg���ls#6Z����Y[ܺ�A�[��4,7uu9�D)���*��x�������#�{���ûOm��t�"�Z��9�J�8e�\�hͤ�)hi�:0-s���s� ��`%o�f:ݎ��NM�M�q�z�q8EE�F��}�t+���r#�� �#Z�������~̠������e�\M��\v��k��ea�/��E�㦫{Y��׺~�rʿu��	�u���֨TZ�~o�[��퍛���ߝ�9�h��/��N�'e^D�3�S���,�f%wq�O�c�hpn"u9��yM2f�|���ڼ��*��g.E �GN����.��p�S�����8krL���Mo:��I�g:��N(�������*����##Z�t�n���;�o��J5d-6����.y*�V[��u�zL_��@i�r�\O�=��h�KP�'_(�� ��r��#mRL0w�j3�<4Owglqo�����^Hm�]��}b.S��j��{!�Y!���?.@'e}�W��	�W�,]Ty�4WG�̡��yM!�$�`�vJ��K��AB�^���7a(^�F& �k�坠��@J�����
,%hv�dk��Lt��Ws�,���-�Fm��O#6���m1�}B�Np�Z�Qt:U����̓L�:�M����/���N�J�g��QЬ޸Kuܙ\�^�Zmb((a�>^��83Wn���hf�M��Z�!0_əw�h�h���ms�X�]���eh��˱f�L��n�u�T�=�M�U�r��a�4��Nk5l�.W���F�A�������m-J��o1M�U��D�Fp�W��n��)��]'���/C;�U�څu=���P�"H�����������)�+�\˘&�*a0oƓG/p�������:֐OB����������]
z)
�O`ቌ���()��l�dʹ�4�"�yH0[�\%��ں��J�K0�4��a8�-[Z#�E���0�^����a���q��ף8B�X�����z������;�����<"�]r��1.6Lu�r���;@u�K&]-ȡ��t�WpݝkK ���sc6_i��G"pU�M�J4�v�wv����}ЋW­So���<� ���E�&�Տ%���]�e麌>HU����V��4{��\݁�.�WO�9�Nuj[E*��V�E��N;]�Rw�_L����Jr[Ɔu>�c&.���,�dn��p� ɡ)[��N�ʻy�W"	��+8��~�4g�V��-���m�$�o:�6�n�*��m.@�,��C|i��5�w��W��B�ٙJt
����CP����V��}�0�t�`��rs;{6����W��m}I�%=�Os6v�Bn�ι��X�u22�7��v	V�z�eJY��i�zpW����}��m����O	��qܛ�:싛����W�}6LL�糲t���JģT�6�%����1�q
��q��
V&1M�}�;��Q j�W��#�����H\�|���-2����Fĳ..���t�;� �!p9�J>�VN���7t�[ܒ�yf�y.1:��l����>�m졛�3*��*Umƥ�,m��v�����w�mn��\�T" ٌ�h<]��Їr����)c@�t�� 5c�0�t8o����֝f��uM�"+:�
@�������C�&�2���O�u
���؝
�ns���ͩz�q�l"Ef��eu�+�SUmkK)Z��H�c��cfՌr��ӕ	��7}u��;z���k��p>h�GUE�t���؍b�%�c QdG�q	:���=���i�U��ԃY��ݖ����\jwcӶ�o3a��s��ӭ�k7uܤ=�sr�;���g�\��&����X����O%����
;�ouI��ۈ/����+1<FJ�#1���ض.�4��:�X_H̨y`/�2�;����t.<�����*<�������w4�_^I��Dj�
Dk)V���,iKk*F�D������̦E�.+R�UH������T��TEU�KcAJcX[b���*(�%2�*�TE�Jň*ʋQ�(�ikE+aU-����!PV�2�̙U
1`��YmAp���PE���ԍi��*.��E���.`6�ie�*���l���E*���Q2ʙR�`�J ։Z�(�Q*奶$PKl`�m-e�(�J��G�Q��
#Z*����W�a��-�%2��U�+���+E�V�����A�+
�5��B�*։��&*�$���Q-�E�c"�VU��DUU�UVՋimDYm�Z���+
��1Ph�V�R��j�,U�Q
�6ʉmm�QV(�*��ĭQ���QQ�V�Ҩ�U�6��e�*"U-�JUm(L�J�
�
�Z+-��Ģ��i�U-��dU�Ke��eaA�c�)iH��s��~�o�z�iGn]#2N+�<�T�"�-����켚��5nX`��:v��hL��5�AɊ#/,�Q;s�#�ͽ���[
9-Q�����w��M%o%�v�oz1HJ�4��W;J�ê�w�Y�z�l�}�>�-޲6��e��g�lg�Ǖw��K��~���pCA����:�����r�3b�i9�M�;ڟ)�g�\ ]���,�:�df	Y+���܊�����<�aN�i�Ѯ�iv��.����Oך2|��:GY� �d�{��;�v��V�-G��;��>��ה-�Ԋro���������`�u�jI.AU�e�-�2��Q��)�u��S܂�5��z��޿���c2�/h�ѯ�|�*�Seu]��V�Pfn0�������ˊy��N;ˉV&!;&�0��\S�Ɖ��/�q��m�M(g4(��&�)�r)���ڬ�[g�Ud���]>�9���
�	��Fp�·<k�t�x�U����Y:bu�彏�+i-�^��v�5}ʇ2�G].ӽ�z��\��,c�fK��*�o�a�YC㼳�F�x�+&�2����v�ϥo��[CU˫������ft�J^��:�T�)F�>)��)�5] {`�bw��Nzs�����'�����x�z�]���IZ�H��}�񱕦��/������Y��$�2"%|��%����U,�j�$�8��%�F��g�y�K]����Ӫ��7'ޚ:�`��6�
fN����_��r�7�S4a�7�Z�ks�ޱ��*��g,�|�9���ۼ��$�>��D��2q�W��n=����t�2k�-[]qr��)*�x�\n���jz@+��}�)V.p�k!�e�gd�؝歭(��U3}-�V��\��xD�ud��s�j�:�u���q�4�򋙨*�8�,[���t��M����]�������v��,-?goo>�;/u�P�>�\��6�:�(����t������V-�^���;��k����'�ϻ���Ӑ���N��{�����'���J�KñA,���Һ�2t�Ȗ�H�g��u�Ϡ��/���v�߁m鲈^�\�Z�B�z��x�R�s2�J��7sx��/Ju�ڙm��Z��mw��lc��2���2��\/zd9�T땸�G�Vͳwe*u5"r�֖zt�ĵ^�x�����ɬ�v�=ϋq�n996�	e��lr��Gn����r�!v�i�ve݃�ׯx@�z�.�Ƅ'����u���g�X�<�Q!k�y_�l���lu�Ϳ�R�/{_��'��Y�U|^h0���\;=i����i��nM}*��n�p�[�e���扼淣w��)��}M2�����Wǰm����P<�A��Õ�x�[�s}C}�G}} �jv�'����Y�Ci��i��5$�3��1�Zq"������{>;�y:�	�����J��l�φ%K��2���N�&!�/�ǖ�j4r!+r��I�Z�&gO؎�OA��TЧ��#��M�Sؼ�' g�`.@��p-n�⹒�$� ;�;��sf�35Gp��)�Q�zƱ$�5�5.�y��{v��)��.�w��߂���O��`�NwL���T�Ub,79�s9l1�����Li^Q�B��/�3�J�=�������9��CzPz��X��\�s:�I���8q,>���s4����ۗ��ю��Fo.�5�BQ3ǖn���XT�չشG�	d]���:;�D�b�;��n�V̏6�Ht�r8�+�[���ӛy����+��*1,l�q�����-����Uƀ�9+Z���L⹹�uz��Wu�a=���]yWZ.]�f�I�)��#~�26t U��'<�;}Ow0J��k��tk{f;�Z7��@�pŶ�{���ə�w�Xɺ�Z��h�;`�ٿ����W3�K��:���S�ހ�cM��<��a����i0����Z�7��_��e��6Q2�!@�M�ޙQX��T�q�G>�s��z����N�Y��x�,�GĦ���'��'�n�t�!�ai�	�N���N|w��݂�v��B��l�$hi�KR��q�nk����N�6�nCO�#���:8NU^�^�&�Ü��)�w�:r��8�gb�BY��u���nCi��Y� J9�KZ��1ԡ�Ioo�ǽș�޴2�B���#:�9�E�s��J;b�7��.��C;�)��jE�١�B&x��s/4`��9���N�+�[L�-�""��h��i�pheF��Y%3���g^��Y��@)]Xx�IQÎ�d�{8��k��$V�y^�������25�F�r��\�h�g:$;®;Q�A)����(L�#ϰgGT��L=F�zs�{���k�H�6�Kz�}f�L!Ӵ��:�V����*J�䟙РJNo�Kx!��x��UԷ�(���۾q\P��2q�g��6���8��@�n�L�
�
��;��!�)4Z��Q�T�{N.�!���KX�m��t�B� 1����m���	E�{��x�Ȣ��M޲6�-dC�M[=A�r�')Iɺ΂�S�&��w ����]b=yS�T������г�W�]k�W.˩1Z��Nũ���:�_{��g�o�}]<��+A��7G�jÎ*��s�6��|5�t#��zKS����<�O5��[�ԛIR]6q�7�
w���\c��]��_\�]@�D'[>�T����-X��Rm���a�n��eҭ����W8�}�"�T��莫�����Z/ ��XZ����t��v[�����.ʋ�J�\,�[�]�[
�/w�r�e�T��L�.[�r�w�3������C6�n��p<N��n�f>���JKP�;\�W�=���u��Orq�ls��{9���߱x%�||�$��)X�]d�Eȅ��^�|�tse�<���zC�e�6�7��Mmk���7�s�������3��EaE��r�z0�Wo	��T�6�zrp����7G�%�V�=��X���ֻ�jZ����YT:f�c�i,�Yύ�gπ�g�3�R>��}G�<�z*����p��1���:V��ks�ɜ��/�{"��=Dzs�ޣ�y��׿�ZO�W�nM�X�S�e�����ZF%srk��:^d��Z�bWiN^�Ի!�(�	=U���q�܆������:I��jS/g4r�r\�-�����'ϣ���ώk�^�=�p�Ȇ7�7�<-*4�qJs6Q��$��n���)	4~j����+�}��\oj���z;�9�&�dPSw�gNQ�A���G�a�FZ�pd�g�M���>���+:P������Lv�o6֐&-�%�ay�:��Σ��N�mG�.}&�9H��J	z��=��F��iW�[�\u��3�%�j��U���Y�Qg��@$ٛ���I`S����J�8�#h��7:�8i�M�[��w�	\���G�#�a^���`��4��.ѓ/5H���i�t9X��&p��ꄴ{qW�'��^�WO���_#rVS�+��z�
6/r-��\R�2Vp�T�=�����������9�����oӝ���쇩�0����P��W������{�h�>�B*y^Vxy���ԏ>=��G�O_IȺ|:r-; iϜi������k>�>��}y �6leF�`�{u�|�,ͬ����U`�1���2�~7���:@��v�^���~Y�ߩ߳����.���yx�6;��}~���o���B&�
��ϣ�X��-xK¸u̚�̜�����C���xO���l{.5�ݩ[���9���+�)��Q�Y~�C��Ȟ�Ώu����:L�q;���JȞ��0�=�3����dq�ړg��@qJ}�����J	��ޯfcG��+�UƠک�Q���{'�����l{��y�x��Z
�(����*�Վc��^�(MH�ݦ)�ӧk*��"0"���8]f�K��ڂ8��ح[���)^�{�TX﵇�ͤ�V)Ш��U.�8�6�z�qo.���[��H�����l�N��k�]�ķ�Q���[�%�ś�z��il��0�CDM��;5��8���O�U���cL����X��MCq&1�����>�:�lxy�{�]�U�*mx�u&�8�q���/� ��s5! &㪒U�yp=�_��jq��t��y�]ʮ��O��*���f�7��~��T��u�P��&'��T8��R�}��
�dX���f�12����� N׺|k��q�<u*g�k�L����-ą�#_SvddI���1t*t�P�>�en#���z3������#��7�=�_L��o�\:�A��Й��>Dh����=�(�d���K�OA	�Gy��5����W���؆/�m�0&�`к~�Ł+���h�fUn(JR��B�D��n����}z��S�k�'��2�dy�`��=�L\tw�dɛޣ��^����P�C��C0د.Ν��~#	�s���7��5o�?Dà�W?���O%�yK�O���%�99��R,׀W��C9]�E��� ��Ig��i��M�1��(@V��\�Rw�G���)����g��^J�����؜���uí�#^�t�-O=�������k"��D묦��у.V؋F�u��Hb�nC`�Rΐ�j�<�˻c������y��MT�J���;l��g^�~�'Q$.����Ό�L1��i�+iEJ�Vk��i�h���)�O��^,��"ޛr�<�IN],��������߈�q�V�� �s�3�,���i���T�_������^{=���I�5�c����r����M����lE:���=cX+�y	l+�/G���!z������*���J��[�=蚧/".���떫���S�=!�~����ŵ��_��яnT�y�o�+��
?��ƀ�!�o�(�N]W�Ȳ�XzG�%����'>�G��o�o�u�p6����l�2�[*/l���w�o��v��00���+s�T�Ϭ��Y�������'����Vث9�|n��3�C<]�E������'��ˋIv���	P�뮪��S�E��v�@r=��l���<�o�~�@}�0r��e�*����&�����[n��}���3t����b��)3q^����Dw��>�{*z��j$S\	��-�H�nx��H�Kw�}�������C9�Ru߱��㍎�Q�2=�dQ�W�Jp�31mu��U��u6a�O��˨�d�QC�U�'Ká�K�w�U����c���}U����{j=[}�[y����è} e�z�o.Qn�e3!�����K������+.9iV�(+�bD���;��4�ض�`������8���q�K�C�[����1A7l�&����ޛ�$�����ړo��*�;�ȁ��&�f=ɹM��5�i�u�����><���.���~��DKP�hH}�x��g�T&�Y�U��G��>��~Y�!���೮����԰��h.ܱ��;�R�>�����ʑj���RȟeF�L�p�ñ����O�(���D���Y�nI��>i�PϷ޹�V}�zd�l1ד�}�R��FˁU�|�?�cW�{��r�/��~�[|ڳ�~Ln�^#M��?7��7��g�7�P7�o�' ��[���'C�W���;���Q���v�v�$Ӯ���/�7�k��iő��)���/z+������zA���+G�{w��7�߶�|�{R�zz�~�1r���W�:Y3Y��!���+>����^I,�L���/5��e�������W0�ťw�@���ɚq8�)rO�c�g�λ��-�_3'�[�q��R�ܢ�]{��Y�<FǼmNr�20x���*6C�?L�'\���T�[P�b�w��=QK�x�6g+�|�&��z��׭O���3#�Sٔ�]�b�éC���P���+����a��!�w�}~�4<x�?q~w�C(�20p����C'�򏡗e+�u��ji⬇',�M�$<��;O1L�ܭ#�[o��Ы�-;�ɽ"ocL�GX���,5}m�Y��g;(�F�һ��@@�8	,������Mt�]s��S��;�˥�0{>c�JD�,�9Qr'��/r���v���r��v�A�k���Y'>5���<�#�m�拳�q<2��ipq/0h��+���7a�J0a�gu8GGk;_n0�k7�w� ]/M���W��f�/%�ǲ�ev��.٪�w��K�,�0e�A���O�؃�	99��Z�ۢ%Z���e�����.J��u̎�郈��	�]�CwG6-+���K+�R��i��k#ʯ��6T��1H�dD*�����G��n�-�:u��=�m�p	U{I�]O�mV�˜u�j�N�ݣL���c\GP.� �%�����p�!)u�~v���F�G�F��$ZR�:h.(�m��t��a�Ҏ��+.��6�lE]vX��%M�}a�*7B�YK����n�ҫ�Sgz*��_)��u���Q47�n�º�f=&�-��V�B���c��5b��9�]�n;�o��n�j���1�)�|n�K�Bx�ق�;�띡����bo��d����շq7�{�LJ;h�9v"��i���ѷ#L�����ۄU�S�4�B�W:��l�~Nt[�bׂ[2@��ΎΌ���|�i��7�Ff���^�=�%b�G2K]���]�mk���#�Q�L��I޺�Lδ�� ���vA�'%*��m@S��ͤb�;�8L��Fge�N����}:9��?@�=�A˴;��}uff4���k;T*��I�\��W��ˆ�Q��{�z�_E�Q驽/�!dJ]@�<��� 2f�|��'NA+S�*���j�<_,鲵�!ԾB�7�.�;`J������Ṭ��V:W�mՎ�X�*�Ý0�.Wi����rV�+�TãN�
G�2z����f4�9M�aÙ�]�D�g"�]�@=��]e֋��]���Vxs���cJ�>W;��]`�Z.�"���L��;�>I:�0��I¹��fk����Թ�R�Nj�а�ӵ�B,S^�]��K�� ^
�@���\����Ww�?v=n��U��[w4	�oMo��Y� �v��gDҕ;e\�$���y��B�׳S�Ř�̸;g�w�(�C{�Ԭ ǔ���u:����312Fj���ҥ��C�	Z����I�/w����u���^n+j�	:�'WAq����;���+��;F���;��X�P�qk�ޱӯU���@cRݛ���U�[��;z�CnU�}�z@:�[QRz51�mt���2ej�wVad�IF���H��J:l(�\�TI�zѕ;��G�:�Dl:����cG]�|R�hqE�o"���uU��Օ��(ѣ�h֭j�EQDX)-�E-iZ,jT+F!l�+F��-l�b����D-�Q��j���E����E��PjQAj*�QKK�e�J�(���(�m*Tb��eeF���m�
�q�4F(�(���Ҋ�eeJ�����TZ���1U�l���s#�TJ��H�U
��m�kPUcX6�EAKh6�UkJ�1��QB�((�Em*
� ���b*�T
��c-�*""�U(��X�"
Q ���bU�X�&eJ���(�QUj6�Ueh�DDTŨ"1��P�1TE�e[h��U���J��d��mj,Ub�EE��ڂ++F6�idTQiZ���+iJ���[U%K��J�8�"�(� �h�m�(�(�UX7.*��Ā�iF�)bB��b�*X�J�Qb�E�-)��T���&�&��L�|��mIN&�Xa@��i���g,��}�}�ƴL`����|f��� vX�6���{H�giV\�*���(#(i��D�:����Tm)��ǆ}m�MdCO<F�P�dx���#ܲ�Z��!��4���q�h�������
��D�6(�^TG<���Z��_�ON��cC�ʇ���Er��S̒�]W�i���0{mp?n����N��A+���'W|������\t߾��3~�q�I���B_��eq�eu������[��b����"���62SCǥ��eNɬ�ue�Q�rX�j!�U5^��l�xWO���]2~��"��]"���К�f�c"�4<+�E��U�ù⒳�i�����v/,���jG���3'���.�Э�L6*��[;�a���h{'ޝÏye3��;�o�,�lit�Ϛ������(k�P_{޹��5S�{j����~G Z�cȭ=��Z;��2}���].9}㞜&�gd=OلF��_�f��G����� Ń����R�xP�<Aƈk�����^�ӑi� �N|�NgO�c��v�Oz�Ο1q.����v�-�����k����]a�)@��3u7?j�yK�+,gS$ϫ>Y���N��J�LW���0gݬ^���YJZ�r6�4����u���W~��DX�6�E5�]`��7:�܍ 7��I"̑�^)��R�z���ч�.�
a}*���yb�E�4r���r�:�58�=s��;fWo^�i2&���e���%�c<X�G���^I#~��jr;6�w0;�^�~�^M(p���{�~��2�~�y{9j��Lϣ�8'"�I�.5ߛv�l/S�ʺ����ES�p(�*~�OviD�C�^��J�Q�dz,щLl�D���_�ϼ��x�g�������Sq���N}���f�#��Q�)�MS���7�t���\W�/u��}�~~�<�)Ey����U���<UDE䊳��"�T�q�3�����`�m�M5����ϩN�<lx�n׆ݵW��*R�VbK��3�NP�S��Nf% ':�%[��\e��f�!��t���tR��W���P���A�z���S\1۰���� �Ҡ0`&�RԻ��8���5��ܟ�-{��W����%~Y�z��
=޺���sL �P���ǨMSvdB��1�ݚ���KTo��*�9�Q��cc}U�{ã�o�g�����|*�� ��t�ʰ����#C����ꥩf�O���o/��O}*���B�|�����y��7�yC�7��8�4z�Z�yv}�������=Ʈ�DZ���˴�0��\��w�hVĐ��+�M��-�� ��5� x�bɥ��_v#ã%��ݢ1�0�\^��j����}�ZKچ�K�񭀂�u=�sjM|�W]�J�d�PE��,��m�
�;x���ܜ����q��}�@����$ |.k=G�2���z��!�fP����~�D�q�n�j�r����P,�z�~�Y
&��;t"���j�����u���'>k3�Χ�ʛ��|z�v�v#NW����l�K�Vj���ౕ[���\�
�v�����
�]��S#ˡ,����^y���7�t���_"���{>�n��o{�>�ג8���u;�L����3��p�k�_w���n�Sݳ��>���Bc�Ş��w�ǝ�5Z^\��L�B��C��z*�� ߭va{l�&�����x����R��@2���<�m
^y^a{�����:o*�g���T����/�^�Yx�7�h^nLF��a��AK��F$���8���������[Yw3{}Ns��(��a������>�ۑD9Ϯ��T����I|}?k���Y�#>q9F{�����w4=�o�Z�-�E��Hd`� ȇᢕ�Ⱥ����-Ʌ���d�}�����cmA�;^s���o������ψ�9A, �C��W,SaEy�,���b�*A����m+����zf����v���3����@�������TK�ݺ�䲃����F�c@k`�<����`>�o%z7P�h��������g0�Q)A!*��gKM^��R9'nI(�j�8`��F�G�'�J�~�c·�������+��T��U3>UPs9Ң��Q7�Y�ը�����w�P��q^�Y#���Dt{�8,�{*{#�lUê���.7L�n{�Ǡմ�#ӂ��U�܌�)�9�E�jԝw�lG��lx�=��(���}��y��8�=�+���ۢ�ѵC���(4'h&�擥���u��w�T�}�����ǆ�U�A���{*���Z�&^ ;�\tM�w�:���^Ϧ���f�c"��5�U��y<�	������|����2�W�}��I��G����&_�PT����T����G=cK��"N~9+�n !b�B�����B��k��?;���3�����$z�ɣ^߲`���J��W�E�?Z~�TT]��َ��g-õ͑D2	J�U�܎���Z�c�I�{��HY^o.�j}U�i�Ar�sϫ<��mj����D��}�^۞�Yl�A!�=8�=�N��#a{�g���ِG���wtcw�B��z��3��(=��b��uvUzU�WO��lt�]+��r�3���_S����_x**��u����z����R�d�<�a[M�m�h|v]��"Ń��\�HR��g��>�@�	��1T<Y���,]K��πɰ;z��C�r敹�]���ʻira;���=��i��K�e�R��
Z�S�Oq�X���n��\�����or�*�e����|�e\�*��Y�rc�LЛ��AK�|�i̟�<^>�c��cn�gvY�~y�93#<�z�m���S�k�9�.�#0y.�@v�(����T'\���1����n�o���.1�s�I>�+�n��g�Ϟ߱O�mm���۩��)��7�J��U��e�M[��J)Gy!�9]Hg?fCؓ�������U�^��l�ȑ�$�5�I����j��},s(��fTo�ꛯM���m�ɬ���#cʇ�#|hxr�|��?s��pd]�Z<R�)bFd	�+�Q��T���)��y��g�M�ا�~�>ƇG�����sдœ�9�9��'�S�G��e+2lМ�iy�tK��ϭOJ�_�9�\t�*���r�Y���j_�;D
���j���>BjG"ajB��������}.ཽ+��{~��[����JV��T����������=���3�{�fs����>�� �-�a������@�IV�r��"��cs��C��'7��P��4��2N?�S��u.H�ii���S�j�����V�v�d��`��Ft)W9+��V�^�w�:�DS'L��6���o�!IԀx�f޼u�R��v����B�諨6�3}�k�M��SK��k��R�%n͗�ĺ��ZU�����r'jw��s�Wl������e��Y���t�Ʀ�/��K���)��o7,�S!�uǔ?<��������d�a����=�CwRT\on�h��7�&^#ނ6�k���u��.������l�k;!�����Pϣ}^�q(Io�X�__{JJTu�\�P��h�<��j���yu�9i� �N|��t�v<��c��}/�=k��r�R��+����K��H9�Μ�yU�x4�
�Wh=������²�u2O�eڟ{=f�Y;�*q{�ԯ��W}�Y�k�s�J���Mi��]��2����Ƽ�:Kf�t�����ト��3>�W�	�T�����Q�mڕ��qNr��s���
{*����)�`��Ǖ]�]���E��(���D��������g�����f�����Q�ܻ�B����`��c�I��`���릗�UK��}�0�D�_�g�ǃ��S�[~yUܚ�|}��kr���%
'���=���4$�"`�ɚc��W���7c=��W�M��>�=���+:��Ψ�K�®r�|�>�m����j)�It�d�ܑ��	*��ˁ����Kju4vй��Y�n6��.hٹV�A��iB��1�t��æݧ�{���R�>�\�@�X2�V�5���캒sĒo�F0���M��LΕ�n�C"�g+n�o�>sJ�X��\��=�U�	L�Y���Q"�j���KrnJ�J$��Q�Ă���4-��%R;^s�����CA_{��b���tBjy~��nu-K�Og��!�g5������z,�A)�^|��T�z������I=޺��z��\:��L̷]�'jǳ���L׻�[�פ�>r=���Q�(��c~��Ǫ��xw��H�{�fsվ:���o/���C��.�1i�֏|=BG*���Z� d��~�B��g�{����b�dm��	���E�:���R�}�\
�Jd�Ez���^�Df�U��	��B3��[UW�~�g���-��ʟ(3�`X��֡.--�p��!p�+c��b&ܜ��:\�E2���;w���&�T����Rj�dw�{zrp���_Ƽ��MwY����dy^V��V{|8��o�v|�vzv!z��ls�υ=�fȁW�̫_rӗ��f���~6k�y�n��������#�.���y���سӱN��:�f����9ϴ�,�����
��qV�Ｗ�R��=Dz z�ND^��Ϯ��8uy�{~�K�����߽琖�����f�ѧ�t�u�N�c+:�OR�R\����Y�X�*�t���{�|�4(�R��Wf��|��V�H2�<Nm��<L��W�������6^��ǡZjp7�5�\�X����mPS/�����$ �iwdaCJ�Y���n��'j�Y$|fue�F����������m9Xh)r~輈d���*�r�_s������.��O������l�_D�C^�rڢ``%!�l�!�E�y�˹a���qޯH�|7&�j���]��u�c�c<�=�l-����߅ih���2nC�J��]RB����^��^9�Y����9�0}<�t������>9�9�[xJ\�ɤ�|�0`/�C���G�]Z� /�+ij�����̀�}k�"�;����:;�b|FG�]Oc�r�F ���*˄���hb��7�I�^%�ٟD뾑�)��w�P��z�d��x{ޡ�g��S��b�D�����T�j"�[�.&X^�6&��̌�)�9��]9�S�߱�m���Fg�#/��E+��MuR?~���YRL�?�j��GRu�rQGZ�B7�Z�reͽ�9A�S,��t�QW�7a��ܰoÇ��r�n��>+��	W~�
a���m��EyS��v�M�s�ՙ���'D߄�<n���~K�(�����&_�PT��������:^�t����_��q���X�z���0��8�Q��Y4�8�� ެ�:�@q�4��.|U]YQ�&G��}Ʈ��������y�T���+�s��.Ov`�7���lI��ge�w4D���w=U�7W���t]�I�U��_� 4ҾW3�� �t�v�&���#$�f��#��*ɋ�cs����s����(���d{��<�j���E���/T�f	_D�n��u[��z�}�/���9*��;!l7��9��}A��h5^��j���ߊag�w���ķ�?����Uo�GO�k������qd{i���lB��σ����tu䉴��u[|�z�k����B�d1�uvEG��9\+��G䯽�,��g������} �-��&�꓎s��!�j�I؃�(FGf�p�A�ݐ*��kh�n�|�i̊�\��=�K�r2�"�˅O���9�����v��~�R�u�<X*��F����eDf׼w����f��w��w0c|�I}I�=�s�~�?�JR�]v�C5�N��{��E�O����K/=��z"�qÉ�n���������U�^��l��4�5�Sg��T�*1�7m�O�+�)+�!� �yT�^�Ŗȶ�&�w�ʇ�#|hxr�|\ `噭[J(ُD�#bnF�z�����D�^d6��|6=��7�z��zw���|�G�<3������&�VG/7}{�eg,W��Yl�:�[Gu>�\��/x�b�9אl��8��Y7�6�w**��4eI���ڏ6۝]k ��Ὀ��g+0q�9c�i�-���/�!����Or&�ը0wlA�S�1��S� �\'�w/��{�� ?_O:Y��tjR8"{�A(�{���f+>gؤʷ�VL��&c����� NW�}�x��Q�G��FG��lPb�	�n�T�f�Y����U�u^��Ѷqv���#ѝ�/jzq?<s��Z���}�Ӥ����8��:�T�ԏ��m�_(�t7w��i�ם�c֩�s`�����Jk=C��)q�>؆/�]ӡH0:H�C<�*�.�K;����O�	c'�W齺^`�T��k�#��2�F�~�D{޹�����?[�ʙMo�zR���D/�N%\3���˯	�ņ����p�|Y�~OلF�?E������wy�׏�WZ�e����,�ǸV���%��}@��t&>ņ�<�R��g�/j�}(�=���s½ϓ�[�"ϡSʗ��$�gNN<ۭ,��tC��p�w�:w&xs���e;��׮f|�9�د_�����>az�I|mNGf�N�v@�z.����wK�=��o^���G�]r����ښ�9J�t6!�ƣZ۵+ax���uc�)��#d��[�#�����$���{4�>��}�)vjR���t�vY+�[�[�71ᬤ�C�&�M�V@Xu�Ѝ ,�>�)���V
ν�u(+�ی�x�,�K$��y�2Y�"wV����V���Ց�c9*4���}pid�3ow�6&ҥ�^�v*�M�S{��-K{�����"���9���v
j,!���"gR�Q^WVE�v��v�b���]���aނG'���p�Xz�'N��P��v
��{9����$ћ�� bڄVh�wbj������ԙ׍w�C��P��v6�v�s� g�����Z����vY�J�P�Vӱ1�ᮮ���^�uz��5C�E`�J�pR��\�x�J�d�rf��H\Ԏ���칥v�)���U��:ͻsb4�$He�I�`ذ�j:��r_Z��u5�*ܫu���Mv\.j�.��r|��P�ֱ�jZ�ӗ��J��{�{S8I�:����X75Rd�Y�ׅ�[K0"LF��K�!ڶk5A��Uv�kC
�����Y��,Sew���t$��<v�W�ݯ�+�V'�N��@��z�����S-p˿��w-���H|3���W�d�4�i,�ɻ�[�ԭ?s�iNs�0�b��<!A:��t�&�CZ��5c2�
�[+����g(�M|���z�-_2�7#m�PC��Aȩ���Q�3�2Q���s l��[��w���ם�!���S�V!iw%���tT��g$�HV}#s��y�57�#f=*<��db���"*�N��*n�l>�wM����`�!eXQޯ�K<�8`�� �b7�<�*��̠�9�!o-%�}��G�سv�ӜH�5ύ�I���T��pVּ3E7�\[���E86%��9�{�f�_'lf��#���P�Egq�n=8�v�����R�����6��Pe�\��*a5��^�c�9:�%�n�p�Z������I5��CvT*U�+[/V��ܣ��\��7wg˯r֦�s%�"�fr��2�W�FV�E��wg$v+i��"�h�|�7n�5�]���GVL�yG+�[��+z��NB8�Ѕ�B;��}Gy��B����v*�)ʸ�)�{�_Z�t��1�4���({��m��/�E�N���롄V���J%q�U��(�|�-��x!ҕ%8-��=���m��f�%�p�Z묈�V���[M�#�9|����gI�8�n������	BZ"�~=̣`k���t�/�9|���G;w_1����
������Yݜ;^Q�6*Otx��y
Z��E���]���l�&[�S�:�vaR�3}�ٌ�����ZR�}}�����b��e�Z��i�OT�n�M,��zމ��p�Su�)(澭=�h�E�90dK��|�]5E�xi��ĹW������k�{�$�Ю/H�{Zz�u�9�����6�vwtW�K��`D&L��=��ɼ�r��+TI��C�(P��
�[e"��U
°Q�,T`[c����TeJ�QC�D��QD�TƑTU�"cX֨�B������QJ�"�`�#b�e"(�DFB��[j�U�kjX�l��"���r��2���b�E��֊-�*�e�eVш������R�����TDYR����"#ZK@��A-,b��őV1E`�,U�Qq��UH����B�b-IKj��VQE	P�5���K9KiYkl�Tb1EF(���PQEUIl�b���%aQ`�ZV�ы��DeeDƈ��R���X�*+iJʎ52�ETTF
�J�Z�A�l��DE+��Db"*"���DJ�sY��mUA`�ڲ�U����Q2�KJ�*�Z���iQ6�QAE��h�FQ[J�[(6��˖�h�cF$F�JP���m(����[iE����4H�@P�*�Q��ڰ������Fql��wP��+�f�fwP�o���+�=�wǹޥ̺|�ǭ�{#�C�e]^�x\�zs��l�;��t��1!T/�E��2�z%��j����_���������/�#���JŮ����m�Ӑ��zmW��M� ~��*�&�ϲ.�ʣ;�u�s��>�H^��ǽO�:�؟T��kVQI¼�����\xᑞ� �
s1>A��+^�l1��ъ}�|tí�̛��s�g�6I��<]���H�N'(!hx �9���}T����ˁ�U\���9��[^;�ɩ񲳧~��~aw��#�jk��A�Mq �ؠ0`&�R�I騪=A1QCW�������1{�pX�|�/>��j��W_�=�� g���Ԝ�ۚ��T\B2�ed�쁹x9o{9Y�^���>���������rи�����{�ëd{���𭜺Ѕ�hE��h[�k�c����hMSv��-[@��T�3����G�^@xx���x�\uS���Y�m�>ٟ*�70j@�{d��`�\�:\1l���X�?+��6uy}�U���$-̱��C�ƔI���`�`� �7N�3�^������~#6>��-��i��䭀�?D��(?���8+��(ЗA\�__d��	3��|�N��;��E�x�֖>�ͅwv(�\��ӭGu$�y�p���ӷ	/8T�4���JN�}a�M"�&�SO�W]e�}5���s��Tk���=J��#��J�ՓgV��$��{e�*���\��>��� �н�9'�U#�xs��MwY~��eo��8O�U?�/S7�9���<���{~��w�9��¹�g�ej��ɣC���CK'�Y�s�����7�e���̟T���d
�����b�N�S��ΣY���9ϴʰ�*��	���q/K�S�"�t_��;�f-�O�*�w�y��mS�����V�<�kG���I�v���m���qS-[����ﰸ��G�9T����8)K��E��d���*�r�_�������g�O���q��������/����S0�ܰN�-;W�E�ͭ2��6�w�P,�z�O��v���߂�R��"-�C"00���R�9��$���mM�v�ڴ��-_�;��-ɏlD���:w�k���b|q�����2�r�0�P�U%ί�7w�x׾3ۮH�س xSf�;��y��6'�d{���r�l�s�[t�3�a5�QKJ����W�zf8Ґd/��y%�ߖEg���$6#�]�����pY��T䈷�I�HE�J�������v��M֓m�vi=�wa�&��jLypO��*�2�R"ڮ%������D�����5�����f����W�M�^ԥ�n,���,�������cY�p��@�,��.Ғe�v��]p���[�9��}\�:�� �F�<T$%]#���D�(g5jK�[bz��b}i�lg9]�O*n�̼ z�E�]�R�l+�o$ؑ+ʮvӵ�z]z}��=]<$��օ�U�z�侶2 ��p�Ε��}�$��#�;�R�MT/dMS7��Ѭ>��N��	yޞܺX��W�My�y/`�8��*r<��o�zd���̿eԄ��n$T�3���/���f�|V{�X�>�#��NC#>k�=;��(dk�������(c�'��E�
��d}�Z��_w��Kz�g���ճ�U�:/��y�*di��G���F�����F�.g�����m�0b�n�ԃRtxUS�!����Y��t���Od,�@#I���ǃ���E�5�D��׽��J�Hp7���!�o°wЇ�W��6Y����AW�7�[���������FYɉ�����5Y�#����^I;�P��ͺु�"� �"���@�s>I=4{��Ů�e<�Kz7�3��p�S^~�Hq~�x-�v��ߟ���D,E�7��oݞ%f�M�-T�'o�x ���uǻ5i�G����#Md��	�5��ókL�`�_}������+2}����mlU�:uZV�ɚᝢԐ%5u�fM� J��w�>1{y�Z�:7p�%�X��R���fк�VVC=����[h���(�̊�As'[�/�n��ϝz��J��7���� "��\�{E�wy�/t��]�\=�q�)lz&�1��C����4<x�?�*r}�ej�x�`�rY+�U#~ g�+� ��i0t��LCq�
��KsF)�_�T<�C�ǋ�.�����{yY�>���ZB�#�D��t
s5*��g�Sa��s�>�����_�OO���g=�#;��B�ɏ'C�ȏw�+�����'!5>����M�#Alw�05g��ܯ�&���V���6�tA�a�Y���e��}�������qWPbИ��h��f��uT�T�T}�N�Z�C\�~涧���;�Z��]>��t����H#����'&^D�X�D7���X�w���lz���p��xx���Bk=C��)q�~���b�f�[�Qt���]Yu�ⶽm��f@hN��z�o.�c�\=׎G���C5��2=�\��/���dᛮ�]9{�;eA|x�D/��5ciIϧղ��p�f�9�O����>L����1[a�Q�񇱝�sh�����z6�Jwl�r�%f����%rn����i_d}׽�j��,���N�FQ޺��]���ȭ�ۏ�k1��9��5qc�s��ѡ	��@��8u����uo�5Ϯ,�ś5�ivL����o0��AW��%(�s���g�+A\N�5�=}/.�ç"Ӳ�mϳrN�o�����yiI\�v}�7~;>��Rgגw��%�UR����A@��AЛ��&ܻ�u|�G������VwX�9��3q�垝���9��~���z�I����T�`w`�zo���|=�;�����M]iuo�=��g����p�LΦ�I�T���CˍF�v�l/S�m�c��w�t�k;Ϟf2�x�����n=�n��N'�l�D��'�~"<��x�{!�=�,�7x��:=�HǷ�-�� q!D�l���.5��Ij_`�iu���Vӓ9��Z����X�|����1�N����r�7֎G��#�:)�P�lS��A�Eҵ�b�e�y5��zgl'v{�F�ݣ��T+3��s�])�G���������'(!!��Nf�B@M�RJ�����977���z�a�Wn�ZZ�W�{'�ߘ]V8,��jk�D9r���ȃ�J����Q���Z�Q�q2��k�qw�UIt:�A3�y���;�~@�{�d���T��=v�!�R�ߩ�%�;�Z��|nN����0Y�Μ_F-̮He���v���t���v-YR��ٻ(���<��
ᯪ*u;�[/1��s�^>���8�cN��m������ʜx�:���nN�1��t��atw"ӷ2*މ�Y���g�emz�ME~��I� ���rШ����=�ޣ}##�����q�9Zg���t��]�S��{j��	���hM}^����V�2zU?�!q���3�z���Yx}u�wod�wd�a���YB}h�C�6���]��M��S��sZ�p�U�2!�X�i;
����5>�����KHې�{�Eࡑ�W�߯�H�;Z���Kd���c�Ba�WN���z�aE��ﲮ|�)Z]7�;�:T�'�ʜ�~��VG�^���' �ցu�y��^�wMq����n�Ӕ�{Q�����x�#�M��ν�?����o?\�S��l�2=Y�S����*�Zs�I����6�W�l�{P�{m	�����~�S��ΣY���9���L��� ���������]���7���}~���D��r�q�:X�V�<}�a#&`:1���{U��g��v�H�3����3j�r�p숪s���Yu�9�ϕoU9���#o}�!6dd���f}Z�t�>��,�:����D,�Nv�Qr꼆Yw,>���1�ퟴ�x��,�<V�wݪނ����V�n6z���Nn�ȳ�5���]�Ed_.�r�V�)�;iPJJ�j���C+�]�O:�-�����md*G͑N�`5%[�:�Ř�FGuùqiMt9�,�u�a$��(��nTq�"qC�;����-������E��Hd``b��X�ns:FFڼ:/�Pω�2BEGy!�9p<���ؗ�gNǌ׼;~�>8��|F�YFVNPB�A��֏��V��ե5+�r=�ȟ@j�Cc�1f@��l�V;y��CΏ�	���]Oc�r��J=����5�� S9�{*f|�⁙��;�)����6ߖEg�ؐ�Uw�#���pV���_Vd��`�Ww�¯bu�ߔN���c�<�}Q�nt�)����C��<���K}J���5��ņ����*��c��(��*X��u�QAyU�Zv�}.�>��%3W��z�V݃�����~��8�����xx+�'��#��ȉ�(p��@��6�Ok�&i��ʟE{-ov�I(���y+g�s�~4�U�n~K�����j�>~ܩ���^�\h⻴囿i�k�=�}�{(�߉�dd5㞝~w�3_�g՞�zd�ky9�u#��ɧ���&	ʞ{��a�=�}�!�:�N[����<�BT��9�b�a��'�U���,*��|�G�p>:�M!rO����7�_����a��é���Y��=��/1l��+n�������gЖ����Rs:�-����w��P(�ܑ�r�A3wuG\F	Ÿ�$2��M��m����n�}�]u|ou�q4T��7��.���c�a�8~@�V�ν!	��]=]/"/o��-��i�dF�YاW�wP��3+okޡ�˹��m�� ��8���+F|��SY���L;��m��?��>�9Rv�L�K���ƕ�/GH4^)��_x/yX�߷��4������
�K�W�{#�M�>ۿo��3��/�:�k¥E������m�S�l?S�����K T=��TMg=��o������K�}�vES>h����:�	|u�3��νj}%Vٛ��۩�Ήۂj������>Ò�;� p��5�S�yb���Lswp��}~�4<o�C���Ǫ�NB�c��v�%������*���4��}�$>����|n��5Ęƞx� <f�ײ�C���'�R�ʓ�j����~Qm0d�W��O�2`�w�(P�f������8�U�H�"��oir�f�]˟D}��*}�dVW�-@�&��'�T��7����8��8������K��w+Ĭrgaߞ9�W���z�#��##�늶(1BfTjB�7�q\��}�tdQ����Y���f�ʴ���h5��,`�[»Q�+�c�z~4x{�i0���%�.aɭ�`�f�Z\�����3oA�6�����λ;�;�;٭��׫��W^{���R�9���]�0j�C�4�{�.P�y�ԧL������j�=.�5�;%�<s����=�> ǽ�3>�\S�F�7I��q��xz
=yM�ZE^Õ���f�*�df&��3�����L���}3�����x���g=��t�}�+�HL��Ыf���ܵ�liT�k�q�j�=����V�کsȓ���:��ܩ�3����c�T.C�m)9>��Ap�ﯙ�Ni6�Ƴ�.�F��Ͻ��l�M{�C~�t3}^�>���a�Z0� �v���z�^}u�9��T1Ri�Ǧ����It�3���ΟJ�{��ϮO���ג}�Μ�yU�~�� T/@���6������ֳ�ü�z _Y���=37�g�:����σߡz�I�S�vm��B�ta z/���߯{�d�VR�E���۾Axx_�f���	&�(yq���6�J�^8��DevE5aS���F�ь��G=V��RP#���Ϟ���i��t��j��n�0�ǭ�̚�)�r�����H�5�v��[C�1P ���MQ��u^U�:�~���}~���qC������q�6`r�4f.;]΂����iW<�]rj�ԫn��:<��W���K��b�jY�R�C!9b�S"$�mG�nn���r�G�f��/�vH�x�*V�鏢;���&iu-o��;I\�9ձoi� �2��B��ݞEp8��e����[~y[�T�[j9P���2`���xLt���m�69Hͪ�^���|f�=��zX���yO��o���{�#�FxC�x �S�����'e`6����*镳�Y^���"ߴ�NC��������k}��-hr�1)5~�A��?fa�r5,L�\�w�w�b}}| ���w�|�/��Tu��{�d���]IϽv�C��o�vA����U��C��&d��l# G�t��;���oTa���c�\G�;�o�m���O?"���7�9�f}
�¯�TC>_���S����V�2a�㼅�g��P��᜻[��Ǭ�3~;�<��U�o��,[w�0�@���&�n)��t�a*�R�3^ݜY���0�rRxN1(�~~�A�z'����5���7;P�M{D��}q��;w]����u�oq*ɋ-��~��ft�ߓ�eN�T���dw�{zrp���Y� �'j��w����mf�7��ϴA�_��ȳH�.K=&t�ߤǝߎ���υ>���{�'m��G�ǈS4���ܺ�K�:�w��E͎N����z0;s)
�b�b'�&�p7�v�I���#����n��.Є\'f�Ġ��>�]X��krc1�(����2]����4݊@5�6��ݴ��T��oB�|uv���h8�r�@�4 ���,�˾��/i+�;��]"�W�4
K�ݕ�*T�cTڱXs�Kթt}$��΅:�A$��&vkut�Dj�Z�Kz�4\���=��$hPJ�Zqb�}KR�Ы��q|��[#�f�|�1����h<�i��>��Q�]���Gr#N�jQ��%PRV��WU�9�0�U`5[\�M�=&��ZӼw���F�dl	��������e�c=�r���u٩;��Q�����-�'"�XT����2�T�0_Q�jgŮ~X����"hd	f��
گ^�u ͽcP68um�.��%h���ެ�%��9ӝw�Q�F���;��&L��f7��>���^K���휉+2	7�hl|Wt}�������Ŕ�ԗY���qlA��0E��[Mr�b�j�����T�PT�
d{M��#vh�+�� ���F	��vst�%�F$�7�@+siZ�*�2ʁ���h�"e�޲5.f����ܔ0Gdb��IJu3Y]�͋-�OK��\��y{�p�^�E5Sө�evh�!#K��ŉ�b4j�a�J㛟>��V��V�쏕)�k�6@ �J*i�,�ic��q�}|�o7�����}]v@���M�i����]�n��YJ��AwaTDәϋ;'J�{lQ���;��*j�+������2�T��[��Vu��MmGCU�*Hr�d��QX�f����F*��y`���� R붸���k;�[&Xkn��sH�c+�R��x�×&v­NX�����&�C�&N�{Mй�QB�=7QŖ2=�w�H
�7�tI0(�O���!��[�]�үq�J�wS:�5{�E�i�(\���u滵/h*�ݥծmPa��O#\6�X/X&���u���q�H�^�!�y�L���UEY��owD[,�O�x�y�u7z������O_\Wz`n��;����j$�5.c�L5���h��3`���x�+�v��+q��&�A
��ө��L��3mYEYd�xP�7�x
̰�V�Jkg"'�9;���G��Y�־C���e�U���n�u�lꕮc(24����s�u������0�
����v�]f��V\�4d#,.S���2f���aM1�+v=atqN uDe���V<"r{wiNkW�̛F��Ces�~Y{]X�f�}��>saxLL���;��m�WiqB��a=��X��^l�:��|�������mN�oR�!6�jw>Dx���<��4��j����sBf��e���x�#��ɜ���mn�t�gv[�$��_9ϓ���4h7 L�z�_up��(�����8��2�5Z�j�l��#�X]o/�v�6�G��^vJ!��(��#6�A$X̡Dc""F��c\Kp0PUE�aE�DQYr�DLB���8�`�TJ�"�*��`�QX��\�Q�B�X�1�+X"B嘪*��U�����[imV(��R��Ȉ媂��VŊ,Q�l�DT�hJ�mQA�H�A`.\\�JԴ��Q�"1r�����j[QH���QŢ�TQ�X���	Z��1Z)�m��QH���p�*lB�V����X�ZةP�(1Kh"��Y�(�V�A�r�`��� �Y�[u�A��iF*1��YmQ�Q�"!mAҥUU�EQ+�&&�e���mJ�
��Q�)n��V�V%+hVʍ*�T̨Q-Ƣ,A�keh��RТ��K�QE����Kh"T����q�B�����P�U�f5imDYZ����EUR�YP�RԴ�[[�`�J�[MaDUR�2��[JD�m�*�J�U��*X� ��T�,T`��t�E�'�|{w��O>��-�!ɰ��;�I��*��]1Յ\yu����8�ɝ�)�� ��B�:�;I�kg���M������ �9ʖd��&��Fĭft?��Y����樻��i%lu�+���>�����֢1��p�=
��`�"�^�N'W�Ǖ:���=���>��V���*nq@�$7���KW���m,ߑÍ/	a-��pe��ܦ%���d�O&I��<˜���V�r+��=�x�V�(gdƪ��]�3V
�Lצ���|'������D�,�ܑL�s���V����'#}�=���^�>23�$v�� =��+�.�զ[R�-�v�1�ݾS苪�2�\RYsϽ����5Ǎ����s�6+(�ϧ( ���-���}��$-ZLZ�]�@�P�j;��)x+Wp<[g"��o=�c·��>#ܪ�I��)L�E��B�Q���ҩ,����D��� �?Z���Ĝ���Y��bC�o�ឯ�b��pn6t{�'jg��E�N��~C��Ũ��!�2�S�s�.��5jHBv��0��F��b��&�z#��b���Q�2#��Dm{韔!5=0��(��o�y�x΍˨�l�؝{y��o�����;�97��wLk���di]z�*F�On/��OțB�/:��(;�А�I\.y��b{DM1CL֗U<�+���P��,\�P�ҏT]y�b���$G/2w
�$����ǈᇈlTcqe��ջn<�����A:$W4I\o��9�A^ʞ�^Y�s��,��O��r�GP�m��P1��Tm|i�.:,N�zO��i���Tɬ*���y<���S�n��½2}�dt����H�T�4��1S�S9~�����1'���պ6�c���p�^9�~utk�������(c�&{����!����!)Z$:��\H�D`��Y�d_S#�wЕ22#NvB���G?TϨ�Z~~��l�e2�-
�#�3�OnN!��a���g��at=7?�:��Z�v�#N,�j�N��
.���`[�#؄y�E�Df@?���=6�`3ᵾ����童�]m���W�i�~�l�{�5�[��׮gȣ��������>�l���(E���C�K0�����3�QN~G�����M��q���5�3��/�7����o�����߭ڞ#b��Ϲu���%�*��y>��uxK%�.�S�t'fuP��IoLA�ۤ^.n1���~{�S�[�eFO���g{�̞���{�e0����Q��0�8�c����O��6#Ƈ����~T}q��6�XY��7uzk6��.��Z����$�-������h9�G\6�yy��a!T��]��lt]k/>]VS�sWg��*��4�1C�`<�:P��;N��e��KK���2���e��}����u�`�hP#5n7*P�4����(5�GZ|t)�{����{�[��e�e/�|RY�!�>��!��߫�SP�\�4��3�<���5x{�)^ ����&��Π��[N���O�"~�
0GxVA�s�s�>�x{�����[���k�jw�7�g����4;ʇ���i��A׍Bjx"{�A+���?G�=,��f='=Xs���V�o��/J���ϱI���㝏W����3�w�(��_�)�)�����Ρ1�������f��Y�=[�����Q.�5�;&!�<s��@yǅt�������o�)[�p��g��������WUg�EOx`4$#N�Ūh؂��y9���5�����H��_�d�~�����;٫�^�x�Khv����_��^^&E.���ף��-�����d5��~y�:gh���K�����Xיc�@���d�b<.��#�T�t�'>�V�ȋ�ç>�g=9�M�+m3pG�@���=��;�����?y<�#{ދ��W�A����a�Z0� �'j���yu�&*�!2.�g��wק��/�n���4��NgO�c��v6���>>��{�fN:��T14�)@��2��)wl]�ṫt2��hva���������s!2;,Ц��R�Q���O\�D�U�ᮢ2�n|��;5���|��Z����MvK����u���	��{�R-�H����Ʒa��vLǣ8=����;2��ֲ�nur�M$��W;��w	�[#}�=37�垝�w�,S�w�/^I ��J�ͺ��ôؒ���'��� b�@�Z,q콻���o�-��Ʀ�HA7ACˍF��jVG�S7Q�(��ǜݾ���G:�#) ����Q�Y�2"�8�1�b>�>������a�pG�2b�KL5�l�(�q�o�,�;���i��ӟg��T��������=~���{��恎&��p�#0����l�z�z
�����y�x�ZB����t$�9�����Jׅg�BB᳞�o��j3��EW5�>�zL�yO��o�6<{�#�Eo�8��< Rȥ#�����}2v�h��� ��;��'���[���_��j}Oײ|����yX��u����Ȝ���8y���=�ޝ=�W��������M6� /��wg�"�=~Z�G����z̐=ު��W�9��G��s<�׺�u[2�Xt&��2 ���K��3�߭��U�{�u/�T��Y��B�53~2��~E���|��a�^[ǡ�<f�մ��U?��~~�0��x�����;g ۔�]r%��9ق����p�3��U�طhr�Es�� �ڹ�o����A�৷��^��u}�O�X�t3.��LSU�tOWc돨Ӣi�E.Y;�rajB���Gd��m��~Υ�zK����p��f//Nv��l�Q�S^��E������X��#����]��G��)��o<�ئ�y챆�{{�[�My`��zļ~YP����*G������c�P���Kd�g&��,ßo��3q��;�壹�9{��Z��0�����Η;	�2�"5���^���߳E����]E���/�����y��9�M�����M{�{"��
C�x���I��9���;��s�υ=��� �{j�u�qq7��7�x��5���^�~T��>Cu����A�5���,��S��|�9����BL��v����7�*V�G�o��S�C4פp�x6�����uK�!�8���#�|�=uR*��{��}rȚ��`z=��-���%����Ĵo��;uIxc	A���t�?r�9�<�2hխ~Z<��-��l����FB��H؋���mdq��,FDr�.|G��F�w2��a���7�f'����*;̏DY7(=#ג�{�����[��������h�"ʤ;� NF��e�����K�{иz Q������Yˀ��KralO�������x؟��s�6+(ʦjrʶ�p����b�u@bu�8}^�u�+���\̕.�t�x9�ª�;ʕѰ��̀�%j{V$��wQ�� ��O���kx��kS�5��to:w^��-<Ṏ���m�l�9q��׺���o�jqԳљ�8��L�'7��t΄��|)|�e�t�6�zd/�[ڊ�o=�c·��>"���L;��&s�5�_D�Tߝٕ�0Z���f�%����l=���ICm�dW�֐YdgeJ�{
�������({p&<�=��9_D�"�����}(ǡ�ҫڡ���1�Q��F�~3���b����(kb��9�g��8��U���q�]�T�����bk�ʮP��"�Vu��V��(�և)~�����<�z\�yX�z��I��H�gΜ��9C��@�f���a⺳({/9T�,�����e�{Ƴ`���<�	���̩��w�=���9�ٗ���H�{Թ��F����GG�N��މ>cۀ�v��0o~'!��׎zv��~��R���${�2�k&7܈��5��g\_eNyO����n������[+/��3��dyJ�s����'vb��Ǹ$��2K�\��l��5�Tg���5��E׶\��{���M��+�Y ��i�S�F�=��:ty"�o*�^��E:�p���Y�g�p9~��Fxc���ʈ���r0�W��ȟ��.(�d��xU7?õם��E�Ϳe4j�<H�z���$���
*�\8!d�b�V� VPπg�9V���αn_[���q�e֙��]u��N�9 ��N�w����ً����C�jWv��yέc�:C#��2�R�n�]]:��*+7����i��;�cӴ��}#���ޫ��}���ۮ������.�'�WO]���W�"����L��O�N�m�=#o����O����G.�#���--���x��ۇ���|�x�� �j=���Ϭ��o`���݉?>���[�=�b�J����1~����")P>��?cC�Ujat����J��X� l8�`���Cؓ��������{T��./�q;k�ĸ+k���V�ٕ�H����T�cʡ��T�zwXc>��&������޻�Z<�+3޶9 ���hx�r�gEk$d�Lϗ
s5��^�E6�x�\ߎ���/y�W#;~�=���w�SӾg���*}��Evz�q`1�()\
�X��~�����U���7�4�ֽG<ӡ>
��t1��3�Rg}~x��M�y{ֈ�\W���\C�/�&d؏xh�K3i�LJ�Mx�*�c,אg��qϚʝ��~x��Ԁ�����̼��&���
���E{�U^ȑR����x߬dZ��͂�����0��P��\禥!/�F�XT�U��=�י]�+9Έ�\郘�s;k���ep�uչ�p<��e�� N��Z��+%���hүJ�V�w���e�,;sw�5I�]��:$��ܶ�pz���b㷔�����3�>���0�v�n���w�U�(��I�nk$}�;�H{�3��	��\(������Z�"���^��U22����9wz{�|{�0���=�*,
��d��T��D,A���8��Qy�ņ�8��4�p��^*緽\||�.������I��(��PϷ��r=��{�hψ�
�v�����J��=on�o��W�G�
}k��t�s��4�t�w�;���}r}O���A��c�k�NhTǀo��w��z���vy�~�>��h�V� �W�;c�9���|�ӱN���~��N�$�}Ԧ��B����˺U���������\v@���W�۾A�~�nfn55�s�T���<��k��~o�7'�����3�1#�����~���]@��^OdU=B߯�hQ'�#U藑������exs�iZ6vW����=�g�b��8�ޚ�9�: ��O�ih�r���X^S�=->�������|cu�QƜ��Z	��<�-�)8)`H��
s5<���J��74s|��r�-`�Fv�c"߯&��g���yO��x������<vo�<���� ,S�f��d���:v�>��!}&��b��y�����p�.�k|/�z����2�Y���j��%{���P�g% 0s/�<S��w�c�v���V�^�Dt���.$�e���9��T�!�����x����4 ���Nwh�ۑ8��bD�|�'�8�O�'e�6��}QA$r\j������ci�V�yp=��i���=o�Ӿf��򡠯u����4�!Hύ��Q����O���p*M|<쁆�x>�w|�-}���3�!�޳$�~N�W��gb��a[�;�5]5���G"Kp~HІ�J�/��������Ǟz1O�ҥy��k��`Dղ<��3>�\�hd��Bj��M�h=��:���y�G�}�^O���c�~���z������]�=`58L��3�MlJ���e5�)5�r��xＰ��-%�z3�[#!�X�c�̡���
��=�5{E �7��N����ݾ�v8�2��+=� '���7�3`�����:\�~̩ȇ޹�׼=28�������u#h��e����=���7ӵY��p��[��Z��ЖzL齿I����ls�υ=�f� q썌��/ї��7�>Y�S�x������7���O��r���g�i������ܟ:�.�Q3\�ΧG��^k.�nV2�(�NG��|6Y���#.�x�����fu!��Mw�����_:1��E��O��8�ݺl���w*$Qޮaw\�߄T[��u��W��\�*��6ug������qr�tN���5�C]^���ǪSh�x��J�Z�(�}���X�]��H;
��`g#3�Ή�nJ)M��^/Gz�Z����ao����(dpȖߑÎ��A-�~��Xe�o�*���a�o�h/N� ɍv�{���zF�~������X���Df �
s�Z���T�7{�z��y.��S��2,���z�^�=����z��ǽo�l_�O���"�Gn��tT7�EyjL��'}�,�(Ԩr�zb>�Bv�.��#���������b|_�ϸb��D{���j~��2'����s�j)�jK����NNYy�#�l�V|��o�t<�׀~��Xz �^��ɉʙ��&�r�s,�*���I��a2cŹ��+�j9�ICbߖEG�ϟFffoƑ��|8@���#����[:�(�Aw�^�5Mّ�S�s��J~V��Ϳfm�̙�a���ߝ���8��U���F��?(2�S��;(�\O��]��q��I�4����������ʞ�5��>V<z������x�D�vG�X�^����]���,m����v:��5��W�e`�9	݉�ik���\���<_섒$��	$I?��$��	$I,�$$���$���H�HI BI�0�@�����$��	$I���$��	$I?�$�!$�$�!$�$�	'�$�!$�p�@����IO�	$I?�$�!$���@�����$��$�	'�����)��X�����0(���1 }�^R"�R:�4�J�*���R����R����2UM�	T��5V�֖�P*�V�$**��͘�%*E4h[h$�26�M�m�ƕ�L�ٍ��mb����)I,�Y�e�l�J�dHhڵ��Lmm6$�;���d[f�ֶ�YMm�cU�z�K�Z�J
��Z������h��œ[m�f�kd���6�6ʶ	Zm�d�4)K6�e�=�G)6����S*i1�SMj�eVZ�ln���]���Vm�  �q���e�.�<{b�v��e�2#�պ{=y��m�e]�xuUL���7�O*QNs�{`)�[�ۀUS�;{� �OO{�]��z�{isյv�Ͷe���׾  -�wT��5W���j���@]���Q�_(��\z(��( ���^�:4QEh�s��
 gWF�  ί��
 QEw��(���QD���-Z�m,��U�}�;V��� 0�>��{U�@Ѷ��y�5n�uC��v󚧢���t�Ъ�n��8������W�i�S����`���"�����^j�ٱmQ)�� ƣ���[�ٹ��F���c�+J�k��tj�y�:5]nռz�^�h�i�.�حk�owyk�Z[]�ӵc��tr�۷o[�$��h�{��l³-E5�k��v3k+� }r6λ���;"�m*�]ϫ��ښ�뭧��n��k�t�
�Kz��'���v�n����M��ڍ]ǯ{X�^նRʽ�y 5��[�{hR�ۺ�9�i�L�0�J�ڳ�P�� ����ҫm�����w�K�w;���-v�m�f�����J�֍U��o�k[m5���Ss����h���݃p�4������Q��*ܧ��me��=gzz�Kl���4���mݪ��_  w�}]�k��K�oIG�QSΛ���ݺ�s���f�����H��(�4�n���3Ow���M'm7s^��k���*]�ջ�o\���K^�x��k�j�OZ�L�hf�L���l�� �����Z�n�]�����n�Wv=��k�����xS�r[�������й����V��n���Qz[6���+שMV����q�mUm�c=�s��a͋�g�f��G��5m��w;�Q�  >v�.��ڦ[�ӷ���ڝ�w{ �U^�z�X�����-��gVۻvԸ��۸V
;�U����9ӽs�y�nw��Z����w�^ͳi�V5�I&����   >緧C}�w@���uC�{m'n�/^�[�(�]n�]۪V�WN�ys�ֵn�nu���a��-��xڽ�V��jz�=kѪnu=7�v6n�h�]�rں����4��JR   �{FR�� �j��&������  "��	T��  ���eT�   B��2�j��6�M<S�����~�����'�zn��?Q��N�e�Fh�S�a=4�����_W�}_U}��?�_W�"
�T@QO�Q�"�
�tVES���������е ��0���Й�x���@���xE  ��*�٥<(�4q�lMk[���Qb�TIJ��d1VƆ��˺�Ҕ@y[�ʈb����W�d���/@qnb܂ڨJs�I�Aǌ�TJ8���{Ij���A�p�+V]�6���c�0���{gV�TC���2��VQ�쁵�pv��X-�7`��2�cKꎍ`M����m����܂��2��H�ʲl�������e�nV�-M�ic1����v�<���@֍y`�V�*�b�9����k����Op���"#Y-�݅v��vR�H���f���
��EDjM��5-�xB���^���ԍ�!�+)�#�����*7bP�dL�N !N�E1�S�[FM
���p���,�����XΠ�V&҄����rb;�FEZ����/*���yCF�&�l*�:�,���e��@	�ƃ��7F)b�lol��j26��N��n��c��	��]6>R�`ۻ�׸��[����G ��PN�Ǩ�H�`P�d��^�5!��f�3f)v��e��6P*���K��n˴��K����R��P�vBa3Ƚ�fb[���6!�G�Q4�[��v�#un��ԭW[�^n��+vc���1:�[!P+m�jF�B�릶��7�V�*Pm�*C�������g�Һ[b�b4�ML��Y�Y�y�i�$݈Hn��V�[Ī�֢��bQU�Y�-^4�h�6j�S��h�A&��\J�B����+����*v;�칗�E�4j�ټ����8Bek��R��snR��:��Ƥ�Z�]�ժ��=GKY��[�w`�X)Q�q'W����� ��b��K��X�)�2�_�KQ�G��ȶR��n
�x�Q�f�fm�BBݓR��6Յ�d:��R�A��I�2ˈ�(�"�1f�@\,Ԁ���éPЅYJ���Mxll8��ٺ�`;��r[CscĔvv$Պd�v�9Fޝ��\O.bT����*�ɶ�-TʤPu���ɇ�&^���肅9)b�xK*�8��0��0В^��Xś�!��]��Wc$��1�pc���&E{�Kc' 30��1�mM V�V��[�e�j�ј���݈+2��裁�ӊkY�!q�bcYBnB��[�J3�!&S�桉)����
b��J��hӔ����Jv+h�od4p9PV�[�%�[��Y*"Mո��7%#Rl�aR�%<����R��efe�VҺ@��j��z
HO�c�Z�8r�ޘZ�E/�`z���*Yuy�D�����{Hn�����)R�6�f齢��t���FA)�h*ǢL��yF��Tsc��T.�E������3K��Q<sD�v�
��k1�d��Rʧ:��JX64eI�Xkj��:����M��������9�6p];�Qb�E�!tS�����A*x�kJ�cI����d��Z�"e[Pb�Y��k5eՊ�a��I��,E,)���C)��T�6�ӌ-Ot�lL�sr��D�U��&�β�T��0�0�X��Ew0�YnU���t��F˛`�ׇ��&��G]n@���6]ŀc�(n\gU(E*�2�Xv�izK���/0��e�(VZ��J��Ҡk-eY.4雒�6p-b�X,��lͣ+*�#��4a}on�h_d��ځ�m|m���b���Cp�5#kpMU�������R����Ʋ���M�RXjMUi]��VoD��\�b���z7nP��1aX��rb�Y��/Aj�Im[�,�4+R��S�DB�ʪ��d@v㥘����S8�c`zU�֖��*B�0��^�ӱD9�욽���jH �p��E��;E+�
K�Hr����fe�^f���h�;���&a�H�Njԭ�����e�
��>;-�J��^�mpJ��6���!ję���Z����Q]�bt�ZrrK�u1���X�"�i��R�]5NX�*��u��q'2�JeB��reͩ��h����qj�Ѯ\y�N��,����i�����cr����1hD�U��Xԡq��l�`�Z�J%`�����.�MĢ��7W˨�i����6o*�(�<[&�B�S��Ss]n�xu���HK�S-�����㱟>�X�x���LHF[��22љA�3r4���8��\5�eӹ(%Y�������UwAIK�STn:�I�����Hn\��*Q�)e�E��gNE��mJ�Ahe��bA#g1Z0T����}�	�����\m8T4@�c���lk{���B��F!%�d�;m=YCD 1Z^�o[��rJ������vh�.�bX	9�1�g��oB�˭:�c�.�9�F����L��od 7 ��-6�G��\�ѻ�,V���Qj�!7kJF9�A�Ь���P��a�rUm�B6S#.�X3F��-i,EcCl^��gl,�%�XQ4)=Fb;Nkt���b��ǈ�BL��[�Z)P�#![۩�1 6زw0��+\�m�(řYa���{��T@̦֍XL�y�
�#iԨ<�KmU���qC�5;�Z$fE���O��f��nh��(���A���8��B�4[ոtkr��2*�Lmɵ jõ���n�EH�'f̡�\˭6ڻ�����p�%�+����!Sˠ�����PY@Sߋ��xn7����VGZ�р$��\�&�Z�U�/C�GS{�/�{A<���� �Ked��*���3Fm2)�c	4ʋP�40JA��j�oe
n�y�4�X�r��hpQ5�3Vɻ�[��YZ,nf01e.��)�
J:2�Ê����)SC��O��(�t��Ke�Q ���B��&n��&۔p��}��Q5mM�H �r�fVٻ�X��72�
rT�ڹ,	�-(m,�"���ࡂp�=Ĩ�o�c)��5��呙����!��7V��Z,�r��إ���5�J�{tT�\�Q�֕�LǻE5�X�Ks�(�3��`����ni-�s2JW��c�J��CXQ��8,�ιf#�3u�5�u��q�4��a^�^̐�j����=�$����be��,y�5��y��Q��Vїt{���$��b���V��`M;�*����ծ*�w)B%�nH2�aZ�H����h���ڎ��r��]���hd,Z ���S��J*����t �YL�V�iݺz.
�f��J����(+��"��HL��@t�/b����t��Kf�Q:*`�6�6��������;����[�u��{�'�I��/����T�����j�k�����i�)PS���ʛq�0�c��Qe�ɳ�ֽB�K��W�<wM]���S*���2�S�ѵ��.&)1+Z�uxs(֘�!��m�	"8�Hob��4C��BEFk���-��I$!aL�yqZ`�<�Tm	a����X`;ݛ��v��x����z��+hʻ̤��2`oR���Hj�Y7R�m\E2�|26�U�4�,�3�$�ʣ�U9��F��d )S[��3��W�\�v�ф]-�%�+5\ �y[�֪��"��2��R:�7Кs�w�%�U��>r�ՈR�1�:(����ݺl�����v�%�C%E�nٽ�̀V4$��R��L�*��U,J"�0^�̬¯c@{A��+V ��ѳwLY��K-"�(���*���%�GH�����U�[m�z2�M�-lZ�,U���T�)�:ې�okIi�K>�ѓLe�/6򅒂b��c)mK*���4ٚ/�w:
�Z-�Rj��Ӛ����/	����O��9 ��s��r�ݒ��3�I9e� �w��d
�	lST��n����iKa�[&�q���ViM���.�IzY�YDi�&�@[{B7H<��awI��(�S슱����nfǬ/Iil�9rG.l&��t.dR�Q�X�.U����4��XE.5o���b���[�"��x��%^	�Sޑ��q�+�8��`p2���b�y@Jo+u(n��YX�����DԺv�'�ii��j&)�zv�'-�ףd��z��u�" `a�:��]���č����^��L�����Ь�1�f���Lkb�N��J�4�&��U��*J�����V鲦ֹU65��.ޥ�9H �Yl�	�Yk(k����c �Ǚ��ȣf�b�j*4�jĖ���&c�Co�ֹ�ۇC\�
�澟6�w���sdB���E%�f���T�b鿱�R�����u8�5)hMiZ��VmJ¢!�LB�Ef�⒰>��ˤ�(t�{��JSn�
���H\˨d�G2P�ff�7(K�f��HD��"�)x��+oNX�[h�e�E��Mb;i:L��#l\�thՌ��66�,��kkJ�^��J�����H�<"ְ��F�8ڳ�1��/5� �0Yi��Ш�l�,��I�.�[	b��lK6^�������L\�nS�Bv�C-Z���l��"�蛦�h�d�B�}��#t�`I�u�U�Ȝ��ڙX�<˕�)E�D�eLiU�WsYi�RZ0�F�i�^Hs�HVL�e�{����R�P4dM	&V��*J �X��b�d�m��d�fűn�8�Z��;�(Iw�7`�뽈R�X�t�N���Ŧ���
� W%���7���K)�n<��h�1��3PY�Xϥ�B��6
�'�� ���J�rk�ކR���j^�Bf�&���`Tާ� �s�j��{v�ml��bՒ�)ef���{IMFi�ZT���`v�u�­��m��Ԗ�X荻l���a���6����uV$"�5��n��tԩ�d-��WWM�J{�E����j�����
�򏧼i�?Y���/���������D���������ʮA��hQ&��B�MW����&ҫ�w�	6Y�bX�ߵd����iM�Y�SH6F��Ұn+3j�;0^��,s0�q�b�6�jK�������b�+TU{��-`���Xd�ua�X�sm;�E�� "÷��3n���5"�ڲ�#2#@+T��'�b�Hk.��u�ن�7�a`G�f�qӫ�f�,=5QX6��5�-#�!�C��f��������/4�5x���&����y��zL�F������ɥ|�ݬpKqb�*Ax"��m`y��i��h�!V�Kh�2`P<�`GtTY+	�^�`�/r�O���������nh�L�-����n�g([�cmT�@`0���7�\H���㕷[���� ���(m/��O�7)��cA�� ����v�Ҩ�����̹��SjU�ݤ�F��1�w�&�����*,����{�"�q,�܏A��X֊29J���J�v�kD.ݝ�坴��ۗ/7Rt)`�6�V�ed�5�����S�1��:����a+B#���(��c.���e�i8�fP+Ŵ쪶�F�h8෺�۳b��j�h�������x��Z5�e]�,f�)�+,\c`��4.��J��u֬o$���̷�!�fJ�Xr�Ђi7�R�uv��
�4��,$kJ3B���@�����=��Tq���d)�z.�M��L�ux��c)��
�'�N��S�!t� �)㳮�֝[t��)��7X
�Z�y&�����*,�vo�����6W��aj�c�P�M�~��h� �3a;�-�W�є��A��i��a�pQŪk�V�f�����eX���4bB�Bb�+T�f�mө����'?f�l�ڳ�jőS)��-�Ʊ���!�e7 ЩV	�$f�B�Z<l�x�E�	_)p�_+�Cl	(;؉�av
i�0�޽R��+/qQzBm�2;�/ :�r���6K��ޤYL��P{#��cGԡ(@��z�ŋYx��n���#E6�O&�[��u�2���"*��h�"�.�I˫o@t;Kl��\�K�i`��V�ŏ�M��Q�u�w� � j! j�t�
�0�V�{�3{�Oop�fE1IL��+�ͣ��HӼ�.ʺl��Bk8�^�@�YӁ!>��)����۷ux��B�53k>F�z ���tl.bA�����H�:)(q�Vd�ZV��f�Q%[�\��p�պ�, �-+�2%��՚M���=T�L����;N��ܶ)L�AN1Y�F'cS�sN�ˆJe
HS��[����T���IL,Jf�&mAL�f�ѴR��1�[�����f���y�F\MjqN��	#{VL��԰�m������ȨLNP�ķt�f��1ZU�E/�f!XU:���mY\1[$eZ��w��u��.���&гd�X�f��Z�h�3��SE=F��R�k.e�sQ�%d���Q�/2�Ѝ��+:xr$Ȑ�H*�k#�(]ٖ�ܣq��h��^��`�I(-X�C�u���
�F����j�N=�)�$P�yM�<��6�&�8��� V��E�q�L�ɹ&�eYq9���X�u�.՘�(Z��k���dWtܚ�iA+m��� e�M���9��P��U,J�e��r�NcKq��+�(���)LV�ur[���Y��߶ԥ�(L]j�BB����ږ,-����{�^��	��n�5����9rA%[H\ҵ{�è��dj�.��¼n�[Q;�S�] �+C��m�a�G)n9cEf�Q�F�!��:��nJ�q
,�K��$&�sN����^/E�u	�Ĕ~{�'�r�u�+��1���η��$�e�mK��|��p7`��.��[�ĝmc�F����Ӄ�@��P����fWF�.�5!�0���_*d�=J�i��x�U�p; �_eΞ�ӕ�� ����׹!�ef2-T&��#Ҵ�Q�٭=b h.�J�M�|i|0�ק��&�ǿ��zQ��L'%�EFY�Gf�ٴ��x�MY������+s.4o3�s17���r���(�C�L�GcdQ�A��};���&�+K6r�תf^�M����'��8�h�\�;���ll���Ke�� =�@��d�h�����/ZǮ�4�\(���6WH�m%���~1=L�}DL���t.�b7��/_76��n�R��V��5%n�5>�Zh��Dj�G';�i���2Lb����Cg7�$H3���xj㾵�MR�Of���N�"�����N/k���
w,ڌ�v�gX�Xv�����^oS����c�5��z�s�w��6&ڰ���^�!�u���:�Ʈd�Թ�@^�U� ҸZ�O��֍n�u�g9Nu�?.��n��c:]��Sn�A��;Tїcd��o�4��aU�/��Ϻz��Y�^c��Ϥ�MY��
�l8_v��\��r��m���Yy�~�-�t�f;K�u���2�oB�=uӷ��ɺ9�TC�sO�X�d{���yf�4��[�\�C]m£z�m���"u^a���}Y�(�l輋���"���*��'m+]A�an�W�j�ͺ�h�0.nNn�7lRt�u�'3�w�R������퉉wݗh����������7vz��6�N�zS�u� Ҍ�Ю�p�;u5`�j��m�G��v���j�64oWb�D���h�ؼ���oJ���x�4�x�Հ�6�2ɭá��u�e�y��;3�9J�,<����{8&��h�@�>��	��Z�rӀ��][��Eh���{9�V��)�P|�3��`�{l���z$�VmZ����l�w�Ï(%Z�n�m̻��	���U܏�j7]4��[��j�$�Q����e�R�N���i�Z����S���;�ZY�M��&���y2�ӹP[7`���]�ʦ�n4M3���g%v�fZ��ud�:mF��Kt1����6��{��q.���p��{z[jI���áQ�]i�^?0���b��=�U�h�<���Za�,��B[��h��CJ�mы7{9ص@k6;L�)��0/vZ��8�X���"��贸W1[�u���Z�KDUT��+�(ثd���e:��Q�۴q�P��U�
g��Fc�˱gj/�6�i' ���0�u3�����~�>����*�9���[���k�3�N��*������㏸d5����G�Wv�9V��ͱ�ѱ'MJ멋-��y�7�;�yw�Ā��tֻ��s��$n�)�wdw�uZ�B8�ۮE�� ��y�A�yS(ڪ
��JҨT�޸�S��=&�̱,H�� ���B�$(�P(ך́��7ҌA�jK�G�.�!L�-�昶�[z����6Gsϻf���7m^7�QiN�2���=�"x���x�1�P��ܱm���v��q֠�>��ֵ�����w���BW�_4�����vh�G>�1��F�/i]~���ۓۆD�lsS�����x��)���X��4<���W�}H��]�O}�K����J���Ull�8�����:��������͜�@}x��]���|&��m�^��;;R-֮�q�s�g`��ȓ	�M�6c~�X��:�b���X���bۺw�D��gk�:������<��2�����Y��p�;&!wA��7gM^n��siQL�u��ig7�\܎I��Q��٫�ѧ��5I�vf;���i�����MYz�b�6��&��z����	X��ߢ��ݔ\{��1��κ����rqq �Y����lg)]�j���,ン��]�;�^��%�t���N�����KŃ�6i�1�������δ*n�q�{E0�Rd*�������FP\��H�y,wLr�뷒�Tģ\�]�Y��V)��N��{��Dd��;[wq��9�Q�}vLt-��3�6[5�����wH�;ً�с�����{�oc}�I��}@5�+OV=�����0��h1�Mi����ٙgx�|X��]���8�`��;$�*�+���&c�������jZo@�G�;�N`9�cLܺy�p�B�8�����<{F�db�e*�y-�φ������&yޖ�+>�'��.�k$�V;1>��SF0���,Ddk��w��[��ݶg�Z�@b�wT�ǖ,���ui�j�8�?vn��f
��]�i���Ӧg�na��HU�P�=�H�z
�� ��mm:�2m'[��z\$�E��]*Tm��&��I�t�ƔC;-����m���G�xb�0�T���܋���ۖJ�A���Y���GaJɇ��r��v�؇��,M���Y�w�EA�d��ljh�ǅ�ݐ�����!w�6�Gm:h��u��:G��8t�i	�	ov��[+����n�Z:�έ��������F�ږ�>n<ˇ5���[j�ޜf��L�T9P�jsOUť>�����Y����wªfmd��=޽J����f�Z�Xu:�n�m�2b���FQkh�:.�N�w��c%=�v+�yk/�.�M"��w�Ah�F%r�����w���<Li7s�ɏ�����#��5��{���H�k�]��޻ w)qA@����F�'��u}�F��"؜�E�{ݑ���*��s%�gY�D7m�Zi:�U֡�k�s;kYm�bLCD�o5ކB;�++Q����3e���q����l<�id#��:�S^��\��T�5۝{�.V��{�W.�����i{tU� Znt�Z)���{S����P�Ӱ<��n"�)��K=�L���\�v�:e_h$M���7�Yewh@��ޞ�Z" <l;F	Ds3���F��X����m;CqTQ���hqLЗ��&cO�Ɗ{��]2�]m���=���*�E��L��N;@-���o-A׸�Q( �����4s�f�u�P��$�o+\)V��[�կ��#*��{�DVT��*r7�����P��{�_���Ř�]p���9�rR�s��;q����
�mһ2�HK.f��61ب�ּ�I��f�c�/#5�Bi��CO�]ԩ]��}V4��56�(�y$�ض8�0���6�1.�k���>땗��&Juף>{�%��v��g_�5st4�S3�,U�wLg<V���A'�F�WZ�i8�1Gu{OOZ^f�mNN$�1xu�L�Hv�l�s��6�J�|F��7-v;䝼�C`�X�޶���27]�T���d���3������j�z_����w>-�m汆���{93�5v�K�[���E��%YOo��4�Z�P
;�e�8��]���X�2��Oh.�`8	��\w+�`�"_�����T��f�S5��q&�t�{[�pń�@�g�4��7��O�} ���3D�`{	���u7ltn��w[��X�Gú�a�
��-���_�_ʛ��I8�lO�gl�vڥ"�l�rU�{��=$�|�ɉ�r�qgj
QuI1�	'ؠ>���Y��թ��V!�g��V2�H3�s�,�-���k��φn���qČT{
J��X��F�C��@j\ ���i�e_#J��:t��3i��cT7"WN��V5�'N��ɹu��}�G��2%�<��,�]ut7&�Y���{u�6M����+�04kڷ�!�����o@Gr��u�9h/Q�>.�;��n�ںs��v�,o7�n$6J���P,Z��Ӎ�Iu$C.ޜ^�tJ�[-8UfShoJ��Ekt�dd�:M�[��)#��]e[P3&�o۽�H	�Y�w[/�F��]o����8��u,�LZ�R=	_b��?#�V^��uE�RfK�Y磕�h���v��6�մv���	j�f&Mk����X+���J�s$�TT�#Rޠ�dN�2�a���b�T����u��}i�YnHx=�7�J��)׍1y����;����=�N`��e���01����8�V���׹wT�����W)��[�oHi��*�G��\�*c	��� T�j��uL���M���˙%3Z7z���T�ݶ��b��Hũ͵��~��֝�8[�8��_YCe33��b�ѵ���	{� ���=��6N�uKg�_�`8�ך�*�m�z�����y�A�/�3�Y�ݍ�W!^j^{�IY�͈{�"�;$�r�1�_��3��ݻ���P�D�A<���ŕ +�d�T�An�	�y�K��Vl����d���k���.:ǻm"w�dǾQ�C�����+uJ��|Ic���ú dk�M��5e�
�WE�W�n�j�-��c[�wj9�n�Bj))<����B�
wQuh ucǬ<ʻ�+�ST�ҋ���gf�i�m�XK,��#7.�kd��������u��+v�V��Eۦo��gV��c���9�m��"�o#8|� K��E'1~�KaýڪW:��<P�8K�,iN�G�D��|#'I��%�\XRTwkf.�ܲi��{
����ρ��\�jNW�tƗ�.�K�������cT�wN���̛p�0��"G�!��/5/���*{��w�:�6��[�fN�Ht�q`f�*9V��/�-�fe-<�U˙u!h������.%l�.��]t?=�s�-ly!��
$��\��.,�^�	J�]N�;�fMI���9K�۫�&s��nh;JP֮k�]���Qj��Vp���{�@OAY�rT��9����!GaZ���U��H<2~�B#��I)���^͋�f��ͼ5:e�<�{9���op�����(�$IEXZz�i����[���ڶ����9&�z�*R�}�mj�`3}�A���OY/�j��즰�!Zܝ�W�	�c7E3� �X�����e{r��p�zX&ʽ�ElP��\�: �`y��K�KK�v�`�c�T'�4<� ���������~���ܷVu�J�W  XΉ�r0oa�~�ǴuK��r�]1FgYq2��k��&�gf5�/��z�qِ��<�q�j�wl��n�K��[�%�7����z'�E�n��>�����#��e�F{.6�"��|VǖV�6d|��,��]F���^�6�r��aGm�m��v*-�=��e����´�L���y6��u�y��f΂��]���Tdv��WU֍�I�P�'�1�%]��⠆T��8;��6�,�eK O�w�{ksw�݇8+���h���(�njM�4:
;��{],b{:�R���0\]�{[X�A��\��e�2*ߦ���:�X�����VSՐ�4c{�S0���pՋ��Vr;)���7�-VH�^�$����hwL��*�����H�*��A?��<nf�]������e��ˑ�qgD2�sA �R�����f1m�I�h%����=�.tx�v�)��!���_f:�����n����G&/I6e��-��!}��c8'\�2��Wn���x�j�hI�83w ��Tx�-��͗�(րďz�H�3�-��g%�н���WW.�ֳ5ڽ�ި����G2�F\	xU��<��v�6�[�r�3�}���(�mK��!�/���2�7{J����yob�����,��Es=��o�Ӫ����5��:�..�wS�nNGv\Ў��>�V�f x�G�k��3�s���HkV���}z}�Orչ6�p��h�S���U�����ym'���6P}�����pyJT��H�w��0�U�/�ܻη��Y��nmqk<wj�us]�������ɸ��P���@�����o:���]-���^���);w�h�w;;s(�H�oഛ�bU.�2�]D�:x��KWA�ڰd�p dHQ��e��B�^<�m�/c���f�wI�,����^�-��O�̓Z��wۃ&)��q����:'���T���gh���Z�G��� c|��d�]gI�Q�U\����7���0JBH;73D#l��8�]B����9-��;*f}"2�A3��Y7tQ{*	�wI�TGx)0S��2�v�آL�J���&�Z�f�0�U���g���p��nBT��Z����-�޾O;xM&��y��鹰wN�Ń��Z���v�k��[��T��n�:�Q���g>��00�x����v�V@�5wgm����&S�ttz�a���
*�f��q�Pll0�P�c�&fXK5���F�,h�j��~[��":�F��v����F�Ș�g�Yy<�}}��E��:|w8�G�X%���^;D��e��GI��v)�^��/xf���41e��l�LÅ��m�B�b\	���N�ɻ�S�e8M1 ��4��E�N��8i�9o�p���+�Oބ�A�=���8�iM�]Lp�ݤ3sf�b�}[��
a�:ٮ?�76��'\��SЕ���Le�v��'{h��ӹHܾ=/iG.gf��2�t��i4SL������F�̕�r�򼉳|��R�8f3o���͕�-�7_,�@�k&_v��E�(��|��Aܻ�!Ӻ�9H:齒�q��qs�.�ނ�ݸ/���>z��pQ����\��>�����Ώw)[�w@�q�sD���#`���c��������P�]�J�������TA_�zo;�����ι���DP����g1:{�K������C͵ 3�n�a'�i¨�zrƴ�-�-<u:o�"]ݝ�ć.�;6�H)2�wgd'�&�nfx�J{ेO�)��֓a�<о�׵�<L��,�\>~c4�l�NM��@���k5��)��гيۘ�������	I��cU�h�^���m��d�w���:'�W��,�6�P��{
l��I-U1����763k/;�f �T�ê�Q����o-�ނ�HP��X�/�o7^�.ӳYR�uN�k��5�;�:bǃ2̓~r��V��B��YQ���O$4Д߂�W�*�՘�^��	vГ8�Ԩ���r�շ��	gnv�c�4�ɧn5C���m,�j-���Zo��N\�ls��&�/OI��������Z��e;��8W��qᙚU�f	�{����H���s�lU���v���N��챭J�|�qB���X�R���a�㎸>z@���h[�Pg*L̖��b��7��dJnI�AuA�!���u���T~ŷ���A�gq�=�muհ��u0�b���]Zm����S���� ]w� ��[5f
�a������Qє5�F�q���v�B��m�jo}n �mo6��Pn�ȡ燶�k��em�'�v�-�!n���א��W���3���Q�3K�M+�p���H���m���`CosNQ�-���`�s�柳gȂ�ȴN��A���=7.T��V�
o�#\on���t�ͳ�\�\��g����rКWM�\ւ=�D�����J��emF����w�e65��ː){Y�Tz�B����aC�k���"�q�B�V'%�4�^gf�t3�=O3	�&�nӁ�_yx���� �}<����0=���u��.f�[���5&텶f*EX-5�_�'���5-瓗t�$�dv]�U�w�t�g�1���r��H���܌Cgɣ�٘�����K�����h'��n)�
Z����)Y�F_Q������&i���,�غJ�+U6�f���x�)ص�W���u�qa�Ǩ���1�s<SdA�Y�|g)ƫFvf�&e��ҳ|dY�^_I��7���ɽ}ޖt���Y9}p�/����䁆��� �T:�1��ċ����p�R��gl�T��r��O��o�O8�0����Wӥ�;��N�@2�.�T}���P87D��~͘�p\�	D���ѭ=�������Ū�p$�x�V�{�uK��zd�e^�+Q8��`r|_^�pc�U�gh��)�V����O1��2]�}�pW�ŞCj��7���ӧ*}��+
k�ŋ�Z�xe��3S�w��q7]@��r}RL��av�N9�]׮��T��+퓬����h
fY���$�v�	A���&��;+N��ʯ�R�?f>��Ir[Q9�x3^��e��X�y��*����Y+N�@1�$�`�W-e<tr�^VBM�Gh���
G@Lq+^�����o����
䖗2�ޛRN��n�%�����2��̭t�{mZ�����A�9��׹YV��Ļ��������cyޫ��FA� A�y_K�`���Ю�j�c��i��Y5�W�5*���v�����S�k��w,�G�S-F;7���`� ��TNf�_����8��5V4�-�
���<M��sH�[Y�Qɔ�8�L{}��G�۝�$
ƯobX�x��i.�V�8)�Z;�nQ;3��-���Ձ���'��Ie1xotľA���0kv])լ�ۨt������wE��q���I`4�6:��u|���-��A��[W�)qol�=���9�����[ۼ�5@��\���q����ݳ7���E�jv����k�96r�g�O��@���KE��u�9�}�����̥[��Y9eM�:>�np��{L��Y�3�M�F)w5��iGr���R����j�>�gd���::gR��ǅ�G=%[*�5׸d�J�V��)�S=b��� ٚ�oMUp�Wy�ۓ/y������\m��"'r�J�e�<q	or�@\�i��م�l1,�YG�r��B��ˎ#�wPsA�G�\[`ڨw~�U��*�DwL}���ޫ�ȩݷ<7��#T8�EzY�.���N��Œ�P)̻Y�|$؆�08Ǽ%�n��iX�;14�����Q�>ng��26��od}�t�'��+G5����;[Vv]��´"�p�A�bFȍ�ZWe��P];����G��ac�^f��T�J&'y	g5U�t+n��� |�NC}�E���2��H�^�E��ۥ-�n7FQ�ͅ���i�ڒ�~?S� Pc��Q�g���/��ȱC�R$+y���F��M.�p��2ɑ��]��I9mvobU�8�t�N��)�r��#y���WZ��"vN;��f��B�9 T�xtw�mV��2��A�&W H�|�o+B����s9��i���Щ�.�=���a37+1�w�P��<cR������]��w��n+5uіo�
4�c�\�@�K�!���v���^��������.���!�#�=5�޼�t��X<X_�5%�rO�/�6K��78���-�ȃ���B�`�N�L�31ǲSH��LեU�j��j����:��އ�-�c��L�{�Tsk������f�ۻ��D�k/1I�A�=��{�]|A�ɮ�\3�is`����nԪI<�Db7v� IKO���jF��9���o��-���^	���ѳ�/�k;���naX�4�F���X:��e�r���b�*�(s<EG�RbE�j�"l�r]Y�;����u����9���Qݮ��(����[��-�Z� �3�)Y���e=�8��v�4��ׁmZ5bg
�q����㜮��sQ���i���c������k����Jw�,�z��	O5�ې��c���y��:���H)�R���j��H( �5�[�{ð�۸��jC$�g!OvҶ�&5[��&�X��'q`�wʞ-�1��5��E�D�l����h�Ţ��Ҋ�@�l��G�&2��g#���κ�M�2Z%<�1���J㽧jR�Y`�s�R_5TZ�Z�I�K�yL3ټS ��-�A�ӂ��[���[�76]�miȐ]�>v�`.��[G���A�#���p�,���y�J�N��7H.����c(�u��r	p�6;*Ѩ���d�]f��m_V�	��R4.���j�:�[
���ڕ����rg'Gn���
�+Jup����~��1�EnK�g�6�;��r��S�:�끣�:UJk�����[{�i=�� Rk�ˀ�֓�"I�:o�M��EXݖ�����]���d��:�]�:�>t��އP�{�]jAO�-��X�'�>���������)����`N��T	�]}W)�V慶�5k8�"��rܝq:�.���Pe��+�|dI���Ni2��Y��f)�/��oV �+K1]�E��憁��d����^Đ��RD9��D����{�%�r$C^����i<N�;���X��v,�	��U�t�Ak���h�7��M �qV�-��v���b�~��
P�cp�.�U�n�x`.ӗf���\u{dTg����yω�&�ɣH��L�M/*Y�}Ȼ�V�!q�9'aG�!���	�γ��+X.V�������ӹ��Π;R�,�<-��Z�0&���� Q��׼即N�5|BR�3��6�Wo����Ǖ��<��x�J�H�4�`w5�h�hZ\Y���/�Ȼ�p�T]��ڙ;�Hi]e��*-=�`��ԥ��B��lu�;F�oiRr��uv�Pl��@JF
Uws�g�(K���۾�]pR�RӗF���61�Q�y��XVz�T^mճ�b�o]�����2�E��D�2�����t�J���[�%5˝q����I)y����5b�{Ґ]4s5���Ǝ9Z�9���4���|�ji�w(`)��4uYwʽ_m�lsC>�!�w����X@�lulF�����ǃ���m�v]�ur���k2�ʎ�R �m���9K���&"~��2bH;g)rذ���g�a���KjAݽ�ì�ӽ��uv�qKյ3�t��WP� ��]]aY��2A���h�3ܙM�3����o|� �_6�#rlb����G<[�9V��^c(��W(���B(7Zd�3�b���8'�M�9�>��zs��q����;V�o4��f3�k���*`�a%4U���~�ɑ�����vz�jM�B�c���Y�y�(^����dl�(�=�q�wg5͇l�
�N���b�@75gކӺ�ĉ3��'�K�
�E���P�h"u�6������T��̓�3���:62���S�h���ndQ��et5���0�=G��n��uB����y�Dׇ�<OK�Pf�=�F��xF��j��|��ی�zJ��P�M=�)�MnqQ$r�Ps���{\�K��o�OJ��P/΍U9�j��O�y_'�/-�%>z�b$2�T�,_hږ�.���t�悆@J��������[O��2��T���ԭ��
���ĳ3u���8�B�m5|�����Siowv�۵ͤ�6 kn���ͻ��X�Oz��ЄF�%]�PK�s�9�w���D7��X݃*v��χxL��`�"�C2�^	��lwB��2!���7NMW�,#|��*yJk9�G�B��a����4s9C��]��m�<��Ѿn�否^�9�S���DX��Žy�^_u+�W`z���������/�!��F�u�ǘz:Y�n����5�9�ؓ�JG��8������'Łfn(D�WM7�A�w�����3Qt�}@�]��jg��1K��&(-���w�]J㗀�N�rӭL��tNHS��	�����-�����cr��"�
�M��C-��V�݌�u�.^�ɿ��)�<��t�?G��䷨S��a��־���D�\��r�Da�l�E1
�9W�)����7���6 ��;r
V�n���h���/D���V:��!Z�2��(c�ݯ��K���7�u��ag3(� �r(}R3��/Һ�ۍ�y��!�:����=B�w^�i`�0���swZ��wt]N�ҟhd*yᑮ�0���E2(�c6�dC��P�z6gW]"�s��"�nv,E�8m�
��7����;n#�A2�^�{���@u<���(���w�{c��[��o:>H\~�*�)�P���9�$�Ѩu�l]�!7�M��7����zԷi��U�r�w��5F�	|�v�m�x٧���/./�����%+6���$F��TX���z��_=!���
�!^Pjem���ei��#��IhpK�̐��]�%���d�p���)�O���%=1�>�xe��A^�s ��7)�����E;��5S���-��G,K9�`/V�;o�)��K�'Mbn�+�[u��;.�v�x�a栙��	�wiǵ�V�[�e}�A�&��/�z��d\ų�AV6�0i�nd��5b�N��Gf�}h�lD�\�	kgf��b�\��[%��@�Lح��̑��c���s�0�|+��أwfպ�r��P��ު�C�`��sC��s��Y��Th�[��/zJ5��J>��H�s���ud:`�2�\n�#��
j�s����V�Ĳ�8�e����#��<���`�g{��|q��%R#u��Qnf^Q�hY�t�W�ن�RR��LT��(��JPf[�x&�P�Bv���^�۶�
F���fE&j��x�B�����z�����w0��:9*�~�K4uf�4xm�
2@�Yiu�.����ܴ��:v�=X����ߜֵ��XX�G��ry�P�(q FQ����;J�u����˖'�sqZo���D��Z�)a������sH��nھt"�y��>�8u��l ��AW˷7
��4�rP��t����յ,��+)��6l�Ӎ�l��{q�T����������s��vCS�d���Sw��+�l���n)�5n7w�{��.�|�TY��%N+,�J�n���\;t���DC�1*���[��z�e�=���Ei��P�b�[d�|�@�^��w�V���֯��K�Rtn�4�3n[��^S-٨��fKE4��N�M�B�!�܀�aŴ�wr������45`+�CSp��&���	��f�]�ɹ��+'v
<�5�ʇ*���5����Q�7ވ{�qu󒝔�=�(p��gY6��b9��(�&��J�h���f�,�̵����;7�0��,�g\=ˍ����6Ԕ�k�9�� ��tj���Ǽ��o����se�aՏP��������	Sޠ0��C9=,Q�m���*l7TV�����N��铚��bJv]<9�o<3�m�ޙ�,���6��g5PHf�}�=I�����C�l��;�{ZQ
���f�KOf��X��5Yt������{kӸΧ�2)[nΥ�^��ޜ���tx�]1�*}�R�[ݬФV7�T0���_X
��d�9Co9�1欣��X�ip��]F>mQ2����M�,d�7/Z{��do#z�gw:���s�y��k�|���SN�{���)vI8m8;����]�y�!��Cf�٣���B,�07���Ҫu��s"�;���ɫOu�"�氙������}����66A ��hO���{@VT��1<_6�=�����3_`��C��$���Vѩ��R��Ʃ̡�}d�%�xv�,`�2b"�7�����h����g�W\K��8g+��S�;އ	���$5d�w��8Ys~M�!c������Z8�M\��ԝ0�Ӟki���v�s�]Y^�J��,']4�ü�8'���v!9�{|��<��=nZ]��e�9�(�;U�
ˬw�;z�p3�
#U�=�ەvb�J�qЛ���kǯ��
>��;�"�P�c�ߕ-��]+Rf��!�t��3}��m�m��;�wo�|�&����ٛ���nP\-������,">��V���z��A¡�
�W<h�����}��[�Vr�*u]�����b��ܙ��ǨF�#c�<�����Z+�..�L��aB��6:�-Y�:Z�MSS�k�N�mg޸YNQ��.)Y������u���QW����R���<C}f�rx�D&��Yg��<�<"�{�c��7j���4<�v3]a���u��T�Ի�ҹ4*�V�tS7�h�՜��7V���սV_��料k2��n�D�t��y�V��;P�-�28��Iݡ�q��K$������*V�N�G�u��M����>�����0Gov̫D�"K���H����&��Y'��B-��/]�4	��z�k���� �Q�eEA�MT�D��T�MD�QMLUUD�P�MUI3UE���TIUDRQQ0MUMQ5U%SEMU�T�DI4ED��AU�N`d���eA1DQR3��3DT�VfQSUT�YEP�SA�T5K%QU5%QQDQ���E��ALQ�4�QDULKTDU41AAT�E�UT�U��UfL�EEQ%5�EE13aE�3UI5e�EQ@UTT�%���MSSEFNME%UM�DDUTQIRDEQE4�4�MTTDLEPQIIIQ2PED��R@QAM���]ޙ�߾��y�����۹���ĵ��/��g]�+l��ˊ]Ͱ9��3�v�P7��ֹs�9[���A��k�jjc��xk�kP?��)���CLGɇ�:U���T�]o��Wl��jw���rn����G�����O@:�}H�:��P�JI��Cp92��0X�⪡z��U�!�uk��*����ؽ�n���z�j�"Wh�W���_�]Jv!^f��	��a�.Ȅf�S}c��=��t��xz}�f|�g|��<������v7��}��*�C�b��3�'b��qv'���[�y~�9ĸ)<V��}�{��nz��:�>+���E�=� /�HT��w���Qoܬ���{���t�t�&? �9���×WxO���dz�;Қ�E�6)�s�]6'u�T����`K�����C�]��m5�ǭ��{}6�N����ݵ���h��:>r�0	#��43#����<#�-7�I�&����O`^�bd���"1��Z<��*���Ϛ����4Л.vڔϧ��;��<y�ȗ�o#��H�U֪hJ��(*��'+�@��X�W7�����.����5l�l�E/�&�kq�u�7�vIS��4��w�g +�o/Cz�w�n��5��f��!{e�"#��P�Һ�H*Z��7'w�L)��Ѻ}G��ۻ��,�l^�B��z�Z�#SEl|�<�40�=]�t��gS�/���3��{���k��T|P��u[u6������u*���R�M�0��\.�;��<6��D|�}�W��	8��g�1�9xo��Y�]R���q����`�զ�Ӟ��/�05=�s=�H�M�=����� Ȗho�J����E�k���)���/�/��7���\ۙa�6�om��=�k򎽕�T��D��U�1 �^�&u�
wgg��7�SŅw$�3�:����B4�w��r�����Ӝ'����WW����y]�|�7���+*���vX�y�dʼ�ɑc��ׂ+���jY��!��(u��w�x��9~]8l�v�]s'��
$�uL���|�}Hv�RVʧI���%��%$���Ƕ�R��� lN�s��G�P��We���6����jS<��u�ό��O
/�nF�G̞K.��2}V{��J4�'J��8�תu�].����E�����K����ĩ�Y� ��!hH�|�㭪��g�n%|�u���'�@����1j�U��U�m�c�z��r�.�]$����39"]�OB|�t��Uo/P������/��R��.].[�3z`W�r��d!c(�n:��(���8���K�t
y�y�78�@�ˠC�swM���u2�5v����X�as��<�uc�sa����-�C�;V:'��\�i5	!I���v���Bn]et�����~G�kO��)z���/�F��\�����z���qp���c��_�3�t�kn�f�^½냏V�v2���� ȱ�R`�;*�31�2�|\��x1��[:��/`Q�l��Fū��;�ex�^�N�7�i>�C�v"�6��3��c_sɐ�n�J��u@�)��)�w�� ��T(v�*x.��UU�h�DM���%�a��ƴ�r�|罼�����uԁ��L.'��#(k!2�+J�2�S4z�]]A-
���:w;�O��,��5c�a	��Rd������b]!�hmX'�`q����z	s3=c�v����ѭf����<���F��-���5���&]�:
����'?um/k�/5�@�� I�V�:!��3�[jmz_�:�Chps�g�>�=0߃nˬ���R����������0��d��7�O����A�N�L�=,k��Hg]bx�7��8=���fJ�8V��I^uf<�l{}X霂0�Z6���Ei�Gu�{Y\�K�D���&��ve5��|$fp���e=��{�D���v�-̘��ݕ����C�%y��/:��NA�|����R��g.��	 �f����wY��=^�B����ɂ�Ba�7�K�T��du���w}
T��(�����w���[e�}4�!��ӆ���xN70)^�%}�xo�P^	:W��U]%� Z��������d�T�讨9P��RL(��["8_�;<Iu���N3�mdi=�&�{v���u��1�I�Hk�M!L�D�)�w�O���f���蔗�:��G�:Ƈg��kO�;�u8�Ep��xh/���;�t"C�U^�>�]�Pllճ��;8�y`�6r���&	���^4��QOv��9c>��l7�0VR܋�c�o�����G˱�`�<�Bu��յ+Fb:a=�ڭ��C%�2�/��� ���v&���S���m���L�\~��t4�\_t�+����@�J=�p�a�{����z�5���I�����ju-�z�ϙ��s�!�8&l�����]�]>�p4JY=W����x�/��l���)	���<��>eI�dЯ����@��=�.^�n�m�3�k$62����c{����,����CI�}�FfvҪk�\����f�ΙNߐ~������ʺE[[��~z��$��)��/56�j���&�Ҳ3p�L\��b�㲴X��k���&�z>Y�lS����@ҭ�o�nݾ-��wԂ������򃗹�������/�f���;�6� ��z�|�t럎����������Ǜ;��9����o5{��kO���z�o*�M�l�rh�"��u�(s\:�����@te�6^�����F�k��ɒb�&rO���0�s�C�����W��]�]"��B'�w7I�x%�_>�;�d\�H�A�DP�x؞��Tw:!�61�|�-s�v5��+�`��wNϝ��J��E�.MB!-�x��/N�c�\d�Jw��FB-_��W۾[k-{]Ndy*�N�94P�d�ϗ�Ő�nk��w֧�	��C�^���/m��˽�iq�	<ǥ_yQ�B`�	��̘p�gL$��1���vhh�t�.N�2c�����q�� \��c!������տwvg��w�a��:>�7���o�m�V���^{�����K��G��������p��]|��W�{�o!X0n���K�5��{-'��#{&)�δ���,u�uj����du�\���A�vWh������J�nˠۨ+z���CV�R'��g2��k�K[}y�}���w�pyy�P�yٯy=z��"��@���[���Nɯ���������]�^��l���A����^�s^�Ok�	+���S�I�z6���_�W3a7ap�3���\A�Y�t{�d{��.�ݯ+B�r�e��~k��e-�Ŵ���H/�u��.t���5)g^�Tn�����-�lW7n�;���_W������+�HP�3ٕ��]�ܘ��n��s=�Wt�>�Y��m#�|X�v4*��r�W6X���x��}�}y�u����gkY'<́��Z���Z�����$l�d����V�sm�{֑Y���N�	�e�\�Ja�,��G���fߢ�zߋ	�;'�7�q�]�YKz���-�"՟L䃰�P]֝ظ���7;B�t�6����!x�t}&��v��r-���I3��XYN��#wv&߅R�-�zZ���UܔE� �.���X���H�Gt�E��Nf-	౸��TR�YK�\�<�Q��!<+��m[���j���v>�QN���+Vqs5:�XW�������n��l�b����ᾜZ����m<ّt�]:;�Q	z����.u��������_ku$Q�E������x�>���X8$sg�~�o���y��G�_�N��^qco �]߶���F�A��!�z�j�"����Mb��wav)[���u��-���z�wBm�c\ǧA����E=#d����y�j��n��v��x]�-��<�^��Ͻ���&=9�{�V�Sֶ���3�C?W�`��Ҳ�7�).�%�\�$q{�e�����o �Y���)G���޳��|�y!O��}�����^��w/f�]�5��*��kf�l�g(�G�S�@K�B����<^W���F;)�(�5�݃X�wn�����g��OT~��kX�lzV�\ͮd�.���S��Vm�����&`�x�'���tf<�N>�n�m�T��Z�2�:m�:���ԯ:�K'��Wd�ʇ)�"�`T��4�z}$��� ީX��dCZ�u��]��s��S����Er�f��M�C��B��F5��pʴ�Ƴ��r���eZB�Bv�8��2e�,��I�i�;�|)>�ƭe\lwG���ŕ޾[���׾�$˛R\ձ�]���z#��$Oa��i�>�N59�y��r[���}]��s��5����8Џ�W�~��CV=�>�(���Ȭ�<���;]m
�e<�w9|�<��#��G:�x�����837���$;��"��6+�*^��7�=�����O�3��x���o���^~��n��D�A�D��x�t�_[��/��f��N�:����k����v6�E���
��95L�+�g�Oe�]�m熹����{9�2g���4�a���6�p=wO�	v�i���s�7���pހ��Zخ�-��˰;�R�#� �zzK9��z»���y<�'z�]4{9}s<�;����<�ӎ��	��F�>���etο�Web�{6�ʡ[�8��-+}ʙ��q�l��"���!,=9�a:���`�(e���"�7�{PIf���(c�6�gw8��6Su9'��
�X8bI}���d�͘:��o�n�^l��ۼfaJ�mxy��i�v���f�y[�^��<)n-C�Z��yo�%\,BDˁV�㖶�\cs��s\�MU���{��ͮ��V�(E�9^V��y�gzxHY��^f�t֩�����/g*qdq������h��l�Yxg��|�Kvmȟ����c<&=�r���0�~�N��H��g#�Mzg����ȣ��O/�񵢯G2�����鎤�	�<�s�^�h~��4��~g�������g9}]|��خ����$�L��f�ҩORR�Nփ�c�j�In}w������[�'��Qusu�c�7�����w��\������L���vE���u�(s���t~�e�+�/��RM���ڞ�wO�sˊD�L�a����!C�:�{�{=~��18�m����F������ޙ+�� �+Y���5���ܥ��(�G��kpI�\�XɝәS�+�ܞ�dȄ��v��9u���ʒ�4�b��ٳ��<\-jJ���;�'�-���@`r�/���uJ����4������]9Z����+�x��'��]GPbL�l�Y!f
�`��netSu!�����=�fF�����=w:̂�w�L��cw�ow�c�5������5�8����ڳ�JA���g�;>���uQp맸�F�e��cz@c��G��g��5��Q����21�j���2�\��̘�����"��Ly{<�{��[��ф����7��ȧ�vz!S<�:����3������f��Z'�vOpg��^�彩/1d:B�V��X��^�B�#)sCV_��\0yl��n/`󌬎v��hy��z	RX��W��y涯|���V�![�i�����Â��Rׄ��&�����8�O��q�%O|6�'^;T�S�c�,��A늜鷁r���ē7�M�4sT����辤v��|+��V����8W���\�m�Ukgv^7��{����9�"|�#��luZ��O��D�Q��r�+%Us��VUB`��>�˻�E�ط��8�j�ӗ�2�-��Dz���D^�a8�;�B6Ej�6e�W(7��ǯZK6�Pn&n�]޵WdA��V��G�Ȁ-cz<p��u�д�qj�:3�ab��GX൑�7E�sD3��bb䏴D4�%h�� Ԅ�T�SN�S�޵�8�tյ6�DH�1ՌS�-;��6��(|���ͱAK��x����4�%G.w��L��2ՙ��+3�[�0r��Z܈3�j|F�&k��ӛ<y]M���*���g�6��1��Ǆ���w�0�ź�U�P]s�)�R�M/1Ε<Ƌ�w�t<�ͭ�~[g{S�#��8L���3qp��
c�����N��(9�2�q%%�.��ڏǅÓ�S�?T������L1C)��\3(��έ�K+8xuQ.:�֌�8�a�Jʱ���oOk��fN� ��٢�'k䏟#�����Wh��ڜ�n�Ի��c���<�|x��z�!�me�\��ZY�w�pY�ϻ�����5;Dx���7qsq7��Y--u����hY�3$�>&p�>���0����T��pk��vH�n��J�!������a�w0��,��Z�ZŲn��(��)������5[��R*�FW��%�3��u�:��*1ı�������:�HK�^v�oyPҌX��O�v��c`n���Y1M�4t����r��*�N�����ȶ�sm��r5Z6k�������j���w�>D�ۙ�g��v=}�J�k�	�#�*�dդ�����9d�};���]���Y�m<7����Yj�RrrQeX��9
so.���.��Ճ=���$�s��.��}yf���P^l����q2�wnSh����JZ����#ڟ��n�9��-�R���i�B�������kw�2�1�m����x����05�3y���<���6���acI�A�;-��ޯ��ч�Eghװ�����u�(��uoyu8�U���h(�2���*�D1Ǉ����Q���ʾ��(�!$�L��F���|4��6;�5��d�-ɦκ��[o���K��1h�[��x�f�=3R�9V5{;o��;���-����t�d*e�8o�z�׳TyiQbaw|�:w�WpJ
+�s]��=�*c�����A�����p�a���_���aD���˛&�m�X4oi#[7�����2��m-��z��w$b�N�H#�A���[��δt�����Nd�Ft1���U=O��ڼ�Dn�Vظv����/�7�V�Z�n�w�k��y��	��� ���;�Ң�1Ov�еkA2��,f��m��.uc�E��Ж�J9Ҵ3�8�Wo�v��kh������X���9W�x2h��ж�軎�h�*�b]�������\�����1�^V$�Z������	 �GĐ~�BD��QDAKMR�DQ%PUTR�1D!	AIDE%UQM	ILUM EE44DQTTP�4�ATEAAҔPSLIP�R��T��4-P�����AU@�QHD�EL����D֧&�
j%)���(�� )32*\�2���*�"���
h)��*$�3�h(����	

R�B��a�d����Ȉ��L�
�(�*����(�&���b()"ZF3�r(�����j�i�h()�������J"�"H��R@h�@ Q 
 s��^^J�������ӓ��烸9c,�Ư�J�Hg�q�E.�Ղ�%�[��.P�;��O����H�����:S��S;�{|'3��s��K;�gl�b��a�0_�����P3�����o�:?2�Ν֞�^|�<N;�X�E���n	z{�ux��q�4Z�_��Rf˖����χ\�q��2-Qu��}��߫;v�R�����e����|7!k=/��b/_w룬%��>�	��|s�����h7d�5�7Nu�oo�ڎ��{�ٞ�k�wJeɃ�<�y��*kb���.'��<���V����f�ڐ�s��]����9��T���s�M7%l��B��k�ÏD^��Y���Z/rC��-mʹ�׎ϖ��{f��	��V#�'1�΃o��"��:�����bY��ݝ�V�{N�>%C�o�5�we	1�ϣ�oFg�t6���JC�zl�3�l�z�?i�����Z�������8Ώ�3�#��u��{t�'�F8�cT5]�vv/-����L�V�vC��ݲ����<���{�������&��p�9x��UqG�%��F��4�wM�t;�9��V��*:�A�;h�m��\:�!xyU}�eb<Y�Y�ЛC���ߪuw�e��o����z�߻���Ɵ�ki+�*؋���;��_gl����<��c������M���p���i����mV��y�G\7��c��=������7��~/���N)�Q�G=����F_i��ghٲ7�i���5l�K`)eg��B���:s����q��oE#�|d3�Z�:�uw�]t�A�1��B�ٜ}�#�|���o~�{1霢;Wu`�w.Vk�N���V�uaZ������Or?_�^�ڜ����&�~��j����K�4]�Z���v�������2Wg���ک�`��:���a垅�X�x�EoO>���qk턠�J��T���{g���� �^�e�\��"Q앬��օ�ٝQ��{�<l^��T|yzs�KQ����Aɨ	�;%}��IT�K�k�cz�h D�X[y��tNY@P���&xN�>i���	p�}�Ou�4x5!OtB���2����v{�1�-
�p��U�6U�'|kX۴��QJB�Cȏ�#'��w�Ra�}:�.y�蹷�9�؞$���º)����� ��y��<���y_�t���.�Ҍ��B�������3¢�d�Nd�>}�S�Pk����Ww��ol�ҩc�؎0�p=8o՜���8����2���s�<��=�}s<���3����i�\�eh �������̭�m��x�y�r1�����8���_Sȱ;�,�W[��ۼ�r/?{�g��ݰ6ǐ�FP1��9��f�����%O�F$����tɫݽ*>��/h�r��}{�|\��qׅ�;s�y�n�e'Y�/)nϧ�Mv�|֗�h����~J�g�@���^����|z?`�G�=7)O}(�;]�ض<�kΤ���e!����e?8�ΘI�N{^�s�h#��M�֚���6P�ݕ�Ъخ�͕��bOM3�M�
ĦՕ�w�b���������S{����!�Gp��`��W5r�}\�C���0f�B��<H��J���o�y�k-m� g�*Ʀ�ܻ�>���z�96�}�V��(0G]k�)W���I�co@Ue�m����RR�7��� ��]����tv 0��u��/���^#ۯk����I�2�1��զ;��S�����[�G=�.w����زf�g�@�Y�;"��w��
��3���2�@y��uH��O|�7���5�Nyx&I��K��vF���ww�	�̗��y��N7��v�iɸ\�uk�����d\��"Qa�Eꠞ�H�̓Ϟ�w�]@e��OV���ŭǟKQ�2�\�����h�����&�;^�F�'��}Ț�6*l���[����O���%�`B�Z��fD����f_N4/D�ڃˉ�2��w�d;��|�^~�仔��惻�{�rx{���y/p{�rWQ�~�g��
3�^*w���ۉ���>G����>����:7�%��2N��hJ%���w'G��r�W}�iy�!�nW��v��Ի���z�C�;��^�����^��v�� ȇﴁ�������0{������G%��[惸w��v}�	C쿟:�򼗯���ܮ���w��:�'!{�����ϵ��^]����]k�~���R~��ך9=K�9�{�<���ٿ�/�r������ty��q�<���>NA�bK�=�^������Z��wtzg7�]s��z�����=�ݣ��FI܏����}���z=�����u��K�+^���=7�<��|���K������y��u�!�ˣ���g|��d�߿<G]��>΍�$u�HB����G:<�ió�)��|�s�T*�9	�u���@6V{6>��9�y�u�7^����<7���Ǜ����⃃��C�+�Ր����D�}Xs81���gS����?)�G��p�:f2�v`�6��� ��}��}�Ĝ\��׹���:���y������X����GZ�r�FO������ڠ�.�뿴���y:��<�zǑ�_��:�?|Ο�׾>��W�yZ�[༻>��}/�~������p�Z\����?Y�w=�|���:5��~�#���t~��r^AK��4;�g�!ΰ>�}��7ݷA�/߄�s��點�뇝���a컻��t}#�콧���B��]irOe(<���nb�G�wkJ�#Pn
G��?}��?}?[�n~]�=�H���>�;����2_$�xn�rp���[�r����_�u�܏�ֺ��>�~�'%����=���:���!y��ߒUY�{�����~�F���u��FHp��7/=��ئK�9��C��C��4����^��w?K�δ�+�~7�K��	��~�%�~�]q�5~�����61�=� ���q����?=b}�ytk�%����w/;���i�u�{}/r���}�[��z�7���^u��<����t}���~��׮���H~u� Q������;����y��1]��_h>������z��߿i������r�'��C��_d����k���4u�z���>�;��������R����Z��׹�r]�K�X����F#�}�Ͻ�9d.秽�7&��䝟sG%}�g?i�^�~��z���<��o�������Ͼ��7/P��|��=K�ӭ�<��}�Z
Wpo�.FH��%�2_u��K��:���_c��Ol����ޔ��z���s��������꨽�a�}g�?�~���W�|��x���)���9����~��=�K���=�ɒ�w����?}�P�_|!�{����L������
��v��.Y��Ӄ����k�e�G'�S��L�i����ut��y|�Ix�@�
�]�>��Bꧩ�ޗ�%;gZ�h���'{�����n;,N5�i{.پ#���\��o�?���*�:�K*�~g�o�""{��{�z�~��������_%���iL�Rty�+��?ގI�G\枡�'[撃r�?s��7֟л������+�����p���t�e���]���O������~C�~_?}
��������|=�H{=K�;��%r2O��tr
WW7�!�'���ܾ�I��Д>���u#�}ל�o}�W,���~Z4E�l���}����uw/��X����:N�:�r���G��{�rx���z�s]��B�$�����G��仌���4ɹ}�V��캕��5��9�����w��7/>����/^w�˸}����#��=NA�g���'RnG�_h�:������R�^�^�䞜ގ����3� o�~�)ۺ+=߿u��ﾌ���;�r�{7�y/��w��|��,�R�=b>܇��5��|���X��r?������]��� ~?}��k��8?{2fN��~��?.�>C����'�^����9.��|����y:�;����\��w�����pt��K��5��|���X� >�&�f�?q]�*o�s���~$!�
�q2%�2y�t���9?�y'�kG%��g9��rOo�������]ir^H}���Ϛ�<�G��w��J�_���i�ɾ���}�O��B����7/ђ���仌����2�}�y�+�>޴r]�C���{���}iw#���Z\??|3��{�6?{�WL�y��G�)�k���:�������ҿ]:�I�w!�y�'%����y�;��q��sz��{�~د.]}��d�u�>�/c�`�������}�\��J7&C�)8f	�K�����x��>�п]k�'%ߘ�noAܻ���xs�)�:wּ���z#����ݎ�^��n�����z�>ѧ�x7�<u˲:F˕��j�u�<���#�,��
r���m��s��w m17�ڭ�ͧ�	�캇/�"YMa�Uႍ:���[��N���?���7�w"�ܴ"���έV���:6x� rwϋ�$��۠���552-�5�UW����}~�{ߖ��j�_d�?��iOR����+�~M����q��pP����a+�;��{:���_h>��������ry}&��������������x~��~��p�]���{{/R��}b�7/P�o�G��/7ޚWp~�Z\���{��d��� >�r�1@�C�U��C�~�������_�)��������p;�w�����^�ް�/r>�y���=���4��������K�:�P��񾴹���9/ђ����������u�s:��{����:������|���u���w'`�{/�=��?J������y�?K���vo�
O��=����s� ��߈�L����>��v��\�o��~>{��}�Ͽw�sP�}�sX>��_��؎�5�z�%伃�oBe�z���y�]NA�{��9+��f���
��IA�}����	��-��������g��v_��^}־�^�^��+�;�'$|�Z]��~`��;�����r����wy/r�=�H{��;��r' �y�<�W#���仂���]���w�ןo��߿f��y�ĠԿFA���JO%�o��w���s�W}'�Z_.��t~�ܯw���R�S��z<�Kܛ��{�GR�N���H�A�������~������ǻ|����@$}����l���������d�s��^�gr�������#����G��ܯw#��:�r?��G�Լ�p��w�n�������~�~w�qu&��
�~�B��tsz9#��y�<�s���Op�_}��0%�_��ײ����,��y#U�}JG����Qp�Y�99�a�<��>��u�޸���y���_�����C�+����y'ZގGR��a���;����7/%��7ހ��=��z\���`�d���f��{���G�'s'�I��[}��y�ޘ��,Xc�뫕���u���Ԫc	���x]Dic%�k����h�[-P
�B���&�Y���D�֎3�[��塤,W�0�چ��H���.���f�➻0���dy:�N������.�&�v@>����G$o���Ͼ�K�?��7����'�J���ܼ���� ܼ����H�NI�a��#�/��w����y.�a���y?}�A��3f����:������������>����A��F��|�<����X������A�y	�ؔ;�q�������r�W�w�h���><��߰ך�_{��sμ�y���^_K�ؾJ�g���O��O#%�NA�k�O��r�_`�x�9#����&���O��P�^y��=ҙ/$֎�xx������ˎ{�oﾗ�~�U��/���Y��z�ZL��w�\��N���2]�I���9�f�~�q����W�>��;�����ǿ�:��?&��ӽs�g~��a��x��K��P��;׷��^���z��{����#��^�u��_gz�ɤz���w'�0O`ܼ�%~�s�k�O9���w~�μ�r���:��x�I����w/%����%�Ga�4}n��/:���^��>9ޑ�:��}�rGpoX��{��d���_���<���|:��s��~�^zp����}����O����J���I�������w�w��:�����\��~���z^GR�'Q�\Ҝ��zyւ��~�������7�Vwy�������<��>�C��9�X�ܻ��G�Gr�?��A�%ww����y^�N�ynN�~�Ԝ���u/�y����u/�S���߽o�_s^��W��7������\Pn�AH���r2�sp�?NK��_e���������{����Ow�e�A�=ӹG$�0�B��yٟk[�����f�w��̭y�z��>����M	���JK����A��J�O7ޗ#$y~>ť��C��w/��~����w)���w��.��ߴ��{�5�G7�u����c�۾��]V���T��8��v[�ά5u�9��T��]��
>������wV$��QJWN�P���nt|����+�R����fgh髴��ɫ܂��!���X�.��w��(�j�q�O�L������������9�q%���t/�W��#���oGR�
C��4����:>愡�_����Wrt�ޗ.�w������^���N�ܦ��4A���*6��^�O{��m?�C�>�>d}�؇��_������d�AJ�zw��pRo���>�A�0J%�μ��%���.]�ﯴ�w��;ﻙ��}�w�3��ןu��]ߧ��u&�wޏ'�~���u��:��W{�B� ������ty��q�=s�=ø}����<��}=�^���uל��u�石�=��k�o/��ڗ�|����_ђnG��y�P���z=�����u��K�+���_ ��<�ҽ��Ò��3���9�w���O��n�!�y�[Z�O����?}���Y��?�`�d?��:u�{?K�u�w+�d������ڠ�.����/�n^FO��;��u��yJ�=�~���o�}޹�~��}��y����G����y.����^J�g�\��_`�d?���k�?K��X�G�2?u��)]�4��R�����u����g��w�u�����>C�����'7����=��G�>^�����B���Z\��Oف�伓pu�S��.�XjW�9@B?��]韖g���ok�?zv�>w��w!Ͼ���ӑ�<ҙ/$�����/$�3zy'��ܾs�J�}/?b�G���Z\��J'%������ ~?}�$�D����w������+��؞��_.���r�2C���;����}�2^I������?<���=��Gs�<�I������#�#�@��qH_�d��{ν����d��I�1��_��F+�?GR}��ϰ9.��/�:��y�}�=��u�{}/r�����9n���|��҅��j�M�����W���7��BM��+F͝������u��_���E-�u������'(QU�R�������..vݼ�9[��<�aJ�z�v�,WQ��cf�7�d�XDaJN�=0h�^��y(�'.�3�/o��	�N\�{����>�E�c�<���&H�'���C�P:����
J�wӄ/��>���w=}������޴��{gߴ�_dz>޹n_�?X��%��n]��?��g����W�:���~��)]���Z���{��%�d��`C�~��b;����zNY���zMɫ�y'�Ò�av�V�L�V��ߛ�@�����?��h�^���oC��_����4 �^�u��w�}ir2G^�2_�%�kp���t~�w/����'����Ё����_��@�~o7�_���}��'�ѹO�u�h�NJ��h�.����4���
z7�)�=��a�^C����2_��;�.ﾗ�ߴR�|M��D���ށ{�]Wߨ�z���}���iL�Rty�+��?���rGQ��i��Bt�J���}�	C�?����.����.w_}�.�W���C���nw?ڦow~��~��_dz���1=����������|~��R���\���?�G �u~9�<�pP���ܾ�I��G�G�4�*ݥw1cGۿ�ϵy9��}��;���.�qi;�����'%{����:�r�����r^�ܞ��<����{�B�$�=ގAJ�~�����Њ?|+'����i�Z���_��p:��~������{/^���~�αr�e�z�{����X��y�u&�u��c�y!���/�u?~ |!�� ~?
��?Px��}�z�w����;�{��Gҽ���G��2S��h;���{�7�=��z��#�G�>Y/�w#��O��ܯ��Ԝ?~h���� �ެo��^���}������|���Y�d�j�}���]�нA������<�K�w{�;�H�uδ�/p����I�:�)������_##��u�{��]g��(�_�W��9�*��y\��"���G�jł��4�F�r*4r�S�5W���
�ɿ&J6D��ʏ
�c|>�D���[�����c��qG�+kL��"��Qɡ�66�^�֛o���e�E��C��L�4��Os�Ӹ��%^�j(U!������yr��iV,bn�@^�P]^�JDw�_>Q������>���#�<�:.[�Obc��k���š��eP�����ޔ��q��[���ʪ}]Lqtm5f��2��]LjWR�c�w�mV� �Z���!�q�	YtW7��P���D���� ��l�aՆB�M���a�2�4�l�c�{j�����!�h`P��U�Q	k��ي�jsݛ]l�Us�o4�'ǖ��k�s�?K��x�h�p�G����I\�F^f���'qMw6R����Ԇn����.kwh����䁬}W9o,X��!��r�(=Y;B���Ґٯ�wY�\�ӭ�`_ڴ<z�w��m:!�2�3�a�+���Z[3zЀaC�+8I/�r�v�d�a+/�'����SU^:�+hgٺ�k�jزE�L{�T��Ġ�����i��<�΂1JR�|�u�6�ڱc,&��Ե7�G���{	�E��x����'��G�+��B������
䄷,9�Z��6k;-��+~C�6�I�qC�wWv$F�w�8���ʍ學V�-�}�+HݕΚ[�	��{��6d��>��P}�v�D+��oI��]��3E�MZ��RA��uʰ.�84G]�F��eg\Z�z��	`��M��~��0b��k(��<�Z`�@���Z��77)_dfj�,����raAd�:�{��U�uƴe������|�
h���oZ� ���̃J�W�u+q�m�#�W!W�{D����I��(O;��dnZ9�M��?�D�����13��e�,c�3{+��V_wu�Jg}������g&Hfz��O%߄1�Z3���Z:-�vn�ԑ�#�>%�;q���a�giJ�uL�w�][�L��2Ì6����Uɢ�İ^|\#�2kevq�Et:�{zl�5m�;���r���jî�C;D�7+�!��G��r��:ν�|�f6#w��}����H�+���s|���`����$��aWm�����Wָ]Z:�|��]
����`�y]I���wuE�2GA�c�z���w�W"�M5��o�ϯ��,��Ds}f�G|&'�ܳp�T����x�y&tp�v[�F��b��m��8���'W!�ә0�:����Jf�fu�"Toj~ӹ��Վ[�n�]op�rtPحM)�+j��,����:�R�� #w`�wa�`q.��
i����^���ܕf�[�Cn�F�s�Q�]?����~�����>�L�!h����(����"��$��%��#%)b��((�s1(�)�
B��R�f���\�����p�j���)
B "ZJ�J")ZB����J���j��(�2W$(JJ�rP�Ȥ�����!�Z�i)j%)�L#$�r��*R"��B���"�J@��3C,��" *��r\��1L�*C �B���s1i
2"C2̅�2F����B�2W$r"���2��# h�!�)C!rs1� )�JJ()2T����sr�#$b�Hr�$� ��2J
((^�ִ.�n��ws�<�gu��<�z��u\�J���4w[��Զ���d
����p��D��*�njk�vu��T@s^}��[�[���I�
��֨<��(����/#'�~���:M����G�}�r]����k����u��^�]u��y!��K�w1ߪ_�9�kw2��Ӷ�~����?}�Q���u����P���7.�$:;�CI�w=;�Bd ����W�|�Z9.�!�_}i_/a��]��m�g|1����R���q�>���k�P@��\>�B{��9�5�����ҿ]�I�w!��i9/.���S%��w���?�������/��׿��������_o�־���[���C���ǿ��'�����2�I�0O`伎���~�q�����־�r]��[��]�˸>9����k����^���b^��=���?���t����-�ˠ��e���
��3�I��}(�ڽ��;�z>}-�V8�/�痓$œ9'��h��x�y��5ߤ�ןG��
�&�����n{����>����Qn"�D��݇�.-����z�d�ͽ�gvO33���=��}-G�U���/�������N��fL}���<�&}��*��=W�te�=��r>��C=j�y�j�k�	��ほ�����՚.;��{މ��M�8pI��!/}�{�[9N�L�ԱR�W˴���J/��C��:�LE�Y$�m��T��@ݼ�1�Fy�zH�)�#�J�g]�!mY�1T�R��b�+'���\5�u��yc]Wj����Q��fr���{��p�_W�U}U_��&�g���kJ�1�u9�G�+y�w���ɕ� ��Q�钷r�����5���63�)�zs��m�z!�q��n�8��9���/z�p�EO{9c�S��{裃��2�ɏu�n�F=�|{<�|�W���r�\������{����3W��}{�S�28���o�{u�9.̚E'���t��sW��<r�9a����Y����w���>�G�^��[��T���w��Y��R9}��^�g|��z+86_�.k���0�����~�׭܀>9�E�#��g��UlB��͝bOr��@��2`�ғuu��v�s�����#����}O�<����M��l��,y����e�>���c7��yH;]�u�<!�;����tօ����c��77m�&hu�����毾�&,9/���
�{MH���29�*8QOtAM�*�]����f�7�N`��{%�/^�u�Rq�e�}fm{�k���'eoy�Tn��L��{y���b�t_�d@��b��Kv�ﳸƤU}-�'�[��x�
]-Sb'�;��M����S@��V������;���֧�Q���r;�q���v�>�;�d\�H�>p�,����iͳ|��r"��n���{{�Z�bnr��}��l��-ˢ8%�7)��z��k�WeM���τ}�Y�)��2}EA�~ *���m�͙���'͇�ɛ-O;��&��f�g�",��V����/�8��mv�@�󎐑0�J�<�"��]Me襅��a�5L�Z��Xv �7;�f��4��g���1���m�/E�a��F��,wc��s��z��c��}��'�[��ޚ���=�N	7Q�dg���|��}�q��08A[�<�s��/F2�����ΟJ �{�z�Қtz��}��^@{�⭉S�%��&/��-s~6U���V�W�߳�2;�r���6G�RyR*���z�||���� T��/8�-BV�gAe�����wÚ������r�q��v���r�#�_�X�B^�}�6B�9�o¸f�� ��5���R<�6k�d�a�l�ݬ�j�)�����Β�<�淕�ȧa�����)9V�LpN�W�슒�γѪ��\���U��|{&t�sݽ�6{Ӌ�8:��{=K[>�Q���N�=�'n��u���и;7�a��9�8�����Ue1y��jk�j��;KSM����Ug!{m
��y&�1�3���Ny���Gi�q7V*(/�U��F�����k�:w˯�G��2N�	�e�y&a��~�����IyϞcl��k,X<��k|�z9���7{��g�ծ$[ـ<�2��߼����9jk�C��4F�P�.�������<�#���FA���D��Vl�Y�%E��p˓e���x�:����{�w�7Z�r��^��s&��lfw�\v!O\�6x�ꎺ�(y��a���^
��wl��Ǿ�p_P������E�+D�����3���:2�i�K՗�ٵ�ЖR�x{.���1y?w�1�	���W��0�ǧ�S��>�ள���L���!�c�İKdNk_��Skof�Ɣ�X��*�b�\����+@|��`�����=[ϙ�,�ɍ�ù:Dز��-��E�\*��9�R��%��|d繄�꩸+�N���w{7�zn	��=]+�+�<���}��}��R�aŷ8����QS�h�5S<�'c3����zu_֢�\�w;zʤ���[�����V��{k��$=�bv�T�o(S��+3��E����^3\���Ҟ�1O{D{�����lE��G�d���W�*�v���ǽ��'�Әυ��Y�8�$���pOU��O���.���⩷��}��v+0{¾�;���d+�'qN1�I&���Hŷ�R�N]�;���]<�^q����UN@\z+86P~1���nN���.��G��o5�(�ou�G,/������._!\��g���>y�/���:}o@:���q���+=����;;`�b���\���ǣ��̼_��^'/ɪ�}�kn��L��$iDvݑCx�q}C������s�S��q�;�֟A��; jw���_�$œ9'��h���}{C���v\�E\P+|�ܭ��r��{��Mho����r^RY2�M�
�"�q���[��D]�<��fk]��T'̟3�R~����笺�&�j� b6)v�JT�x+h�S��q��݋nS���GtNV�7
ͼx-2�p�#ax<�?}����b�{��_����o��}�Τ��-g`��/W	�!07d�fwxm�N�ͬᰧ�<���n�^{9�5Y�R�s�%��J��p^��0��q��R�^�/,�Fc��m����B�n/I��K�l�܏��b�ޣ����7Yy璈�����/�	v4L/W�.v|IG�8�O�z��4���l�Z��Wwv�O�wzJ�� ;44{=�gs�O����J�E��3�}���ϸ��x�)�zzo�����]�H��cmM�yǖy�&��EM�������C�3�?{\�C�b�ٕ�m�.��!f�����v�-�ɻ�LZ��oJq{#��9��;����$+<=>�s���K
���=b�/Da�p���Ptyh��Y]Ե���Bz�gݞ�6VwhW�!S����g�~sjv4MaR?j�v���Pw�t���j2#O��5�;�Vv�6�]M���{6�f+y�M�Q[��(��������sav��s)v<��ҭ�_fݬl�0���񹷼Z�CCW`�L7�Z���;��9MeE4:.FЖ���Us����@��_W�UUV�s�����ZZ�A<�ӞC�4#��hW[B�b��͚�DQ�3�L�r׼�o�ɍ~��z�M�>/{�=3�Go���|_�����U@�6��@�,�{:�Kss�8˙��L�̐>�w���_̾۲�}4i
Q%�qG����6d�;�^�<�42sˊD�霚.qH;�M+�]_�Xu�l���uϗ�:Z��wM�\�e{I}�\�{qILl�{!�xϯ֩�Dl<s��־�}�3��5��Z��(���<wӋj�trџ[�,O����7Oe�{{�����^=�AW@�ޑ�@���R�X�n��96x��:�/qyG���8welv�ӻ�D���.�w{���(H�_8��<��aǢ$�V��:������v's���Ǔ�{T��8�pa|�=8:�/L7�����*�Z]�R�`k"��X�^�<��r{�jy�W-Ѧ�`����6�c��y�T�%<�,��,љzߐ�pn]�w�Ωs׻u��+���7R����b���;���r\U݈�w{�zg���s[�#hαs"�ݕ��쇠S}��|>.�p���qb�Y������1����3G�q���jK��;5��x7Ϝi{�3�5��Pp�+o���gн�yl����~ۿZJ+�u�ȕ0WOG�_���mV�{Ņ�^v�~����{�c�_k������Ctܝ�1��'탯�'G�&���O!H��wg�_R�:]��8��܏��=�t{L\_
s� �Og�{ۗ��Ԏ���u�֝e��L�Qk'�zLk������\$(O���8��O�#��9�����Z��%s�+����&?�ʹ���ɹ:��_�Nw{�P�'��,xT]
z�<����J�V���q����;s'gy�Zq�of�V����Ű���W�N�3�Y7�y�=���d�<	~�]�����y^���5�gzdZ�	����+Y��*l3��KVҙ�[�ABt�R����;�[�Ki������z�
�*�S>�|62��1a׵�����T��oX�:�z��s�Syx��;����e0.��c���k���u`�b41(Owڮ�S�^���+.�8�6c�z�q^�+�gq ���S7��M�Kr�����-gg΢�r..M��wY⋜����v%��oɏ_NW��+z��<��Q}&G�J��
�����q<&�&�c�������T�Z���VxV��?|�Ľ���ܔ�L/�B�=�]S��O��Ӂ�n��9_Z�v�������y�b���=��۳�j�p�z�ΒuƗ���\��T�;a��N���8���J��eoWE�8e;ʲ��,�k�$\�Um��wv~�7���Q�������쭏}蚺�B0�Z�_���I��Aj��}K�׵G��������a�tr�~h��a&��f)�7�g`ɽ��N��_goA�^���dq�z8��g�����mD�1㸏��o�=����{�\*�8�
\u.oT~�$����7c6�g'���O�X2���j�!pU�p��)���鎣��X�l}$6H�J�X1��ewbK��;Oa��:�U}vF�f�R1�����(esgys���>��WǾi�"���F!e=�{Aw^�+���y�L����BO�^H��!��Aq��w f莫��Q�-H�p��u+��&�;����a�g/�}���>�=6iԀ�ߢ�l�|���ڪ֮_/��>bL�4�qL��Ӟ�c5���ٽ��o����N�����­���g�`=UE*^V�fo�]�b����6j/o,'b�#HDv�vF�s�k�%�vx_���1�O��/o_�gO~+�w;��5}2LY3���"��B�l��&q��e�*{�p��z��*LlKY������	�!0;���ٚϽ�U�ͺ�gC��6�oo}Y�}��rB�o��=�*��ɋ������v���)�6Dֳة�x7���c�(����}a��"^7q��w�1�$c�~������倣Ww����7q-���>d�X��i�.s�-&����8;Ŏ���r)���y�17-/<�[t��7f�6��;^�g�`��x�(9�N�o��vk��?}��^co��J��~�708��������B��W�fh�yo�H55�gw}ԫ��;�P?kj��,+Э�����d��������mj���t͖{,=[0,yt�3�t�;��;0wF;'#k=� �B���u�}�G��,���g]k@R�K��.|���y�*i���L�S[�E����R���[��B��$�	�X�z��yX����=�W�,GZ�4���&�G�g<�,Κka������)�x��)Ҳ��]��#j�e��=ϑjDp�	��&�ʈ�;dhΊӡD�	ҹY�.��D����V�n7ޤ� ���=�r3�w(�I#ac#���Uon�\ۮVE�IVۆ�j�v�0G��V=��5թ��ʇn�E�ʭ�Τ7'i�y�w$a&uZx^Q�^�1�����t1�&�)J���.U�Veؽڶ�Y[͗dm.а�JZF]l�7�_q#F���Ò
��7�LjIb�
Ξ\�����v'o�P憋�e�r4Fp4,Ó��z\��2A�ԣ���L���B�g�\+ŗ����٧��޾��ۙn+�Q�]�*>�ɮ�nﳳDûBD����Xvhő�<�¯K�#:o�	g�Qç�ͷ� z�LP�R������En,ֆ��5��ۦ�+U�`�]�1�)�i�V�JS{t�Pqv��D�%���}�y�i*Igצ��hmk��r��X���e lL�.�o���[�B���B�rҭ��.<��g�K�7�M&-v늨�7��g_6Ҿ�I�$(��IBތ�v�	����7�N�Y��x'l�\57d^�wS�yQ��R�F�_�P����O%e�kDV��ΰ�xXU�7G�N����3F8��̳O����j���ʿ��K�}�Փ;�,j��G9�*
� ��G|b� ȧZ����%��An,892��y�%g�vv�ub rW[N�v�G��O'�Jl�R���uA[3i
3�s�@'�mj+3ζ�����[}!���{�nF�>{��e�Y���^NI�eց��}$+��b�u�坮����v@�W]s�\�x�Y�
�2�G@{�; �N�9�Kyà��d��q�P�]�@>����+:��-T�6qE���@�geg��Ʀ�lT��k_��=0�X�g!�"v���s�k�Q��nd͹�' ��ܔ�tT�]�)p�{�d�wrg?�ӊ��\�N"�1��C�;R�������s�����3�ò#�oc�N���`A�)ڶt�����/�\�������oX�W}c��=�����ٮ���'w�W��[�r�HO��1p;6�1�1f׷gfw�������۹�&F�Mӵ��r�x2Pla߃��c��A����K��.%[]u�w��zp�"ݨѾl��A��ىc�޵�q�R����E�-�î,�3L��oj�"x�r.�/l]���Y��w�y�G��<@���a���Rd!@d�R�4)JR4�B���`�%)4)@9RR�H�d�1�!Y�@��%!C�B�� U1M#����d�D!B�I��@AB4)F@c��йd�.A����.@�*S@�RB@d���IM)����AB�9&�Bd	��HV@� R��efACHd�!��M	��#�`9)�d94��d�P��K|w�y��ƿzf�vnP�.b�i ��M4Jt՘�u��3l���-G=�NS����O�4hJ�M{�^��O_�諭��3Ly-�ܘZ�}���׳�n{��q��7�NT/ϭ�C�����!��x�o%O$+|T���S��wdq��I;m`1h�������K�K5����5����T�L`�cgk�/\A�Qō|�1�d���~�{;q�����#�	������گ\_T☭������-�j/7��`��6d��M9�Z��1|,{���g��{0�ne�vU�W�;����bgt{r}4�&����zg/�;gl���>���=��{�v��V�s�{^�:�ϼ����&o5�	�ْWOe�]�N�E-'�����ղ�������X���y9��b�=5�p�X:?JW<]��i��C�j��Y�\�}C�����=���v�>�;��"��`�+k"~���oM��o�������}[;[��e<d���U��s�;f[Զ���s�͞}�!¤�yuy;���^պZ9�@�$Ƭ[�õ�N��/��1��a8��<�朧����M�Nᩔ��ᰶt�p��5y�c��������drv�����tL+k���0�)*����|>
�o3������뛍ţɨD%�Mk<lS�j������eIւ�M���昸�?O��Iq�)���͖���D8u���=s��_��j�v��9�տk(�Oω���󎔉�J�=m[_Î��W��n����7�rJ*�'�[�$��q�wN:�)�9�N�|�/ɠ�o-�{�t�����<�GC�i��V���ְ�'�y�|�(zl�Y��K*��{��<�V���հ�Yy�;51��d/}$2��A��+��.�?>���7Ҽ�;S���N{��N�,/)zEj���ϻ�Qǽ�k�W[�/ӓ��>��d{rgR+��9S~���y�@��ֆ��$��/z�Y^[I�c��!Nt�Rzog�^sB��>1���\����q�OӶ�n����^���$*x��N.s~�}�'��0���y�S��h픚ك0��5���QLs��)�qռk��In�J��*�~��)Oz+}�Sf��J;0��.0#��mJΙ9u�̉���Pu��X���\�z֦�`��_n�5:y*])7�Y���K8i�N�e���>��� �~�ρ�|�~<pY��*�+�Ǜ;���7ӌ�3����k �����AZ�yϚ.�Y���b�k�#��ܺ�;�N��������w��O���s_>��pvI�>q�0�D-��|GO.-wO>R?-�Įy<�=�������G#��ȵ`��|�;_f�|�=�e�P�i��b��\��.��ۛ]ӤןKY��-��\2��"�Dֳ��p�.�'3�-8��y\�{L��y!��Rdx%[�x9<�<ݲ��*մ�3�ݧ���PuwR5�P�������ܔ��0�p=���Ҭ�G:�H�C�ȋ�{ro�͟k�p5�&�g���St%�#h؛�Jz�.�t��Bkǧco���8�/Bєw��W�*�V��g�χ�-��:��͝������Rcӂ=�5l_{k�[t{<����:����b����j�]I�$tD��R/[]�pnX�m��|��g��'c��!�v=���h��V^������|W��Lk�*�b��F왵z�,Q�ﳹ2���9<H�y����:n�c�j��p�f�N��n���2�W��|nݸ��� >��c�n�������tLV�����eD������h
ؙ'aV�=/sud���fj�K���t������Ǿ��/�9/��6���j.�F��$n�m��)���;�¾z�s��bI7��_��{��s6��7x�����Y�n�/�N��u%�E}��Q�1S{����yx]�=��������fΏ8W['_���͝I��+��1ϗ�=7#����u���=3e�0���­�����t���T�}�����e���o{ύ5��'b�$iDv�vE|7��\�i�Mx�:�qy�����������?w����9���1d�M�+e�Y��pU$�ܑ�{��*g!A����H*O9V�~��r.QK�t����05t;Jyy=v����g����)��Z�R�s ��ϥ_l�Cj��	o��R9�\Y��f��]4i���Z^�9F�iU�uc��@)��D�_�}���`tF�QR͢���LXK�OGN�ܧ�d.
Y��q���g;�7{�l���j�lqR�,q�2��z�\�w1pc]n�����M�09=s����ϵ|�Kh�Y�_S�h[ܿI�����B��}����3�(��ev��~��:����������K@h����
;�g�']I�U��n�ɾɹ]��k�|�1�8��<��4�d@[�{�C��	�y�l�.�׏E��{s����k��8ˉ��A�������c��c�	�����&��-��Rj�b��G��=���Cy�f]�^���S;��y� ��KsDI
~7����ǯd^�_qfG~���[�y�{㷁��5n�%�s@}������ƣ�v�r���Z�+.צ�mN6����>���}����^w�)S��Z��{̳�WY����&gv1���NB��Ԟ�4�����>1��~'g��Q��+Gd����rz1�B���0禙��f���Ζw��ص}Vq���i��Y�c��R��v�q�}øf�{u��F�=q�{�I�9à��H�/S|��#V�wy�s;��_]/K�o��}F�W��p\�	�ɨ���n�Pb�x;��f����6�&�����$����'��W.����A����޽1��x���W�rr��z9�<��V�}qWF|Ӟ�_��\�>.^�t�[��w�&�X O�����P��*/�����?`u������;V%�~tN����Q��Lwd8�� �΢�Y�\����������f�B�W�Y�vA��`仺��=��\�'�;h����u�olo�k8�򗜵ST�>�q�ƪZ�fδ�/��EI�caeEk��J��E� �������ŏ��KZ�ot�ц���ʒ�Ppݰ{���>�:�$a��n�B��O��=�5u�_�,�zsϗ[#�m�yt�{��uK�ȩ`�]u`a:b��R��^;z��o[�uJ�Q!x��<L�{�<^����]�8���):�R�Yts7!P���nj��Nמ�M���^�5<{*��>U,���<xd�s� ��z�½s4[���u���k}}�D��U=���8�O��'=���p_�P�\�����Fp�6��n��;I줎�ӭ5;E���maLرDg��g�x������(c��L�-iCX����!�N�ey.�=8+J����r�4���7�9���2�P��X�N|O,n�����4�l�c�|��1�)1�M�"�S�K_����t��{��5�r�f�R��,������V�kB�V`Lt���J^u�*��V��[�뇯uoG>���*
�Y[�Q�<l�Ҟ�zE�>9��+��h���^�s�p�}�gGi竤(��%eez8U�Yk�':�cS�N
�#6��CB�Zi���qܞ{�;%,[��"�k�J�~)�}wp�
"Z�$��d�k۩HJ�B`..t�2��~���>:�ܺk��;�8��(��V��W���$^jJ��<�ڝTd��,�{7���G��S��(�:ǫ���YI�U��}b��2ڦr�Sk�T�x��g'���n�d�ޭ�`�˽H���3�<��ETd��F�"`�g�:Z�]_{׊�+�Rs�N�;�e�ꃯ�y�KCHC�~���:��y3��&��t�$��������zm�uj��D�;:*5�<[��+:�3���U���~��2�x(���b5F��l{Q����w�yz�6O���+F���9�֩�gXf�/��������YU��jR�؟����^���:��c,\r��l�&�'6�/���g��凚��|/}�7�;<��}Y��"�8�<�A]g,�`�Lc��rT ��Jgn�{��Z�GF{��w�!O;W#�v���k����n���m`�����U�h���>^���᫷R�T�ȵw]d���xL=AjN��VYo����ޞD���]�F�u��b�	ҥ���D�����	���U�
��B�|��$R�p���z�|�7��m�`���{^x��X����҉A�&I��.ޣ�^��V&<k=��Z|)'��6����ˏ���K�N�y�����<yjEyǔpJ���>�i{b���t���o���i˿[��Y��Yk֨@7�0q���<�JϥE^9����?/-��:ջ�T��%�G_�(�o�<����skϳU�����;e�>�"�*�Hd�{���j�1e.�j�i�϶���B��6Z�IXxb倿��	�/x������3���C���{uwS�|����-U��gO�(��#l�E`���)pNW�0�&������{��f�w��s��1�k��L���`�p���W㴄�
��ȡ�(�V�铛.�L��&���}3{ɏi}<����i���ާƧS�tz]��Y�Uq�9�����z=<��2jY�r�r:J��v�����5�ۼ[a��;B�m?q�6�z��l�#~͠�ffq|R�������w�vN��K��Q��a�]�pEv�s��G6ν�a�Gr�\B�3�?�Opz�x�`Ol�:U��n�{Pv�ٺ���W���br�~c+<���x���,<���|��z��&r+��@��7�;�F�y�W��"������a=�<e
y
����iϚXγ��!��;�fP��]��ot粪�Bů�1�Yo�l�"��#��'RA��O�L
zV���U��X5��[h\��[QB|ʏ��+u���C�UWJ��-�-g��n�9�"�Ѻ{�y���]^�ܶng���2Xc��|9ۇ��Mւ�B"'+���5�N��P��mv;���H�=d������T`����)�:��L$�!���kE�U՛�IC|���N�xgf��;��:x�Ǿ����*��@h�*
��oj��%��6��{PY�Z9�å휆�z?a��my��i��g%��>+��2+�U`����+;Y�	ҷ5Jؘ]����{w-9[�S�u�WYv*��V{.3ۙ߳�ʀ�u��#�_��o�!�9�Y(iR]���&��glǂUa�kY�m���`����ͤ���-2Q����Da��ʧj�@/�����*��n_n�ǔ�Q啜�P͜��ϕN��iOMȼ�z��7碩�'�_`���lc��Hʭ.���IY�omPT��W\6��Hw��_Y�ˆ�qs��v.Ώ>'��S^�"}ۛ�W���)���8꯾���p����:��nK|e�Ӳ��Ɲ'�غ���_�0ln���z��U�����4u[쓩OG��OF�0��?P�$Q���z�Q�@6mJ��C�,u�O����;w&ǚ���c�ɟ6X/Ř������9�o��qy���V��`�j�ȺI�Q����z��z�`�hC<y�O�ƪ�'Y�^���_ŭ�,=�'X���Tz�Ņ出I宏I��Vц�󬻾/�#��l�q���u)Osɔޥ�@�"�o6aЕ�m_eo��K}�]ﹳGҨ��k���X�b�3��g��8��_^�N*���?d^��z�d9���rY�}B2��^\٠��>%�����@e����F������r�4��:�m�}\$�/,����Z��R��\�$�.�*���P�Fϯ��ڑH��-�t �4��-�i�J�m
(w&"a_I�ı�����n����������s
U��m�ttF��aW�Wy�>�n����bF~7Fw�U殝ay(�c�cu��`�!��y���<��F��
�JD���ʌ���md�@GP^d��OH��cw�ؙW��q��.�0Zh̑���;��* YA֜��ک-ʹ�?��6�i�Q�������@��T-�=�����JE�[���	cgf@�U�Dq1پ+<>wz^r����sr����X�岸,�N��|��"dQC��=��&�b?�,�0���
2�N}������5�HnnXec�<�aZ�Q<�ˬ�	;�{_�_m��&��$��u��*|]����FH�!5�\3���;�F7o�F�Ji"G*�]�����.Ti����^��{��TH����h�6���E5vP���}DOΛOM>�8��b�I�bm.w�Y��K�۬��t�f>E��	�z��Gbc��q�n�šr˕}I<�)#�	@�C���n�y-J�����][L��§������#��~�!�`���4/��b7q1�7���:ُ�{f�zТ�ك�,�{+�fe*��\sq�Pho2ƽ�����\��G��t0QSݑ=A�������%=�����he��	�kޓF�.��b��Z�Y����l�m𬴻�ԉ13#u���݃�!�iiH�L�T3�gu� �I3wY�된8��N�F_A�Y��g$�k��w˸ƹ`r�}G�k��ؾ���`�\`�%�K�|h�;X��$�M����A8�ۂΎ�i��
 �{9��]���-wUX�G3��P]Q�ۥ���� ֛��P�4.˖�,�8��V87	G"�_W�4�7<���滁������u�*P�E�f#���Z,��W:�(�W}�R�*֔a�R�`��H�F<Tx��LvM��Z ����c��n�d��K��
�6�q�y�Q�:gnn�uMY�Tʹq1���e���5���Ge��ˋ�u,tʚ�L�*� ���V�89Re�ZJ˒��^|�ѿ������^m>���85�m�=�d.�Z�����>�mi��5�`��^���%���`�,T�W,R��j
u��x�jT�u^��)k[T;�i�9˚C=j�YL�ˏ��9N�q��վ�Ɗ���p\�~}\�4Ҋ��w`��a։����zU����0���K�&N�R8�����y窞�b.���k��ε+�jS糾\[݉S�B(����{��o2i��ۅ���.�+a�e	�$�?h�{/-�)SG�N����6hm#�ɽE�>�i�L��T|>ݚ��}]k-�ЂR�:O�ʈ�N%�{}�V|F\���F�����rcx��v���$�4ݑ�*Ïݵ����uu�{pw��b��׸�щ�[ۅ�7���نr�,�*w-��n�ُ1��b!�-s����Ϛ����	��#)M�bS+U�w�+Y��&F]5�ūm׷���μ�������2�P�JG##%�� ��(�$"�%����3(�2C%,��L���%2��
r����2L ���"����
���i2Dȡ2��!r\e�i����,̒���́���2�L�0�3��Ƞ)�!
J��%���Jr2rT2����(�ɨ�J1S'&�,Ʋ ʢL�!2ɣ,��ʨ���&��r�¢�C,�#0hȥ�\�ɉC,̡l�Z�i�F��r���r(2L�%&�L�
 �� ���>�4�)-ě�E�k���F�l��<.�-�X����Y���¸�H+�gw��u% ��A��n�w�q�(3�Wf.G�o�慎BW����'��fnמ��^�T���x��9l�Rf0s�,��q�6��|R���9��09��]�v�m���P��׼6&W���x���5��/�A�2>��_	B�s}�tο���jq��}+U^tyT����~��q�D��T[��k�[=�z���1��HM�zjJݮ����Q�Yu���q+)u;u����S~y�����\y�	��{k��}YX���D7�Ռ�W^�0f�j^��/}���mh�ʹ�i������%���S>Z��Jex�)��;dz݄Z4��6�������?����+P>��͂ŀ�X����u�5󔾷9�\O��S��Hu�y.���۩��ׄ�F��K�Z=)���� �p3��R�P�\L��8�'9xu۷	<;��q40�l��e"�t~lt�w�&�b�F�ӷ�P���Go�{cW��OV���=K��*�E
���v�'a��S�����s�J�9V�E�՝.��|�]I��;;Vϴ2�q�7��;9G��=�hUb���mS)��0Sܺ��Y��pՈ�P��ZO/�$�ہXg�e��]f����3�t�*�җu�:��X�d��NɅnM�u���TUqw.�|,oTеgq�/C�n�V���Po�$ȵβ����S׽H���g�x	a�S.���X;A�D�` �M=Ae-O:�z���E]�WT��"��xmq݉螛�92ɇ@�l�D�y-����I��=6�ǣO�
#�'�A���I�_������k�2��(��`�p�f3�d��8v��՚�tG	�K�%
}cއ!z�&:�0�&LҒq̽��V�������H̗��@��2bu�I]������ª�o������!�*,2����MT�<�{!��w���4�K�R��A��*,��T�U��(ͮ�F�����=�s�EmcUg����,��j�����D���I_t�|�X��w�z��Zg\C=�R�TDd�W�x	ބ	�S�tևb����D�Ƙ������0��U�5����9QZ�|�10S��|��m6)ygn�n*Z�&�ok�@֡�PÇ|�uX=<���p����-�Sh�+�kF��{��n�7但D�a.yxu��;��"����[���\,���{i�e�߇�jwG,���L"+V���� ��:�UpT��«u��<��㙷���%1�2����Iٽ1S#6Z�%��y3��>�����>}"��[�R�=Vӏ�dvs���;�@C��5��J�[4Ӧ{X7FZMpf��n�ĝ8D���Ȼ}y�w+��ք)�}�0f�����|.J8�	/i��5ol�o�����ە7�ۑ����)ԇ�y�x�E�+�*��ޘ��`�˅�Ts�1s�'���&��7ޝ�7O��zEr�����^>GH��)_i=��������(��w�+�?tR?e�v���nA��5&!�#źX}J3<Mv����)v�hDۜ���	x����r|���Z��_<gJ,��;(�����U�S�g�'N���TTj���jf�Zpn��^r��Q#(Pӧj���ɵ�w�L�����U���1D�*�{�^)�Q|7����W�キx ���>�_W��;>�=6�K�ΜX�p�^�8)�U��]�px�~�70����X>~x��;���-hJ_v�J�ڍd7�w	3��~���&fi��缏�RP�f�����"'��UB����-r��UYja�
�7�A)����ˏj-=e⃵�5*S���p���U��!\�s���-ӆ����
)�r��7iG�U�m��MF9ku����5��eԣ����\Vc�������Xf�Q�HT�[:�������u�ܥ���R����޶.�.)���3�)����v�Źef��׬�Kfp�;h-C��V��t�1�^/Ֆ�@�S,��&���j�m�I�g0��_{��[���ϻ�
��CE*
{U��'Wԍ�ch�=�𚮩�ޑ���)$�+7ۊ�����>��S�����<%agk>����{j�v����gr��q�#��G7\>��{-�{s!�rF���!{<�:����Y��$��^��)F�V�_�Jsˎ��W��h]a���m'G���E�Bn�:zi���<�矟�_��\��c#���żl	h��Ä��8)����o�}�/��3*���TX����o;5u��QyC���8#���"����J��j�C�s�x����fO;\�R��;�X"C�N1|e`�����T>w��6��;ˋ�/'MC<{U�U��~���\�b�����Xj�T�^veLUP.m�]oP��؝�0iZ/�^4N��N����=�ˆ���Q�:;�IW��!X�X��a㒦ׄ�HO5a�z�Nz�~�LJ�csX�A�"|Ѱ�Ԩ�U���1b��cH�]c��u�鷮�g>�1�z�r�T���_Vk��aҵ�0j��]���͉�7<=W���.La+����%���;�M�����\o-��WAi��`GY�t�p:�W� op���Ox
��� |��̫���՚"����kf3]�i.�Z*\��NP��D��%_wu�9�Mx��L���ʙ$?�{]U
<�;'R�&h��Ck}�ʅΜ6�e��˥��z[�9�+	��<3͇AP�_�~�Ĵw�I��`����¶�/��kR�f}�t�-��%���:��*�n\>و�`�$P�^�y恵G~,^{;�ܯ��	e�7]�	���l�u�ɂ��K�A�JI��p��bS0��/ӡ���׬c[�s:�B8|�6˥˃Z�n�pw���7_��P�g�r��&���!���Q,�1(po��S>�$a�E�{+����=u��"V��<�s��n(�H�h�`�x�j���7.�ˬ�5U�G�K��-����s���I��7���N�����u�H_I�ν%�3kƚ�s����N{iޑ��Y�[7�k����ҽZb���-L��1b�����=��O��!�f�JJ>z��L�_-�����+
�ǈ�.��㲥�9�2�|���zE�(�0X�=>Tx]�,�t�'���ۃ��|a�$~Ҟ�Q��\;��y[5�;	��Ӄ��b��jӘ�P��%��\[Vom��juլ�o]�0�ݖ�{:ae�{�ȇ�FQy�4X��A(�K���Ԡ-f��j�\Ң��@ų�o]A�����|꘨VVߗ�#����*�$�&,_�h��ͣ���`NzW��8�ݪ�tv�j���3y�{z6�@�^����&{�w�`Qk�W��Kf��R��:���^�Mi=��\�^=���^�=�HP�0=5��*Q6O�:8��ȭ)���[RU�e�갗R:Jr�n����oO#Yn�J��s7W�-���ϊ�����v�'<})-��x;F����S�{�'1�ˤ��������^U�A���h���E}��'x̑�~�Ŷ��{:�w���C�奕�8�ץ�C�U�!���>��ɖ���L+�ɻ��1�g�?8�osݘI3�!\����Ͻl��`�*�P|%X[Y���������˙&K���x��Ӄ�t�c%��%���ub̕r�~,���L�����~��lYٻ���<�����tA�ø�x�zZ$����a��!�|9t��l����.~w���=z��Ԍ�@[�G�ߤ��/�$e��Gе��*��r*3Ҕ�z�W{�r衦`��X�nm�v��#y��������6v:��`���&��+�-�YN�����e�.��|��2Ѹ/h��x�r��zV��kֵ#j�0o�q{�p[7i3���:�*�������Bn�������e����>l�bA�(�X�O���p��-�P�d�<�&w�z�ϸ^�R��#�o��Og�l.Y:�ZD���͵�^|�ښ�kF8���t�����C=��x�io,v�d��^�}�����kԥޙ�}Aw��[}�ǂ�=*p��q0�u�3��\�| ��M��xWz�wC0�8Nq�I֓�qJ��z
�z�o�C'.�dR�`�P����{g{����������0U�Vl�Ƀ�b��HcD�%�����0��W�袼���u黎a�xw���%qōg��a�h&�NT�1^�\&���#oe�%>�b�ry)7�_����5���o����V}2�@R�����#n�}�)�ִ�3�D�|�z����Gj���f�vQ�y!�wW����=�D��B�@F��<����\�Y�L���${� �!0_Lg>��������zg;���,'Ny�����{�e{^�s���d�w^�g
a�#�-w4�ic.�MC��y�LR��*����Y�:G�M	/-'L9wQu�ٕ��o�⴩u6����T񳚤���ҢG��]L���*�[&ڂϻt�{��G��4S;@�V�oZ.e�T�G��ۇ��D�"%*�R�/E#��Xy6�����[(2y���םn7������
yt)��|u����ׇX=]5LSҷ����VK=C���9�[�ID��g�b�Y�ږe��5���XMJ~�({��7�G%t�9�iNG^��/s��yVmA�=��
�΂�B"#x��_���T�X�=Bx?��y��װ�k��S��]��5�ʔ�\h����
�z����l5��B��竺=��o7����2��
�$�������邩y�4P�`���Έ��P�ˡ�6^j!d�r<'�ӝ�kޡ��~�.�F�^g�Uߜ��6�oo�uV�+�(xJ�����Ca�5Om��W�g�FlǂP��U����zV{-���y�:�B����S�Ẕ�T�2,`H�~A��K~��X�t�����������L/��2Q������q,]NΓv�G�6}ܑ����G1�L�mp�u�B͒�b8)����oÙ9n$U�e��WA٥a�g�P�ũ��$c��A�"��g�CԮ�*�/���E�u>Cؠ>�Y2R���^���gv�;0s�JlRi�Y�������=�4�r�F�u�w�^<��cy��N�d��0������>wڕ�{`��J�B8����u�௢GK�?P+�/ȷ����x,~�i�yD�q�a���ܕ)�}{2�����D<h��p�]`�,�mN�|�!�6���.<k����z�^X��������2�*��K��b��V�J��fTɪ�+��V\�22u!�/+!��zMi^g�gfV�u�Y^�f�(�8I"hnޮ�C��=\']J_O5����7�`��]�^�4٬�����FƠң{�E�k����34��;(g�x�m�ܪ�8�ۯ��O��ř��<W��gg��ʙ$?4���P��^X�b�uS�W��xOnv��sd�c�4�[h�E3� u%a����<2$E; �_{�ʤ.�Wd��+�ܽ鬵��vtk|�Ko�L�<�C:D5�^`�.�0�~��(w>����#�y9�<t�{ܼT�\"cՁ!4��A������l�,�JP})&s��xg��;ٝ��Ӝ�wx�w9D�<Uz��e#@r&�cW�Kef�ἡ���w�["��1����=��W+f3=��T��@9�t��]h���@TRVy�ww�c��V3�+w�X�q�h��Zõ�q�\Vtѕ+�s����{������f�sg�/�s·�#c�BN��	���-Y/3������r~kX���*���t��u�h�ڭN���[�n��4�8��}����ת,������q�8�ݬ-?6_k���,W�܄��w�a�|:�#��0�Q�R�Ɋ-�H]R���y�����m�鹋��P�x���P�6LOMzK�]b{.��t���`���V�](�V-=��g���}������*�q���������Μ�6�}W����Qd�q�מ���!�2,-	@p;*`Z��S+��)�`�B7�D0��"�{#\��~󷚯����0&6RZ��}v�6�Ņ��}�g�V�r��9��x�{���>*����ߪ:�VPT�->�`|bKG��=^^�_*����au���z7�"�}�k=8%��7��w�X��72���Ӌâ+GG��E��$P���>�]�+�k�~ט�=3��k�2v:�f���zTFơVG��mWNʛ�����eN�0_��'�dC�<��Izmf�[ԏ�~�<s�Xj��.����`!�^֟��Fb��o7f<�� �?}i�P������V4��9��"�Y陸9�Ș`� �����W��`Ψ��5J�}F��3�����i��b]�7��gtMε��dm!�tK�v���a��P����"����X�ʄ�{vf�!%"Jl?m���AY����2{j'�ü�,���s�d���9��6L��Q�ۡ�����j�:L<�oY��t4z�l�C�]	��P�>���ݜ�#+����"&��*ǰz��̣k
-(�����ЭJ�yQ�=z*�G��#9�n�������Z=s�*���-���5��\�g�)z�5�#��5]�vXn�K��(3Q٧6�������-x�S+�����Go!���G/��ݒ���+V�w|8�)
��]`0�sP�Vf�G�Xv�����GH%�Y R4C�=��,˂����ȉ��tn©p��K(�X�1d���Yf�j����֐{�t�:�}	�!�)�܈�V�[uգ�2q^����`�(�ѐfo}������?nF]���j��tvh�69��K2@6��Rks����1Q�f1a�s���\�}/V�&�c�j&�u�K��Z��9��G4�B7�����c����,�Z�ya��/�K�p���h_����t������Ч�C1D���V0	�**�1�N7�3P���&ؐB�X�6d��4bj�z�]����sMS�N!� �Ԛӏ��2���H����������[H��6�A����>=��Ԁ:O�����ֽ����ɴ5�1՘��̆���l��YH��(�lB�N��aRf
��o$��JP��B��y�-��<n��r�O���ҕM֔��ro�qVX�h�H����fu��9����j�U(ilF�WE���4e��bw=���b��mZ�PV�O��J�v�fX�N�d�ǡXKfj ��pv����;��$7M�Q���ț	/p���<��TsT�u�qV��^��q�("&�
���!�s��j��t%G=��6��]9��i����.$��iǯ�{�tV:�5`jto7�{�	����/pw�Eg��D�������� ����������}���T=�����թke�$�̖m�s�Z��$jh?I�-�3�Eհ@�\�9.��H�V9��Ƥ�b(L̔��:VYf^8:�?A�-LQK֍����6�m�J��ڼ=�6�|c�'`�Б|����I̓y�g�a�u�����'�פ7\�5[u�+�~�H<�W?J9J�ė����LĦ�ѡ�w64}��%��^Ճ�:π��0�kc3�EC��>L�w�n^�634+��ٛ��0v9�w�)K۰�fp��j0������S	9��{/�ejP��|�ܛV�_}�G"�@�g)�H����0W@o^F{���!���;���Q��{P�բ��;�k�5sau��8�^I�iͤ�;}A��e3W�j��,
%����u�?A�(���*�k$�30ZJ��,���E�*
UȈ�2��2����22JD)Z,ƀ�"����� )2����
V�2P��2F )��r+$���)�"����2B�'!l�(��F�2�&�J�3% ,�"�)
�'&����h���2b�bZ 2��� ��(bJk#%(ZȠ0���r(h�"h)���"�(� �
��(i�!�)+!�Z#�rr����i
r� 30�����2��+�A��$}�����m,o�|��P�e�/�,<&���4�{P�/�*�����8���\�E�8D��聮$1��9Ұ��V.~E�c�l���Ēh4�C�{��(<���t�y�����qK=�Շ�3��Iy}�� ����Z�RXR�:�@tE����J����~ó���֏�δ�X��wr�aΧ�6}�q�YU�;k��2�:#O����@��U��|����ׇ���;L֯۷UަTi0q�$h*K�R�A�yQep���_o�ǫ���@��[Y�{O|��+��lwEF��0�,�D�\Ic����Й����[Pmf(���l?r]�]�]x�V������2W���*x;b����B'��a3|�Un�x9CF++5:a�8)�fV��i�	J~����v��T��j��J��}����gvf��G��W�y�y��f�����n��2흪@d�P�@|눁ޡҰVw��ʥy�/�p�y����_��������6��V�-2`��\���J�RQߞ�	7�]�H����
y�&�v}�-X�E6�2WN�{��R�#h.&��%�<-1Ne<]v,�&�ՂZ�D)$}uק�/��`3�V@�p�O.M%�t�ڼ�:�Z��ϋ}b����2D��.��Tzy�VV�7����Je��)NP�g0�+*�h�68P���1F6�N�swp������|t1���j�b�gv���[�6�5�77�t���mA-�KR��X9H:��ح��!���&��o�v�Y���`���|.���b�CHB=]����L�<�J�����.��颟J�<A'H�TG���`����,�x	�F�h#����g_V����^��K�:i���G�E�Ѳlz]J(�
x�P�}{2m:�t�ٶ s�yQ�����fMsDT�����5�E��ク*vO�N�6��=��a���c8��4�4i�C�(�6=���PWi���K#�bZ�l	��~4�4i��R����Q�]��t��t��P�.ɸо���M��B�����T6t�B`��&�g����fZ�x�BKz�ٜ���/b�#jC�Ռ�jy�R�¼�U��O�X2�&�^uH3�s�<���O�|\����"~̞Ƚ>��,fwLHy�4Wҡ`����d����[n[���{vu����#Y�:��k՚s����=p浶C膓�\��f�@<�{��<l	D��S{Ef�3�Ύ/z�"��Eӆ�D�z��-��R.:�!����7����������i�.G\ᬎ�r5�o�$�;���y�`^��g(�Ѫ�k��4�U)���^��sn)�����z;.j�sq^\.�����������f�ɏD�T
��<	�\\.�t�����}� ����iHs>~�U1q��M��d=X*a����J�:�|�m:�`����	���N���w'r����e���9H��hd�i��� � ���u�%�=��9��0�og�����ް�62����2�jf`jf�<��E^�=��tp�L*�υ����2��}7����y>h"���p�]e�f/�������y�b�}N���J�y��o�/���k*���$��Chy@���a8�C;�5+��V��DY��\�؏?GW���T��τ���|UmӢ�q��Dĕ��}�F�u\3NNF�=�m�Qoo���5�w��U+08d/�654��U<k���)��ƑU�;fn{��E�-\B.7�4������<W��g`0�I�*��UB���B���f>�K����Z�yn\���z-�N��-��U���r�yx�eVD��}`�(q�U�����Q�zg}���ΘbGW�Żm��!�����|�;�֊-�����a9���\�w|�ڷ�Z7h�Cφ��J�]�"μuF>�O��V�&nn��y�Jݘ`|.V���:�ua?��M]-ﾱ��\ \Vo�ў:o�ˇu��̴������U��ɑ�!�����g�!��5(�ج��{2h��⺲�֡����i$NwXi}u5�$R��%{�N�6LT�����RL�p\<3�W��q	����n���n��z60J��C�eR:.+��G��/w�9���)-�^c˼�j]�=��<鳞��G�g�"t�#~�>���>!�������gګ�aoݔ�)gدzn�|��������'|F�"�}��P���Rʡz={�s	�o�y�q��Y���x�Lz���q�\�W��HRbzk�K�Z�ۖ��H�12���҆�%z����r��y��0z�Їn���j�.Ze8U]n8�Ռ�n5���ʲ�o�v�ׯ^�J=�Z���H�>���!z���2,-	p#���jfcJex�)�zK�x{{�Fߕ"w�{��x��`�*�Pܤ�������T�yJ���-�X��R�/�w{ҧ$&N����{���݇��:�V��Z>=>��>���3���Pβ[5���b����W�;��.����u9r�C}*^4���A}χ�h�R�����+�p�::��\����+i���)�������v�]�y�-uv ���ӹ�8kv<����_���Ŕ۵���{�5¬�K#�g�f���hyW5�:��H���k�������z���>u��L�=5�*Q6O�:�;Eu5�_�V��aS��;�ث�ϙ5>�C���Q�铱��f�����'��T2�:O
�'a��So�����C��}9>��4;9��0����xNB�~[ԏ����Xj�ˢ�]O<��v*=~�k��ݸf��W�<D�b�r��n竄�(uʱ�ps��"�6�e�C�.���2��K�Yi���;��I+�F��(X�[�l<�t�o�:E���Bmh×����o�u�N8�iϔL�ɂ�Ba�=*�W�٩��Y����8���{�-�w!�������=���c��I8ݕZ09�8���OM��xl(���I���^�u���,��6(��v���{��r�pݰw�,���%ש<H;�vx���p3	������4R���O��i�o7קK�yX;��K�s	��tN��OJ'<�Й�yW�4��<�wt�	��3��J҆��0��VV��8����Ɛ֠4Pq�Q~��d� (��D{`���%6EVG�,��[
�\���{a�](��n�w��3��̫�%�j��/t��js�P�WM�#����~~P�37&�gA�>ﶕ!3��'juy*<��L��lpdm�\�T1�"�2]#2�LMU�v`=J�sUl��]9>p��j_��i�۪J��|'�~5�K�+�ì�+U<Y`��'U�a�8U�q�W=�;����&��i����8}>Kp�.�ڥ��A���� �m��\��o�u����=��j����_����\ӕ׏Fق�/�͖��g,�9���rQK7ܸ�9^��[���j,�>�\����3�NT�i˛,v|���@�����^~֦a-�I���vj:��&��a8M���<�bc*M]Z#��l}-J��`;H:��4yyW\f�{t�����Uc����8i9W��#\�_mrߺ��Z�U(t��D�|=��.�5�~�5��~�1U��B9}TGJAD��i�w�XY���F'��G>�{޸�sa�����0G숡�\z��.�k�*�,�Pu��,e����ƽ[طr��f���}ڟn3��t����"ho�����N�$S���A���M�y<�պ<j�9}�L�5窭���*�7�g�G��s+ ���o��uH[�Zĥ�]@��kGl޾8��r�L/Y����f�w���91�9��i��D�m	K���ߏg�W�sC��c�1;�z.݆��v�̱��ݦ&bc���Q�
u�?.���v��+���n�OU��,�>g��R^~}��s���=>�*/� 1�u�E��I3������p�0X�⪡{א5Dt���J�!��[���vwթ�����!g�����3%��N�pS�<*u	vD/{0J�}��}��|�`�*w;,�����_]GZ�%%�ݞ�y��w�,�wUbS��OI����is9{��1n>��~~9ĳf��LY�3��0~G:�>��'d"��ڀޭ���<BB[��>��\�ǽ�u����<'J�����#�=i��������f�=V��� ��;��}6'u$�������`O��;y1�J�X�t?Ki��c�독��e�׽����ok{Q�у�CΏ�-3$H�X�����f-�r��N֒����p����z�x���,}�h�-L
����i���f�a��A��}{=��T|u㝓���}S��V�G�T�U�m�HX���(�S.��f+juC�qyx��G�]�<����{����|\��Q�<j��ULV:��	�;Ǚ���T0��5(9�Q�V},]`�Y�9<N�^*���AL&��Kiڽ�u'a��NњWw��1��������n���	�tua�,�[B���)�(ZA�d�q}�\ZC���X�nN��2��z8WWZ���+`t�b��𓸑H�uj�����,�;�^u�μz���/�:��l{�$��7�
ۧE��V]��+�9}|�4R���b����3q>��t���Yʕ������z�� ҭ��u�a|k���)���_��	�ǖb�pwne��&�-�a�� ˝{+���/�%�������e�<��/y��������G��u��^1�,;�S8�ua��=38�D��AS��ٻ�z�z.��++*��S_�']���L��<�:Ox>��+���\|%B��(�߮!g0�.���e���|`(�1�3Td�\�}K��>���f��¯	�}��鹎�o�^��̨���xO��:�$a��tlp����<�x�:1A�U�ό�f�R�֡���oNqp����O%�Cѓ�p7e�,���9��תgY#�YD����$ʾ�)!39ⷺk����ܾ<9���D��-�£���z��#~�>���C�;�^<ʛn,��~vz����<b��
�Zt]q�\�i|<�$�&'������B`�*�t�Iɞ���[c�Ÿ�m�YW�̻0Z����A}+y'ٹp�gBjN��k��b���LU��@Vbb�w4��c6J�K3%lKk��8RG�\t��2��x3����f�2̗�#��D��E��Ó' ��V�#/Yv�5��a��y�蔎=c}�W�K��UI^�o�a��.ZfS���]�"���i����\�/MŠQ��^�{9����~vQ���=U�KE�6���8x�0-L�waߋ�����7�I�w�U]�.��܈����.�Bc�Xϥ%ᄺ��J�Ү�����xcyS���ɤ�M��eM�>w�mzS0�+��h�{j���w�2I�������� }�q�M��߯z{7��u��ۮ��b`.'�ћ��sHV�	�d6/S���u+�$�Z��շ0�/e\�g�����lMF�������3u{�6%��m"x�	�ˮI��|����<��������3.�n�O�z��~�<s�K��ѭ���7֥0�w"�oS�1��(Jt,R�= �K\��	�M8"�Jע/��9�z��,ڊ�^:����8�ٲ���\��
�ɾwD����ΤN�L�%�y�wۈ�:�a[}1��^�%�Wbjx	��_L��G�t�
�~�Y~Gg#ŗi�ϥ5E̺o7l�רP���hծ����_�5�����[]E��p9���x�)�G�����A�8��lԖ��TR=����o/�N|֠[r�Ӝ��zX}�Ծ�u���ڕfp�?{����j�A��e2R�Yf��պ�O[��N���[e�M<k����rʭ�N��UUX:]��P^	:�؎�O�6��T�أ�i繜�d�T�让*�JI��Y#EHM���D�O��r��pZ�j����+�ĉ�^����p��n� Ԟ�cu�&�3�I�D�-��x��Ԍ�7ȥlk]�}��>�X����i3�ۄ{���pm��05+��PQ��W��|��٪�C	�}�'f7V������ֻ�10Mfu�Z|+Jd�Z�}��팕�T�xJ�Em�G;��n��䓗cd�&zWqu���v�{12��7i:�nZ����{(�x�I6��%��mG�=�[�u3�S�C�>Oe��7Jա�ʫ1_���io^3�?v�N�;�-um�Ě�qq��<fzi�R�=��'��F�P�	�s�.��sp��ct�zd���YFZ)y��5`c
Bno��X�ʓWV�4Ͻ��Q�5*׃����v���Y�wԂ����#�z
�t��aJ�9Q�y0৫����|"8��ݤ3�N�W��w_�
A�U��e����,js�!���"�Ϋ��y�ט9,N9|�;C}�p{���u�-de�9�6�+f�m䜕�C���r�R�_?���z._r2�{��L䩮��#e��]4��M2��6� �����Y��y��g\�3!�;�-q�I����h�R���}��⩈f�6�m���cWX�E��G��j|?/�(�1]���.�M�V��qV+�F!֮�w�B���4�v�R�gNð7SG>�Wٛ#`�{א�I��LWi�ri����%cȘz��&�w®�g#P�;rg�sh�Q�����;v��7�:�vA�Z"�����#�}��� X/E$�7η�[Ä=�/���LL� ���eJQ�vsZ�d�9�� p;�)���"k����X�jk;�-�K��x�u��/��^>B=��ܦ�t��J����9���o�H��'|�#2�o9r��$y� 7���:��[!��s�s��EN�wLh���v��K��Y�ЩФs]X��a��q�Ѥ5I�9;�/���!܍p��������ٻ�kv͡܅3��CS���En6��ѺC���[�b��p��S��2q��h�]�]}��z�?V��O�C��9�d�-fo�#w��:�]9v�5�r��r֕�-�ܝ��;!Y3��ٿGMP�
8w�-�!�·���ʛ#8�Y%��-����"֗q�5���c��䫺鵜�df��h��������M�d����):���r��'��M��0�[���ҭv�I��ʐ���w�p���R��X0��y�XH�m䠷���(�x�#�aqйۡ�Sz�"����P���w����n��&}��ʯH���eu�p%�%�e��r�#����w��L�pl�^��h��wE��xjc�U��g�їv�B3��لz�TH������!sT��q�:��%:Co3��\x�>o�fU".Z�u��90 ��.�2y�좐��+���-��i������b��UdE29��	ꔒ�}��k��M��}������?g��B̦�in燬k��kʠSr^9�H,ud���n�On��t� 70�euZ�֭J��K�u�u���-ʾ=Bm�s���ƴdT����qhn�ʕ;�nl�X��1Vx��Wo��F=H�J���˵43	�6�P��P"�U���X(�	�O#V1iH,J��irᡑ�4+�>�.��i�_I�K�6�PIWt-�q�ݲ�̙����AvgQN���k��|���W����$Έl`�K�$?F�����1\W6T��AѡZ�׽�M7D�՛���O���J���p�ZЧz�,�n�懠�D،d����vk{.1eӳC��W��3z�0�͌ҙ�'�ۆ���H��Z�~�T�m~י��}����4�GRd���D�4�LEP1�XTDIM�d4��!��-4�U!MEAAA���4�UDS���-%P�T�R�	IM�5@USPѐeKTU)KIM�VbRaA)D�QI)DY@Y�Y�X�U�!MaeE9�%9@`QMe�dPd9QU�eKABS�4LR19.@DQAUCIfaaUD�XIE9N��d�D�d�eX�ED�CY9!T���Yed��Pд��FfMfd9R�5KY5MS3Ue�MPDd�c�U��B�4| D���g���W��ʷ8��F��
�0u��J����I<y��;�wb"��]��
x��^:<Yl��Ze������5\����6E�p.��̑[����l��8������fo �s�����o��z�ͽ7���L�b��Dl��k�> ���"��oN�2���{���㷑6�;k|�M}��S*�Hj�򓦉|ф��Fo������z�x[x����Nw7U��B�jE��n^uzz�PG&\ʘ(=|�K\�9��1f�M �q{�n�r�h��	pg*;+u`b��RL��Cp1T#@�,F������Q������>FD/��qfu��+�|��kVf	xay*Ӣp8-���g�860ڷ�ݫ��\�z���hO)]>�X���=+@�|F`�*��ʫS��������3$�E�'�o01�XC���:�=k%5��Ϯ[+���J���(`��/��ي�=�tmI^�r����3꾽��O:P��D"�ׇ��9���g�ԡ�R0�ώx�.�9k������5�c� ��/����e���<�|m��X��@<W�����ڍC6Ҙx5pE@	��K���wZ��u/��%�]�����r/(ּOL������Ky��vR2ZgBbzeu�9�<��xdv� 7�8*Y�6Uޕ�쨢讌����x�lܨ�'��h��諗f���֜R�p�/N�<d\�lvU#���=�OJ7��8H��Q�dr����'��4�����]��Jtq���"�C�I�C8Z0եʬjf;���{Bl�ژ���ۣ�8���-l���*�����;�<C��P?-�U���N�g|-���c���wb���
~�_�\�g৒��������i:��3@E�X#����q���5*�Uc�B���n�%�ދ7�j|w�#�C:ĻcD�@�3��4{�>Ih�i
ֵ�h��2m��c8��V�|`mf>���<�3`A�,��4�h�Q.S�L��՜�&�E�ڝ3i�{טr��2^'6ᇋ9����^��0�K�D��������Xaƪ��.������L'�|},_��SCdi�x��)�Y�����3�xdO(X!�����X�is7��mւ�iUQų�w���d�L��o��)�g�2����lZ߳�_�p�}�b�.LD�,�ˮ$Ӈ��zxv�zC�b,�Iૄ��R��x|�QHq��{��5�_]<v	\��Zl�
x�9vVRW������wme[ӛ�u&�t�Z�<�OEJ��EKQ�ݘ�Ƃ�V5S����;C�"�t$�V�8���=Ou��r_��;�$ܺ�Q��/rV��{]�ֱ��56���0t	,C�]�|�Ѳ��t��w�Μ�WOy|�ƭ��e�)c��������ȥc�]p��'J�bP�~��Ld�!�9�,?>�KTY3{&���o������j�s�誫\+dA���gI�:*���J�#�X�U�F�H������}�C��
U�3<��޵(�8d�0�@y�I+~5n֭�4dChDwʞB��}���}��Ǿ��8�8��)�UI^�X`����r��?.�k�)!~�+*a�r�i>����}cvkBǳc�%|d^u�*�V���p;*�fpiL�\=��-������r�x��zP����&R�΢��K|dK�	sԩS�U�6���/H�gsm7��˹o|��dD����aUxu�f�G\*�&���Y�p.8�����F,ܘE.��j�,;��;�V���>'!.�����Ŋ�!�!ZW��2V}}h�u<m�a��QNoʹ�>�Ǡ\��ڒ���,OVM�3$�e?�������@~񼩣.���u�y2�Wkh��-�iy��2�m;���۫�K��U�5�;'�{�JA��F5���x�K9����pZօ���y�^��x��P�86x�ǒ3��V��cv˸�[2ë1I٧�]{3�de7�᝭��o��m����j\��8�>���=|�ݓ���/f�v���W��V�3��^<���F��ޤ|+���*����Z2�Y�U�V�L[�M8�E�B
@�f_�!��"�BmM�Yp��hq9��Ec�^%���T���_���^�ge���ȘP�l��s�5_u>�C���W����i�����Z�O+��<ft
6��22|���;}r�]X��	t�t%�K����jܕr���z��5��]�1��X�r{O�r�ZU��s�q��+�Z$��xl(���o��*���ۜr��G�]a�7���\�^})&9d�J��|� 󼪩�WW|K��\\�����Z�v�d�G:�\c�=��\D��1�.
d��d�=��Ƕ�v.�n7����O��
���hq�m&~[���������*x;��-jE}�Q�
�u���9Y�n��6�F����K�jY�ֻ��L:ϝ->�ɮ�Z�Ե�/3J<������MU{m��<�o\����^��z�<j�#峵Hd�S�f@r!�L�]EG5ouL�W�v<�!�����N"�t��T_Ң��_����9Zc^�̳���}}����-;�>(ٍ�ѽQ�«���q�]���h���\�B�q��f��td�|�.�4>\�X�=�s-�[�[hLj�v�nf�;���z{�[�����r�8tk'eԯ|/P�T�C6\.�#�wk�~�ǽXG��8|���T�i���s���A!��]�oz�0nޣ�WI��fg�E��.ab�H{N\�c�,���u��3���w"Q/c����O�d֚_e�+��
Bj����C���&T�����X��p�}���\wo�a��u^�3c�u�!ucf�<p�걊�z};(�'��	{}��yeJ�q�&���&�$��@&]�%G���(Uu�MeD�b�l�n�M�:�J[�3�����.W:-����3����Al����_Dl���0�8�+�����:����F�T�_8�cI� �9	s��	�P�\�e�Z�"��'��Fm�m㢪�`������+�{�#��9Z�<OJ�s���U�n+�2���L�����@<T:�꧟��P�s�ݚ�?���$�C���TvV�:ȱB�����
�*�re����fTT2,:�X�ew	���$������	P�bP���{�3���~֬�����V�৴|
��v�v
W��?k/�S�:���X��>�۴�y���t����Jب@�B����*��|uk˄'�'��-K��u9�U���퍽b�oػEg>
��L����f�J�`8��wC�"du�^Δ+Y:�+r7��S
gG_�I=�L���͂;�HV�@y�-��ӫRP{��V����`�C�#�=���ٹ��X��Q�>�H�eu�����Z`��ii�;!�ԁ^V�ڢR�ޙկ�5���B��s 0�ϫGL'J��Äak��U���Y�����i���}����MR[���Fr�pxe��[&�Ȳ'*`w����k
�>+q���]�u^n��>hq����{��~𾭚��#�<�f�G1�o�׽X&r��jH�)�(n�ћ�7��c���M�#�a&�}�-}���V-L�jfxF��e�ۙ��;��׷$������^*>+���ꣷC�,u!a�*�E���3ki��~�ejܞ4m����Jcױц|�/��2���զ�.�T�P�L!� �0�cU$�����կ�BɧyG�sP�w�gY�������zN%(�q"��x�$�y+VDp�A���Tig�u�G��{=���mvׄ�HO>ɕ�<�3�B�U����, k���Î3MZ���n��F����ZO��h�Ǯ�-lY8qhQܢp��A��2i޾�,�QV�feø5+a�']F��;TӁe���0�r�e^�Λ���%uh�]Le��K"S*؂���U�*�9^�X=�}XI�;U����5�7����m��soD�YC',7�b�9d:����E=�*�N��+�{������0�{Q:* b�v�t���L��24�+G�������-9�ʇ���q�q�ؽ��9���S
�$���	�v(L�'�"��<5�Wy\��<D��Ƹ�d+o�r@�,�0\�5�Z�Yߊ$��Һr�bA�!���lE���XT�v�^ӼY�\�6��{��uP��� �Z<0Kꘑ��Ѳ����;��;��R,7:ss���gsK|�{X�p^�`�g��	38�냖O���C��^��u�0�l�=�x7�޺��7��^<�K5��\��@�����ʕ{;�A��:��p_K�VFB����'�H����b�ғ
K{g�&�@����&��P��bzk��u?����O�y�w�����T�	�}�0Mg����C������.Zar����Q�u��Ԙr��o�ծ����^���b%f&=�>^u��p�����!���u(�;�8e������{#Z�+�
�r��C�����qȮψ[,Ow�-����%�Y̿u�ɺ�ڌں�T��,�B��+@u���:��-s����9>�2�s���c��w�Ul:歷\;6��`��Ѹ�fr��R��i�2�)ٚe���N+�;]��7R��$R�(����K+�gRc��c>�xa3�j��*��X�E���kn�_G}��Y�=����ܬ�<��fkdyh�{j����)����u�;�f��}]�@-Ѱ� 7����RN�0���2���
tb���zϯ]w���V�����R��{$^[RU�,OV}6�̓����T�m��bW��BVE~�����쎜���Pڀ�M���x���'�踦>��Wu�d/�[�,__�X��ՕHj�>�����&�$<�<�-jT��!�b��L�c��ʙϭ�6�/�r�irƙ�۷�s����m귏����g��9�ȘP�l��?q|E+٦�c��mN�у1T���'ki�9󵞠���iʊ�8d�p��p����DY>	:��[ؼjF4��n��&�s��w��Aܩ�gXg�dY0?	I6����
T�$�&���ƍ��|�<��5縲��$�}Yτ~,�oK���3�RL�$h(	.�H<Hw�o�e30efl��Q�Z�b^"�)+�o;z�y�վ�����D
�*��E#ꞟe�^�L��hm;ݷ|\7�Դܬ�+Xg&�ʕѳ��F�|kR�W����.�q�;�P��͠qWC�����D�%:��)e2�����
{}M}ޜ�ΛE򛣻I,{�v]//�n�H���7*eg��Q�>�0�T�tK��$mu�W��|��?k�vr��x��-hB�ecC��i3KO�o�=���:=>���O��b�e���[=�Ex��wAb�U��g��J�ۯ	�ط���^|����S)�]k^B:�{J�<��넷1ğ.��Q��tN�>��g�Eç���jW��/��i�]i;qJƁ��H��K�{�����r��gݗc�+-�*�|8����s��TB���hTU V���}�0n����5�r�ٙ�Q`�u��+��2o�E�B���!Rɏ�c���5.�	�#��-AH{�p����!77҇��bc*M]Z#��r�u�����ƹ�L�7ԣ6i�
�1Z�?�U������S.�y��o���b�O!����e��zK�y��W�����=��+��pU�2H�^Q!���U�XY�S�`�,���I��������>8��H-��+荓c�Ԣ��0�B����۷���dh%=�3�I�·I��S�'tu|�+�X���no/����w�V`��p5��t���/1��g'Y�%-V*M�f�7��
�M~�:�A*}{��k��I���m�B�Fk̔9�F ���\Yu���3P��O���1�3�-��ΎuH���=S1qzv�4=s��LR�����6Rt�"���O�N�1T�Wݶ�d��?#�������;6���3&���^b��r�eEA.ed���@κ�PTCQTrlX�N���wG*��P��ځ1�Gegź���B�gxT1WB�6��=�	����~��tm�xXS�UP�4�+��%.��κ���H{�7�)��sQvv�0l]�$ym�3�]Q��6"�����ժ�xW"��t�D��@,��Y%�����\�n�{��yU�:���Ž�Έ�_Qa��k��E��\/������/�Є�9?j����1�F�0�p�|�!�Z�X�`ϥagk>��CsT8
���~ϊ�2��H����!K5dw�[�5\�Ι���[���Gp!��r�I�v����cqj!�j��oܞ��gn��'�,�bξ(�!ڔsش�G�r�2D��}�4=]��-����^��Ǯgdۋ��^3O�7u�$)�갔������V�*�婙��]�d~H��Z2�\W�n���}����'h�iB�wO��6�-x��&M�B �m4/���x�o���cg�+EA`��8�:c��X���[��*��'B��VF�¤�,�us���R�r�Y���5hs��[�+�o���Bw�9 M�'����ۓ*��U�����+YO���V�[�¹���U�������v5��Ϭf=�.��5�Ғ�� l�M�447��7RռÍ,�G8:��z���^R��oWu6�f|0+�斫O�ǚGlK5B�^�K��[�M���:��5mb�T�XDН���h��1�_�e(g�
/S���)\=�Gwb�"m㦃���˩%�#�]m�����Q�\�n#Y]Y�H=e�2-|�򫒎��kAEu��f���z)�e!i�יb�iǨ64r�=_�`>����m5�b��5й:�<����3N�*��5� ��(�lc
<*a4�+�.��m�ZǦ��-c�u:���t^»b��
����]��P��k`�SjtDS�X[��+��N�9|��ԙ��ф����pv��G�>60J���1Y6�e^<��alG���m�ɢL!��/j�%hN�Y�R���m��V�h�����Ѥ�V��M�Q�Du�`/�s��1��C�K���lCg�2��q�������}��[P��1,љ�mJW�� �Gr.o�h�����oǽ�7�Tz�V�:$��8��⫲�7��T��AKh)��F]��:*�3����H�P	]�ݴy�����2���f��ֈ�5��3��i3�K�b�9aE`��;G���+\Of���=��g�h� ~]q����(��J�s}��1�)���k�p�>u�݋�1�й�}�����}���Y�!u�tpIeI,�sI��%�w�9n_g����x�R�ʿ]��_�d�S�E��Z�3s�<i�A�nIXl�swRT��M�#3�� U��%�@ZY����;�\�*��=�_B����/��(;&�F,��;�zw ��ҭ���ϻ��jɧV�\j����)ӗh�<Ϋ�!�����ʹ.͌�/[�F5ӗ�H�$�����3��2�qP⁜�EὺF����'��+�{A,k��S��0v��������q�K E#2�{�5�*��ʹ��Y�n��]�g(�ш�r+�L��3gs�p4�$n>07�u���Kfm[]a�#Ǻ�0ax�qm,�q����yw��bqА��2����Y�J_H��a@]#n��O������-�V}��B�r�l�c��H��I<�ޙ� �3�9R������.<U��v��h䩶uU�ee���60w(�V=�\DKݴ�Te�+��2Y�˚[72�k�YxiǕ�uv�q�h��ċ5���EʂZfGF/���}��y~��}��z��U�Q�)AC����TfdAJ�EEUE6FI���FHa8�%L�PL����K5UTSTdJ��SE)UE5E4Y�TSAEfKHPSEDNa�TQ%-4%��Y��QT,�a�MUY�T�E4ӓ��MAYaM�DY�I0d9P11fa�aEACUE44�T%�a��I$�QQTEQUIYffL�.A�AE%EDTe�f`U51�f9��AQ1EMe�TU%4�bKM���E%T�e4MN`̊����{xwgxq�fC�qUDͅm�EJtl���ˎܠ:�w�M̭ !���+��|�g2�]k�Ը�!���9ul�'U�ޙ���޸�Ţ�OM�Yu���c�B�E�
e�[N�$퍐��j��nV=��O�*}ٮ�[���Dh�8��%��R*�Q��<��d��;۸��x�7������9�
qs���1�9xo�Qf�(�Hm%�5��è�4��{q�	��>Y�eJ�f����\�%s)��B�iV���9��9��I*]��}K���[��2�L�EA�;�>�+'<�^˝{+�T��H�%{u4T���vk=�*qd�|y:t)��-�D1�F�J�����8�:���~�DQ�I��٘o����V��B��(P;)2}�<�]v�z*�O&E����/�����g�Ŗ�;�����*o+�:o�bj�1�(�5�q��r�bA�.�*J�T�cUfD�{M_9�\�}M{4Yݥ�9��ځ�h�τ��1#�tl��,�W~�J���hD���%�8��Ϥ������6K�Rf0p9e�q�LJ�YS�
c�{���V��q<��GU�(��Ղ}�OPz��+�oL��F�S`�!V(X��������J��}hYo���0��- nʔx�շ�%�)W#�ϵgq��oZ�z�1�p�Q�cZ�+���ۓ�*�m	О����q���_^z�޽�$ʿ:�5T9�U!�)	`�/mW�K=[�x;s���}VoA�y���@^tyT�I�
K~��*n9�Y�c�\�iy�I+~5���6����u��g��}�5���mFp8L	�=�/o8J�oG�SM��b�_xe�l~|��ZU���L�!~���U��p�[��f�x.�+*X��A�c�><vT��������[7�oGrf-����­r�z°�Bc�%��%ᄿ��	d7�����糹�0nX��Po#�Ց|�/���}����a�� ��Y�pv�*x.��Qh簞>�O��_��1�����o���':����T�d�9oռ#(k�n�߮��K�p%�/B4׽Q����uIT�F�z�Eӹ(�lL75�'c�`�s7V���nL ��K�7�K��|t3D#*�TUoT�u|^+j��qM�S��NTo�ָ6�d���Wx��֯{��E���**j�뻠~�$�T�Ŏy}t΋mF�o��_{�`���2�Ơ�^�Z�Tp�s[D�&�*�k���7��¯�W����K�6�EO�ݮ]z'I�Ћ����f�?FEҥ�%@�4�])l�tи���ɻ��8au�d��'���yW�̾������v��k�g}Q��a	)�x�{�"���Fd���y3�<��}0�7����a�_o���*����=��<�17Y���6���Jʼ2�����w��������	|��.��;6�V��yR�2M}6�#P/x�����vS���)!��Uh���`�ve��T�~�F'����|T�jd�u�]�ciJ��:E���"�B�RL�T4W�G	]��	�F�n^�75-[S޶I�=���yt�pR)v�e��en��s��#�����.�pa��iw�2��S��o��p\���	~����Ff��xm��1�]F�c�VH��җ~W���ǯ
5;�Y��="{.��յ�1Z�|��gZ�Z|(��]uj��q���aX7�K=�p���gB�/L�
��'�L���)[]^;��X��20Mfu���\����;��Nۺ�+��]�k�Aao�C'.�g�Jd�jV��o������T�_A+y%]�ٱ�?aU~0&���r&�r�}��N^�1ܴ':�md��<�0t��X4a����*�>*�A͒17�}kf�:��{/H���%�
�q���k����j��h�a�
��|���l��.���eaUhX�pqk.��3�ߴ���HN�"&u#�DUx���Ӽ� 3�7^�2E��7g���V���!�a�@ǽ�,}����Q�>F��K�Aqz���.�"�!3T����#�&-���>V�P��U��ru��T�e�������(��h]Xٟ%ⲙuK�1p���*:ۋ����"����yߴ#�
�W���Y2������Uq�9׾Q!ֹ�'d�xn��қ��[��m*{��g���L��_�e��G�&��q�}B�����K^�H��?x_<b���a��b�9���\}8��<*9�+a����>&[��ujX8�^Ŵ؁=��Ab��	�A��˚�)�Z�O_��Sq_�=V%�f��~�4;�h��k{��5��q��E@���R�pş%.�	y�Gep-�u-\/���=�����sy~�����7fa��O5d�$!��Y���J��4��9���(<:u@�m���%�m��{������pS0�"|�p��!t��g�IA=�g�h��1�zZ0hH������y�*��s�0�`�+�T�"u
F�<J��6����8��ע����jn犘/Z��GE�bH^��ǂ�.�Da�x!���f�y�K{E�����8w�-���{����"��K�^�0V�ި���2��ӻ8�:̯:�\^�Q�Yt��=��Y\q�d�y&vRG����4�Z�{��]r�ƙ�	z���E`�r��t��o5{��/uwV��!�Z�X�`��T0�+sT!��^E5��^��ʰ�9��i���B�/ԓ&_�b�������-�dY�����N,�xuN��U��޸��"բ2|~��^=�ء_eiN�b�%�LϤH����:##��:J�0���ћ.lj�30����3�����eS~�u6�BY��&<|=9�Av�`�{��6��[��M�B�r����S��]-�*���uP`�z"��[.���3Gn���Z��仙�V��ĸ;(߽��b�Gj�����qkEj�U�B>,�Ux2��y�[��Ƀ�V�97(�p����Bq����xo��N���K<a��C�V�c�+����B�[�C�C0��a��\���s��,2:#cPiV�;y~�J��x�d�29���x��<FW��|����=a��Nm�+'<�S/�fS0�UJ�I	^���~NΒ3n�]W>��^}bً-�E�4���Z;���8��{�u�/�Og)��V��K���;w^��J���2v�Tyk��:�/Z<}�ް��d�L��ҽ�=�ٛ&�!��L�VP�Sq(W,?z]�Q��O1�{����D�>���^s��M{��Op����i�2�s2�fU�g�i	Q��Ǝ:�y��w˓�%)y�cS+
7@��nU+�u���g��*���n���MD�ޣ}*ډ���a�X����ZYf�F;���Q$V��5E��v��*J�苾-ˬ���.=����aT�Ї).������1#�tC#�e�;���z���kH���[���a߾�Vi�G_LT���`�Yu���*bP�X�
�<r{�w��z���s���&4ώ�Z�
��<f��5T8;������$A���u�](�{���7��#�/I�x�y`C��,S�{(���fyOS;���󈚟y�I�e*��}8�a-�\¼����lu����͝�o�δ8_4c>�ɩ�W �i�v�k
�E��������/W~�"�/-���c�ܵo�n�o�f)Y��m!�2,v�2�B�ܙv�׭���/�Wu��cJex��Ok�^��2�aXU�LtK���0���}��m'�T~Ț�c{�a���X��R�3!��q=�Jf�b�+E@�g���]��o�����|�B�k�
���nXw5ª�e1�{�_Dr�h�Y��������a�Z��|�K��6v�O���y�c����&2�ʾ�ո���W�;�׵���Ye�.�aV' Q)A�ƀ9�܅�+�����	{ސ��ەV������<틇�I+�uOipi�n�#'X���v���>)�e<uupsd5��j�ʩ7b��	�o�⫴��1D��mITv
+���N�>ȇ3t�u���W�9*���As/�GB�m O�xvh�4Z.���M8fzP��j'y����;Z�}5{�
3�����T�]M*�!�O:�c*qɃ��wo��CV�[.w�:x�֤�Kx�s�hq9��G�z)��	��`�D¾�l��6��}BÕKޘ�(��	����V����wm)～�!�({M�����r��XR�%�4�*uF���j-�m�D^�HWP�]�C�g��u�:�=+Y0?JHi�,�сͯ@kʳ�#��p�Q6�8���Th�a������Y��7V7��>���^JI��Y#ATg���uG�2���_�e�,�~�}h�+�;/���χ�]yD�K:�\c�=������zO�J���S��Ӫ��X�I���|�Нh�x-�B�Fz���g|o�?���v�\�U�kt+���Ήe�y�f�3��B��nhW%�̉`����ee^<�E���Fm�2��~
�p.��V��XzK=����Jv�2B�k��-�vJS��Ɨn��a��ӛv��W�hX�NryR��ۦ�5IcOw�/+�rǾ�V/j���0v+|��n�xM�o_�^Y�±���fe���{9�Sb�Lyj���>+�8�V}���vܷr�����J̌�1�l6_���zؓw�r9U��_Ovcۗ�A���N$3D�]R�#P�V��\x�0��׍U4�w��M�7��%�d�idD�%w�k��F��u4�xd�ړ�b��5|j���(�F����7�ٲ�h���6�O���P[G�H�c��MP���9�y-��m��݅��f�0fE���f��6(Κg��]tк��>J��]R��|/s�x��+:Æ5~�s���˸����&]Q*<P�7U\CUDs��c�|{��mm�C�u!$�6��2��Aw��G��r7�+������7H�Q�,�O�Oj_��ܹ^��403đ�'-�ɶ^�thx\�y��~�v:���.�h�wIyF7�l᝾���Gz�6L	J�6=A{x�Jt�&�Sҵ���w��~��i�3�ag�eك/h�nGt�1S�o_wX�e7Gm��J��,���g��cF_T���ĆV�3�u���&
KE>�v�Ь�
�͹�]i9YZ󙘄�TV������Ȭ�D&��5n9[�VQ+��
X��ޙy,ꋛ9]���L�}g���3�b��23gS���o�V���2��B���<�j��r����:Ϣ������~�#ُ���|p�<�!!Bt��5�����%(�A]j�`㆓���j�����} ���~�G �(���o��a���"��'��||w�HF��א��^'�z�.��2'K������2���E�����f�8Q�h̽�g��V��׉���,͓���\�/���U`����J���t�n޼���m�ٕ)u�C˼����ŧ�
�>u��⇽����[����pe�ǀ+ؼ 
��;�B�v%�{E�P����z�k�<\����/ �ʘ=���V���i���-3>�"=�j2*�S���.�>�X�w��]�2Q���Y�8K񔎊c�Y�����(u��� ֽ��n�Vh�Ӌ�kW�]���3�?P�M�>�ɪ���G�|�ڕ��UN�R��^�p�+�Զ��j����1l��,���Ա�����/./.24�ؖ3芭)��j����	�o>������-��짛���r��w�P�|3��=LF�{�H��8��a䁃�@�bط�`C�d�ڱ?���]-�c�yS�훎��ǜ��*.�n�r\m&Z���Yh��޿.ndZ�����֢<�f���Y����G�,@5v_7(.uÔ��C�N6=�&c<i�v�ѼεպF;ؤ�N+�v�F���;0$�����ގ�ӫ�i�9}1��9R���t:z��xp涧��&w{t���V�ꣂ\[���31ݗ���+s��T,���x�	�ν��WD��3�1^��a����+ʵ�Aa�z�:�t�R���\O��°O�G_��e�ى�@�����
����	�w���n�!�ܪ_]s���!�R����E8�kzu�3���W-z�fμ��2�W	P���(w>��eI��!t�rϒ��5�wg���Rַ�ن}܋7c����H��$��
��X��:��#HS��k�K^V��ꑿ/1�w=�:��E�UNh�%��uJK�T�0w�,���N�&%	R�3<�����6K�T����Cg2E
������j�pwEUI�\�:��=�l9��I�:Y7��x�6ѳ��j���wT��K~��*n,t}\|b�0�����਋CݟP�r4���*n�sp>��$�k�</��	y��Z��^Kr�� �c�&)!g�{9�,�m�V�췑�v�A>[��n��3T��U^����1v�I�46�$]�Ҕys�2`��gL���f_���o��f�1��VS��Z���u���T~ū)��T�C��с6u��� fT9ܳ ����_ӧ%�ĦE�.ʨ9_!e0{��|^��|t�U���:8�q������1P�i�^��v1�o����"�\ֻܸ+K��u���C�:�W#f�D�$o1e>��c�w�W^�4�C($����BZ���,�v�s�E��f�j���z���l�[��W]#��i6�����m��ʯ�W���t0we��C�⧹t�f�%gZ��fos8!�t�a�%�9�B��S��j6i��|���붛�9�䞞v9(YG=��F����uz�8���/���c$^�M,�ބm �h��S}ҳ]vkqQ*��t��z {�مG�'��;��>�ݒ�c7����1���f�½��T��qNQ��t��pp{��ħXU�E�]]b.k�Z�]�l��,���#���7�"�/I��,�y.)��ض,�0}H�vIYiX����[��v�q�e��v%vǋ� �,��;��0��u ��Z�A����#X�{$�m����ڻ��o��%��x���2ou�Aos\n;���A)�C�S�X���+��Rg�rK>�E�M�bA[�tFR@�ԛ$�s���JMlIA3�N��߯�kXB#U̗֊�`��
ybYRi�w��;���
��Y;}�r���Δ7;�|�ӳE����3�L	ZhI1g��7���Ð]h}���k$=��|�Г;ژ�s������.mg	�T��Uj1�i�d�ۣo��:N�kV/`~��S��Q�0�* P
�����0��q�����}����u�{NZ �z��c�AXƊ�.!�ns8ə�Ŗ#Z(�]�ƷP�w� ����wiHj[�f���jq�������q��q�<c�^�Ԫ���г2�8��J8���r�]�ne�;"��&Q���Î��;5�ÄrU�z�]��#����,s#�pM^���l�f�O&�1�GɊ2-F}�G���8���4枚{ex{�:0��7FA)�>9��ˣ���hP\�j�a�u.0�ٮ�a�̽��/�Ty�69[�Z��ζ��A7%�k�J�lN��o��@�8Wn��K�֬7o�s�^w/��}&�.B�[�[���ݾ�(�1����*Uw��e���̾v�T[j��υL�M�*�\n�B3Y�t*�5��wdB1zmM�?1�)���|�q1�wkWI�� �{��d;z���i�M�-�����P
�n����V,X���7��2�ũ2+P�F�,u]���g����b��"j�""#0Ȉ����b�22R��
"��J����)*,���&�����"�J*�b����
�"f���*���"��X��

J�$�B���i��(�&��������ZZZJj$��	�̪j���f ""`����*�*)h"����(����hjd*��Zb����"���")�&f(�(�)("(��* �Zj"�H���	����,�H���"*"H�\"���i�"��R�)*!"ja�
j)�(����&����(�*�
�
$�(��!��!�fii(���
b�%����
jb��"Y�(�"���*�f)�Ƃi"���((�����߭}��կu�Ŷ%-�f��><�S���U�F���z鎥����.�^Y���3UBwV	΀�;^�Iq����<�GfR}�"Ww_��©�M�^�5�	�&�qC):v�J��æ������;W)���x�՜3�Q���7kѬ+ob'ف1�+�y�p��k�׼����ᖓ��\�A�wS3>iL�|\����(Fܼ8tO�C:���K|f��%D�B!��ӝd�S�3t ��C�v<�p�'.��\Ok�S0�xA��h�_��fx���j�s��s��Y~��=1%�������%}�d�k>{u)'X�\Ok�G^��Z�+���6�[�2{�n�ɠω�wL�Z��H��?x�>�VW�5��}�z��-%ORmɤj����A��m)��wHuV<K�[*Q�/U�L���§�#��G���zL3=dYk�Uy{����MR�tu�,���R�j��z�ʆݼ�ީ;�s�������|����9�1�OE=Y�<�̞D¦'�Q'_u^�oPc���<=2T}���ݯx�v��K�E��}
�a�,���.U��2��t�:f��r�r�8OoO�uZĊ��`�ې���$|wt��ZN��G��K/�oF�c��SC^S�p䏰���=g����7:3�6�M�f� ����Ht����L�g+K�
�b�r���Ϭu�iC8M.�����B%���c����(V���P��{�6��gj�MM����t������Z�Y�a���,���X;�#u��u�2i�-�MH��>�i�%���u�Jȍ<6]Ax$�iW�M�S�;���I0l=��,-��[��߱�D������.��߸�n{%��k�	u��x�R{E���k�=;��~��P
��D�ŲJ�d���0vx��-�B�סx���ơ�5�f���I��^=ә�����֠4W�yG ���VtD����C����%�l�W*Ǻ��L.��������]��cHi�r�)����J���8�9-:�������[�b:gϸ�wZG�wv��C@w �����	�Z�g%���+��=�.T�5uo�ڸ�n��N�U�䏼�lt/�B�oF�w���+�IG|�Iϯm��5	�QM�oL8+��H��U�<�=u�PM͕�#Э��F����s躂{K�Q�<��U�j�zow�⋶�ju���=^Ltunm���ꊡ�������e:�ucf|���e�K���:�=����2��=�����q�*Ř�xa�N��%�F��~��v���v:WҤ����׹|k]�Cr}�]�jϦϊ��|%����7A�vM����
\��ܝ.4:C�s���z�o(�t��G@���+��f���g&=��הZ�CL8)��>7dˣμ�Q��A�:+�"���Ո�u$Y�{u7��Y��M�M�7N���f���1W�-���銏�FɾwR��zsފ�Ў#�nǕ{|Y�(ij��r�׾�Ξ����X��2k�|c�N�<�Y}��{�7O��!����Q�p��HH�Ao��sS�=����ܼ���z�PFo��þ�W��K�����J�I�b.�@��.����� �<�P%�����GN,P����Af�8({�;�o;p��uW����,D*���U+w�,	C�v�u}���y���4�8��lj︾���,�xYy�i�8��r��P�dB��lE��Ԯ�V�JJ�-z:=����}P7|Fgt�U棫=)����Y>c�F�<J��6���NŲd�G�j����X�U ܶP��zV���(gtC���p!K�9�����0�+sT8h����ǩ�3��`�0�XmB3�0~G=z�'��Tf�=V�����߼�:�J�[T̤JJ��3�~�B�Q]�/�K4���`K;P\4��%uA_L�|�n�)�y�=�(:�j�,��J��59_7[��C5����Hq��hԚW�n�]}G��1�NT�2�S��C[t�Wcrv��ΰy��,}��.�S�u!.m�>�\�|�>8D�T/]�
���ɞ�=mpb��6����X��͊��Pl����u�ۤ
��x����c��p)�%x�����*��������8\�0i����繝���i��ks�#A��}{�T=��➛R�]j��C�PF�z{�,�fzft���s�V����fS���c���|������m�����-�Ħu��w����3�e��j����f�9x��5�hU{+�p�B�8\/+&���>�}�ᾝ�CD��IxzSHV�M���'#�>�g*W3v���.+j�-ڭ����|Pq�^�*]�.U��iN���soD�Y_d�)"����Y���k�_�r��/�%��ck��'���ų[��di��[�9ʪr��a�pw-�3������3�zy<�8n�/���}�<�]v�z+D���c��yI�O{�i2 z�5�Wy]�SR�Ve{M)p�D�K"�#]Wۧ+�i91�*>�i�2�=´�Vع�҄�e⽝[R�e��M�]X����9��:��K�������P�)����k����|E�;�@��˺���G'��+{��V���wvG�'�k緖� t���[ʚ@}²�RF�p�KF ��6�c{���;�.�}�rb��*�'�I��^J�RO��G���bF�腍�5�S^ܥ�d��{��ީu�ܯ�#�m�yT���ꐒ���1���.�9d���'����Ǥ^��=n��_^�z�������.������cUC�.���\�>S�m��;m�x�}��x_=1l&��u�gҵxi�yT�I��-�����KW해N�(x�����u��v����;�Ǹ6'�ͯ3���>�����&{����F�)�a�}���z����Og��#�q��Cv�#�p�P�4����^綘{t�g=<���0�PDE▂8�T-L�iL�)�zK�y��|rxߊ�E��U��q�s/\j.�PqZ��fu���� ��Y��~��r���.��V��nu\����5u���;�v%��-���{G��j�؏�2u�����	�3��x_^�BO����T0�&����V��͎���MlK<&�RqH�/(W|��:���ǎ�[wI>8S��T��q���&�K��z�0�gm_�:����@�c��'�],s'k��F��y�5{����]h",�oo��������$��U�؎dܓ�]��n���H���l+lB��9*Xc�������{�ezr��w�#�Ci|	�X���G���t\S'�fH��՛��3u�^�3u�6�
yoR>��<��KR.���,���R�{�P���W���Kv{�j������/�{-!9��G�z)��O&s'�0�0�7�蓜ƛ�
[���w�XǣN�b3�:�w��i��RXבz���=�×2�<2d8pLhŽ-1e�ݯ6 �;Vj��>	:Pu�nJ���Z�Y��3Ҳ,��$4�rʭ���v�{g>N�[x��q�$��Ｋ:���%tF�PZ��4�����u{�]R��P�mVu����.�ٌ�n;�
���#e�Ѻ��<6���^Z/.�k�(�)g]D=�WNy﬜��H��F/�����MO�q��A�l��Y9��xK�����nc��7��X�����^�æ�;4=U""�z卭jE8�2��t�F�/!a���b`�׾��S��M�����l_�ny ��r�*�l�����e��b����0މ(Ky�����BԱ�x��$к[W�N�1������z����o\��Ƴq�=�~����:�{u�F}/�OU�3�e1Km�pb��l�2+,`�nu��q�o��,Z���R�9N����b�®��R�����{����k�N&n���n���|.)^:�
�����á����Jd�����U���ϰ̾��|ܼ�0U�f�[)+�^X����5�p^�3����CȈ���N�L"������@p��w�m�J^z�.����/��ċt}'�_172N���ܡ��à�5uFk�Ne�Ԯ���i��#�������e�y�̞g����w؋���^��N�2zƘK���i�� �ty��V���U�:�_# ��U�������ȇ�~�[˪��f�vQ�	�x����H-��*#d؉{��~]�;�����6G�E�F�h�GQ�k};�X�ӿWF��s���&)B�b]����8/�tq�ۖo<_>#��M_��.�'Q�A|=�|�]9�➕���u��y��0C���c�Ȍ�>�ϊ랜s�h#w�X�Xi�lwE�S�Zԡ�ځ/:��-�u��"_C����s���y@n����P��x��X�o���X���^��w�nmv�F�е.��~Ƨ�V���	ܒ[Ɖ���5W�{�l����'�xߵx��Gh�}�^.%�>�(]Ca���r��ѯ-�}��)��:~'%m���ԗ�c�f�v�r+V��[z0p�w�2zm�p~t9�~%$*��/<;�Ε4NwJ�a�vb��v9��~����K��V�৴{�Pò��|�}��ԅ���Ӎv���7�fIsq�����P9�DԞ4�>uf,p[ڬ��'Wԍ�x�A˞��"+�ׅ�ޅ�2���l�tu��c��y��/�xq:�@��.
�n�i����5\���^���{u���=��a{H��U���[>��y�r�>��>�e��*����ǭ*Z�jdL��g c:Ml6=�dǢe�F�>v���\:���{�,V=��M[�s��}qt:���v�X����;��p�����#E+<*�o�/鴘�	���c�ƽ��ټ�f����/({ jfGa���}{�T=Ytp��Ԭ��AS�Ժq�u6s����9=R*ʺ��Z��P��b�����;�x��yx��Q�i�eB���ђw��]˛х���r"�P:�C	�5P�slԯNr�`��dd�C:�ۮ��;��$Lw�zj�g>���tx�6CGq�.���ػ�Ѻup�8'#�ޖX�\���˞�7�yP�d�毵�g���oݱX̬B����f̞s|���;��i�+��'OVۺ)[ytB^�������
��$�-�o���ͭ���k���r"��ݛ�G@"�]a�6-
rh�/�,Z0p{t��=�%�`��nm�ca���(1�O�6�4�iW]���m�f,i�[A���nz�T,�u��{���2sgÝ��&�V�Y���R��J�������w_������obJ�[�ا���̧ڶ��n�������U�h4(P#](O�<�Z	�KW��e}�|ϸ�l�y�թUq����ϺD5�^g�QV��[F��謖E�C]�˙�s��L���)�u1��9�J$R�oW�9�n��,*��ROO�p�bBbF��Z�{��p}����>�#2���5x�(f�ἪVoD.����&c�.�6gcy_������K-]��Ue8:�lQ��B��nx���j�pwEUO����4�:��Ř�ζ�h@�w����;=Z���u�g�@�k><�\���Io�xeV�l���2[�����%�{�3v��em>��nƩ�Yݻ�]2A6etkB����o ̞�w��|����ʃ�<-0�Vp��q������ͽ�`��1�+�����Z4^d���r�]g�W����%�������Gde���Q(�3�����Z�0֣Y>r$M0levY�J���6�ʺZ�}����@۪6�nq��ɦg}�]<a�����gd�<��f<���|�]��q����]�'Hv��
��D�w��>�jfg�)������zE�(�|rx߈�qCEi�\����֦�1�N#���a3����U¼;f~����r���ӂR��.�P_N�i���~�ս�GKE2��靟%��$��?0�^ 9��ev#�@�� �p�U.8��9���{g���]�?%xk!2�+J�?��\�N�Eu<Q"�ڒ���,OW��5�L�Տgi<ޞF�wod���n�Q�<%�F�N�� �b+GF��V���U�G�d}J��[8����nUr�g�Xj�ˣ��@��0I�S�/^q@�[�L�����媙�.z�_�:�KC�_9���z)��O&re�̥T���z�	�Ve���y��6j�
�����W��N�L�%�x"��!C�NTU��21L3��5*]��Y��m8=����'���V��WY~G]g*u�:�=+"Ɂ�RCOe�ΝU�g���:�i�~����{�h��#O	��-I����fG�����<����Ú��K|�����7�[Ɖ�Ã11����$<�7��DuZq�,��+����͎�ehBc�ymb���ݒ�hTv?dn��iM����9ʸ5ir�|������,`��T4!G�[5=�y=9�r��:>�T�Z�J���vc΃ltҞ���OQr�R�h�.���K�R�V���C]�k ��PU�Ȇ�+�\6-7���F��Tַ���d�*�^.2��oq#zg�&ˆ5T��Ϊaw|o��t4�qu�,�j˫]�����6�.|(���;�X`��H�DI�ڋ!�Z;��lR#�\��ӝl��I�Gt�Om=�S�ruW����i�r64b�t�	I%a<��'9��wݤf�ܗ-#�h��g?��3�p�5��}4:{b�1yi��I��vZy#�I)m���ԣͧ�CF���R���X������6 ��FsFT�k��dm��Kd�������Ք��Z���w��ʻ@k��uk�H���a>p<�So�uNȘ�z��N$ŋ�64��֭qt&=)�)Vm�΅RLtbK`�}�t5��F���:��"���n'�����$1pG�w*��L���_c�d����jj��q._5E�Ju�+e��vm��}q��R!��}���dS�4�<wٹ;J{���W�\|,��%Xmf6 �hgmH��C��2Q{%�a��9�IZɫ�}�}9}w�������ݺB��:�Y��ױ�p}x��˹I����9.�㛳�}D��Q�Ɨ����52�xz4���feƳF_c���4&�M�NA*�GN�V�#�)ee�h���_l4����j_.XN�	�a�S{��۩Y8��e�w���FY��Y��Ơ�ގM�=�[74���6Vx��I��������c�yԻ��@�}��<�5s�Vo�ٚҎKG)'�o]�� �[������yK�u�ҭ��������Z�/��M���
���l�w5p��+�P56�o�Z�Lȥ:瑒2�P�8�t��Cˁ�[�1�7�՝�����q&��-�ʽJRw�V�5�/��[s�L�x�n{��7M�kYDon�"�a��V��iC�i?C�ґ	�7h�kA�l�'������Ww�>j˂86��-�����բ^���U3�~�^-��`k'��k� �/�{���n/��.�����p�ޝ)=���m'i/���Z�F��2���[�j��b��$Wm�u��A��n<-;4bo.�.-�z�L}�B�oX�F�i!YU�p��Akg����z�p����兓�$ǐ�\K�r-k=ܻ���[G#�?g��]�6⾈ƠI�B�ӻ��w
90�Z�`���4ɦORcaYkh��
mY������O� B�A!LT�TMET���b(��)����h�)���*��(�"**���()���&"��"��2��*������J����J����&"h(!���(�&h��"�*��i��"j�������"�f�i��ɒ2�g2�¨22"Jj����"�l1"*��
��
���3&I�0��i���*�0���
��"�h���2Ȫ�#)�&(�,���r2������j��*�2�"*��("*""��ɨ"h���"�*����̈����ʦ�*�)����"�(�f��*,��*��b�"
�,̢�,��"��J�����r)�h������ ���$�*�������*&�p�$���h����*���*"��b��bH�3"$���J*�����+� �I$@�~	�G���;���qI���=�����B	�����BILWj�F�%���&����͹F�M�K��%�IF���X���9�9�vH�W�]z�x�y�yUS.��������n�H]�ø��Չ��=���&�&������ʍk���f:%�L��,�/��B`�*��/}SC�<�h.Ku�����A^/�G�3������ʌ3)�WK$h����-/�i�����}���z����Y�3ڐ��/����P�Y*⇜N���=�.<TBgfc�:���m�e�t=[����[�JK�痃����1���o�C'.�dR�=,��<���F=0����p��=Q=�7Jա���%c��\����/x�W�G�b��Y7����͜����v���J��iOD7�ʽH�"�!u�S..4��;(w���]�)�H�"K�rR���n�B�`��M�;�ꊡ�������e�N������DVj?{���Ɏ�lͭ=U�)���vQ�O!��������=�D��@V����ev��������z�
|*��IrB`�Vmafo�eg���L��_���1��ySFW聅!�+p[5�v�@�{,�4�ˁ�����]ܶ�7���x]�+=��|}��,�	�{��DR�+X��ݮ��hB�ۮ���Iv�K����f��H�ۢ�7]���;���q����}�Y�il�v�v�WU��7E{�y��0U�-qׯ�*ׯK|��&s��qeP��{�Ȇzy����^���}s��LR�%�4�>1u���0>�+��S��p�H��'�:���C����.���E���8���fJ�7J����9����Z�#>N�V0Xh���wE�/��-g�Cݶ	{�O��ڻYY�rgk�MyVmNX�~��=�*�pL�B�.����5��k��9T߆�3i��%��V}��t����eA܋�`f�*��^J����o��a�˲!A�6"�qf/oS<<�Ӭ3�Wڣ����>��y�]B�X'�*�C�b����g�:l�g�vq�ֶ��6���IWע�Բ��?nu���I/�������U`��x����Qk�j�����q�/_� �bx|�
�}��9֓�����G���]O�z�����L��/�)/OL���P@+�+l������C����cҮ>���{�%����{���y�o�O�H�g�ܣ4/#��踷���-;ZJ����.�7}��81o�oA@��d�a�JX�y��ySr]�j��8w.r�˷��h��]\����W��x��@��Jw�(�O:�q�b���Ol`����&Ԝ��i��oj�t��*#^�^�;�w5���S�K"V�{�����U�bQ�Tj�۫������$scA��}{�MP��ʏ���/BkQ	;���\��&�������=��u����������M��^\^�G�X�[�p({ԯͶ���\q>��]X�!lX�\�U!�T0��5+��)V\�20N�3��/��M��s�cx��=��9/�Ն�^Ј��tw��%��搭k_p0p�>�~�<6�����TMA��@�~����l�V���!��wu��]tXF��Y��f,i��~��;��ݖ^\��tk�3�S>j����
�^[8"_��)D�b%@�����^}bً-�H��w�e`�%��wc����f�,=.-<�:���zfq�	��7@���x����®�����j�w�e� �rڨ|�۠�H��Ia�.�WJ�m�E��,��$�u6�͗��zr.�,���n�A���?`�O��"��K�A�JI�{���%�t�G`r���%��f�_"ʯT)B�g�#�w�Οf�ἪVoD.����&gU�3�u&N\r��HJ�ؘ;xR:J��㯞�k�����Dv�q�0�ׇ�vI(�z�CS�� �z�#�����>��T���������N��l���*��e	w��*2�r}=�ќ8�:�ϕ�Q:�:�`��2�b�.]&e-�:T�].ۺ�>�:Sġϟ��S����eC���$�W�e=�R{@+�a��[�t8;2ۗ�s��xPwxA^m[:N}�CK��߄�FϦ�/?�*�*�+|�]	�N`ܬzW��4�gAw,ۃ\�i}�$)1=5n֭��^��X��ڗ�K4A�y��I�څ���Yj�8b����G�ar�0S������E���_{��59n���m�u�0��K;S�Z]�8��G�VM�+�xv�8��;����r��zE릷ڭ^��d�7d�v�"[�=1{`�{����Ic;).K��T�Ү���Jƾr��d>��.+t%�^�z���x�O-�CH���\Wmҩ���Z<����� sP���|e�^���4���l���?\��N��Pp|k���d��R��J����c�R�����o�Z��u�X<����ĺ�zf�5ޙ;^D9���K��Q��;� W�P��K�:�E�ea�؜븞�o�b{�!徺^�.W�k����=,5HL�:�J���b�Ӿ�&�}5�f��Uz��;DC���]���`�y>\�/q�w@�Nz���g�7d��
��f�%S՚ρ�(�yr�vR���P��E�����C:�cգ�٧^�ղ�<���P�6�ho�,��������}�S�����c��T�[jmz_�:�X�89���OE=Y2�\�&_W��}˹=���^�w	b��.��r]
�<Խ��N�L�%�y�x>�i��R�_�lQoc�F�DU��}��C��)x?�itE��G�[����������t������5��čj�O=�������W3H���	���異JfR��I��ab�}~�x�R*���v��ݽ�r��j�7Q0V�t�y�pЫ���6_���l���������x�u�#��xj�!��k���r�\�+��U -s	��tN�-�zQ9��Ж;<p���ɔ�n��%D����|)��U��5c���C%{r��<�4�����yG>3)�V�����l�W�ɉ�=����V�Y��k3ָ���[E2k�3����i���Z��w��4���BH�ݙ�J\��s}�ͻ���Xt���M��I߮)^��]�[�� ao�B\���T�.w=�#�\��n�g2��OJ�:&o���Ha���䲥�;�Hh�¤��k�$��P��6��N5;�S�eqbOI�h_(=G:����،�/���k�ӂ�]ƺ��.�69."/eˎ�vp跮-B��sB�xM�l<D;�c'gQr��iͳ��R�{8$�����!���w$���73�;�v0���]�a54��F�&���.�uU�?�V#��)��d͖;�?u�|�x���YL��Z��)V=���7�75as&���C�N�1�&�����s�U�֪�`�y�.��%s5��݁.J�)�T���f�vQ��4��S��^���&]_D���̾�=�����)��i��I�6U��i�i�pXY��'eT�<������tсx-h!�l�����mo��,�3捓�U(��\aB�-}]t����6���C��;�
>կǛ3[Z����}�W��ax>h�[���I3e�dZޤe�[\P�a{m[����������k#wmmA=s(#�K�X&<T�wE�!�����{{P%�2ew�ҩZ�V���a.�-��v���JI��b�*�h�,E��UCY��.Z<͚oh��ܨn���&�����^�6"�X�~U/讥;�y����
�_K�!O	�*vQ�;'���?=�rJN}�!�wg�o5
����*��yY�H�S���`�ЖpQE|��b��J-��Yg1�nq������X�& ��j��f \�P-^��]��=�]d������ǂݷ�`�]w��v�++��`}��bG���_v�A�Um(*����L���Q�݉���/��\�T���\fsg���{��;�t�e��u�1��ּC�d��/������/��;!d�� ��m��>����6]�Yw]���z�Di�v@0cţo���L-m&O�Ό�G���]w�e?S��ӷ�;����o�0�!�n���ǋ��k��%�.V=mpϡ����EoL̹T�rJ��]�{����\��H�ϼ�f������mI�W��kj����dz�w�bʜ�U���d�٫��Z<z�����33�a��h=��b��FMP��ʏ��W+�P�~��j�����qvU�C	(Z�ނ�ge��̧s�w��7������WM���m!l6�ζ��ʆ�^]���C�@�{���}�T0��5(9�WS��վՋՇh;:���ې�A�&���#�?���I-�4�i��ӫ�i����^h>L=V�_^;ٱ��ﲡ�%fl2��U����,/�qr��3Ƒt�<�{���Ok:"|���n=���'�z�u��N*�}峆Y�<5B)�[\L�N��˙pA��^I�z��]�!.o�ޡL�^-)f���͖_bc�l�7+��5�j�C����Vy�b����
޶kp�ćN c���gºE2�s'fwb�.Tn 7Θ�z�9�{����P�������˳r }Vi�q��*vn�9̡��q�y��Nϰ�����xx̉i���~v"�^x 79�TF@6�������Q�Z�ByJ�s�+t0t�k����eq�
�8��pLD����os�)���}ZI�H�����]�T��]:�&(	/%�)'���xk�-}����y�y�tG{ѱ�e�B�p������m��>ͼ/�ʥfoLT��E:S^��1�kϑO3�(=�Y5~��_	Y"'J��/*���:�C6s:(P�����r�*7�'W{�X���l��2L������z�zY�Cq(p�T��O��t��/N��^�W��M��-���ޭ3�t}\|b�0�C�BHBC��*�d�l����!<�7\���V%��mע�=�A=KhC�]+���oՓ���V~]�"�R��l{��"�Β�y��{L��91v$yU?R���b��&;*�jfcJex�S�鿲OJ��{�Tߵ�|�����g&����
ë��ؖ3�/%�R��k�l'������7�Y#Z��t�VT�on�s�m�®i�\i#P��gY�Iھf]c���btrOo1�~��^ɇ�sm�X����EN�+3X�7҄ыP�F褯^_�ޮbf��JU�V(���||{v��x�r��z���L�9q�Le�#����g^5���G�_��v�����J<M�ǾIh�~`'�� u5�u\F��ٵRe�7�X���[S����zz:C8��̇��|N!<U=Eu5�o��)�����j�,��S�!�nj5<&N�W�f���]�ĺC��ڿ��u^��=���y����&���鯏E|�N[�m{�P�xNTm��ayÏ�a�S.���:�?#>s;�$�ڼ�DxU2�>�c�b�P嶦ץ�C�~���s�����SՓ-��hVm�i���}�MJ;�|`�6O�Q'�/��s���']�g��ƸW���=�{w]ro�/�T���v�A�ßLF��.�Rl��D3���8�}�GfW\��Cד.����'�͸���5�&23��mW���{�J��I]����.��\32JƉ�~Ǚx�M.��i׌{��r�x%$��,�����l��7]>�d���-yh�z]�9��kʹ����:t����_1�I.�y�MAL�D��J����И9hB�}��}���k�)5{�(p%~Ș�s��֋�`^K��CNV!������Xv=��&���� �Hh�3[H�О��:�ݶ��]N�t�e�{�gki����@�ol��uP�E��VN�X�O�<-��r=�nd<�ފI+J�մ�זJ��R�n_����x�֠4W�q�~#��w]�n3�9̏�u&�>sby����i��&Ւ��n`g�qu�����
��9�OG�t�s���V�l)�f܁ڷ~���X�̌]i:�+�<�+��Z���`��j�I��-����f���>k��q��t��x�mт�*�6Z�IX�2�,��ap�(�5f��7�no��\��OQd�����j,�:�mx�%v׾�ك�Fl�Z)qh�>�/=ñc�f	h��y՞����S����؊PMM���~�/���VJ�����!^6��ޖN���n��ސv-���|��u�eB���N�1O!�������`׎���#�͜���\�dBٕ��	<GGJ�C��u]��f�t#�ׯzS�f�i�[��gb[�k�;K�b�
&��J �8��D?.���m��l�/��]��w=����_v�l��������-����f{}�th�cG�-�L���5�TA_��������( �Qt"�
��W� ����"�
��W��* ��DTA_삢
��Wb* �����* ��QȊ�+��TA_���
��W�TA_TA_�����)��-�΀BW/�9,����������0�-�� P�R��  ���H P����*P�

�T3%%"T!H�*��� U�*IQJE* (�,�UIIAU�@T��QU"�D��"EHT�$JTI�I�a$0 �B*�;�-���t:�T-���m����ͪ����j� ���J 9�:�q��l�Ff���M�-��J�k]m��R��-�E�5�j�ٖ0j�T�JB�ER*� ���(�8��   �   �3� : ( �  �5c@���L��J�m(��c5����D�"P� ;�r"�f��C�R���T1�UEXMR��\c
Y��J��҂����J��Ҡ�B�B�� ;��UThԀ6�m���#mUU-��ERŪ��lڕQ�2�Z���LA6��*�EJ�JR� ���JfjR����С�5m��`lj��E*5E%"����� �S�j*�ՁlLd���J��0l`
�H��`5J�**�R�p �
]5dJ�b��� �(���D I�4���@���E� n �3B�%L��	@�*�klkc ��
��B	�IT �
6
,�(Z`QPT3V̍��$��-5H���   ���JEPL� M  S�)JQ�6����M�)�I��h 4hd �J�)�`Cd�	��`F�D�� I�2�CP�2b��S�H$�H4�*(ѣ�A�`�&���@
5�MkJ�j""9�a$�T" ؃ �A��r��R���UB��ZY*tQD8�� @^�DTB��C�JB�*(��%�\��V~����,!�@H��^
"(��5�AQp�,�B@AUC'�ׇ
k���ߗgww� QC.(�P�\*U��7Q���U�V5;�٣B�M�����i)/.Z^���SI�Jq�.u��wC6�Z�+X��aw��ZZX��-v��W��6H׫RW�DP��!V&mж��G&�1fm\e��qk
��^�x6%�:u*GlL,�n�H��v��I� \�����$���6��˛j����)s)J�%^�҈Yf�D�U���훫���ܔ/,c �kc@�G�Ӈuk�Z���W�C�4��r�ݽ1��spc�e5�\1ݪ�k`һ����fbê�o�x�[��P��"�X���S2f��n�L�bY������b]�/S	ܺ�6)-�Ǥ E�O���6�f�<1��f���[]F)��>U`Te�S	,ZY.�A'p4�����:Q<�6��&֥V͍V�ʽ�K�L���r�m;��Ȍ�m�-����31ֶ�B�h�V��]>�O.��#�Y$]�[����Ku�5ZN���utԒųB�2�Aeܠ%m����Z��%�ݶtl�Fa$���U�qT����J��f�֛�4{�	�	T,��,x��])��or�E����Z5���t4�Xk7-��ຘ�cf��4������9ךE�ݍ���$ൊ-�oMj��f*<aG�hێc[w�QZ�.;*dJ��V]q�Z^3�I�.�sG8mm�w��C�X{�V�Ӫe*賃h�c�$ߍ^]�jDmL�m��F��nڭ���Q¤��jٕ�E�X�M���'�VE�k��W�kL����HRy�n�3e�[R%����̶��w��:�AQ�][���>ëK����J^ս�.��Q4��9&is�ඵS���{F��e�em�e����݊�����ljOVf�mY�0�i�7��7y�Τɧ����/Ku�5�zZ9N����w��!�nC{WZ-z�8^Qx��T�U'���T�'���t�Z�nd+2�[RL!�VI%���:�=�b�����+���I.�s�Q����e<��pԎG�5��[���
��bη�@
�[�
��#.��3�b��fR��9��\;{tm�N��Vƪ����j�ǹ	�U�a*���Z�u��&����0Xfd.م;b�Z�̶�L��[���S�4�˗qd[Ҋ�U�*D|ޱ�m�hm�0]�W,�f���!���2e��	�I����2���*��m0�Q���3sJöuA��YW�-�+���YA�0,���w��ޅ�]k��ʏ)ƚI�����1���u⫬kM u��S4c��m]XR-M�̰����p��
5�-m=���vgÐM2Klo�q2�v��kkhe�apm&�=IVn[j�,��Mez5�駋)L����X���K��8���v���@��N��t�YD�A�xs��Ϛzy�q�ln�K��vh�x�b]aն��ą�z�����%�N|p�6q��ҭ�V.�f�ۑb.ЬU�m�An �<:�U� �ɥ����&Z�,,�n�8%�I�x]�2��2��: ^��ԧg/NF2(-%�LYyyB7�`��f\T�)N��X;��z�2�=���]��L��B��β��mwP
c�w��b�0�Z[��I��Fi��0�K6���&5<7N�$���擮��
��I
����^<��ş�\�5n����.�3�x�Ņs��9��=�b�a��T��������$�5�:�N�Y���(l��v�l7�ub��S!f�z667����<` `Gr�W��5�>:�Y�n�=8�w�q��̭��*
��vQ7�#N�Z�ٵq��Ǖ�L&� a��ˍ֭��0��ş8�l��e8�5P���yd��T��Ch�2<�oU8ow��n�/>@�
�P[A��E^�2j�z��U��Z�A��k�AX��lm�+
u�5��ZdMH۔�.I�F��tT@�WL���ʳ#�[�(�B�"2݌ԩ�v !pG�[W�����eb��KH�Rw�N��耳h��tۣn@�d���6��L�YEi&�k���76�ʕ&��S^
{+n������ m���d��������"�[�QN�#�#�T�n��n��.^�3�BH����u]�*Ú�q�Q(s�A�]%M�]��ަ���n�q����X�ɳZ�� $�[�)����ƍ�d�uq"gV��*)��ʕr����B���GI)�*a�͔~�o.���f�"�a5��t������C2H+���]^�Hr�i��k���d�i�)4���n��죕���nM��d0^�mbx]��
�9��c��W�Є���!�D�ٲ�Պ���[՚#��#�Q��0�w(l�ڙWYe�
�F`Cq�FU�`��:۰�?`��y���a�mZ�i��Hѣ̳�Pd�9j]!�&,hlkwsfŅ᳘��Qb�*S-`��Y2�63p��6��w�b�!��2k%ad�M�t��ḷ4T�N`y��vj�J�0�S���n�6�8��f;jAy��VҷZ�M���|%��)'�x��kc
���f�0B١j{�Xj³�w�.�^nS��!�G
d\��J�m��;���a��k��\��b���\ʷ���X(����r���ەu���WEZWv�@�E�<�w�	���I.,k�}�V_:yt�*)��sVU���h�
�YSm"����G& �dB���l���२�dT��;-Y��;6���Yd���莮�[u�ݒ�� �ľ!�oF���X�,Ø���4�5�i�q`]��=�8�n�&��;XjZ4�Ťn�҇%P�+4k��38�M7sj�a��$-��Z <�EIleؠ�{��&5�mY�cb�,��p1�:z�W�i�`4�����{��M[����b�U����ۊ�p���lc�KN�rI>�s��{�:�iwAXcqw|pjtFR$�T���������	À�n��K��.TI�-칏c���Y���f�̬���zŝ��b2�2��jn��td�z�X�Ęp�*�ސ�"���	����7X���ن7H���(��QJ7Y�f$�\�W���^h�Ոؚ�4v��U!t�b�v��.��h��9�_7��^�J ��bәFl�<x��@���>X�B���������+7�B�l&s�n���{L���,0�+s~ɘ�E��w5�WA�c_#��������;��v�^��fn�h��8}�e�y�6ﱣ����Xe<�N���X�(�n� HZ���C���7��$Cna��A��+]RD�3[�
����8^퍣�I�)pŠ��#+( ��Z^�4?����taG��j�Z@��}g��*/Oo���c4��Ҧ5�,������^��.��÷��1��-��&K�[�::N&��B�֥��FY;�	�����
�W����i-�%CJ��V,x+�Jv͑BR: �0PQn�:� �k2���1�Yk��ҫ����K�xp���VfI�D��Y�W���wɖ)ޱ˂m;ç�N�$x�^TƔԄ��]\טkf�M ^XV�n�Hm��8�&�v���P���hԶ�˺���@ǺY��t4��.��2^��7m��*�$淘�慩���aBA�cP�]�i�mK��w�PH�����a|iX���N��k�.޻�ִU���Q"C��\FAtκn������u,Џ&�ͬ��[���4�v�[�u�%PX/c��cyg��n���jKUٲ�ҝn���3g��Q̱���*J�E�g3TT�ǚ����v�𴮩R�.��yd@p�KyL[�C&c�6R%J¶������gM��aJ[���cLU�Afn�H��k�Y���[���#W(�T�W���m6���EV`;�Ib��д&���䧘�6�Yt2��0�<Q;)��MET�ႝ�
�&-yI^;kf��:����3���m�s8��VoJp�G���̥��E��1J�A+H�[����Y�h.+Q�tCGRg/&6�V��m:��1m@v��^ؔX�l�T��T�VM��̨�����KXBfɁ��2�&��E�d�q�G4aw���[Y(]#�ܡ�$&��S�р�ٗK.������'q�h�c�]�2j�U�խ6�@B��VMm���lc�KN�ܶI�/D�c�HR�4C`cwBX8�j�}�c"����n���Ƃ�h�$m�{CHp)�+��}�G6�Fi���ū 9R�ʄ�Z�	����!]s�60H1��q�mk�I0ƔM��+Sd��y���|1�7$Ȇ�ID�.J��I�ܬ��n�j���[B�ˉNq�yr������x�Y��
�����e�Sg-�ɦ�EZ����/��֖JF9�:��,��8�DǙ�5��'����;��+qn�#ǈ�i?62^�`#Z)�|�A�W/xbGn������<�8��#��ڴ�,�3�Ca'��V�_,���%�|7��WJ%�1��5z��/3����N&�ʋp�B����k�XY��~�F��<��َ��pǻ�e�xJes���v�3W���܈6�c�e �s�G���7{���徆r!t�>��]������8]��� ����ΟI v����\����Q�暧jѸ�]�L����-�G���w�'X�����U�V�JP}ي��S!�7���nK�R�G0�QhK��u���W��:ʎ�	r��W8�Y-��ZKŔ;��Щ��<�T5[g�]&���N�a+%2{�L�^.�x�㒢�F`���wDv��|�-��{���F���0>�����h'�;��^��N��r��|��9;g[�&��ԥ�Bu�c=��<�3H�#GI5y�[
sy��7Wv X��S�2\�|&T��"LX�r��tn"qӝ��8-5�1H�s8�Z�����>�]Em��A*
*��ػ&���>	j6��kC�|�Vn�#��;I���*R�	���ΤL��m�fMʐ�OJ�G.�z�)��,u&;!����u-�ڂ� E��9L�\�<n�f̬�t���o��Ǜ2�n����WNA(��颰S�F�n��Ǧɺ�\M`].�[�9Xr��ޱ����b�I����|��`� &��	.61�P[�k�b���"������WJ����.�T�wS��=l��{��YTV%OX���k�|�8���.+���&�ab�&��\&�\��R�Ě����]��]Wiv"b�$���F^�2��ï��N��G_:��/Yuwr{O:�w�7w��2�Ր� iQ�{��	x�/���A��;yRzZ�{�"����,����R�vI.�U���y�s������Ԭ�ۀ�V&�p�qA��=����j����H(�����:u�����d����}�*	J[r�^q�qr\���.���c�R�(�%��Le9m=;(H�C;����¡�T���v�F���Œ~ݤ8wC̖�9�/���f�۵��n�c7iJ�\�r�t��J�W��1���*p	t�������KE��5{zy�Z�)�1.�DgH ��:��rК��'H�R#٦򹗧~H%.�S�n�C��;��N��M�
��餮��Y7��oֹ�s鶯wRvo�F�V�V�J��t�V/]�5g��ۈ�"�)l��K7(=�K��ȓ/��e�xТoL�k(B���nw���79@���@���U��q�<t<�����趖�n�RI�����ǚ����h��W1���j�]��#���[�k���<���X�ڻ����@��2��E*W���܍0r�v��0��ܠ�Z����GN�U�v����J��*�t D���r�b���j�JzVa�΂�Ųb:�N������Ev3\/$�m��:�tV'Qu�)���*U�(�s�0��R�9���xE;��h�i.6M���c�YC.]}�Z�o�#���PYPHM�-���־�m�kLΚww�W�M�	��j܈Ɩ$wpX�n��b=�+B�)����[Ղ���N������q�6n�X�*-��杏��� z"e^躵�����N��8�nw>���e���s {�xn�
�����j+�r�3�Ӊ��|�R����l���()3�����x��Y�^�W��R��4�Rn�%�
�"�9��A��¼�|�5)��Q�Of�K��*v
�C7�F
u-j��8���u���o��+�.&7YO.�YV� ãDfb����"�὚�S�GB]Ȧ�nS��i����"�����x�W��G,T��y�RW}qe�Jh�2m��M�m)}ςÆ}�.{\�N�ˊFM�%F��}���y������]1���3C�#�Mu���u��7��ԮR,JW�a�9z�;ۛ����vD����"n�c�TH���+��� �}u��3��X"[l�B��Z�x5��r����f�!󷺎�y�D�ak���*�ȯ�17�`��n�uӍ��F�q�}��-@�Ūi��P�kNI�Y��t�����K �]�js�����M�%w�4�Vq���
s8�y�-�:�j�`�Z�*�	����Fv��sl�x�	Q��YJ�S�K7+�^
t��/�,��5';]�ef�\Sz�Ky�����n+�6���KE��+,rGjJ&�'p_$�V�0u����=[8,��q�z����0L�X�5��6�N��2eCo4mV&�[v2n�v���綕\� 8fŵo_Vs�1�{�4��sQn�`���wJ�-{�ͅct`"o�zx��|��G~k%����|��j�aOK�DJ�С��b�q�(�k�uv�j�����c��Z=\�p-�B
y�q�S������*�epTSG�]�G6���Z�ڱ�@w@Ë8�|�X�Ț�-�#�v��k)n���2�^���<η0*!ݮ��$>��˔�v*�T��+!Υҷc���;�"��'w��	qG�c��x�R����;�ۦ�;�����}�	"�7��#>�ZZ�ghf�(��L�^����fE�Q�:L�( �f�#xOnU���[W�0D��N��=�jQ�����Q�ne�5�����e w[�:us5�Z� +v�uU�[�[���j�L���[�c��^�m�[k�+h��ﶆ,����X��˩�lxk�e�E�&"�yW��QM�n���iN�@��y� :�m�@�[)�rt�O��KP;H(�z/.����K�5}c�f�.l't:�w0���4�4 ��4�'wy��Z:C�\z��NN��s:��mjZ{��rf�+��ͩO�A]Ւ��9WA�,8WU��S�甦z��fb�"�)�7���V�ħ]�[1��2
������r�P5���s�U�c8��ݒ�%H��]٥\݂z���L�E�I,��1�Xz��� ��Wb�BH%"S,���,^�f@��@�ݠ���"�3F�V��N���Y�����yMVه.��V�JܲX9�U�H�=W��ho*����-����=�v��pR&q�	.���u��ҮQ=XWa�{�(ԭ�!
��Dλߓ��f�r�p3)��*��x#�w��. ���7}�1�� k<�S[��PZ�U�2���1kזY�tQ���{�(!�"���ձ^RO��̕��
V+]X�q�-�2�7�U��#�x��,�lI�[W���	e�W}���z�D$Fe�7܆_`R�-�f���Q��YE���l��p�ؒ[�����r�b
qQ�a�&�1��r�V�p�D{VV9�#�͚��9u`.�C��u����56їۖAĴ���ڤ���B\�ӳ�SD�9
&�a��;���ZZ�v���`�F��Z��w؊���pN�b���1�Ϯ�eN�eEr����SN��9eoD�hb�8ܧ;����f.	,` �TL�}X���'1�O6����dn�en����؆.�<��)q����*�`.�uZ,i�Ii��æ�Q��t�P�|�Z�h*9eH��4u�ax�[9v��k�:��Uӝܔ����s���L�
%�`�D�n�7 nD�18;�.�P�9��(��'�t[,�H�;}��Z��HK�w�["���I��T��1�S6��y���?)`\]�0�RI�x��u���pd.؍>�7�M�/C#u�ղv�6fP�pS�(���#�Dj�n���޽�$ܝ�#ssFrb�7s"�el�Z�
��&�L�	�W���F�½��W�A�Ɏ�y� T\[������a��|m�Y%v+{a�o8:��J�Ȟj	!�-P�%��ƶޖ��,� ٣� ���2lN���j1K7�^R��5M�\2q��35��cV�ӱC��㵦Nj�Θ��dwD晱�!W�H���o%��f)t%i��|j�~�u�c3�����k���i��[�_N� ]&�p`�qd����g:�|�*VH��nknjٗ�N'}��=�{h��V��3d����"k�&�8HR;�IIW�ȷ����A&��3:��\�7beIRI$�I$�I$�I3`2I �$�I$�I3�<�7��r��j٫i��vF{�EBjH^��ꀂ��3�����=rJG�K(�G����qm:��}�ܬ1�6����׵M���9S=g4�L�-ueթ�V;���g�����q}�(�r�],:��wg5m<�$�<y��;N��H>��lkl#���_+E�y;3Y�'+Z�[]Ԏu�Y����A���#[��V]ٲ�I���B��� ��TV%X`����5qs9��;9f�^��N�*o6k�Ƌv_V3(�u��ڬ����(e����5��F���
��C{$�h�2kv�eH�[�+�=��Z_X8�l�p�W�3Y]Zƫ�gגe�V)I�o��;@�X���um�<����K71����vH��f:����W��A��=#����;>!��إI�I�C����l��h8N���k��+�ݣ�>�������-���0���ȓ���45�rL����H��we�Y���]�}|W`@�|��u����k8*b��32}�u(uJΠ�����ÖG�Nu��zdn��jqF;�pV���'V�T.�.�K�J�⮋]n�#����
�/f�Ċף��-���0)nnN�wG�3yJq��R����%���$�Gz�W�7�H�u|���ֺWfז�rd�7@f�*��d�j]�{Rۄi�'r�q5��R�7/3���ͮ�n0�����rgP`���Y���ד:�Ă��/�/
����C�3$��QeB� ���Apt�7�Υ�/q�y���"�`�S�Fi�/h�|���;7a�1�h6���jͲ"��Www�k;q��ױ,]u5��Ϙ�:�d<�e�aWG9+�]�;Yu�%��%�8��wZ8��ʊ�;2n7���[X7��6�"��dS��T�:	����IPY�}��v�>�y/rH�yf���5V�)^l�V�˜ľ�T�@a��8c�D�e���P7�e��'E�=kL��b�}��!���^l�ŧ$Kvn��<yzR��wv�9����];�U�hh_���i��L�b)\�:�w���϶����� ��o ܗH&���Uy�R�ЇR��\�<v���b!�|k�A��ӕ���ڸo@ʻhL&��*��f�܍����b��Xu2'p�#;��y���S�&�Sv:�P)����žԆ��6�J�:��v48b��y,8{/���T���n��N,b��;��;�xwv�;|)�*�U�h�B��l�~41�gi��I�����m�Ć�dݻ�xY4��V����I�8҇7e��ٽŹ���e���=\-<ݢ)QВ���Y+V՜�ӣ�,����&�L��`H+8M�n[� ��9A���V��7k��Qw�'{lbH���뗭�ti̓q�0��9�g<�Q�Lm�$���*ż|VGa6�;��}�E}Q�t�L���R*���s8
Ĩbѐ-z������!�c�h�~T�\�l3��za��m��F%Jţ5�N�ً����j��^�-�Ƿh��$���yܢ�^��Π�-���! �\7n�,�*]�*�Q&<�24ou�������&�_I��,�iY�"
�\,3؂���G��h�F��n�����\E�U��M��)ѩ��8�^�SLD��JĠ� N�]cc����]1O����'g\��%+�8�fL>��Z��4d�ߌW��a������lea���|RF��.�Ţ�8�gN���,P�ɣld�.���=w��,���г!"bճ7��{x�գ��Yg��xq�bN��� �r�t �։�P}w��4�%^�s�I^���֩ĵ�7�u���e���V��:F\�����x�i���ۍ�)*d:��]�h[�.Bv�K��u󒲏+��$
"�fsO=�u����A���z�P���`V	�B#ضQ��4�4˂G�f�u�� �L�1�X�ق��{��Ⱥ2��aZ��T��,�<�Ѿ|/�W����[����g�&IAL�c�v���{v�i���u"��t�"��⅄���o:	��"F�������F�$�� ��Vof�)IJ�m,gU�J�P�\������rd��-s��I��u�z��+��{sD���:��aa��9 ������X��@�@���m�i�[o�93/mM��d���'n<�8�&o�9Fw'u���Q�\�rV!V���Yb���o`̶���KW��G+LN�t�,��j��C��	�]�	-5��2���2����X�E�8���+1�J �Z�㥢];�֩�	lK��u{�v��T����kwԬ\��ꔍ�a��S!7PTz�H��C)	�U&3;"#N����ܨ��߁�W��"���w�-����oĢ�hO���y]�x ۙ�>k*����ݤ*q+#�"���W��bVXU���|���gR�44�Fo��w�����u]s8F��r���RSz�U����Iaձ�^�y
pmJ�Ok-��-�'RZ>��D��'#�4�]F*wWdf\�e��P�L�:Z��-M���}�ݦWR�;��9SQ'1VЂ�����^��,N��
.��#���TP��i|��Ð�v�m%Xneɕ�6PҜ���)ǫ7o!���`��}��gQS5�X�^+�Y���A�%l��ľ˺������j`	�C�Ρ�R��
-���2l�ʷ�sVD6wx, fi��'�[+㮺���i�a��tj|�#+�����xrSL&���j�5�����r�y��G��΀,<��j޼�3F�(�y���o��V��wy���ւ���2�@���,P8�9>��Fu����t<2�M�h��e*��:����9�"�7��v��YfM-��` K̮M��Nowcp��MT6�a�/������ʺ�RTH��]��R�udZ��Kɷ���zc�I��]���qa�1%�i�,:9]���4����5EnM�kM/�Y�������q����6En�as�p��WJr������o/�E�>��uZcS4�sA��z�5���0�M]�/5Cr�e��zܺ���Kák�8�+�pK]|5(�쉁�'3�^Kdʾ7n�8
��FZ�v�U��֖�rS��a��c�8����Bi��(Y��𵮘0� e�<ڶ�hO��N�:�*W�VJ�6pu��Eh���hVh��62��WΠ�(��s���{��J�L�:���]ZZ�Z>���on��v��p�#'	[0�X�f�6넢 SjN�k���!j�oXF���%#�]7�1Wp��N]��؍j]�>��s�U.Rs	��dD;�r5����u���Ai/3��\b]NP$��u��@�����\PS�T�����XT�Խ`<�W��Ŭ:�+zgh3�x�)p7� �s߻1�x��*ޅq+�,uu��ǎ(��H�C��):��Ub�D��wNu^9֓�1���ؽf���k��o��yXHe)m\���X�:��8.� ϬitZ�أ5� rP��6��
k$r��R��N�;
Y��2�ҥ����0��2�S�R��v.���-9�iA�����e���Kͣ�v�71VȨ�{J^������{��S6�T�֍�v�Xt.T��뒓pS��SCF�#f� ��5ء�ԗH�*_m��;�^�N��C4�Hf���S���{���,�R�f��|��E���A*ki�iǹ��X��^mJ�(:��h��̺Ԃ��O�|��Xps�Ñ�~vU�ե�-�=<W��3e�[�ֹ�v�{��J��6�Ru:�DaY�^H����*���:�֡٘��)�s �<�-�����x��d�(�ڃ�cٕ��A��9iڐ�eb;1`�z�"W��޺aJp�{ԑJ������������ty�-)�R�ų&�SD�T�`Q[�9�incw��p(��n���P��Z-�pܭS>W�`�KLc�wt��e�P�g*η��-Kr譹4�[�ڲ��YҲ��V�j�-���vY�͝&��(�Ǆ�YQ�Qv�+��f�j�5w�N�)�>�蓫���ާee���ݔm�j��! tf��f���ޘa|Q�3.�S��pЎ57/���cT��ޗ�]���%8-_A)A-��^�K&Vo	\�H���o$��͔�]A�{Z��/x�J�7cwv���_�n��˭��;.<�J��Xtr��2o�g(�wat��iD0�]�3��aQ��v�{Ze
�͡Ws[#��a�U�Ą�,�[w����}u�tf�	�$!	"�_�� #�x��%ξ��	�?�j��_0u-���h��a�8C��PZ6�#�i&*Y��9�������۰)��ZX���O]gU��&U��y_Ъ�nΨ�á	C��3�בV��sv��A�0q�z3h8K�����q+M���\흦pI`�@�y�<�{z�Ⱗ,�����N���w(}��WS�jW�O�@�a(q۵��c{��5i��3�q��WГ�E�6]
R�/8��\]v�c��l��Q�.TsZv�yV�.�z:ʃAŕk*̣-n��q�h$7��x�P��U��s{+fu�=��/��A}}�r]�����S��%^wX3�o��
���O*�4�Sf$�⃭n�՝ty��<������z��\����ܭm(��kq�˔Φ��{�R���#u�qy�}R�ʳq9��B��z��l��
��T� �m(��EU"�X���j6�TX����\clPT`z�����|�����


E��C++U�b��YZň�*��5���P�!����E�aTP1*j��ʆ&�`�5T�լ�A`��a�S��5.�s0*`�EDFL-QH
DH�a+k
0X--PPY�l��`)-��c�a��(j��H��"%@��c��aZ�UD_�]5]["�4��(��R��AdD��E²(bL���J�V��r�ȬVbE*���u��Fء�
��忹����uo�o1������-vN��u[̹�[5t���rZ�����'2��������E\?���-�n��T�ufD-�������V�V��}@2�0t�,v���uۅ���]�B�mFC��E���绉�H\z�i0t����1�C*e��1>�����j��R<U��T�`�׻�V�]�ŉ<�X|c�!X[���JڻG����Qr6�B��Jk_�H�Ɋ�]������|bi���[�(}C`!�-L�O5�q3FbF�nٕT��:�p[:�Q[��n}�S1����S��Um�u�/�r���z��3z�N�PQ�U�-�N�1İ�j�Ag�|'�%{kG�r���4��¢���>U��&���R
���܁Ӄr���D��K��L�]r����a��SZ�)��8툭tx���e"m7��F���D�յ�0n��^���t(�͡k��x��-��0>A�4{'�'�
����:cD��=�]���-=}ϰ���z���y��f�Q�tv�y疢��Ff;�ytSJ[���zI�d4'�]OH�Bcx��CW܎�k����SH�I�&hI���2��ש��^Z�r����:G��hԵ�Z���h�-��Q=���m1�%�p6�_K=]yŷ`�o�H*,�Ua$��α.pٰ��py]-7�;����K��b\��bŒ���uo�G1$kl��z]on�N�*�BxK���hܫ��6����� �6PѪwQ�0�RI\i:#j���������^� ���� �J�&z7GN�4ڧ*�D�Z�l�淤��E|������y��9��x���=$�wı�NR�*N�Q>�6�p����{�u�=���tJ��ϖ<�RG#fKk�p��C��ɳ��=��_�pҶ�m��}o.$�h���1m��L��c2��Nz�>R��^-�^We�,V�6_:먻���Q�Y���CI���æВ駳�վ��)�ڍE@�׏lkla�	�d��I�mk���rp���Bhj�pV���ymǽ�y2�[�JVk�R16]��@��j��(�d�[\-���ͭ8t��q�]���#G�WfRXî8�-�W��<�яDح�Q���q������L	ޣJ��4��[nۉ��%Tfj��H���+g$h+vl��X�^@���Y�A{Ӭ��ĩP�)���H]��n}��랿o�C��aJwܯP��p�U�2�މu��c���5�:������������3.�w��=�V��4��'��iH~�u4h�-c�C3����K6Rvy�!��7����^=��8��ꕒf�vv�ӽ��5YB���_\�I�e%����ߝ1)��j�_aY��@^�PC\K7�G����7��K8q༎���bd	��y7b6�\F��i}݂��L�|ҥ�ae&���{�U��4ȦZ��fxG���`Y���5�^҅E�����}�_/��Xki�Y�mҨ�����X�K-���1���דѐ%f��9P`�ح�P�+ca��w��RUV�C�l���rFO�O�:��EuM�(4{57�蹈#�P4�Ǫ��=�3}������ߗ�yC`��߾���}��K)��O~o�ީ�Sn3O�Ll����k�5U��;��R�8w���G�"j
,r�	/}��x�߷�k�!�.��tڎr�pR��t�H٘2�k5x���)I�B�b3y.-c�U	�B(t���6"\m���YT)��6hl���Q�N�C&�hoK�/�GOV���χ�*���:Nf��X�E��ɘ'I�� �W9`����tZ��a��x���XZ�k�ed�*[}4��+o��3y��}P��B�.fw�^`5�Z4�ZV��Z��_HfDE�B��Y۩l�2O���O�}t�>Ѥ�����ypp�o�XDٕ1ꫂ�m���P�'�GH��~7F�qb����?�K����o���YCѪ�Z�\kF�p�`��|+h�*�_8���<���zn�=B���{q18���Z��-�ko$��bl�iҫ2H���!g����y�nʡ�[t�~';��RU�ө��ɆO@�)�;���]@j�:6����Jyyy�lDM�P�**dpS�2�tXrVOE@�21��7ͭ��f�L���"��d8��uѣ'�n�	fbf��^��2��M�����WǨ[���K^�G�t͐�`�	ʵ$z�(L�t�D�˅�����v�3��3w��E��*�'�=۠ǜ��k���h��B�ܭ�A�6Sձ���(:W�Zl!�s�׆	B���Bۥ���W@��4v�i�J��.:���*H���̸���Y�".�h�����F(j�eE<)x���yF�X��Y1N΢�����)E��g����sc�1	K�(�Y��ܒ� ��[,t�D��PQP�ՓP�P��з.h���&!���� 9謔5Xi,��:(+��G��lZ�ܾ�i�xz�שV ��� �p;fK�a3�ûݛ�Ĺ����Uuq���}�j�����6��u2V��osN�#!饓1����\�" ���L��kv'2�2Ӿ�=C��@�>F�V3Q��n�u�kg���,�j�q�^<�僖Q gL��{� 7b�����{����+�j����Rۣ��a=�&^X����Kuj�+e#1#�_��7�� 84����#�/�2�u�����\�)�6Kԝz����FCr�L30��#[A���b���Zj��+%�zv��d��'y�Pq��$7=�}�Im
UЊiY�S���=5��gE&W���\�֊�v��Ы�@�È�䮼�
���N�0��1��E��~˿1c���������:1��ڏ��`u�Κ;g��k��1[.n{y�^p8)�S
z���
9�62�������'�;����q]KuaeY�󍈁Q�E�Q}/ j��{8��A�^���Q�\��� �\�Z��:*�j��:���eֈb�oM�Qnr=0�u	�B8@1�MzzE�ф�q�uC�U�[����i&�m;��߹>Zy��WpW�Z�W[@�^��̆��~�����fN7�Ä<�[��(�K{c�c��>��-8�aނ��.#�u��o��Uz��V�ΐ���gJR���w��by/=�W +�x�n�`��1��ÍɸCg�O����ë�gv]�(�PW�Q� Dח.m�V>�'��Ֆ8Up}z�F���t����a#�o7�Ɛ�������/X�y��j���Y�R7$�׸O�G��jz�õ�u|x�Ɠ�>~�ءr7���xp`���v�F�����lP�&��{��o�1��J�i�-v�/�ޡp�5�<�?���m�>F�av�eq��g��صd�f�m�[D���;,F̆�Ǹ[�_&���O���(�_՟o��)�d���}��O�8���#��P�I˞+��u?H�1���e�z��=*�El�]�� �s�;�Olޕ��E<`������e�� z�V��y]&M/N<օ;d��q1����:���y/x��?���v�R�2c��ÑS#"��Σ�y��~d��bͫv.�����-k�J@�dN	@uF�#eu]T�\�Y
^O������*-c�T��"�GW�t	)�c�M���5P�S�DH����z�a�f�C����K.Vn���z݊T>��\NG��u����ʣ,�um����7���ꪺX
ѫ�atT�˃�^�>~w���S 0�a�6��3;�$)��yDݫ�j�c)�=\�'c`!e�wV�U�^N�8Q.�b���@p��jA���qI��5�v�A\%��x�U��
�ֆ(8�eOl�`b�-���,רČ�"k�l Ts�ݟ6��gI�{�#�������O[S�~v*h�4;�8n���4��#�f�yP-�.�f�h��0���;K��{���o�u�Α=Z-�^���5�
Wyٚ3S�}s.km�6޸B��ޗ�E#K9��Aݡsb�/�q�˩C�Cw�Q�]w>b+����f�sh1���s�CS�;t��;��%\xf4�r�2(�D��.��r԰�G2��;p[R`8��ݒ�I�91��Ý�:˩�����oV0���m�?�q���sɓz3uCYz�`Ğ-�9Cy�t�R���κ��t�CgXz)Ł��g!���.������Vc@nU�%�+oc��7�/�����x4:V�~{��q
��m�H�T�+���jV�x,	��7��Ӿ�{Q��WCL�[��-6���0�� �YM	ՀJ׊�:)9����B�r�N��u�$����f�ҢU&��5����U�X����{���1q�{�f���ӱⓓ5���;/#��M�P�41�ڳ�m��C��'��C��g��~�򙆐t��f[6�3�i^~Y;��TzY�pΌ:T�On\ʕed2���{��Xә�]�pu�V.e��&�A���n]�K�{ϖ���d���IZc;�D4&�Ն�N�6�'���7xI���p�Y�����0\T��jvv3w����C	AY�7��P��x[��f�x�@�j�zO�.��w��v��ٙ��}��a���p����J�E�'t��;� �f�ԇa��2��Λ�t�S!4 ��a�X�RQ��kR�qn[�T�ֵ���rlڝ5�	�<�w7�\�����ޘ{dIْ�T���y�,p��(�3��|�`,n}�f�w��VI��kEE.�"j�G
��w/����$�1�2;�[b��I'Ԃi���� b�N;�,P�}�<��*U�g,�����%i���c�B��ߜ?&�}�#QE&!�1��ũ�RȰ�Kj�F�)�P�,�ImX�4B#Ac����R(�mV((���QȤR#&5�
e3%\)Q`V[lU1��2PZ�)RU�+m;�L�H��*c
ʗ)r��h��AI���,FZ��V[Z�EU�bTb*"��0�e����	mX����%�b�D@b[�
�(�5[�aRfR�(����+�1�Ee�E1P�r�`��E-�2V�e���ZEq��LJ�%���*R�)f[��}��U���>�R�9�~�����E+DG��ܝ�gɮ��"VD^s���ȍ�| ^4����2b*?u�c#�h�[��;�C�K�¯Nf�ė7pGG��_{�p��R�����3\�x�t��v)��i��H0T��*���e@�~:���&P�S#诤��}		�O3���)��6|��`�t�oѰ���p��!2��0��$���C�Rb���^�Y %*,�d��[�Lh�َ�]��m�ٞ�u"��XR�\�}Պ}a�8� �[�n�S7�[v�D}�����/�T\)�¼*�n�v$������6���G�Uz$`���U��/�kFP�n;�X�G
����r5<P�p������v%\��&z�S�ŚV�2�u�b#��2L8(̥񳢑(V}W�ܕf�:�	"ccVlш�p�3lP�\f�Qٳ�ʝ��
��Ƶ9�'Y��(����;��zLK	S���k�9q|v��@�&	Y�9M��2ڮ�`�������eY�gAX�о��wHW��H>����&�`:��������g�Q}�k����ty}^.o^o	Z ���>F�9���
��-���ت��P	E�Ҋ0"0������_�3n�{&�.yVR����nT������s�󬝽?Fz����=��L~�y�ӷ�/�m��
@̑?��ӹf���V�;��L�/qh��L��^�Gr^tR�ó�UFb�^*>0X����xU�]8��%N1d��^�06挮��h��"��ۉ0]�⳷�YP8VO���t�ً�y}��^5��i��q��^@O|�k�	�� �ؠ�3>Q읡������k��/��S/wb����:�+uֈJ��v�8j]�=���p��]��H��j�)�ݟ5�\iw~*j�͟�b�=��7V�ٶ"U�A���q����+/z(lg����ۥ�&��*�?@ �8H�0�����Ǫ	n;r�vu'�r���/�*ѿPr�"��Ƹ�D�ҫ�S��/�W�O^c�y� �.�rp:1B]b${"�v'�hϟc/qQ#kK�����9�<�=���B�m����Q[[�u�r�c�ر3y+��j���m�@B �PJR��;2�q��Sj�<���()�P1����ua���ǃuC�<�h��<c�!rwv{���t-4�U��)�g���n�l`�C�uxf�����4!��uCMJ�@�X>��H�|��G�P�H���ٹ����?v��Sz�y&f�O���Y���e֛}���F�����a���U��V����*��ni������^h+�\�h��H�h.�j�w�w3K6���@���a��ӗ;r���g���[7�U�^~ȯ'0�s�����2��a	���Q�ᥑ1�/��l�i���Ͽ��@Q���Q�P]W��Շӥ�y��Z��Bn.uu@O����d��S�����Am��[]�Y���3� H�"6�PU�F=^�B�f�ɧ �
o�6/��o��
R��E��ΞB}���2��r:	��ϑ��)��[T��m��������@�f���r	{d��-��pa��#b�|�j����  u2�S���ȬQr�l�?����_��}��^��<5����&�;��������,�V*�Mt��Yf=a:�D9o��#����i]3���t1�я��y&&)]
�MȾ��d����v��y���b���x~�|�������z���3�o���+(p���� M�3l��8�1�Qu�wcf�Ȝ���[�#{^�8_��ݙ���{��(���%鷈�7!�T�9,�M�`\��M
'�O�� ��}���~�n �P��]=fsg� }��(���`�x[*�g޴�8kh/�U��A¸JӢ�K�5�%�k��4�:M��U�G��l�q�B�R��/��s���<5�3B���4Gu���(��.D9.FԊR7� H��>e���� L��}:����~H
2�`jև
T�W�j��>{���+g-c(� ����z�D�^�≬����x!�A��zE���hp�`�o���*#fk�6�A.d8� �X�V:(�'�������B��6;�,�����p������L�(R�R?��8-�������qᵇF����;B�q+.<O@v*���7
�^2�\��UՊ}a�8��Ce����?� ��	*�������[�2��(���:2�^������]�[���S��1_Y�.���
]y4Z���لQ��D����Q�u!�� ��_�vz~w�<W�|������O�Ӿ��9Ms�r���F�.i�n���^���h�'�j��ŝ(�>�5荐�^o�^�~lߔ���M�p<��Sm���pyۑ[�k;I���وP����H,d�56:Ep�lN\�Ko����|��Ik�M0GU���������f##���;{I�R���y:�*LG�g��{ưV�5ܾ�V7�O¸��?Ay��/}��STt���!"ǲ+�Áy�DT{�P8l�)V�̪笫�+بX>R�
��<���U�R��Ga�j�\�˸� >�~p�Dx���R�+K�i�JeA�z)�ۍZ�g��E.�:Ttl
r4t�� �F�#E57R�][��3��X���mp�w�K���n�L�KYw��e���q]�n��O���'�0[�ABYަ޹�0�[�o�͠WL�ܚ�:�0��_������ܯ_H��;����u	s����؞�c���M�'��P�V�p��\�
��/�,��E@=;sXTeS����/3!��K�:��N�0��1��Dt�e�%���p&:�	��6*��}v�C�CjNʈɌ��ӭ^<��p�@p�@�9�^��Ǫ;K�,h��0��|͎<���B��_p��j�g����v�@R���|�JTA�w������(y*�/���T���2�h�z�% ����+���ؑ�N����M�^� N[��!�@��;٦����i���p��	�X ��I�>�V'y}�| C��R�+��7֣Z]�|�r�z��,���#K�Q�B:DZ�J?4�Z�Ф�i���ۮ��vI�<�.�P�͉up�N�ڞ[/2mUk�� yݜ-��~G�>��«4�UJ8<*Mm�>'��Y�#p�./l�����!��\hh�&G@��l���3U*-g��P�[y���zP�B.�t7��dbT,�)I���u�C�f��{ʹ��
�T+�+4�yo�ի�t�u^a�)��5G�O��Ոx�*�&U.;��0\4�Տ
��n�}˓S�P��n�ټ�K2�T�"�M�S�>V-G!n#�>;^�hn͙1dO� ��Dm��7&=��ِa*��=Y��n���&z=F@�:~�����\�.'�CÒ8^���\�����L�;�7$� �Lw�Y�r��RT�i:<�@��t�Qcdl]ϔ�W�<|+8�4��<�Z�}�p:����k����]�=ϊCmG� ���Ėx���?�$��b�!`�@�r�#�Q��F*���T���j5UQ�R�Cdg����6JmȒ�c����g�a�S~ޝ���_i�P����2%�|��Č�.bl��UC�"+)G����[�an]��g/g��i��X����}X��7���9nCKjpeL9�4��e�dDf�}��^��_+��
Ѥ���T�jg�D������p@�"zN��3[>��X�j��߽�������Q-��v�U�\�UV&J�X���<�8�n�\&Tz"��i�W,@��҇z�m��`���%�$�W����3B�q�(���)��?b��@웻�>=���R��+V��z/'�\a:�C�8l�ȺR���Al���p�X��Ck�"\D�`W���O��y��{a U兖������6��W��1B�H�U�l���J����h2�l�h��1�Ǡ�b��P�gq�_6s�='hPwd4�[Fx+5�+T�:U
��=��y|[zE�៣�%�l�O�@�e@�#fk�С2D
�؋�ï�J4k�{���2F�Pt�lF�2,G�@תOK��Y����&�}2M��k�S��z*>��W��(�����G_/����x}^f^������.���T:�O�ԩ�c�O���o!pxU֝ �t>�h�C����8e(
+[��Y��b�`�[g����?b��i��Mh�(����ދ&R��f��G*�P���k�ӢB�Rr�(���+�����WUî=��@����U�C��
3�T���b�S����3P7�b��5X�����/�*� {�3=\����҈���(8ݗjTW�}v� ����[C`���u@P��%P��ř��Qi+��Q�u#�5��;L��5$��1�d�l����3@�jq����(����.v���3�C�ۇQEm~��u��D�f���{ژ������N�U�g�M݋ڑ0� ��3ra,a�=K�nG+��N�F��؇Wm�6嘬�t�2�0��p�Dv!t��n���c�R�J8z�1��SPs-�V�[���GRd��Vv=�J�S���pb`-�����Wh@CճN9�jڭ��>�̮}�^�/�%޳���*9��#Ȝf�C�+*�	�xɼQmNt�Z�(<Ղ��p�b�u�]�%Ffu7Rh;eҜy�U�v�|zf3��K��2�_"{q��<��8o�:��nE�DNa�g���"�v�0���xW,LI�SY�����k��w�ù�^;�ޔ�ɏBݵ}��k�un���KG��D��>o2R�"v��,zy2�f_U�\�|�:�������-����E��h���<]���yܘ�Bd���I v��Za	K��N5s����m:Ҳn�0k$�)�r\j�b�x�}Ϯ��/92C�x쩈SqÛ}�!���:ܮ
�[��.]�!���^��\fvY|��v�-��,�b���04Μ����ս���>
��[�9�H�X�i,�Y�������߹>�
^�u�d.ںym[���e��9o4�t��3F�-열��1
�E���}�ep�nck�ACK����lnn�l��n���)�����ܾ۸���ي'����ް5� ��q���v�1�4N�֘9�ǻ+[�u�1[�����M��]J��Žw\����8���&+�|��ɫ#7%ɐ8���:'w���<�A�u%�*Ώ��G;��}�;6�1�����,q�\���?Q?8q
)mxٖX��\�X.[�X�1V���h�* �T�dDn\�����R�����9K+s10TĬen�W2\��̹q[mAEQCe3T̢ QPm.R��F�2�Z���cb�U*Z���A2�G,,ƪ+��+�TJ�*�84r���"��X*����X+�����cQ+cX��EH�EPX�ŋ�����**�
�R��R(�%TX�YkAR����UEb16�����µU�����R�"��U���� m~M�������-h�Zɝb1��PIW�	G��n�|`x{o�$�����עM	1+�)d�N��5�@̔ �!��e��K{�MV3_�*ʳBZ��P�zڰ��`�A�d8'
O{b�a�b=���YZ��$Q'억In���Ƈ����ڹV����`�:+4�ES7K�]l�]o/�������O,�RW�J�AC���H,����ͲcP�ˤ��S;��iE6Ώl4�Y0嘝�_)
0�
�I���&3�J�ߞ����9�[���z��PY=eH=\`c���T��í�t���������r�l1�}a�������3l�t���+��n�U0��,�'��� c���	��VO��Ag��eUH,�l��a���B��;��H)��a�t���d��2���H;�TY�+�ۻ��Q�\xT��� \{ɈvTXc
�a�٤���ۖ�a�
�����La�
/;�)!s�h��!Y�)�uHD*���*�~<u/��Ƕ�*��<�H,Z���H>P��'L9�H)�+7t���S�RT���[g1����AHg3&�*�w�=�^����}u� ����]�:�a�
���f�
�+��VuE ��(c'P4%�!XmP��
�Y^�(���}C/�W�e�TX�M���X���MKiX1�i��x.�.�B�T{m5Y����Ix�8fQ��i�n����Fu�O��W����-q%��=����ͺ�Ö�\�wvd�;�8_�����׬����Oû=a�����L�%d�Z��i+�YH,�'3�=�L6°�XsT�Ϙui�
�A����ɞR�;��z<�����μ���/4�P:J�a���+'��z��ḏg��`m�>B�[�b)XV>g=��Ad��(��;.a���w���ι���{�\�߳\���冒
}G)��u��}� ��Vi'n$��a�R]s4�`������9a�w�&$|�і(
,����o5��{�}������Y1�/�
�Y0��f�*��0� �;�bt�}���L+�Nϼä��+��Nj�Ag��Ld�*M�:���s��r��>VmĂ�U=f��9�La�
��*A�C�U��*AL;���%a�Y���J���Vi �l��s��!Xx³_k�<�/|u�7ߛ��y�Agl�4���f��ƺ��Ω
��~fӤ���Af0�b���Ad���P1 �CFX�gl1�SVbO����'�ȿ�f���L� ��4 �Xk��
öu�4�_�_d��H
/���H)8��H:�u�i�L>�Az;�1�I�!�h�"�R}�z���3��yל��g"��`+��y�Nu@Ă�^�& (�vʇT�� �g18�bAa��3�J��s6�R�
��^���ל�ǯ��=�}�O�|¸��S:a�i��s(�Y`c&�PR>R��γI���3l����w@���5݆$Xm:�Θx¤7��;5ތ��Ͻ�����+;d���1>I^��H,�;������+�Ձ�R=�& *�8�H,�2�)
�6ͧI���i������{���h��N���؍7���QK�=]��ٌ8IG ���N^�]���=-�}ѱ�l�T�'c�J�C�P�+5�q!Z�3+z����:�����[�n�z�Y8���H)t�n�LY�z�u�I��n�v�$��J�R5�7E��,1 �d��4ͲT���"�}P>I��i?{��<#dy���#��:��Agz�����q� �@�1���\H)<UIR�a�q%d�Y�vq� N��y�u��κ羼������a� b�ROR|��x�;��&�I�{@�$�U�5���כ�u��}��Y����Xv§7@ă�܆�m�@����V|�|�*$���,�Ag��(}��B���LHr��|ɌP׽k�����y�|�o\'�&ص �`s�L+6��SA�ea��5�LH,��d�AH{[%bϓl1<;�bO����q��g�QN T��o���u��־���8C��Vq;a��Ag*^S���̤hbLaX}���R*OMw�$� �G,�t�`��KhLa�S�����Ϲ�y�{���v�R�t�*Ag�ȡ�J�R��G��T���=d�Ϭ��@�4eH)�&�w[�+a^��t�H,���v�����{����'Ɍ�>�'�����i
�3j�$�c8ϐ�N��
�=�R������Ci+6��SI@�	�F�?�t_���b�{���O�bC�`z{q�2V���$=a�Y=f0�=L`z{q �L115��1 �y�]o�w޺�:���|��JŞ'�8h��!Y�^�H,;�Y'����(�0�Av�Y4��*Mr�?0+mHn�S�ha��V��]߰X�<�u�B�/V]ȬG�(f���j�j�V�0��V�l���B�9�����L�WZ�b��K[�o_5Y��K���ؠ}5P��n���c���ޏt�~H�{�}���$iϨ�IĨ�532�`�SY@ΨL`��$%f�%@S�H(|��s�&$l����l*�S:d�9�7�������O�N�*<�Ă�>��R��ۦ�t��R�2c�'2���O5̚H>Ra�B��g��a�,�RY｟sϯC�y���p� �{�C�0�g{�b����wCH
(T3T�X ��O��!P�������z�P�T����>��p<#�v��ռ����Dx(��2xʐY�=N}� ��S�f$Xf앋6�3��AIP����H
,��,18�RjeH>�d���T��N}���~��9�}�m����d�ݘ�ݰ���1���@Ăͧ��O����1��X,7i�&3�h�a���Ya�ڤ�Ͻ����7�/�IRW���|�G^�0�
��*Ag�<��E6�]}`bAN�YH�HV��Y��N�g����U" `� D�
,�m�{����#�pY�AՓ�Y�T*CFfY�|�3�Xb)���Ă��隰��0��{:�1�Vo�d�@QC���=�+V�����WZﾴkw���o�p$>�8yI��j�U �=��H?S1���cXbAf�?SR�N2�i���X����uC������5�s묿|��[�^{ϵ��g�L@Q}Cbx�P�IR�P�hi��+ֵ�Y�%N�H��P̤ćv��]���v_��
AOU'n$�*,��|�~ξ��{�0<k�7LH?P6�ֲ�ä��2VqRT�	QH(mS
A�GtY4��}I���YA@QM�|�AH)�<�s�a��nڈ�Y����;���	��4tP6��,�7±;K���rs�
gN�z0(����K��E+�SdvU�=�d,:�T��}�=�p��������{���]p�!P�XW�M&2t���_Y7���
AO��3Iv�|�T��Y�=C;� �R0�H)0��j���hj�u|�Y�����\Ă��W��2T0��M=0+'^ٌ�'3�߷L+
���++%a�혪�Y3�1���4w��
�l�c=d�������׾�޽�s��{��x����)��2�Y`f���7�8�I#�
��Ɉ��0�
�@�^X�wE4{I��d�,�l
�I�ۤl
����Κf�^��9�w��B��_)
�IϬuH)7�<I�6�vjɌ5��̂�z�u�4Ü�Ă��T���1�����X��|�r��{�{��{f�1��W�,H,�n�H
)XgVi �3�²_,�M{gl4퓴����%v���:Ф���$�*A�΃�&�mP�/6u�w�����=�`�t�'7N�R�����
�&j�l1��Ă�a���6�PS]�I��I��'3쓾��T�|� ��J��o<z���z����aXj7L6�&v4��YNk!��E'[��}Ciצ�����`L}"�#��?4���cf�(���@ڳb�ej�q�;���F���K�eֈ~����=����:�o�O��m�1��%ɮ�}�N��H���V
Ԗ�^5����g*eiu�U�tQ��͝�C3��bV�c�T.��Q��Wv]����(��cM&3��fdl.�y2w,-�k�Ѿ3���#}\����Rud��ū�]�n��T̏��� �e��f*��v8@�> (p`�u��W�
��\E뭦��T��R�F)�=��U`,:����_y�U�,,�;�^�+w�:���\���P2!�L�e�Q�/���L�vI�s�;
��~�.(A�#�E�-+z �H���2#���2`�렔�&!�B<������
)��Kb��3�4UfԸ� D=�Gq�W��̵�:��וm*&o&�u�@M�nxt��b|1�F�zyP)��vn�� \Tv�\{cb�;��s�I&.*4 k��~ZpX�M`�C���[wXm��]�tl>T:����b���F��dP����e�{����J��C<$Y%Ǫ�_Lqt/�k-�e|S�b�B�4���iBltW}]�2�׽X�ǍֶG�v`��v�[��A���wi۪�Y�����xu+|�u��7�Fv�qV�ؾ�Z���T�j|i�2L��̵T�5��2�/6'���S�P��C�3Y��*�8�S4�[q�,��z��V
�J����D����gk}���}u��[��ڊ1��f��b�^���X<k	��c۪��/���aoo�r=�+Ν�fTY���
��.RU�^Z>J2L�{�gF��Թ��C�U�R�<b�=���q��39e�s��J�����b�z㜘[�c�m%"�d���g:ꯛ�ˏ �`ȩ��@���dl\yf�Q���1�b����t�]p$1�U"��)1�\� �X��㛷Caw���@V	B�혁 ���8:DVS�7>���١Ea
�W��v���G4�0;|w�r�^�*ܳy��Z@��{r5,�<�1��*���fm�\��9	2CU(��L���r��� SZQOd��X�$G�@Q�]`t(
,L�����.�[����SI��Ȉ�$l#+���顢�<`�AF��y������*ɵ�i���+�H�Bhu��3;�U�����J�v/�7��O��e�m�.�k��m?t��f�.�w�e���@,��2c��7"�.H��f���q�hY��K������u�3H��4E�khQg8�m��o��3y��_��	�T_IFW-σ+>f��a��9[̽�\��S��']� ����>�� p���J�0����5�d�0AXf�{
u��-5d�ʵR�_Qշ]���V 9��NC����ݕ�<*
��^];MOW����g����Y\����}C�G�c����T,ޚ�6ެ������,f�$�w��/�D���9o-�W9�ʊ��i[����F/�"7�����i���X�h*"*d=.���U���g��/�}�
[��-^�a<[�&��\Tx8p���^�^������dLْ��Iy��H�����Łax
U]��3,B�kI��`P��e:�� ��,Nƅ#�@:���uM�Qu>thő*��b�s�r�#`.��^�*�����dՏ(P|}��@��"��j�bݽ�=�̧�����Jϥ���+�U{���xA[V@�A�����;fnw`�ǡ ��t������~mSr:9>Qs��m�盼�U/&�
~�� X�>f��ʙ����d���y�-�f�hFɏ^QA�yO�5����[��˛ۻ�p6qxW�\˴��#;:���r��$�WyOǇHCip<H�!��"Ήo%d���I�B���G=%	��t�2��T. =���;Ŵ��*>�nzd>���A�0'���$Ȟs�v�/}��Ɠ��X����=�Z��û& f"��C�ʻē~	�f`1s�}�kj�9���-����G���&b-�͝���n��� ջ�\�
4e�˜sى�s�񝋋���l,�X�}���1|�/���%�צ���!�(�#F*�>�&F������T��[R�Y��f���0rL1rP���M�@BM<$�=SS���v�E�B�`��n�(Y5�_��\T"+�D�Ʉ�vwkڲYr#�'��D)�ʓ����I��=+�@��H=�]�|���X��=>ٗ�"EPFl9qj@�z:����l���r���m@rM���`c�!��osz�lo���%]vw(�cq��M�mP#v�ᝰ����h���c�w�(�n��yV�ͩ��4��]De����4��v̳75�էL�@�ov*��.��k�)Zt�e��|x��A���_ABm��@`�%꺆:∈չ�f��|�ܧa���%�%*3�Y���6t>�)�WC!u��!�"{r㮼7�h���x61|��3������8���%�u��$q�l%�T[͇9��y���U�ٝH�y�:���[��_Ns3OXN.����Ʉ,R��р�ڭ�:4Q�`��br	<SZ�)(��7e͵��9�z�Z�����X��o[W���tP�M�x���b3�,,��h�uNޔ�'Z:���N���[��`t�"��4qVJ��o'sCu
(��R�R⣮�*ʎ�>���8���ǟL@6��e���
Ís���7�'ݽմ�U��rY�v9�v\;Y����ƺ������DS&�胿���U&�׽բ��Wk�g뇤y��KеWt�9XCN�/G�c�=��9�jǄA]nYVC]�AES+���k*��	N�P�ݴJZnd�0^�w�Լ�&/2=���F���=Qp�P�v6:�&ꗭ	3�J�=4�C�ux�~Wke���[RPH+���s(����V+�m��M��1W��ugXӛI5o�T�"�����bU�mȘbK�3e�����w�h�	�
��\�6���䴽5���Z:�
B��:�Ȥ�l���tո�	v��R�׃*>��d�'7�fnڼ�l���GѶ���j��.��̤��VV��Q���+4�U���}�TȊ �%�v1&�^Ĵ`+Q:0�Ԅ�3�Oa1����ש�Ы���Ɗy�:��oy������}�����1墑HΆVE-����TQ�X����b"#�KKTZ��b33��D�e��A�(��X�T��D�����T1�q�Q+H�b�"�����PQR*("��Tgm-,����QK�X\V���ʖ���cR�[+�$�(��-������cms3%�Z-��!��*�Mc"��f.%(�mTDDEL�U���cs���
8�����
��ѲP���VN�T$�(�����G�{�]o2�v�B�ă7��]B@�#�hЈ����n��t����ñ��+w�,��d��H�0+� d\t�A���Ƽ��Ԩw7ܝ�3.2*� ��3�["��t	'����\���k��ԡ�oY���u��@1�PѠE5��uf�[�go��ܾP�����Rg�#���}�Ur��>5喽��Y|�y�3�<��|-IsPd׫�..){>���X�;���Z�Q��bF`ڃ>�q�Q!As��7�z5D�)�w��W<
��huZj�x��b�񬴪�q�C¬L�Z=�h�wyٮU���~�?t�*�/�<��qF�а�C�Ky]�5�����!�۠�k��8Ϸ���Y��g�}�";n.D�;�l~��t�t�bi����Q�pG"�{ܖ��sx*
ŭ��-7���{�����f�V-��l5wa�r 2﫹$&NZ�Z/����ө�����>[�PQ�W�c�R�Qjv}g�����E�+�x�4���*���Q{#b�|�j���b�1������j�R�F�H�R�|><ja�K������-���g3�͉FO�)+:�Z�t�ҫ���3�h�9�I�|b�jĎ�#� (�ݮ��RW�Eю����.�c%Rؘvr�Xt܎�Z�}J�����],=����^	���F܇��n/eF�@L���:EL�o�=�L��E@Y>�b�_�eR�#�V]{Y��<��&����(�ۣ����X��&v�*�k��5��K����t��H`�*�hC�0�j�6�ƈ��PVЫvO*��2�n\���M>^'^��S�'�IO��G<��I	��o)5e�W#u�k��z#�$�:�oF(MƴչR�C�j4h�zdP�I����ێ����{�YE_Y���>*}������T@�����qy=�ËWJ�|R���
��i�G�U]�gEm��@*��4|��W;�m�=��V�E�
2:=�*xl�O�@0�i��;7KI�!���^�L�p�X�Xc�ʋ�X���`�G6�{\�N�,�q� mHExL��cӳ^��8f�}doϏ[�OE���>��aɃ2<!ˀfN�Ԋ
}n\����Wgp�]����
���
�Ϭ:� ��`p$���dp�r�J����3��N��j���XR� z}'cB�q}��s��Հ]ק�i�U:2b�}�A�yl�zh�N�d���G��*���h��(�z{Ǧ <i ���A�<(�wFE���D�ݹF��;��m�FBaͤ��=�)�42�:	Fdq�N�	�4ԋI�$�6�Z�7�^X=�튑�p��j�,�[�٫W���N� �>�� �S�Ŵ�d��ES��jj��qJE�&���;��Α{ZY�'fbL���G�$�葆we��Q���׭_�FF��S:v�H��i�3J����f�2����x��<F*��<��A�����8>���~�������A�a�Pzs��J�`ʊ���R�.ȉ�'u��Mu"��}�7�.;��|����h�;&�L�rI��� V	.f��ӡAIs� hί��*T.�o5���2A�`���
��06�Q���L�L�9f]5[z�w��%v+զ�ň&z�������890o:��'U<z ��f�]�G}Ƽ��S�q�Dj�Tp�aq��~��K�y続��ee���D�t���hu�l7pٽ7x���h�)֝�%!���<U���J(��n��:v��[���.ێ�ܦк�����7�4��Y��ͻR�LT��p2���܁2^����f���|��>,k�G��3c�/���Et��e�T����5"8O�8bdGM7Bܨ��E\��s��t<�n^:�O���Q�����U�����_�����{��^U�L�����q �i_4�`�ʥ�~�������x#N���eɁ� �����
=#���t�ȓ�s�w��_{��P<����P��f�x���N��F�ook���~��z
"��G��]���Z�=ڀ�#�H���2��;��N|�Щ�K���r�qV�]��z���7r���j�k⸭��ve���)I��k��_])��~����P�Eg=K��.���_9~�2?H��2�q%ۅ��9�ꖛZ*ս嵓c���O��\����w)M�oo[����XE���{�]|�5�1�6�9ch�бC+j�#���ϟh�H�ә׻���j��F�5a�2����u��蕺�:�e@0���ؓ;���UyWa��n�8��Vv��ؗ��{xSt9�8�4?�sJx}!t��^�t�$O����6�ۜ�|��O��詑���I���MpC�3�G^[�v��z�J�ss��'�C��^�b��q�^�����Ն>��{͋�">����������0觘y�tWۣ�3t�S~���goo�������^�$t	X��F�Q��mV4��vF6�=���x�y���2aKF���
<�F�G�B���yc�#���+�^V��Yb�K������R����?��k]�A���;��ʷ���K���uʮl�]f۾WNWm�QR�f4)aݤ��b�A����c��h=�A�i���D�m���OQ7�V
c����ғnEl}FUW�(�.�_� t�Bhu��7����U�f^O���P8����������ƫl��g�������#�\xQ_jdخ�KE"x|�|]x�B�5��c]CY�����Lz��/�ƴ1A�Z3F���4EE�W�7���<�`��K�}>��#����&b�=մ�w\���C��<�遐P�M �S�5P�� �P��P��Cx���O�IXˇ24R��zd�P��Jod}j� �[{�}n��U�ɗ�Ј"̃�B��^O�'����ս��*�L�e��
O����
���#�W����HR��OrU^MR���Lt0`ǃ� �Q٘p��b� d-�,Ʉ!���`��1Pvi��F.Q;Y���є9�驖rr�����K��0f�		M�s��͕���e]�;�j��fD��j����
�z��`��@�ٟ)�zp`���&<l�MM�ٞ�+C�?22��p(9��7aC�<g�тv2B&*G���A�o����;ʿnu��.=�G1�yt�vF���U���'�a�IWC��D�x��<0b�:�"{_w,�Ej0�\*�EW�W�l�$�K��Lx.4����:�&z;��P\`:~�`4,��G�����V���E*��֓��*=��(&jz/�_i|���H������}���*d� 2}����FkdFm���W <�����b�<։��`��v()�=9�J�a@7A�tыJ����љ�0��B�(�k��1�,�L� �~	�G�*�H����_�l��u�-�.��fޕܭ�I����9�ʋ����E�f=ܥ�
�l� �=|╛�F�"��������O{vz�b</D�;R���)��/���.Q��$^�~6#�^˪�`���­R[A}�Z����s��Y��*�v��GQ�ݐrL�b�#<##�H�U�0K��:^��|ь��_
���i�9>?�j��0n�)9Q�9i��&'��2,m���[*0\��nۜ�$�"M8G0�[I�!���u^�& P-M��0�z�a_�_�8��L�u�m�q��DK��#��Qb=�W!)\�ƢF�+n�u����JTt�?:�t,4ˇ�����gb$���f���� ��vu	�#�hЈ��n�ʷ���]�{�7���A;�&yw��l����*��c<6���x� |��Su�;�][$�R�U��ېNg��k*�]�[K]L�>N��b�2�U�,[�dl��̶t��@a�Ք�.0	���Np��<<5m��ݛ����ŌJ�oΜvy�J�����.a�l�<�!�[��:�MP팀b�PT=}j63]��:���hرL�#�	��Z����=p�0�t?F�A�Ԧr���]{�dݜ�֟rW)�Z���tp�O	���-M@7��qp9H��]�궙�^cf���K�#�X�RU���<>��ʩk��d��ֶ:�ϥ��N��Ç_�j�x����yVT�q��ެ�f�ZiE{�Tn��R�|�+Ɲ�aE^�QJ��=\�ojN��&$t�1�23�ʿ���M�]{�#T�I@�+����}�gz�nz(L�nk�P�� \vF���PV�ü]� �?y)M�t�N�>�c�������v�7���]�zת�.<���7GOxn��"l��o�2�faN��N�e�fT�F�(��������ј/%#�cw�tB���O�����!y3��ܰ�*6��	��ǒ�"�M�KtY^�J<����]��!mͮ��n�wcm��o��4Ǭ�8WWy�q4nM��֘�a����.Xy�W��Y�H��H��e�����o^�0@-X�;О:�l�����0h�02[J�^�s��#^��9��<�+'�s5�w�v����2�1�oRw[N&��ׁ������wj�&�j�quH�˖������s;$#�9���`��g#����}d�tiN����t�g,g
zC�G��ή�Yu#9�JAMRG)a:УG�
�굽w�KZ�*�W#ˊ"nc�pZ�6<U	R��Y�coyes/J�H]�TUM�C�@\T�˙���F��M�����kn��{�= �_�3����|.��2�X"����f�bO���Ŗ��G�
yM6Vbvo+
�T�.r������9������s��ܳ��&�=�N����T��ώ�V�����F�����X1rŀ��շ��<*�m��[C�=�;��ȝ��t�sM�fQ��E�r���� �'k�
R��g{3*��,ORr[ߜ8d�bX��8�GX��P�E�h�@�۾b�&SBb#�h�tI�4���M����r��U�2XY���[B�XX�9�������WI�5)��X>�̥)�̾���/���m�5��X��y(.*n���ݔ�Uϴ�ܼ�b�E9��5u���JU(
��]	r�Y���[��q��TF2s�i�=�;';�h�KB�G�`�WW&��1�
�=;%�!1��X���}N휴�vo{���G�;��#V=%�J����Qc�6UL����V*5ib��ֳ�UcMa���EX�TD�ETPb��V����R�F,UTLLXi�
�a�Q���������IW�A�9n�LTMը��F*B���Xj�EC�`�1Ln�TE�:�C�U������"�TEUu[CQUQq)R�Q�U��\� �
���K�(�
����R @�� �9�N���*��Ĥ�J;l���7)�K��6��WMD���+M�"k?~���w&��?�{}:� ]i�R�b�B� 4���ʅ����,9�䷢�aK�X��R���0H0'f#�t��P��o]���u�o��B�Pɇ-���x!n�G�E�\F��㶞$^h�����/r�Z��_LC�hDH�(WJS~��{�{/u[)�>(M��Y?!�Uzy�Z���V 3M�O� ���v�	��i����ң�
݋�	�W�ʦ�`R8���2�Z|��?#V
傊�L�+%]/
TL���3���"�r��b�\���!�o��)Ϯa��-�hY�5h��k�^�|�I=4)�HB���3�lߺ�\`2���4���Z9x��=�����!���.���8v;
�����������B��ޜx�K2���8W
�Q�8k�9[�%*��	t��fvGN]�u�D� �z��Eaw�	&�u�KaOXة��YFU�f?r7?C����b���/~	��2�`Y��
B��c�%N�I��ip;��_'��#`)��"}B�5�q�~X.��{ML/&yg'"e�rT"9�ܛ��c�R�*&�ţ��U\p��X�AG&�oPV~��8���xt-:+�r�'��4�8�˥i��/2��;"`�&�:�O��s�:z	�� 8!j]�����s�.:(�����X���Mص,E�>���j�EYwT���c@2h���FT�D%(9�tġ�,��t��m��O�C$�'*���ӓF\:���P3�A���E3�ɻ��謝�S}"�O�f�����MW�J�FMCr�P�xK{A�DNI�s���6Vp��Nz��	��φ鳯ß��VXg��^�N����V
@��e��X�|�]K��Np��G'TVv����Ho(3�ww�(�p�!��3��腪z�6R���;�0����|NknIxk�
�P��U��w�O�կ�k�E����~~�WAz`�+�=C]�2� Q`HmX1*kz�t���9��;;�s��G��S`u��(�{��^ɿ;ɇ��M��C�����{(��!������c��x�Ѣ�{��Ȟ.����&R�|3��=ꐄ\x๡A�s� P.�%gsIO'�X4X�5�l��`���'hp�^_-�M#Ŷ��2����w[���,
��lg�H�>�ѳ�#�c˛��sW�k����kB��ө����5�E�{J�ᙹ��,b���j�X�C�v&ˎ�	͙�W��s��d�r#d�6��+$���ت�*=P��9���f�_f^����p��}��z��ϭR�Հ�nRj�̫j10�T��o����\N�c��̰	�K'e�WL_eŒ�U��'&nV�Cvn�
`����	m:��Qb0P�]/��d
}��>�k���3���	���s�2�|%N�l���BC+�3�{I�Z��3��k˦vuق��,+A�(�g��p�c�P�%ïRZ�B�{;���j�/V��� l!�)0���`tD�D��{�Qjr�I�{n�9�+< C�1|ho��f�EJsN�V�z{�p*J�r2/s��T���|�0�O���ف{�֡|��fw��ZH{"�Lnz�Ū�L`��^I���uy%�&�_�͚���aXj��r�۴~�S��g��*�|������������,�LW�*X�xl�WDؑ�0�ђ���/���L��J������iv,�����;��T�]�o��|(�*M^�Ok�U��	��*�^�D��lBn�U��X��y�hkpmL쫘OaΦ:톺�۔@�	�K�G���e3n���z!rFk���v�h��=�X�i����0`�Xٮ�>�y~.B3�ʋ9^�׊��M���q1�>(Fت�8��1��A^չ���s��ϫٜ�T��0�[ED\��}>�(D@*'�h���ǲ�J5G;�]]4�usTzEÅ
@QA��X���pQ���'��wL/��x.r�HU`��� S?,��0��.�C1�����~���,E А`N�GE.�b{M<d��j��"iY�_�U�Ʌ-�6'�,G��6�7��+o�;��V�&��xhԚ�Ʋ"�hDH�(WJS���zzK:�*�Y��U��}��/�^�J����� �����D�&�Q%�P�36dT�l��H1p�(>�W��U7; �[���6˺2��+��9�t��k�� 1[I��ʷ�A�a��*bBl�h�c.ZL	��b��\FӄY٦�1M6��%QZ�����f���}=�G�0W��_Y�yh��e�/
q�8�7"Q6ë=��`���dc�"����kAMP�FKA�F���uaܱju>�MM�^�� ;��ß"k�֯ �Ⱦ!������޷w��T��|���������yȣ}`H�V,l��)4bltη��"(\�j�*G
�ؤ��p�ʵ�
и�5ԛ���^{�����R-H�:FL� ���43�~wt�U����	�uּ��؍�d�$s�#�Nn����p/k�"��cD��=
5O���3pJ����T�+�]3����Żg�[��%�ʕ ����|ꛟ!��W���	�E��ڵ~��*�8�k�d�2S�u#\�t5K���S�yZ���蹷��sQ$e'x���x�v!�ӛ�$�:+�[�n�Mo�4�i5�D6óa��q�鍀�d��=�����R)�M��� �i�����VE>4j���(x^Ѷ\ w�X*سl={�Y���n�D{vX3��"��Rr�8>j'�x�������ʗ���� �U�
���ࣔ~�+� �?{�:)H9=��]�b娝��R�Q���_p__"�(�����H�5���f�5���ݛJF@B$d�
C`���?k��Y�����3�����߷%Fh�$YT:�F�N�躔`U�M�TإNVH���2�ZM�J�WK�xx�X��>b��3s����'�)�~M�(�S�}�{�%ic��˦W�}�C����&uYYh����A�3iT
���n���o*��@ӡ��b<.{�i1�;]ăD�:���A�W;+I�]�T�Õ�F�ԝ��h<��x�6:t�#/��I>/(�u�}|k8��}jz�d��Drt�u��x��ohY�=��~dЌL��w��:���>E����8�$��"��y+����e����/6C��AQ��D�U�n�B��T�l��w��$�C�ȀQ��2�v�l�R���v�E�A��{ѸUM<�k�<Ɖh��B+�q��r#kx�g-���9���)�*w��H�B}�V��5��2���x�����7���V����Æ�@C�:�w���e��k,{�3����37RS���c�"u40�D��&���7z/��1��[9��G��/e��� ]_vrs�:�6�n�em���ыV!�S�y�{�us�w��5j�NzU+�m푕�����6՛�/Iڴ��ʬ:T-D�B4ELbo)O�
�\�y���(�C�R��Ote�Ƶ��J���r{#�����ܪ1&t*U�F������\�l������ԯ�e�6U6���Ò��δ�^8L����J�����*{�쉭�V��E��;��		��zky�;Xo�W��E�u)���JG��Ff\^�Yށv�y��C�{�Ű��! ����Y�j�m���g���W>���L�k��ld�GVĹ37w�U)1�H|ϙN�|��]c�B2���w��;Z�<��dG�8���}"�(p�Me���6�[ ��r�]CQHT�Z�ؽ�<bm�O*���*l�wl��Bִ�ZC��'I��t�EX������\���tEp��io���&_����jU�x��*ǻDJWz��kI���=��R��]'�|��l���Knu��W5k��ҷA�:��Fsft�`�>[�7"�	xJP>{K�>կ7��[�71���x�t��f�V�ec�o�:���`��=c/
��D?9��z�_��*�;R ��=D�Z�P��P�}��x W���^��;+5�t��H�����7Q�@���r�:D!�C;O��������*(�| ���6�#n����Y���q�zw*���71=��B�X��:�hGc~U��m�_w���\�Sq3]WV:��-7�|�c�e�w������#���j0pq�QhOQ���[�_&�T�����l�)��L��m�)�ij���n��ې,�x0��Ư%7�穬�y\�-"�_f�h�5�p����M�ީA�
�ꚺ��J�n8�ۆ���9�y�X�2[�٘o�\2Ԭ`�e���h��.0�/E�y�Q�S�.���yަ�L� �74����E�^3\uV)g{�k���Puf�S�ֶ�6�a�:�ׯ������^k�t(Ru)[�g=���Z���6�?T3|�Y�璞v�����8�6y��w�ڙ]�ofa"�2��-kQ�\�ܔ/�F��sI�s���j%eI�^�Qo��N]�EY�y�D�ûǐ	�׽I��E*vTZJXՕNvrZ��tkg{��ɐ��aB��f�d�:H[3;7��nQ 4�Ą�m�.Bn�}�Fs+Ee��jb��r��K��=�7b�{�V.�ԙR��]0취�3%a�^��B7O_^�Y�t����jTle�1�e;K����E�R3w��[�fm�X@ �1�)��ʧ�R��.�^ڎ9�]�;
Ԭ�
ev�e鬫y:�HJ��V�V*'(l�rt�&�kv���g�m�6��Ayi���n�7z����W
=:�:�_7�	f�SU��Ɗ�\O	�}n�)P�"�f���^8��f�E���s6ۡ�Ą%��6Y��ˇ�	cp:x�tVr�I;����nu82�%�J���b�H�=U��a�\��a���n�{|ށ]Z��Zvl����Z:�h������5�,�ޜ�㿎����ȩF�5]]��j��ڣ).:�Z�z���Q�܈3,��U*�v����Yu�"���2�+�U�%�VEDH�mH� ���kD�6
*�U���-U��V�X(�K���*DEQ�\��0b*,���"��SՅX�Aq�F"(*����+LVT���*��ED�Em��KiiV
T�E���U*T�V��5C2��*
�H�#"ϭ�ƭJ��b��\�ՙ����YPXe�����/�����gཛྷ��2�a��a�fŜZ�-��C�LQ'�D�L�2���{�a<Sެ��atޢxF����W�]e��-�s�~��/{�G�|�Y=�#ӑ���^��ٔ�Q�lCH���6�=�x�k�GN7�����FnէS�a0��⢩k��=�4��QVOdl���$���8Hu��D)F�r��:�.�h옚kV�a�·Qӈ�E�;F���٧e�W�k���0Ek�KTa��f39�5�|BSӰ�ړ�Ce�&���߮�	Ķ�M�����Ǉ�t�}��e#�7})f��3Z���!+gF���o[	c1��������e�R��i]���q����\C��y;h�)D�*]0���1�
:���U���'�;^��$Ӝ�[��0�'�8Ek���+3lT-Ď�����f����Gfu�N�m��M�⣨d��p��uq]�*v��u��y�7Z�n7�C���āö`�Jw[�Zʒǃɋ��ſ]S��ˣmY"6��Q�Us�Ou�:gk�T�	�Pk���7R�x�����a�3����h���p}�96����*-��{Q��,�2﨑�s	x[��q�P��6� �b��T���.�S磍��.�F�u��u>�x�n%�^��2�����MY�����*�"��3�/`Y�nOZD�Z����o9&5q V]/9;�D��'a��C��"3F�7g+{��r)7C�����n�0j8K4�ooV�{=�x4S�u`)����j�P��h��m���a�Dۻ�mU��B���C��g*��WF1��8id�x�� �5EV-c1gw9���UK�)鮨����Jrr۫#6Ý뻦��ݬ\�KveR�Ѝx���R�����I���θ�L�Is�L�W��`fHl�o�$��Q���[*�gWW��2w�qk{�~�Ĭ�au�\��K�Π�c=���$��Jx*_�����ճ�Kr��eFF�o�}�w6���adF�u�f���2��70����ܰ�F1�^9���pF���'�n��;����ډn��Bp~�9�V@9TFfJӑu_���9?���]u���ֆ[���+�\�V��;Шs>��r8d���;d�d�|`򮍓��8�[k-OZ�nR	�l��69��x���	�U28[x�=�-�bI� �=ɷb�wp��E�r�m��6��0jR">�W�W5��% �W9:�k.[k�9"N#*c]�|U�i�h�oR����V�V2"R��
yOk�X~B0ĳ�6c:t+�eU&�muۻe>y��o��~������)w��jý-f
'd���L������,�I�N�ܳ�*
����@��Ȯ�sqlk˯��v�E'sW'��'���}����^aj�kNoeq�/��n��99��|�|�^�E9���GЍt���H�Jčџ�g	m�B��\�����/��;[9�{'Kǳ�B�
xk%��lb[}�;r�Cuv��4��ݩd���"F��H��{��li�CkS����ْ[JBޡ�ݝ�pF��>���n�s\��e#�����H��	��[�M�]��[!����&�bd)�x�^�s)�b�]V?I�mS����Z�7hb���8�^K#X���j�s�UجP����t� ��\��^	C�;� �j�s��J�m��.��Z^t"��߅���g�pQj��̏�&�=[K%F��J�h�{J�s�f�3�x:��Ѵ���������\�Z҄�ޤk|�8�^�]�"K=,t˼�����k�i[;��K���ꐄ}��(��e��a�K0�ïoz�J(Bɘ�Qlѓ�R�e�L�/uV_��孵�:�7�ٕ|��r�v�'�f(���O׮��v�!.�sWe{�)�۫����o�r��m�o��<rp䞫��v�/^Utq��/�oD8ڨ�9�Y�yO4�)��0%'{]z�$H�3];jb�S�4VS��xg:�'�&u4B��U�Zq'���^��i6���|H{}aOP�j6���*�����ĩ)Y�����6��řrkQ�Ypp�����׻Y).Z�s#�r�ɬ���P���f%ް�u�KUv3ٯ�SU	���Ҋ�5̱��Q����5�ǲV�@ZG.�"J���_{����ş>�tk�:p�郞,GJ�S�$�F�yX ��!u	��G<�h�FݬE���'����$$��p�DdD����'�ӿb�o�6!����w�a艻+��%�/�"W2�v�l��Ewq�z9Yة��m�R5�!6\m+�)�@���W�g
��\^KA�,��Y�-5V5�ΣY��VB䓖c����v�l��8x��Pn%��M��;)��*���uD��ՕV��.�[��ൎA������Z���@���P;6�rچ�(�#;��x��h#�B��~#���)_f���`-��鹏d�e�Y	;e��Z���)���b�6np�h���z�u�CR�=��X��h����9��s���&ӧ�]�:���S�}:�Tr�O����k���<�6n !T��gz�8�I�E,�2�x�����z����q�b�G��:��N�d���?�,���wf|��lvua�$��kBພ��ZGE����s�S���;VRV|�0w��3
������t_W�m��#�u��Bɑ��ʯs�F���QEا5���&�R}0�	��B�����6�E^��U!H"l�Ua%~p9�ؤ\����;d�Ч��W9�'*p6��sۓ=Ϫ�gR�*:�TŇ��0�sZ ��m���_�{J�t��A��K���3�خ�e��Hn�.���U��Y����&��jfM�6�(􊽺DMg���:���|�Jͭ&L_#R���[�Z^5ՕS]�Z޹��%z�ӗ�Anѯ�v]�!*|=�%&�<vN�+�=��ڦ��W!I̮���X���'\������N�f�L儺���9��Ҝ*~b�jwE��"l�Q� u+έ����ˇAN��D�+��ym�n�������֯�7,	T�>���f�)s�����N����{�9+��>��l�P_A�����5oѝ�'���F7�U.������o��TɅ�́RzIka��g&�ފn���|��{ �J3��2�$]��+N��]�����$�+Ͱn�AT�Q���l�.h��U�oL���;P]�Ibu��8,ِR���oZ���Hϼ3��q��9�x&f7�U'���u�M�e��q]J��\d���N�J�rʻ�b9B��9���gGp�8@��� �R+;�˸�靽�tc�
��P��l�F���	GQtK=ʰ�]
�:�p��ӣ�O0�f�j�h�n���R���I햤y�{�̶�[8���鵩���V��5�7J�z -�s�^>*���cǤ#��Iŭ��_�'�>~㞩�µ�ɝ���/����4{Ճ7��D������-,�}o$��ޝ��p���^�2*2q}YT�=/g"���
����4�ؖ�λL���/��%�:)�o�����t$���:���j��ƕu��2B���_e
g!��F�+Ol�o%*K2ե0^t�C�'섘)չC�]ƶb�C�f�4�g��@R�����J�n �v�������|�Rr��r�YkOi��Ih��o*S�B�u�R�7z^�pP�S,�J�,�h���8bLч���{�����+�n2�>R�_]�bս��pJp<�#"v��3�-���f�
؊k��{HX=X�r�tJ�Q�G%��	�.�YA��j�۶S�m�v� ���Y���ˉ�EѓZ=}2�{C��ӻn�5$vk��Q�grdW*�Tr��U���.AgP�jҾ�u�β*��i���,Yoe+�e�v�ğ �$���8�*Ň�j_X��E2�"�.A�[��l�eɺm}���/d�y=��cyr�Đ�.i�jW�,�ӄ 
/1eCV2!�fh#{gJ��ˬa��%+薫�uH�
��ʽ�hb�|I`Ԭ��Tn�#W�]s,�Lei{�#3��*ߏ>�xD#m����0Ӿ������FT��48�I��-��Eb0�i��1ʸ����ݧ����݂�����=�MjJG�:2qB����&���ǅts:�2-�y�4¾�Ȑn	+hLn>?1[7#Z�%|����i�z�к�Es�d�l�X�h�c6���h��z�r�۲JV�����F4d�����/xYz�5yؕ��+x0sc�w�"��e;,v��;'�>OMh��.�\�2��Zli�٨�����:�5�o
{]}r��X�k�r�KpB�`����ʰ�X�:�hW_g}}(�t�{5�s�{���}�t�:�^�DR"�(�rՊDk%zJ��2ʢ��@X,�Zȵ��J1J��[`Q�F((���[,A��µQU���+�"DB��C
ĹTXT�UX-Z�Q�DQ�d��ULA`�¨�N!��ШQ�AHVT+�%-F�BbDI��YX,X[V�Pj���ł��k,(t�i���EH��U�陖V�!X(1�թ�Lq*�*�c

K�J�eJ��Z���CIYwwww��"VR�aD��,<��L�!̓��Cz��j��.��\�%���{V��'5�.g������/C]�t�ɛ�+�qG�d^���qpAd@��:Q��T�p6q�-�{v{eW���=��4'��˦/C����>)�H;�*eGSrzA�m,��:"E"�K��m�1}퐗P��߫�N�a����k���2U�i<Ew��x��9!���Vn�{[V���}���W[r��0u0%���m����Z�6��|
�9EY�h1Z��� =��YJ�:>�t�h����B��!��qf�i��*��7��97t�Si�~���U�ޥ���pT˹���\�Q��>b'N��Z�s2.>��I���զCC���Π��=�9�`�}�h��5_n�ů*P��9w�	G�n�x����i�wؠ��z7	�Yt���v�W�<�������Yx&y�9�>�Y�&D�ڷ��.����pC+k��.&��ޑ���NM5T��<V�.���J�ҡj5"�
�9y�#&�c��9?���s'yZ���ڊ��Z���~A���F��a<6U�خ�O��(��y�Q	�Qd^���/5\֫\�q{̝���Ar��w�.Jjy����w�<_V;���}프�q��c����NսG2�Wm�u��f�$�>JO� �:�9���M�u�u-����WV�m �Z�E���9�
Y|�CP�	���]�7E�|C�e�b��'7���E��d�;�j:�X�g%%�W*ϸ�z{2]ѿ��-�����u�!!$�����-@�����o��x�[�m1c�oI��N��D�㞐�f�8*���
j����%_si��\p���GXT�f��YsM��	]�.�6�+!��Z���q(�/p��i�R��H���\������׻��Z뇆�6����q�[���C�l��[�� 񙊧{�
��OIT1�*�r6�a7�U�u�g�v��+7a�ޠ8T�0���E��"l�z������5��rj��m��@���g�;�Lڮ�M��ƆCM+�j��c2�����4�2��COA��޸�x`˒ ���Pru�����~y���|{s�ӱ��X�N�֥���xwY��%f���C=1����=�D��d�"�i��ܖ��Zn�9�O����]���� ��"��ˌ�7�y�,x1�������*��߲��@)����a�������&��28�=h��_��C��31�AS�b1�)tZx���3����+Ѫ]5���UB�,׬���=s�ɳږ�x"8f���J�'/bfsV���K�7�-ތ�K��1j���͎o^>�7Ƽ�Q���o�4�m�)��g]v6^u���Y�[�� Gj��%�	Z���1$pL��c70m�4kVzǶfܫd�����cG0����N����\�˚�<���Z���n]L��l�kpoQ�F��Z�s����q��n/�a�nM���۽C%ҧH�����B�/�#��FoHxx�t��Ь��oR5(����F��L9\+-�{xd��w�i�q�wP�f�:wf�0���}���<���p��h�!Y���4��=ְ��1"�hiK�͞$����_Q�pYAkD׊��r6}�����>���+*X�ivY42U�^V�S���.��~t��P�Vj;��J�Ύ��AᲑ�,���j}���4��_se��T�r��)!��zױQ���@��]�� r4���#��Qf{0�4�P�e�ΎS:*�����)l6i�{��ݭ��j󌦥�ƭj���Y�إ'2-������Qrn��=�p��`�x~�Uh5)w�RV�..R�6qj�ʁ��EC���T���C�:(��9z���i�%m�H�o�����w�*��&�W����P��1���6���"p�������5�:tu�	����I��l�q�6�^�i[,0�K=���Юٕ�k�ܒ�wu���e�[/7�l�^w2�,���{��gz�\뀙EE�zV���[t0b<ǂs�[��Dz�/x����Ly篧}=�O�^oL=�:����=���v�m�{�R~���o0F�]��F���m7Ć�q�Y��F�'
{��9v��P�v&�:���m�p*8Ń`�����/e̹��[�0e#{�32���9<������7*L��)�2�gD�Z��-���R�`��v'��6Ĺ��E�2'q�+4��c���ɶ����6|��?N7M�Jd�2ε��6��$���$"�q����u�OT̈�A9��宵��1;���ZX�W<-�8cS��p�oS��,jt]��-U�y>#�ހl(�5�U���Ί�j�y�
�ߵ��
Y��&����o.�q���1A�ߖa�]^lܔF��4ڢX�J��#��H��Z/��o�C����¡Y�˺[�_qX�U��\461c��d���=�6�23��%W#!�g10*�;B7pT�X�ܮ`p���F�p�j����M=����}wu|����n�'�v��N�v���n@���8h_+Wdg#�!�Qw5|k�"�d�	�*a5u��7����}He�$���P�ǿ`�!�6xѫ޵֌~J&�'��穖�����մ,e���QL�����9�{n�[����\���0�{��.x1y4M����g���F*�&m��x�p&�8RQ�}5+�3}�׆*O���u�<�=�XV�}�9*��LN�:pq�do+0粷_�7�K���9>f�S�s����g�9ކi%�_rڽ���.�Ѕ�Coy��_llه���u�x���c͍�\�&k�i�N��ݔ���x��$i#.ɏ\�:�PNƴ�$�VǸ���Ҡ(�?=�~��C�؉�o��,������^�`�3���W��e̩ؕD{P�s	���T��e)�Ҩ��uժ���!�G�O%��T�XT���-U�ͪC,ļY�i�{����U6�V>e_L�ԃ1f�����}��N�cIM���=�sk���7�Xf�R�VM�~���$�ൌ�z �Yf'���f,�3ٱ:�e���I�Ox�U.z�*��W�/O������;��$��2=
��\OxhD�;һ�`�OϱMa�V�_�S_`�u����cm![�m!�v#8��J��rԭ�s��=�SQ�c2�w��Q���4��<X˩�Bx:���*���X��3{���aI�: Fԩ��"��S���Z�.�u��T��2��/����q�[�\'Rn�����yI��X�D�z�8$@���<S��t_b��S�sz``�a�O>o{��Y61R���0v�6����rS�Ѐ�W�)#�d�N�l��]��y����--gnw=	�xb�M�����Q{��ABBݯj��4v#X�}I����Kėy��b�{�tO.�����9H��䧳=�fj�2ľ\%���xǖW2��q\�̵��4�L8Yw�ne^.n<�wo���B�Z:�f�ֳ���mmqӂ.��6sX��i�rf	H�3z"��R}�6%l�gu������ǉn�m���v,0�^&�CYk�;��F�������� �nY�u��{���T���q��M���s�(-��,q�R�m:i���\}���n����t�oqN5+,��q��I!���t�Ǡ��d�J��FXV���9�c
�3����w�R��HN�z99{y��F�U�e�X�; ���S�[|�ޕڥǁQ����:�AҢln����,*�iP�;Bڴ���;����>U+J�Ǭ�1Oy޷�M�4muoe�k�*�Y#P̾�tL,�A��x�D�9�����[6 峽���]�軭]��}m�Q��VT`�Ws]��ڽ�ȣ-=�.*�S0��n�{PV����;f��v2���R�>T��h��ǳz�%��z�bۿ�nej;\ɵ�X��d�ے ��A
��p��`����gIfmX5�:�V3׍L�v��e;�����IWR��s�M��Bc��=�74�	�&���.ݻ֖�r������|�0.��A L��]l�r|{���|�]�A�v9U�f��8��NHD�޹��$Q3����p_@���{|#�ԟ@F3i�ik��3H�����XL�'�^-��O*5�n'���k�S:�ԭ�Z֔V]��u.�R �[V�ad��?*�;�A-�Q�F�x΃�F;��c��ZP�#4Ve�:�����Q�}�ٙ�3p�|r@w�(�e�j֮���ӛyG�/E?�h�����A����GiS.+0H��q���:����3{�����~w϶���Y���Tb�E���0�+	���*���!�KAVd���(�"�I�R�R�Y��PeV8��I+V�J�f"�5�f�P���VTQm�PQՅ1�Ƌd�Ԃ��1��Ѩ7Y
�\-�Ա�bQXT�kЭVam�ZCd^�����+1&Z�E֔���Vc�4F�
���U*���J�W,* �I�0t�b��`���S0\��
�:���ӌQ@=L��ĭUce��kI]�-�^,�U��sl�9aj�����d��]�gv�u���Қv{0���'�F��L`�{9�S�A}78��M:�s�|v���o*l�����&�E���E¦�Z;{�Y�x����9槪�?B�<�C��ta����'��.A�5������;s���C���z�Wy��8����j�y7��:v'��6)rq��yՋ<���yE�#��z��5 ��z�����:����٭[X��;�$M*�W5��IQ�฀���=Gh�lS�T5��ݺ���y!���$�B���g�垺J.{V�{�.y�:�d^�֜��@g��u�c��z:ԑ�xK����s���c��k�Ӧ-4�WB�戞�\{��OT����G8�kpm��C�9�W�T(�V�2�l�S
���UtY(ർu8BB�+K��w]m�xy��_��5�ϫ)<��j���,j�����Įy4�at�i;�-�}�/��0,�'p�M�Ml����*.�����j��K�\�����b��������O�M��ŗ!Y�X�����:3zĂ����7���o��U�����GR�j�_��&1�n�΄Q� r�W���D���W�١�"��7wv��N��h�O��ם>ų���|��H���+3č����A�j���1��b*�]�o{!��,���1p���]֘{OA�7sy�8�\Ofr/s�ۮ���,��nX::H/��䠉9K N�Ν-6�R�ӡ�����˧�8�n�<�ps�\gs<�[�D�&�j_]&s5�CN���0���ڑ�%Й޷N��;P��N��)�<��h\}~��h.p�U��EoWc���RU6H�5o�]p�=����I��}��B�3bp+��xִ�n����6��KC�CH�����D@m-gx�ll�\&�S$[n�	�5Af�q��(��s�SZ�j9���zv:7�=9p�l�ᐛ��Ex�Ǿ�'�>�_�*hYR�yX�|�)a��և
T�w���&g_�+iV�}�R�$;,��L�ܗe�&Vh�r�7r38'�]�� ��������څW��r'�*Ⳬ�k&έ����9�J�Py��c�b�����E�z{g1�g���x���s��yu��;mw��{J��.=9 5�3N^:��5�����R����[���d������Q�$ ��5��Թ��5�E	�U�L��Hj5��ND؈퐜�t��#'��Mf]��=5�Iѵ�:�e��H1{�=ٕg+yPŷ+5.���e�}f��C]F���t}Bl�?_�ʜ��O�;8}�R^b��]���l9[�Hs%0��-��Bun��(�lᩣ7�.NPr�'t~��r�瑋
u�wۛ�u�� l_�͊z��I
��'έ�����w�̆(v�	�Z:�Vݔ�F ��U�e�5��~��i�1 R�m������N&�f��'TgN��a1=�e������?eQ�V�R�5�bs�S�fK����&�oe��6M�1+���¶3��_�P�6�[�Vs������yu[7]D���ři�1���1������_,{ܰ_d��Kv��+j��U+u���=��&�J�`&v{�J`����ø8H܆8j٧���S����ٗ���6
���᠍���u�D�}�d��Xܸ9>7�wKop$tb�/�XǍ�o��h�:F����1�{��v#�8��.�������p��j>���mP��2��c�7������]�8oݚ&��ɶ�W^8�f������J$4�"�Z�z���߉����{ˢ�F��m�hmƛ-ձ�� �1��P���ъ��Pk*5�R��𐌎�^�zA�g*�[����砖��j9��hС�M\t�D��iVC����GC�a3C�G]c�L���me1�����xL���V��l��ށ?Zr����}������J��v�:R�2���HVn1�V��`�x-'*��N����.��D�n���[ċ��YtН�5��B��.;֔J��絳]=BVG&�T�ܝz��Kkd�:��JvgG[��N=�0���p����N��n�n�=�^�iӮs]�j�`�����r~�Y�0&~���e�N�+�ע��[�9��U��^�\��~K}ԍ����ڔ��f�����B�O���/��>{x�،�W}���%Y�P���W�R��K8.���gv�NNI\�{����%�N�O:�y����w��4��dp�T�i=��׊�K+37���p�E�E��`��ݨ��)�7ȾiP,_M@��-=��b��I��\S�QS�$�i����@��Ү��=�!��7]z�>ߧu�>Pn�.���A+2�#�:2�*k�Z��`��I޸[$��b1*衴7�d�)�#앷&A&�NV}ڇC�of[�EU콄ʸ�MS��ސ��K���O�>J����Ĩr�b����>�v����W��&��F�_`��̻�4�5U����l�7��2�Z::L���J�&F��ĵ�)L��
bԭ�`�UF�1:����q����|�1m�C��/o�H|����K2��x?/r�Z);SK��P�"�QD�w7��l�#�����@r��ɬ�l8�U�Ƴ��_��9ݾ3�#427@�,�j����uC.6���4b��#x9��G�6��ڣ6�XX������\��d���-
w��DL���Q(^��3x�c����ac�q=z�%�w:�SkR�}��U-��=��ױ�j&㽩��`���w�'���q\��ŉ%���;�V���Պ�:`qMZ�T�R�m!�FK����[v��X���;-�[��9�|������[.4Sޡ!��e�#o\��:E���Q���vu��/}8bi\ɣ=��)q�*�ϝYt�������i���a���~׉���:�'i�vs�Gɯ,�v�-�N��V����ї>e�ԛv��m�֔I�˛6Um<�yؽ�����p��v@�U��}AT�u?Y���u��Ä2q�J�Y��ϏQ�x\�˼ۨ/��s�$C�rv��&���v��$��S2�,����b�WR%��M�Me@��F_*{��)`��.	:�8���nгC78�{nS�E���[l�:�ɠΝ8sG7!�p�����:���~�.^寋���bңN��Հ��#u��様����7+���γQ7��s�wש�n��L���ZƇI7�.�b�����z���)-����n�#֝�+�LFM�M��7Y��>���K5B�r\�[{��OK[����c��5o@+*y>��QW��5`���2���4(F z9��O#�ѻlpfox����$�,�\	<�ps�k"��S�mѢ8u�qR.u*v`D#z�z�
ڕ{�	K��݌1QV��`Π`�e�����g�<�h�v���wq�X͐���.7:�u�����KYO���q�f��a�ˬ��,#N��X�j�4ƫ��7��d��һ��Q�:��:��ع�X��Ď1���R���(��d��.�$��]��DNR*F�GX|���j����s!�^�!|�Ab�7Q��}�'��u��ue�r:Qn��ۢ���J
��V1A�Q^��ժkss ���͓�^�Sͨ3r���<�P+�N^���f]��1��TW!����)���AX�\���a,�Cf��N;2��;�ۉԼ�Q�l0z陊V/Y� A��0�\��p]qt:(s�HFn��T��f�룏��֬WjsB�UvM�oT������٢�ʳ��Z" E��Y{�D��N��7m��v�n#�,�X� �:�,a U�R�<t��M��׿l��B�Vl�*V����D<��Hm%�^�,鸜�À�t�֫oc�p]�������5�rF�Q�h�MP��s�fQ��|��QQ2�u0"F(h�}t�S1:1�R.�TF��*����j��)����Y�0s��t�4�&p{,�F�U��V�Z��;㵶�	�{ڬe�h��Vd}o�r�׀S�M�,�T�r��\b���m�Bj|�n����D��x6�e1Zy��P9)֣�}����@�T\�f����[���eN5o:��/K�7�=]�Ucz����Ws{ȼ�FѼ�V�FZ�|�E�Mi�u�+!�Y��R�ܭX��M}o�����*���$-�7Yߠ���.��$����Ci��������7�����+���ۧCU��Ԭ�������+h,X,���B��J�Z���k1��$*��dYQQB�4H�P�b�Jł����CHi��$t��kWC*Lr�
ԎJV���k!FDk�
�2T!�X��%`�Q��eKl��J��

VT4��ѹd�2�Jm�V-`*Ɍ�!Z�ģ�T��m�V"�*ԩZ�,(�E�� P�,
��TRVbbc�EX�%a����)��XB���燿i�����6ߵ�����o�s7�,��=�A�ò�
R��ٓ�.P=9��6q�Ż7�&����5	�#	�/��仾��؃�7���j�TuеJ��#�{�i$Di3����|VˡY-��9Nn�7cH�W�#M�i�ҚW�(�LU}f�4m�;��*ڹ�:��{V_���0�	�������y��<�I���@t�bxlN:[H�l7٭�ۋ|v�7L��ڡ�O�t�n��:˱F0:ךd�!�������������dG������nM>Y�LQ���{���K���#'F�DL)d�L.�HI��4.ms����O�A��a��gn_x�ȯ�P�v�]��Ǒ�u_��w��%�G�֩$G��Pf@�Q�<�u�eF��s��S��wV��f��6Q�M-�'@�&=���	.(N��pLn�>Ü���r�~�={^m����>�9s| U��]�����[X�&�8F�z�3cL�K)���ʡi'��!>�Um\��k\��������o�ȍyi����}7r�#4���*Vڧ3�۱�ό[����ͽ��d閦*�G5����hݱ�tn����ito5�w��.�o��؟wK��,��H{�	t�;#j������]�l�y'7{Vw�fU�z]��4��}&:�ٌ�������, �`����1!��7�+xM;D�]B�Q�\�VԵX���6���l���S�b֓����%\/.Fg�7�ʌ�Vb�g�n<S�B>�Z���)�+i%�<w==�ǀrx���\*!�K�����S׻��ω|yR�����y/=\�{�l�����S�,hDm�r�"�c'��ˬ�.��{��*�OG{k��!dRa^s(�2\�+�<=BI7�jr�}Q��5~�Υ��\R��+֋���i������dm�d�.��T��1d�[�|VG`�~�(�T�<&�����¹z6+�W��m̄�4�l���;�v��Ŋ��L�`�My��C�ǐ`W��g�,���pf������,��CkQL��Lv%���tsJ3�ĭ�lg7�n�{"�m��2�5�]�+ޖ93c��ĎJ�D����0���/�w�۲(�X�h��1Ƿf3�������;(�R����8l���a;�wLE�<��ETC�ú�:mY���x�AN]�2��?xҡc7�u"&�JK���y��WR}o}���C��y�T�v���>��C�
�g�h��L����Qa�����Z�Nw���Rn��J���V4�GAU^;�u�11�j���wAF6滿D���d�5��M�u�g;:�o�Q�1Ӝ��H��x*��+��z1]�2� ��&�YWLi�]�A�+z\����J�}ÑnE�e7J�vv�ݲ��ʧS6���)Q��v�O�q�6��u��vB��[��)��q\�����nO�6k�v�&B�nE�F#}����-+I���|Hݱ���d�T+Y�ۯu�=+G~N���Ăx`�z�̘�5��T��P�ҷ�B��X�B�O��w-9���n���9D�]&ևõ	�&\KT�D�x�Q͍�ȊeS�Ds�"xG+�����[�׃�hh��NS-��޽�{Q�^�}ך����Y
�\�w~�6��͞����sS{���Umt��0�`�R��i���y ��L����о���+�U�th�N���F9"�h�"�ں�3B6б�:�M�7���M��u��iƍB�2�u��Q7Вk�Q����`�ί���ݼ�B�P����G8���������$/��x��-:a�w/�� ����z���!e��^�dtwy�e��^n�ht��B7O�_Mɧ���ާz�*�)wuFN�$X�!�W�ꘇ�WS%�� 6�g�Mg'���4$��q�s5�����6M�i&�xW�}�ob��\�r���z��J�$|܂D�LO[]�Z��R!�x����6���D2Q�vg_s�9����w�{���Kt�=��L5xQw ���8;GVѡm��Sm����*���<�1ʭ�����u�P]
�Ʈ�u�u�h��T��ӽM����f$��I����8��Ś��K�͡�f$2�APHҨ�Mra�s/S��q�^�ʼ��ƫ�__���D�gf9rզ��ᾣ��ߚ7{\�.�B^�Y�1ɝ��!����z2�⮢�=�����t��VA�7YhS���jQ��:2nr��
�/*̫��+^v�S��YB=5cM��%�R�Vs��5.���/�9RH�@��O/<~�+�/�Z�/��j�{�,V�n���-q���N֠��2F��#a�G�a[�A��T�K���"&�5�v?x�ԛ��v�f�3ר��I$�\Ӟ�٢+�Ǩ��P�_:=wj��}�1Օ�1��v��8i�g" �Zպ�YRK��	���d�9[�r:�T������Qҹ�S����ȼ|[Og�ހ��NK��Ԛ�bە�n]hY1�*�v.l��/��F�,�.��T������gy�(EދuƆ�4��r�v^z�x�L��x��	n�h�T��R:��wo_"�!�7�O/��FR�K6(�΃���}Y�P4���N5kiV
�7�\��W���m�J-����v���	�5�,����ٕ�����(S�[udeb����u���i��r�w,F.� F&�<Y����p��q3{.�����03�y�tVm�㔠�ɴDtWoU��\�Q0�yIV�tf6&k�q����wCO��48ӱE��C	�",gf�E���C�Zma3���w(������rr���U�o��j�5�W�˾��<�'9*�WJ��!�6
�;�e����Oք�*OM��&��}�-�|�)��ks�B�F�BDb�\��H�� W�έl���3$������6
�vv�/��ݵn�B��"��`�
�%̒%Q�G���Vb������8��5o��T��Թ�����i�f�	l����Xy��T��iZ��ݩ�j*FT��5����U_K(;�14��*�9�$p�M#z�w�蚵�J�.8��i������zq,ט/z����5.׽��:��8#W���ڕq�[�dY�:\S�޹�1�g*-iȦ�����*�(���D�pR����i�]�S��璚��M�;Q"�X�vn��k_Lr{�Ǎ��뭛�3�X�����V�p!����L;�"ҳ�ΕYTc�5��ui�t(��dŕ���#�}������{���X��1VV��G�B�_&��}��/C|�Wgb}æ���޹6�V(�+Ql���z�6����u�_�����D�7e0�P�k.:{�@&`�"ū��+�bˣN�Ԏ�m��Ox~�Z�U�zxU�������v�>y8/�[$���۬U�1NZ��iİ9�U�һu��4��(&+a�9*n�~�5����٩��T�f
�S{�z�D��X�<���	AKq��u�ı4��5�|%�h)���,5�b��˱��H�FN�+��K>ㅮ6��*�t/3����]C@6;$U��ݢ,k�m�����	���������rwYA��D16�w�eY��E�بv� �y�k��KSK+l⫡ˋq)���[��4��N�S�q���a_��k&�Q'0f_}�T�˲s2��.Ɛ�����\�feL��F0����4OaYX�k��Ú�-٢4��q����j�gv7�tmؓ��t�z�l�s�Iɕ+T�Y����s�V��{���|P�Ӂ��adX��y˳;>x6̭�ľ�i�s-s�#��?vue����,I���b��X�5��Rx��y[��}�(��%�!{��i�CxZ"Vա#z�mQ�|�Y2l9VƠ�pQ!�	e��Jy1��}��S*�m�6��,����kr�f��oj�D����s���:�77{n�9���Y��9k@ov5(��0.�$CV��&�2f-K��P�z�������³O2�]8�KɁ��r����#n�bV�[�Z���>Cr�]��lu^�X#X�񻏝-��[����� WnLV�r��R�0ޱ|��o��mQ���F��;��|�3g!��m���B��V���oP�TT�i������w�6��� �z&L���<z[�܌�l�q!j�]VW%ںl�2����te��,�˹��U��&�J-tmgFxL�����B�@F���B{;cn-�͕n��g{�4���p�zMv__K����NkZ�Q)!^�񫯪���yl-�@������$1
�)Y ���.QVK[R�<��j��A bALe�
�*��+"�AH�`�@X
��P��E*B�Io�bH���T�t�
�Y(�JëLk�(�!Y�E� �QƂ��T#j����J��-)*�V"Ѭ11��HT�&�a��i"�����m�C���V�Y*TR�&#�E�Qլ�bB�M!�&�5�&21�"��>�2�:*z���z�j�n�3l�(^j] �]o8f8`�EI+1�ދܔ�%X��ӥ��vh��X�,l�bsQ�N�ƾ��Xa�>� 'MaUi+}0�@}��mqU��1C9=m�ҽ]��*rΦh��9�ht;J���V�iU���H�,�!��TH�T8@�蒕ݰ��a+���'�n�6{b*�pv"�	�wxywG�x^`�҇J��|w+ѫx��\Cٞ4�'�(��Pd��ϳ�ՙ[��5S������,cr%<$YJMF[�K�xm�zޝKa����+�-Gƕ���n�ޣ}e�t��Ð�+��Z��n���;bd��H���5{	D����k1Q���m깼1=��"�P��`v%�l��2��-��Bs͊(�G�k�^���}���g�1���*
��T~���·��(5�7��z�R�r5u���Y��U�˞v��f}G�]w}��G�W@��F`�E�Ĩ���P���үM�+�8bJ��D���ȴ�d�@ �p�zPmbڕ5k��uS�H�q���"L>� ��H���۩bqj�|�U���*��*�O�v��l��UV՘�V�zƎ�I���U1�*/.n�͊U6&��ȡ�O%�0t�H�*�B���f�|��x�&�~�<1�_'x��)�ͣ�q[k�kK#B);�b���ɼ%��3��l��c%��W��Y1�9�)s�|恭��K��(�ҧΥY���������ͻ��K�<��8x*�)�57�¨��);�&���8%UM�oE���[3�m
������b�'=cp�e�QOk:�Go<qu��G0<����w�4_E
��$��d�`�z�I��V�p�ݳ�t��2�C�1���t�۝��Yi;'�,峫L�Fʥ\͞׏�ˇ���b�~�J��h��3O��ǜ���1�t��q�+d9]t�CM�ʵ�j�4���2I�6hI�!ut
��S��)o3�𮘺/y�HRU�<G���vKMo�D�-\Ir0;���͑�J���VǺ��vA�("�qС�%������f�W*uۧe&��@�j�N3���u�f��ݜR�.�oPz�[�ē��&:�:5sV��ʦ$nЛ��O�"��(:���9X�:�k.�mX���U����Ü�{�،ҝV�&��nU[�!٘z/�\܃P�whh�5CD��R����VV��m�EU;N���Vr���]�%d�nS��egu���z�##��h��' �ǆg�/�i�u���ZDٕ��s�VSF"�b�N;=��$#\�|+pl�(|��]��ײO9! �^���.�E)e�v��1�%[84l�Ot`4n���=�Xޞ�������P��j�oI��gts�e�D���Y����q���7;;���4�u̓w8�yH��v�g�*7�˹T�t���Uh�;[0+�6~�[�^��=���6QY$�}{"t�j�%<:v�Z_�1��6��y����Wu5;Ŧ�T9졵б��mߐ�^eZ܃�s���<��F��f����	`m�\�Y������ņÓ���KHʴ�>��.�^[d�j�CH�/�L��6�r��8�9ٶ�3��,��t�3C�u�QWM�X��*R���N�Ϙ"��%�0q���1ny�����w2زV��;cJ�ٳ�a����������+�.�bG+�:�T���+��|�h�M}w��~���Ry��>�i�����r�%$=�ĩ��ޫ}���o���+(�h)$�C�ι�rǻÎO4k��p�ά��dc}��A�X�-Ǿ��
�y犏�<��y9:��v�Gp�M�F�o�咦�,S�����|��^��]��^�n�J��JD�I������T��B�~#�U�5��<@���ϒ}~�~��� g^�:;(�m���vpWu]6v�>�U���{z: -�����s�7�ZT�,�y��s����7���x����ˋ}�!����b����^Oғ�K)Q˧K�Ϯ���Hͻ�����[���Yn�g�܃Y=��/���y]
��3]�nr��k���R�3�s��Xە�w&��}�l �4�1S!ġ���Ol貮9]�8U�e�b���=���nk�UXvc�5
V�����g8�i,���D�\�M��F��j���:'(.Q�%ޒ\r�\��y4ګǲE�0�n{�o�ї�l耮ɗT��<�{G�{��5�w�K/itOTo`f�M��#$'s�������^�.a[U}F��=|*c
X)�i�cyvsKL� Ӽ[x��o��x%*���?,������D�Lj+�6�0�a/�2R�y��^�İ��9���}Jƙ�:/�8{)*����.;|M1��w-8��6u��lf�ʉLiZ!j�=��t���Px��C�+2*���Aq?b1�{m�6��9>�q]&Du�-WqIfs��ck�Ѻ}@|M�C�5�u��u�Z�"�9��י$X6}%e��X�N}슈��z��9���
I|��;Y��/|V�>a� �u�s���oH��|�@��׹�Y�K�猪��O=u-�3��ʭ�t�'�̹g s�\턕��B�;2��km�!]$��u���>󹉈�-��o�qJ�5Ӻ�tv���	�r��dF�U9�m�I����Ϊг�Swq�;��T�o7��.��Sg�v�n��s�If�{��i7��G&�p�N����:�ġ�ge�����)������s�5$�k�b.�z�
�Epz�z�B<����)�j���i>ewV�0�r�b�>l*�u [���	o0%
*j�g�Ό���s�[v�*��m�ݭbݼ=�+������y���9�a�����B�m�	�	����g�k�	�-D��v����xM��Y�l�rKjn�[�8=�"Q��f���k�.��������}�g��л��|:��\��0y��9��)[��{k�32p�L�����<iS������m�Q!�r�Z/%��7jrZ����wX�JO���ș:�<��w�B�v�od��t���t��S�?LC"0M��vkX��RЪ��Wh;�0�V��yơù��؋x]ﻔ1��T�F*�ģ��펬�k��CYYG�k[ZvW	��t�G�����
_A���}�C��V��[m����&]*h7��d���8�M�%GX�SV��BA��e�'���m��2C�٥�<'c���e�2��斣��9{�S=�v$�+��0ܖzr�U�sP�V�\�_�AV�.��ɷ�*ŗ��Z3���f�����#B�Zk(υ��4)lٗc� '�y5�I�>]5��U�p�5Y������C�c��J�r/��D��T�Q������8�f�n%�rʷ�+�V���,leLk/�<�����I))$�G�%DQ
�=��(���
`�(���F$#��,h��g���
{���h�z']��O�icX�
V�-[�YT-Q �,,�/t(�|H_�C���g�f����\(�҉�;�X�"�xdٍ�m�S�xm�P{�����3}
�p�6 U�$kb�E��>fdP1�*�QS�JN����<�P09�::�h<�E����<u��r\�� �qW��!�8����A$J-N����	��q�'���=.P�k�e�C��=�a��(r�D2���}*�a���T1i��s�R	��?y�4P�4>����J~��R��pV7�����q��.u{�a�Z����@QBK�tbz��԰R{+�U�(�!?S��I��V�D�
�M�\�=0*&��P���X(�!�pSH�85��ki�{�.��#>��9��h}P8;���Y_�=�3�V�����������ƀ
(����
��=�l09!����J�
�m7Ш�����aN�|�:�^L�M�u?���� �֯G ��<�M�5Ch��c2������t�ɻ�T�>�(��ג#J	m����aW�E�C��B����9�PNFٞ�k��y�ȸP�]_106UEE�0uaD�A�Rn��>&C��PTB�����0[���+��
�R �x����U��zk�7/r�MY1�}��DQڇi��;�8)�DE�	�;�1�h�LOC��?xk4�k� ��m�T��Yj��T T��Bz�c�8��� ��7)oφ��-��DQ������z�'��E^~�2I�D(��;Y�S���a�5����P����N�tC Ȏ*ƩgK@����̈́��+��=p0N�hG��z����2�b9���;]�QD0����%�<RT6S��"��mݛ��z�n#���^�q,�ڗD����E����|ƠoC(q�o��˨�E�<N�ܑ0��:��87�0h.LB���T:V�0bH�P���9�5������w$S�	XJ�p