BZh91AY&SY�3KYۗ߀@qg���#� ����bM~��        ��J	P
RR�$�B��*�
R�"�U$Q"����D���Q)�b������T( ���%��SkJm6�1�4X[lj�[f��+l,4�i�[a+L*���j����Jk&���m�)UEm�FkE+Z�66��  ]�-��ZeM��	�$ ���im��6��RZm��-��lbSmFڢ�kUk�	J��&�"!��H6ȪU�(����kClV��  A*;��@5��������Wk[vU m���ֵF�Rt w`��p�&���U=LZȦqܪ .��e����S
�@�  �����t�9�[��V�������o ��[m^�����闻�㽞��m���^{�l�ʹ���+�斍RT.w��+X���}�O��1}]���|�Ɗ�S[}��Z��Z`��kR�fT|   -��}�V��Tk�{��������{��ʔ�m۾���w@h=���_T���o��R���o�}W��ڪOs���4�մ��\��ka�u��ݔ�*7���JJi��5lm�ųM�  _|]��֫n}w�})]�v��þ�^}
}5�kY��<�����]^�^����u|���}V��}�o�7̃��9^���{3Z��|��Е>�%}���[a����`Ъ�!AkEfj����  �^}*J�����}��R�Zm�w����ݮ�s��yR�������}}�ij�w����}2��i�����[��]��n��kJ����z�m*U*o�O��}`��n}lU*A�2���ͩ5��m_   �{��V�kwK��w��v֚��y�^ʻeٗm7��7�J^�Z^+�vh�!�=w��4wt�=�V���]2�xg[چ�IWz���Y��]k���֤v�mNz����4e5��*�5�  Z��_Z �o/<��j������iT�1ӐR��n��kZ^���)V�n��dV�*Om@{{�P�y�`=P($U��4i���  ��ʕP9ܸ�>�T��j������mBю�w^�R������UD�z�p�h�W�b��Gg�;���;��`��E�l-�@l*�Tf   �g�}��z�z�����ES�y��/A���ǧ�k�۽�P7��/l\�k�������P�]�n��U�:�{lf�ڳbPZ��_   �5UUM���v5J�����5���vԡw���J+5w@�Ǩ��hw��P���s� �˺�R�     �   ��2�*Q�0�0���`O1%JT`20�0	�L@
������200�  M�0���IET�4  � �� ������  h4  �F�I�Ě��ފ=M�z��e4�D�����D�0H�?�������*�v��h�ˍ�Κs�wiY[v|0u��;�� {����PVAS� ���+�G�������?�x����O������j���TW���>�O��$�!PU��?������O����S09��e3)�L��fS0��̦a3�L�f2��&d�3)��f2���&d3!�L�fC0L���&e3)��f0���&e3���f2���&e3 f30�̆a3)�L��2���&e3�&G2��̦`s�\��S2��0L&a3	�L��S2��̦a3)�	��f0���e3)�L�fS09��Lds�L�fG29��.`�s���S09�0��M���̎ds#�L�f6a&2�̦e3)�L��4��G09��&e3)�L��G0��d̎e3#�L��S2���a3L&e3)�L��S29�̎`s�\ɘ`s	�L�fS0��̦e3	��f30��a3)��fC0�̆a3.fĕd3��f2�0��3��a3��f2�̦dg8L��C0��̦ds)�L�f�L�fS2��̎e3�L09�̎e3���W2�\ّ̮`��G0��3	0�3(fW0��3#�ØI��.as fW29��.`3��29��.as+�\�2��̮`��̆d���2���.es2fG0��̎as�\�ds+�\��2�es	0f0��3+�0es#��L��0��̎as#��0���!�2esL.i�3"fW2�`ȹ�̂��G0"�\£�Qs"�s*.ed�"��0 �\�f\�#�se��(�\�+�Asd� 9�S2� �+�s
�eP�C0�f©�3*&dT̨��S0�fL�	�E3 �aD�"��3�)�3 &`T�
��0�f �)�Q3&`����Ds�aQ̪��0��QȀf���Ts .es*���s*���f\ȣ�Qs��g2��̦`s���29��!�\��2d��́��0���.as+�29�̎`f��G0as+�L�� �.dsfP�����09�̎e3)�L�fS2��a�`s��f2��̦`s��2f��?�Mz�����a�ZO��
	���!Ӌo����O�� ��������M�Pz�G$�6�V����52Y�%�$)Pg�ot��Ch���f�QcI
F�2
�@֭W��?:�~{���.��B�tTq�b�v�c� x�ߖ׭�b�ͷ,�򢽉$}���o�ӇJ�a�)���oV�γ���z�d�7TQ��fi֬��r��n��N�e�r��i�2-�ִ�L����Y[YiL�4��wg0B(m����5�r�f�DrL�,h�C5�fh���6�d��HB�]EI5d��<����dAh��Ū3�mUn0�]ȓ̘<-ܹ�<Ƕ�������ua�c�Rdy<7�Q-&M�jT�F܋�r�-�a�4�h�"غ�e���q�%��l���H(�7n,���2��h�IB��.y݉����iE��9�V ���DƵ�o+�c ��YlJ�%��4\	h8�Ř�q�P+"�9פś��6�JR�(��T�;��EV5���&k;�M/|�"{Um��#�x�����b��O�6����[����
�h�&���d�R�`������-��X�o�{�<����+�V������ŀ�����TY4��/�r�X�w|<V$N��卥R�A5��x|==�ň]�^yg�&�Z�.�)!$�����T�3&�M�T� i�$�T"/)��G2XS[�4�8��Nj{�eh�j>َ���}��=z}���W��p����R����;�ۛz��o���X�in5�Z����L�;JQ5���Y����nGMY×I�$�.ƃ�2����P�ݶm�=� �U�g�2���=��!P�v��f�2n�d��Gab����\zֹǋA�.n�e3B�L� �N��(r$[��4s��Y�gnLM���[�F�L\�wLH�3��蒧�ſ��Q`�jDnɋc}K�o��������k����o��Z�T�����k.{ua�ЧN�
�Ƅx<���kw6��L"2�\�yݞ�4�'�)�,ՙW�����/R��V<M�܂�"@ʭj�^޽R�PnO�bZ�6�����Smʹz3!f���z�À�1�֓47.�kXԻ��l6᳚&Ӽn���qAz��N�,knM��,5&�긋ڔtŪ��d`O}�^�&�������~�5-����Yr���f��o ɋ`��+�b���p���'6�Z$C.�*�*��8�F��w�^>�����"3=��[cZ�`��nۑ0���+Z����q�ڛYO&�NZB(t��Ք��{Y�V�ۘf�R�-� Fs��I�����D����T��mʼS���?DƼt��a�hA�[�0�z�z����+��,�OQ�%��^{|��b���Ai��WK�<�k0b��:�p��[�9Xʬ9b@ӪaÀ��-�6�_9o�v�֡��/�dSU���-IMf��@��^K3tI�b{��e[zsl��U�Y�ۀ���8/�!Eɪḿ��A렁�[p���6�T��L�
��lm�襯
l"S�����r��/ajx��on�5�#���]8�'���Z����K5 ���<*���QëI�nK���5;�f���3�o�=��s3;0��^5`����z�jI箯LE�2y1�����r\~$8	:ڀy����8�@�p�n-ʡNĸ�ة��a
�Q��H]�J���)S�I��#K�d0j�h9 ���Q�v(�U����wZF�q�������'��(��v1�A-�<�b"<�d�<���r���-�W���e*���A�b�4�Z�ҒIsW��wn@�wb+ �'�n����L-�#6/o��';�����_X|Z��g��R��}1S�l5L�$@:��w/���(ڨeb��SQV-��8�1��ݮ?_ ��6�*{=8C�n��K�XB\.��ah{wԗ�V�Ai�z}��W�<v;f=�oo&<1��u,���OA�4�A�q�v�6+4�X��+ݬע�Y��_����)DbeOC2/5�5M�n*��=���bڝ�C�d����x��_7���$�)�Q	W�훏D>Oi�ww:%�n`#y7�+��+jLifֵ1#��n,�N���F\;���Y���CZ#��u�)e��ѥ�9|Tl�|��T[��L�#��s٩���z�\N�u��WA�A��+M!G�e'�t�<��]	�i�׭0D��(K6� ?��>߷4Ь>p�s�(��v	��%yx��mep�{Z���䎕�!4�h��w
c.�4MK��`�{p�nm�ǶL�����`�,X������4�7&���C|���T56v�X-���C�P��7,����6E��|/��n�ޛ��%i�
�����<�R$D+aڷ��|�{�/)��l�E55� ���K���wRᑻ� ��E��af�B(����R���OKbG�F)��*Q���ygд:Ϛ��%	^YR���B��nj�EdZ�i�jw����BJӂj/6�ו�`��]Ȏ�jԇ��>8�1i�:��195f�Eg�I۰�Sj2[��;%B�pW���Hp��w#r��j+V�W4��o�ͻ�
�O&	+D�Fjf��Ff5�h$��K��#[PZc%�~/8D���ny���O��v|��Y̴\�2CE�L+)y|st�M�s�S��ў�fL>�t��+���A�y��r�f<B#�C^�m�-꽭��u[)�[=p��3!X����љ2�[**|m@z0z=�ٛ@�m�|O���h��k7f��	2������ق�-کq��6lժ��~YZ�<�������Dm�Y�F�_m/�7��sUU�SM)�tT�4(/-����T`�5f!\��5�}�op�:�C�J
���/��	Kn<���Ͷ�)�d�EL��$��2�
2�����>�5�۪�n����^=Y���J��X�iBQ���X*mXʤ��2�1��m�9�S8/C;L������(ա����bg_ȁ��"En}=7hѪ�ϴ��Rn�3*��)�9�]�����ɮ�o��(BXv�b��'�٦�=ǁMX]� g�j�k�\����q��!AN,�-f��>x��B�(�S�� �������W�&�4�vd���'�2,8ײ�}����/��5^K��)�L��� ���|�B���{������5}[���]���aӺ�Y���Y���U(�p��Io*�I���^,b�?�6<�^�`�E����X��`��neЖʯk�׳Nlmq��Z�
��R�Vt��vx)�$��S�&eO|�J��trB����bA���5��aY^�^h�b+q!`��T^ѿVae�.��� ���N{`�i&��hc��ܸ��٢\n��tV"�tnD<=����/�g%����D=�Um`��!&�[k	ђ�;o��<Fd�K�Îyb'��0���.��Bw��aن芋`L{ۃng�=t���E�A���{���B�VH�H��/�IK�ü�P�e/%Xŋ���yxS�d&ܼ�1S��������Peww\	x$���&)�E�@�i�d���$]�ۨ?g�or�r�����ǔ���j��d�{�B�Lk�7�b<g͌�Y$��cd���Vb�E�z���l�՘n��#0
���Wӣg��l�P�T������$`�4"��V�j�6��RP�ݱB)5]`�+X5��8#���C�KiBҞ���:w5i//�#t��uYt��X�ՉT��5SK�7���BԴk	�f����v��Y���Fk%;���"�ZX�����=1iX�5���@����p!�kh57��͚�]�!�N�U�&�⺗Z�X�EE 5k���"UOv2�/V��,;�JS���^�ׇ	�S3s���۸�ݶ;ᐍ�w�Bȕ�ԶRTkK6),^�>���#�Ju\G��3h����[�~�h�N긞�T���6�
�ĨF�%mS�K��M��n́�u�[��-;ݹ���v��p˔	�P��#]Le ��Mb�lX��+[�	�|�����"L���c�R��bi�ʚ��*�Yt-&�j�y�Ig[$�<��V��7qS�^�/[j�^Sm���@�S5�B���Pi�[����������e51���X��f�ο���V�2��Ow��f������n͓w��r"���ɾ~�!�,H�۷n�גO��s��G��ֆ������h��wC����5�9Z�E:
�����Dɬe�~xő���<����q��q�4���#N��[�e�0�ן��{^E�$30<�Fм��%j��k7�:!i@Š)�&ҴY��H� �{wj��瓠�Uy�Vk��v	���e_]	ǾPlt
Ne��|���f�2T��W���sCIY���uC�g�P����.��Ph�B�E�C��_<���q�� �ѹ3)���Vbv���+Vº���7J�����0h���&�g�����'�3sDwE5yy���<rO0}�X%rX��Vav��(2c�IǗ�06(�bv�Kՙ�ž4�����RF-�̩�d�E;��3v�>Ն��M����A���ܣC$����÷KE-9V�A>r�c^1_�&qչ��H���l�20�]+ekA ]fUp���Rl�"����sM���7ln����2�#wq�ո�U��f����3i�|A�m!���ư8/��9�@�C3}�{�`Nbc|�i=j��p��H��׌G����f���d,��ڛM�.ne��&hG����J��5�F4,~l}5
h���]:� ��
���[�P^Ɲ'k43�h�b��"������7�����c�K$N��M�$�A��y�0le�me��]��BsL�a�����Nbېa���V���b�j��i��Tn�Ǆ:B!u�l��j����V�Ub���YWp&�S�]�3o��g��,y��6�zM�o�x	��qţۮ�t�ձPNY�!�P��H��R��uq�*�Yp#,��F��CB�7`�1+�:IJŪdIfmZ��oڣ��?I��a��*ǐKMoM)j6�9�l�k9�Zz+����2�+�=�k?nS�b�������^Z��[6Y8��	izn�l��n�(��B��{X+�=�����B���fqF.�'ټ��+*��Wi�����4&7َ�1P:�ĝ�n�]�O��<�0y!E�Zv}�r�T��)z�,A����t]�J�ލ�֛5w3T2a"/AmQef�����DY�0a�*�����s3�)Љ��d��0Vҥy��X��lzS�3���U�j@�籿Yu��9Ny(�(�7I n�M��ɚ�^���ǳ�����P3r�E�˓t��l�*nP"�Qzu�t^�ZY����S$���xO@�}�1�}���
��Zyeپ<��̉���4�y4�k.U'�݋�9(c�'�B�ᙵA��]�OCb�솵�I�=)��߲!r�ڦ{-v�v�.K�p��
t�WXdJԤ'%ƫ��V�
۱^/^m�T���{x�k����@��Ɋ=���� ��;<��Qk� ��}"g$☏�<�Oc5n�x��
���v.� �aTі`3+��^{5ID�cɕ�E�+j�s=��H'�Ek�ю���`y�_��p�}�f]�9v曵��*����uY��Uz�,8�	߂i���~n��tm;�Ura�2�WP�}~тOo�Y�pƤUn����BkM��b�H�X�j��I�Vb-�{b:CtŊ=�սQ��Mw�K^�,x�y_:�kW=�Ī7�b��f:E��n�������0�����>�V�L�p���U��FÇ�I�hSf���lx��Ǧ,V@tz�י<겄ݢ���������;��{t�#�ݛ����V�%���)����%CBor��V3�����&�>~ͻ7_���5��%Lr�H��Vu����&MYB�tJ	�B>h.3��K۷Fl���
��ãfn{�[�,z}1�R;��Й�u"QBk�<[�w�?�{�4��lRH���YVn�tA��e�>Ju	A������!�H�Npħ��������c����Z�sHB^O�{���&��$���3%� ��PW�����^E��y<��;q[XWh�3�\|(\nH�}�IY�y��`fz��"Wv�3g[��B�xI6�XʗܩttO.v��^�ޏ��y��_Yg�����$<�<��ʆz%�ݶW�Eu�׳�{;�%`g� rWƞ�!�ۥ����3ԃ��'o���T�r��S~O۞p?dP!��+e�)J�5㉒����#ʎ�=I)�B,�-����f��(IIOmB�����ҵbH+'��<��j`�Wx�`��%�V�m��z�h���`6�aa�l���[;������z�j�v���==��)U�F�����ӻ�dw���`G\��/,�z�V�o�Zyk���8�ꕌ5sv�a���C"NzF�sH8�un�V$A�3˺�/$���0j�gc˪�ɒ0�R�+Lt�iģV'��jr8��9�89�K�z���:C�^� s��Gt~�0�����nZP��YAA 4 �� C=���}����=��feң�~�-, ڵ�i���%K~J"��6�r�ɕڒD�_#F�P��ۮ�&NW����.�j\/� @`�y�z�Gp_n��t>p� "���&Dm0v��N:YI�I6��K�G�����W��V?=���ߛ���_����x`ߣ��{����m��m��m��I�jrԸ�G�c+El"����S��K��b�[,+e��w7,iꜢ��X��փN�	�mf1xͱ 2�����X��-��JA^�S�W]��fg{��1��i��&o=�ګ�<u����&�.��go�{;�qaF��Z�><�<2��ؼ���o�Cjk0A5
[W��nDD������K7aY�r$	�6��N
{�L����[�KҶ��"=l��7Θ6[��`�8[C
���mù���j-�;;�1�u�[��h��I��GٹuՍ�$�W:�R�4������T��͈��Z	��X��X`ȷbFe)	H|t��F�̦`�f��b÷�Y�T��r�G{�M;Ĩrk;]	�^��u�h�����<��vw�W��j?�ri"����ƃ�*�)"V����$l�{ ���t3�R���H2��̋�D��l�.��1��>��έñ�^6����=-��1�g%�I��1L�7������[.��grA�k���Bkqo<[쬺d���C����3rPϰ�~�;Oe�v5ڽm]'1��4f�d��+�x߻<0��L��j�IW�M34���p�&S��9ןZ�a�-�q�N:e6�Ff�uШ�rs�*�r�V$�L�!PnD�U}jz�S��3�W>[n.>��
0x!��a�����ߦF����Lt:�QW�k�7u��ې�q:в5{3i����lX�Ɩ����u]Ct���ں�n{��v�51>2��).����Wd�z��[��� �]a��[��1��LV���QZ֌5���-gv��A�{���~v �R&*��"��������r��j�h���g���j/���;���a¼�uq�ԋ�r��;<G���}�̞`8�"ҟ���Qi�l�f0򣚄�߮���d�РH�,b��j�l�]Wz�8�T/�#�K�#��w7v��,R[Jd���*#��#�t�H�t�R\+��xί�(�˕Q����|���Z�C�z�|#�q�;�ݴ�~�Q��X�[�Ǘl3h�#<�w�7�3^�U�%�Ow�ok%�$v{�{	BGtA�c\.fn&ta��H���/�+~��;0�����c�ON����|�{��g{[/ľ����/R��̛ӻ�31�G��8�Q�&��T�"u���N1i��8]�df�.��	i��)����.�5n�o ���\��ؒ#4oP��[�j,�U�*�*��N',]��qT}��!K3�s+�Iޒ�����,-Vs*�L}���n���
6ܤ�
��.¸���6���R�!�^��C�W�o,��;=�΋7t�˧�"��B������6i�Ե�R�fC�.�
0�V@0��sE�nV��Fb�x�\�PC����ܦs[.:w6�w=�zN�0��ﶀ�܇eQ�������Hz�]\yY�ЬfiT���}}�B1�_t+���}a��0v4�wJ�d=���5{p�H��.&X�cU����ݶ��bV��Sǜ
��c$��~v#��`��Far �wi��P�:_�>i��ю���f��^eZŵ�50�$���J�Ҧ�)pva3� <*a]s�/�>�I�R�rn�f����g'�aקY���Y���Ӳ�7I�,���]FD� �V��:�����yi����P��龤�����{��&f�&��h���Y
����I�AS	U��K��k,�f�Πs���l�b�:8`�����$Zً*�d���6Tm�t�%�R��b�����9�u�Y�S�O������&��0�L�]��Ls�tgr����.���FY�iJ��8�mTȁn�mQ�F�g�p��u�����$H��kCwӮg��÷;�#����|ཧq��o��:����'�oaQ��_�ل 3ANJ ��^��,wH����Nb#��a3$���Y���o)Q�f���5��ƽ��0��M+S�U��t5����!o�J7��wi������6����x��/׮����}/u���X�*{�i\�i�Z�JxD/���{�IY��Y1��Bm�1h�����i�1��j��d-���ϖ����E�|��_7q�J}��o6��%<�կ�4Ƞ�"�a�c�����738E�D�R� ,ؠ���[!P3�|�A�B�:�kC��3��F)ir�8)�D]0�3��19���ޜjě}��1l�d�e���a[܇�p�p�����屰'`�;md�%�1(�f�"�ý̒M-H�+@���������ޯ���f�c3�8��ӥnmK����g z�r�Z(%e]��ru��S�F4K���=c��xf`Y������E���)_%�ž�\�c)��w\v'��v6�vΝ��2�g�d=BX0w�q�wK5*z�C�|=���L��Y����-�\|e�e���%��"=�]�A�Pv����]�4��7�ػM��<�ȭognfv�i������X����d���u�M����"=g�1�F�y4��Wy׾����$�k�v��l��U@�+�������Z}�Χ>#T[D{u���"�V�.�� ��${:)C�Xp�<���\�=U�"C��2��j���E�p�g{#�H3��=�9�(��z�d�`�A�q2E�Cө�7���^r�'j՞g��^�岱��zM^���Թ�2-o(���)�nݣ�ᛁ��O:���x�*����5��#����awc8��۾��E�&�[�,qt�'��ڬĮ&O1`��]$��O�:My&��R�F��9�&�ǕS�20�#��qc6o�t+��Iܺ�O�*�R[��%Rk]Y2�����`؎�V��C��R���Rb���@7�#��lz��#I�wGX�>�.��}���W��I������,���n1�;��,Y�*��E:���2�(,���ɳ&��&�[̱�4�͗;o����.��d3^̵�F=�7Tݍq8!�y�m��nwO�P���D ]��X���+9��\�Nk���Vr��w_�?f%�2vX����5�o|�4�,�L��n�ܥn|��r�D��`5�/�����ve�T7��_b3,�7>�7_n��9�?X���Dʔ~�{}�H�ssvZ5��@�>n����C8���1��u�gMZ=���E��� *;B0^�C&5j���µ���i�e�MUk���Z�̳Ŵ�"3xe��@a87 g��։bSkgVs�>7�Β󡛜L���oniV�Xcm�8�����R�˂�����6�4��$�<��Rh�q��C]o��~�j�O�j�{G���Z�v��k��l5ٖE���#�pfyfK�L�%:����Ћ�E�<tm��i��i:]���5m�v�����P�y�i�>��n�;
�It�'|]��D=�3��,o]-���dɼ��� 9[
ؙr��&�3�j���P��efFqlm�-�Ǭ[�`ܚ�F�Z���6��&�g$le�+1�U`���\1"�)mn�`�sǂ반�}��u�oS'��5�5^�D���d3��\W�5d��ۋ�P�c-]]�����8:����Mmm�9�b[u0�Y�ro�-1�t4��+Z�H��:�OcΟ?Q�2.����r%ڌVg]���Z��Z�Dwn::��<����x@�	�����&ы
ʷs�%"�v��w�ٯ2A�ِ�K����zw��-��3�*E�Z�=��dC-����Jp;�eZo�ĩɣ�P���&Rn&7W�9�xvI���l�g`��;<�b��bG�"�[���9�t��M����1Q�������Ҽ��˂�O����ccnN�]'�mD�:7Mb��܎�ʸsQ-���N�f4���xx�	l���F�'��΃UI�mUں��Q��&,��wpe�;�W�Xc��wۯ� ������.�'�,ں��.��w�/v��׷��)��[F8F��m,sٙ�ݾA��ذ���V'+����v���s�f��:�c��-|RJ�;�SV`���`nzA���:��\>}�K,�Q��wEr��^C�t�Hi�NM���p���9� ����5d�N>%�oh��N�|C�c�DxA�9�����8NP�����)��������t��-��}���;,�wr��{��=�;�b'{;���\<��?�GEug�2oHُ�q�{�0�Y��9��I�	�!�5bj�7�=[�D5+�y� �5E�y��"�&@�K$�L�@�v��0��,/��x�[ؓ�r�z�����D��:�f��!�H36�������S�N@�������ܟh���i�WE��ɠ���������,��[݉rC��Vx��/n��ӆ�:�K[�6m9q�$>��9gX��T�4�ʧ�|8U`�r��Wj��n�k��^�+$Ҍ�/�Xf'��j5����� �:�f=#a˱��
�h��Xʙ��Wq��0qd�P�ݛ�bf��(��.Q�Fa�˶Y�)���yײ���ԙ���c���@^Ψ(_T����O6��=��'�.�����k~��w��`gZ�t�����tw=�GnQ�w'h#y����Y���i����<=7��j{Nd��U���Y�B��,�Y�G^�U��wMp��L��>���e��Xs�Л�����l�A3B�ou2�G]��K7���]��~9��z�L����\o�UCU��;F��C4�p� ���E Jty���o��{n:hv�-�lMkEOk%�H�l�z�\؞y*���E����ĉ�{h��(���7�9Q|��{i:w��2�dNCv�O��}���\	�7�*�79\��W���f��k��7�N1��F��|0��7�=���%�-�{5����缒�L;�v���y{c�����~-�&���W%o���Y�5�[���<�J�\b�J��.�H�I��%����|�n�l^��	���,�Q��Kձ�\u��=b���CA�;ʵ��ƴ���J�Ȋ��������s�w�!� T�l1�go���"W���=���|r�R�<`�
�����l�����6"k.������:�5ah�=�X��]d �B�S�VӤ\�[�d�A;Un�w��r��7w��I�v�J�4�˔��{�x�^��}�'yqΚ{b�b5;��({��l�.x.��rt����$M��K�g��m�Gu�S[��owJ�R���t9�nBtAr����h�n%�(m�[�%Y�0�0 �;Y�%���.�%��1���/t�M�k-�cǊ,�L�`;0�w�kk'C�.���ՠ2xh8*��L�S��#�e X߅%�����ӆ�>ˊ88\�KƎTu�m���Y�A�{�>�o�a��E����D9�{��T�(��������,�"�Y��k�5�V�Y�I�+�:���X�7�\5y�y"m��`�{,�L����3Գؽ�f�Z�Ayi��%�j�*'��jkq�0���6�?1w�%�e��ƿ`�J�uԽ.�������4m8\\-��n|�]4RH�QZ�]��ġ�8!%7��,ا�7`�Z�9瘽ېM�ۈ��r��9��
�R�rV�)ܗ��!�A�Z���i���M�No�p�O&b�5Y�T�q`�j(Sv��N���J�w�A�[6z��
W/����C� t�m=��L��/�ga�Ĕ��G5���ސ��3��d���8_)Ж�����1�)�A�Q��+��Қv�DI]K�v���p��q�;k�N�6�\j6c0��UD�2#۲�]t��s�;V�)4@ތ8c(RY���v�eim���qt�����*�C�Ļ^�����)�xծ �����o/l�Egh�9U����%�s���H:���H�}��{��������R!�z�7`�x^(rd��ě�7ËOԉ�#�gM�q��+�-,�Ӹ�u�o����P�i"�٩M&��=�i��Q�fŒ���v������a��ۻ���CKһR���1
 ̤
���"��Y�[�����c��;��<�c�e�q��s_aVm��6����B]|�8�I0�k#Z=���w:w���Y��N\n��&��2���6ِI�739J�`�ŭ�ќ����2�}��������Y֙"�h�Đ�_��}J�mx8�*Im�f��"�a�3� -ESȔBI�B��Be��h��QHR���>
�S@��B�
$��T���D�	W0�4���b[��	�v�BBm0BE� L>h(}[���n�4�kri����P%/PtQHIƀԨSAڀ�QL�P����J�D�E�	d@B�C�du2�AR)Ah0Ujp��H�A�R�P
Ir��VR O�F�Qb(I�^M/!�V}��,�0�B)."("��%�O�
DS�)�@���T���fr�z�E
���A��F0���@XJ]\�$���*°\a��A)%�4�	H�Q���T%⨑�Bb�H�L�@�)@J��UQI-^d҉!^�P!J��e�� "?C�l��� K��Fcp�26������M�u\���j�7���E��������!�~~���������?�����(������������?��|���NY�O&��������T%s�0�Y����<��z/�<Lb*̹�h	3R���@�t�LTT��C4-��F�o�7��-�)oLWy��,�tΕ�T��
њ���J��Va�q�>��fR�q��`�4!�(��$a*�	Fqt�'U�
�[�e�sF�P��OZ��K����nZZW�{Rж[�:�i�����D9�����.M�_8��:@C���ٚ��Ok�B#쨥��h��_���5}�!3E-9�a�4r�Pm��2�#rn-ۘk���K�ƍ�x}�D�����y��w�vg;�sbE�8���;,l����[��6Q�q�@��?F59����d~�����6�Y�����( m�-���\=��m��/��U��v;��H�G;-cv��Oi�0�vo,�b����FI�Y6���o:H���5,��^;�`�6��w�lʄf�FnֻA�p���;ݩ1���}�sx����{1y��.H"w6_%gzR��io�/o�1�X��f֯W6)V.�e��tay�_t8/o��ϸ��v�vV��`TUn���$��ɸx�ـ�WKN:t����T�*�]5�VM��TVjݵm-0#1#��ڐ���n/�����B^�I��sD.��	�غ����+Ң�}C���BйYi�߮eU��4;�^ ][��`@������ǟY�s������^�z����ׯ^=z��ׯ�ׯ^�z��ׯ_��^�x��ׯ^�O^�z���ׯ^��z����ׯ_��_��Y�ׯ^�z�����=z��ׯ_��^�z���ׯ_^�z���ׯ^�|z��ׯ_^�z���׮z��ׯ^�oG�^�z������=z���ǯ^�z���=z��ׯ^�z�^��z����������ׯ�z�����ׯ^�z�=z��ׯ^�z�����z��ׯ^�z�z�^�z��ׯ�׮z��ׯ^�{��w����{�����wE��uK���oRˌGEm���]]\�|����+��1�	�t���&��<z�Y�C�6�����	�k��Hk�2GT�Oq�x����#_Qr�2�{ƛ��z�gY�c�+	�
ڹxo�=�!8o�����[ =��Xݽx=����fr^�Ȍ��'�m��p��"�ɩ�9幚�s�>��Mr͇��(q�:��J���QO`��Dٓ�k�T�Yw)�hb��;w��n�|@ٺ�7<�cR,�>�DǑ4s����Y�;������ͧk���-ވw���L8�_��@�x���a���v[{i�zX��*�(L�N���j��CJ�4�R��
6E_�o���LL�M�B���V*��	��F`rc\�j�́&�͏<��l���� !F���۹�o��34�uD�s<�É!��3;ӄ��fs�Z��N��}t+�8��|`�������M��E��* ��u��ZYY�����8�r��B��RZ�T5�]��3��k�~�����,a��v�������I�c��˱󫏽�4 ׺�&t�mC���Vo&������^����;�؊=)�;T0L��.��g��0g;ʷʝ��s�L�7��ѕ����6�W����o��4h��7��e1�^����k�����z�~�o����{�sׯ^�z�����z��ׯ^�z�z�^�z��ׯ^��z��ׯ^�z=z��ׯ^�o^��ׯ^�z��z��^�z��ׯ�׮z��ׯ^�z����ׯ^�z����ׯ^�z����=z���z��z����ׯ^=z��ׯ���ׯ^�z����=z��ׯ�^�z���=z���������=z��ׯ^�z�z��ׯ^�z��ׯ^=z��ׯ�ׯ^�z��ׯ_��^��ׯ^�z��z��Ǿ�w��������w����I����W���1�N�!KE�U��n��{��Pպ���)AuN�:�v�t�(Em|6!��f�˨��og�]{J'��!�9x�\$����[�'E�|�a�G
�p|��|�OD��R;�\���O]�	���]'���so�+��򫤲`���]���w��{3�=�����V�g����X�K=�#�"c]����9Y�a�����E���T����rl��bHCf�)��~��7AeL����=%���}n���4tf�������j�kc�݋s���T%�f7��W3Q���&;���B�x��q��՛�2��[9�1��B��u�&U��+I�c�ܽ9��w9V!�^౻J态Ҡꮰ^u�A��&�;c_u�}�x�;l�+G��q��]��p[���	�"��I��>��Ϥ-��j!�R�Ź:�)�q�wf<�����\�NWF� ��� �q�̥�wz���NVe��dy�5U��p;�͇+\�P��/.1���ɓ&Gu��t62)�����n���-5iܰh�i<sl��W�$l<��^^9z&i:Т̤�z�Lò�q�ȠsHc)IbܪXj�Un�� ;���%�3w3���������"�#�����p���.�v7��>��r�9;ӄ�R�2����2�˺/���Ai0��BfS�2Z��!.���7i��u���Ot� I�&p����f�Hr7�n��}��;Q7¦֝��&�;pM<8����΢L�����XG���Y���ؚ5Gj[��C{�ͼ���9�c�P��W��-�b��W��}�+���a�?j�yn�d�k0��4{awk6��]���ݫz���(<b����wy����)�7\��Dy�@�2?2���`�'x�ɽ���u�����|�n�y��v�����]��S,6�6�._nB�q��;SX4vL}}�F�TN��P9�Ee)J˂t�Jj�c�ξ�����b��L����Z�L�����\͞�$ i��*v�C{���lX���C먨�Y݃/��x���7��`)�aD.cb��E�|��x�ݘ|���t���Tk52���ERb����X�*U%�ݬ}բ����rw_��m.#�˪�܁6�γ������s�W$T$�bGT��	���Ө�ՃQ7hڗx��IE���r��z�[O.2����hOӊfcqM�,.`�pߥ��0�j��
�Sh�xe�����p���ːR�d���Yօ�LX�46r���7�.Ņ�c흻�a���Y��M�E�B �@�NW�2�c"��n\&ZR�i���a7/��1 Wm�P14��>ۀ��>�	�ƹ�y����b����r@�d�9� �%�q54��xq��X�i03��D���c7!)��2�����$՘�ۿ��O_@�{s,}�*��==��)�FΗs$�2��S�M�h�0�3�@֏d�\�o��[��h�����t%z�H�-vQ콳ƕK�&���o�I'�> ���e�����(�~!)�BP+q�	��O7Zf֨��δ��U�ϰY���Լ������x�w{Vj>�4�����*�v(��LD����W(��ViZ��r��	l)�(H�!s3u/D�L>&��%e�7���d�]���".�5b<^��RtY���ɚ�	��sؐ��;���L8��dɭ���咉ȔI�Xw{�9p;y�����S�-V	{�
���Č>��H�c��͞��Y�7��V��|%�dƴ�
P�Dn��w3���7z�v'ȓ�_�$�'�>)%n�u��Ən���fh2}��ͼ�Owvr�d���ND3e�����=�����;vի]���k"�罟f���q�<�^�[��&<�c�S�ý��i��1��P��Y��ʬ�U����۸.�#z#&��`,X��+ٳf�yse�P�#���>L���g ��Bnw+�{�gB������y�84r/ү��E�t� ��:{uI1�^�u���V+DN�e�h��'o+i����R}�����;���y���V$��I�S��h^�-
�ٶjܶ�X��6���Yݤx���Q7�|>��98�^ �k�[>�'o%�"�M��MyӁk����o�I6��ٞq�_x7���QW��� ��\��ڤ�!������b�|���3s��,U�o8��\��aZ�Z�8��tpt��a摾Bbô����yT���0�K`~��~��[�&ol\��b��w��g`�ub�!U8�y��#];���ؾ�j�,��=�/	+��;��b��AWݚ��&�Y���cJ+è'0��9zp�'�f=X�Ҧ�%j�RZ�݅�)98L����2�w7�:�ƅŋz`��[=���]@α�GqwNw�L�`��(��i�������5�}��ǁz���`Hvz�
�������j�C/�{O��<�Ҙ�6H��2-�GW�'��Y��������p�pR.�CD���{qQ�H@C��-5� ��0{�ǏݡmDn	���[�cv�i��f>q�Bfjs���Ɂ��Թ��CB���8z��;����Y\���}��z�V��ތ�J��z�`;��;a\��wҕ�a��;E�"�Q���!�h�96ۭ�8v�Q����D㓡9:��
�F)�0"�S#�N��J�w:��&�^^�P�������[�4|�3U�|�Jț���{o%��X��B��{����_��,*��/��Uj������̜�F�<T��y����;&�L��H~������ ǶN_�3)�R�o��"-���'����7]�X֫n�*�q���9jd�Z���y��j>�go]Ҳb�9f�Ʒ�-�[�����tE=*�Haݡ>7�����^Z�m�^��8;-��͹�,`�\���ܹ���[�����c`\TzV�v�Ͱ��k¦_�̟5����nxv)�-�{B:N���fkOWP�x��7J�P��W���@2�]��y��W[,qؤe�l��Dģ$Pѹ��jњ�6a�F�2�m-6y'��]�VmmI|Q}�pv55��+uK
q����}:�I��]�1~�w'�Z������w�S<�#}5��K`ozS^w(�lX��2�je���f_U�f0-�BWݪI�S�Rw��G�Ol^�eeʾ��x1kr�hnqY�%Q�v��Ĳ����ƶK[��`Fs�57!�Vt~v�1=�������<N�${D�kB�C�V�ɛ�}d݄��:�P@�(d�d��n��f����=��Y�y��i:E������0��;a��EHJ�ڭ�t�8Ӭ�K�<VO8/�i�9�L&�� _`塕����uX
���krv�=�o�����';�Og��"M�C�`���X�\'����]+ڛ�CNCy&.�mW��d�gk��B�kr��(���裞�1��E-�\Z�Y�9+�V�z��~	�/���nO_N�<@,�Y	�ё��؛[ָhV�4q�n����(xD�A`�CU�]�Ft�Z�V�{�i9�Z�2��,�7�C�μ��9zoY�y񝲲o�l��_����Bϸ9��<]W��Ꙁ��8��B#�:��|�]�Ɛ���"�
>�tu�[}<�"�
�(n/ӌZ�:����m�um�-�����6)t�X��w�ШE=�V'c�2>�M�DV�N�Vj&6�L�`���E$p��zG�v�иwu�T��Po��Wl�I����� �-}�0��ǝ�3�%1N��>^�YΌ�zX��>xφ�^-�Hvq�V�U���J�[�}�V��Z�v�T����{�$�JJ���&W�ܵ�\�K��X_�s!&w.H?F�;�'I���<�O�V���7��$��#=�!�{�~��܇���E2���Q�p,���N�[׀�W4��Z拈H���R��\����jw��o^�p�����,[�ݮ��f�ũ׏��1�5y)of@]���y8$$��^��6N ����K-�iǚ�`4[��ٗqp��F�A�{|<Z�ԛՠ0���]�{��c�'̀6����an��U�uY�W�����ƻ�f�.\A���-�g�g�>�P�r&*�
�(�m�=�%�wG,��$���-kM����Z�p���i�upT�c��^#���U���z��#�_�հ��5�*��[;�/6���rz�� ���o���P)Oy����1��B�'�o����OJ䘯$F{jٽ���=Ǜ�yj]JvL�������%L��I9��R�u�PO�p0�gEzQ�aԭ&�i�����}=d\�V�]�P�yv��z�p:}�|p�imh�����-���g.��N�WI����S���³���1u���"��(b��xt8��uJa��v�a��M�9q��]�+s϶�-���u��X�k�nh����{x;��&�+�-D���-{[�x�n�/���8!d8�f���
9z�MnmES	��������W���w�����L!�ekD���^���	���+Ǿ�����{`��Ի+�`�%�N�\����Sp�۩�^}Mp%%Y��)�{�h�ѵ��^��H���Z���X�i��{�U�)����|)t�z��5�8�Q�ٝ 1�ws�`ㆽ""n??#����ͻ�?]�ג�c��3*ӡ�U_ ��;�_l������P�J헷�\�[GD�`�;
BKdP���s���1Z{�����f�xf��H�����zW�VF>�Pk�r�fw[+�[�V�!3��� ����S�ǈ)Mu�ҢƔ��jl��z��Á����Dm�5N�e�ĭn�ʹ�xw�����X�v7]�]DQ�:㗽m�c��@����!M����m�FRw�T�TE��hh��8[��x��?������/�S̱3��v�-Fp�E��W��͛���'���W�X�I��j=��jl�͸n����n��Y$�%��Vˉ���%<�ܪc��gw��ڱf�<{�
�t��.T�+ٛ����2�;���bS6�sR����;���_6�G���O��ΔqY(��8��ힶ�痍����~� D;x�b��%���нGC� !���N��@-ի���My��S_c1{M�6=�%61J�N��ҩ�������=�{����M��������O�/�������χ�<M������jO�
GnBd�!HB�b�,���:0YDțQ0�e��l�S�f�D���Q&0Ӣ����O�@�B!��e��G�W1�k�)[c���_c��V�Eڪٮm!i��j�k�
�(����ɽq-�+kD]�ʘmJ�p��X:N�v5�sܬyܑ}����B7f���-���f���:���-���ȼ�egӜ�-�.G���~^���ܤ�Q�#dp���1�^�X:�.���t�=�ذK��{O��;�v����]�;���)�S*����t0[�r�X�_^G�6�}�~7��8�}��da�3!�e�`|�f#[����0<��na^E7�)�o
&̘��-��#��2�Nd�ٞ�Җ��Ӄ
��=�qK���}l!�q� fA��
�ZQ��ӯP�5*�&{x�yv��N��Në�#X{��W�R��K<=�wmk��a:iG��|��3s0fB�v�e~ho�	���'#Z��C7�v�zs�0���H��$[7�v��f��w#�d��m��=ٓ�ԫ�~��8mp�J�K�h�׻M�\�-����pi����6����'�ǾO�S(�5�sT�=�	-�ƹ֛�ݹjv1���!���Ϝܺ�qѵi�����x~�L���m��j��	��5��e�0������)� ��DJ�����ǘ�q5" ��S3��w5�A'u&�����Ph�YTT���fFH�a�&	��%��*�P@�~L"H0��y�h�H��\X�/:�2Pe�ב^�E4g��r�P~BQ��m[�H�%�dN�(�'ʛ�)��d��q)(��dAKĔґ$�0�Š��,Q��6���,�O�%Zu3T��r�T�b'[�Lm�*�i.Ej""�w�s�sѴ�
��g>�>�O�ׯǯY�ׯ^�O�����^��4���Vƨ�:�-l%UcE�(3�p�5�_x�-{�m�8��h�� �C�(6|�Eu�������z����=z���������������(���Q�g��U��PVڂ�7��1�ۅ�b�-�S4U�ۜ�ͩu���Eys����N(�Er�r���50D�Κ��1����*#F�������uk��lp�;�y�\�����<ƨ5��<�ERUL�ꩪ�m�cUPTN���Dr���&5�����5[i#N��7
��f�Z1U��.�������4bi��lb�1�79Ö�9�s:خsE�<�*-��O���9b-�\�c_�c�E���刨�"�8&��Ī�Z�l������01�)��	`�t�,���߂��1z&�UG�0�
0A�B���#�ص~q�^n� D"q@}
>��E"� �A&�q�A0�a�� @ˌ�d~E��I��Y-������Ucr1<�q�
0p��9�OG
�E�y�xcU`#~>$�T`����JI �Biv�F��D���7�W<�����Dz2�!4�M�qC�1 $,��'�3�!�d)$*�xMcA�ϓB{䈔�D�5�~jo�F��&m�)��5($.�1:�Ֆw-��bARA�u5"(�s�uǈU�;�w�.�W
��YB���M�B�E"�RA8�l�B	�������A�����n�w!`�ѤP3:���~���WG����m��c�95^�3���yǙ �P�Uu�f圉*8����٩��b�s�p��@h����@gsz�m➇�]���+�zMߤ;�ݯ6�4O�.	��I��pr��!q%��4R"b�ۨ1��q�;����]��v�swV���Y��v�zk)�J""@_[BUp6�+�d[�\���59*�T8��\�<���{I�h���c������R�<�`�M}�t��rչz�2�.�z잮�<��?>��9�qj��C���]K#�k�d��?Lr�K5��f2b�	�᤮j3*����e�7��R��'���V1'f-�E��j.��X=���D�����Ye���k������k�.�CS��G6\���8�L8��*���1԰��qs�̃uJ�0��BP���vbn�k�z��
Nml�R��%���}�J}�c�������	����%�dt-�t 9'�8�w�g�+���{g�p3������u�3ݴ-�+�ᘖ�elZL���{��>!t�K��}�Q_YOs��G�о������g����M_���e�;L6.��sP�;�=zz�r#��h[�By/v�_^�}��}W�f}�d-�E_T�3j$��r�3˰�ӽl���x1�ǰJ��l�o�Z!I�ν��"bu��F,p��j��_'��y�ui�uV�|�tg˜��"#�X�70U(k:l�Wb:�D�����u�n�]q�_.�"u	�wl�ij�ׅzd��χh�T]�89��Z{����B,��#���;�=f�6��{�1=��<��髁"���{>��mW5l�#�,E@x�t�< T��X��.��V�<ZS����R��'�0Mï�Gc}��N
�H��}�n����ևI�<�r8�I���kz��u1#y&MH�Ȍ�kM��ۘ]�n wJV��K�}�+;>��Cz�'d��"xw):j*pYwa�h�Q���/eA��EM����P�E(�շh�r������~�}�y�[�fr.~R�(����>�z�������ѯ1�\)���ڨ���ڶB}��LcC;q\��+Ҳ�"�<� �4;ٷ������i�50:�����o�'�����O�ra�{2c�z�7$��b�{;��v�tI4>��u\r՜;� L3���=�����i�����h�Л�˚�R��J��.���k1DR@��P9Zc��<qM����bYЅ}ٛ�Lc�{F�|7��F2߫:���yQ})�@SSS��1�q�JT�L�K���F��l�7�
����+�>���]�.�5��s�b��/�J����	�D�6>{�mC�e(���글�<HM=p�EX�.���gn�Y�<n}&�b)�M�W��//)�.�#�Ѿo�x�d��S����OW�٨fQ����tb�%VJ��ݮ�O�x8om���+�aBƷ��/:��^yn������+�mW(���n`�͟m�������
�`����a]���Aŝ��#�����,{8 �d�ɣ3����l�־�k:�\Q���iz�sc������o�%����6�zq�r%}u��v��0]���E���z�7�w\J��>��]�fC�����|�t�����^F�ph=b����> Z��7���N�p�ː'��j�柧�54#�@��A���T\4Ζ�p���SQ�g�o9��y����庯+�N��?.���\��޾׮k3xO6��}�#�� 
���H�����{����m��\(;]��#���t�7`>��>�4Nko�d�mǈ�Y����	̉�&�_7��9}(U�jv�8�n�	�*n�����>�f��S筍��O��B%H��P㌸[�1�2ݬ��ξ�c���\���5.o�ߍf�5����5��u����1?r�LE��Շb��4�IeO-�$���+Fww<���'}�31$��B`��1�_-�wJ�@z�-��i��3���q���oPt����h�@�P��7���z�n?}/{��/|�ɏ8.K��;6��l�><#'�@��9� ��bfx2���@C����v/尐`�/tוmu�
af*�7����jc��IN�r��3���s��KF]@�79���%���&0֙��qO�TA���ܽ�z�篷Emh������"�p�z�$
���_X̪�"^-��6������``�%/"	-��>Be�krM�ݝ������j$�O8s_(�����$��6"9!�k�N\f���p�}�N����7�R�k(p���z�]x+����xP��G��=�[���!�=d�Aj/�����S����_CݓB*仃��$fDA�oo�Mb�:�GT8O��}�������k�p��(}�V���j�몡7�{t2گ���o c�r>�DF�>�W��f�Fm����u�.�$����έL�]�1�>�7�v|b�"M�A��q5�D��}ceژ�C��û��|�ڮ�4���{��>��qQ��D�îk��UU�<�;V#�U��Z��E�Eq5pv�[�	�&�+����7�'>!���}�o�U��y��L� ���I���R��@�9;":U�8=�b6U��ċm����ë��<T�{��wN�@��/�kGۛ0��9H����v��f����)�V�+O�I��j[�t� %�P�T0c�U���T�s��	]��˩�\(�b�������{tU�ي�f+[jp�p�$�i8s�h�����Y4�؈*�<�n��|7���uk��X�r(�����~��M��~}��F�Nb֯>z9�o#�RȎ��d����z�|������U����2b��{i���|�;��K��m�N�(Ó�j����U����q��LuQw��e�M�Ck��T6���Jܹ�]hH�b�[� 	'��&"��*�y��}*��7�f�ʢ�;ە��.a�M�����B�mG+��7�����삻��Z[��S�������|��n��u�D��\�C股t��'9��N����*������dKl�/v��Cx�ޮK�e��K[V�y�;�/�j��Rc�z�����i6N�	������F�\&lج]�ky�Ր^颋��d�8wn;��q�W�_�wAk�y�#����7A�����-CD��j'n�DF�눡|{�_E�F���A"N��Ii��x��r�t�d04/j��|�8u���Ǳ���8q��>�i��嬣�S�3"W�F��YDQ�fc2��uoc����ͬ(gp���4?$��.M�5ĉ;]��A6ђ5G)�hw�m�o��-�E�����~>>�8mWww4FJ�Os�[�0W`ٯ�;n6,\Ss��b����J�7g�h�9e7���޶��לxJP��Wn:��_un�I���9���F�M|��7�|A�$w&8�i��Toe����T1�IS}sc����u_(t>o�qͥ��b^_>��Y�Zl3;%7�v/���k��w���t�108bH�Z���s���@&�M��&Gu��95���s{Z�;O�@2.&��;�n��E��w�������ߊ�.�W/#��۟oۻ�'��d!0���5�	\Tryv{-bϩ ��@�Z]V���z ��Ο�}����������ȸ:s�������ԗ-���|\GI���v[B-dLB?f�Sp��F�=����&N�[��nͬk����K�b#��Cp�Cj�j���"k�S��X��Uzb`�B-,{�F�\��ko�w���5�}ҳ���.�4�X�<��#���ʽ���D�WQ;f��&�CM�XZA"�ko�wU���Y�z������y\Z%��2������U]��.�<v���3�7kAbU\�%o_ �
��������^��|ƞ�*����z�#L��tݲ�g�>���P>�7��ufg"�u��t�D���:�������ӟ#A�CMF>R�5:��診�t�.����+���$|�~aU}��쭷}�"�Yb���坡@$-hƵ�����cD��(J �v>��w �u���Wo��u�Vh��1�b0����n�s2!���pQ���ųose���t.\�tr�'͜;+���&���hA2v���Ndl�TU��T/�Z!�L��O�C&-E���~�݋�wϹ�?�����2;t�f�rKuA�o}p����8��P�)_w9|�JΕ���9��xh�[ft�pv�ˎ[n���
���D.ʋ�5I��4�6��<����Y;f�t�4��d\6���W-_Y>�om�/V�&X�﫱�E,�N��b�ȃA�g?cbnaT�H��?��i��N��-�.�N���+Ё��B�{�;�x�����*7r^��F��'���U̝0���m��4�;wM�<!�!�γ܂�uSv�ѕT�^)�u
��"- JD$ȯ���;�[۷`Uq8��w�����|���MA�ߴ��W\�'3	٘�T/z���;�����9�]���Rx"8����a�����"�,C��A�n��m�Va׻�
�Dn��5�}� �b��.#��֙�HD������) 姚���(N�9:��/R=�GR�9Ŝ���VQ�[o���-n'�{@�������π�g��	3d���v�Ӧ���|�6�*�*{�pm��WÛ/�h}fW�Xs��c�y���a��z�k�7��A\��g��p��E�]�ŉ���'m�h����*Λ�w�z�ۼl������B�زka��B�p>��)���=��b�����>��B��[?t.������+E];��U78h�gy��v\��#`;��d\��o����@A�-���1��"�D�|�91W�!��9Z�׵H5t��ٰ#��ꅯ�`�hn9�PFS{nYLc5�����C7�4 8���o���p�3����Y��ڸ�@=8s^x��̛�qZ�(Z38�o��ÊG��8�;�!��<��P^ �~ϳ샻n����?4�Oz��:��H�\N��ú��������2�����Q\܂k��[�}�7�n:�p�]ۏb�4/z�ՔS惫�o�;���$�����k�;��@7 ��D�ΐ� >�8�6	r0��%��ƃsƁ�3��l�����<Xk���@�Œ�Z��-ci�J�/��*{�Ns>Z��=��q��G\�#$h�)W�t�����}1j����w�a�&�c����'���Y���Y�,�k��)UD�5U>��90��1�;���.��yƛ܆���$�ie�y��%���ݤ�m�|���_O��8Nb�EA��W���EL�u��5gse����s�����D�����ugX��*�觔�)�v���,�+�N�5j��[n��ي��{��j3�}���������{��슁7���?=����{=]����m$eV���A��56��(9Qv�N�e�E��X��X�g8#��Q	��O3f��cw'm9�X9�3�j�f}�
s;�Wy�B�Jf��
(�٣���<GW�,@k�e��aT�g��g_��r�[����2���[��u�r��A9Q�L�q�P��%���� ���O/��b�Ly�W�H���lՕ��y�z���)�s�G���k��{T{�^ȧ�n�o��|.��w�����Pk�!nb7W����E���`�4n6-�$���R��<f�X��/�V�,��>鯭3ؿ}����(.@�&��p�����3�����z�=a��o��73�6��N,�P�tn��'3#V�!�z�����J�pn��o���D��#ށ�1}�>/]<����u�5��{Vj�/O���2o;c�6��
�c�_y��3��h�8]��B�r)Gw*��qγ3�ajP�1s�˫�eѾX�C�ѝe=���_ nu1��7��LZ;z)Oή%��p�Se+1���$l�2�p��*�5mm�>��[������ V����u���;n/c�d�vXm8��8z.�6��Ǥ��Ot���c��\�.��'Rv��g�X�z�7��ah�n> x��H�̎ۑ[��K�)��[��f��x�z�������i&у+&��h���g̃Gh*��Պ>B��,5�^`����rII��E������\x ��̋}��Ⴎd���MU�!�k*��Z�wgh�����RQ���N%�V��X�0"�a:qF���'����=yl��V]�ܥ�1�.wG};Y�#`�oa�9v���&�����Z���g�������Ud��G!�#�c�N�y��+=��lѣr���+D5��q!���zG:���^���ߚ������Fr4��(/36�Uga�lB�v�3d���8���O�����2+əÑwE��Kc����^��վ8�!�M����W]G�F3U�5KG��r����h��^1veԩ��^����V[����CW�랜P9��'k�P!H�6�zG˟,���ػk{��{7��Uީz��zcp�pSw)�I�G�=���[�����8�TY�I(��4k������W��9ݍYj�3���ic���F�a���u�#X5fd���T`2�kS<�ˬ-�.��d�V���~	��gu��˕���<9I.�D�}9�K$�sgݝq��˼�F��p�1��;u�$���ر�,���P��V89� ]N-b�B8����h���D���Lڋ؛[2$�����W(g�3vEEVL��Caٽ�r~��v?Fo���ɇ�oL�l�-�m�]���~��8 ��^ �Ä����_������&�7g�єi	$��P5�f&<"I8"x�)��>�"�p_�l�M�sh��s�W.p�(����9�*�kk$F�����\�7������z�z�?�����z��������?a�ϛ��ˑ���9���9gPm�J@��r��f$�!��ۑZ��1:��mˇSI��		d¥���F>����b���-QT�"���+�����}^�g������x��<||}~�O�����?��8S۞C�,�81��[�6�m�m��j��3�bݎ=�"#��v�գ6��7�o-�9�8Rys���mj�����,��nr�8c�8D\ŗ5�m��-���7.`�dQ���$�A	�!2�G��Y&�l����!%�H��l�[!�I$|�i���'�%�P0���ȸs'*�c�5U�s��d�-͋��	�9�TDr��s����
��gE�CLgRFƾ�Ky�U��w�ǪE\�LQW9�%��D\�A��s����幚(��f
�)�-�sO&��*��TmUSE8�km�cU��Dl{�{�E풮��y(���MU!��^�E\��4���fъ�)�uQUQ>l�:+5UT�Ƿ#��T��"�<�>X�
�g���& �
&��s���j9���*-m��M$�T���mnl�E1�`�1SQA_Q���-x�����S&�lj`���
D�~$�	��]P�W~����Kq�0]�},��-#3t~��7N���o����;�q���d��ws55��}�?��z���5zX�]�9����f�x<pݬ`�=Ћ����e������u�����2�^����鍶���>����e�/V�oٴ6]�s�E�-��T�7��p�^ʹ���S��@֧v�u�χߓ+��C���O�������"�~|�k���И(f͓(1�Sr��T��]��׈������(ި�V��VC�h�伀�$z��s��y��=�E&��m�Xb�t���nD���������S!k��VT�E����{��[�'�|o;G�(#K��K�ȿ1�e��<3�ʙŝ���4�c�.��dU����):dK�x������ȡP1�>O��qm�Rq�klI��Y���ɩ�J���=�A�)��|�����H��勺l������<���T.�[A��)���޽ԇ��t��Ʀe7��Aw;��	>9�NV���a���L�p2njp�b���K�}��A�����B��&hLpm��i��v)���- u@�%��&((�,���^ǃy��>q�ǁ��,�~l��lW��q^�S��Km�޲ٞ�E�}��~\}�&�cftu#��w4��E)¦^	LX��zqT�^�b�I��=���Y�f�+��=���z@��"���NS��iZ�m,��K<���9܆\�UdR7�C�������K���ʘ c
!�)UqyI�e�[��������_f�T���G��dʞCpگ����蔀��#,TWҹ B�S�~_A��G�O}����ז3��Z����ڇK/弰����u?l�_਌cH�ි'W�̏[=�>y�n�q!ﶇ�����Z^��k5c��=]Uq����S�(��A�2��h�k�HD]�ܨ��4sM!��YX@��	E���B7�[\|�j>�(0Ӏ�_��Ҝ��t�P=!ƨ�Q]u'�����P������F3����"c�u =�7�6C��pׄQ3E�v�9m�S�cGy���cwkLR��=�hk}{��h������xu�>��Sc |��u�� {Ȍ��\�ĕ�J�ט�.C�gBc�������Ӗ�x;]��`0&~����&�zz��cp@�l��w�\���y�����Q>A�X����p�ز��e5#�%=����ϻ-*م�Ga��7��ݻ�w/|�a�/��i�A�Z���L=�΃~�*��ņ�S�rS� ���dU<t!��ӝI^^i����!�I��b~r��6�+���������#B�ʤ|����P�����8���p�rFxU"ಹ�ț�SCu�=\n�N��N��?询�|��;�lP9��L*�WV徿��KtV'��y�a,�#�8�>�1W/\�{n�($L�NVl� :��JB)�a}��n��}�o�A��9:�ܨ�A�b�M}��e��o��%"C�e� ���{�����ʾ�g�7>]����e���!y�~���M�F~��i��-ם����ȣ�o��'�,��/@׬7��g��Q��iwMz�7���ds$�G�P�[�hI���B�ge��ÀC*��6^��Ou*L�p��[i�X���oyf��u��4��������*���<Ð��� �y{aʷ��l�;��9u��{H���ǥ�6ĺL�G�c���4�O>�ߙ�����B�b��!���A/�8'�қj��!�-�00�M�~k��O<���b�),c��m�H��A�0-Ɛ)�y��a�ѭ�T�X�^bHx��u�yN�)��ߛ��]���X-�4|���$���sS��p���T�Z�jiW���tN9�@4@�`��.�&5遭�/MxZ�2g t�Z��^�K�xh=s�=�q��G�y�ɬ:���4�xF�?���B����<�S����~�s�4|��V���{5j89�r�^l�(�Y�b�3����[A����4
����?p��z"��@u��[N�e�ܯ{�.�V��{`8��3s�a|�CL3��<��'�}�Y���Y_)�#?jD�
G�+=�,��yO�**-��T!�˅Q��5B��ȑL��"����j�&wU�K�`��9I�A��'��vM�h�Gp�ko+[n�=���+[�u��@D�N1�'�k�N7\�`��Æ�{5sV7]{[92��H>���U>c6�Ք�"�3"Z��]ʭ��^�?��y��;zo�=������4�O�&¡�����G=�,�QJ�l|	XxL�"ˎ��f��&ie%wvp��o�u/i�l��j��^��^n��Y!
��k�7n����tSG��:�,��������(z�k��q1w5�`K�*�wb i��!k�t�j�Q����<���Q���I\�ln5emm�&폪�B�⊏g�c�a�#��u�~�mk������d&T-��Ln�c�i����=�λ������z׫xi��Xߺ0��	��mԆ�����k�4T�����r�Ֆ��hjw�k������K��3��+Dl�*ո����@�$@�!�,�����-�u>�r���̙�=�)��2`��S��d�qv���6�yQ��5Qoڷ~T<���M���.�Q�k���k��WG4����JD�4��K��ЍL��9�X���_��� HMw�����Bdg�wnfn$<G;43�~n^��L�Հa�}`nRwGg0>��#c�Z�AcK���A���(���I��t�S���}�ז��._~���QB4�	��t'���j��.�Te��#��XWC���O<�K�Q��*�U�X�#4(v����;N�`�żYbs���A�,���S��=NP�6�޺�E��c�h�CaY04�u�U��u����r-����3P�a�bJ�V��8ɀ����I��>�̛�������������Xw:�Fq�q,�ON��#[�{���ֿP���S�Z�_�׍��	�X�4B�	�X��vg�iY'8�Ξu���)���?]�@��t�tGyL ��*�Ob�ܛ.+u8/b��̝:G��k�O���J=:�LsO���cf}8@tg���aNdf�]O$υ�7ڌ��,!�>��b&ߏ@v���<���Iz$G�mb�>DY��!r�� x�����uV�%\���t�Yw����z(����^?v�M��wk<��;�������Ӱ_E��b*I����c4.�����c�Y_�?�0|���+���*�j�}�6��W�W����](r��DO���>�m�zs;=UռCu����6���(P��*!�tǟ)z��.J������f��,�qv��D��=�z������ �l�?{^��ёN�0'�À�*_G8��T���Y�x��҈���H{N����.��4��{�V���@P�V�ʾ��0���I�^�_Qe����LX��y�\!���&�9��&%�{(���*Mv �Xkތ)�8�Hq��Ŷ6��Wr���q�LM���fpݱ���Yi_j��:���s%�cD��Ğo0���D�e���;��z��Ml6C���f�3.����1�b��N�m��GN���[b�2�qإ��
�Xu�"�cuhd[2�⌽�*�L1$��";��������m�]�3C�|�/�L
�3ݒ�ϯ���O��dy	��x�"�Sn��q�<id\&(�{�P�b�g��ܖ����c�q�����0C��0W�]�3��$�^S��^@��0���ˋo��G�)GG�_q�L =/I�" ���/����=q�%�v)���-���bӁʈs�]�j춣�ڇ�M:��y
��a'�?/O%d}��M��?�!M3��U>`C�;3wb����%=�9ϻ���b���<c�*���tYzW�ء*�� 1�:H]�"'����lL��YN��"'��[�x�b��[W����?5�lx���W>�UV�H���'��>��:�v�~48U[��E��c�ʩ��i;�6��^3%�Qx�Z��0��u�>/��!݀�� ���w������O�L�6>@�L#��ƨ	G���B6�i���'���D��6���kr�u=��[�"�m���e�YA ��1�YF���� 	����^H|~�ݦ�Q�/�� x�_���m�߷3;�35��U�?Vg�ƫT����D���/tZ�~�R�^���"�J����"����ch���f��4O��Z^��˽����: /�{Cފ��<G+���R4�z�ya�Z:�|q�N�텬|��Ћ�~ۊ��8X@��T�8�7�w_� ���LN�n��;R�i��ݬ�xo��AQ\[��Y�w��7���+kQ��'u�D8�A�kͦ�K�{<��#���zyY�l��G�[��N�͉�.�}$�,����fρoе�i����6�<zE)�$hؿ����j�˄I?WW�GSQ=�� ��FL�,%u>�͌!�Z�9�z0�V�δ�ޝ9_d)��%X���]���VMؓ�]�u����s�ȸ��22�'ֿa�ըʂF��(u�FG�^�v�L���|����'7���qD8
T�LO<��-"���!�:�	�N��J��G���l��"�Т����Q�x����!7���u0hȸ��o��'�-��z ��6��o�E�!�G!b�kw�c��H�r�C�i�p��Ft�D�_ӆ�6�C)��!�׽.�H�J��{��Y�[wyE��r{."�ųS�I%@��/�Be�"w 0���~g�	���m.#w=¸Ի�u��qsݜ���B/׵:�-[��'��4�/-��������R��a|rJI�n՟a�2��͎շu�Hfd<���T쉺��«�O<���	IcC�Ӱ���>m��C;[a^X�r�P������Hx��5��z^S��"��2[���E�Ύ>�;�"G���\�/��v7�gs�������8�Tc��}�cx�A��,�F�K:E����5���}�˖B�j1�up����T�X�M]i����F�XƿE�fi뀅����uN�H΋r���+�]��e#�k�yLG��o�bUK������????2 �Kz�t�Y�z�0nm�`5��|�����˽4-[�8���V����>=@�k�]�__�ǯ�z�y��*(�W����$!�Ġ�G���P�%��׈�_v�A|�g����3խ�~Y�]����\�;l.�O�@��4��9�"]����H�(���& %��f�;�K��y��������s�����8N�K�0�עf]��c]�00i3`S˼ �-ޏ�T��R!KZE
�$�ҙzr���]��{�ֹĤa���7�B!�p�h�#(����9�L�CX%x`��|���d�(��u���<C K�r��2�5������G�(w!������L��t��~4x�ˬ�ll�Eƅ�1�{�H����Pp�h��f~�9~f׿a�j�I�%G\89�6ͫ)�����W��0���3�B9��PϪY?P��~�D�}_eD�5�[�Y�`&NŴ!ύ/Pz�	|�kOr����<r�.�N��M<4�3��[HO�%e	�ظ��θ����ΘU-���;[�.t�!�6#י@\�@I`��q���V↯~@l-���P�y1{@��;�{GΥ�\���"�7\��qXFy.Q[k`����U�~���ˡh}�O���:�*�{j�m$�B�#F�;1�ј�U��.4�z����+�A�։ǹ���^�H^����^]��x:lܾ��������ם�w����G����NB�x�PC�y�x{�G[U�ԇ�\p����|�Ϗ�K�xz(�m�"�E���>��}i�2f�N�[���[Yxy�.�.C)�"U��}��EL-��,���?.,u��TJ�/��R���e���l}E8b'K�����=�N��*�*2���pJ it�~mV�:|�1��{5���J)l����&uy�H�c��������T���n���#�ۮ��q0���[�����:<�5 2�q���cÚA`��8�#Xw�ǫ�k�zb[zv�[+�Y�	C�kc4�����k�o�����tw�Ұ�������~���P��XV�^)�����N��䷕�*���u�5����v�p���`ʉ��C�3�ס�όu�޿0>�G����%��!�/krD
�{�s����{�^�����D�g�M�����e�zK�"�(��y�@�|:%�ƛ	�\f�z� ?Lu]�n�(zCs	���D���/m�b�z�ﻺ���s�r�#���m�-��9���L�v��마r�Q� �\d��d30���U�ׯ6����u�}%�QW^(��،C,��k�W9��.����d��i�P6*�+�KV@���|E]-0z���bμ9�r�Bn���ٍ45�	��/�< �Ӆ��w��<�������(9���bJU��h��eG�xG@l�;פ<�h�m�f�#��u j�E;,��G� ����<x��Ji�B�i�hR�)J���&�f�{��^orY�X����"G�&ڡ�mF�� $���,ѭ��V�?I���9V�/��rwѮ'�Rn;jjp^�u�C�\�i�ả�y�i���:E%�� Մ����9�j�C����K*���3���	�=�Ot�z6q��YZ3I�Q�1��|��x/B��������5�R�x�T,�;�Γ��h�r�Z�`�������/����O�&{+���Ҵ��ⱉ�y�ٹJ�yh�o6/ Iq�&>��D��K{���S��ħVH��������A��Uc	[X�v���Q
��5� �fDOϨ��0�\c}�`�@$��*|M�)u7_;m�װ�Kg3ϫstVDBN���}�#�˰�>߇������W���|i/Y�a�ݐ[���UIǸF��~�p+�v{nx���\��A/^\�G#���@]��#���q4���Np�h)��]�uچ3�u��'P���b#y�(�/73�T-r\�6�?��z_
"��t����-w�_8�u��sz�!�`e����ez�k��)��i�oJ��}U<2��H���?������Z�׍a.iV&]�SZ��.�sFi,�%ۜ�S!B+mLԒ�f�הȯ��Z�f�e�IgV5�$vEfv�p��҆�ΚJ�#�.ݽ,�7s[=�Fg�}���w	þ+cəl�Gy���Db~���.�Y�:h����$�7�o��yR��y!ϻ�U�H	lΜf���=g��«v��6d��]i,�v[�]�T�?���w^l�$����<y�砄3b{'$F��!׊	�۵׫��h�o#��W��t
<9�
�炆,%:S.Aֺ)l�]%������zl�z��7b,h�l?#�JI!�P��@�D���e�dXO

}'w��������mV�0j?��B1���r}��F��yqW@�=�����\�.��u!{Z��#���DQ,�x��mf1qLўȭ�f׋a�'���v\}�e����wB�U���"�e3r�w=���3�����fe��6V�{y�O�Y�,C��m�|K�|�g��s�J>A��F�	��-��\�(V����dPsE�%Cn�����2�
�������z"�����O��ӽҮv׎��W{���M���oF�B9fN�ʢ��Ś�ViRs�Sɱ8.���2�q���'zj7s^I����'��}"��{��z��^�}�%wJҶ[�5�yE��)h�v��K�M��w-x�!�Ȓ��'�cFn��ǽ3˾���	�q��{ښrU�U��	k�	n�f�d�Ik^d��oڂ,2��KPnL���ދ�M�cF�۾=IҸ�Q�m�G��lV|�J5�'�"���z�=�����c]���<3�v]Y77��y��۹���d��έ�n��=�@�Iga�����u^8�+۳-�ưݸP�/U�y���z�*E�4�;~��uv^�H���6���w�2]�'�>tO������#nqˍ�xu�J��X�T�5-�J���Q'�e����Ws0ܬ�r�����9f�i<h�З�+���H��oX��I��s�V��PR���)��2�Y��4[�_p���~�D�x��(n�-Jo��7�hU×��f�9�3��;��U��qu����h�n83)�C�k�-�S(i�g�sHkz��*����<6��IfƗe�%5�b_1�w[v]��ab�)�ze��ʃۊ�a
�ttHv��P�t�/�s�l>�"=.n�~��e#���k]�j� ��}�e[ƞȎa �;��x�%M���@�̉����?akt��"���� 9��U!�+��(��N�(J�W��iÕ����Bi|��-r����3Jy��h�s�����Y�3�:�w��c��i[قM�����V3{Dm���y�xn�=��܏_Q0�r�a���8op˱L��o-iVt��;���e�ay����`��V������,&Jf�d�`�@b�RF�&�kđ	���p۩F���`H6F�TW����Ѝ�YL�<ٸy�F�-�x�_���Q?6(֊J(���j���qPM�L���"���b(���a�j��9��ׯ����~��z�^��������?�����X������uU|1�b���KUP�h�"J�6MZM��"��AS���g�>=z�����ׯ^=z�?O�����?��������~N�1km�lUh�[9�mb�_M�-��[h�-5A��|�-6��SDTsmb��4��A5�I��� ����F�RPֶ�AAIAL�c�j$�"�64Qx�E-E�V�k4Z1h֝�(��J
.`�DIQES��%�M`�3�9�Ͷí1QC�k��{�b�&�|M�g�)�m����tMQ��h�1���Q�:1�;���0j���E�W�4L��c��h5�+I���������6*
�o�F�$���K�.�(�Bhb\N6t."b��H���{����.�RKFĎ@��¬}�ĩ���r�Ɉ�O_9��n|bj��plNB�𠑅;�^�4��8C���W��A5�������2(�LEe�Q�*M ��BA��[[�c��	���'<n>�#�-u5J*��A堡�Y�'�4�t�]O��2�$��$N,#��5~�y�"�x,4�^5����u��i/���!:t����̱������XaQP8G�� *Qk ����wG"�p�{��7�� ���L�l��-G���K:'�ys`�,�oa��9ץ�D�e��O�}S��>u�ٴ��hA1�bn�ҡ5dbZ�_;6�Ϗ������Z�l/��#4z�0�����sc6G���Q���<��D�����9ȃ]��v^��m\��H�����ZP$�|ă��	kp'��;=���'�4�Tv��qm.5�8c�q@Y�j�*����g��8]�dԮ"*����e���1�\�򷸏pb]}��!�l,����5��z����]��¼�՜Qp�#mhoN�~�ˈ
�q��nJ��pq� ������j�吙W0�^؀�LRu�ȔD�L)�"�k�C�ELZ��y[}{�r$���u��P��Ŭ*���E����4&4���?5�WC-��{k�.�؎q��_f�wHc�ځy�ew���>�Gb���g��!�P��\��>E����eO/RPs7&��ٯ7�ߗa�����c��s�[����[U�9n٭/_C��z���ʢ(-T.+އzޫcqCyh���}�u�g���ƇcL��ދ�uc��I�wlЮ9�n]�G.���h���DWw�'�ئ�f��C����z�h�{�C<g��Ǐ" ;��������������ƶ��`*��"��H�����m'r �a�O��F����C,�~��e�-�	볻�{[�۸u˲*x�X&m�t�niy���<��~�<;�w� �{l�p�M�%³3��37���˃T<0@r��7�XO\5����/ʬ7<}C��?RB�܅�z��=�<�|�u���0�����"����s�4.��ITXRΞcV���<^���먦�V��w������=m(. �`��Be����g��r@��LbK���'����'�ǚ��큫Z�ls�OQ�=Y�{i���5�X�u��'�W8ס��^׈����b>ʝ��/(H�i��qUy��f�`�Cn���#C�O@��3���8D �A3���c�~�j�RZ+��҇�������Oޓ&�:�L˴��-��l����K��P#�q�ֻ��j�/�-e�|�N[��N�1�gt�C�⼃�"��i�L>��< j�19��(�У�%�מ��o��Ʀ�?܂��o���;7�������y�-|�>����F��q����=��]�;
�?n��`tʩA+��f�n	F�J��2yw��?�?Y��(���ӻ*���P��E�UWh�8~�mX�_v� xg��vwk>����I�3w�{z��Wǆt�! ��@2E^����Z�V�7��}�}��<N<x�P�P��ϯ��~���_��#�l.&_~03ǈ�a'w_=/�z��Y��>d=W��%��[�쮎�~,,:b7������<�PO�;8E¨[�	+�20Lx�&h��U'H�����F]�o(��5�v!���xȜ��+<���h|9�f|�����4���27F5E���Ț��G	C��-�{�Pe_����LD��]��1i�P�K~���jC����w�(5���y�� �>��@��~E�����钝c�F�0���2��i7��|� ��eƝ2)�>m_��k���p��^��
��%U�~ǒ醔�]9u��)�-5P0i���>V�e^����>�&�����ˍKZ�Nz|vtY��j���^�E�-eA`K≎ca�^e�#�ϐ���k���G�^:dGG���Q��OI`Z��<q��*���ML�����_'v���:>=Z�}�>�t<o>�":kn��0����> �]n��;3�E���2��m˘2G^O.C�r)���u�&�+��������]@A\9�/��<�:���r�(-���gev�1њ���(�
(
bF�s��9� �I��a|�a��hD�W�����gK@����]��ybOw�F�o��y�/c�o�m|f�os�`�J՛�[�գ�a��l���޸������Õ��)E»<< ���������{��W�o�jC���{��"f۔)LJx��6�3�עc�A떗/���`(p0�n�&Yy��5�҇�6�A~�R�gג�r	p;���5$8;��W���-��A�;�J����:�6�ޱ���aTR�>����*S-#�A?��_�ދ5g���,�MׄF����MGC��
��{ʺ��!��<K��~q�K�Q T+��+�q��/h��.��J�c6�gờB(_O���Ŏ޶��@m�]��z��!i��of����E��
vg���o��漹L@Q���TՓA���d��<Nd� AP�6��$r��͜�(��x��U���-�X}.����V�)�TU\3�÷y�����2�U�xJmoX&d��2=J 	D����FcսdL80���
L�Y�c;�33��ņ(��N@B�ΰ�\P��9�3�Fi��T��Dv, P���V#\�߸��p���������e	��Ϯ=͞b;`��1)�;�讑L��(MMP��yx&��m��#۵��}Ӓ���g*���_�)��
E��q�&R~b��R�pYh�m7X�˦��E����6�����A���A����a~�`8���43�f>6��ص�f�ٲ�G�K(MD����U.�[ue�Y��}�9�ނ�B�K�U��\;-�6�&�0K�QQoh;����s˾Wat���X�����I0�R#��(������<UA7��X��{�_}��ou�^ݓ1�[N~J�2g�v���]������B@��}u=�=��}�7�L��^5C�=|��G�_�%�\
>0a2�K�\�GPFi�'Ǡ.�B@�?@��3�/BJ/W?%�f�aS�ĪOY��2��ywQ`.��^S_<��Ҩ�g��C��/Z@D1����{6#2�^Z�<Y��̉/KҀ�
b��MX;���11�oV��^��~�I�����������O1�IYs ǵP�Z��Q�^��9�è�e��G�L�:�>:�����㽸!,�u]ܺ�>�	/�?ApXTe����R�Y{��;i�=5�� � �N8�hBeݮw�#z�����~v�Ŧ����PT���zKTT ���2T3h>��ۆ��dt���ѹ���a|��0��.]�|�Sj=["R`��}�`2"a��Q�^�Z\�����y3o{zf�)1��/2DP��}���sd?B:�4�{�x5�N����laz�cQ3;f���jCݎZ�Л�I�Y�lN�q�a�Ƈ���[P�T3g���ԎT�q9�������g�Ƿ��r�}���6���I���wu7c�����9zn�3n<�R��$AI���:c-oD�-�
��z�{e�k*�@�s��
�1ܑ��鑠�N@�L�ihI}�6���V�AR�m`�S�� ���� �z=�����=�r�!�����^va^����uV��PB|��xi�����|��g/��ݭ�笝�u��s�l}X�7 �m R�,@\e	���ɦ���C}&+|�f�_
���t�e9Q��zoX�9YX��_b�:b�:�¢D3�5��.��h�ƞ������[F��B>uz�����Yz/����o��Rq]8ñ�����HV|[_R!�3qg��7>�ј��nJ�9���t3gi2�2���n�MX�����9RWj���3	���\\ �����WO9���|hra8���q�i�$�/,����Y-3�a��k�$�J�[Ś�!y� ��ח���pH`����vB��%�tّ=WԘU� s�^9��a',u)v�!���(���]����w���B\�������ϒ�]P�4x޻�j:���%RoΎcG��XTO��E5���j��i�o1�2]*A@� x.�ZDuLezg|֘���	�Z�-��$j��ٛ�<������_ S��yb@z} ��1���ҧ�~���Iw'��֯��i��1�&sfm;����`�n�LL<�;
�uؤ]l̏FX�����+z��r�췜ͭ�X/ �Pߏ��_�-��u�z���=9�_SPov؅���`�ԛx����-�M\��a�V ��y{���^�����QO_��
q�ǂ��/sqR�=�v~d��5�hǄ�29����b�g3��;G��h���e��c1�ʩ���\���ȭ�{�>�k�<�րYԘ�\�f�s�&�3S{E�+ˌ%a����΢��[E�_����-�C�1.���0���G6@�q�����/z�/��}�F}�����{�0K�n=񶝕�u�J��9�!�8y�)���oMB�1�����/��׊�r3抷��2q8��'������3���n�b�z��[S�69�v����մ,���~U�3���6���a7:%C୭+�����:N8z��a^�]��[�J����$?0~�	��!��+-��U$L�q���f�(�=}L{N��0h��[��9^z3��[��)YE�+7�BOA$�
����Z�9qqB�]��#���ț��넦���m	��܊[h���ԊV�HB�O{�,�N�5Y�P��c��=�e��tCi�( �L>�.�tȯ�E��wT�P��-��qȻ�=�-���#`l�&��8/�&�_Aw���t����.���d���w6�v�S��Qp2�e�]W��!f`q��а|�NwYH���QFj�"�f;c�=N�p��6��[�d��	^w���)�^�e��w�
�9��<�����¶��8�ow)F)P����}k���V詻|(��R�G� <3����G������r���6�uY�P�S*?ȑK���C�ܾ����;t�/I���r��
ֳ#)D�.~��>�Tj�:�hI�;`-�#���������E57;<c�Ɔs��y�H�ޑ!lnW�E����!CG��������yC�S�gʒ��	}��?�GG�8uO�Ķ E��P�����-����p5��� ���a(%�¸Z���d-�>�@�9��]�i��Y��lZz2����!���L��K�)l��4:�/�Q�F9.�okv�3�E�v����x��x���sg�>��&�m��?c�%�����7&����I�\ vWtWݡQ�|�\!*L����P����Ғc��3��S~Pp�y!f���K0�DgU�M�S*��w&������{y�}�p��R�k��"*PȒ�7np��}�ܠh(}pN����ӡ0d�l�]�ֵa}a��r�W��w�����)*,G,G���%�X�/I��Q�T��-��7V��|eỆ��֠�� ���$r��l�zǶu>���,���B��{j.�t���ћ���o�]̵o�F�Ç��VM�]��,0{ܾ����n���ώ�T�)������C-5{K�*v��.���M��Y��9��x;#|�C�RB����9��^d�D����.���T�;9�_��]z�}���8��AN
1	�l�Q����^�y�<z=�{� @��|]��5Sˀ��z�����>��af�����Y�Rm&nci���3�(�f=z���nͼ�>�x��bp:ܮ����>�o^fHD��sϖ@3�Z��LK"���d��JV-��e�O�����:��l��h��p�ԣ����&�8�{��|�&[\1)Տ%"�N��k)���^0��ƽ��<_ѹ"i���V:>_@�)� M��]-!���	�M������k�},�ۺ��O�xW8E�S��e�3�^�}�虋a!�"me0��p �A������6w޽ċ-��ڭOe���瀹d=��"y�TQ�,���DCwۊ��V�\����Jr%��ȝY'�NM3������/A�2���"
">c n���׳.E]c>Ө7w^�S�fFz�c���G��p��¹���l˻ �RF�ti���웄OVwHam��2A� �<ö��6�`�4-[�,8�߆�ǟ#��fu�Rؒ�Y��P�����ok��T!��
�@�#ǌ���D&����������DC��8�R8e<Y��mٚ���r�]�rG�N��狩]v
o�:e�"�`^��V����{����'8��١�W��ɛ�F��+S��.�>=����WD�����Z�vx�5v��(���>	���v^�В��ƳB*����|4�XH@���������G������.&��Q%thCs�ui�z����A�S)�|Q~����v����C6�ԓ�3��.ʾi�{i��vu�W��듁)��,�(����/ʇW�fl�JBh�ҡ6�)r=O���\ ���5�%P�����a�t"���4<�0ds��>Zm�(r�Q�ܐ03���A]fE��yW*����]�/-��O�U�m5jQ�4ɂ��W,� �׳e��S[�^g�ӃW(�W�'xd�r��A��{�a]�!Z�w�U���}l.�zN!�	�~E��)O�bu��m۽���
ay�����!t���?)�,ȩ�����^��އ>�������<��S�+A|�̠F�c��"K���C�.�VTxAo@Pd]za'i�����Z�]���L��BT6��e��u�Q)̈́�P�'b6@�'r,ï�w�_O�wɗ��}�{���i�M���o�,���e2c���|m���
[ʂWj���=i�m��X��)��՗���b`x5d#�{֍ڜ��ٟ&9W���!x
��G��R�7ca�r�Ϣ�aŷ����`�������`"}���<ZonqU���vm��|����T��,�I�T��D�C{�ÇU k��Yp�v}F2�Wv��Q�7���Vq�P�ws���G�C�2J�F�*U8h\�i�tƽ���������I�#P�I5��j͚9�C���B�<�M71o[�ɅY�O�������s�MKq0�-�|^���k:%��x�mr�^˂�{_�N����͛�N�ne��F�Ү���љ�6��/H</.�ȷ&KO��v���{�wٓ�<��j�N���?�)�'~�n�ܺ��nIn�HK}��q��.��{WFK��a�����Q���5������Zv�<%�:ޛ㓀�%�5��r]�5U�3/�z�s�q;o��Q��#:�YX8��<�o ���j�V��Ѻ����ܾW��{h�煾OZ2�.�����M6(���ދ��Zf���┗,�:��E-�S��s�I��b� ���˂j���cT�,��}���7nޭPDd}pa�駬�܈�*�st���ti�vo+x4ը)8v��Avw
�u:w=�%'�W�0w"��r���G��Je�ʥ�����[v<�kù�A�cZ5o_p�T2��lNh��,`X��"b�g{[��y.L�#�j��K�\�Ƿ@���<��y��"�C8��b�
{��̖�ǐ![Q�łJ�l\u2Z�����P�[��f�򘦧�e���{p��;
�T�����[r���	���s�ܭ�΃�a�u�+v���8;zM��i� x��cI���x���h�<�/8s��C����:V���n�{{J�S�U����uй��ʘ�u�B�n6��i!H�1U���ӜI��̇�5�}t�����`7�[l զ*� �M�u��c	�Deݟh��p��y|��X�X���#��{s�E��.ܷ��7��[n�d�^Ǫ�+8����j`מ<�N[�Ӄ�^�� �_�x�X����]��`�%v�[p^M��-��Ǻ�V�Qs�F��C�����w-.�s�"���ٽ����WGWŊ�n��$D3��1-#q*�-u���e���_e���}��T���ޕ��[Wj�W'%0�dҵ7U�,�VR|%����x^�h�>�8b�|��u�f]��Ig�"p�3�ׯ6��o^i�b�[6����~��ؚ �c8�Ec"4��0mb��&\�,I(�����){K�b�,�������.�}}n���ُ�>��}�l���C���Bӌq�.��q�蜬[-�ڷ�&�J��6�0���#���_�ʧwRc��k����~-dS�<Odo_wv�o��������Gē�A��$A|�p��kl�0����^Q4{��5�9��������>�z��ǯ__���}}���Б���墭�:�I��jh�&&��(���=z���ׯ^�x�����?O�����=���Tp�sMEڀ�-��DL�0^C����`9�<ڨ(�
)��i�UE:�A%4�_{^��s��42���"�����6�"�H��SETQ%MTMKlj�+N���CTP�by&�4b���A������&���j9��9�b*��JB���t�F$�h���4h�L3UDEDh�i�ANک�*�
&�:�`2T���9��kon��ίv�&.��	fn���X(-)(�l�lꒊ)�6(4E�DX�KcD�|	b�m޹��׮��i�f�֌������p��g�'-,ۖ��m�mK���4��Q�9���\�X�������z�=�G���^�o Ul9Ϝ���{��RKyt�v~��=W�Ȫ��Rh{._����$���H��fl��E{"<��nvm:HEm5�C�I�}9�����Th�����*�
9�z&���~�i�${&2\�S�	����LQH���`ar/MW��9m]K��Okr�T�dS�{�:��y��V\�+��<i.���>%�E����$�ח�������Un8T�Yi�Co��k]4a25��U+zGH%}������Fw5#hsŴ�����]o�a�'��v��)��bK�0�uɈtE���l������zv^rlw>̾��ڣ����25
"cu�='������S�3c�CȠ�{=vT��fqh�ީ[7I�4��`w��<�W�Fb!}e�R����Fd{��yʨE�3��68fZ�����Լe]/�
uIQtH�G�m���+���s"����2�UV>42C�а����^��!������c7,]p�X*,Ň(�ʚ�ܟQ�#��Y_P��S�A��)�ŌHn֑�U1y��|��M��ٷ���@��x~��7�ǈ3��gӿgg�~��?^�yԽKVRY߆�|�mn��T���L]����7�X�T�1C]�Z¨r����IpT��~~�w�����O��ǀ4�q��=�{����ܚ��°u�a���Sm�!7y��݊�`:?{({�ڿ�"�A�XQ�=ҜK]������RiU��B8 ��+��W�H�ļ'<����%%B�:s�YMM�Uq7��$��+)���oH�2�<kBYS�K�L���pE�w��Rt�"�f�i%I�?E�Cy�x�y\Wvn�=����h(�s��U=�`�o��M��y�.�#0����c����WD��Qlq���B��4�շQ<��M���y	��	�#��}�F���g��H��̢�'�49sqO�P_�q�ƗK&ԜKGl�����Ι�8������w��ޕ��n�fH�R�B�A���>�=��xCj�y��*KqA��;�_R	���Ѭ&:n���j�Z[�J�M�	U���+^҂^��8�j�e��枠:CrxyCNJ;I��zo���N��2��QLxt�E�S�g���bLsI�g���V��;���.�Tݍٟt�Kb�.��Bg�E��/d#����^�(Z���i�(�W���M�D+�wy�t��D��C#d��udw�}������5���}9#���E|��6y��q��՗��4̣{���1��AGА�c��P��ﯟvE�dV��n��2��F�YU�f`���%�0(�)�'�dd���J�X����-��#�*�����c,��e6�.(�?� >���q�ǈ ����y�۟?_W������JQ�1ʭ�c�8n��C�����@���ܾ2U�A��q���%��2n�Idw���Y���d6�e�Z-}�L'dIP< A�L�c�)�|�oF��C�U�4m�+��d��}v�+RXJ�!C��q7�rsM�5yg��->A@��Ӕh�/��M��F��v�l�k�+�Q��k6���Ɔ���m���qYO�JUa9�FbݵL���l�W���.���2-��oH�5�"Sq�A�R�CI�X�}@՚�D����L�z�`��L�芊@��1�=v������p.�b^Y/("�er�?��z��Cv^�e���W���״�Ѣ��Fҡ#`CQ�/���Ltd�zЙ'�1)�Y9�O2��4����	�|S;;�����u��.=�n� �<��>,V�$����=0�o��p:��L[�5���g�R��aE�5b�ן#ϯq���b�:2�J�Gހ�/�B�����u���[����qɈ��Y�^�&.g�I�R8�}�F��M#���,�q���v�bCPePuLFdU����Pg��y[XN:z/X��s��Ӯ�:��5q��Tm��T��:�q���=w8�~��t����h��w�*��i(5�}��{F͐������2�΅Ym$�ٙw�B3�Tἡ�J[�쓡�� �����xG�������$�Vf%˅8����=OD�oU�U����z�r����A�C�%x��X�5D��375Yʳ��,{㚜&[����작G�t�V{�Rp����W>�U#+��:н�yw���e��/��
и���S�"]�/����Bչ�ì���Y���j�~��,պ(��ՙ����͇���#�`@���tƇڠ?��3q��a@��y�Diƹ=c�ǏE�B=��}��xו���T�*�D;]s��O�3�(���y��'}�U�-��K���I�^�=����A�6�7�^�%���/�z��b��P��y�5syuL����e����C 9v-�I���o`3uD������UQ�]�s�"ЄDk��W��x��{+f���2���Ъd���{6�nc.�b�$�9�=���~��Z�T��!_XO��Wj���뙣�6��=yP�Iw��d���`�]�������m�Q���M�����b%�񟒎S�e�����+q>U���7�>�Skf)>��M����m?�}}��Ļ��r��4��uu	D�"\�/0
5�[���^�.���H�� �r�)I�=�����e�=��F4��v�ц��6n����*�.��b�1*����!}�^��<��L���*��Ǌ��	��ᾆ��?9I�_ӏ9���G��ut��o�����C�EN�0��>��\�+x3�5s8��P�>wǶ<��Ju`h*�)8���a>��5�*8ށ!Y��l!�x�бʼ�Я���]gos�y�p��wC�_j�N�����E�����6��u�����գkəC�� �-��,k�w��}�S�옦E��	��K�m�|��*:_���{ݝ׹�y4��=�a0_=K��0#���
��<��*t������E='��-i���ީ����}��eB\vDE�Y�W!��T��t1ϱ�O&�2x�u�u�4�w5�z�xX�yL�7�"@�ʐQ� A_x,;$-"1?@���T��m���;�.�[E,�k��v���YN�l�{	A/l�������+K��\��j�@0���EX�h\�Su]Q�moZf�^F�����R	O�V踌����<��{� ����J��'�8�Ż/x>L8���v:��3$�yޘm��Y�q`%���f:�����*�@��%�x�<�7�u�]"�h3O��Ҵ��,�˞sVf��ﺃ��w��!~���	�����'͂O����݉���r.M�ƕj��Q�D �ol�E!�Hi3�zu��p�'zr�)Ʃ�y!�)E�U��Kb��۟߾����|�� ���x Ҝx���� -gnDn�*�8d���0�^�TPl���v���ϻ�>�CO.�R�H	�g{ϰ2�0���m	߯o'=�	ߡ�H���
�n[W*�Q���#29���\�2]����i��}_����GZ�C�.��J��G�m
ݾ�M��@��>J�Az`��^�/�{m�Z�U�W@�JN8z͜a>���5�鶉@�����r����veRFj�
����G϶ja�v�-�!2�Z4)<#s�m1�^��xjkgk@Ŵ�~�\�A�_T.����6�[��S�i�j�Ib^�JKΒ��V��c��e4��7���G��*����:@|��C�'̘��@"o�z{�Ru�`�I�	����d+�Q�F�۶�\g^uo�3�~�t��cA@p.DG�z��e������K��EL�EҬ鼸�^2��&����l��r�¼��L�D��3�0��쾠B�y�>b��Tv���Y.��˰/iAb�?70�ڂߗݟ��"8F����rU�R���ؼ��9%���pb�0�=^jVc�v�0���..ZϧM�\�kXʝ���5�.�ȢF���<3��{�Y����/���������m��-�Y�R�����s�B�n�7?q�Άwf�p��nC�UUvsz�L�hM�чl)T�� (pR�`F
߹�y���sc�/������w��<x�{�V��{3[y���6
��B�(am�,��v7�t1����pK}c�=�6��x̀��k!�G��R݉�7h�C�[q�({켟z�������`|�K��g��k)Xp#�R3U��|P>�b��:!]z^�Nt�%��m"\}��]�)�Vt�+�T:�x���z1�X�7���9,���W1y����
CO KI� �b9��BӞU�Z�}C:�;=����I�;���=��yWw	-���{��f\���b,�GX�t��x.#���(}4�|�J��,�k���\�O�Q�q�}�/�j��ͻ��f�ʅ�Mg�l��ƸS�e����Z[T%U����9sZ�q��}��:��@�,:��P�%�^�'��6��<�ǬG4���6��`@�EwY��ѷ�?:� [I�s(V�σb47P*m�-���c�ޝ�C��t�G���o���7,(��ov�}A6��wɁL��pM���Z"f�eM^�S�H��ɣ�>}\�7�Ŭ�>7V�Y�b%�Ȉ�1�j����j�Aq@��E�1-�BWs[d0�UA`�m짷��To��pL��kȚria�U���ƘK���S3�`t�T�N>�[��s
U��/~�EQ]w��
�:b�naY�/ʩ��dgL���}�imNsYxLPB�����QaE�K)V��{t�]qN*]� {�G���<x���ǈ R�"/�����_��7���~`��Xk����Jҁ!�ey�L&
@��ð�c��1l��Z�y�6n�Ğ���Q|C���9��&��#rD�(�O���#�,���x��!�s��|j�۸���"ݷQ�u@!�Q�Bc�X�%�_�Qa�D�����ض1 �'�R!���}�Q�t�;��n�N�eD��һ�5�`�^�_�������.VW���v}���L��ή���.��^��[T6s��X3�N�ܐ���K�K��pY��n�\D�.ܢ�\S�f��m�D?��d���F	Lߢa�<��G�;���Ck�󧼪�?\�FŘ��G>���:��4(��a�i��:�l-��mxJ�z���,;�^5�<Bk�jn��d�.���۱Xkl/�mGuhh@�m v\�^|�-��������t4{=XU�������]��5��ȖȈh��-�尽��>�K�,�~Ѱ�o�8\Z�؈�7\������-��Ky����	x/��f,K�pp=�{g3�.���7D䡅b=�p`4� -F�V��+��^j�/Vɵe�)��y�y�dor".�i�j'�=�+�ݫ����풬��$k>�Uen#�����U]���4kL�>v,�^f�:(������轊��H�=�� l��=;7��6�����}w�ҧ<x�@�P$��ޔ���|9���O^�����gљf�Wt�v�!�r2�[Z��<��������ܭ�|w=,���8G����S�w�ӂ�q�2	+��CsP�jFCt�j�"����~�]�uս���p-�<��x�@���Cݽ0���f�ƨI��z.�F�j�*nz[^������={�e0�	�*��J86"|�L�g>�����o}�x؏vf�8����;��9`�>s�����T*�Ҩ���Qp�R�D�"���q�S����i績�h�^��n�C�tS Y:�d^�s�&=)86�	��qs6]�of��"vw4���#�mw-^`�y�p��e"�2"�Ȟ�4�`c1V�SM��~=��T�PE�29�)	9F�2ܞ�!65�d��$�^�GC��Au�(��O5�).G��U�AD����d��(�y���'���[�L$��*h �D?<��t�f<#�_RaU�'�Z�˔_�ky��մ�_�4Om�r�ܷF��OމH@܅j~A������Լ�a
x�:4���_.�������:�S^AuU�V��F�a4L��(j�	�O����i���%��-�+�@̛%LLb���{���ꣶ�� ��4��p�[����M��I�n�mn�ʻ��w�so�7�p\������}��^j�i��Ʊ�=�G��ן���{���z ��y�����Z�ᝲ�ө�7�Μ�@W��AC�i�!q�3����
�����ͅ=x5%2ⶍ���=p�ͼ�Mc�	t�v��$����a=�\�C��Ә#��,��)7��Ѳ�fj�b��ᄂ���wNt��T�?Mk�1�;޳C�|z�-A����q��B{��j�\�Hr3��(L3.y��;d�*,(bK�&|��L��鍅ܰ��cUl��Y=���E���i�2*,�^m"#2,��;����w������9�ݚ�ob����)��4��X�����E�i��
�["
�$�:euGr�+f7�xف�]go��i�)C�"�m�P��1:��a��yI�Ǯ�ܸ��.V�%��*vUD�;��Hc/n�a ��(!�WC���؂��8E^��)�,а��D�t3�=$��{.os{X�M�t2�H��D��%ĄȌF�'xJ�-{��[՟FH�3S�Y�����\ ��t�0=���[dD�G�k�u�>�^����'6�,T$�]�6s���qE�	0�+��9`�!V�z��a6�1l��ѹl-K5�7�{�AZ�/"�� ��N�E��`F�u{r���-�<|�Qw��fM����h�>@�f����e�$n�vyy���(�nh�4E�
btA����H��y���j�ŋ��n	���]s��|�;L��wW�4y��cxf��=�Zt����r���y��c;�v=�m������`�p�o�� ��{ኟv7��������4.;���'|��}���)ؓ�A����g�UF����.�G�	��Ϭ�O��4���|w8C���;��$�Eֹ����3�هb�gg���M9��&h���%3#&H~f�����2���ãW,ؓ�#�����VE؆�K��wոZ�纲��7Ӈ��[�r).�\y�T��e������0�~�>?-�<�n_��s�3;�d2�d̎>�ϟ
��hԺ�s�j�Z A��׃R����zBܘqǆ�����Uo\��pG����W������ިMB�~�D��\�9��P���$��*y������b�g{�f�(��~�^#�W�_7��{��se��Omv"�;I��������w"��\i��XC{/Ev8�k{Ⱥ.��ؔ'm1t{�	��"�ٳ��n�U�6��˼�/t��gQ�V��i����{n�u����2�--)��`a/�U�ڷ�\^�oR��kQ�IL��ea~'���5P���B['ײ�+�w]Y��j�-�Qԓ#3d��.����t(^�mm���"��)��+l��e!7hX���7K7�nR�2&Ϊ��|��{=���܁��b��^��Vp��vE��KL�¢�8�ץl{�eg/�O��V��i�/���2��>0�-��_=��&�y�Py�M�}���#٣}�g��sF�,_`�/{��<Gy��<&����a�`�ϼ=���va�S�����m��}č8��_%�z�T5�n�\�pq��Eۃ���<_z����m1*��+vV���������m��*rcU@.6�h_bJ�҄�:�:/�ʜV�.Tx��	�3',]7z#�5c%d�g��t�<��S��<��"�1�1�qm{��v��n��6${N�/U
��*�͕tk�|�o�)��)}(8�U����M���p���[�9J��_u��Tޔ�g����M�2���oI\\�l�8��#X7�/F���G]i�1�*rN��wz��;O�a�#t�ħv=�X���Gv�a�N��e~"Xjb	�d�7�>�Ipk@OVE�	��b������9�N�[�m�����޴bNI�/�}ϳ}=c[�w��K|N��ؗn�.Ʌ{�`BN�~I���yy��x<�}3RB�s�� �_�U/�c��ۦ�޻e�rHXv %�\QHִeس'�,�l�'��0�4��8�eF)��Fˣ�P�F �$ʤX�����C�u��(��r���֊)���F��.T�DRr4SQmmE4Q�s��������ǯ^�z������������b�)-�9���KQkZ�HV�b4LU|��d��yr֊�\A�c���>?O��ׯ^�=z���ǯ�������?���i("Ji�gb�R/�:���剫d���)�y�mDQMQT�%)G�RQUA\���UK�3��f�B�W6�
h*"��(�1ִS��\�>yȉ�"�q!K3Qglh�SCE%V$�E�"��$�-SESERQ^�r�"��ls`�����%U�i&j������DDT�Q5A\�o��-U$Qh��PMMDEU5ys�:&�5��UN�EE4��4W�IDG69"n^ێ�)���SQSM�ꨤ�����#4�Qq,QA$�"�(x��DK(��)���Zi�/p�W2�7svSڵN�v�(�����{`���u��e\~��by�xA|��CKn��7!�vp���;=� ��T0�P)0	�o^���\�����~����Ǐ�Ǐ���A>'�xz0}/~���g�<O��C�r���7�p|�I�����qC�Ot�N�xd\�.�eYg[][`���o�m�!���+�w0֑p:���������]�{�(�atH��������=�Ύ��1MԴ��9jw��*8$B��Lvo�O�OmN��y�x���{Em�0�Wl�z�Qi��(-����\Y?l��G����BI�^Ӟ�B�ֻ�ǯ_�Pg��N���PR�vTe�dkJGs��@��y�e���i��-c+��A�ͼ��p��9c�{��6D���"���V�Iw�uN0��Lo��UJ��Em�}�ΐ ��2�w�E���y�6��U���Gb���׉�O4i�{{%^�f)�;�r��=v���0	�\-9�BQk$^�G7!�w(�M���sl`���f*�AX�ۛ�����Gj�1B}y��lX�wm��`O�LK��X[��W��E�Uo�0Ԟj�9��;*PK�&�g��i�}��雅42$���a��2&[^�	�"�nL�L���Om	'h-�Mh�&.v{4Jcm���#r�O^�#��4��Hy�9\1��
R������o���1q��'ܴ�h=�]��3Y������v�
ֹ?tY�mg=c[uN9*�j�}n%e���K�I���MRը��z{��`?b@���<P�Ǐ)G���� f�ɺO�����}��U����ҘuiYa�9�a�s�}*mA��IP,G4*)�y3��Lc�v��=}��OQE�Π���|/�^8����!������됷��ư�N��+p�M��/�ez��>b�?4������L[_��ɏY���n���&�Q)��Y	bG>���zc/�_^�׫��5_Z%�B�("�Dɟ����֮ff��"\�˞
��X*��hu����{�| [4d:ٮ��Q�"��!<�^k�Q,���#�W<u�]!duYWFt�Q��"Nq�W�}�N�i��)]|t͕�����	���z�ܓ0��g�	E+���lc]P2��7{�O�rQ���%�Hc�Kh�3�g�R�%F��Ɍ�,?G�K�
�=��1M�Ǡ2~�y���{��%zX2��J|�}ٓ	��ҽ�Ms��_HE���}�Lg��SYsVi�x�$O�6:|�a��3	���G(;�^�����/���HgҨ7�<(95[�AkV�齻�ݿ����ץ�ga����{�9n5���F<�,E�6u���=�ӡ��2 uۗ�ua��!o�>x$��A_���5�[c�F:�>Z2�v�3�e��,w~����7���xZZpO�T��ؕnJכ�o�NR[E�^��'�0w VmZ�����ɞݾ�8�6m+���mv-'�bs�8�u'ق�?����(�Ǐ�iF"� >A���*�2���R6�-ݚ1�3�ϭ���D���V���9��',�H�ޓ��_z�.��ݜ����z�)�>zv�:�G��+�{��.4�����
�g��Y���ˣ^��9+���h����:i�" ������@��Ư+	��%N��`p<��K}��fm��]ҍ�)���͠����T(���	�b��`��:"��=��"]�CN��;V���`�5�g��t�Rs) W�G��s�>����Z���{}�}B+��yڼ
�yv-�S�`�EM�}3���Ji\��2���(=�jzb^)�Y6�j	>��\���^~�	B���m}�|I]ܫo���Y6]�er�ʒ�XM�k�� �]U��T$�Ơ����u��,�8�T܍���F�� �|���=�U��� �鮮`���A����`i��j�����8��NMs��s�:��ڄʅ�B��TXw�읝��(�L<�� ��&�s��P��&�Wu����

�-�����%9H�F���b��ȳ�u|��}��&� �#/����əۭH`R��g��TR�-Fu�ARS��*�O��e��1�����^��k��ɟ�|E9�{T���O��;h�����3��&����@�����C��y�@kP<ba��,(%��V33���r����}��������>$`y�����O-ҧ�0߁U��9!Ĉt�
�n3�q�Ll�]�0m�)��H:�WD���g��g�i�c��"Hn`@���0��P��Ђ淩ɎNK�.r�n�����h�/.k����ԁQ7 ܱ��k$�~�,��ϟ=/�!�{�-�y"z�S	�vI�waHS�g���*�g+�_:���-�J}P����J�n�L��w�J�'B{��h(ޜ�j��;q�um��q�غ�
:x��u�O�Vt��H(|P1��֩Z�� M�V�N�q��Ekd<�e����B�Kh^ص.)k��&Q{����q�\�\�.����]��M�������w<AZ~K�Q s��n%#�lN:F�P��z�-@�Z^Q��o,��x�7���
A?�G���0����v��TXQ1%��^�3ޡb�Gz8;���EOou�lW���yJQ�a��<�B�����/��l|~ܘlM%p�Q��+�����IsÁ�ؿ�7",�ڢ��c��$�,+��i�r����5�l:�ً���Y_A���g!��V&L�uٽ�_���z7<	����N��'�rWL��1���j7�[U�H�0��Dd�u���D���]0X��q��3R[����ۛb:������t �Wb�&v�/r�hN���ep=B�R��#�Qzss�?i��#0��ǂБD �A��H�F#�EP�C��$�w*���Y�������^����B�#^ii���.�RTX�">a6���הU;�Jh�,�9{�a�нCK'�_{�z�#�HZ���(1�W@�Rq���:��A���V��>��.ǂ��ӆ�J�-x�t��YC�O#^��M�԰��%6�2*��B�ؔr��|�odF�C6��T(�U�o�Y7����{�Lx
<C]r�j�7��x���(�	���@��F�:��-Ӟ���V� �e�U%)��^��k��m��^�ْ\�ķ3 ���52$�ޮ��mk7����GFr��<��0<��C!�\���9�y�W�%kJ��.�h�Y�1��t��ؓ�gH}�3���HD�a�~�t����g�/�,�If��^Mߣy5��B�=/^&-?5���P����<��}����k-D��^J�D�ff�@�#>��
�VG��t.Ǽ�Ҟ:�TE*o7s����-�7`=6����'�� �1{�b��8T��0��yä�%���v�2�a��R��%����T�~��N�"�t�WL�C�&o�[:��֣�X�;�b�S����ki�CN�w/B���g����n:Nu��os�O�<t��%��K{�yPZ�w��t���H T�7}v�� �۾�8��p���)�>�����ٽ>��Ͽ�w�?e�����AǏ�,L0`%]F쓆R�ƍ� �M ����'-H���<���Pj:z1��k�ۥ�nvU�U�����Y������J=@��� G}w�Ģ�Ⱦ���y�/�f8����(���|�C���������ܷ�_Nh�<hu�F5BP<�;h�m�҃��^�ڪ�1�>��0ٙ�t� ���ci�PKׇ|X�{��������Mv ��>(�C#�6����ҫ݊	����<�U<4��C���̾��5�ì�������趨r�Pdb����*�'繏/o�{s�G�_\���>��U[tM}~���M�L������g��PM�¾��u� �����ǂb�z�E��=A4.��#Q�I��ɩ<9R*�I~����k�9L{U�[9?	�Gjf�q��K��	u�+=r�Z��$�s2����>v��׃��,׵�G�όc�A�b�\����W#�^B��g��^����P�/����Xz���������%�mȢ���3f�D�ȸO��y
8!�/���e�L��K��C��R��[Œn���甉^���8;�b޻]u7}dm���H�XY����q��K�`宕��]�.}�{o��͘ �%�涫��¾���P��P�y�9����!�y6�c���V.���^f��;t�׿��{��~~~x�����0`�jI�H����s�R��� �uI>9��Xn�
T����&WP����^;��pa ��3�|R]�B�r ��L �E��}�|܎e/@����)Ӝ�m�L�m�G&3Zݒ���y��\���r����$F�˞%���]��/5�"���^�t���D�ۉst�����u� ��.(���A�H��z�D�t'�Q��4ky�TSU:gg�p�pT�����W^/M�3W%�{�48_����B�������!q����	k��V��E�[����\�˝�$gd���c�
��c�a#>�I���^����4A^ЁC��x��`UgL��3U��}L����6�[%@k	�[��"�&����ܵ kb���|��Է���M�\}�>O\/"��8L��A��v�@�K��bĹwtE���g�9�53WE觘;V;���I�Bp��?DǼ�k��l���"�t���l�~�q��r�O�C��',�ѭ�X�έ��dN߁�J>bX�/GdE�O�W-�AY,����/������J�"b�l3��&a�r�iSB�IIF�9W�0<u�H	[�<:�CݾHr�b���4Ų�`j�,�m�Uԡ�ܘ���hP�C&n�kdk-���n��U�p�d��w�ǭ�uGl��)�̞W.��
;T:mL����{\��@�'�߽�������f`��R[՜Ho����ٳ��,�)��%ǡ|c�	�"Z����"6lnX��J��ٺg�d�&����踆+��r�n2�*���P.zË�1"|����v㝚����ݛԒ���1q\�?��eտP�r�L	�C�Y𭚿E���vU������Y�o�S;H�@��������%��Ju~�h*�'b6q��r-��߶*Y\��ĭ��ݹ^���Z`rl!0�>��4�3{q�����f�������8�)i���w�s�V���PDƑa�_x8����0�Bȭ�v�ʞO~&)�urim4K�[�1�/�޾��
3��{��&T ��&<x�B�_*���$OW��ȏ��y@�zjb�Wj��[�,��Q{JJP2�����	���:~�<�|a�M����4�����;і�IQ`󣋧S�?����(*�+�a����ng��*�*i�&�*��ᦚ��e"�P�^��zW=�����z�[��ۨ�2#���9GoR�ب�4��vMᦞ�����6�>/�����<,�W뭦,����q%��s�D������cV����*��(���5�h+��j7q�é�{/E�Ep]F�b�͌�P.T5Z��2���7kDP][;�_ �
���D8�s6�<���'���<yǏEP�So6ac����1�)�^�h��f|��A��D����=�ݭ����kU� #5�m�hkq]�C��٭���&U�t�א*_H-@��j ��&	�x�ǀ�Tٴd��1$�a��ѩ'p�]^+2���4��s=�Bw��kꖤr��<�}�g�����/�3i�l��Ĵ᫧���]k����Ɔ@/_��r{�x'O��� �z2U&#<���mA�ReG��G��I1��\M^g:O�oF���-B�r�g��n��鋅?j���q�ߏ͠r����̋��;wK4��t��"�i�ʂ��0�*���i)9ށ�:�FLT9F)�5�(J��Y^�����_���QU5g�m8�a�"a&BehȔ��G(Q��s�=���M�n�=�ʧ���֔`p1m)ĵ�@DJ�ժ5��$�����6Ė|�Ӝd���=�}�D^��r�8� f(�e5"���ċ�̘	<�@"o�{�! ou�ݳ��sUk��Gؘ�EP�dWˢ�
WsP� y��C�B�8_gHv��3�k�iz��� =3(	����"��3W`JY����2"~�:��Y�g�B�퇨"�����k+�MU/���N�Q�-�P�(�D���o�uq+��[�0���7G,�2�
�9���Y�G;�/>D�{ǳ�yF�� Ս���/:y�O~����x�Ǐ ��V��o�H�ĜK��lV�aa*��0��.��C���HP�$R���[A��9%�[6��U���B��Ȝ��FH�3��'���\����İ�
�e�����X�9.^�>D��ڙ�����	�	�a�7�л%Q�X�ޞn�r`b|e%�~�5V�Le��޼�^�?O���t}'�*bN:��E��0w9z�7�V�w"#�ÅbL��b�r1�>��F�ܱN��[�3�,�D
d�*�&g�D�ٳ��t:�Ƨ��Z�l��ȿzZ�Tm^�u�g�L�;������L|�:s�%�@���t�>����;7��o����$���������~ugtO�~"�Da�C�B1\D?�a���o�tK�k�8���L��{�_�>��=!���o�t"�Š�i�Oz8c��"��D��B�Y�Q�uf�)-��ĳ�3x���y�����3B{���*�!���^�ܩ����'~�w��N���s���ZZx縲�+���z*�1�qF��Ƀ�<��f��$+	|Y�^R�SO����v-L/z9]Q�d�z]��d���ܰgT�E��2]H���]���Oq�=j�&�݊�����J%�
���yh���ѹ�ӎ�{m��`�����֭2�v&��a�1�fQ�q}�P�|�"0��b�]��v��@)��x��Om�����o�xn4�7���(�:h�\�0Y=�"��5�0v�A�A��>�ʁz�-�F�٭&r��n�*х��>�Jl�e��n��xM�{r��?��yQٗ{�:t�z����n��5�7Jx����V)��7���>fj��gbZF�y�o�נjk�ؖ����wv�`j����C+�6��X�f�w��O~�5�E�[�즫���F��kk�>�1�a\����]�;v]���V,�K�JDl1�jlw1�R;���q�w�k�7#��w4�=<�rg}�N^�oRl&b�ǅm/zy8�d�;Nx�[��%�+�������N4��g�$����]K��a��s�����P�l�e��6ЛR�T���315��mA�R�M�᪛�҅rZ�}��������غ�W¶&��=�2*Ԭ2+�Ϗ��=c���ۋ��tx�^,l��Z���K�N���7/xW����o[[�W�]��Xp�E��*6\"zNG�7ܶn¹!�d�d8�\;4�;GY9û�Au18�6��U�-�at�;BL�Z�%[o�9F�迩�?j������ҍf;�dr��^���*H����'ݪFs�9��J�ѫ�`���y숑�:�L ��2���@[����P��+�oVi�
��rp��%���k�@y	�+�� �����juVu�,S��:[�C�39�J�^p�#_7�<�ѐf�<��t�.�����\JY��nCu�Ԕ* ���Փ{c&��0�)��:ܼ�Em�t�Ƴd�+J�*�jy��]��	��Z�-t'��.�7�9 i���Kn�u��6��[u��<���Qw�J:���w��[�>��޼���m������=�|�R2L�������V�Q"�i�ݼ��ۊ�u�+��ڝɦ��g�����S�A-ܚ?$�fi`1���8�H��7`Tə�xX�4�j��6jk��e�fݵ����Y�{s��g��FrD�'��&4��#F��k���ƛ�[a�'0���sz�;�t���C����o����@�N&���N�F!�x����{�����G�[��J��X���)��x�y�u�W�:8#�HIma2�BJ{*.wۤN0�����zM3Ҟ��}���Z���yX����T�pUΫ8�o�g��f�$j����SR�{��o;������ �||A����1Z�E| �ƪ ������d�f-��b��Ǐ�_���ǯ�z���������}���?x�͘9h�����t�����&d�
������C�j�k��s��ׯ_��^�z��ׯ______����¯���5EE%W�cE�|69��1�Q4QSTBZ�41kh�D�TAQ�[LQ�s���5��P�Qz��E�ۻ�PPSE5D�b���(���()����b
���
����`�DZ4E�TT�C�[G6�*�i)�֭���1QSM��ES4��h�F�����+ĐO�9��&���p��&�(��@A�QE͈�����*=�S�(�b(����g����j���Ty�Psb""�_��)�m�@ �	����K��7~5��2�ɝ��V
�4>+e�VP&j�i��i9R�1�v�I���|�	�Rn7��ݭ�k��ƽ~~c�������� G��~ � ��Ӟ�]:ލ"�}����Τȧ{-�Xr�D\zeCz�B�+ڈ��L Ŗ�B���*�2���{�q�&3�8E �3Uj�� a���I1�v �\�Ҧ�f}�z�[�p�u6s�c/J�b_=�#V�1H����*���aMM+J*�._�
��ZS�t����Xݨ���˾��8oE�N��N�z%�%X��&��"}�B����~w�\u���N���U������JI �Q�|�C!���B{��k��C�J��Ø����zT��0檡Z���n�G��p��i�g�c�ٸ����Mǣ�9a�'�YH�Z^��m�S�\U�h{Z(o�Ǡ�Y�1�b�|�B��L  �U=v��U�e�O�g��l���ʈ7���v��v�[�ZmP�T%��#���r�!>�W�"u8�ywM����5.���i�Oڪ=��P؏n}|A��L� ς�#�k��R�U�_Jӑ�_H�,�CQ�;�n�^�����Q���(/h����k�'����qu �Ӎc�'�RU@�ʭ-4�۹�r�L6n�b�/uӲ���q�$�g������ϥ ��F�T�[��f;U䭡�|�7l��,X���[ ��Ub�'!ޕ��c�f�`j�M+K{��z��������1}�o�n#5c�z��&*}?a؀��x��<h��Y�3Iu�b\}lÞ�ᘹ�7�C>�S�~���&���{�Y|�!U�	3�C^�ԪjGh�ue��g-��(�6I�w0�C6��=��>��K�0�ZA0]���^�Ǽ�/����?0{*\������h�J9'�O����dJP<���}�ʔ���M>6}2�0�7�*݊���.��Y&�q=���Y]M6k���g�0	��8�K
Ȱ�,�+���k&�ۏx!u�x͝��lT��g�F�k���^�s��"d4�͗]�j~�IE�@��6�ڢ��'.�5E�`;�0�-�I�c�}�V�����P%�D	�r�n*a�8f(( X����ƻy�Fk}[s{��9 ]$�������>�u�	�Z4)X�E���3�q�?�/(���lG�L���m�i���_�b�\�"�p�V�mj��&%ؼ')t��JN.�8��sP��Q�y��/*��b�s��B�O�	����]F��E���)�NqM�)=�9ɧ���9.Mᢵm�z(ު߶���c	���3�t!���ȭ�Fw*y�����PD�㥥��7��t2��p!�0-\H3!�� �0sv��������u��G=�^���~E���Nw޻�#E�Of\+��(�M�(�������w�Rn㺒5go,��lj5Iߪ��V�_��i��LN���R�]�c:,9$�ߔ�+����?�<�=�)GOC*r�Nu�w\E��m��]�k���{���c���C���}�B@ꄨ���z��P/�.|��)a���rղ���cm�ok��Xw�5��Բ����ԥټ�<�:FLb ��Bg����g�����9�gw�r���-��.�*��]{�u�O��<eX�x,:��\�/ּ���c��P"&bO�==�z��fh�L-r
�^�K��njK�7����X��闇7��X!��tx�_+�K���ߐf�[��z'3����MWwSĮ��ΉS���w�/e�� ;�_�	P~a1��!��Z�~jo!�7x���|��xվy�R�]�]��;�v��wL�z"ϫ�YMOܥ(���S�
��do6��NS����3u�K�;9c:� ��x�v�tE����]s ��	�"����k�lp飻�`�����g�kl)���s�BP*5�fG'��s��\�(r5曍�M]1p��Ub8�c��]lY��m���p�����.#f����c�� ƽ��e�aT�p��8�.b�̵��������- d����xpnT�J�&���'q��pK����������?�E�<�.V8ʧ���ƉH����}���FP�-I���o�0�X�ۥRWL񞪹u�����j��v��m�k\Wi��]f�ZxQ�b˧X4f+4����e�X���������� f+����*L���|�%ė�{d��컦Ga��)ʭ�����x.�7����:ol�:?�8/�W֤�jӿ4$���Z�~�2k�4<�D��bS���8�y��BO\�=ʱDYF�k��`�eyM+J$!g�̘	<��|kݐ9�^g�(m,]�gݾ�N�[������Qm�q�t_ r���(�s�z��]�銨Y��vi���7U��r&��|�V�C���lj�&�|�{�'IuF~a�"l�3�R�=Jz�Vf?v��٦*2�}"M�0�{��b��$�]��r=Q�m\R�'��*��/W�����{p�_ɂ���̈��-;�Lx�i��B�F^�F��	P�u�9�N+W�&fʵ�G6�;�M�|��ca��C�7펿Tg��_�Sz}A�TwU��ܥk���N�c��g3W���:���AJ�C��O`i��x.��P�u3?B&�t�g�xCs��qƋ��{<�/ږ?�������&�P(���:9�xC�NyT��C�r�-�a�k٥1�ӓ>!a���ox��&��8L�YD.��#�����ǙH��2����:�$H���(5U�[��tȱ���7���!\�Y���wz�Rv�����M��DH<�J.���B�����J�f�����o���~~~��8�ť}��Z���9����=->�;+��tg�U�=A#�%�ȴD����q�E��Uݚ��<�]z]15�A�{kC�0��+<�WN���0�<X�`�MSUt)t�d@m�Z���+B�|�ͩ���}�"0wO���ϋ9�$&�-���ޯ5n
���΋��Y�4�xǢZ8>41	ƽŗ3���/w���ܷtM�0W�^uD3
}��EdH�}w~�{��Z�k<jca���E%`�6��/��#���Q��y�.���w�7UV��ZYq��"gP=�V�o�!ٜZ`�FV�������UN������=Z���cB��,��a�Mb[�HS�ņ�YMM+J>�$zD�˨=Ɓp�9<��*m�h�7#�x�>V�x���M<nEC��6lGd��.��!���|2�	]1��Q�s��z���iq�O��1����y�O��RO��&*�t�U䨰�c��s����s�OQݼv�fB��8�:[hLpm��4'��0�Ŵ����2����\��s������.���2�L�N�/͒�;���XL8��K˭�z�Vsw2�ʣ]��Qn�̢��`�@�cH�lk/�ٰ�'�pv'!�VOt{׏Fvs��7Xݙ�ߎ���j�9����j��f�/-n���=̳Hg�߽�����ʶ���;��:�t�y�N1�a|F�#B#丽T�I��"z��a��62o��Ƒ�p�<޾����`��X8��z���q>t�%�1Q5�o��[N�(��}.�i�,��|��`s��
��8��y��^w?Gު��6-"cഈ��o)����5ِ�O��bj�����^�����y�W�Ʋ�F����3�6���b�����r�0*fo��&s�>��3΀�d�7������a?H�5�>/�娽��"h:��g�I���m�c�#�oŘ�o��;��r��O9qw�Z����ص�}�b���aߕ_#h-^"��q�~���BO������f�:��'�ΈC�zx5�۞��8�wJ2>kM�9M����d�z���?!�#�l
����l��m����Ui�w��x�8C:b�T"��>�g�6���SZe*=�ڑ
�Q	en��1ƃVs���o��ٚ,#�[��JeI���qp�o��P-�6T��SZ���<sv���n�Ƿ[˜��-��|p��}Ǎ��l0\�R��_F���d�)*(,.�I��n������g� ��-�?7�&�m���É� a3���nc%l��Vd뤃��\6+Wg=���[]�f���fm������\���{�a@I!��<��yyy �V߾�2�\3<�$�P�#��4���k��I���jߩ|i˞��Q��4:����U�����2��!7�B�u'ҋ�d+�Y�=	�9s��d#�R�� T��vm���������	������!Yg��B�/�8�9{�+�]2��x;�LT��kj!�Ğ���.�f�%�	�����f&D�cG���ߗW�R-�2�ާk�J
'^�����:�{s�f'�tG�O>=�{�#k�5ʒT%F<E��>��z��f­�=5g.�j�B��՚���[%�bZ�����	E���t�5
JBlWѰAd&nrjx��w��*��:�3_1Ʃ9Rӡ-��5�qŖ`X%�Y�̪�ְ��l�ʣ11&�Jڌ�zo�)�'`��	>l`��nS����j��8�OJ素���Q�$�β�n��s�9y��tI�RǠ@�?���3_���r++����n�3_t�-�?�;��\�W[d�oVfJ�
P/��gR:A+��(��Qk�LڼH�n:�e��v4�]qئg�FX�e��@��i,lJ������}��sq�՘�n}��a�f�#7�k��U����2�r밮����|0p���T/Aڷ��OuŇЎ`�V�7r�[y����,NZ'3YUx�����7[���"�'��	��^q���z<=�öug�|{����ݯA�t=1��-���yw@���g��RՐ�Y~���7Hm��5N���N�
�y*Gs�0n&���TL��`����$���"�ō�.<�9,_�V���'�+�eP����6�?��&9U�y��m�WL\>�3�;��)�Qy�/�Ģ�yO��+��1{�X������R���PcbU�/�J�8z��Y�T�7G*󫮦�C�E3����r����S�Ѻ�a��b�2*�hRt�&^=��Jξ\�׵�ט��Zd�S������m!����x���:ͤAhyy�!�Qk#\jʞnY5��-��,��fT^$ư,��#X}9��QMM{��T��[Y尃j���Nt膪Ojn�Y��S9��j��l�'X\I~W����2)t|��$NXMq4+�#Hz��B���w#4�������P������U�C�,�`�aH7E2��\ۖ�p����Mu�����������Y'�t.=rD<��'��K�1i�b��t(~n�q-�>T$���.gѶkb�R�.�N�"n�6� ��;26�D'{��6�dؼ�˖��9m�臺�d�ڨ��znc�|�O6��.b)�N�$���:��n�b�o��s�铗 +G�bѲwv���7��=����olH�,C�o��F9��8V%t������������MϤ��2܇�G����B����?0֬FE��זF��*ϵ�r:{�o#)����4�&L��P\�|�	����>b�m{m�f����>�] ���x:b����Ϡ��,�����!��H�}����"��g��ʺ:8�`��,wd���@�[Ɨ�	O�^�1� ��j�{�g�38��E�)I����L�h�9�ށa�ɔ�iz]J�;l����b��������(�����ء(��xL*�[����i�����1r��V�f�[#������^�"��ӱm��y���Z����)����}�w��ZGF�(��&%U���6��/�F{�K�t��K�@�f���Q�M>YEtѭ�\�[����,�,G2�o�Ľ��ElY�ܓ^L6�E�&`�
�z�ً������U��͛ʆ�+������,���;~�)0�`M��"�Ogeh��=Y��z�~a3b\KT����B�Z��n����r(D�� {�4E���@L�wR��ҩC0��a�
.$Q����N�9�D���J��x�K���巔So�J�n=�r���lQ��;��z�砥�s�`�v�k}���A�����\��Z�D'p���*�=Ǖ�n=ï��^p�b�/O////���[��ܑ��MNc�q^�\M2/�!��K�N;4SRi(C-����M�lH�fMfq�u�����V�!���~�,��z%����E��f��K��0��׸���;�3����JG<�H)[����rL��}KH�lrC��RO�a1W���*,:�+nY�k��9���]����0G˕�����3�1���/;ja�ߙ���Dau��[�	��ㇷ[�M�ȫBګ�/�W��0��t��<�b�!"���Nнt*�>�5T0��l���v��R�3�T�w*/
�	@�w�%���B|�=��j����X4����gٟ��g=�@�-HB�������ǕϠ�H�ش���Tg������W�T
r��Wfo/�&�xb�]B͹�Ë>��Go��̈S��f��]K�s}��I�	��Z�#M��h�S���}Ck��K= �O3L) �\���k�[�l��WGd��=��h$ܠ�"�>
x�Oc��`&J��A���g��D��0�X��%���>@{��'�b�-�nڍ̖��{2��i6wxrM�%���X��w[t��x��T&�r�fvz)چwuV�~t�Ow<�p\���k(����X&�B�V֒��jip�^�vn�&�5��N���>�#"ᔟwxh{T.�Ncn�ۇ+���+)�(b{�4f�of���ꊇ
6=�V���� �$Y�cX3}�����s#�y�^��w{�q)�ק��k�ӛ��p�r�:Ap�Ŕq��%�)�2�����^8�{ ���0"���ԇ�m�P�Ȼd�cۖ��ř��xC4��8�V�0�N�i*6�Kz�Ǒ�p��EqL����Uo�>���2y��V�3��2�#"d �%�L��r����XE48�����#��*��Vh�����x�ϸl���.�����|����o�<専���C<�.�:��4	YBww[ot�O;d�p��]���m'�;8,{{W��g�}�3��R���:���:������Ь&-i��+�K-d���#;�i|)g����xe�0s���F��<��1V�)�c5���n�D�'Ӥp�7����i�D��C�G���\B�S^�Qm�0N����w�>�G�ݔ>ia�۷�� �Hbʔ�躎gӂ��B�����%m��\*�b�jLm晗-�$�T�Y^3S�E�� ���|;�a��ȥ��h��ȡE{�0X����2��~~O~m�H�|�ia�b�x�B���egbR���a��{�3�p̑a�Q�j�me�hf�d��G(�'b\[���}��rM��7��Y6s�����wd\U4��+��	�U�+NCS���/ows-�-V
���(�FoB4Ce�l$i��lc�!����Y�+PP���i�Ȁ��j�A�=�h<�F��y/��ˡ>|}��4(R/�Tsv]�?z�M#�>ػ��a��N��[V/�|�ή	��.MGf��ok�D8+W�[��ܜ�� �Y��̯5y��I�}�vi�|Z�δhL�P:ެ��[Y����n���,uX4W�%��,av���6mLw2N�Rഽk���z��巧��?er4h�N9��������2�7��vS�dC6�ϻ�f���f�k�P��>�
R�����Z�٣��ƹ~=�+�N����y�ǝ\��N�!e�Rc��'=��qz�����㹕�� n�ٽ5������:^�dшP�2�hu�z��8%�R�5[Fb��L�к�U�#�]�Env�9���Z/9b海7-*�qι���1�d�s�����{��G�r=Zz/.�3^�Au�;Uth͛L���fw�\1yq�b�au���CbV%)�C����z'��w���ԩ���H약��y�cC,,sQ4�f^�26: �c! ��A10ZD i�\j �pO2'�N(�Abq� Ę&JY�,�	e�^M 4�Id*���&�(J����lU��UMQDC�G�IS'7�x����?o_��\��ׯ^����������Ƨ���"����U����ۆ�T�Iu�""*����>���_��׮z��ׯ_______���~|
!����2W�cF�"�Rd'����4ST�T4Q11K�{�olLQ\�AQ\\��y�i51HPy�-5EX��i�b(9hb(���"�1�\�TrM�G��5�5DE��!5��*��I
{oR5��\j�ɣ[��X�.gU5�T�P��h|�[�r��( ���������Q��)��crϑ���j���9��h�0Z������������)���EQ5V�cgDE4SQEMDM�5䙨�)*��mEE;%j��*
���j"�.�痀DI� �"ø��p��A{0b*���߭��/��agr��Ib�D��\����Q�Eڥ��z�ӹF���j!o"�n�#���ʜ]vY��"!b�"ɔdi�A8�P�&��Ӟ�TTC�P.C&(g�����?�{ߍ�D��ٲu]�oD�g�m�>���n������ү~2�0\�Na�Bko6~̾�-Z���'J����F����t�&^����؞���l�j�`M!����������KDޘ��՚v_�X�6(�C2nj\�[��{X]��eO�+�ҡ�W��mT��uK��T�O��wY��4�|`��r��<ӥ��=4[�%�oՅP��G�Oۇ+��L��r��y�-�W(V�x(�~,B�R��~�������>���hȕR��aLNd�l���䶗��>�n϶��Ba� �	��8�Q�(p�[.�ZN�}g�'ʚ����w)�˛w����޼�9�� u���]���2��D�<��GAr��;��H��.�s����E��b	P��<�]�c�4t	����A�/�ʡ]�#1��(�]�Ô�B��4FH��7���g�8�
����Z���c�g��_�6��v� uBTa�)�Gmw�s9��V�}���Y�F�����;d���E�%�r.�
��qrPCV��x٨4�5W1*E���~��~�U�c�ܐ7���osS"w����k�ލ@���q�s�=�R������כ0������
>�D��p���b��s�ZF6�\��F��ձs�z�/6ɡ���7�2��	�9h�U�v��k7��=���yN�����������߳,��y���u��o�I��x��d㋲U���U�u�[ksK��N�zI�����Φ,x,>��qǪ`as��B�x6������^�¨�s��<��.1�M^�� �!on��l��Ltx�u��=s�eq��:P,c�={�e�獗��N+:�0���P�H��z�3��3�p0=��Qk��߯!�FFu�.��r���_gZ֯2�K���I���5�^6cˌ%1��g)�-v����К��� |�>2��*c���%qλ�b8�v�m#^)�3_�0$Z}� ���u̬ݮ�����1%����4��+�ƟfBOB�=�B9�O�6�w���L���H��vVWh��2θG0�pr\H��^�{��[B�|yHZ�]&��5���p�r�hw1���]�7�iS�c.aX�xB{|0L�ByOm���XO�xJm�d&B��c�[O<߶�k��~��я��w�Q,Z��@�6Q��GC� ԅDzC��k�1��l�)��sk��F&��q5�A�Fd!WXv�]F�	;i�>jq����_Q(OM�q�+����j%b�!}�8�#��gn��:�_�V��:��z�-ȇ:�}��`��?�'��i��uE,CR��:����{�?���Oׇ�����o�D����3��q���j���iX���2����w�P�o�6n��;{ ���Ju�x:�����Se$�0�����s	���0-����b�����,��X���!O����s��醣R���T��y���NZ��m|K}J�|^S������O���3�&���vR���K�&-?5���P��nszk �l�@��ല��$�E��m{����U~��N��Ɵ����5�Q�[�Uz#W�V��r�f�ʉ�i	=|�D�@��=9T"��O���ϧ�P~�9w\˙�h������ooV^��L��Edz�mj�@��T%�wR��h��>���2u%��\l�/�v�%<�-��;9��G3�,���܊��W�gp�m��FGp�Q0ϏP/���H��=��o7��D�"ٺ'ܺ�Q'��Q��jJ����L�uц��;��s�f^���l�)��=J�����y��:�����JK� �_Y���[�>9tҠs>��puX�\�M�/t����C��ʘ~�/t��W
%�b���+�֩�h?�E���~7�������}�(��3}c2�p��9�z���2�?��履������|ٞ�9*8Y��O;~�(�%B*�����<�t�*�xf���Y�s^���=7]�.�Ce��2�g��Ѩ�魸���.E�5ޕP6}#o+�۸-*�阪�< ���N4�j������	��ٓ>W���qS^�9��l����M� L2��������Nn
���OreCf��K�w�wAI�^�l_O��gTrQ���B��۹�Ԋ�y��.�i���i���y����$A]7�#�}�M^jH�t�Q*�$�P~k`���l�0�i�U��=�p��h)x�z@���P'O����ƥ��q��,��pө(�~���<��Ao�:�M\B�G]9f8lV����6�R˘qOQ��xe+�=|��7	�|�vʞ���[����*���m�S�3V:�dĜ�3�/'�#{�w�A���\�htcAv|��C6.��ɆE�QBSl\�àˠj#��m,
g�F�H�U�uN.GU��%�l0���8�M���q0��ZQl��/U�%�n��pUw���&t�R>��m�i�x�Q��1V+�K�1��D��&��z�cw�Y�꣱a����[�r��C���˛wƮ�+%�W���I2JE_�߀��zUZ�`����˖��l͜�3UW9 [���_���¹h�����ޓ+z�}����y��Q���.1�y�>�p�����>�x1ߘ�_VPG���0y��mס�й�g<2am����}�|ǇL:\k�~d�+NOb]@��D'u��鉻�����|bL�m�L��e_�G6�f��`�G7n���-�9�Oe��6��%������;�@�ྏ<%&U�&��c8H���jRѵ����k�G� ������9�`�BcϘ��w�n��Ǽze�U����nή�/�����Я%B=YK!{k��lvŅ߳S�7��gw�Kz�w4�%zE�F����EJ�$q�Ǯ>���2���T�T��iٻ5y��u��y!g�"��<z:T�>�[��
��f�g����QW��-MG��p	k/u�ksf%�X��g�P��p�Y��~c�a5mg��<�;Ry
h�觖�E�@粄���P#tģ�챊i-9}�bb�/�c�s��<l�r����O��Ll�������rt<�!J˝?FgM����R�Vc�8t���f���
6}'���^."qM
=���X�?��������7����Y,���)��>�ȑny+�!@���㞡�CT��TS惭��K�w��R�Iѭ�eh�s��������S*8t4�	�ýX�<������,����|ڊoi}���c����
ܧ=�Ǳ�0�O��#�����rQ��3��+x���nQ�%^�%�v�kb��veé᱕�팣��8�͇I k�ȩ��h���\�gr���g��i���&�m�,}
<�	��뀽�B^��Ǉ_ns^C���ge�n���"�'��5P�������[�(����31@p��r�ڑmB���S�S� �e���{�i�=�=q��'���"���}R]�_�M�1�'g�V�K�k>��T��A�_�t�6�}��xBtY][�y=��/t��W0ǽc͈*U�e�n�D��y�4+Z����I=ո��v�O�
7���w:_�
�]dj�Y��"ϼu��ٳL��:b~CqL��ӧ��znl�nRw�c�ℋ�E�D��	^w��=���<�3w9AM�;N�.��8�Nb8&���3IUT��{�5��?+��痗��U�}|f6�
<2���Gg�4�Myd�t$�:3ມ�AgǦ��N���oԒ�sR��Z����^�蜨Z��=����o'=E��|�E$�-zg�e����j@s0�ߦ:z|%"�/z;|ǫ�p� s�b�r  ��}m���sS�1mh�-��8���w��7�o�e�sd���֋��hm���Ϛ�O%P��ګL�	�xq�N�H^��1fN������Q*{�%~c�Z�R�\�]���n{�B��L���ǅ��Z��/63��u�bsf�p�9����F�IN�8"c������!̟K����!��kۙЪ���;�KRD��n�F�X���^���|7��*7����6ʟGv���VEm��۶X�m���� �zҾ��ϻ}nc��ڪ=��׷��ޘ�S(�?�٘ƈ١�p�e�*�.J�j;ZH�}����:�Q���zk�,�I�.-@"\dN!e�Q�d���3V���T������Isnm�� �4��KytoQ)�"a�Cg��!���V�4���<�o��x?��<X9d�ݙ&�v|�54��	���g����#�y�#�n�#$X5�^1k��":��G�r>���ǨGHm�j��熑l�$��X�/�Q1(�V���\q�'�_>�f!�gV���J�~�M��ps�覟���e؂)G�v�g�M-UyT�ȞoW�E yd�A�i��h���ћN��wuk��[�4�lW����n�A�"�@]��*�[��vqw?f��vn�^ٟ#u�-����~�����Y,��D/�]�~���A'�{��OMd�^�¸��c�c�IW�8ӛjn�@�j뱃'�O�2����MC'[�]�w]ԑ��S����xR�$���$\ә���l����3��Q�μ����\��آ���8ﰚR���B3>;w j�U�;�=v��b��{:ǁs�r�/xG��Kn�'���z�%RI�7�.�v.ٝ�w��a��Z-^S����F�ә����]�؇j{Vμ�p�]'��y�{2���&�V�Ԭ�N"�@���D2Ѓ��q��6fa��n�i��w�p)w���(��}u+��槆��ӈfy� q��xw�١����v���Y�W���l£�}�@//!��nw��V�ft�A*��o*������@\	�r/z�S�u$�\�����r3f�A�={וUx�@#1��U��`B�G@�P6�XD���}��E��dj=�˲W���l��V����凰�7�!�>T�+�.��U���>�dE���=�d�[�i�Ս g�k��l0]Ϣ*�M���ŕyg�fH�%ʓ��=���T���iA����Y�z�w=0b�q�
��d�;�%Ģ2�����.+&�=�/Ֆ�eP3��X]�GY�
��S������7�`�p��ʲ�V�ؗQ{�Ҵ|/oM��(�l�wG������]��9��3���rJ���;���]D�<04��!m��֚����u9t?r������d<���(nT�󩾴'4���C�=��-씄���(J�o����A[j�-��h�^�Y��2[(�";jn�)��jZפ�}���F2xg��$��''J:}��^NRUℸ��fk	�E	̋p˺����v��)�iyX�x.צ������{+�-���^�L��ht���o�g����)um���C{���=t��{�///{�@���n�b[}U��S"�����:|U!!.��Z���x�jIΪQ��=g�7 �0\8vf�u~��Z���.K(_!�(�48�z��-���Y�;gt��2n�X\F�
g!\M�2��f�h��Fh��5�yx���y�oir�̑�OL���!^���d������:�P*�M��~FV�4Bǽ�}��c��k��j�n��i+�(�=�0��_8�V�1�6��ݧv�=�a�T�L���|�Ng1�!��a�]GD�wU��2:F��f��{nx���.1�����1�l!��{�KŘs��s0�p]?gЖ�E����ڮ�ѧR}K�N�R��>g-m�kSs�都�yv��vC��C�=E\r����Vw)S���zW�:��m��>�l�	���8a���'�^[�,l���l�|3�p�I�n�Ɍ̷7D���F���wvz�q�Bf��'�H�SxN�b��N��j�ʶ�Q�q|�ZJa�T�Rm)��
nQ�s�,][;�읜l�N�t�[���l�Rq4�>)t��s{ 4zA�h���QBe�	�c:����2��n��.������;�ꮋ0��疪H�f'�x="���[�6�^_jh���S0�0Ty\����=gohh�U�I�u�X[�P��g����wY\�R�H��2���-��&�����{k/��Gd���|<�^�z���k�/V�|2���ݞ�+�{L�@'��JV��~��h���[�r��XJ�|N��ޓD������ϱD�D�;��0�r��bg��Ww�J��w�U��ޛ.	"瞹�;��w|�~�w�&���4�/`�Aʫ�gNz)xέ�ZJ���绲h'}OG|��.��Z<����6nwP��4��3$yw�Մ�{�h�jҥqH�S#3��F��]�[�� �ݚ�Q����
j����{��7����IN����f�����w�;��{�xއ7��)M�c�����n��K1n�!<O*+g�����!Чt��J�w�C�Uٍ*3fYG �1�aفm�^��#��K�g��)D���v���K�!t�bǹ��]<��vYn��si{�5��ʰM���)�̫�(��/i��L��.��A�U��n���n<w��� ��<��T��ɛzn`t��Ip�TͺI�g�ɟ���!Ӥ�����\���Yҁ�K�o���v�k�j^i���Zj��"��
i�nPiܚ��B�6��p�֠FX�����6=��J�����=QǴn��X�/m=��^fM�r�K֡1k'j<���t�e�A���{�|%�[����(f���N�w<�I���{��Y)o�`���D�	�"@��l����x}d�-��~�š3З�F�޻9]/������j�ͺdt�Wun��%��(R���X�G��
���lr�x��g�`L��{tHY��2l�����-���D�f빍�9�;����}���=7�#wth��Q�C���)���#���.;�^�GT@ɛ�9}�P��&@��s)�	��᜷�?k��f�aB�Cپp�c#�ʁ�,�Zf�;Yl�"T��׏�<�fMUn��6r��:��w�͡��TL�z9�.�٢�WAm��)��J�m�%j$�*#`](�����[ژƫR�wg.��k}�W+2��(�;'/QFE#R�l^w����(o��(m:%�^��s�u�^��L��P��M鸻G�$��C��<9����N�!���ųzo"p�w�q77�kNs�Xt�Йa�N�~�¨�&��Q@P�QUCC1E��D�h5l�"6Ƕ(��9�������Y�ׯ^�}}}}}}���|>�T|��e�T���U͆J`�)��3PETTA��������z�����z��������ׯ���S��A�G&��������
��cr�[��0bf�Z���)bhd�Ӫj�ӂi(��rP�V�Ickh��o�6��Ĕ�itQ�5M���pQZ�4�M"�ÇB�nmk�\ű��
��_O3�ѣ[b�N1��1Z��% m�'�rk�b����AF�)�ѧZ
&�kmA�A�*��f*���m>ت �<�ָ����U5;KcMS�m:�m5�QV�<�(�T���:
Jǜ�Cͩ9h�[1x�(��4U���cV�kE���I�9%'#F�����(����/��:`87���s��
�|��j{�]�מ��ttN��_M��󚊼�w5jە�v�i�;�ظm����^@///�{(����Ļ�W�G�K���ꉇ.ށ�5Hp�p�������]ΐ�'��fq����H���Vh�c�p,��U�b���W�c�sL-����~MHz_�&L�A�&;��6�z+�@�]�.�F_��m0�.�¬o�uJ'gRo#����1��YN��ϡs�X��T-02�'q΁`=j��i����<�]��FB��+�U�wf�'�G�i����-���z��P�MC�9P���z;��m�G�\}Ͷ`�ڭ;��ge���|�;V�����/b�eg�;��Ʈ�α{|�Oi��p�I�.���t�m��������R�Ž}�B]����NzQ<�BJ�>���)��R��.�6e��Ow�{5�N{���4o�e�S�er�+�Ƃ��TK)��\�}`�����_(ާ��ۊ����نb�V���+�n�zN#��	�e��_OnRY��I�9^ݻ*Z��-�ב%��*��V�(�ױ"rq���\VJ(��4�_a�jf=/)��qYz�D���Y��a��B���/~yy�W5g[�$�� 9K����=\Z7g���^n�^�,��[�Y��2`�A�;�Y0Y6�j��@~VW9�N}�����Sr�O���Zl�ҡ����1���j�G���B+��@G�����Ƚ�[^���5s��;�mt�L�q�`�}�=����k����%��Ҫ��fn�^q~�I���9��*_t��S[#}�t}��w�A�������b��Ნ�-�C��|YG�ʺ�4�#��bf)i?:�7�Kf�}�W���KN�v��$n@y�"��������g��8ڶ�=���=�v�f{JY�������</im�f����&|H.VW�C�;�+������+�EH�w����*o��i�/_�o�&�2�G\�쮾��1j�|%�YU�Cf��ɱ�CJ��˟��פ��Ӡ���ß�՘äk�v�M�R��;��ӑyՠ]a�*��p�9��J���l3��d���0��t }��o�7z���huI {{�i=�������񌮶w��s�q/��ŹV�;�j]��;
��\1���z�;=ȔU��m�|�H����yyy{�T�]7�I�}�݇d�;����+xwEy#�9��ͺ�j�����6���w�Ww[���/yP����%>��qָ��5ގ�bCd�¼���rꖜ���RA�atya�����)]���U�/�����:_2���ɤ�h-�<x�Qջ'���0ו�iF���U)�o�򥨆ȬĠ�^��ಠm���P=p��8��{�;��D��{��,k�m��³�����=�M,�Z !��6��ƌB�>�ۋ�8{y��z�i�	R&��ag>vܪ�s�=w�<퇳L\��E��'ts]�c"�V��6�bz�3IwN�b�9mhf��r�ܡL�6'�I�����!���{j�n��rR��Ѥ��������V�견�A�՝^#��q�8N_k2�ҩ�-�ݔ�0oM��}_�^A���D��hBӕ���o��Ф���1,��j�5�>]gszz�v_N;rv�Q���ry��}Ϫ^��L�����Q�ق�����B+J�h�X܇�ӗ��Jԩס�6���ˁ,�GV���-W���ʏ��=.���û[�����ꏳ%��ؚ��D��`|��uGb4 Za]ٞ�W���%�����r��	�іF�@��:�p8�K���N�����i�"���>�H�c�h�,�\:�s����gé�{!���`�Ϭz*�Q}���H�{��Ci��ww���c~q��迗sG��mP���ြ]J9�\�d�n����S^������W����T�
���6Vb�,Z�w�oT>�����}���窕B-t���e�XnC���{�d_N���qCf�D�Oh���=N��Ja n��8�~���P,C��#���3���;��aT8irdss�
:���h�Zg�n������x&�>��'����}�ǅ�H{��ֆ=��2_��.y��䚯>ZܧYْ.���!7��Ӽïa�6�]��o�q�I�;�Rn���m��5әܿ!�C��MP9�Eaĝ�n櫲�?*�<��^Έ�?23���}�i��b�\�;��%]����ӫ��_g��Ո��kmy<������ooOaj,]r��:8�0�2L�G�sۜ�~_��ۧ5�l�����cXÀH�����?�����l���^�Q���f�)�-ۜ�VMz�\�Y�˥�|zz|�2v�bO���f]���2ǂޟ9��hJ1�W�����qN�sܽ��W��$3.f%�g��ٵ-���6������wKq2�u��i��ſf����Tt��H��v�e�pFl0�`�H��"��.j�(Z�'�b�|v�O[����H�����)�{���/�1�_BwP��*��'f��DU]��ͳ�ې�;���w���{�t��<v���80��/� Ԫ��os'/WV՘�my|V��q� �rI��=zm��2sPub��NO-���W1�����*U�N��$�"H�[ 8*ٙ����f|ء\�_uі��r>x�Z3�,1S���{���g��yT?���/+wg&iFh|ug�e�2�-�E(�`�o��]Ϫ@���Z���0�AS�c�������jg�e-N�A�������e|�	Q�;Lʭ��*��T�::�9b4��\�,�����8r0@��/&��%,�����bp��	�It�WB�h�|�й�8.�s�:���B���x��j0|>���}Q]�Вy�uF���fy��ԋ�s��M��1���򴧳)ka���ך3=Zp���C7Bңܑ�eW�+�-���S8}V���Y6+7ďh���|����$���G��V���4�06ҍY #BUA��>�٬�,��>��99b��k5�����^��\D�2;�%la*[&I%
z�М�V���|[C�m��c���{�\�jx*�<[}�+��i.��[-"o����k�ѩjOM��e'�����؃��ղ/��i����T�|կ[��'jI����$=�<MS����m��d?�;��ۼn�Kix�([F���E�^oF�w�]�����>�ϡW�o�	�y�|e��~����I�o��s���d���G|n�[�3o��O��d2�ed�Yܝ���`��=p�Ǣ�g���`�pw������]�so"Q��lø9�X��.��W�_���r1LD����r�$gs��i�3쎒L׻�S-Z��i�r����'ńE�]B'U^�]��s
QbP!��׼P�
&���{�ڽ�����ى����m5�EX/��b9��8Q�T��"bϪ���/Ҕ$�0����yyy0.Yz��%�5l9�R��y������5���Ԉ�a|���W�����ݫ�L�椫j��<���]�pAP0�Y�j�p��ucy�޹�`wt9�������k���d��c㢔�S��`hWB��EX����Y֗	(�Qxugvu���j�%'K�FEe)��9����(![�E�-�ç����=��m���"t�C�%A#�9��]2�oz�,�����b��<���(��	��m�.(���A�mP]�74�Y*�{q��������U�a�'� V�p6�Ɖ�i#)ъȻ竨x�oV��μ�����v�O~�]C����pH�n��(�7:��یk4��������5O�t�}�� �%�k�
w�{��^�m��ɽ��<���|ֺ�-���˨p���� ��0B�����sG�ӌN����&0�術p�V�KY�{,�t�3䨤��_G��⧦6OT�v�:8�+	���$i�z�>�(�{m�-)�ʡX/�l7||����-����.`�%h�2XhޡT�4F6��S�(p�� �@?����;��w�OWn� mq�2��c���!l���Y�Lo�gǧS�w;f�0�G��a�r�L��lI���G��B��;;��������-Ja8�{�osFb3�5W7uN���x>�����ʡ�����--c"o�1 ��� �"; V�*~����{�[.==�N�7f^'9)��S>h�8.>�<�@��@gZ[91�t)5��ri��As1�sȓ���~���|��䓜�R�Ťm���ԩ�ݜ��;�f��v��Lm�tr$� tQ��`�FC:4^?����:E�`�!n�87�N���-�]D����T|��x+�~L���ո�|'o�d5G��m����d��o�*!%�+)��Z��>e��7���<q`�-Uqh�Mw%��wEIC�*$��yP׸�-w��h#=B�X���r�뾛��Zjv�3�<F4�k��7v7p���Ew\�1�H\'�cVn�7���$��;�/�{���T^�1���[�3���(��:0;�Z+j_!,���0M�cX����g�S�Tܳ(~�� ������f�oʺ��ˏ�%d�(1밽A.�O� =ü<`��ٜ��8�;�h�}�E��9���P&�xH�O�&��G���&D=U�Zn� W���7��մ|ر+e�x2�6e���[��-�J竭R��b7OE�n�q��D�݂M�$U�J���B�]���d��b}�y{V�71
��p�%�T/�G\�=�m@)Z_OG4b�m��̠��(��k&~�У��)κ�۽p�w�A�GB]��,���v�u&v�+k��\�.O�럼'�~WO˪�������ߟ�P���![��=�������O�Q+�F	�f+�\¯�
��v)���c�t癵�
l~�y<{^�-�Ƕ<�0��k�P���
'e4D���W=�Js�������>Xc������J�8㻢�٣c<���t�qN��ɮH������t*�t�1"2�v܄�(m�q���[�ԫH���`�VVnfQ�zw�2�5(0�_�����}������3�{��t9�G{�E�5��0㫆� o�;��>ٹ�s��.څ�=�dx���9��1�&��{��?���'OR���W�z�%myd��2@�A�&;��N�s{����0�\k����.�E�ѹ>����Xy�Ycy�7o=ކ~�I�K.������+\�0��0��q5$�T������L�y"�=%0�S�/2=�y���P��l�etHm���R��5k�vl(w@�g2^�9^ٍ�Y�:g6�Wwou��5 ����/-M�9��΅8��?G�tn:u+��VOu�J�L/#�eR�hʯB7 ���әl��~IM�cD��fgkw����B=Zt���λI�%:n�Y;]]֧궵��y��z�:u�+\�:7\��2:J&5.a*dω%+4��&��A52�V��vd��}#\nKc�>�P+�F��H�+aӫf�f�@��O>��z�6ǚ�B|�Ljپ�>�[�@8����tz��N�x��U4�>�(U��m!���s1!�Ի|�W1�ov8�jj�ey��s�gW>�9����Eݏc+��ћ�<h�Z��������e<�?���w)7���n����X�0w�+�9����.�ZÆ�u����E���W�_\~�ݾO���K�,�Y� ��{Αe�}����vL�4��o�hǑ��b�f��sٛy�<`�J���,��U������iYu܃$ލ�5,�OfvZ���[f��똩�]�^f��
�|���C�z�W��������s�1Mu��_����v�Ь�*���5�/(�ޱ��Ϋ��8�vjiiF(Nf�)=��F�

h�ͫ|����7y�K�sK�a�FN���F���ר��hw��g�	Ѿ9�=��B{\��OX%�g��`��	ίxn��t�;n礙���H܇	�Wj�H`[�5F�0ܮڦh�����1|X��j r]NV#~ٍ�#�{2�x\HR�9Ȼ_P�ٌV�\y�39�ŻǠ���2���a�����G����'�걪�@X�Mc��Vu���1_	��/V0xE`�e>��z�F�Ա�Yw�����V�-�9^ה� K�L0Z1W�u� ^�L}����wp���6�:����:rf���"[��T�Q�u4+�/l�nVx��ִ���p�c+x�:m,�h�]L��$#q䧩G![����eӇ֢��7�
ۍ7&�"��I�h�mk��?�U�mb���U}���M5��Ҩ�;�/�r���LB^YJ��5��=,���G�F�+u��Qޜե[Cb/Ҏ�s&:���
cx̦�k�BZ�m�*�rⲱ�|��(c^���Y�<�������S��oN���m���Τ��h��Z�����up��>��=�Kݾ�ħP���'r���.׾ѷ����zez�5�P��	]�{zzh&�=����;���,�o����WɎ�%i/�G�׃��>�I��t/ٓ@\b�p3�i�s��\����v>;�G��ݱ!b���I���>9B���<T�C�� �<��*�_�ndΔ�$p;J�52R3��V�δ�h��=D�r�;ރ`�}і�zDx_{�����Ѱ�ڎ,�=ȄD*����P�ͷ�R��C�˾w�b�-�νbp5�ja�ԕ��R�ﺁ��}G�&-�]K�[�l�.�����!�ڛ*i�6�>͞�x3�/J�Y�G��U���b=��h�/��˹��QD�D����VR�u����c���G��Iv�׽��G	w�3q�rשSq'��
�黫3#��I'����fC޵(Lm��#�@�ɨ
f�˥\��&D�;($3;�vkĝ˝��
��P�X:X�p�U��h�����eʭ����漉�� H ��
l @�b�lH�?�?%ZZg,d����醔ca�"���-��"�o��pb)��&�w8��|d�O�9q�6�Q�b���c�sb��||x���?o_�ףׯ^�z������������
~n�3��Xӵm�-��9�V���Wqˆ��Ǜ��Z�A~<x�������ףׯ^�z����������~G��v֓g٪�AF���AM8ݹDslTy����s�z�o6+l���;�18��b9i�j��֊m�qᠶ	ֵ�Ӫi����GX��gNӽ�+�Z�ⵝ1i��VƦ"��F�R֔�Zmj���r60QZӫ�\ع0�ڭ��1���G*4�s���������(9��y�nsN$�UV��Y+nsj�Mcb�ѭc�9'ˇ5TΣ#`�;Z���4�c�ݚKs�E�Eh�h���ZC@E���ι��ϲNsS��xSr�V�T[Z-�փs��F��QÂd�0��o6�AKL~T��G��S�%��������݋#i��F������w��@x���/i\t��k�Z�9{8��'�W���Ć܆�$A�]�����z]�`���ܸ�{��o���"GWG�]iEW'��3����c��+��hz�ϱ�����s�xt�"��U�H����q�{�h6�|i�q��oV�J`�)��^^��#� ��=!�iWq[A"jiS���R}���O�"7L\��N)N$�2�?�*}.��gB�lVyFx�I�T��<�MdFI��1R�0��8c?�I�˄*l�壤�L��v3�a	�zß�z�9VfJBP�^WXg�����L�e�-��d�u�<d�u֪R��o^���W�77�`�#b�O�0���͸����ʿX�^a�d�K]Þ�]��}9X�y��p����+���VN�����K8��.ħ�u�6羳���	�a}v|!8���������6x�T8ٴ���D�隘.�^7o�w4�P��=�ϕ׵U�@}N�-��\!�j�mP]���<5�i���T�g䁻FY���ڈ���9��b0����*��p�<���t8N�3���r-���-�x2*�)z;x���kl٧d]��;����5i�[��C��/����F�EH�&Cc��� ���Ml�W���_TGe��/8�mR@��:���:��϶�`q&����[��묪}��k;gV���^�f��^���xp�����{lͫ����4*��=�OÇ��Om���=��h}B:��l�	hݝ&�wv�y8M�<h6�'��!�=���Bޖ`n�^����q�K�p'y�e�3B	.Vl,���T�w7a�q��je����Gq%�WW|�.�lV����'���	=��F���*3bĩ�&�NQ�7�6���`fN�o{9��P�؈�G5���K���1�ֺ��NVw�^ұ�Mng@����pQ��kG�*�z�/��y�Kך.#Kݛ��t���/h��`B�~�k��d\���y��'�U�ƒ�z�}�s��GLw�+��C��>����+��F>q��B	�qu�tO�ޠə�Ne�����R�^֛�篊��`m�RF+m�?h@]D��nV�[��}�E���ڛ0���y��U{��2E����v����}3n�5�nMW�m���03�c{S���ɕ"t��yWLKP=7��N��:l�RE� Yh��{�[s�c��i��m1��_P0Pk|B[z2�J[\{���g�4z��Q��/=ǣ;�����k��|��z��o6�zc�F�������T+.,�|la��
�'�.�21�7-G�0��;�n����M+u&@g�@z�����V{3��C{��>f��P�m���z��!�D3<^Y~��*��ZІ[�DI���j��Ϡs���}̜yO�gNn��u^Y�\�#�.�o^�uWJ.�H��5O��r�H�ȑkؓ�$f�{n�3{v��G��D6M��Fے*ۥHH����r�-,�Z+y�r�GX�OK�N��J��F�����gJ|����g-碫�;�W0|���j~	l��y�_�����]��}�/H��k�ը�����s~��1�|���yD�I���R����M����� 3�2��r}>�y�#�̽|�;o1Z�]��ۯr�����*�%}��v���/+���o^�Z��Y<��S���uԟm�Cyy��eѾ��=��37��g��g�X����D�N�t4�x����3����Lz^�	gjw9��f*:
��Q1�yl���<7�@^3[3�~RO��K3O[�Viyې8���{�XUǧlu8�B��W�8��߹N�\T��E��p�a�D�O��Q)��ђ����XM��/1�ɓ� [����G��s��C������_0t�rA1�W^h|�ɉ�d�;��^S�@�?���_��uF�h��m��m�ݞD� ���g�~�I�s��O���	��n��OG�ac= +w4%�W�F�D���B/�#dO�wX�iyk%�XQ���o���{W�G.�Gy}�i�+u�+(��yUy��n�b�3J����}yjni̍�p�=_u�i���k:��<��Ss79]�+FF���Tәq�����DL�o�*��X?���x�-��y����b�dz����rb�v]Y+n�(�e��|S"U��5)���C���e��>&�18O7��l˺�r���8���wj�(�
���QM��8��u���!�eU��抹�������1v��m������������[��]�*v\�Ⱥճ���zP'��J;��K�=�S�ˇuW��=sl����\��0T
�'m`��޹��6�=z��wR���$�>m��O������Ms�r].�q�W���Fk|��l�^έ�7�k�itOc�jP�y�w"���'ѫf�
�G�q��.�/���9�A���&���Z_R3��p�ҝ�6C�ʢ���M��\�n��sں�eQ�%^tH'vM�2ԇ�Z oUn�
�q��5K���up�0Y����b![��o�>�y�:_t��f�9�mC>j���j�^wF��y��k��;��\�|��ܧh�^F�+����Y��g>��鞝�kP�!�13�:�}�0ǅa|��z���;�OE�zܽ���z7�,���{E��g�;�#��D����[x�0w�u����J.�۬���e����|�+|�ck /G�j�Sn�b���{!�s����^<��r�>T��k��h�ݲ�?nVg����)=&�dM�W��,��m��{FM�|Q��>Q,����So/Fʍ*]�o�u
�yy����굴�,��O�$Q�y��D��9�й�Z�N���+��/7��C��5���ĻϽ\7�~0+)��/NIV:Ҡ�L�N��Żk��G/ �D�\t�ޤ���i*H�f��t�1�z�e��R;[�L=֙:2��`S�^�z2=,ǒ�zHW��dR� ���5�(Uvۯ5��V�zF��zeߤ ��O�B��(�Y!��5�]��=�r#��w�LT���ۘ�F�K�s���[8�S�EH�� _&�bñ��XX�<�-q�ɴ��5���t\|YJH�e����r�l��ન�[���£ln��-7+��l����.#`��ͽ��6c��t�S�B�y�i��|��Yx��T���sZZ�$�.P-���#�T�7Z��^���Mlb���P�[>���V����:�2��Ս}��X5��Oo	��	_mU����p^�����c#ם�ogv,Wж�Ǳ*������7d��\��:�9��=��e3�}�$j��]�>�rgk̄*�]Y�v�ne�	�# 	�b9#s��
cw����ѻX�<���;U�{���-����G+a�@s�b��.�i�����5��y��kn�ף���H��+&<~��
p��{ݖ���9�V��4���F\ݹ���C��|��]TLA�`|�~��rϹ�x�W�
n{�md���F���SK<>�t'������F0���1˲���W{9{Ӡ\�(��<��s;�f���5I(M�=�c�f"�c�s��4��f6�����vC�@4W��Fe���?�`��$F�k嶎�ع��6[��z�v�MK�8l@R��&��f���|GH*�vN��Nv#�����_P>������/�@O�����'�v�w���2ʛ�2�[������MORӍ'�*%וjgň0�R&�{bg-:��/7=�"��$�����<��u�t���8@�ޠ"Ns�2a}x?�_�y�{��hW!�4e~ڻ����Z�X��qI
��zfK=�6���t�j�_6ٽ��u �MHe�b�Ӏ\Ǧ*��;&���%��z�[���7��>BԟA����ĭZ6�(�j^+E;�}?Oٜۜ�8OFlN�XlD��.%	�L���v���$���E�Og��ڗ{���9}^�!��۰�^�9�V7J��At�B��:�w@q9+�>%!�l�o338���7+�G���Q�\[6���jK*�>��R�C+z��G:��d���G'��t̰]"�lգ]���f���\Y�8�s�M�%�%ԅ���p�d>��A[��e�t,��3&���9�8�ֳz7��@�<P�9պ��VY����򟏟5�ٖͭ7j�o���+�y%���]g�Z�=�IWG�V��^��sR��0ۊup���D�ʼ�����*�6Q�Է�ӛ�A��ޯH�Xh�lB�İIzC���ީ���h�R��a"���>�H��A�&=�!�u�{���ձ2w��q�kѴ3���=<*5h�?<����q}�~����Mgl�t�lW�v�c*Y�T�Tk����k^����"�V�.i�R!U�،�������x�ve��~&�1a;�W����a.����Z�yMco�<��6�K

ff�r��Ŀu�u�	�%���f�5���ef��t�:�w��AM���~����
���zt4DF8<hEG���E�;�b<��zJDMOW�2�����f�w5��g_]���"	p�i�״�ݞ��<ý�f�q��okw<���#=<æ^��F�';�0�iIKi���Ĺ�lB���Q���K$$�7�W��w���u������IsՁm܊�r�n	.�����z�T�}eN1���H�\8����,���xJCɌ��qd���+���a�4}�馨
�.90�
�#o���ISu��I�d�����J~��ؗ� �D+]W*��V�T��-u����{���Pl�+;dw_O���5�H�G��Z���"�M���Q����{��Q5*b���臭^6�s|��u�R�C��c`W�TO\��=�-�⟁'�Q�ܗ�pYS#�tPk�N�] �W�m_Ͽ���\ט�H����SZ)�](���W%֌��n�����;��f@NȮ�LQ�}[��S�#�o0'�&L{���d�	mI`���J挦ٝ���,6��� �����κ{�0���u�����q'k�{�7��ts^��q=��b��#1ϰ�>�u{�-�&�M��m�莾3X�噟�2I��*S�>j��]��	G�Q�i2��t��lY��K��w�s�<��.���9�7��cڙ��xm�p�b��g�JbM�fl,��A�M=~!��y�j�@�E��C�P�A�QU[��Trw��=}���\VZt�RO7X�����*��Uz5�0�1�cA��=Ѻ�|��ɌW��sy�n��R8���cb��4���c��'����Y[}��$jv��aH����n�$p��N����^,Eh�����&K��ݏ=��̎�dV�3�ɄB��f��釡=�������=z}��N}�)G���"��c݁����y'���1覩��G����'���Z:�%}ȀK��W��ϨY�����Ka�5��Q�h� ���rpZ�)T������[e'�z��J]N�y��2�,ƓV4��M�`�[t����]����OMq%�}D��$�M�,'�t��M�V����縮������2�VF��	{=;βԖ/?=�a�q��@b��ʦ`�
��7-�bˌX�z𜷲��dY�M�<���c�����zO�Ua�l~�t!�����>���t��l����!k��c�J!�����ͧ�2tH8��N�7�o5��nL�!�z�+�xE��/�!@<C���.�qrޭ,�Ü�S��!Y��������x��<�p.�|"��MJ�Z�"�2B��݇+r�75`��v\�5~��Rj ���m��!��I����d�Z����V9��)�c��ࡺ����W&e]>���(��1���<dN��W;Ox�r��ⲳ��묄E��C�Fc�~P�.;6N�Aj5ק\NoT��D��ƺ9;l⻄ziV�M��\��zѱJ�$��X4�p����b����`W�a���y��E�[��������S�-!�3]�[9^-@��kW�g:W�#8&��Crw���L+��7���;z��5�r�9�CF�kgC��//����R&n�մSwV% ����q�1��YkuT	��% ��Bz�����۹���g?��-OO�F3q�J�8����u�0ɘ�#����n�w0���`�q��L��Cy�`šРW�L����j��r��,dv��'�1ԅ������X��sO6�f�)X4�j�R4��E�,��t���}YBy�X6�.�_(x ��^��k7l(p���V�S�Ũ򹂏J��=b�NG�~��\�\-v)��T��#Vf�+�tw���w��ǎ��ꃀؘ��w��f�[��a�f� ��� ��E�y�jwu�E�jv�M�:�u���͹4hf\�ۋ����(O;���.Z�/�q%L���xQ�� ����ɺs�:�o�zm�@?Yo��T�^�� V���5�d7��s`��>�9z#�`����~pd��J��3"����і�7GV��"�ܗ������+�и:� ��M%���:cD�����B֠66�O�ԭͰ�J�a)�-�{�'E��޽[�n��h�=a[��]�c#o&�R߷�w"S���V����o-e�5�D��Co9�=�h��Ь�,CC�/P��{==�@o-��SkN���ì�z2i;�o��3���ԃ>Z)���ps��ն��Q��I���=�U,�ܴ�A�JZR�7�[�죳;h��w0(p���P)?�RunL��x����ie=����Ʒ���wK�OXd�|��0t�����Ĩffh@��	���wF&�:S��[��{�E\���m�o��e�9Ͷ/�y��1���>'5p�&j����������~?�����ׯ^�}}}}}}z����km��a�����`���[mm���h�%j�1[TPQc��_��������ׯ^�������z���}�9��p&���m��Z1m��Z��s9�_8c�'�.M��V����E�֍�ƹc��4bB�v1����dМ��y%ͯcǰp���x�1��(��܌m�b���A��4klڸ^s&嫄i�J%�����[�\"d�h��9�U[c�b�m��i����D\�̀�9h�c��4�Ak4m�r75Tlh4r�Q��*�b��:�1<�T{f�p�7<�9��D����y�N�[f�lI��y�4�j��ڽ����j�
�����"�g��瘶�Dx�j�0d�����5A�V��nkVε����֌T��TsncMQTPU5U3QL���ܱ�5�����fbf&E��o4@��gw�"�;�ۧц5L�#j�s���nA���UN��jf��/][���7f����Syy�އ�3��Ofк���x�]I%T�:�֗�/]� ��Yu�:�&�v.�t��At��ZM wJJ�r�M����w�i.��%�=�෉����dB=O�8�>Gr�	���7�>�tq������U�^��η���V�4���F�!l�FȭS>�[�Q��y���L�E�u�Sa�\��`:��~oC+vqkC:���w��g�?u�w/l�ܱ�oey��,�K�z�,�=j�'�Lg��8���܊�}jnl�&�`�M���}��8�{́�;�^���m�o���؍�nk�Z���x�& /sG"8�}*��[]�s����>�b%��nx��ӽ\4��mBIVklvY<���I-�:(���V��n��� '6�_�F�D~���ñ���E`�,�t[��迗9SU}T�L:�ބ��h��qe�W�n�M���NBs���N�fI���?l��%����'gl��;����iƷ�
pȜ*Q�� �Y�{�g	����}ޗ�j	�[Z�ݽ{Q�m-���f[v.�Pw��e�+�q2=��bC@��Nmdmlo��~����6�pMq~�ڿ1c��ߝ�3� ��y��+./�����ͷ�C�ŕO���g����W��kc�G� [��sPF���~Gb(��_nᙽ�+
'��,߽�h�QRk�i���A]�3���x�]����Y�'�=X�3�C";(��4|1��A�T@�������UϞP=��Й���Uۘ}�)�#��E�_i�(�la* ���5O������26S-�l�*����x|�[�������+�u�:ܑW��I��oO��j�mo^f�L}�[�+�9]"��2��ţ�,����<��gz`9�_C�筌T�o:�yt����y��7��L.�1����j연g��g��esw	��q.��>:_��7q�B9�[�>����naS��-O0�Oһ�^a��.���Z���*ww��K>[3}��	�xS�|*�4��<��ד�A*=���sY��	���	*4����'�ٟ����`EH+�te�(�>�1�,�9�Z,�6�׎�۽�g��B�M�{��������np7}��c2t�.��X{��6M�
1A�w�^�D�UG)���8�O߼|}��u�nq�ʼ��4X���`����l^��H�~rGsc��x;��X�����'aN
���]o�g=>A���d��\���;R<���E�;qf��-\�o`�]F�Vt�Ks���g
���h�
�V�-@�2	!�<���#c��wU�̙"�@�o���A}`<#�jV�l��2��}���P� ��Z޽,����H.+@h~�_3��IH���k�sD)���&&�v����sG����R��yz���%bl���O��9m�S��OWt��*x �]m"�ԋ�s��m4UL4�nb�S�\���AYLk�|��#ۜwo�K(ʡ�{�9���^�"'3B��w}�/+s�	#B�%|�
�nC�Y�ղH2<z���2'�}~ZC�:�]Gud��X��G$BP+���2�Β�Cu�&y&��7�HyҮs�H��xEcY��ާa犩$���9��$�ƪU�gs�y�UK�*�w�um2�(���$���Ռ�������vΔ�kA�B�v:�����:��d��*�6�5�|�7�{��cx�
f0����?��'A�����������ucY�ztV؞
+�����`B��4�w7����s|���r6
;{��l^� ���-��Bٚ����8O)�3��u����Α$.O���jT��q�sx|���J®�Q��s��w	�%�W�(����L^���G:���ʹ}��� ���,yx��!��7�!�p���ox�A���MF���ԣg|GBa�#>���<��|����\�d�ay6��Y�͡�N���]B9z���n������j��Q�+��� ���h�����^ǉ�����m&��"L�����{��K��w�r B��ώmQ��+ex�d��{��	O7X��/���i�A��к6)��N�������@ui<��p.��= �N��>>R��Nh�o!��Y�Q��]����̪S�j�P$-�����[M��~Թ�@��r���1�M��{�Þj+�l�=��ĸ��S�D$�S?L�?P	MI�T�:�k�[0�X�����(���B-��&�a2�{�R�[){;��`��o�;U�&��Q'�ϧ���C('�\�|�ݍ*��c=����Er��%^H�o�hϽ��=�ha41t@��v|�D+��Q�g�Y3Sp5��@���Fd�ikѷ]��ӛ�^���u�j|΂�����,@S��'�U3D���O���Y�-Y��^�tc��SL��sN�����m��1�����a�4/wY�1�i�Q)z�$���Ht�t�vSS}\&9`^ �M!�C���]6��.%�L�˨�[1���\�kk�fnU�=�[E������c³Ц�4m�����>�1�.��ĝbzL��:�m�ݫ��`s����C�����tkzkUO��Ď�����ՑX���\v��˙Úv�k�3|z�q�Db��\��)7�˪��!�i�m�}��x{�6�g���q���۔.��q|���|.S1zH�����]��gn ��f�<	���O�fg8�\g�M�n�B���`����9?di'�a[�t�vn�h>��#����D��^9�$Ndo��p��p��A!D劆�c��9/h��=B���x��u���:v�7�؍y>��R=�f\v��������g!s�k��MEZ���]˪Ѐ�K��]���T�;$��=A����
aÜBY��$��f`�DB������
��B��w�r;/���w���tQMM�t;]O/3k7'�������9
#ۣ��M�àf_Ex�"|Q�Hw;O}�d�v2���z��b���1o:('�(�{�\	��
˴O2a9��̩
ͣ}��0��Z7��E���@��<z�oXJ����,��"�Ѹ6{g��Z5�8����VE�4T�H�I�*%��iL=X����5(�����E�k��g۞Y+���S�A�I������4�*�:����S5�s3����i�H�b�ޣ�6��7ͧI�0�$T�$��[�[9����Ww��v{*�}hYm汘�!@�"l��v
6�qW��$��F���N��#L�]6����i�47Z��ㆇ�k��Q���C{+~��H�yt���۫���I�G��D_s0���{+����&*�N>~4�ه�G��'�wdݡ�]�#�o��)�iɜ���h�&�$�V�A�V��湳,��B)u��D`����^����_i�X����>��,��C�h��J�`���ƽl�tq��%�6,�KMw6�r*f�⩂t|(p�ӹ�æL//yuW�>�:H�1�甸<�/�z5��S���^������\���K�P����Zc�◓��ڲ����[n���)4�����q���[?��+[ܦ���6������a�_t:�'�hH�\*�aנ���E�:G���k}��mx�u+
�<V�V��g&;����tzo�ǂni���S}�Gk~��N>W��l�ô�� ���Ǧzw�n+;����0p������ %��Z$�0<3��w�Ә��W�����'oU���t�
��F��ڠ'�L��90�6՛��3���N�G���g�� �0��<����94�Y[����Y���qU�����<�`��8y�\�as Ŗ�ӅR�(L�=R�"��.~���܈�]bu[�k��H�{��=G49�x\���e����Ӕ�4c� ����sݗ4w������׼3!/g�yJ9�%�[��!4oS�no����H�+��
-M�&v�=�J������?N��������S��br�)m�(�@��/-M�9���P�y[�]��4V�v�~���I�LG�HYܒ��g���&E����^����43r���"4䭬��+"�n6�d�zLlj��"E�ƽ��l��]����D!/��8�D%\E��5�i)ef�blg9�ow�k��
A�;^���T(�g`�\߯Ϙ�¦:�%�#�1T�$k������Α�m&z@)ѤU��K;tw_K�4�R�=�U��x�ՙ��(�F|�-�(�=i�u�6'���H�r~F,v��M:�V�c����}����;�~�^=ڔ�+��&6A����N8�e���ޭ��R��L��gK���Α�c{ԩ���(�x$MN�R�}:3q\�Y��I}��;���`?�\Vu*�B�Z5�k�=�W\�=�R6�)M'<�[r��J����5�4�-��]�(�\:���g�'4�Atz�uэ���o��A�J��ye��\L�z!hՒ����di���c���z4�W���8�wJ�P)�j������+��È��w���o��:�����3�G1����Q==6-�uo?�{�~���k�g}_?L��vwm}�v���"�ׁ�2<�U�LH������V�OU�`�H�l��O(��Aoi��G_�"�����Eщ��co�9f@tWTUɫۺ籺Mse�
��ײ���*�i�\\�ְ��|+gk��r��].�����Y	���(G!�5}���\�񔲵&ۍ�<]S�5T�[˺+o��n���!�
�h�8�3%Y<M��ȭ����LNKꬋ}TN�`����{�P=�>��3A�
��u����Qӵ'a�C^�٨�8OVк�R�y#*�#3���W
�;@O��x57��|����òn�i�Z�M�WKKt�J�I.���"�.#�Z��9��.S˺��e��9qt�{��	-n\i�L�ˉ����� ��o���/z�ٍ�E�.���c�^�l�ח/0 ���\S.%uEК��We�39B�
�6j���n����*�W-�{���	�f�üj�t��yyi��8ǲý=ǇR2c�3lX���|�i�͹µ[�}����n��'h��^<�àv�07-��m�Vwp��yCwa�����<�5���u��k%O�kt�r7��ߣ�f�?��P�������{�f��ȉ�.�'�¢L�V4x�8�k�!��>�:����幸��$������{ž�a��HL��
������H�S!�"�MI�/tו.� �?8��R���Z->bR�|*
�e�P:��o/��gů@��z�F�]@�k
K��Ӈ��w1����z	r��g�36��t啑.	P��x���Br�W�TLB��1��C�rj�l\��Yk1T� kC��p\{�
�i�����r�sھ�V�{�:z�A��mw=:�#X8�a6�W3�� z���It�i�3�3jG�}�ķ��C�jL�נ���wx~~qw���������W�������(
*?����(����QO���8=�O��
�I���a�a�eXeXdBV@� !��!�a�eX`B@� !�a�@�P!�a�a�a�aV � eV �U�U�U�!�a�aU�!�a�eXeXd �!�``Xe@�U�P!�`VVVP!�a�a � !�eXd ��aXeX`@�!�a�a�eX �E�!�a�eXd@� !�V@�D!�a �T!�a ����|���BVV@�!�a�a�d ��a�a�a�`XeXeXaXd�+�C(�*�*�*� ʰʰ2�2,2 C*��*�(ʰ�00�C*�*� �0�2�2�2, C
�"� °ʰ�2�2�0
�*� ��Ȅ0,2�2,0,2���FFĩ�E���A�E���f dp��
 C  C( C M2 0�2 � �C s�C(�C �M0�*�L��4 ȨʈL���aP	�dD	��P!�&	�P&	�@&f @��@Bi�!�P9�be	��H`Fd�P�T!�	��	�!��L�M2!C*�*��2�4��"�9�8L�C �0� M�p,0����U�P!�a�eXd2�0�2�0!�[�?���������RdP&O���/�y�����H����G��O��'� ���u�?S������������UE�� �/�����*��ĕUQ_��?�� z�|��S�P����������������?��q%ߠ��D���������xP�+��"� � 
*�(�$B  L� L�B H�� � H?� r� )* @�!" JȀ��# B  @��,� B �� B , � �� @(J0�2,�!*�J�!*��@��B0�0
̫$ R�J��@�����X������O�PTi(
��q��?���g�����x@������*����������?�?�y�O��#�����������?eETW��P�bO����r��+�UE��!�����E���<�*�+�������|_�>���������^�������8�qQU���S����/|TUE�C���`>w��|������|��p�I������w�%ETW���b?�?�������ߠ����}&_?�?����������|��>|	>��������S3����2����8�~���rw�u@U��?g�T]����������O��(+$�k$M�e�{0
 ��d��H�ϛJ@�4-EZd�-4�$�Zm�M)
�BJ&�J�m�TS@�Z�D�T�
�6ѡ�� HER�(BU!dY�+T֖�-�m��KY�9���[m�[[EUU��ݺ�[mm��bʬͦ�����!6��ݕU��mKAh�E���ճAF٦�$��T֚Z�֟y����m��j���Ƴ6�mmV-mkkm4RJD�X��wwaJf��(@m��F�&&��m4M� ɐ�ږ͌�������3i��N쵙k[m-��   ���[}���Kt�SW��j�8�=���G��΅�m�i�/[�*��Jr����'�݀����/:��N�s֞��v�j�]���zk�=�׮�mO[�x�����M(�w��S��-� �J��-��O�  �q�T��	_l�����q�'�U
	}��ozB�ԡ*�H�y���E;�m����S�p�)ӱt�k:�4���:���a�N/{Tm�kmG�5m�=�ikޮ�xҝJ�;{�^�ݻZ�MT�j�Q���b��   s���W��J����{���N��ml�yc�X��:������ӫ�k[�u���w79�+o]mO;��`�u�����ݎ��+<���m5/m��{ܕҺw���
ٕU��6��E1�ag�  �}���j��W�緸]��X�p=��ީ��5�sS��PM��Q�6��tu�x�S�����ޫ{�=z�\����]z:���m��lͬ�mM�V��  3<PP�YZ�c��z^�Pyݞw�U;��ڳm`
;QmT���^�]�[��F3�(QC��Yj�ҵ�e�T@f�i�   Yx����͸P7XN�����Ꝭu��Ѷ�VQR�&��*�+���s�u���2�b���<�J����,M���[-��7�  ��k��}{N ��f �\���z+��里:P ����@wW��@h�pz 
zgZ  r��� r^�Xd�Z,�h`���Z�|   ����;�w@� \�:� w�7�C@{�p�;�6�UB�{��B�Pz�� �֗�^�{ i�k w��jdɔ�lض��X��  ��>� [�7� ��#�({�n  i�7�� (z�{����1�=��@(t�{��t kG���Dl�k6ڂ�mhU5K6=�  ��^�h�=ހ ��&@��ޕ�� {��� �{o� �� 
��8 �����+ǯw� _ E? 2��M4 2���%P��S�2��   �~�R�=M�4 �!0U)��  �J�ª�CA��O���~\��}���c�������_��Й�1k<���e���~v�+"�K�(Oљ�m�y������v�1���lm������1���6�1���m�cgm��������+�3�+3���p���Gn wir��Ի���A��[_iR50o�ks%+&���%f]J���4P��ɫ-Ve���3E-s36���i£����b���e�$4��ni�HP�k�ZΨ��zB&��.]��y�V={�(�Q)2:��:�d��v�-�)G9��j��"fޜû���
�6��H%�Y ��Qh{�i�d�(m �{�2�Y���Y W"I�7H4R�.91^�%A��t.��'6ũ�2�M��*��vi0q������D�0M;ķcövm5Z2�I6Z0�f��&ն)�O4A72��1BKY "�m�h*D�+,��@���ZLǚ�u���RG^J�pb�,��3�,��%0��C�6��50�וy�U��,kӴ�/�Xn��vN��@����d�3,nS
!-!`�fF�I����J��[xp�Q��::l#W��F��j[l٣pfI�(\����#�U,j�I:e�Xm�c��:�GF���%i�JJ�X��xa;DXk)���XƢeѱb���6�*X�-BhmGQ��YX�F6k��6��5m�-H�&�Z��u�ѦrYy��8X�Q�D����{A��!;qޝIY{�[�rT�^D27 pb/j���Ɗj����I����[I	r���x�(��y�rRK(c�$�cv����D/n����,����T��Ta[�L�̬ci����t��t,��j��؝q�1�]R#u/,u��A,�bR- �o$Yv�x]i���k�_OX<�枽�k9x���J��A �-Z(S�DYKYSsn�A�n�`äN�c{����u-&�36�YRPfY���7@�r�*7D�u��Vn�b��YG�;r��Cl�-��k������Z@RČ�]�ۆK���p)�@w���Zдe�m��ߚכ��"�Ȝ�{inm�³q	�U��75�X`�6Ѽ�(P����o,2Ċ����iQ�h�Ae�
7F��07NDe(�ѳ�f�NYn�nef1��N��� ��~Ma���"��wXZ*�V3M���A���1�je����댙H���Z��FK�i�LĄ)	�Z�.�!&u:������X znBu�,N��ڙ�n������'�#��o��L-	��6�0�NQ)	��5��.	v�m��I�KIw$�,���(��� �>��t��ѭ4�J��)�
,Q��N�Z�-�4n6��1�X�����C��0hUee�[V�n]��B��su0�ZE@U���^7��ٵz�ڱSL��ۍU��anȨ�niɻs$$�S��2HQ�V�T� �6M!b�[�	�GFT�Je��eN�<0^Xѫnܵ�* �؉UM/TJV��5��k'����Us���6T���/ ��
���I�h��	Ym`D˚j�[���6�V�[�Q�ǆ:{4i�1ɁQqIwn8e��B5J�=���ɇE�*VJ�YX�C� ,X�F=�F�JV�n��	�5�0���Vcg�ȪaЬ3-��Ռ�vd�YgFl��i���t����љXr|M�3��8�4ay���M�n^RLh5�6�dŐje��3oZ{�J�8љe��-$^M�(�n�]���nT!�5����Q\�oor��x��eV)�ʂ�:�I���.�6�f,M�wV'Xah��JQ^I�9����VXvr`d�ͨ�i��-c/u�-�.�6��+h
�^m'���n�r"�+yix�$�
�h�Q�����5{�+vZ�^��<"��4:��;��j�W#m>��,B���Ȫ�2�T�Xi���<��-�	m�ٻ����9�6����2H��6�-�b��X���[��Q�d��e�+9tr�j*���hzH�H�`^��m��ڽSy��f���R���ӝfR��� �:���f:׷q7�����t57mh��dD�F�{x�����8޵ЬIG�&�����n��kX�1*&�4%Lᖯ,C#6�Pq�r�V�ac�2�:b���%�7#�S(Lؼ.�M ib�;��� Uw[��g�.W7�P��kMC�d��JpY1غ)Yp�Il���2ex>.ܼɠ���UK�e�i�� T���2�@W�F����0�%��[FIB���4o�ٚ�V�=�ٔ�e��&��54�ͶMe;Umn���r��èm�%��y �z��-�īr6jXԲ�����C!�P�^_ڧ�)�F�A�r7��;S3a35�����EV�{K��i�pa���
��PA��� R^K��q9��l�lˊ��Gq�yu�:�k�M�;��f��3�\���� (��CR�yl}���wtv���)d��L��C##݅)��ܺX�3�E�PQ&��1�m)8¨�VF��{I�d*P��Ї7��ފ7>Gxa��.�;��v�j��SL�&��u�E�n��w��I*e��{�5 �I�z�-nk�P��{F�8��I�Qn�KJȭ��d��aM=EӖySDV��j4B��E�5ι�m���@�;'�u�#����/@՘�L��7��l�w��֚Ѹf[;D5�V����wB�!�6�dȐt��ףr�[�a
��8�Y��Y�oeÓb�E[�"���wtm��r��&�/Dg.ٚE�EQ�,���XB��6Z�J=P4�l�ˁ)��m�"��͸
��/��Z����ӱ�G���v[�U�u$�w���*�)��d���6n!jG��� 5)Y����r�[B�̔�Uq��t��-��ׅ���a��U���
w�n0�נ����Z��Ф���K`�ݚܕ�g�V�2���f<�[b)V(��W���+*�,�q�<CO�&!�L���N�F�%*�P����ŉe�\�:�xn��9��[*:j=�> ��m���yH>�g2C2�]漡���Ww�j�FH[X��;5��9��ڐ��Y��SaV[���{J�i�Qݻn;�z�H�`����]��q0m��KN��nlQ,ʃ5=R
³u㩙�V&h��bb�5��i�$Y�	a�x��&L�V`a&0�R[�0Dզ�toaY��+�U������nZ��s\���LD�̧5�1� )#8턎c��S)�pk�GQ�M�����Sl1p�I�[N��@@�h�z��C[�J3n$�.��M2���r����`�8��|�-,
�/������N%�"!ޣR��bD
��ur��U����!ۣ�w�Qj�j`^G/��k;j�h�̹x�`�PF��5U���z���SK@x�a�h���,�Jxv!i�[�QȞMf��c(�kѳP�[�%A�]�T�70+N�g咄���tJØ1Yxt1*��XȦ�V1���I'f��n�VX�2Q�V�2B$7tlx�o*�j�%��݋3[�'t
u*^\K�,cĢ�@��ʹ���lT�&Wb��8�Y�5 ���,ۡ��3n�^at��h=�b.�eB�aI(�i�k2�Ӻ�6�i_2�����il�5��S�v-ճ%�h\9������S�x�[��X^����n��90�$���4�6m�H� ��^�m��+��Y�wL��B��SX����b�]�ŒTZ�5�i���ym� �C�E f;��J�f���Zb�M��S-��1L�h�Ɇۍ�°k�>K�#nrӪ�P�o]�1�wږ�%;6ۦ^`�Jj���.���]k*a�
��C��ujQ���J�o�Q� �\� ����7�sp'g��kf¬�չ��,��*,�W�Ȣ��a5{�-փz��ĉ������1LQ0feɘ�G�Ҡ�CF�� �k*]l�ѪR��k*���G���Y%��_Z뗝DtJ��'c�4����Jۚ��mamm
�d�L&�-��������$,�Ӳ�m3OpQb�GXUƆ�V�_�Z��V44��5�[(;�m^��\�5��t�h��i�v-Eu,�!1V�ط������nkȥ
Z/S;X[�f[V��+-��P�H��2��4^� T��ml:Z	X�.�]Ǭ�$�T6ds#�b��{Uk%l�)�a�ܓb��w����ԼRd�豲��H,���+,�І�skr���R��� ��e
��e�AB��(�Z�:��31�,�wd-�ui��2�����OB�azkyq�y�J�e�In��� h���J��SR����j�O+`��h\;�36�(�Æ=E������B��N�k+�헨n�oa�2,˭��溗uRj4��%��yLů\���u4u˃r��.J�I��#L�IS����BFm�ϭ7X�4g�p�I��j��al���ACbM����G"��~ � :Z�C7��xX$\�0DtXak�޽��V�Y��Z�i���^���ΐ����A���Q��� ���5(�[jՒjm^;��f4�0h'R�f�fc_�#z��ƝjҜ1P�����s>
�AfT$ix�7y1i6�)��h��������l��P&��Fw1L�q�^�[t�Ua�M6�oVI��X�j�Plj��&d��/YN�N�PI��ڰ����@����&ѡZ�+��76��t�����A�Ӣ=Z�r6k!u����������۽�P�����p+TX%6�������{g&�'Y�#���ܫ����=8Q9X޳�+IJ����us.�Ci�ڻ���̊�k#{e#��֏7ON�[��ʭ��H
�T�m���)i�E�j�2�V����ֽx�k�Jn'
�-k�)�fH����yy��T���ҭ�xP7m5�������`o-��J��T�Tԍ�t�,M��i�C�V�ǶH�>:��]��.���S"�N)��ݫ�cg'ҷ#���g,j�q	1�-=�B�I��`��i�+�a`�
"M���!y�s �;�vZx�E��2,�3>�e��6�e�:AJu1�%���2�Y��D�ݬ4p�x��7Y˿��6�*��Yݓ�-I���u+^(�̀���<BL/q�VZxk18;���4T�΅�����ɺ�Ud�,Ӗ�^��oE<+nHC9���ڈ�9)3fl�� �����̩��n�j�a`�b
�Z�;�E�Lf9y4Y��J�d�fe-$cc^�ۻ�O
hH~:ܥ7�� �4�m���vc:�+��4� �b��HK&�wR�� ��JÆ��V�,6	��B��X���7�]���xa�Sif�Ĭ�D�dE�C�1e5S�B�5��w!y�n'���h{bPY/+iMt����ڏm%;�����R��Qb{��r�sT߱�v ��y@],�BhV͵��aT�,P�U)��l�Z�T��$�čM��n�-q��k�xӔ!�ָ��w�����8.P[x37I�C^�QԖ+*���J��~T��>Y��@�N�	7��$i��R����\�+dW��������ˢ�T��=Kc���@ٳ���ɓ	���j��7��e�Qݫ%!�*�E��K��8�"WB��Q��*,�d�v��9Z^|��z$���#Srj�WVU�n3��ⴊ�[[s6]l�� #EM��H��ǳY5��/�Sմ+A�EbX�CF�%�s�w[YQd���y�NȰ���*y*��K*:[X��tp^n�nK�!C�fj�p�yG�"��`�oZ'd�R(�ȳ���=��bh���o��&M̄W�f���We�{�9[ۻF�0��ySn�x�ު�̤u��Ńr����U�֚;��B�� c$%�/��̍��]1M[ӵ5Yyc������KR
�5ԚVW+l< m�tEk�(b����[����M;w��ծ���-,�w��;e�v���Q�B�#�(\`��	����fY�w#	�PӼVn��6�kBSŮ��O�
�3vIc���L��K+( �Z�sh��St�Pdl ����Ų���T�	-�uŶ˫7j��u�G�@oA�c�����ð���d���J�n��'R�q�)�X��0˓u������E���+��BI]�܏"��V�衷�KsL�#M�۫�xa�GtS�岰̺֦<T���e�*��jKI�3%F6�`�Y,[ۺ�@gɺR��U�n��q�i�P�&�r����Ay
ջ�B�hSS^kwN
n��y3-�����Ij	��2U]�l�Ú�2滫��61+iݸ>Z��z F�4;� ��&��d�������2<@��!yv �C���f��WF�wo27A��72�1��,;�%��D`3#�F�6�R���!8o8%]J루����dp���oQpU�V�ͷ���Y��Xz�H��M��t�����(�R�����Tӭቍ.l�Y��nY�j�U��@��+�$]:z���%yXX6-�m�c/Sb��d�f�Hԕ�܆����K�\E�p���� �����sIF��Н���Nff��~����$K�ۦ��n��2y�e�:y�L���<沉ӑn���B��v�B����y��K6��;$�VP��dA�keK��-dV�l*��`Y!�,P�.Z��cq�O+*?�jc�{�+���.�!g��C�L���������5P4�ƞ��WV�h�d�ǰ �8��l"Ϊז���o
�����6�3���)eХ�������B�V��L u1��n�9���VFi&�SQ�;��S�%�O��	eibe5��[�5*��l�D�Վ��p��j��l��L�Gc���@>W|��]a$�I����$N-��Ni	���S"ӭ�녲s6ɸ�b�������mli,�\w��-��"�X;rV�N��{�n�G���2|h5.�e4�66�e:i�9�1�`^�E2���_w!���)fV�x��l��l�3*�^hG^0��<�|�ouk��陸��T�t'AQ�5K�ٷwFqͧ(��e`�V,�j�]*PW.=�e�����7��:��c9�"�))����֓���ˠV�F`�q�1<:^��5,�������1����޵~Ƴ�f��m�핹&�o�4�si��4���s�Xv�e��(djY��]��t�����C���^=����f��!�|�^�ԎG|��
K�G�-�v3�Z�	��ZL*l�j�Y3k�<�-��o��+���v��3�yzfŧ#��(溾�n��QB)]6<E*����4_ml$B�ʸ;�Z����p)b����-$$�%;�,�؃�ή���x���D��,91(���G�SStV�4y��mL9�����h�cK�tɆ�O;NL�TyI�j��tG �/c��2��B��nKꈍ�R�:M�d���es��� ��wS��B�{���U��z$��ز���&PP��7�L]u�)��� �r7H����e� ��y��Nm�M�Q́�۠���7lӨ�������Dq�sJ{�J<��2ct�m���[v[�{��T�+F�W���CΝ�z:��Mw�^H�w���~ܖ�����f�	�T���Ť�CdT��Cq�bf����e��c��a9�ѮZ[�TO�Qe�5{��PNlʷ����;�t��#�����l
�NO��z�Sҥ�M'��J2�/3��9�ę�=P:5d��o7-	��:��ѓ��8sd�{��&��3 ���5���C'GV��Ըi�o:��8nZJ-�
�t�[��(�>:p�.�f�[X�oM}�a��Sh�G;{�\D�H�{�wZ�^.��b|���m9L����k[����na!����+wZ�br��柑U���*ی�Y�S�$Ĭe�g�R�m[�yK[����Eٺy�R����7H�5��,�Ge��Ɂa�j��˩��t=����M�,���v���N�f���r���s.ئ�K���	��JX&正nh�Y�3�цb�Nc8w�T�JL��t�*v�� x�pv]�]�-������\�۳����W��S�{��u�܀( ���XmG�Z9t�c�`5�5��4C��ۉq�v�I��H
��|w*muu'x�M�\�>M�D��ui^�tx)�n7;*.+!�n�Ѹ�~����ޝ���ՀuN7B��@\�ŷ�t���(9��'��uY� ��6�� ��33p��q�)��?���>�S�U����Q�}���X�:��]s5�������z�Ԭ�.S�4E��ڔ��oI�Z4�Ƨ<�]�tfG�kqG��΅WR��*��ާN�`��R����zr,�l7�:�����V�����)AV��"!X�S�盫�Ac�	鼞_#�ம.im�Oe��[[9�����v�a&��}�AZ��s�h�$�����^` ���R�Us�zx�)v��:���N�h,8�q�ޡhUJx�.�2Jz�7�[Uk�3)�Pځ� ���)C�Z=���������R'L[�f�s��Ћ�[|��$lC}�#��hL��	�I2��/wu�jaϤN�7ˡ8Y���e"�����ţn��^����CnTɒ�H�
��Nt��h.������ܶ-gJ�/�����6���4�k䛖n�FR���a��6�ݑ�:�f�*�v�f�mf�-멏m[�
W�v�Ęw9����t���B������ ӡv1�fԾ���$�-�:�^.Ù�w,w芶�XFL·,�f�r���;[x�[p"XS��an�<��eS3KPq��]��L�y3\�f,M�ޢV�C��Q��@W�!x�a���3w{4	���ޞ�H�\�/�¸�(8S�5�6�2�B�b�p�DԻ��_Dm̫��Yo;k,G��Y�Ʌ|��f��Gc����q��H�#x�]wj����S� �ɺ:^�o'cFuc����ɮ/芩+u+�A�&q��L�ΧP��.��QX올*MδDE��V�M35ZEn�C�F�튙���g_T�ym�b���"�;��3��,bZQ��@����w>���oJ�zN��<� �v�'��^��Ws^�\� ����Y�]�kkY�F股�7��þk���n�A��S�YtK���C�Zb�Qa��+j���Ӿ�f�!a䯎ecZ� � (ENK�;A���	���t[%�·c��3�9"lO���J��	ս]���^��/6���bU*������r�ȸ���&9�I�&M�oij*1����r�8��(�ej뫤9��3���3#NfFV�G����KQ#Պt�u�c8��W,��� �b����)���-��GW\��,n=XwP�����|2�@�aT�va�\O��o#b�g�Q��(�K����Z�$.�Ĵ�������������E�ء�+��-��j�3�FE=�ϊO��Ò�������:[C3a�A}�h�A�.\A�Zܔ���]' Q�UŠ1�!�΃Ek�g�G (��ռ�G巯y�T�����d��{��*���v��ʑWejի����g5�[����	�E���}��n�x�R�H31}���	�7�(v�Z�+�������:�
[\:Ƽc��5��7{d�C.̫"�7rs[���_ȣ�L����%��_�OV}�-Vq��ty��~s;��(��}��L�q��p��ŷ��6_@�|��	��ң#��Cڪ0p��S4<Τ�S��R����+its�w:4���!���#�!��7o'S�.U�AKW��Ѣ�'%�w,ޡC$dvT3@س��6�z_ʋ���|#ط~���rV�R�%`][+ԙ*kN��YK{�0cV�ۡF���r(WVE�"h*bڻ���>9�b�;V�Mxj�ݕ��#2�b�
0�*��FՉM�]���}�$)X�v�`�}\]��;R�q��������қUnj�r�>v{�m�֘��wp�Y�s+���ҧ*k��kB{��4���$3���ectI�7kBȺ��ؖ�z�K�4,������&�����Ǔ����q�� {�y<�iL�t)�c�a�m�8�B��.���b��V"�K[A����x���X���~ʁ3nEb��rATc���k�'��y�Ƭe?����r�eǝ<��c풲��f	.��)�����a��C��As�W5}��cM&���SL�S���͝����ۙ]�).~ʹ����~�sD�^�\���x��E'KO*"i�g����R��IG�7v�Y|&㾤s&9Fa!<�au��n�ڬp'��B�5���;U��:��� ��uyq�8>�R�t.A�^N�縦3J�w9vt/zR/8���j�����n���*�s3w� pP���x��̻��eM�.sqVǁ��V���0����VȶÕjŻ�)�0:˸d��e�O����wc�En���V�6�,�;���y ފv��*�	�a�����1�"L��vQ���Ѧ6VI��Xz�o5o1�g�!-Y]6] �f���9�����-WJ|Ʃn����s���® ��l%贚"16��ڑ8�ƃ�ץv�j��N��z��H;��-,������pާ38�ޭRhS�I]�L��nR**�BWf'���L�*@>g5�5$^EYS;�Y���x����B�+�m�shJ���y��Ì��ͻ���Ϸ�
0{�j'qT�n��7� ��j8�)V�����v�cb�p��h:z�D���e*�l gX����$Ry�z���z�
����^��)���'csQ�٧��n�V�Ш�ʱb�&��79�n��vC������0*V4Sܱj��u� �a��FR܄d�5Mv�0��4��9�I^+��Xٽ�Rҙ>U�8��u�4GN�.����w���]��w!z
�Kq,��+y��`�0�ܡHf��s:ai^ĻP�O��"��z"�]<:ó���eϹ�ȭ�8$#���<��E@�����ca|�l-R�Pȑ���.mg��X3��v��8S�E�w)�<t�^�
�r�o6ؓ=QL�WI��U73dR���M2� Lq�;?A��\m	�&ts�t�1XuD�N�:�5\��}��,cf�Z�C���I��3)�[q������hc͠o�����朒�vD�����s�^��r4�ޑK9$��k���p�K�Z���C�:��/��+��ʼCI��F�v	{:�S� כ�o��X�JF9z�96��m�����I,�ȋٵ���M�z�Cv�㶻��+�sWt��Y�ߵZpS�}��h��Et�V�I������91-L5���Mah���괓f�C� ʂ�g�`�8���r��QP�T����Y�#ۛ�A�U��=w��\�A�ؤ��B7b�R4��!G ��ʛȉ,N����w�+�q==���H�u� Фȫ�WJ��ju1vy�+�4h+'9�:���gv��WwF®Z7����Rޙ��k�qU���Z���)HoT:/0-S;�n����Z�ũ�Iugb�g>�LL;�����V�r
�6�3����n�CNU!(�[�R�*�y�E`Ű<��N��G�O�r�Ż$�Ttv��]<�%��	���L����;����-��&���e19(����x��ZV���`'�����w����������QP� �HjX�3r�yvq���Hlɑ�W)��+A��[cO��X\�aN2[�jL6�L��Ew 圅��u`�T�.�hF�I�+K�o8Q���-����ՙ�r�_eM΢�al�M�SIG�����R��WP7�0�gT��-�t37%r��v�XY�^��m=V�*x{�;��kƹ�pF�:(�P	���Q^��t8�N��u��76[����e5Md`���o�+yG2V)�Hr�Oj�gG)�|>�'x*���+Q��dq���_E[��9.KM�'\#;m���(��b�:n��/AJ�H*�3-5�e�Y�o�uf�.����J�L֛��>Δ�8.�+�Ɍf�޼z��]�s�ou�s36^LoT�{Ee@��eh����rv2�i}-Sr��z��Sۗ�۾v�k��t���۵����[ڬ	����^a��X7b��筲�o>r�.l��Zs�=�N
����J��:�S�I�p��MA�S���-�+�ppP"��t�R��r^�ú7NZi<�Bs����n�.�I�mXֳ:�N��:ڧ&��b|�Je�724�����p�@�d8)��x5�mj�r�Bw������cN4�-Lb��n2�]��J��k;��A�w��l��u�Ï��L�l����a�GW�gRYs���JR-�8	5օ��g�W����t�z�9�ҽ�c���e�e!��H���/]��F��TFJ�w��|�fs@[�vA�ϟX7	�'cm�㥲���O�mfgp2@��e���2�s�
�ifi9��K*�Uc�K�wTb�Nһ F关��)��7y,�1�Gl���xGM\I��p�a�.��NS�q_0jEySW]�٩�1e�F��qKc�N��N�pڽU����"�QnO(�}S���+97�|��I���Iu�����e`�`�����{GMa�W�XYf�#Em�|��[wi)�q�cI�]��Ak�K��Wt�u�垦r�dҦ˅ؙ}�j����;�t5cbɴ	�2�����UЇ ʓ���^kg[�J�,N�4��"d,�%�q�B�Nuk����>c7;l��U �e��V$r��+Թ�{Z�y��o2i��\�Aѝ�$�=ҹ�l7;y9���rU�lZ/-f}��E8��3��lJ�C6��u�|a��]�[�tJ!�b�L��ŷ��$[��ݓ�*`���f.i��9bT:�ܾgT�A��fM��6�;�[]�\�V��	�3�)��A�-�#��W:�u�iB9_sd�J�s�Z�BN�a6���h�ԩc"ZD��\je��x�kZ8	̲��hغ�m��N	Vp�j�x���ᕚ����0o���]�
>0�i&�tf��"E���u����wC��h�tfD[��s�Qf3eX��Y�`O���K�>�nj Z�vl��Vɼ�U��e�����*��/	Q;A�����f�*�)�B+4��mk�p-�F<{�ҹ"�Sk�>�®b'k�
��:�t�쀶�|���g7;1�R��O���+���콓9Ŭ���8w�+�}�;O\Joo�[Gdyм=er�I��2�[�wj	�R�GX�lxwhkS����W�C(�@�U]�0�mg*J��$�͎*�Ĭ���S�d�eKr:&��^b�sr��g_X[.wG��)j��`O�e�*M}W66��d�%r"sd��{y��^(�] \�:˒\�Zn,h9S~�2��s%�x�E���i�Ú8��/�y��Q1���sa짽Z��qv�e��iV�#}��ӽ3�j-u�sZ9V28��y+u�':���v�����7�:�{t�D��w�ú�n$�(�7j6��5�+��h�ouJ9V�oY�L1/���"-\\b��F��w\�Z]�[�\Nc�L�*yk�׀&��av{���'r�Y���(p���$+!2X-+uڧ�M,YQ�re���+x���D�&�+��N����lU�C��,{���P���V:�b��:���7��u��eK#29|�һW�2��7�\��.�iwK+��G��=��Kt��J��F��qI�Tec��s��vF�vR[��ǻӪ�oV�R�Py��҅l��˂�{G���V�^*v�"�v����)��d�on�B�u&��A�I�e�w�D�əz�H�����1@S�ؼ�5������0�f�f�"��~�Ya���~�"$�T��1���v��-�0�j�� 4�7���w'2jXZ��@J7�l�ݧԒ��ED���)���wݪi�U�N�q.�ռR��h���Y��b�TЦ5(��}1KM����R���6�ė*���O�u{}lg>�/�Uս5Ƈt�MR�S�AGd�t"qčn���PXֲ���%y��d�w�:�gk+���o/n��XS]Ud���{n����g푵��Q��Vu�g)�{%��lھk����ޚ�))��k+tme�CqC�M��3X;z���/�8�6v���1'� �<��u]ؔ�#��.���mb#�6+��!��U��d�TX�� ڝ�K��m��3��.��[��Doɻǹ���g]:/>��rnlw�����״%�P��p^|3^*��fѥˀ&r�� }�w%sn��S�w�
�Ct���Ee���#�H���
�����0I��K�U��w]�s�T�eU�hWX�}�jP<<8O��VƄ6�N����R�a�v�H�zݡ8Xu��lM�������(�S(uCx���\�Y�m�yCE���!̺�Q�Rʔ�h_H	A��Gn�A#,Ǚ*Zrg,�v0/2f��Mes��,]A��2�`�ڇqQ�;�'�[G5\�Bݕ��&�ڙ��Xu��>��hg!���蠡�}X��}9�8�n����9շϴ�ʓ.�E�0��HՌ�z���q�*L�8�:���XdWB��R��z�k	Ę�;*����Ǡd�5��$q�����2�\`3R���6�iުq�͗�$eqۑ�*�Mj��VB5�:�ڕ"ܖ�WL�&n.����G���б�Q}���[��Ҋ��f|"�66�2Wf�ܤE�.�D��YS�N�Ȁ�	�yJSW�s9D!Y/�5'�}|����i�	�vql�]��Ү� \� ����݉e�Y �X�2���yuHY�5*�uK�s#ߗ)Q`�,���������غh�Q58������ñC�tQ�մ�p�!���}�e5��!-�Jj��)�]��vR�A�Ƀz�-��r�l�;R3��KcXz*ʘ�GENכh6��h�n�ؐfevl�&���F�Gl��wN�f�e��1.�jP�����V�f��.�S�P�dц\)|��_9���
[��)��2����:�ݱ��+o���[6�䤔�.�a.Y�"�X���;_w=�^iȬ������7)Z�a�#C�0&�AC6��x5_e��=�41�ѭ�;���J��	2��t��е;���%������qu�BY�T��.�ҙd�wPV��-cX�:��}�扷d���4�c!�3J��<��������_'�P�S���*�JUo�=W�hHC;1�i�1!�mg+xֳa.�$��Zu���%+�WQ%Y6Ԃ��h�x�S�R�2�yv(H�ev�nV�;�Y�RtJb�����ѝ���Z�olL$;���\�D��k�V��#*G��!���]tub::��'��7j���!�g5r�Qćf�0��hl*w�A�ӳz�MrS����㦮�<yղ��L40^���+��
�a���Jq��/�����#;.��no&+Lk\�3��2��c©;�\]`+�6����ZL�_j���R�M��X}ZY���bH���7�8FA|�@(�ώʍ�|,��d�itߢ�{�<6����yp'��5�Z�԰�\3kGkm�Un���Xz�K�S7$��qU,�=�֣Y.EVsr-\�4��{��9�Ik�ƺ����|��z�����(똷�<������F&�g+�i�s�]8�#��Z$�3��}�0��B����+�Mfo�}|�=ܚ�e:1�1�V&�%q�|(L���m��ßme�N�ƴ4Xtחfa�[Y�M��!��,s�M�9V!.����70h}I΄c���q��V��f�U�ԫ��=.}Gt��HƷ��Y�eij�X;�N̵���儍:M���m��z]��r�v�2dBL�G;Z\7{Y�"��ࡋVR��]���-�J�I�vK:�'b֊�w�����'��t�[��z">�:AG*f�J���T�"�� �2�$��S�`�r.��N�x#���՞<�� �ɻ�ۻ��O+�yQ����p�I�ܲZ+hH%�V�on��z.��x�SNw]�I�)DB�����8"�ϰ����q�Z]�K'�EK,C�-7�c����5���W6L8B�k��/����G�%6�S���xMv^rX��K}���ն�TvG�	[�u��f����S6�u;s���Vd�0�Q��kU7�풵is�� ޜ��M�`�h\�6��;��7�7�"a��_uu2��+�{5uh���d>ך�R�=;���Y-�	I���5�<2EJX�j���6l�G8)T�ʨ�؅oZ'n��ۆ����%v�X���g�YY��������)�Ά+Q�Y��a������B��Q����]�w�^������9j�[�P�-AP���,�9O�����ʼJ����cD����cʉ�� �31�c^G��v{X�]}{wÒ�Je�hY,�P*����n�6�}�Q>BN�(s߭>!)y�i�;��3s!3hN��kV�M�e�0pȠC���a���$\\�}6l�.$�͗V4�z	����@�yr�7�{�i���3/b�j��9��a!�7=�-���x���4)m��9�]����9��Mfhʸ��yyY::����P�6���ݞ�n�d;0�='�ނ�tq�|�`��J�A��N2-�Wg*^ę40��H&"�MANA�p�e�f�띣Ë�k��J�p�e3�u��z\f�ol��
7�"��&�5Z�/���勋	��D;{�6Q�\Mh���XBh��.�VhлK��e3;&Tzw��eJڳs)«�BU����A�Bm��z3����<)rAX���q��fh����{�ނd�ilV�wE�������Ӻt�Z9�ɋn���֡U8���Q=5�"��D�eC����[�3��]�č�9����a�[._l��6���ہB��հ
̽�P�,C�e`g᪬�i��Ku-����Flyn�투U	����9�R*u�5�</�U̞�<�QA����K��i"]����N���Κ�����'��Ź(���m^Gi�zLE+�ٙ43��%Hql�ܭ�B:T�Q�;�t[��͙9�r�DW��Om����fX�ά��T�����Κ�^��6���WLih��V��i���3�M'�:��h<G��>�m�\��t�#8`rh}����D�a�5zV��|�kqR�N֨:��]d��)esy�iP��3��X������`��i┨���&��q�ݩIS%q�=z�nj:�4o�P��h�$�e44j�e���b}s*�������G}5n�e�:�l�1���k#�/0����ĕt�횅��;n8�5��ý|��[;�^��]>Z���Ԣ�V����*#-t	�d�lQ2q�ȝ/�>�y��}a��vD�{�:��N[%���ݬަ5n�GF��wwk�q"�Z۱��G��F��X�a`�0JȂ��1�''e�W�ŻQ�1�y/�tt�Vl�����x��Nt�!�k����N����{�O�m�Ӎpz����%Hn�J����]�'���r����jNc�4�]�׉엂�VP?dfvj�'b�ϔ��Ɩս!�c��Z�x�2�_LR �h��Ek��n���Tu�kv�@��,SsZGC-�;�����6��X�v'0��ҶWLO�M6�Vu��*��t����HhR]��dw����ʔ��O�^-]�=3K�j�<���ڴ��ؗ�U8��S���͛�.�
�vH���͈6���Z]���q�^��r`Ͳ����3�w�*싲��5Ykv+�V��Ni<r�����̮4+hԾ4��o%��g%1�Z��q��<V{;�T�CJ��X�
VVS�T��ڧ-Lyci��7ي�{r�=e�S%G*Zv2�(��Ԑ����w.m`�����*�;��T�:�t�_<��1�I�i�q��Z4C�N�Pc�y�Z��,$]K�4����o9jX+�va�Uu��EY�7�.s2Y߃��[��v�5�b�[D�i�{�1�5�Eշm���lr��e�q�]�u�Q���LU�9bz@����汱6MKVl�N���i��JF�L�.���6��|F��i��C#�*�T�ѭ؛��\����o.ח�ѥ���7gnX -Bv���i)����nR�/,'�	��v�YkEm�Io!ѠV�G����/�O%�d����Q�o3of"�H�s�c:VsyE}�+6\tv]w�C܍���K�T�kO]0�{�ڝp-�5c�0�#;��O�_I�z���Wv��uJ�yy�]W��F�Kq�Z���z��WE���4*��pdn�����Gf�)]��q\k�ڬ|���IP�J�6·P�N��K�N��M�5��Jk[�W�B�Jx	߳.�
w���F=�9��.�,[6��vy�;����<(����^���ܐ��N��on�6�&�Uzh���, �%݇��os~�=�2R�@z�VtgF�eŷ�x���09<��hT;��z� �l��쮔�'�j^���d	l�L$C��G�kʷn�r:	ǌ��d�w�M�W��%Q]��P��z&l$V��I`�o2�ݤk�=�6��@řh��Z�*��kp�m���ι���Y�xs��
��{6c1�L�ڔcٖ��JiM�&m��;�M(�ʥcB���:z���ZF��b���m^�7e-&�7X�6\ �,������k30��su���$Ԭ�k�N\��4�g �k��+V�d��������4��o�lN�q	9A}���I�,�盖�T��v��;Fգqg'"l��1RXF��WZ���,��4�7&��Wfm�7AQ�ī3T|��K���M�1Orŋ<�����Pt�i�@]@�䋧�%F^Whq���t�a�j�\�����^�� 6�NMX���c1�'�խ؆K���=*�܏ ��V33L�b��`��+gVApް��P�W|9X�a��8�o��Ь�W\��te����
�¥�9SI��`p_٢�%h<�No-�{yԔu�o��I��v���@�h��;m��������3ف��/.�ܙ:�Uǭ4u���'�1�n��
��aȬ�%8�����R��:���Va�G-L|���{/���T���ʰ�ڇ��	M�}���K���!��L�ݦ�̲��E�ᙘ��e��в����.}�@��ZK�������"B�PÕ�5x��#6YG�qf��Y"����1㥽�����M��}:�v%��t�����I��|i�y;f�Nٷj��'ob,42��y�`E9�T�w�-i#o��7�ohV#�w�Ǵ�
��/U��N��[��	�`]��[��Z�� ��<H�	eLTy�Գ�($u�Ҋ#rg�_{�)�Z��tgrkp�A{��ێ��P^_P�p$s�L�퇋���5�+�u2�#;N�/7�&�w-���{��IO	mn��:�D�CS@�v#)�]�o_R��m\t~R|m᧖�ʬ��d�$ԻhTa�35�Zw&��s(Y������(��MIȋZ�Ʈ�RW٠إ�zv��
��#V8
�Qe�]1����Xr��gJ�]on,�ie��0��N{r�Q�R�֎wlH,���T�%���f'WZ��@�]��HبA�e�ܑ�H���mf�n��e���i�)*w��<Πӓ�"��R�9opԉ�cM.����n�>�j�ZBО���/ &�6,�B_�+e�>l�5��f̼4n��@��$n�X�+��bc���������o����\�
N�
6��P��
Ƀ s�S����H�)Wv�9^f�j�Ӷ�_­[N��?�^��=�I���E�:V(�[�Ɗa4;�u�+�w��N��f��ꫦ�t��B'�:��ڝ�K���q"ť�e]'�LXf�
C��n^*lpz�vP@;6�f�S��Ӳty��<�Tb��J���9��9�� I�C���ʹ��is�Q����47u*=V�f�
�:��F5G"�T�X�x��r�
]=H������x��Sbs�5ҭ*�\���)���l�+�X=�Sd��o�����ʕ�؃qp�zڽ���SX+�GV�y�7�^e �Z���6Z�>= �Q=���n�L�L��6Ҙ�A�3����`���8�f��e��ik&#�A�Q�A."���|��̽�+f��,}u+;+�r�w���RvH^=����3��.���pټ�*^�[iX*�Q��Cuc�ws��Oh��/�)o�Q���:����-[��|k�n��-.� Inլ�M��-�Ҁ��ف��K��,�IJʶ�3G&��l�:�@u�̵Ϟ]�u5�Q\ַ�ķA��,�0�L���>�ɽͷ7eP{���s�7+��$ �z��e"��2���ح�,0�o.��;K�����ff�|[y*��JT�}�&۶�B��F�[څ�;V�`|�+����U�:Rp����ͫ�����R�ƺ��f�6�P��Ȇ���4��\xt[�������M��h�]j�f�^��6�gTq��4VW	�S��˜V��cX�VQŊZ�՚�3�Y��f��j��pe�)L�7���
�y���^hsm���Ş�U�t�F�l<0^���7��0o6/l5}�.�辋�=qCj��BvX�e��Elu��ЎY �Ѵ��Z��f��¼�˅��3 ��3c5V��t��Z'�����qr�Դ���y�{�޾�o��L)Q�����
nT/�[d�D���Ψ���p=���ws��a-��b��Sw�u���enI�[��Ú�\�)�r�I���-��v�ی�}iJ-t�xw�nl�̸y6RZe�ŗ;A��Lp�\�^���p*W��a�<KR��k���G�/cܤW���W@����U1�9�xe`�£v!�o�Xޛ��fr;̢�f�
��}u��r0)�;e �"w*D���'�i�NZ��-X�{�I��A�;7b�L���}Dq�-�ϱ�Ş+SS��'o����Ӛ�6����u!.� �c�WY�v,���:f�nVr�l�D�r��!���3:�dբ�++�k_#�K�[��#��-�U��<�P��t3�pmX�N�u��
���`$��)
̒n�>�̨��tʭGV�૔g8�W]�;�G�v,h�u̞]�lYp$e%C2��ﴊ+U�K�P�
hF�a�X��4gQ�p��x�WT7��P��t���E�]4��d!ٗTK��t6]G����]�4	rlqMrVjp!2a�G;Q�j+�{ڧ&��f�O)�z.�Fd���z�)�TԤq��������L��c��v���NsFD�Tʒ�:T�Ր$�7W��݋����ʯ�d;��<�]u%cV��آ�a.�D�¥ �eٜ |J�ʐ(�h�
�RJ!EӪ��RWB6�$�*�!��i���Y��Y!�A��G4̴D�4̪�D��*�5�����I#J�6Z&jj`���`\����Mf��h�"i�aT��B��������ÕU)\�J%��T����Z(��jE�M��TTe��J�Ȱĳ.�Z�IUe�iY�ff�DY��ILCi��	DtYB����.��PP��X��-��r�Th��a�M%0�,��
�PP]."RW
��sL.E&h�C$�H��RJФ­I"�C�f$%������ib$��8Vm-,�i���"�9�I)��:	s�<m��_<���:łdusut/^����B� ��]�G��^�����rK�ʤ�|���r���*����&w��%�z�3��S��^]ߜ�����@���+p�,����p��q֊�ގ�om�l���F��]�w�w��z@!~�o��:���C��k=��12�hYע��ﶭL�U���N�1��2���;\pxV:�z�^��3^��5�"��;���O�l��h�V�O��~�ǧ�l�����	�"��fƗ�T
��q��S��PW�τPtڷ�:AJ~?q��o�`K�i�Ĺ�q�;�Բ�t� ';⟽��Hf�E}��o�a��D׼��t���`�Y��v��
د��w�R�2��}�m��)�J��1����S���%�4��\��}a��ς��@t��𫡜@U2u�{��b�t=�ܱ)�9��w���$�нUio���Xx��U�2�"��(1>��}����x�N%9o��]V"�fmGq���Lv-�
��iW�ip
��������N%	�Y���Y�v=�+!.7]���������:�.q���(҂	%4"����%��kL=}I�OR#O�q&��[&�)eLT���C�����=&u��BmX���J*��G�G?�X.���t�9M�r�Z��J*:gs��%�2��	)��2�c��D�����);�5���`ed9'L�ӆ�j��L��SbRwbο�uZ�Su�r��Z�#�IҬ�?f}�ʂ��6�9N�	�	6���m�[�Og��-�$�9\�]p᎚������u�K�Q:xU9�t���&3��k#��u�}��C<�T}��kCˎ5	_ˮ �I5h2��f02bx�Pt�,��b���OI�v���vS����'�@T�|��R,�Q ]�h��X�z�����=��uíG=���{<��(��'v��8�b |rO�V�
���;�+�i윆��<�jq����w��y%�n���z��-U�P��Jy����b�:�o)��-kE.�N ��j^\,�Nf��vԠ	��UnßU�O*mm����.��pY�F��n��5�{��1�!��`F��'χ%�B��@̍�NF�Q�a����<ۭ9�EWk��A#/��|�s	��K�ӳQ �r�m /\����V����r�T���\����عq����ˡ��'vʭ�w/�j�#�N�\ U�������V�՜0�;���h&��E�� ���2A�(Om��t�,�ҹׂ��v����Ů���G��ё_g���diU�o�X�7��l���ޮ���v�䦥�ŕ�F>jT���b�VZ��v��0�\(d��F9m�f�,W�h$��r�n�|AJ�z�o7�yN���W���ߟ�1ޖ��ä��T�auEk����j���[�L������i��U����� 6��*���²�T��`{r*�4ۤ��Xn���/EJ�Ǻ(v��:zIg�F��U\it��s��ۖʖ���qC�g	g�pn1����>���pq2����nqd�	���c����`3����Uk?\��y�a���w*_ol>�Ȓ�W�@�$?�*�zۥ��\�(\*�0\5�ь}'[��p�a�y�%J{]����T�'�F��À�.�2�"��R����p��>+<�qe��M9�m��7;w�'Y�;�頄��d�� b~0��Z^d��B����r�&�q{Ti`t�>Xj��s:#��;X�n���`��S$��<��4Ŋ�17i^�F�7�_-:�4"樸�Ƨ���71��3���ր��$kɂ'�au�:�<�案\!O�g��*=���ӯl�7ʈw�|jLT$��)��|�FEB� cۖZ��o��IK�ј�{qP�_�|
�KhT��R�Ɛ����U�Ə�g%Ir�\��65�umn`[�v�	���dԩƎKf�H���¦N]��h�;3���@ۚ�6m@;�����h���!���Y��$ٷ&�҃�j���n��އV�7���>��f��LE����*ᗺ��7�T�L�2ۖ5�~�Z��(������N��D��ZO:�K��OΗ,yyH`�5e������39ȅʮAx*�m��㯵�`�������K&Pc�s�u�/q�5Au����z�$s�f��;`�߽�;'!�>�G�a�[v�x�ހ��1�W��;)�Nu�Zn(��E�Iv*z�gyǚۚ+_;5��u�g�DIc���<��vkF�#�.�����{��|v�X�`M7)�3Wܔ��zpM���(cj"~��\�b�&^T���n��ְ-.�1[�l��5�-�n��y�}w��\x_�.�y2�bc�(o_�:Z1ܦ{>�\�3�-w=Zwx�VE؋\���k�r9�t�� C�?.3�Q�]4�7M�
����,g��2��*����<�`�N��y+]��qG ;�D���GǄ$��_Q�������J	�-d�JU<9�,$l���W�w�R�,�=Dd=1!=�o�P�zr f�G�T9U/��q�_Lv:t�϶�u2� k�7�����*���'�3i�Դ��Nۮ,M���v޹��<�fX*��.��
�\�u�]�k�O6�&�y�SiwqXd:��}�{W4l%B��}sx�7�ׅϖ<�{Vz����|�j�������J��FQ�Z��Sy!�*����n��GY���1�s��玤^��F� �΂4�G� 9	W���`��MN֧�˽����3h������d*vٌ6Z99���n��~,o$x�h��a��O׭qj����ˈ%dМ0���(+S���C"�e��)��'n⌇O��}�;g<���Aޝ����}ग़t��E����m �*!����2^C2��B�]��o65��O�$�	`8ފ���OITh��N�ďa����+�o�����ʱY;=�c�ߣө);p ǫzP^C3Cl���OP?-5&;�}�#�y;�9�{Z��N�����ɛ\#7z���&��A��n�s"�P�+��5���׃��P����9��J��J<�E�Z��
�xb�'��k�bV}���9����c*1��<I��bb�o*�ݏpo���~t���������}o*����/~�~�!�m�܈zPJUc6�1�S�Q�@k��X���7N@b�`@v*�A����t�R���&OP�o��^!<B�6I��0E=�Osx�֕z�0D�ј��� ïz�M5�\�3��Cp�N��,.X[[���aɛ`�ķ�pZP�B�z�.˖i;}��2̭��զ�OF�L�T�{F�p� A|��A0Q�b=go.)�]
���]�!z$�7�����aw�1��+�fJv���ŉ�_R�Xڠ�X�@���֥�s��&G�vK�KY&OY�V�G����WN�
$�C���W��
�9do�q�V�|+5�Oy�[*��� ��{pقԱ�eh�h$�D�L,��Q��k���Zņ�fj�}cP�/�P�8�==�RY|ph�6�u��e���(҂	% �Gd�4�E=��gL�����9�|i�0ZZ�#�5'J�����W�����˹�J��ڗ8���l	u@� ,��~`�N'\8c���sK��q6��O|,�0(:���S{ڣO�»���F�A��X&*�7F4<�5	.��ա�]"~
�l=1P�9{�3��r��^�xl{| ��Y�#䍳�F�s��w-�#�)nu2T���y����}��f���0	�N�)�3�=?*=��k�u�b{�Q��#�[/=��Qy�o�����L�7��3T7��t�=5��C�(5n�U9�u��a=@ر
���a�&�v3�2唫_�/$�a;w���TsZ��!�8�Qɼ$�#h����Rдv����EnN���	����WU��f������7�lǑA@�Y}�%�5Ҧ�heԫa�0ǋ!�pk:�T�v�w��)���Qټ�I'#�����<9ח9;�1���M}n\���#����{%b��^���sέ�5�6)�b��}h�Bҧ���0�����%m|EKy�o'o��ɺ�r#VR-�N����A�0���`9�HX�QK��*|�2�oV�Y�^R81ؐ���Uw��w��)iU���_Ś�R=�u�U����E��^*Ҋ3�5��õ�x�Z�������p_��q��l�0���k�?7�隧�0�WftY+��M��J�n��@	�櫙u�����3m��*1��<2/�$,7]��3�z�1���[����&ղ8�Cن�t�f.�7-���_�p�w�x�z�:�A7K�ey�e���^l�S�0X���ʩ|�LP��k�>|�i�v�W��*���S�p��$ nί<����R�>$�+@_!!�U��n������5�᭦�>&��K�g�;�K��m��{5��]�)�u�p}I�R�|d�2���Ug���*!k늸t�8(v�b��;q���wRng4D�Z�vE��ֱ���u�9a[��ׁ���>s+1T�e����&KDfĆ`�3�ګ���V*8@<P�4��ٷ����Z��:I-��[*�ô~[o��9zh��������墲��J���2��t��\15�fǼ�Dֹ�7Y��́��WDm9���B�*k���)�o�V����Q�����gwi.�E����s99��Ϝ�`7�n��U�%L��1��@<X��:�!�dKf%Ջs�Ҏ�͍ٔ�cR�rz��[��Kϑ��:�H�y0D��.��_e�n��%Nsgd`�LX�Bq�j��s�zfL4��%3�����] YP��z�ۇu���-���Co�,�R:�k��]�*�7��޻B��yO7,b��jIBwm$�ov5�i�j:/�ʁ��\�r^�4>���B�<��lp�0/����ҙ����������+�j�����WZ|N:�X��Ts.����*
ca����7[�9��i�U��C�2;	��b�5�]��;������^B���&=J&�$MFG�ɥ�^�݆���1T>�5̀C��7��_:�0�Y�$��p��J����Β*�����O}3�X����l��6�;��,�3��b�o���^�-�v����l9�wdf��n��TJ����ً��R�\ڗ%,cze��qm�<����mϭb*駒�[�پ���%]z#��&�˖e����cí�璕 %=j�8���e�y+��WV��z�����M��ak��z�o�of�&L�wH�te
˸(�!u����_ ��LE�r��u���^�昲m��{2[�]��JvZ;���g�
���uM)��+���R�{��>�
�;��Z�jN*[�^��n�&�na�j��%��oO�b��i,���C!�>b�Yv��
�>��jr�˵�$��oJ�x�7�C���Fw�����l�J@	�Y�_�]U���ޕ���nv�o>���i�U�g���f�9�rDs��y��o�R��0��$�����Hף�V�[�I��<�xTe�O}�m�Ȁse���cRn��û�h_���Cc�����މᾑœ��R�g9M���q�<>͈K��2!�VY�-�����0fR��f�V���Z�5�~⼏�#�h)f���q�����;\��-���$���k���m��g�ݫ�q����	*ꕗg�@؈��@�|��^hCO��F�}:]'�;4龬��N���:��� !����+�cl���E�c�~�,��O�t�=��ic�[��)A�d��T�~-U�|�(&�;�!�J��]"*zZ��v
���_�onrn��`�=z�G��|��m�y���ts������ɘJmbX*H�����]N���L�y��+V�+w� ��xS���e�y���pY����6�-�&䌲�G.�J�z$8����=��@97�EKn��ϝ�BE�R�ly6-�+B����� [����e.���ꖉӚy�֯낦��V��e���)9���&-V��p�������m�4� �ٹ��ʖ�>��&�熟��Yf�3��uc�G;�`��n5#������(o���;��4Tf�|n<	��_4��]&V��]�d����Ӈ�^H�q�wm1z�]#�g	J�7���<+�z`�Ѐ�$��8ؤ=v��$��wӎ���q.�1c�k�46�֒t�Fx���ѯB�R�Ȧ�Zo�Ҕ�s;vl�����],1�v�{pً�j�앷�`8LOȠID�+��m
���	Y����.<�fI�Ĝ�H�J��Ie�φ�Ck�p�f�p,W�B/����4����Ew�-s�ց�\w�����DSu�e��]�q8y�q����B�ĵG3�:p�<�V�'�Z���A�|d?@0�O=��e����p�O%�W�i�6�]�Y�+5�^�T���Ciz'���K�/M�Qo��L������1'�f��u��j�H�QCͮ�b <���ZS�QE=�}j��bic�n�0�c�c��t,���cE�歞�v�`$m��j [N��-�.��W*j�*��uo8iY!�5�L��
��eLu���b-6��6շ�E���2�֩�t��{ɼz���,nRAX�e�����9��w���V��IQ\��+[��o�[E2(K���m7�e�������yV�32�[o��\{�zq$WZ���=�,�"B�޻7��1 i$AE��َ��v�8h)���efG*Xۼ �����<.�Q���)��;U�o�U"��fl���%'*˨f�l�#a/wU��;�N��Hc��^@rkZmJ��[u�y}N,U/`�Hc���6a�8`n+*��hK��觌� ��ּ��.���w"r��V��݊� ��XPE켊[C�mt� �n���QP9�[NX���h�{��R<��XF�C&�;����+�7�/��Y�5�Uu�j8��r�!ݣDq�t8��	�h�]�ʻU��C2v.J�5�˨��A��݉A���G5�^���t-b��pc�P�4b�����J��	I�4j���h\����n-��1�`ݶ�Q�W��,��
�/���-7�|u�Թ�tp�ܳ3vs���89��\s��v���\
�/UtU��vQ�΢�w=�����:�`ώ*K���b��р���D~3�F_�=6/x����fNzۧ��m����d�ĞTjR�����I[ܧ7{b��ۡC&$��
1��P�y���8n��F�\���^X*��m4y��5l�4�.��H��X��|�a\�E�圮n��Rͤ�n��\�\�4K�H$v�s�|�{��WR�a8o\��سDj�_+�S��>J�鋅�
���_e��b:ĕ�AMV�8��n^�/*0��gS!�8�$6�D@�kc�tt�G�mw ,Ȏ��2n�����a޿��
ԯ@�O�Y���q�򦌩���
U:���(���x�OOpL�0O�t�́��f'[M3�n���ז1�j`���7K^=q�'��[H��=7z�Q��c���ĵ0�wf+����U��޽�E��d�� �{��m�	2u
*<l�Gම^�t�E�)��z4�̕��T�0�a*}��)��*�+��I��m�r�H7E�b�u�u��sۖcru���&5=�7�I$zUځ��f��(��A_[mqᶪ��\�t2��Q�&�ͅ��`�o�f�Ǉ0DX��/�L�^�����+����ON=Ӷ+�j�v>W�N�{�?�&��� u���ˍu�2�X0���u���f������F4��`�R��\��ib�Ź:B��\u�Ͳ��$ɤ�e$��=�/���e)�J������`o�_"9Z�T�����D(�#�H�(�DĴ�&I��f��TEK%�Q��*��FS4H�TNJ\�%+S�p�@�0��Ь3�$l�2H�r���QF&�!j&T�hȨ��:�m"ʪ�$�s
YRsaT�:KN"�p�͢�Ȉʴ��0���&��"U��'"��EL��T�ʢ*��d���ej�R�AUqBE6PEi�KP���Tt�b`�E�h\�dF���"�����U&Qv�QY����Y��PEkK1UH�J��kR�5(�2Zµ�+4���0�B�8�T���������M@��ː�e��M"U&�,QB��Ԩ�tْ�E"!JI�΁R����PfW9VHb����Pb�D��d�9�Z�i��I�� 6�k.m@N�a���t������T�YO,�5f�[j9Իz���l�wkk6�@+''}M@c�u(�.��`����J s�)������_������©�}�ȡ'�97��ul�w��h��$����t|�m��o(r�1�S۵�7������>����%�fDd"'w��O�ifD	�_-<.�����u�����,�C�CsS���fr@��$��d�y��x?����]�=u��~y�ĕ Eۈ4�Yf�A�-��	#�iNM�<����r{C˽>w�®��FON��a�vC̫�e>^:�`�C(��N��4�?%��'M�5����k�/�	7�$���������C�=&��|8\>�s���|Nw���ǅp.<}Oi��ט?.沣����qժ�r�,�E�����D	!�n������o;QH`I,3{`	!���>׍A���9���ù���\N$����q��򄇷z>x���M;���a�s������R���9^*�ᠹ�1C=�9�Y�i7���x�m�ܮ�{w��7�/6���ȶ��\���CQ!�-��f�8@rW�Ă@���{��93ȳ�#���x�$�Y�����3���Ѵ&��]yR�i�W7��ɼZ �;^��Q�	��}p�+��������󿝤���x��9PO��A�x�+�(0E��+ve�����]�������Sz�*�M<`e�2j7ֱ9�;`JP��q�E�̱��"�$5��
�9n'8����]��0��8�\�8�C����<&_��ېP�������?�-��6�dY�����`	�G�؆n1H0E���[���O��fu���g�5�-%��F�}0��K KMs���<@�RZ���@r�C��n��aw�?�̟��	�]��M�	7������L��i�E�!G����{̚WQ5}�3�Y�����x�������}���}_]����7i !=��,���̋W>��巗r�z<�&��y7�/��!�\�:ZȒ�[�(qXI��_Wa�O��R��V]����$�		�w������_W~�iI�3:Kg&g�K[{��0$�řj�@r!E����%��"�"��"�7�����Ǯ7�<<��ʞ���P��8o����]�h�Uq<�+��
ih�7����tӉ�P���Y<�N觻�u|r�c��WE���u�Z}إZi��/QG�G�}�c�n�LO����x�l!(mҳ��e��I�[O
��3���K^H�ِ7�S�����"�;QD�_�B��"�Xp�"6"`O�,Аn.X���f��qD6��@[�2t�y�C�Ȏ,�!��>��An#�#H��@��P���ӏ�s����I���fr0ol�!��;��sQt�3��"Ο��|vSv+ ��9�����L�p��@,�̭�m ;n��6�-�0$,�Dn����@��JZ��%qlNG=����j-d!�'�HI�����7{��rs�	܁�'����nM�I'���pE�����������@��Y� Ia;7E�Y�kn�k O&m,�6ݛ�|>�Q�U;wy��,�r�\��<�A�-ɽ<�?~�����0����?�Î!ɼ�(
({O���~�.�����7�	$'{w;��n���}��S[2����@��t9�.:��˟����9��-E�:��#6-e��8�H�frî!����#�������}�ǋn~���:v��^r�j��?2t}��{v�7��r�E�G�x_�ذ_�J��������`KIX9Y� I	{�4,4��GC�Z��Y���D��������7�'I�~�����xO��������|�.��}~>룜.#��:�'yA�ɭ;3�OU��1����M�>'!�5��X9��� ��0%���w!�[�A����Ca�@Dy��q�s�Sk�<�{IĞO��yO��&�/G��4,-ў~����M��o5wތ��S���o��������<�]-�d�ibf��Zrݚm-e�o���n!�c�a��!�67\ia�x�s {y�A 	���wi!���HB���W����_]�;����O��cӼ;�n�c�zC�aw�<�}A�@r����I-E��Ba�AY��i#¡�H�f��@�	�}����=0E�ކgI��6������AޭX�>Me��,�d�g.G5[�	`(�#��@Ih,��փAߓ�r|q濓�aw����^8���90��x�ɼ?�?���͎��<E�n<@B-e�Q�i,�Ci������Agj->�\LK9lV��,A1��翼ֶ�(<���ѕ|��T�,��(z�,���w>�f�aý��G��#Y��;hb��ۼR
vH�ys���8����%@ZѝY5Y�{	�d� ���V�e�/s.������.s��ϔ�A���.%���}���yI��� =w�'yv��h6`�������̈���Q,$�D�zpro���8�Wz�N���rz:=��<�}|;����P�o���Cx��О����z��{�u�����U/��HE�x��4Y��r<7\I�dO&x_@i I�#ژQ-ř�7�Q4E���C�o�.��w/����<������G�}��(/����K3�٢��k����=��s��;�i�9��'��	,Ă@���0��L��[�@����z�m���~���I�S��vh6� �g$��ez�
"r�E�V�/~�G���+k��������	�\
o�矎��ԡŚfÄAZ崳$�i�sH`I �x!��[�2t5��%��,�-�D0%�E}��"�@r� 4f6�^]�f�[��ǔ9˳�	2�O���x@���8�Gx��nM�	�y��?S�w�iE�K��T�Ai,Ȏ!��W�����|��~O.?8�޿~�xF�8� ajɹ�ǎ�|v�ԗe�f����������{NL)����yw�~C�zV9\HI����~�q�q4���y����3��$ q�����8�H����m#Ÿ�"�yӻ}\�e'��W5�����`��Y��-E�����5���XCqk._S#`�iĘQ���9�����99�?]�	�]�QO��L?lxI���܁�q�"�ə������f�r&���̒�7�CIQ��6�Q�j�:Y���X{�Đ����eχ[�-�����w���I�\
oކ};rw����N�m����x��}v� $4�bCI���o�=�wvj�fxYD4��Qf�>���4�r(w�i!�-$y㡃�� 9 {a�[�dp���t�C�OWC7�E�����6�g!��6���'H��&��"�e� �82O��dE:��ͨ����poE��$<x�`KYy+�{Oi�?8���7�������q�+g��@��04�Q�An-�"��@E�����Dt�$I���$/RP=I�.��|]��fƼ-5z�ؓf��+L
�2�M��+��_�D���T�]J�H���|��ӜŬ�t)�ݮ繽c����v,r.a��󲜣�܄��R[Ad��ָ9G^綐�6�
�mY`�k|����tɶ9�/�b��3&*r3/2u��C�,�[��I�94��(I�$'����o���]�����x�:w��ɿ!}���ݑ%�$5ѻ���P`��\Ci���qXrw`�Qa�9`�O�)5�u܇������+��0$�bA���a�a�oA�w�}|&�O���ӻS�b����hwY� �@r�)��,�Ih-9n�m]����p�������%z�r�d[�8�Op,�dV ��S�Q�Gn�;M��:k��9�c&�.��y`VU����j�hi:�7X�������\a�LGK'������W�:�*���m���	���h-�g��Lh�ۨI:�8���ؐ�g��l9�1.��xT
��	�R���Xԗ�/e.򓳾���e�����<�W�va�ⵜ��Tĭ��;�s'��9`&�p��g۞�3��&�������g륫���/����^�z��\AN��ߛ���>9K�ʕU�/z�;�Q�5�O��5}�	� ���"U���@xX��[9�!�-�z|*� �������z.[�t̻g��>�g���=n���tW��\��([�K���#(�cxU��]+{�ˢ���J�,T�^pxL�]���۫ZI�ў.�U����w4ΩW�M������k�\;��g�S/���)�**_]p�r��tr4/OqCo�u��q^�:ܥ�:Է�od�٪��9��z���9��(�6���ۏ���u���u��y|�s5 $�_>��r�P	<��̥(/ ���/���{��_Q�X����(O���#����a�چ�/��c��[|&2�I�P=��2إ^�-F7�f��$����Ѹ�P�5�%o�D����םP�|\�/>G�9�����TpVv�JlAC�P2t�y��㮩3��|j���%��;IҬ�?dN"q��;��X�s�խt���'���� 9�a $�{+"8�P��Z��C9��������ܻ��㩤����^�ճW~���48�E��B3�3uL֏d
��.�AE�t�&4^��pJޮVk7sԉ�f02i�Z�ǑB1�� \h�Vˣ�W��)�F��ޣ�)��U}!��
�Na��6�y�4�,!�/7�r�g���#гЌ��C���8
�[K2�S��v��>���I��i�"�L�=��#8�`wL#��ꐚ���ԅ����2�y��_pp-5�yp�����~d����;7t6A����v�	�vf�˔�eb��\&�Y��2��K��k�cMk�t�4�+G	���~P^�G:�$+��Q%c��]��u�r�ɶ��s�=ViM痊��Ь[~Y��)z�ם
���@ӯ_<�iNB�U�Hs��N���H�^������P@�6Ӈ���%q9�� [R.O�s��Z�f����ɠS��)������t�59���
��n��d���9�d�6�08|W��p�k`i��-����3{w�:7���9z������X�������*�	�y@[���/�Jd�t;*Wl5��&�%��X����-L0:
ke':#�����1ql�0���k�h�O(�z�{=�ͮ��"Sˮv̈��9.\�ʹ�[n��G��/L�zb��2I��-����oR��/P���.],��k*+�	��`��`2��r�YM��pP�"$v�����	vr�]�NH.�3�H(C��Ϫ�򜅓&��c���t�3�Ns��uh����պv� o�����~�c�W$�Ep
������\kn���Р��`K��5�FlU[�s�[�Z�Z1�M�nc��P������}��a@��Gg�T����b�ݹ2u\�D[m,�)�+��|s��C��{0F�9���)�����0JU��l�B�}`��s��W9(�8�#Q�{¾�I�G!���|�k�m�n�M|�IB���\*���~kb<�&��+|(,�\�U������`���~�yO�1�f[ƽx��O�B}<�*
uv���5��	�-��!�J���ָ�5f����t�d����h*�v�%)msP� �k�����A��;� #���f�Tx�"����)"��1��[�m�pb��2^D#ZBu��o"�dl�ʻz��nF��;��0�3��0ө���I�G���h�|�vd���F��J]*���i��婮�Q�^�b=gQܠ��`�5k��K����U�/�����{͠�9��;/�pM���;}#R�t}�_AVz���S�V<�]1z��W�y�,#j[�8h��&<��;^�Y��=&m��wlW����b���nb�s����z��j��;=�G���j��؟�MP!��f�[�I��J��5����e�U��Heŀ�OY���t���;�o%>��X���>�x���l���\�� �-�����u�l1xcE���a���[v�-\u(���ˣ�✇�pvP
�mDw9�X*)�e��<#6$@�2k56�_]m�$em�k�D�b�T���
���YK��,bcҷ��C��@�`�C���M�Ί��[q>~�.�Ǡ5�ҏ��ߴ�
���ʏ���)
����P'��v����kO��_��+RMRk���@%�ՇPW�N��ut>K�i�cݡu$�Q�/p���Lyᗝ��뿂���6o"����C�xƖS�c�|Gnک��f�f9���w@��ކ�<�rh�c����v��e�A\�x�c�Y���0��m�����Dm¬��ʗ��ۅ���C��燢VWJ;�<IUc��M�7!��a����ή�\���BhV�-d�P�SÍIf5���=ꑷ=����I���V`�V�sG��n��h�}�m�Cj=p�>8�����,�L1�z�#�;������"-$�C�v�d4r\�����(��d��`��dH�2���7�26wP�+�~���u�*{�Et�f��&�(�{PZ�Ԏ�Q�*:�tL_��Sq�a\)���������0)V�^=�V�,��\��g}?Cn��_�˓đ%)�����^%�z9�Ty�)[�"�,�{K��(���nN��2��DV ���k���;M�c����Z5��^��f��ۏ�ܛ���
�)��F���a���`ih���6���,�vum��X��2I�3�./�ٌ�P�wzsS���F�25�s:!��bms�ld������ط�΢'�����;���u�Ԕ��	8Sǫ=w�A���v�_0�|HF�t�����!ڕ�q�����oJ�K�ȇc���Wא��*n8�4�3�t���WYڣl�s�x$7�n�9{x�H�G/ik�n���`�����C
y�n���#�S�q;z-v�)�H����:��n�-q�
��ԉ3��;x�����UU�y�mOD�P\0Bi�(׆�H��j�3qpO=Ҽ'��DRN����!N��� 27o�t��pgXo�(k��P��Tn��^â�ڸ]�� �s�G3�eLUv��8���|����\:�N��6޸/}���8O:��Q��Z]8��kL>�jdVf��WV+�/�
�yo�m	��2Y�,��ʖ���9�izIR���������.�Rc�+���9�W�S8�b�h��Pق�P���Z8M_РIVu���</�����9\�P��o�L����D�g+|q�,�*��S�a��؀z�n��o�gN�%r�����J~��b�*��)A�	k���Rt�/.i��쥔����(���Q&]Z�aW�c�� &	粲#��\��r����+��
7n$[z�nvs�tx'���&����`�&p-i�n��rt�׳�t(�ͬ��6����Y;۽��!j9�(�f�z����F��-����"(�w�	o��`�[�uM�;��>NX^j�|� �z�׸�8�w�k4���6�XsQK�v�.NZ�m�<��)����QT�f�:MT#�R�ܗ!ӻ�ˮ���iE��z�>Z34���S���讐�.nL	�S�u�ʱ� ���� ��{�؎W����W�v3f���>/vd6�.=M���Pۮ�5p�`	ݰo�8�~�F�TV�
5���ոx�����N����Q�7�/��N��O��JS&M�?{ ~���S��
1xX��Tjo+Z�r�NŜ��r��P���~�n��8�꺅���~D���:M��5���r`���H���`F�Ux��e�[���Â��l�^Ogh�Bҧ��$,��`|4���{���T��&4��E�ܻ�+O���ٮ���lh��˯�k�l��`M��N�5YJ0F���O|�V�X�����ĕ\���EWCg��m0�^��%D�~��=���uq=�� &>��<�������p�k��,��f�n�"#���]��O�W��ݍ���#U�Y�(m� )9�/b�|¿������V���
�8��,Z�Ԭ=�ĳ9�L2l*,t��cb���u�T�F.�7-�.~����zt+�n��#����`��V+ 뢪 xWIG����Wb�v��ia�v4�X�M�)7��Qʩ�r{�J̗&��躏7���6�b���s�����NZV�;���Ia7<��V�n�J�Y�N����uT�m�,�*J�"�j�p�b� ��-U�O5Z0���nF��g��"��,æ�uh](�Wύj���e��ӝY���9�Z͙ K���Uv�)(��R�v�ZQ�3�����	l)��q�kn��������y`��&�4�(S�y�*^��n��B4-E�R�G����]��-5-ѽ�b"�x�得�Ҋ��/���X�M��d�<��8sq�=o��L�\1t[G�μmp
�&Hk[���v�����ԃ�+n�*�/�҆T�Z7e]+��p�<��yؖ�K�9OV��R�2w^$ݹ�ڷY����)Q�+Q(�ْ]���6͋I.%�t0w-�;���2�P4�\�,���[y)?��4��r6z���.���Ԩ����3��[�*Z9��✭�:/�B?����^�T��+�^J�ol�T�v��6�@ޑ �����
=���݆3:0��|T���u��+Yb���
wj��.Bu)tLЮ��oW��St��t�(sU�H;���s�ȳW+�6�K�7��>�t周]�.���@�[н�vq���)�M�{��;�V�u�n�����Q�k�9uGYm�z�(�&�$Q_l��b�L�=�8���:��;{�}:�gh�0���K��,��-�־�Zk��#M�-g�z�f�x+N�O&8\�@!UhPt�����_tv��M�z�\�W+2�N
9Xs{7hS��)}�j�3������#*S���*�*Ywt�fpoX�RĂ�/(���=f��aZ�Jwki��A���.�WJv���$��VN��`VR�����	��1}�wt据=5H��q��G:3�4�����G�;8+4V�s�aW5�-"\�	���v��@��J���*�)J�69��ÖLiqȇn̨qF�)���H>)��aË.�>1�r�=�+�BTۓ�s)J���o���G�A��4�o@*��P���4�E�"k�%�j�=]����0���>[A�b"?EOV���c�nK�6�s�����cz^��k��4Cs�6i�wM y����Eú~ۅr��J��3G$q�}�	jX�Oe�د�y��7#΍usҞ��Q��"��r/����zYPSh��7�m�՘��5�Ƚ��=�[b���T)D�J�*)=ɯ���}���4i�ɛ�vB�c����Mvr��F�(��faܱ�k*[�B
eh��#8��%z�#u�>n�L��u(�d�E�g�4ݴuk	ѩN�̘�����7"����P7�w<��Ć�ɎU�b���+�%Ӽ0>-6�b��%w�k���P�K�)���-p݇�{+h�:�I�j4R7;��t�5x<'�3�YX��g�BbS
���JXD!ШU6Rar*9S.�I�ͤ��I]��t娖�d]dUȳ	@��fcE�G"�D�����q$ډF�������
40���:��J��L�TQ�2*�e
�����HU�B����H�a�6P��q+E�F��ŕ%�Uʈ�(�I�(�a�lL�qeuL̖��"���U�DQI�i�!�)��*Μ��EEfRi��E��Pf-(��Ζ Eʢ#��)K
*��V��Z��QfDf��)YV��i�&Uh%	r������� Eʋ�V�b�(��2@��UW#����F�Z�l��A�jHIPh�r53,�ҫ#��֥�R�f�'J�
B�%���(�	V���VM*�TTVu������19fAreUFbfHȹBeU��i@�J��"����=y������K��QQs��KGD�d�XDV��e�SPД��*�ҙ��.��P�W��˫
�tˋz�v�W#������V���f�b����[Z�,��	:��CO�^U�ֶ�z�����kD��V�_>imM�JF-�>:��A���ν(DB��LEV�Gv����eJ�l�ր^R��]P'��]���N�7/�71�V#�J$�ϸ��Ɣ6V�a)Ӹ��OR�H��-/�_$�"��膎9��nw�w+��'�<*�dw�{{��Һ@�D�xX��)��ƥ��6�Ex?%<OJ�43^�OL���=�e�����"���Ӯ��wM��2��1#��nO3�䆋�Rb�N�����Q��C̥��y���[Q�����G]� }f�v]@�/Cp��fy���`��F�Y[�n���׫���C�Ј��/ '��2�Ս����Ct�G���qE{٥���{Uhf��W<(?��Y��7LE�'A��,Ps�ىS�Ч����6=�w]uk�p��VX�ڸ��y-v.Lp��ћ}l@�E�A㪃���x[�THˏ���lH��+�IeGWTw�,��-�ֳ��Y߫o2G���{%<ɫD��Fv��A�h�&n��2Ǿ����û��fK���n��^��I{���)>�9�s�k��S�/]�>���[Ցat�?��e�ל3��ປ�ִ��D���]'����� �U�eNｱ��
2ǳ.�7���C��T�g�ױrs�G�<_�&���kT��y�v�R��rP�X�K/�ST9}֗Y�����.�mDOs�e���2�����٭�8y���F�p�}��Z;B�RYF��ھ^t�:�Ec�s���0�s�����p��)��@��]�"�� FL��3���_��,a��bZo�ȹ�v��Y��j�c�C!�c/�{P�����epQd��B<I��Hzc��imc�)m�����)z������EL��r�gl�����B�j�R�W��j[e��fK 'bE�]���X-v?-s�C�;
��*�G![WfY���;�D^�a����HU�V�YN+�"�!;�����+���C9_D�!��@b��.�5�ś�F��z�L��"(޼Ґ�Sԅ��i?%;(�M݇�����Q�L��.�*�˅Tqh�~�Ǹ�{@͉��bO�o���9���<ٳ�"[먷ts�<Tu�B�j��=�Ug�Sk�q����������Ń[4���j�C�g	wR�ds�H���ȫ�-(��.��])ܬ�����^�W�%L�ʺ����S�%N^Ař{[��^� ��D�×3�B���[�XzZ@VV��i�{>���6k�"L%T���f�>��3�m{si���Q�q�5,��@jqDF0�DLF��P�6}����\a$��,�Ζ��d�J��|��ϓUrn0�S��io�'�GD�6��-r���2���S۹{�Ŧ9*dr���-�3\%�2��Qԝv/���lW
�]͇�g!�k
�N���6���#"�F9���OJ�T�'M��3�S��%0�Ťⵜ�Tĭvv]�
��зke��S˦,&]x�5p�B(.�|~��j�3qpZ�:��ꦼC"�3�i�gc�强M���N�'��p֣�j
�M�y:������p<��5��ͯq>Pe3��y���J��鎸n��7�p�k���8J�~�0N�,N�1U��"��3+;���+ �a�!�2q���˅OR���:�����-Ⲭ3��Ļ�:������&�9B�3]�H.X_ûn�-S�J��C���{FxX��7x��zO'�`��T� ��D����	����܏�:*uݷP'9`����C��艗^f����<jza׵����OkV�m�hF�l�y�|H�i/q����V*˯�h�E��m�zPʏk�^H�(H�Ɍ緙����5���YV�쉶F��\(_��:�����-��p�z���E��*��T����'�\���J�v���́�`������}uL_ҕ|QA��Z�"�jw0��S�������(�:�����p��h�r�^@� =��-u��P�Y�.)��;/8����{͆iQ����S��԰1	��jZ���HOǝp���9��Ya��5(��o�ӱ��� �I�h2y�P�`d���Q26=�A"E M҅�G.�=X���h�|��4�cJ����8�����[£n�d�ͺ�^|�C,!�L'v��8�~�;��Ҿw� �M�YV������
���Ҵ�I����	Jdɿ�t6&1Vmn�Yx�I">��1�M�U���G����[�a��t���[�z��<��Zs���W���;IG�n�=[-��y�(8h�Wm�X8W��,����:9e��}��雓&y������**-�0u��Ca<ۭ9|J���wMK5�Pc��q5���O��)�Pؠ��U/���iS�1��hhs�_���� 5�������TL�d9�囟ٗ�f����$Q�M[��(;�{o:�zm>�C�}.r�֗M.��n�Ռ�S�{ϩ0{��Ǻ�g�O���8ox�I�D՝b�"�8�`�u���<n�����jG � r�b��\�i�� ���:��`��W�k.hI��i-��Iغ��:��B-l�BN�E�=��vLTB6O���mMU�c����u=Ǌ�G����왃,�4F�AP`߱��U:�����n���"9WE.��RtJ:�:l%G-��k�=xU Q�˳��ec0=np�+o�C-�$�CFi�СG�*�Ye� |+��J8.�^����Lv�x|�>�A9y����םծ�Vp���;I���Ty���*�8I�T�����\5%KãG-{=P:�k\���wX3ִa�[�o��Z5ŕ�6vF�H���N,d`&.��=���q�O��Y�Mݞ�ư�쯐�z�✺��)��n�Q��������H�p�`ל�1����b�]��Z��^d��|����'Is:!��9��m�q��D��3Co[^�{1�&�%|����4�@�LI�(fF�L��5.�9���&�2�v��[��O/8�`ށ��i�<���ا��.m��B��U��vVڴiuel���YB=&����Ɉ�sӒѬDq�vqR��x������̢�,,c7�3\;F`O���x��V��Y|�۹u�����9��]������npՀ,�5�����ꑫ��@�1��^�Ա��E0^P�*3�I��ZS��댾 3 �meU���V����S�[�ď�>D��㫒���BmF�R���M��&P��Nr����>�w"�d9�nX��?`�2E�c��e+��k�Pzأ�Ib�_>Z����4_�j�Ws�"����(9ٶ�(W<�Q����ĳ7�����O7ys}�R���)�E��q����o�<4��!�s0sc��𿟲�Fj�^��Sr/s]��P8k��G���fq:n�*������@�,c=���܉(]�d���a�9ݛkr��0�yח����v�w�8-��ή��>fy�1�m�Zd���������^��+��jf��^Z?1Ri\-����1Mre�L{�e^c�wI��:�$����5hD��3����*�}1�,P�~� ��r����>�2V0N��r�i�
�7T!��R�3��a�����>%\�Q��!d��o��ץסg��97��N�g=k4�������j��^������ޤ;%���%%"��,:�XP.��b�՟0=�2#�3+Vw	�����q�u��%�6��8�׸n�|��i��Қ���v|َ�M W3�[R̕��8��4Cy4��Ի��5�a9�wZq��j���M�ھ8�u�U'q�G���k]ڍ��0�b*� f���W�������ΰ�Qg`l�I�^�ܑ��0��$F���fe���f�]t�5���l��:�*��&@r��g�p��-uñӶ�g���Ӑ1C�+�8e��3;}�J�OuR��o�����$[�M�x>a�O�����Z�|w�܀)`�����y;�C�<���@#5��)ͻ�@�;2BWx����rj"���y�t�����EvRi�b�����3��Pۮ%�2��DF)�R�rz��������N�vqk�[��s{�r�b�۝�$� ��ͳ�``���`ix��ۂ�Ê'�:�Eh(�ɚ�N��di��T��g���1V�B�wzu9�a`چ�=N�4o�]���ˬƟ.R0)����g�τ_u��pGk��3��Mq���{L^'���\��i��W�s��iM�����Cn��)�!�4ؕ'*ښ%N����ֲ��ow�����Z���9��'1C�hs���Z��0P�*�}�<'�����x۲�y�!v蹀�;q��b�xȓN�7m��_7`pYS2u���J&V��ɲ����ʾ�ǽ�y�C�W-��*)I�R;6����C�\.0p���'K4�4��+��:�ʌta`�p�o 6c}u��.\/
�3o�Ê��9�')�xT�w,
�Q�oy���'2�   ,��9��S���"�������g~~X���{���&-7���P��/_?vĠWcN�A��InLM�O|x1'��֥�[�!<,c[_^���p����W���l��+�Vo^k�nR��4B�@h7�*#Nz�Ƥ(��7pقԱ�+o�*�J���J�+��|��I�X$���$.�rH�%�F�B���o�CRYzph�7j2�Z�,�y���dr�Hz���gP<�WDA�'�B(�}ܾ�m�}���p��vWqu�뽚��&�{s18}OΩd��i�6���Z�`D��	� �/��S7r��m�����d.M,X�򚿭�g��u�K�Q:{�T�θ�⾄P�� <�p�G�z(<�hqNg&�q�;�gp��o� ГT��s���30���h��U�!�TBmV�h���maS�F��;�'�9o
�Ja�ͺ�^}ֆ�`	ݰj�.��;��I]�E�*�ɟ��,����|>�ߤ]�x?�z:!"�2zt=��ęם�.b����u��%|GKxD�@50tބ��6,O/n6vE
ή�]r [쮭�(���6�٣�3�b�C$�q܆�ݮz�ă�Ò�>n��y4��.��p2%]h�nW\�n�kk�V����W��N�sRޘ�<����z��|3 � ���y��y�OtO�;I.���9��p�A����^��r��̳N�!y~]�p�Z�1k������k�'�.T�كRװi:VA7�e�PC�(!�X*"��1�P�)��֬�S���=�U�ѡ�K�25� ��0����y�Zei�9b/��s�U�<�DɆj�qv&�a!�;a�κ�.�8�%O��o�����_��qؚa2g�WC~��̄��u�V\���?v;ϽJ*����&{[L����m'\#�O���k|���OȚ\1���giXKNYf]C�3�~����P:�@	�u̳�N�aY|c4H���r�iŴ����P��=g��0����M/EK�o�1ׅR��e�P"N����w:\���f(g�K�Y��_(�uOQY\<�
�LPckӖv*c��Iw�a�]���7˨��Im�����AR�`3������P��4TP�K�p
f˺�i!�g�6������C]+�o��04F�8s���8�Q����Ju�^A˧r���Z���+��M�*������A���qL�Ů���z�J�]�vm��RA�Q42�)J2St]��{�A���S�O9��Vd���2«��ĵs/�s}�Ό;���f
a�����<�9���0��o�����w�\�u|b���|�0 ��u��������gx��]���>��.��|�)��n��^�#Uz�AyU.̺�i�{���'��"��5�l ,U03o�����VEFV�W�
]$q�膎9��n!�r:��� Zv�1z��Ɩof��DNN,�{�4�?(����o��LY#��9���q�86h���y��uY�&{K�{�<X�%DBk�x�^:v�)��ʈqOY�$��S[i�mnr���a�޲�|�b5�B5	����a/����ڪ����-�3%M�	Gr�é� �	q���Bj�E�L�w��}$�N�1Z=T[�V<�] ^��BSة���tefg:I^oP���|4\F�����^'A���;7�P�~�����~� �U۴[i{r9������
1[�������a��_����{�����^��hv4��#THN�p�|K�G'����3<N����<���R����xɵ62����4�^���B�}����n��>��	�����Iفqմqp�v�>_}nz���[rno��R�k�'�t2�v�.�����N�r%O@t2Z�$-t>�VW���L���� ��B�NN�5�s����׶�|e��2^��[�b#��R��h�Ђ;�ޭC8�묘�Y�eG"�t�
���YLe�����b@uTa�1R�*�5U�V��id\ ��z�%�<���SVO(��&h�N([��S�GMf���/$��g�x����t�HRS�]��/���Ln�Ȩx��=���L�����=�=Jܸ��3O�J�E��l�y|��8��Ե�i;�Fe�}f��X\Q�7X�2��`[}���W5@ck�wV�r��|�x���E�rc��4a��:��ɚn���oB-�`��Sөq;�ԯc�ۦ���l{���Uq,����)�X��\��hf]oV\n*�#v]+9pme���t����\��5QΤ���V+�����+q�����0%�.g>yx͌��جŠ�E��������@:���X���5��:�lŲc�]s;�M�����s8�S��<�;F��{@�gg[u;1�1�(�o!�z�#b����>=2��$b���5����+9u�bȶ�Q�;L�X�t���`�p�F���8;�� S���,J���H��e�s���gq��.����	F�5�Z��d����������Z�`�w��*��u�hg��B�a�����mVJo!Y�|61-F�J˹�q�LN�;���R��t\y�:8��mӻiU�D��nq���(�5b�3�/�i ��v�L�q[�Nv�N���Gie����-�خ��U�:!�x�NZ͵���n�*Y98e[���
ǡ�l��v�����R�mRl�*�z�^:�#�����G�ݡ=N�:�7�s	�dA�/��ȣ���c��\�x�c�kq�oo%E��NNt�%��t��V��lи�����Õ]�[�um�-h9x��������h��2m:2����AR<���(���͵<� ��}+�,	����h���A8�
]�A$�D*�K.���T�2jTNI녒_]���|�I��+���;n����e�ț<�Ь�ù�b�\O��,��C�I���L��|"2a�ۭ��h �Z�Z|PEV$�:��Y��dX2�Q;��Np���yڪ,���`�/�Q�q��sr-b����X�Ǽ]_=�+�^������Y[J SZ����+�ظ�\�{�`�9JkB�ZЫO��;�wt\�y��
T�o+�͜hf�t,��>+`��'Yu��y����ʳB���;�YP��76����ܥ�N��n�T#ͤ�� p����G;UC7�cq`RZ�~�4�ͱf�\�����k����Ȍ�\�c���S��*f��efח,;Wl��������,,�s�<�l,XZ<�Q�}`�L[�˺�e��	����5)�CT��YE��ӄ�ڹk��D��L��J�
��p���Er��(�\�*s�r���̖�TE�(��TD� ��H��E0��)
�Z#"���QQEp�*%ThR�9Q�KD(��`QQDY��Y%�I4fͧ2�ԨԙG(��Tʠ�QT�"��\��%EȎDPEUА�UZ*�I
��s�UJ$p��J�E�+��p�J��&#�JT:���D�$�Ue�A�Ud�K9fjF�]jb3�\��Z�QȋS�UE*i��2���Vah��g�Ԭ�*ȫD�)*BBوuYTf�E	�H�!DV�S9��u���DET\��er��M4�UUkJE�gj�r͕�dE*W(�e��r*��p�!"�,�&Es2��T
 �V\R�g"+�E�9I��I �� ����SY�RiE����>3yV�9(t�L
�T��D!E�j(c�Im�1b�u�u���h��C\F�v�u�Hc}������������#R�
�S��ʞ��g�\�7�#+���Zx[�b��8α;�VJ�}�Pf�%6w7�ԡx�k��[Θ�Z��<#b��q�B_��KJ�-z�>�ڎe��Lb�"fg{gm�ʄՓ"6�u �	�2��0�"����s�1�aʅ�Y�\����F{(��+~�%l'�R���/9�2�6��m֨ײC��z�엷��!�V��g5lV,Ky]�e���ԞA��=}�a2骊FY�7�S.9�H���8�4�|���>q(�˱ާ�����_]��%_
�y�q����v:vٌ��o~�\�>[?q��R�
��{*����b�#���@�� ֙�L.5�{P��}\f3XȜj��_l�Rh}/��|�rՖ`d���p��� \�����}'C�^���a�I\��\�ܣҤ�>VG��~��q/>fX��1:c�W.O@!����r�Tt:�9��ه)ңQ�2k�ረ�yld&���"������.0�-eu�Mz&k��ܽ�yZ���������aYe'2wEͼy��Ɂ�2�X{WJn4:VJ��{`9f@��~[���,A1U�V}�3&;=�����V{x�2��nY]Nj�uһ��F-���
�Ҳ�O���J�UȠ.L6dYӾr�Φ+5�30a��s[��x�){���Pe蛏6<���WHeSw�����z�t���#x�a�ɽ0��3���-KL�9�ɖ!�����Oʥ����t�f����k�W�Ңj�dz�\�L������7.����As��RÕ=u�B����F�5��jx�k�&n. 6I{m�Zm��k���q���V���k+c�X��xg
��$C�U�a��[&�U�X������'P!�8	���s�<�d��{���<��k�2���:+�*�䖔�}1����gg�~�����| �3�
E�KطLB�����ݝ�#v�Ee���sY|�nI2\I�As��&��r4����]2n�a�u�Q-S&�A�\��u�ʞ��aꝓGA'k�L,�=S/��+U5�����k6.�S��b��\���"�O[oك��l~W�qAb�:`�0;���\u�u)ip2T���S�T���z�ʛ��R�|3���N��}��A��L@窄ʇ|�V��߷eA1Q��6v���*,vFJzoS��˩���˨�i��К�<���ջ�g[����)��!k�%ՃKo�C����H�R�#��|a����Q��t��5g5�� �Q��J:6HάC2��F4�/T}n�ID�}.��,��Q$g���7|����k����5��}_r�;��E|�uJi�;��>�E��&��l��OR���ZV�6�i\3��c~m�W�m�"������R�O)aжA�SR�2�ҝ}xm%��6�6-�
�˪�w��\�/&�c�䶆�q�ʠz1-o���od�N�d�A��e/������m{Ҷ��p+��W�h�ݵs�{ӓy���h�7GW��=�r�$u�KJ�rP�?_/V������b���R��l�� 1zmw��Bz�e__��یN��L�y;�'.5��o�f*8��Mؕ)\�B����fӗ�*!�:��vT�	=k���yήol]��Ev��);�D+S+-��W�͸�����*�}��2߫Lط�<��'Mjx_k��|<-��^u��㒂�O�2���UD�ʉP��(��{�6|Ϲ�lϡ��)��wAl��ލ����b�3������YVa
Ǎ��k�3�oC[b�0]�i	�^����b>Cj���u�#��5�����A7V����T�R�ܺ�8��ov��p��V2n����I��rX��vuF3%�ɪ~������~�نF���K�y]"����3l2ϞU\��2_\aH '1[iB�#iWvj�t�XǾ�NF|����>31 ��=t�Ue�DL�GV(�IZs�wW�%>JĬp5�[��_�C�m=�+9\
V��T�>��޼�c���T��:m�խ��'�y21ڌu��w)̓~%�>N�{����MSy\������տ}�O����/���q��63�3neLWG.yL���k�f�>J���[1� 7��'׿3Tid�7���\8�y{ll�j;����o�~j x�W�C�c����Ϧ�V����B�P�4��Gl�4�ޛ��k6�-��opv�D�v�f"�����o��jgyr�<u=o�ٳ�n���M��-4øeƻG"S���U	�{n�]�d=���2b��o���_�-|��j�E��6�]���}��~�Ŷ��P+�O3�"�ݝ�>~�9���kv�O?m3���y����w�+�+���̊�/%GR��BI���[˒�ݔz;�V����r�c*I[�2����B[��+�,������-ܼj����,�H�1�VE`iUn��T��`�H��ﾯ����rk�t�Nť��k���Z�"�m�p�[�v���j{V,��=��(o�6^��#"�@z�gVU���k�Eޤ�]�9[���ȹ��9ε�o�G����v���J�?��1�7�S�OY��Vَ+3�j2�Q��)<y�����Rk�I�{K��w��mN�f��{}�rP���V_'ӽ[���@v��妋���Tc[=uc����UK�9��T��֬}˻���a�+�cb��{���_����=)Ub�%.E��{r�6�2���5�Y���s��-����ކ�=o�%��_(���qeM+�D���-kz�eA�guIn�K�L�B����އ�9b��%e�����y$����';���s�w	������t�s����х~>>�Ҭk[tZ�s�5���{2M%��;5�BD3���~f<��n���tv_��a"0��O_���f�Y�F�X��oƢ�R��N5���K7�xJݦ�阣E���84�,n<�o��Ⱥ2x�չ�������F��Z�Dv�6�(+�M���gS��l�G1^�	�n��Mw�A
���͋mM��}o��Y�ff�'D����U}�G�S�<���Y��g;��ڇY�N�G��~W��k6�P�����?����ڄ�L>C8�6�)͹�E��W�D�=��R���h34���y�k�[��!��.e���\k�r'�튈�㪞]�K�������o�\�xsPs�jy��v����;�5F���4ۍh�6$W6��o�)�8�
/�L���e\�^��M����b����r��͑y� �&܇]��XW����uBN�^��t�s}o-�� S6u��,��v��5c,�F=�N�r�X̣�T$�O�zϞ�+�������g��X�wiu�/�OZ�u��;�1�N+y��T=:���u��<z�<�A������:��{
<������kz��F{�K�ؙ^=���im����g9�&9�U�tc�߆(�֚��h��ߚ�Ɨ�u(vV�k�f�F�L�l�Deg�~s0g��;ޥ�e�ͣ�1�s��{<�xu������-��Љ�ͿL����(u+�@�t���y�j^�1�Rݩ��-��c�|v�˻�x�;R��o8�]l�֝��.�*���w/�`JG��X7s�D�̶J���A��5�Ƕ�f��>�����pUd:|Trߡl����=��ͷ���`鬼�zʶ��R��=>����!�w�6�̸��H���Oh7tjͣ���'�^�}﹆�zyi��V	� Ĭ�ذ��.0ՠ�q*�����G�J,�y+r�ֻ����黁a��zJ�(���VĎ������+����O_K/w����}���;N�M"|�Iw[f���}B��څ�q�]�K�P7]�Է��$�b����C4�+]Ob����R��V^�>J�k����MJ��Қ������3�8љ��nl���*K��H��z�<c+���\�V�/�r;V�w0�>�1x���f{Rl��oh��ֶ�^(�p�Dƺt��*��y��#]��g�9�n���u�_8�I]�f�I[p�Cn�9��\a�t�[C1��q[m򫾉�W���.�+"�@���[�%�I:z�N���t&���E�}f�s���~oi-��G�V��%�B�mw������Ú$�_Jڇ8�֐���z����+�=<P�j����C-^r/u�Q�|V�j!w�j����U��33
So6wo$�{;wj^ջJ^�'պgm���w�����V��i�#6�WvN��Gcֲ��J�R�ev�W���
���z�G:X�i;���w$�ѧ�u؇E���e~�/l>�Ss�<�P����<��Z�͑�*'��k�Cۯg���^�qs��Ig��_D�ʕ�(��b���͍CJ�PǍ�n�n��֗��e�Z\�����V�k�6�B<��G��͘���V^�q��(��IV����m���Ϭ���>2��3��e��Sy�!�ύvv�k�-���S^�j�O-�o���i��Vr�����n�g�a]�D�kZ�<�N*u%Tur�R�\4ۇ��C�9_'M�@��3D"b�L���V�\�Lo�:�u§�_9}�[���u<g#e �U�L��O�5�=��.4�O��L�"<�3TM��_��^��P��=H��.�w�Z��}+v���n^�) ��$=T���7�yݱ�&R�o�9y��8e��f����pv���&��%�oR����#�Q}86������L��" �k���X%�t9��}�Rb&��3�n���US�ʧ	�מ2��K3>�3�V9<�|�38{;N��"�!u|4}{W��GQ0�n��s\�Y��R}�f��a[9	ۚE���ꁷ?�k��5P�+ƭ��\�;��Lˋ�I��2�]���T_�Ԏ�+h;����&�J3�'�wL��.�+�fԝ��Tjӆjq����\a�t�I�b��k�=�3���#�~�]%�.���of���o�j-�;m�GV�t�3hf���ֵr���qo� f*����e�:�Ծ*^ZN5�Ȭ��3g��w��6F8���޿NZ�̣�"nr����jU�y����3_���y/8�8[���=޼��ݞqc��A��޴Ե����Vpu�N�w�h�kWW1p��\�ϥ���͆������E\K�6m��T�Q߁݉�rbӴ�_��:A�D��Z|�_>�����vt�Uf�Ӻ�N?�e�dFmi:�$���s�r�<�VSGo =�j���[
sd�F�_BOij�������	��(^W�8c����]�$<�3X��	�f�V����Y]�u�`],�7pv�2�R�C�j�2S�Џ���#����{>�1�����r2��T3��}�KOn����_�[��Яzk&����s�N+��|�k��~\�K~��\+U5Sۇ����������{.^�;��眀�^��sF�]T�;�(���iu�]'K|k�/�1n֢k�/*�����sU�8^����:��XS�oI�	h���Y��sL�3�;�������'���\�׹�}��9���|�S�﷞��9���AW��S���}���G�A���4�2�6-��B4��,�q�d���<���>ƶ{�����f5&流!��.f����.5�B9��;�@���f:kz�Wr����P�ܜ�o&��mDw<i�=i0i��q�� j�<UCo.K��E��ht�[Qۨ����%c��[_wU���`��2 r��ڹ�|��8��P6�Nu���:E��ŋ�].�[��}����h���x��"�㕭a*f�`���w	*L�E����n�{;��a��[���m���0vjz�)��%�j�_t��a콭%��ɒ,����D��l�8oS��N��2��2Gέi�y<�OB�"�ܲ�\�
Fq�0T�W�U��^�N(W^��^m����\�Ύ�=�z��&�5ע������2��q�%@�'RKg��g=���Z��\�lM�����Yd��k��Eb�/*%��(�-�*��T��̾��c�%nMj(�@��VRF6�3�����_^wdb�ζ:A���A//igF.wl˺f�5tdY�����r��ވ���}�4��;��Qkl��b:�R����6[ڷ��&��.�<�c��ד:�˼�ڏ!&8��[��0�4�i����P�@��G8c*
1�W��3���Qo^�����ˢyH�w':�h����T�N�yr���vl<��B]>�{H�Xr���;���k8g�eg �2�%��>����fE��q�e+�63��X�z��="���Rw�Ǵ!�B#Q��o&.���}���сM�syEb%+&0�������pt�����ɯ����*��@kΖ�3l7�vdu*�K�Լ����E��oZբ������r�>I�!��Z�oQ�T�	V:	�՗}��:cI-�Į�Gr���^�j����ҫYz%)��!�㱋��$���|G�������4F�;7xT����D�{$��m/�L�t;��`�;���:� �3�K�3�s���A�ACZ��^n�q�]��669F�o%d.��ßh��1�%��Vv�V�ؕ�P�\��Ӡ㼲K2���y��@�{F�t�\�VѪ�ɹ/	�E��ݎ4��e�AP-���-��2�}�jF0Vvk.��ڂ��f�M�-�}�m���f�!���\%언uf��4��=Yo�V�i��J\2CQ�<��֡Z�9�ɋ���V��Zv����ƈF�p
q�f���`�m��eiz),	Ew�u�X��1�aĞE&���gQ*RGv���k�,5�nf�\��l������]���wH��$@�Y8n���{2�E=�d���d�%�Rء��q�]���wKt�[%Z:�ue]%Yyӯ[9����9CB�f�EVu�K�r�[����$üd��	6������6-V˻��6ޘ_ �Y2�n�՝2��ϖF�r����ɷ�I3w�j�PQ��e_v3K6�4hN9"�3"�&c���c�'%6�����.�v[h�4;K�yU�����+������F��klܭ�7vʶ���u��j�)���͙aV���U�I�v�l��wr)
Y�u���@��?�N�����L:��9y|�4_H����|ʜ�7C�ow1���S:MWbx���ۋn��B��P���q���qt7�r^:�@u��@Ȧj�k-�r�#�s��0(|(U Q ���V�"���Yh�E���:t9r�D\8ED&jjVHdl�
֚I���Er�M0���UI,�ȵ�DP��"�T�.R�'N�(��)@r�(�9�̣$�254�((�eUZʀ��鄗"I*�j4�.I�g��U�h��b	Ҋԃ�ITQVaE��E*����feZȊ�D��U��Ҵ0Ufeɑr�*f�Z[M
$�P����ijV�+�3"2�UPT\&QjDTQDT&QAgK�!Tʹ}�p�r(J�"�H8T��xg�r�+�+S�.ZEȪ�����0�%S+��s$˗�EfUr"��iE�9��"e!�9�-iTTQ]  ��@2A{7���.��^��T�ߥ��HK;��4�����R�Y�S��U�p��w%�&�5�Tzb�-[���I�������َ���Ŀ����n5�9g���w�����P_L�_M�����3�I��K]�J�QX��]��OZϹ��ƽ�w��e|6����~�'�zq:��N��U���4:U��Q�͌�����q�z�ƶzō��t��]Y�]�֮</�˟�n�\�}.T@�CwkM}M5K�ޘ4TvA�%>�^�\��v��<l���K��Tr����l=ު���]�a������D�W5��yU��WFQ�p���e�ͨ�^�m���[e���ֿ�	e�i��+o�XS�
(w	.�TyĢ����mg=K��=��-嵭vC���'M�}��TU�V��9�Lu�пf�rMr��<�/;�_�B�c{��gjR���' #�x�6�߽��q�o�W�L`�n�TL,�V�ky��D��3��4�.FP}x�u�w��'6��`lv�o�������iC��\6[|�]�$�eef�}�gA"��}�����3�-�X|a�WF���c����������h4�A��OI��7�*wEM���_`���:��s���؟磌ꪵ&��S�����R![��Q�騕������ĵ���6o���l�Ǧ�y���^p��܉��b�[=P
�x"������j,o��Giղv��Y��j[�D��x��k��ȟ�����Nˡ�l��z*ɚ��S�߁w�^�mw)���j��7F�8e�9�Z���:`Zځ�����*��b�,�k�y�'���Q{V�!){q��5n���v9�N^��q8�0sr��Z��U��rso��X2��:��vT��ֹ��Ǜ8�R�3Z��rT��fP��M�c��;>�*yŕkE�Y�E��o4�R������T�s�����ҝt�B��}�7��!��c�JI\�͸oV5��V;� ���uTI}Q*:��i�x��X����t�,-���o��g.��"��)��Oz`Ӊ#quy�l�77ke�o+���>�M�ZV�ci[���m:��/��4��r���Z��`�R��j⥜����w7��B֨�*w���W�9�b�{��]�(��Pbqh�Lw`)����OT#�
FC��ntn�%`;�^�` f8�Km�ٷYS������� ּz�C��΂���	h';(� ��Q�O��b�P�"VK<r��v�A�����<��w�"UwJ�9�qI�{��7��`��`4��Wr��_9|���5�{Ù1�{Y�YO�szߓ�|7���:�ES튍x�;�:�w�=M��_�=���y׽��c��=�z�\g6S����.�	��Q+^\qj^�6v����z�W)4%�.v��ض3�0���E��+��s��eҾ��ž�7�kl����I*|����$�w�.5�q�	���R;@��8��k�\V=���6u�|g�o֧^V��~�ɪ5���6�Z��q�dOaڸ�9{�9�N�.t�L�p*�e�}+0�y�f���[�����r�L��fݙю��SWiO=K���n�?}P3D���V��9��r���{N.�zr���]�u�)s�5��q�Wvn5�um�o6ކ�N����K�Πs�Jшr���O�;�x�
&耀�x�T䀊�4yO6���>��n��B�/����}�	[Ak-A���5pv�꿛�,W^�8�,���Ǚ�`�BȜq��̾f��ﮯ=QU��.*����C}]큽:����B��y��O�ޫ�z���N<��\�wn��;kǥ���n���[���c�ʢnrUK�x6(j�f���K�ʉ��}��<����E���{Սl��Xnǒ��c���h����N��\���:�jA-��)��%�낳�Yڕ��:�0ʯ-�s��d��<�1��s"����5o��i��jJx�.{�򓗎����DG2̄y��M�y�E<��1�+���]�	�.n/dm��𜽩�۲��5[�����t�1�r����;MI�+�9<�%�9��ڗdC�_<g)�%����p9��gb���!׳4�ǻ����Z��J��z����:�5�!O����FH����֡K�OW�.m,a.[�ji\C/��q��F��4�7��hf3"����IW}�y2��� ���Z㥫�z��ZIut�U�!L}�+*����U�����tt�/%�;��2���_oc�AG�dQo�2Á�M�w��Tro�
R���[�1W�Q�gb��i���շ)k꘍��s�}U�GV�r����hYz�{�[��C69s5�o��eƻ���VR���'sy�r[#l8�eT��\��5�MDv����5F�&
I=�Er�qƺ�����q�r���&赸��̨��j/�uZ0>�P�w�՘��ц���B5��ng\Y�c����.������9z�W<3�-�k�ێ����[��z\/~�>��z�պȚ�bOY�.�
��]�N_z�k;*^�'�s��y�����d�<�6����ڽ�7���T�_Q=��A�͌�}��Oi�;����GN���,�����u���z�;Ωr�uz:����ԣ�Zy�4�&���⥾rZ���6�t���َ�2ϙ�⪇Ӈ��N�i(T�Ȕ�cy�[4'm�>K�%���y�b	YC�eYo.���C��{�ؤ��W(������em����Z��$��:39�ܩ����}%��<4MU������3�5�2m{6�qk��6u�l�%�{c;9���n�x��Bo�q�R�`Q7���lZ[����U)�mܡIV-*�YT$+I8�ﾈ+n�̖���Ѻ�m�k.���{ecqA,��?�Q���Ԏ�����=�x��͝��ET���Jyqk]��g<�z�7p,9_oM�wV&aA�BzV��yp��GbW_-}<��\#��!��O�2�)�tV���u)R\������Dt7��-wqWR�_BM+����� �;Q�֋�_�����@�W�޻ʄ;v?:Ch�;ˋ�i쨘YU#��U��Է�=x�{�-Z�l��xq�>N��V�T��u��K��[�Yz�n�s����Mn���Mƴ.25��!��w%ve����y��kZ�K%�]���rri8E�ہ��+\a�H��g�m*���u[C/�oe>򓳰����[�(��f����j�3���:���;+��W:�y�HȸY�fq��+v�׵��x/䞵��q�<��n�f7nXNv�]���𫠼��"ӝLVH��p�b%��j�Ko�3p�3�S�V3ӕgA._Rgh��F��gWV^xo`f�Tq��\FN��U4�.т�,�抜�\λ�#/�g7�a1�T;���	�����gb���6�r��UW�ϗW{����*/��⎽��־:�5-o������S��F[������귵�i�S�y�{z�Ѻ&P�|v}r��t��*�̱2�f_md��k.��\����}�m�ƶz���\W_Gm�u�B�t���.y��+��Z�m���~~{Fs�LU�fy��oWS=��&f��ĵ�҈�q3��+T�kyoCy=i����b�3
��6��x�$	f��mIu�W)E;փ[oC^�v��P��Ң���^r�>���ʃ�.��]j�K/����Z�MUvΛ#��/6�-Q�v����{>�fKʄK'f�R!S��Ǒ6қ^ƌ�J�ӯ��r�9h^�!�6�Ӫr�Y�P�`�騕�.70�u.�y�>����hƟ4���8¸g!:s��3G���+g�sm6��#G�c]�����wNs7;=�3��t]�A+�kgX҆�����P;=-�|��{=N�Z��C�~'���J����fJ{$�����qI�X-c��a���E��m�|Q��6g*����ZnMf<�pl��#O��|��ɓ��q���k�}S��:���$�l8ƅ�N.&:��w�]Yr�v���Gs#��s�.'�M^-���Tm8g�mƴ�\�e�e^�|^��S�9b�����|;Y��W;�yE��d��}=^;Kݍd��E¼��G_kF�y�T�a��bU�`����`����s�Ύm��3}��.��ך�r8kr�X�͈��������w�}ј�=�}tb��lf�3����f�ݥ��s�v��n��^�Dc���nQ懷�����%�0ۜ����7	?�8��\+�ϛ��_f�{��z+{Y����w4,����󨞥�U��[_D���\.����$*�{��W�����������Qz��#�i��ǺA�R_TJ�T�{O������3MM+�����\�7���j�a�-d�!�)TD���Z�Z�8jĒ�<=�S�v��?:R�^곘:�\i�x7g�ǀD�,Vy �]v��2���f��͚߇3��HR�t��t�c���9l�e���pީ�W�0����l��Ӓ��xw���nb�W%����SZ���ĉ�L/uv�>�����O7�\خ^�;i�-�����uS�A�uC�=�{��.;�AE�^N�ťOs"����=��=k�އ��:���aO}�?f %�夰��=�W�_'���f��:���r�b��C}���;N��|�S�.j����U�K�{�j�Φ�\����y|Z��6�i[/��q�m�T9�5����]J�U���˒���H�,���[�_n�P��\�|����V=�/-J�x��KD�=��셠c��-�W=׍E����=0�e+�6ˉ�Z�k��Y}`��Q��fr�}XB�"�}�z��Lƻ<��l�Sm7V�]���v8��[x�3Qm�چ�s���xj����^�n����o}��c��4��\���Z�J^�q�}�Y���'y9z�eD�i�!Իv6�6f����Ĳ��J�^��Q5���/�OZϪy��ly�œa�t;k��Lcs9u=B,�����%L�=��i�fލbGzz�e��n�}H,)�������4�*�D��u��YO٪K�����u��lk�JT�!�L�dQ�p��B��y�+�z�N�"X�ֱ�nbHoV)�eX[�Z϶����u���.��k�5���ʈ��W�Ob�G�62^>����%�Ra��,fb�o��-{.hu�wx��*P��#�ZcsW7��œ��׾��mO)�ފ��0�AS+�>fS[e���N9u�`��n���J�h6�v6ި��YY���*���*ʢOu����R��[��j�q�MC���j�����+���?-�����(-[o�>�["��G���n�"9R�Ʊ�P�gW�8�r�@��d@��,�kT�?L���?ϓ׼WT-},��Gn7�)�;�Ry��A�/�;���'~D;��wT*!�/n��yQ0�&����5D��cs���f��ٙ��[m�"� h	�ܭ̸ҝB�۸�z����In�&p�]��3�;�r&�3�
�sV��}��+@1z���[3��^�+j潵��'��\2q������wO1<�Z�6-�,҂��\"����G��LT���z�Ww܄�S��q��6�`�Z��2�%ڕ�X֑��LF+�S������܇iG<���z,cB^n�V5�FVn�Ә.�����O8�R�j�q�!-l:$kW"5zTd�ږ�#�/�����N�]�v1�4����'V���+��n��ZR Ӈ�y-[堝�*7�H�lc�'W ���v1�#����{�\�[��R�o�3o���6p6�9�����$̵|4)/��J���IOqޒ㶬D4��'2M��
u���ɷ>�K�+�vf5��
܈-Kz�Mq[
=�(��}X��؄�xɮ�(�S/��y&S
��Bi�2:���7��TC��7щݬ-Ja�n5��ɒ]�����yܳ=���A�r��)$ĹWqn���=<�!�q��-1h��IJ(\�2��tR�Pʔ�����//�z�:5�}��r�^�M�
d�&{�r��W-�v2�(�j�N@B��X��⻐�Ɨ�>T�8b��;�Fe�Y�cjp����z�e�+�Ar[�(�4Z��Q� 9ִ9�;%d�XU ˲��9u�t��ՙ75c�Ccv���
�Ntt�+w3���w]ms�0�*ޱjm2Y�N�IM�%5kI󕧶L[AL���G`괙���v��z���Po��h�-̑1�Ƚ3\�������sP:ʃ��ow�D����@ٴ�09��W �������%�rp5z��nk��P ]�34�#Ьe��lJ���\æȓW�S�7��x�:4�g^��rG���e�I�pY��gvR3�jx�\j�;����;�}cf�ut-
9�R�,Io��s�B�E<��+d<5	휂wB�:�扬F�<�������q�<b��Ϸn��IaX�7[>�j`�s��3��O1`��&*�9���լ��뫬�w���Ԏq�3��i� �8��� �J'v�,:�f�q"J���i��pe:��lj[�Y�����/�j %lѲ�^*�_#x�vE�B�R�]ϑ���mnEC��}-�ҭ�J�3��.���1Cp՚��pd�V.��P �NB����鍝V�Σ|�� g��d��
�N�j˦�k4Bt�ܸ:�0l�-[E��(���++T;O����Q�1�wi�v �Yz %�bGu�B�ɾ�+u��-�����{\5�=�"ԙ�ҼJ�.�W4=��']q�j���0���80ML!�{q�ŧF���c���M���.��!K���M�"�3M�;ڵJc1�}�R�3�.�mC��*�Zcj�w���08��\Y�zx��!}vY�l�*��)k--�sF�k�k�j���i��2��Mu	�6��ᡐY˔d�M�Bح�A�&��rur���TE�]�$�ךES8�s�ߏ}�Bzf�wK�*+0���*���.iؙ�V�5�*)�\Ďr��B��d�U�.��)ȼ���D��"��EA����	8QIYJ%ʚ��&C�DUW<�G��Pr��T	��B�'4�Y�Q�9�ʳ���9�F�EQ��Ԑ��p��jG"(��f����"��TW�QUQQ�J�B�(�1�u��UT]!!3�#<,��J�wAС ��#���\��B7v��)�'t��7!+�'/1�9��(S�Q:��)�+����]�9��f���Ν(����&P9ܹTEQBH�r#����`%K�d3dRl���y�jETH�S���.UNe�h]��9�A9��YXu�/<(�Z�b�e�0���db�V�3�����#��X���*�$�N�DvDD��8�r�ԓ�K��wNhP����T��G���ۙ�3_Г�r�z����&dy���f��'TDpt���oVZ���d�p�O���U�}7.l�����r
���P<����&&�]��:��~�61n@wL&�&��Vd
v��t����Sɫ�ڎ�q��Nm�͎s���c�uҿ{3�"�˧Gy�gvTp��6w��6���\%/o�N��L�y3;���["���f����6�O��Fbߦ�T�ڟ}{\�
���'�N��.��*e�a�=H��7Cw���2����TM�c�b����Wc-[�����k弍u�1��ٯ}�O8���Ig�6�yK�������w�kr�:I���3=��:q}�R%��_f���1����U��z�dWg@w�;�޶璭���'Q%���B��\6�\K��gR�*�@ֲ�[�s}�z��sSy\���U��_%JWo-�o.���i�W�.��Ռ���.ۊicԩ	kf�Ȅ�$���5�)O/�h5�C�a��x��j�s��l�M舸��3�Q�:Ky�	��v�U]��s���MwCN�~Ϧ����'�;F6�m�L�˜qvU�Km_Y�mt�uv�S��*uӜ7piM�[�]�n7&+�3��ena���V��H]�þI���5�җjK�U���G#OW<�0t��k�=uS���O�Z��֩�����u1��o79��:{�|��r��3�eJtw��%��︮���M�4��%�j�J�l��Xm�n��}�=!u>��µ=���v#�]����&s�.eW�	.i��6q�l�Jv�x-��f�mX'�9
�އ��Ʊeh����Y5��A����$ö\k�r'�������t^JN�W9�S�q�ʂ�=�����ŵ�sƚ�֜3Pۍs'�I ť;7ZԴ���Y��L[_�R�*"V{&tז���g�^9��o��yͩ��v�^8v����Ն�o�T/��39��5�Ks}+��}�D=k�DE��W���}���Zn5�9�~~�6׆et��Us�]\��ڊ���a_n�v4���5�&�k;���_�<}���ƽ�us�`U�s1m���Y4�h��j���$(ky,֨�y�:������f��~�0�v
�Mc�����"C��K�W\�r�m�8Y����[2b�u#.�:\��d��	�'#���c����n`/%k��9}UFh��*����;��T}�}v7���)^��;�ZZj�%�m��_c[=6s48�}�QHgc~�FX����r�}*T���-��"�j���ntL^�W��J/�\���e:�47`򯤾���l�}��oCy���i���\��~�W{�j=�>�6��u
̣C�g�d#�)�/[�
1\<5u\;<���mMk��-zt<��|,)_oIP`w	���j�B���/o2��]P6�Įf��ˈKZ��:�3�e-}��n�a��K��UB�V�4��1�[�寺ܴ��׹�h��3���"-��}D��NTS�3���X~V�{�V�����4��_l��oc��9�^���y�`YhC�Ct�����\]x���3ys5����5
�K;T嗷ٽϪ�;�iȖ�L�� ��rV��rok����r�&�췫��X���VYn̪ѭ��c7�18D��w��Υ��	sN�ݽV�m����$�".&5T��-[��v����^�geɷ��ǻ�oKI�׷�-}������y9�g�9s�1��nT���ᄳ�4�Cۃ���!v,�8�>�{k��Q3e���i7���D�!�k ���Kd�]<��$�iRkf�������e^�ɺیN���P��=�k"�T���\\��f�iv�]��ZQy��j�E�F'�����;���|;��*ڛ�<�_f$����.����"{Wj�������I�Y�z�^���V�H73��\[з����=��we����M�T�:�b���p�ϛ��}�V��� j����/4���ok�ƵK�v&?�Zc^Q��J�T�ԩ��fD�Nw���!��w�rM���mz)��R|�Q��T����;+��ۭ�m��y��+��¡ho.o�%��Vu.«��6~*|����c^st���mb]�/(��n�M-on�އ���[|,)�hYx⧉3�٫e�A\�m�	����J؅Kf���k]��s�6���V_.�ȴj��l2����~v:��&Z5d��
�Ssٰ3�}(�h��y��1K�f,t.B��k����ź��v�&@�r�(`�U��Ӭ�\�s]��L�W_ rҙ{z�+��[����#w��YV-c1�栧	��(�Y�Gk�+��oSVd��:F����ߋ�=꺠���1�O����q��}���sk�`n�\��4�z�b��Cy��BD2�^�f8��<ٿf�G;�N,}�˖��=��H��ob�ۚD)�����>���>Ҟ�U�c;�[�Ws�|�З��i7��l>G"S�*�� ��ak��P{W;Og����K���	-��4�N�I����R��j�B�dRױfr��̽��ĭd�����VM�͎�|����	�o��S#je�랚�u����{�a�gWҳǗ�:��\BR��8f��;S���'����\gy�+��ld��ј�����Qڝ^�;��������V��R^������y]�YS�{�����̋|6�N�����zc�2p̮)U�J��8=-@n��y�w�n��Y�7:�yCU雇�w�f����ת=���fsv5'u�<���]zV_V*gcJ?)��H:����?+�ۆ⮭~�����s�Tv=#690Gq4֡')krV-���T��
1"�Z':9MM+tUa��TV���E�:�n3\\4]^���ז���jka����oL�~u+�]M��ê�<�_f�7�������pU՚72�21�d��v�Y��N�OB��d��)
���m�/��L��V����,����'dD�Y��wj$�T��j�+�\=����&��ɲ��vw<�]���.Rr�([�Z�+���JDw=V�iJyCA��U��}Ww�hvɝ���z�3��M�
~_o(������\*}&!��lg�p��U�D�M�9�ƥҥj����3��妡��h`q�yOG+]�s0�n�sj�gs�rҶsZc,l6��fz��|Y��%�:�o�W�."m,a���6��!���8�����^C⑍X���W!X�5�^��+��c���_d�jt�P�Q������W:�{�Wwvki%"6�*��
�̹O&��sƚ�I�'��f�;Nb�	�*�s~9� ���yoi�-݊t�j���ȳ��̥�Յ�@t����^C��*+����V3�K�fE�5�9a�yj�a�)=�e7os�`��G"��M1n��p��[��M�d�(��*�_�����:�>�V���@��;�q�y��ԍ�W��|6�d�Z��K���3��yo��r��k�a���mjk���靸ok�Y��c��o�f*��xV��h�u�xd�Or���2�]�$�]�z����sz�3(��1v-"�$�'�v����6��n����#�8���!�޿��Tc���X3o9�u��=�O�\�	uM�T�(�\4���}-5q/�m���.��C�޷4�.Z��|�(��U�è�"\�J����}������UY,�a���SBy$N�I k5�\�ҕV �.�s>��\�2+�Q��4ObB����^���u.����K�Z}eg+�aJ�6`�!�!,�K嗷��q��\��M+K�}��5�C���E���V	�O��(�l{_��1�D�kY[9���\�Ɯ�ı�_>�񜯞d�4K'ֽ*�]FX혴��d|n���Z�0��U��M�Z��5t"�P� ��凼�����*�n"0�'��O��c.��NW�Pm���X`��ω=��T�+iM��V���*e�T�̰!Gf3�Luǖ#W��Xo9#V⭫�=A�_��-+g5�C}��9���z2j g��R�״��>J�k߱��8�od�w�qIoԚL>|�1T�\�d�5Ϲh9���\2����	Z�R��Jz89|��]�s�;2�oY�����ޥ��.�F&�D�v�B�z��ҷ��[�3U-ձ6�c3=��0{'�����4��q��Fr�\a�t����v�{3�Y�U�Ē/�.Y����ϡ��t����o����ہ���k�5Z�E���QGT*ͥ�m�cֲ���J�/�׉T^դ�ΌN5��垸ǵQ	�NV�܉��,���;�}G9U	6�>�]��X��R�\$���u�i��Z�R���{{M���~�K��P��MJ�LuQ=���͋���/��\�o7���o�M��/��1�z���T��]^�g�I��OV}�<��ZN�c>cZ�{V�c��|F�fD�&b��M;%3��yY�@�d��Ա�1�R2.��j,b� Lr�d��p��M�
1�h����X��"�J�*�{V9��&��s��e�����㷵��&�:@k�<�*�P���itq$���Q������ߪ��zt}�����Y�����O*�����2��w�$��7��6���Yˬ��3J���gd���h>U��NF߮׽�UJ��|�z�ͧ�V7p,(��yjD�"�A�M���#��3D�o�����Kf�Jymk]��uD<�k]W3H*���+V�Rs��+�r_�|���cϢ�_�ڨ{�un�����oQ$ߟw1��
�ܸo��W��{v��&8�l(?V��7'�cn9Ʋ�9ܘ�����۔ΐ��h	���n�Ί{�;}�]�砬��C�<�k��p�0�Ȕ튅l���*n�[������'s�}nu��^M��I����Mƻ�r'\\OR;�m���k�����7��'�5Fl���+�;.;���'F��N�����<�ѡ;���^�:��~����Ps��)$���ʡ�ҥzͰt�E�V�؞�dd�,{N���%�c���7�E�*^Ji�O�jnY�����Gfj�n'r57�.�o�R��fA�^�����´��]���:����`��A���w�nu�'��Eܤq���BXֳ����eJǷ�j��\%/o�N�ʡ0j�^�Y�M�:󶩻�ˍc$[��F��J����j�������佩w����4$���C���'y9�.�
���T���:P�2��Y7��M��f�ݮ�.yãޞ���3]o�n�yŏ����{M-}�C��G7�Kq��%l��ҭ�6�D��ľ�oF5��V;�o;�8vT�Y��^�]� �yTK��2_\aH-�Gͷ���|���
�U"y�m��r��������U6d���zˈz�R�]M��mڗ���F^s��
�"�=�R��)��^���Vҥ���V��\�!�P�W�׽�D���ٟI��o��r�E/'�4�I��ܿ�V�gn63�3��MF#���dḥ "Vk�Y	jy0�s.B�(��ul�x�p��YJ��޾
�U���I�廚��tx�j�_N��\��]r1��/d�I���$񇲷8�.�U�J��()�@�`�d�f{�H�p��Cx�.^�nOo���R��^��4*9�Yq؂�lf��/XC��Br�\?N�f�rLN���st��+
zɮ�jeE�\�'������%�6��1��U���[�G+��T��P���fEdG��GfG.��Wt��������-�]�������5�kO�����j�p�[v�N�[ޞ�`�,�/�`r�j��y��e�em��0�{�-8�%����'����Aֹ���ɩ��v�l���ݡ��+����8Z�7��}����YQ��s5�|��(�V�KT���(V�hM��,�����9��T����F*ӡ�?�+��u
���ccկX��Vj�{ukxI�T&C��g?���Tu�]������v��P�W׌���Pggg\���\�"�ɛ��ͤ�͚�LJ&|�xy��1XϲVf�m'�[}}��V�F���f,��V�8��+�!ElS�.!4:�z���)�3�X���R�sm-����8lVI�r
Ҝt�*�8�m沭,ۥ]B+z�T�Ik��"xuۂ�As;3ʤD��s[�)���ki��c#%jʐWj�Q
Ty�X�	t�v�ֻ�>s��A*l�z��ҮW����Q>ڙ�^�\6iC�ױ�ں���<��j=��kso/��F��9|%�r�r�)���[��0��Qv�;\~v�Rd�IҾ���x���p]ڲ�o�
r���G�r�p��λ��b5��0�ҮZ�_-�T���B��6� 	@a��塖n��A��闥�V���}.�P4�l4��V+C�s���Ƨט�xT4V/�bJ0�i]�r��/�Y/r���:�1)�ڽ�B�������N��5zv�#�	i��!�*r�lj��*�n�0'l4��>G9#���ܜ�'�d\�R��LuC�۝�Y5�˷���鳝�/9��S���]ن.��"e#�z�
�q�d��7�F*�*q�-Ak�Ql��	5q�yWk
��:@r[0� ��J��T݋Y��\0y-Z8��G����Ӧ�FH;����y������r;4+eҐwK�t��/��s)�徊ʘ�и���[g�*�XO%�ˡ'Zܘ�7���e�-�
�'��k�נ�yn[i�H�|\t�����;�I��̎�b�Z�bH��o�!��7J�n٧�T�Q�'I���^q'����0��g�L{\�I�w�Vu�q�4����L�r�wJ�@t�*�֨�u�U�7�a =��c�.��g���2�4�t�I+ ں���Y�\�˥ء��mj˽LE�IWE�f<8'&ͮx�Ԥ҅����+K�p�}jش[��ʽQ�#u�׭��uw�mf���r��ҭJ���3ZfNxp�YQZ�ҧ[XAʪ���rws�r"*�D*���C����uY��s���"'�r&\��E�GGqdNK�P�	PUUr�\��Q�ʊ/]�¨!ZAr9ȼ�T貂�·.����Az��TwD#C�ҁ�r��UҨ��[9^���P�*��Q�z��2L9+��K��Tr���%�:���9����!��\�[�r��T.We�R:�QR�Q�c�p���W*�R'%�eU��m&\��V�\��GI��E��s�AUEQ܄���DQA%K+����ĮEG�t��s���W*f�"�Ԫ%AE���q�q�Ȋu�҉�	rr�E��&Q�L0�5�&:	&!͕��r��	3$�V�^�+U��oeJ�C��������;���9Juף'�"�s��Y��2�˻�fsf���o�]�Ȱ}<�P�֜擝g9�B�W�oe�M�^��cl�C�sH�=!p�5�)�։�׹��j���Y&�[�|���%�\2�;gV�Bt�|f`�w�Z�m�kf�[�m2�*�/H�_�ڧ%vMGju��B}E$�Pˍq���ze������7^�]Щ^��t��zr���|{$k��Nv�s�i�-�Z�R�k��F�u���,	�
�mO��(��M�r��r�އ�moܢv[i,6�>O������[��x�[�u���n���}�3D���7��Nl�OsSU��+��m��/k�Eޤ�]�z��ܧ�s���O���ov�ёyo'�E봲��E�y�j��|�⧜��7[ׯz��N�� �����������E�=r5������ꁊ&;ϛ���5��8u�o4}u�3;��s�X���j���H�>��^Q�.�����ą|������K\����:B���'oi��	�L�1M٭JZ{c+ȍ�xI\�j�n��S}����*{ݳ�+���B���\i�k��Y�C��Q>��<�*��O���k�/:��y���j]D��Y܏QAub���D�9W�����ܞ�O��Z+�����ⲱ �����Y�˔�}ɾ֕1ί�_݉9�4�&+Ό7��F8���4K��WFQs>�&�f�&��!R۷}o9_>��qõSOSۇ�����C�[p^7b_o�&�E�VN�ⲅ��g}��6[��_bX֨|3�3��J()��Y�ʻ�.m�X�T�?L����P븎+�寺ܴ��y��h�x΃MT�m���}���y썙q�+��݊F���/v�&D��=&׏�kC�:Du����Y���fpq�lS�sP�<��j%nMn�_.Cd2�[b��s{�	�/�����#��1����@�rJw3Ap^�{r�q��ϝ���Њ�q�:�Tj�`�n5�#9Z��; Zڀ��\#��C���M+�q<��ם��V�9:یN���m|��F��U�4fEy�|!���8`�<��f���뮖�"������̴1=�G�3;L؝����y��G�Q����5��"B��nlv�8�q�.��gi�[b ����8����ޭ���m�ѹ��՗�Z��5�:{}x0b�)��JM�E�l]���#y�v�9�奪�R��a�V^J��y΢/jե/n18�x垼{Wy6�q��ic���o"5Jp�̯���Y6����+�Ec��K�p�ֆ��}��n+��֐���7=O8�0ܣ�|=�uI�k�6�N�O�BE��u{˔k�Ç��\��z'�O��z+{Y��Q�A3��\�=�Ю�v�sgwy\�[�b�k��M5q�6�U�l���t�:�Fd�x媖���Z�rU����U��j�K����>>ӟ{���^wY֣l�2�q ���b�Y~���f������zXߪ���D<ub�z�8yK��Q����ǻ��,��z)�O��^��ԭx���;�<�)+��9.�};y�:~�{>g��p�8=;�����U��u�Wx�..rF�:��7��8�]���J�T��E>򸫈�yb�j�@˦�kg3}�۝��7�E��!��{}R:�wlS$�@ �Q#�`�\����F�].���pK���	�G�qMX���2g�YsLo�t&����]*�7�9��8�O6��t=Ӡ)�6���/p�d&����iÀ�Y�6�s��C�uv���;�z�i`+$�KT8�ʇ�B88!���	�'�'5y�ֳ\U�Q���,A�Jݪ�r�C�^�v�|Nq����h7�z���Y�V�IaI-H�GK�!U���T`}��Z��Ϗ���e3q�B��U�+ޟ"|s�L��3Z�߉�}*l��Z	Ҕ���Q��mW�u�Jp�Y^��s�h\WK�W��o�Dzߕܘm���y��6� _A�%]k���2oT��u}�J�=쓾0��xb�-�^�i��6�䪬1П��\c�L�����Ƈc�w����kR�>���N6��=>%@>q� �R1�T��m.�UΛ>���a��q�",:C�a�#�{��y{ܪ�Ê�LE�������~��:��7GuӸ��#!�8ut�����_]�� nV��^�)=�UKI�z�;�v����_��yg%r�p��/Ct,w.�ۘ)WV_*�^��y>仰�Y(���P�Ty}.ix���[���J��F9���Ϟ�ӷ2��,�y۶}@�o���-+K+�7�T�>JG��,�]�KԼ|�S���*�;��	�s�突E�0-���wvg{��j�gFT>(I-�!��Y]�E������++ԇ��{�k�We���S�]�+�iAݕ�{۝�MN�lR��ۋXl,�K��[e�ػ�BS0�s"1�+���P.΍ܡ�"[�u��T�V����Iّ�+pZ�ٱ��+���C���ju눋����/HU�h�r>V :��Q�Kv܎�q���-��<I���6j�b�R7S��<yb��FG�O�w�d�s�2w޾��R���+��'�(5��,�<ITf	>U��fIAx�yQF��̵��=�~�>�����m���î�R�Yj[zg�x��� SRX��|=-��~�ՙ����]P��v�qW��֑�3�+��N�t9�7LN���r�@����V[q��[=V��+� } �,fx�F�*Ac�[f3ӽ~g�������UW�Ie�FzfjRsu�g���|C�@�F�42+��;�σ����m_������/�c ^�|:;׳[��ݚ����W��̐��������n(��V����N���w"�^'�*��v��n�J�5r궀KEF���.+�'�����TT���!��tf�>6���7-��{�݃+���ի���CJ�Sp�~���qލ����@�|F�kպn(�>��(�8�t5�Ԯ'ʏ�����otͯ
ނyԏt������|�4��Oq~t5h���ԁ�XU��V���MC�S+�r���ΧHHkyr�l
YZ8.�h��&WJ��גӥI���G����L����o3U�M^�@�jqP������V�u*ONJp%^��mul�	�Γ�1�E�i�dG=ٹ��6�5bP���܂`@������͉����O��_���+���Wȗ5�0ߢw������������ӌ�;;���_���]����$��G��&Ш�[�U eƓ&�<8��^��{�ޫ����1��Ҫ�^I.�}�\���V}�;�c�E�����,��,��hW���ϥ2��M� �G{�$�4|�W���R*����xj�C��U#,����dOg����(��]Io��I#~�S���L7��C�dK�B᭩G�<vJ�*��>G~��&z=����<���k���t��}}K>����T{�3�,w����[<	=�L�#�a֜X�;4E��o]k}�=���v���z�U��~�R|_7[�W ud��2�\��A&�U�^�����6�S�==:@<�Xϖ]{�"+ޤ&�=^�47���ǔ�*����US0�R���zM����J׏t=�d?�t�q�)�FXW�h!���<s��}��'�}�� pJ�x�n��V�~���v�*ْ�|���P$W����ڄ�j,#�~t������l�Z�v��LS��6/����>[e�\Y�$��o�r�r-�6�e�55�x�'}+)ۭ��tr�A�v*o��lcRj���xR�s��Vn�-�<�0���t����B���Rޥ���8�5�����\Y.>N�bRu�"{������~��Y슷3�	-Ă�}FBӔ��~&C��V�+|wq�����jM�z�>����ցO�~��P�3�o�<�5��;� ם:���3�'����R+O��T;M]��}�d��@��j�_9󺡎5c�/>����U�����.��V�_����Evׅf�Һ����w�25�+�o�����Foz����������nR��#�'!��ᵡIzpK8NwћHz�λ��7^�������'�ا���b���ZԸϴp�7�u�<|N홏*�;��W��9�v�[ T^�_�s��LDo� h�G�o�ݛy����-��[�y�c+��tUvE�B��*��Qc�d�Y�DgC�yS�=<�5�wk�{�j�ܙ��{�{θ,^�B�κ�˜%��xk�=P���R#|I���3��;���ϻ����|}(;���*�/V�_��ϫ��{#ϱ�3���ԒU}2¼�*���'�coQ;��[�����E)��Ϧ�_O����x}���g��q�֢��,���T�]��5ϏٲU�3+ 9M�ecW�a�ٮ1��sgj����ޢ�]�*�]��ԯ�'g��u\�2)b�F]�9H-�A�9Ns�L}�98�;4(���X�B��V�O��]�����r���o1(�����њ���S �y�6V���RH�f��ᜨV��:�wof���Է�i,�>�,	QBK�7�i�C�V*���ÆDyS��>=~��q~}mޝ�W�qR�n�_.R}��œ���'�X�)(�[S�.�};y�~�}^eς3���Y���ww���_lazR���;���(mD�d�A:����X�CF�y\R���_����Y�z[��g�{Ӵ��zxi+��ު�)�\�@M<fu����>��W����my�#���v����>�Ro޶ω�>�~����h���2K�-M��h�W�k����-��lʶ��{�+�T�:7���>B��W�7�O�>9��>�k@���.O�M,��wJ+7�ʴw���=X*vS4/�r����|n!/Q��w&/�߬ɷ���C5���չ+�=�5y$������v.au�%�嵃b��M^m1���3��w"��zdO���C������ 
��~J{�C�o�d1�/T��GER�^�vo[/:����4"�2�m_��ך���P����f��c�ӑ�uX^�����py�0�����zN�������7��i
ܬ��B����A�䵆�*��c��t��3>�&nlnSU1{1U�V�f��1�v�_��[�CD�fQ�K�Ntb��!�S�N�X�.��:���}>�٭D�Ȭ���̃���qƎ
ܚ'�iY��<ɠ���d�f֙�[r���[�C"}U�%���)p�u^�s��emGÛ2��N�=����Yϯf��󇫽���B�K��~ �ܑ��ȕ����=�劷�}�}�<1�:�5���4ǑE�=�`��7?X����������x��~/"+��{#޾f]���yp�8����jP3�VhY-��>P�b�|��9�4<��.�"�W��^�]��@`�=��n�Z����=[�.ڟ�<I�3Ơʦ/�H�UO�yX��;޽�����n��_<��X����D.~�=���	�2K4�U� yL<���n�P^91�IT�'��<h�$��W�i�iȇ�>s��=��=��m��߇��]|��H`Cs�6:�$z=;G^��u��;�c��yTR��z�9g|W���W�\��][5p�Af�AWB��*�W*u5�<��~�_����|/�F|���H'>��8��_��L��~��'��w�BU�vgѝ@�mo���r�Y�莩#}pG���E9�@�7�Dk�m_��+>9��wĿtR�\֍ɮxr�F�T#z��f$6�Ծ��01���}�/�������?J ����.�����>��0������f�j-�/�f����X@,oXW��Sn��j#�^��;,ȕ�-ޣ��]��;]&5�.��u3R�S}ne:1اF�s�S,�r(�r�}�%��<e�D��z�T��Q��M-�<�i����eݎ��~]��u����I�i�{"<n4躁����C�g�QR��NE�y�����}Sv־��Z+<����zurn3ޠ=7�_�����jE�r�~K 㶥S��un���Tl�}�5u����gY�G�>�q�yp��V�����g��'��{�������(��z����߮��{R�z/�N��>�p�f�f�:���s^��'|s�,O{��}�ߍ���!C�wёW���Y��Q�^���� l�w9GD���]L
����ȗK�%���{�Cz�ޏOu����{�k�O���c��6����s�}�ȱu�Ze�<������"�y{<�q(T�l��Nέ�ͬ��UzQ�WW�����7Ϯ��d��aᨃ=P��(�9�ّ�kѕD�W�z�]�QžIm���yϛ�߯�ǞW�^R�dm$�Q%x��Q�"�M�J���x?r��s]�g����Tǳ�>�a�t�n}����yׂ�{h<	l�$�,Sjk�;d��u�w((H���g䁽5������s�p�r�2�����5���GC��᝷
�Ξ����|F#ۂ}��U�{FmN������j������[:��L�K!Mn�<�u��eg.�md%}���G�^J̀B��J�[�҉�:�օ[-���c�X�g��0�`Z�ݱ�p�� �C+���Ҹc��7yT�U�%;�L�J-��z�3.��5ڸԫС�����[o+I�5w���3cE�|a�T��"��E��3f��uB��r(V��Є�Z+�8���Ŭ��-9n����(�w8^U��M�h�W �um�
�hC{�Úw{7��JIôM���2�K2
�gsfVl��JV�Oz'�C{�����R|�ۮ��I�b�;e��ci��e۫'��dػ�Ij�<3.�&��{��GU^�pW;�2���rcsi����(�t���7�j�:e-H�t�B��6�3A��wİoe�攒�&9HS�)����k$�6��}��8df佾I��G�8���C�X�&Ԇ�,�]�!�����3c��7zn�W��.e
{0(:�G�΅���'>��v���zݭ/�r�W�KvT�Ӛ8�n�c�{F$���-��S�$f�[v�V��ʺ�WZ���<;W3�v�����neN�;.z�)ʵVɭ���j�l�t��Ԋ�����:���� ��h�J���B�lՔ��^�7p=n��:ͭ�����'T4�"ʮ눴(��ڻƻ�+�3C���0�"k�V��٦��*eB%ܵ�oŽ�''"+*�Es��R�� ��bXjT�b�Տ���m������Pf��.BvWU���,���<����h|˜I�����]�E�>�dԆ���s�m�:���𹔰���F���j��u���'�tW$=չd��8���ʌ⧺u4oY�wɢ��Y���$;Bn/��'ɖ��z�����dI�*�H����Xs#]�L���i�}Cx�󨹃����7D�al�q��	��"]�/]�Y��w0�$u�9��Ǚ�힉b{0vf��M�J�ގ�8�B�De�AN&�iJ�+"��4e�Fl�2��'I��w�M��Ǭ$�mӅc��w�f;���u�R�IQ�
L,���ˉH��/��VliH��ɼ�wg%���I�ux��]�; sS�'I���;�I��B�b�Y��Y���{�Mfܒu�Yu9���4���Yl���.���jsWGow*Fp��b��j����.��E�]J���WtZ&fN$��	���5��3XB�i&�WI݅�%��/�`�� ��CyH��Ʈ?*�Ei�VQa�P�������줫�έ�D���y����2��ɔ;z�B���%��z�ޜ��K�1��vG$'�ԟQ`�iG�b�ݧxf���n���L��;Dn�L���"��T�O�*��8Q�H��W[�r� �����9�䤔�t�B�	�Et��E��9�ЫB��ܓ���Y�WQ(-ҵ/D��H�)l�"�'<��!Er�*��T�Aʐ�\֗ ��;��Q��d;���((�KrԵ�.]����O%��I�:�j˝F������G#ԫ���rI�
�+RT)����i�<�{�-.T�Ny�V�eR�{,��Q3<<���PD�Bh�KD�4�ՈN�����U�a���F���a����RT��\�.V�#�TIz�r���iyk;��w,-C�r�
8��u�)�P̈��ʯ
LY+N�Jjf{�����1B�����g��9�B"����E�Z�Ve)���1 I�HU"�kH�~J��@�T(��|����]�u�G}��.�j��a�Chat��1EL���/� �n��\����3d�x�>"����)o�p��)9C�qL~���9�<ub��q�'������=���V���Y�{}�:��yPk˖��1�*�e�#g���W�(d,�~9^�!7�Z2�[G|��W����X��d���
�ʫ��oj[#ڌo�d�i��Pd@o�����9��
�}�A�W���zw�í�yGLMZ���u��3ډĨ=-��ͩ֨lD�b��u�
@���]W���8�.��\A�/�&��I��[܉�x��['��z��V{"�>��FIh�� ��QȢ��Mt��g�(���R�S��{�c|���o�� }��^ w������~���3�n
�O��}vR��>�����m-�p�T�v���J��?;�7�_��~���C5Cn;�6d�)�T�N�9�/U�/sU{�g�9��zt_�����6�J���0�_��&�=>�z�롳~�e����[ט�ܹH�fY�,�W�&�Z��N��s���m!��d7^�~���>�L]�I5,ZGV$�ܣ=�W��ǽ�uKֹ*�d��R1��S�UH˝$���;���z2�4(=x����y5g{
�d�v�<�'�1ѭ%�g��:0�Ǆ�͍:���:�ȃ{�j���o��3=�V�*���Vׄ���s{��*�j�rv,�{/pڬ�3ke�ݮ��tt�zV!-$�Vv� ���h:W�%Ҽ������վ�#+�h�d��\�yg#f����>r���#}O�w�`כ^���	���B=JE�U۟UD�[�]�9��s� {u�"�|�{�v�Q�S�9����/|먬��%��xh�T,W�^��}T;�鰪�Z�J��}v�l���r���������y�q��}�o��֤����m�C�y[@m�W^�^C�e�T�s#�漍��[���Hn�\�����g���� ��Oi��T"rFw�qZ�;ܫ����E�H>�<���H]T�9�x��[�_��!�c}�|w՛����ǁ����[䁿Gw�=Z�<��|k�x���`�}-��Yu�o8P�OסM���K��?n����U^�^�8{��'M��~��Y>:ȁʌÁ0[�(��Y#Pѩ�{SV�
��C�2��ZM,�ﲟg��O���RM���H��ݱV�K�D ��<Cs��Y7)V_fE�������\�Y��f����!Q���9��>��OV��z��Vx��9�XRKSQy���Td��ʌ�x����~�*O#�8ˇ�Tu���oޟ"|r=3�'��h��H�֞���kޣU��������)�m�	W�{ݝ�jc5�����b�F����r�ۃ�z�є���ts�t��z�טە������^��o�G�'{J�G%�[�������+T)�W]טN�L��e�2���
4��x4�'������wjE�ј����g�f5�U��T�4'�a��u>6���\?+�0��+�����}�e�䗔���a�F�)@��T��0�D�1_K[z2��M\f�p��2�܍\*}���U�}��\�ws�}��=p��Zn�T9P���A�b�Hl��Siu�o[D�ײ�M��ޭ��W%WZ�%/����'�tI��uęީ�^�� 8<��ڇqY^F��n=~�;�۰=����%�ǥ���?O�o��W�K�����o���z�
����~��;��AӤ�9�y��O*~F�E򤲽�g�Q�DQ�%;.B�+�{����+}�����o�6�������wF��e�5����zgFA>��86�#�o��V5�
�/Z��3�~*}��m�3N��Fe���j�#/lǡw���"�����g�O��rWf��iv����sũ��o�����s���ފU����a�L���x~9eSJGj��<��,C�X}���ζ�n��ۚ�G����{��uǽl{�D����I[a���P�Y^�V���d�D�����������L����;���z�V�^<������υ]�J�+f�
�;A��-�����9}B(��c��{�̭5��7;5s��b�T�B�n	.����4��N����)�R�ƍ��Cө34xǆ=�|��T�+�׺_wb�K�o��>�=���������=�=�{UH��(	u��j$�7#3�޼�w�j|j��-��<��eX�8��"$7GNbԽ�)w%�|WK��:buC$g���wRsuj���^���@���1�P�Rz�1����;��&��\O{}S��u둝7��{w��}E��0�h�����&-�O�r�����dsj�q���:����c}��\��ډ^�Q�+��\U���M)���b�_W���E����ǮvG���@s$p'|���ۜ�g�|�R'�3�;�̊&xzA����;jWzۊ��x�x|�*p���}ӪW�5!�>�{hdC󫓏��G�~��23c�r)�*�����FB���q��GVfs������S>�Ҹ�U�>o�|s�~�=&��]xO{�t�ɛ��x�����x��g{j������ʷ�/��Ǯ��6�^���6W���j�乯i��o�]㑾�𕟿_i\������8����݁g&���i�G����L�(ӣ�S�t])�:�X����p
u���C�T���!��P��T�ɋ�/�]ъ�g���h�o�0�+���������=u��Jsk8���:[Cd��+��-ub�D04j,dYjD�\�0��0�]���ū5�m#X� ܶ����4��r��kBܱ�,��Mf��k]vH��cɊt��8�pg�I��S_�Z�r�g��'v�3(O�b����t�+L�� �����<�Y�f�k������E:l���Ho�������hY)�;0�z�� 5s�V��s�=��ef������|�����z{b�Ly�W���ж��u$�ߤ��*����o���8����S�]^�>����o�U��z}g�O��{�=�9^u�^��]9�I����{���u�隧?@?��]4�*��}I�x��\>w�9R|_�t��j�}�V��ig;�vh^����q]��_�4}�@�W�x	�)@�۔2]?���	���������Rt���0a':�ȳ~��][��}�Ww�@�(� r� 8���J��e�p�ւ�:beo�glQ={�ugg<7O��:\M�}a�H鞑�S�XH;��e�΋�0���>F��F=q�^�v�wm{��dP�n�~��"}�3��߽��.=Y슸s>���d����&_W��)c*%�'�w>U�{�|},�y��ϓК�I��(?�k���o��~���gȨTq���Z�bh�)%�+oA��w�WZ�'\8�ҏ��M<r�S�'�N��r^�=���>δ�ŋ�E�Z��;���KR?�*������kp�E���펪��w
��gR�u�|� 9Շ.��u�'wڤ�[�nd�na7̎*����L�/nqt���PL<��9�+�
r�z*y��p�}����{!��ɿ�_y'R;�	��j�5"�#���J~�[}7y�R�K�9>>��8���{k�%�Q��"`noDRռ#�O��z'U}��{g(y��Դϸw�:f����P|�rX�Qه�TdF�%Rި��޹�>n����J ��{W��y�����U>�4��o���~ͺӜ|N홏*�a�VW��9�v�[ {<���nQ�/ �勜��U���ҩ^���W��צ���k��+�S��%U!8�(]�6c��}G+�z�F��k}�]�},�x ����^#>�u�q�W��h\o�u�s���2����O=�y�]q��GbĲ�ѓ�<}T���(� /�t�}U���Q�����κ��ƃ
A�G�vew�/��|I�l(%��T�SNBr�ϋ���/d��[=�<�	mʨ�{%K������������ĕ(mT�9v�t>��p�!�ckn4rR.�uX�˿	���;��u^<v�j�8�?@�,�C<ITe�1 �H��l�L��~�k��W�5�n�;
�t]@��`uγIԈԢ��̻AL՝v�z@��~x����ݍ�曒�����mww�Z1�m��^��aw�y03+������lm+�I�]}�U��N�3���sR]��K67�胵���U�=f0ޝ���\�4.���q�p�+g%v������]M���GJ������a�P��2q���$��Y�u��`���7�[�����s��}�����:���&����uǮ�d�;�� x�x�h4���ý=Qs�}�jW�@��^g�5F�!Q�߭����>����QR��ɑ���]��sEMV�r�s9����Xw�����"~�T�\T����2�o��Tu���oޟ"|s�;�}��h��:
�ۛ螪~k�qvr[C�d�����%aV
�OxП��S◤�(~Wrb�~�%��"b�U��yY�smfo.�jZ&2�d+�'��>߄�TK[z2)ϴ�l����5r�΁^ź����NWe��WEM�G��AL� w�^��S|*�k~K 8ې^�~z�[G����z�w/c5-iJ��w�LO���[yh?L�J��3y�������Z�m�܎��0y;��=�u(�]�V�aK��g�|���+�����꽤�7^�w������~��;�t;��:�i� ��Z�Υ����(+�ʭ2;ģ�e�[�Q����/�N��#�ێKը�a��������py�{D^�B��Ў�%�B�s�*�+����#uN�.�m�-�torӱ3���E*�w9�i
��Ͱe�7n���l@�k#n3����YÎ�hNl�Ċ�K�wP�6�g�_4�L��*���p�\����k4�M\�)jn9(~~��������2	��*]�yM����|��x��S�z�&9�d��+�$��{䯑�����8JW�c+�g�S>FY�4<�4�`����N2c���O5b���^C=ʛ*}({�Z�[[R���:�3Ơʦ.�R3'�>ً����r���vq�������k��[9��Q�z����x'$�P�P0�_�ʡ�k��T;��N�ɿ5ض�<}S:9���{n*�t��s�O��}�=�ڦFs�߇��]D9 r�U>��������X��0#Oi^��c��W������q�����+�ꑝ�f�>�͟85!���P�܊���+�����@Q�O��C��qKm�a�lt���W=��s��A�����k`l�xg�S���:��ͪ�4?rD(���@�<Pt�o��P�s�F�$��/�f�/����{U*��ͽN�痗����9@�`o{�D�OΠc�:�OY����2ɭ��ǧ�f��Q���q)�dh�r��p����<g�w���(oH9���)�ڐ�� ۊ�pj�_���
.b�un�.U���G����"�jQ���^S���G�)m�c7�_�Ύ��L�D���.m�q�'������sa�cxi}�9\^�/�A��Vq����hF'u��s
��R��y�;sp4��}�h����B���1�~uro�M��_���f���*A�>%P8���7f�b��\�ǝ�x�,�p�}^���i�ޗ��.7�9����z��{=�_/HɖgV��T��+�nw%�P8|}<��Ю+)�����͕�y֮K����o�]�o��%o�(�58=#޺J)y�z����G�y�#Zr?�'�l��(����{��.��mg�n�G�l�j]&�~p�����Z��1k�U%U '�/ش�y┈�'�Xm0�w���/���<�s�[�+���Z�^���҆i��/���r"������y�W�_�@��}�G^���u��)z�� o����?��ǞW�^RmH���<j$��PB`/O{	\3}�f��e�Q��}2�_q�{D{���r=��:�Y/m�z��Te�>�5o��a�L��j�YS>���O�3�X�|��s�)>/�W�g�{�~Sk�;���c�K���i��I����p4��ި2���@��C"]?��	^�Z2�[G�5<d��B��*��w�t��	�͕x�7RP{c��u(���N����s���y
d����q�^�t��1��17�jz���a'+Q�#GQ�ɽ�Dt�,���@/����.漀��꼔�7%e�U��\鎂oz��r�܅���[k��W�=�n�w�T�>%� ZdL� ��#,+}�Aq��oks�)r决�ή���q7�WH{R:g�D�u�rrl��N_dc�k�z$�׹�ܮ|��FW����~�<}(�8���n=�W�\V��L�Ih��#l(���i�5�Y�<�ȴr��~6���IQ�z�>�� ;��h���m�ze1]{j�B��ze�Y�yV��t��:�E]J��6�_�/mǳ��w'~&J��@w���N^����7�����k�$G�#�0��;(u�8�JӢ��{^f��i^\4�U�k�W��'�}~��I��{�Q����@+6�g��f���d�WkC�����9�w6P��^����@�z(��W���]�a��zt9��ό��}|,[�l�/0��U;�����R#^����\�58�����i�P� =�����8�{�/az�r=��6�n|�Iݸ3�waL�����pz��a�Q��^ -j��^��2%�c��o��d/u�q�u�U%�����rG��Ozw�*�c8�Sp�t�uǐ���KN�D�Q�Y�塹�Զw��J�i�V��<�xN��ӻ�5+�@��Y4�uw;-!l�]�p
��n��]t*���Z8a�wF^I{Y
qNYK&�4Y�ƥ�XmR��9�,fR	�ܶ0�\*_LY�V�;X-�.:����nv�]C�T&c(���O침ɓ$�+�'�[��`�;JN�G�wy�#+��r�������tQ��f�Y}z��-޷Ng�":�j��U�)���r�G��f= ��.,Ø����e���\�E�/P���q�p�
����qh��7F���G�e�T[Tt�[���n�F�0��X���q҃R��7*Xo�*mG��vH�C4զ��X��ݴ㿕Ò��ǚ30�4�X�c���^P5�B{�� rf�����w�]I� �Ɯ���!�s-��X�3�oFӘژ]ٶ�]�����tG��γ�Y�.����Q��D�Z����Z�u���ۺ!�>�{��EQ-Tk*��^=|��g���I����ú�Dc�C_iskr�(��3]�5�9�(�ٵ����n5��mK�ģ�t�p�Sy�r���5�7.�u��U;vs�\�m'.U�x0�6��L�֠�y��j�wY��,rRz��|�,��:U	�Ǽ��c���ۺ�bU���&Y�N���r�L0e��ViZĵ��no. ���S$�:ҹ;R�}�t��k~<F-)T���N�Oe��1�a�S��l�]��rʬ�`�Cu3�mr
��N�]�mvЋ�B��Q"&r�w���k#�4|���Z�<_F�i\�eng��n'�e;�C�\A�PncR�h��}}W��T�EK��8�Ρ51����L��ζ'ce�eWl�&C��#���TQ�qT��n�v�"�Cݔ.A��$�ViKs'%y�Ӓ��$�ǲ�Tv٦�Kb�i<z�XX��}�M��N7ѷ4�;��ޭÿ9�ds)l�I\IH�貂Gv���{B���k�oh����2�ZJQ�a����8�c�Li����Y��:Y�f޽���G�'�.�<mB��
���wcU��fs�1�k��A�w�r��f�C�꺽l�͵w	��($��ř:����g���s�mC|jL�֩^ɨ}�(j��a��bf>//;L�Q���]f0
Cg8�0X�.<c3K�I���bk/��x��nT���C<z�k���@3�R�R�K�|�Г��4��0�W�$e݉Ґ�\�z�a�*��#�QT���l�X���T��[|CtQ��l�j��N�m&9Ν�d8� �6,tsn�T��-�b�+��dp�1��v�y��$�*K+.!�6-qQ}����y�;bڼs>��tt	�:�M��rIE�u �!\�+��c��
ꕃ%���,˥lA۝(�El1gk�wn�W�\�h꾕:�r�=��,���,��sP��]��sR�"�5�+��U��O}"9Nuw#��<�(��YTVeA٘U˩;��u6U
��VIJȳ3*,���u�d�Ub�H]�q4�$���V�Z��Y�<ȼ�J��52���ww!ΐ�98�bDY��#���;�E���%a[U*�T��S�%˙�dJ��k2�̐ꔜ-j*��֕dz��%�U�UUUD�P�QFaAR��Ea	I�{�����{�w$
$��TՒ��X�uS�9
ʮa&H���M6!�*eVD��WU#CB�Ԋ"���=5���:k�r�8zU9��;�E��;�����.U&N��,�(�FY�"rċ9Y�J<t=uhEn�DT^U�]�M��Y �2���赇TL0��s����;�㮮�FFg��*K22X��ES�C���)!Q$��Q R��#��{#��{�7u-���J������y�w�QT�³:�ߛ�m���#�y��U�N�ÊeM�hE�mU��ޚ5�-��3�i�e�u�*�dzG������'+����\?�^W���z���{+�}��Ԡg��%��Bg��|�6�����������N{��yH���b�v����_kHM�;������>=}$���&�,\T�B�|��<ub�z�8vɷ8<������6+�o�Uz���~[�w��֨U��}%�Y����l�]TO���� �˾~4u$�����^��~��+~�_��Bt�����r���y�h.�`��%J\i�������y��B5����*��W�!�v��o��!��{}R:��v�\9�� R�ԫ��a���w��ȧ:���1�#o���o���9��/�OV�q�����Vx��[19�)�ͿJ\��'�����"bS�*�_�e���*:�W�>��'��zg|O�J�8l�'M�!��\��G*�H��'aLǔ)��.{ƅ�^���S�iz�����>��62�8�����k���O�e��xLdoz�*˓�.a�������N}��2�M𝾼ُz����JL�Ol�5
&��U�����L�y�Z�0����r��iTkŠk0��O+YAC4^S��1YΧ٪#��Kqw)3d���Z�ʺ�m,[�t�\��+6n^h�v�����,���J���l���\����^������D��^:�j�HI����+��;�T�F{�=/-��J����R/�C�o�d8ې^�ú�n��DwEP��`�m�r��m�/j�Cu^��<f�4��=�וC8��@��.x�o_���pUnM�-k+=*yQ����O�n3�_�D��i-φ���T�{����v��.��U����`�V��p:W�ea���rgN�%9.�:�)sK��~��^�Tok�=WF$r�>3�6�fu�.5��}9�,{��*����+9�~�FZ5�c�T�NH:�B^���{�^O��;�]�}ݓ��O��Wu��?_3�}t�Y�R��x��3�n)�eF�B�����u�§vz�v��l��0�ȏz��+ԇ�Au��Y2�Y�O�>�*�����ʭ�kz�y�����z��b����G���g�O�w=�G�ަ=�}��qd���P0�J��y�u�y3����uE�kY�нFu�����]���.����'�{>�u�7�U#_��=�~Y
N!F����Wy]�wZ�Y`
����ځAO�VBʰ��w�qW��֑d�ңޓ�{}R"��o�:�)����']�a�|����n/?V���%w�w�Ro���Nb�3h���H��'
N<-����ծ�h>�넯\ݗ�@M��(�;"�/�[�j��]��r��\�݊�7�����Ĉ�6]uj��6&�T��ڱ]�*���s�+T,@wbj�cS�4��#^��pG��p7 �3"���>T��u�l�}�޿2v� ��ھ��7_{�=��kw����,�!�����x�#>�+#�צ]��+��.Y�/F�9�g�=3�%�Ld��E8f}&�S$5	�1Q/��d5�OqN��Ƿ-�^m�P�ޢ8y�]ȸm׉�����R(��0�Lk��S��z^k=N�מ8<�<�%��g�E��_ٷ�i=�~urn1�������>`���F܃P�Ĥ=����T�����M�{F��s���t���Ϸ���ˇ���F�P������F����
[>];�嫔�2�@���l�wY^u/I�yO���s�7�^:�����B��k-"3Ҽ���:��6|���;�7�ӟ��ϙ�vv�P6t99'D������,����8��>�s>��5պ��{��@��z����;����n����� O�b�+&��S�<��N�
�q��˜�sG1�u�Ѻ�/��^���~/"�Ho�����>�G,�)Y�xA��fC�W�^��<	YCm�'1M����ӆ���x��;�c/-Ij�4�̳��v��sz=pj�16t4��9KYŤ��*�J���cD�Vv�~�P\�춳:��N#"�җir�Z/Q��yr��&SK���A�`U�*z�Nj� ������0wF��%�3���Y���
5��{�}�~�<�+և��{h[[R:�x뫗�bgn�x���w�MW�A�����>����L<����}���=���+μK�A���s�������z+gkU�Nz#�����g���G��[���}I��:�O�{J��O���>=��U���H�V<�Υ�~��A��^���8 r�2���_��Yt�r��Bo��C@��7���ey-�w[z��v㺪�g���W������f@�,҂*� z`�J�K�FXT�aO�/e�z����,�0z6���N��w�=��=Q:]S��3%����/N�η���{�7Vjno�=��},��3Q����ߝ0���D�<gG����\ǫ=�W���#$�_	�l��K�u��m\��+����9[�	4�GZj�&��R���C5�?]x���0eW���oe�����bZ?��ϖK����x��]/�^ʏ(~wrq��d��@�ә{�*Әͬ��yrXe��}�j0��V<2��c�����T_i�ŷ�6��]�:�����׹�5��Y�����-ELUٓ�v���Z�JL�ԦÛ~�8e�1�N��8�ܽ�֛76aU,zz(�50�.*������ݡ~s3u��͌<�d����L��{\ b���q�T�ޮr�i+ŗ��]z1.�ݜ ����z�s��<\�K�e�ˎ�\=O����R/��yRֹ%a�����T�N��:N�f�����Ʃ�uْ�ǹ*����}���P�No��edo���~ͺӜ|N홏*�a�e{����R�Vn��~�Mwa>`�t�����^��w���X�{�(/�ٷCqΓ�A�x\;�~�"o7�Vk�-*K*�o��S7G̕p6���d\�R����}-�tr�{��:�+{�G��>��������Ȝ�;������dz�}�tNW��߮�����S'f�W{���{�R=cл��|2Ԓ�ߎC{;"�KF��ym��[�]�O���Y�G�?\���=Ko�����}K�Ϗ�Qaa�z�H<�"��J�/��s��Պ[D�^�ՆW���:��[S�
P�G���\{����y@�,�3Ĕ��}-�hj��y�o����x�\�N*�b����^����+cʎ�q�'M�_�=�$��2 r�3��J!V�w�k�+:�OU�o���.y��v-������|���黣� v��u��ث�2\�z{�+�9�����ϼǻig����Pȝ�/T��V����Q��i�W<����c��ՙ��ٮ�l>��P��"5��2ѹ������mwX��\���!�OhTv�U����΅�D�.��M�Z1VR���n,�1<B�c'J��]��7[���$�� O�3:�0hL>+xLko���L�x�zz�{ՠV�?H����̞͙���F_�0:�r�1�{�B���ѹ�_��B�����M�{��O����)����J��o��_��ƴ
��<H���5
f��K��u�Zj�S�%�#���Uֳ+|����av�>���xj�B��9]]1�at��-m�Ȋs�4h
gԧ�:A�wS�}���`�+�]��޻�q��=3� w��+M��jA���d��;�C}�C�Ys�kc+3<�%~�}E3��޴8_�ח��W��k��MN�{�V-{6�n}��w�!ڧt}=d[p��j�|��*Ϗ�G�'����\_����W�꽤�u��9�=�/��#��(�xfy����:-����G�&t��Q���T-��fW�
_�|R[j�i��@lMN�u}�b8fs^M�T=��T�-2	��_��?!���^�o���D.�j���fc׋�5>�(}N�/+��{ޭf���9g	H/�,]L�d2�����~K3�3��]�y2�L45q�e';��2���7�ei�8�~l��vH%!�6�œ_��^��'��ǯ:�{�j�AZ�����X������M�D�{��8�`�qK/q�Z#��_CA�ִe�	`D�4лʡAZH��6VjW^c7ѧց�����z}�νHyau�ŵ�,��x��a��T�z+���S/9_iӾ�}���fex��z`��5�<|ì�r��G��t�������Yc�+=�K�	�{�]��tA��uѕ��e�˷�Ν�O�>s�=�G��T��~�����{�6���o+�&} t�I�$y�
���YV9�+���z�8�w�q����U�\�
7`��5�g�ހ��li�|H<|��*�&@r��~(fB2ѷʐY�[f:�l�y��z����Xr��}3�M�޸=���K*Io�@༦�E9��F|@��LI���F=�<���&�����O���������Q�*��p��MB�!��OY��}^��>m���l��{�Ύ����Ϗ��ס�a�yl��w�e̶��%�nO��y�H�cxz@�t����ƾ�6��}v�F��y޵���K�=9�gj�n=�/ex'�W'�O�L-#=�ېV��.��:NeN_k��S�'=�>	����]:�7�i���|n3�.C~���@zM����Z������l�^�G�N�w�;���*ܤ{�O>�O_��-8}r ����)�7B�qt��'u-��%s�]�����/╃ˠ���c�V]\�geʇ{c��Ժ�[ĵ81ի�\yYO�	Xv�GI�ðǔ1=׫�Js+5)�i��5s)��'�_�gC�����*^��4��u���.k�a��OvM݊��)w�ͬ���c܎l�	�ޭ��fp�㓟�_����:/�S����S�գ����[��w�]/F��ԃ��5�+�$�y���
��E�mT�T�xyB|��d֕��}/v��>��u�,�s]�W����=��A^^��O��z��9�u!{��H��p����M�vTǔe��̊;����*��T�Ґ���tB��9���c�}Hxr�����#����f���U-��RO/�O��'�q�\��2Ѻ.e��G��}�����\{�r+μk�����w���ʞ��Ľ�5�y*�ײ���K�;�6XC�s>�˷4+��q�'���Vr)d{|'���u׹�wr���Ʈ=�Ӟ>@�,� r�2��
P5��2]?�z����C����'�zW���>����\}�'J�o�'}UL��If�P@�F@��-� ^�z�?w��|�ַ�TP���6{��t���x�7te�#��=�3�"[S�P1w&Ϙ5��׃��k�v�H^���M���^~*v����A��zO{��E>��=�5\xt��b볋y���q[r�|2f4���Bs���**����[���U��=�5ʼԽ5�P��`Ә�T�vE�uӒ�57�ӫ�G{7w0�6[�cMq�t���E��s���׿��G{�x�6�Y9�;c�҉���o���\���p�}3�d��X�@��n�/dT��<���K��>�&'�:2<.r7n��lTu���H�Wy�Go�ڢ��1H�*��3woym�����3-���%���񴽷Ȇ��n#�&�<ɾˎ3�w��i۾�v����j��y��)L2���p=8=q+N����W�m>6��ÅWUu�8�
}Z���.�>�C���S�~\�t����I�KZ�L5ckC��i�,�8uu����L{f�]׵�ϐ�Bۼc�{�3_�w�7�^2�}|,[�m֜��qcʠNi�r�\��Yu'g՛�*��%��,�9��_��_�K�^���})��X�s�ԅ�n���t�֮Ζ߯6iR�J���_�p� �P�+*���{īLQZ�.%z�#���o��s��8y�?`Ѷ�>���Q���U��_��ipTuW.Jg�1X\�R}ʓ3�S�L�2��Q|���e^��rI^���b��QB�$��aP���*g�b��!9��^/8���霟y������_t�S���6D�=�{�����w|;R���-?w����8\O2J��:�W�{ݽ��y�^�~�C�<��gse�׀(/cV���U�ޫy4XS�pcA"����k ��h]��%�&F+x�Wf�.�X��)�}כݩϧk�9�]W�ei�r�����Ȃ�Q��Ze����^U����υ�k�y-��Kf�[^�Ik��>b��w�C��8�Q����ǻ��`�,�<ITe�0
D�����"�޳�(���>[����3���xP��?^��>�2����d�+��Y,� o	�)2T��
�Nuk��2�7����.��#p���>V�s��{~��&���q�b�j6#<�W�����5�I�W�z}@�$#1ޮ���b5|�G\7�l�ޙ�>����h3ܤ�oz=�}_�����Z~�=
��s$����w��D��!WR������1�W�&/��uf��رrk9j��q<R�H�dG�h�~$o�'�j�5p`��=��o��.�?B�_�s4щS�z���;�U4��}ܮ�ſ?Y�p�>��bc#�"�E��.a��'�b����=�o�|��O�:jhn����^zk��~WxO�R>���ˉU`gxE)�T5�%��m�Ԟ�w��_]g�Z�Ʊg�Lg��-2;O��z��WLsu^㑯�<g=4=;=�U���ۡ��5�y�ڨ]W=<��ꍰ%�V�1��!қ�����˪������d��5�e�R��7B��������k�]X[R�8�k���3�\T��ړ#v/��2��U0���x�DB���N8qe����Ü끼s�2Lڻ�+h�h���Ǖ��Z9�,R�>Ш#�^��l�9[��:!���Җ_ث�-��B>}l�cr�; ޝ@f�%<�P7�q�F�C�����Rp[p��)�ڗ��-��U����7�`n�t�B��D��c��8�l�V��ٽ[]Mk��V�+�-\�T] �n�����H<8���u�3��KV��wx)Dk�l@����-V����ٗ!}D7�/��]��{5��IV��C0f����w�]���t�2���2���m5�w�PgK���dC����YQ�[ۙSa����bW�Yʮ��˫�����`x�Uu�#6C8��\�C�� ��u���v�S����M!�����@0��aE�2_` r�	��s44u��V`U5������o��(v��zŦf��Ň�J��C�1ȋ�wmݵX9���k�-'ٝv���{henA�e��٘�f� ME�;=�*�0'�g[��v�����nS*�hkc�[l�4��۱BQ��$\�k���kih���CB8���]�`��o����d��de�B�u��y���h�`�}�Zqee%:#�m:�Y�kVF�7�>�eV�hT,P�	���jM�Sbgs8��yr��6Vuh�wL�LViui�:�7g�w6�-V��C�^�J�y��F�)���|DKh^jꊭ�pF�Y�n���6��j(m�S��8����)��%�\�G_4^�,�L27[9�ڙ�>��K'r�̬s��خ�5���a����;G������hm��Έ:z�r�zZ���L�.��m�4+��]�� ��D�m.7�
�
ʚOk���M��3�_(#u��kh'dkv[άN��#xB�쭨��]WNm�t�|��Ȥ*���[�*�m��Ļz ���Z��P;���_<3�g
�'����������M��o�ev�/���\g8��/K��kf��
��q��r�˙���G%LuӬ"�<�1$uv-u�[�oe�^Ҍ+x7�-%eb}ˑ��<A��2,Ř�8�\����F��ݫA̭�Ԋ7��XՐ�%cO����kW6N6���$��Z�n�3�"��ImSƹl�[������p7�1�-ܳ����,���_E��і6�Y�{��oE�L�~���[}N���k�Ln����]1mU�ٻQ۴�S�{r-2��4�:�_u�ղ5l��{'%�"Z��T��A�{���p���%9ts�L�:�Z�z��΢tĥ���| ��'%�}6�&���p�Nk����A|�U�wd�۟\�y�8l� �b���oh��@�=��@�䷮�[�rN�G��m�Z+��1]���	Q�{j��c�ub��	�)�$�LETWZ���3�hDeW�Uvl*ȭRWqp�s
�0R�L�#*��	fu�Y*�*I�D).�^z�%��
喜�O't�qqNf���h�t���H�L���,���I�(�ʼ�ԹrB�DM+�L"���5$��S,DQ4�I�"�0�t)4MK��8Tr���*��Ut�Fk1U)-#U(�S�&�j���Th���h��J�UP�K�d���X�YVdZ����R\Ԅ���*D��	N����E�UAf&!X��:ԮI�*�
J��#ER! �4efl�2+��u5��+X��KDB"�4�$E���!R42D"0�I%�Y�8cNVZk3�J(VbjӫB�K0�����f��+%,UKB+�Vi,�)ŖKC+��l����|����?=9mvkd}��%�y�T�6#���3BTG�9V�]�Vf_u���~GX7\�=Ǥ��s���ұՅoy.��gD�#���j#2c�VSF����6�_�u*�.g�O�����UA���Zm��`����i��C쭣���t��Xd���G�-KB�K�T������{��d�S�>�-ͽ�N������r���.��kD�؎t�����Z�g��Sge��_)������SQ�]�ʷW�����_�`ϥ���q����1q��H�%+2�P3ŉ'ȿ`���)׈*���u��E{�頞i��C���܏z��+ԇ�Au����ԳC�=�a��_ܲ����X{<K�Ƶ,��=S-����<��|��{���s�D{��z���PjIg���q=ꙍi^H9��ޕ�Β�	Ƃ�ʲ9]��Ü���R"Yӿi�'�uǺ���ڪF�� (����}*������8N��@�,	��@����YV9��*���H���\o���|�&��+^ޮ��{�n�mǮ���24��(�=끸�����o�ʐ^�y6Vg^Wg?:���^�0�ur,��|��ު��,�*��� p^SC"������{&M	�������)��C���4�u����t��<�oT8wZ5�b�@��ᴳ�l����u�[wٴ�,أ��wu=X��^��Ⱦ=o�AC"*����n��
zţCm-Q�w�pVS�r��i ��Ig����/q'06���݂��*��D��{9������r�:ߕ�1�����9޹-�r�@���H����Gr���r�Ͻ�bj+���f��W�Q�{5�<�vG��ͺ�>���n4躁�+�'�|3Ɓ�7~)���V#����EDN��9Ex�^m�◲�?:�7����޿������s���Fw[9�3=˗)ސ}�%�8��ا[����9�/��^\6�U��$ǩ磖d����{_w���%z5]
�zFL���(���r|3~�zN�͕�J�߼��m��]~���4�4ǾI�s;�	��_i�ߧ<gNC?�����·'$�ߢ��'U���")
���;�޳��+��;������U�Y޾F/}�u��wn�ʁ>E�s�����p��k�������a� 7聵�*�@��W������~/+Ԇ��{��ڤW�p����]�����ƪ��^���]G\R�f��Wj��������s�����hxt�^�������2��6�$��3}������ω>5���*c�F|��p7��y}^ß{���r=�򛗟1TMy�8z�~��Z�	�͚�ra����	��n�,ӰҜv����Aj����ʾ�n�$wkN����������<0K��;Ad�W��FNN�ck�S[�K皲j��;z5y�zjT�a��Mi���/��I�d�R��ʙ�!�U����]�O��?�����2��UInbO�2��q���!d�^�ȸ��W��ժm�)�F�(��U����@�Yp����R���������ӹ�`�{9��IE�`�FӾ2����'/������ݳ�>u�0"o ��[�����+������v�f�+�U�3<ǻւ�:c�6��G�K��o�'���\S���!�-�<|}�ꭞ��ﳩ��<k��n�q��5w����<}(�8�'�����dUnIf��n�J�<�+�ٟq�w�"FJ�tn���P�SLTu���K�+��q&���I;��-�����>�=��>6�P�#����UԿ�B�|n��{!����D-�uG�3�>��s�_�'њ��Dx��s�i�ƬxT�lr����J��ڎ11�O�(��]Ig�6+|���}�N�y��G:�.U��S}�ʛ\�!�_��}�F�b�u�]7�36ߒ�~d�}�W��3��x7>ی~��}��񕾭�*��>'v�ǒ f��a8�mފ�宰\����lK^����H���S���#��;�V�����m�_{���d6>�a�)�M�z��}Dd'Ҧ*=J��ҋJW+�����Mr�H��9j��hً�̻���tظ�`XO�NBUvᩲ�+��r�WbY���t���N����*���2]z�n�ޗ��c��l��}�t6t��*&<yc����W��O��^�3D�\VUi�/ī�L ��#���^#>�Q��!�W3�k�Qq�Q�#{U�\��:w�p�������	�H���"�ؤ-�@W��@W�:^>��j�k��u�]���}���(�������/|먡�jI*�e�Bg����)��r�}5��}�4��Pw�YEv�%[>�}tQZsޟx��;�,.�ei�k��`@�$����Z��h�b�����5����Պ�s�C��8�Q��y�{������|�P,�3�|���A��4z\[Z�yI #����^�Z�(_Ο�FDy�y���GJ����߯���|R�~|;,ͼ�����XX�U�0�I͠>�U��4ny\W���Nv��o�Hq7��H�����D�����7�W�d��d ��Ćfu��|}hL>+xLk��m��}�>�Z���H���}���ۙ�@�[���Y�Wd�*IjG��J*_��_��B����ᅙF�䝧9�Ut]��W�<gX��m�sũ=�v[�x+���.��;8�gK׺�����<���Hn[�b�'V[r��]��1�g�U�xgZ�Am�Y])曉LS�47m�,�����۸Aǝw�i�a�L��"�]��d7V)�L�d���O�G�w����5��ċy>�Q
f�����^���1�jX�Nl��y��v�>�7�H�?+�1m�Y�m����@�|�Q>l��V!�/�B��=,\��z�U$�7�z��M\f�%w���U"ߤ9�G�> ���Ei��ѵ �O�K��:�*��Q�Y�nҬ�m�H��W�t���o}�lpΫ�9��q��2�=V==>��(�URi�v{Y��k����>'hDn�>���#qE�:nK�ε~꽤�7^�lE�}�p=��c��Y�Ϡﷷ��r�o�t;e�����^%�;.-��{���f,�]����F����QO�Q��z������Ϟ�ӷ2�A<T������)����.c}��d���w^�3�5�
^v�|�z��ϫ��{=��c|��g	H/ ����w�̻��v�|璧�}[!�X١�]�C�����S�Y^�<��Fɖ{�<I�5b0�[ˋ��ͤ�����p���n�|wR!p�;�Ͻ�}��#��RO�� ��]���}����l�Gѷ���x��̗�:v<=Z�Vy�z�QC\+;Z����ܫ+�nl��Q`��]�n[���ٻY��y]:}�W�i[ܝ�;�S�ͨ;@۶�n��Y�&Hp������Qtj��oC룴\C-Աg$v��j�άQ�d��>$���%*�Q���L��s�n*�ӿi�9>s�����rC�9���k�y��O�~����h<	�9 r��,	�u<[+�U��;򸫏W�#V��<I��M'�������}�N�~�\��][5qdk�qU z`7\��P�E�j�f��];�%��L�Tl�!��W=����)�!\�L�*�K*Il	 ��4c��`��yX���T�=��O�����VG[j��O��������Q�)�=qV��MB�!�$PÎ�ʤ��:���-Y���~�F觳K���村�?+���>���ϙ�����RVQe��vݮEw*גw����^TT��Ӕ}�y�������ԛ~��޿��9��%�zv<L��3�yrZg�;Мm�>>%l��;8�w���w�ҳ�.7�&|�����W��W;����'ٷLO?T����d˾���t>����/Iñ�+��990��&���]5����^�<g�ǟ��9����VG���o���Ӑ�㳷?���n_aAגz]?�$�i�*־�U�7�*���͇ebk��j71qm��>H��+����R̼�Q�&F(3�T�����0՜ܦ��0,��fe�ˢ�s�N�`���-|��^7�-�r���k����ځ�
ٸK�Put7�k���b�����-�-��~�D^�dxdK�쁑/׾+{�M��o��Tŭ>Kޠ�o��{�B��
٭��5��:=Ji��R�l�5k��^^�>��W���R�H����3�=S�L�W?>��Ȝ����S�F✀��ڡ�\������c�"�hx'Xτu̎U�ǟ��N�ǣ��#�sĞ5'�4eT;�(ϑ��&y�S>���q>>�h��b��O�sԧk۝ʏ�{�Ժ�Y�%����yL<��nb�}I�x��\/b�9?e�5ט�e��$�����RY|r=�|{ڪ���d��N��@�@>nP[瞻ת��v�=��k]P7Շ�MW��ã�6���*��d���R�3:���iA�A�<���7+%O��U�FK��䗱=�<����|����}��2=;����R�}���=�\S�N?�1�PY2񥴰�焁�0s�Q�����j��,#���ldz}H�g�3���{ޮ��^��4�̬����Khmz+Ц}2�%#����QȢ��_����b��5~�q����3B�߯�EJ�t7XEIs&��ʊ�=箼���;w8�fg�?
���A��e��U�q�2����f�F��LR��g��=�_���MS����Tf6uUd���M���x�f�Y =�����8;�S���iؔv�<��w-qB�F�������HDS��8�@����+����7�:ϑ�*pӢ�*_�ѵ������d�(�~�OV�w��Q3��jy%���3T6�CHFS�vX����Zt\S��wڣ�m�Z;�����Q�-����Ui���^��>�wީ��4͞%E�|�ևy{s3p��b���)w�����v�k�����{�25��zw�|g���X���n��q�;�CkÞ�ט�]y-줕zA|a����:�� ��W��u��r�w����c���u ��sTUυ���f�i�܀�����wl�<5����eV�Į����� �J�
>�Q���{5��*l�.����B���.��:�+"��a���=�Ɏ��-A�R���u��y�ǅ��=�4���aU�w�>U�������AZ�J��XUg����Bs;�3�MU�W鳹���þ�>��>>¾���*|�=��F�ei�k���A�,�Έ��uwo8�ug>Փ��!��������ϛ��i���\{��݅��ǳ�Yc�*�~��J���J�a�s�I���*(�B�k�o���CEy���'" ~g_�<�Ɗ~�Ra�'Y�Ո���v��Q��꫚���-����Lu�����=#]u*��p]4z�/ ��ǧna�t����P��M6�w�:��լ�w��>�֖���n��9k�����i"�J�q�U�+b�:~�}^eo�*���鿟���Q��_����rĻ��x���(ޠ+�ҼUd#PѸ}�qW���3�;^G��z��e߻L�P
��t�����k�7���S$��D�4H�����j7����m��C�ԡ�ͷ[��=����q��=Z��@�U�5qd�*Ijl��2�HU�K�s���|���V̡3�o�=�+����ۮԛ��|���9�|���l���>�S0ՅX*\�����M�����w��	��^���/Q��w&.!��2o���o�ڠP��>D�d���c.6��J*�Y0�����z�z�ǥ�މ���}�LrUV��w"�����z|���+M��jA��C�'���7�_"����	�	�0��n���ͦ4,��c����3q�����^��&�����t�j\g|�m�����v���F�����7E�:nK�ε~��	o0;^�1Y��;�5W}3�oU�r=��2�ފ�^�V��/����x�Q^%;.DC�k�^vJ���dqj��-_4�};:L�[y�i1��<!�7[ɫ/e�T�mn:s�E&{��{g���b��wyK�{<pz��t��q��3	����Ke�b%wuw̎�gs�"�ɶR�>ܤ��K�Bo��z��`�LwWu΀7� k�u��Uv��S^g��V���{n9x6t�)�ꇳ��uJ�;��1w��!�����]�TOd�[ݯ�)O�� �}P6���^���7�޾f/���r���X�]���i�w�#Wy۾Y첇��yD2���k�������O�dW� ��kjY���âZ�>0�՜��q��g�c�2���h̖�]V7��=�����#�~���.=���P�8�w{��Wr�'�'��$���8�a�`����n*�t��s�O���GX��"��Vu-��w;��mt��{�~Ȁp�_9 r�����@���ϖU��|��◹{���&s�ͽ���I,��}�G������\��M3Z�Af��W� z`7\��Co���6n;g��۽�����%^=^��g�z���g��~���UW�Ie*�� g݋���;*������{������+#�W��G��Ϗ���P(��CS�p�{
��be����_^ ��%ي�ޥF����ZꆹB:m�b��Է��nF@�?��0`���1���6��m��m����`�6ɶcm��l���{l���`�6���`�6���`�6����m��m��}�`�6��1����co��`�6��m����1��]�cm�6�1�����co�cm���e5�Z<v�^*Ř ?�s2}p$m���W�i
�Rؙ�YKZ����$U@�*�l������*�M�A�Z��Y�f�h����U3iSF*�lĤDPɓ|���wu'�ug�sgn��p]�W5s9\��s�v���6�5mI�aV�6�]��:��m������\Эkj�297[�V6ֵ�%��R�Z��w\&�u�@����3cjj�͎��j�u�]0M�ӭ���)�[V̚�]ͬ�N�i1E
�ťR�m,�&���;L�lj��wJ�V�ʥ��[Mݶ�9�i�e��   ��}�4zQsڹ{6mw���ԏAݮ��މ��]�K�Eu��ׇ��n�=�p4=Q��=����u�t�Ѧ��p/g������R��iF���톾   �}�q��l�=�;M�{r��Ol(�yz��(��-�N:(��4i$�rq�E4QEo�����(��(��;�$��(��#�n(��(��(����$QEQE�x��_n]i�MYVM���6}�O�  ���UU]��!�Zk&�����v����磝���:��X�G�WrG�Z�N{�*��wx����ۚ�k\׵U���ֵ�+W�er�ѥ|  g��5���y�����g^s����c�{5��wp�"��n��Ӯۮޮz^�ݶ��%�=�	/4���������ٻK=^������{�׷U�ЩN維h�/wj[j-�NZm|  ��;�v���{�=٪i�u���5)V�ǽ�=�ڝ*�����k��v�ut�V��m��[i^�&��[ٹ�VZ��vz�Pt罵�z�m���3��f2���3fm�ͽs�JR���  c��/���k;��v�����Wu׽מ�[j�v�Ox==m�nT���g��tOs+�׷aU���νڷs-�n��\���jۺw^�ݡ��a���۬nt�8��[f�ڥֺj�v�Z���  ޮ|�i��+�V��S�"M���ѫm����޽���vU�ǵ�R�m��=�{���-t��sw^4�Ǐi���^�
Wv�/.���s��ko�ouS��䞔�b��e��֗N�[bo� ������l���p��@swos�@�����S:��ܡ7���ӵݻ6�k�o=�󹭽��T�k^k׻ՋY][��v{]歋���y�5ۻ{���f�Z�p�e�v�����  ����N�Ԇ�y���Un�.��Wv嵜ގ��yT���wy��v�W]�����%�O^�z��V�!cs��ͽ�۶���k8����1{��+e��ՋyZ덬Um���٦Ŷ�m��  ϽS�-kl�t{��zum[n����oc]A��=z��{m�59׫�R�e�]k�\��
{ںS]��{���R�[m�s���k���o4t�Op;7W��Wm���O 2�	����$�T��41��MT�@  S�A*T�`  5O�M����@�J�M1T(@��#����r�������0���������5���Wٙ"��n���{ޏD{�w�c��zW�QE?�W��TA_�"�
ʢ�y��n�������~�G!��h�)+f��D���J"��Ғ%�����a[�d�|�'�����q��ۏr��dy�`�M��1y"�)^�KB*��鞑�O%<fTˬ�ot��z0\�'{]0������p�q�A$����<�a`�N%/v!��y�L�k w��+v�R�#	<��o��Sɲ��� �̌Y@�&�C�W�&L�[�.��[��T���VQE��Dj��=��hY�K�j��@�W��V��A�Kq�.�j�ɍ��k������,0�&Z��I�^n��K�ȧ��6��ֻ`�a�me�(%��)'2�
H�Zj]m*׀5����
��pŪ���f���g&��m���Se�w6�)5ն��SN��v^j$�KP���B��4���ʵdB���)�t-î����N$I�x׌�Ń>G�:W\�8P�q�phQ����L��>�2�t��[�����[bj����rc�t�W�ژn̉��[R�b'CA�U��:8n�Q3@,,���4ܦ�׈���{Zd��ܬ���Q��f�3d�K���Fnʔ� dݤ6�+��r�lDS�k΢41Zel���jЖ��Y�!�qhc4�y)`�q���hg-l�s;|��C�yf9��Ū�
ٕ��j�}R ��fM��)�Vf	(
����/)V���P}��� &H��J+)aƃ,`�'00��9}�O��>-�{�`�!�������Y��q�#��cP�,��e!��.]��\ɐ��iY��b���#������Ě:�`*��N�2 �e��%�SC�)�X�k�oJ��)�֋�Dc�*�-.^%�[���b!���銃EK��N����r�����)e䧲�c�IE����"'�=�E�{�ic'z6�%�����y��*���[�0�W�E� w�B�&��C�ٺ7&:#��Z��(�g3 �5�BlO#�P��/N6�@���,+�2�[d��n�	jo!.�J4�� �s���*�ʣ�id�aX�cִ�ɲ�8��h����
�Tڍij�T/@�kLF٣X�r>p���:	{nmҫQs4R�ݜ�ai��n�:c�7d�z��^[K�LM�캖m5����mӠ�(j�ރX��+u���pĈ�F^��tb�+��qa�{��6�W�)Xts*�U�c��w�a*|�2.���T~��MpK�+(�Hdr����x%�ww6V(���q��9��
vŚEX���E�Եi톰U�oL����Y���G�g�a�Z����g##�kv�uI�]��$�A��B!A�/U�+h*����	�K�)�Ghl�`xMf�u�l�&R�E�LF�F7ml��w���Z�Y+�#�y����F��B�NG��gmE`md<��H}S2��B�UU�d*	۹�[VMC��,�*�jљ�2���V�nH#��vfn4fmGp2�mi���c-�i�a�zz���&��܆J[���h���l9�������Z���oj,u�s`ӎ�qS�[��H�e���;dnU(���{��rb�����m�)@I���n���n�,�&UȮ+�^��ă
V��~��v�3Z4LgD��r=ojM�m���q$q=H���ݦ�Y++U�D+օ�f{OS��[�l-��ꍫ��'��]9��&�f��{��LfS�
I�H�Co���x�Lh�h3��U0�jj�)1�j�ae��lke�U[h֕�ǖ�"��XI��C��c�	�n4K���-��dC�nX�&m�l��e�/h�KV-E�ٹ[���P��!�.�qA5iX�u�H����Y����]Ф�A�)�q��mXehY�9���� e��he��н52��o&Z�m ѣ0�����P����
\dX"�����N �SB��e��&`�L�&���ř�f�ĝ�~P�y���$&}y+Ü�>м);�$�Ď�{�5�eJ��D�E���Ig$�j��� +���	����M�Y̬iJv�ʸ�#���ۤ.`[*V�n�l���.�҄e����ճE]�`�P-d�)�aC#A�z�CS߮��j�)6JˍK�)Ͷ�u0`��tn�,��T1%z"9R�ܼje��U��O&�n�S�w�=)|��\�,'��ԫ�x�0�	Z�R�a�Z���{����`�-�>e�-�۷C����{�Yn�eҬpTt3q�G�[FYW�饗�Mܦj���sZ��L�E�H=
k&��wygF�IR�S]lU.�9%<,�j��
^�,�5wcRx�	Ȓ��PW�]�l4goek^'7,QlmaB�B����GGlx*=rnK�	��j�e��^}���cܬRV&����4T����x�2H��n��Z0*��@DHS��Vd���H�䭱�X^°���Z6�ɶ�O�0�*�h-Vs�M��ZJ���0ܲL��lTK�i�Alm�u������mB��z��X��� f�nlZ��g(���(a�Kű��y�%�g�Q��`��%�bݛ���k�I��8��ɍ����¨����jQ(����U����9�m����&�%{Ѿ��
��vln�W��tVKWb�$1\j��:�9jf�I]���݁W([y4��.�j#���{���(��ݹ(�&aT&�Ҕ���V�� 5ITک�3�Vм:����>vn�@b"X��T�7��^tr�����{��N�;�^f��=ֲ��%��e���L���bm�l "���7  o����;yMʎ1*#a�N�["���͊%��ѐ�L��bm*FŊՒ؀PVV��.������&�-��1J��Y�Vث�ɢ�ە4|�ZbC��x!��/o�~����i�e�\Up�J)&��Ϸhfk������(!�;���E�V���u5�2��)L���1����Y3E���v�Xߊ��QN��z�@�H3�xa3%��EV���J�yHhڏi�eZV�]�jMcB31�4�5��ޖ�*m�%Ke����Jz���5q��ʴƦcګ�L=:��B�'�A�q�21�hP��IHD[��\rm�o(6�#�$fd�q���w�* �A��xȞ9��8d����:f�wXi@ �/�t��*H��O��Yl�ɦ����)�����M"�;�1z��sUX{�����GF��Ӆ�hݍt·�oZ�e��TP�&�)Se�V
�׀
�T�)�ѷ�A�ю�k�S��X�nU�4*�C��M��b�܊^VP�ay�q�i�(���4vL����L�@��[��)����s.�F�a�sA��#��3� #�ګ8��%W�2E���U;�rk;C�ȨJ$�-S�(�1L:<�V��(��-G��F�O���n�����珧aѕ���O)���쬂�ٔ$�	��&�en�R� oo1m
��V��Yq�-�&e�Y
�Ԣ�w�4j;ę�X��(G�ӬVW=��;���U�;wk]��1�u�EH>���%$%[�
� M�N�l��mBU7K�/1P�4%��^�[o���V�Tf��$6$X)�9y��NW6�e�!*0�ŰrnZ�t���8��b�IH��ʛ���0�3����==�s�j����^N%N�����[R�m�"^�rQG-R�e�TZ��ɯle�ݳI.=�}$��N�i��-57PS�Zu]h�cT���'��E(C̙.�黸քQ�p��ϓ�)��}u�h�]�w45H�!�^G�'<�g�Սbt�t�1���^C�I���5�`��Q��={&�3J���c����c�(���-�{J�'�jւ��z.�i�sB@�eY����kE^ N<�Wu�����W����4��([�H"�đ����;�,�jf+e�J�ּaX/Hm��m��B̄�J�5)�
�䷻�`P�~�2��ԫ6�Y��+C�e�VA�p�ǡ0�L�A�k�L��A�Ƙ�(M(�'�����҇  ڸ�\@�v���sin�mU=�2��hT{���&��&t`
jI[s%=�ƻ�pa����4����l�tTjd/5���K�u�R<��ŧBeQ�J�f^j��M�T��j�\ �]�����4�Gt5D��ᛔ6�ST6����A��yxJ��s�:v��:M���ƒ���b�,��7)8��&�$[pj���]�v8E��m��t�u��ʓi#���{X��k�'t�Sm4����2��Vp�R==	$��Xw�s�i{ݜ��!�1�Q�/�$�q��O���r+����6ZF'n���#�ݤ���/.��ofj!a�.�"qQ�����"��;ks�Ԯ&�4���[tsC��[y��a�,r��Ϧk6C)my!׺*�k���̻��%ui���Œ*tkB"�&Y���7["w&�d�4�Z���#Ol�	"��ʕ���CT�:ש����q9�d9J���ۥ�ҽH-��U�וm��	���
(7�⇷�^y�qse�saT��u[4��׋7S����\�&�ug��"��k�R�O� ą��Р�Cf*�Bb�Jn�B:�5�1|E�����in�F�&�X�j<N�i:Y��6�a�6�	I�1�P�jҨk)Ҽ�zb�q]�{��-U�$.�F�q���@i-wf]>Z1ˣr� U�5kN�CYWD�*^]�ku	��Up༨�k[j�Էp+�-�� ��,�I�t�
���(���m�I�r��6����vӂ�+'��n��j`����Tl&�Q���A˃.X�6u��N;o �ȑ�Mˤ�ͬ�ᣘ+T2n�y��A�eʓ�{H�-����y{)�l
�ܖZ���k7-X�H���ݑ�X�׎I��9�p���L��Ӷ�]A{w�m�v!M-w�15o.�I�q�S���7ML����%B���q�FC���Vf��	4���6�15g�P���N�kkN��\���Vc.2s ۙ�T�d�t��^��=��hR�/`˭67F	(3V�E�5�2��0U�{�[D�ݖe���"�vE�I�d�Pj��H^-D���HYL�fG*�uV�F��ĩ�WN!�����A��B�o]�#�µgh��������Q)���\q�̛>Ɓ��v�t�ڜ�b���֐�Ojh�GI�ds�7y硫��>Yf�"�Uɬ8o����QQTo\����ILW�ʼs)�
�����Ij��e�E���K�u.ي�hRH�(�ù��5����ͻI�,���jQ�����FF1=�1��������h9*֝J�+̚�� S9/k&�RléBX�j��M��D��5�H���+��0����daԓ5c
���#@�.ց�ڭ��M�����Y��r�k�l�w�1�Y���mK���ɖ3Lȱ�!��P��%dI,GR��K��L@�yt�8�w0l�HJff\rY�}�e,g�WӚ�!"�S$MHi|n'2革�^m�rw��*{���2w�p;�1�BГT�[��&ۻ�of�"	��&(Z��ӧ딈�;��t��.���ghҕ��e��e�(�R7���!��F�]ɉѹL�$vs6�Dɭ� �2��ݘ�)h�D[��c�Ա�!�x*d���;���m�,��S�)Tͤ����i�j�f ��s*�`bXKh�
V�B]�l�ӺU<�.1rd�Z�*�f�h)XŨ�����p�0�*��J�-�`Te�^%0�`V���[{v���D�k�"���.��&�k��٭��7[v�É1{m�j�aI-0�vi`�.�ٺLj^Z۸��7������5m��!���3,�+Ef	0�b�kP��
�c�CV�Z*=5r��G11�IՅ+DFƅ�^&���E뺼.�^�2ք���N-�%i�Ԟi�>c�҅]��!��A[�a�e�r�ӷ(St���������|�g	�V�{���/z���q���Ķ�``�Vk&�[�Z�8/^�z��Z����T�Oni'm�\�����oԧ1]^5u�3��sH�+R�_��bj�4�;�����M�Nl��3^!YN���'�S�ҶZ,��%	m+j�8FV���ffXV�"�0B)�[6�&�^��S��㕸���t6����s2�{�ѹ��A3�j�kD3���Rڰ1i9� �MQ�C�� �v�/�{�"��X�ϥ��qٺ�-KPC��QSl���3�,'�h�#�5���Tǘ�ˁ�U�q&ʘց�0�f�쫘�4@EA��$h�x6�W����V�T����(�8�pRk���a�\�e���]C�1��rP5�Tз2�A��QT)�+`ha�{r�4�85J�f G�x��0��Z�Ӥ��
�;�v��,W�<u��H���	
a�V��-1���e� 9�m���v]Z&�@��SkaHǁ��ӇdB�p^\Ռ���,ٿ,�]�3F��l�X� i��Rb�Md6H�e�VU#B�Fm\���Ƈ��Q��#�D��q�g�|��sF���1�J��53���^Ye�+`��l�5�L�����ͫ�we͌;�i=��L
PGGqkªf_֪�m�Uddf��{�Mz��Ÿ)Qɗ3)X�P��M�+)�xPR��^|aj�鼔VX�(e�5�X᷸c��,X����[f�h���L���۞"Wn������y^��M�L�G�pV�J2eL��4�8%=���"�*�Cղ��YJ<��6��ݮ��z��p��C� ��z�����\F.��),��h��G���GL�`
���k#�f^VM9�^c�@
������]%����jt&9i��� �k�^`3�[�=�sȇ�-��S�z7^K��@�2MM�D�K/���ŗ,S�_wJ����Q�ŏ�2ͫ�����և����Ɇuqo�5`j��!��6�)v,�]m��a䗻$��vt)��eo)5���o������o���WH#��[���/xx�ex>h��u�{��qZb}�n�L��A�o���Ԧ5�cV�k.��Dv�����!q�^���k�k��o~�������l�����1�K9t�<�M!e���
%ٹ�Nc��[d:���aZ?t��%
�|�_E�|���Aqᛱ֪7�ul�{�[p�5؎����H_S!�,�셋��Q���)���`�=�����:b�6Y�mp�R�܊ZB��.��ˌr�i3cDJ�z>�:a��m�H�auS�������Fw{4�B�ywQFa�푌֜��[Aʿ��X
�xֳp�S���om��L�"���p�M��+�-��w�u��;x g�˦��=<P�{$�I"zC���w���֓����am���11�F$z�� 6V���9��Z�X�Iml�\�:�Ӣ��C��[{i�+������T!�6]Ӿ�sGL�6�r��v+�kY/^��i�эq��Fa�r`8��p!u�
�kK�ilN)m� ȉ�3�ݏ�3aR�Z�Q:��\���諓'��"�V*�HT�{�6���{Gjс��d1�I�W.MEF�K�6@g;k<���u�n������{���m��sޤ+l�4$�oEZ,zЬ�yY��$2��4^'fh�*��c�N�"��h����|x:���L*oT�X�Jl�U��8�Yy�K�+6��O��Gh�9b"}�P�y-J�ט ���^���\ىc���~��Ʈ��eƖ9MK��qQ5��+�����Bg����0��l�i�U��i�%T�W��Q��ׁg�O�i�~�*�������E���f�R|�M��HY����_G&^u��L	c�γѝ��-�$�=*<�<n�m�T=5Hv�Μ!.����x�d&�^p�EX��'���\�[�L����:�f-�̈����S�:9R�%[�y�۝C%�Ӏ�}C���C���G2<��XYRdj�I��آ)�A���
[���t@�
ȕ����f�n:��/�/2�N��L9��̀)�ð�"z��x�L5 �=)�M��p��I;6�u�abOU�.�Du� ��Yjח�H�_��/eݔ5|ǹJq��˗��Ȩ�DN-��g�TX�D�kۮ��z�׌%rP�YP�U�%�^/�C��R�&v�����;R��9�����3�ù�pǗą}XB^�~�U(�Fм�+��ski@b�6�4oJK�֭�{��L��ý
�Kj��EW`(�o#�6�%��7¿e�\�����y�D�ъ��U&H��0L�Vc�����\��۽�Ir6V�Ah3-�����l�D�|{.��l��Z�<:q�\ۡ%k���09X��aRb=*0)>�Z.��u�-�B<�A�7t�#.��7/R�otV�BŜEho��s_����|F��o��Ь��Hy��9�,X��K(fim�
�FV��<szMn�%�[G
V)�At8.� 8ӱ<{�Q������T�z�*Y7O�a6L�'QFBҔ�>O���
��p,RE7�(4�3�Z� W(L��g��n�R��!ѱ�W/WnIl�uU�xX�Ml���Mz�ܰ:�]�$��w"/�ǺV,O������G�B��-�)�pr��}!:��K�,���U���t�}�4(����;qN)�nGp��}����g����!�$80NN�H��">�l��:�Q����4'�fq���ů���O����臎��nʬ�K۷[o�n�IK�R�a��OWu�<W�.P
�L�v��Z�B+���$jNSD�zY#�;�)ID�&�mB��H�Z)������Q��hfs���S��ۭՅR�+{��i|Mۜ����6]f�5uUN�����I��Ï0Å�3�`�^�KmR�A��.���c���5L��Rm��wf8p����.g'v�'/���a�f�S0Ȯ����}
��G{P�f��7���}��|���6�>�U�g '�u<b��-e�f�p���vN]�ha�9/���Z����]	5��1�72�\Eϊ�ED�e�|�WR�qn��o�p㣗�<����+P��Sť��t�g����F�����%.��J��9֨8� 0�/(P;�˶�� O�W�'���@^��˅����uD�����p$6�.�P9�'tX�%fƁ8�``&f��.�˄Hc(o*g1S�Qͮw��D��U�E@T��Ԝw�ݖ����Н������u��M��PŇ�c�`-�fEN��F��|6�P.�/.hIN���˅�(䢭˯�2d������/QU>��H���-�s��ӗv��O�bO5G*/��7Iw,,�Q�����u[�����.p�y�/ag7����@�� �Y��g/)a\q�5ƧN�,C��^ ��[Q���P�сϣ�}�"�(0A��I�$�rf��gyl؊#hPÖ�Ҟ�4��&I�i��y�`�ulRSLX�ޢ�������Q�]��,�7b�r�"��J׶^�rK8�n����[#���=��Z{/O���A��ⱑDP�"b�f�Nh������wn�T�����1�
��["�HZ�7M�?v��`�uӏ�@oa��/���x	�@�(,Q�Z��wIR��72<���S=h� ��^ݴ⸴��D9����ų�p�����q��7�<A�]�xhn񦜘1�=�D t�ιQP%ۋ�Y��i&i�C����$���z�3�3ŨLa�u��H�T6y-CQ�N[��˛���%aV%��L.��%Ѭ7ϴȝ"ɭ�h�J�u�r��|�w���ā�̴�v�q",��n�<;]�9�4U�:�e��E���D�"�G�f����c!˺D/ |�߅LV<��3�װ�S�����U��)�77x�`�>�@��R��	QR�W�x��J�����j�x^*C͖��T��ZcfgW.C���Q�6�HKU��{�c�����e1]Kئ��.���@�m�Kms�,([I��˨�_n'J1�v���Z�޶N�Gh��ݒ;�j1��l��9%��e���'s���ս�x�jBAp!��L�*g-��;�o[�H%6��`��������6���,Ce��g�w�/��6@�{��}-h���{�$T-j;�CR���r�����&�^�:�P^�OY� �qg=
^���<Kڗ2�iq���[{]�.��g�����@]S���뀱�^���|�d��X�-��1�<=�՚F�[Iڠ6�X�����:��4�*73U�7W4�u+].��r�©���L���I�m��ԑDkk��G{v�s�3��au�
j�Vs�]�s�1u�h���ޙ*��t����T��V��N��Jo���n�1���S���bnV�-c�1����;*]����!��vei���e�B:}i�<�j0�Ϫ��Ș��֋nZ� ����r4G�$��E*Z:{�V�j�K�NL��T�%�43��@�`�L|��w3E=��h��W&L��]�e�t��1�,��cd;��QF*�q�ǹN�I�01V��� ��}���=3���%����<�dդC���wn����Cl���3N`�M��(����d�Rţ ���ηA3"��S ,=��e��nS�%,��{hu;��Lq�֬r�|� ?7]-�u9���;/M逓�ʥ�9��(mm�������Ƴ��\�w{�ʛD��f�@ON���w�F��}��I�Ԧ��U���V���Z㕺�<���G6�/��cG}���K�>Sx�'&K�4&7���Y���׬�_
vS?c\��N	�R@��{֌:ӧ��߁**�H�n��7����u�\�w�gq)ٲ��^J]��Y�R^��ubI��@�Q֊�y`qA��� �0��N��ݎ}��V��S���h�L]��X�*����-`�q����y�ɵ�]���0&�ˠ�C���"��d��-Ma���������F��D�,�榛ݺ��|�L�f��[`����a���`oc�C�kQq'J<�t	X�7��;Ġ��u�͊\��vf�߈��HJ�p8�|̻%��xdE�F���X:�p*�o$V.�5�l��٧\�yo��/��'�����ln/JF�*���rΡ�eZ�C%g9@P�����q����y]x;9�����t3;��I+�ĳ/�YLK�.��v&˽j�!�����N���)B��+�;��]W����&5j��%�W	�Z���v<=i͓R����oXy[�[\���c�X9���P�R۶i�M�I��H� �H��k��O[��(�<,�S�j(-�ç��b���F�������E�����\�ݶbטFy-�ʶ�zMZ��^�o�5z��Y�z�@
9�Tv���xu���Uj��q�=�c�������1B�P�p�h�H�2w��tD��F.�<`�C����˾��	a:7�OQ2���'��h�Z�ޝnn�����-p"��Ѱ�-�e^��^[��\�u6�"*�wҥ�X�Z�ցu�j�r�}�s�	`inﱫ{O!��߆��si4���m�'��U��]./�9�f�\M�7��U0ɷԈo(ڏ7\� �Ti��[Y��-�tr�n����mЊ�̩�Bdt�i���<&t�����`�"��f�\���E�Wޭz�*n���I�PkYw�3�sǍ�xM�*���f�JY�����ٔi����cv�N��6RR��r^K����*҉���[莍4��B���ҫ�-�V��ߍ%��$~�O�ݺ��^�,P�{d rJ�Cǽ��������i���US��p�瓊7e*��]1\���;��<L���iƧ+5P�^��c��iv����C�x,4��nu^q�
|��*����Mcn>�v��v��0!�I�R%i}4�<\�z��:��ɶ/�=�=��%G�*���W5i��I�r�#ٙ�J�� �Z\�1{�[�;�����FC����w���-t�p�Z�쁫>�I�l'���^ݖ��}شL�a��^�nud
�h�ZQS��}��N�K�:Ua)�tt[�f���Bt2��)z*}�q�}�g��0��[�s�Ӳ�RgV��F�>ŨU���u��ѷV��
=��:���	o�
�e\Y�˭��Ug�PX�-rC�8?5�#|�q�o��\�f�=��2��������
y�H<lva����#\��8z��v�ū$��N�0<I��_T�o*l�s毷�jD�ƈ�������w�E�ֹ�V��2�2��]�!X2��p�y�uH`����&�?�i��e�]�.�
���J�Q��B��T��+�
=Dl:�L��k��o�ЎG�[��V�_/��2c���u8Q#i尷7�C����._[<Σ�v���q�d�u]��)�u��/�^�Â��t�b��b�Ghm�
U�[��K�ȍ���6�1�ol�P�Oٺ�:���p��㸶�u�O��Fo.�M���r��s��\��& ���Ei��󞝗�&*5�� ����g媭}q�I�G,a4E����3���A��(�����üy�O���J+����8B��Ω\v�5���T��O^��9��\�ň��"ժI���=�.���Vɻ&f�<���u��OfN��}�ԫ�v����;�M�9����O�;�މr�A�^�c�]�9v����w)�u˖��R#��HuѼ��a��k�9��0��N|�`�� Y��ܱz��m�Æ�iE�����(���I��k��:�*}X�t1�w4�V9��r�Ɛ�:i���{�H+9�TO�8�}��Qr��)� vO����ɾq͙;_;�jJ}�����/g6{�]vS��W��Z[���(\����>f��qlFJ#fS#:S5_V�U(-�-q�'2����d�:��I|�D�:4��Ws/���z�=�,�`�d�hOa��~���!��P#��zv�p�[�hӆ��iu��=���yh)#�ͱv�`�&��S��uN�<y�D��,�I��ʒѷ���W��i*�{E�x�3|��m�fN�C����̭���mn���R��X-���QH�Q�X��̕#���W�!�潐#�������k+G�f��55����L��v-�t������zo}�Ish�M�p�׋�<^��^��{<�m��e��-�Yˈ,�F��]��p�����®����U��3�������;܍���5��K{[:��3ó<��b�� f���ȹ�-�W�]G�/����A��A��y�mЃ�Qɽ��o����k/���mL�͎�G���[i`%�����},���.'	��#����T�m7��!����콭ꁧʸ4�R6�9����j�/$6��vv㋥^��qT�t��g�-��:.h�tʂŻ6�;��+�y@���K�{��z"=����ޏ{��{�k_B��ٌ��f�~ؾ��D����	xMU�=8z�el�qy�gh��� �b����h��3�ev̫L��7Z��E��jWaQܲ�ڍ���{ae*�<Oa&B��'��	h�����Bz�q:�,�`�6�S�H}���tG)�X��\�h�f�#�"}����͉�b�f���
G�:��_Ǫ>V{�.<]�k�kC0�>�(��R��N�{:@��@�|����Z���=ȋ
�b%E�w��G�Z����}�݋L�ie>z-�gOnrD"6��n�W�:x�5�:u�HǮ��pofv��^@3�\��i=�*��ʎ �e"��:*�}��[�9�$��jn��\0��� ��e7tG}�z�Yි'0j�W�wdɳ�hqH��ߞ;<Rr{��XA���7�p�2"���`����N�.�@�s��cl<�Y�_90��]L6�R�oj3���[ܾ|a�>�uؼ�:i�Y��w*wئZ�gk5ru�(A���F�����k���GM舾b�-���vo���앷�D@}�	s��v�:��8����H�k�hx�`*���I��ܕ���^ �U�#S5�0�>l���3Y��)��$x��h(m*����t��QY_v�z��d��-�wu�[�j�I���"����s�]t��j:�嚾�:UGt�T=Vwց��I�9���b%R�׌LIx�x
P�x[�)F{~��=�Ro�A�O���l��\1����f?= �Z�
�$��7�P���ܖ���`��uB�(j��.�����;nR��y���}�������gO�,*�xpg�0f��O�,U}�W��Y�o��2�r�Q���w;GG݃�'�ֽ�/��w��b�s����VC9�S���\�b��:�`���c9�ٽ�!��s��SN[V��Љ�qP���<���,3N9�kO=W_'��Ź��N3`���7�LVX�QC������ݹS4����4�8�H��Kh�� Jo{'��y��0��_f�c�����Fͽ��n��k�we0y�4+^�1X�����S)�P��d� �^��X<��W`�v$+�'=��.�p캰���zوJؕ�|.l�7<4>��Z��x���k߲Ћ�+��T��%JFn��}��L+A�d���^�hX&>.�#^��c��Z&!�����֗����8�Kv�"\����zqE+�v��%��L*�vu�zÐ��i�)O8�wŴ$�1�󾰗�9��즦B�90ڔ�dw�����#��I��U�ѽ8�u���[jv�)��E��u��g4e�,�}J���-�,�Sg�w��`Sg M�7$oO��j�t9$�7K�p�뵢�s7�V���]tAT�jM%Xӷs^��h؁F�"3���싐q8@֋��qTJ-7@����o��F6�.؂j���N�K~�.�+"��)��2z�E�m����7c�A�l�J����To"�uM�άۦ�J�u�4!c��J�ʣy�Bq��,�;n�;��.�,]��b�[]svg�h�  ���;�JY��"�j!D:������_7(��{* u��}y/jelJ�y&�3OK��l���.�7D��}M��*�gvj�u�phS��\
��sn@-#6j�����d��hQ���^r�^<��x�{�2F�l���o��xj#�U���h&�`�g[d��zW��c���`��J��醂�ٍ����rȰT��˕��XH*Qsmʽr��*/{�g�=�.	&&Q�%x�x�B�@ϝŻ�D{�E�+�t{��yϯ��Z�t�rMj����}J�i��`�Qvu��>�QR�:I����sy|ӹ�]�F��>�L<f*�MrN�����T甊���4y ���7�e2t$�t��wEYۋ��`[�:0eH��	_�5�V�C(WZ7qP��J�l�w��c#Q�{Mj@d��h��,R��H�!��x���nݞ��޵��-�/�2(����Vr�z'�F�z�LU���b
DI���ʅ�oF�i�B ��U�V����޺��{7Hؽ��͕$Ă�c7/�x�p8c��.Ǣ����Z��]��J��k�� �m��q���E{�on.�1��2�{��d�k��k��n�\"����+�Kє�<�*��Q�)�s�#�:5���f��/OM��e����A�A��Wf�74����љ���GroE[%dxqeϾ
���=y����Q ܙ}��&+�N���M����h�o�����N���]��$�G��G�UwN���e�'ae�_�7�7Nr�XT�)���ﹳ�
����rZSͰ��p���^��o׻j�h?Q;;�/4���ۚ�W��|���Yvr���8��D��ȸ�=k�O6�r��3��\�Ы0:����)e=vM]l��>^!d�=0�������]5�5�7���w|i�I�PÓ�v��|�0��Y�5�_/{F��K;��(�ս�{�4*���ҶW��w%��m,�K�Su"M�L�i�=!_W���|��?waz4�]u*u����O��.�՛}ז�nSF��ŧݻ'�7�Ŭܑ��*�q:�"�R}��������>]`X�dٷ�M�*!�m�z�)���Ϥ�
k�H�2���G0�=���;�K�(����9!��c��nuǷ��i��1L�,鈙�����[���*�N�Ck�8�;wE�J�Pkt]953\�x��0�:��8�S�]m�iM�vѼ��9��>u/�?b@9���<!�rV���3��j��$}��� ������	��d��z,��<�z[�v����s���]�>�a'CQ��kR������[�o%�x��9.Wt��~�����:���I�T���gu����(��\Tc�|ú�>";4��щf�}���)�����}{��.ya� �Z��z1��\7p����\~�J���Mm��'�R�P�֢�",�ӶbЭ�0��i��Pa�[VZ[�!9]��+y�LܖC�X� ʄ�D����s�+*�`vn������|
����9w���eu\���@��m���և*eI�4��t���l�#�_H�<v�(R][5n�A��EWj�TOea��r��o;�E}r�·p��tfз�\����O�؄����#o�n�ET�(ۺ�X#�$��W30��]m� ۃ�]Z�9�a�=~9X�б���.�[ ��u,�@y`�p�4U�П3�p����8.T�]v���ir57�,g@�{�����ރ�Hm�/U�it� ]b۪����rRܡ�=��
h��i�8��K�,�Q�ky���|�J]��{�k�����l�����°w+�Ua�g�6_��J�N	z��8\(f�.�aeʙ�^c=P+�[�f�4 ��(
��r��j
t-g֠%�{7i�-�כ҃���6��gy̔���9�r�[����{���e����1F��7X|~	��g¹��P����x�e����Y}��h�Bo��)�Uu-�d���UKS�Z��
�݋���,Q���U9z�z��y6��9*����ѱ�ęE�]��G$��mb�[jTs+�׽���oy�]��.Za�@/hz7��|�C�;�|�^�+᠗4��ȴ�ϲ�}@p�&,�T�t�+\�O�� �pXq�
,ԧ4���.�vVݫk_E.@�����#�v��F�/�-m����ը%0�&fWq�"7����^�.
�W_="C[�(s;M��ڈ���0�ܦ+o��v\v~����YT؏t��3���S�1<��!N<��۲���Bf���!/r�5�������nɁ�a�1JI�(o:Z]]�[F�Is1�:������Ǉ���p��m��}�^�_�1]zN&�H8٧ź�-!��YV1��{�Nuܪ{�����&m��!V�b�'�A������|�*��Q/�N�����^*r���탞{��v��N|E���q&G�Q��&/x�lʎ��R)-��Ҿ�
��X��l�Q0[�Ӝzh�Ǫ��P��f ��$��F0 n��Ήvhޞ��UƼ��M{7�L�����Y3Mo��ɗ�^�@CYnA�6�_'�w�oد��[�ؑ�i�)�p�=A��f��B/�d�������]�j�	�
FqO+P�iJ�[V.�.�~��W[��{��.w*D�e���*�Ma�����Ke��"��fp@c#%6�����P㧕�Gw�ll���Ⳓ��{oۥlze�y������6f93���R��O����;���>���N��y 5cӾѧQ=���b���采:��a���]\ZJ�2�])p�̠*Y\=f&"�9A�M{Q�)�=�����\y�dEM�;�(�s&�V�y3Ժ�ME}��Z��C���Vg3��^�肫|�l-a�ª��ӊ����	ÁPUb�V�HJ
��-
��ʻ��O�\4�c����,��1R_1�^���֘÷��qP���w+��u�3�����jvʆ>4�2�!�
e[��ɦ��%7HR��{�Os�̃y:�%0/"��-p	�`{��a�}ӈ����������"qo��[�{SX	s���5v���&���X�:ߎ^�T�&#����k>�3������d�XY�ܻ�
�Z�hS��trB��5�L�F��۔|�\7�Üی�u|D?��P<\9���ʾ�M{����1w��Vlq
1��wƯo�3h��q#�B�ۇJ㷭�]�9��~�9�oك���
�t(�D�
��DVЩ��x�3�`���.E6�KVT�3��p͊��P�9՝M�1+�M��Y�sy�{�k�D��;���L�m�*���5���)�5�Y����?;v���N�*�^�n������?���t���������N�d�kMG�Y��S�+nU�[���nt�;�sc�gP�eW��t�M��	��w��&��z�8V+Wa>�.�րK|g�O˳�{�Kx����嫦Fq��m�ʵb���G�-NH��k�q�o۟m擬ѱ���[B�m$��ۃ��m�]+
�Z���w���)C�o5��;i=��}m'; C���(�&��l=�� �ި��_Yv���O�Pe�d�z����]].���WǪ:mb2�2�uN- �d\��ۮ9�wHWG��Ǘ��;���)�2��#՗�q����ޕ���eHZI�뾙�.��z�Kl�/v�^���nK��nL�r���h���\y�M]ǻ����Ų�]Ya�)�-���r]�)��8���G[
g ��k��h8Z��T�iRW���~�ǂΎ�}�T��Z��Vn���9�j��}
�׾��[wz�s(��X����z�!%�CC�T��B��r��U�6W�w;�����-Ӏx� ��'b���3Y�d�f��2!A]�v���/M�	�&Gs%�3��Q�$]ø7�s}��&����Æ�k-�}F�2v�6��>f3�B�����Hdξ\�3���ۘ�G�J������;(��f�uL_FN�w�(6O\}� ����n��ܟ[�&�;�%R�?"+B�0<)�h�8r,Z!�q�SR4J�ǂ���6�ٺ�)p+�vw���,Z�M��5v�J9��K�ҧ��5�\�b�҃
�ں����&[�ɔ�}#�ڸa��_i�e��G=fr�Fѽ]�䝼OM��C�����{m�L��/C�\eE�������}DY�)�Ư�s�kf�D�{!�Ѭ����JI��͑Y�.�jj��� ���}K#��`��˩��𲲄v�|QC�b�7ܻ��>¯+J	CN䙈K������B�>ו�|y��p
��L��o)Rݾ̻r�=���q��T���_M�ֆ��2^�R�.���&��أ�����avU=he�Hm�GjڔZv(��`Sp�V���5Ҳ ' N��4P
2�9\�T���ѕ�����3o��7.V���H�.���M�;f�{��yYI��n3��/[�:���)a�Z9 �n&��*����i�D:����9;�W�}��
�T^V�`WV:'
���	��!$�v8P�جg�����}���%���w;z��0�l�ض�?��L\9Op�����K��0�+h�)z�Θ����#}��"j辰s��q�o٣�6�{X9A��t���v�ζcC�#:p';Qa'zl��ʛ���t8=��0��%�AMv왋5�.e#h�ǲ��m<�����~=�g8W�BL�T�H��t����&!�x�]K����������YZ�Eފn���1j������L��{8�X���*޲�4Ă�ux,jT���-�0���s�{��TP�����yH{����C�<,�>�M/��j<�N☩b����.()C��,��ׇ�^t4�#�Ќ�wEӅ���<2$����xF��c��Zh�.�R�%�%� l�!F�g�����/�یtYj�Vr��C}9g��ɦ:7��d0����e&�T%���I���G}�nZQ�:��k�+S,���<���v+\�yM�_uE��J7TI#\A*oR���ҧR̗�!p�^p6W�ev��|)��.�G�Q"�ً������ �:T�Uk�#���v�o=r��+� Vh�\���ˇ���螋ӑ�kF�ʼ����B�lFs��X&�
���
9D�$���y��N��l����,�r<�ܝ���Ẃ���t,`�Ȱ�>h�YK]�:�4>[�
��q؈���ɷb�:��������T�z��I5T������%��> ��
�Ե�wҍ]��p�g'd�)̨���9G�ˤk,CXhZ�O�#�j�\����%#hrr�w&
s�vոhj�#�ھG8f�$�2�:�$�m.�z�J=�b�
�7D��Fj!o�W����[;�u���Z�������k��nz�nY�z��rWu0�iB�f{�L]i��^�{;�� =b
<6_��$��/O<�s�v8���o%��laumO. 2�J�5o�3��X�cJK�$��zS\���T��ڔ�jǨY4^:ǖ�]�1d�j��3��*����F��9Mb�U=9xH�é܅��?��bB�.W����M^b\M`�SKܭ;S�t�Dr	��6(k�/�xu���-��չ�$�g%�2��w�\�Z��L9��I�x��T	��<7�s�Zv+R#8L��ovӫ�Yln��z����iQ'6љ2\2.�-q;��eS��Z칌�,�E��lY�v�'��
�ŉz�Z{�Vw"����\��s���Q?�QALZ4h(��h�b�hխ���Z6�Q���lm(+j�M��k��L[6��`�4kLMUTb ��m���[8t4�A��@��Y�*�����*��նt�%QT�ŭ͵P�QT�`#mDi�Al�Z�bh�ggk%�PQQ[�6��Ɗ)��ɭ��:)
C�A�֚*�Ŗ�b�Z�֣f")�Z�d֌���ئm��
��ضڱ�Lj���b��I�tTZtMcX1TZvl�$VэS��"&(�����*j&Ū4�䈪�-bb�����d�E�Q�f����)�Mj-�UV�U[64�6�M��"��mAUL�A����i'E��6l`���jq�(���i��0D�"(	��;UF�E�b�"4X�
�uZ�UQCMPF�AEb�ESD����Z֋h�J�m��M}C��wu�翗|[���a�='.��z4�
/��i�([��=)sr��x�p��3����o�ȏ���Y[{-b;*��^z^e��
�?�	�҂�{�ʁӕ`�/-Z�i�]�C���e��ףAԶ�$�:��zjX��s�Џ�y:u���4���t9�7T����a��w6�����Uja�+qP�;�Hi͆�4��J�/�a��uT!�]�ZC�m�{w<ŭ��r��~Q�'�MJw9O7u������N�Rp�h���NG�kv�|ٛ.�L8퇓����(̺W�N��N˥��o;J`��]���6Ҭ��X71���
Y�y!Uӥ1���e(V]4D�Rn�/)���-��JY�g��7�o�[�Tt^UAX��l�ҽ��&v���O'�i.�蝷^I�-h(x��yn��2�ߥ0�N1gwV�L��/`��K��٭�:���55���QM�ܬ�rE�廸��X���g\x����q��׊|�7}����ܽ�%���۹�������nY�N�+�m�V�s\#��;�1CW4�됬ϲj���5���}�y6�;�\��a�� |����,�w^�s�FZW�]
�33��j�+�i��T�5#7ű�L<'ʰ�y�9��b�]��m���f)+�nz�P(��ω}�}R�1=�!KI�b���E=0zFUfp���_?o�o�!AF����\�\�{�dڻyP�0^�uuG�F��Ns�̖<N�Qt:(�h9^��r־����7- m�q�ِ��C�YN�Uw�U^}eӑ܆��r�d�����ƽ1��Ҭ�pw�H���(���I�7�%��1�����#��2U��M\�l��������l�����m7[�:��2�zc����y�^�-��{�`OKW���%�=�{�w ������Tv����Ήq��ƨ}ݴ�Z�����J鋬�~݇U���F,>���9�����坘w%C��<:�v_`�s�vc�u��~��sg}���c_����#����i΂�zh�G8��;�]b�F����x�#◂_`3t�������_)��j�3k�@��X݀�b���t�V��5��w����/5J�Z�ݏ���Ѯ��Ǻ�ո����&,��Zsx�+��'�-Íz,�5��h�g}^���n(�F�	�X�Ki0qy��	䥮C6�	bQ[�\��8�Y�o�ۮ�̧��U�N�cB��Z.ݨ�ƽf����'�߭��=v�^�t�"�[�ͥ��<��Z�P��5�*���c���Jc��K~-���+x�`X��xо�-���`��gU�Λa>����__`��zT���)��y��pYy�R��j*;b�jv)�ʡ���e��Λy�v�sˈm=Y�o�("��\���~Y���?��~�Փ+7#��kGL$�ߠ&���Y���4��ǥQ:���)I����F4&Y�n�Z·��������)>lVvV���c�r��[�w��v��ҥ�}uRy��7{Ӱ�6��VWDf�oc5{M���:�F���)2_G��@��������[Ry��c��U�n��j���fUNq;��r�q�B5	�hN�fSǺ����R�7/=]���Z^�R�"6QN���d�+Uv�{������~�ud�U׳�f$qڴ��ϑx�f�]g���{�o^_�����I��bs�`���#�*xd=g\<ss¬��r��7DV�M��f�����@�I,��ν��1-�O˕l�E7L�,VNä�t���q^�>�ڤ�4]��@�[����}�̽}4�Õ��Ey����+ ơ��������!jf
��N�r8���|�P�BNEz��_��OW���{A̹���ו.��3+���7꫽ỳ1�Mzq��A8L/�t��u��W] ]�YO�J�NN��(n�m2���Ә�*��)߻�����,ka�Z{O%�ȶQ\!ýuO	���B~N���"�s���>T�{�S���ry������̘�m�r}�w�Uhq��n����mV�by{�=]T���׫-���W�1n������M
����������v��.�=�B��GUΑʔ�Rj,m���U�˄�[���*yz�(�ٗ�u3���*�ͽ잪}���q-�{�4+�S���B-��u�z�{F�����*J{"u=";w���{���!�%�OfM�����$�ʅ0�q/I|10���A��g��V�vNԻ�0���3�-�o[?M��+�	�&� \���OU�:3��qnC��VtO@k;��ٴ�{ç�N�E�����.�m��>.6y���X����=���Y�R&L����ع�׮�f��S����#s��|þ;�4��������o{&��O2�s�����~��AʷC��M���wh�C��� o�&�d����.�s�����Bp��W��VE���tcU�+�FiƗ|�>���[����N�.al:h'��b:��i�c�|��7�ϟy��8ot�s��FWw�P�����#���>kUX�6�N�^�p�qڃ�jڸU'!���zm�Pt�ᤕn�s� �F��s���)n9��@$���D�X�ӭ򛚧u�ó��hɄ��+�:��j�YT�_n��q;�Q��r�����I��<>'zi�����Nͪؼ���:16����;Sh5u��k�V������4����|�z�k�)��2�y*�������#}CÕ��&�*�y��=�<���	+�X�oՙtt�������!t:n]���R�}��ڱ^,���0^�G��/�-�Y�:3���*�� ����v�y�\�+��3�ם9/�VЦ�h��k��{,.�������V�bN�U��!���s��U7��\��e�օCǙ~kv��ۍ�4�e
ZK�:�_rT෡Tӂ���S��q]�����W|��Ɵnz��W��_Qx��n�-���żf���pU�|_�Z�AMׇ5sG@����F�u�Yt�%�h���O�"TLN���зXiƫ�B,�
�wK:f��t�L��$Xe�F��	l��v�6�V�u��T��ҝҙնy=O�G+{;�ޜ�ނ]y�y]a��?{�u4����;]��8ƄȻ�+p��y��w�.t��L��並z�$���|{"��K�{=�R�k�Dl䅷�ʺ�<�.��.j7/�M����p���9O=L.���O9�뀝m�7[�ΜjJ�Y��y�����d�w](��wY��4��ڮ@%M���b��JX��x�ѻni��#-u�m,�xN/�{�0m&�ov ��KǠu<��4��[��;��86��{��4�/|4���U4Y�h	{J�5�Ȃޭ�+>����b�����/�c5h;�D��g�}lt�}��T�:�Dp�ucݙz1,�]��?&��y
�:��Z�gO�m�݇Nj�p�t�=2�B�/@}�뜨�NCb񻦨=����[ys׻|B��Y�깷��y�_s}����l&�W8��wF��-Tlc:m��t}hz.}�����_O'i�?Gv�+��}�-�N:ӷ�SJ��0�1M�Χ��讖[�T�����k��v�N�>�1n�g��(�噔�Y�<�N�Q��X��+�T\m�Qs�,)׉�d�A���k�${+ks�m�o,�W��ݭ�1X���N�����uY�u6��FwS��m�~��7s�	������l\�n��9.��s:�n>8cb��r�����;B���|�o.��m㨁#�,�;=z�Z���`�q��+z���ӎ���飅J{3*m���=�� ���)-�$N����X�]@�"��{�Y:v؅|�Q��Ҧ�5I�o�9A�&��ĎU�<zyb��*�@Ka��N�ٱ������'��!z�cܧ�����'��G��^�ޱ1�^���o�	�T��}�Ng<��w(�x'����S���HYo��V�s�T��ؓ̇���-�'���3O�j�5�C�M�;��*�d�/lY��B�t�gR������qK�v��|���S�v�]sǭV�pV�6kݗ�r]���c����A8�B�G���P��/>��s3 �H�x�{wc�p���_u��,	�l:K�^����k�F����\���k^�sMXr��p۷�5���l��Nu�N�\�r2e�{����/)mC�ڨ̎��ڰ�EBp�)���°�{�:�J~܉�Q�3�޿�uw�0n�f�5�Ɯ�,	�x���:Ez�V�]�d��k�.ڶ7��'��s�nߧ۾��A,jGeZ�]�Ⱆ���H�h� �dߦ_le9����;^�g�+r{;a �x��I���ʲ���rJ�/\��[Ԯ�'����t��B��U�c
�G�����xa���W���b���suK�&���- �/�h�Ǚw�$w�e��|�bg�����Ij��>�]C�k�h�Ŗ��w�+]zn[�V�͞��8��Wi�݋�{1�zaw,��W��Oܪ����e��E��H��W)�mJ��9�!'W|�m6�ry�K*���	ۣ����Y��0�4��U�Wf�<����tS���bi�K[�%a��p�E�mY��H��4c�b���+\~2&�3�8����Ϳ'�J��8g5�9P�{)��ƺ%L��F�s���B��z�'ɻ�)(|鉯�#d��ީ��K:��A(3���'s�܇��ݺ܄���ڬk��c�E��,��T��W���Cb`jtc��L�{X�e����w�)�R��n_y�^vK����.��C�C����L�RSY�ˊ�<Yƀ�y�Q�ۃ�k�s��n�o��:����4y�Y`&��=�N瞬��Gs�u��7��MmK[s���TC��,�т�0��m{����m�X�Y۩�M�T��GS좦2�E��^�uh*���4v]�2�-�`�[�z�Ó��
�h.l���J�WY�[��Y�3l�j>G]l�A:�|m瞵d��6g�
�[�<3���=��T���/��{�ɭ�ie��zƁ�ND�����w�:���elBp�2����i7Qq]�>�H̦���%b��w9K7]Tn�&lؚ9l,�4ʮ]�p�UY1C�ŷRұn���N��KSN���=��1���Wv�%�����ћ�'ښ��X��Z�@���Ϋ*Z�4GU��[�p�vx��������_�ls�{8TBƃv�k{��w�(.����ê޷I�s{�v��)�����J/Ӷ�'YkZ�䶽��yFP���矺�[a�੘;b}MLV�Evkw���Wɬ^�i��kv%��M@����.��tr�V�Õ�'(䰢�A�ƣps9�J�1D��=���z�j�����e7�F�-6޺�T�_nΙڗ
�c2�]��w���ѻ���j�z��(r�ѱ�a:�\�c�Z�]^Nf�c�1�WXF��z�#[���g s������gm^L"b����0?l�=�>T+�=
>��ۀ_KA8w��xS[>woEy�R�oU�[M�h��P��̉3N0Ƕ��fN�~��w�L4�18�ī;���m$N��,�}�Ű��vl�jZq{�`�^�T��_iJ5��fu$U��VXU2��EC�ws���� V�p�2����,K�6滰�n8^i�A��y�w9�������^�r���x�p��j�y&��9��wk������>�������b^e�7�dw���0r��!ñ��;HVN�u��s�����*,D��:�5V��fu�-`���x�O�:�coFS���jF��Vp�Y��3r"M�i���yCVt�fҔ3�"�*YڋJ�X4c�:=�.�3)�q�;�[��D��cyOlI]1�򑻫�siV����",�ܸ�#.�/��'p��K�R�rf�&a�.��A
Í����}w�j��JJԮ[}�&&���ndS:��
��q��W��^�Eb��Î�Pn��9Y�]f�ũƜ;A�%�[��弽_v�yG���Y��{_9V�#m�+���{hXE��w}�Pf��Z!v>V�u�x��Y��u�)�ۇ�V�V�AR�1�u*j��ݼVxq�8����+7w�d+��)͵�8w75��R�Ѝ�e�_!*R��ޟ�I|�f��.�]�"hA��-�6w�0]^iKn���-r�D�w�t,il��+�>�Ik�ҹ���Ug`�"�-]],,�X�y5wu=㎂��� �%��&��w�di�pւ�rR鐄f����vos��7��(�o���%�m	�NR�%F<�������1��ׇsz�B.00ʑ��k��+9N�k#v��G���ZFV��0og_7���k�1��4`��֜T�LL�Ͷ�jp��v��Ci*3�%��j��۾"�Ҡ����Y�gEL��PX94�Z� Jc[��=��/(;"^���{��սǴ�y���e��4ū!�P��߁�ށEL�j���3M+c���C�k/n�e��/�|�_fi��Fn����].���5r�O\4�/	�(�;��ca��re(�ݺ�T�<q��<ߴ��������zh�*�3�Tj�M=��a�A���e&m��&)6�m�q館���)57�0p$���\I�8�oj�g�M�4�����;�e=��q%^�q�`�c`�ܽ��W�$��:������HM��f���G��4r�A�_��݇�H���N߈0�)Ug@�h��V	�m]z��x�TGx'ny��(^WuXx�M4�M��ط��&9���פXÛ���_:����v�2�j��.6���k���& V���sE���ڹSԍ�uL���-��0�
�՝�
d{�ð�maT̓}K}�����w�q�����F��֤��cQ���՜EZ�U�"��F֧l�kv5Q5��i������M��$֊����PL5la� �Z���cEL[�f���lli���4�jq�S4QTAV���b&��6�DMDΰE2D��Q5LMF�EQ�U�M�QT�uUERQQ�EkTV�clE�Qƍ�%U3PTE�E�:��LS�Ѣ(�4i*��I�kZ��*6�ĕVڂ�)���
��Fء� +X��c&�5TTPD[f(��""�IT�0�ْ���d�����8��)�-�Lŭ5Fن֢k`)�	i5��l�:" �+X�M&��Ei�Ӣ�`����b��j*���54TMTm��(��Ѣ֝)�ѪMb���J�6�Pj��"��EE4li���* ���X��m�Q�TF؈("j���Y���u�7Uֹ��=�PD�i��/0�����=�Nx�j�F���"�#���K�5ޫ)ElV���,�5f�o'�$>���>�of�'�2��3���CFR���ӑ2筷�z���_�N�]uŧ��w����MOy�\EF��jo%�?G��uu��\�Q��^�����$׊I���}�Cp�T�<�L�/l��(<L��}W�<{�7;��Y���{ES�2k��c��8�m�qչP���+ �P�����'�I[����NHQ`���q��Vv汲���M��4�~�6�
�'p]gC�G6���&b�>/����Ii6�Q�NEy���;��#��-��QNT�����]�^�ow�{o�+�OmG	�N������N�X�4��g.�i�����p��1�[sJ}X�N\��ǩ�V�(o�������L��=�wKK�{�Z�ˉ���|E��k��m�O*�6!��ӱz�j7d��s�i�qo���D���ܛB��n�C(8�����b��x�ך�x�اP\ �y9���Օ��C*|���������<��3��m������}��m�����F�����e�5�qtCOUtJ�8�8���l��g��|�倫Ũ�iٙE`�jb����j.w�DvL]����3Y"ȶ�%,��G��"����f�w�OFΥ*����D���T�F%=8Ԫ
t����qK-�l\�螨9.��&I-��t��:��z
������/6�;�	��=:�u�#�B	g�겍n�un%��ڨ��4�M�5��)V���Kڈ}g�r8M�-�O+21mt)�LFA��T���_ObO2�zuVm�9�,R͊������o'���!�рԆ������jG�=����	�o����qՋ/i��;�󾪈OC���0yug�:;o^;P��j*��{L��L������ߓu�~�n��B�+5y��Jچf�F��s�^����-v暰�m�s�P��sP�XPԯk�_9ǻ�x�T���]�hV)�Y+������(]�4��Ie3�{#,��/|2���/�lAX�Jfv	i���
gy��W,_a!p�Zǟ��Vfkt�P<�:E�.:L�2�L�x%,��s� ��8
4ג���aM`*������[�a%�wն\��%�ep�W���m����;��"�8Y�y��C����-�F�V'r���nN�Q�>��W���8���ju�=5����	(�d(����nK��ܔ��etve;�z+S�j�����*]�;��Wl�%5���~n2c�u�U��?\|��t�k�+jJ��������/S��T~�K��������μ��6��͙ʘqs<�:W:��6ڋ�s	:��M
���e^'wuf[��SJ�J���Νjz�eu�j��2;5�~�L'9��e��܈��oҰ�b�J5�t���"�nw��}叮���.c)��y�!KS���"�=W��w,����.�(U�-�>j�����s���XO]S���y��E�/��n�.7��s�85��ꦉL:������b0�j{͚��M�T�>���9��qJk��,�����iG�^��i6"`7�n�f�ݍ' �%yU�ָ�h����y����n��6dH�]�x���^V-[�|�K�Y��v�R��#oR�R�K��f�i��ۯR�s��˔���g6��H�@��U}���������E�� ��۶��ZN��j��ԥ���^�zOg�rʸv�[��캇"?�G��"��z"���B<Ǽ�Y�����f�ܭ�[S�.=W�O�;��Q�9;���������'ӎ�<��!�����<����ܟ#�p�y�߁J�'�x���#�r�΢���}g{�eƏ�C��}��=K�s�G�OǜZW��w���~���!z�����`Oܷ|>K䟠=�/��^����U}�U1_<Ύ�:���6n��o�q���R��\�4/���z�/�0���}�\H��:~���>��ï����w������a|��=�=�����ݿ�m"���������R��|��N����/>���̯�}<�ѡx�is�����_o�?0=�{�9���I����=��E�t��x�#���bW(Y�	�ﻱ����zuR<G��9��)_}�(<��y}�4=K��߿e}��x]}������댏�y��?2{/��DY����X�1��a�s?pw�V��X�w��쿠������<�����y/pR���u���ӿx��~u�ߊ�{��_%|�����F��{�0{�����őn�>]��#�+��"=�8�}��;���\!�s/�W���^��O�p{ |�e�4/��������:��?���^ 9:���|�g��|��W���vkww(��U}����d�G��y>�� ~8�~K�/ϼ/P{/�W�����<��9��~����|��Ye���d:��{�T��u��~��sa��WШD��Zl�����c.�;az5:��Ѵ*6���zr}gmazJ-㻏�<�7���B'R�[�������f����]���m4�#F\��uaNz��c��<D81w*9݋��;z��h.�n��l������)��z�ys���������y�����_���_���8=��o�q/pR��/P{/�y�� ��rq��̯��ߜ��=��7�Ϧf�pL�^�)Ə{��^}��=\��_�z���?��z�N0=G�}�N3�!G�AJ�|��_ ������gG��>Q3�T�rg��w��鵝�X��rz����#��_!��_}�}����@?�u:^��N2�G�{�x����9>`�
W��<����N�0w���^o9�Ͱ���G�������)��O��p{w�M���Ͻ\!�?o��O=���#�}8���|���:_�vC���rq�%��!�A�}J���V��AF5������z��z�!�޸�|��?p���>}���#�<ϰ�y�|�����{���į������	�6{�K� E��}W$��h}=h�߽�F�{A��W�>Gǜ�G�_m��s)����/�`����O����ܾ�̿}���!�7��|���{�_�C���<]1�
��P�\n���~3�|EP_~�~�4�AI@u��=pa{���s��_'�8?K��S���<��z���0�H���?]�������^��G��x}Y{7#��:��N=�!�{�mD�{�E������-/Q�������#ܾG�r{h_'�xN���}�y!��hb#}�O�{�=P��J3
�}��f9V��.��=��"#�jc�zǽ�=�s�>�Լ����)_ �ϼ.�#��I��_�_e��>?2=��|~���������=c�7�gd����W�p���N�13F���������{�X��|��@{�M���Ǿ�~��~s��|�.���M/W0|ǽ����H��h���'�a��<�ksn��5�j�%���[�.��r(�ǐKAk����a8���d��e�=I=7��8f��ٮ�.w����������/��p��0�y�dG��e�=G�=����].���RK;���lt���|��Y�gW���"���>~�_.%�^��y�?�߸�WF��p{'�����|���ܔK�
������~<������}���!B"&��/��7d�Z�W].T���.�ߘ�>O�~Js�|!��/�};�eti>u��R��w���	��!�F��p�?a��~�y���W��_�t>Z~w3�������G��^����d�C�y����Ne�S�8�=��{��=p�S̾����d����R�>>u��F���x���A��q���Iٺ�����Kߟ?|W�};���쏑��Z�P�:`c��'�<��s���_a�������{�����_�{'/�p{ 1U�a|�z��~������]���}�������Oe�~���xC�{���޻�S���W����q��w3��|��4|�'�y#�C�����>�YϦ����7v�8�Ո/��?����_�~���>�|���>���K���}��_���������3Ծ�'�W���AB��ߟ׏n>�j�8����n�[_P���({�<�������`�c��#��{/w�=��a�_��x_d?C����K�C�������猧C�=�[x�E�7��8�76��6~�]��`�}���(^>o`�^�Hw�'��{�=���>���K�{/����p���w�=��� s��t��z
�4��qO�k�:�� �{D{C���%�98������w�<����{�i=�˨<����~}����x=���|������^���}��O��h��,���yǤ{ޡFT��~�����'	���h�?��:>`�~B�i=��N���_%����4�������~C�˧�Ӯ��g�)��c�c��Om�)�&�VI��˽�\+�xq �1	��@A��5��7/yV������`���daT9�l0o(O�����SDN�79d�8;"خG{�FXU���mW^pz���h�{�$���l�&�bՐ�7��z#35-�V�Ž�4{�{�ϣ�?��O{��q+�s��A@��|�C�
���/�����������G��&#��|0G��L�1G��<��|�U�V��s�5]���B���c���X���������{���<�������A@�w� ���/�0���`z=ȣ��}�!�X�S�����U���}��%�s	���$=���=���/�8=��?@}����_������>�̾��|��>� ����K�A�����!Czr�t�}����wм��u'{z��y���>�}��+������e|���|��?H}���PSϾ��u/�|�)a�:H�x8�?WL1�^�w}����_`�K�C݇�z���r|��/��}���/ps�����'']p�>����d�WϷ�%�
�rPy�)�{�=��,�?Z4S����,Z��U��E�����#������ǌ>@~����)܇���e�/�~���=��;;�!t�>=y��!��~p{>b �ڜm��5
`g�z>|6���2�:�i>���~Ȝ�|𻜯���i_`>q��a�uA�_%:�'����{�!�>K쟻�d�"$����톗�d��~������~��_O=��%�O�����K�~��+Ľ�s�>����}���y+��u�0�#�u%�O!��ݮ����ٕ�ջ#{>��G�G�D�C��rs��H�>~ϰ�:S�z��%�/�}���������W�y:���q�rw��u/1���>�������wф\��}��I}�#������({�D珸��`�ϟ��O��p{�����p���9����/w�z�� ��<�{��z��:���q/2�<�����]o�vrw\���w��1TJ�]e��v�p�Α6)�0�&S۲%o�-NzK\9��g�wJ�����xd�Qk�\[�X�M�.$�R��uEa�cFF9���_LZ��xvS ��Ʃ~���X��c�j��\���DG�����xn������^c�8��/����N���%�
^{�?A�Ə�?p��{'<y��sry����G�y����{�p�W���z#�{C� �m������v�c�9�r�=#��菡xzG�A
}�%�t�#����/�����}p�%�4y�#���ǜ�{��z1�����O����خ8�~5�4�����5�[����{�>�y�{�2rc�C�'͓�iI�A���|���^��9���)��rw��>}p�=�����{>��1�f���؄��}��{�~����+̞��p�y#��y��ι����]'�N͓�iAI�a?A�>O<n%#�q���+��w胴/E>�P��2��_Nu��G��r������)�;��߼��/��8=��ܽC�H����~��/�8] pw� ����㰟��_c��{�C�Ǧo��cw�ٵ��:3��AC�~ZO���)������_{��=��z�����_���ג����{����|�<H��~p�
��y��@���ƾ��18~ǵ�+gW}�cӃ+ԝ�0wi^�䟥��S���|���:��e�G�}��������_c俤�����y|�����F�k��g��b�������;�:
׭�:ӡ�q�����e�?9��|��xN���N�ϐ�n��|��^|>K̟�>����"ǽ� u}��W�ru^T:H]Iw�=A�>��J���ѡ~��á�:_�|��{�\�2>@~��ui���a�R�g}��#��9����{�[W��G^>�w�uiϕ�=�� 뼔K�
}�����������ܺ4/���t���h|����. |������?e�O߰�� 玾�;�>�V��	���0�ȟT;,�;W��p!�_u�NT��/�;�7�o��s�P�,��"�3;���a�����
J�֊���:�<�8�f:x�^�!����r�����@
�ɛF�.%G��;"7�����53�:��)\�x�����G��U�2�B�.��ti?��pw�<G'~�s/�R�{�Py/PSϾp&��}�����ןx]}�������>K�?n����{�z�8 �>�z-VwY��!����=����|��}�쮝ï8=������e�
C�}�:��N��~�%R��߿dx����.����O�{�DJug>��>�]B�Y��>��_/���e�S��}�����C�|��+����=���p{+���\��h}���|���=�!ԽK�ﲐ�zDD}�O������{��}�}#${�{�C��^c������'�!��}�%�Oa�9��2�}>~�_�y�g��+�|���h=뇨����1���N��MO�1���(���g�|��{����!��=\C�_#H�~��i�W�i����7pq/�R��\/�=��+����>��ǜ>�7��'��p�?|k�j�};;x��=�<?c�|��X}9��:��?�|��^�?�?��z�N0=G�}�xϒ�N�`�
W����AK��\�����EnC���{�r��J:����������q̏�]��|����K�?�%�x_az�8���!��������4�QĽƍ+�c��<����	��B'��fGW�9�S���P�=����|����{�
i}������'�y��>]H�=�p���w/�=���#�}>�!(?N�����;���bTTLf
;d����\`���"�}E<����N0y/q�>w���_:����)��O�}���#�}��{���z���z���{��8��9����߾��{u�.��+'�!���#����l�pu/���G�>G?2w%{�8���e9;��_%������'����ܾ�̿}�����7�=�_#�~O�O��e�����eؽ���;�UL�qU�!cӫZami���ny�i�lZ��d��ږ%��01A�sR�����~���%(�����'Y�����Iw�;���QU�p|Q�g8 �*<�ۊ���9w:\P�3��(���W�4LW	��Y��ϾϾΝR����9���#��d�� D{�DiAI�`;��}�B����N�䏓����}����|���:<��GG��{�=�������弫S�SԷ���p�y�E��c�B,{�����}���x�y�/�����秃#����'v��{��G�h���L���G�18n_@�	����qY=آ��;���c����=�� }|���y���/y���}���>�4���M/�����>���r|��/�����|�ǿ���E��<�ٱ��㶥}�#yG��c��{�>����Oe|�{��_!���xM�z��O}�O`�/!��~#�<�}�th^?o$����s�_%�/�1��|����Z�b9�K���=���1�!�!������O߷��4��<��Oe|�^����(N|����^����xC�>���_a�<����>߿vs��m��֌v~6���H.��!��#���ho#ߘe8>g��^e���xC��/�>��ǲ�4��8=������� �<�%���'�x��}�~��Le*�^����5�U����G�{�Gd��}���̴=_`>q��a�uC�Ne�S��:�e�$��C����?w����I��{+���p{/��7Ө5��5��G}jE��~����1z>��ǍR�:���U�^C��.��������<�<`�W��s�'2y#��G�}��~������|��?|�����Ĉ2�}���q��f�" �y�����S�θ��_��z<��;��y�޻�^%����Ŀ��>��P�<�%z���H�����PEgR�{�'!|��ͮS�9O}�!c��q��p{ǜ�0�`�ߜ��iN~������\��K�׾���@uV��}��2�g���'�W����< W������~^Z����8:QB#�P=Ԗ��*�p�1F,p��O"�����4j�dO�����Cn��V�mv�p��e��L���t�o� ��%�7��*��{@������_X�z;GsW,λ�Cæ��Z���z0"�7��˴����Z7'{|�W���4�z_�6�R��awG�|�ڂ��昝Y�Y\ts�@��Tq�	����
u��a���NWܞ�H��&�I^�βh�$���j4{��s5'���;�@8gY���y�%�u0���##{��Һ}�&�N��Υ��0�,&����*�鳲ȹ�=�&leM�;]k�B;fi�˵�����)�-ոJ>�p/��Gݺ�{�	���Ik+�!���u�h'Y63�vB�h-�{���b[x�V�p���Y��0S���1����p�qUL�R��]�h����e�K`�)�CN�'�t�b��SlIٯ�g��|Ḥ���b�ȁiac(���C�ʺgF�̖��fl�����y�˒��{C a�J��0�X'�nvt�>��
Ûa��mX�6�u`������X�,�#��%���{8w��~��Oވ�oi-(p�,���|ٺU:
�
�d3�n>���z�o<w9f����۞�%��*fY��j���\h��f|Պ��!gU��Q��kݡK��ؗZ<N�.t�����G�I�/-��K25r�i�me��U��ve!�J��^m��e�pBs�#9<�X�(j�z	�n[�L���잨q�����_��L��_�����fo�Y#ܝѵ�J�c0���<���<������ۺvrO)JU[������]�Hd��q�jR�uz�ׇ/hU���:���cEH�I�Hw ��j⚅	�pL�f��6s�ZJrn�+t���%�[�6��rV�Y����n\D��Y�^�*�|��wX7'>=�����l}����
b�\ >W����f�g���1�X�<��,�}�� y�ٳn^���n}����ɶ	o���jes4_e×�����͙�mv��lS�J��y/韂8�Dߢ�ݺ�2�a�A�U� �S��V�������ɯ�/xq����h�׬�Ճ�K㖤�i���t���6����}0]�T���vZ⠠�z
h҅BZ�۫�ݘ�a�6��L゛頧1�}�������|���G�[+�z__m��z6ڵ����Jiĺ�/%�kR�u� ��!S�ZuR&X�����}���Q�˭�N��:D\(W*���.kA�dHG�V߇Md�u���6���B�< �uzj�p�pG���!�M��0���OTz�����"�aBo3m�a��S��� [��L�CWw�nq}E�-|�ξ�����m�̻�+Mi�EN�f�d�k�c��q�]��}��&I*�"�h�h��h��lUS�����EPU4QT�E3DTQ�i��("u�*)�����������4�4h��*�M�E4�`������$�f�	��L[[I[�T�TURQE1QPIQ1A4R�4�RAQTT-T�5ULT�m����"J&	"&$���8ъ�*����RAEM%51$U-Fڢ��b�&����PQD4Pα�m&*
��jm�LEDDQ$Z�V�SRk1TI13Q4Mƪ"F�)*+m1�SDӣP�RTA�)"�j���h�� �(���[gD�N�֙���]:����mSQ0D��DU�J	����ML���4E�Ql䨶�ESlh"���h�lT�4�Ik:�V�����;������+m�v���X��z���{�'��x��'+�]���$�;��k:��*�� 뼝�D�"�s{�����Dc��W*�ƿ}D��"4G�Dl��"��G�"�_��N��\?�����ې_Rݫ���S�Kk�O���H&+�?�V�m��g�59���Y֞=�U]�M�s��������|p�XN�����B�41���4�oZ{�(�3ݭ�定�Ť���;��-�E�Ӣ�;��N.O�3O�v�C��B�Z:	�UJ�[�{V,�yZ��зq�v%��E�C��X�n����U'�Vי)R��w*��z���쮷Z>���:�p�.6|�����j�_N�%	㐧�y���x�f��>���뾫���t�8R>��]syw�����_M�&���y�5��m���yNjt�n��J~~w�^G�\�����qF��I�s�����[�SO�-���m�c��p]w�&�0��R}�d�����w�ki��؃��v����V����0���V{��,�&�	�	Y��Y��J��Bċj�1O�r��J��C�*՟�P5�}�AK5�z����\�_m.�1�ǖ8���1�ozQ�}�XUK����R�nK̷Go#��ewnwf�}���b�ԡj�8�VG�(x)1��ӸV-�udח�5N��n�ORP�������ޞ�4��wd�|2{�U�9-��X�ח�޿��C2�\6?W�kή�a��Z�bև<Ţ��u�}��W^g�y�)e�����g��o-��b�Y7�E�Nڤ�e�hU��r)f�}��oq�Լ�&U�j�Љ���`�Ss]*+�S:�Nk"5��5�K�Y�n�'���Ъ�Y�6��'(亂�O�A���Aj|S籁Q�	��Q�ĝ���;_���@��az���u��#�$&��qd��=�0c���q>�1�9�GD�ë�	}�~�����3+�΅O�'�$?v����˾ٯI�{�̗��X��~;:
wm�����Ү�,�nh��9[j<��w��A�s)֪���T>���D?D`~�K�;�Q�kΓ$,
C4YkP6�Fڕ������G�(.�1ل�	�K���1�8�k e��*8n�/Z�gVO��N+Fh�|_�&�Cuu�g-&���E76Dѽӽ�4�omT�R�=tl�EkJ4��)� Y����ϱ��I�R�@�TcT�1Z򸥝�>��^�Su�n��&(�f�{R��<�/l��!}�g2'����f��
k�e�05���/����_e��ᗎ��{=ׁ��2d�u�����gnk���Ḝ��k�~�`�ǳɮ�Ν��8B�v�y��m(�k8	I�P�(��dW�>n���su�szs3���H�].�m��w܀���Lrj��}�7I��L�]�\\b��o��?z�e�o�m)��J�)E�v:��Jƅ7�E�[���~my>H]�sl{���9VA9���+]EҘ���6T����ր�G�]���v�ɫ��v=�ꞓ&��KQ�~6꠬�qQ���_�S½��P�u�ǎk:�.Oq�����v�ӻ��A�a`�R�֡ڃ騛^yۣ{E�G��獤Ӷ^.�N��=i!�F��ց�J�����7�$����G)������oPZ,Q�����g�����t��z�9Ւ����3�X��j�cf��`}�d�?a�sƭ������;��u�GwB3�{ޏz"�������8>�Ԩ�N9�O�s��
����u�R�<�f����N����v�x�6�>	���г��Ѱ�h���v��z�rk��z�ܢ�2xs���o3(	��Ӝ�9�;��'R�����y���G�{�S7�υ�`$�4�<fN���vk��ٯ/���)�zm�b�a�Z'U�\�xz�H��o�<�S]*�����+)v����<��zI9��p�\���}���v�G|��I�`!:��O��iҪ�S���#�W�����:����;u^sp�Xچ��Ϧ�+U�0c�I�S��GOV���
���~sM\@r�����c��K'ø��{r>B�Yr4Y�|����鋬�q��^�@O�mXr����ؼn������Y���^c�ʷ;�ܠ1�۟���7]�n�/���N���3ұ���EV�vI�/��;��N�?C�=�����,��7c{����Ւ`]�нU=�O�%�gʫ�@�Q���k�B�b����)�%��|5c<���ʄ^˷k�]���y&����󻩼
��8�#��p�X9�+1g{Qf:+�����}�}U�|������$�O�b��2�w�VV:WY�����[ȼ����+��՘Ը=�e����_��Nu�-�=<���{��<��7�7��9�ͩ�B��9�S��~�>�%ͮ��<��Z���h��陥����Xv���s�q�q6ڋ��tS��Ч�1�,�o3ctK��6���]��Z��R��bC�%���l/N�PS������Ȧ�nl_v��t�l��T�p4�i���AӃ���	
�X���n������;�sZ�*�˝l�٘l���ak����\���:{�*޷�%p싹�y��e�wMwT����|�;�QcN�;��I��WS1� �'m:uUώ���4A>L�c������p����Nΰ��n���EU\XJ���&�q���Z��YW���;����Bp�.7ݤ{j�k'��i��nY�y?�S�:Ǘ��M�!�{v�Ě�d��(k�/ާ�E�[ŵ�,�
eȋ]�˽�#�^6.��[�;�#M�ƜŖ�0�x�N�E���d� f��y��j;:!���fv�s}�<\��U�qx�eE����#����m~t���D��ld�im��,s{Q��dSu�-�3	yX�۹u�� Jz�r�x�Р�w�Ol�o�����sMXr��u�q-��7��"�6�S��>�+u�ۄ�Κ	�U��1Lj�e%w�������U8oKsn���$�ٷ�=={`.����a�)������������ y뙥T�W�yF\�ge���qQ��^hd�t�
{�+����I�9��yxjz�e3ѽ��޵�EF�cQ�o��q��Nu�]�=�Qv
��Ĵ����Ҿ�z����ۍ��U�bևC�Z.ݨ�|k�xT�c3.U���5�~8�EҚ�qSx�������ж���tj�v�_\cf��r����uօ�5}������.u:��]�k{����5��j���ײ�m�t�m�%�ʅ�r�K��O�A��⣰$)j{�f�f.z�8�q���f��O*��!��S��o�S��v��1�{��l۞���Rp��^�sD& 4�>W�+u�l��qt:�(�a���+���@�={̷�c�v���e��U�ͮ�h3���n�h}�V9][��S[��J^�0ӂ)/߳�>���W����Ω���<�{�z^<60bPrU��GM&*�jh��Gf�#<�rei�Г�`3��ӛ`	����:tQ�--���oB�F!y���A�e��^6�"0�j|��\�Y�#��غ�P�mS�ʪ�\�GV�c1��y���Okw�t�ޫ��j����o��]�8�姲_+԰*���s��
}Z�W�S�o��Su��0�3�/.n�W8:�����Fұ9yh�˧��f�u�׳��������C6���Ķ�v��8����5
��uW��U��%��z�c�<���O�Ԓ7�_u��+m8��m�y�S��C����Q�2��y�1�Jw3f	���dp�8{�X�I�P�(�'!�y���h�J��z��H���i�F��Ν��?Ol�e;���w���p'�QP�-�6q�kU�T (���1a�\�2��U�wt����	bW��|��ɢ�����|n��i�P"�"5���T{pox�lW�l���ם޳�T�-����q�;]]pv���J:������z[�K��K��WfWSA�#z���M�I�����=���k%r�/�C��Q}!չSnWVe(���u���,h7k�JC�jqZ�M�y�Z͔�;�Yb�Ed����ano%A�K�:�\7��[k2zy�����k���ϧ�ot��}A`���TWf��QRq[Gfv����5����O��{��g�{U�e���k�����q�Q��g2��fZ�r*h\��:w��M=YM�1�%QW+1-έ|V�_�����-�rJ̢����������}m�Y֞7f���bnf���H[U�H�~;<Y�s�p�ZZ���޵���0��7*ї��F�j�p:tP_ZN&��<���c���:C%ɬ��\����-㊜oK�~N"0����r�԰���Ry�V��j̡ׅgEUd�&����z����2����c����8�!:ٕ�#+��Fv@)���Z�Q�Y*���Z�r�n�2���#[�E6�zk���k
�+-#ʕ���%�\ݫ�u0E�z���I���o�dO��K�D`�.GUŹ�l��WD3��5)��]^�y���xG��Q#��j�E�����dd�ʜ������G[�=�N\�U��3Y���m��fݺ�9�T��h�})����J��8i.��o��C]����z��5��6'"�{Nj�.�>�W}�4�:�}�����C�I�~���ݱ�[�	I���Bp�+͌bf�Ym���Ҭޮq��amfO���׮﹁8�MFU�n���N�_OU��a�aE��d���]by�\Tw��|�ߟJwo���`�x��z����o��7�f�|�sŢ��O�ޚ��+$*u)Ed����rն�ܵX�k�K�`�k��bևD<Ż��uT����VeCŖJ�޹�ۋ�Ci�7���yW�uw�M
���E,ݶ�ktK�)��r���l�.v(Vj�>4-��l�?l�Vΰ�\ƺ{ M>ܦ�^��s{]n��P��e!�lK��E�Pbu1]� �>��;	���x�{������M�e�/5�F�2ϳ��*_a�7��֮��i����P���ƋG�Я��eKL�Sv5�� d�.VNA˞�̬��}�fv���eR���w��͹Z��#��I�k=�ښI�0G��U��R%����l��]�o��_UU}\���im�B�}�ߍ����]A�U�uץ�M.��k.�N&{9S�I�콞˞�Wڛ�Ù����E�Ӣ�;Ж��種*�7��"��)��U�.
^k�����݈�;�Bp�vu��ݚ�C4�.yLԜ���[���}�_.�^y�*�sq��<.��<��$"�Zr_��e(�_!�B�u��7]س����Yަ�f[�sP�)���X���ܮ�C�<c@֧%���S|5�OU�����ۭ��v�����P����bjjC�j&�5+f�:�#j����w��+.�����=����^R���{P]S�V���5�n����԰y˞�ǆ=�����a��N42[�w�V-�tuϊ�˚C�pJ�)@�7��
W:i�N.{��o�y��ޡk�o�q{���X�Q�x���T��*|#���ۂ�+7'S���I�9M�+
:�v,o�R���oC� +�����\�#h�vt�$f]�v�2�)Cl���}��M��c/L9�Ƃ��o6Z)�ƭȖ��Ts��Y\L�ڥǫڏ\�Hu݊f<ªަ�g%�d�
�O}D��-����`����o�\wh'����*�+x��SgD��E�����"=@]���Z%4 �|�;]:�Om�6Ҭ"��.��)_
ܧ�{K
q#��������\���Q��JAtkWA���1�X+�.�	l/N��Ѿ��]xe��!G���p��L�z���{sT�m�&��g0����\Y�F�sb��+���lc$^�?H��	
�qP���-'�8�{)�X4R1m(�OL�s9��4(�m���w�Q���,-�]֊���q��o�^�����ɒ3w��D�g
/{*�;*����/q8�v�#�,PS�E��bt|s��՗Gwظ��8��Qn��*��	S�����N>������nam+�n��|0-+�Y��n���{;{w�<+Sɩ�.V9fv��C�B2�ÙSH��*�[����Z��xj~��	Q�Ժ>3���r��k;��GOe��1P����4-�S�ڊ׽&>H�/z�z�'�ґ���`n`��'s�y��4�}Q��2Ԭ`������2���;�CB/��M7\2���"��<���]Q�YC�'{�z*���/ݡ��<^q�-˦�uZ�[��~t�V*9ܼ˛dc@�����4 �o�6��)�S��z�7�9��"
����ݫ<�z�e��<��˖�ɼ^p�`ʦu�:��ƶ0>��n�L��ĭ�q0.�2�"0��
F���wFr�M��x�����5W�S'D�V�Q�bx3��uy�\5�=ݾ�v�MM�Ƴ�U|�,�2:מ�K=Ȣ4�Mi�v�x1��-��F���ޖ�̠���m
i���k&hhŻz±���}Bt�� L0q�j�hVϕ��j0$�c0�W[�-!��̱��"|��FN;�{2?h%��.#(Ê(f�.������@E�E�꺸ˮ�T�GZ�g���h_{�u�<��|B��pg��[o�ޟ�<V2�>/Ef��2Ν�&t"��2�T�
�;��&u�2��m�DlMjħYC�4�'��orp���R�QQ�j��q
�%�e�١�9%9��T�a�O"�d2��d�b�ش���a�؅>�1��9�����K��j�&7f����F�k�P�N��v
��ylw�c��T��FL	U�oO��a\���6��L5��ړ#ބ>�Z����ύ����3�v ��n"���t�������Z]]����u7s�'N�#V��#��T~��{�`)I����x�c�ͅI{��:�#'��Ѥk�y�ך��LZ�XB��<ylA�d���mH���d���4�������\��u�DwfэZf(&	�*����!�Ѫj�m�V�Y�b���X4ETTD��U����ŧN����b���(��b���b"jcZ����j**4��f+Z�:
�m�EZ�[S�m&��ѩ�(����&(�1�&(��QUS%PULLQ3Zu�QDASlm����S�$ES1D�T�h5UUPD�LQE[��"�j٬ѭL�Z��&"���	�b)��6�3:5E$M"����lTa��(�uXu� ��њh���&*)��"��S�Eb�ff-:��"*�4b���DTUKUcY�5�**(��("(�(b�ѣ1Tm����)`��)�� ����|�����}ʍ�+��H��W�0��u"�r��|�=���u�y�s��=��ߎ�ҭ�e�[��1��քt���>��>�����R�湵?�N}Y:�)�u���*�-�{Ϳd-��E��TV��u9��$�<�aw�����=�-��:ˈ�Ыi����RC9oj`�.�����r˔��-��4��UAX&���Q^����N�E:�pde��S�WN�%յ{�q�7�q��-�%��=�u�����9�f�Щ�|6ƫcsY��h���s���0:Aw|��,P�l���i]nl*Y9�v����9I��`�9���o�Ɲ�d\FÌ?{��T�7��|��\���\&;{���}���kςT��S��#�D�3x�9R�����g>�|�V�ڏ�����y̷�f��{����/:~ܩM�oT��3���)�z�A��Fs���̫���'��;�s^�3�<�e�z�a��#o�f�t��v�㤸������;6����eR�F�^eG���ZqOQ�̗�#�������Op�۽=wá�=�����5�O_E3�c�
$��)����>_n��s����}@=ɣ��Y@���%�o���|&ƌ|�b%su�T����V\�S�C+g�H�]x�;�MWBD���=�z=�ۯ{���wڻ��nu�q-�3	P�)�ԭ����t�M;�V6q��r��p���5�s�p���f^, �ak��<�\�Ag�u��ۖ��Ҿ����u0�f���NE41���ŵ�WL�d�:�U��)0��!�\�U�0om���N�a�?�������� �Q��1��S�jU����n�E�V�g�+��Q�o�58�ͼ�lFj�Yqz�� �1ƻ�Yb�Dt^Ux�uJk%���Qq�����)&�nkY���w�W��k�$���i����9Y_U���bV����N�3!��TS��Mm�O�")�Ӟk���pL\�+gҒ��B���y{�н{�~B*+Ld$�ʟ&z%;�0�E�Yn؍�M��^�EZAY�b�.q;�z=Xǽ]5��+��W �h�@ߖ�f�������5Ú��?p�..gbɑ視cu���������Һ�,�^dbO+\���Jof>�Yt��kP��q�A�~�,_L)�8v_;�x!iN�i�_��2��K��­w�nOX8a�'�,K���s���2�9�Fz@��=�K�������Qm�f��
?Dd�7�頮"L�r�Bٖ��L,SR2gn��9��Hф�%���Sy=TZ�P�TC$ĴKyv
T�˩Eʳ�R��}D1�C�&u�UB۵[�^�Yx(=�W���u�2;aUp��	�>��o?��xO��Y�F$�ϓ�i2��̖�,�����7�2�E�Oc�B���v$	�R@�=&;�.#|�ij�Ę����c���+J�ʖ1'5�a`s�2��;�(8u�L[�$O9<M�
�p�Cr񑥬�ݤ��EI�~��P�'�M�c-ջ��z�i��Jׇu��^�t���sK^õ�yRD�u�3ge��}U޲")�"��.³�,o��Ãu�Hw.1����D��孪�w��pQ��EϽ�!�PP��s�7"�
�(p��� ��N�.�[���q���_G.͜j���} ��2�ʸ�죆��w�r��:���;W���٧\�O�Ɖ���6���s%2��i�2g�
t��j��Wo��w���5��W��R=i��V���V�)���4�""�qq�Oo{zw�x�i�ʣ�y���9{g���&Ko�]�g����*�<��P�>�i.�w5�;MMO���V��7K��ݱ���=�������oJ���՛��8��r9��H�rjgbR�=�G��<	<�}�#�Ւ�Ȋڌf�p0R�H����	_�d��FRՖ=�-3��v�yl}~hG3��=#	��5�JX�H�m��v3B��YҸm����vPc�Y�[s���D�M/k���܁���k� _�er�\,�]=9�g��y)���fs�.ǵ^�Ow�J��:��e��KKF����bq"h=��<��s��ڸ�w5	�O=�3P�f��E��Yi�t����J��]�,��Q+.=�9{7�ޅ�3L���]������+�C̬�G��K�a,�	,��H��뺈0#:�6����|�W������nC�!��������d�bPV�\��L�S<I����Z�~X�uγ��h�f�)HmԷ��tSV���}�3p��b.���:�xe��u&���qYҲ���F�s:5�dW	��9��B�c8�S�c�f��vbD��੪��I�o���or��Bp�Z�t�J�r��)�v�Y��i�zes���%���ޔ��`�_�%��t�����
YVc�����\��S}�Y��3��[��$��W�k=�[��i��!�Z1W�t�f:ϡS��Қ܂0�v�"���UqN	m�2�LjГ�N�{&���h�.�|(�b��mܾ�,�O���z�Y޵W�����}U_UkN)>�<�f��n���bd���l4ұ�Jg�|߆�S	U���39��ⷫ��8���ם���L�qĭ"��1�^HW���*��[e��i����c�mO�qg�?b�}�3�>f�-�#���Rq+I�j�ڇ6(0��zDW�xD�^�F�s���rf�[�C-���t���}���bog;>;Y5�T��b,'�nu�횭��%�	2��l�\�^��a��m�#�:58�˅��6�u�' =:S�ۋ��S=&=���w��V��zQ�[O��Ǧ]!ze�YZ"zl>��e�*h�����b��U9u�ʻե���eB��V�0Ve��{�a��L�L��ί*��v��'���§
��y����zb���4����`o�֛�[hXR�W�U�|��=9ޝ��Fs�#��Ü�|X�.���R����'�243�`�K��*�|T��Yr����c�ȡ]�^>J��R��F�b�S�E�1{�}���P��x��6|�� �m�A��t̙�\�֭��J|�!�/�rip1=]6�b����[x�_*Xa��6�ѻ�;�n�#ݹ7�;����gkNAF��R�$3�6�,F=�V�>��3��O �'Y��9E�7
�仵�G�����Ej�`��|c���]����xZ����C=ݭ�[��W��L�qS"ze�<!2�%�]	�G2
�E�x�5��_�]���g6��:4\�3�CGf
��PW��1]*���c��<�/!�r9gpe�3d���Qe޼�;)�ْhqp�H��������â���踟8�U��ڹ���oBt�,^ߦk�\�=ӮGbŘt �|��Vy�+7�l���N�^��G�bPꈹd��I��#��c��ܥը�g.������E����ZE�:cm��X�}e�Gx�y���P��I�ᭉ#��2}�������诐�������pXci�݆1h�&�VJU��t�a��p{�wӯ�%��(L�k�9Svyf7�V;��W;2��ţu���F�.U�Qw���'�c�r��E��֤����eX��Icu�'9Ą�	��#�G^-���R��3��/;�`���Ȇ�a���t|�\��U�졑{�h����F�`͚0��$�ƶּ�ħ,۹OA��߹�S�l�J�7�E�ZB��h���&:���5z��v4��Z��n�l����a�p"g�D��ԛX�V���A�-u�����݃<,{{�۰��j�t�O�xc��ZQ_7NM�{%��FP�'gE��ח#�;�g G�R�k.{K�r���/��裖X�z�\���C�p�����?ϳ3>υ�N�g?����Cc�i^o)�����ʠ��.ZW�J^u��\)��zo*R��<�$b�JL��eE���w*��0��j���u�t�]\/�M�L��L����̢�0��t��D�r���1�+�K,ߕy3Q)ݱ��-9��c:秅d����ó�K��u~�b��7�=1%������� m�;��vIf�����i�|%FI#gMuT��3u�.ypu��(�Y(�F�=4�eS�c�^�C�
���Ds���t�dhQ�o�����kN���ֵ������f�J%��[˲�30�j�Y�)t�dd�:�*�Ӆ���#\gm񳃳^x焠�X��E�@��p�]�(9yn�9~�+�/7�zTc�t.p�t�1�a�p���fX��٧s���DӔ�4f0�2M.���{Z�)wӍ��-Հ:��z��	�z���'.�Ӻb�:Ȧ-��/WV	�.�vz��K�QO�,Ⱥ���nO��k6�����E�rh�[u�fz���̙���/rԱ�x��_qr��jk������X0bg�ħ���� �[uB((\�w}Z	�m� ���p�6W3coxLO��.�#��ɹ;��Z��0g\4��M�.���Y�҈�bS̏�W<ɭ<|rmq�P}�W+O7J��k�w߫��ꪒ��$�պćq$� :R/� �L��UQ��TF�6.7z�5�°��Ƈ$�_r��@�}*����8y�T-��I�u�z�^Z/.�੗qp��8=|�Z+"8DO�ı�;<�(����9�d
�q(\���'�M�[�;��/ğ�d�O���_E'�J&�Eg�:�)�:ԡ�� �����p-&��1~�)�*��/���	5Kv=�c�~,�5�wL{�V���c�\w�>����q,��n���-�2��g��>"^bS�[=j�����օDɧ(2j"�x?�7����>X�xϩw����<K����L��06�5�v�㜦!��5(�Ge΃Qn���l��-�q;(;�N�zt�цz�9x�V5�g.����Ճ=�l��h��Ѷ}���V2�5n�$s馻���|Bx�K&�����WO:f��N��q��S����e��҄>!җJ��W���7������
�:�ʛ�R:��爪yQ���ֆC�9���*G\B�!
��mD�d��=���[MJH+�ͼK���g1ۻ��O�cL�ͦ����N`	wS�Z�l�y�@E轝N˗��eU;�]HF�eoi2wU��B{{���k��t�9�%��ɀ��y�&��Ļ���
��4�C�-���T/4d��U�UUU�lk
1�*(��~�q���<�t-��d�&%�Ԅ��''��FU+]�)Ue�����;gĂ<_|� �
��x�� w)�+�.�U�wq�o��=e1�w�9�Լ���r0m��lUi����W�١-�}��Uq핢�עW�nyzC��4�X��\ݜު~�k��6.�X��z�4�ZWR���w��ޠL��m-,Í1/.����F�Wd4�1l��ʭ	�L*;��P梡��Lg�	�J<o���ɽ(_�h��-��j�z�R	^��;x���c��D�q+H�0�לȆ)X%\D������-�얽�g�^y�k#����23}�+�ܨ�=j8��TF�9�A�DY��u̼����S���So��[3GWM"��z�w9�'���A����
m�#EF�둲dJ./xoge7���B8cR,�@,^E�ɖ���.D%:#S���Z�ogY�T���.\�J΁�0�Y�P�z��Z�}>����/+�S�%;x#"+���er=p)��̵;p���	:�ֲ$�q����V��9�!t��?���}t�X0��/�V-��V!��Ҝ�+f�����-�&�^WJ�IYFH�����S=4+���=]��A�k-[�����1�t,쌉�	ƭ�9��H���t�;�%7��"=7Vo-���hփ_�O���[�k�B��5n���[<G��r���X>�9";h�隯�zhc6�<�s���d'P���5O�i�;U=�0OhOG�yV�]B���~�Biz�Zܔ��PB�,"t �=*�3��X����w*y�d���zRX�D��Ub�E�A]��5��Y��*&:�_?R�,qD�\XS��﹚
oމp�tf��Ho����6{4֣��\X*��`����ʰМ�NC�,���B�&y�|*���x���1�#=�i��i��,x�g,����vbA������3��s�pb����P�շ6{7�]ה��t�s�GX��Z��CP��D���dx�J���
��Dn��Z$�J�8P�401�3�}=s�u�A�I�LJe���ٳ ������.Q�g�Lg8�7z;�g�6g�S�6���p�$!������5ӕA��f��m��sYԸ�Ix��x��Π���0���.9�M�,1���1�D���|/D�%��BÛ��X1-�����q�T�rn�!�Xa[u�b&��\c�6�ᆟ_ ]�=�ݵS���� ���v���/��/f��ܽ�S
��>��Fa�@��uS�B���i`�7��� Rh�u�Z.�I�F�47w�K/k�,2�<�G���4����}��.p�u�G%���u�c<FN@zI�!�+����F�4��Sp�Om'YNeuUrI���-=�ΡX�m�tl�z��:p�&�t���˟;"J���8ٌL�J�˹�lv
��w��r�k�:��v�,�*K,\g�,\��̅�v{�N[�w=����;JeA�D\���S�Y�7l�n��4ȣ1�6�MyW�@�'�ɰEz�>DWY�\�}B���>	q[w)���Y筦���4S�2Vp髬�A���v�귁�)wӜ�	�GҔ�W����*+z�r��{lJ"���@��u^�Fx��u�}Y(�׍��6�=
�b#��7D�,l�ܾi!L��okz�f�
v��!�R�h;Sx]�cz��u�ӂS����,[C��6H��z�+)��F9;��B��O+::��Fy��pu��$����霎�8n� ��W�<勜Rnh6f�[yf�麯[F6Wу�V�۶�TJ`��N�|U�qIr���Tv|��M�?i ���\1�������g$�5��t/�Q.;0elE�t�=.��:��W{xϸ8&˻wm<92.�2�Y.�>��e���!{�+��Nk$��b��+.��睏"��\aꄥ��..��1��Rw֪�Mr����d:X�k^��)�Ž���ݻ��q%�B�ұ�On=���t�QZo1�Lf��os�G�a��|��_��n������ �R���-��b��U��辐����d4��Q.�O�ҩ��u��؈2�i���f�{(��x#9����ۈ�X�f֫ON�"xu�E0�ۦ�ܵdK�1�
8(o���#a^��C�_u�]���gI����5��y���APr��6�i� beS{��A���"Gu�t�͂�?W)k��Q�㕬���!��D;ܠ�G����)Y���!~�]�a�=R��L]�Y]�F��R�bU��mC��WJΤ��K.Y�u�N��]�YG� � �pr�1��s���Tb�sut���u��W�A��M�:kqq��ԣ�uG�N�����svi�ڲ"=r�+Ä�w�ٻ{4��,0���'�w�z`���\�<S{����F��T#��V����7zY�n}�\�	�֫6p����s���Z�Ë�O]�#�ّH�9���|˃G,$���� e��}�9�M[�������4��»& �����pG4�X���b�{��d�^h��I`�8w�������|s��Ͽ7ftJ�J"��ђ6]D5E:t�U1!m��������35RE3SADUTQ3SAUE0EV�4DS�AS4�TESQSRTSTSQ;�������� ����A[����&���*H�
�����(���")�uABET�i������4UT�}Ƙ���D�M�AUETU1G�51�1��E5DQUE$�ERTEQTTRUqi�f�"�����,`��Z�3��&#��(h)"�(j��*���"�+N	(���""J��SEL�ESELATQED��5��*�*��
j��0SAEL�5le�&���
**��"*����� '����\7Q�)ķtcFU-�G�r��T\�%A�k��r�J=�iȡ��|��:���ty� ����W����m%���uX��5T�z�Y{xGun��[,AN��$�E�;�"���ܠ�K���$��wL�e�gҫ�
��k6�����|1�	[Ή5��A�N�@�vJ�0����������K�#�����$�w f�*b��Y.�{�h�<08w��s�Q���� �����`:���x�&�7(�b��w�8W��52KeՎ�)?<i��]}"�މ�=����<��G�X}<�T
8sG�]�;��qM*�z���ٸ�{3�#�ݰxƢ�z��w*���XZo�#r)�Ӟk���	���6Գ�n��B���ѷ3��^�]0�v�<�ɚ����<�i��cVE�b6��=�[!;9Y��kvo��v=Yh��I`|bKG�?0(uė䌅9��X���g\�r���#�,���p�T
�x�X�c��9�U*��'<b��DV����藸���#̑�L��5���}��qg.�U�V����ֵ�<�L
�f��h6�]���#�)yu�;68�˓'w٘)K�:�eeu�ܚ�w�S��*��GE�Ǟ���{k����I�D�;��{�I���؋�Qvdo� Ok�+'A$��6�Б�}*��-V��پ�e��ϵöq�J��=��c�Έ&�ӫ�or(dY܁���G�t����L�T"�]D'�\(w��^F:OD.��x�@�0��I��(Ps���xgA�6^:�|Wq6X:V�=|�W��EC|�,d<t��C�B����b@�H LnډR�e���1˱o�A@ ڽ(o,kuc��;4u_�Ǩ^�˳��-��)���\s�W���%����Z<7�4�dJ^ �;@g
�+�Ndk.i�.��E��4r*�e�{ߚ�����~UqL_�I&g���߮
�xE_vU5���70�^�'�h�t��smo{g�[�# Rrpכ˸x��,T(+zZ�y7�S.��u���'��p���皳}[Eto	V�tD؜*l? -�]�r��a�ʭ��].^��sƌ���׻���r��7�p�U9cA�.��"�����tLc����Y]�xw23w��Oo���>����&§�f*���;E�V�c6����k�M����cF��<����r�圌�M�)�܎qӈ��g��V����^ZD�Ë>�ك�S�J�t�-��L���NŽ޳��!5#^����B����{ƻ��ʋ�:��"��q]�a�٧�fڇ�F|���"��X��6S��3�g_��5�w��EF�rWa�}�_o�@��FA^)U/_t�8ֵ]�"*���>���we�j�k�zz���E��������n�c��<�}�:4V�5,�GeN�j@�WKd\-�s��)�B5��@���*6vv���z��/�a3�r-����p�!�Q#�\��Le@h[���i���zl�H�����lPm�O�y�/A]���ǎ�e��҄>!Җ)P��.�D�OS�ݢ�P�ZS8̙^��Y�xn8}d:yQ��R����sM�ʑ�eu3L	2%{,tO�s��kz4oc�b*K�Ur����q���<�t-��d�BbPV�\�.	 ��K6����{��Et�[Z���h!�XN�e�Y�R=�@�,W�r����X���wgQV��K�JYch�h8ړc��J�h(E�������l��_��oH8���Sp�L���͕��Zz��U��z�4�ZV*W�Y����,:������d:Sj[�cץ�.���C�h9}\E��bøYD��Bx��S���1�kJ���ņ0�9�u�D_KZ�nl0��ig<����o��3	C�1O���۹�x�y�ٺ�_T��َbJ�I���@�l�ˬ�RTʉ凐��!�gP���>�6c�Q3@����{��^w���_,��)t2���m?=����O��7��a��$~Yn�L���<���eL���φ���:�F>�D�Wi�d���3o���
�ݵ�U�d�=���C徭.�oOϧ�_r�'��d_���T'��j���@Q�uD�����i�Ŷv��������+�_U�����X԰l�aM��Ga�CVF��/��b���I�m*�P��Y�rDP�	�H��
���P�^�0�/kl��芍N*1k�M�F��������3�d�x�e��a�n��%t�X�����'�J�o�E��c��s:��V1�%Zλ�7�0b�v����>M������tSg�YM��iC��ʼ����'D���Lk:��rD�V�
�%;����ƥ�ʷ,.ȧ�a��Ax�՗����(s��D5��:�'gz1(!�elz%�nt �ҩ�c��zVV鍹�#��t< (�%{Gl�&myb(a+E�%OԡF��T@O��)�#���u��A{F�G�q�{�Ч���nN�^BF�f�캢�FU�'.��t�X�G�p�M&^�]d�'YI����� �k�Xy�i���fr�AC�2]��Aኈ�T�γ�ʦ�5Ո��vG���NI�屷΅�{8���A�r6�����è<�Z\k<��1K�}}S�i��p%tCch��c��ll���\�7�Z�`�$�n;k���I��$]\�v���i�����`��S_�����������}�M�U�x�ŗ�/���r�C0��$C�T`KQ-��B��Q.���<#��,V�o�U�SgT՞p��T3�lhȴ���-3�q��֥b���
���� ��F�2��ܥ�Ia�΢��N�VC���K�� 6kH�,f�:��^��3���=ِS�+7�wi*���F�Y�P��Tx�y'pE56�,��N&�ŖڇWv�z�2���x��z��b�`dTc� y��#�ъ�ف%bJ��LՃkOsR�z�^}��HL�"#��{r�7��f��T8l6�n�t|1�	��IyާG�ӫ^[��YQl�T�[]ה�z�Z�d�{�iu���֍�M@^Ɲ�Rc��d�(e�բ6ڵ���u'��c�{����X���)��G!��<�TN\�,t�J%�p�(Ɔ��P�ms��o'G�iյ�ߊf��Q2c0��pM��ʠ���\w,�wq��=
�u��9[��\�B*�탍��>��Īvpg�ai�Ʃ��sc0����t��Q�ާ�C�@�1uy[���Ѿ�����V��.����d2�V*���=�{6����sDkjl�'o���ڇ��f�r؈k:�f W�^�d�<2�N+ǏQru{���;��!�͘��_�/P�7�E�m�}0U��p��Bf�/��ݭ�i9kk��~���%�U�C]ATVx��v|��Jwlr���cUN��Un�t�nnݧy��b���Q�l/�%���	���$$��,י|a���.�{�ϻB�.��V���	cQ���2`#��9�)jc�+G/$;�݁WYn�=�K;�F�k�ZG{[~�s��s5�t�B0�%�o䷗"��u-C����Yz��R1���[|G���w�&�%t͖%�e�m�6sf�/�#A��]���Z��g���|���g|������̱�<6�P�p�ǻ�kH�;
�s7O+�h�=����H�_	�F���Tƭ��0���;�N]��ylX�n:�r{h���8�Xp��k�&�\C��!��ı���{�3�꾱뱦���ux�tK��ׇJ��uqL\C�$�s�6�^Z):K���Ŏyla�Vf�L�sH�%�������Aһ��ް)P������$�ޅa�s�7*��5qp�`?������Y�1��:�5������o��8'�K����(vU���	�b��c̱�@ibRcq�[sN��C/�ط[V<F���v^k�v�_{�Z:���ݼ�6��0bsE�vy��0�v��R�ϵ����^�/�"[WPm��Z\�]+�p�QS����	Ġ2�w�r�vʶ�W���� d�P���k]�.�q��N�Y9e�JG�S�E-jȶp-'���n$\v�]�ۚpu;���{���IO|��nq�S�Y;eFV�c6���k�OCݤ;�΢4x�v
Y�jאrOb}`�Sז:}����^K�^���Վ���:��)�Ku՛���5���*�u�ʼ��}S��o��,��J�C)r�\����#�h��b��"�;G�V��̖��9��WQo�S��&w
��\;"���B�R��F���砺��*z�ć��3�z��U��ϩ��K���烼d���K�9�co�tx�x�B�t�b��j1�Y���wᵮ��M@�Ꮄ��q,=�}d:��E� ��Ni�]�#�U�A�=4%���7����v�%��)���EuT;�u��"��}d1P�зs����A_�ː�m�7���nT����JgI�쥨�L�g�'HK���:�ե���y��]����5�,_B߅����x�*�`�m�ǾŹ�Ydv�h�X�|�ls�ݦ�
U.[�����C3=7�϶Ӽ5E,KW.Z�f�o}����INJ��.����~��i1CV�I��@�f��Q\8�W��'{8P�{\�Z+n��(��p��S���LS���r������V�.�4�M+����hK�Lsٵ2��;����2�K�s�h�@v%��Qq}*�H��.�ë��k(��$i6�xs��k�T/�#�pg���͎AL35eU�cg,^�WLvT�d9�G`_��^sQP��(��Bx�����)����Y%,Dm<�<�Ok�lz�Hw7���nl0��"'��sm:�#�<M��b��L�,Un[~ٕȑYw��-x��X��'m��}�cj���T'���5DmC���W��u��5.RW���c\)�RXy��u��g^r�t����cg
o_��.u����j�P\�x��y��DpޘЦ)��ըCn��g���7�멏!�JtEF�P*,E#��:��v��5X�-�œ��X��6��V���ڪ�V=*�>�'�+X=�[)b���类+���9v+Z��׾^�l�<S2�oN�~$`���YT߼dx��u2fu�N璞���Z&�iS��Ρi�Ʃ�Nۖe=�.!��~��a׵-���.�m���ĩ��U���u�5���l��c+����4,&���l�B�ӛ��y-m��Hy�~j�7��n�U��.[��Jz��y��fE������]E�i�T1F�2i嚍�3��Ҭ�rg��m������-n)�WڰdY�a@�nzGh����)\�+�x��槹��r��e�G��{�)�ke>�+\0[�k �ȗd�d�Q[D!�	��~��r/����ҷ:%��@Y������
����a`N�`���KG�HV�K�\a2���,�]T*
��E`��:�pwN�d�J����"���u�hċ��9AACג����<B�K����ECӞxA���5�NvS�1O�	j�9"y���(������\�Z����B[�N�
M"������Up���:nK�72��x!��P �Ԑ�y�V��;�ԲbojW[��e�����u��n�t"���٭"\����Bŀ=w��Z�@���o[���
����©�B�^��{��㘓�"���a`uK�D'Cb�XcF�m��v�}���wS�ݍǢsE�4Ԕ5��QC�2��.���w��r���F��qι6�ٌ��*�#y�á0�j�P!�a��Mۃn��3�7|�;�|[-�؈c�C��]+��	m�3iGa�S����ug�r����y��g��3��đ�򘚈�KqJ����̡Ζ7�]�3�!F�%�-�x�^W�g��8���1�%^}��bE����.�d�n`�u�5)�0�MB,Z�s����R�!}]ï�����.w&�Q�Qez�W�k�%OX���"�ѳ��8ӻ��Nס�4�}�o���2%�Vr���X�v�4X��N�4��)����5=ǝ��氣�E3���*Q{.*W��ֽ�}3>Hfe.����7�ͫFG����5w�H�5����|�9�ǫv�ܓ/�SFM2�Z�,r���n�_�Ʋ��iT�66ai��j��ȯb���O|=�v���'O�yl�a���
�Z�*��W�p�mĢ���+�ٜ|�\�UdW���1��;i�t���`}�8VE��"ω���KG���C�����~�gŵO���E���Ι1LwSӏ�����a��f	�u��Bؓ<Ӫ��]_��7N�3��w%S{�rek��.��^��W�2����1Q�J%��Kyv}J���<b�8O:rWWR�#��������1�v�_{q�93^x�Aқ�G`�(�4/<��z�s=�lr���*5T]*(\D��(�c�5��wc����y甅�9����N�g����)�-�{�zGOw�gP��V���f��׹��%��),'{a�;@s;�80�ܑZέ�g���ɽ�i�H:����QZV��Wn¾�5�b�a�Ǉ��<��E:��`c�{Yq`$Dy/�ʤ��M�L�UΣ�h<�o{`:�x?QrNb�3x6��"r�E�t�;���p��Հ̡:�`<-� ��j�N��S"����GUt�jר�S;o).R�p|kt��F
���G����c�9ol
lS�n���<+�6��o_mQBƒ�y�]z����Ťօ�'l���t��eL@wJ@T�E��KL�Pk�-����;�R)Sa)��R����yW�v�,���OtYE���)QԺ�86�@n����s�}���Pm������	��(�H֒r;�\ؖ����x�T!�ov^9�Z�[D����;�J��^�v6�n&b�[X�^I��*�2����4��A:	�)��X������o�����2��/hl��<DMޗ�:ς1�fa���`��{��ejf亹��<&�^�#�|�E
��]x{s^җ{�^}d'a5�]u[��5����>�V�'VpLbS�f�m�5{ 3��k�u!C�i��:�=:_;d�2���EWJg���m��f�!F6/���v���.%A�r�ʄ@�4B܌ڐ!��v��>t�o���H7{�ZJ�^OZ�����8_l7,�a�s(�y	!]BڻvHX��1G/_N�{�9�!<���<�JT�H�'+2Ӻt����el����A�����9�ۗv�@)�
�c��,�ڋ&��:s�i�b�8֎��G��eM�5��,�CD���g�5<��N���ŹwN��s�}�l�S^��z��ƋV᣹��\�r7�uyҸG�nWteL���,���b�;�d���Ê��#���'>X������祵�u��|������x6�h-��ڨ�ݻ@֑�dfǂ��@m:��P]�e���+�\�Y(���G�U㇔]�E����D޸L۩[sDpT�KGS��ٵ�(e��Tl|��$�V�!����a��.����5+�Ds�v�[&��&{����o;���W8n���=��VT��cn�X����n�����Q�{TO,Z� �.�=���>�Yl�+�W-�|Nr��Ƅ6�式Y���b�r�c�dq�c0�0O:XV���aw�i%?o*}�x�'��ܱ������y��UUtn�:�#�8�33�+��i�3�8S{q�-qB���DLC�x��8$R��9����o<���eWZ�)��R��k`����[���ht��Ų������iЮ�D+�Y+�(��%ȕ��z-����Ȥ��xR�9nP�քxL��<��g�ǹ����8ﻂn�-n��b��׫:.��ӣӝ�bo����m�j˻ڏr���0T��O�跚~Е�)�WV�ʕ˟]�ߢi���`���PDQ2ETQMIUܚ�%����$��!��`������ �"����J*���*����j8�q�i����*�j��" ��6(*�h�����bH�8��LAUD�QDZ�E%D�D�LU0�D�QEDR�0��(���&���mEAPQ\X�i�j��
�����������J
��DQ�����������l4U1SS0W��$�""e���&�X��5DPTU��"��J���-��*)"�����)�*j*ѩ�����"&�*
�8���a�I�����LREEE��Jf�/��.{�+tќ�.�a�x�� >�4+څ�� �|t���=ͪ�z:�y4u��|w�]��O:�wɨ��Y�G���OW_>;�C�" B�o3J5�a�w�*�ծk8���+M�>��j�Eb��t�\�������}�t�N��[��.��Z��2�x:������2�[�YnQNl����+�5�Ѓ]&�E�P�ߝ\S�'9�f/-��TX��-�0y>y3�q/_r����Ԑ��tJ�	�H�6rp�7�p��%��ԹᛑT�T���6nV>���NNgC�~�tA�N�5
a�Bq(\��'�q7�p��VѿMO(�ャ�rǳ_u�c��#O׳��NY|X�{U8W��d_���������}r[AΥ{��O�saኳ��_)�Z~5�1��)��z�f-�E��Q]"^䡻l�U�&M�܃���x��)�.:�mMW�JK�<|2�7���]Qc��zJ�E��Ϸ&�O[/W��d��;<$.�� ۯ,-zRV2K��sS���x0 �nv'!v-�f�z���=�p�ON3	�Ӟ��Jʜ>B�r�.�+��1i��t�{�pt���İ·����N���/�9�K8S��G��Q�|��2%�ѷ�ᓻ�F^O��|��)��'�fdC�,���'^����[�Ͱ���IJ�h�s$����,y���Ë�ƹ��|wJe����˵���4�>�Qg�K��%Y4Hq�R&��1S뇞
[ه�w�N^<we�����6t��Os�U�@-�Bk9�5��mFӪp�E�D�(���!�<���O�����j��1���`ޛ�kE��	� ��DkWr�5)�2({�m{��s,���s���-�5�l��[���{�s�#�m�&��Ѳ��fZt�����c��MA�� �9��']k�^�Z�����AV�ս�!S۸Vm�4�é0%9-+���Ϩ(E����k%W�V(W�6rL�[ؗWρ:��mp�k�r�9��v,x,Lց��ZW�J�/S^ɀ06{`@3L\��eL�A���]BĪggèu��q��c��&3P�$������565yٜr�>��f��q�\�!�6W�"����cjUb�0͘x�F�;Q�d�����]#�ԏa�7��o��鑍�	d��� z�pS�oKGt;X�97s��Uw8wa&�f��Ƒf:�Q~����u�(�����djqPik����w���8��<pW��J�ڀ�Y&c�d�)�}<T+_��~�^��v�'�!���H��m&9(�2�BS��L[�sm�Y�]Tu=%0j�F�ʔ|�kŖ�_�"20���wդ=}1�ő��1���<4�Eܡ�<2���ky�g_>��ӧ:l"ڲ4Tkι,E�^��`y`�mWc6�"�
?a,W��.�v����sn.9�j�Kӌ�;C�p?�ױ	Yk�~�ӥ�ǥ���LO��ܯ+�N��{��]�&����b�+�oN�Ͼ�[�|T,mSW�m�8D�#0��R�i�eg<��i#��)��X�)�u������g��-1x�>�ط,.��#�ZN]ڝ��s6E�C��N*�N����B�w��J��A�D�|X	�X�KJ�,dUe`)�o(�s�n	6r΄!�:.m]��J�"�AAڇ�~J(�n#�Θ��2EF
�W��{Z/x��!Q3^c,��P��G��r�*����~���k�&^�}%�����Ba��^�K���i��f�"}�����V�X��L�Hz�Q��<CVY�˦a��l�{�:�%3��d�F8*���E�����������h����Z�m	A�P��;M苣�xQG�N�X*��������p�,X}��}]o������Ԇ����:�_�ǰ�Z3��I^\R�a���:��csmp>��b���U�W[��:�nP˫�{����{؆��f�x��\7:I���jw��kH���/-�����2)���Jޯ�%���;r�;� jR�ôL�``��R�����/��ױSYk�mR�i,��DLO^�D��I�Г�Ր��GB.���٭"\����+6�8��z��Qv����E !든�I�UL�㱚%
�tx�N����0���.9	����Qٗ��z��IW��p\�g�J��}4�4x���.:�o�P��e��]�����^nX�|$�y�vv�}�={g�����C;���F�'Z6}+P�6���U�d�	K0�jg]��w���I��Ap�@o���/t���]ј�.n��,�q1��Wg�-��]4�Vo�m�)⃽ڴFx���S�-� ��y��U����ڦ���E3�4H�St랍������S3�b���V�#w�VdEu`VS40Z֬�{���^>����U��ܢcݘڨ;5��tĦ��U{�`�cU���wp���iT�6c��j����s�-�[Y��җ9����32�����-�G�e&KJ�����Y�^Lԧvî5�Z¬��,�9������U�\E�랞����E�'�$�yy �� �~�d*��;�9�D���h[�7贼nQ�rKx�Ky{܌�x�XD�&S�0w{�Ri�6�6r�;�>�^c��Y��Y1u���9ֽ�J��Y���j8Ý-��gkܛ|�&i���u��Ohb���i�i�y�5��u�G�����;&�n���Sc���^ӣt�0�-8�J��a��f	�w��C��Z:S�c�[����f�y��C�.�$5�cp�=�,}�V�)�����Xj��|J'`T�����K�,�G_-̱N�Q�r�a�R��}Dy�^���3e�W*�_m�6sf�v��:��}۞η1�#�˃�x��\LLo\��6z^�Lj؇5�+��̰�˳k�)�rF���j��sm���/l$�ۆ��6�&����Br�f��7�t�t�cS3za(b�������'[ޗ�qwlޕ[u���a�$s'RJ���g}M:ær!x����Ӽ�iks�}��Ɯ�J׆w\>6�☿<�O2GY,���:�	9��H1=�:u�咰a�֪$��
êP/���+���P�]�ŔIa@VO��>Ҥ͋�y%���2������j5; ה�D��s�2��9Jm�f�/N\o52vNɭ��ZQs��DU[1W���d�Ō�S�E-j�b��w��$U*c"���t+5R��f(n>A��·y5E�������D��lu��h�N�Ц�c}����i�׫q�qa�
wtlǝ�_��`�
O��1K
�ɔ7�ul�{҉r����l�>�a����I�#�pԦ��;m�����y����n����%��-�u1������x��gP���Ġ�rļy��r��3����e1O\e\����/).L��ɋ�����-u�ޡ�򜼾p�y�{��,���Lt.��Az�a�n����j��9[��t�D�l�:đ���N8�s���"vPW�\,��=9�ei�[uóԲ,2�p�e�6ϧ��A�ެޥkze���0'M�!`)��1>�p�w�v�<�0��U�-i� ';o����g�e.u���UkJ�p�t���\�<#��}��.���k,6si`�fdۿ1��S�����l$Ȅ��WU�[Hz({�s�x���/�����@�!պ1j��
�Цc�tt�(��I�e3��3,'HE��4�O����i����;r��ںi�W·=�N։گ�|:�_N��J�b١�.���w}���S�R]��5K��� ȟ,�|�Т﫱`��bd��\H��K��9M�o�ϺZ��y^[���{��Ԗ����DM��P%= ᳩ.Y�YtzFBb5ʊ��x���70z�;�P �c�}:���IC����5�o�F��{X�rux�j.���}|tw�����vX����!���n�%�3�p���t�R���>��c��{��܌�}�e�P�b^\/�˸_!Լ��"��X锒�E�;kee��_�`�';��~��;��:��Z=�ua�0����p��[�cjUbv�݌�C[�2�[u���K�u\G>�8����ּ^*��+c��}�@lN5'�+s��X�'9K�'I�pX� �O��W�g�{kו�μ��<C��l�aN�c��T���'q)���cM��4<��B��:�m��Y��LK��1�>���z�ԝ[�Oj�~c���j�%e-����y���X�~SlkV�����MJ����f��@�Oq���'�!�S������[M����]o�õ^*5�vwĈ*�S|��7CZ}�K��:H�qu<���il����S��aa��S�e��^j��ɗ�^�qV�F�����,�\)zе�9!�����p=5YZa��`'1a�=�ZU��7��o^��x`~�аlK�T��ꒉ���&c�J(ߖ�PO���R���H�j¼�-W�w�i���d�[���o�����1�ir��}�y
,�"L1VHN��݌ӎw�dw�W9jy�,i�y����2�,w6�c��[���׃�!
��ј70�<�%���}*X���ʽ�`�.��r��v�z\�fΜ7���^۾.����GH���9I-�!Z�FU���ڲ�MÚ��l6����G2�98���؄_��Xy�i�R�b�)��o�.�ݬ���;`��ђ�l��NS��1���Y���r9g�4�����,Ĵ �C=C�m�W��;ߧ��|K͸)�_����27�i]�YJ�;�\��(_���{#�U��ǌ�KP�h��9�<;b���'�y'Q�!�ގ����5�K�0^3]oE��Ftn.Gw��HQ�ҬR|����MB�Ԛ�'`F��f9����u(wXsU�v�8�ʸf�92���y�a�)�](w����^�ʤ�����$�]�ҷ����Ҡ�K;0Aq�v�_����rF�t�'Z6}5P!�a�T�ݸ4�
%����ƿK�qi���A��|p��܎��m�����g�K��s~�0g-mx�} ����L�爔`AV�`����-<���x�&�(��c�L�2�7q��H�sv��1�}۷�m	�V$]}��kg�9�I�w�f�#�>��.4gt52�E��Qu�6s.X��֧��2�����^ue&�:�ƻw�]3j�K逓��!�0�Ɔ�f��R�x��������Ƃ�\�ޡ�]��#<�׃�Ŋ�}�%リ꺰+)�-kVCܘ�;槇k��]���$���3w}sy:���.�J���5nX�P�wϚ˅mC�WZ��E�̰�bM���p]��}|�
^��!�n��z'պ)+g�/%�=J�=U��Qr�����]A��d�Ӓ�y�w����X\�������&J^����%�����z� s�+�9��U-�3��=$N��l�4���'KN>����&8N���OMq&x'���Y�Wk�u��t�
1!�)���C�aYղB���*��)��|'x�5���D3ID���C��G3�S�uM=��6:OIAĹXmK�#3Ϩ�O6�P�t͖%�ʵ�]��њ78ڏɎh�����N�#��<%�>і�Cq=/�tƭ�5�)�Y�1㧆ٛ���s�ewd����-��9��@�~��"O����	���hC�o��R����~hC=���}��>�3�cb�5t8�s�	�t�="�|����Z��\1T�u�-��z��Mze���� -[4��˚K|��eּب�[�7��<�6eݒYq�c.V3=V���ҩ��y�UIw.��y�����4&q�S+�Ɯ[��c����e�5�)��Y҇�S\r`�L�v4�;X��s�5����Kc�UԯyL���p`�;4�5�uQ��ܚ9�>7�^ヽI*}H�,�ȫ���s��;;2f�GVr�� F7��{��4,+�@L�[�������I,w�������J�smeZ�N���]V��5�(g��: �jvF '@�@[�[��(f׸(rS�me��q,Ӕ^�ǆ���X�\>�V���T���#��I�FN�W��&�f��@C�w�/݃*��f��D��2����v!�/ո�����\�Hz�E"�Ok��u{�$'�8��G^�b	�W-��U���Ip�]O/1�P�;LWRV"����V2��N.kY�\y��S�J�t�-�6�~�ӦƭW\����R���%��9��,�fAQ�ޒ��C	+ɘ��9S˾�')��Oy��}�a��n��}�g�J��m��.�OUwj�6��P)���[&������\<�R��g�	z�����19�.%ש�/7'I����o�Hz�;2�&a����E�Dז�a�C�!�ʍYO��ޙ��oNN�ĶpP9�͛��eٜ;�>�2��}aiwsقH3ޞ�v���K� ss��9�H�S�iA]@d��hU4���hcyԷ�"���^�$i��X0`�38�r�`383�����}�V|;�)�9Jj�,��jT��y9�i���!E>*��9sz�R��:ơ�Mj�o E��Q�������җ����D��B6��s*I^�"�^P�����~�v��V�B�tS��X4�H�Ӄ��c%�[չx-<���+��a8��l;�7�� sR���Vk�ຬ�b>�:�=�!�|.[0��ܝ��^�D�x�����W��}Ş\��`R�
�+���E�޸��BJ;eK̪n^��釤]��2��5�rI�*7�Tǻ�L�ub�m頕���U���{�{A��	+�V��(+hD��¢��e�)��T0�hJ� J�a�M�w\�t-頁YFuq�V��.)rխŶ��Ą��"���|KDo��q8���W���\�{^��;w8 	�6_h���qBY��YZ"����ϑa֊;ē�7}v��L�g�a�m����9���p�[c!�[��j���6Ռ�������ĩ��dǀu��\�2~�)��7��Mb��΄ZNު���{	�3�v��6�3ݹ�k޵{����V���,�-�H��|�o��I��e�x�ћ(j��ݷyp�?K�N���˞���
�p��bf���ا"B�y�-�!�r�\�W�}�r��]��<Qx軯<S�1��YqrS4-�Ҳ��������%nli;:�]-��έ�r�d����S�}��x��s��!8<�X� ��j�]M"+�qKof9o��f���b.(t��Q�ק����%�M�z�G?��t��1�4m1�;5F2�h��R�|o�|���H�#k ������d2��� �. ×;K�������/=���-n�}zb���!J��	�����=���{&`Fa��2Lm�����-����$Np�4��b�J�/4�=���&s{c�%bȰ�|2�����}VH%_�Q��`�#B-�ª��=�X�gvN~�|���Q�Ͷ�,�j�+̗Z0�1&\-�f́�Z~i���=3Z�}��,�3f%n��n�ݫ������3M���=xu�[����*0f�X�ʏ�Ӵ��l�`�,���{cqk�+4�\��N2���aiV+I/L��1�KȺ'eZ�Q1ɥnu�J[�<�D
���G\��5�#VЭ�<{m���I0���ohͧ(S��a���B��g�vM�8m���'��:�X�n�F�,�R����pr��7��G@�����}���� BS��}>p�o rM]`�ぁ�5��:���}C��U������ˎ�.+���e��\<{T:t���
���đr������1!�GV��#���  <E��L�EIUE3QEIɱ�"��*�"*��b((�&��f*��b"-f�
�����`�	���T�I��ITD��Q4%!EPQQTIBSCKM:LA�K�KEUESUCDUE4�A$4���*�I���ZJH��:�$�*���QEj
�i�	h�����(��F���6�11TF�((�tDTKILI֌EQT�QkMAI�IAEAPDQF�N��ĄZ�αm�:�6��h�D�mB*-�QCA�uV�TQA}�f���n�@=���R#���K�ZJ����E�S}Z2�o`��x��^�ї���H\�&'�J�����%N��۲��(exQ�:��U��E���b�r��L�Ιx�V�̆�^�ޙ�/P�WR�(�'Rh��3��3,'HK���:���s�
�����,�@���L�Z�{g!�V���zi��u&d�$��S���f;�쬛�mS�Mj\l�T�s���3zrܻ1"�)�b�ׂ���@�r�i]J�-(�O2MJ'3m��2��u	� Z��p>,g5(wz�C��:;��^sQP�e|,<��Ukr?/p���а������(o�du��!�9�°�8+�9�4^�fh�3��ˡ�IV�P�`;�?+���.��cٷ�^n��70Q��2/��P2�q�%+z�Ckgｬ�~P1�qםji��o�����7]�a�[�u��7y�}���kd�if�\�n��6Ց�]�H�AΫP��pv|��c~�u1M��T6��8�X�^���=N*2ֻD�C��x�N��y�"��;%\^T�p5��L�v�����xa�WOJ�.�UBRN]]DMf����f7*u�i�i��	�E\~ޤ��J��r�,����#�^!��ˡ�����FMf��R���O���
τ�WI�k��a�:ls|}N�P>� x�����hCp +{�v>�K;��x�#ر��Ձ�uB2���1�[���/���Z�g��2����1)v�G���B��f}U��^�U���N�fG:��`�K��s��q���U�4r���z#�<�]#��BkI&3��q�L8g]8��1ei���k�
u��;��S��}n�U�E�CMI3�D���v��J�"�AAڇ���QE�n#
<�B[�ھ���wO:fh3�\�>��و!��PO��lߦg��DvL��J*ԧ~ڰ��~m�o�<eJS}(��ݑ9kY4�dw<V}�i�
R,X)��((x�~��-���"��cB�S���0˔�X���Y��W#�q�Ti���Q�<Q;G�Լ����j�Oi�cO��
�/*%120�:�<�����Zæ��s)ڀ������gN���eo���`�8{�i5'Qf�r�b�6��՞sw���g�@l֑}�����vUҸt��w#��K�'N���-+)NN���i�l?u��'XG���÷cq׵��ƅ�3��S53ff�V�m��gtK��ۥ`V� �X����Km���t�*u�޿�H����n]MKJj�fA]�{���=:;�I��}���u���U(�bs����B�U����*�_W9�E�;��[�^�.����rˍMq��.��|\�aW����f݆3�D�>GY!u;�(ue��Y�A��s��ev:�3�̧�j��҄U]�!���Աk$�|@���Y��Jc<���O`Υ�ͮE38-;j���g
�X�؝^�R���ƽ�.�Z�8_/Or\��1����SqzÛ֦��M��cb�j����jv[,�R�r����D�na�A�<�+�l⧶1�Q�P�s�[��Qf��%�w�VOM��)���y+����5�g���|��hM�ϼ����x3�^��Y��ƫ���J�\(��Īvpq���))�M��z����vxS_g�ʞ��/گZ��W�-Ѐ��(� y��fլ}���G��\Ou���* 4X�M�U���g�XI-�?0+��]��k&���2�'9*2 q�$.�,���p��	CQ��aߦ`"�����=U����f<��:ou�`�鑤��0��$.���p�)�̯j}<�LTC<���w�°Ю�uu���]�>���zצ祪ԡ������[�#^ْ3�w�ߎ�YɅ�w�^�#	�m����k0�{mt���_Mb>j�uh�d�=gۓ�%$���U���<U���
��J�SA�N�냐�pRMvKV�;�;�ø���J��L�w*�.V�LFc�#޼zߺf��k;Q�|��T�u��wE힣�v�t��N.�(Tr�����K�j]1����]��;�;C�m�u��l׵�g��sW�<l�D��'f;�!Br�P�5��_g��]��L�?��J%�{^�1�LV�ˣ��-��)�x$���'����#���&�(<t<��×�n�[''���5un�d@uQ��4r�zy��1~��I��$v��e��Ww���P��zf��y`gF�r�4,+�@����ܜ4�]��YD�2�E��7�
�WTYE���Ǟ�b��J0:=��D��Q
a�.	6Q>@�a�{��;�r���69.�qk�Բ��r��9���e��,h5�T�QZ�.+s�S�&1������|��w�/�eB��x���_�[�4�7\�g�^:��y��a(s�� ���6�pp�S&�m!��u�C�-:�mJ�xdK���^���P�М��Q�Y�{��R�|ַ�~F�����2��l>A$���\�鄑�b�� �r����oRx�s:J[�˸����n���^���N�����gbu�/#�&{�^ݛu�����+���9}f�ݹ���"٦�U5�)�+�>��~�{����<��֬��24wն$Ju��94{}��!u���l1����A�<X,;��Wʫ~y/%{�d��+Z8;m� \��%:�Y:zs��ei��F�RܭX�W��Z���{���:	��g	U���@���L���^{LEx����a�/:T3���1��&�l����u�ok˗<�Ƈ:R�Pު�Yص(���Xz��n�0 �օv�T�����<� ���t��ʑ���*4���"ZD8���򥴯������Cypw�g�L<�`93��{*����6�NG��j�B�H	�� �����%�[��/J��+qg3W�<�b����
y��˲�]�ف��\_] hN�Һ�z,?N��ܻ��n��X�] �p�j��t�s���ޜ�.�H��.ͺ��V���F�e[���سv�й��.���2�@��M-:��]B��]��:����r�S���GzJ9iCwQ�x���ib&���k�XY2�nM�B�du��!ۛ+�i���NE���@ա�A�.ܾ���º�,�r0�s�}���S�sc+R���c��P��x��祧x���S���{�󶔋���ص�M
��9���nhT�øz1o��u�
1gL��^bs�+8&��/�N��f�*%tkh*�o�����:�i莲9�/���`b�t��pwdq�'����)�#�۸x���c=�DWGr�&��dQ̶�c&
Чo'9Gj�8�Q�K�n�6���D5�m�8lŎ.O9�uڷ0��lk��'�η^�w����	��xP�pՑ���:�E���7��xn<�P�=L6��=����Tf��]�ts��m�!���LZ�\KÈ�.��a�fXtջ=�~Ֆ�u�P(���n�J���b��b��k��VV�������n�F-���|�t�s�m��dQ��WE�����V�T���Ȳ���U6j�h(3Jd�Em �"S��Ρi�j^��dfoWN3YGt6�l�·/3{���8#5z��� ר@BuӁq�PF�B���`^��,���/�Ao�z����T���Lm�n�f�Mi�[jgԨ2/�PPv<��<x�V¯����5����c�	%�`S���f��~�0�W�Ci�h�)��-�!ZvǮ�<�:�#�}������D�sK��G�D����؄X��λMXR�g+O��W��cՐ� �Sɽ}��RW����ySjt��.e�����y`��2�ߗ�a���Y>����w�{1$i>"`ǘK���T�Ϳ�s���v�4V1q�d�;�S�������f�݇Ri�ytk�����?qu[�<o�\0u>}%��9��k��/*��-�\���g�����2�^e�Q����V�G;	�7��u�&�x��ҕ-��|�яO������/�ylט�K�������*r�G�x7y!�<S�5�wB�FV���ءP���؞���:��׺�C��`�݅���Y�*~��ġ�N5�gQ��C��� EƩ:		����ƽ�%�'��uF7�S�u�s����5�Ӗc#�V��M��,1����}4�4a�J��.���D�ur.�Y���{I)��pIl�S�P-9�\7Dh��XVM�� E�������q��4� ����eB�������NS꺹�R�N�'�E�'�s���P�~�RAF:��\���a=���H�ک�1�S��𺙎qGE�Q�����+��-��Uue<�w�g�v`k��ED��G�4�˨�Via-���
:+��������dW:��{���1�W^���'�>�^>��σ�x{«"��ܱ�U�ho.�����S߻e�3HѲ�Ob5���
�l��-�$��d��J�j��uQ���'*�$�2�z��5�dv߯|��{�S=���I����w��ӑq�[��dW�rVa��_=,�ض�p�81,w��l}�z^��Y1�۽���o�-K������vx8E���S���a�}\.;��ԽK��:���B��BD�$�C�IůNtcS�d�p������t������YU��=��ϒZ=[��s6�h�R�D�J1p�+N ���[/�8NV|%G�0�"d�Է��}m�c]W���x�I�9�L�W�A��#ah�XV������_zp�{���0�?Oc=e��>�|%2,�J��6�S*g�JP�SW_�s�{��͗��y㒘�@�쨶�=栭�ށ��U�.�"�<F�K��A�2ݨr�w�+���V�=�m�X�{�v����^݇{���C�B��p �yؐ'ܤ�& G�ba3|-�;����
��9g�ͼ8��V3�)��<�i����wLPsq,w��H��M$����׹B��xf�vd9[k�Q��qs��˚U�Th�nM�n��y��0�y�6�I���u�Un�jU�IwxE$��V|e���67zI=2¿T�_��# T7'{�%{�zd��s�t+��-���</&E��^��9ӫ���rJ���^B��"'�h�ۺ�Biܔ��60Ꙍ����e�5e5�"�];�IN�=�:���c�;+�$�+�^��e"�����ʸ�y�_M�b��-��p�H�r@�s�����T�ü{��E�I��Q�-j�x�k����`o������DM�	9�G%lt/]�$��vþ^M�tL�*�nR�7B�R��yt��S>1ڸ}z�0��@��p�������G:���!����y�W玐�"���/�p�Z~4�!b��!p��v׻11x^R׳O{[�6Xt4z�����/<�'��bO\f^T�qӚn�P�m�.Pr4i�Ė���0v��������� �+l>YS�����/�k@ɶ��V�65j��^;�,�Y����Rf�l���vW�Y5�r�g� (���up�t��0�L������#��R�o/;I�叮�Fa~�tz穃Qr�LEt�H��[&�����T>�R��d>�M�H�pj�s��.eǙ���O(�tx*����EV��p8W�Ԣih��>�<���b��T�q����r	�j����g���Y��ϥ�0�ɚ`�L�I/_]��4X\xy�x�y����������H�H�<=5垵�)�ơ�:{(Ã��4'Rh�)�6�����2V�/2�Ӕ0�wQ��Vv(:�S{!LP,^z�v�
5=�s��޴�����kCܻ[\Em(�¡=ҵ7�L,��7���D�nq�LTo��752�2�gM��;�<{�T4\O[�w�I�*ؒ�E�"��_yR3/���-�]}�b>��~<ˡ!�yʲ�<�"��GQ؄��I��NO^�A�v�Ӧ-V�(;-�uw��@�Cbc*>�Kf��T��pC��=�ىN]��W
�e�̷�w���7����O�j��7�]��#�ph�4�ʮ��
�f��ާ,Ft].��)�\�%�UH�[r�G�I�w��<�1���҅�v���TC�9�¿4�
2h4�%�{��+�l����d�\G�]h���b�J�W�m-�GiǍ��rz��m�	rU(ybL9�޾�ȴ&�gn��2��Mĭ&��6�lPb���9��穋ʆ�g^rp��>��������.7�R��r��u8�<��;>ZLGM��<���e�G��/	���LS�ƵZ��9����vz��ˁ�N��N*2�k�M��g��e���6��V��:͸�̾cL�r�)��^��A?e�{4ȸ���=6CuB1l�,i�q�s�r�c��4p����QI����=�R����d^�Ȼ�a����o�iL���Aܧv3=Ρj}�o�+ǡT����"��	��U+���U~�ϣ��6�sfmHe���R�S3�$��^ֆ�'�b���*�=�����"{+�Z��˚8E���jN�r���5u���Wr�L.8d ��Rcjpu<k��X��+.��օ��{��G٥���-jًY�o��Vp������Q�ɠ|�ZC�B�U>���=/@4�;��
�]��ՌH������q�rx"���Ȋ�ײ���b�|��Q<U�9��ku�т�'R���\��:�6����/c=�J;�h�z�{��xj�ג-<Z��7G��7��E���5�(g-8SfṓZI�@�8����	C̀�0�gcoؗy{�X.��zoYϚ�"���16m�]�Mn-�&nfp�m����̛,��{z��7o�d����jf��[&�*�V%�ո���R��G���5c��`=���l�"���iVX!�j�+�S����rW0�]�oj�Z�l�������u�
��u�^�균GՑ^�CY��L�������9t����R���o����΢`S�Z 
�J^�W����]�t�w�U�;��> =m���CZ#3���6�2ĬQe�'L:>�����k�B�c3���_p�\�y�lY1S}a��3���nmӀ���KJ}�n��ռ|��t^ӷ(�fK1���Sh��f7WggEvIb����h��n��ss�RPv�(�͹6��rQ�p�R+�[�2�v�LSf1��.�;r����Н�}ꕏ�,U�h������v�q]���
t� hcY�I�$�אX�'���_��6���B
��v�{Q��M���	�Ԋ홈�lJ,T�� KY��%���q�6퀝����v�ۏ�o��;!�V�V[B�.����6�*����=%��k���N��(�K��nU���_;�i�0��<$W��U5���}� ł��T�
����,֝$���y���β޲Ky��ƾ�e�y;^�(��O�	X�
��X���P��NM>���v=���U��[��P�R�1E!�^!��y�J��z�!\��3��'��:�=�A��� A�j2O7��Z��N��xUų�ӎ�����@���7�;[�*@���&��rhsrُ�����(�5]̬��=�x�yRO�����=�y�vXIG"���^���]v<"����������e����ui�ms��N�P���N�ޗ�9>;�w��Tw=�"�-p�7��U!e�V�֏S������,�����ͫ~���i{���^�/^'�����W(o�w�^	��sݥ��\4l�[����%K�.c]$�{X�wJ�c\(W���e�_�����&���%ҷ-#�C&��m�h�z4o}s��!�]�y[e'S��f������ԟH��A��֨
�ٵ�t���LN�Akh���Hk�&#Vh4ѵ�kB�lX�QDkZ��U��j�M&�C�&��#X�6�BS6��A���J�lq���M:LF��E-U�[b��풗;�4�֍%h�h
Дcg���:��9�[d��UET�[!��dК��mA�)t���.�1)KEU�Mm�))Ѣ�&�њ)֊ح��i��Mi����3�litPѵ�[d�1R��%5IZ�Q�M1٧ZJ
�lb]�ɭ:Jj��6ƍPSA�X�Z�)�DQ�����MbM�5AA�&�+�>�"�OE�}��%y)�X&d�) N�Wݚ��Ɨ{8	36��v�4�/�G�����~���fv3�1EwV�%/��JǇr�����E����}GN|9��H�!�Ѐ�o_�D���t �L�=�ܗݎT�M��tl8=άOf���<�2(����X=),g�T
����f��=�=5/����Kl�{�-u��x'���N���1���aXT:�&��S=�>��xD-<�]u����"\L��l�'Η+���98���؄_<Vuه*�Y�i�ۊ����f]�f_o��L�˾��̕G�U�Xu.v���y��n�xݔ�*4�H���k���'Rᚳ������(젯����K���Hg��9�2�.gvc�V��v/��e�Q�al���=���#5�X��x(T.�W%�����I�6{�1�5�t�QrWm�(�o+�.浞#ZE��1��W`!~ ��N�RS=W�\j3D����n�OH�����׆��cF�`���c�̭=��hl�y�x���x��;�X�]�h��Y��y��\�`�����PI��)�(	�Gb��4T@wRŬ���,��r���d
aC��c��T��o�z+���:�4u&"���{I�ض�e��-p�����׽���U��ѣ<�Y���<A5)��%��ː�S��#�F��E�N�3S��)�'��a9<���f�:��`%�wʾ�
��^���z	w��>�ŷ֒�6p��N���W�ԗ��!���n���Q	�OD��­�NU�:����1ysA���e��բ3ǆZ��j� E'��1>0���n�j�;�4�-<뉽�8X�(9��%�p�(�d����Յ]X��h`j���5ٷ�䳛��Gu{��Sg�Zu��g�>�W��ȯk�j��!�����ᮺf�G�s��Gێ(�_WgiAC����ݞ�{l�;b} ����e�&��LEl�����Q+w%�&&��(�s��Jwldt��h��"��,&&�,��,�ݜ���-q�.���8*z@qNX�$���-���>�N����P�r <s�`#�l��qFwYF�3|�NYs�C�,)s!(����L,+I�c�>Sa>�r}���U�3=Y)�Y��x�S2#D�:N��'x���ऩ(l�XmK�#1����
�Ģ�K7y9o
�:���^��ּ��t%������v�a$��A̧J��w�J����y��ƚ%��<��9tF�?rCz���W}��@�A�ا��R 6��xme�d�C��ďvIF��T!U��i��Gt��؛�Z$�ׇy�vetw��}�%MÚX�����M�XJtI_D'
�Y�)k=ڴ�qU�����=*Rw4t'��|�`[��
��ϒў�����B�� ��b@�R@�0�ȾL���r��%UI�
R�<�4\GK�5l9��"��)�G+��8���\{
E��ұUt����2X�^���@��B�i�#ә���e�:���F��nM����a�$���+Ŋ:�Gyf.�U_H�K�"j&P�C�ܡ���I'�e�e@�' F@l�97�h�X��o#��I*����$���Xk��nERk.P������V6v�#UfMi�U��v1��t+ <r7sQ9�G;���5*X�ʫf*�b��7E�cRf�[�@֓�Eޏ��^9h�^3R���=ْ���-�J�/�p�O��s��șs�MM:nF�:G��8���7�\��į+�ܪ�SeO\g�VX��L���d���dS���sh�����,�
�jg`?VN�qq;Q��Jwq�S(����!u���l0�7~�,�9�j���=��Z�N��욷S��6��҃�N����a2��\:��1;�z��zr���9�)	qA��&�-k�73,I�X�gؽ�^����Y�ש�o�wn��VS0c���k ��&�vK88�����t
�Hq��dga��NP��ʚ���KC�����/
��ơ��]�Y�n�s��� ���%o��H�,����Q�Fٞ�����P&+�2Eǖ�l����W�}p���bE������7��^��M=��mҖ��;���B�Zhq���E��2R&��K_Q.q���_K�So:�=���s5��t^	v�64���"XH��]��-���'FO{/���2�<��nYT<�t-��d�bPV�\�-А'���(T1���0�z�-�C���bLw���~'�qb��+�8�X���wf�=4�é0%;0�D�b�}��t��v�]*��h;t�ϥW�[�w��_+�c:����س��ļf����~r�m��Z@z����Z���7��ʲ='����*�C�*�;ã�+:��=׌����i��.Z!��L:�'D���烩M�k��0𕸆�+3��Pxq��+9E\e��i����N�}|@΂��a��UBV��v�D��j�b�����t���/˜/s@�&^�j�3&	ݭFC��^N%i-I�lPa �{>�6Ӥxm⺧����* 0�հ۱`"�����8�'��B�?m���Ie�t�s6��lA�uX�6��iVn,<��a���:ɝЇ��H�@cb�O:&��r��6vetd�L��s\����6>r8��a�-iX���U�YR˧P��B,n
�Ò�^\ً#�5��������ہp4�VF�םr.���j�_k_:���i��Jg���ڮ"/kl�	N���b�k�M���<Nx=:+^u��blu����\��֑��4�yX�k�LO���x����n�F\-���z���-u�g)�=Pz-�8��fq�x�,o�[��*��P�3M���
��)�q[H;���p`ܧlj��S���mFч���N�ܱ���t�*��R�BԠՁB���#�Y��z6����ۊ:z� �S��>S�x��w5Mξ;���6���3ґU���U��fi������1�u<��$��(�{d1^	��~)Ӌ�s4<��C�P�N�F�)��9�uy����՞s��3՗b�]�*������W�.�<�c�P�S�5n���X��rD�]�2r�Y-�Dd8�Yؐ,��%٘*��-Թ�[� �X�ɍ^Y8�+ƻI�Xr�}^ֵ�7G_H��;��5�h6�q�({FTK�)��ԩ��.ٱ��NSq�f)دx۬H�hP��mJ�x�U�0SJf^�
��Ɵor��N�9.D�ꕎTO3kQ�T�e�Oy�*�t	o
%oҽ�Tm(n3^�<(�N���kψ��Ws�PM�{����&��r5���U}��]g|�:��xM�����G;��t��j��6�C�uO�jWI��B�er\nzZe'>�Փ�/X��.�أ�����:U��٭"��q�W`!q������ͬ��s����U�'^�&b�����r�<���MM� :��8228��ӫ�,�GY�IC]J�8�X�p�Fq��Ë-v藖�>��n��K��5�����#�~n��^�X��p��������H.� ƍ����~�0��.-�����,)� 3�5�G9\d�U��!�Jzԫ5WH}�p�@�;.}xd!��졗�V�����N�5�����L[�˽Ļ%eE�+n�+�i|�\M�Q���n�%�p��H�xFIl�^mXQ�Ձ4m�ʉ8wo#1y<��XY��G;v�������^����2R�/��'����@U�x�EN�y��-�f�����C��#Խ��M}��*zdR��V^̱���T3˨5ǳ+U�>������(�p�ɒ�Sy�Ӂ�Ƭ�w��J���n"�_@�x?]M�Ycw���˛p�f5K0E�	ēp%:��T�m�,���`��ow�/,�Ҋs�;��Խnz�F|��jjT3Fz�n��W�o�.���Y�RO鲥oy��)���^�)�Z��|}4��b#�xG�_e����4��Y�2����\?�+>z�_=\ nI	p�K5�0�t��>����U�5��m�i<5���U(Y6N�Z�7�T�`��3 �葱4ОY6�����e��p=W3+*�7���$���eE�yXx�%�I�]�R�f]KP_�\�(�b/�QDK;Ӹ$�8�*�%Kd�X��P~��W���u���P#�F�A'`�A�n�9N���P(�:�PV��sH�̖�,����7���z-�xkR~s�*�}�H�g�L&r�N]���P�tK�\G8��V��Lj؇5�a`s��9vv����)���H�O�o��ܳ�L����:n�Ur"���
�[�ǧ1������4[rh�70��`س�;@(1�g��5��$��rGY��xRt���ŎuYla�Vf�K���:�Ӑ# B�Nw2��΁X�>]�Q|��<�J��5�s�6e�Yu��}h��ga+F �'��4V!�n�cu�J�����%� ^'nR�[lٮ�K,��/ğ�;4��vY�\<�fB*z���'��ă�;q[Q�ἤ�(�pr�0䌫�w�˴k&�M��=x,߫;ݕ|�Oq�JX������{�E�a�z��D�㧠���˪U��V'U����xYF�����M�.��Z^���կH����|�-���T	�;zb8/�`}d���q���ƅ�.�nx�� G�_]�V�W�ֱw��]��ڌf�p0R�H�ǵ�w<��[堋v��V��l�܈�F,qКA���նE��
������ [A��v`���Ε�u1�m���������L�C]���;�^��Ui��S�*�u�@[��f�<I��`�V�T��f+M��DOS7��+5Bys���E�
�J������uOWx�x��^��)�üJ\A� �=���g�<ǔ8k5���r���4<�І�!Җ)P�˾��%D�M5Ǵ��aaj���gc5�Dkި�Ŕ���|'�g����m3L	2!$8����C_-�/׾���U��*����o�#��ˡ�Y�p�.<�,�(��l8qW�^Z��lr����Ν`��$F�OV�ĴV�Ŋ���l�<�
�}�+a�Y^^h����2����r^n�c�|�<:I((M+Ր]{>�Q�ڙaꝗ����7�-˳.˲2���F����5�8&�"�m0s��.�2�Y�c�J�TJ��=�������J�U��vS����.u/c��Y����R��;ET鯈'9#�w=�_A���i����U�U�8:#�*�y���<�g���f���0?7�
���4t�J�J�.��߭P�='�</L�����17�����5�G����u�x��4�J����]�F�Y�Л{M���3�����\jם���d�#��Q��1k �}�礮;S(1��m��dz�@D�7�\��m���ف�m��P)8���CTFӛ�F!���J�N���-�gB[V���O���hnK�y���RvS'_z��?S��+���F�a9�ӫ����v�R��	B�BL�E�}r�^�0�g(��DTjqQ���7糬�8�3��N������	�݉������5R�uK��J����b|D�o�E��c��˅��0��c'�i<ft<Y*��Wx��[��p�q�q�;&�ȓ�(!r*�5}4�)��+iw��轍��Nk:�4���j�t�avE=�:ps5z��[h�^��\�^�e�T��S�h��e��´�,
��q3���f�������FF�p,��X�JETkJ��8H&�nkK4�����#ʻ�t��{ㆉ���M�y]wʡ繡9
ZC�:?,�+^ҚGaR�XS��V�bЍ�HP�=�p�ه"��s��m�'�<��PC7jkh�a�cY�򈓊澁gWC|`[C�����UԤ^�+J;�����Aɼ'I�J1p���&^Ie��!O���.�����1�����#X��U�ɦ��:��$�3�\Ux�H���\ʰ��Ӑ�K4�uа��s<�T!��t��ѽ�I��_�S�h�G���(({%Q�T ԩާ�3�;�{Nxw���^������g
�{�El�48��Ԉ�T���%��u�B��Q.���%�r3���h�^u�l�\�W.ZX��9���T��x!�:�'Ƶ+����
���螖�;�'���G=���9u��7z; )vx`l֑t��&d��l��_ԧ'x؍h���EI�Y�nZ����q�PBjm�XR����1�j�0�h�$!f����M�k�.�)V3*_��������p7�]ˈ[;2�u�7$`؀
d_��<ƽ��ڷ+_E���r�CGCh�n�g�Po�%{8XV'X����Z��i!/�6��CL�Ӝ����-��+(��X	����ח4��vP�ɤGx���S��G	So*&pw����(�h6�z�x<+�s5g*�؀�ͩl(��]���˩��;:3�Z�<�n�4�1bF	��`����Q�u�`���sQ��kq7.wJ�G�
�M��0G0n�A�N��
8΋�0��=��<�I�^zk%�C=����NMz'5-��
c��w^�^����s����m㑅��n�5%�W�Ǭ����c$v�|%L\\�`�s^��hZ�wl\�r*C��_�<!.�0��U6w�JF��Vi�g��`lH���E��n�+r��0n�$<5Q��va�����$Xn��*��2����w�~>%Y�)�r�_sI���t�gm[�ò#v�;;SWR��~����>O�s
�r�jь���Հ�p]H�=J��6�ԣ���7��q.Ջ�k�{��Y4G�w+685J������F�&)Ф4�m�\wh�a�V��*f"3Fv-&f�
�*�ԟh�:�0��
2�w�I�|EY6&��B����%�e��Ҳ�
N&U��,�V�V[Ĝ#g'9��;�B��6�X� �)�-�U�c�B �7GkM��훬�}f�#	���t�s�X3k�&�dA���� yKhv�t*�7[���)�JH,�2�v�ʜx�,���w�y���NUD��4�wY�l9��7����&{���_R�D�������'����ơ��w$Lb|�\��Z�ԩ�ݝ��`D�w���|��3��Ɣ+7����L8�/�ι�Y�4-u�E{\��o:�6����-<~d���:���Fj������j�8�12�ȚT�-�\�2������x�ƪ�����]@F����;�ǵɼA�����$������ @��Zz�Pm��6)h�%�r�q�k�,#;���l��1ر��Q����@ͧ׳WJs�1Cǎ��W����Tx����J� g	��Y��m"bs�\��J��׷C�غ?�� �C�'�\�N��M�Q�*oJ�D���?fnK8�rn�l��t��ZՆ^L�ky���]�2��V镦A�8"�OAӾ��V���v���R��la�D��h�]ܚ�Ԯ��3[���XsH�8��.q�B�gB���Csc(�]�����Κ�(k
+�.�9�I����0���9��*K���n�t\Ӿ��\�r�##y�R�Ԭ�(�K&[f~W�����,˼`�V�V|�^m�
삹�J�ݛB�ٚ�޵�頔n ��u��yR�'�w��/a>bG�����qf��ڡ2�����FM]�����Mh�f>ည,cf����Û�L��n�4	�<��=��}�����e�R��i̓�p�v�k��L��7����$xE��p�������|-�X����㳯��ş��KKZ\Tѭ��4P�`�Pb֩����� ��.ح&���euF�֨�b1���Pш�T����Z�F�1&��T%�lb�cA��(JӭiKm�AI�i�Al�i'gU���RPSIV�b�X�8���Qkٶq��Ŋ1��)4�h(֫ƭ��A�&��U0��-�N��hE&�m�)�h�T(�cmITSl[ZɶŢ�.�f0P�sA�dhj��CA�QLl�:4[5�������	LN�m�(ꭃF�CK��[XӤ�`�jحmgA��0�TD��MQ�l�&�Z�!�-���))
��R:b5M	i)k4:u�ST�5ZMh6,�$�Ң5=�*��y��̆�.�C8q�6?v��Q7���3&�[wZwF.r�5��H�9�rb���qb�]iý�y�,��3
�M��w�C�����,\(9��]G
�H�	l�^<��2��nә�խ�; ^2l֬��1�u����dp��4��n�.ƫ�������3�։V��Xa���iq*�����5LF��ʪ����D�4ٝ퓴M�{�N�^��"�~��s��%�T�3�)ݱ��-0�c9[�=��V&�tX�����5z3݋86l߾J��^�� gd��7d�P���t���(j*M�[U��������:~J�O�b�Ǣ+GJ~lt�K�H}�WY�$.X�"�sY;KX�]w�:��S҃|kZ銄j�f��h$�.�J��Ԣ��\�7���KN��T�*��9��;�{���;5�xJ��#��y.�"�#A��]�(9c-چ�c���Q{9��-�:rP�nk���Y�2ۧ��!�!wp à@�R@�C��j�9*+m�n�u��Qryͣ�x�c�sY�3�2��?[�,9��7ް��]��s�$��;�T;ujjf�t���_OCS�أݶ#Cc��O�Z���hv�-���e֞�]�_L�k��[�z3/����9���KpF�)�brt�
����s����ڥt��¼���'E�닟EQs�v.�}��W��BxJ>��.J��z�7A���l�$�R��@�xev|�q������n��,�uQ��ܚ9��)� ���S��澭�$<�I*)��\yUw�r��3�i�������3�*ez4���Ew?�9?,r�p>퓆���,��Ia@Vs��nER0˸�^��V���1�ʞ)k���=�gd�t�"n% 9�/ʸ���f�}��˥���۞4�*|tS�@�>�N�gV��X�N���(h5��"��dO�lv+|��W钐�"���/�%�z��:彚�'���Έ�^^̨-���=|"�|no\K>�m�ގ����yRДhǸ[��r�U&M8�A�Q}(^̸g(91��N�3
eV�1�id��u��:�Nfu��q�y�b���s86�˝�n��-��m�$��)�b0g_jħ��z�yٵN�m�A����[/�ە�B'	%��j.T	��L�p�Kdߞ�
���.,t����z��Z�=�o�U�B�j�gM:8pb�h��Jo�4?�.$e��Z0��)B�J�����WvG3Y��fy���j�]���/w�l9�F-Ѣa}dS�eu:�B����f\��o���;Eo\D$�vН�ѝZ܋�nKM\�:�V���0�B��b���0Ҧ�pHX��:[�zŝ�6��'(we*�$����m=���R:��}d*�ʍYO�|'8ߣ��x%�0�	�`�L�I#�9��"Oc��IםJ]����}��^>S�M!�y��:1�r�<9��!t$��3��_�殩��m���!�Z���Rߖ:�ՠ���ü�n/w����ف��گ�챵�S:�O���7\�@��-J���9e�lЖ�>��UǶV������7�-˳r�vwB�zA5��b[`ꧪ�
�*6�Q�<��&��\e�q{����Ӂ�|ԫ�[��f���r�-ct.���c���xS�t��&����].Z<���]�;�6�Y.G/�G�]�V��.�a�"pV�a��uT!���L:�O��F���x���[�\ӊg�I}�u��{���#3��W�ʈ�P�*i-I���-f{�vOl8��Pi�	G�K���ؐ\�՛lf�f��/Jo�jY���bog���Հ>�t���X����j����Er��xT�cL�X�6�X�ڦ^��p2�Q��F\-v��{:�:vs`9�j�P\r�|�@���Rk^�2%��7^���My/��wunڰ�/���t��n��釀P17�6�2������e�`���Ȝf���q{׸�z(���q�MfI�WWeH�T�+�GhV�t��
'w���-���=Km�o��K^d��"�'g��yc�ջ>�U�/-�yt�^�"''Cd*�����*��m\�Xa)s��m��i�y���_���jݝ�Uf
�Y���lu=�i�ǹ+n���t�"�S������%+��Ρi��5O�vܰ�)�H��g�i�U���ʳ�sv�i�D��-)*�v���^�O�:��]gzy�dQ��`8=�c=V���}.ۗS��a��D�8�쒊7�B>�-K�G	�m��A���#F�kEu5���[�}4���4֣�2��*��`TC�UVМ�W�:\��Y�#i�B'wr���aCØՉN9^���޻MXN�b�fr�
���̪�qR�K����E������;.����}5�yL\9	k�Dv��@��|�CP���Z�0ϝK�Om�W���绽�I���pqgx�ёm]���Vo��!܁c�Z��I��P�]��K�����Fsk6hl��r�6\-u�Yn�vz�g�x6kH�t��:��j'�IL�$�[P�kvb�Iܼλ�f�`������K�^e���ӁS:A2�qw�B��~=cg-0�l�BṢ�&r�s�W8�'s��#�=���;]՘��ªv����(�l�C%&�K���y8ۂ���Y+��#~�]�C;�M�S�%�L�����Bt<Rx��PCjm�Y�.8ؚR���:��H�s����"kd���L���
P���\]������p�J���V'f@pN���wZ:v��T(�nsJў�����\��(��
b���5�|ݸ6��c>�|�.��T� v���q�7���bݷ8�;�㜎5�.�_�I���zv �����+��
���!�Z�A����?.���f� ���Q򖃞j{���b���.9��]A�5#Ի�mK�V��p��n7l�����Ɉp�7�Z�.�F�Ƨ�_������h2m���Ʈ"�׋��M�ft#H��\3����R���E����#r�`�<�twp�D��w0�FEN�m��L�Z�L�W�P�t8~�,�J�f�S�`s��3�[�=��S������ջ7��v=�e�ϥRX������`
���f����'KO�y��MZ��{�2`�a�7��8�E��TD�[�Y�J���FmWBC�
���Dr�7\����fz�"�%�f�}�b������1��]˞.Q��4�Ɠ���Z�8�;-J����܍&���m{-p���5��s3��u�f��^�^N���5�s�k�H1�Hݡ[hY��zG����w{C�TY�;2f�QT��N'�]
'���և�	f�ëd����Q��p%�� �L̺���W��r��G랑f�L��d��+{����f�5�D&#��x%�W���I��(Ps��w�s�&��Gt(��'C���\��9��o�e��n�ǔ�ߜ��� Lr� YU�Rĺ�~Ne��}|�	B��5��˦537�3��'.��E�b�ë�b�L5 �s�b��[��n�c8��OORr1�lT*��q�̃�e�:�f0(�����t�s��k7+�z�ьg�UqL[�$�s�;˞$����#M��$�e��]�Y8��\�汽Zq���3�prp�7�p�Q%��ԹᛕHD�˔3��d�%˦Dݽ�V@y�m��2����X��tD�
_"r	޼��א���Qq�ۼ�2���v]:NM���ydmk�d��rƃZ��!kTGy�I��@E���j��WB5�C���D�[��l��aS�b����VN�q;1l��`�؛���ۅ�cK7��e�D,�'���v�Ìݘ��.��rg���QޡW:�]�<��i�g��uDH�{�t�W�e�����)���&\~o�E,a@��W��c�)7�W�ً*V�0L���������zhƕ�{��e_W=�(�ty1�Tw�#��gG��_���f�/�Z�����lO}-q��-K�����ߨGkuJX�x��T^��&ږ7M�ei%�N�����ќ���Ur���-zRV2�`/�,��m�$�P�ׂG{bA}�;;;�g��j��/L&V�������,3�\)YuH�>���Qu�w��h�ɋv���ֲd��pv5��!���HWw�O���u�:�M�|t�(ox]�,�ٛr����C}}�V��
�'9�RK��k�!�����O�f��}���Hé�`��2%S|��U��fn{p����SG�>n�U.zMxc(=��C�п;����Ġ���\:������n�ԭ�d�p���,��i��!˩��uR)�A|X�<�{g"Kt꣨ɚ̧҃zwr�h�h?mI�1�'�%��`�lЖ�Y*�����[8}Y�F_�ΥA&\�P;���У�r�}��c�OZ�r�i]J�/�c�	�7-�� j5/c��=�;�6�h���=z9��6�¢�\S�"�梡��$��jIk��9M�k�����)�C��o��W+|�-�t|3P�G��&3g�UZ�Q�R^
�Cq^M(:F��tm�Q&4�B&�jxk֑=�|^9 ���!��TUéN���I> �N{�������7p��C���N%Ӣ���.\푄�Q��G�Ʋ�x_!(���yP��k]��aXsH�p�J�.�c��8�4:ا�kl؞�CkJ����Lbǖ�(}�N�%v{����P�J�Z�3|��-fJf-�F^�u���ri0��*\��f�v���t�o�jX6p��og���:���^���:�1�fܩ��V+`�W!�xK3�p�����<��/�`�U���g�{"[���z�HP�q�r�7�'O;��<O�a���^�'Ֆ���[N�ZY|k��71��b�
�T����7+�F䞵�v#�u&\=N��۝��4���X��tStxU��~�ML@{�2e��������6��p���wc3�B�Խ٦P�t�$h|�ϩf��Zv�V����X9.��{c�Wel���������b�z�j��u����6�Zy�[���m�}ڎ�|&myg
T<E��C��%A��(��!
��K��#���6�f ���*� ʮ7=1����B���)j �l��rH��L���e�|K)��p3�����u���t�w����0;�0C�f�ZfP*�Z��t؇>��k���\�zw�vd���[y��+�f��t`Yt>�\��f�z�2J7�skuu�;
/(ri��hBipv�Nθ
]�p��pGޯƢGY�����g���=��͔Sy=�v+��ZR,_�39g��%ٙ1�b�U'���pl�9o�]�xZ唶\�ŗ�-�W3�r!�T_!�08"v���عD�<"�֪���k{KAy�}�_�μ�=]p_��B
��c7�=s|{�u��A�Ƶ+�Rq<
����ü�ae�1]�+:�-y�	8��m�^Ր��Gd.��l֑t鍷W`!b���7��ӀjwI3��ݴ�U����/њ%
�Tx�BN����م��.9ؚ�3|����,@8��XP����r�FQrt�u��.ǳs�x7g�c}�%wW��ِ�F-����W�-��{��sv��\���l�)��p�nS\7n�ach�}Ή5�����`-'���g����N3��r8�k˹�N~�4�}Xd!��졑�4��D
�����1k&�@���&�s�����ȁU��;9vս������Ǯ��p��am�ױ��d���s��uaD��}3A���7��6}ņ���9���q�y���Ely�l�d���͜y�3�39����49�J�6��"�P��Ch�[XS�5,�}(�����8�|��W`��`�9�}���Y3�l�ћ����"|y��3����k%�|7��4�`�NU�b��[Ӂ�]׭��O��{��E����}v��cYq~��R��A�±�b6\��<�ر<�l�����{�Bh^���Υp ��BoԢ�_Ӓ�wľ��E�L���q}&�]�,�Z�S�G��P8٨���?I-�?0�W��B@�-��2��tQiR���c�e�=U�g��%�G�a�L�FI�w�R��JEh����I{����u���)���)P'/��q��$k��ȫ�a�^>�kY���(�|�h6�]��G#��m\��q��׻�k���p��S��G�z�hb}�6X�ʵ�]�����?B4'_�u�4k����踩~�Tx\J��,bfty�|�,e�Oc�B��p �;�꾎�7��%����qx�Є$V�oW��u)�[k8��1Zo�˳��nذnccf�^`��a�!c�wz9�$��H�-/
�X��������:8g���mr̦:ϓ��{Z��ϩN�`�,F����ޤ����]L���]�v5��M�$���6��-�og���i']�K(��~��x�Vv���V�d6%f���ӌ�9E���m��nr���,������:���T'��6Hz�ђq��nonҥ*_��TA����Z�P�6��Qٲ��=����iUv\�ʅ�|JtU7�Z�:]���6`u�ꇸx�e��b��}��}����;�	�yb�������Q�y����p�QH^m>�"��&mV҃��w.��+QU�d�:B�>�.PJ���;KF�S�H�_�Ab�#}��w�����O��יk�N�5�i�ΝN�H8������^����9��^�]E5H�."-���8�}��Be�42��s��BuW�,�|��w��la�6Ūʓ,��<�Đk�υ^Q����&���k*,��(v�?ЬeS��}��絶�w��X�vLm��ø=�؄yC��W�MW ���Ϣ��k`ـ�Ef�1t������/`�m� �����XU{lL�j�pj��5�!ⷖ:�N�������V'�k��:�c���ӑ��1T[�".��m�'Ҷ�����"�d�7K��A���o�;��B}��=D��/۔�0e�k7�L�.���NA�����y���f�Z2��
�pօ	��ʘ)s @�Py�_ q�
]5�ҹ�+���_!���F���j�ZtDϙ:X�xz������,�[d=֪v t8�����ƪ|JI:���J�%�z����bn������u�cc�w:�f��������O���v&V�@���52,�C�jV�f���nܵ߼����rn�I=a���+1�[�T���HS�vDi�I�7���2w���� 5���>��R��J�`e�r<��5��T��Y���G��[��1�V_��9c>�۱m�<k*��\t�{;^Wqr�B����	YE�v%�o�"W��n���X�i�1Z��G�.�y������c�O��'�fV��A���(d]�\��,�:t�fѥ�T�G�\2��JQ���k��g n���Tc��>f�BW9e��"����3P�-2�<5��8e�q�o^B��ɵ¶��&��Y�p�ZMB^h�� ����ɹ��x7��g�ܬ?$��vA����iͨA�YX�4�]�٪�|BX�ל;&�׃(UL�@��q"[��X]�{��|#!�-	��LQ�kx��Nbh�oU�e����Gl��7}�����e]]t�g��Q �Q9��'�x�:��XG��e�ۯE��u���┕�^�ؽ�k]��cGh������l�K��x�E(%e;�����ت�Y�h�S1�=�V53O�.����^)Y7T��.�I����&�A(8��qW;�|�<�6�NW^��*���51G�e�Mn+:�W.���郣��՝�
S�aںj�ZT��[�N��0��/aV�Y�%��6����l��Z5�������6�KV�"�ډ�4���5�lִhj4�h�!�E)�ETӭ:5�Y�R�C�@b�ֵCSض�h6�Q�m�i6�S�b
i
m�A����Z�(��m�vΊ�R�a�V��SA��$l�h���Chѫj(��4P�R�f��m`��4b5��V�"&��"�Ŧ�XM�S���M,@�V����t�)�:�!�%$U��T!El:(��(�f��ZhkF�V�B���c5���JcѶ�����Z(��#Hfm�:�KLA��t�Z��J(i�C�v4QMh�� �mEPh4SBQJMCm�l"ԲkMi�UET�5E�0DѠ�IE%%RR44�MSW7ۯ�q��w����a�׏���uSqi�Տע�����;���[g�1�ك�f7#5h�]`p٣�]��%����.Ó���߆�8�"�l7'7�p�Q%��z�^Z/-��w<�W��ew-�Oc{,ŮTA���Ja�pP+|���w��Sm�5�ie��x^)䜙��JiFvo6����8bщ��Y9e�JF�pZ���ZM�:'��n$����/�B6�=|2���n��;�T��,��s�9���d=WO_���*�D��Cu�hѮG92�)�l�S���5Y�Ao*B�9��e�&�b�e��v�WTX�x�ޒ��x�1�yR��A�c+i֗*����p�s�C�XZ�61���u9���x�U��x.���:)�tVUھ��|�^��V�-�L�4���YS�B'D��˖V�@h[�����6�z�{G��nt������\<�e��|͔�6�c:i�
�1Z�4Ug��BМ�`d}��Q�i�!��t������o&41�Ny���Q�QlK�a���j�t4��`�X���'�w\�O�H��ꞷ^��\ME���C9]F7�S�?5�!SQ�1�[��R̘���J��ܐ���:��W}�TۦCE]̶�i�(Kۏ��{��e��"K�1,�{ٳ\歛����v�؃:C���󳌣=���5��z3Fn.�i��+���1��muHuK�r�7��z�,nC����9�jb��9y��t�����g��!S��T�i��X���l��b.��ЗP��z�d�Z�zPqwӵ[8%���I�uP�YAB([4#A��eW�Zw��>S�I�t�s�p��rV��e����{o�v��X�=hR-++��]�w��L�)�Vn)dT�z�F6r��q�t�g��C��:;�)�^�5�Q&'ڄ�.�-q��*y���X�/{+����'�}0���9�°�ӉZC0�l:����&{�{�>���=۷��+=�beR׋��.
ݮ�pMF+lȰ�	ĭ&ڢ6�ؠ���~�+k@�����q���f���'H�z�[���O9�}�a���XL��S�P�ہ�T�.L!�u,�E��Ky�zcC�
�]j��	fW���7��׵�\���b���E��jwr��wf6O���	C̱��m�����U-��X����0�!Ec�#���1�n��3k����ʨF\v�@����mhΦ���i������dQ�bc3�5wEv����S���K5��-��يF{�`��]�ݮ��%#����O_�m���x
wJ�rt��x4v\3ޛ�7�c���M�w�]:]�_���#� 
�W�ᢞ�Uʵ��r�����Sɳ�EsN�)�޻i�X�>.�R�C�5��Eq/մ��Jwc3�B��>�X���Xcj��;����z��~uw`�i�uK�{�>�� +��9��\b��:�T���S����a�r�8��8��g��	e���PH�ka�Z|�RޥC�\~
I�(��7����	^��z�7;�ufqb��SߌWD����h����lz�#�0tw�Ih���(��hN]�Ý.V;��t�W����O���SS���"�<Vu�hċ��g,=��ă�u.v�s(��V��7���J軌�&D��b��KW�:Du���j%��u�B�u�K�g� ���ݝQ�$H�g/���v�ŭa��1��R��w�`A�1:MzO#ԫ/^ޮ�5x����4%��tS�G���ڙ��������:�1���B��`�2�����Q�WݸЫƪѰ\����T.5�P�rx�$�h�0�:��!�46.lSEӝ�����*z��7z��"�
x�
P�]e�]�f�n�+������by;�3Tmq�rj��2����{i��2t�O�x�.��u`�W���t��7yxx�n*9������9f�B�����{Omn@��*y�=���쫒���F�WCcRoD�.��ۀr�����x��盻*%w�d�}F�˅wRq�Xr�WbV���Vu�œ��q�4�z���}Cۗ�yYG�P6�pMۃn�>τ��2N-3	��=���
��`2{�U�}Qe8�#��#OF���p�Nq�i����c����<)T�$��?e��3��f�����: �-� ��yKA�j{�󾔧�l�����Z'+�n[�]�^~}���]'�����6�}]X��	����7�����ʠQÚ=��s��O���^�M�2�Z�,r��!n���q�e����S��!��j����b����5���=N9�[�g�W�L�UqԳ�Ѐ��Qr����'���� R^[BS����~�Zצ�]�ޝ8}��ĭ�Y�8Ih��@W ��! V��7d�Y���Kg�z��L��;���>��ųL�FI�u��Bؓ<Ӫ
�e�Fڀ���]���W=�#���鴋����p|�>�m�5
̈�$�vA:� �1U�E����/��='��=R�˗W���p�n3g&k��:LG��R�Hp�A��΅����)��"t�|4��������W�����i�<�R�5e[�kl�ir�H�f�T��М}u�D�u\y̹�U�x�$�(�X��DL���B�e
�_�Â�%Wd��jP]כ�0�<�b����X��b��gIk��2[�_K�a�11��ICg��E��C���o�e���Od<�.���5�&�H�[f��:�m���d�I��rС9c(-�;��U1���0�1Zm9vv��D~��`�o|:�El�fV+Ǿ�4�9I�b��X"��b^��u�&a�7��*[;O��D�m[{y]��{�%��<#�k� �c�μ�;Ԓ���~X��R'�� �Yb���^d�ͷ��=�gnb��vÛ��qx�	�Ld
���o.���$��+%���!u���>�ܮ}so������9%1���J3������x+����������������)hq�bkV�\Ed嗞�cA��N��"�/�`}d���]-�u,�I3Ѷze,8��҆�k�7~�c�e[4�7\%;YU�u~2����]�|L�fR�b�QW��f�Y�!��EDe�I�U誇R�\tf��8/դA��I:��O'ZY�;ۭm�k(�.#9g���Az�c�r��]���,�o0�x��z< ̓�y����2�WQ���G�`M����`��%W��Ի�ҷ����$�퉀��J1w�vn�`��h�AeĨX�$u���Np��X�J����Y�����fjyu3<F����Mʱ��1[݊��^�	
��nD���͟I�N�L{i65��U��	�ӌ�ei�n�vRذ�\)Yh�>>Z}PY����}�2��N<8���$>�)�X���'�{1��Kޜ�8ۛ��* �C�J;��Ύ5wT�Q�|��m8�p�Q:�Kq����*41pS�C	�6�*GZl��W�ՠ+�_�Ƚ/����pF�"�Ur����sϬ�*r��7�sɉA_�à��q�����^EGd�)α�X zK0��<2�f�����:�ե����f�<��ܾB4�g�a֫ս�!S���f��|s��3�iz���P�tmBXx��p�ݺ$n�3A:��mparS���4���z)J�*�٠��KJXUqLv1�.rgu��.{��Z$����U��U!��0���9b��^�l�J���].Z<��C���L����gR�/f������tC�6W��ӉZEØckΪ�1k �yk�M�z۪��춖��72;�E�JuL1��l�t����pM{�dXtT�<�u����u��/^�n%s��YHZ����!��\F��k�[绯���Ej�����d��9x]��AOpg(%�舝�W������!>g�\5�ZjL�a��,�x��=W��^Ju�����:���VO{nל�o�����3�`�o8�[����>>�AT�[��U��&�vIu����4�Ӷ�o�j[8PS�p�zd~���z�:�^�WqgG�~Slm�Ќ)��w(W�������\JtEMk��I�S�yN>,�4���S8�W��JÁ����J�X�J5R�<l{.>�'���5~�%Fz�Gz�VIRC���\7T#-m4[���[������rM3ޓ�*��`��N8���{�)eZH�2:^D���Aߥ;��Ρi��cT��bܰ�=OrF���Ӝ�¼��{ݙR��GpL��8�y!���wϻD��΄D�|X�)�`��KJطLl�����W0�9�3�U��*�a���(��7�����N�XUtb���yH+���N9f#�����>��{�UL��!ت��hN]�Ý.N�g��x1wV�N��/�����:Ӌ��lB/�+]���),�g,�PP��2]��A��p�k,��'�gq����'��&5}�/b��%���]�h�Z�P��Ġ�r�s�aJř��
o2�4�m�i;ٖ���6��~�Z���J���?P�h�l��"���Z�+о'5�b;�����f�dV,��ǫ�*��Nn��tM;����وls��䅆�����E+a�D9X`f���ꦬ+û9�؋<Wv�_��Hg���OD�f�Z�>�3��-0x!��!�Z������ٹ�˸29�,�1<\�P�X��$�ڱ�ގ�.���.�1���%eL�6�13՛�t�@x��5'U~��Ƣ3D�]��I���fx:��!�46�:6�ÌT�e��p����,���u��ƺ�v�^�����:�Ke(B���$o�>zWve���<]w��F�%u�gҵPWf�����;k��]'��}Y��װ�ė��B�P��:Ns��]�HŒp���3MAS�˚E�&�\����g��m�)⃽ڴF�@[L�o)`7��n�����e�g�u�=�%�8���.֔�M����4#$�5�4`[�g*8tM������)��>�����w�9���n+tĦ��EkhyvX�[���47���yJ�XtEð��?
ȴ�G�[�n��9�eu����3˃�l�Uh^��*��V3�D�WL(���B�&jS�`q3�3(��E��d��yH�vZ���P`�@P���ݭ�<�n�L�z��Ȗ� �x�*jE��ÿU�Qn�ߢ*51ꡞ�фD�i2Q����h����٩�B�9
G.��W��Q縴�Q�����z2�y�V���cwN�����</}=<>�J{J��U��I3�/��k�/2k�f�����n�v�������0�'KNC�(j9�q�d�G	�u���
���͎��hX�x[�j�K6�v�Hz�cp��!�}q\X|�C�;ū3�ȎJ'`T���1[נ�dPy�4
��o,S�J���*V�LFd>�Cqv�YT��<�8��do*O�s|�+V9�\C�hh����*�11�Qu�X��xn�cV���7�2÷.ͯ<�.R�ҋ[�����4��� p�@�@M�I�!�hP���&��n��Ծ;8����T��o��ٴG����s��7��׵K�1�8pu�9�4�ԚW�:W���bX�[N����y`�5s��<���r�uO	�Lo��8T\7P��:��-�g���~�<"j&P�40#P�w]���3e��+.TI��
ʁ���*!�8[��{��,R��Թ�sbC͙�Z��Y��!ŚW<3��Vo�Q�; �58� �� e7�qW�G,�CP�]��+СcNm+]� ��-=�i�x�j5+���2�tuֲM�ἉN�U��$1��ӥ%%���8����;��e�m�f,�rt=(����~��jwh����z|�'�dL�sp�}�=��;Ɍ��6�}-���޷�����\ı�M�x�����E��sƟ�?N����်���W��d1aa<�^��o�]"%���=�X�]+��L���1��u��TemF3p����k�M�/2��#�z� �1;�+}�o��7��e�hzj�2R\0�S���o�'��
�,ʜ|޵X��ʭ�������n��3����g���<�*����ߟ�h=:�`3��{�4�}���U�E����]|, �vPE9�]����Ӗ�p��՜�\)Yt���K�A�<�j���ў؜��|L[/I�Kdۖ"|Sۉ��I�<9��u�C��Rh`^4!�<�1Od�}vo���~�_��U:SyA��r��Z%����O*40�Ay�5�?]������S�&��ձ<�i�i2!$>^��<-�g�C��vC9Uw1��)T�v�Q��q���6D���	��#��А&��@��x��N��]o���MZk���UE����6ᮮK���> Ӑ����ӂ] aӟ$�kȡzh;��sk�
�+��* ���W��* �Q���+��TA_�Q�+�B* ������Q���+���+�TA_����"�"��Q���+��TA_�"�
��W�QQzQ��d�Mg�'a���f�A@��̟\�!���)@P�E"�>�� $   ( P@�i@ ���J�
U  )@ � $6�VZ5C3F�Uk�(����e�50��V�iEi�Y�����em4cZƶm�f�k$�EYm��U���m���R-��e3m��/���m�@�if���ѥ,�����b�Ԧ�!��j�Fڱ�ҭQ�o�rKDiM)�T���mVڲf�4�6�ٶ��Z�iV��5�q�6�U�x   �P�=���cOm%٩����5��56�(43z.���z��v�t ���Zt���WP =n�*`l��n���
ۂ���ٳf�mlm�m�{�  㾠-��n۾�ιP�4���@��\��)^�����^Ӎi����u�M4��\�@ SP�:�=+Fq��t3���;;�w�T͒�њɖ�j�#M��O�  �qB�
(P�Bνx=
(P���An�� (P�{��xP�
(P�r�(P�
{�n(P�@(P�y��
 �B�
/�R�N��嫵��U�����֒k;��l��m�f�թ��Q��  3�C@fV4�5���wVP4Pf��Ty:�mHk�dtw�n ��iN��r�aӡf�&�Jt������R����T�J���FK$U��e��USlլ�  o|��ꭝ��ۺ������4Ц������:-�9����ꕩ���ȡG��m뇯M4��V���з�ݥ(�wK^ۃE��)��^��j�U�]3Yi�hN��  㫽�N�n������t5G��5��Th]U�@��R�ѱT5��rj����w9U:�U�V�mmt둷�\{��]W=�{�J.̯<�Z�RV�ə�T҉[� 3ڥe46��4)�����@}mw�<��\���qvV��h�\�Bښ��s�TZ�O[���Ju�U����lt�5�h��;6�ʉQ��U�ekd� n�Z lvpt�(�ٺ� ��qEn�P C� 4�X j���	�h4v����f���6U�4L-lU�
ĭ�  �(P{���)GL�\u@�V ҂:�ݧh�;u�� Wg\($n�A�3�@
ݛV�f�e�A���v�x  u�AG�� ��ث�4C�;�C@K�v�ܰ9 8�\����A;�w@��h| ��*J�hF�4Њ~CR�� ��12���2z� )�A�RP�T��*� `@ I���*�OD �)�����_�?���WP�O���>�Mz�9A}w�~|t�'�/���O�W��� IOw���$�	&�! ���B��`IO�H@�$! ���~���s�g�h�6��E�����5��.=@^V)>v���.חqhK���e�����@�C��Iݝ6A�9���~�.�5aF����Am�wڍW;q�jq5$)e��;[�,j��ycgKp�s��t�Y�'�4w%V��g/h�)��7ڱ;��]o��u��R�Q7+N-�%:����t��[�^�km&� �mٚ0�_�zd�,�8��Z��Ci�r㏞��؁�K��
�����[��e ��4�`�7���gs"���oԶ2;D��@19�Ҏ��-�p۟Cv�-�Q���a�U{�^�F�޸���av�0*�ڱ����P�G+Zu����Q�OL���"����r2���(q3Z��e����4[��]ֲ���{{���םY��Z��y�*����S�{tV\
�'y�ѐE>sfB_]���z=Ά��wZ�1c���WJ�!�=�%��@�x��o����{�+�Ӛ�f�s��d�S"2��ynXK?��%C�n�;6�W��,�],�9�W���5�gh;6��� �<�ۮ����I�c��L�I4	Vj�J�x�K^�Y�[ڹ�TN�2]<f��Ɖķ%m�N�M�8^q�]S���B�hC��8��E��6���ý������N�zʖ���9�����9��;��őv�9=�Pn����y�5���{o&�U=f�ȠJ�Nꮡ��H��/9���&�j�\�7��)���ᵰ(7�a�թ�E��\C�0���+	��ԇ^�r��D���b	o<,&t%�.0��D�$Y��I��淁��2n�x��́���%�<�ֱ=$�w��d�{s,Yǆں��E�ѦCsnA�'WhM׽'�+<��������4p����X�:q\?W�P�OR��p=�E"�����D^5K0C��W�h/�I���Y5 4� �tc8�K����\�Ӭj;�ά2ma��=8���t�r��!LH6�-a�){�A���F�γ3�����pT���j0���|�@��3P��#,��Ktf�(q{]��*_M�Ѯ��k���h��9�+w��drw�酳k�z2�3��Um�Bvp�xk"�ُb�����9�M�+W&�hǬdQ#ysCғ� �#[��!�1�����8�VPq��BQ#U�Ɂ�6+��wR�Rr��/q&���@�*&Rٹkr�J%IbR{�����f�G6�ST�a��p����weL��㴁9�4S �uan��b;�׉qd����{)��iqM
̅Td�qm�:�6VǠ��1�]M���~8���wn��^s�貎_1%�M�D�*�Ԣ9d�1\�yn�*j��f�!�*|J{a��tn,6,��g��:��x�x�8j��yK����q�԰�ȸ�Z��7��EɁf��P�t��H�s�";�'�U��U�vc�\�\?���1N��d�n#�M�Ij΃l埍Er��H@���YF�|H7���3)F/%��;&SaCtʫ��ve �+nB5$�B+�!K]ԝ=�.����+y�Q�V��!��]��8�mX�m%k��%����r&Cc�V�Ϫ�M��6�Ӌ�t���{��ɪ]ymN1�,�I��1��/�os�V�ɄYL$a݉z٫)���rH	z��'cŤ"���n�d�ŋN��q���HDv�C$�sY�N����KC���X���@+�B������i*u�g-ӥL�ב���N��ug5hpk�`Jȼ����m}���Ѻ-*�'�����X��v���Lo-�֠�oDW=��'��D�ʋ*�D�ڝ�c������#)����4�X$5� ǫ7I��Z!��c�.;�%|^!����m��^�cS�r(�g��Z����pF�&zo^��bc�9��%baT��"i�7��b��N07w�٣8K�b�.Z�+
�&�v�ZĸI���|-��y:���m&&n�X�P*ҝ�^rvCz���\���ػZ!�N���eZY
�%`��&�̢�i&�dF#��;�(0�whlMyc갺�MF8e�3&�v�ۥG���ٻ�G:�վO9�<�K��������h�\���nw����xTf�xw1�$Uve���W$mW��^�uq�,[���7J�Ϧ�ĭ��;���w��N��WOs���GdIa�!qB���2��'����5Wܵ�g-��eܝ�Am�%���2K��N^���n!l� �/p�կ��y�k%�����r��A������T�e���|�}����U����7����n;��-��7�vD�z����u7�\\��˹�6f��x��(���Ǫ�z��ǣ�0��f+�Z�y}8�5a�(�ـs�Eɗ��&*7n�㗚D>跔�`sQ$xn/�7��;���t�>y��E�
���7��uMLr���1u��b�,�,��gi���Wd ,�r��L[Ik�|�1��ܨ:Ԝ�Fˈ��/Q�-�%�뢉B��y���Dy��u}�l��n��f��0��L��ea ��߁.�{��i(���2%���軲q���4n��.DW�6i�+�Q���02�F�Å�'Y��5�R�dl��"'���A���
�dO��Ȇ�h��9n�A�'L� �F�2|���2���/i]�P� ���B�mU�-2�1Z(n\�8C��Un�-f��!o��/�#^PqTeC��(�Ea�C
)�$�d�y��tQ���E��l
n��sЂ]p��It���j]�/��f�f�:ؑ�x�b�,
��9���bٝt7^�A�-�/4q��D.�Y��|1�P�ێ��:�O��;x	�s@cW���[�pM=Ȳ�������h� �k�,8K�>�j�;('�	����S�3��lO����e;d[K���QcR��WI!�ж���F1�{x�$]Xڛ/p�69�dJ�,��5�V١���s�����pcْ�8B���4NWd]K� �:�^�0DC�w�D����V�������qj�U��J���W4��'�
���x��4��j�12��&aL� 0�2����2ѐ^;����'��'wwK�!S��jiR�əs~yH��OA&�sUAU{\�����y%xJ_\�Ad��Aхw;{����\��)y���0k���賹�9aEe���̣%7P6尨7�3�$:�ӝwz8����h"rB�t�J��oA�]��,h̭�T�l����ܼc8��]�C�HɊ�}�@Eoo�u�V�rw,5k}��=�;	x�h��>i�
�:�� Y�v��z�5�5n
��1bA�| srF������,�޴a�c��~�f�ȎR�>;�EQ���5���WH�ǏN4u�S|(<��.nj	Ǻ�c;w�ĺ���L��q����+?	���}sNp?
kD��JǱ�卍���]+�sF1>90#-�����4�� � i�[�`|�s,os����<��sْ�a��09���h����aieF�H~P��ɲ��Ӯ��)g��<l˰��C�>�X�u�ޅ�����>�����7956��\H��G)��@��Nu}�l��7b_2�n���}���)`�b��LɖTgX�=�,R1���r�ڛ;ܶp�9Ǳ�]<���ӗ��v^g6�$+]ɺKY<�����A83{���vgnE�p���y�mn"G�^ݙ�� t���	�ۥL@����� +�Tﰮ*'v�j9
�w%����N?�����:�n���ƄR�FZ�SaܽO��\��f���Q6��5���[�M�B��KLtD�	mΪ�\��s(BK�.KZ�#��Ơyz�oB�<Y�F�ý�X���ٽ�)2�.s����L���!��"i쭡 \7U�����m-�1�f ���z��5�.�&��OK]�bP�F������B�B���䳱�!�lb�GS#���������E)�ܴꛎ�[�a�.k���mŗZ���dZ�b���qwk�O{�6a}n�p��N`-���;��!��o�bѥ���đ/7��Bn�L��fmY����$�,���7sA��x%h|:p�:��lZ/B��Z7O+HUS�^�^�u��%��<���U�
�T��Z�� ���b��^Sتdk�syjΧZ��d�&��ng<̬�]%�("��w�a`��q���wb�8� $�ȳg��sI����+�j��=��k�vXz2�D��T�c�Wێ|)[�xJ� 7E[tr�'�@ e-
��Z�k�Y�-�t:-���#��6q�-%�R�M�6�2r,-[��Ch>��Zӳ0@؋'"�@a[U��B��tL�{H٧\% ��,;\�(��ݧ-��G�b�7c�P�@��b��yǯj'�����.���9�r���]��gqňnh��<Dw�a���ęG�T�2��w,:�AZee7�Y1`I�"��Zi6k�.T��׳Xl�o`��#�zG�!�l獜|$��B��t�� �AYt��8����&ν�C��
c�s��{S�R!�M[�ڑܘ��L�T�(�ׯR�JҥYW�N�����)16�D�ûy�e(`�����v�$':�G���^��.휗h���G�c�kr�ؗgo=j6y0��w���m+BlnI�pʃ�lܣ�n�=ڑ<��W&��mp�.FN"�:����5N��˴e�J�B�=�$а��O��BZr�̆�g>i8;cCU�wPev��r�y�-
*��"��w
�\5�(�m������{���%��刍��%$D�0��KdS�D��t��9�R*��f姬ޫآ��f,v�R���U�7���:1Ɖͽ�w�&�#&=�q;��&�!kFG���B+9 ;�z^#~C�28H�[��V춥��5��q�e�Ա�Q�.�;���Y�2���2u��3-��2������:qY�+l�w�p�&-�м�a�e�lثɚF�Z7f�y�jc��7��6f��ܩ���HN�<���^�. �\�4Yw�>���]|H1(�ו��s�^+}g��7U�Ro����4`P��ɓ`���7�Ɗ99&jtI���4��W�X������y��F�ﶁ8��Z'\=M_U��X������:O`��[�8�Rj��;O�wF�c<�{O<�)e�Ü�]�6;h��wf�A�L�I�!k�Uk��b۲�����D�S��4���RW'�I�g#�[��x'�~�����gL.��B��Up ��ĕCd�l!b������l׵m48Nv��מ��	�%��Y;�?7��yi]�g<q$ ���e�����b�r�e\�Fۿ��j���]e^�C�;un���y��ѫx�s��}��w2��$[q�U�#��a]Ļ6LE}�X=U�;#S9f�́��p���`��hU�|{�='(B<$Ց���L��0 s�Ȱt$&�E���I�߭]~`���Q�'
�.7����4��{�����0��Z	]S�r��U��f��Jv��`����bTɫR�2��\�sy�j͘v%�ݛ��"��jH�)��%��X[i"6i81^��kU��*H��vDU��t̬����M�ob���go+���\�x�.WU�B��6�!�ha�C�	��,��,�U��WZ;r#~5���5�e
do����2;���-��P���^�Ĵ�^�\����p�u,=q��<�C���L��7;z�"�[�Rqv�EiG7F{:���t��\�t�w�����s�0���f���M�&.݅��}s�։]�K�!�dZe��q�c���1-͎j���N�E��Z�m.D��-�d�1���|��9�U�q�2cc&̹Jq V���"�V)XY\D:Ogjb�pF{��lO㽛�`=jk���v�=��H��=�
������k�G:H���!ө�ˡ6�:N��YIJ�a���eP�h�֫����Xc�0�!`&S77Yn��J �w���&�IU�(���t-�\��˳C�qY��	��QgM�Z�L\�Y�i(渱�<N\��6�[Pn<�*Ǹ�O���02K�a?���#�{\�!��­�M���0��%R��7�i�X����2�h��A�l��Ūk��^�;�h@���*P4��7�ƨz���Fs���=��5�y�q�]Ʋ8o>�
֏|v([��Kx����-ؑ���Gc
}�nXx��\�e.����l#Nͽ�6�Z��_oq�9��vZ�$��{�{j�I=*��W�䏖�u-����3����ͧ!�"x}3J���#VhJF孤�Џ��^b���l��l���ڏ*��P���Rd��܏C�1ܐ����&hY�[ߣS�t�g"�A��S��2.ݼ�<���Эn�vd�7:����02��.wvp7K��X�/wP��!q2̓\·c
`B����/A�:�.o<7{�.���G����pG�Tݒ�j�w�=;7��v}H(�_�������;w.�x0����Y�e��#��;�\�Q�u>*���+��]8��oR�y4(ܡ՚�7:u�W�N�y�N7]�O6xN�j�̍'ٺ�y���f��:�Ԅ����KO7�چ^1�c6^Sh�/E��#�����]���M�D��K�,� ]8�1�$�ZVjgɞ~e�nL9����[��F���C-�/Y3f3���B1|�]a	-�y��q]e�*q��:x�T�a�K�Ѿ�O+���(��]�����%((P �I8m�����n5�<f�~���ʚ�Sǥ���&�����Nt�������� ��u(�Ln'}bZ��}��\�/e�X�_S���ٰa4�r���]vV�rܵmeL�<���y{Li��
��4͸ܴ�c:3����p�z��S�����u;�w�E鈿��sX���vJ'�2��{�@o|��������8#�9��-xL~np��5x`��Qg��
�LTr���K�L�Z�?n*˕�]x���_��i]�:�s����s�m�?r��yu!�K�zL$y��^�J���&�:.���%;f�H�GWGW��%$D�=|5�4�n��s��Y�$B�_˺5�l�����wG�loϥh�n�s�Ґ9�U��:���ʼ�f����m=�"�X����;0�'R`���>��S�2仏�Ħ0��-��W�-���!0?p�s ��N�Z�z�JN�v
�!'N�s��|�V�f�OJȸh��;U�b����մu��G�������E�9����X������^ol#rMzL�Ow�l��>G�0�Ҭ�v�������!y�_kI���q]W�o���$m�vVBz*9��V)+X���.S
*��Q0\��XsA���!]��-��sUq%�~��4w^�x۶�c�'k�}�x�4j���*�iESv:z�Mx,�(������[O�����Oۤ�V������OR���o6���Is��X�'Ee	Q}��G\�2|L�¢�%��:�p2����	0&b| �=ؔ�0�/o�*�b�ˤW=�'�s�{�/Z�E� ����o^�k��=�7���P��3��=7qa�
�04��Cb����{X�wTr�.��ۥ�ƥ���!�����L˭J�d#��PW��u�T��u�z�<�}i�Iεl��
�m����X�C����z �#w��;�}�i%��6-�����$Gٽ�֕N��@��;oz��$����U�0U�ͽKp�@�5�5'+u�Ե]�r��u���ո�o��M��,�;y����}6��O,���7o�U�Ӵ�'���	8IL��];[��Ğ9|��Bl��:���:����+�gW�h�x���ܼ��l~�xlnd쥍L�b���6��y���N��Y��̹(- >E5۫.n�DٹqF�@uNӶ��$̞ɽ�Otsw<���ю��ḑTl�ΘU�wV;_�5�n'��p���7bBo9-$�x���_z �E0WZ�S���=��]X�H��;�n�/y��H�m;����s�h����N�V��:�.������7j�έ\F�z_�殒:�'�=�QQD7א d�lˈ�9ɸ�9���-G�-���3Aes1��s)��u(#Bn�ɦ��c�A�$�r����t剧�j��D��GG|��N�>���Ky� �'���/�*����_3�Ց#��| X9*�K8�5te.���g�N3��x+ޘ
�P'p�V2�s���B�z�%�&h��m����6��0���>�3�P�vB�D(	�|��=�pFM�9n��a��Q\s�r;[ ��}��1nٚ�寽&O9�]nzGN�y�UY�ͅY�*���5�ր��]��ďv�0��,з-*�̼K|<%]Ӌ�8���8�?���gh�&.'*28MW����:�S�|^��9��n��E�ecj�)i�}�\L� ����Cq�b(�^��r�#�xj���$�[	����)�Ԭ'���E�/��<[�i߮jd��E#�P��xj#��ItE��H:��獫3=y����nU�a���O���h�T����2)���7]>���:���+�+�s�Wv�:5׵��;B8��\N�.��fU�|���梁��n�Q!�'Q�I:3�1:�*YL:U}:�]a�.M�N�m�L��L��s�v5��]u:1D�L+�N^�J�Z�=FdB[}2�v1��>'�	�My$����/veh&��oy�i%��Ԭ�����9�����������(
6����SB�L�I��m�u�>B#�d���A��6���=�������ISn��3�3:�oYvy�/J<�=7�xe,����ӎK̢��ɹ��(¸,kȱ<�=;u��E�bG���̸�ɹ��n�6������s�r1\ȘkMEK��cܩ��m�k��N��a��L��%�.���Q��/����r��Y��[�>��f9�}휕�I��l�Qw22��h�;'ek��m��%G��aʔ�Z ����fR����l�e۫�Pޡ]�b��J\V &�fU�s
ųW&j�i��fʱ}-�[]��� s��R�K�����<%:��")�;\�S-� /(e�W6��F�h�F�WOUrV��ܹI"ͽX�^n������}�����(�|���yl�٢ۊA8[¡�9��Ks���[� z�����E�WA�&����À�mU�{+ګ�����6�37S	[�kS[�z�Km6�ZJ�+Qbʼ�)� an��9��[
?��k8̤�{.�t����j2Ԑ����qv�;�s�RL�<����J�l�{�W����	8�zպ�+��X{��1	Y��:Z����ҭθe��j�{����)_p泭�|�켺�}/U]z!�b��$�囝�s�c�У��]ݽbY�J�˩ٴos.!�#���}�K���j��Y�e�¦W��|�z���c��f�(*�R�>�B�w+�����́�%���h3�jr�Wa�n�Vu�5�q}�dК?�}���@j�Vvf����Q]\�����[KdDY]�K���=�͢Z�S�["MX��%�2�ޙ�^]�қ������-d�dgk+Ot��]J���L����Pb�k��-�p��Hk{0�p׎Ҝ����dK8�-�qVf%&�S�+�s`Q��֭����%]8���qFx�+H��v�\�x��{O	�.<{�&(Ǎ�^]_>ǌ�J�X^r��ʜ%� �dU*S�6�N��1�i����f>nV���?e2�ԅ62뷈hdR�r� s�"/�&�H;����"[��DL�{'B{w�x)�JM���A��脙{�4t;�d�=O.��݃��-$���4����Ĩ7��юa�ïg���4m�9(�v���S˽F{���g M�Yò7�{t1�n9������`{�xMf��!�"�͋9���Y~���1����7�/�t�'[6�-3EM�]XP��,�J��ࣤ.��Z���cQ	A������k�]�i`\����iSq�]tz����c��������}�����W�Wy�\p2����)҃����5כ�-T�I���e妨�e�P���K��<F|��s^�4oT�t�q��x�Vf�����%m=%`����tjhLR��><�"��C]4��|"���ð�
��΄T�
e<:��՛�y�`qd�7��bw�Rz�.�Qu�,���7�ve��3>7:���� Q]櫘���ԭ����ۡU��Rq��C ��� M	�&�(��/��/"���Mzݒ{x�� -͏x�W6�Q�J��^狄+���ٴ>�A�޾,��c�]\s�r��'uY�9���Ǧuw��ݩ�k�X�Z���*��e����Op�:�ۂ�[��ΰ��������w�*^D��CxI2��680����[72]ΥMm���F���&.9�c�k�w��u���)�:�YvJӽ�q}|��^�#N��ma����r�#�j�]GW.�s(�V\J�/�?�����AW,;�Dy���1����呗9z�f�L�`_6w{��%Y�ᛮ�k����{^����Ьh��2��^�����7)�簎^�p�,b-�����sK�⨗	�NU��9�mM�<�R
�᫶��A}2M[M�4�|1�r�<Yԏ]p��xm��bϳ/=mb��K�A���W)�R���g��~E̤��뫆��a.��+�^M�Z�)��]O�����G6�5C�!��jgyN�!�Y4���^%�z�Y� ���%w��CS^�;,bO����z_Ɋw�F����W�]L$��p��А��b�k6늣�Nu5�.�|���՛B=�����Sr������$v�~�F���j��~Tx��T�3Ͻ*1!.X����c��b��q�OX�\�
⬊]��f��[(偼�aԝ+f�܃��(���圙^��UV��O�+͓>S�Z��7(m�톤bd�j;	�B����(4���-�Ц�S`�G��|�ٵ� �1դ�Lj@&W�H(�:綦]�6��їt Ö"72�b���{�>L�~�gO<�:6IE ��{e���s���Z�.\0��foQ�xļZ:A^����ʾ�C
��qu��2��]L��J��|T�������";݅r�4�5KF�j_q<�Ͳ2��<��F�%��Sf|��a��.��`˨�#;���fź���h��A9���:�tlC�#��-w2b��{-٥�j/��3$�u�w�����~H�Y��|NZ��2k}�s�U��1Y�sPU�>�ű)�3h��[�%p)�\�ywv���7/��r��Yt�X�K^vl�H�f'�ǸSj�B��;M؃:,��[K[޹J	Yϴs�;-VT�`�$U�+)�.�ӽ�gP�D�E6�~�xGSk˾|�ܯ�z���%n��Lo�8w�0�{�'K�`� O��J���~��E�=��]���Lm��*��՛Z7�\���J�06�5f�ԭt�gG�r�-q�j���`��M�sk��,oAO���i��E�z*��4�\3FR��i�&��C�Q�r�+��'M�I�͕���[�P�>y�m�1����'��۬};��(����O/G5��S�1F�}��sf�߽t��	��@?M��y�<6�-������4f'�zJ�էJEN�Z��ηɝ����or�a�q'-������#�I�����L��L5�&G��[�a���&��������Oo���b=��b��n<[Ba��gA1;b���"�IK�չ{*�!l.���mժ���� '��T8*U+ߍ#*�]A��z���$=&�-ҙ҅7˲j��H3 ����)?���m]�ޙ�kXoc=Wbn�a�*aI1�!�����P7hA�N��}Y0q�t2�v$)�kNI��3y��T�T�u��\�蓑�UsM�	��0����m��yj��	�Vova$
��u����;l�!J!(M�/b��#� k��6w�D���yT� -w��z�+���h�3�h�v�1R��b��& �-_q���.��.�tM�<��� ր[���v������k#V�%���5��	�	+V�;�
S�EC�bn˾��F�D�ǻ��JO�A�^U��8-�^�Hr����ue�$r��u�����G�2��6`Z�U��e+2���j���y��P(�j{��d�5�K	�y/��(��тu�\�N�)��S7���&vj��5ǻR��i)���H��O�94��{��АƏr�)��wl�� ����⫞Sgk#9G_7���A7�l �+��\�e(A�JX���A��F���r�h�Rzʚ�M�j�U��q���(�"k�ڗ�x%��(�9�6����{md���F�\��'0�i�5Ղ!��:7�jd=��ī��R��q�6.;R�ih�������L,��Q�G�2�."j��]�}�+^X���[���/31P.��cih���V���DQ'`yn��cdP���Y��g%1<�`4e�ɖ�Vp�8����˺Hq��h��e=��*�{ӟf:y('�i*��J`��(J;2����<��b�)�ѿ/a�����2��v�~��f��}{ń��L���z΂.��.�
e,������NK��7�P�h�m�}#don&��,f�3��R��$y21i�M�\�59��ܣ�*dB���\��:7�F.�����{Q�
�
��ݛמi�r�/�;~�ܰA�sU���q6d�T��U4�٨��ؒ��^��3��;�x�c4�P�C:u���!1o]7\S�ֵB��f�Wv&��X��._q�������/�)����m�MZ;v�\��!7OF�m,
�*���o-�:�h�;fV�cM�t(Nk�G���͝8���<���a������[ {��j:��H4S��>홯��V�~RkcY�\ъ���V�vʸ�4/���`Ggun3�����9۳,�B٦�(��'q�Q�Xd�.��]y�f\}9�cxze��	g �T�`�˂du�]�P\�ec�y�	t
=K˗8��F�a��ٯkt�O�{hMᶶ�rLD�=3^�:��q}Xެ�lE|�&s��X43��x1k:�b����)��z2�X�T�=7����fTr�{̀�a�R%\E���΄�ÆP�l�C:;� ��[wN��*�9`�nБ�3�ũ.�&�)�]��nh�l ֨�n�ʋ$$=��R�-����
�]�V�xξ�&�iZvΈJ�od�R�r�I�{���xxx��B�5�����n��~�]�xs��l�u��j��:��Sjb<z��T\6�FU�I��zky��#��X�_yW������^܄�`T�f��7�}fU�W��A��6�����\�3p����������5��}�ĚoN��-,���r�pt2m�3Wf�&c'b��bFܾ�����vQ��%[�ߌ�7�;�d7&yd�,�7AB����pCe���eh��}Ȧ�"������G9LqE�}k8�ވqx�E�ج�hj��T�@��lm:ܫ��6��0�O:Rm��GɌ���c:���rh�7'��|N�z�]m'�H��kh��D�e��%�F����qt-���$�C�����6�N��*F�WiBP���
*υ��04Ĳ���y���6�!wbC��;�=�3��Z����}ΝE.in?C���mt�
b�R~Yα1�ŋ}������$b�N�@8��ڊ�ܺrG�F�E*�{bFj�a�0�O��Ӳ���-DN>�tj�R�Y:1É���,[z8��'lH����r�|�l��Gu"x�n�I}ǻ^��xخ�����F(�{n.���}��ZA�F�pr�66m-n�tq��LGm��|v��rC�E��/���.�<��j���Ϯ���os�nE�^'�.�kF��|��vE5���* �a����(Ա��{at���=۲WA����L�`��s<�lD�}���b+�d�m1���4���;h֮�z\�����[Mx7��������_�2�~�9�����g���կOR�vB�d�9�$����좨����7^(�fXI+��T3geaλV2�>���wH��ɠ�v�[�	���	YXtJ�x.zMw�O[���� ;[�Q��Y�F�;��;�:�|�R��4����9G���x�du�V"���^���ǜH����˫�����`|NNv�>>3���v^�j{����:'��P��}���и�v��Q��Q����c�ڵ�	�f��m� �ns9���;���Z���њ �DXxD�Ҟ9'\�Uq;�toX]M%�^ڷx/�yZe�y�Zt�Jmq��R���	嗗KNP U�yi��tҴ��Y�J�v����;�ǽ���#LF��U�f���ѵ�"�+�m�d΅p�ٲ ه��X�'N��99�����EF���e22��j���f��f�|K��3}����7P�ǝh��-HM�]�Rm05:��u��X&�-$S�SlR+LݫW��u�D�EPxJ*}��q/y�M�׎�dzk��y\iV�@��1(ls�S�RcpN�>g)pX�lB�<�#6�Z�gm-7E��I#�.��[��ϴ�q[�0M�R;�
�D���ހak�W��h���ˢd�9hl�&�Ո��f�H�a�(�CЩv�㩃w������\���:l�+�ukW�If��[\�s�h�u����S�)�*�٨��Zj�^���Z��X�Gifŝ6K[�8���և]W�Ŵ�4�1nOM��xd���2��q�j�;|����5��w�ތthb��0����j���^�����ҝ�5�bf�.��ȶ�&�6��b����]��s<�QNn1��w���g��'&���r[���<�H�4U���B��Gm�`Q|�y,����ܕM�㙋C�����aU1ɗ�3s)q�Wn��Y�w^.��12qn�f�%XD	�,��2�^��+1)�w�pa?n����|�̜�_u��)�t�V[v���:������[���$���T���O����&����X2B�Cc�}\^M7�S�������&�+9p��(�Pޥ"u ��<��\��}�ŘR�{���ny�{��jEՂ3$��T�E^}ѵ��AE�ɻ��}��xR��H�p6z���;�i�[!��*WpӹLl�a�ݹ�j*���x�`��[�}�+�(�����ͥ��X-��<�F ����V�����)I\+?Rq�=��0]ԮH�c=�Pzlk*^� $h�DHs�l��R���k�_sy^_2Ye��C{[�Yr�}��8�]�s9cd�L�c�ysR|��K�o�Uh�B�؅vu���v�h��(	ҭ���\xb47!��Ȫ�f�LSP�+�г�jJ�'U*ɚ������Na�2qD��W��=��yG��+�YB��R���BԨ�`�&������W�����ذ:���n����0�+m/n�gf§t�)N�\��d-�E���Z�bz<��ܦ��3͒��k�==M|<�s
yJ�ۋ|ޕ��7�u��u�Wq�L��[��H�6������YÜCGP�E�;��v��Z#m?%���F^����ݢ�XG�ǘ���=�y̋�.G�\`T8Rr;_%���2���^��L4{%�F��k:Ҝ��$A�5|.8�Z��j�)c�ԇ9uw�z+�����	�r���ێ�~v����Kͻ[ۭ���D�\)���G�۴յ΢�3v5�D�Nd�U���m6�#o!U��W,��N��Bη��O8k��'��ޚ�FBzX��}��]h�ňmn�T0���*HkY�qe��x�BL���.�v��޽�_��({�������-���EY��t�}V��<�0�G�
���X��g{Ibw2��u�2�0��;���ؚw7R����:Cv�#���B�8(��R��J��2.���l�{�o�������ZP�}�|j�]:��XIS�÷D�w{���NOx�.�˄Of��=^%a�|�T�uԛ}�s�Jii#�t�Nduu��wl�0�(��i�A43eY�'sc5a��Y�8�B�xK�.x����A�h�v3"�A{|�������s��=}K�(�ؘ�K��5>弊XD6v(u���v������e�[5���h�)����)YS;.�Z�ʄ���:�Oػ{:���)We,�1�<��0ݠ���Zj܆�Jzw�ֿ;�]㗹n�O�-�*�����F.���9,+,*�b��],8Fb]
C�\�N w4�w>K�&�F�O@r��L��-�����Ɠ,�Ȯ��>�ٻ�];R�Z��ˋxKt�x�+:�Ij�+�́��DwaѮ��v�.�"m��!8���{���Jʛ}��|���i�)�ǖ;�Zj<k��~��
EGSkH�pnٌ�f��elF����ݽ�/�����L�e�0�޹�r��K���Q��;N��%��B��tD����f�Vہ�ˣ�}�̚��{�a�������>$���p`�pA�&�+m���);�7N���Bf��A%PM�G�4�*����R�ݝk�"і�9�#��z�H�^12�j�h]���&��n$b��m��k�A�)����n�a���{��lY&�k���0���.�)&����Oc�]�/�&�֠�+���'w�,C����Y���D4E4�6ݥcS\���<5؊=�C���V�7�Z,���|3�-�H�jͷ#���δ#�ћu�3z�ZYBV��R�.*�,w�!:0�N�yK�Ɣ6�jv�&,[�a�
)݋s4:vA��6��N��x�!҃wh��yH�˵#�~����C�Oo�9v�E83Y퓞��]���˟t�n�����Jm
ZZ�д7W4*�pL�<��i5���EKK�e�}�'Mh㳪���^e
�z��W���g9��1fƜ� ���cX�E�6c�7�I0��Q ��%W�p���,l�#9B�q��w�d�53.*TԼ	�;��YwNZ��mV����]��G���Y��m����:����u���q�Z�p�m<����hb.�wm�hb��	���%F�7K�50�+l���] ��zv�Nzc�5�捊COb^+u�3=�Y����j��c�3�AP�#�����cwr���`�c��?�oe�-�I�W�EJ��׽0wv�@���Fb�g�A3����]��@u�wpJXE�\��[Ym<�ee,�PX3�$�t�U���cu�Re�	휎 ̬���LYO6�2�G��t���(V� �D����G}�������[|o��\�7:�^����8����qr;ݺy�a���|Ck��3�z��F뫻��֜ ͗e�>@J�{˃���ɱun�4��kIC�f��]|ù���ŵ�#D���J
+G�tУ�S�Ҭ�[��E�ȷQ42��r0 �;�\9}"���,%�� .��J8��wok\7�=}|���mw(]u @o7.�n�3�6c�vhz(�6G��-���ڑ�h�Է�\ۻή����up�]\��i</3R�s�%s	I6��������I�����Ƃ����G3ɴ�ו��g�,L�|9�N ��"�;b���Y���]f��h�uA�P�k��%��].b K�Z~v� �y�E�ݕ+у��C>ͽ�<tz����1���j3{Hc�np�z�p��uy�����5*+���њ��ڂu݀>IN��7���t�]�!�.�g%inf�H�^��kǵ|c�
nj�|�=����x�L��YѨ�*��*'f��R�l����<���;뫛e�ʂdA����@�7�Q�U# �(�j����`S ݇YCb׃|��.��=\��,o�6�	�(���a;��i�Й�g<݄��p*�5��ݤ;r�b�{]����-��ih���8�wY����� <|�n�݃;�)��ĩ���<i�܎��V��F��Lv���>@ې1�zv4������t�*�W֏wuș�ѫ�sh�m��
��\��t��cS.��Y�PGi�Ħ1|-���]>�ɣ�W��&4�*�v�M���]��k.1�r{8R�����y7prL�A�0%���eR��7��n�^RR�w��L�O�Ėo�j폗*=��������8�$�]]z$}�ٓ�aK,dt�{�ͦ�5#bިŦ�3v�+p�{+gg%�b�xw�m[�l�v�]����?m�1��}͊�'��zCKχcH�-Z�=�)@���Uzl��b���(��:ƶo��xz�g�pƀ�ۭ��sIo��f�ܭG7��)B,>.T'�� ���lFu��Ӕĩ�;���zd�/"\�s��"�0r�OX��ƚ���1��5V�åCI�^�t�g���ow7Dp-��<b����>�˽Z�lF�ԇ�o%R
���3(YDI.��*�o7\�l�QN�I�ecE<W�o��������|\ 4�ZG�1���ɑ@=뛚���\!M���ͷa�he�9�@0�T�Ju�*K����f+"`L]pɿK�7�/Y�P��31LB��M+8<鹩o���A#IBy]N�-4�>�����PM%l6Zwt4�]��u',�\%.�y����'Y�e_�,r̰�x�j.�7��7�t�]�%�f�sT	���[����Ћ�Nu� 9�q���Yg��Ə�Н ���n��8q-�S4v۱�.X��=K� Y[F-{���Sy;�oy�^$imB���IԒ�*�@���n�H��;cG;n��Lx����	�枮��[������eO^=�����a�6c������iN�@�rp��y���x�|�V͸r��VvL:�i��##h�w(��կ�Y�7�^�9P�ŜGv�R������s�T鸅ND^p6�Q�[��g���E��pv{�HR���$E�n�y7�]5uו�]��PI/�؞��^�S%�}�"v�Ş�ޝ<:�P� 
���E;�1m�n\Ս��A��?��>�8l[DIxn�t\��ܳR���f�7X��OW������F��[+�*kP�X"�1�`
�ެh(
[H�F,Ѹ���dH\��8I<j�����nf;T�L�*�ٜ*k�OK:�խ7-��P�ɞח�Y�\��a�
��<��s�µjʍ���R�-������6+A�'H�<��=�h]b�C���.^T�l��Y�ź�s5Y�M������+���0e������[�%�y@�y�Bj`��Kί��d�b�z4��g;B�u��e���3pP�Z/B���z;��e��5P�n}·���|�ǩ���t�C88�v/��[Ϝx� ��k)䠝1�k)�ȉ2�w��<����r����.�|z;�Z��ܨ�ɦ3��F��QRa_�zfₔ�����˳����H��3x���q{Я&r�ѩ��A��y�����lI�e�z�p�iq޷�ý�9٨�Xr���(�j1Z56�9;����ᛘ @��ԏä;�Y�zŸ��1־WXi>n�\�ŵ�t�]Z\�gٚ�BjW2�ȑU��ɯ�;֩˴V�y��[k��S��T�еl���oR��p�X�p��z�PM7��ow�F�Z�Knс��$nH��0z�՜�����^�J6�X�/�S��7�6���dB��������ѳZ����N��[���cƒ9���ܗ�,;_�y|u)w/>1�:G��i�k��>t��6絴���}f+�k������d�hlS�Oٔu��B�Y�E\�=}���rz����w;b��y�;���P�%��\}.�z�'��_&�7��}���Q#�2ۖ1M1Z��|�w|[Em���b!h�ċU�7s���ɹa��M�t�,���`�njXR)������F�N��1��ݧ���ʠ�K�b���μ���fJ�򚮟&r�oEXp?D�>��{vv�З"�V���d������_}��8&�*'�^lUy̯fgT4�q�A���N�j^a"3��8��|�p�P�X�@{8�L�3��l�fK�o�W�6*<[�ð+A;ʳ\*D靘�]��E�;X/bA#���\l�=�e,rȫ}L�FndI���c�ɷJ�)�������G>�K,����Ym��j���Qc��59�wq�^,FF�0s����[�5����#�۾�MtW�=ۑ���	�ۯoO|����.J��A;R���̩gZ<	��˦Q��򿞜��]V�Lǜ=�J:w����.�k���䵣�.�9�ܓ�s��h�j�9!�jg��O4ST3M�z;f����G��>���������a����r.���*��ѽ���S^X$��#R�3�-H�Y=� ԉ['+N���wck`��9A�+-��n�����.׮]�{8�����ቦFd����Eet�4��-2kqb����j�[;+8!�U���&q�̮�<^u��#�|3Դ��.��Ա;b�svk����HS��p����P�>�&<v�/�zWV�������u����\���x�8�,��a�]pL6��һʳW1�$��ɽm�$5������tN�(�Uٺm����V�䠹��^*��&B��Q���5εd�W���L�[�ڒK`�"��P���jԖ��u̳��&j�����z�Hժ�un"%Kj(����mU�\�X�V���pq�*�\�U�Q�A�h֩��b[b�2��Qm�ƪԨ�)na��Z�e�%Q��Q�,m,�ҵZ�э�eȥT�V��-F%h��QV�Qk+m
,VرKmK��-��SiJ�VЫm�kmB�*Q�����֢ �Kl������J�����Q�V"��X���)meD`�4V��X�R�UDkUb�F�X��U��mEUTXʭ�R�mT��+EKQ�j���-U(5l-���-F���-�����[meAB�(�lk*-i�J����mB�Ѣ��[��mRѰ�Q�[D�iKm��EhU�4��ֱF��ZıE,j�Ņb���ŢQT�lJ�U
�ڵ,4��e���J)[jƖ�Z4�m��*Ej�Q*Z�[m�0��Ե�m-*V��A�`�)+�/�'��W�D��E��iV���:��b���ͽ�n���3�w�U���Y�R���՛c�݋�)}��C��r���	Yr��j2=Z���a]���v�:��Wْ��ط����L�{��gZ/�����J�zD5C�nu����Պz�J3LI6s����׭fRm�Mzܑ>���Θ	�۬T��ܝX%5uF�\�=���r��᪳��^��@�!J�.�>�p�g�]�[��4V)Yّ�IevM��$OC��|�zK<��%.�M8��h���A4���^|���M�v.iTѨ{{Bj��^��������2��p�Y�4*k�#F�ֻ�WKN�����ˬ[gȱn�εb��[�~j|�7HɤЭ���j}ۤf�1%�;I_KW2|v
�,!#��S>Þ��5�ᚼڴ"�S�
IPQ��.e����ǉ#��������A�y��t�m�
�:����3�p�Qj�N��s���ԅ�f��F�Bط�yi���*p�4D��F���W�q���,2p�Fme֊�μ�7�\�vglF/E���x��;p"�Q�-w��x��n�"�Anf�.t�^�HH�rj������2|�v�l��>|f���M�����}B*�x��unK�P���7XW)��2)�r];7���먨m���W-��;��91-	3@�~�!�q�7J���x�V���Ar��r*:W�9���R8�L�Of/������:��8��y9�q�C������ީ'�����J5'z��Se�Mh�,��D��h��v�е~N��x8�j-L��O�s��Mwz(i������U�q��܄j�Bqo��,�&�Pƍܡgn�N0�[�y;r�9�0z�n�Դ��)ydy�P�O\�9݄_��uY1�u-��/����`��9������ ��,��囘@#�v�ʡ�m��k��O��tj�၆���a���&B8�K��ދ{ʦ.D�
�4�AqǬT�C����I�t!M��ՅM-20��:S��D]];⮗������]	�F�JP�@Wx�a�yj-?rߢ$}X��߄�ƶ��"�],���+���8!�`3m׌VؑYs/m�au�7��k��F�������`���CO]��p^�<��
qa�SB���8�N�չ]��U�d�D����hT��h ����[{����q�P����s�ԍ�Ƨ֓�k��Dֲ�{V�<P�uOOt�)����{2�;i�UϓWQG�Ƞ;�S)N��u���ܳخR�fŖ����(E�U�l�Z�o84�=�QU^��������ц�w��L���q�ЗL7�ɣ]�M��B$��Y��]�-�TXG�����v��:���"=R�'H&�q���.��Î-@��wc:�Be^n��YQ2p��_��`ʺ�54�g�	�	��g�(�%(3
j���{� ��$��*�o'C^��Vq�A���^T�<�p+�hߞ�3MW��2rNB7I���w��N���.K2ufK�U��sWS�K"��v��ͪ͌p/ M<�1���q9���
��Ý=hD��=��J�(q�����P�'Lی4܊q^�9��9t� ��s��wt�p�N�����T���L�WZm�S!a��vX�O�o_��S��:G:�klz�~����đ��2�2D��u4x�>�	F�M�,așӇ�*�g!�c���,{��:���-���<rT�
g�R�>�Y�e��G3�G�n�zbN�g�x+��7�K��N8ٔU���@���͆�t��c�H��H�e�L����� �.�:�|M�����m:P'*1��ݗcq��ϭ������Mq�SK���v㾧:�Wk��-Dj7W2e�g	���;�	L��J��^�J���I�F\��]�k��ݐ��b��\J
�W�����ǡ���<�{��^3mN���М,�!�#�8�����v8ד��Fުʋ�"� `K����-:㞙��2+��Q��	�iE��ӥ��i���QT�j��s��׺�9KU�����'ۗ$Ձ:I�yz5E	��U��Dz�Q����:�盦^9ۀ��U8����͈�x�bw��E��# �DJ�LA��u@���`���q�KYi�t'd��x�ݍl�I<�0�3q� ��h��F��t-��DaUO�t�m>]��{�Q�u	:�՝�Ώ
Ȧ�qF��Ӳg��<`I�+ό�'��U�p�BiָZ�a�&m�֎>Im��>��MZ��U�����e��7Q������4D�A��Y�P�/��\ԝ�`�G��}�Z�5=���M�@�����;]:E��ؚ�=���ep��/�\�jtO
��<(s;����gM��B�f� �f�th	*�[u�&KƦ&�:��D��Ka���A�{Y.U��G�
X�.g���~��bR���k�3x��F^� ��m!�iU�@fw�����������Gu��V,��a�ɼ]��]�)o7|�7�̠l���������:�%)J�mܻ��-���kx�$^�j�n�ss��CR�q���$�G���ް��`���s�0v��B��Μ��=�	��&���|��֫:%FK����J�B�x�(M�+Z��6�F'���R%)i��-Ӧm��ã�Z�O����:��CO��A�P"��VK�:�*�6gZ�5M�g�a�zdW4�2�:�q�9��6�Z1B����b˞eg���CG9�#�Y��(�R�P�-�p�������ȧ�֙x��{&q��z�#S�ԝ�51��_�h����W:G�n��畟B���Ũc�亠bCRo��0�������f�z8�X)eP�.Q��#J5�!񽮺�x���Y<�v�F�����	i��8�@�jQ!�Ѫ(Lצ�T�v\�N^����5�*a��G��$v�`'!��x����wMb%g4��F�5E�ô�#�椇T�3%;QJ��1�!���\^��I��	f��Qe\3��E4��؏�(��Y���_[�ȑ����sW|��0TWt�~�ׇ��t}ao욯'L"�Y�bCF�K����3��ґ˕]@.�����;��{p�pR:�����qim-�d�oQ��o�C�m�ӵ+��#�rJ�+ie�����\�{��Ts�G�4I�#�Y|}�\�>`�j�Lʇ��{��@ߜ���tvA��|�X����ĉ�KbF�Zyxs��ǫ��T��ǅ���T���5��ł�Un��$:~������t4��Ź�gvs�G�,GL).�	�8p�u^� ]��Y�s�W�Z�Қ]<�3�>n'*���;2w)Vm��M[v2#��_�N8��"������W�_U7Nng��t�)V�R��]�&�p��U�����ȭ{Y�~�	}V�v�dߍAh�5.�MV�>r﬎�8l�ٌ���j�W@@�����k4��0���6"k��i�N���uцp��G�;�̞^���s5��#�P)E�4��N�N��S��[S�yy�������^�r�z,��N�4�A�2�q�Ni�+A�*�4-Zvϙ΋P2)��E���Z��b��J#2H��Z0hX���:�HBE�����@N��,A4������d�9����I�$ا��du�H�؄�F�Y�04���/��cP�0�.�=�Ib�k+9��t4��e����eKp�L�w�ѧ�)h��U��=D��<C����[��cV��9�q�*�;�%�Dɉ�y8��U� ;���<���˘�0[�[G���͛�ڝè9�T�C����`�)��f��r��ؘ��)-�!�v�V�S�:V2�@w9�I8A���ʻ%��.�۽u�C]me侵:�T�}K�CRm_Wx�����.�Wm)��B2*�r���{}Kp��ޝeM>�yB��J"��7��hy(���;���{CuY1`�@B��{=�,pk5�sow���#K>[
��;��`*y��zh�����qr��9��gc�gI�����Ȫ���Ip"CL�Ԍ*� �մ���t͎�z���&�_���\�Hxbp2��xv�94d�ӡE�6iL���^�𶾈�nS�>�ȝ+7��6�\�N�&([����I�#���"�ĨS+>��h�����-���"Eڬ%b�7<�mc���7���A؛�Ӛ-F5�p��ˮ"��a/�/l�(�V[:>\g�J��y�E��O^%xv��"2������B�uy��o�
�6ܡi����p�1w�\��M�8�_,gC��x�=�,�Y�R>��^lk�{r��ח���[Eh��)7��K-b��e5���냴��]�ᙾ~�W�]Z4�k�dZ�^��)�e+����*ͦ�Yu�ݫ�34��k�r�9��*����9���)d��PC��&�t��/؇71�c�hM��C��u�{F���kegQ��U��k�ݹq=o�m;�5-�V�}���!杪�ub%ʖ�:�E��2��*�����須m�^�ܯJ���J�5���&��x��
��MS!�&��GӾ�!u2�sE���o,>8�p��d���!���F̉�`T�@��΅ĥ�q�i�[�ַ�����&n�y���e�+}\y:��� ��R�8��	����`,�
�t�Ơ��h(��L]�����4�1t�~h�*�ӈ�xڌ]t����(�9;���F7���8�	Q"vQ��8�j8�
���Aq�Xz�*,R(�ʀ荨*�m��gTɦ��j�F�"8��3�E�N�loc��A��Y�r5E�8B1��K��\쫎�Ww��l\o*��ՙ�|�uE�r�T�#Ւ�a��7L�s��o�*��%mA���#N�:��a�P�L�4�B5�����|E�q�es�5�����\�m��9������雰��^cʨ��o�UԺ��Eje��j�f���vZ���R�V���L�=%�tN�(d<0$��z3����X �;]jJ���xp�����k�Ȍ�*ej�dG�ؤ���nR�<^U�]Rm��P�lWK-�
�o���������b�>lsz��Xͩ�Qn���nh=p��݂��@V�;d������L3��)�D,.�@�j^ߒ�Y�WҮ�\�ȩb=�NY���>�2=N�"�o]��U�3��"^�*�ɝ	�銽����#*�ϔ�+3R$dÃ��dc�§��v4�ӯVd�a��ń��{g����*6��k|����YO����3�@���S8^��L�Τ(o{z�Uo4l$o���r��c�{�Fg���I~�㣅�A��Ud��Z�t~P�>g���~��ʇO D�����'��k�M����1ϫ��t��>W�kU��>8�N�ֺ�@�����&'�L���f���W�}�&�Hc``<��
Nq�XE�Ӧly̅��9*酁�#aP�'c�Ud;ګS�5�>��֤�]�Z��:x��_������W�P�~N�*�����|��H�ۺ�U��ZԎX�:X�����#T�QF�}j�F58��WV;Q�:�[����'�-��Y���/�B�T/�!��f��1%���k�#�;F��+>�x>��q�d
�pEs��<�e|�0L���7��4��q/<�x���ۧ����'D9W�������mY`h�.�P�]η=s�K}�{�X��	�sY7����^萛$uאio��gMZ��_Z��;Uc!�/$_U�w�P�ƹmNC�*�;�3t*���;�e��'��������R�w������
w��|<՗y��Jx�yE|���=k U�D@4��l8��KIȩ��ѩ�w�vykط\���z�i�5!��^������0��F%	��2v���Gh�,�k����,�?_�r�I��	f�����VC7pDSN���"��<�2�8h�KS���u#��i��=�D�k��x�ߟI�\�)�`�`�V�w:-	P���ҕ̜:'��æf�V*l�c�d��b�y�Un�$�+��2e�y��w���@B��g�<�J�0|��!���U�`���{ݪÅ�3]�V�BB4�Eg�^�h�Øw���D��Ae��J��i��#�8'W�0�V$afn�{�{t�Br{��y�6hMO �i~>��_\�Z���H[~{Y�&����#tD�b"�s7�Ns�3��A�v��Ű�mC5sT�G ]!��8���6}CO��5畦(!6u�
AI��Z��w7���z��5�YB�V��i#�r��Ny:�7!��9�4�mWZ<�r%�˖�ܲۥ�(Tkr⽫y�����wF���zFN��Q<���}�ϵh�;���V�z�V(`e�6�~�I�d�ja�=����"ҩv�����
;�k����g:��{�<��0�B�v{j\�}q�q���-j�X�����8~>�jL�:S#���]y��y��j�4ݛqI��<�;官N=�����9A�T	��|o
��;�.���H�l�BU���8w�Yx[��O�t�M�����3c��v-7B�J �;�q��4��x3Q��;�^ѫ���E�
������@b~�py݁29�O96�T-��4jd��4l�+s0����M>".��R�\ܣ�U����v ��3Y�{o����t`-�˲��%h�p^�9]S��}6&�E망/�Y�OptM�4�![P�h�}��P�u������<z]v��
+f��Gjt�U����(�� u�WKD!�#;i`�kȷ��#�]��kr�P�eԮ�Y ��y�E_{+���s���@E�t�G?L�������9� �x.��&� �۩��ȹ��e����Ci=�)������1���������0�s�<�<�7(�t�s�}�x}/�z*���J���Z�1����9�*��6jT�!��s���an��^f-"K��9t�X�{�,w��+'%Ұ�8�oT̰(�7�{8�}"�bIt��;�>��9��o�j�ag)�H�^w�_wq�66A�-����(�M4%Ԃ]�׮W��穫�LB���*'�����}��yÏP���Jgd���ӯ���s�r��[u���+]+�[g��4����'O"�����M@��}G��1���b�s��|��N��4����c�Q6�kQn��u��-܇uB0,�9��F^���ҝC���1%yl�<�+2�Hpms�K���z$��])ʱ�/.�v�N�ѩmقSMx�ۼ���_)D�ǝ&6Eu���zVn2%���-� 5Ջ:�s�/���Sa�O���*��b��kD�o���a9Bћdf]:a˛yҞS�1�h�l�N�Sb�+��׊����Z�TJ$G٤��ʑ�|ӷF�u,Fz���^�\k�Av��<�h�$�InŸ���m��vk}�g�TS��Ф���t٥N�L8��X�A_�R��������9q]�s	�M�Oj4�NUe�\r"w.�P��T��-3�t�2T$ư}٤�U���n?�[.��ٛu!Q�N���Xp	�v�4�4�X����v2.p����e2����g^��K�C(��@�Yv�Ҡ2�Y�(���s,)̓�t/+���f=˾>V�3
��+ӓ����)i�TϢ�'Y�]��;:�{�'���>��K�$�B{�K/[�>��m��\P�yuk:^ܭ�q�^߼e6U�կ'i��&1466ƭ�TkKJT�e�Q,���"��eV���h�i�FEF[[eUE�kj�ikX�Z�R�E�U�kAkVԶV�J�h��E"�
�l����h++E��Q�X)PF*ҕ���Z�0	iQbT�����E)kQ�-F�(�R�[eX��UZ֠*�imV�Q��DQ�kUE`�1��P��*�X���T����jت����*Q�,��+V�Xն�m)Z4�K[h�Q�T+kjV��[%+K��EE�b֣m-��b�ڣj��ePP��R�ċV"#�aF%h�km�QV��((��[m(ѵ�@�R��V�ZU��A��ģE��mB��4J��Jլ�[h��
�$���-�U���kR-m�`�V�Z,-�6�Ke���Ɣ��JYUU*���U	kV6��jT��ʕ)h�Q�FҫZʔX�b"��ajP���F�TKhڲ�Y@(l��}���q���坺��N�u�G��
f��D�d)�?���O�s�}o�F�>�b�����G9\ͻ��������?_D��5��^���8��4������B��;g��+v�{��6�7גH����	�����v:}"c��T�-O8-�F��'tS�1TFmn���t�h%d*�f�mՑ��쀬(���F��503�IP���q�tY�9����Yo*�V��c���gCL�(�y��Ԡܳs iㇻ�(��S�Ra�k2��18ۈ��}u��8�IU��ۺ���b�T����v��CZ:�גI�mgy�8�;�ֺs\8��n��T,W�K�[�y(��w|T9܏kuY1e8��+g�mv#�{�{�l�`S>p�"ܖn˞p/Q�,.�pt�5��ͭ����Y	]��Ͻۡ)�/�;>��U+�0�x�p �<�8�.������jϭ�����S�Н�{�>�L���L�3^��n�!��?]Vk�㫚�����u���u�V�Ş$�m��9��`����.�s�l)��F4�Gq���Tn�t_Q����,͊�sAҹ)�I3�d��d{'��7n^�<�z��EH�n�L����Ja2x���=�ҷH��⼹����-�.U]=�vٝ���L=xc���Jԭk�f�&"�V+=���9�+m��U䡴��*��8y^��<c�]�M]^��^Ÿ3f�q�m3Cˮ"����Ph��V�f�៵��_�!���*��,����
b�+�����@:x{>��z�x��:�n�O���|��d��C�P!JS���H��j���gCw�����ޖ�DJn�Pn�����v65vܽЦ��x�;W����������r]��S���P�B�}�,ڵ=���Ϊ�oScq���]�6-V�S{�>� Hs���0$�`Uq
�q�:j��Y��yl�sڊ�{������|qF;t̓�b��"�s�Fȑ8��4P4���r�ع1��E���&�T1�7�^���|c˱�E`uKa��*#�hB}��Y�6�Í��ck*75�IR�Xx�E[�E�J���q��єV�q��ȥ�*�a`���EK.����bߝ_���Cύ[3=,�_Sp0Ҏ#���;�݄k��B/b�d��-���c��}�1���$lq�Y�3��U�ӥ��i���J,ا#T"�j�wZ
�HW�����/�Ʉ�畘��S�����F��������I/&;�D�ֲ!Ɣy�r*hw;;6.u	��(*\�	�)O�|^�s�lI��T�����_n�FN@5٢'��d���r'�pokT�g�����	>��N\�1(��U�<j�Ȱ��Ѫ �r�T�+!Y{���v��#�G;|k'�L�Z<��˖��m��b�S"s����ƛx^��)�Q�q���wgcSъ���}א��ο>�]�g��t��O�&��PW���=��Kj֧Gم?,��~���l�pg�|�\UJ+F�#�1Ǥ���	��&ȧ�|WR���p`�Ƚ+^<�Ӯ��X�}Z�M�]ǣE_XDV�Sp�]VX�e�>{(����f�h�gf���j3-Z��d�#AD0�4�ㅀT���C�:�fH@��,Zt��1m:|�'i���h����s[Mи��:g�#\P+X]{2��c:б����%']�z	�)Yc����=��+}b��"�H�4,�;��{��~�l4k���g3���,�wӳG�n7^w�N���|��֫:%F=4#��60�uIe�*X�8�;��5�4�.+;B��m�n�2���˧f9��aP��N�^��6[���u��VƱ��*c%�p��xoC��O��:�bv�:��e��3�N��Y��2v����\P�XyX�����U���M�iMr�:�L�i{�|'��>�d�y ������D�[V�2�u�W����ꦟ��ӧ�nQQ�#�Y[q)E�p��x˅z�W��2��6����͕��dV7qc.ˉ��J�J�6%4$h��dJx�zE֭�`jq�(�{�;Q�U�dϣ/2�OnTN�K������X��Q0�"����>t����5��gЮg^�v}�Jj*�MlXކY��α&�ԫ�y�,����&�H�.�>pXDX�Aj'�88V헉B�%�!�qVW��v��lR�cZ�F��~3A�5�
0Ȝ���^��X}W�v+����v�Мg���Չg��yx{�� o��b|�=γ-6�\�ú��o,�=��D�O�dr��H���Y���Ug����TN{��-��"o4��l�'I���H�jF����*4�BhZ����.�/��-�욯'L#"���r�䝪\�}��	@����R���(Ș!]M��c�dׯ;�r�p-��K�b��K�={��f.��)Ϝ>�r�����)A%��H�8p�u^�7j���w�:��Ê[@���V'C���גӓ��:�@����3�1�,�zK&Q�qnhn�-�a�5���f�u�^"Q��[�nW4p�Ϲ�`���V_ZC@�T��Z4���\���^����8�N!6�jڑw�+��W���ۡ �8��0��Xk����ya�Td:*�K�7#�J��j�݌���=3�q�La�af�媬.����y���\v����VVy�h>��*��͉5mVDW����ˤv%�PSҥ�o�ܷX�"�(�z�� �C��;�7ޙL@�.�7��ˣ��
.]�GF��DgaI��R�B��g�(��K���z��A��:Ɣ��E[��z����^Kގ�`S�/ચ�u�ׁҥG�*f�hy?\h���е5�:y���{�`]���`s<Du�h��>��:`!��q�^�!���;u�Tzf����\nsT&�i�{4:�n��p; +Q#�(:Q�tr`0gԕ���^���s�a��H�Ģ�������l�(�u���Sa�f���G�ѧ��(����М���o��Sat9��J���t�&�����y~��b��W��W"6��sZ;+�Y�����ν�f�*�~�!�������<*��>�xSq�b�?z���(|�+8�>�]o���ߞ�^�=����U)�H�y}tZcݫ���w�hB��i��ĵ<��KF�7�w'w�k���H��-���)֧d�B�	�N+�:Ɲ��@�H�ZD)m3D�}��T�N�ڷ9V�k#{��K�7e�ݝ�_�����I�1����?k�U'�E�v\�z�U�k����+���߲:����^w!&�K���>R\�!����5^z�B�<�/��\M �Ř�̜�ѩ�'�4�2(CB��.q2Wk�0Oڏ��E�0Oj"���>����M�@����̮uΏe�[�t�D�=<�_w��%Љ�WS��igҧH�艸n+�qV$Dͷ�5�[��1�Ն���,f���[�`�ˮ"�v����-b9�epes�yc�MN�N�|�`ި~ő~���<E���q�@=P�y��;��ȿ8�4m�P�7�s������Z�z����0����MP�^ʾ��g�z�/!�-�q�ȭ,U7�q)��ؑ��ul7�����Y�VQP��/Y�SZ�.�Y?p��wtw��s
�а�_.�JY�t>�MH����dN�q�8hp�Q^�[�U�*�UǢ<l��j�֍=Xa�j�
=ɾ�q�;t̓�b��!��#����1%a�}y=�z>�7Ƕ��_on�JR�q��n��n��M�_k����c-*r�_���#�߷���h<
��N5��6t��t�X^3f.�5���PL!r��������Ә+��Dw�()���Y]��j>3X$dw�5G�3�߫꽗86yku~�1j>�6ܽ*l�_�ភ�74�(��W�\����u|�v���k[~@��R���B*�"*�iGT.�ph�+\���g��p�fA��N�G35�Gm���0�􎞐8�!��T���ȵB���|��s���x�F�hS��\td���E��eAjD2L�K(̓ӥ��8�l�Fb��d�#�L��֢1����o����ՙ�$��j��<�]I"=Y(��{���z�mg�,�b���09�/��KW�7C��L�4������XP.51<6��׹���T�-d�E���i��%�v7L݁2���	�:��!��yB�&�"f�Vr��7V��N�S�#�0~��Bk��/�z���I{a;&|����h���=����Z��"w/�m��P�FX���ocs'�>�vcz���U�2dK�@�F,�[6�,۩�&p!|Ok��v�X���J+Є|
+��S�k1X�y���{�-���E_�LU�4��u��ڏ^�3i�<��>�6�:}�p�s]lA7:a��xӺ�s{�];�{.����W�=��������PZVJ'V[�9Q7NU�i�v��K��`�U��DGʊ���CW�3ݝC�>L^U��H�h(֕Hl�9���*#e*�D�v���lX�W�S�sv�=Nt��{5�5a���3�5�xLV-��^/��[d+M�l5��	��9���`�Uf�`MWj��F�7��Ud�V������7�����ơ��ż�2�:gC�ƪ�"��N��|��֫:%F��&�z�P���~.������N��p�>TU�J"�p)_�Ф�u�9r�2F��䫦y�#`һ�O�>e=�q"�P?=�����f�zO��(��еi�e_�R8���8�;hf�%׆���Dd0��h�bx�#D��2Q�,ek��պ�jq��G��ѬT�ueZ-_$�U)�T-E���B��D8��ʇ��<�*����H��ѩ��
���5��j����g3�5��Ӱ�Y���I����x�`/�ǅ"}BD�v8,*z�5��Ǔ��ü�f�tK
GqN�'�a8�6*�ZŨ׿<��|k����Z��k�Yn�7��X[�yB��Ҝ`HF��.U���^�2�k���e���o^��X.�L��p��40�(M�#�������ɷ��>�u���w+��33�9S�Os������A�У#��K�pR���U���n��0�Ȏo}eP4����/C|�[b���L��Z��b�"g-�Wq����`��o��
ӿL��$�`��U����$�Qk��}�ߪ�2�>;D�V`x+���fF���E8v�	q�D8;צ����.$_:V��������3{��4���ꪌ���e[9t�Hɚ�p�<Y�a�"f�
f�0�"`<�u6s�'o;�4�@/,�u#�5#ː��Bu3&�hV�7�i��*��n��@�`��%����a�梩Y��[�^�prb�4�؆��rBL���;���XK�?%YK<Z8E+�����M6�k����5x���z��T�q�pﲬ����ȭk6$���Ȋ.F����6�<����֥�+�q #&0�ƅ�S�t���S��f�o�i��DI���ގ��"3�kS�u/y�f�0���RkaJQ�<*���TG?R���]z�����wd#5K±��v��Ob
�B���\ec��3l,���bc��P8�4��-8�+�VɩՕ3V���6+��m#���S<Dsni����jV\|w�PxE	�3�ڭ��b�	�-PNI+U�%��H؆�����/r�^r�Jtm9(^�a���50�����T�Kv��|��>2fA��2��4]�L=���U�s��7�{m����Λ+W0徣8��Im`q���x���������G7��jb��w�7���&�Pƍ�ۼ"��
��GD!Ў���S���o���i�B��R��Bf�61�3a]y�6a����g��[�n`Xiލ=F2�s��Z3����p9N�R������8�I�����/�@'[�Q'@���E%bf�8{Ft��ݹ�v�Gz�`����ԧB��(gM�7�QW�w�X�[��*���cv���ʾi��yja�P HBY�RHFA��T*OD��F��Q�9t��$��4�D��%U7�LL��`N��s��n|F�.O��F&@z+i5x�C`U孻��ա5�������K��J,�"*��)3k�0N��b��q��Q��H���V�ka���vy;G�g�ޛ���>�0 �E��w��%���9��ꊳ��Cmw� �uI�9��N)9NK'�uD��k�qŸ�%�Mm-�0^T��j�����w;�9VR�[gU�\絵�\�4�3
j��&�j��˶㎃�~ί!I�ȷ�&�����ޫ��Wf�S쮅TTI�u6���K�wC펩�0�!D^>~��p��Jɳ3���Br�{��O)B��˦�Y�ftH��Lqvu	ڽ}��Z�إ��>�nn�,���j�7K�Ov:�d�o'9$|�<��}�$�f��R�j�5Ӷ�޳�)�@q�'7(��AQ��B�K�E�j����ȹ��Y�<��)v-�R�	m��\�b��N�}�f�?IϷ27Z���p�G��5�T/����w�P����a��+�"��sB=ԡֲXnȶ�qLr�,ﳩٯ9w�ֲ����M��>��G4{6�q�|��q���q��h��ֽ"j�ʾQ�F��;�̫u"�N��SU�m��]B�;�{��۩��f��gL�O#�S�B�����z^��}��1��Y���u\��sSK�m�fWA�)���kNw.�uU��d�E�F�����Է�#���K��I������9�1-�+<�ͮ�I�G̸���yzj�^8��Ľ�Nb�v�k�v�n<H79Y��w�J�D��N�e"�/�{�;/J�?������� ��.����lv��Z:tQl׵{�q���]�@�����f�U�^HT�nJ�5��f>[��Wka��o�1��5u�;E��Ϋ1��/��#5h,5)����W7�W����}�ӻ��)h��/-�d�Z��#=w���'-�˥���ot\��oK	�UA]��󍨹��ʚt^�=�<{�y�T��{$P彪=X�ں�rh�6�T�1�{]˞<�V$��;X�l�o�WY��PM�x1���K�7Q���|���9L% �,�J2�_f�w9%]h6��������V�*�z�9i��=�p�1!�O��3>�KsVV㤑-es��Y��P���,,hVʼ�	�c޼݉_�^y+�@d��1R&��j�6��Cx/PDc�5oFr��6V+��o�2�?)���(F��x��H�&�u���|䦳��Gr�[�3����ɣ�ޯD��pV.�4�V��l���@�U�����CS^���L��1׶�v�
.P#L<��&ݣ/�p��ȯ+g�ب ��O�'UچC'�xw1V�$���S�H�J���擸�"�5��i��G6�F�Z�v/��2n��u�桊�7����e>[�S�g�3��q5�|�7&r��t�X�B7si��j��ˡ\�&�;I#�=�˝�y�В͉2�M��w=(����N�W�S�
䄵�4�4'�&ҽ�z�Kx$�QbzН2�r=@���]��W��]`h9ά�Uѩ���u`����28aǓ��ۉգ��������S������O�=��F嗎W��$m����
~5�L Xf�1t�J�C/-V��^�g�.�٬�s�sY�ae�Q�����6h~u����J*�o�y+�����ڨ�Z�W���P7f^^J�7q���e`���[T��R�Q�cJ,-��-J�Ғ���V-Z6���,�Z�Z�l�4��T���*��Y[iP���X�)klbֲ�X���B�iT���E�V
����R�B�X�+"��-mb�0�T��Q������J%,�Z�D
�֖��B�PA�U�E��kk+*R��R�**�%��U�Ym�dV���+m�V�R���P�FQ+
�B�eJU[Z�YP�jJʋ(�dU�B�"JԊTE�l����%XV�,�����Z�V�Q�eV�V
TR[V�Km�-k
�R�k%kZ���P��Ь�!cPF�eU
�V����і�)V��F�AJ�dD��B��J��*�(X��*�TmJ���-���"��V�)hڌ��լ*�-Te�IU��DVƊ���m�T��J���ZS� -�Y�+�o-<c���躞O�3�K~>/��8�N�����e���K5XP<�5	��D{n�~ �fmk���pg�ޯ9�8����d��)
����?�<�4��v�̕�'��
AO=�}�Dⲡԗ�?}d���g}�J�_Y��|۳�i���sʅ1G��A����8�i���w��|���f��CH���8�Sl����{E&:x��bz�3���䟍٦�Vm���oD|�Sg��iU'�T���_o�+�T-gY�8���Q��#�}�XzϹM}HVg;�:Φ�7�{�q<C��������i>ON� �d�]��a��CϨ���,��z�"�L*w�O&��|�G�p+�Ņ<��k4��k��}�I���
�졤��%E� �f (�2q:w�4u���=��}�+.{�sT��9��|��4����|Ɏ3v�� ���S{�@��\�c�����쟯�ԭ� 2 �ʒ���H��o��i��P�O=�&����ՇPyqiR��~�ɤ�6����
���w�i�O�v��3��+�&�M3��d�g̕��e��W�M`���˔e��<	D�QqYP�%�t��T+<<�C����f���m�aQ`l���m�a��C}`g�a��!�ea�%C���ܛz�Ɉ���%v��$�v���y�]��ƾ�_ �}��Y�C���aY�h�Q� ����U'��)4θ�S\�k��a����m�Y�Ă�{�xÉ�|�E��$�x��1�����z���Ay�F]�K�_g�>�1� |�����<ݓ���,6¦r��f�q
��.Z,��a�
��"�����&�XiE�ɣ;�N T�Ce�Z��/)
�?}��;�##�$�gʇlW���O?�v�13���$�ĜK�|Ѥ���:��{���*A�;���wa�<��u6��ViXxr鬕��8QI��Cީ2��'ua��1�Hxo�jq� �H�na��fN�d��wK���N&�+�̨i>d���=;�6ì+�O{Mm�q��O�܇<��S�;�x��b�9��HV�Wg(��i �"�3�
�O��A�	#H�6��ɜ�Eg�m��HܲT�f}ꛩ���ޫ�v��_+��\`��G��]&�J���I�6I^eh�����L�D�5�=�bU�6� �'4T��e3V��]��J���D�L1�����),��<���/v_C���XF�oV$�ߦ�N.�E�����sͻ��Ͻ��_�H6�L1?[6 bT?��O��&2y�b�$�ޠs��*�d�~��� ����3,�6�Y���4����]~����q�Qa��+|��㮾���W	N��_�_D>�$�>�@��>&!�ɫ�����N!���'�}�E�'Xb��ٴ�B���1=�aXi�N���w!�J�d�;�\���:�ۆ����w���>����'��wd5s'�z� �L�>X���&�s�ud���!]�P���u1���1����M���R
c&��m��
�w~�$�<a��b��&�<JΫ/l�Y*,;��wu�����r��0e�A#�p�YH�����̚Շ��riY4~��8�P�مd���f3�1=d띰�va�
�d���h� ��%|�����QH)����I�'��u��ش�r+�Q���w~b��3 xA�d�|9�����a�|����E~�i6��14��;̞$l1TY��T����N�c��Cԕ���i=B���}�vB��²�����~ܳ�o�q�Q@�'�}��@�������m<@�<g�>��o�B���g��x��|����`Vx��bB���AM��bz��!���
ŋ18�<����u
�9g���ӑ�6,��~�R� H'�O�N�y���B���d5�,�q�����h%z�Q���u�h
/S���m<@�?s�h9��^P?N�����I��c쿲g�1�57E1��Ue�ˮ�i=K#��?о���o�����е���������'SHJ�>{�M<d��ny��)+�C������'uN�ΰ��XwV՜d�N2z�~@�s	��ޣ*=�?c,�S��
�����rM��q�yG��Ag�5M5��QH.����'U����B����04�0�c����<gP�u�E=�SL�N3�߲�������'� Fm������t^^s����=I^'�Lg2�Cĕ��t;܇�8�f0��V0��,?#�Agۚ�4�����`i>@�1�3�Xq��!]�}��8�0�6���y��=a��:�	.�xk�S?o��n|�`�QZ4W�Fد����W����ŏ,bi�������f�{=�DTQҺ'�f�*��r��x��y�6kv��oi��#�m�a�{\���y, �tuE����=�w�ɗqY��RV]0�a`c9�T7g^G;�cg�=� &��H'����E����LC���m�<N���:�I������i�a����@ĜB�f���N8��Xb��d�5�q��[�$�m8�Y�}�D8wFbwrk����q�#�y�0�)>O��AgRu�Ù���H)�o��|`�B�nw�5���5��J��S�9UI��
�S,1:�J�ٴ��>d�I�`��T�J��U�؟����|=���z��	�?d8�������~d�a�0��O�������8�?Xi��CSd�$��_QI�I��VOX|�������ts�U��Y����q�"�i�����H��bo^�|�����: ~=��H~I^�Y3Ӽ�!ĕ�۝�T�!Y�}��{�B���������A|=�:�X
����ﹷ��{泚?g}�����E'*L�;�tÌ/�8³��gSH�����M$��ܚC��1!����IX�i��N}�SI:�g�S��r$f�w
����:��k���|�{�z]w�����m�<�Lq����XmĮ�xeY�%@��1�����C�Y=e���4°�Ry�:�H,�O|���'�T���l�t�z�@)���'��#6|>�7n�Oտ~|k��
���s��uRW��풦�I\C��$Y��ՇT%x[�g+5�&'Y=q8��t4��*z��n�HVa_�{����i��31c/��co7�Wօ|M:d�1��s&��Q'6w��8�ꐩ����Cl��i�<;܆��?!��Y���f0��T:�$Y��Xiq�`�Ԩz��N��h�@�=~פ��G�EI�9���c}�|�gC���<��
�o���g�8�XNs4�Y+W���M T?����/�Og9�l<gɌ4;�x�Y�LM�QI�4�{B}D#��{�L���Kޫ�˾���;9�%b�� |�'�+;�ԛH,7���6��|���
�{E��;��Xmį���6�?2T�;��2~LM�xw�m'�~�&�wO;� Y���3 e�n����/떸M�Y=���˛o��U�F��ތ�[�]Cs����F$ǖ^"9�_]�M��<f��ִ�=��h�p.��V�۰�mN]aGF���.�����Qc��F�o��t�m�����H�q�&M��w.�BU�Rni�&lKv?x��:�����	F��O����]$�TR��O\`�B���g��0�y�C>J��5�g%z�S����:�J�/�uH:���;�=�� y���i�ϙ+�������%
�~���F�zL�D}�G���*b;b��B����]5�}��
l��ɧl��(xj��
$��ɤ:��Hxf9*�a�Ŀ��3�c:��E ���k>.���r�<jI��j���$"�$���x�?0����q6��+��;��(�P��4�h��+��M�B�����L�#�������.��)>B��
��g]����{�-�wK�;�4����;���,1��x����Af�|��|�u
�AM�纇��=N!�=���X��y;�<@�T��vO(�d��4e����>�xH<���.�| bS�eudus����TqS֌����O�������/�N�'X{~ɤ�!ܲq=;�m!Xm�r�����>O���$�*,�N�E>d���<9���&3��a�J��Պc?*H?z3����+�Ko!�k�U��<	?"�����A�7�2Nya�'�����C�f�y�3h
)�O�|�{�I8�N'�;��HV&��&ߙ=�4��w��u��2k(����� �M��,����3�����.ޕ��$��ė�&3qP������ͳ�1��E �f���~C�b���Xu�"�0�y�|�C��y�}Ԟ (��o�����I�y�b�2dԏ9!,�T�i����ů�'
b��q��i���Lg�Jɩj���>@ֵ���8��n��g��5ܝM�x��y���
�C߳���C��1��&�d�Y�m��"�"����j��;t�y�0�3|�b��wl6�ꁈx^��1 �5�L8 c���Y*,�%E"�������n�I*e�G���)
��s	�u1 ���eI�%E�y�?�?g�Y������a��'`�Nn�H<�m3���� u+=�܆�l�RWL<�p�)*(q1�:�$�����8¡��M$=�q�L��(�Y0���q��*�����l��B���X���l3pe���#ؽ�̡�&�^�+���wb�����b2WCA�[�e'���*�뮖��ɛ�&¯�Ҵ��Ҍ�wz ����wtK�'6ʇ\7�ۺ����)��IB��Z�_un�������J�Fu=U����e� ~����7�i��Y����'r��AN Q6gp8������^�4��B�w�4�Y�i�
�AJ�����z�Ę�ՇXb,��~a۔�5X��	��FjIl���A����1Eo�h�|x��<}��ɶq���@��eaXVi�Q�s�ed�=>�M*��
�a�ɤ�g�0�}���٤�o�,�i �d.��&�(M����w�߻���Ċ q�t�bi���=N!���3�%b�y�a�R������,�����0�
��C��~Ci�Sú�u�1�d��s���%E�I�y�@Q<}�"Hɸ�q<��jj3��u��i6��ð��3��a���R~N�$75�?$��O��Y1<d�6y��*A����|����>J�Y4��*J�;����S��;CO_ I�W)��|is�6��{R2{��>�j�l+ӽ�=M�2٧����V���N�T��������!S�?0����SL=7a���]�ny��R
z��϶h�VT:��g���6ê�gX���{�7�{�����ᤩ�3��w�<gXTR��6�0�=C��m#�Xb,��}���c�]5<d����Lt���gY7��?�L?0��'���Y�%Itat����ӂ�wf�7t�̖=D�G�B����rI�:���i������VgI���C������w�O~f!��;�)�%b�7E6�H�C�P��,���T�X(�A}��E��-P������R,E�o����k�I�*A�;?fI�aP���o*,���4����~�GP*OP�S���5�B�o��I�|�����>I�4��D4�2c�Q~B�Ԕ��8[���>׆����=�t��q�B>#�H��(�,�3����rM"�S��ǌ8�2~~ɯ,�'ua�?K���R��ed��q���|N T�}��m8�����0����4�|f��|����?���.s�ݼ�5�=f�+�t厨��&����eC�K˰݁�T+4ẏi��;CL�
���٤�8��6�<���,:�N�V@�T8��ɷ�����S�S�{rm}���pt�N�.TUGJ�̲T+V�uq������, �;=��it�[�x:-�J��̧2]>i���v�8(�D6�;���z]p^��9�!�z�]iT�-�X�u�)Yܞ4����'�F��^��y�p�zv8�쥟����d��*ަ�:?iH��@��P�����Y�C�[a�
�CG*���d��U'��,�M3�0Ѯd5�B��ny�a�u1 �{�xÉ�|�E�ݓl?2H��}-�R�U����}�Ml|��%N��i�La�J����g��b�H��
��-�I�+��Y?8��=5H�=d����� (��4gp��
�hl�kS�}�^MÝ�`}��O�g��g�Ϗ?R|�&$����8�O�7�H)���>��P��<���񇻰Ğ�M m+4�>��Y*)2p���8�!�Re��N�É�� "������p72��7�3d)�{8�PS��$���a���i?2q��=�p���Y=�5�<�Ag+�ٮ�9���!��Г�eC�y�7�B��B�E�S1� �(���H�>`��+d;�>������%g�1=C�i�A��bt<̟0���	���&2}j�$�� |s�4J�gY<ϰ�w��u�g�浓��AgX=� *�*��P��,�a�>��`t��g#t�{������B�Ǽ��a��L@ީ��&!�
��Ձ�Xz�CS|Èm �ɳϷ����@���i:�g��bzw0�,4§Y���<IP��9ܚ�O\a��~>�3��~�g>�Z��J��ߛ& (���S�I���ud����q0�?'S�vLg�?8��i���Ow�u�� ���ɴ����8� "�'�9��tc�g6�����J���sI�RW�C�����̚Շ��!P6��_�rβT5�aY=q8�Y��=CI�'\퇻��XW�&�}�?2W���jO�#��eF3;��Q���O��خ��{��*'�Pה�a��m�a�1 �_�m�!�z¢�Rbi����{�6�|��9��ΰ����RW�u�{5f"��+��<ݛG���{jN�_]�b�b٭��n��
��
����C�|�|�C��@URq6~�i�I�>q�9�0�ԅC��gSl?3�bO���0�����}��Sl1���(��i �B��>���[����>�x�ގ8#�`=���������r���3G~��r�퍨v�[,�E5}Q纃��6����ì,���mؚtO=9��"�L�l������BW\<�<o%o����$������ͬvt�����[��Kk�]~��&�w��Y�}�����Z[���G��c��.� H��
��p$�
����N8��s��ҽd����u�h
/S���m<@�?s�h9��^P?�a���I���`V|�C�o�߶��wx;���{�W��"�Sht勦���h�Ý���t�&�6��|=�&��TY7<̊u��!���wg;�zw�:�h�a���ݝd�ִ)�O\O�㟿|w[��(�v��҈χ�����Q���¸ó�<��>a�SMd��R�/�qYP���HVw�`i�a���\f��1�aQN_�
�gXbq���4�wa������N�������7������g�*ӿoz����Lg���i=I\3���q
�a�9��>a_ڢ��:�}�d�@URgy�����l��a���vy���xì�bϳ�Ȼ����Ĳ��h�|=��|@G�	�j)6é�{�!��1 �Ow!�,�:�w,�i'�Vk�>�̛@QaXh氿P1'��Փ=���}ἆ�6��&�k�d�
.�{=I�ƙ�ό��g�g1$j����!�+:r���'YwI��p6���O����<H,�N��9��QH)�o��|`�B�w�ghLa��\@�TJ��U&?2TXk,1:�JY�gk����cy���m\��#���2w<ޡ�
��Vy�Nj�2V�f"�d���O���!S�N���,0��~g�;���� �����v��Q`yˉ�
$�eN"��<��Ʉ���!~��^��u�$����rc'f��Vqg�*oY��?0�޽��H>Xyy��,�
��ߜ4���u�=;��P�J���]�*O���6k����>g{M3l=G(�%�׃������u��AD[}� UϨ���I��E�X_��]0���ì�bi���b�~��)6�wܚC��1!��rJ���g�H^jG�G��[���uK'��My�#�l���Q��%�GaY���|�L��⯼�;�x>�U�o�����w���zB����.�9fv���tGL(]4x���7���s(8
ʉk�N�����s�Puq;�z���C�(Į�����RW^�(�6�����=׭Y+�ˡ�c�/:KoT�)�b��]sm��1C,�1��۴+U����T��;��=� &�p���ȃЗ��5A�`�6HhЩ�(�Qـ���/B�^�Y˳W�g�%�M��7b�n������7HɤЭ�n+"tG�U�x�}J�Cx��J�쨣�@��+����Շ
��]�ڴ!(�]2$���yR;���XOP�����;�ż�辨s�w#}^�/����C(�+<�4�Bا�yho�v,6���{����=K�2���P�~�����q�sT�g�b9���^�z��n�./^Km*1,>��+nq��)�6�p�Mn�#���AJ.6i��IʙW
d���ɟrch5��XӁ�\ec��Rj0��R�f���`���I�}i̫ܵX3��`�,)�T;|hZ��S����x���v����8��!#�s����5cc1�QsF�����=6�I��۫#��
��GD!ЌGf�冝t���k[c8X��P���h���ͅu��m�E�p{]�]{��Ѯ��,ܦח���-���nR��D�Q5wK�/��`^�t�Uum�����h𜖎g��~��xV�;a�+"G�ƎEJ�W������0�N���}BL�Thb�)YN���y�+�daԌs�t;Q�����b��|d��wFZf������_}�}_b�tι�t�~O��%�;��~&�uj��t�&�W������blҵf	y�ʟ��&���E�|lz�y�F�C2zfK�U��دKt.�T�3����ױAV��tw�n��� Z�퐴[�Q��}K�fৼ!B��Z���8T*OD�J7`����K�NF1vu1ۜ��!���c�
��g�:�m����D�2��58U�Q�SC'r��;��g���Uvk���+��
qa���4+��)�B�)�m,�߼G��`��ǚ1�#ޙo�����W�n/z]�~�I�!8'9Ϭ�;*r!#�^n��O!*�#6K[y��ы5�|GijKjVͺN��{6h���bܳ^]qv&�u:o���&/��Ik�N�-}�>�-��nős�yT�i0�o���;U[=�qb�F`�.������Z㈗sG�}�D'^�඗��|5jۋ��_�����=LA��Ԛ��s��1�5<E+ݣ��t�6�'���&�ӂ%�zϲ����'����'M^Q�r���#�yf��n��f��!W����b�'�M�`�����#=y��]�p�-�'`iN�ػzѝ��1�����s6I${n�M9�0�t6lX"�D�1�Rɸ�	<�S f�2���a=�Wd��^*NC�r��k}�A-ú� =�VlP�P�9��g�6g�孫P�k�m� i����dN����
�5�JV�	�88�f՞׍rܰ���d*��2�C#ɭ�mCv�1N(��tI���{����)ood��p��,��LJE��d;�r��Q^|g��R�-�y��*\'�=��-��g��n�,W���#�=0���E9D/_M(��nh(%�S^Y�f<��'��H����,ڌ]t��bW�)R=P%��T�}M��J8����R�|�n���gޞ���l8O{c�o슘2�(Њ���J��GT�ڨ�@�o��rX2�n\�cA�e,Y֜i��Y�r5E�8B�]�E�bufE�'����O9W,O+��#����u���T�0WB43�ꇍ�/��xKW��`1^�L�4D-F�l��0��6>�](n� B��fPgDn+��~�;k���17L݉�a����������T�oc�(�UJ>z�BB�Eb#
��:N������8���^�N�� ��������@���4��Z�N��)�TΔ[��SFV
/��Wb(�L�-v'}
������&�a@�t�{s�]p�2�L�r�R���9{��g=ӧԝ�Xb��b�{G��#��_�`��=����,��5��]u5���-�kqf�W��on�]�%Ƴ)v�'��ٶ-��L�;	�z(tuG��t��o/_q��'t��X�SС����;�1���`#����#���(�v̜��]�z�m%N��u�$�e��e�ʶk:� �K<�����oIz.	xĦ4���}��r�����M[T�T��UW^�jP��m��u�l�I���
<��-{{���i����U-Bk�����h|g�0.�}�$���$��LB�S��j^��)�KJn���>��aI�����Z6�0.�h�no+";̂�NQ�n��\^{.YGh�׾wcmc�t�x�l�+�CbY�gΰ��X�B��$uxY�%�[[�Y`�\q>;���gz���r.�v��{����T��NcNj�h���}�ʲ��Ϥ���a�V�>j��5�`���)�Օ�,@8+VKڻ5م��ϜȎ9=�&e�7�)!���WǞܨ��ʾñ�͌N�W@o���)c�w���4n-L7�+��ܒ��3r�{���V��UԬ�#1᠓\K��y�Ĝ}���"oOp:��-Ғb�I�o�/(������O�T)������]�Q��r靻�2ZBX��+���흕�#�C*N�q>�<����B�Q��z`�/`�9ֳ3EIMV6:툧���ו��2J�n���/�E�S�aS�=Ν�Θ���k��`�^m3�!屖��=�*O���f�q������g{X<;�;����tSY]oh��f�Xg Ί=���� �4�n���	J��DR�������c�qX�L�V���âV&�O*r���%9�[6]��ˑ�"*�][��t�����'��.�3��B9�rwC^�Y�����o��a�p=.g��]J�M�)����Bh�Y�ecJ��!PN#nV᧽�4�̧�ֈ��>$����u�Z�!@�w�k��/|��;'���y�����>Vs�K�?.g�ĭ���7��2(d�ZP�mf���;$wϗ?zQ�r/����Ą^��=���B}77�ӏ�DםA�zw�UI��n
�{��ۋ!�(�y�0��{���5�~�ut*�6Q��v����T�� �۠�sF��\5I�GҠHgV�ty�{QV����P��:�<�oh?r��21��<��_[���%��:��$]mB��7X��.���c�����:y��1��h�ܩ�q�'o@��Q&�A��5�֔��%ө�m��zS�N�_Tn�>ʜ�ahݽj��o���> �A'����(�V[FR�-R�X��m=əTmP��ڹ�e(�[m�QD�clYYYZ��iilU��Kf5�K(��aKh����2��(�j������V"�Ad*-����T�ejQ��J�TU�+RQ(ʋR���e�V�cq�Qb��VV���EKl��+m�%E�J�@F*
�Zʂ�b�*�%�,m�V�T[iKEd�T+ke�[+کR�%��Z�Um�b�U�mPQRص�*%h�!S�*ĭ+RR�X�Q+R�Y+iVV6֘�9`��+`*� [V���)kH�*�*�P��Z�ԑeJ�m
�AE�a$X��"�+�E��+���%BV*���"�mC-����	X�d����ԥ�X�aEP��/	���ƽ"7��*]�l�1g9˸�l�\t���OX�u�:P��vBUe��w �2�������܆��܉Y�����S�=u��2eh���0$��`�,�{��F�ӭq�����vcz��Cj.��豦�o3Ϙ���ő/e����ߜDh,�&���p�,��cIa݇[Wyyg5k��^���0SSe�n����ӄ[٭��j�EO�Ӡ댘iv����q��L��Ư%~�t߱�;z@H^՛�IN�ԫv<obK����KY�uDs��eL#�����9���U���I��ɔv%VY1��N��|��֫:%F3*����<��*^�V�7؏t�!#&���*�D�*�0R��)9m͐�:d������r%뀛���Q��bo-G��pus�Hi�U���Y�\JQz��3�0�m����T;JJ�iw�����[�F�8�f3z��'���GT����(��%�C��㫇ZFn�*NqC�B>��J w�[��Ze�>:��#R#��D�{Odj��ޠ��g��yH��Z5�+>�y���t����&��q/�x�L�A�������s�x�_;HL)/h��w̰� )�:�Ѡ�f��� ���z�,��gީ-�%��t��E�%馡�5Z�◘�EyXR�£�U�p����]9��Ѭn�[�7�s�Xj�=�t��U"�ʛIA÷J��Tw������a�oy��u�P�vQ��Dig:�N���Ǭ��3�n�R��nd�+��C_;p_=�x��|>�!�2�ղW��|=u�q�-�HF����Y���s��n1έ�K`��B J�O��=S'a�l�oOʰ�ǻP�G��g.��z� ���z�n�bw��iy��LXK�³���i��|�L��⯼�:�ׇ֫]W���1Krk��b�`��ɨ\�<��~,�0ё3|)4FW��Yz����Iw��7!(�&͎K��/^��|��C�2S�XϡxW���Cƕ�R�)��`��9�=$G^����z=��o���2RrBL���H�~�'��w��]2�>qj�2A�4'�T�]:.�z��Sq�h�����e7#>��)��fu�6`9�jەq�Yi��Ȇ*扢	��ʊ��W5Hqt���S�W4L���1F�E.�ݪ�h��V��W��2�����-OƭF�\K=b �R��e�юPSy�4(r+7z���Ɛ%b�=:'����.�c�vʈ��Yǎ�����D�k�)4����ܽ�ܑ͊{h�Y9���C��ȅā��i�m�[�ua;����U�wAF7�Q�E�3{a7[�$���ã>�3k\A��������q�m�*&r/���V�S��q�\e`}~3Rj0�
�jvi#s�d�����z����4��<�	P�>4-Zvϩ�tb�
g����`�:}"c��ǂ�owdn�2�e>K�����V�5jC5�!8xzm���N1�#�Ud0�v@H������+�pt4����E�D p��@�9��ѼYC��
�Ϣ�fQW��ȲŇs�;k*@w�{���p;5�8�~�*��+�P�*|k�ThΜp$ߕ�qw�y~��`��Q��O_WKu�L�DsRěnjDj�|4�̗��MlP��]�<E{:oa��ߤG\ɫ��k�RV�;�T��.ĺݏ[uY0�
�R���
���?�U��l�.Δ�6er�[Ր�UY����t��[l��`3m׈�).!��MM`�*/��<#��xm������R��fM[��8�<I4��܄EhV���b�hЩ��㏏W"���huu���P��t�3g�zE^ո����,BpO8������:l�\�Ô=5��2��ν�N�P$����I��o��n�u �s�e˖�˹����m)ed[˺ܫ��.���+��WI�.����*q#f]6 LS^��_f�MwHƖ��u7s�烳o�j���`v;�q���f�˩�J�6���  ɺS���j�bL}�ʙ��eũ-�U[6����ȗ�5�E�,�W\��ٝ���yv���֧v>����*O�Z��~�0���+���yv�q�z��v������������@�ɣanP�4U�:%��l��hN�ڙ:gmײ|>���Ø����}�xJ����.���w��vr��UKx�,���b�I�䫖��P�'/���G)���G��{��B�,ӆ��Ps��nob{Ϡ��(a�ɪM�^�>�����}����uL�V*�2�C�ɰ�����r,�>�w>#cT ^y�����L3k�J�=��# Ft,�����	F��6����E>3�^ƭ���<+��̜�y����k�Ag%M���.����~��AU��ߔ�_'2�������k5p)����`[˩�
{<mF9u�1����.vg�i��ri3D���竗�_i�7s{
�;��;��ꬨ�L.Q�I�� �G�<�����ܫx4F�['�k�7:�串uF�.���2aT�VZ��$���B����T5v���̴7��:�$�f�+پ�ŬC��u�\�)a�
����_>QX�y.�78��,s���K����wY���O�t�N�\)S�J�P��z1w�<��P[{�U6�aÿx���{��8R�*��Qi����T_�'VdZ�|�uCfv�\��b)VºY�c嗇�i��� VOQ�k��u�nYv���0���7C��L�-�5��#��l���.D1�t�c:�T
�,��Y-Ŏ�q���u��f�L�Cцb�q�ސǅ��d�ò�Vo��r��G��'Lj���Ot���zUi5��w�yǤ���=7�L�>�Ή�u�S�B�?@�+�@��6���/N���+�~���o|��n�A)�h\/�<��2�����,`�Y�P9Qa�����"�B5���N�uv(��`��Ev/�!7"��_��m��ߑ�KB�����m"~�aU:/�.�^b
f�����ϗfHF��#�3)�7��B�`ޠ�Ѯ�IW���p��I��E�>��DWUq���K��)���O�N�yU�3M�&��*���s�;�a>W�p��+�S�9�R�ۭ�dɫ#E���(���8j��#�=Ϭ�Ex\
W�)9���"��w��6`�C��A���N+d�D�\|���[�V�w9�o�����q>8�b�UeH��x��8�#Y�=O<�]��6W��q�eȽ�jג���	���L偭�3EР�f��]gW ��XEֈ������6��;Y{�7 �1�4�o�����L\�}�S�����C�Ӟ*酞��aP胱��d��^����M�g����r�Jg7:1�Y�j۰ʰ�� Y��V�X�<tH�#�L� 5<bX��&�K��Eev�&�^��N8y��(�ܝp��|��d)=�#��>��N������.z�bdq���f���5�yY�+���
4��=V$כ�Y^��F�/ћ�Ѱ��f�{����W��C%��=f?N�g*�E\;Ɲ�Ov�qƲ�,���U���ִ'�ȷ�3I��~�F��E�r��:[�jB7W�g�+ڤ���9ٱ
�!&��N�D�!#YT[�<;L�G�a�S��){!�;+��$a�jq�p+�L'~��V>o)���º?xQ�i����h8�r%h��s�Ձ�"�E�iS�|���T��j7D�y:`�64f���p0�`�|�{5��-��_�]���%����dмx�^r�p,5$�(7Hɠ�����؎>����c�VwE̬�n�5-�{�5�	�"<���2N�o;!���hB��mM�K�W�����
�dI�~�l���9�{K����ν*\�D�DnA��G���Z��
x��Z ��Kn+�м2GIo�f�kQ��<|�>�UN��Z�S�ΰ< ��}M��ك��,��꽆n�a��p�_�jЋ	N
�$h9�ע���NK�R]="��q���u2}R��})g�G9*������Sq�#�X�ڲ����P��G��/���^X���,GN������"O�B�D5_p�҂���9������&�C�ܱHڼ��Rs��i��P�����s�Bl��iH��p01�+0�wA�Jܼ
����݈�	�oa�sN7^��7��)�\e`�_�U4�ԏ�-NQ��s����
��ꌐ�@��tҴV�T7�E$�0�:1F)�":۴`׬t��H��%zhg{�\��:sT;�M(	�fR�vHN�	C$ӊƍ�����	Z��9��Tm-p����(Ԉ�Q�����Fz��61e3j�Ϣ�2��Cq�2UY�U��iQ�{��je����5���>,L����7O����a�7�HuK���=#a�L���M;�z����5CnGj��OL�p��S[�B����Vt�9/ )�+��۵!b����M�⭭
�:o����3"źC(�}sW��b"��{�wf
{�T�uf�Ô�8�Q�W~sϸlf�fi��4(�"�� [!U��Ҹ-u��2X��Z��<ޓ�����{RĘ[���ҵ3?>����ꦹ����4fGl|�d]Xw|T9܏hn�&.��aS�J��T>��e�ݾ������N��va���V�W�s�,.�p�
�����C��fۯ*K�d����苨Tfnp^^��K1!�_�](ɿ^*dp=*yt�N,7!PЬχ�P.���|�ͣw�-������h��a��&+�(�8p����Qy��y�L1	�/��ʱ*��d
Zzb3+=��շ�n�>��Mԥ��*ϼs�p�j�ߎ8��l�n1��/�-���7�]��{zV�,v]2*ۯlCF*LO�{�(�&�+��Z������΁6ٺ�����:y-v*5��	W����Xp+�h�{� �5^3�Y�'a���Rc���/k������{QG��:���`ޤ�dK�S�}Mҽ���^����4)7��%Eb�,fk�v�Y}|�-ۅ�lT�O�;s>㝳J��f�`��^s���s{��q6�H�b�C�����S��z�"E�Y�aW�\ld�2�'o��q�ۦo�1Z�+��e�\����ڮ��9ڧ�ޑ��Q�������c��&���^g���ni��6�rg^�=��eA��a���.C%��KO�/7�����\���l���WAo�w5¶änÎ���-�L�(F:�l�騅�0`x�I���ʾ�r/�U|  l�1��'J#�I{��Ex�#fD㎺�(�ή%(��6��*l�m�'����7��w��@��6�S�d�6��p.R�G�Có�r:.��W/8�&�ÞڙG竨v�~Z�g[��L�~�N W��P���4�0�\UPs4�R�y̥�W���{�,�+qW���E�",+��w��󍈃���7Y0e�Q
��ң�Pl7P�<c��Fm��W�_�����z�QF��Zq�6R�2�j�Np�~����ՙ��B}*yH��
����x����[*�I+%Pl#@g��eږ.5R������b�d�6�i^×{��`��Ｚ��x^ҙOHU���㏴��]F��3qb�m���wr�rf��\�L��W1|!��p�����D9O�t��8^�����.�'u����;%a���
EՆP��}��������ќb��wT�Q���%yM�)="Ȧ��Q�uYc �Yau���ߜDH��'!��p�ŗA�J��:�D��7�6{�B�Z(	��"�ٺ�E�+�D�ߑ!�R5'�.�)$���#V��7�o?=�OOjupr��f���;D�8ɚp�Qu4��71��h��O �ҥ��뫳]���J��#ᴁ�us�姷�i�ʮ�1kJ�&�ZW��� ���cW������m��_�h ]����� �t��lM_���B|Μ��ep9Aw4�;�����#>F�?[x%fW7�lX�ޠڳ}���6ջ�5��@����g+�֞������&��Q�tTCb�*�q#Ӓ��^�M�5H(�*�ȼ�^w�N�ckM^י�#��؊��㫂�z���Bn�z焄d��n.�h�ȖE��J�v��!ʇ��jR���k����o��c����ã�Z�O��8���$4�23�Q��[�5�s��ob���H~,ʇ~�V�ʷT�8q�g*��p��U����7����'@���Z}��E�qg5jݺ�jq��G�Վ�@��t-Ç8e��'�u�P�wOr�ث����lG�`D�>����;uƛ�ϡ^}���>���bM��K��Rǜ�Mg_:aV#�B"b4�T+��h�F�hgH}jGqW�Ǔ��O^Y��vo>,_]t�o����6PBx��|��}�Xс{
q�-r��0��Ԅn�&+yE��W��.�%�Qm�`�u'm��q��{q^�'��u/�Q�e���y{���N+;h��ãzf)�9jU3fv��dn��;�@�W���9�*D ����b���Q�z������:���ʛل=��=Tv���M򃢭�)|��8<$�P��؝�����T�&c�.	�܋C��?�x�]|<&��hu*=�u��(�ڱ��U��2_[�d��d�<�+��;�eұ����$�1e`��:t	ֺ�u��y�����H��e��V��,���P�I����\G}޽�n�N���i���ʢ�G{k��཈ 蝦�s̬���6lۓ�}�ӘAy!���~�ii���oM�z��NkRo@o��g�_�/N`�n'�r���7��`��ȊD�弜=��IR��DWn��Ѹ�Z�9�iF���\kq�d2P\1'�{+TF�&�!���՛%I|(j/��WQ4i��=J.��f�s���'������Z�ސ���<�Nγ�0�t�y�BNx��>���������(^(����i<Z�c�Sy-���IYF��M�^�N5��s�J�'�R�����ӻU�)��pn�5��j6n畉������>�9�4�.;��3Y�9��]�B��ݓY�Y8���7vH֭�ύ-�A!�JN�r��ݛ֟o��ͅ=�~[=��	W� k���n�}�ڌڢ��J)u�J�}��s�� Eu�l\���J�x���y{h�y�0�$�e�k�l�ȕ��om��u,���5]ڪ�78��d�uؗ#]�&�<� �i( �V��e`hy',[�F�f��vڧo8��4�Fr��$};�H�tٜ�4ˍ���f4�����6�Y4RC_n��٣�$"d]�vN)�1��Y��|5��u���!�K�xJ#�7g���+A�'���MI^�-o���%*T#���*�K;�z�����( ��ȫ��6��j�����e�G�X-a�"�!C��(�g"8�y�On{��S�l{/c᥄�jH�
4�9y����_����m�y�f��ڴo�(ݼ;�ڡ�Vy�vtw��/3K����r��έ�.ȑ��ZS��1,w��)X�;J�����4Z��r8p��}[�0b�<>����ꥬ5�5-4o���}�j4 UvV��+:̔	oM�\�d��HV�#w5��r�ޝ�Ki҆�wW.���.�ai�wd���u]:��0M9\����pӱ�2��U���G˻jȉ${N缷��������h�\�U�M�V!�9���w�:Ek{��Zk7 �қ��l�C��tNk��.�f�t�T�u)s;Dl}�)�j� ��E���&�Ƀ5�4Y�.R
�c�Y}K�dC̾6�'X�L��]�oz��}D_d��V�*��)X,"�Aq(��)YX�b�B��@��F[B��@��E*T���lY
ƍ��PAcl���VcʡR�jJ��j"��((T�0-��X�(��h��AdZ��j5+eeV��+RVT���
�#j��`�-@��6�TXT�U`�TЬ��Uj�j�mRm�Q*,��V�VV"B�(�X"KeDE%KlkH�E�l�3)�ed��X,UZ�F�V�DFQ���AF��Pb�m#lR�ŋ
��Ki+Z2�Z�
�T��j�J)����clY+[h�*�%�J��mTZ�I�ƾm	��w�,طQK�.�o5����XY�k]�N�K�r޼]\��z��9y�7_�XK�3v�!ٷ�蜃}3��1G{��������E;�Ӯ�� �^�C O��bP�~�i�G�a�S��/�{��r��][�U�q�F��U�~�VC6!�`��<�+���F�'��hx��J��ۚ��Vs��ɱ/�������̀�MB�nɤ僄o�6HhЩ�(��Fpܿ?F��f�Ag��9)]����)\d��b�|��ԒnQ���[Q~n����ek�p'A��ݶ�>���a��Å����U���5c6���
���[5�����7bV��`�o�.Y�xS��XK�Q�*�Y��Ҭ,ȻU꾪n8�Ç��+8k:.�:�P�v��pta}��X{Y�&�5Y��P�R
�k�Ȼ�<������%Rȣ.�g���ͤ�ƍ��)_����Hå���畦(&�׶M)�ӁbcKz�߬�\�ʻXb�|�j���A�yAؕ�N�M�n9�4�U�S���T��5¥���1d�,�%����ݣ�|)U3\4?�r��)��B�tϸ8ΌQ�g���7h��5�q�~D�'�A�9w���]�:�ub�y�� d[ޏ!�"�U��z۸d�Jr|SB��(��u����mwh�Q��Uu=l�ѼYC�c�;*|�,ds6�&��j�|{���Ot�.��::�w+#v6�$�ֽ������1џ_&������6�h�R��P뀜&M�X!�i�cF�Xm�uW(uqPpB�u�ˌ��ӡH�gx���F�F��L���/��x��쿽��{6�^�ޅ\������}����]�ΠT�Ə|c�j{5�~.�_O�ÜoƐ�}j���'y��B�*����lBpD���W"/�`B�G<`����^�z�/<w)����j������.�S�*���z۪ɀ�I��#� k��\ʔso�����r��r��U�at�;��!��K��e��J��Ef���`�>{f�1�_t��}ŉ�r��6mq�x����z���e��"+��狜��7Zif��J�i<A*�<*KQ�5E�*	�m}Nܾ��ɭ)9�G���G�@�Ӕ��t�7��^�>���y;*DBGj����R�@��*0�j����^l�n6���y|���L^�]�\�qA�K0^Ԣ+ n��=�*	�s���3������%Q�]�mu�f#�`�2/-M���p���	XO��ݮ�c�kf�����C����v���s]��o���nx�kq����+��A�m3-ْl:�V��bf��jsZ���yCҊOK���-�;�.r������~�c��q����[�Qk?x{����������W�.�uy
	�ȿ8�4o�r��G�[K�_چ��m�8a�l�eM��h��u���n���`�%�N��>��^�k�{k�+LR�q��ř����hs���7N#�V���/�9\j�}�/��������i�1V�����j ؙ���pmGsEh�YJjéE�t�!�m�b^�aK§P��o��p�J=xb�6�73�����*.VCs+�H���Ex�#fD㎺�(q�F��t�r����x��o���3���T�v��>L^+��:���<mE	�d������#(9~pPo�4Sh�J�s��m��ڎQ}�e~�N P{<mFyˮ�xq����ύ_�&�&ؙc*�N�w�ԁ�E[�/"�q�oa��#\�bz��;�0e�P�<6}���2HmWN�oy�
�%���f�N�o{��QEW���Z�麰���.^%�-
�t�Y���G����0w���$��Ϩ��g�t��;p������%z����M-������("<��>竟�J�c�;�cat�(�Wl��t�=��A"i�g m�~�Jo���<n{�~��{6��K��u�8�2Qc�ե����D$���nv�ۻYZw"�[�Oq�ƍ�4���,
.��-;�U������f��Ok$�~z��i �Q�B��}2���8��●��v`��ʽ��M�"�����a�L�C��d.us
1�p�QTi0r&��7�)ET��s�)�\�ror��Tv���Ӳj��!����dW�F}
��@�R�O�|s�sMƽ*-�����cx��}��"����᭚,(e��ju%�EdE}�r�}��xvk��`�*�/�3����]�21dlŝ~�v4�m��f�@��,7/#�;6Gy���Ն�dI���q��3aR��`�8Ϭ�6��W��Ք�̪�ך6I*�m[����=Q��z��������5�%�zE�S#*=='%�Y�I�
n��MR
;R�,��u��u�g!q���h�q@4���t.w�ۣ�I;`����i��JW���M\�O�^Ҳ9�i���ݎ�l��<5�m1Q�w%���??��Waџt����uʶ$4��H@��)�M꽊�pN�7ko�\�J��[�x˅~|hZ��2��#�3�da���ъ�<xׄ�8x(TR���At��5㢨��5��,��{Gy^�|�����U����P�ye*���u䛃{޻�MᎰ��Z;�☝��	����]��g0�]��尉p]���ഭʐ�2�mm�D���#�A껭�]���+!�b~UW�W�+�:�7�V��Y:`�ŝ���uE�oЏ��҈�з�.���*�����/j{���o��Q��Bb��P!�Ms�o��h�y�gЯ=���Q��A�"Oa�m����1�~��v�6�T-��~�`�uB����N�w��DڑǜU��ǁ�*���.���d�Z�&cqk�)�Z�F��~3A�5�P(�~Q{*��-s~q��%��@f�T�L����/�v_-A�^*5>G�5(�grd��@0+'�ݖ��,V8ɭ��9��]vNC�0E8��Y��7~�ʸd��ӫ3b<ȅa��V@���ˬ奵����H�����w޼o!��MB��w���O��cF�OR��Rޠ�1�w[%V5��t��˘��*l�b�d�εc�M85$��d�M
ڋnobQ�YÜ��@���Q���3�bo�Z��y/�eZ�5�p�X�B-)�Jd�.�n^N��w�=ض/w2<c{���{�2#��_�N8�1�R�#3v���-��0`�x�2�����W;�g���-�'������B��P�K�;Z��y�i��n�LY�� m�������u�x����)]z�Y�i�.�����ىn��8f��fE#�o�Z<��yNtK�ov�;�&��~f`u(�&x�~ M�����uY�|:k��V��bM[U���mDH
�k�Ȼ�3�֊�J��WUzsw�B�k���54�9H`��p)�W����D�r�%{��JV5�*kS�%z\]�=4l���:F�
\ �;�����u�w�A��X�ڝ3�>�&�;��2k��Ɔ���iޥ�ً��Q�qҢ]"�������}�9�!��}V���]���S��CH���Lͅu4X�*���쐜<��	�&\v4hr}|jwS���:��ם�Lw�0�0:!�P�503�J�U�lb�f����70E��/ym�Ͱ����{HZ;�G�H�^��շ,��F{�z!���N+ҧ�|+�TJռ꺑���;/3� Iaۮ.��/�A:؅nB��Bҫ�#$=7cǇY�KH�����9�Y|�^s�`��3���%uc�u�nU��x��ԥ�
��ws �yz�<���r����VX��U���R�	������-m���n|E��Z�1��O����==ek�Spe�ة�=��Gz,�ٍ�u���	�Y{~��F��5`�+��*u�r�h:�Wu�*ZVc*�s�k���jQs=���w�g���`�l�l�$����L�;{��oL�,؊�d�4�b֚ʑU���^���xr�Ww�s�h����BjF�G�i�4/3~��Sk��qa��Л.e_N4'3bti��Ћ��ի��<�B�+�G�h�D�'���)ۗ�}	Md֕y��:ѭ�b"^z٠UR���D���[�Q;��'�����2/�KE"U�x�dg��a�k��D5�t�O�u���9p�[VPp��<E �{b)�71Zs?yFq0f�A\7ۑ�#�ћ��J޴�[U�4��@���('O"Á]�F�ܡi��Y݃���qw��Gj��u��c��f$ ^���B����oS߲Y��t�v48�&�����7􊼞�8���+R#OޔW����`U�m/�e��P�k�m�nE8�O�M�����4�۽�J�w6%0�Ȋlp�qB`In�*��W���D�!q��o��qx�&{j�!a�L�}�����s�09�����x�#`F8쩢��.|��J3�������&�v��er�P�)�}</�b��'��}	1Eq.ԥ��?eFIH�X���&dnnmk���ڕN��۔��"!"ț�ps���4]����gQ%,����'m�$ͨ��1��1�2i,^���}4q.�~v��?����q�ߏ��>9��uf�MPnᾁh�]�x�ԩqt�<|��=+R���n%ղ��"	l��ǑrSz��/�<==�6���ڒ>�[����2��t�=�6��]0���{�]ƫ������KnI��]���U�J��Q�XW7�� n�4;�I���p���9���0綛���Qy���T�EȄB��l�,��Ҏ��v�i��Y�r5E�8B��yP�����Bf�8�̩ܵ���#`�0���&9WRH��G��F��뇁�e���w�8����b5�kpbw��oJ��U��Nut"5F5	���S�V`!�������w��3�^�:�ȒyB�(�G�ϟ:���;���FO�t���ɂ�t��̭ޮvP��m�8�zK��vMPN��`�4F��$p�j�NjiָsT�Od�9��!6�����d�&�X�*�u�q�5�e���8�M��͇ѫ�Gµ���j�& �5�OD�C�˕��T���V4�ӯW�mV,�� �t��kbk�7{��]��W�[W���3¡ϑ�(F��L4��X]xfS:o�օ�ސ�f�0$������	�Q��٪���.t�^s`㗽\��7ë��d�2���Z�nM�lz^D�1g���®T�zn��Wz9oR=3;T֨��aTz�Vq��q����-�;�w�wB,�~��GG�ޞ���+Ą��&^���#;&V|�N��,��D��K`#XP��*�]J�X>0�>s ��υ����U�B�z�ks$�N��/Ss�]*���_�VtJ���:�z�Ä�}���qBuV�V8�ш���ya���"�eЦ�n��t����9*酞��,*^�;�!s��zS�����3b����7[��V�X�V��U�T�8�20��+F*���f�5��"oo�Qx�\�v���� n�0x���[�Ƨ2�����֝p��u�uOlGk������ꔈ�S
N��:����2�s�t��XV}
���7�>����gi�٧ñ�֕GF!%�����f
��.!�%�t��|�tN��ʽ�\Uü_��>jɩ[+�f?:�E1=��E^FF�Vƴ'+Q�>ߌ�~��T
0���KƸ
��Y�"X���h�+b�"�s��Չg��//cuz adB�,�!���"�K&q+�������}�`��FtA��,�cw���nV	��N��Ǚ�sl�Js]��
�b���E<=(�`�w#����,���w��1��c�Vi�}���i9�j�)⫦���HzR�m]�W�Z s݇-mBb�'���L�����$v3����[�עq&�P����6wwr�����D�V�M�kё!�7�S�c���UmU�=�{�
�x]�u���ZT�Q��BmuY��x��}&�ru{��H�̓0����u��+ZR!#ŀF�`��x*l�t̚���*���C�#%4'*�5�4��Gnʸ��w+S�������Y�*�8p�b��d]��c!�3W�V�XJt�t�3*5As�L�^����%��w��7W�5~n�Dp>��	�1�R�#7[��f��x˻H�� 5y��ԋ�FU�I����Z=Ʀ�ךPw��Xi�ux(�
��7<p�ԫ�S���1�Xɪ�Y]Ψ�v�M��֎^�ZJ~Ǡ���k�TX|
�:&6�[���Inܮ��ģ�P)E��8mϥ�A�1Pí��+_��}��ix��Cu�΅�8����9sLE�q*.%�(
�Vvϩ�tb�uWJ���.���v�����\]q�>4sǮ�bSQ�!ߕC]�����,r	�d�[!�Z;��}�D��b�UY�쀑���F�#�5�ҝ�D׺������zh{���R��筚J�U���gV��v�ݞ�1���2�g&\�\��J��]���Y0R�B����7Y��f6j2�b:4rЯ��[jZ���{73L�Xd��s)�>W�Yg�T���-�1a����GL�/{p�ec�ۚH5=՛xph�M#)�yz̸H��.x��r\ ij���nc3��ԕ,8��4f�ZKMraPs�,���C/�M��W-��V{/=��,��6��9�����kh�a��(�3��z�mA1Z�rn_���q�CᬐY}�wV��|�C��Z�+iݜ�+
W���k+8��|�����]���N�#�m�p��*�G�S�Udܩ1jXN��;]�N�R�;�\4�2m�� �q��*��\9�>G�{��޹��,N�pY��S[�A]�Ɠ�g�6��ܗ�{;l���5��]��k�����m@�BN��Ӈ�ԖC�n�َ����n���j�ͦn���D�n���ۜ9��TwE��;[�����B]u��'v����jA����u�����.0�w��w�_K�S��53�yK�dY]���m���^�}w=ɭ��ݵ�x�G/�����$s�|���&���@-�U�t�}�|r^���GC����kctOҲ\��!��9'�C��<�L�'���\��̫Aɔ��
�&��0��`���ݳ4������wV��cV��G�b��bX��ѕ�&I�_�/}�	����TB��ݭ�N�]����H��x���ll��oL��k+=}7*�	;S]�����d+�ؐ"#�e1�����6��4�/ѓ��d<j]��y�K=������ebG4���n�[Èy��G,�aڻ�
�bƳ��I���f���0��w�t�&"���#��V���8�DtU"|��{r�[���,�سda���J��P]�R�яw�&��A_R��a]tZLB�
&�������8h��^F�=`l�����˧1�4E�m�f�
�Ϲ�K�e�-�4�Q,\+9d�Otcy:vsG0������"���]��kǡ�6�h=[|�Hy�h]��;���֎�x�]�#�A���ٗhjQÔ�s"����4���{)� h>3�iC:v��25���(7�V�����a�W@���0��[�V5W%�[�Ϳ#g�����L��}�x�JE9���)"J_�p8��\�	�j����8���su��9ڳ2;b�׷�!r�jd��kJ��*��+�WZ:�gk�ea�)@4��Rp��O9>j���Ũ�1��./�hbC���m�j낞*ܛ��ړ�Mc����(��k#A=gH�0m����Qf펽:Y X�Y�����hS�:��������u�gT�/�����J�-�y\�P��ؔ-*Y�& �Y3�V�U{j.onȟ�)���i��6Ĭ��+mEDF)XڲE���m�
���U+*TV��-V�Taihֈ�ۗ&2�*UT*�b�r�S�ի(�+
´IP��T�l��cXҕZ������XD�+h"�jQQ��¶�-�U��R�X�����[QH������T��Q�-`�ʀ�X�� ���#QT�*
E�E�Aea[h�ŀ�VQ��m%TAV�F,Ej����`+ZJ�B��Ȥ�d���c�b�AIPUY��l*���B�mX��+*
(#R����J�UX,%jc\J��*�FP+*�d��������
�T+Q��F
H��F�m�AB���
�Z���+�Kl��^�}��}�����U�!Dj=���u�>Gu�%wBwn�/:'8���1��S�g��v0Q7y1(�p�����ξ�V&r/���3<]�n ���n���(��G?��$�����E�H��sƅ�+���0�PU�Yb��l+����{�t�od���ݚ�R�_���ƽ^���j>�U���~���N�o�9�YFtV�p�J"�]qP�.<��VL�L�J1z8�۹��&�Xg�=g1�U9�F�;#��;/%�T�~�z�����`wA\\���C��d��ݩ�ad-l����
�!��V?�`�j�{Hɡx���Sk��p�GD<�۸�Е��|�	3�t��s��fD�b爽*	�mDS�?'�}
k&���==g�%�ࡲ�����B�$�K��Nʺ��h�CK*R�H�g�9T�{��K�VÕ�hv��)�m�g9�N����Q�mYc�|��V�hOݮ*	K�|�� �)������^����ݨ=>���ft,A0�m.� ����p+�h�{� � �xϴK;��4��者v��}�%�OD�%�_NQ���{/�0Y��`�2Y�S�}^};Y�.`�.�l]���<���ٺ���!!���h��.S-%4�v��&:�s��l��YZ�^�,}��4�t
��U�{�4S�b�S��7'[��)��]= 
A1u7 l��,q0���k�읽[�Q����9�d��c}�$��*��D�7�ovHv�`>�~R��R��3���ȡ��=��B�,ӆ7"i��o�^"��ҵ'1c��
�ޗ��_v}'M`u�\.��=�o����~0j�x�ԇ��^��my�Jo,>>ێ
��.�_���B�V�K<y%�>u�J�
���5Gr�۳�؉���\�ߟ�Z+<R�d��&�_{�}�?�#��n<�a��"�Jb�}��Z�q��q�����]8��8Ҏ�]0����nT��\�2�<c�{|�p%D��1V�8iG�\�ün�49��#oUeE����LQ��.�q�<��^�X��x��ŉ�tG�����ҍ�c��QJ(�s[�O,	/�>:�%:V�߷�i�����̋I���0yʿT�#Ւ�a��(�Szym�̵����ܜD�:��m��`1jY�t �D�	֠��O��X���3�a;�%x�m��9�s�z�:f��(À�w��u�`+�д\:*�g�����1�dkZ���������Gt_B��W���杒y\��S�Om�Gݹi��ҟI�N��6�"����#Cn���v�V
����T���s��H��љ��[�5&��2>���9Oy�u��g`-�lr�CP��*��s�^��<c/�u�W92%�]ح�f�/8����j��6l��H%�V�=85u= +<�잾��N���Ê(fO�j݆EX�nɢ��"|�C�y^�x��V��'m8��ϙ�B�։0��3^��p�T���v4���՛!ך�,Xn���v�p��wi	�r�;���y؍�ZO�T.`a�~���fS:o�օ���@*��7�;��G����.�3���v�d/��Iy�0!r0�X��mg��&E7\l��p��v��j4ޛ���Ш�8C�W��w�>U��j��T`ODM���!#&��h��j��6�F�oR�W$a�;B��M�aӦl2;#NWH��{���u�!������8���}�5�]��F<�%8�ᐏp�>4-'A��R8���|�*p�z�Y��q��H��p[JJ4�W @�<b�"�4/�[�Ƨ<�#��\�rr)Ç��I��yQE�uVQ�=�ΔEu�`(�rz�"0(��MS!Ms�l~X��<����Xn;SX����P�W�B���r�����Yj�{��X�N#wU��D��:�@�gXv��wB=��Z���D���y�^Z�=6�P�"OL�y
��y)�x�p�{ȩV3���]�dՅG��κ��,�3s����r$��s9b՚��bW�A�IJ�����f�H~y����0d/G"!����WT:F�:`��^�G[�*��{5k��̐i�:o+K��v��5�+֥ �Q���0\#Sv(N*�%������ݮ.�E-�cR��K<\<�=���y�(B1 !8z�N�Q����E��=��"C
��EOt_����3[�ߪ����ê�1m:�6#̎�i".��v:iN�s�80������}�J�U�p�.�/��-�'pi9`�6	M����m�k��vm�Vp��æyM�����W����V�[RHb��#&]�{7� �V�b�����P�9����bv��U�p��^�7j��C�f�v���9��<o�\S�.�7:d�������&��\#�s��N]*��w�P�=Q1m[i:޳���W�,8��+<����SK���G��3[����/Ơ�����Q�:VOu�K̚}B��ZnP�t`G8�+í�<q􍈗��6��C���?A���7Q�	n���A
�<d���ɥ2m��.��[��Z'���\���	���b�ʵ��W�f��R�'t"��ǤM�M�.vzr��Q�J��G2�ŝb+�u��s�gY�� ��[P+��FV���y��)�s��B�uש���U{4hJA�I�&��F��^�ά�f
(�4��n�Nà��a�ڮ2���S�yPΒ��^/ä�3HT�b2c��8��4��>4-X	߇â���}�	��u�s{����F�ݣ�G�6㺦�*���nB5تx���|���{8�'��#����VC#n%:"�(Б4&��/��-C�K!��dUnM1֑�c���b�2��n �y�vT�r���Gx��@�~���NtSJ@��M��N���M�ΩkƬmṽګ�����V��$д��E�FAO{*�O|���v�E7���~��/��ߊ�"�����y(��w|U˭��s71�8�!j����YXY��ݾ�H���/����Rz$^K7`��ƣ�d_���c�
�ĵ��d�sw�"�1sWG3�2�*���>C)�Ԍ*� ⶐA�y��c�s�qx��t}IV�9OhV�!ƱX^�����@����]"�j]%c��;�p�}A�\W��X��M�2�4��e�gB$C��/w�4z8k~�W�[� ����}ޏG����jI�"\<��#�jxʼ�Hu�%�}M_]�$��e9�Y��h�$`S���h1��l���ڏ�Ҽ��j[ɲQ�.���Sp�ӂe�S����w��lg&���ǌ�� �S�����'eND$z��>�K�GqImny��ʤd�[;�yEf&�*����-��٢�5�E��2;*u����Wk��q���'_�"	�0R4���o�f\���/b�p�ʼ��GL [ί!I�ȷ�&���W���x�0��`�/'��7õ2D����4'gm�Ti�S뮐�gV�0]��E9t���W�wj�dӬ:�O��.�q���al97�aE��wN�Xdqۙ��P��Lێ�eg.�f}y����;縪|n<s��W�)R6�E�h�[t�:�<�]V&�8�~�H�qu��O�N��!q�z�(�;t�8��w��tI�Dw��6|$N8�4P/����og
��Б���s�M�}U�7�^��ϩ�uZ���T�'�ʞ
g�PO�D{g�(l��k_r����m$�J��*nQ��Q�.�p0�^��
{<mC�;0��3��'iU��3�[Z29r�S��,�@����b�[��"�q���x݄hs��F��YQ3ڰ�n�R�;��Q�w�3�Y&$�Θ�Ҕ�T�3f���="���fAa���&-(�,���(=5���2��-aAK��>UәJE:,푃�Rieu��]^)Hs�l�.�ɜ�7�8��ݾ�*�˳�ɺ����f�n��c������ov�j�b)����~P�kg�����ӥ{��e(�~�#TJ�: _�;��Y� LJ!?7w�1��"����㰺Dw��h
?S��{L8-��C������>Qv-�:7H��%�W�nE�j��Pp# Bt��;�St<UY��w��
�V8�����9�����%�v �3v&P!׋�	�y4s��WR�_ȸtV��rs7i[�3IT�}}Bk֨Z���Gg�zK�	�5A:Ca�	6E4g�#��[�������%��f�}=7kX��ɏ��)�Y>�}a]�M��[VX�C,�e�o�W���}��ӱ���\�}�D+AD0��i���N�T0�S�W{6��6X�7O`;2�E��f;���!�,I;�<Cnkbj�݌��3�F��00ҙ���7��[�X�+�L�C���1UuC���5n��OؓA�Փ)���V/���*~��6�mx��NluSoLs&��F1ʬ�,g:�N�_��/��G�T84q*��u*�P�G�>pֹta!sr�(��`w�c�E�sSm��]��J�pm�l�&�j��-�ﷶ͋c$�|,&���Ϳ?[��q�bGD�S��O#����h�qIW�՚�gGtM0fX'�*JL�j3]ڝȬ*�=�f�	���;��P��TܣrM=wC7vt�Ƹ�Dp=��hRs�&��:tˈ���zG�����/������ܞy�^��EG�d�qemĥ5M�da�.�4-XN�)̣n9̌1�i'zض�.���yCJ0e=�N 
�S�(C(�B�պ��S�G��3'�C#�𮄥���oS�u�v�<R����(�*9P��Lx����pm~�����Ǵy֣�5�#ʻ�qJs�Xޏ��=T$q/�x�"2]7O�8,]���ϖ��8w޸���Č�{�8�sǸ'݁��3b��ք�Q��f��XсỎ]���s<�L7�M�.q�)�y��X�x����<��2P�aQBVe�FiW[����-�
G�D7���Q���0E(��K7��UC+!���G�Ʌ�{���bn�c*�]��[��W�p?�׃��
������׃���3~}&�v ���N�:GX*�".�G.��/9[W8P0�q�R���(�!]M��t̚����V�5�)@#���FvV��[%d�o�M֑Z�7���V�7&0��[cn��0��<en���x��nIB�_�i�a���e\���OLރ��Em(�����E	�{\�T�L���5[+�^vr�f�73�c����M�A(����'}f��:���,���f�T��X�����&㏦6K�7�B2p�n�U�3v���p�f�u
(qzWZ+�n.ņ�pCJt�ҙ:���� �W���wR��#�_��EO��οe��0�87��CL�ճ1��`��⢼+��4H[a�fĚjn#x\��B�U�(���lu��-ʥ˘u<S�5sT�gH`��;v�M��4���ZJu�z�DP]�I�����#8��Y"K��cT.%��` R��N���:�q��s��hdQ����y�p�
{e��p?���:T��E�K�t� 	P������_C��l�o�����/�����\�6:=�c���(T����!������*��8��9�.�L�c4:�w�Xp; +�^C��C��5�	��K۽�^Kړ��)\��#W���Pfo��y�_�2������*l7,��Fw�OD RӔR1��鰬�;����X����CH_����w^�:؅nB��^�\�E��#�l�
��;g�kk��fhz�ݺh�;�.���d�;�	�T�ҟm�J���p޷c��4��zTEa��w'\������c�d)���Q��V9�o���|�\��Y�w2�p��0�����K:Q�t����
r�]��x3B�$V�g�.���2G�i�jGWb.�^�x�b�][��K�����c�ܻ��V�����eLf�p�1>RHF|}�z��^B5��8��YO8�
�B�ݓ�e��.�y�19ZX�j|F�%��e#SR0�� ⶑ�x�<R�.�mY��L�W����yCNC"�;T��O��;\(�֣�b��T�ګ�`���O�Z��۹�Ž2{�ض���&X����9��eM\M�̆�ꊛ�R�J��g�"֛l��7��O���m�a�(��c6h��Ֆ09f��DU����SFncAfw*A\@վ^���{�:L��d��o���#/*��#f-�W�N]�"v��B��"&�^�Q�w-�&|P�:��N�ڜj�ײ�B���`�,�k��M�����Q�M^ۏ3}�&��\*�G\c3a���i_E�Q�1�v�(q�s>�;j�,��q��ӎV�'2�(`�R(9�zCqY�}�H������H{��|�U�>���w)V3 ��'�N�4s���dl3���⦯T�@���5Y�ß��D�vS�)xt{ip5Е��.�+�.�̾\�����]X�!�O_b+ggE�(����h�cs�>'��s�<=WӋA��(��)mݢ��tZk:fU�{x8����(��W��ǅ%��m�̍���9.ɑ���I5�VZ&W"J)�NT���<]��(uv����<��c�&��䵴{|����<�RWf��j���$8��kwY�T��:��Ko4��W�E#]RkB��r�6Vxx�V����Y���M�1��;�d�r�E��C�A��Ro����k�xe�Vץ^<�,�j�{ѡ�o�r�Cɚ'x��g������o.δ�3B�YǑ���2����w�����L��Q���ꛀi�x9�W���lɄ�cov_F^NT�x��zI�8'���q�q�C̣�7�v/v�i�Y+$ͤp���~^��L��Y�R�yoU����ki���&�	j��bƭ���.���܁c�7�/�ւ~�Mkox�EQ@��j�9J��Q��5�t�Z����t/z�;j�fǊ�h�%�y��/\�3���I���͞�K���ތ�U��əz1È��!)u���h�oVeu����f`�x�7��0ݕn����>�E���?^�A&̔]�ׇ^K�]�ײ�y�ҁ@�N�.���5Z[F�c�����B��q�c�����c?x!�G�(ˠ+x2��%esj�6*ܤoT��b���Q�`/0EY��eK27�����/��'�9�0�>}���}�Gq�=��}�C&p�/$8�ĺ��%Z̫y��wgGw.V{�Ïe�r$�{(��=|�a�t�[�@��&L�y�K�DQ��$y��.�y1K���]RE�U�V��`�)��j2�n4��H?���u�u��nn�����{��`�\��87ڃ�\�1;�loqѦ�&�Gs]d�՜�v����o���!p�d򻚊C���o�]�1o�61���Vc\�0�=���9ԙ�&���}���W��̬wS%)�sDIԝCa�y,ᨬ0�:��br�>��Y��dp�>i?��5{a�ؖ8�>�zm��bvK����8���Vʽmӛ-��xB�K����D���&�Og�6|���vv������d�6Č�R_]oq3����h���]�X�đ�s���Ê/�z�I�~*8�����Ʋ�~�e�/���H��&{�����S�M��̬,���x�Ӥ�v^W�Tv]�p����td����)�R�y�:u���aY"2�x����O_NluƉ��_���V�毩�W�1[)�%�xR&�]j�[�y�Ѕ�a�+
�Q�#�r����q���j#7��=�Cڳ�|�Մ��ҹV\Y�=���l\.q�7����s��eĮ�J�2m]��ʗr�_�y�ַ�Y
���b��Y*���X���*��XƲ�T��VT��%`�Q�T`�b(�


��%j���
AH�5Z�ڢ�VH�-�b�Z
J��AEU"���*ł�"��UJ�X(*�`((�JʋPPX,�,�X��"ʕ����V1$PYAk"�m�-k
� e���l�YU��#�b�m�C�ĕ"�E�b�H�-��U�D���PP(��J�E[P�IQT��`�`��Eb%J,[eE�j�q�Y�)i
��� ��
*�j6�J0Y`#
$�PX(!Q���,��U@|��ٳa�<�B�ևG� due^�tRa�'�3^��A�����;��LN��5�W 4ۢ��ἒ�g�2aI�gP��S�_���f� �� �P�7bHM�DP#���<��
���]x�$�v�3w�cbq�(�岦�F�|g��RuKa�8b����߽��-�
}�M�ɥ�������X�T"Ԣ4_M(�t�~h�+\���g��p�f��gD�Ρ���Ȥ {�[��Gx��T��(_Sp0Ҏ#����x݄k��b���!~t2^e�5���\td���E� �0���0!tϺD2�W�N�l��]�C�Ot�uһ�֐���㒺tX*{��w'��W�@|g�aj9W�D
�G�^�5vP:N��n�:�vg*"oc5J*��e�W��(\~���EJZ)4俛��:���Y/5�̴oô�T�=q{t{�;]d���雈@��� ���W1����f�����x�wl�͜�يqb�Ud��]�&�E8���3�3�=%��;&�'Hl<�!���\1q�8�x�]�	Q���f'�Th�͊�蚷a]�M�kj�!�C�@�F�x�wn��F���Q��^[,��'P��p�N� �7����T�{3��>�71nd'k�T�����Y	�]�8R~��<Vn>ژ����T�:��&f�3�k��347�Cz�R���VjZf8��(��vZ@�*6�qɜ��˹:<K'2�e�&�@�8��tNN8yS�kيƛ6���d Zj��"�tZ�ɜ�܁Bu�������9�,=�ؚ��dT��24F��00ҙ��2��yօ�e�
���7T���*h�`��Y������5��C����*�c?(WԱxZ�U�1�u:�(>tJ�I�dv�:j�8�j��3���N�ߓ�|V�Y�*0!9C�ߪU��ح�#ֈ���q%�tZ��u�E_�%^���
Nq7XE�Ӧm̎���N�r��zcrU�e<q*�|�lbd��r!�*�%j�p��x˅o�V<��U�U�x������~s�9&�vq(���xEǍH�#�� CS�(��J��N8y�����ǒ.�6�+��H��ɧ���B�}�(���X����!H�t���;F���rCF�U�^m����D�G[�v��Q��A�&��q/�`�"�C+B����]�g���Z�9�k�*^!c�|�aP�qI�q�	�`yk W�J"��"�VG�@QK5�G��{R���U��T"�D���<)p��I�#X6X4V���yon�q�o'>�*dG[2Y�r8>A�a�O��=#Ѻ����;����6S5&����u^_#J���;Ng+�Q+؟u�أv�]���Lіs5V�w'P�vͼ���n���S���<�O�U��x������@����#�ճ<=�Jg��~T�i#���28����c%8Έ"Tw�	f��Qe\2\͉�I�G�N="S�=ev�^?xQ��hMuay���Ȝ��>���#at����욵��G!�N-*�u�d�`8|��
��LѠ�0B�T��r̚��b���	�|�����&�<cw���B.�d�hV�Xnobn8�bF�p*�8HF|-��]��-���T�;�j�uۃ�i)�!��HJ��Y~�un�x���VO��\��T��q��^�oV%x���z��T�v�,8���e7#>��*���bM[U���n���j���6�r\�D�!�7錨��D���C��;�l7�4���6"o	��|��\�Z&i��)�VÝ�a!�[,�LZ��B6i����܆�B\R<����Hulno{Aܫ�G�L�_�4����t�8��5H���螭{��4�Q��E�P���LJ��]푁+�w-��ɹ���#�|V�V���:�oz��T��F�fG㙯]��w���%ޙ��}��o�R<1nC��|�sjn�:o"����1��� ��ԡ��$��<n���E�Y�5��bn-�Ĺ�E�[������t�ٷΡ�9}�G��޸w\�Th�]4Ħ��C�܄L	�:�b�w.�؎�e�)6/#�s}�&\w��C�udpd��ЇJ4$F��	��y!+�z��i�a��nb�c�m�ǔ8ʩ���ٔU�n ����囘F����
;��s�q��������p9N�R���5ծ,gN8l+���<�����V�q&�MQ]�gF\6�͹�;�Up��Hi���zL��S�9^�x���[u\W	u���U9t�rO��ȭ���tˈ�t,*u)xQPUw�DqڼPn�\��f��g�Fm<"Cu&Z�_)���u��U�ͷ^"T�$2��&�aW 8����tȁ��xDsg��=o�o*uA3�Ӑ��hV��i��k�0J�|��(�&	�m(�vqU���`�˙���nTov:���Ǖzo>�~��0 �E����_X�
eND${�KEz]���Q75f���sV�f_(͇�"}w���qŸ7f�q���,c�`��DV7^؊�Fn`$U{ќ7�ϱl��asw6:I�oyϳ͌xGG�~}��
�H����N�6�I"�Y��2����^�����G�9u�]vY=,�R�(�y�h��Y;7�RE�t�L.C��$9I��n�u�zR'��-����jZc�A����!u��gEm�����K7.ێ#�-�W���<�p+�h�2sjtY�}�]���e�z�d%��;�FR���Un��/� Y�ަ�dK�ɽ�9P���Q�~���i���bG�<4�^Ǡ���(�],^��kC�U��4���	��]W��K��*:v1�Hی��A�+�1����u�"hT�:���H{��"�ty�QF�}�x?l��&�p���!�&�����n��3ح�޸N
���Z�F��٧z�uZܕi�J��ϕ\O8�gM�/A��A{��:�K�y)�Б�WQ.��D���mB�v��=8����Q��h��"ӡn�/��uFS��ez�D�ƔF�ķ��qj�i����"���G�p>��*��*�9�^)E`_Sp,dZ�!TVþ�v�c��7Y7���z���`��bô�u��u��Ƅ�d(�u��Tzt�c{��t#v4R�:�y���+�P1C�s�+}w��N�ȵ$� ^�QB`�0H��(>�[��n��?���qgH
ʒ�|��c��v�|@���m
�\����IG*0s�~c�9{̰p����t��]z{�*��G}=����Rɖ�8�ٸ��ʃ�#����t�Wv��,m�(W>��Ɉ�z��tq��mf��]n�K-wA��(��Ot<n�x�E�F�Z�u�C���+ʊ�KE*$iȗ�`����'���O��(Y�㠋�\�~��3���?i�7L��ep/���p�`�c����L���yԵL����Z>E��V�T&��qV7��q�=%�'d�'Hl{(B�<�o�Fo{�E�+y݂KH?���,!8tĹ�Q�3'�V�"+Gu�q���,Yz�sY[�1fU9}��� !+�l��W�@�F
\F��*p�{1X�~ͷ~��/�m�{+)G*�3����(?.��,��"��lM_���S�t�����J�U�׳)�9���8��B�]ʳ��Ɖ�5�@+���T����_q�/Jت�u*�,?_��vV�AP�r�zowj�uҍ���iU�E�:�:w���|SS��=�bu�~�Y+��eg��w����Kt!��2cz,
sEa�F���J����n��Ӧl9��s���Q�${B���ؤ��߷����}*:��Cc� 0B<W�J/Tۆ}�$�B��	��I滓]��Oe[�Y��ַ�����<��@.���F|&���Jڹ�hv��8�j�t!Ea�PL:_Y��f�D�+8�G�� �96Ag.������#���J�6���;��</���va�I=W��c�n4���j�{+\����2x���x���8�]:Y!�u� ^�{����W�@�1��2�4.�7E�fi�㕵��#0�ކ�O?^[�
ӡn9���B�
�`t��t�t�A����+�Q�N��7u�k�Z_��_�Vt;PnQ���P��:�L�0ez8��`�b�W8�n�&2���FF,�J]z��'�o�A7�"�##V� W���y��k�s(e�9Μ��E}����%ׂ���CPfz���Լ�=���c!�6�_�h���|�!#�G�Bq����/g�@��0E(�.��u�,��({s3�U^�ݍ�����>�9G�(��/!2���B�x��ׂ:�}�3;+��H�k��ٷ��S@\��'� ;�W�6HbD��
F�x�(τ�y
�l�9fN�yذ_�'���z�%˱�[3����"����=g�/
�<>Ek4�$"0�oEW���+kq��m�G�ޙ)ۜ=�l�;��r�ȴU9#A����r'�>�����~J��x����&����'�[B9��[��^�s�
�5]�_=ǖ�oe�CW�7N�񻀯z�\����+�b�{��9tɚ�u������Bt��l9���{o�e�L��ۓݼ���rg3���<H!����bP�b�%�eެ��s��'ŇU�U�ߟ��G�Ƌ,gmYX����Bثk6$�Ed��e�X��\��B+2��Rdy��ʊ(�@\� Y]�Ψ�v�M��4�̆�:���O��FR��Y��'�S�Yz�p�Mnq,���@�lӇ�ש�3
e��%��B���� >�v4�U�V>�Mp>���(���_3\4x�8&����:��UY�;����lk4-Xn��8ΌQ�g����`Վ�H��[LJt��Eې�qf�̋�sEj��Q��Q5�#\1�N�L�`cF�6���8��(���J0��e�T�x�C���UL�/I���z�fQ��l�,��m]y�6aZ�:��eM��F�V������L���fw{yL������]�����8�IU��ۺ���lBpD�9;7�:�&�mrj��ЅV�UI%���ySτ\EgM�7J"�]qQ��	����]��&:�y��b�QFEy	F�}�
��y�<�^��d����j�{��0�ǚ-LU�gU�^5�(��vʧ��[�
�ZJ��$�}}�J���@.b��kV�0�Ӆ �X��x�JU��2��Re��{���G��H;}�#ݎ]uk=I�vͺO�����Nk̰��%ё��f6�7�9�JU!T9km��l��ƔCƊ��I��/�U�	��
�7R����\�ie��M��M8�܍j~;T���&gk�0J�|Ŋ/IPO@V҅�ʊ�b�ȷ���Y7��7��j�E�ԲB$����>�����9�ꆖW��U�.�ՙMn\�;.���'�I�3�j��9�j�In]Vyq�~���Z������&�'���qܾ�䴃h����u)o����Fᲈ���n8��@�����n��ƫah�7��Ԍ��4R�e)�z%��;���ʍ5B�{(_P@����`���^����$u����	�#��St�0�¬u�36Zf����1��U��nrKL�o=�@�������6� 4܊q^��77�=���P��c�R�Ku7p_N���[�ʪd�o&��ǓO��q�ۦl�˗�گzʌa7��^��Hsr�ܷ�~�Ba5W	PΤ�����CJÕ��vB�*�C��j�:s���M�zTD/T91u���د*���V�<����m�
�u+�օ�P��طF�=CI�\�0Ύ��;�.N��}P��颅56�6���6�<,�-z+}E.��+�u�\�b3sj�eCx�f&j9�y=�ˁRC�I��vH��UKIim�.��m[E'��]'�����~��݆��-��4��J���[�z��Q��l��]@�5�Mlo?�U=W6���Q���CK=3�Uڰ���{q�o:�Č��~V�Խ\�V��jӨ�^�b5^�����/*�(9]�a,�6�]��jv�V���CW��i�� �yG�]k�V.tT���OܕD���8��U�:����j���gϝE��]��W�ХOxn4F�1LOb�ID�Ү�v�/l&&Bhc����ް�S����o?Io;��J亲��w�Wp��v��u7me1��Sp�	�H�*����ɯ7Y�Q:��c1��˵ur�!\V'go+}��#�� ۽{]�~{[A�2���\���N?yF��cæ�K�eb@-��,
5��n�Q49�P}��4&�!*��y���=O����<���q-�b�ܟY�qN�����2d8f��H�8�Y+[�m�HY�t��fk�}S�Q��t��븰��ẟV%�Eǻz��V�q�a�\Ftʼ�J�
3�n�q�mS�(bj�(����I\���O��n��-	�v���3#�2Y�;'|{���A��
�ħC+G%[s�S]����^�1c�@�&XW&�T�i9��l�R��+�4K�-k6n��yn��F�s���5��"�3���7���
�>��/;_E��m�RH���yn2�]nD�÷�8��KF��)��,���n��z;Y���s;ž����#��@��]A���t��ıZ�iKʈ�s6��.�w�9����a�u,������:�hޅA�92ݒqLK��*�?Z2rћN۶R�O�/"�p*i/�3w;����d�{<#씭�����
�I`_f���fȵU����#�3�ܥ��@O=�afT�������r-w]����V6�2�b�p(kk���ض�����ɰ�r�%�`m�f���(M��1	�C�U-R��3`�i^�`#N�=c��e�o6���Ƚ�Rea{��>��� <��0����Sg;�z.��R5�\,e+$�j���X2%y���Y1��[;U˽Ͳ�#5�%��,�Y�P77v@i��aK�C��ٕ�W'�6����v�mskSO7;�۽)wgo�\��4-����t�m����`�����K���|�͂��l{4y�Êo�7/�ɳ���J�ש^_5���5("w.�^�QY�8��w�dA�bm��l�]%��w�6�	*���f'2L�2t�芣h��I݋�G[  ���Y�/����Gz{��\�U�Q^�;�$XR2��A�"�Y�9eZ4@�rMTN�N�^���ɮ�CA��z\w���Y|�����ǽ<��Svw:7�=.e�v����ʔ���j�M��q���罨BG��J�FoS��78�TF�r���+Aݘ(P25�o����X�y�[&�ǰb]%�S(on$^>C[�fJ` �\�da�a{��ܖ{z,%��*�[`5�.�ծ��$�1Y�7f<�o�{�\Lw��f�ER�_X�5�.�7[ѣ�[�����ڼ���E���	��(g(�n���n�^�\u���;������ޓbm��T�R�����{������3����˾o���=�fY�]���Te��.�A+�\����>�u���=Z'��9>����[Id!�U���W<��=�u3gL�9�?ok�}�����[�[�&��lvo�"$��A��IǊ�Ȭ����y.�(E1>kK����Ҧw��<��t��ⲧ:�Q�sӚ��7*[�VMfW`�'-*|$�\e�0��2P���"s��'���cb������T"���X6�AJ�J�%�P+(�A�1++6Ɍ+r�R���,X��%V
EХ�G2��Em!D*H�#j�
6�֐��
�
��bH�,G"�m* �YP+*)�+A���C*�1��ed
�X��T�,�¨�)J1adQ�H�AE���)d+Qa��b
D`�d����lU"%s)��R"0�cjL�aD*��E�����B�h��V" �T�0Jږ(�X�V((�1V-e�QV*1U(�9j����f[*QEH1�����CLL�TDUUdY�ŐQV���b��}VN��ىE;
�2�dv��ǰm��A��3\ ��L�kR������G%��'�4�{$���:**ȫ��C���]iC ���i�Lcsx%�ۮ����n���wE!Y�%�҇j��lƗq��-�inR˅R}W��]M�s�a��OV�y��u��Mﺙ����k��p;6ޠ�����S�����zᄆ�|��a�t�;6wj33�
�z����H�8p�}���]��c��B�>VR�-�<zZ���Ih4p�-G���ȧ�M$�����^���ʚF��q���_RrN�-pt��D�g�e��Gc;�V���m[���4x��z��n��N�����FJƙ���V9�}w�U���OS�s^��e�^�,%�N�����N�����JԮ~���gZ鰯����u'��ϫ&�iT
.���b��i��SaGm��^�b��#QZ���[�4����:��۬i77;�����/H~�f� kU#��Uxo8�\sjl�ڼ��9���U/jͣ#���f���u.x�{TC^�h��%qc9�T����vW%������_K�5�0vj��ɲ��Sz.�kj%@�t�&Ů\'#%=�L�\���<偽�G��������d�Q� ��܊��,��"���J�m�ě�:��V�Ҧ$�Ǚ�Q�x9�)�A�j���bC�q~��4�Ug1g;(��q��@䟓!�1�@�Fc��F)/���ۈ��˫��'�/����=7O��Mc�P�8��|f$hs>�Df6�75$j9	�\���ͽ�ز�v����>�7�"�	V��Y�{C�����]���ov�Y���}N3�ﲅ�7���~��V{^}��|��Ԗ���a=�͹��ʻNh�iO194�Q�%�:�t�:X�ni�^L�ހ�r\�zf�R�,�Cx'%P�|-���;S�1�vT'��������[[�L���\��7��{T���ʇ��:����~�o���n3�b����C� ���ze���Hˈ�n$�.�x�e6��5a�C=^m[�8�~Q�|�,�*cL��^�X-r��ǉH�ӯe;��p��q�ЭPllG
 
�ΰu��bd��v�F3���(�V�Љ���+�$�m����|Wr��n���n,��:��E�<���D�B�N�0��h�Cf�f��%�-���6��[���5,t���mԫ�)Q\��J��tڻ}a����{�:ۨs�ֆ-��!��s�@���yQ�>��v��{)_s���ҷU��wC՛�,��R��jq���ҩ���ګ:��Һ�؍��Cɦ�:�7�d�W��Ƞ-:�H#S��	�Pz���P٧t{P��b��j]\����[���SL��ǐ�"'q@s��m��V�q����C�ή�Ԭ.��<!��:Fb@���7�ok}J���uٵ�����ԋ�{n���݆��I���������b�<������F_r�w�$Dcc�k&��^�j�v����q!�,���1""Ϛ1G3�ǫi�����jqc�#�+&�ݬ�^S}�(7��CNsWH��I޸64M��⾲u�W�W����Vt=ь��BrdW��_W���c-Ӥ��j+3}���Z/=�����5.k��2�e��/8���� �ХLS��X��v=ގC����ƹ9�b�b���ыm������|\����Ƹ����u��{g�	e��NM�Cq��w�������@T�����ag��]3]����[���\�����>����d!Y��:w9+�K�o��
���{X[I�7N�t� �ny���{�+8Ba�sw�N&�>]Ӛ�k�/��=4����;v�qZ����͵E��(\e_X=��%#m�
��P�\���:�xSVU�%a�Ʋ�C`�Ӿ��a�W7�v�(����ѥ^������r���˭��VHɞ����{i4`ܙ{��/!�����T�)�����}f2��읮n�9�L'·=*��Zw#2���I�r����t9��~\��c�{r�5y6�-^��Һ��<�[7,Zu�
<��`sA����ɣ�b�WL�k�g7�uu@�v�N�IZ�������L�A�3G�w��������#�߄��VtV'��u+\u������	�#&�∻�Xl�V.ױK�e3�����rbQ �]��z�>�̳��Y�QlmsJ�]�κ��׶-�V�����ΚR�Y躸:Q@]t�F�ރ��+!��Q���c9���J��Y3g�����4��wfWOv�Mn��&��.��3oH��W���iVs�ǚ�1����x.:�x��I�&pf0\�SFc����/���v�jݪ��mjw[R!]����1s<�\�^��A�Ƞ��u�K�^��{����;��3�7�j�oj��T��0�������{[A�24=�h�>��J���]m:����5x��-�c5�W�]~ImԷp>���Y�+*��t��wmee&[�KR�oљ]brf���%�Sw��N�<�'�{^�j����TmJM��l��t�%H���Q{�\0�������~t���TXFf�Kp�r؂�շˡ=�l��>���	P�M�=--�Ff�cyT�+�����A���L9X��dm����0l�q�igQ��Q@�P�˴����M�]C=@6�ۇ��GC����!����2){ǯ7Ubj�;	e3L���f�Q�7u��T!4�M�gv��19�,;�^)�Lܵ��Ԯ`����ƏZ��KJ����fs��7s�|��4����vd�<U75�x#�{%[��Ѽg�+����3�S�J��wG\��$���ɔ"r����u��HM��o{�)���M��a��\כu3�^ަë��ޛڸ�9dgv���r�2�F*�םO���:�}Ԟ�>���@:�U�F��JM�|�B��^�@�����c��nq�����Ї��A����F�O]!����A�C7�h3遭T��+Q������:�f١xH�3U�J�z�LN��i���uf��=��Z�U�v�E�����i��1f�1+��l`�h�HΌS�Xy,vc�ٓz�i�}'u㚹��yn�{U'm	b�j'ɡ�^n�(>3�<1I+x��6��سv�"��홆^z����U��\�;%9!_L}��U�-Q�L+�+��F󙽭�H9�x�α8�]���o�oS�vR�޾�tln���Π줘��^��/�S�/ՊpOH�t�#7�.%��l_:j�t��ٶw�����)ʻ��	9'�1v����z�,H*�|x]MࣸG�`e0�Y�𵎅���]�rl�4n�;�j�Dx.޳ް���3զi�r��k�\nR��C6<B$��1OwuN8�����R�h]�(Vҩ�3!���˭6���:OiQ�]䋢��vo���&��2���FKv䪸}W$�VL�/��i\��Km�Qo����Mלb�mls�.�d�>��*7��.Z�[�5 �|o�m�٨��9��N�Tn���H�F�h��1��[청�S9�U�Z��њf�:�����ƝcG�6��q�
=�3��yva��{�(�$p�r�s3�u���T��e-l�=뙺����m��1�]�J������Qa,,�lWj����W����X�`阀f�p;�۩�fOo*��n�W����CK��7T�U�z�CT����j��f&v*jӡ3���EN�P#j���#�Պ���O�3�1�wJ��v�S�>�k5U[���P2'�3b1��Cb���{W5p%�\M.��J�	}~mQh[��WT
�=�h|s�U��'�,f�����뻠9k��x���MH��/Z���tfD�g݄=�l�	��@�W��p�PI�+9�jfS�֨���Nij��\�0a뭇]@)Q�M�OPV>󬶕j7�	>{F�y�n)hv�+�s���JG�t�uo�vayIGU�o;vЖ)1 s�j�SqnF��7������Ϻa���C�Y���n��]��^;U{�݆��m��[K*�Za��/�ʽK�wr����D�g�9�J)��P�����Y���B���wOkBꐾ�`-�ڰ���j·�1���Q���NM�B��_<���M�X�6��Z������&�i�+$`�qˁp�Z�|3�{��Y/�j��I^7N�7^q�7��{ǀ�Y1�y�i��Lt��I�S<qoZ��3���Mj��7^q�(���kz3��Q�~�Q��o�'	��/������M���ϔ���Z�-��b�ϻS�u���q��C�D�J)#M-���au�)8����)�R�BxNkȪ{֙y���AuL�2siGe�����S[���{}S�����c��:]�S�F��ueG"��[HH�)���[�mSM%����u�y�q��Q��o-[�}]#�I�]x tQW�zE�ű긻b坚J]�޼�]�_J=6-�%C�t�i�f�m[S1O�=�����z�c��=*��sBҨV
+���Bg���US:ga�v�J�ٌ�`ίg[�Һ�z�=��nw֝@�/j��H�<��x:��r�����Y�@��ѭ��V��������i�X��;-�w|��8�_�7:������7C�u+\u����s$��9}�*���Y��k�������V$d
n&�mU��n�U�� 5z���w���#���)��h(�a�1>��DK�~��j&�ڭ\}5ð�T�-���u�1��,�-���n�)񨑡���>����y�`��j��y�NIxjB�5�U��ٴ���1M�{=u��lM��{�����U,�䃜��Iӳ��w���+o٨*���	-�Է_VD��+��8���opU���s�6XBzam;���7�q(-����g:w�O('�z��&�V</y��x�X,~�D0�2�+�d�����iW)����cZ̕�䃇[q��(��v&��:�ɭ�޻�H�`���'���P����сyq�Br�6��/�8�c��_s�h��Y��W�R}w9G�s���޴�+�����*�p�1���zU��XK��vv�*��U�wb������5/_c�n4�����>��� _.	V*m�1E��l��cɗ��؎��Ҡ�jܬvvF�G�vȁ�f8@k�Q��ke��]��Ut�#5	���6�ڿ4k�=M�v��;
8�ȋ�a:���Go�mya�ޝ��''�%5<���6�w�z�����~,�]�:o��'�mq齼�_��e\ij3���Y��x+�u~��'���d�w��{c;�'f^�b90׺�׾؍zF��9�Y�[�4����J�����v&���u���D�a遭T��Sg�;(w78w-g��ܨ�q��˚n���0�cN��f�1=��p'���Z\d[�q�[��_V0*��[�Cty�1<ΌS藊 &j��n�k<��s��S�>Y�)Y�*��0�
}��+��C�W�)Mi��V�����ўt���*��D�Ȗ�}�O&���mƫ���W�֕7����)gTa�ۇ�撗�ga���U�p�`M����'5L��nVu�!�p6*��IH�7����Ia�ު����k@grΒ�l�>�}�W	:S��ѧ�5�x��}R�⹌=4L|�G2R��]��ygHYV8�
�BZ�`<oi��GA�V������K�*}K�;�W�P{���]����@�uZR-���HJB����9��X��L1Pc�2e�N�]�/i`���(e͢Y�'7�)`�7�/�-j��X����w6&��ˮ-�=�=Z\���F t��8j{x��6yY��`�D��(GLs�蝦X۬��߅t���I����*��+��u8��6_�pY�ݓ����3��ċ���2��kL�g��B��w9oM�R�)u3���+$�u��=.��@^��w��O�&�j" Ω@�Bu�;{���{�H�����<S�=��H~Eр�g�u��h/�S���b́FJ��/���W���zG
V��'`��ޑ���7����>qw{������C�v!��4L�ߤ�Nd3���A0Wj�����/y(g�Z���� �L��f"��+�c��jpo���{ Q4Ui�^(9 �ڮ��:���x3�Hj�o��A�I� �t'9��аz�������@��<��G��f���+F�!�}�q��;�hk��BY���G&+/�7b�� ��.��{\]-���2(ɱ�:7陭���t��j��q����f�|H�`m��� 8���u��r�{��iB�WN+6�t?4�#�]N�ـ\���C}�/>K��F��D��=�n�"�,��D0~��˸�(���2�鮣�]�C��J��<��x8,��ZXz��RVe�ЬOU�[��7� U]����[��6��M�}�5r��pn#˕v�t�!tݙT���:�M9]M5�be�<��X��5u��7�cћ ;f���7�y��<��z�*�w`�m��`��@Ȭ�˾W]C�P�g�5�*�`ݛ�JR�t������R%��ąN����]��I�Μ��ޛeS��A*R˺=�3.>I �Z7�mq�_v�y�J��nܬ[����9=�*ߨ��|��Ф{ɜ���>8	��Xt��,��w�B�U؊FzY7�!7�һ\x��RT�3*::�6����؀s�+�1���W��I�ۧ|�NE��*l��{�	��"��8�6`���οs�:Խ�u,\.�l][Dm�^9���.Y��i1�h��Y��p����҂�%�=��&��:��θ�d>�/m��R�gS��u�dP�^a�oWN˩w��*(�Fj}�M/n�
`dΠ�{�~�{����ǻͥV(* ��2"�*�Q�ED-�"�+�����(�B��#��"""��YS*(��TUc"�1�3
�+TX�G,.2��[A�� [b��1j�REYU\�be�P+�
(�b8�m(�����A�VT+�Pm�D�"�!R�Z"��*�[j0QF(��PQAb.2��F[+b �X�PV5+"!YPUF�)iQEIB�1
����[*�m�*VVL��������[EX[Ab��-E��E
�"�Ab�fS1*�PX#[�������[jX�څ��J��c�TEUb�"��Ĳ�H�"��R�´Tm���UX��R�T�(Ɩ�-.P�U[j�@Z9Je����\�T`����#-}��^�����w>,�4o^g>�r��[c������]�Bnj�Ѿ�,܏���`\6X�[�{Z|8�����d�Ime|6�$U�걽Iߚ�y�C&���|f'������Tl8Cg���vX�pָ�˷�/��n�b�����G�o��d�^+7�/�r�C�uy(1Ȍ�W8��e�o�oS󲕦���j���\�s�Z2{w���bh7fF���	S�J�93M�\Jqs���5�v6�OB����R�,�յ�-�'/����Z��}������m�Ӽ��M&@ ^��7N�7N1f�mt'�z�d�����#*S�4�B��k���T�ȵAD����\�t�;�ͣ#s����Wë�=���K��U�L�"2)%C��c����Əw�V�8��'�xf��+�o�C��	RZ�*� RFk���]6�}~l�Z���Nh[%8��\߻�¥������ˣ�ѥ��'��������wb�Fw���:���[���BFh��ޙ
��W�C��:�(����F�Fw�7q���ע��wĦ�Q��R Vm�x��\��je>�[{R]����\�y`d��\�>}��_cv��t�\Rx����mp�y 5b�W�4��\˵20P�+�-/��M;װw��-:��x/o��&vD7C�8�*�98�*����Č��~V�Շ|�y�a�ȫN�PACQ�n��PX���1�!ͮg3�8�;]��SUB�`���"B�CV��ruڧ}���)�K1-�$(�Q5���J��/��Uv]�!�1�f���z�Vvv�rcZ"�_LN�Efx[Q5{j�y۶��^LG>��x}M���<��.F�i�pE}+�WVxE��o&�e�j�n�md�G!�3�����+cnU�n�+��ϸg��r��U��W���Ok�o$J�9�;�Q��l%�P	����V��&�ՙ��F�r#2��ɧa�=P�%��6"�_��C�yB�ӹk(7Kw<��&�x��b�W�����h��LڐR'���m�%˫�������7N�7N1f�w���BƤ�&w7:�qv�FX�yu�M.�+���v�^>v��]���p3�/z��"�iǠ
�ܹ͈�����1ozbG�O��q�jr=J:0$9�l���{Y�J�'�#��lӓn%��!�t}�J����f��\����sZŵ�ޓyi�!���T�Lr��J�p��%�6@>vܷ�q�Mu����OL���+z��(�������� c�@�yp�t���i�qL�F��֦����� e�>��Î�V����P�
H�ҡ}JX���T#�G���U37��fl�eI8jz��{֙y���W �!��m�ң`�K�i��h�ű�z�Uk��isҞsS둙O��zI���˰C=�V�i+���+h$�:�<Һ�z��Ofԫ�f�N�\aق���5������~�#��c�U@�U�5�i+X)��_Xn�F���u��^�N��aD_�3�s���*�����R��:�mU�:d�k�V�q�Y|��3c�X}����}د�2 ��Evڭ�NT>Y��F��`&&[C���FbxEՓ
�z�⫸X�(3g�������ơ���Ⱥ�l���U����
���^��6�Vd��aG����k�>+�v�Ŵ˜��֡{���ZV����J*0"�z8B'pQ-s�#`J��%/4o.��
����V)�\}���X���g�+WZ��t�tյ���6�^��A�ȧƢt9�f6#������Q�=�Ư6߶�U�.�6�v�(6���և��5�·�h�$�qEU��q��Z��/����qM�e����%{u֒���[��ױ9"Й�5N�vr��U���%�]!	s�X�����%������ۧ�"E��;ڙ���'��F+o�c�o�W>%O�%��[p���	X;)�;k��{_���}|u9�Yw�q��*'���2(vȁ�Dd�B*	[�k�: Vu�l֞{��5Y̹N�To����^1��eF�*b}��`�Mf��UE�oTܾ��h�cG�ͫl�����,J�����_ݼ���eF�$�T�����V�U�i�z�[s淳���v�Or�T¤_��H��L�J�j�����:�}Ԟ���m^zڷ73�%^,C��{s�a7�����8���1�d�\͕�����z��<~+��/`�}��;	ɍ�s8�<��-ũ/��&���ý�aNF��ۥ�n��؏^������fr*��s!3`�����Or�m�.�vjY�9i�NrNw2���W�8ڦJ�vcQz�gn��WZ�<����\�8�gk�'Y�F��n�Zd �gLj�ub����2�j�/V���Q����uu���5�˛@4�+�3j�ج	�u��y�h�8{/25^:��{u��U+���ؙ	��˰d4f'��щ,
��:��;[���3����'�{j�z��4%���C&���|f+�̳vR��j�^p����1H�Ʈo$]��x�Ս�B�bq��b��:�}�)���{�G��.���̰�,��W8��k/���L;�K�s(�����&ս<�F���y��M�Ί��*D[�brg��Y�n�:��$�V�6�-��Rr�Cz��VD�y�P��
�%���x`�q.n��[=���VvS�ۧa�tb�mls�/�+$p�����9뭪� ׺�l5��,Z���ʾ�̇.�];E�����%(��oݲ�V��ߎ��K�I]�8��R{#����/\xNj��Y�'-dt���R����w��]w"��+gɆJ��+Y�<o��<h�)u�fu�{�&'��1;��_r۾�Z�����RX����I6��v,
;c�6���*�3�/y(�l@W�2���"�U��M��i�o�~��Q���>ZRvq:Q~�x�c�d�I�j��O ��_�)�#����FTMU����#����l��ew��ʑ����>���QoԹPFh������>��l�.T�oJz�vҨ�/oL�L�n��yny�ڗS}b�uWE�zý������+��>U�y}{���iʀ�ب�zg�Io�����^�{�1MK+��q�v�������v\؊i�>A��Ty8��MYXn�}(f�� l�G
��u+����T41��v
�"5Lj������Mb	Tɨc�0�l���+)��U����BXLi糗�5p�:n뻒0gc��F#8)�p�b��M���e^;Ucv��9��y�F"B|���Ǒ7��L�^�gDq��I����C�h���4x�m����=j͡h�zjұÝ����휱���ola�\�9�赑�n_��z6�)�S��ٵv2:r�����T��̆Gs����S�����W��F��C��܅��˜O���nr4�D�s<1ȌY�{��_)>����LաE8x���
m���V��&�Vg��ׂ3)X��,�aRQ��8�cW��[�r�h�*�T�JXܬ���ؗ�t!Y�WPN�"��$��oZ[�tu���9=W5v_m5`ct��tb����u8#i)q��-Tjl�e�V�u�KV'�U�긖� vS�;n[�c�k�k��D�;�.�*-c���"�l���2���\%^Τ��j����躧�ݑ5S5����<�x�ە���H�Hv��n84��i:;Bn&�J��J1֑���U��R�l�=�W�a�:c���`�b���.�:��u�S\�.�o6�}o��޺�ҡ�J��\д��a{{=
C�umͺ��s�jm���]�B?b�|��WV)�����N`P�D�C5�܃�Йʖ��Ӹ������B�}�2�JQ�H,�:f����M=8v�v'aF�JJǂ�F����c�����ivض�gs8L�|�1��ۮ���
���EŴ��N6��	�}/u$�u+7�}M�͠�M�o=i��Σ��;�OW}�iɗL��`/Uv�n�J�STZ��aw^��cGOt����R�i��x��dHAg��$:���p�K��M��
�C"�꧛��n�A?@�s��'�@��������Sݍz�`iG�jun,hGg!�Z`���ј��b�"^;y�2�7v����4k��b���WJ���v�b�mĽC&����D�C��wz�Tߗ�ydV;ܩz�j̅x��Ϯ�P�ʬ�B�ZY^[]��r'|՝|��@K��,d�{������X�ׯw�lΦ�Wv����W�swy"�=��PL�s��\mdK�e������o��PZ�[�R���5��od�r��ȥOûV�>�����	��*c%��[p���	:�f��E��hTF[}֭�t�;79.�a��l�9���`/�a^lM��sf�X�Ϟ��H��y%jA�3�Iy��;d-�4�B��m>�Gy��8Q����BQւ0��M�;(1� �ۓ�ʫ���m^V��rCi�&�E�n��l���
[I�<S�̀(Z��&Y���CkFQX�\]�r�>l5֕�Z��W5	��Lt4��0�jܬvvF����l�6��q�5�#�J[���\�hk4������>3���&���yG�aߡ�zԋ��ޛ���p�����f���5<���ү�OS�r����]e�彳�Sp�+�9��<��>����CU@���}*�]7}�T���4\
�cqYO��&e&�d�sR��S�Bm��^|���xmë�j�1Ӳ{�����`�ZdHA3���V*�Z�FV�7��!Ns�]6힧a����#�emF7��g����-9ǩ�r%��b_uf��~\%��2��`�h�pL�mM#=u�H��v�^lٸ�-�v~}�;�N��s�Ju ?t�"�4��^ε����}-#Q�G��MػYW��n����do�xb�\��jW��2�k��S����[y#��i�����
�חY*�Cu{i�֍�$I��N����d���op�۷Ԧ�����Nwo�)��Rb�˛���J�6���w�I_�I+9��V4
y��Z��dJɕU����0k�i�[�8[��r׏�˽^������[�"0�օ�'�)mvU����ՙ3#NT\h��Ћ�)]'�s�{SȚ�v�0󥍫�{y�N�6�;Z����kj#W��ٖ6|�R�~P���)_�t��l�����dP����cy�dcJ�-���2v���a�2[=�&�,Q�N��N�ʜ�����*���D1bH��v�o<z��Ɲc\��ƥ�`c�e]�N�4��W��<�n8ϐ�X{r�Wq�m_.����TY���n�M;�'��l�~��ó� �tALC��5�{JؑXT�]u۰�BČ��aީ���'�Pz�k֕E%��4�4cywyۣ���G_5��X������5)����ȴ���!��@#�c4H��z�B��c��E��K�`;�|B����QE�������w��]C�:��re8���`�n/\2�8L*�ͅ�k�<�I�����߅�!m#� �s�fQ窊�z�I��h�F�Y$�X�mi�*��4�R�A.-�CV�n�h���RǪNP;��J�p<���|�� ���}�F*�1X���g��Dj�m����ɼ�z��>v��b�2�A9���|ú���$��F���*�1�8\
�i��vp��9�,m4��N�I�B.��S��n˅�9�X��n���Y �gTi"^C��k���������\2,>��DD/N-�w}�ٝ����Զ)`G��"
[�ʂp].ZD�Y�]�	��X�����WK�v��S�\yH�K���&�
�o>�9z�>����mܬ#��+����C.�F˩[�o�hU���H������a&Rs��$���z`y�U����a@�`�N��X�fq�r���w�6Β�ph���a��M�BE���p�|�W.�+ύN��lЕ�"�ಫ����)���},wpY��q���Ś'&,�Ǌ�vZ�JΆr�$w�Jn��5	���9n�)F���%kL�r��ᕯ�̀e�+�,�O%}�vi��ͭ��Ҏ'�m"�'��Di<h!�[�_'O%ɮ<r션�d�c �j���P5e�g�ks���^P�u<9��m��D2�4~���K�`���ͽhSa���
r���d>=��Z���0��h j�s-�`ńQ��C�V�IŚ�Jl�ah#�V�c�X�x�	�z��;���w��mB����NG��9���T�ܫƘI�fa���k��k7;e&��z-��ysø��87���pO|��.�w�O����ʉC~� �q�����&��)�vq�
O`�_�o�.l&XJ��Fk��7I����~h������t��$�B�+�:]�@��5��:�ڱR�+���C���b(��.v��T	�%�X��#1�{Z;�
�-�G:m�a��-�zIf_Dh�[����'?��#�8g-�~�11����V3�gN�~�n��u:����<�}�DOO�n+�|F��x^�j��GR�gOs�c.�2'��mU5Ӓ�?.+�OK(݁�S�[���
:V��ݣ���]�����{�u͝�D[��ڨD�e���0��.ܐr�˫�e�@i)��4	�����QKM`/w�분�]۬J�ъu��ΕbOt�Y�ն���Yg�0�gtH}�ʝ�B����J�=g���+���#��ۊi4+M�peu�lu�I�K�ժ��/�-f%_4��(e��Yz�ёj*����.�\�Ht���ܡ�����[+���}�ް�����.�,��J���p��y����w���EY�ʬ~k�eUbV�nfL�26�R�p�jR�2�����ʕ�V%kS�3�V��嵨�[Zc.
��qR��E1�fQD�+[��R�Yil�XQTE1+i`V��Llb�.%�
���ʃJb ܴň�)-�4h�9dU�����(²��I�T1*�"�V���1��Z��mQY���QQ)Y[U�(�11�Db8YEDPq�*�h�(��m�am����c2��j6�T*�D��)�e���0L�QLV�nT�U�ܸ6�b嶫�+�Ab&\LT`�%j��EQT*(R+Z�s0�´Ub��Fj������kb�jV�����`X��PF�6�\�Ĩ�֠���2�V���VҢ��1��Sq,L��Ks.5RҊ�.R��elL�W(&��(/��((
F�{����^b�a�����g#.���⻌��N�9�-�;���'��Qox�~�T�Q���n���oeL�2�d�$ugM��zq.]��SUP��sb��Ƣ�a��m�i���M�*Ǩ!�w;���c{�:�ݡ�mOxCA�ޫ�]v0���i�W�~͓!:1X/�Sqb�mV�B\@��qSj��ɜ�̥D���-ߊ����1#�?m_"��t��T��6�+_���=���|���5m-�-��&����|h�x�^�K�W��>��<�l�D�uy#q�_V����>�w�k��=�Q�0=ѬߠF��+Tus�ْ��["��}Hm株�z�Y^n���ȗ`�Ю�%J�*0g��,'�B�w�ɧ�=Qò�i+��ۧ)���%e�J.����3��{�'L�u#k�:{@�}W+��N�۷zt��S|
R$N�Z["��Ǘ��c�7�Eف��*�=��M��/LuP���6&E����ٗ������M�!H�G޼"�_��(�zI�0����vb�fȎ��ҳ���2�ݮ�X�KyY���;[�82�{zv�kU�(�w��h�v.����a��Vͅu��y�`�+�}�;�����E-�K&$:;�iSi+r�ێȠ9q��i6�@:����跗Ts�w�����\���h�4wB}j���1�8tAt�:O-ZńoN�mr�]�/��S����]�VJ��闝SM*�eͅ��H��Z�d=�}V��OбP�ل��U�o�*�u~����V��U<n��r�b����Le���׮j���X��^��ݴ�ܾyk�R�Z�M�%��6 ��4��B���>�!�+��h�F��u`�g��Ǝ@�M�CN��_9�Z�����^�O��YY3Q��bW�����ʼ~MR|!g6%4-?{���]n�*7�e[��n뛗,��u4���D��}W�I�jX�Q)��M�Ey�:M��Q��n��|�0u0}7֯]�w���*s��ES[�aB�\g�~ <�>�T߳sJ��f51TE.ҬY��nq�[�ws��1�a�HqNa�O��m��̭]}7��&V)�-mݽ�.ؤ�
���#��� �b�[�z�#�����ߺ�3$��&,�p�_H�`K�c�	�<�N���?tM���?+�s���xc���bq]���{~�AU��ZKg)�	�[{N�[S��bzѓۼ�u�4ݔ',`�"�s"����͈{��W�-[;/[sɇO)�[���)�J��}�Tϵ]�M�]ny�9����z˖�ͷA�u�����V�C#�1���'p.]"�[�UP�Eꄗ��I�Î�aF�m��3C�p����p���k[�s�w34��_Rw����+�4y�O�YT:����3+�,�Z�r�%�遃�.=I���5<���m*~g�F�e�c-1��ɹ�O���L*_��xf��'�z�0����j�g[鰯��z��t�;y�-��7���&�*��/lu	��CUE�nbp��MԾT�ҩ��m�H��>m]K��__���i�!Pθ��K�E;�᥮5�O��#4�j��O�RBM�K)���n'+��ҧB��VU�cݼV^�۞���Ξ��>�΄�8�uE���_�༊K9K
)��96\��2�[ɦ��U�NV������6Lc"ٙ�xd�bS:��n�qV�*7���t�/R�9d)��w���i��]a�T!�v\؊3(2�*"9B.��׽9�f%�ą���:�it�˄��ܦ��.����f,�]!}�쬥ٰ������o$ZQ>�ۚ���1�͘�>"j]���jxίo�91b��T�%]Y��M\�v���v��i�]hB��l)/)�i3�x�V���U��b�j��dp�1�Jĺ�W{M��3СOsD�5}+^*3-��So+�k��=�����ё����;jյ�V>W.�U�1zx8��c�\���Mʶ��x=����O	��oWJ�fs�8��-�]lK�gd��\�t��tb�����!vƮ�u����A{I>QP:�E8r�F��%����Wۧ�n�5F*�euيξj�FFB~�#r`[�����^Τ���ύ#�DoZ�b��:z�U!xeiQ,��v��ڸ�pD��4�S6�-ǔ�H���]�ݛJ߹�n�nU9�y��\C��EƎ���9)���.~WY�^Jb�"{����Z�2[�vG���'��\gV�<[,�V7�uKB��J-���kS�V��q�{J�
[��D��W��;!_�qC�a�zP���g�ζt>{���k1���g�;'�L�kg��6�:{�\���;��j�`�Ge7�:�ncq�U�n��M�^��7�@'�PU�ZU�/o�=����3�r�ל��\fK���<v�ՁM'��u�V�@���� ��Y�2�#��C�Z�j�����8Յ��e5E��76 |�.e	��Q�y�PS�>�c��U!@�Q5��������+�k�0R�r��r�`���L�f���J�~��n$Wm���l�Ӓ8Z)��rGu!�9=B�h(���bxF��*{֯]���p*�_?w?!��M5��jz�k��EƢt9�8d��.�{Qjb�eUT����Ư6��ʼ��7ea��A��g���՜}��+�]>��	��r�%>W`P�q�/^�	�qH9܎��(^y�󞝺��<�v���K��|�Q��~��_?�D���#dG����x��t����J�-+�i;R>�<��t��G7Nթ�`)p7�]˸U��	Du%�%�:X���]���h�AP��������ױ"xV�έQ���j������B�1W\�ȧ�Qò�m%x�7.�eI�qq1f���oL����u�o�
��.[���}B�ge;���s=����m�5S�et�+�Ό���������_�ϳL�gJ�~pj�*`�k9:��ӽU�3��%�+��\���E����Y�����]qv[|�,=�v���.��4{;�	��ÿ1��tT���y,�Y�7�.������"5�%[=��u�u~m*��y�4ҨR��ɥ��.��Rk����9��x�6{U�|����=T��Nh^��1ob��$�.5K�'��g\�	جUE��5�%wRű��B��UZ�q��k��7X+֙��{01�b�H��QW'y�Y����K�-`�6Q��:|��­�J_=�k���Ŭ����Z�%�3M��%��c�����qo�c�t>�
����ֈ&��]�i����l'��iu0c^�!�3���n��uwh�Ҽ�R	��S/4IJ����f�%
pr��[<�������eR�yz�ΰ������c�:3�co�BݹΉ�hȘ�3M��c�1����bd&�;.�F"�)�hĲ���rR�>�7Z�W<�Vg��v&�ڭ�m� �mD��Ksq�|NeMmྪI��z��7� ���FcV&��W�HR��꘺�N��N�ӽ��uY[�{���qwJ1�+�}Olf��^�v���q��D�Kc���ݕ��k"h5fP���Qp�ng������Y��[O]c�!ݕ�X�11��>�n�PoV�>��y�P���T�Kv&���1ϥ�]�O�MEᱼ�vS�ۯ9m���.�~{�E��1�V6�.~e�{�wn�A�a��KIg��v�Ҡ�l�$r�;�"�I�����6,T'z�9#����CW����>��>4�cG��mʾ.\lh���dz���yBhKi���w}�=[�&=�z��6e���l�Tp`ŜH�i��u��'#�}��ұ0w0",v+ᝐtԋz,�2 �I0nJ\-�7ݧO���Y���"�R�;�%j��|qu�+ЮhCSX�7y��<�ˉF2R�T�/���Ʃ0>�q�HȮj�V�ߝ���^���C;b�ί�\��?o;�o�d�l�����U�r܋��`_s͝�N���]ܧ��[��2��E{�����װ��s������W�LZ���%ub�*�<��7YB�"|�0Θ���wM9�Z������]P+��q�v:�ԗ�ߋ�A�e`Q�2�B7�ħ��u�蕹r6���y����_7��wV!@���εnOh���>�Vj+�.�^+󊽩�m���^l��W���/k�մ��8-��n)#1�G[�M�+��j�6�Q5�k���;�:a��\�ݪO]bU�MQ���8c�Fe+�J�ٙ�L^:������Xڦ�j���z�׶��F3kedF��;��{�y�q�>#�g�5��)um�#+hܙ�����q1z�4j�=�7���S-\�B�l��ۧt�!�s;w�}K��8��������=��5����Ng	V@��f�u�OA��|����Ys����P�pY���^�@$s�/LH9&������^L�u�典0�Sk6��Ț��<%].�S���^NN�9����Sj�����C�vKV��n���s�����1��#NC�d��*��hU����u�*;Q�����ԩ6͵Ǻn,B�9�-sO]0TZ��lu�$n\{Bg��}M-�u&����-YwJf*i��2��K�0vBG��:����f�L:kE�>���U�MhV���i޴�K[=^z鷰��L�G �!�S��|���>zb{S��/�6��O+�4�uy=*��sBҨ��{z���Tz5,S��pu�g�2d�:���;J�ZN�Rt�7���(E��^����>�S�uM��^��+�zq��됦��]���Gu��y����=�D��yR#qP��Ec{�����=ԛ�:b�O&E��e!%���b�@�J��t?��
�]���8��X����	��3��KVWN�*��-y@�����:�V8\��	H�<u�2�3�O^˼S;N]��xM��X��m����{f,`ҐRʌ�U[�j���(�P����&�gB�_�k�t�64q��,�s�9vn����t9��,�Yk���>��M�.3� h�������)��y�щb��~ǔ��:N��a��d�n�)�dp�C����RO�fB��ʥus��eo�
m�=�ڰ�L5F�+a���n��
�Z� �oH�U��ʾ�6�"�w������+V5�?�黝�,�½�GԭU����J�92=����I_��hb͎�b�<f���q�z���Ց��x�
��.[�;=W��cn肳�����s������[���1g.��o����������4���!zUO�r��O��<<��+SIXV;����P��*{_+���a��ח�qv���j�e�/WEӯ���u]:��&�=�$ I?���$�b��$�8B���$����$��$�	'���$����$��	!I�P$�	'���$����$�	!I�0	!I�H@�XB����$����$��$�	'��$ I?���$���$���
�2��H�hG��������>����1�  NE*�� ,�EH�)UB*"H��@��E �  HQA�%(�P� %T�*�    挘� ���F	� �"z%)Jj 4hh�ɦ������c�2b`b0#L1&L0j��	R��bi��F@C�hɉ�	���0 �`�0�I��F��O�4h����mM�2��������w�p�
��hh���'��@�(*)� U�?0� �����I�IAp�c�HA�
��Ai Y"��Qq��5��w@����O�V�*,[�U�M~]4.�J����ǎkBM����ZX��h_�y�Li�Z]A���ӕ��'r�P�m���.��*����͒�O]�"��k�%Z��]Tp���bZ�%nc�0���^�`��2]�{`[�m�b�l�S�A7�]�ӕ
f����&8�:�^��A��ҹ�Z-�#�T�x]�y�i����]k�Z퉫R%V�+w^�A���`�,cHn
�kT�j4�i9wT���N9�x�&e�yssr�AV��ĉ�
�ۨ��zj�'N��/sF�U`ݦ�:����bڭVN��4nMz��խ<KU����- �P�kJ�cl���6��U��-\�B�%+���O71P��+VT3��O"��׺R�W�QԽ��:7.n����p���b��vD·c�m���]I�Wd����f�ݙ�s1,�۬r��ZUlw7i-ͽ �x�5b�����L�wmob���m����_w�����o;mP�gT�@�UB�ۙ��\�U��5�ՒZ��m���-C-�Xt�RN�mZNB�qFT^ �j�hnIT�Ԙnt�퇱�
$\��e�.�NwX��V���*�GS�l�uw��bcku2�.ef��kk�VKo*��4���{X nkQã�1빖��;v�02u��Eu/{k�<�sxN��^B��r��u�v�ĺDo���)�����lW^!.����de).%S��ȕ�5g]���f��fl�i���T����T�ڂ�8��Zp�Рݩ��2O鲒
��q�ԥN\����"�5M2��qb7�!N�Dꫤ�Ӷ�o[S�U%1�� �:���������y�`���;���Az�TN��;�5'��%*�x�� p]��8K{��i��N�2^�y\�%�	�t��0���;4&���+��N�n�oi�E�r��������#�t~������ +�)��� 8��R�yK"�����o)�]gL����J�*��IB��*a�l�p���b�3��I�����t��-H@�n2$H���DB."�M�F�tB,���תmg��(�	$?F�:W�Lb!�PQ1H b7E3T�6#��.Z����"�
6K���T�~�Z�n��b���V�tѠ�}TI�Ŋ�sF�� �K�tŸ����/�(Q�BjG	$��:i�R��Z����C�XX,�?�H*Pg��,�ׁ�Y�~4�Ħ4��!��� �r@�U�B̸�Ʈ+!D�8����ѣgH6��	%�?|�A�	?i	���$B'�d�	
,�m鲉?VS�=!5����l��44Ơ�lR�):�|�e�F���/�Ujb�i�#��C ?1kc�:[&sZ�J�y��$�'؇�އ�Q���G�+��q���L���.$e����J+`��˼t����wx)¶�j����淑�+�$��5 $@	@j Td@�4�Ӎ��;q�-�����C{�Z��S����'���qML۟�7P_�>dO}&���A\�����~[kĕь��@9
��K�v��?<��g�����$��$36B4��+|ǏW���+��E�@��>'��F�$��}P����;��M�7��޻�"��H���'j�]=��͸�|*�
j q�5:�n��21K�Cg�����^�A�l�yv^�E�/ �\p��	 I��\���ݴ���h�Dlt�����ݘ^[�Q�*�űq�J�r.8r�.в<-��,����sp���7c,�ķd��)��&��+mh������(4#�CJ:rk#yKOSe��⦝M:���_Qչ�����yx�#�e� 6�ur��3p���ڞ!yx4�x��C�<����B^�+R&xk�K��~;���
�U��x���h�7Z�櫌��|�uF�Q:3��9.�h��[�(�l��|=�{��A���M�m� �%᥵�E&�d�A�5'SE��v[u���$[}t��N�z��/��~��C�s��]�j�I�ӹ:>;�8��*{f0nΈ�ˇ�:;�I��k���b���6cVz�ǮAo.)(G��i/k��#��R���� �ȫ��!`��;32� ݑ��\\�i\]�m�'��r|g��կAƴ��J�7��Xo���:���z�ߑ%D,�}u `����^F���8�\�e��9����;�3�?3������ծM�
:QO�̖~����?��<F�	p'������u��c������(	a)@�=,���%�)�0p�	�Κ� �s�X� 	
7�ݲ�/���1��1U�sr�{G'e�T���-�x��=A���`��o+%s��߇?]ph��>��W�G���."�b��oeA~��6n��p,�L�K��ƇJ����^�P?���Bd/�_,ى�*c8(c>+w76��M���h=����	"4�QyPwX�v��Tv�`��]<�4�-�HZ.J��+q8pF��0Jm��7�/��N����0b=�Џ|�???w��F��`�֟���D�S%rU�ɕ��Hd����w�/���Љ�{��p�r!�^40��{,�L����'����O6��f�@�SbT��
��W,��$ϸD�A�N˹ݐ	��h��`, ��Ƴ���H��\W���=J�}��J/�ByW���:�=|�ul���IaR@�6f�NM�
;~�S�]H���"��K���3 �t�UjI��6 
���\2��Tϕ����ǓR�ag��R�oQ>��6��:4����+2��w� q @T���J�����L�N-�o���@o@^7�M�Qt��"@@�*gJ@
�@A�-��{�1��b�8�g6�li��'� d�]�`i;��,��fgw3ӱӼ�a��d�u��T�u�g�#��~s �T��/ݝ���K
ta�T�k��+ˉ���g�<�_K���=��3��w�$�$�.�����ɔ��Qf�r���&��>�	��^󇃫)}=�ۀ��h�7��.p��A0�2�ٗ(ۋg��o�"=�ů��_U-��j��Йy ��(��-���S���5��f'��k-�Q�ӱTuݓ�	<�����Q�-o�г�Cک�|�a�~��7~�*⢙|j,���ocZ`M=H�bH�!eP�ï7I�ms
g [��� �Q��k�2��T����ڎ|=Z{�i���9�[}�:/{��8����m͋n�?\����;�sp�@��gi��v�Q�hw�$s�v{w������f��!�:j,+�u�R�)�v�y��=�v
�b^����B��XH����Ѹ�N�U߽��C��=�םQ/p��pC���Q�s�I�9���v���q]r��wګ2�6,�[��j�Iԫkqc�.�u�N����n�~���ۀ���p�i*�Ӑ2NzZqsX���X����MЈ�sTu5��.��yݿ�q�����j��X���p+!_m䫾�O��7]C��UҎtsK7�Ȼ�?;��]D�Yү�#
o	ŭ}�B<��,��7�-�3�ac1O_��w� �޽�=tG[����G�˾]|�}��.���F�E^LԬ:��]po.(�
��yu}�yw�{�� �~W�9����A�r�B G #@_�����ǂ����ވ�}�?�����}W��f	k37+/R��0��������[���'y��Ư��"�����)�(V@�ھ�O}��z�J������Gݖ�=�����5��$�q�'�}�{�;7}3Aӕ� �h?�QY,0~�v��f�����G����|_;�n>ی��*�*�,G�׫�����(O(k��z��UxdP'dDĪue�Z`+5�p�1�e��$�+1�,*El�]B�P��i�J\4��ZY�U�e�J�nb��f�K`��Z�V�c��)�~>�G����|���=�B�0E�Jz�ĐmVd��&���h���ѡ��]��y��}r��kg��?ረ�S�r�l�2�K��t�D��P�uuhr�$p�׍uA����;�w�s.rj,�b����KM���#"�Kۅ˪�e�b�^r�g'՘f��ԡ¨��ۘoy�d�d�{#.�jD�6�Q���=9	��f��MP=gB:R/9w��������@?W�������2�_B���[3e��<������i�]��=�H�;��˺*�N;���v��yJ�lKsKTL����y6k�]��e��h[@OD���z!�w��jx4�pD�S��\p��|�v6K������DQ��3kTP�q�b���ݺ�e��u7��k40�\&�.�+m��ꇘ],SJ{���z=由�D�H�����}��I{;��*[�gh�.e�쭔����6�&�����/T���+\'�v�3b�2��mӌ�k�jcr��NnL����N��*��pz2M�5� �I��\.K�<��t
�ط�qJ���8ũ�.y���l� N��nc���Uh,�A���q�;�x쎋�s�z�i�����]�zb���H{t�\Z�%z�]��*�����듵#�����FR]�Hw{��)	�����Y�B����y�km1���l	�	�MD�E�B�K�X��Mu�x-��hT�oX�b$�!���%�P�)h���O�r�J�콅84m�<��������gLl#�(��w���a(�&��O!6�bs&5W��.7W�6JN�S/[p�JRw�u�ynQ��!޻L�o%�0cN��nz=��������AP��xP��w�"��f���Dox�ޖ�q�P`�d�P�	�F���"4G�D`��y���{�s'2+�4��s�ｕ5Ҝ��Y�,�����doH�T��G�c�3��=AN7'��Yv����� �#�Z m1M�洱x�q@�(���`�ŴM�D7�f��u�i
�bVu���q��/�������H߽�B��57��o �
i_d)��av���S��z�>5�n�Ogq���@Ҽ���0�m������R#7���ܜ֊�t<:P.�#W�+�g(�΢�oH��l+�ZWS���Lêu9Y�iB�R�}�'.���d���%���{n���Q�������8�i.�y�}��n+'��};�`࢕_il���L:�Él�7�j%���4�C�y�+F�紷2�Ꚗ�e�qƘ��nm�}��ج��Üd�N�U�޲�N��-�S��F2KT苬��yMޗy	�ë�%���]���G�yoW&n�ژl�؋I�P� ��eJ�lGfe�G4�iv���1d��ɸ� :�fC��N�w:��[3�������wZ�.��T]m\ͦ�5���&L�\���9��9h��nkռ�����y���z����	1���>���\ⲅ��9����y�9�s�:룧-�S�jwV���"�"K<�i���8���j����Χ�A�ʹ�_.5U �f��,@�b�b�G.���ު���;�\�.&�|�)=z��w)# ��r(F,{Z4
K)�H�f�)��eD�9b0t��1<r�p� n.���7�`��l}��F�+yv+h��V(-:a@ЊnL�8R�j��mBqj��\��7n�Vm����&j.d�d^��N�Si�^����'I��h�ا
)�oUlc�K S%�7X�FG�����<��,[oTh����$�F�PSn���bs6E��������cZ��/���*���R�\	�郑1EE9�Vzw{;����I�	��r�HS>^�KU$��(z�O/9���"��u�a�扴̋U9%́sf��<�_*��	�]���ޟQ+s'��6zffP�0�:���ṛ++����rQX��*	j�5��m�Gݔm�#���󤮗@�	h����8	��\�dtI��$�</�:�>vW�ꤾ������.�&4d�u_ӯ�,���v�ɳ/�G,����w�rüC�,��Ɓ���$p��߮3�ϟ�&�k�o\u�W]t6M�S��n�D�$�I/2{�V9x�J��YisA8ٔ��#�Rw�T�u"-��nj���A퍙����������t���D�$�J�ҏO�����Zr"���BLȭl�MNZ�Z����,ir�lQ����֎�Њ�hH1�t�-�����R�h>�
��zJI9M`�t������/	�׌�Ҭa/~�	c�@�˯뱶��q�X�x�Ԑf�C�˺�SMr
��E����.������/�"�UE������8�f��=T��]}�b����d������x(Q�梢���_����$���� ����`�E��N��f��JŠ��`��9������g-��H?��P��6�f&�Z�4=,��q�V�2�H�p4X�r�bkyksP�.<��C�֢��p8�WQ���%�?X�O>�H�6y|`s�L��EO�����G��{O0�9wiEE�c�3���',%��� �����4�wyx�cܟ��O�;ü=�s�F<�����x���)�owh��y�x�\6�>ć�@9*��	�J*/��~�a�/��()z��>r�>!�b�B=���谈+�;I!�lH�f��5Ec��5 Y�pM��^�*��aC8b�q�=�*�㩡}6����\Eܰx�^{�z��EE���
~���.�; ���}�ur�2u���N����é�Jgg�F���;8���� Oq�-�u�6O��0"��F�=*2z�}��Q{W�h�	�c����O��<�s�p�V� ]Yb羍��Ӯ���hw�����`z��W��kF���ӹ����ut�N}]I-ʻqr&��ըtd9��o B�~��WQp�Zz\!���/��~6�c�� 랇Ǥ���Ъ���Y�=$L�`;{hp�0�o���.<�H/�!�
 ��g�����H�
��� 