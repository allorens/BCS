BZh91AY&SYA
�݋_�`qc����� ����bF            (���)���$H��= Ĩ�H��R�PJ���U*J@��UCZ
(� PmK` owP����c@�jIT֕Vڒ�
h Ȥ�I$�JH�қE���BP�R�4��	ᠠB"��0dJ�P���J��� ,��"��AET����@GM"���$B���UJ�R���BȪ�����
($R�  �褁� ���w�[�V�J�oC�����n�bu�%�Fۻ� �����&�R�lҕ��]�z:���]u�N�
�b(��H�u��Sl
��I@ 1�� h�}K�h�nR�u�{�R�Pw���V̅zh��Ò��RO�9{iJѡ�/8� vʤ�'�^�ʴk۵�J
�N窩K�R
TS�$ ;ȃ��	R�	c�� =.��O8���K= zcǗ��6�\�Τ
�J��ӽܥ(\u��*����o "�^�B���餛d$���@QRH�҂({|k� E���*�U�w����Ƿ���A{�� z����z�����'��ʞ�m
.��� )US��xzRT�N���TU=P�T��R�$����@�{0{�� F��x<J���m�J��;��*��u�`��
.twR5��F�΂��[ew��v�M�S�Wc@S�<�AJR�wH
V�Q3�wn��
U��R �k.�\4t+�R�C���
Z��rW�����7
�=̑y�fs�T �˺DU(��*�zč��� 8P�R�z��E ��J@ {�=�  {Ua� \� �e` @��2 �K�E9�q݀���n�� 0H
��ED)U*��) u��;u8 
9��� �{]p� ;����X �6Jw  wR� �  m]pР���	RJe� I*D}�R� �^a��� 5K98 �  ;]80 gx��`EVݡ�(���t�撔�����"J��I}������@�ظ 9������  e  k�W: u�*������P(���         ��2�*��4�`2b0 ��1))J��0�42h�aCjy2
J�F       j��L��S�`Ɉ��#L@J~�)U@ �h    D�M�$����I�$�G��1�#�5>��O���?���f�f��}��rZ����/�����7���s��̭y��@@k�iA@EO�@U��?i@��O���'�?��������O�� 
�?�I$����W遁?��/?�?w�Ӂ�?{1sض��-�b[ضĶ1�[�-�m�lb���-�-�l`� ��m�lcb���-�lKb��lR0[`� �	l[`S؅1b��-�lB�L[b� �!lB؅�`Ŷ1�l[b�-�lB؅�KaLؑ�L؅�m�[�l��l��b�-�[ ��m�b�-�[ �	lB��`�`�؅�m�lض�,`�-�lض��!lBض�ؑ�[�lB��`[Ŷ)lBض�-�[�alض�-�[ �!l[`S�l؅1b��	l��0`�-�[�)lR�%�)�lB���`�-�l[`��-�lB؅�`��-�6�-�[ �l؅�ض�-�[��Kb��lXŶ-�m�lb���m�le0-�S ��m�l[b[ؖĦ�Z`��[����-�-�l[`���b���b�ض��-�m�l#�6�-�[�6ĶlKb�1��m�l`[؅�m�[Ķ�m�lB��m�l[`�1�-�m�lKb�؅�`�2��`���m�lb��6Ŷ-�i��i�lض��lK`��6ĶF%�m�lb[�6���m�l[clHĶ-�-�l`� �%�m�li��-1-�l`�ض�-�[�[0`Ŷl[b� �l؅�c-�lB��`�-�l[b��Lb�ؖŶ%�b�ضĶl�Kb��6Ŷ%�m�[إ�i��1b��l[`��ض6�)�[��`�-�[ �؍�`��-�lإ����)�[�)l؅�`��-�[�-�b�-�[�%���l�%�m�[)�lB��`��-�����i�lb[ؖ��%�m�e�m�l��0-��lPb�[؀�@�
��V�l c[` [؊�[b�[ ؈��B�+lAi����*6�P���U�"6� �
��R���P������T-��lm�S`S[b�[[`�lQm�	l` F�-��lm�lm�!l `�lTm���� [Z`+lDm�-��"6�F� � �(� b+Lm��Q� ��!lTcblUm��R0E�*��@� �U���؀�V�"[cBت�Bؠ�F؂�@� ��6�@��U� ��P-�-�-��l``����آ�؊�b[Kb$b�l@b[�
��*��Vآ�[`	 [[`�[Bت��P����-�m�l[m��K`��6Ķ-�-�lK`���m�li�l��m�lb�ضŶ-��`Ķl��m�[Ķ�m�[��`�[���b��-�i�-�L[`��-�`�-�S �%�m�lض��clKb��6Ŷ%�m�[`F�m�l`�-�lb[��-�b�ض�-�[1��`���m�l`0m�[ �%�m�[��m�l�`��6Ķ�-�lb���`�ضĶ�m�lK`��l`��Ŷ-�m����Ŷ%�`Ŷ-�a��4����V���U�� W��7,�YUen�E۩t�Ƶ�t��9n�â"������.�w�6B��Em4�R�l=�%"�ç�͸ՊF�T1�Eی�t�͍R+q���B�h�M�gaB�+�M8E�mL�9�6�0%P�%;x5$Š)�E�Њ��Ţ�	v��u�D�-Jf�l�d��ʭT5�F�Y���R��\�v��;)�X�+�']�AT�֒�E���[c@�:�z�hT( )��WVHZ�L�t����X��.���in�y�cQ����]�u���v*�շ��K��n�ܕ��v�:�wb-b�2T�L��vpk�z̼���-n���M�ȭ�d�ZlZD"^�x�
�T����U4�����ҷ�a��k����lJhեj�����,�a��p���p�/���]R�-
��㎈X���t�ͰkkS�P�-��֮����x�*4M�#ن�^eM˻Yd*ۭ����D��{P^
U���-�X-c5Mvy.E�5�ݻ�Tڴ��[B�2������ˉ��ɯV�E�YZxXUIVi<��	t�:����-�P�1ުj
�i
Og�����Yf�/]��u��G^�w�v�K����'&V[E:N���wr�j��^�*�t��#vj0XnL�iB�YU���T���Y�[������85n�G��e9�;"�(*S7f���q�N�AX�a��f�&�H�V� ���a�2L(Щ51n��wA���.��Ś!a��T�1||/_]V�ܙ�G����mFV�AԤ^�i*��/l��\I�r4Dr�J�њ/a,�㲁�d��Kौ�4�cv뷀���^�1��"����U��
���gj�s1�	Qf�m6#�n�k6h��g�+3h�Z&�$���.�oNْ����T58l,�9�*A���DnKF�J�4$�V3oѷ$�*�\dmF�U��4o!��
VP7BR�P�ٌ�z����u�M��r�E6�,$/7^ޙ��цR��F��g7m3z�S �o-F\�nKKPA�c�B�i�V�L���A9&͛��mE[��ǚ�"	���2bh����Wo�G*�νb�L��� ���z��-i<uXR�h޺J����F��-�2Ҽ������)�Яx�5b�m��IF�驂1C#��@�,Ż�t�d��`;�B�����žXIɮ�b��Kr�*��6�:���f�]ߚ��:VrZ����fÉ�A۴��Q�Ok*�s�.�f�5�R��e-a�Y[���Ǘ�K�ۧ�Ŕ��ȓ6:Y܌`;���TިF�M�u��Pǖ`yQU���U4��V;���l8�5�c���)d�a���nA%P�)Z���g<u�� ���B(���r��e�Sx�1�Sp�����]�&7�'�=j�J�J��*�`��
�d[d۽B;�������*�)�oK��UM���n7e�Rt1�(�@�(�7��6b���Y�
��\�%1EV��e���`=Xa�Mn�W�ՅX;�1��Vե藖�.�[n�"CE�h�.JV6�eVra��L�J�Icr;t�rQ���-+kD�b��z]��r[�!�7P�6������e,�J�!�B�l�3SB��z�nmӃ�O$f�T�h�X�SoPY(_���a�	ZX,�(�d@V"����j-;&��ny<���h�ڕ��+p=f�q^٭Z���c� '+ub���L&;لMYy�
x)�7��5)q��3%j^�Y$�[K#\{��uHc�0�W2Q��[Z�ܹ�̈5��D�j�dM��I����~"֝#s��U�����َ�޷R�1�Hu{�&N�̬JKfQ�"V�9v���]Z����M@d ��j(-yVd��#{2�U�o4�C��o �hr\��*�ĭ�,ҙhXٶ*�"n,@^�����cc�6He�;r��q���IV���f)�c���i�n��W�����(�.P����Uf�t��:	*)'����,Ͱ��d�03Q�W���YJZ��c��c��Zzǵs�4*�@ �KO(��tM�yF���Y1�0�q�kk&`����TN�[�J�=�3d�fL!"3T�v�i�ה�[��e(��P�W��-�U��)�$�uQ2���h��{��S�yb?^�%��q�zF�x��X��[�]����lj8�c3,i'��k1]jD;��cX��V�+&� (�M�e�Ѳ��S*e���[vF���*�H��ԉR�������ȝ4˂��b�gB:��ik�q�8��ZTtR��	�P���ݷ���l72�f�mf �]K�)�3�r����9���jjl!iMvRB��m��ĝ��Դ3FRPEJ���Spi�skF	��CM^�Yr23pZ ���9$IL�a�jeioZ��f\v��X4����iKʥ����FK��O.�C����+�/a˭���#K0�UJ(��˺̭�-�ǘ�Omi��f� �iѣg`�6K�-@ �;�K���j��S��2x0e���	{��"�6���wgu�c�Ӛ�*H�-\P!W�.Ձ��d�)ށ�����:Q0�pQ�q�����M���Ҧ����^��-�q훸A�C#f���[��/��%A1ᙂ�ٍ<9m���3T� ��7KZ��]1��,m��k*�4�5d�x��{{�D.��;EhѠk$��+h�^Q��-Œ��f,��U��3h�K3�Ti+mf��]+ͫ�$Q���Nc7(bL"��A�ҩ-��-���3P'R��`�n��J�wIe�%Fi�l����)�r?8�N� 0v�;�sb�Y�9Ou����j*:��dj�Z�퇔k7a�m*f��v��Xˡx�b��8aGuyV��2J����K3��wYM��H(�o@�XR ��6���h0J�sV�V�˽(�LM�K]�4������V@�v���"I�%n8���{9�P�v����6hi;��gsm�`��T#/%]�Ȗ�ej�\�̶���@+Cд4F���өCw(F��X���k	4�<�S+F`5�%I��w�3]�.�
�k4,ЀQ7�6��b��y�V�Zƻ��xњ&�f�	Xm#/k������X�e��q0O��b1����֦�(]��V�dܖ�֬@�z�ڔR0u1��knU<ȞG-���Q�q*�:x��v/r;����ic���x�*�A����7wu�X�Z�ЧN�^9�[�G�&86 �I8�u6���TZ9N�ַ��9��K՗��xl�Wn�kJ��� �Q+uͬ�h�)��s3�LiV �G��G��fai��f���J�x]!RB)�6Vn��F*�q'�oV`����ir�e��X�+ii����xܬǹ��F&�����1�&e�
�ӱ�£^Z%ޫY1��f���,�If�#��;���Q:4��W(73M�U%(�z%��ΝG)�
 d�����b��W�
Y��(6�Ƒˎcb�#$�T#dI!��d�R+��!�ʴq�;
7{w��|"�%�"qm�Ek��ץ	(:6�@��1ͭ7mjd�K+wKjí{KՏ �gMւ��	�":��-�6���h�N�Ԭ�)�f'����0f�E�0��YWh���	Jȼ@���j۫����n�e+Jޕ���A��ː8�1
իҴ�"-�jR�N�L��tb*��Kkq��B�̓e3��%����e�M��:�,�T���Wn�X�0�nY��u��Y��)kcR���cp��!w;l�ݦ�jμ��Ȏ�&EZ�H��ʹ�-a��XM@`�o  ��(�p�'�b�aQ�Ǹ,���*m�*�ʶqB*�4��1�{��L4��5��nK�t��g%�h�8TqDe+ ə�z�X��Y�v�eଽ`�rO	ez��	=������
暱�j�5�'r��!�f�*Ga��+�;5�WV��H�<���q����Q�
걷I�2ʷZp����8��Ք��G@2��24���ԏk2Q�w�Y�t��*��vc�{�[I��Q��cf���.�U�2Q �[i��t���۫k���̽EE{0�SkkV`N�J@��M/�/n�̺�e�I!��X����VJ�"Kqc�̖4Ք���Y� ��1d�K]��	O)hۂd���4�*����j�h�@鷁��mk0-cT�x���@T/ ��&���j�;.�-۷��/2Rx���Y5�Y12 t�2�G�oe5�G5��by��S�B�e�{���F��ܱu��Q�2�-��ٵV�R�+&8�*���(��Ēr��f\ec�N=�]�yV�[(��8D䥎]],e�y�.���[�R�^%ZŗJ�eJŹ�t��X��P�BG���Κ��if5djɈ���Vy1&�mk�w֩Aq姸���,�d���h[ضEY��֞�%� t(�j�f���,RCj=r�3lk��8d�Iʴi�ݶjKs|:I�� � �^�����eF��v��-�ǔ f��Z��(iQW��6T�Ƃ��6�[E��n䲳M�XI�ǆHj]�F�&�7�+�6�6�6�ܭ5�T0a�γ	Ǚ�'^�bʭ�#ZJzR2��[2��v���f]��0���5�^ۆ���2�l�
�@(�ܱ�w/^<�+)љ��n��\sc0P8�Ι��=�����B�ʕ5\M�ma��MC/}�xN����<F�T�pa��D;ȩ&X���[��/%��Ʋ6%�C]�Z��дpɒ޺F�[N+ۤ-��DP�,��6��b��T4�c&�����%y��rS�ojR���M���YjTT&9+.�f�(�U��MK�X��R �Zkbe�ҝ�u<AUض���^F�"��r�q����F��֜ʄ��B�q7xېb��Jj�e�,<ܳr1j�K{��C��щ�`'^k���CN*�n�ެdS�
�)RT��E�$���2�T��֬�[�Gi�ׯ�"ڬ�2��(�^���r�K
;[�e1��J�m��f�ؕg��x�Y"˲2:vΚ[�`�)�u��Dkb�'p2�c(�Q��J�0G^��n��Z([kVڂ�b���m=׳B�z",QQ$ó<\u�R���y��c,ڦ۶����wk+�i�k*b5 ��4k�GRJ��N�hW8�T)�f4�����V�f�.�n�p�kǛ{��`Ak%@��ӑ�+H+Z�$��m����9j��U<d9���!�]!Z�n�y��
FuP���9�^^�h�VN"LT�Zy�m���7vG����RlZ#�5n�$V��c<�US�7g"���C�h�g"�T:e�è�k�̷I�e���Ħ9Wx����L�������{%��f���Zn�褖]5�]f���xc�����j�ђfؠ�K��PE�����h�=��t��ܩ`���ձ��YKm��hm)*�n����;J���ڐ��ح*��Oӑ�0�f�y�N("p�lI���퍹��Ҷ������P�n��JfjްwoI8e6��x�����vXlo.r����L-�s�� q7\t��fe)�w@�ʇD�`�gd�3Me��ĝ�/Mcċ*�4]�W�N�P�Z���c�T��)�X�*�ya+Ux]���
q�+j��f��h�]_�E�栫 �ʹW2�NvN���������{{V��ń�L�O,6qS�#FmSy��o�Ő-R�dx�I�hfzG�.��V�D�iT7�E�n�QQ�h�1�2��o3�D�t�)E�s�kD�JӴ�$�X�5"�[k@�Ě��	x��[Y8Uh6	��.k5e��ܜV��{[k9,[J��o<��mO���_]�J�v���MZ\嘺�j湮E5n�$��Z����]҉0\W�V�Sr��E�W������-&�r�6z��sOQ��e,�v�S楡"�ʫ��2Z�NC{�6-ks�o^MR֥��A�_j�%���Vj:��j���_t�������w;�p��Q$�*I�z�'��i,wW�c̴qU��.���̺�
�Y��mWm���D���Wm(�$�Sy6�E5,&f]�-��6�B�^&�t\�t�����e�UhھVӥ�P8��z����6�E�kAu|]Eֶ�[�Z�K�k�<�j�L��� ��sQK�*O�m�4��]v�A�+T��X�s��\���m;x�����B$���&�1>���mCܡ�.ڄkV��-$�P٭;Q�sA�Z�j���6Mst��b�;x���q[r��U�'+��v�峂�Y��-GV��kM+���;��zR:�֥���i����QZQ*�Z�D����T����S�5���h��q4�O�K�`۶�(�.Y���[�}YoGg�a���(�N�`�N�a�X�W9i4i4�%-K��4�#JD�T_9��)^���X�`�x҅��O�bۃ��4���qr�h��(�,Jm-P�ڻX��@��,C#6��h�ܭ#��(�+�Z�V�jȜV�I�t�]KmWi�mZLi��Ӎں]k�]*ʹ�;j��OV��K��o\����:Ly}�	J��.�U�@��54���mp;ʢ�\�%֞��z|����ҾJ-k�eU�sN��Z@�#j�ı%��gk���#K���S���8���\����:$��A�:R����1d]K-bS����E9m�h�uC\K����ҠTZ�jV��Z�Db�-Q�]��9�[��]�\����ط5�MD�:`�����R�1F�k9o��m|������v`�Z�,Z�V��^ds-ZR'ʱ��|��ۘo��zlЙq^�\�i��T�'��a�5�0��!�/X���;�k-Ŵ���|�m��X��E����?���B=ߥ�~~0t�~�W�[35T?�u��}�mm�=g�������TO8��5������T��&\W�7�[u�Ͻ���^&�O�s�x���^N8�7�$���T���q	n��ay]Bȕ��.�k�;GX��r���y�̛�_k�]:�.n�v7����Џ�ҫ1�5c;I��x�aɾ��V+�{�c�1G}��yAS4.ݽ�\��*<*��m�nN:����׻˻=&aS;:�'WW]�kG+�'dw�T?#�H{��Q��a�;���H��%ε��|�i�;���F�r���l;m��׽&��*���uY��m�[��WٚD�8V[�Q��X���ٮ�JO��kS���P*�3�V%�8ଽ�Y���p@��bw��} É���i��=�JYm$���9��St�2�Z��cO18�&2fX�D78i���v	�e嚑c����}3�\�f
�P��0ӣ�-4��*re�
������ktrj"����vΈWS�hn�J]US�p�'3�v/7��Z҂������LGʉi�r���{�usg:���:ۙ�j9}�y�2��НPX1b�#&���w����^gP�ɛ��@E���u�͗�ާ���a�_��Y5yS'+��ѧQ�:�;�8Rv+���7L�mp:)��q��`#�J�Ybq�����닂9uº���l��5Tp�M�w�f��v�<I9v�:��҅�q#�����it�ct�w}]��
.�����H؋�!��f�p:O1˶\���rSh�݆2��gNn��˴�t(S&���4�2�)oJ�+��su��?C�M�8з1DLW�<�1>����uv;�E���]v���������oEy���[��bI �GǸ�5a�&檵��Z)�nһ�ܣǬ��Kielˏ�֊u�"�Hf��#�FR��R����)���8�2��u����yϟ^t��p�q�Y��]�ˌ�Oq�wCIiз�ye��L�S���%�ݲ�l�O��긦,���;�7���N�qޝgWf�v�(��ޮ�$��p��f������o���j��[�v���
�j	��-�*\Z7��,ƏX+���(���t�f�"�L��+];N�՘�J����u�)2Nöz�*��Kr�݉�p�܀��}o��<��Y��l�X�.�,�P淔�3n���qEVاYK�<Y�7�L�ҷE�M�����c�թ���Synk�Ա������1�3Z���k���g���7���4_bJ��R�렎�0����43�E�t�;A<8�J���uQ�d����r�:d��,[vx�ۡd�-��a1����%��;,@�u,���������r�5Tx�s�k,�Ewo{�S�]U�g �s��-sK�q��m�4MF��⮞�'v�8.қFK�tF�αe����5vlQ�+�z���6��g.�����
��{�k�L�p�g{V��4�x�Դ� YF��Nw�L��B��kKi�zn��&�������-�k#�cf,A�a&���_`Lc8��$���CAw� a�҆s"���b�7X��X��%�,���Ү`�1[�CiL��#��B��L��Rؔ�z'�m���{9�x�n�(M�GN��i�O.��E>*��7g;��We�9�6�
���� 2���{�1*E���n��6p��e9*i���u�1��]��1�w�X��wi�EQ�X"�v�u�o���	il�����/�����Nt�޵�K6x���{U�c���~�f�Q����_en��Ye0\d<����&���nŔsu�;Y�4H�{S<��j=mc���dNwZ�b[�C%���[�KC�\ѻ�/�c�J�w:X�;K��x�g-�b�Q�T����Pѱ�����y:ђu�#���Yw�y�}*[�(��tn�x���%̊��9LbfXK��ɹ���<�y�pj��̹-d!u��'�S����F�us�e�*��٪��Z��2�\�9aZ�J��={��t���\�T{>�1��mq�":5Q�<��wJ�E�؄�<{�ٓ-��fB�7��a�2<aٛ��h��f�l��dr�o�T�G��i�%�,�[��BR/ri��
ÃtV�{�����d�|8k�7����H�0F�����r�˜���r��Ê��\�]�.��fj�n��7�����+i���\�W^t�es�ᅠ�3͵�=�<�X�8��*su�휸�}7'u;0s�\���rq�se�E�;Yy�&�TY�����t\��,�:��P|@���b!.�2*���y��S����7G5Q����f���'�����n]F�%���9:��nZ��{��.P^�q�[clm����2G�K��~5�t���{���cF�&du�>CT���T�^��+g/CΩF����ȇ'o�T�r�޺�mR����m̺k��(��3�a{8�sH�-+�̍�����n���V�E���x�Y9_*Σ�RV:}���p����D�w"��҇�xor�R���n"�nRy�+�.Y��q�]uq7��&��ru���V�ږ��VW_+-q�D��&+	�Y�RI15]���c�w�-X$�ʎ'q�;��������Tq��]ȹ�-)�>���75w��Y$����s���R���D�dׁ%�����5�}��ݧݣ���H��i)Y4nu�j�����3��m�o�=n��YK�,�ǹ�6s����ç06��ҕ��7	�qkJ�zTV&>���rx��=������u�2dJ�4���1����6�v�GG��7���[�5Eۘ��x��\pJ�T;G����ԫ�X�ht�������5����)<�?>�7�����y�)��r�E���T�]�C��ԣ���^��NVK�4�:^ƺ	T/�I%��1���R����zz����qx�yON7&���`�\�8�{Jjo�,�vc��(f!x�L�6z){;�vH�d�:�ٮڎ���AG,a�1�CT�Ҭ�!:���nF�uS�1"��N���:��-;����=��VN�p�z^D�/#��6h��Y9���8{v ���dP|��+�fav�'*�E���<1���.0J�����)��2�p���ŋ�<�fqn�Y���m��N<!U�m���sښ(nL{8{E9.�B���76���oQm�D���Z��a�3���u\B����I���m�i��2����"�e�UB�ӍlQN-�B|q �[F�E�&�t!���̦Q�ks8�s3!��F5=�_U��\�= թ�X���C�\W��R ��b�$��\õU���bz�'�D$TM޺�u��6��a�"Uvo0kmqٗC��l�M*f��]�.෈҃3�&M��"	tՅG�[�cǔjy��-�ݽ�+�O�5�hB�`��up�
P��GW\�k��N�9�y��w�蓨�}}�)�r��*�84w��Je)��.��:9��y(iu���k�9����8c`w>�/.��ɐ9�N��c}� 5��	`<i��.g];��1�TX\�&vq�^�J�һI��`X��$��c�*`�y������Bv�x����{-�F�����L��؆�7mV�l�A���y%ɯ@:�hm[���&�t�5�U2��ގt�K������X3X3v�Ƈgs�xK��<��#IGp���w۷���uod��J>�g]����[�YY+{d�N�e�w.��)����\XD��ua�Lb�3Q�$Y��z��-���n�>9&���=C`�4X-��h)�t�ӥ[[ڞH��l����JwE|Z�2��0ǫ��@w��؎�Flnv��T�-�nZ�d�{�lC�QV,�v8_&��P��U�����~#NTIS�C��:�ɽ1WhJ�)v���nk���9t� �.�{FN>�ߪ�c�J8�5�[��}����L=��b�S��W;5�]Ab;]����ɑk��mѠ뙻.q�h��E�1T5f]ҽ=9�ή>��I��0�]��n��0fX@����x��֚zb�*���9����+|�#{{}WNN�&Y�Sהzm�p�=k��!ϟJ"VV�+��]]��El玫0��խ
�ɋ����ڌ��v��P�)���,�Yzn���3���hh�ض��,-��_��N���������\��/8���x,�+.#u#:�B��/t�4��i����8�V���L���T��s{�zj�m�t���������$g��u*���4��9sY���m'Cl�?�-��ca�
�G�O,��u;����ySF��}��䐷.��n�_}{��K՝�]
�j�p7d.f��ݏ6ژnԹ���Ut�REm3}I�FLr��.�KF�z!5��[x�Y��e��l$�X���r��I�ɔ]U�u)wI���8�F]N闫�L�W�|�D��;8*U��}��o\��ڙWOL���gW.��f�h��
���������Kf���=}�u�������;���uZ��bz�����rc�\P;��*f9� 7�\��e�N[[ӡ�5e=�\kE�L�q�Fu�>؅Z|��ڰ���E74J �Qk�*GX5Z� Y����td�}�'&����T�I$	��U[���캂�e� ��$Ḷh�G�q�7�@��w�X�h!���{E�{��u$x�o{��Rg��V��b�Y�p�X�w)�p����e��;m�ϻ,�|�$ee�VuNc%�hX#��,�VEתQ
BE��gw^�e��/!]P5o�f;���r���Yԩ'S��1�E-�v�9Ohԥ�N���k8�j�=���窮X�4#ӭwd}2Ά�m�Sn��ƨT��h.\Rwhm�;̓�������Z{Q1�%H��s�9=��q���q##��f
�s����Z��[���1�g�pc�u�l�r���Q�a��"]_4��.Ĺ����%��y5^�ާ����WuGg�l�b�|(��*��5�)�/(8�bC��U%z;2
�|N��Wөh�w+��-St�.7���xѴC�;��B��ٸJ��:z�R��r��jۦ�s8e<�DNc��I��ܭ����L�o�hB��	!k*�۝���l�;��>�'�.ڼ����H��EU���}A:W\���;+&�ָ:j��د3`�fWR�-�]�SŴ,[MSw�.��c�SW>��[�{���J��bkW:F;�U/V-�0wh:����L2�H\�/6����cWK��fG{C7^K}&gk����N{1뾸3 ��J�L�4#6Хj-5�\;$�	\Ớ��u�2]����p��O����KT��<�9�u�*���o13b�4Ӣ�[������.wbU���Vt7�DH�(��e����F	
v���;f��6yڈ�A`�.�cYÎX�[�Y�`���ݜ��Vѧ�6�����v�:#Z u�� \u��w:ݼt�K���v�}ؐ�Rm*��˅�oc����S]�W%�P&�6u��'˶2����m`�/�{�q�՛��.2�j9۵+�a�Q�����=�qh�����M�4o]뜻.�W��^^���i�n�<X�Ia����k	����q%S���SN�E���.�b2�F��3Z�]���L�-�c�F����zi��21�i����`�n˫'V�:�
��ZɻOU���7�s9�*g1��}8��siMe�+q7&mǮ�'��V^�{�ʥ�`��Ƈ>� �\_������z}9'x���s�ύ��ܭ3��GB�s�eK��!r+uu�};�G6o�%�$��B���qT�q��m�
�y��J1�K����T�;�wϺ֘Xl�uT�&=���H�]Bu�ˬ�K�᧮����@�T���;l��q���;�������W�{��;Gr��r�!�HJe�`\G"���!�Ԁ�J�|�@�����p�Z�L����{���R��C�C5{��µj޹�+�n	�V��˱9I�^Q+-Z��%� <��>��vc�� ����]>ME=��7��;$��	5�!�%E'��Mr��a��D��n��a���Z�����:�>D����DM{�ԇb�}��7��wt&��\)!Û�hG���@ �ܮ�4��b�Z�y�;tX��.��򒪎@|���y r/y[��\M�<���#�Qاouk�d 6J��w5�y����@���ET��P�)��7.t��3�����	ʐ�P� >�z�e3�7�mNC���?��t�(*>�����w?����T@G�������������?}�^Hnq�&���5��o'w�xP�Ⱥ�.ݕ}0�[�Cj���&���VK�6�&p[-�2�XZ�4�nnѻTCȫ U�Z��s��q�LQ�P6���]�^+!����� ���33o{Z�y���D����&��_L G8giV��Ν3���Rٸ U�1ez�Ѧ���Qe�u�mZ����V֤����I����G\�7Yڅ�"`OG]�7�Լ ׸a�BFO���F�elw�Ou8+WoBj�`�PFmIw�6Ւ�ti�0�'5\-�h���B̬2�D�n�8����R���_"��"�D��
���h�5��Q�u���z�@�h(���H�x�.>�霨�Q]��CQ���Ġ>�P���6�[V������ג��r��P��f.���B�]���s瓪�'78/�#�6s����{���iW1���X�
���U��]N�;p݈ZÝ���k"&�h�un���1��GO{�e��+�϶�	�l M2b�bH%��J�Vm4F��|��u=�,sִ�1n��6��3�0�e�JM]��Xy��Yh��T��S4R[0�v�ƃ9��/O/?u�z�q�qێ8ӎ�qƜq��q���q�q��q�qӎ8��q�8�8�\qƜq�q��q�q�q��i�qǮ1��q�q�x�8ێ8�<q�m�q�88�8�>8�N8��8�8�>8�N8�8��t�qǎ;q��t�ӏq�q�q��q�q��q�qӎ8��q�q�qǎ8�N8�85W&�5���u����.P�[ ��Ů�E��.�3,�<r�i�����܍+;�؇t8:
]�^������A��*D����v)D��ɗ���e0��ގ�r�7n����u[*ͬ5V��z�&�;&���vn����igv��R��9j�k�,�t�^Л��;�ȝM��cqN]ZQ-઻3Շy��w���F*<�|{8T�ͣtk�t��Y;2q�KY�Ml˥����:c!�kw�Ud��M�Z!zfhӽ ��=:�
�����]�dwVC�Y�F՜�J�9���ذ�I�hK�S�r��y�����v����_<n��퇹�5(;|z����=�9J�S�*�i�5�u;�h�,�]u�V��|YX�]6����.��"�tU�-��M�p����6��8io�Z�Osd��|۞��fU��c���
�w,�D�>���p��,[����۳�J��/r���`�m��V��ty���dSH�S����*���	��v�+&�.<��}[NRz�[4ݽ��TA�����Y�,��U�LT(�H��bRpT�k����pk��兙7��ޚ��q77�O�M�(��W�0_�y��Vy~s��jgz���q�qǎ8�8㏎8ӎ8�;q�t�4�8㎜|pq�n8�>8�N8�8��qӎ8�8��m�q���:q�q�n8㎜q�qǎ8�n8�8㏎8ӎ8��m�8ێ8�n8�8���q��8�8���q�q�q�q�v�۷N<q�q�q�q�q��㏎�q�q��i�q�x�6���w����{��H���'^���'Z/d���ز��:�Na�n޼�n������j��5[i���+NiҬ��lC%vM���s,R͑�efk�\���C��u�<��wu��-�9:FL���s�õ(OK���Q�a�n�?�0�����ۗ�3�T����}�b���gJ�F�y�u�t	���06����u*�IJ�ح�	��A@����e�z���t[���3�P��]�(��W�w���E-��c��l�0�%���I������9��i��\�y�N�����*��fq���t�y8܆C�����3�����gt���Ю*rwnm۶����>;�msǸ�y8�$��X=r��6/5�|;l�f;ެw	lj�O_o�O/��#���hj8�U�๏\&��Z3ln핔�+5I��6�U�X�{�"�_d�s��˕0�U�*�3fW1X�!��W��voV'j�Ф�!(�	���^r��ni\���ɽf��{YdQ����"�-7
���;EJڛ=��yέI�`��y;��t�6�Tי3�@Y[������s���0<�B��C2��
8	t-�a�YR�Y��R�T�^^�/m�Ǐ�\x�6�4�8�>88�8�>8�N8�8��qӎ8ӎ8�8���8�8��i�8�8�88�8�8��8�8�8ノ8�8�88�8�8ノ8�8�\c�8�;q�t��c�:q�qӎ8��q�q�qǎ8�N8�8�N;v��q�q��i�q���:q�q�q�q�q�q��qǎ8��;�s�f�yc�Hmo?t����7�����s �l�J��y����`N����]�6.��K;KY����3c3(^������[�ח��мO6
B�+�.�9ͦr�v��ݜ1���]k+z���"f�p�A���u9q�W�'�c�����Fp�o\�؏R}��e��\�dR��[��g'X8��_[�)=Z��ڳ���p�UU�9:�Ɔ�.�.�)�G�.
�m���,�!��t5��5tB�zxR�%���ҥF�3(���h{�F�.n�2V�^c�E2�dj��Y<<����G��\����}���B�\�����e^��|�3��aԞ>�t����h���)B����ʰ�c:�p{j֑�U6H��I8����{ΰI��UX��7:sy-K]xO[��W���7\:������!"Ή.s�(&٭t[}�U�+��kYxu�e��D7t&鬔��&������H��k=�����2��p�q.���Mpu��G.m9�]GӇ�rO#�v6�Lu\:��+�"ⴌ炔K�j��:60u����Y�V�ѭ9][������-�=�]�xˑvAؚ�ޅU"�U��5lRM::iF��}˕roWvIy�7���3h����ق�[�I���f�0�\I,��Y�H���;Ut9�feM�*D��,�c6s���՛���,+p��\_`��	I=�ɞ���˖u�(��;�˭�����ZNeu�V��X%�{G8�M:[feHͣ{\�n`ݺ���3v��,���B��%�p(>);#I�����c�L>
ou�,eb��1��
Y�2��,
��)�����yWQ��rn���j�ԤԬ�֊ZT��E��颮�u��6wiU�:ŠC�je�=���5($ܘy7���B�+e�^�[��=�K����;o��F���eO�q9R���vM��̡��QND���,�g4�.���E�f��(�]Գ���f��7�]Xe.��Z���˃�6��F�0�;�#�y)k��&�]�Jy�pIhލ����c���=�>���Z��ާ�z�,�ȅ��
�f�01Wv9�ٮ���s�;h�*�{rlɻ0xdwc5��E6;'��eM;�)��X�v.U���# ݦh��A�s�Ε+Cr�Ҹv�<=x��|���]�[W��(�g��:)����Ƀn�6Q�AC����.�RX��![y |x[1Pܹ��m��@X{�F��x��k����b�^�I�^���TD���ѷL�N�h娧>|t*IA�O�����v�gY��~ �A,� HI��9�{���	�gk�ԒwZ�ܺή���R{�΍>�����ޮΣ���X7�.��Kf$���ˣ�M#]!���ET*�h*�4�sD/|<^U���!��]��\i EG{�7o��pK��ޑ�٢��޼Dؼ���gs]��Ur��W:��k�"Q�t�ܾ�q�b��%�*�7��7Up��*���t@������ThS����>`�ۘ[��ʪ�őo�/0�%40���=����I<��!Dn���S�B�eJ�z(�\+�"G����jl}F��Sokf1�L��cPR���t��ҭ�*7�ƺ/t7�5v����1�o	���+T�����*G����j�8��*�҄gn\���^��1�m5�߽I���
*��/6:�xé>�/3D΢��L�CbJ+�^�^ju�A�AJ�g^��*��F���p�F+��Yt�\��h>��HM/��W\��ضj���pi*ʦ�i��)hP7������f��.��/K^��'S͌�51}�6xo�\��S�)J�(�PT���o:�T��ՅXC����5w�FT&��W+�pת�e�%١�D���&���|�ӹ/��)���[�k��s�pV��_K���g���k;"������0�9�X <.d�D�Ymi�p �V���6nd�A�/yKy��)r�]uҥ�ƖjS{`�l�GiA�=�vo�%E{�Ak�0*iˡ,�w���v��`[�S�-F���%�ˋ��xwLx��aǸy�:
n�uFRH_J�X+��\�S����RL�;yպu�>8�y S�����lq6�y@�V:�nMr;켝{I:ɢm������yZ�
�ږjlӝ�H�s�6Q��Ҧ���)!�{O-�:���茲��]����{yA���gp�i�A;7ǽ�Bƙ��B�6����-�����=��I ��,�G��U��Sv.LD��ŴKt���� Lw���c,p<���r2$��Ut{�Jre�v�u�8�zL��e���4m�^�V<�2����pzL3�_)�*%���힉%�[���%L���
���nƂ����Պ���;����:k4�Ŏ �Ӿ�'Q��Sq�@��7ܬt+������V��C��6�y`��o�K�Y�d����"�)y��iY����2iJ�U=/����ga�M�J��\��/��17�5-��޾&�C.�3�u�mN�Y��� C5��T�ke����{���� (H�x����\���4+=NGUqPŗ�BTr`J���k��&�O��؆c:Y�U:{�'`]-+�\j�-c8a�l��SH�X�6�ʛeҷ�'���}���TUhQ{��f7`�];���\�VmOM�EA�U����gPgl6'�b�kq+�)�Z.�*��\�_��z.ܒh��G���f���s�O���W$7�"rŜ����(�U!����غ�0������r4���^-�Y�u���6�j���Crc�	�uX��ǀѸ�x^V����df�L����op���E�T�ْ�	�z��U*n���c`�e5
�r����"=*�󽜥=Z���$z��f�Ҭ�#.�A�+!!�\�{��/B�(f<��˹���H&�������lX�wP�{�������NodC0B*�K��Z��UWW)�Α�=�,�o4�un�/E	X�9b��4��B��lX�2[�bΚxAo��R�+��<t
���e��]K�I5w�7djj�iB��7����Uۇ�����U���g(�**)mf�2 �����o������^>X�ܮ��w�d釨�T8�T�˃�X��÷��-�х�ݴ)�
}1z���dhX�pP^R�.�T2��v���P[�I���`���v�7�.�%R����q:�Ǡ.��aV�ʷ���@-�u�˧�˥Y�cU��j��l��*����9ԡ�sTu�7,�w��{��%��&Y�VA��Ζ�,�)o'�w�ϔx��I���A�N�Zf��n�]e@�d�W]t�%�y1��d�
�~'z+����^}U�C���'v�v�ǉ�tNVޞ�UE�t�.Kj��k�_�"��;A�2�ιR�U'b���|!(T%\�����I�u�bn�a��u�UGgZ��5p6��I7w5p���t^��V�69@�*�uu>o��17=b�X
֜
��Xf-W�|�L�v��=��@[��f��eh�>�ށ���6���9y:�yur�8�� 5\�
Cg��b�ų�0O������ٰX];q����H74]Γ{�{������N�T�ں�NXW!)�(ZήNY��LKU.����2��[��v�cʱ��[��"��r�L�De���/1P�"Qnjz�u;,��2N��alsS�"h,i�2��nh���@�S�#6��*��)`=�27�P9�T:�r��$Z��\���[��g�־��������U���
.����`��	�T�c��J�rѾ7�G%��qmш�u�sQÑ��yKu��-e�di��ذ�8�C^�X8bU5�|�Ab����.��/�WAd
�,%��T;����X�ZtE�2p�f�ts F1�۝9��.���̵����͇�=�۲���k��v��L���; D���
uk�Q����L{�ǲmf�!k.ӯb�"�,��[��r#v�Ŏ�Lg0��u<��;K6j�K�r��Kw��%��'˨>,r،�g.�0�����z6�R� 3M�J�m{����G�f��{R�����F����8��nj�w�p����>X�j�0�S˩�H�	�w�M��E��o�7��TM�.���GDGa;�\m&v���䋑R�����Q1����=tko(��a.��^���-�A67�6���f��7*G���)�S��5�.�j�3;�ͣާ!�+�s!�i)�=v�j�6i�,Uh��ya���1TƸ�(��n�7u|���8���x8���z��3P�I=�;�K���@�v�8\Xk�ҬīiK���ٴ�_ZGMM[t��v̥��\t]�i��i:���.�5�n��E�W0��Z��V��B���]�Rr�-��Y����[Ot.���Z��T�v5![{����ek�:x'�=*�]wt�a}n�.����o��&��w�s���˧}}��Sw�+#i��_z�^�ݠ����N}Ԧ����<�vs���?PW�?��~_���_��!��� #��������QF|O̶Ie P!0B)@L-0�e�b(�i��G"1H�B�_���N6��:�D&�Bd��J9uUU!aKH�p(�7h�dl��8]
b���KD�D���Q0��D���WФ�	0����A�D���N8�1$�2D��L	��(8�n6�e�
D�!�
L�Zq�˜_0H2#D�X��4�-�.%q�K	���۾x������{���>/{���������5��c��v/�P�u!J�L�pcU�*-_�Q2Wzx+�˱ʫ��9�<��ccz�b'Mv*Q�Wp�WVt��z6�%�]���[���M�O7��ep���r�V�Wt ���J�^��]���Y@q+5+C�G��sl���{e�	a\h�ё�C
�N#�Z���"oQ!&�K{�����͛�Z10=Y&�yݤ�g1 r�q�w3�rٰT<�љ/��T̻RwV�;��]i]�#h��X�2SʈXc�L!�d��U �f�ҭ�_0F13q)����̚������έ�+�V�s)7N��<i-��Wd�}[�W�dĭ(ϸ�=�.{�P��m݅���	�� &�-Ƥ0]�r�I`!H�7���`���F9fx�������Io�4����6��
��x��sɓ�S�ZF9��a�yy�;�6nh�.�{w:�p���s�zE\Wpn	Yh��e볼�Wc����"T�7vG�kgga����m�1��XE;��k+9�H�MaƲ���c�y���D�ڲ/��V�;{M��8J�xF�O	� Fc.iT����E,RLέ2
uU\���ݙ���׭�]g��<TX�w�������[K��6�Vd��X��	�;v���jB�a%	�|�	��e7	��!@L�5#!�m��a_6CP�R�l�I-,#D�\PH �N4
��)�Tp��B0�* �_a�,4�DE-4�F0Ď4��%�
L�:�CU-"�aGD���HL_2�H��%��Cl���"3�U,�-&ZI4�_Pm%��lk���
���?S%$�ؐȔ%@�L"��	&Ù��f�j$R\TD�$2W̤�!*�d��ArF�)��]����+*�h�R�J#D�!P�[B2�$&�aBI|bL�#��%Q�Ta�K�1��]N@CM�	%�Cҍ��2��D�a��3�Ԏ8̟�8AeF�-�&�OиC����"�_:dI	1�<� "NQDH�Bm�Ql�p6�aÔĊ���J�2\�P�؆,�(��)�Xi�P���v�7n6"$�H�0�(�
�d%�aeى�ڟ2'jD�#�˪ K"E1
��P6x�*��%��!-
R4h�OĂ~$;�>;	:˶ݶ��*B苸�.'I$㧯�>>��8�ׯ^�q��뾻뾯��]iGG_[Fݠ�J[��9Bs�/���aw�ZCl䀻�X��v�8��x��8�=z���۷}���Y�E�'�]��w�Ӭ�.^k��w��u�����$��I�8�����q�z���N;i۷n��MB�yT� B2Qܜr9p%�9��GA�8�	~n��")zY�Rԥ>l�-e�����~��.v�s��[{�7k(Zj���k�؆|����M�U�{�陠Q^ra�		X@���H$|�m���왧��FM�6�Z��2��wWױ/m.��x?�����������6�[r|���x�wi3H[[���ϛ��I���=����io�Qw/m�݁N�:�{�纯���duӜsm5�⼫��-m���Z]^���������uZ��w[A��]��|yl��[Cc��+�m��V�n^z�]�w�.>%��v����ۙgH��zyĠ���>��t�����xGZ�Z�_����qXݺ��ԯJ+mM��m�����YiE��=+p����;"��r�s���_��z�ߎ󽵝��ü��e��2N��dg����)�Y�a�(P���`�"m��d��1��&Z*�A ��4�5�!�D��Hh���Y'��(�S��n�a��,����6�|N��;mjD���Nl}���NE��j�i�� JH��5���A�B4Ԏ���E0�_L�ډ��f2Њ0��4X%�p�Th�$�ID.�5�*�$utCZ��j���0Rx=n��"3a�j��m,��v�	��p�o����v$��]�/��/�g}w���}&��R���e��߫0%f�'/�=�_uN�}�y��,38�;IEL��F���o�&�]Z4PC��x��u��ttC���S��<Kz����k\��~�\�!�v��m�o{WMg{��㇡�]��u�n��t!�ܺ�4q�_l�&N�6�	(j�F<�01�{漾bR�}��s/I�:���Q�l��e�ϳ�7��28�������/��r�3/m[A�9�7Fq�����:�ƙ;�'�>�s���>�Wʬ�v�?[}�.չ:\�`�m�C����<��1�1��1��s(e�zzob�V}������*��p#��z�F\�;�dloN����0g~I�e_���ʘ\��}�p��'���Cx��)��2���Y�Oo0�w����w�*b���g��δ6f&.�һ���4.`�Rmv,9J�6q�U����6W5#+>���~oW92K�oQ�xq��\c��+��Y��<���G��w Z�fu�Ô��o3��^;F�J�a�ϯ�w�����޺ɒu�ČL�h�v��fk�������c�@�i�=��l���tN4v�S�ʀ����%������4��?^�z�Z+F!c��}�W޺�ֹ�/Qݱ��ݲ�@<|~���x������i��g������O�ǩ�����׷�����}���fG�3������	�NyQU�Q�����۟q$G��h�~��Kk�٢pnp3�̎=�y'G��be�3j���2�����g�=�U��V#H2n`�[#�#�_/s������<9(�[�zw��A`���˶{�����W�5�>�+"��;�2�?I��x�Ϳ��Q���#zv����$7)(�o�RُQ���9��dn%���k|L�����A���͍gP��3�l���^
ݸbL���w6	:�x�l���gr�A��I�(v��&���.bf�� س*�2,�np��Z��R�;=wL�w�W+��թB�V�5��>�a�*�H
:`h2O������:!�\}}���I�o6��{��kz�m�)�Tov���J��N�u���͜�$!�3�����gna�և����~ݓ�إ���|>g����v{O1� ���l�v�3�<�6�۰�{��" ��D���¿1�%��cgl�֝y�q/ �ܡ=��c6C5���Es{l�q���$w [�y����uϾ������4�.p��vV!��R���}�e{������
�S��)���}͑��7V�0���;:2=����~a�|�4��Ӯ��Qׄ�I#2��J~���C�t�s'�t>���{ʄ ԮkQ�����E�t��Y��*]�Zd��ӆ?T�ud�z*�<��A��Q�t__��Hw�5�<g5zX�Lƾ��� �����dD��a��b8�Y$��c��A1�:(UwTM���h뇷�9s-a��#&j0�0���g�����z��/A��J/�י3��컺u�b�0�f��iWR�L=�9��$�H���^�݉Ѿ�+��[�\#�S.�
�;Q#���mh���߂�ɢ�C�1����t�u�������s�P�>�����_m���(�b�'ós��1��' ����o{�b�a���3�,�9�nq�,r��%E�'�JW���������s(wq��SP����;o��zM=3�mܕ/|��Wa�o�w��U8W)g~�=p�wcձ$�;����]��[r\�1�d�s�-Ǩ�n8�#�4`��@��f�� �p������VnȺlכ�ˇk~�Y�9�i��Ч�ç�`��}љ����|�3�o�[��5��\WӒ{�s=��v�"��� �s���ˎ�ȷ�Ľ��۽�}��gqI���ܡ�ݝ�_�͌�>��^��}�ڡ܏*�Zα�g7� �wn;h��Gt�S�y l�z�f���~�Ƴ��#�?����wW��$�{g{'/i�7�Dݼ�y9&ؽ�֐����� �q���d�{�g+z3�z����`��;mV[�T�Ϧ���j��<�$|������������B�`m�B�=�5�Su�Q<]q�4Ab��Tv���3P�wp� �v�F�p<��J���Wg��U6�� ����Z^��2�+�ɜ�W��������gQ��ˣ5�eWL�o��`��r�](R[�����U�"\pŔ��	~������p�
���}PL�u��d��u���cm�����|�՝���5�M�1�n�J�������P��~�n��XL�ݩ�cl�n_�lO>V
�y}�^#��$G���Dȉ���q�s�q׎�l��~>��=]�I�xe]���^pA�xL0k��[��7�%�7�8��zdɩ��p6�3��O�**%�rXV�m�m��ꆣ��N��#Y�g8�fh5��'�oI�9������ǘ�|��d�����K>pb��9�lX7F�M{�X﫾,Q;>i$�M�s����oVL�9��8'�^(��*�fA�q!�h����]�Nm����F��,X�s�n+���J_Y������匭ˬ�/�8�}8d�('�� �������~�֏���DC)}������p��x�]*�.A;a�*$�>��ܧ�����<bl�Oin��r�L�u��Y4Ԭ9�Јt��@@uƥc"��$[��%Uw_q��9�	�/g<\0�nh��"�w[�J��b7nbͪ%�7��o.ީo;� �����f
�7��PF�\�/�o��7��sǨ/ӑ�7!��K�d�2ѝ���_0fr�6�ȍ�p���o��wdǰ�Mt%{y*�s;��4����AuU?7��>�~�9S��w��۝_,��ʹp���TDp�H�Ծ�s�YR���� a�8���;ށ��ت�7���}�O7�Y'�sg�e�%� ����륗�}w�#�3\�Ț�>�w�w�p���������!��ݟ���w�h�����ȭ���3�2(m�ĐM���>{89_�7���{�t�Qv#~��i�����3Tz�l��왉��o_����g������V����[ƋL���=���|z� ��D�>��� mp=�l<{`���x�xo1�A��-��10�B��0�wM6�����?%P�%]}q˝>��֠�����ݝ�n�R3!<s�����g4&����$~&�C��D���,xz�U�ڱ�'h���YI���V7�G<�(1VU��S0�YZe����8Å�bq�K��M\��z����<<<|��Wu��Vn�	I���Q�k��>�����B��v���	�K5��s����b�{3~�v.ϰ ;�n��>���^o�u�g��C��t_W�urq�,�[�%�h�3�5��m���q&�ƀ9YQw>�ڭ�G�a�i۝�z�w'|�����<M�4�=$��u􆶬��.�^A��/9wY��`�Jw���î}2=W�4f�f���:o�s����N?<����z.4����N8b6�� x�/�Vw��U�ۥ�ͧ����qJ}�]q6�o*��B�_Ӯ�Ȗj������Ҏ����m�s���Jr�����>���_�2FP�C�w�1Yz���Ml�j�.���w��ʮ���58��f{��6�Po��*W��:���?���;�Z�5��Z����ÞN��X�X���=�}�I�Y\*�x�[Y�\
��q�u;:�ĳ:���l�|;m9����qW/n��q��]�y�v�_>>��TUEIU-��t因k����ٌ�*�Me�qDF�j�2q�p�2�M�;%��Ar�`ޅ���o�������9�?|"�m�k��Z���:qQ��΢�^�	/7sqov���B�?tWi=��X*��@��C`����u��Vq9���E����k��X�g�'ܚ�ި�1�}�I�	��Ս�]W]ݛ���>�~�"�����(OO��E���؛�{��g5����M�㷾Y�n�G�tu1A몐�;�U:6���u����5t������+:Mz{��}�o4`	P�>|��B)}� �~a��5���y���׋�6I�$9�]��e�x�� jo2.8�gy>;������mz3$�{}�i��~��W:jsA_g������S�t���`�T.׺��zz���l�ۘ����_�_w��V��>��e|y���bN?O��ϭ����`�(�9���] l5���m��{7�;�.�7�cv�WY1𩻚��꛼N|U?�'EP�����3k��N�T���毛2������d�%���Β��7�11��B�q��k�o{ݙ�C�<�;��Kw5�"�eX�n�=0CMJ�5�����UUw���P�f^���+�
bsH�+�7y��	�\''hW�ƕ�A����xuA`w�U_f����oP'�Nߺ'�4v�Ǜ��d9��Z	��m�Db��S��Z�{���N5c����״��]����Vv���i4���~.+r@�1Y=#c{�No����;}��&�og��ɽrw�����s��U���|�kz<��8���i���ͱy�~��I��n�ͨk=�6�ɖށD&��Z���h�W6
����*CȨ8:����{gc�X���oɔz��Fϸ/g����A�J�g:���C�m�{��wNH���sǳ~�s*��t6�EkU��D���=Z�{���{"�{�������a��(K�jj3>t0�;4%�q���o����^�P6;�#�x�5�u�_u|��rw��'J��Ibwe�wnK��;�Ή��%���l34���b�Ѓ�:�����{ڮ�K�MZ��v�LY��.U ����~������|�,�l<)��_^܄B��_8��j�b^Ūʗu��4�Rֵ��y��"�֦��{����F	t�D֥s2r9�"�0윖���>4�L�hY=�� ������vkh^{����1����ᯆ���� �va�o/`O���.{���T�ϳA����Q��Y��2|F���3�Ͼ����7A�g���L�n�_S]����`i������{���,��nd=���['	��$���dw^���`cv[d���tn�#��M��t��+{_z@/�	���>=���v�����b7�}�`<��v���1g���=.Na7ާ�;e�{`�l&���`��z��a�>�Ȗ���.e9��}�wiߛ���Ϗ���6I�ɉ8��������O����Cʩ����yw1�E���}�Zϟ�����hGI�_u�̡B.��_wԩ�QӸs�}�t���ܿ)x�i��=43۳�ע����{�{�2(���_�*<�I qv+�����YNN�����*�,�ˬ��w/C��:�����7�_x����t7�c ���K�tM�"�G����Kz��f��ilb�;�f�T�\��^^6LƟW�!���'+O�7|��R���~qy��YO�[
j��(d�e�n��
&��-�9�ҽ���f띉sN=�yJ'�8s�Jb+�JV�!oj��j��&㱜�iH<��+�ɹʖ'��a�T���$weN�)���ם_��?:�t��~�#��.��'���]_W&����8�B���[��d�<�0c�s��g�k���l���˓�T�!��A���P�wN�)�����WqN�O1���\�C���i��ړ���Y�B]p5N�Ƌ�5DNZN�u$��fÖ�N�u�ѝ���S����j��3t�y�ɼ�*e�g%!�؃]���> x;l��g�3� �$u6���4�#�n���TD��G�Ĥe�ؔB����lR�'7���[�.L(�0���ټF;����r1KÔK9�U�������v�u},���Զ���I�4v�������*����z Ӆ��f.��X�v���1������$@[��íIk�����uC9a1m�[+GM�dL90�'$DM"b��4��R,,�CN�:��cZ�X��ʥ�|��y��a�o�Ge���;����h�ݙoeƉB���aVF�"c��	&B��^t�ƻvd�Kh�hq�r񬗶�­f��c��7'v�M5�l�jqe���]��կe_l����e���H]����sK�L�LX՗�Y��.���S���js^�����n���>�j�y'75,���0mǚ�*��ϔ�=���Q�e���fV6��!�;�Bәy�+�0����dg\��;��]��8�J䒲*:-����3��v��.��٩� ����P�7α��l*3��Jn��<���"��z^�2��l(l4��Ηg�n���&�x��[!�t���9c����~4*͚�J3jiyK'r�).�M����"e�
�G�L�Y�1ڲ�sV�F���ˮ}/��O���x�X���.���6������*s����J�v�V�'�t%bS�p<@�6�̨����X��m���x�>N	-n��5e����ڶ�+��F�wrUdO\ڳ���E`���#�+(wB������\�ٝ������z	��-I+�oC$��D{'��u3�%�ٚ��!����uf*�t۬؟v��%���%(�״͡/~�>��{����>��X��-R�+�%�Y�x�8�����^z��%�s�G	ywך4䃰j}�]3_,�3`��12��H�M�*�n��@'��A���K����Q�j�{bB�$$��!��=q������q�����_^4���ݻ�	�*#'E�u��S�[Z���*!!	! �$$�q���ׯ���q�||||}}}i�o:6��ܩtT�����h�������8:;������{��]�߯���q�__^<m�f��Bt�YY�ٶ⣄�/�*����s�\�����hGIq�%y���n����).�m�DA}/��m�E	ܖy{j���H�:.����'��!�~k."$�����{VP\Ir[?�~2��J���ۇQ�J�V�w�N�����9���}3�_�u��(H�����ݿY���:ď�߻�ꐤ㻈�+��t�:���+����QIRG|�뎊�u�YYBtq�]u�:;��_����z�G���W,t�o94���R�&���/����\3���Z'm	}!9s� �Y����^�$Ox����CM/u�s�{^k=�W������ߙ_A3��\�5G�U�v�r\Z�M3>��h}1�khq-a��73�-��@ CxK/!pZa�.p(z^��X�����ݒ�� �����0�ȵ�t�E"\$���E�����5�D�`��G4��
<!�,���1��Z��*�C$����%M����͌YxsF>^.@~�{���h����r/a�c	�.�|�ف�p'ё��[�=`i"SY�Ϝ���0��wvkJ�O[ኚhw��`41��t3L�y��%%@w>���9�fƅ͔0E0ɋ��"���
!�=��!��$`�y�<���羧�/Ü LK�䌁LR�������^�� ��z��b�̈́�OŬ�3�m�d���"��gr��a�~p����"�c�/�|��tg������
l�֑��� Ǳ�Ǩu�h�u�z32���Y֐����z���弅�06��4i7�`sޯRhX�QRP�Ú����SqLe
��VZ�򀇼>a]ٚ����}������zO��₿�ŧ�ުO�R9�@�-,���!��v�Ix 7W�Я�1���{ϋ����P�GL��>����=��ʏ�{�ò�� �~_�A_��ᦶ����\S[5_S�#��ل"�VHH9*Rl$�=M+��a2\}[7�|��x�ϵ��>�w�]�>���lԝ_���"��@)�1 0�3[��	/&�K��X<�U��\z��S���2���������`y���`�PΊ){�L[�0�j�?��&'SI�Q���^�il���zS�}�-��$w�q��ub��ٚ�x��i��S�R��y�3/ P�/Z ��a8,ԉ��o���?_��1�s�{���ڭ�5S3���\���'�7\<k&�Ϟ�=#�/Ƥ������}�g~�6L���!Wq���f:d�}e�Bg���U�my��[�Z|�8�x�5�%���j���}
6%[I]�&o��3�ZB1���@��
��L�VHlx�B������wb����6�+�ن�K���Ju����XiW��2��1��*���v�=w]",n�.G]d�p�9�U�x�Q�x��O�:v\�_˷�tKz��̀������}��O��ű5�zZ3(/��-qC�4�G8G�椮P`(�!�"Ys�go&��EÁ#�'�{����ѷs��:	���w�m�+�õŞ�n�(���_l ��@�TWV��1��a \�C�p�h(�c)ߙ�R��VO��n.��ac� �m��$2��;`ǜգ^�J�aM@�[O���n��ߘVeI�$�Vn��G0���#׷qPý���0w��%�A���b_W��=��n�[�+���ߜCg����U^۸е��J���"��É�N�v�.Sx6��h��p���K9�kx,�0v��t��,�O�J����<+¨W�S�=��(��/�����;�=Ʃn�����N'�w1Y���|ؑ+I&�4?�����@O��8S�ư�	���z%��
�))�-h'$S=�2�&�+���}�ņE0C:F� Oy���G�<�C]��K�/X�nʤ����V�Jӏe���M%�j �����q8�y��0ס�!�Z4~���>���^]���U����@�b�_gKͼM����^ �a�Z���������WvV�A��AŴ��^�M�Zڌ�u�/{�ܹ��3�r�i0��<��,ܦ�k	Ac@.5;�y�����vag�2>���:9�qv';.J��oj����AU2�O�⨰�]<�mY����sizw�0��4�a�So��SI/�� =���S�
*��lّJ�:'��'�s�`�%�*�m� z�k	��0��S'45Z��sK����8�f��,Z��2����M;�P�/�Z���	���rUf��垽ށ�N��)_9ÿxq�+��ρ+}�Q;BWC�>9�	RZ��>��o/ӹ�
�����#���i@{q�q�nפ�@DK�V}צ%cБp@;��>jyY���	@��w��\�|7J쵧6�?G�[����ȨRub#|�`K��%�������Z����Q��h<��z~��;eX2gc������a��fs=�>�{n��;f�3yW^i�X��x
�Xr4橂N�W���9��d�x��4��D��� �$<<����9E6��0�㰙�F���:	��i�;��6`��3��	^	<�.�������.nv���p��c�u�zo&��A���m��K�W��/A+��{��o�#[�ɷ&.Z�:�B;u�����vt�2�g��?���Ĉ̝��ؗ A�T�h�E�x^� ��x����lK�&�]�Wr��J��m-s�tS�Ņ�N�B�C�Ͻ\�噢S]���7��������E4�ݓ�����#q��
i�S�;�l`�s��{=>�.��<'�K�rl�l��!
-�7���x�=�[Ù)@O��پ, Q^P�L��/uu�G�[빞پ�{k����F���C���I��~M�,S�ye�#�M�nc�ʈ����������j�l�9C)>���j��Ł�Ȃ�;����S"�<��?{:��i�Ξ��8�T[��]u�+���k[z�5��0Qb9�����T)Q������;K��.i�?7����0�Ʉ3�d�J����Hx(4{`0tŦ�5���X���34��k���Uz�YE%^�p5vk�e��&��8xQÛݝȣR���d�X�̚�d�Au�]x�L	,X�f�0VOյ*��W@zǠܻ�4|\=��V�4(g�o"Lɱ֑�WZovu�/fZ���jf򄚼�K6�����v�ߛ��g��NC�Ldc �1�*(H�"�	�o�<�9>|C�}�(w$k}����+c������1�G�8sj�0+�\��!���M#�4�����Ӹ̧j��Y���|��x��~�F�G�T�s��c����F�/�<��E1-՚ٱ/�Úw����q;��X���b�޽_(;��@���	KҜ�Y�=���fAM�.o��:�{t�͈���j�a�3S޸f+�W>�8�6o/g������	�S�Z�;��<�����g�wH�9��4��G/w�|&s�0S��	�L��{��y��B7��-I�h��O�Ȋ��9�p�}�c�[��o/ Z�!����v��~����^a2���3�ll8�����m��Ǣ�����4��)�<��=>q�˖#�ꔨ���}�b1�eC��}�������x�	��� on��n��R�X*����-/g������\zd(��&�|k�?n�1�ɸ�ň�D[�i[��Z�D�����Wu�̤������Ç�q��U��մ��C�m�>��+^�>��bX��-L�*T)?_��WC���S[��0'Ss�/ڭoc�˿ff��ܘ�ŀ����0�y�+:7��Ǽ��j�'sw�T���n�&�����TE�!��-q��on��μ��5���[B��C75�,�s/M5�B��i�Z}��T�����։'пcU)�4%B�cCP��� ���w�u�׿>!���g�a0�y�b��:����oВ�L���Mm~��c����y�M�`�.�{;��˗�-���ƘTX_�_��n��0V��3{�jԾ1�&(t	7I_0��>�ұ�eS��4�;߀�ԁ�@x,'n�ty���}9Q�=�+�>4~�B���9�=b��n�=?]���Gc��'���p�z��<�^�6i��G���Yx.�Ѩ"'�cZ���z�q�y���N:�_ch��5�=q-�'`�l�wX��ߧ��(0<�l	�����[�|׈�H&��/o��0��"�T�5/l)�z1Q`.�2��\d�(�R=>c�llV��D�O��-��d�|��v�DXv�5M�64� K3w׻t%��/�R���<k-p/Ƙ��u�a�Ú���}�9��m��Y[�����ޯ��C�K9�y��������ul�+zX�/��ON�>s^��`�{�|F�[߀�/�(�XvQc��0����d�$6<�f�+�$�qoC1j�΀�y�*�´W��wo�ϭL��"R�_x-i�����
Q�.���
�h�|ѡ�k�� {�x�[�w���ӈ�	@������h}�bw�<�hM9-mD�}3{.�>��1
$�[���Yњ_q9v]�`q��xG~ۭ�l-J�KÜ�V���GS���7�a���b��e�)�N�r��9�v����/��TV�cB��4"TRD��n������F�Mlc��wr��T$(�GRIp�7S� wP|���,��D����->���yX�
��ң���;�����R��_��}��g8�P�}X��^(�k��S���c:y/N�����#YD$��k�ti��%�@����@v�m�>�?,�q�uO���w� ҧ�ּ�Dv�ځ.�;�HKV�Wn5_>-��8C�ZB$�vt~�E��|�zk�-c�v�� �@�F�+�E�5x�{C�S��U��ƽ#;�3��{!��3�VS�t�ށ��� y������4?����x�wV�"Is�K����U��L�j> ��p[Ϗl�����] ,���9��[�9�}t���ޡ��<@ݓ%���o�{�Ԭs$�������M�+��Dׅ�z�Wj��^?�-W�_���2��9&�'��b�v\���Ix����'���M���iyG�
�f�~w�� ����s��b[]sl��C+F�^D�l��m@��'�w��*����0�^�t�$���Aq�`������я��|ݰ�RK�3l�n�v�卛Ex��%��K�uBL�����c����e6�����Q��8��Uc$����v`M�=V��[�v�,��JWfiJK>��^�s1q쬙K�1�TI	{���]������?t�)��V�����f�5䩃�"�GYΏ>к��+p"���ݲ��>�*�`��
�Q�,�b멬��w�o7>�_��ҥEZi�*1�4�VDdAd2�= �Ix�W��|C�T���&��c��㋎텮��U���£6|�kN�<�^�`e�m��@!��ġяJ�@_��T�:g���N:��ֽOL�zzR(�z��|e_)U���;�`�:`�Q��%`�	�~?�-m�O|�ϒ���{��X��V+�������c�8@�`z������G��1ᡴ���{ox�(i�2-�+k�xޚ�a�U8γ$i0�7��%0̰E6���c����`39[�l.`�q!��iTe$�y�̄�$�'}����E���{ sHF1�ߺxW�~�Ⱦ0s�.��C�J����bzp�^���ݓ��#nJ�vH��9O��q%�\GT	`+�T�k��Ǽr�ŽC���ۮ5J+�n5�w|���j��W��|<3�}���P�KS˄�d���	[��3>	�Zp�ʷ�T�R_ ^!�wW������Z�L�VQa [&�"O�o�R�i�T����Wf�u6�w/ j�u�r�,R�z�&�:��V@^PR��+��^��F<v�D|��g�	�w2W޽�ua��B�5�=�-Ͼ���<u!���o�������x�^̢9�KX��2j�wT�39k�(�pr85+�m+V(���O8�N�h	��;74��-w}�nCG��u�(��s1V���y�̻�5�e��4��4(1�4"�F!D$  ���
+�E7��q���$����=�tS �]�L�������@Q�k�m�6��k�tr^ �0�P�'f�kי`�%�fs4�t�L*x��7E2��C����mw�q��b�ߕ�pn\�fvA��r ��ǁm�/�J��P���C��[�I��S�,w؞T?{\]�Ӵ��|h��������48|�M7��m�ۺ����ɤ'g������a������5��ښm�a6=�W&����Kx��5��l���W�_��:g?O7���������,[e	��%�,�^�#i�t�/�_H��;?���a�-?t�8�`h�ZW+_c���Ԟ4�z���|���U?��}/�	��׮5��{'�y@�Ɍ�a1���V�
�8+�<�����^ �5��78�3RrS�T<��4; ��;EC�{�R8@I^�!mcFu�����/X3� �\H�R��K�Y��������K��2L�G��S�n�X�[�8�۽�؏/���|-�`A����'���'ߕqT��{��[�[�AI��@���:�������_���+��6=`Ʋ��\�D��1��Q��O��;����VYc��iB���ba�T[���^uilcP�Dj��;�_mR��hc[�m�}��,4#���zS�yL��~r�����c�?OX�(ƘЅ@P��� %A$A �D�{����x���g?;�}� Yz�x�=e� ��!4������~�~y�G��1%BOnq�B�]Vi>����{L�b�O���K�?�����
I�B˰��v���m�Lr������6j�x� ������MH���2e�	�ԏz����֫�E���Z$��.Xp��v�y[�v:P�lw�����}�}q�c��vĆ-���J@2$��������o��j�l�it֚��> �p�D덇-ᕷ�*Ϥ�A�Si{� ��%>ʂF�[\?�ge�$�+�n1ncT��y�����c�Y�;h��xG��W> V��X�]1I�|(����^�J�/7�4��~���:t�7O0sI�G��qK��c������C�ƀ�s��ꂼ���~eїZ�K.�f`�����rc>�i}���L7�p�������Ѩ@��	�ʔ0*���3��q�Q�k�zZ�9.s�,g����6�O����x��V�������ٚ1r��-�C���Vl�]<^n���U22��޶q�v_�6�������ɕ��^�_Xj��	���2�Q�*�����_L������]��gE��k�B,�Z��S޳�����X�^]Ր��|��\�P�4%ە�p*�뉸�>�8�n����C�I�4ѥ�%��&t�T�m^d������*Jx���k9��F.=�	qB�r��@�D�弇
����}N�i^3�rs�3����R�HpY��-��H��z�61�0�E�&����n�7�&�gb<2�uEp��]1l�7(�+�(�u�Z.����=���=�p�"P̀�����b0�i楢Ѿ��rK�#Dѷ$��y���o2;��BF;�Q��<�Kn�s}`?v�kS2v�L�-���8Pzq�TꃪZ���ݙ˧&�K����^Lf��!�ں鐻�K�p�!zq-�#��jU�,�]�8�cS
�n^Q�J�SQ���e�df)Q0m��"#��|���4HX&�(t���8��Ձh�n:2��Q�6v^�|�6̙�蘹��haGkb��Æ*G5!U��q�HY��]��;���������_<��xa�i��y�^Ǜ���.�[�hX��PLd&nXZ���,��͙�is)Ue�jiҠOMG���&��㝱�w���
�SY�����W��X����u��(E�(��K��/����9;�3e�@�~K;�U���U��Y���4�x��L��I!�P.�1Mˢ/�m�D��>���Ф��q��2\ۇr��K�}��}כ���s�5c�o��SXo1�J���2�V
��Ȓ�Ɩ�.��/J��� ��:����\��ܸ��p���֏���0&SV� Ę���De�8%�s���v;s;h@T[����F�2�.��G+�軏�q��}���|���d\x`W37D^c4Izp�%�����1���6�'�Z���ZS�*�	�����~�s�$<���DU9[�h�����#	V:�֫��z%���iwB�l��}�ь��f�r)ϗE[�+B*v1��`�;su�.�z �#aL�j����
�=��;.�.q9μV������Gbˍ�m�z9^�ٺ�syZ���}�6���i����Ì.���G'fe�'����6*e���x^�r������l�ˮ\i@wF�IØ�=͏9�3Kˏ���o�S9 s)d���1T�3�Z��kT��Q�z���>I��m����vVIԆ̑���k�q�a�*N{�k��6���"�5j���'t��B󒫘34Q��祮�D lܮ����%E;�����$M&"�צ�gv�� ��\�+n�w\^mUH�e�o*��'T��i@i$�d���9�����}�\�>G�sͱ;��s]F��U�S��^�� {�{�����U��t�q�mA�*:����i����׮�_������z��������o�"�Ȑ��j2H&�B:.�.�N$��������Ǭq�������������Ǎ��{��r%�Ui�G�^W�uo�ՑG�S�RH�=t������֟______^�>>8����o!q� �FIA;;��ˎ�+��~�ӣ��8ȸ�.�u�EAE�v]_q�Y�HEwWg?�������]N��_J�:�(�J�qqI�_w���g\y����8���,+���ӽ�v�vWfۣN�8�
�㨻��ugE�q�\uE���ԝ�\w_�:�u�\'GE�ڲ����uNtwq�Dq��#�����h*�tZ+]A��1Qi��QE$BO�-��-$����3�,��	�	e�Á(�x!����(���m���.�l���V��
�]]G!�7�U�G`�\RnE�ܪ���ʜ�T͝��4�
>0F��wI��%S�4�)`��	�(�B؍F�L�� ���$��B-����A�D)Fʒ����L���@J&�M�0
�T����PT>4ƀ4ƀ4ƑT��+ ������}��ߟ*0�8<�,;IIz��oROv��ƌK��/m�!F�$K{��k_���y�7���9;�fu��϶����v�j�{Y>C�]�Uȯ X������T:d�'���03w%e���S
����&��eO(U��O^û߀���e|�H=L��x�^ #>��4�mkC��_Y��/�+��:��Dcʎ̞Ģ"�7���w`-���`p)�� �1��/�ސ�D��kNtd<�;Zx'8 �_�q�q^o���[�x�"�Z�7"����0��K�Cń@�}���x>ջ {�
�[8[�<M�ǒ�/�ǖB� �=# ދZ����Q��/&�]��U$��9�s�s�D�Oي�[���ޤe�!
��x�^�@�����-���Ӭ�c����8��dSD�M��F��`̂��]ňx�>��K[c6>�9�7^���FW����Vlź�O�/e��^5�{.��Q�1Ml�By:��I�Zώ�o�3�ǽW�Π=���Fw-od�s!�g{��C`�|�m�kFZ��çz$=�^��T?y�C*�-���o}���i�J������qD��ܭ!�r��v]r��jԚ��������+�6��}�C���A�*�ڣ�e�3Da䧍���|��J;��>&G�I#Эq��N���y*���mpT�;�},+�!1�&˓���^����˿�P��iE)�����* H������u���=�g�3���?6�LP��|&���ٮ�^d�a�M�ㆼ9ק��8a������f���f^�����)��JN�b�X�^�Z���P�����T@mx�����F,�Ƀ�\�����5c�T�*�)���d���Z�B./��za�gw�[�������׸-�#����T��̋ץ�9�I��;'���q�e��,��@^�����nRh�����f��!�0ea�i���皤�_����	�,5���\�⠗����چtvZ����?����b��[?�3���9�6'�veu��iH��*$Fn�|hda�YC5�34��C��{{_3��L�� ������?�?��j�a��Ï3�ퟸ�"��?6;��f�;Q��W���v\�?�yh�c�)��k˼y����Tz�zZ���6��l����E�e�2Y�.ޙ� ~F f��^)Ẳ2����ɪ�Y��Q��.$E��.[�[G������z9���}���>��r�=�ݫ�b��@_O^;�mv�������"�v��qa�+)ݢ3E����{�d�އ���X���9�[��B��3Ɓ �H����^^:C/ʾm��H�J�~�P�-2ѴJNN�M��k���]�v,�RVV.ƕ�z��^������j�'�"�Zhii��Aj)����G�y�{KE%���r���K< s��\L]�^?`�щO��z�819R�hx���%5�[k��r�p�n�7���?^���Ņ�OJ!j�<������� �{�ű�^"9�A�W��2<�7o@�r*����/֭��R�aU�>@3�mw�1q���Ҍ�{�B�\�*���u����`'� �s`�LW��Q�ؖ��{^���=����=��L���T�eZfoy�S��gfggwB�t�SFG�j�I�7D�[��(x)�d�y2k��3��0^����š]�2n����"-�4Ö�2] �%�(�ahԀ���E2���Q��X-A��iu�i׮�j�����߼�cE;����@��cN@/���-�]��ā�g������~d��_���N�� KU�7�=���p����X�/���/�a��W�G��8k3ݡvv|����T*a/���T3K�e�k���^�g�@RO=�@��������_�LKb�L�d�ѓ'xJ�E�=}m�;�E>�f�/q�\�9/R�\xG�S��TFs�`���Bި�����b�չ?_�ViĿ,p�'�A��D�a��^p*)�ʚز4Vu�$)�ic]v^�@�v����q�V���wJ^�GU�ʁ"2�Y�r�M�˸���ݘ]3�x��Y����es钍l#�(u���p-��pwZE�Xʯ{��S@ SC@ SC@"k��|�uYꁨg��yc�ʡ��_[�Lzu���<x��Q� �J���1��j�FmtV!���P�&8�%�>H�ח_|�G*e�x���/�T<gX��A�ʘl�K�I�W}=7ǽ�~���� �׸,�?��Vz�?�e}����j݂^��x&]�����1k�!�v�o-��|��H�!�t5��鎼O�����>]�P�ݐ
���]���q7uEb;#[��Ȳ��y�7ϳ���H�?!a]g�z��??��ln��G_%���a���:��(��3f��+Y����.d8��^t_##����)�S��|u���{��<��0²|�Ω���&��%=��
�1�[ռ�n��AEy�dZ/�;�<Ff��+<1�j��+r̤60�i}�9����Q�ej�
����s�:~��Gy�0]8�I�6��w#_��]L&4����8k�~t�<�>A���&!��ƞ�:�}���-��g;��<�(���6ޡ����ƹJD��R*9�H�'x���|a1Zr֘�л.yo��).o��p��w�}UR�$����F�RT��t����
�6���[lQ�,�Y{O\�슪�.T7��Z�D�P;���ױ�WX�(ʵ�9�igѾ4�P�@�����*�]>"�\�J��b�}�e'��U����������{�{��(�44*��҂$BEAT$|�����<������u+/�����7ǟMދ%̬��ܪp�w�]mR&�"a�ݞ��ɶ����y���Q�!���*(6ȸ^��W	�8K4m��ȅ|ps(k�\b����|/��=:���su�����CˣP�bΛXÃn�7"ƏemK5P��\�Fc�J;��,g������>�m���{r�,�;��vf�b��ӭT�D�T&�}���I���=�1y�}
�FֻH>"wù����EM�zѾg�L�-��t�XW�4|��
�/�Opk�FP�Zj����<>oK'�'�<�����%�T���땸N�N��C�-@C��.�}@Y�S�)8��i�{�@:s��i�����o]+m�����T)�ҋ���?��	�m�:}��0���~���G�<x����?�n%��m�.�C�4�����ac�Fc�S>��&;��18�c�׎��.�w�y�=g1����޶�v���w���a*@��z�PnF��5���6�kd3>d-f����v�UG^zs!A텍��=q�B��<)A�{�%r�`6�����֑��IR�b�ѽ�AB?\e=54Nw.����f�,��̔
Z�w���ĖҽA�]�Co�"�WwL�9��\
/��IJB;p<�ޅ�J�.��.H�36��]k;s��ja�����^%�4�~��Xd쾽��W|�*�����J��hhE)���!�~w����ߘk�g��|���za^���^���N�M�Y�Az9X�uc>��qD=��^���۝]Ja�(���\��>i�uY��<���FD�B"3|ci綤�Z�����GOw���
+��������yKCC����u{f�;~���W5��T�)�ll�Ǧ��8z$=����؆R��ece��?f�|E��F�2X���9@��}H���N�o$f@��0S��06�QZ�ӫ\"���B����hε��/��2.��e���7OMs׃��?<��E��UV��}�\�<�m�Z�+�h��}}o�w�S	ۃ�,lܤ��Ig\fjxw�>���MWkӢk�U�Iva7�����	��N�(���H�3���@�9�����M�n�/^�ܵ0z���-{w��9��s���z�k,0%�N	=+��C�0i�u�[*5q�����xI�S�����`���OF-ߕ�/��D��_}�Z��5�?.�G��K�3������@����][xV)�Ւu�	-&�ӱ�P�|.�|�W��� ֬xNL�0p>xg�۵�!A�
����n��]v,�;�8E�k� ���v���!Q���(M�*We�p\$��I�"�Ei��*1��U����uD������EMUL�VXff�;X���=v���&=�P/t�`3��A��)0�\L��v�B�e��j�\�� �^�+�%?v8�\tD��tg/���	�$��00J�5i����R������o�����M�Pݟ�%�O��-��^�_o$��f�b<�2�
<%�q�pR��j�Vk�s��S�Xͯ������}��|/��w�t��|��hp���: xo��L�c��YUa��B�ܮ� �EH��JE���cU��A�����9����;5w�-@���b�|��Ɇh������+�B�Ōzbd0uO��[%b��\ٌ��m���S�f�K�Z�]!1XdJ~���(����߱��i�򃃠8`��c�ڿv^�OfT�����y��R�CTcH}"y��ŗy),P
R�w7�@k�:y��x�-���s�����u�=���L��|�!R/<���ϣz� �5�>��%�n��䕦^�כDfL'*Cr�]J�5�����'�����=!M�/=�Ez��%uEӷg��r�Ҹ�!<�|ǲ�򯻯m^��dn���5�K�U���M}ڨN�����f�u�3�4�7�"���RU.Nw�c.�!$�$����4��ʼC3taum�U%VRWbR�����'�}S�V��u⮗��lE�b��ھ
����ɝ\��W�����E)��U}�d��3�r�}`>w�ޘ���^[jnBm΁ܨpl���^����6���Ed�s�E�5kQ��tɄ5�v�}��t0txc���L��r;#�{�-������Ty����	���c��v���3ٔ;���ƙ�I1�a?<?�u{>��]�1-�N��zXem:e��Z�zCiQa�B��T�/a\5R3^�n���� �]]i���g��̷1һ�c�;3w{<f��{�hm�S��ӯA(�z�O=v�p͚�6	ٝ��Ĝ�cPv��B��|���L��R���W7S�҆��^�-��gf���NO^;_��p�
Ǩ��&����A>��fϽ.}�0�Xͯ�]�����4��i6�W��?~u�ݙ�?���^ĝ,�3\4�(�?Y�a������S����mO�v���=W!fT���a�00oF���Y~^y� �
c���<5��ߗo�7���w�ض"�#�39���<�k%�P��=�s~U8�5x���l�zǶu="��0��,:/�Itc4��w�DR舘⹚���sw�|���J^����b�P�m�w�$gV�NV^��VڛG-�\�;|�};��VGZVdY��ǵ9��	[-s*1TN{dc�Eb��Qۺ�6Yz�V�O�eH_s�*>��O��� )��i����5y7����^%��^��6\ȑ����:��w-���i�� ���6��s�a��؍�`���.�OCuyW0E��i�?vf�Nm[�MMJ9��m����D!i�1 �8���4���(�"C�Fi��T)?P�ƛ��s5i�ԛ�����?y�K�^I��<'X]d��U� ��x.���C�8rӗ;,����/��ص�!>�^k���z���Tj�dH��ʟX,��q'��$���f���1�����V���^ 3�Nѣ`N���sW��.��{ضQ�!�m���.o���F�S=E��~�j��Ǘ2]	�>'����������Xw8}���P��T��z���[�'�< �fpG��n��YVgP��'�(Y��C�Q���X�$�VQ{�g�9�߬�����q�����'�Y�V_o�؄3�2��kc5I���RP����^��E&�Ƀ C����0��}l�fE.x���5���zx��J��p�2:�J�a纖K�z׬L6WC����-� C�"�AD'vT��v�'`�|��S�k��4c�ڃ5�stqv$�Ǟ{��KT� �>�-��Sۭϋ-jnfM�s~k�o�,�t�)���W�Y��>�����&{83h�iiK��k�(iYe�ݱ��C�*Q�=�Ej�EBs�^��L#˗���������	�����jhi��������X%'z�c2�6��kt�N�)�=(��0�M���ч�t�$>C�ޑW5{O��G��d	�נL;��=�"��^��S"\�%ѣ!��:�zjyC��\v.����gPُ��Wu�#�8�� ��F\ή���>�d��(���7�rcmuJ��pE�y�b^�7����PS�����PJ�)yHn͛k�hΞ��al��g���ܤ�'���7нA@A��j�iE�l{j�u���.���|�n#�ֳ�W�!\�x{�˅�h������琁��<��U}�\xmn.�����:r�d&��>z���P��צՑF�������++�t�^}����-����v��&,K��*F����%?X(AW�IN.�gn=4*��o@�<�'�r��o#�������PlO�����c��o���R&�s�=�"3M�C4c<�l���j��Eu�F�\ք@A<��"�b��f����:.���@- -/#h�����G��{��f���i���l4��q��5�u�	�$��n�Z3�%�CuX�jUd����,���A�:>(>J��6�]����S�dF)�L6�`�	��$!?h׆�fܝa{:��71Z{�M�9�Y����pq��Z%��d��3Bd�Km�֪s\v�d4��9��u�>���F±f̀S����Z��x9o
����{�S�����p=�	؜2�ԬV��t��jJxv��c��5"+���Y�N6�ݩt���˽��N<���!Y��+����0�H8[J�����8._]��I�V���1��&��F�fN!Z���4�l� ��������iA�+/�v�H��`�N���"�5u^��Z�\����f]��SC�|2���=���63�w^@��%B�7�/fl��[J�م
sp_`vkh��6/�t¤�	&�cyх쐠�=���x�a3�2��"k1o!O8]3�z���L6n��3�� ��{7*��$N뺍`����p�j��r�M���X�*e��M��h��(ճF듋����}��Ǳ�cK�u�N:y��̴2�֠v5��h��!uDk��e��,qm^(�媵�9a��fcR�V�D��"��O��a�Kݍ�+Ԑ��;��YWL3�r��2m�R+��[Ul�����n�9�ǅ�H���JQWG9�UH�Q�^:~~-�.;H��]ق�6t����8ӝ�;U	�����T˭�~Bv�"{r�/O\S��c�c��������Av�nLy9��W蛓Y��[ut�g#w�60!��Ü�dq1!U�w���oڮ����#��EdݡD����ts�^*���\�N��Kk6�}�(��t�v��L���w�6�	���.�����řsp�)���6��$�]J�����af��Wf���޽�x*%��Q]��c�>���J�mu��G�Y�Cw�dZ�h�J�����\:U���:���gt<7��i�v2*�t�U:��Wբ�/�LV����;��!a�*;S_�%w�S��I:^7FL!I�(���B�MrF�&*��8��T f2('Io��G��鵢�1�V+֚=_J�}��_�9I�ׄde
��)�~#�Rͪʵd��G��f-�N�x���Y�9d
�)�{�Iw[�M�L�>����Vu8��k�J�d��Pͽ�OnH�ۛ��fe�}��JN�hOh<�������e��6d�lqݙ7�����;��k�ǀ�yPb�*늻�V=$'y��.�^��i	V�s�Ge� j�/n7GZۻ�ׄ_J����@�W6�s�r����g����ۆS��2ֹ�����[�:yG���b�~r�|�O�L�EBH��2�C�'�!''\^_�u�z����'^������֟______\q����׏:t��"4D� �5.��U�y�yw�vQ��\Gp������^�|zӎ8����=z����ǎ���P�-F�AQ*��吗C#p<��#dL��)"�B�P$d
z������ǭ8�8��=z����ǎ��BHʠ�4��(m[k"�������(�����k��|���^Vm�ʎ(��k��Y\Vu%P1�;�Z���5j/�RگN+��.���묫ߛ�⼮�V^wVq�e��Q�qv]���9�#������≵_��������'�6����u���YvWe�wm�8�,�:�ݝST�d�
TBdC�Q�A����Ph��@����8�N�����ѫ!���4�g)l,����[��d7�&��~���N�P}�}��e�9�������U1�)�����<=�b�ԓ1Q�1����1����fv{��i��پyj[�)=��ʡ�W7�5��zRڴd.��u5�k��퐼q!�x���	�7x��ViM�,*�O2�������}-+�`�����]R���ɥ�x;��%~:}*sͭ0ȥ^1'�Tm�77)��u��b�R�[�G���;�0��g`�Zġ�Hɥ�s~��9�����T�_i�I��ve�-�6���/�Z��<'I>�Y��c����N����-��Qv��9��_>k)㬰
}^�f)홮�٤»�(��kס�,h�l��ױN�G���f��y�*�"Wh�����` �/B;�I�����=y��a�l��>�c���I�c�馡d��)�; �u�!�N+���38��2�N�i�[�����VhZ���u3_^>��K�C���h�9i����nE�tn8��QN[����P���?�!>wr����W��H��f�S	�Ѱu�*���ӡ��t9(8��6q����s�,��m�#��>4&�r�Y�Y!�FFӊ��h��v��*Zd�\bq�ǌ�\�h㰋�ƥ��.Y(4�_]=ĝoM�0�ak�����u4q&Z��,�|]U{�T��{���x%��wQ���GX��U�·v^�#�d�� ��i�3ong��:���_VK�� {�z�
hiB��hh_��>����w�ߘdO5�29�,4)=���K�>�z�����v�cH.%�W���71p�.ըg��z��/�I=wE'%�b==�a�*�eyQ��U�Z�X�WG=�j�imS_x3��x��c��_��2���S��L�$�0���n�OxҺ�p�&�]�΢�@�	�3���=![�����3��KS��;�R�ׯu���i�,7qo���7_���mO䨿�5�t/�ǎO�`��O42��a��wk1�0PS!��t��~d	��9����t��,n0�|�X>$2x`k�i�y�#�Y~&�)���`�3Se�D�qDc��t3�YE%C��O�G5uZLf1Ϝ�F�h�v} �����+ȏ3�n���k�2%��������%�PK�TeR�g��2�-�k�^:x�.n.��-�s�v�K�6?3�1���چʡ�<j}�>�r_�|z��9�3�&�Wt��ĭ�v{�fHt�$�z�^<ʄG��`�|�'��Ƨ�,o_�PwOJ�P��RU]A�$fGJ���w>x-*�Z5يlҐ�?�V����M�@#m�|�w��%�✆�!������J��ژ�JÃ��wh��Z�k��펎��w%J3�=���H���t^Y�|��k󙜯;r��ߡ�hi@���P�,Ky�I�4Pٌő1����;xC�.��cT��LT+o�`�*�{���a�����zG@���ï;�e񒬐��l�n�/ڟ��E+���y���g���E�pR�q�k��
�A:/~���O��_�Ү���.fdշ��'Զnwt>����U �1�����}T5KLϸ�V�k���'�����\9��h��i��ݤz��s�@�]B��W�%^p��]A�o�Y�z�Τl�w�Xqm�Md���狈m9�sV�/�5�"�:p�a3�`v�0��W�)6�1Y����a@�ff��{Ǭx/�xܻge��4Z�drfHL��%�Ϣ�c���#�;��v�1/e�V�P�6��tiz6���ͧ�n=���=����{�`G�z$��������b��s)�$���nqz�o��R��ݪS7���ٹ��L�p싇5��`[H�L��P�C#��w ���:�C#r3sS�c�6Q��>Bd���$�J�;s�__c��Q�0�mzc��K�L��	��%��HU:��}}�9/I�R9�iyG��Ot�l�>5c����e<bMN��/"NI��M;���������Rx��a[狞ˍ<N�UI�5��r׭׷�o�.#���)��c:�X�f��e_p�:�)٧�Ϛ\��.V�ϻ[u���讦/C�+�|�V����z���@��44+ �w�7��w5^���p�xeOS^�W�hU��W �flk��{��}M#��G>BE���e��T�90z�vL�L��4&�ȍ��ޔ�U��/7JG�T�̗�mz�"�VFpl(Ot<3?y]�E�3�~k�J��o�??yr+<��v��#+S��W�����{0���g��T5]aSI�N}ϖ�������AX+�N��wU�u�^d�y�@�%c=�«]c�q��:�ui�U��Up=(������vz@K�e����R�O��F�A�׻VP���4��`�vM �s��E��9�O��Ѓ<��MOi���v��giÍ2���+%�>3�Ց�aFF���I@@���Fupߕ�c]q>и8���l�^����u,�sD�'�[�FN1O��yh�	8�{0�A�����d9�T4f�ȴGMoqϮ�zw� ��@��f=�|p��m��&���7��)���:[h�
�9wj��ƾۋ��{[ ���.u>i���F���{id�~1�dX���IY�W�/��a�ǚ�O�4�1�����ǧ���mm���'�}ұ粆tab��!��S�V��%������-���Lf��]��0��ǭ�\XB�$J6�p��^e��_����<��N�C@SCJSCIM�� -��ҩ,�p���%t(ߥP�5�Ʈ�Tܽ[� �9oR�"�a'�-��� ;2Eֺ\�Ps�K�"i�FB�qqO�l܋�<���	l�-��j�}I�Z�j�X|]�kǏ5��J�m�Y!�%:]��|��A��ᄌ�V��x�ɅVS^�.����1 �����GG��ڎNI�d�`n��.���vk����yKiaz�Emt��m��t������u3����m&U�(��X�r���i;�=�䬭��k�sZ�`�<;�N���p�ɶ�XL��k{�+�%�(NIN.�*,6�B��O7�&�ɇ~D�L�n���\PO��Y�V��(x,;a~;Bo�k*ỗ>�b�;ϑ.��3�j�������euE�Nf�/���0��s�����@&о%�zc���������ze�Ɍ��q�3*�=�E�,��ź'���	�� ��^�9�ՠ�xU���1������v�R�S�3^�E�wD����G=�%�P-��<6u�K�mP�^qy&����A�BX�"Ы��Ս5���R��ÛS�P6�1�*�wD7aw�����A,Y�<"OF�E�x��Ӡ)�\C�f�T:�T�KJ�2I��>����6�~�>�v���|�{��dם�ް�q� SC@��О�f���Yx�f���[��C��������G�Y����yrA/HפĘ
���5v�J����r�4��CX%}�s��|���1��ϑ���e��/W�̲F\�oI�w5(����'jjԉ,�ѕp/�����>W���Sg̔�
�(|+����9�=A���g�&VgX��̉��2z�c�{�Ц]��u��$���6q����������aBi�]�Y랎��8m���֣���(Ik����\dx�w�G'<����z���{gh�-���\&h%fE.��9�z %;�� �_[P��z$��%~��0==�oe�Wڬ�Z%aB�i�#R�}��|ú�j@��ה ���yr�.�	�t�B.t�)�.�eA%I�s,����u�~�g��:�˘/@�x
ȈL1�/ѡ�*��������3��?�V��ĝ�WZ��
[��
����]$���%E�y�z��ǎK�!��\e�R���x�=�>�r��Zr�������ִ��9�k4��������#DV�3�S�N��I�%�ES�*����R_5�n�ɺtH��;��5��I}���
ζ��&}W�}���0�D�`;f֓�O�?����\+�q|ʏB�4 �s��Tk���O�`|�f/Ed��u+�m�]��9�]��2��y��q�j
F�������9��c>[��9��5�sk7wr���s��V�6ɔl�X�q�t�%�XCFE}�ʌ<Zq�y*��9�=$��3�Ly����=�1��ެ�ry_��h�T�;־p��}�̮�C�����ڸT�צ��f�ф��7=˰��m���-F���h�O�����綕����I�F>�c��@�H��\�T�N��\ʹiHgjB�39�9���s�V��qO�Ι��/�8.�-��X���͑b�t,&�	���3?�i�68�ZH�ޡ����s�Sgޞ�Ec�Y�����o��*h�J��m�.���:|����/���6"������#�kJ=>��Uj�r����;�>��ڍ���8Ԃ(i�w/b���xlhg�L�{����.<);,�dFJ�[�&��{`ֹS���zh>��{��� Բ-�m(�o�/�3k��|�<*E����xpg�[V�i����ҽRF	N!M����������ϩ	Mv� �,�OIt��v�p:�u6̛֨���d�*��u���6"X[��sn=��o�|85��O�=��zݭ�܂p�p*�������(�!� ��iT��]t�[p�9f���c�N�p�%�C�]N�dJ;�i�w��>2������^��
�4U�6�f��6��ṇ����b���7��s8�h"b{,��s��ɽfn�ܟKO���CCM �=�2�+�����z�?�|j�t�)�(�O`�<�P���:�4R�����w�[!@�=Pdf�ΞѴ���PFE��Mmb;$Od\:���0-���O��2����
;�����XEb�i��N��h���\8IU���~n�F��Ú��/N���Ƕ-�0t��G�Љn6�1(�[<�xנ�{SP}�]Q�i����1i������zi�����Ŗ�7jں|eM��'�ۺ�}�^�q>��X����ĘP���x�2���w:lw^�!ٙ.��/Xj�)r�dG�Ld.�O�^;ڐL?U1G#�6����'�]<^lR�W�3u�r����1��ӡK�� k�gA����>�uP� ��^�g�ejx}ŕ��l>җ�M1����^��8��ߣ�/X`���_�?(����D|�/�s�;P�۸~r�D�3լMR�q��%�%�lç�}�A �2�ҍ0�j߫L;h�8�8yơM|�C'ܾ����*֏L�h��SV+x�K��v����5�6�a��D�o�!�89� ���Ve�|v�~3��A��f�Y�����Sc���ܯ�Q���`��j8m���)1	K~tR��v�@ɻg�찯����QA�.����6�c*_sjT�������������� *(y���w�Vsߚ.�Tk�ź|�1��Z���z�}f��t�t� ��˱ljO��x<5��g3�ү�noq� �L����x��eE4WA.(^��J�H�m��t��$�J�����/�������I;�����j�S
�\�ڏ�5�ݰ�u���/"�U��U�ф�ڜmk=�Gc����5����,9� i��ό���|ܔz�`��'(ľvo4�w���uLNM�4�ĵ[�33-u�1��iP�
Kg��}���Ci�R���~���.�~�W��͞��Uܨ���V=�1<(xk��>\}=�}%Հ��P����7"�t���	�ʭy�J��^�������!�����_@݃)��� �V�Rz"hW���ٮ�8���=F��M�7(�xxc���=��A�l��M��_��`Sx` 2�P�~���v<�ɼ%����]e�j��W;�b��B z�J���X�W�t��6��»�y���NogSKTY���Etߴb�M�dN��yƸ�C�9��)���7m�W½ش����wE�)��t,�hi�f�fjb����)�]4��K���y���.m����� ��=T�����Q����(J�²�k�,^�vʸٳ�'T���[39m�l;�ƄToV�0�m˝Ӎ�Z̳�~!M-44	P�N�lT�k�a���lu�[k`秿E��@`��C�W�XS�	����D2gn8�����&_�U�k�Rq@���eA/m~��@;�0֫;5����Q����y\y��t�|��ۻ3qB����*Ga�]�&P�hi���Ǧ�U�����Y�1�	h��lr��"a�ʷ���36g����tb�ñ��ᾓ�i�C��j��9�횲Ж}t)��a�й��VE5�>�#��ѷC��`���qǳR�Av�V���8���g+���K�x;���{��ݽ5[�@���p�!p�܏Q�v�����gP�ЮG����]7tůLW��0A�8�w�	)��t�<7��!6��/$z_�U]k����>��j��>�T�����͌a�&*��:)�Ψ� �-��͇�ͪ��ύLMǳ�jG�&V��O�A=�Bޭ�^��3�R��q���uV�������Z�M
W���C�����C�%:J��R�v#f���!�M{�)ES���bP�>YV��J1u�t��n�nZqV���p
{#����PU�ݱ�:��]O;_��*F�(VhV9V������i�i�s�\w�W\��"����ifW��
5�j��<�{$|!�K���Q�.�Z�HȂok�x&U�~7�F�Q6�X`�:7�!��GM ��&�����eYqQ$=����ݨD�e���b�%�lV�z��;-<�0_I����9[��筌��A���(֭[vP�j�H7��H=v�L={f����l*Ɋ^��O��wJ57*zvdOCT��LO��آ���v���Ӓtٱ<�[�d�b�u�l�9[�K����peD���f���*9���o��z�tH��-��n�Z��H��BqV����m5���8�G;&a���4��ָs�����+X��Û�v�Vqi����A��kY�\�Zk�%�������@�;\E��rZ) ��Y�m��׳K�Ӭ5�>�x�<H���8:�X�W3����w���A��82;[�Z�:]�B5��x7���� ���~Y��x�!.�:e�23oWg�7h�h�ժ;Mc�(Ќ�1L��>R��'��vrO�iŚ����}Z�+�
z��̍e�B��Jhr��oPr���az�NDr�TE���h%j��l��\��t� HIƍ*�Xɜ!:�h^��6�;�Zp*2��GI�j���$�GںXþ���w�t[{�,b}��֙:�m��k�9�#PUۗyv�^��!:���Ru�Șho:X��t�#��(����J�Z�񽄭�9�;��/DMomYd!8Q�Oh���^5�I:Uφ�}S3�[��	<����ۺx��*�VK�=<;��*ܻ���ݦ��%��ikf�����h����yo^�T]�>:5��^6e���jޗ���k�Z�Oo�X�gd2b�Y�Ўv�"���6Sr�7e���E�v��&��x��#=N��9ks��&m�ưL���;m�J�Wc�����-
7a:���a�q��ME���~��؉[���x	aD��s���T�y�c���b-'�f�
�����K��b�������.u"��ڦc��ϩ��F�+̺�=`ڹ;M/S�_0���]��x/+'a�@�v�6�N�@�N��s�kP��Y�7��w���u�����WI�o9k��R��]1�|�s��wg���z:�	��mM�="�NUܨ���vW9�|
��5�t�0]D�U\G�q�l򝥼��uaT�2]m[ոpv'b�vK��A�G�������9ڄ�$f_S���LNX�^N�\�V(7]�#5j�*�+x� �D|�q��utuiDe��η�޸����q�q��=t�������5I� �Ad	E:}}}}t��델�8���������в� Tj�N�tBH2z��j����! �J	T�m����Oq�q������_^<xމ���u�Y�j:+3�:�+l���yY�wI���QV3q�ge����(����m�c�wiyg:_>�q�P��'ar]�vTv�Ie��\u�we�ݖ~;;�J+��mfqYvf}kE�C6tM��U�_�|Y}����4�Ӣ켯K�����t����:Nz�wY�n�dՔ�n�;3:8��.:���������r�:mgVw[��>��Bx�4|
����SM$�4b!Q&�!���/�nG"	�C,O�M¢!�TQ��P�pI/Y��w{P��yM-��\(���e�ɖ�p�wE�c�z�N]N�%�i��(�hkEI�}V;_NאZ�KD(��Fʐa�"���W�⾁��h�X-F�i)�2J���B�(�T�B�FfC"e&+�HiȾE�M��D�E�S������&}����p���K��I	�_�HSCHSCH����y�_���3q����CgS��f����bX�i =����k�?�Cx�{���cEl���2����,����\��<<^�b�{o8����w�����-�-��]z!0Ɵ�F�T�B�.	y���<��7�4�e�N�<f�ַ�W��1���6��6�;���B#���m��}����{h8�F;�_ �J��$���'������PN%��ٙ��'���ɵ�F�֐N������	��>�3��rP���w�V�Ta�֣YE�w:�������>Q�ìl�2t�@�5�I��W���|��+ ��1�\ùB��},^��+�j`f�0�V# ^�YbMv�D8o/`F�0	�;3U>WE2��Cy�S�L�u�~l�6�oS�xӽ7+z�zᚼ����]�[�2{�վ˔_lsǥ���&Nlc��a��Y��ح�igw�]x8��G�4J=69a��%�1���zl�	zd�$6.�|N�Q������s�^�#��};�����b,j���g+�x0�E�7�k��]�F\��,���p�+��/*��+�9�J�U���=+�Ke[�m^��R�r�mְ�S�p�",4M ��4%~x����6�5{3���q�z�#p��W�W���۽�b���[�1v�֛�e�O$|�V�y�}>�CT�����}��������ھ�=���s`���n��I��|� �*�NN��"T+�:�ƺ�(ى�靤xr�!�ӛ�#ѯM-��nC$�����3f��=�����ݷj{dt�(��vI�<�C���h��^b��*-�%y>qn�ـ��0d�� Jt�b󋼨	�j�?a�|{(�:��V�U�|<�`���~�{�z[�`.=��g�E��"ǩ�C�ݷ��ܙ���\5��~~u��ύP�i��aX�E����*�dŻTPPaݐ޺~Y��iKqu�����.���ݎ'�.�k,@ز��-�}�]�o���eC2��:;�i�;�s]
�nʔ������&=a+-��@��z|�<�a(��X���d��m��.��!�b�o����`��eDŧ�e#�s��i��r�V�i��9�s+�c1.9C���A8���OD���U��\�fe�z7]���1;2�9�Rj$c��}^��}���)�O�_�����j��F}"$յ�����B*+(�ӱ�S�N�ȥ	NI�ӵ��U��O!n���c���,������[����I)�֥CW!U��י�&�T���hjFZ#X���fЛ��D���<^\����,
���)*<���q��6�M��Sg+����'�y��Ǜ�<����A�E'̧�e���1���"
����f����U	}l�W=zy�s#Y�^Ӗ+w������r/����|ޗ�-y����ACB��~:c��L�.G�[�+|ǆ���5��;+\�i�{�@;\b�3_3z�q���ƵB�<� lW�$�|�Sݬr�P����;-P��UoZ=;���87�Xh��A��ۙ�鯺����m>�uV��%����1�)���Ռ�O�2��P��\��┻J~kױFT?pN#ء�W/�AP%h�}a�՞�:_8��?+�b�Hnb�!�Q�.eH�V1���@ �g%����ϓꨩ'|$z8��\�M�k�7�z@�[��M�����md�v�4�lmj�h.��Q�g鎷
5�ϠE�y�p'�-��>��Yg��<���}�VJ�����m��?z�A����5hХbU�{''�z�<9�!�S�<y-�ރ#z*��#�^��=��~���0���Ơ��;s�	�] �B��]��0�zhXN~�G���s���gm���T:p�����^u.�f)~�~d|���n��΅�v�缥�c��yތT�]7O���J(�Cm�VX�s�[�a�Z����X;�.Hܧ+�������3l��l��	s1��4��S��Ȯ�������?��q�8��c�
��ɾ�{��rO�5�4���*��d���)=$���c�GY�g�OG�\�=>Q/,9 ��D:m�r�Gr��e/*L�����A/L���09�OV�k��9��я{�ﱡ^�X� q0�Ѕ�����"㷬s�K�/��X7�y��63ΒC��;�iw<yg��v23ɤ�5�>Hg��9�"�^����Ǟ����uWyMG�b�*��Z�q����GＰ��ĻU��c�
�B$-aN&5���;�A�C^!��
k[�)W�$����{EW�Ъ9���,��u�͍�����78�(���:l�8$����B<K�;2��Joi��W0/�X�\Fo��� ���Z|����;OOm՚T՞������!Z��N�O�y~�"�Pk����G���s&���^y��F�3~�C��,�ZZ^C����H�.�;<���tT�$w<mm'�7RU<T��#/Yن8���c�k��q�E�O^��zj+F��X</��ϴ3R�}t!Ё�Y����ndGtHB!a��X��z��c<L��Cm����g��:�ȪRa����C>��VI���8%�e��D�0�琪u�Y"���-�y�=�{��b�`���waOGggp<#���g���a��}X�ΕUT�$느�妠��������'U����ɩbQz�g�{��������|��Cc���
b���	{�0��uP�s���70챖�{�>�3��j�C#� ���-�� �5�g����6��2�̲ۋE�+�5BAy׶@���Ik��*�^6-<#�8׌�=�C[�1���ތ8����)d�| ��!��?��:&��y��),(JE!�Ͷ^y)���^5�4�x��G�5�2�|����1�Z(L�1}��[ώ�zj5���i�5C8t�Nc*v�ʆ���w�q�w0_XX�X��	3�iƨ����> z��ޣB�s�l:��5ʩ�3��~��ú`�A�%� s�"���Y;�C�C�P���M�1����5�F���wzX��2W8�_�z����PXǫ˨��W�������d���4��t.�_d�]�S/C�uS��=v�B��a��k(��砲4��a�ǀٻ�׫�T��0󛎻x5Z���0d��p�jA�̚W�w��[嚪.��c�R�}����ƶ�Hh
�I�:�r-��	A;I�IjT�r�qA��bܵC��v�]��7q�y��ְ�������#��H�k�n�u�qa��5�j�UqW_�i�S��ˉ[�=gX2�]3rm��:�S���uY�Ϋ�<�a��;���|'0�4+�1�}�a����<�Z���"���^�O�L�yԒ �L�����{�ݗ�9tǅ�`���8<��^�]�i�[��ϊ<�纲ै.��ؠ�3	�Y��{����}��E75{��&u��<C�4:N1��}��"p��_Z��]ۻL�VA�N�`��_x�Ā��m���:o���eѢ��x>��e��xi]��%X�]K�z�>{���_fN�>�o��͚����V�I�Uܫ1�T�7�&�寷:G�O�Dd�����y���Q��+���W��`��(��ٴ�-;sm!�]�O�Z���!6�o�j�=$����ڭ��O��j�Ϩ�Mg�LVD�7�9jj�ɽ����V����C�ռs�3X �����΂
:�S��_ �C{+4'j!fK��j}�SiuEM6�T�U'��kU��2�|j}C�1�����G��4J㞣-l.,��t�(�N��/`�zh�ĤS*\i5��;$OdvL+<��p-�BR23�m�U�]��ǽ�FgCV��T�L&��rP=m���5��c3���w��C2�!
��3j|IJ�3�d�g
�vc�81��tKG�M=�$���q��g�Ø�"�*N����y)�������V�A��]&9k����o��y���=`�>㦃b��S�8�Ƚ�$�]1I�EJ�bU��=w�O�ׄw��z�L 5��mgWp���#��L��B�_���r��1�a蘴��R9�9H���VSۡx)�2���Y��=H9A��G�?4'C�H����Ly�n%��
�fW<W�ςe��>����u6�kGVg;=�j]��ׇ�~��Ƈ�p��Xw� ��_F!��k��zUy@�%l6e��Q���p|�y�*�ҹ��s�]A��ă�~���΍�[Ծ�M��� oZ�Fm�#7[Q�V��/ �2װ���z�O4��zt���3΁���O^�+.���!�ѫ�m���:j�5MO��B��E���[(�z\=���:�t��A!�J:˼���9�c���{_��H	���;,ЯwD�������a�Gh��VWf��3���>28�nw�|�B���Z�������\�Q�tc���(E{vIz�P�dyv�{�'�yE�[à��ƒ�y���e���9�\��`���4��\����^~�y�Ut��^�3��%�2_,�j�������5��nQ2��|�02+0J.�wu�Z�S����;l�ߐk�R=f�HL�G�]"�m6S;��SA'��fY��+,�Z���ZO"����gx���"���X��	�����6v]\��;߇�����>���LV�ސ�}�c`��|~iw� ����_�:ơVP�����n��M��\5���a���� KMk?V�����	S��9��:�=[��|�ut��@�c7f�ҵ�(Ӊ���C!o��hcnu�j�lZ�%���jꋇ�U�2¼���}�]�|1]m�)��1za'�g�������C�ߠ	N�2�'`F�0��Ы&.V��wi��6�+o ��At�O��cO����{vU&9����76<֝#r2�~���X�e��g�\��`M�+�f����D5��y}+g5P�7��&)��z�#���v;�ܸOF/���Ä"O�>�1A�����bА_�Yx���R/���G�<DN�h>�S�e�i]�Nr�yd\�{*�a����7�ن����و	���/%�=b�]!������Gur4�J��\]�U�4�tz��g�}��ZO�z�Ǒ��m{���`��'��
j^���H�^�.#�OR���m+�U0�{${����[[w|~K�v�ɴm���zW���bhBc\t�<�K�C�^�jb�{_Y�O�iq�?��K��Y� 0Ղd"o�¦Y;�"�U�pt�P���F\z*�ظ���̸WS��!O=Gk�@�Oe��Y�}�E��W��xxW�T2��>����~�'U�:���-{[˚��c3b�]-��n�'߉C���~�'�*i0g=�Ӯc�q|MCr���&�8Y�&R�rs[-�.k��՛R�@!��&a���!0i��ی����#o�WH���UoZ'^�Ny���kOgh�J38堇b%���YX���u��u"��E�v}�r��Eu
}�.���r\�c�:��A�.���HH��^����x����@fp��9�Bp��z2z�oMV4�:(�<*���v	�v�.5z�s03=�� �]4�mA�ai�B�˽��s�D�p]�+K�K�3K�-={�d[U�pbr��:��ٳo��0��)���1��|��b��ojЅ�����-M�������Ǫ�ec�I�+��t��T�Zis��}G��� �3��~�k	ĵ�B�%^��I������(,-���#)�*��*c
ް1�f򣍕�)ZLO�X��\g�<lV1�V}���2�����Q)����3N^�f���P�]�M�7����(=��p5��h����5�"ȲoZ¼����χ��>D:��:
���w�ˇ���\��b��:aNvA[��=�6�X����iK��T'2�.��]j�bb�#��B x�U�E���X�7Y�e�c������2�M�6{�M�h����s����A鐗jV�l���'7�����<�����Gx$���t}�-:aauJ.��]{;}�;;���HL���5��ٔ�]��'lg"�ܑ*��x�+����1i�rrą��2�֜KGt�h�i�jWcfN3:*��&y�-ig���.�`�֟n#K͘Uݙ{�1��J�s�Y�Kӹ�6wD�flSF^�ݿ���;#`#���v㇞� Qy�^�,	�X�
�^��\������Zۉ�W`A�-�k��~��A�y�b�Q'�������~Գ˒ɞ��u�m&����^�u�Ǫ��ǀ����軶���d�n���[{��GU�+)�׫4����Kʭ�7�|PP��	wN�����%M�~k��슮qg�#��|[@dni��ۻ��4� �f�`�����+�����xh�I�,�]��������>2OB^������Ҡ�H�7�Fu�C/�>w����d8�ΎR��'7��fj��f~Zy&`dK�e:����=4=�_�����N�w($>���D���d<��|SS0�W@���6�)��e��o2�w��
��z`4/U�d<&<wS��Β�Aā���ŗt�xi�\�؂�v�S�.��i3Ou�S��
On�4�3��#ʶ[�6����͜3[M=�<���*�[x[�};&N��z�2I����z.S[$��\9���P��^�{���jݨ�3�'GPV��}2m���[���rCg���.��U�#Ko4��XY̐Bī��J�b����J{���i@��
+:q	ǧf5��9C7���۲e��h`Iu�V�Jy�7^�5�Jf��)ʶ�#�p��:j��^�c#�;:�t�F���F��׵,S�9�5�p�qo%,��Z�1��'j��r�+&j�N�����s��]�Y�!o,wZ'h�K��놘}n̷q`7z���n /⊒��	�zN�)��6��ű�������)�+���c4v��+I�� P�bm!�u�gn��f�9wg��9���k+��P~���d�:�Ew]���v^Nd"����!fT�Y�v���u�����d<H$e�-�7�|�G��۾�u7kч�s�m
���g@D�ݴ��j�P�An9�l���91��+4���6�g�9�$(A�^��+�Q���g�w2>���Ah_rgw���I����8��C��%X$[n�TTCl����"�]�;�����\ٖ�q�_K�q�s�V];�#.�2��&"���q�{ݺ%u���ZgoJ�xxA	cwF�t�N���|�{���Vl�g�����y���f����FVo�V<�'sm��O<`�{��a��
:O:v���T��J��}_"jRl�R��y>ʛ�*5,WUfu�5V%�ݹ�(�.�]%�w��Yc��_Ez_-�Z��i�����*�	I�Fe��Iz�vi�H�3^�S"Z,�v])��]����{{���sw�T�	����b;�t���Ի�O'�9r�3mq\��%-T��g!������ZjV^c�5�H�u	s,
�N�c��u��䶦����PYP�ym\�9sYFT4��d<5k����&�:bb�S�S��}�z'yO.�i�)\����R�AVj-�W ��-����Us ;C�U��SM�a�:��'���F������ȕ�Ἃ۝⼦��Ls/_�9����]�ϳ�L�� 
�p��΄�"hS�r��1̬�	wP�p��.r!]�`�w�_ug�iq��ʶ^�ܨ/V�	�1V������T�Z��M�\���S�����2��r���e���Bny�ȬPӧ�;:�ʳ��h�L�`-o�T;1r��T���MN.�/H��׵]���X�g��h��qЋ&7]�68�*���E��V�K¦
r�������2Τ�83|ק���}��$��*{TH��㏯]<|z��qǯ�8�o��<l�
� ���fŶ[���:�êa*���'`u�����>8㎜q��}qƟ_^<x��$$w���/�ȼ";(�2EBI	HU�M�}}m��8�q���i�Ǐ6����ITm��n{e�YՄڢ�B:���9;�;���'m��S[������w>K�����ֆ��|y�e2��ڷ;m[Z�vt^g^�\Snם�M��~��
<�|����N�Zh��:3&�6���ݍ�����m��n�g6���􋼛ɦ���se��������dB;��[_������5;_�^�<��BC�m�[��v�Ȅ���,���z�-H����^3�k�[��nw�u�{�����(^�yg���h�U����Y���8��<��h�����<�a�%ȎK63�����	�R)��-�ä�"�Ҟ��\�Q���ex2iSV�<�a�(d��w���s�G@�v��OU$�<��a�.6;�}�@S�g-�G�����J�s���@.�D�粌�+T���j;Z�=���{w�x..�xM�ՊD��%L���s�8a�"K���[+	*�z�4�v׵}lu�3�H�jJ�=���?tqiM;����e5�M��皷�����m�(Ϩ%e���%˶?�f�������6�`��ǣϞ"Ksz��n�p!<��5ϟ�%�?h05�Z^F­ڃT�bZ�2�wo��m���VD��.�A}��}I1��
�{=�о��攋�g�y��e�F�3Vf�߹��X�`u4��C�>!wTx�}۪���cܮ�����5����r鿖̮�ڄ���gP����&��=RCŎ�$��@��y�;E�__ϝv���sR㗎���_i�d��&'�X�c�O��kpj實Ph��AX+��N�^�VAF�Q�q�5�6ԧE�+^p���J�{�	���\6�|vG�<w3e@U�j�MFv��5]l����K��4x�A>I
6��g�4wj� ���y�u����m���W{{�9R�K������2�؛��y쭮V:4��[3s��y�����m��o���>��b�w�������bk�`�1�a��Fy�������;��<3�y.��ɉ��ո'vU���L���zۯ� �*8�v_�N��O��Hý�"+�T�k��8W֗�fs9�	�	��T�w���4���Mi͌�8u�#v	~@A�ٮ�a<E?��3�Eg�N������j����	��d?��>꿔as�QMI�qt8�Vz�B�e].������CVM�H��<��ɶ\���홹|�U�#/��£ .����,��##�'W1�]�Zڽ}�q�����9�ޘ�u�����\؉.,P��ާ֫�Y�,�1�ܞ���
�gǆ���hn����zѩjP%o���'#A��y�νF4ګ��E���u�iࣼ�JvFì|�)�fy��7k��'I#R�$�6cJ�����\o.e����� �_�^����E<:���3"���JۤRz���q�:l$y�����l�{v��YM١�|X�����W��?�������$+$�N�q(�2�?];��z��#C{�z��l\���d����d�	���EjNi�˗�޶��3�oYer�b-WHZ�ϝ�<{;�uK�&��=�J�� �Qp��`�{��(����;�e[��	��4�>#��{�g�k,?�۝5m�/rZΝ;�wֈ�t�����\eN���lk��ط��Ӻ^e��Mj����EQC�,-������s0��+�x	օm�nT0��)�Z{��',uq��8���&5��Lk�xw�6��l�g� �[x3 z��Frq�-�N�R;%��v8�,-to�9�T+�!��G�?�%C �|L�~���B7T=��`�����qF�k���7�^:����*	{kU��vW5��+�*]�<�X�s���b��;%���^{� ωz:���D������3����ֽ�0'hC�7M��6{+j_T���~}J�W�J��	��4�.�{ϩ��(8����ZFä7:�w���G+�]g߂�z��Ǿ+��?o�f�UƘ^Po�(�ì?�.u@��(5����	�aJj�K�S��zT4z��-z&�L�M����k��P�/mBbyɮ�]p0����>:�;fe'�����7![�Pэ����"�=���)t��mLP�a��,r���������؞�x"\!��q>�aB�|5T�j��p�./e�~*W8z�m~jx�0m�������$�A\������[��6%��6/ۿj���mù�{w6.*I��'��r�a]�{fR66�:L�;}-�hn����=@=�s����`O����-5׽�ݼ�oI�-�sL�-�|�(�̽�������<�a��A�� ���R��|5�y0��T++�~_���暾�b" �&��-��R{����u��ܯk{�Y�b�.�S��4�ʏ�|��i��" #>
]�I�τO7s�y2�N�^��1>v�k"��#�L���_j����i8����~�} �u��+��h��e3%�B3{�ۖg\�xc�v=�r������q�w0^�È�������:������XEc���%��H��˼����s�~���m((�kU�/�.��v�"���L�X��(��|e��^��w�PX��ִא��3�Y6�>ç�˕}���̘>�i�!4�xO�1��;�о+�x�YB]���c��L�R�����
���j��9�����B�
�C�m��$Kt��s
�r��S��/��z^͇����p�9r3��f{`0g+�"@�[�GW�$���u�Gld��]	���&|�{4�=/�N���z�ÚAGo�h��a7�=�Ma����r���#)���R�w� ��jC𶮖�@c(�X�9�}�} ڧvk�Z���w��+�Q�*���_bվ�Q��!�lf7]�-�{�bĲ9׻�36�n����iDN��n��ýe\�P
�L��͕�uj�ӎ$�Պ����^��p���|�ؖp�j��������Ͼf����p(t��h�&��i���_�C�/kkډ�ӯ��Z�k��y���6��u�|�c,��{}p�ϣӑ|gd
g�n�q�-.<Q�;���!,���4��{���)ut��	sk���ꃢ��MHK�}Y]�iN�<��K��;q3��
�XjO�����v������%#�ʒ�`��0n>�.�^�f�._3pf����쾨���6"T,/���U����K�N����C�V�<Ҳ�x3
��Fk���Ż�5�Ix�0��n�z����vg��H����:��Zu��s���eʳ9��ie���.(������+T�UyG[�W=���{w�H0���k��&�%?nך�M3t	2�N�)�`!5]Bd^�"K��K$�K_���ȟv�â��u�-��O,��s3mCFt��î��6z�$�t�&�hl%rÚ�1����eGa�"��rs�`�>u1l��4DCA�l?ܸ��z9��[ׁ1i�`?��=���.��ϿG�v��7z(�Mim#��%(%��Y�[��-c��ˏe��Ȱ�n�4�r��cD�9��{�b���q��AY���2����n�L�������=��pmwN˓m���6��;N���I6�w\q�����<�oz��Q�ۑKri��Z��xy��CKO�=L�q�}as_��dz�%b�vP���p)B��vN��ť5ﻯ5W�)(8����$'�H��[W�1�RS�Q\���2��v�S�-�Pu�̽k���ҟ1�r��A�"�H�$<�M�u�s�rx�gm�i�3N�ḱ'B7���-o?H>oK�Yk�lR:�y�t0��E��'ob%h���KP����%�>H�#'rRznp_��W�v�ƹ����`/B���B���ژɵ}S}�58z&��,�v�
������E�yD�p�6|&c��5��~���g�dyT�߸ͼ��y��ǹ�G�O��堄g%���QPS�=5�8����Ѝ؏~�[{�s�6^�J�z֊��&����i�}k*�KOՐ����-[�����������R���(����o�bD�������Z�\����l��[;y4���D��a�wk����T�$c�ꦬ�[�q(��4�KK�8��G\ƽ�֕_u�>�����+��_�����ٴ�߳��(f�\k�K���2�`Z1$�1t���H~�8�v|���#�=QV�8ȳU�.��-D��B�D.���K�e'P��V%N\a�{�{�BJ�d��8��y%�47,���gg3F���ޓeF��u��9ot�{:��S��� �e)[�F��Π�Ó��|�v��c���EF���J9�{���k���sWR{�?��W8��}lml��pco`�&V��\�,)�{�m�^��yS�Gp��qE�n���t�� ��kڹh�S��.?�k��+=	)��"%JN.ۧac�yM�*��WT>��,��h��zC�E(I�C��j9��D@�+eU'1���)��η�ɨ������z��z��H�?�GW�׎F��F(<�>��I�$�p�m.r��a=�`-N:&)�u��,�c;>�X��R����3�/�3�[^���1�h�d�^���7��f!�I�P8l0k~z�=�3):.X���0L���>;7�ט:m٨Ǿ�+���'��Wq^K����ݓ��߸�,(Z~���\��=��4�׆8`�s��t��j�m�����ͬ~�)M501�E�^k~x����fW=�����k�QܚdS��p��cj�j������39L�������-�8�=��;��i��X�4�SO���ж]�9����?VAϒ``�	�����Yk�;�d�.��]!����ܼ=�O��2��k�ٻ��8`���.���'�<�n8~��%>���7R�}Yj��u/�,Z�͙�+�W�qW�,�G�$0�]�j���>]�ku	m�7yܱv�t�[��;��d�s#]�juƺ'�gn�!��7�z���k��ق�v�z���{C�Z���Q��:�Ω�S�XdT[#�f�Cĭrf[-�)�?��`��%�;�'�U�=>��V��1:L�q�|:����P��������L�e�$I>z��"�ThZ���o�8y�N��E���|t��#c�����wN�{g�fd6#��
�pj.�.��	q5"� ħ��g8��AQR����0�m]�V��ơ׷D�(������}E�ϼ��A�z�������@L�t����1�g�j��'��nW�q]��I-{���Å�f^4�^�	H��I��i�mf24&|�EF?i/�<���<��z���0L�Q�|@Vx|�[R���B���W(F<X�cG*��i#v�Y��Z�;���j�%�1�9N�����(=���=�p�zO��a�kf	���$�Fwj�ٽ ����y�,F�C�gιi�ta�Afa~}�w�ʭ��nU�1y=�� ��2%�j�|fzb ����',O��ִא�*�����R�	M%�S4�4)�\s�ʼ�c�"��B{� ��ۍ�3�{-��<[7}��+�5�'�~��y�{�60��iǞ�M_hۄ�e��l���8��L�䮴��ު{�*in�1gA���wb�E�w��ɽ�����0�{���YM\���D�CƐ!x�σ�oi��i���9�H��Q��Z�e	eg���m�ك,���m��u�ƽ;Ƙ�X/s���Z�<�$��ZEn�{d���u�����K7sHS�V�����/����|5:�F�/>y�G8�T=���_a/Q�i�t7Y�|�}#ʺ %��n:�vc��~�RG��L:����K�鼇]��MO�t�z!Q����<ʼ��4; ��=�*3�R8��sμ����4�Fte���p�q3g�l˔B>�}꡽,u�P��*�;Y~ʦN��>��w'�~���o�~2�1����2}n�ʂ|_�w�#r�A��T]�8ms��Mo��'-Qt9��K�=�ֆ��2(R�r���z����
��_���r���)�n㘙=�4��r��:���evl����ax�������vG{W>;m���C���K��]9�� 9N-^Y*����馞�fA8�X&�c�E�4�F�)m���y�̆{�v�z���i>�*We5Ai���@kZ#��.�� ��N;Z�T͜�6�k��P���8\vɋ��T�.�Q�yw�n[�zr�b}��"z���.���{(�˱���TTغ�_u�y;�'��`���w�w������9���,�b\�Ȥ����*������ȣ��y�Q�pf:5Z�s&���:kg{�S�S	�
�l�nv�����t��^H���{���{'�7���Dx�2�D�����4BA	�t��uVj���I[s��6MyvSf��9N>��޵n������inOWН�Y��b���m�u�i��ڊ]]����{�����X�G\���ֆJ#zDB":6G�Ԇ,�Z�ĵ�������!ϷR�+���x.�mt�=��#���L� Od�,C\I;&�<�h3��m�3�yn���M�M&��L�,�oV�V3^�~��4��4�w�6�oF�2a��l��յϫh9��3�/�k+�6��M6�;�;�L��5��4�^e��-�@9n6���tqc��ǀ���U�8�{cbg.��h�HT5�0�!�
�z�/壕���}������x6����];112�E�}Hwb6�Td�W���OԹ
Z��ҁE��J�t�nǾ���t�m���������q��f��$���k����e�5���|Ǝ�v'�x��].�%�����W�e���|���\}#r�d;�X�v0P�*���"��I�(�����P�.1OW�7>�;d�a�[��SE����[��T�J�S��xr��w b�.����2LV���h�<�Լ0��Q����4N��/�mm`V����<\�,�2��۝ۙ�����ݿF� ^Y�m��ľ��o)�tZ@\��dnZrnF�S�m���$"z�6j�l��wv<��_�1Uh��ߔ;+��ReU�5[�1	��s�Ac���;ۆ�m�)-�-�޼�^�\��N�pv�wv�*駙�/�E&�g`�Kw�G��7�޽x�b)M��|�ȶ�I�0D���M{���,���նt���}E����+��e�n����ӕV%f�-�
�K��o(�:f0 �G]�"���%wϺ�Rol�kx3�De��O����fϐS2�3��v���JhcD�"�oP�=����Ǹ�l$��t0`Bi�EI�X�/4`���p��f��j�;Jਊĵ�FnΧ���.�%i��p=Ce��]�r�q��Փ�G,@�T)��Zy���=�E��ط#��%�d�Z՗b�����P�1 �V�X0U�l�|�rx+m����Р�Z�$��\B�3&4q�髩�T�d��:��b̽�C�b}��@
��_)�if-\�mԢ �0�m�V8�u� MX	rX�L�2���NQ�+��W^����Yɢ.�!��'��s���W�g.{[�l[�]M�iЛ9��.�d|����A��[�p��n^q���9�(��.6���Q�2e�)�Qe��y}a�����&��Sz��<��x�yg��OVMC����\GfV<ح�%@Q�����\'�4w�;��z��(*J���k�\���e�|�ò֯Bg_J�R��%j�9�΄�CRsF�hW\^���	�����س�?��>� �ů������Q�5X�K�	fv3w�����g`w���3�Z�+�[�1N� �܎^F���W�"+�*��DdC�#C�����2^��ob
��2��o��,\��z����%�K��x4����v#�ɪ�YD�wƸ�{�w�:�EÏK���d������7�9�oj�=(GPJ���9aVݕ}�v�lR������Vc=��4�Eu�FA���&,+sF�E�@Q��srk��Bz�A����X`r��0ed��q��\�f��ű��#:�B˅l�O������p�n���]Vdr�=��'���
(Q��n+:�.62�K;#�n$FC6���oq���^�N1��nڳRUTjT�%B�Q*�4q3Y�k-�N�m��
�UT�RJ����}t������8�q�����۷ms{tTE�w������μ���J�ud�UP#�}t�����q�8�ׯ_G��nݶh�U$���ff��׻�Y�le��W��b�hٴ��ڂ[6�,"g��7i� ��X6��ͦ������O���Ks���8c�m�k��/�wn���bY�Ͳ���k~�{څ|��n�N;5�ӯ[K��h�p��{�v����rN�rJXv��a��r�뛔�Ŷ�G@L���@�t����":N:tVMl����>kW�/5$�8ND'O��{���-o���'$H�[�����R��~,�q�3���[����~ϯ����>�ȕj"�7!l���H�BBYN���I�bJE��$�C��0�xkz�:,��;�2�V��x���U�\��.��p9�8h-��^%"�����"��Z�+sm�B�%8���1�j�$D"q�)�E)a�[)�(A`/�)?�IBҌ���@Y����@n6�aBP�H����@�L��t]�,����ʚ��*�ZѨ�1�F\!ɗ^��q�
�������߶����^4*�8�w,9�a��h��5w�@<P���<�F��N�5��N��G,�f\<��ʋfاf���9�jg���|N�'�rۯ.�sCm33���y���N�'h�u1���Ėz�ݟ%�$)R	o�h��b�Y&Z�n�:�a&�P���~i\�чG5����/�B��s���N���SÚY��>NJۢ&$�gs�����ϼ$GC���S�����i8)t�<�|{3[md��ޙ���8����K`3�;�8�S5�C�=�k(��).*�>���=�R�Ou�5�]��Gf@-�J��B�7���K��`�Ȏ��y}{P�����Ũ���H��y��:�e�N�f��S�W�Q�h�u�5������v.�vi�'��q���j2�� ����8ip��\<f%9C~�;8n���?!�ʨv��I.��e��|��e��R������X
z��u�S����A����Yx�|�~!�;6Y㠰���[��>$l��V*���+��>��e��Ǧw�UU'�uucXl��^|���-��}7ui�b�X���5����0�ᓮ�I�������ͮʡL!�}��o7��o~2M��n4�k�U�Q����~�MP�\��r�
�u^׺X�b}d�V�[������y�y.�Gi�^	RG=�k�_���W{��1���ǖ ���[s�Q�l'�^�X�[�^�y���C��9�9Xz��o[s|�H�tUPz�M�wT&�=Y�2��G�{�h1���x�h�9�`
Mt*D�t鉞�ܺ�R�; �9#���L�9�5��q�V��g�\c,WQ홭������ᙦ|����I�6+Z��́{�+��LZ�ܸ̚���ڞɟDԫ��3+�E�t���{t���Y��x�7|�ɚ�p+����z��p*���T3�2,�t/xsg�c[թ��f7�.�hD�G����0���S�lR�����T;JC/��z"���]S����ǔ�l���SO�Mn�q�1�ܹ+�X��[��32�W�ޅ�ou�;�6�%3S��>�\�O��X��%9�����tu�\6��"۫�/��rԇ�L䜭r7��"��6my�iZ�g�ޢU;�q���ɧ�%`�v���6=�٬O�#��T������_�w�.�w{yri��O���>#���7Q�9޻% �ҁ,���w^]q�JU^v�����e�hq�H��ޥ�-��re6ֿ�Hh�ѺXMH#
��$��)l�+	m�����y��wt��|�2��E�u�F��j� ���>��^�%h�*�t�gl�_K1}�fj�{�+d;D⥁����`8vL#�}^�h�<��RI 7��ħZ��s"xM��9�OKJj>YA�k2U�#ۈ�1�c}+K�5��X�89㦷�a�����ڸ�V�����{}A���*����l��ms�)y�{�D�7�&�ƦA�37 e-�vt�8�|�2�2����x)�5(��[TzH��Ύ���鮐�9�s�M�,�/c�c��yl�{������"A�d�f���++[��GYCñ�o���@oQϿ-�NG�9�_s�a@C=�/+M���Ÿۢ���:E�$�q�\�OW/��a67���;=NWj4X�L����C��ڙ� �ړGM���4��yWL@��١g�I��Yͳ�6��֊;tVXY�E�d�v\8-�һtw�����7E�.�!�>��2��N��|��O���<�a��x6I�-��ܿK����2$�n[��T"�7Q7=��-���c�у{r/;�5��Pا@d5XQJ�7z-Ez9�z.�Q���[P�B(��Q�`N�̵7��C�33p���I֑�J}t�a�
���l���`��9��2 xR�Sӗ<y���5���O��'oٗ��L�Uޱy�[�7��pܛ;�vq�`]]��k�IU)3>:}y�ަ��fA�KiAr�|緸9�01���
�GG���ʼJ�IT��te�*,�513��q�����K������lM?���ݞ��R=�}�\ 
��(����^���T^�ꗭ;��vf�D0mٮװn�S�O�s�+;��^�ұ��V'Z;x�籷F�9�Gl�����c�7��_�k`-�q����X�]R�@;�跒S�/B;����f�`�<�=Ǎtv���Čm}�n���j��]�z��%m}ތA5�ե�����'O��iD�m��D��oB]	�|�9����Y�N&U*X������6�/h��E����iUwo
9�ϣ�xcA�H������QFtS���y	6�w
7�fҝ��:�c��z�+�¼<=�jx�S��"F�*�p�9���k9os��U�,�aA�Y=2�FL�i��Я�iLNo4�w�M%S�-��3l���Wx���Q�����"'�m����j��յǺ���쬑�3ϼ�s���S�uH���k��YCu�1i�[��*�����ە��dXv�|�Η�-�on 5؂�
g&͉4�{?�����a^[q��E��ݰ���)�z����>x���E���xV�H���U�X�9��{{���{ <�yn*�}��B�U#8�e�JmHl֛,_	��V�=p+�W��HIG�K���#-r�8��2�+m�s[G.'(�抄�خ�Q��a�^��2q��xr`�WS��\��}ٛ�i�Q����\'l*Fw6<� �vǉ��^��
�]������t3{*/"]	���fCZ��O[�۶����EZ��W�w*'��
�jF��ߘ�{�p��}+�\��,�@Z�屬J̅tl�4��	�EgeV�[6{���k�����)U�����+9��i=�xb=/2�K}��t��y�@Pp깦�����c��Bm
ȸ���v:����o0�y���-����]��˧�;2$[��Ϡ�����͌�0$^[7Uy��d�of���O{X�%�ۥHH���U9��l�������'["gCt�l���4���?Nxo:�sf�����9�J�!�O�{G���~�~�j�nRE�.ڐ�����_�W�]g�����,��A�u���@�IW��;V�`�hMP�Ԟ.ͷ[���}gJ���/��zj��*����vF��ZI�ׁkvC�Ve�hl�i��ba�Ӹ^K�E{�VT��>��Ž�J���3a6��z�.ψ��k���Ы��5@p�&|Ion�F^A�Om��@����׹#:2}����4��h�|��� ���ߪi�ԋ��l���pڭ�9��; �{�G_|�l3��3�+����{�~���)��UW��d��I�&�bA�Q�y~�[{]�ս�
�M܁�*~\���� 싢��y��Zw[IHqJY{�]�p0��J~<t��i�us�_P �^tƕt�]N�L*���Ba��m���j��X�F�����)Z3Z�Fs����{����/���]�oC�5q�Y߽<<<=C�'��w;]��RE��<�wXr��]���}+����i���tZ�[=���֋��FY��G����p�s�q|����.n��ʉ9�3&EM�Q��ݻL{���`�T]�����Ly�:U�"��|d�x���Q9�z"fU��1�J�4#��v�B�p�^3��&ؕD�`�����sV���Џ�û��û�N�Г��\x%���KS�M3�@7	��\�;I�Z�UŮ;4qx�7u�)g+�7��<O���|���+_b5�i�4ս[��2��t�!��{��Mx�6=�l6����h�h�q �I�x�ٙ0��}��~��wp�Y��ܾ�"�ɠW~敫����\;�#��gޮ�2�KK6h`��כԮc�>�>}�Y��`�״t���}k��>�J�~W�����H\J�S9�LN��q�Fp33#A[8����ާH!N������1[c{1�a�7�n�Ơ�vV6�sH&�8D�J7GCQ�d]��U���xrL�jk�N��ZQ���>>�n��F*}��xh�0!��ۙ���o�1e3�̆�m����k�b���֒�����x�[7w�Rs���x����������R�o5��Q5�=�y+w�h)�ٓ�q�ۋ*)���tbn�:��l�'��r��g���_�Kz��>�\���Y���b|��,�ʞ�r �H�F�@Y|�1�u�lr��ӯ�f�����=��d�c��z]��}���;Y՛�_^Jtcz������R�i�h�f��o"�����Dg_��Z�3�>�o7�T����࠶O:�J`LNGi��{5�'��Ւ�e�s�!=��7"�6���v��OC3;�K	�i�t��J8ۛK��˛���q|�x��1��6�:��_f{9[��uZPD+�$�{hxގ2}sNg� ��0��O�O�}trkz��z���B'�Nʫ��7��Nx��v�H=y<���:'W.�[���^�u��b��nD[����d���b^
���N�T����D^i;]����s,�[.NP�}˭���K��݃��Գ/'�����Ի@�h���M�{6{�B��A�+uՈ�T��5`1o���)�e�M�Ê�)֫�F�w3��}|�@�5s�2ubd=0�l���8[''�L�k�U�_�������U�<�,�0�����=�7'Z�k�
���a�/�RgA�sx����=�HaBƼ.R����>��)�a�r���&y+ˍcz�"gms�ي�=�5��1*G�n�R
��!l�8l
sV������z��\;���#��j��Ɨd��9��C��R;�/d���>�[&5�b�g1���MRo�֝y�7��l$L��r� �w�s�O����|�vȴ��}��f�{0��L�I��>���5\yH�w�M(UY3�3g���kV P������̔�����l}[\_��0�ecU���̛�CI��tL�^��-�7�<���r��p6���d׸�ه��Q���Yb��Y�7YXF�e�g�[�u]^�)P�`��E�w,�P2)��s��q\}��ڨ$�tOH��fk���pE�煮a���**���<��k]�j̎f�f�H����6	�AO��"^��U�ӑ�,�(�pt�f%�IR\����8�3Ȓ~$�}i�y֪k��ۗ���"�e�fŢ=��Н���ܴw��e�j����ω�۝u��.�wn�pv�;�*W>Eh�a�m���D�Ը�H�
�y[�&[��L�G߼�<<<<=_����j�R�N)}��O%H&�t�ڭ����;��Dn��{��k[��
#��1}�)G�6�WS�T���fMq:�>�D��ܮyV��I��p� -�4���݇�z�`��$���68��f�I����%��s�������o�⭭c��G�(�p�L�ǆ��^�, ��Ԗ�0�r7�z&#!�3�K/Cv�i�j��ܷR;2$[�^K���(���r�j��.��c����7JH�m>���oR3�h�tؠNH�����X?�>'+�LHܒhv���Ԗ����a��,�}a���.�[gWpN�
��E�6Ѫ8z&���yW��})�z�`�lQ!�#VfR�O���O�k����U��Y��%+��)���(Ξ}7��a�7�h��Cy���Tv)eOGڲG�Ȫ�vǓq�X}�]��t�1�J�͒i�a�6>��S����lK��lN,�:�m��z�
�W>�uJ&�t�ɖι�C��Z��-άʻ�3����9�l�w&��,�8�S2�V�x���M�y�3�D�E ˺��ʃ�X6�<��33^�]u2���FS�[C�#�C�&*˦A�4�GV7a���'�X��38�VP���v�F�cZ�¯���t^��Z��r4�"��ngY���ff�A����
��G*���&�[\yv_k9'gAJM� �@�dY������U���s1��;�́S���ǝozaʊ���$U��s^YBg�AQ�3f�mp"u��(*���-�x�0�(���O�sY�rVK�2q�o+��{��lU�����T���'I���L�����v�����l�r'c��t7U����
Vޜ��Fq�V9b�}94\9���ݒ�s��hplu�ky�M��S�7CT�3^Þ����F�ۘ���p{Kh�en];ow��#�ґ�.�m��y���6�IH�\��P�[K�vR���ܘ�A��W2�F78����v��h�l�u�u�v=(_8C
��X3'��ba�2�b!�ꛎ��k�F�WMGSEٵ�T{z)��:������yW(E29hFd����s��%�ץF�����wd�Y�ڨVk-�ʑvZ1�����0<�tx�ȋ�L��n��n��Տ�`�~����L�[[��,��7nw
N^k&֢�8Z;J%^v�$ZB�@�A�R^��
����Y���}�]��-�EN��,��s�`��a�}�0M9v9Lޔ2h����r#H��=D"��T�VL�m�b;;%�n����Qh{W�jY�;s�/T�y谺8:�����L�b}�wf��V�����C_(wC	��R��I�t���{Tބg9Y�T�0����C��!��-��^��Cs{`��L��ܾՈc��43��ҿmv�1ܹ��{�ѼCV�҅r�h��<�d���vis�W�e܎����J��s|�i�'�B�)��k*��OgDe��A;{�8��m)�yT�C.t֎�KUZ�
��#���[�g'���R{x;�:o17K��o;����ڶwQ�&X�[��4�Y2kΫc�u�]u�36�5�nωW	��Z8*�U��s'.X.�2���t3ozWt�4��ἷ�[�R���M(��aR�$nR�_!�Vy ޫ�}N�b�)�
W�`D<7]�DCOy������s�g�s���i��1�]���[�Ϥ̚侚I��|0��{9��pܚ{6���R(]Iu��I �@�$5��O�$?��M��J<mӪ��I!�:x������q�=z��}|v�ۚ6�ԁ�ZGTRBk��'9�޶6�O�Q��HI$5^�<m��O��8�<qǯ^����ݻoA$���T�Bꤐft�(���!9m�$� I�Ǎ��i��8�q�ׯ���n��rI7���,	$$���ӑI�?�����Y'm�*�X[k��$��[b�$�����V�kw�U�s�rJ?�	'B'�[欂,m�Q%s�^Ey�Fu���ä�����ܬ��dTGY�fQmڔ�ܜ���;��ﯚ�;}=yΈ��9�bsl��󻳼��ͳc��pv��t�[j��=��Ĝ�;(N���*8���Ί���r��t�Pl��r�i��AڕUm(Q��q�l���n�,���;t({�u�_����}������?�P�r�I�;O�~[POn���goG��;2ɮ �f[��Z��9�Y���r�Uu��3��1�;��4��m���|�jL��d��k�-�x�y���A}����,rx��^��`v"zP喪j/;0?+�x��3�p�go�V%�1�����$�7ė�O��y~�]�t���n-����3�f� �l�z*bg�]swg��J��ۅ��,��l{7�7��^�>�=�����m�?�#w�	ń�2�xj��Qy�1�xs��E�+�~��r)�A��,�%^�i�0,���s{��Q:��,2�õ]SNv�W^�/V�sЕ�\K9tl5�`=ՍM�w��1x^�Gk�*ɴ�)J��j��d�<�C3rn���4ZJ�g��mAq6��b�h�AT�z�E_���Z��x���=��r��x+�㠸�U���ν�w#�K�b/e餝�n��J�e����&wse�VcH}�������۵Y�����LO�ۂ��`uuh���jR�=�^ș�[y�p���Z�����f3m�������Ym<0/7����xc�m��1<�ˇo�=:u�����a06�թb4�Xn���wu\�����cg3e��	�y��B�@��ܳ
��e�ޕ��C��P����"��^0p٨x�>a`���|���d�}6<�T���hn#S�4ЩЋ�.*�.�O������t϶+��������-�a����Ǹ��3]������M'4��0>�<��Z��=A��D�XT�nFR��0>�qΌ�.��fJ{���.R���z�^�{c����3|O?�ǣ�6�7v�l�A��ޖ�'4���RC�Ɂ��M���~��n����r]T��J9&����>�j�+C������6@ܾ~�tqcT�F+j���}�t��1O���ފ�����܋�z��]K��%@E\����xj���ݜ��v:�.r�i���8h���/����x`Bv�F�tvbB� �9M;�;û3jt[�ѱ��Ҥ�:�}�oj���aה%�o3��;N
��\�ef��0k{MN���i�������*Ê��3��g�}ϱ���ל�|��v��٠���Qwy��kR��r�}�I!�c��IG��w�{��r��<ߔ�4��6|�s�I�#u���L4�sx���+o�Ő�X�T�E	���DWj�!HJ����m�]2��S��n ��x�3��L�DƇ���v��f�R
��	[�_�k�{vni̊�1=���{jc FX�������"9V��6ƏJT��AI�j�$��y}f���÷�(zA&��`ʄ:�&sF��d�Ǩk�* �]�x7����!M�q�|�O������t�Pg�(~
sVz��wJI�X�S��p�bj��	����������xnW�["8l
r�_2���S6m\���O��'���K�[�Yϒ;\x	Oݞ~�6!��X7�GC��''��@��q�][���k�k7\֠��]һ;�[]����FAr0�f��k�B@����>�~� Y�U�����[�T��s�A�d�Rfaf	�$���
�2#n(ߩPؓ��}�.�=�ی1Z�����Q��ز�j�r�����������ƶ�o��1��$��\���tڊ�eWx���ghX��)��W�Jy2��e�ԱEj�K�m�|os����VC���a���]���A]�v�o*�S�;�%�/�~>o7�����n;�䚸*�5��0��� ��F�dQ�\�m+�ϲsv�˗ԍ�g�{��/77`1Y�9�)꺄qJ�dN0���n���L��A�]o2���θ뛥{�������o�����1;��Z���[�t��>��u�;��%!�D����s#E��#2���ru^f�Rk�M��P�����@J��{�Jf|���X1c�-����RO`s�ݬ˯�C�#�<�U���s�Ҫ�H��+ԊZ�����;LXf�wv}�o֚�3�ޒ�삳.Ŷ7�#�����j���T=ɖ�=�����.̐:i��=4΁�Pm�]py[���YE��zF�S�;[�.P�t.�QRa��ᖨn�́X��eBI͎j���:�v�?HCk��m���ۦ$L��og��y127!�#.�l𺮳(s�@���]��<������۔8i����8���4�ɒ������C__�ʞ��NL����B3Y�L���N�Õ6�t�qU�4oQv'Ww�q^�#�d�b�ԬI�5�xi�][.-nr&��}�5E¿yxxxW���s�_�/��F���(U� ۞7��J���#�y����<��3u�ʙ���1�	G �@��F6EV�7}�(�U�I�/���,����xb:o����C�^�bbT�^2s���+��ۏ�S��n=����z���i<L]������&�pͦ�]>��:�G�h5v��5�0m�/;�uSD��L̾��k�<(�~ɛ+H�>_���-�50ڻ���T��5�|�5��;��x�NW��N�=tɠ�46��]Awl���1w=腽�u�)�WC�L�c���t�x��vwc�:�b�%��*���X;��>��&�E^�1��žGvIIx��M
�A��S+���gfj�>��~�����L4��ݸ�<�ZO�#DA/l�`l�e��xN�˞C��]�-�AK]���i�+�OL`X���U�����Sv�WV�[Y6�����ߟ9��;�<�і��u���$)O)n�P1K��>>�L�4�׀D�#�6�|4l̖�ʼ���+��gsX����w�/��5*mM�J��v�]8�˼�Ng[�W�_�������]V����k���yJ�\�{,�M[�s�b������U���M��qc�/xj�߉�K.�#��v�ji̊�t���j��x��1M������塞5��b�_�f���Y��]Q<�)Sl��_��D�[��l|�a3]�%�n ��` ��+��K�͉D�9W�9� �\p�Rr�����9����ɍ<�E��Z'�~Jp7I��ښq���=�M2{w$���[�nf�#���>8B�1_�྅>�`W}Y���v���=��8r������{��L*=�_�<�a����h;�";����鹁d��E���K�����p���ڲ댱��-0�z��M	S��&_[�CN���"=�ù-�
&����.����s�F�j��2������@�R=̲}u t���5�e{��@�$���:Ci�}�J5�*Z��hsST��ޔu@)s�u��\�ڸmu��/�j��Z�o*��
��f����mv����!��2�$ ��JY�9�ʈ}Z�4lK����S��t&�joT\y�{2��BU[�6v�w�>/;r���
_��>> �5��Ϧ=9[�bؾ�u���W��Xl!�[Mj�U$�g�w�`}TW�
Ʒy�Kb�o���[ �;��\���T��V�M�xf	����
���+4!�(�o�\�4i2���"�P#'ydDQ:Z5��@=bV<�����A���(��4/<VNM�~Ɍ�cn�y�yh�rN"��F<ղltS����:#�'T�����d�Ƶ�����n��vx���%�W��-�&��u�e`��:�m3�7�H�h���K�Q6��Z��Т��؅[�!]iA+�A�{Ucٗ+��ʲ��מ̞�h�;�bF\h��c�L���Ot_��kzL�(�Q�;�vl�7��]��x�E�+�l��o�������R�b�W�㖿mT���麪�3R�ĳ�3��<Do���̪~���w�!d?\*��x/���u�66@Ⱦ�9�3"���<c�6ɐ	���p������d�]",i��-b:B�SC*�E4��cz������W8�dX�h��J|��W�N�s��㷓�^��Гܣ�^�ƻwp"6!�@��7��v͜i:'���<�*��������XO��=����|U񳌽�yַqӽ��yȟ�}��|@> >��F���Vvj&:�.Tl,���=����e�̐������ܗݰ},��c`�ښկ��┤N����mq�բ7�i�^�n���@I�"3��M���T7��Kw��(UX��U��M囬�Ca�w�z`hN���m�{ԫ��hs����D�=���N�F{7����Ȕ��e�݇gfr	�:��㴯�:�lSc.�Xƈ���ش�����lI��Ƿ�v i�ա;:�B	H܋�Q�wkE�{���lwqh`�E��}�y�=��� �C���Fo��3	��zfu*h��O�L��F?Tol���|��< v���5�ٷ�c���p;��o&ddQ��9�*_ǅ�y{[W2*�RF=�z|CHJ�H	t5fZ��TKH`wG����D�ԏ���,À�H��d����׮:I�ql:��1i�$�Dqg/�1�Dr�!� V���D�S��|�n�k�l�6�� ��7����prvkZ6�8P���a�r���F�><%�;.b4�X��R�{Z���ǝЭ\�=6���}��S��WUb��r8�5ݧ՗Y\%�-rQ�Z�?� �7��'�͎��lv�=��J�^�R��09���#o���m5C�H=��OQ���q�3� �T�2GM<M3�G��ץ(�8�54���kH��,��˻�cREHrM6Ro`ܷR:�$[�%|�ֻ�8��ӡܶF� Q�rW���)_��$N�6��U9�35ޚW�-��t��igfa�խC� ���6疜��CjR�:���5�2K���\]�md�j�������z(�~������ы;�'��ű��t�G�$�a���3s�	����ò�ި��E������Vj����v�*�ޯt�ζ��N%{���f�C0��KƤ�z���zv������q/�'3{I��Jy1kz����F�q�Jg�Uj��# �����dhħۀ#�_�4�����p�beJ�_4���;?K�:�{Ýr�,_R�~[}F���T�O���]A݊������d��*_�1����	5�dqǶ�\̲.�3�1�#�T�+�2�șۄӽ��iq�x��5Q^�$�g����z:d$;�����ͥ'Vsꗳ�Z׀�0��y��x�o`4O)��=�
��w|[��H2�8��0GN�s��/)�������͞�b��ö@y6��o4�qwM�N"c��$�X�6�]w�J�������$��O�mdg�@ABiJ���f]�{�i�w����9�Bzh15������yFG@�6����5�^�@��(F��z��xy�˥�=��\��4�Q��s^��|.Ǻqo.�`�F�K;��_fV�8:��%K��G'�n}u�s5l��oyC�Cd���/''< Z�]�[�������:YhX��؇H킉�)��}��F���;3Π��b@G�A*�ν{�oV��.%�� �I<U�c�eeT�QYL�S�������Z�&��
'69$eqP+�>��ܺ�Ss�v�f���<�-n�3����=�}�^�UH[X��m��6�F�=S@���R,޵]��k��:��0�R��J
V*�ʊ�VY�]�تb��ֳ����V�a� tҵ�u�k�^ܘe��VN�����5�b��|Od)
�#�
��%�/i�2v�[�/;��s
=��c��K���o;��-�F�%p�cb=�%�9"�6*����f�]ۋN�v���6T1����e7B�-�v��+�T���ִU>u.��mP�hp�F��zKn���ˇr�ƌ9J�k�զCbջ��N"�m�\[6������V�Ua�v	5�i�:���-�9��D�%����g���p�Ǝ����+��(B5׷ݯp��V(qa��F��L���v9��Ū=���$�M�w�;���6�GE��凇�������Q4�+á_�#��ݼ��C{�^\�$ 0�B
�� �`�b�����
�r�cf��1lY�+ُS���B|+GZ�KG�c}+6�aWqc#�b��a�稪k.�.��a���Rv	�F��v=}�2.%�s�2�����Vd�v'����]����%"�7}�ݝ&q�G9��70%�,���)ڢ,.��,ѩёk=��}ڢ�@ѥ�z�,�]��20� .�����gh؅����uf*���W7�d� rf��G-41��T�8�1���u�8ym�������U�q��.%8���q+
:,hhQ�(����-ZF���vo�\��W$a�J���A��u��p�PZ�W���5«u���OLz�[�����b+��mgsR\	���g]�c,LT2C��G�Һ�'�w\�N���Ѝ�A�2�d�\�Ţ�Q��ʰ'ӛݦ�R�rrǙ�ay��+�,�`uN�>9�=����ƃ�x2l;gX��3�w���d�ܺ����a �F��@{�	�;:�k������r�zD�"R�cY�<C*gpokC�6�oMo0���[�R[�@�e�RѰ6�lك�nU�޷
o�U���,�c_1zNhơ��_
�*=�ӧS�l��}jh���p{fN���V�|�<і�v)<ۮ�) � �r��.h^>�#�.�)��i�bja�ռ��w�$&��U�N'Ug$*-��-P��6�׹W�G���^V%�y��4Tz��`�V���TM��S�]b�M�v��)7����r��J�]�K�����{�5Z�,�L=�}�M;o�yB��J�ܧHt&CyW|�U[*
��6��\�o9{�e���a���x1�/U�bY�2J��(MKj	j17��k|��W���j������h��;�gg:�2���k��d��q����X(��q��G����`�Ua�� �̒/͢��:ߔ��%A��j@ؕR06�����<|}}q�|q�ׯ�}x�۶���!D˶�iѦEE��O�=xD�% w�;����}w�����8�>8������n�s@}����W�����{Kϯ]e�Z���.��N�:|c��q�|q�ׯ���뾻�u{���l@e͖�g	�q�'�Vr�E'$rtIΔYaI�I��yۮ+"������g�ݏ5Ĝ�'Y���]������Ʒiru�Da��[7M��C�Y�Z��yڶ��/:���I�tw~,��n�rw-�����v��7{v���7YE$\qtI_[���}n���!��NBu�E!GC��iٻ5GR'n�E�Q����el�|���k�A�D����6BD�b2�!x��lI&d�!����,�):4�F����Z1kF��-ӴOnn���Q�ԥ�qK��t.k�+����A�k�����f�H��������IA.S$8ȩ�-(���K0ƙJDK���09i���Ӑ��Yt"D��LRq�2lڶ�!$AD��H4J��L$�(#e�PF�gH	R
UDB$8>��������OKn��V�%%�W���Y�)9�릒^�WM7fЬ�իKl����Ϯ� ��@V(��F��.�����`�F}ѐ%��xsJ�K2�oV�;�T���RD���^Iݓk����Yw����0�ײ�3)[�m6�u�3j�ę3P�e��Fj)S�����7�r�t�;	��<�y��ő�.�'�Jq��F��ϵ�gq�'O�P뚙��UZ���&�Pr� U*D���'��Ɣ�(}�0���壕�~���u�sv"�fc}�n�J1��V�b�Dk���v�M{��<+5�J�����X��Fr����@�>v���q��Kd!�ؕ#"�����< ���"yTU��;2�V5��hi���ň���=ڧ����*��t�rc[�����;=p�x����#П�\
��5|}!RWj�:ٲ�׭�6[:�q����F>��
�Z��L��D+�^���!gq^L�jGR��砸�~Hw:�gJ9�E���?Q���-J�B����a��ֆl4:�e��3��f4{�ʎ�-�v�c�������֠�)��17vuf�3����&,=ï3=*��2���y.�=m�7�ׯ�<�o7�F��$�C��P�����yO�5��e��4
2�[z�o�9�:�s[�{3��_u���U��.���f��/��t�Š�	z�����v�w*4��n��R4�7F&��Q9�\��A�q\���ԝ�����C�jG��8e�6��+�9o���F��h+ױ��#\����Li+�ܭ�{ag>Od��st��۫�ɨ��N[����	�Sǣv�n�KZ�ϫ�a(K��c�i�֘��j0�G��*�"�N��<;��Bo�0� ߺ���T�{P>�9������fk���D��ȹE ���ݽ��޺�9M��F("}�>pWS�nﳿ{�ff���R"�إ��\�4�|������m���w�7b;�(�2-.ڇc>�F�|�n���9�$曍 ��W���W�b�0w�Y��I��O��d�;+;���uzִt}v���8��vI�ԥ�|�ö�zI��Ҵ�{³p���rA��̂�|~ Q�Ň�5UҐT���T
��.BpY�,5��\�է/	쏝]��*��J<r�.���jxdꃺ֗P���T<�o7��l�����gf9�E/��u��H�p;����z�3|���`z��T�k�pm <YH���1=�'�'J"�x��t[��f�[l��2�;��A�3V�J��jj�[^���	K��R�hP�9-ymV��<@�n�K=����꧟���f�Q�U��BzL�S��[bMTo��9��TTK���X�9��Ph��C5�뽘s�����q�A��z��U����&���P{�R��]�UhN��:5 ᱛ�I�s���R.	����u#�"Dz�s��S��Kn�8��L!I��k�q�|��i)Xn�>	-���r�1Ha������k��oTq��}�?\>��P�
�wHܞU�W+�O��ކfef[deƇ-
su������� $~���j���X��ypa=��uD.�7v�P2e��3��|I���z
��QpP�k�l���oe���N�f���77�B��=�R���R�����^��\�,n�y:�x��Y����4,i^ܪ�s��J��J�<����%�km*�;\Yد�'����y��\���x��m�6�ey�Y�|`���!�q���V�)��[|�ܪ����kkx�4.�U���8#7<�_�
َ��b(h���.��T����������Ǻ�W�]kdu\a��$s�'9�=�19��cg��ѕ�P�+��NP��>�&�~�3�E�cF�\TڎוT�eU���lkh��kv�S�z��w�ˀ��S+�
v	��@��j��#4��	ۜ�{��R���pE�uF�2�3��%�F���cח�t^Z��ٚ�@�c�TnKY
#�YjJ|/TI����.�3��M�ltu���cuϯ��ݫ<�2(Ϻ)��hw@%������7Q�r^{_��a漽T�4#t���� fҐ.i����t��o*�>^��ژ|�n:���W����)W�N����d������Wb��1�l�+\4��e�ՎP��fa��ыz圴��w*���`��B���X��ON50X��D�v���*)h&ʹP�t���f���d��w\n���]�ڮ�Zyj�P�Jv����Fm<�z,.�i�%˧:�ݏw'4(~�x�����7��aG�|S��J�u���ei�Pmvi
N��PH�2n*���H����1�f�jnC�hR����v�TO%JTyS����^#ޖ��n��v�K@V���H����L3���WH�(�g+����g��en��>i�f&��R���5/�-�h0�@Lf�%�<����ǹ��w��cz�u��|�-K�Cにv��HW��=�H�����!����G��V�2�?J3��B7���m��۵_b��������J�Yawm՘�J��\Q~������v�=�0�-r���]�*�r��w�vbH����wWrZQ3 r�雑��3l�:ʭ8�pJ���<!�c1�*��ҧad����3��y���sP��;��y�{(�=Xl�k&�,�؜EIj�e��9�d���O*Jw��эTFb�tWO��8��9ׁue�-���lWˮا(S��!!俅,t�7#8�+7.w[V��p���*;N��d��#4��;rۡx�owZޱ�k��n��|=X #{���'��4�Av]vV`Y����<!��rwdX����71>6�2_Z�6p��e�p<$�L�ޞ>> <;�i}��/�؉cH����/���r+�������5M#cyv�/_ 9��^}��(�4�Uɱ�O�2Z�;k5v��AOOeN��|���Zo}}��A���z���ɤ�8�3iO�����6������CpU�y��h�b!RPR���[��3kQ�)�^�>�G*/"_h�b���-r#��<����oW�d�zUYY�^K.=q���\�U��V� ��O빃� QŌŪ�j�u��S�����\o3O���P߶���*���L+����y�L�ͩ�_,=�l�Ӣ�[�'�Eg���k,(uzV%K���`͆�1�m��z�ڙy�
1�׏�v���
}�=��P&�+�s���C��tejQyNPgj����n�b��H�[1����B�s�ģ�]һ,�E�T��u�Z�n�f��)��|�H%u]���X%~V�c����"�X�q�p߱����w3O�5�h�8j����`T)
8\n��MUʸ��Ӻ��T��vx�=�:nwK�3]���Z���kNQ�D	�fuA��8��롒���1�`����3��ϭy�e����|��/�x0���q����6�7���SKt��dFͻ��m�<��������|�������>�ѕ#cN�zΒ�����^j�K8��)�l�˩��m�H�^n�?jצYORZ&+i	$��j�\�v󫞽�������:`�Ps>�gW��#�P�+��p�gk��4Tw�a����˹�l�N�q�ag�zv��f�^�CvS�m7-�W/s[�h�R������ޚ�}~���]��eO9+ms7k2f��t��������}@����4���'��}v`�x^�3���j�][˄��g�c��7�>c����=����,'��y꧞�hO�TVV\�S�Ln�ݳL��Q�>���v򂽚u���k8Ae�,Q5}�*!����E]�q`$�p�����bM*�ٓ�Oi�-��vKGFE����z�6H�~�`:�,�w�[t�Ҽō=��,�,{�2�m�.�</h<��q��8F�1);�K]�i�p���y49
�}�oo<����2)z�}FE�콙�z:�F]u-�f�h��=��[}���W�� �`�*Un�:%mo�C�\���n��V�R%Uq�f��}۴.Y�k��`��I����H�)�[��]��vx6���JH����WOG3�\��w+����@?�aMw@۞�+���Kp7Z*ob��!�AW���q���K4�W^���]�a[�Ǯ�C�����/p`�L�˺f�wsI�w�,�s|�-,�սB �=ڪT΁������>�x�7x�]����{>��p2HC����Dw��b�/U�ox;��BI$Vl��r��um<R���������ט>�cۈGD�m.����/Hpj$��K��_���6]�i�~��� vv���֦��۲ G��3=.��h$c=�P�e
�E�s��W�j�Ĺ��:���y�̑pon�Ύz�A��L �቟d���pf�ѝ���<?�-+���X��]��k�:���-�����X�s����K��K�f�nG�[tl�.���V����LJ$D�1���k s$#m��msކ�
�",N��v��i��.Ԅ>[��|W����y�u\gd�|�;߽�>> <���j�~�R��!(iR�$5[�rVfnҢ~���H���5��P�u��}aW��6�}�yi��V�ҿKni]�{L<�t6�Q�K	�����BP�M��/Bi�m�����Ҫ��B7@;m��Ĺ��B��I��{k�ը]g�qu-uh�!UqJ|o����-��SOu[|r�2��E�Q�\k���D�]���c}./y����tu��'��!��2:�6v.�vR�~���m2���
�9��w�	ޏb�M�x+y��Ú$�ؓ��e��3^��O���.=2����G$G�ʏx�Q��&vks�F��]vi츴��V�����-��S�����÷�p�$��4���H��:ߦ�sqn���C3������;[Eus�d�2b���#��w>l��,��F�>�gys�O$絤���1�x��{e�5��C���d;�Ǫ�"#+����}���L7[�h�8m��s9�ܬtr����ѓ2��E��n��_:
���Ώ[��x��\��u@W%0�����ea�ŹI-���u��w���b�F�s=[�
�ݖ&e�9���sX|�1�S��w��9��������	�Α*_$wP�m�����1Y¯�*�A����4[�K��ߟ7�2��8��q#r��'��r�q>�;�!�0R�+"E�v��=��ć|���� �?�B0�![���GD"���C9�N�w]�[͹�s�WO��8�����`<+/o䞩�Cǔk�n��N-��3w��03�m�22)�FC8A����X}oM�uj�6�Ԯ�tP�������f�h�y��߶)ύn����.����]�Zޮ����ڄ�*�/��н�5�"e"�݌�(���S��p�kl�<�k�`����a�T&ѩ��z�YڂTr|����q�n^*��cstnV��K��6�U��A�QB:����EX���ؠ�wU~a�2��j�='��W��;UcU��V<���\n�Gt��6��9���b��9�\��wh*��{�$JN����G���U�v�iq���ҡ@�[	�Y�8o�D�An��sN��5twB��ǽuk���Z*	��oI�Iϝ*(F����2��lU!��|�>����sq�e�˖rv�ٺF�t� ]t��|vZ:�
�0�֐E1�A.x���z�
<��\�N���(���4�zhm��]/��=�';̥w�Q�բ��/��6n�ޮ��c�:2��ӹ��v�m"���o(T�6�W��[�c��B:�[̡Ԩ��*IS�zNJ`�O3(��G ��.�읃�.fvK�l?�Ȇ�!��ӓձ3V��Y8�+豘��0Ļ#]<�*wo5-^"ۭ+d�F���V0l�+��}���n:�E� �_]`:B�m�kI�[�>��z�x�ir"��5*���p8�ͭ"����z2t��sR�UAmq�b�6�I�F�%�͵O�KN�Ӓ���o�(�Q�k�0i»<�g:�C2sYW[T�2b3r���¶�F#�Ѳ�J����ۘ���E��8�]��* γu���'��Vu5�.�+4�x�[�I��Vd�Fq�j;C&-�G��;�Ӡ�|ZIb�e�b4[�������D�ecʙMW;;�e��~W�X$;B8��!
�����(���t�X�ڎ�..�·!�x"6�m��M�ھX�v����1V�ecm�c}xON��g�gg;y��]�+d��Y��N��;��*���*ءe�d�  �ǉQ\j>�u��������~��e��`�����Ԯ͖�����{��@�(�z�d��o���S��X�1���]D�vR�N/709Â`$��.�����Yg���Mϻ��*|/��I�wZ���H�3r�9&t��4���Mgٌ��<TL]/�<��O4)7,į�;���3N�)��O�J��|���&V��Bvnx{�oN���I]��[B�3���j}-_����7u�|P,���k+�3�Q}�iK��U�)u�ʰs�<������:�Is*����F.W��,�[G����7*\�3ۓB�D�R�
ER�z.�ź����X���h��d�Ѫ�K.�v�GT�R�����"����j�hTS�r�a��]KkLqU(��|�S�7�/^ea�S�\t��sxQei�׬�Y5[!�@^c7T�wz����b7�/��'���[щ�ѽ���G��6����c�_kf��ݮʱ�7�,��F��� =/���8Ɇ��k����R��wEжM��7q�%��j�B�;q1���!;2�YTHf�Y���)vjgW.�Wt�_���Y�OMCحu%���ɝR�q�}��3�u���%>Kw$��;c,� |�[��ʃpd>� �O�>�
^w�Gw��U�u���w�� ��<||t���8��ׯ_��x�۷n��
F�d.7*O�y�dtQQ(I	��}}t�Ǐ�8�8�ׯ^���۷n�۪��T�#��C����o�u�^����x��ARHD$d��=}}x��x��8�=z�����v��j,���I��˭�	W���E���(���xwfv\GG@v���#�"W�c�"A�"rK㲣�:3���y�tQ�rO�`N��e��`\E�W�}�;6�G'sγ���r!�) ���x]��EW-���s�촓����������ؗ~��B�r���agY�Y���=^��w�k���:mvDVbQ�b��¯��G<��� |�Q�򣖊o-=�_4q��Tʫ�꒺���p��u7��ǝBjj3}wX(Q�h��ק�n�"qE� ���x7�� ��E��ׇ��y���Fg��Q+�DT���Z_���ޅP�8�*$ٗ�T_�/5-vzGu%vܸ�����udf>� j��)���^�cI���0��(�+n��EK���YϒszQ���w�T.�y��ܚ������Aw�̥��tYV�-�*�ݳl̮.�}إ��g�&��ۙ���N�zz��D�u��J�ٻ�B,mA�z��`MV���:����g}�=�,�y�Sq�)��1��{o%��ZV9�s6�����=�{۵]���!�������sv"հ\B���{e��awh�;�6�o6��,vA<���:C_���a�{Qx�3]�s'H�'_��;W��,�o.���Y���\��q�8�`��m7rs�ڲD�}�_a�v �Gd8�d<�4/��{��7�'�cO �Ƴ�(�=���V]XşG�e%��iX�	�¬�C-�H�WY��zu��g�f���_^��|Sܸ�������B_�Ri��q�Ŕ��`ͩ��W7�5ڸpt���F��mZ��̛��u�VL��~���|@> {�}v^�$���GQ��NCݣ^���U����ׯxe\b֚�'vzEL�^j���z 
�[t�kc>�g�^�%/w=B,���,���퍆��\%�0f蓹�uҧ�O_z�sNsq���7av%��Ô	�cºl��D/�m��d^RC�a=��.�B#�]�*����ݫS7���譭N;=�\͚�O\��.�����D	e؈��2£x=�7C�r���{���)\�F���?�!jo[i*��RD�j��݉���j�n���..].b�u���*+�7k�˽�q��d��!s{,���t]�=���
���.��@��[<�F�,�� �t�a�l�M��e��z�;h�q������h0�����C�M$T���m#��j�U��
�<��Y��>��!���]j0PCXf��9S؇3.����xF�ܢ���mϑN����āw����{*w��Ej��TAC*��cO��a
�J15.�7���Օ�͝نug.3(�D�ܺ���Ek�ϱsz΀q���7!�V1�|���W�WxxxU��q���w?sǻ}�\.�V�{��j��X��nT�8W �Ew^���CK��ȸ�}7��ǫ�u��p�ޞ�g��b��Y�sME��=r)S��y�e-�����u�����t��ެ,��o�!��l8 ������)���`�c�j��4;���[��y!��V�1z	�%��n����2�~^>���p�m{o3Qh2O>�(ϱ'�&^�a�|փ�]A��;�GA3�dt�[��<V�.�6Wk�o1�I4D���^J��}v�P�!?���8�zJ{���sj����^Ι�����o��M�{E���,�f��b�ȨF;��Q"�<��N�_���o��R�sIۼ�>���6���ᗪ���m���G���a��i<�j��r�$���ew\�#�}�4v��5	�6�3FI�H��h�E�>&����;�.��>z��T�����a'�뷆�^iS'#݈��[9���K�We����U��5��__J39ڍ�Gh`T������P�s�#��f�Uu��D5ܼ�p�6"GX!��D��]̗��^y��>�-�c����׹�k��}9��K�n��[>�f[�`��:�}<�w^��j�\m�b�Zhfqw�zIVR*�t��tw_Kڐ�p�pX&g���C��KV�&�s��=@��ZK�uW���#r}]���v���ZCie�xf�F�y�-�;˟E^Iݓhݗ��L���a=LL�0�~u]1]�>guw$�@'�1J��s�Tk���7�q1�wK}(l��`U�N<
�9���uG���0���0����r�͠��xe�UZ�~}�ig���:�
��l����ܛ�ˮ�wڼ��$�9�N��3�/ό�t�A��0�nc1}1m�6����%�z.�Oi�xçwfwU��h�ci�h��;>�W������dxK�kv߬��v�X�)�R�0�����͞��fGE=���;�TI;��2P��ͦ����k隥�b˼����6n<I�h�B[µ� ��n.`അ^��cRӣ�y�N��#��}L$cf;S����R�[��Q�z�Y���кk����{"Y�<����`�ϕ�����z��81��*D��6+8E�33$QB�;Rɹ�M���E��ˌ��0*Y�*	W��g��M[�J�J
�[q�bc#������9*�늉s#B
��zY��)�`ֲlA�n�§�cz%�K�Ir�T.�ګm�i��Ӣ�u�:�Q�T)��w��0�۵�x�J\*�>���S�z�E�m���!�J������� 9�5��t2w\����R�D�\;���=p����I�
ؚ��ܹ�Zn�tF��=
�t
�Uer�r��5�:5����
k���'��p�����n�F�ڜ���e,�ٚ�Ȼ�1.�k4�V<�k�Qx�N�:���-��zb
s���um�g5��V>1ٖ��{}�]����� ��Y����^I�E�Iۀ�U^�L�f��zb��e�`��z6r��̄�.GF̖}{�
\;Q�������͍���Mn?�����F�x���]V#��7��(�.���f��}WO
[��W}�u���Rw:q�OE��y��7����><��&��U���>Eһd�.���m��a�a�v�U�뽰����c-��r�a�N��d��}�\hx�x��H:L����L�ol���v�?7
�N�W�F�'���I\v�g8�,��lծ-��g���"�<�H����Fgt������;}�h��=���Cb�=[���{P�37H���fk��Y�"������>����߸M�Y�X�.�p�MUpy��B4�w��쎭�E݅���"�B�x�>1a�O=�87|^<��߳u38��>�m�9ϔT���z��R�.yh=w#��&�S�,r+������
. r���)e���W�����{ʂ��+h����ͪ7c������ws��` ���6C&��`�Bk��K���^�Ԥ��h�7�(�xw��Aǘ�q�H/o��!�Gr��tf.�Ҋ}y�Y�Dbʄ»��s�r�i^�5�ÄB.��Ⱦ����%�XnG{p�A!���8�:��Vb�g41�9�8VM#�-�%]e%�S/�ޤ������� �'o�|�Ye��;_K�������66��1�>����\�p��g_e�x���/��X2/����8)e�A�Q]ѻ<��]z�"����n�{{��џ->=Q����7�������V�|�+`�;�x9�jZ��F�K��C�	�����+���gt��˗5p�����{�Y�!��*�*���%�֐�O��n�^,m4?�����]�\��C�	t�-}��^Xx�J���'$mmM��N��6Q܋/9[�� ����v$ê��w&�j�ٶx�O��f9M6��قxͤ.�A��&u��t��H�U
�t�P�=P�˫/BJj�F-����#gU��j��Y��}mQhط~�;,!�.h_�7���:�'�K����7̃B��䖱YdO����3x�T����m�P}��÷�w�ыx@��)�jEd���<lmu�rL?lss�FA�֯>%s�d��R��g��s�,c�:oŎݡ��J��\1�q����V.����Vʾ����B��ˡaL��j6�}f>���5T�D7��޳%��\y˽�pܛ͑rM9�]^M#�7�y��ood�dN�{T>G�z�����88�4��9Lj6���:���=��T�a>n��#�ܥ��3~�ҕ�RG3b�C��y흾U�v�F��S�'s^�����-����׸�g���aU[\�Z��:�����m�ͱ(�4��v��K��w�CZ���a����=���~�I���|rLө~���}���u�����_�ƞ���L�f�E�����3��ǎigH*����gK=�马���cr�"�C�EV>��`W/#	�U�^�Z_���m,/X@�i6ж���5@t3�������n)��^�.���Y�vҦ�ESx�a�v[4�C��#�&�����`N=e�\0wh����Vw8�;ssx������ 7�������Fdz�L�~����P�ne��]�2�	���*�����kk�Ԋ�Y{��h��-��������",+Z��o�~$-�V���Ed�$qY��7
[)�`(�k@��ڈ��>᧞:5&���uHU�ل��A��WTDiQ^@������β���H��<|���)�Y�����]��b���$��v����do3�����
���`�~���G�9�w4�g�v���sm��Xg��|3��/��g��KO��\��ΛTF�)u�,x�u�̖����c6�c���#�ToWp�Ely�Rk�[��U�zQ"4�@��e�c�ČWGy��eC��#GD
	��ꢼ���Q���cA+�F�NKU���f��;#i�6Y�'�L=Tʳ�V�ԕН�w�jFM�U�s�<w���L�)�K�10�t�]/	��̇���qǚ�c�Q'���uу��cƢj���(6�0�\�UJ���}�#�F�#l�{z=+�#��Q� $Sz�%?ev�܁��auut�D{]�n��	=Y������a#a���(�t�:�֡�l~ج�;a��~k���o��gC*ɧ�.=a��]���	�V0�Π_��1���k�U�g�E���hV��`ڕ�ڐ�ۡ�8���|��h��FX���[m���vK�\��f\ݖ��s9xH@�#b���m#4�����?@�|~?~���o{�w�E�Wǣ�c���ã�#��:�+b��?��\���s��:��\m�
��o7P��v�"���>�h������r���`�r���6)I��m����A'k�w��f��]��}���&='�=��A�e�(�<Q�v��q�IV^�=Ϗ��dQ�m\��&bx4�N��229H�Ӽ{����ʿem��y���������5s�������:�����>u�M׫v�6h��uRD��i��]q�Gvz��RS�x�ok�e$Q��="�7����9H�yH߹�xf���*�z�m�;Xжb��7Ts�9B4���!�R0_C�R�H�닺h��v�b��6��_)J��ё����O}��^�����s�I��/�z]�����C3�c�; Y�rdn�ð�����߸�?���ٵ��G�@@k��
?�����$�(������ʤ㳕����`�1�D#X�T�0D�# X���F�A##�V#�.�\s���*�\s���0Q���# �R2"�#!"�DB! �P"��20D�AX� ��B(�Bc�"�E!�1@�DB!�"�D"@�@!ʡ�X�D" �@B!�@"�"P�A!�"@�AB!�"�1@�@B!ƁJB"D )��B"�D"�`���B"(D 	��B"�D"��$Q��B(D ���B�D ���B*F ��D"!�$B"�D"��B ��W8:E4�D !�B
D"!��B �D"�b!"�5B��!�F� ���B �A"(��H�* A�"���B(�A"���B�A�w`���A
 (� B  A"(��B(�A(T�D� B* A"���B
 A� ��B"݊��*B*B
�BB �a�D")��B�@��D )1�$B"�c�A��$�F��$bF1�d ��%�`��d"�FF1"A���B 1������")T�Dd`�db��,b�*1(�bFF �a(���?���G'��B" F
�"��)$ wB����<�߸?�o�����{��������g�_��=?���%S�?��u�s�>��U C������DE�R �
��h�`| 1g�O�E�4��}��� *���������H��<���?G�����>�D��?�U@b! �`� ��E�$��HE`� b���  �"B B"E` ��@�B"�B ��`�F(�!
2*������H�
)"""��"��i�( " B(�$�����"B
��"���@��("!""!��H@�`� ��*B"(Eb!"!�$ �X E�DH@`� 	b	"(�"X�@�A�$�������������Y�'�@dTI@d�}ÀW��ߏ��	����a���@@h?u���k�O����'��C��6�g���6}�� ���!����_ޞ@DW� ����z~��*"�����DDW�@)��P].��4P@�pW�Ma�Q��X@����~_�� W���U�����?_���k·�����xx4��*����� �������6'���G���?��?/��:��z<�� �*�8A����H�h������L�~�/�:`P};�DQ��C�N}m���
C�'��(+$�k,����xĻ0
 ��d��HS{���V�#l�M��m�%&�)4��
(� ��Q
6�)H[�
1T��*�)J�F�MV��P�*U�KmkU���H�!R�%TH��\�JPJ������U(сQ	E�N���ȗF��L*;,�!�*�V`�RV�֪�m5j҅WZ�y��Y��[�*�mh�UPH��.�5��TR�J�Sf�١���mT�R�+M*R� Am�j5	%Y�DJ�P*�v0���HQ�  ���u��Z����L��cU`:wu�S���N����[w:��N׶�ݻwn�c1]2��8�WT�MS�����:��]�:�M�ηcnT��ݨ��.�*��6�����k�  #�}
(Qv(4(y�À�P�B�
�V�(P�B����{���:��u;���uu����u�v���S��n�u�;��]�J���.�׎�SU�ɫc��v敻+�sm[l)ER�kR���)��  ����V��UҶݶ�]wO�[���eJ�c���к��l�Z��lQ�{oЗl3K���S.ݶ���N�mY�����Z֬�ݴ9uqE*�(��$�J6ԥ�  �w��]�r�����]j���
Wl�o]^���w�IM��n���y�������˨�^�����v�=)T$�%��S�  ���֗`s��t�XU!��TwSF�Σ;b�jپ�{ö[+E`��1���(\��s�mUJ��骢֤K0#I4aBO� �{iW�-�tM7�V��̫R�]���p�6�A�@���,��z����׼u�j�Q]5�7^��  �=��)JE)��U��  �� :X
 `� �ܦ P �U� ���  ��46&  5` :�U� 
@ʤ����^�"�"UAU+�   !� 	�@ w��  �  .ۀ  գ( h�� 1�� ^�G++J�5�  )cFR���**��m���  �� KT�  �p(]w+� �q�  m{8 f� �b`  n�� E�@:�.OZ�)R��^�ڍ6�d���  ��J� �� �.F  ø =����  ���@,�8  =k��Pg��� ��8  ;���	��RF�FA��$����j��&�����D���JJ�=CA� j��OJ�� �$�JDM�T�  3S�~>�G������{w���qV��r�k��곴�Ǘ_��PTI��b��|>�|>}��ߞ���kkZ�~�j����������ֶ����-mk[f�UU����������g���O��3���qoYiꘈ�����)�����1#7'� �����&^i�u7�)qh�Wvn�Ct��.�2��0r�ׁnh4.ؙ�=�3�lm����y�H�7C����52�|����A�Q;��<g���`�	x'n�G�_���C�+K5�a��oN�Nma�U�9I(m�v�ai���e�B���"u&$=�gz8d�xl�,���/Zɇ��"�<��̘э�R�Ҩi�F�"Fea�O(6��̀�Сu(SJ�
�{
���Am�O-\��Y�u��!x�@mJ�^�R1B�ti�c ���^Y�kL܊�BW���tw`��F�[�h���%�	Aɻ���@��(�օSY�+�RX�,^#[y�gEk�'�=s&�?v���!A��7]�l"��8ͣ�]ʶ$z#-\�,h�VQojcr���;�Tv��d����tf��E{E�mH4��A�)DՖ�)[e �eXD�I�J���Ynni�DE����m*�5�l���Г�<�k5n��MA���p�8Mk{s;O�<�6�}�Ճ�rK��L;�1��$��ڼ��A	n��h���{-�E�����TQF��X7eB�.J�^%��L����?�F�sX<_�,�O6�����U4 n
+]��
��	+>tv&/�I���gq�C�g[g��vd�б}�a4/K��X[�r�R�2�p0�^��e'���a�P�9k�L�^�If�uԈ�6�ptC��rqx4��38<�֍V{q�B�2Z�d����h�����D��
���d�>���p�ϸ%oNʺg���7W�97;qL.��kB�X\�&ƥ�
²�,ږ�D�Gv�@��m�2�7����à��������.�s��tj*�5oh<��si;�)�lTҔ^G�X��Pr�ڴeX��J��H�w�P%IVP�`l���R:h��7/[70m쑶Fa�K!cĉ���'��`B���T#yS��_uj��,S��$fm �2�i_b�n�6���.*yB0�FH9t�J�V��@V�F�ڢ�1v1��LCĵ�:�`gC�p-���p�j�"+,��	k��q�ݖ5��t5r#�D��t+h�Ӎж�d��>���kP�%[�:A�A�l-d;�n-�-���n�S�*bW����TP\���ƚ�4#����U�jJ6�;�U5)6lBb�w�Ǎ`Lލ��nZ���t--��y�]$�ܷbmZ��}����*$��:w4�y�!�ڬ�����:�h�ފE�U4�nJ5{�խ�b����e�7Ϧh=�=�_O��Ly��~@�λvby�di�̶.R�ϔz
b�MN��ܰT���T�q�������@����6K�H�3�V��#y.��a��c-4wE'�[�PV�^��ڟ<	Ӻ����4��կuY��ӤR@��8F��溒�՘���
6�㳍���]�FT��:�+-x��c8�ˣ���:]M�6���u����r��J�x��1PLR���&!̬ǎ�S	�ay5�n&��E���0ݢJl���y2���\�H� �8(�������{��CpI��8p3��1�k1\����f� �3/PC*:�[Lb��aű��o`#Dd*ʱ��{��YۗN��yBe�m6�M*m_k)�2��0b�5
�r�7!������v��i�ʋ oV�4�r]�udn:n�B�U�e�P8N����{X�
[��6f�2�E�t�M��� h���I�WwrZ�M�vY�	��#�uw]-�JY�F)`n^��֑����sK�f�=�,��v�R<�r<81S�waO7nk"ƶ�-[w��� n�jFn�,�T�$J�!�++e�A �bwi<u�y��Z���Yh*[f��s�L��5����sm�Q���b;�ac�Hn�f�embPS�t+9���+X����J���IC)�i�0�щ�.�][j��A�k���
���gqj╱^�R�oP���9n�`\� 5�P�`^l��6��i;b�.:���Ҽ ��V����2��P4�`AF���ժd7�.�{��d*�4�dʧwY���01.�K�m$p+ed���l.�{�I;�GG&У�� uc,���<���F�6	e�@m�gC��䶍n��I��-�CI\6Qx[���f�󠺞�z��Xt+Ͳ�u+ i�۠�EJ9t�'r4u�(�Y��M�ѳ��ț��`	^� �t/%��R�4izi4�*�t޺����v�,���"�Fdˇ�����Dp�R��ע�73Z�ى�lB&�iyQ:3b�EZMSW���z�X��X�iS�M�a,�-+�^��n(���K(�L��Ǧek�X;f��K����݂���������q�u�u�i�v����Wha��V�z���0ڷWz�֤�N+#�f��Wso`Ʀ�������2�sU0�NG��9�0-y�f���~����e� ȓ1�7R�ʰ�K�I�	8nẁ�+t�v���c ����W␝��n^賭8�頡��C,E z�֝hn+x�[Ev��X�ɲ�j^d��o,�΋��*$3 �y��;C�ȷ6𴴋��[r�j��|�=+B.�F��=����[�N'D������y�%��)ږ��7Xܰn�Ա7sV+P^:Ln@)
��&���S�E�A���ht��,,�]��ha�Y�ڰ+Jd�����h,'>Z�[r����-^n��]����2��CV�v�=&��&D6�{F�L<� +�V2������|H�
�L/j"�[Y�Tʳ�����Y-�G�R2�[wu�0����B��Z�v��{EMב���G׃4�v&qF�#2v�����c�Bo2%BM�I�&3Wq�f��-bZ�P��du1����4�ma��b�Zv��xE���d�J�@��AB謣[ٛ����'\3���f�
�&���3��2��J�"�I�8mAv1��n��-1�(��?f���&?g��g���ĄLB�[��dd����r��ԓ�z0�m?��1+v����mF�7�[�	tĺ���nn9VM AN��h%[�v�0a��j�*V�n��ƬH�$�t2Rh\�2����½J��ӈ����y�i��<@���]-�)]��,j��i���4#Z( ]b����Z4�&Bj���J�\���{H��6����"͹�3u�K	���.�=��3 ^�SYZ�iƢ��x�Y{��,M6�T�j.��{�q���f��׷b�dL�jr�J���pm���$ۺx��B�m�C˘�Z�[2�漐��p�ӬW�����oF�0���f��,*.�A��"s�B�����Ǌ��FhTX��x+ց���[�u�;�����>��7'k�W�h�>\����t6fv<8M��N H�mb��G^�(&2aT2��)-�2��Ѷѯ�nM�]Y�\�����!�1nl�Aa	cW�k�;����׺a��j��-��i*;Y��a�MMY��������6�6�Gt��g�5����x��V,�Yr4a� ��IV�jF�lf���x��N�ԝa��SNJ�:1����:m�z%[/E�N�M�����aY�����1����ě�պPf�mK[&���I��M&�Y��f�?�F������y���Nh_jˡI�!�$�63"U,*���vNB�-4�
@ا��Ҷ��d�T�:Qv�M�$v
E�gT�х�F��蓧V��;���~ai:�x��I1��	vܲ�P�b�Ѐ�SBR�h��5n���JG(� �k�=����!f,�e
:4kF��*9J3(���kP�d��"zm,7�S�+���`�+D���t�R�0a��0^U��]:׵�a�c
�n�ȭ��)d*H��~��e�`�`с:V��V�o�Eu��`i���b�e8���E�7db%2��%v��G��W��1�R;���ԥd�Yg(�ϔ�3������a&!S粞3��P#n'J�H)��LV�
����ڏ%�a��e�֭0i����k!<a�Q8�T��z����M�D�4�^����W�����f�n�HVe+��Qal$�J��m��`�rQ_+�k(*�u�+.[i#��^�S2��ք��٭��.f2���E\tm���.'�KV�mp|>�*�z�a���m(3a��nؽ�s �L���?�嫢���e��;N4�jZ�p/�#���%�(�wfV�<����b(�j�n^m�:��K�kX��n���x\GV-b9���QM�GI،�7��n�]F����^L�KA^2��j\y�4�f�m��<�4K�pc�P:���j(�����n	��1�0�9�
b�܏l��>�Cv�1B�t���h�ȸ�zBKt#�!�U��軥w�a.�i.�L���i�Uv�#rG>n��ѽ��dRּ��l1�6���.F�n��,)[�4�p ���m�� �����[J�զH�"�%JZ�Պ�m?��ڃ7�-���|���ld�t�ϱ:� �܌�[*U]cݗ�Ӭ����Jf;��)�j*A�;�����o��0t>#DFO����{��n���
�h!���S��1��zt^TT�7O61�$�%��2+CZ��g�;f�%��b�+mŗ��V��ƨ�Er9�q�En��#MBh6]��ac�1�66dU&6�
èe�1eа
t��fV��x2�o���'G���f,
ܓZmL�,O�5{`5/k!XF��bH��u3Q{�th�8��,��p4B�\��KBҡDa�C�|�t�c��D�7yM�[��-��@��]Z"cܽ�L��R��U6����mb�*nc�f�Ա�f����=����/y��k+>�0�U5�s�,]�4�ݍ�"��$u��dr���4��Y���14RU���/���`���:��4�!�Y4��P�t����e�sCg҆��4�]fS�"�z���E$��Z(R(
8��V*�5����zH���I��tMiV�R���+J	�-hef<)�Ͷl1�Lӂ�^�C(* �,�7��7N����eŧV+�&v1f`&KںG�����Q�m�����;�J�B)K]�NT��dˈ�N�>7r�⽩#f��7`�@\��h�����D^5D'�aԪm�)�ia�U�c����G�Cx��.DL��Wr`hэ�f�kld��(����F6�Bm�XF�xf�OQ.D�p|7!���v��yI�c tr崲����R� [Fh'��v�\�R������I�d��G�6ð.�k�j���4�&�+~1f����,Jď#W��@뱑!���9��bjͷ�탠�l�D�>�Zh=V�m��g]Cw.Ӑ�ay[���$�N��AVm�W�ҫU��I0*���TOF2-�ZvZ�ś���;�����#��䡚shZ��4��i�{ݹ"�k����*f�v�)ЮҩaEc�0�J��h�KX��P�)GlO&|�Ҡ+D��.���1p+����4g�. �'���8Sa���
�-[��5�QC&fǙP&5!�JTq;�0�b-ۥY��)�6i�C�Ön�[�9B�ՠ�o �Z?(Pɜ<s휓����vI鏟(t��KSSJ�!j�z6�Kj��KM�P�˹��
�,SkE�m��iWE*gn^l�~�˧��[�zg*Z�aZ��<�H���Y'�T�Ȳ�X)�m�o.ທe#�LE"^�vFJ9�a��N�x���`�UЩ��0���	VA���\��u�_��Z�v��lIF��-��v��$�tC���f�l�ХL�����y�b��-���[�f�֝�q�R�ɏ���{����z��g5�1����|���O+4x��(�d�2�b$��",�����ooZ�J
]HŨ�S�ͨ�k�Uk�3(���S5��٠���j�ؚ�VⶴS#)JүV��,��T�	]^& ٭�v欁@َj44'�[*챒e�[L�1Y �{�;�v\�H5J�v���(�\r��֤{�oY�bD.�J+I��X틤
�� P�(�"���ֻ���0K���A'5�w���YN�.;�R�%3,�(��Z�� D4֛6.�"0`ѡ�6Ykt�&ڃ��7���r���)��In�b�h�Z����'l���SuE+��)E���v��ۼ�aǄ�LtYA��r]�7뻧�I��n�T��!�Y�-�ɫb���x6�Av�˰�� �"�b즕�8[@;�0��i��B�̬�d�f�B񣩄F����X���jn*�엷�X��:���:�N�M��.�L�i�p'�TYov"
�8M�{ �iم�-A����w�h,��b\ۺZ6
�{��;�A��MZ�F�:e��� 4_�hTD�̲j2�݊b��/Y�ct�\�2�nfc���N���""#��4�X `��sP��G�Q���G+5��'n�2nmb
��)�N:�t��T�CS`0�u+NT'6�;�dVŉZ�OeG$�Ǜ�P:�а���;�6��P;[a�Y �yʽx��Y�6T��2S����g�V7z��cm�B�a��l�;��$��[��/&�K�y,�$)Y6>9i�ɢ^]�6��mB�m��ww��,�ŏ���G�V�2���/���;OO'}�/7�m(�N�����$��l�x͙8"3�۝��FCǐ��{��u���f�e�Υ..�F�.bz�a\�:Ggn<(N!��w����V��B�'}��{w�z��Q�EJ���'�{�x�j+ٖ�p=�b�e`����}�QW��)���@����ɼ����S����w��nt��=���a۽�}������a�Am
j�ݺt��c�OwZ0�϶ʇ����=�.��!�^�� �OA��-ħ<�����`�=j�4'.�T��Y�ŗ��͙Cy�4�13-k�s�Kun���k헙)	�V�s�·#.nw��:��.6@�9kZ��=�x���b�Yϡ�xM��$��];��)�
��H��.��ԳK���2K�pНVE#�^�}��Wt��U���$�9W0��"pq �����sm�e�o��N�%�e_ U���{�����,]����ݾ��Pb����sHՌw�1GgJ;ot�b�kk\�����lc`\�m��l��vg=��=^��KIyU���A���N�x<� (��m]֩��[-m�ǵݷ�j{�,��i�R��>C��x�1�ܭ`�Q0���˘tR��t]�Ե]��������z^s�����]h��:�[,���Uƚ��T|QW���|�&oD�`�1C��+T�aq���p�	uwU��>��{ћ��5�$�{|�qF���M�
��M3�8֞����n7
����#�V]mZ�Q�1R�{)i���6T��泟>���P)�oMܰYr�����\ʖ�Ɗ]��8],rgl]��K�b�َ���*�J�*�
��з�r ��p:���TzmfP��L�tD�T����"�k�Kf�r%V�T�������j���hM�l{�)���2�ӫ�=�>ܬ=abjԾe;f��hD++R�����'(���]�wt�@�l>WJ6M�o�k�	NC�9�F��;5��^q�|��S�=F9}m�uQ��{S�R��J�ʛ"�״z��ܜkw7)�޾ܴ���ḯbC3���0Aͳ�he�!_F�q2��,tU��Ÿ���DQSzQ�����Fe_�����Gժ�K�+y(��.��*�Ҩ���b��=��qLb�-�N��J $�! k���C���y�q-��ˆ�h/�,u�6�`f�Lܛk Yk����%`��d莅���x[e���F�8���l���h��(���Ծ`ro)i��t7սB��;��w���:3���Bk4c,����v�z�oAd�Z�(Mچ���g-qR�6)��e6Q���u��`�	��Ў�j6���s��:\�[��u�YKt�P�.C����bc@މ�k���uaE���*J8���9�ݎ���v�uA�go��P��Z�i��ok�z�#�pZ���{g��seZ����(S��v����v�rV�U+fu�,� �f%��������Ȋt���=�0�<v�ثȸ]rF��P��\o�T�n^��ket���*죐\�{Ƚ��n_i�t3I�R�X���'ʶ6�F)��Zw�;{r�گ�Y�kuIm�:����̗����4�]�vF��,T�B��\�؏�q��Ev��}�N�6���%�xﴍ��7�{�Jsy�C�k�g5n�@�z/�b%��a�8��.%�Vl�of*:zW���ߥj���T�اG%/����_!�_u�i�Մ
�z*���R3U� ��4���(�u��jr�������U+M�6�����.�Y�V���5��'t�l\ݶ�˲N�m��y�6f����3dٜp��k8N��k ��Vj��(�ɺ��f�Q��fP���m�7)`�d�G/��K�T��t��X.�UjP�;��5��8�}�k����d��ׯ���������Gpj��>.��쳝Iá=�ϵ�WP���C%܃��u:�lʀ�R�hb�W��<�kzJ̃�k�V��ͅ����v���ƹ�����I�6��HWV��i���{z��p:�cB븫���'�sMj�iy���Y,`1Pӡ!�]p���f��jE8i˾��
�Ѫ��EP��_�;����t��e��ݝ��u�er⻰�F�]�s��V���Qz���>aÐ��Q�`6{�뻂��A��u�G���$��{;��xV�rr�=R�e�v1�EF���z�F�������,9ݡ��/���W�$*1M8G>���2����˗�N�m�f�����]�M�6	F�g���1��y'}�L[/w{��ķ�VP��:�0����}�[;�6T�eSN%�y�E�ټV;ǽv�\��A�=�O���y^Q��|	�4k�VW[x�X6�X6���`��Fki�cYw*�s}?��˩�g�?X�XBǳv�V�85\���7y�<--��=v�E���ٷ�+�A� ��~�s7(+[Qn1j)�Y��v�R�9�>�袇[��C{�4$�#(ͷzh�r�n������4��B,�)0ж�Ў�Y�N��z�Q0à�v�=�{U&l�*
)����o�L�w������+��詀�]�����X���W�ؗ�%�V1��7n.�0vs��JȦt4�E]p�䱥8��%�e�n�53n����Ā���<wzj�`�U(;�0P����w�ٗ��TѴ��KW��M�e���H�����J�'��v�{LT�a�Æ�.H>�)Xz_+G[��.�m&9ҭCJ�1���-y{R٦��q����!�po"�]�2�r6M�fZWvjk�໱�ۜ������N:3b��uolb���]W�7�E��	P�Y���V!8�;�ܙ\&^����S�qtn�pnN4�g6 l�,����̬mev�ʹX9�ۊ�ze�qכ$�)}���5�F���بJ��Sum�=|��Mu3k� kl�[��!6��ٜ�J,=Ǉ\\-�ۤs�u��J_f�V�w+�63.eL���7���:���Җ�u�9�)���A�/�b�U�w�Ď��UA���N���X'Σ�Ԅ�v�u���6e�;�x�o��zcsm����e����Ra��v��Ws�t�{��<h�"�݊��2�D/�gyr̜#�u��tb\jI���ۭ=ź�E/�@4)�Y��)D��A���)	۶B���T���{*�e�=��v�rk
Д&�b���\��쾽�C{����i�r_"��I��j�ѽ�5���/W)S>Y���v�l��f�gO{|����:Զ�8�R�s�U1l��/"�7Z�csb�3�>��j|wb�\m���[A�;��h���+�
��`�pV\�˰ݡme5��;�y&(�.��A{+;sM;����麺׳�=,�7R�o
�"�`�S� 3{�_D�c�0%JsaH^��5maKk�}K�Z������W��m[��lI�;t�*͟Y�̏��C3&8�
���#�WC���Gpݵ5(M�����\+{���2��0�#��=���W�@�[��y��5���#M��Jb>}���-����d��)c�u��p��N�m���|�I��󔷑ٝ'���ފgk�9�N����dݩƙ�Y����.yC�w�������VcvYE��I.���+�������i��r�r��o�]e�F��7�m���Ө)���ͭ�Ӯ�X�5u�Tf��P���J͚*��8k�������z�kVJ644�7����%���uLY�Ʈ���WEJ�R#\����u�h�8T�s���$o��x��[�� �˘Bj�}����Y��=�5'�}lEr�ħ�b6��b�^�h�<n�僬�����B==5���ռ1�oq��Dov9;� �����Y`�xU�YV��|��'/�4�q;���wܞ![OGuk�KFwMm !�r�<T�����K1�P��b�B����(�M4v���{���U[ ���Voi�!+�w�������ǙBhu�<quI[�kV�z���ZuP|��̽ǐ4h��/CqDw�Tb��K����f������y�-� ��K�,v��lh}�K77L`z�U�Wfh���i�+�`\��ݥ����j��J���\ՌLwvWG��QجӁ�8�z{b�YIe�p�N��2 {�_Ctq�T����q�3
�]�����R�Y�P6v�AY�RŁ!� Λ`&KA,�P5�53{N@Ջk�h���c�'�f��'���X�XF��{-44�:�S�k�}vh�m7N�^���������i�[Llʴ^��5�v|w��p���TXC��\�ȃ,���2�G�;đ�"�%�͕���={�p�6�S��F'ۖ�wb��U��J$s�A���V`o��R�Љ_d�j6�=��`F�zx��*�ޗ-�5�=˷��q�v�oMV��֛�`��yk���FE�ӆ�dV�G*���c%�T�yY��q)�[ mp�,��8����	Қ�9��[���"&üg��8'���|��;�&����?B�:յ� }J'�6K<��Q^Gf`��^�ϰ�l����	n��ڪ�h�B��n�s��)X�������npE��PR��^�ا�8�`�喗���{��������a��bnX!�0}}+;4I�3E'G9{
�0`ۋ#���y���Ԃ��ONgQ�[����1�ʻ`�٫	'KEH#ł��>k���ޮ\v�d�Lh�{Nf7|�q.�lḓ�:.X��g4�E����Z�z;b��[j��_��)cTL���3�8s�i�T��b1�R���˱F������e2LT�Z�����*]����w�E�^l�E	|�}y�Z��
j���ws^bќ�O�3-�7˶э,�����M��&ʻf!!�s�>΀�n�
���Mb�=���;p2ӗ�k�\+9�wXB5ι�j�D������Hc�q�jLu9s�ؔY0A�N;:�j8�	��	|�F�"�W�I�ĭgm��v�37B2���$Ӓ�×�f���2�Ȭr��[\Ɂ���'�<��~���9�U�V����VC-K�I]cM��S���֍���ξȄ��Ǆ7�M���	�[���*fA�xW>}����\BTOX��͞�<�*y���Pa5Yw���p��7�P�ܖ�۩sX;���Ky�hص�VL�:��N�p怍�)B��e�q�wܸ	��̼1J���`�C�ϖPɵ�b�/���Ի1^��vL�W�ET��/��{�H�f8̚��Y��6�9ε)4��j���Ū��k;9��v:��D�	k8]���3�z5c�����2��u���K���|�*�W�v+��7�Ck�.��0�^{��@�#���CX���{�/Yx0��/`�Rm�>�y]+kQ�՘E:�\�ѧPi�We�X��L��f��� �ڳ[Fv��r���C�Ms1�x tc낝�AH�k}��Z���<lt]����]�L��ޮG0�0�GW�: l.��2� $�74r��tn�V�Bj<�[X�S�i�V�
�V,-�4�dՒk��nt&�]�ÎWVP�\�������ҵ^��z�^_n_h��_=���;�m֫9i�����n\�I+�������\�'�m�T��1��H}��P\��V�X��@o��pjn�9��g*�-�%��V�H�ZS�gw�Wt���1��+��K���l��ywV�8��d�BN\.i�{Q��D���]���.�R��s�C=���O������=C�M�+`���L�FMI0c��Z����
r�|i�Z�G,	ժX�y֢�З{��
�X�� Um��o�MQ�����^c{.s۔`��N�w������
����a�(���f����/��uh����j}IӼ�7x5�{�v��GWhHӹz�����yf�Y[Ȇ��}��u�H�,	�;��J��wJ`�{Z+hl�T��\P� �j�����aV�;H�������˧��x-���^�f���X9�s�`�{B&�q-�q�7q=ݽ�CN�R*P��gEZ{�>��;��0�Ȼ�4֮Ӊg]@��dt�r���[Z���,@�_.���P���&q�xx5���(^>����nJj�����]�#ʍ͔z�Hc��
�\8$ޥ��.���R=�R�#9��7v:ſ 5ǂ��9�6��<w9��=�g/XE��C���������m	�0B{��+����b.��o��]^�VA�-N�R����5,��k>�%.��'n�����QH��-���
7f��Q����8r��l���)vf�T��d���k��1IRa�b�Op��L���k�Z=�\.�p�-��P�D���W�;sB���N�|zeNsՑ����Y'�R�n30� m�@���R;K�܌�*�ƛ�-]jO��֋�N�fG���i�;=0v��]�SPwf�bCIɕ����k^�d��;��Z<�F��9�We�p��I��v3�Z-zG��Sj�ϨU��+�f`Ȇ?��������Z�wd.[���Y���&���)�5�u�ژ̤�"�uaΥ'/���\q���"�V�|���Q*�9U�=7vBA.��Z��qJLV��v�����-kJ}ؓ��.��es�<��Ȅ�����s�Nb�J�]�����V�$u�G%���Qα�����_4�o7k��ړVVXwx�r�ڬ79��R<mM�)|u��BH�k;_!֭#e�cw�Вo�8����m�8�/6l̜6�����2vM�Ԙ�`��|u+�ʳ�X{�f����.����*p���Jt�x�}a9M�<��Zqu��ӯ;��������KmUV�����km������ߣ�ႭQ��-
z�Z��ּ��挤��2�7l�eUe����=19jl���z�8�$f^}n]����*8~�t�jke�L��k���i��L]3ޯ��~�7�s篇 ���`�aF`�z@�<F ���ӭ�N,IC����_#�5q0��p�][��#fY�p��BKZ�g+E�W���<LeJ�h��ޜ�P��I䱮�q�E4�f)˰�e��*f̼R[���x%r�n��լ�^r��t��w;v�l] �Nٗv�/��sRw�)n�@���
����
@j�&���s��ThW<Ы0��̈́3��;Hs'|c�B34��
��W�p?{r�#��b�$�|�㧍٢=o�Ӣ��"t��tnoU�7�V�QWg*�I��lD�3V��qM���.�˺ګ<ݎ�ut������K#�u+O��͚�[���=7= �����p�V�^�O~�
���̝K�h�Li��@�]mIϓ����a�ڥ-����4��`�]gw�͒�G���ʷ_.c1\��ͬ��V6%����J=HQ�[�Gm��eˏW����w&Mgsҩ�`�N"�̻s:�ʦ�:�##�2Ϊ��Cr҆�����T��2v9��iXsnXᲯ��B;��i����=ۖk�'�;����&�E����g|o��� ��f�f�w�ID��'/���6j�Z+
��nR�jRT�����CCa�+�����Ȟ�l�.�(����Zs9�#�Y�/i�Uݕ��?m��i��7�sec��8��U���8.�y���6�]Ƿ��W9��)%Y��Ǳ���lm����O�K>x��e;�%i�8�R�JS�R �6�d�N|��u*����]O�݂o;��H)�s?X耀ķ��7|�0��=,ի���=�MI�ʳ�3]�g� �1�sl�>��=:�x���#�;��d�ƧdG*�]��Җ7Ore+�A�MhwL��m�j8�:�af�K:5����R]�t
�$�Ļ������H��=e��V�񁇯:���X'4�˱�7x�(�̴��r],�r>���>���W�����]X�js��`��E�,LJ����a��4ˮe�J���0��Z�ՙ�KFq���$v��ݩ��h�܏Ǘ\��Rڲ�:����]Z0^�]E�u���F-.��	�n�V`篧��1�)����KK����ެ5wU�'�k9n�Q$mi,�)m�nWK�v�)ԨD�\G>�Xj���v��Ysw���$���p�8B���2�ŗ'���c��RBd�,d��ߔ'��Ќ���[�f:��՘��kdS�$��]�:W׀��D����|k���Dl݊ve 1.�l���9@�w�`��wZF:ܰ�ʃ��_Dզ�j��i�<]g���-Qme,��:�+�EW�j��u�Γ8�$ wWש�P�k4s�r��Ae��[W2��+-g ��Շ��6��8�r�b�n�A	ڬ���ZLy������؜}0v��X��V�ts2����b�^tsS��If�I��;�v�tn�J�m��¾
�φ�]Y_K���k\]0���k�����P�����Y #��\�jpܗ,h�h��9��i���Hbh�w{V�:NmĺSt/�hK��4����E�A�aR\�s��z�}J��ua�['��;�	��Y޾yo5�ܽaF:�R<9�h��l���TR���7M�2c4�L�iǶ��|%U7�+�p�T��"ʷ�Q/�i}`�Y89�L�}ӹ�}ף8a%���rWR�q0�H�L�ZNt�z�)*׋�����U%r���B˨��{˃���]�E��L
�)Y {��{�lEz4'ADn�Rv4B1I�MTu���VL�N�56��Vk�x������셲��7��֛2M��Yi[A���]3(R�_R�K/O=���e���.�����K�s��l��[s������e���9�}�0l��ܱ,�wJ!�0�,�����[�Ni�R��zQr3���V�v���,.]�`s���d��#1�4b�4s�86��n����������P���ṓzJw���\r��s�Skt	 |:�E�R&�:��+ى��{��x����!�חF�؎fWJy��ʴ�\�`�HR���ܛԾ+����&�oԷ�]� ��5��ir�H����1Zw���9o9b�7���t^M��w�yj�j骷{i��o] �]@u�]5���+U��C�
PAd<=�m�Wh(��v"��n��Z�_,��B��#��{p��-�F�ؖ/�g���MW�u�V�m�܋��&�d���[�a�n�6�D=X�k���|�u�tn��A��u���U��˼ǅ�����m��y��k��A*�J�ͦm���b�t�Ш�P� �#%'t��.�&&�e����袽��`ûK[��龔�M�W�QB�u����~;��I���,����������Z��U�#W=�������6��Ԗ��&|�|;Vq��P*�i�0��5;�EwM
�fiَ�1tn���NǪ��p7^�r*n�B�Z��㴤�|��NPUoyXhu�-Q|;:�\!*�6v���{"]yd�ے�g%k)$�qc��h�!t����6�],�����=y	�g	:]+�4Eչz8����8b�T�\ �U{�x1z�{��8>(SW�,l�N��{r>�{�Gz�/�%��R3�,^:D����]�L�4.����`T�i	 xd�[�7����?�ц7Z�N60�Ҡf!����.�Q���*��L�f�.��L	�P+۴2��+k�t.(�lo�];jIDj6��]0fs��r��[�f�u���^�s����l�sv((��S��9��[׌�R��n��2�=�G��5�`�/u���oKV&LC�W>v��[�Ʈ+���+��sj�]�⒡E���Q�8M�6����7L�]5$w9L/!��X(DVs���3V��cZV]�):yd@ɭ΀��	������]E;�Jg�u!ڸ���(�ۥ���\�>m�n�N�o���!"�N!�#�ѭqp�������r�_*��F�c�,}�QO:v��2=�\`FM��#6�M[�8�#zr���d2�������5��mv��n[���sTp�#!����{r�K.�u�"c�ȭ��6����q�9n�}�ei�t��zsmW3��fr�=��e���s-\������]�s��Z�x-s�={G]Z���	�R�]=Z,zm�r���(�!{�}�աэ���.�5
$��+����1�� 5�r�XZ�mT��L�%ep\޺�Z��V��|����4���.�=Y+g$���xi��8l�*�Sc�~�T���[zv�܂.́��.Z�6��u��7ȹ�0�d�������d���H�4JoF�]���9�����;�ޓl��o>����ݩ6��iu�n�g�i��L��K�5d�s&cֹЛ}��\9�w0J�ݑ.�.N�d��o�k6�6�/0�C1kE�U�7se��3ˇLsV▆#Sb���wmNr)���$c�F�K����Iۣ��ǵp3�X������NT�)f+�8��,���<鹣`;q�J}�,���:��5i�i9�o�;D����N��P�*XP�0���.E��s�d�29��J��	v�[A�Rrz�p�������%���k�]�Vu]frv֨�֕Vm �0*��"�6*��+:��d��X�7�z]
���b�T���F�W��I���(�	�ݣ����Sp�5kfFe��d�U[��7��e��V4��@�	��x�q�#uL����ƥ�G.�g��R��x��*�Uԯf| 2ئ3e4^R��a�
<ud��7a��]�ŎV>O~��ɟj��f���CL_2Y7*ckF��ܚ5�6t����,��@��[9�&P�N`ȇW�-���r9�J�>�ts�>�xA�w<�1d�pQ��)$��u��Z2bu�˹�8W\g*�۸Ua���b���tr�۷����WK���a��ն�N#8m�m�s��B�]孀1����iɴ䋖�uu5O��}�m`�k�[�P0����]Ϲ� �u��je�ʐ+��t�Z�TU�f��˺�q�WgXt�ԋ�Nͫ�ޙ]���(;-͠���Sp���A3O>e]�[;�r��T��5�=ڽ�̃�0�Sq������"�Ww�@VF2�˨�r�@r5xL����[C]YP��Q��妝^s(�Y�ڭU�������릺����2��f�٘�V�=��[���}�L��1����Ǐ~ub�o-{���pN+�,��Q%�嬃�� �{��}�Px�otξIy1i�2@�sШ͕k�[y*!0U�D����/�u��BWj��D3��F�E�f�cle;Ƿ�Vi}�lYڻ�>u�L�C��v����F���V`��!d�͹r�m�t�T�&7s<����K��b|=C-�L��t���ޗ�n��e'R�)��H�蔆";.��V�Gt¶H���ӻ�v�۠P�R[�T�p�q�6^��W(�q���-���xʷ|��6.2��y#ܺ�a�7��:c�WK���\V�]��S���z��d��kR�A}cۇ��U�3Io8w��݊�]H֎NQ{�r���q|�U��i���[VRc�Y�u����q���}�ЉL�|DS]r��U�j¬�A����&�O�	&�f��Յ��d����oG9	��n�5o�k��e[�ܽرt��ͬT�Ք�����D��<��Vg7�L��k�gX��|�+�*ֳG��M�.�tֶ�Lb��%�w0�.�x���Λ.b$�XA�;w���k�ᰌ�pTE�O��!;�"�ۓ����ZܮY3Q|��
�{n���H])�X�v�Ud�`�4��nŗ�\|�wt�Э(:�9�y����S1�:�+P�Kwr��K>Fu��dAa�C�ic�Ŭ��7��;5�`T���HD7������#Yc�τ2�4P�'�Mv+������H�8�$`{Z:(L�|pK�"�7�i	����:��,]��F��ky�'+,�ٚ鵛�ҝ��拮)���D&��U���H�3�c�/��=ۛ��eks����M���@A�7(�[�3n�h�6^Ĥ
�_q4�]�]i|y����Ӌ�¬��l�r�����T�:U�`J׹��/F[��y�Y��J��:�s��:5�w�$�嬕Yԝ��%$yv�W�#%F�`�C��n�k4X�Ƿ���d\���R���Ů�:����(OcO:�H�pJg��vf����e������E�ȌCCf�t>��W�*5,�=��	�Ы�7���g����O9jyz�%�����j����u@�Ժu����
�ۍi�0� Z+4���f�G|w���f�m��r��UɅ�<�5�mM�r�o��h༥�,�+�;D���V�̤�k�o�u�E�b��gGu�=|��v�1:���< 6l@o�]ܝ5.�z�����ڷi�Y�U�LM,���i��נ�ܧP$�|�D����r
�T+M�Ř�f�Rs��D��㣬�k�q�r*�� qF�R�ӓ�­d���-ݻϝp�@��!�ݻ	ކ�#[�9��1}�aT�q7Z����'Qt�,��;%:nR�.���km���+X]r��u�D:�5}C`���.F;s:��E���-TT��S>��<��{�}�R����z���^��m�,v�i�Ğ\�*岶�foE��z��c��rug;5�6���XD�h�O����Fp�TӳKW]���ȥw{��طa_GS�9��Ƥ�R���>tM�xl�d�ٛVQ��'"�0J��tڢy`w��1�vf��q,�����Sf�����n�6sX�b��]w*�ϲ��6��k�/zQ�6go#��kF����	�g�7ӆt�A�I_\����ڽT#˸��.���.ۑ�ht]�*�\M����6�Rv��oxu��PY��KN#�1ӌ#�9�
$���WM���9��4u�9O*��:H!��[Q���q�BC���S�(�*�uӬojհx��&2��;s�ra�+���6�\;oz�jq�աy�����˳;������N��Ӳ�ӥ��y>(a\��������=H�������چ���j��.�'U���*�ʘ��Y�eA���$2C&i#N����/���b2�7��M��9��7C	��`g]u�,5Y��(���I�vI�
�5ZffPIZ���aX+�0���a��$��C���F���j�h�F�>,;���5�ٵ�dcξ���'ø�ԫ�U�ou���o;u6ʅn���m�G0��ʹM�@�A�<> ��t���b� 
���{�e�&�v+T��e<�]7,RWEl6�����k�K[ȉ�i�v�8�g"݊Z��}NZ�C���k/t��x�\r��I�A�lZw��i��Cf�]�m�TE�D�0�e<�%�[tWM�D�Mn�����p|�Nӓw0�� u�b���
�4��]�Qk��7f	b��X:[��n��8��`R�.ܷ����JL�ӆ��7dCPQ8���>R��Kf�"���ns�+z��Cme�ŧ7uwv��h�h��p��7/o4u嬥`$���;�ofwK�l��j������;���"�T']C�r
;5�O�:�h�-s�W�9ml�!�Ǚ�-��Vr�b!X@�����2��3�@�����$�guɝ4Eum�ԉ��
�\+2q���Z�9�E�~��WnP��v��_W����`�����ۯ[x�1{�_���[��cv�j*�{}�z���Ziˀ�/���ܹ]���>cZ�+���1���H��X�vui뚐��6-�̆a#��%ݶ2���\i|'+���ƭ��b��w��o2��Yi�z���K��߉
}���Q�u���Kf��Ɨg.�	w(*Uh��l�ԠET�ϴ��sgI������( �����u�[���/��p/4R��DVg9&�\�.Ƈ�s����B�wI[�����Z���N�"��o��hV�o�Zٽ$��:��LI&��k�4�D����:��%��@+5����/�޻cx�;1���p@K(��s8�s��eۧ@ݦ�M�FV���Y}��uVT[Cu�
y�0��@�\�nK.vg��yXaY>h����}ÅM��c˶��ɍ7��f	���[��"�<��;j�%����� �]m���YMfپ㗈r�޴���6���C�Ξ&B+H��$���U�[��p�1GO�P�ł��9@ٕ�#ݰ�vVe�),�T>�ywR;
�R��h
ڌQΕ8���C\��˺���)m�u'mH60^n�w��֡���8��9��g(�]v�'*��zEX�[�C����e��ZVx5��*��ut���#��`%��gv�;46�%�rg6)��p��#3gv�#s���$+�Q�\��˕�Y�T �h
�P
���ld�	)�(�1!���s���,������ۡ���$��&R]�C"Q� Ad��(ɂ�;��e�&���aLe(��M�t9����1J���b2&$f�L ��d��l�L�E)�"�����t ���e�P�;�ؤN���Ҁgv�i�̀n]��u��v��@�6I��hT�$� ��22b��捤Ƞ��
$��5�$Ę"�Ƞ˺���wI�2�Iw]Wwc&e��@đ�EEH4fX�Z#A���K6�ɠH�2Ť�I���5�IQc!˙9��߾w�����＿�����p�O���n;i���n���CJ���Y-���]�vKġ@:oyh�-α���k
X9<�IM��*<i�X1>�ֳ@]��T�c�P�_��E+ιSwZ�����Y|6Y��o�\�ۮ�
���{A�H�O��Q�#����Ֆq���ea����+n�x����²3��7�{ܨ&�0�6�U�LZPW�h����K���k��&[]�u2��V7!�x�y��Xh���\�ʴ�����,m[;�Gg�JV+�_s�о���p���e�l}�؀Eg��v��W<��}��P�ޗ��������3�# fa�=s�W��Ud`�t�Us�w�5�]U�OUՑ�e�g�I�8���j}��ۯz�N��Ҵ�ɬ1	���}�'k<����V? )Y���%5�Z�#�ƅqι�;���OV�ϝ�\cn-$�#���V��#^��WPЪr�ه�N�OA�y���!2��^����.<����U���Ftu�� ���uҚCE4|7�?p��8����<�F�'�%n���|�>>Dq�* h�_%�q6����<o�H"��PEQ,�����gg�^X�fQE	�Mx�/@��0��z&��}�o8�H��uuh=׆���,P��0��Fx<uflnҶod��J���cÙ��6���v꒬���ú�V�u�b�η//�<�޾w�>?��A}��zJ�]�+W�؋�3�0�R�˱�V;��[2��০�|#���?v0Jkݗ�j�牤+ԨUzf?l�����C�����(b��t��>�o������1Y�>!�73{HOǲ�Ҟ�6`�Q� nА4LA�@xU���Ӭ	Ǯ�K�P��W���j�Z���%a�ߩ�S0���ƶŋU�U�׍�\Ň~�����V.6����-0$`+�Or�9_���i��֎!r�@�Ub���Dw�|v~���?)�i�pu�>��/,�ں
�3�su�}>�0]g�[����ʥ:��������tb�C���+�<D��Ұ�ߚ��=��Y��{D����/�N	.
>��+���U��T�d�i>���2z����V�5q��7��V�#���hX�{�^��R
�xN.�`�6u����w�^�o���t��Ĝ�~�vk%5[���`۫|<}�0:�m�Qߓȥ��^P>/7�a��<��Z�~��Q�K�`X�!���E*ﬨJ�,:� j�e;���wT^���E����e���`�\�]o=}�����ڊ��{/CUc��;do{fJl�W��y�+啕hyS��6!��S`g]��M�rY݂��!l4�Oڕ��>����,�cYS��%�yGwQ��[l��a����Jٺ�_׸��L��c�+D՛�ܥ�;՜�C��^�y�>���ע�N��!{S=����,R�C��"��.�2�wU<�z�.gν�;�;�`t�<�*�z�#	u��S�qX��B#�g.����<'z�uWN3`)��!���>�#|c��\:1Y��ܥܝ�蟺�wW5o��he@.�%]�����߼fJ���+a�6�?#|��*���Xu�HhΥf|�zƬF�q� o2*f`��Jp|�Օ��WV�.2'�g����.�oy���/֜	�z�>���վEVPT{��w�����JqwJ�=�}����ep܄[��XgT\,c��J`��頄�< �F��T
��w��y]�����K�}��g"��Pf�4`�}AC�_���m�ܙ��Z=�Q Q�o��#��O"$���W�s�v��#	5��.¡+j���=~/ w���+ͺA�Dv��r/o���Qz� �m����0qP���o�ڬ�1�4��]���prE1vR��=u������q�Y��'-�Ј���sA�=�<�nm�3=�5��7�
�'�ZY	ڼi���ՠ�vu7P����[۝����w*��X�\�g��%z�wv�qO��6a���x�W�r�Z N�Au�E3���)gYQ.WZ&Zw!�-n+�e>�6����ڬSiY�&rEu�=�xwklV��K���O�:/eK�4¯s�rgC�ۅ�*݁e��|�]����mp�_���V"�9PFT�.7W��^��p{Q1^��w�>r�|�Ч�D�u@��2�c����
b��Bxo�z� ����yu%�Y:!�Tp�UHO����O*$e�TA���6:ݷ�3��û|ڧ�[��=�v5T��.uM{�%�p�W�q�Z���4��^����]��������*i�M���Ǯ�OU����_<U�+�������4����Dh���Ghm�t��܊�_MZ|Z�����|�1N��ehyQo��U��C(p�r�&*��-AMPd�����g�bZu��C@W���i_��SK�c�s�Hh���cѽb�ඩO���B�V�D
��үmR�v�8�$�7�"�!��m�&ReV���,��PկJ}�E4w�u򲝡O�{�.0~�sz�oޔ�8��UU�EW�R�9��p�g8�����N�{���P����D����J�x,�K5�խ����λ<�Gn�H��0x�_vP��$
�T�i͢y��k|�:f��O"�W)b�ֻ�1��)���ٖ@������_���L�y���Dl�Nwi���1|�YЊ�D��k
�rl��|F�^*M�o{/X�ܩ�~�Ħ�Ef��w�+��=c�꺈�ā��w:"��t+g��y�^B]nӔ%��u��#
	�=�!)�KD�F��6��u+o�¾S��f��j����W�_���J�����x���u���Q�d�M�g��h�5�{�ش����+�w=�װ�׆vi j���vp/�^u���mӭԿ�I1:�Jy>u���������z�]T��u���+�(�i�_˵�(W�WV�$��Z��:�}��mE��$GW���n�I-Ux��TE �	e��#��k���:9�hwF�n���:�t�|��WEU��R��ϵ*I��͎UC/<ť%Q��#���ם�@��������v��=M~.et��/�2U��UՀ卫gb�H����X�)rY'y��	��OΗ��xx�^���3���;�j�Gݰ��L\iHb���e�8ǜ�K9�N��]�b�},��ٕO���Vx�ޚ�k�z�u�et����u*K
�W��L��jl�K�Ձu����1Q�8{��5��U��F�}�<�c�j���WO�̹���|���Fg���c:����r���p�t��5S�o(����\z�����N��AY�=�(T�|�ݍ�5:�JTL!E�9h�"�����W�"pV����� =���� ټ��O�6T�k�=��6��{§��]^������\�$��Ylᵟ`DG(1I�&R�ӕ[^MvTsk�}*|]T��Mh����Rwة4���gA'I� ����>KE&��~��[�m{��l�Sg�|��3Ǿ��R�=�t�"�l��7�AN�_S�p�Y1�7�#e�t`��n]�����׀̮��OMl������~�0A^�-��7�[�&����=�d�?QX�k 
����`�,e.�@�Z�t��:'��F���z�u�ꦜ���w��KШ��`�#�=a�-�g�Ǯ�K�P�VX�I�t����{��ڥWX�d�$��^w�NQA�4id�(����9��+�W�z\�yM�R�c�Tw�(��%Dr�@�F� E��0	�v�����5R��F����S^ӌ�G�r��:)ݯ�O3O/�g�9����p�<����
�
��@J갧ӆ��,%��ޣ���\�$h��do�������{�z��Z{��E�Uؖ��OZ�z�����@`X:�vqҎ�-�:�IѤ^]��1�ӵ[�hd�ۭ�ѫ��1���ϭ^F����sp��.ud�j<�#����,ft���c~+�Ǩi�z��I� �y����[�uf����{D�F���d�������H���i��␀*=Y�K{ǧR���G��D�Ճ�#G����B��R�FF�Xc�������]7v7�+"=�7�G{}�}���O������W���ݾ.:�*��8��Z��݉�)�rݱ:QPWc�L���8ؗ�{���eW��9���:Ga+E�UDQl�:\�ǵ��}ٰxt�{�z�R���{�ثGOg�����v�ى�cڇ}���U����X���������f`�@	��צ&k���:���P�9��v\7��0�[�y��*�K�z{u��M�S�v�]�ﳮ�Vq�qx+L�f�?�G�-v9[�p�ج�H��o�.��䨗f�ɜ@��O,m{yt(Wma���\%w},S>����y�~�*'x�Ȋ_�ݹ���rBi�i�N2�@�O	�a��T�|���+~�r��Aq�<K=\�VyAR�up^N�0ŪTpς���9E��{�����@{��S?`�J��.�Z��NI��V�y�9\�*�؟B{޹��Ի�اp�~��j��w�6�F��JR�ٳO!r�:%��vu��8�;�U ޳{��\�t�n;��1�O{�=އ1Yy������:2��υ�kL����1r@nЭQ�,�e�ܾ���}�A�ۜ��3�uGܨ�p�`��48O)�S��
�@z��P�p�B�4U�ͭ�3��쩇s׻��ɒ�}A��_����H��&(���� ��=�'ϥc�̉��S�Cm��86�`Wl�}Ä�
���|�}�9����r�L�Y�H��V\�׊�m�ǽA+�<����U8��� �鲪�6�x	v�v4pei��<�y9'�ڵ��]����
>����ӈw)�J�m�п�":f�� Q�*;�.��np����,]��j����*�O��Z+U{`Yg漮̦xW�W��Xb8�L�8"����#�xE��36;���dp���qB���Ч�D�t�(�:����p���ԡ��bՠ��蚯/6YYj�}��+Mǒ�!�T��#������QP~3'\VUi��d3� ���>RY;����nOh\����J�Ҫ�n;kQ��a�	d�9�L��h|�j�J�_�a_f=
��/�S��犾��b�Wnl�������4���;{��Z�^�a�1���,�jcU���u׶���*���GDv�n�i��ל��	�Y���8�r��3MV�3��szD�/��/z"� c�;���h-���%��s�ZX�[���S0vbj�,�OT7]�|�k	H.�ݵ���E՜�u.���h�r��|s��o��?�VtJ~LS�;�V�������;P�2\�pɊ��>%ک:��?e�z�Ȃ/{r���Ҫ���4��>@W?��6�KYԫ��\⭱�h��o�k����Yt�}�~H���LVQg̢J��ʈ��m��.�&F�?6*�:���t�C���~��|���o\�-���0���@���:>Cø�Y�ͼ���\����i��u�Jr���3yW�i�^�#k��b��="�����@ՙc5ķ��y��30�\*}D>2�О65<�N���w����=C'L훧�l�n�pV�=.�ڶDeW��G��P�(�+��/+FK�h�XW��s]pEuP#8�I\}C@���
s��gr����t�=�AG�8<����u9,�t��d�3�����x�2�V��{��0��c��˘Ug�+p`���ta��vB��N�C��·s�ɥP:*Ϻ�GBTr���91��ꆂ�|����iPzSטf�c����{�t���V���|��9˥{��{
u��wm�����z�V�rû�%���o4o���k���4E���:Џd�#,H{��@
���TB���z��Q�Og7��wgbW˹��v����]��3]�6�7���h�>՜��6��;���ǫ/�/a�g�8�Ͻ�~FY�c��6.Ug�����hTbᴇ܇6�z��i��^��z�r05��v���yX���({�2U��UՇ2���� )jv�⮽��c)��b��y��F���Y7*�s�+�����}�71C�n&#��	'��b�_ߐ�����U�wRg��� ݳ0����ٔ�x���4>���к^u�}e/Y5w:�3jf�{��l�t_-�3�[|z��{%Q_@��Z��J��׀�g�!�k�^�������O�υl�y豛�OllgE��-���ϲȈ�)2f<^L��y����y��)W����<fU`��7�4HF�y+n�����٤0si,Uk��}�;�p=ܵu6&�nӡ,�6w�E�y�l���ӃDpڄ���EF�ǼH4g�e#l�q�J���^����|�˰�ׯ>�-�]Z��ٌ�>toO��μ+����[͞���(qa�z�Ί�(W��}��<)Vߞ[m��i�^�1"h���nĮ9�خ�|�t�L*��d��\[h�si�ET�r�v
i�w����9�7��=��0/���Ь6��0ч^s��=� 8ma2P��8xS��x�.{@b���Tr��|.F���6y���{yd�AC8���`�AX��G��M�z������Z*��GgVK��v�"[���꘥�C��nӉ�Q�9Ǥ�d�V�
���7�Cu][S�"�#;���/;m�g��$F�o��z<U�	�G����}F��"o8�Skc�5(�|&9��A�$�^�����ޗدwYuSrѕ�>�;u'b�H����oY����e�Gn��{�C���x�g[+��;��8�c��9V
/5�7���]H$m��h���i]�D:|V�B汷��v�nŝ��lP��+y�_[�0e]!Z�@,��eռ��jv)dt'b�pŚ;uq�5�D���+�A��@��[5��"&�������+Ú1�d�Q����o���b�彌>�#g��BB���|	T���5�k��f٣�֍|��p��b�oh��q7P�u{���H�Ϯ-��1�nGeI[r�l�mB1&M��A��VA3�������k@���Rv�{�{CQܲ�Fe3��tf^�{/t���uu�&4�:6p �e�o�>�!R:(%[��Xv���;�y�*9ܝJ�൅B�"����7�u��캝�U�	�"W��Z�^�?ttI�x`7Ϫ�c�WG�e��o�Ӽ������&tN��m}\_���aڹ���;xP�:��-S_b������(�g8J���39���qs(ؖ��wx���ltY���ʗ�A���>_# �9ڐ�]��\[ j�5�`�=޷��8��kx�F'fin�����ܵ��fV�ѵ��
��\2���ۥV�IT:��h�U�N��
+dz���GK���Ê���^�}2 i�#�Tox��j,�إ�+���0v���C#\vJ�;,U����Wc�knv�FWp�Xʢ)Ҵ��\���L>�Y�7{T2��W���^�b���X�"cF�O�{)�JΘܺ�t#���{k�k.�2�ǎ����81��W���g�l�����<���y\9�^�N�e��@:f��N��E�n�y����0'
�ڔ�c��U��z�4xU�|��k�/TF=�x�b��4��]���w�i�)Q��%i�7c��_�H�7Zt��W�ҍ�8^�2���r+�+��x�ˎ���d�U6��u�����*{�3��yJ���W��\(���C	�����H����m�է�*l�Ґ��qU�fT��rGmvS֓ۗN����Kpc}�-t�M,�\�ѻ�{�3̎�uN���D&p�qf��n@som}��;� �4Fj��;�xrJ�P��pW�VN|�D3;v��x�mW#Ƭ�;�O��5��r|� 77 H3��5s��c�Cd7w(1�R@��I&��wv%I�܂��d��sB���롌������Dms\��v���$Ӻ�m�0�Cr�R!e��.WP����Q���w]�����$;�S ��C���2H�X.\�M&����37u�h�(�H����RI& �::먣	59�;���QC�����B0R#��)wt��u��e9�Y�5��ŝ�.]6g3�A;��C5�\D�E;�b�wW	4�&"���e	��@h��1�*��k$y�%�jm�B���I{jf����b/�*�ڄM��D�po>��A*)[�i؍b(X��vO$6�!{X�;��y^���y�=�����+����O~k�~�KA{���"�_��������u�W.m�nr�����+�η��m�z�?^��:�6���=�ܫ���_�>����6�{��Lh[U�~�Ci�P�<>��H7߾y�����/>}��צ�m���_}�_���h���y��w�۟*��ׂ�r�?��sWwj�<o�>y}k��[��o��W��5��-�~�zZ�nz��>[5����w�Nf�_�"#�}LC��zm�ou��W��m�v�����=��.o������<���sz�>�_�Ͻk��~|����V�������m�o��x����ס��>/����w���ǯ��?Ҳ�*ve�6�q���H��b$8GW��W��o���5����|��꽭�\����=|�}W�Ǧ�?>}�o��\�/���}����+�����j幾��J��}�M�����*��k���w޻�y�ٞ�Ҽ=�]m�������(����7�S������o�w�ߟ�������^��������ߟ>���okţ������W��o~��������ߝ^�z\����{n��U˗�?����=�}~��T�8� #�LX��@�u�k��7�nU�^�.���x߭�z[������W����o���ow�~���\�w���߽����ѿ�>���v��p����P"">�ɢ<����r�g-���S�?U@�x�
��APW�)+����x�k����^-�5������Z|���ץ�����������m�v�W�zU�s}m�������Qo��*�7��M}D|�L�{C����n��9����~��z��K�ߏץ_~�����p���^~_�}k�ױ���|ߋ�~+������~y^��^7��W��y��h�U��=����������z[�\������x�-��湮_���z������I��7>x�G(e�����]�og���s���n�w����߾o�ޕ�K���5�om�ۚ��~���������7��/K�ǋ����޻W��[��{�:����h���{���׶�/��z?��
���l����uo@|"8DH��ڼ����{�y�ռU˛z�|�������\�޾y�h/������^W�r����~|��~�6���ϋ��m��6���*�^�6�^��m����um������{�
�/�_a�����-I*��S�륌����O\�H3bQbݷ���K����%��tA܆Z¬-�,��2T���{�ϵ�2��N�-������kNv�@��x�u��#0�6`Ԁ[%u�*�F��mArV�����!77�,���uoVV](������V鯨��}LRG�p��z_yݷ?˛��m�W�-����z�kN�]������ս��߾j��Wּ_￾W���W�~|��?Z�W�^�}��ήX����+o<��?�K�����Ϗ?��o_�����oֹ�7��y�_�~��wo_˛|�ߞ�y�����ߕ���^�o�w�|���W�Ϟh�-�o���ր����"�����!���������v����6m��т$G�8*b0DH�����������^>+�y�ү�湧u����_/�}z[��W5��ޕ�_�w�}m�|����o�nU�w��~z��s~������������-���?Ϗ�{G�5]�g���T���G�H��C�0|c�#x��ǿ�<�������y�~�mx��~]�TE/������v����>-�W.W���[�|��x���z^��>����=n��"0G�,��u_�G��=��|������v��ۚ��ok�����Z��J�s��������^��\�^���^�|�\ޛ�ޯ^�oO�ү���wv������j�9\�|�����z!}#�}b]���F5{�9�v� =����ok�^/����V����|��ƾ+��|���W,/��}���_��[w�~o�|���W����/|׿ε�x��ν/M�y�s��׶ޗ�|=7睷��>��>�L�5�]4e�K6Q2�č~��_o]�߫�x��w�~�ڼo��o�����^-���޷�}k������K+���_��^U����^/���5�W�s\������_[x����ﺈ�X��Af�\��:������Y�����W�w����wo��r�~��^��[��n{�������o���x����ow������s|[��s^���h�|������_�}yoJ��������b>���69/Mlj��wC���|^��W._�<��{o��o���ޗ��+�v����W�O{��W����[s~o]�������{\�W���ߟ�|����|�|��o���s>}�o;����/�Z��)A��N_�+�[���|I�s���zZ5~���i��Ӻ��y���x�5��h��Z7����w�/�߫Ţ�믫z~����������W����^�|\߭���߭��ү�����i��νPՃ	��7�Rå�tvoQ,p�Ż�q�4��d�3U�X%��F���>�mZ��c���;�X� 2��b��:��0�^l�ΊCmX�b�h�b�	�puO�Z�r����-nE�Yo]��v�
%Cl�6�k;nl�-)�U�e'���۞R˩�P�^��������>y^�6�y����|�����oO������^��n���)�׶�5�^���+�ܼ^+��{��ε��_����W�zZ7���߭��^6��~�Ѣ ��DAJ��~gm���{W���q�b1����^W��`�� ��Mz�������>|����[����/߾��^��n����}���~���>�~�soM����ߞ^�x�����=�y�ž��DEɍ�>�>C�ו���{Η^f�x���5���Ư��x�Z�/�������W��/�>����߯[�>-�]����s�v�/;���׵����|�y���x���]���o��9�DxE����>�{d��2|�{ �����ExfyHT���D`�4}�� �[�{�ޟ���?z�?=�����?��~o�[��ۻ����߯��AW��_}{[��W�N�ϝ�׶�����o�{�~/������<#�">����f�H'��{����������oKs�_����?:�c���k�_W7�����m⯋��}}m��sQ��]�+���u�/ޯM�/�?7�Ϟ��͹���[}�ƾ�����D|�1"<>��i�]��NY3������|��]k���w+�_���}��y�_��om/�ߝ��\��ם�O�o�y��/O���|\ߗ��5�}6��}�/J���{�z���r���]}���|G��nwb��2�����|�{������uzU�����/����5�����~k�^���7��y�׍�x����7�^/�����y�}_��i��sx��V����c�>�~�w�}��n�</f��߿�j�^-���ͽ|�+ſ���6�o־��y{U����������m�W���������j-����O�ޗ�;W��76����o���F���#� ��˽ثz���Z��F�u
qc�������ߞ�j�x�WƼ_�߿}[����~z��ֹ-��U���������������\���=c�����:��f�ssk�]�z�/WO�=���!C(	�_T����N��X�`�0_�黰�4Cܢg�/�4�i?���G�fL�w2B�8��mV��³�+fq�ڼ�܋�.�'DJ��vJ�MQ��dY���L�$��QZ���HJ�w]�(���O���T���9�wnã�Ff�V�c� ��Z.t���[Z�C�T�u����6�f���L�諭�`�.�ZS�F�N��� ��f��L!��<=G�~�r�;�+�� _��e��]^��P�}r�Yǟ%�ъͬ9Z���@Q��8<���<=���\���uLb	����-*��o�pCn�NhuU�2W��ɇQ�b;�+p`���ׅ�n�U�=A��A.�)�����L慩UѸ�����4��3Co���#�@��/�-YfqO�ؚ;ェ?�������/�0f���{��w����� Vw�<�I���
о1p��*�?�#�{��y���g۞`0��#Eo�<�DF�pb���d�|����`�8���٤��=LR��lk/3�!B%+�����g���꯶.��Z>�S��F��}�ⶐ�94uYW}[��k4yg>���Ȫ��ë9M��>A�<瀌^ޔ�����'���U�zq%_o���k��v�q�8Om���������P�)�퀶b6ݯ>WV��q��n���6d���*��|�߳���]��$���g��ЈΉ�~�ô�k�zN���cA��N7��Vo�.��;]�a���j����+Y �M��8��*:;8^��dܣxem���*\K��a�.%��y�����pü�_enН��J���uֈ�sk:�M���#-��՘k-�ƻF=�(ʿ�����n`��� �d��f|6�J�+�<#���I�B6��I�b���a0�$�~��.��UBz�7g(!}w�Fϲ�̤��ȶo���|��3�z��R=��+���V��~�6��Y��w!�H��k�yL]LǑ�����G����?���A�ߺ1W�y+r��O8�f:
����RxmUX�UW��Sρ�K�<J]�>��������.�{�	��^c&	&�GEfK�$�H�qW�@�;����nz��	oz]k�O9f�}M
c4��A/�28#0�IV�*őWD�� w�4��l�kG@�[D8�u)6x�.�&�]{���aI�J�
�kB_�c ��죡�t�(�h����+!�����)��N����s�=���8o�]ީ�t�&M�%@ydZG��WU�:�(n_�����x;��^�
��X�����_�n���'�/�NIpQ�慾�hu��6�{Y���<�ǁ=��E�Vd��ƿ��Y��+�&U� ᚽ����#�2j���6��r�˫��YZ�ъ���5���W�x�{l���P�Oe�tԅ��^���:�7q38���<�x�r_*�+A�KS��1�$�GIMA=x�:§RI+zs�xS�ӆ�"�A�4�Y9�C�ۤ��Ћ/U�t/Xy����X���^^����]%�	��+=�����ְ{͝AW� mgҭ!\�+�m��
��![�Q�WN��-�&VE�\E]x�D������7�+�<D��+�o���j�⽬�D{�ϴy7粚��.���;epy�V�]J�W�{Q���Z�Ţ�N����Ho����^���IϘ�^^�@h���,��j��)��o%	J����Y��aU��t��olcK��w'kL`�'y��Cr]R�D��qx+L�f��/�N?C]��y�U.��V�:���Q:��v�>exm+�RZ�F׷���+�J�>��*C2���ݸh��g�4��~��y�~�^�+(���~��i�>iWN��N��k��&�+�0�jf���o�$����Tx��f��#�Y��'fǅYo*�φ]���_��a�,|�E%#o���+p��ݵ�GM����@o��SC��;@�F�=�3��U���������V$8:%�S��K�����:��$ۭ�����D�u�՞��Nd��Qև�=4�8�Kϻ%w7]tgI���9�f�e�TE��t"[;)����4��{�˻̫K�ǅ) RTXs��X�țg�����x�*�;�u�Z�M���ؠ�o��,Qٴzh�|�au's��2f�3"��}��UW�S~���QF�p'M������
�:Hi���vJ�.����V3��չ~�2�\�/o���ב3ԇ��"3 ��:��t��\9�e��j��ϛsL0�:R��,N�T��)-z��{}v��N��b��|���"���ӥ��Ĥ�q�!�r�����V���U��˅�N������֑�=�@��c:.`/�y�V���n{�uי�{֭$t�[��ls�6�0sMߪ�3ho{�x�|�w����� N��`�:�������h�G���"�מq"M��"��Q�{~I�;ܨC��'��ͱu�<Fb!���E���[��Ŏ�<�=����G|�r�����R������.;R���{�������^��ם5�l�sٞ�L}	�;]�;��~�uW�}��(Ep��]^���Z�7[)W�o_<�p���G���B���W��p���:\���^�����>EA.�׫�њ�v����3[=n�5.����=��T��Ѳ�������u�4k{8��;׮����|��}����dc�|�XB�$d�/����\�O2��㢎�ru��@.��Ow�D���j��K{S
��={�* ���vҁY��F�{�_h��U�ȵp��R�^�n��Wu_q윌2���Y۸)q�ZK*=�k����n8�����e�9�
Q�hq�&�[]Q\ϧ���R�Q`2�+��D=m��u�3�S��gw+�.pY�]K�
�.�S'�����{?�)}�Aţ�@��̃�B� ��p�y{�ެ6�}+����B��B���'bSG���`�6�^2�K�]z.��(�	�>�2k��꤀�C5С[�Ee �uK�D.M��'|_�	,z�K�v	���;������f����%�(X�6`-��t����O�_{���.=0�Z�޳�뚽�������L�o�꼧Js�i��Z�Ҩ 4*�py9��T��ڤ9}~��Zi���������O�����'�!�GMңx�1Y`�}�a���nW#�����D���u�wu]�����R�ҳ�3Co�	�Rz��`��[Kw۪Geg�d�RS5}{�a^3��:��[�hJI�과��68W�w�3�ZPxZ���b����FwMg��ľ�JR��\ή�<O�7>�"x�9��K��,`ݮ�V�ӊ�5�ú�2�4F��t�I�m�"�A�!� �E�1������[�ֽ	��C��Q����uZ� {��S��c�,t��=Bw�8�<��%3�kj����h�=��[��vʼ�Nn�#�.4���ﾪ���p�����v���,�;����2��w������������w{
!7k뽦s�bΩ	�kR�߻ǘ�L$1xU�N�W�.�<8���x��
���D�X�Ϣf�S�;�����.`�+�s>�;�T�vG��{%�h�:q����z��׫;����n�g�������i�̖�z\�]^�߰t}�K��%���C&���ӂ����j�K�d��ﮍ\ヮ�/S���AԹ��$#@��R��};���X�{	���q10u�9w�Լ}U>��.�P�,�L���v�Z|�EaCD!��\!��*�{|3��ɖ�
o�n����AC��D��r��Z���nƌ�
�cy��[2��OMl�;>+}���S�^#�ab??{�t�������/�� #�}��¶��1���}|�dg:v���o��ӓ�{�t���q>7���J`#\D΂���tuV*5�s�j�����D�oIJ���B���%9^F1ф�Ф�Uo�gN���Y�"���^6�����VG���r�-���'~&�&�(�f�Ɂ�/tR�^�Pְ�'�|��w�yjڦS�tw��ҋf�7C�y��	s���@��OA���wح�U����6��̜%�}��\��a��r��y�_��ޠ�v�X����dY�6C#���������!�'V���@���q�� �	fIj�`C��F��R��U1#�T�5;{y��yw_^�u"��:Շ�k<q�X}�����wz�Wt�&M�%@yg�V�^���Պ��z��}��ݺ������S��K���/y�r�af˕����~_q/�)P����'�f��c;�I� ��ʅ�(�t�d���?�z͇��~5>c�m,�7�\�E^$��Gj��}ZewU� ��<'m+��q�u�I'j_����:�=���\L��3"�R���(:�nQ�E-Ct��߷�Q�Kݰ	�!�������'��Nj�;��xN��T�ª�7�k�wbU"�W��{�ثz{=�&
ӬĆ�n�P ,�磊���rWQ��:Y�;��}ŊUL�o��pB��\�8Tb��>�Ws�ά���k��畤l���V=)�ڪS������/`)�ò\����������7Fc��ѳQU��0��- 뢼6��%�D�׷���+��|�_h�&J����kP��z�_���cW�݁�ei4�뺋����H�Z�B�7J��2|GDj>�wܪPC��p���S���i��]�b��6�E��Ӈ���Ix��4��JRs�4���Sg�ӆ��C�=|��V�wΚIʵZj>��+M��X0���7�z��EM�͋ձq�.��-������Jϓ.1�nk+i1�[��{�J�O6D����E��I�vY�y�(�)��p�:��)�~�Rr.H�բ.(�M�t��1B���&���I��B�n�n�M�>\��R�Z�'����4ٜ�X�'�fv� �rF�|��/��|���Oz����hI��N{P�c_Y�{�.砃ʈ/sz�Y�*��sRv/t�l�1wwV++S�d`�@�@8i���Fes�;�2��s���5Aۇ�9lU�%>j���"v�)`Jd������޻�,�I�g*�j�ڽw��N�b����{qkR���=��t���Uk)�9V�h�˵����4��F_t�}ϳyD:9�M�	+�ϵ ^k�G�ϺV>�����ՙ7u^ �[�)���N��Е��+r��TN��u�b���诜ζާ*s��-j��N�s(W�����-e�Mm��@� `F����V^�b������*��dv>��|����4���ܫ@s�əX���z�:��ļ���>�)t n��+;w�i�ˤ���м
�Oy������o�m�xE�%��ۜ�ޝC���.}�k8��ʆ��L�����ӻ��u	HJ��n��x%�`�cX/��w�(�p�=r?ov3s�'ſLV��L�2��4����݆�h^�[�UǢ.���֘�VoM�@�/�d�R����eg�\��967�.�#���(�ܛ��t��2����i�-�ȣ'&2��~&ޫ��A[�$6v�Sv�������� �Ԭ"���92}�7;5+��\ǫ�36�>&���ޙ/��]H�W]9tś6pE/7����s�.{�g��a��dӌ�3>�PA�]J��{{:��Rfwe���1m�k���H���\��nt�����&�;��JJ��,�L�]�D�K�w���1ZWv�����hy}�if�ɻ���Mb��4,��]4u�����"���3�m�LH�n����n�����W]cKnrskd�'h.H�I-�ќ�K���C�i��5W�{Ȃ=#�VEk�+��3�� �eJ���ZC�-e��c��NzV��x�,H㼠5\(%}��ToFR���V�Dr���>����R�|v�!�le�;�u�PO�7DE�m��l�ik�.���c`�E��j����J�!yX8��ë��>�[O/�(��)t�k!r��,�*8ǝx����P��f#�r`��N�I���t͠�O��fG��vWl7�Q}��K'`o`���Z u�:���#Mu�ç���~�?}~����!���&�5))E�b˱����I���(Cn��;���`�(��ˬBQwu&�ȓDDd-�Dd64�wIN�3HF��C���fTȯ}�-r���<��\�0d�iT�u�m�@Ĕ$�(�6�5�"���G:�(��h1<]Lˡ�s��1X���ȥ�\�F�\�L�� ��mI�M�]
(ۜ�o^u�A���6�\�-�M�4�����b5�t�<���%�Ad��O�9��ly�.u��Ӻ�W:QF�P��Hs�d���h�] 7�Єo<�<BFg�v.�P U���|{Wi�ɔ�%�/ir��������"5;��9���w"X��ռ��.�i��V��)��-�';�����}�}_}�\��]�#չV��OhJ�~B��:�Q%�7ꫣu��p$��g�}xMA�����>��!��}]^`�D�a��aQ�M�'#�Y߫���c¬��ٕO�þ���p�<3��̽���ћjhT�J��G*x�-�#+�48MG*�Sq�
�V+�VJ�����(��y%O0�Z*W��3:�4s�[���6xK�����8�W#�J�A�<$�xo%�]��V�4��x�0�� }�xB����� �|Hx���}.¡+D��K��UZ�X�N��?M��-k奏y�H<H���ů*�B�l5x�ćw-ww��ӳ������ļx|1�+��j:�� ��o��䈭`�4�]��J]+Y�9�!<�3�����%wM�o@c4��*CJ��*�k7�VA�+>S����vς�?���^�c�B(Iy��o;�9>��ɫ��K�1��c�)�LV��B����v�h�g��WG�s��f6|��42��������>-=�@�=���g��Н�H�_�����C�#�\�L�ӊ�e�n�F��rm-�y<���NW��� i/�X�������hqfgPϲ5��aS҈k��!�z�����Ѽ�Ρ���:Y�c�W�g�����]���Iwuq�t�㬝|��T���ۣhP8E'�O�Sm�g5�(@�HS/�m��U�W�W�#��+���K?��V�7����TfOhjͦj��^gD����qr���y>�G��Μ��5����9%����4�6#�=���Gεy��~�Y���x�\�^�ا_3"{�F�+L�PV�+�t
��x�WK���N��q���7�=��)%]��"o��lؼU	�Kl�Ɋ��w\��~�G����ݥQZ�O�^�)��i]�̩�0��5UkW!YSb�!���B�{Es>�)�b��v�8�$�7�5sۏ�J�g,�?���n�敎�L�"���Q�B1�h�ҷ��yV���l�zr o+�1�b�J�Wy���� ���]J�!���0�KO�v%4Uz`�{���Z5㧇
��sr/��=K%�ӽut$�����r�m�T4�3~U�d�i�&���JcD��]r��u��M=���M݇(˳�5A]1|�����Gp�η�8p�����y�K�O��vZ-�®��w�>��N�~f}��B��E�JUz޷��̅�};.��M `~6�)�;�;H�p��V=�p�G`D��v�W-
��Y�3u�f-�(�hKէgl����Os��+<��R�e�����B�g��m���w��h���]ԵKq^�0�������gq'e�)�@��AO$�'g��	���� > ��K��ɗ�yu��}RK��3��T�a��V�_c�ɇQ�b:
�m40��B3�f�W�����7u�/V���-�x|"�)@iY�hm�8��0K/~��F|���m�sfP�+@��X	F���@֊�",��Q�ݳ���z��*��a�_!F����:-]�~���kM�*Ǿ-`�B���^v.5�O���pv�����Dh�(}.�ZK�5��M{Vb��W����W�DvI�f�j�r7���	���%h�so ����P�r���.��%�)�G;O�ݛ���w(������)��!՞ VJF��q.qYx�<�xWi�F�ȧ
�s�]������V�<�����
�TN
�|��5�|x��%wr��>^� # _Ѿ��S[�̔��]^����e%��(�[7]T�!qȜA\w��,�C�P��8]�[��8���D�o�J\{Uor�k%�3u�Û��cr��`$�RX������M�8��g�����<lAb�_v��|C8"{u�t
���B�(H��\��Zf����C�~��k�0��b*&�}V�*ƙ� �W��,o5y�i�GE},S�(���ښ�.��6��t�T�.y� ��]��Vgn8�&w	�t��s���X�Βs픐m9�An��CT_�_}U_|%�p�z�-�G�Wy�@��#���+�b�c��t�;��(`����p�uj�6��rf�X1�r���*�!XܩG��@� |�k��Q{����p�u���d�wX8�{��M����$N�����w�}%���� .� h��@TA�ƅ(��ײG�t�{���Un�fA�Ӭn=u��#��'$��:p� �]:ϑM&�vn���b���B��90�i{��{���^8v%�$�Fp�=R��G+��V*�坾�-WNȟW���� ���꣋�o_��Mv�fa�.�������<���H��@�M���\��/N���6� {<���uF-��k�����Y�u��������oK��z��WZ�����ljP2�\���B2��Dm#]�AU�f�f�|�ƥV]��+iӓ㉥���rzx9	;��_rT&8N�r��>Y�Vut�v�����7f�|�{Mp�e����\��Og�J��+�WX�èͳ�:�E/�R��ޞϳ�7�+�G���؜p����z���guɎ�W��E����h
�@]�/0�V�{�袮���`I����[��f�#"��=�׍1��]��ڷ����e��e��o�Η�7:ә��e:�zb��͇7|{�(��1
�n�Sú���i`��W�U��a��k���i��ﾯ��S����Ƃ:�� ;�z�Ϊ�@Y����!,z*W��~ǌ��XN%C�z�*�]j�K��#G�3<ta���*�j�򘡮�������{~sC�3�0'�|k/;�����sg������GT�������,W���y�gx�f\��]f�U������V_�>j�K���z�:�+�]�pt������x̕�~��puw���eM����}��0<w�T-�Mo��c�}�I<C�xkJ�?�Z7�c9IM��u+F���VS��j}���=fh�9&��G����N��-�U���n�5>s��12�q�.���e�r�wJ�ůi�����3ب�u��Ù�/~f����{����W1]��9����eu��*�G ����6z]��	~Σ�I�KFL���uRsS�W�=�r	8ީ;�d�r>GiB�Q��x��[�v	P�d�R��!=���X�p>�V2��w���+[t�Ԉ�p5ʼc�٧g�ou!�\�4~S�.�/=�O7~j�Y(])O	��T�L,����Nȯx�r�^��d�&/��ϧ�quh�f.��a׍�ݿNKT�o߭���N_֬�3YIs��nb^���#���=Q����;,�u�H���J�Vn�Rm�E#�y0���������|�>�&d:x���]>������䈭t3N�c��/Yr�p�H��wz+;ތ�Sʅ\��%wB�Dt�%(�U�}a����Q�"��Ae��/+��kz�2v;_���L�����B8�%f����P�1��&+}M!WY�	�{M���Ʒ6�rf���*gWy�v��1�0W�W����Zk��@B��	�D~~��THά�VWd��3���=1{�w-M��z��atmX���xc2�x�w'�>Yx��5+�_I�(#�YB�N��]�;u��"� �.���c8p�	�1}Β��\G�ma�/����g���댩������7��s��W��zf���ai�
��Y\#�V�
��q�({F��Y���)(����U ��B�vK��Ɋ��w\���ﴊ���7񵎬����mG�
����G�=ȃY�E-�c^މ�2�{E�7莇���Q�,�(��c���7�o6��~$e��]�L�'�nwRÑ�B1���#��-�p�*��\[Ã���Kk��
�Z���;t���2wm�Yң����$帪����]�v���9�j
�h�z����-JA^x=�݋ily�lԧ�k5���+��ά�mN�YW&N�m��u��ӳ][���Ĝ �U#-w�w!�3j*�O�,��b��}U_W��ET�W�GԀ2�ĝ`HC���m>~ф�Z|��MY���tۮ�w��W몼�j��91 �Yx��B���x�2|;�o����
��xD�i�oOiʱ����\ݫ�h�q3#��'�w|h�<v:������^�꣸~�f
��4��Z�I
�4�RZ�a�5̜�o�%�њ�?3��ݴ ��g��G�����M�v�^a��ՐzM���Կ�����Jw�huU��J� w�0�FɈ��mG	Q9��ͮ�Е=��dE���"c7�hwt��>Q	JJ�3CB�09L��n1��֪iU{�}Y�U<_4-����[Dc�b��n�Ԟ&�P
M��m}ʨeg=��y�WR��i��{ɛ�]�> V�F�k�>V"�����G�y���ճ�o�UL�45zʯB(��{�qJ6��E���M[�^Vlr3���r�nZ�v��ҽ�S7g�IyԕS����%{�F��}���Ƌ�6r�v��"��P�+�����M͸]u`Sm����A���%���5�Dbo7�*�"o��5����ůH�0���f���������dOޏ�;*vh^�Y��u�⮞!�%r���3hdX5�魝�����-�$�k��S5��s������}1zg�.�U�P��A�R�2%To%?f��W���r������U�	�4���)ϻ��k�#��@v���*���ؤ��2P[su{�Qo�:>ܥ�h������d�#�gE{��B��Ҍ��"��Γ+�J���:�&	wJN�%�k~����za��=�����$�z�
��iP�fRgY������)u��+��wa�%�	?ep׮���ծ�i2�{���w"D�j�pQ��ܻ
��ϯl����l��B����fl%�Ei��=���z~�ʡ�dK�:�̭|p[�N��]�;���}4�C�.�{o����7��7�x���t�Ut�ILk������KyT���Y઼� ��+���VW��!^����#ƌ&�U�)�t�pu���3v����E�4X�6^��e`�����x�]|��.�yW��&*3��T�Z��svQT��B�|�ｚ񧋚�P"�8�������fP�~8>�>���t�p�.;��	���D�EjJY�[R�Ḱ�1,��N.�ag=��M��d��^�f�p���`��@f��EU.��.��]��pE��`w���k���܁zg#t�}��MĮ�� ���5o�Fo1�ܩ��������Y�����ܐjm�}�U}������z�G9����Wk�V���: K���R�;U�Ú���xF�=�O������V��V�D�%�G%{ь��,���#i�Ϩ*�½f�ax��o5��y"�.�zN髧S�"���eQ��:�k�3�N��>�'�����]�i(����^����2N�u��R��nZ7��s��ٷA�K�~��v��ݰ	� \/���Y髢�v�K� �_{ ��)`��TS~wj�5�w���;���r��������q����?���^�,¾,_�Po��L��W��t���"��x�a*�6����I`3o�>x,ş[q�Ë�Ԗ0����v�E3ڼ�c1���kD�Y�h��E��f���z�۱��:'�t�|��y�����N�=O�#����^��檝��z,�{�6{��m*U!�soyt����=}hɾA�z��r=�I�o��:﷗�+�K*ʂQv���{O_[Dή�ݴn����Ӏ_r��Ln��)қ���8��]�+B�&�=�v�٣<5Wco��,&�o�R��Й�5g2��h�[�[CZ���*�Wp#�:7@�
ڏO}m��*��ue�;l,[ۃAr`�� r=�q�7�(���}_}T5�}��գ\�G��{��,�[KYؽ���'C���g�Y�<D���A^^f���$��C��T�^����_Ǘu�#{ݟ#�G'beQ5�ƸA,�ʫ;Z�3]jх�{ƒ��<E(��M�x�&��K�ۗk�/x�g+��K�����]r^ZnPƫ���:K���ؖ[��#�;��[�6���f�p)�RT���.=��1��w>]�^�.����ckNG���?U���I�~m�끕��zhf���aM���p��VhON�׭�A�T5���~�<��sf�)�~��e��_�o�,�ūu������J�{�k5{��*�ߗe������ǎ�Y}��J���gX�̜����̢�#3�&�Z������1Ns�fA�8o7}�,�)��U�<����8�{��#�-&t�b,����x�͇ٔ�Vo�^�N�bs$�Ǚ�oe��w+U]	�Σ��n�#������Y��#R�h @Bl7���<�a��&o�Go��}Ԏ#��Z푋�{.��;V�7)��-�Z�T�Vnt箠�÷WwJT�\���7G����rƠ%,c Z/�xт�1&��S�2���׎bCe����;��Sz���ѷ.'�eI�j9�����}t����%����rW7
�[b�WR�t���q:�^Ι��BUh��Z�lm�˸��K
�� 6�oVg,y]�/y�i�i�y�ɂ*Y%X����]�n�;��V�r���o)P���C�7d҄�|���;3��ܵ��p�o�Q����LQ�k�P����a�J<���l4����e^trZ�$���6�-�dT
�j���ұ@�8J)����x�mق������F
-��)���So(�Ao8t�^.[.we�E]�Nk����SUe}۴q:�Cr ��V �]�4�05�]Y�0!��=��[|Q�\6��»:�*��a*��>��X�N��-Ӣ�&��N��4�-yC��|2D)L�m�d�5k�f��њ�o�\L��ύ,�<Gv��p3|�%�PX��L-k�[��ZV�'�G �ΰXw]a��]�r�z�D�w@ʴ�y�g4�� f���|�ҭ�x,�g[��FJ��02P��VV���$�.�粴B��3���A��Eubxu���6���*�B�2�>0���(�R����BE�Kd���܎�D.<���K�L}�>{:���םБ��V�[X�pV5G^-�ȝ2��h���:��g�"Xn�J�L�}W�;a���|մ+x��5gb��;/�vs�/��],�[d���/ek	�e%gLe{OE��M�o�ݮ%��;˨�Jռ�k�qF4�]����� {2᥀	%ut-=�"mE��)!s���Y[��\��L�)��-�Nm�ή�h��8x��XT��pHzZ�ӟjXh�P�V�`jR�8GS���}��c1��ngu���&#�q ~a\�{���u�����x�;\� b�m�E5N��[��m���c������8�5�vT�w��sk��Pw��`�3!l�ZsD�KQ�p,>�zܵ{0vV�|�5��!��[�Vl&�s�c�u9�� DTw5���Y-`Ӯˇ��ʿ�!�Brfq�+h¹� 3���������$�Ƶu�X�[U|5��a�Եp�;���eAXHvo�G^gŭ,p��pAlS'��5�bᖨU��� �7PZ�μ�7���C���6����Tï�QJ�v���Ԟ3ϳv6��M�����Z�S�F,����Hgm2��fv�G�b�x����]�R,RR��<'n�[=��n`B�������fպ��J����t��"�Y\���Meܧi U��Ux�q3��o�̮��f];p�=\��us������~w竿ߞ�<�^ۚLx�����uwv(�]ۨ0O:����������DT���/���e�eδ�s]62P��J��/�ι�D�\5wqw\� o$�ss�r��"�̼vh#&ЖH����hԞ.����b���x�<W�4n�ۑV�'+�n�QQ����Ҹ���v^9��k��vwN*8$:�ÎN��j*o�ή��,k�p�r�M����r��j�X�9λ���r)�S��&�,I����r4b��J�^.o;�%&�����n[����q���ĳg����F?B���9 ⻢�";4un�Q�+|��z���M���Lm��e���QӔvj/6���1�Tʹ��������?Z~���Z�_t���/'z�ߺ���=9�������-�펻��R�Uu�4��^�=I/����`q���R�Z��9�;3����g��{�OV�z�1o=�9�'�[��gS_W��j��zn��������R�4���{n�ss��G힦���3�^��y/��W��Y�>�f����z�0}QU�l�s�_^|[\���w����_j�*�!��fr�*qo���?Sb��+�)���=*F��K$@����h�v�:suG-б�T���x�j�Sׂߧ�&�W�ƥ�e*7[&����h��
IlT)�52��H�b��<�N�O���������3��>w���x$���: �seg��'ZG��Cj����n�{�J��ى�N�:�zsmݡ�J9��z:;�4vv�_l�qQ���`�W�r�rSsy^[{��&���8��nz��t�bm�oF���[�����5}�r�u>���T^t�۫p��{���+�`$��o�9X�o�>�R;�f��cg2�1�!2ʤ�[Xѓ��΢;sgMN������:��YڽꚣӬbX+ڲ�v\�|��ܳZR���lb���.Q<�8�V��T�=���0&*e}gҒ�K~�V���|��4�zS�-�βm��5*��@�Z'���+�ۣ�T.���k�]�l��4=l��c�����A�����V�"�=.ytݷ���\�{d��*��V,���Щ�r_.���xN�R�7�R-@�q�U�'��5{�C���n�֌��}J
�!��A{��_�"��SO�\�$�E��Ч�t}h-ஔ��<��{��u���E������ӗ�I"1�x�k���g�e���֌UJ�>�ye,���{n��N�Aw�+[Z��=�Ɩ2��$����6���UNρ�]F�%<���w��1����|{��`���)Ѯ����{�&׸�'^��¼��q��⹫���*�=vٵ]�.���łS��4�H�Y�c�>��keA��՛F�-�.�K����pQ���yW7�c�P1�i�].�n=]ݎ�ߺ��b�c���/�����R|%� �T�V�w�~a<��������k���y���^|TK~��{���'C왎�Iu0?��3=�)���r#��k�]�h����������g�p�������ݗn�wg#�q6�`���:���AA\���wm9cW�ϓR�IM��Mg��8�D¹
��q��Xz�w���hz��=/..�{ým]��:�jw�UCn�>#�ŨN��m�+~������#��K�|���a���-����]��3� �b���8_��Bߢ��Y�ش%�+.L�t�o�v���K��㹳5��[\����~p��S��~��Yg�j��y$����K2gW��'ή�ޗ۞��߫~N)�z\>����G���l���:噽�9���\~�9�J^�s���ݨ4<�	;�D~CҠ��݄�Z�u�9��=-�Ҟ��{Aݺ>X-�`�"�aX���E��~�Y�JD�e�ZW�WW�fI{�b�:G<%l3�
��]֭=�:S�H�ì��\�-��_iv�f��&R-v�v�[�u�{2�s%;���|�g�.V'04�v�0Z���o�My�N�mmq�4�|�� 5ݻ5�겙�K��N����;!�������G�������.gF�*1Wי���Z��K>/l
>f��l5�-�/]��'X����ouF2����kn(����떪�O/���RϮ�~��{
�c��I�L��w���\��$����9��=�/ j��>TL�5M��<}��<�8j����4M���O�ZϾ��߻���o���s��Y�v|�f4.^x@*а+�Ϭ��g^��v/ppr�:�s�����.��V+���yb���g"�O��<$��+_S��s�@3�o��Uޟ�׍X�]�#ߜ�tm�ӉT��;�=�b�z`����L��:t��9�y���.D��z�3��ަ�}Nx[�/ wr�k+�e�^k�9���/K�0��w���=���>�t�j9RS����6^|�E��_���j�/9�Æ�ɩX{�w=�}�ѷw�[c�f�=*�}����>˱�Vb�~�<�g�G&-��Q8z�[<R��u�f�`�/"]�h�
�n���i�Bdm�Go@-�����I�	�Ҷuz���u2T�[.�ǎ�n��M�m��Z��Y�*�m���y���4j�M �6[�c��-����1ohi�q��� }UUcLw<�Հ���[Xי|����K���1�hr��9�]�R�6��ja�Ӝ�ݫ^��=��������O`�扝��
oå�}�t%�?�/-$o��@�&�v�.! 3*
��3:�Q[[�[���~Ε�oPazS��h2T���<_ ���ߗ�gN���=^���B����.�m�^*k^��[�[��xH+���+������z9`�����Y�z+�~�k7k�g9#8�md��|���-Ek���SR_}�E��C�X��Z1U+�J�T����ݡ��_�V���Y�`S�qK+��a͜���[���F���k�%��jޜ�ئ�	 �g�TϬ����nw���R�''��	)Um]vnOxIU��n}SK��Rρ�����)�_]6��'Ѥ�G犰�bo��C[t�}$<����`���<^Q^�~�=(�f����T���gY��zl����lq�v 3�:`j���5f�*��{��	�T�^�ޙ���bK9�ǰݺ�&Ja�/�O|/��700��܃6�i�_:��'��^�����[ya��)\܃I�Pe�uv��DYb�,S�T�J.������[m�}��b:��W-�P��UJG�����<�j{Vn���>Fvw��_������ǫ�w\"�&�γ�'�}/e���Z�k�ܣ���0�k����prE���"��C���1�Ш�5(">f��B�e���;P���}�9י�:���������zhf�T)��+�}�g�oyx{��bC��������_,שL[�8!�� �%z1)ۯ	���c}�2��S��Ә��b����go}]�n^;6;2?|�Jg�y�N�-��ߧ�Z�=����v��+K��>{�r�<��4����9��1��1N���o��4z\���uw#6�rwi�[t�.-��u1��⺽�MMV|�()�~Rw�jC����u�>�m��;90�n9w��AG��x.�t
��cɩ.d�\^����>��BB;��W���[�e�M����S�b��QX��`�R�a|-�*(�`Ɠ�pZ��}�shVd�+kks�dX���
�m	����9��3���^�˷�z�L��=S[rv6-�8m��fX�Y1w]:��3Z�Vk3�E�<\Y�lެV�S���}�|ʃ��´��_����Xs��a<�}ŋ����$�s}B�97;_=�W]��@��g��<ˮo�R��{e,����m���������f��DA�3۵큪{[�}�IK�9��}&����S����6i)������vݜ��۟'l}諽�NG�8��2ϟ}��Q��V�O�W��~��&Ve�\%��׀���ؽ�Oz�t>Ϧc�]G�tv�(��������	ؑ��������.�oRC,$�3�뼲PM�vM�}�;�����'�����4��������5.H�1J�^��upR�/�+�J��XOEz�U4:�_�ฺ�s��/ͬ��n��#=��k�B�z�~��8_��b=�mdC٠��[�|���8�/Ir���VmߧI�� g�W�)}�4w��h���y�Z]�䃇ƍcvd^�9}���g&��YAܮf�ӋC�8��w#F��9]���N��R������>N��٩���n-՞�R4J�I�ŴLY-�h�ipoG�n?Rf�4�������A�/�����{�2m�j���N	YX�*��v��x,D��Ef��K�~������3[�� J��O�؇�ſpC�l�}�_�)�{�Uu�ŧ�tfD��e�f{�z�5�}�M�+[K��G_������~�������M���"��5�W�u�|fخ���>�)g0uE*�s�pw�����p�}�y��ݑw�����9�y[��TY�+����R���4�Q����^��1��f���9��Z��K{b��1g��Y����t�{��{\�����\�h���|�8��UJ������;u�iIsX�_��~����^��Z�֡h�K�{�=Ѵ{~��v7/�9�ce��\n��r}ex�O�^OW���օ�����-:����&�w'�3�Av��گZu����`��C:�����pr�:�0�9}uU�y9P,�rK+��#�Sy�~���h���w�n�E��b�>X�1̭�j:T��W�2f*��>��J^�^�Y�}���c�m��2�u�wV�c2�^u�Y"�5�\!y&s�N��$�;6�Ļ�ĮW�l	��޲f���ƹ�����ک��s����k0��LL]�k�j�ۓ�������܁N�����!�3�wO�k�h�&o��ʽ�1��x=2�#� ��nu_�ۮt���9Z89��2��i����/-�����/��:���)T��HV�Ym�Q���>��)��#Q`����y�1z2Z���3�B#���>S��6��\�z:;ރ��E	�Om]S:&��-�����8.wgֹ�~}c��?9�w��O���Y�kGr|������ށ;��� �X��>���q}Z��Oe#������?;�<��մ!e��v;�O 2����������� fuM�ܟ�j�Q�>�e=Ȉ���>T������|d����..�~��z����+�����N�s�k]�z�ҧ��ܱ5N�W>.H�f��Ծ��֌�K /d�8���^U�s�;E���d���jjK�'���ߝ����Z1U&"7y����}rM��ë5��:w-�K�����,vMj��~���n�������܍��!u̚k{�8{����:q�;�_/.�� �Z#�4�#{���h��`iw��g�Zp0�2�qv��e^Aм��D�	óIr�;{49��ĵ� ������g6��F	y�~��5}p'�qK+����s�O8�sȾN�S��歯tĔ���' ]U,��`��1=���nv������7�y�T!2�����a����z
���N�xRUb�ye9�=}xk���F�g	(��lk�{֞�/�{w���3��N��غ��S��6�kީ�y�T�����$��{s�E|�Iy]C���j�V��R�Sr��l�^�k��Jnƿ�8ܨ�8y�}$�ϥ�L�F�bW���:�^�7�&,��Mu�֧^���ϛR�H�l0zhg����yf�-!��N���:)��W�4zW�P6��ۓR�Nu�f���;����(��L{��i
~��ٮ�={����z�謋+�0]�-����9f�Jb��4.�Z^���r�`��1g�!^�%���}�)X�hw37K���O��?r��亍^W?� z_V
���V�6.��܄�0Y�0m��Vkj���2_S�և3���r�L�v�w�!﮸`��x�j�����)�5p�8v�+����9+K�k+�L�2�wѺT��#)�x��:��Z��Y3S��O�ʄ�7��p�@;"����e]dEQ��\[���,��àH�\{[hÚ�-ԝ�Iy9vKsݵ3�6,pp�U��좲P(9�R������N*ˬ��SU�}oS�eD�E�[�Ns��׬w`��LK��`�s$g-lҤ'��J���gF���}Bg=���[��-�}��\8���w�큟��R9X�醎��I�7t:��1���]і�wf^��"��C5]�LxB��J);T!vu@���[ae�̻ᚂ]@��mm�؅dm�]�O.�����Fp��!���.�7��`'-��%\B�&��7��|x�R�qS��Efʽ�Ae���\ŷ�z���w_Mw|t͈U�p���֍J�Ǌs�vʡj��k�c���v�Ƿx!ܵ�:(%9�����@�-��ŉJ�3�u���^$STB�w�� �Y���w]:��3y�:�y��4�9>�c;��u,���n���.ݯ�qQ�׺���k��(���h�n�v-��Tλ)��g���/eK?_,wsz���.�6Ԉ�ï7K֏A���W{R��2�d�^�k�d)uɗ����wNƆ�t�wSp���t)M���.u�����K�3]!'ې��*pOB�TSilK�q�ٝ�{$M�@�����;��i7��Y���a�D)V������ÛWٻ* �R�aqӥV_V�Rt�'�ԭi��i�n�6�f�N��<�̕�HVq�VWyȱ�U:�Ve�S|��rl����*i炆3׺ì-�7wIV�|��q�Yd�i\]�X{��f�Z�t4<l��r���k��w؋=��+�f�[�VכWn�1j���a��nb3h:�6S���k�e���6�Fb<sU�zcrl�g9:�..V�z�������x�K�㔱Vif��&�)e�CN}m	V�\gI���g>{3o�Kv�oNK�� Fi
���"��b��
坖r˨l'��6�9|�5wݥ�EBZ����u��:��V��n��>���L`.��ٸ�#�ha��*�;+A��r�>����ஹλe])��)]j��!��X�a��)}u����04D�%Y���1r�Y�x�����+�ų�~�����qÌwR �[yW�Xx5��vA,���=;x�b�B�� ݗ�k����_v�� �� ��+4���a�&b�v/
��蔟C}Q�]�gQFڣ��V�Yo��x��]�浜>��}������;:^��]7��)���8�R�e�:���L����PL`��\����� n��<��d�V,���_��c�m%fP�.�ъĮvMTÙ8EH�����ٌ��r({9a��@9��S/5f��,�)P�VU�t��Y�>���}���������h�1�������-J�h����+Ƣ�c@��/(����m�Er�C��X79�̨'u\�h����LX��;����r+�rܹ˔�y׋��ڊ��]ѭ�swv�&Ň:������\��r�;��1;�%�Z�q�s�w;;�˓����]��݅�&9�����wA�tX�v����+��w�nsu݊��2���ǌ�ǘ�Fx�u�L;�4\���!ٮ\���N�;��tܹ]]�j�]�k�swqk��9��̀ۛ��;�p���wIλ������W���.�\���$��n^v.��s�tGwW-��G]@EB�Q&��ma��ok������wF�0N��[�){�u4+��ih�j�뜟M�\ u�y�y�@�r��6Z�2t���S�����}H��=�{F%WeO����7k�fW�Ғ�X|�ͯy
�XQ$�>�p ڻ��;��:��z�Q.�{'WuL�p�+���xz�]Nj����-�X9�55X�(4��N�Z@A;����a��op�Nؽ���5���@�,_�P�����W�n��n�Sp^�ƇLo&����l<�t�<j�]�+|��E���.�;�N��W������ԕ3��ނ_'��*�*N߫�Y���;8�}eP-�Ǳc
{����<�,�����-��J6�ox)*�Q�5�}xZ0bz�o����ś��G�����:5oM���&�^�1���U����b����̉�G�s�J���O�{T�-�����;�l=&c�K�Y�����H��������PF�����)��x��8ܬ�}��I<--��a/�A��1�RJ��}����=�ܖ-}�tm
6��5�WVN^��T��`&�X�Қ�]Wj�S黵g��+i5+B��c��j�zk+s�Ք%� ��+�w8�?��`�o',ﺦ_K��-�{�����B������Q~��<����D� H[w�q^~��r�x�Դ$������{b��Uz>�1)U�n���Y󽖀���Q��k�i�Z��Ǵm�1w|�䗌zk4��OJ8��O��A��}+�6���.yd�3tP��k�qǪ�ޙ�J]�$���_`���M���p��pL�[��f��gֹ��*�����?.�xg���y,&���G�PL�i��!��.��y�"M�\yҵ.�������4��!��w��#��=�������P�}XqmZ���#TS]ڃ~.y���n��)�=�J�u���~�:w_�'���0W��U�s
�2�y@׽�^G�y�}���F�	���9�{if�T�h�����պVQ|�1�����P����Z��7Ҝ��I��&uy��4b�U�ʭ���S�$�0�n�%[�Ø}B�s�A�;u]x����!�ڊ�֧����A˕��ΩQM�Ryt_l�$\�푣a���\���s2*�.I��w��rt\24%k��vq���8����!;�u4�}:F��d�dҭ\:e�ܛ�n��ӈ��UULk*R�����u�\��ҕ�b���h�K���OE{�Ϛ�n�3�S��?���� ��iNbz鿕��윏g�d���md��gvݶ�-�=���O����"�Q�I��g]6�gb�}����}�TpS�X���Q�.g
Yx��x�M���
~�5{�Aq�F�m�k/�z�4�W�=�붣��&g�Ge���1W=0s�w�:���t���ޑ���gs��$��1T��������;�x������t9�oK���OD&ך��ϒ3ͬ��RT</���jl�F��8�{,/7�������Ag7!��o��:��|�Mm���9��zhf��h�=�N�G���|����6�[�E�y-�/7ţ��9�w��h�g�NΛR�2,Y���}e�G�i�7��s>��j��|W�������u��!?u�lo�V����tWH� =1�|�h�)���y����;��V���`�CN[�R�a��BT��es�m�R��u�ṇ�������C�� c6K�Y�+{R��.�����Ŏ����gu7���Е�X�Ɋ�f�����ri����{1�������^iEWE넧�����r�4������~��9�i+}�I��؏B1]�8��I�}%�(���u�N���\�{}OF�;�����&6�Q�O�諾V��rE/7��.�m,�K /W� ��sF#~��I/����A��k"�ŋ���d�h����ZSև'�j��q�:#���Wyd��{l�`O�qHt���<�ێ$
�0�Sr�4�[5�a�nf9K�J�{�|�����Q%{��zk;�j��`H�fg;�h�{���V�2���^���^�������7��s^��w}�c$F��̩�ԓ�w���w�N��������v
b�������������C:�Q�}��<���{q-�K��U)���WCۮ��NSW�7�S�6��v-��W�N7)����g�O�[&^|+��Me�Z�gF���3Q3~��L���U�3��؁ �÷:�
t>���6���W���]��=@�0�Y��P���b��lw^���1>&DS�57ϙ�w[��e��]��p��k�3��k�������A��{v�]�W����l�ﾭl����ʫ���
r����s��~��/�T�����;�3�]����?7F�(�Q6�@��'`��<�o�sVu�uN����E~˶0�$���f߽V�VOC}����H�VD=�����^s����Y��+}幨$�Ҳ9;��_`����b���~�v[����^�V{��fdɛ3[axΧ��k��������zMg���i�6Ù��;��R�Wt7��v�Z�S���%�Ӻ�d�{�Ck*�j�:�r����E2���K>�55\�(4��N򏐽�*�����罎v��^b�qWأ��e�@��/ɨu�~���
��4�)'w=V�7}9��rM�s>2��h�Z��cڡ���D)opl�������#h�<������R�����y���]��ոb�/�җ����i׺tV��/:���[������Y(OP�"d�f�����1A��I�ǌf�� ۛW��O�%`++�r�ۦ��#h���\���	'�wJ,r�y��N����S95�k���RAY�;�O��s��7r�FÍ��6c��_S�NTyyR��e���hY�m��W^��g��U��K��ɗ��[�A2�/e��е��nv�:5�Wzr;%�>�i��&�y����y��LL������j�)��\�-�E��=��'C�v�GyHx�L!;ǝ1��[���oٟc�r�ڦ;v����r�F�,�wL^�W��wغm��� Z{V	/e���
��υ��x-��~�/W�MKŔM��Ƕw��%��F^����9�Ш�/H�c��y5���S�.�]�Wf?W�,�0�Y�&Z�Q@9���~���Y
��Ů��^V��󵾬�ri�=��zu��f��^p3�H+���-~�Y��6�y������%w���cK���E�כ�;���3Ю�xo�����=�K	�͝�s�n�(߼g�M�۵�|�&69��j�g���S3��ޞ?K�԰�Qy�<�X��3�^���z���-���*�v�d;ы6N[�R�dr�gzӀ2�<F��⪲Z���+4Ž�-)�.u
�O,�9S~�й�:usvV'��"�K{���x{)nꃖ�pNA}���2Wp|��lU�7`�P���i�s��7+8	}|M!�y��k�����9iv��`�)`�����y����]���!�u�����ߢ��~O���������lE�.dX5VƑML��=�H+��O����f���y���ͤ���>x���mT�>�q���i1�L'xZ���c<��m�AqE��`q��UK��Q<<���ʎ�缽S�����L��)��7GA'l�?g�9�/��g��� S���o�t��,^��2ʆ����V��~�=S�'#ʷ���n�̛��y��aʯ_cpv�/��}�c*6i?x��ih�^ȱ,�[���~��:�\� �Ǚ/�1���G�6.�����y�\7N��1&aOot��U�����wBH�*�x]��t�
?R���~�'iՑ�3����������eϣQ�*���B�<�%���;XS�vU�=�ºu�Թ]%���t5�����i�/��7n�pь9�ŗt��m��x�o+O��c�ȶ��K�'9������O+�M)��B��%YS;����+F�p�n��m�D���w��ƻ���=D3�A���}Ң�$�X�u��ƻ�;T[�u�T�J)S���bK�Rot�ϛr������qtF����v�}]�CYT�>�ywm�׃�X�:6�ָ�$���V����Ǯ�zAɛtk�{`6�<�.k�u��u�&u�����b߹�����%H��#ܽ~�������&z84�}�)]lC������kT�#��m���I,���-l&�t�w^��{�w����ҕm�Q�Fg5����׆S՞����#��7��S�;�Ƃ��s�/j��~�����UB��K�	�He��޼��V'/�뵎`�j���rE����9�t}j�vljbޤ��U�i�sޔTϭ�Ϯ��︱cSR_|2H�≝W�흃S3�w7���~x���w�k]Z��)`���j
M�y�l�[�W-p<�V�� b~{KR��3UJ�>�&i�Y��.��������z+��E}�fG+�����X���6����J�/�K�"�mD���o��*��G>���M-up���+Y+H-?���V�*��n��Xq��O�N����`CWWtJC@�Ť��8�
b�t2̕5�^�ꨭ��Wp.��VUo����>�c�W��'^�*�e8�~~�Þvu"�'7���v��5�W{'C�&c{S���vG����~�u���Y��RBef^��Qާ��ؙ��I�T�{�fK��/�Aֵ:����jL��ү�Ϥ{MX�����z!���γ�'�K�y���s$��%��Z��.�5�}��yo�y�X�y�j^IM=3�ɘ�f��G$�w�9���sV��φ4{-5޴����篥ws^��&h��=�R!�W���w:]��ůԩL��+"�ֻ��KϹ�_��Z����lKym��7��bސC���/��A��)~B��\�5�,=��VNWU�J�nj�+�y����'���׶�eD�e]���y�E5�wq\������v�ZqM�����g�;��ű6/�x6
�*:˼���6J׺��}�����T4�F�0>�q&J��~+,�>\_U�]ܮ�	�/�E����Ñ_��%�J�ynF�@qbk�0�eF ��ʸ9[M�\�g���5gu:H;���
[�����\-�߭W^3..�_b�{��n]r�m��L���K>���g���;Ϣ���KP/�+�{��_���I����&m>��}G�>�h���ŏ&���r�8��m/0��s��<�t}kF*�`�y��b�l'��Z\�N�����S}T�J��:J�ܓ��-�~]n�U�|��e*�=��ڀ�AFgt�ܾH�5��s�QԳT'��ꞑ�N�M�/�v�%�ڢJ�ivH��SKw��5G�/�{H^펾���:5oM��&I��1�Πg��=@f]�{�v�~�Pv@݉�/q��;iN�[�=���Y��z�Q���uΞp�:��^�C^Yn�V �����M��lv���=�]܍�W�<3���>S��\<���M��/]�/ WM`��)ďd�_��<�Orx{.��|�WmS��G-A_��
��Lr�*:mO��o�j~<���z,�|��<Z�X}H�����}v���gq*��<j���S���;=6��&`��v�ʒ\�C�R�{���{;}A���=%s|��Gk�̫�f��k$���'^vN�c�ʹ�I�I(���t���ŋW�cimg�tc�؉��U�j�]$ǲ�v�&я�X��G�%�jF���6�v��^�jV��z��b���e!��,��(���ᷢ����]�7�{��/�Y�on�\L
U���J7֧&q�o���� sI��C}Om>�Yt�5e�MK��j��1�k7tZ�:pŊ; �����a /9w�w8A�e���9�L�/B���b;�É����E>OI�GO_]SU�ݴք7Q�kKԹyw5�����X��껮�p��W"��M��۾ �,\�^�jS�TK�%�t��6@�K�d�Z.0��=�BvWm
�Z8�gI7��U+�]����5���5[WR��6�*���t3R���8`e'�iA'L"Ɏ!�u��`��U��Y�h(!�դӡn�(����n���W>�/)�M-���o��R� /C��S����q�iv\E�[yi�.��VIu�k�l�H��ѩ3p�^�K���{���C�+�g��o����^������>��C�S��jr3�=w;�5� 1-���|��`	�$�0]_4�nq�,Y�zT�y�����s�*8u�Z�z�W{Ɖ��eB(�E����oe>õ��\���r��%78��rr����]�\s�_Fv�uk;V�Nb�Zج��"�`�A���M�m�}�Z��#˶�T*3�c�3r{F�����8G�O�����$���k�Gw7��}��q��,���Ы��m������^@n���2-G�ɫ�wfʻw��WK�:�&_e���uа��4h@�#�B6�@R�n֜Y�[�,Z��=�ov�zgE9�x���R�[��[׎��[�8h�q�#2��9�3;hG�թU���FFS���;x~%���]|����.�Ɍ ���m�h��C�/��;.�v�ǰ;��NX�2[e�6���{7�1v�N�k������Ǽz�7S��=�jNn�7���ų ���9n��;�)�hv:�������!C�6S�5��暡w����rs ��/͕9��zWe��z�K3ITQ�$���Z���r�.$�c]fZ���q�둰5r�|�]$j��u>C���NB���6g-��_��..m��k�eN���[�:uq���Ib1���}�"ۺ�Em���:G]oUԢ)-������<�tdm[�
9�jxe��ح�W�`�;Jަ�=����TnЫgk��ᣇ57�܈�ݸ(5������_b�0��򭫢�캘�tŐ*C���Y@k�9��j:��n'$k䶺У�*ע="��hF�/�zO^��	;�� ��]ܲk��ݖJ䆝q���tN:u��;��c�:�<�^;��uԹ۹���<��u�y��us��]�^w�Ν��s���wm��;���͋��r�vŎ�r���u�s��˛��n��Z)ӭ�tf��Kp��w]���ss��nl����wN]ӷ:wq�',WI�'v�����7s�s������Yw]�W2%\�wv4[�]�nq�\�ؤҮ�˕���K�.kwucEt�k�d�틎�69��Gu����W)ݬ�.j�"��9�\w�]�Hh��f��ƒ��ݩ�wvEw;](��4P`��W0��+'wX�Qi7+�.��5�a�+�6+��ڹF���?����_��hY��uF�{�0C�%�MUrldN��͆4ý��u8�ټ�;T�G����hˬ�y;��{��k��i�HV|��m�(9���c�`�q�پ�l�ך���c���4�[s�X��hp3�A^P�}�8_ޛEk�]�(�v��:zʗ��������Y�������]������{�ɳ$lՒ����ۻp9U��lC�󕜭.�G_���y�5Ν��(�ʥE��*��Kr�^N\.ѻq\�;�{}��,���%�3p�3���r�CN�Wܧ���3U��x�ns�����n{�uz&�����}G�x˙��rǧ-z&4�"�3{��<����%��`赧2�6�ur�7�.�=�*��{P�8��Ԗ��Db�A�,q��UJ�>)��R�'��N�����Y��1xZxɽ���G9ɱ�C�xKN����gn�9Uz�>����ye)�tڵ&�#��N��=XM��]�wY�X��$�hr4�pJ�ئ�Th5~^طަ]36�r�Q,�&b�ЬW�]ǳι���o�����;{�e���S��f^�n�͓OQ�"��W\�R_^�59P#����_4��4�0O���Z/e�j�vJo�<�v��'/))O��
�Ȧy��ژ�;>��7�S����ixp��.�c"�v	�+��wގX�τ�w��3�:ϩ�b�����a:�[Y�_lr�&K�w:n�wr�o{���8�T�L��H�T�J+�dm�u'r�4��1���V5x�5��J�Jse�e�F�μ�pŖf�=k��ӥ'���F*��ދ�-N�%�E�me�nTߡ��~g����%ӭ���O׵�ڜ��z6�faw4�=z_����约�yy�rH=:V��x����]�ǯr88Zf�ګ�:[�<��/3�>Y�:xӞ��핺����x��MΎ��N�ݕ���d�`Pi�AK¶!��{;-�vr�Y���.���qEe�U�S��yH=K�~��ʞQ�E�FgTM�]��xT���md��i;'k��ۓ��@��\��"]�;��'���f췍W����ey*ḋ(�(:�M6TB͝��m�x����x5�9���z���ib����@Һ�[)e�B�ȕu'l�͝��rs3�e����ߖ��hTS��h�hY�)k.�jݘ���RU��z8��
��GՕ�H�yc���-�3ԽQg0F����䋾���9!�����{�k�o������9Z�G"�o])k-���,����I�QD.w%��ř��=���{�n*��'�b�l'Ԑ�y���3x�iUY��sW8<`�kK�z9=����j�Y��=[�f&���(.S}/w��w�4o��($��=O�9?C�!^��?��|�
����^x狞�W��,;۞����=�^~؟F�諽����f7�T�1�:��h��c^�rQ�����>P�z��������K0z#����#�VɃ=83�����'�wނ���_9�SW�����CM��I;垗����Y(怺�s���^估߯({<�����m�hIH�AÏX��o�ŌR
�1jC��s]c����Y�e���X����{vL���b�f��`�}s8����Kn��®�F��{�Dy
�Q����P�2��㦮��R���FIWu��l���}�]�,�kpM�^�&ZU�>;9#�q�b=�e�(��0YӻC��ȵ��OV�|��HN�ג���皪up�#��zQϜ��Y��=2[�dY^�Wi{�²[D=<�P��:�x�o�R���/��}���9}��s��<�
�xlR����5�� ����wۚ����O�U��|���䰟K���k�	��
��ȡ6d�~^�9�����=���-�Q��<�/��7��sˢ\/�c;�˭б2�=�+	���y�f�x��������sSU�\PS��ۃl�V�j�Zc84�m���]b�_�׃����;��רּ��,r�x��z����y�!p_g�`�۞���Zъ�X-
��f"�w�Y;�jfI6r=��gb�x�c})��$[��������R��v���Z��ʷ3��}R����}q�*k�,��B쿡h[P�-�ixm���}�)Kl��F�n6��/�=���p��(j'篯s��:5�E]윏d� ��L�~��+,^V��֫y�v�2ެg�r1�I+���w{^�e�}��9O)�L���:���/ �8l缳��_x0�.<	�F�r>���t}vw�X�o�1�Rڇt iH`BwUe*dz�ݮ�뮆򰥕3��ǚي�}���p��U{�V�#�s�(z�X��xio��/psާ�,.���H�瘨��r3:�K/�;<�������N7{;�=�N��9*k�ײ��}ՎOr_��v�Xhw�5�w(w��<��^�j_X��\�s:���K�"�������<r�O�#��h�y-�������mݯO!2�޻����C3��^ܢ�>��ǰ�Y�*�;��s'�_�����=�>�z�}x�Je���g�W��/�z�u�����k�I��,/U�{Ui=��[�^o��GO.-��e�ú������)>�}ْ
=�����uֵ�Ws�ذ[���ǝ>Իc���m�#.\�)�^!>+�@������}��#�*��8�'�&,i��B�EC~��)�����ƫ�)�^�/%���m��9aͬ�!_L�"�;���v5��z�]���e��J���Ɛ�gNru^�& ��4�Рn�4
s���99̇37��cE�|/�����;i;�.1ΞXT[9��8њ��U��f�fR��|�t�w^�*=��б'Hqqc���x]{���@ʭl �m�����T���rE/7��t}k~ͤ��{`7�'���~�I�mY�o{��ϙ�/��,_ڝIz�-��]�ϹvJ��u���ݳ���﫷�`�d���\.�z�{�������OS�ty���D~�����b�SҒ�u�¢x,���S^鰭I�(#��A���b��v=�_!6˧�I���I�;O�:�ϩ�To>���l�#����q� i�5Dߎ��k��Xz�`y���^}>s!rVU[�3}��U�X	�{���}�����F��!�_$��*�< �2�m�C��yɼ��>ƒ��h"���TV5x�MG**�CΞ�2_}�*k��B��ھ��X� n�'s�j���r������ە6=o�h]e��'����)��4-�^���m1ro�ol�wm�ל�������5��w'vAOK����2�I�K0���=�>���G�ot��ֵA.��Y����*u+����x��x;���:�n���sz$�EQ��S��y}}�<�������^��>�{��G�n�`�Ϗ��g�G�M�5��'�ll�zZ��v�����}�h�d�um~�l��~�]� �ݟ[��=���Um��ʼ�{����|��ٌ�~r���y����wΔ��]b�|�3;�ɷ�{۞r�����9�wo��
h�(�Ộ�:R��K����8���ks��;������|7����8�W��qzE���3���;i�Mw����zqz�uNn���IL���9���ς���$��sȬ9ѻ\c�F�̼�R�x����t}�ז���gەg����.���m��Ya����N
�����}k~�T����1e��qK+�f"G]����d��mh[�|������g��O,���N��3��w��p��ʕ��Y{лmh�`���} ���`��*��t�g�v�W��:z�yW��;���k�'ѮW{'C�3ߪq���72ٚ�k)�������f^�}��쭠�d	뗭ze�y�j=���t	�ۏ��{[�6���)m��`�=`t�m2v��]���c�ռ��u��7�,]~(-Ί�����|�&��0��k.��}��V8^N�Ї7L.ӹ�lfR/2rήi��)	��ت��A.�
��!-�P��UJp�w����ծ�ؽ�T�ٶk���z������=���xq���J�U��o�oG[��c�X�ǂ	{/ڼ�YCƟ��u�Z^��귺O�����v��[5��S�B����Û)����X+�O�}nu����z�9��N�1"�YVVb�s����͊Q�$��7����jl���z6�}>�>���]^�C��y9'L�}}���x��pC��`r����AJ�[�yLL�w�x���q���VH��<��?�ף���p)��-Osv��h(S���8t�鳻Zl�j�z�k��]�����~����K�P��T��oN�l�����3!誅�5��nR�`�j��qA����oY=s��^��^�p׹��9'|�tՇ4\��[t	]
^YJ\�P�R���-T=��~e���˨ix���t�HK46�Pf�S�Z-�I�d��+5�]♵��5r5�����>yJ�����P[��鑮��x*B�3Z����7��������:��v�2�g5C[�:��r���z���1]�A�z�߷�s�Ч���Z�^-]<�K4�
������f���A⽀q������$Z.8��[\��;.�R����j�j~�Öak\����m����}��=�G<�ȅm�Oz��y���X��o ����P�S������:5�*�d�{��걎T뉠��_���� �N�>�o�({��Ͻ��}|��{�m��n],ķ9���u$��ܾr��������Sp;f���qO_-U���g�v)�C�'}/e�-k�<W���%�V���2>�� ����dj^}$U6�4|�se`w��SC�����Jw��܂xM����Ϲ�y߮�nQϜ��@����a&B�ѹ�&��V��'C��v�s�>�x�%2�\�W�/��P�~�s��+�B�W@h���(����"�+��Y��
������o���]n��ޱ5�1�`�l�;k;
˘īF��r���v)\���F���gtP3�a�2A3�V.˭e������v���s5���o'��JS�bo��h{B��l-�ojқ�g%����}c�5���8!幣�X�(�ۜ&�.��\ir��Y�w�d�?����B��|d-'Ɣ�n_�U�y�I�Xe�ǡp�.�vڦ9�b}��٢�<����xdL�4vt+�ʭ7G�<[~�ÂVTS��Q�h/)�
�ʄ�U5ȁ�Ju�q���b��7�v��>��>>ɜ�tjJy�U�=w囝�:6]��8Gzpp�����0
t��w���;�b�5���g	����٘�Sa�u4�= ��8�����l�}�T����+��e:���19>��P�K�7��7�r){���]aqgI.���Fz����7UK�ԄG�w�#\Kgr���6���cEkclwllt8�����AdeK6�P1��}P���n*g�3��*'�����Bٟ
R����>����g�ͺ#�n�Hۆ��y3��R �5'�L�D)���r���*�������D��M��-�g!L�=�'#O\=w#]M#Z�P�T�{�=0��U���+=+�c�ժ#�޵Dq�8�c	��Q�8pQÛv���r�mua WQ�7����΃[�B�`�Q7x7b(-YFƹ)�2U����Ԭ��ǃ��ir���e�̼�',��o��lӑh�39�� �-��Ri�L�B�.5#������*d]�X4M(�,T�6Z����F�.z0�ÎQ&#�����/��چmd�ٳDvT�vr��ө���=�ıH�#���P�tY* �tԔDMW(r\]�KQ�3w�]G+O�,��ѡJ�]+��|'�kC���!�-=��ۣ4��4�J�7Zkr_Q�U	*]1�S����o(�j4p�i^u��݄�\�2\"�uq�-���ެ�E�K'I�l��ݳ ��W�V�;H�����)8���2* -
X����i��;kr�-��ZF`�N'���*�΁���7C��|{�e2�%��j)��3���s6]�Paz�܊�9vK�|���p]��6d����!ՍB�+nWB�nH,�nQx���e�xj�G9���m��H���ݬ�$)�O.N������z�����L�x�>��qn�J��c[�j�گ�AM��m�n�.��s�U{���wkeX�=1�乻���mG�u��B���bé0������cC��y:�;���3ek��xf���soy]q�q�ez��L��:M<�!�:'^H�W7.���n�.�cuK�X�wj��N���o���x�Q�C*��l#{\țy�,�ǘ=6ؕ}�Y�0{�9l�c�5�,|�su�uq�`���9Na��k�(��1�}y}���-�u���w]����Jw(�o[�ӡ�Át��Ғ���7�6�r-�q�v	����#M�L�۠��h�}tlU�i�zl}x�\ݭ�L\��Ī�x��U �cz�b�
�͝���N;ó>�+Es=���N���Cr�1A��t/Q���4�Q�EA�U(��)���S�7\�l)�C�*�ѭӏz�d�rT�w�Er���oX���n��|��q���e`=�#Mⵕ���9�8�Ku+���qxx�7w�Һ ]M�ڻ�yCipY�6��Mk+�yН�Ar����7p�}[�;ļ5V�`�)�lء���{�;�kƹupO�ǚr��v���� IͿ �חh�zȥ��b9��|�q�w2r�i�̦{��VS�{%�����3:�sV+�P�"��Mrm ���_u�;}�o��#Q޴��Nm,��q�φ��ٹi��w׽V�n��wj5Qbn8�U��2��P��*��On�ϲ�Y�`ė����ؐ�� ���������D��{9�tN�g�87��(\u$��n,X򎡩E8w-S��b�v�U�Y���{(>��Ni�ⷶ���aR2v`�tw��������.�20��}��
��O�[Y�/#�=�k54Aeii�4v�]1&���n�s�	�0:Ը�T�W�@~"�sn�IF"���M$.\Ӻ�F��rط#��K�5��;��7��W+��I��r��܍�\�L& 6��b,�wwN`�v�s�s\�;�(���Q�9u܌��U�wwsF��Au������5Nrgs��r���"�M�r�j�5r�2�*:c����ƒst�ȆXɷwc2b"��%";�Id�n��6��ܮܹ���]��wn뙎h�8Qs��]wp�n��ۑ�a�]�%�[���ur$����X���wsr.\�Ws���F��JKer��tȈ�tH�&�5�r����6.�Τ*wp��\,ZIGuҊ�)!��5����������?V�+�։���ۓ}�G>M��R������}*u���<�q�F�гw}N��>Hia����q\���ʼ�GH�~ٱP���if�IN�.w�wv�32�I!z�z7�y"�9��������dк��wc��R/S9}e��3����l
O�>�=8}��y�%�}�l�E��=�2"�ޥF�횽�ou�B����K�e��k'k�<|g�[}3���q@r��)���f���,�b���g�����=�m���;e��i�y=ӝ���t(����w�x�ho�]@�u�g� ���.w������ݱf�k�m�F��WDՙQ�����@98�P��BwC�ΆLߜ�x�Kt/}YLi���L0"��%7y��4ΓE����W�;��4�cq\�F��'�~��iȓ�����Y�6.B۹[W�Z�qDM?��8R�N��-��}�\�Jw�s���>�a��{�^2�`�dEG�H7���V�צ�Q;��ʁ;���VMi�� >�@nr�t�w�Sn{b�`���V���v��c�I]�v]�L�'���0�џT+��U�─���1��Pʹ��o`�x��Vχmd��&p zF���\�v�9aCb8�}�C2�`�+�����q�w���o�1>w��m����CU����VsBٺ�=\~�X�.��-�(9������)}��88�����}�-�/� �y�T3RB�=�ǭ�w�W-�PPD��[[&>���o�ܺ��t�����;a�[|-5�C��'��J�L,���7TF�fxu}\h��m�ڝ�.%���4栠����E<~�O�)�c�V��=;%#��ޙ�T+��R����O�t>{�;�6�Y�f��K��H���#�C+�!�J>�{��kYyӂQP ��+@i��g�)�-�L����[���uzb�e�9h��p��w����>���u�R0��K#�w��GfnV�+}�{D�)���@�.yt���9߃ڴ�R�Cu���N�����ɻq c�o8Do�u�2t���H���-A���rQɫA�<K���x�!�_t�uNµ�d�����dU�����$�>$x��to�+�kf9�3^�s��ףnv�5�ne�/���ؖ ��ցI�o�U��.#�K鿏��^�%3�k&�<�{zkyw�q�#����7��+�7��2nt�|�P��W:��NA�c���{��է9�m`�8�{����b���Q�yp��W�v���F9P�����t0ؿ��������?,.��ƭ�G�/6�,���j��A��%�d�k���a��lk2�u��5�"�����rʕ���]�Je�C���Э�s��c���u��A2Cj�6�ܷ�wse�0�'���Z�M�o�['.�P.�Vȵur��G�H��xuM(\y��������''��;��.q����^�Γ�<F��3�u>����s��,׹��IY�<�����ʼ�]�]K�ZrIݳ0���a�VS�:��H9oֆuR��%O����[6̈́�v/v
p:��->���ۡ�Γ��3�q�Zo�)��(|�DOx�:��z�a�{Р����r�.����;��֫h�,�%d�a�����˪�)���N���Gl���*����w�r3���#��=���B�֫h�$�%t	��1^��u҅�u�G{Ǵ[�S���Ag��T
�VQtr!�l��P��V�^��r�H=	�ˋ�E��M������|$��R�N,�
�y�2<���?Qg�6��Mk0��V� ����iz���˛.�O��	�"�����x�f��;ё������>ڍ�|�["������\&˄�����p�4)���B�K��_�hQ���*�R��>�~^>���F�x@�<oX��L�{��xx��z�F���Ы�N�\�B ��3*�CҼ]d	���M����;�-,X�L|����
;�,��*��|߲���~b��}�������oQ��:��ŗ�nf�flX�xAj����
x�6&|�>��:8���#���S+:-չZiD�N�,�nv�zҼ�.�i�4(���:Ύ���E׻�{��l���l��ι�h7�n���f��URP��+���=!:�X�$�ze��:�'��֚`����r�tm�|K9gY-	��d��)ѿ�d��|�Tqݧoo�$�;i����֗�<�BIu�I:2y9p<�*���:@��A(ߪz[b��[��O�h�%���\	����z2��5�Ϊ����/�:
f�`�1��kMׅ�:+��3��e��p�m@��pq��W�o�������?E��[�h�����3�=.6˹}�W��W1�\7V:}-��2�Z�}D���pwj�S�!i8v4�v������:����)�|�q�T�N|�1���uLO�5�4Zy[Gq��>>%��;:�Uiw�?o�68��~3��I6Γ����}P�
���3�N��w1���k5��O�-��I�u�'"��u���ͭ�*}GD�O�J�#J��\��$|�����F.5���s��[1���IQ�wΧ:�ޜtNۈ3� Ζ.*eq��R덚�*�79lVCt��u����i���Fbs�wU���1�f�8
r�8V�J�'��o>�L��D�P���U��R����h��or�v���ݳVES#r�X<��Xƫ���J��G���a�U��zE	��t����=���;��#R�45J�Y�{n0i��/�a]�4j����Ϟ��n��_�;�9x��a��RS=�ꥎJ�B�y����[;����h�]^�c���TT�=n���[\eJ6�U�@���Q���S<9���Q12lK���������A�/�_9ϱ��~7�ީp��>�%Z�)�>��f}��+��V���\UK�7��[qG�w�L�=�7'O[�r6�գV�P�n�TL��բ���̆�_Z���>�s%
�k;���t���=i�3�&�m�O��wlиUU(߫��8oǪ,����G���:`s����@,ugz�+�]l!�_Ye�����F�0_��-�iS�1��W�����u�5SN�ǦH]D\y���+�j�eQ��"T�3)|$���˲���8��ĺ�/-tr+|�e4rN2�W,�F㌒����QQ+պr(�v�aa��Ǟ�|o���Ӟ������E��������q��9������l��R�p�����H����(�ٔ�m��[T^�ˏgr��jt���	�D't=s��7y����h�Т}��P����:��,��+)j����Ne��{ev.�w��TJxt^m{~yB����ֈHr���/�Q�
�z!Ud�~�8<���^����3sg9W�j�9�k�&U�Z������ �'�+ޙ �Z"t��ͼD�`�[�^�h�M�~�"���S�N��O�����Ω��	8�g5�1=���௟�i���I�٘�2OG���:����eS����N*r����d��l�2߮�Ur���ni�v���1=�g��z�*�{�U�wR����g�fT	�(\Ed֛�R��@g*�F�>y �mϽ{��;{*58�NE�q�LkYUǬ�=�f�3�.g��J@]{T�ҨO�����nFs�變�}�qn�]����o�k*�Q�'Ǥ�4g�ї����N��a�@8�̻G6�	��A8uc<G���}9MS�+o������'��T+�y��ޡ~�[�؏�炿el�芜��Gd�5q�_�9r^8�%\=��g|=8%�P@��f�z���>�柀��؊�m�B�Z*������Z�q�}'O����;�F����δ�<}{j��Oe�.t��2�L�<y�ׁC�μ-�pe�l7^�1ֆ���t5"�@އ~q6UR��*h�|D�@��E�ZZ��;�!��V���ߚu�|~ȳԵgC�çyԠh���Ή��Ǭ$�x�ʂ�e��C��'qsx�21w?{w˽ꎽ���+���cu�},#��^�^����B`)�"�wlnN�����C��3��˫ج���{]0�F�0����ѥ��Y�$w/���ox��O�Ρ��Ĥ�M׀�u�"�US���$� �.�DQ^;W�	�S�-l�#ע���z8�Φ�K�q�ۣi��^|�0��l'����V:����G����S��,�A;��5��B�-�/���sc����Ft�L���@y�#T6�Ά�\��9�c���j��W[�=\ww�I�v:N��;��?�V���˅��c�8�'@ﾄ�ߝ6���2"�h�J|��M��X�S��w?0����x:�˼g��ddjt9�?M3\�im;^�U����2��jI;���9��)��E)�we 7-���Z	�"�LhQ뾺�y�9{"�vl��dv�W�����?{��n�x��sk�ڷX?h��Y��6]kS�5}}�s����|����C�tǗKy:=�5��q�V�셕��m�vYZ���|s��4/���{��M��\\G���*�g�$}��ǽ���_�Nq�\I=�C�wto�����^���'�ͭ���)��#�ޙg�)�������7-������6�=�H��Sgq@�jS��ٻu�m��`.�.9r!9X�9`���)N>�ޮ�8�"Ww�(�xf����9�%2���ҕ���|7z��h�������v���fW;����1ԭ�GJ��.�uyԳ�A´Qw�_Φ�}�[�SV:��;�0�m��ɼ����ޛ�A�p	Qb�]p��|�MW���4yÔ1|�E�[j��s��=w�Kz���6m�0�\�ǉ.�3� w,�H�T�x�f��;ё����ᑃ���^�J�G���Eqׄ�j�C���x�f=JT|}<��M{���ΪC{�;�	�^����ׇ��z�F��B������� x���J�ucV���]�+�yj�v⨽H�+I�G!��g~s��nw�ͳ[�(t��|H��t�������g��=碝N�ѹ �s�f��[��|K+�3����h�u��p�)ў������=³}�HD{�������S�j�V���u����&ӗ� *����=�����}Q�<��8��bH�)ɸ��wX�a����z2��5q�����3��мN�����==v�˯C��@�hI\N�m@�,�'��/h��
��鿨�/��4V��{,��n
�8����n�z�M�Fn1Յ>��9��绔3>}D���pwj�>���(��t�rL�RQ��vG!�fvE|��m�YZ+ms+�Y-[w��v�㖎l�QK�v��!��+Ge�.��:��p�n鑫�@n�<Ġ������B�'sG��˰�G�37(䮓���mv��]�E�_P���S�ܲ`�����}���FuzR���{lb���r9S�G�S�{x��8�����闆���N�tux�Y�֎�6���zOҠNr뇊���2%:�8�To�լ�){S���||��w��ܩX����
���	�u*���!t�F�V�p+����{a�\o�;�a���C���y�ⷔ�U�˭.,�>ve��|X�����HG�6h>�Ү ���Y�6z2��M/l`[�g�{����W�s�G%�L�Y�OW�a�����7U,rWR]��;c������$:��<��	���;A����ne�U|f=K�te#T�e�j�.`"���x�w�n%�V��5!������=ꑭ�0��p��K��/ ���T�+�����q�ki�nF��N��6R/�ǷR���B��{�[��������Z5i�	f�PG�-LlL�N=��J{/���4�؝�3T�L���]�Jv��oԑNg�M��'����3jqݺ=�]���m.t��=� {O���)�;��՝됯�[d9}e��3���e��Q�#v���{��.��I͜
���1�Zѹ;���,`#h��RC;oZ��4iE�y��)����fS7��y����f�y�4@n�:��к��D�r���{W�h��pu�p��<ᬩ��(�����m#]Pz�]7��oՋ����������|�����4#�����5��ꐇw��=L]#��t��-���ե�"�_����y�ƁP�e�����q�_>���;�b�gj�j������7)�R���=U�B�e�8������ ��`i|��8���l����񳳁_��t�G��-@l��xr���$��5e��5��>�+�9��M�;�'�	�_:3w�@#�{}-H�ӹ7�v����M[��]\6K�p��Z5����t�zc�8�g\���?^��4Ϸ��ڥ��_�ֽ��k�ST���2�F�b�(踧,���e9o�t�+�ҝ�ni�vk�%D���3���|�;����=ۯų���N�B�&�� >�@_�x�:�<��ɹŌ�K�.��ݐ�B�T����:��8߫�Ƶ�\r,�=�³��B�u\n������v}Э:�f�؝̮���t��ħWM?���)�9NWBkn�eT\I���Es�FW�.�_���kZ@�3/}�A��=e�g��k��#�y�	��5LvJ���$�|��'���&����"4�M쏰ܥ���q83+3�b�4�̶��2��AQ�=ո��ĆW�E���R���������\Awm��ʊ�|>ʇ�����]1�"�Ibxņ9�JN�:��Y��}z��{c��y�r�a�
�9�Z=1=��]�i���L-_N����:,<��Y��f�y���.u����>
Z�+�^�2Ⱥ*��Uݡ���˅��֮�6�p���v[���v�VF�$�*4�r�8:�87�Ⱥ��T(�Rk�_�y*�I�"�sE��$wmۺ�n��l]D.�xC&���N�n{��)��cWR�^pb���an����V�f9{��x����O����]CoS&���o\Bv����c4y���]��`r�Pf��b��c����N;/���
m1;��'�*���%f�a���%�n�.�ZVNZ⭧b�O.�[+P�Go��v%�v{-�ui�n�[��������n|KI�7VN%o�"f��܏��hy7��fj��M�+_���_)��*���[snᕗ����uY�:�*`�e4"��B�\�8�:a��`�{�q�_`�\Vn�Ec�/��7���3-mM��]���/���i��#��X�D�Ks�c����U��E,�j����;�V�mRbǵ���w���6j���Jޱy2tV�^.ٙ����:N�w���l�'�b�����Yv�[�ih�|��2�+��$͑�v�f��h��GϹj���hb/�<��X�ζ�]�mh������v���fI�d� {ZE��[;b*��u������N�������os�V�c�\��p8�\�k�|��m�d�ޭ��݂xv�tT[��No7k7`.�r�y�M�3x�u�]�6��]�{�0�jCu��%�%b�+ةȉ�s�eG	���N5�g-�"��nA�xsCr0�������4�S�N��+����*�kZ��Y|]��<c����:x_A˹Zꔖ� lu��72�T��@۝R��l�"�3xǯ.�]J�.�Ħ�-�ܐ3��w�lr���[,S����zVd^Y���n��L�&S
y�bwGL,��k�k�����j�@�H�l��y{ٶSĞ��{n.�(_rEg̏�v�1wF
w��V�RWp�V��ӱ�ya�3�k��T9��X+�t�^.�V�oMˬU��6��BVV��d����H��:Y���f��̫}Le�~��K-���Jc��-"�m]�Ve�4m�|�.���²V%�ׯ%M��6ê᪡)�V�uK�Ǩh�)X٠�x{:�lc��A�Z�X�
h�tv�QŹ�@��M(s�,�Uj��t9�����x�s\T�B���#�^��O+5���P�)���<:tn0t�4���-M+{9�roE[�Qb��T������*H����E�b����<�U��
�T��U�����K����+"V��U�q ��>4I w\��Y6wW+����.].](��i�N����':e͹R]ۢ�������6䓛�&+��.w:*CWM�;��0:���:\�\�"fS�ΗN2�qu�]�%��\�wuwv㮛�滺�!���E:\�w"�sq�	�n�����eȚ��!��wwK��.:��wL7w�������;��]��3��s��$�k���
r�΄�Ӧ��ur��D;�]$n�8S��ne�p���B�뺸$�]�%ӆ �"�u���"\�:�f	����H�h�':9�1r���P�0sv���wti�1�uwk�l�l��2��wr� aI1sq3u����L ���.���b��g:	���v�Br�Ns���r�w$M�FI2����Wtn&hw(�wG��e�d�!_q���]yc��08i)�4�5��7"��Ui��E`�����h��F�����Ό���̥.��Wia���M.�S�>�Y4�^�oO��/I�=Q���k/ zpJ/�H����1���ϧ��,ΜSP��f|�J��b�y9ϖ*�W)_�]�/�ü��N���ә���O=��v��
L���*���"O>�ρC���Ȗՠ���֡N�T�V���g�FK�Km�O�»Wr��7D�@�ΤT����3��n8�%��'nwvU��tU�~�R�u�-�<��UN�㌒��ď�.�Q^;S�K�j����J������Q�/͚�p�[�m��^C4�hN ��|�����L��g�c�q9QW�*���lwQ3ڴS�zv���i��v�<�%wF��S̙7��>F�mǝ"��X)���C��m�]շ��ށ��8�Ӂ�T�:'�P�+F��������N%�U�����[sT�����NG����&v����r	�LwF΅�zt])�v����r����sW�MǐQq<��p+^#VӸ���n��>�N���}P'tº�~7Jt�� ��~�a�NSߝ9P^G���un~Ƌ�ȋԩ����p���^��������@��g
�����I���yv(���Y	�}�vfaT!Z�;M�mB��:�Q��]J���)m`��cZ�� �u!��Cr���p���plH	��b=zszN���o�W^x�����|�81�UM׉���gb�B��ӱE2{��m�&h,�$N=k':;��T w�l��<��Lyt�{^���3�_	��e"wOX���ɮ/���Y�}��
���9q���uDiT}�U��+�H�);�{9��֫h�ϯ��ƳML����Վ��gzB�~bg�_�2���9��L�����VQts�n[=����8�|�П�)N�������˺~�Xk	3>`ŋ���U/��,�
��^xƏ8r�(~�ϗw���ٗ�H��ޅ�p������e$�|g�L@=Ċ.R7S<9�BŚ(\*N�\��&S2�ǃz����ͺ:}x���Cv�eK7���z��
���f���{!�p����gqs7�6�Ko
���N�<M�]H�wv�ZuR� S�G����H���瑞�p�e?i�	��b�w��q��gc�>��~�V3Jfd��RWN�ʯR�_���`k���U��:7 �gx�.]N�Cr��s�3����h�c$>?{���"�����}&�G�h�9��wE/�)��Y4:������W���!6|���n4�r�;mv��-��jRӯ]:(<�J[�~ֹ�^�A�li�U�6��9=�_2�����E�u�bH1ާN��:f���vٴ:�s�As|��5�h����.CsH����п��i������:���1p�vd�Br�y�`�~�['ԁ���_�z:��iв.��7s��>��oFE)zj�e��gs����tq�9�����p��c�.� �;�ñ�P<�s�wL)s�z(�/��4f��TNZ��5��L�+&��A��>9�f�Յ>�Nhz�绔3Q'h��څVS�[�j8�7;u�泼��l�4_�{�}�~��T�NG*c���b}�k�hN�(�S����eᖂ���n3e�g����~��Ui��<}�@����"L��)h�CyQ�ȅ��o\���'{��v�TGw��>Ϳ���:y�82�:�'F�NC�Ѐ�iW������m��w�����m܉���6��'ʨ��.ۦr��fXʀg���|n"��z�h>�Ү ���Q4����Syn���k��T�8����oMeS=g�=Pf�=HI=�b�X�.�
��p��[`]=ڿJ9�(�������!�u�ip�k��\�>G�*��z��
⌯���4��/){�!f^�J��u��'U�s'�4_�q}bje�{2��>�W�	�J�<��"�&q�2p�B�n\ �� �c��:���x"�DV �x�7�õQu�$���C��\:f�v�;�þ7]�3��|l�c��b���5���U�� �����Y�^�i�d5:����oz�kuL=�IH���|q��y�����W��J�te�㝋n*�+�9
g�nN����m��F�:�,�.s��S��܅��-$�í��@��`+Ƴ�^%;H�7�H�3�&�m�O�o��d�USdw���uƃ�UU>7�#�ā��M��>grc���\�q��A��Y�Is�dA��V�Tm�K�O?��������SN��2B�2"���:7Wl���{�BE����������*�:�~�K�fXhT`�e��yn�K�6�
��=��ӂ�{;�}~[�/��z��˴����{|STm9�*@iQ�F8�ΰ���ax�6l���=�^f��'aqG�����ˇ��w�S��bwC��d�ߝ x�O�O"7��b���)���t�W���zN�������gT�񌄜W3�e��}������ߦm�6�;�N��z��9n��<�98��c�l�RrN���Y;{(	���:g���;�=]���:~�Uc/{��:�H���͝U`��-7nءmT�8A6<��ɳ���w�u>��s�f��M���11"����M�U՘�6uu��-CZ0�Zs�k�z�B�	�3��o:�l=��	C5�镕�#7�uŤ�ԼLn2E�=�`3��6_+W�l8و���'P�x��*�q�v��!��>�|fP���d֛�R��i1���:��R�|��u	��P
��>t������kYUǢ����L,�u\ek�׹�6����jMS�c����u��l[�dS�r��	�U+�$�!q�=P��2����o�.g5����v󋣐72�\Ub�qo��ϩ�c�V��=;%Z����|h���U��X����y�]K�GM#Z�<=���W�C��}p����e�V���'Eۈo�{��ʽշV�M�
�3�$9�h����'*�࢕x`Q�]�;�>��ڢ�ǁ�S2"i�����Q��o�wzc�����U@��
D�Ϧ��(z���0[T���gՍs��\���-t���S�Kz�'���v�*�Mo����H�+KPat%�V��8T`1Ti�B]�g���"�$�����gB&�m׀sn��UN�㌒��<d�S���ݩ�rN��G���V5��
�Q��5
��tm�\�i�<МS�`�Ъ���_K��?Q�5���V^��=f����_�c�YU���0�ʖ���NUq�vL��{$��wuF���z��]T��Ǳ_֨�=��L���ͺ&��ҽ\b����n�mL����a����!;���,��1���CzvL���gWa*eww�����NM{c2��yo���?A�~סϢ����������I]ѼS̙7��	��t4�RɄN�r�����kޟT��yj�F.>�tk���S���s��޼�Y���Ƨ��*���z�R���g^�h�E��a�|����ᵡ]KӢQ�scg��˼d{��EO;{~���\�"���\�zy�^[Q:_���a�}$��a��wL+��~7Jt�@Z���e&wX�Z�|�j�߁Ϛ��r<�>��6�n7^'��0��ިW�ZFù�-+wd��:&��y�W 3Ϩ���\��TǗN�7���z�\kU�{>YZJȉ��q��8=ٙ��3\t�Q��>.�����\�Ҩ
�*�g�$}�Rw�=�:5��=y���RQG���Mm������%�	��WL\R��oL���߳��]�gʚ�}����� �.��qU��(��;��O�k�_I��=S����fB�|����:CbW��h�l��s;���EK>6���{>SZ�8�̣��J�>q"˔��L��h�����ff�I��k�EPs@/��x�=/;^L}ߕ�or/<]&㺪G�M�������E-�f7/��i��'�Ҟv���4�"G�F��L�n�H#<���Np-��.��c�����=\&�jRS]v_n^=�x�YK�b˝U�gD�$�N��w鿿�C>�u����8�̳�DTf=b
TO33��įiλ���y�&���-]qWϳ�W/��'^&��p��
��͢ jj	7�����S~
�ϼ�1��.� L/�����#��sų��ՠ�n���kaUT��v�Z�˫�3�� g�/�@�ޖ+"������gx�+�]n��ܾ%��3����p��Z��0&�3Z�ԧIVS�~�!tzh|�	g�i}����ԅ%�tb�N̙����Y���r->���
��u	ȢW.ODu�>����X6��5{(m}�w�7�\��6G�R�7Ѿ@��΃M���9`_<��~q�����0�p't¸�u�n����{}|��Vt�SB���yhb��5:�9��g��s̺���;P����"�g��e��n�v\)�Q���85�~�3��x��Ls9uLO����'��w!��L�r��q����b�Go��~�[�\Q�O�*�>�yǵsʚ9�To�_���R�^����ƕ����s�yRm��p�W	�~cX����p�߽�������'{1רbQ�b�]�k�]�1(A�Ӆ[����v�FW�՚q�έQqa�X⎰tC4c�6��+rr���ǃ�4�q�46�+U�����Ă����y�����Gǵi��j����t�b�PKGF���?rߴ�:�J��\��$}����K�N�o�w@��o��{�/Rۮ9p��P��T��qJB={4hU W�u�����0|j��讋��)�'IȊu��B��1p�ۦr��a��	'��"�X��鶼*K>���ڷ�yoE��'x3TKgq��~n�zzmpY�R���U�@���b��g&c�#��h�;N��6=��2�zz�<�}:����qz�m�wl<�%\B�)�Vr{�cv�Ƿ����zi�+�i�w�2���yP�R���{OCrt���n�ѫ��{��y�uo��]=�mȝ/��=S z`7P*�s /}���E:H�s���Ù��c향W��V���@��[��S�ޒx�9���R#�ς��n�ԥcW���M�D�C�/Sَ�pv"2�YE���^3Q�*�t��i�frD{��/���3*��br�x<�}�Y�*����T�K������sR�j��|�ƁP�e��t��%�v:k��	_�y��˕���'z�)X݊�(�ghsv:���v�٥��֠��B�u=�H�f��\<�k���SyaS!*H��u��,zΣ���uo�5���M�]us��I����]����O�����=���JS�3mb�3�0��^���������<�<���q��
n���
hmǜe��������U5�N��Fn�F|o�Ul�����!(ה���O΀ro�wHO����C&l��1wo�^�2n�kM�����1`�N��9ZN����W�I��N+��uLO1�W�>9���O%�o�^�����M�Zo��N,�~�b��ճ�S��NO�x����GUr�nd@6��70M]�>�"��iH���{8׻u�7>'��3(N�B�kMҐ\m �����d�y�*k����!�S��.�s����'��q�m�Ow���F}P��u\\�'�ܚu�UD�^T���uP��@��\��źa�S�vB��	��GĔX�������l�7��o�ԐW���γt\f�fxu��V3���ڎ^�MS�+o������Ǵur�[����鷠�Ng@���L󘸩u��,�F��ԭ��9��Qވ{��+ÏVv�:VZ�6��pJ7�@�Pg�G�iLI<��b�q��ќ���¶/����j�����������8St+��u����gL�x�р�oA��o��G
�����L���n\�&˕h�i�3��.-.��i}��Tѝg����q��<�Jl,$boTr���VnԤ��^��pa���sE���Bf�uq�g?m��ۅwl�,�A��
D
>�}5�
��~��~:�k����`������
�xk�N��n���v�*�Mn8��H�H�+KK&���wǶ����ۊ��d�.j�Ϝ��^3:-��<�E\*�u7d���$x�Bs�s��;�����=����L����S�ͺ�[���*!<���u0�K�MF��Yss��e��^�M��ޭqS���+N��B�BJ�#̙-�W	��,�ݘ�� �K�]h�1$?:���(��NqS�tJ�b�+MF����u^1�ĩ3=��2��Et��X�P2ڀi�t6ӡ�Ǒ���X�Ф�86��;{<n]�A�`s�zoo��.$�׭C�7C��f��?\W���u�>}$������a\VS�N��_���r�Ҥ ����_��/�Ty��>~��6�kr�nP�����^�V���9�i~N+�G5狢�Ol��r�"��22U1�ӱ�xs[\:5��=�B��P�DG��42]�,蘳=�s-Ε�n��>�)@�I3��h*�s������WS��_[Ͱ��=�-�����+
e��Oח9\9X�w�e�U�oI�l��;"�4}5v�C^��^�vo�<�o����;����JĈ�N�3N�	ipަ,���M��un��Qv�UӼ�y����K�θ�+Eln�1泌S%܊b��f�f�.R�W7���ᦽ�/�x��'���v��+��<u��<˫Қ��E�,�P�\���ns��������_uv���>��^O�iR���:�[�@���;ºr��βk
��{����#iv�0һ:���S!�=��_o,�����r���M���N��CAq�=��%+9����ˡZx�X�_�,�ͥP������r�n豖�;PΤ0vlq^�)�*uuۏip�ܹ�J�oI�`�Z�r=�O��v^��T[�wjn�^��i[k���L�
��+3]�A��kB3p�`�fn��J8s%�c����8���!u0!a{wb���|Z���@k�a�ͬ�w��n��:�B#
�ں$ �sr^0�J>5!ֽ��<�b�rҴ9C��j52�n_a��H6��v��cf�N�5�O��5�٩�ۺ{I۵yEnj��<g�+5�OwC���ha+khh���.���^=�����.�������ˆ5u2�ͩA�Ӓ�MY�X�Ի�*����aꖺ�Zǩ-}���#��um���s]46��[���m���(V�?	{+��O \�n���=�P��8��P���~�C/5�u�PS��b���]#�xOf�f�]�O�ES�7~?N�,�]1fVg;�^桋�!���p�����E���氱w�
Y�跠�O���ʶ��y�X8Ktv�Z�����MO�ۻ�����aR��=�Jq��|.�����"E�J�<é�hl崫(�R�?7C3.r�n�������.�Ϊ���I��F��Y��,�I���e���^��if�(�E��uڬ�j띵�n�ӄ2�JT�R���$B�ՉY����)�n�"M�S�˨����}w{���ޛ�C���L+V���(VM�N �o��|Qϖ[m�P=4{F�t�55u���9s�����U�N�e�]ER�X��b��k����ś�iAt#׏"o��`��>������*�`�� ��mv���Ƴ���j��W%�1�E�ٹǔ�O_a��4�
ݹ�A+�k$�<uv�Z��d-���	s8.��p�9�r9!]mX�
8�8�o�wGo�v�Z�>�<�_g�t�iZn�s���oT�\T�d��tz�mi�(k^u���Z���+��A��ruҘ���Ӿ����缁W]t��M��S��Xig�#t{�v��
��ǇC|�e�5&�`�{�ˮŞy>��F���YV�@!4~�aGq���B�%8&�%��w0��!�6�s!%\܊s�9�ˤQF)��]ۉΈ2�I9�wn��LR.wnK9ۜĹ��2Hd$$\� �3�D�r���Fwp�CIs�;�b��	s��T�#@��")���P�̦�ۻ� �;wXF��!��]�9t�����`1�1s�wq��a&�.��k��L)%��$��wn�wq��5��ن���N�r��М���.p#7t�@���lRs���b�]$�����Ɛ�h�W42BfR�bB)+�2 ��p���*I��tF�.�bcI	��K��\4DI��3F#��t�F�%��#�׏=^y���ԬY��8J���s$ut�0���N�A��{:,��f��JeYFE���@],�p��v�ؼ*���-�_{�u~���3�qJ���>7���Ҩ
�ܫ��WP���Q��~��f��%�^�:����yW^uGC�I%�L��&|�L����H�7�Y�ҪDg+(�8ܶx��x��E��D]Ew�aN�XʭFק�i���TA�?��T�p�/��2(^xƏ{�R�n�ǞM\��pwиu�ȷ��������~�5�Ï\�>�x�����H��#u3Ý�4p��6Dܼ�^�(�˗��t���k�����>�u��n�C�ʖn9T�@�)P0�7l:�Ts�B��p6{��})vp
��ވN�<M�u#n!��q	�K��R6��bMW�mK�4Ɨ�T
���]g�ax�x�/G'is9��؇>��w�-�c5j8zy�����d�<��Ol�s'C��O�6H��]J�ѹ�����W˭Ѹn_�',G�zހe9�J�½J��7ćY]G�!w�z�T��4.)�i�)�����ۺ))�;��R_�tX�f������d�nz�@ur(���S�q�0��O��]��Qxk�P�J׻���i�e��2��/Ev�wȮݬZ��n�̡�B����X�JB�PSYi�~��+��Wn�a��4��
��Lʰ�˲������»p&ྮ�\�F�����rq��;%�{��3n���A8�4�L]�J�"4Oy7'h��C����мn���nX��<����n�~D`����C�^6+��7;һ����bs� (4��o�w�4Q�S�_�S���:��ҙ���{�C1�v�����gH�ʞӯY�՞�o\s�������؍-��r�hduU/�ʘ�|�X����Н�Q��	��wn�e����j�����Pvt;�ʭ6'�aP3��~�S\��y����VL�z�ssϧO�3zk�u��;�,c~�����&|:�]JC�Ѐ�
�w��w����:�[u��!oB�U�q���}�ޣ�m�Ow����>(]L�7�#�4&���MC�1;[�'w�A�* ka���6{)�ئ��_Кۦhq'��|h�R3�G��->n��1����Uoó�<�v~w�5Ķw������V���R��<IUf=�jL�ܾ���Tt������9��Q5]m��r�d?Q���H�n퇞3��#����[[���NuR nK�>`o�<�ў+�#���\D�}�
�g�v����܍��]��6biL�=�/ټz iT�,`Ń�<Ó��/h�U�����p�m��,�\�9�3��1?oB�Dc�c���X]k}����</Gd��G�4f��hm+��m�C������tA\��N�mm�	\�	{c �s;GQ�R�i�uBx��qU�L��	T
�'<+>x�gz�}��c>s���{o"���*~�5��p�q*�)*�֮�
fe��\	�>�J|��,ugz�&���7��n���OV�V9@QVZ�|쳐�u����;��SN��rD{�LV�W�s�}؟=7��w�{��g��[�O�܎	u�IS%�2���F�@��.}�-Ѹ�$�7�����)q���;W���b�:&{^鐴�8څ����	*�7��
m�`x��)��qu�ٙ���X_HS�9�{
:_�����r�p��{J����7/.}�w|u9�X'R6.־�������)�����R��9,ti��YLm�R��7y�ܿ\,�������gw�	��HG�3�3�{�ڶ����'7��9����3�s���V�	O��91xs��xo��,Bv���s�q�B"������q9�}�U��1F�����~��e~T[�Y��� >�kY�q_mTކ��n� �3��"��,����=�������\k[u�"��+9}P��z5Hށj��rZ����v�%���bī��<v�ö���/m>{@�x) �q=�a��t�Unit��͊�T��,
qj	�ľ��\���jS�aO��S��Ś���if�8�d�݇8nA]���"�;���Fg��o�Ċ�k�e������Fl�����:�J�+9W75NX~Q��*���ʡ�sĞ=V��K��ΰ[Y�GM?x�9Q�2��E��ٞp5Ռ�8���閥�t*��A􈗺�f�N7�5�t�M���Iu>C�u2��Ժ�qd�5q�[Ӟr^9�Q�6��L��k�zFP������8X�S[���bY�*3�& t�4Jb�g�����Uĥ|4Q\�l�W�H�Ŷ���o�-�:}k]���;�F�,�B�*2�H�_O>��P��'��A6������zf�%`��l~�5��%b��*�TS�T�F�� .���u!���Q�TfcQ�1�5�L%Q��!�MR	ˮ%�3:7�n��ǑW
��OJ�VU����̷{��e�#�9E�G�ڽ�h���p�[�۞��� ��F�
O-�}\b��>��2;�K7�}[SNUL52W�x��^�T�v���i��ۅ�+�7�y�&�t��J���W$0����*:6^p�"��
T�c�zp;�*{N�[,W�ei�ޗ+�]ߤ�[�K��4�99�쓷�����u���O+~�Wo'P�X6P�E�͢R�ѷ�A�W�̐�;��S�Cn>���<�&�=s�U�Q�[�|�PWm�д�9��oV醏�8�X�N]��[�N���h����t匴��N=��I#�r��6�vF���*���} �n�o��1�y�'�l����
�^�q�����,�$�W��iR"�8����f��#^N�t��Ue>�N��>�9��e?T*]VY潀�5��6�O�o�æ]h>�T��}�4�F�V�ͺ�׉����4<5��5}c]۹�sX}��'S�ڬ7E2}q��	�9u����FJ�<�w���;���9'�7ȉs����×
����ޫGT�;'G8��4gjӪ\�aP=Zz��s�eI���Rw�'�J���ه���J������[E��ze���ς�_Lm)�Fg�:`lg��.���e����m�@����**�G��;��x�r��r/���Ǯ|P���U/��ɠ��x��R���ɽ�Ûà���LnC�}6��ֈV6�x��'��<���H�u".7�{�z�\���Q&i����4P��n�s-O�Y��:�t��۸x=�#���ߌ������fxٝ�<�w=�Ѽ��0�Ҽn(��^�wq)vp�S���a:��=u#m��i�K���]1E3UGG3Y o�7����|�
�{nތ[ı�h��u�\�!�Gq���/g5�hk�ba]F=Rl��:��mmb�Ƽ ��Ē�!n�|���>���ݕ�5wNw�Kd��ǃ��7(w�9\b�1|ڊ��g�mp���������}>�i%�0�$x��@�������B�N�8�s�#�9�h-���썖��\�Nh��ys��t����R{���τ��S�X܀S5�w�B���7/�g7�����&ߏ��h�W��H�lր��1��)Ѹ�_��b�R�ň��N�~.�7�C�[�S�5��Q�7�z5�"��F?;!2�k�1���d
�����0��O��^�����q��Ign��sz�o;�W[�F�x<2;���N���nX�Q8v#�6�T}�,���'D,��Up^]�g�q�0�=�{>�p�[����S㚝g�S��u"�I'՚�u\L�����O,��Q��g�=�
Ⲙ!�6r0�5�~�3/O"Ǒzꘟdk�h'ُϜ�%�g�{h�fN]:��uN���GgB����p9�&,�_�\,��@)΢!f��іjnf�n�<�d��r�f�Z�kE��Ν&��-h�#����V ��V��-˜���R�������O��#���}�'z"��]xв}�A� ��e��)񕴌�Y��ϟקQ�qhM;����4H��ظ���x][|������ �)E���Т�换�i�U�\�yr�b��L�����dǎp�'v��Iv�WNZF����i�����7�6�Ĉ�n�'˺E38��;����H��-U���o;͛\�m����T�_�����[��6{"�p}�kx��kn��}_��F}\/��x��V|>ތ�E��.(�J��� y���g�C��h>*rx(ۙE#ę���ˊ����v=�f�%�8��Tm�g��X�}&���s�����D?��Q���e�J�M���W�[wJI�����O������3������JWÑ�{OCrt����cc�*6���W�%
=~r-���q�tJ6��*�@�@>g�o�{Mg�x,�S��+�z�ofʛ���h�����>�nw�UL�ߕUJ7@]B@���B�%���(�z�Yv���)Z��l��l���a�_Qe9�D���F�N�Eoʦ��X�����J-��Y�3�Z�s{����4�S�V�\������K�e���h	���yn��%�`������ot7N�W�f�r����C!%WF�1K
n���
hm��p"��z;9�Y�ʨ�;��gj��j���܀�+��������~�Ly����;�9��M��P>ga����B�ޤ�q����v"%A ��D����M��6�2S42hX�j��o����2�Fl^�����Ru��N�(y��mw7��V;����q �3�<�g2��R�������c�7�I�ޜz�o��)���6;L����:o$�h����G�����ߘ��y x�ɏP����*cn*V������n]B�zc��z�^�30��yD�C���y�Ấ'�?~���L��$��?�h��E�:6������[;솽���Fv<�e�8A��p/��#�74Ϲ�{v�ۡmΓ����'|xNӋ�V�72+�z�i��z'�>�y�:W;��*�>nlf�'��eW���} ³���9�>ػZh"�����(��q��U����6��Ф�r�nkm���w�=q�=�	��}@G��;M#�Ύ��q�&���4fa�W���z6e��.��:G���閥�t�W�r��]����,���a��$���$�Dπ���L񊉗^㝓\j���>d2�OV�KnY��^o��,��o��SZ����(� r�>`t�4Jb���f���V��y�=����%�R�kK����z�q�}'O��N�^�=�f�9TA����y���y;��o��8��r�t�"�%| s���c�<���]��ۻ�����7�@]P$���9���u�8������o�`V�VO!��/]�7�KhWk��
��]�S��TB���`~b��;G�,����H0P`�-�D�<�ի1e:n�}aI�٭��Z͈5�q\���&3�(e�U���zQ��Gx�*�q�P�ks���L�(ܽ��Y���	�)��^��d�95H(s>e�p"}�n��w���O$��~��;Q�>Q'�\8�ާF豕�	��3ܺ���u��f��<F�	�V�|n��zn	�|���/Aq
�Lx��0�ߥ�!RS9G���W�z��2d�^�7�+�/����s�S�Dd%X��c�zp�63��LU���_o^\#oվ����^�W����ЎJ'���@>���ߝ1^r	ꁳ�kB����E�Q�w۾v}$`�ʲ�<�ή��8�w�]K�25:�=�F��D��{�Xq��� ��7�ֶ+�)'�63�3��}��R'���;�]v�T���*|�>��"5��'yT3~n�O�0O'~d�ȹz�
�>��Q�Q�\�u7U�G�>��\ �����*������;!�_�kH]����z�i�mwP0�%U��`���p�uVu��|�&;Ys@����'c��y�ʗn9{8jS�xu�ǉC�ς��}1t�#Q�Y���&�=gӶ^�9� �+.�z�Q��ޛ�%�{�\����z�q���x�i-p&��z3U���E��[�A)9|��[�wǫ:���R�Z/kan`�h͜v��Ϭ"zW%�����{\n�vn��<��
�Ӕ��dn94Q���2�_�讋��p���e:�뎚��=��ϯ���f=0��T�p���|�g�����~˯c��]���0j�,b~�ϮW�
kD+u<xx���π���Rٿsf��
:�Ӭ/����Ś(\��G2���E_���m۸x=�"��(o~��s�韅Z[ۯ�.Oմ� ��]Zj#؝���t)�|}��o�z�F�;�B�K|<�]�~^疫��Q�3���4�č2[���u��;���≽=��9�h;^�U�0��37&�z�?F߿E��U�ҙ�(oT��6H�|&�����7�f�]l	u7S��{XG��+���2׼J.!����+���S���$.�U��>f��a���U����*�mST��Ýr�t��G�Ӳ/����ς�بN��)��'�>��P�z�d�Y�+o��S7�hC��G:��}F�zc'��x��wB�:
fۖ����y�T
��d�Q��;��	x�Pk�zf��jQ&�㳖_�wK��ܼ���:|u9��V�s�懯�\�����c����xv���O�ɩ;����tg72��{۵�H�7��`��l�wt�*�!c�z2�i8�d����˪�2���)�IC���ٱ��6�s
ur�N��H�W2�Gj�Et.��⻱�(3�i2_K��r�E���#�?s�e�g�K��3o8���w%�j��*ie@keT�U�*o2E�u�t:��Q�{D��H�b������`o@�j�Q��W;u���	�<��"�R��j��?ڌ5��t	��l_<�m��9����
]Ϣ� ,�k1���������:��Fe#u�%�N�����yV"����!���S��9�9����t����;G2&�A`Ia	�g���o7O��8_�)qr� P��W:5�Q�㷊N�8���׺ɭ�A�=�8��ꅎa1Æ��+,��V���MM���;pP�g`�2v#��v�z�|)���w\ؙ5#KOn��5�2��u'�Yݡ�e��FT���eι8X��!˖v+��0��dK���#���Z�[u8��\�Sk�w4�!������T��(*�Z~�c��i麚�ާ���tW{O���呢J�H��tE#S�=��\ګ5�Ct2gh��q��\�j��X�|1(ç\�����^�6󘠈����S|)b}�)�`��6�^�Y�� ���/���[֐+}l<սqV��k#DWL�w�宧�q_�v��Xs@�ӭ0k���\7ya8�hh�ו-6".�[�-���ՠ4��,��%�)��!�N�h����-S���R��I}�\=���x��l\��|�϶r!>�Y�S�v�J*�9���|�4��KB�H�oe0hVf����?__u�J+����,e�_C��ۚݳE�2I;��Hi�Ճ�$�oX���'��n��E$��Z]���Xڽhb�����1���.%~F��O�ּ��
�4 ]XA��A�Y뾨�`Mv�|P�i�]�Uϋ�T��L�/�D�[A%Ci�p�]w�:�{���.�
�m.L��ö��ӑBy�t7̦ J�1X�Ȼ�������ˉ�J�
4�Ӽ�_9�=�˄Khws�{��靈��c�n�GÏ,�#R�˰�U���۽U�=�Z���/9T�M�Ǌ%�{�p\Ò��������[��,X��9gDm*j��}���sv�YT���n�A[�@�,���knlcp��b���|~ nD�tHe_T��t�8���u�+vH�i�/2ĝ���b<Ťw3���\�3yw(��0�`��L(��:�KW��Q�EJV��|L�ָ�]�X�8�;[Z�-ui�O����X�XLuk�oqZ�j�%I�@��Nv���/Ep���P>׬E9)�5x2�'ۋ��D�m��}�����y1�0�KK;,��Ꮔh�&b�J�}ۮŠ���Y���G�t�V�pp[9JO\rY ���"��)"izWw\	�p���fDbɊ�@f������$�0�"H��r�EA�·.2L��$1n]�]H%�	"�k��qI**H�����JM1��.�%����wv�K�B0�&JHI1�!1�.�nk��79#%� Iww5��C�Ps��$�Q��"JD��&�d�r�˘\�$.n��S e�
L����`D��DS; ����p�K;�.t��djûr�Ȅ�Dd���H�Ww�w�!h�&�20��
ɱ"��ɹWGw0R(cw�Csv���9�h�tAP(���������=��ʔUYk;e��u��u�e����Bb�Va���ΡGIf��s��T������M�mvV����g,��޾���$���0�:���h�ɳc�����zRR�3�ꘞ��A��;P���q�.��^�V��J�i���2vt+���<�T	�����3ȁ)m�����'͞+�T��y�#��Y�s�֋���t�QP���5������a@v��OvC3^���}�쓕�\J�[��:���|�芌}�^9g	����5>_��!�xk1�ˬ7G�YY=�j��b�i��q��Y����g�������"~��H(���b#}hx-����6���?A򌛗bI�d!�׮����%����C��h>8�k���GPg=#�0�i�Z��slk�m�%�~:�џ3qS,s8�`�gu�r#�����D/��Q�bǘ�xmL\�O��p9Mٜ%_H���,t�����tgǙ�ǷJW��N3�=��ƌ�����2q��<�.YF�ͻ�������D��+� zBU����_g�x,��"D���UO�����ބEa}��;���'ͻ��hj��F������qJ|��D�n3�^��f���ίd���=8!�7������{S�)��h�R)w�n����kk���V�`1J�h�Q��4r���;z6)��1�к���,˥��_˨u���;a;]j#�q��\�ɾ�=9�[*ה�I���=��a�[��bH=J��{}�]���\�.v����r!��%�����;���M:7�$.��?se�ʺ:&��o}���=�#3&����"7���\$���,}�h�\
�����zW�7SИ����d����먨���q'�ʸʅ�����A%5G�K
n���
hn�ҡ�-���3���飕�>���x�6;iV鐴��:�����U�ڿPK~z1�A�p-{jwc�o��`'t6ӡ�7~T�G%����_��F�J�t��y�ʺ�k��O'<]t�ߕ��\I���c���ꘞ��?]
���f���I�ۙ�:4�[9��5��L�"�|?�5;�]�=���܆1U/d�y�sL������{�Zq��>�0�D�9�&�L��ː���wУf�i�:��s��"��<����Oku��r�p�ֶ�E�'�:}��}�+�;x��]g�F�{��z�ʙG~� .��`��*���*���L>ȧ|4{9��G+�>�8ՕW�/_M�]z]\���I|A��ȣ/����̱�UY�8��C~�1�{�0���ѓkb���i��.֢.Sqge�Ej��Y�,�CC��a��C��'	Ƒ��R�-��� ��Z���y�ā�F"���ֲ�g���f裮bq��K&���o�u5|*h����Ý�)����-N*��ɂ�]�7A��|Y��t��Q9ki_����ӭj�и^��/.xz�|>�Y3�1U:�U�F���<�C�Y�����p��a�����M\?b��^|=8%]$F|���h�ē��O��s�����>Rj��-�2�k������޸����ه�mK6��ʠπ�R [���뮯xW���B��\��Fr�	)u��+���^�7]���;�qW	�K7�"P�X�g��n��r��4���ר
'̵��쐅�ɫC�y��3>M�ۯp�EmP�wN�q;����{dۙ�|h�x�<r:�7Ex��	��Fw�B����n��ֆ��^�a��W�$u�L���gУe����7�Y�1q2WM�M���b����7�i�30��]���d3�g��/��ݖ}k�&J^�5B���Bȯ��zr�cӀ��po�I֊Ұ��AG�����9]UOu
��Ī�Ìn)I���>����y��y�'���6�+�zt-�w�31���Ed����j�ѽ(c�˼3�O�3S��nͣ^��+����a|I9�0�u*!l�UK�n@j��i�j�1���X7�ʘ};����,N�]�����_I�ɨ�<��CT�)�ݭ�Jc��i=�M0�hI��4���wGs����X�1��`�Z@i�=�+I���/Zut�ښ����܍����C�y��\`�w2����eߌ'��n��;�������uR����3!��}�բ�ͺ^o`����]=�]>��D�30��Aݨw�Zo��=q��ϩ�3>d)TǗN�����ǐ���4i�����a�[[E��׉��7g"����V�����ޕ�)=ι��ݍ��Z�Y�7{=�;}"�����Q��b�V�ᗒx�̡�O�Ϣ�_L\R��n4�=7j�hv��V���z��A�.�[�ʣ�Br��}p�!Mo��i�r"�H<��B⧫��P����G�b�}�r�DU�VK��Av;ck�LnC�}m��	y�Dn�P�L�mU~���͈��k2��1�T_I��{���c��x(z%'z29Ĵ}��Q����-Өq�2���]�!`�5�-,Ϊ� m83�'}@y������[wr�g�9O���3Ǿz�F���lu��ݗ��}��#}RФ�g����<BS`zW���Z'\�������OE�]�|�*�b#&Z��G��uhͪ����I]7� z9�
ʕ�����giu���A�ܱL�]m�U�M�y��X��ϸ��n��;åe`M�Ҏ* X�wH.sh_^�=�Wj:|-\���ҏ,����13�Y�6�xR(���o_$G��ݡ��l���]�uo�g+��8\Һ[闗eZ���D2��}��/,�5A�.�f�3��UvMd{�tU��ng̖Y8�LN ��f���tn:d����X��O��R��L/O��6rUum��������GZ]wF-$��p5��TlW�в|�S�q�0���S�J�wtd��j��g���zR�i�(fr�$��NB�l�50�+M��P+�yfOgF��=�'����e�=
u��>�	�:�7�Q�+��CEF�塟G����N�3�h)��'4=s�ٔ¤/:]]�)�˂�sN�>��gv��VS�tV���O3[��C>�~)9̄Y�T�5��U�'7��p�V�܈j�:t>:vt)ɟ��2t�iP'-��+�
*[뽾q�=�DU��Ku�)��o���޹ݩ���G����x-��(�RK�����3E^-I�T�{�z]r0:%;l���.7��q��5���p����_>(7��Ď�������]<Fl�>{4^�pg.x�o���N�>ȅ5�a5�\z�z3���z��,�4�{ۚ�tҏx�9^K��W�A����q-���A�E;A�ϕmpN���di��گ@�	�apz���D�th!_�eҟ]�;��j+,&����ٲUoȬ�=�jl����M�wo�uD��sٴ�иc��-�٥d�Wwf��Ě���N�SjXW�N���=hB�<Y}tK�{en��oS��Q c�}8껢��㤗Pf=`��wFR72�#���&���>d5:�~����k{�r�d
�:=W��G��*��Y�8K� SR|��A�F��L�YQ^�J�H�F�P���y�R���L�>�H�;تF*��Ў	E8���@�@>�<+^>ݾϽvk8��y����KvنoԴ�7=�n���û�h)��w�������c�wg���_�����g<��s�^�㓴Ϝ���C��M��=�c���TӣĐ�/7}�M�f	'֭u��Q&X�ϫh�Q�W�¯��� �:�ͺ�[��
�Bx�
�nLB~���z��L��?{G���=���*W�h�����N��!�Uto�]L�n�-,��W����z�e�Aׂ�'p*9V*����ϧ����!it}V��z��dw;�4�/����~��������>�n�mǝ��9 ���%���K��R��:9���-gj�0�t鑔e��ex�%�\k�by���i��$���3�uD�
����à��I��[λ)~5)ҽ����<�}�Z��^��B��;Y�;Vu��j�EPYq+b$�j-�K 7�7�a�o'���vw�T\�ˋSv2�nnf��V� N4( ��,ws���d{�������Ҳ����h>w{`����/|��m>� ��8������^�9�$���gݱ���ƽۭ8���{�˫.��o��xC������	��l8��֛�R���@Lg+�GK�p:"U?)����5��k[u�:8C�:�q���ʯS�8��c���
\�S�_�L�U�S��(�L>ȧ|4{�t箮�����J��t�m�y<I�R_3�qF_��r7�,u�Tq[Ne{Q��U�^ݾ�{��U(K%��p�[|-{�h������!�B�{�&\�+�Hך]�Ob��:.*=�e��� ��.9�e�~%����B��^G�ӂQ�]$F|�:x�iLlTS�4��[����yힾ��y�29��~}'O��\N�wl��ږmA�A� �7E�䪞����WP4��Ҽ�1��Z$/�.�[��׼M�w��EjsR��l�VzOq��oJ��%�� x3�+�V��L/gz�!�MZr�������m�^{u(7�T�]� r�� n}G�)�̵z���i~Ǉp�}�D�W���W˭Ѹ��p.�8�;�`Z���hF��z�LR�x��g\�}�����W3�HܼΪµZ��WP:�r�
����d����:v�5B-��b���1ė3.k/UܵHt'S�}��w'kT�:�y�qL: Rݵ��Z栒:G-�xw3r�&]�k����}��uΞ���NB�3Z'��S6�cc�J��W��ة|v�ƕ��|�B�{���<(�^Mto���-Qiϙ2nt�ZG�t,����� ܱ�=8*T���ୌ���;R�^̽�l�[TqU�o���ÌN)I���p����t0�^r	�0�p6�/[��ѹ4ݟ1�v����4����η�Ѽg��}����s7�ٴk؝�x�=۬8�I;^���7����;��uN3�}��)�:�m �n_������O��y�>��~���"u�����v_oN�<ɻ�t�N�O�;:wj�eV���2{e 63�[�����.�>�^$̻�(���{X����?�_�O��\F���;}��ۤ�ˢ��G��=C���uF�@r_���U�ntk�q9O�!ĺ����7���(�(��Ǯe�3஦_LJ!t߅�9|�TN�R=�Ԛ��|���
�;(�9�r����Mo��i�k��e��g��j�U��Q���umU8��ɠ�;c�r�'�,��p���\=�(���%v^���-�Ś���\�I5�j� �l�w�W	��f���ru� &�CҴ����f�9[?�ӳ|��׌��bv��p��N>j
9�����E���Yߣcq3��j�u
�d�\�k�!u���~x��<�IB�D�yu�56�<	KӶ3�Y}3�r�
��S<��T��b�
N�s����(��p:m�w����TN޵��k�.�e�"���z N@��#q3O���������S�3�v<�������|]�Q�[�5GG��E���O�uR�� r��Y�lɂ�R����Ϲ��u��!O`FIh�Uޭ��9N���ՠ��F�)ճ7*��/�J� G9�]R�X��5�.�y��G��g���IQ��$[�|K8�u����f���Gc�H]p=V*%O��y�v���Z2����n��X�}F�s��{�C����$�S�p<�*��N��*!��&���3m�W<�ԭ��J���(�O,×�^���K�W���o;��J��F'AL������7�P*$�uJ��9�ީ�?���9RƅL��Z?1�)��z�G���z5:��
}=^=�bg��5K���{�E(�8N2�]�D�������v�_Ք����<�n_����pf_����17���`g�n�	����i�mƨ��C�gB�ʯ��2t��T}���p�&#(8���ce֧��F����a����,E�NI�)�Cj�]%^��CǱТ5� �N�����1Q�-��9�-MЭ�Nv����V�z�-�ȋ3��|˾\�����6�ճ�B�ݝ�v���ܸefp8/>U��9��]	MZ��!��g�U5��}��^G>n�7ؽ~gY̩�od��2�W�g���tw>�e�@:�q~3�q�����1�}�n:��02S��o���}��������g	(g,3��Ղg��d�ė�T\�ӂtϋ���z�f��Ү ��\��t��u��B��1p�ۮ;o2}+c��ܢ�+��zI�ct�A�L]L�7N@�q�� �y����Z;��H>ȧh>3x���~bwo_��t�&;*x�$��@���H(d�c��YU�����CS�F�(zz}u��b�_R��)l�oNR	��8JD�}'�H�4�n��L�ŷ�a��<a���	�[��g��'�=w#o�uh�g��PG_L��	T
�s��9�SKk�˷����pY��a��--�i/��};�f���Gc����yVLyR���O\�廞�u/�f���u����;�!_'h!����r΢nw���El*�b����n��h1�S��9�A`n�T�dã^���r[t�[�u�LD���w������?�kkZ��kkZ��mk[o�mmk[n���m��kkZ���ֵ����ֵ���[Z����[Z���孭km����km�[[Z��孭kmֶ���浵�m��kkZ�ŭ�km�K[Z���������Z�ֶ����ֶ߻[Z�����e5���ܠܭ� ?�s2}p$��8�ED"P����UR"�65H�DP�P"����2BSZ�F����`�U(Z����bR�����J�jֵ`�R��$"�T����R�IUla!""o��WZUHIUT��4�J�%��-�CmZm*��5$[��h(UM2I�RP�4B�QZT4j(���E(	[dٳP���ZF��PR��eUB �UU��fu�*�*�ŤU��J�M<   Ǩ�Cejh)�8��
��`�Dm�`�qu�Z�C��N*�
�h����EZtE*����ns�Z3Z�R�EI��$�   ���UM�s��Ct�:�w���=z(�F�(��{Ǣ�����=�   4�`���Q�   
 ;qp�@  4�x@ j���R��Km@&�ƒ�o  s�h=�m����w]��=�q]V� �i���֪���ձsn�Lr2�kUKGv�0��mһ��iJ���ݹ��S�TJ�T�̈u��  Y{C%7��k9K\����nGtU)[�]�K��(tmt\k�.����M���[v�2�n�ٰ����en���T��5�km�T������¨C�%���  ;�m�=�ѷ�һf�CY�[���!�+)��u�]����Muݪ���4���;bC��ݍ�D��i�n�  ݳku��N嶩t:uD�4��UR
��  ����˙�C�H�T�]�wNVԶ�N����kn۫n®���Q�m��m9���we:u��]��tʆ��k�vt��Wu&ꛫ�vd�B����*�E*���  ����-�붝��KXSYs�lK7]]��d-��uS;f-��`si��4�e�[�t�;W;4�t�V�n�u��:�镮��R���n���R�5���	[�  9�tғ�1�s��
�Ӯ��]m�m�]%��Ji��M�����յ[�ոY�l��V�J�����v�[;����s���]]���L�]�!���*�+u��l%J�  ܶ��GvPn��n�*ڸ���v��GC��uf�ݻm�VۦPќv�Mӭ������6��wmU;[Uۡ]�h:��9M�w)RJ��   7�U5�L�.�wT�[�]ۭ��;v�]֭ͭsD����ss�g����jݶ����t���՚R��]�Zu�l��:�d]+.�[� E?&�2�J� h��$�%  !��ɓPd�  E?�SM�ɐ�T�I�*�� h �J�UMH@2x�Hc(�%#t��W"���2�	�)� P�����\���c|��_�B����	!I�@$$?�	!I��$�	'��$ I@$$?���x��������}��j�c����JG.�&S׵x�:��*���[ε�$�(����â�Ѡճ��dϢ���!
��Z�F�c��݆��I6:��۵���N�xLfթ��((|�נKF��6��k~[f�=��O(�кh#:o�W��s��Y��E�L�Af��wB3�74[���v�P�EdٻKP����ܙW����8a��� ��Z�v����T�ˡ������h3t3~z!2���
f�kS��-�M�B�wW��*�����6���KK5К[F�8�G��+ \�finѤ�Ƞ	�Ja��-��˵YR�`��vv<��*��͎`�GP�2*�k.)�{�(wsRCl$���;����+JE�P+߶�K�u"�~��`f����yJ�ܴLѵ���p'^�7L�.�وi�'5��sr 5@��[�����oe=�L-��;w�jHš�Kn�P��:~��-�)�� E]���(K?�6}�g4�n�Р6��AQd7���\��*�j4��9���J�X�����3\'^�
���V�!�tct����~��h.D�bE�� ���^�-�(sRp�]�t!�F���,�ؕ4�!�l�j�ݤ"ғʴ�vfՌw��]��њ໶TJ��4৵wG3%!�7X�-���P�q&�v+l��^!�`�@��+. J��iD�����	ӛk-�$gH�FjSt�B��C1ݖ��h�aD6�aE���;�-]فu�[2n��ĕZ��T1�9�oȱ�g�лDX0���Xh�i�D���r5z��ˈ��bul�W��UH�����݊@=
fm�_C���?�Wd^0�[��^Iw&&��2��*��7�*�,h�@ ٸ�B� a�z�`�2f��A)�y*������Dl�����c&%-	.�A���୚���뭍�[K�zG��1)�h]�\�t6��ӂh�*($�1Qeddy����	պ���%�se��n� 7	�Y���)u���u�<�N�Bȋ��<���X)P��t�/UnY�m�Y[uj��Z{�3�dV��[��*<Wx
Q��?1�Yn�U�mX�.pvX������:R(�@��kь�s6���ޘ.;���N�v�9%�ڱ��̻�=NK�l�!��b�QS);�a�jnc���tn;�%"n�Xe��v��4�6�X�����b�E���F�:pф⑑�N�e`�h4+4tPj8�Cj�+e5t��\�y�p�� ,�^�דS�Z �uۜ:�m�2tҩ+O;-���Э�3 �LY �Z�`�xZ9��00���[�2�ݖ�v-�a���!����%�
�7p5��"䫱��t��h�Gf��fͭ��)���ʷ�daEf���9#��	��������b��]�մ�f�ܼ�O]��Q�yB�0�)1y�.��G,*u5Ի�5����4R6����lӐ�j�9iU�;X����zmD�0Lw,V�[uJ���9����J��jډi�Ʀ(`0S[����U	31ܡV��Z0�^Q�3���2%F"*�*�U�KU�}�f�G3XjV�X�wJVV&���Qܘ�PJ�TrV�R�C�E#��f]qZ��w��9YR蔆Ԏ�m+4�łtV]L0P���iX�dS�[�I��--0�`+c�ui��%n���4�rl��e+�7d(h=�)h�2�,Ձ,b�l��u��lj.��̫H�ƅ�qE��XDu�n},ډQI�XF�+��O�3 Y���3#J*tүjBn���0!R�j�7�f�>v�n�[D\,�	iV�R�&D�!�)'��n*b^Lv�:r��5�6�a���ދ��z	�ic(��-M�9M�opU�Q!KbĒ��͛E���?h��6A@�Y�4��m���j���S��YcRm�@��d\Cid�fb��p��=X>��H^y�)o��(��gf�-�ݶ0��DS���� !ܲ-�ڴrP�:�uqU�m��q�&R*�zA#Al��<�$.�(�b�@lL�VG�[�z�ʽ��Е{��u�G��&�[��a`��B�7MV,�9H�0Խߨ��)���Y����ެ�
L��oPפ(��ICf�5s��U���s��\��[;�� -��u��Zqf3�<����(B`k�n��
d��V�VMɨ��NQ�sEnl�1M�ɧ��*ل]��f&*�k�hVK&m���xU��#��B����ˬfȥw��M
����#�&Ֆ�n���Ӏ醶e�
�����4�
P9�R+wk�*a[�ɻYF�'�n��/c�@�]=ۢE�hU�j��z�dQ�l"�ަM����&�{j��71�I^�mi�b�(�����0�����Y0�H��ʷjj�h�7(c����\9�Z�G�@���G� 0G"���F�>ԢwE���@!�Ko��	�f��ʃ��z��6�{���+h�*R�u���{+�x �n3kT�za&�ߜ,%dɤk���Ͳ�^K��%Na�sJ��f� �-�ֽ6���t5�5�6�[���
S3&e����if���Ӟ�C3�`�4�W;)Xf-�ҁ���Lqn�{z��Ytko2��uv����0e��4�`��_(��e����A����#C�5-���@+�eA���fb��Ahd�0���V2MV
�E�]�e4�������ۧ��$����MV"&Pv�{�Y	fc�͙i�n�ø���m���$�*��tcYkl(䬚�7!�%K��.�p[�I:M�{a�ܖ ��'����4����`��2��U��%�hZx���;�5V���%�I8�f5�M����J���C)"������*#H6�Ë/+Uܢ�ىI��2�[�G�8�#bjw5f���6&����+u|01�Kt�*U�YO2�5,JGF�+��9W��k`P^���Vc�o�I00*R:�*�Y�&qaY��nᶤB��ұ2�(��Ֆ��d����Q�MVf��f��m�L7��ݖX7J���Œdj2���%j;Wo&��&ʩ�p˒�@A�Jm���ĝYf��DA����2m�b$�F�w��2I�c^�7N2�{i�p̬)mCt6�(˻ѵ�	�z�aVz{M��1k�(��In؎��ɗ6���Y2]Y�Q�K!�G+OIٵ�N�f�f�)Q�ɇk)�Y�hF�%/3T����X%^**�u36^��e�"H�j�cqP�m���g-LYB�jy���5�-FM�t�nn����X"5b�$O~[٬̻�W��ir+6�j����IVʦ-ZĒ����^_�i�B�/Ӛ��J�fe�gf�B��뱐��	Rá���G1���2w6���*��Q�.F�^L(^^�x��1i!܋2��gʳ0���2M5��T5b��sLt�p�,V�,�
��Z�x+qQ��p��u�cZ�N��L�eвJ�V/0$R��V*�vm����o��Ie�)pLr}�h���/ Td���Sa$���$&�#W�qA-!F��A�������'�%���&�:������cբ�m��{F`��P�J-A�ù�Dj&�:�Y��L{�R&�L,�/-exb-7,5F��,E��V�:������r��B�������͊J���V	��6uY�+ug�s3H/a2jl�n�-d�T���]�&��[���<�p<�tP5^M��
gK%�`�Y5�o�o7Su��	��cHeF�V���Ve$&ظ���w,STh\U�>:b�by�N;e͛&���p�`��#2�ň��W���޺�$��A�ܺQ�iꧩR�[�r�ZT%�(ލ�ł���������S��Z&@�m�L���ݮ��Nb����.�7Qś���Ղ@vj�"1���9�9�t�`u�o�e'5 ��]�!g@V�չ���.ec4%$M�CJ��X�*Xyj��n��mjF�[���rm�{O)�I�H�(]�sC���+bY�C��]?��X'r��C�)����X�3�� b���t�$+���>e�T4�Wh�n�Zu��B�ly��)�ʺiX���9�t�)���ͼ�i�K-�-H�����n��V�� w&^ j��⥉��q:�k3d�n�+a}��R`������e��+.��� (fb�7�¼̷v���m�`L�d��
-��`�¿��;,�i�K��-H��9��5j��i����N�O)VSm$��Q�])tM��cGY�3e�pGNf�j��
��8��29s+*���n^o6�T5���Vc�8X�)����2�;����^0%�bfޠ-�{NM�p2%ܭM�N�-�8S�;aA�q�WjC���Z���أN���r�7cIˏB�F5p;��WIc`��1�x~ʒMۨ�U���1$�ę���G̸FK�e��,h@5�V�����K4���Y�����C.�nf�z��)�q!��	��[$���t^1jTX��/@�7�<�PJQz�(֩�H�?�]o׬��� �d�j��f��mW+,���E5-�a���fQ	�	)���kI���-�I���!�ҪJ,
��-]���)��T]�.�4��Z������d�xU=ɓF+��%J�;�ڌIB�����O^���>�@бŘ�f2�^�N�Q9��@����pQ���͍���F)9���JBdR�@�w�L�/ON��Y&J��Pٹ�)��hV�m�w,�Oe�.��.��B��%��6�d4�2�4^*1a��6�!Ok+���W�@؛����;(ɉX�1`ʹ��PM3����]Zh�@Y��kX�d����vC�{�'��ҫY�+5tE��oYzS7��<�,��۽����nHwlC��	�Rw��U,^�<�C6�\{L�*"ͥ���,�T
�<oLIG��ݽRPuwl%���p�f-)6|%���wn�񆴣C7r� *��Ze��:���t�h�d�n�֌I3�-�V	���`�V8jVo�e�X2M��7�jI�N�쬫���)��R"���Z�X�aX?Y�j��I$l�v۸ɳBm&8��M��d��ݳ,4��wEL�c&B��X0S��m���%��6ZNZ8�CKh_�A���kq��E!vw3�,��V�`QT��ڻȥ$Uc�,C(|�n�+�a�2���x@�����ʩh���/(xkp��`�Œ��^5u&&�!Ix�o�WB�P�ic�{�(X
��Ym���&tH �ӷ��m,�M
�ؔ�X2pd�n9��9���	��h>�X%F��'�5��w	�(7���7`���F�p�-�j�=�t���ԕ8�h&�M��mY��9L�S�T�lC�iMQb�csQ��8��¾ĥ�jҩj尷@Ci��t��H5��n�4-��MS�����(D�:�[f��P;���M��v�^=�	�lˁZ������b�.�J���n[j"ڛcDN�ƚ�2*+.ڴ��ԑS����Rr`�4�qa����õ.-V�{�RQenGa�%�cQQ�h7{F�Ϛe�5M�X6Z�,�	'���9��`�uAZ��,a�v��{��&��]�
�ϗ���#*���q��'yKʙ����k]�&Z+X��W�n�']��l��MHw/��N�m������}��Aj��+=UU$0I�5c�6�4�5��U���n=
�\��+�e�y��E�z�"��A��]-c�<A�J7w/�D�2� �bD����)��a��hF�� �v��	ԩIC��fһ�UV%�4�Pɫ1ax�=T�ɏ�&%���N����m����G6[#pi�V��eV����YB�)^oMWMhZ�cDq��Mk���{(�3㶁ևŉ�S�2��su_ѹ���^ op��a��[MFԻyj��ee��*�Ƽ�byiR䙂�T��C/���f��/m�9H��W6���Ǭ���%4��x�tƠU)�Ed�D�sK�Z^��֢�*<��{c3,�(�����	��*l:��i��j���� q�1Di�2�޼�;�"� Ʈc��7�6��b�pR3R"n��؃w,en]���`�ޫ�-����&��ӡY��N�R�v)�E�b7���ǹl�9C*h��Pui;4.�j21�����@�1L��d�>:(⡭61��E	(7s²���ž ���X	�2&��Z�b�/A���H�A�2�+�e���^�,�V��2!���% ʵ��F!��ϡ*H��(R��]���i�@��&;n��\~[�	{�V뱪!j�������9��U[!)� ���6��T�����I�j�3�ֲ��CX�kR���\��ۙj�4����Ax��b݋;je��L����p �F���#S��%n[	La�GM]��5��U+V�Z��u ���խ��B�d�Xd&-ݭCpJ%�K���6�?�^B�ň�X�%j�Jͭ3E��94�P{�Y�۲��ڬQ��kEAu��`R�]%���U��l����LV,Ӎ%n޺�f���$��S,�,�.%"M^"v쁂��$���
 AC��Ѭ�Z�Ϳ�h���)R���QSN+*�e�X��gp�*Z4Y�4*�{J�+ �4SE��B�Xo3�D!V�$:j�+rM#-"u���E�Ѳ�)`D3{�F�+�D�$�$C	�U�#8t	v��{�mԤ�cK�5��Z��}@�zs��D���[�¤޺*j蹇J^^�Cfs�Z.N�����c���inؾ0��:}ܞ�Z�| ����:^�F�%�gN�1��zf������3����I��C��,� �(a�:C�!"���k��$�|�����5����SV����S钸�z�w.{���	��+˛�p����YJ��ҋY+@'�j.=�����ݵ�mx�����\�Y�^d-evӇ�nd�뷨r*Tj�pr�V������%X��)s�*��N��YgQ�[�w�H��;����-�7�t�d���}�i���Ӯ^
3���0����}�y�;q:{����ږM{wO����F*s41�_gQ������ge��@��9w+{VXH,X[�W�:�b)�k��Z^��Yc�r:i�k��9�c�K�D�=���mҤ�V*���!b��g\��� �U�t;��N���A�ݜ��λ�ܴ�S�`����j�W"�)�89�p�u5��i����^7̞�\�M�!��qPG3(}�݊w��u�ͬ����D+,��sY��d��܂ȶ8_R�lKf�"�N�+	6��K8QY�D&��e��ת�m�;�V��h��&ovj%�99]q��^=Sd�]vvWB����/�,7�"1:`���:t�l\���p�4�>��Y���D����Î�xN�Z����dv4�����A���ͥFf�kR�9�	v_Da/s�ҫ�R�[�AڌW3x��)�k�O+c	�����ϯ4�`������ۤN�tԴT+�9�ܮ�4�j�0�+e/�dS����ͤ�	橨Ω��{�B�]�3MB��B]^�\H�Au�F�b��z��5Q�e5�d�r�<�;�}D�˩:�M�D�i���g6��`��K)q.�u�k���z��f�V�U��R��D6���s'Xhkvq�Lo�y
\��wZ�v�+���d���ɔ��������s¨�<��9|��j���`m�9�oE�i\y��n��LV��z�V��#z���6`�Ȟ70
�,PD2
-k��άVnmΡ��|\Vv�� �� 79�_ƅ����E�ò�a��e5^��7�"����'r���h�;�龜f��a�1��F&���*�����w���5�K(l���<���K6����z\�dE��m��[D��ڥ���v��v`8�$������5���4�=��L�,}GP�F��o=k�r���J��D@a�]R�؝�
f���'I�Y�n�=��f`R����w8 �EK�|¶v9�Ԙ�2�"��PO:�z<}�T�\���W��G���7`f8h��~�Vͺ�@a�8�&���b�"��!��E���~Grm�,���5�=�f��
�On�[�$wtLb�^nsSx�N�ڥX�e�K=݇�����Vc�@�� ����n�ި����6gB��C��zÎʑM���o��O#��,u��;�=��t�WH�Z���r5X�e����sD���}y���d�Q�!5[G��ƶ��~oiyxg+���c�r]4cⲗ9�r{�4��A:�Nt�6aP�c-[���\	�q�L�;�*lRM+t�]j
��af�L5�A��Wι���۷r�ԫs���ʹ
@"6���(9��[�U�|�V�ʘ
����gt2�G��evD&��8i�]ܖ�QH�rf��\�{(kU�	�'lt]:�h�̮�j�`���-V��q���!Q �F�viǝ�z����8.���6��\�uSSQ,�R+lo.Z����k9>Ô��pVV���pXsU�pA6	�2s�x!�'\�1gLE��8�t�@�W�kn���+���sK�bޛpֈ���}�tݡ)��o{�A��c-gU�Y��79�	��|��D����&�6ǫ�
��iɬ��7
I�U�����o��:��x6n2*�1u���M��[G
���˝6gN셝��� T����5�z��(B.�J��V�CzysUՃ6��,�aw��.���
�=�ק�&e���� �V���tp��r.̭��/���؛�e�ĥ/�*B%�ч����S�ށҲ������c8�@ƴ�/`�T��@�=N!�h4�Z�+jǆ���(>�1bTD�C�$���Vs�u�j�/Npa���'�%+EC#�7�'
2.餮�u�\+����Jtb�5�I�{��Kn���F[����C�=x:ӟ��ڧ���q1bp��ދ��L{S Yܛ�KN��j°%J������/�g�^�S��t��*C���U,Hn纕bFrl��8�R��^�X���;�pq�}����H��E�8��Ťf�1ݱ`#��,;}W�Yٷ8M	�7��8 ��'�.aQ��뜺��@��QH��Q�gT�X"+x��&'�V_|p;�+�Օ�R[��y:���bIt�b�iI�kTXWm��w)�el-���٥�Z�U����W,+]^^.�7�i�J�0�_N sY��e��/��N�dhl.�و���ӑ.[Tf�����v�
4��&n�x��\��3�خS�l:f��N�!qN�ar*}:��$��S9�]d��˦3�
�	����]_c�7���v��l�D�_=�xY3ss2eqeN�ue���l5X;�g]�V�PNå<ݽP[+iQn8/���ڐ9��A�]�m&�����mgq�׾ikp�0=cL5��:�����1:st��Q��Y[��?
��h�*ǵ�!o�9�w��#�L��)"Γ���jT�ti4o�Zh�pq���6����Y���-_.���0���6��}�RL-&�����i��3��������p�љ����M(9�g%����
x�b*�F��&Y�؏j�6��߂��u@r��*��)ϒ mةZI��o9N����*ʮ�f���Y&�peE_Un�β����O���]K@��i���+��V�m|�T�T!�]�+M��QŶB�O�(.�{���g���{b,�K���_T��E�o#5����M�$$�X�&��A|�q��RgG��g�Pͼg*�*>�if'@���\0����aQ��Oyl�U=׫7{����j�q�XaQ^�(!)�:���gY��:�l�Kf��J��#�Y}�:z���r��ܫH��:ժ����5�:5�)�ꋏ��ʎ��iU�����甪c����@Z�����T폆�,^�]�]]h ��^,�Z��`<����a�ڻ��/�EM)Q���g�A1�3J<�`|����̓�v��ư�_�9WH�"��R�����S�K�����^�� 첔��9�;�[�+��G��VF�iC����;%"�T%�P�M�$�c��ξ�Q�b�p<�*�%�/����Z��$�R�c6��c)�q�z򰈕��o�f:�'{�%G]D]�����D˕�
�F9[�-��l�u]�jU���Z�6R�m�p�VѷS�J��fRj,��b7���6/ ΰI��w��]��ޖH�Ogr�$v�'vj6���ZtۺS���maPi=��2��E�D�*&�I�Dv�hR�qs�W���7qf=*�����~�x�Y8U�t4��lQ)���K9}t��KjT�w]ud�I2r�s#!�ǧlYP����2�s��E��vZ�:�;]o��^Y�z�h:-�n��2�V�:��{j�%��:��7ܳ�q"��M�n��{ɽѼh� ���0)��}yY�60b[��\���
�<�z^t7&g-E*��
���5�ZpŹwE�v/ywa)�����;}:�M���.
u�r��׵��Y1�Z\����\��`#:��0�|1u���>�HV���a�Ut.����0̨3ò���ݔ"�����'tS�K;r&���6>���!���p5K�;��4���f�D��q�r�L��a�UD �V�}q�޹9gwe�sf*<�(�Ω8�*4��{�R�x�Q���屨u0�b7���gEh[0W�`SV�9VѺ9Οm:��WLn>�p�p]k
�D��H����t������ mv�;�y!@n`\�rh̨�Ae�n��L��� ��.&wֺjZ��AZ����>���Z��XQ��<qa	[Y��ś����`O'�)W,�����KnZ�{��Z����^��n�7t�7n��aX|��7��4�%����e�'C���H.�y�+��z򖥕���ڍ��ԝ�}`0h�}�9��&���6��*��9+U��n��.��:���N���f��R�r�5�f�G�-P��˗Z�A!ye�f�HɣP���a�Ʉ0<�R�������񡗔���Ԁz�)�M%�u�s:۷I63�pS#��ԇU�`�VS1�GYS�'6�Z�wGM\_a���E��K	��p�I�#��,�hlŕ+�t�J��Mˤ;��^�A����q���z�Y{�@�@Ȱb�`�޴��Z���̡-�4��k˷�j���<��@QL��sA}W�u�P��S�ȳ��E��/\$��enl��V_R�)�i�F�8V�X���X��h��pT�Dv�C=Now]䗨���װ���ː�A�h��К�:��!dV+z�ː\=�Ͱ���u0�q˭�LS[�V�gmL������ϭ���t�c����9y�|�_25c.�k�r��es�^�E�t�ӿ8݋��\�(�s�
WuE�U��81��D�˛\B�Lx��B������\�`��5�$׻\��i�`�ySDE'�[E�>�Ĺ�J;y�c�٣,��<�+�${��v�}̈�%R17o����Ɏ��ng61���x&�Z#8fAa� �a�\�l#8�6�
3��Z�n_^5'���Jl;G'�6(���X�xnlU����m���֪J�)RWkq<W/Mx�p����N�F�L<��3rc��J5ʁ��ϕ���E팧�� w�3�̕��降��	ƻUo,B���2���9�E�����n��R.�A��.�ȫ!ĸa�8�켽EK�v3Z���]�$�t�rr���TU;Ƭ�CA��w�oW�9+�}]S�f�����>�&<8�Z���1�0�]דM2x��42�}�P���t��f�IB:X��+��޽'���t����,�+y�E���D`�!�Y�-�2��Ò����u)���s��+�-V��|���g�lR��4Xc����;˧8X����u���F��f��l�ܶ�.��9Ε%m�9��+O'[֨�EhY�4�����B'�63:�ݺ<`��m&���"6�)�Q�9%���������������d%H������W?��	�����nb�,<2��u�q]��Eka�[�)��+L{���ݍ��m�k�h�ɺ���D�͂Tך���Y�Β<���[7Y�n���*�t�q��`����MX�oq�@*t�/��\��o�	�ĩ��Zw�í���);뫄��=ǡ��c�C����o�������vVq�ԯn��x�E�����Z�Ӈ=�v9���Nub��[W����eh����<-i�&��*�o�ӓm�Xsp�W=Y���Y�8eg�Z��iw
LL�P�&
�ˣ�^'�a����v���3Y�)sȀWi�Vq�<_3�\�1�
����G�ĥg��l,���jU��E�eh�ᡗSNd�T�;;���^��e�D:�l�gHi.A^R#��٩��s#}+�q���Ҡ:��/�4�P{
�{���]�Br�sf�ma����R1�.=�Y�[��TdҺ�6]��p�Zy{�)Z�nTi��*�[�Dq���ը��Ƭ�`���;Ҍޙ����QV�)��[an��������B��ޙ�B�������ژʭ�l�םP]kh�j7;t�W�v]�AAwOxN��01��(�أ�7�!�����B���M�q֏h>6,M�/��[�R��7��S8}sM���/p�=t&%�:�������B�����:p�Ys�)�W��\E�^��WSD�Z�u؄�����e�WS7����h82$Ճ{a��EÃ}5�c:���o2�Π����4�[$e=�]���\w	Հ�T��!�7:���(�p,&Z� �:��g-�.8��bB,ƫ�gX��<�m�)��ٰ��t�Ԣ;¦�r,fΣq�(��i N���L��j8l���``�O��:����A��^�]���@���"����SeB޽>X���e�7�o�).x��Y3/�#��8�JBu���B|&��}i�:�ޓz���k�6��P�|�[�o,�8�xSM��|I�S6%��E1rY]�/��]YO��7��)#yPS�hAy&;vi�m�@���Z�D�bWm��[�u�����3��������G��'_(���4�ș\Ȕ�>�:wi�(�b
�b���<Չaf�dyGQdr'x=Χ
���\[��Q�Sh֑�[W��Lq8���;������-i/���-�1���oa�9�apk��qT$�#/����ܷ����{#���1��2g-��`]���>��m� ݙc�u�s+Vb+���}��R��ؕ+0�G�"�(�;�-�҄]�bnN6���*�o339T��`掻���z��e+]����W�vo�����N¥�1�lMB��k���8���x{�n)u��+�WS�{�Yϔi�������^��it�yB]�b	i컘-�ݲM�33�J�N32��NξWr���%�u܉���t��|�P�o���K�	޺#���v����Y[�96R���_p�:��{����� @�����>��;�����Y7�3e�f�ٕ�!�6Ƽ�T/M��&�6d��Ji��[+,7_6^�I	F��Ύb��Wې��K*�6���5aY��&ۡ�.���t��@�>`D[Q�ui��םf�.ꆠ�;��X*��ޔ���lN���.�/L�7jաB�5	�`�e|��	���3b�t�X^�D�e�[Y�����Ӕ���W*�,P(��q����z��篯,��'8�KCs���}ح*��V68�l�M\�go�B�K���h�s-�����xOkI���,���Q1O�_ �n�Z�g=�j�X��xUϸ�p�eVaw�t{�,#�%Ȇ)_8)j�m�t�/��ʸ_X��c����\۴S��)]>�N�@Ԇ� �nں���on��-Uu%4�R��Xy!Y*�{y����v�3Yr��:��]^n}�i!4-Wn�@@8�i�q�v���/2�t��v>3c�^:���A6���AYW��^��&�am�Y�wPz¡ά_�G�ff�̙T�^�������.+���4HR�-�G�s���.���mM���z�N�Vbn��k��^k��Yjj�M�od�7)�cSS� BYll��n��.ź�-�;*���F�-�%�pn�V�s�����z�����kr�	O�.���a�޽iY\�$�8�g\���*�:���&(8񜱱J�|.º���]4�9�nd=r�\]z�Z�s�3c�b �J+e�K�OnwWnO�g72�MЭ��]v�\d�ɑ���� �:�_;��v鵀T�����%g`@.A���R�����6
�ٺ��-�r�(\��f���-�|{r�Jq���u�p22�v��w��5ӝ[��&���.���ը��Y�݉�#��
!j*��ڛk�O
��vS��`�)�ƍ��)�0q��p@;�K��&D����ᵪ���L �cĵv��w�X؝քX�d������֞�k�5�}c�z�<�lc����;��j�X@kE�O4�Q��[���ݵ,�!3(�����Gc��7�5y������5+�B2��t��L�U�����U)�o.��C����w(
2����w��Yg8���}t���nKm�m�0�Vv�6�]H=ϋ��*�1,|-�(o\y�n(f�&;��݅��޶��e�e^�Σ�H5���ҳ0V�����c����K���;lU�B��nꈣ��Jf��t`�ZZ�b�R35j��嚥��I�����S}w@�ẕLK��4b����w�.�c�K��P��!�Sߍ,�����f�ܧʲ���TMC������΅^Hq�u�ˬ�֧�;�;���,4�'�+�.�]qw�o;�.�b��a;a��A�hl��ll���}4H��$
�ૌ:���۫��P��\���BXC�C+�o$P�Xrhc]l�ݾ׳'��l]8�,#mG7���L.�|�4����t8i�'�*+ݲ��$�t .��lH7T�b��U�u��*��6�>1�p�j:���u5����p�U�%�H�Y=����Q�qlޟ,wρ�%pL�%�d�r�{d�vl�[E��� ���Ʊ�����I��|]'��X�̫�_�;�	�G��!�Ś(��kw(�uw�X	d�&��B�}�D�b�Y������������']v�F���ءν48e�B���먞�y������clwpή�4{�3��ru���W�{%h5o�>�ϟU�Ms9����˝ �2�F0�fe\b��4��r����K(XYt�l�g0tV�am.D��Yyz���;�Hz�r��tz��J+v�]_��\;QU�+8�~�>]Fu�kugU搎J�"�zXCy�����f�e��f��LTa�H��c���0��
|k4�l���)Q=�ۏKjձ�#smڽ7��΄��S9j�ЧH�̫(�K0a�f�]�y"�Ƅ���͛�P*�1�l�2��6Ng	j��Y1S����ɚ��%tμ[��
4�)b5/���";7�i��C"�s�^����,2���#Tk k���ڑ�s5��+�]��m��/6�n^B����n��چ'S�)��Ν��ҥXtw>�f-�귚2����\f�J�3)̾�{��Fس@e�{�������h��ҳ y\�g�ė���ڂ;p�!E�wtf�i��m\�q����+�^�݌�ެ�s��J44�7+~�o�^k���l;�0�ۺp�i7Y;LG�egd�A���EW�����9f���Gv�g��m-�Y�KY�s������k�����ep;��:o3�F� ��xx��\l��]f]�:+~�:[w�
ݸ�&Xރ A͛��V1�9���X�ȝ>�a�}��R��naux��J��4�"U7(���:l�Y��Ô�Yo�;�9C�j�0]7�:��K;���#����{hG�N�d�S��{c2�I�Υ����m5s���W�b�r��g�vWM�z��ʙ��uʺ���p�c+��N���Z�U��c��N���]��tGڽ̉�� V�r(�ι����JVU���"��֫UA+�0>,�Y���Yh:��m�0>"-�6��ݥ&�{)R�Y�P��ֱ4"?B�n��th�3y%�u���$��Ã����膲*mQV຿��v�����u�#ԗS8��Uu�H��V'��P���dN�jf����Ɨ-��k������ժ�\��ܛ�<���ڒ�l���>�8�b���deA$�Le�XL�[�+���$m�$;�-w:�T[{b�f��oI��[�krNo��2�*G2�Գ-W&y��C֛��L�7��I	���S�0�F5�Z������rj� w,e������m$Z\��(�y���8
%�]�Jn쌳֯���Ӻ�Vi��ΨI��Q����ZX�j��í��n�s����y�(��*�˵/71&`^�
�	�;��K \���v��P�Xn �6�k��'x)i���Dy'�5��;��B���'jA�����Q#Cn���W)n� �.�}M�
[��w���\c��Gt�_-`aV���GҞn|I<��O	qB"�4k�vV[{��Y��_'�)��r^�[��>Өc�g�h#A���]-��K�o��:�j4)q۝�#�gb�W���@*�d��Ns]����ej=��_���ʙ1C8�D����?q�l�ս�^�[�-m��/�����rc���Vo� ��$:�w�0R��R�gJ��gBXN�hW.�*a���Dqt��t�\�p��6�����\�Aa�9f�p�5)���c�x��{YcF��֩�:Z_Lp��z�J�ܓ�E��P;�r���m���S��\�@t�p���V�"4�s;���8+i�|���:�$>��4v��*[M-u�)�l�t��[ug�lu��"�,[���1/h�D��z��۫v�Z��ɛ5'�Y�����b���Ɲr�`�U`�{U�c<��2ذͤ/�#�5ѡ�a����[�����+/IԨ-�P�k�6 5�� ۡk/_�xn��f�״)a��pIq\\����N�W8v#o�����۵1�?uhT�`�|�8�$��ŌMJ�NL�˄�ɗO��M����d��R�gk�������ب]rȲ�=�4ҝ���L�)�ֽy��]��G<�V��kK�E�gO^S{���C�1|gToT��YJy���")����V�3�!�2�_8�I�qD�i�WL�D�R~
���	�O�*��N���j�2K�e�8źP{M�b�b[XNk��r��z;q�F���߯�3}�4[�I�]��i�k����� �!���/,u�Y�nv���;�E������kr�3�W`}IS��1É1$�rU�@wie�gL�W�^_(�)"K�NY�����4�kLm�5��1>N�2+��6����^��}o�K���9�1�����O�z1f�H.�7���X��+��l��V��}�����c5n�WX$�f]�4�G��p�d�n�����	g��ܤI��
<��ذ��e��j��(i��Մ4/��32�,�	#��5?�+��.��T�PrN5&r�X�s�'yt����p�Sؐ��f�t���-�.:�m���{$����/飯��+5� �S�9W3bM��4�.J��!0�j�tĥ��n�z���&c�xb۔�N�s��(*���=�f�u���f܄���t��2��
/���i�/FQ�7�.-�݆�)o3� F
oR�c|-��;W�;΃���@�I�U���*v�\�w����m�wxQJ��C�af-�L�v9�G��{uZʍ�p"�O-oN��U|��#��I��\�@�dK���P��*����L��cg�o��F����vl�輢��15Z��)Ҍ�5�G뷮�J��Y֩n:�)���Fܙ�r|]��T�(Sd�_h'4A�r1��7���z��-e2N�ݿ;����� [so+�u�sr��>j�3C9	�p5b5�gvw>�9���7�]��vY*�%ظ�cF�˗�\bnn볙AA2��@]7�f�u;)RW��ȥȵ�X�y���#�R+��@���[���-M�"jC�������9;؉da��!:�i��r�Hue6o6L�ek�9t�Vr��u �۳��GM��]˰)�*��\��\kO�Z����
�d/@7vu��R8��Sp�]��!��X�����a�_K�����SӶO�������Y�LʰM]g5�������-F�\]t!}��+!G7k��]Y�7��3���W����EE[R����H�i��pAWÝ�!͵�v������]*��AL�P펻)Iˎ�.�@�vGoQ�-�������D���e@IA?W��W��Sr��׬)��_7Õ��f����� �Y�����3t����2n��.�r�#�҃,�u</-`�ur��R������:��lKɊ�������e&�oF�3Vm��v�|�32� F��V3�l��Z.�8�kl<Ok��MݾۼG,�I����@wV��c%-Sz��ь�C2Έ��)�:�J�Dv����95gS���Lb�v_d�ب_N�	F�Ec�����T�z�R}�v�:�tl�����t̶�ٝn�j��hpe���۷\���T0p���ܰiU����'�+�շn�̲�!cv�&�,����{�i���J(݅*��׍ �I[b5�2���n��"��T7I���}	g`ќ:��8���3�۰#u�uj9�'u��!�)�`�����]ܸޫ�9-���odfi�/m\#���{I�1Y���5����b�f�5�w�����cKlgn�D�%x/ �'n@��W!���W�y}v�}�Z+nmhN�kQ4�ajޡ�ǝV�8�i�q�fFm��u6���^��5�s��8�,��n�N��,�
щ�}yڗ
)j�]x����*שP�s��z� �l���*  �tHQmf�l:�鼁@�ֿ�-͆6{�a�eF2BD��V�Z��*�gˮ�qQz��]�/��%������>���atغ�̝d>gTx�eY����7���:γX�\��SӏP�̮�)�.�aH�fq4f��ۼrĴ�z@��m�C9�+����v�e�A�#dM��ޕw�rN�_�r�ݻV�ytkq�\aG���dWJ2N 挢_YY��8�8���{�֞���q���:j=$8+S��>Ӛ��Y]�*�1)P�
��Hӎ� ���_a+�R��[]�+�B��+t�:��/E�Cw'q�OG|�FA��ތ�8u;!���G ܮ��8އ���ܥ�K4�؞sa.�Q�Vf���D>q�3��x�s�w�ܖ�K1��v	��֬�F�=g��K;�^��g
�UD({+��u���5�/0��s5z�=ގ�@幽V��+/��f��,bԑ��ܱB���2V����b��يh�'��5-�%�aodB���R�JQ0�ZiX�F�7��/T+�=�ܮ�԰3��[W(}lZ�ƝM�G4H�����}�;س���j�ac������m߫�u���D�;.��\`�5��̲����20���'Z7�擽���[�b	\OJ[gN	3��A�4�|�k5:.���8�l�ͅK�ҸgU`0�>a��I�M��7��;MQݽ/xՠbQD�r�!ZMw=�w5%�OM�NSG����t�y��!�ۈ
���C�w��Cx�g�؂�s���,�ҰI�˫N��O��&7Kj�kK\b�TqZ���)���a�]yec 1�J�-�k�#�����7x��c�yc�e�wʕ* �����X�2�oR{�|��ib�wU��nʽ�_Z�i>Ǔ����������ƻ��"��*v]�H� ��]�]�L1�]�ճz���fHB�C1e��I)gwv���"�����ߔ�8Q��Z�p��K�|��]�O9��.W|��害j̒<x�&�3\�Rj�U�gK�A�&����sNR�V�#��ͫ�M;`؇3�j悥�b�����ن��읛�ZQ�bv���ou�5�)�>ce��x/:�b�K;�ԭ� �y�6��x�O9�鵄(����N�pQ��b�R�s���ݻUk��	�#vAr�S;�nS}�&���.�"cdFD����Fc1.��R���0T�H��I���[�`���y�m�ˬu�Nȭn�p]Z�Sw�t׽�.����Zf�,CŻy	{�g��1��5l%0\��qe1M�(�.�T|�Sfj9�m�E?w�}��꯾���H��@�7L��%fJ�m˶lM1Y�z�d����HIiP�_YZ9�N>L��F��.B�Yӥ?��|Ot';x9�������\��nu6ބ#=|X� ���:�8��H�y���6��}f*B�v9+{L�/[bKGq�o��L���/b뤑"�m��Q��ZnK�S�qŋ�*䛸8h�c�e� q�O�Q�%M������.	]���Fw\�dM�7�O�6��:�W���3:��ڝ��g1J�g��OuM�	�������5�����u�t6H����ՆL��P��wfNK�:�%����imk�[��c.�͡�ڂJ]tdܠp��yՏ��Tjg4�t�]��j��*%�����ؾwst��!td���Xt�=�����o*��Rgn���{�X���0w.�-�i���������֣]�Y/2�
s�M�v��}�[\�j��U�"nXɮ̵�x����aO\\���۹j��Auv��� ��G�z!8���>��]b��),}�bñk%rZ��O$LJ�{��fl*�Ǧ��m�rm������uY�x���ݺ��2��)tY}/���)$�m��8eԆ�c���wi+KI�H㼛ׅ��P@v�b���/��l��y��U��m�k!e�>����gN%xR�}XeR�K�z��l��g:a��%J��H�X�Km���e
%V+Z���Q�P����Im�Kk-B�ڶ�Q��b�X��V��ԥR��`�ֵ-�V�`�V ����b��V@m%J�E�@m����J�V�ڕ*J�XU���%DB�J��[kF��cDm-*��Z�YmE*�-����R�m-�iV�b���im���QEY*�Q-�F�E
��
�F�ĕ��4�P*(�P�j�DH��F����U�l��KT`ԢֵZ���VT�ʅdZ��*���l�VԴV
�b��V�֭Z,PUm
֕��QPe�*4�Z���[lJʂ0m�,J�ث�����[A�k
�U,D-����bȰ�UQ[KK[J ƴb�ج[D�+P�ATR�%J���E@XTmb�U �k*�Z��[F�kc#j�)j¡V#iieb"���*��)A*QmQ�j�b2�e`-B6մ�%R�l*VT�
��3�W5ʻ��\��ZH}bZ+)p�n��3W4o�*�Dp%�����M}*�嬀���U��ԩ7.�q�����ԗLƛ�*x����ݳq��ƻ��}u
����p�!�m,�?f�9��������Ѯ�s7�yM|��;Zj�X�x��½\:���曞���v�N`�����95K�,ӡ�U3ښݘ��ms"o�b�6Z��x��xE�07�B�N���P$ە���C�c��[��5=T�u���P�B�w��{����`�t��,zc�s�}<�t�r���f��e/���Qu�R��J��}����)CO�GK^���zmL��ؼc�Ȼ�k�\���z���l�Ee���ަX�hͶ���M��"�vJ�G�]=���^ג�j6��?Gi�5��o=c�DuLƶA����[�+h�)_��<�g��ܩ�v�����o�����a�؞�;qQ~	�^�K9����.)�<�q�����[��~ξ�.�Yi��wRg����։� �
h�GO��1�%G�����VsS;�47�xড়+ːj�{�&��Qv��H�fw3����`o;�_R�"��e���6ݏ+{f��={��U��k��`�Ul鏩�ȫ93$�y�n��
�rگ��]e^�sa�H浮��靵Փ<e�K=@�yK�g��_�!�|��j�֪��/��t~�5gF?{0�OKr�#�*ǥ'�k��9ófyf��K��fq3m�+؞�벧vI�zw�����ɢ]<޵T���z�iT�SQ�c�������V�y�P�mW��|�x����;ؾ����&^}3R��p׼*w����s-���bQ�5�w��-o�����S���^΍u�Ȇ��֬����{����+��|/����޵V��t�{u�;�����Uut��oc��O�bB��v�w�q�*���t�Tw�xcw|�u�r���G٘�yn���4��x[�S)�uv�ǧ%�~W���}<����N��v�����@��҅��t�@�.���to��/�3��vK�f��+ q�/O=�".�y{Lv�|���N��Z�-�k���k����+v\�4���Oq��8�3�?�̧�q�lr�;$���͑�t�}��\)��p�-8Z�V)N����v�J�,��۽Yg���0�|�1���.R,m��5o_,�s�s���١V��c����nz�|�X��V��f�^4��:/�{�h��z�sO:��G�=E�lb{���v�Wʉ���W�/�{��挧��k�Y��k�׳�ҿs_�9����D�V��x�K��9}~�k�����չ�g�������:U�y����g_<j5��y�����J��tY�ݳ|ԝ�V���^��Q�-:5z��nݒ66L;�1?	������C�s�w-�������;<Cz�ra1�p�޽�u��p��<�6��s�&l�;9���}�hK��%K�u.j�{�'Z�q�L~�������y<_��53g��;���C���g5����\[�y�ES��E&.C8��L��{����K9�_\�ݍ�q���HNb��+:��nXז��� �e��^�=���r����s�&���q��ӛ|��Kl�(�'�n5g���u���}/L�5���L��}WD/����Y��&kT�����!W��`{72�	
�
��ʍn�=Nu�w��-�P�M�]��\*k���r�w����f��OJ�])o.���B�����E�Z���;�p���v�x�1���5��ݛy{~r.�s7�yQS8E��he������tg������v��q���"}���t�@��95}/�g�E][!׾��\7s�z�õ��[��9}�ܳ_{��Hd�[ z�+�󘣆����(&\�z|Q�\J���g�q�g����%1�{�n�y��l��(zu�@k�d�;.�7�����:ͩ�޴���>������zV$�����o�r��ڇ>��_����w7���i�ڔUr򧽨u"�Շv����E(}�{'n5�a�G�{��mV�}��Gl�n�XO�;lG|��̗��+��ok���>�k2�ǳ\�\~���5��a�|e95E�ɑLz}�����Y���=�=q|\����o=�U);K���џ�Cx���2�e�V������9ΞZ��3X�� V���E��O̎�|��D�����ٵ3�Z�mH(Ȉ���U�U�P�+��YD�B~2�v�Z.J��[��U�ν7�:���S�9f�ZΙգ*�3i�I	w�LU"��GF7���f&�]�����]n�l?����?�kcCK}��V�`Z�x�/_���u��|{܏;��>���	�����I�[<���ԝ�o�y�딪�?]NU�&�=�A��Գu{;1%seil�l�z�������S�Z��_��U��5��;h���Y-��tf�g��;�JN��c�wt�c�x���ޱ��h?�Zܞӹ�qٝ|T����A�C}P��r{�{�K�WF��̅Snx�^�^W���s�2�)s�-k<l1層���5|�]���O�s�jA{J�����3ug�~�8��k�z�B�pߟ�s�\U�L��
�:�mW�֮�Y��o3s�v�W�2�t;���R��
���=�3w`L<Vj|C{�$y��/R���N<��R��g�^2���Q���b��#��|i�QY���*-O0�ʺ(/n���Y�׌��2 ��j�KB���Gj%fǿ/�&RgZ}��}L���/,�z�*�~��R77��%�smNw�w��u���f7�0|6�e�[��,��f��Lhٕ��!n�]C�]�c�{y��M�U��{�k�\���{O�f�)Ee_?V]�b�s���(�b���Uw��O?V���������|��^�6��f��4���]�g�@�����gCF�.�>\=H�z����&w���Ͻ��o(�vaZ�瞒���78OEW��,�^�K9����.)�c�ě J���V�r�=W�=���ʹ�>z�[_��8�׿Q�׿r�.�J���R+&�j����Z^���dz���/���-��֪����qA��im��e�lx���>y6�s�UN�ʝ���bu]�5FN~�c�ז4�[��]��|get�u\��.gg�&w�}��EgӮT��ݡ8��y�k�r{���4�x��������9�}rL���W?T�5�^o#C<�ٹ�5��� g�9k���ik�c�~§�fg�x�+����km�m<�-�M�f��h$��7�'8��Vg#s0,y�x����
��mu�mQۦxʹr�Qq+%�5_��)��rr��۝��İ�����v� #:�-���9L.`����{�.��-�`�����̾��i7x�6��$Wl!����Ӛ��Mga��2��#���^������]n��ʏ�U���\��QDx��5d�s�u��{/**g��7{-[�?VA���v�
�K�tJ����"�}�ͺ�?V��z�s�g�N�^�/sǧ���+t�wg����U��Ԫ��פ�t�t�@�.��1�rmunW�]�8ׅ�>�����~�;��o���zP��1���YKŀy�����e�Ew3��Զ̙��/\yU�J��ϥy=�{乽ͫŕ(]{~O�,�)���ꯦ^'Pz�Yu��[�C��(;�AtY��K���y-@�y%��}�bV�sy�.�\��)�W�A��|Wz���Uj[�75�;g��k�Y�w˳�-�)�;}JN��<ؼG.#8_���U}ˏ�θ��O��V���	��\�̞ɡ�s�����uK�����+z�vz�i�@3]ц��b�j ���V`�����2Vl��ߏ����(�Ʉh�9&#|g)`�� �D��ޏ#���:��I��o�r�*��܆X���WOn�ɪ>4��3��H�ܬ7B�Z���۾�#�۝Y����gtv��]�ͬ̕}^�]��9�c���ٕA�y4yC����\q*˭��.�mx�&�hU����k�w���c�짡�<޵noc��x m����;�u��=+�5꿌͠��Q����'u�xu��z�)��,�+^��������S�]���t��-�U�?tx�gG\/->�֤��g{��sbqu�/~���9�]Z��f�sϏ����?6�W{Ϣ��K݄t�}��y{~r.��yT����.���{,={�{��O�ۧ��5w56�������)�ͺ�?VӓaW<ψ�]�'���L��5�>�xf{���._�{��HT�Ҫ�=�{7�_�+��A�9ȻdQ���|=
5�w=������&��{{G+W�yk����O�!�fQ/P�{���//У��Z��i,��׻.�r�
�G:@3�nS����qqt��8B{Oµq��`���4&h��ak��~�fR
x���>��SV�m���wY{Qq%:�+��F_
����V���F����ek�mQ���s�N���Q�d��5W�c��w�쁇��]õ7�%�׺��7׼�;�$��A̱��Ee_/k��Y�F�}��nw�ə浭�z�/G�{��OuU9�ܝ�mVo%�~�sR��P��]��o��>y}J��«�5��+\{�5�վ�g�䷋����c=�=n#<�����t���\k�̞ɼ��U��l�T>;�%9Lo�^�϶p^�}�}mQ:̮�g6?mΙL�n쪇"y�fo�o/��tO��Og�h�1Pѵt&�N�r������oշH���Ć5H���~��i��R����~Z��<���l�k�{�;�ϯ�fj��*T�������y�J��v�����w�D���ʝs�q|*ym��t�U��|/�Xw��]�N�ʡo�ϧUI���"�>3v�ʽ�E)��ɇp�usb�_��Fd�ֻLu����7�N��1{:5Ք��*�RV)�S}�Lz��޼�yyb�\��ZĔo7�~����nh���t6k\�og�����o8�ӳ��U.�Bkv*��ԫ�vŨȓ��c{��;�X|;{]��ˠ�綋����7�)�*����h������\��S�p�|�����ns®f�����T�'c6�$��8ue)��W���(�}��U�6:=�N�j����K�`_t�]oj��{�>�{d��7�ձ�2��loz��U�t��z=�w:]�%#ʱ��7۞a��n �P���&=�J�צ"����R��>�e�`�����4%
URV�K���p�x(k^s�o����\��<޿(7�j�mT�����ӧ��^lv���ә{�^{mҿcT�/e=�*������/���z�j�"���}��ܭ��'��9k���=%+�5G�����;f�~*Wo�C�]��S�n�L����X�j��~V�ޡU�ΕVs�=q���7��ڗ���h�����9��Rv�y�("����ѽp:��1�s�"c���1tޚ���S1�*h~�$fa�h�#-�'Y���K��k���&���n���� �r^��sS>��M��Ŋ���d;|�\�(���Z�������M���u�耫�[n�u(^�p>n:RDo3cK/.���ʽ{2��y�\х�y�
�jR���څ�+�I�S����8�_G8��2�2�B�:�7K�V�4��$�1������H}2Vbv5���Tf�S�p<t�}�J��qi+8��:Ky�KN;Q����][�(ͭ�� ��f�b�ێU�V�{�h)\�ۣ�E<[k����d"�q	i�]j�C��*����0LqD2п/�64��lB�G�pv��m�c�]��k��p��=\�f\L]�N�$��Tq��f*E��aNw�:�������B�����,ZN<�P,_v#X�-
3j��ƶ��}ե�YC��Er��N�{����u�N����3��Nq�ud��Z�Z�� ���[%�R�>z 	lɘ�د����:��<ұ�ACW[�b˖B#z֛4��v�,�Ek�UА���`r�b�����"�l��C󽮲`h%��\L�p�R�YtE��;�����u�V띷B�S7WEX2��4�.�qan��h�n��=���l��qw���|h7)"���[ɍ>���g^;���A���.�^�Gru��%�;���K�㗛mc�"cn�]+��Y�5��L��6�l�U�q��D����q��N#:�G2 ���b�mj�n�R}�-�B���cN�uò#�8�#+~�Wr�2���T��;�B�NG�ԜHV��/S��Sfwv�_q��v��$@Q*IGsf�ò�q����B�7��/�T�F�Vuuk��T��C��C/���6*�Opg&��t�5��m��f�c��9����ܮ&���F�u��bi:z�	��r��;P��p;MK�U�|��"��.���Qu2��zk~��'��*�=�<Z����������6�.�L���D��V�5��x.��ʗ�eH�.��R��NnnI,JŇ�;7��*��B��9@���鹙l�X�����]��/Llb�o� �_j�BDw���	���sO�;�ا�wo5��y��{���+��oBJXZS�z�tk#��-9NjӘ��17���)���k%pܮ�[�{5V�vsb��x��mV��+�%~���1�:��b#��U����Ew+�)[�h�R���\�0���-ͻ,��9>A]n�öp�K��VwS.d�� ]��B�Uʻu�]{�A$��Q����f��h^�F]�շ+q�0�SU�]*��mM1LZ���_s�-N�b����vn�7٭��k�o���:�i�B�_XG�<�B{\T
����X��3��<�ξ�-,y3%'Ԏ�][����ٸ���7�����I��~TX�"�b�lQk[e`���
�
T���J�(��"0QB�V��T����b��l�XT(�Z�@�*T�Y��h�H�T�V��A�-
B4�²���"����Qm�P�m���K�ڵ1eQ�[jU`�Qe�XĪ�m+D��T����b�+b�dP��R�XT�-�����"��EU�PZ�em���UH-E�U-hV#
�Ƞ���"��Q`T*��-[H�Aj�օ%KiUbZP�*VU`V�Um��cZ,iKcmTYR�l-l��UBĔeeҌ-���)V�6��%`TYKam+QIF�+YmPX[A����
�%�Tm�J��+
5��J�B�-VR�[J�V�VXT���R�J��KiX�����Z,RZ�AڒժJ��)RԤFEQ(����QKJ@�kb�KA�*-�E�9���#�"��0�k6pˆ_v:�VF�4ؙ���0nu�:��!y���'&��y"[�rW��7���aW%�y�����l�}�~��������	�8�B������SK&k��mg�U��/�	�2��o7�U57��q�;Ǘ�RglB=��O{�r_U��%����C5�\Gf.-��N�/��j�y3UWj�xק`8�ә�m{j�ޞ5o����9�֖��Qv9�=���`��uwꝽ3���3����f����s�_��p��f�����e��7���#c7��4�O�����~��os���������g�cqP���·$0���Q�g2��G���.�H�t�@��9^�1L�|DU���>c���fU����߽k�X���Q�zK����h��jp��k�N�~�'��+�J��L��Ϝx�Vw�gƪ�r�޸��f�[҆8ċ�t�t�%8���E�DF�z����<3���=��}~ȟJ򧱍��q�9��δ��+^��/`�j �H�!�<�x�Y߅�$��u
��
E��v�`I�廷P�L+tҀ0�-��]������ƴ���ˠ�M]c�U3����窍3�>�c&�����ɻ�<㙳�����͌��T���ғ�Ȣu�^~�g(7�1�(���7ݕ�:������s����;{9M}Qc�1�ϥeq��D��ұ�e��V�#輪��0����tG�{>��<���;|���~�l^#����Y7�k}���f�r�N�|���L�d�MێMܷ���H�#�r������u��$gِ�j�K��]gG�z�ɳ��h���ڭ���\y����>W��j��_*/�������t�c���ɱp��
E���_��a���ҕ�ܤ�L��M�����wg�������_g����oJ�\�׉�9�]ݔ��a`-�A	�T:�:��}c: 
�cg�y4un�i-���J��{��]yS"�S�5}/z�Ԯz�`M;Poz	�陷{��.�J����c�eF��佮�yKʋ�p��4p�E�н���Jtv����$�A���hغ���-ѲY޾���@uϲ����t�	K�N��S�f+:+"q��&��e��'X��Gpv��u�>��qN.�;+ħ}�x�7}��[o��´�!@)G��YH�1#��:oT���;�Uط�޿d3����?Q���z��N`�ڐ=�'�^(����9��~��O{��2;k�~˕q�b��/1��!�"t�@�;�9�˱X�[��q�p5=K�W���U�㛾<i,���Y4��	��ï'���T�}Lv#����^,o�Z�����B�ٽ��܈��P,g�2�h�
�|_���gnE�(��}�ٮ�o�\�+R���{�r`Y Hz�zآ���}����ܯRG�=����yw�[��yFk����sw�W^ӱhC�}�2���_j��%c�R+޽�S�N��ܺ��Ѫ�y�Y��+y`�پ��!� �����=}-}�G��+9��=q:c2zo?mżf/�_�7�i�����m tˠ���h���&u���Xu'�X�I�N�N�d+'Xl�py�$����~���`�?{ܖz$��W_+W�}���|��y�:�u��Ęa��iY>Aa�i!��ek$�L0�a�q���+?�u�̝~g��9ݍ˷|�F��mvV@�(���t����Ux�Z�ϖݑ�yx�����Gǝa��9�T��ug��K���1O��U.�h6҅TɳG�9��m�8ܼ��ڃ�`t��D����叆�nW'Z����q���i�v��Two��}�]u�Ԟި��~�"�ֻ���&Y4w�<��XO��+	��'��	&پ�Y�8�h����,3i!�O&�I�fMP�e����l�H���W�Gw�ק[��X�s�C�c�N2q�r���t��8���&��I���0�|w؄�i�^��&N����d�
��+'X}MUA_p��+�Vw���>3��;ly��I>a�x���q3Xu��Y�̝I��w8����=�z��@Ϭ�L�m�S���N3I;���y	�������ߙ~�;��p��ɺ�?|���*J���2q=��u�l��5�y3���̆w�N�y&�0�w8���;q<ɦ ~9�I��'_�W�U}������~��e~��S=�z��&P���fL%I3�$�8�ɐ�'Y6��.N�m>�C氜a�j��W�C;�'XJ�a����'�N=����}Z*��g��_ᓖ���ޯ��Ŀ}E�|�����Cl����d�a�wfL%I3�ԕ���C�d�'��Bu���0�a��>I_2i}�:>��(��^'��Lr��?y�/fd�K�h&XL'�o�:������m��AI�&g}�&�'�~�>̘2OrȲsV�I�N$����Bu����.��u���.��]ۙ�O�����X���g�M�|�ܿ2Jʇ�� �J��<���{�'Rm���)>d����L&5�}�0��=�s)?;`f߫�U]u�j�@�������oﾤ�m8βe��<v��2��\�	>C�o��$����̝J���b|��6ʇ�{6ɶMM���$����'���_m��Q�>a��3߈{!�fM���L9`z[�O'���4��L�S�e��<����he��.���O�uN�ɦI�?�2u*S�b|�̛�_o�U1��}�����)U��q���W��OT��yA�lA��k���Xܤ�f!�L�3]6��������;�R�c[u��[v�zt³m����� ޾f�$ث-3�Q�Ӎ,کm���ƫr�Wg���4��z��cl榎
%蛾�����*^.ѿ�������	���o$�)��Ȥ��I�u�|���$�3W�e��,����!�O ���	ĝB�ΦY��>�r����8}_5��}�W����s������&�>�I�b�6�o��y$�[��m�M$���(O�,�JβO�S(u�o;�y��,��q'Ry�;����������������_�ɷ���\���:�~a�O�:�a=�`�'�m�'�ױ'�8�o���|��hq��,?!�Ő��d�jb�d�Cɠ���LQ���#������ү��9�I:��T��!Y6ü�]��a��by'_�O��q�>v���'�O&��ٓ	<�ա�VM���<�Y ��5c��U;�����~��~�v�/H�����1�e6�>}1C̜J�����8��~;�HVN����<��M�'�q�	��@�O�2{��2N';�fL$�CAl���,g�q5}��Gy�������/`|�̟�ئM��k6L�O:1C��2
d�'�C}�$+'Xg����&Y5;�I��>I��'E!�߻��X��|��_�:�;P���f{<�y�(O��+'PXz�:�i<�`��I��5a��	�k6���!�c�N����!��{�oL�xϰO3̟�e�7���:�x����=����ۯa>d���dI�=��&P�,���Y2b�ԛI�j`��d�gVjI�dՆ�|��kx���|�ڊ����|���O~���c��G�=�s�2e'<wx'�N0�����i�G�� �N��~ĘJ�|��VN%d�(I�Nf����d�~a��
����|F������;�y{��n���[����ƘI�l>�4ì��=pe��6��XT0��7;�Hy�k���XO$�q�2a*I�w�+&��œ��_�~�GG������'1��6,�mB�Q�F�1V�����
Υ�N�)W��b�¨@L���H��o����-�����m�C��%��U���up��߼����m6��|��3���68V\{�s�QU��-Չ����il��n�n�n���� .5���9���w��t�e��$�i���d�+r�a�I�6a'R=�B��M��S��'�3�~��I䝿�&��w9H�q����x�������}��g����~�q�>d�N�OLП y�՚~I:����<ɤ4}�<�*V>���J���N��=�
�Y>J�g=�
O�g�������;q�~e�������_���N��I��LXq�ğ�����3O�̚I��,��O!�oa6�a���Y%L��2u+!�P��|��;�>�1ﱌ����?��[���׈)8��5��0�����_�L��dR~~`d�:�������0�	��0��I���C,�A�~�'�<�Gy��,'�}�{K�;�1���}����~��|~d�VC�`>a�M�I���8ɮ{�jI�MOo�nL��~I�}Y�I�T�0�	�|̤�
��O��'Pu�_�o��1�ow����ݺ�9��ИI�����������J�j�Y<ɷi>5�@�&�m��o$�@�7�ۄ�ɣ����d�Vu�|�2è)'(�����|[�߳�s�w�>����$�
8�6����	ĞCX��L'X~��2u����c�I�i>5�I�m����O���Ԭ�I��Ő�̲y9��|sދ޼�������{��,&�������3|�Y:����'y��Y�w��O!�wܲO0��`�'��Om�:���NC�Ğ`m&���ٓ:�\o[����Io��W1>{ښ��T�����~���N��L$�C��hu��d�V�q��:�C��$+'P��؞ݒy���Iǩ'�m�$��O��O���~r�߸����k~&'S�{Y�<�j��*N ��i!�N���	ĝMf������a�N%`g��q���~��$+'Xw��ē)/wX�׾���;�CU�<׶���,)�v�D_j�g�����P�x��vfQ�'�`6�]a�c���U���Xx�w4�Q����#f��޻�	�
�A��շ�]n5�%IA�8��ڲ�+�_iz�X�N7)c�k,<��2fr��@v�L����ɛ�ɝ'�UU�}�B��#<��+���I?�m�'��OoX�&�gw�Ʉ&yg��8��`q�y>0Y'u35C��	�h�2q����0@�N?!���߳�|g��k���q�08���qǉ&Rw6O'�4�O�a>fY99߳0�C^޳&P��B�q+&LP:�l�M,��<�5a�d�e�e�w��O�g��ﵟ��zd�ć����|����`|�S��2|ÈkؓɦN$��P�C,��d��k��2a	�_$��Jə�Xm��Vp�ӿ�������8�_����+�i��2M�$�$�̆f���Rm��4�̓���2��`~�O3I8����`'���S���XO$��~�0��k;��~����؟��u޿.k<`����(��I�Ơr����d�d�CO�'��I]�>��a+<���O�<�9��Y:����b��5�`'��>3Ͻ�~�D�?\���!�s�;����ݟd�ea7�"��Hb��I��l�L��4��u�'�2���Ԓ���,�0�M��4���u��7��g~ﻻ��ֱ�u�z2|�n�,?2x�?d�$�O��ٓ��߹�N?�3��8���~��?&MP��O�:���ɖO0���0�B�ϰ��&�d�LK���בj_��T}����>d�
C\�'�d�V� ��ɳ�~��&4{�fK��y��E'�l�08���~3CI:�i>L2y�R8u�"�=����ƿ}T��+�@~��pI�a���XO����ed8{�O�u�iX~�� �&�5�}�2L2k��$ۄ�)ĊM?0a?3����tr�.�~7�{��w�����!�A�|�AV$�'�P>C�<��?`��a�SɖI����$�+!�}���d۴�� ��h;��lǹ���L�����~���j��VW�Q�q���&��J5)��U�a�@�#�*L�ʯy����0K�6J���؞eյ�呜��x:���[Ìm���Tք>O:�9�`݅����)fLyW�x�1;���ݠT�j[�V�5�H���a�Ή�?Տo{?���ﾯc_����[��H~M2~O�(u$�*gVa�\��O �}���d�T���:�s���$������N��~��u�̜v��^Ğ`m&߱�����?W���{�����zls�	��a��Y�,�f�Y��Tά<��gt<���Xq'Y:�5;�Bu��h�py�$���2{�	���s��ۮ�~�����Ƽa�I:�ƽ�<��M���}�a'RaĬ�a�1d>fRu��.&��k6Aa8�VI�VO�I�N�M���9��Og>o�kc������O��O�=�`�O>a?�*�|���bN��f�{�d�$4[�d��C�m'Y���I�:�͇�,���,:�������^����ϳ�]�����Ͽ}�g��M�m��O��
��3��8��&��IǬ'��b��N2h��d�I6�޳&q�է���Aa�ZC�m�ɠ�d�a�c����;�5�}�}�]>���ǃ)�I��Xy�����c�N�y�r���t��8���&�}�i6���N��u2����$�	�4{z̘ABd9N�Y8�×}�>��Ӧt߹���^��^�R~d�{�|ì�k$�e��;��p�0d�O�0��ql!���q�O�q>�y2ɶNO~�'����,��kz�f?~�(~�թ�~�El������P+����eI��m�����ff�y�������̆�gP<��9���Nh���&�|���ĝM2q��돼����{8ι���w�N!ğcX�u�ٓ	RL��%I�VL�̛d�Fl'P6����'e$��C{�'XJ�a�w�?$�I���ts�}������\�u����&Xq��!P�&�Y���'��&���&�'�~;��&��7z��s���Ru�l�r�4'XL��i���~��J��H~�ק�7��7R�W�fɦ�W=�|bn�w���za�ͻq�ft��l�b��!�ơ�"zvHXM�=֭S��ME��TOΡ
7p��k��huj�L�����G��nG��"�E+���ȷW��C�����Z�����]�Q�ҵ�� �]}��oO�}�g?�̒�a�5�I�	����'PX{�u�h,��AI�&{��4�<���}�0�d��d����'~~O�hN�<��@hƧ{3�[��̪Ⴞ���_~�~�,�C[�<�+*��<��*d�py��,{��:�l�~�AI�&g���L&59�&�'�ĊO����)�i��?w����b��W�p��+!�!�4��d�$�r��2��G7�O���0y�T�~��N�Bh=�O�u&�P�s؁�M�o߱ēVo�R���B-y�J�����^����~�$R~x�Ͱ�	��6�Ry	���2y��~d�2u韰I����by4�>gwO2u*����'�7�L�z��`�c��g{��=u�2m����z�m��s��8��k��I��&�F,�$�+3�I�&ux�Y:�ɯ�O��'�]g��N��s��I��}Ͽn�\����w��g�����&^��9�d�'7I�X2|��g���m����&�$�O�P�&<�ŝd�2�MP�$���<��M�8��<ʛ�5�=��ƿw�7����8�L$���cx>M0�a����N�0���Y<�o>��$�m�`���q��4�YɖN��L2M���hu�}wxa��ﳭ~���{����o��C,�J���M��N2��}�
��=�x�y����:��~m����'}d�	��$�N�=-��m��hŁ�2���u�ӎ�����η�g��I���6L�O�LP�'�2�8��������!Y:�=����L�׻��z�~��I��O��ن'G}�Ʉ�Hr���k��9ۭ�ϵ������P��Aa�`~C�N���	��M6L�N:1C��2C��d������3���ē,��<�o~I��}�N���׮>}�_���>������]�ǈ�9꬙����b�A����ue���C��Ŋ�thz*^��7��\�L�A*cU�a���e�OX�~��h	�7F���~:�1t/t]���*c�5#ʮ����\;�^���ֆ��>�t(V�z߳�[��^�1hf�Q����aͩ?#�}��gl3q�����2N3�絒a	�Y�+'XfZ�m'����q'S3VL��f�P�'�̆��Y:��|w8!�0׽�=I2������n汏��=���9���<O��M���T���OOw��<��o�(L�ΡY8��&(I��f���L�ÍI:̚��O����ez���u󾺧��3���������������8�sM?2e'��	�i��2����d��dI�4�ٓ	XL���VN%dɊRm����a:ɴ����a:�z����O��g���}�߽�zI]�?sXI��>���<�;�d�O�7;�B��M��]�$<��4{?�	��?fL%I6��dۤ
��O�=�9Ǵq�}���������������,�g���ԓ�h�aԕ�M0��c���a�sXy�w�뉔�AHk��*d�5�`�����2�y'�q�d�V�3��W��^v����~����v��&^�{M2|������ff���I�5?X��M!��̒�a���$�{�O$�
CP��
�Y6��=H)?$������~���s���w���g{����'�߳&�M��dRm���`q'����:�c4�<ɤ�a����'�����&Ь5�`�$"������Q`��i��\̝��k��~]K,m{���Eg�|O�r՞�um�$��篲�I��0�u�i�˕��To�k���w�ڞPo�c6Q[|�=�C�L'}�Z�7��76{b����-�UG����aO9�o�����1g�h�	�ș�������ߪԂՈ1n�rcas�XG��狜t�6�Kw)������qu�tGN��N<�ٓ�qY
�j�d2sn�CM] f���t��3�����/��2H����&���%n;����FB6�xǇr>�!�u�s�^-`�
��1�8J���q�0Q�+�:9�kk���mc���%)R�k���_tU�]�$��u�֐i�ʺGnt��J�v�ܧ/r�Ϟ�2v�A�I���܍��ѵ�w1��!�iC��L��V��]�DIGu�Ρe�4�mWJ��V�;�Wua�'�k-�i)dR&�=��6��w:��<�ҐT��n�e����,A	���=��d7	\�95vR���q�)%y1b�ep�	���[�q�n]�ͽ͒7qc.���[�i⡂$Ǖ9��˺äcW�{AҌ871Z�m�+@�;��j�O��T��,�UڂY�
X�*dG�m�WeӽjЬ�|i������<�$)��݋���b,X@�6��=���!3�+ϱEV��F��nν���77(@��m�T魹7Am%/f�疫�n�����{C���(�ґ�J�O)��Ԯ���t�ڮ����6�y��,X&�5��+p�#;q���<��9 JV���� �g���Y��Gch�+g%l�l�f�%jz�(l��Z,�a]^w�;�Z/��A§Y�����g�)9m�����<�RȾ����6���'۸!�L����q�DfGu��)9XB�S��I3���(5�W�`2Xk��
��"M��J����9d�7
?kI���7"GNeA.tK)#�Ġ���a&���Erj�5��)��|o*V���	�޹ՑPM�/�}ܹ�y�5�1*-���큶8g�P���;9@�u"%�)ݨ1>�ʮ�d �s���+���ù��p�SX��0AK�5��n�v̬����v]J�̓���a�}.�{E�r�����0l"T�����s]��ٴ��N��l-AW�e7�Ye�io#�y�O�b(s�0��Y�l#O(�Y��/�Q�JC$��/1&
�{]�W0_[���36R�&�����_���XBhq��Vi;R�O;���U�'=��F�&,`�5Z|���V�V^�_픵t�8 �fPI�%�n����kr��di"y�w���Zw�5	�o�1�a����� �+KT;�E��(�ܻ�f����[��r	�� �W9m��`��*���'Q�tw����r��⺰7����|�)�{�c��v<�I��"�)9өYz�j4l�ft��r�P����6�ۗCt>,�z�
*�T���1CI� ��yv\l�O&��=Y؆�;���Sf��
9�tW��Iۜ��$�T�F�;��o5�E�w�3�~�]�BX��́^v� L�g�f�I��W�����܉*�xږ�#]v��&Nҙ�Y���0���R����q���>�յ�I<�1tWo��T���;�� 'u�Lx��]f����Ú��~ �)1-�P�[J��c-
�V-j���TX��%�VR�%TUXQ���YU����m�#AJ�PQ�T�jʬ��@XU`�**QV���*��@*���-��¤��YieaKdm��jT*J�Q%@��eU�J��$ ,X�V
�RH[aZԅT� �"�,J�ETDIZ�H�Vm"�VѴ��eB�EY+�H�U��Q-�Z�((���(��
ʪ��aDFTZ��[j�#$�QX��V(*�"�eem���PD������5(*,U����b�(�-�Dm��Ap��Ȩ��*5�`ʑe�����-���U"��1cؼp4g5}��1��=Lh})sN���K�Ź�W��zJ��Vԩ)�mq�T�3Wp����ok�co�UU}��U<���^�غ�W)՞�kg�y���N9��'n[��g�0,ҒĻܷ}��s2�ꓣ{�,���\�L���~���S��r���~k�����j��ew�O��G�z��2�9̿^������/rp�����͞<�F!ê��~���/�>��o���ym�v�G��!�3Z�Ow��UMë���W���5����e<�3{�Jt5{W�po�w[Kw}>��Os��Rbɚ�?�j5s,��k����bc�ˆu���nM�c'��1��N�ʛ���)^TȕK�k�<j��;p�\*p��,j�sQ�� �}�8}�6M�S��*��9VE=
�f�~��%����'Og��s"V�b��e����71��d����K�=�}_��Yr��.�g����pB��*k7'�.�<�� �}�3C}#�N�
�M�z�6���9q��E���ލ�S�6�G��ѿ�ֈ��h�y��n��<n:�W�>��g%{
o(Q���-� �~b�����QcVn��-<�Q���%l�Qe���q`�a�o4�*8��h���k��f?>�UW�U_W���I�(��˯�w�Щ��Ә�T�����o/�Jc�������9�u,�����u��)1��Y��UT~��6�N�e����ܞ%w3��S:}����T��zVm=�/���e|���g�o4�oҊs�|�)pD�v���ӳ}~n��.��z��y�>OϢ�=�)�7}I�=�ʴEz������6Wl�xnn�Tg��/���g�
���Q�>���{�߭���&�.��79���:ϳ�o�4�a��3��tj�J�lu=p9В�K�h�<=yG~�+;�S���z3Y�m�
��	gS�o�w�����0�^w�������ޓD�����*8s�Ͱ�m�$")̭8v;�]�d�P�e�vo�=ޛ�fmҾ����fu��ꭾ���8L����f����d~_ؾ���tS��U����S�\�5�<��Ogfd��R���i�<MC� 唺�#�G
Q�3���=Y��q���/��nGY^o%K�I���*�����FuPy]����8���soK�{�% �skT�y.�HV�����E�,,u��vv�b�[]oDX��z2�nI�q
ɡ��PH���!�����1�k�pz?}����3��ٞ��~�S���9���]y3����kX���.��q{j�����o#OmA���7�"�`���ﺃ5n�y�{�s|�C��ڭ.��Y8hG�S]���Π�)|j��^�_���Ǿ>��{���'&���c>"��;���V/7�iPQV^H��{���������t�}"t�iWJ�Ә�3㓫��}���xR�]��p�ݧ^v�D�7�juZ���:�?��z���Ut���I�g�=�{�栟|r��z�w+}�����������&?黝R ��r�&���D�T��־�Y�5��׌��J��|�/eS��rul�Y6�d�t[�zMk}��7��l-o�c7�G�|�}�탩�PS��R���4�ђ�?R�����'���F��7��۹�xx͢�����}��nN�:S@��_�䌝�s7�vsOW/1#���59��z�(�9^�]�N7�d�=^V�s�ި*���� �ïnDEa��Cvs]�*^�z]tںT��/F�5n=�t�5t�A:��x�ɜKb��ŝ��h��hf��MsA�I]������ه���I��W���ʋ�g���ުRv����T�^*9m��6b��'��r55>��O�M'@�&�s��T���H".����סt�KSf��Os>̄��w|3��z��j������=���=�g�����'��o>�:�݊�毯����c���֩����1@��9�U9�z�����S�j������.�6.溧{2�mU�N����6ގ�ޓ"�4���>�O��*w�u�	4��ܔ��u�˳�� �Ͻx��[��Kwf����b�WF���J^S_9�/��e�Z����p�}�a��n���]�+�w5��Tn�������UKʊ��.��Τ>�m����w���!���N8�e�t�]��Cn�ծW��1J�^ӈ�b�wg{=�s#��J3s�W�^k�ȗ� �s��{Ew�.r7��K���#"g�A�r:w�8�+�qZ꛱�Xhv��2F�h����p��4��-Yk+��q9}M�n�ޮM;Ǯ�%����hi7�R}��z�8�#˜[Y��j'j:μ�ze��١Es=ݷ�����p��R�bjO�'����꯫�mk~�x��������Oo���/�>�6�f�[҄�>�gd[��1�r�����������+Y+R��|3�j�q��:���]ǽG�v�^1ҏ����zM����3e�����#r+="�I~��+gy8$�>w:����w��˼�rK��2Ǌy-��w�.��\���q�"Uc���Ծ�H���A�G�ޏ=�rY�9�Ōe���4օ�����p_����̈́��.t�fy�;��Q�]^���eI<4d�%��z�nC��Q;�+���gG��;y6S����C˽<�[�J�'��P�D'{�ê�kD�UW/���L[{�$Oː���qV6�޹|����j;�Q���ö#\�BM�wÉ�e��-էy��x�w�l��n�JLԪ��ɶk�s,��yp^��nVh��M)[��˞�����L2�k�Ǯ]�x��J�&%
])�V9���`�Q�ϲ_@��U��[�����l���3\��^�9�i��⺾���/;�U�R�_S�r���r��t36d�2��,���@k��u��o��99s��������9�痿[��m<]o$?Ϫ�v5�wO�d���2%R�sƠώ<��^f�=�il>J=��[۬�.�^��w��g�Ⱥ��)��$I��YS����E�4���e���b�,�o�b*��;>f����g��e��J�Z����^���!ݭ���h��n��
�D�`·��п��VY)ˊ�=K;�|xٞ�ml��t_7��͂RT�j^r�uƻ�z����t*��B��K�1�ʞ���/�ܭx��_�SfM܋�{ܻa}3zp��Ig�3�T�ms�^�.v~��{O��i�j�su���'&��v���h�cr��Z��Y���?U>���3@u�f=��.�j��� ۓ6��pٚ��<[e�]�Tz(z��|�i������*��g�w���gb;��tK՜�Zo<}q�ӣW�R��§�gVg=������ӥa � � �j]F��t�Z�C�g�c��7���G�A�B�%���֦�w(�g�}V6W����b�OVW-�.�b�-g��Nv�䅨�x&9wgH��/��{qN�����.�rg����BVԳ����_}Y�= ��^ٺ����j��qo��^�8w�[D�V듁���If�^�ǻ�����xLc�9щ��4OnNmQ�b6��5����שa����㧷�[y|�_����^�c�ޛ���;<���)G�
�1Վ�q�s��sU�J�Z�;����ls��\�~^��������g�ً���{3ɴ�Ԫ�%X{�t�5�=\[�z��Rs�{�R.�vx��~wOK�:���^<��_y�S�Z��V��]����ݎY�Q�ӏ�s�gzc�}>{˫��Ss�437�U������9��qg������J���L�ܩ�9=��F0�V�؋�k�|�WE%;ow1�W�{���:�?V�ҽt�(�6��3��ъi�=n����'�������f����z���Oåc��h���݋��#���R��0�z|��V��b�X�����g��2�5m���4h������b��O�z��]{=���R��xm
֥k/e���u�г���(8�V�yW���mY��Sq0�6)�WGt�][�X���.�1��������{�S�8o~�z�^��W�w����[҅��aI硭�̫�x��\��V�\y���ˆ�j�mJ>���-N׮L�ۥ����x�w�{2eA�d�~�Atj�_��\��x��U���~
?.�Y�+�\l�~�.XQ�|�-�|�\�f����^��X�B�h�y�V}���'��L��rW{tG�*.)�q���ޥ'iy����6-1E*-���.{���y{�9��O�\s�3�h~�rA�!~ ��Y��ڛ9;��-�ǥ"�|�/�����w�ɶ��������~�V�a��	�ڼS��p���L���6�����W�\\ɡL���|*{b���f����f��1�a�Tk�����_q��٥�y�w�O�g7���{����T���A���!�C���gx�j��o<j�h�#��o9h	'w���d�í��gp?-�s���k��6�(�њ�X��w�c�m�x����E�|hWi��$��N��8��U���AD�k�ʳۇ���;��]*)>}��hL՗f���0�Z� ��rj�=�P_pti%�ms�j�.�U�U}G���\�/v	?RU��L����[R��yMS�"��^����W��H�6��ng����[ֱ��*w��75�}Z��R���"�&���|߬CV}��\��r�k��Ջ�}�jWzL��'����pP�	7�4I]+��8���)���k�P�=K'��W*�ȗ����s�m�CGS�#�V�7���(�B��{�ܥ7���u_x��Ƿ�AKM[<2���XB{1�s&��ȵ-�O������IΈ
��L�������B�:'�߭9�Ncu�}73x՗��7��g��{u�1�B�έK�vei��3�(�e癯	���fu���/1]3#ھ���~]���:^:*Q��Bz%X�Y*��q�`�ʆX�a�C���0�{9�yM�΄�Xe���<��#=z  ��g���ߋ���͛�v��G;S7=�^�k��J��
����ܹB�u�Hʪ�	ɪ
r��ܛt�׳��LO/z-ޔ�ݻ������]Ic������v�9��/Ko�=���B9��ܣ�xb?-y��S�r�4R�n)k0�)X�Nq�]�ދ�Ɇ�H#Egᝓ� ���&h�������n�AH�Ĥj�L�T�f*�͜�О�u��������������o=�p��u֗��YX�@�i���s��*��gJG�x�}]��&��ۦ����ߏ�{��w�U��K@��<O
h�\�Q*����y� zd��}[�<Ѿ��aOs�.�.�ҧ{,p��P�,��F�po���sFgu�^R??vzt��[������-���q�{�C�e�X��en���N�t�Y77S4Nw`����/u�Q�@�ZX�������{M_�枬�0Ո�Gb�*o��4�9��>E��W��~h=p�xUq��;S�Y��Odw�����(;��#�!�w�_�^Þw��M�{!�1���B��S�W������HU��`�>�~��ܙ�P힅#�N��zz�K��`�4p�I
��v��O,���)�<p_���ՑK�Gg-�ׯ�O�:��X��Y���ϙAА�w�Q�P�)ݜ53�w�}g�'�GZ� ��߼ywMԻ^�8=�BS:�*݊���ޔ���(`�Xӕ� ѳ9Xߡ��GUUD(����-��.��\E�pԮ�� �U�;:��2�l����7Q���g!����Y�r�x��;����[w�E��n�q����f�06��b8@��]��,1���o�o�z�]�3]zU{tb*L@}���q�����D�L%��|��]� ��I2���a��JgioC|�W=�eru5`����ʓ)�33���T}�vp;3�(�I�u�s,�v��i�u���oQv��X�*齫/dofmEz.wk��B��Gyi`i� .�t�ږ:�B�Qb�-k8�㞴�]�/z������E[wX^啕��ˮ���4��@�[���.֋�U���˥��;�<���w���dt;q�]&�K�v�0�V��ر���I����8��Ї�V�{�V���v�����M��lc8���èm�`��ݴ�n���΄�v0��D7/I�τ��f,
o3�t��U����A
B�ޚI5������hf�y��'�-��ms}Q�{c:践�Qq�ڐ���x�؊�rb�t�eW��tU�t�n�*�J^o!AD8�J���Ҷ2��-Z%�_q��,-Hr\ڊ�����8c�o�Θ���wY��;���a�q��m	���<�B/΄�ބ���o��|�#F��\ֱ%b,z��e����8���]A|�W����O~��s���X$8K�3dw�6��Kr]�&On@�����an�����)sp��⧸Zu8�T���z�TjL�Qm�r�[ݢ���j&#��׃�0�����q툰3	��r���D>��9�03��De���z��5�K�����h�#��rb͹�|��ˍ�ڗ]��cQ�Z�p��Et���1X�́�ȫ��ٽ���Y�p�NU��'���Kɼ7Wvɫ��ލ����KOH�.%upb�W(�薦lC�շ��\5o�v�[۞���{��-�n��W0�N����R��Ҷ��J�]N��T�2�$(�a\�7�n�"�u��Xʲe:ʔ��mf�v3{8-J�Ǚ U��7�r�4v�]>#��ksqȮ�����;ʼ� �U��+:�0�����eB)�L������w�σ���^opf��pi*��G�f�p�Up�w����DTѥ��e�\1�J��$��d��7�Q�ΧAAű�_HB\����H����+4{�hmm�c�9��gb�n�����{��9<�9Q~��ړ�������SK}W2��Ď���,Y�ð��w[ʰ]l+V\�m��<���*YˣDh�.�R=ř{N���V�*���"�Im���p��0��Mk�T��KI"�5�F�r������ፚf�	g%c����k"��q*"Z�Jfc�:�Ac���:��a)w}:��pW-���wݬ[�=M7{O��A>*���-hr�ū��$�@:��-��՝�2E�����Zw�v��9��A �H��U_��\7 �ԩjثR��m��T�h�BV�X��Q-Z�B���.1�0F1,Fa�m�E`�*�q�a��1H�DQ��cŔQm�Upʊ
����T��f1����"*�Qc"*�DUEA��F�Ukh�Vb�F�QqB���TTDQ�)�5Y
���j,QQUUX�QQ��ԍ�h�Km�����H���E[J�l�A[QDE1J����
��[aTk*��$�Z� �cE�.Y-�ja�E
��S����#��DUH�b�F�f)`�
�1ZرUQh�T���lL&+DURV)X�[A�%kmI�U�UQEU��X8�"��1j���Y'&�St&��/F����g�M��;��K<�s��{�X��r-�'v�iT��ծG�*ͽ=.����u�� -�N��=s��[��+�MԸOm�2�|��R��J��&L��:L�v�����^��Qc���_��;���*��8�MWf�dg�D�e-^*4�{>z�����ǧ]�^��O�z�{$Nq�g�ќ|%Wv���x𤾣x�RYփ���p�Z��Unfm�U������w��,�=C���{�,
챇�u�^�a��(-b*�<��=���Tӡ��l��k�J�*���c��*�ʛ���Ƞ}�7� �,^��yK�BoC����=�����j#�od���:rn9�2���p�����ؔz����}��y��{�(�E�>��կne���,}�!���~��J�e{B������"�;�U���d���.[��q���\}����.���چ�I�yK�]��@������A��tZ~��S=����?�{�%��þ�0�������"��ژ)��eK�|8���>�e�^��)>�v]w��;;( C�qq*n(�����Oo�:����N:꼢Vt;�4�4v�zR#1�ݙQ,�W>ïK|���}z0D[U��8����	WX�I�dZHX��(8mCk�0)��R�W
�3ab�w�Ri[ޠ��ٙ�9���ڗ�D��r�\B��'�;���� �k��'��8��wﾯ����w�,��]��.~�1��'��>7ê�N��HbsP��5إݮ�S���\Y�i�=��]� c�fp!T��k��O���ZP�س0A�zQ�WaUVXدV$�p�i盷���0\ܙO=zz�7^Q%}�wRf:U%�z��@h_C������`������1V���=�_C`S�{����	�F�d��r�R*t$)��,1�l_����s��Ȧ_�ak���g��r�p4�z��|D��ǝf� U=PZ6l�;}o�y���;_N��d����}�9�>��6�PLo��\4[>�W��s�h:ū���M����\O���ٸ�\��h�K)!�;~�}b�W�Z>�Y���z��Q�lD�>	����I�A^�}�p�M�
�W���f����������Ѵ��K����K��eǝ����bCˢ���nfA�����������}�B�9�6�h�}ƹw�!�1_hŀ=��`�=��N�bz}S��Ȭ܇f�,U����#�{Մ�#��}|�6mK�V�9�E�8~��.+��[�lcPʁ{�߯�ٞ��*�1���Ǒ*� �S����ݍ�ц��\Q�Η�@��9*�Aާ����T{7( �1���C����L�5���v^WR�c-m���}�O�}��_U�nW���q�A� "��ߍ���D�ʫ�������!���z�5�_���Ƿ�O�0l�q���y���٦%	���3�7��+h��W-���f=D?^��)2	TNխ~o�{����[�[�M͓�=��;.�MJ�W�@Z[��Bnz�->q���޹׾������w[KsGv���{�	�O�����]�x��DК�%�4�!��\�
���;z�n=�b�%tON}.(5�}��ʮ�����A�*/R�+�����HU���h���S�˱�g�G��p��2�hw�*j���ֈ7���U��F9e�.���Ԡ��}[Ք7dޗ��7]������t�(|��j�������%��
N�IdV�[�/��M�Ʈ�?K} }g.R�&���|'Q�.�������e��(A�n��;[� -��T�_7�>��&����< �݁�Nye^tܽ5<�����n�﮵����C��y4�^�0���<u����A�g-�G��GC��9�W������7B�Fo:o݁׹ gni=��cK�v�v�[׮��=Ŋ����0�&:ޫ�r���M=dE�{�����4	Rܳ)��������:}���+ep-m {%��rw's2�='�l����Wʯ�Wo5v�u.���/��м�, ����gt�+yt9x���{k5�������7TܙЛ�����VR�Bġ�i�L���L���	�hv^y���qhٮ��K�w�,���Vj]C�E:9u���^�%}S�A�w�|�w�ӣ���	.H��������	r��v��^�������W����~����P���EU$�4�k1��3=��~��K�|�&+�(]#�L�ąŲ{��窜��N�)�nS��k�dht)^��^r�0j�WZ��K8Q�/+��%���lĥ��l����WDt)��Wm�7�U�]t�	E��'=��=VUK@��<O
h�\��D��t�9�T�ǁ��@��������kx�J���)��r�!P,p�e�7i#���w!�mVW�O�Y�_[O�*��2���0)�x�L�+UL��9U�J�'b��}v�^v^giy�.z��T�ᚐ0��X�3��\3�l�`�/4�Z5bL�������z���&z-y��R�*�7.���!����k>J��_ᡉ���(pi�=��G�7�4�����ՉeqRFk�(�Z���(5ޮ������`�;����i*��U��ۖ�a�1'���9�a�1��\z/�ZfIu��x���"��i�浳��ޓi<{и��R�%�����93��[b�8*��x�=�~����'QO���훵h��q`�\�:��5���h��ʽy��
s�+�@����T���S!ixX��L��ž#(���v*N��S:��W�_WlA�� �d��V�3s/ �[��t��b-zb��|����!��
���[�s�y���xFe��5�^:?>��X��=ٷ�<�5+^���ڦ�i�iέ���2P��;� ж{��+���������<����,���|��,Ԡ��oQ�3�ע��]f���ɷ��>�th�#��/�3ƌ�W)��^_�����UK(�X�5�>��-`����{�2����Pzo��ůw�~j��Ӽ�Z'F��w���Z}��x�-B*��-:��:�t2���8�1�Gp�7����/�U[�8l�؇��]#�s�%�e�>�*�+�����<o�1�(z	'�s��+cİ�Kjq��u���zyK���)��|X�7*�Q�b=���>j�;��u�RB��p,i7�/QS�lqw�^��z};�#=lL^Vu��B\���5����α�����U�LN�>Wi��+-̺5��1ݾ����8Z�j�n�����8�:-V�VjJ[��!n�ָ���f��;�gTԙ���V�I���WyCh�`wwrǖli� �>�YA#�ċE�=d���;�!������}�3�+��s�a�I+3�6GPoaT��Ϟ�eS��C��ϧ�*j7[3��������;��y~0�!Ҡxt&�q�U�vU�ӛ{P�����R����f��{/���T��O��V�^�GP���4"�'T;�����='��.�s�;�sz<�d#L���OJ�(p��ٜ��<8'��U5QN*%5���zey�\}�%��T�G+�wcI?�f���L�ã�#+�Ǌ��4O*륞UY�ybT��<�u�o�E���w����=�c�'K,��ED/�^C\����H-��Pj��0A�w��1]�r>w}YP���7s;���8s��=��~�E��K�ߍ 6��(ȓ��Ie��q�f	윌�{���./q�*{g<"{��׮hJ� �����~��`��:�].����KMi�A�g���_R�NY�ϴ�0�?9��+>g��[���y���U=[�(�W׷~�f�u�󰻲@j���^��6����{+�ҙ_
��{m^�\��,`���m�OZ�ٴ�1��]�*z����q�t���"on��L�S�����K���҇}�Uר��q�c�c�I��qQ��9]�e��������ǅRYKU����a��L�;E�B�T[�5�����re��Z&��}�UU}<�\}�>�ۂZ�#j���f���aW�%��O>U-W�p5�e��~��N]1Rtg�k^��z��]�1oP��=Iyp�|�3ӟMj
�|�Ѻ}:l��Pi��1��ty]f	E!A�2o[����L󫫥.����Ô���[��q��]P����ۖ���N����w��[��]�L�`���u��<م}�S���N��{�p�����Љ������i�tx�'I�3���J�V����藸���U�y�}�����i��T]q�������D�:����C|���IrP	L]���Қ�xJ^]f.*��V�_
Xu��ב�*�2vpC>y9�G���EN����ˡH1]B�%�uu�b�Xh�����W����[�nqw_m�ƽ��|��b�O輪�w�
���\�>c{=d�iT��~;�}�=Ѫt���*ƷNW[Pkکk�<��x�t���}��͚�j����݈XU�q?�'�]��W5�nO��\��&�]uQqۭo��5���B�h�,�������~��7M	�
>�)�2�D��wx��#tm�Zc�|�A��ˆx�.��$�W�:��t�㕷�^;��ez�l��/p�n�ӥ��7�yG�LŨ+��(�P�3�����ʾΪ!��M�f|o�B�N�д�웊
��hpWb�������}���|��^��8}��u�x� ߻�. 8K���C��m�h��C�Rt2|)f����v_{�=�wp]*��e���_��>���K�E��|)}L�< ����~�ԁ{mZ��۷��<��`Ě�^�g"}��A�];C�Y�Ϟ��(*�[t��+h	�;�u�<寏J�^�o)@�����D_�l�;�[������9K����|�}8�3Qī�Ux�2��Y�̡ઞ�ԼfV�0>0�Bs���4��מ�V���"ٹ��xOL�l,ԥ��N��W2z%Y�%O5q�|�t���O���Y������pw�*�G��A܈��!�� ǃ߯��~f)�/e-i�=\b!�v���!h���p�'��*�1W�Y�a����u.�	�r�5AF���ӈ���k������WZ/
Ͷ7
��܇�
۷�P�#[M1��jԩ5��y�.�t���7��o��!��U� �&�}��v�3��E5��h%�H��}7k`����K{��]�R��zEf�hY+p-8
�A����b��L^����Xv���9
��[:WNe�|�gZ����`�6�Q�Ȍn 3s�s[��ҫ_ڶ���u]eV�������5���m+o�@���i��V��9����o������\���e��o�&J��&��v��b�[�>����3�g�@o5�ߦ�*� ��r<��\�����v�ֆ�jZ���ŀw�<C*e�X�fV�ϫ��gq�=ٛ�t��&��t&�0�Uv�C�]��cH��|w#�6�9�s�����ˏZ��k�d�]*"���Ǟ���v�4�GR��8v��0`������V���z֟�hɳr8�1x�uFpĥ��>"��P�>m!�V%�W���+�~ŧ��8�����r��~�{D�͍%�=�)�L��|FR��(sdq�H����ز�Ui���"<�"��չ����4`���<�Uzd��}P��H�;U���(A�N��Ap�t�Hly��Ӧy�;6Y��C��z�[�i9[ΕU�2Pτ���v��(r�CR��L�O	>�Iw3¬9�0��ߪ�\5('��C)�襽)W���NUM����{2�X�ڔ��_{!��z����}&Tj�jֻ=����L��^���cHW��k���T�퀑��ZJ-��Ezn���DZ(�t�r��L�����U�gv�=��M�e��c�s��-���gM����ƍmǴ/b|�۫�[n�->2�����d�i��3M�w\3z�l�F��,�,2:�x���S2��w}s.gQ�{���ﾯ�|\�=�F��د�w����H��٪�{0m��	t�Ŋ�+��A��m�N�8����&c�;����^ȷ&Z�FM��\�w�o�x=ό�+��u�^�me!@-b*�����K<�R���O�yv�i��q�\����^�"��=N�������ˮ�g��Z^��yK����Ǖ�A��7�dVg�NѺ��Ք�\W�N=��:��qs3��=ӱ��p~�Z/&Iv�.'K���%��r��	d��_�
p����?>�2���{"\���;��Z6l�њ�W�WJٙp�C��,t9UtX�A��u<�Z��Ϲz�\�2IB��W�-�)5w��g����2�p���E5��ˡ@E�@k�Ai��R��Y�^�Ke�9���º���]�/j&��r+0z����<��j*��Ы�/�!��c�e�`ǭ[��Dgf7��������k��où��tz�eqO�*�N��D��Nj@5إv�cQ{r�zS�*H��-��;:{�����S5[�����q�uTx�T� 1��<����^K8�f�"_.�م�����B��k�הo�:uoa<��,b�q���X|S.�]$�ѥa�Xo��PW3�T�b�*��k0���=DN���	:n�����l����p�,�x���\ �/ega�v������Gn4�"y}�Ǘf�0R�'�v��=�,��Qt�n)`�ĳ�ڲ���ݼ�b�\5��;S:��θ)����雜�su��C�N�|�� OE��.S���U��}5l�{�G� ��4d��ۤ�09f��ڙ7�60�],�yvy-S��>�nm��n�j��<L���5JT�z����wj*4o2�f�`Z�M[�v'�U�Sx�ȫe��l-v�XїJ��[���Z���i�L�0�c�R�p��\���\U���0��4\遭̰;�W%�'w��*�AE�b3@�,;oOgr���# ���k�����z��xz��65=����p�ͮ�����1���b���j��1���j�2�p��x3�3�yn��M��o��q��ú�_(�*����o)�ӳs0U�t�9�s�����!���v��OM^���R��:5mt�����'����ja���$ڳ�*�V�]��L��r�]��<���i���[B����i�|�Si۾�M�O���7�vT<S�p�罻a
r�VN��J��X����/���WVWX��Re����{Y��\�,Ň��^�H�9z�����X�t��X�P����1��:#)'��w����Xp_)��&��Z��ǫ��c�4�^�ihj2m�(�q�X���-�E>b��yu�p�}�f��
��>����nӻņe���m�a�nZ1���RV<����9�z�x�`��qiNK�%x�l�Kw�A�F���p�&��X������v;����r��)��-v^Eolo<7���ϯ2�ZC�u����RǏe�9�rt��j��'B���ޙ�Y��VS�mS�b�wL^��􉤕ݸy�<̑u�ͳ��+��"�B�m�(Z�����/�"�S-�Qm�_��ZL�.2�S���{6e��@jm��9޻ɚ�3��i��+�is�B�Pٴv���Y����cN���Y����hnQ�EQ�)j!�ĸ-��V�
��\��s����ś�zE��eb윩�����R�_#+�e�fn��7���Gf��H��W+���_iy��-W-8�lh���Y��,;]�D�fBm]η�`	eսk�N�����v�;��5��Z�s�%��� mW&�z�E�71�#v�G�1|�!y�})���3���s���c�e��,�M�R�ۭ�ٽ9�0+�S�U+�d�ԟS`@�2�����W�������+����P:5շ���ӄT���bu�s^x;bC�
~���;����r�ͼ\�5�6���5����c#J8Y 2	�~?̣�`X�Ɇ"���1l�X+J[U��
1���Y�)�X��0�0b
-R�GQb��mm����b�"ZUbF�*��a
#ha(�1jŢQ0�,[lZR�	�k(��#R6�+m��Dŭ�Z��1�B�e� T����`�U�ł�qI�U1h"�q���1q�bEEGL2����ŐX�Q��0\2�+UPm+V�0�Y���
�b���Lb��1!Q+QjT*T\&"�ˆ��b�ԕ�U�m,U�k���b��Ū��Z0Ŕ"+��QGpa`�EDL4�1��-ZV[*"���EF"�DF�ʕ��iU��.0P���Ke����D�*ʭ[eŸ\����-���*+Q�
�b��
#-)P�,cYpՈ���J���G��p�X�FV�Dˌ����W�3Ue��Clk�<-�g�3����6�b!�ݝd`���N�A�0�<�	�w$�{��Ԡ�QP��������X���<��$!�Wa��W�r�}��/7b�O}M�W�f:U%�z���\fF0񘇧{6x���r��\B_�-�r�P!�a��:�%��Xφ�'q�TUH�Е3̞��
}��N���z;��{��5�',��XC�]���Y���x]n'�z+5~���B˹"s�E�{�2�V�)W?'���_qϧ����cl�u��+�����hJ�XþM���ێ�d�o�	ᶬ��g��6�%�SϕK^��֟�Z�$�1Z�滮{�ww^���1�Jo�B�����3�������5�ҫ�6Y�6��G��C(߱t���3�b9*�J�WWK��Xy�r��ª���=�\OO�f�d�>�%�v�����[��c�ͩ�	�R��֯�;�\��� 
��l��`�ju3��J{s��b��=��.'���BC��|��
'����ګ7���]�H�4���^W�J�����r�I��8�}I��c��m�7B�C�%�@i)����Ѯg�^]d�D���L/c�ڼ���D����vkq_R6o�v����YdW1�g�aL�ow8E�L�(/�[ט�����Q�S��&<�r�N�֥L�#f.����G��lf����OYO\e�q7�8��|eZ��O��R�M�ev���ak�U}U��-��Y��h��do立8 ��T�iW�.��=���@X	n.�a��u���2������v���[�\pޏ�I��"�+�Sˆg�� �T�M5�N8z�d��W}{7+뜁�Ʈ���]r�[�:�^�-p��U
��w���u�O;�ರ�Y�--�n߮�Tԑ�y�J��kTF��6�_����_S^�O�
U����o�8gw����z{G�I�R�z���~VO2Fß/�E"xm�b�?�����I���j�j��5�<�x-�BU=�+h6FS�̨ǮɁ��&�I1WH�)	e���5�u=�t�&���A���UG�d � U],'<��:n^���W�+�Ƿ�%��9Om\n�~�ص?t&�����0x�yJ/���2����0)U�d�'v���5��ޗ��{�k����?O�c4�R�<6̮^U�X�0kؙ9��Lw4h����wSd�����7��XSl{�2�%V;�6�P��}~U̞�Vm%T�2&=[Y~�:-�R�#í����/������#�;۪�ؿCWj�޻���ף�uh�"8k�غ�
�k'f�&S�q�I֬"���:d��%�j���"�nʹi�����uK߅ǥm>�ڸP��E�7ҳq��I���:�U�
}L������e�D�t�������w�Si�l��{��4���#>��~�>�k)�W��Ţ���VV��\���#�l��{& �N̤m�E���-��%������W�Ϋ~�L���T���/�7J�7�}��܇�}[v�(X�@��՛��IJ3�&Ry��=[�A��C���L���v��aT�as��}8\�~�U��K@��}AQ<)�$3���G��c���]�|�U����W��7�;�Os�1K��crw��}�]ۄ#�}�
�u�qMz�.�� �2��-D�V��"�_���>3}t��P���ܯ,�V���ڦ{V�Bt�t#%�Lɡ.M��U�xvj�kF�)�Ny��5��t��{;�I����V'��S^�OܺK��������u�q+8t��.���U�0'~4:�{q�޺w�9e�s����2�\��yJ�3�d��/�V�YIAʽy��Dӕ�w2{w됶�Or{��vhx���P���dRzFQ�UB��w�L������W�e���^�DZz;��TL�u�}��6�l���u��*� v�t*\�N��;������Vǧ�Dv��FG+/��YuyQ��vΜ�j��u��N3��j-�Z+�o"ܫ"Еe%k�|L����$6.���G�W����O_�H����ȘϽ���7^Q*�ێXt7��'�����vp�K۽��V���җ8����nљ��|O�N�K�ثIϷ�*>qJ&4�L@:�-`��ye�׍]k���7�b�Yb�V2r��o��?�7��Ō�����VQs��3߻����5經S��h����v�\P��{0iE�{�LO����!Z��ex�c��Z�s��O˕���O�@k>��w�4�:�����z�
H�^7IHW�փ�r��'�/f�w��g��+�&(�yV�nshh���s�%�]�0��uiZ�O��P��p�G��iK���p�p�����K����q���Y������dP>��o�A��ck]���F����x��X*U[����̲�� �\N��}8_�ܝ�0�:mfW�ӱ�}Q���9߾��'�ڥv+���P��ǶYT����'	�,����/�����~ҽ��Ϭ���"�><��`������e%[qv�
�U[�G]����o�9��G�C�����	 N�D�BQ�7��n�rSK�ک�\_{��^E��?�F�i���b������/Q^�q��z�J��7�P����ͻ�lqL�֡J_=�A�*r9WY�'Yý�K.���g����ً��%G�^�+wWR=���sǻ�<֝o�׮K�: h��dSU72�.,�������؊��1e��m�^��e%Ebb[.un���o�\��K�|8{$��V:�|�z�hp"qX����=�L�]�w����懫c��ϓ��d�:Ye}:/���h�na��\F<PnE���<@����iZ�~��n�X�P���e��Bj�����ֱI�`�wʟ��Jq��C�%�������	���>�Y��x��C!<�����j�vM�p��wl�����Ro���� ǣg�c�Zqw�v}uZ������%��Xτ��$��\�D	�̶f%���y���=�0xe�jį��qgz���j��tD���G+�}�<GZ��x\����ˋ���!��;p�lRe��K�9�^V�d1�~�	��r��W��\yMU
��\�gCF�xʮ66�/&&Q�P�5\��Y�7��_W�%��Ɲ��N��B�AM���z+=<���_sz��<�|.�!����\(U�;��o���j�r����Qh�>��p����Wt.�:壔̧�{�rA8�ee�B�|�n�+�)�5��n�VV�[������\�8�����Wر�TT_w��rX��K;��6f�s������)Ж�-]S]��a3�c�J�jR�+���Bl�`ތ~���پ;g}�<=΅��pi9(שuӠ�3U5�}V�d������M�9c�y���N/�C�7���M���h����RKG��U=^ :�tw>�G�k��W����f[re����Ή Y�>�.��)EFD�=�փʳ|U(�yw!Uy�?���{�!��K��8�Dyw�R�N�s����z��O>1�	� v��o��V�a	�v^��F�y4f0��c�&K�~�DD���y9�G���Fv]���Ю��u �XR�v�f�=ͪ�54xe[���^�-p�I��"�*e�L�	7�k��l���P��6z$��d��t���2��Qg-ӟu����h~��4�9s)�=�fT7�e{�������SBi�$]9g�WpWYB��� T��ۯ=�}yt�R�矝q�k�jb��K
;Sܫ��ʸ6��Y+�F�>:)�6�9��(39b�E�xZw��,���Oix����'C�"�A�0�=�S�Ϋ&�E������K�/�vxl��Ր]k���z�X�^�E<�y���x-�{�\���1k��_:iVTI]{+ظh��V$HP��.��g���]�{H��|��<\z"������C��#����h��I�3W��P[�L�T�(-�Yx�ɨ��I]�u0�v�X+Mu����߾���Q�i�nͶ7���D�0��T��WKʜ�ʼ�zjy�������8�y@�˯�Oj������ii���fu����R��<#*IΈ
���5�{��Z��kY2V�mrڴO��;^�����N�����Ln�J���O��z�e�&L�[�W�c`�rs��S���4�}�ac��Ϯ��W�.۹C|tS�~U̞�Vo�\,��>�=4�� h��Y�f_����A�}S��m�Á��|���C)r�\���\�g�D +��qyn�S�3J��+�r^~�J��i����}U�.��4eR�ʳ�a����r�p�/e�,�:y��'��f�4��3b����s7&�X�_d|G�[v�(X��Kl4�s�c�S�l��+$�>=���秲���"��U�g&&�����c���|x_P���Ϟu�~SW{�^��Ek*�J�w��y�};�}=��R�x����?E�N~�ۼ�g~�u��<'5��*H"�A�K^��^��w�������d�o��͈��?[���nu�o�!j+�}ݐ�i����F	c+CmU�dBU\�^�Z�~�F��I�e��(];|Œ:�e��ضR��,t�~u���	1`��:�Y֫m�B�,���3�t߸�[�a	5�d��;�:�z��@�3��t�0ho5�S|f��P��gy���[���y�W�nC}���9?4���\ef�a����/R��n]	�����-�u�N%gV�N�]�����oo6o���{�5y@�
Pt5,��pR�yJ�3�dҭb���[�bPp��R��`f��������W��>w��i��ޑ� �B���/kƥdC����`Ή{�љ��b^/f�=����%W�$6 ��l�ޓ�]��0�֩�7�fۊ�lᢧ�e�����e��D��k6���4�V��]������;�#��n-�&�9p灗}~�ˎY��!3�c��߾��¬Ԡ��oQ�1��[ҕ{�Z��M�a»T�����:A@��pv�_�9g�f��AP�𙸘Y��^��i��6o��1���xo��TE�{��ޑW,�9\X}�*5G�"�ഋT��ʒ�ì�n��rKY�f�Lmw.�V.�ސ]ﶹ�5U���1�g�E[���K
�=5����]x�EM�Wڔkݳ_�<�cb���(��$�����ǩ��ۚV�/a6���@��r��V�T`�!�n�X�����d�����3I�BY��hUY{Iq��ޝ�̗ls�&`/Y�Y�}q��K3k1<uvvS�֑��ᕻ}/4W!������[X�j���t*�C��ʽE�[S�ˬSy==��@��o�@%��AC;+��N�yj��bؾJ��H��O�U�"�'2ν�Aθ1�\Ͼ�y�q�B#����L�Q˱���}~��O�Z�D3�|ۇ�M�(7������s�Y~|���*F�6�7���=�p����xT��u��"�(�#���*�cH<���J��sl��y���ۛK_dk���鏻Բ�]���*u�MM̺�'�*.�<��b*��L�X����g����p���+��ó�	���
D�.����	�5&���/�Ue��n���y�K������;l�6�PSm��V;:Uw5������ã�#+�Ǌʋ�Bx�^����F�֑&���q�.ǰ;s+�t�zh{��'8Y����U]�F}νo�
�#���[C�)�F�_��*
�H��_|������^�y�z��(���t<L�z��g\a����+(�L@X�τ�mY�֠*8l7>k���e_*x�z�I� ]�\��ԼF[���_Xô�E��u��{�ɸ0��˙��Y+hr���wJ��%Y��U��4#�&p��r���_`����s4X�M(Ӊ����yOM�$��/����iB�����:F7�v�z�[ţ�'lߌ4����w(y��}�_!·d<�z��=��_�{ꬡ�����7��e�����<�<~�v����F���b����9i.�YFF}���ƙ�"Qc�W�� *��
�-��1h����L��GA�,��ba-^KP�c_���W/@������)���5�xL��(x=����ѽ�_���>g)g��6�1W�I�y����Z��[Uʇ�B�*�/�n�+|����X5��릷��1��<�I�G=^N>�����^9a���iİ{��}��Í|�UnfA��nk�$������%��χ���;IFbV��2�@_Ժ�}��`�&���l���㳯�k�Y�V��}�+qX�^��H|#QQ�|O�9}h<�7��(�yW��,���+�JY��b�y��H�>㪽�4���w�d��p�޿}�OHq��(%1w�p�&�{W��{cr�5ߖ��[��.ج�z�oڸ!�'m��6�t�f{���t�`|f��Of�>��Y��uu�}�"�U���qA�~��|��e)�^�\3>w���Ѯ�d�������)VF;�1\x�2yL�|��rE<��8q��4��jx��.V���������T��)P�
�ot���ʋ#�����Q9�v�Z.��eNm�Ep!�+0|�.]��:�=�s�唫&����N�t�-��yϷi]8Rݕ��ZpC�YF�G>�j�pp�]������W3ji����A���9�����L�Vq�\�l똻U7��9��h-�"0t���\~��d�[R��ͱr�!�SɃ]��032jVP 
W�V���~]雈���N_F�1�t�V����5ܢ|n#k@�ǒ�C�u��4�g/��K�{ǥ5�԰�
��*ҵJ�_feu���%�|�+��{�к+a*	o�j�}Vv2�$�L������"�T@Z�g��w\�~^�wW�ME��'��J�j��]��ЧK��	��뻫1.�ir��[�"y.ae�}��;�yMS��6d@Mn�ά�Vg�c�:ef���b�oON�M!�1KT ́5�Ś�N�>����</nX�b�]/�J�K&�v�*u;�&�-�C�W<��ց��`���<��26;���g�Q��f�<�p��lJ7���C������M){W���n�Hs���脄V��Ś��5y���'��M ���3w���v�}���u���p��C�ZӽJ���kr�j�c�m��W-06_u����1iΗ ����}��E�1m6����rS���tӃ��y�'8�
���5���C᭮6mq�>��wV,P�i%Y�8�� �Xxf^$�,�)[�rgZ��'�(��pr�73����J�R]u�V������ �wK!�)���S�[u{*Q?�V���s{@�1͹��\gD;��)ekv/�Kc�� ]�}�׬��L�Gݶ�Z7���ʄu��j|��ӾC�E�����AfҕK莶_U�
7b��w����j��v&�ý�6��(�';*@f���k�)
����w%��Ne��eϒ���s�oE-�V��2[�J���Ρ�>�v��K���P�޻A1�P�`Տ�P}��[Z6P.��ڍns=����Y��]*a�;w�]v��{4��0��!���������q�m�Y�,��pI��n\���Ta>Ӌ<�k�����ʲ�F�T/��wpʈ��M�Loz�b��'8Ә�>�-�����jN��S�8�nS��L����͜לfu��`	��v�<������ʐR�W�9v�Þ-�)��o��ʚ�"{b63]���e	Yx�&���n�t�6Ԋ�BҸ:�s�N�Y�R�U=��x�����0��qTSdc91�����gKFM�;�>���c��];�蝔GA�͎">���B�Z�gY�x�w�ŵ˝L�e�=��{y��7��QGHZF,Ui����<��VeB�f�(�Uqf�eVʍ�J"-b�0�
%�*�[���V�(�[bQm�,E��ʑ[J)*XȈ�l����l�p���QUE1n"V��J1�m������­�Ѷ%-�U+iK-*(��Za���J���EQ-�jE\\���p��U��U%�f+F�[h[�a£PZ��[Acl���"T�l�m��J"��Z��ʕ*��\b`�V�-���0��*�j�Q��k�L1�bZ5l�6����.��cYiE�Ka\80��aj�Z�E*��J���ᵩTY�cU,��,�%�[cX�6�meE�F�m���������I��j�e�j�ÃیL)mVb�4�qG0�JR��0V��jYcZ��TJԴUKkF��R�R�R�TŘp5Dm-kJ���#eRH�{ӄb]��㹗B���V��)��&l�c%�����z�88[��t�n��g=�7���7���cEz��.�%O#۳�(R�{ݽ�]������W3����Y�t�u���k����9s&iүI�}|�������W��A$���D��#_i�{�����G��b�^5Л�u��=�$k����5eK�n5K�ݡ�s�|s�wM*�і���t�6v�+t{f'qR~�)K�*c��Yd�7K���HH�P�rǋ��M�gU�����/��ԓ��/�j��v�9�r{��aB���β�@X�� ,�t�<�Z���7/MO:���lkGV`H���왼� ��Sx,<۬�>��3+�o)@�U���Nd���x3f��e�3��{�%����J~�/S�t]��NxӘ�p�q�YKʽ3(x*{'*n�;��]�?m��F���[8<4J��������/'�	����7��
�t���|M'�<��l�d���R��VF�����.*aޱLmV�?Vv;���됏�[{��(=ɾ����nǥ_j�~f)��p���p�U'��8S�>F���砸��^�r��R��իJ"Gs5�v��pDՓ:�Xl5��,�΍~۵ە�β;0<վG�Cʺ�b�\ ��T�2�
nB��U̽�Q��'�w3 ]�-��wmL|Q%`� ��}�Rx�k<6�G���p��𩋌=�¨��<֑�m.L�[d͸+���<�ɷ^쏈�w+nޡ�b��9�qv��ӟ7ڧ�H�:��%(hX풼��<�u������lt/�;�L�����~���MY��߷�h�P�N�`
�}�iWe�Ī�&���D
{�!�+�ȼ7�Ӌl:v1�6Hy��k���0��d��kQL6��A�K^�ո�s}E�Uu+����+}�g��x��ny*hϤҘϧb���$��X��*6���F��GF�H��LIÝ͹�zw_TM�9�l���sX��v��*x���_9d2W�/�׾��*�'}Ae�Sd޼��k��88o��^P?}
Pw���G�d˂�Uuת�(f�����cei���97d��#X��m�,}�;��ȇ��A�ͦ@��u �B�g���پ=	��Ι:,�����K��p�lS�k�%{rCc*RzNt@n�6^3�y�ǻ����9H��r�E/WeśX=q<Z:��O��v�So�LNuPU{��B�]���%���QB���Z��*ed�D�p����k=�cb�[����n�D��q0H��n�9֐���߽z��¹-7�7)����x��J�*��ܣv{R�*�F��u������;/�nu6��VHX�uF��M��ѿ� �������s&g6�d8`�꾀`͚���V=+��᷊�\Lo���,g�%v���A��ivTػ��Z���Gݐ��{�%Xp���<πٕ� �����ff�af�d^�L�9���{�G�z{�oli��D�E��݊ͧ�0k*k��?��@|�z=�6ʡ.�~t���E��5�b.k��z	�=^Y��f���2��&U��=��鬚��u�e+~Pic��oZ���c%o>Fp�Ez���x���N�xt���q�|��>�����<r_^���S}��-yٵ7���y���1��%|X��a�YǸC
��pc����.��z.Ũ����z�����˞*��p�r�m����{
�yo�ƴ?r�^��q��e���p����5�/���UvM̶s��K�X�r�ӛ)*�k��S���8�ե�ڝ�W��\���q�Os�,��]��Ё��Y��ˡ���:��bl@����m�O@�s��"}:�]�=���!�phR%�J�O	�5T�F�_AzJ�ᇑ�&\7LP��p�i��b�/B���yVK3�dl�7�v��c��0*��������ul�qo�O�A,����j�m\a�xO�bE�w�umӾ�w���h�>��S��+,��7��c9�Vٱ���}�u��;8_Mݏ�7�L_����O�򥃝E��uSQû����x7��64FW��A��.`W��l9�o��g��s W�<�4ŉS�����Y�BN�Y�ۮ��ʫ������6�;���V{��<'i�g)����	�(�4V���xg���w2WKX|���J$�]���̖��^xf�9z�j��ԑ�}#;��
CC��_+b,�����`�6�=ϯ',��ay�K4�3��M�t���=��Ĭ6|�J�@^G���*��_��r���;3V�~�O�>綸�:<"ޘ{pO�yo;
��@jy��Z�u�]���{�f y93S�{�$��	�2�0;~3�S�>s���[k>�p�}<�T��q���Z���������.�IKΰ���)=o�J~>�Nގ���>f�k�+ƚbf*���r�Y����,e�o�蕷���T�3�/%�%]Z�A}����ª�̃�����f;�Ƭ��Z~�������P�ڋ7��ϒZ=�
�� C��+�]��t��Uck���4	�UJX`n��{A�Õ��i99:<��@ow�<�W?Z�]Z6�֥4.�u��0�U�\-f�WX���Q|5A��8�Y��Z_e�dz���&eg,;�5S}��U��P�R5���m-h:�x��Y��\��#��7q�<B��綧�ӑY�Xy���R҉�ϙ�>Q �~�������F����ƏW�o���1�X�T�s��T7�DjL'�"{L����ӵ��Oo��/�s8"��g�˅I����^MJ����{+�zˎ�	ʺ����g���|�)�}�f��J\|��Z������|�Nx�R�O輪�d���7E��qI���b}��|H�=Cyw�c}Zϣ�㛃�C�lL{i�����3w���SFY���Uq�䑿�5�ޑ�Ӟ��ߜX�C�`xv*��J{�j���,][4�Z3�vQ�ϜU8��z���>����&{v�"���{Qf���qv��X��ƒ�g.;�ʫA�H�>�f� �*z��d����UW/��c�c�s=�]�"\�Eͫ�SJ��9^�D[� !��U � U],/��ʼ�g�|ZAm������|��U�|�`�%�}SOf���်�~�C�8��~'z )}U={1�������U�U�Ս(ht&�<.�'�%V���=ݒ�N�c��^���)��'{n�#2-�N̳��AC��I��m�z����}��[]�-V��\�i�r��sJ��̟Q{��2ƼS0.̻�'�,'C�q<��W;���Ļ��*9l��/��Z~��h=��Y,ԩ���]b�C��
���e����g��et]��6��z���堏dƃ��/��&x�d��0WP�O��I|8w	Wp��ܮ{7:�Y3�j�c�ýFiо�ZLU��C,rޯx�&�a���Zm{[��sYc����W�e?3�����/F�R{�)*���>Fe���my�_s��ww�y'j�)n$z��%�����������_dv!�3�~�C�^R��Std^WP;�iyz����� �}k�2 ��/�z/���׳9�k�ry;q���m^+ _�m)rh�{;:w,C����"��J%L��w�;bo�a)�x�)u�}+�s^z��3w�8���|����[=�8NF�ߜ��T"�A�K^��ņE���+k6�5��p��CS�x�;���j{�&2v+���,�w3�E�\?Q����s�qټ#����m'�{�W+�_K�F�w�.aʋԩ�9�t�Y�W/�YT���PXQ���k��j��j��n'�؛ti����+V�sB�]3�aG�rC3rڟ(��I^�|k��j.�Y������ŀ.�mv������]lz:_^,�!�_5��e-�U�y�Dz�m�*�� �n��6͍�M�.�灳�{X�)��{q뻠2W\%�z�ה�B�K;C��\��*�ϕ�J���ZUa(�"{|�o6-���s�S+�o�z"#(A��`��l��Pf��� �>T�:oLy�F��uҫ�ߊ����-�6����>�yD����B���AoI����jn_A�ۧ{I���>���0קըm��<6� �%C��4�b�'y���ĝn\���8�s�������A�,i�o ѳ9X�Ƽ&S��P0w��75('�oQ�H��]����g\�OЊ�{�|x��?�v�������*��w�5[ouJ�^b���-Z�K)q���KW�ʍ!^Ǫ0k>��w�d���vk����U	u����<s׹���)���1w���^ې��bu��=��鬩�N�P���S}Z�3��a;Y3����z���f�U��t(��(g��g/CU�8��wxeT�OOh.�!�ɓ�+�P�xw��,1>\^��o)w�b_��KO$��z��*u�����R� ��W�aU=k�i��9�����$x������v�qܱ+7#\��V��i���t�/Fߤ��yZM]}�,!f�zl��FY����ed��Ӱ���ڙ�SeP;tWJ�/8���=Y�^<�6��s4��q8��㶞�׏���it���.䳢H��S��'�z����U��F�4W�͸{���oaTÐ�r�Wu��G=�Ǹ��B��؆|<�T�|��n�y+��!���*<<�sc�s����YB����9;�L@����=C�m�|��~C�kq"'}��0k�(-p�	z���,̝�v<�T|���<�د���ip�U/����3��m�=F�ۣB�#�
YCkZ}׷蹼�>Gp��n[&�t���}��v�vS70���lk���+j�K�u9�r�����O*�r�������{E���=��Xmߡ��)��cR�sǆ���y��cb���������(��¶8g�C�o�2WJ���J���K�\L��w�d<��Q^K�O��g�)��>�ڳ�@T
�����%��P� Z
�����u����x���V�J���S��K�t�t��V�fXc�7�=�Qw�{�7����f)��_k�X7�Güm�<09U�0�� �Ry=���@j�����!��[��HoL��ǔ֋FIƀ*��+�U�=�[xQ�����d$G�u�-35�IF� �^�մ���¶�9pxJ���U�Ғ�[�����)�%�.mձF�=�2*P�s��#Dݻ\&'ug1��bf���*v�jY]X��މ��]V⬜H|�����¦h�	��g���tAYVw�)ʍ���G�ػ]��p̹��f��a��$흽R�^��kP�ֶ��+1WK�t0W�����|� ~:�]A�:�����n������ٻ\7eC�qW�[yK��`���h)������_�{[���]m����\\��xq�~0F`��VL��ʫ~���Y��V���O������.~���07jJ�Y�W'x��+��j*����ո���Ȭ�,<��Ș�y,L%����3�W���b!�y�����x�$h_1ֽ��Gko���1�X�ás#��qP�ԇ	rP2�GA���n�=Пx����yJ�0e�~9��c�!��Ѓy9�G��e��+O����������^�i�]
�
t,��e��E��`�Y��}-p�T��R)����u�셗mj���<\�!��`�e�&���%�4��U�X��zVbζ�׵-p��u��Y�9w<�<��V]��R�o�||:�W��E�j"�خ��ꬁSUY|v���kM�;���YH�'x]��B�F��<í��ە�M�2��`��v���G���Ս+u�58pk|���6W`��ܙΐkY*񌘱�Gt�nC�Es�5�i�Ve�M��Na�`|Agh�p����m
5|�P��O�2��(Ɇ����,����S/�v�����2��J�c�Q��N9Qz���6'4e���3��2�?u^]����|��;���v"J*��#��ͪ޿xv�m.0h[j��G.vP˽^^���݁���U��X�%�W�y��# H o�,*s�*ܼ6��`�⼽ĩ�:a���!��ļ Ϧ*�eU�gҵx`/5����>�7�9ei�vv��U���4^���h�ٲ�αn�j�=�'<G������*�_/j�l�q�2W4��L}�x�{ᚉ����߭�t�)�ȃ���.K�yx?�7��ய���W���k��Q�>��ͬ#��4�e������>\;�iЫMi1Ue�n�z
ƀE�_u�3�ݖ�^����#�}W��3�k)�.x����/F�Ԟ�A��>�ϑ�f>)^�JTS�z��ٳ��[�)m�2��Br��)Qs��O]?���ꆠݷ�lѫ
^%G̅���~�5�W��[e�jOU$�pX풼�	���O*�S���z^y�گ�W�q��&�R���%����",6�ղ�P}}�R��Aq�U�H��
(�D}�:
������χ,[����kL��B��ڝ�#�\U�Wq*r��36wt�Z�j��;�ԫ4ǚ<��+N��������	��v�(2���b5phO���0�l�,�n�_M�[}�P�1�P)�7Pa�b��n�x;L�Ӵ��w#��}��	��r5����`�,�!�����&��Ꮊԁu��v]e�طz�ĺ�W::��V> ˰�6�*��+���y�M�d-��w�r.����Sl�[��8���k֋��]���K+#��zl.���U1;�A�g���B��r���'$c�y1���4jy��oXw]Q��Z"�l\�:��w��-=��ĪV�⳨h��Oj�8�&L
�h���v�ټ�xW-��3j����>�`��Dn��G1�[��3�g.E����޵\f(�#�
d�G=
*����V������X��3���G@�rw�@�*��{�0�\a���M��m�k���*3�]DKï�;BeǏ���:�aJ��[Sۼ�pe�cR��n
�=X�5������v�)ξ5A���Y�I]d���^ƞkzyLS]ީR��Pώ�W�o���禳D��Y8���Ot�u����t!��+���<�X"�Mjn��oUXR�[ob�u{��J���\v-��X�ٗ(���鏬ӽ���
�5[��ؐ�s��eIgq�Cr�d'L��Y�K''q��Kz�]�j�sߺ�Mh�v��e˚x�7�V�04M�r��%g�-A��ui��&���²s�^!eTu�.X���d����>�-=2u�؜$;�����S�a�
��r�*��t����ǭb3N����1e�ݐ)oe�pU��\����<Xs[�U�=.ޅ(�YO[�;�V�M�X�7��m�\���������s������LPFz�s��|��>���V�����P�Y��Qڊ5,�dl���$IV���X��#�U�}]X�q��S|��pU���+�7���MkK��CzuvX�3M7}M�S�a����u��\���+�Z�\�ar�^��})��a��Q$��W32�n�u�Tv�n�d��u܂�s+<���|�C��l[��ui���7km�x�����Iռ$[Vp1B���B�]W��֮�{<��y]�5ㇵj7�T��8jZ�_Xg(�VpУR�pL<���1���3q�-�1�1J��R��X�2{Gf[��I�cN�o�hȘ7����:x���Z�����f5% %)�y�F]�I��T���־!����';�y]b�`}qQ�wt�����ӗgVd�2)��A��f���8l�K�wAP��Dޙ������k����ؕ�r���!ݜ�Zz���dYwL�E��P;e汙�Zg_$vK ""��4�Fڬ��cq+L7
��p��Q--�1�)bQіZ��%����ť-[iF�c,(���b���QUUTih�ZU�jѶ�����ٌa�KU���5h�AJVְ[X�#1nm�j��(�U�ElbԢ����%hJ-�c�.1c�jR����B��QÇ�D��XV�����T�F�V�-�j
�ʖ�j3����V��Ҹ�1Z�Q�Zʈ�cZ�-*P�j����h�Fֵ��m�F�-�JRڥ�h��eJ�E�J�EJ+j-J�4��Q��Kcm*�l���4�Ŧ��+J�E�m+l�kF���m�Kh���1�-V[Z�E+YR�T�)h-�)KFUD��0���p��%E���m�mZ[h�Z�P$�4(�Yg8s�e6��N-���S���ʡ��ɘ�`GUu�wB����Rǟ.��Y�,]�@Y�!U�L�o�@�Q�ya�/��6�����I�m��S�İ��Uz��X�A=�!����ɰ�o5<�{<r���\���8>F�ߩ�,��\������[�w��cl��¤�mqW��v�B'�
��̮ÎiLNIP��#ĺK�xϕ��]���s�9�U쓽��w:����̏S�<οq��.a��˘e�]=��ˠ��*��i����J���՞�5�)�@j1+8a�Ǡm]q�-��9���y�<�:��4�&�ɄOZ$��u�-x���w����6�:�հ�K�_�Q� ��Q>��G�.<q/u��ݙk���������u/�1�gn�V$�
�����
[��^ܐ؂ë��z���)f��'˅��m۸�If��ji��o�<-��~7�F�e׉�m��l�癅^)&kX�RThy6z��|G[xݻ�~P嚿!J��;u{o�,�f��ƶ����{�=�hO;�K��J��Sٌ��{c�43�y��*5^Z`-vy��.�T,����o�vz�V�5�⽘� *v��ɭ*T�=7c3.�6:KY:�6�u���IxU�ͅ�Uh\K�����qV��KS=�����Ŕ�u�[�3w��h��1�!��e)IV�Kw3�C�G�,��\��t�4����K�a�s�������ec��f�Z�Q�+��Fd�3��d��q�ڝ����M���b��y�3g����Y�O�δ%��n��12����tT��T֧u��.� ��:��n�����3�:���9F"���C�|�ӫE�bs�T�*��]�^�L�vwj���xm3��ު_�� ϋƓ�aB z���1�5j�۞GOٙ�����Ss4��R��n��h,����3�z������Q+�䒇��"PoaK�5����)�_o��yON�y�⧟b<�T�|��⫲ne��]��P,t&����ر��z2��n�v˷�I�F��~�*���(���4WF������R����.�ƹtǽ{�������K���e�^����]4�L���p�I��{������P�=@��d��%�el�ΡW^f�߰F8�g�	�s��U��ުv�v3s�P�����Ec���p����1�����D��B�5إz�lW�i�sX�N�Y��ߡ���Z����Ԯ�\)�c��構˞��f%���Z�fi���8�L�ZRT�.k��sX���k��].]u�t�;��m�0�R�i�v�X��uww9�[V���tfA`�_Wi�Lt/;����l;la�j���У��hwW��6�ىE7�z����[����:��u��0A��D �vVXد)9}�ܧ�ZD��>h��zZ�k���[K2�36آ���C$��S��
�r��!��Jؖ`���gֲk��s���Lz;�xewDIU�R���S�!L���ŝ�lj��tD��"�i��������=�~�ﲕ�Y�z����Y��[� /n *L��/���������"O}k}��g��l����2�_�.P�Y��{mW����P�Ǳ���T�ɴ��}�Y��9��s]��,�8�����j��Z~Yk����L��[7]�e*^\_'��wL��cۻ�9w%�yºe��2="޻7k���N��o)w��{�!��)���c��k@k�^K��l;�;��S;y�W��=<>Ⱥ��Q��VI-��6����]>6Z*x�Oݻ�w~�ܖ1�`�ju3�����>�HtL�EF� �L�������%��v���;��4���#~�~9��!���z�},t�=й��ݸ�o��C��n{򬧪��P0��p�?f��F�be9�Z<�U:��)�`���¢�r��%���n�RIzxz���_���2��ڵ�앇sf����]c�M�;t{�KU2�/���Q��O�e�Y��׷�v��tέ��4ܦfU��771�D7����Mv�j�@&<,p{���~9F[�OQS��1���ڗM� a��Φ�W��ֺڼ�dڦ�t�K�w�bmz�->q��S�������\z�T���#v	�7:{-��sٚr}�Pd8 �f��9� �7��p����Y�t��mA��x�E[s)��3ǋ�>�s%���2������Od2�/R�>�đu���خ��1�Y��2���Cj��zl��5���0����}�9U;�5c ޡ�{��q���U9�-x���Y|{�o٘�k��mtk�(Pa��go�Mk0t�Rt2��+h',x���eO3�Ƀ-K����sY��d��kəyz<������">�����
��d	`��67_�6���e��W�rK���|�1QWVD6��֚�w֯K�< �̮�4���q�kT�H1�lM��z��m�b���5�v�i�iڢX���d5�wLo�:����^�c��5=J�U�Oo-��Nz�����������&�g(Qϻ/<�xFo�ӈ�iz��r�Vw��F����A�z���f1$��_�����CQR��S���8��9|�=�٫oi�q$~{��v�hĥ�\ՠX��r$��&���g=��Ȏރݸo��8u�N�y6�����N�c	S���u����9�]']Ը��2���{�n�]בs]5�;V]*�gmt�x�w�[�R�׵�E�{eCZ���%�������^=��D�w��z�ivOv\dg�G ��<�k)����P���U{e�[̻6o��:��]�`��sw/�j۵k^�y�,T{��ܗ[�;�<;J�7�}��!�3���ckj��g��5�oMJ:.���՛�yIJc�J����9O*�|�v0���l&{�5�e�{�o9�nV�V�:(�pJ��U]T"�����Ћ��d����L*~+�2b�k|���Rczw��}� ���T�\=f����Y����yC����m#�w�P�XUS��S���]��c�v+��,�`�_�E��}K���ɓ\&nMwckҨ�~�.�{״����^i��sXɗ0�ʺz���UNY����\~��k��t#|<��pk�0Lb�J�\{#���tr��/��P���I������w���{=�k��!�e�\a�7�%�b��@�֏f�v3i�$�F��j��z��%�D��.X�ڠ�f���z��ʑ�۫�0��9����w�۳WC6CC@U)�X�R�u���-�%��3J���rX�%�GAژq�w@���׺1�X�l-��F�j\zq��&�����"Vv�ԟQ�r���uq���b�NVC�M��]#�8�|<\��/
��ΔK���@�ޖ�o���-�����-�9�h{��W��.,��U��m�0�R�����/��^�'4��<��8�
���u� ж{��L5�2�U^+qpJ�Tv:>�.Ry��ųx��=%�=C'^�[ҕ{�d�T��x�T.���,�{0m�j��FW���ts]k�ך��8{��#kr.ߏll�v��X���2G� >
g�{
��%��=,����5�o҃���Cq���A���	t�12���EOMeMjw^��ٷ�U�*Z�O,��j(nJ]�0�n*�+e!K��y�W�K'C���&�������N�xb�%{��{~���S}b,[�{K�b�!,��c�j�2��m�{g���gL⬑�>���qs>�����Oi��Z�>Q��<g,��4�����^?b����ÜVK��4y���~}�g����Ӆ�b��x�웙l�d:T
��/v5I!��6�;�p�emldV.<Q�~\�{�W���+!�X�n��`�8�@��ʸ�ŏ�엉�G��>`��iB�N�"��N{m��B}}�1=�t1�{�G��W�����%v����K��%��CXw���qI�jun�W�d=�R�9v��g����p�Ts͉�(.s���8�\��;�w�����dSSs.���z���>7ޯv9��b�(��>.��Yl���W����;�䘙R���38)��s��>�`��Toj�zcڼ>����D��R�_y�\hz5����%�u�{S�:8�e;m�$��q��%�|D�-9���� R�#��G�u�봻��d'N��
-�.�3���d;�#V��oO0lmIu������D/��7[����5�5�849�y�L�)t����v�$��
*��t2���VU8��ƚ�c]ӵ�(�:g��A;�d��l��Mu��oeb��[� k����[A�ܦ�&��*��40Gu�tz��y��%ə���3�8��p?+[���:<"ޘ� ����}����
�O�	^�u�"�L��W(Cg��"e3���獇\�x<=
߸��R����=%8��N�M���b�o�Z5����ƑT��}�˅U�:�+��E=�̼��%+���W��Y��ӫ�]��[�2�0��ЄZ�8f�Z�^�Gf��ƳH�;���^��Qc�QGvk&Ѽ�z��4T	\І�qr��[��O�͘�iU�t�E�l����.��������5��AF�BOgfLA�Գ�6�{73����r��o�E�tǷ���V'��J��1QoJ�~�V�2���՞�s��<gL�_FU��oň��S��씺�]��r���Ė�]��v8��}���f��� UX`�S�0�8�b_xʜ-��R�EFDĥ�ûY�hB�t��ۜ���4��M!2�2B�~8��i�w�CS�өב�^�6����I�ғ�|.5�{�+��%�fY�˲�ܷ�[���/��2��}8�^�I�ܢ,JQ���5x+^�l���P:D�����&�.E����̸<ܵ��a
@�D��5�zV�������3�~ A7���%��Ӓ�o*�,o��G�B(�K��9��n�i'úu����.����T^�I	�z�خ��1����f���Y�}�6]���;�Zݖ�"��J�e9e��N9�^�T�&�}9�-R��;�LVf��l��zr��K�%��,s�N(&g2K�o��J�I��,��	�)�fT���-s��R��=N���C;���X�b�(������b��z�p��^��GM�5�
�~��M���_l��9�,wҝ�*�;T��]:���"Q���M�����f��k���X�n�Q���.��oyں]�c^��������3��S�kiC�����#*��Q��D����H-�;]�����B�ݙ�y�����u��:g�!ס�+�l{}IA�ͺ�|2���u��w:.lzD�竳x�/�����`��{��钐�n�j�<S�iW���hf��=u&2�z����WSX��f֥�2�Ɂ��(ײ� �x��.K�yxQžG�sոyX7��X�kO���(;�9y�����yjU�^��=j�C�v7���=b��M�5~�3y`�4��6�z U_���沟�����þ.�{e���;qO��wL>c�k��.�2Σ3닁��_	�2_���\�6�Ӆ���Jd�is���f�������ib�|DkQC:�k�kԯW����u����˲}�#��vL���x�?	[����=VT�����h%�H��6"׉h�z{�n�"<V�ӧ l�l�[�U�ퟫ����=�K�0��Ϸ��A��h��b��F0B��~�-K��\�i�z޻������Q[�gxj���ڹ;Z;�b�3Cs1?�ye�3��0�1ꚬ	\�k�t�ƣ��gg�n�9x������)�ժ��4�Bq��[�r6�Ɖrym[�={^8f�V.����O��Ο�b�Zu�-�6����0OsHw�r���3+��9�1��]�Y*�f�軐�q/��c\�����g%7m�oN�y���-��qW.��2�yWM�+�7��ƴ�y-��|���B&_^��&9z�	j�����m����Wc��Pw��y�����9罯=���NW+&�8/�P�ϒ��V�7Ɔ���"e;�c6��k��71��o����ā��i!Pe5d:����Z=�o����?	���R}��d�,g�G����=�t�f���KK�Q8z�<o[^C��類����̙�k�=�睋3v����Ǧ�޺U{�*)���P�Xӝ0g�z��C9C�KA$�ݽ�&�oJ���}R�c�5�-[Z�d^hc��W ~���@������]�â M���Vpy{�v�r�j��}pL���4�;^:$#�	�F��e=Q�Y6-��/�A��G�r�9E�����v�~��{��ZG���T=���w'j����]�b�� �v�ؖRN[t_YwؕL��pdK[j�#�@�f��,�{��[��7�&;EL
��`e�uۉ+�WQ6��&nl��5��gR�I����mi�X�gh�g�c5�D�r�fI��f�u:�*��w+�����@��"���s��X�]�Hk�ފ��)�(zN�9zͅK��
��f �ܓ��B�S4WU!�ۧ�*E�󄚗����39M����	F�P̭	c�-��@j�5�^���9A7(ܭ����To��+��kU�X��6m��I;��6��u�L
P�,!�!�����N�&W#�g��k�*΄ZJ�y�t�2�P�X@��NW���%��6�j��eq쮤��w�*m8���s���9s�d"+N��{6v'���7X��B� ���^2��=���@�	�xEd�����AR����Glu��۠�ڲ!���T��C���m�ՙ��T�H� �:r�]f�ڊ$��:G�j��d�[��y�lV�Ŷ�U�ݩ��yq�a���j*f���ԺuYẑs�i�=�������+��~�V�����
�lR�V)����Ս���i���� ^��X���h�Apu-�{}��8Iv)�_[�n�.�v�Mu�Tͳ���)���J�z(�M���Sv飵v��?������n�8��ڒ}���j�l[�Y��\��1����u��4���^��e�zJ3U}(�OM^���YmIj-"���q�OCݮ�һ��%*Q�K+h3w4b��j���I�!�6ʏ9��VI���t�}b�m��� ���+-���Rq���(�ެ��r�����6��������*�{<F����q�n�ڸR�[؛W�$SHz�R�cq�b�3�M�sF��O���_p���7�:6�옩�º:��°�J[&��Zߒ0K�&Iw�ڇ{M��:gx����ڐ���Ɍc�5d�ѥ��aPpۜ�㐬/89�I�D�����f���A�T�Xk��:�\��2�}�ýi���̤�\ce��Ti����N�ݍ���6P��U��Q'w(���`31%��o�a�����+��+'YL��1����v6Pr�i��m������aUnY���L=�t�\�Mme��y����v-s��WT,Լ��-`A���Ho��X�6�`��4΋f��:w2�9>{Zi����
�tSw����x����s��EWM�;����\���R÷��\س;Zaf���rޫ�ʵ�N�2SL��XR�����]��㴭LR���nA�2��i�&��Qj��ZOv��.��=�+1YL;���x���c�a$���n	��*sO^Q�ŵ{v3�a�3���u���l��CJf�t��&��w*��9k�U99����w5D5gU��@�ֱ��҆>�8J���X� �����x�X<"��id������	(��Vҵ��*"��m�j,D�R�ZV�e�U-�����YTU��Z��)Z"(֊���5DP��-kD�Ym��m����kKYk�-m�EYm������+P�mm�A����ej�R��+h�-[iQ�R��(Җ-b��ET)iim
�[kb�al-e�5Z�kJ4��Ԣ�"E�ڵ���J",e�kZU�(�JYQ�TKkR�-�*�X���Y(��ֵ`�iQ����-��£jR��J5h��4-m$mBҶ�F���Dmm���[YX�V��e�e��V��J�F�F#F�kZ6��
%U-��Ҳ�)iU�JT�K�h�ڪ���mKR��DQmb��A�j�5��ZQU��(�ֶ�(�mk��)h��hZ
%Z1��)�U�[V�+**��*V��Ģ�m�jR�TUm*��)J��`��[jU�
���)m�Q��Rڢ��~ ����վĬ�w(�w2�������,$Q=Ҵ����L^��Q�\��y/U��t�s'%1�f�g�L����SRN�m�����w!k?c3��c��b���B��� ���	��H��"���o�zW��F	Uת�7��u�P>�)��J�Ɠ��U���T�p�.m�l`��/3�a����v3�W� �\�&2h���&us�A�z� �I<#�:��p��y3c��o��*�þT%�}<��g'��V�9�l�vC���;�=}׷��dx{�:Ɛ�Wu<��u�W���%�z�k�!�5ã"�vVWJl|[Jg���(���B|]�ulE��U�°*�i����Hy�ww��7�*"�_��&f>^n���Web�0Ե�aþ\������E]��V\|\9⊈���5�<%��˃r/``� U�K<
�ᶩ*�*����,O}�B;Ҧn�w�J���X�Ou�4�P�8���jO�̨�dx1[�Ycb���k��V�rHs���s&���\Y�S�ٔI_7pR�t2���S��È��;�2��ol�uW@�i^���@���?[���7蘚O޼2l������-��X����Q�p^�J�Wi���xp�W���
!tK%0�X���p��(}n��+ݘ;�I�z��33���_F���	Z����J�y"��h�
�r�-��=��\�W�v+�`�x�;��{\�ET��U%���t���%b{���g�Nr�m>�K�ͩ�Rތ�-G�{��.�R�Z|����� >w �T������Z��u���
/{�x��O.5�y����	���_$�Qk�x^:0<~=�)�Y��:��u���{��D.���-����s�xNͿ�\T*f��Ϩb��C��B�Kz�*� \O�vs�}-��W�p�pa�<��&�n�S��g{���O�̫�4����]<3�w���cg4�u�+��U_<�=��Q�5���~_��H�+�n�r�O�sz�g�=���q��ΰ"��
���{pP���ϭ@:�"��z��)�R�y#}A^.�G�]�]���{�y�����e�H^wO��S��VT59�xv���ʵ�ӽ�n2ow�{�iT�� �2���7����X˖¯Kb�����~��w�_s�N���q����O��m��
t8V��4k{qj<3�<q�P;�&�G��Xk�m�M�y�͠W�%��+�]XS��7aX{ߢ�`ԭॽ�0�iL�n�G�V�%	tj�S�V�Vok �kUΒ�p7�v$1Ԁ��=x�P��͍p2s������)�:}g.�N͘���{`�r�^K�[gG-��֙�`܎��Ǥ;f��|�^����dq��j���X#NJ1���;�����ylq�4W{A�!/��K\4eIu�\1SH�J0�S� ��S�w���]��E�~�A��4�t��,���6��7�b�o46���=Qz���+'P���T���n����g� �&��tX���㷃+v�(t0<���ȭ����mBh�����ȷ���uY<2Q~*�_ʻb��,x`���� ��C�(�����U˾��H��B��P���!�����>zo,Uq���^��`�3����t�>׳^5�n�"}�ו+�����U�d�=�-�i'�߆o�?�ݮ�.m	yN.�\\�ۊ�Kn��S2���l�����|`ѣa�C���2��s)x7� ���=+��ϯrM]�wv�-�����p��<M%T;À�.�\����_�W�!HOXN�0�y�y��� ސ ���*=�}��<I��êk��M��V�1X�uC;S����F5a�y���a]�Z��j�'Fu`K�vש���ȋ�O�Z�۫o��)�i��8��:ޕ3qż�m��kK:�, &�m����ccǯ���ύ��1K�ĥ	@F��������;f�ꔞW+|/)V��}��%t���l����*�"����!��;���u;*0d���
�K,��u�[��=��!�g���z��P�f��]zbN���	��&T�D��}�u7�v�f��+ٱ,�%m��=S����G�o/x�P�	0���ҹ���ľ����Ǩ��f�o���F���O5aIu�s�����e��
�	dm�hT�
v��;ܒ���2
�����U���;C�����:�W�ev�4�'+�NYgD�_$ۯ;o���#�e0��҄��ͷ���Ox���`d���d�AS��O]���c�*��y���6����y*\=�������%f�i���Кy��9�����pP�>���n�^�G*=�M!@d.$�h�K�6�`�7�_2=9A��d񾱲o=��x���j}�-��=�$*	�+!��9�w���x;��%���$�(y�w{5=��R�m,TL���lg̠�)�9�KU�2���S+�w�43�ه�������D������G ������E�9��d�*Öi$6-e��D��ܝƆi5/��)1ܜ�]+>p�VK�����;��y�ӷ9�\���F��4z�:d��kV�v*9Zl'���)���5����(r�M����5Ҷ������o�|ΣKv*{�*)���	��9U� о�[!�CPzV�H�l���b�9�kq�0����V�Ǆd����9%�<O��vX˸���&�zk�����j�;~*�
�mC�B/ׂO�HW���Ϧź`ws��C'�Vl^|���V-ƨ�a|��w��C�g��9��bg��`�F��Y	]�ɥ�%�Vk8W�N�I����;��u�^�me!@-`���|��p�3D��I�o<u3�+s}*�G��qxp��j�e|�'���ޥ7�)Tb���y�!�<n��*zY�N�ʄ{c�3���Ϧ�*��\�c���<�a�W<T��<UC�|�cx(�EM�f{��k�[�t���,m�\#j��x���C��ϧ���n�i��f���9ݾ��U����k���l^ת՜���;C�Tu!)Z�[���o�XX���p�8�UÇ��;|���k���3��45D�\;���Ֆ�U�°.���kK�ʗ��Vѥ�^�C��f{Cjx�����͈U�Qi�%����!�%_gp9�C]�3�����a㗊k��j��`ӷnC�Nt;Oq\̬��5m�'BG��"�M�f�����;t����n�K-�;Yx�#i�g8�F��c�.a�d�Hٝ39��m�{��\�l�]��:4)m,I�Ե�8z��%ƽ���N(��{;mt�M=�+!�c|^�]�{��N�։sP�j�6��_�S\�*xʔ��Ϸ��e/v �1�z�;�i��8-��u��2�g���UU�6+^�C�]rrl���B���L���g�2��yD���J�I��,�՟8�ЪFw�b �{+�� �[��X�e�u�Y�0u��eY����%3xP]�h=�Kg3i]�9|�j��dx�$Ω.3�YV��k'���|b�b<=]��ʡ��-�^j )r�~��Yz�|w�	c����a�y����o��b���	�e���ǲ��>��ܞ�����kD�ׄe=�[�w�\�\~�z8i���a5��`�u��Ϋ��\�&Q�iRv�AW���}�L>�`aT�PW��Ѻ}�g��+�ǎg���v������g�I<r6.�r5�%V���2���ce�T#0v|���e��ø�8�h����l.���ʦY`t��*^�hS6�v�Z��[~j���o�Z��vR��Y�p��8� ��ë�Q�����5��dl�ћ�ն-g[��Ry�.�x�R~����T��Lw�W����tot�����x�7׶�/o�݋���s|�p�꧷�q���SO�p�7�H|U;ٜ�o�:���k�V���3��N��.2G���j��?N�AS��پ��^7��D�v�|����>��J�%��h�6���/*���W`����lVe=D8(<s�ˣ�/#.��w�;�nx#���89��͙�T�����d�ơ�>��{Y����8ff�]�6k\>��C����O.�S�
�We�&jD�#NJA�)/=.)��=v�l�3s�݋��}�%����hϤ��87�yJ����ǟ��r������o��MNܙ�ù{�Q|+)�Ҥt��&��^�O�
U�)�CkU4������/Ǫ��Or)N�� ��4t��ii�Tl�.X�ݣ�ˎ�oA���	s����T��}��ŏ�Z=~�+.��D�J���Z�ё.�pu�7��%�,9�;���xR󇒏x!�@���	���,���j:/\�=����UXi2���0�Wa$�,�ioSd�Nx {S�=�|#���ɇu�/�Ud����H��L�Q��Ou�3W.Py�L�8v�\��|2RޏOD�M�`WHv]��-w��R��(�|j��,�$%���T:��w�5�/c�#���M̨���6'.u�o7'T��1`�W@�ۮ���zX�zf�X��nW ���%������Ns1Oy͌��%�p�u�(�u�=���u1�0hЪ�^�=��je�����y�CWZ�9�R~��{�Q��W˃���Еgu:V����U�%O5q��ˆ	��	s�E�;�z��K�z;U��q�yu�FW�Oiۇ|��N{�~��>(E�I���8�x����o��`:!��AY}Aq��3!2�()|\��֓�V���\��J���Lry��\gy[�<�b�����z����Ǳܧ��rz����M-"-�=�/l�t/�;���vQ�@(\�F�H�+ٔ����e-<I�ȭOX`u7��_"y�M���`��O��8c�*�G������7�ymM�=#U���k�X�Eִ�o����y���Ô���wB���7۳�d9���X�	�K��j�
��X�C:�ؗ�ī��y��\�V2�Z:lr��q���Ԙ��U��.��)���7�)�X���iqT�G
��y�@9%�n�ضpU���Q^7o��DSv-WZ^�Ǚ`i{]N��ɮ�_d<[�ӝ&y�%���F�x���*���d�{K�.,
�ϻ�45��5mK}�K8  hΗ;[U������k�J��ܺ	�!����yWpJ�막Y�Z{#���4��RYW�i�ɝÛ�Ԫ�Ԭ�Tc;��5����RPr��aV7�h�YN9�"�:m�i����`7Ƨ1o�όj��HT��*[Gp�=�,I�<��BH�j�<6M^gM���E�L�Z��M����AT�ޜ���3
e;�Ex̸�pS+&�*��Ɯ�Ϣ\s�J�7���Vm�w'��4PU���GR�g7�=l�C��۔�i%w{����ZZ�pߵ�1W�R�|6=�zR���L���'�C�C��x�;w�rL��X�}�)@~^�s���1p_Vm�s��W����z���d��{Y����N�H.�e�}�*5G������*}�Ǳр�.嵏�ո���&B�|G�ϩv�՝s��k�Q���}&o�%=�ٯ(4��=�`������yPDO����7�z��Vǌ���������C\����Eˮ�dP����"�#�	o잩s\��K����[X�ey�AR�OJ���0��e��2.������:�s�ʴ9����ܴ��1��9�r�V�ۂ܎�fq\�����-6vn�ަ3�Zu�q�ΓkT�**v�\y��w;T�����֜��}�w�x�'��f�j| �n��a��"�s�e��E���1��pi�<q�c��M���9f�ͼ;全:��W�e+�Kj*�z���:���C)����{���;��y~3�,���А�x�.������c��S��Rϩ59��j�
�۸�+�=a�|eW�D?��41jX=���秫�9tofv��n���,�K��v4�G�މ�[�
��-
|���=F���Ю��{楬��<�.4=U8�dl������k�][��%�n��Z;>f��T^|��?Q:p��C�sP�l�T&*�wW���n�7w���nsg���*�E±��i������_E�Pe;�DS��_g��B?7���:�ڮ#R���}��/2�fQ%�Iw�#'�ԧ��0:�Ӝ3�n���ۗ�{؆��¡�ܦ�9�I�ǆCWtD�Z�**�T�)-�'2�)�ڲ�<�`��U��q����U�gҵ�Q���\
��t_ۉ���_��<nǾ�T+Gl������0C̺e��*�ؖ��3���ݼ4��ܮ]��J)C�7S�x9�������Ψ�]
T�l�MJ�Z`}b���g���Y���w^�m]l�Np��rG^&��e����4iJ�Np�״��E�/i�Rc]o�r�)�9���c�&t�׫���a�Ԥ�f��&�hn�A�>�k(<u�+�t0v]	n���%ny�A�n���3)�ۙi�`��Fa,�@ηZU���H}Mw_2n�'+z�6:�E��M
�6�U|*1��(�����3L�6Q�0�Sߎ*�(�q�'.U�-��&���4ϴ2.�.���:<�n�O}����#����ʎ���p�"���rV-d�t��w&W��F9�mIf�)�#n�o���
��2���k���$,�Z�/������tQ:��l�=�\�Bh���KL�xxݒ9�R����hpz�qj
�e]ؾ�z�����f����@|j��t��O>,�.P%&s.��,�:���NL�ak)�b��:�I=�V��n�+t�K	�8�<��oB��:��y�d�U:��ۖ���)tsې�w#�,�<䱛��wFY�^+!�j.j�ϻL�uU�؀2�t�	`�B���{b0����c����Q q��LӽA;�u� �%n��p5�M�se�rMQWaV6���e��i�k1�%�sy�r��1E�K��C��ַ�D�m�6Y[��d��}Ny�5(����ޥs涮��٘fh����ե�&S�Ar�[�U�VB	��J��wa$������i��pb���S��`u ��(�X�.KF�yO&Xg��f�$��6zVgU	hZ�T��B�F�L����s·4�45y�]��#��}zE�f����v!kx�V��k��eլ!�6��mF�ʈܗ!��x�.�z��P�T���ʬ�/!�}ע�8>��^��������D����'DN��z](�Ŧ��䭻�?�N��{�+���^Pq���=��Y^�F���vr�YùQe]0Ma �``���@�j�]�mo(�ufe����.gk~�z�*�s��]���_-ީF+=}@4\��_a�����wX��J�彂 5p��5��!G�w\gl�U�f�1]�[ci1�̾I�o�^�35qP�L�nU��	r���������h$3o�u����q1���\k�i�0vu���p�v:�B��h\�i�U�u�IO�(�
}�:�FR�������\���2�Q��#"r�pNv�=�z_+�-�[��hKmE�>��
�{r^<���f���|��U˥�zY��$�t.Vq��,�,�쨲��,�����H�ϸP�s�ք����v3��v!}�K6�S���97�-�+wJ<��A#��eoH��� 5��L�
��S�!�Wbޫ��Nk�L}T8�H �O���j5VԔaQJ�#j��chU@��-�m���J��eE*բ�eAK+F�6Ɩ�[Q*
"-�h������(��kUZ�UiF�K*%VѰQKBŃT�(ڕ���-�X�Th��[ZԬFQ(�Yam�h#m����2�h�DQ*�h�
ڕ-R֭+m������K(,�"�)mm�)h�b��m�U�-�KcR��Z�h*$��-��lX��m��kkiU��(�H�[mm�Э���Ke�J,+*6�R(ڵ����-b5���*�-�Fرj�ը"U�V�A�[JJR��6ŭm�Z�����[kXUeJ�k���J��V+�Z����-X+h�R�,���Z�5��T
�"���X�
�J�Fֶ)XT�+D[Uj%�)Z�m
�-J�h
K
؈��Dj�
��Z��N:��kZA��q}�%:~���.��]�V��V��,su�;y)�pڥ	�p*y���"�kzؖ^;���v�ޣ��c�t'9�d�����v���j��5��y���]F�>V)�J��D}�^&6�]/n�:ش���7�w�Y��G�ׂ����?y���x;o���G�=��	��*ҫ1^�"V��{=�:�L���6,����cW5׵�]���u�עm�px|�)tR��V�m�S���L�ή����
��
�_s'�Lo\OO�F`�QA����g�s<�ǳdF�%�4꽿<��X���O0=^ *���r��
ƦU3��-�ⱪG�i�zk!_3��.�*��w�*���7�b���ˌ������=�k�VΧ~�,5��b���{=����mW��8��G{��o��C���_�e�Ϭގ�q2�尫�ج�5��}7\U�9=Z������2w�����P:D��� �+Ք��ώwf��\��{ٳp�h��Ͷ�qޏ���eTȧ�z���w�P*��U���7�-c�h��_��NzX�F�Չ�]r����:ڃ^�K\4d�Y�)˘yLP!�z���X�ffw:'|�FPIYg�|w��4b���!�x��rۥ�O��Yd���/�U���S'�Y�������ó��YOJ$���g^T)̩
{P'��>��]��f˷x��4�^�t�IgZ�`�g�;
�Z���;��Ԯ[e�������g��	����]
�ht��6���;����oŞ�tpo1փ��W���xfnK�����;���FZ��]���������!���PͶ�.�`�LO���7�q+"�C�u�*}���4O����YuK�FD�R�\<)�`Iv��i�<O�!=�z�u�����^Ted�[ *�`y9啟t�~5=�~&3u(<�i3��E{�Փ255�I�c�"
ՏS��z��h׆���+"����#6�,w�9�k4�ݩ�4�ӎc5��`!���3)�C�=���M��x��B�e�!=���q��I�O��f3<���e{�h�0�R�3�E:>�c��fW����y�;���e���{~G:1�x)\�~��ں�u�-�RՀ�*���"U� 5kGE�ees�i�]�-���^�ӽ�7���m�LA��#����h{��!����''(+�!����fvn�3ҽӯdw�ʫ��9���}��r��oP��BŚ!a�/�*�5��!�Pp���ز`�l��_Ղ_��b�T�{Or��[kW���Ц���VZ��i�T��F{�+����J�7a�qL4p�s;8�"4kl"�Jd�AV��'��n����$T�1�� !.��D��wi"�?Cs`ڂ���q���s�����:�˴���V�1��bp3�n=T��~@��p�(F�	���{k��M��2}���I��lM�N� U<Չo���l��CD��N����]V��^:�v�n�w�5;6H"����/cr-Ńt�?^�bU?k�)ޕ������z����7����|���,�X�r�K�`!�n$'��Ҟ�[9�W�}�RVzϯ����Éft9�4�*��R���]	������e���>V�������_0pӻ��/����;�bR��.#9�P����\J��W�%x�ck#XoW�uy�����m%�=�>f�5�H-�F5D��1߈U�5}g��v���>M��)/�1�X��r�KޙD�ܐ؂á� ��>�`j��(@�(����W��wG�x]�7�����-R~�H�E������4�b��Ң����|&�۵n����q��_�S�]��V^�g�k⡗��y�*���+k��c�*��mo/o }�~��7��XL,ib�_m��_�jp&+�%e�(Wb9�;��nYh�r���{�����>�K�((��5�Y�z��!��lX���m��ejƗh|�����?B��3����ɶQc{��C:�ϗJ��,r}R�е+g2$����y�kz\Y��w�ˎY��߅V�|<'��pū�di
�,Ħ Qgs�OI1�ѫ�)�ć����Pa����/�ZG�>�X���x���Ǜ^��6ہvE�2׫#&��v�0<;6�G���g�vX�މլk)
X,!��y@�SC��]�u��Y�ݪy ���r�1��eu�X1�OOnE�R����[�z�� Wx�RCװnf����uyu*_Jg8�[��
��pe;������Á�m�a��H�<OnMW�焳�lgI/Ji
�l*�g���ϥ���5t*���^2�4U��9��W����y��C�	MƐd�#^.�z����lU�g��Ǿ�7�jWs�)��=̠	��.��Ժ$Gy������OUE���T�s�;��A����j�Է�=���;�O��8/T�xs�=Du�AmKY�=��q�r\�
�X>y۞/�ޥ݃e�NߔU��}�L�ã���.Ƚ�1�	�_KP���8��SCw�o�,�X�b�U�;�AwRE�G✅V(`�����וi]fS=����Se�h
���a�bK�c��+t"7j���2k�ڦ�Nb}��U�+��'1���X̷��j��$�r�A�9��]�*!*��Y���0�-)}N���.��JF��t�m*H��-��Ξ�|4u;���sOS���ʗPj�01ߊ#C��]��u��
���W��RfY��^U"�/f�<��י�2�*����B���Ie�]�W��3����)dؤ>��鉢rW *8d7*���U&K��X߫�"J��)QUR*t8	��[���O��0<�-���"r�pV��e�@r���cJ��-6&:�㜰��a,!J���]�ƖOz0���.ǔ�wu�8�;
{-�~P�y���U��حY�)�B�f3��@I٫���y�5��6�ɯ6�Ǆd�U�\:7g�*Ñ�kOe��綘V�GW��7��c���1Qĝ��{������#��%T�PVۿx뜸g��+Y��F��[�n�g21'�&}���uԠ���q/��W�1�u���f��&A��s��z�L��2I4ǝ�S^�cT���5��^�^�]p ��ʧ���3�F%�ckך�ݯ_h���=W���ϨHtn|�����'�r��yVo�ϔ@5�\d���+���X�(�#殕E^X�����	Xn�?��EΛ���k�=�tPWv�g�m��:�6����b�b΀mQ
L=f�@3U�K�vn�{�gb�	�:��7e������ݭ!5_^�.=�W�,G��6_��y�\��=KxB�tY)ۧ/X��c���p�T7˩$Ġ6S�毃�Wc.[%�Z�Y��m�����nߴVODGOj��Rs��@��yX��0F"�Sx0��;۞��R��n답ӽɲ�ӢU�~9U.(Ƹ|꧹�2)㞞\3��� �� Y��
Oպ�1߂�*��e.G�*i��f\n��2�F��n���{ ��z��o��S~��p��2N�{9�d��ON��0Sy������n�*n�FS�0��W����Ճy7����u!�Tשh��~VJ�dq'��W�4X��V\;x3u�|ތ�&{�I���.̼��Ǐϊ�T%=�+h&�i�W��^�8�>��]R�ю7 VX�%����gb����y�kK4�>��b��R`���j����jX���>zo.����`��١:%K���T�3���g��<��U���Ϸ�
U~�)	�����MJr�Җق�1���E�v4'�V��_f�Pg���eev��s����L���4�\4/�_��|�#�xS{)���G�#޵�c����du�B�{TK��=j�Mf!�=�PY%�����CSyLw�2��\IpŨ��s�U:���'�T֨ؽ�`sn��z��N�X��y|nѕѵ�&_S��o�R1�B����U͊!�c������g���b~KFxˋ�b^��pWS�n��o����������hx�d
�-/xv{�&�t�����1_��)�w4bO?���D����J֎�Kyʼ]`Y'���g��ѫ+xz�_xF7��nS� �;2��})s�]E���%y܄���Vs��E��ٜ�劊_xm�5>�b�M����q��۷�x(X�����Lgz�A���7N<�溰�/b�z��lxS&v�97�E\ �o����_d}���^(��p�(F�u�U��8���Kb<��v��G�f�#�q+�����D
�y�!�]s9S�����e�O��7D&�mf����28�%g �e�ږ��]�L\{�n߷�e��]�\GGD���UC��LQ�^)G6��Z�h�3W�ZCFL�%��M_';�:�-�v�d͞�l��;�n��F}ҩ;��m9d2�����>2��:�<J�b���\ٕ��C���b����O.��G5k��.
U/)S�7,��'~�|Ġ���X�g_�Ow�^nJrK��r/��޻� G�!��\�0�s���H��{�G�|�k���Q��9M�$�U*���9Ԯ�#!|W\k��2�Ygx�["�NE6�Z�ܦe���ȸ�Xܒ��R�y[@�6��.��k�^�vqe��X]FX�bs�3�{�j�4o����S�XlwQ��$�A���*_k�9���"pۊ�롘&{�~�W�	[�1��"����wc��}P��*�[�2� 5||F߬�f+�/n��v�i�����[�B��`��l�y�I��pZ5��tI~�J�����}BacNt�4�צ������x>��~���_!J��_�{��afł{oQ�
��J��錗^� 3��H�<s�$HD�L;w�(pd�GJK��މ���U�jꭾ
k^��q�/{b��^[7]OUtހ�Tݙ�vKl�>�'j�(z�
��aԣ9�à*Z���1���^��g��Uv�����oy��:�������.���������BL�ޱ����̝�Cc׀�������Z����X��{~���S}cFTb��|q��繩�D���t:�ppD��S�"Aθ2����p����A�R�X��A�R�.3�wh�.�LWb�]���׶YOӱg�U9�� �Z���*��2'�9`k��#X;Z]�g�.?Qse/N���FV�G~�N��hH@q/{n���/�\�l�CY�~Z�py�]����͗��2��p[�ԯ��LU���­��W���(�:-��l�Byo3M�$�����m+�}<��{�O��
�9y����w�R�:��
��Vҧ̜4��zb�ӭ��r^�ߨ@�S���72�.,�����2�zz���{��(�GV���I����m.[Ǵ��R��m`]��xpO!�;( CK�S[�{�����::�~Ƕf��b��:[��������70����\~��T'�WK2��������r���}���Uy�ac��Wt\8{�w���)N>pZYU.��i����zvfw�{=�k���
xUY�b��9U{7)�W��ʭٔIM���Rt2���V�����{'�c���G���&o�`Txd7>kG��Y�7w̒��
&��r��Yݍ<{�]	]�,�8�_��	\l>�C��},�V��O�~��̭\�~����8T܂�қUݙ��-�����B�(7��� ��S��o�98��:��V�pQ��]t�:���	����h��n��7�ᓯ|�2/
�}���tN_���O�a{Xn��rJ�a;�����sU޳�*�+=�	h�G������og)r�u��86�ݷ5{Z���i�CyN(̉����P���!�
�a��c]�W�pq�oc����kGlS��V���á�L�&�IvۆV���A=R9�:�z��'~n�՜��R�y-��
�.�����|=�02T�PV��Z7O��R�e{���BV��i~}�DWެ�����4�:��aϒ��W�1�2ߋ���^�]2d�{=Oe�Os���̱��/\�+�nRV��<�|`�x6=�UY�jxr�Pr�>Nc�}o���fk��	��MQe����a��1D_e�H^wO��>z���&�E�o:gh�J�{=O��Mc���s��]Hq&%��-�N��"�9t�n�3݄ly�;"'��w_
�}5��19��6��c����t�	L\���/�]�9]��g4<�T+�V���ݿ��P=���<C>��ɗ�s� �����4���~��K̋ +��j�YY��*�SNS��ײ�;���\�����A��~���I��/u4%i� _�Y�U��~c}Y���㶆�&��ȩ�R��֝"<gy�SW�,�;S����W^m)�J>p�����ٕYp���֌#�Ӕ��*�;t6���}Mm��-tw�a0\E�z�^��}��f,�z���֮Ğ ����VA��� �@;2����u+x(����xFd��#ut�J��&
J<���/TΜ�$X��1�Y�oRŪ�k`�_u�퍖$`d�yF�4'���]	�4�-U��Iz!�2"����yh*��\���'*�� �ڭ�lH���n���܀��H����*.���#y�,:���EVQ��Vm�$�k�3
� �������9�`�u��Xw[��z/�.�,���4٣|���)�������
�#�w5�g	>�k��i� �g[�|�5�r$2���R�8�v8ɔ"����K�6Zy����Dh�u%Mv����7��G^��>���T�%��\	��m��;�	�uLY�8T����[[��r���=Ɯ;���C���
�c���uf� 	��Q���+��dt�ܾ� &�gu�4_*�-Hi���([cm�&��ħwp��	�%�w_WK�٩fm�l$~NV�����:6����%�I�#���'i�P��g���cXsr,��R��6�I�L�ԯ��YW3�ʗȜ�ڡ���1lD�v}��f=�s����ă�m�T��ٓL܅.���ژw����/W\�+��+a��ưwm�����,S�@'�@K+`;M9R�Zf[��mN�|��!���fc��U��ȭ�8��R9������IK�.�5Ļ�I�_f���73�9weՍ���X����lS���h�w{��r��j��&ૂT@�=u{���Foj����)ɚx�����y�J�I����p\x���s��<���y}�w(���W�rװ�.�,ʰ3A̜�m���t���V'%�S���oj�k�V��)P9B�r,u6/u��#a:��_��<�әC�C��N�&==����ي��"˓�R�3`*b+z����5m��Tww�����k;H���K�R-�W�F��
���V�
nǇ�I�
d298��cwKν�z��<\G]�l�ɮ���y�}�0�}����B�R\����n��)��V����t:�k�e��e��h���w���F�[����E^U��n�q㮐=�:n����EM������tĻ6���Tl��f����3��w�SpT�uO�4�X!og(�����¯hR��v��7Z���O#+�Q��X�Veo1S��X*�6��]�of�e�t5��㢕,e�m[�:^�����R:6��&�V%�"����.�����Q�ԓãw���n���R*��Πޣ�lq�J��̱�WU���m՛r�Iv���:�FY��p��2u���5��+v���䣧��l�Ό2:�o��%�;�AX��^��|`�я:N9ǵNf����gF�\tm�W3� kt�kO�#�-t}�Z�[�qϲgᶰm
ʕ��Q+D��*�#h�QE5)mF�PZX#
��h5�eB�+��*��BգK-(�%@�TQ@�V��
�
�DF-JQeAkkR��(6���A�A�mTj�cK1eU������b���+�ҔA�("�k+[b2�J��ёF��֫*�j"��D���V4(���j����Z�Z֢�TF�eb�UjQkE�P�Z6"�҅����j�VЋm���X�KJ6��Ԫ��-E
��bԶ�*ZUB���V��E-�TѥmTK�*T�kJV�k"��V�)RT�U,+
�b�#UP�-J�X6�V(�AV����jF��Z�V,EJ2����m��lh#
��,�T�lb��*�AVQX�E��Ҷ�R�AcT,%�A�TQ`Z�J�ڌ���ֈ����-�h��`�R��h�Jʊ��2U`EL�!Y*A�	Zve��.CM�������6{�IKPޫ��s�^�u�a}��>k�c��+8�yhۯ7��nާ���l{��):��T��9Q{2���d��<&]I1X/Ń���)Sމ�o$�L�hy��ci�^-�6AlЁ�e���u_�GE��֙�)u�ݵ��.܋�yZ�W��W��y[lh;���q� �OK�/*�*=�&�]��Nk]9�~�l���Mx�}i�4�7\%�g�qU���;�2f������x�F��3����D���;l_��r��e���g��F�Y�J)�_�c8�fV���d��wݺ����}�Y�f������e��|����\�<�'�2�� +�}�k<I�2�X痳��훫�I&��phx��.*�e٪�n�P8�����]r;�#ծ����bt9��~&}�AK��eOS7&�zsS��P��۷�xh�ki�3�����3��}<��[9ٺ'K�W���D�U�w;����=POU߁#�����1�A^}���t+²Q"��M*�mq>f	@��b�]N�{��a���;((��|z����&���;�,WMyy�]d��G-0�|�>�f��-b�ݩ��8�k\�Yv�������)��ܱ�	�1�k���7�fa�������D�������(d���C��u>�������R�f�=~�i��%��Ă!�Q�9�q��ذȸ���>��¼��f�n���x�-^�S�l9t�u�Uǥ6}�֣@�3W�ZC�X�kg�}]v�޽���uh#KMP�}���zV�+�Q���siT��ts�接_>p����x���nh��s��ә�ӭݍ$�ϵyh�3�������<srɥ]�L<ϛ���Y�j��j��Z�vys%Wo�2��;>f�:= ��e �v��c]�B��.Z8��nș�)��oy��Fpl����}k^u��]n�ƀڝ�P��*�[�2��DF�����='�k�q*v�*ze��~�^4`��7=�Өҭب����QM̔2��u���ܶ��9��/= ��e�g\�J��jǴ�s*�᷊���g�>���80�b��W�s��}��z���֭Z�{��`CxUl��2�q0�6�3O�L�˙�1mE��5��.��d�̖���ҏ;�Wy�zEܤ[�����*5G��T�-1Ua@�]�n�9��ᠪ�%�x-�m����݇�KCJwݴ�y��ʉ�"=)W?�����e:��׮���:�T��j�k(Z��1�i.�p�aZNmi�ލ����B�K�\Fpټ��qQַ�d����Ɓ�Ɩ�k���6�=;�z&uN�w�/_<V�P�=�JZ��nfz�T�Q�Ϸ�c�>�r/z*�b�K�
�5��z�!�foV���=��4�-�����1�����*�q���U�C����g�8M��[��ϝ��Þ8O���uF�k0��/Ȉ+������p�����{�颩K��� ���.��J<���x?I-�SHV��|�ô��*��b�5�庚v��o-�F��Rw�����=�s��=�袴�^�<���	HE�u��F��c�o�=�r��D�o��zv4U��S�����ˡ���6���b"��cҳ1�|��f]K�ɱ���g���2�I����τ��j�B�����P��xz��_�cW;he�|N�9f��^�'�eq^��=��r�߄�w �(z�.٬�����ɯ�o[�W���}fq�>J����;X��J�	ÕWE�S8974Kt����k���95��"��N�BVB��Jg���+�Z��'ٞ�I|�
y
N���^�5���{I:�����c��P��E��z����Ns{T�A��}I@)�S<�o�{��L�,�Z{i�yz��O�K-Ћ7 d(E��ōֳ�F�<ʒ��ͨ�*:%\.V�y���|�k���2��f��Ǽ��#w�b��.���ޞ}�/:L�E��U����'�Z���ܦ�yɒ�^,�V�%^e����lqoM�>/ڻꬡ�*U������{Ѵ.��6}5�Z���Lz�s��QX�Vr����霙�5�>UoL ��� R��}],iٚ�{�͖6���+2�w[(�:�[]=�=��;��,�9�?U�����@�Oc�3麫t��/�g�5��N�J�ֽ����YZm<q��g����ڨUb�k�J+кT��3�����US�A[�Mh�>ߛ�f�oyl}S���5�&Ɠx_�.L��z��:����{�ᵓ��US=���?7~��Ny	؜OU�({&Lc�/ɳ�W~
��<�T�x �����w���ac�)���oҼ�%�k&�OK�X��BC�m�t�'�r��yf�LQ �\d�ꀩ�{�A/H=�i���DyL7����Mc݅�Gc��]Hq��P	L[�;3��:�에v<������^v�{����8!ns�P�����Cg�EB��[A��f藞x]9��m�����mo��b0��M��w�Zv )='�pN��G6�M���V��>[�ӽ�p]��i{6Z]�f+�� �������]sW�;��Y�s���dn�����{����8�͍6���δ��aHȾ黱؋m����ߟ���}*���F���r������<C>���T�����/{����%s����m6x	],�/�Llk�\5�<x�c�>��hʑ�P-�x��=�����0��W�y�D8{��Õ�LԢIi��q��Ӑ<�}~S'ݫƺ�:���Z}��ت؆Z�X;����Ǘ�J��$�¬�=�P���	YO������:�5���3�X�����K"��r木��S��`�E����V|�{��29��:gkks'K�aB��y�
�2�d � _t�<��,��ub��Vr�3o7�=F��0�g�s�8;R��ES�Y�}+�������]��7�=�u�Ś��ڮSfi��G�^�z��ze�������f�
/2��E�Wj��8�	�L������JR��v���gi��=Yˁ��ȃ���.�*��Lo�,`���n�]�̭x��ԂSY�.P��\�я�����[c�zl�W�1٦)���;��"��FׯD U�˙���%};mz��4˳��:�J�lm �|�U�,���Ǣ�CI�1�22��1p�^_�j΂�=�J{u0�]IcrR��u��8<!��=��ghcN}��җ�,�#v����9{������&B&�:�73�%�#�>C8����Pr�q�G��]��vZ�dzi)�>����C���j�v0A���T����0�o�����;��d{y�ɐ%>����
r�݌_�6�k�8���@�C�A�R�e�*����1u殱;��U�]C�Uc�J����>��ER*�;��z��_d}���7e1�w�.����'Mx��/� 0WBEFRiWe[\O��{���@�y�!!�e�N�B�2���Yk�w#����v8N�Te�E! �v(Д���F�Wb��7TeNB�>]���Y�æ�o�5����=L�y�F��5x���X��!�n�oN�l]O^C]<�w���}Q6�����+�F�J�}�)ͥRw���,�M��a�@�U�r��_b�v��6�W�����>�c�����f,�;;C�\�^R�畓[�Al�r�4Zn=v�Y����;9�^��� �x��4<n�w�*�����m3�@oHA�Q$*w�z��w!$Ґ^�#����6.q�#zy�oÃ���}x����Q*��Cc*RzGK����f�`K@y;"�h&^<�(��EoGg;wLǻQ��^ԱX����I��S�j%�-d�t�f�8�YB,8����+;� X��H��h]kw�(),S�҆��A�;�4�C����	]�1���C���sn���pj�S9sa�E[��9�H{d
���f)�츳k\O2��>%��a�o�@�:��tR��
~Ñ�^s�\�����`͍�Y���8�x��<���k�ݏ����,��U!�'WH���UuTl�]�~�۽~P基=V��螪�L*͵8d��^N-�ܖ�zof��L��"kò4�y���ٝ���W�\Xz[�Q�XVEPt��ɩڭ<���v8�	�8�0�r/���{����C�=�}�pȫފ����Ǖ*��3�uˍ�b���9��ju	�B���R�����1�0��늼1Ʀ�߲(K~�OvB��pǝ�S|0�7[�����%Ve�{�@�9�2ߏ��37o'����=7�4�^��i�犇�5{���/�=�)�"[
�r�-��;�M�}�s}�c٭,�B|7L�'ᢲ�w��Ϝ̸p�!��v���;������#�3�{3���n���oz�W9߼X���u�ʦ�� gs�	�բw���U%�q���P�z���P���pei�۬�7,(hb��_�t�Q�*]�-r�{ٕK��İFe��XcJ�mI5�-�X�7�Kpi��盄����N��0���^�5f��EĎ���k�ha�}���<���Ҿ��V���%��{�]��([�y��Rs�$W�������a��jusW�5W|��Lu���Zd�3��f/tw��"R�/1���>qb�9��p�3}y���j��@�]n���yCss�p^����P�L��v��C&�{gc���X�7{,��b�Y�y���;�B��?D�]�M��[��]Ւ���&�Wb=��-�w˯�潌fP����3�,|��'�}B�7J�@�t��������t(��s�J��11��9�S�c��z�xo�҅�H��J��S~�Pz�!�yB�xVGݘ��y[|�X�yƓ�V�#�����sj��l򃙺^׷ۈbN&��G��ܭ��'����[��u��h�Y�0�����5�{&��s�f�L�Ḵ
x�W��B���J�^❵Bv���Q�f̮��l��CM;^���!�7]u�]�- f�9�"*Y*S.|�U�YۙB핸��6;�n��	]�#�r5Ms��b�����uWItF���l�[,օ��,�Ð��Ü��6�,� ��\ud�m'���.dɧ���IC��cVs�Jw��y�Y�o��x0�Q�.��z�U���W�:��L��o=�l�J�Cޏ)�=�4?nS�t�-�Q������F?o�.�s�q��xX����M�M��MݟN�7��0��ͧ*;�#���s�g��Y�>�~��'O=�y�j��ʧ٨�,��q�RXw���׫��+�ev��\g�3�qo��}�{��Rbɚ��SWS"�e���SU�~և}��w%�'?�Vu�]�/^]|7g\f�a����A?or�̔�r^��^�K�yM|�]t.�޵or�\={�o%�����u7ڳ��K���ʮquK��/*&p��4Y{-}on�{�����f��𾰦�=^�vG�����S6�H�rl*�B���χ5��P�+���"��7��V��fr^���"t�@�t��9�e3�~�4��k�z	����hv���/���\�|�ը2�{;��'�"���{qo��I�`�ܱm'�)�B��wGZ���l��e=��j�ۺ\Obt&� ���ٽv�Z��hX��iN�V��<n*R\"����K�����{ǒ�>�7˥\�K�{�ݚo:X�&=]+��l����ڂG ݕ7��w#)��Qy~��ϵg��%�[Q�k���ϴ�tM#l���⌯\͗�uO*�|7�(7��Ld�U���ej΢��1��m��>ٵ�hG���rٸ�{�׵^]������H���sv�+��{*�gQ�5�u��k���ru+�Ϻάf��}S\��w>�~�Zo�_횡^f=���Վ�tLoҺt�7y���E܏����Fk9ڹqJy����-�w�9����'���_?mΘ��4OnT�����ޫVm�s8J�~x���xu]��\�_�y�Cy�{M�ki���۫h��S��pO���Ʀ������� �z�[�w��<��zp��vb�LB!��V%ܵWF�<�}�H9�|e� �k�:Ϳ��}�����IO��$�	'� IKH@��B��@�$��H@��$�	'��IO��$ I?�H@��B�]�$ I1H@�X��$��$�	'��$ I?�	!I� IO�H@�`$�	'�$�	'��PVI��l��wAM���@���y�d���[��8 �        �        
   �T�"z�Rmm[K���k����&�6K�NlM�٪�Ɔ��j[EH�-֫����Nۧ�Ñmk5Z[M�-��"md�V�jԶ�ih�5�mj��EmB�Xm�1���e��ݓj�c� }�m�Юz�������7���뫳��y�����=�(6Ŧ�3{��V+jڞ�f�z��1ݷ�n�o2��m�+< m��e��=��Z��J��;۔��Z�zq.n�ݽ��b���ګۛ�U֦�u�*�gY��GwQ���m���-I��� ��@  ŀ    {��    {��    �,��p��b���T�ۻ�ʵ���k�j����w{ٽծu�ޮ����[+16d� �ot�^탭����ۻn�j==�^�z�l鱞����Mݩ�eN�;w=��cRT5��S���ζmgp�6�[f�� �n�5ۻU�����P�n�ݸ�F*�n��v�lv����nǀ ��z[+m@�p
;��b V��ۮ��n΢G:�:�����b�M�����x � 3,U�D�^���Q����AU���Wvpt�f͚k��SZ�mg� m�J���&� α]�3cl)ۮ�
P����� �ց��;i�m�kK5�< oZF�6��=wݷ(SV+ Z�6� ��wp��L�v4�  '��iUM�E]���]Xu�5�gw .���P����ح�7s�>@@   Sm*����M A��� �{C
R��� h     O��J0     	�B)�A�T�?Tb`��0�#L$M	�0�SF�P��MG�z����F�A&�!��SP�ɉ�i�0d2����v����ki{v떵Tҙ��Ʒ�Y�l��b����K��uH�ޏ�׋�!!�jK �	$�;""#/ޟ5Z����a"����W�+�~��F�4n)"�QQ#�D*,������n���A�QPeD������v02)�v���z�{�l�I�U�K�{����Q�e�d�축=�Sn���ܱe���ˆ5��x��t�Vƕ� �<���;��M�J��s�`gvD�l6�@IbK]H*A��нP<p�s�H�Όs��rMZ����<(���xNpx���7{�r)G��v@��ࢁ������J�Y|��ݢM2���LID�MRń��:�w+�v:�\�s]�6nK� ���3n��F<�P��|z��k���po�vI�޽�*�Y6�Y�t,�qN�KN��Ƣ�v�8Ǳ��_|$e�Wr$����r���w���] K����б�g��Ӿ6��y^��RjT�`	�h��u�Ma��&���l��=���`KD�"i'*ܚP)$
��o�FZ����T��ٵ1�b.�FÝ��RDf�Y���{yj+(��d3@{tS�ٗ�k�wL�Z��\}�BC�q��{v�	, �$��eծ^�!���ìok�AF�	x�Y̎�1�
���1� �]���S���#7o%�D��i�t�b�����7"�hf1;x=����uN�_5��9ɶ�6-���n]QD�n�כ-�9]�P�-����]��Pr�0�ފ��>��9ӊ�����RY�*��]Qw-�:��:���ަYt��x�	=��#�Y���]�ٲ�lVH�ơ�eg�Rٲ�Ƚ�d������2-�`M�˽D_,닭��q�������C��xgR:nܘF�2�%\ڭD	L����TrF���:V�6�y��xַ�ڄC�Ȉ^)�q(�ߋI�qj���n���z�{_p�4��%��q%�r��'x;�7L}бݣP�c<�r;�G
���}Ǒ8~9 �u�(��+sƸ戭}���<=��6��������p��4�����~��4�j}h)U�����V8��Ùub���,_Kn��jFo����Q��>��>f��& ��@z�Oû{n���yCa:u���'"�Dκn���Β�/VrBYlk���zV�����#J��\�-���l�;�9ő�ƯaV8��;��V���/@��a�7R���Ү�ѳ7w:����jĪU����.7����7i=��#8�l�\�@�D[ƾ�Hٮ=�ܹ����s^@]zhe�wn��ʻ`p�Y:��잻OwLOF�6AӃHr��Q�N�\x�:~�CRo'�mط�����oSoU��	����a����b��1-��sߤi�����޵��Jw��kqi�9�Vi�V�&o]5d"���X��z��1������f7؀M\x7S�v����3�5���̮v�S7���Gg;�Y\4��V6e�8R�ۇ��e���������v����~hV�������;�tH����9��n�\G �O~�}T�S �Ӹ�F��{�)��=l�w��_����֠W.&�Z��C�����@���-��Zc�8p�|�L���/7z��ӊ�4s�ON�F��-٨S�:�z�g  G�F
�����{L���7vۣ9��mAW��u��76gW��K�4��db�������زU2婰�l��M��^�8�{]b�¨h�k����;���[���W��>nw�x�Y�m#��c����񣲵�dCK}��l^Y�0.K|@�-]�	��c��#�ݻB��Gn��n�u�G|FN��E����AP�{�w���p��XS�����4�T���^;��#��f�vc�ƥ��w{���.��uc���Og-�,g�3n�r=>6Y����[6�2>| �Eœ`I`[τ�s��kW��6�g�ܶ�\��O���zP�J={A+c��\*^O��='�mhz��߮@;f�9~{��Z�~Ov��,*�Y��{#�eY���v�n��	����ų\�Q���˺]�E�e]ڲ�=�SuQ�v!97�6�o�� ���w[0����w>�0�u�ev��}١���Tec�@��S'�a*7���=\^g2��;�t�MDJ�o �Tg-���4�f�;�9RA�l��&l/R��`��'n�:�)KG}N��V3�W(uL�@�_���u�R��̪�U�J�w擷; �X����'+�<�����b�ij�5�R\�[���dt2�	�E�i=�%��Q�u;��wGp.��˷� �V�4���ktwE�u��iX�tؒ��S�Րl�{b�ܴ���
�͘D{�ߒI���8���θ9�1�j�S(����l���l���!Ӽ�8�3Gk{�Y�����4�
�3�$���ҰV��������>a���Ϙ��Y�gaA�ըam�='2,O�eM�`-�ģe`n��i�������ѣGvi�1J�gsRǬ���zbs�wZ�3]�W J<�=x��t�c��w�#B�z�p|h���p�Q��wqoY�f��b�J�\
ZNɚj�����v�9�k�`Z8-(=GO�~��Wv�7�쯢�u@���$r�uR;Sd����b�q�����B�x���%�}�3�3� �ßtet�Zx�����!���E�4[��7{HW��(�Z�;�`�lNY�.��9�kGy1{`� ͛���o�PB�1�)-��_�j��RH5C���rR<��D�F�|����`k!��z�/:�e�>lUػ�<5�b�RF�e58��6����R��\K: ��ݶW�U�Me��{;R&9�7q��-(�����𙼐�;z���#
ޒ��oY�Fv=){�N�]�����dOS���(�M�r�<8���vnH��7�p���P�k�e�ӱ�Q��f�j�H��h�x_��UĢv�l�:Ϊx�!I�o[WO�^JyK�xҴڬq����
e��B�v�n�{�X�Kk�2w2�z�-="Q�a��x��p�I8(k�o9�KGn�ڦB����m!�̛���\��j���=���dv�ˇ�I8u��Z�qD�+��Fǃ:�JA��k9�q�\��Zb���Z�F�xt^���e��:%c|�J�V�Ż�
�w%�z�e���h�v��9����7����>ŕ�ٴ��y�r4h�P޺s�௹�4��nO�Z��b�,�0�m�qҚ�$&��\���p�l;%j!�����k]��hZqM�0&��{����ZH��6ܽ��rl�;Z�(��c��~�r\�:GJ&}i�Zw^v�w^��r]��9�cԆ�D��R�_F�t���S}����}^�ܣ1��ANb�>���X)hn��C�蛣)��+9h�\Nb����ÕS�U����tժ�:�s���=\��ܷO�՛G4���CGB+�c�t���&�X��z仦a��(z诱i��N<��4ܥ�M䍐�QbB�9&�V��z"�]���n����
�n6/i4���T�m�r����w����7�������^N������e ��w`r黛r���Nd[�{�w���.JvP��s-]��W�N n��C�Nr�ƷR��f���w/����Tjn�oO�؋\�X����r7Ft���e(I�#2��Dw�2�zGڱr���4i�vm�F�!f�s�h.�qc�'=<�j����)Hؘ�ד��A0,��c/�����
�F������}�z�'w�+��a�-�t�9�p}1��U���u��Y�r����܃����;:��cX��Ґ=�š�Ed���]]�Z�͌[���AѲ~?h{����%*�.o��U���.7sk�Z�ݫ�iױ�<i�`#�=u�Ō�9h�Ww��Z���1p�3G�����.FF-75��9�	�'s(<}@�Bm�"�>;���8�3�z�����Ol#.#aV_��w-�&���r��xޏ��u��n��y[�{��K�wI5�'5E�HU�Ǿ�K�v��p���p2l���Q<H�>Cf(�oUк�UE��R�s�?����k����ɝ}��nX��j|4�I@T�X��nF����)#�;{S����[b�[�#�yW�-S��f[+�-o,�)*^vѵ�}�mR�4����/gWW,�f����0�ܻ��d���coef��L*����x���j�BR��G���6N�N��kc<.�-������k�i��ڭ���:�
�|�RE��:΃m�OrԺ=��Zm�iʆ�U��
�|����2y�:�\��@��w(0g(Z� �mHU
�/n�,�kV�6��=ro�a:�Z�[`��6ӝxl�ɲh�B�����>�L�6y���\~s ��C�jTi���ڏw�q��},p"������F�:ך�%��vՌwY�7<wFE�A���s�����՛��-�6a�Sh�O^mfWq���
2�ח�ً.�R��.���]GP]Y�g=�XL�F�������P;WM�/֒9��Gy��ה�ִX�=iy�d��̚�3��T��|y)1-ֶ���-�+�c��/x���`.te��d�`Wd��p��-��R� ��Hδ��v��iȜ|�7�.�4�`T��|�j2�fi�g>��]E��b��v5��u�yT��9�ʒÛ0�/��P}̔�j��v>�7][�m�8uh؆�*�&jp;�,�ؗ8 ��>����/L��W`���5���P;޻o��I!h��t����-KQnOg��P}��0�*�p����/F�{�]�s�uΗ:�W10}��@�޴���N"v9�����
�8��Ҧ�Z�y�� �e7���#�.����6�mL��F�؜�c��
j��8�f���c=�񼖳���v�_ͱ�>Z�l�;.���==���5LFӁ{���52�/��d�6��Eǎ���0b�\��j�!���o"��t%��s��Jx��5m�=���\�ě^�R���q����z/�7����7xZ3us �NE�/Q�U�htY��r�l�g0��ڪJ��w_G*R���������c5��2�� �+���z������y���ۗЧ�UM54]�2\�ᱶ�š�d���F��R�Q�b�u��&���]�k�󰌘�N�>y�����:*ެ� �a)�N��hdw=�/?{N�xy7�>��l�f�S�.�)�����.~�Ս�#��8�ĕ��9=�Lh����ߙV�RO��p�~I��+^�m\���TX��A!gMl:�7���R��T�,覦�Z�|:�8.>%v�f�7u��,*�卝�i�@�u�Z��@��U�@i���J].huӋ֒��T�nSZ*=��sc���ύ�ɰ�2�=�wN���
.T.O$��h/<�'	}��p�yd���R����x�dtU��������:�k_ќ�-Mue�F����dh��4���N���<6�[��2��0���ܼ�`Q���^�}Wf��ۣ^T�9��6XX��Ɉ��`�a�9k��b
^b��VR-Ǖvb�Їyi��*�Y{�	Α=}�1���v��E�mR��@qj�seg�^x}�,H��ŕ�.{���`�6{��ڏ[]�['q�SJl^�oW������T7�ZqU����>u�	��oei�Yж#�I�r�Ws+77H��X�	�']������yg��yꗏ\�(�=X��V�M��/{p���nTՎS64�wQ�y�l�7������ְ�JEW:����P���q�Q@��:�[��7C�;��?c�^��{@�7��ug�� ��v!�p1);�+L7g$�v(�u��"��I�{�[TJ��H�̲�kq��"��k����&����_2�΢��q�=�p�.�i�́�*-d�YiM�̋�b�2�S�2̣ �+)SYݗ[p+���hS��M�au�P�^8�ۻ��nLR��"S��'��p��e˭�)���I(R�pرR�P�8mW;�m��U�������a�f����7a0�f���D$�7u�ї�;XG�>t��R��ޭ���Ƿ����+μ���dyyE��S�{�k��_��~�)o�n���U�{e6v�;��9}Z-5�g0
6֌0��b|e��WS��:�R�ӽ�Zɾ��dg�|Ǯԓ%���#�Q#�f�'_\��eQ|�6tB����F��L����$�6oZv]���+#&r)ޜ\؃;X��<�F���
�^�e�Jd]u�27/�r��Z�{XP��ԭa�S��e��|���D����.u���N-����<�����n�!�p�@�DC��j����,�P���<~	����=�4c����G5��$f�P���kܼJ!,����V4�7q�J���[7ձ�����x�x�V�3"����WmiK�*�*�$X�]J��[�Ƨׅ;ڊ�d�N��,k��HMpU�x����eK}���/f�|�[|��K�`��Af��u�j���y[x���h��%|��yv�m)��߆�.�, ��͎�;�Zva�'�muEDl�zeL5fT$��>έn�;{�U"��g$�HJ����k��0.�D���.�u![�#�Ю�m��5�ģʻk�s/E�~Zo���Nv,�>O���Z	�]��ᷣ�5�ݑGk�W}��{n�÷O�8��f�D�e��pU�)@^��e�*��{��/������DT�f·1��)Y|3b��^�wQ��Q��<Z/�{���+d6H�X�����wQ�أ4=Q�{%so�셼�1�Oc-��Y	n79��Ӷ��qr�����?e�A�X�Y��~Q�ܨ�ä�d�N�$�����R��q۩%����ڹE1m�v�ä�k؎Ь��%���'�SV��M泡ze�l�\snT��;�y�������:�i_$0�o��&�쥐W
>k�9�iP��<�OR�C��W��[{����y�CCRe��7Q��j�j�7bE,Y�9*Qwm���ֆY��1[��g w1�oB1�㶬8�)dT�b*�q��s��ht��󒹦x�.��ڝQ����V5�Ž&����C�Z|-U�B��I�/۲����[4�����af��Ӵ0��;���+Wqzotm�}/6�;a����j~�[�7�ш�!�߆��_���sU�}̤��Dq���NX�	I�g�Y��1��W84�����BLǖM��r;�Vl��,��ڭ��ޢW���R��� ���5wt���X���}�X�,�7>19)��n-��-;cUp��L�(���`��J�����P��<�wx�S��+[Z�8a��HL���^��:`��Fyc�MAr��.>��E�2�����r�5\�1M�5]Zw1�V�x1�}|C(
4^o8�Z�XP�_N�׷6K���g#)�ԻFP��
�_��mǡ�
9�V!�'rr�k{CGn�%Vj��}~��o{ �^�Y�:�r����W=�m�6 �&���]����yk�}N��C/�R;��Rb'���'�pf�O֮�N�<�ܗ@�[�)V��wpZs#��%(�3#օu$�9a���w=p����%�`�7 hڃM�A"'��*����j%Ba��ӨN���5�N��,u,��S����>���$,�p^D/`@-�^��Wez�ݡi�K��r��642�=���N�`���� ��[��/.��wL�0��wj��em�q$�q]��عy�z'�x�y�[�e��w_V���H�=�]�i�1�uO�V}�kޫ��`R��"<îJG�k�+b�ܫڼh�Fu��p�u��f�u��=�Я{��V�1�����7�YZpl�.Zt��Cb�:,�j"�"0�o{L�T�c��,-O[ƨ�)���{nSە��c%��6�sF���ȕ�;�P��;ɕ��q���|����;ϯ�zͽB�u���=t�yc�7�I�b(ܐ�����KiH�|�X�L���lGv�c����iY"ηУȜ4�=g��R���a�z8��oN32FB���rH�*I$��$�G�F�m��m��m��m��m��m��He'8gnEnvl�M�����r(u�I$�G$�G�G�6�m��m��m��m��m��m�$�I$�I$���E#�I%AsnR�iB�L�N��$2րy
�9x&�x��*+G�m�@m��A�ʶ��b��j�5����jD'S��t=��`��H�V=��J�2=�pv�D��@�4�T_*0����O:�ض�����}�-���8 �}O�RV�q6�\�%"�����O�+��J�C��/���8T��$$"��ۉ�!�=�Iԍ�8)j�H�$"�j��Z��T���,mz����-�n�c��f;x��i�C9��j�C��6�b5��U,u���iw��7Z�دr|�xy�����L{��g�儡�dL�����(������V��GaW2��e�y��z-���gf"����i�Q ]p�zK����wŋ�Y�vs.�w;Ń�����2p�ї.��j<
2�Y�I����s�w^�{�A�<p{꼸��+x�ԝq���[���o�)Y��eQ)��7�����Lԡi챏f���</�z��]7,3���u�`���PU��޽�Y�jI�k���yjE�^^єE��a�&�4wV�v���x�;[�Qu�z��`,�VS�um��=��8��9סP�0r����O����d�)
������H���"�;����JNs+�]����]�_,O���^��m�g�	@�ɠq��ۙ:hteG�nVb!�oy�r�m�Hz�w5�n���x_)���o;��m�8i
���F��c<�����p��4�-Y&9�n��G���߄Y&7���]�3�k�p�}���f���
��'df1��g�J܋\	i{�C%A��o�e枣��A��Oo
O]}�w�հ�ۧ��%κF�Ji�0|s)��]ќ��#;�΋��lʽ�*urպu2�͖7HX2���t�ĩ��
V3�M{4m{Cʷ5��G<�d��>�[�����+N͜���;D�jM��ԫ��\b�7y1�1i
��i��'�t-.0=���0�=/��+�X��P��z��yr"�6�֌X�m)�9�)��2D]0~�4VӤ�}&M�Q�������&)ڴNGa��w?zQ�7�ɬ�:ý�E���@��Z�����~�هe�&���w �:¶���3�����/^V,I���ڻ�\w��i\��/�\��S>��~;FƟ��f��f�u�b���t�Zu�ԯWi+`wԘ��gr;<�r�[��I��ujq��:�Y�+gv�jE��I�Gr��6�\�L}�qS��f�_b�w�.�
��A���Np��(��77��-�u�����(�H��3�R�a���I]9 �rv�]7|"�ќ�1N��8c;X%,�z��{1$2��yiZnЭ��js�v�;��ͪ\�����k��"�Mެ�%lp݂�L Y��T���ɒ�����nj���MVq�3���/x2˅+��d=�Q�r�f����=@ݛ��L�Po �R:���h.���_*�d��V'm�s!_gh��<���f�>�F�cF�h��uL���k��h�o����-ұq'\�ЏU�cA'9;�{b ۳�S':B��b�T8�Q��7��]υ"�[-�m��\�FڶqZ���%�>�jۭ��j�en�P����oa2��!�0�;�v|�D����,r婳Y�N��� ���8u��V2��j,��pB"�2�h���m�3��.i�)�Î+�wt���	�.�};��b� ���EN��!q&�7��{�ݞɱ�'��>7Z[\
�R)�Ӝ(Y�J�1Km�l�l�L�w2E۫R�в��v��k3����s]s��kX&��*<*X���R�O����<+�
��ű�Yդ�U.�u++m���.�=�ɗJ���� ~��`���M��f �{K>���Bv�}��u4�5\�}v�j�s�x��6�Hm���[�`SCs7�NM�Y���:ۀ��z�-���Xj��;�]l&^"�M����i7BL�W
�N�]Ъ�S���h��k�x�`�{�*z�\ᣆp�N�^N�J���Wq��!%�����_v��nKMwG�Z�hP�q�r�H�j=� ��C�7�����m�F�a��w3s���Zf��<�;��V OmY�؞)4E���ʴҹkL,��s�^jU����sᖮS=q���G؄N򷕎`ߓ�x�p�eĸK�a��N��wF��x9�=�r���㔤Nn?B{��&rڸ"8_? �޺n*~<^ۏ�`O3~Z�kK8��*;���jA�֬�:�Lu|		*ެ�:�hm�x�3�1||W�a����&g#�8�2�:��d�:���#2�Zyʹ� �Is5Cj�֮����4t��rji����3���uǥ��%N��f�|>�����3֋�s��.�E2��-�sox:��
-p�ԗK�<F�AS�s�o��G��1����`W����C�7���s�/+��GI����~ye�QZ�u:�h�r��5��}���0�0�vÙIʼ;w�"p���MG)�̷����]��趀=N�^��
�S�!�3GW������5"��3��)xc���>V��p�u�֐��6mZw���j�0�q��ݪ��&�=f���h���%�=}��Y9�����,p��eq�'C�R�C0w
�J��Q��B���}w$WX:�-!1"��ft��]��O���ʜ��M����M�V괹�&z�,�v�0�d�.���]��wk��ۦ+��<\U��_0�Y.3�<�{Mk���M���q��Xw�-b��6�P8�ӿt�*�Ok�F�Y�2ݦ�s��N��]����J+����Y[�c�:��}7��e˺��1 ��tL��w���A{��7d������qr-7*+ӻdS� �wk�o(Ė�: ���g�ܙ�-Ȓ#��?������{s�;v�]�Y;{���y-�-�yn�Kŕ�*ڛ�Ǚ$����������X6�c��r]��qn[�A]:V���V�*�� ~�m#4ݵ��z����0߽9���C6�/���\���۾e�ɛ�`g<�gE�(�p���|�p r����dы�{4v��D���*�����]PẤ�!�پv�jͤ��{7x)��{���ğ}�@���#�b�k��ip6F+���z��f�{	�=3fM��NK�����[%Zˬ�E��Oe�nt��4�X�����jo�r��h�nv�86	ch�ŷjѽ�Y� -j&̭�V���w)�iϝ=�5�d7�]M�%�Am�:���131,u��,ڇK:L���֯g8e�7LЁ[Ul��5�͔�o�o���%�>���p�p�uY}���C�d,���H����x���6��N(�OJ/|u�jkˑ�ӽԤ2����']J��D6��	G�z?{#��s�qR7i�K��e���[�y��4ta;ǲ���|�'�B�<���[� A��r��^���xzb�����lį7��(��἗�	q�ufoi�p(�(:�@�4%'�HG2ݝܫ=(;���b�@+KP�N�W��{�kc�r�&��8it�^>�HjD:�'�U��O�5�C��\]��zQ�o�n��59&p��zd�&9��9���D����g&�w����ܬ́Z��"/���,�u�dߞ��5{x��Φ�v�Q�Ǯk�Twe����؉tX��VP�L}��^�S1Aٱ�8�Ȗ��"�7K��^�r��D����t�2����hX�\�v�0�nv�2��Jj�-Ȁ�"��~�W�@�f���fݧ���|�-�&K��´!9�ݯoxT�zuEy��Op�+Qm� v�� s�Ml�{��[�^���B|�ݻ���]�(�c�Ү�o�s�]B1��]uXy��z񭙴�n�<�EX����r�׈nav�,m~وh��|M�<���O2��~�9��P{��%&݌%�
���WGi��k��@�	��Ǫ�=�;XV+���Z���>�tv��uMg4h���֦N�ñ�ұ٪�w[���d�M' ��S0�onB��.�y�I}|Xȅ�xf����&���.�^�V��J)2�=���v�y��rX1uDY��Ι4�\_oh��mU �b���'�:����,_/]g�-�ۍ�+�_0�;S���bVY,���a�<e��^�iX>z��}<U*�M��K�7�p�Y�ag��ݺ2^�ؽ}DZsjZh����6�˦��c�F���$j�{��g]�m]p�k$�GK�A3
�2������3d��I���+�KP�Eu3s�I�L&%PW���L7Z����)*}��6�+״F�V�X�g�.f9�����S�y�}�S�W=╯���I�؍�v���I�wf�����I��5œ��h3�o+�9���^{���M��J B���	�`����J0�5���'�-L�w��7���ժ²e�TEG4�uD�򆊒�n��o�L�I�/5
��ǉ�^�ەas��4�����p��Z�ED�p�l�J���@�[_e��d�b��^�צ�5��\�]ꮬ�z�6Q�J�>Vq��ș�����L���!���{��x�{;r>���]�\2�m�;�H�v��9�T����&�ͺJ��Қ����Z]�/`ec\�T��E��͈=�͝ℕ�U���[S"Y��=�3U_Sg�b�����w|�%�;��åw���l��x��<�)F7�K_<�w|]Dڢ�v��y�Kf��i.թ��"�u]��v��t��\f�ޣ����5�VN�2v��`�N;�,�gK���M=�����S�p�9$�H�HbO%�U��L�͢�J𻿎���bbKJ
���+�cp̕X��Q����+�0�n��c4�Q1
�1bϒV)�h��E��efGƉr��j�E�b���+-�j�J��h�q��Qb&�����
�o�Tb
bQ��DA�wq�"7��k�DE�d��D-���"��6
��PTQ<n�b��]��F�ATQ�U�A���1��ۧV�X�X�QE*m��JZͲ�2��5*VQJ�$F�Z���3M��*�Z�*8�� �*H�i2����H}��foxd6W�^�8����䴃��h^cO#�D�2�L��7�rW|Rﾫww��������PyH��#��C�3`�ѳ\>�W��Ɍ���Ş�3��F��aZ}e�����.z�gS�����/ۗG(n_k�f�o���~�QձAx�h�Coد��8p�tJ6W�=����L�5b��|q�Z�TN%|m�>��V�Y�$�xo�������*)A���v�TA��o;�eD��ߏp�����z�^����<|j�S�Eٓb^�O�	F��x�zD��˯x5Cΰk)��S\^ݹ��d�SA�ឪ����-��te!�'�^��R �x������{E̨%��MM_S�Y�ye�g{w�>���K�zl�Z�IvF�	(w���a��T4{�\*A_�_�����S=�1Z��Ú�F ���b^]��*k�)�Mq{yx�+{݀��l����9ӰcpԬ�CS��r�Yu�ml%�s�����g�/�����)�b�|�m�w]����^q����?^(t�����O`��u���Kw�^~��Z��i���y��p���y8H��?`?Z#n�:2�<@�dg�K�L�(�bN';����a����	���{���t��+�OiDuy'�/��]to+%/��x5>��u�c>^��������<��sǩ�ߗi�{�v>�p�|����}H�w5��c���S��f�{�j�Y�K�uQ�κ@?���{Ĥg��;���Я/��t�M���y�B���}gsٰ}��C�p6<�UR��s�41Ֆ�J��t'� �����*Q�1��B]v̗����R�º��a��IEY\(.����hj��wM�n��\I��Ś�>�z�_�մ6���J��p��ݸI�N��ξ���D��r�9���;0t-�<�sOu_��x}���`��~`���Dㄧ-�wk��ܣ��zķwq�]$>64V��M?p�طS���I�ćՅ�@��)�����y�QC�:�Z�ޞ�lzk���
�n��_���s�._ŏ�}wn�����{p����뻣�n�W[�Z�� cD`�*��������
O��~!�zUo���[ e�/���:�}}޽�7�Z���ʙA�dpE!;�6���g�/,=��ؤg�N�4Tf�P��Uq�/�b�[e�(x�slV[�>���r'����*��>,u����E>|p�>f�,�y�s^�L��QsZr^��J�B�U��i������ �8�2& ���$��-�s�mcu���sw��\}K|�.��:z�m)|�S�W�\��Q����z��y��wVm�lu��i��m�2�gT�����#���+���L�������{��p>+���6�yQj�ݛ��LZ���vU��������0�+߽rŚ�	��h�F;n����K��NMv��}�4t�:�����xh~>⃽f�����
1z�Z�a�Adg�֪��r���?�ǝ��8Jƛ��蚙az�½u�/O����Ј�o� x����[�F�DA�w����������z�;._�	i
w�N՛�G'��}ޞ����;����},P�����Ǿ���>��}v�f�����I�z�+�㦼.��z�~�Ƹ�0�ГE��|�l�堲ϼ"7���	�Aa�[����� xl%;P�3�=�����p�m:��G)�|�۵g���5o�U�~�$��w{h�n���q�A�����8��8/�s��H�O�h[�w>�F��ܼu�zX����n�Y�X2X��1T�3Bj�^H^�l�>�P��U¡�c+�ܶ�Wfq@�x}7~����y�r�A�|n���_�w���?h�mW��u2�L���g�ƕ�<U1�n�
>�kѢ
�L<�G
�Q�N�ؾ� �^�����l�Ҽ��M;��j݋Y��� ������`��D!��h��ឿ|�=�&A�~�{z�)uz*������a]v���K[C�l��{;>^�r��쭳t��+^�(S� ����#�vϷV����༥|��/�pۡc������,�+ 7����u%7��]��N�5z��Nr����i�3%�{��W�����qz �u
8@,"/ޔ�"��<�~��:� ��s�1��%=�\
�t��@�s��X�K�:����yka�]`�C�踽�h��*�3�����=��TR��WT�d�`������^��B+��Zi��G�^p��뭻��U�҅u�G�6I�����z���{���"�/ܫB{�\�s�&�S�F�Aʰ�/U��/���_/O}N���q[��&�oЎ�W�+��԰º٨kj��;(]V*�³kTY�_�,eOp��)�+�w���T7��-�x\k�"Θ���Ug��F�O!ឞ�|������y��}���<kRE���x1��-گ	��}r��ҧ�ϸ����w`����KLU�Z=U��дZ(m���KƼ5�+˥xƇG�!�ʌ����v}�1 �����o���c���=�_Z�g�Vy.JI�����+=ʃ�#k<7ðp:<j�����\�0/Ofn�֪,�s�A�d��h�'�续����[�ݮ���������X���3|��Q�t�C�s��vȧX�����;�٘.LU|�*;���p�T�k������ʃ�!{����q�M
�RG<:'���z�d�����+M:G´���TdR�+�J�Y�_{Z3'5���?a'<z�Ρ����3п����:�^e��G��m���_��
q�w�����e?j�9A�����}����#�@�i����1F��
�j�n+�-�B��o@�Ӟ컈z�QɕS>�/��K���h)��@]��kO'��}/G�:���{W��9��s������ݳ���,{��Ԫ�j	Cˊ�����z8���˗�c�����:���v�����Ϛ���[��P���s�=+��[�1k{��7M�VQ�a�Β��s�S���Z�a�jvz����b(�����q�GB�~{��y�(���c�,ע:S�^�m��u]�6��m��ZٿN��98�K]��*�7-X{F��LD>��&\P��`�Vs,���X�.�׹��Ѧ'[t��+��c�(�,�ůN��w��P�{�lkU�X����~y�T��<�M��ƶ��e|��s��ݴ���{���i.�x�X�l�͉�L?/)B�N�g6�ϥg��H;[B���pO"[�w.ꇅu�%�����|.��ཹ]�@�Gx/%�ۻS��n���MG�1�Ǩ���ւ�V���u���g`�}��ܜQ��-���U(��,�K���A����(4zK���o�(���N���.�H|(�т��8�-�������5鳣s~�j��Qhf*�
��P�[�ȑ�ހ�s�5��<�����?Gr�:e�� ����i���.��w��r	��(�&P�(4lbmY�j�������){5'�v�.��	za��G6>�����	+(Uŗg!�,�0Iht��^�N��.1���.�X���^s;��^�(v��罾p��K�Yw;����W�X�$Ž_(~/U@�ˇ����A�/>��������.�/���L<��m;��O�z�{z͹r���2=�z��3~�v�]K���¦P�ھ����zmp��j�%P�����*3�(��4�>4�X��=�DU،e�ЪZU{	����~��J���
�߶c(����h��>��ض{u����`�
�c��S<>T���3^������T�\�\��z�?U/|�'�`U��E���r�0[�������[C��=�	�1_�)��?]u�_�����>���Y�$������o����q��{>�}<�>��s?T�qI'� ����7D��o�;鏛8ҟ�r%��"	p�A{J�_��;��`~*�W�(��P�l�u�&fq�U�i�b*N�^`7�yCG���7J��A*멃uwM�X�Z�R�+�r�s�m�W^���}�G��C<����TW����<�%a�$�oz��U>sW�Y��)�s:?v���:a��3ȿh�r
�̴2���T��y�lK�{������wRI�.�o�1	�x����&@��Pu~��W4�����]g������=�ឡU���R��nP��Om��!�ӻ�ߩy{������L��=Գ���Bf���m吏������-Tz�Ez�
�f������Y뤮ؿ{����Ol�uS�2����,+�w����D"9Q�W��c�l}���?z�-B6�G�f�ݟ{�u/u�m�������:�����S%y���}�<����M�J���x��:\qҒ�_��.�uk��s��b"Co���`�Z�sf'M�O{#P{}�6�SmmۅF�.Ŋ���#��q&��w���"��ܕ��Z4��3���In|>��F;I *5�v�i��H��R��Iʙ��T�m8#�.s[�����5Z�[r�%n���}Mu
�*lD�`ᖸ�9�ڮZ���f:]Wa��+9:�f�R��t���� �f��ؐ����{Es�-�j)u����I�횠tw)��b�w�4܋弜�\�X����T�����_ӻ�>�����#����x.X72����+5+y�,f����$��Ut�+��#�Q=1�#�l��:�㡜��oV�V��r���pJW,���D�����������N�ܒ���{2��V���Q�eC8X���8�Ʈ��7!˫��(`�p��[Ro1�%Z�;a�6���������ߗ���C]��)w��R���X�:+v��%_gj��ID��kWR�o@���z���S�ٜ��n���#3���@ɼ�A�˾�Vv�.SV�����h-���}(P�m��e�2��;|�9��R2V7Me�ɠ�C��,F��[n-����E�o��J�gB�CX��<Hj�������(����!�����4Q��] _>'�-~qN�6:�R�&lO+�1����n���/V�%=[��ƪ��.��TC�5�I0�e����e�C�����#���7�s�N�C+�_;!�`r���I-�w]�V6l��lKo�4f�ŗ�1��Э�U7w \w��r�EH�����Ҩ�־p��M��#����;a��9[�Y���^�J� �m����."�вx	��q6�m��M��}�Y�|��$��a���~Ϫ�k�PP�ň�-U�mPTZ��E�m�b8�TmPm+U������啊�*+�,[O2��Q��ڂ
Ȫ[`�F������E�Ų�
�FZW-q�J�eH��V"֮]�X����UV ֊"�X�J����mU8��Ք�ʘ����S)`��AT�Q4F�|��4�x��1U�P)Z���++V*:�DAT1(��`��T.Z���U)Q-��-
���`�D��i(��b�9��W:'�?k�|���9�{�^��d�߂��f��Kn뽾��O�y������y������i��7i�E/m���T7ht�����P��Η�����<�8��Yk_|L��:��o>_^���z�/����t�}�!1��Ք���T���Pt�s�-��n��>�mL�����D+;Ȉw���o��F������'�����t��_��2��2���?A�a�yt��C>.����ky%�2�U�f��Я/�HGH"��R���Ӻ�d������IX��~Ͻk��BE\8�t~��L��ff����g������%/�_�
7�R�nv��Z=k6�4�ʅׇe{o��p��]r�XU��J�B����(���;W�D�w�a����[�}O�*��6
����Wytk�TC��<�e�qު��7��"3l����{�*Y����"��|���ۮI����;��έ&/O���?�^��k� o{��Ё�"%��]��?����I��o�����?��L���t<;)����R�<�����z����WЕ��T��LT��%:��CO��O؅�x�b�6}}�―�
b�ɯa�6�
��>����:��Ƭe�$��e^c�٥tn���YK���%����8����aaoW<2>�}(���.��|*"8xY�~��>���}~���Ϥ�ȧ�|p7�����[a�EPZ;�~��.p��j{��{:^PbW:�@�|�Nzy������C�����a��P�>�5��W�r�i���W�C�?T��=K�b��/^$[��;^��U�k�;��S��];�7X�_�z��u&F��rC+o_��_��|O��ib��:hإ�N��фW*M�5+�}�x��"3;up]\tݾ��xN߻�K��ף�b�n\�K���%��\��7�~�/�
�R�)��u7��* �tK�UP��s���5i�ظ�}/>�)]�@}�5r�燮_=I2�*z>OӠ�b�X�X�yq�C������������ώ��f�^1=��H�7���]22T�
S�y��Eu`�sz�<�����>�և�E*O7r�#Lc��|�/�w^�/�׾.���b��
�����(y��0xIWK�B��75ǀ�}�������^��u�X�'����;s��a�7�3G�F�Q�kh��Li5��z�������~}2%�fg��+<bZ4�%;L���Y��g�������d�����!�}����CDe�@e���YB�����ҫVb���������o��}t��>HQ�w�� ���y��e;=�Ҵ���֒�7O+����kK�ƨ��?!ٷ�����j��X�2��{���=����8�mr�GC���*̾/{2O�PgEfG�|y�UW�d��>���៛�*�0|��.�iGZ�*�nC�-3T��nڽ���4AA�9��>�ڷto��D�}s��'��^��k޽���+�k����{��d
0�����M����9^~��r��O���:���Re�|�����b���>�B��f�����_?"���WS�����n����Uչ<��֌;{#�]o��i4��9|ϟ9s����0;z��>�/[��x�����X��yR�
Щ� �e�L�t�qwJW�6�5���x��֐��MZ�[QRdC%�����O�D)f_rR��K����{��uP���xj�)�*e��=�[�l���������s�����m��y�75�|��צ�xS�5�ݫe�'�+�Pvu[�u��S3���k|\s[��W~�'ә�jA�R��{<u����:�����hfL�G<7�9^ӭ�=��}��=�w)8��(O||@�xѐQ�^�0d��?@5\ձ]�������	�q���{¥��+�G��5�	�:�7y҇��C��4��V|%����v4Uh��c�ܽ|���'��lR%���P� �~�u��8����YJP�~�ދ󯑆�4x��ZhO_��e�6�t��7��kzI�3l[���!x���V]W�mZZ)S��5ὶ�l�{i^�d���c��\>���
,kyWVn���*��~���������nx}��K*]+f�
��;Y�v�p��қ���+!��sAe��q�����em����.�n/
�+�.�X(bϽb
�Kê���
����{�Lv},,���K3�wSl�#82�G��R�F�<w ��TK�22�m[��y���ߩ�v���lv�f�����MS��;l��B�J^�ԓ��k��UU���)=��tj������fm����<;����.���]J�|����^��U���PJtj�O��U�
O����w�����=I'
w�}��%^�N�Ny@������2�|R��܉sX���/v׼0W���b^1w�(!�#4T�����n��}��۹��.Tyv)	n�����\@C~Z����uO> �uY�m��W������9J��>�+��:����/��gޮ�z{eo��8i���
@{�\@�w�sgo4��!2�є&�@���a���W�y��UV�x
;�z�t�2������	��2�u�U����m��P��:�SB6AԷ�==~���<���9���獧���؏i���m�锒>���4pJqpP���y���;�t�J��ZdU�E�;�3M�ߛ�~짼z�w���g����,��V�ht�NR���Qj)-�t�z��� >o:D���~����hQ����u˖������LeG��Y�c�ΕPR:������8Ӳ��57¼:����Zǳ���W^{�e.�
�ᣜ_g�Wɕ�ƸX�X:
���l���h����urݛ���)X�9H?8�b��=~]�=�zH�n�+.��.<�ܜp�K�w}�u�_G��q�E����c�b���T��A*���}���P��}~���1!���CdO9]㠻J� �_���~��E����z}�v���9N�9~Lg^s�_/G�*	�tʒ���s}�H�xׂ�:'=���U�FK����t�0xu�.��|����vϮ��, x*�cZL[��
?Q�'���b�����sN*�q���`��Խ���	�ĂTgv]��t�����z�G<%��/���XJ��#��f)"���!tF��x՝��d���8�wz�_Ͼ����n(���U��a�_�ik��ѣXi�iW*���߬B*�����=[�o���́����G�,2~��������׉C�4��_3��b#:��/���Gb�"�\r��ͨ.����
��PR���u�N�� ����=��{���l>{���5U���[>*gt�Q��F��'�RG�鹑ǖ/�t:V�|H�=��yr��y�kHW��<�������&��<x���_7Dt>Zs�8gs��>��r���(��;L��+��=���㩴|@u�+��
=����{���K��ľ�,��];7Jτ�UӾ���tV+/�S]yt)�~��g
�Z>`��';0}�Ꭳ幛��~s7�0J��K��X����F����y^��[��؜��C��;����VdI�M���wrn���m/wl��<dKx�r*�����������.
]������?�_��Nr��gG��y���{�$����!�y�}(P8@��y�p��6�$7t�M�3��/�<��M��F�-S��j��K�M=�kx���[��$�wKە|"�R��Q?���+��X�&��|I���y�=�:�`^�p���wzfPB@X�yu@�Ү�3�NX�W��+���G�z�w�WP~�]�Y�7Լ/M����O�#����	�5�ϚPU�	Cp�{�Zj�W��Y~v���˧�Ǩ
?3b�,R����R�>>��,t#ե�M����X���J�	�p�\��?*�[����jZ��h���^*���5f��X'��C��t�<;��4i���ی�wB�`^�G��3�(u�F�3P�?��$��/Vه���2����ٖjѪ��ce컻7���e߶�w��|>�|�MQ�����u/ �(x���������*�iO�V���/v;��/�l��F�~b��|G]eJ��7�zW%�˧��I�;���0��_\>~�y<�Y���s_Y�ۻ����=�)x�Y�b�;��Z�^*P�Kì����}O=ũ�;�˯��=��\)���IXU�\~����5�}x.s���P���"Bg���� �/w���x��w�~W�'�ߥО!��:=^�%|�#}Y]���O�۩{���y���E���4�@��eg�K��V���)��H)��3R
u����R�!Xu�LgY*A@�*����y���߽�ﳅLa�bAk��X����$�hT���k0���1�큌4���l�&�V��Ǭ
��. (�`T��R[}�wyΦ���~��_������~�� �;l��͙d��'�o�H>P5���a���1*�Vk�E��*~E>C���l�Ɍ4¬��נn9���V(���f�_���N�ΝȎÑL���*ƛ[�]�ˇ�wm5!���bڄ�+��8�uz��4P��9v��NQ4'w7�EV���m],W;uQ����q��A�tj\�O?K~�TS�[���x��S{�-�=��5�ӽ��ۻ޹�(�ِ�3�k�����%`�&V��{w�'�n�1����]4r�9��Ù�e@�dX�G1>��8XM<Qt��k-f�f엙xz�w�����\2�wE��C��aKG_]ئJEj]���7ȩ3��ѝB����RQ�y�ы�¯�ۃ�ׯ��<t�.�7#��si8��w��$�*��C'\�k�|&eOvQ��=�To���ۋ��Ȗ���7�挭�u�G������eC��u(�Y��g�S��sܓ�i�̚�cg��kgp�k��T/8�����3������۰�3ԕ�������i5=_�9�j�?~ �-˝c:P��]g'����K��r�bkqQݔ �M����t4�@)�NAr�X��.>2]���\~�y��l�������܇f�c�Z��������9�պG��J��G��Yr��F���D����,��i�r7��~�+̎\�P�>և�Nqʷއ��zEu���
А%x+ŎюN�����x�Y�dq����r��7����ij���r���ۓ9Wi�u�\zd#��vd�x7��d8m<M�Wx&X�*Xm>�6��K =����8P��F_�ǐ��<KU�[�B���q��Ѷ��;����Cy��������ݾ����0�
ȒHuB��rƚ�Hgg\��R�-�[�l˖�|{]�Õ���)���&��<�UM��M��m6�m�A<�_\׿}���tg�y���/��d�OX?��-���W�l��T�DEUPr�d1��+X,b(���AATb*1UDUPWƌU�Z1E��&%E`��UQ`����,EAjX"1D|h��\���ƱDTUE�̘�N�EY

�"��DAQDSMJ�J����"��&��m�"(*$E6�1r�
�	��DA�Z��,Eݧ��",`��T���TTPTQ��_Ur�oUU�4�Q�\�Tcl(�(���ň3IAA`�:k�������O�!��˷	5\$U�u;�S�%tח׻+�E�w�_}_UV��yϹ��`i ��)�L@QN0��4��3� _�
���0����XbA j{� ��5�'YR�l�d��*&� ��{���3�s]��s��x���_Ư���
;I���a��bAC�?8�PS��)18�P��&3�K�&�f�z³l����AH)��b�AM���sw���?w����@��g��a��L
AgX~L@QI�(bi�Y��S,���P�$>E
�RoT�Xm�Oܲi�Aa�*�+q�N�_����K����¼��>>������@Q~`~�z�RZ{�>�+]�9����S5G�!S��q��ɉ�O�La��1�����W�y�y�k��J��+��OS��I���3��d�!�I �P1E8��i<@���S��C�,8¾�+5�ɉ�o�/���~���~�:�ALI��#'YR�Շ��f2T���wH
,�N3�1 ��`f�:������
f��I5T��������?~��������d�XV���O��R��*J��S�,5���B��>��H)��&�Y�J�ìĞ~���J�;�|���<���o�Xi�H.�x�$:�E�T���f�!��Q@�:¦�P1��Xk,1E�ɬ�� T��Z �HV~M0�'u������~���~���`u��xbAO�=q��hzyC�m�{a�<=��J�X~qE����RT���Re��La�l՚H)֐PS/?>����{��@���XT��@�{M0�
����Ă�O�b)<C��42u�[�v��XuP�� ��
����*W��|�~�ZR���Y�b
��x@������G������w��N����G�Mi�nf����$�8�m���ի�:����P��Zb��ߴJVݩk��n$W�ſ�� 6u͌��U|7�O���i ��}�i �*�IS��Ag�K�~@����c�P:~�'�U �~@��f�d���[�=�ou�;��=H(J�Ĩ
/�%a�1�T�l�5��0��I�
�S�H�ì*w�o���&�l��(�Xl���
�s�<9�s���d���?��~@���R)
��a�����<jOR��R�gn�
A��N��~�!���4���X�(�~L�^���~��߻��S�RT����3�=d�� �xv�H(
g��@��f��bx�~�ެ4�l+�'S
As�LE �>�d���T��W�{�{�����XqY� ����
(a�LO��d�嘐ua�t°�<��LH,0��E�����$q��wVaY{����}u��ߵ�d�Ԃ��T�J����@�5����)
���~M$����Ĩ��1���
�{CܱbÌ+'̩<B�/>��u���?~�����������������Q@�=g��I���!�
/���M&�*O�s)t��a̤v�X5!QH)���9�7�����y�v/���k���9�'�����o�& (�xo�M'�RT���yg�LO�H,>�XbA@��N T������=�\���<����~���
�AH(�k%E ��.�42u����Hw,8����A`m�:�@QO7@���0��a�VM�Y�0����?}���s^�>IR?n�Cĕ<g��Y���i
��֨�y�Af�ɉĕU%B����ԃ�!_{C���H(z��|��!�ֻ���.����P����V���F��D�bc:v��,��!^=�ɑWAߒ#h_�o�.�z;ZA�2�|��f�"��
w�����������S{� >��3��.�ɉ<a�m�AH=��������a��1'P����0�O��bAf���a��H/Y:��R�~�O�+;����[�~����&���~�0��֤�}��Ă�'�t�Y<��>�u1�{CӷiIP�J�XqT�)+%eH<��&��g�����߳���!�$<@��|��ē�<g�!�8�>��'�4v�ć�x�!�;��_�}�~�߹���O�T����3l1?j��V��a�gi�u%H:<���*|�,�Ag��B���~���N� �<�1:�U߿w�{�y�s]&ӈ�֤��n�Vz��SY@�R��J�S=�
C��rJŇ�*h�q
�G�H,:�E;�$u��/=�~���=a�P+?O)�H/XoT4�R���߶���oT�aX~�O�T���.$��N�H(kt�hLa��^����?yϿw�R
��z��%H,�hzʝE%a���{gXo�6��
�]
�Y}�bm��l�$�'�r��1�|�� i ��p�sϾ�����~�=�N��+&�R�Q�i���A���M��CI�����VM2��8�Gw���4����V�
$�*ACI+�񏟻����u�����@� ���rM~�+;?P�6�̰7�Ă��*�偉P*��,���0�:���ˉ�Q@R
Vh��4�Y2�os��]�}��~咱a�����+3�LH,0�솓�����1��^Q@����$���&�
L��=`T�N8���S��@���(e�0���e�3C]F��r�ޞ՛�hC9����X��j�k{��f9ݨb���N�B����ì����p�m�i��y���w��,(eh��k�0�����I����o�T����(�?��<d�Ă��y@���w�5H(�b�T7l��S�����&$Y�����@��Ă�_}���{������~����*b~7I���C��B��\k��t|d������5��4�}�7�rT*AMy@ğ��4yf"�S������y��s������I �ra�aY��LC�J��T<C��4�@�״Y3t�C[�0�6��)<���8���H)�O&쟝$h{��,�ӭ��;���g����ى��5�(����f��^Y+3�bAI�+��Y�,*y�$ިc0�Qd�|¤�?9�?_����>�[�
�P�^�*|�~Y�����Z�HVaܧ� ���� (�{혜d��� �@�cr�r�1RT����kۮk��{���Y:ʞ����`bA���ɦ0�6�H,wqE:�_���S�R?R���4���5 �d����1<@��{��W�w��߾��������R�0���+4v�H)��7�CiSt�X~a�>a_7`bIY���P�5�'���Vq�򐯝矿��o\������2y�?{I�?0ӊ�:�̰<jA��j��gSc
�P7����C��0��H,�Փ9d�X|��$�O����=u{�?}�o��E�6�P1֑a�/(��1�XV�x���.�=M�I-�G�3�B���ݏ��>�Co��A���f4�gR���{UЍ��?	�;��+����
�ԫQ������m�y�%���>��l�ZN�ǚ=��ѷ��b�Ge��]�d1��K�WT�3�ܑ��M|se�t˴%�V2��\e�\]>������]$��~�r�x�C<�A��Ax������r�d�Nnk�w�x
��}}y��\���w�>}W�]������ߥ��>�<k�K�U*||`���˔�ڹi����^d4w�?m�h��&wl����5��r�^�N�<��z����r�e���>�S.��ef�"4�wBx\�#��������϶�&��Tv�x){}�ZN���b�/Q����W�J^�g��?E�����B��~�J{����ƥx!����>��kt0n�(C埍��#]�F�`֚�r�|��e�F��(��}�ߐ�����c(B3�	�������n������K�E?A�k��z�?�|0`�8���z�y�ژ����5nX����b�RoU�*;������=|�jM��F����H���p��(T���R<0��VM���rᏲ�0��f�~������Q������ѱz� Z�ׄ:���z~@����{��t��r�.�����?%�!�䁼�`�cR��enC�#���ж+�ס�X��3
ח�)F�;iP������s�}�����3���8���^\�U��P�>R�m�C�o��=/����e}��S�>cSUC�b��x�U'��_~oK~���S�h஬
V��;�?7r�#Lg�\.�Nv$٠})��yhZk�k�N�����E�wJ�˫�;���ڢ< u��
+��B�c]$Ÿ�\~(�/{ٙ��n�AJ� O|UEV��~���FпuPO|uG���f_l`�%W��||>���ᰆ�`/�
�t�^�刺\ʤFV�CF�Qĳ>Z�����[~�V��{��\J��ۛ�RY��vvu�1[j�C&��:9n��WH.�ֹ�L�}j��� �o���]�> | ���
��ܡT������Ϩ�b#:��/����Vv6���	ಶQ�x��n=�
Wo��\#P�{������(���p��4���R��x>�]����C�BX%m�Vj6٩�|���x���M,0q�'������Ա�ٱ�59�������hZx,?h�4(:�TQU?��r��^����j�*���/s����|���Π���^V״PB��?A��z��p�Z<$5��)��s|"���4jx�H��$Qb-VY�h|�v|2
^�ʙ��C�쾿!K54��B*Z@�p���6x��ޅI�tV�l�@U7��Hc��Q���:j�]��K�{{Wz󅼯��x�����=����ڶ����%�Wy�4,�r�}k�J���
�o1s���.�x&=��8/{I�^c��@>�׽;���U��lK�OA�t#�x�>�$24�W�1�:W�{`����޽5<tS Vi�㵒�/����ߎ�|���MEg���EO�B⡱^J�Ȩ�RƸ!U_/a�]k}�9X�ĭ�_o���RS�E��n{��<݃�p���Tj׼�;K*�8{����*�U��ɞ��=�
q�N�ԞO&�x�Y�������n<����g{����n��/|t_v����w�����b�����jb���ܬ4��_o�������7v��s�<j/�Uc��±�W��[F� ���ř�y�۩Գ��W���T#�����Ua"<}���~��$�����`��'�٢��&��F�r�,
��g��k\{�r��R7T)��ו/��ak�e�խ�bEaԍs�T���E�6:��4h�Z�,b��M=���T�E*��:%���#�9Գ��om�������{��i�ߥة��{�ee������mu��q���)<k�/��۬�PF�t�xuR���?OT����`�Ӂ�OT3���d
��n�xW�5��\>�0�/�Cc��q�~c�d�Lg�.��43��nĪ��Bz �/o� �Aw,faño>Z��2��A[���xe2tǴ*�J���5���rwtr�$o���3���+ާJP�q�?Z�y�h{�uoJB{��U_�A]V�������r��7/����,O�s^M=4_��\���f���&�k�s�#����)��7E�|���{^G���<~����F��T�����1xL����.��!��P9ؾ���Y�R��c�X�ʥ{l��tu�{B��ѳ���rQ˸wnf���axSՄ�T%}����vE":��7��N�#S=qtb|
G��E)#yV��l�κk�j��o^o���˝6'}�L�/G_��W��ޙ�!N��T*��;��Ԭ���.�򼣾���_2&�}����~6��W�ؔ���V.VAp�^�o�О��.�������a�~0hl�o��}ޓ)�/��J=�Ѣ��W�q��驭O:�ѹ<w�{}n՟
7����]�,,x+{W���'�6��\پ��+G��
r����K�~^�`������U��^-�����v,�x�9]��u�-�|��ѻ�^^c�9�D)�&�J�#����xhh�Z���P1!���+���x��}Dв��'�H|Ʀ��8�7J:_x�W��|=�e�y�$���>����^ܞѹ��&�ǜ�tgB������o;�۪�r�+��x�bkXWI�W#|g������Ƌ]u�%^2� p�!�OK�Wf�����n���5��S~U����#�i��4�하[�[r���%,j����h}�vq�q�O<�6uH¡{��9j��)��3�[I�qԨ*�d���l�-�ͮi�e����z�#d4�Y��RI�`xy�y�K�vlۗ���F�gʶ!��%%RǶ{��֛Z����d�u�Q���B�G�k�B	�����dRh�5�]����+���;ЌE��n�Q�}���{X�Z5�#Մ=J��D�Qqۚ~��c6�o*f��8s�bG28�|��gja+W)Q��ӗpQ�<���[�ϔ'�o2�oE�Z�z��Z�:E��p�r#Y�&X�8�-�u� )�X��w�,�|����1���=�}��l��7�^��!���Fs������'\����s���*̡s�9Fԩ����=������~��qg8��4Kv.��������t��S�=d*���`�NV��\�v�q��\2Ew��H3{"�d�1`���t��ɾG��~�6��9�=��3�ú8�4��rR�Od�'��XZ�g�/�[��\(��Sz���·�s���*�� �R�j���]}K���4+�)cR�!	�lμ�}�*��u����7�� ^�baK������&�a7s�{�����ϒ�F����iݷ�7���/�.��G��s��eR����A���r�[÷��:��M=���ί��;���񰢛:��&xɞ�y�	��x来�I�l�fL��fw���tlQ:U'��d�.�J�(FQ�e��2�ݽ�%e��7�̑����zZL-��ft�9$�H�H�t%��B#V9w@xo���)���r��UX�D%G�*���
�YSƊ
�UUb*&�D�]!Dcrʂ*��&�2Qm"�UQ�(�(*�jn�C�D<J��QE��TTblƨ��
ɪ��X���UW(�#�b�ɫ,U�Y�Y��L�b)�3-�,�&�UD�4�lXys
����QZm���]fJ�B�X��.:�ۂ���1��n\��>k1վaLFcS+u�\�Q�K�`x�v���im���4�J�Qm��Zآ�Q+O-A<ә�S�y��*�AUe* }F� c��6����AӺV�����.�C7��8�l+�i����6������ꪧ�foO_m�V���\5b�&���?.���/#�N��x���s�8�����3�}w�����u��\��y��go���e^�����>��1��2`��s�{B+�׹��Dk�g�e��{��U�z������>�
���W�"�ݐ��~^�����.��(e���{�[���ҘG+�hLK�)���8Pt�u�����c��f��u��{�[NL#}��[픽��t��j�b�vU&|>T��^�~���ٗ50�ٗ�.��xg�P�����z�����]=<�a0��탽Ź�\k�>1o����7!������� ���MS�b\{y���a^�ߨ~�2�xg��w�G���(Z����A��w�WK�M�]�l�Yꅆ�ׯ5�|��8����sJ��w�.��z������p���rc%
�����U���X3����m�u�,�>�������%=t�WwHؗ_�}�\6�����Z��.8+E��V�X��OD�
����) .���{�����W{����{{3)���9}�B���*x�H�@`�~U:�hL���ǌ��ߢ��}҆e�%�9A�?W�����d�S��H�r&��B]zV�K�1�=z<N�ú�`�O��8�m�~�M>̽{�3=^yB*�]{�G�`��>��Q��莬R��L�۞��<O�n�^<��_�k�� :Ȩ�R\k��G��Wu��qE@[���Ooʾ�̇ACr�M5��+痉�w�ɱG�mT��4W��3ꬕ~���g��O1��R�T��VUj�ɕ��@R��E�2�u��D���%��|����k޼��g��q!���E��C���Zʬv里K� �k^?6���vwCR%c��}t���۷��$1<5��[�|>� 36D��t~>g�o����o�J�	�~$W_�o~��R�O��n��V�ٴ��3a��_
˪�>��s���Bg��sr��v-��*���Zf~8��g��.$�<�?*��z�!��~�����
�J߇^��|�V2�p�۬�t���� �����I��2�~��om�� ��雍)��}~�'ETtU����ѥ��^+Ʊ�K7!ޞ���"�4���B�}�!���~�����޾�����.�'�~�M?��^+Kv.<�'�������Yz�
8�7`c߁�w������i��}��pt}O��nh���Y��"�ԩ@H�WO�*y^�x��x�ϩ�|V}�����V���mɆε�6r��"'�9��q�v��y�w{2����kj�o��]u��wXƚ�%���o]��E�Z4��-#OnX�諭��I�S�w��wI�6ܧ��&N����/��מ������hX[�_��W����P�r���L1��J��O����/o���w�����D�9�!�G߲����
 Q�k b������u��wޘ����⇀�繅{sq��Ew0�00����oe��N�cg��*���������_w��x/�Y�x.���HF����.�G�X��1�����:4u9����$��^�ޙ,WzR�-<#^�T�R��++�F��[��]x�d�/��ཞ�P���xz�0���T7(ʾ;�u���G<�np������r囮��P#�����!��k\��o.�>�QО�w�l����`�^~*�ƫ�u�`���d�ăH�Y۔�8�'�r��+lv���+�tNu�F�T�zV�f��m�^�V,rR�˅�f�J�1��Hfq�䮼U2t�eޭ'��W��2�H���CC<�#��.�u���X6������x���<&��^���^�t3'�:���ϧ���YNg�7�Î3!��3��<<13����P}�!�M	GY��}�d/+�����e��������s8����}���̵��O^<`�׽���]#�����>u�0�WN�iڻ�7��ǿ����#������/|���C�oD�׽��m__Mݾۗ�j��NJ�|b�?����u�����󸂺e�����A�r{UK`Q�������<<9�5�vv�?4�)�c��7�/_���Cٔ�k��}b"2��lk��J��+� �~��^ңB��q�PO����k�sO�K�DY���O��L�SA�=��G@°��; �)9F�a�/aT����
Ӭ˘����-�M�J�/3�p�1�HϮ�@[��l�vj���$[O���{�M�c�4/��T����{�Wv���](X����/��h�������A�Av~ܚX`�9�Mb��.Q^�g�2 ��������p�c?M��p`X'�����Wh���X�8�i�W����|��`�\�v�qYK��տH)�T��~�ġ=���Jw�V\�B���
����d����=N�X�2�F�`��ᛈ�}^76�Z���\'G8A��|6��43�1�|sƕ�ѷ�Y���S~���>��]3%[�>�^|{)lt؈�"�6�f=Q<\q��]1�=S�OA�t#�.x}�/�K�U�6���k����iۺ˻�^U�e
����s~�ne��������z���s�H�:�-�3��Z��:6��&�EK:��~c���7ɝ�
���]>zq�R�r�&0���Z�ĵ�C��Wy0M����U_}TѶ��+߇��U||@�"�/��^О�{޽dWSu��в��%�OZ(_���|�@J���JϺ��������1�vɗZ��|T0U��Ƴ@><$4�3�=<Ǯ��*ѾQ�����J��T;7����ʫ�.�y�Y�4��M[�uxQ�������S�G�jb���~8��&���-�o����>��Q�L?
x����V��>^4�;��N�h�W���?u�=���*��&���J�����T�v9�2�G�>"��|2�a�k�SvSV|��q=~S��"䕷ɡ��!���g.�3^]�K��5�klx+˗���.�L�?b��_���/��`��#�T�W�R��d�˭3��E������"�@�v.b�|�e�U���i�}6duz �V�v2�s��9GO:L�h!u�w�[�YۜJ 9�s����}��=Λ��U�+��~����$��G�y�^���mVzx�ܫ��z�^�+�&�ԕ^*�"UOGBz���|���k�v����4灸g���g���:	2Ǭ*��>�%�k��G�T5�*�ZU��P�և�W�{MT��]�ٽ�蹄 |}�Z>U�3@!O���履���y��
��Z�v}�j�]|����ϲ��c��+K�O����~�[���b*�EF�������y{F��_�A[�ۑ]}r��C��q#QTe�^�
��s\k�y3�Xn���Ʃ�Z�Vpl5^��S��w۾˛~=�f�}��B��BE0l1�g���2��^����G��]R�:�g�wy댧z�l\��ƶ�=rmc�X!H�a�A
�\�Ⱥ��R��195����#)�{�nvJ��W��&�`��UU_lH��ɱ����Y�q��P�����g�u=�C�j��\�O~R�X�<~9G�>ˢ=��]��*[�
�E�R�`����3�A�����s�2i�*����>��Ȥn�~��>���'����u�X$R~?*�n����������W*���M�ƺ����"w�_?J잖�J+Β����Y`��P<��U�b�CF�����	沦����j,�����!�(i~�N���k홊�7�/��RQ��W�u�g�;߰z�������s)\�uXP	E�z�᭪>�hJt0J�\���8��停僉q��ОQj׻��~�Jr��˟����?nŮ����}W����藺�����9"s����9���h���J$=ve�������n��+vC�!�y��z�?Ͼ���O>������ⰴ6{��&��A-���6w�nkn×�۟9wSb췧S]眒�����侳���dcf����:�d�>�:93v93�w��3Kc�O{G�\��tS;��|�Zy�i�*���5�F{]rX�����}�6V���~~��'q����̗y�8j�ic�'ǖ"��)������C�� �#��p�2���.mm�s<C���$�����=�v���Z�xEgf�k�+͔�so4�x]��;˶��:L����n�Z�{=�O6/*'�^�f��5.��Y[�T*��g�۱�(�b
T�ܤ�z;�n w�,�h���N��\z�uw&��Oz${��'\�+GL�1j^Z<#)
�Wh�,*�/{���9\n�:α�M�t���X�`�����]a5J�� ��,û��M�>5�5�/�����5���	���X}f�������N���{���q�w�{DyO-�����:�J��b����>D֧Avk�\��ti= Y�q^��t�։ڨ�b\�,����u�}��Jrnwx��Z�p��9��hs`^Nyý�:E�z��_��3%=V�Y��;E�g���1{��x�#J�\����d��'�[:�o�������J�X�q�+�r�Ӓ�QBÛX��������VG)Qůz3Y-7}д��h�������,�"�-9�n��x�{�{�0��e�WF\˙Gwl��l�<�{(�C[ޓ@����p�yy*�H�'dŝ(��mR	�ON�a72J�-�8ԯ����ANИ�M��fҰD�\*�of񊷆ȎR�a��[�ܭ#�J8��89oI���)AJ�5BB6w���-g2��$�#�wv��`.3Ps�Hl�fӟ#}&��U�4��aS=�!\��1�����Ǳ��x��>���jS�<�߻:�`�}�j�M���_<��ۣ�=�6�5���pz����H栴��1��F�>��CR�U{�'ڷ0���MiK�8�ݢ�ӻpI09Wu���9����	���U<�( �f��|׎nvn��ݕEnF�����|�Oo��MZw(j]nm��l�����A91&md�i�)g��1Yr���2FMիú�il��$�$�I�$�M��T�nU�L�h����*� 1�@��m�-��]�(cUQT�ڬ���sUɂ(�����Y�\U�J�$�kU]arD�ET.���YYn��u_��X���ص�Үa�krᖔU���5�E\���1uHi3�Yuh�TEb\���mo��X�m-�f!F��,���j6�m<�\D�,D�U6��,�J������J&(��v摺����JXƖ�Lr��_,т�۴�V�peG0�[u�(�%��1pVR�69��ҥ*ѣbe�b&&1�Ӂ�q¬mզ�E��.	P�YP��ٌĶԶ�Y��d��t"�[PSyq��h��D�U��G�̚t8��+�B�R������x(��i�yi�2cÎ�\m�֞��w}��m�JA7ojPr_��ݚ���z���X��A��>����d�{)��k�U�_nw����n=�Nb��be���ă�dIJ���r@�+R��q���4���W.�^aʫ�N9W��Q�MWC���k���\66�v����<t[�ϪJ%�c�,�}�V������/�Z�uٮ�\�Ϯ��;�G���s��7�\����]A���f��4��V�%��B�^.�в����CA���մ��"f��n��i����ϻ"{�?=�G~�ޞ��^����}ACg'��p:�Ǥ����Qv88c�٫%���ũ�I���ӱ����f`�ݑ�og�� ���;�N��wv>�ޮR]~��U���3����|��Wo۶/.�S�~9�>��ь�Fq�.���;ݼ�����=�EF�����.���c6���+�q����^��G�4s��r���K��q�c)%��F����TO��/$�G�|�[�����ϔ�Ys�}�%I�>�Ό�aj]y��b�yu�NԼޏL2���<*���<�U�-{�b�g
�z���ޭ6|l�+��M4�bj<\��ȇ!��oZ���Su�f_����W:T�(���
��ڵڗ��.��^>���ם�x9��O��ֽ.,^H�e���V:�i8�.�N�c�z!?�^�؍�">���H���}Dx�NZg�����Qj�U�^C{{�s�o#���Ϟ��s��>�5��o�^̈�q�'%�c��v�#%���}�Ν�)/m��u3��wu{u<�=�^�Ja�y�r[�6����e:�ݽ�k�_{�Hd���j,L瘮�+I��Ʀ�ߝl���1ljgd�v��U3yv��{�0w��w�^'%���Ye���_ԖJ�B�e���92%�3%3_��{��y�}=��no9��<�����k�����5�l�У#7V��c��_�Q���cqt|� ��5Iܢ�x�����`f��kh�]�AYtm!�]�����'m=���7|���`������Gm�ƻ����}��9z�3�J;�K>�C��>��T��'A��{�V���Oщ�u*��x'����bM>�D�~� |�'ʇ����m̿O�yN{���:����0��ױ˝(�
���[B`��M]��k�.�GmH�@��*r6,͈n[?m���ǋU�9����(��}{��L��ƹGCFMV@oћQ�&d7g�YY)X�s"�hm�+_��t����/y�3�Z�z�Os�{bܑK��{s���ת�gP�B�¦z�ߺn��[h��N8�*��%@t�R�3{��wTx`��wa@IX\�d�¸����N�Oڅ��+�ٛ$��U�����ɷ)��[&)�����[��6[�;�?}N�-q�}���ؘ����GeL�x�~�i9���?})~O�����~���fb��˻Zo�I��g�p��O�����j<tt��,)�z��>��)댆<�����:G�u����́�is�u���I�@��4]|�������z��/��O_��0�@��הR��r���8l��U��Hq��m�םQ8�y�oٛެ�]�g��B�&�Y��ŭ;�<�����X!�#5��7��H����1���gy:�&�Q�^��+l�=k�ͬ�}u�ޮ�h:�-��4�S�mi����/��3�����.&�z��wh7Gṱ�N]+<�pj�/%��ؕj�0&�W�[�}���tr�Kͯ�w�+��>�F�3��S1G}��	��u���ڊ?`�7�{�3f�o�����_�b��2^.��.�:��tz�f8�l��l>�����3�D�ߑ>^�*ܻC���Υ���Vn����/T�vxb"�R�8���u�\ޑ�l�x���xqC�G�dOQ��⧖�nu��m��mk8ҁb���L�|����O:�u�M�yHH�3M�����*�hLѴ��)�*$^��K@�㏎�����n>)�x�.�"b�Ϫ�T.�x�������kc`��A�$.�D8B�_,���$�qo� ����1�Eݾ�oۡ��zƤ��^�5��Բ�%s�����L>krY�������kv���Wͫcq��}r���A���l��|W�_���m�����ō�:2�!��Q�E��m�J�dk�q�?e�/�ʰ�\��G7;]������@)w]r ����Tb���;�ݨ�8�!�����Y���uMkq�
�i�u�s�T�'�|�٥6�"u��zgC0���ж��z]&�eQS�r�����I9�_{��$�y�ۭ7�����<d���u�ud���9U�t/G`B"�{���\E��{�z��k���
����l���~�7�"��Npl��1�S�=�o�M��2���W�/9�����V����2xk�yxG�TOzf��e��ػ����~�G�Z�����5}�-���P��{#���z�3��(N�#?c�9*y������;Kt	�ϧ���V��[����K�I�'�}[J0Tf�V7;����ѶS��^-�S�h��>���L�\p��H�}�^��w9�P�%t
F�Ǚ�F/���G�P�F��V�3Bw?RkA�s������8c��q�f�7-�\�z���W�(|��Y��)�E-�c�����W�k�
@��χ��͗�wo/um^��Q�Ҷ.p���v,�e����shdtc��aqA�
�����Nx��z�$�Muc�N�C2,������O�,����Ymq�3]�'Х��19��iw���Ue�Vx�أ��[�ܾ�靴a}�H��2�)غ}rѿL�\�{�[�Eq���q�x�n�7�Q�4��;��z%O{��S�{moa��/�͸cSɤ3�,W�}O��i]wrsg�8�i덱agyv
���y*�[Ԟ\7K^Jn�bT8e{,H
���x���n��~�ȕ�iwi���e;~����o��<��fvpuK��Y�#�!�W-)�	(�D���G,E���PwE�����R��H���!FuJ������'����/���U��+cq��žw�kd�}�xxX�8{�j�:�ʋc�-�l���&l�U�rǨ��QJ�L�r�Ukg6��(����*��_gyd4\��g/8��Oj�.Rv0NE��D.�C�,�a�(���e�[���K/'�u����PE����sa�2l�7�Pj�.!�����O�UK=鏧+�=Y���~�{�u�c�CF��g��{�2�e��,WQqN��⺦o�k]�ɐU�o^����Q�)�/�����J~�Ϸ�+�~Ֆ:��千VЍ����]�U�]���2R���;�ud�"_9H���.S�(R�es����%�.�[f��E�mQ�Iv.J�d�^��y��*F�v- �{�f��u �����ܱ3��Z�0�-����͸˓ܘ�ȏ�\�BQbյKDKw(����$�i��m�_�2BpӇa{���2�u��/��5�!��X�Ψ�[[�U�f^3/D���j�ɝ��jrsy�T�9�,U׮˧PA�q�y ���W;����g`�c�u�+D��}�@u ��g���>��h3�ih$b� ||s��}_���|�d3�3�{�nֵStG:�ɗzJ�qjg��pg_���Y����F���\P8��ѽ/�D���@�&s	��X[iUڈȱa;8�q��+E�V�rX۵�5��%Wu��]���;(��!�	��{	�%����e[��IGF���v����vCv?w�^X_�0���EM�sDX7:�{Ϥ�r6���E��KU��WHpX���W�zr���}�K����\
�5^ẀrN��Y�Ps3�u������'�n�V6��b��=�=�W�bv?eH1���ܝIݷ����<����X�|X�EYɽ���ѳZ�b��u�룗��N�{7V�H���DH�·A���C�
�*5�#}]��޹&<�,��Tk����P��Vww�H*�#�:u2u"������Hf
9L@���+#�{�{ϼk�pT�e�8��X�c1���-}G��w۵���iE��ijQ��p�֜G2�yj������^�g3�q�z1,�v`^���\�t\�Y,�HS�ٯ���b�]�c����^Q˱	�)$�HܒIRp�� L���`Y�k��鍴V���#�����8�+{�3%�+5�֬F�+J�*.:�aU��5���.[�0��̠����EQjc����b
[b��Fx��R��m-���j*��]��6�&j��4�P��4�wu��Vtd�D���b��0�����a��F-���b�b�q<t�5Ji���b��pˍ̹��i�SJ0S��N'�t	-�ɻA]4EQPR�咂�T�̢6�X�DQ�ҬLj�B��J�a�h�y��cc�10���KZ����UF,UP3�� �94pS H	����#Wj���p��������%���N��0q�ǎ���}Q.Rn��s�(D�O�+�}�EJ|���ɓ��cn�J��陽i�X�GQ�+;P�`�Ϣ�l>�yƦu,�m��@Ȕ���V�쩏c�񳺪?>}2��FE���jw�g�4)Eݟ,�ƅ�fE��s��k�ͩ��bQ��g]>���R��#����w6��z�*�3Mbh'43f�>��Yŵ9_���)՘��@Q���a��6�%W�K���j�ːvr�^����ڦ���&#�vE��"�lm*T�H��?n�hU�TTmѤ-,u�JG�+3���]Wgc5yZ!0����]ͽ���He*��ـ�w�E�i=�cT_����K5x_~�8��X�@f�U�[������O�;̚z��bѭ+|+W�7�WI��F�4�N��bEmp�5P�M��;ǆm�O\QL[�%e#�BN<�,�����_�
��q%��(r���L�9wm`�N�}X��jxA^Ț����`�Nu��I\�}��]r�]�u1R����u��5|DL���|��霓�ۿ&�{��۔\���VJ��������ga�?2���_uh�����N:W�ڜsE�-�zM:��u���Ȇ������d�Ďa~˭��mjI^{؆K�¼�zwnN�~�l��h�$(�~���޻��}}�5::�דu��oc`��WdC���{:����O'�a�bU��i��Q�'�NTd��w��q�X�)R���+;ytUpAOQ��,����~������K��^ܺPh�w�R�vE��oQŝy�:L�{~t�ѡWez����Y$c��J�8�M�k6��,T�U��jV�j�ڜ�׈A��ǽ�]���|+!��>�矸D��݆�~�1�H�DLE�o�RVc=뺛��^
,�/LS;�v5M�ͧx]�/��lSn���8Ҋ�3���,���e7 ��`�5��w�=�R��}�h�J�s3��cc�x�n�����ś$VsXs�<���z�	�7�{�4��r<�9���(�<Im�_G�d$��F8����e��������|/�;<�'z9kq�'r/|b+O\l�<q��Uv�G��ޗ�Zչ6�2%c�Ֆ
�{)-M^CAO��r[�lʁG��}����ؼ����|!�籟H:YLw&ron˝������m�o��IMq[Ū'�!�$~ѽ�=W:�)T��\�U3�S,N�B����:�J��;���z���ד�R��,�x��|�u�#{7;֒���%^�6����Q[Ԩ��CD#ǐ.$�>�/��ڵ���.N�v:f��Qu��p��X�t��$���o9u�.�j	�;Hұ���n�-�7��;(�+��j�VJ�q��W��t,��3���W-�=��
������6���"��DGV{$k�ðZݸ�g>�����Xپ�5�|��7��q摼����]6<���}���RL�i��96�|~�'{�����zH�w+�O�Q����7��]J4���Vh�>��n���2�,�+r�o<���w5S�����++Y#�Z�L�2)����=���sX��*���%Dc��P����u���'�^�2��I��-*��||w�8vς\�7�ܹ��ً�J���j�o4�����]�z��� e��P�S~��~hb|��_��!V0��{�_i�E�g:J�襁x�=<�~�X_P�!t�E�m���	�|:��yj�ި6�({_7�u!U���ȍ���Ҏ�fs^�� ���(��*�f�m�:�ع*@^`��Ӵ$@��8�9��e�l���nu�0*�G�Ò�q�s�jLZ�ʪ�ۺ]�
�kMu�K��h�Ω$Ss`��W[Xo>�f��ET�on��ne�͒�j����E����iu~bKQ$�O|k�^���C��8�f��ʚo�+�IϤ��w��R�wp���i�j�r���ݜ���j�њ��ϯgu��t0�l��N�FP��RڻmK��!b���Μ"X���-[ p��V��q�I:���}[e9�7_�M|-��w�,��"&��Y�f�6'�Ŗ˒V��g�Q/z,]�.��^Kӭ�
�S<��bϻ�]��'J6_�ݽ�{�f��/Y�i"�I�Fi��;է�$��X� ��4�����`dy�~l׵f�D�-���>��/�ƶ��Rkz���T��.�X����g>juuA�L�Vs��{�w�Ƌ��I�va؄�C�~��8�����7�K�
!�
����C@�Ǭ�D�/=]]�<[ �>���;��+"c5�hҼ��[}{���b�K~Ex=w���߷D�nȸ^v��=�,�o?!���{Ї�ڗ$&i̹k{�=B���u�S$�Z��z������{��ՒV���_������y����>��ʱK�{{}�%2�0�߇X�����xW�W�g�_�����3�mG�^�p	������|ѝ���nP�7*��k�����ϕP	�C(k���ևl�]jF�ۡ�8���-������o���X>I���ɨFY�dt����1���*Q�i%�'��%�|m�yM�A�F6L��E��8i�Y�eZ#��a�r�ch�m����vļE�v���R�z�9���g���v�-'���f�V��^� ��f��W��3/�$)쭻��}�Y x��ɣ/Ǳ��k����>�∜[Fol-�"�pՐbP�&o=i��|�;�%%��
��jz��,z���J�]7�MI�๡�=��]HUh���^�T@�R�O���wr��H�����d<�`V]����+�/"p�<��j���*K�Ѱ6/���z�p��=��4�hc�/_zz�w�{R�IE5�%��M�ʜn�����\Nz+�3mfo)�N�svڥ��,�U��#���:O�7�n-IO �G�cR3R�h���S��J^䒅�JOǜG�QJ�
5=Qv��w��]����P��\UǷ\����w��}tW]��>�zWNH$;n[�ԵU�Q��'}���+T�\@���{��
`칶%#��L��c��\��'�I��sqG�����Sy.*�/�UUh����[7|`����$@����r[��鶫�5e<�56>O��rONޥ��z���mM������*�^����Q�9�Rb'�������g]5R�j߼�i�jڲ�J~����Q�b�Z{�r��]��ء������5�hw*r�Uk�Pb(h�Vcz�a�h�s�֩6{P۵�����w�,{���}+�K� k�+��gU*ɽ6�t��}t�P����!h^�w	����n�I��ȋ����|]ņ���_a��j��ʧ�J�|3M�4p6����ܑv�ز���)TL�Z^^�V]^���(�3��v:��4ǫKtic���{O��N|��;�%����L@�ڟs�I)�]>�Ե��ye��6�zaھ糴���q�æa���nl�[WV���v��1V�ic����^B�e�KjK}�ٝ��yhD�\+���W}�
*�\<r��[�����q.�2��LJWA�vGt�q7��2����N�wDȑݐ��,���F�ݨD(�X��$Z�,�����./�[d�Cr���Z�{�Sn�ƶM�r+��6�'wZ�f�P}ʲ�9S�_c@=��RK��R5���G�F{6�x]���U�c�̽��W\zE��0b�ל)�CԮp�5P�H��գ۷�*�X�c�D2�4�%�G��n*�!�l@;/	9����\�yٛ4�ZZ.NM����`���s��m�cNq�L.v�?MM�v�ٜ+nW9Z'r���Ŋ�ט�n��C@9 �vqX)T�W��3��c����	��(s�{N���]�,����đ�m��� *R�9�v��3:I�D���,S�Ȫ*tx�����f�z��P���X���&V�� ��M�L[�v�]���j� �����C��΂$����<i���P>r�on�Y�������Y�n�ŋqť���y�ѣ�q\����/���r?Ş���c�;�������5y����GA�q�Hm���/i��)�����8n���]VF����$x�t_�C�&:v�|�ِM�6�.�V��w9:�i(9ᵖ3@w =�wb�7"�s��d�3'uu�3������rH��O)D�x%�˲�����j�ڼj����H�I#�I$E9]y�L�s�˭��^���s惘"���*R�F�5X��LCYUƬ�8�խ+Z�Q}n�D�%T+墊9J��EPV�q*�<��#�r�mZcm��U��l��Q-�r�QZ�ƪ���5�1�<pAuiQEQB�J��"e�Q���T\E�bC0|v�٦n��LJ���Jc`)��%b�EJ�|�a�Q1�U��T*#*�h�b�h�h�E���h��EQB�-�<@����$r�F-A���*�)Q��V��$�4Zʕ4��հ����*ր�lX�����ָx�����D�ʛnQ{�mcZ��7J���%��fYގ�.?ʪ�q�K�w��O�������u������ML��a���Sq��Zb��~4O�m��2��U6�5�g��3yquFU��)��a�y�\�t{��DZFukVl:����]�~����x�ȫ�^~���g��j&{����)H��=�8��ҫ�>�	���L�y=�-?u��O-�,���_Ӵa�#�R������	���i���0���^�x��r��~���X�ؕ�0��4�f�r�|���PG޼���#�I��A���^>mC��>� ����E�N���V,0��R�ғ�v�����Z�Kޞx(6]0I^Rt��p�M��7W��][���eqӊ��`�����1q�{1�O�7�S��qZ����ٟKo�jWr�S�z�������;6d���󛋣�B]�7���}
oB��xxj������c,f�s=q��+�Q��Q�E��'w/gƨ����y�w����L[�ۓ]ӭ�۸= |r�����ԏ��DW�:x�zv�{��9B�]�5���q�s ��\�ĳ{�yuy��=�ჼ⩽�K�ea��"��?����<ԑ0uն���fG��oL�%��sz�Y[Ѷ,,�a�>���pPy�y����i�H_{����uOA��i����ν�j̻Վ�A6ɡ����;��>�+냮�c��f�um��-�k��V�Ex�[���sz;���&���(`���{�yh�zC��s�̏��/���/��_<dSfT�ضS�J�i��v�?<RXm�kJ{�_��$y��oC��6���N�z�Si��x�M(����TT$���
<*�fE��꩎so��2���ute�u|���ө󩕗f�|�d4�}H���p�w�r�k�gF�bכ��}1�!O,dcT�z��S"��O+�[3���}��E�ٔ�U����Sb)���xwfm|"�:*�=��m���y{���hdt�+����b�<<d�_�q�z�����ݳ�1�1t��n
�Ku���}W�kG�uG;p:CI5� .�Dn�e�f�0�b�C��z����3��)3kQ��n�R���Y��Eu�0tkT�ggLx���3ljFj+��t�j�{*��qkg3�b�|���r����h�{���Ef�����7(K�ȳ�ZK�=�]�ӎ��� �X��+·��ygi[��=�k:E%�]������S�m7��D,�tP�}w%2�Yt���F<�&�mޭrh�f��Ӈф�6V�:����֬\�H�Bb����:4��+={�D��d��Fz����({_7�w/0�x�ཞۆ�\	\mi1p�·t{>g��!�'��`�*�{a�{��cqS�zg7�׺&��ڔ�Kᧃ��ե�kz*W7S������U���.�٣�u�q�Mːw9H_���U���E,׹�5`����k��vS:�_g(�em�*]u���u���G\߁g��CԒN6}'�<���u®�r�v��_$�v}\�����$V��{�n�vf����2�]�Ք�#��.Tl�ܫ`�bMʂ�Y�f�]|ٮT<�{������y;.�8�J��E�ݖYh��ʽ�r);L�rE=�����w�1ޥz�N�$��_i[q�)#?1����*�2�<)���V-���!�*��ϴݯU�&(ӽ�)/:��:����u�M��'j�LU%�,oC&��A����٘.L��&T�e.?��v��S4����}5^�]��|{���6��v�/�F��������m`�$
5M�r�Lݾ[��F�2�U�%��ʡ�2<�|,w��Z��.�ޜp�]gz����mF$�zM��)�'�2� (��nK���YV�/Ԫ�~�M���^��?*�,h�u�Ҩ섦��\}ܯ�rz��/J枅]�:{6�YRlTvM��/:Ӎ���b�Eh�{C�a��dI�n3r�9�GiG�V�mx�}�1%�=�>��ɥ1S�?Jdv�gW9�"Wݴu�1g�\��K;5�qzK�Y��xM�޺������= #�k������up�ԅ9���"r��YƯI�m�X��5#(�<����cs�c�߽<+�ת����
�5�<���Î�x�8�G���P���w�Jv�����Y�]�W˛xP	�(y~��X�9uqc�~�] �u��oz�д�m�qNz�S�m�r�}��v���[)�ôNW�V+��ƕ�1�����SS|��r�w�']�+[�����l��Tʒyl�8��ͫc�&��#�}b��Vc���=76s�]2�]u����0p ^{ɩ�2S��p!����u!T4|J8���b��PzԢ�w�N�fTv{�� -%��%|ώ�zx<@�y���}~���${�v�+�Y��;
��ީk�	-�=�Ɖ�}�N�s�����Y��A�d'���jǱ]���}�k�ͺb�ط6".�dc��yp2��NtS��G|j)��߲U��n��;3So%K�
%�:���L��]i��u�7�HƦ��i��v��L��|�s�U�5~�TW�Ҽ��gP�.�fޤD�WW��*r�=腅��rމ�e����hg"�O��i�0Y�;�ԭ�1^���o����XF���y�������wpdA�YƓ5�[��Iw���&�s:ŞA4����bq
�v�a����K��i� �^]�^�;M�v��t�������(Y�3hb���!~�_&33U�2��wt�
v�\�4����;Θ�]߾��ts<�R�l��$�t��ŁJͻ;9<ސu����,�`��6W���ھw���+�:��)ɰ4<����-Bl�$n.u�>6s��G&�0B���aܼ��U�z�ds����}w���.�mzY�.��9�뛳�{�R�y��#ʱ]Լ �Vz��9{��l&��^Ul`[��Y���+�����8���[�1��'�U�7|��eD��Яx�������D���Y:b)��=Qx�mp"�k����e&}��!���~��[{mh�%�81�3i=�q��͎傌u.�w���{e`�w7k�b��ojjd�!KKڰ~����sOR�%��I�����Q�^�C�*/��{>��4�T7�P����lm�)��3I�;��W(���w=�N�R�&H�L�An��֔���e)�w�G1�~��o=r�q���R={�q�n����pN����9�&詫2���V��`S�]�v^�O
G-y�=V�zM6e@��Gja�ʆ��l��żhJC�h��6�:�J�Q�Ï98H���V�f�V{#�Ɗ����3u�c`6�6eW[�ѳꃶ��]�sb��]�t��qV��vw�W�!�/?�b��+�l�Ŕ보�w+kE���%z�U��w��8z�Dm�M�%V<�7�X��p�ե�D���A=��Fr2�V��6�4��%�V��p�23w2v�'ȧ�c������"+
z��v����3}�=���m�F��n8Ri��@.Ѡ[+�V�\�)'/�;2[3Y�Y)��WF���F�J��d�2�&Og���wk	�ޥ��Mک��yd\�u�te���>p����͚wLdU�ipokV�C�V,��,�{n5X�v�՚P�=���dI�|�K�Am�h�0ک��igk����*�s�5���`۶C9��w2:�&��x)n9�e>��߰�v�g$_0s6�/��]kz�G(PhX"�cc0,�B/ȏU*�2��uh{�K���H�u��9!w��68i�0L��E�ų��,��P�&C�|7 E��F)�_���f��Z��CK����y�����}�z�V��_u.�i�P^��Xq�e�\V��7��\�)�X,*��w7"�Oi[ţres֩�����ꓐ
�J�7���G��p�5Mx�/avx��]�}�K����s9[�$6���j�VE��Js�Tt�:��������u�G������=��f+��Tԋr;%��fel�8�W�կ�>��~J��"�Sʌ��D{�
ܲ.Y?R���3pm��n��'����r�VP�OE��Q7*t���XSfX��8�M�U���EZF?��U�	�f�Gu䲸���G\v�NW��ba��|��ہ��	w�v3z��� �9�]����|#M��9,��p��׼R���4�#�W����r�#�I$�I$��O�?=�c�u�XU������C��Rj���Z(�X�TZ�QAT�Xhb*)R5)
�kVТ"D@kQ��Z��B�Q�PP�wC�
ʔm�mR��A)J�i2!���͵1�e�UUE��ciX�(�Rڵ��RV��b)Qk����kK)ieAk-��Q7�8-�eIZ U��1B��J�m�A�Q���\#U�WT��ʱDE�
�-�*�-*+cj
U�+h��������N��m�p�m��ik(R��jV��ű"R�.U!m��ke����Z�Z���d��,�:t��#�7h�ga���$�p�|��������W+Z��.i��w�)��C����k�1%/����c/�|v+�U�>͇�y#g�
���s�����j�w�^����r.p���u��6]�]���:�BR=o��+�zL�f��������X���ӣ#�uz�cz��O��
�&R/>hU�S��1뻲���ܽ�=���v&���*����u~���Q�Yn��2Z�]�ֈ��l�*���%��뺾N6��r�X ���-�5�r���K�7=Fnfot�v�wp������=s����
�O�5[�ž �#��QU��pmp���մ>�}��]Mk�}�)��p�<0)����<$�Q�8�L��x�(/�F�0��c��/�)m�lK���NxW!�GTN����P��gG]bS7b��"��SWj�s�?ub��~����ۯ�w9ۃ܄�|��~�ʽ�`��srY��J��1���}͐�PB��A�ȭ^k�P����XT�lm�tB�s�{��o6G}rǸ:f���Ť-p��%�G^�4�oO���n��[��o��tv��H\���\������]NY�p&�-5��b��;ʓ&D�񈙜�˫�'��6^��m��+���{3'����9g�
��x�������Uu��f(y�	�Oպ_���^�G�5�H�{�W����������3��A��z������2�D;�l��b�f_5����j���;%��q�&I���m�:ڿ>�dg"&�j�Y��"��jv6�CB���6��]��,Ź���s�ɩ��n��@���E)�g��y�A���;7q���:q(2���zk(N!,�y�^�l�O��M��� ��%\2��Y	����t�>��A�#�4�<��ѻ��K[͈\r�0@��4pSs�C΂X�����R8G��2z�+�$���5���p�u�x���G1�P��F�vSeT[rs3o�\͉䮺!�*�43Y��Ñ��ro���h/m�k��Vg���g#��7]yJ��#i��߻^��Đ��Od=�I�t�/3�*��,�#�9M�5���>џG�v���ح�n�c�V��>�r�q��J��yVB�t4*�DV�tf�f���|d�36�Z��<	���
��!�ߞ������*{E�^�U����b�-K�}�Ժ�;?W�]�Qs��ND��_qϯ�����w{���Z#�T�H���3٥�]�^���Leߧj�'��0w�����T'�r;��y�]���K�x ���
�+ǲ�e���onm�R�1����|8�&��jIo}��.y5w��粡��a��1N�ʓJ��T&p�6�z|�J�}���>59����4[��zS<~�T>�L�����Yt]D�2�PۜfĮ���v�l�j{2�m;~���7��j�uJz^lۜ��� ->���{�w����
�wd�Z���n�_���z>}h�D��T8���㞸��t�LY�&�\�pr`b<�T��φo�+r��=�j�(L��ȉ�[ͧR��~���:���^�Nr��r�k7���$�,;��gn��E/T)�����,�K9(G;�y��!s�y��*��؂�nr�X�I��,��&�[cq�ָ� �7w�&���Si��cq�U�rVW��׮��M��;�?j݋~]��Y�����6[֣��vu���{��?sg�.����czn+Fl�N��"���ow�ɉ��/n@m'����͌��ͻ�ǋ\��k�'���xZ�!�b�x�ۭ�0�;Ί�l����*��2[�_z�����.�H��}��ߎ�n�g�������U;��~O-"�7�T]�T-���|�Uv����G��ePޕ6�u-Yֺ�E��sN�.��}Ӆ��S�����v&������c~��\;�;(*�o�|�ӻ�FB&m�'�pH1�D��ub�g�Z�=3�m&�����;���0������;4�{$�)�g�x�uE\���!k�6�s��ל�J ��wW�˓B��l���2{*�=�zR�o\��@	FCVd;��7c�+�{2��Y���]���zw�.`�6�wC���J���c}l�y��z�@)n�[R��C��[ӢҶK�<��b<iF)�i�eB�� �'%޾�ϫ�"�&�g��B�G�p*�G�Ót[CO�tq�����a���*�����M�Zu����w[r�_�>9����l�����`6k<P��Y�����Ky���>DW��ϋ!�����c˧��P�)_����DMﻅgf�ufH林
y�B"�}�����ނߦu9�9�ip5�����1?v��>�{���9�W>=�m���)�+*q��͔A�71�<�y���E7�� �ܸe��,ۃ��iX�.���r9���>�(����rX&S�m�i�;|~�o�w�s�E�s��c��k��t���۫E�I�'6(S�1J7���W�)(��:k�w��dٽ��w�?IM�f}��h�"���큑�j��{����]�s��8|o;��7%��
7�;��E���"���g6͕��FR�׸�N�SRwk�ȕt��{CՋi�9�P|����K���aPu�X*"�v4E�E+�-���຃,c�评vQe=?;w�{����g\2y�H�����Z�x��!ֲ��ϗ�[R�K	��4�aWM_�=���]�9~7~��="r-�/QY�I[�B��Cʧlo=�'~������̓ �R�pH����>�����W�RW�-x�/3;'-�/	�q8�O{��Ξ�^�1�ﲽ[���<1JH���^֭�O���}.^+]cw�#���P<٢�]��@sl��X��g�]�,����.m�UH:>Q���]�����Qi�[��m[o:�I ������{5/���"��m��U���C�|=�%jNKR*g�u���Jm`��������m�L��v�BPz�pya��yҒ�sS��a��Q�ھ��y���Ԗs��;�������@pU���y{]T���%�bd�]e���?�EW!��i;��9�jd�9ԁ�zu:�)X{r�oNp��}�c>b���~눶��y�����������:��d{,oO8ŧKveL{i�����)8:�#Z��,+m����c�vl�;�]{E�^|�}���{�\�������Ә�c��G�1*�3{�lc��kF�Aq�9ol��Ke���s;H����vu?nYT7���nI2��; �z�6*]��Y�����Ƃ��>W�1t�Ub.��7�sdv�}��!�c���I�/�,3�������������\J���[�d�7�ө��V�bl�E�m�4������M����C<���qAǩx3�d��^���lR�V|��)־�f��rsy���l!�
1��s����9h�NˇgI1s��oMzH�āƾ�;���#�%�G7s/ü�h�x�쐄�g�r���R1�xG�j�&ĖY�}&�5��\�y��k��Е�
�l�Ȓy�&�\e�W�h�Cμ9i2&@�'�h�p;<|\��{j�K&�������r�BRx����&&��p��y����z<]�U��Ԏ*�
u��)
�9�ϧ6Yt�ފہ�g� �k�}0���|����X����k�i�x��@��x �w=U�=�]7�8�U�dwBs�Yِw��шi{�͌5n�Q��0���.���l�";Hzf��u����6ٽ�v�՜�3惩��k������<+��6F�\̟m����N�݉a���8��3DU.S���9�_u�2�"�Vs���G���f�\N��a��dѶhs�����ox4�:��J{oXl��3vU���L������@��$ئ��r�	����n�!:D 5ko`�G&��ښ�y݌rl���6��ӈ�?wg�K��E��Ex�P#+O:3
]A^Qnhu]@��o�����K�4q�-wV�Fe +�J��,ξae�>�Rĥ�)��j�6vz�;�h����M(���Auu++[4������N�U�9�������1�5R5��Ł�h�"��թ���5��$D]�ǎ����	�3p�ؔer۬��5j��A��(�]�6̫��2n���M�h�ɑ;l\ խ���}\�5�G�����-�tu��=��G*�]��C�f�2��7W�����-�E�;�������L���"^%��9Ղ��Բ��J/X�z]b�% i����YBuˣ��zz�Xe��,��d���9�r�;yr��]=u!w\=z�=�u=v_/H�I#�I$ESڕ�k����x���.gƼw�X�j���
((���QM\f2�kh����U
�DUX����QJ�E�&+���nZ�PUYXUV{��+��(�
���,X���*EEV*�Z�*�b��F1Z�`����ͦ�R(�v��H���P��*�*�Ɗ���L��b;�uB�T�m��Y���(c����1*��3,FE�bQ�W�
�L�A�`��FQKJ孹l�.[R�*�ʊ��kmiGV[r6���(�1!X�����
�X�q�(��a�AST.�wXLQ P ��=�;~�����|�z�-��N˼�Z,��V��&u)MZi+^=�^ioy^~�ƔCB��Ϛ?7s1�x����8P����`�K�`�=������vgNnX0����o�ߥ�&�L�7_��ݙ�c��R�ҝ�0-���Z�n���:eK��x�}wBw��i���^#XrnT��N�G�W�Cy��Q񙽚�����<B���~���2S?zs�嫺�|��o���;�^�=u��:���h
E��,h�7VwtJ�*�RJ'�ZP
�(:q��S7��!�Z�o)3�m`�\4<��9�Z���3��(a;ğ�g��O��V��r��P����	�n ��uN�a����N��*œ^ y��[�!�X���o�H�@� ���().e�b��t�W���,�_ �v}JJ�<���>���y��z�&����!#C�/H���쮻��Rg2d�\�x�\�SIS+U(3�Hn�r��ˆF1nFD�j3�Q��9��+�!=՛b������M�lb�̫Ӌ�5E	��DN��X(�w��P�K�i��2��qŜ��(��>��{G]���J#�*ч���(�s��R��C�X��CV+���܍t�W+n#n�iyWB�u�3�����sW2V;��)���Y��LT�8ByV�>���.�H�e�ʡe9\᧊� i_U�U�F���P��^��G��x+3�`Z5���Z�c�\�M�[�saY�u�iJSVৗ�bt}}�j���}��0��m{�Un����˾͓��Y��a�ƍ��z?��=���V�h�G'���*N#O�'j���W�\��,�IFտ<��3z$�/ >�
�VRi��uq�O�#��緻�+ܒ3��i�Dc\�^��X&__�_n���'�3�)X8�z{k�m�R�w��׭*�������}�U�\��3�r��'�(��D;]�8g�g���9Mȡ�2�3l�Ĝ�������
�G7\����Mo����\�H)0�����a{�_r�$��Q�B���W��^��@��f����d揑p���H���kav�R���p���K ���D���n�e`Mvvj��ۛWݛ��޵��0{`Bt
Nb3+��S�긺m�7�b��3:�"�ˌX{�~��^�Wȏ-O[�us�Ξ�r�{Ɛu�v�:��Rz���Ӥ�ղ����H�C�_���(g>"uw���F�nϬ��Wpx�E�&�[cq͙���{�0�Qɜ��Uۛ�u_
&̺�+��E7�7w�E��pmëv%��g�������<fsH�&i�ո��3u��av�EM������;��ԝ�c�6���o\gM��O��3 C~�i��
��y^�>�Ȳ��n��;7»Fs
k�@�qм�nn��Xz��, �5J���띉�� �;+��z6���ݝ��L�+�p���ԛ��r�F*wW��b�._2��/�w<q٫��O4������4Ѫ���a��Yޔ�9�su6���t��������!={+�~3f��Mz�A{SfTF�]�7;�)�X^Ĥ�(&a�,8�W���2�u��7�l�i����_�!3��bP�t�M;7~�r�3�U�+�p��MT� �u���7L,�]��x�돨��/B��9;�A����>gu��<����]px`U��k{�0�9����{�K��~wL=�7��B���;���j>�]>��KB�.�"�n��\ˢ�=ɻ}-w:��950�zש��{9�j^���d	��uf�",�٪�z��q٬޽#A۵����ruN7�Z���ڭ)>V6<�9X���wf;��o5/<�*d�j<��x�[3�	��}ä�����W/|M�9u����z���}��k���oW�b����+��W�L��H��Ⱦf�t�^l%l�y9=�7�4�i僆�E8�G��ּ�طm�5����|��=������vr�i[��])b�\��m��"E�����n��ލ8����cɾ����2䃁~U[q�]��N	C�+��]����Q�H5�i��x����{k'��U�m`�sû�36�/:��y���A�ʸૼ�WOy
"�"+<�Z4���A��_]dx^��va:�����w���;P�k����p�磻9"�DQ��(��A[��w,N7�[r̼MT���^��i��C�>r!�{vgz�Ŀ��m��/�j�ץ���!kä�e�!�}��� C�ɝ�su�K"���8m��@kER�
l;X�j����<�VH|Ŭy���v����_z���&р]�1�4�ۂо�;vw���(w[O��H�o:+�I��.u�MJ�G˚���N���L��x|+V���Cn�鞅I˽Z&kǵ�W�O��������M���Rs�ȸ��rǁsm{B�{�*�lّ?O�'���~�`DG�����Q��V��U��.�1
��8��F\�����>�y�=�� ��B3�>����_Wht`��J�z�ｾ�S�ܼ⨤Mb��ʍ���`/wS��t�^��	]�Jﭯz���K��3��K�/�A.~A�#·�I{wlm	흋��t�<�(�6B]� ��!V���UX���rr�FB&k���'˫V]���EU�]2���9�*���!Fep[@��U8�r�Ҏ��G�fơ�~Mb��[���ȗEB�q�_'wRh�CӺ�E�\���������ܷ��K��B���x���;䛏2�N�d��dY��nu�'2s�ز�e����/Zy�w�zyj68u2��|8�Ym�Ֆj����,BɺΊt��X�t���YM��_����zs�-I�O���B�Y�h��NQY���q�sD-��2��v�'�}^�;���vEE��i���ЏuH���t��S-b�"��BoP��^����t�p�`�t��[��[m��*�u^��j�Pl%�o�]r7�i��яiCr����7��r���ħ��h��ޕ������so<�����w���ᝂ��=U�c�Œ�lY��k�d"�"T�4����vF��[��K3P�#o�щ8�p�y�~�7:%��b�|M���X��W>�<�vNS��nU�/aj�2^� �_��&�)c�bF�n��ڷ2��;�Ig��o�|�z���] M���o	7��InN�}��k��A:�h�*�k�tjZy�
���Ӆ]]�c�E�w��t\��4�V
w�G.�Asz�Oj`[ك�#���GQQű���k�5�w�`����q8F��)��*�߲��o~Q�E�ZU�̯d�n��!���~��_37�wZř���*�ε�'-PCo�v*".��XΡ���RˇZ��^�[�$��᝔��$r���x�:�+��+e��}&���u��U7��K��{���je�YsHΫuڒ��tW�Sָ��D[�)~r����������c)H���'��}����ݏ��{Yټ����=6⇺��V�+��T����T�]��Jۺ�;r����t�U:��{�K��W�4O\'��F��ac�o��Y�@�n�����CM͉
7���އ�拸�M���m�7�3���:�`o��A7[5N�}ǆ~���K^K�ĽFM=X�6,.�{�R-��[|�R�%=��*1zH}3 �u���ݣbr���K���{�Kh���r+��#��D�,q
ֈ����٧n���(.�fQ��c `��sB=u,��+X�3kk#�l�slR��wBY�X��y�QQ����0��7ܬ�e��/[�ι�=��n�9o�Z�<{��\B~�����vT�hZ:�[�:i�d�����%`�Į��3�����!cC.^�X�%C��k�"*�ؒ��w��CW<˾�&��Z�P�[�e:�?U=㻠������%g�摲�;�Ң,��n��e��;����w}�K��I�HM+�	�^�FY��k�׽}���LU>'�}�o?Z:]|��P����Q�u�!N'��!�2�s�ӎ��o~i����38��e������p��]}����{X�u��m��R�����"��؝����}+@Z�v.�;��ŝșS]�)g�oy��|Ʊ�I]BHgZ�Z��!w/c��Ր�����J"Z-��؆�g,M���s�	E���)lv�|=���ŷ��@�mGy{@κǽFh�u-׾�[�a�;�D�`n���ڪ���cm�;U��r�w;Dn�"@�1�LGR���c'=<�`�&>��'M��w;��N[g;�2�ll�S����Z�˶�I�I$rI$1'����d�bR��V	*�T�u�[�1U��QiӌSְU5L2i���R�2PMRU�q�J��t�鉴�[TTw�В���PH�a�"(��*�"�q�(,��ʪ�´���7qUUDET�ԅj&�E�jT�V��%m(�ter�0\mX�mk���DC�EUMP�\EDiJV�.Z�mTaYPU�Vaurb,U�,�HfZ��k`֢���c��i@�*
"&ڎ�1T��(��3vSF-��LEY��Q%�V:j�������jZՂ�hٌ�e��kIl�1A�Z"�Ԣ�����b&��]ZV��Q��"���2�ҥ��F��f5�(�_���W��Dy��㆕����J/w]L�uq�����Gd�#ξ<��;�O��u����Ǿx�Jr��
��٩'.	ԅׄ�t�֔��M4���7�I{b[f�W���U���Xm�ɖ�
�Mf5%�Xa@�����޺�;�y�ͻ��;����d���d!�V���;�b�z�^�n-s!�c<Fۂ׹�4�܇�s�১$�W�{`r͔F�0�u���Iov�G�rG$O��C/�@��k2�w(Uϭ���s�o�m���M��6��y�LL�e�;s֣�魕��=�T	S��rb�L���h�9A�@�1�B`Àq��Ş���I����v�b�����<BKQ-���\F���]��S�s�N��[��JN����+8�����v�T�04���ǧg���
ՓK�]I�\����[c����s(�o�)�ʽ��so�/ʝ�[ޟC� �#��r?BU�xM�X�C��ގ��F��~Y�|����J��j8�V{�N�K��8�>��E߳;�h�N~��}.R~��#�������y���A�7����0�o���lG�,T>�7��K�%�[B:�Z�h4�Zc*��O\#χ���T̮��ute�R?[�"�o�$�"w`ms#��j���u��9 �K�' ����K����j�@�`�3V_f�4���$�Ӣ�]��uJ����z��� /��<˾ޑ�B�s�����;�h�gf�ʯX�S���T���a�Doaŭ�K�1�|�d��\�.�smӥʗ�Ɯ�\}x$xP��f�7kF�v2����Z|l�״u�L��vz׶��� ����?>Ԥ��|�I��굹�[�rǪ��(������2��(�ajxb���������**�^y_�0�k��m�o�����o�_N�틕U\�[$=��^�ԴF�=V��*��;X�<�#�=���v
��є��t^��ju�f�n�S������a=����C}��u��v:.xu�t�B��ס�Y�۞rˣsw�l �Q��Ԇ;`g�k8������ݳ��剋�\7'�`��(���-��nާ<���FF0��	��`�b����菪w�%J<*���)�(l��m��	��f{핦�]��z�r^�Cm��Yo;���ۢ�}]�ʏ��]�䓱��/���멕��Yo��=���o��t�q�򮊀oU���ڿL�s����όC2^sAGJ�,�Oo�mMn_1���>c-����w6��q5ٛ���ނmp�����.�E:���yCٗ���.9�hhK�ڻ���>z��R[0���F��s�{����T���EG"T�8�+6-Ǽ�^L��Un��7�M�#��[���RI�#O�1�Wm֛�,x���Wc�IE$�r�dɛ˻+xh��S�˟z^�c8���A$6x�ӝV��%<����7��'�x�WW��F�7����Ү�$��xk(u�8�ӭY)��<�؎��}~�hj��S4+O�G��4��_G�{���'x�`./G�s�����ȱM��̓���kc�6��NU"ho^��^��6��r��6�*2���`��B��I�k��pa�!k�:�)n7i����v��)v{u]�G��۰;ndR��s�,^Tw]�Tfs�;����ű=�������b��0T;(���Nn�T���op��n�U䅋��qnv�^��:����j,���ާ�z^��I��Ծ�{\`/1�.��+9�9y��maJ�Y$��,��e3��ȫ��h���u��Q�7��V���*���5~����M]cm�w�(e>�٫/��B�ˆU�aG��r����qoڰ�r��X��DZ�7\O���@���}�O�P���t���0V�۽�A+��J#<5���3_ţ��f�;/3�;%��/L���66�,e /�+��J�T�����9&o]2Г���ʜH���4\�$o�hj5�I��9��^�v�%��O\�ܧ�!	��w�h��Ab�/�x�l�|�_s��5m-x�&�r6.N��ī!̳�%(���[����Q{��۝�<+]�K!3�%����z@C�Ȇ��x�w��ԁo�^���6)�����5&ut�zlRji����y��}*:�_��1yG�kݼ�R��B
�E��L��ޤ[�2��5�'8��i�ߕt��o`���u32~'�^b�n ^��J��K�
��t�W�&�Fu^.�݄��z�4c��噾ޗZE�����|�7辳9iq72���XiqK:��x��<s�m����Lwl���9��t��s.|o_Q�9M���xNgE�D�Υ���D'�1��k�#�C$��Fvǲ��T�k%���9{1 �N�W$�lSOK\��f�MӼ�}O
_z�j}��u��f�g��"L3�4�k�~�����h�Y��t��`���YAP/��z�㡥�w���I$�~�]}�"�|'���j�Pf�j�V��$S��q5����=_x5��\hL��u�������^����@ȦF�cV aW�]k��3ţW�#��	�<%�����Y�W/?}<P���=a
���e��̱��/��l�X�Au�(��eJ�=�x
��[��z}��xB�������<}%{�պ����L�){U!����z����ԙ.{�nrv�E߼�x}�uj�݂k(p���!�;~����1�z�������W��c�.��eu��D��y�Q5z�����������wviMt�N��l���S�D�L�ٳz0�i�]10��l�9m
So�nX��vl:�f3������L:^�}�ׅ;�r�{MU�U�W�]Pzr�b��yR�<`��X���?*�v���a�}|UJ�WS��%4��.�<(U#LN��vV2��^X4=:3޳����CK�G;�h��>�Lm1Gb�,y����/�Wv�/'u�̜��3�t(tk�\0/�k��|�a�hj4W��ݽ{���޻�%��^��wʹ����c��_ư%���@��F�=��T�y���l�����}�EU�Ax�w��A��d�|�A$�W�y����N|O�*��^skpu׮�
9]6@l\��{�3������t�w�̗��]�y�3����#���q��{0dq�R�_���Lx�gY���{s�ᆹ���S��A7n�ݻ�W3���.�ͭ��{�Vlb�qǖ���7��9wL�7��5�
����
c��L��4+~hf^?tOwDz���fJHm���=vL���s	P�6�jU�"+��kՇk<�e?d�r�yB�7�p+�������|�S�+�P����G��TA�q@��Z�׽�Bm:-j����� ��G��	����;R��|�$���y�4�����Y^��:�eT����;��t���T��+�]��
V�����]����.�������>��H��d���S>�;O0���jλ�y�P��|��>�����\��=n�f��8j�x}۴��ϸ�B��C(8B�K|�%s���L��7�������;�!�Ȟ��!�����z�xD���]N��Rk���r9���p~�enr�>�1��={9�<~����cp@����z�Dzx����U�U*���^k"!�Y�∄C��&�D"��YQJ��(�"�ݝ����P�eY������1�-�m��ZK����	z¦K�b�R*$�*D��QI+_���
�F{H��#_�Qc|��r���1�ۭ|�z�B!�RUp�(�+�r�1��}��9�57O��R���^J/:�E�XՒ4?��4�ƙ��޻R�&sf�i&��®��l`�L�6��D?�~O���]�l��II4��$B!��&���:ꈪ�Iw|u��d��g��̞H��g���v���0v�J������G��K��z����.h|"�#箙)K�����6��V�z,���o�,���_9%���GRxԥV����sיL��*O�"!��8Zm���{]�^��f�;p��l!$��D�$�:U sd�7�ҡk�1���FH��pܟݓ{؈�C����R��K9�<G"c��-�����1�*W��i�0q=*9�1�:����>'G���ڽi�g��ý*Z$B!���m\s>R83w��GHq�]�"��N&|��m�cB=;��v�g��;�V��'�w�u�}�N�?q��z:�0�D8��IEk���%y���&�L�R�x���v�*Z�2�"��=h�D?�O��l+���V�VG5�[��$���j�X���>H�����U�ETQI�^]]VIGͪp�ZD�D-&�	���n�902�lmʶ���j�%�qZ"m̔��3�ZyB��KY&�d�\��k��3��m�=nǋ�ܑ�#��dW�����Q�x�T���������&��?�✑rGOY�M쬕�=T����'�q�6���G���ꑗ��|k~�hD"���:���J�4Z� ���Dk�B!i>����>��6���:|6�o����<��mF��Th/���x�%�ǋ��=�pt��o�3GIT{��eV�w���lm91�/	�8D"��GZ3���N����-ݞ��e8���uTvTYF��v�nz�����0���TI����$��OAq�֍�H�W��z9͝�i"	=OZr�L�#y�w��31�Y�I��cK�o+��p��J(���G�sz&�SI���H�
$�.@