BZh91AY&SY�U.g�M_�`qc���"� ����bH��         7����mݴ)���i���TR�V���Z�+)4�;i �$��ZP�U1 �,��I�iB۶�em��VP�l����։����ZV�1AAm��R�IMj�Z�ը�A	&6�TU��m �k�[M��a%�dm�Q6Ј�U�f���/���3���3f�i�^wmQ2Ɔ�۲ؚ�l��g9A�hL�K[mj4"TTf��A���:�֥4`M5�E5���aU&Dɶͪ���dj+�
 
�Z w��Ϻ���-�����l��I�+�]��j�0��6e���:t���3sv�iu�����]N�i��mN����5B����)��i�B��o   \x=*�Y�jV���Î ��pQB����T��Zi�L.�P�7vd�
�-�qҮ�
�/p�
	�O{�M4�ٍ!�l�[b�m���֪�ǀ  M{�Ҁ�k�� �JGy�z�{m��M��6J���!])�����AT���<�mJ���u{ǥR���m������{7{��z�z��mc[+jwgb�U�Ֆ�  ��BUUS�[� Z;�7�W��Q�mOsv�a�+z�w{ S�����<��oU}��hPW�����Gz���zhz�O���*�K�]a�B)�5��ģ*��  �{��(�}w��E�7.ڮ��t4{�С*��m������k�=�\W��Д��{�;U@�*��}窪� {�`�J��9�(�R�cV�j���Sg�  6��T��v/\�+m �m���������� 5UUv��Y��2U�3��(t�^\Q�U@m��MR�U��(n(�
S&�-6j��F��   ���� -�g6�ulhQ��
�C��w i��ݧ �b�������y��	�p�7T�ʩ�jfɦ�h�K�   .>_`���n\uӠѷ-ڠP-�hP[�� f]g  ,��@i�u�� � .�I��ƛV��ֳ�|   	�� 4�� �;�� ݧ j�jw�]�@ Z0h�k�ЧL� ���@t�L��C�GdUsdجm��V�V։�   -{�G]h� :��\��҂�;�t�Cc� 8�pu����p �v�]���9�N�� 7;n4��      P�� ʕ%F      ���)U &��  	�4"��	J�� �    ��$�J� �  �@�SM���zG�i�@$��B�F���S�O���m#G�<����^�Yk�]��޲�w�V�9��M{�뮞�y�6���u��~ � {���v��}�xx_�A?�@U��W�C�?����_���΅X?��D��W���%O�aAU����?��_A�v�d����9��9��9�`�g73�9�`�`�y��9��rL�'0s2s2s<�na��3�����L����̼���/2��/2�0s(��'0!̨s ��'2̨s �ȇ2	̼��2���*�2̂�*<ِNd2�̀���'0��"s*�ʳ�"s*ʇ2	̊s ��'0�̈s2��
s(��'2	�s ��/0�̧2	0)̀� <�2�̪s <���&`�A3 ��'2!�s<�'0!̨sf�Q3
<ȧ0)̊s*�ʇ0	̀L��'2��(s ��'0�� �0�"� <�'0!̢s
�2)� s
�0�� s��0!�s �ʇ2!�s$¼ȇ0�̨s ��'0#̀�<¼�L�s��'0�̢sʇ2	�(s
�	2	�(s
��2	̂s"�0	̂s$�2��
s"<�'2��s(��'3�*L�s�ȧ0�� �(��2�*�0�̈�"�ʯ0�̄�/0�s('2��(
�ȁ�
�!̠��dG�3 '2�̊�*�"��	̊�(<ʏ0�̩̀L"���*<ʏ0��ʬ�̊�"<�/2��fU�Es �ʯ2�s��̦eW�3"'2(s2)̌��0�̂ȯ2�̨�"��̠�*0��(�
<ʯ2�̬�0 s(��/0+̢� 0̂� ��̢�� �Ȝ�,¯2(s '2̀�/2���(�2��(��<ʏ2 s �ȏ0�̨�̙��2�̼�̓��y��d��`9��y��a�b`9��y��^d��	�9��9��9��9�y�̜�̜�3̜�̜�0s'4�0s0s2s2s3�2s2s0s'0s<���'2s0s0s'0s1�����2s2s0s'4�0s'0s0s2s0s'3��30s'0s2s2s9�a̜���̜��s32s0s'0s<���d�y��9��9�`�N`ᓘy��9��9��9���d�d�g�9��y���<���0�'0��'0s0s'3̜�2s4�2s3�<�0s3��3����'3��'3�Ls3̜�����8?�>�?��}���~��j�bT/�WYOMy��|�9$Yk����-V�n�t&\��lT[��m�kذ������o̤��R�T�Gd��0�hO��$]��EkN�G�b�����Vo-�Sn��9���3uC�v�س�ܨ��5����Y�r�c���ڮ�=�A�ȥ�``T��n�̲$ղ��L�;)9&�^bd�˲sU�dr�b'�7�-���V�ݤ��ݲ�r���X�ٚ���7\w�)��hGOn�b\N#wg,�ҡ��pJr�f�;�5i�C1�g��r�*�'p��Jؘ�~�����W��,�i3���0��[0���mj��a����<�
��ǰ��t �D�,$�q���2~0�����^ˍ�I9�u*쿕a<ɃYT�85�t��̎��$�2�&�Jb��nq�v��=0���Cf7���(v��M��˒n��(f/���·c�
v�+Vv��&�Zէ�9٣��h٘��TU`��М��U�N������!�(Ħ����d��j!^�F���z�޲@��#��hÖY��:�`2�j%]l^=&jD�^ӽaUފ��n��Z�
��
��tD��Rn9��)�P|)y}���[���`����(��32:��Q��>wƖ�|V=c6��1�c��1��db�Ƭ, t�%H�^���a9�%���fTɻ��^*@[ٮ��3Fkۋs��"�Z-�L�P/��\�۷�7:�-V�kV B�@Zڴ���ܕq��wi���mJ�ݦ��Z��ۄ���ԝ»��໭�(�bFk��'j�l��� F� �"�0� L��Y�Um1(k]f��� ��G��Ř5d(k�N�ˇ��b5R"de0L,�L�0�F���������WG�OY���0I�6�7���6d����[�4�֮зx��	V��A��R�X�+*�tXf�k�`�bS�u�u�Ѽ�s#�����Ѩ�ي�=�b"�L��Y�f�vZ���K�i2��>,!��ZYn����b�3`����3%�j�e�w�J\��ְh�תCv�M���J��(��@��$c�����X�T���X������4X��U_Z�7O�%Z��Yg�օzꛆ�
� ��x�m���Ѹ4���{f���e2����n�"[uq��g�#�쥙�^��#�u�2AN4D��y�+�7�Q뛨m�20��1�d36o�V0�! �vi[����f��s�v,�a�i��mBE]���-����U&;�y�	��d3JR!^î��XG�ö+/4�M;��x�nl��!�\���sN
۸2��D	��@�)�v�,�T���9��U?e=*AI�!h��9޶��6ѵ��$ARkW6i��Ń72���e74A�.Qg��4�^��C{����aZ,:O��� �۽��LzA��[ WI�J��ڌ�a%�R���M�*�HH�YVC�,��3�����&�.ٰ�e��"�k+N&��M�ܒk�maA	��^�cյ,�*����
��c��CB]��R�mk��h�hZZ�m��V��m:��Zs{4<i3�oM�Y(�����/Qu�5�I�sX@�1�i�MX[A�ve��t�����7,棱*�ڏ]l��~�m�̗fcKn�&�2ԣ�欴&�����u�S�L����٫D�-&5��-�co꼽�Pv���Ш��r�A� �Y��iʲ�(^[yA�WL�c9lj� `�8aN쇗d�5�/`$�K.K���dfQ$Rb�ѽR����ִv�zf�OX'̤��A$���&��h�Tr��s
#Pk�p����D6`�J�8�ܚ���h��a�\Y���֦u�
6�-��	��h�����w5��%H�YA`J��m���Y�~�wt˰~��w�u�a^ ���,�&�h롅�v\<&�*
�[0�U������n]n�ox+
ʓ�i�{�y+�oH�fVc�P�ֳ+YܙVɨN�����0�s!�S$�T�)^f<S�{E���O�	 ��mhw�r�77bxރx���ϊ�Y
��3��T�(iУ����éZ���oR��Obxe1j�ÛA��,!�n����kl�z4��]cuterV.X9��L���u�͡3c�v�"p#L�-L
�nސN�%H��8�k�%]]�7����Ҏ�E)|�#l�zq�fs8���S�w,$�e�8)!Z�h�H�T�f�����L�Xv
"ힰw�|֍$vZ�KI8�9o��ӣ�YYPnH.�O&\;���!bQݿ�43,S3V5r�������B��n6]��r��.�T����Mb�S�+eX�ܒ�v�*N!Ѕ� �0ݷ�-:�L��U��Q�c�
��*���Z�ˢ$$�^lw��"CCc�����oo"BW�d�Q+ɋ+l�@�&���H��c��WM�ے�{�nt��*���b����fn��Tܷ4����6!JE;+4Ḱ��y��X-G��h���ܽ̑5��ö-��3#�I�,1��=�{a�˩QE,���E3�M����R�J���c׎O�gv]��SZzM0a�!�-�T���is3Qt�˙��$JJ��d�q����mД����ʇ>��lɉ�߶�� ��ˑ-&��� D�CF����45�s��3��޼��6���j/5�n�-Y��ayH]�Tӆ����m��b^mi��I7%�`L9H@(�V<hh|�;C�6��+Y����v��r�I��,���1��S\1�h�e4b%Bn�MLצm
J��K:���ۥY�[t\��Pg�wO�Lhourie�T��T���ɘ-�͒��K>�j�H!�a{CV�ۚ��7]'�`�dK��"Y& ��`�f��[C c��x���5�l%*Q$���ղR���vPŬeG��"��W۵�C�g�+_���8�T�1�&�E�-4�u>����lb����F+�3m�(bɪ�U�/aP:J䂶▙�L���۳yeVh:�a�k�wy��Nn�Q/�f�խ�ii�RX��ޡ�RO����j�[6�P�K�Ό�vKWcK[���Q����G�@�km��R�f�f�wE��Y�	����v�,�VBsRÕA�Md��(ˌ�=�4��������b(����T�y2�F��b�����/-�Lb���2i!ʒ�Y��ҫ�ݽ���M��h1����⋛/d��|�,Uo�����}�B:*���AI���2˥X�˕q��\Jm[�R��.�(6��lf4Dl��Fc�;�!�Ґ����2�eǘ�q:BE2�wT��L��4$~W���=dRԭ�#]/�ŦΡN�/�x�������	3�Bȇ�6�:b�1���Q�f)��Ga�u�e#q'�Y�ȼU��r��f��'ݹ�Z��Ɔ���貅3��C9��Xk]�`݉A���dHz��G��XU�]���ڒT[Gl-)� 򖦱��e���R�ۭn��#.�K)KN�ǅޫQKWl���IV�`��0�
I�Ֆ���Ś3nJ!���ͳ��a�rB�f���!%�w�MZY"Z�1��dφÔ��5\�wv�)�"`:3
uqV<���j�a��q"�0��L��f�����F�n[�cspO��^(7.�Q�^BY�0i�t�0L���B�D]4��J.�1ֽ�ȯKzv��y��Rcu��@��
ȞM���ə�w%i;�L�ڬ"�BDh��,X��J�1�8�B�{�
�k�v(Q�ma%�:`e�6u���t���^8���;zi��y��a���B[	�F&�&�]��E��Z���k��T�ۣ�ݛ�s��	ȵ"�Yu��+V�,�`¡�2�����JsMQ�!�Й�.+�HAr�\Gb�m�o4��6��Jc'r�DUY6�(�MQ1&.�۶�?��"�3M�����wM�K�D�#�g6J3?"�H�VmT16�f6(eŕ�fZ��v�7p���m��(!����1��4H�-ڊ��f��&�ٔ�쐒n�҄(A�sr�:xu��Z��� �hV=;�$԰��3өS:Mh5#�џE0������A��WVU��Ԃ�"<7��Y�zU0�#�1)%��=�"���P�S-��Յ���.B5켤�٫&�wW���t���E �A�Q*�l�KR"X6k�&ź[�jnQ-�J���Cq\w�7F�gW�\��gu��!�z����#fHֵLǲb�pʡjP�Pj�[���b��.�Fܴ�� �݉i�r����ٺ�2cf�CN�kE�*(�p�8(�<�:O3)�A�(�r)�V�1�Gt+7,�Y����7F!�ƎU�3�T�������0I�e��n�.�!�5 �+D�[CuJ�af���(2�-�wc2c�M�j���_hـ�V�*��"&��ܱ�P�z�s
x���ͽJٍG14���Jv����.�v�݂����;�f��&ʰ�(���$1��Ph����L��vY��0M��4Y�n\D�vȀ5�)7[i�Oa#o2���
XGY|0|�mf�j���<�J�m55�E�����e�$�1[����\�dڤ7J�?=���^�1��P� �;�>O����A�l��>M���%Y��-^63H�мsi@����V��o�i�VW%]a9��:Yq�U^	�k�Z��U��6J#\�"���R6f���2�͌�"�l&��#�i�@ɸ�g#Sr�ytC�tK��������D�[���컊n�O �zp��p�lO6�7���t>�A�5�˴$ZM:�&�{m�Z�ܱZ�l)��2��ǋ�bHF
�S���-�2��Q�O��9X�!#�Dܱ��Ԭ��mPZ�%bƎ� m�0���ͨ� �T0l�8]��Ur�J E����E���LXӻ;C\�m�f���j��&2��E�V��n��̗4̬���Te�7!��`m�Cߊ��[��;7vl�4;�V8 d4U��VTKm3��b�ޡ��
�H�1��$���A�z�U��fD��trX٥ǭY�[&m�;I�`�36���o\�N�m�A� �f(�����V=A�A���(�ܱE���Ccw�8;�2�/��svM�D�PD��闠�Jm^olelR����ˬ���I�.�8�3QVV2���h���PR�ʵB^�&�jd̽;yy�/�+!�K3�Q��cDP�75S{���2�cѮ�r�Px�;\��]����rA!���*��C��B�gX:9a�i��{��eZ)���{��rV�^ܤA������2��cpV��B
X2����@l��eB�$U�49gl���j�xY�Ui����kn
�c�Ri�۠f��L`�/75���{���8-E��L�e3�.���wb�[R�jd���k"��A��X�?0�lor���^��I)�I�m�d����E����9&`j�of����m#�H�Q���M\1�ۖ���º�w���vu8�4Ǫ�=ͷ���h��u'ma1]�ԅ+ŦR�e��\5�
�D+r����L��Un����1�ݩ���V��Ȃ�DgB�����-͘��W�z���e�YL�����5*
ꖺ0CDڷFc@�t�h@Vϰ��F-����NfH�ݒ
�4�z�4E��R�*��/�kڷ������Y�}ذk�8w.�H4�tX�����cKu\9z�wa�V��n+�~������������y^|� ��g9��v�hX��m�"��1�;+K�L9��H��#{N�9A
5����7��C,�ɢzE���P�e���V��3SF���jenI�n�V튼Z�m;X���;
ɇd,��ͺx�,��.�n�w�ح�[��pn��1��tB�eӬ�j�7Y��KAőQڍ�Zڽ/�]&������.I.6ط��i��eb�B�<��؁�w��r�[@���%��|�c53X	x/VS��Qڽ8�L�7o]'n�r��&�)d1����s�^�`�^%z��ѷ�j��3���`�+���K)-`���̦���*%&>�0����gdu��e�U������Ɇ�:����(x\��{���X��9�f�tưd�V���v�f�7B��w#bh�x�(����8ks�Ԛ�{ͪ�T`a�Sp'$�,Sor�d�aצ��+r��#�&���1����B�	��1��ґP�Ӻ[*��:I+��l`�c` 
�0N2�t�-��V:���j�#�۴�ɗ�1%l��Cs�9(^Y�Sl(�r-�e�Y8���FU0n˸��60��L����Ƿur����v��A�$��z9�q�f!xGtC��ȋY�Ǘv���o���=�Օ@�e\��.� �.���'DxQouk{7\I�7��n��$*6��y�KJ�c^9W�[�K�Q��r��uQHX��`�5���`�-���1��k�M7ӟ�Μ{h<ŉ)ٸ�T�����B��S�Q
wc��;n�]IO�Q�S8���E����B���D8a�8FKo��*��րѵ�gf18�W(=�3�d �ojrW�qkrebެ1��A}{�,�q�\���������I�w��u�35�<�����W��wJpŮ<����QL��%^����]��@�N��z4�B��Q�h�ʶ�x��\��հ�Q��w#Vl�W"ߎ@�� o��KՎ�uCj�tK[ڄ�S�^&]e �&o�{��͐��戋����X�Nς���1��t��;h�t�@�&����a=���um��B�R$8�e��y��k\�"�>��7<�l�e��>���>�ZV�T��~�}ō���P���c�ZU���[�b-�u.u�O�%�}[�w�v���}����;��5��3�I�k#��`hf ���e�h��L��3�5����}vsmq�t*�ٷ/���'���b�����P}�����LD��߀�������:��^�:v��eteӎ��އW�71I4��_����E�:-݇��r�[�K����
�;,0���Dz��YGej��:�����2�k���nsqWz�M�����88�iu��d��V\�N��`�Y�+4���U��8�e�:���`�Z��z�XG�1�	[�#��n`e�36nM��p����C�&İ�1<�B��#��ċ�gp�f�.ê�Z��<�;˄Z��3(�98�YC���(����iY�$�G��U��R|r+�vQm_N����U��O��6>yt���b)l��% Πhڽ+w�7"M�hU���3+�Kt�����:�	��c�%��b��,���05S4�J�t���!�vt ���U���K��ع,}e�o8��^:\1U�/��kV�f�V�����b8�]M���X���Vt�S4�:%;��f Y������b#����Sv?�=ʶ�VM[~$-N����}�c
 ��1ks��u(G^QU�ĥ�V3�kدh�e�uW�e��x)��5F62KN��^W0��V�ğb��#eA7���s+���+�����c�u�]B�/��P��Y��^\��cv�`.K��A>��u��ʻ�Jٱ;�רs��-I|^�y;� �2��v�QX����!G�U���Fj�J�ѐ���ѵq(H2~!hЛ�V"��QYeۚ������d�̛Ɛ��5����4�e]HW[�q�c��9�W&�#hv�ք�����[��ć[��3�)b]iWL�Mvlf�I��.6�kq�Z�uX��RQ����Y��&��QlF�X'vI]�0����lL��f�D�G��quǇ��◂U���𡘰�����9�霬A��T+��T��q��m�s��<J�5�|�ao$�;�H���3/U��%�okbW[�ˀE�1S�0�bY�o
�^me��=��J�mGݢK�z�6)�E��v	di͘'E����fSM�f�[���i-�܋�.t(��l�0�ŗ�5[\1�Z!��B��o��k��8m
\��v,�z��-U��Q���x�ǖ���d[#�V��tv��,|�u眦q�zn��u[���#4���%�MI���V3y����[ֲ�8x"2�e��0�v	��![�zy���+ab�)F�ih�[��`��r��4N헄V��+`�ISخ��3[b*�Հ�%Qc��0au*7K3�p8(��۹Ln���)�ܰ�8�{�>�n��ߛ@��=å��R��.�S�2�}/����QW)��N��Wv4��[�P\U_0q��ύe�2�P�)@�/,b�=��R���<�; v�W��/�T���dԍ
뾙�^�6��ˏ�"���Z��V�dK��q��qL���oEQŠ����.X:*�G3I� g���x_:��f���91�[v��d��'����)�}B��Y���a�7�+-c��͢�{��#����/��\�#�;���_���h�J�����J�@�{	��Y��5�;D�6�x��}��}ul*�e�P�w�5b�����@p�ٰe�Y��"�����oU᷊��ؓ�c��v���f(��a3l�ՐqV0*�ȗ����Y!�Ti]c��y��"��Yޤ��m]��r���S�żz�+�մe�K�B����A��q�P��[:�7��ՎR�=�e�f�h�˲�_p���'�`NF�W�[�
��ٝ�mG�u��n��oo"Z�龑v&azoNbL	�/�Y���K]{���M��ٶ��b�
m4���&3u{d��N��Y�K8�yǤ�l�;Z�a}����kt^�]Q,�4Ʈ`�=�ls�����9WP]���.6tinT�@ٙ*�f�P��d�ݜ�6��U.zu���gH���S�C&&�������5���,kt��t+{�4]�]�L��ZU�Z6�����M�2�t�k�oy�%��U;ȹ��\U+��V��X�,�2�
ܔΫX 8
�r]N�7�nZ�;Ph�ue����Y�$/sTk�+�}R��i{BL���/3F���ˮZ��N�9��knnn�2� *����{ ����S����Ç����w���vkQת�"3zŽ�������VM����t�F��31e��]�8V�Ek9�9�tO�q�niy�At�V���L��B3j�^�X�{
��|}��*_L�GWB�^.Y�s̸���CFq%U�c	��̺r�6����r�:x %J*���L&���̷S�f�:�\�-p�;NH�ɩ�v�P-_QH}6R�n�;�qɯ�p(k��0�5��u��J�M��4^s+4�)�ggVA�퐩�n��Dv�s|�5�H�P�rsNKJ�֘y����_��Rx��
� J���c��7*�{��v�6V�۠�R�s.d�7�����U1�b
��m+ꥆ���-�+Q�2�l]|�ɭYo2Դ�4���A���;�s3N=��&J�VJ`vrx�l�P�)�3m_M��V}x6��7��ijƚ��\�)��I�enHNk�����iCoS-r0\˶]=Wt�MS,�˟l�[�ã��譣3���mNwH���V��(�ɂ
$�f[]N+��i��5�ܖ�l�4�;!�������T�j�;�ؙ��N�J���Pٌ���{���Τ%w!:h_#RӺy���7�3*+��� �lL�i�
���͖p�+	nリ-��=X�;p��Fn�Yͭ����+���+���.�:Qg2dӓ	�+б[lP�^py��J�N�);zC�S�WG^����VU�r>����2��{dW�9������GtI�X����%2�m<�v7.j�f����Fkh�NŮ��d�CT�I�m	��@�$.�X��!<�ӸOŘ�$�y̬}�]l6u� �Yq���Yn\Ú�ǥ�Hά�E�������wY�P<��1�]�����huƬ��t�,*���7��E�p�4�V��3���hu+g4����t�XV��ݖ�n�Y��n�}i�A3Bu��.�n�����T蹷	B�d]���f��-)�8V�C��C�Evee
s�HwH��[���eR2l����s��������
��)ц��k�Y�͡Fݩ��Ժ��;�S�O�s��;%v�c�EJ6q��4��$]ֲؑ��]���Պ��0�D���>9�6u-}������AӮC����2��o���Y���${,m�3,I|�L/��3Y4������IzT6���K-ZCj�y�;n�ӳ��F�C��9[��gRְ]h�K�(v_V�l��;��E��ɠӃk%[��Oxt�|y�V�u��8�xS��t�$�%�����#�9��B��U�/��9�Ĭ���EH"�sN�6��(n<�f��bNQ�ב�g1�}^�;Ou�n`�4"�LD�6\���pw�-4��!J�SJb-���z��iU�7EI��X�O��)񵵡u����)�Er��	�R��Fh�s[c�C�nt�=�*S6�ZDuxW%z�ý.����u|�*�U{x��\C�OP���K�\�I[OQر,/�N��e��F�+��#��Q�Y�*����i|�v��l[p�8�v�5��M	�样������D����hV_vk�x��8(?�אbV5�}�NӼ��l��i$�VJeǉt�.�[m�Iy`T&��ki�y&�;�o^b���Mr�u-z�nZpM�b���n�s'#I��%D���S�˼��e�֡4d��S^&�����m极���&�f<�L�9t�Fԁ�N�=[�}*b�hC�]��F��F1sw��U*L;{y�K\��X��G��A�����/hƲ�v�.�*}��lW*Rח˖c|%�)�ի�uL�Tb�֑ӊb�� �Д^S�c]��or�4�(�#�}/w�^nD$��A-����&16�!Oa�٫��n�ͼ��2���s�-3��9�J�1�X�V��1*
��nЛ�]t6*k8�-�n��UǣF�lS�j�L5x-֍�%�g8^\�UԗT\4+3�g���;P�
��e�]]��q�{����h����!XU:{�B���A�:�FfЪ��u�D�a�fK�f�v'C[5.:+�y��ްH�z�󜝠����y���̋x�����b���qǷ�],4�ӑ6>�B|q'JIyQ��{b<���Y���o,4�k���Ȱ.�و���d����x8N	6:����r�8�p���f�����F���l_��F��ؑͰ�@�)��!�����ӧ���"ЙܭPk��s͗�ƮO}�lf�d��f̦�N��9+��Y9e�U��V�Q�v6���.>���mY]�su�Uؚ��=�ޙ�c�nu��XY$��?vP�h�=	�H��K7z��/�Z�c���i^�v����pН��(<W ��*c@��kg; �m��ۭ�ЌB9�̡K"wKU"~����Ϫf{��j��3Jv_ &$����Xw����'���U���,��x���t����[��̻���-�e�.�Sq>����3�y.�\�;|S��u���N��A���
Fqnja��v�h���YÃ��f·N���=ӝ��=���R��`Yd����`r�sM։��)�t�J�T���^�R=� Ԯ�7ˋ�<Ö%.F��i���o�)ǔ9v��GzA�7 ���@Rw�g+F���]&#��f���m\
׮��(�������T�|��w�=+b�ͽ49ܢ��"H�蔜s�{)E�Ws��c{,���69��T��l�u��^�B�<@!�*Qc�ʂ!f�ďe��uA�ѣ-ԀPT��䛊^TXJ�Wcڀ�z�('[km�0mL�Ub�Y���_h�$͆3��tiY�lT�6\��]>|�}W�%bX܈5.ݬ��-elݗ�Sm�ʉ���ס��#@k�%����.Q�l�m�	Z3�^��.�X;��әdaXŭo�'��)Gy.=�3o��o@vfҮoP;CU,�Sf-v�GaS���@�bb��f���+S��P`���%ч�5�G���""�D�T��\��P詩R�*�)��b�Y��sj�` 6<��X��E{� ��X��wSgs>��G4B�P��5�V�}k%������ͨ������b��\��Zz%�m>T8Yur��%���޾$��Pӡ!A;oASU��.���':|v�Z#ʝ�ʤ�1t�vBq�w����h��H�KW�᚟[x�wL�J��R�� ����k�mM�!YC�sj�qR�m�� �����૗.�-m�ލ�.����z�2MM�H�M�؃��ǲ��IC�X�/�n�R�F���m)�=�b�ި�7FS�.��@ݽvnK��n��q�4;�.��,l+	�a�0v7<���:�Y��n��������%r���ط��6՘)-�\O;�BW�B�w�(��9P�(fڦv���#��cJu�@�.��ޙQ��ޭ�R�u��[��7}Vn0v�3(�J�[�:)nSOOܳ����f����eɉLx�<����T3oA�9��4�sc,.K뿛׈]�)m�o��ؾ������0:���u��b���{S��n�sv˱�I�F<ŹA8�I���C�� 3�d*K&,+ssA�w���ء�_x�)��	�ul�kT�gS�X��V�C� �u���d������ھ9�q͸�E��5:�2��}+(�[Ӌ28��a��>�]`/K�x����3ĢD�fi�I^��uk�!-a#6�NX�N��
�B�L�w�PZ&�+0��4r�����lţ��jh��s@����Z��w{jv>��c����v:��"�5b�2�@��f;�&L�q_t(��y��m^͢6��ɏ�f�W�m�I��כ
q�М��	��uf�;LC+7t�N��kP��{$��,��6�������;��(r>cGf�������P��C�jsڵ�Mݦ�a��V�Í^7mS��R�G����5b���
�3vUJ�8�P�OHw��HpԴ�t3X��=�)��w��Sɡ#�x;6�A�S3EBX�!�%K�bNt�vT�d�-�$��%�#`޳�υ�;���\�xr���aLRD1�r۔������S	ܡM�S���M���1���6ԢH�K!GQL��$
(�.����0l���+�A��0��q��"i�d��(��I��m	jAP�`�R�"!d�b8��P�(eHVL_����h?�G��)�q$�Q*�b�N�Ē1��h'��qh�A����펍yi�/���>��$Q
!������
$�F�'� ���!�M�Э�əM4b)��v<��g�b����^Lq�v�GRb�c	6"�,�����*����_�R�A�BS.2]%RJ__�5u)��0�M׉��B��
(��n�?�&������b"�q�a��̅ P,���T�I�M���(�YN),ڈ�֡��6k�a�� �I_�_�m���A����ā���k����ty}y����QQ�?����⪢|���~u�)�s���~
*?�����A�=�{������a��\*�L�Y���V+�8�9�Hi��zwA�b�Ue.��]8��Y�D���5�q�x��s��s��U���Q���\담�n,+:�c�y+�Ro��k|�J�Aܧ�iy!�cenH&��:�3�=y�N�W%���i���6���;+RO�]j�9V�8ػ4*n��V�N��|��b� bDb�2��lVHf��V(�\��Y���V"f;�*��3��Ղ�M,-lW]U�>$:fc�8R�T�M���ʕ�M���K(dl􂮗�.�ӆ�f�*�Q��9{�_�V�]x�M�	J�#F�U�y��(�mk��D}�6yRG�9~u�b��k��vEԥ��y3X�-ou�>MBމ6�W��Q.ގ"����sq�\	��pV�GJZ�o`�Gu��_�u�uGi��M�n7�G����9�bFiퟤ�+1 ��%��+zkp0k�I8�)�Y/��^eu��V/�d�d��;V��:��n=�M-�UA��%��B���]Oa��_Sr�9��5U�ƶ�f�Q�E`vp('-e�6��<�
yV���%}�x�-���җkƓ�{����z�����D�ʞ�( t�8��������Scl�t��A�F3��Od�g�w$�?����������������������?O��������ϯ���������������ϯ���������_______���}}}}}}}__\��ϯ���������__\�����������������������>��>>>>>�����������������������ϯ������������������}>������}>�O���Tz��f���یuke��v1�Z}Ya�!OY���c��-oyAog�v�����T{}����U�H9�;Pg�U���J�޴wOqE;�^F�(�]�a�W< h9�ս##_�5�����IF�N��d8������B���MȘͱy��]|�<qKBuT�2����

��רVU�ڂ�۳��X�"ms;Y��e�E9��Cb�m(e\bc��5��IT"�ٷkfv�˚&9��s�WV��U��>ts
wlf9�m����r-�����S6DjD:�=�t.ےȡ��z^���oֲ1�����[���b��u��]�%���3�6��[�e�Ɩ���+�/08ԤU��
���Un��+o:��$Lqy���d��#7�\jZ���@�j�a\1hbĮb��ĝG�j`d�_m^�;+@�=w����+��^GW]F�vu��)�l6+�,sXޭ�i�Xb@��gX�KE��lƵXvTm��ׂ�%sV��ĸ{v�#5n4�/T}���52�HX?i��w{Dq��:�&��vf�(��wy��}L���Ŗ�}�.�������[��I��Z�a��R��q��j�=�u]���q�2	Xt�{��Ĭ��u��
�-Y����E��/���~дJ;�� �uk��wh�\�z䃑=+s&�$&O�?O���������>�����������������������������������������������������������������}}}}y�������}______���������������}}}y���_||}}}}~�__________���������ן______����>���������|>�O�����}>�8k�V �5�/Jb �f˜Yc6:�B�]wߓ�>�5��d\#/t��&�R��]k{x�U:L��*@�<T�#��^Ǻ����7Hh5�v�6&P�͌ts���{��&�`u�J�ǒ�	MaZ5�H&�^��wD��f�+\p��蛪{-w�]h.�5͆pCx+6���u����h��V����)U�]6�M�O:i��2�ܖL�Y�s�2����к��T��Nn
��^;��c���A����Aڶ���4�H�F�$�o����.�=[�/N����\�qO�t�>1*:�֮'����e�[��^�fe���9(:�BR%����gb�qs���]8d�I���R��kjS�������un���-��ᫍYFL ��q����W�Ü�:�*��T�㚃W�qo2�I�[Y�>�d���Dbi��n3*��c>�7��&S�P��+�@:�I�l�7�H��u���-��`�����U�7!CH1�uZ)���ܓ	�qu��b�ܙ3�M�]��o�x�����]����ݘ	Ka3�BL �{,5�[�b���1dgC�}#�º���;�ԩ���c2�l�T\V�8�:Cq|>?�������O����}>�O������>>�����o���}}}}}}}G��������������������}}s��������������������>����>������������ϯ��}}}}}}}}Y������|}}}}}}}}s��ϯ����������ϯ����������ϯ�����o����}�O�����>�O�����-dc&`��(�Sqd;D�T��Ք��\	�4�[�ǹl(�˦��J�Ztn!����t��CֶES�dZ퐟T��IB2PQJ�s6
����1$sU��'ڄ�(>��Y\�ͮJ��R���6r������W@�Y���]pTOS{U��m��S�]4�C��kl�tq�ݺ�h'�.GY��r�D�*�� �Z��o^�`Zq�֝%ݧU�����2��!�(�����i���}msci��gj�\�d�pqػ嶻��_}�֘q�ʻw��w��������}��cj����ٺ^Xa[�ꭸ`±e0�5Y\6xJ�����۪�?}JF�F�a�u��7���η��&��N1y6��C��K,�U���u��� t��R�0�u��進D�c?~[�ݪ
���O7���S+�8+�̙���L��6*)�en��:����#.���h.�z�6��*吠�y��g/���E����e
�X����C,��B�=����,�]7w.B�����;3�hM]�S<�WM�q���v�(��[z��U����aserF5���2�,t���J�e��6�Ʈ��wO��u)�H��S���	c�G
g�������@&x�U��[�Y�*'�}}��GUs׬ݍ��X����͵}m�I;����A�fP�o���ݵLtZ� j�����w�	�|1��έ�u �����|�h�ߥF�Ѭ�*��ܫ\٭�P�/��-Sv>�5�e�W���d�f�jͦ@�U�~��x�M	Ya�j��R�V��n�s�n$���r���7 m�t,�|'+0�+A�cA@��р\�w�v�B��:��E��΂�@�	���4��)�q��A����{�7�(湱�ʾ�Eou�]��Q*����9_g��gj^N��xˤ��b�dx�>�í��5ǡ�BIu���=V�DحĎֿ����hs&L��h��Gl��ά���r`�T{ic��$[��o&�8!��!{��[Ս����W\�t��wQ��Qv�Yi��:���R}��"��Y�:')�j�T�e��!��9Q<��ח��u+� ��=��WB���X@�\L���@�]�"<�꼬�,�Γ̮�����jۣ�/�R��^k����	x*Pѹ���z�>���NQ��+*r���!�y��CU��҇�	�
�8|�a[�p�a
��os;��--K��+�k=VD�+�2���	�7�p���*���z�I��lN���J�aô�:����h�}��)Vl�Z"�.L��BR�P���أ�(��~�P[��:(�՗��k;F�XlV���ՆU����]1��Xwtܵ�X�
�����x���I��Lt�[�� a�Vԥf��*�����,u.;����vˎ��+jcPfVg$v�RX���`��a�j=s."��X���ь�6HX[{@�B�a�+;��!]k]�Zػ0��e�o0>��nl���G4��)�0Ҫ��F�N*�E��",,�����;��h!�F"L
�PN�-U2%�X`(����[Ob/Bg:�n�f"7s4V�ĩ��+]qvs�ٹ�A�h��Nr��X��P�K8��	-.��Z��#}C�KCi6O�9U��?��U5 �(�/0��7պ ���d����J���rL���'�tQL2���챢7�*}o�#7�%�7i�vW7{��ݐ�[F�ܡ�˛�����Đo�K-����C��;㜟X�zU���hlB~�����ٛ�bzAP��*c��F��tP:�WW\*���������җ���1ǻ��Ӿ,�Bw%w2�˭���N���y��e���ȕZ;6�����*,�4��2 ��x�S�M"]㶨wb��1�,��d�»Yi��ۮD���jk��MD���ݶ�{>�2��\"��X63�V#��9F1�}���q��t���Vǖ\��sy3�E��^J!b��F�IO-��Jk#��)�9��x�Ztn�a���;x�dR���Z��KF�<>ƨ?��t��z�Q����eo/-�3\�K�|����uN�:7�ޝ׍#��"M�ƺ�>J�/���R����;�����v�jΥ��;���嶏�(�T���^UaIެ�m��Z���i���6���R�A[AU
�ėY���#a&�I��sVڂ}�j&�V��uq�#:��b�Z�y�ew�C�Y ��݋�ute�<�n�f�]|�[x#�+Q��7K�x�ˇAa��Vf��)s�� �vҜ�5}��P���&�G��܏#����zj��.�3c���+�b��S:�г6�"�E�:QK��������~������#-�KuD�&ssxZ�%�\�[��j��rs���˩nQ��ƶ�� ^�ʃE���������;�(�|	܏����f��W^	Q}����Ww��x�J.q7�P�̶a]��}'tX���sl�Z��z�n�_\��eBn`��.�5�{�{�N`�Be�7���ɟm[���ط��K�5�OZz\y�B��ŕ���ݔ�yN����;O�f�;{g%(.�J��^pSڏC�%��,vF���后R��V�����2����B-�nD��u�̷���z�[s�����J���6�վ)��b���g�J�'\����N��[�!�\�Ro�y��:2���=�n��E�=�U[��DoN{�)d
�ls�Bc&^,t
���ƶ�0RJ��g%�GHQt�t�z&9th� *�W5���RޭH��d۝�w�{�p��c$�i�Y��Z���-��"��������*����UCK�t�Qg6��@�M�T��Zʷ�vԊ�e��p��@pd�F4n�C����YA��V8��kMW�t�CuY��^ƟD�n5���oM�z�X��m�]yr������q��8�YV�L��j�T���_�ʝ��h<�����/6���RwЂ3h���퇷���]��P�NI,/o9��1�0��3�nN�Wa@������:�;0�Pj�y����`��,�긦C�se`90�q�]p�JKs�����+̨�lX3uPx��T&�����j��"��q�չ�0wH��Ǜb=�+��Na�6.(��^�m`��xZ�tg;7Qh��];N7O\�J �)���"cwUc�'�50�E�rܛ��;)3ǥ�D`=ܭ��*k^㬮��!�g����bߍj���|`
Gn�^��{��>�M��vQ�9t$�5�
��}]�ߓ���v����9� �J�����a�����e�ddWiB�.=���_-5(���Wt+� C�J*�
���G�����є��^�v��m�:�=������xi�kS�C�,�6$*��j�n
Mt�l�Y����\��[���np�r��gi�:C�<�l���b��D�L�l�%�z�+M�2�4o�in�5��1n�3M*6�:s�M9rn��VE��=<Q�Xd-��k��6{+F׮Z����q���")Ϯ�V�u`S
�'y1�ֆ9��y��F�<�I|�aF.�7���T��ݪ��R}c��p�Yr��*S2i����J6��<r��ks�B�<H+w G���-&��!4��Vf����bB�N��Z�ܖ���c�7/����:�r(��Y�s�wv��y�y9l���<z��W������\Z�z����v�oj|C]�{�aK��Sw��qM*��8fKo"3l����Y,.QՑ�kݱ�����s$èЗc�Y�Ek�,d=d)i4la��Ѵfee��*x\�[��(Rp��!�qE�Np��n��kSUdܬ
�EN��R��䝘�,sr��nV��
=|)��P�ur�3'g�km�"�^��Bq�O��_7t [�VK��Y:&�l���y��y��q�4V:�;*�n��;��ھ�/I���GjX�R\�K�3�ZsWU��� VR	�f<�c�b�xG;�[Z�&��W1	��tb�x���Wp�p��m���wy�^��2�p�����B��B���jO�<�gp�x���T:N��t�����wֺ���CY��\�%r�߮ØvCW	J�y���6��v�\���e�N��l!���u���_T��vFV��L�.�i��l�(��M������omU�O�{r�7V�4�� �Vy�L�˻�>�Bs�)������F���i^�nbd����e�pg�3����˘J;e�s+F�5`�x�iL㪻�ЕY��0�Pu�/%t����\��}M�9�d��3��6��wS5�ֻ)wq��s�CJR���U�����Ζ~$eWS����f��s�L�,���)�r�*���o�K�3���Z�(�m'woZ�}�ޛ��d?����>��ڈ?�h`�u��5*�8/iAy�[��r=�Y��kE����,BNe%��K���*Q��nWB/������#<+�[��1�&:4�N����z-�Ѷ`,�o'[l�UWw��
G�>����t��.�(\K�ٴ��zi����l�b�WN9:r�{qWk+�q<�(L�����(,H�,}{���&#�:wk��ܺ1mh�L��%*Vͮ����G��~$A ������˯�#ď��!�z	��s0�G'ޢe��HL4�j�a�N��N�2�P4a��bh���)	�X.�(�X�m��(��.��*3J(�01$jG�O�g�?��?��R�۱�V���0����s��&�u��7�!�Z/n��<��.��J�ҌLB3�+�d�Q�m=�bX(^a�Vw�h�)Қ�珞p!7EQ���Z�����߄����So5Y���MEv���s��;ZB[},��J�ұZ���̌�4P���Ą�q�-�{n�in�r;I˨xkd|A�!z��T/
|$Z�U!H�����˲�n;�+*lr�iڠ�rvf�i\����t���)n.1�Al�����#�l�e�va젗U��y��' VÙu�ӔiSGp���g��u�b�8NO.t�l��A34�\�0�vff튾}E�>8�nS����E!c��Hw"�����ةB��T`�Y���z�;yWb���f�g�o��\/��KF�Œ�n.'[chE�.V��Xo�Z	��A>�k���@4�۴����߮>Q�,e(�m�S7hηթb��2�ʿ�䐲6����fˈWb�έ��ؚk7a"g'���1�۝2��V���]�X���CW"N�y�ù� �|*܉ԩ��;\tTC��u�:z�X���{�*��(l�%���ѣn�H�Bo,
�v���m��KT葴ܴHҤ�52J����E�ɔ�Qh&X!�*b~d�ʪJ�T�d�Hn�-6[)6�m�P�Z�I`�$5	���\,����8ۍ"�	P���&8����Ia4�2�m��H�!���0����,�)���(�L�D�D4Qr��C�$�q���:��7nH����^;�Y�n�&;w:�4k��MwbƢ���������������>?��������� �n;���h�'�;$Q'? �� T{��	���.�]ۈ.�8��:�7Yō\u�����Ϗ��������>����j(����]��'Vέ�[Tz6���Oݻ�Q7w�Nn�S��۱l���;oǟ���~�����?��������o<<{��]g̞y��y�v㞏6x�_6���H��^Xu�)���y�KT�Ji�1	䏗Gv��@���!,a�M]�7m]tp�R��JCcEB�ڥ>�v�]cwc��x�m���c���-y���;��Z��<���q��n��$ra��/�2FL&�<�F�<(����m�;P_�0�LI1���Sd��@�v��ۮ��h��������y�LQ����g�q��iػyh;�n<<���Yx�y��bhi�Hs#�����R���*�w��Ƣ��w��u��S��W]�����M�"�NAq��󷗓�o3������j�!�3Z;�����֋���b�:��o<�6��"Ƣ�wc���-&��Z�#���w����A�wn#�GY�:1D>G��.(��*�c]m�zcq��A�4WX��h��;Q���l��ZB�j-�Rjcl�X�P�D�M�
����;l��xk�V�T��W�k�#_�j�������m�L�����ҷ�3��qj�q%Ф�K��su�)���FK ����2+��˻��]u�n1y�lq瞋3K�����v$���I4�+S�𹎯c��Ӳ&��h������y���Tߏ�Ū�5�{�����ޅ�l	}= <�y�=y�v�L�S�}B�n?���S�= t{Ց�u�	>ʸ �ꩳr�i0J~��w�l5~ ��`@i�s�'��Vtk�{v	��'������-�kٱ��U��i�炙��=��&Tc9�C��:�>�?V{����=��8O{����7c��>7ٴuO�k��j�����my)�qC���an�7����~�<�����s�|���'��l���� C�~K�[[�ߡ�M��IT���Y�1���޽����H;�����׌��vXk-���<I����E�B�lѰ~����}������w��<���wd���RζS��U��47���_��(o��%x��<K���+�g;��wO:W@�2(щ�5�hf���.ؖy9W�걎&��~:�������z�4;!L%�X0���woǯF?�Ҽ�w��t�[M�K}�EEݲV��Rg�H���4�)�.ۇHh������f��ج���
��w�RboC��K_ɎTA�}vz��y?,^���3/M>�Z�bz}���}��]�|� ��!�E�L?����`�,Y2���g��o��?o/��keol�9�Ug��:E����.�f#|��^g�b��L^c�ͼ��� o
�k�i}�;
�ӴF��A�Ɯ��׹���T����WG2oXU��V�s������H�;��/������0��Zߟex��^�P��sg��l�x]���\���b�ArH$�%����*�V��o/��/��T����sZ�*�|��v=��Y�qON���k���T��z���^癓j�t�Et�dge_Iھ��U X�y�g f��ࣼ]<(�v�y�����(�3�u�h�5�i��odX�{x�N>wb�Fh8v�Vz�j[��6�.�]��՞����&��5�w�#�\1�Ou:���i뒐p�'Ύ�����6�r�`�[]��b� �����?+�l�u����L�KL1Vp4R�%wp��u�j�2t�X'�T̎Y)���=Uծ�V�<�ls~�<�W��6��y=��.�h<{0�O{w�ן5����G��,{~ULm���}�k��s@~��" �g��F7FdՐ�8��:iy��݈�Jr��󝖌�yJ�riO_���璘�rJ>���1�=*gU=�˼42���G��;�t��-�ʛ��^�{��Cך��=�2��T�{b�Ko�ז��#]���1�E\W�s���d V�k����2{����jw
t9��]Ax~РH¤qO�����ٗ��)��5�y_̸�#B�N�9��+>�*e;דw��h��z�L�?gU�E���3�ƒ�$��v����ˈ�� I�~�[�}��*��_��oY��S5�
�����X=|f��/7�P���I�q�[^sN|q./k}������'M��ž�V���EgA7Ov���]��)��DT&��]&��׷�:3l�
f4(ms�}r�n�V��f�������-ߓU�:�c��R
�]���4�]��u��z�mt,���S��3Hr�-vǚo~-�w`}-�C��^��x��,쬿����[����<;�@�`��[~ԃ��è��+���7�W�9�N����z,��_w����AyC���=��
�īN����I�������8.��}���;��6�k�Fq��9s7��[i�=� �-èzoL�Kx�{���Kӗ�7Säݿ{��3��O;�*�i-�׊
e���E��+��ᕹ]a��(��z*E�8s��G��gXc���~n�l�����k:�[�+���l��n/����*��:P��1T��A��=���Z�߆���[^��yV,�}������l ��t��,u������#���'�m�L�<U�YwG�J��Q|�no��~s�'�L�|�&���tg
������_�����9 w�[�����tG��<^��`!���1�	� >t�ハ5^�<pf��|�WWV[�&��WS�(M���*��:P�me���y�W��:I�=��֢�a/S��հj��h�{�\�����<a܍�M�FDBr�s��7�<��^� �ۛzM�\�v�������XC�� T}\��>�^Q+{��-aiS	T���Ɣ����n(����M���HC�3��ߟ�߈ܤ2�
�2���MN��Y"/_������v������{�S����qo��u�Ƒ�*K+']y^ؿ��_��M���ᡷ3V�9�=�K���Rm���k	�HP�ns��p.E��~-b�� շ���W�QgS�^�߭C�M�����;޸�%�@.Gh�_}sdvtzn�+:�����b��w�M�H��ҩ��5�"�_Ԯ�͞����RZi���M3���W�*w�W�����;4�C�����2�=
9����wA��QzT�����JK�K���|^�CyN��:����%�t ��/�r§�o�u/oO�q���gJY3��ohwýO�)�V͝O�W�$]�*��
�uqz{h>�v k���<�#��d>K��O�=rmS����O�ۛו0Pt�������MA��2����)��,�ݨ>�Ӕ�B��.$�!5�|�LK\��0�߀:Q���Q�(y~w�������D!~Q$2��җ�ZT��呵��)���	]ᶓ���U�+�6���}#�s����:�)������2'�B�e��nIW�;*�������4=�O�d���w{�C�NmA<��~(�AN�J��P�*�py��d�"8�\l
=o����=Ǭ9ݑ��F*��{ו暇gwI|��nlɮ�;��тW��e����}�{�o˨�<W�sv�1{ݬ��j�����_D+�O�ߕQ8hMUK3���9T{�̊� ��2��*��\��NKL`�O��Z0Ѻ
�J��}2�=er�M�U�����n����6��V��@vh�D��#Ev��xxť�o)4?)������&���X�2��MER>�2T�
�0��{|�VC��ipw3E�puƲ�F�{�����/j��g���z���l���s|���^8g��W"T~���k����+~�焙�����g���T�������X��\F��TV�M����W���������yJJ���[T�(���-���=�Ao���Ū���1�F�RHv���X./�'��]N���>/t���;0B��PS�|C�0;�t��L([jOp�t�ٕ8�Ϸ+A�ݮ��ޭ�f�ޡ� �=v�@N��au*��u��d��ﳰ�Z��	��k�Tw�w.����0�8���.vCP=Y�tc���f�U6M���n�+<�⪛��bkĭ��1�|.�Gmzw�2!��O'�/g�ߦ;�y�｀k��ʈ3=WJBU�p{�Y}��<q����8���F��o�&y�~����[]��#��<�y{��7o��{"���M����5<��5����S�����S����u�K�r8�FC^ǥι�oX�1��h���C�=�x��y��k�s�<O�,i��� �\|"�7�~r���I�ju�o�ǵh��ܨ"�	��;/Iܷ�p���롺	��	<z�)�?7���b�������߻�)��k6���5w�#M\���cN}���X/��!Ձ1bz??3�]�z��z<gl��[���rA=ro�����aE�7�M�"�7�U��,x�aZ^{��TG7�.(r�˥z�܏����-� M�}� ���;#�BpU%/&J��1ҏr�1�ծI�vf����,�2ʼ>�ѳZ_1��E�q���L���{����S9d�agi�r��j�I)[s4Ux`�+�r�n��ɇt"ܩ�Ņ�Dm	Q�.�~�z����B��s����;�_t�eH�蜃�*�t�rm=�{y�s������;�A�Qa>V7��~���ϟ�5�˜�S���k�[6�(��r��j��-�>�Y��8~���"�T�r�{�uZ�SX��zo�Bǽ�9���=���KY�B����US����d�!��LDQ���V���ϫ��x����3f��l��k����N*��؝�S�'b����X��u����v�������	��]�6��@l���>�[����a7C��GO�Ĝ���\��q=�,Վ~���^���8&Iͽ��!�CMg
�[FW�r�[+�#T�Ù��-��ϗ�%�)v>��{�Ur��U�`��ڨ�n�����{���V6xʊ9y#��nєܤ��Y;��,Z�a�v��Q�`�`7��BvV��z7�M�{�;�)XaM�Ę{R���`̡Y���:H�\�>��|Z.�S�f�����ss�*x��{��[go���D�
~�$n"�Q9�~*�H*�5}7{K{���%��ӧ��w}�W�{��+�>��~ߜ^󥷩�k��\������;|궫ޓ��Q�`pñ�g<lvz����Yĩ��kȚ�-oF=���jzy
�O�S�8Q�x����y�du��2E�g���i�5^���[�3(\J<=��}���g{L��녯��Q�G����"�׻��W�2��q{�,���|}�;��jDe�^��(,��R��{����{-OҨ�2��6f�*�s���/�2����k׳*�5C��)�.p�
��؊�����ýʉ[=�po��("��.dl6|�C���{sX�Þ��=�}�H�����ֽ���2X̙�^�3z�/l��t���:;�b�O����<�xzw�j�>(���K��U�ؽ���SMX�����I�;�c'��I��+�����Ay�!4��0�R�ˣgA�/I�(����q�M��ѹ�)�u����&gE�>�d�V�,����΀�"ν���)	�\��n�j�QnVң��T�;*�����^�qj��: .&8��4��쿾�y�ǻ`�"D������]�n�>�H<Z(�s8G^��'���azLŎ��=�[V�}ڐ�I[��؀U ���+��z�u���<�uF�F=�LWM���I͝5;��3y9µ�����j���>�y�4�!n{�?)4{ܩ��;�zb��{�ןTܭ5�x+l��+��z�S���Wk����V�:1Dyy�������7�iմ:ɛ�'������VK�6�^W�>>���L3��y�6����i��,@!�j(0�~�f�r�Tu�]�
;�7��||���u�d�����靸=5��8�Y.��u�bI&�N�s�#��fD��t�����+������<��h���9=���2?�Q[�ʟ&PpX^�WO�Wg�?a>-��2��}����"��ϲs+*�\�do�� 0��q��}�>�� �u�\�&��+�-�����=tѪ�Fvr)c�-�D���\���̫)�[K�M�ѕ3�y�Kz��"����a=�p�y�@.��>� Zii��u�y� ��6�����!K\�w|�,R��I���ŻA���������҂ݛ�6���S���W��L���-�K(nY�W��ӧP�Z�wD
%��Jy���戫)[���d`�=�s끎�Ԯ=
nF�2�3f��>*���
r� ����N��i��a*eC��b���׋r�t�-l
�U3*vK]�&1S(���
���.� �V�Z����ӥ��Z[1X]�Fvo���Ƿ2c'�i�)�j݇@�����A�S@R��ώWv
�r��5��=��F'�+v���Kt�17N4�"ܸ05E�VN�TWE�>��[3XF7B+o��z�w�tH=��{��%q��l�Q��Z�1�mѷrģ�
H�+�Ž
I^m���b�3�9�N�r�$ʙz�q�y�&�Yӯ���/�"~��U:��@�g��hu^�w�J��y��Z�����U��T7'|��v����3�>,#���@<Fi��EH��X�h,�n�pN�#z+xw*m�+����l��g��#/�s�;��tJm�܇^w[�X�¨>-���/LRe�!��<����dR/X:�*Q�ӣS3qt�d���ۗ�!�F��,5m��mfݼLF�Q��5/7`��.�;|Y�u�]kq��vp՜M7�[)��N���Z�,�8m'v��Ϫ��B�뜳#�v��s���y�w���v�Ÿ(�O�<6���O�p%�N�l��u����b�D���8w_<GC�2䙹�S�^@t�e��"��1e�#=�ܷh��s�c5s\E�D+*Z#��
b5���-�	��v���*37_Kp�K�,>+�v�M��c�aݸiZ�RX��g|�Y�&��:��z
��l�,�{�Z���+��Q��E�#�个"���/m%���Nw[`�GF_^�����pX�uo|�����<{F3��lui��40�h<y��8ȴӥ�btMH�/�����L����{���C���&	���B"���*�3����f�"mq��wn�b��j�T�5��s�6�0���7}6��Xx�ÚŻT^V󏳺�1N6�F�ҩS�(�;,e�O��5HR���:���Ub��Su�Ҹ��15;��ԫV��N�D�,�,ufS��򚤐�� �i��f�ڇ�;��k6�vFYu*Z/;Y8���#w�,��ҙ��^,����P�96��d�W�����opb
�Ƨ2�ۻ��+,2N-�#ᙤE���w(�b7ҟ`�A�u7o�����|(<�w"h�&�͋9��5|��G�Oeeu�E6��Va����o�����J&tV��Eh�Jj$�:�bf((��ut�"]~�o�>?�������~3���|~>u�Ah�N�7A����l�j��kf�m:���i"&�m]8�5�;��~����~ߏ���}g����{����`�5_;��'�M�hkcd�(�6*���h���������~?��?��ヸ�)��4EZs���UpmV�TT��ђ-�TN�ן/6�h�ڊ��i�q�(�kl�h��=b�j�j��f"J��Ξj��T���(65U5�(�I�hɱ��(�kN"֢(�tEl��"-i���V���Iε�m�h�`�E5��&�UTZ�DS�S��ѭ�f�N,F,mF"�tDla���QD�%DѫS�k$A�f��"�"����F'Q�`��Q�kjMj����G۳llj�ZZ��3Y�U5j��6u��[(f���\�̏�i'I��Q��늒�p�[�ٻ\���4U�`Le������_�����[���W�v� xO�)��K��aёe�� �Pn�S���3����`��͑c��\-ξLf�m�PƘ�^�ဆBl�`+���f`1h̠�4ϱ��t���PĦˁ�h�WP��9yrj=Ц��2`����w����E�w���m �~�`���������`#��]��P�ae��0V��h��VL�P�������z��������p"�(�o�@8�u/�h������Vy���;��(ٺo"�.n�h�{��@�����5ݑ�y��ڞT��Ph�R-�Q�L.sx��2�r�x��ރW	����t��B��Ӏi�Ck!�d
d݊� e�����m ���!��:	�#��" �qg���b����6R �ط���#�z۹�:��P'7�R)�
�.^��!����ʨ��S9i��B@��#�����3,�l��f�f5����A�M-r����uP������M�K�i�=ʛYsQ��O<?��M����
8��f���vE�,��s&8�Rp7s�P<�j���"�8yh�ZSqp�(On0�-Fc����>��ܙ���E��t?�����&Qt���5�n��⋛��,�t����^�t���U��n_���}�"pR=[)L�Ǵ�����U�v���3��B�Q��g�<W��I�w��{5[��%�J�v���y4(r��+	 �"w��-4�IV�s��Įu��2��Ɉ;.$赜ƨ?|~��7��f��;��Ž:��C'�6߹e45+aO�ǲ'ܪ)��X�')��H��xO1�\W�]1K�W���s�ޏ�w���y?�W������ 0�������j��eu�|�$����ߵ���z�3;����dU��0�g��P��~�]��y�+��˿=&�8OҰ�6!��~�����b��hc�y�S���S�]�{?�GT��O���ס�kH�m���l���ҥx{��S>k�6�M���>�j��}Ϧe��G�ޯA�.5f�cKU2�P�dA�[:������DG:��z���-P/0�W)��g��f��������Q��I��>n�.��١_�U�t�u�'U����I�@&&��a؟M�_e���'����d~�o�0{;DڽV�2{�t/����3N��E�J��;�m}C��8��?+�S'�@S��Ĳ�[7�H5���� 'j�(�����Zk�	�m��.��)��7����O�T>9w��b�Vzx���ii���?i�M��bo �a4a[պ[���1I��YB����]1>݋�KŊ�:�STX]p��4)��8#�����xi}.V!u�iq�3��;��f������z���)R����:�T=6�^l���;��9��C�:�;Ȋ�gx)�%��h�ls�m`�΂[�����s���I�U���CcW�j4�(���#��G��� 2�6���6�_C�"ƑM"[O�oߟ�G~}����*���ɍcB�$���<�k�yO�nEg[�.�c����ة�ca�[{���h4[z4��;$�3��H�aZū��u�o��Q�
�͊�S�`�sqAx�����1s7S��w�q>��"J�i�!��6�ъ�K�#����x�	׻.9�m��X���${���ړ7��͖���ɗ?z\��z�<�'QBs���6��;���@��XO��Kq|*Ty����	J��hi�ٹ}���>`�¸͍��R�=��Zf�;�-�^Sȼ�pɗr�sH�d�9�a�#U����"�C	�{�;��^ϧ�׼�bJ���j��r�&`�X��@�4+�I�ׅ�\'��	q���|��u�Wܪ�UR�l�,���(f��4@c����!�9��O�X{�R���/qi��b�A���&b�4�����7����"tLO��P���Zo��1�*u��Ϡj<���<�{����q+����j^1���&��T��ߒ'��}��3ʄG�K
��6��x#*{��ؘ�ˊ�EvVœ�~}�j*>�y�A�\vt�y\4×�婽w�)�����F�n�X���*�ď�~���9Id��śo����O��a�C�p��.�ʮ��?[�:X�>�W�!���G�G���~���o0� �ͦƍ��jd�Kc!� ����,��f��-^~�gt��˿�|�dD(��BC�lr'�'�����N8�����;F�r}f�!�GB��	N0i�4О�f\Ј��c:'���hy�[v7�m%{5�!�xME��}Ɔ�hq�e��A������-���L0��e�T.��7���wh�$����<~���/�G��}Tl�x?��K(V;>�n���.̪{$��x���mA�*K	6l����4:�_1����i
m�uKꦓ�Ĳ��b���B0P�2��k{�܉�s�o����>cϝ魦��
�����j��kbz�L��s"���Ɛ7��Ĳ�[T�'�b\���>�h��Z�s����uqA�=��eD���.�!�}-!�tsn)}6�4\zC�t�=?D�L-���M6��V�r��蜛�֢����ߨ�\gA<H�\���w�~5��tBc�dգa�҇G�qv/)��tsqP���Ҡv۞�S��<&,��Re�@���2Xw���4ӵ?[�*Q����L� �\���	tp:�ܯ��g�������=���cz�ӳmv^�ދ��g{�6'�$N��$9ha7ttǬK�zf\��8g��hԧ������/�U�|�^R길F�řQ�rv�u��̎�.�O?�Xz.��q��.��4�j�4����Ɇ�n0<�a�*s�h����Ǝ�W��� ���C��_��b���1�f��'%�T)����jN�v:���e�z��̽�7�F�{�?����o����"��,���<�6�Ɉ�Hd�=94�[�l�������%������G�y�t�CM.�k���-�X�ӱ9���v\EF1- s�{M\p%xm�Biԋ�l�����y��z2����F��~~#��>ڿ~j�o�2f� ԫ��O�����-���`-^����Z�ʽ�37/��3��nL�A��<`=7�l�C�^؃lsCO����4c�e��X��t�CH�a(���`�-�O�D�b`W��E����!�$3�xi��U4�_�}��F��E��U��3=�7���œ�2]�^�o!�n�G?k�O�
���-�Co|�S��_�Y�9��ǔ�4�U�"��뵭��{�p�S��Jfׯ���;gXH��N�^�����?�*w5�?���I�����͂�$z]�A<]�^�-B�K&�+*�R�ƭ�������i�h�	{g�-#�k�T�3n�㓨�7�Y�m�CrIo-��t3m3����'*IZ�oFI�sca��
o^7L�+]��x^K}qĵ��C�ˑ͊�n6ۻ3UI��,%�.zـ2���5zݬp���C�i�}n3�R�f�ĶD�#4b�ZF� o��_z�
��Վ[��������+:GW���\E;�~��߱H��Nc݀T�l�k���E�:v4����O���[�ٱm�B9K���j5��<���4�z4(�NNj�{\މ��9w~��O����?^>�{Xs]��k�R�	��������'�A�%��O��}���}���mpw��I�c����Ԯg^ds�����C���=t������K�>���Y ^���M>��v��%�r��N�I�5ЎY�G!�m̿�̄!E{	[C:`s�}m�&���0��@��P�'-y�"ݜ�FJ��X�6K����[!��e�	��5 ���[%���B)�_ݷb44Q�$B�.�EC:��&�cF�Ӛ�G�m��z��Ȍ�C�Qa��4'ߗ��ϏmOl�>����l,��_]��I�ֵ+|�"-��(xn���}�-B\,�zO1�F�t�9#C�t�ړZ�LP�<�ғ�AJ�����N�+���K/;�\~N� 93�BC���d{�5X�{�2:��S�0Xc�I�:ٷy��������1Bc]'�~��L/0�]��/������̟���)ʙ��;�A��������wE߷Xw��Q���[�'�W��sU^��;�Sn�FE���*�F�uv8C��w��Nz.��(y~m4����w	��3lu�59�t�6��P	k)�'j�9��/>GC�hr�+X�۱�}wv�ѭj(�"$R8���������� �$r�����+�$SA$C�|�}<��&]�4�q�-^"��<������@��M"8����/ӏ�Z�瑝��+�c�8�y��fC6��8�,���G3HJ��EC�6(�y�k0*�$�w���=w1�LAͤ����qm��W�e�\�^��k��k]���Ừ�zNT{Kȉ|mg�:�t�s*X���^[�/��	3�T����e�������^[Ɏ��+l#Z��ox��/�W��C����3�n�{���14[d�έ�.bZ��O"�5���67s�Z��QI�Ȭomل��l��

�\�]�P�o!�pp-�cM�5�)�V9f�S�����j�i6Ƒ�¡�ҳ٘cE)^�0��_u��G3(i79.��F��z�ճ5�~�c��^@�꽙����Ϫ?�My��e׼"ۧ3;����L���l�g,m�3y1\��`=|hP��K�Ļ�w\m$���߄�����(~�ۻ4<���^�&�	����z�X��A)[�@J�����۽<F�ML�6�G*��5 =7/L�^�<�ȹF=B�q�$v��_4Y-�@�O���e��j���-�W���{-�>w�1�>Z*=��=�z��8]r�A�Vؼ)�T7��04��.�u>�����CtIJ�y \ɔvK:;7Wl��T��`
��LoZ͉�����*�Û�%m�f���vdַlwn[��j��u��aYX�)ǟͳ���__0�8�8o +�x�B��{Y������0K���G��ػ�&eY�t�j;�e�%�jF����Z;�[dkrهΏڈ=�ȃD+�}�(����|��)���ow?�qh������Ec�Vfay}Msނ�^x�F�i�lSBz;�`BTy��~��9Xag���ܕ�(7tɫ�m�� ���s��k]x��x�OT�B %���'|�:�}��5g��/�ۯG�w�%��TS�[�U!������ŧ�n���	q��%t���B��l���k�P��'Pq��9��;`����Ä���mq�]ônG'�nr7��bBSl�KB|��O�� ۳"#8Tfs8� �{K���l�(&������C3��Le�#	�͵�H��]{zr�T�<�e�X5W2��㻇ǵ�>���ϥc�_/%F�z�5O-�S-m��O��UNi�
���i�������&`g?�u�Ugf�ˁC����������{����e� 9���)����"�<�z�X�c�ɥ��:F������
��Sj�%��-f(��f��*<cLX�b&0�۝fɭS�L��*�핀�H�S�_K2�	�J�&�Ӕj;x���ر�Ѱ�K��+�:�G~���x�U����Q�Ρ!��v�wrnDvu8���.�s���TL�2a'9���h�ڜ�^�?S?A�Xm�?����|�[���5P��7�,ЕS"�4��7�6�J�>5#5�Tw����9ec\�WYSc��Q{;%x&�N����ݐ�4���酏#�I��4�*������g"��%��ꠢɪo�ʃ�%s<a�x�\����P��C &�,�Ω\����5<c��O����|
����U�-����_v��������������\�m~ǆ8-IoJ؊����A/��	Y��^�y��ױ���0m�.�9�$���B�:���'�	-=�A}<h��z�饖5�ٷ��};�Դ/.��Q��Kc(-�T�c<�����͐͞��(�	y�MR�����u�c�`�ћ�o[)x]�c-�T��s�}�ם�AS�%5K�� t��-w�S������Iv�R!��"�Nj
�1����='�6lAO{�}���"2���I5,��C����D3j���O�zܰ�u��|`��#�8e�l��U�7@�֠�\��cnK����1a�����-e��z���xf�]45	9%�\aQ�͇s(;nٗ�k{B�<v��V�?0�0>������8���)Rd����f�(�\�/h��x�h�P��ݝ�h#ٷ��:!J�&�*�P��s�]^���M�`��xNp�}M��+�P6.��76�3%�Y��G4"!��-�\�aĎ}~�|��'�0,2�0~��@����2h�)�����3U�˾���X��?#�4�_�}��!w3��K]v�U5�̣ӷwY��z��r��N���]?�ܩ-��LMG��o�(��ME0%��_%p��r�A�oj3g��3�G�܇���ǌ0���sM��j.�~0��9�#��Dp�T���O�*w��J�.�����V�,�����ǯ�1i�ɗ+�l�*d��s�v��&e�w�	]��o�x��q��<������%z*qu쁭VvBm�wE7�$���ޛN�`K\���݂����
szR��ͱ{����͜�<�b����C��G�1����5A�_|TZrsU�V�uGlFT����ȁ\��e�F0�)�� �7�m�3`}\������.��9�|A�b�yĻ���[�z$�\�8MOֽƻ̋����<�ĵ{z܈�q?�3�x���
��O���lo��Q�˙yT�7��>8׼V����|Q,SG������;�?�lSyG��4�6=^�i^ë��>c���.��X�=�SenK;�l�����#����/�wb35��3+6�':�4�9B�j�9FىmD2�f�}���N��:�U�77�oVW}q�t���h.�������;��df��&�y�=��j�7���alw-�C�yc�5�l��e�s=D_d	�r �Y6-��xu\5֩��Ԉ�̭s�K �`=K�aξ��9I����j�u�Oepp��S�.��]ˠF�O��3S
������{5�x|��L[�F�u��ř�2
�L.yu}��\��a�5T�)�n����ְ��n�j���fl�f�r��2�����
�C���gC:��m;����.+� �Q[��bG�����w���N�(r���ی��YU�$�Z��ʂ5ٻ�����!���l��|e��G�N��V�|ѫ8���W�a�*�]D�mWR}�<�`���
5��͒�g�rfI9<�F�X��R�(���v�U��B�6A��f��-9�gK?qT9CUjoG �Gv�32���u���5���Ǵ�̽�b�hgm�Bj�b;ٲ���QA3��u�ggrc:���<�u���B��9/s�N�v��|�wVh!Ғ}5��P���U�,��ѷB�(��9�Q�6�j��38��E�~����㤜/.Ú�=V�(�����U�<9��ѹ(������ѷ�#J�sр��4��\-�	��	�}�V�x-_l���Q^bﭟ��(v=�nҢ�f��}�'>����h��|ģ9put�IًpY����hQ�&�4!�9�)�&���ф�yA�V,���YE�}��ͥ���QK���}�vz�۝Ou��h������3���&�αw�'kwHO�@֘w��	�u
��H��s-�w��i�d�%�4��}���p�7��~qL���:���^���-\�^'˞p� ��d�rڱ�e��4[��]X/���hN�Y#;�i�t�����unCv�K�g�Z�C	"��T�#��t5�R�qY��E�y��;���;B��,��K�N�3N�D�)Sw7G�WLW��[�sE��L��D:�(�1�(SלzWnvُ;�9��*=;��7�L�ܣJ@넧�"��^G���Y���[��ƚ{is�^C�R�k��Z�l�������_E&Қ]lse��+d��?t��W9P�%u|�[�s'i3�åϙX��Eb�;����D����X&v�k��d���X��:]������n���pN��\a@Ԧ�f�E�wt���	��2T8�X˺��f�����Dn�.`���b�Op�z����!�X+��wI��j>��һ�*[��<=b�9���j-�M-fgl\빧�74�.�p[�o��zU���E%��a�ĂWVؾ읒;@������ζY���jm���mM�CJ�;iû��]td��;Ȇ8	*��]�R]��kFwu'��k�wlF��Y}��i��gU�HM�E ~��"�GR��
C���a26�U��b��L+N�L�̀ F!@�r�d��/;W���~����Tm��U3��4��[-b�ƭ���_ן����~߷�}���������j�#2��Q|v3V��T��FM:�Z1m�������1��ǟ����~߷����Y��~?���Y����*��h���o�c�[�:kAQ�G�������?o���~?���������AN�kF�:��T�6�-h��*�SC'F�#�]�:6��5����)�Q���l���MQ����(�AF�5LA��Mv�����Pj�E�SUc�i-a�PX�h��,�9��R:b��Q�B�ژ߻���EKhǻE߽�A�1����6űm�(�ƪ#gA���#mL�j-UuVڊ�6���EA1m�J"*#`��mV ��[m��j��Fڤ��&d�-f�&�+�DM�����(т&�F���X����������M�=3f���2���7G<^� .�tچ�f�;Ʋ
ͳ��Aeb��ónK�/5��oZ��u��Y����#!%��5
 �Te��&B�B)!@��2�d��?��a�e<�X���*�xr�g��e2�k�) ���i�ʭ�����^��7�gg�B�Ϟ�O�/X�~ʔB.[L����)$��O.fA�5�Y��5	pp�{���F�&iap��ܨȶ!gH��&��K-1j)��`K���l�U���.ր/%ĻD��s�F��.����j��A����hwy�m���������\�!���خC�ױ>W�%�+_0�]��*�Yy��{v|սY�Y������DF�z�h^>́��H˵���KQ�������T�����-۳�/J��Z2'��i�L���K�oBA�.���"-�R��y���ty���OB��2j�x�������G�u/EŵwH�.ѻ����F46��B�鈯���2�rNcD��}[W:� B���J[%Խ4���+{�A�0�f)>���E�kSVX��i֥j����_�/��=�À�����ϟ�J;���:jl�˞�(��?F�=<]��ۈB落��	\�u��\�
�v;�h����`0^���سJ�b���I��h~�ܺ��� c-����[�n�LVƔ�Jz *>���hX+�=�2��F��9Z�=n�	�����}[-ⳅ��L����7p��O�Ya��QyY�jT�nyg�8��W��]s�9�*�f̔�kk��۱Q���bEe�J^�w���"��0� C ���y/�����F�;�ǻ�������|��^���SO��@��O�P�'꜐Cqf�����V�t��mNC��s�NK<��ԣ�k��͓�70����ޝ�.vŘ1j4ۙ��ۻV8t�j�M�/)�z3фý��-���*S �(4[��q�kCH���xK�4T���o�Ǝ���/�^�	���4���w�N�9Jy�JNKCܢ�a���j�u�6�ކUFԻ:w��a�m�1��6�P�L��/M
��F_����O����}�s�Bz�@��Zr'v�g<uިa�����;�1�������H���g�IoH'x��5FC�u�K8{%S�����[�����=CL�:��ă�Pl}���a0����%�o:U�k	�{���uGCح[bM,d2�py�oz��T'�x�����H,#�@8�:2".0��ם]ޛ��9����pt�E�V�;���n�����vĪ�S��/�2�y/ؚ��#�c�S����������8���%��&ޚ;#[ɵ�lt��`���4�3M	��<J�ɇ9�ǫ+���s٦�>*H&�{�Όt�.v�i���`�l^���.d͓sdM��/F�ˬ�X��6����-�p]@��î���H2����:������c�| �\H�8�g9T΁8�Y�X��w>y�7]G�w���?|�>�=�{������0#�`0��[���WW����y���s�c%;�;�xz�=6w5���w�?�"��#25����NQ���*0a�������Π�'�@_� ����L�i��m�V�Zڅ�	�xq[�Ϋ ;eZ�����5n>���~��2}}��u���͖d�M	���y����w�}L�ꬫt�yC�Tr�@.���^�Ye��>{��%�ܿ-�9U��%"�O�w�r�t�^w�(��I�sBD�q�5y
	к��a0.�T�GA��
~�<�Z�k��خ����uL1���Mt]_7���$(���[�,��_�y�����(���u����2�[i��uW��q3w�n5G!-�3�G�l�kT� �5������5���m={�-������`���������:K��vO�������2�-������*�?Yqp�l$�ô(ɚ�$�-ֺ�y �B�tX���_���$3�phLsxG�!6��L�ڂ��IF3���ݛ�N�.m�6�A/��!B�ӈ\�oQpͽ!�hh�m��Ey��9�3���"���t������M�f�YSa�	r�Ȼ�R˄9/�ʮ���f��E_1a���p������ENQ����k5"0�]��M�Ywx�����C��ގO���#bHb�ɇ혋Q������K{������(��U�N���������|�������f���ʓv�1�,��z��q|gx�G��:|�ÿ�z�ٿu�N�v<ִ�D[��u��B]��z���A�O�ꖳ|R��G���������e�P�՚9̝�@�!�Y���]0�a@��Ѫm/y��9g/����lۺE�xk��J~��'�f����d�,C�'3o��j!��؇n�xf�n��CB�-�\aQX��s$9|������rg ��Mj���I;O[����p�,�ZbL�*�2�^�d��ُ�����f�x��ʙȝ��ݎNЗH6�����v(���W*K~(=V@������Q뾶8�*�P�M;���U0����0��B3~N��-��>ߑڂ �;m�_�5����]٩�}y�v�]�7A7�Sb��Fc�k���U� ɫ޵ɶ�)m�v��X����7(ו���������ri��z�C��З[ClDO8���v�<���5�9ok-QI��M�E�и�DEB��/y��(�r�,�m�h�1MmP��m{#�)�F��Py�?I���E�&^�Ww�h�U�\���m�:�ݽ�7��S]�W=eC��ոfl,���+#k�FM�Vwp�5��j�դo�ғ�:��:Lg7ݓ�a�[�k�;�WJ�]%��R�Ih�]%��9�x���kv#�;��r����H��h�����>��y��w�v���!�X` 0���ox �m�!��%g<���׬�L�qt���/��#�z���_�axC��K��?-�|K�qF^��C=&��n��.�͆�Htl.���yH:�,[C�Ү�4��/��g\�.Cs[7��F66w5�J�K�.�2_�S��εi�E�2�r0��پ	�o����H���]ʫ�;��v{/�k=��-����3`Kg�Gk�e�iOa#%����}����N�$<�t��F~���s��cs�T�����yN�ا�y�EP�TXm��hOV�|�C�z���y� D�����̂�}�/n3���e~c��9�:e	�T��1X�y�F�>�$��쎒��� �=�*�y�����:b���K	�pD�ݛT&��nm��,��a۹�u�$�.S�xw���ʣ�9A6����&5�Tq�hW�5��M?SS��a����R>�� �����'��k��)z8��> s�⠱����t�a��,]�?���3ʉ�v��.�{c�g�j�Z+�ԴӠu��5��g�f���̕L3���WD;�C���7{s��Ʉ)J2���Z�����/YWZeM�7"S�-YY���e��Z�N��Ah��u?��C�?��ŋjJo�����o���ވ%����-u0�����Ի1�)���W�G��/?�D�FaG�S������&aq�ǆ�qM~���R��K�Fm�2%�t\;�M��w�Ċ�7e��9�Z��O+�#��3��]��7%�)驅�[�^l�ee�bU"n��.�E���U�XK/��y��.N�c��_��_/|��w��%66��1�;�ebnU�;ʎ�@t�Ie&.�V�*M�;j��om=����t�Yş�]h�y�y�'+O<������/�{��_=xnW�,X���z��;�i�����F�m�N �V3�������W���?�����>�q�e���j�t7D��ȡ�.^]�c$�>+Ւ��z��˩��#{M^��ܞ��	���8�o	=R��ኔ�at�my)Z�(憣��J���r�ڵo!��6�󧈦�ih���@-��)�l�4C�uj�e���	 �(9�`�KBEcL�v뷺���@s�f����θwt�����P��T�3�ç�3�y�����~�c���߇zx��ܘ,��;�&7��	�|�ʄ�~U?,|G��i�Gy��yjxG�x��+D��;'3�	-� -�8�r�rr�Έ�Rs�{g�4j@�̖�4P�9�U�ˠ���O���9��-�Up�k�^��k�2��Y��딇��c8�7z�cA諏[�g9�Ɣ�S�K��Y�ukc|b#Ą�~D��������|�>����;�o���O�V�5H�CZx�4�]�oHx�w�р�	�-��W����]y�>��6@W�I������{ӎEBzA?{�"=_��w������>sbz���fe��J�U:�ΘXkm�_g���8����=٥+���5,�,�(�=��k��y�L��щJ��_/��M�|���+&�;j�$�*w�K�gxH�!)�w��3CqVbxd�Z������K��F�@�9�����������u�k�,e�:�.���H�r�KV�Ov�6�*:���0�W�a�k����}��S�:==�*�5�]����9�Z�@�
h]�"�D���R��F��K��M��1m�(�g�q�q#������r5�u��3+ŵ�)�%��[C���R�of���b�ض�k�P������溴�+�IZ��1cDq����`&��hxL'�e2ԦYs�ylEec
S����ƊN\v�P�SݕO�ʁhD�z�4xZ�5A�nx.�hJ�7v%Vܲ-�̆�6osG��r�4��X�z`�UFr��JS�|g��8e�|9��73r�,��������C���'���4����`�7pY��1��Q2�SW�kU� ������_
��$��c�P�1i�"j"�V�^��*����2�C!�
�aAq����5ૅ�r��ڃ[P��v	���M���0C�R�
���1�Z4F&�2��c�W9�h��Tډ��Z�E��1[�!?�`mŦ�3�L��ӛ��FD!����U"���l���v_�_:��Qg��(���0���w$�2������T�oֽ�����I����-�.�i��]EQ��c!@w�3�!�w�1��/����_yO�Ъ�(���Թ�&�����^Y4��U��`ʟ>X5�H����5�&�v�;!�#��0N�w�l��_`sg"�^�!�w���;�`,tl����>��{".:'�7�Z�urmz��9f^R�!5:�>���	��9�^�>1�R4wF0�B�1�׾�U�s,͂`��dM_U�b���9��$��4*ɖx��ߤ=ӄTV�6�����4�U��ؚ�r�Q��ܯD�o11E�x�K�qii/�f~��&w�����g~��_��eK4*_V]�o,�f��j�{̑G���ި�S�9�থ��Qc��O��GX�/Ĭ�s\(���Զ_�آb���mJR����W�f��5F�j)��S\f�uV����.����L�]f�z�E�?ϔ�K�|D5lY�Q�m=�SN+�Sr(��b�ةܕ:5�n��ޡs�
Y�J4*�����0� �H2ҌwW� ?�ȉ�����ߟ_l9�4���랩g�qL�`�0�M���lS'�}5�,^�͏�D��]�$r�I_r��'��2��?	^����������^��Mt&<;�n�@J{"�a��>�d٠�ާ�K(USp�ف��&�I>?)��O�_��������0C藚ӈk��:��
Йs�(���H��$`Ѕ���U��=���/vd�X�˵��^���K��߃E(�1Gs��R��p�[a�Y��;#2CY��T�hχz����cW��:����cSO���\s5�l�p�F��0���"����~���`�M��P1�Q�bz�CH=��n�3�w���xd���IT[�S�7��ꈙ�T�ݎ�:D�v�s�c˾v=�@}��H�q����>͖˵�-l��u��tr�U΄�2� w���8�������	�rFK$�=�cE6P��wg+ok\C�n�n�^�K��a�6�}#����� t��e���-��)}2*���-��69�=[>�Q���O�6o��?g.����|8#k䰚>`�RO�B\j1YދN�0,gs�N5#"�T��{��e���n��[e;#�MtOf-F99��`W]����[D�&�am@&�ڽ�]:��_9N�����>L�8���A��D~7�6���E*�t!chw�g{+�*8�H�
VU-)��b��Y��٬�w.��c�{힭�֠ϝ�o��  C�<� ` ���@~���o�?���?;���>�'��Έ�^D,$9��$o��>�����+�CZbs2z��-w�C[���r�K0����1Bc���N��_0�x�I ���
�\~��V�잷y�ҙ��>�6�h���"q)���'�yw�����dFT��S��k�2����V+`�`mOx�*��.����f�<Ds2U!���:�����3�缋u�_����CY�|�����qMA��=�͗pX������Se��}�w�G%y*����}M	��;5�����P����0&�,�n��)�4�*V=C����'�J��mOU�Y���2�h�EA����W����+F��e٘Ht4m������sW��[��x�p�-�9��b-�ί��'���M��n���zeԝ��kz���v��/\ߝ���;%M����͓��M��ޙ-��J|������Y�B�\�[㸬��d�S�]���3չH[�ۖ���"�Z���6]��3*0���9=i�e�q)�ʳ�6�:k6��O�z|=�x ׹���M'�)0l�m�$�kT�A��{ju��6��Ï<Д��vwq�n%:�|���*���$�U�u�;��7t�����;M֧k����R�I��6J�ΑpŖ�[|��w|N�uΤ�b��k�9N�M��p�Ƨ0,�s��.wA&�5}Y��_R��XɆ��2D7h�:Z&u�:�\pω�cG5��m�����G�cB7v���Q�!�Y�AE�� 1�Ji��P7���v]�`8'�E꠯hR�P2��2�Y��ϴE��gwz��]��>���p�u�c�W�	o�e[�ۭ^�t��i7�BoG<�ы{�.>���5|�R�9���X`��l��#��,.p�6U�6�s]F���\�N�	ӖM咣�@qj5����t�`lv�l����!���4�-�Dr�#���pWQg�b=�:h��	��w��n���Ak�?mӭxc+MlYȩ�{�k�5��ۤ��D]�7�ܹ��ďZ����H΅+�g_ݸ��k����$b�۽�+�F
�����������)2�c���U�/x������<�E"un����E��\4.#w�T��qo.��wI�3���u�{/-t��v�bV)A�qđ�δF(��dy�/�H�N\��G�՜��,��3��o�`N�J[1*l����c�WPcr�)�� �����|�2�Ƈ�3~�MHr$�[D�*w�`���D܈+F�l�rۧ�:<�0d��'J��<�n7���%�S-
�t�i�Cޮ�W*fR��ٸDa��b�7�@�!+s�����'�]�L� ��{k���n
�j'��3�u.��\R�>E�5V]�ޡ���ʻ"�u�D�Օ�T+\�c�ZS�'�}��������l�j�e>���ŏC�=P_+�5vtZH��`�.�%���7wE�L|���G"���֛
�e�:����K����G0�W��%N�����}���9�ʸ���/�ft֕�kxò+'YՒd�5��c��a��(Hg	C���Р򎕋!��a,��LA����FJܬT2ʠVn��M��o�S��M{�ÝZ�.j�Ҭ*�2�l�l;�E��kQ�$�VO��R���2��A�gr���,��8�2i`'!BL�+d\������fT�Fч��[-rz�C|��O�D������[F�o\',�կR��l���ba�Ż��P�;�xB��뭓[��7&m�%bTmھ �R�f��Or����x�6��l5���r�4�HI��o۹��ow'j�l,C�Sh��2��ٹ��n(�WӰD��3 ���d����J~$�H6�UF�b*��"�*�U,lf���?�<�?O�������������~8붡�����kPp9u4tf�d�(������51����Uf�?���?o���~?��������tԕ��֊�cTj���E��5�Zӊ
u�c��DPPy����������o���~?�������b6q��1ML�ۀ�#�/ͧ�b������Z-���(��%D�i�ڿph��	�:���jDo��G8�-�cf""�:"�6�Q������cm����h��V-2V����1���Z�*)��U�Mq�Dlj����ѭ�UC^G]AQb5S��$1Sڧ�N�;[V1;62ULU��ت����mh#F���b����[X�&�*�6�DTT�`���%1b	)�lkU_;uD�m��8��[�4ch���55k�����jkv;��{g���!��cf���P-�L�{/1S�I[4*�Sw��3�(�iX���o�����P�eV(�`o{�{�]<�7���=K��ױ�E�!�̦L���f������+\o�	����Z��,�吱�����.��.l8M���y/9��yF�8�Jy�%��"1��s��m+�\���y��׵��ÍJ���	j6�����1@Teĥ}7��2"�ʤ+��<���qh�����c��]�z^���3'��3��܁m0�N�d]��wWݯJNϙ�^0V�@A�ln�>=����0���t_�~� �Mp"��>�O��~&^jm�>ʍ�����^j5_g�b�Ϳt�BkH)8�q�k�L�F=OT{�"=��Z������������f5BUh,�V�sܻ'��s֧F�9GX�*���~�O^�R�E\����vɶ�9Aj�VϏ� {m��)f4����*�8��h���Zl.~;_���^;�cA��7MW"��bZ-�L>��MC!��F�N����E�0�k,e7���v�hR�]�C��7��
w���9�	Ó�_0;�xЈq�~�G���Jd�|��3�/���r�WrkYJf��;���V�}���J۝�<�y��x�IV_oE�ν�`J(k�&(�0	E3u�}C�z9
6�v��y.x:3na��]����\?�zE�Ɵ����E�f��	�`q�/�7�wm���>a�<y����y��ޘ��x��X~;pJi��&l&�Y"m�Z.6(W���9is��|l0*�6Q���b�;2����ݻ�m�z�6���u�V���,^��+Jm��#uB�,�T��3.}�n�^V�7&��'��Y�i�{!y���H�g-���b	U2/��J�����c&���d3G����U��[����Ѓ�p4ԋ���k�?G��ֶEvtC2���y.��'�M��g�q;�j��*-�b�:�\Kzm��rl3�D�.�|#�&�p���?{T�qO�x�J��f���9갩�>���v��ǌ���d�=5ʀ���w�����'����xc>�<�ׁ]��S�
��o8���B�4�ۨ�\���Q��[�֡�Wڇ�'�$�;ڵp>��[9L8�t�U]
��*D���`/�'Q�*8�|�/�w�2��@��Tx�}�w����,JT���c��F�hhmef���������o�nOc������&ʣ��޶�NR�p�����$<���r��1^Ǵ�S66y>���_���t'f�|���,\�5D.Wim���E�F� z����)�ܕ!ʟZp52�E���RM'k��W\�f�Ĥ��μ�2Ɨr�U�l;�f�c�J;yV��A���Tඤ�;�˹�'�)��R4��w@�ڸc���].
���2��]o����rM���]�,��ٝoN-Ǳ��lFĉ0
m6HI���߇�0��X`R��U������{��+��� &[�B2A�\��>M"y�>"��y���Xp���4jr��yo���(�I�'�7Nz_�T���@�&��z�'>a����5�
����"���U�1��h�785�~ܴ�C�drL_��Bj��	EԺz�����P*�3'��G%��VkM}�旔L	��}�^� 'Z��̳3cg��.�t�a�)[σ��9ٵO���(�g1�?��zJ���c��o������5�lz���^��Bf�Ԣ_���3�鑺���j��;�ejU��<���s ��P�h��[�W�-@Y�b�?rɖ�[�*I��1)r�a�w3{Ua8=�~�5�f����!T�T{�Be���/bV=�Z��S��V��z�3w2�{u܊�Ƕ�wVE
݋c5�8/Ml�C���h�N(�p��G�P>0���������P�٫l�W���`	¨^pɌ`�[��K��=��°��9}��ȶi�,L�C.Qu]�uN���A�78��c}���~��1���P�g��FwHɯF0ts��}��?%,v}u�y���>�ꥹ�r�ɺ�ރO�ǥ�|��ڵ[G�)�ȝ=F\���Q<��ӅBŠ��J�k���-ա����X��]J�D"�f���zu��N2V�f��Lf��w�����c��=�{�ʋ�� �,<�xx����v:H�:�*�@�/�j�]���Ry�1�$b��ʹGlo�i�YB�x�-���{?f���~�>����ݰM��@f����Weϙ5�d�Lc���w���n�ҟ)�u��Y�$��%��L�#�9���8}xdV��F��[>�=[&�j�{V�vV|��|��c�Y� Jɟ����U�:�ֳ�|5���4����z+�L����=|�7k��&��<��ͅ�6�yݛ#��]�@�e!�[�?�AsKO�kZl7�d膘m���b�vC!�|LϽ��s\X�1�Eٴ�x�:�_0�x�Y��;���;��0�.��a!�ٻ ���K�����}�|��Oz}��n��W(���cK�Z^0���vk�5��e��䰘��I��ޖf�},�c�69�"٫��$��yřp����*]���iK�3
m�9R&2
x<ۊk���
a����[�����΅6���s
x^�&�p3�À�~�Ѓ�k%��147~�_��b�R��@J��!�?)n1�k���5��|��s�l��'
YG�cҸ��p#������$M�BQ늜}(3�h��Ti�Ք�'t�)6&�v�`D��D�|eNb}�Z�?��M<�]�5W�!�{�����nL�Ɍ�9k�"a��3��������������q��?��� 8e��7��o{�x�M���eB�P��{�T���n��2H��P�w.O�w����C��	&{�Y�0fd���﷥�s���tk.|/)��,����8��,�ax�˴�oF�[L?I�츕�{٠��
h��R�P
q��aH�I�R=>D߱X�u�s~nW�:��� ;3��tm9~�Ս�Z��۵4J�P����`;�(P�:`��yeϼ��Vn����T�-]�k������Ô473���A�Z%�=Kאu�c\�;!�2�H�-���g�7?�-��NI��ؓQ�ߖ�]]�y�=,Ǯ��������6�)�՚f�a���Dڮ`���� !������H7٪��9� '������6M +�BY,ҫ���0��g�����5�U�ӜM���W�1e��W���D��zJ;�e�����ε \��q�����:�/S1��a�-�%Yǋ��<��{o��n*���CZ�΋��A�Oɍ-w�R�J��. 7�].����p�ȫM��aϟ �t⊌k���1�UH�B]�����f�c���	43�zP얟t���b*��YF�
im-{r#l�ш�Hj�>3�t������G-a�D�v���!l�{�sk��N_�p��q�qxrS|��z�K?�OwIV���:�!<�W7Ci��Nթ���/�P�FOЕ0	�| ���6�p5F��D��"2>/R�_O��S34W5,��h.)����֙�f���(��{Vpv5�*���c�3���������'�y�{�؎ �31w�M.O�4w��?���JWK�8V���;d$/8����M�:�����P�ER�(5�|���w�v!��`��lJ��y��SyK�E�_��l@w�����]�FF���@�D��ׅY_�*ݶw|*�56A
����ף�c��hoit�q�D��`&�K(V:�x�"���-m�����E��.=���m��0Lo!���F,x�b���e�՘��iN7��Y�.�,��ڽ�}I��D|�|�X\ڙ�i��*_ �0C��Fh��3��2�n����٠��`��2�S�gSv�b�u�5� �j/���� D��l,|����_�A��酂�SwS:�<�d9Gs�8��-���q1P��qm2�m%C�y�LM�p_t�\q��]��j9�8/-�`�]|��x�Rz���'��*V��>arl����M�:�&}�{��}N��ul�i>�0���c滶��p<k��k���lU����ȷN�'Tp	��&�R��p������y'@̥yV =�WG�/,5#y�o].S��u���R�R�%�}���׫�Pa#��u�t��f�����_r��ڷ�3:j��t���֦����nn�����G� y�A!DDox��x���%ď�-����������*��"�U���u˭B����-��z��Ld��s�R�Xo{D�֝�2ލ���"&�^,l��R���ƚw�WS^{��P*:<��8џ	j��cA���^��_���n�^yN̟��R)���Λy�~�In�&�g��,�;T�5��T�1��vDJ��?i������B��b"~�R�H���C��,Z�m�?�$����M4�w��o�r�ʮ��Yؼ��h}j;k�tN?ǟ�}�#��*}j
;�[fy�yP:"6Eu����a��u�Ev�v��̓�`C:�d��.0��c�>Q�ьc��ŵ'm�u�7l�;<�g�y)��aNj]=xs˾� I��_&d��ks{�(>�����Қ��3��.���[�;PFm�2�-�����WP��ٵ3��)����v
UUVi�Kx�2���&��N��
T׳��Ƅe6��ZQ�d�a<��/�^�yj��z�DPs�S�Ժ���AQ�n���_�O���g��u��bYS�Y2۔�zCc������MS��#-�{�b���Wʟe�]&��9�:�6��4_$+4����+ph�4?5%h�.���A'���`9�[�^�;|��'a�H-O+OdD7;J7wg6v.���'���{�|Q���"a�ds <��xx]�9<)�C�)����s\�+7�<Д>�Ŋ�`��ػ��k����C)�k�>ˎ�&\��Sm9������KW�!� o�4�B`�4u������&��5zv��版����^s&�lBQ93���,�a�ʢ���z�[?�
����d��iDd�ҭ�c�"�(fEHf��2�|�#b)?n$ޡ�*��ۓu'��4c�DA2[�M���u�K�d�o~�Ƹ�.ף�uB�:�s�g�����G,T��/���kb�)y�,4��%��З��q��&�E���P��z���r�5�%���}sA��L��R�j�ڬ{Zܶ� ����}�ҿ�D���H5�Y��^�}��z�Vs�-�cY������>ڞO��U�t/j�%yλ�8�6~���]��_�������x��ߞ��#Lǚys���b��ʭN�[�������0п��=Z`���^D-"q�+Kπ���H��߁3�y�D�j/y���k"v	���Ɓ�x���xWʟT�������C]�WkE{Xi|E͆��9��J�;�$!�-���oٖ�ph׮y
�4+���8��+H��E�k��;Æ��N#��㵰T�[kt|�o���l�Ͼ�}�&��^rX�W&����!�.\�o ,�c��������ʤ�yA�1�;}�;�Y����t�� ` !���a����< ��{�V�Hg�qT���[�[f{>��8�a�0��&E�J��^��g��(��o�6��ϺwׯB�|,�l��"�q��+�钲��8�� ,���r٩��G<�Kp�(e�x���Oܵx���q� �T<�
c��%�����N6�;n\3PܡЭ����g�J|��܅��3��	���z\����蟰���R���Hy��0�j��P�u��_�Y�ю��hǠ�#�\&���&�U8ՐPq4��"��9?f�??%�r��^�y�)?G��"�-�;h��9{�-�����<x���M��Զ�͝�Ws��̨a7��4[{i���L�٫附tZ�g
�3Ed��6��2�ڑ�$�h7�bB���;
��'E�g����rf�����1B2��4z�����lG'�q�E��*�R̻�޶���b��k�냷0�\e�;�@��<��.}�t^��<��#L�=�.�q}�E�4qgޠ�V���t������Og��	��8��w]"mL��X�Iy��"Ga�.?PE��OONc0����1�����w]���AnӨ��t\���y;<�`5r�r��4��i�N��O�ͼ��^�cV����*���^n���
E2.�X]p��NYҜ���%�r�}`��f�}p޺ᄀ�ݧȪ���ן^������?���E��g�"y����0o{��⒉�z�3y����Ǟ�����G>�6�T�T��Y�����!m�|��0����~u����[�s�{	�gHŽ��8��l�{�PK��RXO���^D��\X�+���_TP�����R��c�倛?�x�g�>�ޟ\^���-@j�/���q�h�]�oKö���OW�{W��wk��l|D/��r��y��uw�h�>7Cޜ�9&�H�\X�c��/%s�q�շ��Mb�����(?<�Q�?XVz0gצ�66�b�WrO�1�ta�u�`��n��Wv-e�/�*ZҌ��~o��k��<��G�H�����拠ڹ
2re���-Iې�G���}�,��zQ*�ѭQ&r|B?|�d�Y��q<�5e���w}���8!&vq��^�`�^ℋ�}7�\����cG}IÀ�/��?N�.��6�}~g�VPy��,��E6�3�L1Z˓!7�}�P�V>�PL��jT��lٙ��	��Y�Z���O�~hBMc�~��y5Qm9�X�Κe�)�zVl^)�H~��jj_�uO8ϕ��흝�|���po,���V��uƦ&�>�w>;/t��V5va�n)�͆0�N	!j��:�s�ȯj[ؖ�Ő.c��":��ۦ�-����{s�$�Ø�N�\�+'!���"�+���1�QуX�<˖-����\�k��c2v�7R���f��K�1V���$���Y�u��C��$�q
l�<�F���f�LD�3�#.g'Y�LOv^̰C�j�	2m�u��fڻ.�:ixͷ�C(v-+w)[�eo&��Y(��]:IE�!���E��o��j
�����4�M���1�z*�cK�p�.\��h�;�e�_^�V륚�s#8�&�f���r��Q;�W��A�xƪ*4��O6�7�{����l	9�[M��Fem��>O����J�ؿ�\!u�G3F�7��ۚ��!�@�+{(�I?��T����r:X�d�5<�>��1��	��V���ֲ�j
H��3��v\�hY��rЖ	��&�%8'vef�j\C^`_.%ݭԖ�F�М�����J�6��(v���͊�?ǁt_��A��_>h������Tp���d"wiH6&�yP���13��IetI��!�Q����{Lĵ�3���N(u[w-ÑQ��fi7�>bM�XyJXP\M��v�b�t:;�����5|��Fj[�{$��V��ݩ2qY�/8���$˷m펅	6�ZX�ԍ�U�M�b�B���H%�.�	��(�ȑ�Z��d�����;�7)��Q"�V�gG<[Y΁K��m赢�YT�7E���x�+U	R��0��1[8������kor�jIV�0��u. ���A+C>i+Z6>�h̢ɒ1c2%�k�[�p��$2�plsW׎���b�a���H�͸V�i�M[��� �ݨ���#`}>��8��	<K���,�������V�.6�D�ڒ�c���v��挾�(P�fʫՆ�9���Yƍ���Y�T2�CT���%��T!�߆��
hα���_7�v��S7�Z�vVv�3���u�x�63C��p�	���3u�vpLk�L���6��)m���i_Z��\י���,�
d�B����e�y�3I��38ˑZ��2�+a�*��<ŭ��փ�L��>��ݎ��k%��\WON���àG[���v�V�7�E�%�q[�^jcO���ȡ��oS��vG�����s�k(vh۷�4��`)�i��=���u���êl�q2��T�۔��y���R��8�ӏPb}kb�����)��m�p�[�o@:��ħp�P�{\�pG�VjW
�ۚ�pѺ/��&�	$�vh r��4��h���Ǥt���e9/���U�Fr��N�עl���+2�r=rV���-G���k(_w,ƙ(��9MP"f��	��L@�)���b(U,�) ��$ULȚ�E"q���:<�͵�ݏ�(��TQ��Ehű����}�qU�������KL�s��>?���~�_��������~;�:�hѭ�A0�y�Z��4SU5E�&�4kLF��[bbH��O�Ǟ|���~?�������{�h�΃EEQ1���"
��GmD7cTA_�<��?o���~?���������э��
���Q���&�ѥ����b6������OI�"�h��sAlꔡ�)�l�ɠ���MF�����)*��u���Z�ݜ�q8�Mm�TPZ�V�h���c5�4;*������آ��b��&������tL5DS51T��EUkAD�QDQ�ED:3���DWZ)�(��W��	�cME:�QAUi5UL�QV΀�md�ET�T�Q�bq1��
��h���B6�QM;�m~w�ǞZ�7l[$�u�C���w�Lp^�oF�M�VT$���I���_h�h�:RqA2�=��QDb�c�sB���5�)}���~!@��	'�i�K�Iwmݭ�(}��20&!��A T^l�W=u��������߈�'�;�\�6����W��y�b�t�dR�e�qE6��)�V�myN�k]Z��l`���i���x��p�H� &�z�Gq���j=y�����7�����;���x^�g�Se�M[m��}ޖr� �!���DB�;����C�Ğ��hT؋}�����P��A�9}�R|m
�i)Z��*����g���O�^��ד�{IH=�,s�*zU5/q�oMޓb,<����pj����F75�w���6�<f�ò������ka��gЅ��ޟ��C�����T7��)���p�	���5�n�Ίy���fq�����OjD�0���QJa3��E6�ޚj�R�qG3��Yv�1�v�����ME�N\���]�ԝ��6�Y2�������^|-�<�24�cg��2-��L��v��za��a�q�6w[�+z�'�K���\l���dQ�$C�0*B�/C��#V4��w.ifk5����AnfǮ�B�Fd6����T�t
"m�"埃����r��A�[�&�i1�P��d�M�,��=��[��87����ęYd�W9r�f ���N���j���}�����A�@U
 
�^ҏ�r+�5&��|�m��`
����,�7i��:�{V��2���*�S�`�x�~�?;�������	 F�O��\`�)o�&j�3�J���pZ�p�>����k�ť��5�ߓ3h}�������s�j�x����mV��&��v�ۑ�Pш��� ưƐ����'.�vn�V���<&fi�DB�&�>�oS�t.zQ隊a�Z=u�,^(M&nt����.������fl-{-d.�[�����5e��AT�F�F7�Y��B��y1j�.�V�v<�D�!��w�F�ޟi(U�m2�>�<�y���	愯�������W֞ݛ��N`�ɷMp���ۨ�ۮ1I���E6��1�;�V}0��G��E�3�ö�?C��F����]���)�37�[r���Z�:b��)�����*���v=S�{a�4x�}�v&�7O\'��n�����a3E�hT���F��b�E'��U�j�����S^���ʶ��bޅ�|��>�بE�>0Zg�+�#��N��A%�c�[h$v��A#Sh�(���HS��a���	����|��t�k$N{��l� t�v\��'Č�u�1�m�a}g�'��/n�<[���>�i�p#}1vn^çk|�C1%�Lni9Y�T�s7����h���ַ*%��
�7�
�����b�}�P�+n��Ų1�r+z�����$�6��)cΕ���L}�PaP�|Ʈ��`�9i1[�C�:��"���5��=,=�� <���ox;y�{����s_�Ty3�g��.gO��+��$���,?=�QO/��R�^����c��IR���~p��v8�ӗLisu�;>������=3��y���#P0��uW˺��A���Q��YSS�,�+�iFE���"6G��?�L󲼼H:p$N2��?�j����g�F��X����,ޡͯ�[���Ǡ~��g�xS�t��������sߪ��s��ݛ� h� ʯS?o֨@��"6z�����g/�-��{��KWDSBx��d�p�21����o�/W���.�9=0������_�����-�M�Ztͯ<Ds7H^%���I�*̔:MWr�MC�6�hS��g�H���ڂ\������-A�����6:���]=�+����ւ���]ހ*rO�T�:�?��#"��L`f��枘d�^�glER���17(ӡ�����M����Kh�s<�L;hjj�vp����>y�l������w��5}Q�ѷt�}4[��-{N��o��#J��ce�
݋e46q����C�nn_�nv/ń���.��]�;�����/8}�cl3"�˼%�]�{�hk�x������h���h��Vj[�b���ht�v�6���[k&.P��B��c�_H�gJRƮe�vB�&�u�jv��Z�I}����C�`a�$ �㾾|/ԢӊP�C���[�43���:D�锟p%>D߱,�6�۲;Uɗ���ϖ�2gwy��|[��h{��q�'� ����}�g���˟��Ho6�ҞTt���lf��b�g���F5(V_�?j���R��K�@�_Ja=�%���2�.{k���|=�}F�P&SjP�ƈQ�1���" t��8i�ۂ`&�|h/���u�a���n�Yֈ��F\,�4�YFKP	?��0�Qg��`�"����X���Q�����a��ss�dކ�:��*�W�K��Z��U��=ύ�D�B�Z��oKǆ��g��B��;%,����+�S1�᡺�$��U�A{��4���l&r� �O_L-�e���?,��_�����R��q/ؖ����3͖c���MHQ�{,��O�cV5f�{��{�'w?�@F��̎{��,"�[vS�;-��`_3��*������-m�a?�֚[P����c ��@��<�C��S�.�($�na��ڱg�[�:9�,,���qu��Ͷ[tCS,7ΞC��BA���[P�[�C�d�g95�C�ici���i���x-��.��	���/�m "5��i�o-3Me���׉�
��Z�:݆�I��Ɲ/ڰA/7^o-( C�a�]~v�,1�o��_�9�`��I�Hn!��g�?Am�$[y�)�>g�fi�=�}xv��L:�XP����U\m�6�a
��Q�}�^�T_���E�c�@�M�}Q�ccG�\9_=�QT��}�?���e�-f��{�G
q�N%][aQ:��i�g�6�Em���;vF*����i�{[9؄��U�a(~h[�&X@f�0M���T)��P���bYe��c{h%�b���t��l���t](�#�yd��׬|y�׼�W��_z��]��f����*<l��lsy�In�sl7^��/^C��w4ԋ�!�J�<���=�6ız�5�]�|U �EZ��j6���[�%��&i��N2��Gk)x�2ʲ���������Kh�#kB�g.�ax�}1x�*x���"��5�%�EJ��sJp�7�3�����+�⧞�g�D,ӏ�M�B�v,��
����vHV�7��L���G(d�˘��}J1���;����i�ָS��C���T�a�(�M�1�-N���E��n`�F�٬I��L�h+q�Z	�Y��^eNsWc���%}4�F�']KYS�;+��Gku�$����S���c�v��5G2��H�$�g�]���ǁߕ��g���I��#c0��9ܚ��b��{)�\�`ξA
N��:���)���T��ם�'�#!�¦a?~�7����1��c8��>�#�%�{�N�^Y��>�馭�J�k�Z!ez��uĪy����M��2��v�s�lm�25���<��W���\wʱP%z�7����&%>�u_U�qW;Nk����vD]	�Hީh~j�k@��|�9��|F)�'���^�KJ����jBY�fgb�곌�21���,�b����+<����T!�m҉���K�%��Ӎ=]Jۡ��ȩ�o.�d�//�7�z�Xc������T�p�a��lT<4�ygM�&�����i�:�s�	�B�9�&1�d{�E�;F�v�a�e�[H��=R��od�.k!j����^w��(�"�����(��j�*=T��m(�H��s1x�c���a(���c�F�.��Z��h�9T�3֡�:�$�V�埭���b���G�P䲜_�ٶ�r��(�zƓ�=ЋK�r��ynP����s��mo�st I��+�c�`�w �j�*��~w�޾7k�{R~�b�M���=�*q����i��4p{��o�WS����Q���&e�~s%�{7�+bRY%�t`P��.�s�*��gU�V���Kp;�Y��y�c��@{yT���c��A����$�%GUg0RS�Sh�s"ܬ�W�J#"qve�����si�q���<��.�mt؉�mh�z��龖�WU��(����#� �p����GVsBU�����>�y�s=饯���bgب^,�a����eA��@U��������q�ߌ���kx����29�q v�Y�h�����4b������i
�P�7"�n�e�Ukt��w�|���&���l��LCs@��Y5����uJ� ���*L������3���Wx|?45$l�4d���3��h�'O��͘V�N��˔ɴ^�9�.i�3��N[�ٙx �;~M�B���Q��$ZX�	��/�������q��s�/�]��9ҫ�f�,-i�О�l��r�i��TW��Z��a7�`�����}��	�F�iUF�����IT	t�Z[���A���i��tQ���AӉ��;�>���P��*���PP��l�֤cwF��~�o^&9�T��P��s�i�1I�Nfb����Op�A���:en�eͿ�ۺk���]猎)\��r��;o��5F5�%���.���PBs����48����/�U4_췼�,}�������e5upK߰�U�n���f�i][(�$�غoXW�i�o���{3�R�����.S��*��wR�ҍ��o�����P�.��H<����WX���Q�<�!j�h�&�^J�����N��Y��`Se�ސ\[X��w%��y�>��W�y��K{�<���� ��S�,y���<�z@��%Eӟ�9�����_���?|�M���w��2��`#MO<6+-RU�Wq�ϼcYˁ�����tƣ=����.���Uf�Ct��k���bqܧ�;�k��$}DsUJ�p>k�?��WB��V���Q���>g��ܟ��ӌ62_��u��H[�j@tby0�xMm[����tƘӛ��INc��YP�G�v�|��kv�C��/��V�ڞ�syVƴ�u��b�*-�n�H��2��y)�&�+f�u�r,l��c�0�5n΍mE���ߘ�Hl���x��2���Z�C��V6>�[�G�]�;���M:�ml��������O`9�|�.6^^}�Ŗ��_�"��gL�1�V<�{��:F�
���a� ��-\���݆9�BR��(v��kּ��>���o>�K�V/"��-;Ķ\be5ZA���)�2Y,s=�)�[�ͮ��Y8�P���{z���\�X�o��]���~UQw�b��:qGa��1��~'���k��]�C�̛C��-?���i�@n�����Z��M��Л ��j����߳+�62��[����C���K������on��ք2�p�x�	��~��S�%�}9���k�b�$��W��lPS��P��GQ�֌��c9��'C��)o*��>�yߚ����yc�o?�?���B�����ޙ��V%��+�e�DL��f\�����!�<5�_�6Kz}�yX�>X��`��P�;΋?�m^�M�J+�z����0i��1�ʐ�:�8���^ɣ���^���w������ðz�,	-�Wc)��A{�	v�d;:}f�xy���������HQ�?o��gQ�GiG����{�kP�gG�[4���+�J�)�W~��~�?za��Cg`��lymrφ,&�k���$s�e�֛_���A���a��+��c�؉h�� 2*��;i|��u4�E�dӫ���:���,e�ܡ��#'�-�����7�N��W�^߯u��W]�me�.9�|*)y�B�n�V�)�����P�{]�"q\�;�7QۯU�yo���퓽5����mA��s�775�d���t��f%�ZU������񏒶ȹ��������R�=��-ٗ;5�۽5���{�5-�s�xwD&YI�f���tM(:.��R-\�<�ω�,+�E���g��Ís�qt$�D���[�<��$5��P1��o�&܁�L�H�B�5��,��<k|���+��w�;5�i�w"��Y�V�Y��9�__M-Z��>��<MV��^o�w1L�3z��5ǫn�r��S��A��%�j��ȼ�N��,����`ۚ���^F�Xz��R'�x���0�x0�{�� <�� f�-�S%%���s�>���I�Ц�U�6g�M�Lz(�>���*]��M��Y�:�LN%`��5(;.=!�vO?�?)���S�$��|T�~hN�ǠV��s�9�m�#2�5O̤�g�Pǆ�P[�g�/4�J���u˯�dn�rN;��[�{Ht.	�>fn���#�Yq�^	�z�^_`Z�-;x��,QXS����g��&;7=TS�ݳ��X�B�@c��o~*׸��$O��VS��QC�c�P�)���3�t�N�����1���់;���xƏ�����ށC�"�%���c�y���pe���y�ʻ7�֮�3��[���}q�W�"�zTꅮ48#����X�_>?�k~��g����+�-|�)=~����d_���P��8�����_�t�s_f������ ���z�d��~a:������5˻���j�"?
��Zo}c���C}[��������Cd�H��(���_.--/4(�^ߌ������׿Q�+�36��Pt�~^���r����F�ބk��iJ�C��"Y�Mi�2��u�典��'��fl���HLj��(��h����%���e�#e���5��S �:�"ٕ���X����V9/�A�fp�=&�AT�]�=;zn���I�%��������TT^��aH����vL�!:$^n��HÚ�0�>N�MfpC��.�|�:n���ڭtfw6��cj�k��p��[v�nơ*�=x��hy9��n�J����O�R��N����݅hN�[���2�7���e�-��z�sKd�C��y��
��o>䥊�����j�-wig��d��I^����"��A�����n�x�J��0@{�}g�~ciT4r�|�LGo�c�8��5���w��r�WQ�n����{��9�wCtԼѫVKd<�2��ٝ�N�Һ�քZX�#E�	�krv�!#�h�(��2Q�+����S����)zg�S��sw}%�=�+.��Cy�lt����(��ȕd7�[r|⢬R��}\����Z�)�;����c�����k��S9�#���'/���t���T2r�0P�<$�ɐ�V\��u���H|FO�f�Nfoҥ]��弼���l�_n B�Y�QF��X��@V4�S.�ɋ1M��zC����t��.��n��v*`k8$�hzu�p�@�s1�o��-��2J��\�H�
J�SE.�d��㸄���� �m�[_��а4�0�3KH�Z��Q�j���pWۀS۠�.�OTb�C��$��T��{k���w��^��wz�m��SAt��,��$�,�����`P�í�6Z��#-e���B!�e�nZ��۟' 2��RjG������"�˰��i�;TEܢN�67/���٠��$w�����w�v�&c�*^���O��Z�P����Pk�vgv��ʉ��L��ѥ;9w;w�0ɇ�o5��YHaJPb�;):�0�_<�\s���+��W:N���e��L*�[�ح:.Pՙ��`M���ZW2W���)a�#s%�!���h{�#}�;�Qp�jea)Μ(Ŏ�g6��Q6��oJ"Ka1��>0w-�.���W`I�I��/��{�C8S�kT�F�G�[���YZ�e��UϝY�j*�^QS�TKk0a(�w83��	v��:]���,;���2��Q�AO�[�"%�T�U�n���|K���b���]��.7`Gh�(6h�v�DԸ�#��ܛ�r�v���Up`�c�3���2�����cx��MЩ&i���-r}�+)����fP��yR#��L,T����2�E�!n��7CX�mk��6�0�$�v�n��L��.�� ʌ}��s����`�mV����%Av����KSY�o<8�"�*"���ECK~g0��&�G��8�
Ѫb�_�����o���}~?l?�����c��ږ"&"	4���U%Ec��j�?����?o����~?l?����1T%=8�ي;m?�Z �b-�$EDh��(~?������o����~�����u���"ֈ�����]i(����)Ӭc!�j"*�&�Ulb��b�������*#cPljt�"�Z4bN�'ԝA���4�W�Ɗ��"))�:�A���z�ET�T�l[
�75��f*i"J)J���E�k��փ_[�o��LC}X6#�n��A��UULV�k�&N�1W�j#�� ��UUhЄ�b��m�h�����IADIMUDT[&��$�t�4h4j�cZ����و�(�
����l���9W�U��'mp��LCXצM�g*�]�=Wro�b�������y��C�V` � �������ϗ�� N��������К�L���<��L׫���1xF1ؑQ�S�
���t��wr��$o���Ew<mى_�VO�b+b�Ɨ�P*};7���&b����Q,��3L��s-�䲅bSr��R��P�����E/�1�o݃�������οZ��C���y�$��)?_�H���*��Y�|�V������f<oq�Y㗉�}����)�Q$M�?b�����O���(���7+�*�����r9[Oq��|��yq���`�M��}
?[�l����g�wf�ˠ�zO�ҡ�>Vr��^=�3��bZw����Y����!�ɔCY��az=	t�}nz]5�C�]������M��2ZM�jݺ镻j�W���fxف�R,:B88kܮ/�z�	��A����ް%���.((K��E��=)�>�����$XKa|����X ����݆�E���vEֶ��Wo]�gP�;�sxm��hOB�Ϥ[{��H9L~���<��C��fx�/*��W�A�WwZ,�?�bC�'�v.��*�of�_*3E<�����4�L$97�GWݍ��vaf*:�BYO `����(�M�1�� ��b��6��x��xp�q9��F����O�B0�^w5�(f��Uq��P���X �-di��<���|��U����\����s�y����]pS�)��H}�&���tW�yt��',q�9�`�TX���N�5lվи̕����㴽�v*;�PXeB�N(&9�r~dN���}��۹��W9nHSQ��0y5��_��H�։������o�m��.��dXe�����i}���W=���w��?y�/U(��P�s����#��|��G>U�ݐ��>5���'?�}�o�h��Z�)f.�N3P3t�*��Ϳ8�������ϒ�B��=���ٛr����-	�nE���v�0�I�w�[��þ{��8���1��{`1R*�E����p�=D��f��I�e�#n�z`q�8y1��fm%t+N5y��LC��z�5��:{�1�L(F��y��]
5�����sϢ��x/綠7a1�1I����U��6��V'�f6+�Vnu�v�A����C�q)�4��bٱ�9�'�	L	�b���S����u��e���Zw\�p1ߚڄ�2[ͷjq�2��g�}�6�<��2S�X�"��}�p"��k�w�j��`Ɩ�SZ��r�`��x�t�Kנb�cH]�0�����$]�fW��=/GiU2O_�Ԙ���.��������:[���ҙ`�|GQk޾�����e��s(�j8�o-���v��~�GuK�	�J\2A�qV�S�����@��	�Ґ����P<*�_I�=��"�,�z�����M��y�N��w!5O�Y����p?r�_~�-e��2j�}u�m1�Lo]_T�w>)��O6�R��zsA�О�/���W��O���ڥ�gҴq�
Ⱦ�r������C�H�Γ.(�U�,��.T����_��Q4���ЕЕR�#^� �1���{`Y4*�v�4��a��(���0�	Ja!{�����@�6�<A��O2��{��n5z����2}��Bf4�	yd������U��i��Z��>�P���
�u�M�k@�w�i!�Ͱ�H����ɳъ'Y��r
�ps����?~J6R~V�g�����u��D~�	ߖ�h�?z~
^yTG�O��E��Ɖᣡ���S��$���nA?H���S2U)�sR�靟d@�C"!F-�Vħ)![�3!Hn�+'D��@7���`N8,���IO̝�o%x�9� ���J/�]�ꏕ$��q�²�ޝ��6�9��]+Zn���ʀ��E4��̱� ڊp�3g�n\<r��7/��3�=�>K�T�י�],���Z�ST;7z�_�r���B����-�5���(s���#3"� �����#]^z���8L���o�E��Z���lxq��N.��2C�.�2nj��Z�X�U�l�Z+�|>���uJ��ݸW��O�i����ㆢ)��~l�a4<s�Rm�6pG(R���y�W��O�ʩ�)���C�9��4��ٟ�t��QB�1ނ��3����"_�F%��XG����m���D�Zh��?����o�%L�CtK�S
w-��Jh�жvfl���L�l
����B�ֵ�HՈTȽ�3mֲr|�
��W���P�R.�e�X��>?aV��cU楕O�XL�3.y�z~�.�X�R��Um��Z�f-�Íg�D[$��VD�ERy�뛱cgL�H�2i3d<�N�3�~3����O�a(��*V�4'ǜeF�}�8Hw��-��p���4S�D`��ҌA{j��1{gn�S���dA*t��:��F��Q�~�=��Fd��ZU�wB�x|q����lBn�'��]�`ʼ)�i�n�:��Q�ء߫:�j���۰�Ц��~���0}^`��	�b�?>�/�,�,������C-Ӝ0m�DK��}Lf�z���1�y
&�5��p���4��<���
�x��j�X�7�*V&WǗֈ4�Ȥ��E]e���B4^D(=˘Cn�O��:,v4Tn��+4���0�ev8�Fڮ�0F���i7�e\S��\4�M��T����U)���&pH]
`Z3�t����EW)Z�PUԚ��y����:=�=}uꯐ�7����/m�M���~,c����N��oHZ�@pG"q����+�Y���f�:�{���w�m�h��x�s��O���ˠæ��*��2��׍~�t#Rv���p[V38�!�S�8��\^���A���N,����n"s�����내`�Q"E�)�����ٗ������Io3Z����J�(��{�̚��)��X��4{s%�F,���aL其x��Gs��`4��;xw9��YQ��W����>��@�Є?S���ɲ�l�g�Y����Y�e4:�����Euqm|8��rz&�Q�_{A�����#.&b��\���.�nӫ'j�C�Rn]'��=7��^|��ɬ�d�@%�Lm-�U�Sp�y�����܉�/�Zr�4���1���j�HS���D�{�˟�}�R)�ڔ�=`NC�Ǹu�����P䊶,���G��my툕R�>�=F1��)�qC�*V�N���B���p��a��"���r5ݭ<u���噜;���Y�J=a�>��3_@f��N�`r1`�����;�h���A��9K�K�/T�>��sh��vU��c4Oc,�L���j��VHX����7/�B��V�Kge���7���������þS�<��;k�	Mgf:�<��5Mk:�{�}�/���p�8��r��n-�dG�g��R�kG�� 8o]�
�6�+����9�WaxC�#��L�b����"i�D�wT�sZz:$/�L_��-��Q�;s�sg�#���jIm�����=�_d_�rg����� ���
�����N�f��su&��|)���g����9ṣ�Q�ȶG�Ɗl��wl��Q�>�众EՐ��n�:�>�F�~JEW�޴ó�؞�l��r�i#CS�x#�`�,��w�>�O�U��!������40�a�e��Fr�K���$�C-t�F��Z�LS�j;8��$�=�]|� ���'ҿ|3���t���ۣ�_�斟���p�
ήg�9�<[,�
9�.�z^k��z���Ht�ݚ���P��m�]䪜�fNYI�W�S���S1�,��\éB�`��~�	��~�K"8����`_��UڄXE�6������uIp�Afׯrl�� q��Tt��C�����x��Zz���� ��zǷ��~R�L!j�i��ಗ�a�T�At�%}-�;*6�C��ŋ0�Pgo�5�W�9ZmL����16�2�NW1��"�W�3�4����j��])kԥ)�=�'��ݻn\9RB6-SEA�g �D%���0�U7wA�i�}�#!�#(i�e��g�톲���n����I���P�>� ;�Ix��f���G�y�q۫���F����]�r��W�ɾ9(�H�%��:�I/�
_)枘@�oW�Cza6�WB��D;�g�]�4��稿s1�>ѷ��w%� �/h��>ׄ��7`.y�a�O�1exm%9�/I������C��v�9����7ٵ�8ޚ��Ӳq9fRN�4���=�%>�S�I��9�j��P���e��r
ݡ^&��g7�bhn���=�ǁ�~`�q9�u۪������Oݔ�81L��
�l�9q��f�b����w��*�e�82�隨`m��=Wg���+�� �b�-5)��y���-�ոt�YV��	��tO����#��z��&���m\�����"Gb���j���f�%����cX���EШ�A�����]�ٗ�LjhмW�z^��q>���.r����+�I�ge��Q��-),$b��̓����p���_��&�uLU~}xQ ��iu���cK�C(��]e���z���c����𧎆h�x�KhEV^O�G:��g��t^*�zƓ�aQ����~zo��~0?��g|��ڵ�F/߈c�w"�]M�+O�9^6Kͻ*7.��{h�0�:g�y�X��8���yWw��R�J�x�om����x�ڼ����� �ٱ<;.7P�O����y{hmi!S�i����[m�kѻ��4��|�8*`��������§xW;���6������Q����5ǚl�z�����Їn�:6�vmztdO�oӅ�>���n���y�h}M�K�N�_��ﲸ>�r達|=�n��3���3�a�@�r@��5U�����e�KT���b�ݗ�#S�X~���@��%6��q�hW7��<����5�ϩ�b�r�ș����SƲ`�>_@�ME�Ɂ�;s'���5�T<�� ǈ��^x.��6���u��"�*�+=W|����'�h�oܪ!�S�n��	a�D&�&BmJ�M�=�{�]w����]�������IY&͖��%�A����֡M5�.�S��'��C��ff�~Y�B@�4�7����%\ުs,]�YQ"ݛSϡ�ݚ���9�P;Z�q�������oStd�a����5L��yl���
z������,�w8ԋo;ݮ�->��/�S��eV>���Jr;"/vL�s�t�Y��Jm��N6�ކ��\[L�=�Ũ�fp���zn�þk.Ȕ��FLj���g�=(\�Ɨ�ؤ�ɵ� T�}k��"�ֻUÉ~"aŞ��ё��+_8�!7L�,�1�՟�oa��Q/j1�����Z��gތ���<i��L�B�a�㵸su�[�7�'v�@�/Wh0��빏�j�%u�-U�SI4��v��A�Ϯs�g|?��Y��^��٪"x?�	�/��_�2��\ޯq�T&�YZ��s����Gs��Ws�{
��r�Ub��	*'��C��/��G�D�����ޱR���(ֿ���܇�C�Y?B���β㌵wB`@�#+�V����܅?��U�)ˍ��t�k۶h�Yp� ����}[�(���%}�����{Ơ� ���,~[�����t�^x&ݱ_��������q����a�y6:`�x��q�SI��s@N��zB�����(�>��p�����c���n�F�ɘ
GBOX�ۆ��#Z��bz&��2���A����fXR�V�Sh�Q�m��(�����JX��V;67��z�M��n�H-��"��U��oikc��cjO�Ojzu�yw�/������|Xv������Gs��b0�l�z��`���O۝|�ۥ�coRu���r�*�N�T
أ��*��R�oM��JEy���7G�V��ě:7y5<$g�L���1-u��P�yE�G4��|�&!`�v�����^���ۙ��M��hni؛p�8�d�tp��*3����$����G7+Q��FQ]m�8k���hBd��4 ���+&��ft����r  �[V��xZ]��]8�쭍`��mn�z��8����O{/�i�f�<k3�d<x�/Fu���7�u�0�sW�E��6�Jݷv��-M��H.(��mr����x�����l��#z�S�^0@����c�:e���Siθ��������x<3�:�d'�֠�O
EG���;Q�[9�1k�y�\�C��)��3g��h�b~�Хc����fȭ�ul1���&}�v�kY2���d�w�%�Y��=����.����}!�1)֠��db��}ְ���_ZA�T�^�Tvf��{��u�"w1}_�����"� sM�2i�.��K*MLX8� �]tBV�Ax�&.:5��GlT8�wla�N�GP���B\�U�.� ���m�e�KZ��fPƼ�;N���%�̒�}?}����$XKaw烈ϼ����ʹK�E�s(��k[���КE�H�ʋ��y�=Z���Q�m�_����0�AN�z�u��ٴ�K��~+yx�C�Q^Ǥ�/)ƛ'��^m�����6����}�=Z�LS9z��kN���+ra0jffj 4�0��[> 9�ʸ�8�n���4+�e=�h�h7L��������
,��d&�2�x�*��LKywt������@.��!��&f�s �+%�k�w&:`p����gqNM�B6��5mv��Q�ۂ�Zյ;y��p>��)&AG��;[��&�Ԅ�����R�Q�Z4���Tb�x,��;�[}��u�-t��r]����c��}ȋ��18}�li)QT�+�C�Xw��&jx 䞢ޱ�������#z������pT��́fL�<�	��Z�J�E�)50�R"�
dd6��j�E-�pr���7���P3.;�	��K|a[DO�ZJi�*� �;ժ�z���1ػF��|�_1r���z�ױl6i�XTj x�X����vɶg=��HnpZ�����vr�8��1�L��+wd�۬=��_ʋ�[@v���%p��J�������ۮӏmoEM�D	��a+��cF��4]�@���:�W�z�A�qxf��ٕ�./]�v�cmfj7�����Sv!�L��-���]� ��� ��xJX@HI��xm�Ek�!��,��I۲���7�+�xEs-�=ˈT�1�ڤڛ�p`9�*�Ð�o��rv���E��C�:�
�7���R��m.2�ϝ�;*k�Ҽ��lrVk�������{������p�ЩH	�2@9�E6���G�aη�^�d�˴L�ν�ŀ%N�7��8�E]�f,��n�<A*�Z5�?u0�;����ö����I�:C��F�cN�ts1�	ʥvD+e����FE�]����Kp�2\A:�ʀ`ӡ̞wl��c����W-��#B��\n 2���c"����æ��;��P����dkH\��(�w����L�.��'V4�NZ�9��pk\}�k3��wu�T!�ܶ
���7��f�O!wP�c%=7�nA��r+���ZÁ�t%�Fj�S�w="��2�t��ۆ�v��`��@��!�����^��t(i;t�[�mWQ�n�c�J�BK�����V�u�k{aJG�U����9^m-�3���y���M�УAL�]��C�Lt5�圸���ċ������M�F��-1/*�]\'r-Q��;�5C�S\����D�Bp6x�ܵY� ��|�0�w��s���5;�q���r!�I�V��Ucs5�"��C^�a�����j�o;E�j�c�'O3���C�v:����VTYa���pK��	�H�N��(�A�.ZQ�����{���z�%�rnh:4]�{���a�P��p���2����;�!ő����W�9��ݹJ�N��1�(��[�� rmn�sgryB�gD;��~��
�,�`/BUp��>jvq�d�V�2	p�ڇ��gbt+�[���ob0K"eeh��>�4��ɧ�ң�%zPA��d�-�{��ɰ�����R$tC�3��0���
�q�Vi��
1Fg��qQ�鲿D�!"�L(K�
?����(S,�QB`Ӊǻb��"�&�&��Զ�R�[M�S�UJ7��IT�F�����PR[+�N �a�/��MWZ�ccW�:������������~3���|�;��%v�U$E�
)���E�L�I�MEQQP_������|~?��~>�GO�Pj�][��KM�F�%��X����h���:�[f�V�E��h�w��>?���������~3����{l_1�&��)�T}v�+Q`�$�f �����b�z�.��yb���[i(������f�
�����&�/��x�
�����I�jkaѨ�b*�"�N�BWTW�`�F)�l�@RPW�����4i���((��q��~�1�?�v��f �-Mv���jtm��b�;M}N/��*�+�}w�ݦ�m��u�RD5QSU�f�mR��VJ����"	;��j(��$6��F>���m�������Mh�g�(���֠��h���*&j�b���4j)��ձ�(������&���8���$����;q�Q+�M�	<�큯s+E�.�f�
��Z/L�����r9ʪ�1��yZ4 ��Oq����X_/�ԭK������$]%Q5
�0�!���h(`&0�lUBiݪ�����,�d"-�J�Z�
�M�]0�kER(5Ԉ=���>v#�����q�EZ�]���]~�������1?y,�˦���N��1������8<��x��7E���K}I�/�HP>���*ĩ�ܟz�Jv�'�v󭯴L�6�y�v4�ql�]�3M}��ߚ/����k�NX�m=�KK$�����B���,h^[��hlc�Fc\dK]Ӑ�>�7:���d�v����L2'�^F�.k݈͸
^��\[�^q�dކ�0�PU"n�V0��nf\�=�%��Neh����DV�a
��g�����%�(�)��#��5���d^��'�Ŕ7��t&lh�"e-C��#�+t�K����oN�����8LY�iVG��쎑Ρ6֭d3��h�x�ܔ���W�)b��vfP�3u����"Z�<6�����_�'���u�A�|s|�s����C��~� ������bVr�ؓ7�¥����Y2�%�2���zǙ}�
�!n��Rv^��G^�a�鸿�Z�G6׽XT@k@T=�׼!��P���%F��}ڦP����j�7�M�b�r��n�����ltA6zmvq�;�5Қ���k,]8T�f�Q+�3>����j5����U�K�+jd�:E�/FmGe�we�t�4�	
�}R��x��GM[*v%�n�نڎ]�W.�\��� �V�|����0�0�wv�0e��t�F�׽y��YR$v2�6��X	,�y��0MM>���.���?d�P����vWw��4f5fM���b�;�Y���7�}hЪ�r�.(Y�t�?G����ÜkZ�h�S�y�V��X�m�ͥ�G�V��H%|�(ߔC��?����*ƕ� �$���.��y>�4=?����A{Ԡ��]�+����B/���f��>�ք��1�����(��v/�ˎ�֤T��z�R$�vf�:6��v׏:i�C�q	�Vn/k�83�ݮF�����Ls c%�c?� �׈{�5��0o�����)�S+�#����-�y���STP������g��8SQ����x]� ���Z��қM@��)��O�ZS�3��&�؈�꒷���5 �.C�0*j,�_�����/5{�O��[�:h.ĿuY3!��F�ڡ��b���|��Z���|L#Ú�\[t�)�bZ	��!lQ�*��|�+����[f����ܶ��y߿7F�Xp�c��f_�w�?q?�>��|߮3{�j4������0D�,^��)J[{c)��D���E��u��((�;��#�l*�����}O�7���f��q������͸U^�CifT�X��`h�妴��S��#�/�_kکj��L�뫈��jܞ�������{�Yp{x5��-.�Ĳ�&�y��en��n_^ٙr&��9�*6Q�*�>c�]���&�od׵,U�L�w�k�1�-2�(q�)���`S����W�MH��h5�j�:�KY���$Z�N�: ^�.��?8%�3��E^7^t�ux���.&�M��w$���Z�ܿ)���a���Z�HyT�|�bK�1�Z��siQ�.>����{��|30��NGRa�
��?i�W�/��F�i���ߪ�>���޽FDh%W'^��j�l��K@LﳆI�z�Bm�{�G;n������,%q�G�?�ֹ�������2��Ł���.2��;z�	��6C�v[��Ԣ6�/Ѱ�ЛU���}�*z�l�����L'YOR8���w�#��`7�o�2���z;�U^����h�����s�nt:��2��P U/�b�����{�_Sh���iE�/@l�:ki�1�}^��N�j�x��b[1��Ϳ�#h��ܢ �l$�}ܝ[�ږ�]��x,l���]�2U�R�h���n��G�(�pr����	���V�IO���°#�J����h��Z�_�(X�p�9� �7���{y(����xŔ�ʴ�o���oK�W�^��>3Ӽͻa>���S��y)W��n]n]��	`�W�����]���v�n��vŞe�A�)��T�깿o�N�Qҧ1wv+v�ոIC\��{���l���2��d��Mqs���T�NL���R��x�x���O6�X5#���=���@;n�;0|MXd�z�W7���NEZ�i�&���o���SFVPF�(�kj#1Z��^1y�[�K�tt�E�ּ�I�a��A������v��ھ*��\�V�� �m.ޡy�6�c�p��>�8�W>r�+��Mߺ�wHn��Yi.ڳY�d�V�1���F��oOr���w;�u�I�b�8�^lu�����D�B˙�=�H��Õ�7G�#��(�Q#����2�-�Q��ޛ~a1���W��L:8xF�o�����H͹h��y�>Φm8ø�_�֢3�_�đ���j}���Fp{}b�;��]|���+�4�����t�����@���L�����Wu�8��`�ͽ�0���Ź*!�.Ĺj0���l��S�yr�̙��M�b�<yW�m奱9��Rv }���f��y�)���ک���$��g\�E4����F�~���'�}���Y�;ERv󋽓u��]W�����r�&<�������ܻ��+�	��c&���u�YӚyg{2���4��9&��5�Q��-�O3\4�Y^��z��Z9�5;r������J�byb���	�}\Y�A���Kl���7ܘF�����a��}B�f-�~9CNT�;NcT��꧵�����7�5�:ቅ�d�e���]H��vƎ���(�� ���[o�}��\�F"�P�m2��k.����"m����ZS\\��y����$���G���3�SBƩu#Sjg�f�bڇ}{���.�-�NE�uo��U��y�8�&$.C7�V.�h�㡬�
�D�1�7��+E3��ϱ��
 L�qV/NUwLiqW�j��e���Nݻ��X�]�mJ|���sEG�:��(����^F�����ޟ�=;)����Z{W⼥�?�׶�Y�^fN���\�����Q%�R;�λ�ݨf����;��~�B�n��v�']F�]ÁZ����#~��˫Y��D�[�\Ď�'vt`3��"��T�r*d�s$��x��b�`k��@q���幼n�wڸ~V�]�s��V	���̇W�C_\�Q�E]��wd����U>kgd���T�h`c&0u䞊3	��x9��2�l����5q�R�j�@�Keᵰӥq�*��4hU]t"��������wQ����廒��B<>�P�z�X�|�Z&~���w$��L%�C �j�����=��a"R��q^�/��,T��7V-7|�Dy���iܮ�OlzѯU{�Q��i�V�T)��nTh[��VkGS<��ɜ�%?�l_{������|��m��G}����h�<���T�<Yy�����=��ށ��x�����Ĥ}"�'�SN��)�ﭺ�g����Q�:��ǏHm�-�\k�5鍃8��Q�g�|���i���i�0&���z�������m�h�c!�n/тN�!�����ǧ�gτTU&$�ְ��F�~{��j�m?B�r"j~OUޚ[:�a����S'+�����+���eɑ���Z���7t�g],���hW]��ӼԼS/�8�&�+4�
��yC�)��H+�nZ�g �>�?��/݃��v���$E�t֠]��r�pcY��B�qI�˷�{m�����2ŜA�ؽ]���π@k-�/�<v07�\]7{���rCg��h�e�c!b4���ｂ��~�2�M�w�:��²�	��Q�b�����LWF�����|���s���mz%�z=w!�\�>MJ�Vq�hY� ��z���\ӝ;����r���9D��K2�S�z����'��ވ�RNw�w*̿c�F珺�[��J[`�o.��� 3��/�ɼe"ǣ.g��4��ni���m��y��+�;������g��N��Ȼ�ٚ^<���B_j���ԧPk�N�9:��C���N���V$��wDJ�U-];��5��cS���k�K�Hn�V���0ģ�B�ME���:N�����=�������?���?�,�n¼�l��v�n���οf�ܿx��e7�8�����f���՘���g�|�O�M�"�6|3��)k�LA�����y��������>G.�`�R�eAVkz���wM&b{y�K��m4���*-���55\{Eٍ�;Ĝ�����"����~Ϲ��M�Y�І�.��V㴩�MV�ܟ>�l�[�5�WGC��(y���g��c(�T;������Uw8��z���?���:�_��2�}ߵw�=N�A��w��5�dվ�/�� ���q[�FO����߁-w�ͭ�1��D��S���nҕ�ͤ�\��j-�uA����>'w��+�ɳ��E�Dl6d��d��t��~+F��q�o)��S�9o�fp�n��(��3����- H4��Cj���5���xB�гۘ���?:���dC��N9����pHW)[�)�B���`5eH�/��&ꛭi뛖#d�Um5j}�ޙs�@�#<��Ce(��u���KY��
��s|��S>Cda�f��z�"ʩ⦃U���wҳږB�vdͥ눞��-Ѽ�j�V8��ʑ׹�0��u�}���kz}ί}ܖǭJ�=8��e+��xοD�=���N�+y�e�I�"	�����5P\�TE�ƴN�5�j��T{:��D�o��W0�f0EwfڹңD�� 6���	Q��K7�]�N�G��"�|�)�Z�[>�Fq�q���P�wyPCjo3�fe'RF�ΦQ{	M �AL���H�3s.n��ƺ�w�	�|�p�f�l߃'�W!�h�
*��tgBY@��`��Wgr�0�O<v���q��	��۲Y�/�સ?��\�:I���t�$gh�g���]��S�u֦�WC]��� ��������i����u7<���:N��.!�rR9.ux>Ͽ?����\��,�RA���=u7���Z������ƪ�~��T�wW_��zЬ����ѽ�fܴ��ԭ��آz�!�DB&:��l.[��D�ˡ��n��7f�5�fP�Aľۗ��Vr�k�y�?�{��2�9 "��;u,'�R�r��Lԛ�ӂ���^p5|�����d3�L�=5�#8���A�n�;W�C�˦�܎����ә�l�Ǟf����<F_8J�B=HĬ�ar����qc:�Ι�W�Z�m����2�o�]u�`��:���S�tf#p�|<�`�2���Ɔ��{7B�hgS�J��ڗ��9�����ȏ�Kk���(���d��v������9ܓn�� ��c0�p�b�s�5�t���<�����i��7:e��nJ�ZG��dX��\n*-hOT|�7:���7��iw�O�Ӯ���x�'��,Na[ۖ��t?]�{̘�Wu�i�]#2��;Af;G*|ȕR�a�ob�rj�n����2��R���z�������'���r��=�f?	�Ih�(]���P��K���"���U>�(��B's��J���7�9��ټ�[Vڤ=�u\97!�ݑVv���+'6g53��x�f偽�%�f����G*���ږ��Y�K^a�����s+܆wE��gI)$ǿu|@�=����%|��l����ЃOs��s
�v��Yn�����g3p�5\�	V^�l�wQ�lf����'�{����B���~�ʍ-]W�TӸ,6|뷧!`�W�ۚ�ќԗr	�t�2-��xT��M�-9�޼g'�|��{��P�����F��~�}����7���oh��DA����{� 2˺�4U뻶�<�>n����jyW�n�P�(=�^��{w���]>5�<�C�rb�VB�ٙ��rݡ\DE�[��G	���J5x�뜎�p�#.+)�}�Z�3L\���u����X�.����sF�7�e���Nt�0��*�uz2���T�G�:�΢�+�Z��m�{�6t����z<ũ�te�"sJ%�A���en٭i��etO
�Lq��OT��(oZ��h*�N��i_eܘP��C�"rٵv�{J0����R�&��A��}�]J��:��Uνݔ��V�2��i�mF��lr].�;C�GK��@e�g<��Are�eU�(�l��}������H�J{�}z�.	.i���%,�)��y�\�a�:�uˋ��ݤݭ��^��wMn'*]u�;��ԣ�����3���@�	V�cT$������E�ز���*���=��R�����Jn�kk[H1cf����Ef0�Ω��	}2���w��FS7
=�٭X�F�Uԯ,�`�o;2��!>*ic�-����KfV�O��9IN�J��	���&�D�E�eQ�-�9[B�J�y��m�5q�$��iYGn�unu�$�����Z�յ�í��Pp:3NPD��Y�8�E�5��yh����y��9<ͺ��cР�gnV�[jRΧ��ޕ�y�"����K7xJ�Ĵ�i�wx��8w�k	 ��x-�	�r-TG�{���͆ɮ�V1�/���m����&���t��N�c|o2�DY���t\n%6��}�E��8�����TN����a$��}�������Bۊ]���)ܠ�� V�֓hV�]of��s��SڥZ������L;�62������n��+��?���[fev�b�os1�盱�|�_Np����t+���*�XLH���͝�{2���k�h	0�i[��T$5�Xɀ��ARw@N¤�w�3�c>�+�T�Ĺ.j�Cla;K'*��D��*.���l�,R`��Ǳ�p91*.��|������m����hw%�U�c�'%����͔9Z$�v��8j."��g��b�ӬL����sሮ�s��8��B����V�٪�źh
�oQ��q�I�^^�2�x�m����xJ�)a��-�1oT<<����B��:5��h��ɾv�5��:��B�˃�(���o'��Q����`3>���]Dv����-�z]��#���uvM�RJ8�- q+t��#s_�js���
��V�;��`�w�\	�뮔��(xqm�n�A��[XaA�n���'�N�I��������[uyu�H8m82��9��5�ak�$��S��W/�T�ȡ��
m��m�G[%C�:Ǧڼt*KxG<w�Kk&�M�5Ʊ�U��ʎ�N'�r$�09D&(���7�����প�q��!&��(P�$E�EE��v(������1��hր������Ei5�EU1PT}��?o��������������Ǒ-�PSTTU�3C婨�:$*��MS�b"���<�����������s���M=���?6j�&�����ATE���E�"h����1��?o������y��~9��wx���$OZ��Wl�m���c�QE}��o#T�k��������v�5cbhә���1��ڢMf
)5�����
�h;`��'�Z�7g�j�����i�c���ΚѨ����vKjf"�-��]y���nb.��ݴE:������S�i��4�����ѫ��Z�lj�����ٶ���(��:��Ӣ�&�*tj6Lv�4A[e킢}-�j���2X�(�U��Y.�	[m�F��:����=M1�ߝ�x��%Iʕ0�SIB��ťnv��sl�ǂ�q�͹�eB9<5J�nP8��p��çt�SE2E�*�9����SA�ﾟU
��z6����Hǰ��H͏>�o0Zg��PZ�K	�����vm�Զ���%jAȩޤ��������E����}|g�Lg�����u_�F)or㒒q�*B2���C�t�]p���R=��m,&rC�_f�nn���wf�F̆2�Y�.͓m�V��uKݞ��a�����{%�:��s�tq�EF�l�ܐϼ(Q���ZV=c�x�eL%�"l���]��1����V.�~{��;�gL��ᗲ�w.��k(;�7�[� �9x��2�%ߴ3͙ɱ�͊7xK��:���d�u��QF^�r�{����C����F7V�1��L���}9�.�(Y���Ws����l$ET����n3:��Ϳ}a�3�U4x���U�SБ�%+j����ISig�Ͽ?w��r��%�f[���O���?
8\�q!�<�vr�z���4�ěc/w��W�Dm�.� �g;2�R�#�C1��"S|	�bS�}�Gi�>�֊�k��آ,�.e3�c(',K�����n��u��ѵ�9N��w�oX/B����i�r�l�J�"�ײ����R��U�)^+[������g�co��Pk���+�Z��|�6��xϹ�Z�=���Jf�?o�� 2�5]�G�be���;��#��9�]�|��-�,���t��&tWu�in;��{����:����O��ޟ�ZlTP�m���0�`�6޹��.&h�N��E�y�≚���{�׻�����ď`ӗo�^��^7j��+�e�S+�����#y�ٹ�U��|sc�H��!�7�O�(o�Q��6�_�p�5L�{"�^��|�Q�y�o=�=N����1{�5P����c�+��>��$uf��dk���v'���dOL�͙F��c9י tPu>0֧�1۳� A����}�=U���N,�\�C�ʝ�ɁA�<�r�x��i������|�	3�+��� �5�?=SMj��6w�sS5����K8јc�����(��p�i���1`\L�g+����A�B����"���̳z^�x��9A�Ö}��84ӪEL�����3�ݝɯ���1�L��R������N��A��'���zN�WH�Bʁ���#����R��k���<4CE8�39��8��$��y㔖;/�-3ؓ=ȡ�qg���Aحw;hӪ@ul{�"���C	ȬM�G+�UE\��>9'h�FN}��6�[P,��R��m�Jo�U�R�d���r�[Y'w} H5��\.'�t��1_��|��}��J�Rޜ�YZ�Q�h��c�ںפX*��s����{�m⭎�CU\�M��*�$�������g�'f��[V$���on���K[����9�|/���5�]��zg&nw�����;��^V����P�����Kn�Gq�d�����4f`��h�gF��d���H����Ǜf����5ۮ o[�[��u�_��`GҜGY&����w��]�q�wO��-�l?(��Y;��J�|��1T'�}V�,�;Aj*@�O�)�z�1y��0���t��es=߻l�of�����N�ޥ9���wS���}�I����l� _n�כ���e�\9u�h��� ���w�:
��;4�`8�^u�x���i��@K�݊���sq'&�<�:�YBm>f�=�æ��߀`MoM�������`�!�"���.dn�t	՟��"���I����;�N"�[�x=�������ؠ
���hXYC���9�q�n�8�Ͻ��g��f���f��ń�@�a���T�\���h~����ƜEq�Z(��4g���U�ɺ�kO��\j�+op���YID��-�&��!�x�f�d�o
p������jgTo�wn틨���z$��k���i鉹�����F�.C'J���"
���'�;<6��j���L�Dg~p5�x�e�/j���v%�0��mfV���=q��}�Ý����7f�&���oE*�x�#�uL�}-��O�vf33�Wn�6�&WU��J�f���c�E��b���ŧ�6��B"n�zy����������u�jqy]܎Uw�x/����@/K{�eޢ��Y�4���[�f�v軷%O�B�{��m!��I��������ݺ��e��f�	@�!�Wb� ����C���ajUۢ��ה�SBK�kl�#���[���+3�2��o�6S��t�Z%�6ߧ1�]�Om������	���|����f����^�+v�[!Y�s5��M���}a���G����5_eC�l�ќ���G�����uj�_�w0m�[E�=qN|�u��ո��_��Ƒ6z	�Z�"Jc=���T<w]���1ۗ)a�$k�g�:����#�-��ce�%X:�|�-�g9��:�z�\o�zxxא��އ�w2fӏ��(����c�ۏFz�R�v�b��y}��Q�0�`������Ī��ړ���b�ג�ҡ��1ܣ��^��f<zCn?�4���w��ײ����b��԰Gy�*�Q{��������v��o�����*�Ө1��\e�m�]��5�fZ#�up�^+���d�d�`^c��7�.�TP鸨`�\�-B'q2��}�m�{�����qWe�U�}�F;�mJ���YK'Y��Ò~��7,�<#�^����Ȩ��Z.Wf�:�)�y�mK�o��U��b�6Q�_�~���p�
���I���t3x��+A$�RX�$���>ä�gP\v���P��� �5�jL5��H^��V�:���|,�a<y�^�s�b��y�>t̕�^U�ҹ�g�H-�����%\�����!L���v�}P+��/X���OV��D4I5�����z���l�TagX�\ڧuI�ESz��l�Sx.��^-h�W:�]��=�o���BY^d�JP���n�UqIH��+f^�a����zC0Κd��p��׮v[`J�T����#V��ǆ�cͶ0��UsX��i��@�k�I,X�����,�� _sj]�m;�ύ�Tde����:��m"V���x����k�<6�3�G���q'nA��xe]��7����{���n�>*����B��!oCm�,�.�l7r��#z2�:v�ē{�=h�=���׺F� u�՗Q��ql0��rl�iU鞊�5Z����OS�x�5{��d��d56����x�o��*>�HJQ���ER����@�;�� 'o�J�y�H�%÷F�.�ߌ6W�5
��m��=�bIb�*�j1��&"�m�Q������M��f�=ڐ�{!�T�=N��OMA��F��S����db��5���k��z�,��s��m⺧�T�~f�a�h2H0�>����?:�i���ݣ�u��H���T�n�f���\�{ֿn��=F���7���&���N������-۵H�&@����
��I�Nw���+�I���5xfJ�qB0ٗ��ͯV�:q�:܇~���vU����E��n�-��.����=�bp�Ro�e��6)���2�<_*������/^"N1��)�&f�O撼/x*(۴U��C��F�S�܆�v�kZ)��]3\��{zLr��d�
�	�B�mzy[�{���J��H�qZ���\�t��-���tr�ET��5�2����PK'#�rޯ��v7:��sݶ�=v�u6m5�s-hW%�>ޑή}ܖ׭Ioo>�Վ��2�7�;���wD�@���ȕ�v��z�:}��=>�32��
J�^���|��%[�γC�j��ث���1��j�ݭ�W2[����@!m�^�a�f��tN�֩)8�g���MF�[�gG@d�ڜu����u�\��Mm�*�+��wQ;\��k,h���
�^��e�R��:ܫ[�֫ǉ����;�vQY��5�>�������:�����X}M��9���A1#�f�\�E��m>CP�3�4f����Zf��'j�d����c�[!s��z�H:w{G���ؔ��
�ii�Q�+z��S���^�	k.�vm-��MQt�����M|���"ϧ�W�nwD��T��pD0G���|���t���;R-��w�V�}o��"
4'��g[��c���:�h��u�L�*������//�B�_/>�܍Gj5��R�`V�X���t�x1F��\��K�dA�a��{#̓K_�b`���$�T�{j�$�p����{����tQql=��b-�U{�c7�̂��{�q��<��=WSE�ihiYu�v�*ml]������� ��؃{�!�F)ص�/5(��,r�Ȋ�16���/V. ��'�$%a��_E�~�.���s*���>2|��`U=��]UYJ���LJ(d�&n�wn"	y�K.X{��u�?']��z�2ko�z�_t���Ob�ƫ.�C���!0�{�`�z�zz��@�w�^�g5ұ��?	�X�%
�֛H�ƖM���1p�YJU���D�\r΋ް��V�N�.�}���1_dF�l�ױ����
j����j��{r�]�Y^2U!�ԁ0��`��4��9Z&���l��0����{\�۫�M�0:_wp��>��~�;�����ʧ��~���Ň{ �i�BWuBͺoO�t�\m\�{����޿5���5�]���^�J���Z���ʞ歌�7�����=�c]��Dlk��Y��$�|.�����lrl;庖�[yPM��������������Z�CH�Wپ6�,�3��GZFK33G;�J���mҶ���d,#Dl�s����F�ǟgd3���ս�pT#��&8[�&�i��wN��k'v4��؝��T���=��ΰ�����P�߫�o�����t�5�]�1U=�Ȧ�'y���b�x�B�A����i�`�Ј�0���3*�g�m�� �9/l��Y�'�
��{#�ʠ�:��Rk�c�է��2��~�{��4�	׾W]��'�Vo�:� �^V,j�����+�7�Z�o��[�����ן"V78�M�Gy�:f��1jJ������z��������u����:�!F�2�9��6ν�]��Uf�� <g��c�w&� rSs~َ���g�q��y��P=!�t���[�W�ɾ�ZO��j���3 ڑbɜ�m��������l@gOj�xa�2k!E��xPa����;H��2��@8c�>��`λj�Ӵݥ�c(�o���U���ε�����>oLϥ�`���.��yF
���po8�e��&�GEf�U�z''����!pӴi�R6[�d2�G���6n!���&^��L��'�9�P+Ȭ��̋T��l=�G�~P|BHe��sy��� �x&��YB����E���-J���b�S��6�n)���ff��{_�z���3�:�&�a�k�wJ[�J�p8�,��h����߻%�f��+[�3f�K��8-��F����*�%K����76Vf���Rٷ�%������{�W,����@~��/��S��ﾗ�����H{Q{�^Okn`ה2PZknf,#n�>�>ޚ{�����4�NE���,9�Q亹ĺ��K������z�*t��Ѳ`�ji�*�,�˦�n�:O T��CLs6iT'4�剮����+$�yt�^Ğ��o�\���</�
�iLF%�_.��ұt�\c%�vep��&ÀQ����b�$��/�v&wym�ÛJ��<��X�2+�+���aA�q�K<�z�6l�H˓�$�$�GC�V�J��]_t���r�jܧ�W`B� !��4���e3Mi��~�	�+bBW��V�Ƅ:Q��ڪ�ۮ���#��2�<�qq�Ĥ�0���٣��SM�Sx�W�S�#��u�W��ܝ�%��[jPO+2��)�R���1�+
-B��_pmܲ&�������p�:�+#1�U��p@��Ϯ�,�Z��:����P=u�T.�<��n�e�Ky7�,��m�M#�wqzm=ډ�h��q��O`hA��t�X��w]ُ6��Էr���R��"�?����V�Rykx۱*�ᢶ�i@2�-}&c�R�Hud�����t�X��/8�LW���!u�i���&�Yk�bZ��Nڙ�u�%#N��"C�7w�x]�Jn��Mp����pn	[�/�夢����J"�v)D1�X����s&�5��w1�Bɸgf��H�\�Q�� ������8�ӌe^9w��Y�"�1���_m�ӡ���N�0�3I��J♊>�Ywk:�� ܇hD+�''x����wL��r�2�G�4޻��.��Q&VX#Wn�u,mMX��h���y�mN�I�b�et�)�зz�͍T�\����c�IdbP;E+Z�؀��ǵ�[��c�:� ���e�W��F�����.)f�һ��7����t�ٕ��=l�7�ռx�q�ِ���Pݵ�[m����N�@��wd]�-m���&�:�B(�#w�uj�U��n������E����څdB�N*J��, RT^���Pќތ�N�P0Ђ�SwyK�m��"⮛&Z�s���vWLzc�L��j-���n�Q�ź��A�(�/FqP�u�dd���:��ݭ��Im�չ�K�y���2C���p��(3���Z���vi�U�(���d��u��V�P>�|֌GH$@���D�Fݗ3,�t�mg1�%���[F���Oh�'_h+D����7��0�\wnp��ݣ�5+��@�f�m�We̕6,�N_=��]1�� V�k�	X�<�o?�[9o2��B�25f�c��V��#�Ct)��<��o@L9y��K�]���P��q"1k�V9�ЎYJ���+jg,�Zr��De�U
����P��&9�24P��TP�͗�#1��S&վ2cڸ���H! j IB�,���܁��1K��ȿ�Ԧ�`�ā�Ȉ�b�(��Q������w��yz1U�kZ���7�~��g����������y��~9��{¼�#��E�tQvvL�b:y���ѭ;��D�y&h�����mX����w��!c�f��v���y�|~?���������y���y��-	|��i�����6�[�������:��
nݵ���4�n��q��s����}~?�ǟ�������Eq��Ek�i��]/Th߽���]�����z�.�ݻT�g��E�]����h�j�t�U��us�cPn�6%�H�n�#Sh.�
h߻�k�X���1���y��WF��m�n��������:۸v�Z���4b"�k��q���f�F��;=���;��]��#�u����6�Tv4uӻv��Si��ݎ�nw]Tuێ�*;�]Q�[]t��o���P�7n�5�PRtoݼ�tW�u��n��57������٧F�j{������gu�w�Ӯ�"�hꈍ���lWAA�Ɉ*�x�;b�n���&�m�֮�u�n��qkk���#PG\I`�� �h7��CR8E2���#D�E{{�P��hR��6B��Eq���u#2�7|O9}��������>��mn,����!�NQ�UX�$�૵���� ���d�B����E<�ES��%���hrҵcR���drz-������P�g2=F�Fa����uJ/F=�"K���NG=Vm,�z������S:��k��J|&���W�[���,2!���M�铵�4��35	��zg�}�5�]ܬ���5���21��|37�jd5֟40������FuV�r:��ri��c�Kr��V_�Fi����+�'��G���2J|#�ȹPkj7�z�ێ���$��cφ��L��΀׾�X��#�P���a�Y_7���0��z㿳�����bl�}��U��T	ؽa.�\`M��ގE`�*��նH5��b��{�Ͱv�-b<�e����>x�k�Km��
�elf�m���z�3�4����ވ���4�ȣ�;�!d��ݣܩ����O��t)�y�TV�u����6�̛ŨFn�M�*�y9��������ki���ל
CN���(	����@�&Қ��/J���WJ���c.�|�CKXQ�ܨ�{��^�{]����T�9���5X������#Wj�\4�{��9@F�e�ʽ�������M禮�,t����-��|�6����n�¿W�]�B���:��ӆޖ�5s����)��@��$%rVLĵ5ٖ���5�0mt�A�e;��:�l�� c��,�Y���j�g����m��pzz;yN/^̻*qzhv�Ԏm3r!�<��{�|"���=Jr�����,��]�M��B�,�7om7���9IZ�8�^臉��ވ����s}��#^/~>�
Uꮼ��o�޴բ!'�۟5�8����L��dt__�ȳ��+M��R)�gy�8�Ğ	���Vn��w���p��<�;%bg�c�RS>�=�I%ܼ�^��ʻ�Ʀ�[گ)���OOn�J�'Ѣ�x������S5Y���RbO��ǃp�QgMwފ/W����x���9#��>�F���E�5�����E�d�2*p_L����7������l�n���1�m�&S�2�܉�Qֆ�r[k��ps��o�H��&�=����w�Gם�'��|/ϕs5{}��Vk7�蝱�^�&WEw�U�Ѯ}Bx-Vtǯ"�k\�؍�Ŋ���| YB��NB{!�|�.ڏ8�<�������ea咝������PI�$��埾�i=f�K��{I�8w�L���؉� ���ᅟ�YA�|�P�9T�0E��C#YR�8Ь�V7Nmc��d#5K������V��z�+��#6o���M}͒�T���>m���s�b�7�n�%B�Z�wv�^m�xbt�K��o�ԛ�C�ǚ�=� D�]���{g�@��\49Ή��f�hL5m��5�e����F݉��jY��!��{5":bg`$��2O�*Բ�����c�G'z���Vy[����W��1Y�B	��t�xgp�����O6���t��=Q�����J�fJWwv��O�3�|���`�8�ӤS��xܻ��^!z�:F���e��8Uo��;V�`޾��bb�t�u+b��N����!�+�@�ߨ>�*��+vä��k��YQM��y-���1�M�TSO{j]"���h�J}�G��X�\�J=��g.=�$��)C�=2�{A>wQ{��G�����X�K��f�Ex:̰���
��	�NC���X.ڗ��@�uВ���L����kz`�m��R� ���Vb]��;��r��0GPꆧT����G�{�_�����m�s�ov'�����m�u�u���Md*&����5��}�l��������q�K�+u���S����e���r�g���TH�jA<#K�k�A~��ڪ}����(��[�۫-#�l��l>�|�r�j�l*e�|�v��������I�A.{�m1��q��nz�w��<��OU��W�:�PtMve�k� @����7F\|�o8�W�o���Y}q@Mɻ��ww�O�ς��逬�?��<��׼������h��8g֮i"�����T�ρ��9�_`�Kݣ�鯪��ٿ/�/x���Q{�]ʹ��B=�֚���)���4U�b�~��|Vy�˯�L���=V ��UtL"ڕu!�F��:�:m}?t9�C���r�p���+]}Ef�])�m��{Sh+�%m�r�c��n�R�dw|��_���hD��o!�d��3~sFN0u�F\�[ �f`�FY�6c�!�*�p�ڒ�]�4���˽�tﮫ���DKe-�hjF�@ 0��Z�n����	��a��C�VwBb�5Ƭl�C]��7��(d��f��5�A0q��;�γ
Чm�Y|���!�DIM�	Q�?	�U�����q�m��Oi�W�����0������6��+f�Jޞ�}z+7{E���4�i���	?3���&)f��N�|�H�F�X��^���y3g~�'+��1�o�܉S���-d��z���]�˭u����v�JX��6z�f}��[;���[ٲM\���$����E�/��H�Q
�Ӎ���]����ۛ��']���լ�a�G�n����3˸_6e����n�V��_|J�{�pc�!.Π�ݟ2���mBF����=[�3ì�R^���Et6S�����P�ܱ>Rr56jz�y*�ͦ���xn|����v|��fv�dn�}��c��Ƙ��eB[]k3�E��׷���p����X�&�5	������������.H�������l��/��ݐɽ#��<��I����P7צ���E�~�qL���w.I3mb���f���Tv��uS�fv ����e\ŷ:�&!Q�B���1+L�S��������f L�n=��:���,�x��Ƿz:��2������R��������z���ّ�z��Y��ޠ;�JHm!���1�,5Tf׫�\��w4:�g|�fU���V�[O��62�6��oH�^�+�Xb�c��8��	R^l��xј馯���:Y�ma���4�Q���J.���-(���RT��l�������Ԉ�k�����P|�1�="�!�}s"��Aǻ���a{�Q��u�^~�	��������='��Q�$��a`+�F*RS7�@�xiZ�����f�2�h�j����r{j/�ɟ^ӼLzC/fHd�L����s��˻���X�9����h�I6Q�L�����f��m%�TU�
�Z}N��5r�4WW��oV���h���32���Vm7AYar^&���B�ݮ]�f�uK[I�@O����WBi"�y�
����y[��Uה#�D�vT���
���c��kx���kC��P(�W-�y�V��rF�������5֌��|�"�4��p��̓���{p*��{g��>���35S��ʼ��ң4��y�*��0��im��>'��ns���{׭��4' KKw��`�����]�/Q\l��LZ�Lh����:�^o1.��\�n�䳚]Js��*3To%_ﾟU�GeG~��fݺ56�ȇ�B�a�R�����I,���mb��ݵ]��
���E}$g�Cm����P�+��{�Z��<��SZm�7�WWo����+��2߱��mHo6��f#C%3s�={yE������ƭ�w{}�KȮ������	���a������ə���$M�a�	��zV �7d������K�����$^� ��P1A���A�g�`�Ql��:ۼ�J����^���9��~q��H�j8r�K���Zٗ=Kf1�Xz���/�=臵q7ʽ�=�*#����f�V����-��@
z�U=��)�+ԗ8�(��k�Q��w����1���30t�.nNp��{T�{N_�獿;_�n}(+���`I���N������ͭ�e]�y��5~;��b�~�ڗ���pP9Dĳf���R���6�v�ƞ����3�PdP�DO��Yk-��oMe�z��ɛ1!x,;);�"w���U%9��oR�u�-������B��5)K�)Αe'[pG�l��3|���W����������yz��C5�i1�\o��O��#1#����d����:��]!����3M���5O���νu��mH�ص�wa-��+�9��]U����0;����~��1� 1L��ÏO�ڞ��S������&��[����] ��׹6B���0k�yz�C\�%���D�d��D�./��c�0%��<�֋�5zx�&�AO�i���djޯdxE��O�6%�"Hy��>��)Y�J)A3��^/��D5g;f�w(��ʚ�zLѭ��N�@����2��vՄ�b����C�k�^1dm5�jM�GI��1f����V�E�w��S�Ց����|l4�����Js�hs�%z�y�ӎ��{]٭+�ϼ��u�D/1c#�B�ܠ�ߌ�(?UO��3C޺�d
̋5����yA����׹~�&v.�z�9=��Z)Η��(-���3��X�P����iyi�m)���Y0�]���JБٕ`]���Q(�����_q*-��f٬�y=:.�|Cq��U	N�E������(i���Xg9�D��Nc����VHh�(): ��~���<��[��K
)!6��b`��{=����jC�C"��YSb��?˝�j���i�SŰ���N�/�|٦t�	�k�����zo�BI4�N��r��F�!�uu��;�1e�c1�EEHl���i�L���=���C)�˨L�[����q��ur�U5)�VBrU�*�;OF]�)j9ks��`[�\�P�ӕe���[�f��W<���e;���FG��	^_�[��q/c�&�^;���yU�\��ܠ����k�	])E�f�O��z�&�yG����'�z�^v3]�:[�88�\���-rv����x���[�G�9*n��2N��<��S7��Gݟ};)w^ܜ�{6�ũ~�` �\K7̏��^�tVU�>�s�	�D��l ߡ��9&��i����}U��~���Eⲋ�s�U�q��w�[���3ZA�:^emRl����~c�^q�f.�*@��{��{�Moݺ�)ʗ��E��=y��,�/�9����-xJh�k���jK���j)b�
\����;T��j��o����t�,�m�ۏ�+O�۳zS��a}���gjN��7�=�uݓ�����gnM���:����?���S����.z+��M<��'������|����Ϧg��YIR�W2��i�=9x�:�{���m�l�-3��/�r�G�N���"�ۡUI���]���{��#(��e'�/��0��H��>��υ�X��xv��n���\�h�~W�nt��[i��w��r:꺡����ղ�&�͡�(�q�׃x��k�c,��<G�Ij�]O�~�-��ϏO�_��Z���:�q<VeZ1v���-!2w��	[�{�=yd:��;ӆk��۝�7b%���hU7��{��*�<���-���\/ &}>�7ݹGr��tЪ �q5\�������:��=�׭T�̽u]M{M�$�EZE�
��j�������QrټfCkX�k�M�C������N�Z��>�|#���HF~�V��ѥ�����'���;X���|Q%Y� �SJ��D'���3SM�q�,}+��fS��*q4kjԤ��yx��7ۭ�̛mVd�-��r�{�-�`�h��R����h\ƪP�͌S�D�|w��2�]���i¸:J.�q�g5w���f�̧MC�	W:����c�h�ms��b���H|��g�_03]�h �}��MrW�_ge������nkyB�؈��=�r��R�{��lV��,e��AC������R�9кF�n[JT-/�=7���wg���9���[cP��T�l���:����J�
�`K�����>��!�Dko����h�*��{��^�S�
���}�A�u
����j�ǏlS[�d��lHX����=��j�oL��y��p|w�7�3Ոmt\t��.�.��-�wCsH���kM��Fjw;���^7`��s��P�n�RĶ���f�Y���a�Vj�ዜ<�'�B���1!�����ܩ�t	�M b�sJ,n�bg6�w㫚(ɷ�A��_Pк}��	YS��wu8��yj��48����ʠ���hj�s�����vG"v�l��Y��n�b��h^
K�-�c�S��n�|��]����I�ԭ�h+z�u���������/��w2��:
��S�%|�����]��G/5��k�f�P��(r\z�>�`���`ٱz���Ȝ����g�I������e���e"�X�s�T��
dր7���%�o�ؚ�8��Ǖ��UU6�|Jv�d��D/V�Ŕ,9����-���(���6�&�yՄR�ɐ�Z��/O��h
�ŽYaoPoz�=fG�z�~���ZXo%<htƊ�P#,JX�	��vP��u@_(�}(�0�4e�ƗnvZ=O�R��_�n���қ��V���Z�n�����o$�no�Lʽ�&� ������]���頒6�HC]�Rh=ME9��
��X�
7�V��Ɖؓ�o$�f\:[�:׿�	#�n*wp�WT.E|m����"En"/�����Gkq�s~?0u��������4.�����*��`�9`���t,uqpУ(p�+���X���>��Q���2S�ԭ^��x.��&��>]Ұ�z��2�f.�7#-}��(��B���4����.l5��f`J�G28�i�`VD��2u��M����d,�e\KXXcqj+/7jV&���3+vV��g��T���ؽ$��E���Ǎ���F�鎷ytb=��Î�9�U�����e��QҒf�]q���k���s�l��Z��syAgPĺI�o�ܶV����X��0��"击
rJ�;1�Z��宯�[�e�FV��1: ^���q��2��W�4���ִ����v���5�1T�ݎ��w[����mmcb-�����u�cn֮*�Z���_~�_��������~<������u�n�jS�u����J4��un�lF4u�غ��l���v�w��_�����������������]��(�wrV��w5�]��q���=]��u����ӭU��lM���c|g�����>?���������q���ηX� �n�[\]���ֵ��8�ZMtnرZ���s;gv��<<�C����ѭ��wpF�un�:q��y�wK'n��`��݊5Zb�l���^`��k\�\DZ�۸֢�v��wm�pumłz6ɺ�[wj������ƵV����Ѫ>���̇Z5�m�[D�h;L{�A�Z(��wuVvZy�5�4wnۣ�h������n#�؞�v�G~��7v믉yw���xv��u�;���]����m�N�Z��j{���E�۞�z;j>��o6���&'f;�;��S�n��OFq���,n�����j�N��m��u֍qŜU��8������@���%eoj�?�t���{��п�ye�;J�G��g{��v�ږl��X��J��Px>��`�$ǐ�{�䋸�f���rGj����섬�}i�V~�H�V��1|s�a�̜L���Z'�!֣ۧ�7BYi.�3Xn���#���N�Q��ix�|�b��yG���q��-�ګ�	h[��uf�P���=�o�_z檷��vwӝ淌FD�)�1]�W����Y�$�7��+:����q�/��1���
�|���7�x����%A������&(�f&{�V�$53ӛ���zF���g
��l�}�7,+�yܥ���z�ް�ʉ}�M�����O����S���)�h��a��L��u��ɞ�ot�WWt�V�B��E���m{�Fn��ב`-����v�lx���]��h]W%Ɠ"�t�[��:}�h���}f���7O7�0�����׭��υ�aiޒ�	@�D��.��e��h@F����#���u����{����������]��Wv�+s�$6ELJ�e(����44|�Lt�k���p�
Ԓ� .p���L��n�I�����JR�jhjg�R���x*�&����J*�:Ww)���S�if�4u��e�Td���ށS{ѽ�4��������|�D����b���^�H\A�� �N'i7�|��V�
�̗��ڙ��k1粞+�����isF,K28���M�<�,�[�ܽԆ���]���U<k3�9UH}��2�a�vA�ܶls��T���5q	Ҭ�5=GqUY숐:Z�P�r{� �z�^�:�#������*�����D�9+j�d�wQfcз۶�Ӹ����]W��5Go�!��������5�dk�k�:�|1V����[��'�b)��޾%������l�r���"x���tm;�4r�h���xy���x�k�C��#[�����'�y��<�Y`G֬W�䧔��gcz|-:w �{���'hq����S���,0�pm�<fvb��9�Q}q-Se��c׵}p�oT�I�m�t������Z��9������2��������V�y���5?�m�y�s���n�z���̛;���9�%�n���|��`�G�$iX����G������Hb��YR������v6�y�f��7����\|�uŊi����׋@.�%j��Ժ�~k��#1��?�J����g�b�^�*�6A	3!�^���>�'�~�Ml�)+ue�GUdJ�������I�o���Y�?��%1
��t���)�|�	�����0S�q=4�tv�=̟0�O�Bh#�=��2�:�l�tqڐO\eC�6W�ᦨ#辝�����l �|��:��5��4$.��0�!�Ϸ���5�Hf#���SGV�j��^�Dt��fC�C""��b�N*n�.3�������tşn�i ��ƝH�m�3���$Em7��6g2��<j*(�u�T��LP:S�7���ke�L�ݖ�>xʨU��V�	�[D��/ՙ��m�M���HJ'Մ'���A+�����ݢ�uWH��A`���;��'�HRbO����z��R���b�G�,8a�e��\l�ʬfz�z��w��5Tڽ�uhr�k��K{�!Ou�nb���b5Jz[h�5W�mvI��]L[]�;�����bu+ �C'AFn�qy���yMj���@��,�ܼY�%�2��>\��v�[��{&��W��_^nv�t�&�3s��"+��ѽ��	��z��xa�X�J���N<Owȫ�ƕ��o��8?�j�}���Wnzk��o1����d�V?�;��
�F�~�:�g�� f,T��1T�q��=��z��/kZ]�
Y���[��ʽ�$K�y1S���rgLp0)�'�M��
�)��s�Vu̲.��ªj��M�A���>0�VL^�k��-鎴b}]��%ܲ�Q����<�s��V�^���v\���N����s�ߟ8?����Y�@yV���t����!��ė�~���_�~�av7�#y�̑�f�[��8\��!{6ʽV�y<qsy�&}�����[.�s�hX��=#�������4V��ޮ���bh �vϺ7Xk0I��3�!��6�foz3��ɯjt/� �t�dB����+���;j�U\���P�� o��C�~c�%w�>�b�d�C��r�F�����^��+��i%�E#�����$b��=ީ'fZ�8ɼ�_:x��6����Z�Ó��I]d���-�w�pӻ�K\��V���6���}�`ܴ���@,_ŋ��5�����(���X���]�}�-B��3��W�c�M�o&�P����۵ҖM�������4o3�*{��S3���2o&�(
mЩ�����v́�g[�'���uӺ�A��z�i�D�J�H��К�G3k�q}���3<%-�;\VV�,x�N�122����[5Viyj&�5(�͡����k�7��d�eV�w8V񗌢p�k�Ƈ�A�K�V�����LG5� +x7E���R&�U���r��̕x�_XZ��Gd�3�T�4�Z���=���ŕ��|<��,�K!WZ�Ѧ�DĦ�1Ouݸb�'+L!�̻��/�i�S��Z�۲����r�P�t"~2Wm��w��Z�W�����T��u�#<��G@�����=җ�'"/��'N�[��=��l�v�;XvW�>�{P������ScK۩P�K�ެ�"f�:e��=�]%C`�tࡕ�l��0���A��7�Rb[�]J�Y%��WVD�>�]�;|�uSםY%b}���y�#�no�J)��v4������j��e佮-��^�d3�O����X�̯�3��4�������������f�Ev�Rs{y�bɵC��{�ԥ�ݺVY<����>�� �c'�`8ǖlL)�[���r¼�T�ha�#��Z��WI-�[ s���ʃ�}���{�&O��e�S7��ý�6�[������^f1��k�Q�(#�ʯvӻ�(��.�6/������Õ>P0ڛk��<z�7��L�{��]�Sp�.n�cxm&wG`�m�7��MɟE�{I�j�`���t��y�Gtp3�]3�@�@I]n�9S��k2��}PXg��GR�u�Y�ܺ]���N�:Pp�b4���77GqUV�-�檙���
�m͸c�u� �����uYm�7�㒕Z��W�̬4�R{h����Nh��ν�}Mj<'��\yʴE�Xu�}`n�y.��i�9���K��/U}���2Y���JQM�G9�ю�;�s17L��y"gr�g�细�ںYxc�L>�s#�|�aX�����v&�!ʹ���@�M��Bu(��8c�V�hV<Sm�j�-7�U��vd��;���*�X[��fC���?��ӛ�#T�5��$�,2_��?$�0���V��na�u��$�`��L��L�g�߽]��eR���� 9[d_��@�tk��I���!�&�l]���3� ��M��r��Pj��W��d	������
, e�6u5A�r��4����t��ffj[�<�*�������4��٠��QM�R�d�{`N�@ޯ=�'T����]ӊ�xk�`��9�v�����U*h��rY���[d�"�i�Ӻ�ҟ�/N�v��B�q�1�]\��m���ZS@k옎�1����+��k6Ѫڏd���}.r����]���@�������WP6�}C)5&��G�׮W���K�^����_��ZYC�횝������0vT��"���E���/
�����M:z0?��v-��3�S^\��lI6d1���v�/������^�*���q۫���t8�[�irg��+=���B<�sH�@:��.��4;�^u�r�rȃ�` �N&wB���oe�-��n���:[�`�@�B]i 9g6��u�v��-B��n���	�l,[�, �������*�6D�.��̴V�̼#GFa8c�r�@�x�7W	�v�l�T�ic�/� ��2c���W��q��^�S}q�w�֪�>�uR���Š����|��F�a6��O��^�;j'�t1�.�I�u��ATrBw��	�x��U�P]�y�iC;��!�v�Wm�9��y����3�[5?{��m�<�W7�`�F\���v��ٰͮ�.��ͷx��U 7U�{����J�:� �l�1P����z��z���/z�!8^=e2�9�}�np��5[��`�
3�Ǉ~��c��K��(�:���Ɉ��-�kvyr�U�j��4�����u�G�i��^Y��4���;��T�b퀒��<����L�B�z�g�{�d��Q�G�~��:)�Jޛ�^|���9XO@i����%^��N	qЮ�=�d�6^L>�z�ߧoe.���� Q4����3��[Z�MVig��>�x�0ey�?��y�R��/Ъg[:7R>�i[�e��*%���\,�>�2 쎸6�[s8�[Yj�٣�q
��5�P �I?�:i��n�W��N]���_du��Xo��EEF����@А'�=[�����&��]t��u�V�^t���f�m��]��˸f��S�$�HaS9�כ�����B*��ʢ�t��5=~h�7�T��D5}>�f*pm~�U��v~(��6u%]��>#۞=Q�X� Gd{�Ct���Cp�܈�e=v�&c}����8К�������߲=�t3�6* ����u��^��z!��}u\�dh*���T����EvϢ�U�ͯ{�j�6�p:�Ť@*�2���tG\�Y�mF��v筭'��5����x�G׏�.��	�>��nE�X�*����������n^�3��)�"�MU;�6e�rYb��(���Z6���s�E�Qq0�nA��n|���@=�}Ma��&�	����;�-���[t���>��U�X�E�q޳N��:�21��fMH>�ΜY<�]վVW��i�zU��KNjY�B�Ǽe`�,�S��m<^���KҡcE�p&M�ywCt$lțɳR�������C�N�����:�e64�Μ�v��4�j��,��;
O���h��:�ǰ��p�*j����|*�6]�~��Z5�L޹O{��5�㇬T�]d����5�f�p��: �ǎ8����r!lv�y�+7,6� =�f�t��=gS�u�w�qU��VǛo��y[��L��(B2��5����%B����#Op��u���;�]����BL�)~�֦��)���{12��~[),l/�j�u|������S���[3��vv�ڧ���2w�����-
of߱�<�ۭ�(����|���Sкs��X��t���Vp��R�+N�8Ӓ;6�y�_�aG{���z�3x7vM��N0�^~Pv��ye\�>��L�H�a�����L�c/�hh�:0��a�N:�}I%@n�?�}�����-�/����&?Q��{̝�G('O�]�����@K��F�������|y��隮����3Ů[.���O���!��Yx�fDM��ػn��{�-;�q��:�ue�$���E�hF�7���՝dHg]���ϗ������f���D *��ʨ�����y� (��dQ���/��T��<�}p���IT��A��Hi�i�I	D�i���10����2,4ʳC
� 	B���@��}�����@T��@�C"�wp�  w}���T�!�\!*#�8B@�$B � DB @�%2!�@!	T�!A�@!�@!�@!	 B �$BT �!B �$PBA � B �	�@!	D�@!�@!	D�@!	T_J !* B(!*�B! ��(B	@$!(��@4�B�J�!*���B�+2�!(��(��*CL�H@��
CL�HJ�� �@���J2)!*��0)!�#!��0�*�#�?�����1���b��4�(L��$���h�;�7���/��O�ֿg��__��/�?��H�A��?�~��}�?��!DW�������Z
*����@b�������������?����@��`���?��������������D���?�?�?�b���@E�R%RaR%T�Q"%$�fE`�bE���I���`�f�F	F`X$F	Va%�bA��A�E��E�A���A��b�A�VeHFID�bA��a!`XE��eQ�!U��d$YdYIFQ���`ed	A���iRf�e HFIF!@I�P
D�JJ(��@Ui
AJJA"&Q)T�D�T��J&&)D�Q"Q&)�Q&iD��Ra�!����o��Q �B�E������������xx�|���nT@x?����<p'?A�AǠvB>?�
=�� *�އ������?%W��_�C����
����?�{�%W���S�<C�x/�?��w�#���|�<T@o��w��Q ���� 3�:���y�lp<���
���?���P_����Q U���~�� (��#{��@��a�OO������$���DW�>��?�L����?�������	����QT_��?���U_���������!����b��L����z	'M� � ���{ϻ ����D<>Nx|ٶ�ڰ��i��Z�6�ٔضjj���&֥��e�ֶ�hi��TճU���%IllŶ�6�ٖ��5^F�&MJj��2��-U6�j�%JkUm6ɭ��jԖ´�m#���j�Ze��m*�
kT�cr�6!�Vզ�6U-*-U����m�����5��f��JՖmU����iXh�mZͥ�o��z�i�  ���J��u����43un�ۭ(��p�V�d��uUFq��T*���jVvU���wh-�6V�(����^!%-lw9ږ%��� �(QE(�Ɗ������0��65]��i;:v݁;��[-c:(n�B����jڳ�ҭu�D�em&���w� �`���M��颹��tA�k���9�ͪ��t��r�Ү�]�u��v�m��V�RYb��� UOf���'m��t�6u�5���P�WN�s��ukffZ�N�gCK�6���K�&ƭiV�f�  {���z`4�[V�60��ӛ�5L5�eA�ӎ�����:�ٻgh��jȌv��4�*�X՗� ��]k����8�]u·]m:�@�v��.T����f:;��Z�����uR��[l��[f�f��V�x �=5�j���ݨ-�E�� ����ݷ t�n� ��� ��A��  �rSYfZ��l0Q[< ���@	�(�: �0 tgB���  뻮  C� ���h�` i]պ9-�Y�-U�  s�� o, �;�ۀ � ��t wn@ ���pѭ�  Y�P��ٱ�E�Y-j�lx  g�@�=�� 	�  �j4 kv �]�@�U�� ���( ; {�    S�)J�500 � �{�R�S��� �10L 	�S�bi)T�Q�b`L�b0�)�CIJ� �  4    � �4�=4F��mi����jm��J�b�@      ��v��&��ٚR���+|8�4,^�6��x��V1�M ��)8Rbkj;@TKNy��d��QED�~�2�UPE ;TJ)� QED��:|O��c�?ğ�C�#|C91��cc	!��� 6������I� �1��w�|굊���n��DTI�Õ	��:Cb`9xNw(�$N�g\5�-Y����:ւ�b�hd��>�-�F<���Y9���]�ǎ��C(�m�*V-;x�&�w��pf&I�d����i�i���ca묱u�l��_=N �&�v�LZ�7n�7P�QՅa���P��!n;Ov�6�'�j�c�H��5m�N��$�7�|1�T�00}j��qa,�:�u�L%ZX��@�"J�g"kp�1�ٷWY����N���t,��	��e^\CQ��7t�����ږR�ȧ�+o*�z�7��!���:�HȆ'��׶r�X����J�,^����ۑ�ԄG^]2(lu�!��m`#�P�5&��)�����m�n�J�yD����`�kī6h/]�y�^���De�)V��Y���`l]�B�$B9U	�8�"�{�L�
��v5�"eKe�8�555��b䕻�]b�^�Ss1��I��]ҁ1�^W�h��ǍU�b�R��s
��ȩz�Lf��.,Ǯ�a�ଌ���%K& ��̢�"j�ur�ֵ�vDcf��f�iz��������6M��Fi�z�'A��I�l1�<���X��a�۰6 T�md3❹xi8���6���F
�e��,�� �6��Q�u��H^YT�KT�BN@���wp`3K;�n�u4��˽a۷(��P,x�Aj�Qܠp�X�x���>��]*8�� �U�E�b�%ѼF�X�q�1�(���L�u��U�r,u�2= ZWv;Й�oZ	��5D`aH�k`R���p���'Zv�ñ�f���U�����Yo65[ec�Fj�ܘ�TUo~V�Y �In�:�Ǵ�Ww���l��[�4����Īٰ��V�mfQ5#��a����<���A�`쐀+�s]ғ�\�d[��dn�f��̈́tL-s74��V�StsPq�ML�Ve<WCZ�=��Z4]ӰSjT�ҳ�XVjSF���Ģw���@����v�X��*�P�41��l�m݄^��Шr���e�PRk�S2�Ʒ��X�\�.۩ 3	j+Yr�	�,,����nf�)�N��7�m�w�J^���Zn�0�B鰲ЙLX6t�z�F$�e�0�X�D�1`��y������Z,DZ�S��v�l�dVe���t�%�ސb��j���UD,�kh��e1������0j)�7& `4#��V%��[˧`Z:T���$kG6V�CQ�kX��Zue=��rl��J�[+�6��!L8�)�Iu{-���Z�`�\�X�n��x�Y�+keة�(fadn�T&�F0�@d'Ml��r�xvnд�B�
��j�z4����H2��-'cPb�ηOg#���6Ÿ�\�V���0Q�E,N<��'��w����FF�E���KշK�)  �[u�?�-���V�
��R�M7xs0�{xp��d�r�\���!�1��*_�>�%C��VJ�e��b�c��^?�. Dc�p^���.T�X�E!#5�#Xl͗��:���ݻL��V��`e�J��p=�IDa��Nb"�c �<�:�KX�5��a�M�ѹJ� ���Oʴ�t�����7 ��=@�]�"����y[3JĎ�-����\�)3��.X�ydQW��MeŁ�j��,��.�
W���w��ax&Lua�;)J���D�|�]7�HK4ʺ�[B���;�Ej�YZ ԭ:ۭ-,ǽ@�Z��NU�%G�K5x�A"�f%�n�����4�� k�v�S.eP��:ڂU�A'�O��@@�.� ����V�����<��1�Q�XGq�7�GL	�!x�ц��Œ��j����3D��i �`@<Q��47diCJf�P�e�E�x��1�)Za4�Up�P��Uv�6,
e6�2�w��Rwy��E��h���]D0�DXtE����ܣL�"�q���V��!����J�B݊2�217^|���B��T�4ilMڳiK�j��0k����x%Y@�F����]\cr<Oom�Z�I��ݤΘ�y�N������Dl�e<�i�9A"]ɨ2eD�P�������f�%�Z�P�y���ȯdE&+؎���N��2��&�2 ��t���G���b���eZɷj�Xh�b�� ֍�Yx!����s�S��O ��c4o��0l¬	!Sl�N���z�H�9�X�$��c+;LM1�sm�i]��@/�Ve�:�Lǆ3i;XH-	e�nb m,Е���	R6k%��2򃶈C�U���Э��n��xۘ�Q:+�i�[H�)�06��fDْ�im�S[�`���ȅ&S���WV�.�;�h����,�L�������{�aʹ ��Rb�4e9�P���꣪I�2j�`,�Z$�NXdЦٵMI{WYx��8��.Ñ]�ǒG$�T���0E�7z�N� Й3VU�ى9�-7��o�2��"�pL&��f�G�7�	�C**����]�-�LctÖ���)
1�u�Qإ�:A3E*�s/U6�{6U�[����a88/0�_X�`�XoM�nô�vm��3;o��!N�&�i֧��r��f��f�R���[I���õb�*�� �G,8�*�T�&Ic���mj�-��Z����ՙ�ҙ��h�+1n���!��6�@��*������3YT�x��x!��"��{Xc%����Ө�Ѡ�Ȩ�t7\�u�U�����Y�]��9���R��n�Ʋ�ҶL�XʹjXi��"���\;sIuw��ݸrV�U��@�R����:r:⾑V��{طJŶ-7z��K�~���!9�VZ�5�W+&I�B
$ 1�&ilc-�-�q�iۉ��Y���}(e�=A`�29:;)��p���w5�2��2!L+8bd�X��7hj�
��j�&�5�nلt;8�W�iTq�mnV��ǁm�^�2�R�(��Wu&�m��J�įCa`�sr�{4! ,��L����'�:���rR�ډ���m��K��E����Z���~yC5�2mJcGc)���,a{Nn'��ui�շ(MՀ���&h�Ŵ(���Ӌc52�7��%|Eb�� Vbb�L���V,=݇^����wm�0hS�����ypN��K>�J���:*��Y�r�k��hn�Z��J�Ǘ3v^��U���1(!������*��Y�^� ����sh(̳R���7l�B�ۼ{yVmcֹn�p��h��Fo͊���3E1�l�
І���ٕГ:2�(�o"Ɗm*��f�p��{w���B�X�`�pGi���2�9����l�d�l�N2��T:e��`2
�*�uGr� �O.�ybF�kx4Rh��Ӧ�s&Qj"�jf�1��.�۽X�ـ̷.F,n�q]'��L�Y�Z��̱�uk�!`�0,�9�oBДД3N�.�,)�����cMb�z~�r��cX��g6��r�͢kZ��L�m;�2�P[����V��&�)Q��*_��6i:�����6zզ),h'�j�,> �2b��y0lgJ(�Y�c7*Q(૕��Sg�d��^�<`썼�3昭�5�$�TnƬ�YV1f�T���w7))�jڽ��(��,�J��q�"�]f,�[�n�J�\�m<-�n��- t�i�:�fP��H��-��e��H�u0�ʹn��L��+n��]����B[�cŘ�X�r��2LL���i:6]��v�z�N�,v7Z���[L�r��ڵwHkP'O9YW�hP���C]U�ѵ�v"[�6՛����E����]6�$��UȪ�V��������2�ЙUj�(�%ಁ�\?mŷ�v1кҮ^�4�d ;ܲ~����o2����zL���;D��I(�v�"f���X��,�.f�I����[F����E`�t��[OI�h��]��4�`��!eH�:ۻj�oCHeڬ�Z�h���E:�OM��'� zC�IL���{YCY&�A�r�ћ��֢ѷ6�S����,@.-9-Ȅb�jYL$a�����G�G8��j$kXF�wta�Sov��wy���ȩ�4�ƙ�0l�%̃�4^[CU��1�X�l�1z�F:��i�sU���h��,��aV��c]C/f���m�Ύ��[*� ��oB�[h[gU�uyj-05�LV<.St��teFMmj٠�t�V�ڵ���䰄&��BeYW���wkNS�
-���v��Z�AL��+ �jm1�<��Uۧ�h��N��`��:^GF�4+�lI�4�AN�R�2���5���E���4�9Z�-�����J
����м��=M9�)ҭ�5�n�ۥ.��G,Y8YTQ�07�l����XN��0�1|�τ���t�1Q�t��4�چ��ؔ��+A"�����a"�]���un�v4�{�-ʎ]Jk+!4k0�����u�4�Di�R�,�´v�n	osYoQ�eܴ�dL�pX�Ĭm�Rwz���J�a\��	��;l[�R�fR�%��Yy���LP������^��
�@搁�܌A��fTV�jnQ��Q�=�W ��"�Km����m"Q�zN�T7*��`U���T&fH��趉�B!��
Sm8ɫ%�F�'>Fm�Z%����ˊ# �#��x��
��+����_X���3H鲰j�j!��F3��[�bM���St�~�N;a��;�����L+J%˘��%;s%�!»כ��0Fbl�������h��7T�A�K$u|%X�G"�m�6KA��#1ᕁ��"j���0�&¦Y�Ct[�c���xs<�[#��0\��Mqa�6�(X�Z�Uy�������2)�IHuv!{f��zT�%*����Q�2���*b����ܻO&�+N�ڄ����6V�to����i,�R��w�*r�cr.j*�q�&�fE=�^X�F�NkݺzC8�8�[Ŋ�Gl���u��r���rÖH���vDB��\�4��U�#Od�5X}E�V��j��R���f���GEݭ�ծG��J|��t�wB�b� �`�1�� ���o,͈/��r�Js�5%�lR�Σ.n�}�[U��uAJ��\	��*
��h*].s�1���`���՝�W-�E��<k��V.VVU����;����Cm��K\�:�u�Nk�}5̂V��{��n��	�٫Y��( ���B��g<�o�X�x6�"��]wa=շ��c��cjRvu;\n)znQ�sl`ZH�\}��z��;���wh�y�ZK���Tz9����'�{����O|�n�Z�GC1]\#
�f�=y���Ղ��v+ʷ�+�tI ���u��PD�$�y�e_o�^���앵�[��ʮfӤ�7Aҭ�˒d���fҼ����
}�L�i�v��J�
]c����a��H�|	j�'V��ڹ��f����&VM��gf�W�ܣf�'�[����'coMZ�4�'4�Z۷W�����k{X�9qv�E4z����>HJ'9����;-�z{�oq�x2܊�๦Ut8v��,gu����f*+���Z��+��-����qVѻ$]�gFu&� �3a����d��%t�Kl+�q��N]c�:2	:��Zԫt0�l�F`jګ㴗kd�wh�m��u`ة9.�٦C�{����j� �j��u���[�Fk�I(�8�N�v�=n�����Y0Y�ӱ����mf���o��\�o����r�f)��]���K����j�gn8N+�E�v�\�e��R��Kz�YR���
���Ve�/$���un�t�lV���a�]�&+-a���w���뀼t1�����9N�����c����G�z�NX}Y�+L��V{�_"E!�SU����k�8�����]�\T��2۫��tT�W�pM�ifm^IB�5���2�.,�+�w�i�2on��9Q��۴4eݳϮ�(�1v�D��>���+�s.t�U΅ܴVE-U�q��T�?h2��QʶTO8�4���[�^>�i�d��s��U��@��{�}�3���[,xZ����7+ I=	��e�P��c`�f����0���J�x-Q�}�t��iӠ05Y)���I��t��w7��4���Cc�הb�v�A�4������i��_��*2�x�)��KUvg\�v԰2��n��[��ͩ`��x�19�����Xe����Gv�t/q���x�*�_W7���.����X�������Gi]5�d̵Y]D��V�WյsK�μ(�u���PN�!{tb�;0Wk.�|LW�Է��Π�S�p'+������]�p�K��O*=��@{/h����n4�Dx�:Tw����B���p4��m*�YC��vk����e��vlP��x�V)6��tWS�����v?��O]��՜^��	��(��M�nX$���a��鑜���j�:��>�^Q��i�vf�'�u)"ۮ����� ]qV+(nx��^�P�k�K!C7 X�t�j�;�iZ�[y�n��SK�o��3���hv�켘>I���:фs�o3W;��.��2�p`�w����o͈'��`��G�-�hX[)�7K1�C�`R	]fhw��VW���0�Ċ��.�$�]�s����e�I���;ORL��ޚ���Wls6���%@�<�wr�H{��@�j�⡛-�9�����.��{���v`�w��2<��-a֓z"ֶ2�6�Q���0�D���s��3)�Yj�H��o5�\x��z�fU��CH[�`;�km#�]�!�� 
L^�՗79�6��a6���=�dcvR���gZ'H�zgN(��=�{�¦A�����'o#��z���4ԣB�k_fW
P����ķ��B��0���g,��g$�7�Cjm;��$lQ��<�[P�#2w`3��*a���Z\]�m./��(.UQ��N;�N)��\�a.Z̼.��*��ØC��읧���5�r��[�|#���*�e�Vq/E�m��m^Pʉ�J�m>���j!LP�9��/H�Ԝ�����zjm�ujn�C��1�Ӝ�=�.�#���}B���i�Fj��f�t$�;#' �mөn�5����F�B���-7�b�9hV�L�\�KHO�޾�Ю�c�h@r�puһ�ŀRK�r��"���)���)�X�՜��*eY�lN�Vڍ��%�\�k黯;*@7����5 )�ثF�݇c�V3N�</0G��GF��-U��g��ͥ��I��.��\3�w}@�q�9*�mVJ�@<I<���Q�N�*B��� 
s�C*��3�a`㸫6�{V*U�_�����+cO�P�*�%uw}��\&���"T�/j�т<�����G״De��齊��^|��~yvڹ�����xv���Ҧ�Z�"��.�MEÄ:�i�-���gR�᧶�n;�X�T]�]aꝥ��wG����͵g�t������|T92�25�� ��\M.�\7��:@V��K���<���79�fk�:X<g��1T�ɡ��s�` �n��ǖow/�r���:�u��]G�!�;�mp���fu>���t�n��&%�wZ�u�%wl��u�YaZ��a���g�n�1��ՑI����'=���yR-�_:m�iNo�o_\�2�7`�o���
Qw]�/�p嬬x��|��v�Tn�Y"�����bk>�����<�6�(�����C��gW�K�U�v�O`��M�3�f��5҄�j�X��W\��"gb�� �|A]BKa���*1���_o}��Y7_^���>ډn�w)v�'�^�0�+u�p�VRZUbTnN�v+8T{zö����[��]�0>�}h�n���/��:�n�;��B�'��U�:��9�����ge$r5�b�Ø*޽��=�'/����Z{(��%�;��Ӯ��U������7.����PX�A
�#7��6�@����WB���+]_VJ�z��X��8�r��UT9>�⻌&��*��]��@[�L�ѐ�a�{3�#���u�����[�L�H;2^�kwiR㡮�Hh�+���ǐl��x��!q��Z�T0k�p �������O��Ǜ�C��*�9j�Y��hD��1V���.�S����u�G����C���pwopu�2�
qܨ �oec|5����w��>�F�*?�vBSāX���l1�b�ŊbyM�,�l3n��t�R��:�k!���Wۡ���Y=�m�t�3(�JczU"����IY5��\Zf>�����Q��})-��ԢI� �f�y{Q��%����Z7���fΪ)+�v�L�ZluV1Ab�����ne��7q�a��H&�z��Khl�v�ݶ����)�TF6'Q�e�������*Bg3�\lVm����Cw�Y��|�����a�6���413��wzF61�o���nؕϟ'x4
� l&�^)��c3��h@ƺ�3�Ы��W]�EѺ����9�*��E`T��a�B���i�j�
�������@p��2y��O���d����[Jk&���1]EY���r�3F;��<vdRb��&0gV��	�n�Cĺ�ygcJ�-	(�5��mg��ff�A{-��:s��]�"$L���*�s;�ǳ,䮬��N��C��=�cF@�<�+�ݝ��:�� .9�i=�Y�s�V�R����@��S��WB�2N�Ք�a}�l��O���L�R�{&������K�����oQaJ�_hG*"5�-p�-�o0�=���e��y���HwYfVU��/r�
p�Vm0�s�.��Wc�ac���к����
5�P�Z;��ҧZ�!�g��O>�k��;HF��J�Р�ͩN����-��j�t�x���u�qF\�5��?<�����r%��$ZI�8���ͼ��t&����a����׵
�wyA���ґ�n��E4�O0�WȺ�H�8��]������Ղ�{A���.ݡ�-̢�#��:����;][7j.p+搛Wݜ�\�Zn@6&�u%�-������%�V�5f33oe�8�D�s];���N`r�b���:*o�J�3�d�+FT-���<v���غ�r3Xwp��;y��_\E�v\�(��9>��h����������寥�� ��k���A���:����<Vk��ݼ{{���%c���:�.���5��f�'�oz�9]#|��Աݮ��x�5ܪ}+�U�Of���u���G2���ξ�:������<_n�B�i-��7i>e�l�)��s�&�q�b�K��˛�1���a�R��tm��f��TAw=� �T �6m��E"Vh�/xբ�>���V���a�cp�"�Wl\�k��#�nt��;k���r%���ũ���s��V�˷�j��0M]����+��\��i��nN�@�Z��2���z��fb�3��WX.��S������Q.=x_L���r����;��.���k8mm��y��.�gWtԏQ����<��G-�&�v�����Z�7��"֩Cλ�?7Z��P'B�����D�ɮڛ[{Ą�ʔ�zn����45��^N�r˶��ԕ���R,G.�hU�j>�N�s��<%t���f����(4�*�oi�ໍ�g+g�e�I�߶��m�նq�*+��*vdYʟ�����:,V��6l��㏇�{g6jNor�ӄdeH���7���o�1lr�kL�����~�����F9�M$��(��� �i�
k��@�LN�(����͑vR�V�*�x��;��n	aΎ��h�s/C��z[�Y�S��s^WT�N�'kr�MY��G�қ�M�,S��k���Cg����{��&�өt�u:��xMe�譋ҷ����M.�[�t�Վ?eN�id���ތ�][j��~����S�娇,<�ܙϷ:�
Ngoj/�`-n��n�>��TХwn�Ѭ<��db(���(E������ڳv�B�3ƻ����)�Vq��\/�a�[Mu�ѝ�ٷ�����< v�]~�2"�Y�G�U��WOt�Q���r�J̺�����^���̫ӭ���!�\��rp�B 38���J��UZw�����o�6���# iN�uǍj���ˢ��yv�y�u�^D�Í�B/kI�f���{������a"�A����X:��o�k���h����V,BR�:7�d*�%a�J�ޝ�
&fe,�>Ĵ�὘a^5+`{NwW/��\.��A���&����A$r_fȋ͙}՝&ޱg8`��g�v�;� ��XJ깼��$���*����#	<����O���A�>�ʍ�=lU,2�U�y���Y�[3	 G��u��Ӕm�7v�{Q��A��J�Xkn`��aŊF���ƀr���֯�顱���kx��l��.�i�ʳ{��^b���6�;קk$]\1	��|�t	x��[��6jgv�YW��;'��AW�0��m�s
Pqi7w��dE�W�R-*�9]�
$N��f30+�a(�;r�Z�e�	��ם��ջh�G�)�f6"z��}yKl�T\�ȓ�5wAkOF�a!�JWY��]�����V=��sQ�Z�����cZjc:��j�,U��֣��ʇ�ظ�ͧӆ��0�l�m<��k�:�ήTš|�G9I;�α
��yQv�6��ҜeXx��C�)�3{�s9�>��9Qƻ1.�����{�`�*2��؞I٪h���FTc66ݮڔ�2$�A�����K���6�����)Mh��玴�>�eD�
e��7 [ԕ��;v4u���ੴTX����R6���4���/I��� ���Qv�*�_���WMwp����#�*��cN#�b��+�\���W����4.;5���mF�`4P�+�chܪ7��5[mQ���g~�$��M�r,�+8�4���n��e��et=r5O6>y\�^��|��g�c�]f	��os�a�R|�\��	 �O�Q���9���S��me� ��k������Nq[{-mۤ-nY��"���3#渒�3�ԍl��;z>�=�nglͻ��p�B�m܌꽚���K�2��g,`&G\��IC:�Ž���Gs%@��E�Q��zM�Nu}ao*��)��$�I1soMv �(3盦 8�h��%��W��N����5���]�B��'.����⯠�,��R	[x���((
l�ky�Z�0)��U� *�pьN��AV���,��
�uo*��T��bJ��_R������t�(,������| �J�H/��%���#nvw0m�i�Ȅ��)ؼI���}��j����ʆ'�ǷT��[���E�������R}ʂ�ʝ*@�*�r�Y��g���Ֆ��Pʨ�{�V߂�v�-�6,I�TU�r ���3�����sr9�_G ᝼f��!���5�~��3M�W��ţv�.PygNv#���V�����s�dbԃ�L�7a���j��趢I	�]�f�}�X�s������ �&ѾOH�Ӷ������������r��l�֯��[�e�օ3hI�M�qt�n�o���Z�5�`۫�[�*m�v�[SD�n�;|�<*��҂��T˝�������I<+>�E���I��E�@',�a-62�D1�FS�;Ë����ę���w�>-Ӿ7MQ�9u<f]w�ձ�p;v�X�>Th�E<�������N۸t�����hU�[�]���ͩ+�L�Q�40[vo��Cjn�Iݔ���r�;��S)m���]hk�+��>��P[ V>Z��:��Ю�IW]�ҷ��͡�oS�>eJ���j�9�WVc�O�sW`W�b��x�d�ܶ�-�_P�,kL�u>C�.��� {�����x�X�ƹc���h=`�5b���q�vН���@���Q�*L���p�b��9��Y��N*uL��z�-�-��&�a�݌��d�����e��t��k�XҒ�,�W��#�ҫ����A��� 1���F�juR,t������Щ��he���p5c�v^/�l�(��&�	Һ�g��΋.�7G�}�:v������Pљ�RT����"��ޭɖ�s܊��xبM&\���hv���Z�P��Ѯʼ���XU��f��[���pU�u�	�5 �]���#��}5�n��2����.r�1�t��a��Ej�U����&���}��Uj�
fP������Ήc��p#�jv��wA\Y#�̆�
��m+�j]]i�i�bl',I
j it7w��&k�'�b�}[c{M��qm���.�낣\����@�Nq�{����;HB���]�,��U������k��x ��̤�^�m��@6���Q7�k/]�kqɾ!:�m�xfX�WĔ;ǎ�Ձg��&ڼ�k^Y2�&)lP�;RӼ��pڀ���K)�Ƌxʑo`��Ya��5s�� ܦI�@�wy�6�,L��o�7ZΊ"p�m��QRSWwDˬ���F�iK
,;����k]�y�&�:P�Z��`�G���۫�͸�w_em�ם��[ ���5�Z�y�,-�9��ńWq���hV��G:v�W��+�x:��r�W���� b�[��GE�|z^ �fC�u��햖#h�`Ln�Y�{|� ����2�b��k��ڵ{��-��U%���_)�����t	LH>�eյZ^`[+�*UY�H�#��#i-���+�]��G�|�b�=t)�\�{��K��Bmnk���1��݃nQ��<R�N�mۇ�⭭$�Z�T,�%�>Xwrs7SPV�9�-7%-�M�*d5j���x�i� \�+QD�%Y�cYYθ������'v��t���eH,W
Ǻ���pg��	�N�������g�S��K�Y����8�֓͵�a��U-��U��a]��a<{���)Eۧb�֊I�8�0M,_!�r���V�"Q��64waާ�YY��b��I�ѷ�W�,����Z*Pz�6U��u�q���c�\n��]�Y��z�8�9�n���n��7�z�u�5�L]͡Du�O���Ջ*;�Xl�N��ݎY*=I�]�V�i�}eC��O�fKa��]����i���+D�[[|(V�Tt��s"�Nڧ�3;�|!�Ws5|�-�x9����ƣ<BX{���&-���w-΁�3��v�H"��B�:a9�H6s�������Si�F��h�*�4�厶�v�wQzI��zf�n�>��%u������'mn[�J
�2{�kb�Q�Whs���d��}������3���t� ��6r��5��v�2\��<�]��E�Ҽ�z2�y+c�*s_tR��AwS-P�nM�$��EY��m�/�u�Q��h�q��Σj�'&��MZC&Y %��*�W��nA٩!5{���G�Z�-���d%/�e
�2L]D/��Yt�����m�)��o^�_�B��K�H�;��Ы�\��2�YhVZ���6��e���yҲ��O8���ڱ��,�V�ta������h�	�:�)G�Q{���IP��u����h��<�o��ٌ4&��5�z�X�Hg�8M]FS츖��ʊ���a��[�?�[������]��(cbP �����&����R]NőD�:X�K��u�tMmb�0��1gS{�0+�A��s{�1kNNO �*�j��[,�t�K����,�;���ˮB��9&�ר�[���P1Vnu:�;�f����B��"�Ż����@�&g:hЕy��7N��3[�j�3p���y��(��e�{�Ӥ�9#�6��Wu�׈��Kn�;�v��0�3�VZ`�]�Y��֪�X}JΧ��ҡ�������k��PkZ����@��ܮO���X���.!]���'w��Wo]V'ʉ���@=YE�����O�腢@�����s�`+rR=�b�lQ7����o����z��V��� �L���6�ԩm4��35<Ň�#)$�,̲{n�&�ى[�I�a�Y�C:6����	���rW�w�F'P/���b9��3һ�8WCs��������p�]�91e�h+�� �5����7W�"h,�Y���sw����
�.6sr�����(�B�9Z9fO���*�ؘ�14V��G�O��M�cw��^Q2�/�C��Ե�2s�ķ1��vƭR��!��Sq�*Jt2�V�i\^h�O4
"�\H��*���!x��crs����[p��ڝ�Z�{�z=v��
�7�PVo.�)�:����˞h"�Ξ_�@��E�٥N��vWS�F�+.��*����3.��{o7.ƈ1��|�#�>,�!�}ǫ-T+��Z��9�I|,Y
�;n��^�h��38/���u��N��8� �ts�\K�+n;�.6J��d|!�Vus����H�nü;��)���v����8iʒ��"��6ʕ���6���_�9ӫ���R�s,������.�n�34V蠠HdY���v�Z��3��ȃ�kݡ��Z�x&@m|~L
����4�0@o�Sl��t��� |,�����箋R枝��p����Fb-���.����5K�=b�x1;O�o�cc"�_�������_Ώ�H��A�����@ԝ H��?5v&��Ǡ��S��V�h���mÏol���v'�_.<]�8���J`�/���7AO��� G�\_ ��ʹ�p|��X�WJ�h�;�w*/��D^���ч�R�\��ʗZ�a�-�Ҹ�~�����G�E�����q��u#AԮ���:m�;��mʘ�U%słvx @8�Y=W�Q�8�F�
z��V��W��wG���q�e��=-��r_k����:�͞ ���{�����m/mf�\Ņ+^�c��p�{����>�ܥ:03�8Tެ��n��sg>$m%�z����,�7�ww`����D�{|*�T~b�2�������X�@WlƭM%��5�*�_���MY���i�d�o�Z���>���s0�r�!�-���1��g���I��ׅ��B�32�%ͫWEUՑ��f�E��,����Y���	K���]�B� �
�먋��=�9��Q:9���G��WV�ja�t��d����6�Na������9:�Lq�XP��!4,�H�e븲�竩�w��:��f8]Þ��(U�%7u9{��ȣ��N][��DSQ���;��.I�7'������sF�-'*w1f�'�R^X�N�%��,�C�nn�zzH�뎓����{����\�EнY8�1����;��	:U���q�t(�/V^EM�ʦ�2��)�GP�L�̮RT�bt������9r�F\I0�Q��d�HNP\2�I��5"�V��I2�UL��X�Y)���հ�����g
(�J9Q�L�J.,�Bi��Rp���,U������x�����~���uzȕ2��RoBV	m�8e�k��dt����ُp=sUQR�$�>�ȿ�}5��¡@�~5��V��Z�΅D�*C�����I��`	��׽� ����@�Bg���&8�.�.G<κ��iá�5 $n$��
�D�N�D�O�1R��ً&S3O����ڵ�����~��08�(0{]1,�f b�|@c�H�Jq�^ºOir���z���L�^�]3(��fG2�d.b`p�����3��d�S���pTL肽���b��0/�C�������]&�;1�l��(=��pO��
�Ȏ S��#4��_��ޱ�nķ��>����]��wD]�ŢG�*��E��T���~ϗE���wH��٧~��zc��ntXV�L�*�~U��Я> z��Wf��z,�
��!�Zj���E���'�D���:ϼ����I҃�cr��C����]�
����� �/Lȉ�,!�r�_J�9���Ћ���sJs�3�1wcI3�.������y��H�Z��_-4��ɻ̡d�t�v�i���X�%^u��UV�A\��8�>^z���jQ6hi�׹�4a�H��2�'s ���Y������P���U+:���Nv�k|��h�9�!S�;5���Mv���?���Ҭ�nd��Q��{�lb��ػ�]S�
�����^�QQ?gxj�/��׷��a@�*�H�@�����8ؔ8 q�^��e��;�_�Ƹx��������E3���P� }c��eQ��I�쑎��q0��F*!��#�ϼn�O/Y�Ի"�����d͚�l��6��TQck�4LN0�+���~n��XW����}oR��޲����u���1M�'�.ܰ��"�u�����$�7Y�9o_�X�19�,ó!��j�u��' `^5�5�= �35]_
~9�q�9q��C���wb3u�覼:mL�,���m�A�=El����Mi��ԨnJvK܉��wP-��^�>:�Rw|��9�m�nȎ���n�Sb
�����4igَ��j2�U������T,�l��ݸ��6͏��`��jN�E��b����XX��u�|=��S�$z~wP��N�P�����C#Le�ua�U=���{"Nh2v��K!��}���Ă��x|���QWf���'n&87��(B��k�T�|��dS���d
}*���u-xK���5��yL<^�ō�r}�anH��	�˨��; >;�~�O9Ը����t�wBk�b�X+�cg  ;f���=��Kf7Nş���ƶk�\&�8e�(E�[��\:�
��3��E�>�p��k��@�����Rv��F�\E�c>=<��I�'�&b�A�[q���w{{�&�:�%�J_PpK"s�a|M顦��b�:�Uep�R�;i�n���<!TטUf*8�˹Ě�A^B��]�p�3<�&���iѧ�����X����tLJ��Q���(8��'��3&����Dt�ɻ�\��^e��	:��=��krt������{ʓ���T�8F<���VK����n���v��U�� �*H�P�$t�A�8���*���q9n3�:Tj��0���=҇\B�ю�1�b���F�u(p
��Jcxs�y��<+Ex*�n��G�����5�5���ɢ�/&�X	5��1mb�lLC�ul� +��~��,T-�L ��SQs�t�5��;I�5�t�����`Mr�5��ʅ��<h����S8�5�N��}r����i�|��q�<�@�����X�S���;���Y����jS4�kJ�������R2n�x��g表�;�T;�׷5�wl���q�{�ᱥ����Y"��9~�P� gN�����^��y0�������l��#�-G���ϸ^^"�D�4n6�M�Vn��@t�%�Au�u_%�~G���ɇ����{�vC����`�C�]��t�5��Z�܃�aKy6�;�FJ$᥊N=i���q�l��*�g�+5��5h�5�g}12ۮO���鞥Rq����օC�8D`��lE�ڳL*��sb�JCd�Y�Ǹq��ű&�gsח�3/x�a�?#�"�j�j��Y�J��*evOʇ2�z+�14��˪�Ĕ�{ME�ܑ~#�WT-92ނ�RŪ��D���qP 1t+Է>5��j
_x�Yj��O��Nv�)˷�ٔ#h�U���}�>�i �#+�x��Lf�^�KN[���c��v/��E�`���Z���A
kښ�n�G_�t��5���La�,"XK��&��^�L�{�r�L��`�>U"@�E�tⷐ��Ys5"ց1���k�W,�g"�Ppra#F
E�!��;���ה��Sa���r��St�v0��;p]45k�'P�R���m;飪�,<1ֶ8����EZ*){GbQ�Yt��4U%������@�64`sz�$d5��{}�a�ր���:9�G�=u9ŗ������h��ZlT_�� �U�[���=��Z�8�����D4~:�T]��(��\O��x4:�Y����7�Q�bܶ�6_8�Lpub٦lOܧGݒh���ET)��p��
p{�-kxj���i�T�T)�EZ� �"�a: ƯnMu�K��/2��L¨�����
��Ü^���AN�қ�쎊�|�Y��S1ra �w�Y���~�:��BZ�ё�u�3���fh�d�����.�CT�a(��ۘᚧ3��"�M��L̒08f%w;��@��4��@��.��*����Y��m?�7:_��1��͢b����C�ʲ/{|�ê�,g�~0�cE̑ȁ��:��`L��´ t�gvE�>�̔���[��#P�wj�YD$K<����Q����aj�b<��G�}nK�٥HQ霹w���\��t��NGz���u�J�m�άz��`�YJ�b�����=AV��0O/#O��3Y�0����s�jv*�`#�+�3��&MgU�܁C�#���9��-�c�L���&+�Z��E`������G��d�7#�j����wtF���-f�h��6����~L�ǼK�P ��u+�g��6�rk�Tp����� Gi#��Kf�	��U/� ��8�ry\���!
G��s0V�%�DX�[8 }5���W���y��B[S5���<�Cuxpb��>u�X�L}x�VK�3F��XTs��U��7���$f�>U��t<4X��:�,-}<��g��t�G�S�RP�xӸ�iV�h�PO�xGʵ/�G���}�`p,E�'B�&�,���9���Yʦ�N�;}t*�٨C��A�h:6[�.�*{J��E��ƗJc��KbNm� B��I%6��ڳ)�2#�������[�п�YYE�V;���w�;���ѳ��(J�� ^h�	��Ӧb˒�+@���n۔,%��V�z���z�U�^5�Vy>5 ��
����h3뛆���{=����t��i�N�ߧf�:U�a����'��$Y,C�ћۙͭ�k��GiA�W1����GF䡊g����a(����z~���s�!����E�AOԨ��1psk��Z�V
 P�ٙʚ�M,�tq�>~� (��N>A���@o���zJ&��o�G�9��m��D�؅Pk�C�)W^��^Dxp��00�0�}��0T�����fk毐�L"[ r>,v�B�юȷQ1�,A��n*�ꃙ�X�R��,�����&:^�Tp�a�BEi��ɣ\�|��	%Ƙ�S�
 ld�Q��Lgȁ�~51]8u��^�J��q�b��/T��*���ʅ��yQTt|f�Y͢/ֹ]�"E�ac�x��[mF:��ӫ��5�Z?Z�������v4�����mz�,��eoG�o���t����v��s��E��d����� �{P���WKB��m0î@�W}͠�؆1�ڙ�f��1x;�ԛ�t�ύn��?{F��b��{�<�����:��P@� �X��@��5��LG3E���5�*��K'��F��m��k3V� T�QG�$��ٓ_\���W=�EZ�:Vk��0VW���C�@��e�\K�'����8ߧ��'֫�&tc�\r�N��;4��<�T�DV�M6���V�F��,i��}��f�'�̉%q�G�F.O�!
��?!�G*���7�5��)z�)p4u�!Å�4��?,,��A��=[y)o&��[Z�ӌ�*UDWAp�$h�[���pl��8'�5ay��Ǻ��E��
�0����7r?n�
�D���f�%Q�ȇ9f� F�n�Mf�B��ţ�[��V�޲�NB�����b�3�p�]˼	���ҙ:�li��ǈ/�.�IP��v��nZ"��n�V����\�ֈ�>Zz���]V� �����\�tH|@���23�%����z����ƞ�p��c��ʖL"lh]3��Cq,R�aXs� ĵ/�q�10�5U����q:��	>�tۨn]C�b&e�3"c��t^�s&��H� d1��51��Ɖ&�|��g���f5ܰ5L=ï���53^��6>����ޠ�@�|l�#��P� SȌ�b7�
WP��m�Pl�z����㍈�E�]?.�"�f/�I�U}1F-�
K'4�>T�
Nu�Pw�s��9`u1J���ġg׮�kn�B�����*�N@��Ry`"��>Ӛi����4�������ڇ�G�%�>���)w�`��X�x��F�%i�a��i��ڨ*»�~�jޣ���ɪ�2ҭ�5^ 1���p��s�/�W
e�-q�\ͦ3.�L�q�#��u��g��
�G]��ب8'k��m�X������%�F��*����?Mi֣Di��ս9Â�=��.���֊��:�֫tY�����r#ne��r�j5�A�r�鮫�%,���C�M�@Tn
�[��+x0E��A� DkExG;�����jΫn�N|5*pp%9̐7K��U�w���V�Τq1�5*��
o$�-����[)�e����wn� ��E(HZ�3|�Ea�L���Ǟ��8]���ƜEZ�8I����BR��nڜl�a���P���(� Za�������+G`�NQJ�\��g�r�ѽg+Bw"6����9۷F�ϖ�&v�1j�BӬ0�up�(�z5�uIW�jT9t��W�,p����Z�ì�$�]W�e�g^��e(���z������ �Gh��Y�Ӡn���3��y�m��u5�}�3�,@_eLQF�v ؔ����.�v���=���c&ݓ��+������<��!��a蘈�.��n�����wn9�T�v��h�e6��6�f�=�Wg\�C�������a9�6�s��W�2�wD�:4�.4�X�T���J4wnIFd/eK'��-�՟[9* G���hPnś�]�2�����J��PG��N��_�B[�,KvTB�=X���r�Ӝ�˗TP��Ae����&�|\�»�T((;]4�Қ����0���|�����_/t9���A{�R�]�+
s:������Đ��"H\m]��0sw�]����%VR\f�&�֑�.�m�E�r�5;.;4E^s�-��h&��[Ib|n)�I+2�Х���oN��g(A�#\��V��+g]�{�&L��gm
ֈ,��R�����%1y:1���=)Q�As.���v���U��a�<��1k�}/o�;�5A,ޮ�X`R�&�Zih|��69�ŕM���y�!V�cSD.{@��wtf���+l�E�e�F�Y�e�n�A;�W���rU�[b����E&�nt)%�t�ݝq�붹62��f���u3�;>! ��-_]���:�e�t�}�c��tE {�����U�kx�Z�)l���/[�p�J�,�����BC(�΅A[��e�#h�d!���Y�$*��B������
��%@��Y	ȓ���T* �)*)5"_�۪U��	KV�F%�"��"��K�*�Ri
��r�J-N�E�adRI$Q�Dę+H4����haY	�5�D#MN�59Ө�J(H�$Z�E���m�LL�9q*1.U-
(��N4�V��	�!AQQ�N'ILC9��:�������B
YD��Ep���$!"�C�}�����u�<�lAIε�<&��c���%�cmk���5g7}�����4D����
���|]ɿ:M�<�#������w�<&?7�ܨ}q&��z��}��Cϫ�a@��GxǄ}C�|DB�;#�fP�,�w����4���I�P���u�������Ƿ��0��~��𓴨(U���=����pO8'y:7����$�zw����W&M�����y~@��|�C�E���1"D@��ޏ�zBN~��{��|v���@���~]؟,��}���S���ݗnL>��:�W���=FC��{�z~^��΃�DH"",A`��������m�0�� ���{Bpx�����s�q>��';N���/�<�av��ܮ��M;��&�~��DDA��������}4�;.S�%p?w�7�<?�=jۓ�진���?#ǻo.���>w`D߯�s��~ ,�����"�"��X���#�7#:nS�^��$�z""��DG�ň���I����ώ��s��()�C���ߨO�oi�.pra������~����I;J��|���\��$D�8b��R�˽���} �A��)��$>&����ro�&M���M�	0�G�< �?����s�^,�\}�~�I��"-�}'��@rN�u>�V���u�/LҐ�R
F0����5��+�u¸x���C�F'�!����@�#��&����&w��)�7�$�P��>��9O {I�t��E��/=�̿zB􏾀"?1� 7�i4��o	����ߺ1 yI;�ߏ .��8�~��%v��xM�O�|����0�S����]��>����X�G���u��=9W{���@&��w?,�@Y��@�vS�;þ���w&C�<op}C�ay��xL.�=�S��w�k���=&�=���Н� �����W�zu�~�,�V6�t^�.�W�J�2�*��,*/��V}�q��N��%^��
h��q^-�x�U��6�<��seWڲ��'1��Nt�[-�-e)K�L��*�l��k�(v��+33nq%<�(��a%�~���U������|&�>;rNһӴ�_�<����0����Ԑ>$������C�����]��M�	����}:�>� D}�\W�#HK���^����|��O�|��\{M�!�ěϸB��aP��i���%0��>�>�1��ql�}�y���B+	'���c-O&7��eF�����c��{�y^�K�,o
ܩD٠>�G�V��-�xk�8ԩ�h��M�����\.��h�W�	& )Q5�q�5,t�܃9Īv�;
6����q��i�p�T+�(,��I"P*�d+V�zO,!�<&"�cjUD�a��Ԡ��a�<���ҭ��?L�K�����w{;���@clq9��jaMګ����e[���� �bw�P,��WB<�x�2���R�C�b�g������[0�F(��=UX�|�C�/�j�Yȶ�=��u��yS�|��n�RT�.����v�c����D�;C��6��Щ��J��M�)�铲��d������7����-s{��}�'���KҼ}=�Z�x9���2o&��,j�q%�Sn�	����(Ļ6��&w{c/r�o,��HR��Jzds\nV�ah�*o�>"s%�K^�N��)��rǪ29F��0�0b02��^����A~��hy/�U��3�H�Q�uG7j���g M ����%�n��	؝�c�\�yo{E]�t���WV�O>>�H~�;��vhJ;鵂9�n"�1˖g��OR��O�ڦ6����҃z%	A[������\O�{z��V�D�����v���a�5�oVcKs�����:��ϖom>�s�@�%{i����.���(�&�g�Mc$�T�+�����Ý1Nʜ��SlQľy��<�d�׋�Lv\�*�A2���J�RmZ�{�X�:�/��x9�ƱJ�+E.��ױ��.�wb�Az��D��{�f��=�Y�u�5!��U���a�_?��ڏ��V;f�K�+�������EU�A8[�I��v�� �S��p)5�WoWD.��aj�?�9�d���P]�tq�]�B��s%�g�'�p�j��Q�<f�����k*��hR��n���s��a�C�Ֆ�=�����}�{N�55S�3lÖ�(�L9e婉w[ڷ�v��&]�rٵ�k(]��NP���z�y�0v�k�^��ϩ;]<�`��f�3!�q;+<�ە���ȼ���:�S0��:L�V����jW��@g}k zfw[�7�X�C�J�=���zq�m���P�E]�7T�w}��6���6����cD���S{vn�����!˷�V�E6*�aU��!�#ǀ���R���yԟ3i����t}��Y�ڮ�G�W�6�uJ�6k��sO���}X�>zg��m�y�V{(��E��o�����U���9���3�b�:�������?T�H�UU�h�xOtV��֎m�V�`��cHҚz�տ�x����Mӥ�K~�=�S<֯>4&d��@�ޘ���MyN�׆���"C��Yإk5���t.�B��{'�rj�v6 52Z��J�@s	�#}#��Q���[���M��Z�p�� A@�gu���x��F����q�Vj��j��v4��{-Ī��~�P1Z��Al7��e��"q�M��m�P�?�^�X�Ю.�f�ځ#����翼����@�����R�ۈTXΫ�����q��y(YY+��q����Ħ��怜�R�jF�]�'sz�����$����S�^u�t��O/fi泓y�����_�'/ m�@�u�񚦘ه�k ��SK����(΄~Qsx�J;{���v��7�Czr�]��Q�F��n�َ�f4G,K-"�c�b����d�qS�K:�3�O�]�>�[�Vė��_���{��2���&?H��^�t
/�4���/E%���鵘�y
�Nn8�ؓ�g:ioV�Z�8�˰I�EV�c��0���ٞ�y�+)�+6�h��-��^�W�V�7�� ���z��\��@v	)u/Ot������5���f�oyA���i��\���^J�,�����R�=��B�˻��M`�K��u����Mu�gf[�X�~Ȏ��4�^2ߝg����.p���H�V�n�V�,�J���n"��b��A�N�:yh�;�V몫Č��W魲�5j;�\��j����XM��q+�6cq���g�F���-��ȫ9d/��P���ڝ�;��{%�Pj#���a}�u�Jʫ���OǲA��A�Ⱦ�}�ƴ��v�K�����`�!�}_9E=q??w�-���,�}�r�ZG�x9G�%�Vv�]��{��5��cʮ�2�n�J��Áͭ VFKg��v��r(S.�"��7��T����Ϙ���ia�obA�<�I���?l��,�r���z��t4�I���5z���"�L�8��۞q1�9W��>�XV�*m��:�·h)\���{��r�$��b��^7�/�Fpw��e�t�>���֧C�k�_��@��Wùu��9�Vx��&���/��Z�t#�*�Գd]ޭ��S���F�iyP�NȔ(�\��ۚɏ=�����nNx��<F�g���Q�/殐���~~��Iw+��V���5ښ�kҤ~]}]i8ߗ=�ʣ���<��(/{ik�ӫ2I엵s%;|Ӟɧ�5ƻ#>��W�5�]��t�<����{yn�P�ڍO�Yt'���;(����n�ӯN|6{y�����e)�*%�]��l�|� weJ�[m'G%��s���rs���pUFE3�9sy�=�/���������Ts@j���vvf�Z�
N"�+E�Эv�HSØE��\��Z��E���8���ô$�v�{r�L��҃Z��D�ΰi����c3���$������_�F=�TZ�#0C��Xd���^'�SBo]��BsE��(�޺����~�菧/�y� o���+�35��bѷM�Q���u�Ϋ����;u�������
)wo��!��A��-k���sT�|�w_?et��� K�W��n���8��3`K������U�uΈְ^�������K���gzMO���}��t{�~��N���5�x.K��r����V�ݯs�NEzs؁^�n,��^O3ب窄�(���_�t^��Gמ����zl��Cu?'0.2�t�;�q�x���n�9�}èq�;w����V�.��z'�����l�I�M%c��g��e��2������v�e��S`�Þ�=l#^U�J�f�Ln��x��8#����&p3��nV�<�
�A��<� ���ja���B34�%-���-�z�u��s�O�)�i-�着���'y^F�\%aW#)Jr���PSkv�S�{˃��T�J�v🷣)A��4�q����g~�^�@�f�A����:. ��݊�O^���D��Ba��	UY�Û�\E��Kp�^Z��՞�g(Q]��>��V����`�j�� 6�޽t��#��P�0�d_^��eX�Ƿ-�5�Q�/�����z�5q��TvͣN��\�ݹ�;��V�=��oA�]:�c�?-�-���7��)ةc���y��N;�Q�,�6Yֵ�2?I/ӳ��%mС�U�q07�7��e�p@���<��<=ae��ۙ�籗S�5�ۻ}É�܃^KEFd�*�igv���jK�vzS��m
vy�-��3��5k��u�ZR���&n���@D�7
Q=��Xz�Z/���Vή����=����lì�ڙ⩵5׹ٛûJ�ʝ|�)��)��'m��-���k���]�ܧl�(���R��.��O�eJ�E��{�,�u2���/!��*,M��eX�u\�Ԫ�d�Մ>�u�9�%��S��u�y艂A�q=���o��v[�-P��tO
�
��W�l;�G���<��|�ޫË�7:�MGt��>�XP���i��-�y#�q�n��A�-��ޛڄ� ܭ��L��
76Ҝ-��\�r�et�pnPgL���^��慄*�a�1�+T{�\:=�S/kY��apћ�__'���t�$�m�4�o�#\��Ji��%�2k�=T�Y�����YH	��ý��K��2#W���zy�Wo-�[�g4�u�d�#�9"�c��w�Y�XP��s��5���v!wr�(�i�'>׽���mn��&���(Oߺ��:?�W�:_�Ϸ()�[v�p���=m1��4�A �)ݐ�L���ɢ$�`閶�X�ֺ+�Mށ�K���k��M�5�pR�p{��.��Y�ͮ��%�/5�(z�=�:�=Y�o��9��ڎ0�����8fT�':jD,\����*M�6�0P&d���{����Xi7�vF��x���1f+�yV���C�|�nZ&�qu�X�}��
�a�"Ų�YM����<_[�ȾpB��o�ٻ��sU���,vOԘ['vz�P�{M����ok)]ip�}(k-u�d%����}2���FP:k��6�g<R��+���>��2m�r�YV^�Z�` �L���w}�o5�C�b��:���1��i�-Զ��Tq^n�k�Fڻ0�htص��v�gVR�8���V�e4;��W��#x�j�mK�o5��R[Q��j�c�8����)��B���E�;�4� [X�i6�L乂����Wi]Z�ͯE{��1��߄@ �Rufĩ22�L���DT���PUDr-L$�ifEmdJ�LDᤥiWRY�L��*�"�"���E0�L�9�N��(E"�hA�mPШ�+:t�-D�+�$���:\���Ad�̅�50�)Me� �#0�H�(��Ue��m�A��JfhV!(��5�&VL��"�$4)0�ԓ��Ih��d�%V�E��vE*��#�GY��euE�!j'Mh�"��B��+$9+.�I�*�ZӐ�'Qe��?���Ϸ���V�L���6m���ޗ4��<�Z-�W9��S�G1�����O�̗&���������ӿ~���v��N]���T#^}mM��g�k�����=������B��Eң�f��Wp~y���j��)?%���zT��a����Bm��y�+�<1�^~Gxg����n3o�ɥa5ܹ�T�!�s��[�М���MJ�+D�V�纗2����9��y�êX�"���4�۵���M��8<��
1��8$��\.���R��6�;��Y��pb+�1P{f�ۂ����R��-��iH1i:��%�s��["o'P۷���7�=�{9`�����=+�v��zB+�6��Ϳ����~m�����]�|�ng;'��஄J�':���Z��WT(^���Uu�׹!澺���v�(���F.݁obR,�@�0�T#��r�V�[YOz[ޓ&�⪾�����H�����v�
3y�_Fsam\�\S�m� *�08�
`Tޝ2ռ�\κq\�wo<,R��l�q3�2`l�l��7�R��u��_
>�
�ϗz����ٕ�tw�"��ED//DMz{�)��8g��Ϫǧ���'	�5Ssn�~������\��A�BO&�[��3�C���(�欽K9��4��j=L��QeM�����uL��	^��ʞ4տj��a��J��i�N)����W:����Dg	�X��ov5.�>���H�?>j��V�vm�\����6��/�G¡�s��S��o�[2�2d~�Y%SE*=V�Fj�!���+:qq����άVM��s�,�{��%�<9뻣��p}�щ�0λ��k����;��3�\�\�A�I�D}����t+������wm!ޕ��t���K��r�;�	c��~���r���D�f(������٣��[��
&A�<��PV�.�-��M歼�s����?u��x�eJ�0�4�4��T�2n�]�H�8�O�B��3G���H�9j���E�x�Ž�qk���w}Z���
��l��ܝ8����V��py�x���W�=�d�-Oj۩���a�ig%`A���1��U�=��
���Y�gQ�[�9�N��ƴv,�{�����c����Sz��Ш[��Z����V��ܭ���j��E֛��F��|�w��o�2���W]
r�h۰�Z�6�VR�휅����7I��S��<�����]h���if{y�ң�qcx��˫kq��-��kZ�L�]u{�Y3�;C2�3�}��m�-������X=X���+�	�=~�fv:��!�;R�n�7W�dlmԣ�8�KY�劻W��v�%7����}�O3[	N�T6,��b�R��޾����pه�+�uQJzyu�!��l^��wj)ش���zb��mm�Z�����T�5DK��ykjs[��<��̍�wK�g �p75�\�.��y`������m�@6���)���s�����r^~�jWz�N� {�����<�'���M����pk{+�qP҇_s遚z��s���&�~�WW������ÔLr?,LWGY=���*YDv���U�أv;*Z�n��N�ڐ����v}œ������%�٦V��d�wSA8�q��uu�Da"��u^�?�fӔ�yY�ǦAյ��IWLg`ML\�����D}��Z�7���cbc��F}Ќ(z�lс����;�m�{)8�T����Db��5Ө�y����a�f�	X�or�Κ��y��1�(ֹV��0�ͷU)6��y|�����MŽ��";�|V������w]��U�P[d:|~]R�m����^�yOI�ߩ{���>ij�ץf[h��mL�7��8v�>no{��}��g�b��E���!���Kv��TҜ�͹;_y%Es4��W��>L�s�wFo7n�O������Nna,"�?.Ψ�f�e{��v�m��Y/����k�!�T4*5�����[��C�� �tw���p�>��H��e�~iL{é���F�r������ʶ���#@�MsR����*&��%�z[���T�Ӕ�����7q�v6���RȌ�s�:����>�ﾈt��t1ocNB�}])=�GoӖPV�,JμI��rw��T�E�t:����{��u�:��5��U��`_nv�;^]K��#�q�7��Ӯ�:�9/:po�rN�g�r�q�ja�*�8z8��5Ԩ�@Ho;ܔ�WTuy���_0fه-��r�R�ChFƜ���{��XLl�uY�ji�y�������qM��y��ӵ�c��G+�P�+�J?��@�J����Ցc�^Y2��E"ʯEh�PNk8���h�Y��Z�#��RY�.f�{�'5�r�Uѻ�;Vߐ�B9�=[4d� ��>�^������M^T @��Cn���C� ��V��;=uR�����`H6��r��� Z�z�&�?Pܙ�4g�%�`m��ϵc�'�ﮓ���<j�C�N��^f�dr�gFl6����_}��}T���q��r�����T����*��|Wnk�RkV�oܜ^;��+c;ջF�5��~O�=�kZw���,.K)�;��gWL�
���ڡ�_5}��R'�1�X�|'Vۊ:þ+��h��"���a�:�Ln����B��6/z�߹l�Q\���J��˧p��/;�zR���>w�=Q���Q��l����$�ZK���\58�P1�t$��t�)�n9�Ap�=�}�Vc�|����pz�lJBudt�A[p�o&FL�O[Ow7\�\4�Cو�Uw��e��|�q��u@VZ�|���Z<����P��[
i��)�z����lڊ��Ŏµ�gN���,9�oS������Fc����emz�DU�N��X��4�u�t_^�*YJ��hwfv>xX�p��"]��pL�(+D��G�tD������>���=����c�.a����;�>���Fm�Y��_�?sVW���t8���1���1��ij��
�YjMi�	�b����xF����}	awY���D�9�<jz�c4c�ӎ)~Į��CH?^������zs
�T�\U�'r>�'��^�+�*�hx6��G�e�=x�mS�V��'��=�{wf�uL����s�~�u�uu,9�u���|ME�M����Ҕ\��_�{Y�F�[����i��k�+j\���^J�,x�Ee�f�̦%�o�/��o�+
������y.-���5{2�W0��U�ɍv�)u�C�jhFCVgk`�� i�n��;�ӫ��f�u�#��02�X��:�y�h?<��T��bo`�Sq+U]m�9��Y��ڽ����J���qZZ��N;c�C�]��v���>���N֤���t�}A���d��tq�qT��B�P����N���gWS��xӨ�
7[.뻍�Y�����b�4R�5��9|���k������-�}�� ��,��?gx{hH9ձ˻j��,�Iu�Y�͞����7[�(;-��TLt#
jS�`���o��fU�ʉᘏ���Nu
���c��w���ع����S'�]�w��l���Yя]���9u�)'�{s���Hmi7�>!y{d�	��=u�5�;�S�{\�1u|�>�ޘ;�tTK�(A�w�5��Nn.��}�_�{+���O���(��V�d5�{���{Z-v�`nl�$���$��gDpeL�&+2�Ք:ɮ���x�z���{�/|�=s����Ng5.�]��b��(Հ�}��v�ȫ�'�p��Nq�����}�D}��u��bg��~��8�q)�~\��zTz�Xb�f�&��y�G���g�Ҟ?'�eoa��3�ۘ�U�GҗH��dx]��qz� ���oZ
dvgv"�9�i!S�Ϥ���U"�j��
��3���;�.�^>�zb	6�s����U�ew+���r�
t/EKl���5�:9.7�������s��=�Udnr�ap}��y��w�b��dt��[�z[����«�U#�R|�y��kA��7�\���!�p��J9����y��{˟�;��5W�>���	��L��mV,�ows5��j�7Y��M�vy���E�_���<b��O�k�x�˴�H�&�q|��v�g>����(�T��j�(�aޙ�ɮ���ۙ�oy��t�8.�qT�%�b���%�u���.����֪����������OF�8i}K)�����D�kt��Y�mm���Eybd�[9�"��G2�=ø�s���>�q�w:�:��9t�%i\���%>��#���՞MT�2���+3����P6-8�n��1Y�����k_�E�7�Nc��/%�:ח:��e�B{��((���ǉ=⯂���)��
��$������Z���<����)R"m8s�:��EѼF�mw*��I�n�h�hażS�#(^����G
�E����#{9uv����U�M�:�a����x�h;��:C�l�|�U�ʫXT�"��\�去#P4��Pf��rWZ��4X.&��u,���A9)�w-D!��oZ��z4�I��!�5nLM֮�{�2s}��CD��!��#nx��g���Фk�ޝSt���iu��Zfa�����-�X�\�.v�Y�6�"\��!��ټE�y�qE,��o���)�解���)��Jy˽�F��F��=������6�Yc�T�=�}�Ց;D;Y�%YNn.�&�47��	�ޞC��w�1�h���'�/U�j��;�w�������ȩ�e�Oo�PI��]Űۻ-�jA֧j����n�^��{	�>"����p\��Wo����Ǯ�o�7���<`X����Sc6�Ǜwt*+�f�y�0�`�zb|�ͳ�k櫮���
�Z9>�s�I/	�e�6[�w�P��;�mٙ��{{��aň��v��aCڻk�KC}�ݜ� )�V��D̰��x3���#�t��_^	���T��7�^�z����e�=<���,V�s3Q�O;6:��N<�ؼ�
.���'d'LUf�8��P�;���������~~��Q�}B°��� ,)�g�T9Eڕ2g[̮�2⑳a�w�E+�=l��K��Qi�2�h��e�^�w~�ោ �|@ ���-g*�V,�*"↝M��:L3)E:]Nj�Q�g+��A�	2C,٤�A��,�k-L���E\m"�0�%�Z��.p�D
���Ҩ�YQʌ�hT���\8�,4�DBT\�B��$vEQ̌#9@\��(+��sHT
.��Yȋ�2B�	�(�&kJ�.�((�M"�2(��Z�$S(�#�Δ��*�%i�ȹ�d�HU�[T�.Qs� P�Br5\9ҋl���q{S�#eF�*(�]0���'L]w�#r�jw=w���y�ܻ��d��[�g����}�}F�U楮l�!KZ蕣6�c&��Md��}Ԉ]e�rz.�c��=y���������.R��	79�ɯ��7�]�}�n�U2x��~y\˸��BRu��o�v��.h���b����㵝���Y8�4���c=�z.u�)�b��-��G�7'b��u��\��f�z����`2Q�?��Z��Pt�{���G?a�!|b�N+u�W���<��ƫy��އ	e���r��}[�_.\�t�#zȇ�u�@�OV*)50���abؔ������4���&���8�X ��
d%0�˞���(���ۊ*�⤵޼&hB��Ew='�n.ྕx��q4������j�b��4R���n����2oV�+�%I:	0]2�����y�h;S�}Z�ӽ�V�Q��]�p�����W�U�RI7��h���]|$���8�?�V^����l�}Ф_@��=pV\o`��+U�@�g��+G&�=w�����(��B��PwҮ�:��S�+kz�˦���Uoz�N��t�������-^�MMD�kj20��Wec�J���=8�Ԫ�wQ��:F��j��s�������C�fLۋx�7�J����Dp�kE���=jb�����jhm8�9O:�+�(֮:�~��+)V�ar��a̍�f+XǱo����5QF�\�e_&��Կ��W��`�ioX׹�]�&��?ua�ͮ�ߞ�>��Q5n�#(�Tw�w��[y��]�8k��e�,��f�� mҫ��Ngm��)K\�����Ҹ�b+�E�Аc�
��&w&.o�/	uԚ���Vַb�^8o�����Yp�޼����W"�_2���s8]�'ID�]E3�l��
ޫޝ�������k_��x���٣�)RV�@��C\����Em����r�&��W�.K$;'�ғ�]�o9-�N$��~���5��.�*��%泛�5}��������pV*25;�]�.�uNEpV�;�Y΋�\�_@��Ӝ�~���V�}d�m���8�z�{·�Y�19�z��씬����:שgs���A�s�k�܇C��>�5�ݻ̹���r��M�Z��O�C�L9���5�ﳦ�)-�.^힂N��a�Z��[����5$�3����]ϒ��������f+f�Ǫ3�Q�\_;������ƙ��^ܨ�LB(���{�n��s������t�bŐ�a��m*V^ׯ�.���XEѸ[<�y��2L'e�r[ƹ��DG�M[�����)Ъ�06tܻw�o����� ��d��ۤ�kok��5���ge���*���ރ�a��se���񗜪;����q���I�1/���4��3��3��%�)|�q�ö�QewQ��{�ԹӣV=�nwx���b�9^ɼP�T�qh;e��hKz��8�u(T���^>�:��W�����\3R���+u��
��m<�t!���0k}��'�P�+t����9/̽���G=�'L�*}
�'�*�S�_$�rе��OP���݁)B���m� ��w[��qx�-�C��M�*6a�<٧�B$�5�� V�k.�Y�ŗ�-��.������޽��)t����" �-b�� 浶�Mš����WU���2d��ޙ٥� ���9�<뢩Yu�^�|[@��b�)������k�;��G^����#�u{�����z�۩r:c�7�$����R�{Z���&���ci�W ӇЏF�Թ�n�����O�{���M��ǥ��*��j���P�n0d�ז+��j-zQ]�����c�����*Pz�l6�&
ֺ&֍�:k��RmDý��楀A�V�4�Փ��w\���\yQIS��mvszx���V�N�y��:�]r�ۅQ��u�.I��[�����#�ʩ��Z�+vf�Ƽ�V��C�=�w���n��a~^��{<ӓ9y�!Xΰ���܈^^�2P�L��d�S�O}΂���sحS�q���/�;)�]� 7&u�Ug��a������
�#�t), �v������K�m/��������^�3��3�}��W�U���������El�;�ԛU{JI#��8�TOk�Sĝ����_S[��s��v
�+%�K�)'�/Yq�姥��4����-XU�i*���)�o9.]0�瑦7�Y�F��7+��,�
�&ҟO�רk�P����ܪ�'ީ��8��I<ۯnP�;!�B,�Ǯ+T�M#��q�����<�P����p_C��}A��Ԧ���`�d���p�NE$��0/jZ`vsa�����E*��n`ں7{ٛ�:���]Fc���G�*{�7���^�w�/(Z=<��KًԼi��P��=��N�w�Y��D��巶!�grB�6`�㞡b�GF�9s;4J9�a�]�o�l&�O,��(���iĠ2��]B�w�8ʏZ�,�|�97��ӵD�t�X��'�Q3��;�dm���&��?}UU�SĔ���U���9?R�V(S]�(k74 c��Z��7��͌��{�#c���_F�u�V���qomi��n��Jsy7s\��<��mۡ���e���M������k��[WYװ�Ltm���Z�ql��*o�P�.�zlUFq��5u)RT�����+��Ϝ�k���*�nQהt>Y��B�����'����gv3�����vv[3[%5adw(��@�����x���0㯦���
�8�Q�#�݊]YCUݝ3�ݴҳhfŰӠ��尩FƜ�	u>�;i��E�s�7U�+�1�`���+�C�g�r��"�Y��u���ժ�+] �r���[�2���ia�=wdK����bE��N#p^����c/��};���ՏW�}_|��Ν�z?SG���n9�n~J>�9ϥ ��lf���t�]4��j~r�i�?#��eF�ol�����<\߼v��k������;�*��y1�ep���H�n)�$p�����c7y,�Vި?r����f�Z�{� q\�n�&�;U����1�tc�u�kLw;z�[��ԥ6�+��위�>�]���������W���ҥ�n7����������0��!�f�����Gƞ	���:w��Aq��W��h�Nn%�{�,U�����7��9Yg�ϯ�i^{O��MT|u�)��A����1^]�xNДZ[켱��FGV4�쫜��Z^{K '����R�xw����|B�Eg��ֆ���F�c��㜺����7�}�-+F�������깣��}�}�}Si�O/2�/5=b;�:Ȍo��E�'a(L]-��u�=�̕�\7�xTʺ�%О��k���
Cžn���2_�Ȭ���IE(��B零�����r�Wʫ�
��G�*ij�=<ي��1{VLm�[�#V��r�kW��v�)�����{)��ٛ���9;�����������������S����q��|ݿ���^]��料�����j�-�1�R��=c�1_vÅ��s��@=��uY�4�vx�
:��{Dm�'��y����ϫ�����KTw	g!�ޞ[^�Y�{�n)w��\�=�n�����)���!SR_JVD򻏷8��e#]B[J	��r������wV�w[M�vPW3	�g�}ïe����,�O(V����cƄ�o�<��m�I^��ggG����UW�GS��>��&Y��~`���?s�r��#�aX���M9���"�Z��<����Υ_T8�l��z۾����7�_N��J��e�[�����BE�c�Z�qq��^y|s�n�*<d���=�t�T�=;��|����zt;�ԛW����$��QZ��v�x,���㹇jb�z_Nrg�
�^k�U���m%�N�U�ڰ���YG��0m�Qֱ�^�Y�1���pv�Ù��e�G!�05�?��1'Y���?��;����PoP�G�����'��E���I�C��pu��'ξ�����$�K,V����:��O���:Mi��I٧zpqs;��	[��^
2k���IH��X|z��f�Y�ۘ���d��1��2�R����&�t�> YX� �Vq,�����ۅ���l"8�!������zs�uP�S�Ţ��g%r��ے��mq\���[zK�du'!���+{:h9G�L�����]�<ީ�˭¯��k!5g��l=x�S���2�P�Ϸ5>KY��]Ƅ��U�n2�[������q;+V9F=y�D���[XR�M�<�,f0��%�t6�t�[�� @��V��t�J�.8�r�Q����h���
:�jK�ᓑj�*��Q��l�ܰl����<��srv�ES�f퉴C�۸u|�����-���]HƳ:�ͱ��C!���kG*5gw^1�1�N�wV���k��*���'f#}Ɂpd��w����]����\9�;:N�s��[$x�s<"z�̌�����S��珲�b�a�⛚Me�\:��cEHr��lT��;�E�����w]Ꚓ�a�UЙ}�ЃX������:��n���O<��UaK�c)��lSyV\v[���f��j]:OfS�S �O@��-0��8/���H�d��Ѳ;�|����$˾�ح��1�k���^��˜���TH"�h;��-�u��-_h�us5�cA��*������t����n��wυ�"��Ҩ��ŧ	������Vk�w�|7:�*�����P�a�ʛ�]����k�[ɐ��G8�`���ֳ�W��~��l|���3'K�9�j��e,��b� ��;𻟳�)�u�[-X�U��2��NP;�͗K6�5��N�=.=��\Ս��-��Ǻ�'4��܈s����5���
��ecه$����\9c�B	�X�$�ӎ��J��Rls�1��{{J��Ph�])�z������N_s�i%����,���H>��8 ݀�����b,�ǲ���r�fݺw�"�&�fB{:�}�X�{X�������oIV�Ϣq����P��sZr��+�8_sP\�G-3NŘҗy�+�c99�5u����  �)QdW8���j�9@D&�aW(�H(4hDVd���l�Y�V�"�"�4B��	\�e�.QJ,�����9�K(�!L�L9Ò�Z��!@�
Y�H�Z슉�M��4�B�UTUAjh�����l��Ki�+J*�2�VHUjQg@��0.TuB���̀��eA(��Ds��B��cHJ�2���t�4Ԣ9�I��3"�� ������W""
��*\,����dVeG
8p���(��霈�TIf I�O�@��HBŝZ���I۽�]]���d�#�4�p��B�M��e���J%���є�t��ﾯ�k{�S��S/��"���O���SW�U�������RI�6Ax��q�9��c�נ9k�Z�����8�{����_�Pg�}�R�z���#\|_tR�y�npt�Vzs��&�k=�Iʃ�<�BԈ�����=��*�;�=sӓ��(S�u�5������7'Z��'����O2��b�0o�zs�<��z�+=7��|�s���U���X������Vm�=Z��N:p�{�ӕ�1���:���m�<�什����^�>4��ٳ��f!�{yҪ/cz���J-��gt�-J��#C���OM&6a��S^>r�M� �W�s��A<�x�xK�F���_��rV��iKj�n���x����Va�q7]7����:�eU�2���`�a9ǩv9ɮ�Pw4���������1�着��cg��<� sʓGgm�5?'��Y[�3���)�Ȯ��5�(}�U��X�L�N�p82��-���p�l��(��|�\t�iՄ9YW��N���9K�Z����?6���ל���A����=��j{<�#"�R�s�-�pbC�ρ��׏&S��υ'o���<�˗Џgxz�������
U����T`����{{W5�M1�/e��J���Fv���w%�u��u���s곘��>�{��oT���M ����׫�ӂۭ�m&�^愪�~r���Y�Z�<��G����\��N��J�3����{`��f��ޏ�)�ep�R]=��v������ᕊ��=g�a^���W3H����r����q&S@t;V�uz�[�n5�{���;�˷��{��7-�)�������ܝ��G߾co=sd�����!�]�ӈ|���^�����L�O9�{>�*%lM�őr�j|���k;�Q=%��V���Y��c	�5��7�ޜ�vM^�t�	����(�
��̮�yV��s�X�n=�&I���>��b�R+sUO���&���
-���N񼞡r�*vQ�ʤys�:�8h3��^��s��a�J�u�arݤ�(�к�Jg��u��7��Ob�
�#�=Aj��[���>Xث��~�w9G=`�^�bw���L7�X�#z-�SY��9ލ���Y;t��F�c�?G�6.��r�	���>f�*�8M�t��WI]Gh�*��om�'�-�Mx�zK���0����"m�)Ij��Վ�h��,J{�켮��&�r�y�k��G�\}Y��^����DD@�yڛ�������w�|���3z��[ʡq��z�������NY<ܭ ��y�FX5צʹ�p7k$x��S��W2�Z�tT�#���ɫgvk�~��Sy�����U��8���r���|}�0a�$)��H��쳾]S+�}!��o��R��%�9�j����j�Ϩ�WL[U���n��'K����І������zqC؞�n��S�U���[ʟ�;w(���366�T�Eֻfa�έ�O�Ӏ��|����ߔqЭ�]b��2cjh:+�&ow�Qc�������xΝ�u}�$�P���!�2����|��/G���#<��%�����=ʹR�$0�ֹ5J�sn�N�\m:�Ҫ�Q���5��F0��j�eJ��C8�9bW,D��������%�W�}_%�s��W�I$,��S�ȃf,
�ĥ�}�ЅP�O���������T�z�?W���5��Y�=5��d��j�߳���ڬ�`�w_	?jjj=�<�ש�9���9�8$���t���?J#�\}z�\OT�T��Ҕ��F�SR����Ƨ:�$�
��>槩{�1˸�0�r��y��Z�'tX�_7�����z_�Pg���+�U��I��&�nj�b)�"�q⨵3�Z�u�F�����N+���_rY�?��:�.l������w�ԧ����>��ޮ���f�o2�L]% �W�=�NnU��� Wx�K�w�jFr�Wo�D�w!ŧ㵜pۛKh��+��*
Ym_�P�>�Nz0l�J+����ute驺E�c�0�CԲ����M]ŞH��������;{�ո�[�~��5;�1P[d:;��<��_���=���^>�\�4�n9�^�&�<�$A��aR��������K�7�r�����I�j6�e�ZӚ��QqL���G��הVī��>]o=y���M�����1^�{��~���p�;|�ih�v��_�j� ����Q�P�5B�)�0���׾V�R��=��n��p�Q�ۚ*%��Uq�>=���N;�V[��+;c�1%�1}=P�����1� �j��_f�˻�8�5]��#>T���q/�����Ӧ��̋�bja��3����r�Lqa0������",��i3YtU�״f�y���kX�V�K���l�ݢ<w`tI���ֻk��(��X�ՅV�hV�e>5�Co�Lb�=��Ndd�f��r�v��{v�ޑ��:9q��+ﾨUz���O-��mdDӺ��1F��7eE_�+�ݬN^
Xq� {w@�v�+�ZX�D� ]�������ؤ�0V��7S���s=�� 2vb��w`e�<���F��#9^������WY��M���v�2����в����A^G'i���iQ���e���.���׋��`��3���qS��p�61��OE۴�y�>�e�2��^0�Y��+j����v!��n��ʚ�<(�R�jz��QW��(�k\�	�ҭ�6:Uu���&�@��^����{�N�'��eN���yd�H����E��;c�g;�M�ɫߑLu��״9^��燕e\��k������}�^�����������:��滶��V��O,Y�]L��_wv���4��}ډ޾��F�羏� Wvj���^擕ft�Ar��|>��	ucR���9�wص�����C��˞��T-��ds�qC�B���↡^����/��O%53�2m�C�ܝ�R��n�EGZ��6p�f��5�~�Ƽz�Ѵt�xh���|����:a�����P�U�w=F"j�/X:2z�����11d\�5��q����S����y}�A�A��M-d�^����:�c���N�q_sLR�+����u�8���9���m�����Y�}��r����
��A>m��2�ՉC�쥜my���:o��)�YS�@	y��r����?m`e]kVE�5��=�Ԏ7��5Q�yݽj��D`��+n��4Ai�f���)����z�3�r�����^��a_r�|���\*�X~���lc�x{哆A���Щ���mJ�\�{-�qhn}UU`���z���７2��d��͡��ӵl>���ŵ�+{���;�z>Ϟ�!O�dlm�s���qǣ^���6���+^�0�s��˩[��]��bۛ�縌t�I;��v~�ijɕ?rԋ�[�r�F�Ru�Lg���0��֫z�j���o�2�5{���'��)�V��;(ĝgC�|��Ku�
p� ��ʄZqgR��c�ؗ��M�S�� s���6)�q�9���,��[҃��S��W��y�����*���Æ�����+&gm�B��rٽtҰk���4�a�s@{9�n�6�/�*4�v,�wv����B�+e4܏C��'u��)�jGlڸ���}ݴ���F�������r�v̹FT��\����c�x��w�7��r���������[��~���U��L��Lntiu�c�H����XwS��P�S�Ⱥ�nb�,�g��[�Pw����X8V!d\�����o��$V�s]p��?�W;�e7�a�����:��d��+b5Hحf�D_���]={i^7��:,�O�ۥJ�m���6��1b���A�L�Cc���鋱Lm���5�0����C���މ�Nn���oo���a���Qp�9��s�J��~UW+"J+��zi1�=7i������Z���Q��sX!)�DI!���ֳ�4����k`)t��\C�P��V�*����Zb���]#��G��E1xÙ�/�ՍDI<����ʳ��0-����]N�gB�3lD�M���/+h,����^���׳�����Xpp��R��̬G���c�R%�3�$�j�$�GK��Ҝ�!-�m��O4u::�:�$Z;� պ&�AjӚԐN�JR�1ܳC�k�]�_U����),.�(�b���L�P.����e�&��-�y$؝c6����Q��+�
�D�ԋ:6<�:���y�b�F��*��E`-
f|��s><��oѴ �$b��V}o�c3��q�X�z֢��V)b�d��4�Ц;�ۙjҧ{׸5���W>��t9n2�I�.n��0��rW�ޣ!+�ͼy�z"HoC��T㤅N�-��eܜ���9Ջ+�pi*�\��G!�De�t]\�na�����g���ѣ��*B����.Y�W�p;ՍV2v�&�M���m�q>��Ju.Oo��I	�P�`*ϗ:�'zrg�*�����X��8�]�oQ΁�fp�o�[W�Qx��Nn�d�tR�Y=6��@с�q��R�~n�:'�.9Yy�$��U�{�6��Q��$ͭ|�f8���}3�Ӿ�{��@h��4lʓ�e��Sx.�^��E�:U�/��Me�Y�5�+&��N8WYZ�aM�lݨi�xo�P��y�s�`(9�g[P��/a&�!�@�wAa��ih5��/������ �Z"�f�0��MvT�AR�0l�"��c�/kw�Ҳ�b��٩�Uצ��Zl5��b����#�tb�j�R���lEn��Y�^�ޱDγ����v�bu�J�ɋ�|�]O����K�S+:bi4@��U�ڽM�֍�dPov�tc6�K�JJ�+y�����aۻ�,mc�%;����.֤S���"2���M5�[�]�`@F;-��bN�(�YB��:ۖ�oVN��{b픫v��W��Ŧݸ���Y�V[+zk�^Z�x �3�t����ĩ4u>7���y	��ƨ ���(P'�(�f�$ ��$dD�I]�&Y�\�G"L�%EY�G)Md��fȹ� ��*��¹s��h�UY*)�BeQV+f�*"�'eQr�C9W+CK�Qa�B(���)VS.E���ΨDTh&Ug4�bT�9u@���k"�Nr��JF\"�.M*)"+5���*�`r�Fl3�UPG.RMT5aj�,6��L�*92�2
"�YC4�����HBAHr�"��I$�d͔��QAE�Td$]��d�ʎ�$@����W5���r�A��.r�;ԫ^��Ի��Nj����Ի��VH�ʁ�5B'�_%���>�>w��;?��Ev��9F�6�[��^�/nЄUrZ�J��0_�
��Z�
��sf8����/CW���
��LO��"���A7�j�Y�Ѻڗ]�-`�}��	��t���5�~�*~��^5y��)�z��c��Ov������i���jr-l��_h��=�̯z�V�9�bm�YĲxֵ�5�6"��J�{�����LC�:z�ʍZSo�Y�d�i��ǻ<u�3sO���?k���L�	�"�h��V9_��m��Y�-�	���=��~.s{��Y����E��j��K�+7�V~�7٫��l?G���O����\���iݨT�0UΑ�������נ���-�F�$���\v0��Qf�z��)f+DϦ�c�k�dƟc*n�
I��	��tXf�Hu���6A�]Q�{��x�n��J���~����2����s��aޮ�{7��>~���Gޔ�SG�>��Cj�$��#�h�u&�9�N1`����[�{kWEF��ƚ�g�:��ؔ�.�UR�cfw]	�o]�|���p�E7.�º`r��%1ED�q'��EĹ�y�1��Q� ��ruC�a�ە5��%��6�;߮D��i*��`-�W�e���y��O<��t���2�ĕ+v�bjr�~�6��䂜����[�����i�]�{ˇ�z����ݑ�a����͐^#
ypq��lTsr��l��ӽf�i�4�[�{J���{R�.|'L�U�ikY}��J���k�B	å�Fn�gj5�I�݅�u��x��s���f���ʅ��X�m�*=͏���O�(�����U��;�h�O;z8�t�S��γ�E�ȷ86o[�o=W3�3ᴽK���eA��Xx<|��l-�̡N^��4m�Z�����{�9�}�3wSK%[�1o���n��U�e�A���q{�6�k�J6^�O��y�n{(M����K�p�K�z���?w�����O�8瑛ŵ�,�J&�i�<�7^�����c�gq]��U��q�t�i
������������yī�ϨO�ʲ2���gґ��	�6�[L���q��]\�Hܭ�]�j����xu_S]����GZP��&J����C6���A_�3}�C��>T����&κ�K@	m��͙��:����
�� *?>Z3���;���f�w�.���|سϔA��m�hx]<�����"l,�;��Q�q����Q�Ъ��_;�s-�O����_C&9�0�҆����PǙ�y�%�&�V�
��g0�9��ž�����5R7��9�y�/�����4��]ķM�ͼ��*�Z��m�5� �Z����jj��3�K��j+�����md'n��ѳk2��^�u/>���me'VFZ�I�[3\�Kv����*�Z\nU��P�2��G�}���Q3Q1�&۩�X�4�vL[�i�jGl���E�{y�WlZ�
�Y;i0���|��gQ�{-�k����n9��7�yZ��S{~t=��36���!�f��SO��W��U���~@����|�]0|���x��r�ѯ�cn��K���N߹�����-��΃zm�=�3�������^�����>�'�[щ���c̣� {[�ҭ�{U�9���%L�W������^�q��l�}�V{�6����%q����H��T���J����o*�Z�������:�X�u��9���n�����w_Ð��ۚ*%�.�O8(9w�j�=�k�9;}0_�~�=Pn4�&(!�[�W��+�W�0&[S���)��s�ݻ��lr>��W�mi��H���4��X�;Ô�ZwP6@�f��*t�ֽ��Lߺmw�C�>G��}NЉ)K�lv_%J��P���-j�k��|��d�I��[� ����R�,@V�:��#��>�Z	{ˉ��	�em\8��Qc+K��i��ڳ�y�&r]X� �eN6*��JMme�5Q/,�Ԍ�r.VH���!�Y}���d� ���H:��G>an�Ю�2�Oa;�(j��z;��n8���'Tsjw��s�c�y=�~�ӳs���^���µ�2#u|&����=�x8|�t4�|:�>����iƻ:9��RS�\�7�6�;W҇^�:2��8�x�?W��ͱ��=I��G�jj�۬F*�L�xLJ].��j*��mع���뭛r�#�#��MT@����y����mO9����f���3[%[����R�.b8�V�eNV����ιS�[<���&9<��ݩ����ڟ��;�h�o||�<_zy*���n���o�i	��Ҩ>���s96%����ai�t����]��@�䟙����m^�1��B�w������v.�K"�+Rq-o���ۻPxb�H��ș���&j*�+XWU扑�N����Wt4��{C�W���ꟺ���8n�fީ�k%8�JT>?���j�N�RL��'uQ6�����#�9E�o�{����9��=��ocOk����N��E:s���v�\Ȝ��x�^}'3ӽ[������z8��v⹘L��{�s�M��פ�WE���ۋ�JR���S>q��G��J�nC�{���p�T��yQZB����~��u.�oy�S�{=�O�����qi�G�~�X8��ո��%s֭cV�8���v�F��FYU�r�'`ν�5i�����������f������k"^��W��d�T���#�~�ty6��6a��J�x;%�@���Jvh�39v/�F��t��)j�l�\�k'�dN��]��yrΜ]�u�K8���oJ�_�C]���CCH������=!:ߊ�\mw9s-$��lW1t/:�_����O)�gk�~��S��5�O�g�t���sԳ��|���50j2(pS�毶{�[��V�/��k����o�ggSX�ﯨ�[�ɭ�}�m�3�_Oc�V1݌Rt95��Pz��)��M��C��G^6�z���yF�[p5j
�A����V�X�����6ğ���q�8n5$ɮ}0%g�u��t#���^_����*�{Q�)���-��;�j��s��U�J�@W1��VqX3M��8�)�0�qUw����p���X'�N���昜����S[O.�g�ϼ���ʹ<����`�ɫ�u.�����k(3���6i��8U��ql �Y�ʪ\��6M���>,��NS6��;�roF1��D����9p��IC(�v��[mH6�80��Χ[�z��5=c�����Pz���,|:���M楀D��������,�Vġ��t�~���gRehݙ願��8��j�u<�cn�6��w���_B��\���}�g�(D�?n���y	��Q�����w���i�#�6�?w�}��lFq��{�uH�y��C�J�U����J+��z��ލ��m�S�VJ�q��7���X��,�0��rr����}�Nut��AU�_�QQk��|��;*''U�3�Ow[ҕ0�`'?u�h� a�M�*�N�mܯ{1�\�b�e9Ԫ�I��G�j�*q����E�{c����4MWU
@.n���]��u�Jk5u���[��k^��V���@d�}\)��n���WjD.6��D@�o�;�9��l��مt�&^�+�;̀��j���eD���#��<{*������b�������{"�:I췭r{�Ѹq׭m|&�z^�:���R7S��(�=;��=^�*�+�`�iǿV�~m1
�c;B�<��ҵa�p������
O�n���+�1��n�|����]8�si�U�.-�K��`�i͝���ȷ�S�����T��ռ��g+��;Ԋ�r��[��𜑮Z��z��^�t'ʵ��[�5���r�{���@��GEq��z�������q�ޞQ��.���>��坃��D��ۑ�f�� ����~��Gx�_��Md>�#�5˺��5ܴ[WiG���ֲ���t���>7o���(J*������i��B��&��:��%����{�����7��Ku�A籼7 �wKT(ب���\s���P�4Gl���CB��Tڲh�n
'�M��9[��*�c.�p�52����*�W*�:�Y��:@�/u+�jD��v�ҹy����.��p|�*��a�fu��gou��!�ay`_k�ۖ;�`9d�i�@�:"��rtØ��8z��Y�n�A�pW܁��4�5��[���ʺ��8304�щ�ݴ���PWX�]bE�>a��&�Pū�^X���d��'�= .Y���C�FDto�]��A��6������s�{�h�
�oU��JT����ո��!>��%�G�������1�T�8l�pMk-��ǹQj�����K)��%!�of�:=O��ǖ[���|	������6�F��EQ�ngS�H�*s��8�]D�=��%� 6�u�V�ih!�׸��4��\cE�u�Y�s��}Z�5�
asӔ��X9Rw�9q�v�:y�eg'Q��9ϕjf�s�d[ӵ�ق��Gm0D��Y�*��ܮ7hb����f6��Hn�����ќU7���pM�od㆞�z�\K8��喸�h�,dv��v����u�h��QӶ�t���P�U��2����`�G���x�*aHe��WE�mǵв)P��s���J�g&gϻn#�Ƴ��ެ�KL������_R�nbN<6��D���M5���ǥ#��^��(O��8Ý�(��|b�Ƕ��"Q��:��Zn�r+��z&�^%�ً�ƚy�n�O��牼�*�j��n�Ʀ�޽��i:��\E]gQ���O�X�/m�#��y��К�v��h�+���ue�X��]�R�v.��|K!ob��m��Ѯi���,���9y��$e[�ŗ[ϴ1ݶ,�����������`.�z*��@%-�S:*J�Ь��E�,=zei����c���Ov�.diX/E�F�p��W-W��n�lG����(�5ˎ=�of���C���Ƞ�y|�St�5�q蝹S
wu�B/��ݜ�[�̦�u]'d5.e��w�� (_UZ>�l�HUd!$�3.�R�J�"��@�h�(�˂Nl�(��֗�Xbt���A5m�'hp������
)+�W.�*AI�
�D]T�����H��($9U�2�$��ò�˅PPP\Ԃ����ɤQUgNY�PJ�v���.ʪ(�e�ʙv\��Aˤ�fB��9Ver��a��숺v]�U�43"�W�r�EfPPP�dP>�
�Iw��ε�x9�Ȼ-e�ҹ�����n�\�^�q쓝�~�w�p�aO�Rh��_C�e]INO��NnA����\�)����^dMl�nҮJ�!ˡM����\�`�8ݚ��Q�<��uAW-މ�ƇI�v���1��NW�DS����c��=����%���fnP�]��eU�=)����ꭀP/���af��
Y{w��.4e��]�p���45eMu�/��f���O+^gJ�<C���-C������f�o3p��D�y��6���7'X3k��0ud&���-� ]_V�!]�ͪ��h�v�7��]�q1�1*R��SO8��+c�n�=�f����x)K�[�4�A����#^��P���*�1�p�x��ڮ����PV�;���uͯU�J�V��z���xqkx)�օ���b�V�B�����`��(�o��Y]؛��x��.�3����fc�u9��v�%]�q��'���Z�Y�v�,�t��Z5ZT99D/.��yT��>�y����PY�Zwl��{P�kGu�XV^����g�z.a�W��;^��IB��!	���u���=�蟻�f���W���{/�3��P4I�D��9�y�]れ������O��!��\�gي��0�d���b�	ruLEsWۿU�i>\�R������WW[�X������7.���(�sV��oD��2�=�J~�ʚ��Et���l��S�{S��v2\n��F��ӎ��1.N�.6
0ӭT�����bNh�F��E�qJ{�ў�=���d�S�L&���H���NPa�\څpK�d}Q.�J9u��[��	��umw*�j� �8[�e������.w81�D|87�V����eUj�K�jy�º��s�1p�è�.3
�3�R�pN�j�S�r�8n]՜��-tq0�2/��m-��w35 ��~�����4�t^�)�����ː���Ե�WC�Ƙ\=�فs���ٟ.�꒧$�hS���'+����ˮ_*��tAv>�-TYR�����#�\b��i��wc���+�WʰX�an̓Ãr*��c����Eϰ�a;��aH��dh����:�W|�}�펀}>�*n��^������d�����Vp�&�S�5-�=k�ïqw�u�/�'*����#vLg���4�0�O%��xc�k\¯�Tf9A��O�"����=��o����!ԥ�k��>U���~�ԫ�ە��M�[��e	 Ǉp#]��d��	+�e�Ƽ��5���:n�};���k�2r���*�n����b�fK�ң,���E��J��r"f�;/�<�c����4=>���2��2f�L��Ȓ|LVmڷ�������O��W1�ꉆ^��)���b�̦c��F<ܸH)mxw������Ǡ�*�a��"	��.
�MB,�z��e�=v������LfR� ���y�
����B��k�_9!��x1p��Mֺ;��=B���X�>�fa���b�DO��Q��Lc%��5Bm�[��a�_ $@yU�H��aW�;��f��-y߶�R���+��8���1��T�p��3
�9�z$�MTp�9(e�N
��u����I�2���J���| ^'�b<`/O�������+c!�`n�{�%O�a�6}ϵ��`bu ��0*5W�G�Z��u	��ɫ���fw�-�s�^4}�U�1Q~��o�}1��`�>�6:��x�B�#}��w ��/ULb\��y�c�-S���X�%�;�G������.�@1���ل唹72��#b��OP��;t"�]���Z�!�J��@P3xJ��{���x.OzGf���]�<n�c�����9t���f�#��fy5�/��F��z�O�Up
�﮺��/	��/��'ٍoz7�=��x1�c!d���Wk�@Ԍ�vW*������:ӓ����(m��e+��w���tp�t�8��A�+�����9��U�u��Iq����0���W>�2/�E���s��/&%"}F�c���۝�oW�S�T�%x�3�ݓ56:���0W�q��	�u0ǎ_
§�q���q��b|\���L\��A����nP�^gt�W\�y�w���Z�g\!Qs�P�W��@�1�b{&/�3v+5,��1�Wg�����%�џ ��j@�L)B} K$Tx�˼0��������K�*Q�U���>����$�cGA���ٱ�*p�\E�p腖1���nK�ORL栞��k����&�o�"�C�����"���}xQ[�Ǚ���S� ]u��C6��ٗ�y5;��Q�����-e�R�fэg9�~�+�O���Ԫ��O�1�'σ�}Q_���_�O�LTN�����7/�����&��1�nc���ǅ�u�O��>\.���$���Q� n��Y1�h�x������ex�1�+���z�[^��=y<+}�s���ueB��U
�R{f<3���4��TӴ��>�lu|刖�5�F\t����&a�\�zo���3�_Ve�n���^�^��Eۘ�X�i�
�GM�\UC��\=��z�<��ط��Ǿɔ�:��}j�pR�'��Z����U��C��Q�*:(ڂg÷���g��|�����	�Y�7�x!Q�lR:�q�ܙF.�F�N�Yo�����C���;�lK�_��Ѩ����RƼ��6=��O�3�����Ga�0��G���/&d1Sި�+�����!:��n�2|�E��4+����)I>�7Mڌ�SE�k�)�jW[���jfX��7(�u����*�K�����x&�����˘�gwq�9�b�Ko��j���}ZszN�z7�txUת)y;��i��A N�t���pd�.�N2���b��y�*�͸��G��a��,Q<������1
@�p#�=S�נ{���xz ��C1��^6J�"��;ޘ����\J�h��ۡ��T�Y��}�E,,^K¡irbc���p<r^�I���y�o�/WEyYb�ިsS�D�`��#$ư�=�<}�����	������^;ހ=btS��n	��hC�ʉ�S��]C�S	UO��V+&�/�-U#UP��X��Hh����uVn!�&0���k���s����A�G�=8�����d�X�] Z�#�����m������]���Ն@��a�j��k�Q���Ʉ��D*�(S6DL�k}ӝѡ������䏰���8���p&:|�o�#<�a�b�x������n,%�F���)M�!�c�(ֲ�_�j�ةU��ܮWQ�/Br�pܗ���B#n苙�����|v��o���}�x���l�K{!�[�`�}�������{,o�J�����6=��!���ͮ1��*;�7ѽ��f_^j>�|��T��r&|�N����L�z����JV����	]������P�8#��z�q��O�sP�Mt�L�����ay��{6����S�|ԡwU�u��0����NN��q"��J�Y�V�;��K�-�s����z6ϴǧΰT"��_M��:��e� 4Y<��#�DW1����KKB��8��B��d������j]1d�b��|�>Y�/׫ں��;����p�tU�TzpmLY=��Lz�gO�#f��9���)�� 7`�>��X�����>0�'�7K�/���qFq5�Ow��r�	{�p/�<$�����LW����5P��?\�~Ը�<}��1�G�� z���\B�u�*��TO�ˁN}�����kk�fdԬ���.�\���"k���6�|%=�r�o�״`Yӳʷ��ekaݙ����y<���Q�S�Q�Dq���Wx謰
���\�N^b���({�%<���aPs�I����GN�|Y����g�;��-OO��x���'��z�� /��z|=���O
Ub�	M��c���˥�~��A��9�>�O��@�����>�a�|U�R*�}'O�jw��H��mu0�sc���p+��5��U���g�z���'��w��k������N��B����;L5��+׻KG��Oޜ*��C���C�\{���+���'⧠疞�{�P3ף��}�B5��Tn*�|/?s�ʩ5[<�΄���?mի��������Tdt��6��<'ri"E -�5�Vy�{2�0�lE����0FEO;��uK���ك{Y�?\�{�Nnzl���T�=�g���luL������=/v�q��<H���׊s#���"��u���`q����8.����R��s5�\gj�,��{ObH�]۹v���E��74��VOjt8���"a�j�f!�.���LM��w2l��u����J�yU��%q�(:�������F&���l�j��	.`w����@��1�)��aY�Ū^��*��L�<9����E/z��7����� K$;��O;����c�&=���Q�Q�L�w��<@A�Qc�So�nۑ2��5�>н�Pe�[�����UC��L�L?A��3���=���ާ7��V���ozv)� !l��FŊ�S�f�*=1��ǅ�T��_������	��������y��Gv1��71�َW5f�ō�� %Mx�G{+�V��ﳵ�߽c�_�KS�P�M���'�
�NL-�T+���j<6�̹*8ܫ^�o{����4�}�p;��7X.:�F+T�QA�UC��g= �����}�X�C�3�uǼ|�Z:͇P��H��c������ W5���u��],�Ƶ�
�3����쐏Ko]p��-u�0��W���#8l��ˀ=``��{��WJ(Bv�=�"�ݥy��khs��������aam�a�'e��M�>I_v����O��S����_rj�a|��R�(t/4��[xEf��2��.|���ڝ�eF�e- >'��/Qm��B�� �w��-�En��$���
�&�-Ѭ����R��ª���lX&��[�/�|p������{��l���!�`B����L����,��q��T�U;˶y���75W1�v��t6�{˯�⽮��WI&E@���FY��R�O&:��lWL�5�I&�1�#�汤���x)�g,!��Ŷ�;�/��N�!VZ��a]���0��p1h	�[骈.�е�]tݾ�2��uԋŮ�'F���1mpgn�ۇ7��.�6�e�G�	��ħS��]�Jv��C�vȧn;�Rh�v������ե���jik�kU.*�J!����a����u.diՖ.e�-"k�=M:�fCV�]d�xYss:�;s�8�YZ8��J%��T3���e����zU�j�5˕nV�3CFtr�.��Q�ĝ�GΆ�d<w�wz��> �)��V�k��e���.p�5P��sˀ��� b�p
c�PZ����<;1k����R���3{)6�V�hc;��'Ê��YW��rSǅC٘�T}�![AE����m������.t��\��x^"�S��,��ߩ$a
�7{ו��u�gNOD��������ǎ�+k@ �#PV�A�d6X!��o�ꗵ�_M��*C*h�x�-7b]���:��+}�T�|�	`:�f󪮎8y�gMr�$�[ŕmR%9�!�*D�����km���8�:�lT�o�B�����s{��5�m�C��c}���4�f1�8{��Ò@�;�7���0]6.Df>��\A�sE"����J�9J^nR�-����;f�;Z��J�#�7"�ko8�.�%*�C�:�E��i	2��PD$�J�� �S�@��\��sH�d��qPN�
�Nub$�"�uȭrs�PF�9�E^E�H���*����ePS�"�:T�e(癄T���EEA�y�=r�%Aʒ�+��UD�G�s�\�QS�eQº�Q\�P��ܗC��G'
dT֓�hg9PjU"��$�  �>7`���*
v�����uN�Y��=Y}4�4���]�Q�X�t��(T���x��8�{�?R�4��	�<u�gZ��J	�Nj��l�O���ob�Ex����7�p�~��&��jϑc	�Y��:�h4u���wY��k��'��I�O<5鴐@�J�ꔈ{ƾ��k��LoN
���3��V��2�z�ky~��v\x*�\ �j	��$���OΝY��׊�;u�b��E��X��	�}��\��T&�CZd#_,�\JOi�w}���{9�Cі}�TNTr8�T1��e3�G�S�W��py>,H�3t��Ҽ��
 ?F=?nU#pJd����z�k��T�Fo}�����}�+��Ѳ��֪2M��K��H^����H�՞��e<��&���*�Q�"�~���M�:��zG�V=j:�~�\<��h���'��
n|��1�s�^w��o,;u��~^�=������W�=2��bl흨����X���K�qa��n�L���i|&�����4sAR���gU�j� �/��!�+݉twO��UbX{��	���T�AJŽCf�����̢}�D?h$y��&��h��/��4���ɇ^�56 <���ٴE)���i�Ѐ���"_T����Xg�<�<ղTY���K�� \s��c<iz`�1m]a��n�W���^�V����w�kM}e��C8���p'���|g�cyN�m�7���Y��yF���8�'�a�/�<<7��KUϧ��IgC�?_��H��o	�Pw�e_��x�O׮�U���L�ߵ�S�ků1^�S
�荾u�Т�f��@�s�8#�_�ܣ�;��*󚱮7����X��LX�zxV��o�����2J�\/jі�.��ֆC�ϣ2c�p2U��#=N��<˼2F���և9������X��=c���@>
�P�1����PLԖ9��{������o��~u���>A�<Ǳ�v��[.�6irÙ�����9C�]�E���n���� @o{������Zp�i�U^��DYt�C^P��L����ك��_ZU;�x��k�d��|f��f��.WY���{p����*t0�ρ���?�s0�'���{FW@�e�9�zz� ��{z:��+j+�|.��@C�wg�j��������>w�B�� ��jS���»���9#���(X�T= וw��ˌ�E�J:ԁ>�x˟P�����F_�*�S�����ow�G�$�Lg%B�>5�>œ�*�hDy��u8�a��RQf.�ɿ�S���p�(2j4�'�\z�� W���3����2L+��Dm���f��Ǟ�9C�=f*�Ӄl�M����x05:���透�񃋽UJ�9���nث���5�U�Xb��D���S L#��p\*���5��ֲ}�=<5��
��D���^T�d獏[$E�X%�qض���c����=1�-9��G)�68�A�@Mo��C* ty»�y{>���;���^]txW��pa���V^�j�aov��׀�U���ɮ�|;2����fL�K5ӌŘ�M����:2@X�KU���x�s�C1\n��4-Ejت�ż�/HvP�����P���dŢ��L�ɐ�[�xQ�[�>;�R��W�鎯��'�<��Gp�<7��yH	�ңNu������ӵ^���)��!�:3���'\���1�g�ש�t?^���9���Ň��x�<��R&	�b��x;�����������u,�^W褑���eTp�+��B�.����S�6{��lzB����bo��O��=��عu��56H&:쨯��¼;>���uz)EF�����Xg�A>��,���Q�� 1�B�d=��������Ta����0�̏x��\�P�0Բj'��B��D��{���|+����E���P��a�>�Q��.g�������C-K��_���%����|2�ؚ6,Vt�k�ʇ?~�\x"�׏���ߕ�m"���h��X,�O���q�����B�&�������N��w5�w�|x��B�C��E殾����y�aq��]@u'Xw3��˹��`��g>9����Ybu�����jF�]�;��;lK��~�vh�q!��/j8M\՛�X�t�7_�L��w�g��-f��s��D,L>�
��lS�<h�T,�*~&�����ѩ~�����u~�zǢ�k��>�Q��	�F_L^)����*�� 9��o�6�y�R<��ѥ�����Q�{��E��C8'�@u68��W�/ٷ��޿eǮg�HvO	�-��n
�N�O��^���z߷R�����P�@dT��Yh�y3��|8��Ca�
�3����aE؊�<��wy_�/��7��;�aeJD�xmG���ޜS�<�{�{��|�{�.c�\!|�_цBS�0���TU�����T���ޤkٺҰ�E�c�,��%�γ�νxP��v+�P_J����2�?5c�'�ax�{g*&���:���e3�G�
��S�����̬j�0��д �G�W&�#`���͚aØx��l�8���UsF�:r++��<�(l�]Ӿ3�$b�ބ\V0�O�-�V�nm$�vk۝$xt��6��w��1%�t�����[4�9�r�%2EG��q��G�8��s��yrίF���*= H�Bg���L*��F*=��r} ����{����0+�Q0Y�"L+م�&�f�FI��a�(���ŏ��1���qw R��?yϸ��4!��b6����w�]>�w�8��ْ��'�$B��z	�t��xn8��=��;�S��T}�N �QZ�<E��̲[,TrT_N�Ɋ�\d{��3��{�槻ѹ�#ч�c��)c�7�h�x�/L��%��,j�G�e������1e�E��zg�TG��՟k��r��>9�`oO���b�l4����k7�������{"�YB�g|o�|H�>���Zڰ�k��,�˄�/m��Y�_�}����F02��/zyɘ�l�G�@N��B������ǹ�H���S�d��d3:#io@�<�����(�խ�lt��kB��M�����u��&��o���0�P����K��}�0;2�dh�
J��/J��g*�o�z�h�[:"w;��yТדP�W%���Cܪ�kܼ<�{�h�=�Q֦R��1b}����k���'��Q&C6���z����%�����Qf;T��V�����1���^i�'-�5�e��rާT_��@`����O���uG����Y�S5u((�[3Xߏ�����W��1�s�����:*���=8 ��0�d�<�*P<fo��V�� ^�:���g���!�T[Q^s�p"m]���!~�{��diEO�x� ���p.%� L*���9"�^�=�:�_����c���%���x��>R�<��X4,W\�7%�d�}{��q�>�3s⤱�3>1�l��TM9��I���}4�/3^�ǚ�8&�����H�����G�8� W��`��؈]�'�%��\I���Y��R�Yj������(��'l|Z�=�⵲7X��W��raOw9�YwR3B��r�1W>=Cj%1�X�S�9�W��u�K�0�U��a��$Ĕ���kV�.C7�[�lit��vĚ���j����xM�������N�TW���/�G[U3ՙ����h�s̯��C��9𪎚����R��=�����F��͋ٻ��]�hN�(O�����Q_q�L&nJM��>�@��ՏY����q�"u�{ٵ�a�Z�ѽr9I�0���\,fq,�Ş��=�NgѦ:~�L!�����%��*����i�����>�ԛ���u��6Bٍ��Qg��p�=���ʶD�wNsӦ�����6F3&c}��Y�G�t\�:�W�΢�������-{�I�����ǃ�T�tN	�H���b���_Y��CIB�y;[۞g�v�}#��<?�e�~�N�xA�`���2�L ������1o]W5ޡ�c���T>�P��˨R�$�`�eC��͇&m,����/�{7[�	[���d./k��G�����]"֪:����0�ŜpN�4���YD�t�C��el:N�S�V��s�+IEA���w{'��w�)9�a����ɤn	�� w�0�v�7 # �/+q��o�R��誒&�b��רL-s##ސ����@�0ԲW�����iv\[�c�jb�=6}>c�-��a^5�h�錇�O�;W�c*�	�,��P��N���[ ~�lM+:|�T9�^��E��e�]k��5Zia��B���
} U�&�j��]@��v|<3�ԀZ ���<��>0�����9�!���j&�C�<@�&���c��"�~�ݯN��y�x
��c=t���/��YDg�S�E�����w����o���3ᗾ����.��#LؘNpWd���'ќe_{Ҵ6,�UFO����K1D�\��ȼ���x�Gl��N	�ͩ��={�B^��?.�)�4nlUx
=�CȰ�f=Y>Q��
�6=���N���	�v����m�ku�f����ݗ�P�f�c�Șu�/w�p+j6�:cMi2���9QD^���2�J
�z'u�[��ڎU���,���4L��Z�ק�ǽ�>1iD���d�<�H�V{Ƭ���S����k�Ϲ���ν��9t�d���_���	H�!�ޘVW�z�+��c՞�滝�F�L1�9�H��\�b��6�Bq�B ��(��^���J23�{����C��5��l�ɅS���]PƲĒ�Q�#�ñ9�3���U ���y�j�C��z|6	�<�G�=ɔp��	�Q�Tc��i�{ڒno}�G�j7�-6N'�|2M�1p�&=ސ}!�xN�o5.��`,���c��|D�w������G��SD�ro��+�f����G��"�q�;�'¼���1쯕X�y1��p�!���;<��<��������>����xxdG�4G��&������u�����<}��'O�.c<m���fa�-�)t�u��#���F��T^X�T W��"y��e"1�xu++�a`W�h1��{ee[O�N��(1�+4���6n��L�����HD��Wf�(�#��f57��=���h�Y:�7�{zk�N��#�)�VqV/�q�<��[�uSAS`wLT�S���e����fż�P��P�>��SX�e|���o<�ʦ����-�,
��q�f�΀�(o����dԭ��͝��v9�}�,�=�rq�֣�|����G�KZ�ht�M(�r|�_�	������6�js���ݫ�е�Q���w�A<<����]4�Y�&��:����_�[��o<��Q5�tĴT���.��b]ώR��n���z��t��`1�r�sU0��3����8@��eX��k�J0���˜ױ��.n3�x����\�O㼯�����g{{N9��*4Cې�u0�+���<�OC�t��i�r���l@�w��2KW��wXEt���K�]�|,�c��[�� � %uN�I�й��N�\�IktW ��������#b��,�4�|�^ւ�g^��m.��.�4-���E��qgi���H]ބ�W{70+wup��g��f���[����*��c�����.�37�Tթr���6�pj�T̴�5[Y
�&�Uj���[�;]���A`�;W[؂�zp����i3e��ڜ�V���Js���qk��E�g��8R�U}O�C@��A�jj��
��N�Ke;.']S�v�[���T��`9�K^=w�O��We�kX��a�&��-e�J�^�z�u��W��c��2����N?r>�7��X�Y�����.|��z�X���iL��S�b����ح�=ټ��u4��*�[��7���P��y�rԱ��P"���.�h�.�����^J�	Z+sF4v2l@f�&HhMe�z�:��:�u�2vS��faY�q�
����s<��7ޘ6[Z��Nʾ�Ԕ�w��K������D�_L
e�C�EE�"2Р9ۣK�'
�9�9Dʂ��ȳ�N&�9�	0���UQ�\�Y҉3���Ap��w/s2eU��*+u��O%u�%�+���{)�J�q���´�S�nNy�R�6DA���W�T"��N��]�TrG72��r��(*�������B�PE�'p�)����QP(e0�#&�v�t��
eU�^�*쫗:DUE�^�r�RJ*��"�	"�q���.Qr<�U�£�n�N��9�(�$�*��0� �9vh.��*��Q9h��s�i���o��56 ֈ� �Z��Ӫ:��n6���6��v�uҭ���'�&�n-Z�W�w{P��?���7���� Lw��oT���E�nⳫ�s�����E��c�>P��{��!��#�z���1P��{�0φ[z�g8~�+�8LV��>���:��;�x|��鑣��F�Vm%�~�g��:=�{j2�<��.��C�� ߚ�Ɲ_��x�O�ƶp��W�^{�`�=R�x�Z:�����
 pfa@� 3�@��0+��紝Q�ϣ}0��E��b��1�O�i��@�˺�z��i�y-�P~��ˁQr�U�v��?k���Ƈ��&y��V�*I���zO����	��^����1�,8hV|:�c�]G��Y�S8cp_yM{���9�)8�2 C��PeΆ �8^��S�H���H� k=���F\�>G@�:�P,�yD�l�yJ��+j<υl�,�\�*��z{/+o�jw}*!)��W����uՕ؉��$r#F�\��p�q[�gc��뻓�MW^sX{��z��S�z��o�I�9`����s\�����6D�_JB���+9�k�P\g���9����z���P
�fa]�u|�)����P��j�[F�`}'�A�b��O������HDyO� hX������c6�](ՙQð�˨L�K���3�|i�¨a�$=���D���r���Px_�8&��Mǋ&�8��q��'��>50$5����o-��b^���a$ǡ�O
�sY86�|+����`ju������d뜛����a����ai8ҨV���>7o�E_���Ҏ����*����=�X��ly�NpG;*�S0�yR���/���g�G]�w���*����D��jax�q��r�(a"��׸�������ٞ�U���?�Lvo���U<0c�X�)^(�r�}��ևn}p	�T	��}�o��U2*�3��g��c�\�4/y?܅�k��q<7�����PtO*�d+�n�t�]��+�����-��O�N`a����Ä�T�u�&c�Kh��J���C1�y[�n)��g f�y�ݫ��ټ�:��<Z{n�H*��Y����F���ø@�|T��f=�N�c��E���B��5<���u
޵����痗�2����mT�'�b��l�Y$o�9�u�������L���xġP`�Yu_��`�C���+9� �s>��t��l�D��"��PU��}~�!� .�O@��i5�)z=_���Ǭ�ᑹ4���;�,��TOԽ�.UG+��1�N�/�}˗`����$plŅGU	�Zꇻ���x��H��*�ʿs�G��NO������M�W(���aAת��O���s����>�]W��{�G_���l�����6,W���g&~�\x^^vON���{R������M
�|!�D��A��{1�h���7�)h����P~��^1_ye0.Øs�C��Dب}'���]q�Z�R��Q�3�e�Qx�����畠j��xXK_�Ŋ�>�vǐ�A�᧮������B8t=�6Y���[��,-8IS��*���<ZN��^�)��rz���k� ���66�X���֋�bb�:b����4r�M���m��ﮪE�⛌=����ˍ�D���Z:͉NpL��h�ч����v���`o�&��UB��C�ɖb��}�t��c�����Q���M���ꌟ�P���ݿ��
=�Z,^Lǰ�u�^�z��{����A{���1ӹU��QT(��uP�@ȳ�5g���8�ޣ����#�)�W��^M�33�UQ�dwM��2�fB=ꇢ*���^Jg}�����I~�f�躆7�x�us���u�&����! �r/�=π��kr�	�j,���L*���8�UuD[�*.e3gsɽ���~O:'�M�+�� ���V� ;Ƽa�d�4Jd��o=T����f�+�Z"��F�'�+�0��/�,jR������>��^W��;��_Tg+?rC��h�׬{5�^��_L���9���̉�]<'��"���`[m[W�rJ`�����r��^��mJR����4V����u�� /^��i8������\�VM���M榹���2D�a�/O��ʟ#��|�ɯ����V��;x�z<��{���G��V¨���Ϗ���&�|+�9�7ǱMy���.����'f� ϶���Ҧ.���>��2"az|=����(���8k�����m*�W���<ɨ�@��G�2L\
��
��v��f��^"���eF��������Lr�'��ߍ�#�K�,�3wf���-�ݺ"ſN��C�4zc�5�f���^���>)��*��g{W��F5�&*6��명7:�N��"�GG��:�"缽�\�{��Gd����1�1u	��]�T���L�;����.��~����;�:�VO?��pj�ޏg��R�W���5��z�_z�V�{�`U��&w�򨟭K)��ᚦ���HJS��D-v������g��:5OGL���rӳ]�Ֆ��e�+�4�D��*�K��gEN�\]@B����R.�ƭh�v�	��.�l�]<��5Z�����Ek�]k��V�iY���^K��o��K�P��Hp��3��W�g?B������@bCB���U�qs�f��E��gٞ|�[�5'B'����DW�PeΆ �8^�����q�ng�z=LǏJ&�O��0��5���%@A���>~~�[����'��_9!���T�?
�Q*�aU�|�Ef<1�8�w���"�#�<,WP��rY�z@^�1��Ϩ �G�xwUܪw���B�s{R��1칍�U9uƽR�B�>5�>œ
��G	�ԫӾ�^�r6��޾��J�Ċ��(x��\{�`�|n��̭S[+�����O]I1]s ��VN��+��OG�u ��?LñT��"�C��C�E�W���/���b�Q�
f����7��[J��\\{ۢ"��ֱv���k:�+,��n<�:}WDz_�ɇ\�9���;Z�SC#�᧝٦GL}e]��Wπ�kv��2����2�sa�I��}�xڼ�S�Uwu�]v��+���ڔ��� Jռ����GW�� L3�١����KEG�T�&w*PPE`���x��,]�hsT}x/_T��s��#}8,Rs��
��1��G�W^f�h
�\<���C�sLv�XC�G��1+%��X$sk�\���|v��(�&+��NV�-yV�Ti����_���C��,o�K�/L�L��� vz*�Ӗ�}<6�͈��I�]��)ƍ��7��0�H�<�UH�����o��g�U}����Pt��,g�G.��ʡtxġP`�Y3���1nV)�
�Wy��X���=^�&�
�����U��1�r�yE4n	�d+9Z/�w��#�;S5�0�,la�j�� �zaE/z�
��F�狫qw,��dX��(���*ʐak��H���yx)����4�>��e�v���;86%����4Q�s.��vVm��S�T۹�p�Y������̹�5��E�iY+I���r�:�Z:��C�m�;?0�?��Z�z�Gk�**�UY�Tz�yULMmA�C�U߽��<�ULM���O�����(��)M��b�gO��ʇ��tw��?.�\1�P<Y���|#π����ƍ�+�ڎfh�z�m�Nmk��w'G�Nd�=�чG�o*�Q��K
���PL*3[��V�֮���F�v�g��چ7������ڎ�"~JpW�Q�3}*�ug��k�VH�~�UG�.g��0��L?�g�X�GZ�2����@��u���c0��sc����_z���2�U����"�X\w�M-�³����2?D�v�͏��)�ܤ�7g����u\g>��c	�ld�v
�ە�O|���
��������eߌr�G|v@޺�tR g�{�3��v�a�������6#߹`uq~uX��~��#R�T����&d!��s&S��1��T�gp�W��L��B�\���M�$�C5�R����/�r4']�&l�P:���i嫟]�!A8�J��nT�7��͕��e�Q���;��	ܸ;{y�i��~è�]Sc6<,/\�b�-�[N��Fa\şg��X33u���	�2�N��X��y�*���8ߕCnX��;5ל��Nyґ;�����,{�.T�bT�V�
'��s�T�&Hj�����d�>��|��_{�j��p�4K�`#<�� D��m�+|2�4���VڴcܤyMğ@��Z�zL|�|ja�¨sS�D�6tXZ�Ei�Uwx�r�M��EB���z�	�(�
�#א��8�"�s�>�>Q�6��L�f���C�,���!x�t{����7|tx<��^Ÿᣂ����'�P����E� �l����q��7)�X�f8?��e����C(j0��ƹ�P�e���ns~�>��̨�~�"��l�D�h��L-r�2=���\��@q�b��jr������vx�%YTQ�6�霬Ioh�cz�D���0$t��*���:����2���K����$�v�`޴�v�.rqr��x���km�Y����c���j�z�ǘ��4ޟ��u��'	�ۛ�adEβ������-�D���k�'���Q����B�7U�_j�Ip�1���v��*?k��}�u����m��UFL����&3��eGCޝ1��2���W���6�w��=��z�ߡ��\�H�;c��s	_V�c2P���M3�}�'7ͤ��|&���H"Z���~��M.�M�?�Nⱝ����q|q��f��vI�8hVX깎�W������������B)I�'�2����'�7<�PeΆ �8�wT��������K���@Ώ:�_Y� �(����c]1����\���F@�u$0�G�v|\�y�p��P*]h�3
��총�=3>Ի��<�ᨌ>+�&&1�g� /q������g�i�T��#�9W7 ��nݦO囔��
F E���r�D�H9��_p/�n���sY�]�ӟ]v�䊮�)����'f�`��⯍q;t��?v��`\o��s,�L�$��T��]}��;"����t��B.����/��a�ި:�'${b����4�ِ�Qj�M�Ys`)�L��m�8���$��.�7�N �q�@7�QYgc�p��]^�]bsv�#o�>'{hj�uq=��iج�h����:l%uq�͹+e�CJq=x�F6w���u;O=8���(ےF�ɷ}hrd{YZk8���v��p����u%�"�ƪ��PRo$�=�3��@�2��{��v����|h�B�V ��Z�U�*��TU��Ü�q26��k9=圷E�n��.� XĒ�ͳ�u
�;Ȁ��6�ºv��`���^���F2Y;t~P�L]n����h��섀�uo�롕n�H/�����;�ᰳ5A:�wg9\x�4��4R������=͇k,k����X��u��s3�f�p�R�5�#��E,/���(*ÁJL���w6;�Z(�1)*{����N�JN�51�\<.�z�M�D�s�:�:zlf�����g(E���ێ4��n�_|h���s�%H�ǛI�a{7gtS����+���hBl���^����fq����I!��Z�̾����%�A���=N"6��v+n��^����ziY�s�{�G��)#b(/t�]��hm^�w,��D��hh��wi
�=-��3]�Q�hloudCa�oh+�V@����и��X�k+7,�M���`�ƾ���f�{Z;:��Mw&�ώ7Eu���L�L�D�[ԶŶΨ�����´��8L�޶�ά�6c�v��A��Nݙ�Q킬j�;���5�k���q�������3�[��5�b��y���c�-�GKDf��j-�K��I#O��`��w����$���8��zg,i79�o
��g�*_;J�-Q������?f*X���ѥ��^�BpmLS���$��[C����8�fNdZ��HsRD\�x�vT���r���A9.y;��.���q�51u�p�	J�'R<���\��������z㇆�y��DP �]RJ��ێ.�{��i��";����0�S�9�\����x����Kr����֘�t�+Ш���@���;��t��d�t\��\r�p�
��̉�
m:��S
��]ps�	ܼ���)<��B�a#��ٺ��y*�Q;�]�b�H�=,p���e0�s�8JH�ҩ�D{2''!��)*�Vu�t�2��֚^xxV�fV��YʫwOTg�u\��KZw]=���)�G�XE�,�uB"�p�kO:r=(�^x�����s4q7w�0�1DMwp�L��OW-3�HA HQ��/�Ҥ��ux���R����tT��_:���o�{K��ٚG��c��١��rޜv������g��+��^5P�j=R�%U>1�~;Ϊ&��\-��f�9��ܬ�~��7>pl���Pd�a@O���XH(eg�=���i���\B�$��x
19��j�
���OGN���{�V��.�`{?���V��a1�M�&�xi�|��\Ǯ�ev^o{ `M{j=��@	�|=P��T)��%bc8ݒ�a3�C�4��7w͵��#�3�o�>�"���<^S��3���UgE�
r��o�/����Ł5���
3��:#�7��#�����1�����k��ՓˈQu|�?%@?]RjC��o.��ʦEYf#a�)��:�����	�[V�"F�H���Ӧ��{<6�.P�Q�3]7�~��x��B=��U�f�uꎴ�1)8,ߪ�O���y�=|Kk$e1"iw�
¤kM�b��OT��i����3m�]��de^C��ru҆��նU��}8+�F��8�f����:]�"�́)I����܎�e�Ltj@�Q|��U_8�C�(`��՞	�u�:r��(�Ǝ��o�j������Zx�F��攽`f��r�,�u��*��
�Ԟ�<�v���%�cBF� Vkō�(�ı� �zc�tg	[s��iU�� zz��B��Q#|W�TaVj	�Z�{����ĉκ�^�n����<I��S[6:�0r:bɘ��T:�Z9�������*c�Q(2|�=11�%������ ~����+���2�!�ܘ�Y���yS�@q��S���̱�	���������W�僜���=���1޹��<ρ�>�����xҋ��O^y{VϠ��]mB��uB����j<7����ٱcg����t�6�F��\<����dŢG�S0��s�x\4�Ϸ�Ǽ]��D�Ա�]{��خ+�
Qy�Vo�ķ4.@�"��3-G�f��y��[��y!��<�����p��e�K1O�25b���y<n�1bZ���,�;@2�*�n�7՘�ΕU��U��jY�c�ea�t��}uP�/�p�cng��A��;�y;#����y[~�cH�cɍǔ"F�ɞ�{Ƣ�E�ɘ��jU �_��}ܰ4;[4<��Qc�7*����_�;.*��T�@���®�8qv�?r����i����pQ�b�Q�;�
f�=�~'�gV�����ıns[��ǧ2�ǼU�Z������x1r�14�G�Ү��� �Y �}FD�r��>��P�amFD3��&�'G��}�K����q�= �8�(�f��?nU#ꪋ�8��v���y5g��� m}�Q1^�x�� 1|@Q'^��)f\V�md���W�G�=��1Kz������z@�^�I��S�7�[�t|��	�뗼�: ��
��1:Ǫ+ޑ�����@Q>g��1��r��w~p
�eT�\�w�IEm�4.�8�l�LjD�����{�E���:w�u�H"j\3���>��0p��o�����z��7���w�6�}��]�6��}2�	ܯ�
X��|�pס��f��^�.��c���dG����B�/���==��OrI�����������7/��� t�c|m��`2�
�����V`�����-'9�� W���rb�&:����,��p9zo��������Ռ�9#��{ڰz�Ꮉ=.����ƹ֙�������{yDר,��d���^>[ʰv&6��0����q�;��
=����y�p��,��i���K�)����*�"��x����|�J�Toau�=�/���rَ�(Tx�t�C��;��/ʅ>C�\��7@4f.���O#a���ao*�E��S&=��Wdoy�p~��Y�v��M���Rdx�P(�.���5f:uV
��:TneۊGoq���蹹�Ǚ^� 6@L��Tȟ��t
�5s�kī칏��n1�wWS��0�}X��@�OKjfG�a�ʢ�ڋ��U����\ #��~�S�c�~��	��p��p��	�Őr���=��l�έR8��w#
p����L��r�>�G��:X^=u,2S1�Ȉ���.t1d�v�	�qt◻w&��w�:�>�I/LI��5��u6�<��@�}�.kѮm>�J�G�υ�1\@b�=4����X�T ׼jS��s�ph�����>\+П�:��DL"��B�B�1>�Q���x�H��t��{t���;˩�\B�G\ǯ��=P���1L�g���O��ےjr=��绎7æ%�I�*���2̓���Pd��P��G��w��ng>]M 9�<},�s�
�"M*�
F�7��\���I����s�^��չ�X��`z=*����,/7^�쮊ʵ]� K&ab���4��~�IZ����� o�:��]L?.�
�����Tp�%{�Q��{5�,.�׃�����z"*�ΕMPu�ʹ}��b���49\U3b=��b7zˠ��!�n!�=B#+f;���r&v��:����冺�B���9:��1x�֭��o%�i�P��\���ƻ�[�s�.c�S�:����q��L:�C=k�r��8��h� +}P��Qs,w�i����[����s�N^���w��U��z@�Fc;��&)T
s��#ñ�ugT^Ob�������3C�V��e�j@H�Rۊ�s�f<�k�#���ؼ�{��b=s���u�:��y!���.���ڑ OƉ��K��oy��C��6:�g��#�x*��AU���f�@;��7�2�;�+�z+n� ~4<=�b�B���
��c�>�y;�MȺ��t��>$�=��/��V|�ɤ@c�|e�9v�]O ���9>p�fo����!��O����Y�BaTk���K�:������)�'�0���M�����"l�Y�&-Ǔ��]�o��&J��(�
�3���'ߤ��\~��f��2�M��(ذ���~�����.��31����Gv��q��j��&�M���;��8��Ҥ`N�[�HtCc[4���}H55A�PT䡳sK�Y��+脵:�������^:խ�����%*����T9��׌����*�"�*��5�}�{�.�Ѣ��3���@#>1}� �y�>����W;�m����~4W�ãN��n1�
���j<6��1�(P܎�#�Y������G����ݔFx�q�(z�UC�sӸ\4���TO�hH0*�ϓ�Y.t6?L@~��m7^Us�ׯ�k���;v{��rnO�3��k��8�~�Y�������h��J�MO�Ǒb���Μ�׫��Qٱ����X|{�
�>���_��:��7^��튟[�>>� XH�,����'zp_/rb�Σ����v�/�(����{6�p�dX��ꊋ-^L.��3�����b���d],���f�<��o�Ѩ� k��Q�'҅|Oi�1��-�r���.��G]�=&}�Żu�+�p9�0���x�e:�.]�u�vQ�|;i��M��m_:Y�g��=y!ܱ��me��]8N�z]�
��4u��2����qQ0vQ����lE����X�R3�-�������R�T�V������+�F{��@�.I۟����L��ju^�x��T4l�1�G��ai�nQ��Xڰ�{��OޗF9��z$��� z�μL)>G`��ˈꇸ��=�ʽ^�ϐ#�X6t>2Ll{��ǀ�l���`��|Db5B�o/-����?eX���*'T�3WQ�?z�L\B�>,x�x���ޝ~f�t���ۋ���2;�X�Ɏ����Y��k� ��Tg��)*�Ȼ�(��Ѿkk7ܷ�=��C�H��,ҟLu_�Ǉ���t���r<9+8�"�e,+���A��B/JF������p�p;�C+�5����L^��-��"���yҏ5�`<�x_��Ur���&��J�j��<.���{<���ﴴ}q�#C�v�jX�Wx��tOX�_�z���?Y�m�7���:��p��//�T�߈��7N��VD��gED��8�&��1}B���!��ڼi���,��Ƴ���qQ,�K7�VC=cv�N}�*H�y��ѽL��d/\�}����~b����ɍy1�gJV,���v:�w�)>��ν�zO�A:m�G@��4����1�5�G*��Աw
b�瑎ϧ��j}�yj��\�V����Hjn	�0�CYܪ���ƖT�i
�[���O�;�R��>��Cz�EX . $s�2$�@��ab{#ޏ%�`̜��	]�q^�uⰟE3Qu,T9��_�O�!ۘ�s������O�m"�Xl��&�b���x 7c�����(-!���L �ד�t��=]u�X�)�e�q%��Lm{��C]dz���t1U�_ziQØP�����f��z�Ǽz-�3��{�;��d~�@4,Tu�+��qXL�]Bf�R�$���/�j'�t���>`��l�*��'�I��8(^A�~�\i��Ps,G�n�}/zZ�	\E]����Ք�f��j�왛���d4�n��� �}��G�*h7�`�\�|���wl����P���ܚ�@v������ �j���jR;���Rnu��ئ=�'����s�$���<��67nP�>�f�=k�^5�3��>a���צ|��W����u	���:O
��g�Y����pi�=���}q�ޖ C��͎���&pF|�
��^'��S�7}���s�UC�YS�d�;|9t�z�0hIL)�N���2{=���z#�B>8��[�`Ģ����1��b��I���G��槷�,.���K��,��袀�U��6�s���q�����{wʽ�R6,e�e�gc�@H� -���N�c��^+�9�Ǔ�9%��}��|�U��,u�S�玨!Q����ж�L.�z���g�r��y���٫���V��G���Eg��PC9��(�W� �8����ɓ|B���Ɩ:�pJ�Va3b,����)�?��?�L?��S�12���_��6����UQ=�).J�*&��zAwW�J0͉g�$��y��R�+�" �*�g�I�\
�*Ēa"""��P5�^\!9u�[iDneg)������F�%2���m+���MA��n�O���kp�8,4���0�/|I/:�h_-Q��V,P5fY��5�%Q�L�\�׷���QQ?`��
����bV�3W���N�/��>	�fO�]1�h~GR����������)����D�=�#@Kr
z2_����%#$��j@��V�3�І�w�`<wub1�+�G��/4� ~���DTH�ќr����,  L*��(QDl�"�E@D&+�V(M��!f�����o,�j�MG������������h��5I��\R����%r6oW�fW��>������0����_�UDTKz�s�(���4�$��.���B�d�A����k K�>�s׏q~�SȈ�n[��n�C٥5�Կ�����m;�DTM�Ā�1���1��k�c�g֒gt�!�#� *�f(�UQ=���}�$���A�,g@�q0,	�����uTTK�͔��!��4#l�|LGH�PD�č�y�.��S34��b`���X3J!{���e2����@��J�(��4W�ᐻӀ����9��`H��؇OC��?f�=ư>�3x}��(	��xk�����@P��%����!=����R�~�f_��$TED�:�����b<Rd�{�Hb��"�'� ���F2h��e�Y��|�M������/d����$�w�R (��s�H{G��ՐZ�@ȇ��o��x�h`�Wqz�,*"�s�p+`˘S��i<�]1 ��$�fN��٩�Huɇ��KE��K��`HQQ?��6��7����Î��*'�rM�p���ol��Y�������Z=ԥ��� ���"�խ[��.�p�!7�7�