BZh91AY&SYӽ&� ��ߔPy����߰����  `[^�  z(@_n�����$UO��:��n�|�tv�F���qUs6�J���TRh0;�A@ H�.��   p2LPh�vb@b�@@ �E� 
dI �0h��`Z��w'�(c� @VP     >�)	R��HǪ���c@	��& ��0j���*IHh&�@ @  �	��I��4i�4�� hz"J��1  0F&�  B�" AM��i���i�h2��@HDҩTd 0 &�`<��>K�D/��@AP��U<}�( ����Cm����F6�7?�ԁQp@���A����a�X������	vJ���?<H��2���a��v��"�"x|-I4�(��A
J"�##-�F�j��DpB�I��~jIe
����w�i�>����|O���y���%���c�z2�q�=Ƿrm��l�,2J�666�cz�淮����f���3X!�޳Y�q�np�GX��1������ꊆѱ�ؠ�8-l�)�t�:S�<�[�<��v��b�-_G"��F���Cb#��b1�������c��p[����E)��h��'���i�*Cb���c�X<o��~SX��<�mi���B#F؎�D����-/��It9�y�["i		��c�(�6�clZ�b��z�:�X?,-_�i�����&�Kb�,V��c���Z��s_��sw_u�\1Ũ�#�/\xs��� �g���\��Y�iu��j4s�!!�����7�m��s�u��O}NX��o�=<\�Ln�7�mz��jcŌ�1�rKF�Ճ4�5����p[N��Z��qb�8c��y~�M��'�d������o}�{�����xs��3X?x�%0)��q����]��!p�d�����x?�pZ:F�cO-���Z��i�Zx6�Zb軈V�/	
Ŕ&&qyjx�A1h�����]^k���%�.�	�&D�pHo�o�ݢ&�T��#�)Dm4���c��Z�����c�G�F��n�G;�5MT7�?GVG0�`��O��E?#��9�+	���n��Fu�S�Ŏ��m�f��t��g��O#�x?.�Ga%��p$��Ā�	<8�hg�mK{o����|��F(G��[�,j����=^�sʱ�Ksʣh�ءN�lG[��+ky�pPtsU����Zq�����8Z�^x��y����y�y�y����q	�k�Ʊ�q���u��d�,k���;K���zKԖ��/#�þ7��/464�h�9\#�eT�T��D�y%�Ix��K|�/%:$���1��#��p���3�9�r�/)U ���ph���~��>h��=-4:XO� ���ȩ�?���Ӥ�_�͝���ad���i������3H�8H��JEX,��*�S,�?��ܕ�����w�ҽ�B�^��~��~:�=�>����w���b��h�{'�2\�	�q��0L���}.E��f`��n�6���o���I�#����o������#�3������Й$�Ujx��t�fS`��d!�t��dz>J��~�焯Ma=�V<�%��F�
���9Pq��N�h�n�Á�� '�e�-���6I������5ң(�h�o:��M���Z��:�00H�,9�5e�/f�?H��>"�l�����(���Hᥡ�ru�?�??5��	�S�OϚ�gJ$�n�9ޜ��t���p+=r��x9w�:Y��4
R�yW=��S��v� � �C�ko���́
h �f�g�S4Xv3�ҫ���� �6�`=�B�ε����T�И���B�-ó]�z�|�^Z�Rmı�D'���Ú�JcB��c/�ź5��g���}�: w�=�(�Vx2Y��m�6���c��Yh�g<�C.w�y�N̜l��*�(D�YT޷ܵ�<���h5l����81���n���(�Z�V�n�HH��)ev�&e6�7��'6\ݷp�Ξ{y	�
Q����T���pҚ�M]�sJR��F@���Ud�ۘI&M�b6+(�R�i�<�<4W`�{! �F��# �3��.˴�3J���I.˵6�4�k�C�4�%����x8 A�Ѫ���B����$���{.:��p��q�D%p�_�ۙ�[K�m��H���wq��YE��\�e��u��ں5u@�,�����5��y9˧ c���v.����t�W٪2l�%�C�?�9� �,l���!�E0�8�L&CJۺ�`�e\P�����5���b���Я��0d�ܘ;��Q��S@ �.���p��|���scj1f�X�4��f���l��o�>�ÿ��'��x�������x=�{��4$|�������^�o�
� c9���PL@�>,M(L�>h1x[AP(��YY�����n!�jҊ��������N��q�kl8AZATec��KB�+-�6�eh`�$=mQp4-N1v�``��l�Oͻ�X�pL��������wh�Fɩ�--v��sti�,28�+MT+	/����S��Lm���{0�0�Q\�FCyV͚�vM��e�pb�:Z�}7O�M�s�ԅ�#d�f�dN�{�&�M�+E��^����7�͵�țryݢ�h��s�`�*��F�1�SV�֚ %���O�ք�'�	J���0"l�4�ǌ����iM
�}
ǑbEZy��B�MخW()6~D��@pS��ݶ�܉���r��u	2#����A쀌Q��m�F�π����m� �*k�8�zm�#��{�C"�'W�Vvk�JK�*��1x��{��|#��~�<�� ��� � < fbs��SU��Rs���� �� ��� �:  ���5���[�i�4�ƚi��iw�`  �*�� `P  ��k����c�D�a`���m�|��� h� �(���  z��������bBp�in&�$S��U$�J�#@  � *��  h�  @��I$�I8��|�>$�KQ��� �  UT     vw�}�ikl�	x�|܄��B�k�M�S�'ēM$��N݁  �`  
��`  A��Al�}�80AڪIB���w�@  �`v��� ` qr�$�$\�\�ISI6�0�Pmd�z����"���0���ۏ/6�`Ndd<a�� �0�+�/�|�HB�	P����5�B�H]T�.�R/*^U����+B�!R�-B���Z�Q�*B�!�b
��������7.��Z4}+]K�r�婌Q@��H�ץ|�"z�@�do�����buv9bL\yQr�Q:��Xk�B ��AZ�r'#�r$+ &JBQLrȨ1�c[6z�UN(�Z���y���uS�ע��[�UScp�2�E�ʭ��6;l�Y��ީ@R�+U�I��cD�GI�P�S�Ջ
HDL��m������ỻ��>��kZִ�&��kZҊkZֵ� ��kZ҂�Zֵ� !�kZִ"����A�7���!mP��Q�I�I�]Ȃ!�a�����ȱ��m�z�E�g�܆qn����{u%4����|Q��zCE�"�u���8��!I��P���Og3�eeY3Ï+��hnlD����J6NӃ"�3H�2�E=W=S��ՠ�1Ng�<�q ��Qґ�qQ��zF����z4h�F��o��.�˳�>�4�rD���h�L���Q���#�.���t ��0��e��eģk^5V�q�n*aV68�l�sH-8���PS��V�פuDZH�a��U���u(^%�,��F�im ����4i��j+kIl�4w�GoIۇL�F��*���ܥ|GS6m[_-��ƚѣf͔h,�>�`��M��K��6E�H7}m��F�_qo�M�E�Y�f�6s�|�N����13���"���ny�D�m1Y���g�gϗ��.��p���7���;fYF����}z��k[My7u�����sU���ʹ�dF[���*1�Xw=W����LX�J�J��j��Ѧ��I�99Y�OX<:����tnra�n�: �0� 
6�bg��RQ�i:���ZDF�'"��9$�l���h�p����x=�gF�c�>�O!�D�	���0�,�3�8T0�2h�Ǎ��G����xz�c<Y(�xp�'�7=O�<?��`��0}0�8CfC�n<,�Sp��B��S�������w�}�:��Y#PǦ�Y~�A�j��:����E�+��ZG9��9@���X��k��>�mc�m��>ۻ���{�� �6l���&�%���9!p�d����y]��zHN�F�"ɝ�ٔ�C�c	#zc�C�lp��LK�=*�iiƓ���k����,����n�^��N���Ǧ]k{2ʼ@�Tr�6�j��+-@֙�^�Rd�dឹ1��V/>h��yIя(��h�R�L\(k�RQ��SW�����F�[$_ �19)ka]���c�X�k�5�[8�I�yq0�嗶O>���5:Ix	���Cr#��%��8��QlS,`������ۍ�`&`ڹ��	sBxb��ܭ�3b�F;0�78v� hI�|���N	<<��N��'xdv���vC�ѹ��f,ɨq��9:v̧��R�GL�A�<3�-�|a������n��<�����n�#�p��d��!�%Nux��32�3ø��$_�E}�B1�,bV��T��⧂5�Um�!�X9'�<$m4~�8~>!��F�[��,����Ӊ��4ia�.c��.K��U{m[�p�2xך�x`���!F�6�� t�j/	��:HE�Ha����Z�HfΖC�f�>�o!�33 ������d�NEr5e�T=q�5� �e�338#h�#dM0D�2*፳X�oIZ�"�"�P��ub�,"\CI^�p�h>�י�[F��a������I3��؆Q�>4U���Ih�4��@���#�v�I��'���4I�)��1͍��V�Y��8t��r��N
��y�M	'NT�(""�Z��!�ы��<jI�յ�$��.x!%�<�b��[U����:M���bi0��ҡ���k��I퍑�͞(�h�͛!#6�T6�]И�vB((x�%�.��b�]���]]Fݺ�r�s�kA|�J�:�}�D]5�����$��h:���xc6F3�D����h�-�O����#0��3���Qf�̏D�	���v<�D����g���������=��0xh�>�N�&�!��Q�F����aD���A_g=��h�Ok^���ޛ`�́
h�e��Gmy� s/��&��md-W��[�Z��.�C�^QQH��n�)z�n�؁a�7v�
�xoli���xԵ�뀦��m��C�6�n7��7MoFM\�e�X5�ƚ{�9���� �rJ4�緜hӓv�vG	�Im��lCU/mȗ&���j��Ze�T+[�X[�Ԯ�FH���S�mD���� ���~���Z���j�e�}m���ܤm�H�۔�A
��x|
@�L��(�lV�vIYpu�,���a�F�m��:�̫�B �x�CAɁ��d��Ӹi�5(:�ͱ���L�������"#2p�63��K�k�'T:�A�q.#�X�?���R�f�~މR�a4��@��PU�6P\���p��p�A��Ջ�Z�R��������/y�̉0=�r=�f%�i��J���lj/�gF���4>��nҰ_"��:B��F��om�5�m�2Ý�:u��
[�b�4"��"[<�y-yiL,h�GI��8QF�D���$�hmGdCr����j���,���:X�հ��(*�Pw��	�>4���P^#��"Z@Q���]}$oi�P��[m��F�H;�l�(���;���o*m��%D@D���Po�4}���A��pÊ�b�iPoG{^vnU^���*�mSM�w����>0U����4�W�4b��(�e(��G6���eZ=���n����}�����&3*QTQG�Kk�Vt��H����m��|��Du�*&@��,�D4O����agɍe�<��D[P(����o��yh#<qe"��c:cZ�-?+�X,6b�])�W�����å�i}Sh���R�nեZf�ź�"�wxnGM�ouX��������9'A0�li�k�"�E����:��]K1PYȃ)U�_|7�e
��m�"}�m���A�qt�0�-]]Z�D֥��F��l�A����jQ#!U
�&�Q�6݅덍R!�]M��3KJ��ڠ��.o�⳩(7�R���}�.�h�1��@�-���6R�ѳƾ4A��f��x�
����4<:K1G�x9&aVa,�`�f���4K�S�8=�&����Ş0�0��a�߇�	��a:p�!��4K�&O{,z�z~zo�w��fe�]G�����ŭ�Qͬ~u��zq V��	�nx�m�)�ۖ�m��m6�m��m������d!���CA���_�������7�16)����p��ta��Si��h�<pz���l��t�h�T@Ѳ��:l��!��W!`��|���͝���5t[ڭ�`ģ�¼RK	0�a��sa��Y�a�p �ֆ4aA�}��ڳ>(f��s�HIS���.�I���X�ʹD쑍͸Ȣ~%��RHB8ޱ��ҹ���.�3O�_�����|^0{��Qa����h��|�ѳ��a��N�d��aE4��E*[6CG�͖3��V�q��h�a�1�VyZ��M���f�t����40٥�_6�d0�gxi��0Tb(4Y��!,���h4}ߟ�+�*]P�F�����g�ѥa:ߤd`2���Y�lv�έ!n�mh��Ƹ"�,��h
D+KSӥ+6Cf�,f�Gw`�~Xu|���~u$��U���T��(kZ)Kg�JFͳ��\���3H�Tx},�E�]!�(�h4g�W\ײ�U|R�n�&�,!AX�bqF�v�-�����6<`bkhٳԸbp��}���l�`=�l��_.���هh�K[>^ �bȏ!���$��4|�����e�����pw|����fE�2zFqml�Dyiq��g�͙h���S���l�Ҵ1��l#H���������Q�Q�(�D�H����l� |����������EA�CMq//͟!��H�H����d�l��F�A�������T�1�ԫpaj�s�)p0e �63����/Z����J��J�겊6�oO8�h��6��>j�SD��w�_�_�g�M|=�W���>�D��K0&Ha0xQ�Y�Z,¡F���f��q�'����y�(��<<�~<Oǉ�������F�E��������eht'Rk�yK_��ʋl'i�@k�K���9\�Z�s�	KQ��Q;o~p�/{���fn� !�����8U�@�n`��X$��yw�zy.='�x.@a��-��A�&���}�n�W����S�jJRf��\.� G�Yz�r��y�Th\Ύ�&�Da��d��-�9�� S����m��m��m�-�ܦ�m��m�۟�1 �0e��8��Y�n�ұX��Ml��mM���;T�=B�h�eNM�ݛŉ�G�G�e�h��Imb��,>�j�Í�Jϗ£�����k���a��I4T��CT�14Y���8t��8Ϗc.Mࢅ3�)6p�4m�,�N�F^��G����s��:z�ã>I��ӡ8M�ߔz�(�p4w�7M�G˫������|�{1h���vpx�ǚ&-Gt}G(⥬�\]]-. ��$B�(�l4��8��s�ccح8Y�G �a���-�����13��P�#vw�p�q4EH�v_��J��ֺ/��||B�4����J�UET0�ob�2!Э\<X�C]�Jq���3\<���A^��>���!I��-"h��J�TFί�+08���;)u(�3f��
Z:��8tCE7Pn�D^F�o�G��F�6�4qC��ڣe"�4���7*���Y/,�P�Q��K�δCᶍ��>(�t4gv7�b9^�����9
�"0Ҥ����D�ŖErf���&>4�T���ʌ!�ty05K��$��G�)q.��j!�ɉ�j]��� `FC�Z<p�:����GP��l�ͪ��x-R�GDmm,Κ_+*QW���Gˈ��Fw���jaY��2T#1H�!0l)�]H[r�+��nٻb�KK0uY8��ZnkE�x�94�V���ucG�HnՇ Z����G=��ͼn��8f#]X�^�zL�uiR4��ǌ�T�c��:Q5�od�#gxx��KԸ���O�ZB�v�&�H(�M�f5T&�Uz�X�iL��h�Bwf�Z2"(�Q&�{m��.ꜻ��ը�z(�Y�.��n�m���5�M�c�m���������a�a�����	��`�0�27��a-`�M`�|8M���l�<>����<|O���?'�Ӥ��l~���"���a,����]�7�,�v~b<�zq����n��/Y�������`8+���?Ze��m��m��m��m�m��n���{��ٲ���;b,�c"��+J�|���
E#�s��
���~?M �|l���ZV�Vh<�U�"�,Ũt�񢍆�E����&�Yj�R\Z:��Gڳ���k��lm}t��X�Z�:l�%�,P F��ZᡃC
y&W�x�t��d��cq���)\�Ɏa%*e������q<[]A1�oV&�laZF鑚FQ�Z[,�<3~Fȗ�*>>qp�m��*�6iyY�����Y	�lgg�2�m6�[Y��x��TU-F�鯞�h�N��Zg�F�E�L�Y�>궨�a67N컷v�Yφ6�I�a�及�:?�8|Xl,�ܕ��I5Ob5L|Vh��QË�Rf���6��P���}r�z���ѳ��h�}Bvp��o�KI�D��{�6t�M����CAf}�=`��>.�"Y5�I��r����l��"�_WKE����h�kmыiR��g��9��ϕ�h�Ta��Y��Q�dϣy�����Lѣk��qm�q�D")�lp���d�@��<X�؁����3�<�1;���Qu����ښ|0��d��t�6��>hѿhx���u*��k�՜6��0�|{�a�&���ߗ��ph�Z)L���im4B�d3���w��)ܹH�Ո��pdVB*�8���#ڵ�8Xh-uﰧO�H�*���u���(�h��(Q�[��ѣݗR���9�|�2�hg���T�&uZ8�e#�8<C�R�������ܔ����E�V�:�+g���.���iZ��\���:�����lf��հ����y"�C��%Ç��K$�n�1�l|L(��&2�0�6K�L!0�a���VdoC�a�3	f��0v>����8W�����O�����<V�I�pp���C0t<8YT�������9�� ��W�ʢ(�e��3����i;Y�.6Eߏ�G��b�[`��AHJB矵BqӨ�_��6�Pdr��GkL���sH�wז
���B�-��e�m��A�Mj�"��Dswv= �Æ�����$~��N��ۍ�W���k���酎*�%�`�2F�M���i��$��r�,C����f�v�6$��=*�\�ؔ�/� ��I�R ��{}��m��m��e��m��-��m��BQ � ���!�q��e)V�I�	M���)!\�0t����n8ISD:��I#b"3Ɠ�k�ǆŠ�<�U���PΑl�H�ܙeT$�r���:�����:h�l,���"��[zTgN*���y��q{�ϣw��ݎƛ��R�-�00�R���g��&����R">4h��h,�}rm������b�3���DT�}��f���Ӷ��<��^e�H�ຎ����qh�ņ�ǡ�z��M��1�:h�z8/zF9T6��7]1G�^I}�l-��+1Z6�ZZ�<o���s	�|�{�Gm���Wd��q�;�1�߉(�oX����s�����kk��ϐ��~��>¥Q�m�Քukgn�ut�7r�.��5�0<//|kC��|k^ZKqm�q��#H��[-Z�F��C8uuo0�Hッ-�΍���{�<f�ьd�h�|h>
7�2���D�����[䲝:Ig瓟/�H8�Y�E�
,EZ���vI#r6�$�,��x�y`��④�3���k,���a><|||rg7Ou���� �F�
H.V7�ǵDkQ�n�U>�J7NFhy`Z�׼�E�f������*͑t�4q�ˢ:�l��ar���E�� ���h��x����Q��k��RA�vXәQ8�S���/�I��xb�Es�x��p�ɟ*��F��Y��9��G#Hэ>��a,�ᢨpڍ���>����Æ���
��fǃfL0�p�މ�ل�d0vQ0f&��q����t�}<W��x~����ό'ǉӤ��t~��∼Q��ü9Oސ��L����w�%&�<�ј+��3F����&5��yO�[m��m��k��m��m����m��(�03�>��p���j..'m�����|p��p��`��q\4QI��]�Э���P�Xp(�Y'�8�DO(�7���ٵ�����F��� ڈ���gM#"���R8���G�͖
=�7�}P��]�"���U5#`Q�eq�6�p$v�-h�	Z��\:�-�-E&Q�+hj��ķL��v�I@�m��#�"���g�������c��#���\4�A��M^�G�ZGQ��Ŋ֍#\^-(�p�����b�Þ��uR(�E�G<Xl(�쁳�l{-/Nъ�P�h���o��Z1b<t�;�#�6��f��!������6l6>�s:i�P�u�Q��hi&�x� ����L�Y�sK(�<|�L�:���Of#AҼF��qm�K�!�"g~_��&�)`:��p��\(
	������wnI_P22I�<E�E��%��<���f��ݣ��՟&�- �_M"�'Ө�J�h�:
6k���lѭ�`�1�#�Qkg�[ޒ����Z"1��b�G��u"���p�2!�����m�Q���>E/qF�n�E/����Y���uPn�;���F���uH��c}�>F��Q�RD4l���5{ Q#�N4i�M�����J�+����a#y���Z3�l��5���"�PbcK�{ ��Z:�Ňux�ū5v]$Z#3�c���'��	�+��S�!�=S0��a,�1�C�	�ɃVae�c�d��a0|������3ǉ��x<��x��ߩ�x�}�/�,�/йu^�S��ڤ�^<j�MbG+'n��ډN;Ѱ��ϒG�u#2_dfX!�'K���D����vϬ2`˓yJiE�vc�p�����ywkjJ�[�z�(j��u��p\|j��Ʃ�^NcF�f��ɹ)ϑ2GC��MR�gl�&�L�k�wu�������6�4�x�E�"�Y��7-`�;_�\U�#5��t���G�v��qc���pu�(KPD�,h�:7���zhS4X�����c�<A�i�)G�w���m��m��m��m��mV�-�������g�Q����KjI#�uuTF�n�m��覴��HXە8��*��r��vOW��ƻ�Ũ�m���M�iqe���3���S�(s�Y�:g|�+��8�u�=.-�p�[^Le66�8����F
s�<�D��R�`�]�}#�k��:��hh8|Y�������f#Hgɲ������D}�E��<,Vj�`mmD��k(���!��ݮ���%�É���(b���"�o�����o���_/b<�e=�R�lX ����0��L��rv�VF�[Diƚ#��,J�ZKRcjZ!YDH@ȗ�x��g�̫�,�;=�z�m>m���83�G_d1���
��p���y�H�M�9!�/��h���l|G0��#�⺸'UQL<�o:x��*�ӾvBG�DY��04oZ��|r*LŴux�1{T�dsjы�tG�χ���O��|���Z(����(�Y�}(r���ȋ>\��{M^�"\M=�WW�-#k</3���l,��~Ќ"������q�؜�g��e�����j�1S�lAP֨˦�]BG%c�2g�[��'iyMi�C���t�凳���:t�N�w�Op��6ӝ.-!��Y�����N�7QIL%�m�b��6Z�!��]����l}\^ �|���Gܐ��wd-ݩ!K��5���>1bi�K˂_��|B�j�y4$$+B�B��H]T�.�R/*^(ѣ�G�ύ�a��a�tٳGƌ2��Ca�f�]ѭU|�ˮ3�a��h�=�g{���tf�r<mL�d�w��k
�ǀG��*��W��j��W�R���Yo3ǝ^i-�')�����Cϻ��m��g��U�,�=ZI���/V(�&�q��p;i~��n{���c�Wg�j[d�����1e�˪W�/7�1�<�~y5oex/S���y���eۭ��{+خv�.^��A��4�H�N���ٗ'(Ps���ӡ���>�=�x�O{����m��m��m��m��m��m��(��ƍ�F�VbT�Z�v>e+�vW�/�K��u|�1mmQ���>F_CE�(�Xw�4aЮ��Sy$UYE�t��p��E\���i<�����/Z-Tx��p,�3[�E#OuLnA���|QSk݊�l���AGboNsw+[�`�xLA�1��"�<847��êͯ}D�ڣ�:4٤Kg0�^��R�/
����p��g����,�;�hh�Ҏ�V�།����=�a�Ӫ�ꪘ,�/�Y奲�!�Zm�my24Qг��T�c^>QR�]Gɯ#T|8��u�=�*��%���H��CTG�͵g��:M?F6�i��4��3�l��K�d��}G|��h��8�uo�GJ9k�>E#Zh�GW�MuER��t��9삊�+U:��KS����{6��:�kT�X��R�cnF�&l�Cϋ�1��Kj9㤥�`u�R:�sC�¥B�F��<���4t�
6pn�q�(̳�^4�Ү�����}�8��x�kX�mE����QGϾ���mǕ4����ݚ �4�_h�2ۓ�v|��ZW���^��D^^V�7KȣgMp,�VǢU8bIǎlDi�n&�f��s���W0m��������-&s����r���{~`~���(���UT ��}���gڿ�����+�:���� l B�Lд��/��Q�&ͷ)@�-P�!HRu�`b��A�
�!��JA+�!��!,�HA!��0JA8��J� A �+��V		B	X$X!`� ��@�@�P��V	`� � � � `� � � �`� �	X $H0��H 	! ��B!`��F��v	R	$%% ��V	Y2�BX!�	 �`��B q10����	��H2�:7"L��


) �|� d�$�!`fv��ـ� � &C! �	�$�h6�vHdrH $�`b
�`� �� $��("� ���$�
jjJ�("H�� �f  	�f ������&�d���"`	�a��X	!	!�"	" 	 $�bH*��c�%�H"	!b	!�f�!��&	�`b`&�&���HBHd�� $�"&"	!��	�`(
`��	�&2����JHh`���B`&"	�&HRa�d�a	!����(HF@��`d	i�`$ H X%`��FBYJI%� �BH$ ����!`��F	R	!$H$`� �)��FI��e���'&������H��2d(�S���u��y�	�m<���ޤ�/�4��FWϺ�S-����bY*��a<C7�3�E��:�[Eh�\3�q�p#����EaX�vz ��s�Đ	�+<�ռ�0_�ZG�� �S"���D��[����~�s������	��VLķ��ȟ��)�;O�Ɛ��h������P/����0��z*9C��"{�g������fO�9_��$�����ռ��'<맓P|�S�������6^x�6&h?w������ܘ�����.�ll�`(������e���JQS� ��8��0��צj6�o��~���?��z���O��F� �r�� A�� � $!����m�
�B�Z�?R��~����y!�Ǡ�r�0A�}�'�)?��~�����$�
�;�kzV.4���JK�(�����ȍ)V �#��e͊�L�̻B!�l��,/Z@�֭��u����`-�H��h`�
`n�	3߿#YUD�&�7L�p�a E��>�(
��Y_�����3m����}�{t��vz��B�p��>�(����Ϸp�l��P�6�����9G�0g��q�lL#�&8'ÔND�xu��������t�&НKП�=( ���~���߃����?P>?��O�0&�E���p� �:<�R���t���"���sd-��r/:u�&��$q�5�������'��a����X%-��kB@$��dg�����8�w"Ð=��} ��W�ʼ�p�DGǏ�w7	܊�766�?K�}0|]�F�qP�V T�-�"pL��J	�P���@P�?!{��>��n�'Ȟ���>�`����}��?G����yS��S��Fk�p�㶼��ӡO_�T������ٷ�cܺ!Ox~������Ш��jn��߽�b�|��щ�ΥCG�h�#Hs�Ca"��/�����)���4`