BZh91AY&SYP;.9��߀`q���b� ����bJ��           x7�
	 Q@H �2V�I@� 
  (
�P�@P@UE �(   
 � {`@�-��՘RJ5�%J�� 	&C@ֵ����M� R�4ձ��mL���kOB*Z�;mj�+�l)I\�A���TU�v]�SMh�Mp  �E RZ�
I)-��5�l�����T l�Y
4� :*�(
  ��RH(4��� ˵�@j�F�  �w  uv �`���� �
�� 
$ �PHu�*ER�zR� ��핥n^o5��GN�麺���lw���^���^�\{��ʻ`S�M���t��ښ��םz%���v���� �#=�8=�^�@���z�f��͆F�j�J��R�<���{S��M�/<w�%�g]yx�)Z�x��C�T�u��T(KѤ���JP��Z�7�ojV̠/p����c���m��w���GM[�|��҉}�}�z4(-� P@wҢ� �>쐭�������}��nr��>�JҕT3|��B�������P�_N���OT����+}��ѡ�=����i�����!����jt��}{}�T픑�TР�֢��j���|�E  á;����n-��[����t�ך���c�h2�;7wv�+�٥��A\���;j8��5ۭի��J��*��Z�T�Tt�r���;+%[ʠ�	B��$�*���JP ;����	�u9�u��lj��ӃM����]ִhk�]����[
�ܞ��Ƕm��^��
4��9��UM4�;��ۻ��%�� {ڙW�:H���*�Ɗ46�Ϥ�@����47uN�Eh\�}��+Kڽ�Tu����U�]v�
*I��������i�̕��v�s��(7a�
i�hh�[b|�R� 7��T�o�����:F:(�����@��-ºT��j��ظ���5]����� :9��:�Pu�ӣC!��Y��ҥ  w�� q�wr�x=����"�Ek�ۀt4v��t�p�z�g�( R�Դ���n�ت��SclMfED��Wϥ)  ��һMW�۰�u��p�V�n�
�gu\n�W6�@;f��v��˂���u��u1�����  �T��QH S eJUF` hi�� j`bR���      S�2UR���      �))*�jd�� �`F�0��%$b�M 44  h� D�Q�RJbbOH�"a�2hi�b~C����ψ��W��Y+�n�1~Z� !��N発��o�������e^�저*��i@EOԨ *�����(A U���O���w�ڧ�X�RI$�-
 
���EO� 
/����_����'�1-�lK6���-�lb[ؖ����m�l[b[�6��F�m�l`�ؖŶ�0m�lK`�ؖĶ�-�[ؖĶ%�-�lK`[��b[Lb[ؖ����Ķ&�6���-�l`[al�%1-�lKb[���%�-�b[ؖĶ%�-�l`[#�Ķ%�-�lKb[��Ķ%�m�l`[�Ķ%��bS�6Ķ%�m�lKb[c�Ķ%�m�lKb[��Ķ�m�lb[�������-�lb[ؖĶ4��6���Ķ%�-�lKf�Ħ%�-�l`[L-�Lm��Kb[ؖ���-�lK����-�l`[��0-�lK`��Ķ%�-�lKt�[��Ŷ%�-�lcl2����-�lK`[����clK`i�l`[���%�-�cؖĶ�-�lclb[�4����-�lKb[�����`[���Ķ�-�l)���&�Ķ1����-�l`[�b[�Ķ%�-��m�lK`[db[ؖ��%�m��`lm��T� 6�ؠ�0�6�ؠ� `�l@m��T�*F"�[`�lm��A�6�F���T-���T�
6�؀�`�lm��F��l@m��*[`lPm���A� 6�R��1P�"6�؈� b�lE-���Q�
��bl-���A���Rؠ�blU�-�0�
��R؀�Kb#lm���m��`lm��A�
��؀�b��Dm���6�� �K`l m���T�6�R� �`l m���A�6�M0؊SKblm��T�6�ؠ�`����
6�F��`�lEm��@�`�[[b+lm�-��#����"��"�T� ��R0Kb�l `+lEm���Q���V؀� �آ�[blm�-��"60Q�(��F�
�Kb#lDm���@�(F ����`l@m����6�#[b+lm�-�A� ���
��K`(�V؈� �6�M1� 1� m�L@`+lTm�-�U��� �:`�[Z`l@-�lb[��%�m�l`� �`�����%�-�lKb[4��Ķ%�-�lK`[ؚm��%�-�lK`[���%�-�1�%�4Ķ�m�lm�l`�d`[�Ķ�-�lb[6�[�Ķ%�-�lb[��`F%�-�l`[�Ķ%��-�lb[�Ŷ-��1�l)��-��%�m�lKb[��`[L`�ؖĶ�m��[���%�-�l`�ؖ�1�6���-�lK`�����6��%�m�lb[�b��6���-�l`�)��m���m�lK`[ؖ�Lm�Lb[�6���-�l�b[�Ķ�-�lKb[�hm��4��%�-�lKe0-�l-��)�l`[����-�l�b[�[����Tw�A��ܯ�	ػX��.���L�	���VnA	I�M�K-�/�n��a^�HT��+�M�Tk���\M�{���I�X�1�Lz�^JZj�� A�(YV)T���tm���;Gܻ�Rb�Z5�q�7��7p���W1�+�t�@���L-$#�lL)�Y�q���E�ABC��ݯ�b�@�����r]I�/e#z�!t�LͧG!U�B�Qj��:Mf��7�JE�qIM	�T���%�n��[��5Va���W��� ��k¦0��j�T�WꖃJ�DX��ieU��e%�� �{"�I�D��j�㴅��"��d��b�ZY"ø�,���b��m܆�C0�9lN�+=�c�j�j��ZU�{�Q�]\ݻ����ܤC��ț���w�R2)�q�l�7Jڂ���H�؍��`r�0��j�-�nU3N�6�:Y���k2�0�-�sVU���cIl�������m!��/�eU�+
�h��	�T���T[
1N2�ŧ�&�9h��e��Z6��5��R{���p���wwN��a[�chTmc�4��r+6�k��(V7xQɚ�^mь`�մ�����alB�m^mX�8R�/28������Ȏ�{������TK��ӣ�f[�FL7Q/'n�cm[�skV=��KJ�Z�@��N�W����yy��m�V���װ��5�^?[�w.y�/7A�e��/^��y����o�f���7v�jwݮ�.��W`�j�������;Me���-�\%aѱo���)�z�%���u%��Sʺ��vd��L�{Z�X��!�(a��EW�+$b`h�8���a��lkŪ��L��o��	A�:r�n�p-.�a$�����[����Z�W#aT�m�<<��z/�ӁЬYB˦�c�+e*)���5�z������n����i�����,2p9�CD<�t����p\(�`���Q���WamN-�7L.�T�I��"�0,9U5V��X]��G0i�Q����N ][5�3m<wh�u��zĵ��͚�m��zƨ.�Fe8��T6��F�]㬧�*�tm��\��:ӻ�wV�/1m�xn�!eX�hR�S�nk�яwJ;��f��6D�uW)IXI���KLHse�(�m�8�`�r�7i�6̕Vp�P��p�Ԉ�M=��ʩ�a+���R���lN�v�LAU�^��V�5p�+d��CMe����'2�!��Ҹ��O$��j¼:�=U�i�ä-��U�Μg6m優b�ѱ��7��iU^�k���Y�d�w�B���X����mGQV�*R��+,6�JћT�#]Fª��X�:p��W�c)5cq�f�x�d�eś����ݙ�	ǒ��ֆw#r�i�$�Z���]۵��c-V㠠O=6�7�m��M����)I%f��*�J�Ԥ4�pE.�&���Z��on2�o���Bb�U�K��a�Gz�/c��+ja���)�f��6Ϛ9EQ{���t/ja��kb8�(���R�cN& ���Q�"�+��ܽ4�sn�il��;a��:u
y���{.BĨ��f�n��f�����P�V��+(�7�֭i�Z��5�gR���ea���3(���|�2��%�vJHR�b#�:�1V<WA����$�,�s+�v�{)�gV�3*�F���F�Q�I�n���x�U������q�m�{�\C=RkQ�)JB�̴�0<ƭ�����"�f*m��VN�w�9��F�0@�ڕ1%�ۥj���Q0�#G*�Q�Z�A����r�m�5#Whbؘ&ᙹz��=�ʶ4m����$��1?7r��-�r7�k44솮�	{r*���M*��_�h���ʃ3��TLS��V����H����n�Z0��g.F)�%T<8Sa5�-�A&N1���Y��)aݻ]���:3oB'H�E�WdXDe%�ӛ�����pQ��$��e�PQ��rS�US�e���#���
��\���:��f�ڢ��0�M��p8C�{�/+MA��۫J�m�RɹKv�U����śV��t�[L�MU-�/H���\��)3���)�ݻ�yQͥj���*���廴#X7n��-f��J�Wg3R�������܄����	�')YoK��VUդ�Ui5(��k(e�1SMmf�)v�i
}M���74m�1�V"kEM��0N5f2�L�8��B�5ɋk
6�~�t&����t�d�j����y�͋�FV�B`�S%�3P!/NB���,#h��̢b5xu�YyJ��yAߓ����Jޒv�u7�Hݨ�LN��pVe�r���Y�i�x��}[w��3�E,���Q��V��QX���Y[$�U����o4�{Z\�����[�zl����s(!��n<q�zq@���zCt�՗WOk�c	�����T3"m���6�Q��醋j�f�)PJ�m!�%VM�/b�=�/SӮ�Gv��qи���7e=�qI���iX� �d�s6��UyL`xҲ*�,�6��+R����7�]�d�YAl�X^2/.�-/. �����-�֋�hb1�J����*�ň珦�9��ڽj���aܫ�F�ּ2L�C5n��j*>S��0�^��h���7b�2h��a,����=��Y�T�)d�,s���P�T�k�7�E�5�R3.��e�^�W`�Fe����9���ɴ�P~6r�r��4�,��˳��D�Ѝ�H�eb�B�,	d:R�Բ�Ե0@�QxuKF]\���M'jeU�B�JA-H�J�h�o1��˕�ȱ��{��� ��,D�=5iU3S6�g�]-���,���a7�y��Y�w&�[�u�����PFWV��Kr�c�d9��c3o)����i���J�t�LV)
�e���R`e!2]�6�fDNӱAٚ�&	{�a�UAF���h���si��!�˸3"��o���qʕ�S�T�	d�t����eǭ�����ا��2����Z��49-wE^hyzi��F�����ڃDwrG��ޕ��7j[{�P��Yx#�f5w�jk*��̨��m�˻�1�깭������V�[-�TΝ�۴.��z"�wr�*�3hk��
B�Y�X���K���V�HQ5VN�VY�k9��[7RwXu�(`snO`��>�-�����j֫���Go"�s%^e�4(r��C3��4lµ͵)���^<I��V��1,�4�Q�(�Z���A�IL��Q-���9�)I1�Y���[��f�u�֪bc�~�Uy�V���;%շ{��R���/.Q�:�5�f�����8n�5M+.eC-��E�x��c�ъi$�Cjfc���V��oV�.d0l�vw)d�� �[b�X V<�A��Rov\�����sҴ+�u�7r�	��ݡ�x�S"�8�A�wZ��`[E7ۖsF�R��iͭQ��[Ÿ1P�DmVP�.�n��oU����s}����wr���a�茕��+�*�m�ӄf�kJȯqf/.��+y&hÐe)E2��c�Ґ��Lͬwm��,��Sp�.��(;�݄�j�Pc4c�1@TD�����f���y��[��Q�ő6���/O��1�RN<Բ�aB��;C����vjg��c�n���P�x�&��(]�H��*��Ψܵ������+�3vmڥ�P9��C�z�b�$UVm,5����Z�*��I�I����2�J�Q�V:�Z�y��ڬ�����
���-!T�Bl=������%�.��/A��RwM�{�]��i�"	�V�-���6En�zM16��Z.��~��������Ut2���e
@ѵ�����4��6�/յu�tyY�C����0ڃM=TjZ"��d�;ٚh;f�0��R&���â������˲*Ӹ��nЩ�1�X�Ц^A����/0�iҍf*��9�PM��`�]�;�m�V�5�2a��S�Z�ӧD���jɢM��m���;�V[�p�!�F�5��	�2�mʻ^.d��-4	̬3���%b�õO
�w#T�K:�@�b�E�ݺ����#��Hj��9I�����n���d��t�!� �G)�i8�2�QkK�&�����st�*�#v��̋#�whY��)3f��k�UOn�����l�w�n;����2��ڒ��RT�܃�Z��{u��+������+&k�[��9�0�Jon���m�d��wY�0�b�C��P�T�w6����юr��MUi60-[�+SJ�;�.P�J��ù�
I��L��Z����GfS�ZE�f�d���x�7��ycciH1E��[�Z�yDVi��ܷ�y63�!���.����QYR�&f�5c��:�R궽{[Z�d�Q��ň�⠱f��қE,�
�7E���x�9xf�Wi-��͆:�hԪ�7ۓ`V��rK(�RA(�tff%�-	��xJ�Y�1-pHE���;�W2f�sUh��^ظ�ѩ�a�m���.�L��(���[FM��V�K)M�IҽyOYD��K��t�*=��V����*��^��2n[�JbF�]E-�2��1�ٕ*]���k���V���ܻ�bXo�,</n4M�p�U������۴�5��"���^�E^�7��"%�(��eY�͉J4c9��{�lLT�B�U�6���L���M컸��bKj褭��5c�h�Snm ����2&�k�JX����mM�"�%T���s!��L�v�
V	��	�#q�[W0V��5XJ�R��T��V�R�5z�S��<ي��r���Km�l�o�۱�ciKC6�N�S:cJ�M�Eon����!Ga-��>�T8-N��,����ؽj��'/cB����V%��`�DI5�0�Kj+�J�Gɪ�E�]�4�-nݒʽ�]j�%�.�5�ʍ�cR��M%8�Zq98�)�&�Z�t��JSnY���Uh���K��7���`����oׁ3��
9�k6ӭ�4�VCp�u�a��k�+L��0��Ui
y���͙��ʙZ�j�Gum^�����N��m�U��F:���U5�F?H��V+���,���6q�ŇVS��i�:���.-+QS4^<�AFX����C�cn��q)�Ա3tfePW(��1m���8�;KopZ2N軴���v�x�e�$3��T+�U��	�0�*i��]���T�6�:GQ�=S�e������Zk;Tw����AY�J�ք��1������jc!<n��
�L-Ƕ�e��m��u���Z�^M��������l�v�%nX��a�K4�e[��fo��Yb&��ƅ�7r�+��F�8ů*��8D�����:�4�׷(ͦ�i�Xd�H�0�팻�s�D��Pi�F�U�Ŷ��
yg"�أzwsj%"��܂	ĲR�J���7T�ĸݻ:�����Mm�h�U�v��;�%
�Vpf�	эcD[�7j�I�q��-]g�˖u��Li�h���DSЭ�r�^�f�J
P���g����`;�j�B�S�1k����ztS۹u(;1no�J�P(6H�a,�歹��*�A���.�1�ka�kNR׫/*�RP�S�r�,Qc&�i�*��Sh��8X3+7��	э�.a��0^��W��D;�U���͖�����ؽZ�Zr�g)�T�i*Yԝ[&=Nl[��e#�]�6v��i���KZ�fmnY�ѹR��]��W���BF$�#��&���р��%�͘��ce�j3UT�%�����UcɆe-��1Jڤ������N��d���T�e���髮�l��SƫM�s.��J7�ۛ+7���.��v�i�bE2�-]K�U2�Gxd5)�I�H�M��i<����no�B*��i�V���{o��$(4���WQ�����B��ŴT:ۭDTUZ�f���eU%��U�$vU��Wg!�h'yx����Ǵ��b������E��U=�����QjD:6�"����F�j�oe.㰸ze.J�i.1UX�'K-e,rb�V��L��;J�r:�Ӵ�JE�ֶR�u`��1SxYrE�0�M��K�%���Z�Xs5�DiRoej�qTKrHv��ՕT�>甆��[SC����Z�t�Ԙ/�őv�U<�E�g]e�h;�4�V1f���5v�kiM�l&뒋u*W��^�C�@e�2ďC�qdJ�y�h�y,�Ń8V���^�6�����,���S��A�W��.Ujx���A��ܳ-���Sa��fwM'*.�Ga#�-D�I*Y�T2}u*�r]����I�V�&q�หjk^���m�P�wX7��N+�aո����U,�.�邩R'b����+YkyN��"O��Gl��J�]��
�U-чV�d �.�e&��Yj*[&UD>ɝ[�D��]�2���%�!�]��%��s!�\���;-(�As(�ծ�ݝco6�8�M�ɥ��(���]y�-��j@��'�m]+=x�9ɂmlO��`�L�$֭C�5̊��`�T#āi;U�㻧�ڢ0�ͽJ�)KTwcȰ��F&s!�A18�[j�,Uj��R�]̢��u�Uc�e�Ԧrb�!�'J�NR,��U��U��w
\�j�6�jqp4�T�Uj�(�ޱM˺�v�*�R�bԵ(�\���m���k�輍����U�˞�Oe(䧋ԛ��M���V������v.��-k[����8b4������^��%�ywWJԊj�Pp���,kkj�l��S1bLip��-R8�V�;�6�2�ͼ����xrcʨ�jȺ����P�u]�ڭF�yWjt�+m&�IbX%�5JI*�`�	#�V}����:��.|�U�g}������R�Zv���|��%����E��fIK[�f^-�O.�U�Wi$�
�F�U�b6�'&�cSV暆U�kta�d�/�'9�{J�@m�J��+o7�:�)rM'tzMX��\�l�αqڻJ�J��I������J.�y��JRZ�U����;�o=�f�i��o�.�������zT/_�����_�O�q��Zw�--J�w���n�ˬr�n�!�$��6海�8f�x7�_\����*Z�9v�a}t��\2���e�VԄISJ�
��B�>k�
4m:�)�`T��Ic�A�c+��5jS&1�e���S�o s9L���oڪuNǷ�J�9Au�vZ��I�;*����+�J���[������
�ʃ2���$1�\,��ŗ��Yr�QR���5�q�sJ�����^uRU�`�)��^� �Xm�r�/5S��\�P&I�MK�gLXT�֪i�Q����PCM.�}��	�*��UJ���W�Nm��^�BB)�ץ�]8�Q�����X���n�!T�͙��o-��7sLO�PF��f��j�L��,��tvo*áe���v�.su�4�]���EQX������"�b�w0�W�15,��1a��A�������q���A�H��X*�û%.��UVRy���,C��ۑ�H�n�5N������Ic4���5�6]�6k(&���N�mhԦ�)<�FnI�fĬ�S�xS���fª�\���d��rW1ʍ���U��m�Ŕ� ��hA�t�6�BR�m�����8c�=�)�ˋ%+�z�y9jQ\o��ө&LOE#تUga�n�Y�-R���2���,J�#UWD��Y�j��X�`��^�QB%'�=K�J�$-�N�ù$�C+j����U[,��m�dj! ċ[���b�W?��N�*勪���0g�N�9��aŨTCTT��F�ϲ��sR��D܎����u��%W]�.��U���q�k��0���]X�lZ���Z^�@�Z@�P��/�goVYWS��I�kkv��_�Zq��0�3�l�.<Wc��6��\��o��љ2�A�T��P.r�����gSڌ%sT�ՃwE༦]J�f!xc�r)�/�e�2,���+���o����\�-�4�KJ���̖��m��Y�Q�C7e�ĵ&�j����n��YYkA�u|m�V�� ��A�\k�i�
��T��c³^�u��� �y#m�o�uL܉��.]�=֮����7���w"���ee8Ywx�v�5t�\��wz��]A&ʹʛ��P���Ͷ���i��1;�Ws��(�\X2�:�[}xW���%)�.S���j��Dk&��2op�՗���:�t�)\'Kɛ�&!�V��r."�3%m�om5 �*eʗF�n*Xy��8�Kój�vͬ
�˖(n�� �L���9;�$���֑dUI��V̍ �v�}i��7[_8g֙�,5����Z�جUV�?\%�oU��t��>+�0��U��#Mr5$�
Y{�#'4d]#����<_#���N�jb��������l�}�cfX��έy�x�y���k�N��C6���^ȇ�6�,����ܳU��)o���}s[1d��>�zFl.;n�0N~�V�r������ڝ\�n��+�%�7��9�ytJq#%-�&���m8ʷ7��8�噗Y[��5f�ڻ��\z�m+3x�cǭ^b�F���r�����c�*�E�ܤ�j^aU'�f:s.�Ȃ�]a��������)Z��aRF���G��K;Jf,B�����l��.�ُ;l!@��L���yS)̘^�BusӁpGvW-�z��*���M�,�T�H����5"�s9l�������i�����[f�Z`'f�''R˰dt�;�S21ٽ�=P�2��Ed�4+uf�NI���[wU�.B���)S=���N$�Y�U�*�s�,[D՞��V_N�#����L��w�K�A0�ae�QV�rL,���oW4�n
�w���*�bxZ�=o�Z�;����Q��i��7��i�Eo��p�+X��+I�نiƃtiakKM�-���,�1x�dl}Cn��H�
M�6�*<����TLUT@�M,��3Zr�b���b�Fl�-h�KۥRm-�**�G��+����f���.������)��[QX�=��Ի�5�Xwl&5�Ve��6��T�V��"H�]e�q\��ř־b�t��1�+��s�ʚ�;�n�6*w�r�U�[EQ[�-o7/_(�J�v��NI���vp�L��՚��Ns7�a�{kρˡ6�u�2S�	�{�ǋ/�ɱf��u�p(jνgGG[f�	�)�78n�0���o�����L��b_R1��(>5��\Z���z�NU��<���c�P)��m����mL��!X���ʼŏu���T�v�Ek��=}]ND��7[=M�ҩѓ��L�xz��GD>�кٻInU.t�K�;e�zfki9�+M�x>�w�rU׏W<�6�a]�X�V/��s �Hr�d�98�L'��i�WC�\YrfPڨ�OCjq��(�zBp�f�i��b3W���ǩ���>����Ub�f���������GjȤY�e�X�K��\��kV3�����Y�$m��x��uR]����Z��X���,�y����1r�(�ҷ!HL][�Tb�X]64�#r�k/(m*9�Pָ�pۊX���
���]�J�u9vK�w�fv5���έ-��3�D�h}�a�:��>�ҽ�DX꛲�ڋȮ����ہI5���}[.*=W[K�e>W�bH��L,�V��E�D�����ژ��f�'�M,�~�D�)"U��X�޴Vیt�+*,No5[�1V�V7+�T����Tj�N=o�K�B��/ws��nSlt�8�J�VKⴌ=vO;�k5���l�+���q���m%ͳ��G��ۊ۷��Vj�l�e����Sl��y�+_T������1�*�)Vw��v�8��6�qX:zS����X�fe٩�1d�ږ{e1�5(���;�hܬ}]F�z�0c��f-�m̻�����z����/}0όDK$#���yU7�-y&�ok�Z�3i�GC�-[�}���P]�Ԫ۳�ݒm��LV�����hmQC6�j��N��V�nֽ͓l�W���t���T�jJ-��p�]��v������;Xm�%DP��wM�݋�1m^�k�(�n����h�T�f���L�LiЖ!�"!��`�V���-%2��A¯i�U��� J�e�D=0ҕ���p��ɱI߭R���6P��[�ՙc�U��wj���jn�](ɑ�(�N*t�Y�f��M:u%��ɗ�m�IW�.�G-FR�B�d�̇��ȇ6#��:�%�Xˢ���WW�hw�^�N�Ƹ�	��i�!,�2쪬���f���16ni�kP���Xp�|Zs2�NRY�j�ب�/���4���|BW6C�n���9�{qP�crHZ)���4��X5�J�]h#$a��u�s{��d�R���-k��j�X�e�v%Tê����61�t\	vf�1D��[Ý�:F"�c�/X�i'�6�&��0&ch�Q��]4�>$Zm�bf�u^7�/���7Ļ��#(ͧV՛��9���Oi=�J�o|y��N�����w��Y@���/Ams�r%�=U�b����Rɸl��#��X,�g�7s$�d6�F�=�V�r�9d�m�����D�	S	���jS�h�r�#3����c4���J�!ͰH��[��H��\�Lm&��I������P�X5�R���ʍ�f�0��h�9�[�Pڸ��B�F��F/o[�U���l�k2�p&�C��}�.ʹ����.��wƺCG�8NJ�]e�h�(+�0�M�bbK�Z�+�v�@J&�qK�=B�5�Yj.�.�J����!��$l��#d]���y��|BO�jء,V`��Wi2�MU����o�R=�.�C���4{z2Aػ-
�6�=�u0��M0�>��4���'��ۧT��u[���.ܻĮ�;z�R�R�#,���*���B���2.f�4d=�%�uL2p�Ո�w��h�MO��Wn��Gs�Fw�	��2�]��8���/-'�.��wn.h��t���Sg����Z���f��`]�ҵ�j��y ��7����l����.�8R��of� ��#و�{z�'q�d�P��/%V>Rf..��T�l�I��a��I�lU�46�`�j��a���hj�Ȫ��N�[-�;���L�V��l�e��DfK�\* az�S��{;7(���:�����j�]��|r$7N��Z��;����
��B+!Z���$/ZB;܏��Z�8�ѻե��ꂚx��S�v[�nic�*hYy���X����[�*�Rh��A�fB:��t��1ɪ=�\�s��o��F��ڴ���h�yo0�f|n�� Ψ�폣gm�{����%{I�rX��o�N�un�ez)�ҕa�ݵ�'v��n�3�Kqۣ�!L�t�)v���~�X����e#ӭ蒶н��V�<v�5E��e��O���IEͬ��Qc,�2���밇%R=ӗ4m���vr�U���g-�j]�E��Z�����V�MPY<X��ou׵��N�x%c��^=p�]1ol*s6��˂-}a�E�Lf����do������"޺ǔ��e�)*Y�V놕X3S6�R�<������5����h�{G+�:j䱍���P�TrN�\eB�%�	�Y��,�J�dS�R��%ŪM*qr!MKt���f6a�EX��Q�Jݘ{u�a�F��-V���,ի��uE:�%�D�����^w(��Ǟnv@z�mݝ�n<+C��R7(��4٣����ԃ�w�Βؼ|uwu�A;��_��z�^r�]]�+h���ꚘO,����TM�ZrL�H�q��ZZ��q��N�a�����H��]5��*�R� D]�={�[�^�V�J�qM��ƣgt�sV�θJ�4w�y��R.<���W{�*�Iھ�C)���P�CX�T�[STT�u5-���=�k`�N�l���##��9u�oF� ���^z�N�v���QoTݛ:��<���-hh=C�n�7&�����5T��P�}\7U�Q�}�H}3�Ż�W]m� �c��zj�Y�-�x�#F1ү����V�V��q�:��4u3���cs�j&��n�,����۪�w5Nqr����d����t�6=�֗d6p�uAe�}a�����}{��n��ugn5�`V����w+Qy8T[Jh��V�@Ծ-l�v�L�[$ŹթZ�Γ7uУ����na�sn�y[��o,�>��$=teϬ7�m�^k���N�3ٻ��T�:���퍧[OxU���͝�r��Ӿ�M�5i���7$���:��	*�ޝ�٠R�
JL+�YV�/j�ZUc�x��[��]��
J�|�ޓ4Vdrz[Ji^���ɽp�C����U$gE�Ι�x�v69Н�L-�go�(w��E�F�j+is
��+�%���2�Ӫ��+4����hm�ǯ5[T�۱Y&e�W3%��\�Un�%�ҝv�b�Jm�]bzA�u��m>�(>�8��%�)d��M�2Vb+#'/x��,�F�F�-��Q���o�%ldЛ}Yy�b�΃�U�{m��������;5}X�b�5K�r�ٲ�X[RY��	��P���P�up�F�����F>�wJ���O_Ir���#T��j�0���U0sc.�����!�!�r�g,���e[6l=�) mQ���)43k�m�l҈�� �������'H׳o�/fSl�n�Y16����hˣ����pJ;Q�V7��{�F�pvK�+",�1QWۜ��h��T�h�ݯe�]7�_휛:�di��N�7b�M���j0�aT�n�6|SQ-��YVlDA���k4`�I�Ƹ��J�LV�nj�ћ��!����$��̫&)\�|о؉fp�H��̷w��'��i�,6nƊwi����ϝ��z跈⦯v�4$��.�:^�Nl��I��nj��r�<a�OS�H�aTVñ��5W�����Y�N��hW���(_IW��ᖊvC��cv)�iԔ�d68�s�t�6�	�Z�_LǖLU뽴|��|/V��i�f�)x��J�;Xo0�u�ѯWq˝�u���'-���RjB��H�s�N�Xڱ^R�uCc���vet�4Vm7"��K��Z�e�m��Dަ�m��]�i�e�jy�ږ�iNbN�m���ɺ���ڞ������������ �H-����BV�8�0{�G-�g��)qgV�u�Djb�.�<��w5;�*���#c�q�>����A����u¬���t��_>���#����OOZ@�E�=E�:�8qc�C#���>����I,Wz ����x",�i������ZGs�'a�ٹ�j��s7�7Hv75$�����{���2��VC!pȵwF�����=����g���K^��z�*K��O'�,���ʞו%
V�]�{W����7Q��4��gnY��v�����hI�ΟUD�,�{ކ���|!��Y����֧6�TŔC�۴�t��� �&�$	�@U[�F{����V���"G�(媽zE���&6�&���˸��F#�x{7�2'��<�4$�f����$?�TE~������QC{��������>""�?��?�}�����}�z���_w릹����Sܺŕk��U�l=���\3(�w���5�ҡ�s$�Qo7ыl6�6�7=S��E]��'v��s�2�,	i.�1��.XW�uG�V��7�=��A�1[��6�m�vVK�r'��tf�Tk����0�+����.����1;yx!�}��*��iS$e�}�q�B[����=�U\��wy��[������Y������ـ��2��b[��Sa�Nm,�:3����h��V5���:��ro4�sۥ�%�Eӛ����B�bSM�UY���w�+�u���b���)��1٤q�cn���U�Op�=�!�0�ʍ��e����R��Ld�+�Zꪅ�7����[�[J�+/S�1{�	G.�!ŉ��R
)��*��K2�V��Vg��B	�S=�YEe=E�pP�gKב�T�WEA�Oӑ�hp��'w"<p�j�G0�a9�١.[��!xŌ��*ʐ�0�ٜ3nnq���|��j�F��#�"�@I4��R�E��p����o9��{-:ŗX���S�q���w�+�_f
")[���8��ڰ�N�:Ime�
��ڋ��V��޼]�%�$d��z�uJ��9D���"�Ǽͪד��6���ˑNE�%�*\֭��+s���ӷ�^<v�8�8㏮8�q�|q�m�q��q�8��8���q��q�q�qێ8�q�nݾ�����8��8�q�}q�q�q��8�8�;qƜv�8��8�n8㎜q�q��qӎ8�>��8�8��q�q���=���Rjt����PJ���	��GޣN�Pk\ȩ���j��E�JA�k�*��4���&�sΨ6ȩ��g�����.��qݬ�+�j��p���b�F.��]��ʸ���Zĥ�G��)�����qNbK�I�]�̾�Bc7J>YXrެX�m�O�]H����h�'{���B���6�u�xD
�������	v�b�]=�Y{X�]���1�.�vs�f���Ʀ\�u�AX�wr�L˗f+Z��jT��d�4�g�WL�QW{��3�� �o�Z��!jED�X���RYng2�KԲB�6\�p<r �Q	pӲ,R�:�/%+�8ѰV&�XܷLR,]�����ui�p��#KLbrh�RP�E���m��[32��v�ܤp���U3r���LMg]>�Ϧ��b/\h*��iۅ��z�⏲ڷx�<��8�:A1��~=Q��>Yt�p�8
x�j�7�S�7cTm�CVNɋ���v�y8��ȈY\����
����=+M�T�+� �Z��-�κ�rq⏦�&m=���]H�U�R�z�+;CͦU	
{t��f�m�]�Z�f&���_'o��b��zV阰�Q�\)�t�J4g5�;�Daց�1�Z���Lh��N,7�7U^^�˞�|}|}v��88�8�8��8�8�;qƜq�q��qӎ8�>8�6�8㏎8㍸ノ8��ݻv����\q�N8�8��8ێ8㍸�8��4�8�;pq�q�\q�N8�8��8ێ8㎜|q�m��q�q�qƜq�q�n0�.0�l\�R�*J�B��%���c��e���ժ��slnl�f��=��7'�{]��V�N鼖0�wm���WYQUmVt�V��s����~Q-*g�cd���Һ����ңB�^9	C�q���4x��/Fv:��٫T�u�1i��/��-WNֵI����/]�D����RÉ��5�nn]����7)٘F1�Q��!z���=�Z�sٝ;^s�޽�M�7�n�o�\f��_M�ipF�4��m�v��a�����m�qu�"�F'�.�� ��R����o+3*�wa���н�x�ý�ȳ/D�����%e�T{�Y·S�kFV���F�����1wVܒ �o/iL0v݆w%\j;�xCY���ҋv�Y]uW~ݐ���LE�ݏS�mY�k][�*����Ǘw{��l�;oy�bguئw�e&j�8�z����E4�\�ں�*e�K�D�65��B�x^�檬ǷL��y����`��gLI[�%M�1�m�$�U�ĐgPa�5�(Q��Ws3�p��an��0���B���O-�L�{��@7I	��zQ�}�s�\�v�$數�}!�Ƭ��dN!�WoMc]��-�R|E,u�226(����ӆ�i�^�\aӲ�1��g����gU�wm)�P�n�(��;��yy����||�|q�q�q���q�q�88�8�8��8�8�;qƜq�q���N8�8�ݻ�v�ێ8�8�8��q�q�q��t�8�n8�>8�q�q�q�8�8�<q�8�8��q�q�q��t�8㏎8��6�+\�\ݞs^��9�7�:gN�	(:1�<��ܽZ �p"��e�vlܖ��ria�����5[�[tr������$�Ԇ[gp�ٲ��S�ĉC0ȑ��`J�����('��.-�s�⠨�L��'�c]<f+vm�HF\DJ��۶�<��Ԩ�x���=�h�;B(�Uv[��,�f��ӶS�&eZk�#V�]������M"M�to7G6����Q8̬���Q��=ףS�R�{��I��Û8�8-[�c5fmw]�6��X��ǗC�+h���3���f����"�$k;�.`鍆P��z��\�U��m�8��]~�s{�̌�c{�gx��4���ԱSq�����`c"^F�5b��7m��R��.�������NK<o�&�w����n�lL��F�'��:k6%\j:j��ޠ(���At]uZ���o�v��$r�z��0�'ÞI�GQ���j�V����Y�S������H��wY�`Eၷ��xG�$ヘH�)]̪ۺu��ꋬ}�����!-1YqH�lK�ݭ{��\��ya{��xWd��=�u�u꼹R������1mڗ��-K"�KuF!m[�7[����=��>�!g�v9xycU��g6�;٧c��j9�zAO�ǐه��o#l���m��ɵ�����Jk��G��������}��c�q�q�|q�t�8㏮8�N8�8�c�8�8��q�q�pq�q�v�۷m;v��qێ1�q�qノ8�8�c�8�>8�6�8��q�\q�q�q��q�q�q�q�x�q�q���N:P�~k�(����+=�!���ܴH�U4�sU�����j�0��lV�$jٲ�g3wkr�B^zby�J��j壬�/J���/�v��sn����81Qއ��"��c�xІŎ�d_IE�k�V�qW�ҵ�����]hA�7Rwk�˩b醰�H ����Л���Kr^��mY�*��T,�QӐY���5xi�;C�
���W�Zn�ᜎ��j��9ۭ�qR�k+LW�w:P ��d�9�i<b��l�K�w�Z��!�I�� �e�*)íi�.D��+�9�f�����⾃��&�{y�:��uF�`�+���n��J b��,��rͰ=�5��+C+��J��ȸj�|������j��VEs��h�人�k������l��K��*{��32a�v��m ul���؈;ZF���'��䐧Z�ڸA�6��N	z�N\�.���9X�Z����*�V�8aF���D���Mq�_4�b�;���ǹTm���S)�pOu���4v,̻��Y�8wZu�������ѱF">��r�IVj����FHd�.mD'v�[gO�b;���:�MU%�uI�.nqzs{D
�u�0�Xܘ��F%��1Q�E�$�%M2��]:�,B��>ʸM1el�����h�N����<7��T� ��-���nǽ<��4�����u�����]�Z��QQ	nda�"H��B��IU9�]�kzN�V�u�J�:�xUֽ�s�+/X��s��*
Dzφ7���]7�u��I��e�A���9q̝Sw�b�e�l}6<X��̉��޼]p����C���<��ݕ. �<�|�ڴ�v�=T�����yfge��~�oS�Q���]t/�>�7��=;Xd��:�j!���9}U@���ixثQw^��ݱ�-�4eK�Z����J�I���XLB"�h���3_	E�Ϊ��"6L��e���9�!M�0�M��W[�zK�/8Vb{��w(&JiE
H�7�rw2�"��U���М*�k
R���<*`ޡ�&㜄ʕ���M1xl&y�����Nb,&�(�c�����[baQ���Ԩ���xx�/�7N$�(^�c;�K��,���n&�6�l��WP)�oq]����K`�ܱ��Ǐ�>�#�n���7�rd+��(�3�t<�lE���hA�dQ���0�l-r��+b�&���H�]t'1���z�d�[�W)|��+������qڛSIC{8�mqܤ/r�OiTf�8i��RƔ�[)Q��%�V�#32�5k ]���h+o���b�����@��_��ڱI`Y�jB��N+�'7[�hs�2���T���Q�X��I��h��xA�)<3�uIZZ[$^���rb��æ�ѹ5����fޤ��P���mV�Jm��Yt51qN8�{	���/���[f�n�:Zǻ�&o�ك3���Wf����K̇�J�{����ƏQ�{Y�� �P���Z��6�r�Kr
ӭ�0�q��w6Z���A�`��@�V���dGͮR'�%Y��
��u5j̠a����Ӯʾ
�"(�FU5��F�	IEPɝnJТ�(a�i��.B4��av�c�����j�ʘ�-i��Ʋ��O��6�lǄȘ���m	���g�>�
��m�}s�"%�5����a�F�mҭk\xݴ%iY�:�r�����;�XVI�b�w���z���N��F��]6t����V�í[ur�E+�j�NnSo��Q
ӭ!�!V�x�yA����i�J��/�븷(e<����Iãa�E�����sr��ۉ+[p)���L�Rc]HՙIz�"�5NRHV-���v��U�!�'�3s��n�5�\�t���=}x�V�hJ:��ǚ�
�f� �,`�\�^`�*��kH��N��nȥ�UX�6s�G%9��ө���ܛ�Z@ l��.۝Nmn�۵��vY��ԫ�zY��r�̏��Px6�N�$��w���Lu���P�)�݀�$��x�f-�Wq��f�9i�-է�L�Qh��Z�&c��Ka<�t�b}��e�y�O+���Be\��;����P��ñ�JBź�AⰫݣL�]�CvL�iͺ��u�8]��G���َ?.uW\��h��D��f�\�G�Y���V�VcY���P��<Ą��ȃ�QeN���L��T�hI�r�M�ƣ	�°���u&���'3�𳈻�w��$\��Y�J�Щc�c�4Z���amvs�'g,Nd긖;-��M�۪u��S	��Z��b��5J�����)����s �oI�ͣ{:�7rukkK���d���A�#�#��v�vW�������I�8��V�_�<�5fY�x�;.e�Bs���vx;�Yyԡ�L�����[TLwƦ�;k{�r�ִ���f^��zљ#&� ��۾��Q��}y�Z��ڢF_T�M�O��p��앙�MӜl,]j�m��[λ)Rt�q�IM�
e�6���ܝg0"�CFQ�d��u�v�+���̝+������6+}%U���' k��d�l�L��V$WL:�Kն�ckx��N����,+v�4iWAk(�έ��W��\3^e�2%Ѷh�]IL	�v3^(ñ!��g`�F�P�(�ke�pm��r�y�hd;Y�V%٧Q�7��Vu�n+�0�Ŋ��R�5�������ے�b�6��ū	�E��n �C�j�Y�b�d�N�6����l�INߩN,�v���Z���xU�g�R"�J5�f(��Dd��78�jm��e��%jOW,�$�JM%�&sr#n��L趜��!؜�]���;�����׫,�R��d�U����b5n
J-��Ёt���t\<��Kt;;$�b;�Y�bN'��s�t�Ї�5����<�a'��L�b�o����]k��@��zf������GjڣNN�z ���L�ږ(�X�I���D:պ�Tf�v�MJ=�ۃV�)����_�s����g˰�Ӄ�:hU�]Av���wb��f!K���n�1S�Hr�W�)c7R��op�k�<�(Ӻ%���L��aÜ�{?X$�qp�|'�u
#wf�5U}��#e�K�v�6�ݨs�m�o{n��$`i
��V�s���+0�+8&Z�v(f�Y3!+i*�sY�6Bn����Ξz����ݢ$�5���]���|E�5��9˘�V�p�'jf����s^ۦ���B]}7�l��P�o�3CU�ޅyP���*"�/Mѫ˘��rW������.�7J��\'P�ޠ�PU��P^Y��C�����d�����+J	���A�S��ٴEKj��z�(u�!�P��"���"D��҉��1m�YN����bwpU��a��I���VEB�#�x�>��C=ԛ2�������Յ�Feuj�vg"���U�˲IۯY�ܳ5/(�y����y
�X��\N�j����|��l�Σ]%[嗄�*��Vj�����l�:ou��h��0�$h0��B��V]���1��)Y&�V�L�|�r����+�3mV�6t̝yc��i�X{k���g�֝����v��p杭�5��1�����=Ħ%p�bw@ʳ���j�3�����^=�E�bR �f,S7���8�c�Zpl��g:�&F����X�p�ZsB�2�5��f�hG�ɧ�e1gR]�������e���a��;:���!v�*������E씎[����x"��bT�=3ܧ��"j�^♦������W}'k�a�H��*���SWꬮ��p�X[5B�TKb�R�юȽ��Ġ��ZFʰ�k˱��q�XWt�5�1�/���m��/r��{���M̘�ވ�I�M��5Q�Y{NQ��ާ:ڪ��B&�e�5��I���ة�����z �����o�?��޿r��ߟ�
�w�������R���5J)���(�A��ʠ�EXT`�DB�Rڈ�d"ӑ�l��Q�,D�Rh�T���(���P�K���h�d�!��
$��q�D�4C^$����:�\J+��	��\6AeS�?QL�f��.S�l�D�X4��L0�$���9dd�m�W� �SD�*2�EzE$�yE�$`�cTeJP��A�SH���Hf�AD!*�U3IF�@L_%v���φ��G�*|������N��� Tkۙag3�o[��5WG�:{|c��J�Zz�mˀ��k�J��8�,RU�w0U��R�f��!n��w�s�d�-�M���J\�z�H�M���9�f���uU�����3*T=��:���]!v� ��I.mnk�(N�XtVp�C�L!L@�库�c���*����Z2T��U��N�8d4IS)���11	b��
U�㚥n�UL��e��+.أVC��oYUJ���a'S�{-�b���.AY�/d��d���w��̌'pD�rZ��94^�T��,N=�2�fۧr�-�Y2U��_7��ϟ]��F��Ej��'w���d�� ̊�˺��\f��;��%��WM�ǽ�v�����GS{��vs7$U�ӱ�B�CLj�"�z�.�S�w9��Wk]�j�ˬ�d�Fp[���S�����-��K|�u�	{�u�Y2>�[�Ck^�Ʉ��6(g�K��	�j���o����#�d�'��|��l:aۀNf�mdnݔ�N�:B.�휘�+�Afu�;��璙��u��;:���x;!3�Lf�uz!����q-�]Cz��RS������z����h�����7��B�IA.���C(�R�0J�f4�RFOUJI*b
3rRu*�J%�FQ">S-��)� �!$Б�& Q�[%8�hLЄ&��I&�f�8DQ3Q��qD�m� e6��R��e%�R
6�>`��K:�F�mӀ�ˑ!JI��I�L�ʅ�nE�
�q��8 J		%�d��,����TTm"Q!	��k�$�.D!��m�2�l���FI�ē�?�6�m�I��Hh��M�h���l(��9 8�m I����Q8���n�)���KT#�@��b�����	,��"�)�@1�: ���	4�,�JE6A8��N$-��J5���*����E�f�A(��Q��q��J
�Q	(S$��i��E�z�Ϗ.%�ˆ1�;�wu�
RN������sQ��kU%T�j%<m�׎ݻv�۷n8��r���j��I! M��.u���2��7e��RT�N6�;v�۷nݼq�9�*Q)���2,���ܗwB�w7rRs�B�UHT�q�q۷nݻv��q0ʨr�N��UUT�O#�\+����w������t�J���^Gw�ʋ�<��]����U���,�QZ�D$�F�Zz��׏�v�۷n=c�T:J����SP�d�5^N���E�ȫͿ�ƍ�w]�\��ka�F�ܷ6�-����cZ���O�W>+�Гss^my���u�j������T�J�R��S]�\�dJԭCE�y���{��8���G�^��]w����|w��ٗ���;t�N���{y��/N��z�K�ޯ\��t������z5��q�'v��iBD��HH$T 4L/��Ӻu�عN]��ݹuӮ��]<��]-���\�`l\w9�r;�{Խ��=ݗt��n����H�q(����:s�E��뻹W�o��r�]�S(y҄"f�8��Rs����~���$Si���JMS� bA���r0ㄒ�'
`�^_]�RN�S���!M���90^c�ݥ(�Z��VYU��2��R[������֢��f���=����H4#�9�@�1D�i�$0�QAG�'�m�L$!B�h��H�|�F8"��I�`�A�L8(DEl'q���(x�-�����A�.��f�	��ZI�M7XXH �vT���f/N/X��v�$Y��Tr���9M�*���~�7O�����^o_gZ6ͼ��j�j�;�|ydu��b0"�Ϧ <$ݷћ�'�����]��gcBivG�d:������wP�B�0��4��ʨ������4���.C��.�^�A�xOeI�˱0"�pf�����q5+�%/;]��Sn���3 ȋ��������7=%�\)�v��TVsSi�,}�o:ܫ@O��B����;2P؜��1��.��x/��)ո_f�͌���%}���3�#+�����|{�%�S1��`DL�b�oʀ��N�+����uֈK�����Iu�ǧ/�Ԁ�ɩ����7RP��f���b�M���I[1>����2��f�M�L��>������e%Vɟ��X8a���OXP�3�曼����M�l�*�3�ɸjx��Ό��tw����K��+���.h7�6��h�8�+"��c+�[Yn�J���ִ=t�V�t3��\R�G��V���]6g��B �.sـq�C�c�m]�L�y۳��J���Ml+��9�m؃HS��Mv<��wX^:ݎ�g�'�P1��\�{�r�ښ��Q��{Q=�3����s�]��:�oܭ꾾��yj�N���=��������������fgq睴|��3����y�g_����8�Iw��2f����;]�L>w4d�@u	ʥ���s�Lv�|z�v�}8���$N�da>�&U�������'0KT;z��x�;h㘳�T�Wf�o�w�����K6�GP������]>�"��'���Ә�:���|ɶ�淗u���ْ��;<�N�{+�ݳd�Ƕ.�v��kT�>Uq�%Ww8΀�	o�6�4�Bہ����Gڠ��*�v���&�':�SK��n�������JeB,V)����KA�sv$��Ϫ��Ξ������MyuJ<4\EZ��4�n�r�\�:�ch��QϭJ����a5�5��y�Hwv�6���N��z�y�d� �2�{n_@0�_U잫5p��^-�y�B\T�޼��pen8��{˹�<���/9(*<lR�c{��ٱ������ݤ&j�Lr�9��1(Ď*�"��ɓ�*�I+0��v��])vv4���lk��]�lG�]m��h28R;���`u`'b$��Ui�q��n�4�[_ gn����}q��<�{=Hr���s�iD=�bvt�O��%kv�=�j�֜-L�ջ�� �SUg��ɛpWY���h^���M�7qR�N'�՜�^]p6�׽���Bn"tWqx�{b����O;�4;����t��)s��}L��U�GS�39ପs�ݝA�-w�ć5�3/7J��:�d�4�ͥ�du+��(��bwn7�x������ތ��0'i��a7C��;Ƴ;j�<O��Ĩi�`�W5#N����� �aL���ΝF������Q}D��jxr�E'��"�#u�ږu]�T����#㪎Ϣ^��Ң�&u��0`ɔ��wvpFz^�!@��������s����vӿ>F/�e��Fp��ee��W��\FZ\��(-��׌���B}1��w���֮�Ͷ�f�bxs��VM�4!\�W�۷wk���>�ِѿ ���w.�u>� ރ�=��.�u���!�� �~��s�,u�7�UO�ݮ{�=�n�'zᛉm��d;�ê��0.��Ha�>Z)�C'�ʌ4���N4h��y&'���D�����fN�fՈb�1�����F�kU�.~��*�bJ'FY�OLw\����3\^5��Cs���1����L�p�Io���o7U1|۬n��{�
��	{�W��MW��>�9���a�wg%e匵¹⧾���j��θU���d*^��Ʌ�>ۉ�\J���p#H�HyWΰ� �aN��}�˰Z��&z�E󌼕u>�a�m�7yT�������ub����HÒWL֜͋����w��������nO��TIѷ�Zʙaˮ����r��/{3WRIןv��e�W/3�έ;ic!j�����.ޠ�I�r����(���=��r��J�7�wYDx�ލI&&.�Y�Z�[�zN���	�!Ja#�a�,��Ƙ6�Z��o	���_x5ź�{&i������5�Z��R�GW����#@y5�sy�=� �����v�`+�:��>�n�٬PmM=@��y�!�1��t�T�̑aE�1���;ٸ�I�����xv�so�z��ʢt2#���Ȭ�7|��2�����B�w#�~�{�9�.��1�� ��j�Y��Ū�V���v�a��mp��(v�}����֎��8�{+!D�W�����3�#B��ʐ9�1}�%⫻w<�x.ɸתvNi��7�e���w�y�42|= ��@�xUqg��ޫ���]J��I��=��U���qW�y����d��!�	�!׹p=AMwX���)\�v�{m�N���;�y�������:X���t'(i�jZ�#-I�V[w���W�y
��������Y�lt�tk-L5���Ldh�x��w�hk7MN�݋�E�$&ni�ˋ��x�hv��T��Zf�����,u���a�J,�q��i9�BSx4"�MDO��[w����i^5��ΰ۫��L	�+z(9���Aؾ��w�s<sB�҅�Be��0��>3`g6�,��u��%h���W��nH��՞�r�%�y{�u���ܔ���Y�6-�Fk������X,��!uH9n���b�>шfFN�(�m:Z�\����B1�!E��']�C��b���N5�3���;�T�NT5n���C��q�/�+�aݺ���ɼ4I�[cw�-�{�po`wj�A�-���K�_�h�]�Z��!���wl�ޒՊ�2�mz�k��Ғ3qߕd�Y&]�齼��7���5Z;"1-�P�g�B�;������������w)�!�{���m���"}�$`y���_0Rez�W�m)sDڃ>2�R��긱��WԚ�iP�c����H��j��r��w�)���������V�5�\$��DB0��]崵n�UF��h��ձ4Y}Փ^�7c8[r�,��y��y��>���1Efk<"��Mƪ���Q 6Q�n��j�>��/Z�ܼ���P�����p���5��cX.N�tv]��c�ؼ_Q��w�@s�o!�FPS��ˮ�W)F�u����)�l�c>�*�x�}�w[�π���[s��C��h��k���fw��B���U�U���>���o�Mc����h�ȝ�����~��Ni������-���G�k'�˃��ҝ�|:W&s�yC��:_&;�^-=}
�#�������YF����j1�7�}�Q�ݰU\2��g���b�7���:b|�z�O��OW��tzg`�x�Y*���Qq=5(�设�=~��V��{���D���
�!�G]�����C�m��S~#�H�>��&F���C㏕؞^Lڡ	���Y�pg�s#H/�.��'_P�������;���|U����1��r��y�;�hE!Ӷ�\��o�P�X۶4�r�RlP�P`�#M.Y��iYWYaY�cM��Ǆ�+A̳:�Ż�1F��	u�2K����o�u1+(�hY.T�md��AE#47����.gV"���̨F��)Y����z�մZOlG�p"�D�nu�z6ս2�	¤��N����ˉ�����i��X뚡,bɥн{�t�Fn*���wp7�c\��K����ǲ{���J�W��	�K�`��	D	���w7Wt���]�u��u���}��-63k��GӔa"F��G��C��[��XܦB�p�h]_]��v@;�%�}��-��R��x�{8�^�}�g�(�d��$��n{g�f{S}�]�i����}��zW7]���{�E�����@����y���-�l�J'�wwGG�Y���j$.�k�5�O1ե��j@�����YB�������s�Sn7�Nմd^ �nk{18���3:��fMn���]��L^��^S~�i���<*�L�R�}�����NR�&�6�"&.G��!�u쟼��i�ԥ���J {̯1��"Z��1F��w�tNެJ��w�����͵�*�Nڦ�I%�"�S��"
x�4�ɗKS�MV�c��ms���bȜ�)'1o7SW�nnߣ�(�٬���x���� �{�4�)���	����7b����r�����s�+	���U\�����|�����������ף|j*���'�!C�1�븿L��c�I�'�9'L_����Ǉ��
�<�l�.斚�k8������IV+�I�&����+�:B��kqJ��xַź�8z
�Z��%@w�ӡ��|��,��Xi,x�Is��	ft�I��n
��ۂ:��$>��YA�`ɳ�ʧ]n{%��፬=�����8���+�dq�9��>@�	�˛�y����]��aV�}[��^�8�s�lPmM�(�ʭ���s�ϵl��	�$�n������h;��v�^�b����}�G��5�={h{�^,���`F�ݼ��}�<е�ouZl���ʹ>}��n�f��N�*8�r�3����`l{J��0x�v��ogߝo��sߩ�x����#��j�vU�WS�oK�*�z�)C�ܬR�{n��F�՜J�b0ƚ��Ď������]�9VIN��l9�x�,������g6Q��l�syɜ{�MlHF�g#mU��-��KG^n#Pv^"H~�}[��&�^���^D���2[�a�3��'O}�X�<�/4��
o��z�i���ӑ^Q���H}��h��|7��R�=Q;I勻}��"*��	@������Ү|��^���3������=�N	�y�����Z�aQ^����u��Sn��X�ȼ��<���C"�<�o�;�r�a���@Jw��]�ʱ�,������"Μ��u�E3��(*+���'����xl�/�C�
��f�>)C��Vb`L�������e]V��uzIVWq���^枩�z���Φ�]}����!S�	����-[�'�I|j�m���E��n�]>�[ܞѡ ��Rt;��'vy3����?}e��>�_,�}EAҟ��!����\������qOD���Uf��Y��q7� ���&�Z'(�{�{��COp�R�}(�Ƅ�ջ�l	���2gyU���Ŵ%_.a�É�NU�ѥ���/�4�i�*}V���uw9�s6�&֪ε�ry���j�f����neͽ�/1���nIR��hAe��Ve�V5�������.z\=V�ġ�ӂ�]�Pl��wrW�ݞҦ<�ar���(��i�#*Y�n�om�x\�y����L�7p�9��[rX���Щu$�/uu���D�t�s��L�\s���od�H��ë/q1t�o�)�-M��=ŏU���nT�-�8S�[Ԇs��J��OdH��Ju��dݚ]��&eZK+�u�XdMv�t���Y�����g.�E���t%_):�g^
�ڃy	��b�ja�t���V������U:�4��q�Id�#ښ4&��2a�g=qwb٧p��M����f�;����B��f �M;[�y�����V�!-�[Ƿ�b������]�Ń�|O�e�՞\�Fc-�ޮك��[9�Y���E�m��|�
��n��[�ə�$rp&	omC��+�T{u.5]!�Ҝ�2��z��H=�ä��t`���;��H2/��KJ��ˀ�)�θ��V�tԲ�嗇&���s�!*8"�q�{R^��J-�}�H�)�gO!P`�~�F��S{7�˗w�%��97W�&�ɲ�=�䗨ʝ���;~�H<����˰����˻z �2Ӫ;p뗥�6[s7�,y��i�Q�4Ħ�/*,���YŞ���1:iܟ?�Z�6��kM �^�	�Ξ�Yeg�k�9�yU�nG����6��-��#�]�E��y���˼�u��Ҵ�Qt�*�n֙���^I�
l^d�{(,��k%8�8�),�lҘj�r��W�Q����v֙�qe�p���ֽ�'�t�(PѺ7m�i�#jh$t�pfV7�R�]�O^;��2R��P�7-0���Uh���۫;��bF�"��ޥ��!T�`$lb�;�j�fg�fΗ��w|)�;��YV�ca�k\ݤ�:��kdē���n-�kv��� ԍ�Ge+[F���|�v��@����-�QZw�]�zN2w�L��w2�=��ZvZ���<����/s6H�bk{z^Oo���b��s��m�wb7��z�$�i*q�66�foٚ�! �d����*vۃ�U&r�`܁I��҂/���Ӡ��]�x��}7�e���=gh��ʝ]��i�WJ�;�[����zk6ݾ.w_J�����EYt� ���Q�ؚz�MƧ�6��޸�d�<{k���4�-V��UE!�lF�:�Eh�1 �8D���]���j*d]O�nk�R�n��7��]�t)U[Z��gX($^d�BI�%���U�TY�B�k3�xR��8O�G�ĢRH��@$�\��v�]G;�t�]΢Mˑn����n�v���\q۷nݼx��ף�!ڒT�*�C������ݜ������;�9��N뻲gu����t��
zێ8�۷nݻv����$*B7@�wB�4R��i$`�L��2뮻��T!P���z��nݻv�ێ_�������+�Å�L\ۈNڦ�d���]���<��T$�S㧯�^�x�۷nݻz�q��냻t���rR�]s��������feB��%�λ����d���t�����D�������vQ���4\�s�70BQ�2DN;�hJI����v�HCa�PӘ�B1�ݝpP&;�@��"B0��b':��.	��{�����A����N�dU�y��BH�CHx�J,0�-��>�}�V�����[�P��;Ľ�l��=�Q�5��Jn�LfZ��1����4�Ӹi=Yς�TGޠ�����Cۓ;�ә���苷�\�W�Cd�����%�qh�$���N={O莬�go)��򘁑����6��c-����/x���S�%�v�,%�E Mi�H�r�^/?(�mh�(�%+w/;]πN���:!����>����s`LG<��Bԫdʼ�a8����cjD���y{�;y!�k���x^@Y���SX�5ag��;���O��p=k��ׄ��%_cZ���N�����, sɮ�7ެ!{dp�(�E�p��<7��D_���{�1Y'�o��Q�j�1���B�8k�ހ%�~���G��+ˈ#T3oH� OB��$���Y��̉#����3|��i`��x5�;����K�	H�&YL��;�6�C����9M:��3�ыw�wi��C��`��� 7�a�!�>����a�Si�/^���
4�{�XF����\Tv�5*�����<�c�O?30p��:���ۗ�Ej�k��C���KG���A"���Zfч����4��Ũ	�_��k<f�GO��S�r��V���z�Kg��g~�xt�M�Q��e<"~�*o�g4�����U̞�|P"�=7S�a��k��y��%�f�oe�zf� ���`�?=�jn1��ֻp�\�R�
�v��JsN�����ͨ�;�hڼ�D��ĵS"̭���ז�:�_Q�e� �ޯx��z������=�.-�^@	=�� ��6!�����\��pr��X�}��^�5R��`������N� K�; o<У>��^p)�3�A�L"�+�h����ۡ_��DpbV����vh���"��&����X��� WO�-e!�;��h@���2{�6��N�2�.�`���k�[�R�����[?��Ǧ�W�σ:�X�y t`�DT��[ʢ5��'�;��X��F���P�`""��L�%�/�ׅ��]�`7�;xi�d�{�|���!�d�P�E����$��A���x��~Z����_`qW�q43d�;�>6�77f�Od�C�N�!�{�Pŵ��}�x5��L�T8H��,��&�`W���F����S���G���{]�<�1������(w��ht�!����B�� ǄXt�a�ޛ�Vm]��C ��7��X�<6}P;�-�]���v���Cuk ���e�Sz�Ƿ�������s�}��括� �.D�����"47[�8����IL�xKo�E�k�.@w$�jyw�,ţveE;�y�������t���9n��캸�zqn��(Y]�X@����������#�ib��^�����GG[���h�]9�����m��˄�m�"��F�ӰR�ܜ��RG-���;�6�[)���||@> ]b�h�m��=�L�7��Wd���3����`�;Q�Fhrعz�����jڪ�*J�%���Hs oF8�������S�	*�AD�S�{~Rں��&���ԇ����S���	�o`��g��O�>���j5�5���oB��<���LSpI2�. f}S��}{,����F�ױ���zv_�mD��0��_��pИ΀1T������s��PS	}j~����c�� ۀ��7'Y��q ��x�:������m(8��d^��ۥ�9:��z]��&���x����k�¨Z�熳P�Ż�Ab��7���z6%v/F�O?������tw�#�
���X	��@�mfn��w� �eduD� ��8=}<����`ߩV����kO=;��󆇤�H��
6�n�4)�چ �!�,lL`�E*��c¸��r��
`��f5���9e�`�媻�OT�^���T��?���"/�	 s��8�������}^o2R����rޓ{]}�����!�7�~ Aj��,����T(B`+�11��t �3�,���H	���)x���$�����K��؁�Dƴޙ�6`[>�0�q�.�	���,���[f�~5���R���u��+��b�50�T�#���EY��PU�L'L{�W��Rv�>4n�+��W��,ed���/K]��-:�\C�`���oJ����̭��1��5�9L͹���i܍��MkX� ��]HT =�1���9��~�S$��nk�ޠ]�����L�C����y�T-����5k��ӭ�+�*'-{���pT.�W�S�آ�\���s��&��n2�5{�-����i��t���foW�?�<:Q$'���� U?Q�R�6js��dȶ�[d��x�P�0[���"�p�vs��E+��=4� <=��m�(�3ƈ�Κ��#�E����>��Mo�|"�^�՗OlL�ǽ������>y��pq&�P� pP���1 W��O�`)��[E8��	��>(��E˚���yL��+���u{�qr�c!�$t�q X��2.`���G�������Z�{� �±Æ}w�;����=�bޢ�œמw0��ǣ���!7�1̓�ˈ��;tu'�C��49q���襞���|C�)�4������	 � d�=����.J�����n�m����>�+ y�&L��ZJ��N���C����q<>:�\�J\��q,#����k�3���4� �S?=o�/����(������"��3_@z��(^�:���q=���t���*�tɑ�i)��v��^ ����E�06�CM֯E��@���32w%9ׇo͹2�3	��0�`�u�{E�@������N�=���Q��ы�S��W;��e=�F�3���Wgi�S䜭^M��@���!��W�<P"!x�Q�R�.D�"v��e��3�_2�����O����X`�R����q�vԵ nic�*/\O�jU�☇��'O�Ԭ��� .����_���'-A\��Egt�@��Z�3�\�^�[��t�6Y�LU��������]Z�	Z+�"$�[Ϸ8]KIp'�×2xOD.���x{��L��xDugZr�C��Ɖ{�{_�J v�`�9 �~������]�]�d��QF����`��蚒�����l�_U���� "�Š���~�cF8�;�?Zɟx�u��R�W��7�ާD�`��4æI���yX2G��M�� �H!�y�*M�ˬ�n2���6�rC�t��r�Uc�~���tg���~V������ʽom]\� �M�����!�M4�-ఒrOU#��_XK /׃�l�={ GQ�
"���,�11�?V��U�^A��A�M�ɩfW�K3T` <0s�����!�RȖ�`+�t�����U�yĬ�M���}<,(E�����%��.�\dk�\u�����7-�,��Nժ@�)�$�z�ԙ�W��*v@f:q�>�A#D;���a�s��]�����'wJ�J�LԢ�;DE�e2��4�sfY�v-i��j�I[��B��抺���)ق�{��ny��l�P��tr��f���
���f2P�Y���
��ۉ@��q�.�]/*�|��Z�y����\c�1��R�I�eJ��zZ��.a��½��ʧ�b^�"K���(��Q���=�;"���`�6le:j�6��A����4TxcL,�j����tӹ�P�j��� 1	��	:2�a�OZX�ƿ�����Vh���×��n�y��yG=��x&�W�D��p,6��-Z��/c��Z����M�'7Y*�f�"���y�ώ{��{�k�r�IXW���&֑G?��C�|��-uz�T�sɴDVd�{�Nٲ�G��`��¶|1�8S&3�C㿄x�|k`����r,g����>��;�*��������ob���K��S�������)�c��ȣ @��	P8B�8XT}'��L���[�&�ng�ף�b�ə �S�����5�g�ǻ}N�Tv�O��?���4�-GՑ�P� ��50/c����M�}�cx}���G	�8�B�b�j [	8�Ǧ�W��8��b�O�YvVi>�Q��gpԗ}��p�W�#�O�<2�#��K�[���:�0ؿ_D��7�-��c��b�-a1}W��u݂DW=i�4�J��.�q:����9�_G���?-_	ΈR}�K�f�l!Η��w�v"��`V2��d�&��=�U�v8�u2�N�w�-�4\�i��S'��3	�nA� �&�zb#��Ԗ�vٽ��nx[9�������[H��e��æ��ZKQY�r=��.f+	v��\��lvX�'[�0>�i��I~w�+^w���n-U��[��n��R�w���i̘�D봻!�v9���0��^A�L4��֞�^�Ǖ���5W��a�������_sS5�P~_V�g�tm_}�x�����!�Y$1Fm��*����K��>�����T��#�9ӥxo�03E��B6u��:Om���u�!������S�1P}^��m�)����ozVb�7F� h���p��}��<��������t&+��䴄}�Y��g���$�3�n�=������:#����0����
�l�G��6w�]k���s�z%�����א�?��^�"����͟�o�a'!zg���9�c���L��Iv�B��<�,��@{8�5fy3��^C�z�9�JQ$_�Ȝ��:���RǛq�a��J���s"4�2�E{��0�*I{[�L���ZV���덚�����L��1�3�ޭΫ6��_Q{�x������zb��I�T�/]�U\��=e�0l�.S�+L�øfd��|Oǭ��.㩿��{s�<C[5�=K�s
e��q|T��O1� 0�ᡰ�����F_:x\ĺ����r�%,!�V�}I��AJh�$|��<�Iz��Ǌ�|��\9#��U�t�-O*K������e�9WZz��-��u����ֈF�k����L�}���9�+�Rg�`�|7^׺�PO���)���jB�h	�<6�V�Y�/{��<���/ey�c�	��1�Է�3�����)���'�S�N9"fsM�����]�^��p�p����Ҁ��S����8���5�zs��j���ծ��Mt.�0��L9g��~���"��H���f��t¼�o�>�b�F;6!��s�vE���1�&%�ΉO@ݏ@q�t<1�9�+奥�|F�O0��!}�GV���瘌�����;�>�uv�"�f��� �'��ӯ��^��mƥ�S�(Yخ�d�@{C^8Q�rBp�p�������Wt:믇�{�>�7�r~�S�(��Le�q�)�=��lԁ�Bg���=��S2W����Ѻ�[V�pbr�36X<jo\:9B_7����N�ǻ;��m/��Ӧ�����h��h�����KFLy�{7���d&P���Ϸ���3�@{;}�n,�ݴ?olԪ�Zfz��_Ý��n@�ʟԟ�U�ڞ��td�cuL���$F�=�Ĺ�\S0,��B�6o�=���8�[&�s��&O�ԝ����rf��M΋c~�y*�G��s���v����"����R�R��ẆgX��LV(�fw=�O��-��G�Lq��x�}���o_ʚ�(70w�LC�4�Q�E¼Ovv���\��{!��N5n�.�^7����d����a~��2-4�H4�B�@ȩ��������~|���։\����W:�xb��QLh�I��[��/�H�Σo8�J��5s�=r�����P�7O)E��y����9T�u��1���_��g����7=�H}2���U{��Dk�/����L� _H�Wԝ�����Yx�,kˤ�z9�9�_Q�؜�{�W�Nix{XkAp��<��Am�=	"9�.�L����O�gy���z����Ҧ��&��'yk3�����6>������AW��s�A}��g?g��[�����0�*�a�w���e&��1�����+��q
�|ovs`�\|+��"xF� ��=d�ȇW�����J���<yiB/�h����gӏ�}�j�3����$B.L,�����n�oR�@z��Зd�n5�B^1��1�`'}<��;0w��|<k�4_�4�+G>ĸ+��~��w���?�A@�^���ԋ�����0��b�6E�]Ӟ���z��A��7�FI��.�`]�S��bZ�����C=���5d�_
��y�O�HN����;	�d^�g%�g[/��,*Ϊ�����D�W�doWq�=;�T_m�e�p�(eF�U�U5:���t�I���Z�g{oEʱ��]fZ���6��:+*��Z�,��1��T�9�kgBcUӲ�r�j��Ip��˫l���C�����H��H�-4�ȁM4����7��i=s��׸q������P��$O��)��ǟ��yj�T_��CGf�xM>���Jٮ��􀼦Y���{P�3i���Y�M}ꠢ0!���E��KJx`L�ð�>�q�˄D���`�BoD�e���ǂ�WN��z��q>��\��:�X&������C�ޥ�w{#�]w@3}:ӱ'�_g��t>�ϓ ��h%Ӯ,�F:-C��#i6@m�8��G�E�o��C�����(����:�;�<�$�J��&��������+$��z�lk6�{@{��<�q��j��'���a����w��F �s@��;7/k+>v�G��=1�Y�e�0�P��?=������<q
�+��O��_�n�T��I݃"����g�c���^d�^�[7��#t$.��̆����
4ƾ��L���lK���{�^.[�
W:��9�5U�٦,��FB`:�8�sד�l@�w}kg`���\�!�q:�l�Wס��X�&_��5!�-3k�}�V�)�f��ϚC�f�>��KU'|�;�|/�Z�{~]ʩ���s!�{�c�U�+u:�c&�Cv����l��Uоf�:���^�&�ooU���|\[@�7n��a�T��� �/��]�t���D>�W2m�/�ǖ\8�UW��*��Ϸȩ%!���q�V�I�A+R����9�s�f�f��s�Sto����娞��(�a�b4+�y�n�/1H�6�Y���	�!�m�0���F��jvX�Mܻה����A-w��N�ִ�
|:LwB�
F:{��c�͓gb���{��:��ZHQ���ׅN��5HTm^���f,[�k�ۣ���\��I�lԈ��n��aΛbeT�o/���8_Lˈ�fd!�\�Q2��4��d꡶���]f��6�nC��Zۜ��nh��QmNۋ�ij�����vE-؍��d�[��6��Q�Y���A�Mi�+:��Ti�""���ji�GD���6]J�%�Fv'bZ�ۏ(8NK8�6
5s�d��\�v/J�x��y9�4)�N�X�v�R�U�l�k4l٧j���A]dfczV�V�0U����Սa6����$�i�`ے7UF�66^�P���Hƒ�rS��45G�o�hA��*-2�S��%�+D�B0o��4U���`���w.�È�m]s�����V��LL���%m��;`�Cz@Nb���4˥��Թm�ΥEl�I�@�ي�"VҫT�C37Z�UY� �;p_N�/K��̅��0�"D ��bJC�B<i����S�)��~�,�����Z#룼���4⾾�y����2ބ]v�yf���$\�$��w��j
P9R�T`���:=�2U�����»B����$4�?��r�E�����/86�{�)��n;�.l=����{��U>5�mi2?J7�`�jr�NP��pv湲���:*��y e%�Mk.hv��`�TW��^ڧ[�,^�}2�3���nPĻ#H��k�4��8��m�bJ��Ьd��h򝒠Ɇ�-��+goḑ٧�J��;;&a���{��di�E�t(
�j<q�u�*�=�<�Wd�e����w�7ːX���B����R���,����W�|��s�ˋ���S�B%A[�6
�Qv��|��m��GSܹ[9U��n�(3�[�iz#�zLwa�l�Ui�;�St>�WN�t�x�Q)���f�iCOV���J��u��B��M�p���Pʋs��L���dm`����e����~�6���{u�g�h�)T����0m�%?c<���EQ�z ���YZ{Boit��&�����5�r���;K����fj����e��L+!�R���vn��E"NN3�z��{x���Yfa�؈f���k�
�{��ʟ��	������@��\���2�2@DE������I G��ݽz��Ǐ;v�ǣ�����������u�f�κ	1�:���D���N�qǯ^<x��ǎ޽�~w c	0�\���K��M����(В��23A�&��%��q�o^<x��Ǐ^�S!�}��%6H/��q۩����{�0&��"���q��x��Ǐ=z=revD�#B`�i�`��$�HF)����",h�AF`$�2:�J4���\$�F?W�]��'ν����Ba��$�|]A��vf�%�C��ё���PiȔ�
�C/;.����,�6���D&2F��LJ�J���׾��y������Ē�J�d�c(�F�a��M�pJ6� /+͑ˡ��-<�q�kv`��[��--�V�ԉ5�c�R.S����f������6IOw�����9��M�N����@P^N��L��,Fل��(�#�2�(��a�PH4�m \j�m�m�!7���@�E��A�M���L�p�����С��@$��I��hP��  1D.���ֹw~y��ϙ}W��s�$����ܳ$	�rU���f
5�;c�z�-�`Jn�a���a�'C�k�7E����r}a`��DH�]}��,��/o�� �"�_Ъ<wbI/�{#&�Rq��K,�l�5�u;���Mt�F���lVvr�G��2$Ǆi�x�
߬L�d���4+��%�Y�a1�=�Jq��'he[��N��z���a�_'��-��=��mX5�u�~uŷ2�gf��D��'��P�[�5��,��H��%�?4S�����	��[{�d]���ʺ�Wx�Q�̤��b�hˌG�/�$1j	d���<��!���Q	�HW�މ��ܢ����;2lG��tl;�EE0.���ЕL	cEu7�޼c����C�7�Q���Պ���f^У|ʰES�gN�>6������||�_ ���i�Jr{�,��3\����S(�f|#O�
|.�y��5;��~�N�G&���5ޒs�_�2Й�y[�.2��dM�e��|�
����#�~_�7�A��k~���껺2�:D�'���G�^��S�m�#���R����ɻ҄f�1æ���|����$��yqՕ�p�DP�Ғo�R����M0�Z�:ذ��Lic�@��ݠr%��p�i=�Qꃠ�{��B�qUuJ��7��f�W��u+_B���@�4ҋM4��HH���+���s�µ������n�q�OÞE+���\��ަ�n3�Ƙ�BO��T����S�Em�%6��f�u�3r�4�ͩvB�I/~�Ⱥ�q��S@�V��EzUDdg�6-�Nw(:B��;���4D}�Q£��{� ���*�<0,ܢ�
�Ƃ�P�Sø�ȋ��V}�A�K2�`�X/��UL�;�&v:��P�{[�\�i�0�@xB�tY����tu$�M�ie��W�� �vH�9�D�wjE��������s�r@�C5D�0���c�wk�I��i1�9�0^�R��F;̎���p���:h: �tP�'�*�8��Яk?Q{��]w�^g���"%�C<O*.��v�P�N�,ZC9��4!0�<F[�;1N�dV��zw���7���n�KW���wn��i�DK�@�pμ��\V��1ua⸐��p�.&�)n=�yr�n���
�z�/a(4��f~����qC׌�Ϙte���}�mm��C�3�p����%ϸB�NC,�Ɵ�6�չ��B&���.�}��c����cA��*C��)S�E�z��r�׾�����n�?RC	۪��8�)�l����D�\���l����D�^DE��}�{�Ҫ̮�V���MI�eI�%�)������ŅG�a�����z>�M+v��-��w�nUA��Ы��H���M�4Ь��4�*E"��|�����{��{��*��\���(S���_~^;�_&B��T�m�����om�R%�NQ��Z\u���Ͱ�su��dH��aAi�Κ����7���=��Ԥ�]���U|��+о�YlKٗ R�`�F
��f��� j����=�g<z�.��0n�|����l��GLW��B�2o��=_���Hql��n��oF���[��OWDC�����}>��2��px�+@��L���(�a^}��^k��Ɋ| �؎��싧V����xL����]!_Aw�y.�!ʥX9☭��;��]���-�7��ɶfd# �E�O�rD�H�����t@��_-���2��X��S�ȭ�Ԥ<�l��;���g��`/��_0>馼"��������]�P�`}3��i;2�{�I=���bЇ\�4=
"~۟��B5�Ktz:�y��� C!��F�<
�w����Eu�º<g��P{�Oa��P�6Xe�A�"G�E	���5�>���j����<"�!���eFĜ1��-I�U�C(qژrvzKCi��;;�T���uN�ͿZ((�z�r�me�li<��K
Pمt�f����e����'õ^�ۍ]N+��`�MSY��ޡ�-aeh�����<��M" ��B	M4��J�ȨH H�H��7��>tJ�S3��yn��S����K����a���>ڇ�r�Q�;���0��?lTz����3�W���t�'�.��Gd��cU���H^�.>��gC��xsq�C�C�K)�<�ؓ�l�k����Ӑ����O�I�-=�|d�$6@��a#6	~,��=P�w������]�)�3i���c���3�fx�<E�4�~=�u
�{P����
y>!cCz`��i��^�
צ|�^ƙP�{��4,J4k�H.G���إ�w�f�ux�hSro�@Y�,��*q�j(���/��1�6���U�1=�R�W��{�v�p|Ŷ�L��
�w g�8�)��H�5�Cݵ�!�p�k��2N!�[��cQ���w����)�vL!���5Ii1���=���̬*4*��qel3�q�{�������S�T�У�<s����4h��g�0������(ǁF�[o\�'o,��#�Me�
�.���qM�
��|C��������@��T���&+e�Op���m��Oj�E1Pԣ;���a��m롇X���)��&漶�VN�a��i�٦l�Q��C{:��7���$� ���"�h Q����l��y �،����E�RS7	h1lj"�n�#��;�k���n򪐃Sl:r����5<�T��C�A��@�M4���H�AR4Ҩ� 1B�x5hk�������Z;na�F���C¥NKrdbn"А�Xgu���a߽uV��z,��>����
=v'�*�(9�Y��2_�!]�.3
���e��E�_E뢚7��4�I�#4�'�<:p���=�i���N,�Ke
��lb����R�x�fBc@�����m�;�׶v�Ϙ:�\����x����2m�W�D�5�,dF�&��I��L{�Uڟ*��N�كJ��3�>�ǹ�g^A>dw�"�+�p�Ծ�M��^��4s�+}z}U�3��[���[?�x�[Ҷy�J�;�MVh.Ҫ3���:X�÷���E�vO�`n_My/)@e�L(��r1�zT��v�Ǘ��K;Q�� 1$^4fDi����?D�8�J��D�)��Th1��P�V���X��;�P&]���z��ºz��1� ��/��ߖxC�j��쑥B`�f�ou�N��8e��^CzO=zq!s0{GL4�ִ�֢���!�q�"�@'��Ȩ�jB��Y�Y�̓s�j�T}5xs��
�n��Ź$7+��3f�άlgW�^��:b��%O<&�g�1�^�$GK�U;�Q�9��yT�l��5P��u�Χ��
�g0����FԪ�����	>�I!]�	�>�_}w�O�>��!^��%��m\༗�7ń��n!βV5�q�q����8N+&�7
���97��˜�sr��|抯�Q���H��F�i�E����H��/����=��3�}+��k����)������qwǵa�=:�j���i�z$Ә*���6y�5���s���sb%8�༗�Mm��������t5劼)n8V*g�$���_xs$�"O^"�(s����O�A�q���8��64��M��e�7���!���}x�]���h*�\���dPr��VO��
�P��RG��s���1�7�el4u����M ��LW4	/�&hP}���v��s B1��~�Ƭ�z-��V��kP�]q�v]���'�1L���Hy�b������5��m�6��U޹J��6�p��l`=q<c�5"wC��U�<���7(�NX�.5;�q�r���=ƶ�^s3�����$)��;c�Hz���U&GM��|�fqUm�V�y��r�"SD=���q���YF�;�A������Jcs['�dR����ǥdW�:�q_dt�}��W��U�=W8E}����iw E|A�%��H�"00���0O5:G.�}rn��s}1�d
�M�ŗ�'XHp9X{o9�jNK����H�MµUt�\�[qy�8{}[>�v�����6�)K@���^��sn�O�6SoE��j��٩;�g%nƱ)C�W:��Y��cu�He��*qT�ʓ�B���� ��B�+hTi���"Ȭi�Q
D�(H����yϜ�~M���۞�+E�R"!�߀k��{&�q��>; ���̍�("���	��¿I���]�ܟ/��v��w��Œw��-#63���L7c�x�a�ƺ���� `+nک�������c��LUǈR��˒E�)�E��A��3x�����K��i�D��]�d3`��B.���M=p̄�x�/�}����CB�y|S���t?T��}KA{~�~g��x�d)�;���Ͽ~b�d�����*
3��C.t���^�TՋ-wd��{|+���@��DX���l�U�F< #A9n��)���OC'��'�j�;a+�;�<3�-l� �	ʖ*��v�^������\I���<=��(�#ޓNN��*;7����2��l}�7�S���&PTϓ�}�~�{�|y�=�C�f��5f����3�g��K��ڽS�d���! Y�Fu������b�S�(�g�P���s������`z
��u~���P.@�LL?X�t�-�6��]0�0��yMu]����t�"L^'k���gD�[8nj�f�-�vwZ�e�ɨ=vWA��L��yV���ߠLˎ�*�����a�����<���ig�L��7�Y5λm����MC���Ձ�:�fą��}��o���]��`��1i&�>Υ��z-�q���������R�$����ݺ�nݺ�r���+m��""�
2 	"7��fw�^�y���� �^頃b6ؘ	�E�4�'q7�z�ū�m��C��,7����VԻ%C�P9���}��t�n�	q��x.����j2*�A��N���9��S��)���W,zt���cv�b��ʒ}�&?�ts�A~��9�5��?	9���h�r$���@L,~*	{����&FP [�����~/&�a�Z�l�Rm�bX'��B�#�8�ᑖ�}�i�o����e��^�PNT
=5�P�\�,5������.����4<��ע�sU?,�[~(ܬw�@DC�\^���y��8="�w�);�>V��6���,zO}Q1��O�'�uk�����>�+a�PT�Je�Y��KS�Ǿ���0�[�o�"�9�1:$W��>gMLq�*��?ZkP��;��wG����ye�!5#GwӚ^;������
��碱���ş�r�}<�V�
�s��z�$ߕ4Vd��1������z�l�v��l�zE;Ň�a�z��UD��B�m1���/�ݺ��A�%��l�W!�d`w���}(;�3���m�o���i��Y�f���o�o^�st�q�����Tc���ܜ�h�Pp�-e���#:�MiFVԱ}g;�Eյ���2kV��'����Qu�4���H5�H7-��M۵����[UoG�����K�-����tT��x�)��4�E+@�&A"|���T�i���	Mz@�1Y^�WNߜ{��cռ��6�{ �O�S�#�;���KlW�w��'�	|ʀ��M����1,���z>r��T3T�`�Yڢ*��t,��?e���rԘ�{����2��Ej%;(�Ľ�����R)�U�[�s��]��{�P��k�F5H�!Lgl�C���t�8GS�؁Y��tf���p�&yw}�}��cVc@�C�sj �Yz��y�� ��C�	��d�g��ަ�u���U+w��Ѽ���X�׸����#N�lS���R"���ButT�(֑�r8$�.ru+}�\�5o�-��Q9���6�sµ!1�)������?�������@�lX��³�K���}�13�=b����z2&�,q�7��(2F3���>�����n�8h���M<e���̳s5��HdC��뢾�9�SDNU��mi;Tz�}��s cOE옚E���nK�<�����d�p�L�M	�=�U�ߤ_���!��oŎ	ގ�{'L��
.��8o,�#�$��=ؘ���hr�k?��^�E�S��z���G��ۛ�m���N*�ʳ��.s���nm�d�uU�'���zz3��ʭg/:UX�p--!ʹo���Y�E~#63'z`.1]+rn��0��0���U}�<�����4
�#M-FAV4ЩQE&��浨�cm�-�Z�ff��� �H�1�/�!Y8ߗ)Q�����3������wV�~�{������l#�J���;�B^����o2�)��O��û8"�������P�yA�4P��>���ĭMq]]�5;�#�[�~���*��[�]��|FS�C֤���o[!���Ǆ�;18n:�jպvd�ўL�1̋ߧ���.-�b��Ł��W6�d4��G��f:6o 7��j]�}���Dv����v��K���D1�=���s~���	cEuk �v�f6W�v�M��Oé�]Z��ř��\�� ��@~VxӋ2.g�{>>����YG�I��1]o������L�P�:����R�^�ޏ(2.�0��y٘X�a)��Ն�D0��{{�Zze_"���^ȉ�Et�|�}�]�6�w"�F7�H{hN���!��p��kJ6�?�7�1[�>��������E�ƅخz�q�f1��9�c�l��s¯3��5�[��f�Ї�7z`�Ӵ�ڞ/��t����9�g<����z�+�j��Y�5�K���O�t��.UE�&i��w�b��o:k*����Ʃ�Eֲd[�ۻ]yךB���K*�^���Ss}��R_6!U���lgǛ{tmk']��jI{�v��i�I�GD��n�X��t.7]qH�7x]E��j�40�q�mc۸�eގлS�BN�l�y��ȶcS')�9�g=�U�7u�{ڌ���R�&E9Bmtt\ݕ
�s�nm5��F�'r��ڒ{F��
���gUcQ��]�XMS�#Hʏ,�7{�8J~�d��eQ̜����CR��Pi_r�p��]v���:�K2�BQ�u��3�J�+h��7	%xA���UbBÃ��V�Uh�K��X���I�0�*I�$#�)�E�W�:KaV �`��CF`��oB�^���ne�֡���*��=[�s��J�gef�u�fu�{�\��Fee��me�qI����b�l����S��t�U
��0���s{�Z&g<�
V�TV���۪����[ê�mATQ������:�j7d�J���5^�p�!��ݛ��x��)m��p�F]JV��>;̥[��]6o�Δդ����1��Re�I����D�4J;5���_d34��1���.9���x/�F��]�C�Sb����0��Z3�6�r�&���%�&����F�<v,�!�y(��R��T�]@�`�b�1�y��"6z��` ��Zp�N^8�~ɑ���{,.��X�f�n����ݦȫ��e�I�?eu�6�gv]j,Ú	bկ��Ng��2�ʽ�s;��t]���c�Ǒ�*&V�W="dw����,����s\�K[e�j��Y6�/][ihZ(��&Q�� ��bQ�ÍM��]uؘ�5���Z�q²�&����겪�f��y�_I��멹����W(�a����!U�=f�%��~[�����Zo7p���8�@�[۳�̡U�1���N]�J����8�C2��.�eQ�#��$�5V��m;���u�������Qo����¦�.01]hH���Ų�)\��[9],ΪnS{rU,λ�n�[(N$�
S��R�5��!�g�JKj/lU�ܽ)d����f[��Y�0�D�ۮ��v&i�����pXR��N�C^+$4�����t��ʭ���H�q�E7)Zۇ�ge�*��NdZ�EY��^M�7�zVt7��Z͔���19ut򦍺�2�ִ��B���kzb�Ǎ��9ȯ��Lsd��e�-���=Vn��^�_!r��
�£����e���}M�.�΅]�����m�����{k&ʔ�<ٔ��dʬg��h3{,J@����dQڷV'KZۖB7/Eva���A�(Wv�}kR�ʘ
Yϡ�k�LW�r{���l�����'	�L���$# L�!�2�C(���Q�!�A�#Ǐ��z�Ǐ<x��ף��!!$� �'�Sʧ�	HA7uԧ��5#�H�4���8��Ǐo������ߺ�I���6$���d�(P��e�2�r��|ݽ�lq�=x��Ǐ=z�2!	2M�d��r{.���	�\�E0�hL7�oo��x��׏<x��ׯaH�W7K	�)���{"����fe����D�I��wu���!"O�\�6+�מ&m ;���dI)$�l��sL@��L��
�E�R��R3F���(ĒY����6I_mv�;@NWD��)M�l$\�)1�lCd�&�����
)7��_���������w���30�R���Ō�R��eۛm�r����Fu��
���t�\�#J�Hv��
�����*f���~���F�i����iR�� H� Ƞ�	"U���%K*l`�~pq-lC�ɻ��hW_��0��=�;٨E��sj��ߜf�qJ���28���Z��|�����!y��L�֞��?A�p_O|U-t���L�by�gO̭�V�͈���B�q�"$@:�1�Da��;.1�Y�P�ndۅ{<��{��;����z�yat4�/mr��-����n��w��K��� ��z���iB=U���d�]��'�+l���3ȏ��C�;���	���擰W��zAw�g��H����~-oM�/�T�M�U,��0̋ͻ5��TXV�Iz�v�s?�����<��$��{Øe-�ݢT�^�7LW@B��S=�萜*��^o�y�9� ���HX"ڞ�ݜ�bo�l���/A�T������@t/>�7�.{�
���S�أc.{���p���`�Jո�ʦ���]�ڋ=��Pj���D�_�wr�W|}J�=�!��f����1��|�I�ᾯdW��s1�2Q��(Y�c�����=ƃ�u�T^��o��0f3N^����\�����Ȝ�8��[i��W\ȁM�Z�ً�{QrMj�6��e�ӗ&;>��Ki��wn�5�ꫵ���;rt�7+w�$�L����Z,s/P��I1sX̨3����h,fBWb�cSj��hV�EC�|<H��f���F�*"H�R
H���k�n�Ͷ�Z+cj�U��� ���D*����։ƻ�C��S�)�5�B���z��V���|�ҜK\)���a����,�����{}���%5i�N���1�[�U�k�:yJ�X_���3ks��w��*�Ě��FC���8K�נ!��@ۙE�3��#S��6Q>�Üŧw/9��{������s�1yڢ]s���\�&�����"����y��&���y`:c�Fֳ6*o��^/�2z㊈"DB3�G��Bm�5�	�:������@zD��+&(�3�,�Y�L�b�C��ƽ�X�=��ԧ����S���s����U�RTs�`��}���΃fj������9�^�<�H�~Y�M�.C�^�R���R'�.�VX)g_=�ݻ����r��S"XȎ4XP�R��r^�ϲԉ
�F��#c��9i�-�ϕ�����Z�5K�=0N������]�{�իƑ}~�9ʞzprء����/(=N%��}|	��C��S�[TE�r	r��я���+�@�q�o[Nhҕ>"m����ƂԪR�(�ڥ��f�7X���jxo΍�fH�^�j�m�R�ǻ����3/wx�`�4���8����7N�*����gl��[T�s���V;�s�Y��dT���Y����6�{�]�y[����} ���J�R4ЅM�����ksSv�m��)IDEY�D�$ >o�7~�MSz�=�����V���*-:�n��K4��;��ȃ��u���"0+����&����X=� ݽL�i�K��K^Lr��Y'c_2�CH�h���_W����,�O�����z��c'|�KN���Id�42v^�gs�ڐ/�P��<�A7:�`c&H������f�+,>0����zr~_mk'�����9j�U�b�s�zl�R3ݐ�$��G�{�����0\3[AD0C/'��x��]�&m�,�Pc�&$z�v}�Д�ܥ�V���ct{c�yk޼d<ݷnOojR�v�ԼO��u14E����3�`�)�}�	�@�i�d��SL���5=���x��]Y��UZ�}0�}q>�B�/�D��̀ ����'��>Q	��O�TYu{��d����Fy����D(���c�g	5��.,��We��Td9���x[H��L?SQ�:�V����Qoq���ofA����/dAe��y�5���sw�E��������G�Ȅ�Bc�m���f����[�S}�!^�<�͗i��Zc��~D'�i[�#Nİ�;�?O��?�Q�~	��uf|Ͱs%�mr����hVJzFu$�=�d�g�Q���ȃ�{Q���3ܲ���VoN����Da���R#ў�ب�VMk��
s��� �Uj��A�DE�M�����ۆN7�r�TÂU��Z��AV�e�@��V�S�K4����~����ƚTj��J�F�E��0V"H"	�o{ƕ��U�eX���ʞ1��A'��A��L!�݇�FDb#0Et�ӆk�f�Sko�nW���l���2'�W��Lv�,��>�N+��O��|�\�ݩdb����xU��X8���p��i�5�ïpyj�N�����=K�dّJ���mk��Z�=>	'����g���}'��T}[�1Rp�V���v�<�Ůt���%�kf���f�in�y��˘!|�%;�����q��`H=L�4>)��i�ֺ�c���d#ѳd�#3S����w�k���@f�W����"�o}�_$GX@NZ5Y]6
��D�Ý3է6�&�}��5 �]d!/5�E�xl
�FWH��I/I@^(��fp��i�R�V<��HfkRz�I5J����@_��'��w�E���%�ƣK�ɐ��-�.��Q���ɦE�e!�t�[Qy�W�c9t9�=8&Cz�p�B\��3����O��"��^4���b_Lm[O���e�����ވ�b������}�A���)��vl�9���Zֺا����"_�V*{����E��sN[�>���p�)߈w��
����h1���f2DF��c�P��^�z���G^1��t�NP�͹�ms�j�ײ֛e!��^�Pˋ	<6i��%�9vkRR���g'�&���Wo�@D#M"5&��W-Sv�V��Qm�X�@IA���g|������ɐs��ը.c��?Wݎ��=C�S=� �����v8!�w2f �ŷ���Z-l�"۹��%դ�%S�V�6m��E�*�����;PN�����&z�%��g�9]��@��*�,J$C~�E�4)�+���v�®�r{�/z���۵���� �|S ��q�Ml�����{���i�d�g�����6�ٮv�D^^��.����+��!���Ê���9m�K�����/�0����B,��E��F1��v��������agZ�
��L8����Hw`�|"m���<�[&A��V�TXfq�֬Y3c�x����Yα���^ݑ��9ZLj>NB��zx�T�="��|�:�
�(H"s�x�������YRu�% �l�(,$f��C����(p^&�>����y�|6��z��]ٌ4��LM�T:���=�g`q�GA����DJBW:{k��=>��Tj¶;�����9/~�fȭ4�V�Iza۱���~�<����V�K�Tu{�d�UP�-)Zyr"9Q�*oN-.ے7��ف�h%FZ+bgUM�����j-@�刈��"�__M92��]��;�u[F$��)��j��mV�˝�W�N,�s����V���I��?_U�Թv^�x��u��w����+M�-��v���V�Unݺ��-�ZƴU��f���E,��G��#\~xh}J��dS�g�!!
�O��y�r����S�C�N#]A����KY���w�)ᶇ4g(!���}��{k�<�D\.ym�I磟�x��O�VϺ��ꯔ�%�X���Kb��SX[=��2AԸ���/��@��$c �h�u�\��r�_r�a���@��Խ�!e�"�J��E|%��1��P�9�n���a�.��Y�۵�8��\[�yu����c���]���	ę�;B-����0�k�Tѣ�N����{�H�S�5l4��������h6&���d3VA]�K�̷>2�۾��6�ʣ�@f���1��D��,ǯ6e&�1�mi��l�L6nw{Xu�)D�2jZ�p�.`�nz�������~et���Aw��0�`�R��A�Pm:ʜ���w�L3W4�بr~�-���;�G�Q�~�jc�6�@�����/�tn;�՚�L=��f�n;��z�/^�d������8����hp��u��&֘�B�)�K��܍4�i�;��1Q�W�N�UU���Q[��6I�sw#"g�e�S'ы�=x���d{�3�z�F��{��Ȏoz6��'F]'q�"�&�	��V���/F��#�gK�27(������Z�9�h�>�O��Q�"����M۵�Y���r���d@Id@d@N{����������=���N�,qZgU��5jBH+jC5����FfX��Dл�h��}c�w=r���������F��a���{��*V���;ݳ�R���Й�f/�)���J����R�J�^���tc��AQJ;ܩZ"s;:}{�|���H��0z8И��-��u3*s��vu��/��q��8���R/�ow\���~�h��0W ����}H`����Nj�����#�/P��]����>���*#�HV�I^�ω��j!o�'��ƃ�k;�C0r�0:.Y���,�ܳ/S"Lg��W��g9n}Q~���	__S3��x���p���D��8T�1Ǻ$ӌ^��%�)n�s�\x����yyz�
�	�4��|,}�M㿕{����Vh	�l{y�x5J+�ٌ�2K�<ӯgY�F6��S��9�f͋�N"��R�6L]���:��)�U-"e�u˯�raг�G?�=c~��Sq�dl��9�%5ޙA�W�D��WN��z/���=x����;wju� ;6����4���Ð��m۝��(TK*�$��k���j��˛|�_�"i�y'm�/Rշ�w��i��X;{��Ҥ���NYy�J�L���Ъ���;��@ߦgތP�̧3X�,�;ǐ�(޸������޵՛q�9�v���������Y{n�6�ˇ��3��*��̓�D�񥨄����Z����j��[��EF��QlX�5��>�����d�r��?8+�qg��3�q:���ИL+h�6����\�{�oa_�:�z�^�c��Q��� ܉"���Bf
/<L@�~�n]��4׷n��3��l�3����ft���TO�ʞyh\Ú�E�l=�[AG�9�D�*WT��}��ڽ(�V�!�l磰��z�){���'��+y��6�����K�[Rv�u�t5_|�7��Z,��'�Ľ�*%����<ףzU�W�d&0�⣹�����d��Ooj�u?n+���'3�^�<˞�9nQ5�z[ށ-�#v������)T�y�J|�|�<� S�9��l�˳�wg�w��A��"����+�VC����E�+�F��Q��?P\�mi60�}Y쎱'��jc�.(����z�d8�6����#�
���x�Z��N#�d��̮�%<rY�@W�{ȋ7��ӋM�i��;+�k�K�9b�Ƴ��7T<��|�-ƊU���N���77O'|$�vP>����'W��f ��"�'�)W�b�yX���	�/_}y%l�G�������z_-��d���Fv�k����d�3�y��b��w;���,O�֎��˲��W1i��s����΅���/w�V��jur��j�v�D����v����Y�<�:�XZVՂ9��m��32������?M ��J66nݺZ4ݝ��h��H �� H�H)���|�T�`б���/P��Ϸ�������&���{jME�ѦTO�-Od��������� ��M�Y܉P�K���ߛҋ�]dpj�t�'�?�4˵e�q�5z�zv�nF���zw���*�BO������	�"�@]>7k��_;^Fl<;��r��5"�i^��Q9�^�dg�����Ј��u�p�Θ����Gz'65�>�ye���Di��uUjy�n;�]�����K7�\�и�xBz<������.�EHy/}��RV'�pUű�Ѭ�����r����o�|�� �;r��ڳ�Y�Mb�3/���nӟ7�J���(�<l��C;�¤�9�J��"��+�
��W=T0�w�K+�tq�sW� 8Td�z,z	us�n��W)�ojx��e�Y�Y�k�x\D�2��]o~GՁ(�)o?u+�_�i����G��*<u�D���4TK��la�E���H�����;=�V5�)�C���֨������㼙/�:�}<\_� �1���}�,�Mb~�}ҋ�W;��V�/��y���Q�uvy����G� �3S�ϧF���l�Wy�E �JFs2.�J�3�o+���{����er�Z6�ŧqE|�2rl�Y��GW't��ա�jL�O(���z�<�nj�a>�d�d?f��!Sv��v����v��QA��Z���ō�~�������;-�P7yK
ލc2g|�>��zw����1��㪤Y�F<9��zVf�:�]ΓJk�\_��eA/l�N%��.m�5�V����6X^����E�N��V�x�ۉ]w����f��nGLD|o�nE���Fu{+ϨY����(�Hg=�������g%m�wuC;��	�$D�8���:~�	r���,ْ���.�^�@��%��b��&w�uev3Uhk>���x���@A��4<��{��A��!܍������'��?qU-N�:^�t���2�"�K�=z]_�@�~��������]0�Bp�p̧>أ{���J$�����]�I��rd@�k���N
ﾯY��5B��8���%�j�ĸ��y��Y��Y�ަ�V�2�B=���!�`+���R�ϜT�f�u )�,�bG	�>Q�����VNq�;�#0���1�'���%5�]��`����]^��${f�=��6Y�B�7(����c��KlW���}^�o�s ��a��Z�i��:PމN���0IT.�&���k���<+/��������(J�IWb�`�IMM���(ޫX�!�uRõp޸�t�T�Z���J�mIᅶj��ۋnDձ!]y����u^&N�ѵ�T(`�G�;����>�w;[�����37s�
p0�m+�&Z�����/��j����o�1�L�m�*�bݝԞ������Ԫ��r�*bQ�v���U6�s�mT�E����P��4��Ų
�
���KU/M���1���gV�-D�d��^�Z�z�sv����9n>��(�Y�%�m�ܽ�=,7|jM�q��PDy���6��5��Ԏj�K��r��W�se\W�)����N��:��x�:P���l���]5����� �̤�KIn�D��"J�˯�+�Ko�����$�����p���{��u�9uj5Y0Bs-<j �>wuf�M��Sq]�gu���J�2�e��+21-�ẇ9���Z�����u���y�-8���޸��I��v �Lp>��2�wm�[�t[S	ՙi�aM��DW�̥4�F�:�^ZT�%u�C�T�m�"��g\ɸȻ�I�ԝ���m�w�5��<դ�se�����v���#Y�QBc7 �ox�\�(�]��[��Nl��UI��N��؛�P�I�BZ��iF�{���/E���lS���^��mx���'�,ۘ��������}�*�X{�E����rrO�o�Q1��ܤ�Fk�*G�Laɢgr�/����]��	�w�%(Û��8�4�.�r��֦P!�˻�lT�[����oXv��*+;;��i�h�/�uѵ{�M�C�Ƥ�����-��ͳ�ZO"��/�����%أwV*{B:��Ռ�RY%N�
���\<;f9�ּ����skXo^m#��8��ݹ0&�cA��췍+$�k�i��2�V;��Q��N�%Uk��oow�һ=�T	/d�k��;]h�SZh��Y��mm�?m�(�8��f����Y+U��ד�-�z�c��g�5T��r��i��j>�q̸�����)�E�������ĪR�H��(sgweҬ�hvf�
����}�$���pr`�#mTV; Y�[���}k��y���N�.?���qjpŋ)<���r�)7do;3jR�B�WeFp���Skڶ��ɳ6���[�2�jb��Q��\^0��c�;\�Z���
i��3EbW���٢u|���Yq]Vs��v�f��cm�;�E�Q�{b��N���j��eyU��ά�����+����Cz����y!f^ηD伌$2PD�R���	n4'�0ŵ��텙h���`4�@WL7Px's�cc5�,v��A�4���	��V�v3oM�\sm�����oe�5UUuoWUg���(�L�&BS1c$L�!�$�L$FIB�n�8�۷;~�<x��ǯ^�B#	#!��+{�y\�!1�LL�2��H�t��qǏ�x��Ǐ^�{��BF�!$�$�HD����6��Sfc	BI$����|q�<z����{�}����u���� %o�����	�DB̣S&:q�qǏ�x��Ǐ^�;$d#3%b+B_��F4>��B4�&d��T�&c�f%H$LbM��e%4&@���Ԓߝr@(f���d$a6���	�	b�b$���&)	�bB#>.�&Q�HcD ���0EFg���޺!����#h>7i��]v,ȫ��!�F� ���&̟;s!A&2"�K��21D�o�&�I$i;r[v6�+�`. $��J�IM�I�����9W����$A9T�>L�1�F]���Ք�nV��];w��Q�:@\ΊI��<]k98⨤O���ي̵�/� �{$�&g`_�6YoѸъ	 ��aP�F�AB���P�!-�C��"Rb�� �2zIhQd:-R!i%t���$�Tp����SM;���?T�����+�'�TֵvHU���Y�iB�h�e �i�jH����~]���6Bݭґ�i��e��"��ޫƧ�6�?B�B�����~��e��S�dCf= f̢�<K��*9��w<��Е���{�϶9��o��n-"�ψ��_���+�������.H͐���]�/:�\/y���ݾ�s��(��j����>2"ȕ$I4�2�7M�0t��ȓɠ\C���jʌ]��tLQ{f�E�!������x�|�v�,�(r�5�ð;ϲ<��64�8F��c���Y�UZ\4��p���Lk�h��I�>��zmE�]r4��BnDO	�6E��+���ξk��'�ND�UQݙz7g�f�%A/r��PEH���7s�CD�h|r��9�0e�c�(:ǘv.Z}���e�xGu��O�dCN?��k^^����[���Ӥ 1�r�l����ӑ���Q�g�5ǫ%��5������y
i�6�=ъo��/h_�= y�aaɬ��C`��t4��k����YX7�%'�2�^�fr,!��jz�$�L���kڔ���?��\Vy~?� +m���s�9l�4ri`�N�_m�q*BdQ�P̊���}��#{u��e��V�ݧ��;�8G2')�̥�OU;��/K��;S�n�UL�V.zx���2���(���mɒ��P�e����V;����7QVOV�ۊ-ٕ��_�f��S!E���*,��i�h
�h
#i���s\��w�<�x������!م]m	͂�B5�E������*�-3%`X|a�����\�y��[*�Z?F����)�-J�+� �P��,Q�y�i���k{nF�4����~��Q�
���L�ھ�q����ϝs�%CۮU�RȯQ�+���Lr���=�Y��=rv�M(��w��R|&'�lX�B��>�}:�6. i�d�]��]4b�լ�n�שd����ϭa�v��R���{������_�%H#}��	4/Ed��}��u'r-���O?O�^�l�*4���G\�Ǩu�ty���JD��eb��3ym[�v���	�r���ƍ$���	ʑ�"�S�9��M��� ��GF0��ǯ�Q��oV�Q�6��L�>Y"K��i��P���2~E<�sH�F�ɦܥ��j��D�;	��8mn�笏"�p��w�ꘖ4�=�@^����ҹ��La�~��'�q��y�ьD/ͬ#��տk���C�;0�>���=L{��s[�qu0hƑ;�� f�/�C��W�Z՝�ʥ��`��F*��%��B֛�~�yN%�:�
��˙�4�(u%4u#JC�s�r��[W+m���SFW#�҇�_AΪ�����,{Zq�5�LI�PM�vm�'M�b�6�,��Щ��*.�Z�A��yu~_2��f�$�0~Ϗ�M4��U���<��a�ag)jR�?c��Ƥ*�2��(|��?(K[��qi�,ȥO��7eB%��fC���kI��N;n*��UA�V��H֡��h���3��lʏ�6�=�<��N�Uwʪ{Tp��]!���'>�i9���؈=�8\>(���U��U�����DT��ٙ4��צx���d6�Y��[�|�w�=�F���T5Y]6�p�:i��Z!S����b�30L��b����Ͻ.���s��	�_
W�K�S�5#�8XC5��4��KT	J�Y��u}y�A=���5�2ȁY�C����h��K���Ź,��ov�:Rk꺷����A��؞�rf��������~PHC�VE�M����U�'s��C_�IN^.:�YR�Ư	u{�W�]iT>}hAq�_W�����ͫ|�q;���%���fycy�ۂgS�c�UX�b�t���
�䴊Q{YN��ys����!40a�bY�'(D#�������]�y
K�xpU��"~w���$�*S%8��q�|��������!z�ĳ��h�-��s��W����d^�|3ڍ���D�}�U��MX��
��|�~U(m�{�7�k�O������#�(����JZ:��⋷��iY�����s�0�_V���y�wF��ޱ����Ft����̦a)o�x����x7��3����t
�����C�n��e,�Ϻe�6M&8^K��(�ANh�K�s2��5T������uۥ������l
�c�2.T�#�}nC���E;M�O'��ȘN9�z�����s��a�QP3_���1&���ϯ�����rOC�g` ���=|�b�L�Kb���t5���N�p�ū!Į���L~�>�D��C���$�CP:HO��c��>j)��	�g������ߌ�X�{�oTU��%�,*�/5�dt��U�~6uyr�k�@����-��{�^�fD	�1��]��ן��"�+���8��gCY
I|�>Qޓ�e�s�{x�>�D�ڻ�ANH�uv>�U䙀`�<$Έ��rʭ�a����0���_�>��������&�kt]�<������qe� <z�&��P�f0b١����XbS׊�g�7��J���br�W�c��;J��r��]��I��г�ٟ��C�;?��	���ؼ�u��Ë���o�.����V)��m���xcC 3�A�檁0�2L��*�F6�~H��
O��� �(�!Z�#�?a9�܊�qN��+����ia��)�~(�Y���[k�o���O,;�s���p"�LUǪ3Mf�Ӆ��/v4D�C6�ާI���������ӆ�չ̼��W\#r��ѭҧ8U��_I�C*N�BH���<G���g���z ����V~"e)đ�Tm�c�2-����s��5�7�#�'����x{/���c�CrB��6)��e�w5��d<�yg�XA���P�$���0F/��<�^W}�۽����Pe+��;E�8%�}|�Jnd@�����`>�gA���ÔТgL���Y����v-s!a:_X����{���0}u|�]1�q�bp�Ik�����<��۾�cN2e�
N���,$rQ���Q��K/q�O\T�	��J�hx,�s�aas˸D�(�� ��{2=�0X�SLE�~WB1��Z�4�s���I��g�-��~��UA�YV�׸���^�i��'���;e���8x
�T�R�u����w�9tыZ�q�y�xtsV$ь0�O1���G6��v8$��d_�����dOOщH�N���nsV�wgW܅3k��Z3��^����v:X��#�����?y�kE��W�"�k���]�զ`]0��̡�8^���zU�qTa����u�zJ�ݰ��s{��=Y�{޺&�����1�9�����*h�L�>cvz\7���~NKԼ�T�ź��_=�E�fbv����خ��c��������R��gN�Z�q�.���/'!��U�Ϊ��z)Fc��b�W����WV=�J��7[���F�|����+������KT􍏨Z�mwr%���3�,�q'�`݌��>>>o7�����O7=Xy�/T8g~�"��y�]6C�T\8��i1���}Oz`z-���ɋ7.m�Y���~��Q�5��G&���ώ�Q�(9�[�Wz)���S�[�v?_o����C����L��>���3�<�H^<;�A��ht\O�XT*��/^�I�\=�m��M�Z���ެg(fհ��{J8���>����H|u�F}�d�?�X�.t�5;r��ǖ��ݷ���T.��dP�`�М���nA���[��k���v.}�f.E~��Z��i��Fȇ����;�%=[=�<#�C��d�[e�>�0��6�9%��0y�wu���I^P�x!�[Ȁ��1q�b��7���Mw�Pd��Z��9ˌfNfu�"w�'��衪Y��޺@/Q���f ǇHt���#�:�u��Xc&}D��B���3�qb�~�5z��\8��G�r��$:uŔ�$�O�_["n�^��<S	�cϛD�k.:i�>���nѧ^��n��x.�)ƁF�[\uȟvEê��˷�)�0Ç*��[�8�k���*���Ych�Y�fù�4��h�n�vV3�Tf���^A.�=tT�)I�M��O�;��� &n�����'qaa<!�ͼy���Z��O�iдC�	��wi�.v�F�9z���n\�����
;o	m����y�o7���n��u<^��"�o�g�č�i>��N�y�Q���8�s��p�g��;�����8*�iQ�81���	���3��H���!<�P�
a�^�2�	o<[��)�sH�R6��4�\I�d�'2�n�v�Y�A�?`��מ�B��g�):z�p��U�\�^�!4���Q��79|��y�02�-�멙�b���ĸ���f��#!�Q��}R��~�(���]J����[���K�[n�r�������ߪA��>��$P����[�y���D�7a���޹%U\_K��ޕ+��N)۠�cܒ�}��s����ʡom	��2H07H2�LY�Fj����t�[�SKuަw�0oZ�9��fh�����L<v/�_	�&]�tQ���X��ՕYH�Rj� ���Oy0X`K��P���ʇ|���'���/\�!hs�O��==*#l���5���u�g��@P�ba'�!鬹�����5�$��҈i�#��[ͭ��=�`5,�o�ܵK���o�d3>X����������& +},�~���P��1��]�����\s��D�)J�3x�Hei
W�.$`���+!;J�K���c�1��Z��K2N/sK�uݡ�����	�1�(��;]����f�9 �����xi��L�ۄ�D�ܽX��&��Q��7$���uh+ţ�Cv[}g���OB���z �@���-�,έy��#��j�������gx��)�`��1�~��j�Qˑ�N���Y�g�U�S�+5��u�}�e�8'��zE2SӚ�壭�x\�C��q��h���4�ξ+����;J���tk+u��kW�����{��b|�T����ZB>�,��)z��Y����ޡj�����Z��OlPp0J�6@�rݞFzi:ė�è��V�Ͱ�Шk�z��D��T�v���C��@�EāCu>��}l�Lps���Kt�/@�4Ua��Fk��ٷ�GLue�iם�_�`@A/N�z^=&:�0�o�h�G��p�/�J{���"�ױ!����9�+6 2B���y@��bC�!�"�t {aQ�_�N��:SP}��PՑp�Ğy�M�G�;�8����Sߒ��Yq�a>O�=��!��]�qʙsa}��������%u�pp<��̍��*�R�@k*,*�O1�U�g�鳥�QSC``p�;DC"�˜a,�L��#8�Fz՟9UYY�69�.+�J׿L[O��s	ju����F�#�w�������t �[�������߷v�{wx�Jx��oԓ�q�o+jUb��kk�u[}��ïlR���ͻQ�S*���>���_}Y�Ҡ찮MnV�tw��i�b�z�i��YT���R��N�K��k4�Ӫ��4�n�pU]�")�~�> �{�|,��v�GD���1�U]�H7`�lVeK�̧�G�I:��aw��o�ZG����}��]�Ѓ������H�m�"����v�EjO��
�6=+��"�k�'��Ak:�FwD�^�C�cл��5Z�t�ۚ��g�,���0-�t�.�������yN�!}*Y�1o� ��)�`�>��zJ'��8Ӱn�"]^@!��Â-�dJ�:��&>��\%� 9�P�#�b"��k��7�ۼ���Y�Y+^Z� ���HA����&�z��i1,N��;��Y�$p�E������u�p��g�І����puG.�Pd뇬ٶ�1P�7��ݨi�J��k��p8��`_Ւ�E�����'xBj�R"�P����B��x�t���T��ly�ձ'�<0lˎ"���	�x��Q�>�"u�z%:��1�j{�N.�%�Y-N�[��gob�ǘ�t^��ȧ�x���ȾT�I�w��
����a޹g�ȷY*�{�eM=�<�W�^��l��&���{�����s>N2���C��<h-��+%���;��)w��\���?2�'|ݗ��S��ڠ��d�m9��f���^���L�������@r.6=p<IĴ�<rޙi�\��p�i�2zbt�5I���:	��Q����<̂(y#m�AncT����0#0;��7�y���|=�{U�Ί�,8�"�Y�-~����;����(ps��<qx��H��^f�^�o�K������5��o��=q�O�`�,it�~�'�\>�h�)��]X�=뛫�η�p��d�!X���<�O���*~�L�Q�b�T;��{$sV��w��cH�;[ї�����Z ��t�0#�r���s��QT'1i7�k�A/r�J���P�kɏR��n���|چ�0��0h�"L3�������u���������z�7�oZ�fϝ���{�N�;�5�T���d�cȉ�=��S�!Pz.��K[����{��s0��3��4#�3B��7�~;�h�Z��W���#�@��]���f�|3m-���s����#ci����z��-��׭R������F�]�UYR���녵��`��iE_]��}��H^W�����9��q>�e�80���u�l�.���1��FpF(��@.Ɵ��};�#��+��:J1�1]�ǣ�zi�S;��lK�I���f�(b^�s��<��T�+��[��n�0һU�ڂ���n)�읔�#f�t�r��v�'L��+]v�(�pp��dM�,�QQ���A���|��n��[-l#]&���%<ҪT�%K�\�1	
b��FE�τ�{uu=�(8a�+]R+�⺷W�!�]m��%f`��w4:��S�Z���i�Ⳏ[����^'1�[��B78]��d��;��8�X�W����4y=0��m'��E�Q`�r�*�jV�9�H`F�5{�4Au�v�V�o��"�`�Nc�!���rܥ�CF��J� ����U���r�$=���Ry�^�VeV{D"�.:K{I��*��E�T�5)3�ꐒ��sc����9�NbQ��z�K�F]�r�.zq%�u��5qz�\=F��i��&��U��VV-�4�K�N�$�RVvL.q���݊������u�Ӷ��B�NA�"qeJ4$)��d�f|s�.z�*��"��9q{���oq=&�-	GSj��J5oeBڨF�L�����x��R��8j�4ޅPmݑ�n�]k��b�6�/J��5Q�t_
�(i4f`��uWL�P���*��v�61LܝJ����n�ÝWed�S�a���.��R���E���vx�v�1�Um\ڃ54Q������M컾e������f�|���o�+���5�K�l�y��5�~>�쯘���|�G��Y]�{��#�gU�UN��Z�HM�>���i���Dcr�MC;i�f�^&�c76��N�[�F��E�蕘z^�gf�N(B���݅���(+B��&QuI�:��k�l�~w(�Ř��zn:��z��Z�s:jS4t�0�zS� �����^B���0���_Y�y��wG=/�LUWZhƍ���kS�
;؉�Z��|�c �2�{�[��T�-n%G���W����v�z�=�Y���������l\4�X�Cy���t��X�Q��U��K�k�Lb��P(3�e<�UPIn��K j��j�5To9�oE���R����������]��I��m��.�u ���~�!���V��5�!m�n�r�8?$q�S���)*6R������U���a�8/2u���zZ}�H�rע���yo��i7-��b<1d\���qq��4o"3b/"�@��TKi������7�ؓj��m���Ykpj���z�b���}NV����>��T�a��!%3�]͸G���j�`�ݽ)���b�^"g��h�M`DV[��zr8D-���%?��A�6���m���m�$�Q����6]Y�����[Up��W��r��b�-�IR�9C\\Y\�4�,Ի���A�j��Ʌ8[H;�U���oV�2Vn�ZV"wv���2e\[�?����翝{���}BE�K	P)��)�d�R��q��#�5������x��Ǐ<z���،�(2�5��3L�F1(�1�1���0�{u�qǏ�x��Ǐ^��d�H�  (�d���I��Ƣ"��n�FF=m�qǏ=x��Ǐ^��J��1Il�ђ1F4h)(�d	I$� @�]8�8��ǯ7���{�~�����h3�`
4I�K���ƍ�t
M@$F��D,E!�PE}�BIc �:�0S��Б�E%3n�M\ܹ�H��C"�[��kQX�6M?��*ѹs���a#L�h-ˢ�F�$aQD��ܯ��"L��/�t�F�f2��O�F������>~yݚ�,�5M=Hiy����M
cI���[nq�4���y,u�F�w8���J�M��y����g�X�1�g�3���B�!�)��,�ѳ�)��j��C��=0'EϜ.>0�צ;�:f:�N�u��zbU��ʫ�>ʄ󦵅��9�c\xVK���h14C�2=�\��~���:9�:e�o|��T�qn��z��Y�nN��dU����q�����Ϩ�2P������c���V%.�d���z��8!qe��̋ߺ"K����L��,P����
��� TnO�a�P��k;+��4`��A��FuO�/e;�ޥI9wLR�F�U�9��Yz��QV���n2{wT��E��'"*6���������<cɹby�=~z0�Q(Tb�!�f�r������#����Y:0�\A�</H��z�
sGS�A��^��f</<c��{��ζ�nJ��L�jg}`*10kf�r�~=�H&����~���6Z-�39�����MM��ߙx93?)??g��T6�g�H=D4-!���y�;E�_[.����C���Z�k��d ��,6�n��X�zy�$���A|����L� �}�x�~W9W.�k���uMOOޓ��s�b��M�$��I�S�r����+�ꃬ4�ASz��ܪK-�w�JVWp/(��Gm�R�.���oRȣ'`��$42u-�rU(��LfY�:�rdtR����$�"FeQXD�������y�E)��ga�B&��y��o7����^�q&�2��Ӏ��9�!�<[� 0�g�'� s���EsϱŁ��>(D�&vk�|�,O�D���/�Ѯx���-�q����b���[�D�������\��EFݓmU��7�NIf	�5|��Q(x\�_L�'�2"�Ӝ�`�^��"w�a(�TC ��Mu?O�bv��\L���c��z����R��$M�X����M �ÿ,�~��*'�w@�=�fW\SUy�c+V�����>�w��@�ײ���aDK� C�Z(�%������}g�6Z%Z�Sq�����AxYX�Ӎ���o�M)��c�!��)����z�Ɋ%oc��3�)�^�-�OC�]��ʞ��+��.
�M;���5uE��([�=t�����k��ۛ�q]��yl)��`r��6!7s�C��N�����d���&��Q/nu]��b�d��4��O7�H{hN�z�K�FG0E�͕I�{�eI�s	]��:�q�	/Y�{�iu�xO��%��܉��"���9���`����1��N��L+���훠dKC�Y����7�.-^<ʠ�CB�\�{۬j��Sg�ս�tۂ�,���,�J2mE��j�����Qk�j����)1W:����*m�!�a���qGj�L۱m��)�ʹ�Ư]Yȴ+YV��:��f� �����~����i�)ҭW�畇��t���0��*��UWN�#�=�g�w��1FA��4�O>��^�Ѓ�h�~��K��̉�ŵ�%�Pn�L��&���E�R5�y�=��%��ל�38b�w��9ك{40���it���j��+9D?E����`\*�
�ڠ6<�r�(t3�5����9��Sg.i����F�+k�! �C�n���Ndӎ'�k�PK�o�Ds���R��s��2~��4�F���{�y���d�%=%�6=`q�L��ih<�CX���:���}���[�}���77񡴅2��0y��C3��<�@��q�*>�=Й�.Vr�6k���s
Nz�I�S�p���CO:L�DD��e�`���=>Q��Y�z?��L.�f<�=����8��}#S�%�4�z��"�%D�W �����B��u=�}.pK������(S�#;4���8�禷ݕ�id�+Ț�?�\�j2�0Ʌ��<��<��݆aҷ{�U����=5�r��ǚ�B�#q��ǎe�>�Ͱ�銗�<z�V�Z�F;hg�?//=�5T�Yu1)�Y�h��ث4����z&o*P��&�3��bm��e�F�/�X����"<b���^a��:�V�N�³�u�uN�z:�}p�'f��˃	��20����pi�ܶ�s�*�E�]]��N�խ������y��a�o��첚�y3?� ��+�1�MtY�C+� i�I!}Aq���	�yb��=�TvAț0a���EnX��g��_��L��e�����C�#\�Tx��)F69��ހ%:\:�@�Q�y���W-y@�����A�Jo��r�Q Hqm �/��BO��f���'vh�tѹx��" ��Fߐ׉nO`j�bQ�ü��(=�eL>�8�DPo�g������g����;wU�$�C�������D��G<S�#��1��ޚQ�aQ]q��94���a�"PVԦn���O\��|c���&���~e~.�L?2lil0q#GK�Γ�g*D̙����lП-0�AuR״M�*�=x_F�����r����ڜY��oW����exI��1��=;B�z��LKb��fW���yBײ���vov9�1�%>�����PW��Ls	�4A�o��l}0J��e)�C���;�`��ڸ�̟�y��>�zJ9��'*�k���|���}9�s3��>&����c�KJ��A!r�SH�n*�Y����Oj�R����=̱#krr�o�V�E���@�����)��0�c��xfTK7��ê�K�':I��9����F���`�Kwaj�LΗN7r�]ww�v�bu\���RY�шD��7��y�o7�A���O�rs�۳>�??C�Ux��ޯ^��a����`1�$`���X�c3B����7��3+-o�!z�����馟4���@2/�t|h(���*cn$����έ��B;��;/8�zv}C/P�ƟC��;��/	 ���P���~9�V��g��P͌�kim��3F;*��9s�uᗩ�,F4�Ň���y��>��T�; �t�c�p2"���nZks*��x����I��w~��ա�_VAI@�}p:N����E�F�r�ˈ��2ϯ��mv<�9���ޫ,�{��F�s�ٮ�+��U�W����"�l}ʇ\���w�Y.0 �����{̨��`��X����_��i���ΞE=��O�<�hz�otT�#@i�R������n��O��Bb^�"K�	H�%%57G\��p�Ӣv�u�	أc�<�ۺ��v
�2BDM[?{�0'r�	~������w��O��7��|�(о�\��g�iZ�6bx��Z��������aG�Ȏm�n�.��.�-��~/I�QO@�Gb�T4S��}؃6ܙ}�ZS6cw5Y�h��pʡ2��p��ujkj�������I;�B��:���
��Z��0m\��x:��M���W[���K�.惙s�J�a�.]5�j�►�}º�N�g�ʾ�ښ`F1�&w7�����y;�nߌ��P��f� _Z�9#���]
٣�<�{]�>�h�Ҫ���-aw1ٜ�y���t/!'M>ȁ���Y`�쑴�؃�}uB�'�J�9^�b�>e�IԺ�h��3rv(��ڠ`�d����*��N�;pC�!��aغ/�Y�xv�Pzj�n�w_diH���@7�;$|��=>���傦
�����'|f�<xD�cͥ]��Yg���=z]����8��㭏M0�qh�ƹ��A����!�V�%4Ò�2f�^�vH���F�5��a�3�`6��u�A3\�Cz#�r�un&�)���;Z�j�ݜ {Tu����'c��6�9�*wikN�dg�G�,К���G2����l�3Y<�:/��>t�[�qt��6V�x�{�p�j����w���\��莬����kܢA�{����F�A�FM2�/�c:z������2�P���1w�y����Ƶ��WuỒ�wٵ����4<�q5�a|�sn$\�C�qN���Q����ǰC��䋅�Ce�Asl���X.�8'U���Nhh3��]�F��9�a=x�0AuڛC-֖(:�Uv|��]N��c]]6vu7=]��S���Z�Ҳ�B
$��wP|Q"L_
f����KF*����gIJ,��[U[�^���=c�i��VWg���w<�w\������+m%��$�
�1�hv��3�Aś��>P�g�˯���|���+�I'��
c���'H��U���n��IK��G	M�[�t&��q�=P[�M���	��J��z UE8��k��y��_'x"z�[���7_S5��g��&v�E8�C�֨\�hl����k��*�ml#�;W)���!��_%^�=��v��r��$���9�L9���Ȭ�Ν��E�����w��& ��yD��ir�<ҷ�F�ٮv`��{򘶀�ڂ~��]7"���fN�ܟwc$M�(���^�'��Ԣ�=�/.5'���]���0t�,�S2��KΛU�զlR׮��������@�*l��8v�.XGk��q��P �#KI��������vs�Cb`������X��+P$���qC�+\�%鏥G0��:ݭx�K��9���Ѫ�oз�� !pc�_�`|`an)��t���z��=5���\��O��W���G\t.�!��^�9����A��0�<F\k�'���9x��'O;u���:N�HP�J�����S(��K���Y�tfIx�K��\2�]�p�T�ʍ���Wv�ﰌ�	ۨ�Җ�&V�*q�������T�D��I�e��z�qH̫�웵Wv(N�Z]��,�����$�ӵ*���]0������'�g�/|�0���
�)A�Uز_>Ǉc�D�:�z4�yw���D313]�jY�M,��]v����ߌz�@3O�zn5��.��ݰDxL �'JѬ�bm�g�r�G�,�]�%ח���q����1 o��Q'Q�ȫ�疣��Sؕ�DϛE�S��z�ֆ{u�E�[F�4��^!�q��K�H���'��,����5����Y�l3 q5,�.�.�k��Kd���ɏlQ��!��A���*ElP�Y�B�ϚD��0"*�^5��KN�B��j�vz]�p�I������u�.���@%@�!�Z�iN�ݱ�b�vY*D�j�����j޸@s���%�j
}��ߞK�Z���z���w�~�ʌ$���>f�ץ��ev�hU|��&{��sıOk��׊4�S�W8`.�渀\]z!0�c�w,�E��wsS�8�!�To!`�8y�I�S�\�LioP�1��p���L��|�18�nj=sg/ ��-�09�lȕWԝ����1i������a��'ս9.c%{d.��|w9k�D�ۦ�]Cj[e�|��M�aYX�quiJ�NV���5���\��p�&$ɝ{*�ڽ�S��B�����^��:9��͠���K�v�0CWp���L_C�U�X4��O�����e����g��=×��[��T��2�>gyń�U�`!ϼ��[a�	��p%�ǍT�l�dV�JԿ{���j�sߧ{W'2g��g�7�ָY��DRY�u��+#�#_�An��9���[���o)Z��ϖu�����O|����!� ����#�]�4u~0~��A����o�t����v��>m��-N��}�ɜ}N,r�,D�ШD>���������;���?[{����|�a�O�*7`?�/�V�5�O�sL���;C��{�4N�P�qdӎ���b'(��p����yG۾4*�HO``ӬN���l!�s�'���ꈿt���UYR���d4�>I��\r?8� A�l��r��DJ=0���p�����א���J6�LqO{{�NS`��$��Xqc��O{c�ȧk�F&�WP"|�y�e�zc�^�
�;��U�]�C*a�w�{�U~��9-�����]�{O�e�ADK`��˟��Y�׬��َ`JU9z:jU���ۥ�0dԲ$��u��x��ȼx/���t��h�Bdw���b�~�2��t8q��˶�O�O!�-�
9(�aۼ�3�(Q�H<��W���.�_�^r�/����>��󹻢ϑ�է�
u�צ���*�7�q'�Q�8���2J;GWmfk�ݙ�h-�F#0ҥ)�Ҕ��#
r����ާ�o2\�O�1���*F�P�_���yʬ�C�c[���bY')D�	OH��m�����x�~�����fn��\xݸ�r�w�B�Z�ވ�����E2 *4�����m��tT:�'�"��ľr̨�����1�1�^\.��2�;pcu���;�ԩ'.�\�(�U�9����$�ٯxVp�Yk���y�������Bm��ۂ�Ay�K���"��-?,� �L�)?gMݰ:��=���Ů��^@��	w�8~Zl5�� i�ڪs�j��
ܾ�ޥ�'u�t����<.��`=���c��&��!�dO����P5�����lB��]����2���'��� ��(F-z`��O�v�Ց�4{=!����}��y�k�ԯ^��R�b�r�|��+�$��%.���	zv�Dg�x��<���bq�8�M*Զ�n�I��]�^\����Yznݫ*=�Y����(�A�;*�d����8�@`��'4������񍹵;���%sj:�S�%ѷ�&��z3S�X�k�pm�M�>r]�m��ʙV�l�hV]ƕ^~oqilź��mЙ��+��ޮTގ9OKw�<s�Զk�ۇM�z��sN5L�3�m�<ʺ����f��D�ʛm����Fan�m�L�X��ޗ\�Zej�lPy�q�i1�o+;����"�C��D[^��.v�a\`1�J�$M	ʥ�j��m�P�N#x5*6�X�,��9��T�-��t�EY���Ys��dJ����]��e�U�&;�) ���;d���k"�e���[��]�kgf��+�x�Q����)�WY;�*z�a'�2g%&Bb��j�X�\f���D�٦T���b�l��%���M�c5��6�Ͱ],۳��%kֳ/v)1gv��
����Ap��f�9���J��Lfޠ�F��P��D���'����Vɶ�-캛d���� �X5�3{�x����V�n�Bmo�o�EYtبb�$���5e�C��wv8o���P�D�OA�n����<L"o��������!w]E�9Y3�ۮ�lc.�T�f���`��Lf��;�C5t��0�I)8;�w��X�m*����b'
�:��n<c3y�0��UVp��ԙ���G�&�n8ΜznP��Y�hr���V�+�q(�m�����)�[��u���ޡ��,�y�~WkA��/zu-rM�H��>�vr�M�*:]�r7��*S%&�&��rVCox��@�$bA�+<�\̩��MAY���5����ư1�Ё�^�LM8��bMyj�{<�-3�e^,Wc�����¯b-S��[ma���SwP;x�������vx]����<��U �T'{��Q��tΚҢ��j�Z����ֵыdK���Y���|��&oUj�\�����[C��1\�n�W)��V��j,�p%V9$T$��婹̼�M��s�����3&��4�=ԥ�vz��xѓ�U����h��e_*v��E�pܻ(�5��WM�J�AڳJ���ѐ��;6��� t�����j�a1�.2�T�X\YSe�C�7��q�Y/�S�WR:n��j�ɕ���S].뫋�������8�O���z��X;�6�'�v�t�Yׇ4(�v��Okmc�N2��ٍո�j���"IV`�opv�9gVSC(	�sf��X)��:gvST���"��t�{����h���G���_;F��!u)Jǵ��^-���\�F�^����Xӗ�r�B�㳩��b#]�ԕ����|�A,��ݹZ��:LJt�f��'��mܪZ^�[�Ů��������3)����y��zJ05�?��*�춳��ӫ�����@WR�* �XB�u1��ZC{z#w(*��6�ݭn�<��B1V*�&r$Ur+*w*&�u��[5��"�)k��ߟ�|��"��}7,B�ͮR2�v1�QH0%QQ�8����Ǐ;~�<x�~����Y&�RHwr�Д�F�$�*O�ڐd���$��$H���8�Ǐ;z��Ǐ^��$IBE�d��_�ҊJ"��_�� H�BHƛm�q�ǎ޼x����w����Y,��77I(�۱�ͮ���B��m��<x��׏<z���j"���ܻ��"�F1�%~�Z7ۛ��K$$,�E��ȂW�u��=܂(��Re4D1�aL� ��Sy�;WLowRd,k���HF��)7w+�_��*/wD@��d��(���1+��"s�I!�;_^�ʐ�)��H{��E;�\�C�ع�2K&�-��QmH���Ѣ�H�@�|�$�ZH�V^�S�?%y�lk��˙ݧ4�0�c�2t�&�����#�f.��z:��)���V�89�y�Ӆ�@��`p�*D�D��(�cjU
0*I4�J�����p�$.3e&�Ix� Ҍ��(��ƙ���-��h�l������������#4~��>�_�g�z���29$�D�W\���w����ð�DO���[����no����`T��W���3u�5�mK���rx���x <[�\�O!��n�[w�sP�HnG�5䰉�W�&�ڷS��`��eu^Jn��ˉ6{;��c�$ ���169�W���RJ�c�¢\���1�|�S�MK���>}�ۄ'1R*&f��{�z�t��ڪ�����Y�^3����`��.�����suq�����I��Q�4V�c��s�TH��u��-��D�9���{וR|�J|r߻3�0�,�,��w����DWcŴ�Ջ����Kq�%K��������>�V�ё�Ӳ���\%t ��FR,fɜ*$S�&�l��p�/x�d8~���9���FB�}����4���w�0i�ɩ�7�̮����j���^�H���yԅ��\]�~�A�sք�>������.A�V��U��u���+d�4��k���ݒ�nP�%n#G"Z�u�*����yʹ����S(�p1Yqu7��:�AKN�X�n��ͷ�z�֋���3�e��r���U��ps����5�{}]��	:oi���{����^>>w��v���bŕB��-=�#K���5[�9Z��n��-ʶ�e6$��{ws����GO�C�*b�Ȳ�M/�t�{�_�s��yvҹi���˛��h�O���r2�q�B���'�@yM������:�6��Wګ���j�?�*�Ǆ��[����{�G��V�I�I�
����_j�7�H��sǰ?i�8�>�fg�*�݊7���ҝ]��y�'D�t�y� �Ex�}�:*9��o��0��랳�,ܺ��6AO�)[=��I�O6m�h��4��R:)��&+T��]p�`?P7>w魷�.�{��e���_3٫�I�-m�"�ܝ� �#����/��}�O���t�s�F{7��7���k�7,,ݭX��Kěں7=��l��f�O��؃k"�;�#�ȁKq�{R���	��m={����F╘��)�/9D�g��77��Θ��.Uy}�t*��ʂ���V��u�Rb����M�hL���u6��7x�d�Av�3e85�EN�Z���;���o4^���q�Y���sa{3�}��h��Q�1�Z��������5��4�3�:0���AS�ן� u���hu�H��é��ɠCD��Ǌ㗠�(� r6�4�H��P~���~�T7~����c�n��J�F�<��o�B�.�;��M���r�R�<�f����Y����M��\K�����eR3�m`�������dW&�\u�oR�`���qsmx�A)� �Q���n���/u�j8^{1��k1Oݭ�/��qE�R��E��kn��2�O[Y��Rs�S��=�"���G�ت?]P���-�q�9²L�<N%��I����7S^��o�=��pr8.� ���L.�����0ˉqgAן�s���� Ϗ��5�`�ӛj[�K������&�����x�
���7kHck�����l�-����jJ���S�z�y�o��@?J���b�V�w[��榃#9������?eј��ʨRw<њQ'J,1`�f^���!����xX���@�q���j�X�"��%5t$��,�k����t��Yx��`��:�PI�7��U�6�����u�3��5k�7t�
ɡ"�"�*�q���9RW����M1�P�U9��|�����x��/�K�b,���g�*�E��y{�*z�ܔ��_:���Q�=O3�M��r�9��!TM�GSzh-I�6W�)�}�&6��y7܎o�A8U��}N�����sxx`Q.��y	�ɒ͌�ol�����-&�����[�q�U�ח�� �E��樺�=9r21�z�n�v�9�i���PS�qz�F�c��d�Zh�Z�e�wn(��1�?+�B�/����ʉTh����	V_kG�ꮾ������G'�qp�u�z�r��y���Y``ͥy2����r`;���-g�fZ+���y�+�7*oAO��U�U���եأ�=�`�o���s۫v����D���}~nF���ᮦ{*vq{С�RMlOCwwy)-ћ�o����`����x.���Y�/}?>*���s��fF��1*�d��j�c�{��k���Ņ�m@��jv�g2VΑ#2n\Lͷ�l���5H��u��U����<���2�2��>�����%۝�����WtQ�cd9q;s��d&��e��?/��o|�7��������A�c��ޛ�ᱷ{�8���� �&^m��6��������'7�yP��b���*�$mD��
b�#�p�������8���@��Y���ۊ���[��Vq�T����PnQ{�tO�m���k8��= �g���Q���%��W��=Sj�75�ս{-<v`ԆX��sπ8��5uO�f��{��_��3i�s{��i�s.���;���o�w
S���tF�r��3@��֎�3���A��w����:ڮצ|I��]-zrw|����ס���~S�ѭ4�<Ցk�����8m��JȒ�U��N��X.E4���Wf�ɱZ|���/���;���r���{X��D�{�wFE�K���$�����Fp>C���W��}���ɯ��ֶqMv�U����Z̛���y���Qo:n{�-�sg;w6'�My)�*k�#�I���/��	Ԝ�l�e�ތ�#��Y�0�C����y2Ŕ�RQ�I^AE�����*bF��6��c�%�9`�ѕ9�MM�U"�Y�v�U��fPyFB���oK�YuZ P�Sb�ǵs�:�����o7������U�����f\?�7k���w,?H��@$�D���@�WT���W�C�O^�={}ZF:���d��������1�8�[�T�7��;x�r���f���B�ui���][ϲv{�"�7�]�ѭ� �׵�������-^i��rR�/�<ѤJ�sq�u*�Y�	�q��"�+���wB�����z��T7�*�q�������6��K�B���wsuI��0�>^�f˲;U�M܈ӫ7�8�k6�������£��֗R&o�n�〽x}�N���]u��K��Lj[����|y˞��swӢ��Np�;�g�]�1�|�h��VTE��(�f#�ӽAy�'�H��[�G���_�t�nxp·>�#L]yM"�74�ee�y�(`ʺzK}��>qC��
n]�7�>�J�o)Z��>ͩY��R�,55����Ĺ��s�G���݌���qDN%F`;J*���ӊ��	�j)�#P��"q��jc����f���x(�鍽p�l�oq9�F.�ީ�G'l��rS�z�0J�'�ժv�`���N[�,�Œ��gJ;U������{�������忶�OQmO�������n5}�L�����՞��~1pԅѫ:<�oћ��P���0s�ڡ�v%�`��AW釹 T?D��j��$]�4���6�VS��'"w�*��R�\�6@PF��>VR.^�*�bԹ�&=g�o9� ���B��Ԭ�c�N��M9�kN�+&�ɏL0��y�S����y��D����RH���$#�G���޲{\D�";�kz�z����.�f��[=Ǌ���r}��� ��
���y�ŕ[`S��{��Y�6.��k9��3�I�R�n��p�6��1x��o��pܘղ/��O��4g~2��(�s�t��m�[�	gΈf~�ʠ�t;����~�Uzlޣ\Qy
s&�t`�1����/��\Փ&���|�oC�z�1H�S���}EU�Y܁|��Kz��1xu�q�k�vWt8%*���t�J��е�eY�!)7ZF/h����;J��ڊ����X��N&�qI;fPW�bx]M�6�s�o:�b���f��'7��=�Q�s9�7`@����ueP5׏*�*��~��c�w^y~�;<�;�Ü~���D�W�{�e-��clà�,5�����fD4�ݭ�:nF��Ez�t��گL�������Yͣ�����\�=or��Ȩȩ�$�կ�R<�.-_rP��NߓTж��&���G¾Yq�x[*���c��xb����Z���T0e�{����.�a���)�߉|�2Y�'`rY�=C@"����X�ɫ�`��*��W{У�5��hۯk4;ٽU��^]��[��'��<�����
�}"m��-�M�-W=Y5�Q4"#�� l�f4{=�������1#h��4H�/�+���%�xzfN��opWZPR�Hw%1���ǹ��X�æg�б�q�]�ѿg�ʃ��A��`/8�JUx�L���m��qYJtdev6�q� ]_v�ct�p�S���+�ˣ�5����*W��v*"rZ�&�<�UCV'�4Y��cʗH�Ckr��`�w�j��iw�Tz��h��X�ʶg���|��]3TD�Ⳝ��:��b��ӳKjq5Q���Azr�qj�Fc�{g�>�����������4��˴_e��H�v^���x�������Q�b���u�nڲ��o�hNSѴ؃W�����⣑��I7�������_�u�J��Ճs��#yz�-�%/�Cq�:/�vG=��/�}C7h��W��32��sdk��[1���nkSE4PJS+[/KI�;���<�g{�`}��n���>n����|F�D*��M��j�%ma}9�{������/z�Ud�ȮH�wG�.ǃ>��i��c�y[��hd-l�}ܽޭSRjfZCCC�z@�:ݪw�@R�肔���l��+|�j�c�G�.�0�pM,S���߫�O�O��v��=�PvN?u�FI�)	5Y��Ϙ_��X�@Yn+R��vɡŻ ���׃�B�8�w��8�c�LR��IH���d��s-^m�r�/fA{��g�^E�}�0���5�c{%)����Mw��h�\��<xë���~�ԅ^�Nox�Q�0����b�h�}(Y9�7?(�.JFxhOWz����
f�͛���̹�n���b܈Q�Ζ�೗s��4�P�\��݃�8K�i�@?om�����`�2��Q��u]���ْ!����z�ްsxb�پ����1KY�u�M�<V57K*2A[��9+DL�y��o7���ڽ4NV4Ũ�3T�V�w8.	Y
��T�Q�F�w��%$_gm���ٗ�ޣ���֎�t�G[L�i�pz�#k� 6������1��M��ì�i�=�������m�SQٖ���M�)J�y> M<Oz� .Nm��\U� P	�Ғ{=��|o�_�'�K��\�é�F������>!��k�A
+xvD��[��Q��w�M����E+n�W���NdfO�C���Y�"hnԾƤIx���4�3�܀��m��FRjH���F|������a�k�Brv��i�;�?��2� 
�ѳZ�_y2���f�(l'{�޷�xz��I�/���c.���K��ۗ{ȫ��V��Y�z�"0���5���[�94EKj`�ny��zc�M�M������~��<�����qc�����B*+oT��ۣi�����B�RK״�[n��;����̼�V���hN�*���ż��8هLZ`�`�J�w�*b+˘
���= �T��y>TvJ�R�3#^g{").����|����*���|;d�u��kt�yF'���w�w���SMݺ}x�WmۂUvr�+�Ҷ��b��HQ�7g^�lJ�6�n&�6�Bue۱:�Sf^��f���i�����α��.G����6��Ƥ����&��Yi��b��lC �sWOq$��_'��6���꤅�����•W;b��̳�m��N�rٖ��͒�l[�����r.|k+�w`K��g��.�Pn��e��U�p�,��,�bf��U����e�庄�(屻{�~D���v0ݞ.�N��$U�8F�oj�L���4���]�suP�<�l�L7wPR�Sd��30�;�m�jU��VS���)�]+�\��v��'!�W���-[����i��#�Po�*��$��
*V�GVŠe`od^�e:�b���W:�k:�,���xM��,Ģڸ�������⭓(�:����u�Os�C �\���֊�빗ч��2p�X�R!٫ �S��۩R[b6az-�7e���V';���EH�2��F+�K���w�!��$��:r��nY���Pkd͉�ε*w�*��ޔ�Ѹ���I4�o\���XFrP*��3�
�	j7��jŒ�	����ی ���^,%��ﾵ6�M��A8���U�ȉA-T�O�m�_�
��2�vܒ؝�n�;2-�ë.nˬT�n0u�ս��m1�bo�0�z���5@Ý�YP:�и�g�'//���,��ACMd�����;͚Y�ob��[�tu��G�5�%l0�Ӯ��Mn�e'/��9�6�$���AaOj�[�'�Qm���{�ݺ��c��i�&ԍͭ�n�B�8�o]bF���pZj��Gl	w\�Iybs��6k�uP�0����-��,^��O�oE`e�ث��aTj.[��5@�k�1}[k1�BZ���+��7�ή���KO9�;T����%��ME@T��1-0�:�:�
�:��Q��GM���űP��t�[{�aP7�T�9�Y[*���I1�C��6�m���,���U�Y
R�(0d��%Ïa�t��rJ��ܩ�vjB˂<�'WU�i���X#�UeTB�:�*�+��i�1�u!:�3* lJ����'u)wVM�2�[ˌ�fv�2k^�f�P����V��lҰ����xT�G`K�Y
w4�a�o%ۍ����8*�mS�ܶx@��|��Omū�'L�IM[�&V�=@�x0w�R�f�e����k��(�UW�N�):��ʌ�l���Vs�<�q-� ؉z�!з��4���bh��V!�w��@�-_��%$i����Q4K6�!rM����^<x�Ǐ<z���Fȑ�$~���T���F%�ur�G�v��ێ8�Ǐ=x��ǯ\:�"��hM�#��r��˘�4d"��߯$������qǏ<v��Ǐ^��$$�w�`�16���܂#��W�b�Ww\�H�)6���q�Ǐ=x��ׯ{�ݶ�ؿV����=�˻�Cck���1����3)��^�w���h�_��()(�lY����wp��!��TH�W.�r5�wm�I�vQsn\����o#�+&5�\��[<�1�ۥ��d�)+��s�mʍ��b��E�%˖"w]�w|�<���9�vu����>�-����N�N*TuwR�l�uco%-G"�^5��"�Sj��)O+R�s7%��*f��5����X�1�b�Β�F��5��t�	j���s���c�=Ӿm���������q�oʹ"�xz�in���gN�<�|``|��3���y�Ϡ��]}Ec2�5k2���ğGn��Y�_\�,O��c��)�*�A��1O�!�/-i�V&�;�OUݹ�fqWO��Iǚ9�ut���l����#����(#G��7=�1�Z葶j|��O�������g�(mf"̱��9{�)�h�$�>d�}�2�����LO�j��uݳ��SۚXϝ�sQ�(�*��y�:U� ^x�G�^
~�l8qf��7�e��ʖ.�+TutՊ�u>�gYnJ7Ҕ(�#"7sK�ѝ��j�qY��8]-$�AIUO�y��e�huSxy�Vӛ*M�V���:#ӊ�&�<Al��0���C]:<���c=sO�<������2���gF���%DNn�E밳9f5�PyG�;-���U��v��rfmuRXӾ�B}�
Š�΍���i��M�#mv3�N1�m�כZ���t�Y���5�VU�֋�����bz��E���d����������K�3���X���)���<�_�v�T��wv��wf)�a^���M��]�*����s���.�A��0W&��#z���ۅ�ǊKEB��g}w��M�ϋȼ���j����ùR#�oQ�.��֪�2��N�˝޷5�^|N�k�M3��W�o0[�"1	�U��m��r$��-�9|mo��=�Q3)���R�|��#�O�<��EgfVnEJB���[��Bh	�b�V߯��>ɣ=9�RO�ֻ0�s� �XϯO�.G��.F��-�\=�����P��<�꙱Xk/St�^0��
Ax6_=�vqOܟT������G�n��k��識�.�J���L�I��]א��LMrw��ۘ�y�3�Yuɭ��;u�tVz+=�9�(UA���-��𜙦���5ub��/(������_q˕$�4y�*�u�)��PЋVܨv8f	����Z)Y�n+Kf�ۓ�7T��Ŕ������kI�ժ���,Kӊ��ͽ�2�6L�f��ڑ�	�*��(�>>>>>>�|��}:�ԝR?BMT�ݲ�r7���Z���(�<�C�[X���9���5)���g�n��@�h�GZsiH�e-@׭�6����=/PlN�]f3Cy��"�r
�LyALt��v�ח�C�?,��7�u���>'����_&ٍ�3��)J�=3㴽�+y�L��лy��N�eZה;Y�s�L#�ѝ��r�կ��G�Q/ c �Uft���c;�fYpܹ+c�͡	o�E]���S�O��������0�ˮ�YT}o'{Wq�#���sAd�B�}6=N_��4�yT�UZOK=�c6���K=�=���968ۿ7�g�g�	��]%Ui�#2e.����T����A�^�:3��>E``�4��N6FCf�N4K:Z�w7��\�0ku�#4��7���}ު�*E,͕^�So&A�a��~�ۺO���ؐ��YStaX}Ӵ�e��D����3}�$�
���o9�^��Z�3�v������:��Y�����5̴�NW�0]T�=�o*�1#n֢���:�H��֮%�<�ݷr��S�&j걄񍥮e��Y�.\��0�,���Ufk,윌O^����/Y|ԛ~1�c�s}�ﻭֳ�2g~o��}����,�)��� M0+�7ҵ�^���y_2�)������F{��/���@�g����W�"�T0b��F�%l��8�.C��_t?�?�������t9�Fc9P�c\���h��/�F��7u߰����99Y��nO��G8d(�A��2�����I?iꊹ������ϒ�3�«�U�[�ߩ�2׶��2]����n��K�)��
 =T��v����Ydv�q£~(�=��$?r�[b��,A�a}�
�Ϻ$!6X���#"��/OQ��-��;��p�LW�)�9���t6�M"�����+�%\�
6��ӢbadۿK���ڙ7��[>�IF8�=���G�V���0l��U��>�M#6�]U�ߛe^.Տ�1��k�@J�t�+����jQ껎�۷u=qSo�m9��K�ʥ��[�O� :�B��C:�JB�&<��U��qʄN�]���&�ܛ�:�3T�:��rS[.h����S<,M^��2f��z��&��S�/nS��5쳰
�U�[h��OQ��,k���S�
��q��{�9;*� g�x������i�^�^�V�)�0D7�c$�t���Ko��4����o>�������;���^Wv��#B���T�]�1�t�P�<�F�+����ɷ�%�����n1�l��ݒ��P�)�{���≫]�4(���E�H�2�X#w���5���f��_��F`�Z�3�[,L���sN�k��P��;e7}m��X
�,��0�!���8�p���ld6�U���o�*�p+�mx�����u?�|��Hr�;U-���'�v��ʀ®���8�%CzL��p!��)��yLnө{����ַ�bݐW� ��_/�4?��9�:[ }���68%L�w��.��0kA'*2�#�3�؟K���|I⣮��ɉۯ]|2����S[���$��L��s�Ϩl���BR!��1�U��/C]�I*6Td��Ʋ���vS
��!<�UwVW�V��d��(��nΊ���s�ܺ�/3�t]\�+&`��pB��ގu�[۰��u���7�wer�\^:��̭v�>\�gB���Dh�N;)iFgt6i�^Ʌt�M��)�R^��������ޗ}̯���W&�՛���>�j�(�e!ޑ^���E�L��0��w%6��֞^������-k����W��S�*��6���!��x×˟3���+2>�Zk�ʉ)(*u��}��&���ɗ�����9یF�(Ghfe7$@���ls�Kc�q^(�,�3�l2wЄΨ�����[�������C�^o49Y F�<���lr[�T*�䇖��+9�`M^n����8��)�x#���ſ��bO�S{g��o����k�5U���X����������	ԥq~�f�6�[ ���ф�����C]�u�S2}h�����-�0Ϛ�w���Mo _t4}x2ڽ���z�0;���v��:�;���/�9�LG6�-䳏t�����͛���;=14'�臌�y�*M��#_�(=����+��k�|ky��R�B���\�_�n�X;r��!M�s��r+�''��;$�!ϞO��=�wj�T�a��j��2:	=�v���QԄ'm�[�h�"=&���ᄊAd�$��9�t��Dɖ������[J;���\�y��5��tC���β��ҫ��]8�Ye�ڝX0G�ޏG����y�SҚy�ndƩ7i'P]�Konh�Kd����!�iy���zI ��ޤ$���!�ǟ�2ɳ~|�G���;��ۭ��B�ܸ���uI����>���^���b�,��ťb�g�Ef��m0vVGX��f���_���A��Y�+H��DS����C�`9)TUɠ.)�^6�̇CV$~��h�������wg��m��Y,�Ϭl�p�@jg�2�N��֭X$w!�:yeY
I�h���+.�F�8�l;t����f_Jû2o�������k�Tt��+��q�T^M�9�5���Ck����7��V���
��!fk=�:�:I��ʒ����m�ƭۋ�k~��I��M]�J��*�H.�}�G�C���s�4�q�Ȯ�W���s�cd���G	���uޅ���:L8(�Y|��>�WmW6�MWݫ^-��)�a����	��ֆf�(-�������=Jw��caL�����EuVu��-9Y�oW#��n�F�Hb*z9m���OE�{�6��֍����-C9�6q�܉���/!˷�rEF�����lt�d6�dK�ׅm<ڜіԬ�YצU&E��ĶZ�����繢��m��1�c���9ޚ���x��\�Ex��@���p��<�-�v�߯Of��E�.��
�wF�j��^k�1EwH]����[�v�[�t�p�m�%�ȭwf���}ݘ�3
v_w�����[�1Q�S��,u[b9e�I��>�_�J�2Y`�	�3��\�k�>o2(�%3i���n2>�E��sֽa���7;`Eyt�j/~d�J�yn?��p�к���/3ݝ�_2�K<|i�ߤA�7��O>�Lゟ@
M�Ē��i1�W�Z���\ͼ�;0�s��k>Y�	�޷x瀇F���=�Ũ�����6�$�v��yϫ���<#��Mѣӎhpy�Yr��n�Wq���p��vSߩ�Ǫ�u����* ��f�ֺ���ĳ+o�uR\�P�=��b�@CۿW��J]}ڤQ$���C���n48���}8�ظ���%�b���.m�!�q��Ոc�����Xp+�sU�q�|[0Q��
�T*�ePau�k��o[���^�#|��3�����g�b;�æS��<�.��Ҫ�a�P�-�ݷ}j��vp�᷇��*ɯ~��������ٹ�n��$���p*%�S_p,A�~�HϯA�zSub�<��{^�7;&�Ө
����x�Sy�Р��P(�)7-�㷝�5W������ͺ<l�j�*xŚk��N�� 	�%e�m���4��b�{x�^�㖽�E�toD�z�R��%q��;!���Xz/�E�m.�f�{��>Sh��KV���}EP����FVǺ4�q��zݛ�����b�S�X_�;�Q~�Fz���F��h�֛}���gC`�bs����d6��fw�D�M��[��o;�,��<���v3$IyO������0D�R�CO��8#6�04�&�Y�Z��OB�w<�Z���Ƕ�wR�J屷��7�9���1o\��݂�2C{�B�{��<�磝��SG��u��}th�r���`�3�����+��4��B�o�TF�'\[�gr�uLT�нo�07sm�ue0�7�RM��	�@���>�x�)�t�i1���r�GtC��ΣԨr��4v�!��sR�*:�\�9�ZVݒ9���E;w;�4.��I��>o0��{z�t��E��p��q+Ӆޓś�\{�GH�noU��܄-��X����,�Ե��0U�����up|�?�F���'D�A1	ϔ �7*�3�G��ԕ����qVz&�zO�#l��^io9�uk48f����s}�u	�!�j�X��.��2�:�|��8�e��8�0�o�0��dw÷]��1zs��{}�����a�;���r�ؐ�]�v��*̭Ӭ3k��w<���U)�>>n�^ܭ���:�&=�";<������0�TG�=�k{w�h�m��"U�e��3�ߕ�-�AS��s�ȷE�o=������OK�����+�#cr}�w}�k��D�9K#Hx��}���)��fz�����Ck�}�-�G
�O����3g��(�Ъ���д���F=ћ���P�-�:&�Y��&Xr��Qq��85!wI:�<m���f�7X�@��!�έ�U;4Br@���w�V��v9`���'bk�јN����t�ۭ���?u��O:�^�*�Y�1&ګ��b��]�9/��y����Q<b�:��ݐ�2�(��s+`���B��d���Kb��f���w���%y+
�tu�Dc;���n�!0��ڷz�g��d䍶n��!�Q�ba�̲);
�ʮ�������}��ʂ[Q�W(�ѽT���w�}Gkf8h"N�P�f�n�����aeUx�?#ϱ�0�\���8:�Q>WWx�`��A�K*�Ug4β����l��ݥ����*^mZ��a���#Tu�kk���lV�f!ivv':�3uj0Q\p],�����%Ȟ�V��-7Ocyx�p�a+p<�NJ��A�38��� �*:ծ��M��$�Z��5��˕[
ݖ�[�1��`�a���m�Uөn�Hh�9��(�qPL�l<ڣ.�бs��QnΧguS��F5�MfR��[�k�r�u:�j�(a۲��J��X����5���6sp;[4��Ep�w�OS����zE�ǘ�+"��}�MǗ`��[f������\��ruur�k�vD�N�]LΊ��<���z�9��\���rk���W��ܤ��#�f��O&l����CQ�YG������4��yX��:�x���D	�_|����3��\*'F��᳭[-�Ξ���ռc����w9�Y�J�C��;���$�ث�Erm�����	+�������J��+
@�t:��;V;��n�1F�Uc�ժI�u[�^�Q����A�c���]�~�Q�A��LS�f��5�|��4A[{�J�.�Tl��� r�ʣIK	��01��!hj��sfv���&m�b�e=iU
u��v��
ѧ01n�����\f4'!j�Dn��u�u���lʳI%rk�H�)��ٹK,<˝nv�� ���]z	�sS�}�����r�$[t���뱉�0U��p����Νӻ�24U[IBw�*��+�זN�)���^�R�ʅu;�iS�1Y�pT��Q^,�1=�W��Wn��U��[~[���bw��ٚ�����h�:��b�%m�v]���7�5U`��U�@��9fK�2$(Q+T+�f�^Bk4dg�n�����d:$B��=�6-�*�d���ٲ3y1+ݾ�F����2�����RzOU'Bjt$7�2��-2{l�$1�8�r�`�ҩF�����7�l��9ګ3��XQݷ�6a,�x/aX7�(P�d�1�%�J�B*e�8:r2�׈M�D⹤�3�Ov�����fMW��pe�c;�]-b��3ٕ�p�a��պ�輶����G]`v�73��]�@ȇI�8�ݵ�R��h�j���xx]N��ȹ��Ǩ�F#�
k��o5��9�ۖ��k�CP��o�>=z�۷n߳�oǯZs�����{���0�ۦ77f(�wr7 �Z�솋��m6���v�۷o]�z���āH ?^^Y�]ӱwv��+IR�#U暉&����eSM�z��ݻv��n=z�$$�HTdB��2w���4r�;�F�Q$�-F=z����v�۷�޽z���#�F�	*�FIUPh���v�uή��ۻww\ϝ�߾�7�%˗.gvwg\n�g�����F��c>u��{��v��苄�I۵�ůwE�|��U��u˜����\���N�`�_]�]�;�÷wL!�]#wq�w��G9q�c��]㳮t�+���.�:n��N���˝�y��]���u=�E�e�r��lk���r� Sm���)$�~���E���@�D�ԍ#q?Cp$������fV���]f�����qyè��KvX�j�X��=�ZY1\�!�qn����F���m�A�\&��	�1�QH�D1$a#��M��J$J>dD�b�Q�ZG��	y�|X�1#�H%D���D���>>>>>>�s�����+?E�1��l��w�&���&b�R�`�n)�|��fv���Y��pI�3�c6��`���{�ԥT$β��76tOw6@3��R�y� ��-�ط�0��qG�`w��[��`H��zb1�
�䶊&��)��_�z�{�s*Z�;�`�
��hV�`8%8˕|��Cn+��"��>�{�qIpL%��`�H�6f`;>��L��·&�7�\Qk�X�כ��T:[nz͊�ċ��6f�� ��<d5c��vm�_s��Žmt,���Ur�ROD��"�� �n�
�E>���aC���~)<�oZ�U�W4���}��gp�/m�i��\�H�1"�����pv�|`�_�.�u|�g�뫅Q{d�3�u�4Tc��T���
A6���l���:�gw��V�j���=ti�pί=�PV�]��_b	[�{��׀�	O���|5�YW��]P�R9��Øi�ܻ���>����.ֲLJGx���;|�7%�T��KM5����Q��(�%d�$�/Un�弋	޻�*�e�gb�{�4�����5��!�)�A���s���{�wR��
�~��y��o7���8�7w�:���!\�F;V��7����JTcWJ9�M��{������a�3�g�p�'5"�Y�S�/����J~hd�{�����fJ�iឮT�QT�-��S���:P��]Z�9Ć�K0�o3�n7w[�������=G@l�ۯ ����5�������94��q}�5�X��2���AR�`3_�p�/��2��a�^Tڢ��I�:�e�O^��!GH�35�^�#Wt����� ���^��W��'&=�Z�ك.�`zI��>5��4���U��b�1BVޢ_����7z�I��7M�#���8H�z����;�M���5�A40�E��J����]}
�(3f��B�%�$W�OÝ	{�g��~��#>�ؿ��n�̶q-������͆z�!�{W��Ag��vu]�Z�ECG2��c��qe�&̆��;ESw�10ݥ:�PHظ��Y��rغ�$ms2ڌ���)c&��=9[(�k ���b��9W�j��Kn�Q��ғBKn��(��N�6�mF�UKv���
�Q�|�2359�����9&ߌc�<v�o��OS��_]~Mzc�>�E�i��!�Ej�cS�<y���6C��EnR�U�D�4�" ׁ�-WE���q�[*�vN�fn��82 H)��^j0
�h�{5���+���SFR"��Dc����<��A�ń�j��=sK�M�5�B��;K=^U��� �=fOTTK���+�Y�U_����
\��ݗyj�Y��j�H��E��*X�PS�Tv�GM<�R���!#��s���՚���Ws:\RE���HܷS��h�g�;�TӁ��c����WIxG�HI�!?�X�%+c#��3����J=����y\���T�u��G���Ic�/Z򅗼�+�U R���)���ő�.�ȶNY����=g���
�:E#f����FQ�9b�B6>\�w8������U�S������v�%
CY<��6~�����~\/ֻ��a�p�/$V^��\B�["�Ç|U��~�Y���Wx�R���k�tw��n�Ka����tP��+A�ԍ�����/���W]��㋃X:R�˂�X��[m4����>�.L�mJ��u �?c`>�u��淪 �=u�i=�$w=E���㶙s�֕���w��:Y����8�ᅢ�5��c{���J8c�T����]�Ío�	�|]����=t���9�q?�jafOY;w� U�	����z���i�����QԥPm�j�����d��g~���I�^T�)-��'kzO���<Ȧ��	����p�����������X�Y��lЊ��0dU����t�I
7K�OX�T�V���z�=��g�z���Lȳy�%P}^𼳹��wg�T��s���+&�a�On/R���|�
�[6wJ�&D���������Z��ȁ���j3[�����/�y�ͯ��5�j7�F8%�;���uos�RM^c�f'+x���g�X�PS�vj�MCPL�32c'�6�T�W�1��֍�s�`ki�-S�2B�v��1c}�L�PYچz��$m�S�7SYf�r_,�EJ�>�Uw]���4�f�޷��k���-EUĲ]�ҍ����+u�{IEB��^�̪T�1x�fp�Ƥ+f�dz�L�>>>>>>߳���S6au�Oo/!1�Y�D^�f�㿙�or[��?b�;/�Y�1���KA%*RU6�Y5�ܽ���Kt�c>[8T�=��Xo��[(�g+��Qʊ���`2/=ja�2� �/��P�����ar�+�Fl�Q�R�_X��'u�ѻ۩�1�������EG�C���Z��:)��`J��WD�&���<]w<�Q�%8%t��d�m���!�b�����d�f�ka�<Ѽ��d.�����qJ�[�?��Y\e����օM�|��xI�ub�2y���t�D&����V�(�����)n����1ڮ��fY��fA��r�6\�I�>���W[��>p�k���o姹��K�m1x"{�X��=��]�E�+��(��-�)��Q�o���(��9�����A @����f�SX��u�!�[*DL�n숓�Q�e'�Dd��ޗ���n��LJ����w�!$ o,E�1g��BI���Joh2�^i{�H]m"
���	�e�ou"g�	�ͻu�uɮ�/����f՜���WGu�h)j�}Fڅued̥l�^������y�3vn�9��ڧı�1�oGg�Iק�v���\���Ag��oj�����&6V4Ԙ��R�$�=\��Q�xp��筴�}9}�T}���;�3�h�6�H�R��e8!+'Q�KZski����R�yT{�[��R��#��Z�2d&j�.����a+~�;�^Ll<a�U��m<�����q�a����@��-�\�_nn�	��u�*�8o�P1�,~��'2���w��~���Nez�|$�T�B0){�Zۺ0 �(���݂v'���6�,��~�TQ����t�F��H1Ҁ�祼�ڸ��^e��7��@���JV�4��]��>l�ۯ �_�-b䴳�z����Fb�I���}��e齎1\ir����=����m�m�&8	�?$��ڊ���*�X�s�+L�h^k�1EwH���uMN�:�h��4�f�:#5�quH����W.�d�^w뎊T��RJ�{v
��[Ֆ��9a�q�����c�ɶ\���W.�իC����W#33�wF�V��0[���q�n�I�ybڹZ�zW�N��c�~}��a��|��N?�M�^}3�������z���p��_p@��k�y�]g�ڌ�Ĵʟ*l���Cy�E����e>}ӷ�f�b��܍y5���g⪡l��$�X}�O���؋��D�+�o6����j���}����{�:؝�y�,q
uWs��M���,�mݍQ�o�������.=\�.� ��4�4by�V�B����$I����h<�U��u�葚L�Dwk�,�u�r!]�ڣ�ycwmԋw��0DN�ƾo�	��8
�m{r=��K�9Cw�,;��j����B�(�3���꧳ч�)����vOѾ�����g2Z�Ć"�J�=� �@��3�\�`M� �ǣ�Oy3j��d�i=Le��P���RE���2hΪ���K�� z�f-v�;qO>�Byp���F�+���˲�
�6jD]�e+[L��.�&���o�5�%��Uv��A�{�nI�>�]�;�B�r�ؙi5��0�W��[�,�x���.w�.u�j���	՚y�0V]��������8�b��A�A��H}��y��o7��0��x܆�y�=n��炊H����R7-��d��j��c5�gksdZ���fF�V�׎W`�$$:���µ	�:�w��_؉a֠܉����ѹְ2�Mʡ{�]��eq�tf�3�ƭ=5��V��u��${H�n�!u���|y�hS��͢3�v���^���� �t����W�(0�2�u�F�9�q9��z2�X��i=U4tf�i3\/%��E�w�\o�i��}�����S#�Nk�[r�sk1�[{+��e.��R�T�:��t�+������憁��+�#���M�]k���`�e��KT�d^�~�z@�@�#�l��L�;��4Q��aT�f�À�P*��q&�`�D״ɞ-�>��6ݙo.�.+eL�F����1@�f�y[\Y�	^���������}��ɬ�t�fQ��"�T�(6���x�z�9��ӮB��:��4���I����"�4����\cytT*���ՃV���L�-��s���"�!ڛ6/�����g%WԦ�7w|J�W��*�U�V=�ƥ��o�eY�-��G�0ș��G����l�E�O���{g&�N��v�k꘦�9�* !�jm�:�����Bͽ%>��4�z�5Կ�f���i))�ϵ�V��i}7�́�O���D��P�r_��ߤ��/q��>��RⲊ_k<f.|�Xӝ~y=j�}�ʗwc��%�)�U��W	Q�}��پ�!U�J|lɣ=��r*i�r�n�-����;	�Qcw���:&ȿR��vs����18����HǪ���z��StK����fA��"x�l�o�
�n����N??9�̓��U?W�7�`��3��#A\���G3������0�:K<A���KrW�&�����|�	}���A*5n�2GbOF��?lJ�	JzTV6����y�|���u�Ơ�I�T�nF�X�*$�X��z��s��l��W��=NT{0�]2[�<a�	��Uwߪr>�Y��/���#%b>gF��'4�H�jڑ����T��rY�o¼��8�5��NB�{3��'};�v�؞G#�w��Jc,�'��*�9�����2^�V��Q��M���Yi�鬭J�lb�Z���b�� }�� �o7������o�� �8���F)3�����(����	kk��ɫ�Ҭ�X�7���o2�D���<}Y��5\�ˊ�u�e�֕9���s�q~S�v��_�Jf���j�������(���G5����Ҝ*�P��sV�jc�!X���O�A�F���y��B���
�z1*�q��x�`����Y�ގ5z�F�\X8}�$��~�V�:��M������f_k����+��_@S|�^�=��B���f�Z��jc���@X�6�wuI�v�vg�:5�Uq�B�R�i�!H�GZ}�I6���D��.����GK=�O�ȀTy���ɫ��+��#�<��YZ�'w�Ǯ�����HT��ʺ�μC&�п�s4��#U����p�ffWٟOğ�U<ԍ�T�u���z��U����sn�sG��7�K:���pb�ыt�tp�Vt�i.掣�(��"���Tj��7b���2[�z�ѻ�Ν�o���5}i���i6]�cp5&F7�fկA�N���^��]���6o+���-m�����:�[Ad�W�&^ƻr*@Wy��Jr��d�zj-l�Փw1���<��ͻ��dhZn�B���
wt�R����N��X�Yw�V(��i�����	]�-��'^��9�Zmә��VmM�{��
�����d�t1���]лD�޴pJ�AH4>�WN�u*��mb���z��),nc*����փ2;��1N%ft:内�k]��p����ܝ@��}�2^,r�hި���f��f-9�*���b-��e�̊�L�1�j�B��V��sSm�����i�gMe�n"��F,u'B�^[Wn[H�.�Z0㛅�73�6.��].�nS�[&g==�^��U\�]��,�	Z�F�ObO{l���!}È�j������̓��|���k����N��֫��V����e����h�';F(	^��z�E3x�v-"i�ƚ0�c1�Q򔰩��U0�V8T���+�6�i�œQ��;��j�,ӑ��l-�č/oF���D��ehJ�3{T#7��t�n㱑O5��JIWMe62�VRv�$�VN�d�Q%�Vd�y�U�%�[TMv!��cgn�nڦ�WM0A�Lŋ���$[�����x���=R�'��Q�QAI�/����h�}ݧ6n󻮱O\�AF%��"�_R繝��M߷GgЌr�S��]�qu)�ث�nfY�����ZxlJj�/c���,J��T�\}�IN!m�n΃�ȩ�g����{�-�t�㧼͊W�M�nU��;���ś��G�յ��7ƛ�Z<�>��׷j�"�d8m� ޲2LBxR��&fC���G�19(J��j��RZ��Rۼ-S2\�{["�zH��2��XY�������x�ej�,\幹w�A�ж���S�Ύ�ɭg�^����b�RV�)-y;zg!z�r�cWm&�e��Z�{d���fkI@mF�2��piIP�;̜�M�f=y��S)P�s(�%������U������͐��Eh��p��ͥ[p���csݵ
�y-�\�o��q�����6믟����-�s۶�<�T��aІ&��&�Әܵ��UY��XV�I��ܣ�R�{df(֔�9��{��5q�nQr�	��sSfG#�V%BY��0�鋄F��&\Xj^�)�e����rfWv ����]����:�fWJ�IY��۠�]��˾��V�m۫�����U�z�٭�er}�q*sp����^��5A�P!�@yj����Na#c
О�㶏.�F�qM�O�&rK؃�7�,�؉Ů-�F��Rb�_iQ�Nx��$P!ݺ���݌u��79ػ�PPPr�'NΝ��qd�$�T���n�\v�۷nߎ�z���ոA��s�����;����Lr�ey���X� H%:z���ݻv���o^�z_�8W.w]s�;��;��d�p�q�}������NV�RD�Tc���o�ݻv�۷������v�_�z�sν�ṸGwb�p��v���w��"�V��TUĩ�H�鷯\v�۷nݻz��קaP�#
+��4FE9�W(Mt�Y�W��r7;��w?}�/��뮘�wn���<<�u�^��͹]�77)�������5������0�vu4�+�}Ξ�	�����;��u�s���ww���c�]�]7Gu����n�����wu!�wq�w_�/N�Ĺ�v닛;���ܻ�(�q8�Nu�tF�7S��.��u��w7Ds�u��.qΎ�wS�����#��Q� ��)Wۮ�������om�9Ս�坉 �%T�R��Pҝ��gЁ�d'�X��F���\�������^��1��}��3R��7�����xΩ3d�4<QUO�t�t��n.~����	�uY�x�q�e�9Ͻ	c��}�c{k�ۭ�R+B}
;��M1/>��î�D�x�gr�irM���n��"&y�0�:W�c��B��q�3�;Y��"�|��|�掣Ws�&3�/�Q�y���	�5�&v�lY���R'�Wљ�f�Q���+�;:��L����g�0�y����X�SS�6҉gZ��ecԾ���9�����O1���A@��hF�z�
W�l��۫б��Md5`}�5�}�!b���~}œ��v��Ej}��[3�h�D��WR�gA���#�88'��6��t}y���U��@�)cj�Є��}~���<%!�}k��Upᙫ��I�."�T�ms��ރ%\ƈ�{�U�N$,�g�/����ŋ#z^��nV���4Yd��b�.�8�9A��Byu��'�9���HN�mm��j���%�ミ[ŷ/+�K93�c=�IP�FF�rf�N�v��U@�@�'���>>o7��������7��C��谞B��tn����>� Ğ)8����D�l�D���ޭ�^��#�=	�<�um`������{=R/&%p�1~Sۻ�f�cz"C8���ϟ�®�ǹ����8YZ,A^w14Y�چS�o�̭W�_Ey]�"�BЧVz���M8L�jlԻ᪲�U���部^�U���g�����c���.T�[��ۓqp͖�ut��	���~Eo�s�����(�%h��\[*ġ��(ikݽ���:O����m�_k��c��_�j�{ԯ8��Fyj�ĝ�ٛ�ݜ��^9�޵�,�X�D�Ǿ�*�U���:։�����Rb�^�q���'�U��f�O۽NEma�{��<�yU/Su� G�uȌ��&|���@��ر�}[��(I���>�yP��b�wE��u�'�^X��u�Z�7�3̜��r	]p�8y�8r��rf^6fA�V�1AlD����5y(c7j�t�jl�m��f��	1 O�-)��S���X�9x+R���J ��Vuo{9��,=h��Nn��YFH��ə�8��UsOT�WJ˭I���>>>>>>t)����#s��ٽ[q�l$�`&TD����se�Mܴ�Ǻ���[;=]���9��M�]��!��	C�R�yhΕ�Ǧ�L\���N[�
-���=-��$�^��$5�g���� ��S��7���-�j����£�͘�� W��+����ㅨ�z*Ѭ�t���aIe�d1�z�q�7�Oc�51����Q�y~�k@�!g=1iH��W�R������߸ǭ5I����mp����+(�E<l5�!(c=<��3ò�w���}���!�b|t���������E�eM�9�G7��O\���3[���������XC���P��&xg�,S�umױ>���fs)]�5��� ���gǻ&�хd@���r;�w���[���螊?9~y��j���N�������s �7�WŽ��3ţ3*귈��i����\9*&!�n��t�.pF������ٽ��ݲ�)f�l��N�!������N�����+֖��ZF��&(�*�K-��Z��;��c��G��n7[a��7�S��U�;[����Δ�nL-����ܩD��y��`��2�9������ٙ�5�3��ƽ�Qհ5�߸�!�� ���8rU��ކsw��q��E_<�[����9 ��A�֬_z��J��|	��J��U>^��gVQ1r)&�u�z���Dϗ�������G8:��i�񌾽Ւs��ÿo�
��2x��s��(��o�`�3��y��v�e�.pƻ��k��_k4�vm�[����8:��q
�w[�mMEzUŉa>�ٓ{o��NNٺFN��� �1t��W/R���m�t��Ѳ��M'+�l�#��g�����������&���3]��:m��֩�O蝻{�7���:�m���v1���tO�˾�=gcS��\R~�7z�|Ni\X��q�$�E>�6�O?�.M��x���/['[+�B#�u�*jz/w��$�<
�26)�<����~���0iS���������
��~�]�̀j2="�rf��+B�%[Cc"u���$|iu�f,�r���QD���USg.��[�-���2�p�zRw��ң��2�=���V�V�A"_�'�!��њ�Lt�{Y#��b����������{�_������_�W��5�5힠.Υ�B�h�G[6�Rz�д���N�n�^�h+�KUE�d�]��,�����!�U]�#�H꾻y����_�Q�7*���HF���\�'f��:��m.zuUy�K��/A!,���ғ�yW�*]������ڎy^��*�ho�Ϛ�G���k�O�"����@�R4��le�a˸�OMȚv��J���}�Is-缈�(���e�v���~���S����e����*<�$Ά�8=8� ��QC�.W���[��;�����ݾ��F���fm�0HZn���5��0���#�f�M�����BA�Q�syq#'���:��v|��'z"˕�#�u�%�Ϫ~�g���溕o{ښ���
U�HM~�I0���ݔ�e�Xn5٬J�����.p�(V��T1�I�pC7��#�v��h%\�,�]�T�7m���
����]h��\پ{j˼�iاc�����⾼�|1.h��d;��6�s�MK���u���9�L�Cꪴ3�*���n���s0w��7����9]���y߾��[mܰ��s�f��_�/b�1�?}��Oq�Ԛ9���0��*1���M�<Gqm�8׺A��1��%tYƪ�o�r���C��fgvq�}�[�Ʈ�.F�۾f�sU�^�>��m;�<��Yw�n�/z����%�j`^6R��^��)y��62|b��N�{JD6��ȷ�3mu���d����"Ѽ��p����!Fݮ�E\�S�d��f�Hߟ����ϲ\f/@���������Y�:�ц=��w��_z�ɋ�VP٫'�S����Xs��o~�����#D�� 3�����FKt�dL�,s`�=�1�����AUg!Y�\i�+]y��)�^(�����+��{���Wp�F`�����[� �{��
V��l�G.#'j�:q�uW�B��v�ڳ�/�2GgѡEi\���+�\���O��p���]嬠q���Dս��nѵ�1Wt�W�tO7U��Yo���������t�]��x�h�6ț`��?@'�H�vZ�͆!7x�E<B�.���=�����;�!�V�1;Z��O�'��ѧ�rA��/�Wp��Ӝq� ��� |||||@˓�>�����5qGV�:�Ɗ۩bwq&�dd���b�%"����:)GU����y��{`##v��V� �P]�k٣@kFՖ�n7yu6F?y4���;=!�?����.�]E�0eDfc&w�D�q11F��+��4i+�A�t�Cv6Sk�XڳXp�"����gC�}��^�<�Z�1wU�^����pG)h�[�7�37��X�(�v���6�g�o�
&�,Y;[!C\��ei���s<p'�<���]�=�P�ũ���4�e�j��A�ꃻے�z�B�2������4�}p
�6���Ƙ�(yvw������LV8��&i[�;9�`E�QzGE�u	d'5,W=Q�l��$_/v�=FT�E�.��^�g1���B��������aUF�f�t,�wa�}4/=�Z5��4��:��Q>���T�vv>'�Jsu�s5L��E�M6����
T�ru-�1��E�=eʧ�4�/nh��������ť�IdQ�Ŗ�˱QobY��)��˴k&7�ǲSb�iHgS�3`��Ua�u5�E��Tc���uS�^����z=�[g�����@�u��	�9��+��r.|M���k�8.��y���*��<e��14S	vl:�6M- ����R����ej�SeKm1m�|ݾ�$�յ��g�#��B��x�26T
Y�t�BO�c�Q��j�8��'
��&�S��>b�՚��E���7�]8��b3��}��Ï�Sl]u��؈�����r�����OO��ߖU�@+�1Re���F�o
�����ח�·k�#z���Z���=������A����%����m3����z��ز��|{���'+�5��+k����y�F�7���H��S����4Qr�tH��kݤbj/��}�D�8�0Ô���!6�;�"��*/zk��Ҋ-�9Φ�]~�������@>���a?dV�l�}M��kur�k�<8NL`����j}������'#�Y�J��l�5fB	�O#�h��q}L�����k��G� o��> �Y��ǽ��/Z:z�mF�Y��y���Ԥ�ټ7��&�T4�S:6\��3d�0��7lD�P�s9S����S�����{�^Mok�yg)��N͎R��uqg>b4�"�U��jq�ߑ�*3�_�����`�m����l���63ݠ��V��sP.�Q�~l�{����qR��g�[��?��ߍ��nC;���2⻖��রY�����F�jz&�|z�� �r������/ל��\����q��ٶ��w����z6&%a'X�>垥�v����*��s���{N��v~�0�!�P�P����NA���k�Q��L��]�pW{u�����(��|Ǝ	PBt�+�z��>���r6��re�Z���%B�L�]H�oi��Ƙ!�uW.�_,�:\��0��g�@�	�mx*�@(��;)ԁň�BuI�f^�q�"�,�^�6*���������vq�~�v�{��<>s��+�l��E��Qf�/t�̞	��;�M<�����4��ywW�%k]�Rs�V�v�.��2��%�w�c�խ+��M�ɕ��(��2��NJ5������"6��ޫ���#efp2�m.�Y�������2�OC:�.��p�l�^#����y�׳ʇ\��*\��1��2�_C�D�S���!��T�`H� ���b��b�7�iI�����Ԧ~�J�o�/�P��]�m��-�[�{ʦ��^/M�m�ŗ�gj��r�/aFN�0���Y����C6���ކٚqefN,�do�ϽMC�R7���h�][9#��t�����MͿ,}��X��#���b���/����L;��S�@q��t�i��r�o>��.��Ĉ�;�I ⟻�b��s�T����e��)fQ�w�èu���g,��%4k��ʏ������:�j�Qu^zA�/K*�������Y�=#152*������c���sZ���� ��'q�<���~W�j��t�tW�_?�����������j�hA������A��4U 5A�|=���B��J�ZVmiY��eZVU�f՘��ҳU�b�Z�R�m��f����cSZ��Zb�Uf�-��,�e�e�6ɒʶVmi�����j2�̦�Vbɕ�YK5Yc35jc&L�edŌֳ�,�i�3�fL�f��1���̲�2�d�3Z̘ɚ�də����ɕ����*��Z�mic&U�&2e��m55���e�-�c��fb�Vfc&miY�+5YY��f��3lŚ���ڲŚ�jm2�,c5_3mՖ٨�jV+6�2�X��jfkt���YY�����[+*��l�5��k+5eeT�Օ���VVV��Yb��VU���Y�+5���VV�ʲ�[+-ef�kO�ݫ+5���VV��YY��� �
>ߣ`6����
"�@b( j���R��U+5�R�H1D/H4"�&�Vm�R��U+-j�f֪VZ�J�Z�Ym���@�D @ 0 ��mT��U+5�R�ڀ��PQ �A�P5���کY�����R��T���JʵR�kU!��kZЉ��"���VjҲ�Jʴ��HQ*�iD��RH�Ҳ�+5��եf�J�BMk@:A 1D��[iYV��ZVU�f֕���f����V���VU��5����e����iYkKU�f�_�>�����������( �� F

����
��O�����������{����?���_��`�'�J?�*���?����� �����?�"*��� �*��?�0�@b�O����C���: �����w���I �����a�?��',
��@���I��TUQ����2�%ZeZf�&֚���kIkM6���4��Km&ږV�+i�kJU����զ�kK*�Ե��Zm�kMfڕR���Zm+i�M�*���E#H� )H!���kJ��kMZU��� ���T�H1�0M*[ii�����5iR�M�m��m3kJͶ�m�[6��Z��Ŭ�lm�4@H�dT�G�eU�Z�[l�i�V���mh��V�U�m�|���'O������ �Ƞ"� �H (�_��}������� ����J��A����q���C���_��CG��m�q,���W����W���7�P� �_�C� �`~g�  Qu��u������S�~���K_�z6A��
�'�G�a�,@g܇�}�� �*���?s��?��? �p >�'������҂ ����?��� 
������D,$O�z}�~ig����j�o�?��0���)3�� �*��� �R�?�,�p4���3���UD^�O���"��������`R���d�Mdy�(Dof�A@��̟\�o|�}@R�U
AUH(T�"�P�T��
����QEB	I���BD�IU�Q�RT@II(�
U@�RQ)D�B�
��%*��]aRIJ��JPRT�U��**TT%$�(!"���I�iR$IP
(�(�$��J�R�U$�T@"RIB�$�""��R*�%%Q"QR*�!IJ�i�U!	p  3:ѩK�u�A)֮�÷lh�4ST��p���n�[w\����f��坬Z�JWv�](�ݧS�lۘ;vՖ�����\�[�W:�k�6�ݬ��n�NJQUUQ
B�)TUx  ���q7w$�ć�]�=&9�E��"�����=�+ҩ���j[
xz��k��6���MM�ժ��38�mZ9ڕ��.\�M��)�v�c5��۵Gf�������6��jr���R��$����QS�W�   ���ZM[��8��\�f�v�wwv�v�nȳ�خ�Nܰ�lL9]ݤ�۵��]Ugwv�m��.s	�-��6�J�Һ�J��`
5U���
T(U	Q(
T�   Z��n��Pi��+ ��`P��0�����҇GE���kdX�
\l�4N����Ԩ��($� !Ix   ��׮�3:@.J�4\�s�P ��j�9�h:�TvUj �8q�t.����X��nN�UPB�(� A!"�   q�H���J�ӥ`t:������]mJ���-�k����N�V�t��ջ�ƇpH�"�J$�P$��  ���4�À ]�l�@ ��ҁ�\;��܎  �wJjѡT��p( h�,4  Y,� n�U�T�(�JA�"�� m<  ���� :�u�0 80 tۃ�F�i` ����		����@�`��A�U((H�R��P� �  Y��: u�  �a�  �eM� [�� j, A���J X P틃 iA��*����"�H�B�� �� ZL(�3��[�� twt  .v� t�J�� �Ght vU`��5`  � E? ��J�A� �{FR�   OLS��  "��	IJ� � ��b�*   z�"&ʪ� A��x��U��
8�����
���l�lE4��U;^͓ ����Я��=����ya����j�ֶ��UV���Vֵ���Vֵ�����klժ��^�_~_<��*��jܯ��Ub���h�-�z��*]�lY��wp��\!�c���PXj�;�a�
a�u�[LZ����!�f�԰�2��j�[,M�$QJ���2��p��1�N�Tzk0Yff��f��s�-G�y��d-X�B�WO�������سz����[k\{��V� 6���%���] ���ѳ���~���)&UJ,�t��*�lՕ*W3`�'���{{��Ko*�}s
����Ve2�v����ӡWxfE,AV�e���,V]h*֪�:�t�1J:G�43"um�.��E�0��#�`�W�QZ��(�Á���T�E̎�Gݭ����6jV!�ij��:@���"��F
�%\.�-�f)0�p�u�DX��� ;����d���1��Q�-���l������- �5���0b�<�bV[l�L-�)�'�؋S��;o��ˬ�Tu�O	�Q��yhFI�:�`q�xݲn�]eb8z�a1KTHۣMR��e��Т�0;Y��*����F��c�k뤑R���܍�{��h�׃ ����J[�\�37�J�6\zڹJ����ܚ�(�+kFeڶ����f�%������h�n�D���)��wpmX�F�����l;���[-�kp�5��&Z{�t婀��!A'x#/2���(2�8�[{i�;6�V.��Z�e-7��D^Z�M�EM2܎�j��l�B4P���A��� �#&���Ӻ��]A1�"%�*&������wN�j�ٰ�����v�Ԫ:��)���sj)�#c���S�Ò�饈��xX�o"ˬ.�nE��e��Ue�J�;r�j��5��+n^�1��b���z��b����ʬ�sA��Y`���{���*�JI�hӯw@ڙ)�*W��v�nce��+X���T�u`Y2W�#7*P
i]�ԡX3hb���x��j hi�H�4*�?E<#rg�]]5�[.;��U�V$+!��z�ZL���cm�eJ5b;���ig��ԍc¬����BdT�&`�#n��ܗr��� ���sr�͛m�d�5u�,�L��B�,mi
��		�K5֒	��Ѓr�a�3oT�V�۠"Z�E��n,UddT[�_j�$aT���b���^�����i,�uY�Z�)SaNl�Me�Xʑ|ᴖG�t���
�p�s��ۙtˢQ��\c����E��E�h���Lf��Y�p����i!a��v�Və�Iqkl]0���71�4��(��$T��ՖK�N��l<߳�*�S(�I���ԓoR��r�7�����ЩѷYm5�Q,6�a������d|��+HL1��	*RĘ@FL$b3KU��2��H5{Vi8��;��΁�jS;N�j�{D+ȷQ�6�͇[5�� Ϝ�����+p�P�m�M��m*���m�:3*�X�$B� �U���b]֊Y���9�֧=�h)ŋo36�ݽ��ʳ�O��Qc@�P��Ga�w@].Z��e,[�A%�1j1�BÑ���	e�8�А�-љI�趄2�+��
.���Br�4�v��e��6��G�֍�6��EmFak'2��UH>V\�tR�������4V��c�q��ذ������a�/qY����ƪT�`�*+[yW�h˒�ۼ%F�60�����h�4j�4�`Z0E���5�l�g1���	9��vHX��|v���H�����*�MZ�L{Gq1r^E�n:�Lbֻ�PF^�/Rݤ��L���ͷ�hV6��٥+����Q%b�ypf^4���R�:t��ɀ�n�	�&�4����/Me�j�葬y��""1��H�E��{� 9�%P_`Kq�tA��MeDx����ۥ�vҷ�n��ۧsYxFA%f���Q$V8J(����m�m��{oX4kJRW��#mEi��*�7$�k7E��t��φ椃o)|]�4q�z�׀���{��b�ڋ�Ocgl�H:��L�˄-��!fە7S�R���%�,�ٛ�&�	,T��y���7/%��آ��A'��ֆ틋TT�����i�T9�R/t*�[�2�����cP@�[{B��U�U��˸1����m�yHe0���n={p+K[k]�qY��ӭ"��m�1��2%QF -��cH��>ytQ��	,f�m��y��9 ��8.��������K*d��ԫ�*)6�J�F6q*�j�
J�S�jOv�v�[�ґқ���d�����X��]����l�:u�4ԖY��ƹY�J��y��ðF�dr��e�%�w4C
�`FigA��D�J"�DLB��B��4Xʚq�b��i�Wg&ɺ����E��5��ڇL�2�5�ĭ�\f�+CN��aşhr#���L4��2����tU��S��'Xī���J�f��,-��"�
�b���f,wCF*[I�r�ݱ1K�'+nv�L%{����LpLb��)&sf���c͡�l;ĳ�b���^��
���]�b�o5�x��M��;���:۠,:86�^R��mR��`���c>�T��ɶhĄ#���,Y�����J	ef�m��s�� -�b+ɉw��w�l3���,����5��wk]c���JU��r4���:�ĵ�M$��ˏ]*J����7�i4iM�n��u��VwU��>)�Ӵ�J�,|M��r�X��e]�a�R�v^P˷��-�p��Q�0I��s+L�NV2�45�U�q�u�X�d�^O4֫���h f�V V�^���*포��nj41��m����c�`�&ݼ0KL�4�/7Y�BɼH*���A� ���ާ6�v(�U*�i4��śu(�[ThR�mkb�:����U֢6��SN�On��[3@&�*��@%�Q�b���+��-v��M� ��{��Gw ь���V�� ���2��7X�F��S�[����U��)�r9Xf޼g�V	�v�[��J����4nջD�3��@�5�L��T�ʻ�W���� @㿅�����\wwF�e�9�%ސN&!��+�4��O��%XnѦ�a�iY�cXm�c}j*tFF������\����$9�س0�jnKOa�,x�w��p;i��ۖ��m�o4T�Iض��6�C.=��,�JR�2�@�M�66oj`v~('�h��+Q��T`ۙA���ܓfʃ�f�\)َe�������5)��v���wW�#�f����dTyx�fST�m�'g(�ŅW`к�U�c-��
c-�a-H	7u;��'[�ۄMk���:"8��`b2�ծ��!�q������U۫�KOވt!��hU��Y��2$
���2���R�w�Mb�F1��Z�����6*�[�1�� EՋ)�¥���2f��Y��j�;���x�][�$F)�Y���e[�{�3�e�]@pĤY6
dK�����YMj���2�ߐ�F�P(0M�m��2N��-u��7nh1h�
��`v�neH4�� M	�n��q�V0nRqXrN� �{)%D/�ܱ�ռ9*��a��.�i��v��;La,FNIJ�$�
Y�T̀^�B�E�n�ң 86H�c_ڌ��Ă�9�*^ٽm�1ۑ�sV�s�L:N��5���/&m6�m���4��0��3[�˗nd��7%��+_�j�Ղ�
�n8�
iI���	9�̵Hn��R�
�4�(�D{��p<��iXh��f�M�����j�9 #I��n@�EW�0̏>���{E����|�e�@��;�O�t8��Y��l`���c��/6����2�ZnV�D5�ۖ��-$�6彲�5h;2]`ͭ�м��cH�kR*J�BU�m^5�F�5+�V���U�dƣ�D�fJW����fDҖN�"��T��P�v�'
rP�Wm�k5;����U6�P+(eƔ��r�dN�4��)VF����VђK��\��F�6�-u�Fau��W���6������W��.�6�=4ͷ[w�S��Jx�;��D��Bn�{�ikZU���)l��k��E*�Y�Q`�t�ց���R�K5����'�P�vѮ9rR�ÐR��\ݡ�-�)��Q
�.�*n;�	��H�;��b��m�2��NR�
�T��l�u_Ч������A��Su�-Սbe���++c�[�ȑP���!����6�)SW3T�0�M��2�YKij�P�7V��m��Lh���ꋷ��l׏F10��*ԃv�"��me�(�6���3i!45��,�b�p�q�Q�r��Q��f\�^`�,l,��E�JǠ^,�f��+���T�m*�N�ʺ�f|�����TN����k����*e
P̨�YK1S^ÓQL��R�x��-a����k�RS_l"Z��L�-Nժu�Z���ѩ���"v���Zq�*���
)����ܡ��	�$۸���5aǚ\`��Tx��)f`��
Z1Ԧe��^U�-\����[qިvl�F%�M�F�j�X��P�/r�v�v��n;	�X�0��K*�U��Q�eV�V��,.�9j�:�G�[��дT�/o@[�&[?F
Edw�	�l��{i/��e+�[��@R��&4�+!��ˁ倢�>܅U�+i��:�CD�h2,��^��cv��2٤�˥��N�&��4K�Y�#WI���qSc�r��5�8�j���U�ԝn�9��0Å���밁���Us�d����J׶��Acb�q\OF�[�#
�9j����-��E	h��

7��Ŷ�f6m�"�����RP+2f���-8���Ɔ]E�wRnC�&�:1L�>��-�ź\,�
E/FK�lwNˬ�ނ�a;�v~q��j
��B.�;L��fl;j�ݬrMrh1+����u�fҡ�\�3\���mTv�l�S��Yu��Y>{�V�ˆ\ �/(]�P\S)�;E�Pܢ��v
z)� ���wHӺT���F��f�u����l�����6�ܡ��҂��Ғ��;1ރ�иɫ��{��ws
��`r��(D�ZK^���0M�ũ6�ɺ�چ���+Kv�����A��uyy�`D:"�v�XTq��d�1�W�օ�^�C�n���Hz�����R5	r�M�ʵ�Y[6ZY���1T�J+F��Rܚ��q^M�5k�mm��5n��m��op	q�a�9NT�xv��{a(��5������2X�X��f��,��d��퐧E��pl��w�D@ک���W���z�ź�a��]�M��"���-��h�J/6�Wvtͧ�p�.�9�M���SiX�Sx��7e��"���1�9�W4�y��LE��j�0��L��[-P`��.f�R^U����`�X4�D2��j坒-���R�[0�A��	���fg�Q�D�ɬ�^YL!D[��t����wZx�6Ĕ���l��Xt��t"�ff2-�l9"7D�b}���$�c �˛�n��8��!c�Y�n'��jƱc�{B��qI{p`mȷ�x�G��)�w�mhe�{�VC�h��ktf�*Cj6�*I���9��u�Hiz�4�Yu� )�ju1�j�;Y�GC��P����Y���xY�d��<׷R�%�1,���Od1���ʸe��ٛb�Ef4�aM8vff-�a���ݽ��2]�H#t�ì��)�Nm]d6/K;2Nf��|31�FL��-�l;qV:,���,e	I�KՕ/+%��eu��ϓ�[b�ǉ� �ସ���HԊ2s;��
	�Y2f�;�Y�0��Ӣi$�q��Dn�A���G$n�o
v.�˻��~ӇTU�vk�Tth"Q@�X�i�F��]7ZՄE۽�&�,ֶ��	BGp:`dr]]�*&��i���fhÆR�z����a�С��CXr�`�^�,�e7�9GiX���Kd������d�"��I�L�U�i"�;�f�h�
��A���[�*$��tܴ�`����aZ)���ؿ��;/q\�YM$	i޺��KZ�� �)Z4,f�L�����Bcr�-Ke�+�]�KiY��r2�d��K��\×>�&�--��g�-*K�{�ț`TE�\Jz�D�{��u�2�t-]1.�J�Q9��eaN�\S%�K5�Z�V*k��RU6��/Ea�"4JYE�"��J����.4�%0��!�{z���$������r]�L�bo&�����<t 81Œ'�doN�*��d�kJ:f��r ���<la�ww�J�n .ңh��%��ǲ���w&�S�Y�T�eG�����4ݒ�[S)�Jݕz�4�?��v��2�ܬI�7�n��H4qYn�*�e������bEۋ@C�p�í�j���٨jԒ�1��VV%[z��w���[��f�uu���E`{"����nP 襌�'+1l��̣[X�qZص�Ƒ����
��5�u dP���^�Ь��Cld�V�U��n�S��BXݑ$�����L��e�P��IL(� T����k�E�XV�[O#��1�r�Qb:��߉K��W@$��F�h^��&��yj���ݗ�N�1��$�yI$��������։��51V�w/��԰�cKyL�r̆��8�@+b.�歽�kA��Sq$t�E�e\L[7��R+�����(V���X90P����Z�b�`�a|o���m�;��Vj�^-	O���t��yb��턭��x��I�tc�n�)��I�l�h�n�޽�J�e:\ܥ4�jѠ�ee�GӉ� �o�XY[4!w�\*� r�&����7
�	R��S��⻍�������Qry�w���B�,K����q���4�vPU}�V�W6]wR��5-dtYUҥݭ�ΏX.}�'lp^�:�O�S�U���g�&�d8e�8��۳�:�9�5�KWq���ZĠ�J��Y��;�jԎf[v	�F���ԉ�ƭ��'+gQ�Έ��)�ufۿ�mm���e�%i�Wj����H������.tM<OwG�4�o�m&3�2��лT��gZ��{��)�����i��{�<=3���4��Y
T�*�6�ࠓ#.�q��p���¸v�QRR����3V�\;{	r6XjK[���,,��&U��;�X0�\F�7ٮ��۹�j��K����E���P'��w��*_;^�nT��lS���Mp�ۊ��49Л�_7��p�ߌ]ϊ���{�u��N��4hZ��u���ʰ6ٵ6��j�d�h�U�+8�@�_n��
�z&Ε|T9�fpΓ�-̢U��ǣ��i��NF�\����޺��W��/.��[��/7T��O�/�R7y�w�W	�G]IA!���l�sC7Ş�v��4��+l��k^m����yKz8(P�_A�Z�%e�WV�ǦE\1����0�
�͚��%̥�ɐ9��
��hB��)t�7��Ka}��h��)����%yʇ"�:�i�L�Z]J�4�1�jC���؆��֭�b�ݮ���>���	\]�&rãG&�L��9�˷���Y�'������*�nȲ�o)Bt=��++�wJV��q�����d�Ŗ���]Ր6WY�J5�;�#9�9��r�.�(E�(����Pт��z�W	����=V�Aj"����u[Ǫ:4&D�ƫ-�=Q�\u��5->:xoLKk�Ք賁�&w���S��P�uml��j&�ۀ���(ť![�b�Uy�yu�l��n@"���xL���w���eѫ����(�8���J��#�cn��Є`�j�XԺs�!����x�b�6ԙap�ى6��S�Uf�T�V�K����d��)\��pݓqL�$<㝄����Tڤ�wدA�;Q�Uo�]ǖ.ή�.�R+靘�K�x�X�x2��\w����m)�[���0u���p�v�ݤ�v��c{)�T]X�0Ji�q�4�fXͮ2�gaTN���gcq��k�s�7.�]a��A�3�Ē��^-z4SX,�5�"�ٰu�Nd�#][q���.�7���$���l�o���ݝ�+���
�Olـ-�Z��Z�+p_dfʝ�Xafh�ޏ+�����o���6��٠��e[��OY�"�멼���Jt͑��G �ݹ��{j,W���C��a]�Q�b���J�}�8^�wk<N��09�;����]��፰��rL���c�	��w�ڶ+� ]�N>�^mG������ƞ�w��|1M�/:��18�Nک%IZ��K����r+��*��r�z&��+���Ly�C�]t���ㇸ���
��
�)��`E7&S��^vH�yvpl�Rq�ƣ�9W�C��|m��n�]yh��Ă�0�Ш)�1��W��0u�N��tr�Ӌ[S5u�84��q`���Z�N4���92���X�K�7�l��7T
�_u���R�\t�O�AC��� �V,��R&��aoWhn��l8���.t�����e���B:�	 |��|��m�0�0-5������7�Ց�6z���x���y��QX��i��yV�Kw��;���C��#66=���>���f��g#�]���,�Dg5b�xk���ۉc�9�O�Ckf,���ݎ#���o`���7_t���vè�wZ��í��7���Ug3�Tƪ��LL�_e[�0ǵX��g\]]z��U��W�6���X����m�r�����#P���S8s�b[�:-]��hGk�c�꙲�
s�`�;��
���p%<��Ж{x8Y�,����9*�|7��2<F�I0�[�*9Sv��x��ܮ�w�pO�|i�����[�UE���:q9J��ts�f

���,�y�[����6��q;���X��;�
幕a��S$�Lw'\���g�V�2�!2̅��B�[�Mz"|�Vn�:ٰU��\�lqRa��]Zy���yh�6�5�0���0�w�l�o��`C��M�ɇ����)|sD��jK�)�y�����;���spf�t��+*����U Ԕ�Vu��[,�� ��JX�=�E�� 4����)a��O.��+c!��iu�-Д,�X9,R�>��N��>��oc<w7"��O�*�uq�� u_n�k߄[O�9�/.,*
47���x�=�J���2�V̮ *�w�K<xI�s ��iY��w�
QQ�].����cN�San���5��Iz��)�8�Nac����p\��y�E^h�6����&VvRdju��;a��J8FĄ��=��+e���5}6�N�+&�+�]�+e�/ok���"ԣ�v��;~�[ݣe�JE�H;���E��[2���V,���l+˦1���݄�\Ru�]��,�����5�b�#�X��C���^��s��9T�u��:�ՋB�F��f��/z�.�CJ�4KH�j�o��iuɴ��͙�vi顊��{J��R9u��J!i�(X�6�;N����8\��w�(N�.JB!��V�t-�u��BTG�9��A����b�X�����h�4��'x^�4�6MtT�Wuw��x���}}�svvS����t5'1�σ���<�{Y��j�m�b���SZ�Hi�#��go���6�F��Xxj����>f骍�G����硶��W>�r3�Ng]��8E�H+,cc��bbs�w��̛���bXM)Ё����b�K�Wpma!W	Sf��l�˚ս���[Ӫ��qp[��}h����Jθu�뭮X��'�V8u��������,?�
����iދ���I
�y�@�X�l�73^���"����q=�+>h8UB�f�MY˨<�**w��EER�/�m9��}KM.�x����ծ�Ԅ���MR�f���^
< u�������@]p���)�G����哛���V��t��%S��T���� Ks�k�kw��W4����={�>"�UŦ�^EQíՎ���A�*1+7/U�nF&�
��l������Sh��י��(��Uc��-�m�S9P���S讽��況w�;�<^czbǮ[��ŕ�
S���uX0�
i�
�Tl�0�8t��Pׅ<e�O/������Y`�u��Z�v�q��$�5�'nqGz,ӹCA �3i�P:���3t�%s]�%_�K�/O!�k���۪�"����C^'}�Qy|�^��:�Zo�;���7�|�o&��Z��ٔw
2��q�7��+v,aom;)��j�b�j�qR��@N��������u�w(]�4�)�9Q��D21ڧe[�R<U�ReU�Yu�Q\��J��ⳇ����8U���P̺�B1�)��o|���G���t���a��&�f>��G��=�}y�M�
gM�s�9��C���;��H����gT]�E�	h��9�E[����yZ%�I-(rZ,�шl�u�e>�,B&!�>�jK@�3#�i8-wwU���^���3y�1�r:ߑX����wd�/E��9���<�!{�x�em�n�܃��ٽaF3�ir�NC\s@K,>�q-��Wуk #5�͜�����W<6*�𸒊��w���k��]�rl���`������"]N^5����Xt���ύ���X~6��f��vͭ��}w�o �܏�-b׶��T"��:���J�[Gf�ݟ*�*.K��vkw&�9��w3
��W,���"p���*I2�A������F��n�y�R|�g7�2ȶ7�m3�����m��F���s]�b\/�hr��֚�j��9�:2�$�L; yx�s��\;o!A���:YWݑ�z���0�;:K&�^�]�j'��Ÿ��"�V��q��n�w��;�*T���d�P��ǎe·��#,�h2O<nN��4�l�u��|�p\�d�������*+9�Ĭ^�˵��[�/ZⲢ�q̧i���t�0��1wE�{��K�g	Afᬤ:Xo4KI.�E6tj�X�(5F��o��zW�sVb����(�ϭ)�R�ޑeLc�����<�ݲ�.��\s��a���|�p\��ޓ{���a�qK�#�dmU��x+;U�i����YV4���p�J��T,
5#џr��^����~���qJޡc��i\Uاe�o90��z0����AH�޼8��l`\��2�i��%��)eT�ѡum9��5��o�.��ۣ��NJG��=λ��4)WR��ݫ&�ۋ���Q����2��j�+���ںk����/�W/����{*f���q�j��/�b��<����H�<*s�gs�z�A������X���!�`U��]���Bs*�/9�Ul��9���he]��m6	��-�������qz;�ψ{�:���d���].���׼%2��-�1g&�\��n1:މ�-�T���]ܥ�k��I�0�7�B���u]@�$;v��P��̔Iae�"�ڙ de$��{X�gZ���\���h�-T{�'�.��sw��)�gZSo��;�*�����3�痚�'�%<Mv+Nv�(���R��ȴF�'O&w;J;�����dHW�X�J9��ڈ:��)���݇=�>f����^*p��7]D�X5T�>:�r��,�!�U���Svu��m�0�L��\j�*Gn`s��ր���;4I�\�)9�gku �B�s����r,Uշ�&���"A5k�Q���DM�4-ڹI�SkGl��=��L%wq�*X�Ew+��<[Vr�x�l|�U�j�M���f5*r���v��B�&�}������3�s~)R���&s��.5��.v&�����H��G�(KO/�®�������u�u��uڄCK�X�z;��)�rS�9���A0Y�Q�r�w��f>�{GK��[B=�@?M@�n�4v�^Ω��Y}��n����X5�vҋa�뺅�GȫL�q��]�u��^w�B�lv�v���z�vj�e��1����E0�s�3�)�Q�ʱ�1�i�X��e��ߛ�[����{q3G��:�ɪːs���I��N�}��n_NO��\��pTUl�<��a*���Q�&�����]���F�]̟X�l��xk�.�Uˋ"�T(Ⱥ볬��2��L8�u>l��콾�������Ä��3�u�t�8-��g��T5���I� kv��o3�����ʶ�����ϩ;[,��TZ��"`�@ih'ך���X|��j�Rb;mm�q�x�Pv
��o���
���q��DT5�l�𤻩�՛W��Qi�V�WY�L�����(�p���pY�x�
�2t��::ȲH��U�ݍ^��������xww�SB!�\��xm�]|�w�o1Z�8`)��Ǘ6�@H�N�o���9����c+0�&h+S�;����h��pƔ��0Ƶ!j�o�-`�tj�u��<VMb�3j��wx�ɚ�MRrBL��6��'.ŷ2��0�F��m��0�e����dm蕴RYx��vԎ(s�c��n#[[���p���BUތ:���	��hT�`0h�5/T��
� �t����\��Z�I�]��RU��o,{���[!��Wm4�k�|$nPڧ�7M ���>������y�.YNA��s1P�j:�]�o)4���=��
H�+mS���,b�Tp�0���R�m���cN��u�Ed������֏&���y�X�^�W]<��r���*5��}z5α\ S~�[�ɤ��ꜱ�$3z��Ҙ]�/F�ٕ���[M_Ӷ�5�g��;}�T����k���*P�K��nc�i��l⯷pԙ�ɭ�5���v@ɽ���ʆ����<��m.�]3��s�@��z���:ĥn��W��T�$�ۺ�׺���H]4��L`�jY4*v���b����@r��t>�֎�k�FvS�N�pΆ~�ѫ��n���$�>�VWU�������SPF��rgkZ'$�������֊�G���Y)7[�[��G�u���'	�*v��ǀbۃ�Pl���ʂ?,r���wS���<��So��y����	uo�SK��>�1�q �HT+���;����]�� )����qou1:�lp�v	l��vT���'v���2jz�3[X�}0��|c��+*�	�o\y�Z��Ԉ�Ec�=��bA�@��g�j�u���r�vҫ��tS��ú��۽Ls%�諡O]4	�&�CtkZ^����ʝ����;�=��nܜ�]��������*gu��#����2�_rMo)�շz��jyZͩ�j�	�n ]Р]�s�V��v��<�צ�mk��=z:v��v�ގ^�W+���U��f�C\ԝsɿ�ɔqm�a���(,kj�O@�.��V���;��Ys9'�����焹��՝�[�]�"Evn%ǹa-5�3���S�c�,9�~�<�\�v�f@��/��P��h��NP�sx*;�2���`]��Bt,m�DN:��d�������Hjݼ�o�gnku���c��ԕ�]�G�K��s}ng�~�=BCW�V��A�;gl�14����'
ۻI��0P�7ܻ&ڠ,�-�ZA���pu^��F]�]�-l7δ��V렌��ar�:�V���f90�~)p�Ʈ$�z��+����'�i�ӝ�ݜu�����IX�fcHr<���Y�6R|a��8Pp*n`�c���;��)f]�ݦf�v��s/V.hwd�=`J}�;'r=/�C��oj��ӱ�6�(nr�#�&��.�MW��Q��y[�@v
��2���}:uݜ�z�ܹ#�O%��#$�H��<<  {��=����{v���$���_�m߿Y���m �{��T�A��e	��������*�.�_+��q���M��bںf�ۙ�z��lZP%�YŊ�$�/F��$�F��rp��lR�A2F��9<�c�{)lJ׏�; 0�i�t싼M���áZ]C:��+�3^�r����n�[���{3Z 'gwj���P�5�c�w�<����ձt��1����ѭ���	�DV�㼹��+Q�+05��2��(����;�����,�ợ�j�&S�<��r�V��.�������t�p�C���Փ�h.p���u^"����-Հ��3Mv���S���@!n�i\�z��y�*g���A(�����E��[j�ݝ����u8��0+d�6p]�Q��	v]��������E����w�_U��k&���a��-d�
��������/�+��Qv�]��B���xV[�!@�e�sؓ����x��%�k{�Y�	�I��]dJ�ͷO4�R+�ԭތ}����^�FӖ�Wv�2���FJ�ehf�;��;��k�� �Q�L�cupW=͉imU�%��=����ɰao��\$䅴��q��=�Υ��kJ=�k~��CcK����,��]ǫ�x/qsC�B�·|Up`+�e�hr���+6%-ֱY�S��o����� �v��e���kjd�v���u�0�'PA��L��0u�lHc��FE+r	R��	CA�=ʱW�NY�s8̚*l�Z�r�b�V�`Hr#�˰���'O ���zVwt�f��6�7k�����'&7�`J9�t<���W�KѬJ)r]+t�|���pD�i�j�����Be0M�"bIW3X��R���v���v�.��}1�ya3��Y4�+a��CM�\n�q�u�ҡ���cz���M��qr����P�ۥx�0�c/n4s�6e��0�xt�<A�>�9@<Vܽv�]r�hL�N�"��k��i↌�Pt(����2��w��PV�.3�����]�k:�r,YδSt[�"X������a0�g�n��ջl�SN��`�)�w/���Y	=$�uu	��)I�,Gʎ^ѵRĜ���,�ꘒ������Z���gOP�&&t���9��u�pŜ,�U��HLǴwVoZ���<�#�G`�rI��=��Q�f�ՏLbH�	v@{r�ڻ%��ٴ�Ţr�p�&r�q���b�Z�
=7�s)X�ک�lㆅ��ۚ�E��oV����(>(GJؗ4��,�U[�SJ����0|y�6��R]g�R�N��h Md�\�Е�"��Y]�}� {�\-ٺ����Qz�o6U����V=��}���	v;��X(�8���{!��5���XC�#��y��lD��7.�]f�3�>E`-����=��RR����]��ńq��8��ח�o:d^����L�կ��]�k�L��mͼקu��4�h]��2X��w N;m���E-��ĳ%��QΚ������Z%m,8wK�n�! ��ڂ����JC,]]�Ϯ��Q_�R;�=/{z�Ɯ�*)�>}{l�zw��k��'^��\8���""Y�[}��V2����v7���n�rZ��h>x��s��Vd��p�~ݚwM��s��diw|��7+�9j��/)Sδ-���,1t����a���}!�n�����9�qo�8���	��_��,[@�>���Uv�Sz��\�uإs�zZ�W�Y��H'��BE�̻oy�J��v�R�ws;�]�;�%��H���{Q�}�������X[�s�K���,#��ڛ�4j���9���b}kF7���ZC �'_^F�e��
�ʺ��r�n5��\�]Ap��6f�o��z<b���:wb�;$�.�[���R�5&Xt/n�^3z��+FmC����h�1���4��{�Vu�U%�wZ��΁�@>�Z�/�N�QL�;3W;�f�$���/�m�y|�R:`k�n\�gI�3
�7"��r��X� B��m�v���+e�ݖA�8��R�Y�p:���#��z-@���7a.�+6N�q�f������5��4���ޔ0�R`R�s�r��4��u4D���9�����q5�v�+���pk��k�$����L�vf�1F��Ȭ�+qPݖ%�o���^E}�6�W���+��D�vn���ug�$w��SYZjD��1����3'rq�[X�GN�K��x�S n��b��!��z�Xp��Y/�U�J=�n�����+}w�l��.�� tu�Z�j���eй|��v0�;NX�0��c�Ek��,.�}tV�m��D��vC5��һ�rg,n��'p����͒���BWw,+Z�����(2�b��z��z����Z���%a���j�-G�^�b4k=��C,���I��Jsejǋ��1]RYʔ%+󕴨�q��z���[���$V�KF�I�CFGH���u��*vgq��#lL��|�B�;�-_� j��X���"h�\�I������,�zVv���ؓ�"\e; 6����b}v"W�#]Ou���X�^"7����8��K.u
#��\h����;(���e��Hg 8�����&wi���|sbQ��TәX"&�a]��U�*�����`�&�����K�/���*Pe�z�V�!�fM�c���2�����Ճ��5�@�]�
Ʈ%�ٍ�qW[-+kN;�a�W[Po�\(���`�f 3��a�ϰ�.S�}֦m�o=¹-�rcIM�ݭ5�a��|�'����'au�'.����`3��Io���Ԥخ�t]�8%�*!N�1�Q��A^�;�����>��^�]�՛Iv:5�`�yS8Y��u��&����5%zEk,��D�D%[�yYK�$�l��n�;����B=�M����,�z����,@]���=�Yan���(]�wj�>3�W��:/�J�eqދ���8�����t
�J\$�]<x�;�Պ\]];y��£�6��h��cW��Sm��E�b2���U#�5�ݠ���ӿ�P���l2��]Z�w^=�nV�<��̜溺x���&�V�Zr�Z�o�I��3��.*0ʰo��ΉN���#
�̈��k�a���]t�:>��VV��F#�p^%�����6O��؎&�Q��:X����J-ˊ5Ҟ��9�W�l
l����T2�f�jM�a7�EP.��8��b�n��Y�0�Ø�!��}�t2Nڛ�U��H.Nu��qu1�3��j4 ϲ��X��Ǒ�q��+}YO)wbx�1�u�0u�]��yYA�ѵa�܂�|�;o�e	z��8yft�Yc���@��M%(W*�<���}��&�kU�x��WG(�J5��y�G#&�/B
|{.M�w�Tb��a�*i����ZM�(�*+�x�Snc�:'Sx�H/�ّ�7k4(�v��Zw�W1\.�UAdj���]��I��P���e���2��}ɋ�Y�	�E꾊����<i�'���ٖ�ְbub�t+HPp�૷]��/�����r�hd]	Ϫ׽(f>����Z,Uذ뭈�X'n�)�'�򻚜��ȳ;{`��VyQ��j�w �説V�Y�TǒJ��]A��g���%,��q�\I5�K�����$�g名7��]�����CP]���^�����"����4t�TCjؤծ���'��P*��+���af�g1J�6�g^�x�i�&�L��w�;��2�Xά�*��2�w;�h瓩rۥ���e}��(Wj}�z�|�_
�4s3/�P�/R�����e�ߣn$34�Z��7m���3�;j�Qʧt�f�1�㮔A���J$](�]$ 6zW>�E��C�r��̆�f�IjF`�ԨZ�s�M�̳���v�̢"��*wR˽��/��n��:��Bu�k�Q%�V �B5����K�%L�\�߬��|�b�*uz��R��B%��Ӱ5 ��ީS]3�7��1��a	�"�Vp�ː�W{�kZ!��$�ި/�s!k�F-^���!�_f�{9R;�
�kUs��2�s�I�`]s����t��iT��#83y����(5�Be�x��D�/ʻ�Y`vL3��6�֬��]-��"M��jS��c&���A�N��; #�ۮ�� �"x�[��u]v>�������c�v!I��zs7��T`��u���VlK���>z�(�Λ�mu�� ���#�I	1���Zu��Y�a�9�b�7����^ٳ*u�3�*EN�ӫyˀ���b�k�g8��mV�h��:٫���fWl�0����k5u���"�<2���6�֗$GQ�|z�-bkEg[� ���d���;k��p��u1V.�WQY�T=ю��M�:�	��M�5m��]��qIv+Uט˙��g��k��v��"�h�2��n�R
�Ru�1PU�U�]\Dl�r��(�~��[T��Ժ�)Z0d,ȓ�2��s�ޮ*\��o-Gz44H�u��������������%]��:I�;�S�|E]&d��Qeۺ��6�u@��æ�gQ]")�Մjr�"�j�G��0��_
�m��4�Wb�P��;�
�{Թ�5{�d�rnl�:��:�k]�|[:�R�����J�t�v暻=�tRa�#�{3�N[�m�:nP�3��ԍ�{�F����gBݥͣWݳW���E�u��\�����yu;�msPGlK��0�W�B����!��X�N��p�YLʃh�5��DC8+3~��]��f�g��(�F���Bʜܻ���N�A��׳W	y����͌^�ei9wt��*+�� j�䋚+$��}n�Xa]F
TK�EZed�ܾ�Bʮ�=��[�)��@7���\�u/���J��ىp�����[t�u������ds�"���;Q&�R�նLP�B��X]�t��ǚF��,*��7�)<[B�X�PV �Z���ֻ�����H���P;>�@[:�ԍ��33�+!��wl+IZ�0�U&
N��-���XBj�)��f�n"�,��ڼѻb*��n���7 ӷK�n����e��ڱ�Z�ڸ5"L��zҤ�ј/A`�;��˔҃��Hҹ�oj�c�;$�Sn����&Q7�$W��9:�q���lDK)8�*U�˫��q��S0OL���Ǜ�kw�U�;�������[T�B[����-�v(gn��쭀�/3���9V�
^6ݛޅS����K����Í���֣�U�DP�K�gdo�z���x\�l2�����ڝ�l������A�v�h�u���5�Rޚ,�e6ݕ�F�Z/�r����T�c��˸;,�³���#,���>�3f`B�������{�����M.;�nؼ+fR\(�i��ju��Zҍ�s�ӂn���.�ed�NQѪ�t5����7pݺ*��'�6vô$�\΋J�q=,F;��'���q�����Jf��E�����Ҭ���9b4o8��GjT�Ζޮgfk���r��D�>t�J�9�R��P��;�6[�R�o��9%i�X�ڨL�K\��.�{����sk�d����B�����D��Q���d?.I��^u�>�v`Y6���ɴu@���\u6H9]���yxo���o�o�,Ҍ�ԫ�j�WR�"j��xʹVk+e�I/1�k�+�XYc;/97��Z���(hɽX�N�y\yw҃!��4��)we� �L>�ƙo�������mؤk�[Ǥ%�|满0�����m@y�	��_G����g:�ꝛ�u��3miĵ�g]�Mr�e6�o�vq�@�}�^�a��]gD�4��9v��5��tֈ&�w,_�1̷�m�T�9���c����ɉ![���;5S�/Uo(*g0v���v��g��"�Z�,T=���P���p�{�h:on�D�0P�;���Gv������G�O�U�UjV�>�Ó����j�V�P�[��s���O:]�F���֤G�%s8X�y�Z4�jP��m�x�/$0'�/W-���v ;^��k���KpG͔woeu��|���-�Y���Y���>�����2�^Ы��s��<���n�e�of�	[pbΝ����J��w�Z6��=K3��"J�"�Z������ۙ\H����5�Ǳaʄ�#�R;N���k2���ů��f�9����hQ$�tS�ݺZ8#۲�ú�ݪ2�\��R��V�%<�n�|������v^�eڥ\�]-ͬ�[,m�Iޥ��QĢ���ǃ�Г"�!�ڔۆ��ks�
J��d<T��gPM�+̕@��o��f�"9Q��n��u^�ɢ�SeZVyW��1���E��qH��T�m������tMc�;��r������b��$9�pP�pl+ t�h�S��+��@.e�W#Qe�̹���R��J�_�p^�A�k�a����T
�j��qc7����_K���>�{���rA|��J��Du^��yͶ4�側��}*U��v�cP�&h���o''��W��*�;�K��[of��F��H�:S{(\������Ǝ3�՗�5ח�"=��tniX�����j�,�o��OMh8�&�2��ײ�`�c��U�%�4e��H���f�%���ھ���k6�宥N�| �n��$�mZ�Hb��7kAp�ER����V��%,�u:�!��c�sv,�g�%nk}ɵ6T�P��Ɛ�Y��òU���|�>*���*Eٽ��F���(���K�gd
�:h����.��v\K(���u����#�.��wa��K����Ҡ6�S���yN؜x\��@_
�R�m�����M ������������RK�8�r�h����ѻ�+J�pwiՋFYk�=Χ��\���t�'Y��[��+�a
����[Y�b��,����Ap-CSw3�����'A|�s�� �-/�7؆,N����w�(6�Y���6��QVy��K�Q��ST{�(g_l��:�FZ�LIbk��>g�̐-����H��	��at �������.��@$�_yܦP�+C���0��4T)��p��xt3��ӯ���H�ҵ�������b���������٬^�:9�К�vL���a b�+)e_��VZ��wHn�p*p�z�V�*����=��;�̫�V�����k�h��5}�a]x&1��#�ʕ�]�u��KCS�f+�ʨ�,Y.�-�gs��yt=�J���f�B��Y�)���tiU�l���5qWc�,m}�j�I�%��p�U�c�z������z�s!<p�M�
�vȝ-��6B"68Q.���֌��̷m�r������X2A���c������*�:���u���Xu�r>��ݦP޳ҙ�{�;跨Ջ�CwB��t�����5s]�rVe���ZJ�#	�`dSS�%ݛܦ�"J���Y��t��x7ג�a��r�(���gXr�S{:�z�S�6��Wu��}���ź�3Ou&V�J}]��	k�=^�ܥn
b��H���X��1΄R��,S�n\�2]ܦ�r�;�vc,�Is�$����r��H�	D��wts���0(��r�Q��M�s��6��w3`�w9�\��uɇ9n��5���.\I�;���EDDc'u��sbM��wRA&��˕�&1�c77 �X��D�[��]�l]�G9�nu�0�wB.\�I2N�sw!ă"��d�%	(�%�(��&BN���r��1�J����i" �4J�F,�5�t�`��A�D(��W�������/���Ʀ�*��ؓȋ�N�8����vb��]�$�v�S��>����mQo�Z����㚹MǶ�+ﺺ�^<;�c���>���0�]T;�t�p��m��ܷ&�Q0����B�!Ŧo_�\�G þ�)����[�^G�z��ߎ�lǴ)^Txn�v�~W�v4�:�u��q�Mv�=]�`y�B�@�{͋�!i<�^��l��K��ƻ	�k�v_���W��ϻ�<��E���s�M�0.b�0.v���}�U� ��F�6���;Im���C0+]���[S��T�w6�"��:J�����rO;;!��6kg�.�S��!�N�8��vV
~>�{4����@��(��F��ƹ:�9���!9��R�B�B]�vӘK��!7~+���:<����P3��:��E�B:�OvN�����J�"	��7}W���{'���u�5�$�"�)�M��ftA�U�Z ����vc�:���5����C�=�5ޑ�����.��*�Eɉ�6*�"�3c�Hh�����gl�@zc��z�D���ni����@j�����
:����}�_��
�x�ω�Pՠ�:�0x��
�]p��qo���h|zS�N09�@7F±m'�J;jˋ�z�E��oy*$�S�NǼw��#�b��a���5��׫����ʺ9�һݒ�h9F�]�gE����t1cL6���]f	�K;B��C�ɮ�<oqqX�r�mGu�W����,ژ��ImW��]�)b�T%.2�d�.����m�'a�x:v��!1e�z�+kO7��M�V�`qw�:+6��19�ϧ�њ��3���]9j�YQ��#[{DE�ͫ��1��6_�`C��TGE	.�"�\�z�� p����,�F:�I"(��C�sU��]X�����Q��+բ�Thu�����H~z���>�Sp��	Xs>�5�/t(c��q�˸��ޏ'�j ��I�b�~J�+��8�_{����z1�f�$f/��	'���rڂ*7��4RR�#XD`/s��Uы;g��Q���+*�wu�et[���9���eH�u�2���ˎ.�f#��D���姸o�k0�̣�]M_>��У�1�ŋu�F��Qp�I�th��"b��+�?��gP�~&���zՍ�ӛ�9������5Ѫ�,p�mվ�G\%���z��\dD����f��ŞK/�{yq��/�<Q�L c+�oÞ��J*���w��\ ?M��\�x&4�*�1ý��'`��n�����pX�,[�R�{VK-��0a�B
d���B�l,Ϩǎ�[��=�K��GJ��2rr�Нt�ñwV�G���n���ݰ�<;]�'Ӟ䧏w�֝���,mw`�D��ХK�G�0uud����ҡsGN�P��dfm0�Y�Vу~������6.R]e�X�g���L�{K�=Ce{�``�}�W�Go���`�m�]�A����N����ړ"�ʌ=E�3Az���ol.��������AS� o�Q\���k=�FnL	r�f�$ĸ4`�T]���Y��*絘@��Q3�a��%V����9ۏ`}�n���5��U�|GN�ẁ�>�3�{���N�8"�@�����kl\��lg�Ԍ�\�	pbvf2����%u��­��3��yQU��>]���^󦂵��yV�3��X*ќ͛�nui�^x��sM<y�	�͟)\@����%+qԜ���Q9��PZ1�y�㋺�2^ ��ub�S��/obp6�>�pRtx"x?��ڀ���N��C�x*�B�۝�2�`�qҾA�Qݶ���Lh�,��O!6�V#B�StC�H��1�rĳ��o<��{սS%H���a�O�7�D+��jLV�+(�)�5�ScE��6b�u-��ׁ2���SGy��>[(�m���b�W藜8�>�zzS�ٛ�S*��9�:M0)_	We��3�	���S�s+�P.|&N��t��+�Ꝛ]��:,���h�n��k�Y"��8{���S��p��	�)�yX�s������=��`Ƶ��p���"��k&rEu���~���]Ⱦ(3Q�P_�g�w��^3T��[.�d�LCHm`�ʩ��eD�?Z�vg��f.0����m�/�-H��m5z��Z��tCX�[Ɋ�������V����ҽBxiE����^=�z�=X�7Y��.*��@�	z�
�C{�	�ċ�KPzg�c�;o�w�8{Λ��v]534f��'I�.bS�s����U���F�F�ĸ[���s��ۯl�u���AnԘb�C5��DW�Y�X���[������q����8 d\�U���(�s��؛퓵��h�P�BQ�;!��4��\Y�ȡJy�F^��2��R�,,�l-���L�K-�>���G�iTV��^�>|���Hp�Ī�Z&�S�z�Q&�}K��
�z(�A/OVj���Nˈ� ǅ�fB�\�S��;�ʟPM�"Y�˚[si�^շ���S�/�?.�׷^w>��
���@�����㌭=���8�`z�G�_:�����gV.�wݶ5X����'������GK��{Em��*5˫vM���l��-�ĉ9�\�XɃ���ժ�"���iG�+n � ��+�#���>�Vtwł��㲗u�E!ȉY�{r�m�ZUJ��"����P��B�ў�ja��[$F�,W#/�u|y�����F�3�*��sm݅lt�B�û�mN�bS^Z��nF�'z�N�:��b�f9��R��8��y7߶�3�w.,}�W�?P>����V����������WÆ)]e�F"i%B4�<撗�*>.���z圏�#�p$?i�Rj�x��O��#��G��̰��k[xl�*tZ۾��ȫ��AX��χ���ZQ=�kUk��1����uٞ��{�G�7*cK�>�=�S=[fAǀ���hx(�"5T)=��Y��SטP�>gpՍ-S�uvin��i�ΝE�C�� ki	�g�Ĥ��hF.(Z��������)�z���z�L �i�Zw�}%�0�_9��ۋ;�*):�:����C�WO��v�P�cZx��Q�8�΍l���q��t(�W{��4�w�_x�����<����F�h�z0@A�BӢ��k�WJ`�(�蘞e���Ʃ;����9A�丙v��[D�ˠ�2�u�a +*�����Ad�J*�mM�ˣ}�� �X�����l��x+��}X�U�'�vСP!3�NN��ՇG(�#�b��m+�+��WE��7�7F�&��1X�+B���\1s�!X�.����Yࣽ��z �z�a��}�tt�Q^�s�R:��OHw���23�yT��Cך_ϐ�1�O�|@U��}�Ǐ6c9�0mFuU�R�ƫ�#Y]���r�n-$�uH�Ek���{K�7����(B�sF�E��ٵ�Y19�p7�9)�pw��rU� ܘ��`UtEf��몃 2{^3u��2��v\�G�GiH����^9��(��xGR]p���"�#�p=Ă=O�J�U.�9��B��K�ĸ�n�]P*p,W�%)q��/�%<]GI��>�NÀ��;e�՗(���#kڣ�@��3`LDA��_z%@�u�E�+G=�uɎ�왜�為H�Χ���
c���:�z'�*~Q�0� w{� xOǺ�0$$-'�D(���/�����J�j�ג�\W�f��=S�]�a����;U0��z̦{Ne�����]t����7pgN�
���F��nhɖn���p�#���z�L��";MA��Q�~S^ӌ�k= �H�r�;�cH/Q�\�W�������M���!`:�������f/�0-��*�4u��v�E^uv�{���ჹ*�D�Yq�p,/� YX �[��ۑu+�p
`�ƱVq���}����X~�X�M<o��!)�S�gC}V7F�lml#+�ӕ�)2����i޴ڹ6�o�4��u�ch)�r���y�)]�oT�3�~��Y9���eH�5לͧLEvx���@cE�����/	�<ZU��g.��Y�
�c5�6�~5���LA�n�m�{� B�Ny+��sg��ܔ�Ѽ��5C�]�`=��M����^��Z��>du´�����nS�����{癳T��v� ��߶�vҩ���+���)Z��C��v>3�����Q��	�Ц�����D7AF�Z�Y�|�\^Z�Q��V��Pǵo�X˪��F�P��+&X�N�2�E!	��DW��e�*�(�8؞������1�'��>rp��g/Lz�=�-�����1s���_���.�)�yWW��+ǾJxAFt�w��nNUJϟ�(��e��fY�����Z��;���Y�Ǳ�;q�s֚���Uꟶ �����b�ڮ�(�`�
4�'�π�iB�c�L΍Y���B���W
>x<L�k��]b$ߔ�>�we�V���:��s��Uzhp�J�0K��.�����O�:э/,���;����kE�zu�!Uo���zV˃���Um�u/C�B�����蝜��lڳ���O\����l\�ˣ<��5Σ��젚�}�k��X�5�͞�����q��,W�y�ml�Ӯ�cM���5�I&����ڸ�����5��+�����iP�0FTG��UEM� 
���A���:Ӌz���u�CId:/$񍥊���eNˮ���e`)*��
��H�Iᑵ'�@,j:+l�j��� {ro3���b�@�43�¨���#!�L�'����,{�����Gln䭯7z�,FE@0rC)��񹅞�f�E��K�u@kQC�;���8����v]�x�y}��>ľ��95���\�e�\-W۞�!{�w"���G)@r{��-��_z�J�w=��ClA9uRxz2�9�����1���Xp�xM�8)p�p�h]lW��b��/<:!~�*c�)]Ɋu��hS� N�`��G1�Jv��S5wJ�	ἥ�n����K��������_I��7ʀ�-z�
�7��i�D��_��N��(ڱ��m��v�N��d��t�gA�ʎ_D��� J8��ɿ�U�T<%��+�7�lO?zltS㍜�m��_��6#�7T���/�,ǮK��F�o��Y�y�Fk�A��Wi�ޭ>;6��5&j�����Ǔ�
��A4Y�9����l�Ь!җYP�lYy��ߊ���͕pT��Zg2�����]�م�4+�|�G�=��&�7��Vm�f�T7��!�V>�:���z�ǋ�cUն�[���4K��������@L0ʾ]E�Z]�u�]W~��#�U��
���8�!n�u���P��<�e*иvI�'����9:���gi��ʞ*�Z�ݥ|V��^�>|��}��c=�q����U����P��n�<��ޣ���d�X7��<]q�N���T=������ixo����hu��~�Z��X	ԩ��at�ͨ:�s�L�=��;'@������F]��b*AP��)n(��~��Bc�r�klp�:	Pp��50���F���+\�D����<� 0�^-��i�2g��<��O��P��̘��뮆��R;��uyV
u=�F礞,O�6x�~�h/y	�ٚ�� F/�*~�f��]0�X<6�|>��WÂ+����IW�]F謺r3�2�iH���o�;5�53 �\i�Rj�x�����#�G���̺���]�Vܪ/�X8�vDr�2* �����~FiD�H֪�]��ׅ�V�*��������w�H���l��J���EBR��Y��낣	�N��J�itqA�,�3�|�C^���-��<�rM�]��Z�R.ܙY7���'gn�o��u@c��V��+ͼo:�]t�+�FbֱU���f�E�x�L�*�cv#�|3�#��.����9��!Ob�T쵏�����w��Af�EX�ƕ�yA�i�e�$0�+ʜ���&Q:��ҧ���\��.���RQ_D�BUC.��bRQ��/�\6|-}�o�WQ{���+K�ަ�Y�nN�Lw��?��<���:�ۋ:=�*('C"������	��9���3�$Zg��H؞j���+&���m�����N�ΎunR�^.��-��B�b-z��G��P�$�U�|+��:q;2�JVoz�q:�dUQ�w��,%��blzX�g�$������yw��вv�������-/��l�c��� ���ƃ�r-x��>�=֒|�o������vZ����|���@��7�t�� �HD˩��sC��n���2�܎`CW`l��x��`������J��`�13&�U��T��s���RJ�t^{ԯm�z���5³�X����U._N��
:�k�
���`�]Ȃe�k:���)S�}-�׸H&�@�t���j7}_M���iO�:NN���v�m��C1�Uc+���x^[6}�@�� k��}��J�@뾋�Hߊ�rc�;&f=��k`╸-Up�K�u1�:Ȭ֣��y���[`r�PKQ�����V6�."��jꕺ�c�	�� �YAgٔ�"ugnVv"@�K�D,fI�m�TP�[�r+���|��MΛ�W:�G��W�L�0[��U��p§jvC�`���d7��t����I�ڬ�__����Ⰽ��O�>U�(\��eL�41��U2t}�V��Gu̇*;�ܣǖ{��lQ��V��&;k��w�-d��i(Ty���fJm��[ҳ$]f�O�P�-�-V��k��m�,��u�E��ԡ�S}����ن���
�Qa]AR���J�gtԞb��.�wg]�(S��h#iU��d��w4�x�w��K��㛨*YDη�/nWv�ܵggu���l��ͭ↠�ʈ^:CtA���K�:����׌�L���#�XT�ќb��M:O.�hv�����7�"g��F��a�{��\)��[�(���;�A�o�Q�eZ�eX:���ّ��d"繽ig/�%R��S��Ŕ:��o8���؏A�c�ޝ�Ѓ���bx����I�W4�b�6�r�y}���1ͺg]��kst^�غJ șu\V_*¸}}�����.�J��g��]���ڷJ��F��,S`��phB��m��X�Y�b�}
F�[�mʸ�˨�q���Ko��a`�m��Y���έ��$��k�aW*���ξQ�;��T/P��e%�ݴ�����<��aݪ��|��ߊћ*垌V�s)3:��X7��J��^&[�шb�L$t�3�޾2�gZ�ĺ:5�;{q�{3Y6�_ه��U����µ��N�y<x��[u��Y�"�+Z����Vr�w��;��u�9�a�ɱ٪�'����Ʌ�c�Y��;�˭;/���w�=:���PzmԂX%�R�vK���FK֯�q��.��}`>�������Y	γ�(�in��Q�7��t����U;p�w��H��pi�{۝����7uh�lQ/�3k\�*��"���tdM�<�+�]���W62�XL��+f���Qf	��/r�k5(B��{�{6��
��v����lJA�z����wt���z<�.���jZ�nj�Vs����psD؛l�:>yi��=2Rw/�w�+e�����e��Ŵ�2MŢJ:��m;��9 ���B�[���-��N��0��X��o�"��٪4tg��͹�Nr�Y�:�!�Uy��$yɴ�fg8�E%2���[7�V�]��m�[4��C}&��.�ޕ��]t��-L���J�N��B�e�Q�,>"�eɮ�kx��u���Ֆ_��3�s�J��W������X�KćR9O��7#'�����y�E��^k�� �t�"��e�����}a8��n����覞)�vr�HΡau�v��]5�))���r2U�v��I�t���ө�k�u?�~w�����()�\3��1��9�"3��FH�hB�D�ݻ\�\�%(���6c1�!�ҌQ`�1e(DȠaD""���D뫳b��,���RI3��a��LI�A"f�wwS�(2f(�LI"SM$\�Y)�Ba�2˺�3���s�v�9�\�������)��M��ݹ	)��a����d��ː����ݮ���"r�D��1��$���D��b� $e	dc́�di�ˉ$�r��R�CJn��I��(��MJRS9�� #�����K��HWU.�t72�r���Ը�Tk{,��on5�+���`f�^4�wu-	c������宸Q�ռz���������>c��K�E�A��zZ���5���[�|��cs}|W��Ү\�����_>v��r�{�u��n�����^��:�6���ߞ�1�L 	���~�8�� ���˴}���՟��2=�� {�}U���s����>}�k��wv�����}_�F��7�^i���ʽ�u૜�����^wj�<o[Ϟ_Z�����[��W��\>�+E}�>%����¾!J����ҍں͑�o&��",G�4�?����B%��������w�������~�o������{W.o�����~}�\�+���7���ק��㷍�m��������p�=9 �-ucs3a�_v�����ty@� ��G���:=Q�UxL���Q�.� ����u�����o�߾m�{k�������彪�\�ow��n?;W-���zW�����"�lI���"!�0>���v�b���I��ެ�P|G�}�|���� �G��yǔdt9>���<�{��������������W�_��x�~o߾�lE}^+���}�o_{csz����+�W����_VG�ϽP ����}
�r��=y���1&=���&F�����E�߭�W��������~������O��W��/�kž+����������=�_|ƈ�@v�_}d�� ���~�� DCGզ3��T91�~Y&��7�ߺ'>�t�y�C���~��|�ޛ��x���w_���o��x�k�^->u�^����6�^�����m�v�W����|\�[w�������D8`h�w�8���1ꁹ�tUҳF��	����� {��������6�������ֿ�{����7��_���~����~���_���y��h���=�u��������z[�\��]^u�����o�\U�s\�/����;����BU(� %:�������T�U��-��v�[�~z��n���߿}o�l��"�����zc�{��@�>�G�|\��x�o�w�~޻W������T���#�=��@����Q�	�����5T6���lv) }�F�!������77��w�ޭʹso��oM����W?�����������^W�r�����7ϾW��so����/�ޞ7�n��~/6�/��m����v���~����o�����?���ٻV��z���PfZ}R�,�6	;E�E�>���0�,��r	[�0�|��KgDVe�R��w:=��j��맘�f�Kٷ����h1*�yt���͚�W�jV����m�zOS�V����!v�{}˫}��������CM����zZ=/���۟˛�y��ޚ��o����iݫ�y��׍��׋��׏�{W��}k���}��/Ţ����ט�k�#�ni�#�$C}"�Gֹh��4c@ϟgh�x}}�`�~��0G��>�  ]H��������(Y o���签*��?|�/�|[�-�=�S���������uuv��x������k�x�_~��~����W��[��x��{�ޕ�5�z��/���*��~o}z[��W5��x�����x���G�{� �:U��G�=��L{G9� �g��D|��T�i�������gF��q#�`�p��1����E�����W�Ѿ����zk���[�wQQ��7�;�����������\�^����7ϝ���/}�zZ7�n����>b#}��>G�7�u������+��P�>�����~������[��^.�|^~W���^��\�]���y�szo߿|�~�oW�_�:�wmϋ��W���^u��W��u��o��|��"8G�<��d�rܸPȫ�fWR�Ƅ} }�>��7Q��>�"���&�+��/>����c������ת�W��m�u�o�|���W����/��k��Z�/{�^���<�ֹ����o�������� �1ɇ�X��K���O^���^��MsW�]�߫�x����{�x�z�����#� �ڿl{��kƯ�>��o�r�U��_}yW�η�x�|_�|�^��5��Ͼok���������U}U�.�o�[�O�;�=�� 0@���3�z`��z�|noM�m�w�m��7��m�����U��#�c��SWQ��P<"1:�5�~5�}^+��-�Q���woB>���E�.�U���$>#��*���Ͼk�����m�_������o�{���ߊ�i�����m�o��ߗ����}m����h����o���/kE����?�����sw�6��=/K>�g�������{�b�����gޘQ��U�����xGH�&@ϝxtlzצ�_�~]ߋ�Ѿ/�7z��-��Z/u믫z~������^|�叨ǆ�#  �L{�ޜ9~��� Ǿ�+�p}�{��P�� 伵~��w��;���u��ɞɔ���.�.�#�Ol�|{�:��Ye5S�7��-��tVQZin�kwF�g��B3O��Y;����c��&j&��9�p�o��y'%�< FR㽤�j�v�voR�ɸ9wTtne��˵��䀿�������}�f"1��X��!��������{m�{���O޽�����^����_��ֹ����\�U��-���o���Z�/~^�x5��[�TT/>�Y�?X�ۑ�����}J�ED�i�p����$��C>�DDo'W�r�}�]����[ڽ���������/��m�{�}��^�ޛ����⯫����皼[�<W�:�W�޵���ۆt{��,_��(���?�P�(|�H�/���5�x׍�^/���^W���6�}>�W~��� 	�=^���~��/�������_���5����^*}������ͻ��ʿW��o׏wן㦠R��qe�E9?{� 
.���~/CQo����oK�޵��|{�3�}
�dz��=������*�y��׵���x��~{�o����������כ�rѿ������~���Z{�Rsȑ;x���+�tw/�#�$}+�6{����_o;^�}\ߍ{��=v�6�W��K�o=w5���6�������n_V�>W�z�Z76����m��^5������z[���W�{>�>TA����1�Hw}��xLy@��ׅ~+�x�_~w�~������mp�+��?��Z|�+�^yz6��������K����~^�|^��LC�{42� �����'������x����,_I&�{df�lm���ﭹ������W��{o����������<~^�y��{��\�ݯǍx����;x��x�k��sŠ؋��x������o��x�םx��s|�軌�1��~V�$o/�2�.�� ��_k���[{�u���߷��+ם}m��熁� �Ǽb�~4{� aG�}����"���.6=�N|��ۛwv�ϋ��z�o���F��� #����Ʋ��3���F�9�#�Q�x|2����(G�@����<"=�&�xT�� [�q�zaǂ�+�V<.�	������ �1�h�h��z� �}4.<cޚ���R�����=�/�44g�w�ӋTmJ��_� .�:��v�"w���c�;�<�sq��g�1���W�I9;e@l���*ї�Q�m�q�o:�V���7T�[N�ˏ����L�{)@���E��ս"��4�/�ݵ���k���c��u��ns�s{:��(]�\��ӹɊ��Ƽ*"#�s"^A����E�#7�` �Ny����y۽[���� V @���2�ᵳ��Wr�2���h�S�;W�{�4����Ɨ}h�0b�y]V�I${� (�ZpyL�N�=̈́p��|~7w mv$O�j:g��<_=��ވ
P�",	�H}Pz�I�2J�gn��뚀�+(({��J���铜a6�쓙Xܺ�LgԥⳌ��PE\�W�J��ǃ�~5[5����Ij� ���Y8���p���F�ܧ���,.��3(_���������| �Ġ�Xk{C��L�n��7I���e�����c�6�(�j���~�����w���:Aw�@�ւ�.���+��>��	���Z�����ꗕ�r� �v΅J�c�N��9�$�ܕ'a/X�ɑ���j��{�C,U�[T2�>�</��)��!�g���A��롙���Jk�_�[�����մH^���Heocў�o�}��
�Gk�മ -�� ��`t���}GM��+�-�]_c�`wf6;A}��>[�FQ��6*R��7�!��s��F�}�-9z����~���+q��H�2��K9
���ܭ�J��(d7���e�)���,�g8�9w%[�T��^��J��M��F���J���w�l"�S������B�ƶFlޛ'P���r�䳢-\\���!d�7 �\u���p���wf�\@�
-�NF|���y[ѵ���΂N��T{h��|.�/#�h$˄�.�`�b��S�E)�����CU._H�
4�5��*�r�1��L��^p�R�����Q�z(,�M�#%_˦.*f5���w,-�zw�!�e���b%m�.B�<C�7ˋ�nʕ/�LAw4b(D� *8�ڝ�ߞ9v��O�Xc�5Y���;�ݙ`���ER�hn�#_qT	�wH��&;��8E2g������Fn0ifnb�=/������ �*őD�24���#���gwCB!�f�;��.�t6��u��P��A]�X"�X����\��TWiQ������N�K���%��log\[Z��pt��%���SO"h�R�B5�*��&!uXS�A^��:��⋽��V�`�P�K������^���sp-)�T���e9b+{���+��-}F͇����j{������������;
��F<8]�8n�-�Ͻʀ!Eb�ɛ�F��~z��:����q�7އf�d(WY��W���ba���s�u&{x��~�^)�q������7��m1eNg{�׮��Y}�st]��y><w�ڃ��]WR>��Z*Qλ�9s�T��Qc$䱽ϰm���љ�������*�{#"��V�����)�!�Ua!\kr��W֬-[���G\2xR唋�37)���v�>�]hj�t����y�q�k�{�	���>��QX#|N��uڤ�2&�eM@�����F�8�!�.��00�Y^Z�Q�� ���XyS)�����M�7�z��]/� >�� �J��]0B�������^Ԙ�ړ>�G3c�8y4�NOLk�UYuM��-T&ہ�P* �����;�����(`(���y^��=1��֎9�����`��V�%�Dm{y]WZb���{C��t!�:�9O[v;X7�N�=Aڬ��i��lpᤞϊ�>��SH(�UFX�b૧���Z�������6Sw���2�T�	Pbvl'���񯷰���(�wO�"��.^���&-�֕F&a�b���:�z}䨏q^0E��<&�*���� "<,JV"`�b�U�1(�

������b�iN�u��󭽉��ʃ�.
N�OZ��EANJ������eF�T���E��s�6��[�E-y���نl�z�X�}��b��ώ�������/ZW*L@����Lu�c��.��d���#��P�)����$�{.�Wm:�FA��=x�ב$��t�7@@��]%g�+�7o/O6�2b��s��FH£��:/����Q�k�1�S6��F�G*�X���x�kss���#֑����(�
H�NO��X�7R
N����so�sj�q��0�Ǽa^e��@{������O�c��/Yb�a�~p�Y�禃yv�T�,�N'�5/= D���3A��Vz��u^��PDOd�i���ʀ�:�l_��nЦ�]4�W;$6�gvv
5p�p��:yb���궅g�'s�`�������t�4�,���qlX��å�e�oAm���B�^�B���x*9eD���V��=�׵�%�hn��ף��P����*gg�H+`Z(Օ1|g��y��U��p�	�9���R_\{�L2�{�[�y}�(͉��=�Dr�1�]�"4+x����@���>�����M���n���tJ���	�P8x]?&)�C�ʲ���Δ�]��N�*�vO��������;���u�KC���Fw�" П#54mF4��>@W:�lp�"� ���<5�=�E�D��{@;�#df���Y�X{ ���q�u}�]K�t�'ݻ��kB�6�9ԝ��S���3:�u��M�����8�7v.EaW ��F�"gnn���%�6���Qf�7�:G-�]��2��B=����J��#r�=I��p������g���x��cx�op[����z�Gl��ᤝ�_Q�\�ew�Yn·��J�=���n�S��m��j\��>��ӏ��:�O�>�*�@�Q�'U߫{\�|Wr\z6�|�PH�ґȎ����l��C�gC50�u�yx�hs]d�V��׸3�����S\t�TFTq�R`p��h뾇����o�w���N�E��e��T��J������cԹ��:��1���O�x\���`��w+���Q�W5�Z���v���Q��c,�V�g��OJqr~GI#���Zpy�t��m(vx���o׵�Ih�1��W��~P��'�)@yH@g�ʐ���~F}��2��N�k�e3^�����E�[�!�0���i��i^T�R��JP+8�Z����'���<h*z�,��$Z������s�M�{�l-�����I��|��2���Y�$&yI� ��O�r�=�zWJ�����(�Yk�:bx�~_T�^b�W?V�O���:@�n
�N$���4o�*��B�7Y31�Ai'~�.��:��Ƙr���i8�'>��5��+rA�]�4a����5�v��t왫ِ;iK�B��j�6�Wͺ4l4͛��0n�4�J�2#���x��	��JԲ��5�?� �;ZAJ]i��Y� ���h�-X�o��\���U�߶W�sv>��VxQ��I�m��.rc�V͝p�g��1G�
�]]��*�/�{O�vc��C�� �oM"�3zt�8� �M)�텚��7v5�О� 3�e��x"�ύ���Z�!�ͻ{����ʣs7�u��D�}1���_xc�g�ٍ���=~|�*��3&f��7��:����;%�L�D,.�P������6�&k����m�ɢVw<F���$�U�0����ѱ���/���؇�ΰp]T'F���k9Z���Q^8<#��9u�X垑�a036h��[�ZS��� �'�HS��]�Lj=����R�c /�%<]GIz��X�{ob��Q$�݌!��ӷ�P���ê��J.���8�ڝ�m��c�k�Y�U"��/kQ�6�cvL�.x(�������{���{�
&0.���{B����^Ys�_]� x(��a^�F2 !�	��x�X�(�#�F����U��B����K75P�VP�3i�z�I��Q�|��n�9į|,�1�1�EA,�y�O���$á����w��b9,��O2/�hV�j��k͞Y�S���kuL�z(�{�*)���JV~U-�vQ��.���2> \������$/���k��DV�c�x{���nq�\�˩��+�+7ơ_uB'��pU�/��*�	�<�m+���[�e��dp��.���m}�#��5�8���w|�؈���%����5!8���p�(a�� \B'���;
�xł���Z���w����]$�X\
y�#�󙰝1��dxy�~��Gm�}���Pg�y� 1��ڳ]�X�F�f��~5�x[�LA�u{%u���,�T�t����1˲�yW��S�7בٺ� N1k�`�+�}�^�o�X[��z�m�I��{Y9�r�s���l?C���*�:fjl���Ͻ.1wZ���Uu��_Z�ŋ��ڎmX��i�Y����w%�w��݊2C�T�È�AƣZ�Y������o�F;2��9��7�5�$�+s;7��z�n�n�j &{�(A��"�.˘�+�(9�Nv'�E�W�&:�e7].��Uj&���j�:0Y�
	B��3�I;���Ʉ6�gT
;Ģ��G)�{���]��H��H���\�*��Y���/���W�Ep�k�)���С]W��x*C}BI$��)�J�]�N���j�Y�R9:� b����YBQ��Y{F�X�ZwwϳF9������M+A|�����\�s���g6D��>�ָ��.�M�aaP�]y�*�;�
i�gZ
�w4�+yg�8Ofc�{x�vV�e����:*t�HEa�Np�o��ٺ�ȰwBǣO����QA9L�����t���=���.fw�P���!RS�nL��.���L��``����3�L���n�<.�t���pl��*���a�;dx�Q��v]F���f\,:�t���eЬ��
��VP�cM{Ǯ�@Hg��^R���� o�x߇ue\YtiC��4r��c���W+�m���|��Wi�����\k��	��$���]D�R��l�ތ:[�L���V�\�!�eK�e>��ִ�h�xxݺysZ���R�퓳�[]���s7� �u뿂n�i�BF-�j�c��8��z%l���T�6�ѭN}�sz�ֺq��smL�B,]�ӄ7p1r��A i]Wd���nᠹ0�)K��K��qv��[N��_]�Uo�[�Ai.�ӛľ�Y#�C�uX;x�"1H��4�C��5���qOP�;]�|Nurs�M4�gfј������h��t�'��P�U՝le��p�ݮ�^w@����H�i��mw��S�P�Q�x�X�+w{�
�Z�/�p��܂':����XG�NsJ���c���29�j�� ��u���:T�R�9����V�lmpV����P�AMR�o-�]\'"�����/{��85 ���z�R����K�j�If�]F����;��2��(�+e�g�S�Ҕ�Gg=Q�[��j��c-e�&)ewƓ�Zb�*Tm��8��R�������VS?bx��{ݘ����2ʣA�s��;���Ϋ[��fg4��E������Z��Y��]�p�=֞_k����RL�*Tz�&��6���u�챉����< �Ы+�6�; ǡ�d#M��!�3��W���}�v�*n��W׻���܇'7���.��z���,���WiF˭�q6�C�2���	�2�xA]��.+�kZ�
����Y`��ͭd����R��|t��P����
�N;�p-�#�!\f��:�T[AEn���u
�sd�6�)��`�}�]�������`��I��*�g���ґ��i�'j��̑��$���:�2$����[8^5�x^� ��ф�g7ÞU���b6f�e7r�؀�I� ��CM��1_cׅ5�Mj|�����;��]L�t��2��[�n�iF����*eګ#��9�ou�A���c��&�#�k��\����o��V�B��N	�*�V�V ނ�Ꝼ�Z%����Hp��7��o\ňfW�<��rD�,�,��	������`Ag,N�W�����A�QF��gr���ڰ��5)JSFf� 8���T��Z��?9�)��D�(E;�`�	9�!7F�4�)`Cw\&b&��I(ц#��r�w] �;�&��ˤX b��Rdb��E$�iQHCD0��0�����LbD9s)s���s�F�)��w]]�cH�4ȧ7gur�wuɘ0�]"�r 5	d��3� ��
$�0`�HC���Sb#wW`BI(҉����� �Iˌ�Ww5�r���,&2L���`Lc&4m2�3�B&r�[�a9�bNㄱ(L��w4A$�	3&TQ�$$�`4IN�XI�wq���t�E4��̙*11��@�-�fgu�`�����@MB���v�&Ȅ�r�Gu�;�����2fZ~���z������
�2$}��[�|��ǉ[��i���˛�*y]�6��=B�oH5�}��Y��>�3���ݿʯ����*g6���pE���wүT�:v�
I'�� >��SJ�:������ׁ��q{�=�v�5�xu�Y��.b���}R��r�p�4���x�=�DION��Z�/M��a���CW�ⵀ�yV�3���c���a�n�]p
b"�rQ�vI7�8wH�*�@�Zv�L-9۵�;�>�qNV~��>~pQg�'�c�7/�x��z���w��I3���: ��B�
�P3��wm.(���	L�'���2j�f�ݭͦ|;�'���o��stFF�p5ʼc�٧�Y�����#Y�ޒ�$\'`�**��5�gS�K0MM�����[�3��_�CO���ĥ��o$(�<��u����O$אG�Uu��
f�J +�?X��.d������Ƈ����^]b<U�;#��lN���*�gxhH՞��b;�B5�b��M���2�9��"'!��Bl�Vt-s��P���ެ�될l_���_^_��@!a��@B��R���<.ʉ},1:��BS���5�B�^r��8y�\"�Ƿ�-8 ],c�uV��p4�c��f`�Lj�V��uȾ�̙F2�A��m���bS@���8�o�oU��8�E��P�,����.v�R�N��aVgR�%�ڤN�	X�CN��uФz�q�P�1��w�U�UW��D}�"�\�����M��TiOd�����@��o�Uw����W�_N1�ʰ�7��ED��ɫ�F͓�X����ؿ�!�S�<b��]�"7��'-��t��z�v���z)o��8���Ln��G@�<#��U
N��g}�DT�����ڝJ�����+C�0�H�!��\z�U�J�������
�d��-㺜T��q*��FA`CK67���F*�!]��OT��,�=t��g�!i��߻(a�!��=D�E�hz�(�89�ʟW����3.F��0�p>6���<�6O\t�7�������[ձQ7�'�w���5����gz��<wq�J��6���/��n3x���l-���Q����7U��� �00@]4u�C���s�Χ����z)�f��{�>C�{�gJ;ꭒqbR���@�@����bb>U�p�`��w��<bG{J�)�)�Z�B�7�w:x�Fx��w����)�N.O��H��AG�8<����I�k��W��s�k�h�3��ǒS��^�������<]��#��K�=��M�V^�6�ބR�����4�IF�Cza�3����6�!��Ŗ�8��|;�"�Ml���t\Dh:�K�V��$�`��]��zLW�zܬ���:�7@����������\?G�� >��e��On�L�J�&��P�����yR�RsL������v�
.D;�\q�_<��s�;h�^�Z"wۗ�7��M���R��Yf��Ll��]�R�D��c¥H����u�V�$���aƁ�E0",��SS�l��fP�Z�����K��s2M;]]�w`� "�����?*��u=�|pt�6vnx�d�_9�����o9OaԷwizr�km𭼃�9�-��j�F���K��r� �w��.ocѱ���Z*�hc��j��f�N��v�횰ძ�#*�*�<*���P"���a���������'���W��&�Z#|�Ʃ:�%�#�9jU��c���Cא\{�3ÖK;2G.(��@_���Jj����1����=~|�*��3&lT�5�~j�N����]��@گ:�\� �]T� ���F�P��'#5n�}��u]�S����=ٵ�	3�% T5Tu�S#DW�P�7��3��aZJ6�]K[:��w*W�0y����������`�qz�<����o$i �1nY���4ܑ-��-�%�r�7�x4���}pм�D�׏�_K���j陔�Q�.�퓱�K�P���!�γ@w=:��z��A�T3�vDEv
�;F�Љ}[��ӝ�W������>�\�p��<���>���7�$���΃P
cQ���x�0\j�⣖p6a��]p�x»퍞~���~j���(�}�:� :�j�^�{k�1;U������a�������t��炌���^��mLj��?�����Zl���ʞ����u�$��t��c�M$��)�q^�f$p�0i�$x��+����x�-��l0{ܱrT�h��zl,JÙ�ݘ*�@���X��OV)��N��Tx�.���݇H�g�/����ӌ�ºl���F�ŕI���n��7��b��i��1@.<eU��D���X���: _/-��]�a�]���]��1ا�J��`���UF�9�5�����#%C�� n��X���]�kVm���ě�)���KZ�o80�����V���}8����Z���@ݚ��5^�\,~��u�o]�ȫd̬�����lNl�֓���?�z\b�V�
��ϱ�y����e�aecR:.ױY����vjjc,/{��(w�rR�cEi�A�m^��KV�'��	�zc�s�aC}lf�5��ҮビQn,��Bބ���'��Zh֑�i�D��u[��[`+"�pr�4�G>�kxU�!#�����_U{�&���
�(�T�2r���Q�J�8��ƣZ�00�c^V܎Fɱf��B��9K|�����^���1Ma�P &7Uj#�~��(Fb�q��*j���vx���(���>
/$�O�a,^�Q�C6��e�A�S.]�'I����7n��ݼ�-��|[��K���51&�Dɣ.�Z��Y�n=}��j�͛傗ol<y�+!0�C�MX|D��>�Ӱ_$�A� �<$��3�V�9��+6�YΑ���tl`,SR0>�s�.Ǹ�<L�ʑ�F��JW�Y�!P�^*oT��}����[Ξs�.:r��%$f��z`��*�	Jd��q��P4[��dEl�۝{��C�v l�&τPFlD�NҘs��9Y�yPr��	{y�m������Q�%zl� �GDTI�3 ��g�����!�3��G�tz�� �g|ʦǷ�;�=�=�w�ĥ���"=����ʼc�٧V{����:�ѭ��^��K�Oo&s�G#:U����%�Gf����K43�JK���X�R�ƛ�ِ��*W�����2P�f�m��%�eD�-	.�۽OwٖA��ս"��ݫ�v�Xȼ�Eq�� �*�+1�K��[M`�6./��vD�".�2yx�}�<=���9�{�UeΞ?��Fu�ƣ"�P��'��7�rk�Ճ�м5��ﲹ�0�����R۝�ln�R�U���C��}���n��uĎ�Wl������7O�gI|��x�_����s�k�a�.��.wo�p멹����@�΢d؉�fqf�S������aj��VR�1�0Ta�o+�� V}�@�	z�
�G��'�2j+_��9	i2���Q:X"�!�b�un�tw�`�T0������#}�\瓻�N����G�]�����p�1��rN%����6#�=����|���6���ܰ�c:P4d�����,]d�L��tI��+u��0V�1O��q�e1�įN��'�}��)�(F|�yMh�Ou{ݑib��vqp�^ҷ.pd�8k��f»����1 �����=��-��pZ��XOT�o�p�7�P��������leq���lȧsM�z�:#*}C	��Y�r;��O%�����@���]��/o�7;aD4lLw½��2�X�y�=�
�:�GkN�9a>ɼR�s�]�`S��9ա���+|k�wq�\��yCMĪ�d2������;�n��ta���y��oV�6�4ݼ�b��|�Q�C:PDp������+����W� x.���J\Di��v C�5=sFS�Z�禔��	Pp��50�yQ�1z�D��n�:�8t�w�����F|��4�) 1�A�[㢧»
������{|}�J�y�(�]#������Z��cv���H؝��1��
Wr�� />�wؘ��W��xn�v��t\�(m�u�c�3:7��3=�x�F"i%W��k��2�R#����ߙ�4����a�/��`���x���/Y/�:���V��)@yH@g*C�=t���je��$�ubv��V9+6լ;#l���iۯ
Y�s�극�e��CJP+>�3C֤a�1��I���*'�t8�ST�F�+����du�5eܮ�an(+�o��u����/�
���ؾ1�1`�Z"oz"_#U�Ң (��pOֳ���j�ks���YG�y
��W�.w�,k��K\�|�\=ao�� ��U�3�V�׆���*����`$:�֯E]s���k�J���+(|�.�#��i�U�1�7�p��.����3�+�BS+��Q���_�e�����9���U��\N��v؝����x:��i�����LLi�e�>ڽ���j���
1�p�c�����5J�� O|�!�6v��_'K:�c�㷢P�:���ꓯQ$���pW9̐�h�]������^Si��  .{5Y�9}��gLe$���v5I�������g����FN̮�&��I��è�&�#!lg`t��H�r:�D�b(��W��ٍ�ߧ��ώ��r  �"��j]��/�K�0��h�˚W��Hjl@"���-�qBx�����U�PϚ�ϔo>Õ��.|�W�Ь �v,-�멑�*$��n8���K
�Q�,G@Q��S��ȬC��/xt9Uh��Q���|i�n]�3�<�_��t\n�;�7O^�{#�9�{����u'=:g�a;�t�˜� o�P� ][�N��Ph��8;���V2]k�L�=v��Wu���&;[��my\N�]?$`#︈���0{�$�I�����pW��X�8�pc�Do� �_w.�W�Q�F0a5	*��C��T�Zh�O�lے+�\l�Qoei�Ř�bs/�j
�����=4%aɨ�AX`@��1`r�@��]�\r?���l|�z��,�����t�����~��X(ؘ*S��)��/��d7*V���}D6*��>Ů���m�t]�3]ɑ��r�c�����Ԧt��ǳ�I���Ժ�ޕ!!2�Ɗ<���8��g�]f����M�U�/�2�C�\�\�.@��o�ɳ3�a����f��^L�{��޲�l�P4��M���0����� �����j��������q���\)���}���b�it߉�����R(d-0[�F�V⮮Rٙ�Ω��d��B+��e�O��a��j�(Վ�5�6>W�S�*4�;��4]Wƛڦ9�����\��#>�* ���J�p�����R	덯������)cD�C;���Hu�����Q~��6zp�^S˳n��T����v����|��N��
�PEaj^����O��Daf�w�+��3ҡƣM�t���g����ESFD<�u��u^[�HgL�ƱT􃪶���2����g�k�
�|��_��� ���G,�wY
.�S���ywZ;�Dtz�������,>i{U. h�6��`�t�x�3\Z�b"&�=9�᫽ų�b�v*f�t�S��LIexk�+�K^������+�
b�k�����Xn��8V�uЅ=a5���w��U��pᤞ�+ _P>��]}�n�f����kU"�ô�<��]��>�c1���ѐ���T��U�R��ڌ���9õ�V��Ċ�vv�9»FH�K�^���Dy���ζ�.nf
y���A��{������*�$��µc{���P�ƃ��lg[�#M:֩��e:��6��k���]�C�V�k�j=n�)��x��8�S�� {��F�|�0o�E�b�m��V"qN���q\�S�n���gfw�v��s�e�3�\���*F��;��$,�_��ض���b!������,J�v�G݂
5t��z��
��k�a����ʪC�ʮ۾��3�����:�%S�3��R�ՁH�jgzN"ep{3"�%R�4�l1��^�6�,�ׁN
L`��̓,� �t�֭J��e	��7� ����>Ս+�Xt�ϔ�_1��Y2n-u�ⵝ����录v����u���ս%�b�_�ۮnw�cf�sx�C<�<��y��޹��Vc�񳅡{|��^�Ƴ���ߟv�ѹ�b�c�n��4�~��,^I�ix�d���P�X�d�(`
����ʍ���׽׳2zyv���U9~�J�oP�u��l�Ϟ:۫XJKr�SM��8�R�L�)��}�KPR�˩�oa��0���\��R�ˍ�:���pg	�`��Td@�`{hc��HZ �R�)�DJ�h}�a�YC�D:��;T}L]r��շx��O7�l�+MoB���)�	���yS۾68X��VJ:��5z��ô�k+22�e4,�;v���+��x��b���0�ͽ���G��9&��ϣ��`���Y�`͂o^�۾f��ւ�l���R��yܛ���4�������XЉ���������7��*��;�5t�\o�c�; ���B�2:t	i�I颅f�r�Oi��m����1�`�)�S��۾3������{��fp�A�B@��n���X���ͨ
��k8��g�#p��vj�ܰ;+@���fd��gZ}�5���f�r�9�Cm�O�s]�3��Ś�"���
��=����Ua�W�y��a[z�Z�Ms��*�pn����5��ؙw,��0r}¶E��5�-"
T�]oo����Qh��.��}y�+�3tQ]O#7E\z��5�@;Ǆ�(X{w���ϵM�V��YxV����^m)%�'8����2%?\Tk��p�F���֒��b\C/bF�\D35�m�������G9]PsQ�*�����\{G^�f
���Mj��r�݇Zq��Gre�$ç�pvDj�c_)�z�+{�f̥͕׵��!�Bv���)�P�nWK��s�l;zW#맶;`;RTݓxŶ]1�ekj�u+�μ�͈&����[6��_|��/��{]*�+����6LU����,ĺ���s�o�\D1I˾�N��#��;MD��&�\ZטG0S�﹋fp�u�A�J��(^��c�T�	�:TU#K���y6���>�Z�k��G*��J��ЂR�|r�:9���`Sg `w �2�`� ��+n�{3.�^ji+*AtH�P��,�.Yԍ��5�������ڑ"�ز��#�÷�%)v�7�\����䕬��z�2��i�Z�ҫ:f1˰Ex�[�mZA�b�ϰb����D-��ɕ	=N��꾣�¶NJW,]�upd������զ��X�ٴTF��k����B� ��s���}��կ�wu�M\]J�h�X�꡵��j�˭*Z�+�=�3$[�q6�vEU���ObX��s��s��9z�L粕�]8�����܋Px5)\��Q�:���ǄȹG�?v�7�$��tA��k��xGl�0���B��^�NT񝧿dQ�x�� .��;끵����m�
��U!���9C�`D����8�)'{��/�k�x�ǅ�;���e�Kh�s�Z&�n���z��[�r�����se��Ij��]i�\��� ��l���Oh�*�L�<����֛u������^��޻���y��%1���H ��)�ҹd��`B%�BT���3N�te ��u�!��\�R�)�h��eI%�A(���0&"�$đ���"Ƌ �BM�Xd��I���$��$�#1�2F[���wn�RJFF�nu#cq�QI&*�ܺ5����!����k���E"�� ���"6+$����!k����c�W3(�cK���E@�X�	@I&1b����)2`K2��$��i�Khفd���\�JcK3�r"��#QI)����B5E�A��Dl�`H�b �II�"ų4�%��˻�uQ!I�'�*��>��^��:M�w�v+H�yo���]>��ɲ]-�S�o��-Ax�ѷ�3piG��{u������=q٪ce.A~ ��U��M�l,����-m<������j�����W�tn�F�3�nJ��:���P.��,9�AjMּm`v_`����HbJ5R�]�^�l�,"a�4I~�	��K#��}��;O�V��*�1v��\!4ڹx�J�zo�-�I/ʚ��a���XzWc�o�QyY�=�@�8���j��3��%<ՎΈ����zZ�e��q��͋<k# /"��f�� �aZ�U�#�5���u���Rw!�:�/N�-�mn0=18�T��'�Ё���].{��]!�Ys�}jƫ���˻��!h&�)�OҩɈG�9s��V\�m��wvc+oTAT�?�G�;6lÿ�Q���q?r�R:���ڤ������ɾ:��wns]5�~״s�{��ݜ��BJ<�Z.
]�j��A�]L�%�_vŌ�lmY����!���Ke{�8	`�t���&�W.���yX��q1[��g�i�n�Kzy/�k�x���g��Zg5Ӳ�:�ˊ(x`��i�#�-�,/-��[/�N J�Y�_Nǅ�A̾��W��C��ԓ��F���������V5m�Y��g�0�ޱ=T��ّ2E��#�)�����6n�"z1��t�o9Z�=�7�I�c2S6E�ڋ;s�ܧ}#1��Of��'yK9�ݱ,Ѝ�`Q����U�F�<�����s<�E|�
|�d���c^mn��
�e]eo:/��M)���͈H#�	��	1�J,b���oI���ֺ�\�	Y��;3ۃ�u+���7��?Q�k�P�	E��i����[�U��{<���c�c���U���P9��tئ
����� �xi�� ��lZ�V�Y��ϊ[e����Y�4'��ީ;�+z�랚�K��D���
�#6S9�8{�z�M�	X���a�.	�S���؋����Yz�ߓ�΁�oXzgm;o�!�^*���K�Y�uܺ*"���{���{	ǖ��{����O'^,u�!Cb�H����z��ǚ�k54{k^W]��%d�޷q<O�V�����!�S����<F+t�<]L���h0'X���5��u��I�{���姕����*P�]^�'���v^` <=��/��a���%ƭR%F3���랰ګ�uך�@��g�$�	�@�{X�H)��2{>�w�XI�����9݋�o���V��;Dr������6�&\�Eo��J��n���.l&�0��*pJS�qQ�/��[�9Y�����Υ��մ;�+�)8��yQ�����»�Uz��}�4�:((5�H�z;*Q��I�^�=V��mk�DOA[�g!j��m���bz�u�9��5��u_�=ۥ���VD��k-��{��w��&��Þ��c?{��x�/�e��ګK���mX��=���u=L��gz֮���~"g+>)���:��ڝ�f���L3��=�tT��NOk|����#ơ8Yy*�)�-���|iMB1�N��A�))�g+[�ݹX#�J��oP5�x�X�����@-Ŗ�z�ŽDU��Gn���M��Z�"�@��ok�fZ=W4�������[No�Գ�э�2��\ľݾ^���L�h	z=8:���y/�]�*b'�a;۔�wJ�c�řw7n�1"��z�N��t�:�}��y)�c�6j�����إR�4[M��M�>['=yؕ��V*Y�H#~��pF�gFv���+��F��lV��q�}���ki嘃^�k�%L�L���<�����ܞ%�ٲÒqt7�к��}�V��aX�*�!�>�ϵg��˭X���e�Ch����3U�mZ�� �K�!w��O�K�':Ǝ]�e��8x*9��[u�ʔI
u���M���اjD2;W
���j��:����jGL*93X.�ڭS'-����*�����~s��'k�A�Q���~5+�t3^;Э"�a툎9Q��v�w:tw9�s*�ps�tW��W*�٘F����ՊGj����9�r�����e[U��uK)8x!��<�&0Pk�2��e	]�F%k�9�sq�*
�	�;�mB��'㨥RV���c����4Pk&M���	e\��5�<LE�����׵��F�=Gw��B�B�����]�}	�
ꁬ'�dz�78�c�b��}@��`�e ���k�����f�e	s���䪻��])DX8���z\\�Kۗ)ҽ�t9b=���c�����ZV2w��  w�T��6�}Xv�-=�8^�,%�`\ë{n�u�cf�#I��v�P"h�hrlF��v+���]^�(2�c�y�:�]�����ʗ=�OT������Fu��?L��j+t��W�T�t��z�^ֽW� u�%�u}^�6j�\���imP�ʜ��A��OINs��C|1R�b��4�8��#<���S���ˤ��M�+r�S��.�K7��Rw
���N:�k�l�u&�<mc���mt��7k~�d,�s�I����׫Ԏ��h*�RX#������3�������[F�t�(s�W���]��j�JV*YJ�ta-�f��sҷ�l�������sr���hD��a�A��O	�=+%<X����\�ӹ��q,֗�9�ok
�d_2����õ�G��8�Y�]G_:T��R��$��Q���I5yW=��Y:��n�q�<��#�]f^��ϮUɐ�t�ß"�{����`��+��p"���n獤�1�[�L��:�V<בC�y���*�9*s��e�J@y����b�=�s�k�*�W��[�M罘��Ȥ3����*���+!���_ �y���E���v�Ī�|�@���~��D�=��9vOoU�^�ᗉ.	r�C�9)�����B�=�z���T��%geS�[W�Q�
�.m6a��Ƽ
n'��G��{���<9�3+�7^�Lg?F]I[V%�z���z�U$-N*�ls�5�����r��&�Id9�Xk�-��v+��Z�m׋��Z¥N���R/7�ȴ��oM۾�<�U[�-�z��;X��v�u�u{�N��w��
��Y�kh�)�՛x���]9���I���b7a���V>�R��{�L�{g�V$�^h+�X�O`���������ih��؃=��"�&�Ω��H+��7�"}��%�3ʞ��w�ߵ������[8ӫ����9�8��:t��f�k�P�Qn�[M���O.�W�%�%��±I��d9Ǳ �=�-PY �JE����S4��z�zЂa�n�Js	<=ه֚�v3��~۷������cu�ʐg�3��ӍɈ:�י��vމ�t'�+:���#�j�=��vR���!ITJ�ʉ˨�{��L)�^�a-��ȍ�Y�a��
����#���xL�l�ޘ�$�fBƣ/Zb�{��1��1��!�0N��V�������	���.c���sV�՛e�XM>�m�d#�	�0LW��b��ŧ�ۼ��hܺ���z�/��]����Gy��zgo��x:v��UO	���"�h'�������X�W���Z��H�S����E��z�ګn���T��o�A�8�N��
��\B�;Ь�A�6�2�|-�:9ԕ˻�"y�+e��7&�@��].��BuᇥZE�l�P��;Ջ�f��<�4n��پ�����f�G]J�V3�z�Vg�:��qP���I�E��=9����sJ�TS-�8�c���"ٰ#�*�D�gyb��^����4��rAn��́��)�;����4Pf �j덾>��#���՗1���Vxu.�s��{�,�c�B�쳅��S�Y� =��+a�:ﵬR���t�c 7���n���ھ�3't	m��ضWN"c`�ᠠ3wb�Y;K �ۥ
慭W�S)�oz��9
{٫���T<�sꊜՒ�~�����B��V�L+�Ϗmn^"er�7��7\]�^����F2{ۘ��Ca
��6PZ�ms���|/o�&��OZʟ^/er�� 
���RT�o���KK"���M�V�'��H���J��	OQО��C;�n�*��ud3r�����^m,��ݹYQ<lS��A�P4#P�Yc6t\c�����D%w���g�Z�>[&�	�++�<��,����E�$���Cl`$���,���L&������&��Y�4�B$�$蠖ܣs�tuxUz��o!��;�w��C{��>M=2�����F!P��Q%w�V�'���P6i���	J�Q����^3�6zvp ���"�9jj����++lW76�N)�{[�/\箺���0�j�#2z�%���-*�g��넅��d.�=�4�������S%�֓���M[\�}y�x��t���	N`�%L!�k�{�������6�*�C���w�-�-]z�/��%b2�&>�/9��/+��2��zS�3�6�����7{���6��»�MA���jD�v�f'#�`�gla��U}�RS��i ���G��naL-�F��,Ԯy���U7��)�i�xF�V�n&�:��:�ȞV��J5�v�T��)��;AVU�<ڶ��+-8]V�i��I��d81�sfY��TxL��Ѽ��j����X�j�ׇV>&��
�ls�5�9�ɓ'��yn�gs�R�Ue;��-+c����{�)k��-��Z	wع�Oiַ:��^��jݜ�lD�1ȉ|�δ�!���±�[~��^�(2�Lsa\�;�s�[���Jk&����V����0=���M�b�:&���$�E����u���\^J�<����ծ���b�ݱ+(eX���HzW�^-��,���x_�T�v7^�9İU4֊yݍ�>]'�bV�"�"�66x��j�v$��́�D�!�Rn��S�����F �[uU��4rкQ�w��d�Wg&����Qz82ǃB��yy�/?Qo&�l�I�g��u�i�1i>pSܸ��DV� ��p��ِV���y�0�odk�m :mk��n�m ��b�;�}3oBA��iCm:�m`K0����gm�<8��[�Ͼ���S�Z}����a��
�.��z9��>��=�3��}�VJcu4��.N�V2��0�vJ`�GT�eX�J�YXT�-�a��B�qq��9ek�ӑّSjnwy�Z�t�;^*����ұRS��m_�#�Z�7JT}r��|7ږ#����r�[�Գ�v�R8%�,��.�}�RGr�������i��Xt�q���&z/��m��P��#P8�t"9�eLa�X���3�8���Q��#�w �.G��u��K�a�V����ݪ��b��e:+j�:�+6flk�e.�������A�JL�t}�����Ւ{j�=�Y��V�l-N)�5�WWfW!�E�f�Vf��h�n�͈�wGv�k���^,�����+��$�sŇ�by)��1�|����"���=���1R��^وQ��X���/���L��ݵ����:_1[s�7632���>��QZ�B�`s�Ms�Z�L�zw$��]ޱӬ��M7Ή���rtt�o3�Ql�nz84��A��d�#��Ɗ�RGV�Ӫ�"��K������rb�P�oy����v��)�tni��}O"s
݁�99�B�X�2�� 9�+vw�Y}���{|���f��J�MpYա�q�)mf�Z&�� x��v�A��ý�@�׫,F{�D��z8��h��7o���h뜈2�2[��l��� \�F��n��V���n�ʧ�W1��tk>u/��v�_rJ�_NV7,�xL��X��k~Q��oU>0�,2urW3T�@��ҟY���6�)x�J��3��kgJ���F<n�LLݦW8�^ӫ	��8hu�	����!��wW��6mK�F��1���aI�˽zB�]{V�3ETޓ�38��u�(��z��H�R��lf�@λ
��]����c���v����j�г�^�>�J��-�ۇno[((�(jXph:w%��jؒ@��E��^��fހ�6��J�\C\�$�	��zfY�AN���mkzw�jd�5}-i��_?��gm�����Q�1]:���=
�sG����K(�o�N1��J����	^�l����Tс���g����sW.}�A�h��0(�4.�e�8�2�З��U9Z7ΘspP��ݜ@�3 ��"�x�:�bYq�C$�L[M��5^����*�.��t�`�U�8�-5�D�xwp�e7��
j9���U�D����$�����Ћ��ő�yh�
r��3�nd����曅��n���57�\z��PV&��t Z,�@P`��:^���\��9qŸ�K���~��8�^>���k@VݼR����V�h��Y/��X}[��r`<��!��~|���Kz3d�WwoL3ׂ�5�y,2kiv=&�'k�b�L�XyS��N�v�!U��;5�/N(�tB�1
c��o��8̮0�����k�kr���[���g�t��-���m�"�/p. ga˙��y��\���ub�#V�cP����2����,iE�}���%���۶Š]�uϕ�m򾒳�{SYբ�:��H�Y|9��fN���@`���}:�xE�7�9�:���rƂ�@�D���^u�w&���f�Hp��5��n��������&a[:��bP�7ot�Gu rM�Z@|g�*ZV~��g�Ѽ�}YJ� [���g
ۭ���f�a�e9P�Ք�=LMn�2p�
���2�z��4� 8��Ё��[���x��ww�������d>���ZL{�.��T�Llpn}y������c���v1e����.��7��y�DN��o��QXvP���^�gU��!���� �C��(.��Q�E*;4\x9�Ʒ:�N����X(�_Α!�"*4��VM�.����T��ws;��A[�$Ȍ̤�IK�B�Qr�jB�#hH �F�E�rX�TL62m��1�4	�%����E%-&�#j2bJK	��"�ݘ1%E�s3K��QD������dŎ\�6�A9��F�.�D*BɌQ�D���[bX�5��IF��"K�i����Z1���$КL�	QPcF�%nnEL��CE�Ɔb1�,Y(!�1�h��Dd5�6��Y4cb�5 �iB,�)(-Ԃ�lQI�II�a*BfĘ��BAR�(UT�jY���HsW�����n�͠j�k��rfu��G�*#i����%
���+�Xp ��.+�m��V�C�����V�ڦ9���Ҥ��1�=���u@'yK1��@F�+-6�p���[ث�3��7�E���;C��Y�4�0��/��϶��6�<�7lJΌ�sFÚ�+����.Z��.���q�z��F ��T��8_ֹj��G� ��v��n�X�� s��n�fǣX6#P��u����gz��٪�KI�<U��y���qZ���WR���*����#�����^v�l3��z�~��E9���ڌ,N�~��D8�FS����>��y5��ɷc���=�����zj�N�ai�i�	X�t�+�1
����iLލ��=6���7�OaT5��a�ڿJOKƹcy��'m�Nð�TpRt��\�Dp��yS
�1Ѭ��_W*D��<�l=s���_��f��Gk����f���zu�"0��}��I4���7���[o�3}v�J*�Z�_��u9�e�oHl[Akh�g��V��vWɓ�)��Uo4B�X:cpx�v��]e'�8�>�6��sX�L�N���Q��4$��2*2b���[���w�����]jV�}��� H�]��ƒ[{�Wkv�E%�KU�4��Z�����<��G=N!V�}*���zO��W�]����;�KB i���J�G��M�����v�!���8�+ߌ�7u�\�靫���'�#<�mı��^�ڊ���tW���99�G\#�څZ�4F]K�fӅ��'x�sx�s`&���[c��C���\7V9<����T%޾��+�廕kI�p.a��u����k0b6V���5w�ͨ����\�~���Y�kW{5k��Kc<
|�3N�5������QA\C� ����kcv�=�k�++d�=�H���TX�)�:Mɽٸ3���է��O]�^mv-��������ؤ�@ЍA��I�鵛���:hv���u��݁=V-���	�YB'�Գb�D�����Y��6����pȡ�Cu�4�y�}�����b,עJ��P�׊t���o������V���kW2���D%; VF]�n�k0gF��\��LA����jV�Ug�]�D�w�]��x)MPy���j��3ncJ����Y�:<�����EXU�w8bqEmZ��{�����]�cX����+��_}�����3�KA�Uryj��G7���@>�֚}�����W�b��kQ�vp��ʷ8�0��0�Ԓ�bڰ�=�Xk��������·�DC�{s�)Ű��ڣ��,P�����\ܩD�)�y�γ��@�Ox�팹��[*����6�٨K�t��	
�L�B�{�M,<�⺶"ɥ��:\[����;�i9�naL-�H��J��guL^u�G�5���fW��˗w\"�+G�r'���*���z:�s�X:sR�X�m�3��;���77䓆�XI��xK�fė�����8���Q��&nz��ך=x
W6��W���Nh�4MWFCn$H�8�YK�g��o@��t��[W��	w˘t�ۮ�7�xb��ݙ�X��d�^�Ԇ�W�M��t���.�o��'o:^���"�Ț��F����Aݢ��(���ՌkTo/&�l��������M)�4L�1]$9�x4PT�� ����!G�4�R1e^�C�+U�����ηC_riM����Qی�ݳ�fmn�.J.��%�D2��.4�B��� U�Nw�������GN�*�b��S������9q�e�3�nr�u��5a���u[[G�\�.)ni�.�=m��j�c^mv{�cv�%ezV(���#{��R���[�r{�΅&.J,g�4������;=W�VDU��6 �������q��sے�+�+�Rn��X��J�m��'$�M�Zev��ļ������0R�Hkv��5�q�|��7':8Q�ն�{y1��Y)�k�xH�Uԥ~�e+�ф��f�VtV�S�ѕ�qE���Ⱦe7��Z�t�%�O	�+���epnh˓[�;�'���y���|Y�cz���ۻI�C��H鄅Gjn2�l��9�"���	n�K��M'�O�=�ƺ�Z%T+��4 r�s5%H�WY��
����;���Vi`r�<s�,6�9�Z%S� .�1�����ں.��ci7��[vϷ0&����o4�Yy�`P��h��=��>�Y����e��Į�
U�VR1�*gݓ �G�gT�z:�,��8�v���1tQ+�t�co-�Zέ�S:�u�FVwb�W|�K�Ԉ�C�U�#f2�	MNLV��4�����tW⋛M�y�x��v�E��#A"03��j��#׆�Bځ꒽�Q<�k���
W6�8���ʹ0�U���u�����Q��hS����إ��f�׊]���F ������ua��u��Mh�1����oԶ5 97#R�˵\�d��w���&s�������.�!�uZ[���3ʏop�{e*�784;%:N6�����$��3���<�~kW��yZP�xn��J�Īe��#[�Y[t�Pl�]p����<�|�D��z�%�黴��8����1y�%`�r���lF�F���[�i�q�'r�_E����ѵ�y��QK9�['��R�z'���l
@�R�Ʊ�`J���#Iqg�N�5W�9��SO�V�G%f ����&��g��^��$�=�yY�U�:����ވ����;3�����U�=*  �_n;r��)d�}39�J�(��N�ÒV���5�Mq�Ƒ;oc����D�⮟;���:���3����ø����z��<��0����[��,;ز`�=�#�L����Gf����a�^�Zi�+Ν��B��Vp����Wy&XW�<������ւO;��GG1�a�N�=;׊�i@�ף��n��G��p�8v(G&k!q�ԥw%:�7�cq��v�1�w#��wF���:D(Z�zW��+I�����;���לtD@tgx��q��ϫ�t�H������j'��p9L�V.pF�qb��(�wCS��g$r
�ێ7�+@u#��v�T���QڽZv�9[��=I[U��ɛ���!69�
tW1��rxE�`GeJ;�s��>Dn���������z�,oL,���Û	�=e��5��B5s��̠(f���E�Շ��,GO�=3˘uom�cu�ͬ��0sxLC0u�m��[�aۍ�~�F�-��jw�ˤ��)�LӮ���;��*�1$�����s�yp��8�����U��O(|^׵�g���(�e�S����{g!:�������˕�Ν���v�L����r��k۷�mMH���m��Ŋ/��D���6X�:�<���-`�c�f�K3��=�m�}U=�u�/x�$�T�X�V����ۇ���!8Yy*���N�.By���.S�{������r�K�c5�Ҿ�V߳ض��65�v��9��
`�0��pi�F*(�{���d���2����Y�L�-E��.�V�J:�S���"��x&����Xl&��Y�0�D|�p��a,=}��^�U#��-ޟ>]Ս���}O�O�YDt�!N/jsp�S}�vv� ����[�j`��ŵaR{���f����f7�΅m�v�`5�7�/�s�o��T�HT4�
��:۫T�Q��sڛjlݨ�Н�Z�R����S��;^*���HP�L�]�{�*����vwe�ܬ�v-���y���m�K�;*�X����K�ꢮ�2�W;۝k-q��/a�s�w��EhV�!��OܭH�i��Ξ��$R���'���E�/��%<]����ʛ�>uٺ��s�;ӭKKh�Vq�N�Ʃ���i�&��I�����J��2�	D��w�����b�����nm���A¹�6�y3}�� ��V���f�"a����-��|nм��E�i6�N���[�q��U:r��h0���si'!����
c�>�2E�ܫ����k`�s�ʒ�r�ڱ�h�׀�l-aն�<1Pe6����>��t�^�@{{�b7�[��Z�9m^�,%�.aպ��q�Aڄ�=�j�n���Hlݎb&U�M�����m)�X� 7tր\C�x0#m�TT=Y��͡�S��ϻj�9|�fQ{#3�np��>���{��^u����'�M0*z���5s�y�����ʆT�F=��!��W�W%�!��Q���X�M5��wc|m��8/ �0�V�n,[��{S�� ��t��f��L�P:�t�6��P�b��i�m��n5	��\uK4"J��oԁK�!������2^�qWQ�mp�)��͊��r���)���eL%¥��eM{	lL�3kּ���N&��)S͜Ua�m̮�Z�1��
=mB�F���ٵna���Oo��"���GT\��}*K�m�lS�ӄ���˹X�3����aS����,�S�N����_e����(wn������Xd�큅�+�ׯ��z9�K�rV7}S��k��፞��k�T�&*V*Jd�.#b����ѼC3[�*r�n�������vûK�;�P��! gD���g�FE8��½��W��y�M'�HL�[�:�B�D�=Do"����ܚ(�����\���x�BI��t&!��oER$�^B�f���
/�.�ӥd���:�K��S�x²��	�61�Q�\��& �q�K�+����,�l�~��9�ڬ�,�ɿs�B��G(�����7�)s�Vr��M�8����]�+�l�v;wek�Yld��[�S�)�[��Kvwu����:��OXo��!���\�=6���W���H��#L$���b�5��e���9��N{\�����FgK9I�޶�L��F����0�k���v6���c�M-� ��4��F���b�����a�Cm���v�4�����Ǭ=K<���d�@l�]��7X	+����&:��ܻY}n�Y���6�E�"5ԕ��
ΫU��D��{mt�*1���[���k!۠�cy�']�Ѓ�&k#�v=4L�W����mr��6��2p�S�ܥ�l�ep]L��:�A���xq�9���)865	X����:ޒW�vb�`����Y����Y��;~��8�F�lF�lF�@�u��7n(Tfr�w��/Oj=����.��$��w0	F�yL3��V���KաG�N�s_tBǖCN)���֫M�;+�4e1��H���V�|����)E��W�=��5�5�֚}�V7��aXF!W��1v��tk|'F��,0)'RJ��mBO�y��L��;��}{t�uÞ�X^��ؑ�)��}JQ*1������`BȐ�uWO"�ei%�U�L%P���P���	
��d.�w�XI���z�K����.2�um^��.��~,�Sn�J�VB���}��g4���'}��dk��#�g�Wdb�W��T$�u�V��7�ԏ��FOA�)���+���xP����ug=.�Dˡ�koN1��x�����O��������B��<�Q#���n<=����Ο<N�'�_v���r�U{�
�C�0-��g|{[�9(��ҭ�{�"L�=��b��Q����S�w�/��]��ޠ��Y:$[)�ٻ��%�h+��}Ap<�.g/y*�,��՝�5.b�q"����̔R�B�3�+;���=
���%�f��d�z��4�Y���Zv��걨$�é�[�f�ʹRX�
,�PH3j<',mu�ذoS�nѡ��p=����~�2�e_/L`Q�'�H���t��,�9�̓7;wI,�P�#)�b�����2��G��$Vڔ���{Ǭ8��nk�$�2�Y[}>E���,��]Y�(*7WR���f7�bΜ��QVmٗ��Hj;�(@�E�ܐ4Ua9�6��X�X�h���n��C�u�Q��Zy�f��ĢU��ޤE��\+E�Xs�!%d�c��� ����v]�/�"�{ov�:J��]���܍g8/7w�eu�o�7�hoA���GK]��~V>�9�mX�J�Dz�q�1�;9�}�LuA%.,+&tۿ%�0��)|�<����ݽ�V�»FX�kr��t��¹�o;��OW]�H��K3.��5���3�M���PAx].[+Ar�0�!q,VλV�w^=�[[kf�Hv��ӄ���m ��'p"+8'L��2�*�}}�wώ���P]�\��k�T�P���ei�(��|�u�lT` Խ��bj�w���7�|.�3R�y�:y_`@;�-�<+wQ禵�ixY걼1�LD1�V��[�7��."U�3�<nH(j��w��x��j� 墷z�a�-@P��N��p,���L��n���]�K�Pl�;6P�+	�q�'��r��4⾤�:Q�Pt޾��kD��G�T��q��CK��>�Yp���`u��X�&�Q�qՅc����"i܍uJ99n�r��n#N����:��d��&�#����9���#n�'ͫi��z��ͨ�ȚV�W	Yѱ�rv���X�[�w���.`���Ҡ���y���MԲ���iX���}ו�����nΛg]cy��s�0��)�-Ԭ�X>{�<g�ܗr��;sj-���M���	��!��r9�&t�M�W�)�pg!N��tK;Ϡ��Rݰ��jTb�S��5�wC�1W��Z���!7{����l�/q>/7m��S�����nV9ʦ�!��Ǵ�3D�l!WX&Txn���t�V�]��9���i��4��
P�׷���wn��P��P�A>�n�UjtzD3$�����ѕБOj.�v��ic�v�g	��wi�o;�ܧ�޸W3OO7t�	"�����_�u��Ƙ�-d;�-�:��7z���ul@�yO�8f5�����rWk;��2�f�*	j�[+뙦�#�-L�H&�3B�FR�!��=�3�4@���C����_ޗ�������*McF1`��h�$b���e�sc	#E�JVTR@X�lC)"HF$1F���B��� ƃFc0cPı	IA�R�h��rM��r�0�4QF5�4�" &R$F��1���MDj��!�ѣ2Ƨw1�hƋb�%d�E��k�5&�b�b�(0bFǾ�-snc	�эF�<nIE�*5@�2,�lh�QQd�F�F-%d�Y�%x�wksbyڹbLF�lms��Rh�D�@@�cE&�lD�Bj#��&ō�
,�F
&a"���h��A����]lȘ���\lm����]��tu,k&{Wҹ覯��p/�9^(�T�z��6�o�T�ٜ��ts	��Ox�����(5�H�{��b�w>���d�^�P���+VՍ;G�RV�������0o��%Vt�aWl%�磌�[��.�{���Z� 廕kA4��:��뱺�w���NM�yqVG'�^ְ��F�g�ln����`ilg�|�A͚��3����v�e|��8�F+Khq���BU��R3�ٻZq�x��$]<(���8�u�~��8�c^mvyln���x��lR�tN�ї�Tl�r��X�%�����v�[�r�	�b9di#'�ޭ�̂vS$�����9��Cu��]�V�S>�vS
���u�j�OcA�����R����������C�M>�J»���=�ܵ�l���0���,	�>�]ԥu$��ŵj��B�_ءz��;(�`�Q&��P �'���7J�ѹE�c�pHo�*zr1��9��q�<5�N��5m�ޮ�"�tU�Z �.�6[P��:w�Z�͜�QV��9yb-����僕��/��+n�W]3�gu6/�\殺o�;)cj�����%���g=Ӱ�x��HX�������X
�%�%E���o�X��֦��[���C�/BGO�!^�L�\�_\�k�����Ȉ��[Iu��镐���;�a�=~�͉U
��F��4W7rUj5�:��*�����
�-8fu���E�ՉT���#�N�är�%!��ޚH]�]�?R[Z�0�5<Nlk>S��c=�&#����uS���y�U0��[8#Hw�5�#���90��>ٻ����}���;s�Һ��`���'&M�����V=������<jOkm÷�uzG�������킶��ZL�,l�1�c6#uX�{~������$[A��3t>x��P�4g(�^�>�����ˎp3��fq��/^0�i�@��f{��唫�X[�0��S׍�vxj�z�k���
�^n�IG��!,����a�̇xk���ޑ^$/k�X[�V�;�7�9��I�P���_:^^U�s.��	�5�d�}P��$s�M��
�x��K���&�.�,s!I�]^�.��٫���H=�(������kq��'H�q��(-�059uB��}��ߗP��^�,���k]�sxH|�NTY0q8K��s֬�2#u�^P�&�:7L#cf���(I�v�A�}��ԋ�p^i����ʻ����f Дk�%X�f��u%����o:̘�U��P��a��Ӝշ�%aY��h��bS	mK+:�J���pt��>�k�6i}�r���!�]�ַ�p��)�"	�ҹ[;4��+�[���W�o������s��X�wig��5�GNე�+{~�998��g�wP;ص7M,���g���m����C�Q��^L��?m�j/Ӿ�M].{���
�M ن��m��.��b���R�U�L	U�`t�79s��m^�x�⋛M�q]��l�ƈ�릲˭@�cSS�+v��/Ҟ�f�w�.+���_R���5��Q0��ď}G�N���;@�u5�2Jlh�J+
���Eƫp��Y��5�i�^W֐A4�(t�� E�g�2��VҽZ0>,�����1U�Ό���R��l���B�X�nJf��˟Go�Wb���.w�	=S-s}|�쩢L�V�딑�a�9���1���K"�o@��~�������r�:k��Y�_4�J��aՇ�O[u��l�1���U��8D$�shVf4�lQQ��B��`&�g�1�\�㮨'yK9��P�ɡ����n>��Ԓ�u�����lf�P���$��<�1|���gI���mӽC�X}U�7o��P�������8Q���X�*{ڎA��`w���W���݋�wb+ ��ʉ�b��7������b��ԓ�ݾ��wVu;e�󳽀�V�l��a<�T�(1�N�p���Δ�VD�&o����OL穧�p����bp��q*u�ug\Vtb����\��Uڛ��0���XM>�X�Ӱ�#��:Ȋ��h����KÈ��8���j`���$�z���o[�;iｩ�W
���u�C2ޝ��|Sj�:��e�I�bnp���J򧟺��.��Ƥ)m��Df�yOj��+�����c���}4�<u���Z��]wu��G�ۇ�}M�v�uͰЗ���Ӥ��"є�WF�|3$��݀���=3��D�Y(�v7�����D(Gk.�}V"qN��=b�;����yݪ����*��ۦf��!������+I�����k�^�:\[����;�����/J�Vj�>��].��!8��]U/85�l�D�]v��j̬Q��rZ�h.��z8�mA})����ۦ���n�V�7u��3��;G�+(�ߊN*�c���`jܞ�d���3OWM��8�۸��b�ڽ[^=x�����:�&���]o1���/�8�Χ3JE��i5��E��Ѻ��O_r���	��0���u�]��1R,#g��:�W���Nf���9V�Ϧ�\��V��{V>t&r��[!LUgwN�.�1��Wj�N�}�.���z������w�$C7PA������\R���]"0OYО�����V3�+Kj������>�s�Ŗ�\��r��<4Ln�C��}.�֑�r��tp��3�:[A�j+ e����sJ�C]KY��sF�:����֡��T)mc)5-��{\,������5s[���Y�;ќ�EX!��2��{ϴ&�r��@��{�����y \Zc�s�wz+����p5EQcs��vy=O�I7�K=+���7���F��˫g/#�-ߣi��aP��g<��*�i��8��G^n�&t�Sy�J��JV*I��R�H�7������4��ǒ(¼���V�B%_�;F!��T�Z*Iy�j�'�r���6��f;E����~I��V�t�+^*���B�+�[}m��(�L��N�.���r��yr��v�+2�o��ԍ�$TqF����|��!�}�ؽ{�J�[��E�i!y�wb�s�N�ߥT+�wUka�=h�b�nq0«�u��B5��ZE�r�<�p�`N�)T�`ݬzX׆(u�5vx�gf+X��IT��}���
�F���p�Cc�9���Җ@�{�1xmSD�?z�*5��(k���<��v�x�5)k��P<�������4ueȞ�KB��+x�F����[#W$­B�y��TW��-��H*�i|�$�b�',Q����Av��n$1<�y�s#�M yV����P�>Z��t�E �$��Bɋ��627JYC����7i�%�������:�G��·���na�M9��b��U��"����V�ny-�^g�|�f��J�w޶��ES�x�u0�_^$B���ss���������|g��.�s��	�	�S_5�仾a;=Vp)�xS������ƾ��P^��ᕙ����_wVLl��k���)�N6�7������������{N>6M�t�!�ξ��eܘ42�\ZwY[~�ޡ'Q�YaKL��;��0g����V�g2�����d�/#M�yQ<�S�t�7�L�@�-Sx���\b��MP�y�I�ܸ�Xl4�NxY�5(�IWR͊@�]I`��m�7s:��z�1��vbp��8�>�XV�h��D2�ږV�l���f�᫼�ITve.�]�}��]�u��r�x�� �=��Z2�]�3����b����mX���֎����ۻK s����:��Z���z�yRY�r(�k�,�t�|Ab�߄��^˼}�;=o�O����U�R2e;�ŝK\U���k����㱥�来��=O�q���=�g��)d� �-B�Uw��g��	��3@W�~�(�	�o�ݽ�3�Y�ی���Si�s��?v*53X!q����K��ڙ���ۻu�$�)8�EU%�8�k���0_U�K��x�B��A�C��UG�t�>{G�������D0�X��6�>�˝].ڽL�W9��7qJ.$ƚ#�N+9P�64����^��LC=u�]�t����[���Yw�C%�V�����ls���ٍ�K �f�أ������+���R������K�0qw�|Xz���[|���x�Tb�(J[�S]���:��=�]���^���Y|�9b�v�O)����R�vwIV�B-9Z7\���6�	��	4�0�<�&�C��]��X�.��ksX/6�lnؗ���em�N��
1rY~�VEdb��6:zK�w���='\u��Ld��|k�yk���b�["��E+^[Z�W���]>R�!�Iʓ۽]�d��o�#�^Y^��l�VƲ�¯܊w��%��&k[���;���1<���`T�Q.l�u���Y�l�')�X
�ueKc:XNu��$5wN(E@_!uh��������G��ś�s�����ũ*�8�^L��m���/U�['=f ץ�O+�A��s��.�K�]^�[i����I����R�I��K+XU�����A��Pb<��� ����k��w�%�ҖR����0�氺��}����N�哋��������n��pF!09uI�Wֶ�'��<���L�sԜ0L�D-ݞ�*���;>.����h�}\;:C�z1�f�^��*���S�|�V�1�ڦ��0���ޅ��	��%nYt��8��a���L{�8̎��B�Zj��L����rbY*�n�ff�m�ats�f�\�	�=<�	ۍ��sfa��^`�ޅ7n�%�P��ʩ��ƽ�ܡߊ76RqW���N��
c�)[���G]��MԖ V��R�징�V��Ş��mk�ɱ<\�˪t"�D�^W���=��� �p��Ư6�������n˔�.¥�}V]L=r��,>7yr�O���M���@��L��p���.7ݥa}�K�;5��ɂ$��<3p���l�*���u��J�W@�5`ڑ�uL��E��ã� AIw�ԩ˵�^{_Z�t�oԵ�[{V�����:1J��T���2�;~�o��Y�叺Z��(OmΩ��=�+9OՕ�C6�r[��*���*��՛�6��4�_m�<��;��YP�X���E��!�u�Pkv�]g0�悷��M1S�w��9�^�כ]�Ig�����g?t�i�_�VN�������hF�@�X�EV��'�׻�EX��*�ГX��b]������C7��g=�*��i�E�)����ץ?R���&��ٖ����El�;��$�}U,r�YtY����[8��s���R�Ly�A���4�7K�VWϴ�n�J�������ة��C��-ӿ�]��>��1�V����&��H��1u���z��9M}'@�	T
R7FB�.�}c#��z��M�з+�Su׼rϙ�-��{��r=t�ћ��f��qU2����_]g~����C�m�h�K��u�mG{��VM�z�I��x� %e���a.� wFb��J���u� ����
JV��s�M��#�l}�BA7#GA{�ή��L��Mt�eWb�H!����M�K�K��8C�4��b�e=Y��g>��;��F��a>7������T��oP��P?*<fQ꽵u;����IHe�a��nվc6\J�1�3/�m�U�pR�B�c��n�&�!��-XT{h�v����,u|�^`���H�t��gu��$���z"��̧n�Yk�7�b���=���u�;5k�/�U�<tVws�WJ���!u\���XY�`ǡ1ڣ	p�:��I櫨n��k
��g[v%a�%�Q�U��Wv��+maޫ�xM�:�2�m�Y�Mĥ��
ݚ7N@z�w�:���d1�1ٜu�v^m[y�Ef�"ŋ���e��������j�V�[����k��<%�V��+�s��az�]�ifꈱ���;R�PL
�9eu��G'�,������é��͘�Wl�	&�)Q\;�&�2L����3sАwP[⦨M������]��w���+[�A�����YG���FN�����VE�4�v-�wlv��.�C��q��O��镣��K����δ�	�:z�*6�뼕h�cnas7�WcFYf]n�Awu�v�|�Ѐ��;f����H���������T;�Z5h�s�ho�-Q�
�c(��Ŵ{��O�n�L�,����>"f�A�8�{v�����n��M}��H�;��Z���foj
�Y�`�t�d���(s�]˩M�x3����&��Id[�Q�dNk��)�
�evgJl_wZN�G�XX�г���/�2S�6��շ;ܗ�7�0�`]�q��Z��b����t��I�=��su�&�meE���BX�V�����d�l�R��+��Tw*9T�Vl��f���Te��i�v�w}�ս�u��I}��['��pe,��4�^J�Z�ΌfX����K�[FkW�V�֮7���vo���bu��Ӽ�5��NRN��<�a��M�{�����.rJrG��e��r�e��wP�^9|�8�-w1#�htJ�{@����E��{���r%�Po��ݵ��NJ7����v&�R�Hf��b��l�2�[E���{��l�h��κ�D��������Uj>Ż�L\q�S�m�ǙҺe۬Ed1��о�Xo�ԫ�z`���3��kw��4�)ԯ���4K��������߄4����Wg�Ȳn��ﺬ�%Ëі���^�-�O��{���Rfc��2���T�:i����$6��<�a��6P���]���}RX��`r�E��h��������JG;�Ŵ��Gt�ۈU��;3p���sx�dw@�r�Г�\���L�}��M�z�ݣ�Ie;0����|�V����Z�h:wp�ܰ��6`5�v�>�oN�Co�29T�b�-QI���h�dV5�n_�\f��b�Z"LQl�	�Eh��6KL��QQcb����IF�cb4j,Z�ܱ�"�Z0h�E��*Ɂ6��2��#�1�1d**(�j]���	G7J4^5rw^/$J5�0TF�����Fk�" &�@�QQD�Q1	�I�L��F�!�4lQD&��j-�DX�mj,DP0R���EE@��3H(�1BcY"��1 ɫ�RT�����1{$�I���ʍ��
�z�hn����uEaz���m����ó���r��ޫ�@_	�]���oA](.,!�s��
�.�b�5?�.6c�w�6c>/�mC������몦hzUQF�H\�ϩ,+�h\���Q�
p��Ҹ�" ;;jBKi���,�q����
�<wS��a@LW�ϬoJR\G�H{p'l�K�Td.ɯG�Q��Bˮ�ZJ�/>X��=썲X�1�uz�h9�\�NO��\n�A[>�都}W��Q��lg%W%���
UJ;�Z�tʭ,�	�Ob3C׮=p*;����{~����w��h��U�`� ^��Q�J6�vk�p�k��1ǚj�N|��������wCo�t=3w�� �Kp=>
rXɲlv�����	�mG=�p�>�~��[=4�c98�e����������k�~ ��?������ǉȋ�9{��� �ܜ����+�!�=\�}
���̏{c�����~��89�X�v��Wtb$ָ3(K���+&�e�lz��\�O>y"SNW��ً�D9][c��R�����')Ό�'����Pgj�:�7J@]x�; yP�yRnk*�^��7����1��4�����W{(*����͓
��^�Fƨ���������:��lX�"��A�I:�z�s� ���L�nΫtt�&i*�a��xrR�}�]WB�w0�f�C}-MȎ�R�d�7�7M��V;�Yy!-�5F�a7����|kh�[�=r'</'cz���w��Y|-���<I�Q%q�3�
⌾7E@�n� �{���>}�զ����՞D�X���>��ڦ7!V_�6rJ���$�}3�H}P������5G�'n:�n�����fD����ϵ�ei�{%~����y���pT 9lA�;���^w�F�{&�6���|
Ja�T�79�,U�W)_�^v��'���O���0��}E�w�퉧�S�m4������}�
�=)t�@(m}�w��tա�}�Ƨ;�y��O��{�a��l��.{�:}�(�� .��<�h�QZ_����n���5han��S�A�ˑ��#6]Vu�}Z�0�[8M��q*���%q�@:������=P����P���nL�ʍog.v⹏xr��y%%<B� ��F�
���%M���L��gf�J��)������r�7����h/3��{�ƕܛ^�ɣm�^}�[�>"��X)�r�X���ak�^`��|F)�ǁ�g�S��vb�u.���{⾻��✛��p'm���t<f��k�Oo��/~#��J�?�d)�a���]���k�l��T��}��İF��
�;��Ϙ�{A���{p�[��y���*��|�U��/6S\�3�
�"c���+8�+�W�n�E��V������	(L<k�ee��JpSN�{F˲@�
ޥ�t���̒��0b���\��'�[������^u���V�}�Or<��9Q�4��G��^O�=F6�E/!�0r_Gw�kx���O�fau	��+����O��� =�m��~#�=rlG��}�u��;^�4��W�C/����k����j����!�ݵ�u���=~� �]D"��ȯ5s�[��^%�)��\'����\:<�mȹ�xz�eaf;"�W��>5
�]�9�]��|�W2���)�Tg��b�V��\I=�2�A:�C�5~<{p��zb|G)kf�X5�
��(�q9L�E5p��;�=�(�_I��NϸϢ�=|b��ʟ^�|���qR��T�)�Y4Z׌xgσ�=��A������*��{�7��FS>��:�.(�c(���J��΁ �$T)����>X�Ĥ��#�����a�t��*�2���:��~��+w�}E�D@�Pf6�R��g�D��Q�{qW�����z���Gy����إ���q)��\/:�����m�( ��F���@�W�X&�Q�>@2U9�>��4nT/��7E��Fܲ���>�v�3��S�2hE[ݢ��A��1��S%=�p�������%˼TN"&&�*����tr�e`�Ρe.��;yD�SV� �wl�ƻ8V�u;�ꀅ4��޴�������'GIk��v�J��aq8���vXQ��o�s�-�rp�x3hӕTJRWM� l�N�W����D�X�Ӡ��Τ���f��h�v�[�'/�d3l�Ѝ`�c$\��&��_��U�=P݁y��WJs_ES��rsM�+ƯҼj7]�uT��΍	ˁ���W��a AՏ����ugwu������f�?�i��-�~��/�n7�T���:���;����=^���ڳ���O�g��Q�_wQ'���Y��*��P�ٺ�0Lq�w%���T��P�N��e�
Ux�f�uaV�FG��y졙��>�p>7ިWYO���||#.�#�ٛ�����~%�o���Lk/�X�ty�xZy^����>>%Y�[�^7�>�D�H"\�q����������%Ms b�^g��~����65��tc_T��{�N5D��hF&|$�UZ�q����7'���x�:�W���02;L�WQ�l'~F-�������eQ#r�^s��>�,e@3���L����z�zh>χ���;b���3���n�Y:|E�OO���>!�ӕq�X�eT�-sM��D�: �:����h�J{,_kty�Rvٻ��� �ɇdV��
����Ћ��Y�"�[�=�s�Nuuj�:%�O���PZ�"D3�T��� 19y�˸u�]�,���e6���,g���f���woL�;����L�Y�O��B�{��T��]HAp��C�-��Q��l\�ދ�����5Uc��+a�Ss�tF����ĕPf6 }0�"��n�xs*�TUκ��,�	�ד�Ck��՗�r9��y�M������v���>%" �$x	T
�9H΍�w�_�C7��
��fP+~9<g���x+�8�|�i�����~w#��ћn�o�qD�����^�k�z:m@�KgE0V��΅ʝ�c>s��s;�m�q;p��*���i����"�q	�{=��R��?��� �tкS����r]L �r��,�d��j=������Q�qֵ�՚��/fH혨����ޚ�A�v����ˮ�\$�����֌؍̚���;O"9���Xln�k-ɾ2K�qn���a��QL��=P�j;_��}�=V=�]à�v�5gO��m���v������\z�W���@����p+��{����xk�SU��R��Xv�v<�Ӽ�y�J�J� :)��܆��5�t�G%����T��x��FP�ĺ���m��f�;�!�V�I8�:��
e"���^�;����3qRܯX���V����'�Z���
;1�&��$�xwmFɭsT�8���hU��&�2`�}�]�!%e��4���Y�c#f�T�ˬ<�����՘����k��T�t���ެ��Dw���q�V�#�^Q��k9�ڦ+~�a���_�O�۟�S#����:����\���>���Jk�!�=\�B�~e�,����.Y�{�m�E�g��a�^.�>���ʈ��u�^7J@}q�@w�p#�Ϟ@�Tӕ��#����!|�W�~�-�۞9g	�3;0����R��ƨ1�ʀ�ʹ����f���9���1�٦�5����/��k�#��'�OA��We�r9��"al�i�K�n��+��v��c\@}]�i,�^w	��ST��_�6rJ��<	<N�q�B羚��%�/�D��8���LI��G�&���W��>�!���Gn��n9�2�4���)�<����C�*�n��@E��L\T�'9xU�W��>��k��I����خ��܇U�uk��Z���pO%��������� � <�k`7��C��϶��']��p�	t,5�VHkO��O�j�vh�� .���v��Ei~�0��ۄ!q	5h��n��ƕ�O�kJ:�$Fo|x ��g�����NTN�6ݝ�z>��6�#D��$�<��v����`�֫�D^�{^Sh����ma�BS�3���f��IJ������:�Z,Y������Uӟv�v��k4(�+���3���/�sQ-җ�,�ZS�}z���Y���ߠ9����xu�"��s<	+O4���B���{^�*���rw���5������>�&�u����<��k �����J�rG�)GT���s������{-`������\9��Qh��}�ʅ��Rw�)�E� y�5C������`t� ܱ��E�^�]�xƟu��3X�w�����`W���=��O<��t(ה���I�����;CwC��a�.8O��!��0Vow<�	��ɏz=>j_��ҟ�O~���t�\(�'C\��3�
O�~�MF׬D�d��Ow�;�����<���5C+�PlW����c��z��c�@���L}���&aH$f��p�#����g�2��UO�^����� ��erl�z+*�n(��< w�[��l���l��eW�Y%�\B�c�|߫�ds��q�h�E������Fv��)�q�^�K�;�WE��P�40�����\�����s.��&y��g��{���x\�I�Ixu��^��V���[w�����*I�0�r��l�*5�^w,�)��<u|�=ΗM9��!ۥx���{ƶ~pe~ݸ`�_U�j�6mrdd{��h�v:/kw��k];�p�\ݚ�q̫f�:�z�L�1*�Ig��IۅAL�pV��b����1V�\��V19���%.�Wwel]ݢ١�t�a ��>�N�6b2��51���{xf28�6�ȡT�p�/��ɠ��k�<1�t��΃;i���/���lƹ�Ά}fg�ug�@�wF9�>���P:�=Ā�G�S<9�Ş
N�ls�4{܉\�ND��W�q����9S�m[�y}E�Zf6�J�y��Uy^�k��kO�e(;����;tR���h8s��w�'\4���ԏ_��Ы�n���D ��č3�J�F���䝏uw�t:ț��<�2}]�3����p۴�g4�W����o�����j�U���%t��Kr�^�^�_D��\�����w���${<&�K�ɴ��,�m���F�
��"�VS�u�$�vG���j����,��V�R���ۮ�Wˮ����;4m9p5�5���q/�q9��ω�C#�W���}bwT���dR��W�C��w���w!y�u#+���B�=��n��	��+��(�A���*���zU?�0�g�n��t�g�ﷄ(�X��-�R�~w�.��,�
�.����_�]}@�|n�P����+����C���x�r�~=\VdT�،C*[�fZW��E�ܯf�q��}���T���ãf�p� ����mC0��<����ޯeE�os��}]�>�.�[�W;�K�o���켝�;\$�BK�IeM���b��Ȝ���C�]�Y
[]�{�N���z�eu�����K��FD�S�9ʘ�_L�^��<.��dt�\L�5�s�U�S8Y=q��/ѽJQqE2x�tŵJ��@R���u�ڠ^��U灇�]�]A(��?�>�oN�1���'�t���(�W���02;L�����D'~F8�{2Ѷ1�-^Ec<��Gvc�/�8O��2�@:Pʙ|e�h��}���
�9lV|�&zFv�2^z�J/e�Ws��C����.9�]3�g�=Fa�=HI=��R�,YtQ�Տnx��\�}S��%mg��W��<����;A��Y\}�(�h�%W�c`�(�F�����a�ʋb�g�����r}kk�.��N�s�n���"9�jw�@~6�Hĝ�>�>%_�@��N�?�b;/���F���7��0��/�d���QN+�9
g����ïH��і�Agb�M�$����Ɯ�z�X�;�=�xV���w��,�N�1�}��d�	�m�N�C��h_�����.r�S�s{�{�����6`}4.)N��X��ې��ar��8�|�UG�-UDA�F�]��L�Υ��.�T����;y>
Wj8�%{���u����H�+������7*o��{6�3����s���KEm��E��]��y��Q�ݗ�ɚ��]�T̏�]��SYAB�޼�VE:��ٳ���ͫ�x�V�q��\�ӓq�$>��혩[N��ޚ���뷬�.9u܄���y�k@�h�q��ڢS
X��7|�e��k-ɿ��/�ژϢV׼d&r�#��,)��\7c�ј����X�h�죘�j�M���Vݰ4���P:9�������������鯷����JݎT���Ts�>���5����;�ޜ�Z�E�����t6��������;��.��K�陓9ٳ��:�c�;�|o�3W�ۅ�=4�c98�e������{�p�N3^!׬���,�Lϱ����P�|=>
�r�����}�@V=�Cg��@�N��|��=��&Ñ<��N��o0i~��yU�F���~ʁ/��^7���@Oy_>w��m�M�Y��ga*�w�:��`�)d��z��}g	0���
\�� .����)�K�Ku>l��>�9�;�+�	�$���;�j���T����*J�Qz�]|U���,8l%1����y����W�T�����w	��ST��_�g$��OOT΁�}&:q�R*1�3����RpM��:jw5nc����z�/K�ls��[&��{�9��h���Vp;U��8Ӝ�Fiͣ�h�F�;ɵ��ޟ�Z!۫�J��{WNi����	L*�t�u.��{���䜢V�'c�{��J�Ow����Q�e�
)�Q����\�dm#W��*.����d�K^ތ<���t,V�RW�8`���ѯ^��Ư�����P��K�����	wu�/3�h�R�̂��MIt��W��C��Wa�P}SU�(�Б6�^sf�1rzz�[��&��2���'j8e3J�w��aUdԱ2���-��	e��cx��]��Գ�,K�k��eR��&����H�QS��p�g�N���:�׼7���佰�ե�S)V��j��W'�s�;d��;�{�f^�;�ųD7��X�6T���]W`�k_���Z�e���H�`�%KR b�֚��Ǜ��>�SM�·wzԭč��R��pU>�IT�uZ�Dt\���E��]t5�B��u��%�|��=RF����mhy�J��&+:˒DF� Y��c�b��)l���E�fb�7p~\�v�4̶݉i�}}��ιY79��ۗr2b�;7�<�_���^��I�Z��4ySa�������[u�J[8����ŵ72*��[I���\F藽��ޙ�By4f��3�Ю��q��I�m�G�YP����˚��Խ8.�����q�ӽ�*^R���V��WC	9b��wu]��Q=���řii�FB�V�x�Vխ��Enq�0�%f(:�]�p<*�� ���i�Q�i�s���2j'�t{�Jf�Zb�ࠦk�E�m��9��W:�wE�$t�Z�⩶���u�B�ٯeI(y�͈Px�p��Stl�(�$�S����k%�˨IB� ��������8�cn�h�m���i-g�Z\+r��Tf$��.�9�\���-<��X*Wv�u�Y���iY����W ��]����4=����G�=�W��ޤ#Չn���Q�!<ђ�U�6:�r,�Y��H�B�G!����gqY���b�5:��ۡ�.�A�V�K1g8��Jvv%��gg<�̫ժh�
Z���u��t��ʝ\ıX�z��n3��U��Ou�Em�#��]ne0�WS<���J�H0,i�6�VX��WLpdܸ�����Ω��;wxX������Ԩ�e��s���3^h��JJ�;��2�jQ6� �oVҕ!3�eT��u��vK��C{ЍgT��
z�=�l��hˣ
��Lb2�j:P&2�����p<��A����QL,���m*3o5q}(�b��%�&�Ҹ�+��fs��-R�4Y�Ν�c5&�j�1�v�u۸�F*7�kVPw�����5Ӵ'����#���%	�,ʖl�ˤ�,n��Z_`ڝ/6���ٛI��J_9��0�;e����lX,ևһ��z�����?w���ts�F4d���c��D[b�b5&KA��A V5�X�`�ڊ4h�#�b�IX�R$TKb(�(���K��lP�56��E7(��c-�Q�lEA�B��h.W5�S6B*b��sF$�6+�6���Fɶ1�D��\��X+ATj���ԅZ6��Dm P T��p�h����q��*���*����7�.s�\�`q#����:�v��\m.kv���B�*v�enQ�(F5v���-�2�_p�׿������US�ȫ2�o�JߎF��8�J;p��Y�e�F��QS]�ݣ���c�����6X4
jbI��V*�*�`؎Z�q��>;p��'�=���ѵ`��{��t�Y��Qq�@�Pd��H�Gg�M@Cv;��0�A9����t�m��s�݋����qˮ'��۸��T�G���~��ζ����"���n��b<�W33��]��Y�s��m���E_Ҫ��J㤍3�[N���՞�W�O�������'+z�-=
��rSs��0�#X'����V9���/��;6�����(up����g�Ч8��ߋ��^�y�ܛ��L�7�^#T=o����X)��g]_=��3=����_�'I~8=K��_�x�m��ȍ�w�3��97�.��wC�Q��Ԓ���Nl�Pv����aX{�'U��ǃѯ�pO����p�Q~���wS܏'#�}	W(�/mfO�zzW*S]����D����]a�� �z����S���R���Ԁ�ih�\V������G�>��+(�QJr�����÷�������G�3�@���z�x�}�_gVsr�Rs�C�Yu��J��]RȬ��9�b���!b��Lu#%�u�}/��6V[��S駆 C@S�"�[�;\/!���G�ݣդJ��{i�N�t&+rw�/�����Z�M�>�^ׅ�箇�O����,4_T+���)��s�9t5���fo�qX� �ozȹ�dgʩ�.�7�����y���d��U�}1��C�=���p;��=٧��O��Y���Tw*�]S�L��8k؅�U�xg��I�a��ò&�P�[Z��#�gB��jb�����l�*5����E�')�Ȧ��9�c��Z�f:*n�Y��1�9XH>ft	�BOOET�S�,�
�k�<2H{#΃;���؉=��xz��z�W�n�*�����,���%Q�q"˔��L��,Y�B�'~��2��B˓<�m�xu*�u�T<uzxNN�����,� r؃1�R ���p����������>Y���f1#,��n�s�9�>;�:����whU�T\� ���Ug�4I�w�
ێ�Tr��h�v��$�#�ϴ�}��������UQ(t��M��vX����Q�ܧj�`[u�WS�|=��k����p�[��|K+��/��ߵ~�:��S�dY	V��tx8l�!~��F�h�h�X�$b�(C���0.������Dg7O����v�-���!�����~�+�%����YG��xt����^0ޡӓ�)����u9�#s hpn�
j2����Dq��<3,>G�`ֈV�C�D�/{�{��.=2C��mX��:��=�^+�u�
���rb�9'f�����*������w����a����!�Gd]5�Ѷ�����#��௮�{���N�=�鞭,eKnP��t�Ϸ�c��uďJW��k��y�2�^��Hx_��b�.j�o�y�
�w{+1x4ꖕ�C4�h*��nho;ˡ~�@�W��|l��
�)����Ft��{93��<�p�g��^��K��G*cY�}T�o�����>Ο�눙Xo��ahf���"�3��q��N+*�do�|\�ꇿI�d��M��~��Ϲ߸�����q_��!o�.<�S,��ʁ3�o�t|.���~(��p+y�3!S��y�\n��/�$l�:mgwE^/q��{�r��C(҅���t�#��!��<� ��A��k���bo�R��v�����-�:�p]����.^�g>�Ğ3ԅ�S=�ꥎX�� �b̏!�3V�6���&��eX�#�΀{p���⬮>ӔQ�x���l	���H)���G��'�1�m���#}!��"0�ը�X�K��3��SR�7%f���x�ٱ}zD��e��v��ι���ʱWȠ��9�]�C�;�]lO�e �q�C�_h)K�,QҜf��3uw�s�+�tk��^t<����p���t'�u򠸫ܨ�
���!��9������uL?����j$�Iז_e�2W��QK���p�h�<V����R���)�3�}�7'ǭ�܏_��ћ��e���͇�e��O�G��<�@�U�槅`+MG{kB�T�#��mO��m�N�cqER��.���+��=2Q�$v��˦��)�}����R��[g�_YfqZ�<�'���W��ѷ�o�Jh�z%��%M972B�;f*VӣtWzj�(>ޢ�^[\b�lZ�����P�
=��YnCm�%`r��B��N.�>�rtV��=��."�g�f̹��*�]�X����^���W&�� �۶���^����u�g�������`Q}v#��[�ޗ���1��ˊ8�����7꺇��W�] ����LV�R=�FLל�t���ǊL��N���:<Ⲑ��T��x�5����g��O�3�N+Y�{T�n~�{�3����}C}c�=?�oj��u�^-)���g�P��;����q],�\zPX�!��Y~������+�?���yW�z�!�1�1_ǯjD�xu��̖�U썅��R�>��L��X�ҡd�L����H��z���ى9��P�RW/�=��R�t>��m�&�=��9]n����܏VY�鼅�Nm^�����ۺMG�T:���ų2d/^θn����<�*��#�}�3*>��qY5�R�_ޤ���"�����=�i{�ƒ�y�pΩs��l{�a�Wz��Y�{��,4gj�:�7�)v�8{��P��f�mt.��#G0��^R��Q)���cre�mz�u$�ߤ�4g�����L=ؿqY<����ȸ[T�����!���9l�����^��IH�$���H�b��v�+��� �_�6�e��=<ʳ(��V�u���Od����\-�5�]W��O�y��Q��=Ѿ~�@���`��."�y9�X���c��\|�OI��~uc��(��Tћ�2�.���<���2J;�*� l�)*�>�ρCj;��0�@�(�=D��F�p�d��Wz�W�8n�I��q>7��Uĩ��v��4I�[F�/�at�y���������1�������^86ۯn��UĪ�3|d��� ��G'�B����j�|�n(�Rn�mF�Q�¡�ܺܔ��.�'�I�o�U�f.:d��r&N�>�7�(���p���V|�
�[����ӏ������\ύ��Ц/|^cn� ���?V����
yLTt�w�s���Ǚi��J�W'�}Λ�c�ѧR���y��h�Y����Pi�xMsK^ξ�*�x��.�^wPuۺ�35w�He��O�V��Չo�Mn~��<ğ���J�J�L�<۠5�5C�����Gj͔9U�;���yʇW���l?T����?S~��Q��7�ޘ��qNM�K�;b}��c�ё5tϹ��|�k��T3��	��^�CF�a��p����u�gu=�w%x�6��j�k�l�N���,fKni�+��i箰� ��a��	Ee=7J|�=H���KLu�D�y��DINg�~w�����*�rM�>�{^��z�{��z��,4_T+����d>��*�q�ϻ@݅�(�������d\�db�c˧�߫�ds��~j��d\�<=s+	��u�i�E��g��ѷ�5�YT�����K��<��<˥.)�T{��^����D�gO�K����i��Tf2N���·q3�1,�S��i��]@^u,�)�GeuB�n>XR���ꝏNs�p��|[s�2�E��z��
���p����qd�Uk^1�>��B�5/{�sj�`ު�,����{�X�<��(�#Ĕ��H�.R7T�j����`]/ح~�ܬ}M�4�����!�,��ɗ;�	�)��� ���owǫº�)���Ԟv=��E[T�'��Wx�I95���EX���&�����j݆�{9���2�gI�u��u���e���@�d�Xm�W��Z�����ٟN�6���u;�W3��a�?W	�N��ȍ>��-3 % \�g�s��Ff���3�gv�L�5��io\U¥��>S�|wНp�m�ԏK�B[�.WȀ��F�7S�;V�뻉9���\q�(�;O�0��i�I:�.�il��x���3l׾�UD�QO��+NR�^�.Y�K�@�jP��z|=�
f��*����r��C6�}�5�t��a��uq'��u��OȐ����7�̑�p6�u�����x�>�tB���rb�'f����9OWo��{��}���	��� W�e9=��_�wެ��]�C��xb�V�,�@�ldoE���95A��М�'n9�W��Ɂ��\��0���W�:���^/W`� g
.��<3o�]c�xhp���dwU-+\�i��U�p������A9��|G�0��l�d<��j�k�:7�إE2|o�q�����K��*cY�}T�o���'��Wc�Ý)k��^mߢ8��я�:�YU�!q<v<T	�>�y���@�R��O����ƾ�]�L�cח���Ջ#���G2�-��U��G�[��ܩ��FuF^�]�^�,,鼦n»����v3K�P�kIn�5�3��)���=Ej�!N0�D��]CB���u��w1+�[�[mY0#yC��]mDq�t��il�A�Ã����q��;�r���I��(\��J��t�>�h����g��B�w�*%
���s�����m߸���]q����pe���(I/���!�����p���N���|F����n��1�����s=.x=FsL(Mz霳�uA�|A�C>���qU,ro�QO�=�s��;�E�a�^Z%���΀{p������4�P�J=Kꅱ�M#�=�쫦F�_O1��E�΄�D,^���JߎG9N�y�M�>�=p��4ωW
@����I��(Y{��΀a�@��ٿ���Zs�yP�R��g���7'ǭ�܏K�FN�)���%U%���� î&@��0,NxV��{kB�T�#�m�}��=���ū�Ӿ�n��k�o�d�X����G� w�A��3��q��]�<<�H�Έ���}�o��QE��2{!�@N�EzTӓt���ȕ���Q]������~�O��y�w}�3h�>��q�2\2���#q�Rq���rn8�/���������Ou�
��kZ�m~f�~՗�F����ynjcC=�@s� յ�������`�mfT�ɔ��4[$��ʕ��nq��_[����&J��:��赳wVZꂙ�Ib�U���g�a�����B���u{�F�m���bP�5&���Ev!��\�� :�n�^B3C��*������{c�%��E��36�N�m��o0ty��}�ߋ(חw�`^������t�n}��t=3}>U7�����֫Q�`,����O���C�R�O���7�ڄx��
98�g!�S���ա7�D�q�==���Ń�~�?�_��� ��IcJj����v|��W��>Y�V0���:1����a�g��b��L���١�巟�z�ڳX;���H	��pS����e9W��>��+/ρwm�j��+���o'�=[sƅ�ݰf���)s<Y�����|~G�l�������2<5��P�T���<�u\�B������<I�W��<��W������������##�r;j�Yt�����u�\E5Ln*��X6rJ;�xj�e��nvj�����N`1��]L�1u.�fQ�J��2��%s�\-��I�4������p;��K��*3�G�iL\T�'9xU�)_X�i5�$�`�"��}��j"@l�����W'Y�o:�:�T&<-Vk��|j;���Y��j+��:�R=uoE�r""�
��+����$N��Bv���l<Ɏ��n

�u����t^\0Y;ެL#s��y�UY����as��+�l����}+�FC>�ͨ r�� i�JC{δ1�e�=%�Vxm�����Ri�i6��'��:������W�@�'�mK����1�J��d���J�q�q�!����2uļp2[s�k�yr����W����*{k)OU�q{j����>��CF���P��[���������`�D��3B{s^bY~�9��7�K8k��ȺN�/�s�8:_M��`zy�mzS&��n�ב���>dTL�Nn�>�|C���g ܱѦ��Ox�]/SzW�Gm��Ϸ�ޘ�'��K:X260��J�8��s������t=iP¡�V�@�t-W��`��M~Â?,'%<������">��loJkm����J� ��ʵ��r��5��'�By�9���42�u�y������4��K�!��g�v&�������F}=N�%O\�>�zu�pw�瞺G	��Xh��Q���Q�!鎪�v1G(�r���d�����r�"�s#>ULyt���{���5[G��	�ꏡpne໎ʱ�QA������\s+���A�cMܡ�kW|d2��vY���%宁���<��+t�|�<;E${*�&t���
�n[��#�r5����r9u/� ��K\[g�p�__��˰��29s_)�6�wi�vVm#��R�Ʈ��HR�7V���w'&n�{��h����1r�M#i#�	W��
qyj�d��d��u���^��/�Z�ZJ��.�^f�}�� A�ǎ�x��m�Ge�o
v�>r	������^l�.#G��ŷիfշZJ�5y����A��L(,�7�b��3���&#���3��^0�*}���Vv�<2�i\j%Ђu�Nu
KfA�%6����mb��J����#c�+�>�a�w�I����m� �^��F�w6���wزWu�~���[�op�s!%.e����{H�ԏv����m� �
�4��å�%
��{e����݃�ʆuk��P(zWK��;p�s������w�+�׶mlf����b*:��ɡ���B�к�;��GmN�)�U�Pɚ;1M��Q���%E�oet��FqSE�pnZ�P��E�D��Q��\���ͺ-T��;�V�`�W2�D�ʦ�]�#X��}X 9]"�W�Ɨ��O-HPj{�W�G}sM+�M��Q�}��T6�ݗAC��G������D�e׫��]�Q�:X����8	��^\[x�c�T�j������a����E��+�_7(�픯.�72�zc���)��vԘt$R�l�����d���9��9�0%��hk,O���(=K����Iu�'os ���Ld]doS��aw^ք ��S�:q]�P��Wc��u4���[�ek�l�x��_*�Q쏥���>oc����;�7ݎu�B_t�k��[�{U�<��+}j��|l�LL��,!�2���N���ʝ4X%�$�++�=Τ�pM�W�ٌ�A�Ab�1��3���S���v�	!wb+�u�Q�{T�Ckj���n��+9+s6QU�q[�\=�j\���u�d��e�R��+�p�{]:Ѳw>�31��Ԭ,�b�V���w�f�4[n���9X1`�t.��Ґ��X�g=�]g5�ֶ�|L���ߘ�����d#GLYm�.�J]���]�>�(`�([e�Ў���g]ަ��yt_J �Dr<��:��F���%VՋu)���a�}��t�]�v]�L��M7m���͹{	�8�%l�����Ԁ��˱�.	Y�Z��u#�]��VkoR5Զ�{p��ș���+��`u����+���2�"Xք�ulyV]�wLhn�J�|�O��2��հ.�Ì��|6�N�u��n�Ac,�Q���󾤅R�Z��ܤ2�����M��0屏��D����g�b��5�p#37Hyγ <i�V��G�qO���" l{l,��S�}�[QB������ܶ'w,F��Ė��ػ�sr�5ʍs8��w�vZ����-t�s�wX�]��w#\ֺV��K��u�Q;��+��\�s�.��sr�Ӻ���n%˜�+����������M�.K���Z9r9cwth�%���H��wVwE�9�ܴ��"��\
��CFܭ�+��nI�ME'(�*4�僻�\�S��˛��ns]�64\��.Wwd�r�Q�swt���U�I�wk��5ʊ�;��t�������
��n`r�87�Q]Gsq�]Q1φ��认©M�I��\��R�]|���]�����Y�so.rY���{���yW���o�}G�>6}.\*�O2�C˄��}q��-Zms0扨�������:��$�L��&t+��_LJ#��B٦Vu�^w,�)������5&���
�Y�����g4��t�����A�3�L��T�p����qd�Uk^1ᑡ�/o5�*�xu�c���gn!5p�>*��y��QF��J�3�H=Ċ��#$��N=�2ՙ�^�^Ⱥ^ҷ-�A����h��5��ۇ��>)Ө~%��1��@Ua8�5I��!&���Tu?Q�8�0ѥ�p�vpG%��s�ķ�R=t�Л�ꋛD ���~�r��vlh����wF!D*�zy�0��v��������[>��^�w�-�c5�6��\����y�s�|z�����6��R��{ �w�T+��ܔ��YE�2\ꮶ�1Q8��Tc����z��X�n\�t���b�N�BY�5�+Ʒ]�uT���Bp�y�͋*��˖h�*��Q��"��S��.a���1_J�_�����P�u�{a����׽Xw����q��*-[�Yb��Gm�<5m�	��l������,gQ���#��S=\rgx�w�٘�Y�jM�����{���X�٩,c�	��ֱ�?�ۑD�qU��z.�@:{��Du�wKu�Zh�"ә���y�f�+��:7�gg�ه��M]ȸ^tM���������~B8��T�r�EwHWN����u�V\I��{;ӛ\���>��C��KND-t����:����<�P��@�@����N�L��`����%���+)�=�|n<S5~��2'����TƳ�>�b�<�<-<�Q�e�dD�s+���]�4S�g��AS��YU���QT	�5p�T�2*t�~��w���^�A/~��>}ׅy2��P�'ze�3�����!�� ;`y\
���35�T�̒κ..�}�YO��w��V#kn�в{����BI|}�)����}�8��R�9�w�W�^poí��n�=�E:��!M{�\&�t�Y�O�|g�	'����~�#�f
����!��k��?F��c��l�<������ʲ�,ӔQ�x����Fb���ǏH~>� �v{x8���(�fI����늿�+~<�j|�΀Zn1��N퇟i��>Cد�ѳ�x�圡s {��' �ځ_�����c��Z�}�>S>g���>=p��G�������ow�VםQ�[�&{��uc�V��4HJ](Q퓯�;D��9��^��i���L0�OY>���
l��`F��Z{���d���L���!���x����z;�]��y�t�^��T���0qW��
^_a:�	�ٜ3w!�`�]'P���*�Y���8��f %P js´���Z*v��s��m��RU=s΋>����k���_.���wlйUE�Ar��B�N���:�;nB��_zI��f��G^F8K2��AÖ���g̕��z'��Tӓt��혯�Vӣ!vM^hTL����M׸?"5���Z]w#��KA��>F� ��.CYnM�_;u�on;re�y��5G�n��>G�采ݫ��G%W&�^t����21F�����Xfz򱹋^Nmގ��~�U�懴��N��^񸢼^�Ҽj/ח#���Ů�to��+r���Z���[ ߺ7��c�>iP���\O����=u+��ߏ3W�ۅ��O�98�3޼��@��u}+iMd���{�N2�߿�8�R_ØŃ��8�o���ǹg �
W(�ő�^ul_�Y�f��SՈ����[�;�=u��>�0��ٜ=��劢{X�S����f���y����{��2�O*��K'Cz��'�Vz�Bc���\�����Bҳ��Y�w�^��oek�J�S4w�.ӎ�d��h��r�d��tܛajw����:����):��F=��k���]�΄�,B�Y�m�|k]�/1t ��6pA�n�N�d��oXҥ���1��)F��~�f&%X����������ѱ� ~���ע� �;�r��������<_�����׵9X<+홋��w)���B�2���z#qj�X5�ßy�e�#��>����S��L�%���?fz=��h�|���v�g@��"�R���\��(��+~9�C+NC�(����'ٟ^dٶj=H��(��5�{>�3����t�1q3��}xU�)_Y�߹���W��f�fK������q>�wh��g�Y��9Td�g�Md���z�Pf���Ӟ�������.�1϶��']�����|n۸��4Q� .؁ h��:�#F�1ѱ�;#�5�Nc�L7Q��!�I�C>-�����x�X�*��UNf��$�6y��+��3��gJQLY������_�5�¡\G.�&�u����<ЛО[�ٞ��7Lxϵ{]�k�3R;�ib�k��^�q���w[�mw�"+�2h�n�׎;w���N��U��f!Y��S6�y�%G�Tj���c�l�w=��t�LW��ޫ�]��������qc{0�M�#ܲ�a7CxM-���L�i�{]L�"��!}ܴ Y=�QDC��c)�kӭ>
���\8��E�>��&��i��7��K7�;��H>[Q���6�YZ�Sk1�\+������gwf���,h���)sT�i��|gY@-���E~X?W�.�U#5��4z5�'���z��O�8#��rb��� �z�t����YY��{���:]���y�{4�vG��i���]a�r	���>��W�������K�����3�� ����n�ԯ��/�S���ѯk����]b��\��}�=�aA�׏���Ks��s�ʯ��O_� &3�Y��dd|�����7����=�j}G�%�O�6�=ٳ���ŲMs/|gj6��q�����p;`yPʹ�^�yp�X�7j=>��"&t�Ĕ]�>	zrO�I�C��*e��ґ�n!l�*5����D�	��'�-�3�4ͮ��V>î);��
k�n<��e�A�:����p����qd�U5>΋�3Fd;�����BÄ¦=�t�M\=Ȃ���}E8��� �(�H�x��H�p,�B/�vx�s����¤��9�4{\�>�:t���,�" r�3/���l��̥H*�𜯜������K��)�>;�놓?:�����p�Qk1��?��U�bϵ�A�$٤Fyc��>y�䗼���B�\��ǹ�n�K�}��k�����M4:I���mC'g�NE���כP���F�{;Si���=H�6�ke�g(�J��u�L���M��w).Ч%���Ш��i�=� ��3�ӝ�>Z&�ͻ�j�]���O�b�H��A�_��x&���P�t�P\�Kg������K�[q�6m8N;�=��GK��r��b���+��g��p�+N������%���'/�g�;+۾wG�^��Y��^�+��*�H�YNOB���߾�:��s�5~���^t=κ�f\�*=��X�L$��ܸИ����a��'��0����]���R�k�s�Ŗ�O�v]��W&��C\'w����܋�y�u7	�v��W���=P+��s'��-�����إ&9p�]�۸���	G�͙Ǽ�i
�^Z�ONB�A����g!����=�3>�@�-�t�q&	�'���wXԂ�/f<�)q�/����)���{hd�R�9ʘ�s��LV���Sv3:	
iw�?*��X��п{��Ȇ�crg��d�*���y*k�!S�3�{���r����r���![���3�o*tj��\���t|%�p 7����
��WvBh}�^���;ԣs��+�W�w���#��ۮ4,��2�P3���|n)HG�t���#)s����1�s<����G�V�ұ�p�Ջ|L� �6���Њ�.����jU��J��=�j�e�X݊�W	z�[jv�ۥq�M�*��6�{��s[X!�ǇWr�y�Q�����)�uos�pn��b*�w�I�5ڵ�gl.��#�Z����|��[��;����������v�ct����p|���׮��<I�a��	U����m�IQ}��u�Ӟ3'Ó��A�n�=��΀{p����*��\�v�J��Ɖ���2�/���(\�?������n�xs*�TQJ��9N� ��>�=mݰ�a�t�3�E�r*��7�ħ� ��$��`Xr���<V��~��*��|�|�il�;�G�V�}H��ޟN����f��P(ڂ8�@��%P+�u9�P��mhY�*v��Q<��4*�G7���K�.������몦hzUQF���!u�$����B��>ρc���O���97����{�F�MZd9}e�s>d�&2��<wQ�'��$.�rE�L��:�,�N�E�}��1vP�3�OgC���!���r/��K���E��]@�k-ɸ�$�#��X�F��x�/ٸ�US�w;��Z>�L<>���c#���k΀upݰ4��������]���f=+���tfq�c�7T+�w���?1����5�]߉�|����K軛�a���S���\w�,y�;4����ѩ��M����q�%s}b�	ڹ\V����&�<6��d���{N��-�EQs;5�{k���n��[`i5}��Bgi���(�jվ�R�%!��r�u�TV-��p��f�6ˢ�N���7��Y?b�]g6��$5ћF���]{>K����}ʇ�o�@<t�������|o�f�׷'���.���Fp�>����X>��^0�n�
܏������k�����g����W�V�	O��9+�;x<�!��?<�op9��%�쀥�3���=��}�w�Zu�Y�YP%�B�+&�W	l�X��I+�w�3k�~�~���$��1U4�z�Ӑ߫��շ<hY=�aa��Z��W9��	�[{�J:�ƿ�*����uǍPc���@Tw�&�����c�V_�׮Gzpf�V�C0�«uf���N%ᨃ=P����.#-�Adt�眆_��'�-K�t�2��k�r�=��=ٜ%ڞ���L,���/�\�,�F�#�[��C+���+:���V�3�o3c�zٳ���{�)�2�4���-3�L��iL]L�s�xU7��.�����9�g;~�|}�����:�F�3�,���� l� �@�;<�j�.�@zr⵫9>��^im�c!�V�9���봛~w�p���d��@[�$Q��j/�[��.P4)7�|�����kz�Dq�m4J�Y����]��j0,A�޺�҅�(��#������B��L�����Wǝ:ة��8w���Q�(��-�FuNԕh���;K�X�w�W��vab�~�Ga��(<�������E���/���:������0��ۄ!i5hd�y�3��۟ ����s=�ׂ_Vf�[{�ۢk��#jU\��L��0�9u�7�n��� y�5�U�����a�Vށ�o�q�=3�%��ٱQ/k®�3�7�ku��g��T��Jd��&�W�I+���X{4�e�ڡ������l:R(���a��8'�X�=���\-�z&4�5�Qo�FG+�^w�ͨ�&ߥ��n�f�f�k�OT�]c�஥��])�>>��c�:2N{��6�;x5*�wR��t5�C٦k��'�b�[�o�d�����x�V���@�Z��;��P�=nQ�(���b�`���R��+L����/�=t=�)�>���-������;=�u����ۨw�eW��_ޔ ��ˬ��y��X��K'F��a�CQ��̡�����~ڞy@X��\U��iC�xo�}C]��ޮFr�r=uR����
9S*�l��_r��߳��9'�E��z�P��L�WS/�.��k���=�*�z�{�?M]��>��k���R=Y)%�w�l�r���t�e����Q�n�\}1�ɔ�!M�C����V��í�=0ংt��i�aw(;t�GΘ���`wy�P�-�ҡ�QR[ #:r�t8wn�W����~L\V}NQ��nY�9]����g��m��G�7<�e:��3zZ;�Q�$Fcf|P���R�K��)��+��u�����qȷ	����=��}�A�MT?6#��Q�q�I=_�$�9��p�
dʲob�_��.�t&�^
�;���-ǴYیu���v�F�QD�oz��ӣ^^���1�vWl.qP���Q��~�=��T�8a^��}	�{M����ݡ3�o�|{�o��������q` Y�D�#|�J��X&���V���>ґ�|_��ū��ڡ��OW٧v5g�>��������xNh�r������'�]���ߋ����iu�jc�U7���N���3����k�%�s��ϑ�9�`+�'I!j��`�����5<�(D6��r}C'�{&q��1�:#���!�EBt0�Me9<!�Q����)�z�'&��TX�Mnu��t�Ά�<saF��*1y�u)��>�qXu�L5�2z��-n���T=�feft��#M�a��w�HxT_�.7\�Z�3W�?U�[-��ߖ���薩:Llͼ�l�NQ�(t�Ùk���⍽�;�(4ͩ�n�]Jm[ɫ�=|��;�w���r�2���w��X���jm�\���%�`�y��v�^ uZ�i,���Fںrs�I(��	�>c�g.Z��Z��X��=+������ͣV��]8v��-B�g[:��ӣP�ޛMַͣ��5+n�M93�k��~���5ݍ���kj�JWð�!�|���d']XI��X��C+z�}:�F���ţ
I�g���W]�C��9xڇ( ��������u;Je0�)#`�ˏiT˼�#n�{l+�T���y�[����
.�k�>qU���
E�Lʲ�
�����V�Hu��\VwU��7���OCs;2Q�f�l��v��tÒ�]Ƃ��k�	�{f�me�ס֭��t�j�p\|P�)Y`,���yb���Vⱹ���4>ħ\�K�� �]&c,�,��N$n�o��*�]�n�H�^l��凶�!����0/hR��1�m��6je��;����C ��5�Y�<�W��И�[ʡ�z���'��u�B�b��ۢ�T���\���Ɏ�`�6nQ��󻻘�}Y��v�gZ�X)��7�rS<��4��f,�&[7�FE��*.��f��h�߄���b�Q8��ROd;���e�N�k<A���u�u�*����g1�VDWlZٽ'�p��a�k�ܫAF�H=�wO��r��zp����l�)��d����OU�r�g#���DF��)���-��6S[i����f�A/��.�����V45:����hs�``b��gfQ�٨6lt��<m�N@dׅ�V{��]�� �p����S��v��˘���[]�6�>��P��+xM���hΙ��f�����Z/���ݝu�k$���ḷ���-�f��Q�h��*٦��g6�56a7����J�-:��=��'�z�� ��U3�[��:�5����e=�p[i)�yZ��,p�v\�}i�@������Z���#�j�3k�C�,1�wD�/v������S���&}���U3bks�W3
 땮?�(��k�:���hP�؏^`���ۗR#X�I`Rz�n�\�ʚ۶e���kǴ�qsHd
�4t_[�g
Yc9ԛ}Q���/��ͻ����(i蠟�t�Z�<:��6�f�����@���r���tD��ʓ��s6oMom]Epn�|m΢ ��E�`�1C`��#0��7���um8y���:��kck+VG��ҫ�V��]벴���a;���㹪�'~�V-�ݕ�j�<�� ��1��.��^��IY2D:�W�C�vi�L��+3��Oy���k)b��:\0p+h��e\�͸��͛�h�� W��˧c�+{���ٌTM�1�k��Zn�[���m�M�Vsb�1\���F�J�L �/K�
6���8>����u
�>��(
�� ��\�6ws�h��wj7.�ە�ݤ���IwuGM�h�F��wmr.[�wm��s��b��5�wQ8j�밍shL����nr*�\��F1�%n]�]�9�wU�d�+��T��N��\ܹ�9�s�\�w:��u�,\�nnh�˗s��r�\��M����]���ܷ-�\�(���6��]�I¹m��(�.1b���r;���W,;�N�+�rܴ�Gut�nnrt�4��Pwv�b���Ɋɫ��!1%�lPk�Js�����.�P�W���0QǷal�����0ڭ|r��z�V�;��Mu8Qz�J��@��Wk�0�se�XJU���:��9�4��\Rt��]&�N�X�a_0j�{_�ڷ׸<�A_~�0����r�5��{T�j�2��F��G
��:�,�1�>y^��ف�*��Y�Zds$z0��j�Mr 3Cъ so��`eê��a71�{��9�T��'�tuԺ>�}8y���0ۏlO�q���˫���U��w�R/ߋ��_������εV ��~���hlJ�nǜ�k?p��U~)��� Tg'hN|�&z\�z��I�]	I�����j�����d˗����tL�7xr�[tQ�Շ�Z9�ay�'h=9
��,ӔQ��s�﯀�Tq�uS��Q����.�:� �>��X�qd�����9�9N��Ǿ�}Q�?��d��\�S}~��[��!��{����6L	{����ߣ���R�����Y����<�ѺF��Ю���\r����Z-���qU2�S�gD�@=�s�z��wV�޹	<�����e��0��m��9�ۨ��wlйUE���H �١t�Y�Cs�ylC�"�kL�A�Ӷ/sz��@��������B�	�&^�����k7�:��Ir(ͦ��e�<���s$~4&.��ur��{I�sD�J��(��|D�/:��i��7�m�y�N��U�},�+���[�z.K5Ҹ<�ؓ�<3��-�W�ƴ��;I[d9}e�s>d�7Q�	ۨ�D��'�!v��Z�Q��c]{&��7�E��Q��ɬ(s��"+{]ȸ䩒�9`y�B7Byp)��'&2��S�ϝ���P�9[��(?|�߳����Zc*�n�Z�Uɵ�a��7l/���j6��{ʢ����@����nO�H^,�puүx���Ǌ�]�˅���NB�@:>ǎaP2.��ǝT����t=p�L޹ �ӓP2puӦ=T��~<�D_��T�X�9t��z&^�μw��"��S��Tk�4�3��A���ã+���]?�����(������p*߀�q���N�����u?b�S���5��H������w%�<A��pzT9���hq��G���p�\��Ϟ@�T������[���{�s��!ǜ�w���~���+�̌��/�2��:�g����:�yPʹ��}n�k����_��l@[�
���U�m��xkَF��O���љ�Azdt�ݵL,�����S���\�)0=?j��@�N
��(j=×2�eb�Fѱ���pѽ![8&pʟ��߹��91�U�qY���|*��rruie�.e7����]r�{؆^q��`�*뫧�m�U�w�ګ����|�u7�����p� =�Svwk��bΊ��,9�cÑ��y+^�R󺓿�7��N��.�t���~�^�.4�/�x�u��ϳ�G�m�<�����q���;cl>rQ���q�y���pm9Q�`t�5�-)���y��o��{Sq����Z�oE�s���������>��|v����'v�,��Qf�9Q��	-ueonT�
�`_��+o�u?W��,*�y^�Eup�>v��:�&�~w�;�����(�v7�����}���.��1�@*�pN���{p�j�Eβ�!��ɶ�h�EL��sWE� �{=�j7����/��3:td-9�L&{�&����n���1�n�g�^�.�y���������?Uw�R���\���&�~SI�Q�Xw�aomT�o_S����=��F)=�#=Z��H��z��#��uӦ厱����c+�1W��/XS�n��U��j=��0�8��،N%������n�z����\�z<ao�z��¿ƭ����m�ՙ��L�]��_��pwR����f��i��nⴧyN����k�����p�H�,z��P��?({;hf@�2���h`xz�pR}Po�m�t�^��IY}��'J?s삺��h�7Wg�e8�c�
7Z���S����Ɔc� ����J���x�Wj��x;&
�o(0`�
]�yw�w(�d�M��T7)�4�޾�~F<�����|��V=�J�BT���!���X/���C�9�}Nz�&���ק�̓H�!�S6]��O =Ϯ/�ι��*�<�}��sL��W���hZ���Q7�����U�ӄ��*�;1��
�ﰨ��β�7#K�Cb��UnE�p.�XY'�`'S�bު��ߦP�'Bȩ���)�w���2T`г.&sy������u�o�x�)��˘X���mOx�9}$�1���OW�iV���>aW�(n��)].M���c=��y�gSU�U`��rx���xw�v6w��g�Y��|a�ܶn*g�,��<(\*N�3��w�gn1��i۸y��C�>��S��,w�#��G1y����@Wǥ#tax�n7qW
�gS�|w�'Q�6��G�ww-�j0Т�}�$�+�2T�� �$��=����u��L%	;H�>ґ��xf��ut��\�:��<V�cUX�\J�%꒺n	a�qS�,zgc����XW���E�
.@'�OiǘN��W�����8����u��"�s;>�#G�Ut���)�t��WZ�Sk���]��́Y6nڢ�R���|����F�nMx\�vx��vyu�����z��	]]'�n�$=4�v|�_X���LwP^��q�t��U������o�����s��+"�9�c�e97�L����k�%3�S��ǽ�#��̗eG�����!��Rc�:!�r�y�5�N�*�rxC�>��e$z�Fv:p��G8̹xzW�_�2w�xϷ�܋��A��r�ێw�\d���e̞�ŝ��ݹ"MULԬ�j=�=�N�D��7Ex�ͮ~����ON-t����ّ���TOD�{�j`�[���{�A=�i�7(8���7����^���~9�X�}�p���111�U�N���wk��+s�����+�}����V�.|�Ui���$W�T	�q����rT�y۷g��z���:U�[1�o��7�9�ޓ��b��qR��_Ԥ>�c���F�CDQ���x��ӯ@q	�����`r�i�����7z"���:r��fxe} Θ]+���b��
�ǇTu��>!~3C����rv��t����p}�k�a5�Cb��u I�na��K�c��v,��Gr���	%iqG�+��@��=��}�P�Ӵ�7<��z/Sj��7H;Z�w)PV�Q�6G|�F��(�����Od���q�٪�MD�K[�NF�m�ܮ�A-W�+��,q�յ��x6�#4w�U��R���m'��eoWWn��,����U�!�hgC�=s6�^f�BY�T�S���Gn���v�_W��q��Q||I���@�/j��2Kʳ���<�j|��N�@;Ӿ�S�C�s��Ec�ie�����]�) r�4��C��tgO3���p�_�}�\V:�ٯV�Mv[�ai���^w#����8��d���������bǇTv>��Ëkҷ�����1�9��	���m�O�ݳB�UQG�����{4<}�rp}���GJ�8��1{됮;���9}e��3�M��G�T'��Tӓt��P�sWa�m����b���s/�jھ���z��F���q�S%�|�<��;�:�D�UD������]����%��I�6v�+�����ʼ�^5��hrSR{��aշl/���i��L5�Y��Rm`����Y'�HZ|}8�N��qEx�q��z��gs�Ҷ��O���y�{�eV�Q7(N�%t=z�zf�] x��&6�N�,g��^'��ǙE]�wl���;����w_1� ��]#S�Y�w�����J_���_�}��ő/�Ψb���pl֌��9v�����=}�Zi��)D��ԂgM�i�N���hͮT�ֵ��t��.aѦ�Q;κN�����Դ��ܵY� ���CxRfU��S�1�݃���9t���|��V:�_)]�1�/$b�<r-�:�dWq�}Xr���I��	�#�ݩ׎j�;��8���+7nߧ�\N�����s��(��&vς#C+ȧٵ�HW^u6K�أ��xM�����R{��D��2Sg����q��W�x�L<lf��d����ɜ��ь��;5�ڏK��,���z���Tw*����W��5~����|�n���Cȹ�O�J�PfaTI��G@�=�9}]Q�B)��>�w�U�\�V��e���t�1�r�o�]^��.xz�t	���\T�t��:�U�F�:[��'�O�Ǹ�z����V\7!�d���j��B��/#L�(�� �3�Oç��ҘE4ci7�[C+�{<�'��dwg;]-�W�\�lxg���q���O��?u���;�a�Qf�A�A��FW���18Ɩ��G:�7/�j��z(\*]|3�>w�S��<��'��ڸ�nh�T�O;�)�Y����K'��b~9��[�j;ۄ!q�MZ���������,j��D���8���9��UQsq�W�-�Q�+O��a3Q��P�.�&�{�?A?~&�۠���LAXJ�XU��F�%G#v�F����Il:s��l�J�ѵ����ܠ�s[���k��)}n!�.�('0fr�v�yN�^۾�gK�Bم�����N����/n�ޭ��:�p��$��k�Y�CoL�@��q�҉ͨ
a��;u�R���M�),�Ī�3�%t�Aٰ�^��9M~��>����x�=�Lzغ�*f�����yܖܴM���"���#��u���c�l�(��}Iׅ{�,�T���Mkii�\<��ܘ��\�������9�k���Dʸ����>ܩ��1��'����w&ì���l��e�;���}��9��L׶!���|��Xs\�}]�+)	j{�~�'�7'_�_�s�m�e.7N|�ԃ��@���u*z���g��u,��"�߄�҆�A�t1�)�9������~���>g�ұ� ���[*��
e�[7��U�{���^{��~�C�|�m��s�u'�����uӪ񿨨����<�}���ъ��u~�s�31�!LǑ�
���'�B��I�^I��2�T@�Ф���!t����WW��(�]O��}η\���@Ĩ���r��}P�Ц���^2�E��z��� �/�/k�x�"���*~��2���S���A(�LX������&���Vq����Q�x��}"��gK�f�Y�w�F ���i��c���[z9j��sb�/��'qAq[G:�^�o�79�j]f�:�ȋ�F�U��]���2�� lg�����]�V�\�<��+v����c@�ܑ/�5�+�hsa�77J���G]��u����ٙ���9Zk+2gWw���D���S<9�,Y�B�'~�Z;���;x��N�á�3���u�rNn�����/�"�|f6�t e#詘^;M�V¥��>S�|u94���T*K���*��dk[���#�Eu�p���@�vH�%�pi�*Ćgu�ÿ��˩�x�WNW;�[sxR�~��\��6���wV�_Ҫ�C��Ӥ��9�
����`/�0ԗ�.S��c�-f^�V����,�8�Y� ��4=���$��顿J�f��<�۩�5o��2��8i�Σ]�D+��]ɋ䝖rˁ��G�b����FrU��36�G��
�)���o&u/Ċ��qv�g1���{]?�J�E�:��9`kB�l�5Ǫ�OL'~��� Ș4�[V{e̛p.cރ�0�N��!��n�~��;�׏-t������͢�1r��o�'<�xx<�G�E�oP'�������VS�+���x�5~��3���X��1�]\��~�6yH���3n�
܏-��O+�}Ń�7�����+���ty��q*�����^Ə�Y5�/�O�1��lx+.b+�V��ʝo@�}y���e���G&]*WVt���q���x�n�mNu�^�}R�����ީ3�K.��w��3�J���Lۺ��Ɍ*�\	����>�g*�X!���6z5Ʋ'�rV���]E�Z��T���4��N��'U�W�o�s�:3��>>%�x)9'æ;�"_:eg��v`;����-{���y_3%;L�DSˏn|��z�SǢ��
q�;�Q�߁r��S��+&�����\x���P����+�n�=.x=�5�1i�]q���qZ��m�o���N30�ў�.*g��S�9\-�(���C�-�g�t��wh=38=Rp�#Q2g)O�<���s�r�7�'������te
�,r*�bo��>D.�N���#^�G2+�toV["���1��-��g	H�9N��'��H���L�YQJ�G�*�f�NU�m]����N}���.���Τf��E0pv�T�	L�w��X������7�Ò��~�%���Ν�c>s���i/΢q�S4Ҫ�= �@�8�T�Ky}Zv��Qή���Oq�} ���N�A��Qng̖�G�l:�qW*i�������0��V���Sr�����[�^�L)�m���N�-7fe�:q��D~xxxx{����ֶ��궵���ڶ���U�m[�J��j�⭭km�][Z����[Z���*�ֶ��j�ֶ��j�ֶ����ֶ��յ�m���ֶ�Vֵ���mk[o�j�ֶ��kZ��Vֵ�����km��������ֶߵmk[o��PVI��}���sw��@���y�d���J��D�Q@	(
(
*��
 PR�PR�@  �EQ��BJ	BT()"Q**�B�R*� �����hP�!R����*$(
T��D$�J�n!J� �)ِ�ld���j�I�"��PZ�h�UfĊ�
��   ��9m�F����  �   N�  ��-GZ�Il�T�Y��X�R�  �At����E��35B�`��J�قSM@f6�I]h�"��"� j�'V�l�kCl���j��!��I�X2)kveR��TIb�%����"T�`w;5ֶC�N�ʹ�6u�5G��q�Mk �2�b�h���Mt㥳P�*�
Q��*�5��U�R�%S�4�*������3u�XlƵ@�`��H�*�B@���Bv���2��Sl����j6�QZ�J�QT�ш[�T\tсV�PQ
�ce���*%%[Qh�J�*�����"m�P�(V�сH����m`�h�i�%B@� �
�B��*�&��������I3jJ��     D�*R���M4�4ɠh "�)R*��� CM  ��"���d4dF@ 4 ��@�*SFL�&�	�M0#M�� T�4 &D�mFA�����I�2z�i(i$2*�       *�u[n2dۊB�&�M6Rs	�!T�@@Du���ŝ$DD����,�)H�BD��e���R�H�&+.X~ߥ?9_�����!�Ѹ�����FDI*,���� �$�Q��$�*�ʒ$D�:G?f|���o����k ��c�M�.Z_;ܿ��ZQ����y٥�9T����\�e����֏��S��K��X�W-?K�K�ij����WwtM\ǔ~'U���Qb*ZECX-���b����9�U��Lʈ��z7~����eϮF5[ScR�E%D��2�m�4k%\�ePK7 K=�h�&��t�6�:�t/�C6��R�0D�f�ږ���5V����Qv���]�klV�T�D�KXWz���Q1[T�k�I�{�"�W�2���h���!��;W^PZ��K��IVs9�u�| |����)�4�6��V���^M���8�o
s�%=Q���n͘3*��'_J�Tˣq�YHڬߪ��AV�.UE�l[����e��u����v�"�hD��u�D��ZC������?MW�(P��M5S2��-��Kt�UA��M�{yy,�o4<9��,�V�9��HX�DI�������Kt�+Ǻȸ���s[�M]�Qx%�ne_pyl#�hM��O5԰�7Q㔕��FZ�#�Bjf��u���(Y̫35CWv�K���x�9�Ы�nۦo]�ܳ�ҪX��M�t�jYt�I��Sr�r^`��"�f�h�It�t���32٣�M��$��Xn᢬�f�ݛ۵K&
�[w�"��ch�'�Zv�-*�̣z�31�o*l'6�V�ѽ�+U%���6�:,�db\�71�����*��	N�nnҩ�Q��l;5\Z�#k�a}hL�V���yX��v]Mv��0��e��9GK5[���Rf-�$�r�U�⧫i4�7Q�,�ذ�n躭aH��<i�yյ�͐Y�0�ދ�t��ww�]6[z��[�Յc�e%h�9����ڎ���նu}�����8q�6m��U�aS,����c�;�^�Z���q�k�"շ��m�f�9h�����2��$֬њ�mSd�&UV�8S/L�9�T�,�Nڣ��.@�t2^�,�/2���6m\Jk�5,9�"eVm�Q�Z�m�;*m�{
tj��x.ݺF��P�4I�'DŴ)�����Sόɹ��i�\�qf��n��E#�ˤ[�u�k
�)����V�j����*��nm�F��X2Ƽ̓.ͤ��B�m�&�%mлV�)ʫ�h��-̔DXP����cNÇ@��[f�;է�)���5��m��}Kc�V5�A'}[Wr�S����t�]n��ܻ�N,�IԂ�L�:2c�������
[S�v�N��g"Ǩ�б���{�z�I鬶��W�n�&����	�R.4d�o�q�q��70e�5Μ.��zp���*����^���O*�S/b��{u&O��_k=�ۧ[g�a�9W�Md�Vʰ�U�eٹo#�F�[ʭ�A����v�kX�����A�T��1Bqກ�j˦�!{���c�|Ao�� Պ�-\�hY�X�Z�;�
͔�"-�*cw-Yv�sFM��Zn����ޝ��+��:t����ʺT4��D)���{���ŉ�8VlA�ڻ�%0�\��I���;�R{)m��K!�U��1������2F���IgP�y :�>�R�7��D���h`�g#�!w
�ø(�5�fa�jՌ�ك)((ؠo)�8F�*�)P��!#�,X�4S�!�^^�����N����mEh[�iV0j���7�Gc%G�P��Z5��yZ�U�,*��U1/v��*�mS�Q��n˺[6�r��YU�pe�r�m�ʻ��uy�� �h0�Z��O���T���j�32�.�mJ1"ӏuU�\ �NsN�c�aH:t���{R���G������&-;{'vT0��kW{��I�ap��j_nU��!�[hTj�Zv��f��WW�#��Awv얅�5�0`��K�22vc��U��i���ZZ.,�H,�H�V�V�-�t#�����w\e3��2ݷ��{gs������	�A9v*Μ��]f�̫'p�/�{Mqx��W0�P�6M9W����3-��x������#�*��T��HAf�Y�V�J�u�e;�S1�6�]�cZ�^
�y�&���Bb7".�-�=��13��Q��0"��[�%��ʓvm��+h�9��E�ʔ��9wm�-T��+������^�Tf]��I;bl+CPa����ن\�j��Al[4iܣ��VV���ӧV7-6R��+��n����Z�Q�۩b��T5�H�w�I�xرM��ڰ[+wB��U���W������ʬ;Xu���b�˅��V��i�L�4-m]l�)�R�`3��z)7C�#
�B:���T��mŅ�Uc��]�D�B��jV���-�<�O%;��q�9z�}I�
�W��y�p@�gt�M���-��W�[��`��ԛ5ͫ�w]�S���ߩ�u=g��X��	%Z(����C��X�]1]��gtƄ����YV���Sxc��C2�F�ƌj1�ʩN��8*��,�8��z�'�j@�d5�Di�b[�yL�V�E	�2�F��CN�m,�ue����nG{+�3�9Y�����.�M��ܴq���	���ut��iP�u5�OrĮ�֚��C�uT�����j���5� XT��ͻU�Y�L0Ҡ��[Z��T7.�ݨ ��ٕx꤫-U/����������C��32�P�8^*�znc��]`�c(�����DZ�D�2Jk�7{���X��H������M��Vi�e��]+ks>�d��Uݗ6e�ԛ�k�)Zl�.�;um���%���ca����XS��2���3�1�ΪiVv��*ðXa8n镅�ƷF���Tv^�;6�{[���)e�g���k�MJ�N�`s!�+3%v�]j���������^�n���oM�F�������㙃ww�l�n2j���^��������_��w��"56KZ3.��DSj���0��Y+�1�;8
��NJ��d��E�ջsv�՝
����[Y���N��)�.ʳ(�K�^��lR�9jT����ĭJ��B�S-�F�ɽq��pdJ��ݛ�%��Иwy&ʋ)!^���P����wf���ZM�Ы�M������Q�{t�]��(EYq2����F<_n�E�"�d6&S
h���n��U�vL�n�T��8j�Lɠ�Ҷ[WJ^�N�l��If�r�naj��OP��&Fn����u�p�LUk�m��n�g^R�d�E{Y�1ѩ7V	�V�ɲ5��l5Q@�a�f��0���T�\������f�(�e�u�C#V�n� ��S!�엖3i�;�Ր�ĎU�tA�U�� �[%	Y1�Zf�no��q��*����.�)��Q�%[V̿�6P(��4�[�E"i}Uydj&�$z~�{Ze�7p\5�+�mGi2��퓪�C�5�kU��ZKt���oZ!�U��/wT�`��E5�P�f��Ci��YY"Z�醲��0ʙj������j�i�Pv��S�5�Zg�n܏��Z�]:k]����"���m�\�}�j�)��k+�N�u�6�Nul�����&b�6�P#a��W�GiP��gnܘ���*��yu�Qy�yݵ�2<�4~|�����Ķ�r��b(�J\K�j@��I�Z�A�ݽ�ܢwZV1�/(����m�3�i�����.��v�����lF��j�z�n���[��jȸ��K����%�&�q�bś2��j͛�s
�Ew��i��2��*��c��
�k�1���#�(�����/{:�׺X��^�
K�jtzҰ�ً�E0�x�I�NVj�wV\8��es��r�����{�qŭ��yA��D��`��ڝg:S��F��jN[�l���Sbr�/B|հyu�#�c`]ڲ����ҏ�n�vAs@ɑu*����z�\��+�Ȯ���²v��e�r�ݎ�d�����炙F;�*��B�:v>�Zd�u�9Ș�f��T����k|4*��A����n�d�&o��C(�L��ݼ��;o�ܫ��8ۙ|���Sȣ���֪_싻��<��(	��� ���-��z�����:���P��J�n��w\�,�NQnԽ��W�N���4������n�p��a���븷O"␅�G/P�R�3Ys��I��[���V���hv޳�LZ�P��G9�P��fe�����e�Pe��j�ˬ�j�����U�~�x_o����љ�Y	�p�q�b��
�
c���j��cg�\%��[K�܏J����R`\hPd]��h��B�w�ɷ���9���kF%��t��ƣP���یvNZ��޸γ��y��s�)�l����Zy�׼��RQ��(N��2�[�S�k|0����T�VM�CÈ{S�;��1�8�x����q�=N�˝`���Uz�H
���ǼjB4k*Ð(o4�vy�fta�1������!Ջ�J���˫�\���C���d�i�ʰs��>��[ev�*�:*��i�Z<I�9tv��b�̴5	��se�]�%��8#m���#����3A�݅�����ӹ�f�s�uJC�gRk���Xg�=s(S5�d޽/oUҺ�ّt3�����UR6("-R�}ٳK��ժ�P������-Z�U{�V�Z�x�Z��G��f哹)�V�6+4��z�����L��p�b�͛�ŧ0GVi)�m��=4�/���0i.I�^�Q�-T�!p�GZ��b�p�υِL���f�w5���p��Q���U�0�Ճ�m��]VE,�f][B,�.֔�٨4����&J3��N�������c�0kN��Z׷�!m��ޥk&�)ȼZ�#{�I�\6��KR}�4s����c�<�.*}��D��ë���맾26:eH���F���=�Ֆ����H�'k�w\�j�ڊ�b�zf��6>o*WX��X��r��{[��JKmRp�VTα���mNW�}�jǈWZ�2�v*��ɢ0�:�Jl]b�`Z����e�GK�r<�'J�*�E��:��u;%�*C��t�@�.tiVQDD�,4�٫���w��Q캍�:}x�b�b�y��3lu>em��3��징�f�{Ju�"c��8Y*���\��-m��f���:�_wȅ�Y�D�`��@�Z��2��Y[�{����ѭ�&au�B��,/J���4`�]��o�Ʌ�Y;�� �B3�D�Qcn�m�\Ψj��t�Mb:ُ����Q8��כʫ�N���[{��M�W�Q9w�U�X�aXM&�N<���(�M�镕|kZ��T��^+/��aI�mɑ�c=��:��h�yޫ"��sÕ�w�yt���^�û����ef�!���v!	,�B1Ļ�sS���4�	�X�E2o{��͍�yņ��w�c2�ȥj�����nswC.�쁒zrl���󦮕���9�\�T�Y{,����u���m��ڱ�)*���a�;�:�\nVY�-6eP�� p����[Fy-���Z�0eE�1�l��WYi'�Y�iI*��2$'���#��U,��]�P�o�ܴ]t�c��k(b���XV�*7:�lܻޓ:��X��ǨN�i(F��q�+*�M����xy��K�Ӎ��s&�0k��v02������:�د�ʺ �`הk�q��nWr�a*d�EΛy݅SM�[%K11\q������.���(��N�WUұ`dZI�k*�SL��t��;�J7���@���V����6h�MxZ�G���y#q�e���.��Z������`�y���pY��i�dn^[U�m�V�'k:��-^�PL��Wk�Cwۛ�����6M)32wt��r�o2�Ip�Ī3��o_Hc�yw�79�4���`���V��-��m����k�p7�N7}�u�]}W�[�ʷi>�nv���:Y�/''M��ʲF&8�WTf'o��."����{�r�J��ڛo[��E���Qw�^Ɔ�BղC��2�:]]J�w��n��UdÝ�y�e��.&�t�Z�\�A��{{�l��.�z�+97*TG�����k28K���+���l�/%�nue����JRWs�Zu�!��t�a�왨���[V靻��T�R��TEc�3���e�Qp:]'Ĝ{��J�l�Bή]�����5���:w�4S���Ig�X�C�o
����f�l���6�^����ו3K�E����⸾��-�mK0��kuV�\��w�Q*jk��Jm1亝Z�S��^�NGͶ�%`@qf���XX/\��ܬ�H"%��G���;)�L�Uǔ�M������a�\�@r�\i�K8BKG���L�b�����#�
-�ѦV�ugB8�:���������4!���-:�2�kN��^���NE�t��`���<���TdC��ť�7&�����l������H�'i�z4!}�"oP.2ݡY��+L��ݳ�@���4�8�kZnuE��:z��X:�"M󸡒ks�Ml�N͑H� $�I$�I$�I$�I$�I$�I$�GnK�P<�4�9�g=n�p�obVN�tCC6�;Q�7r��594�;]f�a6#֜=ug-S�O�m��pF��&�8b��H�{ܖ�q˙M\p`Y�P)ZCgXU{�aY�~v*mZg*E����V��ץ�*�g@�"�f#�2�w+Y+�o����n$GU�Uŀ4���)��L֪.��0.GWYZ�������ھ�M����*�Z�A*zw� �,sC���5�3UWd�ˮ��r=ԍn)�+�����<n7˵\m��+me�.�2�7J��KEV��-��n0�P������zX�v�ض�ie%'6�sp��;�0��Q��r�1fw0/�ܫwPm�ĵH9W|�LV&��MJ�do��>x��P�qI�P��;:С�tR��� ��`ǽ{�o���Y�G��'.
����	 �/��=�jU�{�]-��68���5����U���h�%�u/�3Y�!JWVp��9��*�J�L��x���������������9<8N<���Y�ӍJ��J��Wق�N�H��۳z��䌡OS�Sc��յ��=Zq�5����1 � ��H73od3*֝h2���*�+\27SDA
�G�+^ރu�t+IΐnbgE/���VSre޼�R�(*�U�Vv|����cv�SǕ۾P[Ǐo:i\aZ ��v����f�Uy3�6���wK�EM1::��]����'3
U�`[P��zL���g��V&-��T�s�Y�]�����p"��qzm�u{mm]@��N�_2m�'�ko��ϴ����չ�L�:��9(��f�To6����Uݶ󤺥M��mR�K��rqn�y}�ݛ4�
�@�˰o�bJ*��͞iԺ\��twǛ}�o��`x%��������Uk.��S���pc��Ǻ]�छ!:�5i���a�GR2]a5_��.}��S"D���u�F��+�PU�1��f滱��͈�`}��fV\s_j˻nm�s!�OC7�f�S��r����u�M��Vae[9w�-�QT�ꛪ�J�VOv�_v�����᝙m:Y<�۪��=�0'�P�Dw]��s�����.�P�W���wm��Nfʖ裱C����h�ζ^9���e�OML��]��LԷk(Ҕ4h����[Փ�\��z�)c���]VLu(��;\Xop�EK6�Q��Nm�S�w�tV��lZ�}�r�R����.�\y��|RJ�ۉа�[R������$5ή�J�Lf'�A�G��� ȭu�y���b��dګ��I4ΦW=��m�;��,O���a�U��gS]��m��*}�+���)�7)o}*���.�G�������m �&�ge�@�tGrUk�sB�����G����|M���U�X�ŝ���
X6S�b�J��j���賵�"ie�0b�#�xƷ}�m��R�³r�Y�fY���]��쓖\mbA�V{r�t��>�=�X~8kE* �]X�#�@���\.���mR�D�L���!?k�rT��ܚ�P.�ޗ�/�\}F��T��9B�U��Mo"�k(�8\��%L�dE�:#u\�ܾO**���f�ڱ��)_c6�[#T�\�f��[�Ƨ�D���W[v��t]��mk&�\��T�)�V!��]]
����]��D��b*wU�P�i��C����Y7|�e�']d���p�	(��ۇ����a�����,
��Yb�ۻ�F\Ӗ����0��RB�<{�ri��LTL��	<�ȹs�?'&�������8&L�W���o>VLv4MN�N�e�j�
j�V�xIj�S�ʽu�9h�wfZ�hhN���b�V@�����E��k]<Œ�\W2�[��w���ޔ�%����Ju�}&�U��Be�|{vͷ��F��Z�c�ʝj��z�8�����K�Ga�Z��^��nG(�Y�yT��2]]i� 9O����=�3�6��/"�\�o,�ĥM�>n�y���s476�h֍��:k>�
��I����V*r��o7��j�u6�����sI1I6����U��uCon��e��{����἗x ��[ �F��!��/r��vXOY"�����n�|Cc�u�Ru�M�ˠ5ұr����b�;9�&��w&u=3%�Ci�2�V�B\Go�\�g\�ͰNQ��h�i>�T�$!�MD�s�Eq��n]�X��I�ï0aq-b�`P���զ��jhE�V޻F�+�b"���,X��u2�N���N�%C�7�Q�,l���
�BV�w�v���-�_D9L3
�gZ���m��y%9�Jft�p�iiΡʖ�h0��2@WK���UԁӺ�jN��z�l��+�7/�2�;�.��2�UƆ�����V�sp1fS��9ēHR�û*�V�d�u"�a��l8�r���f_;|�H���1�á�YG��&�s�n���Zf�q��.
���6Q/joδ�]w��|�&a�c��^1�B��R��VE�����Ѿ��Y�l�m�UB��Q۴m����c�>�.|E�k#w)YvrB��y�Ts�K�L\��7l`a���$���`������u�on�dx�rE⠱A��5D�	Ο�oY��N8%eӷR��Ey���T���L󂃽Õ��b���9�E�cTYâٷ��*B1�9]�Ŝ���-DTF��p|iRn�h[�v��G[ܭ�a��IV79��/F�Ų�{n��ya#�6͗Q�$0��V!w	�'w�ݚV�+��+l�nF�yvPj�WP	��`�BZ�^V�b��U6�8lJ����-\���H�� �Κ`��ʨB�fh��=h2�@b{R��gZ�Vo�gm����cq��U���w�����Z�w4_�R�j��f�i鬳�mTcv�G����\�-�fǎ˰�M
,�*��u����C��68D�d���z�
#���HJ��rkze�E�.h�h���BM�����F���T�g^���� J�Q��}�]�A�䪔2�4.�X��q��G6�K��}�v�v�Q NcTn�����.Bx[w�@��˙�� �;`w��歚��%s����������Q���='i���T��]3u7-0K2S@*;0*��Յ���.�d�L�w��g-Mm��b�6)�Y'��v+�L��}��[��C�*Q�۹�:ȃ;T��.���b�#l��DlL�W�X�ܐU�s�qV��Th�\��w�;0+�m�kv�N;���E���}֝jf��Uӳ)�󮢻N2�\4)ڽ���Sr2��G�Ӿ}�[�^U:�%H��Vk�6����w�jCR���)�o��
^zt��ʮ����7zA�{A�H|���m嗐Ѐ�,������<k9Le���-�k�yIr�i>4�6�����+/r�]��J�Zl�'zqLΪ�&�ӣo�o�b�;��g3�����!0���s)�':�4���(8sXŲ���$��l��v���ٳӵM�C}D���{���A���(Ϋ�7��ȝ�<�m�_�� ˛����o�ˠke�ۏ��E؁%m�r������,Xv�Z�gX���R��*�e��&_#�����2Th�\&�2Ӫ�V��.�m��*7H�J^0o-��F��;�_e�R�!Dܷ���������TXˍ#D�y:�T�ᡒ��{�x�ձ�F���o��dR{�^�b��Fn�u��R�}o-҈�m��5���¡�	��Ē�:���(E���6~�/�^��sMˣ��:��Jގ[��>&;�Ǐ�c ]��%��\]����C&���7;�%����훽P�q�d"��X>ں䫲�)��Q�I2�m�w�,W,�o�z��:����%F�.�܃{�.����֩s��kU0���9���,�t�A�Z�'���uf�m�9��iH����wu����Z�A�2�<jb�,����d/+ZD=Z���_b<<4�0�R�C�V�����3��0ז�n��םsFt��BIE�_߁�i%>'�_A艉����w\_仰�uN `����tu6���������k�ۦ򃴉��*:�@�q7v��������9�;�������KϷ���ph����"���EA��~��kJğ���E�L�ލw�����͢3��L��yЫ<8gR��{����wce葨,\eGd�4��Wm����y��p����5���^�krp$��������wC��Qj�Z�L%�T/[��d[�Sm��J�j%R�����H��:�']�R�B^AEj[��)*�^�:���ӶWb�
�e����r1�v���3	khX%�e����C���ц�;�h� �k���='z}%�u��w~I�=��yT�Ѷ帥j�k�)�[m�(�s)��KB��ˍa��k��ZP�q�e�4��:.�mV���h�h[j���b���JPmA��K�QY�Fܳ:�CMt#*ѭ
�0��A�Q��ڲ�&5�-)G��#A��p\�˂�h�R�Z�Lq�K�[LL�U���ea��0��2�P�f"Ĺ��eQb�)jcf��*6���(��eJ�a�-R��ƚ�qeus���)QGY�m�����kJ��k��?�:�3�w�ۜ�.mw�L`Qq�j|�J�R]��$�+���y����	���;z7s�pVp�w�F��HF�8C4�Ott�{���4e��Dw:�,���v�*��.�Fb��M�Z�xAj��]c;]n�K�9ض�������w���t����c��)_N	�{����oq%�϶K����1�}	�`R�����ˡǵ��K<��Š��^Z�����̓�+��z�k&yҗT�Iw���g��W�f����v��ߤ,r�5��H�������S"8��❰
�÷�1��5��t��p�b�����[� ؓ�yf"ܙ�Rwo���kZ��U�Wr��Z����j/ݮ�|6������5�F9�9R�(6�=2�큊P4�����,�W���i�j��k٣Vtq��OJ��N8ݦ�z-��	-��HjG�T�Ї����en]�"CFFY����>UՂ'�0�jL<Y�Ŝk�
Qݱz�.d{���~��Ux�T�C-��ԗMl0�>Z��2�ү(]�N�ʡ�Rh2�Ň�/���e�[�P*���r�Ӆ+!t����4�h�&��3o��.��_�ĺ�����3��M�����4�r�w���$���Y�1`tǪ�>�|��?�q�UhoC�ͺ��W4]OZʺ3�V���ʰ���dl�Q��F�������g]c� �滜�}���Umj�]f��*�S��kt�D�ԍ\�;.�D�y�%*ǊgZ/z7��n��G$��p��]�I�l�����\�|j��`���Mr�6�MIgM�['��x�P��υ�Y��Mb#٨_Dxo`��9t&*dWRv��<6��UtGw-���VÏ)V�(N؆��#�Ը����-r��J���缛J�
j�����,$B���wq=�yI�U�l�Gԅv�Qe����Ԇ�qS�b�V욽e
���}	��a.!�k��dq�}n�:)�ѹf������|K�[Wu!�Ъx�W�`+ky�.�W�7;��F��WV>�c���{��O��Wյ	g5�_U��r�3����*�=D�t!Y�����z3�����S�����I>�H���2�����+ו6�I�ܖ�������Mש���5�8�%a�c��!c[�7��{;yJ�\痵����Q72��sp��>�iT9䈭x� H��6�v�����|֚gW�l{�%�9��egq��r^�7�!�p�pO{�6��.�&,7Y���oK{W���%�Tq�r:}�sU�Ln�h���ю��j�4�
'dn���q�d'��u��W뉺.=�d�磝��%���),���^Z��7�<�A���U]7]3����cQ����P��O��@�z�à3�uӔ&`VkK�u=ܤ�[�W(���ڊ�+`)���ڱ��� Y��(4��P�u�5/\�ùbrHq�i�	�Ɓ�;0�|m�ZN�.|]�{���٨k�fh�vm�]���A�d/^h�F5�r�Y��^�������{8�|#���vI�P�G���*���v��zyy���}Z���ltL��]����q����ZY2�2�ua���E�Y27��"�zNc�7�"��q�1�&A�.�{��n��Yی�ɠtL%�Y�E�xCb0�����9i�O<*U���>d1�-�ƅ���OgM�	f��)5ٳ{r�]X�;����nv�	��k�Qښ�1H�
�e'71�@'�U���U~�i�[��<��'���Y9kU���y��M�:��8'��T�B�#F�yD�6{�����=u1QsQN�"EN˲�+
�CE�T�FF��p��c!c��h�Lr��9\.>����طO�
M(�%h�y�ż}x؋�c��oh�k��d����4ٻ}wd%��wF8o5�q�W�]S�3"��j$ �Z=�x�?6&�2�����W��'��Ύ��/��M���w�삆d�,men��gs�C-��cp˭<�����V��!��Q�AD����5�ý��rzM?F}����^��V0�~|���e]]<",�v_��W�U���cF�6�,�ُ���|=�8Wzv���4�X��<�'���T�5F�P%����j�6�Fxq�G�轃j�V�����EZ1-�P�>\澔K�GohhT�gBk$�[�2�:�m�)m=Q�dk�����U�����p�=98:�X�s��#!z��~��zK�X���dS#�P�z���z����M(�5�������'HvC���B�p�p<����ڴFܼ���8B�Q~"��!�����ԏN2�+`qZ�51�[ybﴚw6�:�l��/Q$�{rs�\���$=(Z���q��{ඒ}\Qgo����715�Uk~�OT�d����Է%����j6 Z�� �@����zD, ]�w�|z빝OYB�F<w:�r��#8ߜ�%'����I��G���]�]f�O�<���Y�G6W�T�in>VG[1U'j�MћR��bw�o�W���9�]TyE�%^�Y�����W���^�����f����pH���zR�\Iae˶���T�H��.e]{��Σ:r�q�."���w����8�}FY�iγ�6��#�:H�:��b�P:c��vqE�f���LT�i�z�����R+]��zX��E*��'n`(?)7�-{'��=��sl���^�R��N[��ټ"��l�o���Cڎ��(s[�\������������v�긄��Zw���:oj5���U]� í�Pݝ���Ok�?oD}0'��s�������<"���޻���D��m�6�ns���!�������Qu�;��wewn���G`z��pIi�u��,�[WZ��9RSMY��$R��*���_e����[9u�xMg'tVۋ���7f�g��T����xu#��kNe�4�b�u"��d�W/7GL������˫��w����EH�-�V�n��,j�L��38[��t�j4�帽�6��h�NC���8�P�l��\Ýȋ3�`z��o(z�:�eZy�vgoY"���J.�"Y�����ov�;�{��M��&�۲��V��ޣjvW$���j�L���n��uЬ�Y��*ý��D���T`�}�qZ�T)]�۫X��ɐq�Mf]9N#����{S�?G�O�>�ߤ�4��ޱ�fp޻�j�����Ń��^��-��]w]�G2�0�\�M9Q;+k���i�Ob�R;Nm�^��g�ʋP5n�-��K.���Z��$�mZcj�n#]O�:��K�����xڮD��
)�m��G4��W�DxvSe�7A��-1�g�|��+�3\�wF-���s�Ӡ-�-/c�z�F�}+� ��y�*w[�LN����k駩�)c��t�X�B�Do���ρ���$ �&V�i�����|�(ݜF�����2�X5o^���mp	�kD#�T�����[��y(2�
�u�D����*�ou)v	י�ef���Y'�����[-E��Z��rխ�����[bVZ":B̥EVښ���`\h�2��D��1+**�JS�c+MR��`�hT[j���Tb���**Z4il�,m�2��b��iTY��e�FT�(�E+*QUUR���lh�c-,c��(��5�Y�6�m(�\��l��h¤P���r����V�sr��X�	J-E�m�ZՈ�K*T(�RQ-���1���JV�ZR�F�TQQh��F�Q-�9j�Z
�+X�kR��[J%Z�J�jՖ"!mjֶ��E�������3��j8��Kj������}���G���ii�,k��8��2<l�[j7E�|ydi)8����]q���z��=�ʗABP�n}�&���S<F�_u�j�>ſ���Ggϕ^,���>Y'�}FW|EI_�oDfG�)��з�{���{��4�x�^h��Ga{�N���|m�
�ho
�D���i�|��#�;�l��ɷ(����t�~T��ް}Y��9ռ�|��+D�ނ�y��[���T�x*0t����/�^df�îQu��F�s
]����G<`9J�L��j&;FTN��= �Be�j��uF���6 |5"8r�S"l�r`L»��0뜘F�b�3���,
s�I�_��ߥ��q��ey�N���+_ze�f�'�,��/FB���ji����2�����j�O��n��94:�δH~Q��d{�Gt,d0�^����LC]�����#Z.��^\��\�{�oX|UC�}�K�:�Kf� ��̲�x�_f��z�ސ���E���&p�ȤZB��s��]��֘M	��#���&��pB�}��6]n����ȁƼ��tG?>��
���&.�U]4����e.�m��H�>f�ۦ*�V��l߷�
�k��gz/ �,��v�Ӽ��+�>��F�$�D�igC�I��<����yP8GWU���400�T��U�̦�uD��ye�ǽ��T�]8���p�*S��9�A���h�ꞹw�N�Q�<Xt��r��3(�,wS^g�
w{�UO��|�-��ꃩ����S�_5�^����OQ'|��uq����W(8#b\��4x�#U������,�����Q�]���:�����M��k�׹�ּ�l�!�Ԙ��N���<d��@>�'I�O�1$;q����C����n��,T��e�b�*p�{�V�Q����0�ؔѵc��_s%]����dw/�Um܌kC�.	���K��ħ�3ﾡuU�T��u_T�������':Bg{�6�C�I�:`v!ĕ�x���g]}�;����<�a�@�;@�N��4�m����N�RN����̝���w�d����hI;`w���g�{��澒|öv��l�2Zd�	�l��:{B��'_XN٤�ݐ8�u̐��w�����>���'l��$逈C�k��x�jô����4�V��	�>Bz�ߖOSI%@8���u��7�k�}�|�;C���C�m���	���
@�|��<�ͲO�h�p��	�f}�ޛ�s߽װ;d8�ЛC��$>��I1�OI�N�<kv�Oil4�W�C��0�Z6�k^{�:����@�$�)�C9`��C��� �&�&�j�$���q�m��E�<`q>COi�]{�����;߿{����d������'�����=a6�Rq��C|�z�=d� ���&!s߷{��s߳�d4��'�>݁�i	�� z�Rz�*v���_Y��`(m �'d�(�q�=tj�:�|���&�m�t�>gi!��8��'��d6��$�P��Sl	��I8�x����}�ξ�U�zfds��ۯ���(R�v�E錕sK����g�?K�������W"��G�t4����d��p2ܱ���R]�Ou��W�ʯ���c�!<N3�)�3V�3�'H|�q�@���2M3]������Ϲ��@�&�ry`tɶM��06���I�I���I�T��$.o�Cl��>d<��'g�ߝ���=�{��������O=I6�8�M0<d�	�1��1���>N m�f�|�;ߝ��_��}ϻ�����OO)l=`0�<d�����N�8��$�Bq�Bi0��Sl��>G��l��}߾��IuC����v�l��������>d�!�o z���N!S�'�T��~79�w�9�:`|�2ɆY1�v�(z�d8��;��m�l:@6�ߔ�N�O�Y4Ì��xo�l�Z��Z�{�	�d:d�	'i8�d�� q�ա�OR|��6�XBq߽T��������O�O!<d���	���<�q>BgZ��l��q&0�ZCl#׼���s�Cěg�O@+'�P�$�N{��2m��T�遅��2q6�`�i5罿j���|��y�{��ě{aRC�>a8���$�2C���2��I�I&�<J�x��?7�;������
�>�mK�õ��c���7H�侍�Wf�JiU�,S��)z�X�~?w��h^�O�)C���]:�Ȯ�dY}l�-%�'�"�'�]}T��_�믲������>a�'̓��1m��3��$�� �G��;@�}o��y��s^}�d�M0!�>��2O�	�!��IR��Ԑ�$8��RO7H)8��T!O�ﯳ���{�{��!��8�$�{�&����3�CO�Ĝd�:O��������\����w�H)>d���M�I���������Ci�	����c!���C�$��]����}���`,��T4�ԓ\�dϾ�%d��8��&=0���!�	��b@�'H|�y\�ݽ{�;��u쁈}7d!�)�d0����9`tɶM}I�M2N&���&�'�S�Hl�\��y���p�!��Y;C�&��<I�݆$�a����'tn�q'O�&�&������w��Yֽ��L`4��I��� |ud>`,�T'i8���x� q����&r��ԝ>{d��_un�u������:a4�RJ��Hv�����L6�X���<:�!���$�Sl!�o q'O�<�^߷����~�H}5��q��t$=C�C�@�+v��=�@���m�l5�$5�ӊ��d�TMrХ\���O��[4L��8T�_��o[׎��+b<U��k�B�.�;�w'z��
*9����\��������|NUU;��x�6����I��i:`m�2N�x��& ZH�P���C�|�Ͻy�5׼�~�1���'i+i'N3���Ì�d6��Ch0��I�N&���޽��޹�l4��ABt�c��=����+'��	�d�@�n�m�<`,��0���vz����k�C���<g5Cā����>!ٔ�~��<�]�%�<�o��ڋC�x+zV!:�ב�Y�I���bSx؍�yy+:��B��;�S%.��;��,m��{ݾ�G��� �g�Oa�*J�!qK:N��H{N�e�[�ܼ�)�X�J+�)܈�#\mbX2)�f�F�-.��ގ&:���ڋ�"�*��	�;О}����&ؽ�d����]�&���M��<��.+&Ϳݕ?�Kge�g�e���m�'.��m���=�������ȡ�Gc��d=F�5�L�Iˡ.�5��}�>���˧k/��o�WλZ:�P��|3b�<�s�l�h�.{X˭�T�B�[�o��)��<��C�siw��c�3U҉%�p��4�T����8���2w�>����S&�=�7��SV���\ܓ�SCj�=�<��{�L�0�Z�VTn���ڽ�C���Gi�o���SZ'�v���lJ{�r.��Ou���2���'Ɇ4K���;hv���ݢ��x6�����
�%q��7'�s�7m�����k�(*���dI��W�_T��6������~���<B��2�f7�Vk�9��\R�9����QH�ʤ��x��#L�`��0��ɼ����_d닷NczQ�W�#*]�P��y�SNٸ�b��\l_a�}�[�F��[)ղ�g��z#O37j=������U8o����F����!
U�Â^��-��# ���zm�/>�f�Ӽ�ṡ͚eoQ�{pK,���r�,��s�~c����ֵR�eP��ofe��VGbN��f�?x�y�{r��=؟uq�Wt��}	f;�Z껭�o��:R_��G��JOU���� �̸��c��E��#�8F�$�/n���8]Y�A�f�Ʒ�?���O"f�˲�T,��rU�$Jwt�g�ӎퟩ:KM%}i��^a>љ�ǽ��*@�&�8��L9ʥm�T��8N������z�eR��7 3@~>�� h�04�7ǃ�*���|b&Wd[x���{ѯ}�cP�4�D]�(�mx�Ө,����J/>��Q�S��ѫ��qA���z��_P����N�-��&d��+�3w�r鲇-
7B+��B�1�Z�Ê�{ </��VAC��]�:����[7�i��+L�x.c��Z��'�ZrKJPԵ��m!��������P��kh������(�\���u�u��K��R�j�Hp��k&�Z���jr�~X*��r���V��f��Jɪ��i۵l�WKw��e�u���6��6�����u�u���<���ѝ
xҠ��*�y�+	��ƔX���v����͎�>@����z	E]�.VU��gv��)����J�r�Xn�5��֙�pd<���Ӂ^�w�{d�;�|�7�L7n[�]�Pܭʻ"�5����e���V[T9It��Y;Cψ�7� ��#U���PGP��}�V����ɾ�vr�C���6jL=�P��]qw9�m��1���f�(�ŗ�����={(.�4�z���-���}/;Ϳ��S��!�ˠ�۫�3�y���D0�z$w�b�V]���\�M�̘�t�����μv�}#=�9f�2�Vu#Sn՞ڜ,p�qj���3�J=���d�l_wU�opv�R�qe�*Nh*=�hŧ���Bغ�^�V�hM�U���eyˤ�>Ye-�U����݈�:�c��#ż�����N)0#�ԏs����)`��N�f�o�Y[}\�ܑ���W[�����]�gl�w�ɔu�C)R���]d;�y��cWwR�����H�~��&��ϳ+l�
�Z�AЩ���(Z�����H�sEAȴ�(��´*�D�Zʫl%����	m��+ZR�V%�����*FѣE��L���UEkDB���nR�V�Ơ8�m��I-�%KiYm���µ�ڢ5�X,�R���Tl����D-�QVVkZ��Y*,	JJ�Z��B�̶.5R�32�N4�Ʋ�"�ڌb![i-,��jT��1��RJ���,-i%-�[H��(�m�\C�ڲ��b����Ш5�kPik�����
��+T�EaV�IRV�h�d-�33bd��W~w�uv��3fT١x5��IM��ݥ��8d�O�O��UW���D����?nÚ��%�1��Q�\�-���Bz��O�g?�X��Kk�,��T~�S~�CK�y^����r��z��^�:j6>���&ϭ`��(��^ٸ� �Vό�6�,(=��i���{i�B�E;�8��T�i9U�[���8��k�m��l���5K�t}�T��N�)9j���xV	Q,��e�hĴnr��w��ư%��F+�8��t6�8�UH�&�c�*�י���>�뮔3��>��O����_F.�K�J�f��E�\(�{6i����&�^+'�*l�z'�~��ﾯ���:пh'��kNF��u붺�7EU���tk-F����v��w!�Ao��<��mb`Ɲ3�"�^b���dO|�k�{z���i��3t�xx�k�tq�6�<�G��ƭ��F�y�}y]��6��[����l�o3�=4�-��"�`5p�o�Ɵ��`�lZ�̆z����1���:�J/��fV7�;J��k��v�;�}��b�i�؀S�@�7��xZ������7y�*� �\|i���G��o����F�L��{/z�>�T��ygO!=[H�+���z"=7�����������m�O|�>�޾�v_����t��U��P�q	������}�^DGt���5yP�3OY�<x��J���'X�U wW��{R�����d&�5᎛MW�m[rCR]�(w��l�U���C��qJ�r�|��T%�(л:gãg&�޳�b�5���h�T�����2�Z�����O�F��[9���H�L<G�yj�i�Gm��|=�<,�|�,�2����&���]D�FB5P�볝]ٷ8�J���\��j�v{�_`Ml�Q�҅�a�a$W)U�\8��""=�z�ZV�#/T��f���7��B0��q���������k%�}KI�[��j�z����:��"����5'v-��%�,9Ӽ�P{���}�m�ζ]xi^�g4��k=��G��W�h]�����J���n�i��'JɄsm�։Ȥ�+r���x�qs%m�{��XoNS���,�:	�!�5&F-j'��=C�׎y�P����)�7p��M�d�����M^�`˅�dUҗOr��[K8�pTO�#}^l.ɻ)���:����G2��'>���G��(�\?�q�{���wfi� Pk���gz�������2v�b��Y}�e�K��݀��Tr�N��r�M��l�\���{C���vYj�v"��_J��h)_g�|�m{��f�	��W:|+|�g��h~?*61�k�E�VT}�v�犆���O�s�����}�즸�9�|2�.1f�.����#g����|��� �.�
6v-zj�gj�b����	:��hD�`��̷娭O9�H�ߒlsu��X"��`���b٬�l���po4.P;U�PQVT��Nu�I(����q}�Dz#р�ڷ�i�F�s��SBw�#GZޜ��2�me�;��mTn��#k]һmrVCؽ��.zu�Ԏ6R��x��.�&N�P૭�6�3���r��n/>���E�,�§ᎃ�aT��tu�J�y9gy��ڻ��[+��v���핪b�\�i>!�rc����mwOo|Ue'���Tձ�l���O�Y�7��l���6up+=O�*�����q����pf�C²��ǟy5c��hTTq����T��S��w�%9�,X�E��e^��X�Ad�/,��s?>������ ׉<�x�}�=�S�b�{[���O��Q�<�iY�=@y�y���q���a/{T�+�C�93U�+�m�~��z��0�ݷ���$s��+�N��\yjO��Hk��Dr~�e��V�&{��|�ݞ5����F�Mv�>�x��ʢ���=�k�>��O���F�G>���59��";X=��3�d�%{��*m?Yv�U�_���e���.��� �Ȩ�:Y��Qn
1�7D����xR&`i�ٴ�m��U�:v�sz�J��ҮO���fD6�h�%�n�5`���'�-,�v�.���_}U���wZlu��3��꺫b4Ȍbg)��6kS�\\���B���U>yβ�)�GD;�Po��xg=���{/j{��۬�
8QM3}N���ukڻ�Qe�aݬo@�i�W�������5�=�7�>���
����,0kN�$/;}Wu�r�r3k���Z�J����U�؅������ۨ�K�������o�<��i�7H��)q�jϵ2�?�;�zc:�A��u��*�S>��=0��T�{Uv(�=�2K�<�-�o%�u�',]�U�]�q�C�n�KJ��-U�Q�OȚ�lg#R�ξ��/�ޏ{�˓*���g�L>����Iq$����^���0�NoOoF�:������줅9��\OA�LN�[y��������*5�lF�˶x铵q�)��FToJ�ƴ��ڌb:�0��k����Oh&�N���C�b�����d+��|�)t[�ѳ���W�U7�[��*����f�����(�[��}osz�/4�v�{�+�۔�>��o�b�.���<Eվ�;xm:%�^��k������.�NR���͵���f�
Z�W"����w"�΂��Z%q{�X��]Z���|Js�����KA�������|k&&|V�jbș�
{�!j�t;�{k�ǵ��/��2��H�<Q���V�C�`����ܱt(�uŔ�WI�C�rL��N��f��]Ja���J@�~��7��RXt鎠>�&_��FKf+*��6nzK�pb�a�X��!�v�狑\ٗ�S2 ���C��N1��ò�"��;41Ž�u[�a�����Dѣ�������+ơ�):K�����*�0HRPr�*�̠��G)ZCO�Ӕ��)��ӷ����pk����o�_�7��w�{w��]�쳘(�]^`���
���q�C8ҕ��z?h�~ݸ�}Ր��ӳ�p����m)����CB�*Į��VlI��8�Xya6L$�Lr���+�9��ԥf�{m��i���i�S��\Sm�}��[��;h>�>�;y��T�ܢn��
����q�tfZ�7c
�u�H�t�T&|���.ڙ0>�h�P</$�X�F��.�sTu�
	�t�n�;"��g�o�nͭ� T�m��/E�� �ph�ڨ#�I�l�4N���uI���VF�i�����ՉT�gP����b��|��IT��.����u�~H���;�Qu��1&�;�J��ew]� Z�"��)t6���
����qu�_I����b�J��)�M�f֠�W�n3Y:��س��]P�΢!�16wD���g��W���]Y|gu*�����T���C'mԩv�/�3����_�Br�� ��u��
6����<���˲��=���s!���kc�Ʀv N>{�i�ή�x���B�6�_[�)�e��0[&>��s����;��ÖN�����Ը��vf�N���7�w��4f\�%]k��.��
]3I�bW�]�m�j�V�t-�IuB6��'��73�����$�OZBZ�F!�v寖]�H��"�'�w�9tKj�F��\���-,2�tY9�b�㽔�w:R��;��Na�ѹ�)b����/��pa�!vV;�'�'�
�j��G۶s;Wkv���%ݺ�v:��|�e,鷤X���)-u%�V���/��u|�:���s��ܱ�]볛���R�M>�LB�V�ʂ�Ҷ�B�%mdX%��`�QKiPQ�%������LL@ph"%�m���T`,Z�-(�YUR��T�J�+m���+��ք�FьP��p�IP-������&�$���m���,*6�i�`��T��R�
�6��
�m2����X�����Qb�YLaX,XQ,���kAV噍m�Ed�j��Fڅ�E+V�J���km�����h�������e2�+��U�ڭki*VV"��u�뮾��&m6o�^�	E�d�!�o�0B��N���i_����̛M�S�u�E���GVX�����#��"~�Y��Uj���3�M<��c��D)7��؋�bc�����r�|��#:@�"���
6k��`�5�f
/,�{�"�>D"��+���"$fq�3mUv$�fM��e`�dY�{<f*ht��⩦�}s9�X�<_�陬Q�b�{U�(�����y�^�]�#�/��S��yY���-V��#�䛹�����'@�<꣫)j��+�����Bʯn���$�����Z���ت��^�*�r��Z�C]1�a��Cq����r�b�A+.J��ַ�6�!W١NF��^R,,O�vr���;[����k8ۛt��+Zq_D�؇q6似�:��""=��ι�ɓ0�H�Ｉ;�_.�$��/���옍"���2$�t�U�Ʀzb:oC���+7�,M^��V8s��Q�A�Aq���(�kX�}[я=��j�K�z\�5���U1�ǈ�GV���FwU���N���)0�^��ǥZ��fSJy����2���}oHv�x��#�3�'�+%����:�sgV߷D�P�E_�`�{W��*�5��';��R��H���a�ڡӣʋ���8bOm�1�?vy�8|~�N�W=>ŧH
�"���<�1�ov��R�鯌��A���uoyq����z��xY�䲌�,��9�] ��*.�q0��5��!�@��Ӄ:N=���^�8P����2�������zz�Zg�a�Ma'������Sz�]Eo���[CK�Dn�܉�/�슪���c
U�Q��v��tt�%p�Qi�='�E���c ��5^�*�罓��܀[���Ȁz��XF�Ѹ�׺k!�v��7f1d��e���8MH����{������#F�a��Dp�񲍑�����JYUY�Y=K�n�o���&�S>7k�������y��'�/��,��f��l%�LဏĊ��f\��5�����$�
Ţ"7�W�;;6L\h�л�Yx���}��;�J;�x�9����J����8nz��|;˄vg_y|��p�^�#]n�O����r���{7J�+c�'��k�b��]�tn�uSnQ}}z7�!�t�ɋ��T˒�\b���{ރ�ɗ��'�71_�Sz�i�q���b�Jk�z��K����0���6S|C�I6x�ذ��zu��Iz����ʁA���'d�*5�kI�S�B�<�f�tY ���u�9.�����뮵�"}��:��u�:�٬�����)�"g�H�.�WV���4{���Տ��F��F�,4�B�-����b��P�~�tn�ϖ��xt�F�gM��6Y�_m�V�P�<��~WkM���ƾ�ʷX���։VOg�Y>�@�1���mz�w��D���s���$�g�tىj'*;!��e�h/y���4,��v�_{6���bb�_HwjgWT��hܗ�R)��n���!M���菣W]9��9ZX�s����e�r�7�������c%�8�o��M~k˴����$9�l��ҵi͗;)���ӟ ��X�zqx�����ߡu�Q���CX�gLK�a^�����뾚�T�o��Q3DD�V��g�ɞb8�*��{��0�͑Oَ����1|ǋ�MƇz��ΕmUN�i�W���kǆbf��ء�!-`!U����o0B�x!P���90���ZyV&r�����ȃP�.ib��J�PDL� ]�w�T����L���z�ϭi�9�]|��k�^H��v9 t��r2��^1��������lү�=�ii7�n�)L;*mj�"��a��c�̗S
��y�q����_-�fv.�����u(���I��}�{���Z�S�X3��@�b|�.�q��"���ܕ��*�|�f&`�ʉ�@�!�"#:�6�(�ʓ�������/��Tl�{�S\x���:G�=:�o.�������B�K_]#�t��E�9܉A�M��D�|�I�5�XR���j:�M-��:�f�V<jUr'"c����3�<%w�;H��c����<]��m����AO�x���+�|��l�Ql���FK��� S0GK�0z.8�G���AeW��"�Ȋ,E���e!�ZV�ݪ�OfU2!�p��-"����Fya��^�y��#vy$,�fɭYVT�X��Z�:/��K��z�N�7��~ܬ�ٌ�L��%4�ø���>h1�	H��;�������n�֏}��]�n}�)ɿ�gF��a�o�[z\�b��:���f���(t���S�5�슬��9շ]�K� ���������?[�1 ���o�靯���8h�|��^;Hh,Eş���.#�O�7���e~��P�E��OZ����.�2�Noe�	��Oj�13+x�`F�!T���ln�A�e�[6�x/UТ4�����2(�~�Y	g�������8x_<2��5��O-���/�-�������!�_����qi�>�($�jL��)h��ɓ�}^F��g�Z#=��12�!����D˳<�V�����+�Ʌ�˼U��q�w�WTt��kd�K���w�:��$uM}�5��B�c)Hpk5�Or�⦄-_G��,�$�G�j+�����a�_#���]�67j��ݝN=>>����5��Yƽ�'�޼�mMV��z:T��.ab����Ld�����x=)����3D͡�8�<���(�m�0�3/���a��ˈNP�_0��!�y#�w�*�U�N�my�য.��u�S�Daa&Α�Y�������!�8u�EI�C%�L��*|�m�L�W����G��@����Ij����Jݽr�ӧ��;%�|�B	dg����wt�G��,�U���5*����l�o�dx�v��]n�C/�"K��j�}�<TmjV8��f�G��SnPd35��B�ַ5�[���U���8d�Y�x���{ށ��Lw��̩3�:zl��,�ci6=�3�ԾJcsjW�O���31(EpH�S�`�h�b
��fK�7վ��>"�4C��P$(�g�+���K��wc�W�^�mѝ�$!��#��r+ j�����z<a�n�PY�b��#���3�3��
�(D�<-kZmov�Y��Õ+z���P#cD���UE7oxƺy�F�Ϻb{��Q`Zl��G	?a�Mp���6��:I��.��9t�W�����I�1z"�̝Z�`K���0dLm]]��#X�s�D[��"fy��j�p�e�l���=�Pv�l��y
���Α�v��P�u]�f"����c�K�g�����C�v7Y1j)���Su�Q���Q���1i<������c��z��'���5@|F��E��fGXrQ��N��ۊpj��TC��G�u�kl�@�T9L+�{�̧��Z��t�����Sp����[��=���s�D�4C7�bo�����D{P�-on�mz�j���ѿ�8x�0�Do*��QV��s��BY׳r&��X�Dl H��Ѝ��
4���_���,���6>�dYw���0c�t�&.�����D{�ն�|��.�yLB�Y�a1��0�kz����޳2�oo'O9�߷���1�хۍ��+��`�VV��s��r�⎑�R��� ��[$��ʗVc�ğ�*|��w�uBE��W]T)2�34Ͳ�l繇2�h.?�UТ�Y%����/9غ7�3`��4')VM��Kz}s�
	��v�e����4.n�3z�qۜ�ٗ�ky��a��w]�T�����(��|���0^2N(.�F���U�^h���9]�z��.3ȸlg�c������72a�sC:jy�a�)��f�����Mwjڴ�X
��ML2�ͤx�p])�~-�a�j�EJق#ȼ·B�fZ4yi���Ł�묋���H���˭�'O]�Jgʭ��*k�M̭&�o�7Y��!�W>}���X�*q.pW���I6��o9_%������I_��+ѯ����x�����uo4�M���B�ՍX�6���oqY[��tִ";|��ْi�*cKߋʒ�XV��,_V��w2��ī������E&�}����Z.�R��X��*�	x��F�OQ�q)qcl������i���.�K:waS��D�ƻ��{v˽���R�İ#ԋ�cfn�F3`��+c�����u|����>��"���ðWU��bQ(�S{���K9�4ڵ��6_^�1�"��Έo8c���(pR��%��;CU[.M|���mh�����h�-${��Q�j���@��u�+�]b�P�[j�gL�1l�v�7�����k��-x����u�g�8��PE���֢�ҩYR�bT�e1������+����	P��E �eX�@��f1��Ut�Y�e*���H�J������1D�[E��
&[�Edua��Md*U`,*
Tb��c5�V,��d0`��Y`,�̴]2��
��M$�RE�,�"!XUA�~[��z}�<�uε��/�;َ��KmwJ9"�r���s�����M���b�U���U��ձu��li<���2�g��:��Ֆ��u
^"bIx��0���d^��d�U��fOoi��Jt��7�׾�w�kUH�Q5)�"DS1~���G1�bW��[�%��rn{H������}dm|�[�z+�K�*����!�Ő�CB*{UGJ��ɓ�+ˏ]@���<��ˢ<Z^��M��
�B����xf ��f��Ug���^0M|h��������kJ��~���V�4��C
(�� �{���o�]���=�R�z5��ed���L~Kѐ�}QU5n��_K53
�	9�K��*�%z���_d�
=�H��9K1�DD���fn�y��r�ju�V'�1C6V	�>�5���K�c9I$����Xd��9�=�W�f�A�����S1s�Vϫ���-ɾא��{��txcZ|t��ׇN=��z���v�
��>�
��SRf�('|��Q��1�XRS�C��'��"��˝��Ba��dH��9�`������G��T f*rx��`]E�փ:�b�T�5��G9g���yӼS;��J�{q�О����r7ϺfF��s��&a9P�]JY�N��������):C���'1��1�c�ƣ"vS:2�����V:�
���NP!_��\p�9�Ѿ�'9��a��n8E��)���hx��l����x^�X�]z��A,����b��L�@�\f\ �;���r��Ζ�>1�og>)�p.��.�D���W�z&�\㜘�&b������Ps�l�ɂxTc�[[��;��4���7�����k׈��mz��k�s�QF�=兂,엵�����˥���ӊy����N���#}�^џ��ʯG����.!���l��X�9hBǱ����B�q��ޞj�X3�=�3 :�C�3�ܙ�����U�޾��配�-Y��4F:�"��z��u;}yiT���8}���k���-VXHv�r�vC��t��'��{:����#Ռd��?M�3W՘�f�J�y}��j�(�{��d�W�T� �_Q�qU�	k�~=z��.խ0�b�2K��*��E杖�7�㙹�,n*szźj�2�YW���F@e^iq^b���Z���<N/���Sn�2r\���J4f>�1�&vc��OL϶����S���K}{�\ѧ�7E����m�'�]��K9�;�
,ғ=;1�uS ��u�������@�f�uK�f�%��0�uJ�Ӫop�;�]wO]�t�u�-}Kt�:&*	�SDd��D�k��رSr�ݢo�#uN�qieDA|y`�����>�{�U���w�G������.�w۞銳��!�y{�e. ���Uh�c��<~V���GM�~�f�c$p2�@����C"7ܫ�^�������'�'���ت�.'�^��׻[7�sʒ2��]��%5��L�MX^�yr�]:W���˹�q�5Y�81(��&6�#SjΠrK��J���UY��~WDa���!�8�0<�d�Ld�!z��?��|p������~�>�?1�/��e�"�t��\�	����TU��;�2�]EC���.cdʑ0n)SeW���֦�P)��T��Ӳ��p�{ɦx{v���x���_m��=�4OR�	!�b�������v��d�~�)ܫ�v�ś�f��*��C��O�J��i�$��ީ���Sk��i��Ҳ�t��5�g���sfB����dp3T��3�Ҙً���Iq�N�kMl_�"jvS�.��c�W�hu�A�]�H�y��b�i<�
c_1�<{G::g��U`/��v���%B��h�T�X������p9)>�Oo��#�|�;������N]��ۉ�Ǘw3Q�v��%~{Ѣ�Zq\��NH�ٰ+��#f�sQ>�^���q&mBX[&"�S��h�4~��8&�Hh,Eş�xy�����칅������D��t�3q]��[��`ɾBO^��"�Tڗ^������R������0#e�V�oe`��>���S�����3����(�:1Q��ۃ�� ��xe G�5��-<@Z��ev�Vk�t���/�d��ixäW�ʖ���0���t���:p�D�?C�/�0�3U��v�~3�l}U[ۑQ�f%�ost�4q�����lx��%׻3+���ŰƯ��ZX�1���dA��K��͜�Є�w4j����]ׅ^��ٌ!�EW�Z+(=�D���q	K��5��ej�+d�
��'����0�9�dV Ծ�g�r}�=�,��?h�5
�%J����U
���˂����
��=ծ�L(�ᢸ\���6Dc3Q�3�o�
�w;"��t>4jz����C�4��a�>0bwmtĦ�}}�>G܂�p�M�c�b������*
�Z�l���3C>"Go�a���ό���Wr�z��a�QQ1�9��f����u���#+i�x�+{-����w��]p�쮩�jcdޛ�MLL�[�u8�����[��ؖ��;9���B�t�Z�:FHg��z��2���4<[B16�i��D>�6!�|�b�˿kp�\m��$A�y9*M�5��oE�.I!Ƭ0G|�]����K�u�٭*�F��=��t��y�vl�Խ;�2�kd�[ʎ�E��0��Js�7RrvR���A��\�LW� 𙌚��|Rzut�#�gܙ~C�zqF�6���ϔ#v�k �И�#�uu��P�"8�v����6sheo#��12tC�s��
W+�U�TTV�y�o+l�.�r�8t��{=8�D,K�1����*{��st��9}KͯP��sX'H5��2�V��=j�݄��!����E�����΢~�kL��۵�v�Ԭu)ȘF<���%�C���x����]�:��ֈd(����:iS`����Y)&U�{}��dTTz���̟Syv�#<�;1�Euz��twG$ڌ;�`���'� �Xn�,�WqΎWj���r�lM����M���f�f��[ɋjڱm$�3x����}ͶȨ���Uҥ��:Wf�S~{FL�v2}�uj�G�y��%�r��@�^_|6��LW�mK�<�x��e꺀�;F�"��=_Fk`�!��C�����Nvn+��j��Q_4~���nETC�G��ř:���"ѥ��S�Ey���+0"��Uq%��G+vl4N�=Hy�~:�O=�daE���������A��<&1��ac�Ξ-��Ϗ��0^�8��(��2���{�_�U�w�ͽ�V�d���"���%�_ D�������x���m����^�m{��G���8h�C_H^!�ƒ�j��q?ad?W������f��Z�rY���	9�$%+����}6{ݠE��	ȵ�ف�7�IQM����兜�՜�4.]4��]gr*=oo=��tv�v�=_.�'���(ʝ8j��N��ͦ;/O,�2�AA�����)S~4�*4GO���QWe�UPf)7������2X�;C}��#L�Kv9R��{�=!��"r�C�y�]�x����H�73=��&!�(�Դ��@ܿ]W,'v�ϳm��>�B���^mՑf#|�ɯ�R��YΒʧ�M��[�����qB	���һ��o�-�yG�}S����uV�a�h��R�Q�Y�%UC�kz��!;���O�}P4՜��|(�w��*��pg��P�5��Íic�n_�k�٧�������g��L����/2��6տ����v��<�̃:��T�I����V�h�����f)܄:X%�9���00'"8�6���jn$����fj@���i��Gך�q*�X�}7l��Ǜo9��tJ/p%<��HL��!X�畆�b$�fY�,a��[����j�.�����/geN��iIL[���&
]��B)��R�u�P�ڭ��#sNe,�E.P�]	���wv�Tyw������"��&��ˤ���g�J��7�*�/�-ia9M�um����ϏQj�PW�n�ǟoL�v8s)�b',ku�uM;PP�v�9���KLkVry�75X�PcfT���8�d�H�b��cmKʡv/����Ώ��eDW��ō7�e��L5Yc{3��d�1
v�f��p �b���R��������-�i�����g)�Y�:u^��]w^+���ke�>�3D�Î��PU��zŜw��eˤgT�ڶ��eg*^�:�\t3]^^��4��uk���9e��r�K��WaRK������.�ݚ������l��I:Jj|6�N/�@�G��іi9�NC�S(�^�Ѳ�ư����O�Ũ�t@ز�8�H�p7z�=����2��v2:��T���O�{�WqX{�,֍�:8�M^Θ�=��R�`/�&Cڽ}ό:rt���������joU�Y�m�f���V�k���U���(�U�@�*�F"E!U�����E�
AT
ʦ6+l��\`(�6��DR,��UQHE���,��DbE#�\�[eL@�5�������KAE�eB("�Zf1+��Rj�,Y �(��`"B) i�!�
Ȍ�	Kd�33詁1v*c����w��+��eeV�Y4h�����������k���z ���S.L�?S׈���Vf�7&c��P=�'N����W�ge˕>�Z��?j����g'4A2��J�o^缔�ᩞ#ܭ�y�:EGxl�d�,��������; B�t�T�AD���D���D{*W��6~�u�!R��
k�B�*(��u)М8j�-���4�7���=�s^ᇷ��1K���v�e��l�����M�O�~xp��~Vt����
7U�z��h�Ak�<��2A��\c��	ֆQ����D���{�!�hB��Θg�9Qs���Ӹը�EBb"�s�����u���u����j����%��Rq��Y�W�T�Oz�xCXs/��I@\A�ݬ�V��<���	����]��t\��@�9?>�P���Cu�T�]���.Ya��l��~٩���Wlr������"Z&?#�<�t�5�P@�}`��e����~�QJ��^.,8`�,�{�^�}��<|+X`ٹs��#�@�ʚ�;���o��@�]�D��a��4E}��v���@�;�����jYAJ�"L�*��L",���D��8�f�g�HGM;��]B�����^�1r�)K,O[���j�t�vyF�0=�y�3o-��j�bQv�p�o�Ɓ%�5c�1)ҟL��]��*��^7�[������Z����uu	Kŉ���҄srkC�����P�˚w�v�OS����etLH��wR(���]�UsÎ:�u�k�����:!B��}7wYt�X&t�ٽ���:�W�u���F��&zLž�+ ��&*�b�D%/�D<o�:�u�7|�"g�G�L������䆶�<���6�k%1�D�B:iS1�b}幼��kj�M�g�G]<4GjE�0�j��T��{�j�Z���KM9���������3�B�D�/Y���	`9 ߘgHf��X]��g��w�W��D>�����AM`,�!�շ̙��y7�q�!��E!*��h�/R7T��(�]��u��M���T)SdC�FLd�O@2ɣ�Ƅ\x�Za�(~KX�-j�Fdc�����{բLJ��뎳{��Ks+���
�Y�5�<o^�:�w\����9.��ue3�{��y�:��ʩH�T�N]�q���U5���W^��|r��D���ό��XR��˾���}�Sr DY�)T2=�=���"xRٜ����7�j'�Ĉ~B�<\��.�D��POyw]�]͚
�	��>�#"rL��� ���sժ�Jd�� ���M���x���6��{J2�J��250�歞�9u��	� �)�*$ʕ0w_dX�͞�~�?�u�i�Y�/��澲6���U)Y��C��d��Nb���:�6"���J����_=�Ԃ��0������hY~^ V*�ǟ<�Yl��\]�(��b�6r'g&�a�^z��W�ۜOo.��C��}Ӂqh&>���_c[]72HN��:&���J'���Y���i|�|�#eԗ������@�۪��W�H�~@n&aEGϟ��r�ܾ��	;V��u{�0E����zG�i�=Kkr��Oc:�ź�3z#r�6=�����rzO�����ҽ��(�0�F��d5��x`��xQ�㧈�$5Ů^`�ᖬ�/�8��c��x��X����vz�sj�4�ZX:~�M���, �>6z�m�n�&�ޥäȗB@!�4�h�Xn�؁�پ��i����!z���-,ygY"Ș�������~�_�`�s&Zq�I�0���TQO�\r��+��t�R\G���0�V�*sya8�}���e�1Uܻ�<��ca�ab��t-�J'��\m�a�o���Y�I���}1��)g"�w{	��!�}������١zx��m~|l��o��O�(ЈO(����쑽~4��r��^E�o�8D6��|p�C��v���M\���3M�y������ C8Ѕ>�����iN���V|}�����W�W-0b����0r+���}I{r"��R��u.]��MԺ<��g]��8>��*?D��!�F�vCrޘ)�o�u������fx�=k�di��LJ���g�
Г�4��N��{Jꎚ��*$��3��&$��99����y�vr|��EOk�Ӈ�I�x����,^d���	�خPr�Ȝ�!J`�q4(J����N�li9>ܜQ��/�m���F�e� ����J�ֳ��wk���FeЕi��	�K\i쟟U���V1�á3�;�lE��f���{�L�YskUc�K뙓-�xD�H��=����ش�_*7'��u����sW�Ogh�)��y�������$��V��G==>/P'tD��8���(���*�3P�q
V�>�*��Q�]�p�Nh$Wh���)�Bf��"0z&FdDЄ��ē<�YJ�P�s��X��әB�tʗN��U�K����.vm���ᔼ��T@��9��iM�t�.��rl��|��/KL_.5�zK�WC=˥w�z�s�h3�B����Z4�Ն�L!��Ug5v�ׂ�U���n�&Zy��Xn�`�z�b�S�w�p]e�G'#���,Q�4�9�[%���\J���jӄ��sD)���N���*z'�c:�^��jٺ�"�D>C_�a�0��D���m߳\�*���طOoX��W0��a�b�,�<e)|g���׍z�fωņ�P��Z�{�]������*H
aT��˫��c�4�����8<Q��J�mo<s��=�*nfcX�t�)��X�C_������Gg�9��݈�k�)F�z���X�:v��J�����{���� �c��b������Ǫ�+\O;��#�ZK����ǈ�uy!�H֬�~BI����v0���E���x��\G��W ������➧Y��0��<�j��4[A�t��k;yl(��mC]|f;p�it�H�E�_`{���g.�nh�x�w�J9�U_}|�-S��xD`���f�T�ԟ��z�]^�1k5ʁ۽��G�c���Ck�*�-�ܨT�.u�D��v�&oE�I�~7^���X���R�g��kz�a���یu�8@Z�E~�k���=����Ѳ���9qq��70�(�*ͮ�k��/Xo�Go��,���w�!�|g��,+3ss�B<���<w�����1DiMY�g}�"M*}[�&'D>/�"�鸠gX��d��0� z����|F�C'=6���>N	�VN�tx�,vz�*\��3�%�?#�+3}�t�iy-��U�O�oE�ӓi]��nD���	�G6�.��b��n>��١)�<f�̹],.�&�Τ�U%��q'?*����q,�v����s|*j8A@!3��g'@�Z�ұv��`E �%I�#a��3��t3�:�R��l;��D��Ñ�d��ɛ񀦈��B�V\��m�h��Ц2fzc'�BzbtD�[�s��,�º��oq!��7'�h���^XvD��� �f[�oN�Aʂ#��h��ҠG����H'/�����t����|x�j��BG��bS���=��Mwl�;90�
�B"�3��˚��P�7�W����6 �]d3�[0�2Y��MLl��9�$�ɶV��>(�*}�1<Ø�e!�^:sP�]u�d�� a�)���g05��b^�غ���U�ɽ�����fD�%R̫�yZ�K���)��bL�+r�F��,Z����c���K2�O`���'8_����f��6�u-��Jg>s��n8pqۼ����-/����4��,(�]�ۖ���r�nU��Qk����56��[I�t�9C���V�Yd�ɦP�Ğ��9�<X�5,�y�Q��5�Cz����pCYF�X˭����QL���A��"̭$$�h��,ܱ}y�^:���`�1T�bĺ�"�m��+�9#'9(i�u��$���#u��jۋ:�槮��u-�#�3�v��ww�)Wgg>u�4X������6+K{W\Փ	H�Uz��O�]CD*�h�HuU��	�I<���ɦ������&�ݕ}���0Y7jδ;!��$����y�o#�f]:�w	�qJ��f�������l׹W��>�<{�����J�5؎�W2��Q�Q�:2b$�S��(�E�r;�/��7W��^5�n��f])�;��R�ѢN�'{Vi�[��ټ���XI��0���D�A	[+�Sj�{8�/�c�L~�HcS�i���<����=�`#jX���Y�N</�����'4I�L��.Z�e�q�CS�zGwL���%x���{����V�<��r�+���Y��/�ܝ1�{w�=5��J��C0k�㹋@1I���C#�|Ĝ�\���dѪ���y�_9����g<�:@� V*��^�°� ���Y��AN%a+���!:C5aY%a+$�[m�Krٚ�I�Ht��TP������*��d�!�"��* �-IFc�(DE�2V�Pĕ��LP����	��\�G�`x`��0�s\lL�tV�*@��x���EV����q/����hG*Ƭ,E��BoJ�˛g�t�ڃ�� ę��3�=�3@c�9i*�iTWU�t�⳧��;��:l=X_�Q&�~Co�mq�����a����x��GH�ӈ�4Ѯ����J���D���G�$w!���	��QQƽn6��'����e�H �1�12�A#�$)�aJ��)�jǢ�݁�y�ng�8uJ=�{�a�n3�y�q�n�<��3 4^3�6��@V(D+��1�B�f��]����o�l*����[&T��*L� �g^���-���w�v��{�r�ut�|W���z����Z�gp5�T
e��r�e�lw�w,�J����O��]����덴��P�9h��~�«\����.�-YZT_]�$���蕜�u�t��K�r��P8�(Fp�!L�(dZ�v��>����!txYDU��)~l�L�ڦ!��̀��u���ylq���xvs�Ҹ{�R��s�_����]/Du��b�i����?�3V�SG\
?3�{׷Pա�W��kj��8|���U������{^��±��Jmo=�Ք�ӕ��+�E �񁷯��U;K%_�B6򎚇*{ت~��g�"�ˉם��|l�Ѝq�ya�C������b�#!"�7{i��:}�����ڇ>P���Q�ė8���a�v|gs�A6j�k�>�K��d�ãj�E^l;��l���2m���x͔��l��w�DO&�.����_W������:) f>M��7$] x����;}ʊ��z=�����*}����ީ��_/���Br�.f��</�s303z��<<�.���Ŭ3GN$���
���̳BGo4��R_����BΑ�+!EB�I����,������C�=)��ˁcW s,���Ҭ�"ϔ!�t쉩�lx�T�;�i�Ѯ���W�!OVמ��LT]TE��!�lZy�����!�a@ᴟ���.s���c��]���{]8@\��l�f���-zu��"��^����{�a�ԅza��/q�-���52X�-�z��5Hy�$�k��=�c&6b�5�Dj��g6��w��YG΍23YU�p8pb���Z���ÈZ��l5�������m�n}շ������Xje�:�N~I$��]��'�z�>�y�v��m���ͻ���`iΚݞ�6v7��P0����7V@�Vj�t�]�g�,��ǈ����D!����4���}.����6|e���QR�����g��������F�����?(�YNgl�s(6��f�J��y��]2x�>}�^��ty'YJqv�l���)�!�D)��!AG�o��a��z#a�1R�5���;}���=��A�Y�&�t�^� ���F�`�ց2���7�P��p\݀
Ȭ�IyoOk��Q��nV��+Ɏ9ԩ;sy�O�g>�D5��H͚2�(?�&�c�7.�qI}�y����H���������1����z����bYx��{�������v�,�F�v�5,�����q�Ei����Ù�G1���#�^��2�kE5դ�U��$�.н��_^l�)���#���u��(����./�yJ��|t�30�8�"���'�k�v���{p�B��5^�l�9��U�[�k����E«�f��׳����l���u���_ZYz�jN�Z��RvH����U{ʦ1��-��޸�A���դ) K����oV��1H�Y�"�smrH����}�����?���NG�N�k�־ᜇ#Ƃ0�9݉�u9ʝ;�hL]K5�˄l=f����i9;�.�z�SP��p�����]�"�lm�T����n3T�ފ�#h�9u�%�	EO�[f��!VR:o�3�^�=Ɔկd��9�7z�q�͈y,���xE�2霭�h5��i{�����l�7��u��<��]U ����<�3W�9,m��8�x��T˞�Sp��L4-XȚڴ�~9����A��a23}��.3k�&�U���Wc����C���%�K�h-6k��?�^�ы�,�˱vښ��\�1FV��ڲ�k5���o5���~k�5^�l�b�9u����@�9 �ΥԱ�<���V�u\maU��p��wW�އ@)�~�g�&P�t�~T�����	����n�n�Wj9��$,yr.��B\@l�[gL�>u��\�<H�(�����F�۳}t6�ƛս�����ck�h���k;������w�lV�<�i�n�e��ǚY���W�):�2�a�XM��/�� n��{Z\�# ʷ�ܰ5#6��@�����`�=M��-�=߶��y�B�!O
��A}�8�̠�V{M�죃M�L����u��B/@�z���gif���`{�U��m֛8B<O#7x?xO�q��6��ް�Z�xF��<�w]%�y���o�tp�y�ﵮk(]������V:D��o��Q��{q�{q�ik��"�\��&�ox�#���:�H�e;�&�J{!�tz%�<_=�A���n��as���>� ®-�Gt8�%��r휓t�����y7�MGw/��o��z��܎�4���|z&��$�O��O��[���p�Ш��I���G���yQ��ޜ���̬t��S=au��*u{(��(^�[#m�弯(��l'�'dv9� �g���%�x���A!�|�ٮ�xG��z�꪿]��V(6=���t�+�E����ĳ����g����bE�ñ��J����S����,V@��jr�� ,�)���D:�ʣo�]�Z�7��}j�!�t��{��(�e���#��	E�<�i�����k�,�4*)�:kl��/���9qD�����A��ol3�u=I@�<gx-�2��[��08�4ѓ�m�����8�ˎuS-��5C�Ua]�<k�C���a���\���)QM�,��1Y1�7][�U�ʷ���rV�H����gP[^�W��
Լ���S�nT��y9�ݩ�N�	����v�tpC�u������H����s�.�*�<:�;�,=�����.�F���Aۭr(��_*���Z�4�I�Wr��1/������d#!ǛV�d�T���vX}%p{R���zwh'@�Mќ�:���F��1�{v�f�7D��g�:� 8c���j#��s��Ү#�U�����{a���&�Yaܭw�t�ة�d�λ6��vo�nM������}��W+�ќb��c���"��r��#Xssi�AWVy=Y]28����oZ�� []v�J�@΋vj�t8s���i`��ꫥ�jiN���.�"�	6�+\�X����:�Ee�0�U܏؂r�H�;����{��͊�"�E�?T4cŗ�������{�.І<a+8������]gX����E{qX��V1��J+�:�I$��6��}d�EYh()����;�³1Ji�(��n��P�QQS,�J(�ܻU��;+j$�yO�;���ƚ.m)gJ�a�Sal�\p��ڵ����[ ��9i�6.�6h��&�p+N,�o��$ݭݥ]����u*ݏ3����B53�5����ᚂf��ʱ�`<�t��#2N�#8�+D62pP���f�yʺ`އ}���x�َk��T�Yt���eE.���J�������
��ea��t�=��~.�[c��Y\���LФ���<���� 6�X�E\�1[C��8{s�g�G;^��	����OV�D7�'R�]ugΩ���pB_
2>���[4��aKY �	��p�C
R��$b�3
9��P�.����ҫ*��;
��Efn�g���k��z���O�1��Y����b�,�n&$}�I+YT�ʐ�B���%ek	�%b�1kt0+S�S2���hf[j#�2�HbbEl�V)k+S2�j�C�i10�Z�Z��U"�7��[�cSˮ/�K�c�GD���V���9/`�����eo�y���W1>�N�4C�]zZ����n�hgC���h��^P�Ao��r>wgB<�w�.�5��L���oE��:����_{"oI�8}��$A��Ϝ��x��;��Mu`r��oG����Y'�G�4g����@Z(�ynJNZ��QB'lH$����n4>|w+r?1�pD�
��.J�HQd��;<=�3)Si�����,9�xKϺ�cnα~I>��Y҅�D�R��ׄ�%��9a������=RU���.u�!��9(��1�ғ��"u�������O��6�$9:�\�B��4[i[�3���/��z����ڌ槟w��l+�N��ԴA�g��v���Ԛ}t�;��X}E[L�2:�rA����uŞ��E�hVnF�S�����b�vo m����C�1�4v�3sV)����U�VFyR�_5�����SGo�9�P�LyW�uJ��|�zkK{sx�jבX�WO`CN�����̽�K�t.�T7�U�7���C�_�z�T	k��s�e�jZ����EA�G%I{��Z�a�&w�;�_Q�!�j��*$麸���H�P��4z��W jwu_y͗#
�<M`O�_�-�N��Y���m=]/8��4�eq�h)��R�V��N��<���*�^,m���U�Qr�5n�"�y�nx�_Xny�����SfҊY=u���
�l��/ǽ3B��%�LۅNA��m��E���i�+�n��U���]cKs&��^�Hx�����g�4i�Z+u֋�G�E?S���srv���@���gA�z�9c'g��͒K����B�?p�2��Z����R��Qy�5�h���g�״���5�����d��SV��8�W���65��+������8�Y1�D�XN��z��=S�bh�ҽ��~�NZ��s�G�'��v	 Ɗ�D6{�}F��+tq�E��Ӑe���X���s4���55��[y=o�����Y��@ג��H��3�O��>g��I]���m�EK��7l"^�
�#6��X�BK�F���;v�]��l7F�yqwZ��RZK���GZ�]ޭ��ދ�R��N,�{�M��&�Ӻ�Aw�qUt5z�Ilf�0��E��뢫)<���]��8�r�|���DP�^����{_hV��t�f���1��Y1�jH;L�ǵ���Dٿs4/���5i<+��!�{q�����&�l+�{qW����7�M�c��wٜg�k�]-��2��ܭÅ"���]���E��U+�b�-�_z|{ݐ�1��pe�V1A�5�Q��i23[�|��i����d}�c��,�oL��Ȫ�έ{�Y��*�S�ܺ�A��h`Qj@vr��ʕ�v߷����=�l�!�"rm%^(tMLᭃ.��=���V��[)ޕD�<�܏ɠ�D�w��hy��zd��f
+�NTZT"�͙�5�eD�u:�s{�œQ�`�A�[g]�ۚ��a_٧�� 7���x�7�ZU�\NΏw{�+���d�8��y���3�����Vp�p?q%n�������>9[Cʔ4�}wW@�@�˺ ��s���g�kr��X1X�c-��**�h�ժeћ&����qU�}���K+�N]�Z�RZ�H{�@�j|�k���3��4/k97�Q<j���=dCY�4����.x�'kR�كW�����]O��z��=�Lz낺G�G�~�ɭ6��ܙ�x��&ž�M�7qVW*��;f7V�֤�on�Q�ְ?Cb�v�v1������@������j3��3���_A��uG�m��a��i!kyP�a�8��9x�q��g��+�P:�����/�z�ْ�]��:R�ȋ�����ecʾӎj�%C|d2���u�`���誒�sc-Ńx��+�yѤ|S#�7�Q���o_%�O �t֦��7��eh�˟��ݚ�y�����������D�U��C�y�ǈF���v���m4���m��5�.�ÈZ�'��{�$����kM�ި��LV����y�L�<��͂���-����J֪�����C�����m�����CeSY�R�\Ue;L>���ǎQv��θ6���|�����K��I�y�{P���˶�^#q���lo��r��i|`e9D�������ʉ�"��ī�ײpJѢ�s>l�OwL�i5׌q,�t�˯ f��]e���\(��vUt<7�1�U�h�Sп6�8�A!��mD�uܫO6�'b�Z��Q�G����Y�.��F���	i���<�ｮ��>���I��Txo
ڡ���Ub9�NS|�eNծbwQ�^Ԫu�؜>���g�N�����WO��� �����gP~ځjzn4l���`����]g���9��T�]���]�R�}�&]f���;�ocyN�2�U��nM)��]�%1�N�YZc�K��I�KRM�Ыz2�4<���\(�ݲ�+q{-T�41^fbe2k[u|Z^f�N{T�n?7�>d��Ga)��v�x�z���bxu:�I�7���.�;�gۂ&9m�d��V�㏜�xW<�+�jbp�>�u#N�eE�b�?_�
�'7}�hni�5�<�-;W=��WFH3�oY�)�*�B�l˧�evʺ:�C��yR�[A�\C��*RWX�1R�:�]2�����]����-{ܑ�c����Dj�j�a�PԔt�8u�'K&��#��k[)vZͭ�����5r���|�B���+V�111��H��լVE&�f���t��XMyqd�7{�tb��Z�Z�Ri��PP�8��#]��-�B
��h���%On�a��!�.��4vD�����`q�k��\�-{7#�����a'������=��M��Xs��F֫�:�Uu7�6n�v�F#��jkM�� N��\��V����۱[��r���=JJ�[X,t���E��L�(d�r��SX�|�j�H2�d�9vn�ϒ�YkΥ8�M��n�t,Q��Խ�{b&�\���%FD��z�
뫻�R�KF�4M4�_�nu2�0ي��Ot!��ѽ}���\�U6㛔jT9}D彍�\m�Q��Iu
�ɞ*�j�=�Z�n�Z�9�WG]c)�G kI�'N��{I��z�Os��c���G7s�+v��y]�*Z��u�1d��R-c,�u�3�:S5X� �V�c�j\�^-�%-�{��� Z������B�umC�(�Ι{��KH�g���5�e��ܵ+Je0�)ӭ���5��zn� ��X�
=A�tԨ�\���W)YVE\m�C{�,+������q~d���b�ң��`�0����)�ۢ	@@gD��S�5�z�e��Y��ɽc6G��&n�kB�5��7k��N�!���Ҳ��.#��eSUs.eR���WIMX�*]5�fU�m��0Ȫ���Q1Ӥ��UT���e�+uf�X,nZ��(�lZ��b��f\�A�����nf�iӃ1��V�-,���a�L�3.:u������D��T+�2�+LL2��Q[\����:����ɓ�\ŶkT�a�5��VR�PkA9>��� ��^ޭʛ�g�x�ssq�ء��n1-�/
��f�ַ0]Ճ�Pk'PR9��4�'�^+�ٿ�!|txWN��G�.�R1��Q&��ɡZeq�r{�FK��緑9���t����~%-I��kQ��r�g�E�m�v��I���ن��{�?C�����G\�,�Ns�:��ؽ�Q�}
�X��M�ܣ�[#9��ua]j�>�7�Gz{�Ǟs]�Mw�z�7GdN����p�P�%�Q��!�5�(�==l�G�G�=ΧU���sy�MȺ!q�,�����j�mNI��ՏX7������w����ـaޜ�,�#���TU���p8Q���	��h�lN�<�E�i�W����7(�r��Uج��]��P��6�'�*ڶ6��J�u��n֗^P�S�N����S��'$��E�=c����짶�s�X[�w�Գr8'�E�z7oonT���k�qt�r���BV������8X�O+����<�r��t2k��>:���}{
u�����0ٲ���p}�Bw���no��A��ꁰ�M��V�����*̖_�"�Xs����WN�ɝ��
̱pڜ�`�,~�b�L��W9B���I+�ȑ��"��#�.���լ��-=*SzH�a��<��98s�h�I��[^5�p?��	��M�M�u6z�T��x�""�U���} �RCjڣ�<�`3����L�#��NZ�8�����d�!߳�H�9i�:#^���^D�1��x^ҧ�g��YTS�h88�{er����T���3f����q�o�����{ب?��Z��7�nX,� �~CvwW4�f:y�[D������|�wq��떈w^t죆�.j�ڑK���Ĝ��1���ړk�lj�k��v��T9-��w�B�@�Sd߮u�^����u�=cdre>��|�5��"�h��_�|������<��x�{vvf���ئ,c�/�Fk"�2�4��`b��ڹ��U#`s�(�5�h���>��r)،S���9���%ۧ��w�v�"�K��΢	�ڜj�D �ˤ{�uj\Hۥ��L�!y�Y�դA*��E_�3Zb��t:�]�S0`�%t�?��aybޮxB9�PǌR�s�-���Q��Ҭ�cH���	W+y�X2��$��qi1+�i��cQYЍ�7���F:g-)�M���,��'�Y�k�^�I�7!W�S�"žs�{5�x��qq������3AÅ}g���D�&3���b��׺�Y��<��F����鍉�L���<l�hZ>�Mv3NT�;�/��4�|��cFy��dR���u���.�k\o�(���`ÂqĲ�$�Ls~Zj�<�׆��{̦��T񺼘\��]d��L���0�Z�sh�.��FfD�LK5���V	�-�B�W���3�Y%���R
�ԔH,�ޑ��^5�g����&<IUf�8��/r���3��]e}��}%��b���"�K��j�B�A��Gh2]�͚��sk����oz��6�l��)�[��t��^���g�c�z\�ή,�T	f�}3&6��v��H��o�C���N��ڲP�&2wW{|$,�4t����F��OI���rFwVr�|��t1�v�W�)���NI�(�2�hqd`�ؖ��6��-���|2�rH��S-�Uof��n���#�iv"r�]p��$��xi�qmw��P.,�@�}�|};1+���z��,�Z�>�G4�?]�%�35���Nh���^eoo�i��#���8����k]o7m�]^޲/����s(v�	�+6c���L"w�<�;���&R�y�^_���`y^r��8�_`�j��T�oc�c�7'*������HSTs����->V~[ĺsmsi�f5�I�Q7�N�A�/�s�����B߳��J�Y&�-M�=>���cZz��?���I��qp�/���+Xq�)/����3"}��&��_�I����E����+���Q/���z�%�zፎxA'S��jD;n�E���Qk���w��9�F�eϔl��]��F5��G����C]cꋶf���L��<���	��$^���3�8�<��y�
�ZH�w1F��w�wr�[��{������'���7;�/��x���:��/Zh{[�ukzUV�{Kx����%���a��y�aLL�l�חㅑ3^U���b.cWC�A�m�`�	{�L���N1��u���L�\��� 09/
�ħ,n����cB�p�`ڬy������l�~]��H�����?\h���=�t��Kr���+ԉ�t��]��A�Ͻ�:�O�Id�+��ʈ��z��<�yί���x�*p{�s���])�F0t��\p%��V�T_A�аD��S�2�W!죍�b�f�N{f,��k�VL�ސw�����#� ��Y��v(3��鉍;�7g����s���F}�>d��F�R݉w�lZ�U����v`�N���M���5������S�-t]	�˔��L#�r�q��E���y�y��A�ޯpz펒�.�.�ܽ6�ٽ�xG�i��$s2��ޑ�\�{�=B`N���WH��u9�\�Dtmi�e����y�&/��h�����9J&+�5��=�Ƹ>��{��{qB��Yغm{c�=�����nzz�^�,N�O���'ip�jtWx�&�����R���-��[�TttO��/ޞ�!Q��ZN���VW�'c����_����s�������g��r���c�B��^�"��"E-�uh�R������pn�*XJV��E%�y���CجG�eq�����0�v6Q��u��b�qۇ��@�W@*�D+6����wX�ᮉ(�g>@cB�%4i; �F�N��R
t��5����ʸ�2�ĊfH��GK�]�j"��L{W� ;$ƖWZ��z���j^�R�2S�p�y�*�H�*[Q��ڬ��˯�Y���=��B��]��J��#Y����K���3$qt%;��n�@�\�v]Ҡ��x��TkF��y�'�'���Ŗ#/V�Ι�@F�*�M}nB�W�T��v��ep����|t�O��]�����qgpܙ6�� 4Un�]������r��7���9�����T�Ee���@B�faz�k-.�}������Ӎp���本�v�nƸja�J�F�.(:�IWll��:��n_,�R��.CB8��6j���U9+V�N�#�d:��fв7��t.2��u�Hr�9uU�L�ڄ�\�Z�YEtX�����B�s<p즋p�����e���Y�vvʴ-w,������&��Xa�f��*P��
�[U��J���G�M+
�QT�*�.��uy*J|hl��֖�FCv*��ݐ,r�+��R�m��uR�(�6���z�ƥ(�n��AzbeYv�L�컣�m�݁�;���{�0�2��GU�{��A�}��}�|nyƻ[�\qTKu3ce���n�d�T�J����YJ�ܥ��K�6�YSj�-��SY�Դ�̴Tn8W2ۅL5��m���ƪ��Ls,B�%�f9��ե��[I��E�V-U�3*�lk�9�.Z�k\f%..J%�,�31pF֔�F�k)��\
)i��2��-nfYR�Z�,�F���G2����.�]7-.�J6�T�ID��]�[�x��Z�o�7���2�
���q#+d�|9(��ކi?�%%=�`Fm��pu�E����� �$#�P�qs�N�B����ͫe���E�Z����i��6���qsͅ���U�.艹L(�ATK��uT�}�%�8yv�hU%m��+ݫi�s��w�CV;��ݞ;�b����ʭ���(U�6=�>�v�@��$����u�G��Ye�tU�_W����g��n�{�M-��tQz��QX"(�!���0o'��ԭ�wQZ	e[C=I݇�f�RZ���O!}"bh�33�kFH���R���#ف��r0���a��- �h���<y(�>�#���eSVw��,� �����Q��V��A��?Z<�1��{�Eہ�G�oU������YǽM&�.�����U�CJ��L�<�#j�Ӑr�\��\{�I��������K�3&QY����Aj�)�:�!@w1Jj�R���+U弮�o�ޜ���hG���ݎ%�N 4[ڇuVƙ��JX�
;T_8��p�3��_L[����܇%��J�l��E�;�*x�f���H?S��pBQ˰-������]��.�&l���:�7u�Iu��n_|�씚�Z�ε��J$�Ȩt}G�8>�ׂ
1�^׼��gi�c89�ś~��{k�U�@^܋0y��qTy��+}9���b&1
I�gi��)B���M�o�dOj�(��uĴ\ʰt��N��.W1�#HS���=���x��4Bz�̝�����&�T�U���z*�4	:�,�p�p�vBXQ�,���]1����ĝq8y�@�KU�oV"bO<D��OE聹G��'j�fS�R����I��O�9b�y��� �+��R�!�3���л����햞��Z;m��IC%vν5�p���y�l�0��P�z{-��S��Ɗ��/�5�*9���9oEL���@H_��/����S�t����m�MiFl��5y���V{fҘ��:6w�5����^��a��{�o�1���^3�#|�=0Q�g��\�j�b���W�Vs�^��y����QlC8������j�z'1ɼ2'VW'şG�3)��a�M��M-&u��L�'�i�7<���r�A^�m�+١�]^�G��n�Ͷ+t�i��K���B���C��w61]7b�xa�}[��d�)D��)�Z'��\p��_T@!�PJ�=v�W�uPЌ��_5�����޹杈�fC	���j��=�X<���*����J
��)�U��Ȗ�����E�R���NP�&2��z6,�����5��}�0�1�$�i�W"��Eb5�^�<��}l�0#��v'�ʂ����Z郵wR�
���aDе0��n�r6eA� ��Euc���-v����V�V���Ǎ��\�nuym�t�!U����$���N��Y�{���mk[	s{+cQ�X�7�"V�	��1 �(ބ�U��⍌��a��&I�+'z�&�7��wq��~����y���'ȡ�3hwU�-��N�z�Ŷ�6�=���B�f�����Fi��$�f��B������T�y�wE-��_=�H��X�����X�"p�N�bl�\^�"���0GF��m��5|���F&�j��!�E`]����� *Ŵ�\~���Iӫ��y���)fl�)�0�\�t\n5m�����NI�Y
�f��I���K[Z����wP����e�8lH��[$�n�6�Q\ne�4{O)Ź{����S)�[�
>�»ڮ��_yd�b���]z�8x��+���{P�����׷�_h���R ��Z�f�� S:ϞM��8�Xγ��^�����^Fj4n^�xԎ�5��v��Ӈ<��&���^ޚ�#���b��k[��NӚ:�+�^�U��f�M(�д�S�e�7���u3څ@�ZkM��T]u�7�cH�6q0څGt��W�ąoJ'�'�����@�(o[�Ժ�� [�{ ߋZb�JҬ.ڽW+�xԣ����p�j���|}�<�`�m<^�yg�R�&8����v����lRZ�C�IN��S�f8��W�	�5F���T���Ƕ���3������IsJp�ዹ7��Ģb�c�O`j�dX�6�i�"u��q�;�+]������Q��OqSr�ϼ��a
{�[�v�ɉ�&t�5�!�'4����]�N��VU�ԌB��c7�������eطAk�p��ކ-S9v2wp�'�:�������{C�}��Ǌ�����y����V���6#�iJ�2�����
ʉ�څb�U�n2y��E��O��\0Q�)V�܃H���C%E��uóS�۴�K�Ň�@V�x���F�f�wy7��uR��W��e\�T`k��lM��t��{0����O%qy��}�����F��7�An������J�;���r~��|,~�%!��[:m
ހD2��^a7��O�v�d��<��W������-�}y�(=���Ho������/�*վ/��▹��ǉ�]�����@�{����M��BK#���Ld��l��mK���WaV�D���.6�T��3tnl�o�2&2�#��5k��E�tS�Pf�B�
�ޝ��j"x�s:v۔V'�eV��G �YN]��nV�J=�m��]����1��1SӺ�1ϟ�^���c;G��y������ϔ`�f�q�^��S��uc��ۘTѺ�w�����$�[E7��Nx@�^mc$iTVLނ�>�͂�xO������z��8_G��S�+o˕�G=��Ь�[�E�ͮ~5�SGy�@��7X+a��w����bg|�5�a����~��e��{����Ԛˋޞ��������a���S�iZ��_م�I1��� ��{��d� ��n2�}�E*fzE�,^��_KoeFU��GO��:�עz'�	$P� �$${H� �DA(�o|*U��4���׋Egb��%4�[}��6E��Y�WHb1�ۭ|�zA$�RUp�(�+����g�=���̹���}�R��Ɇ��^u��䱫$h~�t��f^_r�K,�͛����r�
���Li24�$"$��~o�����o���h�"$��Rh���hu�UE���:�����g���̞�}����s_�^;_�t�;N�%Y��DI5>�>6���;Ԕ�ؑsC�Iw=t�H�\�g�WQ��"�#��E��YE��rJ1��Ҏ�Ƣ�+���2��/U���ZA$��8Zm�����l����ׂ&�!$�?U�d�p*�7�-.��z͵\�����2G&p�?�&��A$�&r3T����l�r&9���N/'̌E�J��<-6&'ʣ��#��}0����t}�g����Z{��;8w�K$"$��KISj��zH��ޏ��!��vl�?�8����cB>]�{;z3��;�V��'�w�u�}�N�?3���:�("$�Gj��������=ǽ�	�S�ԧ�,6�N�QeKZF\$I(��\�"I��r}�SaX}�O���9�2�����$�Ц�E�Df�y	$��u^�UE�E���d�}�	U�A"Ih�0��M$su�Ɂ���ܫl*3��Ԗ<��nd�^I�r��
K�Z��4�&��W�\����&�s��x���:�v ��VEz<��J9O!ꔟg�ޟ����z?$�9��S�.H��9ɽ���'��]\���n;�ޕ�"_�:�e�s��_��YD���r�S�r	U�E��/�b��"$���?��~��a��n?���8�|�%����j4�j�H*^)��fJ���wX�pPǟ�:ylo�3GITy�ʭ�6��ciɎx3A$�oj:ќe�u��\�n���On���l8r'�Q�Qe�i۝���2���0��:��""I�IROIy�.<��e;+�yz9M��!N�;	�)3L��q��d��%fY&���/�=����R�Q�O�d����7r�O�.�p�!ˑ0