BZh91AY&SY^���׼_�`q����� ����bF~�      �����25K��m�A���k��[m�����h�mb-m���֦���m�j������%���Qm5����m�:����wӗ�T�-�Z���6����KJ��%6�i�$����mU��Z�f,mjSJ&�1�VƦ�A]�قڋU� Y�Uj-���6A�w| ��|35݀��f��,�ғLV�X�[kJ��l�ͪk6�[Z�Z��2�4�$kUT�Ғ��fآh���X�m�F�&��[KJP�d�V�Αj��ed� �  �fo��Uv;�ۣ�n��sj�d��s�:wn%;��n�vN���t�USV���6�R��6�r]jKwl]ҵ[r��W�$45���[F4mAx   0��M4ϯ\h�N�.{ٽ�Ҁ���[�z���=�᧭k����	P�3�Q�B�S�z��zp�y�A�m��Ww�΀O�}}���M��V���l�M�N    w;;{���݀i��}�Ҁ��:����y|�
u��΁��=q����>����{� >�����}zt������ �M��>�w��@���۾]|����>�X{�+P�f�Wю�m�2��   }��>R�����/�k�)R��|��o��
�>�>�(�����E@=�}���2WЏ��=w�� �M9לw�����������-2��[,I5V�iO�  f��� �؛�"�	��^�ۣ֫9���aGo�� �m�Ү�w�/G��h�<v�%����F禨+R-�k{��5��;o���*Em�ϻr��i��a�[]� ���B�$�=�:�5��v�� :�=��AB���t��ڴ���Jt)��W�T����V���U�r�M��;�y�@��׽_VH������k5���[3[x �����=��EZ�ׇ��5J6������� =�F�<�:�{�n  ,S +U���Ӡ�;8@�n*�r�d���Yl*�Y��Y7� ���Ҟ�%�Ew8\=t �:���n�n��� t�Q�@ Όz ���p��� =ǦūM�Y��V�m[2��  v��� ��� �y�*�ݫ�� -�8���^�T��yM^� ��\�@罳��ho^��2��[Si��(��M|  x��>� �{tN�����` z;#  -Qm ({u=� 	ݩ��4mU��Tt�     
   LMRT�   � 4)�IJT�F M41#�2`O��JT� 	�  4Ɉ��%*J� �   �d�O#@UQ��     	I!�TDh�2e0���Q���z���7�������Y�'�~P���gf�ea̯	{�9��������Ͽ� U�^y� _J �*~(���|?���
 ���$~����C������}�?��*��-UWQ� ����0t$�!I�H� ����_��zG�X����G��/�`��,��Xd?&� ��:d��XS���D�"u����XS����*u�:ʝaN��YS�)7Y��)�D�u�:ʝaN�'�(u�:�`�X�	��(u�:ʝaN���� ���/X���� ��z�=`��Q�!0�X�(��z�=e�/XG��� u�s"��z��e��Y��T�}2u�z�<`��XG�#��*u�z�=g�:�=`2�X���T�*u�zʝe~X��YS��*u�:aN��XG�)�S��
u�z0�XS����*u�z�?�Q� ��z�>�S���*u�:�=e�d��XS���Q��=eL�Y���A�?�Q�*u�z�=a�� ��3X������z�=`���L�eN�Y��A� ��z�=aN��`f� ��:��aN�'YS�#����
f�
u�:`��Y���_�@�"u�8��eN�'Y����u���(u�:0'X��T�
u�==pYG�#�T�*|0Y�#���X���E�*��z�=`_�A�ʽd�/YG�#��(��z��g���s ��z��`^��X �'�
u�z�=c��0/�Q���zȜ`:��d^�/X����*�0�Y�z��Y@�*=` �Q�Q�Q�@:�����(��E��X� 	�Q� /X��=`@z����e@z� ���"��Q�Ez�(�����D���YP�:ʢ��Q�
��AOP:Ƚ`�X�#�E�`C���A��S��E���z�=a�/���z�9����A���z�=d��Y���zØ���S8*����zmTU(�2��]/H��d��0�3fͱ�K�M�FS��Ҏ`-��X� �;̻/L�jx�	Gu,���,�CR��M�׀��j]�T�@!�vY`�Y��^Z���{���[�2Xt�#����)�W)e$+���V��e��Hbɺ��Cc%T���`��ݹ  ��fS*I�vL��Զ�D��;�{{�e���p����ȸV��Z����U����-hP�[)H��јM^!zL�d��+s%��[/v�9�.����6�]xj��CZi��BP�Z.�^JRR�B�#hr^��R�(��ZA�L�Yt`	)��:�Uc�1H����K�OC�y�n�`�e���&Z�U
	���Q2�ٗOsS�znf0���ī-[N�Ҩ3w�غ�1<	�B���f��P�/fZ���]ՓאmHBR���c�e����Mb��A%2w2	�F�U��A���REǂ��9��4,�s���on�v]�0A$*�%��Vk\0CԉmD���Ra��ͫ�1zU�J��˭v�^|��I��w�j��^�7.��6�"hä�r�����۩�nH,[�qj6�:̘�l�1�^a��5CHm�
d;�A�A��ZtMǣ,��ֵ�F����(S��4����6K��)W�a�bU�ZHȕ�x�6�Ͷ^o�4&q"9���b�oHǸ\a�N#ib(Vd��L��4�W����-�e(o$�ৱ���m��l`���UcnI�& �IdNY��l0�mϥ���Gr�6]i��*剘1�8Đ�����Y.6v҆҄���L7l勬a�̈&X��#���^�v2R�q�Ct�uۆc0Qݴm���&��ܗ���Sh�L�-��E'�L��V7{h3J�a�[�f[�YV��w�#��� ���i���~GU�����s�[ye�p}�f�X2�!1
�j8kV@�S�ah�0�L�dQw����˚��֛p��Z��-6(a�"�3ܑ;�V�3�D�͊��]Ev����*b�UY�t����wFT��5�#oqD��;4�WW�sZ�4=k	;�B&h�b�'%
ʽ���KCM[�mHf >����d���"2i�K�/ �C&R��D2'�$�-��V��*���y�[�ְ���]��q��K9L�ۢ����Xt}�)иD���#L]��f]0�	�� ���B&�{
[�Y�Q��f3�0�F!w>ߚB�[�M��T���0Ef7*�Ǳ�R��Ff������H�a{{�5�v^��1�4)�B�ј�AK�b<��&�f�Y/,�e!Vjm!��5�f=�sEcd�4���匲�{a�kM�A�&���aڼ �m��`[���$�ܕ����KP���J�`:5�.���\���ay,f�a[{{z��cf[E�Xt1��M�6��L�p0�6űA�9-|T+��鿌{I��՗d���k�5���Gr�r�J�KH�Q��4%d������I�0"��B�ڂn%x�#[xX6/
���ӹu`g�P{I�]�+\p|�$3Cq��%:�b�����O�˸�ܧ��au�0]�ҽ&]1�c͌�B�:M\.P�P��^Mq�#/%+&�ԙG ͤ+iI����5�2��ԃW�c�ཐ]6]�tCy�
�/�,�d��ج�	�UԢ[[R��]�.ʭ��/��:�#�+@�ⴧb�{�$�A2�g�N��e6��$;��eC��P7����l��Z:�q�2��rX�c+0��ˎi�To~�S*�2�8���֘U�=��唾.�;yJ���j4�SUkw�SS*]�Oˉ��V�^�j��!�l� -r��Cw��u�H*��>�;���u�����Ͳ&if3v]a��,�`�6��0�(PfT�*���i�r|���oj�C�u���Zek�x�7U���4ĒM��HwUN��Y��X���Qõ�$� �&|�,a����
�&��2�;�t\� uu�(�sSl]�pGe^�;�<�oS�J�� ҏ��q�n�,�65S��ڳO�uga��tr��ґ��-;��m]&+d�h,�ujnkupt8u���P���fDY5�ND&��(f曖�Q�[*cn�;��i����]�Vm�Y(�+@�e��c�[��i�E�/*����w[.�.�ͺ�����I֋ь��iiLj�+(��d���B���+ڼ�L�u��
�2P*�b����ê`��+7������%&-�X��WK!a���
"���V�`��s���L��٤\d���9�Jͤ5f]���#\3s�Cs*�a|�4��wl��PE>mҬO:�J�W��yt�]�j�Wst��N�t�1�0SvR��Ԟ�M���O ��.���AQ��$�T��U�4��x>��d,�JkM�ӛkJ+,����[�����t>՘�Kl[�K4���íd��/���,��.��)����2�@�[�%�sw m$�`F�5iՕ�ڔ�%I�6�ٲ��Y�V����SrFr��w��1.����%+r�M���1�Q���Z3F�%YH�m�z�Y[Z�J���Ch�l��1�A2�����ݴ
Yv���m�fV��m�n���Xn:����*��NTO2tXֆ-����U�Z��ޠ����]��JÂ�E*w%��F��Y�Dݶ�[р����@�RFT��ǣc�yM&Z@�N��d�M����W����l1�)!���*Y���牊jR�$�`h:�YC7t�] ��l�;Gg������N����j���7��	9K(e��6��(n��g2����N�*�J��W�[�D ��S�)�[�������Uš�z�W����@P�F\�/#ZZ�7+5\d!�n��RX����f&c10�Tr��l�zSC]�b�+ج�tr�+�ک�C�U��	���L�S ���K9ݬ�`Y��
l9�V�����˼�!�­Q��H�)&YǃгM×N8�ۛ) U���V��ڽt���a�ܩ�5CJ�)|�ź9��S��i� �B�Wu-��]6��;�Q/6QEQ��[>��f��7��"ֺ��{%:�F���Od�$v�%O4hĵk���L������3��:���ێ���Zq�cF��L��%!���]������E[��	b�-d�͕��Y˕[����b]�[��dȒ{f��B#ol�W/ JjH-��]ǘ�-c�I-�j�AOvL�!*,��]�E��
��p��7[�[OtY*�`�iVP2�E@9k%Ã0��fK��I�ȳw�X��'b�-�>��]X��ad�q't�fT喁I��O�2Ɩs-�r��5�G.p9�B1�L�9���uuz`��٪U�-����(PZe�V�\Z�&�my���"u̺p0D���ѭ�
�5�7���Y����T�P�3.b`�4�IE��G����i�	)��m�y�5�*m�WݳT�a�PT��G�̤�5.-ۦ	�+u��Be)�R��Ր�(,��.X�S6ª*xb�L4v�e�il�K.����N�8�ẚ"�wr��H���Yj�lkz� E4��]��l'�ı�X��K�v7w*!�8ʈ<P!o4�2��#��`�5&rTD����h`�����6�)V!C4TP��![z^�g�e�c�YV�r����"�,� FÖ�@Kh�&�K)�uy���)�Ww�T�M�h����O�10��LhR֞�}�����A�;�3B�t �
�1?�3
yQ+w�.�jmـ��F�)iSi7����E2n�m��n�u���7�Y�ohm� �T�e����rd�>9V�Q�0)Q�켲�:����N����(��S�m,b�S�n��@��D�8%eM�$��+^^'@b6�o^f�XcHs��)���&`[����1�zC�.�I� p�[X2W�/.AZ1m:eI�d�媻$`ٺm�1�;��ݨ�Zi֮;�vr`TP[bV�a;��ђ�T�I��7�&��/~A^�GV��l\���n�Ʋ��v�\�V��.P9.�ũiLH6]eq��1^q�)Jr�9o.X�M
/$(��[�O]^���tb�O �n��GQK��t؎�
�(�%Q4���<8Q���Z�/�.cfm<���2��k^Y&6���`dh���[�ЖC+�5cj�0�`F7H�F���ӻCX�9nX�gv��ڌ�GEVJ$n�tF ؑX�)���o�U�Rf��d��ƭRw-��������H�ARR�ul�-yO �@X�L��KE0J��Δ�*US7q,l��9S�)j�b��Xe�54�@�Ӭ43���h����:"-�yZr٦�z��w�+�R��5��a�)�(�
a"���(�#��n��t3ch+(�����n:�ٰ%��nX��r��fڈk�����F�oKwy�McԲb&��f�쎑�2I�;�ü�y�cf]՝�P��X휢T�?=�n��rW�/�V����o�lU�fR��5�Z�v�U��H�Mc��Pk��Kӣ�-�)�,-�t�U8�����Ub�+2������u�lq�@S��W �J�����S�L�+���	HP1Ei`���4+6�T�����WV�L�]xMֶj(��8�*�4�yuv�L�)VUJ�j�̅SH�驊�F!HܘV���ۧ�L+.�MX�¤��oI��0m5o6Zi$�^0�cɵ��v�*`,"����@7��o-)֥(�j�6�ff��:_�5���G $6��0���� �ne�z��Yt�P�A�gm'Nj��SDo���;pe^�
��Q�ڼ��pn��N��.(�%6N�S[�p(okQaS2���:)T����H^�M��+]�]L�S'�d��%��[*�M��E$]��@�m�&�җNbڊK�0� �y�5xꚦݧW B��ysSREU���XT��������ۅ�yElw���ͭ�&�6�kb0��1�oeب��,M� ƃ�9�m��5����a�X���g �eր.�-6�h��cn�����i%z��ܻn��.Ƹ�l��$�iŕe��z"p��9���^�h̅�	����拇+H	�Ж�;&2`9����e��T4��Guyl5jRwt��F��XܡO��x���{a�ȥ��H+S���wg�`��,I��f��J���lm�F�g ��LfcͼܣH5�T�ɬFd�r�׎bZM� G.:��J�Z���-�4��ª
�R�
�:�f6�jR���ql�v�$Ū�ov1�4��э�.ټ8�Q���l�R�]3x�+�)8�ա���(j��>%1%G)�%C�H��u�z7�Z&T��ģOTSEn��d#��a��T�aWD�!jc0�U�Q�D���!��F�f�y�C%����l,oH�٘����p��I�!͸�Ⱦ6Rq�$�5:2kE���� �7���Pӏv�;��"J�tɩ2��ef-,iMЬb��lCk7n%���f�-�IlGi����1m8�^��')�Q��v������1Lj#N��Z���f��Ɋ�ڂ�
)����i�	����i�Z {hK_"jR2�����A�tܳ���2�ƛ�2к4����[��5d�6�nl����si�D�(*5���b�L�k%�vˋ.!�;�� �Z��!�z�7�=�[[E����tݘ=
��s%mկ�K����c�R����dn�z�춊�n�fغx&��¶���I��B�VE$#*��.�.k�%\Ű���#RvosMe��[�r���2�$I�pң��*��	D9ۂ7��b�vf�.�a'�m�A�zh�d���h�m��4Xnh�A�䑫�7G��h�1��mYs.V�;�N�՛V(Ql�#�S��ĒNL�*�s[��b�[�s��t��+(��)5n�٬hh�ݑh��&&�6�]�Ʉ�ʰ�Pq�2���֜P��.;�.�`UqSe�E��Fᩪ��Xo6P;S�
�)��ЛC%w[XN5�ҋq�t�U����a��D��-�eŴ�:���p�Pc�&U��e��zj�:-��ȴ���,Y?7c1&�S@h��$B��`�R��0\��8 �5P4n@�@��yp�yF�Vɡ���v�l�����"�4'L6��'ڹ�m� ���2�j�x�f�7���,Sφ-,��o`��4�GM�3j��1��Q��;W�k\�!U0�⤄��<�bݰiZB�Pj�kn�p-�+1�Zf�6�kF���J�d��/u�[U�Ua���ʇ$Qt\��(�oM�N�0�90�pT����{ XzV�@ݩ0�Ǘ��2S�Ȇ��c�à��W{ �'2����(�2°�F�Sui9H�'ټ1'!'�$�(���)�rd��\4�(�.N���u*�ܚ�D�:L0���6�(��rLk�D�dy�m�!:q�3��0�e���!�1R��#�����U���r�0�'j�T#7�p�Np���W�[:���5�5�d&$՜�Qqˢ�\��$�"
�l�d�5dTTaPrI�D�
�S�&ܾ���9�����+/��������c��"�5�����R ���d�к�l븚F"��O*#4�=��V��C͜��U]Y,��khI$A2Ii�������(vʻ�.�(n�0�76���Ph���"��VU�Q�!�ӄ�2���u|M�ɍ�=@���ԙD���c
$A�R2LA�!��=�H6���� �j�A�����$�o���=?���&�k���ʿ��f~�'b[Vg;�Z�ᕇ���^:'�{���sʘ�L���'TfpC��R��Ž�����{L�fL�y�+�4`\��\���x���LY�UG��̆���)^̟v m����D����Mv���7%�kUN7�٬��!Wu8�'���=���ܓDL�G�m������b��A�ެ��$�~�u������{v	ٔ4�t�m�Szs-���Y]k1f���9�(�mwS�1��+Na��	n���D�wtv�٧���)�nA��w��d�7�<�.��ѵ�;~{].�����6��ݘ)���S�er�Nt�s:��+U���X����d��/� ��ql�mgnk�������Y���w�S�j�$ý������sVu�Z�����U6�`��bl{�e��Ѫ�C�sG*ސ.(w�h�gd�^���XZ��%_%[��V��Kyj/�A.\SA��U�>g.�u͂��T�����}�^խ�h.�����d�넡�{ޫ(���.�:V������{G�F�̣I&�6k)��Z��>���V�{Muϰm�-�P�:����(9B=W.�k{6<��m,��G�(���ґ�컦6�_����{�*ϡ�����/V-�G���P�͍�����Ǔ���'C�}�%5�ɻwu�������$t�H>@#�˄ћ2�W;lZ�za��"��G"�Q�Ұh�F���<qǵ�y(�d=��wX��9[�PS��7�`ԎjY@��Vg�ͮ���^V�Nj�1��t���$�F6��2�T��y�-ƻ�e�܍��v��]�Jl0�o��:��]��W+۷uǌ����K{O=��wI����<wh}+�+e�{�EаTWl�<8G�mn"gF���WF��j�oq��t��r	���Z��w�Í�1��2�u�L��c�қ�/v�ދ��������Q�H*�v�5����ceO���(��S��Zb\sd�LD����2��U �mW
A=Wc�أnEY��[) #Wd�Zkn
�T�)��t���8 Њ�\���B���s��=����)m'{/��V�.���o9�ky�t��p�H=�aN��Ѹ�T��G U�E͠9e�g[&���͚�ҡR�V�`G��gp����R[=M��yA؜�+J�P�%=Iӭ�9/��7@�;�2�a&����`����'t�%WDC�XE6
]�:o1y�;�z���k��L�Jܦ_v:���6�1-]L�݊��n�J�7��*�ޠZ�9BW��
ܲi��V��gJs����r�{{�Hڊ!�a�d!I����}��E|�.���y�Ys��T*��c/q�2� �/_s�x �N������Iօ�]vգ2�m�m�=�"J�m k��=P�nU�|fY�P*���%�jj�G.xidIƛ��p�Ŏ^ݍu�y�ť���W�udM-���j��|��?3/{c;j��ĹV��cJA�g3sM��A�S�u]S���p�`РI��������i��BV�I��Cul�%�K�ݚ ��i�S��L���\���^�����8�@�W���7��l�ʽ{�e@�j�k�je���ei�.���XGA)�kߑtM�u�\�*�v)�V#r�`��:hR�ue��Sw��x�*˜���s9{�7��OU�59v����G{+���]mǈ��P݀�������Ζ�ָR�r�ҏ���>�r��t�+=\�v�V��7�-��X����T	�T�l;o��!�P�C����ƨ�e�K��v���]p	֔������S�*��o>�'�j���jyvNc4G&Yz�����-Z�q����Lzbˮ���lPD^[�����;���rnHY���A���`�,1W����:�n�Eg^���xu����P-Ύ�\uάO5>Uy��ڙ�'ö�;��Nq�D���K�@LV�ev^���xw��m,�x{`ގ�r�b�S�=[Ҁ�pE���ܙ�m��C���䶠U�:��G])T;��a�G��ڌoj��Ucs��uą�IB����#*T�0iB0��j:�ʀ�m�-��y��j`�ϔ��v��b6*ۣ��j�M���*|Y���hp��ۤ��Sޛ�@;�[���z!����ѡ�|�m��m�!�<��K>���X�:x�����sX3q�g��5a�3�'-J�ƪ�\qe��w��|��(_u;���X��7��7�n��4��Q�*�r�;H+�^AF�p[x�������A�!�jf������ ��h��n��h]1�ڝm�v��WuϹ���ջ���L��;�(ے�;H�pG�t�4����FfS}W�Jқ��Ԏ�G���иIم���L��.�	ְq��V��T�VMz��5�tT�P��{ ޤ�k�M��3�;��I��X�COo��w$�F�Չ�/.]��F��K -�ﮆ"�p���������5X�ݠ�t��=Fm�S��0��ݺh&7݅]�v�-��ŭ��O!Y��z�<�O����G�h<8]��p��6���ն��;�ގ��P�Zs�H�ܩ����E��b���M�7s5���Ԫ3OUӺ��b�}1r��r��{wnWw;\֦y�
T��(u;k�(�;CMm�X�����YO7y���s����6��vu��;I�Xv�������;��I��Ex:�w:m��9P�7mF���f�]o�n��h�:5���g���N�]o%)��U��5ǖ �r�z��c��eZ�"�[�V�jV�ݪ��-�ӑgE��u���۸�3{8�[�j�q�j�Vt�,=G��̮�7�v�!z38�U�δ�@ک`�Z܅�Т�
U�h?0�,��*�#[Ea�/o4��gEx��=բN,Ѯ���R�p�#��P!�5p1��m��;x����}�vv�Y�iX��ƴq{}{�ϢB�O)˨�m���{�<�G���[9�7k���Uղ�q5�A�ի��]���R�**�����K��4k�o����7��B�-�S�3����s?o��[�:S�c&wla��}\7,(���VŇ���G ۊ`V����]�<\��*-�u��0�`����Gf����S[��Ā�֮䛴��:�Dt���� {��2��0`o�F(�ϼ*�����Ю�'���t�|����f�tSV�7� ��i��D���5rT�8������ݷ���Ś��l�i�� J�œ)R�
�Dz���\���_^���{�׹���1^���j̱ݹ&H���/.(����1|�Z�m���w�ua��G�[8sm�)�C&^���\Lb�fMzRm�z&�9d8��]�żIV���e�q�z�;�;em?�tO0�R�~U���і�e�h62�7|�)ە{th0�U���L���&_.FSz�����:�eh�X�3:�.�d�3�Mze�P���m]��uM�]��ĸ�K�\�>����,3����0f�ͪ`sN�@7V+�A+�5]Z�s`�%��2�z7q��
��7g� 78�����M�ꬾ�Dޒ�b�1�58��ڡηݽ#�N��t� �C!.Q��M�|���F%/=�ܸH��3j��{���=�6�1��u�:g��2�95�3&����3l���6��oQ��T�uڭ�W�ʺ%�@`��^����T>������#¯t�*[�אC|m-	��nyޱZ���dR*���5� �>Agw.W����i��K8ε�F�Z95m�4ʳ���j���G�;�7)����V[T�H�5��h��;X�Qñ�ȹ���;�:%J��\�#��Y�0�um$�L���u$�()�^�G���R<tiWi�,q6�Ó%�D͞6��lr�NU�ۑ�������Z�`�tN������=W{����=V��9ۆ�W�)�1���L|m��1o1u��*�u:z:bQ[��K���[E���*<���uf���k�w]û �n�/���uo-w���]js6
Bd���aZ�O�(ȵ�㱹:�+��^��|����\Ͳ��>��3���)�{D��Cl_H6l�tv��/�fQ\�K/qоm����𰙻���3�u�0u�lNԢ�>��I[�)gW��:�Yy�C'5��
0��[�6����3��=&��D4�T�;�t.5�\�ljR�n���w��^�ִ�}{��@�R7B��ޞy����]u�L�9[��K��_۲�K���g�� r�k�D�s!N�l'[o����msU+�׫�7Cߊ�]bP�>��tsv�T+��^VfAb�%Q��7�)9=���+A�Iљ���ώ�F�aԩ���K,��-��5l�C���2�N�bcA���A7Ǵ���������U<�A��T��$�����7v�?�܇����r��mR�e1����2q{E�,�<aPs� h\�m1pk�Wcn$el�Z�&���S���H�\���ͬsd���A;.���0��l��P�[�u3w*�4�����@��'�`����V�{C�Nm� \ﴉ9>�P@�y�n���Cٺ��W��g+��1|��;��$O
����z�+�����m��r�NulmK��q������-�l�P����S�i������K�����k,�͡]y'�/,$͡.�}8�����S��ٽ ��u��T�:���(
RJ]\�Ӭ38Jʷ6*
��9=~ƺм%Mk�sz��G5�LM�.�n�P���B+�LFGa�5��ٜ$�w���1��ڦ��r�i��r��Y��u�i8�:_����N}�Q�ݾ�f�3�ۊ��x��W,��	�u�c��C��x��Ѡ.})+��Zr@:� #c�f�KJ�J�DLx��X���@@�V��Z�8{(V��Z**���m!1V��q]�5u�m`��t�'��XvymU�f�B���vO�B��S�Z�q�o\�X^̨ �lFa�6���ti�eJػ,m�0��ˤK�7��"h#s�\���:xTw�N�z��]Xi�{�A(���J�P�n�/�Џi�qahG]�k+�rl�J�#�E��:*��`���}i�"�yp������&�v�z��s��u���t�dS�ɕ�vw�ybJH����b�ћ��ݹ�� "�Ww��/��a�T@rG@彺��f�-K\�)}LCa�ڇ�h�M��%��hcroga��98�Yr�YVo1�t�8-Ev���:�SNT}���HjЕ�{��t�KQ�T����|��N^:7��7�8�z���^cp�"[B�sz���'#�ܷ��>�b�HvY�[�6���O��Yst�������ye���Q��/g_]��-��XtTڴt���(bB�S��o�W[w��n�knFE��.3�F��[�%}3L�� �u�o�0d|E\*�!g���9�"
q�>UR��.Kymݪ�ީ^]�-�-5R��������[��nVr%��a�䭵ۉ�]u��oh�#��b�19Ţ�s	+���rӭW���W����L�tD�o���8���U��FT���P_n��kh��zS�)h�Vq������M�](�a��¬�`�Ծ��%w �c�^(���j�l
��(�/Cӡ]���Ǜ4���j�ܠڔ�g)Ր�u}��mۆ�������D:�|T�E�q�խ�n�c3���N�w;��t�yۼ]!��wCn�CT�{�,�8�`犮���?�>��k�0^��+�'A���vf�PqΡSY�;M�x�>ݜ�m+��nb����)��^�N�h���i�:��@Rt�:ΝLSYɚ����J�1��f-�Te����-��NV�OT�A|{�5����&(J}���O{�ް*��$�+�����u +_k�^2;(^�W�;L�����u�i�
�}��v��>]�y`����p{X�7n���3�jZX��Z��pl��+'T��>@q�7)ڜ1��ڐ��w�#]e�u����}��b�]��d����z�t�]C@�p�x�[���6��
���Z܊����Hn�7񃞔k������&�|h�ńܫn����Q�����Ԟ�ض_ZTɡt i�c�B��u[o+����m������]q����g:|��4,q�+� "�ϻ�9ǂ����o~
�s�Ⱥ��7؜�!��a�o:{�v�\P�Eu���L�]�L�UՑ�sB�7��Y��������:��I��{��d��Kx�gb��o�b�omME�u�W�D.�N�^�2�eL��	+9)x9�S�`I��No!H1�y�uu(y#�Bk{9vf�*�j�a-7;Na�aK��9�vW_X�ޓ��&(|�ؾS�����_n���<�[\4֧]���N��ug��:�s��+��7Li�n��4ᝈ�9��I$��I�����z0��<cX:d]/�л�|�S�!@h��P�Ry���>A�y+�4��S�y|��hOs�C��ɯ {����G=d����䴇��!�C��~��oX>����(y)���H�AG�z�M0��@������O'�]/���|�{�"||Y>/8S䞡�=A}o�Ov��> ��r{���'�XO��u����TP_��?��x����v.��� ������ *������������~Y�w���}��
�U�{����U#Np�o%�� 햷t�v+�^`�fIt�h��p0:�Xw�s1��:.�^ӰVK���6
0{�Io���St±�r�q��n�u��!T0��C�q�:�� d�q�
���J����^�/M��5e>Q�zs*�H:��~Zj��=�|��Ȏ�]5m�)P�=�`����#.��;l�O�"����Ҹ�R=����w�H�
�-�K�b����BC�r�t���s��tgp��гtT�)�`X����}|����dD�ϴ۠�Քh�uպ\��e\��X��%k�`�̍�7J�� 责S0K���0d�x�SFNʎ����)�M
|���x���������^3�Դ�ؽ����ה����α�eQ�2�����CR��Tz�Uw{��^I�`�ک�q��Ӧ�-��F1���7Y[X���j�v_�G�7t8[Wus��M9��3�6�bN�Xk�el�8�r� ���zڡn�s���ᓁ��7�E��+z��O�5P�cNަu�N�id����jbA��/*U� f��)��]C��N�d@����V�����Da��×�}�m�M�Όyq�%8�u�\z4��8yhb���h�v9-w���Y��bx���n4����.��w*YW�z.����'��mve7��w�����W��-���EK'�1mv5L�y1�¬2�L	���^Z���cYL�wC�2n;b�F@��Q4`&�ڽ��w��]��8E(/cʲ�iw��D����9g�O�7w0[��[%*;�Wf�o�����o�73��rI��ҁ1�V�˼|$h�m�pܫ�G�X���d+x�v뽔��J��x*(E����(�k�ViJW���H�>�ItIm�������t�Λ]]r�{��Yպ�9�K�;�:5{���qsv���m!WQ�X[g2ve���L��kn4�1%G-U��3+��3B�2�^�N�c(+�`�֫D���`�捖��b�� �<4�v IQ�t���B��^�V�))y�
c%ٕnk۱|�������駁 <��\CY6󥌡���z���r�8�#�v4 ��Y-Hu��-h9����L���8Д�܅t��i��(��"˂���Q��eX�SYp�b��6�����l��X�w��7.�\?Pjo���E[�P!�l�2&�|����5�Y��З1R�}���a5En�p�HǴhEyI�M��Bq�o�Q��E����t�� Y0*���I�Q3�lݟr�N��Àس�+"�w8|��t�]�ћ�{��j�.�s�PG�*�3qڢ\a��ǠP�L���N�V�LQO�6\�6vX�wT�I�Ѹ�<�][�+V(qJ��!�pefKw5s�)�t!Uu�*cfW̍v��(��v�����.WTs�vH��T,������9+�U��շ8�Y�M,�E�K�ag	E-TS�WW�Z��Z��p�q�ʹwO9��MѴw0�P���κQخZ��y� �y5�u��X5�sst�E}U		��{���\F���5����x�]<�F����J�t5����7A�Vl�dV��[���r�[�%-�ٴ������r�t�V�L�L}k�u���ʇ�o&��lg�WGqu]�k��,�R�6s|s6ۗ;0��th��vyaZ*[��R���WYo`�)�h���r���lpF�޾�,��ά�.��˖o�\k�Yz=��]�[o��s��u� ����|Tt�:��n������)�T��F��qݓګUua��1�m�/UP09e����I����b/{8KUƂ��#VD�-ԨR��*�z,'A*Tx�m�d�u!�G��O���V�cwj:���#�n����h�7��B��T�!��0#�V�eQ�����\��p�*��t�IFvڬ�e�)��5�;�'*V�4���
m- :�"eNR�G�i*�����W9ge�|d�7u�Iɋ���Lv�}�l'ڵ��l|b�4*hQ�v�:zڝGz�]]��8��LF�6��KpU�+���;'�-��������0�y��8��*�+�EV�K���r�2�Z�09|��@E@6+���Fw����l�"sE�\O��	<LV���MՆ��l�&3w�~�
Jz����.��J�W#oT��9����-��B�j���k��q�sV7��&�+�ol.g�mR�:)+�`�T���n���H1�6���K�+,�o x�o_JaU��pfP��\\�W�^[�:<�Gd��$�e.�ÂGB�.}I�l��]�cvC\��*軤p����e)H��B�U�m뫦9��b�7��T��Q�\�l�޶�u��3d�OџV�|b�V�-�(���<�p�c(�Zԛ��L�.��@�6Lm�0U�r�nU�S��M�N4���Z˧h�>O���Z3�&�ȁ�߬v�|�1T��E�O���泃�;�F�Ev�n�ϫCEآ>k>AS�r����,��Α*߶�F�{8���^��	�V��<j�J��ʊ�6Q ��<��$ ց�@րx%c�f)+��+J�y+����FcM�M��;3#�+�αWq����@'��q�ǹ׶@�3����ҰO�`jV�'J� D��ӸE���<ӗ]�<e(k4]��D�ݶ�u%��v�@pL�dK
��T�veMh��6,[�A�u����b���:��J�]�y��XY@]�)0�� _�V[�(��u��Z�F�j
Dp�n��\˹�"��J@t�^SP4�c7�T���Aк�u��i����[ץ+V�l$ɦ�d��ލ,f�փ����@��k�/G�����-�4+>�X�K��i���
�o+-��P��z�f���up���I�<��«�|�儹�#�����%���|H��ѷ�"�wpݣ(os��`�]U��r��V�78��U:.�P�w��j�.C��n���5�R1洠��R���>{j[�ٸ�ư]�Zj���.��n�Y�����زԶ�%�L../E�T�n���:�M9o�&���.#�Pw×��2�aL1�ff�����;���^G�4�K�e@�C=J��kPw-ͤ[��ab��5�(4F\-�䜺]jr�d((�����K������)��C`kܹ(nʱ�+M������B��0@���]��Lhi�G\o���~hKn�mB!]#�0浐�Qu�ݐKpн�\��=d
���7�T����h�|�5���q\�$�웨a�(ue:�哩ٳ�����8O��*��2�H��v5ݧ���q�H�v�<T�RN�f�|j�{�I�l��ڼ�S&U_n�b��FA�6�52m�H�I�e����IvF� >��m�ߵ��k�\Q�[9��n=|\�P�G���Z���f�����z-R�k�*��\	�Lb����=5��V�-�Fv�U7�Q��ޜ�3��%f�3\J!��R���TU��JpP��4��6"i�­h�h;��ڀ���u\�%���k;c��,c�"1�|"����ڪTM�4(�z�`]����oH�%V�b�T5yuF�i'�@ M�/c��Y̟JIX`�<�[ :�<&b�2Ko:����t,�F�k���P�;�J�U�_T�Ǆ�hէ ��6F
�a_
�����)�Lx�v����D����Z��A'Zw4\I�]��9�n�����ذƣ� F�NSm�y-��f�̻!��΅J�qا��r �E��a��86d�X���u�tw0�O�uVFPY�(��W't�>����.��A\�������:Y�;�AR�ꛔ�=4��#�z�:块nf\w,��$ο�cY��![tw%:}�5O���jj�E\2kx��xA�J��z��������?��w�x�\�uʚ��[��Ǘ���$�\e�>�꿆�De�L�e�jZ�� ���ǥIy�V�shl׊�X��͎��t��7�w6]oc�Ə3/_݅��ۧ�wH��N���u���v�)U�Dl���0�
��*����539�zf�TcL��&�Dj���b���0�m2M��o#ۓ���?��.F��̚@�6,�.ʷt)�鍤;J9]m�F��e5\Wm��e [5D ^	u������PU�U�F2�[�R\V�E弔�ƨ�{��<�΍�*y�2���C�t��&��75�}���C]-l��SN�2@`RP�*[B���U��d,b�I&G��Ȑ�S�@L�2�凫L�[���[3�(���gK���ݮ�3�T��n]ʺ��]�d��A%�@_Z�eNψ��-5�O[�d���`�J��l��ܶ(���E�ƠD|�����Ζ��5'�|�Y�;���4;�k��B���u�X�erqYD�.����fw ��� ��dp�X�����d�LsBUh<�a�t�GB�;��/��v�*�mh}ğ)Z����1�5
���6'�w2�8�@�/k$�.�bk��b��Ze#����k���l�a�v���d����sGA�ޒ,(������R��"�U�c��e%���)�:as��\��������K�
�konʧV�ihr"�!45��%eC�9�T=�����۵�%�ҧ��O.��^���F��ȾEM�1��@���KZ����֕*�s3��������i�$���ݎ��/��D�m�L��[j�;JyFe�*�֨�K����~��߭ {��Etz�����r�m�[Q�	ڙE�S������xl�wWV�C)���>{;;[��A���e��g�eWv�UiTtĬ�zC؞�^tW�F�Q�Y��VE�Y]��l�(��t�Z:�/���c��:#�ZףA/D�����z�I���WJ����n�ř�#�kF	G��Ӌu��w�em<
�j�`���T잒�7X�n
�H�U�죎�i�-#F���0*�5n�Ռ�����"��Z!eџc"���g�3�D����n���L��}}��N�S�p�!
!(�n�����P������.����}3E��h#X�{�+S��c�Êb�f�=���[�B]`��}Re��6�Q?t#�����X8�Rs�K}��
��ο��hn�*�va�$<��"��><��C�k]oJ�%_ޒ�m��]ì�GV����ӯ`���A��qf��WX����j�V�Q���%�P�{z>GZ�hy]�$�
�s�@�ݗ3^��
��J���>����4�c\?.��P5/jũ��io��z7w6<#�t]Z53�hd-��X�oNB�b��w
�*7��t�=ֵQ�Q���ŽR�[�zs;��
m�jS�ʜ�^+�h�@p+넱Qԙ5l��:麕j��M����n�:�[��F�E����|��Ʒ�u�t��<kv�I �lY7��F�p�.��ki�h�Ĳ�l��h�怡\G&*I��n�gJ��v��%��<B��<��4�����֩"�8>9]��{�v[���0�eu��6�I��-�����*�P�-h'�f��e&^�9 ���;{)��)�
���
��:�A�!�ԭ�{+*쑂N�����gc���+�$��T�m^�먾2Q�u��əJ�GI������m��i�BM7x6���ffs)��s��ܕH�V��[#�|74^�JP�c0��@�z��*#Z���­�u��(��אط{��RՔSR|�NT��L�r�n�6Q��L*|m����!�[���N�� ��t�Q��v����d��\X�]�v9joj�����|�on��ȩ7��\@�̞�+�^�o�hG;*۟>���O�]]�]P;���Ϝ�ȹ�%�:h�Pw{����p�!n�&X�g"����?Ksm��{�����T��w����(��:��lw겸�����7�`�P��A�Z�m0�ӳ�:��q].|F���t�1�O�Y�c��Y�����*j�9��< �>
2�p��C�L�u  Uб�4�OX��ܒ����wU1�%���f�k���x�ۂ�r�.�wQ{S��L�2M�@��ޮ����k�|�yI@X\6���@�e�f����Mu���#�)Pw[�8v�T�������	��Цm�$iK���(4֛ņ�.��)���ԽÚ�����⥚�1��W�eʾ���(���㙝ֳAC� ��;��.�������7��C�@�'d�[�=N�Jw+��k���1�(n��@����q��j�Q�ZlBB�Y����;[{3��v��Nca�S�1%k�X��g��u�[����Ei����}���ˡn»����*p4b	�i%w��4+���v8��38�=[�*�eB$륥VPS��c!AK�4V�qq)]��	�#F�q�����ڔk�+���a�z�hKh��p��lxCn���xX��J׳K���q_m#A(����̥]niZ�u���feS���]Ө_��	Xq!�CJ�'Q[��J*��Kr�F��"�rU����]u㝹R�ar��B)�sz�Z ��ȕ؝p*��u��}��p���}{xEl����ͅ��}A;��bu������D���A�Ŏw�{;���������j>2qB9@N�;b}aĎ�/����6-ȘTo$���Q�N2�zq��ʸ	������DW�4_����~���w�/��/����'�k�?���}������}��o���}��o������������S�|o����9k�9}�/7��L�	SH��?~?U���A�H�(���D�� /ր |,ث%h �DW�K�[I�$Rm�HK�H���ׅ�7�<6��<<nm���k�m�a�M2Y  �:-%T��ر�V��@ӯ~[�K*
u�o����hN��Z��[�}�
�bB4���b���p*�u,��EN�Yq`��[�;aǤ�:�9���i]�o���R�<Ze��H�-{Q�b�w1B�3t�B��z%�͑D]��`.·)��$�ޢ���s(9�C�*<�,U� $%Z�ІRB����։@�(N����K4iv�P�.[�R
�+�S)���s�d�-*���V�p�t�WW��N�]��[;3�%���6�g]Φ��{r����Ijm ��t�L�U����N:���ݭ�S��+P���KO=�X�Fr��rD�ZScJl��p�p�xq�s�Y��ggph�\a�g�:YUj����M������'73/}�c�M^lT���w��Q�HV�����N�r=����8���\����+�n�Pܠ6R���jt�w�>��Y����qֵRC;4uJ@��x�
S�ܑ:�b�r䎽�}�U�^��M��Nir!)�Ma�ujpܼ��r�GP��=���k�t]��h��LJ��k0]���[�itUD���S	�z�$�
�/��3�����C+���vRb:Е7���a�B�����/���ص���=˥���n�d݄�7�}{�HY����%�i1K�a ʪ_ i.��*b�L&���B�� �e�(4�
�I��E*��-:6�M��"� �l���~ �!��N�N�m�U/�Qj��)PT
m�D�@;m��D�(F��YA�t)|Be�F���:A��'�&� KJ�]S`�M��|çE��L6)�
`�d���(�E�U�ҥimR)�i��H�,�A���	6����"�&��'�I"�U�I� �aG�ώz�|�����y�IQW4kk��ڶΌF�ͱF��1k$N-�8΢�����b�'Z
�m�c��UT豢�+�(�F�6ΫV-�#�1h��q*<ڪ�Z�UEm�&�ư�-m�֍���r�PTQ���&�6-���lFJ���
1bJ�m�A盕SG�,UFb�h�y����ͭ��m�9�f�m4Z�EV���ƍ�˜���ܼ�*9�Q�LDSG1���F�1�"&ums9����)�L�1��թ�j ������$�:��l�/9�1X��:6��V�C�j9�����U41�yb.lT��&�X�f(���rNF�I�G6.X���(�
 ��6ͱ�j�ZmY�DQ2QUlS�l� Sy���V��cm��	��l4�M�l��_��: ��h�m ��-.>���J�P�����VWX5鲟:�o�v�iÇ{\T$Z$M.��6�N9��S���v�g+�A�'���J�D2H<�0�  M*j� �WH�F���Th��:.��f�VU*����ݽ��lu��A˫����N��>�0eE���O�j��5;A�mvPcʾܴ�o�.
�����o*Q}�=�K�c�o���}���^�z�]s';��ܡ��oI5Yu��T����=�G@&�?W�V����뽽�d����uի�龖��}����/�����G�^US+�T~���w���z�no��'���]X��}�r�a����s���ܝE�Y�}���`�"rp�}jg����3��];�`wVϫ�mA���-G�+�m<��;6��W�>�u�������D����;�}�=x������6�����Ǡ˿m
�[���}���̴�.�%]E����%�|OoPn'��S�v�N�f�נ��2a��gE�o_����7-�*f�����	&��^���<�ǳޓ�P�󽷥��|S-�U�=�]D:�g��]�f���Y��e'�z/Ney����y��_��Y�4m?՗�qh�7����cw����,c����n�������᭧���c���zG/�5��^vUr.��j��l���(r�B���s��������7�b�o�V��%>٘(�뗱=\��9C�yÂ��r*��Ӥ];a=/mz}:�}s���>YP�>T:�d��mt9���~;�{�l1�~��&O�LU���k�ק\��\�7��=Ds��S;���١���ݠ�iۂ|b����o�-���˯�}�-��K��=�m�wz�M�;��{��C~���'+>z�T*GM�������;�l�9�(��G�#�α:{�7��_�����[��f��v=<��'N�-w��J��{�ro-�_?%o:�_��W��Q=��X�NvΞ�t�)%CW������D}R�wF[;ҟ�yA羯du��.}�9i�ק�m�d槽ٍ�/b7�1�M��/⶝׼��{g3&a��LGo�:,���x��W���9�]��� �/�S�a�V���s/"�k�����y�8��ݿs�@���?lʭ�yә{oA�wތs���.=�9��L
��cMd�-�v3��i��/�e�r�s�ܴ�:+}{2�ݚ���E�����5�f�����o:Խ�̰��[���1<)��gHm������askc��λL�W�#d����u_^�=z;��Hl鼋6���<�ɮ(�����݇��Ne���ٯ��fO4�����z�ᷳ��@��ݵն=�4+��]w{>�/�ݿ{��ĺ���m�4w�N[�3��ꥀX��=(/������W����E�ϳ� �����3���l`�kު>;��L*�(����K}��z''$���^��-���K���P�T�y��˯�M6�۪�_²:�����>��>�c}�����;z}%��zu{z�yFs�\���|������qu>�K�D���'�ϺE��=�3N�1�jr:$�/A�A�Æ�Lp��&�sI��S�_e�Y���
�y�Y��b��sxr���]��u�}j��~��o�� T=�C0	�x��[[�� 5�o���	�8�w��sÞ5��J^�e>�;�J�w���6>���}��6��:ͥږ�DJ��t'�]@���Cm���w�9{��Ƕ��۰ŗ�-\�/u�BJ�]�*�>rN��nR��x���ܜ�=���J�z
�E]9����	��urX�բt��L ��1$�J�r++��\�gQ]:f����Q��c�{ U��Uk��w�7ַ�ɾ#�[�����<�������9��|g{�X�y�|��52�2�#����z\3��^\��@�W�i߅��y��F�q�}=�,�H��s}Ob���m7X��5ē�'{׹r�E�\�}��z_�~��{���3��3d�S���"�{]�	��/j{�Z��ܟuN��o�X�����my�g؃o�g�Nqz��PM�Y�V釪L�G�{��;�;7��xy��r�����}�I2��yC�]2��Ϧ���(�v!����������m9�7��]���J��{�}�J+Uz� ���{�ꙛL5<m^�a��zѡOg�{تw7���}�"���ם��|��7�3�Ս���r&�P��~=wχ7O^��1t;Z|�oC�������,{��n7���ǭ̜s�I���{��=��T{���@w]b~t�p��ѳ��)���v��vy�~����`���vv8D8y3(@pR�&k����.�w���Ծs�Z944�x�o_)uf�H�la�*���;�봵)�7Wv�5���A����w��1b�}��}�A/B�a�J����?����ƅ=���<�>U+$�K,wJ��븠h���ʪ���i���s��!�Fv�b^ ��0; �מ;��n�������;���_�����Xx���������	�|�����T��x��'�3V��>�X+�]��V:������:�'��{�by|g�E��8����k���;W�]��ލ���{��z�ϟ�٩��c��_�'[��zss��<�ٸ^`3iw��^�^��/-j7�����X};K���^�~�-z�������O���Ԟ�M^�d�^Me�����G�;.�7��0N⿜N�|��?o_ڗ]n�{Q��������7��G������Q~�i�g1���~��ޭ��� o���������@wIݿwVȮ9� ����Ǩ�׼*��k�|v��zƪ-&�!b�@';�e��i|l֨2��B�$��L�'I��FYt���.�c�׳�����L�<|�w^h���F�!�6`�,����&�_�/��ȭ�p�2�]7բ�a��2�179�E���FZ�)�_&����
u��������$��7I��n��om�0l��w&t�ګ�߽���՝�������cդ����y��x�nh���r7�o���Ϟ� x>���!鮩�wݙ[=�91�zO5��$��ZR����s��ބ��zVj�(�h_P���-��.��zzp�wG�Xޭ�F��y{�Ӯ�޳8u���	�K@l� @�2=s�G&s�	�.�:}�ZR��^�>.-}�ޟn_I���$GL�!�@�af�d��	��W��q�.z&i����۾��)Qx��'8ט��/���ɿ���{aŸn/w�6�a��5��,}*p���P��ƕ/ݹ����umw����G�u<�);�b�(��Τ���Q�3ٯ�8��d��W^�M��t��`�ܻ���3�wo��	���귦��f�ϳ~/��7�o�K�����Ժ��@�e�ܯJZ���* �c)A�%�=��ry �|Sz ��٢mg<�듷&v��Z�}����/|����杧���,�tsebڄ�n�v'QY��J�����lmG�m��;4L�\lt�s�8W-�VP�v5�s̿�7�O@�l�Z����T;��;kyZz��?C��ӂ�D�6��W�'yh��;������PU�I�{+�K���*�}����e�|�!��d괧�{�{��V��=��_?g��O�Kw��g�nZ���������vwe�^-VG
�ћ�!��������eo�ʮ�sŀ�����'{��L�;���?�D8�֌��,Ǐ���G�w_���� �Z���m��Dz�My����z�h����Nx���N�ս�L�7��y[�������>5([Uυ�*�����c���3���]�n�z�|��P�L}/{zz�#�0���P}��>�&{�����Lx��Ͻ�Kj{�#���Q��V�rc����0O�Ew��Eg;�/�=�v�3���ϹI��������n:��<�E+�?��w�wE_��&G{Q�ۀ:�U;D�=���˵��jb��\[]fwg���ؔ�F�~Bt[O��h�,{4c0�jkq�*�����~���a^�w���@ig4������G\+�Ն�u�κ�K{r���FWv�N����o��+:r8_h��fY����%����YF����ܜ���폕�G��B�^�f�{b�w�'��-O
c�w~�mQ��b�ƣe��6����}[V�<=�q�������֬h������c+��a7{����W�w'z�/���V�$��NӘ[�:�kzϦЬ�+|���\�o��t��z�
�g��;�_�mP}��������AY���%-��g�����Xo���w3�᧷+��MT�W���:��=�y�|��52�)%�X�okz.����������R|Q~�O�Ԟ>�S�~����;�^g���=��t`yk�'�w΃�B��]V�}W��X��Pz*��9{kf3I�<����o��ț��Ե���Gl��z!�8����{}S;��=5-/��m��h�$�t��,�G�2�T�{;�}0�G��ڇi�z�(^�N���W5r%s8r��>��빍\wb�-�*1�\7�������]��@v��u�[��i�iu�#���_1���j����W1�i����R�
�\����Y�5@���o��h��v
\r�b��z�͠�-J��qI5t�:�Kw+*՗D�������_w�m�w�x�CP���\��=֞��A7w�c��;7�	�����}~- �v���c�+|õ�~ΩF��_ܯ��z��}���Ñ���y��}��=�p{>�o�Ʒ���}�ͻ�5פt?uNܒz얟@�׳�S$���|���=�}z�����\|3q.��N��������B��u�>��Omߺײ�{3�0�o$Y��~4{�&׽;T#����ƨW���w��Dȡ[��=b�L�q��x�Wi��wz��w�ʻ���C�[�����e��o��6'��d�s�h�KGf��\��"������/,ރݎkEm�X��Q��4��m����z��S�{�ٞD6�{�ƎOo��z{��v6y���N�=1;>�ӕzGG���+���Ǟ�c��x7ӏ�u�n<\�!@TB��D9:����.�j&��>��n����[��B/�ˇb����7���+�+}p�L��D{���4A4oN�`�K���S�v���o���k��8���`k#�+j�Ӂ�4��+'YdB��jl=�ɩ-��ג���ks{w�����K�a��_M>�Oj4+vz�xvMt�v�[�Y���<���z�T��~M�S�3�HMW�y�x��� Pw<�|h@����2�2�AcMo�]ݱ�=[>/�sW}R�>�YGޙ�����w��[\l�'�d�Ɲ���z|�� L��յ��D�]��h���	df��2N/_���=�U�`oM�Zxך;M3�۹���u�o1U4?o�l��!f����yߧ�<�w`<�υ��\f��}�v�y���s�=�CҬ뭫~kg{�}w�����*#�=�*��ܣ;�=��􏝼��.A�^y���9�Y>��X��R��[Zv�Jx|��ku����e~��A���=�wc�m�3����&�A�U�o*# �`�
+돵礸'����������m��}�s�{���&`܇��1���'ǿ�>�|����~_�����g���z�}�������<|||}�G�������ٜf�v{|lƷ��<gq�&�Y�a-]
x�[�AW�>�௷�\n�M�6��������@5i��pl��ы^Mk+��Y��*c�{�uᎠ	-�V:Vvr��q���LN�{0ɽ@��6��=Kq��L3�Lw�ځ��Vi�M�3Pb���J�\�(#��!>�C��f[�A����$��յ �\����M��IiX;�b�\I���2���������K˭���l; mkd6+MÔ��E�޺�J�<�N�
MXm��YL�k����Ω�����zw/����
dZ��g��K���w'�eo<��u��W�8���6t�-�YL��:��mZ%�鹵�Ǚ����Q4$n½=��(F�͡���uY:�lr�G�PXqJ���4R�wgb	G���|�o�z��*��D��\+-�K	�q�4`���Of�m�*F,����(^P���l�A򏖼����v��*:ۗ˰�wK�sY�_T��F�&�b�v�^$Ԇ=Uۢ��e�5Ӟ�N��%M�Jly^�����O^�[&O��9}����[�b��S�Î��{�@�]z��+�2��yA���s�]p/�[�(u[����'����i�1���9ѧ/xNm�y8�h�^��'�/)��s��֜�g�|�pͺ�V
7Qdu0v�W}Cl�N��	�5Zb7gh[���(� W��NP8o�e���t�� �oe�}3@��9���Ln�@E\
}̜r��E�D�k�9l��{��m����0j�i��,��1�}�S���wSz���ˡ�z���Q2�9��܏ ��%7а$:�=���U���D��eҡ�w�;�#\4$U�������<un���o�N
�>�Ѷ,�DNT���tx ��oF}/N�ǹ��VRź]�m�=�W˵9�H����56�L[���t�2�Ves�;9:L����Q>X�<f�T�K:������ʮ�uv�;����w�4��^6��p�u}O1;R�G������8���J�����Y]���pR�a��U����F�Հ;@T�f_j8�{��FO@�F��ҷ��J�,U��׃
�\�K���EG�G%^(i
t���]���M��w��k%��u�07�ok�7��ػ��^�+�63��y���0�5��J{�um�z0�D���:F�`ycwqjk;,�$6�K�P�;Q���ή���A��M����.ty�1)����N�k�
��xc�S��)�>Y�I���IPq�O7 �V�a�S�=�T��.��v�;c�ǽ��.��/V�.Ep3A�~�Y�'K���)�z�֧wC��F�S#mm���̓'R9�4�=�Ϣw;��_�OR�.����{u��S-[xv��˽�c���`u�,�;�)\(��P���|+Z�d��*&��cUL� h�?\ܶ�W���i
*"5��I�
)��R�fJ��א���i,b����-�A[gy�ͣTb��P�U-�U�m��U�ѣAZ�9^cT��AQ5����*"�i���6�kA���5TV]h(J
j6�^A�X4�SKE��4�jci�Q��vɨ�+��ipQ[���v��4SEU��6�<���N�m͗��(*��h�F��r���'Jy �N���((�����s��·y�\˪E��N���1[+lSMh]&�2h}cQ塈��������kl-QTQ�CEW�h.o�6)����4r�rM��X���Q%\ι�A���ͩ�.\�:�*��h�G'F8`� �i�c9��#�p��9sU���v���np�C�''l�gIpثX��%c^c̦�փ���Eh�m�y< 9<�\7�͢��8�k�A�hf��O.G+ ���?������ǩ�e�A�E���1n.�X��Ul��T#Vٶ���� Zn��*�RŶ{����U�I�8M'�Mޭ?��i�o����Z8w�"�޻�xh����o�uV�O�a�l<3kz$�f��0H��+:d��
E����sAj�uDW�ܻLE���"���h��$`��m8z�麄�W'VRd��٘ ��k:�lrdq%�;
qE��M�vX��h�ʨj�=N�\��*Y�0�8�P�개6#6q�2��:]u�ex=�G� ��q�?�SL/IlQ��{��὜S'N�wt�g##�a�T��̌��y�*h�ywxm(�Ҝ��;��Q�L.�縘�� (�0�.mAE�]���Ѓ&�Fi��ɖ��W5ީ����G�)D�c��c}��>��)���M��d�������z���t_���~��h%9�w�vX�eX�o�wE!��6j�)�Y29�v�����_F��^˅]�ng���O݃U6��kh���p8ފ��k����YY��obg,#���%�7>и �@�%��JUL@��Puϻ�P�p&,V����R}�k&��p�w�d��VІ��/���/ "��~Z��5�2�"�����ΐ��?�SϞ��z�V�P�2�>x���OQ����+�]��1b�{��ݮ�Js+8�mF3��"��{��W�7´�V�6�pق擢��ī2)]F� �Z�Iט�&�3�ejbٮ�v�ms�z;f�n�ˀ�}�#��x�C�'�L�{������s/[ց[C�`k�g��[#�K�/	�h�^@�R)��6���qO�`7xÍ���k��2[����mN/���2��~��K�x��:|*�n7Ե���Y��C8d��L	Em�6�l�����\����l��C�9�����ޞ�d:��<����H�^PUO,��/6(c�y�j���Mrput�i�
�Uk����\��sP`����#�����y��ݤ�)��H~��ī����Y@�<e���Ia��3��o
�����dk��&�x���M�j�#�|z�����]����,'xx���V4�����{����v��7��&�x�����?������O�˨p���|��s&�[M�<���tl���ۭ�p�$�K1~>��m����C��3����^�<�'�_��f�Z�p��d��a�-<#ze�چ%�8�7�`:�t³��m��':%˯D��w�G��y5��ۘJ�����^2k�n��:�m�^��t�y��	e
�V����$�5[˞�o��{�<U9�o�'v2�&(}u:7�f͍GT��OYhgj��0���[K���(8�嵷y��0�rރh@ j�
<�Z���.u�)G�|{�WSˎt�v�aJ�k��jr�m7sj�˓/w^�o����W���]�������ba���ZzI ����ߊ�y�2W.�s����;4��s�\��QI��3����vZG�9�L��+D�����u�0�Õ̀���E��4�ơ�8�~fR.q��ڣe��I��{�G������8RT���*��mi������˳(=�:��CH���^�>�/�R���G�0�Tsx���.'g�r�Bj�!7>��%�'��}��⯲�О��N���YK��5Hz�i�~5JP��}��3���b~��Fܼ@g{A�J�0]�4o<�cǶ��`��e�K5K�ܽEy��L[�-H�R�n���ڋ����SȾ�^���q�JK�O0�v04u��aa�@iC��%�[˻�@��JT�c���\�~��^�
�*���i�N�K�I���kd��KKՊ�Fv�s��Ν'��^]���������E2|�9�ޱ���q)踠�\��8��P���4�bw�v]�j��˙�ѭ��1���mx��k&Z�D�n�ͻ��m�6�����JNCS���I
��h�E�f#Th�+��W]yP~�uL�*���O�vO�����g���fE x���K�-�b�P�b�N�}�Gu�ad��]���u@;�/+r���J���v���Xo�{X��|�s���'NO{E4,ebs�G���Ԃ�Yf!,����lp���h�1D>ʺ���fvt���:�w�Y�|�3��k5ӭm�!y�����؂���������?�3G�Uss�4:��/�Q�^Α7*w��{�a��핏P�����xYΆ�?8���$iݎG���!���c�S�Н0��-�������Rx����#b�;����&��d���S�ݪhj܎n��9B�℉��X���WQ~��gp�=�+;{_8����t0=�A��ך`P��kۂ�٪�A� %�25�U"m�;�(��O#ڟ�)�����\�$sNdù沉Ɵ;�[K�g`e��P9[ǹ��6��J�N[��ٸ�p��t�Bj{k�k��IX��ء����za�Ԛ"��5F�屫����JG���9��[z�B�T6T��q1X���Q`��2X��Y<5M��Z���3&�uqN����l�&d\
�m&�A�Y���s+�@Xd/�C�ʢ^��'�0��O1)M6�Z����ઞ5��	`�}��y�����sNd`{NŐ��k &�_t�<ޞ�N/�H��p�y�Z0ZAa�V�k���l���s[Ww�m]sh]�_�I�`�mrr%�ڞoM���=ʊvO��v�>����e��''VL�2��ҝ#6�(���-�(��UXHZ�[���gvu�'s��-ܷ��d\�h��;HZ�^�j��z�Rkn� o���E"f�7�boQ۱/��`��e�贄�g8&&�7V�|#�����]����v9J���rD+�h�a��c�,����<�\,^	���v6L�ϯs[X��Qk�����4]��F¦�r"��u�N2���B:9�Z��s�6�������y�(<P\j����U~V{�c�P���<�-�Ъˉ�����o��Ѐ]U8�y�]�t0b�"#��O��Hq�����(cK4_4�N/! 4�*�ۆlF�����F��kM������y{#��w�>������mR@m~>T.�Y+��'9��9��h�R$�������፭@�Yw�20oOV;�Pga~�>����g,�Gu��,cS�
{hd'L���%��=G,3��h�q�x7����m8v��6�j�U.b�VoY������� "]�(?�����v�켟��˸kz]��\�|��z����Gw�SM?c�w��bǲ�>�u�dS����"ৡ5���6�g��]��w��{������4;Í���M�߿K�����S���k�&�e#!gߝe���[C��5[>~7Ժ��*Csv��y��]����3���ɭm̶��KT�<6�Q)�sH��W��,���}���'�N>&��ǥ��cC]!|n�o��*�l�/�>�<HE]�_D���aw������v�6l� AC���q>�mf�;r᢭���؄GH�Ns��Ҳ��yh.�VP�N�m5P���8`�S7��2��qO�f��1�*}�:����ʧv�����,�Fb{��|�5E'8�Kf�9�|�%�ٰ��&�F޵ƹ������@�]L7/5�c��IR�CG��Xk���\�U��%�,�,ڛo`�%-��7\L��>�7GԀ2��>�Ƒ�&n0;Hҕs78\���|��\-��{����i4��5����ʆ�0,�|q��xE�K�b�o�E.��Ҫ�&�J7Z�d�Ek�,oSZg�n�B�l�R��������Z	z	�UH��`!R�/N�9=V�]nJ/�S/�=C�}+B�]�:���h�$�4Il�l��hs���h�N�N�$��H�غ��z`�_�姝BR*��a��%�:͏:�v���A�cF�f��`����]���Ҍ�ިt)c:������ XؾynF�<�n2]C��/�U3����?t�]IV�S�3h��Ld��`u�膠�M5zC�~��gH:V��F�C�;���5��N0C�lɗ�[ӷ:^:u�E���z*_��Ck��x;@�^�:nU�͍�ݯN��w,=>�k'{I��Ytn�!�t�LƊ�ur��Z[��P�q��x �a��Y�l��<b��QC7'n�Ge�����B�H�3�m`'>�._J����u-������u|�a��w��ά\Q8��E���){�<���7�o^�v�؝!�³ST�Qk�ڴ���l#vc��y�6/��!��~|�>�:�bbا�X#�_�0݊Y�_�M�i��w̆��,�ߎ M�3��3�燗��_<9�"vX��NvMZ`�	��ԍn�.5�ˁ��j��^���9B��Kej�o;<�7e������b�" ���cck�׽���N�5V��_�mkL?":�CcͰ��U�����z+�j[^o�k
j�,��d޼ܒ{�8A�j����A��a�qD������֎���.�����b���]�����7ؖu��wQN-wmC	��dh���H=��^������[��Y*��Q��j#�Λ[��N��gE�s{�i���
�@Y̺��q�όF�i����0�=C�\u�s�oz���f�4
�-b6�3PՕ8�y.x~��u������R<f�e��]uNLPÂ��1w�xvXfiv��t5tWef:��q,8׳�fr���a7'��<�8�xc����X�8@�n��.�0{f/:�wr�a�9�:�b��]���㮔�]�̖���C��V�ga������[5��__�_�>VQ�t����v]����a�x�T��N_��[��gDg����^�~���<�`�=}�7idnX3�U��������W�ή�l��m7��bm�W1�˚q7K*��y}$�\Xj�������k8D�?�����⯦�p�o�Tsl;��sD:O��٬4+���ٳ	�d�-)���̃<�a�O�9�!�˭v�@Cy�0f�?�K���O�*)�����x�T2�Rc ֞���i�Չc�G]��F���q�hO\a� �#dK�x���L6��4ɺ�����f>���q����m/v��,Q�o^�M�[��t���9�@o�Dq��o\Ҡ�/g�q$k=��k� �̱h��kJr��:�����_3׻���T����#��|�v�|J�>�ob���vr�90����ƅq��z�0����>;��ŬWK���c�H�>�U��M�'�f]7��CN�gJ6	��`�kh�*���tW�G���[S��pU>u[�ö��t���y��p���c���}}���;�`��;w6M4g����Ɲ^�X�(S��{z��m�J5M���Ǆ����	��OqSJ�{�Lٟ�b�k����7����ZEa��|.;�Hw��c�Mp��z.��9HȟsOt��pCUl4�u/#�����_SS�f��άa��wAOT;�i4Ob�9F<�ȑ3A�-�=���(��G�r��y���rC���N�M����otP�{��J�ow��p4+uc��=N�%�)E
��淀��Z �{�H�r�G'm�ܴ�5�D`�n\�}�+Gv����X�}6_(��9��ga��Ԩ�j��,��o�  �y�{�o=M��μ�X����}옞aIL��%T˟�yV7^d�m���Nz]A�׳P�Tkz��q�P�nf�5���|nE���H����L-#u�ݡM1�m�����z���,Үr)��r2�G��l��ʙL�;Y����P��&�_tߚ+�z�8�?M0W��\W9nNX�
�X}�2��+�ڋb�<(�u��O�Bz6�e7���I0���6�vO����W<mªi��j��F�`���2���&��O��5*������S��ὖ�ן���߽j|j�z�WR��-�q���l�-��^И�3У�Bֹv�6�h/�s��~]�2���*����Q����M��rIz~�©'�1�7e��`�R��Z���v����Ƶ �@0�����~��Sת��&oCt�Ǥ�(F�O�;�ُ��!k�_���CϹ�3k�v>pz&�M)i8�淉&HjS���5Oq/��\�� �����p�ŏDw�20tW����,47����ZOu��������x���?UZt�Jj��(c�gH;��Nu3�6P<'�o��b��^W�qX��*C�_��\ͽ��0��^7(�gw��J[-^kLk��+�iB.�oH��6�U%���C)�avS�ds���1���]h���؋�U�n����$�}�eK�5��:��]k��9ԇT���I�OS��Z�G��{�3x yE���G���X�^ؔ�SY�lC��Ax��;Pze��"HUen������7m$���7�s��롙�nJ�L�ٴ��lb��L]��1�d���5 CWù�S��C�/�q:����b��t�k���mz��6X���a��J}œ<]#��}��:Yt�E�^=\���&yu������i��M�<ν�H�����4��Ks+	eSm����F/LK[����
\�G)]�x��<�M�b쫡G�":���`k@��C�[׉�N�����Y�-���|�`��pa��
^�눚�X6�N'l��?�E5��.�C�4]���d�\1��_�뜕�U 5��b�;f�4�{bs3;o�2��<�gV��Xd˭]`h���z�t2}���f�;U���øE@`�n�ٍ�5z��4-"e�j���id�Vؖ��{v�~��1l�ɨ��
Vϥ�JX˖<�wc_`��*eB�������{z��z��a&�B<{dt3��/)�?��F'f�Tmd"_9�0
����sBt�u�n�BƊl����m}x�r,}����>������޿g���}����ׯ^�~��^��o<x�{������f�[�b>�(�Hԍ������s�n����YѿM�q���iģ�c���ܔ���Ff�.9R���V�8��C�m�:������9�໣��([f��m�܄㻁aA�{���j�p�����Y�æ��ˠ:��v�U�Y�.���/Gp%��})�r��̗E>T�o�g�`���B�i��m�ǚA�놙r%
Yf��Sv��;�BL�Q0��Z���ueEW<ޑ.�,���� bi��
�f�|�]��1@�������<*ۉ�LU�F�!է>t#�rj'���`M�&c;�֕^|P�R��Fm���o��i@^�Ɂ��G^�P��̂�=�V���u�޼����_ms�we0B��{��(m���Г��=�r�*ۭ����|(��A��8��c/*���y˻��;���:�}�_LAJ�&��֕��TlH)AR��U�]\�u�jɧ����0]$�P�{����%��G��h]"�o���ͫ޾[buc>�OJ ����x�y�f�cg��up���Ѧ�b�;�rw�j{Ź��W[ViN��P8��6K�wv=.4i�r���*R�#Ŝ�փֆ��t��2�|zP# -���K|	UtͮVkyf�=ą|DGܛ���Su��H���0��yu_r��w�:r�I���#7k��N�H���O	Z_J�Z��5-
`R�����\hT�)��3F�3����(�o:y^�f{g�}@���ܟ?sĉw5�盻C4.jsa̙CE;���]Q7��b��ZM�>���ƶ��u��� ��e��ܯ�9}))GG,��8Wf+�2�P���f�t�5 ��΃T~w��b2���I�>$����eh��:��z�-)n1N+�ç�����^���:�s�@ڷ�M</*��uU�FtX�=P �V�At��TM�(n��u�Ign�4��uJޤmQ�
e#b�����*VT��Mr�zzs$P���o)�7Yݘ��p��a�V!�}��pӣ81�k�{�;nWNWZ"Jp݋� x���2�jxQ�aD8�Ӈ7�����ͳ���=�ż�=�
�u���m�ݎ�t�D:��>��NW/K$� �2�!�5��]ؤ�-���6<���������ʞSb
�|<'���xOl��������;Xqh�w�Cԍ��X<�=�|�l>�ۡi���B�֤�X�w��	���U�[��"ۧ�C�"h�n�3�mS;ξ�u�o
�u�S�����VC����2n-
ͤ�?�T6v��T��p�Wg[B�>A	Ky��Jɷ���]gLg;����T�l-�(��9��q��;k�wk��X��os�D)VseP|J�VT[��tzÍ\�V�{#�����U��Y�ٴ��H�Ղ���^A��9�X�G<����o�u�Ȇl���6�k�C�Q��uDV�l؂�2cJ�X�:���8@ry͢�~a�|��*9��$�U�c[���+�4�̹4h�k����G�<"�ձ�2��r��IT��|�<8��,��3�͢���
ƍQ��A���r�;�8>E&���Jy�l�[h�/<�p�:��y���w �Ph�v��˜3bЛr��9�rhՋ4�.A�:�����AF�����pN!�՜�`xç�'�gj��r��p���x�'�r�X�&���h(63��$4���h
9:(i����C��CA����E�j9�3��9PX,�4ɤ�i(��U�p�4�4���TY���	��$ZLT�$ccl4R�r�E)EU'EPQ�,T5H_s���劌m�O�9y!�ȡ�:���.X��N����������6H�Z
Zh(�&�)#�̍!�+J\����QLEPh!����M��Z"Z�������nmJ\�Ss"���`hj��(�*�f��ъ���i14�TQF�)�5̅HPLQAJ�c�R𑪦�(o>χ��^�VU(��(��e����'(�X�=i��\��3wܪ��2��R�2n����P)Y�az�K��a�I�U�w����|�pG��w H���e�� �t�%J�K��Q4�!|D�)�h��.��y���<�>� $��߯=�tY����K\�����j�fY� �����<����2*�����?WyMڰFۙьEk�(���'aB�w��5Ɇ�a/L}4o=40���zOނ��	8Pƥ�Dm*�X���:e������+�x�T�0ld2}���A��b"��v���c�q}]�@�����(~�O���^���rfm8���)����o^kè�/�8	�VK67H;�<���h�<�V�~�muMUj˅SpX�v��p����d��`J߱�_�K�o�'}tW�����!��X=��N�T�qK�[c!��;b2:B���N����(�ms��=��g�7��j���v���S{.:��4R�KO]������[P���36j��zx7K�.��'Tۻ�~����;.$T���-P��̽I�Ȫ[/�
�nb����e�e>�BќO��D�@c
`$^���/���U�n<�y�9�=
�nKz<5PQ��oe��t�ĺe�i�[�TW1���[ΫY�i�;8�c�Rӵ$LD~�*�K��~��|���xjC�W���[t�v�妢	�)�:q��^��e#:-��ZX���Nt
R-����>�ޯ{��'����t�"��G4���-Q�Kkd��V7|�?{�ͨ�����jVe��ռ�0��́�.�9�DR��C.a��V��7:1:ں��G`C	�34��M���53�׿�{�|����}� (DT�U��F��y"��=���9H�w^+�j�F�+ke��Kc��_�s�� ��5h�7<Z0��/�8Lb�f[|����{�N�QM���Ɨ]�=9�	�RSz��afE�=�0Ku���������t^m��fCE��ø��4'n�-�]\ܝc�l #ZDdQp��ZD�P�s�S���SG@]�b�E�A7Cا��x���Ξ���TXXK��,�[�V����w^'�4e̜���g�L-vval���'-Bg�7]@�1�a�G�(��=@G�_c�s�.^��b!�>���+NJ�˚���;��7�X32}/���П�#c�פ�꜖�JR֙��&�)�.ʅ�Q�m���`^.�E�6�T{�FƤ� >����I�y�=�)�S�m�:n�t���N��EIhש��=�S��c2��5N��Q��I����v��6^�n�,��əZ�4�l��,�M���,��>�y����뚺.Z7��������f��h÷AEwVm�s?3B��v�O�m�ӛ-TP��|�pι�zc��(��)�>{��o?���KVA��,�G�ˁ�$��YT_1Gwղ�xOT�Qy�=�uv���+d��u���Q]�TL<%�;s�〯�v�v��b�~�G:h]�Ӛ1���)�WY�Wo8������M"%�v��-���P�gyr�+v[y��=Y3A��,]]�_(O>հq�> ~���""P���- ,� R+>|����������޻�w~���clj�Do~U��tG�U-��U%n��sz�Ӡ�P��tsT+hvz	��u�ov�s֊&���e�N��&�LJ�lX����pZ���ո��Z��!6���Mf_As��~�'q�z��]���h�ˬ΄���0��*����yT�u<��-�e�i�ԎI�ҋ 98�i���i��ֻ���Y��;�h�D�MQ	�4�>�R2o��."�ڸ���vd'BvM�����+�2ۮgņ��n�c
�B���f|����l�U%G��sqV�E1Fl;`�*��@��#eW����O18+����sS�m��S����Ub�br�}����ϭL���Ʋ�>	�;�<�����<��;'�}b0X������(؈O%a�׍�F\��y="�@�3�}i�v�3�%�mO7�_w=�w*(�t�Ⱦݾ]u7�Vɋ� u٭�=y�,'.��3̵�7?��L�6�� ����b`�f,ه;�װ�e��3��������+Z��K��;CG��!�s��`3�����cM��ߑ��+}�`�9�X���5J���C@<���ƝJ#�驌^u��H��(����S5���t���:�@��8�-�����hHec玏Y`�;5��n2��S�FI��a�[y��,���B�W:Jd�r��?����TO�% "S@@*D��J#@��P��o0���zL�x.^�U=��	o�.��<�����ꇕ��-��݃��kt��B=�D}8D����P����u���3:�c�y��fi�%>w<{-�>��]_���C�P����9h�Orʑ�V(Ԉ�o�K�� �獖*�Lg>3c��#{��#����9����=3\�6�f��H�dD�mR�9�
CCx .!۱��7��SCB�M���P͇m�ݠ��=]�a.�(y�Ƣ.��f�2���E�#�ԟ���߾�Y�2׌�,� ��4�*9=zj1�,d��fd�h�ة���=Q���+p�h��06 T�5���J~+
&�x�C5�cN�FEC��56��y�K;[���|g#T,a�V�ǯL7<H���ג�e[n�;�I*�i�W�|{� ���N�Z����bi��Z�t�Bڡ�7�z�]xm�0�[�ɺ�K&��ݱ�-�j����3� fɄ��jc)s�͕Fq�5��dc�����6�^&������	�N�樤�x�Sm�1�vә����k%�5K����4?�E5�J]��e>���8��3ԋ�zNK�<ޟD�n$!	5.iU�=���s�(P�}�'���ٵ˅��&�v�7떶�͡-"�J8�]�P8�$�2~H+����~Y����׿x`��d�5��� M��6�ٛ�x1=`���6v݌eh!ᣮI�Z���.6�s��*%�{����)B���4-(J��P4 �	��
СA��*1!G��o0�0��F��튋�˶���O'S2!RA�p<�`&�#�̗q������ F?k��F0���鎆O�pY��gk��J�Y�nP܋HD���w��� b�y�R~���{�[^���!�q�d=F@�gE�K�b�o��r#$���D]�w8�0��쫕��Z��'��P<WE��m�r��0��g��l��x%�jv���KU,��*k��o4R�~�*D��(�\ۀN\�����[��z��|h����wm�Dh`fS�Z~n�y�st�x�`֞h1�t�%�ޑU�W0��О�͟E����|g}k%��C� �؜��GIs҈�h�l%��1-�{:tc��E� ���N��E4��
_�zګպ��եv]���2�^�F:�`š�l�ݩ�O5Hu��=���9��h�������(�m����q��
v�ev�}z+_��	��ޔ���jh�:T����tY��Htܫ�,�O���H����6Q�7�v33���К�/���e��G6tE�'�^]���k�|�
5��i�WZ���n��;��A�Z��팬�v�-�w��[����i�����=Yq�y�A,����lv�v��h+����52��� �a]+˫<��l��<NF=�� �]8�(��R�4;5̮��$����;�^ޛ�x��Ġo�<a�c��-�lS:����i�]sn�Q��ԝ*�4��!��v�?||�^����}�A)H"A��
Eh"�d � �X�BeJA)Q�@oGY�37TQ�ܒ��z��w��I�i���6��Y��)5�Q&3�\��r�e_'g@����-�����ؙt��m�n2\���S	�V��Cը���Ȝu5f�f�Y��Nmi��ϐ�)�G&!�ۘe7 c>T'@/5�i
9<���5�&XRml�����n�Ѯжi�eJ�t�de/�(^�][��v5mC�vկހ6��P�!�$[�4R�n`;��f�U�����8��vF��âg��%#���z��Y�6�[[/X��)�#$O�h}���ȿ��TSK�}�p�,/4����tx3F�<^Ù�N�̢����S�"�e��=9\Ϝw�����;�A{�}[���-cK{Yz_�-z[ _t��<&��ܟ��e��KP������Xg/o.����Vjlmڷ>�4��mx4�sy�^mt���q�����\���e��@-��f�t�fvm��~.`u��j�s��w�-�0���x��P�*zcx����TF�eV?=]\�R���u:�ưC��	��,�;Ί��@�Pżo�mo��e�Y<������f*a�NT'.���֋��Z����H�����y�Av\�����#=91���%e熑�]+ؤ�z�p�vqK��0�?�ggl�}�(s{(�K�ا���L�7�8�;��t�ݡɮ�o[,.�Onn�)�q����߼ ��7�� 
ĢP$�%D� TT�@�@�H$ʅ 1(ҭ@�O�y����w,��pᲷ�~;*2(�Z �UT��|�^7����@�?��i_�Ԩh�M�/dȑ�.�:6tn��miSʵ�9p2S�tAz�wIm��=3�C����y��e�!��sw̃t(rwz�����]��	�H��֧0;\�8�g����\��'�T�z[K�=?7��ʇC��dY����^�Y# �鬞�-r�̄�@Wo�N/��=�ŵ�zm�7����z��CtՕ�������	y~�4|{�K�=Zd4)��N���W���ݪhj܎n���mogBS�\	`[`U+%��0�*�����^˖��A�5�����QU{�\-�Z�/�U5������}����V�?��4Q��Q�X�5kH�ŕ�p)�X���� �f�m����h���|b=�':���Bv������+�x߄^9{}\�7�{z�Zk���M�S15F���3�H�T�1�Y���צm�6^�M#��b9��fS-�`J�?aSlhZǂ���j�������!��yJך���Xח ;Z�	��c�h�d<����;�t�����U���og����������j:�̈S��Sywg���zq�Y�Q���|��q�HQ����\��G�Ne��� w��C=�G�f�j&��_�~'�Z��@�Qa�[]�y��a�Y���ʈŅᆭnw�(��i���̮\`�|��vØD>����������oooy)�h$@�F� Vj��	!i�&"A�"@I�I������}y�������C0����R�mj�����/�CϯOZ��ԧ�ߝEs�Me�Φ4V�jxU�J���]���:K#Ec���q��DǝR����{�RZsnF��v�V�-�֪�z�i'H�</#�-���3�ǶgZ㡜��!6�v�bޓ���dҬF	�%�KS�4�\t.�,V�U��-l�k��3灡��A�p�^�{��d�� �sm�]r�	yd�R����>������T��[�1�!s\�u�.�϶0��<CU��{��]W��S��M��\5fڊ�l�z���C2�[{�+hȍ���O�\�9`8�9���"(����Gu��`9��^ s	��0���l�k~>:��:�����w��CC���(�8#���W�vxȬ5
q˽�,���Y>^jh�M->Y>v��Ec�f���y����,%��0q����gd8�sH����<#r'K�O�a�lA(G@�����A���|j��m���b^�#'�,&��n^ӴW��h,�_u�l���\1�	��'8�/������7f���3{jz\.\4�f��e_h��'��"�з�g0ւzhYҬ|i�t2�J�ٿ�Π�F44�s��Y�^���7���~";�K�gjꑽ�}�Ps�p��rC rؖT��|����{nnr�8���'�ן;�?>�����h�ZP�AI!�a��P�h�������	d�ZQ�@�hb���]�7~�[v����d����gu�:����A��"߇�z)����ׯT2x�	��sM��]��Qq%z.�8��n�x�e{'-Y�qB.E5����.jB�Q+^������M��U0~嵭w�mˁv���}�ٸl���k	��exғ�&ch�<[D�d6�&Ȉ�3��\{N����«<����=��hSf.æ�>���&_5ݕhh�覶��m���8���)����z�su-}�iP�i���67i=a�$41`��w@�T�׌5�wl���oVS�0���鎆O�z�	�s�D.���k�����ӺG�~(�y�ܢã _9:�w<�YCfz�Cg��xޡ����}��'��!��yޝ]4�-��b�nCa1�KS x˴�3�^&�s�������9 ����>��]l��׳����+V��	R]K�~W�)�����ɇ��)�=��y��@�`N[�$[���@M/=W6���K� ����J���e���<�o9hk����{�M�tZ�b{�TKo]a̅ٱ�����P�� �~m�:(�E'�#zF�c����]C�z��K�~����Ѧa��a��Gk�D��x8�])<���*%�E��6���V֭�^:}��\�;,�&�z���y�p��gEV�TP�Z��x[�l9�_q��(�Fhy��ݦ4���u���l�W��ɪ�+��5��>:�ˁ*��D�<;fi�ݪ��/�����Ȍ��Ģ��P�D R�B�H)2-
��9ڮ�d�B'����04'��(p_�(4�!џ��ӣ�_�WӤ�X9��C�|OoKw�	,'7�o!��$���֛b'KiL聆�7��0�'��w��)���J���!��'br��ԗ��̡�R�}^�=@�<|�� K
ޘᤠ�p95�]��x��9�赛,*z���{q���D�`7���47e��;��氝3k���<�����u�1��kk.ӛ�n�W���i ��<������xi��{ٖ�٫�yU�˃m Sz|%��M��1˕M��v�t���k��H���8|��V�Um)�*�Mt&�z�g5ܺ�{0�0�֞�.��.o�n)������L�]�|gڲ�7ֈ�]�5�ɋ�����֎�W�a���{�֩�lRz"b]k^:�f���e��[�.ƪۖ�^צ��ލ�j��ċ~f��vK����j�8n|o1���7�!O5tL�~J�������bٵ�ޛ0;�V[問߰ k��
�a2U�<u�A��t�� �:ak��*7E1���S�4�챶�j3���n|��s����?g��~ϧ����x�}��o������x����W����z��;4�÷uy�٩�5�Ϳ�\�R;�V��e5Z�/�HC�F͋$�x��������bܺ�l%	��|L6�_�q�a�:�������BWd.�����Oq��M��]�����]�5��������A��C,��m̌��J��Z�WSwh��6sP��Fd|]���M9�r�egAd	�g3&�7�̤��!���ڼ�0��X��$�v:n槌X:��ҥhɶ�	�&=�V��Z�����spFE�'A�M��I�)t���7��B\�V�'�b�.��,�B7��0p�3y�3{
=�]�|�x���J_���h��.�Ws�1��U�/;eEXj���w2�vV\�{K����:�LY֬VCHǺ��e"�v1�3i�[���\.N��w��u9�lp������K�rp��6�63F���rR�]p���
�kF._^� �M�1��EbZ�.�m�&�L�&Q��][�LN�G�]�7�	ד�����$�����wWcy2M]�t�79�B�}0��]br<��<Fr�j��흂_�$������6<з!���SX}�8gt%��paP�sw��O���703�ֆ�V]�|T��r�)i��ѵK�ݏC+�U젻*:��dJ�}�u���}��&]m]="IX�,*v��2	����9����t�N�� �iS3�`�β_^|���W7���\b0,�Zd�+��#\']����m(2������t�A�ֶWK�;X/{2s�vU�q�T�QTM�q1����n����6��%ɚ��;��1q�����["��Q�R�[�N���kB���ُh@*l\���)�J�[�%���^VJ�z8���t���U�V�K8��O+��fA-�ʲ��ɍ�����j���Q�޲i:ܵ��@w���p�s9�&)�V/C
h_B��q���hN�Y�Ah�5m)�)�V`���C ��s;�t�|g �͠rս�&]�R=���S���m��LI�/i[�5�7��$�T����DY�;��
f��n���o�N����[��~�gOJ������n궠��������F91J-��#Y;��t,ɮ��J�x ����<6ⶤCh̕n��̥�C��4�˪f�3�uf��T8���ͧ�G��7Cm��V�;Q�k9ݕ.ҭ�D� c]�Mgv��yr����먔�L��2������ݗ�a�n��N�ok����c��q�-X'r�R�m7f��k�vH����(7r�jy"�Υ[��
��DWv�+6n<Vu-v�Fjg��]����줃��6��W��Ā=}�WX�'�[Ƹ������`to�
j��ú�T
B�Q��)�X�7
�#л�:�ۮכ]�9iG���׽�	��U��6)�(�v���K�c\T�*ֽ��n�+�BN�oH�%~����W�@)4h* j��4�)O+j
�j�h��
�M	B��iqihi�H����&�>9ƃ͝!���.���������t�	'A�#JSEyj�(h�h*���4PL;�����щ�@�HV���J�(�i�Hj��֖f&������A#@P�[b���c
i��h��Hj�&�5�ii�:�� *��)ZR���U%i4P�1%4�-	E��M.�����h(�
���h*��JѪ����ţUE�;j4h�����CB4�F�C�Q3F�o\�Q�44�b$��K��6��j�6��B8��j��(i6�@bHD�$Q4�UD�@V�TT�MQHL�C��ֵT#�����AHPS�����$�tcT-1i5LMM,M옒j�� j���g?�������$5B��Q���>ƈ�ۓ�/Lp4đ�P��t��;҃�
��)��t=���j�fԴ�����eEӺ_T�N���xi�Ba&)IB�iV!V$D�f y����n�1|=�[�>1���|��>z�u��֘X0��۪��p9�-<����V�)w=Fn��M���w�Y^.�8yɿq.[�i�j1�{a� �z�_R�FK���]��UQ94oa�";�%�c�<s�ř� ��dg4C�����ަG��\�âq�»��9��/���t��:8Ġ`V���Iv�^�9a�w��$�C�~�TS'Z�ڌ��^�h6J��kp��a},<�t����Tcׂ�-��2�Ǟ�9���m���G@x�	�M!����+�Ѯr=
���L�ԩ֟93�����{��iw�~�'V�>T��4��l��[ǯ
|��B�335W���K~|aB�������rG<�z�1��O7=@sơ<���C�țu�v�œ�8=�}ʙG��:�~w��}�M�-T��v/}���g����uК�Lm��:�c��X���\�(o�GO]$Ʊ�?�������E��ηv�!{'����`;�Fڜ�N�K��$�z�)�g���X�w�Ч�=e1({�[�k��Ǽ~_������$п֗���u��wo��6t�+����Q��_� o���v:�+3;�N㓸YƘ���o0�x���zJu���C�M�3�S
a��[N9�omt�3�xmu+hte���O��A�^p���u���s����>=�o������Y��()T���
Q=s��s�_o���ޅ�X�xIh���A1�r'U�	�s��L 0��p4k��ڙ�߄�-��pэ�0Y�@fד ��j��sc!�]=V��R�-]i�Ě'��bj�0h�Q�3���T� b�3���M�44_l�@�O7�2�	U2�����6��6�9E�����OV�l�v��H��#�Bܴ~YN�tx�����"���=�����'<�[�0��c-���ԝ�D�����te�	S�����{��|i�m`2H��&�_t��i�\���*��Ҟ7��^r�*4�eZ�:�c���8�[�E�k��Ͱ����k��7�����2�m����Ա�3xB$�O~uλH7��576��#<mښ�����i.�/&X��vB���dN�Q�MB���8�֗L1�d��8���Z�ۆ0d����a�,T�u���.�qDr��c���ɟ];�j�O��n�YB��ֺ)��b�@��P�b��p�M]U��T��Jz�s1S`s��F�Қ��j�9���s�}���gLO��?��(�,�iꦸ���������a^W�~����'oS7QA/����Zn�7��}�a��
���R՘#ĜR�a��@P]L�,,3݃q��avK��3�c"�[ٌsh�̶2��7�{�!|�_.�T�^��P��:��P�w�s>�|��>��~�M�%(Ġ�1*3"� �AH������:x�zz���6��rҒ�An�7�&��D<Zk~o�;'Sͱ�������@�
7^�1�}��$�c�8�,}���˸�4�֊x�����q����Tŧ��N��"'��!�����B��-���o��iޭ�����Sr�%�;#a�������'��p�:n�=�����#�x��ދoJ(SI��E��T�+nZש�<��M3B��<zX6��C��O�6M�f.�f; ���;�%%�6V~��ɲ�����k�Jh`�ۆk�j>W)�mzJ��j�v���jb��^�'6��@�z���+�:u�2�i�,
��&�Q+\�t4҉nl�;�����ִm���u^6!�;T�;���C� 1�-���6�c{=iݮ�����	�3dt�r���'E��A�;�f��
�K�l3|/�o����{kF�+Y��tl��=0�~�.ў�!��ku\[���M��YM��ClD@fލtz-?v�g�q�{^}�s����˯4c�M>��d�W�9�yk54�3�tI�/�g8؜P���u&d�r�O%�T;��im
�>f��/��b1�KE��o_�����_U;���3�l�OO�k�ח��J�jP@]aY ���;Ã��}���u���|�6�N�;#�����S�ݍS��zĭg�˔r�C�z����+m4�t{��.r�.\�yM�8-�Z�]<� }kσy������444�x�ڛ�Nق��̨1o�^4��v��n�_�(�]5��.�޹p]����b�{��&�.�wK�s�A�HKƗ��~�"Kϭ@���&�`�Pԟ�t�-���HZ�m���ٜ���w�;W����H]�z`��d��tǃ��0ӯ`Ft��*�����?,����y.�VЯv�͜o(n;L��͏a�ن>���<��Շ�NU�}�[��|�|``ZM�Ѿ�H��k����rJ��s�9��� �K��S�}
Q�>ķ]��vv�{��Y5��5HS �ٰsÝN㽁�XoD<��,L��E7���x���<�ŗ��y��L���[��f`��g2]����h*q��q7� 3Kfޘе�C�X`����v'��z�\^j��m�[���	��d�����!���|�/Х����ֿ"٧�ӳ����#pa���oV���W�:d!�X���R�H�e<~H�������dTk�k��xU4b�¶�e�"O�u�P�h鼤��~�t�%=dpm��s�{S�V�A�8����}�����)���m��� '�{���_�=џ�w��%:�����b��`,Σ��;��C�"���-�t@�Q�[YIEa-UY��+��v�n��h�a���I��V�Vu-��t;ᔥ�_ׂh����)�|U7�,S��D�G��3����u��W���~ҫJ�P4z������{��߷�_�fh�{x�Op)��j�!�j�w��c�}����of�P_�-���SC"c����L+p`Tlm��O�vSMv�"�jچy��E��� ��C�go4.�1¸p����}�i՚���l�M�%����9O��T+E��emF�6�� ����aU����_1��1Қ��w-i�ЗA��\�o�?�N���i��ԧ�"��bzs&7���*n�f�tnpN�N�x�iX��g�ļ��y�!��Ra�0����e���W(1=����혍��
cCH� V=y�:�Y�v�c�C'����uΎ��G���o0��-Y��N�Һ�����s�v847[�6k ��q����Z��r~��N0��E?In��wm�^��;QX)q�xi����O^Y��Jy��k\�{X�r�0k9`�����3��g�m=���(c7��(S��K�X�Q�qK ��*�mj�h�9�1�����z��w����'t��˱�puZ�[;*J��~�;��KF�t�0�N�v~p���!�6d�����m��)C�|��wd��-��HU1�2Q���A����'�[�-ײ���B�	"*5�.X��������QA�xQI�AS�/9u�r�����P�ˎ�L�s�R�^�u)G/���c�]�騂�6�tj>��"��U(�����~.z������}y�=z]����m�P��~����3��|�f�W\жZ9�3�\�O[�zsb9x��5�y���WC;�֖�U�����UH�g4�:K6��y,4�C���E��	`�(-�!���fn�3�G0�|�T�_d^>1�ٖ��iN$�/�g����Z-sl��� �m����E�~�B�W4D�(J�lm(����!�S1��Fݽ^,�1��7��t��{�O4V)	�*��M�j֟
�YQq�Z�������S�uv#���2x��B����\N�.��3�>ǿ����BÕ�#�~ޏU����a��7�͵�5�ԤL��f��ܒð�(H#d�e��85���f'�W��L�%T�yB�j{��x���B�c9���uv4]^�n䌒y�;u[��-�إ�Ƞ�;I���!��*�����L,%S�Kh��3����o���-�����|��0g�At x�V�XpBcC &����J���f��R3M���4a�J�t���.�`�������x�����!�>��mṽ^>Zɴ�B�~�c��X;3@�E:�:}����j��"�ڻ����U���I]C��`��]��x܁���:5�9[��ɞb�[�$#L�C��7�cꈎ�r�Bbzd�F@\)'r�լ����8U�]�R�'�����W;��=�8k�j޳F�̣�? ?0���0  ��;�n-;sU�|w	&ndU40�x`��T������cȏ˕��Q����%���H�.�1�P�\uK�a*k�ˮ���ۂ�Z��]�u�Cn�S,�Ԧ��g���l(���-�O�Bֹv��N��heQ�m�'7�o�dY��y�z��X4b[Fj�NQ�h�+��!t�O�5˷MN��eƿuk����d�0�1i@Dh|����3AkJ����k�ߴ��ǲ޻�����kyNn�����'����x��A�ht�C���ͣ��T>�@�!Fsױ��qz�wH�-S׸�ϯ�e�	�(�Wt�8񡣢/���L`ha<��>���r����f��+���#s��f͝�g�q���Z�fBN�nہ��(H"@�6�?EMʈ�yw֐�w�9�J��ݽ�p� /���\��-M����̗i��c����<V� �(/_P�9��{J&�1v�;ru*�J#��Cݮ<LY�C>�Z�.
x��U��>�W�/=����mO3'����Y.�qE�Gm�s��6��ݙ+8�8�	�<���w&�{�B�;m�j��Sd�R�Z��d��Q,�o�eM>�����S�،p�Ahmwǉn)-��@��KM�U�[��8����ה����<E��:<����uc��ʝ�mM�Ah-*�mCG��AT�뇧�q�Fj�)Gt�]��[��80�S�1[a���P���9�a5��U}UU�r�����w�Z�];"��t3cf6\�w2��a@Mx�ax�z�1I�rL��ȡ�����:�Ͳ4�R)��a*�{k峲����G��"�ڡ)f�4Z�a/{
Rgk��/��mL^n�;+��u*���9E���T,ի,��٭>b��bM<�e�h�SG�����)����xP��B`�l}��v�YC7<��-�Mc�.Q^uϻ�P�z����lRʆ��4F8��j�W�R�S���%�_�&�xd�"�ӵiS�P��j��]!����g�3��U��v�K.|��RT�LӐ0��/^��s�����E3�0a���iO��̱?O��w��gT_]v�*��rY�@~f��H�m�c�`L(<�%��z�u�B�Q�,�k:y�����h�V.N</D����-��O�먀�\
���t�l�|������x�fStm?cO^����R%ŭ�C��"5Lξ o�CO=�nhwf�3I	�th^�=GX�[����uD�G[t�{ejƗ�[�6�.���l3�f��xŉ�s�0�۲%�!���>_����?���4^��_�=ZDX�g6�NTn���B�Ԗ���1]Nr�vkI���G;�^���Yr��Zk�j[3^�:� 0��|��w,��7��Γ���_APk�5.����Gx��Ө�2�����+��a{����N��{��:��}�P�m�me�v� i��<�\Y�4�殈��yw��t���[�b�v�cY�O��7�k�e�f07������ps����.�ɋV�R���'���O cͽ^o��^:O���-������^�����8�N.i���ގ��%�m�����6'4yy���z:�����^��S	ĥk��HMɂ���\���rko������Ek�{(V�U�)�\D>P�4ce3�?���H
9=��jv�	��U^�m;��T<k[v�n.�E?��t/O��8�������Pk��z7�q�+��gF'331�ʼ6�8^.����klB��J�����hV�ҽ��l�YY�Pdny��h�E�]Uu�;�C7%��n7��њ���9oL�u���q~��ί����cSU���G� )�n��M�A�W&�|?sץ�1/@c�y�����L'��1O���]t��tewn�u�U��kR]'\TrZ��	��r��ь3��9�]����W��=�9d�3Jh}f���f��EO��< �xp@�K�齿Jshށw��SM��׶�x<o�b��D�w��K��W���L{�tqXgO�����v�w]�\FL���^��2��k+�Y���P� p"B�*mfˏ�$�M�*M�?�  ��o{;L�V��>(�7u3��nd�^�d%�a�C�%���z���`���x
m�z���~j(R�g+�ptƧV��-��-j����K8�1kgfO����Gus�I���Oϋ��aJoO��+�t\r�-�e���z�:��c��q����`��e�ڳh�����\&���1n��E��v�����:����������!����DaY�D�'5�3Yt!�^L��S��K�}au(�۟�F�U�=�i�x�I����,c�����"}/�~+,���?i?J|��:+K&hU�}r��CU9��3I³��v�a�7��0��񓕌�hkB��+�m�gE4'0D�ϛ#�L>%�J�+��.���8�p�t��2��N÷v[�YK���
'(j�w<�Ҝ4d9���x�4u�V8�v܈�7�{y��ևE5�g���4J�[��D��c@��*!����]��S}"*���El��Z��C�Ou�M�דQm��d��.�e�6q����V��0��3�=��_�������������|||||}^>>>O������ D��a�ށ%����!��wu�9
C�|�٧����tF����b�SN�2�e퍾j��KJ��nA�Q�u°7bՋ�Aiwr�"��+i�}z�+S�sdd"�c�X۳�׭����|>�V`�i4���eh�������ge�\�{](�+G3��N@�u]�h��·L�u�O3�:4 &�1T\���dr�/5'�\�s2�<�G;��gE�n�37 ��r$�;��r/�&���v�]�^��:f��3� �)n_��tu3ft�НHZ����q���f�e�,���gK;��+����і�-�	����7����vUd���S�*�����(���N�J�Į�.�wv����ҷz���R�a�0��L[���a�{`��S�[r
9�V�Ed�0T��6el���VVqF>Gc�7�s}����Q������;����D��+���%�=��;��ju@n�G�{����Ǚ,NT_>��U�;v����ڌ�o+jf֔x���p!ǅ��gF��4��q@6�j��:�*Uy�n�P6��|AЍ��� �5�X�ef��F�W*�\����.r,�3:�
��EL��B4�7E�ݖ�vq�#�yhC�R�ܘ��ut��߭r=����,Oh�n�V�f���*�&)�k��)�J3�Ư���R��T���2&&�֗��Z]i�A�G��y�|��6��S�}�8&ʴ��c��U�p
bNY��Y�\!��:A�+�˝J���RD޺"�mh���Z&e'���"?+�q}���GD���E��w{�Mz;��w���S�R���m�' �G1Cή��K�� ��Eݷ�"�1˥x��Ϋ,'y|���}[�#>��x9ݽ�Ea�
3��,�k�P$Awcd��]>��fК�-�c/�4��F0`�� �H
�&���N"�^����Nר�s��vm)72Z?jN�4���6e����ݖ6<�w�r���Rg��,h����7�6I���R��Y�s:Fe�I؞�����ML���l�.�WAKi�Z{����:٤^vT5��Eu+(kt�]Ga� :q�MqWZ�� -��ڨ��H�+k�yTֺ��ծs�:�;�0}��!�a�?vNns̭�.��o�f���ۭ����%uB�`�\3�����eVN���JF��t;��8����c/��&a2��A��͛���ﳭ�����m�r�&-q�����|��9P_rch;�6��4�w<Q��2	�A]�x����j�-6:+����.f;�wZ/�KL�\�شaL���ҟ>��₲�]F��Bn�4�w�'��n+}\^B�rs������>����]l��/�]���p6N0.�99��F�v_pp%�YK�]��1��{�k������A��-��K}b��@Lqn]�҈��E\lڨ�pl�\�����}�H(\軧v��]����]�Lޔ�H���B��@�� �"
D�h)h)

bH�)&�v4�iK�I�R�i�j�h*���+IF�ER�)q|�G-&�E4�%- PҥQPPS2�IF�E4���)KT�1D�4�RP�4h����
�h��hR��AA�)�h)��i(�(�`ib���R�P��-��DS�ئ���)((*��)�(����)�Ө�*R*
����&���O6Nl؂

)��"J*a���%1�V��E$�F��LKIEj)i(���٠��B�Ѧ*kK�65R�M%SUE5L�i5IEUDM4U��mjCl4�P}͐��!�

��b���!�����*b*�6<z�>���N�(����m|P��%R��J ���6�e�a���J�z	*�]W�r���Y�^�|��I��:��cj������P�W6�.�o5ϳ�uv�p�&JT�tiI	I|�4�B�5D"I�Sa�T�k���;c��9��n�y�
��9�&.%[FL)���	s��?�`�-�,��86w��뇎a$̦@v��s�����`����l���oLS��`�����ThwƁ���(LȾ7�W�A�\����07r�`򅭍��o���&ڕ�r��������GV{]����ᩞ �/|j�!1���/�C�"뫞��CfE��{h���<�I�7�K�hFm�k��P:`���3Ǻb!>�zL6��s
��p��z!��L��t/�[�|��A�%=y���� ���c����/d8��9�u�+9�Ή�[�qqU0Q�zb��-Met����QiG7���|��]���ͧ�9vg騠�N+Ÿf��=t���
xhN�%嵟KX�S��#<єW��|�u���	Ӂ�=if���eD3:v(`źDmz�����a�y�4���`����[�BƦ�pxK��zM�8�ٵ��3+�+̩���8;k���m�1�����9��)gl����]�[Y۵��b�-b��"�޻�:f��������|{p�T7��B�E�٬� w��������
�v�L�C��J!����VzU�X2�]�SeO�(T=��p����t���i�fv�`�0
H������mS�]B��7����+i�	�uoF��@�{�ioU!Vr�I�:�Ձ{���+�}�̀�Z�����\V��T�Cy���}�}�º��;�:|+�c�a�AY��o�6����<X��O�a�lA.*�..��Dj�-�7ESzv�#���[r�|[3!�t��G�\�?��cV�i%]Br��3%W�u�b�݂C0����4�1���yU\����{����&b���R��Cuh���/s��U+���<����Q5�y�QC�&I��������T��[՘A�P�ɷs_4�|��>�>�s��|ZNLҦ���Z�zga��2��;�<��@Du;��	�_&��6:�Uس�6M(�mBjШ���=�g
*+��@���n�6�����?��S[Tr�m�!��	������N���X6���p`�k����T�;j���u���>��C\o�^�ݱ6E���]���iL_�� Z���4�\����_�E_�60.]�	�@%\�i;�+n��f��UʭqHK��� ɲ�4��X��*q�w\��{G��5��v��!��A�j�*b3/�C�6��O�G/A~q͕by�+��#(���wle�dɮ�KT'��9��i���n��֍$��+��kj�e��I�^u9�r�LRmJm��G��i]�S��r�[a'��x���·�L��>�P�<�U�+iwCt6���a��yu�p���u�竒;�Ǵ��/���� �H��7Z�_os�S���	|��F27~ x����в�{�I������#=:\�a0���^K�{���#zEW�J�`P�'�4SaȈ�;�k,w6ۣ�>������r�l��pq���@��X>�|/�k������M�5*����a�'��1�I����1��ےVVk�қHa����D��/=�|���w��Տ�����GJ��C�mG��tI�z�a�:f��=�2��'|<�����+�8j�����!�b�mу���vD��*��xj�'��Jߟ�~���~;Wچ��J����Ib����.�f��<GE��^f����X_s��l��Q��|�]�^��hM�pGS�f𵽆��E�CB����=�B�&*����3p��ǎ��gMcX�!�\���6'�a��VK��Yx=�/�ӝ1/��p���|����}�ٟ��4��S\��KLT��d���▮�׉��ڜ�b��f)>�X�\�r��/WT;��ڠ��b���>��-Oj-)6ƥfxkx<Lmd�ި,�]��ɢ���.z����y�B���n������	�k��a����A��]�ܶw-�"�S�(�2+��`�)}o��RH�5"y�����w�ʷ��ɾ���E��j����|�l&���䂧t�<�E`���F�}:C�( ԃ�ÇN�t�ya�7:N�E���m�]�49�c:ust�������S�Yy{,?�/'/�H�̖ϭ�����5�M�2h�x��R�v�3�/~̹^++���rx�s�tcsOFO��9�WK�ЗC���_8f�Q��9���E78��䚐C��uin�b.���1�0c��Ѐ���"���ļ��zо�L+��7'�����3{�v6Zs<�([���츿DF;P���B`&<��^�@���J��WL��5�j�p��}\����K������_]� w��cͮ[t&�u������Z!^no^�]�)z�u]6��5	�� �ƴ��Jֹ})�����[p0]�8�k��8����ػm�EU�h���4�,~�_7�I�cq(����NY�L�c z��4�Q~fG\�ͭhM�uܣ����W!���9k7�:"�ZApk��u�5��ϯ"z��9XY��&�&�v�؆p��ܨ�@�g��&�����觐(:�)֟9���e�_3�E0V�Řdu�m	ʜ]�ra	fXn���{)���K9uQ1��"$H9�+�k'�ߵ�\@��v �O���̻�d����Z7��K$o%oR��_`��\��шe�n��g�S�N����'*D{7������Cx����4XwF�w)pR�^���o��N!&Gٿj�r���Q!�M,��3(WC�χs�N�$b���'d����S���}_W���-��ݫ���I��+�	�d�
��5�����3��,�����sg�qr)�<Yz���hF�\�b�h݈����DP�G#T!���F����n��r�W�'(j�w ��a �;t�Kd����!g�q�}�՝G�k]���j�QM�3�ScX�BSB�4��ҙQ��h����AL�&�ܳ�ѮFvp�Me�5�2-�C�O|����'��S�D�d���X���b��p�����{��륔�.	��EC|LɆ&�/� �κ�X��Q%R^7�7�9�w�ŏ���es_�`�����u0�m�P�dLȽ~�d=��u#1���V��K<Ady�T�m��i��:��k��s�j�{c��.ŶxF1���)M�TFq{�塻I��7���I8�T�O�:��-h�cC��rМt>��[A�=�"!>��ս�S&<��/=�T�-3���S��\ޡ��B(TSۨ�tsΤ��c�s�w�� 4����;�d��0&ѽsWW!l8�%�;�>v9S-��������C&�4%��#��Bֹv��y��Kn![s<M��x����5������Dt���MuN7]��J�`�Z���9���6B����9J���W_8�q-Y��lr�p]�f�]/�΍"�N���Ӌ�^r�xN����"��0^B<�N]����f5�Iq���\l����ઔ��C�^�_��cA��̚���1��Aez��ĴA�llCi��]�zn2���K�mn؁�zC�l.xf/��Ҝ��dCN����j��Z���K9�'�.헣i2#k�k�\�9���������a"s������P�lt��pb2T#u;�zm
mj�1~�ĺ�s��������]i�3�%|sCB�挦.���s�ݭZ��B�k�%"�w��El��[4�9E#���)��%�5��ˎ�57c���1Yxe5^���e���|�}�R�>�*���)��z��jX�~h��.�fc�ľ�_
�W�yyH��#��]��xӲ"�����6��%5��,�+ܥ3k�wL!Qѧ�A-s��%�7
��t���X�LX��xa+�߂����5 �P�Z����'���xʩ�Yx�������M�mk^��xm��mQ"��7\�w���a@M��쎀��kg|�R�.���5��Ew?�9�����:y^2��bফr:P���yk��߉������O;�^��ɟ����{���A6��v���zCY��N�[��'����]���.�rp���yjן)�޽��m5gY�X��G- h�ʉ���xm�O�Bc]}�	a�m
T�WU㷠6�hx�}��>J� �s�Ut�h��VM���}Y=={��f ��F��Q��|�*�|���`�B�Z�a�]�1����ƌa''K�b*�f�x������b1��d�W� Y�^xjҕsX}��C'�p34%C��Z[@��M�X㎈�n��K���d|�t���X^��>�P�r#�����s�e+����X������B��h��>�:;��pŁdǰ���K�B}�"Kϭ@��V�0�*Js�k�j3��t���v�/��!�M$�'hѬ$B��B^K�yi.��'2T9�n��TH���9�����k�Re4q��M,���|{Q�~u�D:�(�<�Bnj�:&�T-��G%���H�1ώ���ọ��HȦ>Xdl��k������"#�����B>u*+e��5oQ;�)s�А�
��X:�n�ٍ�=DΨ�ֶ"t����i��7��(����ײ"�>05:z��:
u������n?g�=�zq�i�s���CpU���8��3���(��e,�}���l�z_�~t���hS�5��B���FF�����i�g�� ����)���!�3��fVd����y���z�f�k���I^��N�[+��9{���.���ҭc���ڄ���aQ�Q�:Ut̐d6��H�:��#͓w�p�V����+��N�ȼ�}�Q(ܫøZ��թ����ei0>��vry�x��R>�o�];�\G����+�oH�T�*�~(\4�f���]�Һ`eT�Ӭ�5��3[�6C���:�
M}I�Ήr�؜��}7��"���:���	�~5��T��p��c'NKX�M�Z��82��Z�O�䲛�\�+�l���V�#��PIc�ە���cTU��
��+�~����P�h����a2���������ckB�7��U�8+����M�lq`�oȶ�C�&ߙ���sPٓE��I��S��ح���]���z3)�P|aّ=�uA���2����4SA��������Y��������(���m�3�Lg2��6n�8w�1��X��g{gne���^����^=)��K���e�Y���zE�cЄ+��]�����qK��BM��]2�F�����j6H��jY5V4�L���V�R�N�j��a��v4wQ�����b��\�����u��K�I�O3��lk*��s��z��(Ty7�U�B�1��q���.�}��2��y��k�נv3�������� �h;z�TD����9%����w���|��� .�2׀�!jHWe�˞���O
#�{;���t͏Eb�4�I���J���y��C��ԃԮY��P&��J��.+�ÇiTZΧ��S���oN��Rl%7�_}TO��Cx���<�|�[�[��᎒I�������[f�S��T�1���O+�OFB�-�
��Z��Ǝx�~Y�����	��]��&���x]�l1�}���i�8jh�	̪��m:;��˺�X�UVu���v3��grp�B�AE	�4vC���k��D�:������YCO�~���U�=ES�\�o���ei5��6Τ��djy�����?g�����'��[�[�~�t,H��f�;�n�t�9�fa�;W�S��oc�m(@���c��l��;묃4ρ����d�d��T��Y��C��5�F��45nBn��r�h$NV��p�⮡���l���u/��k{��<������b�Y5�V:{�c���BԄ�@%t+V4	�YP>�ky��)�.k��a49��B-��猆(�(��=���g�*Y9��i��U��8q�J��Y�V��by������I�{
&�ǉBDy�q2���'��k"'��m$ڵ���>���cD�����m��~U�&���Qa\�2`W�+���z��+�2/P3]ᇧ�@�2���?�!�@���/�E;;J��j/Ѹ��/z����H'W�~9P`}IU��^ ��Q�[�۷�uިV��չV�o${7���P`��m���;�����ʘJ���)>�K��l?M=[M��v.���
(I��s)�z�[�r���р�bw`�+���﷏lcY����'��ZF뛻B�c4�����������F�O�~�?'���/չ����B���EOs�Ԩ�����.[O)Z�8~v/^j��x�t�d�ڎkmFy^�<��r����	���e~�S�����&��E=���G�l��aL�p�Y-N�r���ב�8PA����K��b!6�2�j9�����q��',VGB�g	ڣ)o)��Ν��ͅ�hj����(<�%��l������7����? �����~�k��:�Nveu�h�Ȗ�v\�Xۿ���v([���FҨ�0�p��L�q�y9!�ox�8N�[��%�.<mׇg����v�����]Di���ҏ��V��@�	
3�W%BdvMBYW8Q�$ܦהmU���e�X[_D_;׻����}�)�rDn�@E����27Ʊ�d��#�#զ�m|[�q��P͇m�ݠ�{i؆���b��p�:n���&���4�Q��]-�m�$i�iA����t�A���|\��޲׿2h1N%�cV�i��{=>�_������}��o�����}��o�������������_-s��q��dL\��^{�����]%���l=j��H�Q2Ha��	k�@�;26u-�W�ÇV�b��[l���l9QjB�p+�@���Ьu��<?C.�T�pS��w]bL�:�)C�{���#�6\}u�ȠcǁE+!Jn�Z�r�1�������\ʲt��&>�V�ġn�PZ}��y��X��ܕ�j�������ؾɁH*��K���:,�����}��V��%��h:�Z�ί�feR���3EeϷ��\�э�+q��]��(b{���j����� ��ݪ�������	�2Y��pP�q����0���z�>Ũ�l�:���`�h'-l�e��[��C���m����&rD�:U���Um����v�hg0���u��1Ru��T�Mp�p]���j��O{.=Ω�R��ˤL�4⾜���Y|WC�1��='�V�4�@yh,���Y֥^�"�mĆ�o��1
���+����LoEa][w����""��vTen��/����gT�Yt�`��Y��J�yݦ�4�����nnn͵&����]3�ǻO>gR�e���'�G3C�o�{�C\mv�Ӝ�T�<RX��sL�����ntVkN�.`� ��Ighw����3)ᬮ*rC�PK��v��n�mi��"�J�!�9n6��UH���oky�6�[���v��Hr2���k3�z���_��U���%��3�����>9�Y�ϖz�q�߮`5Dϫ��W�6�o�n�.;��ø�`}�?o#ץ�Κ�δ���G9]�UnY�����)�HL��'ܮt�t�k��b�޵�u�9Es$bmG���=�������S�V��k��Mh����p�f�9���E-AVA.�b�z�N�������7hwr[����cWu�|zlvO[��qS�A&�V;����C9�!���
Q�Y���jY��N5٘��r=a��S(���O'F5$�`x��0ot53/���zMuEL�򮒒�Ӟ�����a������J�'va�u|B��c�>p5�ެȄ�����U��p~�N�lU���7��ٶ�C�s�ph�XT嬎���t��Q������]buJ�o�u��_-d���A�J8��|%�v���09e��eM��[%̦
�]K n��	5�����vݤR���`��;9���]Vt԰i'VVH9��Q�70P��z�aa�`IW�m��SF��Ļ;��T�zaS�ٜp5Z�]�".�4P��;�L�Z��آ�c�(��ajm�@�ۑ���$^Jp)z���(���K�@��lcS�����[�nU�t�f�J��/s_B�M��N����bȶ:����.Nܚ��:�(Mf�8/4�4���B��`X�o�2Z�$΍3P�DQRLER[*��b
���ii"Z�N�F���Y644h5E6؊
F�)�(	���X��J(������-U5��]ɪ*����
k�$QM�N�������(��j&"-��P�d�l�4D���it�E$A�5��֡�j� `���**���D��1��LUTKUT�JEEEIQETUhMSIAk%QD�DKI0D����LT��m�4+�b���
h�"*�'͚��b�"���>������B���5�A�9����e�4v+k����f�/	�N;��(�<���<���weG�W�b�v�P矏��Q7��E�f4�<�ťBd��`gщU�����G)�d�"W_X/���m��5�L�>��Q�a#z."9������F�CJ�=C!.[4�O)M�Q�&�C*�8�՛�:hۿ��[!��M�z�5�z����Wǣ��0�NA!qnn�3��E�h;uY��8Fj�<z���|���ؤSmʷ_�\:���6�f�C�km��qR�$ױW5c^)�׶h}:®����J�%�z�|�rz$5�m͵h�>)R�8z$��h���.�38���yB��4.9�=fK;V����u��('���*�B��)��.*��:����	�q��w�bh��xE�1l�ɦ��n�fY���s(�ꉕ��-��OF�R�1�U�Z5qܡ�I�����8lK�Bs�¤N��P%�Ly�}�C[�N��V]�y�⓴I�ލtv<�AФ��I���<y�4?<�Pci�F�7��2����J�zt)|��m��-	�lz+B�-#���C6>�� ̓Dx�C'�<�.��l�{����>օv�Pv�����.�j�p�<��r ��dG\yY�к��<౜u��Q��3P�Y�������{��پ?h�{�H�R1�n��o�GOx���]���T��WI�F(3��<��B�U��b�+n��H��l�r��N��������O������d8QCo�L�q�t�e{3�'x�g����P� Xw��=�?,��ێ:�ݚ�-�1����U��7u�G�%n���:Y{^ZJi�8�g�̫�<I��.�gb��^�yz��6�O^����x�w�wK6��3t���W��VC�X�w��U�&�1v{TD��c��S�5���~�RK!�����&�H�C�c&#���5-k��{f@q�v�!��uF<ڡ�5�=􋌄�Z
��)�m�(n�sUqx0�;o�s���l�C�g�8:6�*m���C��W�8|�/��tɞj��¢�W�� ����&�[ݚ<�wCL�lz�2��S���H�%V���Y1>5ȇ��ے���z��]�t����������sʌĦƿ	�>)�2}>Ŕ/lrVK�ò�1�3��;_2�&�ua�k�l�<э��q��qm��)�桛Tn�ä�BS��~�b��7L��2iT��V��g[�¯6/r4e����Ǹ���K㷨Ls#^���5{5Oc���O���.����+/68M��!ظ5Χn�9����y_4X�v�����QK1x������;3yr�x?��s��/��($�{�G˩M�t�f5�[�J�^M2����˘��{/F��	/0�c�I6Hܻ� %���Ԧf�%(z_p7��Ϻ�Q���ĳ�f��S�����`�Ř�<�I2%���+�q�a^��kv�Dh�����O։��Տ��ɘn�ko:�)��@�ƽ�V��
CLlV;;�~���i~�~�ٻ9m��K�M��m�
iо2&�OC��E���<��7Ia+b�X�h|w�e��p�+�FA4J��%�O'���E��W�WC����ϵ��)����Z��iǗ71F6p�k�����wp���4y�.z4§x�/,�c��0�V5.����.�mjv���P��Ψ��xn��~�L����Hy��Lֳ@\�t�'T��1���-i]X���m�ʸ9zcM��u��t��h~�T��F��ʮ���l��
���cCT�
Ȍ�XTٳ�i�kC���W����`�߃��R�d]"&wʷ�\�Z|��l�=a�a�׵��0�f	����ֶ;s����|xH� r�`�
�hO@�>���d��-^b��
���Z��Ã���˸@e/H����65��d^��J/TS�}U0ý{R���o�صQ ���_5��L*��gu��nV��؀;M�񔽜�X��	�y�ƻ@���!xy�)�dC[�����tR��6i�����&��A )��R"�:б���2���l��Ů��|6���fP@��rj�E�d;.՚�5TE�^�$��0>s��G��5}�zji�:��5H����U,7�l� w�&��&�]t+ƭi���Ը�@S3k�]��e�D:ק|i����j��*M7!�ūT���#��xA��1��8[$�1=o5�1�J-�=\ٷr�O���1�22K�Q�-2���JBh�GP3�(�h���'������w���er�n籅M�W�9D�;&�s��-z��P�ì��^.�g= ^L��3����Oѥ��N�a`%S�JSM��q��1�GLg�D[@I��N���5&��EY5V�zszֵ�9�9�H���8�� r{uϭ~J�k��P����B�|nM%�5�(�`��|{�I�c��Q�Iqpˣ��yyN�PYm�H�z��ȋ|cU\�tj,����Cc��1p��0��Mz�[&ԉj�fN@P�',mC���㫄�֓�9ZnK���Q�͊^�s����A�<�W����@�dXw4�ݳT+;�-�4��N6�dx
8��(���_�k���7���z<����$��j����6F��.�w��nI\*��=}Q��uؖ�VQ*tR̾�N�~-�lp�@�;�[�s6��[i-�o���> ����fp���aV��� ���x]w�]N�67�:�;�ﶮ1�Cf����f39�G�i��1ݹ�[��~2��O�����Q�i��h#�k��*�!�t�����/��ǋ=�S��Y�������3c���H2��1���_;��47���<����N���@cG���Q��p7���5�b�y���ɶ�.9tV;6q�,/�Nӱ���(w	�6��6�WE�'��I=/b�T��vu��<I��K��j�����=y>-�Z��ot�O(�ʼT�jZͱ�/%�"U��1��^;rZ1���p3{l]��1�l���J�k�m1[u?z���c�z�}���r�AG
��R�.�����v��q%�3ţ���MҖ�Gj���tmxp:�\�gO�k��GJ�c�6�*Hl������.#Ǐ"c�f	2��gj�tQͽy��65Vm�`��l�&bM����\��QI��M��s��8�/"������$4��o6�Po+�:��q�����].���lc�Ri�����^�n�v��֫��'%�zEpq�{l���ۻ�*2�j��~a{ɚ}"7>ۖj0�f����������m*��oW��JܘP��lQs�{:u����[��Z=�@�eS��Z�3J�K8v��>��\�q�@�[��M�^�K:n�>4	��k�b�1@o�Hti���h�G��K_N�j4馮���e�]�E�!�:�rwp�:a�e��,&eG`��Q�:X/d����m���ط}��͟z���/�i�1çE�K�a��i�&��aR'��X$�'�pȧ�m��h�Ӳ��*Л{�)z���໸ia�A�$��^��cՒ$��j�d�3�>e�[��u�m����gf`��ЅvO0��K�Gu�?Pft)5�C�L����y��s�7Mv�[���8�Vݛ��D,e��Uz����z����.zKv;�>�b(�;��n��LX�U�u�[�M^�v��	q�b�Ǥ��s�A�^&y8�H���0#5UV����0���gjf�'២Rd�3e���]�o�u>a�9��q���@&�I1t�^�:�LE0~I�e�L=�1���G0�@��^�fݐ�^q;�9�`Ht�7�Ʒ{OF��9�˽�����l[*dv����so�S�t?V�=��NVJ��*ySo��;���r}ꪇn9۴�pg�g�6v�h�ռ�3���[�f�r(�ܹ�w�c|��a��cGx�4%�65ı�9M0�����ob��T=�[�� �
�͕�q�����٩x~��2M�����T*����]E�t��Tc���tﱳCut����&~�u�(W�m��+�j�݉L�\�o��Z{��2nA��P�;�gh��i�d�����8���ݨ�K=����gG;�{Q;�#ca�5g�Rn
�]�!'�+@�+��jӯ��n�>�f��v�d�Vq$ԤU�qL����_ş3t�1W^�_��Q�u/B�&�	]
���XSb��|�}wga�0�(���cY����1��?@�Г�L#LJlk�S.}O6�qe��s\1Y�9�F�59��v-�/fò4�+���a�̓;��_��F�m�2�޳�I���Ou�I	�����&CB4�'��������s���8���0�|z��L��B�3F<_s����]V�I �S�3j�so-����]t7}=��ڋ.2�@x�e��7�[����'y��1i�a�&38:ʹ��Sr|uS�m.�n�\O�F�4��XQwl �}W�s�u�X{�ǫ��������k�H���⻭Qaj�W7u���F	���- uE�nj!�mv]����҄�c���.n����V�]+��OA(%�ZS�%k\��A�H뜄О_vOi����XA�3G�G�f`��=ܖ����A���@����l>�z��j�����^]ѯ@�=/Z s�k��
�ټ�d�!F4�� ���G�ԫ3�Ѯi�,�ٖ�;M�F�n���m:�L�p�Eg��s'�"
x�}�O����hC�w>q�2���k����y�%�����.,�B��ݜjթ �rnRB�{��%�`�X����6����6�٧t����+���J+�c5�9��7�t�� ���s�&���e����}��ު�������}~�O�t��ו�-�Q��P���4ƃG����Q�o:L����3y�Ŵm��l�R������>P5�BI��:{��,����#<���H�Q��.i��g&#�������P�Vl �ò`�r�:#�h�yM�iM�~7\���e���OfAi�\����d�����=q�SQk"�8Q��۶��~n���eE	#ڦ���WP�����Na�MVvN��7�_w���`p!���Al
EE1�J����+���I]
Ǿ4��4ƿ'�Y���|���QD�D�9�-P�Z���̚�j
�Q*Y>�*��\ѓn�R����S.����/.̱w�j!�o�A�fL��g;�J���v;l�9�:�h��1yy�ĎȢ�8��qJe�~�+��m�-�a���^C��p��.�B`&Z�gH�Jws#��X��/eQ���tÔ�1���ڋ`7�.۽���L�зU���wf+;בb1; �M�.5Y2���!
d�ߟ��9lN��R���R�z<�A�?�S�����7��eW���X�9�af
g
M�B�����b[&�	:Lph�H�ӈ�[-o��Ԙ���\����g�sƵ���C�{UΩbt=���8�Wv�ő�F9�r-UJK�E�vz���d��8��s�w�w�B�
����1o���(��������׏*%��-��#uګ�;���MY��\�$��Zy��-�@|w~���R%�Q�b������@k�jێ]��f�|���=�~^T��-�6#� ����F��T���6���]2Ɔ�;���!�ܓ�S�����E�	��u�j��t:�ጇ\E5�P*;΋�y~�C��SqfFA��g{YM�nh�Ok�P)�t���SH��4:��#M�C��u����!��<#�3�ENgY��	��/H�I��3�̤�GtbǢ/���	��s���PB�$D��ע����W�O<_IcCY3Rk���SP��W�ٲ��ߣOe;�<�^���V;���P�o�*ퟺ"�����:z�`Y@�(OT�`��U����{�B�}ast���Թ�J���9B��sWH�0�r�Jl _Ch�e�'8�'�b���[����o�ᷲ��J���l�Y{�Sk��:ͯ@���S����"0�gJg2�p�I��	�C��fW��zJ��7:�2]G6���Te�NRV�,w-��wg�F��O�)�>����pT�o{׆p�n��b)��n�];;UI��2�֮���5��n��+&t�u�F)�X��ۼ�=��D�}o���wK[9ھ����m����^M]�k�.����pъ'�7�3��Z��уzjj�ɶ�-�c�dL�[�0"õ���.�pd�Yuº���K��wj[4�a�����`�L��s�9���w�i��O'<�G�u��W2��`%d���ƪ2 �wf^�yke%�E�I0�a�u�s*�t�w/m0`�dR�a�a�f��F�q�*��Y�T�;�c��5&�LW��>��,׻!�ƥ%��J,s�|ژtǭ���t���3�M�p��D�bNT0�$�i�1��GaMXe��Q���3�EU�&[��+-������mfo�����(��/��9vبq����ٖ@8%��L{rD�d]2��]o-�ůwrI�a�[!�ʔ=��M�A# �~�@X�M�������5���}�O�"���B���K�i���uO�O���$��[%�=��������8�h�u��������3�۶�E�����r1L���(��s����c���J|lcg��"6�����cF���d=����w6�P�$05���"�����U�^�v�
�1N��v>~P�|z�=}?��}�x�}��o�����O�����������>�?�n0;�L�o��_�O�̋,�z䥗�nVӗxM�ɺT��k����c^i�n��e��,	1X��ͬ�ڤ�IΔ�5�/��is�d�e�Y��.f(� B������Q7�!�
�4�`j�wwӹ�;���B�X�g�)�4��H�19[�瀌m���5�
��]�V�8M�Hf�HN엥S7�e�6�{�kl��V��HSc����;�Ӡ�l�mG�]�6>z.U���a����\e���@ct)\B<˄I��I��B��ή��FW_.�9cN?�%�~q�������K�Y�U1=Ѕڮo]����4�6�uiZ�seJ��Gj����
S�a=x���N�3����xL|8�s]ګ��7(�%�&!NgFL�Ɩ��F^��غ���.<��ѓ#�%LR��hgn�ل�w�՝�b��*�ԻyHe���VmM��T�3��t/�!:�7h5��ּ��m�)!eήB��7��:e�9il�l��W>G���X��n��si3ϟt62_,ƇW�&��F`�����y�]b�oV;�sj]�(�����xXM�w����q��etlq��,X�3k��(J���k�[��=�u�xc�ٛV��:�W_܊��[nf�\f��8d�;k�V%}���ܝ��q�	���&���#K;���/o�u:��1�t<�N�Y9}�LԻT�h�j�R	�Wv��09��δmnY�=B6�t5�r�
�r�X:�A��w�۳Yov�Tu���l��Rux ���mV�۸�u��&kш�ާRed�%Z���*�Z��#���kx���ua��*"B�m�t._-Ǳo<�3+uv2�pul�(Ⱥ�g \y�����^�Ȥ���6�rn�,7�u�����D��[��u�����y]�tt�U���9m�h���2n��]K�κ��p��!�Z�[�|�&���s�m�6k�d3�&�e���P����pu�DS� �\��� )�ݝ+M�4V�B���[����cp�F�E���H`3j4خ���]���0Q�M���*�}e�0M�Ì�Ez:.l`n��N}�Q��
bm�٧�3�\rd���J�X�`v �����lV�z���e�|s3�����\Q�rmR��sc=�T"u���u��V>ӹ:���1��W��"� <�^�Ep���-���Z�c{�l��j�˹]6�t8��{�7�{0BS&-�'U�-��SJGm��뫑�����G-�|�;t'hyɘ����|�;g*衺��
b����4ދC) sQ��V�/GB:�WV/j�{&6�*h鏥zz°��)� R܍���JR$QSO�7��F��j����2�'.�S4�xZ|��M(�;:���6�{93��ଵuo�h*1J��VM0���_��;MԶ֝�yk��dߏ�|�ED4�0SVɪ)�)(��)�i#X�*��f���"b��b1���6����P�i�QS%Ψ�&��`��*����b"����M$��4�ET���DMT$CQSEER�LG$�\ږ�����&h����hq�h((����(��褢 (�)Q����3CK����"��
����cF�i(	$���5���$i����)(<��&$�*�>��מ|\����E�%�Q_��D"�ƙF����C{uu���@��cO4�;�ǣ�g8ob�}�jEvǼ�w�7{��L���w+j �F�Se�I�S	|�� ���Q�K�PE�L ��t�eM$h�������K�O�����CgT)'ad���3���� �X�Fr<�����LCWG��Y��J�dE0��כ��I��?�9��~�~�/ǂ'}�Z��&��	1lS�oF��kh
�\���b|���^��\�c�ي����Tcͪ$Cμ������3�zCt�{^�Q:���Y����5�t<�W��"]o�	/�<F�W4a�����:����+������
@DY��}��7LSN��_�(u��<�¹����5[Q�ǰWkS�<r6�¬:;��RԀg��g�7<4�P��ו!�h��Ƣa2OcRscPܺ-;�"���13��<��D��v�0��vF�-�j-��p����R�1���4(R��Cub={]"(hڛ��-�̽3�ڬ^���c�X<�͑��g7E�CIb�}�h<;T6�_O*���eo���)�߳2��.�^x���)����O�.��ә0XO���"Za�-z����e�P���\`��p>�qq
���U��L&�����0Xג��(F��q>�p��o?���5�	��zA�oW�n\N��n����C����7H̲�^�0��Lu9�����k��g����o{8���R���*t⼥O�c"�T0LS.��|�8±qF�\͵���nM؁4�P)���sa���� m��)��t��r��x�B�:��-���,;���-� 3�I:Zg��7Ln���)��"�OC���	ts.cS���kH����姭��Q���!L��) ��DB�7Q�k�UiU��b���'��C_%��Q�j���.�/��Y��U�@(f�K��/,��-�������"k��`�ժ���I̽9�u�x[�@6�1�	띃��Z@y�c�߃C;�a��iQ�й�aN��-�v��[эt;��kק�D��0Ƽ`3o;�k�P�"F��q�ê-&]і�gh\N^��P4�o�Z������gr���_�ז0��(x����D8���4<bJ:�{���	�ߍ����#!�x�9��ò�l|%CoD�͝>@?rl�dP)�����r{��P��O�wܪ���b��}#@��}n�s��j�tK�GA���o9�f�:��`3���:jip���0L�fV7X�2�Eo	MT���K;�r�:*�v.���g��U����a��3�,�,� �޸�1
�.+����U����{x���
��D��c2^)�Z�K�d,�;�r��I�¯���X��.�jQ����ۦ��h�J�fw���G�L�5Oa��;�#�f
�ٕ0�k /n��;@Ov���n�LW'e�% Jsf�3��%}o�s��C~�[s3�d�{`���n%�lwU_����j��{Y� N&d���g7��^P1��zǍ��6�uwT��j������C�eMsw�X��{����7���M9�u�Xި"{�Р9��U3kNV�p�6��t5�h��ȑ�e�=�t�ҩ�'+��gX�E�C�8�r�O�CJ�__�<m�����E5���j�s^!�+�7()�~�O��������L�X}�vǱd�c������ �RȨ���""5��z^@��T���Jy���e>Qm����<T>�	���1�z�������8�5Tt�ׯ�W
iBm7�m�jD���7����OeVnG�z�����4˶V��;f�C20*z�]442�~:'��d�]h���g+��(�5�WV�˩x���C�d?��kK�o*7�����22yJ"��_^u�d��<��	�h�B(�=[�1���	>P�[I�2ӑ�S^��G�Pw�$���]�lI�yr{�v+������>�F7P*A���1�J���'ܫ7�]��>�����P����>V8f~��o��~�/ɽ~B-�o�a�.��#1��#��gP:�Z���o ��!i������I!r�e��6������C��'�M����K�y;K޹_���^�5S	�������%�`;�#4��k�N��
�����f��5$�%��I�:r{�;^��w���!\��%�r�ʇl�;^�9��Cj=�A`��s����Vf��s�5|����le��Ax��V������ɶ���y!�����v�#&k�,kL �7rL1�ك�)�<Y�.�!٥��x��a��W�6өQ4*}譮���K�ߊ��=�;����Ke{VS���I_L�h���]3Xv����c+��x����[[$��W���c�F�l���uZ�2i���c�*�m-�Y�r^F����.t;t��l���S�����iv�gd*bV=�a2籊)9���[
2ިr�hi�Zb� ��:�T�]�6)m���"�ڣT�O��h�cxc�%Ƈ3
�yJwX�B�Ȋ�B�J&�h�oiƕ1��d�������������j4^�f����9���fȼ z�ʅ�I�[o[�F��졷=�!���9A�1�^��1i�M4L�D����`v.���<u��J���G�t\���.�5��cj�H4:/!��������?!�¿S���[4�j��<�xJ]K0��X]������+ �c"Ж-u���J���� ��naT�!:���X0vm����e�D�u��*Tv��c/�6�K�qj�yغȓ�-U2C2�}�o���J��؜������1[��<���S$�B�n��Њ�]��S��w<�#��2b�Os�a�#��]�ٱ�C��~˕�oEg'����/͔9��:�*����hO�6}t�KOd=����l}H�m�o��I�k����[-�*fA�@Ǉ/�A�wD�zO1�"@�g���;�SP�v;��~&�VR�VUc�p�y�����D�kv=F*j=��[�W>��T���%3��cbS�H~n�Vwii�����qF,L',ͽ�c��õ���2ˆkn��^�ip�A��:�j��V׫��<^��t�ʣ��$�=�:N��?�UX9;?q�#xE��D��o6����j��H*79��͞�tASp进T<��^zBZ1�|�mr��3D��:1v<4�k��V�MCV�st�P�iP!���w�7$�>?�X��&�B����ګe�@�"6�z]K�u6¼�,z�3��??�6%r$��Zj�V*�\���]�S�Zs���l$K�X����D�@trw��Ѧ%5��a2籊)9oO����������Q��5��� �@p�~ބOy�أo�:ި*p镥�woT�Iϛ����yP��3WK���W�+T�yYz�3 ���nħ�Q���l����P�̽|���^�{�-�Yxs෢��轝�+soz�TQ�$֜U�+�v��)x��qy�0�o!ؚh��{j-��g���J���^��k��K �$�F[$�f�� .S��b�z���`+'%��;�ٱō�/�R��ײ8];b�,�����\�E��c�O#����K��߻��еەwLzb��O5,����\�N���*�-��i�i��(��+h��]��|}�c��s�K��m��n��{�����M-V�rV��ז��e�Su�.��wMvt��zf�=>���ߗP�bҙ�+���ve*��.cC+����XL��.7��͍@MףϝA�;j>y�O�
��&,���:\��sFꬖ�;����;��w����Y^����c�1+����K7�v��U٭���a-lsut�Q|�GN��ͽ 8��C��5>[%"�_&z_;w�c�в�tg�͟�ZA;��v{����;����?����VS�v��E�fcs8~u�.K�ٖr։2 �7��a�i�.�f_w��:q�63�t��J�g^��|í����N����V���o)�U�V�9�/�𗘶i�z:vu�]:�y;H�O�|�
����V�Ŋ�]�Vk�����gdo�N��a���J���'z�|9��,@��Zg)�¤���"���n�]��g�w	�"&������ot��!�܆[��FlS1��nrΓ���xq����}�j
��A5>�05)���\�̒Lk��f'������^-=e���K��[3.3�1�Qٮ��Ct�����O�qى��xf}'�:�t�A��Y�r̬V��4��-q�׌�L�s�&��]��Λ����#b5��k���g��Z�7��_�����֫�y/��۷����k�C���o�)�7����4td�����
��V�%��d�6����.���N��Z������ⴎfR�.���zޥ'�$�Z���Zl�g��{pF�?@��Ƚ)�Gr)�CTs�@Y�u˧�c>�z����N���� ,��K
��wG�ꗊS��?���7~�Cz5�%��t��0����Ю�Ȝ[lA4��O%��!����i��NZl��e�n�ˣ��C�\�hy��k50������o_M�px�棹��,�Z��y�	{�j	@����������8�2	�M0�;*�"�$4�(+S���k��4�F�K��p����$��SCT�m���#�Ra�S�[4��Q6���qcoD=�G��r(�q�1��`jh�s��Xh�Z����)�y�ߦ��n��>Y�����z�����䎙��à}�r��UhE�U�l'�խ�ܪ�CM)����s1*��f=���j�=��tQ��!���v��k�{
����;,�?���l�r����G��6���=j����c�g�!�l���ѩ;Vt"�[�ox�@x�P(��n�/-��;ka�ۼ[��0�z�I�R�hS�|ڶ��$v�~*]�Ǿ��q�c�?A�Q�WT�;#z2�ut���s��I���l��w0��#�XY�����Kf��1tlZ�RTe�H%]6�˝b+��Y6���6��2F�z�����;$��]&���d��kIwTu-�_Om�[@r̬�x��i���0��+�9J�y%��(.5w��ǎ�7�O	"ua�o�3��{3�=�ڐڴ�]N&�2`飱�����J5ZE� ��W!�wZ�kWJ]�X�MX��؆@�8��t�A�(��F3E�bT$��7�?��G�6|����mjo��Kz�����n���!��uۓ�����zM�Q�y�Kkܸ�췞��g����ǯ&L�F�ݏ��ݙn3�[�[�Ȫ#�d�.w�KgwX��w&�@h]:������4a��K&���[0\6�u��8���ci�����+�_��������"��/�&�4�ٹ�����;C�w&���*��^@2���ur�n/��σ^O��7���?>��*�N��V)����:d6j+pqeT��\{��,jl��.�����֫\������f����u,��U�9�!X[S�J��7�kb;��n�e��g�Y�;�Fh����w^4h�����QzN�Q�m�έ�6��?_�Ώ���fQB�F"Y��,�{�D��2�E���o��Fتu��oH�g�Я�oG���Է�bT��֞��Γtﾱ�������L�`m RFd{���[v�*�!�V�z��2��kr��G+�Tt�k���A$�מRr�հu��XZ�n73�8��ૣ}oi�9�5����T�U�����W�<��ذ���	�-�p��p�<,r�Z���mL�fڌ�6��#����yܯO�MD��.�gC߲�A\/ �S�����Y!=b~������9���@���,@1MV���T�i-�<�.�z�9�]�ӻ�3y���W��52��|���jW(�A��
�0��ڱE*R %#sT5������i���Q�Vڥ���ǟ�\�pRη	�@��eQ�r��k{w&�6���qK�#�[ ���W�v�kq�6H����j�pH�����{�xsx�l��K�7���H/^����ZE.6�u�ɠ 5Ds�L�u4z���f�Tp]6�WsFiJ��r�Om��Wb��[�d
�B3[�m���Ɖ����߲a8� ��"��{2��99<�?v7���j��uqsZsb��j��e<o����B]`K��E�����ٮ��_������~�g���������������x�����}>�O�����FM6�zO�Y��z���w�}2�&v��&q�G�9�Ő���
c6�Ld7��IđoHڲ��IΜV�Iz���k-I%��:r���N����%M����l�s�����o�ɵ���<���lt���$�jȭ���{���m�m������`�;1�&��N-h\�v��C���U��2��2)�C������^{�v��&�mj,R�6�L��]�L���m.�j��A�1�s�rt4 }�/Z��$�;�؀�:��.�����s��Ř��J�0����:��d�v�@ӗ\�N��Bڨ�*�+���GwV�2��w%-�u��9z�Q�Y��$Q�t+^	����.�tw�Nc���)T�}4W B(�6��0��{/������H���}�:�,+Q�@c������ƆS���|���y��-]{��촞���7��Jd��4�.������մ���L��F��Qu�-W]��s�΁�9A���5�JRy��,n�kT*�b*ۇ�m!���Ȳ�A&ۦh��;`���5�\��|��p]��λw����R��lk�f]f/�G�P���v�^T<�f���6��M��n�O^K�;�%�d��t,"O9�6��}�a1���t�>��Ρ��p�%D�W��!>A&r4m�9� ��-��/��$���Z���^�7yӓ����%G>�$�\�%��;Nvu�.���ux���g�Lv!�p5m*��
Sz���'0t}H��&o�_hW�Q���ۻW�}��(Mui7TW<̔=�����"j�BL�4�W]� {�{'e�QɀL���wq2���ӝ��/C�T�( �>�"�w�FZ���t��n֬��\�f��Y����/6�{�}э�2����[i��tm��ٽ�8oe����ǲ�лt���GY������K/wV�7�����L�ލ�8�ӗ��ռ�h�g6č8Nv���C��-q�l6跧�3���{�mN��a4!�&R=����ۧ $���YĲ�r�2�gk�*��v*z&:�w�%��{�> �es����CR�]n�X(<�nU�k�gN��gZ���!x�}�`�+6M6�w[v�mҶ��N�c4񥦴�[�8��o#�7lj<݁����2�Qp�ސM[������(�E�ϷA#��8.�&Y�g=ESߴ�{�6֩՟G�O4j�lX"#y�+�(�x�Ia���3����^���gQ�]g��4��WU�m��)��3{(.���)��L����81jL�p�
Wq�|�Z���Wr� K�i*J�A�K� =��TǴ�`�9h׸���fj��8m�)]��Lٛ�4��3�����nV�*\�P�k�h�����}�G�o�#/$�(��v�	�BW5$8�ևk��x5��nT�#�ܻ��Tf�h0�!��\�V�v��7���u�8u�u��ft�A��٦y�&�
�h-�5�EP�M-K@PPPR�ĺMA�5ILF�DUBS6�CSUZ���44�h�SHAlja���c\�j���9��&i5���JX �"j֨�(��*��(�-�01mӉ��Y�bJ*�B��f�c��J���Z6�4�5K�@PD�5D\�JJb�(�m�Eyb
��`(9p�cmF�:F� @� P"�@)��~?/s�{\����2�S�MI��8�K�j��<~��u�Zf��s�¥�K|�ᷴ#NZ���i�f�I���s
�g���{Z[o����;��2�"#T�!@z�o�����^���-��7�.6U�{���z��Y��@}�CbR m�|�0���4ӡKH�n�8?^z=>Ӽ��t�Ș�ހ�~�m�L���B�hi����I'�YSx�Ӈbܜ���I��i��FΎj�$a[C�7����#<�6k�S�����ۧ�����
��JqLi]t�K�_!��;g�E?$bo��^fS�otr� ��J�<�����<n�D^�7�u~��Й�)�=0MM+�OqRj�LN���Ȯ�Sd�I����Fj�Dzʸw��{��Mq��
9Z�4�b��9�"M���-������r�9!
k��ힵ�T�u�ɺ�$�1M�yf�����V�٥xpT���y�ͫ��@�J�J{o���uڡг&���!7���{�Z���>��f�Gk.9%e��u�\�B�oh=���f�a9]��_��.��9מ��W��p
�l�}�#;�{|4}�����N���/&�t�,��T=�wZ$�HS��.��X�o�
�5�*3nVgGg�z�{�o.��u;uq���c`�l
��v�}��i�]�^C��brm��R��V�l�)^1�W?uŉz{����6���WB�h�rO�TY-E.�2=��v�
�)�ͭ���Yeo�Y���^7�ҢF�< �,r7)�Q9�ҟ}����P�[g
׶ɹ�8i��9^��fp�c̳�L����4o&iUg��`�3y��A/s:u�x��U�}	wUX��5��&�݆�@�j���}��m��j��;S�O�	�uӚU�9���=O��y����m�l�g����s6ǭaӳs�m��s�#���&���V�s��U%��m���~)3��Nݓ�h�Ǳv�T�@:���gI�g�݄��n�r�;K;c�ׇ�����^n��æ�3�=S�ؘN7���?Qr�h��;����O%R�w0x�8g��� vJ��A,%�3�s�4(��/����yX	�[7�)�[
%�7<A��7��������w����W��l�V��|�ڗӕ�;q1V��Gǅ'gq�����{�29�vQ���o\��f_Px��9vܹ*�xԦm]gj���y[����!����b��,wUo;ڊ�\��Pު�Y*s��e�R��V�wGܸo.�s,ڧhǎɡﳷ���um���9[4����������mub8;&�a�4u_a��ʼ/�jo7<��2BQs��IV�a��z���wx��ʘk�������X��J�4��䲅���u����beaAK=az�W�v�5���ڏ6�L�z�3�e`5~��ދ߶e��C	�_��fQ#=�V۸?�����96���B&���J���.ݺ;��sM�\1�ӝ{Sv��\`�ڐ�95��D�W	�l�
im�s{�#N��;3�#��A��x�l��N;8�<<M_Jlݝ}舕�8�(�o�_��w�mˊ��w�^��dXXq��.G1Q������aݘDǧ�=Z�E��`a�-Kt��P��퓸̌����pgE�SD���"G����<�"���9������{~�=3��x�Z��pŹ���q��.Z��Me��2ˌ�vn�d�ir��8dz �[�k�_����:=C%{t�@fг�1�2���d���TO��wμF�1�¨��eK��P�����:q���u`��^m[���ܮ[�Jq^>�9>L�1$3�sU:�%�ރ S_uv���^�͈fvHg���샆\�2���M��7y]wj��`z�2�$��4V�x�Ӵ��>�q�KW��@p��b���B��Q[cv]�:kTQl���X�$�[P:�zk��9�|����x�e�U��8;�n9�x�vѦm�����Z��y�h�Ut���Ta��Ϯ���]qw+�n�OU�Sd���vW�[ ���~m��f�B��<�	�V/w��n�T�nöπ����M���/5�i�4�뎊��]豵9%��X͊�D�K>Ϛ����{y�0к�mu�j�*���D f݄�nbK7�EymZ�m�G���y�������y��9�*�h5�nx���ʜ׳a[�yoG���Mcla2eѭCzI�K6���u���D]��<�+�3&���Fn̬�y�3OTF�糹q7ӈR��
��v�����.f��{|�T��Q�sr��?�nQZ���c�1�W�.q�뒬f�;xm�pQ�yٵ�K�/[)�ލ����a���'e�v�����h�l�,��c���`XiY���wI�n����Sl��q��J�{f�S��:A�p[�o2�E���N���է}9}�R��;��>�Z�ow�i�.�~��+*��1��;v�uT���8��3|��恚R��\�2��[�%v&�.��~����8w��K=� ��;�-�٤
�J�]���V��w)�\>�$%����]>��Γ��9�b���E���}�;�jN�OjL���	uv��bW;������F��G�e�е��|Fl>m9��|���څ�5�p�8ˤ�5�<^�/QIm����7:VA��0�A�ģ���|�n�Ɗt��vd�c�s���|�����{��};ўh���y��ƻ���F�ۑ���/�3����jE�0���͢�X�����=+B�Y�4Lm��>f��gF��P��>�|jI.{����ԩLx@_��^Lxxi�y⑼D����7*�os>��W�.	c.�o�����|~��ؗ���c�x�\�?[��j��&�l�����Rp�娌�����,�����+Ьy�#�����rmor��ƽ� s��G�3�,v4���,��֟4�<:�+��:�u�;Z9�w��3^Zy���\{M��m ��gn$�Rޫ�v�4i�R6[:C�G�L=.���C3-N�`Fm��x+x�ssE�j�W=Z����/�^D�1�l�Fa4�M��m�IY��\9���];����5,ͯr̪Ŏ�����L��Y)�&w;f@YK��Z�az8��d�t�� r��T��d��f�{�Z�J�|�t�H���|R��\�l��]u�|�j�-���Fǣv��;Տp" ��y�*�Ե�����Z��5�sWJ�V��5��ݞ��W�����2�3)!\���Ѕ���5�í�#`S�+K�J:un������֭.��OW��������k1m�����B�)�Q/�2�a��=[Wv�E��ڒ&�K��Z�b�2���})�}��VM*����t�9�ڞ�F\��ʧ�;ʉ�u&�Ԯ^295�c�����8��;2�v)�&�����7�p�͐TzWT���1�y�3�WT�Z�~��AT��l�乼*�z��9�M1ӳ�2�WX�A���Tݢ��X{��S��ʑ;(�+��Ĭ��9�Q٭d��n�_I
k�6�R�<vd��:Z��L�m���W!I>[�;��,��}����x�\���<��n��ׯ�:gF�A;5�U���W)�FmL���z�n*c;�:E�@�����9Tq�f������b�i�?��<� |G�'�ˑ��7G�dM��˭�C�,��wn����Yk�`�r�#��k�,x�k/��(�.Z���@�m��	�Qh�ZxO"��`�[#��@�NdfPK=����[�z�W|���5��J��������^��1
Qs��IV�Z���`�z\��n�T lG=ʺ�o&|1r����9fB�	\�+��jF�ά�����.�˻�L�Z��N�v��9�<bP:��}=�,�֘�<�3����CU8Sh.ݮ6�L�q�mɬQ%Y�2'�붤�!�ik���rkx�&��z�Eu-��"@�ڟ5�N�|�Cyx�z<���U`�B^�E�z�&��U�mi�&@���B�ok;$28](4v<��uC�rqצ��)
�W�����o���E��:/�o[��]/O`V�xH�7�Ϩ��1��tn�F.����Yl׀�v{�㏟A]�D��N�	Q���pL��v�^Gu����1�:Oir]�S۷���r#k�m^��J�E鉶h�ٕj������1-��\ZiR2�X<�|�|���n|�xTM��Ub"�U��;*a�B�r��4�<��Iy �%JQ=������j�%ꚲzgx�1{�|Lɼؼ� ������
=�Bc�W���ְW��Q�ٮ�������Ob��Un��{�'��O
�ah�}ȹ����F卯`�iz�1�o����{_^֑Ⱦ���U����@��h�*p�dU��P���{�����s�y�`�a=��M���J�o��?X#:c��x�����ْ׷�+7r�z�P&0����^�O���n����w����p�&"go�����mH���2��56��:O*'U����Z�u"�7.���;K��g��Kg'��۷9�}����o)�����׹\���?���Ϳ���ه��۹.��ކR��ճ�9�w��7K/0�/�`&�a�$4D�����Vk��;�%�
b�UoQ�T��kd�7�����1t����M�%mI�0�V�����5�V��#����ո{'LS�#����#����㍄M��p��A�g�߭����=U5���n4pOJ_ H�[e��3{y�xɋ��W`ok�CT9rޕ˪�-[]um�2fo����6��RF��Q�W��{2��X����q�<�Pf8À���Ϋ�'�����������yr��["��T�~�n��Z6;l��)��fNe4;�a�]nE��E4��,c�����]y]=���{I��nnFq��|^�}&�p�"��s_���(��9�n�K�ډ��X�����l�k=�o�h�ȧ�~��&5���M.ab�VD6��u^b[��7+�甎�ӡ�q�yav��E��z�L1st����ݜh�;-r�q!����L`wf,��k�ͳ�3[=�����vrO����C���n�k�9�:�-�%�R�^��iW����0#�������'	o�?F*5��\�]����һ�j_/',Z��u� �Ѵ����Y�;�LOp�kޭ)�{<��[׹u�����R���f9b��4�-_i] ���t��6"�����aPUm�.���'uӨ��άF��C�uX��7��;:wk������"�6�y�
owuΎ����!�y����q&�f#�ܭ�z�w�&�ڑb�Hv<�ޖ�l���%v7x�ƞcc^�{o�v*XH~�k��O(Y��ŀs�1�٧�׹��vghy��f��s�L�w���a��Q3 .O�m8Zf`�e$��1ё�z�pўێk�><.1S4�u>�l�|��_�E� A�lƂ.P�[W��ެ�Az��fEv��䶗,��`v*w�j�{��[���#���*ly�]�74E�2�������SKg�����]޳\C�ui�ôWU�3RolL�+�".���>1�i���Գ� ��Gjݙ�U99\��ه�8[�|͛-R=��}zb��.R�D���|{���8݊�n&6P=fA6�UE���rf!e�Z�%����C����������|��>>>>>>>>�?����������|}���0+gmeWZ�E+Ԫ�tv8ɨL-���5R�z�}�:�ׄ�A��t2�.�6[����b��Lل�f�t����Mk�,Aw&ݾ��\4�z�Ν](�곴��雙��n���Z��ֵ��z���w+�
�Yڐ��y�b�S�g]`�T~�f�R�pq8�i�S~`	��c���3Qniݘ�/�+p��c9��ܕ>�ه����Yt�fe0��+�g8�%�6fo`�¶������y���8����G0�\���$��3n�Z^N�ٍ]�d��͗����=���l������Dn�ԾG��BY����Bq��V
yY�Z���I����[F��\�%j,���s �\Z�u{��'��x�,]RYv;*WU�8̌U��/�����*7#k�3��9��t��%)ǩ]��8)�mc4�4:so��;�ʃ5.H��šXe�:��5vL/��*h�)�9#tl�����b�^]�����𥡊Osq��!��>I[�X�mp,r+�\4I;@�e��.��"F0�5xjb��5n2��g\���}�����]�L�JS�ƱQ��yp�Oc
Ѧ�
��]6�|;�8�IJr����Y��� �ڽ�yCn�R^j�L��}0�Ku͍�wi����[YtU�jZqfYZ�,�L�t��g>'�)�;�b�b��L[�1�����˴�,��\�;_q��f��3��Gx�vP�H'���<�eG�C����uj���b���ד��+EC�u�S㝎���>��08oI*��K2b���|q���u�M��%��fm>�]�����%�u�ha�"�w�U��GFq��+�-+T[0���r�B�yF�u�uA���ڄ�QuoJ.�=L�X��\�2�v�=��� ����;���(D޾�x��Tq�tT��^Gkv�֡ڂ"��h��57y�&E�K��]��ft�;���"G�e6�d�}o��%b��yx�wQ�h`+�7˭M�]�Vr�&��6�a�˵���悙K��׊�!m�U���j�"t�*K���	��Ũ���P$�1mL�b���Mgx��1Z<1����3[��b�,�{'_��ˠ{5�eJ�A]�GK�_\��� ��=[nb+��;����ۏ͝��_ov��@m/�a�<��չ�^��T��n��Ji�
=�gMv������ث�ݔS���༵-��C�r�`xYQM�MR��>������..g��-n��,��EX���U:D�1���U+�&ʋ��X�D{��б�+?�*�Va�b��#كl�?��K�nZʍ�(^���h�STQ��W1�y�Nv�W%s��c��-��m"�aZ;�Y�m����Y3O^�ىwiq�nL齻ky_΃��?�ߴ|H"�O|�<����O ��Q6QEk�ɮMh�*���b�c ���B����G.�TCs/.2SAr�IHQEEʷ3����4QIW#QEU�s5�1sF�ۘ)i�9�E͙KgG.C����O.T5r�0�Ӣ���.Z�%9�ȮE��9�j�8N�b�g�ʴ��ȸb���'7-��(�Idѣ�b���5�`<�yb��j��#F3��RF�Z�l����<�\*vq���E��]�<9������G"�͍��ִkK��M��Di�Y�T.ssE~s�g���Tm�T���E�@�a�t(�����EXF��l����|���#��S��}+�P����X�,�B�s ��q�9�kE]�fK��J叝i�>��iFsFJk��k���P�H���D�D�P$0M��-�)�d���$�?�-ЦQ���H�a�t(*mSD
T� �9.%Hͨ��v�ճ�n���r�7I�|o��%����p�3�O��ȇ�>���w��g�;:0��H�$�^H����̟Xk�3�܀�:a�/I)�K������y�ҧ��o�ۑ�mg��	w/ǃ��Ʀ��Ko����|޺�U�ȗ��] DqU3�.0�jW �R�����U��\9:Ϣoz�w���Ƿ�����hd�`�Mʀ��!�Wgq�׹a��E��U��wGUi��v��{anę�]"Α��>űnOkx��z:�L��M����<��n��f��ރ��l,2�ɟ��%r�)�?zD���D�:�p�~����z�.P��Wzu#a�Hx�k/q��j^1�&�����f���~��iҚ-}�,�L�U:��2�&�`%�j1�US�n�eqjPY�k�YR+�'l��9�r<6��)ee[����~�#"�_ld����\yc�<E��!ՙKe��� f���A^�p��nq��	AX-n]K����Tis�Ƿ<�B��	{���N2�N�VT��*ҦQ�׃����񻛢ʄ=�ӘY��(�t�}�����ۋ���}��ݓ!�U�ꮉ�K$S�����7+��DK�e���\�D���$�/q�M��k�J*Z�W��K��8���7u:wz��j��YG�*��r3%�s�t�R��v~�u��
D5=�=���sy����WՓ]kh��ݩk|�����4a6o��oi�s�$p�"�w̒TI�a-�J7�r�|,�۬�&�P�cc�����_AH\(�ZiS�e�7.]a�K� ~�f�ǓR�����E��0��u"_�ԹS>4�+#`
]2+x����'�jQU��¶��i]f0�3<p�fp��-@CL:>M"v����+��-����熷��y�r�<)C{c��Sd�[���s��}�J6�r�ٽ}1G(�_T�������
ggǭ̟o@�fq�?4�	ޫ���}ܣ��\�s?�B^lG��Jr�܅��+jі[���؅���x�N@+��u�{�':zk&�@��V��Y[�Mi0y��Q�˕�b�;4���D���@�t�^;J�9�و�|Uh_\Z�S�g�� Ǩc2v"�кJ���u��������N���t�.�W�m�J�(q�i ���}c������x�t�S�S����m��< gP���t���6�6���UQeP�Co4�Y��#+-����A�S����dظ�.Ì�9�� ��h�ʃ�����2�>��Kq�{��;���ByD<��DѺw�3����^���h���=*6��)m�U�z�����\��g؃r�]ɥ���� f%��;]s��kz��nt����/��d驺�v*�X�a��m�Õ�����Ƨ��-N�Q$��o���9cW-�jyP�9UM�}��׌�����mZ�y�d��{k���k�KPz���],�ܗu�9Y���U�V���U3�tPŌ��[�b���^[k�g!�YM j� s��y_��ݾ�>4�di�x[���;�3�]����3�:��!���f��wR�a�������g}���{hM�@
�E��	f�����+'��y���@��c����5ڼ�ޙ��KIVp�TXJ
���p�Ϲ��bvwFd'�����3z�r�R��u�-���>�{�?o����9!���ݏ�I�G@��g����2�˾EVfٳ�2�yX�[[���nym���nF��W{3�\1�̬N�� �����x�=۫/�K�е��H�_Q�F�C��F� ���O�|�7�9��<" �z�O,�$^մY3���;�tV.53E��S��;��^$���WH������>a]�ݹC�d遽!�J�=�љc�$���t�l-y�C�R +�k:��r �{s�P�N6��g�B��j�/e;rY�p���}n�O���J�|łF�6\���ӓ�<���C$;zּ��=&&��P��L��e��}v�]%�7�nb%�'��nK���+%�r�p��u���ݯwp҅_�S4oS��l����f�Dt�^iU����D���ޫAY�ؒ��Ս�\<��~�V���y�I�j6�^�ԉ�,)љ7F�?F!�'�iF��X��z�g���"�S6D��}*�4w�)�z�JNZ���K�g�Q�`� �n����õ�(��Wjӕ� �-�l^Eŋ6u'6��up������u�æ��n���pn�B S��]�1J�Ry���W	2w�r���E�;d��C�Wh�fOmW�;0��L��QjF�XJ�J;+�b6�ە^Ŏ���2�5�N���	�k�eW!��?��v����H�Y�j������Y�����wy�,�߼;�"^�e��[��qHǱ�my�
Wcn��#�훭|�+I���͜�F�I��*n|���M�YZ��f1�h����ns�vټ|��|�~���oر.�Jˮ~kd3��`�����MF������b\��/�;�r*��s��a�gG�!�uZ�,w,FN��7 L$"�=sQ�ů�eB��+b���M�ů�(�|?˼��}Y��\�߉�c�^����ܚc˲�J�[��bV��˸xc��1�[�I��ܹ���k��mҲ�q���u��I@6tV<@��8�r�^���6é��Dȋ�.�mȻ�Ž���n�P���¥_\7-2(u�	Y�� i���!E�`羛·] 4��P��^j�
$�4��ICHۂ������
��B��+H�;�g����ơ��Y'��ifhxZ���/�k���6�T9-E��H��0�>��aWǌ{�������f��{�{]$���>���.1�ɝ�+�B��4�t�v��g{�X_(����������� r���}p��j�<l5��<�@��7��s3�����6��ՎhZ����<�Ȍ�!g*f�
�Rk͊-�kV�j.���j��ɐxS5*�Fv�M��Q4;=�$s�B�9�W�ԧ�e�nyk����/��f� {閻�ΉzUt'SEN+L�J�ԭ��rZq���L�̿�g�gf��<��n"���Pi�Tz֙fVUtav1;�'��h$�l���T��Um�2�{�nhvC-z���X�[%�L�FqS�2��7.p��Լ�n���Q�����/ӿ+�7������"�e�/j��-����������j䭺V��%�%ʃj$��L�Z���3��Kv5��E��=a�9H��4K@�OG�7.\�wXr��?��UU=�)麔��,���Hm�,"��`)�F�}D�ڕ�<f�dP[��m�����G��pk*�<]=�Ɩ^�IN]�U݅T> ���+�Og.ɡJ�q͜Υk��i�<��R�����v�,;��
�ժ�ea<t�j��E��&�"��Z�tl��$ӧ��3�S�.����;iFe�/W)HKw�ڧ$�qr�|�+.��WZ���j�|m�;`1��o;���qW�T5�Y��*�lS��8p��yXyZG����U��U���� v.��<ǧ`VK�_j��Eޣ4�' V�a}�)����@>�a�K[b�)��T��R�w��v���y1+���;�8Ե�N�Ў��y�q��!��+��g*��1�.�������(Q���F��C���wX����n�&_����̨������}m�T|�e��0eݵ{0��P� ��3�P9`//=�78�5f�Or/9��h8���n�yY�@�O����b'Z6�:K���upn��jՊs��`=O �_7e�*���h`Z���^kp�T��ކ&���+�;�,\g8�W�X�[`4�G���.v���t���~ֶ5�e-!o�Jn��xXӗ/3&�t�h�i�qvUv1PWZ���u��^,Do����oY���i�>�]�v�v^�ʯ���Y��̦Q�=z��E���^՝���.����G�y:p,m�Լ�L_�Y'�_��5j�y]�����D]�v��fI��x�q�Ǒ��K)�F��� ��f�$�v)��䫸�y��z�&g��u�U��n�v�qWy�
��к@;�y�y��=Nf�O��g__Lu\Hژ�=C��BFm=w4f����+�5vQ�Q8�.��a�mi��j��O�R�`;��զ�:.Y�;��6.������an�7�u�=ͺ���%��Ce�Yv�p�������Q�#kwg���0L�I��7�H�ݵit�M�F�!��K���FL��\��w�A�B�;�~ʙ���ZT� %�l0Xђg$iY]������,��u1Kx�mȎh���S�o��)�p)�
�����1KiMm"��L�sb��&�a��}��
�}b���{���z,|3���sFD~��i�|��=�5�����_{v��.	˚��k�f� LC�u�	������<5��9C���lva|�Wm`=DTԸ�)�M��8q��nY�:Ka�Q�	٨Gv����r��3�̚d�W���;��k��xv�L��SAe��e%C��ώ�!�����s.x�,�|��,��9Xï���D�N��,��ag�f}�X�ԚJ�R6�=�Q3����-�D�[t���׶s!����v^Gb=��(w�F�f�
�͆�g����\�|�۷�]דӼ/o�*�.�O��zkOC��.lg[@��xR��Z�Kd�3���XLj�;���u5 �EE���YD�����?�ߤ��r�����0Ćy�k�wu����A�\��	(��G���ϼ�kT��S'*��z��&z��/F3gKT�Kp�Kd2흼Q���m��L94�]}݊v=*�I9�C�a���MrV��ۃҹ�e��M��<�3f2&�l͠�6��v|v��8��=���7$+(r0.V1=�p8�mh�U���,0�*}̟w,�,q�L�χ��Ve�ZM5����I���d�۽�Mf�}'p���ﯸ~Y�'��^��zA��&Gxnm��t��H~V(o�TD�eT�f=����	ۧ�����5�u֖��姸ۧ6���.lb�-�d�)�\z��2M��̈́��H�L���M�ջo��!��}�nE(�|�zҝ%���SCUֆ̂�l˳U�q�8H�Ɛ|�î��F���df�z��Ԫ-�knW7U�F�E��*��K�]MlŦq���]����P���:��B��Jq��*��:�C���Ԏ��z�����c����]0t�v�|��R:@��m ��yz!�s�{����G'��H4�a�ㆯ ��ͪ��|h�v�EC�;��fjД́�cm���r�>�S�إ����A:������:Nil,��t^�x��Ks1�ۥ4�M���*�LĪu��͈|ث�9I�ُ���|
?!�w2�������u���y�O��\�S��D���3fo<FB͛�W$��Β_�v
,�G��S�*&$��P��6�6T�����^*�q����yM6&�/wn�g"d"�E�Z}�����z���>�������������x�����}>�O���z������T���JU�{ ��ԝ�^��e���M����:�+�p�Ɉj��xld�$��V��E��hO��<ږ�tT��&�T�w�5�l˩�[�����Ap�2�{�q pJ�ci�S]nM��G�ɼo:R��0�}�0�+�v{��bPRT�@�{r�:�����ڛr���Z/���Oz���۱��a��m�Õt����Y��u7)�'4p�9|k�gB�)�o�B|��Ȁ	n�7�Ew˄��Ŵ��[K:�o�\���g%NĲ�N\�q�Q���kc�H�*Ivr�yRJ��M�ڻ�k��u����>"�'�f	���a�=�Y{487g1ǂY[\�C�^�=Put8�s�f[�_%gs��57;.�\�d(/�Ih�x���`�K�I�Bʶ���t>�����tK��
یj�I��-��)�W%�GJW�4���xS��7u�>�X����/��`c&�Ip�ox�U�b؉D-		�����[
����z�*�C�ha�pm̴������^�+p<w���V��i�޵��m��N�D��#�t쾾�aʹ�(��T��|ų6�b�j�i�e?	�3�qW,�Խ����r	��q	q��e�Uv�s�����$t��Q�]>��29�(��YT-�*_3v�%�mޤ�݇W��;(W�}���:nK�}�|�E��dM���{f��#���\\��e���B�v
Q�{mM�f�a�?�ݷ���`l⹻�Nq�\���V�\ܧ��d�ț�$�%p�\h��ɔ���Β��̒e� sG�M*�[7�ܡ�f��Ի�;�,���A��x�PGk�ΖKǭ�ﴕ˘�+M��Oz`P�s�F㫣���!�#�բ�X
 μ&i�.�L.�0]�������8gXj�Lq���{�t�KyJ�;Y �xd�E`5�P|�;sFw`Zb��;݂�LJk֜���ɾ�g���i��L�4]�<*���rr�}vEdT�J�Cc�6 �Ǝ�K\�w54�|)��uл��G#uƒ��Fﷃŵn;V�}s(�yWMo+u6��]1�U{ˑV�I�㎐Y��`�t�gOù-Y����ce�f��j��l0��͓'9�d��ww��������ҕ�����Н�K��a��1�B��2�g�e+���ǜ�4tHm�>ʮn�����ID`M�%��[su:�-�I�9�Z�A �E�li�[a��:��}�����p 2�ӽ"����.��gVܫCi�P�NTt��e���m8���n�n��/3�$/�ԫ1��Tp���(�ƧC�s�g�X�Wm�	�3j��:���6f���8	��ԹSz�ˈŰ%�z�S(m�f�C�^[�ݧ�ZK���:-䍮�܌wطF8�h���͊��~q��P�܊����[J��Q��cX��QZ�1�m�8���'FƼ�G7-�նڵ�*��s��V��V"��ˏ�*8U1˗&��b՝�Z'\��M�h�n��NӶ-m�Mj�����'�c��\�X�N1�m��4E�����d��جlj4Q�Ub�r�cF֊��64:��l�QQG-�hѧT�79��ڵ[b��F��Qc[	�j��Yأl��kN�m�4U�9ɼ� �i�F�#�Ǘ��yp������Ƨb�[c��1E���16�[W�9���jd�ƃE���[[h(�h娉m��b�\��/&�&����)�4[%gmh�G-T\�Ph�j�W��5���ȫbcE:u��(6s1y�ͭ��_�����K�C�3�4U�'ta�ՍҤ�@�,{4P��OY��D�k�Z��ʗ�
4��tR��Qw�eK�\�'U�X�9`�p�5nC������c>����W,x�a��Cs�U�&�q]�}w��ù���ًׁG�O��1�[������O@�|��RL6,	�̊���w��1�>s�Gl���{Ķ�oG%��۸1�]yPo�J�{�VY�r�go�iy�{k� �V�薋�*�#Ñ��wg�D�r���1G�볯/sE[L���+����p,,��q�1IL�����R�Wksdf��n.L<e� ��2� hg�͵�x�~�c�'����}�9��}����1`S�����ݮ��ik�^p|��nEή��n觪{����ލކ�ٜ�����t�Sz����8����l	:seY����,��IV�����U4�k���<��/��{�y�z��ˋb��a"�T��(R���=��u��X���h嵥��p}W�\��Ψ��6�݆3A^ƫ8V�B+m�b�r��ld�ۊ:���;`����9N��[\o�Vԫ��o%�0��ή\9�2c:s��Z��o�[�$��I]^���ppv���}׹n�f18A��f�y�ۓ�CÅ3�{a�h5��
�����ٙ��[t����uGq�]IW=��gm�Mu/�p|>k�}�ry>ν�M{:��ϭ�nV��]`��=�Z����{�mތ�����S��k�� 7*�=�L�x��C�Gٵ������#z1!�l�s�=�v�W=Z��b�x[a���Q�����3�姉�ܤ���bf{7�U��ێ�I.�+k�׉UM���T7m��!e���5���.�.}�=,��'Y+�GyU���І2��l��Ω��wS۬�]I�a-�G�sW��tm��Ł�׶q�3��jT��܍���4��!@_��FiJs�5�$zn򮑅�ھgv��sǻ7ɽUv�톩9�{fYB
��X8�D����²����Y�w�{�R]˭�3已O��[�C{����/�W~f1$�Vx���.�޽`M��e�Jk��mdr8#�@�M�X�!9}�b���S�j�!��m
�[�$� e"�wD\N*��v�4���Ȓ8�����k�v�G��uSҩ���i�|��R��(֡���ֱ:���*Uyp,W�js:��цe�`4�˿���w�,j\�^:�wn�K�4�p#6<�(4�����Jb	9�z�n��2X�/Һ�`>Y�\�"�����9#J���K�|e;u��j&	��:n)�Z��g�=��l��^��->���,[?��rՄ�狜׸ �dNSG��k�t�gLflY����;�wFg�~��g�g�.�h:h��8جq�@���f@s�˞!gH�/��%��2�ZdEr��p��l��p�Ҙ��Ԗ�����D����4[�.���8r���Ȼ>��7RQ\k�m25g��A6�L�l�cʽ���7��Nn��O<n�ٺ�9Mg�<����V�4T��n#:;�>�iѝd;�i���i�&�0*j,�XPK���������ۓ/�(_�мM�$\t�w�C��*�}Ms䞖t�lA��)���UJa��!�]NU��f��[�R�r��!:.�����%7!�Tf�;T[;���֔h��"�7'Vc�d����V�~-�v��]�6�q�۝R��˻��T���'p�Ʋ�|]��
ޜ7��o;na;5���[�_���Fv�m�3��5�:�����^4��-T ��0������dI֛��1����t���dR��n�z��[�94!c�+�����wkR�9�u�ܱ������+(��Õ�^�q$t�K\��������M�F���6����>���g0��ә�;����Ps�><��g]�g;+�K���;��=��B����6(�'��m�	-�e}�D==��a��xs.�^�;am�9�G�DjU3��5�V�xz�����3j�#v�jp�Av��Mɦ�>��9��x2\��.�J^;7��lة�!�f�Y��ۯW\0º�O��GL�p�\0���F.�:f�n��2V�H�����͡�ڸG6��讒n���ұ�Q�¢�~��]�`��{$�����P�鬖�G0��_�8�%m u2�^�:=G���f 7'��.6���v�1J�ZQ?��3��Yz�ޣ��\��Zr�/��h�ug
4k��5m
u�ŶnQOY=�]O��jX��&�Cu��:p����t�]1����"|@[(����I���X=�H8"�T��Cr�ɻ@j}����m��^#w�}u�I���<��X.}�H����`_�Ŧh٩�=ݏ���c� 5*�"�/P�˟]�έ�;$2�,tٴt՜��݆w�ɘ��l�n��4ΨP�����@���$�[�ц;_K���H1�6�E$0�����Dz�;�e�滏7T1����Ý���#w�,�crH�J��tI�^��ھU��2�ܱ�/D��g�'�K�r���S9c��5�dp�jFF�Y��K�о��+�m�"{v�m�u֥�Gn���oe]�~kD�@^%�{��R���+�k(6��쇝�������0�lݐ�B޽�y�d����V��{%w@�<9#�y{ז���N�!���F���y}��6����=�\l
��UxY��_�>;���#k+v�ȶ��'I��BƬ�f��̯d)m2��D���M�K	�B3�P�p~͒���/��Wx����X�;^��3��C�4�Bۛ&�� �Hk��T�_i9���]�R~Eߑ{An_c�H����K\gϨ����b!ldL7�程��.��+�U�t��`�w-�j+���ܝ]+��V�8�Z����&ͽ�[K�n���}�{�K�Ʀ��f�|�����|���n�Q��bK�%Tl����Z�|^S; �����3�kCD�1�s	/V(U�y�6)�b�Oe7M ��}��S��~/uc���=���+9ŋO"� �B��\s���<��bZ�(��,gj#��h嚈�ʢ���y9q�|��W�Vwm�KK6,t��s:�𦝨jׂ�{��i��v�(��^�{J}F�n��6;Q�a�'v�Nz���1�$��w�z���z�X��^������S羪jw0�-<��!-��M�9Gx�u��+u��~�'���gb����m5Q-|3^ᾜ�3�EbA�jo:�P�+/��mZ�V���P��;�^�3ڢ������Ӌk�kP��m�ً�z,��؃#v��wX�[��>L��?k2v��Yow[+�iĺRrJ'��m1ݒ6�� 5�V�LE`��[��������_%^h�J��tǠ�+�����jй�Xۼ����%;�T����k�sz%��1e7�>y~�]����J�w*K%	8�:G�mSG;��Сگn�y�;�z�'���#�+�ձ�_���M���/�՞i��X�%hc_<����U� ��3�-n?N��[�9���P�LR�!m�Ws fgҘWL�T�Eo̛�`V��|�)��Wb�B/�r|�Y�P�Zf�Y�S�⬈���l&"go��>��G�
A|��A�,��ۡ�I�7B�,��"���R�_)�{���n��%��M�q�i�J1=�g6��=�f�����{y;�b.=1d�������G[T ��8���v�iʹ������_��S�����f�]B|»GvZ�
�2b9��A7�{�0ϛ�������������W�b�n-f��ɼjY��oM��@dvZ��[��vs�x�k,p.}�,�|��n!�:�ӳ� ��e�'�s���X��4�U���p�@�3�ڠ�G�lXǅ����	� ٗ1�t�(ѻ�� ���_F�FbWV��6�5��9g*,��)i��B��H�����Y�ֽ{q
��Y}��[�jQ���~ފg=Q��g�V�nurͦ�������c�w�\��A��
��i�A>(���� ������x㾙�s�v�L��<����|�b�Hf�.1S4�u#e���yc�R{o���O�w_��,�����G�%2*�Y)�4�Þ����VmW9Z��+S66	s�F0���ʜ�����mMVׅ�.j)����W^��R��;v�d��6�l�B�;�}]��ߩ���������N�'��3�'�[.�Nt�ʱN�$f�3�y��[�v��$w]��"@�eA����fR�EVKSЛ��iQ�f�nn��{@0UW���~J��\�շ��1 ����95�i9Í.O@����OU39��֜���h���h�˨1G�7mX1�J����$"s�AZ�����-�WPҩC�tS���}zS�� ����m�#Ǖ����G�u��z�)��ؽ����b;MLl
�3�[s�T*�D�d"Ψg=����!�f��V���--ڛ;|�������;�X��C�NO�^�|��~Şی0�h��lx�,��'q�����T�f��V�cLs.�8-�l+n���;C�ػ�=�l�^y���9X��_�]
�58UmZ��]k���=vf+��=�[h徙����X�@Wua)Ƀi�PyK� �����g��5!'I��.�ǂ�#��V�R��so�y�´0���}ypijn]"􋕳	����8���_e�*P��KQ��Տ���Ù>��vDϣ?hA�:�d�T�t�P���1��^Ġ�'�7�|�;�OE�?H�����(Y�4��,�n7S�\��gA;�7��	�~��0�#�.iu�)K��)��/���>�l�͔��ػu�I��W�Ə��>�FH�t:���y~�4�Q�9�M=��ǌ�5*�:s��M�Q�gF����+���S�Ӓh��iիӔn�WE��������|��N�\L!qj!�يzjW�k����'H)R�����-dϭ[�jdd2F��~�7����.	�ZO$d~��X>E�Ҡ����j[5�z��m{�er�ʶ[-�E�;3��Q���Y�+�~-C�3���2^�	=y9=+0��({}��՛.H�ѿكR%k"���.w�T!�J�)D�
z���T��r��#}��IP�v���t���F��ˢ�W8�վ��`��v���e�E�ke�Δ�S�XW���eQ��U4��9��˺�z������>��վ��˝��b\j���p��
͐�ܕx����I���}B�C�$������=fG��-~�>���V_�A���9\�s�N���f�u�s�i�e�H?-�����熟\�ק�avUP�M��%19����~�����8zd��_I�a�Xӗ��,@e{!K{K�.�lA�ze�������{�;s>n�+s8��{���Ab?�
�}�;{�o����;n�t,Ӑ����-�������̂;É�'.�r����~�N�
tد^����]��W�]��8�4���&���c�a�̲klމ&�#CJX3ddq�D��*�
1�k�Oi�z�ˆ�
ڣ�_~s��u蹼u��]�r���m����B�x��=ݱX�*�q2�qw
���9~���f�`�����;��{޽����������_��v��H(���U�_������*( �,��������J3̋0,���0,��2���̋2��3"� L�0,4��"̫0,�3
�2��ʲ,�3 �0,ȳ
� L!*�0,ȳ�2����(�J�"̃0,���"�0,��,�3"�2�ȳ"�2�Ȱ�"̣0,ȳ�0,�� �(̋0,��̋2����0���"�0,��(�+2���"�a��C pi�	�f�`Y�f� �FdXf`Y�f�`Y�f�VaY�a��F|ȹ�fQ�`Y�f &�R`Y�fQ�eY�f� �F`XadY�f�aY�fU�`Y�a�	�fQ�dY�fU� �`Y�0�D�F`Y�f�eY�fE�aXaRdY�fQ�`dY�f�eeF`d@aH|�C*(C�C"�C
C
�C" C�H��  C  C��s� �UV UXa@eUa� !� !�U�UVK� !� !�U�V@UXa eUa�U�UV9����  C*�*�0�2C��"�å�����0����°ȰȰ�0����x�#��̋0,��̋0,³�+�K�?�_0c���*� �� �����������j��� 8o��a������������ ����ǳ���������~�}��A@q�������"
��H @U����b@�$���4���?��@�~��;���������~��a�П^�O��~��� �D U�PR�P"U@�UP�& ��P!IU%T	P�!@�ITdA	� @��P I@�@�A%UV�P�IT�~�����?��A� �@)K���=���?/����� �`~���}�̀P^���?w������?���O�������"=����֟pW�~H�>�?R|����Q U���!����G�A__�~c΄��*�'������/���O��`��A�I������8�p U����~��!���׀(������0_��|_���O�}{�?��I����ߑ �
�ϯ�������*��=|���}!��zz�Ӈ����ۃ�����@}���$��~�P_I�A��~i�?�x���������g'�{�_�D���Þ�AW_���=?����~i���
�2���#��%N� ���9�>�+�����P��*�H�D"!J�� R� ��R�
�J)P�T�"�*��EUHT$��
A ��*�U@PD�UA��.�����R$��QR��R�%J$�/�v5U*�EUT�AJD�j)**��DAI�%)JPQi�`T��B����UTJT�D$$v4J		%*��j��z ��l�   W��֭�C��m�
��-�U̺٣N�gwv� S�ÝCMS�w5��(j榹�Xn��Y�uж�6��+B�]�5�����j��Ұ�*��J*�� m��  k�=��
(=��@�
(P�0hP�C��B�zU���P��y=ܓ��N�gZwUM%Wv�iG;]5��Қ�t�Wg@�wcN���mY�*�e�U)P�Q �/    ���%�ڭf�n��:vNŻI��v�2��t4:u���ۍ�r�q�]-�t�����v��N�,�T�;��;��u�9�:�-�g�[.���5 ��
U"������   a�U�^��n�\滝:�[����ƭܖ�m�v��m�9Ҳ�i�U�uS$�Y�Tnf��V�F
��#CT�0f��[q��UV��IUJEP��  �y�Ֆ�[U�u�ګ�j��[9NdU�C�U�iε�۲cK�ts �*��6-eZ��n�:6�m��QպPD�HE*'`���  ,u�kQUN�Ѣ���)���Ѹݮ�k**��QW]���LT.��d����SCUn�jK��U�R��j��*���PPR���I�  ��� =�N�V�k�ʫN:6�[�(�V�4s��@h`�([h3  ҫP4 �� �t�T�TQU
P�UT��  < 42(� � Pɀ `  ,��֔6I� �#�::���  j0  5��� B)"�P  8  :����  2��  T�� ��� �[X 
Z�  j� Q� 41�H*F��T@��D�  �@ �  P�F  �`  0k Pւ�X  ��  @PLL
 �` =�S�)JR �Oh�JJT� hS�2A�@ �JR�  Si�Ң�L� �I&�eU&����[:��bQ��ocFSi��@�SX2� � _P\y�U�p*ʉJy>��� xx{��3���@BI�@$�̀���� �$�Ԁ��$I!!���������O�Cv�7h����B�V�K�hҚ½2f�j�yB1"cul��^M�M�.\
���6�)U�ۺ@�3R��f�Mde�����i'yZfK��RN�*7Kv�knj�$Wy�B[kX��7��yv��2��Ţ��L�Sla� 7L�9�-c�xeB�H�Qݪ����TT��Ų���/%�v�;�cU�F�#n� wY�b�ҢYNέ@+�<�
�YA_�Z4������P�z�#A�`�T�]��5�PJ�jV�^XV���d�^�t.j�j�+z���2PYĳX�dq�2̷�^[�kb؆+�b[���[U�c*Ex�����7Bʪ��9b������	;q��3H�Z����P8�s���OP��y�6V��U�ɘBk7.�,T襚�bL��p������b^��Hj��j�Z�!tu�(e�J�5�L�Y8��!-nٲ@Q�;mn�w�c�_�g3���l;t�n��@�x�� ��d�6���f"�m�pLm��9��&�i^h�
�e�uj��ph�[h�QsM�B
�oh�,/m�t��B'R� ���[����G1��1���[h*��ˁGV��T��y&嬭�5�Aji�V1+(*�.�)tۗ����Ve��f�a��vX��S$(�T�b�0�w��(�������Ƥh��Y�m�X5�^�Ҳ�Cf�^M£Ha�$��2�D���wQ#F�I���{In��g�Ze���-BV$�1���Za�̻�R*6X�rTiz
�S�l�qHm�mK�P�ʏ3nYe���,8
�,Z��nA68vf�����9{DGkh�-�:�"�����emG���,m��{�̸n(�W��c����F�=q�`f�}���q�l$�O/6�{�Z�_)��1�O��ZRڬ'.�)*���IS"i�	2���˸�P�ިo^��75@�CO)�w�6�Fi �ٍ\	L�裖��+o+3>f[��k/#wu��a���v�⽑1�b�,��>�p�� ["�-�ͧV��a�)�5��:"���3iZ?G����v�»��M�����3��o6�T�p]4��b`t�d����i�b�Y�,��nKT�wM����0��̭r=�Q1MECPی��U��ʸ]�b͗����-hFh������W��3(��b�S)b,����N��Z�;��B�1"����De�cLu4 �)�z%+�Z^�Xp�Թ$Y�M,ڗut�$U�FlfY��D	71җ��w�T�HLu;�z�)3T1���c�U�P
[���&}�v7!�1�GX�@���bȞS��!�/%������(�8�3pL�Ȭ[�U�S�)]aJ4D�+֭��1��aE+f�9%�%a���ʼ8Uݽ��wt%1�7K0��iD�M@ZT��k��hpbI�am�z)=�`<��z37 k*�A�bѹN�!VF�-T�:9��6��h
;B�b�nɳ۷�;K���@��\KmWa�F�n�?�
Ǜ��ֽ9�ۀlc1�b�Ŗ��O�8
[e����k�R����`Y��M�n�8�t\WQY�ӡ��+��Y u���YVwlb��fbǬR�#��*�T��-�d%�a��ql:��n�{�7c`ۥ��&)�07��-F)$��f��G�wri ﮗS҄�$2Y▬�/`�ݤ��%jԖT�X��m��ʗ�mZ��,�A&�
55�)T���ɔ�˶ȻW5օnh��M�Xa�qn�Q��%�ua��@��Y�U�͛``�z�+����?K�I�g~��B7@��
v��%㡜~��Q�@��߮�TBP'r�I�Zm5&�qSy{���gU+��)�D��3�S`OQu7R%mL���l���Ys(D�3-!�F᠕��pV̗T^̲�E�A:��r�+n�Z��pX�N��b�,�ǶƦw㰙p9A�����55�h���U��7Zyp�=��e��Z�#�ѽ��ۖt�oOۻ�<K7bإ�b�֨�T��!��OdN�iۗ���7��&ݬ�(��)�r<)
�ҕb�M��j�:���Dn뗔��[�V�%��4���a`�hB�bͫ��
����Y��nӵi�6N��2�ee�*�h�y(5��ȼ�o/��ۻ�`%.��@��2l�m+r�S�Vɴ�,t��UT��6ۅ���CkZl��&CX����`��:Wc눭	=σd;ɪ�\fM:�z'�D]��E(4��6)�-�Z(Հ"x��{�Rӑj�F��r�2K�1cj�5�E2+hf،��AwBZ:o!ұ<�ʼ�v����#K��7�x�[�&�n#�a���Z��@��[O,y+>#�^-�/Pν�GA��{�q6�Q��ӣSj�1?��Օv-��NL��LҠ~Z�������6Ы�CtD���N�!��{�,<� \��d�,��E]h6eUxQ@^ b5t/"�a�&�f�#b����Y$n�Qد��t�iI�s[o[��t��L5���V+
�Ә��0�CB�)f�S�ӫ�p})%u&���"�"Z.�XY���Ơ���ݍZr���z�')��J���{���7u-u�Q8��_j��iq�$�>�*�$X�c��L�6�.��3��u2�K�[ij��p���A�2Z�P�В�NkO3n�BSE�1T[�ͅ�[�.��Q��ݩN�Ӻ+�tڵ[gN�.D���U0���L���:ڵ��t��,�j��Y��:��K���T�b���	r��[���V��NʙQ�NŲr0�U;CS@̼�EK�Q��Et,]�n�+[I����ɯo䡗R�-��F,Oww�0���`͔P߈[��f�d��4�dG6���AnU�՘4 4m���PȊ*I���K;"�P�)�y�t��kf���=/U�@���x`���!y ׇ+F|��e��Jc.�ː�wz�b�V $����\DfI ���l�`�YF�[Y������7Qۋax�є*��&k��t�ԙn�M�
�V���w�K1��V4�F�aلhj�s� �̤��7jjy
P0�@�ёh4r�h��]c�K�����݊Z����rj���k)a�$ҕ�/@����UE��b�X�AhkS,���(«t�;0A���֪N�e�l;_Ja��!@�<.�K�W��Vbf��LT��U3x�;@#��o�� P�"hZa�vS�J�L�u�5��rB|YC�q5���[R�k/S wu,�^��&��4���9�gE�;fڧ��dԣW�j�X�x�ğ�gol$�
:���6.) �F�inY�٫i�i9�[8da�#b�G�{y.򵽰�����N�ԬN���F]nT�dc)��%͈��+�cL8��5�J�NZc�"Mk!b��ff�-��s%�F�4�4�����b7a���E ���:�Y�X���D[j�����%1G�v�i,;��=�stI��׮��C�Ѓ�j�%�����N
̆ӭfb zD���oٳ�E�k���i�������B*�%kRMչ��;[L1��0i]�m�ʵ���.C�BN}��,b)�~�34�9{� �� �M.娚��6(B�����pZ5xv*ܗt��*;��8�z���(��d�,�{Ǩbj�TV"�7�ڂ�A9�8�*�4I�x�:�1m��BQ��e7u�xq
q��H�e��B��#����)�J��b-m�dV���2��A	���R�J��v�7d���Wv)K�X3 ��{aY��(�dŅ,UXZ+T,�@+˽*]�ԋٺ�Y���;�T�jb��\Q6���f+L��{�Q����V�ut%`�ɱR��YP���n� ��eTL��
��A��m$*�՜�� 1|RR+�Ѩk�e�ֶcZì�f�*9H�J�c"DV�1��c`;T�E��l}y�fU�꭛i��b�cKef���9�i�:���4��;e-Q82�wxS.�T�L֡Lp�;ʖ��"h-z���eeu��bUx����U�Щ5����Mf��Մ�e�f^�w��&kQ�3(^:�R�L`gVU�XI@X�Tؔ�;���1��eL�V� �˵X��nF�K��Х��-咖Y����ch)O�2)�>��I�Zib��8*+�!�����S�LB�(̓Z�Z�W5j�����(�a�Tl'ra�񚍩[/@i�r8�-�b@�7�{,�PVmXOi�G�$9{j&�����%u*a�l�׃U6]�J���
��!RH��A���4���`�$�ٗ������D��o\��Z�;Cme�?!4Ax�ɱ`PdܥB7mP��n�V$hU�&B҇��j���41 ��d�y5�n]��T@�er�ěM���,#tV�Z½˷��y#�a�j��j`1m*�`� {	��FS� w��]E�K(���n�\�]�V�-̒,�N���nJ�� �r�M�X�kB#U�4m[8Pw5���j'��c����0+6�%���#�`c�^����,jW����,�)!*�ނ�ʨ�GA���d`e�̊����[��EaT�HXv���!�r��h�rkzq���7F]V�E5g�K�V%LX�KV�0�w�lޤ���۪w{R۵�S��t^b�&�Y�����%7a#�@��ɷ�V�(�Y��+�s@�;#�,�tLcR�����nAj��廡Vc&��wi
f��Rr�iz*?��%hͳ
W{n���[eM�������b���fakv��'zU��%���Zy-��X�0[J�q���v��Z���-�Df���"/q6�
G�jD9Wd�FP�E�5�]�͗iʂ��A�̚hZ���a�D;���{f�So��a�%�tMm�ۊ��+e-���X� ��1N�{���"��X�[JL�� �޼ڼ����Y��:{��pRį14��I���!�wv�\��j����$˺�r
�Sґ*Z�^�ض�+HU+ƒ�Ÿ鼠�f�=LiN�H�qI�Cf�X&��d���Y�ۘ�^�[�"Ś �ѫ!:�]���Hh�6�Ǯ���8���1��1�K*PU�步��7j��r��n��v�Tŷ)[��i�f�ˡ�����x�H�ך���r� �v�c�J5��uh��imJ�`X�V�oStr��-ݳ�P p�Mˍ�F�e[{6AR�XF���3u�����B��z��m��hXG 6৙�,w7jQ�v�Ea�[ b�z��g���n!K�c3�˖��y�'K�F���L�)�]+B����>f�WуTsGڕ �.G\̹��Bh��L�n��TLՀ:i�5�'��S>�8�T�*�Ŋ�Ҫؙъc'&eX��n`�e��e�	���nҖEOu�w����G�r��oI�,1T���S,�ŖXm����m?i4¨lZ�˔��wv��X�(SFB芏v�5�vr�×Fj��@ZMH"�M�bf�K�C�$4�/�#d^��M/ܴ(1I��t�
��(�ͺ�I��k������*
�]ފ(�D���k	F)aEX/2�Z�wkn(N�3E����P�@0 �lj�J�5�Sc2b��,ǩ�U �����`��d+ҥlz�[)����6�)le텶��p˚���r<GP����
-�,
����Kz�|�wX0������t��քb��1����oWdۡZ��@�����)��KQek���t�C]K��
e-ͼ�r��G+V�ͅ�h�&�(��
���Ϡz�5�,볥�_V������K�I�)`r�A�(�j���4�����bR��@�a�ٿ8��v�h������W�hM�B��$�u%A�v�:�od�)6[Lk0Iwdf7�;�E;�<��6�e�dk/4��b5�ɶ��J�n�˻��2ܤ┵�۴*�h��8f���x�U�h@����1���ʹڽԸ�Ѭ�1d�Y�v�<n�mج�ˏ#����ة����� �Z��4v��H���T,�3$�k���f�f��ǋ\`R�(�ێ������$�#)^��UQ�>v���Z\�a��7!��r��
����!�6e+JB�Uks N-���x�@Z��DN0vĭB�f��˥K-b�q̬��F<|Kڙ�⡭���0��b֦�:9��˦,���KiP߲-Si��*ݫ��'�f;˦JۀUũ6M9`�����"/D�O4F3)XU2j�`;͡��1�0�Q]��
�V�!�� "�~uia+iQph��x�̉�7eU�7Z�h�3�M������]FhDm�,�65��L��{���f�ڹbۥ�1Ej���f�+(Қ�s끍0GD3�
���:B��(c�5��S�y�@�8r�(R��nAh����g�V*96�D�t+mK��e\��r]�����m�4�r�-{B]:HPf�U�"z\�VN�L������%��5�0����[͗W0�c*ŀ+qɆ�3���G&���[R����e-�����E�+llU���J[�p�4�c�H�تS	Y����h���CR؍�P��5� U�"����H��;n��GfM5��6S4�QL	�+�KU���
�-M�j�Q�2�&Ƃd�"�R���0�k�a���X�F��^�s�Yn��k�����)�^n�vCڤP��(�ڛ ��G�6�j��
(h9wG+V���Ⱥ4�g1:j�ʄ����a�2��Yvb��m�f��v2n(�,��J,1�
��mۡ�&_�W.��+��V5rW��U�����`�w:�i�V��,N��P(m��ik<a_2���7�9���.�3F������!zGm� �/W̚M]�9���;�U��ӫ������9�<h��ng��㫫Vvmn�f
p��iX�h+_M4zcr���wKD k�MF��pĴ����8@w�Ý-QH�x:X��}��Ze���gK��t�J�o+#g{5ӫ�\���e\씛Ł$���/�Jj*j'
��P��>�5����t~���Ml�/��(���^\��a����n�h.�Q�o9(GՔh8�^S}O0M;��>�V� �S�Ҽ����V���
���u���WR�,��Z�=�.�h��c�R�����Mon"R�q��8���M%]�v�����0��<[x��B���"[�fr7��a˭�}�ЛP��:Á�%.��l�ū�O�o '*y�+E��pkz�`�6$��mf���BZ��O^�/�VeM���j��:���4'�#<c;�h+u:���MR�E0��mtő��!����9�׻����Z�����Ywgn=�{|#�ݝ��������ѼU��t�ŭ�̚չgg.;bc�3�#��a�11IY�{�k��BƵo= f���J�ġ@Jb#��M�e�:��\*fаu�)�I5yV�̹�[t�M@n��C.�&g�}&�H� ˕܀���]�7�o��9Kq��n���ZEN�,]��k�v%]���jv�
�y�QV�R9"���6G�X5�d�pl�*�8t��;����K���+6#}�C�����:��M�{j3�ڛ���	�{�q�y%��n��q��Q�7��Q��ۚ(N��p�m�����wQ�s�[��-Y,�اu��#'4��X�m����w`� ܕ�$��5ŵ&	���,�L�g=cub��}\�͸z.$�n�9�2�jG�MC��}��v��� �z�1���&�jYݺ�x�.�v�hJ�ן;�x��*�ohuz�-[
Bvq�1]�׼uS�k%�tC̠oRJ�:bn��^0#R�wuӏm�̮�mTvh�h�ô�i��ڗ֧e%f�����
����NZ��'�{�;���tq�����J�оl��/�>�]%��K��x:޺���N4Rے����.���{;�c&�o�_.3V�Kg�>z��սg6(B�I�	L�o�Y}7x`��,1��2�d��]6�-��뵷��Bb:y��MW�`��J����8���ܮ�غ��[�G�b��y��MЊ���A����*���0ɴ9�A��ЩӼL�ˮ��q��Ϣu�3��CS\|Z-���1È�oo5ƕ�|�f͹(���b�f^Ǖ��]h;�$�=���n=+W_nS���PW�Ĩ��}�3N���8~�3Q7����m���;w�����l��φ�er��z�P������k�w[��(h�RU�|!q�BU̘36ξ�6ے��h▬��O�/sz�sZ�M�E����v7h6n��g'�T50�4[��i�W Cs)n7�R�i]%���JS���,����{���z����û}���(Mt���D�����hf�
�Q�c���7�ͤ�^W[�}�']Ir�F�r�-�emgc���9]>��6�BC�_S�Ӫy!��7����u��UK���yN��x�Ý˅�w�an��,uΓ��C+�M&a�-�7V���Q�1k���S�A���`iҽ����@���b�4	±�� �]�ڳ!R�Y3{��{��ecf.��]<8��8�Y+�F��(���5�cs�A.��.����=ㄌ:С�]��l�䈴�f��d����Z�SoI׊�;��.�'�Vp�x��v�y6��n�V�%W�����-�殥RP���h�����K�փ�j\���i+X�"2��<m�����P�W�۱6�U�L�ģ]"��t*��B5�ؐȰ�w7EXE�#�R���%q-X�/�j�ʨc�k�o�đFr�+cn���'n�i۳���gzg���Ū��d���Y�s;Ri��^*�J�P�G7{[h^�h,6��x�:�S�,[�F]7�
X�ǲ�x��K��d3�a� �����rQ�hr�*I|���T�[7�w�����+m��0�����w��z��N�C���m=�g%���Xx���;-��t��lwU=��o�J�jՙLB�K�Z�Zu�*���-�$���(d5drȚ̖��o�n�r�!�°T�"j�߄	F�O��5��s�˨DV(N�ڝ�j0��n�'j
:�-w(�W	��iJ��P��c:�&V8�]%Y�ଧ��՜�;��n���S�B�m�1:C(j�t��z�zZ��vշ�Q�=Vΐ#���k�#�ީv�ve3�3�k5�J�]�8ɋrh�d�i����i�D����r�)�U��,l��P9�&Q;2���2�ݴ[Y�\@�=7{x���\�F��K��jJ3����Y3~Ԭ�3���;�-�����Z�!R��-=n�6S���Y�O��t`}J�na7���Xr�lC�P�>y��g�#}F0�ֱ�I�ʃGR�b(�<�n�|4�8nvU�7(�i�+{�<�``Yj��<���8�ÿm�T YZ.�Ջ<�u�"U2�.�bywS��OD<�k�GY�45���m1�trAYy���Jj ���fT�c�y�A�qT�������{v���K��>���^���bv$ۉ��lۃ-m䏺�3MsQ�r�Y������lQս��"Gv�ݷ;���R���K4ӜP��b�s\=b2ri`���աrΰ{���%-���z^��X6�`�j�c�u�,b"��X���{P}A)�]u]me�z�Su���W"
Z�):�g�3ZܴQ�B^Ff뜕��yd�O붛���Q%sśW�z\�ѻ��0�]ZF-�2�-�vZ*=h��Ηqߚ[New�	��e� ���9ڱ�h�M�"��6V�7sz��}7���W#/�":`epRӓ���&�C�عht�>��V�kl2U��y�e���e�����Z5��α��rޱ�
�ȅ�G�7��� �&뻩dyYn���8hS-os%b��_��p8됖Բ7u�έ��bwj��v���Z�u����O{s&n�2�I�U��7�b[�5�c�^�S�O[��� ��ۭj���	3;ZU�5)��|��T�>�}��ԴR0��x_[W��9Wp��
�Y�d�}��+�5+oG(X��v�-��:�h�#W��cR����1��F��c�^/�5�k&Y3����ud���f,��y�V �#���T9�1BAD�0�N�k�`�ц��ኑ����hۡ"�J�hh�rq{R��xo�j�\%IO�j\ �sq�"ޫS���!�y���x±�F��T�ح�}��	8V�7�Ҫ��\�N�gU�����z��t�\XB��&L�R��ͅچ��@# w}xơ���Y�PJ�^[�N�2��w��HS���*��I�v�fbu˪R������D���ay�;T[v�ާ��ߘ��Y�(>N������Z�d�����OoC7ۘ^���Q6ur���2ngb���#�x���DV%���=(	O�a��m6s�g;�J��V�m2�w�份��]�8�m\t[��*�aV#a}6�hc�:L$�Sւ�{Δ�M8�i�v9�U�3 �.S���0ۙ��vq�Y��� ��E�4:��U,{N���L6;�y��t�'�>e�"p�ZBֵ��R��@����'T�#��pbѿy���K�ԝ9ۙ,����׊���Aݚ�;r�dvJ�kM�ϛF�`!���v�*��eX�ع��*�U���#��G�ـEV��v�dnDҠ��j�,����|sw�n��s��.���\��љMe.ѣ��A4Lkon�\js�L�&����NΓ.���&����:�O�)ګ;@�HY��2xc�4W�J�+�^7o,��l|�AǛg�f-����+���Ի;@1v���^6am�Z�+�`T���>C��$���ܐ��mK�Í�҇bT�)r����k�a�l#GV�dm��ط��c�.k��+P�aY��^��vm�,���1w9��n%�L����z�a�-�}��3����g�8���o�v��٭XE[]ݖ]�8��<ɏ�m��M�rކ6\4��%�(̨36ȎRk-XV���U�����Mf�ޢݨ��4`ep�#,�}r($�� �{m�Z;�{�wO�޵�vڼ�Jg@�ۖ�WP�6uk�\��iv�]�N�
'/A�'��K��60�*�7($�t��{�&,.��0��$� T����VB��n�ތ��E_Wu��&lx� a?gm�W}��'+�^D���j��K�����ͳ���������ݎK�Ų��X�'%]h&���i>6���xwwA`s�f�n)A�����g��~�5kW���+G���k�Ft��9�{y{;@�M�zY"�	�ٶ��
=�k%u�r�އ���F��Fq��JǢi;� u 4h'%�Z��J����cj�<R]ٺ����f��E¸�oE�<�Yt*�.J�뿭ҭ����h��a�˼$bs6�2�-�M䕆G]�&�wR!������ͅ�"}��Ck�E���,�y��}���}�i���:��%���*u���I�u��)u�mI�ծ��|Ɯ�uX�*�MK�<
�bW��"�I���6i�{٫2e��7nc6�G#��g%[T��aL"�hbK��E�6��PU1�.���
���1���k\��Y��V��q����J[ab|��.۔�}Eꋃ۠n��T̯h��Y,;��W��s��)Jv�[7�j4w[�n����t�E��zcY(�}�����hp�(�� ؒ�e��Z�?h�L���W��b }x���`㮳��7VN&�_,aRnGj؆�]M͚�8Du��Ky0���v����`��`dMYN�nٛj��f'd��r^�ڛ��լv�CSw�'���b��me�{ѫ��3��_���n��h�ER܌��rXK{�+L�<�/�V�h+��{�澗�L걖��J�^䔜�G8]20e��u�e��ǃ��������XW�i��Pw�h�9Xp�P*?��X9tڗcE0h�[w�;�Jb�珹s�K+�E���jub[��e+����(v���'F�o9��`vE7	�iБFV�t�5}�"A�\4�G%1y��2�u�H���rv�ve-X��:>{�͘�|Ǎ����wG
{|�ܷ+M� .1usU=�.˖��XC���f��R=�=��:�W`}��Hy��F�r�{@�}j7��O�:��A��VbY�)^=KQ��ǞNX��ܪ�WN�q�@��]-=��q�ʌ���t�	ۜ���p�TC�P/O=+��9��|Z����✩�7����v�*UtP}���;Wp��J�h���)���u�z�#;)V���5�cU[�֟1���9A��^o�]�����R�V<f!r�M�:>5�����dZ�9o�3�.X����e��e���6��*_i�jw�a05���[����}ع0{7�U���;H��z�l����C�؞F�ⷺ�T�����(��kzt+������Gh�	0�}nU�6��\(i�^�-�H�vU꾮�s�V�pNwJ�H�E��^�#|��6�`�ڭQ|u�z��qU��0{�]�H1�.+B̮�]��yi�2�`���&ܨ	;_2�G�� �Qk�WڻXB蟒��Ot�Y��'M�s��f0�3�!����ʹM���oA��t���Y�C�W�1<S,���(b�ϸ�i.��>ݨ�����J�n7�e��X��.�j���x�݉;����Xz\6n�awP2�<���Z��{�/Y�-ͅ+E�=\��'5�[Z�"��]�Uw����GX�a�֥�P�5�V��J�Nu���7`�*jԫp��W*9ۄ�:�-�\/���.r�:��]��*o+�03dn��؜+6�3�͆�ȱ��]^LU��p�:��K�u���j�Mp�8�X=o�)�w ���k�y�mKD̝�n�*�W�3�����ӻ`;��H�.&n�Aӎ�z�w^[��C�Z�a5��/�|[���D��[�qLI�pHs-q���1��X��U	Ze�&��n�Z�j�������Z�VA3G����5����r�l��uv�uG-av.bE�S*pX��+��@-�1�ޝ���f,ܙ�wWb;k�Y��;^�L�ih�j�qu'f�0K��,<|̛МUr�\�ӷ ��]��fkqs��˴:��R���K�S�I`��;��b�BY
�]k*<��+Q�2�R��M��w|	�K�mQ}�mΌ���o5��2�p�\���q�J63�\oYܽ�/��7�k�,U�3!]��X[��\P�G�n����ap��u|�W>��L�=[@I[��q�Y�+GXbf������i�{I��ٓ�X�fƌ�n�X�]�/��M*z�`�lu+��.�.^WI{i5o{W'%���}��l����%��8{�۔plsdx�t�Ȅ׫��z�{�($~oxY�_[��X�����.�q���[:��x�����%�,�t��*��7�>뗓���������N�	�++.�kw��{����Qi��ƺ��Z_Go{A��f��	TNd��kr��P.���۽�Μ^P���k!c�ή8!k;����#������<I�0kљ�v�t�rT�Z��Gop=�K��9lW���L.Y�>��rQn���Nw�qF����x�{���{����D�t+�����h��3TBI�
���X�釞8�/:�9��' �O����@R1-��[������QOg)p�=�R��n��6��i\��9��as�y���P��c\���GiR��؝��AP:l���O7�u�X�O���.��>��I���Q��8�wΕ��G�]����4���X�ns��i��+��>�4x���&��,E�;�x�p޼V�!�js4	��H��G8����j[4��r�N]3F�]<�*Pa����Z��W�oiuV��a�R�R[�%Y����[�k	I��,vC;��)>Ҁ�
�����i<tiC�Mr�ag>��� �­�k�(��N�d�=]C9v`�uV��=��7aR�-l\�E҉�f;�v�:�Ո�;�rcp;�
 ��}�SW�>|�ea0v5�㧜�:���l�,�&�PW�o�yK��//lJJ���I�Z:�[X��7���{�B8�V��+��$��2��b�R�,Ř�*��cOT�ώ�y��Y[vQ��2i��������Z�(��W����8��W𲕅z�I^bʋt��p,�����GTDD�,nS�H��ؖ�Wi����Q�c4r>WIM=�d��^K�#�	_�P979��j+��F�����5�Ŧw-	SJʃ �%���e[�B�!�R��v���춨п��Դ�ޱ�)�W��[���˸s2��=+Fe'��/'iC�Q��(kflӴ��MU����Tqʺ�`[����"EY�w��R���Wi*�g'u�p�3T�.=㙙Q�����u��y� Ζ�%l�(i�f؝�C�V[��Zr��X��b�3�8C�z:Y�љh���Ŋ�4I�����1f:r�F�q�T���
͌���5
�}B������Y�d��oqqƌʝ2��yQ^�E<�!4)V���c9�nT���5��@/�j&�4-�)�7m^�v���V!JG�uv�f�ǫj�]=�+_7Q5�38�PR�ق�ȫt �m,����+@�X:K�c/�\YM�Ùs3@�( ]�ע��uj���c�hl�����ĹCe��|�7W�����ʔ�X8���\z+���>�]wX�8�Ձ��u�y��ǫ&htĀ��}�Y.�m��qU�.����mX�Y�w4��.Q�s��� �����+�aJfMs�4��Q�� P�ek����k7�̅���i�s:E6���f\��q�@CX
�x0IҖc5wqb����c]A"z������*R:BBV�"�ok��������.�3g]�K����-�OZUx*�;�����t<g5]5�6�;�
�l��[�Բ���}x�ͳY ��hd�Gu�Si;]ǖύg]y�#�HV�����'{ܞM�[]s�*� 5)WJ���\��ɔ�J4t���#��r]��_ku���,��\�=����ѽ;�vz�Z[Y��5��[d�ާ�S�ܵPE��>�L]��Y9��^V���稢��uMڑ ��nhM�uի8��mwi������%k��ιaf�0�wn��:���xw?���)�[@5�zxXˌ7qC����u��<ܩ������jMg �[$�u��vs{�
�O�im�1��⎝�xBO�0,�u�B<��Zg+(l|!g�����h�_C�\n���u�_M�xh��e�vDb�b ��P=N�Sc�DL����՝�Mk�V��X*NW�%Yu1�����
��c�]滕s�ՠ=S���t��#��4�l{�__;G�Y����[\Ȋ*�
�B���o�8ɱ�]O��Q&WY�:��ot��I>7�������A�u��j�g�z�^�Ւ��P9CU�hWU��e*�Y��.�U���]y�:v�rיm뾼����('33ml�4�4���m�y6�������,^n��p�y��V�S���Z�{ݡqm�h0%�wąԳG6�lյ�F:����nS�r�[}Ne=�[�W�y>Ү����]�DMΘ��I4�4k5sC^t#p�[8:��i���9�l��ιZ�tc�N�X5z2)�Wep�$e3+R\1-<1�����:��jBՃ���0@
_S�"�?21bg2�P�e�t	�Y�)S�Q�ېVqkx4P�ٙI�A��ܬ��|�S�d�R�̴��Un`��i,����m.YV7ӑ���:�rN���s.�K7S�p�yAe��N�5�+oY�
�C���Ul�պUewN�p]���0҅�V.`���o$:ns����ww`��b���b��A���ӫX̵���_1�4�]�-	-�9`S����Y��	�o��V4#�|!���<՗x�ȭ�M��Y5)b�t�����g� �c2��i���I�wW��I���uB���ɉ��Pٹx�vr�876�t��ⶎb��K2ґi��dk��b�ʲ+[A�j�1T�6��rzOQ|��ۧYN�F�@����.b_my'k0n!�iXv��r�N�\%�Y��>8%m:�b��VՀ�Tc�m=�����;w���]B)�����z��1%܎�
琪���Q����n����۽��ԮHЦb��\�cP:��0O���U��|�/��vV�@1�fLY:��(��IXB���x�S�8�O���Wk��ط�ec:�g�nM9�C���0�\+���3��+s�]�����7�kYs�v�5^���M}������4PX,���]�e�ƕ�nKI�/J�e,����-�U��񥗔����\��1��vV�`�AG���2��"����r���9��x�2��[!2�ol��=�C{�.8���X�{WM7+85�;:��S�Z-�^��y�+6MUۗ��+�)�����YXr�D�:�}�8w����)�Q(�4�.0�N�3Cf5Rc5�-́���Ҡz���4�1V'��M�b}����9u�û�IFhQ{�	D���HZ4l���R�h/�
=��V۶��à��vsB��j[�&O���.<5w:-��P��7@ޥN�����_L��P�.�n�!�Ld}��%.wH^�Z�����ހRْ�Rfi �� �qQ)2�R���sy��E��ݺ�ݭec�����႞���L�H����\���g��݄�'�b�6Yڌ�/�&���9�Ms�U�v����R6���/���-)y���� [��V"Vo��������ݗSn�*4�Wu1�)��Kn�q�F�m�F�ӲO(�cJ�J�p�����\�RE����/���;��_e�ib�z�Ō�[Ռ�YԜ7��]�ٽ�
yOj��Uݲ��m�-t���k�]j��R����ï%�F!�ar:k�gf7}����`���\�FT�\�*VkCx*졶�&|yJ��m9ث��_Mg�[�,�GՕ&��� io>WoXMn6���
uff�Y3�lcgM�#ٶ�P	�S
�;y��ӄH�39&K]Cz�n��g�L�b��.�C�k�`���'0���m+�w� l�Ø�Q��4J�ж.����e�7l��!҇Bne"-k�0��*9�n�=�w(��Rf��;��};r�Z�]��է��sj3�=�9��k�5`u[{���P���RB���X:�V�x�Q�ia�w�k�;���:wfs��.� �6m\|��i�������
��Pyl�h�W���0�)��ӝ��*L��%[�h�oyet%槫����`�$�
��%)����gf̹	Z�n�K+FuU�Mش4�ţgqQ��@�jQ��L=j�mX�e	�L�@IR�D,�n�����%�W1EL/�J$�Ia̾U1�.+�Etg3��m��Z�d\���[m�;��ꭥ���Յ
�Y]hٴ��:�C՗�2���_&i�3�B���tJ��`P�{�ɧd={QJ���Zojq�6��O���yr��av��h�Vj��AU�gu�ޜ��˙�V����������ka���z�cB�ݴ��@9Br;w�G�B��dc�pw%Yώ
�wf]����Aw�+61k��R�{c����2��Go)��x4�`Ơp_*	�{EL��;�J�Z������:N�{�;c�Z�,D�V��8ҹhB�k5��m�����B\zs�q��V]��Kl�A��G�EͲ�ժ�7��k)<� ǜqg�z���C���[}��n�T��;v���uۃr���Պ��L�9��V�}�lL�K�C)-��$h4$�!�	im9r���x�4���h��]�ʽ��j���	ێ�9ma��(��4�6��`j�Kd�Qز`��fEŚ��ڝrrJ��"��G9�Pc�jp��!P����ݙ�؀s��Ti���6e�h�b��6Xm��õgP4����U�U�:����gd�����|�ҫC�&��|]�\Gg+2n[��G�B��|�uՖ��q	�.젋DœR��b��xVl����l�Wq��:]�d8�.�uW�bU�P�����L��V�f�w[u5�O3����9���t�����3EV+3m6\T�]��j4�Mr{-���CL
��������rU|�3��Wx/����S�&��.x��o.36��,g|�����ګkF�a�Ȯ�CFG�0���Kqj8��]N�trQ1�m�����B[���ş0Ѿ�~�j��R:�	�D�<3O*����kDۀw�;�:�9���_k*�2�uԺJ���wx6�:�(=<OǏk*쪽�M�:���Q�g�\Ë�M��H
}ˀ��ת�t��z������Ύg>�O{R���Q�KM�vx�j��ڧ4�t*�{EjTu`!��o؉�Ë�
��([<-�ut����Gi.��NF]�zj�/�',�v5g�#0[i.	��,**,@�)F�5����7ob�4��.�}��� �R\b�:��\"�jD�����|�����Oc�8�֚�r\��`�hp�C��G�I�r�oR�{MاN �|K��7��������ېN�z�Օ݋b��$%��U�uZ��::Y���ͭz��{{]��
Ϟ�1t� r����f-t���γ]qLW�^�B�6 S�;܅�7$H���NU�d��� �j�ps�%ceb�h=Y�m���j��%��"٩R�U�%����5�P��3�\��X���#���8��̴�̝�΍m/��|������H|��Z9f������{��u:`�7Y���m��OD�0X]��1����{(�<��f<�9�vW黉���;ї�y�����X�L�1�=�p�>V���@�kl_!Jp����-wB3�c��mqKE���.��mҼ�ij��9U�;��R�S����#�����>b��N��sfJ3��K!��]4�L�:����s1��+� f�1S�U�ׄ��IL2�n8��"3]�t�bP=�� ռ��.Z%wd�n�p�`�.�˶�ų�,�$�j��bn��P�%]A	��gs������FzP�AT�����<�B���SGl��K�ڂ��C��T�b�CS��,kMA	�K�+���Χ��[An�2M}si�l����Ÿ�[���8��sk/R��T�m�ċz�e���6��]��i���s1�����/��'8r�b��ٰA�Z�dV)���0��A��e�}]�ؾ��8G�d`Ò���Vu)	æ�&��R���(p\u�ci�'�7/viv%'�T��K��v�j���47L7WY��
8�(^A۪ؼ}��*���,�=v��#Q=����]䝣JOA�v��C�.b�k��7��DG�0;+��w��E#����z��n�WV6�H���aX<����[pӔ�6�d��yIIBeY�ﶀ`��n�p��])Nm���uf�lu�k��[[0�TM���u���̫H��*�v���ȟV\\���x��#r����'��w*Ҽ:9'B.���]��:36�S���,vIMu-m�pd�w��5��Ҕ͕jq���2.Zk37pY
��Y-�GDiރJ�s��%ڗT��Y��P�[5�FV��*O
�
�LTd��L�ÜMgR�Ω�Ɏ�2WNe�'2m�Eԝ�8��-�-���T�M�7X�էyX��K�� �Z�ˏk��ۤ�,a��X�Q�aV����r��S3�2�iy�A��A�+�:"̤뾼�V�Y�ujTn�c����\��^���Δ$�̣���g7�-%.z'֏=G&S�q5k��e�L��Z��V(�*���λ7tSs(bZ�����ފy�9o��>���˪W%�:����X���u_c�(�;p�E��#�<&	�F�:��Խ�I�:��[���	8�qw�{�(��]Z���ye��L�Y	ح�d�!wu�����Nֽ=p���*Uյ������G��c����Ƴ��B����Sl���$5�]��쳫jؕ���vT�	�����+ʍַ�v#�U�Ǥ`=�l �V��@�uPR�-Ԥk8��6��Θ>�kuK���E�d�3O�`'�b�ٵ&j��(󃊻����W���-̹Oh�r�{�0:r�*����7�����Y��-�kVI�R��1 ��]�V�<pR�V��FЈV��(�3{+��y!�]�.�!*�g05fJ�`D��,k�0%��*u�Ζ�Q�F,�ݺ���^�5!7�����i5�z��'y�u�(҃%�6:u��������ƨXz�A�4c��W��Z���M����0�V�{s3g&�8�J�Q���}���d���w�Mt懷:�vf��O��,cz�-F�G%�Dj��U�����Z�f�E�ZnA����P=���Z�K=��� !	%�yv�8߹�k����0�>�:�S]�7�s�SF60t}@�8J*�f�Ss/uCF�p�"������@�v��h�k�Dfk���w^��Y��]nd�?b=rsxw|�M�0��߽�n�4H��إ�|ok"3�%O��͗0��+cx��J�,�`b�l�Q�����d`�`ј �Ӗ6+�GXb��uLNo9�o���̉՝	�7Z��J��YKV�[4g�{��=���w	h!ʁ�t��a���k�ƪQ#o:rW"'�v��K����R�R=��b��&'�Y�����O���7�4�	VU���+��|(��O2Q����6*�����״z�[ـ�HX��hy��۾[�:�飋��9�taB%N�=��1�:ZD<���9���D_.Q,ꚕ�#�t��t�Fv5���B��+����g�7�x��3i���4� �C��(j]|��(]osWR��x-��$�-_B��\ݫ��6����{���4��m����k15s=@�V�����n
��5�[x�v�p��+�i�ǘ�~݂�n1�ѳ
�� ֆ�4�i����}�Hw	�;��Y�6hr�0T�h��'/UZĒ�����mvz`BG��Avĺf��(fl��-NR�O����w����7M L+�{�>q�N��G���8���D-�0�a�U��N����fL�JhV�X9E�ݼ�W��m�ʃJ)[}��jE��U��j��-L�V�E(�J���(Vʸŕ%��*�QQR��T�ar��6��E�VT�ZAB�m��Q��e���"�V�e)TZ��Ubԕ
�����T�+�\F��(��
�R�KQ��]P�.�MS-P�h�U�Xc��&6���aKF��ˆD�����Y.[�
\���F�E
��N8YB���Œ[��(�[X��m�Zŀ����R�[+R�TJ�Z�k[eF��Uj֩Z�e�QTAQ�J�*(�hV�2�-Db�[-h��kj��B�#fam(%)Z�Ѣ��0�EF%�)EBؖ��*5�R�*V��E���°���֤�J[Kh��M5�"akm�Q�VT(��Jʬ`�AV-�ih֊#�h�b�(���[j��V,Q��E���J1�k5�9mZ-��Ѷ����PA�o�]��[ٯ��N<&K���WO��XM�鑺��v=�v(�!��^����<�Xޜ��P*�2x;Y��@��Z�p5Ug�u�t�)
�臘� �7��+q�6+��e��\ ��p��Y���'�S��:���޾��w���=Y�ETk��+��5�<����{�X��E%��t޴�#�|�^���@��r{wtE��L�9rV�#E@��T^Wʮq��Y��a{w�!ZX^x�-9��ͯX} �
؛�7{:¿v#ei�F�0��:�E$; ���gp�Ǘ�?8��P�ҁ���Wo:ێ��G�<���3�Q�����Rҭ�w�Ԏjnn�5����<�ᯱH���@Q�L�/4�_�WY��}�Y�PuC�!���&��~�,���[�c<�[f��uHb63�2a�g3a�����.��L�-��HV���\�Î��!NԳ��Qɘ��n�ʈ�+ْ�H��e.v��QJ��ܮ�w��֬S98T�onX�oI㶧E
&�o�޻���X�d�00����Ɛ��׽����x1�
�r�H���:j�����~d>2��*��#��-��yT�53�F�ԡ۔�i�LI$)�u�𭞷ѳ��*�ّ�ںg��A��}���B�BÍ�WW:���*TN���2~��U6�� � :m�*���#:�]�s�|�|�ՌN�h�;���n(�p��S�P�$U��G��yS+,J�p:���7�T�E���)���W�u.���3��>O>������gl���4"]�����^%��vb3\f&�y[TV�ڭ���y�̥p�=�;���O��h�p�W���u������7u�[s���Vrwo~������рܫ:LpweB�$lj�i{(_<�ʧ���}Xl��*s����{�Z3�V�ChA�"� 6el����xr	H�������*��P�� �dr��yX,fg�MkR��9�Z ���*E#!I҇c��*w@L�,6g�tqqnku��J�#~}���Ý�G��1���BcMx�zr�4���!��?jX�;vk��e-�-������.-x�5�tԊ}>�4�؎qS$�=H֌&��oV�Ȓ�Q���=�u/��0z�+#ο���d�Ϛ�B��e{�EM���"v�H犙��sy[L�vws;Tp����9�Xw\�3{P����D ��H(1Wj���%���ͽ�ų��\$���y^!��7���!�&z���|@wy�-Vj��Gg��ȕ۝C������N�٢�"��-���s�fWG�d��oz�*�=�v��V��b8.��Dn�]㶹���I.�z�T��M�Sj�7XX՜AWWRV+��JC����Ǉ�1W$oD=����֢�j���3c�`�{��v�q��G���B������=�1�^oL�w�v�$Q��*S!��#rʝ0g>�rP̝��tD[;������Iv7�{v����O�`�9���=2R�}f�?u�3��X!�:<�vz��1df�5�e�p�Ms�;TG~5��^���o���/�E�A���{;�,BG���۪@���M��VU����#��H�L�W;QC��~P�KG2��Q=�m��?c��j)�<��O&���U'e�W5/�����Ts�����8�a�=�r��s�O/'_��=�HW�R%7_�A׹QL��$�'�A�֓Vw��{^p�_m��p��i���[aJYur��u��G��4Y�<U�]5���?O�!,�yJ{]���5�,(� 1ڵ���|.�p�#Q=��*���D�`���0PH�T�1b�7�w5둜�ˆ����;�e�)��_��ܚF@�A�Se��F!Թ1�-H���%`ض��m0��H�ݬ���`q�0ن1'HoD:�nc�˘�������i��&��;�-�P�ݦHAx�_��B��\*�����_j(������]<�՗4���o�gK=qKk��� ]ރv�h�AV�<R�߭v�Ehsk���fnpw�`���t>�7���3�[V\�rLu��"�J��R�nk���d�D���0���2��6���Q���;]	ٸ�s�ď��)��R�ĽZ�V#���,��,tQ�l��~s�"��'�l��>ށ�J�dB��Te�<NJ�N�F�l��y��x��^��J�B���?78�{
�6��4AܘL�wLM>Im�(B��uJ��{�Y�c�b8\7�qV�����ԫ�Ŀ���(<�+x��x~Ԙ���}��/f��N[=d*�L}!cSZ�'S�����w3g��&0C/')�";��:�-3x�vC�Nw__JRFiq�F���:�����s|P8�o��"p�;�-7D�#�x�ݳ	�JI5uKh�2���L��V��m�R���:)N���vs�aeuȤ��������Β��t5�%��d���"3Q�o��0�\S�hx���H���#������/�:�Q�5�&�\ץx	�A׉�eд��:������-@ܶiv��P�	*�Sʴ�8�Lp*��&Db�N��pg��
"\������zyWi'[�nj[< {]���4�K	�5LV���V�n5ٶW.�kb1Ϸ1�Rs˹k=�s�s$asW%x���	�I�v+��-�����i%1ʸ��Ȕ��s�T�=���[{TZ,�m3���9�}��Sx���4;콹��T��E�)H�G�0��B8�팃�K�` W:�ۍ��:�P��������,s'����	�'Rv��h*L��%ܡ
�)�C>0R4`��nV���S�hMRģ��;OYc�8�c�u�4P�x'��Lc jqw��1�����^ˊ��h��h���sN�bb����\c/�i�T�	�ЊF���Q# n��tkK��Ā�=��P�.����
��x�
��.�UG&+E��U��s;��pAg�M^){���A �9!C�k�-�_p���GT[��ZV�F�)��^�ːZ��w��*��;U͖���p�I�;������
:5z�y�S|fn�u0�f�֕Vl�3vts�o3>��B�a/�!��8��{O�6���Js�;˱�2	]uV�����@�tH�����޷��+���ܞ5
f�5�3�T�X�u�Uo���o=S:f��bz��pp�`�8�^ژ�t> :��v2gd���
dn]�,Gm(OyV'H;�v��O�v�'%�K�幥����8��\�+Hsض��G���t�B��3k�����v$� �s��e7*9'w�dV,��.�es�ݝ/#��3���v�̫O�ܕ�i�^�U���<}���t�8�=<m����Rԣ�1����z�r_0��<�3��Z7ɓ�q�{��
zf���=g�����W�[��y�|���/�Y���W�����p9�����n�Ş���ʎ֮9��r�f��1�Ν�Q2X�r|� ���]*��^�;~�G�9\1^궝��%j��^�e2��[��#/��/#d	F�z@���-�l���͗�
;{u��!��B*�Xw	�����d#�S/OJ�X�0�i�uo3�{*ݲ�w�E�ycz�vc��U#�f8"j�"�6��V�Ei����$W��ϸ�yW���P���cm���9U�ᒽ�G����青,���#c���;��0��_d�0�X��V*��"�j�3�`VG
���JnA�#�#�eB��6Kg2���j+`##=z�T�,[ϖ�^���/b� CD�RGGJ@��Ϗ��j�x67����L.O=��L��z�ץΡ�,����+�}P�&�rzV�w� ���_�Wi��O<�&����1Qgp���o{���C;JS*�F�+�p p�S&D9�� �K�ۿ�m�{����)�v`����ӹIj�Q�H�#��'on���ȔԬ���������L������9Cnq)km9,��Yz�֙����$���<QN�{���ʊZ�|����s+v�hY�l���Gr�CT��ȎT��-9��]l��V�h�V�:)M�CLu3��N��Ҽ�й��W(l�`"c�P|��c���+��b��|�h����4�Mҷݴ��oNE�ܪn�t.Ga^Μ�*�q#kWGE�t�DQ`P��j�	�έ�<�y�Q��ϽҰ0Ng�g� izo�VR�C��]����Iܽ��-�~��2S�}��i��u]�E�����R��eR���}o%l�׺)���<_���3	�>80���~>AG�s�o��=�)C�5��[C0�+Vh���'g��[~:�l\����H��NW�L�
��}����&W����\kڞ7�C$o鹰u�s�C������ת&@qj�Xq+�*��Җ:c`��?J�s�Ϻ�&��]���*8�yL��#̗���| uc�)�ė� 9ʸv�t�F�����0=��p�Ξ�;�+])�%N}d�)0v��S>�����֓q�]�1{b|벇�#w�gn�D�6*����rwsF����S]��%F�7|��yk���益-"�3�l�m�)Z77�������"���P]�3-`SE��3�w�4�TX���]�Y�%�S�9
����7:M�3�D
�P��uc]k�WR�}�Sr�<����Z��Ug�s�1[r�v �r�;�^��L6v
:4���`�� ڧZ�+��NR�r�rn�y*�,�<��e��ndL=b+����LH.{H��b`�'O6���-\`�6�y��Ws:,��99:U�ˑP��Q��YS�O���y�)�Ζ�|�Ԁ����Q�vExi�>�����Et��3@xUL�Y��}��9���饾�^�N1�o���@T�"S�&�������(B�`��:�YRʓ�{R�%��g��S��D1X�g@�V����>u<�Y��yO��X{�?	_i�k��
����+J�ڌ}ŮƠ����٪+� ?7t�6����d�_Fm>7�4QT��x��9��롩*�t�+"v���W�:d��!*˸y�N�z2����u��g�����2�jcW)2�����,��\umDV*w�h�W9�ƾ}�[y[�&,hc�TNR��X���x��?i�;x�� H�w<+21OFt�:�\1���t�4�=W���9�ؗ 5�x�&�^���֌S�S*�X�¢�9ܦk�s3�����Ŗ��=J�x�v�ǁ��	{�r��i�:^mb�v��%\7חRd��@l�l�̥+ �܊�5����Sͷ���JZf�wmrN?�	��7�����\���W[=����5	f�eK�[��tҌ��Do�jzE�no��K::���)L�5�&��k�q��p=�*��+U�.����J�ʴ�)\
�m�v��s1Ԝ��}w\��VZk�d��%e���Mp��P�F��NhJ�"s�t	�eд��:�{w�0�q�;uò{-sk���9Qf;SZ�|!�db���\��3R�u�N��S̎��h���r���y:�]H�KZ���r�cD1�m�]�b�'���L� u�T�߹k�d��Z�en��]x��lo�(s<4jN�0���3���P�X�c��B��q��Oa���:�~1J~S�Vn�����W��=��kҋ��^}�K�:cOP7Dk4<Չ��y��pQ��A@�
�qt���:%q��2����X؉SB���K]�@����+ڜ���Ɛ��]��h��}�"@v��T�V3b���0�/�1Z"�r�9� ��N��=������@F�Ac I�KH�Pk�-��r��y�/�=���/d/��)�M�����O,�۠��Ƚ��0��Eu5]�^�J/9���/+mj<'P�߮���7`M�/��0�w����Q�+r�ni������; ;
V��o0q;X�`�zQ�B��m����NYc:�Sm_�͡�P�԰���ѵ�^Sh;=�|��n��;���]wa�M�.��(�[�gF��t�Z��ah����U1��b@ޞ���g�d/B��UkϱE�U��5��FY+چ���pfo�3�ƻ����,����}i�q�6hi�F�RW0U��Q��G��-�׼�\жcl�M��.�&��O�k�t_��Tp��y���Ȝ���L+͉%i��&���WC&*�1U�2ΏU
Ⱦ@C%vR5M��Sf���uy̶�ۑ9�q�_���5\�db`�*o�Cb��O<� _:�xT���7X:�lÊ�]<�N��xn��r�Pye�v������������q?���U����Lx������8P��Nv����!ih��c^��ڤ�MfP��EY��l��k{)c��wF�hxa3Q��>�2��*ڭ�t�W;];*�̇����7:�e�����J(��oH���'�ߓǟ<F[83�u����R���7p�[OPP.�_f��;��Z�L���1"}3q5g�[�HD·Z(4�|�	�5U쫵}_)�y�x��O��c�*̣����J�3��M�(VRg��p���V�s�^��*��ǔ4�v'`j�w��GSU���6�,_\���w4VK̸�uu�5���U���B��ԭǛ;�n��	Ʉ����$����YBjp�o42cŷ xuh}�ܛ#-�;.uE΋Q��v�Ǻ?�i��#�����u�X��G�mc,�X�-k���� �hV=��np]�^Y�E�".��M�(+@U�p��_XC!t��hT����+hIL�]���[s:]��I�F7�46s�SrbJ�ej����+�K܁J��n=�I��|��Q�V.`��9�RN؆Эy��3'v�ݲj���Vɏ�E��g���tw��h��]cHj�Ec.��%Wn�55W �}\Ќ�[
�uM7u�F� �ܠz �s��kI_m�/f�lPT�ˢ�۹6��*Ķx���-PǔUj�ID���Jqt����AT�;�����k���7�1C�6���X-Vt���Oz��Ʈ��M�9�u%�=*qx.������)e`9V�������uq�d�"��ˆ���J����Dn7��S0E+h�d�����G���Jݍv��:Ʒ��+Z �NNx�z�Q����*�hxmn�����r+�X��f<�56��Ɣ��Kh�Pin�� �p�}������K�����u\�7�\P]��͙�u(�v��ˤ*J3uLy%vF/~��jM���~��ԓ�㢪ᒅvT.Q�A^C՚��Å�n�_���	��Fi��B�
�"4����U{��R����98ت�,�JGE$:þ�{U��[��9�V.���Jy�S�UiY�J���:}��vC�
�n@�94`������T��E����d,�n�յ���wf�0�J�ۉ"ٽ�,�4�����X�,��lg
�b�jx�۸����&���vU������]���ۥkg�y�<�C��E,�uR6mOVހ$��v&,�
]�w��ه��[���O���x��W������siK�<`���5'9�;� ���ʕ��;]<X��k����:ׂ�=��K6������Ŷv`���ӝ�� a�v��/\���D������w�k[�tf��U�������`u��K*R�;--����u�E1��SH����[�XY�m"{�������z�"NUC���Sw�������<�U7�uT�h+/9+;ײ�!v�A�K��Ku�2py�.9 ����ȱN��ڋ.�*�)�G0�ަW�}�/6���孡��NAP��P���%+���=�5`�QaOq9z��Sn=`\8��M5uY��3Po=��z�I!>�L�v��ܞ���y8��3�������]�!k硒��u8D�])B����i��)FvN�E��D&wV.�ž[V�:��7c�X\���#� �һ��<��I��^�u�_=�߮�[h�(�(�����j��U�2����,UKj�Z�
�1EAD�,F1-��Q�ZF�T��ň5�Բ�UD�ZX�X�1���J�Qf%F1R��J*�Yb�m��ETƆ5[lQQb2��j"օ�`��WN`UD�*�[%VZՠ���Um�*[(�(�kZ�"(���T
ؕK�c1X���C-��FŲ,PDkEQ��mmlR���Q������We�
��m��A#KQ�Ҡ��,`� ��X�ckm*�j��a�Q�U#�QPD�E�EV%��m�kPP��m(�R��UKZU�TjUXƴQYe�(��Xc��U����)Qb�T*PF+Z�i(�c��
2,6��QEګ"l�,-�EQ�&X���12�Q�UQT-�""�Ѩ(�-j$LK����Դ� �ګbEDR,��UEY6ʌX"�0TTA_��5�}��ø��lĈz-�0Vt��(ju��B��]}O�;�(n�h8F�Dc;~ш�hV�e>[���Ƴw`���N=�'qk�ѭ~����ǅ���j�� �,����*��8�O��������)�:���=C�e&*0��7����!�=ͫ>IP4�<9���M�N2b����d��wb{{�kyI�!B#DD��}��dRm
�Y/��_0<f�+<;�5�v�Y���bT:�T����'���P������L:ͦ$�2�3�q�����Kt�U'Y[��+���S�?�jg�OuI̩��*�W�A�f���q�&2l�i�O�T�䞜�m'�VVJ�����M!Xxs5�W��1
�>�HJ��Q�,�'���)�
���C_�������;�7Q�w�+�O��CF	��Ǘ2g�=q��g-$aӴ��I�+�k���SӦ��OɦJ��<�މ�J�d���VbK�Leq �O̙�?j��%E�����ieW����XڏDc�|D|�����>qX��q>��'�fI�8�����V��Y�Ϲ���Ӷi ��u�����sVLv������i�&0<�w4γHbq�b}�;n���b$��R�l�����������i��4�_�;�+=IP?'���ĕ��d�P�R\�~���N!^�n}�h����:��;�Oc�i��2M%C�1Rx}���6�>���+�7�"����5Ik����>����|�E
�a�=LCz��q������
��x�M����� ���������~B�:Cz�I�+
������
��T����g�J�|ܭR��F�gwr��
��'a��4,��/�oRc4���b�eRc��CHq��$��5�8���aߨx�U�C�ěB��{C0���Ho�ٴ%~����Y[A�{�Z ����%��4G�	P�vk�8ͫ:��I��w&���&x��L@�*s�֤�Y�%a���&2~qY<�bN�]�|��׹Hq%}M�a��m ��l���I�l��@"�ˡ�=����y�x��7�n��`"N;f=���4�j���:������g�����?Nw6�U�T����>Ci�3������xs=O�J�O̙��=Ir��J��+:�Bq��w~�M}�VQ[�N*9�i���uճ���yYj(D)��g/Sa����������}�i�4h�fG2wRĲ��5��;�q]�3v3�
�<%����k���4���;�.�v�{��,t:��t����c��R�BX�U��%G�� �� � �>��x�3���1 �ߧ>����� n{��!���O����@Y���ns��u�M��ɤ1>CK̯Tq�LFByqX���ff�٧:������8��|�q0�<�	��$������yw�̟$�}̇�q��z�r�q��O��?2M���xy����y��]��}���L��^��ISI8�C��/��&3��xY��Vjk'�䘒�S�݇Y�8���g��<H/��3�o�8�<K��c'Z�Y+<��'>q'�x��|�}�5�߼���<I�+������=�!P�%}���'����>���I��bJ�H"O�Ɋ�^ -Oڧ�xϘbb���:�r����g���/2c�#�E�� ��滀�����[�Ď�<a�Y���}�����J���s�x��z�����$�����0�!���1��:@�Y�%J�����֜N&0��q���i�����x}­��ձ�X��c��t�%}��Y�x�N����
~f��qd��1��Ag�g`1&Щ���6��+*o��x��Rq�+
�>�L@�W����>���f�����P�۹��FY�l�mRz���c���4��8���N'��!�����hc}�i�T�!S|��?&!�s���6�����Y4�>$ĕ�"ʇ���fbݟ`�Ōz��+u����"4�7a�1& k�a�Y8�z�]̰�O�=q�>̑I�+�9�:�x���'��3ǌ��4�_K�h�ɮRu�4�����:��ڛH.�5��\X�NAzM���
U��r�E��kLNꁌ�Ρ��6j���ݚ�&!�G��>a�I+<߹'�u%~O���I�*���`�HT�B�}�:���X�gu�I�+(Gۗ���#Ѿ�sIWo�z ���"��w��JLB����&�|¸�ڤ�C���I�C�oT=OPĂ���u�C�ia�
�Az�!�s�6�ԩ?!w>捵�Ğ}��r�hA,R��b���@�F`#K0q`�'fL jow���<������ќ�??/*4�6+���za�Ķi���1\�q��7z�.��Z�qk%�"yhtOHrID���!ƗϦ�d��1�ɝKq��x�h���O����{��_P*N��40�+��OMw���*R�3y&�ed�j~�
�'�b�����/�'��˧l
��:�n{C�~O8�{a��'~����Y���*LC���޾���w���>�;��r�3����} 1�h����ƏXm�Xu1��^$ĕ>�����Ug��w�	�6�^���چ'�z���v�b,�5�a橤�B�̞��Y��B�g������P�y�?~V�+�����_>����bG�[1C�G����:f�s߰+ѿ���6�^��i���8�3���wD4��!�����H*����P�4��bϻ���!���/��P�%}`ͣ�JϜ�y�ng�R���1!DG�3V��gwt�2_/�w=�5h��C~���8�R���sF�'P����I�u1�����4��8���w��� �H~?k�J�'�1 �w���nϖ�F�z��bf�o#��}#���Κ�gԕ��w��Rm5�i<}dĜB����i^�Vz�!�+
�����%@��߳ǌ�VJ�!�Y?3��&$���)]�Ǽ�Oql5n���u��lx*�w�>��i:��Sr����$�(c���iR~|��I��x��� q+<�4�L��La�n��'YU�Cs?ayI��_ۜ���{��}#�Di��[��}=������DX�Ì��;'��$�
�2l�����^�y&&��
����x�'���6j�f�/)8�6j��U������<H/�2�5��c8��SI��"&)R�n?zwِ墸�©�E��� �v_p�N!����c�a���p�x�Ԩ|�����'�8�C�9�A����s�����̺C䕕���I�(�2T��f����A Gҽڊη~�*�Z���I�m1��at��~C���9���6�Y����4��b}�'YP�=C;�!�0�,��|�hJ�������LI���Y*� W�'�b"��G�B���3�Q]E�O�|e^Oog��<��'�z����c���ʓ�ۤ�!ya����$���O�_�
���9�]��q1 ��jT�|I������
���a���� �d�{���@�_<~������������h�_-4�3^1i��)Q����s���e���ׄ�h��� ��⍲�-�Sʼ��<�B�(իʉi���Z�̎ۼWr�MƷ]gc(�/��������K��u6z��J�Kǘy+�.��o����X������q�n��ge�����|��1_!�B�m�Y�t�v��1�)����Rc�N&�d�Y�~�i'P��s�56�'��sX�2u1���N���&r�a����x�d��8�����jc������HYW��>���D���|�<H/�ܴ��q:�3�oV)��ϙ���<N!�bA|�?0��6�3ܲc�>a��Ss������sǉ�LI�+�|�Ğn� �0�V��z�o��,�=D�K�i;>��h~IYXq����4�S�w�Y�g̕P�XbN'Ɍ?&�Vi�
�����eM$h<�������1Ru���6}�x��A 4q��O��;[��^�G؁�+;�}��6��dğ�wA�+
���q'�P+�㗾�hT��SN2TYP�Ru��{�J�Rq��n���)
�φ�u�'�Љ}���
Y.�r}� �C������>@��I��3�ϴCJ��+<;܊H/�<9�M�I�͜�4���fm=��i���J����$1ݑ��,�u��w>�.n���7���S�<8�����Ԟf}k���<�uC���%9�fΏ��EF���m�^��+����5$5�>Z:�<�+"��N}�o!�s�#YTcʱ;Ff�
yŷ�y��,KrtŨ���0��8`�5�)D\�@q�j��˫�8�j�g���\��n�y����&]��y?V!ܾ�ߍ�!S��i.�E\n�z&s�����Gjx�E���h�w:0(�|k�YR�_�n,��;���T�{n��\��{������2��َV��a�~��6G�2�㉼����[N �n�F��s����n�寖ES�R����՗^����B���͗��D<�W��XzAo����	Jj��Ρ��݂������/�������\;2K=D���k���}ӢF���4R5~�@�f�b1��6#^���RD�&����k�M����j�X�'Z��f1^���Ӫ�(;<��R;�8W�_Le��!�{E�y�1�]�qb>~S�;��K@U�^�X4S�h��z}�CW�ؿ��Eq�^��I��$8b��sW9ٜљ�N��n��J� �&]�wr�
�+<�܍�"a[�.j�|iɒ��xԗԮ,� s�o#F�7���2Nn����N�@�徴�Cb`ዩ���/u,�!ZKp��CO��Q�O�M~�F @l�[*/Y��nxu׵�C���~n��|o�xme���tҸ;a�lD]��@9�҇Ϡ�A��x}�v ꃣo-|��ݼ�Ug-�Ӏ���b�O��Mqr}��`oz0="���ԕv��8j?=���v�9�M(U�)#��a�qe1�eFP:�$e�MH�q�qMM�mI"�-ۘ���͕W�F��h�0���C��*0;,l�`"b;e|��b�*a5�g�z�6��ru��ȯ.���S\�}C��W^�y|W!��U�7R�S/J�5�Df��;��6'A��kw[�j�v�ǵ�e]0���R�(�DF�an��J��
�cu$�woH�õ���3)ds5�� A#��\��wBd�&
hr%�v��W:��YJvqi^.��[��y��b��*� k@�=��9���N�����P��,1ciUK��:j��Y��~�=�~/l���_V	��y\C�zo�Eb�}��;��x�ɴ���wo��g.@"�0��uJ�;ّQ	�+�T鋂X������_q����>���Ƀ���F�q��ʌ�l��(c=���	�Uc�߻�V�b�y��J<�ؔ:�i�o�gn2g\�Ʃ�u�Z�l��|^���[�g\Η9�
�/�#�w�<���T�<>Q@})� ���㱓::����c����R�̷P��\�2}\k�l��M<xa�2��kY�`.'�/�M�	����\:U�[�q��u1��kY��훸}���ݼs�yq�z2���� �9A�=S@�� �U��a�V��_p�4K�LK�4�f�s\��-�q�p�}���k�,r��d����a�\C!zz}>���Nf����Ƨ���wk��8U	��?"��rDr7D�yJ�'39F��AN�)j�yG0U�%f�7P,^)t\==�xxm�X ��yZ�W)�C֨�,��r�m��)!��@�g$�d�dY��bz���P�Uee-:w"gee9�����\����]��f����#��5�\>��m_6;�`5��1)����Rʹru�a<���o¥�(f�縠�A��tsHl1�e��FB��2T�^�>͚�&y2Q��)�ZJd8����(!�_$��T��d�9��1�=��8����W*�m���Ď�l�&����M/b<H��	�g��lӍ�`(�Ҹ���Jj����[��{��Z�X�]\y>��(	�õ�լ��t�,�j!u�������b�K��	FH��4��
j� ـ&5ĝ1PO˃69��څy����h��iE�jk7bAyu��{�ƹ�Ȭ�B��˸x��ḇ8Y,u��^�d?�2rƪm��3����UZn#J�n3�"�]C��N�r��z~���9ҾUq�]sB��z���.�I�ٳ���+!С��3����Ҽ)��;G�؇9�ZUZ�5}�٫U{KR�@ٯ_";G�^�\$*��J���Uv�2U��@9��M)[���y�8eHH^s|��	�c�C��\�0��_�Wx���J��KºQ���y=�y��F�X0u1�ǳq� 4Wmr�T��&��S���2���:�4�mge�j�MA��m�G[-Vi�)u���^:�V9ؒ����O��´^�D��g�L��^�}��jS/�Yݚi�0�}��k�����l�ͯ��_�1G�����Rg�+�ґ�[�-)��5#�ˋ�S�Cr�������V�߱���P��9�:Ʋ�E�M�;�+��\r��E�U��;���c��:"Vu�y���N��pg@��Z:�O<h�~잩RF�����b|u'� 'M��n������O�_��֩��Գ��������v�r��u̐ʞ*�ы�(u%Hp�T�#:[60F	w���1*���J�ܨ���^�n;��`r�
��g���L1w�K����(k<-=�.w�I���k^��n���1�K��r`�~�*y��+4;����%p�ڒ�t��b�7
�Yu�%�n�<��M؇���S�ȑB��1 .9��g��ڭ��^��͢_\���[�SzQ��!�k���[,�0!`P�XȀ!���?!����n��)oV�d�'X����#fKY-E���&.O+>Tg$���l�g�n\�ܙb4K���{�L��]�w���([�_m�fl�&N�A��3놦
1Q�E2��%{�҆:^au��^CC���s�)��^��[��ozH�Es[�Y�{[ַ,�L���rwr�tʺ#��e�ł�g�*|���w\[�f��;��JP�n;r�!R�V�6�t�����yeoۃ�Q2�\:9�N-3
��T6dL���iK���0=����)U��>�"�Ǡ��wg�ȌR����
��yg�r������m3�ݪ?m�u�m�� RПϺ��ꃶtI��p���\�F�-�@����3������M�nW��]�6^H����r����m�����xk��]�"Kë*��xaS���*#e`�	�}��5h�o9d���{���\��:6��SjY�j(����-�yU��E8�{ݸ�QC�U��."��l�D�F2�;|s\�rX��MJ/^����*�.Xp]�S_�=�ޞq�����Y�۸댙f���3S��(;<��e"юwʅ��Ya/D�X��s�װv�́�+@V��_5�D84V\�&��p:Z81��i����e�ȰBM\=���۪���q�J͝�;fHy3q69���hE[�.j������n�P��Z������W�:#x����b����N�@�嶇L����&9��&�=Y+ӘB���Ҥ�|�R\=�4W��2*�7>21x�ِʄx�Α̪��Y�˜�2��M{k�.��z9fS�0%��.fmNц���a74�9u��i��U�j��`-����
!9�.b~������h��w��ns�{�  �O�f��'+��u� x�,��JL
߂��(����&-y����\ֺ׹����<���QSΪ��폾���Q!��Uh=�� "��T��FB�8����Ef�팚���I�6��wL ��LWԟS�E�+$_'���˂�O7��vX��g?rR<MޚW����g����i���5Z����^z���%�(y��`9׹;�XǒJӲr�I� ��h\5ꞌ�`#";e|��a�T����7�-­��C����Ev�a�Z��P��F�!�{NO�?��+�]*�{���S����;���m�s��uQd\À��ee���7���y���ǵ�^���V+I�z�W���Ӹ/{��i-"T��@	�4�w:�8�s�j���,ک�����س�R`䜄�(���S���*voLF3P�\��vɸ	����i��C���S�`S��v֍�U�9�������������ꐌ�_f�;`��<�Ӗai����(�h��B�+QՄ5;�q�%��}J(Jo���8_�+�-/i��k�
��g�mSGTDP�v-�g@�јn$Epa��N�	�T�Kw���IR���l�q����R�T��tX��#4��NX��{K�� P����zBE�y���Bi�c���{2���������]�J�s�̭�#���If��}�ݲ
��	/f�g�e��Y��8zۺ�ݡm[�)���&�����`�[�H�*�[]����H��^<�f�\;z�o��ש���8h�&:j��W'P�}lۮ��2�R�OD��ͼ�[7��6���R��:&^݌O,a��=*H�a��p�է�ƷV�T��Y͜����u)�h^�.n��
Ȼf)�듶�f����}���sw�_IhJ��޵�٩���1���i�����j��;��#y��ؖ*�,A�����I�uۛ���3KP����r�Fwc��g�]e�.������3J�JmA7t�*S�)ދ(l�=��r�J�XLZ��G-�N�CJ�e^KB!��p�h�c�1HM�x[Z)�|1o]fE�Q��k�'�V� [[E���pr��`�{�(���MU������څ�c�iv���Ԛ��K���
gn�O+;�E�{�4����kMJ��e����;��]Y�e�r�B��a#�C�rnP��D4�sv`�RY�v�1�^���F�껭ގ�]}�|-�n]��χu�%�򭀢�a�F�3V�U�
Ì�"��+J
��n�p�N��n�Lb��0$�j����ut5���e��{��ك
�X����oWd�E⌤�T��Y��E�`��rj�]-gR���j���e�*���Ѓ�m3j��r�7\v�`�5�̍���<�/*����T��i�AK�o�m���w��6;z-|�(��	{S��pz��qJ�$_f+u�B�*�ch���E�OB�ٺ��f�E��������֓|i��*�	p��<x����̰y���x��S"���E0�J��M�.�ꧻ Ϳ�I��[���2dJ��ͺ�-x!�۫���r��R��	M�޳Δ�UVoCF�ͧ��ZK���s�sVݜx+s�wܬ��%o���zA��xz���ӄ��,�8�$�P$f�E�B�M%Һb��WZ{��K*������ �;٣v s(<��j��f�A��-Թ١!��N�\$�~�_mn;ˮ�5o�8�>B��Î���>O�U�6H$1C��� �� <1ٚ��;:�������� �t�B��a�7hc�����-�:��8�\�2��Z�E��]�;���K*�ù��J��f����$�s�ëe�|��#U�ۼޥ��nRHb��箠��:��[o��v�+��1QCI�vyv��q���)�z���Y�� �tб�V����zq���:�TuC�E�-���d��%M�-Nn�������ۼ�ֶ�N陧w���D�L�6�<��m���68�C���o�L��M�5�~��x�J�eU��F �[H��mU�3(([GİA���1H��E�"2ڱ��UF�cDUb�T���ł��m�%aEU�Hѱ��*QDF�bDm���Z�X��eJ�U��G����TX��b�ъ1ƣAAV��ʬV+Qc�U��m(�YUUX ��(�KU%e��ch�EJ�UA�*��Pe�`Qb�-c�s�PUke���*�U
���QX�(�R�"*(��**AG-A��[X�,���[
-�٤�P����(�
֤V�d��Em(�(�Ŕj"��X�Ym��q
�V"��[,b"*�AI����YYP���Qr������ej.��T��ł�ő��*�1�TUV�B�R�QH�*�#�`�F(��-��AE�0m��Ԭ�l�Ũ-��m�%�U��+1����LJ��PEecJ,�AdF,�m��# �������EQ�(�e��R���Y�&U|�&�l��B�1��Zt�x3/v�����l��"Š0�ֹ=f]g`�ǶO8�2ds\D*��ʗ���vNi8"�~�{����v6��������5sw"��U_���=:�7�&�H��wV�o��i�����܎gu�j'�����SF2c*Uގ�8:FS�z��$�'�A�֓B��yX�;�Ɨ)��-�eZ���=mGP��W\<	� �7:!����N���z�*��	ȆB����ͩo���]ʉPz�4����ݟ//���}1񼜬zd739#�ƪ�Ĵ gJ����O]�pP����\@��w�D,J�gCf��h���*�{�"&X�x��z[j�l�Y��Vr���\1�U���|k���jV�3��^Z��UV���ž�^15Y�Y�X��Y,	2z̹<MI�.����-=Bb��7��.2���\a�Lv��W*{��ڥ�\l��#�1�:f����/A����v�y�����]��q�c��m;V�s�lC&|@i�nA����4��Pw���1�^h!=�Vĉ��J�U��*\\i��d+Cx׼��tX|��
���u�;S����a'�Y�Q��v���>�q�	ٵ�%�]��|�>/ι��P��CN\����������CEZ�{�}Cz�z܂�\ʋc �]y;6޶O5oY!"�%��>�2��9e��S�Kw'S��Ō ��Qvr��fn*{�*n�j9#률Z��fN�9o�,W��v�!	؃��������-�_�����6R���=x���UeQ��t�J�t��F����>쥆B�f��]�C�M�u���|k��2�)�o�qpve_!�S�\��^��S��枡}*BҚ3v�k��J%�l�>4�Ȍ��ث�_D��x<�`jΩo� N�	�=��ɞ�Z���ԭ�ɵ��ݴ�o��d(��BH�Ү�g�&��|+�{b!�U��oN���8/,�KK���rƕu��	����C��?�g�v��&��������B�vu�T&H���}�^{<�vS�8X��{4#Q �3�oM��%�F�n�E��ԓ�L��q$}���W�e����$���r�p4C���:c`ǹùvD�p�yO��ފ=��u��9 f\UHU.��W(4c�)�W'm�p�Rg h�V%ņab��[�6���F�.�8�N� Al�@hL�(<"vW��뒹C�mvS�&��q�_�=v��3\�ww����5�"*��K�6����$o*L�!��D�"�i�>�T�1lF�C�fP�cBJ(6KɄj:�wH�,�~�D>�۞��^��^��q����r"��F���Mw�� �͜m
��Y�����k�S��ٝ[cOI\���T��;n��H\4:�/���.:.���k���ݑ���qUj�3 ��{���Y7SgG��Ub/�g��V:��p�U��EB{Na~��kCeҜ�dmX������.Ƽ4�[�Lp�i�b��YrgD0�� ��P��k�q��������G�괦�h":b�]��u��j����{���n�6n�����Opy1�����wx�*|��[�a�+-p���ǝ�}Ќg��N����N�HyY�WJW���l�茢�'t�����g�V�U|�
+�vz����%h���p[�=G{1�cEPE�ʱ=�S�2��+�֋j�p��xT�
���4V�F�k�D��л��P4e�j�p"���@_]x¾��;����'�㰗���+�ߏ��N
u*�ɚ���xnOt�;3v T���B19d�ų��h��[��������l���K�#n�T��;,R��裞�d6W����B�h����[ۅ��4Tcʝ=����N�3r��^��ך�P�y�Rm���Q�:0�3_N��� ����g�o���הCa��}@�M܋�e+�3P=8�5zp�+ݛ� |��h�C�cn�Cn�v�pcX��"��Q�U,q�t�-�4�ڬ܅b]��u��D�|wV(]s�	A	�2�!ҒWZ�����rb���r�R�����ҭ\����fs�|��Wՠ�̈́���{�
;Y�t�[�5��}х��~�p&*w���_#�e�������RY�:��]#P"����S�����k�`�o���y�>m:������}�0�~V��i+�SN�/��|��'���+�� ^�o!������$d���ݚ*糈R�g����|�`IG7��圮4PR���x���)WT�M�p��e��q��_^�0�j0:�cC����/�3�1�'�%.늸UPٿ��h=�'| �y�!��!PMc�rW��V����m(���^^�� �wN@!a�I�������fd�R �lV����i$V�в���1����h��v�g68���\�����c�b]�:��{��%�~�jI^ݞ��߄���JA�zиj��$��5&*4��M��������ږ��o9�&��uuD�=��:q��Ӊ
�T�����;Ή׶hģ��7֛�5x�E�^�[UED���
!�ey�$�=�*qf��y����X�OY�,�a�Xt�����C��W7����N���(��z*J���c��ŝT�u�:�d�G���k;�.�?C�Ӹ��V��e�W�V^9�~�{g���K*��B�c��)XI��M�$��oEΩ�dw��S�M�m�H�33�I���������m��z��1��Gf�9��Q'1���p8�w�#[�/�Y'LT��_1��Ӻ���R]��5(��2UB,�8��>��i� P����?K�3k��,�}�#�ZiM�~��S���v|�X!���V{>��ʳ��[��?�|;`��S=��Z3w=L)=���ƐF{�Y�W��O���(�9i8��L�4.g���AC{���hH��MR�{�h���:����f�&�����x�/�W)����Y�	�\;j����Rۚ8���ޥ����v)���qq^�Sd_����Ën���E	��k���q��r���:�L������q����<	�!qD�۟>�4W��C{*QXJh���8^���+��%&��O�T;��-e����>A�-�`>�Y}�7-v�=����F�V��*�\}�:�a���)v{H�6�Vb|hn2�_�Cf��`�	�ҫM�D�H�iN���o�9)ڧ$8^LLr��&��,as�b�!���9̪sML^F�������0��>k�	9�Å�8�g��X96�K1���:�����kݮ�O��镺hEͦR��փ��rwV��=܍�霃40�u��R��ss6�8�~Ns������8GR����QIoCs���'veR�r��Rcr�e?}��U}�x��ֵ֔)�>���P��M,�tx�����i{��D��L!nz3,)�v0�.�y��Qڻe��EA��7:jK����F�u�菕o�^�������Y��;$"�Z�ks)�׌�H���꽮ӗ\0.�(8FD!I��B����f�U��t���r���i���^�_*oT��S���!�4�׆���P���w؇3���0�h����p�T�?~��Z��g~{i�G_��u��@]p�E�`������ٛ�[.���N�!���HD�ܻ�o��ms|�VO_�&�1�E�o��LV�����_��PX���J��75۸]l�l���������
�����RF�>�>U�/�vxKJ�/���1�N�H��ٮ��:6�@/z�ϩNO+��>�F,f�"(F�L�f:J3��N'85�CxG8s�lGdw+|r5L1r��xm�d���z:�P\����?�U�������Nr�_;X�Zj1�3��id�������u���ˣ`���|9�]>��#�0�[�/��=>�Z��p3T���k?�{��n��l0z�{��(�ʴ�S3�GP��tZ�'������49�0yuEV�F4v��Q�v���n�Ap��kb��n��8��3Gs�լ��-�g�W�������Yұ�Y���*2�������+���]��\�"�b�BQg�W��|�뇟A)�g�1�q�"M;x�{Kx싗T���\潜+PTh��������9����.�R����c"Po��/���2�X�.d�r���ޮ�Ҕ#ne:(d)0xB��E�v�2:��j��,j��J2y_>���!Z�Ì��˝��h@-K�6����#y
L�(�u����]J�)4���NJ$����T��AʚŎSw�+��dHm��Oi��@v<z�l�̓�Lq7}�����t\i�7q��#���Oj�ϔ�6� +��d@�oF<�#v¦�M�{'-����kF5
ՒP��6�ƎD��s�����D\B9`tU����u'<�#�����XV.8B��B�y�T�^�q�e�q�:�����EsY$��J�T`]Qy�VOl�{�u�{S���@��p���V��~�VV�8(Eb��Nu;�3sa�yXj���g�)��!���	�Oma�����$V�t�����²��c�o��g�,���G�\��']è\��☍�	�G
@�ֲ�����"}k�q}c2}�8U������u/��:��uj�il<�偪[D��ou�q�
��WY�Vn̖.Aj��+ ܫ����#��٘:_WV_v��x�!/�2�3��LP[1wlN�� {Ձ[	's,<y�ﾪ���X�-�7���8)�*%��B���������5\��<���!]qy[o��A�^�%��`��˻Sk����S�:��ul����;J��L���x�!d�s7#w���̪�@�pQ��Ih�{˰��,5�Ní^��܂Vz��yc[��י���,2h`.�*���o�2�1q�0Y�SA\@(<7	�e#�nc�޸��H�V�;¶�N���޷%��[F'LD^L�&�x����B.2ep����KG ��B^jdD̛�;�yO+��r�ܞ�/��W���u���J�i.������Ot��\�J-��|-b7a�:��n��������{\���'(wJoY��]C��p�vDޠ�����4̷V*2�ƀt6&���)�B{$h�i	ӛ���cDBDlL�D���6xn9�ۀ���.	�wr����q���Pٸ����%��^������M�^���s�|�ᣍf��(|eN����r$�}��^���|����o�'���3���ŵ�� ��,�?
~V��௩��|4N�������Z��qX�ycC:v���%�P��EPv��}�z�]��t�L���9�8�sH�V���v��NJ�m����&W~�xzһ�3�����'��4aFGi�����1��}V�8���Z���&8�M��т�z�]�S=� �ץ�6���7^��=�ѭ�M�l�uc��1�j��e��#���[�U����#b̓���K�iH&7�W��f���5�~��HWY^a�{,j�����{˷dE�� ��a�M�4�zee�u^�g�	��<�#��#eݭ�U|�{n��n7>q}1���;7�hXi)'P���P8���̊NH�Q�<����$�X���c�;�2��eĹC.2�㰥S�"�P�\���N|�w\��Djy����ޛ�c���"Ë�R�f�p]sXV�cau�.t��<�i�@�fZi����]��%koާ��+��p��|��Ã��񖗴��Ht��kR=0�uܬ�5��h�}�Wp�'�b�[t��88�zj�5;�fXDT.�bl��O�f�����������W�卹Y|���'E�� m�>b�1Q���)%������T��eX����Oo^�b43o�I��}v�}y���EuZ~�s[�Tc�QV��R�����Tzf7�*q���[|���K������^Tm]�o��濈|�-y���Ǻt7ޙ�㦦m��7:뒙̊=�$��>X�U�W��{�u��q���΢~��{-�y®ڇ	�p�Z%��j�о�uY�(���5��͜צ&����:�.�W�eSg`�Oi챈6W��g�<�M��`k5������ۣ�or���w�6�=ҧLH�����]�Ā��!�w���ͷ!W�q�:dd�g*����I��s�[Jc��M��61zbc�]q3Ja����ʄ���֦.�g��9b)��^V��X\���q// 5�BW���t����צ���/�ꬽ�]���K7��w�j������ֳ���`����*C�"��>;,�=8v�,h}M�2,�-Nُ}�r��,B��ֆ��b�@�CST�M��l���#�����&�[�6�~�(��5w�󓺗^���jO}�����L�wL4�#�!����z�0Y����*,�|E��5�`Ň���������k(qp��]V�����^�+�RrZ�p������=zO<�cT?z�ڳ*�P&�:,��/��k��ٗ�g���p��U:�,�^]���i�6^y�˰F��o�Uke�Sl'w1-/�"﹕0���N��m�b�l�
�����f�٣ؠ�W���*-��ս�c��R�\���f�C��!@�(h�6��I���umus��nU��]�XNηl\}3G �}�,H���n��)d��j�l���`����2+�䬜���2|CpB�μ�Gt���̵�����J`���Z"�w���K�ݷ����jb��4�Ix�Z�:V*w0�T��wt+ �1�O m]	��?4�����F`�%B�l�MvL�z�:ݚ��AY[����d���d1Q�wU�b�\��}����]3�G�+�[!�0M�U�m
�w���[��u��imq�p��YS�դeH����1/����$c��s;�gwh��'����j�$��c��Q�ht���+)�(W��䢶��s��0�5⓮���O3k���<���J�N��2E4T����)�]�,�H嚜�as�w�r�G�����r^V�"�BsiglE�@���ȫ�!`M4���t�+�Yt*�ȡm��J]h+��ÊV������{5gkK��95<��s�á;0/n)x��H�o]9�7Z�6�@�f��p�bv��O��Þ�'[.Z��U�rx���*�-I|06�=�t·�8@2g!��A��ŴHChZj�gg������ sg�-+��p�Q��'>�M�l�餻�˺s��7+�7����M.�̍�5|�������K\(�/{�W*�Y���zPY��Y@���]s��D��51�ŀ��}j�t����*Q�,8>y�R,�Zρ�`R��q�8���
�KJId��a�t��R�E"�v.e���W��;N�3�"n��s[�cض��Ren�4
��e�8v��X��L�r��W|nShh.�,L��e'CF��׀T2����'3���ג�1A]�=4,�H�1���Õ�.ؙN��.}.L{��,t��X��,�2|�s��17ɽ��L�Jo.G�s�^�j���N����g<��]�4ۖ�[��Mov��fi�`4[��<]�����7�\��g2l�t�r�'ف�ҁ q�E_�]W�:w+����i�
`\�^��<E��a���b0TT�b9ŮT��uW���)V��^�ɮ���N�9a��W�X!ivss�7�-�e�9K5%�2 .��]��|D�K+�w���Lw[O�!%�ڵƶ��sE�iҥ�:�WYf]�*Ӯ9�ZÇݾ}w\�*K���TH<���CsTom�,�V�QZ\�e�4�d���WGh<j�K��%�4��wǗk��9d���]��_�\.rX��>��s�q{�Z�&FBSFk.�UՄ�z%�.��f��<*�xy�{�z+�QER�EYP�*
���0DPF-�"��Pb�"�*��5�R�-���YEP�(�VҊ���T��E[@m-J
EKJ�B�Tej�(�-,�اQ#��U�i[��lb��,���6���[U�5�,De�+VЩ�+�`��8֥��A
ʶ[DQ-Z�������`��m�#aib�e�V����m
�"2[EY�X
cFE#lZ�i[Uَ���b
	��[J����AT�GHV(��Z����*-�aD��b�eH��T�E1��QE�,PcX([H�`�Ջ6��eUV-����e�q��
-�`UEUR,�q*-K��*+D�ҡcR�V*Ŋ1m��U�8լ�lXpkX�-EA��b�Z�J��b�-Db�[DE����-��TEc�e��6ʑ�@R��1(���ERl
�-Kj�88�X���R�Em*��T��������
�1���Z��X�)��~�O��ۯ�^�"%�@ֺҝg\֐��g��Em"+���f����6������4@�1�
���"���_}U��O��<#�dr������|�6���|��$xT�U�*���*ү|����d��n�uF=Ē�3|��щ�+b ����\S�6�Oo�g>�F.`)�1cJ���5��m�U��˰z�.zf��+
���&xC��э�����ܦ�6R�X�]�/F�po��`�]0��J��׬��������e�Hl��*����Ơ�<¯L�
�:�s8�-|#ܺv{/�q�|�ܼ�yδ���wq�Ҁ���19�$.)>�k��6ph�;M��"��qڦہ�B�r�tr��o��x��b"�:8�ۍ�������Մ;���4��H�&hiw輍����]��{&E�Ӱ9�\��flBș�4O3�p��.�%�[�N���t�Qv��..a"����K�t��!Թ#h@/NW�H�^����.`���ws��1�\�\�<C�	N
ϓ��˸��b6 ��w�WXU��x��	1�+5��=�C����q���0�o&+B}4�r��(`�!<�+���B9l۔dՙ�=�v͖�0ﶮu �VU'W4���t���˥{nJ����r��!�$�,\���N��y�s[�l�$s+T����[!�Y�Rn��ݡ)' �^:�@�oQR�&�����b�K�юw���T��:F�#���`��{����ಖdEuuu��	�����l�Nx���>fWr��#m'sf�j@l�C���-<��6�v�r�)J���X�(!�y_*����:��uRg_�ğ�~ǁ��s��P1�̚��q	]��t��J5vy�a�_/���os�]ضrr�̓җ�ݒT;�׊j4���
�*.�v��-�N�$lZ����X��E)�{��ܴ�6R}�f�e㲐P�@���3�h�y_�c�X'��/t��o���B�^�a񿼧�ov%S��"�_R�p5�5�uHb*��&�!og]���{Hh��]3�2�"B[xH��r%�ģ>}�oD�hw�T�O��q؋."B����9�[�,Fi�ip���_�^8��K�����Qm�(�Wi�(��ER~�w	Fm��W�u�²㬠K��ǀ��IS��.�|�c�����nG*�ei ��-@V�K�T�i�/i�S�K����O����i�۽ڞ�s��ѱ��L�T�g��^��X��8!�����;fE�
�m��h�)�/u���H;�8�v�xq>�]�4v�qwJ4���Әs�׷�Λc�k]��w�lV���������J��$�ԗ�>'8�y�hΫ��<F�]��[� ksa���c�ݣ
DM��[bU�Ꚇ�s�&v�!)�`��Ӄeo����j��!�ϪH�Ν=�y�v�q���)��vO3?p�"@Jg���x2��B�<U��/Ȭ�G�
��ezJ�jD�r�6jd��qL� �t�w_X�
gG��
\J��e�=uV�Ͱ�z��KGw��]���7V��p&!ک�,�˧Q���S��B��H,����p�;��vPo�y>�:+�3L����v�`���;���'�y�\<y`TveD�7c��4�+��"6Ϧ���4ˌ�Z�I��n��!Ww��%y�s�qez�ϷL�G�=uB+%��y�t�h�I��Q�Ycd�C2�s��[ �\���Nj�UY,\}1\�b�9�|���=Am�H���K�Evk�y��)G�{�^��/n_AKO��p)�G�Pc���;P�E*#�����0Mfz��m�:�����ia�l��m�Gl� $�ң�1u�#�0M�T��̐��pf�������%��Z�qY�p�K�zg���� i
<U]���UA����<���C�n*tmbv�wМ�VrҸVA����0��Ns��gJ�7fqN�0�)*�$�%�u:���[���9��y.AW�~��������mvG�.�9O�d�G��7��Ee�y5�n�� ���]�Sy�u�	���׃�u�3�Vh����ig�g�9��B�x���W8����ٜ�f���.m�!}jp�d\�55(S|���%|e��<Ĩ���k�j�[�-��H�m�h�źhܛ��mx��ે�N����� �����l@�9�(�/(��ݡ�9�pL�Vj<�(�;���ڠ��9יo�*�iގ�F)i�ز�S��������Sͯ�L+{p�'P���,v�>�4RwP��Ec��Ig=�mi���;^R��' F*%�Cg����Ɏ�,J�L�X(����{�c]�!�:�X�����F����y{MA\6̖���bWq3���؉G��*�)~{��%;�~��1�^��w�]���R�ҥ[�Ǥ�ʼ,J>[f�i���r��E{�˄�冊��6h;S亙�d�3�AS3�b/K*}��$HOP��E��������5!��1N�����(F
����r�>���f����<�L�;M�.��KS��"�Y�YPb�g�.�Q����o�����kЗ�)c�d�����!d:�W3�Ә\L�j�Sc��y�`�כҗS������E� �K̢���ʈ�����׵��S�7�X�C����{C-Ү\ڻ��ps�v������v��}g�jJ�	�`�_W�W�sލ��8��(��J�_n��㩌�K�D1i��5Ch���I��I��\�I<&ޯ78&��Rz���v2a2��1���"�a�_Byw*A�[m?�V�����5���O�BE~�P{�k)U���JU[�T�{kƽ��À�.3��+������ӱ��"�N3���+t�8L`��1�*'�8��*�R�����;V�
��{o��e���f���~Pj��_���p͵F���~r/��o/���4�N��z-6/���<U�yۯr�	\���q����z��ۇ8����笆�O��Um����ƚܦ�������؄�)B��ӛz���~��=��zv�D�BzTZ����.ֵ�܂��w��i)g{o����Ʋ����Fږ�Ѐ�n��uBO��i\=�Ɇ
��B��M!������	Wã��e.��*�W�7�W�N}������v��kFwL��PB#���>�k3-`��m�	���W*)�{zy�{;�ԙ�|�k�|��gz�Qr۱v�>�K����^����e��}xd��΋�׵�ʟZl��"�+����78dܩ�Tu��(-�3�Gu?���"6e,x�C�[~��������*�%��x�@����$��=X�>�-��3�3�����k��������Ǆۮ�hT��[���q�+�<��97qe�ոٖ�u������9���<�����]�e�D'@V
����������]��ѵ����;�����*�V���䤹:��=�[ܬz�v�U�]fm�Ju��Z{�'�v��o1N�y��u��f$�ӄLw2�>�4����Ex.V"�w�r^����z6�b0��r�ǹ(��q��m5.�7X�+���@��]�*���	δ']J8��n§&GV&�����Mvmb2׏E���~�F(�����R���lΣ��[�S{������@١�xwQ"�q.��4�8K~$�[^y�i�JR��g�=��>>m{�l��?1ygx��Ɓ۫��۲�Hd���r�m˽��_s��*�j�.���nm��cVH���9d��-�Ű���0#�z-���GL�T�R��
�3���jS��u",��s��������UܡtP��U�o_Qɂ��{���=�V�f��7�ܚ��5Pק���+�-�*=��#y�������J4��-�ښ٧�K5��j{�R��V�v���6S�؟��K<6S�s�{Ӕ͓�[�4q��tc������R����ށr�
!��aLgr��Tk�95M�ors]��
T�X��p���ʈ��
\ H':��D�7+4���ww��\�;{5�M+|;���;��	O�a"ָ��Yn��%��o]���t���iK����N�|�˕>���:&S<�)8Wg��ʮ�W5P��	�%�5�n�g4u���z�ZJWb�2��n�dr�D��Grةyw@'�qҶ�Ld�{M��!d�f�׋��)Ii9݇pD���oi�����"��ǷV.��/�A�޼��RE�cr��lv�sc�#7����+��.��a�aw�u�����%Z�b�V�JHإ��A�C�ĽqsI4 :��s�uʳ��s��奛��^@�ΥBd� x��s�����{4�ʙ��)���2�Ü��c'x�{����:�e���5@,�ݞ6�T���}��ӻ-O:���y_P^�d)MhoO/3F$�H�^7�ۙsP��[�Ӎ��J'������c���A���7����4���GGr����55�'[���:c��X�{�mՔu0�o��g�a�xUuQ�4搩�β�occ�����]Z�J��z�R�^���z��{GǛO6������\tb�/p�=_/�{9�m��qv���ꝡ�{~Q��]��ZW��P5#���O�+��v��D,����T\V�QgA{B�<X�[��C^�MM<R�kyp�kr)�
�������hN��5�_\X܇l.���?����x�d��t^ˇ�v�oj,Sqg>��3�E�V�n���>��*��܅_%������4�>�x3��2a\`��"�R���^k��8i��U���� �ݢ��yq��_t���!1܇u1N_��
��V��p	g?��Ա`���A}K]���2���~LN��X�^��~���	���h�r�M�� '��b��i#�ď�2��j��`Ԥ�.��H�z������[g,p|�v�-cr��pu:��{�'h��!��Z����>��>�y�m6�AJ�9�OxBS5#���.�15��j�9�w|�.F��S�Di���[���!�S��lZ��Wn3[�OA]�����H�3%5r{��C��V�_u��w�8��/#����WeA��ll铭X�dʇN�+�+��ϲrZ���+�T$������ؿ��¾/��5d���|E�I�k,�ڝw/w�i�3������S�:�!TBj\)�w�3*b�Ā:�ޕaM����P1h��2����{u]��~�lu��Dq��\���Е��ff\~��W�q�_���^�W�/���0pM����yN��ԧ�ō� ������~��S~>ū�x�f�U�X�%]�?>:0���Z~�������[�SGp:�*��-/Suϊ�Wegtwc�T�:�K��lT[O�)��j7�&�w��~Яԫ(#�/Y� ���L��y�EHt�*A]�&�jR��DJ�j��RbJ����F$���x0��fqf����]4cm�n�+lK��'ե���Ա�=[�
ܬ.�����r.�o0�X�=���S���ӄ��5 S2���8 Z��}�D��n건�׷k*�*��r���������ݔ�����٦j�9Vb��?xV?P������H��d��|��5<���dS}5NR�CE@x[����v� \n&�Z�����-�Y����j!�t5�m�9��ʆ0�V���Z����au����I��۽����X�`�ה��G&��^4��=0nWK�K"zg�Ϭ7sWng9�v7�e+��{ɬJ�����b�fʞ�vl�f� DĢ���7�eRƠw��Ve��Kz!�.�q�@w`}h���(�:ܢ���ħ�~Rp�n�c�g5����0r��N�5o (y_��OV�F�v�Cm�9�$1��OB��Wu�uӘ�6b�й���N1�3�{r)�ݍ���L�~������G�}6�]�W��aT}�=�p�f�e��m�w	B�n%�tH���zo,k��v������B�:1�:B��2�Қy{W����Z8��]K��`�v���c@p�7D�.uׅ124YeĦ}���0˹m�쒳i�F�<�ڑ�I3��q��:�ٛW�J7�O��a7t��u�ݪ}� �.�9�K*�GR �t\�SY��f�-7�,s��A��ZW'�ɢJDu�u<j5�������j�{����:q�sq��3ۻ���l���y���'96v�s���k{����=���ʗ��@�2 �/Oe��I�,�l���e�S�Nz�2cRP����{�1�s����կW�ί4l���	:���A}� b����h���B�_Ɇhz�e�ʗ,�$�i��{Z�+u({&>��EJ�}xj��4 n����⮉v���]��A�Xs1�egM,�GJ��FWA�L��Ow��۶L�x8�`�_^'���[׵�H��Y��z�u�`�Z��e��w�t���,������C������ÿ%��y��"��°3���TB<��ۛ�8�F;5Q��ـgZBu�S�m�)�cv�����Ҹ����Z�J�ں�˼v㰢�݄61]���4����LZ!D�?_shڂ��:�^��)�G��wIS�  BM�m\UއI%�x�f��ϐ�C2^�7��k�(�K�Ms���S̵�:l�v�Fwel�nlɅ��˵��Z���e�܎�վ��t����楚*�w���Aͻ�7x#�_Q��j����Ĥ��R˙]{�p s?h��HM��[I�w>_3��z:�.&CQB�;��Eɗ/pT��oP{I\�_n2�Z��I��Ghgt�$��V�u�%��M���sv��m�1QIڦ��/��V�]�Ɣ�����	�~a�l��܆�:��^g��������(�&��U�s�:�; �}0]�RI�%����ʇ���{�<��i�y�	�سV�B�tq.->ܭCXf���i�v)Gw(|��o�<I�mnd[lA{u�Yz�ھ�/ak2s�Ͷ��0����}E#�a��m�&�[)^]�����Ԙ\�C��C�u��"R6I���w2Uul��`�+-�0v�_Pԧ��^�;m�75�l�LhY�"�n����h�ήn���,U�2d��r�X����!%wQ}��+��?!u;u���h�
���PC�Xz\]Οjŉ�S�Kwm��b/�B�f�v�n��鞄\4��_N'��y��aΛg$�ɣ�t�M�x�0E���)������S͊.�(M���X3c#�m�b�,�<i�Ħ!-��!kh05��R��a3���&�.��u����p�In���&r��v�y��aR�>�و���	_	p����8���J���q=��pQW��r��4�o�govk�0�r�B�2��!4���"�S��d���"(�X5��BѶ[EDEQF�
0`�֬e�V�`����Ah�Q�m(�B֤UE��֠���E�PZ�,X#Ҩ�TVҊ�PX%[QEam��F��UR�Q��K(��+Q�h��KJ� ���TcYUD`���FX�D�G-�XŊ1m�*�R�(���Q-��R�ADb���YQHղ�2ؔ�D���UJ���UVڊ,��AAb++(�X�2�YZ#UTU5
,T`�V�QV(�
�A�*��jF�DkQV
����F�U	mA��PX���ؘذX�U2�F1�%A-E�V�
��ԢV�
����
���*,P��F1��Z*
��EDV��-��-B�Z�*����U�Ab-�QF%���V��Q�E��5�(+"�Kj�"*�0QV�R�QV��Z�@B�+�`�X�Q�A�@
�J�@��v,usk7�4���H@]2�֛�}�z���ޚ�A��y�	���"�����ci�Z�������Cw4;}F�Ͼy'���p���H���o���*��N'g�3Ni�C5��|�L�m�5����5N8�q��rÚ�m��o��Է������a�ﴩ�cu�z��+�f�ow�K_O9�P~P�9�ݒ����V�w+��m�Yu�'nb.sj�j�F*S��y��ˆ�Ts���{��I5��f��=Ը/>C��ok'MjhQ�@Wq�i�u�׷V��R��k��c�:�{����#���l��g��u�8��[~5G[ښ�6�q=py��׼���
�V�J�`���Ҡ��S�
l#��4R�*�/嫝��u�r�v"�P��x�-���k�G�����9��(Ϲ��C�Qs�^�J���X�.�y��� u�V#�sW��B�ʕ��-NZm�m��f`Ӊَ�Y��ү�Q}��p�l��=;��2����q��pĒ�M̳��P�e�J)+F�ډ<X ��A^�w0��O^J[N)���Y�۹���EP�ښ��c��Ʉ���Vⴶ+�V�9��B�����1��ݎຳ�u�ӹvp�w)��M����8~�������0��y�l�׾�G9�t�Z��.̽)�b�[�e�q��a�y�5�"z%���:ba����+.�;��e$��=S'5��٩r�a������;��]��pWh����D�����-����Nl��/z\��3��%co�L�5җ�+�l�_ǷOP����xl��o�k)<FJ˃�o:��A��II����6DぷG�*�GR��?�ϝ9�������W=���}X�c��<�(�cj���p��#���Ս<�;���I�_e|sn�_E��F'����ja��ō��aLp�j�ޘ�|r����>���qڣ�T[��Q���d�6:bn��&�v.wV�d~���l���ᴥ���4	�'��\⨳��G#g-��'"�1�k��ތ3�]�=��=:5��x�^A�J��$mD�5�4i�(�z��/���S��A����0	�`��s)�74�mZ �i�,\F+g(��s�V�L���N���w�rnr�/O5�1/�;Y��^q��m������B��6d�|��V���z��v7~�؀oEl7۪�}��d���Z�ᮌ�Dk�����g�W�7�ؚ�Y��s�����	˚�t���vPrѪ��,�j�6�#��Z�.�&��q�΢�Q��7}�y�Ì��k��KVv7˞)��. \fTJ��
���1t·��w��ߣ5�iy;u�^+&��w�J�%���a��$��B�����u]�����pe�䈯w��Rd���)>�NS��~o���j�{uV�Ì��2z/f��H�kf��6�\59�dC�T�ʲ�3�v����+^>���L��D�.�n��f{:�îZ|��Sb�<^GRvf˞v�Z9b�Cצ)y������w��{�9�Prߧm��ӸeC��[���΍v���<Y���0����m���1y{7�S���^f��;h9��\��)�U�N�L�z�(�D��V����^=�ՠ�EbiU=�r3J�ڭ�&��jgr�lFꀱ7���j�ެ����@F��F���"��u��ق ��(-;�IXG\�\)���v�S�����J�B�}B�Z6��N=Y5�<YW��Nr�G�V�ъ�J�O:-eU�}'�0��lS!\v�T�Z�B���۽�1��)I��覆�%K��{�;���\�ބ��>YG߭�ד�����Glҫ��{�kYS�2PU����N>k��� �궶��߂�SO��N�p��ȝ�� ��ꏩ�.�g���)qbR�� ١��V�b]-c/��hqg�c�U��{y�ظ���}Msߗ�{G�Z;�>���q.G��7C�꟭ӱ���3�.ookr)��=6�jpܬ>RgjG�ޝ�s����Q8�,�;����J1:��6�l����`FJr�vSi@	���F�쨆��1�X:7�y�
�hov�Ag"e�D�^v��U��[�	-����,	P��.~)p�}x�ˍ�`i��n���5b_�sSjZW5�;g*��Z#�bY��5J����=�]��/&��Z�Jbky�;���r����ò}�m}چ�W��o�4�ʾ˻��]%Y&<A&�z2�2-�����~�U����C�e�Yr�ZS�Zt��'uW	�a�$O6���7�{��H;�NfRYmU�u'�e��>�eb7avu8�TVݒ���]a�짊�3��菢"kr�j�[_W�j��>̾)��i|�C6¸n��܃���]}u��bݧm�g7��'K�V���LmB}N��*|�����R��KTo�~��=K�=)d�Z'�--�����ʼZ�9\򠜅�z�Nd�ݴ�[Tm��	az%p����5��]�[fc+����{q��j;�0ū�}�*t�[9oK!�[��z��u�Ni����f�ۨ��m����l�[����#u�ۛm�B��PKS/�d�=�t��=��ʌX��D��(I�ѯV;�P��F��.��.�o'<^��7>�=�iz/������N��j���Li�c��g��Ņ�XV����}r�(۵��M��[�f����)s����b�ʾn�P�ë��
���`�g4(�F����z�޻�Tqо�Y��������f*iT��N F.U�ts8�T��r��B��6���/Jˬu:�V���ck��s �����c_cd��M�c�yCz%���n�:��(j��b��h�F�l���r��@wK�A����<�����������o�˿K-�[{0{w/�zW^1*�v��BbX�ֻMk�s�޽����������V�P�����5o��I�+C<���MR���f~��y]2���4Ҹzo>�C��w�nY|�<�L�. dfԩ��"�;��J�8�/I������� ���d���;$���լ��"��L��Un�`ovP+[���Y���f��~��)K����Tz��u.B�#��������]���8��F�/w�y%pw�N��Uɞ��V��E�I�Q���.x�CBP�3.6��B뷭�YP��N�P���:��"c�=A�T[yأPbP�7����������O{��k�n7�sƍ���~T&��]-�^��"e�no�7O�I������|�j�}�=�Խ֝w���~�N�-8�l�X�Լ�S�r�Fs��d�큊+ۑ�����T��Md4���+k�Է\��V���褟xx�|���pN�R�? ��T-�{�B��~�ۤW�z���U�Ɇuc��6�Q�V :�WA��;}�wR��{@�uNj���x���������m'Ii�[��Evu�[Ssug�����}�O?u�O�'IKbL}ܷ�eN#7�|/��ϋX1U���a�>ڏ���+����>�|���>g����1��{S�6hi{Y=�qv��~�T�m�"]��|��j�y\��hT[�G{ޗ�W�L�rmm�y�}�-��9�È�܅�q�*���A�T��m>]����.�zæ�gu-��y��t+	��w�d�Y�}�;�����w���=����B�r̀a����m.;z�q9��$p�Bt	�p�o5Od7��Jއہfz���e�Զ�C9�;[�J`lt�F�
�|�^.���D���#�þk��̮R΢ӹ;�iܨ�*a;r�G/�,���=���9f��F�j�K:��}�[��?����:��;�5�DHt��{k�o-�'.-���!f��*�Q^����K%rۍw��h�U�܆u�Smj";���΂

�-n @�]�K��˚��Y�n�,ú�l�>�CuwL{.֍�20V�U�zJu������xT�D\�I*h<���K1S@�u���}��<����v��j�:��w	��s�ж65��pe"�
+zS�NpF蘱�ӷ���sQ��3��]��fp��y��N��*<�U���)�����Oi|�����p7��S�*�vn�������o���2�B�4^��B�oT3c�iw+�p뢷�Wkb��b�g�:J������OjS�5����ߑ�������?���j�׊�Y�t�4O�,��Uf1������\i�����p5h�-�(G9a�����-Q�k�{�ŵY�}Z�s�5�,w�zݙ�$G�q)Sn����Z��g��R�V����K���6*-���7��ec��vk62N����R�jg$�A�y{]_Y�[��F�����MnS�Yzѓ}0y�c���g]Z�qڽn%�VD�X��D9�K'�>��4����^0I�ۣA&�P<�8�_+���p:ua!�xQ�؜'و��|\b��-b���z?�J������'8f}<�L���6�y��5R��|����˝�!M9�����V�T�T6V�A��t�=I���j�;��XyT�uJ5������w|3F�]�z�w�)����bۄĪ;[mu-��1ŝ��;�~�@j��'5{�gc{B��S�7�{��@>�^=O�YZ�%d=)pˌ��n��Jr�-S�<��)�og~I��v���\��%ܮ�	HԸܽԭh�����Q��ƥy���j3�Wޅp�uFy�J�v����EZN����2�2�{�P���"V���2���\�l�p��o���̜�MF:�d��j����Sq�ф�)�[����W0��&�v� �x�Y�L�y�aj�Zq2>���=�">�u�C)r��'+�g`�j�
y�Nך�r����j����l�l��}�v���3+ƪz/���Vn�.�wΚ����Y)�7���UEnQ�wT�m�mu&�;7cf�(�]�Q���W�F�,/_�7��͡�F4�����K0V�g��j��92�P�C�;�5Bۛw2[!C��h�a�q:��9�5���@T�&)FΗҷ�K�peDnB�k)_u�˙�D/���l�u�b=�}N�k� r�T�D�k����g\��ռ��X��}�¹�Z5坊�������Ϧ//<�Ý/V�U͡�w�V1������5�Sw���)�n���S�SY���Ci"��U��p�>{�R�O'J{״|y���[m���h*<���q����Q�9a��|� ���<s���[jv�n�����^����U�ۄ��Y���\d%0w��Z�G�T�aV��^՜{�6�Y�gU;�\&�����^�_0�(gY�O׸9.<7yӨ�~�+ȩ���5�1;ߖ��qɝ�X�`�aUVn�F��sŧG���*h^�:u��t�}��M+zm��d��7f�XUSO�������r6��d6Q�z����1t�	bUp_u'�Of�ɕ�ҕ�{1le�mÌ��J͞�@@�n�nL��P{Yi�%�'Y�u7k-8W-eU�6�o��f|�\���"8�ȝ�������ت"1ሌ|�P�F֍��2�v���2.;�T�S���� h��r�	�3&��Em�C��`��r9���b�����R�	�Vy�-P��m��%\�E��v�-ͨ��q�����{��c�ܼ�g=�l5���SOSEM�~�s�֟"d[�3"�X:K]�`�w�BnT����_ n��֗S9��ԙ»�뼉⺽r���v��є�Y�)x����ӘRtv���LN/^=R���nf��kz҉�{P��=I�Ts���XU��uݓ�'�"DAGu�J-3�8z��ѡI��ۍ*À�@C�c��૭Q���.�X����A��=/q
�0V*��ΰ�jKHyWC��jR#o(|�=�ۍ��z��[v�q�=|E-����8�.���Қ�����=ו}�y�w{�yr!_f���'�;��ά7�k-���F�
<���1K��,�����@�m7�^v��@D�_܋�W�Q��f&q:���+y���N�,3��WR�r>Ε�`�z���@�7���G� ��to�ժ�]4u�G�f[)�f���@H�9v���Z�gsC^.d�M��Fv[��N�1φ�L�����}�o��k��J�M���� H��]�]CҌ�fK�'t:-��!�k�*Ʒp�u�(��������V�cwL�'5�O�y%H���b�]5�-�[0V��U�+��.7rٕ}%�؉��ռ��V�g`o���]��[�yYYʕbQӼ:��r7Y����{��ί���t��Or��:��{�١I��E�ۊ��V�n�P@�5ح�l���B�a�H�%���QP�:�-a6�;F�����BKn�t�1��o2�
5(�Dm��m���*��# a�@����j�+�JS%8 Y��=st9��Z���PAYn���_�d�3C��vA�%�5R�ڝ���n��.�q�w��8�f�;OD�	�7��,[��e��S
�--0B�igт��"��p����o6+u�u-I�È8��jȖ-����\3�P�Cj�u�N�v�%�ݨ"��4� ��ݘ����	f�{����D�Ĥ*�^���M�V�⨷Uɲ������|]�����{{wDwR�Qc׹>=A�N��ZZ�M���F�ޥ%b��ӊ��N-� &*��vz�p��J�ǘ���/�W]�-.�k$����5��$@�3��
�\R �<+���J��%�|�o-D�W)ۗ��Wa@n�|�:[��R���K�L5&b�Wܭ����>j�მ�J��Z�S��R��A��|�&л
��˖�Ui��;[DZh#�RZ�ӗOjV��v�7��Bo)�uq��b#/����� �_�(�ΩZ�a�u��5�V9eM<l��Bµ6��� ]�ٷy��|A�c�x(Df�Y�)N�m��y���[jSc�i�]���=�E�^��`�̂=���n��A4��_�6����(L_PQ4jڵ(�ֈ�l�m�m��E�Rэ�aD,b�V-B�h��
�2�F"+-�RUA���b"��ȕ�������DDEX��*)F�VQ�E��(�"���(�mb��*EeX�V�Q�մmk(��"V��Kq�`�D@QPQĪ+�eddDjU`�X��E*�
P�T�FȨ,b�D��1�-�
�b�
-���*��KJ,�TBڪ�5,[KhQ1�EEm+�U�Ab(���Km��m��Q[h+Z�#m��#cEJԬ�-�V�(�k*Ym�X,e(E�Ԫ�4��h�5Q�jX�V�6��mA��
���JTjڊ�F��V���Z�Ue�jҠ�R����U�YZ�@@�?}���]S܏xi������O���k��K���[�a�v��}i5���[+++3B��z^i#O�_Y�7�a2�k����Y�zq�5�����{��8�e�������v	[��U��N{��������#��s5��~��־H>c����ƌN�^���;(�
��ېe�Z�7��uwO'�c�3ڝG*���5�2��.RV��7�'���:|����^�y��7W;�!�}��F�:�z��Q�{�j׉Үk�z-��=8v���ߨ�Xf�c�p���i�.V=��G�S�ڃ��R>0?�R��]P�[AqӊG��e��S���҇��Y3X�����'�^������ߋ� ���l�/k'���+Zƻn�J�U[�ӎԅ�[��ɥ��8��(n�<���v�� 1N�/R��,�TY�VuU.��5��"����������r�Oob�|�"OA��M�s�gT����U�5<z�:p��E���z�EM��[��-�ܤ�l}f���KyZ&2�z��kx����8;o���R�_�hEa�����z����V���#����C���m{��z�l�ERU�-fV�*��{�r;ߌU��2�_s*��/]�F��}��v8��']�*�C�{P����:�C�Ч���:���oMX:�iR�7�R�{��&1s�ܕ���)_�9F�p7pT>o/M���or����������ɱڔ=?;�P�9V!)�Td̿=󡕓9�ι��s���9Ȱ�-s�hX�k�uuxʅ�F9�W�q�Jz9<\2k�����B��ڄ��z_|�!P�G'G>W.x@�(�y"w�眚�}��&/P=���sY��n^��1$��5��0�ki��S�/+��X�a��j8�S�W�������׋Z���V���n��8.�r�{�)Gu�W�!yS��k~�ߨ��W�r�x��9�Y�b��С���\�qPv����b���4!�ߗ���@��*���(�{�q�ڑu�ڦ���9�Lc�5�A?U��t[�\b9n�x�(n'�W�Ѝ]-5n^�[�e�,�v�!��t��b��70P�F�.M�p�K3.Hmi�kqC��'(��5���T�.���KQVc���'�oUu��v��Z�-��B��;q5yWlh�|�q\jҲ�#�C�PNZ}�Q "YO*��\�[�N�r��*��O���W�}\;�%���0V���1�+�T�QQ�kA�i���K�U=vk��~��zaQ��ջ�Lǎ�R���y�S޳��N��6��{�+=;�C�FaOu.ϐ�A1�uȭMQ�B�kCg]e�{�Wk�f-�f��5���N���<��N��S���r���B������K'�>��Q/J��Su8�DkGk��&�[�*�/�]�u�D��m	`�h��tV�	@�&0P�ݺ�ǭ.�2�����)����i������<�
tlvTI|r���v�f��1+r� ����a�o,�}*��CM+�|;����N���U�K��5םB�Ľ���*[^�{C=X�*ۄ�~�&�IW�4��_�>A�ۛ.�J��+ۑ>5��r��1mJ������2�')wMD��3z:]|,�]`-np����,O
�3����!���ytT�Ӫ��2erk�:M�-��'�%�ySݨR��W\x�
�[|;P��.��G��2���N�W�R����ok�Q�V�n��K9ie�������|b��m��y���X�}Ju�{�c;����o6��}bԌK�����+�}�t�ԁ��:�����(��O���-� [�Ȝ����/@��ӛ��y�n����y�5;�������hQ͞�����[�@��u�7P��w�+��ѓ[����Hzԕ_&�mw���-��j�$I|v�>~{+�/^��@Vą�]���<Oy`/�V���};��;�ڼ��At=%�����֫�y�鯯TM�(��x�s�wSv⪒�],�ߋ��<���mX-���+j��qM��K�{zz��-���UҞE��Źilʙ�X����א{9�m�d�]�/o˪uw��EmA^3���/��z}ލo'����O�M��w���Z��vͫ	?���ݷ�3�ؚk$�g�ҵ�֛�Cy���K���ɣzh�i�k�s���z���qXڼ�uV����з:{E_+�8�@��*�j�'J�b���T��ҁ�����ks ۬ѷ������e�F������U\����ݔ��y��ʹ�����IЂ;��7�n�kUNݳSW[k��q�؅q�W+M�U��Y�\��s��R鶮�	Ef%��w�����/=^��X��f��P~��T_5�����I��o�{0��v�[J��3,���d$Y��6����������A.��S�F��5k\��1U���Br�_�!)��L��Bj�"~]�xv���$��&A;�lܵ8���p�S�L(P�� �:�q+^l���sHފ{C�r/�OgS�=��Mp}/��͗�ԝ��r�]�iml'9�̽�N2�P�ݚ���
�H��ӷ���y_͞�&K��2�UB��,���|4��I�c)y{:y8�A�|ԕ_&����J�lf)�4�j5Y��D:P2���Wj��}�A�������!B����pWUܙ�[���Tg����h�p�Ek�.ұj�1��4].��}��Hi��	D�Cr��t��S�e/;�S�mh�[Aq�8��"����WzZo�lj�_MJHk�U�oK�܋!�>W]���.p�d����q�\CLE%�vś�i�z$������F���OTtA��d^�;��:�Q���x�띩�E��#��U{|�]Vm�Q�o�}Ft�Y����h�0���r��y�9�RUA��lb�bl9V6�Q�F,;���u{�J�ԯ_J����T�Ţ\�� ���U�@u�_��Ok��??19���4+�Wt	�~��~O�r�3�o��tK�5No˛��3�k[�+�3SZz�V�ku']�oc7�5�� �҄�}9�
:��O1�WO-�%�Ӷ�VZ{q[9ͤ0�����ۄĪ=�*��_%W=6������A���}Ւ\Ӫ.� z�'}��=���hHj����`U��j�w(&�ѵ�����]��慨�M*���녣&�Ue��BS1#��k ��f�*i[����}Ujq+�q�4V�����Y�W*z�B�ɠ�V�!���S�Vo<�]p���ٜ|��Z���o!T<��
�<�e��gR޸J�<��w[8{Pc�i	[�����YɌOe��P��@��80�>5��b�h:I����]oPS5��<���Ԙ6��k~����ԧ@	�	Wn��⋎_
�yH�tS�(�J�2fQwM�mtٸ�S����-l'@�oF��,��Kb�
�խ��R�]�����U���woT�T���T�hO�pG�U ���O�}�5{�TG�Ӻ���L��y��h��[�1r�mI�N�H��#��u�1o�U�'9`{"r�v�L�_#dO��Yp\w��O2�1r��̷�>L�ߏ�q�+�mHU��O)�#���ބ�ൃ�E/~�e�}��!�,.D���z��7��S���q���Z+ݑR3�]���m4��N�ne�Ԣ��g7Qy9�.��/�ޭ�1�|��Pj���J�
r��}��1����UW���/[�����y��wM��6ڷ|���#k�1p���FZ�@����y�����L��!x��J��{�u5(]�3^�Q��.�z���X�6�,[k��q�J�J��j�'�<�F^ŶR��v�:�\�+-K1r�qI�A�z��lOQQ�R���B�=�������Yw�6u��ƾ���ok⭻�v��*��8=ً�*7V���J�}�c-ԉd;|�S��V�ڙ}��ul=�@�F����#�]�ٔ�J�s�����L�E�^=;�{�"^u5��Q]�j$�z��\�JMa���;[~�y{0��ƆwP�9�mVLl�\�����|>�
f�5Gf�I_�L+{4�J�A.���N[�nU���6x�o����՝�s��.+K���]�]�it�2f�g�5�r���b����uQ'&����{�Z�µ�B;D6��=w��&�whZک�Y[��E5�J�彊��tu�h2ȟk�D>��D�̰�e�Y�8�	���7z�B�E��W[6�������&۞vi��ǳb	*d��q�[���ug�w'���ƞ������7�)�u�6G6z��K��)����}KPɟ���;����c�ޮT|ԕI����8DƸl����SV9쁖q���fo�{Zv�[���*؝��S���(��#aVW�]��[�k^�G_��u"���X��Vj����$V���{�]�u.6b��Xի*�l��9Q��dr��HTު�Hb��3q�uz�f<��GLW�-Z���<��	�K��<���ev��0K�� [υh�=%������0��vp��wt]�Y��S8��K�����O6P�fm�r�=��[��s���ӹ�m�������$��j4v�z��꥛�C��nr�M�������� ]���qp����o5��'���i�6*"��y�:���_����;�vڬ��:�(\Ѯ��s�)�p��B��TC�S#��e��������l=���]e�;���[:�)�\K�n%rK'���pu<�]������wS:'ܵ\�/B�ok���mzX>���y�{.�:�i=s��Yy}�{�7sݙh<KR;;}��-��06��@��)�V�odsP`����4[��q�[�\��DrNS�s�o ����ȇ�U�{t������f'����o�h��lގ�Lj��DHtȑ��F���� �J�kQ.�oOm��٫l���ܤ��)j��bf�z�@v��SӱE��ț�!Φ���sΛ�iB�q�}���o�VTr����%y@k��Ež�e��s�<�%��x��#8�՘M��n�� ':�x7!A�L%�,�RStww+�_^�F�F2�������Fa2�9"����<{�F�����C�A���O��F#�L�b���j�@-��On�>�E��������+��F9���x'p[�ǍA�\:ா��/m�hm.�S�H�ui��6=o�Jܼ�V��b�5k�\r�ЮϹ��#�:����h��� ����hF�l����E=�ՠ�bt�۽�f�J实����7=�N��w�m5��7_k��P_eWV�TE��bze�Q����9'�k��o:�X}7����^�늝�kǝ�t��T�n�&�y�ܚ��_���=K���=�;קǝ��^,E�=�A�C�N�S3ʱ���#��3���;g�����eE�B��Av�{�v�5�ڨj��]���Л�k�J�ԉ���_Js}J������Y�[k��i�*o���b�w>u=l�U���Y�K��
:�}�E�j�����J�2ʷ����u�U;�2c�^,m�,K}��]x5�eݗц�=8�5��^�ɪp1��=�z����v�BScz�Lwh���t*m�粈
�B�^�3�mv֮�*ks�G�`B��e�� L�7�:��E�⅓�RhAW��u}We��v�w�qa6��U.g2���݁쎏�U�8򕐴;�hq9��vgu�T$��HM�\G֣<{��%q]ò>��^i�aΥ�rl�u4K=����~]2���k���-+?ivr�Km��:W�g�O���n�2��H�]dt�O�[Fvr�����ɹ�pax��ŷ���'�(ի�W
뜡{���|�F�.f�fn�yٲ�ow�R�I��h�Y�ގ���]�)W��l�ۥ]4M]"Ҳ��=t�0�gc	o�[��:��f
q�a\&Lj@ɭ��n���[�o_r���@��,�{]�{h�A'�0�j��w�^��}j̟s�
�r�7��"����2��J���Z����f�++�hCzQ(������+b|�=�$ag9lݳ��o��g&)�u�z�h'd9�V�{����M}}���j�����8`�7�r�U4.5.]Z���|�
U6R�x�R�J�2<K,�n.�C�R�^��š�)'�> 7�8��նt5���m�S�-�T���\Tق��4uN����eKbA.�%K��=*�d\v,��&ZV�I�n�����_�t3o%���(���ϳ$3X�.=r���:����A�!7�c\�Z�2��U��Yn�F�5+��S.LW�]�e��+)�C8�����f�=�䅬�t�p_a�5|�-ï��\4U��b����+NR\Y���j�Ȑ��r��9��y[zVR��E�8�[��;,�ޠ
w�`��֬�n��h-t�4aY@��w+.�g==�!�XB
ˊ���ƹ�u��3�}��AT��>���p��3v�K*�M'�EblV&D�_[�QtK7��m;���LzOi��>u�g2��n�SM[Oue�ZU�����Y�ڬ�4d�F+G^��c`Kt x��L��%4� ��%�o��ȧ#Z�]t�]��j�Q	^C�s�h�˔�M�{ȩ��(A��B�4�/���nX�[1�jBd�lYΤ�R���5ɫ�լ�Yv6p���=���#/^�������v�Sq���5���N$�Y���f�)�ٙ~3=61�m�g��_]��sCi�Jc�8Tg�Ǖ\h�^7C�/5�i�y��y�X����һ;��]`'0��Tp�lx�Y6���q��,������zq8];��� ��`��ӝ��rC��֧���ȕg�y%a��+Z�t��T}��뱠e4�.Sx�Oz˕j����}i����e�H짰�s�C�#
 >)V+o���EfA�lQv1ة��I䳧-��A����߬�C5GQ`�0ʲ�����*���d�G�+�a��D�Cop0�w#�f�ٹm�� -V1�@{���h��B�R�V�@bMW��v5:Ԫ�Ss���͵�@r���8y6����������Qݨ֊֊",F*$bF�"1QDcH����AP��ҬEV*�1��5D��1�%J*��ʕ�"�UF0QTUTADEUTEF)Z����D�Tb���(�Q�(�E�*

����XF�TP��*ITB�Ȋ1m�0E�)i(�QZ�`������,E�b("�(��UQ!mPU�U**()Z��D`V���QX��X�-**�b�,�D`��m+P#�(��FA)q*�1UU�������� ��UPV*��*���`�0Ub�V(�d��dU��""�,X�+��D�T[������߶]�[ڳ����Ni��}Uz�V��w�5���*�˙�"�X�Y��D	��]]�&�]K,x�,5�����_��-3<�/k��a�]V�OF���w)l�U���jK{���mdv�eM�8USƠTnm1�]���_t�Z��<�>���eOJ3 ���I������w3
tE���1+V_�ve�qM����7��:�p�M���W�l���5�8�Ӣ��0�~�Jܚ��x+������;��u)tY8b�7;�̶1�7c��5�q�~eP�zU�����'#�D�Q��m'
�6����*��OQ�'�l��`���Ux�Lt��s��1j�Ț/R鬝��&�j���'���u�BX�8���ɘxk���躞�F�X��z�+���V8��n��t�S�2�� גZ�V�9~fW���Q��iFZ�O5U͠/��c�a�cf+��,Ք�'�����5��]�\���qU���b����l���Y˼�9Vv3S��c�b�V�N���4f�K���թ���N��'����@Y��f�o�A�&�=�ؼ�F���>|���I��a.,�G�h<����ne@�y�jf�A�������]u�v��3uW,���4gr1�/%~�qq����@h��8<����g,�@eZr�������w{_�G�2�h��&؞Foi�G�;C�\:m�8a~�v���:Z���x�'�s�f�Ms��I*�.FZ�?<�A���y�m(��i43\�q��>]�)����ʵ�uc���ڬ��ok
&�i��U:��P��췩�w�<�g��-����<���;��k׽9��5�'��r=rv
��N��g�|�^.�of�i>��FJt��=m���99���[��-k�m��F�;#{U�ުq�2����}9�B��,��vr{E`w��1�R���!��ܭ����U�{wP�C{��Cwa,�b��U�i�J���Ny����u.B���C�`�yw^��w�(�����rW;ըR�˘�MQ�|���B�wS<0�����l2��Y�k��9������&OWk�]�kQk_��Z��P��?sg���2%r�n�*>ݭ͜{]/on�H�+�o+jc�+r��$�/�;��i����c �&�@�.l���a�������t��	�V*���C,�h�!�"QE]�n<�Z���I;5���-��8�ǿ��B)���I����y=1��aGιPt�T����J]'9"��&/f�Գ��b*f��{�����h'�)v��; ʶ$n��ޘaz�^�i*�s`���ۛE;�cV���.��P_`�Y�^�Oj�]JV��\�yVi�isJz{�Q�^���>;�ՋUF���V(�e���J���s[W37���p��g��}�6yA�/ ���6A6������Ky����M�i�����Q�j��;���O�ܥ�PSŭf��-ۏ�z��J?Y���
�-\膪uu�k.MnS}PU�\'��f��Tm��=�y^�ި��ғ�ޯL��uE.K���5j��{��97���0/.B7�^f�s�ZF��9�6ץ�-�j�J���i't^t9٨ي��|w�Z���c�㬮_JF�U.d%���\��od=*H|<�Pu��8}�ԩ��|�oo(\φ}��J�E����i�O%�ƴ����\Nܭ��[9«n*�:u�t/r�"*#:��s�YX��w�:�;��]��eN�k���ҮZ�z��;a��oR�<�6�� H�ڰ$�y�gꪮ2{w�T>Zp��>�Isasq��T�r�X���:ew��^5� OS���Ye9��@��q����1��3�R�-q'���c�}���kw�*��ƍ\�w�	5��6)3�/a9�EΉ�+z��L�N��V���Rv��{��t��T12��\=��!HF;//�2��[��T�yw�趨o�F:>c/f��=�<�܏e���������y�E��"��[;��^Oi<��ڧ��}�:&��d�<8�<qN��6es��[�����٥�#ix�F�WSʹ�[VҨV�K�Ik�(���M�7p����:qޔ��s��TV��)�`�$�j5��N�r�����Y���ξ��y�"ߗ ���mV>�um�����.iN׻=�3��]G��������RͨO;v`�(X�,�7��.';��AQ�돳�\׫Z��<��vM=�����M�:��ZT�t x�p	Yæy-�Z�pz�q1n�y���~���;���
�}�9�V�v���cy@C_; 0/�����y'wI��1�u��2PK���K�֮ׄr�Ը7�vn�Է7Ԭb��r�T�B���3Zo���ц��\�i�PJ�[�q�E�=_\j%A�u��d��O`:y��Z��r�>���jGk�����ox��B6���KGFږ������C��R�U�ch�U��Z]Rg����V�m������+�-�@�",f�I蹿A��hҠr�,��o�NG��cͮ�$�v��dúJ�\!(�|*Q6�ڦ�bm����z{eR��&:y��N�%����R26Kݱ0�`wv����P��ռ�%5��א��c�u����g�<ʙ�9�Ԋ�ʞY�ˊ�q��<6 �ڃf���5i��Wɇ3u[A��]n&�*������=�SPaS<(��񥷃���c���+{w�M�[}ë��Z���Q����>�S8в9�֋�4���Vܑ�'������7.��P��N�pH&0�C��q�����k�TY3O�:�+��I�H��qJY��X��z�a,G�2Ɨ}S1��7�����r���������{�v�@��FT�-EN��[�-(��&.�]h�xb+����%�h4���z����Om�9��,[�y���㺵�ؽ���t�g�+��uI���{KU=Q{pZxs�A����Wc���^e�]��Q�������DV���k��~�J]�G׌���i7��Ыܼ��LV�1�+�w�[G��H��Mh���q!���P���[P�3��n5�����~'!����}�ro.�5=����s��내����4���jY쉜zn��Wp���a��e[��g��_ouo{�T�r���?r����L��q����h��Af�"������~T�Ҽ�}�nq�n�L�{/�z<}���2xz6���Oz�8�>���v�>D�U�u�+7�E3r��o���a�Yb?�:��O�~��@�ӚEEχ��(>��և��3�=��㐟�x�<�G�ລ��e��5��ډy������揠䁻2G�e��������}��8/��L{��;Ϩ��XT���P}�[z.9�G*�]���w��5��T�Ȃ�KA-f}�<���^������>̀=��{O��������hġN���}`X�[|,�k"�F�O�|8ݬ�ă�6mvw$շw��^vn��̈́N�Q�X|&\F]�aL]�Kg%3no]7:R�죵��K8�A32��{5�gv�'p�qw2���ܻ=3����YFM��P����'�`���.^���и~�MÀ<�I��M �}d�b�0�h���]{�j������*s�~�'}nM�y��=���n\�yT�R��q0X��#)�i�#=���L���V�y7�#�ei�?
���L�9�3�9/ho�`T<��p�4xԱ�o���_)��q�Y�P<B��d{�s��|������}>ۘ|����c�T�+��^� +�%��w���I<?n����Z؆�u��gA���ǯ�N��9.��H;.��{���Xc6���5˔j�=n��K�;Q�d�}�m{��{����m0�%~��n�|A��Ϙ�o}z}'�B�d����扽�L}@ �����������𼩏�Sڼ�ܫL�x�)_������u�(���k��u�~�87��� ����i�X�֍R�k��?q�ݰ?&gU�y��c��߰r�%�G?_��6�����d�U�{|�|�H�7��*���2���=�����\����<d���Ǣ7���V7>k��o=O�qط;���]�dG{�Q�rKf��+�P��˟�Zh԰$/��z�wh��9fN��~���aW�Cn�rY�3�,o�E�֭�s����B+;gR9E`��I�Omܨ&�* ���.$ ��W\+���AH�(�Q��.XP��n0�U�:&f����r�k
v�����J��t��Y���
�U0&���\dγq�<Ϋ��8�6xlGyי틗�Q>�,�w�ޕ0�}W����j��j^7&�T̰2����Je��/�����ў�-�6��D�eQ��VJԒ�w�'�~2!N�q��+�n	@-���b��N��&=����x�����R��Ž�9^�>\�0����W��YR��BsQ������ n2Z>�/e��S���W�ouWr�D��{Q^���H���QL�����w@\?W��Ȁ�Jde��/r;,��C�n���U��@:���Ī:��}~��L��B~���m֋�̹ R����]�:|/�Uj+s7�ӛ�/�}���<���i��c[�1�=T����~�>9t?e�������!=�B�'7���X�r��N��u��2�11MVѽs�܄����'�?Mx�����`߽����e�5{O�Ѧ�A��H�h��7P��+t¸�WI�/O���Н	�r�|�>&'#o��׉Զ����΀K#�T<.�{S�`��3�3C��~M�x�{�	~���_�Y��:�ە��x^k"ʯ�)�w�%����|&�NWV9����ac>��;V��Ջs�CWs��Ց�kawl��<�u��<cwn�.�-�i�CxM� ��q�K}g�t��C��V+���Rڟ��;z�,q��W^���ZZ�����0��s�$X��,��U�:k��J8O�����k�C�s�Ea�S?����*}�4��P}3q��1S��{�Z�%x�+}�q6��:m��C\rr��ro]��ݼ���GMx��'´���o��:Xq�x�V3��E?^�����Ʈx�tx��������Wg%�^���a�eSQ�ZX����t<U#*��$^%Mʞx7������E��Y�߱<��{jY��%"E�;3	�}���ɝf�g�1�����z�ę�驓��x^b��K�>�_��
������Af�4���6����z��L������;�Tٌ��nN�'�Q5N+�:����L������V+�ϊږ{"��ve �d0%��-n<s���;�1����%�´��}~W����t���^����a[Rˀg�= r�>Ş��諮���)����9����se�_>Ո^7���gǳ���da�]���m:>���'=�]��܌3'����_�Ð\�϶|<V�\K��C!�i9��@�2���~�_��I����WYcH55j)%Y��lud�[�[c��M|�8��k�n�;�*�o+k�v��-�t����d��E��	:è��p�������i9�h�}�1���3^+k9��]A�4Op�m>��Vi���0�ǤƵ-����\��U�;����D|�@?�D�ʓ$O�m{N���_	c��$|2#��y$�р�L��^����~�Zj��T�k�Q2��@|w��ӴwK���F�����@#X�K��o4TQ�宭��݅ր��X��(��gö�3a�͒zrH��������/���
���W�ϓ�Q���m����	G�Ώ/�&��/. χ"h�,�`YB�fkN���ɜ�P�鉭�4̮,{�O3#ؽT\��Q�o�wϙڜ7��!��~�K,M߬���N)'���_�g���X��K���bz/m�P�g�<6=��c~S��k��	�������o�juy��=��ܕ�����.3f�����u0-M2����K������F�9/�+��o)��i�	��I��V}U���/��eVy���~���;)����U�3ށ��"o�q���B���/|�m�YΙᇦB،Wp�#&wҏTj��O�g�W�߮���w��������~��>x�E�w���5���68�`(�}0�r.��:6�SR8tj�KP�O���8�߬Z�D����Ҫn���U�K����-��X��oد�Υ�}��Tt�r��F����:�lkg.-0��v���Q��=+#Y���gF�;vJֺ��68(B�.�݊4 ��d�{{җbZe���Nҷ�t�^r�1����;%V�IR���2RZ/�D��$�VgTQ�z;BCB�j���d��ZN�@�NP���oS�ǳ�[�XݻH���l��d����
eڇ-�4Ӕ�9��dnv�� B��0���Yʾh:o�j�":AR��j7��:r�>���@��7�ۣ���	Qε���Gș:��K���j��2���џ3-�n1���fO�$�UC�m��5@pB�]�Vc�@��h����p��p���d�7hW1����y�@��z��ur�(]fB�����
�� N�t�����.ʖ ����y�z�Q]�q=�]on��2��E����!G�����n���{��-RX� ��yR�i���ΧU�q�豭�MJ�����+l� ��]`8h���ճT�»%ugqvfZ�k�vj	�m�r����U����m`��<�D���r�'�0w!b���k\��e�|�wS�g�g#��E{�hV���Ǫ����\��I۠�p�ĜvuamݍZ���/�nt�4��z��#�N�v�ŗط����^J��TRyn�1��]���f���4��kW��Z�[�c�dקX�Z΁�WkE<ͮ��Ƭj�W9-���t^�h��e�
���5d�e���ZZx��]��D�6]�[V��6�nD=m1x�<�&���w@c;
�Bم��D�ƥf;�7��^8�ČV[���Ĭ:=����ǖ�mh��DwO�ӆ�ǯ`�@)P�y���;]ۄ̺@M� k����/�D	�	��/e��U:׮e��|�����մ��$Գ��u�8Z&8�}��+h-	n0�Rќ{,���k��m�FD�)��]��ֱdܵ��s�7�x��B`6�j��j'����@���e6$�o	V��g�d�yw��Goh$g��ך�f,�U���X}fD�t7F�ˋgT�.�gqj���Wo\9]ɚտ$�*Sh��JW�PkUi�Z*��U��:D�{A=��>��y"`����\���8��q���t1G�)�r�EԌڝ���fh�R��q�Т�/{�C	sGK�Mm�9��c�n�(_?�{��M��s-�KB���"ͼv�Dj��1�M1Y��B� �[����x�`�ۗ.�E���9mZ=0�i����F��HR�xE��	�t�|\,�t��ݧr�*|;��o!%
�}�[�� ���$%Xq�U�rфi�z�mbs]ز�ZS��DmUӋn]ZbP5��wNئ�^.�Ԟ�����t�6��i�ͬo6��N��񣦘�e�ʨ�[>�;V�K;�X�
����DMҊ �b,`��UDQY����b ,EDb�B*�YEPY��J��%J#b1b�iR*�v���,Qe�EPQUd��Z��dQ�����-e`�D*X-edEH��bȱ`�(*�R�
�؊��* ����PF� ���AAV(�JʬEEDX���PUX�B�cZ�"*�������E�l*�"�",TQVU�Z�U�"*���I�T(UdPX�R*"�F,H�**��AT*
���j�"�m�`6���
��UEEP6��""�*� ��,Q�ĕ�$QV�bԪ2��}@|+-�մgˮᮏ#p8����,��M�k1-�xs[�Վ��S��l��\� ,X���ϑݱ��C�|���f��:u�Iև�O�����������sA��^ӏ��Z:��(�c�q��{=$J#b�^�4�ʧ��=xr��9����@Q�#.x$n2�?z��
|Ό��.8�>�]���3��s�jn�*j��|9zl���� �m�Hu2�D�F��e���b2�1q��=w�b�]��j]���r����~��o���<O@n��+԰������-#C}Wn'Sz�<.���;C+ۇ��L{���t.��p�9ޙ�h�����>%��X4̻u���r��[����C��I��\uyc�ߍ������������xvJ���9�?-��iЊ)v��{v��]�k/]Y�D�wNzg�m�
���w㞙�}'"%� �����^�'"f<Eu�{�3<��xp�y׷��l/1��~�E��"�}����iظ���S��yO���=_2�I(ly?F���gj4�MI�}'Y뛨�ͬ茟�_w:�f㩏'4O�R}Pߝ�_{��z=]u~����.��^Ctd�#�5V	���Ɩ�+Ɠ����X�,�����?���3��i^���n���pL�5��qu 1���7��+0҆��%v.��S�/5QB�����eEVo�!@����3!�E�CU�k{�����Od��C�)b\d��ii�x U;���uoh��c���"f�@�\v��I-&���4k�Ȧ�߄^]�Qy�޻?OV��������{Zn#K��r�IM��U+�S�,�2}`}�~�=�l���p8��:�_���/d���t�{�V�+�P���7�U���K�����-@�^��=8�v���#}��/�9�=�%��b�u~���.wk��RH>��ی��Lj!zTOz�l5��/��S�\v�3P����G{�Q��L� ����53��7��NN�o����xʴ�t�Y����8.��y��O�����d{73&}������u⢌w��*����7L
<�~���ڨ^�����g��C�ݺغN�7,u�/V�=����1���C��Np����n	@-3�(��x�ȍ�h��>]^�����M]��_G�Qɧᾦϸ������^� �e����77�zhQn�9�L�jux��V�k��v������ϣ����H��T��v�tW��z3�.O� �؃={$G�|��;�!U^Ơz���o��zs6}�P�+�������q(���/�u#a�S���)�>��?T^.v��+�o�T�:��p6kx$����(Z�h�>�0-�V=�ȞG�,��J���,g:��]�8_(OT��c��5�Ws+%:Zn�M��j��)go���OB�T��P��̼7�q�Wg�$Σ�m������n��W��ՉNM�~���ƪ��1Ny�}+N����m?_��U;���雟z�.y̱�W�mح�҅�1�U�t��K�ۛ�}��c~��h�>��iՓ���_��;ѽ ��Q��͕��R��>�vt�n���(��#�7P��L+��t�O����αt<�:���:� �l�h�URϾ~� Ué�d��O%�3a3y�P�3k�G�I#^x�N��y���˨�}���~�E������c;S���%����e�sq�W��K��kE*�@y���6vP�L�6��ϛ��N��#p���|������*��?G��[���V}��Z?,�!��z�nF�n3������=6΃��[���j����^`Tŋ�=X�U�߱���Lz5�ćgES_d֖/&w�Y=T1Dt�H��}M��'�����<�&�?N{q��O�3�[7V��UC�WL_�3��>	����!��5|ћ����o���Gڝy�߯���yhhϟ��5ѧ7l%75	��\;�)�;PY�!� U�!�~0����j���~�3�*W�F�����|{����n����ޑ�VU�N�P��׼�Y9��#�jd.��b���ܮ���� ���ع����ݐ�������9cs{�:�z ��࠷/���c�bE��C�iAe<�P���5��
Ͼ�j�؊��������lxj���TY�~�)ٞl�Q`b����v�n��[׎�����]����+�d�l���>+�{��}�������dUT�hx-��mw���\π���U"J�d۟3���x��7�Hǡ��o�x����n�̧KؼMq��ۊ75��RĝQ� .>����qJ�Q+�a��x�l�*��Ы�]��J.K���ۆ�䛛�Ss�[��<�gfD��SP��\����&2)�{Hd�#,{ޖ�Z-ǰyH�y[�lk�]�}�}���i��eT`<�M�re�Ā��_��>���_�s��[V�bC}'٘�f�:)�ϡ��oxW�t׍���Ȃ�@
��ze�>�f�q�D*y+Wޯ^�e�������ˏ�M�����_�Lf�5�7΀�8�G�ɒw����܉�ŝ��柬a�t�Y�[�B���87�;�5>�d��c�^fG�{�S������ǘɛ=��>�R���"�ZK�����#��;H~������'Ei�s����W�^�x���C�{՟��i$�"�AǂXƮ��Z���_l��:��^�f�E9nV��H�I+��;�f���7yv�WӫqBs5�+H�>�¯��1��eu��k�]k�B1)�˹��5B���ݼ�k/��'7�s�Q���u%�bcyJ���Wf��	����L_�@��q'���;P��ŋ�٭:���:�����_z�d-������L��O��qʐ�q��Z-{Mw��:�a�ܭ�w��7�u�л��i
ӈ�y�W&o��h���/_�����v���/e!���Ɛ�ǵ,�L���!oخ����r��{�����z;�ߍ���*���c5�_������z�3��{�g)(�9"WA�ȫnc��HZ�ġ�=��q�>���W��4��s��~-���1��\��bġ�,e�Y�9��3�^�DN��T����E�	ʔ=p׽�VJ�3�=V�~�h��}����c����\?m�]�)�Uz6��ǔ'�= %2G�e����^d��z�P����:z�;�O�Tw4UjS����$g���o�����zwT���Xp���f���ɻ���}�55Y���Ӟ�4=����cӴ�y��}��e���Q��_L�٨�4*��ګ�>��_��9�غ�KW����	���J�__�sӕ�������r*U:!���S�H�/@���L�iBj�wqIZ31]"(U�,�|��(��M&�uA�oP��c.����es���r��Mg5X2�F�5FTvi�/����͸��|�st���O��\G�/t�!.�ąs3����M;:zq�S���mN��R�S����U#��c;�Aw��o£����#�լ�NϺ�w�� ��Q�5Tf�}Qϗ��b��gШﾛ���.V����F^�N�F�'^����C�q��p�y��j{ �Gw��b�^�}nT��CGzn�����'ä�k�Vu����:.�i�:2�ZGk=E^/r+|O������G,��I|v�u�~��zU���Uo堧2x ��Ԏ�iݚQ���:��gL�G��K�v$�5ٞ�#�g�0�C�~�^4���E�����x�������]>[l]�=�d?N3�;���}�r/��5�{&x�����y�Ke�(n��Ŀm����*0�/�Q�i��j}�z�M��;��㑿��\M���{R;�!/�s˝�Փ�t��.�`�DUpu5��dι��r��{�cs�~�zϊ�C;Ɵ���k��q��:���4�ҏ��;%��ڰv7�T[��O�,�ih賤t2[:1�י䢧�.v=A�Ȼ�����irϧ�\nr�Y�L�I�T�U0'��@��Jnr6��S���uN�W���_�f�,�6�!�6=Gh8��ݯ^wΦd�F[n�00��fn#������N��D��Z4zs�%ԥ%K�ʑç�$2N�G^Pi(�GL�g��dL,�z^ɨ�l�Gf��/jn�o;L;[�D��@X��,A��3O;arW�	\��c��-���y�z7�|�b��G_�)��7����o�Po�p)�D�a^/}s�&���O��梖�]uz&��9��g�ґ������}dh�����eIe�74N���W���H l�ĩu]wz�Ϯ}���+=�F�%qW�ZG>~��g=�tT}�t�}E����H%w�O�x%U�i����G��ɑ�.y��i��e����yZ�I�ZO�'K����3n���U�yf�F)��(���`�<`�{jȦ{��}+N���m��Y�W��Ӵ�3�;F�;3��s�S�yq�����;&�EG�މ���^&&"���q�}Ǳcn;�xj{>�{�R͎�J&]���.���x��T�-{Ƙ73�v��\en�W������Lm��`W�K�N����V+��d��΀��5C��s�����I�2�h4���C����>�������P�#胲�3{P�[������gܩ�G!��⚓g~�D�r�|���_��Y^�)7,��wQ�m~}��icׅ�xL
]�^���ޚ�Q({��g\M�mΕU��W��+�v���XEu	K%�8S�2��YuiZ!�e�4�<i�W�rˤ����OWJȱ*wP�+ʖ1�_�7%��X��z���M�N�/�v+�W{AZ�O:�X�\¬�I][��wR}���6��;���]8�
�Qp�qY�H�h�W�4{�̫;�a;rt
�r ���sMD��&�����g�7��J�q;He�֗y,V��\���Nu0;#��q�h�_�^�qp����(S����o U����xǰ��I���2�kK3�7�v���Φ�
obRm��Ͻ���ds���?�{tu���dw����)��D��j�}��'Y�g�:������)f�;}�S��s٦��_������\�������	Ce_�|�#�D��'��z��n��R�ʯ�p����ɘL�{�p�:��qL�w��B����¶����"�����>����ޮͅ3�ƣ�k�@����M���q��l�)>/�����~������n��z�0��Y��{�|����$_������Ǚ��a<U�$c�ARg"=�F�ƒ��#<1����Y���ޯ
�:�K���7ג�Q;Ƣ�.w��a/�xiS�����X����=�Mϟ�q�Q��j�/����������	h��|�1����7uMw�W�a�N*k��Ӵ�Y�_ ��ndHy>�@�%�;�\�/���*�w�/ʹ������ã�K����bK�(�x���W��U�̺���ۨ�*�_�}�ky1`����즓��F5]T��7о�4\sI��q �Wm�w[ɚ�^�vG(�����:�:�s����)��ӯsT�[jK���������<����S^>.@��Z V��<�J&�|;A��m��'�S^���v�*s��x��R�Q���QH�<������sf���rUh�2J����{y��K�8�}UJ��/��͜�:��l��f�]/�;��tR��spN���ǋ|�+�m����Ӈ߽#��Cg:'k���p��	Ì�\^��+�G����3���PBN��s;iwb��a�_eX���ls�=���lN�<��qb�͚Ӭ���ζmd�}��ӚF.�����i���>�W��約��5�״�q�>ë"����w�z�˶+&�z�>��:W(&{}R�~�q�sǻ~����^�C�}��H\F=�g�&pa鿢��wr��=�fh	�~纕�F�<���/Ϊ3~k��9�~/��q�O�;����V�"_'�?y���6�����^�@�U0&/���L�>�ԯ�Rw���N��>�~/�E�}��b���f4t<�f�s��<��Ɣr���G:"�n%Ho��O"*�F�o޴=���po��<=^��,��\y�[I�1��Z���&�
� ��t�=����&Mǫ[߶,�<�m	��	�* �,eNTΚ,]]!*�m_������{S w�X��JE�O������.���h��،U�P�.����+��:.���6��[�8�pY�nnq5�8�Hg�O��v�,�c�N��Rۊ�%��߰�9��a>�Z2֬����_f,���N�ǎ�>=�����C��ǳ�CsPO@n�Q�+԰���*`�7�N�ǽ��]��Mz{8P�W�#�?u ^G���Q�t��C@�9ۙ�Qjh%S="��Q����'�۸��}x|N��=�qW��I�=����������:"�K��U<�;}_֧7eNn�/�³��E9Zwl2��7�Q����s�L�>��/ho�`/H�ǀ����f�?L���>�MG/::A�GMK�tG��27�s�<���ظ�>ۘ�Kޱ*N�����U�<��w�[�������	��}g�K�&�����2|:M}�t]Ly9�|�A.������Զ��� ��<��{ڐEGz�$>8rayFV�q�^�}��f߷�s'���{r�ɾ�Y�g��j�g���T�������繂�B�8+�Iӗ-���j��T=Ş۫5�)�U�]�X=H��v}�~ Tb�`_����uz�#Q�δ=�ʱ��ӷI~�UV���O�p��s�K&��w�~\D��Np��Ù�Lx_�w�5QV�}W�I��W���t�f�̀�"���Lu�qݷ��Vݻ�.���+r��8�=����*��yެJ7���]�Sxw�/4(���A�2H��w�f];K>b�oL��:��b�t�5�_Ϧ�i\[jYj
И0�h�R偃���]��9u�[��Y��Í]-,�NLDT�$���Mg9W�G|�\�9 �b�-(rڕ�Gf�ɤmr��F��*8+6.�uF�}�#";��K�!{P��d��ƃ��Gq����T)�s͗:�NƗS�oZMӹ�KǸ�2gê񇸬gk��'n!i*d˾����k��嶶��"�R���N�u���]L\�Eӑ�k�9g��hM.�=����U|ݺޭG�㮺)=}���_3�,�Fup���O!�j��2��y�����:%փ���ed�$���Jy�v,�CR�=L&��NHSD�]l��^��c�E5��cx���5m`9̋���!��sxF��B7e���hcArŏ�,٢��)��S�sv�SXޑN���
��6�U.��v���l�HU�"��̫������(�������W.�����2Χ��ӹ�ݝ7�n��؂I��P�]w[6e���b�D�E'ϭ_/�sd��T���າ���w'V�4u�zΕb
�e��/#V�p)u�N�لN��v�&RLϐ'�-}��n�U��eL�=[[d� ��*�H��o��ҳ�;)cr qEsUb����T��3@k$62�Zr4���i��Ft�]}��V""����+�@�Z�e�3%b�B$�Q��SƜNS�H��]�1ڶ�p:�$X�a�3��1&j�ܼ٬VyA��-��޼Ac�Wӭ �W�J�k�5
iU���ʸ!�7@�J3Bk��cU�ڰw9h��ue'f\��w;��D�R�Av(ҹԯg`�A�ܹ��x��b�!YPs���W���\��"�7�o&>�<;�_Ep��.���%Ew���NU��;���>����{�6�v��O@��.<n�M��*ڂ՜��,�Q���h�%��K]nwLK�v^����D��l��l��29oZ4+]���U1�
�n'W|�5�ۼ��^[W�x泃f����k)d/�X��L11��w˛3�� �%)u�m�qY�������[�+J�{3��Y��&8�ܦx!��Ou��E;r���9+����eAv�<�J�Bjt7Z�F��9�!�&�������Ѥ�pT�w3ڔl$�|p�EE�Òs�[��;�{)ʷl´�����F�P��䫾[�]�3F�Vi�J�L*�;ܝ>�J��7R�fد�J�ة;s> 
�"�B�-�(�E�b*(("���V��*���jE�lR�*
(��*����0X�,U����*��*�*��QQYUE�T[j�%QR*��PYR��*�Qq�L��"*�J0TEbPb*-����jQc�"�QU����"�Y��̵D\eQТ(1�V(5��YV�V$��,˒-�����R��U��E�A��b+XR��`�Q�XUb�am�E*LI1P�Q�,abYX"��ܭ(��J.%q*)Z ,Q�J�lF�$R
�h�ɉC,
���L�D4���-����X8f0��U
�\A�����%eX�f5k�-��wY��� mke<2��3rgS���L���c6��d�����{\ꥑ�*Q����ホ4Swib,d�C�/&�Y��^,Ԣ�pݗP�FKW7�����n/W���ޭe.��9���v��R9���?�4�=�כ=y��|E����>��d֗q�;��!9���X���_���S�\v����a���?Y7�M�����jY���d�rrp����x�y3��v�HW�����gC����1�>�ū|�W���,��7�k��*>1מH�I�T̰$� w�~��ͪ���j=�C���nˍ�)�U���	h�?W��r��u����@@,ߢj	�n�;�j�QT_?q��R+�a�ٍe�}qI�G��>�=�F���xw�mK/�|O ��E�o�&����q�nה`�ԁy����\U��֑�~��g��[��U�.@� \�A*v�>��4}`�O�F|T����x_�x��\GSY��o�F��������5Yj+�w}��y�ϳW�E�r@��>Gnba:��?S��ѐ}+N�#,m�߭���~�� �}Q��C�Y�N�t��kϦ}�����"^�OIh���>���11MV��|7P�3|	����[~=�0���6y�4��5�V΢7�~��Y��]�(1@1�|���LV�"��J�ug]p�4<6V�o�l,�� ��[f���qJऻ�*��\+�S���U	&�t9��1����,�ٓ_c���2�M9�3��[gTI3I��-��wҷ�Db��h����f��
uz�C�]Z9�v<�d��r���@�L�����[��z�NE/B4��0;/t_ez���kJ�u1��ޱ^Ψ��9ܡ�P�8h��D�9L��fl/M�u�h�ř~��շz�sᾅ��W����^�?��/���"����o�ّ�;��Q��a�w�Y��ʫ�V<]�ǸVD�X��Z��ٛ��^����q�Nw�q��g\N�ƽbw�XU�k)%�5zQ�zA/���%,~-<=-~���^���灼�c<�=�8�Wo;2z��ό�^�<h�b>�o�&�V��OMw=gES�t�d�k�5�R12�o�_x)�3ܹw�o���F��}s���_��F����Na=qUƱ]1y3��;���n��W'����O��7n�����9�u�{o��%塶r���ɗ=����j9�M�W�{��:+ߒc��Fu����B�����|�ju���J�,��ec�N��!7�I׷��m�Hs#@��հp�Z�&�E�*�GzR>�I�\}��_O����陙~�^.,v��u�/���(
������Н�n�D����8����t��v��a��m����vڷK2;�5逰��o]�nԴ�\Z��A�����*��#�*�0C��8�o��=׋kCR�� ���.0G�.��ռ�s׽JËs~x���x�vNO7xo~P��@�GP�H��q,��s�XN;U����l��zx��7���l�~�GK�gm6�}���G'�@|D��.	^+D+�3�_<V�{�>�Q�(��r]�>�83rQS�����Ȑ�\�/��baz��14���>%��*��_�����>���gfk�/�Co��>uro�X*���{.���7-�����c%��y9J���ջW콗t}i�=����W~U~9����.� ���*z�L�v�7'�������˦���iG�c=�tB�U�j#K��7	K�	��i{+��	���~��&ξ�k����Lwz���mG�6�g�A_ٵ���;�5��fW=�	�dyzd���:f���v����vi�Su�c����N��2���s�v�?\d�a�8v���m0'����W���*'w4U�ny��Wg�>���n=�{����wMĖΝ�w���,f�ñ��p���휘�7��,��Fށ�ͫ���i=�:����z��S��!����>U�^Ac���/V!��
�;MeҤ&�"��H�X��PЫ�˱�+����	+l�M9���/�xy�c�e���33�L6�W<���/��ؼǟkj�kzr��q_�@C���ޢ��ʧ��g����������|@�g���z�M_�<}��_q+ۈp�>V�F�6�g��X�B=T�{v3���_����}!4��o�燫#���k��;��V������Z;��T���(������Ӿ�Ox��������}�q2��l�⾞ua��ǝ�����5�^��]!�y���v��m�]�z�f���l�*yQs�#q�(;~��쀧���^y�V��ow}{8��y��s�7����,���N��Rۊ�����&�
�{�L/Ur3�YN���$;�yO�P�o��c��[��k���ǆA[�y�!��zwT���XR�R}~�s��w�.By^�=��T'_{-#B�z�/�(�4{�e��o��x󞸉�'VqW��o_#�hzǎ:xp�Gw"ǼjJ�__�sӕ����b {6�ECʧDX�l��-��G�m+��՝��
�郁�[�'�=�px��T������3�>����G�pS2����+=fV��r�JvN�|f<���t�\g��W�+L��5���|���Ш��:���~���`+H���+�Yp�%���*�Fi�U����^�g[�rF�1�0���=;�[I��J���u�q�� �0K�j�vԴ��n�����SC''GpƂ;��f�neÎ.�7B�E;�=2�k8����Z+Ԭ�X�V��%��w����:�%�.�U9�êݰY����y�1Ǆ��2��J�y+��"��������̓���+IG{麆�+t����5�A��u���򺋇��[��V�x᠔��Ϩ����k�^ڱ�2d�ށ+�|v�j�2�L;�6��s�=��2&h���^Y�so����`:�xw��E�o���/���|�D�g�3�=� <�����&�����y���b��q��zo:��3V<%���>��ӝ��}���p��<{8�����SX�4������#�~�h��jY�f��7�mO�v�W�Q��g�a�㑿��\KG�5S�N���{�U]۫�Ɣb>��{R����Q�Z^����t%�x�͆�~�}oţ%%���'!�^Y�����R>�z�=�ʊ5n\�ɳ`��S�x��3���3�UAvw�s0W�W�d���Wp5���xz5:�=���7/���\��Ϸ©��h����� T_�2�>����x�o���_��{�{ެ�Z;o�l,���F�z�p�=#�5�	_�P�j�Yb6��Y����w��M���Q�j!����-���O���Q*!��~�[R��79�`lL<����	�~Gz@ＴǨU�8���E+��"�Qu����WL`oC���p��|��݋|/�Ju�*���!b�q�0P�ݫ�寤0��^�>6�Ũ��u��yi���HU�̧���"��v��^ܕf��jbɇ;���R�<����5���G��7>G۳}���6t�u��{/�`v^��@&u��n��t'Rn 	,?)��>G3�XZs#e������__�s�L�����#�	~���1O0�x׳�r+��Q��\LL/T]"f"������R����\�<6�R$�Yw��=�͘�Ϻ��v'��;�+��Ϩ�w���S�+���U�o\�wQ
���<��Vy��=��y��Y:.#���r=.��K8�*����?�1�^�kb��.���`{�M���t]I�quy�!���R�QF�{��s��វ�"�Y'�\L��v.O9�%G�Q�=�U�i������j;6}������ۇ�p�e�g��E������c;S�מm�/�	^�j�.��ㅒ����C.1ևy;[7��t���r�Ƿ�q�'>�HdjBpFG�q���k[��>�mΔ�'��O�;,^�MiW�O�i�r7�^����_�qYZᇝ³�'������s�\X>��x�=W�ʞ1��k���8�����kK�;�q�@��77�w�����4[��'ʅnw'���p�Ygm��4S�v�,�ct��ǼO�p��ܷ�L_HB�2�*���ɔ��=
ɳk�'a��Hvw=�o�;��Q�:H3#��Zn�+��.YJ�ԙ��XWj�b��Vt��������,�hy��"�	\w�tu?;C��R�'�)��s	몇�_b�cՖ�k��}`G��ڲ65�V=V}3��>��ׯ�r7μ�m����CFC�Ak,���Jw�ur��G
ʽ�9�� z.�p��3�^F�B�y���ν�=ҙka�B��L�,��7�o����.j�������Z�>����z��]�����q�������q���X���O㷐�\����z��'���#H�誑%J�|X�9��<W®��a�(�uFzͺޭ�ƺk|��y���:^S�}�^����46�Qx�;��̍�k�L*��3c�e+��Q�[&��/ѵM�=⋛�ye�H�{)���Z=*�Σ�i?k���V�|&/�bPM�H�W/t����6P�R���N�{ՠ5�ȑQ+�hZ;�2�Ѿ��C��n�^]U���u��}S=�L{
��\=ί�=>�'mR *�{,
y���sUR��v�/.{f�����¿�h��u�t{O���K�	�؆�se����V�/o��FER�$xq5v*^IL�6Uh�m.R��2��2�8��'3��a-�Wn뷴�e�ܤz-j��S=fm�!﬊�N.׻:�嬻۲�5j�Z��:��b����^I\c��_hdЏ.��K�(H5$����f_R(]u�U��(�Y�*Onaq���y����ݖ4̨�Ǔ����7w>�ʏX�t7C�ksȌ�>>�}wmQ�_�He�ȓ�v�v�?a�>��p����׶��=�ᑔeǣ�3Ƿ���:�Іt���G}sB_��w���Hh�ɇ}��,f�Ý��]_��II$6�i���v��@�r�7ݰ�%m�����=�n$�
S0��s���U���t���`F{�T��o����������7���Ol{��Z��3�Ɛ�ǵ,���k�Z�M����ֺ�
*}GC�UC�ɝsx}3q<��X^�iw����b�{����P�1g/a�;��Ss��P��o��^��튦�����)φmJ�<�ᮽ����Z�Y6Y��Ë%¡;�zf���zQ��=q�ˮ|Vo��f�HfXSȊ������A����N�e�������܏z�C���[G��K��XU�L����R)�=�2�D�a^/s�D��Uow�+���Сq��ly��u��?_�=g"%x�8��vs*LlDe�{�fok�A�C?l`����z�4J�#>7w����T�[K���Σև������9���J�E
�7,3{ʻw=��6�zZ�=,�u�Jo����m���9�T��q<�z�ɂvI��	�*8�_J)wJi�E�>��)[�|#��X�����{�/'����/3��w����ґO�H����/�~�z|j�<�ź��D��e��k�37<�x'ٳB��Xp��ơ.��_���㞜�dG�| w�ˑ�y��� c��y7Kz��/m����7V��g���/�t�)���~>���L�N��Oz��z�.�j�ve:(��a��t�\g��U��"�\�b2��v.4�'�*F�{���,9��na�S�z�`z�ʒk�����>��z�����+t�>'�f��w��3�UA���+!^b�f�C˽r�3�A٨^uc��Ԃ+�V�,ev�/^V�Ɯc���^��+ں+z3=cԏ�\�f��� �J��/L�B�PK�v$_��֋��Iㄴs]���U۹W��/*�vju�ͪ�i��M�[ V+v~�g��~���Ω��5��G�}�c"�˸3�}���z�*�M��\;߯�>��ms�MZ�gS��.�V^�_VXF�ox��D�5�Ϗ�L��ӓ����ɭ.�ɝ��ƹ	��Mֽ~���-9�=1�{�J�r�Kw��cm�"<��hd{(v2��5��S�6�\s�Ut_fA��]���m[�2�8��(�t-�HW��
/�_2�9���䱬���]թ��%������[{��W7{���p���gT*v1�w��+�N�U>GR7��Ǵ�)��p��ǘ���޼����#q�vKg"''����1s�,\dγq�<��wѧ�u�[^��Y�NO)9~�^���<2#�|��������r=��,�6������ WWW�krg�Ѭ����.y��a�uT?�qaA��ў�-�~�����)��9�O���v
Ж���W�f���/1���x�}}��ͨh������x�gkûb�~����;&Q��GT{�7;s�7��of�x��|N��7NhTz�7�����Pѯ�%qV�֑��(�s�'E�Az�m��/n�p�u.��^�/���|�0Xu�UB��#�Nf��x��\���jo�.j9�8%�l�K߽�JG����t�iY���2聐��x���OE9�Ҵ���ڝ��ڄ�W��ǒV(�G{j�����?L����
߲�^�O#�:Z�n[�M*~��~ˮ	�GЫ}��1{��yM��ά���׋s���y���[�	>�n���Ďv=�Z3v����L�J<Y��t�֟ium_�N�xZ�Qfߝ�C���np轩��@�}F��v�_�-S�����4`����)c媺�f�Iv���dy���'%g-�n�Ǎ])b�tL�m&M`<�����X��9w�n��5���YxOi���u���ܟ�\��э�+,��nl(�c��E�C�5��,HD�#/k�w��4n��AC�p�R#��E�@BąnQED��*��u�Y��ѭķD�v� ��<g/N���*Z�6�Y��?vF��G{.�}�:������K�}�̰�u᫴�\���1�KFP{8�Ύ�b��������K�Y^�Mw �Z�����6us�x�6!�lM���>�D�;&W\5���V2�ث�5;�k2j�M��CXg����XGU�� iN�
]pa��n���y�wX�.���<�|lM��Hs����ɼʏ7��(�J�E�e24���`����q�8�Å쩶�F�F�6챜�u�,�����
R�4��]�M[�u��ӣ��V۠]�sq05ehW�G��)�$����Ao�,,��L����Q�}��N�ư�&-�ռ:����gZxLd;��Pr��h����x��m���XWX/�gA9&/2���A[H���qrb�)��]h�w��]JBxv��;3��#���7�&�;R>;>Gk)��6����/��b��c`[�^M�v8�&��i�,�ow�����F��S�;���T�{,U��n�� u�������>/�����^V�>�(񰲔ՍbHb����N5�y1A����T1;ں�u�5��N�\�����J��^$�2'���A�����ʔ����E�4��0������8G�le;�����ٷn�f�Q�= y%>��4(�,��^��K���=���V�:�\����Vp쇓�p�����>WX�q�][Dk�[ìEAU���켮��:�t���Ww\|\�y9��t�ִk�pRS�},Q7���x�ӭD󡈲���'�N�� TzԻ�m�wX"�i�s9�),ƪuk-ٖ{&��N���*l�e%�B������f��w+X�A4���eE��v����Y�\սl��v6�|��l���'3�0��$�/�6��۝9-���L��&6���lknS���"���b;ȅQiuǖ��_+˲hPc�(�� E�C9Z�8�/�o�������|ێ�i�yr��U�����8���G��mr�{ʷz��jU��"{�ǣ/�����2���aK+�U�H�>/�Ŏu�v�dM����*�EB�y�*�q�lg"��0㼔9�{��y���TT��ؑ	^^�v���cM:뿭/�X��43�领VGk�1���n]q�7�@��^e'�н
�V,<(̨��Vm���0Q�E�kз��*�5p�!(N5��j�%V��F0�α(n�^_R�W\��T�jfn�`�6���iD�[(e�ԋټV�,��:�b4%6�Z�,e;�K��\��u�JY�8^.2����*�ؙ;8��AA@L�ݜ�\��qc �_��?~�<����P�XQf8��$PZ�c��RڱT���2ܶ
��2�[�����D\faQD1����)Z�!��b�1�T�PLlֶ*1Lu��6��9
$V�aki�DUej�`��5��`�QaVҶ��)mm����8"U�Lk�*[Am*�Q@m��KV�r`��Ն$�\AA@��"�aU�
��aTt�iX���3)�L�Ȣ�m�X[q���V��
*�Tbљ�aR�*TYR�R�)l�jX�e��DĨcX�j*���R�X�UR9q1��Lt��k0��*Lq1�S3[J�ڕ+P����U��U��1J�eJ��Ԭ�X�Y�T�S+f&& �-�����f&"%��.Z)V�"J��*c�� �>,���VQ���Τ�a�6̜�V��L�rܫ��5];Dk�1m ����:˗�Z�Gj�j,��7j�E���وj\r�p������s�[�
�6����f�����׻��T���e�f���ّ\/����0��E�Ι��|�`�[�:r�Pzn"v|3��ۜ���,{�o:X�����<M_�o�F��՗�G|#3�벼�_��~[s�פX"��dX�.U���ֿ�}�C?)z�G��Ω&�T^����v���bW�(���Q�J�u�n����=����)dU1�5���&w�=[��&'9��%���7^߽�CqO�!cT��u���m��\��E6rNa=uP�o���>ꧦ�a�w����ky>��e�y�^�&7�����ϑ���!{�Lh��W��ҙQ]3y6�A��y������5	�+���Zڨ^7Ϯu�>�\�/���ļV��͜��ۧI{Y���ݞ��#���+�Pf�&)��7)�q�A�m?<�ϗ��q�>+�ޏ<���w{Wzx��ǯ(g�f�y�dq��H��q>,y�_l���:��A�7}*�m��M+�7/pǷ����:k�n��mz�`�D�U*5��"��|��W�$���4�f�Y�\��hLq�(�u�!�Oqe�ݸ)s��v�_���]]�g��8�8����A�����Z�Np���w��ޖ�T�eϳ9��o�hr�)�{z&���uE`Gs@h"�wל��(Y[ �Ep"�'�湃�Ӛ�=;��7|+�R�c�x��z@󿽹�030�Ah��L/U�&�r�+�����쾗�}�;��x�����z�_�zv�+#޾�{s"E<�M�r&Z=�z�����]��[�(�#����hޖ�v#P��~���_�zy�Zg@
���{y�Q�eo���ܒ��Q���}�΅�f�y�C��u�j3e�����;�\�~r�����L#��+]��v��a��Ԓ����|�n|�և�>Ѳƙ��],z�<̏},o�3j.zg�U��ڔ����:}���d{~;��~��Ӓ|��Nׇ댝��:'���[B���{r��.�Q��N{ ��p��8����k}�bo�۝1ހ{G�Z;s�/+�X�w��:���[Y��g�zQ��]�_���Ul����u�ו�Cצ�\/h� ��.����~GR&���οTÒ���]f��R�᫡������9�9�ݾ���|�i�.�ӊ{f�qW��%^kg'Ӈ	�eϨ���w�g}7��'�Tf�^�q��K�}�~��'j�7g�y�E��z��m�-����j�j���Q��Y��i̤ȥ�6O5�c	3���֢`+���L��]Y0�.]Ct,V�|���\m'�>�n
����;�Z`�*�諎��[���hV���ssR��}TY���u�]o�U�^)`�v7�_�w	���%��k�)����`M���L�>�+����~��w�M���5�Qy��n���ah���n"R����nY{�"YR���Sb��x${*Pg�cA�^����Ӎx�'�/��3�>�K��������,��k�vo��U#ĶQ%׼1x͉6�V�M�]�D�z�ա��Zd{Θ������/��0�5�Z 8�n�����۽C�f�z6f��Q���>�'�y�P�|��4.z�9�?u ^}�8T{-�����7~���~sw7�~�vw#��Q b>��M
�����g	��M6�/>���|���`xo�UL�1&ߕK��z������RE}�Ǵ�LW֨�g���T)���
��~W~6��0�{��39��p.��UE��W�='ӻ@z�����W�Iș��_�t�_��#�+L��{^����A389�U�~Q���=�{��d�G�������Cī$==麆��ͽ�'ä�$y>�����9�<�7]>��AߝY>t]ſ:��{jǱ��w�g~�����B�p)����z��{�ڥ��I���Z*]'o�+�ˮ�.�c��
۳��8v�<� AٮV;h�	Ф��o��@l٧D�s��$|mI����|�� �y�a�li��ר@���Q�y�ۚ��\J�5��O'g4-��z�v���,)��ftl��Q�?s��r�r| I_��#�Q�ޠ7���P\��q'NM�
i�L\n��w���0���]P�3j�ޟx�������߫YEz�q_o��A��_�g3��݋�Ux�qƣ���mO��xv'e�����\d�\ޖ�o�J�����_�|�l�`�ao�����{���&�+�啼}��<t\��=uHz�kK�ɝ����'7=걹1�4|y<��>mbь,��ҳw��{O����w�w���;%�l�=�L	���b�ɝf��/�z�_����\�G�+ӝv=�z�<<ϸ�zS%_Te�E��beD��⩀��~��>ٌ�=�s��rudmT'g��c ����p��d?W�\��G��~����RV}V z�zޗ�[�٘p=I�'e��j4��q���Ȉ^B���ᢾ~�_��l�LX�258�*�wf����鳞�CsPO�M�zhW�[���F�4k�\U��֑�~��e�>��"�~��7�y�[�]�U�/� 0ڙ\����}/ơ�W��~"=f�T�#��s�FּQ�)��	��r��iخ�����ܞ�C\� ��o�;����u�r�N�2���(�0;����Y,�����]��z���<��W��W#k,�TrΓ-o����w��G;���-��oV�N�i�\��+�yX�t��vƋu��,�ɏ����UKޢ����P����\����')�x�ȃ�Zw����TO���;���egV���ѽꐮ==^���9^������L7��(�9�7P��LOur~��t����6ie����(n�(g��'B~��^�C�9.t\x��"�{Ɛ$��nv:����{����z{�OLu⮓Q���5^:���Lϊ�9޸sT<-N#μ%=��Ƚ�W}6z����l�L��~n~7��I��A����W���/L�FzP:M�p���t]�Ѿ���{�j�Bѓ6}D�r�|���c<l=���q��t���,
�5g�=���[��I�����'��J$���|��5��7��Vs� Nᔿ.?�����g���6���9�{����9�{���x�g�����\��ư��9��l�V�jϪ���&��GGj^Ptn���{պ���]�G���Hʋ�l�b�m��낸~�C�ʊ1_<b�9'0��\��T���>�w�건����;��\dγq�('�z���k��9�u�{o��^Z��\���&�����(�f��vb��y��s�����
�H���]@��#U����:��h{�μ��u�17���I)fn(�l�#�`k����mS���*�������r� �l-�h�fae]�p�s����}V�%�
U���K���>�3�loM�C��;2�mT/��ȣν�x�_e���=魄�6�4{���Y��[W���%ў)����n����w�A�pߕǳ��ٗ�����z�eo_g��t�}ޟq���� �e��L�ٲ���T�*W~�<��F�7t:���>}�)��`�Dc�g�cT��ǈ�1�f{#�6\�� 0ۊW@���>����������^{8���V�\��1�i9���s"E})��τ�\���/�ONP�O&��2��Q�Lz3:�N��gT��zR>
=J��=+���Ƹ~WK�����F=Ƽ���8�����gʎ�&@�j-	�};G~���&O¸[���K�=�]ht�;1��*��U���j�^�ZU<M�χm�fǇf���[&��>�-T�ϝ	���sf�dw�1��g���^����к��-���n�s��r=s�g�w�k헤ɨ],{7������a���;��Dl^S��2\ǣ[�<m�n���N�ߤ2��3�g��f֏\FN����\�т�:}jy_#�r�gױ,�seh�S9W�s(�%���DR�4m,�F���l��ؗ��u=k^��(���O`���B>��x�= $�V��qk��gE!�c�nΖ!��g�u��Yܙ4�y������ٕ��r��d�+��AK5���V���G�,g���_�{c�b=8���w�4'��L\Gz���-�ڇ�˯.����M����c�ODb�Ӿ c���� ?�����w�=yo�b�ߘ��g��x����oJ<�����+791��]g|@��]���.1z��.�hU�hp��:��J{z%��Ue���4���G=�g�g��(<UP�2g}7��'�Tc^�i�S+{	��0a�`]�K�N-x�G��T��ɒɡ����z��d�sᑵ+��yՇ2���~��ꖇtH�yq�j���w�)��i\��}DS7��L	��DT\�H����M�]]��r�t/iW��෣��_���y�^E��qN͞��T�w�q�׏�{W���[�4O��/sk�W������BR=�{�����G��������l�}T�|^�����z�Mz"�h��g~�|��#�i��ͅ�M��ޔ�m���嫡}}��L0j���}��v;v���S��5�_� 6j�Ш���a�Z;�a��6������uB�B�F`D�c#���˫}7&���O6�IWA�1`.3���U�:��ݩ��[����|Z;�x3Jƨ��C4!�h�f�A�	,���Ӧ�]���gI���]��Den��Gy
�-���8�N����E���s��R�W0Zsw8��s�y�+���T���R��s�Z�3�=�s�_��ϔ��o�������|����5>�>;8�ɿ)W��˟Qd|uM�g��T\�2*#\�W��f|�қ�N���un!�\s�Lg�צ�.�)rr���{��{	��n����.��tu�ן�AK�gv��-�H�+�3ﺐ�'VO�N��|�r���j�\5D1S�^r�~��F�A�mu5���?�綖��ͧ���5{l �z��J!����.9�}Q]�m䊥���~�g����v���ڭ7�����`�U�ߧg#�삏V�t,:�����K7�*���o_��x���b7;,e�m¿�Ԭ�i`o�ڟ@����)0�H.3Ӈ.���	)�j{ˋ�U��B{ư����q�A��n��՚ǐ�T�\��)׷�����s��3��h~����s}O�q�8�D7�y[%��l���=2�Ϯ{ŏb���8I>˾����جz��&X�����-�μ�l_���K�q���>0�|*�"�S��K���q_�~\���a�7Ws���1�� #wìu+�Y���;]�`spqK+"�%�#s�/*uq�+gB��um���6��������	X����� Z�^�%>,v�W�eq)����b������։H��H/��̗w�i�M�Y���Oz^~�ژ^�=O�y��dy#M��>�] �>��A�៽'���d�@�-���|ω�3��p&��D��W�܍�h�<�\{�6r#�'�v{��/��k�̺�U�C�ΎU�蝢����|N�����E�@�d�}��7�%Q��ZER��ND�����Y�?N�?9r�G����g�}%���ѯ�S#>.|�g����}��g5�:2'��3V��<z�J�jm�z"q�G#�9Ģ�N��=�r*U: \(-���^�De9��>�5Q>R]��T��oyq^��(m�?g�ߦUzb�ҩ�g"}:~���y5�(�:ja���Y��z�F�{�2L�>�c�j���ǳ�e��N���~���r=�Y�=��EB�� n}X@)�6�z��ҷ΍�������]&�4�O����iد���ܳ�r���wVj�[��~��5�q'N\D������n�;�ͯq�����ۇ�m�_�/UBwT���>���e��Ƶ��^�Y���c&l��蒎జ,_}��r�n4���X���;�=�-n���g�YT�;�Ϧ;�ܻM��NF��Xd��\e��4"�oB�{]Q����x�s(VxnRQ2u�+�*�Iʙ�F�?R�Y��'J��!]����f��uI��G6�)>��M�3wj����#�[�\;CV���SG'kGV��B�j���:��F��Q/ʧ�� ��|P͉�c2gB�
�TM^o
�)��{�ʬ��{>�,�~�q��ǁ���=�Uѯnx���=}�VU1�dTf���&���e�o1�'��&[7��7�]�Φ��SG�-֎���q�mr1qtSgמ�3U�F�zL�o�of�wD�}U�Dg��/&u�ɟ��*�[�~㚥��D_���Yhh��g�K������V&����tk�rl%7P���\;��(+�u�����}�L�x�Th�=���+�\��!��z��,���)�@-��������L��A�;~Y7�cjU���Ӵ�F�}�}�;�zk�������ԣ�� 6B ,ک�+�����v�f��]�fg��+2�q�j�Eyw�
�?[f2<��ϸ�>�u
�W��p`�j�R��Ö0sR�o��#k�>z
���K瞵_<V�Z�kō�{i�N�c;�"b=t��`�Ƹ�;4򚊪=�n�wY��@.Ւ$'���n��9��ؿr�ƺm|���<���ߞ�" BO� !$��@BI�� �$����� ����?� !	'�� BO� !$�� BM��b BN�R BM� BO�@BI��R BO�@BI��9 !	'� �$��b��L���[@ \I� � ���fO� ď��<UTU QPE) R*�*R��T��B��(
�RD%J�*��(DP�HUR��"�*EHR$���I$RPS�!IZe*����H�����D��T$*TJ��
�ʊ �QUDR�AQA�
��h�Bٔ�"�����*T����$����*���E$(��UT	
�EQU**$�$��B�( J�(�%T����   3y�R�N���Jn�ٸku%u�j�\�Ҕ�g:X WWk���Ӯ��隸�n�ӌ`t"�u˳���m��ܩv�wrD����U^    b��(��:���Rj�Ւ�'4�y� ��q@z=h =@   \���Ez(�k���� �(�@   ý� z  ޔ�H�M(AQ	
\    ;s���u=��]����f����sVm���7+��rl��m����[�����@
[����]�u�2،)�c�lR��H@HJ����   g/keRf��ȭ��6(��P�H��,V�A]���:�ƕ�UԚ���Ç*�ݻ�v�nNM�M��wZ0ۻ[i�� B�UB* T	^   mު�M6���]�K�;]ڵ�*���#�S��s���F.N�]5�%�7I4im�չU�5i�nr�ݩU(u��R6em�a��ꛍ-'P��R�T�R�	
�� ]�U�ٺ��#mv�2X�NQkkK�n�uX��a�Zꪩ����]7n�:�\�iٶ��õm���3���M���n�E]ڹ;�U�"�PJT(��� �Q#V���u�4T��\q��X(�w\�B��t�:���M�gD��-���SU9�]�����u����B��ժ��E�K���l��J%TIJ�@kV���  �:�Ѷ�u��S��AU֫�l7aUM�n.:%K;���ݳ�7aM�a��ƭ�5��[NUt�f���i�m�wV�]���N��7T�Wl[vBBN�(UD�RB�  �x���5"K�鳪U�W-���)������n���u�'Gu�ݚΉ�Nڑ]ݵ˴��*+����UIڵ%�]��:�ʸ�픩Ԣ)�KZA��J��  #�{n�J���ʊ�N���s�sw%n�5ݶ͚�݉6��5\�vhs[u�����ۥi��wIKY$���kV�Ӌ:�uuە��� �~M&eRUA���hb)�IJT @���FH4z� )� ��z�  ����T��@ I�
zb�"���<R�Z⨜����{"�*���$ hB.E͛u�s�l�1�?�	!I�?�BH@�`�		�BH@�rB���$�$ ������������������f��Qq��a����V}Y>�V�SB����GY(��E�(��KE*  ����wWDe3��#�l
)���5SjE�����:��0�%��(�uP�
u�8�[1j�LMv���Z+Vޛ� 1��fe�PZb	41,�6�H��]*t�sfeփI����"��Ym�\{��%]� S�4���u����쁮��jͅk�s^(v=U"5���II��4�w�{�h�;��
cX��Zh$�#5n<�)j�ٷ9�ƾ$i�v��Q�v,ݐ�V��̔]&t����tMn7�,m�m*���������$��b�C�
�f#x豹E!���v�Uٛ���'@�n��tV=����d�4U�܊��5�n�;1;C�R�,�6�&�����~�z��bQ��v�=�nc5&7[i]���`ې�[��#�J/2�kF՗�f@dv�Ve*��U{+eЬ�����Q�i�Л�X�Ow,�ZkL��*�C��c1Z�Z2���1;�aLv6ΰ��h՗����m�Ԇ�Q<�r��+x�'.��5�-gu,ߣ�������4���z�]<%�	��D�eּ�j�b��`[��%Yb��Q�����۷�Q���QU�v!�4�]�c�MP`TkmV���˭f:gi]Lì�����XͳR�;�ee�ܬh�h���$�җ%�7D��Qe��iK��A^��ʕv���Ò���gZ��������2�Y���N��Y�Va���Sn�l:v��v���۰��yi钱;ע�7����hZ�5����X����;a����&�jlj8��V,d�Wl�%�PH�Z�� ]�Ő�;���&<v3\X�EM�X��0ܺv4�ۘ����f�ƫ3�z(�VD��.��#��$IRh^P@�!#��+E:�= �X��"���-�[��.�xi�}E��t��Vv�4�Y�Hr��Vcn�e��2���n˭eM����{Z�!uV��3����ɤ(�;�)%�˗y�XԠ�ct��v?�īǇ�B���Gq�@ڬߕ�� 6^R��%A��Т&� u ��cr�]$�3Z��R5`�&�OH�TywW��-Uj�KfV��N��Hktc�nۧL�K
��.�3m��k���@i6�3WC�'r�J*еHVZ�d��g2+�Q�Gy�0�$�!���H{�6 Mԙ�.�]��r��i��ÛeB�! ��O[I��Jk31�⹵&X)�� @ʭ�an�Ҋ�W����%tۺU��X5�7f����:�� J<h$q��
�[3Ej�4���|�*���[�BTp%�+W�Lcq�l�4-�Ǖ^�Y�@�X�1��wQ���.�c�2�#Q�7n1�d�57WMEP��k,	����u���N��8�U�Kw�B�ARa�x��k5E��1	YH[���ۘ���d�P���)���������0�S.�5MK��|�:�4�4�m�����+Ch��;"	K��X���E�Z)
Dµj���������d���)����ǚ�Q�Y���$�Z��c��`����)��q)+Eԩ[��Yte;d�tF�Ck4m�L�*R�٢�%"���fM��]2芊��t��x���Kn�j����5"-�ctJ�)%Ak,ּe͚ML�J+61Z���D�؃�X�TaaB���r��l�j4��hFE:֕dѵx^"#) ����ؖ���v)����^aŻ� ��%Eb��A���ɨު�z��Îm;>�0���JM�wY��Y&)(�f���p\:T�B�,�Ҝ��+SCU㽗�lT�2�2�:u���Ы.	ZE*�ְ�;IJԍU��͍�b�pV���¤ն>ncSoݛ(�b��(����Yn� �wkF�-��5��Aj�<5�u�PB�[�m�3k���(J�;n��+^St��/7511D��p�jIXGr΍�l��i
ej���2�c��h8�nD�Q�.����(��G��9�7����J�ZEKr��[�n@��9{�4�nm��)��	JX� X۴L$�Z�sjQ7N`��E�I�Cp�1bZ6��L�H���
w���IgX7��p�w��0}�����N١��E��V̡1$��"�����
Eb�eKBe�:V�6@��u銵���l�dwJò�­���H�u0&�͙b��e��6�YԪB@P�:��l��YJ���WV�F�]�!�ښ�TL�Za6��1�� mêԖ�K�Qݬc��(�
�zv�z+/e��EvӒ���]x�M�-�d)��LfmH�ܬ@?�	�lV��t�T]������a���6���R������#ݧSX�2�m�w���AY�ݳ
��]X����Ĝ�5tM7�D��sf'�é�We���LV�5t���ATn���6sm,�I5�ƌ�h�d�%E�2��p�(�)�f��R��0`ei�޽�
�3���I *�^c8�nm`MR��������-��x�t��ڎzP����Z3PW���&��O�Z�=I�I�T�۷�b�n<��X`mψ�8��q�Ku&��L�6I�$��n���RR8��xD�Q�J�ʂ�n��xdx��)��tܧ+��8g��n�T ��� $MCCNU�x�0kN�4����8��6��p�*�T���U�c��z���Q����ԡN�������8�hLu�j����ျ���tuK�s��Unÿb0˒�)����udk��v�I��:�Y�1cR��6��v�f�b`���P:T(��L�
laNm��˼fv��:�՛rF�!A�Kt;ː�L�"��s\tp7���f;�J�on)�b�e*�㈀�"������8�U�{`�������ţnK�j�%�-���P�bk)f�y�&�����K����j팸/f%���P��V��Y���4�"�T�G����J���r�dmhڀɳ�li��XΑ��.()4j�o]ʱV��ቦ����Z�8�H�+�{L�)kk'�T[�������bw�bPhZ�8�n�\��mD&B�vƨL!3�ܨ��g���j7�����ѭc#�6+s1S�0`�f�9nh���%`Q�=(VPy�i�fU�ӴԀ̦C|��@�V,�ks1ֹ�r��KVbH�˼��Ze��B���� $�7I�36
�vn-��D�#�Ո)cu�[)F�X�V`j���2��xH!�mLD��ڕo
ݼ;��N����eɚ�ݸ�ʋ5��e^�����	�e�@6V��z��˭@�mT��m�klb��֭P�a�����2`��W����Gr��ZӋX�a{dlC^�3b&�i����Sj�W���9R�`4�V�),6�%\4�+���+9��-1yG�+;Ohk��D������/.�:F��/)��u�t��h�%]d
Ã�vleӃ-�N��HQ����v�kSe�KtV�wBTD9d7V&Zݗ6l��@��+J��SHLUemmm�o=�@�����,lc!�j�̲.L[6ޖ�Mӿ�Ŋ�я�6"[�xuzJNT�;G�βp]jv�] ]��t
�V�1/ZdYjh��}3ˡd�j��-c�R]!.�3&�6��n�j�������p�;�A�w ch؁�V^)L�Pķfe^�3oB	�(e�5��%:�
[u�]*fӨ��D\'s��;�0/�.:��A��j��o5���9b����bh+v.᭷E,�ū7X� ���yV$��b����n�77TW'�
t���)�"Ŷ�,�q�������Y����A�-Eϰ0Ehsm�e
�7iL�M�&�Km�&�v�h�W�p�K�ME�)�d+-Q���0��^H�hi�r�%�	B��eI�asi5 rj�]�ٱ*�mL�� �f*Qĕ�P�ml���W{�fj6��Uy\j7\�9�|.nTtDWjР^��Xq`�Q�$�����c�)�v��Ei�`Ѭt�hiy�o#6�֑X����+���V�U&T���Dv�̹�Q���m���eM��X���*�*�3�ē�L$e=ښ Tq��&��Ye���O ڏܡzi��^TnlX�ܤk�![:�m\n��-EF
�a��!�-p1�o[�p�F1��
xd�ýtg�P�g��v2iܥ�ӛ�աٗ�����U�Z�H2!v�a��Z��Qxf��n�sn¼��Ѫn݄�D�8���!�d�U�֐	���M9�p�-2E�7���S's���9��.��7�`�w*�;wnQɭZ���G, ���֢�Rw�v�ih�4����Ӷ��CPȮ+�X�cQ��U�/oU��ޖE9n��y*�ĉ�5H�%%�V�8nT8�����T�nVf{)�N���[�:��L��nK��b�%�%�i-oj΁`3��a;%�����olm�YK)�c�����u��bN�b��cH��f��%a:�f��%og�7����B�L�q�i�'�
�뼢�i#��Q*H�Պ����f�l��C �`���^+UL�^Fp#C!�(]b&��س+nn�F]�ǃ�5ˌ���X�n��ú�����5��ɱ8�R��r�c�!}/DY�Ly��u� F�M���;���cɯ%�Ww�%n�KoT��9��A�ڒ<eIP�w[��G,��V8����t��H%VѼ�ȥ��"�[L�v�d*�#Tm�5
)���*�6!�n˲vN��Hm�-KS.�CR�,j��
r�%�i��dhmh�����ek��:�B�a2��*�D��^�ť;7�N�����|YJ˃Y��&mеo]E���l��W�=��N�F�3n���Cq1�*ӑ_��1�KfZ�3
���v4n�E�Y*:��.��:m�J�iELo0�KX�s`ڣ���bT�Mڂ"HA�#ѵtN�72Gx�%��M,d�i*�Mj�ki��Yr��^&��y�(��k(�?
�\�P�v�mU�KB;�A0U�%<+P�NRGR[�d��]fǯ�#�4��ʌ%�S�˦Fɖ��ޓ���r�"OM��hR�%��VR5&Gk0Q�)��u��jc��!%,��d!�T�olT6��\��K��+5t�]�f�ʅP���ƢR���5�t���mkw{�L%
����Q*��}�Vjv�ع�3A�v]5$2:�l�Wl�Kq,f�؀�����ɐ���E[(;�j��ĉH5�bJ�N�i�Vj�B��P ��T�^SxqM4��EҌWB!�-�/(m�nmb�&R�����]%�Yw*@w1%����%Rf�SЙ,X�c�h��nŚ��t��Ś�Ze,eA�W)�Ohԥ�+3����n+R
e�09h�����t�[��i��Ws����BF�G���/.��*J�aL�:�k]�A��LA6Mw[��˫��J'I��K�������1\��7hb+��a���lA2�غ@�+,Ս����6�=����V�J�-F�"M�Q�B�E��Zv�ґ�e�Ѡ�[s)܎�L.��d��
�ot��͐�
�����&�M/[Q�!MѲw]�*��@
QU�rIe�SN�k�W�m�0E� j*�k)�kk [�7��E3����z�5a�fR�hP6L!U�CH[�����{pn%2� ��f#�n�͚*ļmj�d�cJ���A��Ђ��o�f�X�a�M�������uK-�ƌ:54�����su_�1�4@�^j��{[l�G��`��(Vm�*Ե���-a�@�]=n����R�o4ʎ2w"���b`-�su� f�,\ђ�{�3Y҃�Q���Zs+5]�9yz����X��FQPn�j@����cd
x��
��e�l�'K�7艅�XE���R��A��Օ���W� {Z�Q�w%n���q&��^U�V�);�����6��Q�Y�`�c�Kn���,��"�@Ґh�&-��[�[��"�Yx3q��)X�8�T�L�b%�o.�o�;�%�דv\ܩ�uv��؍\�PK9m�v�V��+��V�T	��$�J,ѭ5*���3����$Ĕ7G4[��H�v���nɆ����\s�^�ȑp�*�I�^Z�5,Z���)*��z-]ES!&���$I�j,���b�������^s'���k�ܥnG�0�[�Q�>���&�pՠ�������]'�2��#���@�e"�@���q<����֓&nX
=l��skXK(p��P����jKB�IDX&ɉ �v����6��Ztq�HbN�ͼ�L*6�j)�M���-R"��B��5�&:�r㕴�ԓ ��!�n<2����Y$v���N����x�M�m��+ϡ�&�i{[�Â�j��p�2`�bܵ󥱉nf�� ���&X�u���\{�:C]E�C�Bj�f�)f�rY�c[d �sc44�ݏ������r��j�0�n:t(�Kv[�t���������V.��W�8nئ%�"�z�ˤ��g*��eY^��$e�f��FW-� h;���ݕ�X(�#rSL���nR��i�Ͳ"8�dh��Ay(�_��G�dY{{@�a�(ֺ���Kو�� ��,�G]i�ުD�k;cQ�U�v~�>@VJpc�)��T�����´�s4DJ���4�뭤ً0�uY�L�ߩ̲B��hM���'V5�K��p�Զ��vƞb�F�G���џY����}���7ڸ�5�
�5�Ճ3�aM*�N���p�Yմ3�!��U�M����T�Sh�ۧ�`��R}J�&$_|l#�U֝��J����0�{:޽���]Rb��RE]cѣY�{4i�������$��>����@\�1�@�]E��|��y�a����c�ۘ���e;�����.�М����82�0)e�&���.�wI��-�Ķ��Xc8��5t�j�ud��:�J"�������� ��7�(m�X޶��`����4�i ���GUhY�h"�)�va�8�J����+	�c��댎Q�`M����:r;:�6�oF�N�!P����
5�6�f�&v�������g��v^b�5���l̘��� ���J������>o���j1po�gIm����u7=�CQ�z���ݼv�BZ��6k�6Zn���Z�y�b�ת�2��%��'v����pl�K�t����i��R:	�׻4]wNۍ�,��W�/T(�#�P��ՙ��46��G��+�]Wg�8'0�[Y؁�'C�,>��s�׼(3�\�ӈ�V֮f�(�V�8Xe�bl=h.��K�y$�8κk�f3�Y]��ꎁ|��z�@�ŵ9�z3frM�$�;@�nP��{�3.��� :�8��k����:VR�L�uŽ��ʜ�_>�O1vn�j;�X� ��WK�d����p���.X��I>����L��Ĩ,ōwܷ�Ɛ�*���Ռ1&��NS~�x�u�}95�#�&�����<����H<�{�{���q�#�|�:�z�8�Q�%3���(�	֜$vҵ'U��J�[�iP�[$ٕս�n=KMv,�Ϋ�����P*v���HZ�݀1�ӗ�V9����]���t_M��bX�䋖���.eul����Z�ޥҳ�K`�K�y�-{9�3'WDֱͩ�W��{ۘ���Ь?,��o�K��n��/��.(��١L��K�G*{�t]�3�1}��ʲ�mn�xx󜲋�L /�U+h|�v<�n}�y�[br5�s	��Ż�f�	�˫�6��~v/v��N�Bx&(�m
��Y�]�O���)��SF�vp.I�O8e���%k� ���O�-n+�o��=����/�1�!mquݠUn;�'�8�Į�י%�m,��� \���S�����+ ��+��6��n��z�[G\���}P�qq̸�)��/r3A��a��{�l����"A�jv��]�}�0G��Zmm���=�f���1о�@s�K;0���f�o��Y����5<
�!�"���hA���yr���J�,��QW�Q��N@�s-�*.�]�����j�#8�x�����dѶ	
���ǊH�$��u��|%a$��5�nT�)�L @s�K�vn�ڑ+ѕ�WI�cK�S���x�,��C��v�.QMg.�wm�wJ��ZӺӧ�I�%.g�a��ޅ�m��2�+u�����*÷�J
�)I�n��2���W�8R��-��f���/}k���$Y	�&uf�.��}��A�:�)U�p��m3P�/p����3�P4n��9����]�e7�]��Z	�X�:G`��9��k3}j���ϐ�3��,so��B��^�[��F�����@��t���ݏ�-����6��(�V�J�x�\�0�''wR��AU��9s��l�9���'�]�.A)����mM�������������4b~ͧ�'�x��M:����tL��x��:TwrPJL@,wtF7`�
d���J���z���]�֊.j�<����#��E�pĳj@�d�Ҟ�	#o�|�7N������b��V�]��i���r����وg3��֝��x��5ٮ��Y��i��.�J�|-�Xap��pY��N<�ө׍��ҘT��Df�����Y���;��G�_@��qa�ы�Jn�x�3��y���G
[��te�0-����t��=B�ӳ_Toն��t+bDcfu���Ѡ��T$�1��An`���3�O<�v��p���	�;W79-.��H�)ά|t�q��!���ͪ�T��mԙ���}T�[��jc2T�`ss�]��U��n��_�<M��q���]��yB��Gy�/aueh����1���ۡ�x5��z*ZH���/N��,E�����s�s �x[�ef����+w�rwk��a}A���3n�K��zo1w݂9yc��x'��y�m���U�{�c�:H��%�ꭝW5n���̄�V�4(�Sy�r�g=����$�仛��1s��XP\�Ou��`q�{�k��,Մd�]Z/l���ꮷ]x�����Ld���h+�ˑ�,,ʭ���B�2 ����8��2�����}�n�A�0���WK�u�h�6�:����s�ݍ�����ܙ���RP�w��
&��V#�}g�X���l4��+�ݕ���p�B�G��ҡq>��;	�3b4�,�+IU$���7�ٹ��n�tj4�8�ȇ3 �0Z�Wё|ë��bz�����}]�2�d]w���R�:ׯ&��3qv�J��u��w\�,n^(�r|&�x��z+7۸��1,��u���Ğ�$��2=Zi���Y$d.􂆃Y�Iy:���Fp�y0a�y�`��j�/t6�>Ǥ=����O��x�W"��־�H�,�F��K)J٘*'�tmd,�E�l��u�2���gD���`���d�oEEϥK[�_Q�t0�K�[J���M�b�=+�)�ⴲ4e����]������x�+�J:�ȳ���344����]}q�AҸ&�u���y���t�X�2B� �NԆQ�IVPW�(�����]cw���,��U�Ol6陆+�� 5��p��؁%V�bC�3{0%}����|�rw1��j��]��1Z6W=S��_3*�sjv�N���V�����#;�Cgfm4ͳB���Ս��_T��Ԯx���Yݸ��|,Wn��Y��j
��aU��]��wE�����m]�������l�sz�`����;Ho!��c���ʗ]�����՜5�;�Y9�y����9�b�n=�-m��8�l�\87��t�j7om��H�&�Aۥ��P���ՋU׈�j�O[+.��w�"��+�Of�yط�K�@�����ب�+�=)�,��'r���p?�.�Da�s
c����Ӵ��z��3z�w'��d(iT!���Y-}�@�ϭK��� l��S)�H�+	iv�Q�9�wS�˷.v�
W��)�hJ� ��kᗝ��X�"��.�Q���T����A����RV#ؓOn�ӹخ���GuS���ˤILᎀ��퇩���Z�WM%MWwn�'.,��yu�{��]�0���N�i��0��QD���wp�*�n��¦tVe���m�pS:�����U���Fo����`F�+��e�4
�s\��&�yI+Ӓ2����1Kf'�v�)�|3v�&
���bo���# ���bNׇ{_nTR��=����5vc(t����U�-Xk�Z��2��ܐ��뷐���ef
�Pj">���gM�[�orV��C|��L+��и��e�2.w�nG��(&��}��A�1�>�&��m� [�<U�2lX#�s8-(��:��:}�o2"�1Res�v�f͊rS��V�v{����d����FJU��-���:YYIT*��Qw�e�l:ޓh�}��s�F�d<c��{0�(�l��B��O�a��ˎ�tK�,vfo�,E�	�7��/"�~�ڄ����M&���/(���]b���Һ���r �H%�V����%l���N���Y���P��L�rn��	���uw�7OS�bu$ה��Ѫ�)Qԗ�j��܈Laj���j��1�l�r��C��21jC�0K�2ˏP��<�^�᥌X�e�A&�9b����%���vh��g�hak�\�r=M�ٌ��UMbN�������YѴ{w/8��5ޔ�	��W�7�4 cv¹lIA,�m�]�k;Tڭ6�Yߣ�?�8t5��:�샓��v��nr��ڳ��{%@�aR�8���R�Iu�����J��ͺ�`8� �w
��]$0����{��=�]5��c]��D5kZ�����:̽ӗ2n�6�rPc�_l�jkC-�ۅ>Չv�+a�dYt�A������������:`��hG;@�����ur�C��g`�',f��ʹaf��(����Uܪ��N�}�ڻL�:x ��5�����]L�ؾ����u$�z�T�k�~k�U�U�(ZA�ˆ��4]K��V�G�>��Kl����bή��[@l/-�P�*�0����Պj��]�k��`�-�W�	��vu4��h�j�S��Z���c5��V�=T��}��c�Ga^����&+WM@�m�O���f��Gk%���J�:搫����c�����Ov��m<8��F��X
�Y`�$���.�������*�����NM���-m�L��x�F��{�y|������WU�:�R�Dt�[���c=N����J�����#f*�ڗ���JS,�$��N�rڙS��v��b��X�+8��Uֱ�Z�_����!�Q>|�8�a(
䶗SJӍ=P$��Ԡ��Ұ�5�7�mPn��{o������$J����{��P���/�]���b�9���Џ�R�Ev
�s(á�kE���{H��������n:Ѵ�*\�Uɸur�
Uyt%�{2��5ht�h]�������iuX��A1�!Q��9�rZKgn<��� �,�AXuTTfE�dբ���=��ޕd�cb���b_Jk�nlGT��fЙt����d���b��N��9v�?���~�J�����9 �P����)Qj�_u�,���M�}�.�E"&�Y���	�Ӵ�
��$��6��e��vv�ْJ��ds�>��<��Y�p\�A��gp���m[d��ǜ��9w��-�u��>�)0LcN��)S8S��]�[Ʌ�\�n���=[�X�v�����"w�|n�E���vu�[�t��)z�q�ɬ�']6�ޕ��s�Itr��7��93���W�����P۳g"
�-��:�pl]�f*�:�($�R��<�@+�oan�*��m3�:�W���<�J�RdC�5��G�m*3b�� ��X�K%Lس���w@���G	���e�f���n���� ����XZ��`e�QT}]++QǏ�,��pZH�fe$f��Ҩ=ԫmmԵwS�t�h�X�Bl!"ŬD��]vq<��L�䵼�[[�@ʚ9��.x��G72�_F)�|&K$p7f^���>a
�w��Q�����o�<��+yU��Kݧv�eHzd����#�lz��j7[E4�������\[U)�=���<KY�*h�ͱC�2��#O��OBe�I2��3%�-JVu7]�x��A��YF՚W�@��5daF�w1�Y5��=�v�v�ܓ���2�]�4�����70JfP8�H��V]v��Uۻ�ٲ�[swOqZ�@ �=|����R�)��ի�t�y�2A���X,vn��zM#.{�p�1�]�S.���`�Q��ɫ�b��96�w<����7���/u�1�Ozݡ	K5L�V�an�Q�-VK�.�L���+�U�� I�7��ʵ�������BܵZ�x��P���Yf�9���e���Uy����rÔ;乯�+���$�E����LZ��e��2G�e�C:����3�W!��ۼ�z�M_=�������F9�e������5�|�g���������R�MZ�w��M�9ũ#=�]��+�g^�FcV{�P��	�v�tD����X��+�Rϓ�Jw���#!9��w�xL���J,1H>ǚ��6p���Y�Z7�I��x��Y6�zRV�s!�J�#wV@��3]��`}�G�__:A��9kV�����%�8���'�໫v�'�l�wB������u6Ln�Y5ɝ��Ȳ��U�U��t�r�sn%D��`�%��"M���[����nwCd�@�\3s�ev��B���3.�M-|���)�� .���/鸯�#IR�&��e1 �L �q���}�1���5��8^D�鑺�g&#�nms5�ϟ�>��Wk�'d�Ǧ��6���y���q�'vLN�!2c��(2I�A\��2����!hѓ$���jV�6��;g��T;8w,�3�5`��NG�~M����7bo���K�m�,DVfJ��i;�}k(��.��F!�g�oNM�P=�S,V�����a��i�z�xf�-��n�Ӈ(v:DS���vd�vxr��Aݣi�Қ.p���S@��A�hM��֕6� �� �\������w[�]�[���a;�Ȑ^�#;a�Z�t͍(�,g(N q�¥��n�ţz�]��O_L߷�pG���am�D�goY���բ�B����N�6V��
f�w]�t!�B��G7��W� cpW�X��˂����{�]�᧯c�X��ڹ͜A�-� �d�0By!��:�Η����8�Lq��c���}/��}��k��Z=/3zݦ�׷��s��wm'e���c����2p��⇙���1.͔�-��H��zY����y\]΅�/3�4.����#�֫r�o���ytO�� ��Q�O/�s�)E�3��l����;c��Hq�9K�4ܻ�����VEý�R�1F�xj���7>0��c�.�f�o.��7��$ �B��汻�����E�$d��� ku�{g���L��Bձ�s"��!���P����kgn�@�HҴ� ��U�,?�'���������_gݮ�n>6�\i�j��d�_���m�j��XU�J�Lk�6�h�	u�;*ɦ٣F����0�j����o�r<�s�'p�{�Öy���P����t��-S�N�s�{��#v�+�d�સ�6q�f2vt���ޣk��𑽙m�,��AJ�͕'QTRO���[���X}lsLR�`/(������WW�p!D�s�fk���ь�\YAd`���}�䖺�E�B���,X�Թ�g*u#Q������=�>��2���U8D���]m��t{�+i}w�7M�n��+�+f�C�X��y���#Zt��/�����C·�YATt,������t���<���Vf0�{��q�ׄZv�3�w@���3���ff=^%�i|��n�gR�fU��U��̤R�A���̧0��fK�g 7u^�Mkq��2f���N�n���t��ȫj�G��7e��펭'H�[��n�5���,��	c��׺���vp#È�뻺�q�2oR
�Ѡ03ң!Qileom=�/]�GN4�1�����Ⱥ��m%0@춍����`���i���tvg'��(�j7[��V�e�E���{�Jw��|��}�9	��E�v�b��e��L=F��*�VK��Z��f{�c�E
R�6д�Hr)�W��3gm^q:��Ȭ�` 1+�Jݮ�uP�
�H`x�C�Vi$��=��m��w����&Z
�p�#�j�X�P��	�f��6��	#�*�V3(�Ieq�E�T��U:X[Ziha6���џm��lG� f��vb��]h�4?!1n���+h{
su;H�N\�et}B�b��T�K�y�i5)� ��rd�o���=:/u�`��%;Vh-/C��9���;G�������]��$���H�y��7m������-`No>�!�l�W�1�Lgz� �W@���5�X���R��_2���VK7w�\a��ٹ �1��t�>��uf%oUN6y�WFt�ga\�v��(E8��c�T��J�6���;-j�U��ԘҩZ��k�Q��������B�$j ��ú��2��|H��ℭ�j�Y;+%�}ŋȧ�d8�K���;ފѕoP
�`��-����!uӸ]�M��h6P���J��(�n��LX�y�mu��ZhE(�F
v1���n�8r����@��:�c��-��Rk�$S���Y��G3��ڐ�C�C��GL��Y,�ܴ���S�D������׹����Ao5uy���i �08V;=�A�nS��&��{�����&s�2-���J�M�ʕ���-���i� ���hkc c�'�]؋����U�u��%�:�ņ�F��:;���(�3Ϻ��f�e�ì�%s��/�����6���z���k/y�����NK�҇s�
� B��ۚ6�5�)&"�V��&�Sz�T�^�Zk:=Sa�J�P�la��gOb���"�n��]�ֶ*��k(�<��j�-[�#l�x����w�^�N|$*�K!XN���A�[��
Nh����+��M�jT�{]�c����$>���+��;WfM��*U����u(�,V�I��VP�`��V�I`�I
�N".�
��
�e��{��+w�b¼U4�;`�8�N)���Ý��yж!z��R�oJ�7Y�����B�3���Vn|9B�;�`���cR=�2��G�����;���;T�Հr�1_S�^!RYV!+~�Y�iU�xui�m��J�p;�q@{>�jv�XD!�Tl=W@�4i���-N���
��ITZ��H�|���Z�L�D'S��YJ�;0�ӜB�I�#�I���	Z��E^qR�ֹ@�v�����aL����T`�xHܽT��A�1MO�pVs���@��Z�	]�e�s6h�ia;�#�օ�%��EY�G�m�W��ǃ,qe
B�Y*f'��'��\�>t�	v6��*��&�}����;�[��V�tʹ�v>ŏ�jSpf����s��p��)�[�]f9U}a:)h�3P���Q��ص�Wz��Jct���2����*��ۥat�ZS�0�:�~�@WBcOwv�������o�8�,B
*&���OnԵ��&#1��s�uh�"�n�����%*�f+�͐�_u�9�+rr���~*����%�~����[�蔖�^t*���D���o��۸�r�v��@	걧6�Dם�^vSD�!�ӷF��m:7���y �����3����;�Pf�ֈB��ڹvC�5�
�7`h�sPSz�^�L�]�0�P��+���`�]��9�����0.Z��LCN��Y��2k��e;�����zi��:�\�Z�Վ��ߢ�h�1��J�j�Y{}-�)�<0�Fk����.͛۸��n�$�],�#P���<�&��0⇡F������Wuf��毒����^�z鑑�� e'���˺3n$�P̡���@*8�����F��B��IVn�h�D5|�ы�$������1J�2�qI��բhִ�Nk�����|��-WR��5ok�U���ul"���F���Y�*T�X:e0��1���v� 'fnJ9�U�/���J۔�����B� ��d<�$�Ni��'H#�e;d�����KB8�����4�IT�TEg[��^)��0IsK/~u�M�
_,ڡ�9M�o�[�ut���.HMe���&
�G7��<i#[��{������O��0�����ӄ`�G�^8�T�׋fꛤ�Ղ�Ae�m��qa�
F��V�����^��h��3&��3OV�w�(�8J��n�2W#0L�|k���99 $�:4��psLO�CGsͩ�H��%6�0���6"P�W-kf�2��M��|M	tq�č5��ϙ���ȅ��3bFWLg(�\q����{b��rk-�ʍ�s��ǘ�9f�Z6LΧݚ���V�ȫ����I�:���Lc�	��h�lϥ���GK��qP������n���x��.��lg�ی�E��uGK�]r�~�e �� �ϔͣ/9�]/;n�AqX�-�zݞ����4�̖�8����V�к�<�e=�p zQ���>f)-0E�Tٛ�Y�X�2�ϲk�m��t�v�l�m>r��b��V���
�<`�z0I��W>8u�R�j�#P�� �<�{���[��ַՎA0nw.+�q�H��iPM�Z;-o�h�v���u���v-FNQ �va��Du"�5t���;3�����A��p�cF;�	�X� ��K{7-nY��P�Ύ�;���ua�1������pv�aK�d�c�Tֺu�V�7���z��-My-�G�td\D�xl�.��!�ݐ������u�Z/I%
B,�2e
��ں������
��n�Y��CF���S"�b;j�N۾�}+29Nݻ$�� ��V�Qљ].�3q6ۓ�l�֦Z�Cu\`�h���z1�rY��Z�_E�YqT1�W�^4��,
wa7R��f���]$[4���Ea��O�j�z̛���m�wf�
7WU�a�E��R\����B�a�z�1�,Wer�Ԑ��t}�w|�t����F6�V�7㹺�,�����Ub������1c����KUԁ�A�m|�}˫)��6��q_p���P��)���]|���VsE��˔���\��H5�z>�����X�np,�LO��R�͎�9YJ�7ȹ�u�r�����������:�3)
H֊�a��4/Nl(IIKW��,��&���w8��[��w�K������eŰC����e��9x�߻]�#�ZR�����|%�k�1��YS2�:"��râ�e�u�7F���0���(k���e���Q��7\�Zڸ1�إi"����
g:��-O��v��D
ʷ%4;������ #�g^�0�z~�L�%n�U�����Wx(Eo�]0oF�Y��Z��}���!��^1zB{�)�]�|�9������4J*�\���t�YF�����XH����iм.&�h��;&c����/+Rw�J��Z���l(Ap�J[�nQ�IVV�h{�m���q\t2$�ۅ�A�e�`��'��
��M�tӸňRj1zm�qC*m�島[s�b똇���,�v	�i��Z�Qgu���[�;l�s�G����^�q�H��r�@Ѧ���(ް�ev�j��#��fH��VM���
-[T7+, ��Ӟ�(�*e][��8hJ�sn�s6���r���l��M�LjD%�E�3�.QLә�� ҉�ʑw�-J���Ry����ޗذ���Ⱥ*�k��m╆�	k�R��n�k���!]omGD]�:��F�9G!���Y���.�E�<�)0�Sp�( T�h�7nSb��Y���$rq��V�_�3$T��Cܒ��<�Ы�<R�EM$�e����8i���ũ�[C*AV�"��G�9�Nr���r������潉@����Y�V��+NksVZ@P�f�˒�m���r��R�u*7SJ��g7ݸj�E��=�\�c��kZ�}���N�9�)8�v�{���� ۥ�H,%{R��L�ʡ�. [��َ��y�k�Sa^:QZ{�m8C����������J�n��*N�&��B��v7�; �`�|�L�����-��t��T6���p$�1�5�p^�c}��s�A��X�w��*��fk(�@�/��X�K�z��RmeN�iT�n1jNA]=Y���j���*O�z�;��S�N��0;woS���y��U�H�ƸgU���ú���'s����n�4��*�r#$v���`��-��ָ��֬��+/��ۨ��M�@��k�����;6�}�=G�2�l<3�N�;wGhB健V�,�� A�j}tz�9}�&Fp���D�Za�E9�ޕr���G�VO�1p-��I\�D���{��:wI{���5t��Z������w �����hJ��J #y�XU���k鷶�p��lZ}X���[[><9��F�8 ��:�!�3,�l��H�<N@��R5�'E\���IE7*��p�&��������f�]V��*������j�[�r�� ��:ѡ�3������#��b�\��wփ%���W�$��[��/Ve�!z�s�8rWwh����Ѽy]��Q%m�o�'��y�^g�Js�]��������DjEti#4n*U�/�&���h��/+�)n 
x�CoN�g1t�ڕ����p��@��ͮŖ�e+�]o�dΟevw:���}h@���Y2��{sox�N9X޺N�غ�Q����)���Yf�(�˸���poG>P�W��+hRw����7��v:;&��g��1j�o��-�챌�cX�%Ώ�tȗ��niAht���J�3�a��\%��t�q�T���98wj��)���K;N�޶)��ν��r��ݦl�9`6>͹8PjH)��d���r��7si�|��(��d̠��q�w�C���RS��ӜNs޾�8��P�R*������\��5m����Ch���]s���b��)���L��J �i���of^V	y1G�:��=F]� �6�:����c+:=�k�[��y+J	8iv7n��R�c����W!�!�U.���R����[�Vĳ����ª���_Q4�wұJ��j�=c��1�\��W��*u�l����c)_X�����{H�[9d�2�I��!.��r�2��v��v�	>:*�ol"��MN�e��Z�2�n�1�� O�g�#v�TuZ0�{�����P�&����ߔ*�M8ha����d�n��ʖ�t����X�$�ލX�1��<T�ܾ��\YI�Q��ԝƩ8 ]U�B����{o��ʢT����]b�/���S׮�^|Q:�A�FЭwB���Q��r��d԰5MPk(ռ���9�r�X[k�Ø����Χf�F���3j���n��V�#�0M&h�i�U3�p�`�bf]Ԓ�S��˨vf���n��X�;{w�`IbÌ�*�%���A��5)5QWK������f�A7*'H�M�tD�%=MФ���E����k�nm��f��'J0�!�b�&���C�"U�p[�t�CX�i[v�5�(B�6Έ�
uPi��J��K�0]e��(e�j�{��T��#b��Kn�)hHn�hvn��*�kQ���MP̹9VW5��iAr�ғ:�'`U���S�`�cK�ѻ�?'u0aP�tqRX��X��Ϗj�B��Ttuf�� j�Hu��t[�(��"�y����05�]�u�&��8�!�(z��݃�)K�ӧ���ڨ5��)^�c�pmpH1W���*2
��������"K�_-��u�����s��2w0;'ö+i5��$�{_K�e*y�i���U���4he�9�ڑ1%:�G��ٔx@�"Z�t��Y�YW�fD`�l��:JӤ�ظ2h�;��۱+m*���u��[�/���a�:j���Ҫ���]!�7��z��X��4\F�V@���3U�bT--<��p�u�s�JND�IN��\�)��M��Z X�g6���U�\�G�2�4��"�tx�;��bT�z� ������n��UK�cs�}�j���$�	'�:s}�߹��;���!q��|���w٥�} u��,zz����rY���ћ�qe��v�N�ܘ�ߖ��)^�#t����w+�v�Һ��������v����
�<2r�2�ӳSw��-�.���M�����������b{�5r��N���b�ٔ�᥹����ծ=|�U�Y0�|�ݳ4W\M˫�Ī�Eea�y�M'�u���>R��X*���Bʡ�+7y�On�:��̡�Ch 1��N�6�wZ��7v$s����զ]WQ�\��'���[Zj�;. >UR�W�M�^�X����/��t�KR0����Z�P�3S�|nBv*�^U�1�;�މ�n���<u���
�J��8�����j|�ܐU��E��h�m5�R����r�G�e���j�o�eBU��[>�ҷ���\^�Tf�V�=F�Fftqh�+)���뾝,��G��E���0o7�qˁ��ݏ��}Nw]ε����k1TA�H������\\�ܽI��+�_v=s�x/�₻��_X�\V���2T	�O��Q�|�A�K�J�up%WFJ ��"6��E8�,V�0�Im�M����q���*Z��PhY��Mt���	P�y���휶�׶%HȣS���V��7q4��퇟syZ������ҷ��6���]\p ,Rֹ]˭H��khڵj�.��e=���j�˔N��:k���I�Fn������NE�����J�<-4��+nt�7�N���`�P�h��)m�E"1A�V�kX��j�Q0�TQAQF-�.R��(��.*��8j���0KBѵ�"ŶPQ�Z(��ET�TU�UV�EH�F,Q��UTQ��E�lYX(�R��+��

ւ�L�kUkEcie�c-�[U����j����2�V��QQ-���"�m��m,�iA�%X�b�%�F,��`&U\Q���EQDcUcQEJ�TED�mX��Ҋ��b�(���`ZX�X����#�EAT�+�X[h"T���)iJ�jQ� ���(�+QUAT+iF-e���U���JA(�n.0�,R,Tb�����h�U���1J�!Yc��j+iZ�T����b�1UQE��`�RՃmDDE�f��J�`(�!m*X�b(��E#T2�`�T*��X��U��R�*Ԩ�ŭ�m���b*����L0�[QQETF"1EAcR�Z�ʑh�ܙ��\��o|��|^iW�`���dQ�y�T.����[++/%���S����`���_F�s�oo�dnE����{���5�Ow�T?����vzׁ��C͒�c�8?���M-|hj���d�^y��lק�yzQ������
lY�=�\m�D!�1+��A��jSVvl�0]�xf��+;V|���2��Nrk�UD�N}P���� Z.���N0ȃ�t>ޙ�vF��v�g�*S�.Ɔ�51K����rm�IWE\U;S�|�-��C�ȓ�g/�P������K̵fG��%�B��+#����4��D�#�Q�	�^r���֡x+s�)�����Z�
(�ap�,��]�ʑ�3U�����m ��Տ���'������'���O�J��9w�������Z,���C�6/��^B�w���s;�00�ot�aT0xA++�-�
*�]��G�u\d������>
�;�F��9X\e�50�s�q��)g>�c�%�LC�<"�2xޡG���~�� �D�bS�^%���cػw|�{�b1�+�bR�*�P_/ja�U'�A��wӚ𩾿x�����s�\��s��O=�,�M����)��'�3&�,*Z;�iZ�/�k	��L쭊lɽ�nsV�ì	zW��)|�WyF�S���좆������a�u_k�q���x�g�qɖ�m�O;4�7O9�ve(ih�+3cUM��t�qa��a�)즞�ͮe�ðMg��:�0S�(i����@U3��q1[��8����`�v��hl�r��to:��x��'����\d���W�������$եμ}%!gc��(�U\|F�_u���+|��Ύ�<n7ƀq�[;��w�e�M҃rD����Dp��O)�d�Y�g�S��X$��}�H��u&Ϩ,A᭔9��|"ֽ|�G�q�1�S ��]���ݲٯ����"mN��*��_xM�b\~{v�"�3��;�eQ�T�!�);����3pIW��H�U#�����wu��R�����͜�,ϰ"BB�>%u�͙8]30�[:V��;5>�x�C���^CQ��f��=�x�ʽ��
�&��tG#Lj"=�<���誺�H�{���p�3Y{�9���6���5
�$�J9�e%��K�����t1gr<�1-��/v=�Ƞ=�	��u� 5�=9����s�P|*���_���ӞWK�W��i-��
��U���6JYz��cT���u�6��������{Q�]ĭU���	�<�9���Ky����^�H�X���o_h]F����F�7�GR{Q5��&wǍ�bw�i]>��<�[� ���љ8Mƞ�ew#j�֙�\V���ד[ۨ�0�V�C�
�;l���Q͚e���;N�!�Ǉ-�#�vS�<��f�oq�`����ʴq�!�Њ�/��j>g��zhK�k��KH�e����b2Oo=�3�ܫs�].+�E��t!+��:�'�����-�
/�Eg{V!�c$�����s=��u"̜��5q{2P�����5'C���n��>���T�[Ɗ��(a��=�'�z�l�-1�����>9[]z��\׋�8{���<{�,�^�%4�_�{3�Y�"��7~�>��Ѯ���o�N"�b�=t�N��!�7�p��Gy��'�`Zdt|����7�J��Jlc7�:�U���u��ϳ�C~��[�=Y/���w��)}�Py�v��Y�t\bNf��8g=p�V�5�Lk�kZX���FfWB<�oݻ�Ԙ;��;}~FN���8���V&���|e���j���x���fP�J�����caQ�lX4:��t6ܭK��;�~�C�*�eO��!�=�k�3����G7
oݺ�ǾN��}�Y��*��c�����]s܈���z����F��n��m�u�\;�.�
�|�Y�|Z&s���1��ܧh���{���vn����q�[̈́����7�����y/���K�np!�͎���rC�>�9�g=����y��w7w��)>Fe#!U>g�^�����Us+T�k˪xK�sm�9�f�U3��q����"ۮ�^X�F�9�O�>�v-]�t��򒹛�N�Ia��ܕ��S���ȶ��5�n 辬j�O_���l����}��g����O��4�>���t�k�О
B�Bk��W�G�kJ�>���������E2'��qV���({�UF<C,fzg��:w������P���|g�<v��/2�!�U�OUvۥ��ޣ�uS��O���X�5�%?fZ��N��aY��h罨�Vƽ�Y�T�V%�--���yc�T�h�(�~�$���O[��>Zs����&/� آ���S�L�6w7�L��{ѳ���W�h�
W[����z0{%J��Wm���6G��ӂ�����yG�g5�S_��]拉����b�h+G:��}t��It�oc�f"j"D�W��g3[J�xr��\8��P�wr�*��Z��)��0�Q۬��&�;&��ɗ��¹0Z��v�a�2iΖ��M/�8Vuު�e��KQ奤�+Z��i��rS&v��!�މ):�/����9��뿞���S���u͞%��/}�����\ۈfn�Z��k}{K��:������L���>@j�^o2L����y��>�[MS�k�~U�j%�n�v��z Ƃ�{�q2�ᓝ؛��P|^���ڪ5�hw�C����b�u{.�yjm��5�r{���^NIԑ��O���5A��]�)���4	��Z�읯.����3[S�MkVRra�����t��Gԝ�<cy�O�M�w|��g%�r�Z<����'��9�[�h�7��7�G�]��^@Νٴڧk�ﲫ<�mM�&�;[6 �H
�}�9������f�Yw��λ�Ϟ�,p\�VC�3�;|��-�ڸ���W�і����KY�χ��v
�q'B{����z�1^|�����6���S�8�K��KR�*\8�mg����k7�]BrJ�đ�-+U�������Fwh,���V�!�[�k5��M�݅�3NGfK�F��q
��Vg�U!��ž��6�=�m��dɍ��&��Gbe�1u����W\5
<z�T<km>�pg=c��_	�\�h�<L�f��R'��S%�W�u�Y�
{�g,/�8?g�����ԫ�7�uݹ��z�`m�t瑝Bb!�=T�+�Tu��&j�?_�_e�U���R��?��U[*={�{�k�cÝC>S؏q��w���Z;��<n�v^����z�V�I��yhn��$г�y�fa*O�sޔ��ҵhxx!�I��y���q�������m�t��gG.�r�F�M.�m�:\���*;-:���w�2���brsٚ��q������V9��tft�۶���ST�S��T-{�-ٍǫ&R��gH�����)4m7��������%9��ͨ�=�Nd�ĥ[}���xhr��U��z;ݕO��7���#2��O��m�V􈯷����bO{�Π����R�:���ٟ5=�U&��ڤ�5�]⣠��A<_L?d>�!u����v/׽��#	�M�Z���t��B�$B��kj�M��hyo����D�w�4���*�.�M����o�'���]�zl(g93sS�t�;ҵ.���bUt�}9�%C��3U�{���g�: �aR�.�^�+&T\w3Wq�j>s1���neh��p��� ��K}��6W{�O�h&{�$9ڽ�3�q��U�e|+Șj��ЎS�z�]�$��R�/O/���򬷎;�W��}[+(�䑮�#�,D�P��y
�ap}Z+:�^1�ڝd�n\�%��y��F{՛�Y�d/�8�-�T���p�� tb����
op�������K!��>�A��%g�_��(E�jq�X�J��O]M;�8�Zu�N]foO����\����ێ�o:�]�N��IZ�����b6���=�P���r`z�E]-�Sʤ�q{��u7� ���Ԍ��1͍�߯��^Ow:ǐo{���<5?��u����w\2p�󁳈s�3� ��;�{U����y�=�Ӆ�rX��kkҴ[y�2�����_�(]� ZF��۱�u�;������~Ϥy�^���))xiO�}nV���g��r'�����g�> ��)B���`2o9!H�3����=��P�+��j�����"L�B�ذq# R��,�~�����7gI�H[$�`�k�W����,�ձ�wv ��+v3�[o�8�����{H�y����OW�[��'�%Μ_��/��7�OQ��Nt&7�{e���<��ʟ�J�����Lj��jd���{�{�ϫ������^X��Mm*JT�ںr�Q��R�|_�ݑ|���8&{S�u�w����I�ۇ�ǵ	��[�t5\�Ǽ��s�ϥt�2�^6�3���%�6sŊ4^P�ߧ��h%����*�܁pfZ�i��P��z#���,��~N#J����F��ޥ��
{���|�}5��oso~�8's�K��}<�О�h���\�g��R���:�c�����ݦ+���ϰE��O('E�;�"��afk׃��Ck�=�Wzz����|^.Md���������Ez	mV��|2���)ݹd_�����u�^L��6��:��S#U�*�Գ��x_:f
�t�]ӓw\�^D��p��6oa����B��o g]���HN�WfvuSC1n�YVt�$
.v
2������3Wl�쬭org]9�!0�e�%%��p3t�.}�%+ C��Y/gj���v�'vؼ}��HSa��	����q�	N@��k�o�ԛ��
ω����s��^(�B�B��0����=�K�F���fc���������ws4l}2(=E��{"���S��63��ƽ�M�v}ͳ��jT�YA��KzvOk�*�����������66��}W�le_���M]��;+cO.��2*��{<���Z��|=qs���H6�����2g§EFz{:6���p��,a;u��i�*�|��㷔���Ӯ�n��g�\�<�����<�rw�����)^}�]Nߝ�U��H뿔�E�~��jhc½^���gmG���o{�|^WOG5F��ý��;]|��靊����5�Q���g}����sЪ/C��-L.}χf���^��?[��^S�m��rσ�M7�ٳ*�j�����>�IO���6}���ࡱ=d�S�,q��W�	��+�A9w,mqw!�(v��/���.�R 0��x���f�{ibn�X�{����>���(Q�Uՠc��"�U�fh�/����b�h7��<C�@�A�mtTT�_[�u�)]����E}��bQ�x�~�CKG���j\���z�J�a���r�Qu	`���˺�>u����C5�[���O)s��g�h�П["�V�y��� �Q��Υ�|P������Ρ޼H:���$���[};�;�q�"�8/�/�.�֨�x�om�����7�f!|���:��>=�98�����"�.Ϲ_�Ro�����6��]y��f����zW�T��yb�ʮ󕮦��̿���%t�:�h�Mɵ�<E��`4�e<�T]��K���9�jyյ����r��v��(��l�D��5�c�G�?#b�����PK|~ř���s��y ��绎Q�'��z�o/35G��":���;������[�6�/��C���n�uʼ�{���]y�3�s�OvA����9E��>q�y6iUf��������N��N��msT/}�����s]���K}V���T���,�������D�+��A^�ʙ��z%�k�o��L��P��i���l���s�]·_���U�LL��<�j�Qy(��;CJ��pNII�m���z�P�M(^c�@).�2,f��Kb�#3��<á�t:�dx�d�{&��MU���2�����J��*)�M`6".;��㢚�yc6���9���m�bbZ{�8��'f�u�d�R� ��T�,;���G*�㻖K�!i۴��U�n�a�mi
�f'��[/��i����wm�=b�5wX-��9!6���������R�/�L�.��Y{*�]Gв�������I>�����)=��L��ۋOŜ;z��9��z��ėX�݂;��1f�����O̗1:ҭ�(o\��9[�ʹ��ѣv[�&>л[�Q`�M�ډA��Yj��%�:��Tywӫ�гBj�j�s�BҜ�p�w'VDph�V��(��)/��
��(�"�l]gr��<���>ޝ�C#���V��Ǵ�k/���.S���)�r�J͵9��W��j3�An�YK^Ar���؛-$z��4&�T-�-���kk�^��d�����N菚-<Չ�r��|
4�h���G���}�y���ɒ����宮l�+y6�.�ҕ+�K�rXe�mgY��1̽f������բD���QK$Q�0$:�i�ǚ�ܙՂ[���|�����3i��Jå0�4KkS�Q'��V*��ٮ���m̶��,(v��n^p��O���6Y�|A崷2^��}�룛N�"֎�N��KS���r�����Vv�OR��U2 uϵRe���Ԭ9so��V���\��UЇ.������,�0�N��)yp��s��뫘*}Y+�6!=�f��j��e��#4�kܬI�}�Z���V�:��;a��������;�I��|�,�`}am˨�&YۮL�Q}�]1�D���ln��:P�QWQ��Y�{BeKt��
�����{yB��Mچ�He#�N�j����U6\�FT�LpB��Ը������42բ��$��$/�.���=�|��,hiQ�'%f���)�0�u(�+�-�_i��ֺ>�
�6%�-\�m��Q&:�G�TBtʼ뉡4�%�8�S�-e$���5Ta�X]L�\l	Btm�Πg �к}���%�����9�`�rk�V���g����]�6�,���G�����X鎄J���N^5��.�N`0'�ީ�0�И���6"���m� �D�]yV�q�Q��T�¥���V(�V��D ����d���!ޕY�q$B�^64-ӥg+2��X���^gf��*�.���U��k��Q]��R,V�M�ϻ8s{�a�\3�uJp��)/7r9�Vq�Y�3(�  (
�QOԩ�cR(T>��F4Qb1IZ�QUX(��m�����E�U)Z���kTJ�jV��b�j�X*�R�(��PT*4�J�EX�,�U0��TkUX�(�+)l��YR�,Q��,[B����2ڨ�"�ֈ�J�EQV�EYm��b�X�5��c-���p�b��ba�Z��U1eT�(�V����b"�ckQY��-��H��X�("���"*1�ұb"����G���Ա�2������2ڈ�
(��1cF�V("Ե)R�UDA[h�QA-��Qb����YX,b��b6��UU-(���ZX�U��,TE\ZKk��[�T�lÈ��F+���T�UF1mV[U�YRƴQ��*ƥ�(���kl��e����[8a��b֨�U��KU-Z[PDQ��h��TETT(��+i(����m
,�J"$kY\5�Dr�Ce�YKeE�T3�bڶ�DciJ�TKlkb��Ţ(���L5Y+(���*�
+0�I0!mm�*Vb���(��X�+hTV[X�VҨ� �"��P�Tb�B��)mV,-�J��Z�5�Z2�kmb�U�B��X(�UX�����jҬ�l۝:n�n�q��eN�s {C7k�g��ィ:�9ι˚���n��v\��}ݖ�i��k�|�Rsu�"�YJno�,���f�k�MԹ�
���ۂ�>y%C���4���6&Lz�r�e�ϊ}��Q��gh���*�P^x��C��?T��_=�T�[�����hIN/��VR��OkG��,�)�5���`��i/�=�;a�=�Q�y���y�=RY�N��=�qd�k�b�잍��:�y����u�oDy]�Sە���'T��~f�;׶�����[�����a~���P�O��;x�8�Wx�4��w����F�j�NiS`ԕq:`�^�UoR��-�"��;H�����A�����|����2�/��i[�˫k�y�����-7I��]�o=����j�G^�i�pJ-�S�"�H�z+;8����~����o=n����n��L��[��꒡�
� ����k5=�۞�o-��J������5U�2�j����u:�|_�bL����,��F.�ߑ��V�{!}."�W{}˳jZ����@.�h�X@���A�&�K��kC�X4��nn��]����Lf�3��tE�9�y+���j�,Ε}q[\�yAs�">�e���`t���T�q��S�������Ac�&�tĽ������t�;tJP��noϪ�s�� �w�mQ�YEw|������^��8�J��Fצ�o=�ے��S����koSδ蘂]6߳Sq���{1�z�Um�G��������%^+�-.�#ђcY
5��jBs��S7��U����1�|�~������T���H����� ��ڔ�y|��S�����^OTr����S=�p-�.���:�_t��S�1�hfu��o1Q��=���z�*�B<ƈPcE�\Τﲲ�Ǽ��yϡ|fq�t�S�u�Gz��[/l�1Ey��յ������>�yϤYj�j�ԛE�ϧ��:�h�pT:$9�=j�;\*���ld��cW���RL�3UTص[�kj���Ku���%�a��]�]�ηd����C��b�x�d�mPu��B~/U��ز�{LJ��K�ݙ��jĤ&�6�\�1�N:����h�'H.��S�#�nr�(`�����x��ݝ�MC��ɰs��2_+7y�"��f�h��`�sr1zs�=�����+s��E�M��s�!�VӚj��e���0��z��=��'�uֽ��V(5Nj�v��d��w*({��y��{{��fzt6�^hp����_;�ꏽ��R��,I�雯5e>k�z9&��h���d'��z�Ul_&*WP�rn��g�&���S)��e�I�gfk�t�F���U̹�z�<S�n¼��˓��|*�?W{��7[}.L8�A����d����%���Z�u|
�?b�ٺƧn砎�gt׮���Q^}J����c���(~���]�Ҵx�g/��~�xb2�,Mm��x�n�|�����1��N��oVЙ��n�e�-�+�'��7=�������Py��m���9���h�5�J�d;�~��5�9�**|���xiU�e�u��pw�Oî!�f��[�%�`�F�xU�ydf*uc�;�2�.�ͬ������H͸Ej�j�+&��i*�n�Kx㗊\V��d���|�ί�T{�t��1(��]�nm\�օ�A��a�:e�Z.�N�;�d-��ǖS��u�֎��-��g��V9�'E�j�5�X��(��܈�~�5���q�n*�U�N���)v����Y>�i��{)����z��=͞���7�W#�θt.[��+��z9����G�Şs}��^�����vS�7O��Y���US�~����M��lY�Nz�q{D����U�l�k��}��=�R|�*�
�[pWn:X��+����|}�b�^r���4���`k��I�aϩ��M&�5���<�����$｀c�PUnm���(~�n(�q�~_�}�m&g��6�����sd�a��)>k	�X0��L$�'�~cy	�CHi��2�j~��)���2N0���w�;r�:~��>��}��	Ӕ2ɴX�pO$�L5g�!�
�&;�͒u��b�N�N���&��u$��bM0�!��<ɖu%��������u�;��o���z��8���<�T�=��$�}�`�h�5=�@�&-v�y���;����'��|�v�CL�ɏXy�X�E��/~�����yy��Z*��5��2u�I�r��d�.����I���:�%f��d:���?v͠~dš�s+%d���mI<��P�>I�Mo��s�Wi��[�o~��O�0;��'���4�����d�,������<��i"���~�;�$�5=�C�>k!����ɔ7�b`V�l���i���h4�wܜra�ݓ;n�p���^��:��\C�v���Ͳ�O��/l�F1�S���de�L����q�"�C�d4�l���񍟝�y�elz�q�Ǎl�r��[����nt�_m�ϭ�Z��TV�ڷ��!D�\Ff��moX����~�P�`zz���&�u��hy���<�?0���O3�M�!�Qd������O56v�����߱��0�n�R��n�y~����:�O��#k,�'�k�XI�(qi&��ɦ`T���L����	�2ɯP�	ğ~�$�L��	�O"ɬ��'X��g�����s\�:)�����\��s��=0�����<��q����hm�a�;�a�$߹������e��<���M�c�I�M�u�C�$?}�/�7�$:	o���ڼ�����Y9i��`u�ş=I6���N��8�,?{�fI�0����������HV!�O�aX2y'ƻ�d��}ΆL�9��f��Q3^�O!�ﰟ��}�'Rz���
������$:��4c؛z��O�� |ϙ2���u��a��gY'��d����I�}���� =?~~,w甽�ͼ���}^,�p�u�ϳ'��q�2�!�w������=�V�w?3��a�E����I6�a���P�	�?�ٿ	���<��{��~�	 |O֓L�E�@�=5��I�M�	��'Y�48���]�XCl�~��!�a3����i��`�a�L3�M:M\{�ν���礘B���Qd�C'��|�!�O2m��Ƞq���3�N�5��M>I:��kq3�g��̓l�k��?0�	�~������Ϲ���5������c�Ci8��3�1'�&Oz�����E�uôY;l&1N�m'�R�:��&��Bu��}�i��a��6ɔ�g������ϰ߿���wO���:��L�$��{0�'��{a�d�,�=ćY*��.RO$��`}i&&/P>a���͓��i��u�־��|���r�8��ze��WCY�I�%"B���d+o{L��2�(,Pe��8V����|�W�9�KOk/��-�l��՞L�I	[�	O!��kn�.��V��])Bi�:��;ʞ.T��Ɔ�*(-��΅(6���|*�aٝV����OJ9�}���?�r������gY4���Y%B�Ghy��u�bd��Ow�O�0�;�`�*��Œu�NQI�l']b���O$��w{w����8���w�����|ɤ�g>a�C��6�(u���0��d;�y�q
�N��Y'��!�M���hVO̘�=��B��̝����Oa�+����uNVU���_�#�0����7����Lrì���L��!���$�a�s� ��N����E�ə�{!�Y%M��CݡP4�C�\��߻�������������
��:s�2V�Mv�L�!<�ń�?2}���'�7��d�ΰ�����g�k�bN$�'��q$Ry9�t�e��y�k��ۮ��Wy���=��?2n�{���Xw�d��=�~j�)?3l�a��	��jβO�}�8��y	�w�d�cvM$�'��-��m����M�۞e���}�cП u=9�Cڤ�C^�����!���!�L�����P���,�a��Y?3i4�Y�Cl0ɳ^��$�?gu�_��^������f7{�����wp�����a'̝d姳�Bqɯ{�&�~��ěx����hm�C������m׹�d�031C�$�g�he��?wV�f�=���{|�E$�����O�I2~�I�O[S;�>a�Z���Hu���;��u��z�Ri�	Ͻ��I󄟳b��M�g��d�8�s�7x��~�w�g�~���x0Ì���<f��L�g^��O�g\�:ԓ��:��`w��O�<�o��C���=���	䟹��>d�{�̓���9�<�=��g�c��Ƶ��ˎŚd�OLy���CX��2��XT��:ɰ�p,'5�'-�s�I䟞�4w�Hu�����bC�3A�c��'�<��3������1�����ǿg�])e�7X.��*=��HbXGJ�������f`�5��'��N��n����g-�FN��k�ӳ����k��f�\���47�v)��pQ'c֝���sxdt�-b�wt�=�4�G�v��~�&1`*���2�8��e�I�:�\�!>aXd7��Y�I���,�E��6����u���y̓��9l'Y��N$�����P������O��=D�Ƈ������_~�m�RO}|βi��~�1'�|�y夜B���QI:�{b��P�8�l��E�I��1���)���>�y�~D�1���k�eQF�<���I�u?w���a3��'X�����d�:��<�3�`Qd�fNؤ��&^�m��ɫ@ય����xSg���W����_�o�^/�&X�y�W�N!�$4Ͳe3��8�:�'�w�ϙ&��\��>CH�a�d³�:�d��`Qa:�'��q?Wߏo����g��~Z�����!��TæOf��C�4���'��0�d�!���m�$�4sX�I�5;�C��$��{!�O�Hc�I�L"�풿�#��j�r���+6Ϻ��s_7jP��>I�����Ł���'�d��0̚�	�d57A~`e�P��a�g�/�'����<�I���b
�_Woh�u~ؕ]�=z�Y�;����O�1h{�!�
�1�i'5�,4�a=���J�36d��3�i�=g�<ɦu'�s�Cɯ����+�(��݌{ng�iR�Ek�I���/��Y'Ͻ�C�6�C���~dŰ߻�@�fc��RO2q�~Bu>�	�~d���:�2͞�e�a3?SiH}��U�}S@�|U�]�~��V{�{[Y��&�:����$Ry�!�XO��=�N07l���d���ﻐ*B���V̝E3�&�y8�?!���P�I�����y��ןy�k�������4Ͱ��?!�N��Ϩ�u���s���'���w6I�|�!�O���i���'�,=��T��o��'a��b��6ɦNc��>�n~�p���ou����K���eV�+�L����J'�ۻ)gb��\(ؠ��
V5n������D�"yuĽ�7Z5E�0�u�{���:V`t������u�Z7^!C4y�[����zd���+{�]��o�w��H��� }s��#�w��}������{2<���o/���S��y�m~�$���'uNL��$�'�?w����G��C���7�8��q�����i���I�$�<��_����Kw��;�}�O������˪=�!�&��?f�m�Y35�N��I��ĝE$���:��X3�C��v��{�O�M�'��0��`:���Jy�ƿgo��/Ϯ(����~�������Wu�a��q�=�d�6��,>C,���?�8�,��Y'�3�'�a>y��N�v��'y��Ϭ�No��c�v���ǌ]���1��N��a�>��<�2e�2Oزp��(q$���p,�f�Ň�e��,5�C�dɮ�XN2k�O[$��ݓ��������u�]�cZɟ�ξ�7�`a&����u��я`�:��d߱�8�2a}�u��!��C����rbBd��'�?"�X�>I�L��̓��[�����c��\o{���_Ma2�',�0��`k�k!�R~xΰ����'�I�cq2a�O����q�CGlY��gY>E��8��I����-'rו�S���<�6�UU����S��！�{�䓩�͓�|�׾��I�q����a2wx<β~f�=�'��&���`'�T3�b*�:�s�_�U~���nd��+)5�}<C���P_~�hd�i�:�+�	�}�i<�u?fÉ?3�O'��̓l�~�����$��be��2��]ĝCL�D}�K���{_>w*�𯈪�[��O0�h�}i&1z��N[&�'�$ӣ�I:��3i<��9>�6ϙ4�͝a8�����i�K]k�w_�h�6�x��o�{����8��<�:��L"�L�:�dϽ�͒y��lR|��3�0��L����t]�'��̙C�4��e?^�`�G�5�?K��M����Q�[9��:�P����|{�x|�j��V����g�r���[Y�X�}�TLt�ڝ*��9�J;���sU:pt�����]v��0h]��Ƌ{kN&3�b�n/{X�ɂM4+:���O�U�jp������V�jo��1�u�~aS��q3l'��s��i��X��y&�a�d�pC��C���8�](v�wX��W̙͇S������~��T\��Qn=^���q�ֿg<�W�Ğ=`m�u;�y��*|{؇U�y5�`8ɴXwP6ɋC>�$<�Xd�q���d�,Xe>a;�����Lݞ��x�q�~����2�0Ν�	�>Bh�?0�'�ğ��@S,���H��}�bT��'���&�	�{�~dš����ǻ��$�'���s�c�~�/�������}���~�����u&�~Ol'�y�?�ba6�_��i�6�!�N�ɾo���'�y}��I�߬;�$�7=�`|�CG��l��e�������w����/;�_�\�{���X��o5	�C����M0��hy��߱:�6�_��<�!6���E��;��u'����6����؇ud�e����L�{��ַ�z�s�Cl2�	�w�>`|��=�`�M�9E�,?02��6ɦu��Bm2�α쇘N$��VI�o�'�dѝ��@�'m7q����~�w�}�~����d�<rϞ��a���u�����{�0>C�e��{��I�sI�?$71C�d��!�Cha�=��6��{u�q�|��o���=���������a���=���@�'m?L�`y��q>z�mǽ�u��2����̓�a��k��	�jN���Hk!�OȰ�,�<�����������&5����y����8�����d�|2y'm����+'�?'��{�0<�c~����7l��&�oO��sXu�q5��,�f�Ƴ��]�=�}�~���鄜d��b��N��ױ����N[$���a��C]�XI���
�}���q���o��g0ο���'�=��ui�g]?.��s�k�L��G��뵋�G����~���/���Ή[%���ܷ���9�C�r�����f�x�K��:�<bԙ�.�ʖ���]�K�ǜ���ɡ���
S�cV��xu��֎`�=d�*��)���ָ��*��Y�V�������'�wfu����9�
a2�pX*�l�O�?"�S y�:�s$�&�{����l�a���,��|�;�!�a3;�|�~CH6u���Ύw�:�=������{�~�?0�&��ZI����E�yܢ��Y:ɶO['�$�&���u��}�i�I���'�ϒy����&��߱�e>�㸎����u���3��l0�{�s0�O�i�ױ'P�&MO{<�P���E�u��'��c��q�5.1'Xa���	�5�	�hN��?p���W��3���s7�f�:��[��	P�?z���I���M$6� ~�q$�&f��fC̕z����3;E�v�c�~���~���>��c��y1�ܝ��g�޻�c�6�x��8ɖ!��C��&���d�B����?0�|{�Y6���y'̘E�3��J�8�#�$�r�M;a:��9̸���5Ǜ�3������w�1�aS)=�&�Cɬ�2|Ì��3�C�6�XVO&�9�2N!Y���CȲJ��d�,��
����!����*߽�o/;�:�{�����}��s��z;��d��OO���f�o=�:�0���I�d4���Hy����u��E������,�ɯc�M�!�w|����y��v�?o9ƽ�w�T�0�=߱�+wx+	�M���/�N�a2�̟��ba6��{i�a7�i�Y<�$��|�XGG�̑I��~�����?k^�x�Ks�����C��{!�N[!��6����,5�b`V�q��L g����M0�~̈́��2~�gY'�5�'����$�'U�o�7��}�_`��|�����I�&�:���'�����;�I�5���ߙv�Hm��(}�b��~}�N0�d�?$�gٲa�Mz�2O�z���R�}���2�N��T]g��V�s/l7�����-<�H+�V^��q��ˮ�x&8���AY;5Tmb���� ��A:eq'y�G�F
t2	�[����*'�XK<2�dz��漠��$�z�1.�. :87��u;�d\>�1��&�ѭcs{�3:��r�v��|��3��1,�/q1׽ݑ�wJi(�=���Qs�ǹf-�q<�EE��gu���_<�{5������éu��mΨS�Tۗ��wV�ܭ�����L����Df�˭��p'٦tY2����Guf��xIM[u����]n�|ű،���;��kD_M&�wT��4�
7�ue6K���ѱ9�x%���ѧkB�ܕ �w�����n�N��1Q��^]<=��HcĔ��& �˗�c�Юw�V� ��)��K��;�ΰ4moUݫ�gg1e-T:֋D��_n����d��ĺ�wݖ�!l��6�ŋ],$�st��*ݿɧ�+ܐ��ՖG{�zV����VC�=}w�b���|6��5ʤ�͏��n�_R�Zv<9)�g&�$mܰ��vbW&٫���%w����Z|��&f�������kY�	M��՚��ڰ�Cf;��pu'N��A߲�J�wLU�6լ\*�r��I���2�"��I*�5Z]���ۻ�;ri�h�=���C)&����r:�����X$=P^��n��q��vN���켇F��d�e��\��9u/����n����
��bp�Y�ۙ|�L���"N�� ��ݪe`PJ�(�	֩U��-�� `�WhF����p�I�y���-<sws�n���,��\u�\�*��r`�H:�>��j+��;Cp����f�흘��M�	�i�>F�e����F�|�s�]����q��]�r�V䳪�h�ΰ�NH�<�]�=�F��Q���{����ݓP0��J���������v��0�Ԁ��ԣ�ĸ���5ϐ�������v�u0،hFJb�F6TÉ�u'��&��� mX�sUp�O�wJ`������K�yd���T����DXy����E��CD�����4��2p��Z�зL2���X :��r�=�����4�)�Ѳ���W�b�����	�:��1h��GV�-�ۨ���a�T�@"��|�z^\��1S�L�)�� ���ZH�Çu�S����v-�/���lpٷ��j�+��/@���Y0r3m���L����X�&t�{d
�}z�����:��ۊ�e��5����4#Xi$�ț*X��4eM��C{�q�m�;��ռgYl�w�3�U{��<("��8�fHy�Hcd�٢g9�Y�I7�����u�2AM=��0į{5vWCձ����vYӸ�.3w�öő
5��,A�,F�J����J�UE!mD-��J�ci�\U�DjJ�+���XV��Ȣ���ªA+PUT�X��Ŋ��*L!(�ŅaV�[%�DTE-(����,UF"���EQ�*ֆm *1`����)�*��@PR��,D+X,"��"%FՂ�Z6�Q"�0�����FD�Qm���Z�b�E��&0�E��E��-���*��)U
�UTA���mKd��-a�X�1�
���������0�(T�EQ���iT[J�#���Ŵ�Tm��[E��UDAb�-*��LXFʢ1�ȵ
*#X*Z�F�)�E"*�d���,���`���iTX ��LY.(UQAAH�5*�)��QQ��X�*�k( V	Z0V#��Vڵ����mRT��(�Q��b1TDU�AD�."�l-m��+Z�PD���[J��k`*�Z�U""���U��cm#ҥ�����"���X���A[(�T��PTUTBҊ��b"ԔW�|G� ^�os�*o(�s[�\{w�rgJV1kOT���+9]�����4�\u��C�N����}L33�oh�������G��{=�>�I?�]��'Qd�o$������	�'��!�XN��=��6�	�w����2��Qa�$����M0�2�V����W���ۃ��us=\�~��x'�$�&�I�RM���u���ѝ�� u'Z���`y/l�:�~a����O�����~f���W_|�wP?��:�����G<t0��Ͼ�tY>g�C�b�Xe��:�$<��{�>I�Ry�'��u��`wt�@�ϙ��`y=�|��>��ޒ��V�c�>W3��o��O�vx��=AJ��u�Lj�G)�\ٸ�m���g�Y�{cuݲ-�/V�$���u_��R<_����U�w�9�fn�8n9�I��7�8ŧE�[��ue~Ἡ�窵T��@\��w��^�i��'��-//��3Ќ��ub��u�"y>�8x�٦,��`�{��rv�׎���k����\�y/�73�3Tصb�#I�d�}�-�vo	�qJy��Gb�:�i�/���P4�r�t��������ɫ��̝)�8A���[�*����V����r���\��j��kѭ���)�ݸo��<�v��[lkƬ��'C�R���:�Ǒ;_l����4pwT#�K�}9H����$9;m�Eѷ+"��+k&��rYIк�ۮ��%�5�e`�/&p���Wd�F_H�p��{{):�]����| ��g��`������%�
1���/GU�ɒ���\{���>��/|�����L�	���@��U�_�[��(��ka%V��`4�[�Ot���O���N�oě�q�y4��g̚�{Uc-�Y�����<]�JG����g��k���W���^�eu��"v����[�����;� r1w2�����_���ù{_�Q�sKq��Q�rn²���{W�N�n�/�'9e���8��#簡=g��W^ǹ���S�e��T�������W?�A�����d��M�o<u֥i�{��0�_��o�y�ȩ��7(|��P^�WWC��0��W��*VI�3wgd�ܘ-�^�"C��;����P���f��T��o����|{�_zdOC\�7�]ô��ι��ew��(U�'��(���X�rZ]�L���j��n+�9
tކ�Uu�f���i^���y­��i�f����u.}ŊV�Fg�ߛ"�8�f��������B�;N*D����6yL��"T3�t�а{�{F;�]Ī�qKY�Eí�@�W/�;�Oﾯ��ﾥx�~�����Y��"�T�5W�=���喾���IJ^�:3_g���3��5�{��|U{���6�����ٍOt����yO����2��?j��AC���]�F}%T"w�q��vV���ʧ�r�z�C�g��'S��)n��x'�y���=N���yJeh��W���������B�d�4s%��
�<�а][UԼ��{�5Q�����ft�k�sSj��Ӷ��I��jGQT=�uޱ��~�Y:'�8�)�����>��?y1R��[�`n��I8�p�4��/n��]R���V%�]8=Ull���üb�e�2�ːW����U�NІ:�]�m����}�{��{y]o#���X�hy}��(c垈�xj���%7�V��I�s�W��|�R-fW,X*M�o���A8p�W�1���ֆ��,ͿmwL���DQ�r����$��k��򈡪�Uu�T�f��לM=�\ק~ف����U?�8�
ձ���ڞqh�0�BV�� 	��F`��V��������U���$IsFlu�ݣ�z��F�����S�T_���ꪪ������f<��P�t�ޭ���;�x{&�x��p�i2{s�p�z"뭍��O������� z�N���>��Wͅ�v�Wz9�Oh�(#x��7ǣ�.�p����&L�Tg��v�|�j�zz��Վo�v����sړ�ԧGܩ��__Ly�qOݽ����N���}��mr�9���5�>r�ǝ��F.x������3W1,-��T�SRod6X�o�}e��������>��?qwE��2���v��T�>��bl3�m���x�������n����e�	~Y�һ��������V�_55�yVRqUVغ��'Z��:��~�s�t��j�`vO�\_d�}�pM���N��>���>����
�]�������姘~��:P<���8'r���/�"X�Y��K���P_���^9����:�@�O�ggd���N��ț��^�5LՂ��md%r=ï���3x��˷����@`=������v����<sk��纒��:�9	�r�o:*K�P�����R��69t��wn�]H�H�A�_@6u~���諭&q��ON�ο���N�����S^Y2{�n��.GQ��on���4Tݓ�=ó��?��Z�+.�q�}�5����}�U�����u�j������t�oEnw��'� �@Ul��O*����vm^���i����k�[�^��җ����&���.vr��oXj�'��fx��	������$���<����Z�{��⇛oW�MzV�N%��T��9w�4rȑ}�p�ḓNua�\�͌�70��R<�������cν��v��)��躆\�_��z��κ^l]?t�����M�Z�Bm����>��.�����QS��c����)Q�)]j�ʉ�����xK��x�b�:;>���P�-i�uNT�窇;�C۝kh�vlM�p�6uy�υ�e���&{o�)�^�/���w!���w:�|��y���*�����W��J ={[H�O���M�`���o�]Z��4���5*�*�P4�rq��s�1�oD�MVtd\̃|/�n	�Ή{a�hǷc�[��-1)+<���r��3Ԟ]ou�i��%	�9}N�R�����雟������[�x�^���4=~w|����=G��.�I0�2|��çيḷ�-\����~�O��j��y-M����:N#J���=� v���<�ʘ���!_\���)a�U�+NI�V�R��ȽX���~�+ݛ[堸:�"Ե�Ρ%+��;�}��m/r�U�uu䫷�6�+!�q{̬�ms�y�H�I��>��hy��|����ȝ+C�r���}X� �?o?e׺l��'HM���h·�2�?uV�xJ�I"�1b'�xo�����uo�Tʿ3��k����������_M%q�oRo�x���f-�+��Q�<��}��+9�-�&���s�RRS�r�h+�N�^�j��pq�����?m�Ë�Gz����?v��R�[<r+pc�$
^�69���zV�oY��n[�����l�x���7����&�T0gR�XA�c��c7���nݲTR�Y>�U��s��w���'�-*`�̞*�4�"��\7;�,��z�K�R��<�k3�g�1��H��~���s/Er�Q]�-�Yb��:�>��(�r5V�=,3�rǖ��+��W�_U}Vb�Z�[�L�e�ꮏ;+g=6�k
���Ղ�yԃk;��K{��=����/U\�<�S�ꑀ��{;���ʥ���|��W������<U����y6}O�dʑ�Fs���:�=;)�5�~w��8��4�[�o2�C�)�Lk磗c�7Oy<e�x;���<}�Ñ׽Ŀf�LK�=#��A�ӾE�y����c�6�,�#�뵎mݮ�b�7~�u�j�����j�G����ח��ϐמ-J�k�������9O��E��UGz2G��UKܸ���vsxfzt����ח�5���UVع*�u�]^�o�C7�U�,2�7I��3���p��t�d�o����?V��K���V��}~]I���}v!#X��;u�wB}'	Qn	���:��1A$�Z�V���x��y;<�7Ϫ��c��7oe3�[�T���"���{ � �YR�DF�'�tU��Yk���7�>�[ήu~}�L�]��G37���j�Աە��H52g
#��+���VE��M��{J*�� ��5���}�M�N����-Ju��`�I^:��@J�ŁHo:�Q��5bEL�2�K�����W�U^���E{�AZ��슬�<��I�7C��p�'bM�8�7��!�T�ZFŃ�=������QN�㻙B�Jo�}����#:��g��-�,�R��Z�	]=�^S����l��_�I��~��R��o��(���[�|���q�s�����p�5�X��}�s�Jӊ���z��F��1��>���[Ⱦ�9�Ny�7wo9��UN�ZX������_t�m�zs5Ҫ>�U~�'�s�=������!���X�ל�E����O2�M�m�v�j�;k͋��2H�3�e�q�/���dk͊{��w�`k��<7IIu�Tz�g���w�z��V�߷����W�r�z=���s���)ͪ�]W�o)�W�<�Q=�8�0v-1b�V��y�zel׋�̮</���k(?CGy־���q�N�����{vv&�x�N�j��xn�vr�Me,���q�QG�ul���f�e:�Nwwv�rr븬�۪�݌��i��8�\����ҍ'/z�k˓!o(⧇���Ӳ�<Ga}?}�}�}�qF��-����O<�Z����׾��O��E������V坔��E�3<p/\{��\Җ�S�eo���S�����8x�Þ�І;g ��9"+�dOg{jE��c�r�;��󖶱��p�5d����M�/�vm'�lz�}��+}"��jhOWt�w*A�\Rm�Gk��{-%�-"M�꼚w<��ͭM}�ewU�UO�갻��7ԯV�½M]������s�}:B����:��kj��[��\�20v͇�v�;�O��Z�;B�fZ�p�o��|_��:ʱ��[�E��\*G�=���O[�~���_lh����{�yM�[]룞M{|,F~Ҷ�os�xϡ��Ъ�:��Y���݇|�f���׽My9���q�4g{a/�OPxy�Y'Z��g�
������z�~�r��̶����>�M
O"7@���u�z]����#�z��L���3�k��A]�Օ����,n!l���k_ܪh���z�;�]�=5�l̡�8։��� �����gV1|)˦�z������;�|;r�'@��n��=�	�����着�{]���?��S]V�;S���'[e8;�l��rV	3�mG�qVR^��krN���{���j������ϥ�[k��Gk�og�=q�d��H)͎/��{ �=���O����ܦx�,hIF�ΰ��e�W���l0��8���Cm�d�f���w]N�ý��α�w�_�h��K�Gt��^�o���nmwv�7����B�~�+��>s��fOR�ɷ���OE���=�0{�`���VU�:K�ӟ\��7L��
��,{=Z�=�a�F�P�c<}°�<��t��G��(8�W�0��0y���x���vy��/�ʥs��0G��p?��"�\�w���҃��ʟe$����x����8�#���ǈ�аa����]g}��J�e�a=���{��2� F�+o�^oJ�&��=jG�u��ŕ�͂ZTl��>q[��tQ�r�AX��Î󃫣�]�f٬��q1>zsZJ�G���\V9�0RVc��|f�\%+rUA��u��|���'�pr���:�}�;��W�)����n�<kˍ-���j���1rS�c�����"]wv�[۶9�G�t��g�
#
��lAZ��4��j�{;��eWO:N|д f����I3"�ǻk����`��wf��cf$��o�5�ք�巔(ޘ_Su���m+O({�%Rx��U�b�7��6+�gs������uk�F�q�ם�4��D-�X�v͋����R�� ]wgE'b�H+	fvM��g��|�&Y�ʹ@�n_y���en�J�Z�O��wWڗ�_[��a����H��w҅h�C-vf7N��Mh������S1L��Y��}�;Kxܠg�������ې�]Y.�n&��f���\�!�[����X¶�v�GV�hw.b�$(�/;�M>�b�aV9�*d��.c��+q�Fq��������}ޏ}�}��t�xQ&_P%*�-�g��*:�n��Ij�����5�J[շ��f��8 �wK[����ө�`$�#*�����%�-eF;&N�:<��6;ˇ���M�+h�k�J�"���d�J�	I�X�8P��%]�S���۔����p�|��i��c�O(Җ�*��n�Z�kw��Bs�;#S�n�oc&���� ������/}]�fc.��b��N��\'�p3�93R�&#�.�̤,�#�l�k#=QtPM{�6�8C�d��:�]�M��g(|I�V�3�)ZP3�f��b�S:���U�>�&�b���]��A�t��9з�QJ��mD+�7�u�K�qQT��v�ڍo<�t���Vb5��6)et�4��0ey�Z2��{�,^.��޴�L���ô�s�-^`O��LAQ�fe�tp������>���:�cB��^yQ���-�:22T6�1����"���ϙ�]�O���5Ӹ��Ku�{�v�9��q(^��]��Z�1��\�(ݗ(./���N��*����el���]��f.��Ц#(�vsp�%;���q�]^����3������Um�,�:ɏ���.�JT�E��w4�U�	PV�P}|��R;�lS4�aB�\�4oz��w8�.��ZWy�HGCL u�bQ[R�9X�ڬ�ʊ^�'vpS���*,۬��S��f�����<k�v��"���	��<�Ԏ�V�V�$%��j5u�esM�y�u�n�Ρ/�a3����H����"���Z�U`�ɽ0^\U,7٪����(W��l�*���:D��r�3o3�^���/��QD�J�D*1m���aV�T`����m`��PRڤmiYhQb�Uk�L(*�E�������V��X�UekmX�Kj���ek��� ���AUH֫J�UEF#�**9�-)iUb(�F2��TYm+(�VV�-a*�T[h�ƥR�&�ֲ�V�4F--j*��F+m�QZ���jTilZ�il�bѭJ(�EU҈��DJ�m���
��,��Tb5(-�DAE���ڌ��TV�#-,���b�#Yb�-���ض�	Z-L��R�Zځ[�`EAW2�Q�-X(�ŊKh�QFDQ�..WYmb��)l�
6��EQU����V
�TF1�������,KaV1EJ�Սh�PQc���b�-���AD`�
,V�D@Y�Fڳ�"��Uc�*��F(�T�`B�lm�*
*�,����2*(���Q�)hZ�����Y[�X1U�R*��#A,UT���m�`��J�0
�$��Ar���M9q�[�7j�'�\ʖ�p�LT�8�,�F�q輨 ��bt���S��WI/(E>��Rg7E�o�_�}�U}_̗1F�o��&��o{�2�Υ��7�=O�n�K�q�ǽy!q��t�%A����/S�������Ֆ�o�A�zd�I�5;3/�w���{X��\siz�/l���ɪ�œ�]�W�㼜+�y�uǓ���9{��{t��Ó�I"����%�W�jM�ԲC�|8��n�ћ�&�`�^˞���}�f�睕7:]�J^E����o����}��ԜVͬ0��<��}[�3���R>�<z�vW:�����w2�W(��yA�ի���/^ԭ��M���y3�Tc�ʦwJ��+��u���t�b������3��ʇK����;uǜ]J䪴�Ҩ$ U��\�Ƽ5�O܍n{�N���(#�zT;�\�VnE�����I�\G=T�9�["ʵ�/���0Y��@�\���_f�j{��N��1{�g�]]>O���35�8	Wa�ٙ�a�:{����f3ۙ�ކ��%�z|X�� �]C/1:v|5c:E�-PS�].�^䕳:���w�#-=���e���7S|SW�S��u�T��L�F�A:>��mtݽ)�b7���>#/��sY��:y>7{��l���	'��<�e9��N�U�}_W�sj9��9��}��sU�����hC���rE̝�&y{�}$��yg�;X�o�'�]�>�9_p�K�{��/g�n�;`8�6�3�8��^31���g���*�yg��WP�Z��x��K�|^7x�>��h��ƍr�����'	���h��Cݻ-f˘=[A�W|<�&�vX��9Y��?���p�I�ɸcT0ӏׯn/wnY�󻜮/�5�	�'���_](�����R�D��
�vt�W+�I���ªh�`7�����'�����<��ʘ��S�5�=� �Nq@��2P�u*7=`N��쩃�@Y���x�I�:�(,ѷ�>٨*g7�U�a[�G�]9��3/c��:�n�����x�����w������pw���m�^�H��O?�fݲk_:��w_���0�e��I̻=�L[��cK���d���n���%�2�ýI���v��ג�Tw2�V�����D�*�9�H��q�J��W4J��Y�놷���Ⱥ~������"O��������;��b��T�k;���ɀN�)rX;�<^���Y^Xg�W�g����Q�/�u���o'×ޘ���ɾ��6ކ|��C&�v�����J~f��w��޿��jof��F�Zz�1���cz]�I����)jo%U$�8p����:�?��oZ��zd��']�;�E�>���/_*}=�&��}I�T�_���h%�2{X̥Q�ӷmpܔ��x�z�'���p�X嚿��IO*�RJ�ٯ7`w緘�!�;��I��%Wӂw19~��]��ă�8�Y�XS��>^������}��d����ċ�-ܩ[6�u~�}q-zyuO�{@_S��uq}Թ����my5��Q�K��yO.�$
��p9S�8;�1�#��?��k�q�/>���-=ͨ�Z4얻�yѫ�$��<i��Vy���J�J�w�w�N��3�w����{��a�ՙ���&]W^k����(�C���[}OzP�@�����y���v�����5��s��6���ʱ����I�6�̋;t��с���]G�U}_}_Qo�q{�,3�y�Qq�מ�;�Tc2ӌx9g�P
���z��oK/t{�z��½�Jȏz����*��c�W�2��q�Zͻ����O�v���y�W�����y��Zp�����I^��g;��56$�M��/��֌�G�U����Xg^b��etqcw��R�Z�z�gyP�ێ,w�M�t�J�T}xΟ|��ӝ���>�<�����^�>=��2.���kRN�G�T�Q���%U���z�Ul���a'� ��-j�zd��]qT�|�z��_��3]����y�iEB��[57��[�7}�I�_=�=���{��g#�]3N��7�='���\f�'����|�&�^�_�Uڟ��O9Z���B��[�m'GZw/�sc�|UzzHs���ڛ�&j���:.��V{��#�-F��������N?ܽM+��Wdˣ�H�嵀>����j�����q�	�8�Y��h��iL&��z��\�oW��Z����n��/B�[e������VF���eX�ъ���R�{�����M��˸j��}U��A�ߵ��9��};����h��h.�P	N�^I��ד�����^OLU{�����s𯜘� �! }CFw�]U�����\nb�͠�<��΃$�rT[��O#A�'��U��������9�y�wvdex��sSj����"���]H�'-��z,� #��]E
��P��'��'�����eMZ,/�b�m��ڥ(�K��J�H�Aʎύ��� ���W�7z2�Z`�w!-�x�ٲ�s�_���k<�`��u/�!EF�A������-�w�#�	�}��ǥg`X
�}��g���_ɘ_׎�{+�X3��9=�:�����4ZI�^�|�!����*S��ә�ʴ�f��n��?dP�H��3�ֽ���W��F���_{�S�
k^�6�M��Q���1���ԥZ�H;�={K�w��Q[{�;�]%�
f��(��-��0�ө�Vٯv�~�Y�2�g{�ۧ����i$�}*�3V�����2ٷ[r|��m��g���qQM��;�P���6vsU&�v�U���a�rcY>Θ�/5̛Gm�rj)� �1���;]�U�\xO�H�i�2�]T�y��Wӧd0:mV�,����/^���;�ش���ki��V�,�I��{�ҡ��}�꽕0�5�s�4>�����_}_']���ާF�`A�2F~[�=Ədx"�y;=�[�ЏH�(J�����sM�{����c�mmw�����e]���Wq�XC:sp��3��c��Y�������;�z����ﺋwj���^��,�����R���o��yN>��lxS�{2��������yc|�w�b���ڙ�D���ci}�����z��z�(s�皃{SҊ	��3��$�LgA%���v�\�e�+�(�6�Ɖ��'G�yWc���4��i26�_n̢�Z�dWղ�;�U�P�.�p|+�ib�E
��-CC��O��'�_A*9�qӿ;Y�o_�nt�q�����./�%�J�<"\UX�sS|�#j�RPub��Nٶ�_���6T�>+J"5�0n(p�{v���D��
��`.sF�R�r4�"_-7^�0Z{��dʽ������b
"���J��̙�C���7�|�W��6�l`_�����1y`�r�7Q�/��虬Wq��-��7�0y��P���ɐ럶�����7(�93PSS�[<Q�U���z�E2�yq������E�=��еX����CtU� $��u�t�;Y=�&�)w��)nH��"f,=�ݿ\8���7V��ܻ}U_}�3��1MOO���m��8�f�79m����Q}�p��C/*�"�u�Nx���J���ـDq��鈶'��}7���P�t`��tau�h5k!린0�=�tZ??_�z��k�ٽ��#�B��c��x��,����}
o/i�>�y�h����=�*g�=s�����wJ-�tI�d����ᄜy^=�3�ps���-.����,��Mn�x��k��fVJ0��Mm+6��O��q.�8bU<řbJ�/�=p����ލNQ.y�[�Q�P�${�6��0�F��h5�F�ᬲXU^��r�cσ�=<�t[���Kwt�����|��`�D��Ӷ|:�dx������i�t��dV�����{�a~3X�6z<�*{y`�=/��\UzQ�h-,$�����5*}}�ݘ�w�s�� o�ʜ3�_���z�'8��q���p���bP�Bc7|�qq�P���1js����0_�Q��ų�Қ���4p�9ڧ����N��MS$ʿh�ϴ]E��ʕMl�=���7W��me�E��a|'�	�q;(��6�_`��g��6�X]W��X��lh�iǙ�][�I��eɻa�L��I�frUx���.ԇp�*��nr����}����U�2���گjX;rۮ|��|7��"�t�a��y'���q8��?,*���2��J����axJ�f�<����>�)n�zE��Bjҗ�X���_=j*
_Y��_x�(e&�]pp9��~`2{h��zY���W�pm��� .;�P|	�ט�����V<�!@g��jm�B&)��[o�����g"�>�k����],;0֊xzڂ�m��;�f�y�f�׽�_dY�jO%Lew^�u�j�+��X��	�7[6�E���Z�]�ms��+�Ȼ�{�o,�Rs���/o��Lv="��	���U�Z�M�	�H���gw�N�,����f�e��<+��`�u;���S�s�1	=�s�/�:�zk��	�d ��٘�7pt�Η0z�Re8��pS�Z+���yu��]pC��|1L���7n��_��ޙ5C�[\%�Ɓ��B�U6שW�A�pp�,��5�o�/>�A��fya��2c.-*��9%�N�R�����j�a���oVS�W��&��؋�����s҂�{���N�ӒpT^��UɱM�`N������]�D��\Q�,�YX�N��t�tk��9�z�X��|2+��y�+$�-�ͮZ�c�s����&\��N�*��Y�{j;A���Z3X1�,�W��UW�c�yΞ����ځU=��ۦ ���!�ou;���،�ƾ��k�8�����Oe����]��"�U<���jm�����M��a0Q��*����lp|�\��V�����j�,�����P`�k!��U����lO�SG�r5����Zn��O�ai8���{l��kc��f^�NQweYj��d�9�~����z��\�N���^ލ�o+�a���q}'�NG�R�{,p����z��W���*��L�h�w�Jzl�衊�hr�SN7dQ�7���U��26�$:���<{٪C^k�z���>�|'��`�#y\qڂ�[[C(8tY_'�V�F��qf =�t��/��mb>�^���ڼf��"�O���2:��u�:���j.�߂��Mw'5۸�Lx�������µ�Z�XX�1����ϞV@���N&ߒ���R����X�]�p3��G��<=B���U,�@�s�z�<<�p��P����јqJ����ۘR�#t%���P<��B5���Ĭj��y��ǥI�@�=v3�!�6ƾWy/�ob	�Ɍ\�v���-�9�϶�[�]9ܫXJ��s/���x\9��tk;��s�[��˙P���f@h�z�&V���6�wi_�����N׀v�얏�~���U���R��v$oE�^!�W�bP�㇁�^�b��]�Xx���j:�wS�PX��ǖ_y`��1
Z~1�f
�ĺ����V�����-�6�	�9�U9�
�s�s��r�C����WW$\��s�Ҳ̰�j��~��Lq�#֧�!��T0ۓfi��r9�}TN�(2�����B�wγo'��؀7��=kt�}�h̏>�q��y��b>#��
��X�������w���9R����+�*ȓN���2��#3稉n掼L��V��!����ݎ����|KqCa��|�8��)��I�R�1�o���r+�;q-��]��"����m���XO'��:�a���ȡAۘ }��7=Ľ�R�k�ױ`���*;B�\0Q�BB'�>�D�Q�Ԍ=Է^��5���F�>��9�&S.׍9�n^�����00:N��
�HbP�CJG�+i�u�G�v&���3 Ma�2���b�Q�e]���Ђ�AҎ���3`'IfWU�α�7P*��`����s���V˫�����6T컦�#',�ǋ�����M泜����njGS��\���]�:����;o=���=r^e��3)�ȣbv�*����r���Y�:rnqs�|�+H(�Y����Jk<�gg>Y��5�@]�� �_L`^&�TY|\+2W�:����t0S����Z�Dfց;�����7JY��v9nK��5}�8
2���>1�1k�}_t�[�Wd�h��S09�p�ku֋5:�;cG$ �.�,�i鱞통[�pv����%�z���(�u|i��F>̇���v�Z�m�
�ns5eq|/Uvi�3�JN�[n��u����o�n ���A�3C���<SGi�������u;!��X���0��؝q۳��,h���U�r.O7���S�TT6����Y��ErtG-��)�خ�\��J{��zqu=�b�w��ڷ�}ә��e.��Tm�e�+�ɍ�Vxi,M��8����ߓ��D��	[R3ig#X����7�fx���-�����v�R^as5f>l���N�2���]Ġ�4���㽰����-/�Z���F��t�R�㽭�c�Oq�cfm�e����=�R��P 8N5/k"�����Eo�+ED����ڦ��x�Rl�r�f�Z]\�o8�݋1�,-Z�[�fK�Or `H�[)7@�&uŬU	ft��uC|F�u�*� 4Ś����Ҏ�Odux;���ޞp�L)�
�PJ��v�Ƀ65�ث$#�u �y�qz�:i-�����m}�pWVQB;�v��g�Έ�+��Ku�u��d����][�ܥ�̙҄�NW�[�^�eK��R�}'I9ٮ�,�lU�wo�2�V�LA�J�YN�ժ�ib����ntˉ���{(ïi嘖�-{z��
I�d��G�.Gh��V��]�ڤ�]e,��g�Bi�Y�!�f{��.��h���l�i�ګtB�Y��gK�m0	�YK560�)�)"���:�w�r�Kr,�*��/XX<���w!�(�L�eFc�
��VG c�dA6�������S/&�ӫ�����{Eպ[}��X⼈����O3����e��][���ix��K�a1�I�-[�i�-b��3�����Ӧ>�˲�UvD�[״�t ���5�@N�y�s������wi΢��՛��v�9�08���W�*�fV�~��JM��GN���]o�N�z�_&0+x�r���tƺ�p]����B�}�QlIb�9W�R\�����r�S�M�q���	� ,�u�����=�к#�;E��֪u��=c���(�Q���P�˶h�
��0h�+� �Ȓ��:Q�JO�5��Z2펽�B��'d?9,t�\�;�U�Ė�y����9��FN2�-�U��QW�D`��sl��kUQkD��TKKm�b#TEb"��[�T��l�a���V"")��#�V��DX#��B��U���X�F(�EEV�p�b
#��#��(1b*��9�E�ZiDTE�+ADb�QG�EAEDTiQH���ŋ*(�VA�%H�b9h���APU+EZ���F""�3h�-�Y�Eb�e�Aa�U�kQE��Eb(����2
娂�űc ����si�mJ���a��!�V"��b�U"ň��-Eb�Ų�TUr��X���E���-*�"
"���b��lEAZ������(,Q�*1F1UbJجE�QLEPUQpш&u�ޭ�ܷ4����\�E�^��5��0���n��r��I3�?_P��YˣwԞp�H�k��~ %���������o��;nos�K�}I.zpYK�c��l�9+���G>�z���i�M@G�o�k��B������zos���hW�m�(�גgc����PpБҩ��z�ȁ������U֤һh�*	�P}V�tV�N�Ӵ�mj��Z0H}U�h:�h	�;@-o{���(:�{S V<vʯ�4S�w��gW��W��d������`ʸP�Ʒ��\�ޗ������-i���`*r �7�"�x�.��"�H��xI�T|,��o�'���;�e,9˰s�=Rfg�yo�Mzp��'����<{k�A���v�@\+c[aZ��Qݐ���y�9+E� 4���9𮱑\\p���ygn֝���G3��{[��7\9�Ђ�W�!�6�`�t6R|����i��c�s���۶X��wJ��5�GݷY+���q��X�8���\|O:��	�i�"bT���0xÙ��ݦ3�Q�#$[Uʷ>�J�P���^�W����\o�G�c�<*ˁ�P�@m���
�~��46�u��t[]^���YY�tʼ���[c�i��h.G��׳�Ճr��u\C��}-&55���Ј`��ԇwL�HS�G�< �*ܖhrA�w��U�;���`�it��WNSk�ݜ
a�� �u������yV=闅�zTZ�x0~r�'�ܡ�Ϛ���T��~B����jZ���5_��{ZZ�	���z.n}:�!�3�xrI\\�U�W�a�P�| |�'-m-��M��;�m�Z��C�uu���T��3lIxО�U'#���8Qc'��@��Iz�3S*-�8�����ɕ~�8/�F\y:Hȹ�G��]��Ъ�J=l��;y�J�)�,ʀzJ�{�P�t[>�/�`?���X%�]�����1<�殯�h�}��ۻ�2�>!�6������E@*���y]f��hz��t���|�<�ѺQ}�u�p�Ӏ�!���_>ץVҘk�[��ʕ�sƱ�n��C��S�ڼŻ�r���fS�D��6=�J��_�U(	�ч4S���9��ɹ���n:�~�w�6�^��~%	�ͫ�0[cMo�ڃ7���Y��*�U�r���x��tV2�����%�w���/AO�ʇ�pW��A}�0�Oݦ���j�gE���s�!�5ev;��s��B�����txP��%���d��HײQ��ff.�Z
�]�T�4os0b�B�8k��@%�
!c��V�]}��h>�U�J�S�n���e�Z�=��S�8�mc��c,VNX�ǔ�ؕa|/������}����O�{�V��Q�T���A���������%z�� 6xM��������f,�oaԼ�=F�����ڿW
3��X׈�VF5Qx����%`W�A
�4��Z�/}r</�ɏz���\pM���X�4�ʡ��^�W*��oo�]��|�«
-?r@+o�.���zn��Ͻ$�5�=N#ł
�F����Goux�=M�ުu�|;��_y��ld��*��*}.������Xʊ�е�3|A^����V]{k;w��8#c��G�|X�:���h���>�\���!K�jE��a�,޽u3�Ӳ�fX^�����n�(`�T�C骸X��qٮ2�q�!�ԛz��}
�g�ei��k�T3�bpZqs������[J�jޅ�~��ߺn�w�)b�#>�+w��W�|�Az!�I��ϊ��M��M���k�B�`�+�ˍ^��U$��=��n-"SLX��/E�MPb0���p��O�6x�:i)ej���V��꼳@�L��C��C�,{���mv�{	�E%�
��g���Z�	WL˧o���[CS�mK���w��)Nxѡk�����Mi,��B�׶�����N�ԡչ/>�c����5���2qABIZ�_ﾪ����'{�nG��M~�N�9^������v����L�tYM@o�h#K�cGDp�g���ڶ2it�cK̕�!Elz�ڇ)��i7T��L��d��YUl@@O�'��g=�����[E
�^G���ǉ��%n������R.�o}���-�ޥ�fn�<X���)%���г�u�/�Y���P�:<-x��{kՏ��2�.�C�5Csy��.���P�ǙN9���EsT�⸲��`]������p���ι�>�5)I̓���'p{=j�_�|�/�Q�s�3>�=>�S����3���µ��'��ROHz�����J��^�>���9��ׅd�[�{�.�|6����Ȫ�þL��A7gg���A a��Ю�pf�n& �|�D��OF1Ի:�s4���(\�[+��v�zZ���0���B�$m�|��&\����B������|}��uŦ���Kسͻ�*�NULj�i˖���mdI�%��`a�-ӑ�ۺ���C���pݏ��e�iI1�a�u�w�<�3_Q{�+��U�`�,ʶ��ݘ���)��ie���C������\�[og#ϸ:K.�^�ղ����$�l��Es
�:�\�����8t�tj��ɡ]a�����q�?�UTb^j��r]��=�P�q�|dQ��h��{�����%�;�3�zl�~�fJ��s��fLj�J�8iKnȓڻ�Fn�u��Z�T���}_��]�~���'Ǭ�Ofn��^�f}^y�s�^���pf��~�B��D��,x  �_�q�o��,������Շ�s*�&S�^5�"\�c��(�*��o�V���3�ו^w�.���Ph��Ph�խ�%>u������BWk�&%wn;!��xF�F��lO�(Ǣ��
��-(�|�� �P��/ֻ6�(i����TYK{D�p
�q��Y���X49a�Utq%��s��)ih�1�U<s�1�sv�I �~�z����nN��z��c�H�ūU9��xОj�X,�(z��)�����e��S�~Q�,xX���_lO��xi.Au���=�~�,*�^�~�~����o{�K7j%�kәY �C����Z�ǜ���a��]i�����1a���p�L�&f�ד9��>�c.�$�jx��*���:�pʹ������C}��$��7��]z�Fٜ���蕍ׇ�A���v9V�t�V�}�������U�(f���,�iM�k� �����ndt��h��������n�T��N�w����ؗM���_�Yb�a���a��<zz\FEs����{kڰv���W����|�����m��h�:�aV�FO%������(*�� ��ό�6`�UOf\��C*��o��F�;u>�,kV%���"�PkԮ,�tUc��q�%�|`��u�	٦��5����ߪ��߇�6��YO**즩W��\��Fx��Դ9ˉ�ϸ�˘�ѫo۽��^��\�#��c�.���xFPc��!�iQwYC����3�R.lۉ�����;��ˉ�켇�<��D{��y�T�.x�+# Ã�����7w�;Y��G6��{�W  �����vS���:�CZ�Yf��V#��Z}�P�%�6KNn�ɻ��� �|J�b���L<,c>�ArVL������Hj�hS���̹z�Ms�����}cR�'� ^I���J�F�u�����Rcov{e���MD�����-��q�+�ߨ�R�@�.����XT��)K�k5S��2$gv�Ô9r����v;�B���v&!�o%N�^��.�R���4Wc�WV��($@ux��4

Y��n_-��*v_!	r��<91em&.K�i�C�Wp�ܹ]���LO>e���]�VD�u�(Ĭogdś��Hמ:����sw+k.�V���>���P�뀫��0�d����t%��ߘ�y�ꒃ�t�{bCsar�}ؓ��Vʛa��2�U.���bS��ׄ�`.�Fx����k�A\�>�=�y�eN��,f���ln�Z�����)��/%}�Ǘp'd�+3�����^oq��})��,����3�(����d�ǅJ�j������� I}֯k��you�L�r:葒�D]
�1/{�h��C<`��Z� �	��6�SL������'����t�b���[.�w��b颭��\��1RV��)�9����Q��#{%�<�Ӛ�^�n�w��g�k�q�6W��,V��
x�xJGY�YDڋ�E�צK���m�{w�e�:d���C�._��vn����Ƥ���/z�Bߴ�N�����{�Ӟk�8*C�*	��4�OE��g ��TR�t�kx��LB+���v�ı|5���4�_�<V�_���U[��1������+���=-����T���N$0?V��4<�5��)4�6nXXκ=/���"�r���.���Y�ˬ
z^��\�Q� �\m��uk��ȟh��>x�S���<��\�9���{S�5&�J�b�oMotm�=���8ie��]�(�yU�(9m;.�3�?}ZraO��w��D��z%*;A,� X�c*Ձ��F*wPxk�V0�V�e�W�7����S�} ���j����������Z��<�z�'��s�&c�]��2��}��/t9/�ޕ~W\��b���%p~H0j�r��P��Efv����Y"4�Z��$s�F�O�%�q���,�á~,W���dtG����;Gp�׮�to�3ȸ�5���P�!��,j��(tGU�l�^->�V|��m�V�z�"o_B,�pW67�uR|Yơ�#����i
�t�����xN/Ū�_b�K{K5�GՋy�hD��|J(STk��&����u�Ǳ�S>�j{!�Ӆ�zs<a�ի��Y�D���YʞaS��4�t-�T9���C�6/|o����`����싥��Ω}*i;�d�ܷ�^�y�_��AU�9���X/���a3"�Ѭ�0�Iߴ⋽�駼�Љ�@�c�؞ɪ�0oZ�fo����!@�'�3���r�<�k!Y��ٛ���ڭ*%���\w%�to/�]��Sw�;_a/�F:�䖹��{��5���q/z.�L�gf�4�4���0��1w!���s�+O�W���l}�����v/�bD��ꔄvi�g<y�Ξ }����Lu�"s'=^��D�
T/���-��O�gêG3E{v�ⲹ�cs��ãm����ظs1뉼���V׋��P�B�7B��E��-�����dثo&�5��#y{}��gzt����*ĵ3c�zx�����#�[^�=/б�<����7�'�߱����7;��f�i�]�-�8/�ޞ6#|i��m�1gM�}jn��Y
�j<��W����gڰ��Nj|��Ϛ�q��-����_Uq�����J�-�R�)��S�ʍ���<V�/��<��h!R��Vϕ5G�F��@p�f��%�����dҼ`_�����T���Ix�	�P���,Z��J ������c74���I�ݍ@�pvg��gf��Z�W�(q�#u�_��]�*�K�+/(^����O��ݰ��N�ﮈh��2�UX����J�L�'����)BEF��wb΄��8�߶^���p![��ϩ��3*�[��^���GQy܂0e���'��g�P�D�Z�1&�M.����.Y����`wu���{`s�kUt@��:eN�Y��,`�׀@�L�C�C'3^tv�y�=2t}��ٽZ�;�1���\�ӼN,�\�[��'���Hb��v���k�p�r�t2ĸ����7H]M����Dś$�����n�AWt�|ʱ�$��U��_(���g�[O�(A��n�[�q�f��ޤ}�{�3�{C�N� aК%��b��Q��=S)�]{�ӵ^�U�"5��v��SO��x���:�s@E�<62J�]`�U������|�ԟ�]��$�iT��$��?��	��~��i�LV�jR����+�U�qvpmM�|#͟���.Ƿ=3�)S�-ٯ��]s�Y�\�^��"�FyJU�4�>�W�����Syob����er���98��#���*�vӈ���!�:��_]J�ߔ$�oܹ,���.�z�&0�sU�:��t��V'�Ƶu���"�S^�q`�to�����pĢz��j{�λ��A�|��ˬ)D̷=p�1��C�F�KCo�P�@�j�G�e����������z���ʤxJ�ס�ҌO�]��Yr�`��3RF�t/��E�qG$�_�<�Om�2��5ߡ�s�O=�8�T�`���7ꮇ'��o6�
v��Q�4�.��^��{$ل-H�4�i-�XҪK�H��Y�����v*[���v����ߺ-�W��o-Ћ�:��9G�TB�ȱ �biw�k �{eMB���cP������n�8���uu��3��ٛ�ǼJEv�L�B�>�3V�$�2\a�|P�n<{�G�f���.�6`T���X�p�߻8�bS�c)n]������B���֧��5d�no�Ӟ:Y��st�AX���[��ƨ��w�)0��f�:{��";Ŧ������핌�9�����\F��t�`���� 򾮺� "QcI֦WA���9�@�W�Ju���O�&(��v՘�<���V��˫+T��}8�
d�H=o��\dY��}Ȳ�:�Q�u��Ȋ�OQ�=��d�����W�-�P 6m�B�:��%{�㩹w ⻔5�&�BWd���[1�u���c��u�#X��$��u'Q�90Bٰm� ���k�q���:����g9���i���"��/T�J�M˴�L�5w<UY���U���]r���oH�����f�3F�C�V_\�oRtķY�Y�f��}+�V�mp���6k��c^Jhe�v%�w����ќ�BNԧS��;Bޗ��j�o/�k�U ��pv�B�]����XUn鹵g��5��!^`��I�nW&e���[�w!�:Vd��p]�Yl�p�Ĭ-�/1n�9$x*���Z����:л�˽z�O(�0Q���;�δ���m[*�. ]e����'a�E�̕��"$}tnN��8�~�h���ٸp�w-�R��l4.��9��$l6��CR�1�U5�+0��o��em�m*Ru��l|�.;�b��p�Ne�c���r�Z�eg)�#�[Qq.���w��k��X��[ݒ��i�Φ�pWTO�S����1fil�E�2�jusxB��;��tSћ�b��l9m�,m)�'UܣX��v��c�u�aRD��C���E��Tŀ][�W0�tx�>��ۮn:'�0wZ�lsw�;����|��˵6���{��͂,5З%�u�j����4&�
j�'�2�XӫJ�/r%^^�OD@I>ߦۣ��|-�܀(rv�ά_j����;ۜȫjq�E����5O�8��Y��j���X}$�o�o�s-��[��n���}�i˛��]G�L+���P7Gq��2��ƻ:T+D�����]Z�r����W���Exڑ>�	�O52�#�3���[y�{DȦI��p	=����sGY�&ٔ!z!�]P:}4Ջ(�v��Y87On��n*��mՔ�}B�������H��ΜE�B��p3�"��n���6�`V�!�C�0���6Ni��v�����7����P=���y`Tŷyw�H؟mNސ[����d�Z_gJ=��{|)�IM4}gcn��ug�2��u;n�Z|�o^�E�e�� ��o��_J���@AX���E�(�,`�")RUr� (�H�,Q`��$��QUQTH�UX�U��0U��U�1(�Z��DQb���X*
�QXUH��-�TF)�-*�V*�*�EX���b*���X�EPX��J���\0�#Y��V0DX�(�(�*(�����*��J�,X��UQ��PU0�(��,TYZ1
e`[dUȠ�-
�EETb�b�0����mQŪ�EH�`�Ub��Q�A�4K�����X֭J�(��ՌKKZ�+aE]��V�DP4 [���q����"�uܫioi�A�;g[p5{A�QI6�䶢�}�#��j��uY5a�f��/�%��_����$��|��E ?�=B&!R��{�ڽS�c݂U���Q��l+��ɁQcy���7=��t[����-�p[���¡��3�vr��]��~a0�!b�1��'�9e�ZQ.�^��ĩC�����@@�'���M�i�;K"��R��y�^�^���l���/�?h���0Q�Ϝ*��X�C�\^��K�c��u=�	��n������J,%�8�Pq=>�Ě�*�|	z������KL���=��W����/{��Z��3�������K�B-��O_�Q�F �)eg���s�����ʾ^傳x_�J}o��OƳ-�𕺲^�B�JV�q�+���yK±�.)rl6A���^��=J�6�̮>62�C{@�w���0sfNuY3û�`k.���uY���f��wV�I�z�E⮺�0�̕�`e>��.�Xa&��&,��[*���u�����V=5�k����[όC&�M`��\��:����|
;��Y�˲���Q���b������o�ud][+�-�"���ǔ�����a�mսEn�tF��%69Ӥ�W���r�e�W�Ҡ�{Qh�
�`�2���ԭ�]c�L�>޹37�������rL]�g�틓�;(Z+z��L?�����ﾆ�����a������ڂR���:���Wbӂl�eg� u�P~��g��k��5�T=�_Oe��/;�������ˋExtmr/d\�}2���.^9hwux!y-����`y�B���=
C:�*��&8x�_���wѝ�����U��P{������e�y����u�БZ.���|f;zHk��7PNw�磵�`�Ef$�.=س,��j�䫼v����N�C�؁V4�"�����wPxw��f]�5:#��B=3��S/�����ʖ�8�;�1���,.~<����tf��c]����1�qx3�����᯾�����~�B����b�����f�Ө1����<׸�H�Lf�i��L��x�,!�1H�]eL��4EKv<@�q��kso.rOo=�NSvuǼ���ysf����V:,-9P�3�kS�3޾��8�sw�x肐��Ij��E��&3�u-C�>��&�J�GHK�.���t
?W$twix�߼M3AM���dǷN�1NeV��mlر��(mn�oTu�F��C��Ʃ���d2��䨪WB��Ry���]��J�o+:�c�>�}�_nT�Ae��sh^E��<ek�iuE)b�:�G�;��&��(N��q�^q]��*]{������f�m�gy���K�ˬ=��xV3v��S-�Dg��e��\�v]Ӄ�}��|�;}n�N��9��A�����X�T&��3
����C����o��㸬{�n�h!��\٬�����Ђ�W�|ɞ��Y�o��^�<�)��}J��+� ��.����{Tk�ޚ�[O#ר�׭�>^��a���7�Uxht�~³���a}{�!y��jO��5	�3rN��k\x��U����>�/ja�k�3�'5�S}~�[Η']H���M�s%�ootNƜ���J�%X�W�B�y�J���C�bV���Eǹ
7�3,�%K΁��4/s���o��V��ޢ��jb�%��z��\d������Q\Z"a;�G
�m��]�2�b\�a)���q�*\�(�o*[g&.�Z8?��|%x�=��`|<w��g���j�$L]�ҷ�oo�vrsS�.|�	�q�Aa.��6��U�&���h��5��t�wx�|0R��ߏ>�Û�����B�̮/J����R�����)�q�}->=p6H��oJ���ψ7�}>����9M+ ��m]�j�q�=/5�-���:���dR�ѥŒ0��J�j-Wc����5�@��v�-%r��7D9;^�����8�1@kI�}��j��뵂W~��-�j���g�p�Q`c8�SQ�N�j�j�r�H�AC
y(��k%\��vլSu�-��+q�5�}`���T;7$;��s>y2�ʗkƜ�n������k:v�x�0`��>a��>�b���]c�J+��%�&�n��W+���(����0{���"� આ�|��ޔC��֩xz�*G6�|�E�W`��u˝)� �����k������K�~��?fKL��C>ק�����9�(W�i_�V�/e�>����4�K�K����Q�`��T_;o����IC,�y�eϷ���:�j��#�:��\�e�ll<4�U�7��,.�E�(}�Bo���W?ur�7毋��Y>��?��ڿU��a��l���j�Z��gF;l	g]l��fou;%b�GS4��Q��}P�ج�,_��[������԰�ތ�P{�Yk�w��֙'.�Q}��:��,X'�����:2���?��Z��;B�v����;�9e䭧�^>18L�X��Y��X=���1�,�ͬ�Hd@ ���%ϲ��n�����.��l�*fB>��]]�eI�C���@p�(�vM�ܪ�����{�-�~�^�_]�ʤt��Nɺ��y{5,)�iܧFW;�UU^��g{�,�޿V��g��}�V�j��*��Y�g���ê�KC�������n��t�O�珚L�u��i�����r8r�P�P��0��sV
>�c�S84Y��{z��><N�3�ʜ.6'�a;��}\��LrT \v�Huj�}���V<q�/uzt`:��������\}�y�N�	K�^3�R�b�e0i�n�	!Uۣ_y��WzvW Y��_�?I�bևr�óˮ:=k�e�ک�V"3١W�#�̯NV�������{�p�u,?Vb�Tj�&+�ʭ�Ç�Ϙ��"�}���Q�UaR�0�eRj��>P�@�'���=7e5�dQv����b�vprf��5Uӽ%��9<�@%K�`)��p� 8U|�:(0:��վ�x���r7�R�^O�܍_�Dj�9����U��R��q�Cd�|�Ė�Ĉ�1�{1)A��qh}���jnY�\��/��Ecu�f>�`��N��|�NF/E�AK���� W`񳠾Ҟ/2}��;�`z�-aӣf�q�����֨+mk�G�_TNoP�s�<�*�RP�\8U�PZ�B��gUT@����0u逮krY�5�e�B�r�|�����^)/qږ�ܐ&ps�]i��b�-.�*�c�jIӡI�.?�����V��}����
|e�g7.��i;z��N�a�*�Tӄ�G�o�^����|c�_�5|^����~�Y��eq��9jõ�]g:���[�iX	�\���s<��wW��bÔ��4r���E�E�o>ǒ�p5�ߔ0bSu��K|}j�\ض��������<��?d��Wz�Rt2ֵ�+��F4�IZnH�_����Y�;Js{g`��x2e-�>�3Gɍ��֞ex��a�P�+���7�Ȃ��Fyn�om�m�> �ԫv�����G�������E�e��p�ci��W�����������s���V�Ti�d(mgW%_=ǧ��b9����}���#�d���M���u�ҏNoL�m���o���]��yL�W{
�$����+eb�����^�2$�F��~�4Qw��[c�cj�+�2]��׺�x�������+����ꆥ!��5C'�upz��%k�7`�Y��l[���ס�Ƀ7n�s9Խ6#�d��R[v	��L�וt���[��5KUd����^[�-{V2�������4C 6Xߡ���������R��n�n�mMѾ��vy^�޵E�_j+��"sG�@ܨz�<|�΅vͻGc�2�����Ȁ*�b�y���2*�
�]���yus��K��+��~jJ^��tW��{��\W�b�9�Ƙˣ�����p�b���`��i-(�.��{�������J�xd�����3ǃB)���4������>�~�թ����lW��|������ն�ϴ�W�qe��Ċ�����N\��r���T���A��Xf��X̤��tׁ
�e�ˎ���i��K�N [~���8�O��ш)5��6��^�&	��j��Cֱ�8/�\}i�7��&�[O-k�=S��M_��[�F��
s��=���őt��ui�M/L�P�uW>���@���1n>�<��Tk�J��"�ZB��h5���~�,OEg�	����D�%���v%9�KK��0z��\��ܫ:���W�u�<Ŝ>&��g�?�564A+���������ow��b*��\��)|=���{q�nМ`�z�;�^z�/F�W��e�R�M�[u2H�<; �*ύ�αL�j�
k�.�r�[��k��� �|�E̘���ѴV||O_���be�q7�v�c�2�c�Q��Z��I�.�������T����dlm�/��e����i��.�'Xj�V;�tT�Y;x��(ge��Ø{K�\��gl���_��~���:�+�v0迺���Z�ڕM��O�����q]䌾xZ��?~��w^�U����\�(�����]�*ݡ�'��dI��l��j�\�Nj���w��Dp����E�;��3s���.ݕ1QEK�"^�U���LGˠ\��3�Ng�_�6h�`P�w��^��=��Y�#��� uO����?yu鱖������{g{e�P_UCa븡|�P��(f��^5BzT9k�VX�*��&D�����~�[��Y�fHGB���鍬�ܐ��s����5�<�É�t���vT��kn��Ԯ�����`>a��}J�|hXYK�Ev8���o�Yx��������Է3fr/Et��C>���w��J�G4���(�_-j�G����[�SF�����K��=͕��1`М��U}�SK�P�5�hoNyX��/:;cٞy�0$��^�ܣ���=�l:�`�����I"qT��'4���BX���}��Y:�69�*�uɚ�������F��d��1n=�tep맬ԧ5WMJk���N�I�pU��	�[�M�+P�U�\�B=nɇέ�m!BZ$�=y�t�� Y$�9�1�{�8֞e�.�Y��J\{��]<���or{�Ϸ�ח;�vI��N�[�/*�5d�u�J�h��2x���I��]`�SQM>�m����][l"��{oч�{W�l�*̔=yT!��'C>^�C+���l�����x�Gc9��O;��||4Mv����m_�p�+в\�)R�-T�e�f�O+�UyR���T��F�]'K��	[�g3���c�y�­�i�Złz�o��Ͼ�r��m��[q/��y(E=�Z��'�O@����+�V'�Ƶ}c(m���e��������Z;'�M�V=N�������k-Y=>��%S�yZ&�b'2���i_����s]B��#���p�ݫ����ȖlSW(�t��xf��9S���&��OL[N��+�g�8m���!2��%3s����ذh��Ln ��.6=�"�T9�mU��yc>��'��e�a�6������*���Х�eހ��j��i��ͮ;���qX*k���c���&B����r7�Q�>AaVϮ_J:I��Ə
@i�V��"�je��b���ٔ�N�ۻ��\!�ڲ�3�\\n/E��L�X�*U�v^Mp����LԳ3yv���y���b)���ݵ�3<j�� �۬�:Q�L��(u>|�1�hb��k,X6�����[����&%]������̵
�f�;F#��0�Gu��j��M.���5��Nq̤3�b7J�T�U'�jL8�_+��݂�;h�JƳ������J�����|�3¤7�:��+�+��u���.5Z�^�CB{s��袒>��B�ѪЫ�iP�ޣU]pp)�(L��m����`7V��G���o�iD��Y����I��R��j�kpճ�v�g���UK�5�{X��8������-���U������'�g�05�Q���r�!c�T!�YK���@�@M���{��X*����\��I��yg��!�o<�O<�fWqÚ�õ��,��Y�a�4@Pz���o�J�8�ܙ�I�:͋f}��E����
�_F�z�/k�Ks��ĺ�&�*�=�����4�C��x7~65�������/�#��LR���87��륁�J�sx��A�fNz��J����02U/r�.�"�����ָ؞��W�Xxx�]��i���m�|���3;x-�� jRBP��\���d��`���1����΍�Gղ.
���C���.~:�z��,�k+��sFd��u��]�#��PI!�,�n��X����ɛ#k��e@�4q�6���W������P3B�#hT�[:]@���B�\}���r��u,���!�t����Yf�� ��#�K�j��Ce�����N�1�+�rX�~�Aغ"6�#��ۡ. j�oه�e��J����S�i����6��w���`�a\�B�y1b�?�С�[�.��/9�{�:s4��&-%�ֲf�_�eط�i�0%�V]q������$��L9��s�D��9WM�b���P�����6�y}�Y��
��X�ml�u�,
u���uc�O�c�Z	�k����|�tEM�PU����i�35J�/EB��t0#���z�>F�.�cY�t̺�ZU�TE��.�LҔ�J��'R�C �Z��˖s�%���f%�Sv��s4��;/�/>����멷{�}O��Rќ�u���Ta
Sd�2�`l�@_3�Y�bWa�u�`�J���A��l�#\�;2��Te�L�6�ޙFj�_,*%���8�5���9wOgpo3hZ��G'*��-����e�},Ju(�U,��ż')ǵ�6�ܻ�Ŋ�9���x�0�gZ�	���uٸ�C�F�t/x�ݻ��wk������%OVө�`<��'�@k~&�"�ټ�A٘�,U맬���v���ح���0����V�1��@h��↛�ܑ2:IO-��h�ˤ�v��6�12IXs{a�wE҂5zDy}É��Y6R<1���"�P��`���v-��w�*dB-�޽�x-�i��㇬ujmUt���F�u�%�%���$�v9���Ep���:ܗ�8��0=d3o��U��+c�X�?����>�T��[��)H���Nf�*��/��gdѝ-Z�H�Z�i�jO�.���ɍ��KU�^dx�T�Ƶ�w(��#�	���UzYU����^�p�_
mW[��Uڨ���G�@�0m��:����kU���>��2+:*'JP�Nu�913�vK3,UƜ�a�|(��m��X����v]w��ħ��)�*Y}�Xbޮ��l���R��V��k����D�Z����%u��VW8P�,�����I�pۦR�jen25۽��|(
�6V�ԜnĻj�^ڴ�Kp���uҬ��y�Qu&�n
s507(���e����w���`�5�UDV*�Θ0����y:����`ɻ��Ùēb���<̮��65��y�_%��Ř�N�)Z�lTʆ1i,�A+pv��0*�o7{�r�}.��H�T�aÃ{��ڦ��o98�B��h&��񫊕7wZ]%jM�6/xC܅0�N{h��tP�Mڰ���WL]���Pi��]-�� j�e��ۻh�QhVf^4�5/ްF�qڦ�)�8�VSg� uGN^i��o
���*�0�ѻL����g~J%UvZ
*��0Q`��E+Q��*(�-��a��((1*UH(a*�(",QAEm�EDQV(�"� �֪����
���"�[J��e.,**+q�-b��XAҨ���V(���YZ�dY`�EWV(�᪵*,��AҨ5�b�**J�jZ-h��P�mQ�+UZ�U�e�b�h���J2��(����E(�R�XTcPX�Ƞ�)i`�Zֵ�34*(a�TmR��A��kU�a"��ŵ�+Tnl��jV4e��*6�JZ�Q�E��m-J��a�p��V[B�ڍ�%P*�c�5����~�˜��eC����/���1���F�5bΦ���P3�5o���h˦�tSiv
S
�3t:^�|-WK�́[E�]Q�n'� o��Zy����`�#�o����D���l��v����T,5�1\�@���|���q���U[�3+�w)�'#��_�4���tyi��Pp�G���U�F����T�Lv���_���[Q���m�w�^W���Ư�|��q�K�(̮*���r`����D9�6��6���݋1��\{\�����خ}����]"��yj�Z�I�����G>����6�a�yE�rv��BT��S*�a�}O"��U/�6,ӞƘˣ�CPU�}uJ��/_g�̈́�7���=Ad�;=o��?0�'�x����r��6�|�Z.�4���'����Z���4���+i�?:�<v*��MT�X��QXD��ݖ5_��yCx,hg���WG�$/<B͞�Vl"��.�x`�<:L�^VǞ�3�Ҧ�IO�xC�ٿ b�oK=J����m貾�b.߂�>�(STkp�R�
�q1��P�A�Q{�0�곻��^������WU�EUI٤�v�4�N-aP�9�;~l^*7�
y�KA��<KXiy�g����%b��uv�(��Q����7[�0�LQ7���&����Ω��/Y
��;5�
�6�_&A%Oy��(�37�o7��e��.�)c���p]Hw��^w��jT�mW�lB]��z����:u���
+�v�Y󓳶��-I��k�[Y�q$�z5��H��۾���N��*�
���R�&!�Vu���v�u^{Jݙ�Z{���+�M��7{���L�l�\b:���r�IХ��2�^��>���'��3�5�
؅���:��3�˷݇9�\6;�7�oԯBXe*�N�v�[��i�)�A��^:��y�u:���o��|���eM���f���W7��i�#k�}�vyL���T[䃵�p��E�Ƙ��_�Kf��خ������K62�w���dI���P]|�_>��Ӿ'�� �#<&�./����O�|��U�C������z}C2W���F{sl�䏚
Ĝ�6㸦
|l��_b��ٞ�֬�7#���<�t!e��_���9'�:�I��T�T9k����Ȕ���0`��z��c6ė�P�\r����0ڨǭW�o�e+1�p���9�XJvv���\�ֳU��8ĝ���}m�۵���=�b�z�m�ArXg��u�Nޣ���`i��s{�DQ��ϸ��B�c�Q$���=�E�u�f���gw_ר���o�`'-T��k�eŗo��E�w��u�gvM+2���Q���-�����O_5�*�t�v�%�nv՜��*
�X����h��i������>E��Pĸ:��-,0e��7:s���Ic6.����O�P�_8*��8+�iD.Zи��J�멹1��L;�s���B�>�t�j+��J�bX1���2�s�P|*�����%�$���;�֒RΓ�Buz.�A���
�#�`5RVm���)H�*�zIN.�S�+>��bU����:G�:wU�){�F�Ƈ�Be}�5[�z�2�����gB���"�]i��O��ŋ/�Y��b��9��C����t�X��^_�c"*�^����������RȠ��q��]i���0��_eY���s{8ʡ��RX
�mE`��/U�9^R�/��N��^�lT��ۀ?z���5�9�\�q龫f}G�*���3��j��Ey}:�Y_^ތ�KB�u|K�=�����tx�9S6wK�$���x�)q�>s���yֳ��Nϕe�#.$m��Z��R��ܬ�#�Oem�	SZ�	�LC5A�Ñ��e}2��ƫi^\n�AR�����K˂>��7�j�O��ɼ{vz��\����L��4�
�5�F��WS�����W�F��҈{FJ�,�nP�h-�_qd����Q�u]
�)�+y-��A��m�]�s����kr��gl�Ѱ��;�9�lS�a��&�G��KS���_f���(~��e���e�¯K�9T�[3�ܘ���>0z�_.��,���34T��m>�g.�t���7>a���=AP�%�j�-�%�g!��ʈ����y�/i�k��M���+l^��S�Aϗ?I�Xu�ƾ���kne�����WH���{�4�l��IP�m��(,-�[
Q�o뗡��lR����M�ؙ������W��y���f0ᨽu�M���'s�}]C����8h�Ï��Q�e�� [��+�^k'ҝjU�L̿z�>�[��U�9<	�h��L�v�Ԭ�u��MGŋYkǵ5!�od�9W�4�r�F��|Ҕ&C|6�C���l��y<�T/�����>���oW�T��\B��1\����/��+�n��|�N���薁�u�ڗ�䃁�DW���X8�/�[�Z��{R�2��p��5B$�߱�9�/Q)y�b���>8Lp_��N��ȇ���4S�����T�o���0;�߅z�ro�Ȁ�4(���Ǚt�|\�M�����e{�ซ�~^+g���Voe��{�����9HG1J��ӥsN.I��`�Z����ܐ����dȕa�w��Gf�Z�߮�rޣ}�!�4P�d(��Zn�!&Y]vtN�:CƗ8�t��U|#�x\��ڱ+���F����Ub���6��+Z&z�곃��e���x;�<>\�P>Cnd�z��P�<*^\>n�&}����NO]�:72�J�^_N��U��30s�����[{ʸ�Q�y_P^�b{�-L��|��H�i���ne&Sнk��J��f�������5*�T�U���(V�R�Pᔵ�N|8A�E�~��F�u2��t(y(R�#�i��S�蹞8"��GE*�ԫC�_y�J�������IF���!���y�����~�.3��iG�2�#K���%kIr�t��ꚳ�8w�/;�຺z�Kf��%��rc.�P�����-�No�	��T⫧YW������z�1�;rٮ���Y��6��}<C�h8?IUI[-�����]�?8���Yk�|���a�<��7R�/�וX��6°"Cd��ܹ+[˾�1m<��l�Ae�J/>7b/SQ�^ᒶt���s��c(J}�W���Fr^�{���.�iJ8�Xe 6 �uWNZ�A�����(��x�*�]�}�.'�����l_gw �䷝u}�-��Kg��_�����nP�%vTU{���1s/K=c1*�'GGC꼊�wK�����9Rt������ȷ/�m�.[�z)+��w5~�t����k��=i;2��y�|<*���,�񃩴c�K��N��Ӓ���販L��h"��<��1R����0���ij�`��δ��c�窺�JI	`r��6$/ŕ��o�A�]E
k�[�ʔPX_f�aG�?mz�;��]r7;�CeWt�n���$�AW�V��%/&����`���C��x��W�)�(w�̎
������T��5�+�GE�<`�7�eأ�h5���~�; �Ӽ1�\t�qs+Lֱ-�Xүf��R�	�}�f��7"��tx�eq��񚹫�c�%oc�3ۚ]x1�S�t�0��pi�^��6<z�1Gۉ:���/ja�Ry�0����ڊ�=�Nݓ��6鵉�[-�v��VL�<�����5������E�k��33C��1������fi�Ǐr��<�����b��GZa���Q�sZC/�����	�r#��|�_9����s�Ub8GBP��=ŋ�Q-%}\W�����Ii�l�����>\r��&+�E�k^���RhΣ;`�XZm�#ح�ǖ#��a/�$XC�eN��[�yoy"}��_��'\P$:}sWܒ]1��m.��N���V>����
B��O0Yy���j�ܣo/��b��̻e[��P�j��y��nVr5�S���Z��b���V2��ʚ��:yK�M7�j���\*y�R���'�o����-��V(k[�>q�)���x�Ź�P��'��	
�3��>�g��o���)�ޜ����	c�U��r�{U�޻��5[,{�%ZNd�r�i��Ϛ���<��_NW^��^8T�0��4���^������rB�qME\�5S�9����{�;��u���&@*T(�R��ļ��t�>k��XL=��ݻ�^���J{��o��)��Z(�K�GsM�U&�!\���G<����=k��eäRɴU���g���xiٌ�P�:.�W\jP]���uڸ����h��Ƭ�=N/�M�n���T�φ9]�h:�h��b[ V�^X+�샯ƻ^�D�i>��tܗ�8c��&6��k�I���b2=�%es@E�lO�8x���.�*�}IO ݢ�dHeh���L�Y��F^���d��ʡ����^+��0���	�(����>^�M��wv�vc�G۹���[X)R�|�h�� T̥{b_f�֬��k��X���q�eRgj�� ��!�s�Hk�z\�X��w(+k��;}�p�ġmc\֜�V6G���ܥ�T*<hQX��nr֓�b�@uj�.��j�3�ǩ�դK;�W捉_l�x�I���������h5k!�ku<�0K~�Z�WU�z����u)���90���1�>J�E���x��ѫ��Ey}S��Złz�:�KG���׵:���Cֽ5���$�`�_�C`���&U9��C׮����ޘ=c�/�$|עy�w��"L{����}��J��1��Z�%BzP��q��\O��X;�5;�F�;W��3�}p�v�}�+#�h�*��|�.6=EsK��M�&U�����ӳ,h��uZ�V�^n���a��GB!@�#OTLnZyı��T�poz<�)n�oe�O�ɭެ�o]�s8�|�)G�0?i-<u!�>r��g�����{f��u˯���/¤4ա�>�񡾌U/}\���,���jM���.!���¶�������遥dr�a��]*��2���8n��N�'���a&�x������y�w�7ڳPs�k��/�g�״��]�L���m�r�p|�f�،Vf�mbͼ'�-2v�ؔ�]6��� t���z�&�B�p��Г>�Sm���hq;4�W�d��eh��]��|�j�r�i`c��nR<%s���V�ÌMi�͹��;gJٔW*O �O�p�"�W\���G�nTag^w
<NS�t���SpU��ˣ��c�C�TONqC�O�L��5G�v|�I������EV��	��|��N�y�B�W���xn�J_ݲ�T#8�$��� o����&6/E��AA�ȃ�E?����Ż�qm�ho���w�k���/�z�mYɏ�Z����5�U����_�m��Y�~�O�Kzݟ��}l��gz�t�u�r���w��oP�,N���+�a�V=G(q��^*��É(^uQ7SO��Ջۡv��[�})�5�W��<0 ��bfƲ��8�t��q]Jf�gR�9u���鱢+Y��r�V�*����o(!��Q��������h�9A�V;b�{��R�͎�����i�Bm*<�*�ܹ!��Iu�Pr��,�;�T���41�u�2�rƗ��ks^Up3,�cj�ר�½I��A�k�퓿=Ǣ� Pȩna�ݑ���r�%K��z�b��!c*����ӂ�ze[di��hq��u��`$1q��	���ءr�p�k��&L�J�t�[�;5pGR1v��Y�S����Jx\f��x+��)��rX���GzP�2v��74�YS6���T߹	L�y��@Eֱ��gl��sҏ-�)<}RW]7; %r<(
���mEԳ�j��m��v �.�&;��/+2���Fw\J����P�C�؀2|<7�k��ɋ�~��?���U9jX�!÷7-���[��6���w�����ϥ�]�O|����$x�_���=��ÿ�R��x4*s��8�t`�+��:�{m�Ƭ��}���xf�{�Z�M�pe�ޚ�hf��h��if� ������\wNb����E�Mh)�X���#^Z��]���ȅ��I>ݖ5�[�o~�z��۲��"��Dv���f����մc!����b�V�	�|'W��{��;sG��/o;�uq�&�1)��]^ą��A���Ϻ��j>����wQ��Z��r����=j��
QϺXu#�J���*��4�E�"��.y�xѻ�xnB\�l:�2��_��~������VWs�&}�b�K�[Q��W��#p�PU��Q�r�~���w�kF}f3���tVd���[��>�c�-�Ἒ��E���M0/iӂ�A����I���2����ț��}��є�]fl.��aJ��k���U{���|�*�ð�] K��)�*�}ǃ���o�g|�l���a�壦�Vl���[Z��X��ۈ�5]|�έiq!�s�\�p����Z���f���s������.�Hq"��zt���
m�ӣ�y./i��$-��':��rζ��wd��4��.�(�]�'4p�b�,@h��m������:�[d<۵� ��Y���Rtuٔz]:&�v�  ��D�3%f��f�EA3�k��oQr.�oau�V��C����}I��xk�Q ���0e[�V��Z��B���E<pu�ҚQǦ��t�v�zJ,m��"�y�+�{3��'DTg�7�'�ӪCd�_:�]Åj�g�h�7���)�+��0�&�{����% i�L�Mڹ���v���XY�ǭt�fVV�tv�\��-8L���;ve)�X�J�C�dU���6s���>���5��:�w�8�ge��e;����[� ۆj7L�e�����pD��/���QO�;%[�)&V�s��|&7M
Aе����t�s�u���j	��[O2���Krdm��}XSu�����)[R��Hm�th�Y�u(��[K��|�Y5��#h��΀9�ߙjkd�ZŞ����V��b�Ȥ�wV����㏻9.�i�L�-WL<����T���B��Ym>�6����#}�s[ͦ�틜�s^n�����Nh�M\1�3L����ط9e����m|Y����mZP��y�w�R���=ݴqu!��!��b�(���m��X�v����X�FSu�t.�ŝ��4�kx���zL��(u<Vy�	]Yi�����[:)*AV�ߥ��$.�Eh{ʕw�F�n�f������S˭�v�[q��&�Y:�)
* �0�b�]:��:��  ��}��Y[a�%�Z���O`�)�lʘi�N�.K�G�t��+�j�f���+%��]�[h�w�~9k[k�H�Vƀ����8���p���#yR��!�P�N�Y��]�E3��^Pw����(�Ѡ��伦^)D�t�X]�wΤ9+5�֪��u_3�g,��P��O�뷕�4�.��� F��������������N��ފ5,�>�5ћ�n�{V=6�7D��n�bh��	G;�,я/�p���-:�����A������v�ɜ��n���O2�o,*=�T�s��E�Rl�+���e"�h�F��\��"����dZ��_ؚ�Wf;/���)��Eet9D�J�9J�F>LvM0)Dm��fib�O�#�m�ȥ�=r��l����	>Lf�?*�;mP(\?g�[{a/��4�L�
TG*qd�A��0Z⅗Z3�M+��6��#M�Ԭ{_�a�M��m�7D~dz�����5�VP,[��{�ֶbr�뮝q�o�w�7���;�]n��Q�[Db��5�U+[V�-���l��-�1E"��J+
�#R�ѴD��QIF[V��(�PS-�Uj�x�4���
��(�UF�[��j�E�#�Ec-
�����k*��*���Z֭�X�����T�(,Q*�m�h��[TTdR�"��e��TkF,Kkmh�ih�*�c�b��jҴk�c�l�-���#m+,�-��*UE��2�P�dV5�UjUUm(��6�X)XX���V���T�R�6�T����چ-�EjS�?"�E$��$���}�r熳VEDvWj��t8[��y��RE�ݡZĳ�I=�*���+���h:Ӈ��a�<�'3�0��Z�L�X/���!A���gp�V��E��Ϗ-׆`ǴUΰ�x�+޸K���#l�^
Y�9��K�J�1�;>�ks��DB�*�x�JS�fr't��t�yM̭G�S41���B�f�˯_L�㣝�x���*�W�lJZ`.��������Wșq�8���vz/G*EX#�r��ɮ�a�.L].U�(�M�gIS��5�,J��A�.�n�0��xg�r%���mvNj|��Ϛ��C��Ϙ���������:��%������8��zl��z�v-���3�xl�ɳ����5FZ�wX�P��cB��E��	G���-�z�=w8+�j�%W�V
ڗ��S�pni�mc|L�Ǩ��^ʲŅ)��A�C�'�9��-�yS{rX}�n�\"�K��
p;��D1�	.,�^�.G1ł��v�%�k��M��!�ԨZ6��C�'��{�cl��r����A)����.��F����K�7����v�Lנ��͢ �������u��:�
	�{oKKn�ЃOOt`�mG��Л��FN�}]�Mr���Y�Ӻ�`�*E6ތ����#]=�a�$��Z�:E�MYca�B���gd��3+���:J̥%K����X;�܌^�\1�c��nkV`l�U��{�z��`��U'GC���U9ė�\o:��u�y;t,�p7�"f�W�⿍�j+���z��<�zI8�em�n�����k(�l�ݐd�����5�R�*2P���W*�t�X;^�0r�=/��ee;]�������ٱ���g��hav#���5����j��d��lB=���n��P/ee��;ϸޮ��B?gs�և>�z����ӣt�Sk��W��.΋�ȠўR�)0��������Q�����]B^�ǒb�F��M�_m���g�+s��{z2z�Ѐ��F3w��j�EӞ�U�.�~p��l\��\��l��
�k&����򼫰�K�;��R"'���ν��7��Y�*:5������%�PĦu�	>Q13��ނh<:��>2�*�յ*j���[Rfw��*
��	t=Vu����[�K�9�`Cjm���Cn?],!e6"PZ����:ƺjzJ.��C�Ң���%\]�,w��W4�}�S��x��b��ZM�ɣ΀�}z�?k����qCX�����T��W�N���;S�t��,;@F Zl`}��m���gz����0�w�㔻k�e��o�gi��BX��o:����-˧�>y�g:�஛ ��	I)7b�>w��D�;�%�_lמ�~Ȧ1sh[m�z�@3�'�G��
�ge3;��|�C����&=��Ͳ��>0W����4��$v���߄PX��e$á�b���z��*䴋��I�n_�>��Yѳ根���\��(OK�E���刕����t�}�8��kcG`3Z˦�w�^Ey0��p�3<k�QT�fr�^HW��0Q�a���׹ky��pc��O�sgGj�V�ھ'��,����U0�*�x5@k�J��Pc螟yw�C���Q�;LhU��*�ժ����a�^uRPu�߯" �o�jmwL�X܌'B�t@�����u'ӯ�P�^�P�?�e#���vr��1j�,��|�@>�Z<�X��
������ye�u��qz��J������B�U��리c�|0T��i�kOz�u̳>��z|9x��8̚�>���`v<9JǠh�{�X"�Wh��n�ɮ���3�;��}AW�ق��VI����Nt2y�k�G�r�<�l̆*�p��+�lV����
��`�7�À W�V��Z�P㨶�+�;�������4��QTG��m3M�Ð�ܺ��*�?�x[D���9�]�Q�X�>���1|���:6�l�v� KR�4���X��;�񭢓.���ivs��K�ʳ&s�^�t�\3�+t=��O/od�X*����NOŃ���?[�:�08O,�c�W�\���P�(?U7�[Hp#�.P��k�J�Od�%�=rή�͚���W8���#�x�:���9g�_Ⱥ�|��^i�N)��!f�ʫ���fپ�j���؍���������8\Q��m��F�:�gz���f���CiO�nKzHk��튅7�ő�B�XԽ�x�q���������]��G�/�~Bޭ"��҃-X<�����ܧ��
����^��Є�F�w�cX�۾,�m�;g�[��BP�.&Z$����PWD���烮������0K��EG*�=�l�n��7�-�u�o�|�R�<��|2��~γ���ͳ�3��2%�+\b2=����^�����`��^,_��L�"P�%O�[<v���v:���V,ڣ3qe8�J��Olo��%���KKhg�â͵�[A0R8�'��#�ÎwjM�vM���#n�ۡ3̂���ۡ���wVkiA:tKu��To��+�\��.��]CY��VZ�P�Cu�g���<���w;i��&�0�S��ؖ7���T;��v���jS��k�[���G]��z.��(k����`���ܳ��|t��גI����?
>�2���Mq�Є�EՀ���k�(���à�]f�,lk�_��v�qH�{��]�6�	���݋2��J�Ң�E�}�%TbȺ��t��[W��(b�t!)9�op���>fg��mf�Q���Q2���5�Bv��w��A�Ż�ۏaY�!� ʛ�"${J�Ԏ���j��#!�6���!,`��<@�s���5^nE��*cZ��«-_��ǖe�y��r����gT>�'C�P��L2�>�0�����Y��<τ������g:LnF���J�%��pU�Ю�揷{H���J�ܛ�{�Γ+�zr�� ϭ�����J�y�)��z��>Z���RZ<#���蟌�3r�S�����.��+Uz�=���CLEs���v�Y�Ez��WeM�p`�#�����{��(�	�p������!GOe'֤�,�n��7��vO_��[�o�KXY3��T�\���PD�>��r�X�`�XB���[��>�a}7����a��abo}x�g$D��[�l�y���Ę�8<i�@˭{:�rRG����Ǚ�-�
ZVu v[��j8/��/�
XQ=�a{/5*AϠ�I�K�9VR��:�9��B��{'װ��n�0��S�j*�,$��v�-��hoX��5茘�m�q�b9�+y�:���У�w�Μ�����'~�YME^��/�/.&r�qd�诖�(n�7J��*�+�(�ƇHG�i@u���]fk�xo�ۘ���Wkњ�qq���R�x�S�3��X.�ET``t4�U��9cQ���{3�^��'!{�D�ڊ���W�M«��<�|�G>|*��
���wy���%���|�a�*Z�YUBi�GR�7h���踨�P�1��Ӛ8ʜ<��/j	!�bM��N�9~�Bq�Ih�(p��>: �~3�ͧU��ЈK�[�{Z�+i�Ba�`?]��8�sFS�v^����^�U�5l�}��|΄%es@L݄f�����z8;�F��cI\��S��o�E��,dr����0+�O�/w��Â\���o��<{�]J|�D��������l1����Z�5k!�k�^
��͖�ä���횂�S�p�w	I�/�����U�l��ϕ�u�Zpn5�x�wS@Ĺ�*(mn���.�r-G�r���]rַuєF��]m��I���+슘��2!c���*�{||g%X��=�: 7c�n
��K��ʦ���V�8h}O?^<�Lc���[c׃z>=ҋ7w�P��y�;��O�H�egr��Q:;0!'u����p��m_�'C>� ���,I�o�e���S�Ε��W$����y�g>��)3*��9�ᱵ����%�^m�	��N�.nA <6�GV��^�Sʫ��7J��bP��s�#V ע�p=4/�%�ߥdX Pј��`ԡ�s1oW�[�3�;��<'��fm��PTx!K��k�4��m����3�w�_�)&����47���N����C�����.`�\UM�;^�*��߄�]w���(Y�F
��L�޺>�������gҭ ��(]+����eB�ϔ,@��q������X��¥���ݎ�Q�t]�>W�9����ͺU6fR�F���%ԟ\w׾�Ť���=��J��W�3��>x�$��Я� �s�z����Ƽ�@�*�O{ڹ�.͢�3d��T��t2���-5Z�UQ�wz��Jg+�`J���W�)B	�=��=�9~�J�g�S�>N�$�\��u�!��KN&��I��<je�|en�J/��1�!��.���cP���:\6�}��#����hZj��M���2�s	���.ymuǃ-��	ô����Q�+�u��]1��a�1ԴST�
�|�l޾�����2�]1���*���J~�#�Ho�EU�B#~�]�u�kr�&�u��S�Q���kȠ[W,�<�k���l�ۇ�83�opF��]���_������t8~q<�_����BcF�Oǒ���\]r�!�ct��ݛ����&w�%�ʱ�r�(,j�*�:V�q�+�_��N����^�����	����ĵ��6���f	Qrcpۣ�>�+9��[ʼ��x�y�<�XTDJAf��A���d�w+���̕�@|3�z��N��̬��������ܷM#�G��4��\��j�ke>��UYb�?x�Rqp��A{m�N-�>�®=Lk��\ñ��y�*_�w$Ym	�-
���@���T!��ҠW=@GӜ�/�z׾�tޫ�S�AE��Cn�ٌW�����/B�2�."Ό��ר�Y�pcM�C�:u�8q�x0x)G�=���Y��/�t����ғe䮌q�>�K�:'�I`����E�����6g�`b���/^�g8��*���z�/�
x��|z���-�hN���G.x܋_6�P�4�ʲ��{jX�!÷ۖ����X"���Z��]u�wޤ��C�elǠ<d�b���va��uei4FWq�u�;����\��Bq杞�5=���zy�3+%%;IWGѷj_��x��#ȶ-�S��}Y�T�a�F�0����0�oo%Y�q�����������7a�
�μ���<��y��
kY�'�t�g<ҳ<{)̉��<�j����K�5ҋ`�ս\Hg��.�u�5S	�~���R��c�4'�H&�:	z6�'��M0UK�M�zz�+���=�R�S��K,UŻ�?6���c��VH�\��*yCb:��E��S� ���,}c���&%l��l,���,M��}�5~Z%:v����M�T�(Kux���[�5u)�aH^Ǳn�Sؕ�Y��n[T�n,Z,%������(�s�*�Xw���NkJ��Z<��^�};zL*��]���x�冮;�����f=̙=*�R=b�����\^���KW�y��ܮTvA����>Ӑ�y�W�������[��P�jV�hM��o5���o�`�~�p��uF��j�Ea��bN�!�}A3���]�
[��9��ޖe��s��c�ѕ9�
��պs��p܎�z��[X�*�-�Î˻�����Nŏ�m<u1�f��u,k�M5�0]k� �"�65Z�|��)���Ŋ� �@ͮ޶���B���ƻv�=���Jm==x���}�2�G����j�+rY����\9�`@�lը/Xm�0�ڗ2�Q���Ϋ\��Z���
�t���/Mt0�I�����.=�^͖5�6�k������Ǻ���Ń���}���tJ�`�1�C�љ#���vz/ ��*���LR����^˱ۓ�y|{;g5��F^�����Yc*�^m��l�/M�y�9��p�A�'6h�2w	��V��UM��1��0��yx_��k�ߩ�(w��[��[-d[�}B�<F�O���0o�_p�� �릏�B�Qw�̪�I����R的��z�y�O	읆�΂KƤ��Z$tX��0���:k�!9��X��9S�#%����ӏy�j5W����X�v�	%����VX���>���.TF�mАzrF�`��"�o�W�����3�?�K��)��UX��&7�(���o6P�R^��(�\�q��7����9C�����Qw���9\,K��9dz�ɫ}]�㫀E��R��6͖O�YM�u�eRZ/�|(�x� �������&x�}:/����̾�I���N��WگZ�7:�n_t��/gY�������Nʁ֠�8�.:����'6��q"����IQYZ���nϳ1��Ց��5��u%�f��JV�e�J"1a��b�U=X$�/�v�y�����WV��(�:.ԃ��*;��t=�h�C';�r��\�����#�;NH�u%��vL75�E����� ��a�؄���h዁�$�xԿ�%�2en��8[��:���!����z ̥�&�dZ�[�Qåހq��K�<�=�ڝ����yӮ>�O{j�0~{���WVJ�������f
��ĩӳb\ʞ��Hn��O�G��oR\+:O�o٢�2��O.��};Z�k�K�vP��3��U��J��wS�E�ݺ 7{kͻ�a;(�_�o��o�v/�ZK����	p\�FrW�M�Z�Ml�����g:׋K5'uw��@���}���,��M�27�P��j��p�W<�������KwYk³��s+D
���w�Idvx��}�A���]ڍ^�V^I�8��B�KB�X�i��Ԧ �B��b�����'.Z.D��=׫��Բ[U�K�8�M.�<`X�;7#U�y�����-���fS���fi�I
6���[/��07~���o2���Ǒ5��TczV�7��ᇎ.��KG*�X색�9�\�VU��ߺ��:땤�\��aw5]9�������B�Lt��%���w=Es,;9]�'d�V�f�����4f�xw�coY�A�uw�BڽR��c�<h��nG�iA}tp�ԈX���=(�F�����4h,���}G�|�w1Wβ]t���;V��[3�vt!�ŗՒ�Эq��UvRP��	,u���oo�l��f	|n�'�T�<������J-р�i\Á;9�r��[Uܹ�	r�V�-�y@�V ����ƭ��-^˟��f�6�*
�6���H^�Q�Y�;�+��kT�i%ց|l<c� DtP����vѦ�&�3e���F�v_C��Э��( �z��Z����h}��P��)}AuԬ��TZ�������p{M��t2�P������CU�A�]�Үg�ŻO&
Τ��y���L����[��ShN�؉��V�yl��v�v+9n�B9�{u�Vy2��σ���U���V��co��Қ�M��M5�x�q0Ej��r�+˳�f4ʜ�v��ڊ���1#R:{��@�5u���H�2�]EY�mg:��xɕ(vȴڔ.Vs�r���Q%�6��VO@\�㏳�J��L޻�Q�����j�<� ���iH6�)bo-�U�}tǯ	�1|H�B!
C�(֍JEE[j#R�?��)Z6��m�U�"F0Űb�+m+Y`�*-j�DX%V��j����aU�,*+kdT��Ҩ,X�KV����[)m�����4U+U�J��6�[K��)l���amU��ҭEJѶ�[m��J�����Ѩ�ĭk����Ѫ�2�m�*�ڥ��TV��B�E�
�
�-X�cj4*���m-��"Ұ��s�	�Ej�cm��T��,-���VX��֥�e�qp���ZR�--Jز6�Vԥ--��h��jUV��Q��Z��J8j�	ZT����>6�Ԗ'@2�}�R�Z�^QR�]Z�i�}�:�ړ�T��+�t�f�9�e��+���R���qF�wikL�W�{[�� W�b��n]��E�T�-��ԏ��_�V�,�a�2S:�Sg/DC��T̬�^Ώش���Ə>�*�?�����B�md<��˿:�V�B2l�J���O"�}ʹ���yf���u�Љߡt�`��<63鼷��ѣ�� �꽕��d=m`t�Χl���n�C��xP��@[����[c"���Nb��>�sU{~wKkҴ��J�N<�;��ｓ�ǺRL ��W�}��^ۀ~���퉗:z��3�VTו�X���ʼ�W£�؅�M��fVJ0R�_��ŀV�5|���n���2�LL������C�/}��x���up]ǔh�Rs�P�:��|ha�G5`���p=5|�.6=EsK�ʩɃs;�c��!C׳6[N��6�UFPc�HuE�eMpj����cT��
�/�X�������z��׆��7�y��^�qs�W�FA�����Ě�-<�k��kr8��d��̓����!/sr��\ι��5�#�Y�6*�r�;xm��6|`ߥ&<P<Ėz�m���C�;Ry
[��!�ٷ�u�|k+0�ㆼ� r7sK9����s�m�˺ʫ�.�5���K�M�a+U$@-�ոo��\��d�7g�0�&�}���;��n?w�N��d�%y�6� �y��5�����g���w��ߓx�=�z�Z�J�!����d��R։K�j(����G¬~�`U�ؖP�Ԙpӵ�R�J�$�a��MWB��q,�N����$ߟ���i��Ҳ)�a�'��Z���]*��x@nХ�tJ���@ǯJ�������kQP�����^Vt�>�����T�;܃bz��~��基K=�'��֠��A��p���t%������z��T�}~��^��3*{�2-2�:�!o������:[*!����%s��j�C]��7��kJJ�\TO�`�im�������m�4����\<9�ES`�h����S]����Z�X��IYl��ם-f57f��5'8|o+k���u�XD�S�����i�?W���kA~��LY�f��'����(��n�'��Ix1�;��.�{n	X�x@S�Ng(�dOդ++;o2I�^����;����X��Er�1�RV��{lBqkPC�S<(AX�f�m��k4���ٶ�b�,N��1Q�Ҍ��j���6�T<�J��s���՛l`/��"V#�@����z*=�pQ�52��<k���,k<,ຐ�mɭu�ӛH]�����2�Z��|D5��rgR�w���ܱL�J[u�(�'ؕ�|���C�{�~Xlg&�9{3�h��"���h����+i�7k��SG3�/vM���e���O��r.0�����ou;�u�w.�\c��N|�̷���һ�����06H�'� �/���u�h��퉎3y�U�(�[g�+&��7uM�u]���ϕ�6ePX89��:6J��cgݷ,'���R�A�2��:-nv�?F�<���Aϔ~<��p݀y�z��Kid[Q���v|k�]��� �|1�Oo7���zjTb_O���g
>�ԭ��5q���^B��+���I=z<zx��ј�;�!ʩy�T,!��Z.�D�U.�T_:�&�W��U"�f|5Hh�g &�8Ty�Β��wا�"C���9�M�0�^-P��
������]�3ϻ%�Y�G��/g���Az{�W��q��i|�TI�AAMx!xZ��[�5�D��^��w�zb��ބw����,��7���3͠�������Ң���=������㽄-�����%��� ؗ��ڮT�=}����`��ʎ�Mɼ7���n��5�Ei���s5u��l�,������Y�!�6V�z�cǻ�
�XR�;D|��e^u^$�»2�n$���9����rTb`ܮ�Xn�ǔ��-}����7��͆D�XUR���K��!�Y/!Ϸ<�:�%-h��(��Z:�4)��u%]����盍دW�%��4�pԥa�򸲗�b�e�dTy��lW���o1�s�]�/ݚ�����]�����ǖe׹���b�~*����wz����fC��%ʼ�/rv��4u��od��`��������Ѧ���fW��g&j[��������]�v��Q6��z�Hz�j��
�k���b�|�G�a�Seׯ��mfuac�uj��c�ߕ%^�����+�u�ӂ �>4-�Zlr$k��Uw�39���`<��G��V�#�:ߠ����ϡ���Ueg1���r��|Yc.[%��`a�-�ND]S:;���B&����[>զٔ]���1QEK�"^�Pʾ�1ݱ�j"��a
�����j����m`�:_2�i��,x==��-Y���Uk�S_����@s�y���}ym]٨߂g�%�B�n�Ľ�R�5^r,��6(=��%Yb�P�D5��Q<e����WS�!8�,ʱdP�*n#w��䆼R�����%R��v����l�Sl��kZ�'���xO
bbwfiY�X�
�+2�d2Ų����7z��g�;��
cs=NT��	���ƺ��^�OJ|X7 �����1
�����ay��ky}X$x�Ev��ޔ8ĝ!`t뽵��U�/��6``t&gR�˳U���{&�v�>5�QE��e"�\+�L�NE~2�C*;�n��PZ�*s�b��Û����n�4+�ޔC�ǭP940y��ݢj!�N%��}�7�N���b�\�ۿg��" }�։c�|x���&��y�*�ᆢ�	�7���o'f����%*������$
�Y9�������
Y��I��� t{½�x�Ō���_�#�����耊�̞(W�������yj��G*�^T����6�ՙ�ږ	�����u�X+�b]A���U�r�lO��o-��ѣ}��8f�]��ȵ�I>��N���%�x��<��x�5>���(g��h<~=}]c"���Y�t�891�����X�Z�S���9�s]]�e���hAd���r��� o�t6'|!|��u�}��L�z��RY�:�="u�mA�2�x}VugԺ��G��;��ۂ��J�����Qد=�������rљ�����kޏ�x[�+8d�^�(�o�$κ�{;�N�Ժ��b|�ֈ�*Z�����3�v�o(�Ra�L�sFWu�EN�+e��![7�Ls}n���\�M7\�[1s�r�B
;��_S2XXu�f�Pϧu.k��PO���{p&��W��n�9m���9��y>jA�3���L=FٟV�̳���*�b��sV|ע��_>K��G�����ʖ6Ι����N<Z��\��02��ͰQ���T��*.�(!\�j�k���=�אJ�4j?[���O�n�>��S=�8�q0�r�*��H`: ���q�מ[�Y���y�]	��ʦ+�ۃ��7Q��!r1MP�}i���9>P�M1����+g�̳��u���p��/� ���`���+sp��ͺSfe!l�n�x/+����C��w,ʀz�?��U�X��|���v
]-K"�Ϛ𭕤�S<e�k���ow�֫[���3���
j�-��
����.4+Z�)|-}�j��#Jg>��}q�r�7q�7�&��}Cx�� O���BX�KW��IA��� {0(gٙ�=���Iر����it+�Tc��-v�$U���B]t�>i��{ةn�y)���;�_�8߉B���Ym���j�S`l��ioӋÕ~�A�
�+��J�I��u��p_,�op�;J7x������>����L����Y��<�^ ����Y�N���f�C4d|��W�
�c7��܁Ww[���e���<�U�G\Xgu>c��[�)%��$o�G9L}�#�]��}MX�2���p�k����ޱ�3y���W��{���b�e�Mݽϸe*��T��>n�W|�Kk�^R� 6��g���X�ŧV׽��mc��]���eMm#�, �i���}���g�X���PC~�>������<���x[��1���2kZ-��<`.���T!���z����|��0�s�k��ƶ�3���Āz��Z�x��r�F;��`�+K�=�9K���3UX%�(���~�M������:�����;��L���
��ʃԢ]�۶-���U���ࣿ1�/p]Z���;��8 nV��ϴ��K��H�k�بW�o;�>����P�{�v�ļʓ�����	!*��,�� ����<�=b�ږ:�C���6���aײ��cܴYG������)rZN?�Ku{B�a��/~w�^
d�;<�C�{�2�������,�#��L�W�yoM@�!y>bW3�}���.�f	p,�:j�����>��)�ƴq��g�^f��97����8oX�ܜ�n,�������ºAQ`���<��+x�֓9�\�!����U�T�>��`��[|*�t;3a�6��c��`��i7c�$�J�aݩ��Ƶ�Es(���U_N�[k��[���{�����*�9�����N-V탲��D�h5+�֑c���N�w�>�ip/s=�i�W�f�,Y��cU�Χ�17���\+�O�"��<�k�
�~ed��/c��̛�e����+��C�0��Cyux��f[JǺn����֝���Ǚ��=K|Y�~��`z����wK��*+�h0ny���e��~'���^���w$�x�4�KE��i�<�X��/���`{�`��ujWnfŒQV�svz�v�J�;;��3���M�ϴ�>GE_ٍ�ϊ�uW�����xg�`���z��/�g�(�ή�瘳�v<�}:���S�T��q��>�^���F�����38tzߝ��D�p5Y������3�s���t�IK����t-OT�LB�ݓ��<���X�pP�P���Lӆ��@���gб�k&�[y3����*��P�k�����ޅ���l%ǌ�zh\d��|���4fG�D8��9�����T ���u�Cl��:ùa%H�ͤK����;%g�p@�i7:uƬ�_^���q!o���k��{7�0���X��B
����]��ǒ�<|Z���@�y����(��B��}�=�����6�q���Ww���q^�h��C�D>��S�n�ݫ��7D2'�BP��+|��GZx)võ%��H1o��꜈��^�,�����<G;ײ�e����m��lʆ�����P_���}}l*Ɠ���;Js�\6��ɇh���ӭ�CeYy\o�_l�MQ�hPg�'�Y�0e1��	è��>�^��.�O��ь�^5S�\r�4G��B�	��c�����J�z��������ܼE��Ǜ��>��`�q��,��mg�Ҭ�u*_(KP�T���Y�U��US\�75�ЮJ<a��j�qb��]`c��^�	+���@��50ϫȩ���Λ�������
���҈aǭW�"����K����,��TM���{Su�Խ��Nǁ�sG]K���~R�zsN"��z1��0(s��]��ܫ��t�4������t
wU���*���Wn	]�V�8r�*�U=53ۆ�z��o��3w:x�G��t �9�"؞&o��-�
.kEo��h�_n?Z���<�[V�B�M�鼹ߏQ��
>j�8�u-���5�djh�.veu\=}!n�,@��\uY;h�z]�y+��s�Ehu��F����67y�ɇo�r�.�MuN�&�@n���=W�w��ܘ�wS�y��k}`�U���)����̯J�S��s:��fW|�'��}'<�v��WK �_M��:��7��NJ=���^-k��*PP��c���?�+�dô+>s\
�M�6�2��[�I�f-�r���jՙn�d�%�tx(e^ۀy塰v�b�*t�}�Ph�pfVJ�J���OwL���B+U3��>�ւ�W�c�K�ۂ5�`��v�U6Ga̚��ֳ׋߿2���^��g�=:՞����:��|ha�9����%	�O�Ŷ���.޴�.g�f�2��b����1=W����u��o�����5�x#OuQd`N��/����������e����9Q*{{<�ˉ��e0Wӑ��z�}��e>�Z߽�O=[�8������� �vS�θ:�uz�)8*�r�h��eB���S\���m��y',�٘�o�� ��N�:_��8�z�E���ҩ�2��_�*��oQ7
��&�Is�����/E�p�[@��_���^҂��p?U쒑RwU�-Z�%�b_b�>�8���o�MT�j�_^��n��a$���d!��x��eFz���I����+��7o3w[��+�{�V��Z��վ5����"�ܡW(�u��A�4I��q4/+P�{���D���Ku�+�}Xt"y��Pzɓ�7��f�5J��y�9g*7v��|P��m��zYp>�J��Or��oa��s4-J�x��0v+����y�����v���D�[�$�۩ճ�[�y/���r�oL5:�Nf�Y"I��b��9�U�*�d�u��c��Xʛ�����/�
C����{��P�=�_rt���DZ<$]�X�\�-�f�C.9*g��ۆ��Jbm����G�l��/C�#h���%kEŔ�
Ճ�2P%�n�Z����d��nX�'���� [*]����v�XV�����bX��(g�Z�0 ����J���A��n��\v�m�`�NM�V�DP��L�ٯ!�`��Civ���֑n'�]ڀb�z,:ڼR�rfr�L����9g)�����Ff3��,�5�S��R��<fc��yZ#�R.�����ŷ����r��3�E�{�nh�{+�(�z�]3�Nx��UН�Q0p�+�<(]�0H��̛�YM��ݤ�Ç�q
�e����]��S;'Y"B��3!��@G�t�W�Q�ȁ�}���h��sP[�S���_�S�i�����ñּ�`ۦ1��(8tuM�Ooi�����э��/n��k�@8��̻����i!3P�8u޻��3r����ؗ�b��ו���5�"��Pcog%em�b̕)O�$�5���L4�'��[�uh%�W��7Ь�]�j�Oh�iu���iTx�۾�I�t��U����S3.X�sBW5k��P�nSr��9���%� -��k[�̂��gtyϱf]��J�BY޼U���P^�J�+�
@�o�2ۊ�Y9;4%��:�w��A<A0BM	���L�k'V�0ˢ�tC���oH�X���l�	��]�H.KM�N�଺mo
4������^�[�귕�Q��=Տ6���%9ɬ](�,���0�#�I�6�V�X���rs�Y�,nU���-��n��c��V�V_˥���j�\��},��s���i>�8����e�AQ�QVP��	�"u�;������'x���	h���=�j,���Ճ.�T ����6�u�k:�\*�s�m��Ͳ��3g_Θ���f��S��99\2�6��{�k�t��x	��c�Z�\D��4��cK��u��YY,��Q;�p�I�sk���}"��i���_Lu�;e��mvaU�-�Wo��e�)���[���tL�;OA��hX�'��M�w�����tJ��s԰�*S��ASg��r'0��R�weHTμ՜����LYji|D�Obɍ�Ӣ�˞|�2(�R��K��UV,���ZYmK-��,m�[J��jP���)JV���XT���-��)Z*��e��-��/1�FDB�iQb�KD^Za�l��4�E+5ce�QE����(�(ڊ��bQJZ5++PiDZ�X�D�X�������F�4��m���Z�+Z[eh�%h���բ�Q����EZ؅j��JZ-m��hQAb�++��Բңmb�dZ�UUm�����JTb[EՊ�1QcET���iJ�-(-eJ�[b�\c �P�����JW.s\ڌE��4Q����ŉmQ���K*X�)qf$V(��L[D�T�T�DH"�P���"1V�PJ��Z(TUP�>���sS}m�o|N���\V�8,F���	T6�3��3�}-h4�L1�pr�hۆA��t1dٶؽ���T��y������[G��43.��Ϋ�XT��)K�k5S��2j�AX�m��z�[������s�B��g�z|0�'�>p��10f��JKN'���+x!5�˩�^E�d
_pJS���MG��}�a��aT�t!�]��q~-P,"�h�Z)���x�ޚ�&ړ���{���
��k��_�pϷz������3V%Bqxr�N�˽��=������b�J��鞥~��Lh�(���R���R��e���a�uy �瞼�'c�o�m���Olu�қG+��E�/F��ឋFW����	J��� ϩ��w���
�ZmK-��5by��-��z\;��<�M��׈�VF4�J�`e7C�X����:�/P�t�<)7ɍ���X�/�����ƕ�UY�Pt+M�;g�� ���;g=�j�	J5	���.���^ܓ��z.*�;~ite_Z��ԟ,������t�����}�I�u�\��L��[90i���ѽ�����ؗF. �Y;�/o��v�V]
��,��Vo���W�D�{ǹ��4��v�5�� s��>R>�Q-���r͚���-ڊ�����9��/��P���5��l�]����k]wb{xr�蓎�V]�Ϙ���%a&�V9��v4�إ���6��m�A�᝽0�͉�-�,���ϴ��j�g�_��'��.�*=�u|zyIc�q��㊙3i�tz�і�4X�q��YC��}�c��ò������e?2��9����z��R���U<CC��Z���Z���uCz�����E���j;����u��l�w��h�)�ZV}�3l(G�1+���z��M������[����$��F�O��9�<��z%�r��qh���"��v4��������诶���'�Kȸ襔r�,8C~�ƫ�yC��O����I<��h"�ʽ�Z����Ϙ�l�]B�k)�N.��ф���ҩ�B���賤����u6k��j�RFl0D�иeJ(STkp�&���7���1�@)G�
o��ߥmB���s���G�-^h3y��ɘH�⡠4,���Xo�������|l�+����x�����t����W�.�k#պ��Gd��aS>Ӑ��GE)9��({ă���[M.�ؕ�vNf���%���1�p���h��D��k;��xX0�΋�*u�K�7��f��#��`S�Ok�-(�Y;Ҡ�'�ح��uѡ�z�b{��Jx3z�t/#8U��ÍN��u-ɼ��F���k�m��Mw!۫�q�3��tL����SUxh����&1����w�bz|��O�Ba=+U��N|Y|����P�ϫ�0�,3��v���oSђ��C�x�������jZo���D���%X�W�v׭�US5�Êcg�#��lҞj��cj�,��v��{xO{�c���Ұ�C�GZa����w(����v4fG�C83����D�
m�8��}~���֕+���J������]�>�v��.�0�"Le�d��n�0�z-�7s�k��^�<�ȟq��-3sM��%�up��j����z}@�cq���3u���ۭ��H3��vk���*Um��ٖ+��xl�2*jX����u��.y��	�������9�׉���&�G�|/3�
�^\`��P��C7��Pҡ�YrU�,S�Q�x��mwO��
�z��-��yO��	���ʮ�~�1��J������8�]g�(
چ�"==/�͟�D�h�7}tC�1q���������X�VD���9�S+���{�O�����Ҷ������v�������\��=�E��}N���t�b����W8W�Y�!7�/d��-��ݸU�&�e��eNv9Vr���'
����ZS'^���ƒ5(n�uٛ�n��]X�V�S5���!��,�{1��G1�
�iF��U����XoJ!�z��\m��w �A���B��h�x�fL�#��){G�����eT����t��|=�>E�+m3�>��D)��0z��'b����'��C`xʡ9��ӼlK�k\6���C����~o�]�r{�KŊV{���A�W4US�S���?]`�9[�"�!h��-���e���?N�&�~��L�*b��ԥ���W;�	��66���>�%o�]���f��'j���z��o{����S)��\�|o*
�t���p:J�UE�����W}p�{��~{0[?AO.�DÁ�V�NM\p�	5���\�
��]\�f�����	.��켦knMj��U�[�/��Σ���]h*�t�c0��pBX�5L��ҧ��m9����7�=8L���~>j��P���rY�9�_5��zeV⪭iSvR�rl�U�7~�p0!�6ؙ�����m;3�>*����Tt!_.b���]�Z����^$�dQ��X�]#�,�/xW�ӫ�����)��{����ӖV��C��V���q�vsmj@�G}N
6��^P#쫒�����*��r�t%z^Tύ�!z$���݊�ȷ�U��S�z��p��f�P����٫��V[�+眼s~|�3��T�S,y��M�j���7��2ع�qZ�f�֍�<�e��l'����Հ���&�^;C���^�����U�f��O��iU=j�e�m�n�lo�V��T��/�w���q>�z��X�ǭ�5&Vb#ٶÆ�˩.y̛<3�w����Q~֩1>�rNO�5�
$�~/���M�,V��LC�Oa�� ���MqK���>��xe��8��F��w_[�T���.Gſ-
b�S�]�pX�	sGm�z�ga%,�>�q�����D��7> >~h]EW�jtKN#�aL�sV�iL�$o��hϝ��5l�wXFek���p0�G��N+^�!��Hõ^��-X7�������%�[��ʸ�����~���6�Mx�}8�9ZZ�e������lN�G�ê��j�;��w=</�W��Ţ�S��V=3��"��!��Yw(b���'y���g���g��¥���n�ދFW���m�+� R��U2�21����Xw4Jw]�oD��=��|���(�"�]%Y��f�S6�׼�qa�/����3is�H)�k�)�r��w�a��9�j��:��T��.��n��9,��{��rm ��p��B��o$��]Q�̽J��H�(gS��!bg�~o�s�YZ�S]�ÕLv�rh�i�`cO꒴�S�j���^w���$旹^�n�u���>�������E�����ƕ^�PeU�G�u�o��:�.mY�{�\�u�oy�8gގ%Gڡɂ���x���x��ts�*05Q!Ŏ�9��3=x�֟{a���<*�]WP �5�v�׼S1������͏��y�Cr�[����[ޑ"BSUr�<�]���B�:]��C^��b#���
��S���[�֨��&.��!t�U%C�v����X\�b���@E�������U�cJ��.����j�%�y�λ���!*tX�T5�lk|�O�P�����P׏8n��sND��`�W�ce>>A1��W��g�V��q��!'�J�|Po�\N|2�X秅
���ܞ��o/�$M[4Ǫ�iJ�h���i�r�Chg�^��I�
�ub��X�jW�k3B�3"bmg���{y�*pR��`��,bq{!�l�\r���T����)<��}�Ǿ�װz��n�
�vLw��r���c����j�a�n]]��ف�7��Ywgv�lΥ��z�OE�᷋՜[tS"���Y�Yq>��Yz�^܉buxX�i�y!/UGJn�݈������o�4����2iB�<xbH�f��{�K)=��I�!�U]�-|�����u-C�y5�9u�UH�T�Z�z-����̮�G1�g�:�X~h�^�m���Ȁ���QN�Z���#|F�p���$�glkC
��*���&�8�_ǰ�hhX�p�*�{�����o��XR�<H
��nn�yc���@=$R�vi5���nK ���x1�*�GEf;�͡��'$���{;�jxɶ���|�g�Ǆ[�ySUxh���ڮ���Tha��oO��=�<���!��ĪE=�b�A"PWKA��p��<����/��p��;�Jy�ҽ�:\7�^(1����L�G3sw�!�R�vz�ΧZVB�y�J�f�r�� �|�D>5���{nd��N�%��6�e���S������SԴ9�k����<\0W���O%��aLW�����]�*�.#H�5�k�k�GZx��\m�d�4��{w�t��Ex���.�sb"�����m�nʨi���uD��)j������K6U��W��!fk���[n��=�tMKVn(*Li�)!���]�9Ҭ�H���λ;(�ՙ�'�X��j-@H��u�ɛb�<x��V_iS�ۜ�qȅ��<��1���F tԝz��Q�,���"�D�7��:�pe<w}J$-��fu[���B�z1�fy�Gy�ַ�FL�n+9񜩩cq֕}�t~�~.��_)��Mvzj��s|��>��QTP����1{�KƧ���T��(aY���\�}^X�o&��������y�*�9jc�G4�v<��MzD��u�=Y���ܶm���k��c�(�����0���QUw�ȼ�[�3�)�,੫\Z��s�	iy��w���|n�J��U��_�KJ#=j�98���������}B��0�2f�\l�*�1���eP�J�
�o��OӴ�n��eo�0�μ{�ݧ�{�c~/J̪�hJ�怊��_B��(lT'4S��bX�k\6���?]JJ�e�̬�R�Pw�e��1\��#̱�bWs@E�����WHx,�������4��͂l(�V�\���f��y}��=��"��7�CҺ�3���D^>6L��k�'<��]�� ���ՅW��2΋߱�<l�(P�1������pWXȡ��!��Kԫ2�/jёPp�F���5��	��6�,�.�v��[ߌ5�3Bu��p����t��#�K��Q�<罃��'����ٯFV����b�ZhfK��>�.Z�Q��T��F]i��h�����y�Vu�X��ݥp9��on����*N\9z�ϸV�U�-b�=m�a���xz�}1x �Z�������w� �Zo٩�<z���ޕc�;Y��Ft�u���e���7�����оq.b�u�����o:gJث�yD�˛�O}��9L�,��SU���ՇB�A��;}F�}�v,z/��RcoUv�}|N�2���}6��C*nw(us֥�z���US0@�w�r�N�YBP�iڦ]�,u{�EsK�݂u�C=����K�r�+d�5c��uq[#ܽ��֗z����Q��IC)kC���;��5��/hs+mG6��B��Z�u��!��n��y��Q��
$Ïǐ\C'W c>�5,�Y񔗢�&�\��ɾ��[�M�\R���	>pЁjJ/��Zj�C���Qe'AW��i�M���3~ƈ-�	BE~���h&��]O�W���Y�R���f���W�{}�r<����9�,%����g�z|��+�K>|*��k�t��Tq@���F3^��i
���Yv<�^��L�l�}�m3x�>�'RC;���,w���6옳^��+����F��PU���z��GZ�6(�[��@������t� ���^�C:��k�{rv��Tp��� fA:�oc]s�M7��M�V¬�z�� ⡾f��l�UG��)�Yk>�!睔�t��}�S���߈b:V�˼U]p-C^~T!�YK���@�6ρ��#��%i��=�F��grўn+Ô�"��1�Ա��[�ޥ�n��o�������ծ鉡Z�t�"v���Z��G��~-�'��3}D����_
�_%c�*��[�V�������qJ �{�=s��$���=�V=�z�� �zw-��\�t�8C����%iyŹ��uܞg�ݻp���jp������p��BZ�wK��S������C�2 ��z;�S���\��B��N��l�Cx���c*��^]Ə�E��e(Wh��6����ٛ���a�>u�[P��@ƚ��P���{�_�j��P��y�	kݘl��/#٭�s3ܓl,��00��N���i�4�ic����<s�������t��C,{�,�Ĩ�OW%��
���k�C(C������1��.ߵ�}���$��BH@��!$ I?�BH@�RB���$�䄐�$�rB���$��!$ I?�BH@�䄐�$�$$�	'HIO��	!I����$�$�	'�!$ I?�	!I�HIO�BH@�rB�d$�	'��PVI��L�r��	�` �������v�}��RB�HD��)IEY�ҨP)[B�T�!V�Q(DUU2J�����!II�R�I�*�(D$U�=b�%�UQHBZh�U!t4��2UD��[t�)*�R�$��T*�
R TɥD@��j�I)$��h+�Һ�(��*�T���"�J���lEJK����B�)@5�Z��%.�v��"�4*����TP�#�S��ES���5I��I&��[�   {�Z�Jdª�6�b� �biEUS&�(��m�*�Ҥ�c �4�f��F���5�i�Х�[mc
V5I`��T���U�   ��U��5�$k`فCa[lm*Q�«UAQ�eH�ڡh����R��46�h���r��q�P)��6SYj�jUTTR�UvĪ$J)�   �5\B�HP�'p P�B����{�(P44(Pw
: Р
7C�P�B�
 �C���
(P�B�
 ���B�
(	�7
C���qb�J�J�L5@l�R����*�A��R�O   Y�j����K�5��+i[T�����\mm٪S���%R�2�J�M�3%���*�,j -���u�
R���C5��F�7]l4EP�RD#mJ�   nv��(T լ
6���JRͩ4՛*���vj-44(�kM��Ui�Y�T�$-i��fР�eL4�ZZ*�J.�(JTRT�ʭ� �^�֐ C05SVّ��Mee4	i�T6ְ�n�R�F��lֺ\R�m�����iIU��t0%P;�ȕ6h*��  1�hhc2V�5Km�Ͳ4T4�h��@ؖ�iZ��#+hMMS0f�T���j�Tf`��m�e�@mi�IIB�ڛ5����R�� �;��Y���V�Y�)Ah� (��@��n%@V�� ̂�*جk@��������M1�N�
v�&��  ;(�2����6��B�L*f�����`AVЕUT֖��UUV!��&)�kM��A�KlV�B!�  �׊P�V�A��P*��� �h1���m�� ����������U�F��֨�4��U���RT�4 bhE=�	)J�  ~�h�d ��JT�� "{Q��T�C 	��M$D�T���a�� Y��q���	�5�\J��&�9�@8�x�8}�/�"LF�w���<����_��$ I>��BC�$�	'���$����$d! ����?��?��3�>��nڬ�I��x',˺ɓ����k:��Be�s��񬬋J��6�gܑ���F۽�~��-KN1H���K�~���;lnO6�슴�ci���$�>4PX�j�c2�	�ʴ��N�U����u�[QSͨt��V4ڪ��Oo576������^��������8��SLM�j��ù��m��+,�8.;���c�QI���tX�]jmi)�ʖt�ݫ�-U�l�w)�h7�2�E���h�,��x0��{&�l�b%����h*v��B�� �- �
�ܧW�-�ʛc;��I;�0ӃT�%��"[�\:ڐ�5�G7���)�[v�X��P�ŭ��S�x��Y�-G3���.���j,ǰ,Tƫυ�64+[��mm\���%eֆ���6Ԧ�/�{�o�	���PuMH]��+�X-�(�ҭm��hk�q⻨n��-j�L�gȶ27hh{K-�B��zl͊�(��L��י�%�B;�KKH�)H��KRwu�^\�-�%�S�S��b��b�[/$�/&%�l�յqQ$�ɱ6̥�S�i��GrԖ��ђT���E=�@�ֆ;H�R�t�bKE�YCt
R���7C��gE[��%�M����^+q v�Э����t����r�F�#V��y�bX�d�ݭyY�8��x��ˊ�וa�'1�k�͇~���w���Y�`�E�[�u`�D�,�	9����O4��%�b���v΃NmK\cf�n-e��e�c��1��c�0;9yG C��n܈`�y��k/d����a�v	�ETz�=8�A���rmz�4z�1��D�8�n(q���TmTڹB�n�*��غI��ݫ��CIɫi�4Y#R��#����Z���,I��(��������mu&�X�X	:;f�1�Y��[T]�Ь��fi۹�#H��kbWt����K������vԫ�J�h���r��B;Wi��۰h[E���
�v�n )'#����e�j���ܖ]bN����X@Ѣ����h������#Ub�a`(Ф�b;mP��y�VQe7XpV��T���$�2�,!$�Nm�[�B�,�˥�&AGc�z͍k[��4S�ǖ%a�G/qՔ���F�t������LOhZs]��0��c���4�Gs[f���4��2k��4�)�.�r��)�2�l2��nᒑ'���仅f���q⧶.* S���O�CV��wB��@ie1Ę��,L�s�:�j��o�U����;�h3v�l:)��A�P*��oc�2����"6�����r�}���X ����p���Q�`j�ݧSV3���@N���m����J��ݘN����Q/--�Ͷ�`R:EV�T�@?Jzov�퓚��Ų��P:��+����P�T�Z�`ġV6�J�\$��'1^�M()2|d��F�Z�6�n��ƕY�uv*c���i��B��[�5`[V5��țM�l|�j�^�iV�O�l����K*n��Q�ӠB�5i����f�)�ٗ{��%����)����F��U��%�)�2��q�F@ng>��Ĵ*^��yZElu){���Hl�L�"���]��0�%O�#�AUlYf�#�bTV���֥zuc��VQ�me���P^i��p�+k%dXܛ`Mme8��DRZHk�	��P�˃^�&6�XYaSY�u�
֣וq�+n;v���d��%��DpҡR��FZ��n7��n�O5�m�l�Ŭa�h�l��3U�xb�4�R�δ�Һ�9�Ȗ5�Ux�d��s ݊�b_g�Ҕof'-SU�76��a���/N�STznQ�WT��W�0Isoc��5f�m$��[�KM�S�ݫ?7��DIU�@��H�*]���Sr&�kQ�#�G%'�gVEZ.2��*y��\X��J:����ZJ��gmЦnb�Qg�	��D^co�y@���zl�ˤ��Ȇa�i+uH3h���4�-&�
���zK
H聍����f��qܩYeG���0�+Yh����Mʴ��t"U�k����b���yiHb���1�Y"�D#(�vҨ������:�]@�*]��,�����H���K��<T�V�J�)ԁ�P+��D��
��f��Pʚa�Om	%V�cV�h���s"�-VX��(Ky�f,��I��ܭڸhQW���B�Ia�4eٔ.�Kar�)�eS�cp��u�0۴��B�&�t�{Pͥ�(�X�P7!��I�F-��H�:��PVG7`,�B�^��6n\�Q��z���aªlܩ���0�Um�-4���Kf�*�%����'C�r�k8�6�{�`��D6�W��m=E̊KXF޴�bP5�����6����Db��U��5�
Q�CDL۰dC���tU�Khe�-U�*k9�Gq��n�2�a��Z�%k���^��-p��@,�t�֠KЍ�a�|���fX�T3��O+n����B��ݑ�;
@-CViAR̡DI/n-t�3��$���U�6�In��A�Z�|!�@�m��-�q��)1�.�[λ��:�{t�[�jiU�d��r�t�꒯J���&��|ݎ`|%�2Z����ś�;�L��gc-��X�jRqia;��M��r��a���#K`�E��n`�6쓒�c�N�jӌۈ��b�]æ;o��&�}[QqY9Y&��ɿa�m^�74�1ڼ��ֳGIR٣*<���D,2�D�Vرj�T^�5��ǹf֚JR[z�*�x#B34=�PKW[�nZ����qK��+�N���׎�Ҁ$��Y�D�naFdm*MdV���U�����؈z����v���ph���n,;�aD65����5��͔��$�I�M�ws+^�����n��iRQ]L��HUY�{�B� �W���1)f�(e
HMX[;n�[Եǲ�å��<�r"ި��q�����t]��u�
7(Lt�BMS 'fۺuz0�d6��ZyKq���,X"j��c�c��P��(|*;R�cX�
�)�c�YW�B;��v�S���4E�vp�Ϧ�ƥ�qGhiC��oh��vku]f��5��v�-�7���f:�W(�N�bkk �e�[b�j�)�f͈���U��|/n?,z%�e�we]"�%G�Չ)�2-�^�$�e�:i;�j����v��Wfh&����o(^6N���u�$k,�V�n�u�M�C�5�q��m;�+^3fձ���˳Qڷ���eI�`�r��q��Hˤ��v�[X��V�;y��o�#�+)��p�J�Yv�[{6dCj%�@�ͭ�5бxo���	g"�ZS�ܩ�E�erf,��^��^�"ʗf�L`&�;���]�˶75�*��n��+����*{t���[;�A�6㥙"n�6���a��[�h6Y�H�썬�
o�q]�@����ʹ�4��*"����Iha^V�L��ёx�S�0�i���?����l��mFde`����	+��v'��D�ib�����`�ZV(~d�6#�Xk�knɑH��J9w�`]Q�H�e(���Q�,/��H��{�N��Q��3J���c�v�1xS��A9�CMk1e�Ci�SMMɻ/m��eʸn�A�M�1�0��sj�B��Z��tvQm�ݻ�Sq�K�̀(��'�*[шj/U+�r;���x��H;w-'�^��+d��2Y��q���m��J��6��w��PyH��j��܍e�Ҏ��&�+����n�'0��6�o��)Ggn4���ѷWL�� 7�Y�ְ�I���ҖCh'gkB'*�S�`)!�7]�"ƙ.��6�q�AX���!ڱ�c#�TU��7R2��e^1T�tR�LI!�0f�YY-�1�Y�'Yb�/yf�q�\^`�+wl1h�֦k��ǧi���U�nXab5�uc[AL:4ݫ�q�cfnjh8"���׊�!�K��źT��Wt�tL���ϯj��y�=�i��[50��b��$ܻ��ʵ�o&�5�l�hV˽a����"y�w�f7ZP�U��k�ej������C캳z@�h�c�f��NK��ux�U��~�UN�u{���9(Ô���nD�e�Y�Z76�̎6�[��&�)کE�t6�'�-��л�r�\YM2��S�f�^�UD�ɔ~�yh�[f3=9h��:B�����*<���͡F=x��[j��D�%P��mu��-:����a�%�6VdU���V����o*j��eV��2CXׅ��Ρ��h6c:���E��n�R��-Mգ���L�`m�tNjckbj�𜴭1�-���m1
�
�MtDL^�1��4x�r�ɣ,�kub�)���h��ã�<4]�'.��7X�l�ܕ�]��b�"��"�F�pl�@WvOU��Y	�;��ԣ�3&4n�ݫ�^�����sRG��K�d�uQ���)�gv7r.![����Ex�,��m�̴cU��.�����-d��V���:W�e�f9n@���ґ�$]l�ԛŲ��x2��T�T7�e��$�6�J�2��y���*6�
�aB���n�b"���Lԗr��]$I%-�Y����*4�m��!H�0峂b�t"�S6�x#Ϧ^� �vh�i] F��9�M�ܧ�^ՂVG��{�
�-�ܹH-�æ�Z�مf<*"�Wʴ�'7zou �h�t�p��J[&0x[�F�\)�A*"�r�ݡ�CX�xq�[Ք��C��J�7B��ܕ�������m��z^]��P�Mֶkvť ������P�ъ�K x<[o����!E�BY8Dyd� 0��4Ց2:�k�j��"�7�e�s)����cUcͳ3�ř�[���ɫEeY��;9pQ�#�^-�A©B�+��l��xAW�� Z{����xBJ�ݩX/3�I��L<0���Z�
�G+b 1ԡz�Â�jrܙ.�:��cp:�A	�c����`�Jʈ�	і�<�_�C�=��C1��Z��b]�㨍����N䗩�f�Y
���>V��́@�J����Rn僓YZsJĔJ���d[/	���t�th��2�OD��۫[�1T@������$U�2-���c ��nЫH��ݣ�2LÚ��n���-�7Q)��pm�B
����Nm(+P���[�n��ѵ�!����YI��3 m�3B4��䔆S+.�Taz�7W�jזR�[b\�j�f��Q\**��Vҫ	���6RYe��A�n���e��Bjm�x�-d�0��9��vI�vbҋ�E��ȥ��]2M2F�۫���.��֖��蚻�����"�e��т��Ʒ�V�9a�C�1�2�墥n���)@��=ۥP�B���X���V4�-���7v���jj��@4
u
)�i��iǰ�\'j҆ڻ�kkQ�X�ڻ(�*e����؂8s����N�[�^R#N�ƶʃGQMJ4�ȱkb��X@^d��S����3t��zT�KqϘۦm�>L�k6�Xp��{P��ް�Ch�m��.���ۣCde�/ �iQ2�QO
u�����)��:�.RTlR[S]��4����N�@�ֺ�@PKq�&�8�n
�t�N�ƨ1�8���=�+`�XJ4�9H=T4`.4�ql�Va�rD�����L��A��@
T6`ʕa�Z&�X��滭��*Z��%���-\�Z�E���4&ƣ�j8ܰS�YW"��9*�+Bu�$�fį�4�;�Ir�* �Kh�nZ*��
�##vأ�ڬ�)?�n<�	l�M�'�	?�6C+����{���E(�e�H�YcV�']�t b�,#�m��B7k(�ˏ>�*-�rM���`Ӎ;6�ĄjM�{�v]�V7`�;�H��,״���V�Kv�Ej������r���V��ŔC���a ���0�zE�W�n�Nne��nF�nb�����FR�q7*l�1ˤ
��VAV�<Z	7���H56�^LYWn�E��Qb7�,�Lbyn�hfm��w#hk�0�WYP	�ѭwH�O�J�z�o>{�+F�j�
�(�x�s\m免��t�h}��H9�ͻ7A,ݬR�5	���Q$^ے��j4t`L��@�lTA%��������u�T��P]��~t/�goBT��d�����^R7u)�9b�x-�`�Ue۫R�ڶ@�E
�t�H�Ҭ%����c�0\�u��]Ֆ�� Jpn��V0nŐ ���V�5��/��2�LCtS8V�{5���hM-��34+�vt�e�600��M�C5�)
Ra[4��hޟ�7h�!r֔���'�oҝˬ�(CCiPW�!�4�&v��׏ t��{R��0�U,��`�����K�N�����c�٠V1-��l_J�WN��͆�Aw��f���٬�B=tu嚌���)��e)��+�m9���GowS6�[�̎�ۘ�hFP��xC�uLR�mR�Wg1�c�6�
F�H[��階dbt�:qjե
�4BqL΢e�OZgw=nj���a�wuc]��ۊ��hH���	ݬ��ō;��6�̫ ���d�[��[W��0ͫ�۬�t��)��Vj�H4<Q�x5��6�P���P׽���٨͑/-�!n�� #��5Kt�F��m�K� *�4�@�Ѻ��ĨVZ�bW,�32#YxV��w#�M)������$nSquy�ed��5#,鿕�c	�	5(�e꧗�R�8���\�u	+��%m���;�,�˺��4����[K4� �53jr�A��>����\��81���;�KnY�wÒߋ7�[�[�;
Ф��vT����B2:�)�&�V��!3��dw]�_�����Y�aSB4v�ud�����z5�D+\ﾴ޴�,1��U��ۂ�Pv ���K����u}�岟i��HQ��i�A�=���Mh���C�1o:���w��oʈ]3F�k�&!�W�X��,��7��c�
��^;����γ9�Q���R�5G`a}]�X	-����>ǆ�W[ ڸ�����-�1 F�Դ��eW�u^a�u��c�;�wW��+K휞u�}&��%G:>�Ʈ;��;a�ħ�'m��Vo!*q��uvsS8e�[�N���Z�_�)��Dh����T�M��K1��{�~��w)�~7�;^^�D���^��
�.<4b&�R�9�+�D)+����-��T�*��n�6�����X�������;���zp���il�yf��_K7)<����a[Fn�R�!�m���fU��Ms�ʛ����u$��z��K���Y*�|U�o3��S�*ܲ�J˾��E��9��R]��zX�8���=m�쾦��x�YX�ΥC�����FU������c�[R!sm�eN��k��f��ŉw��tgv|�a�q��1��)�rr�k��'��K��;�7�{�|���k�EwsOpٕ;������]�Bc-}�Ocqt/�j���]���S�lVM8��鵒ի���ε܎�U5�WN���&�۽ʀ;Z�5��.��v�w�x�/zW�MӚ�
�
8uݽᗂB�s/�������E�l��9JX���Sh�u�I�*�[.�e��hc9��%-W;�J�+[�� ����	���;6��GrUι�9�er[t�ia�#�v��g�����{��x�ι|��D��1�U����T�u�SV��^7��I��=���9L)Q2{��,���l	H�Z���sڱ�=ˮ؛2�skN���*3{*T�[	D��G8.0@ϭӎ�(����\��$��*<C6����͸�V��aBt�Q�aQ�z�5J�m����4,:̤�^��]Ζ���._�}L�y�����C7ǫw�o7;�RAV�WV���t���P�JS �)��s0V�;���r8}�ȩ0!�B�[��D�3���-*�I��2"cL�7uU�ՃfS�M[��	�]QcݔYn1�O�N��]�g�s��y/��	ot�k�r��S���e��V�Q"��2�8�떴�X�l���T��=����әyL>��s;ce�j�Z{�J}�nr��jGe>����gݬM�;�	]���{W���TS���p�u���m���J�<���=�H�D���ө��Wz�ј����	f��⚶�� �������=���/�(�t���f�um$���}�)��s�W�a;�;ɬ�m��'�*m}�%���wB7�r�M7��d�y{M�)B,�)D'Kabt<�[��
�m�i�]��*5gT�=}"��Jn:z�n�*Ȏ$Į�N����/��5ooK[�b9c�>P-'8���я��e:8��������rN{O���z ;�v1i��g,�4��k�4� ��3�&�g*��fî�h��y�w&F��W;7����-ٛ�5�\�Q|lR��կm�]ź޷�$_
H�F����"̡Ww]�*����폒\���Tr����q�s���<���z�,���.����A����q��x�Ǩ���:kK�۲bY&L�X�k�H���9��(E�A�3	q�k���e�����M=Q�W�V.��A��y���+J�;�/_o4�����:�i�5ضt{f��4��i�pw7gE	(˷uB+����Ř���U�;{��Z��6�n��2)xr<���H��z>�j%�LY�j�!5�U:ҋ\�g/T�Z�s��-ۜ��h`Gw��Z�i�è_η��nC����ĥu�+�<�nuG�Q���s���f\��VY�.�M��tM�k2�m��͸9���	�K�RO_WG�A��t3&;��s�eo'W|�}�.���.#�7N��GB��%�Z안�
Gt\�q��F���r���KMf5���j��d�Vz�J�5Ⱦ��C2�lK)_tXdʵZmLJ9�u���+UoV����*�G}1jh���h:f�im��j�3��[�)�8���vS�r<�AM8�,,�:��qt�kH�{��QS�*�k�NUՍZ�h@���h��'���sb츣|,un�	6����u9���v齅�m��%����åF�����L7��ͮ����1�� �l_V.���4T�$�0�+�G�EtA �v���c�f�J�ůJ7-��ܖd� �[{M*���[��e�`�f�t����6�8�����i3����3�od�l=�Wؕpj*4���WZ��[�o��AY���W@{^�v9�#�u�`��'=lm�|i��:��W&���/u5�kH��y��T�����Eɉe�p�)N��4�$
������v!Փ�,��J�Z�L���u�u�ԭWQ��G5ۇ:�4��mQm�j?t�J�љ���SӲ��XIjݬ}V%�LeXM�\OVm�Ѭ9�J��kC��{)�T�v0G׋ISM�X���Wc�����C�e���-��S͓/co���#j��p�Vv�G5�U��.]�j�G�]%�'F鱼�z��!y#}8%�}z
�����;2IdhX{)�R�Oju��n�ݵC0�]�`�3: 
u��ufT��j�*6*�73s,�`�d�x��Z뵖���utc�[��퓸��{Q(�uw�Sn`Pk4�D&��h���5Lզ�3.����sB�D�����m.�v@�w�����_C!�F\��hf蝰��9����F�f�s�un��(Q�Ңi�uѢ��ޙ�vi�֕N5�x�*oc���s ҅�K-n���{���S��-c�Vd���Ν�����N����ӂ��Qh]{7�M�g�a�	�d}�wZ�����Үr�U��&Q�p�(jq����Wl[ˎu�Ow�rۧ|r�WR�\�I ��=hWae�I�vf:�g0�漿�P�����M�Rh�ZH��ty@)s�r�#Gl���[����.�S����P�nC��N�EJķ�$2������K7Y�艄��B�&;w!|2���_[��)d@h�Ə`�J��/s;�[�y���wµ�UcP�o���e�zL7T�{�:m=�<��0Q뱘�eȡ6���,�q��xV!z�R�U-.�9�ג��݉�c��=������ĝ���*N�"�(8��Q�
�]�Yw;�̼`�SS�J��-)-��F�vY»o&�P5:�㭼N�U���n\*��U�����\���EFB�|���&p ^V�e����R�w����Q�t���o>)���H 5�jl���^��\:��7�h7Jbח���V�t��ּ��r\��*�Ve5Kj��ƅ�]�*�]�����gxN�_v^�����$Q���48��Zv�
���
��_W>Žj&�.ҷ	{�f女2�8��ō�4ay���.W6�X���띆jc�.<I�䨼SRo��^]���9��Ӌ��2�Za�p[�0m˵����s1d�=�k��
�E|])l�X7���w�6�4.ͦ�T+��_z��"�fn,����9�T��B�k'mk̡��©�4���S)��"�JYszbu�#v�T{d�p�]��u��ΨUp�����������3���u�NT�Ŋ���є�Ƌ"�wX!޼�]�K�*MqW��qu�p�\�g.�L�@�Ţ�l�TZ���%<8�'ٸA����_-4�G�#|([ԶcY���bt��9F	Z�"�Nw_v*�W��G�F�K�F"��c}�=et�l5�.�za6�ћ�sZ�:v��yr�œ�<����*v �����`yKO��^����p�d��w���g��C������5a+�J�[�֤�H܃l�D��\=S2�ײ��ŻM�c�D�kr��ҙ]�=�TkcoP;��.����A1V��>j*]%���q��'���}:�Aoh��C���@<�C�������A���� �,F���:�k���u��N� .62�ln�^"C8�or�@a�
z�� �,�΀*�'[��h;S�
zo�s��-|�肬]񽓕饳���d��'P�Co��f��R�bT�}|��ѭ�v���h�{J�#p�%e��Yh^���X�`�i�)@��lb&@"�V��ϻm��X)��%n��S6TשѠ�1�����uf���܃ѤJ4e�Ci�]R1˛4�w.���bq�!��^E�n#�%]
�`U�;9��oն��|�bg�YՀ�ٖʼ�ף-�Qˈ������N͢c�n��B�V�CP��8��tSӴ�V�]2=�IF���n%SC�&5K����.�D�Ehz�i���A��n���:��sR��Z�^uA�m6g�W�֝��_v���9�	��|4��ӏ��$��L�k�Y���MG\�����g8��&��)��R�Xt��\5w�������ۻ����cRЩ&�P��<=�޷��i�X�U(�T�i��v�Ok5+R���a��q�nZF�^�d�F!��Tp����³j��t��;�Ev��1�Y�Q�wQ����Dq�}v� �����ڡ�t���miؑ2�����5��[i����F�F)EL�x;����M:(Ngn�,)�GFl*��k�Ǜ�a�Wmǻz�����+{P�Ȱ�
��[RhdG�ڻ�ke����������(t�Ճt*t:�Y+�<�
��<�Z8_YB
3�#1:�+�["���
�iT������x�tW	�:_�f�������s���Q����2�T�0I�HZ�^J�Ȉ�.�i��:u�{fM�]9�1�R�v��U�D�I�u#�,B���(�p�'�=���!}6n! *b�]��)���R2�,���}xY� ��L6LOs�
T�0�HT��.��y2�ͧ�w�uB��V��f�rժ�]�`"^c+	e=��j�U�Fm���T\{l#�:�c'���1��]�L��|���8�ֹ���Ų�t��o]ұ�i��"��9+ �r�M���et�ڴ�p7���Tק�� ��eη���r��Ign�476ޝ�/6o���ߝm^+9M��)���CEZ�e�N�V0Fӛ��.�;qwj�ީ�KF)ee8�<�N�̙���[˖���\�sT��h�҇7p�A�4�^ݮ�`Il�����ۉ�:�W�}��Lʴ���
47���,�ݭ���Ō�ӛ��P���E�o���)6hk"��L�0��x]=|�7.Fl7>�a�3���V�,�_���$o�ͭ䮡99<�\x{��SV�����:�����m�FS���	�$]G��
9BR�CN�*Y,���yz0ظ;�R���b���\'����w	��vNUC�*6%�gD��~�L����.�3x��;����o�7�
QΫ'����G$5��əq�;����7;:�n�N�ϕ�|���<musn�y�}���J�����8n^v�� ���o%Wo�.�e���,��W=@e]0�(�bv�1�v= �#R z��˳Z:���G��	n�w7��Һm/�ω�F�^ik������Kh%�յl�
���:�'��c8�[�Q:��1�L����v�gs�-v�d��s�ڪ�z�2t��wS�(�*����C��N��S����gpsC�pM\�D�q'K�f=j����Q�tީۜ�U��:`mf�n3Wt�9Z�*`Uɣ�2��˓��^Th�}Ů<���L�KD��w�{��)���n�f �`ȸ��)�-�,�Zqk҈P���eɍ&�+�����Y5G�tU��+��G39�ui�y�9(ڨ�[cW×L5=�n˗�؂�w[��nE`�B����33��w��CT�Xg�\dsm��Z����Wp����9t�(�_!+��Yk�\��KWYZ͠�2� ��N����HMD̮���X�_QM^Wl�n�����r���:�1 ���8�\��*�4ob��r���)So��xb�=KY�$��
�V�yg��Y��"�z�6�i�yV��L\�q�ɶ⾕���y�K�U��eu
K����.����X"a�̦����i���J�:<q�\[�Am�#Λk*�`X�ǽS�����N�wF�2i�����e�6L}���5��9���k�8���V^�2��<���]�+%��Y�i�[J��c[�u�]#O.:o5�ov^�x�YI�BY�{0��G����{����r���(��+Y_�(�z�7�mb��Kuy��u)[��,�:jеp���F��9��\b�Wif�'K����a�p�t���,���nIѺ��Ԏo,�SYKf�'7f�0	�ue"QL�;��|7:g�%���{�L.�� ��:�RZw �e���Za�����_KW�1�AIdZc:\�L,��ok0�	�T����R�k�L����y�C�}
���(�p�X�V�N@�n`v/� �"�"����E�ylB,��f��K]{v1�ln#���N�2�a��a�}G�:o8ʥ�I���re�xG>I-��������W\����T2�0l��I�'&ƾ�NEӰ��|�#�v�[8tد��SԲi���r����F_a�wӖW2���NT��60�|��u]r}���6e&D�f�(��uX�RwU�j����>_~ӿ�}��@$$?���$�;��&hs&���XOꉉ.�Xp����w�=!�3�*f��(��h��"�c�/��\�T�6�vY �jB!�ZW��fs4^p	$�Aۘv�J'��EYݴxu��l8�Cz�1��rovԽ��K�������c` uܘ;�˄�*��G�e��ҕ���VZ�C-L=,��W�K-���v�:S�df���AiP6��c���d[E%���ͳ��F���SU#�x�<����+f�J,upތر�2�y�4�-��#r�j���V�f����Z�(��XB���a�+�X��pt5���B�r�c�gA��vi�m,h���Z [\�JW�mi�q�j��l�x��ebVn�V���Q�;J����{��:Yf�P�f�kn�u�y���J�p����"�&a��gm�S7i �0\�(�]iヾD�i� v�\�F�v)B��4��D1뻰�M8�9��/�wi+��Ww�+��Н]�N��M=}qM���VX�l���ݮ��	;\3�z��:ÈCWd��T���L��^%Ӿ���}`�WX��+:ͧ���Sx��e��g�KN-u#��F��`o.��os�Ĭ��p9-{%�g̫]�� �د����cy�����FbZ{y�45�2v�N:��̂]���"��׊e�cfNͻ�W+ռ�^���h�,PI-���I�ˑ���Q��n1jnQ���l��wc�vP\>�^da^1W$[�SSv��Y@5![���며F˚�ț�EF�nm'O��3�&�u.����Y���ʰ�r��Vw.�H$/5j��QQ��w�$���|����[�D֑�`�\L���ïc��w՘��1��.�6n���*W4(oe�8t���<�n�]����
�%�(q����r�J�)��o}�j�Sv��x�;�8W�0��1u��u�'��2���ޒ�}���U`��V;9�hhIb�����j��e��l���V�q�($��y�&f�Wޣ��3�+��ΝӋ�J��KK]k{䚳V'��d���M9S&ͷ�%���A�I���ߔ͛�� T�t����,��-h�5Ds��K��9\���t6�>t6�c�᧼�>;�mn�%��}��X��Zq �jr�y:e���7펍+2Û�����ͬ*U�km%�k�OF��t��q��0��tp�T����m�%=����k�j5���)ZK� �צrhh�;"���T��v�'`a���ۻC�����ڻu���M���K�����2�_P��u�G�0e�g8J������"�k��������gNaZ�{�	�{�f4�u�oLR�<}7���q#"�v�fb�N����v���X��J��!d�.����
L��<ǜ�\�-�X�N=�2�]9���&�3<������E844�L�ھJ���:4���9�w|�P�pH�:��M�+=�G#W�/^���՛k�c	�m�6��N�˔b���Bq�a��`��RK��#��Nt#sk]pʾW
����{�SMX+qq�ծ�+�,}d����v�z�k�)�M�;Q���i�uvڎ_Vu���,�����v&����u�%��s5&iY�&���\3M#�%��$���e��f"Mw-�Խ1JZ�e��:O4�#5�n�ۤ!���6���R�U��j��1�&E���t��+�6��RR�7��w:�+؅0�͛|�j�LN�*u��O��]R0\�֦'U�� kfW.O�Z�(gfL��w^�*.�\�ŉ�Ӛj���j�,�Ĥ�#$�F؋B�K��a��wT3h�]�[�j�m���w;�|m�����d�[ɸ:�o��OM��!#f�=D>��*������yC 
�*�W@�r�,�6��%���Ϯ�n�A2`�2��y�=taT��¡�����7�I��.7z,z6��j��ې�v�+]Z�쫹>;��m�->�Se��y$:n�Q&���c�_:�� U[�;���='�0��cTb�R)�lu��_
κ�����֐��^��$�Ә��-������.J%�\�wZ�H�������	�4�x�iռ�����kZ�(��[| X2��ڭ�&��Z�Ѿ���5J�=[V#ƅ��7�T5M7ڠ�݆Ր^S�狸�:ȴ1�՘��s�#�wRZ���Y��7إ���i3�Hռ\�;4j1����(��/r�=V���X��nI{\��t:����1��n�u;ʜW�71*OL��t��
_M[|�5ǰ�r�m]�v�ɘ+`��YVC��x��u�d�Y�o���]��{Ud�񽭮U]�tЏ!�v���7�d3�϶�\��F�ֆ1�դ���t�d�%�K㽋����갥�Q
�mkS$�]N����Ƹu���Xh�-Hu�؊�\-ZƊ�\o��+��@7�.�A/i���=K��(,���&��&�wqnVنSX�����,�@���X	
I�MK	W�f��D�N��@�f�`��H�LY�5�c׊oE�7Yդ��0Rӕ|#��t���+��Ɯ��bV,hrt�y��&��x&kr{�Ve��E�p���ؙ`��n(�^�N9F{�V]��r�O�;ҹ���Z�x��/�G������V�#ao@�s	�Oq�k����B�ܶ�|2����]�5x��v)�e���ؐ2e��zʡ�	E@���<=jR�R����r!�von�N:�I���]��6���Sw-��u�j�wc���Zi[v�ݺ-�K$��avɹ�`�ig^�b�&�l��i��;���]k�m8��v��%E�7��Pͻ���������n��Z���Yd{5c�gex��\�'2*�V� �H�ؖ�u�&Q.�rueX릭Jֲjv��ރ�*{t�dKE�r)��d�2�
��84i�6m�#*^�� �=*�r��F��
���+iZ�pY�wu��-����uؕx�d*D�Qͥ{�0�}��ŤZ��[�j5b��I�&V���D�U�]I�0`�DQ[ӫ�(�휺s*�%��
ҫN�3��֙ڈ�T�b�������{֮ �4�G����pf���1�[k&��]]���b)�k�e���|ɭV��sҭ�W�8��T�\�fl/��}��QS�꩙)N�]ڻ�c��\���e��n�63z�l�A,�����C;��8�;��\�9`W$��kO��$��J��p�8s���]�N�;"��gb�;W�����nu'���F��Υ�v�]MU�#�\�*TE�^���'h�͝r�kpV�w+]��V�1QQ�Hщފ@�or)]j����su�9���qe�f���wvD�V*��lR�h��e�S;w��>e��ώ�ٗz�O)�)./�@�!\�鏤��];e^s��*��:Ej��n�Y���ʙS��k�A[:�U���*U�NU�7��1���KԸl��;z�_g�%��:�-e<th�Y��\�&r�m��5nČ����s{�ąDYL�8���R�X��W|7��i㣚����jkW2��� X�b���Y\n8�����H�v ~|6��07�k/P�4�2n�H���*E�M*��R����c�9����/����)��|�
�L,�g�i������1��a����L"Sc���K�YN�����5�t�����1�H��BL�[L�ȭu%̾G,٦u���l7�7�3�u��v&�_F��[#���^�쑎N�m�|�{F�}Ɠ�:.N�1B��=C���D�_sއO5)�籪�}WW+Tn�����X���,z�[�]������i��i
�ř�2�����
��t�	��ob��K�_\�2g)�N�m^
i�AJtsc�+(4FXs��[���d���/�`޾���1+�:�
AZ[�euc���4���7��X�o/�]�/��d�(�P�4q�tm�Xh�t{�G�N� ��۹�Ut1�a4-�47�t�k�n�\�I�jܾsf޾���+V_^ �V���]�cW`z�RlЫ7u$�y��傐ɦR7Sc�3
�{�r䯍��&6D:�A%TaY�Ga�e�pV��5:4Rb��1]d`�	�mQ��\2���;O��u&]�^�7{VX��6�\���@�	qF�du�.3�hA95V�ݮ�,N����5|�o��%��L�� �������8v�m�Sko1Vd�4R�Vn�L��j�bW�xi\�sr��B!6v��*��Zgv��)�X��`+w�HQ�N˅��(A$�N[={�NJ�8er��f�3)v�jޡ���W�#J7 ���>�.��RD��:o���A5��޶��8�U9�]X.��&n��*�ͺ�\C��@��.�aptx�|�5�I�t��o�ǒ���#4�x-�J=�ʕYr��ʲ�fX���g��aS������r͌t�q��3
�{F�k��>���"U^���"�m����`���*ˣl"�aŵx����`sf[���00+h���E]�nWM��
�:�϶�����$h�!Gu�Y@��t�]��d��gbx�Ѡ����Ѿ=oj+9�Z�d�ӕ�<�OI��ڵy���2�▮%�O���a���!J�|�u�����C�m��Z���;En����br���Z&�<�k��۷�5yh��9�JH��"D� �۽��7��Qm���5*�]�s���V-�Z*Ue��:�:���Κ��j��Ⱥ�x��7���\�=�1���}ȴr��a��q��k�v^�YF��)�T�;!c:�V.�C�ᚉ�����H��J�c	���X��_��&f_�}�0�Ȟ�xn�O�+�5XV�
����,ig���v�m���f�R}فv�ɮf�`D��F�ҫ�vô������M�QI�\�<2��n�ط,>�XR�n�jոJ�@���!�+���'�N;�"Lm֭em��KU�l��N�?���mm���].�"��CE=k�C�����t�:�pp���*����n�c��W��T)֫�9�-�t�7o#�;kZ8�]G�̽o^����LU�ά<T��p&a��ke��@���� �F�jnVi�u����Z:-\�7u�bӪ�)I�]C���t�����w��6�=(�]]6]��&n6{.
�OF]�
�o9�%��͊�=�!t!��9GMP�9�RfQňG���u̓!�:��0�!��ˁU�x{WGj��XY� /S�c��**<�r�+�[��zU�� A�(��%K׈���
����p,�F��Ҷ����SU��ib�y�YJK���b�t��,��9��I�[*!��v�3�u�N>0�-�I\cư���6%9�7"Ɲ+�t�x9�mb��ۺ��4�V�I��sim-L���+����u��7+����pm�lV�,�����MjB��f�g�|���j%��4ah6]�vd1�:���������S�,�b`k�#i�Z�ư�[H�v�q,�Y�����$��wh)���nǻW
�L�=k�:��̩p�-�i\4����B,I��{q�ɓ��!�F�����oe9;��ԫ)+bb��R8f͡��69�]Z��	�Fm�ૢ�|��l4*ުޜEW���u��F�>�=���nY.�:t|��o q���m�Jb�.\_Ao!ƶaM��]p,�Z\�U(�ckK+^�Sv骍>�m�Sb�6�w,������Ք�5eA� \���:%�U8$����4t��^�"qK|n*`=��{��7��Q3��F��Av$����A�#r�)��ȳfb�+q�J������	N���٫�����^l���P���]�ڴEi3����[�o�c�.(�ڥn� �aru����E��/^UC�.�ZLBl黦:��<���}K��\�U���JE7����5FKV�4{DV-7���M�H�C��7CC�9�1P�&�Su{x;2�<Z��"ŵ��965�S0�~Iao����rAk��cZ���@=m� ��K��\��r����P쨟bO��j��3b8��HN���.��A�p��]4�g�m\�N�Y���ܒ\�aۮ�%=�蝷����̬m�&f�n!F�s�^;��+]v�q3�MY�wPdNuZ����ڙVP*w*Q��Gu4��WL�!��z\MŭR�������(-�s�� �6u�{�]�Qov�����z.�̛C;u%QN�!��NwG��y�Dް�x�u��>J�6i�ۊ�0p��A�]�q�Κa���u&q�*�.7�e!X��z5_$���=�]�q��J�[�A��5�s'`�6-�6c9ZW6
��͑9J���u�(Y��!pF�e�l� �8 �đ(i��Xk��L���$�\bD�����^eXQm�M^�R��x����gmRji��2�-4�7��mk���5��T��k�6477�.�\���Q򗂈u �*u�Coq�{��S�݈��r��̣n�t�Z�d*��k'��wJ�Ŋ�r�Չ�"3U^���j�, (���6�Tz\75YQ�w�d��!}3�jĨIaX7����y�!�҆�hm�Z{�e��t��K7���N�����vo�i��=���@����oU�N�,��$����k6.Q���+�T�bԸ�w~�4�n�&���:K�u�X�nQ5m:�9�ef�#q�ܮ
�K[D*��SYW�`긷�ܺ��.����ʸ�[ՙ��$�O_u�"zAK;�09�?{��]j��ۯO���$���u�X������ ���vi��#�^ui��
�A[y���Z��g�-�,̇<YD��/�ۍe\�R�*̇uC�֋��q�{��8��0%�F�c�\�0_u2�4���L��V�ތ�����]J�B)W���E���x���gc��&JW]w�l��|%
�d;do�Q��ǩ5�/�6�y�_K'e�ә���# �#��ctN��&we�Ƿ��{C�����4ث(!�3}�*=k!bfJ�8�/�������Nk�b�ʜc��t�Th�'z�)�6b"�� }o%n������Eeg�܁��!�|�7�����l�`��gi��Y�֩����6���vU����̀_J��|N�<�]�3vT��X��!B����d:��M�w�c]�ڦ=6��/�AA�V�j���C��d]��]5d���!NZe#o�Q��D��;�7Z2�Lvk�T��K�5��a����S��c͡ǻ�yn�*�]��iZ L��#%,[��O�_X8pn�{�f1�M�JD�����pewv^�mT�@Gup�ڕA_*ע>�F��FA*��]wy���¬�0�M-P̙3U�����|��$��\����uEe}�q,��2P����)i'�f��t&�*��:�nF�o 
�\E���S�'ܻbs���(Z�j��)�:;WL�Q����7�A�]ե1`h��9�;�34P���͚�A�4��9_2@:�`���(!�p(V����QKv��e�Wۺܷӛyp(�ǳ[{����Ia BH)Uk��Z��m�X��(�jب�m�������Tm��DV2�,`��TKm(T�(�A�Z�D�-�"�Ec(�mlA-,Q��ZV�-���X� ��X֨%V�DUD��*�D�V э� �1DA�V�1EQDQEjX�V(����`�#R��P�++QcX+""	R��� ��EQF#hUb��h6V�0�T�"�V ����QV+l����QH�Db��"1e��R#
�E�
	mDH����2�"�(�ADV"�Q�b������Q��Kd��)iIm+#AR�*����J��lPQa�����PbV,�cTm�F�R(�b+�b�Ŋ�((�*��TDH���U�U�+*���UQV0UEX��+ekDb*
*E�
ER
�Z���"��T�*�����R(��XQQH��"Z�UA�QUbԭJ��[DQPH>$�D�.S�yWV�Fp]��:$�}k2�Qε�x��������Qp��Nx{�)��V�`�N��mͧ�|]�ΦAr {� =�]"�r.�j͠E�]�ͻ(��޾��;���#.��;~�s��9���c@�ɳ�����w�J��+���_���عr�ۡ!�7{eN�{Aр~�u���V�p	n:Y擠{v���usbk6�U[�T��+qJ[�ʣE�#Z��U�W,�t�����|h�+B�op�K��^}��x�@��ǙI�Y�q��P|��C�.��Ukz[�ʚ�.��bus�>O�~��>�EP8���Ԏ�˒�w������i@Нn���O-�sR�;,B��B�^�1Z�D�M��7�
�/[j�ݱ!�CE��-�߇E'm��ju�u���r���5E֭{c�~O���=���Ġ��T���5	�tR��ׂs�
���І=�wg�7�iwrh\��ld�]�w��.E/eR�:����^��[A�K�%�8ܚ	��ՇY���{g�1-�޵~t�ش]g�*kRcO	�{�Ҋ\Q8u#z��.��+��K4�م�K�|�x�^]j�Y��r���f��l�gOذ6�J���E���/��}�m�����iӧ���<I�c��;����^eگq���;��`�*�%8VxcuW3oin��g���O��te���7��Ckz���&��&k�vL�u����*���÷v��.�V�7LZ�e�=-��ny�[��6��(��#*�N�o<�7��.�N��N��L�NkJ�vy��*�6����������d�f�*���̔<ܽΈ��V��,)��z�3�MQ�\��~k*\�W.�A��M�ۖ��J|�3�H�Q�/Eh������Wk�13���vi^�ȸ��ڭ5���N�y��7��ۊO(tr��-P��z����4TUU���HLN=+OD�����[���O�O,Z8lWG"6��*���'7�)��8��_n��S���|��y=�/�?)�E'�7eF����iZ��JU����b$v;��+���oqڹ�iӊ��6�!�@�9�07G��²Mݖz��W@$����}�9�pq+�Ys���gf+ےe��D�렸�{�W[�z/��,,�
56L,��*�ߺ�r�T`4ܷ4�����jܳLܲ
�QN՛��2k�|�
�HWy��n��U�wH��!F��	5ܱ]_�G�jĻr��R_Zz5��ޛOU��']��dj�QT*әmMd�;`�P{�xk���^���tl���j���b�����1��$���x߰��s��h�]�w�-/v��c
&a�]�<Quk{R��Vk��X���j��G]���{Y�'ɭnuU�n�f.u�����[�0�E&5:8��h��5��t���R���}��*V�Tq��e��\B�[��!���T�����sY'շ�;�#)�����Ϊ�ׄj�r��oVx������j��	H�;�t�"��r�����͛�o�5P5y^�)��"��i��H-��Q�{/w�<���݈Iv�
�t���vx[�\�.7���Nv�\�U�Ҫ�[~[�5��`�U�3�j[��`s:T�8��#vzNB�U���K�i�x��No>�U�`'����&��]��vM� ���g�Y+[��b���4�H�r�������
{v�h�X�b���d��6z�4�����v���N�u5:h�\�J�R�B3�c;\.��oN�N�*邱cZ�]��Tj��1;x���7:U��.RU�B[Y��S�LH��R�L���Lt:��]㼨p��&��\��/�+���9�1�����
�L[�n�����[Ns��,ۆ�3z���ክL����p���`���K�{Y^¸|�1N2�x}�Q�J������i�9ae�u�f'g5��mW�9q��+O+��"����EメӄO��+B�T�:hF�q~JG�ݮ�H��s��X���4p���{dj�B���lTF�I���R�Pܸw����֮���ƕ�a�]�C��pV�2Ex\3��\f��w�M�H�9�}3{� ;�\(�d���Ns�١���֑n�K��wU�M��Y�A���I8�Q��8�u<���\?U��[�a�CnX�������^�����ȇ�9�b%bç�k��T�]�:�cD��6Fх���(�~?��.W��-�8�}�tv�T9��}ikΪ�mut�Ի�d��ѬE�UY5�ՏM��������SJ��j��{�Z/��a�S�mc��x\� �+�h���.�b�gNwc�/h�����r��ZP���fǹJX!YW�Wcp��ٿ>�����ۼ�Y�=�cW��=X�3�BD��\�
��t��ۇ���7zq�,0N��L���0Wq�Ar�|��n֙�oQs��+��Z6����,�DX]�2��@xW�ģ]����|)�~�=����O�ȥm���'#�@����2)L�\eA�(�$OJ*�Zġ�%�+b���enr>���-'}�Ge(d`nmłۑv5��Ǵ8w���@s�����J�wez�>̭�n�	��F+6�qF�0�IQN5�^V��7<��P��b3fT&��{�e��q
ޙ.�B>�Zt�������l��:������f��KEBZޤ���W��Bk�gC���բp���	g��u{)��`dP��f��<T>���J"ou�RJ�J-n�iX�d@D2���E	�8��Et3~���Sg�pPbWK
���O����6��e�֍�Ƙ���"
�q. ��,�[��sm��D�wk���>J��g�s\m��R�3�����ib�ouy<�8��H
��"H��Q�c�)��ut�uTw-k�	�M�����mtKp-�F��Me��3���G��GW�x�=2DB���9@�5bY��-d���˖�t�������kݮ�Ŏ/3z=z	�x�A|���sѢ��W��;�Aӭ���oM�é���Y} ��x�����ZcP�9pr�����I
`���2�}��bR�*�����>�2����݉>����̅���6uyD�fےwS���'\\u��B�K���O���t
�К�)䁦�eI��N;R�@rw�73=�pk`�j�$!�Gh�q@ﺾ��(��:�t��)�ǃ��?/��o��'[����+84�1G>�%����l�ð�({]\K���5,�e驾L<X�|*i�f�!^���AF��p�Tv����e��/ܨ��^���/��a՝=ר�ё���I���U���Q���`�D���W��W���=3����������%��Y�pr���/�R�N�86�H�⣪����˿-�0.ڭ>�m_L*���)
�ĳg��/7�a���V'���-��]C����|`�'�'tQM*F�u�)�����#�c��"����ˁ�+�}����3�:����*3��xW^��=�kg;W��<_W���v���Uq����Y��W�X)<���gۊu�%�j��)�]�iS"��t�-��e!Ì|�,�S���<�;�e�pr���mř���B�]�nt�r4ܬ���u��u�.����`���:�F3rN{-<1ξ����Wt��y}W6m�/;y=�aq��Ap�J�ƒ�=WEY;.�m�nWD�e��*�B5�p����z��ڎ���˘�g�=(�>��D��Yx1'����T�օ[ݚ�⟃J��:DW�OtS�y<C��F��S��J�A�n��Q�m��)W&;�(������$ab`7
�
.D�#{���P��<^��Ocn`䂜�4��2�z�*�J��Q>8̧G(١>�b|�F�pЌ�qawSq�Q�^��3ѥN�Ȟ���u��ɦ;������DƟFNV(���*$�iר4�ltM�Г��IQ+B{z�ԉ=p����p�ķC�ex�6����Mg�n��Y�����%^Xs��ɯ�WL@it�46�sZ� ��d1����D��Q��js^�ӧ	�Gf���m.&��)����~y^�4��B�`�ϋ��j��pL�c=��غ�(;J!c��\�G�\�)ӆtM�70Y���`�'�"�0���\�5A�j���Fz�vs{�;���|~�fy?ei��Yû��z�*���0l6��o	�:<W|8��r�<.����{ı������ou7Z����8Ƈ�9����&n:�����R��Y��.#�oL�b_7��J�M���s�uC�!�'n�I�Ϩ>��Ͳ�t���g_�V�|{
w
�ʧ-s�雷^c����wN���S��,
�E
���
�ĭ��v��ϟs��U92�T^t!Gڮ�ӣ��f��V�h���rX:��iw��U�6���J6��Gm��En[���a��i���[n�Z�������u|�b�%@�%�<��%�0�j�٬�Ԏ�ڮ"�Q�29V8�t"�z[��c�Ҧ/ʺ��fQ���&	zvCx�V�O��{S׾�સOW���B<b�>R),v�P�t;\���w��,R	@�@�@�M4���]�%ZS	j[4�@�oa�O���6�!t#�2�����5����;c�Bn"^�~H�u�+���S�����q�H�Q������Yz]E�j�+�SuE�L���	+��,�Ɛ��肫���睈�:��lb���Q�����;��16L�?r9F��M�f�j�t�+��g�U���k��\3�dx�dY�6m���u��u/<��r����q,��
;B�f��
�wfH��}�vY�9���&&'<�_L�n��CS�;���	���3~�[ͫ}U����8�,̻��]��m?]l�|l�:��=ٖX��4�]��w0��ܓҎ�̫��N�ӏ8J�����*]J���ʋ�ɸ��6(�E
�\h��s:��}4��:�j��tq����k��~�E��N�pȺ
T/��Ku��#s�;�3�Kst�\Y����_�X�j���F�D�s�;4:Ӛ�-���p{��%��2+���
̹��f��D,���b�p��6�R1֙5�,���HZ�N�ـ�*� �EGUbT�sd�\{��Ng�T�^?�X�LՎ�UrX��Y�R\R��uf�T��C�L�ѫ]��f�]�ɷ��^n؀��L���FP�
�8Y�~���@d:�`�`�Z���*"щ�ŀ���Ck/z+��{��O%�`6+�gh���*�b������1�4��z���C1���}|���Nx��F����B�T��xQ�f�M�$�{_�[���C-�S��R���P����܊�JƝ�Wzg��g+\W�n�D@��ٜ�9=\Ӣ��	�(�����)T�p۟.Y}s�����G�j�,}�w�o���O���IE�t�u됏�9G|�SP���+���a����x�~b�!����5��&���y��Ɲ-�4W�u�=v������׼��y�=�G�]�@��[����N���沥f���i����W}�Y��������869JĆ��ԩu�3U7Ћ��:�,~ǅ�.=.��<����oi�v������q�iF�8�!���>u�(�Pz�𔲕�>��/9S��s:{!!!<G{�������n����e�w^�)�q~q�z�U���������i��[�]V"���ܮ*�Un��H`�莏s*R�����[,��=a��:�2A\*AVD�'��uK�{۰�P�Q�wg�6#���a�ܣut�[�s8�I�L'}�d@ڼ����|�*X�Q%�#P!�2���GN�n��(�,�rN�e���\�Kp봒����*�b�h�A�l7��'��\ɫ�UXӭ���/��\GPu�mE�Z�ng��sp��0!���]L��.�G�����E��t�fK��X�n��ʮR�{�K��`7aE3gϺ��jFDK[Xfa�;^���G��j�{`��UU�o��c3�6,l
4/�p�Ȏ�r��{s�׹P���a�V(�k｡>��;Fj�/Փn�9:]��7Au0[�"\;��/6�z�$�ͨ3��Y.�U�; �'�W�¬Vb���<t$oE���ǔṻ;�R7F��*.?\藕$�h�,����o˃4�۵�GA륷�6;�et���/��&%��n�`�M�[��
ݧ�5������ƒ�wbv��o+�S�GFұ�6��Tﶶ����vw:�i3�Zv�,�}a<#�-�٢�F���ͥ���S�5rV��d�J����۽�k��z�[�0�Ǳ�	&�^m	'l��5�z�V<���F焁Q}����H퓲�SiM�;�G�J����s�lq�h���A�S�LA�Ӕ��D���r�����8>g)��[5�9��,i�k�sd���bQv���MԕBrQ�[�Y���[�q���dt'�V2�6��twT�B����pu.§g@L�7e�(&��* �f������
w+��C��<�v�B��u5u\��MA�g)]�P�z�e�GF�,[P[�"-J��B���C�'o���yl�k	U�{Yy�����t�v%E��n.�A���ף�n�΀[m��� �\'m�:�JL��f��R�K�U;�.u!=[�宄m;��#�6�9[�4���!M2�as�ӱ��X����q߅�oA�0����j<֤*�O�vJ�u���e�.C+5�{��
��}��=��W��/�WQg-�c�[��:5��m�b�I�ϱp�4
�h���!��y�>�����PP��FQvnV��3#�F�2�%�;fak�Q��U��K���=�LnV�=���.q��b����D6򝫟B��D���+]v>}ӗ#��c��P:z�^*����䶞uc��!�H{���ί�E�G=-\������V���P��q�=t*T�k�:�z,�����c@�{S��P���ۋ�[��;�(�RI[hq�n�J������3/�����t&��lER H�Vݭs&�o�q���ۼ6��ؠ�a�1��:W��#�vᚚ7$Q�����6��\��WZ(��:�Y��E�fIwL�*0p�KS b����Z�qU��&�:�1��8񫳵̫U[��8��g�� �|�04n�C��; 5
{)��}�)���\�(���،U/:�
�qUܒТ�W]�� �l��Q�M&��&k8C�y�������ɜK"�@?����H�3���>8[[�C�iegiE�ƩV%[,%6���\4����p�	1,;F�T)Ю��XŴm,��C&jx�D�`r�O&�7l� u:�:a�B���U���,%�6�q��t�_�V��;z�	k2Ѡ#����L�RKCʰL�sV|h^���W}yYq9�30g`����V�Un2ɳv)�XU!+��Ea]������ �����QEF �1ADA�`�*�,TAEXT�����V(���(�b0UU��AA"	YQb�(�#"���AX��DX��PEQTV�m�"���X ",Db���EEb�
ĭEA�*,T�*(�(�
(�UUDDQ*Q`�TQ���
����,VZ�ETb�b1e�V-lEE��QDZ2��Ad��@c+%X�Q"�(�*(�1�VDU�*DX��+(�UX�	QA�,E*�� �,Db1b���m)m�Dd���*���TAb�"��J�1��*��#���0Pb��Z�E"��ED",b�2#0YF1���(���(�E���,D`��"��D�)U��h"(�X�X���1D*"(�E�*��k*,DUE`����@	�|I�2��T�5�O��
,�;E2b�G�OG�#ӏ��&���/�5��#��Ը��إ{�{?6ka�V����%�|��Y����a���1�D���N���uSq��Yv1S�a���r�.�������e�ݐ�Q��
3�`џo�R�u����{]
<Bp�6^�ZPHr���d�k������[�V�)�u���cb���hm���]s�qBҡ�MCe��qB���98uͫ�Y��W��:������F(�U\a@�2�x�6z�X)^Ю�u\8�֭Q}�������8�%ծ�R��μ�L�w���|��:�:�JG�8:�9�Cp�l�rj�5(�&�k$���^9�8,���x�~/��gc݉e�3~n�� E;����V�\�rIY�qk�T;�G�e���ȿ����E�ϸ�x�˃>���n�p�X��� ��D��lV�ggX��C(_F���,��P7�o~�s�\�΁�qg�*�����_��%ZTAT��1ccҕ��)��\�aN���0z}Zϭ��2:gd�0����qB���I���I���_���o
t���7�+����~4%��|�,Y���%bv��$�Í��_:�����>�;'�����9�;;/+;�����ġ���l5����/{C���^�D7�ǰj�#{oU̖r�v�|���#gMS�(�ߘ{ێrp�KZF9\c�)g�r=�A%��S����!��E�[����)�`���`���Yכ�}�?}t��/I���Y��h�i�ί_�b|P{��=<>�ݖ̈́�^̋�Ǳ�퍕�(C����M7��ȥ�)�gKȺ�j76t�d�2����fp)`�	�������F���T�q���5��4gY����w2(�~��kfa���v���.��ޘ3}/6�=j
Fydӷf�^�Ve��7Qny�
C�p>�
C�*/a��a烹�
�O�i.e{���X�g��{�/�~�l�
��-����:x��AL�Vϰ�Nc �����/��	�l�Э��Iy.Pv'!kn���m��k)�UǦ�nю��D�q��#�e�sk�����3�����*��2��`�t�m�"�xҎQ�B�q~�J6��,SC��V2/n���G��2���i�qz��&��&YF
�#R�h�(��y���.�]\����n&h�+�O�P'���1 �Ød)�u9f��W�em9�7,�etq�1wx����sq�t㑿���d�r�������nv��Y�.��;&s(�c�n�}�quͶ��8P���i�ó��Dmgu.e�v�j3EV��Tg�k`�<�I���ju�=Ѯ�.�^u�I7v5X���������U<�S��!o�n=ל��v�؏��תW���b�c��j��'T{���g�ǯ(8� J������h)�]4�˫�#:�������S)7�J��G�����*\�U����t�C��#���6f���~O�]�e	�Nh�9(��S~�.4��T3K2�������m%CW�6����H���a8�s�´�̑W���3U���[����R�5�&�ˡ���w}E��n=��4��Ní�b��iB�eL�և���)v�D������|�flu�LP�q���V�=�K�T$�Բ'�P:9k�=�����v�D��Q{	�W��S��U�

qB�aY�f��8�Ԅ���
F1�E몇����aM�\����ߗ]jjW���Y���up�B��\�0�øY)�ٱ��+.f�Z�\Vcc��۷,s3�{��O5�eb��%�i����Jͯ��b����w����0�tS��
qm�Y��wE�Uc��d+����B+����7��@���+K�P��oM��X��&�v�C+��ub�Z ޻�a�d�譽�g&��f�'kLC)�[D�2����6��s�m<�;;��Y�:����ݬZ�G.��X�X�����p!x�*9Zz�湷�$^�ͼ6ⵒ�j{+3���C���s�8Y��E)�� ��T2�p�mȻt�i����C"�Z2ҧ�wm�ݏ�\à�F5�TX� Z�c�e���N	V8���Pr�p5�=��g;ʲ��=�@{��m}��Ua՘2�W�W]�B>�):f�줡�?��_jx�0�zwX%ԟ��4Ws��R�λ�+Q㰜(�����P*xM�S�,��{k�Xʳ[�Մ�<��[��썤���-��65mi�n��D2�ޞ�lNҾ(->L��T\�!���ݔ��lf.ռWh��ŀ�kM5u�3���aƃge_;$q���T�Ӵ<9=�K<WF+Z��:j�k#.�4��*}�v[�	O7��i�W�˟_�t�QSh�r���L����/��P�#�8�=��f�ԧc����0�
nx�]'��<�$r��sP�v#w�ZJm�o�D٣���(0�_+��h���lCu���,���u4TM�gm)+E�j]�N�0�K��8�����x�n�pt���Z��gF����vL�r��ˮ���#��巭��d�o�7�o �s�;�vgaT����V���;��j�wP��]B2�f��#�5Y�-�L\�Ρ�sgT�5���Monw��f�^�0e�FL���gmY�L���tN��ڶ]	�p;z8�S�4X 8�I;������E��;:�:���}ZP;��O�8��[�����g����n��˵�Z��<��t��<S1|��I�Ԍ��V�cfh�����%��=S��o�g��ϯ�h6��C��I����U�ر�(թ�{˰ў爿e�!�T���c�]�g����Mi��[�b<Pp�+X:����i��O�6�z�$����s�E ��h�2�n������0nn#�P�P��Plc�EdQ=2�f����g�(㡤O{��y/;��Ξ(ȯ�,:+��D2�̥�=��uk���?�5u��l$�]p��5f�Rg�z�Y�U�R6X�K�ny]i�^nA�g��lᔚ���ܨ��s�\cU��>PoC�^KU�h������
㤮:����6��Z��:��]��.9C'�/g�X\�\
8�X�>x����;(���]S��\r꾴��,�/�UMԉ�n��tˋ�s�;�#a����WPP荤��3 ��0��x�5��{i<����6ɐ�݉K�v�P�o��Mӊ�RZ�)5�J�0IA*N������P��d����q�Ν�oSi<�FSe��c{����Q�y��6��H���7-�Pt����i�P[�>�|{]j�"q���@F�E���/�O-Y�� j#�!\P"Nϧ+���w���%��9^�g�ּR��Qn� �Tl%�q>T�u��gH>ž��bׇ\�o��b#�΍;���k�����ɂ�UϚV*J�7DW�(��>��QB��
��N���[�0��y`Fξ��P�'!�}g�R��^/���|�7�4lw�n����;
�Y��o�HD�֪M�K�`Ify3A�Nk\`��d1����$�x�9v%hB"�B�zYͫ��P�.k(�vK6]��9�\JsúP5��G�ueE׻(��n|�*yug�e��4����O����Pn�N-㗋w����<���7��W�wGH���ڹ�9��I��s
>�VMe
��@�O΍��JE=��eK�w��҉/E>���9�ˤY�q�0���fwn߶�d��D%ʠ�Y��Z�2��=��n�v��a�ȷ��u��ܭ�� �Wo)�N<b�(����Ȅ�'dp/�p����i�9e��n�}�:.����1]ot/G_lO��Wn^��A�܏:bi����Y���:��(��J���{]6Q�;��Y�1�X����t�]l�e�Rы��7FJ����:5���p��ؕ�vv�(��}��Yٽ�T�� =���y���w�q�t҆�7x}B�w��i���M�|���Й�^]�1�[�/�~���z�E����k�Etȣ�Q~�6�۔Q���l�郈X�E�Wd��wx�79e�m�i%�f����9��q%�<c32��NY8Ut6��Qפ��5f@�ѧDն�zr%��mP���+4/I��ڪy�uF��N��r�1��{�u���5�4�W%Uq�/�׺��ə6��}�2o�e�_�AH�������{qÖ�v)��{�K6h�wL��Բ�li-I�8�P6�Nb4����i�H�@W���ew�W;��y 5�ʖ��ř�M_O��C��G���������������Ti���R����}�����k���4���:f(�0˸mH��8�9���2E}��wi�q��AP���¨B�7[$�F���f��s��4:�sZE��8�*i�e���P�S��w�6m{8>�<k>,%�D��L�ۖGt w��;2[�)G�H�����Ҝ�:zR:��혞���f���O+����v��)��	Ι��ycfN7�.
�{%2���F�_޵��9�s@7+VVh�	�up��m7-����޳V:��6��Y�8p:ʱ�N4)ػ)���M���BI,�C���e[��=�ݕ5b�]�n/K���lo1��d�9�OF��9��U���l��Sjj�.�}���X(�����S��@�w]ܧeAq����f��־攜���r1+�&�{���(V�:�/�"���R	�<ͼ�^�ff�w��.ΆQ�T׭]�m����Kl<�홾Pb��tn�b�7Ɵӑ��� �oq�󝾝ֹ�X����Ȕ|�{΅8�-��-�݇�.  �j������[���)�㰝���7�13E�S2��]D�F�8d7�ۑvu�;�V���QrR��t1�_(ݺ^�o�l���xpO��2�*�9>-G`�SЕc�n}R"ֲ�n�٩�a.��dfx/��i��P�ԇ�U���*�k��Ț��{�U����7ֳ���❄m��qz���8�*dg�J�m����D���T7�'+/(j�܍*��Qh�(��6�`n���@����s��)�4�s�WZv݋`�P�mb���Zܡw�Xf�t���Ǽ�R7��GX�Y���{��.��ę���!�,�g�Kʔ�[��Z�}�C|'b�δ�^͍�\�kLJ�Y��],�"�8��m�Ԙ���0�$���"��zMy�H��]G���_}�UX�]%��c>%�6.-�NϤn�qiO�Ϻk�s�gݾׂx��;S�Y^�y"����+H�P5�HU館�;>�����"���ny�5��Ӂ#n�)V��Z�X��\T`2E�A��a_����G�e��������[t�h��F�:�­���ʧ�Z��Է���Ma��beGJ�bo�}�k�3r�MN�;w0t���z�t��%qz��&�I���'��\����sD��>�#%8�Qd,p��&ɵ5�r_n�M,oO�mK*�u�x�I�n�C�ju�P>�I���VP�����6z���^��6\�e4fŷq�{ͨ�Yb,:�;Qa��&(5 ���c��X̚���{��8��bpFgTa�ٲ���yV��
ز%��^����u���#g1ܲ�+CS�}y!��d.�_�P�b��x�>�>��ຝ����;bl���23B�V�@�6����9��:V�&�}�2�_��!^�]k��S��Z��iH����U���/z�n�T5'i�1��4�Q�onK(�ش�-�j�^WmK���2'J�݂Ԑ�k\��j��Y��xG�*�]�"�!��KZ1U�衝��|�*Ω���S�@b������ \m��� ��t�S�6J3�x "O.ު��f����Q�m�8`��3��?��@[����v�����+��rb��ɷ������j�AU>���窸�M�Q�裪%*�`����,[8�x��K6�j����ށǝ��>��凔s��{���Jm�?}�/g<~���`ZO�lnk�9`L���G�zH���鿧�
,�2�۞!�}H�S�>=YY[�Bp�6�k�Xp�{jQ�L�o��u���|D��9\n�Zr,����r��9"�%�dC�,�u']ܑ_�6��U��8�p lZ��VG�\�0p�r�:�c� J�kv�ǒ�x���^�'b��n�*ˑ
4Fϧ$�(�N��N��%����%\m�N�f�R��8d�0�|<ݳ�2�r�}^�@8�]a�3��5���%jB�n�cٚ����֯p� ZʓW�������f��'5�0DI�����S���VHÛb�/�S�v��P��2�S�M�͝8p�N}��F�ҁ���>麌L¼~����s�� 2���ַ�>������1]t�mm��x�*��x�+x,�ס�	���v�%c����i���Drp��_g�]˫�ry���-a��
�*��RՓAì,�x`${:�tZ��N0j�Njqͤf�`��L�	��/2�(�ƙܫ
�f0�6��xz�]N��-������a�f�A��+j�b=�E����'|�X�뻃�[qc����=ݫe����!}�Z��eN�T<���7�Gv�7���dvbUo�zn[�b�9�mjI��
y!�W�)ڵ�tZ�R����r�.lWyot���P������U��;�4Kxf����ݭ�+����@�)Wn�z	5I�h�N�X�o�60�)�wB�oJ��slR�oo%��l�ve����wh&���Ϯ��P�ێp��Od�2�V�OuI�"y֡�K!��v�呥Vto�!X��u4 ��֡Q�Y�>y}�Z�t��/�37y<����ُ����C���hp�1�p�k��ݦ�,�[5��4��um�����ۡl�uZ��P���:t��G7Z ����gL�wN���&,���� �+i�F����>Aj���hg�/�*��E�(��/"��*��W��ժ��&���Q�[����޾�y��H�r�p�ؘ�,�A���&�0�P�ެ�[z(Ny5=��3�Ն0S�W_s�r3�v�1d��B��.	Q��i�s9����z�oq���=�45#�4��gK�$�X��;�1.A�� Gx쩀��ŉ�63}x~r��];\�ٮV&[�u��M��3\@r�\�&L�Ƈ��,���d�!wqJz�����YJ�|bٲct��5��R��xh]��*�w�\oQ�s ��5�ڙ�l�p%�fí9�]ֱ�J�Og�g[�Y
���&�:jTi�|���#Tb�XW�5i=����]�z,��.W;W�׍��uoX��z�	�S��ś�b�8툶35L�*ܺ���m�c�mV����U��f�$��ƙ�ڃ��d�y�k��g:������2��ގ���|�xO�g�t����dT���"[���շ���Y��8���*�$�Y��վn���2�L�d����N#7��@���Qmu���x��N�r�Ba㑭t�Y�5F��]�X�Z1$g	�.�
��L'5i���%�g��;Rr��/evN��r:&f���<.�i9�j u�<�Y�5{5�ݛo���w��K�7�X�,�Xa̽� ��e��t��$���J���Ա���a�ڄ[V��甖p�(p�
삱!.7�9���w�kd�׭i�z:��E�8�|y3/*�{e�sV(�o��N[�3n�����@§=�o�h�(�o^��n�]m��[�DVv� �l�.��W*�N�L�ol�y���8�9�ԌZ:44�ޜ={Wi�Y�_fqK��5-�ֹz32@ ���hl����*�;�8~ލ{�~}�ъ"�0DV"�[Eb���Tc+[R��--���QX���A���� ��QEDDE�����Ub�F(�*���� ��Rګ"1��cUUR�QA�EDU�"[T��DQ�`�[,R�BҨ�������QJ5E�Q�QjV**��"��0U������U`�R�X(Ķ�*��J�*UDKj֊����E�X�TE��FҫU�c"�eE��QKJ�(���kRZT��(�����(� ��b���QF��F*�Tm*��QX���"����b�b��"�,U�e�V(�QAX�PQb�V6ʌQZ����QTF0c�**�AQPTb��b�֨�k*����DX�Q#�[V�"������1EQEb�j1F**""�����b��m+�Q-��
��QEAAT1QX�X��V,��k%U�m*�DbDUc�ȕ�
!Z���E�Q�
*�EQQUI~���k/���W��z:�72�$wy��(�Sa�ok��;[V�|��#�S�v�\2����*18�˳����T�����ﾤ�����Qq�\�Z�=�ǐ8n�l�����p�7�ȭ�2��[�n�Eg,2�$���FQ�sʉ��D`�Ӵ>?:6�t����+����W�6�SUc���3���rk�����i^�)���8�����V+��ŋ��Hz����ÈG�,��Aw}sh�7�6!��>}>�?����s�&��%���ɴu�g��}����*zw����a��}�6�I�H���2W/��kD4�^&�i�R��VN�Hc�}����o���y�y���}��q ��,��E ���{��x�3�1�їVq������R
~9�u��gy�m���=}��6��1ϩ�Y0�c�yg�f}�>Gރ�",M��.�_�7��3�G~���AH)8Ũ|���a��l���$c=O�L8ʋ����X|�|�́�ĝf!�{�q�`q��}��s�o�& /�n$��g����~p�\��)�����+�H���!߷��0�<O->t����O� QVN%g��&!^��}���
���k�'S���3�=dj,��5'w��m ��;���<�7���<���f�ua��`q�{�I�m�M0�9��JÉ��ɧ�CM\1I_P��'���J�d�8�@Qg�3t��&Т|�O��� ���|,���E�c���Y�ه����f�\�!g�}�,���OF$��<��B��H/�y�sD��M3Hby�:� ��)���gTR
l���x�!�i%t���g��6��T���?<d����S�K�86:�M͠���M���}2�T:��퓾s|¡�9��D4βV?��}�)&�CV-C�w0��a��wY��Ă�T>La�*)=�@����͟}����}n�,���o*m[�O�� �b��}0;
d�B)��[�f�j��s���Εc5û��`WBu� B"��8k7���&�h�ᣐ�_V�<���Kh���s�Ԭ�+]I��rVY��NڭK%�I���x����0���-�������X��5�~�<G�ϥ?�W�+桬��i��<�٤R|�g��sF�*N�];7�h|°�~���VM�ΰ�(�*�%��h��T+��&���:>7���k��s�S������H��2�w(u
��l`z�5�9�H/�Zb������>���gS�O{�&�@�+������������0�w�j�f2Q��޷�����/w�y￾�]��(��Xs)&'MSI�'�?0+��,1>d�n���&2�W�{�<E �65��"�_���nÉ�igy�]�|�����x��A>��}[�e�����k�y�uI����������18�׹06�O��J��& )�a��}`VkVx���%~��4°�u:����%y��0��o�M#���#�
�E}�e+�����j`3,
��{�������}��'��
���@�+�]˙4�]��^0�J��a�+9�&0�*)=B�hy�I�'Pߺ�=@��G���XU3p�gk����>���VOf��P���a�wF�
J�y��'����톽�i6�';�3�L�!VڐX�=2�P�A򇆵�U��M��J����c��	����Uw��z� �H�N���?�z�0�/�x�%x����0��Y�K��sS�J������������A���N;d�;�h��4ɽ�>v��|�_����iR_{/��3�~+WW���f��p�zv���go�8����>0.�;�'��~q ���l�i�%E�|�&�u
γ�2�������d���5����i8�Ɉ�0Xx¸���}��,�$z(����߳>�%��|
������a�i�aS��\�u�P�N���
Í�*O����4é�:ʊrw��:����u�4�_y;��<E��V���j'�햪���4o*�{}����}�VLg~�!�RT+<M�}�Ci>B��x���@��Wz��:�+'\g���iEXk�q4�RVh���'��3L/�N�M!yI��'r��{X�_T����2�*+�.�@Qt��Z���L��7��q�L���]�ɸKF��Mu��jҼ�*G���+'�Va3ZZ�n}����j��}�Vp���1��0�W$Kzuc*r��l��FV�In�l`���W8���Wû3� {���J�	�i���ޒ<	�{�ğ{C��>�$ڲ��ü��H�����f�
��s!��|a��7dǌXq��솘k:�=��q���d��s����g;��Ti��eY�W��Y��i���m�O�9�s^$|�_'{�I�x�P�_q1M���0.X}���u�!�q ���ʂ�3�J�q�I�+8�;�ͤl>CK���i=���0�T�X�X߼8�z��(����~`o��>@���G�I����?}�c����d�'����g����%|Ad�? 8�^Y����}�{��>k_o�����>a�c0�R
�S�Yǈm �!翰�<E�aP<=�:d���v��w�4AI����ړi8�I��悸���>g����q+'���|}�#��|W%1�U�}����>�Ͽ}��gC��%�C�6��@���l1��d�u�Af�;�?���H,����I��ć9��V|C�d�;@�Vm<���CĂ�����i������*����U��Y��i_���K����_���c�Xc�����iiY��Z3��R�g��e ���P�������M0�N��Ǯ�>I���<LH)�߾�zé����Ig�Eǂ#�F�X�;k쟢����x����jz���2Vw�LCVq?��1 �'ɲ�I�8�k�O^2c=-�a�?8��PĘ�C��^�1���Y�w�!O��1F4�;t]���{yn����>��l�;>�&�
O���5���
��S��'�.�i�q��s!�m�&0�y����A@�l��PĂ�7��h/V��d���퇺��R~B���9�����.���/�#�@��}d1����?=�����Y6}�w~�L� �̇�T�������M&=I�_�i��\�|��s6�Y�Ne<���Aa��뤜�d���/�|�u�|��y��k�@��׈vwy֠u+7/������I��
������x�^�I]��t�01��߾ԛ�J�}���L`w�m
���ǯ�X�m�O�>��y��X��O[�!���r��ޥ�h[Ԣ�%L���̲m	Hn����s��.�M`�!��Zͭ�������l:��Dǘ�Æ�;ӟR)y��2�`ys���M���PK~�V�� �}z+GJ@��f��W"��q����x^>��x�+���� �h��K�*CSY��>LE7<�c����Ӭ���=�Y�+:§'�ֈ):�g{̞!�������O��@��i<	h��j�Dƞ=��	Ɍ_t��~���¡�t�k	���P�<-~��������u�i
���4�T���&$�u�1�N�__�op�Rq�q?K@Y�La�>ɤS���T���r"~[J%s�(�$�߯���b���{���Y���w06����n��%I��Vx���a�6�)7�tϙ*�ۊÈT����CoY:��~�����@�1�س����'�]�ί�����N�k�8�Ag��s|�r~j);��<jOuC~;a��
�1�6s0��P>J��z�H
,�2�I�a^����H/��ǈ|���3v߾;ӗ~xg�0g̕�E�d�,�~�M$�
�d�{�z��<aSɬ惌㤂�����6�d�Jɹ���AkS}�/�ݛ��z͡�?8�ɻg�,���[���د��ѯ_M�5\�p��<	d=�q$Gl�N��1'�>�㴂�<I��mE�XWgsP6��*�tM�偌>Oټ��c�L����J�aSV�@��s���7G�wq&�J�,P���`�Q�i�È-g�'C���Ͱ�c7�:�"�Xx�&0�����0��N�^���w$�m�����wRmE''�`i��*O�����u
��-��yx�拽�������C�1�!�����������m*C��z��g���aXo^�A�Ԃ�Xz'ud�QHjs�j�I���y9̓_XXu����j��=9F'���u�3�#��� ��s�a6�W��P�Az�<3�h1�8��~d�8�S�T��?2w(nZE&�����T��������u�AG��&?2]Ұ�����o�n�'�Z��Ջ#�#��|(��nP$x����p���:�9>�c>Aeg�3"�Rq7;�i���1 �0��'��C�Ă��f�hmE�P�U���=B��{�;��tc{F���N��f�Q��s�S�Z�V�M�t4�Pu!�q�S�Φu	����3ZGCn�woG:,��2�^^hdr�"�ǋ��LKvj�)\�Ӯ��yb����)�Ҡ9=�֓<�Mq �J�ן�qXŔ�2^�RB��������r�m�js����;��$����!�s���g�+>d��M��w�
AM�w�f�i
�;܆�T��7<�봂�a��3!��E �^�!SL=x�$I:�Ax�rs4�U���3H���0}�}^&��iE=B�L�'���I�
��'C��u�a�q=7�Ԟ�βV�b*�R�{�}���3N i<�:��6��b��SI�Os:�x��l�>J��>ɵ���?xfǽ�@Ĭ�C�����ƠUg���4��Rx{N��������i@�+�����T4�_Y��u�m�a����4�x�Fu'�����>�.Ο������]����@��zЩ�8Z:�!Xi6n�'�Nv�!�޵��%2_iR
Az��z�!R���݇���n>� i�Aef���*)'~�O�6�0^����L�\����;��������>@�)�0ǹ�ڐS���a4�����}`T�f�]!�
��������9���g���a��a�H)~։�eI�+���6è-H�����3�G.o�?'*W�g�'�|>�A������rOɴ�4�!�s	�Ԙ�Az�\�X���6[���L@QM�P�6�Pީ�I�+Ǭ=����+P��q��T�w}P��Y��j��{H$�z����J|4�hW�O9�h����1��w�ܟ'ϩ���<ՓME'��i�Z�ɤ�u���U�Z�0?5����q=a�6n��Ұ�1��S�w��o�<�ݟwĜB��yLI��?0�9�M3��g�>�ܛ@QgY7�{��)<B���w�������2OR~~t����g̕�K�/3bAx�4��Av�G3{~�.��s�{���#��m�ڏ��FQO�޽�#��uRW~ӌ4�ACP���:��Xx�2z˪N!��|����� ���s]d�E��w����
��߹�h|��t���|�8¡�>s�����}����:U����,����}�>�>�@����'�-I���q�ז|ϝ�c6~��u���J��cy`c��f!ӽָ°8�O5��m��d���s������o����甊�nMW}�Łн '�ػ��Mv~9x\��/cy�9I�"��^�}9��n�}  =N�Qu�h�9��9��r�]i�Y���PN,�8�hjm,<��LH;��;1J]�Fqf�G7���G�U��]=�ٙB��;�|�Y��#n�tpr�]�_��h\�V�HWam����}ݶ�BU�{�
fBn6�D��BKk�� A�z��8��z�<g�3!�aXx��:J���&�����J�C�&$���g�_��3A�5����I���wVN�zvɌ���g��|��Т��k��'�wD�2�`q��|�?&ٝ�b��JÉ��ɧ�C�����bi�N3�*,�kV@Qg�N�S�@����G�A�N�R�}qQս�}�^����ɿn�w���:�^�S�a� ���څM��_��w�M�a��4�'�s��|H,�a�˦q�E ��(~CL�8�!�Lv���c"Ϩ�,�#·��5�;����,���������(��}`V[�RW\�w��G�>aP��w�!�u��w���'֐Ro�`i%bԟ'm1���^��u�Af<�>M>}=��$kU�P��5�y
Mw/~�އ�%a��|� ���bt�xi�
��P�?3�Y1�g9�E'�Vx��4a>B��ӽ���0�<�~�~|J���u����PU��2<$�A
 ��ʸ�_V>���R����a�D3�O��HJ��̲~j/��0=j����E*��1����4�Ԭ�~a����4��Xn_��������ڠ �����e	����>���Q�c痟x��¢���
,����H)15�i<d�ǌ
�7Aa��Nv�O�Led������ �5繧�:��A~�6jÉ�i;�5
� ���7����*��V|�SY���τ"����'�Vc?!��9�i�c&'��w;�m��Y<-�~zɈ
k���c
����͡�xî<C�l4°�u{x��B�L���a��H/�nV��	��TVJ�'��I��${�-Iӽ�n0+�x}�ki?&�����?'�6ʊKH�x���lĂ�'��n�^0�%M�a�+9�&0�*)=B�hy�I�'P���oZ�~����g4��4³��m�J���m�~��d��ᤂ��^���7�B���3��d�m�O;�3�L�'�|.eH,Z�������Ұ���͛��;�`D2+���}�wԷ����1U��(�|7�콝;��Eb�51vcb�/�H�K9��ւ�W*�wН�=G�rX�=�{�O��9A�_	3ae��y�x �����j���I� Ĭ�8��5@Q@�T���x��1�����U�CL��mgY/��OY*�;�d��R~��A������<�9���T�&�t�v��|��Q��6�+�m\�}F��{Mb���)R
N�P��LE��Wv���{i��H,���3�*,�9�M$��g�zk�]���w�j~a�ְ�v���L@���hX��'�Emj
���GtG���Ka�q!�8��VM0��C��g���+?0��i�NZAq�Rq�P�}�1��Xq�>g�0?g٦m�Su�����a���i ��g���֞F��ّ����yVw޲�
����oR|�ϵd�x�!�RT+<M��jI�&��1����?0��Chq�VN��&��iUI�)��AIY�ۧ�q�?0+�f�Q�|Y@���:�Øڛ���ye�'��'2����"�X��j�״1 �=��iX~}Cw�8����?w2mEi��C�
���1�d�����04�u�=��q��$R�d��R�!��*'*�7�o�ϼ��Y��!����r��hc���Ny�׉�2W�w����);�E�d��Y4�`\��>O{��a�
x}��,�=aQa��I� ��3yb�ڣ������Y������`x�y�笘Þو��
���w�m'�q%{��
����5w��������,��e�q �����`~Co�
�s�����/&�MnICzo�+�Dx�a��2tݘͰ�c:§�� �q*x���Av���4��@����>2q���z�(��
ϧ;�Rm'�T�s;��>�c���0�P��q���v�������u����K�
K��>�m1����a�/�N�]'��d�P־��)�S�z�';C�g�Xi�O��I��e���xa 	 Fں��'F���{>������Wl<C:?a
�)+��هm�L��J��E��w)�5`�������La�:��T��Ăϒy-��&"�Ss�G���A .����e☌؋�a��-��:U^��o.ezzw1k�՝҉�r_h�J��n�����J��ΠT,.����c�8��$�{��No���M+����\[	�.��B�"ryv��2�Lz5�����X}�r��ޟ�Y���Yx�I����Wz���=��xGWJ|�w[����l�Q���C�x��|�C��>Aet�Qg��4���l�Ρ�)>M�i=gcMvn����&1`�ì+���oi1
��6�׬a��wٳ���q[������g�J�|���Ͱ���s�bAI�;��[I������꡴��x��y�ܟ״�����_a)$�l�M�_�o)�E�So��q&\���N��s5��Ǧ�sD��>�а�Z���]�'\騤�E�}yXQ�}�kˬ0h�	�n�A��Y/ܠ8|/��A巗�_o�>�;��7�3�\X����4�����ؽ��f�jC5��X��ؒv6:�(�ur����l���J�pMC�UqX2P=��Y���ǆY�_B�$���A(�%�3��6��{�h��`c��H?^2��0`�ꕮ��9�_�ZD�F�f�7(t(���:ys�*��0������Ϧ�{����
)����u����G�
�F��s�6�f.Dt�ۑ���@|�nY���b���rC>�9�YQ�j�BfYi����bAMϑ�v��_��j�Հ�y���\m7MGh�:�T�(��h�w�sk'Q�ͼ�R;x��
<�a�_-b�8�l�Z`��we�˺9|����`+��#�\s��A=�DovtͶ5��|�-�Q�}��;n�#�1�J�k�dm��r�����+zoG��V�s�D���˪�rxrwmoR��x{ޭ�����(���E�h+�hS���>��|���j�x
N��0����G'9,�����ӯ����iۨ�����I���N8��e8������ڼU*��/��z=��
e�A� ��B>�����v2Zr	+��[�����MZ�$.���S\��kS��t���S��/�g]�+̌�CU.�d#�Sn/�_Jq�r���z��
C�{�P�P���>8�F��ՓX^���β�M���V���,ϭ:���i�S�ݳ�2�r�s�Z�3����V��S|�VmB�9�٧���K���1��a$g���5�^���E��$��/�1�.]z1�VO������r{b�Y�$�O����r�3�{>����Nb���(
�C����J	��qS�������ϯT´�ıY�CS������|g�/_,>�P�C��lO�o)Vmw��]�%&p��,E�%�����E���^����?Y��Qxw��x'ZX��{2�A�I��u�̱5{4D�n�'g��&8��\U0�mG����7�ڙL�y�qp�Wxh
�Q'�!�n���ΡS���[�;|�s��.����\�1\.;�Z�].�a�sI��ݩP���s��Y�Xxn�GT�hʨ���{�x��+����j��������:��}�0��"��I��0�ٍ5텑�eD��/���\����� I�ê��%l%R���΅�xp�iZ8����#��4��L�y�j�z�L0�2�u�_w5������*���O�{�R��oU�k��"i�~�	��n��"���CxsG;��1�D2l��F�3�J�W��"�Q�
�p�#��Q�yp%��/{:��Uֻ�^�b3_t#_�XC=�UpUSSq~(�r��պd�TRucz����I�*j��U�t{����}+K|lLh9�3������(�Or��a,������[u\�t�7,�@�o���s1jRO�h�Q^����\^P��"3[�]���qb#�<�9�x˰���@mK+�t��$�%�G:5�SU���>�
���"(I��n+�R��)��)g,*Y�{\t'�f������x3��lF�+:E��3�vz��Rゲ˲�{βP5��Ҽ=���P&}�x:��s���*�t8�m/4̯j3a�{�R�НH��v���Y�̖��塀�Wi;�g�fk�١Fǔ�ű���@�)�Y��b�0��'7�����U�񬹱�n�i���i�[{ڸ��9uBeN
�{5�kM�A����������"��S�0V&ouFv3C,vYk(k��M>B��j^:D��-���g��Ba,}y��[⻨R�n�w��~����Dٷ�NwZ2�wk�t;y.�P�T��u�tY��s�r[ˍc��,l���W��ˢ���2�њ	����<�;r������N��]8���vc>��GD�
̇���w$˖�Q����Ke�U��=�tN��`ъ��Y�nv�1�3c�����bQʔ��Q{�b�<�v�-hN�/N���z�*�ou�t��{���E���L��6>G��ڣ|̰�)�����zW>.��H�>U�Mś֜Z�l�/6,;{Ǹ�q=;m���n��R]D�:���*���9��U�l1evMR�֜��7&��x�y��ҌM�g`��o]c;{M_=�&D�kvM�?=��m;�Z�襧��8��e�M�'��J�ܼ��
z��ֵ���9�[{@�{Nd#8k��al�����Ȩ��g�sn���z܆^��,M�h8GR��L�g	L�{��:wu8�9�΋���R2�|��SL��p�k���ėM=�A�Nюbr�c9,Y�!�"��B�^�N�,֎n����3C�gNtki"���O,u,x35"����wH����9�P�­��s2��&n���l�����d�A�t:�b��}� �-�{�9t��sMS���/�8:�`�a�ǰ��>��r����S���P�W��7���	󙷺Q�R��n@&ݔ��r�,&`�]f���bF���HT��*������v=���H����sPZ8fԛq�I+�j�kp�Uʐ�HIg����8M]�$�F\�$�(*�{W���U7JCEèE�q �b�����dl�ܱ]�J�E�:���m��$������PyH�%b��7���]Xt�eF��;P�U{ �l.�Q�����D�:7�yZ�G@)b�K^�xpf�;ʡWdU�
|���
��E%"3
�w������6�vi��o��]�|�Z���y���v�Aw]N�)��U<��5p�(���Zp"A�P):~��讷���e0���%SO�����3s��w����Wgn���e �>=֬XJ�c�'W>w!R�v�f<�ER*��s7I�4�%(Ze��r����?�����V�x��UX�[hS��g;��npY��<�SM�C@�F��P��i���W(����vaiV��K�&#BCDP��0�d�U������4�2�nI5%�|3�9��^�����7��@bW��.�D�cY�Sr:nQ�;�
���qˣx�8��Rѭ�5b�K��r*��S��&iu�綠��(�"*�E�

�ʖAX�,TX�µ�X�k*������UT`�*����F1V1�"b�*F�l*�����V"��ȱV*�(�0BТ,U�������"���*�FEDX�Ȫ�D`��QAb�"
5��
������0F1EQ�b�TX�TUQjQA�����b�DX*����AUUF�� (�������Db�FF*"��#TA�"�TEb"�EH��T��F�F)R�Pb�6�b,QDF"�*�0U1DPU`��b������1V ���H�����1PAETF6�F-j��`�DDQ�UEX�DE�QX����TTTE��H���""0E���Nh��ӓD:�N�dk�3J�<Dup5ox�����Ǒ��%�˲Mܓ,WDSby�Ç�8p9K�#rW��x .��O+��N5�(�./fN��ux�5S��mN�wFN�2%�G`1)�᝗���
�j1gE�D��������#\:qFz��
{���1V�=�eck�ʭ{Q�y�U�U��Qds�D�-9���ڀ�eI�dL���*z�
�X���X�W�V�)j�Smj^�)��4:�a�+�9 ��݌Otx��W�������uf4q�]֪�w�4u���ͫw�43��:X*h_]�m�����F��+f*�U�'��CR5x��o�TdR2�".fs�A�)���
�%�K����)�z�.�:q�hc<���=:ٰ��.����]@Q�ל�]8�(Ec'�1�#!�[�*��TUE�ˆCq."m���s|;�L�mVnH�;�4�U�:-����^�-Y8%>C�q��9h8}ǯ�D��I2���-u��!ه�?N>'Z���n�v5�3�5@ˍ����T����W��i��������hV�M�F����~�?|9�G����5��+�v��;�F��X�滀->�b!f^{�n�@[!���:�r�F�9+�7p��e�5�z(-�/�SZ��ʟpu&����l�����*�����{��^d3��(_Nc����>�7nVC�]���5���1�&9��˔�R�GY�0�x�*k
���R�g�{����y5:�+���	��騳yx���0���x�z����a�^
8�o�q���b���4���cԺ��2���-.g:��\ygWx<�1o�Ğ�c�ɛ�ÄU�?Na -;*�rX��;�o�WR!�֟����3�h�ft��Ϻ�XXTTh�9��uu绵;�d���T!�c�k�#���p��B�i��P���v��;�����{�K:k_s^�h#Bs �p�Q'*(��uP�`^$|4r�;|m����[�a��#Q~�=r氳�pT��SQ
�q>:�1�Iڮ	�_�E��-Y���0-eI�c�g�DPy:����>����P(^��t��E����o�~��N۞��N�%���`����(��ͺN"��0d�A�����jFA�@WQ�r�� �x�PI��=��,`Y�E(�5i�dh�jԆj�B���a7�tMB�檴����W�a�c��PX1�>Ӓ�K8�X_�eY��a���`����6�j�&��_L��|߆w�#�ƌKl��vJ�{�o"];��v�I9��3S���W�0�*4���]��n�h���|+2%E6>pY�ZzD��V�`$�;P�N�>���s���)[�ؔ�9�x'9k�B�r�� ��W�}U�|2y�ts�'t|;��y+[^@��f���������^Z+�h����K���M�$���-u֨��˱����^�{��3~5��uܦ����]�f[U;���2��쵩!�a��A��#Q����ay�ܛ(��6��D
΃���	t=��ʷj�Z|�^����⊉(y>`ȻJ�XR�T+�j�z��ԩjWF�uD��[Ec
�V�����]���@~ٞ5�6z��e
qX��o��%�2�5H��<�ڇF:\�J�g�o�Wq-��#����_�?^@8^�:�JG�5�iq�Q1����L�|*gM�u�!��d����>�"�L�{��|��x�ת|H�%���4~�i�׫;3 Z�ߜ=P�-��,��0��t���"�rh��Ts��p#<rqE��{���mumqKR��ұ�N��QҔ��QƋ�)��/�: ��(����B����l�����mH�܇��:��p�s�J��0��n��*'!��ĭn��c�{�j�=}<d6�k�L�|c�_^�I��䎎�q[�t������H#\���Y�����;L��\<R���pg��#զ_H8�������;��r���� ��%�U�4k7�N�ۻ�B{dW�b'�t���A5���a�}��'X��w�v`Zi�^
{Ü�B��3�Y��vJF��K�3��M���/w�����{�ּ�6�["~��"	�N,�6�T��9y��(���E�y,�rI��[5b�i2��<�8E���������:k}�0Av@򪇏٣=���z��|'�G~W�~���p���v� ����?YG���x�����l�,���0��7p{��f��׮@�*����{]܍C�UK��J;"�a�.u�*���#�s�+��`��F�R�M��^F�m��}�0��"�M�O3#H�^k�V=��7���Ŷ�tYc��UԖ�]N�z��t���^t-�ÇJկv��ϥ��x�����	=糤UQ�n}� Ot�WP`�=�_���>�8w��u�Ҭ8c �ʝ����6�(�L���z�=b���n�,�Qf��%"$k�E3��3Ц�L�Z�@���TYF��o���(�Om>��M`8gڻ���F5zU5U�iC�QF'�)���"�vq�[�*�Y�C<k�X��a`r�6�s
`��e���zckºU5���E|ǝA8�nD�m�^�	G��}�.�L��3 ]99oJ�8M����`GBk���#���U��c�9�Wn��i����b�y����8���wIY�{����������_bڇ��<	k�Ѝ,�uӍ�,�+�qƌ���S0A�T���|w�b�D�=���'�����udO�BQ��ԍ���]��=Qa�Lڅ��,��U�f�͊;%�M��q�yh,�Ǧm!��`LOF:�N6a5���b�ǱH�������E�|�B[����v�����
=�エdVEzS���Q���,��ȳ+n��>������"��]��n�p�}�]�����o��j������a}j����ۏ�"��Ulq䷯��e+Ζ���Ni�n�D�v��#\R�G��v;�JƮ���=�c�>͎����X���a���A�4�{�"h$�ju�X��=g&��CLsw��� �a�[+�M�)��5@O,w&�:�Қ�nr#�R��3]z�jN~{|{�t�鐮(�̪��dQ��S^��,�np��Kn���[1GE��#1���0�=˻�u�UkX6}eQѿT���ក��# ],�ȗ�*����m]�}v0��qt1H`Ś�{�ee��ޞ��6��'Md�e3������A���u}C-�v�;�����Wk��u�Ȩ<�{�/q�)l]h����nS�
�ge��o�Y:�ꎞ	1�r�:�ݮ_N����4+K�N�ӗ6�oR=V��;#���U_UVfp�����K�â��(���y'��Xȓծ��y`�U���h��]J�
�}9yw�R1s���E�T0�{�F�+ڨ���gls3�Q|���f�m�a�s��<V�3w�s����8���u��P7+1a���~/�����P� bdX�ߞrw�.Q};ӥ�촢�����΂<�}\F㑅S<cNU�%�c/{�/o�	M��R>��>�*x����C<�H��g��+Ocu��kb��}]�<�R��0�"�I���W���:���My��#=����0�DdK�x�vz=�{��#�r���O�CҚc=�p�.�������X��1~�h,�(�&�dO#O�{~���L2 �*`�<�B�x:tv�LPy�K�+U@a֦�ۯX|���������EY�MRP1ܣub����6Bq �p#��qD�Q�:�\�;��kb�q�l�zP2Y���v��,�s��ňSQ	���eL�,��NY�c�{u�"�2��s�e4�J�D�J.?�Z�S˿�j
��Po{�6�Q�20�ԋ�#�&{�iq�M�$H�C.M��ou���s�&i�P�Y�V#���R���]K�3��N	Y8��R�s8*&��C
|X�Ta��eܿx�W��K���Q4,�P�W a�s&����L�<�A��s����yP�Ĝ��8{�&�->er�c+8x{>�z�!��af�(���q~U�0S1s�.�O�Σ
un�_�Ż�r���n�$���ur�,2���w��b�,�R0�f`��mP�ؾ[	BKD?d�ي�nP�%-�:tѻ3�0ح�,�UdK9h�Σ`fc�X����߈*�`�p��k�����j�^M!�h�{^O��8"��+��\��FVSa\8��M+��i��R�>�˱���:W������E��SB����;���G�c����n�D1[A��]y�D��M��7<,_��-U�\�Xu^��p���`B��l�{i���o-�q��WQ�b��<���G{3V;��G�QU�V�T����;�b�V�ﳪ��@VW}��#�s<h��D��b����p�R,lK�zٺ��US\cy�ޯ_d��÷}1&��*�`��t	-B�sG�cv.��H����Χ��g/L��n���ۺ������=���]�{�&� 8����76�������vۡ�9[5�;�iŊްv�Jn�8$��I����²���_c��Z��::#�M����� �l(�3޵�3����j�D�h�P?��x	�Q���s�تؽ�(����]OG�T��e�A�QcHF���E�
�"�g:�S�����`[ƛ�jE����ΗV�"�c*w��U��@�9��(vA��\t�wv�����W��j4�k�l$�8���
M
��U\:�D�T&b��Z޾�Jڕh��`��T��	�''>�*�,lK/q�gI��tC�����"KRv�[]�[��1�g~<	�6t��7	�� Zʓ^�+`_@��Zvhh��̷���u�*Y��>����ɚG����?<|����/��j���jY�j�9��B��ژ�-Zt�n��O����}��^ !���_k��h�ڇ8ܪ��Q�2��^�����7'w:���j�Lߒ�
n�F��>{՗W��=WN۱�>�8�5�L]_��`	�vo^�2z�&�M��q�}��aD����#���[��i
u�P������Dҕu�؋q�gzyw�Աz�iS�����+��WL�����ۼ8S]\{ܵ��w���|4�;^ΡE;��:��$|�܋c�Rv��빧�5��C����Q,O\�{�^�h�
��2�U��E�}�E���i�:��^�!_ml��^"9hrnl[LsTu�)&,�P�CGm��1�Ç���D~�Qe��h�ӡ���sL}g7�}�}�]�?{{ϰ�Б�o�_[����o] hc�>0��P�V|Ǜu�aNp�0ӝ=�#VZ��/y��ۤTߟZ1ѹx�:Fd��<P3v���,����[c�jNZ�����z��b�x��'���ב����dn]x��ϫP�ͪ�o�K�E��o4��#z������^���R�j�H�U!������]�*	yU��y���5@_J�-�#�/Lm2���w��s-��͞5p�n�f��,�+�q�cF���\96: x|B�+��⡬*h�}m�����[2��.����=�9G(��]����o��xt�U|Ss\�Zt-���_v����.���G�V)�+��O�:j6S���A�Y�yZJ�eD�7R��m��Z�{0�[�O�3R�
�rQ�u�٩*4�3� Jt0*7TK/#ZJ��Ӕ���k&5q;)�	�`���^;(�T�B7BS����-v5.�(b>^�k��X��η�|���؛y1�o���Ã�1���1�Bcmp5������P��5�-=�㹏J�ٕ�-s;qZ��b��$�wS�k{��P����WBn�g�{Ӟ,�����yP��-��0SV��Ø��j�uܾ����C�:��={��a����n��D�
mF� d�����9Ɨg"5_,�}�{�]螝k�͙%|6xᡷ,���'PvӚځ`7{rE�2NzN�5��aRC׭{�⍵���z�HF��a[bOS��T���0t�H�׷���Xy��vY�=C���3;5����&F�S�VBŎ�o�*[trb��6������m����h��v
�*����YDTf��Q���z��dW�K�,�p:x#9]�f�ˣ�Z]|�����k��LQ���y��np�D�FzrP4-ΔIJ��9����,��׼3��mH�N��7\zb�H&����1yo�EQp�ԛ�O{rvk7�������L���M��ۯ[�V��
�lCt�yU��T
�t�>�&����}�o��E�S{TU�}�덈ۮ�Z��a���E}���n#
���)�����&7MjK��[�bp�W���l�Q�$3�9E�3ƞ��g��牜g��s8�W^����V���#z#I���W����AY�ƛ���qucOet�Z�-m���i�
:>��IT�[�͜�H1XFo��x��P��cL���5��Oak��[��ޕ����K7m'<��i��k\[�9�"�^��8(_hۓ��m�l!.=Օ5-��]�]��̝@u���rvZ��< ��	9�����"+�D���q)�� =ӸhX���ɥ��=��e�2��-���5]L_mm��Gt�1,��k����)� �����j�,<�1S�讟\���v]%%kj"�='H9�_f��
�j�7��[y[��lz�!u�N5�����i�m��˙�+�(��)pԶ���V�IZ���{�{X7]֏�A�5�ɮ��FHwjޠ��^���*��N�g^���t.��%8μ�Z Cʳ.SJ	�RWn�UҦ:�yun\*�N�rWd��z�R�V]��s���w�Q�n��!��8ST��d���3O6�E{�u�v�J�]-�{S���X��7H%|��cĨ��E�8]�ń�o��{rs�m:���þ��A}�9�[�l�S@!�92?u�B���(ݜ��Zn�jwt&���d�qh�F���qg�]���Y*[j9ϲ؟tt�ge>�M�E&C��-/�*En�LN�pc����[�<+����U��K+]��:�u ;GKo�>w/	B�K��L�5��9%dV��K�n������&s5�����]���UҲ�֒��y��g�]�J>���"�2.��n���)����������
��,1܎��6�8]⋞'L`/:�.�nK!KO�����wK�x��:���k��+��1GTa836��Cd{��7J�c�Z+Nl�'%z�%wj!b�/�y��J���:&W>q�I���Eɝ_en�m�$���5>(��S��Yw������<|e+� [IZ�M�
q65��1��;B��ņ���J��j"�[Gv�nЌ0�W
K'���kS6z����<良�k%�\�ܼ�[Ň!yV�09�S�:f���D�ܻB^۬��$�An�N2���ݧ��ۡt��6��)Q���:5�ѳv3���H���5��"�w�����;�l���Q[+�f����_e��Ub�.�q�������:]���OY3�&�G�\��z�l���v^�C��[U�V4(*���(��n��	؎�v*��.�G�/J[��gP��]<���_v�l��ϝg�٧3k+.��d	ӧx�#�h,�o�U!KA��֝/��	R�!�Ͱ��jٺ��i@�-�sP��ÛB�y��{��x� �R�{K�)MU�*EvV'g^iS�w5 �O��'�EE�UA�EDY�DEF�R*�cV(,��QKJ���ŌT���TQV")���kPX�"�`Ȭ` �,Q*(�TQb��5,QV
����AU��b�A��U��1U�b��
Ԣ��Eb� ���X�b�Y*U�2ڠ���AUH�cKb��2ڨ��1*+V
���A��DT��$EX���([bV����QDUDUF�b�)mb��DQJ�b*�,UUZ��"��(���AU"�V1UTPQYl��TTTEX�(��kETX���
�R [A�����QX�Q����DQD��U�X�j �Ԫ�l�"1X�,���X�����(*ȉmX�~�s{���~י����v���ݠ�ֻ�L�kwH���b��loMu��(w/x�{�-g�5h!��*+���]����򪾯�śP��0�nRU�٤a˅�ث B7���T�n����(g���ҽIX��>��VS����y �A��/}�~���bad���
��"}��k���f��zC�A�Ɋ�]ٚ�64��[���Q��SYn9��2GC���W��_�ux-���4V�ַ�R}D��Jq�c��HĖi��輝��k�L��+�n�A�>ޔ�YKT�+ K�m0d�羟i�YRk���vDPy:���s��]�q��N���>]x���4+��z/�n��B̛,�+c�6�8�S�0S1����r���;6���U{"K�1�P>�	1��U	��|�-'Q�� Yݵע숎�ׯ��):4��c���SܯD���dN�/b�ҳ���A�*͎򌰺�������Y�[1��|y�L���眯���f��8��&�mA��8�mynv^D��lS̻�q|��t��ٴ�\������Kp.��^�Xn��a��D�҉����#xs��c�7�;��K��%y5;�;���I
s���V�Eֺ؎�i���＂^$�&M����j��Εm-���Ƅ����;qw
ŝ;v�?��o���	|��8Ef\5͚�JJ�z�T��3p�s/��$R�ĥ&nB+�(�]L�K�������8�;�<�~���B胣��j:Bq�M���gtR������[�G���sY0�'�������kj:.���>`ȴ�Ej���r��>g��h���Dh���ۮ6�m�ْ����ْ��]��5H�D��Z��[Д[�̧��,Y��{��M��g�[����}���=4e�i��#��!�<�\T��ER-t�˲�x��8���\t�)��PۖD5ԍ �WTz���I��A�O(�1�#k�6�gYs�v�E�[kZ����t�<��:8��t�����P�z�'�b�7U).���ܥ���.�t 2�{'̍Q� ���%)ƚ<h��Մp<��: �����k��n�_����(89,�㋨*��pɶ��T��D���f����c��<��hb%���"|M���ÿdR0z�Bk�:Dp�`�$�[A���|ji�;�ߋ]��΀s&;ȧ�%�EPz��]yX���W��o���H�c0`�`eN��It8�ʞ,}wÕk�ψ�ѩI��W]�`�q��[˗)���i�N=��ԬW#�c���]r����2�_w@�K�����b�K�!�B:J�.d}V�i=�}k��+9wV��&a��&�t��6��[7����rf�a%{�H�E^>���tZKx�ˎsH6%�Ӎk�Țxc�:*���^�V�Ej�*�b��@pϝx>��2�ܦ���O٠�)��d9��L!dc���Q���{�Y�E��	S�M到#�4���MFy��v�����'$Vҥ�i�]n�{F�\:�y6tҽ�q������x^5X`כo�`=y2CȨ���]�ñHL�Ƿgc���A��gi�;=�u2(��;VD���Y�]yշxp���ƕ^�b�
Z���3k.�gv�s����UZfǮ}�S����>|a(=��v����ᑊ����g�Hd�9R��S����A�#���f	�4x�d]�b-�>]�V��P:�M��7aS}�Q����b�Lh�F�\�6��«��Lx?G�{#�ݪ��T�-�MX����#��g���gU���z�=��aT�qq�Q�tR���9� �K�_Lx|�����+<ה��q������,7,�`��Ʊ�^��n��Ņ�	�ݞ`��KN{3�wol�'�z��)�0�]&(�9��~X�<e��=Qͪf�{v}�1X�uݹ{��:$��ѩU��ՙY���6)Gݭ��V�V�ݞ,|��a9��fv}���*��<�:ҟy�A�

ʭ.��}�5��u��g�鏹����?xEk�����c.��%���V��+�Xo�:�-��=�!�#�<�oj���`��WIEe �):V�����Z�GJ�@缣#�
um=�Y��CxǞ�y�-L�P�w,��YˤY��K���eXn��/e�E�j�s!�8I ��v��*�^�Bj�k�7���T?w�$>g�js�m�XXN�A��a�GMDu�ë"��f4�}��
�N�2�Zâ^[�4eǳ���9�9����"�x�F�`ON"��*9r�-��R��2X�}P0�ɲ��/�M�E�Xj��S����I���{�_Bo޷x�#w�7��pxKK�����WB��c�fO����Q��J�,�����g�BTS��^�oV1y��Tb��K�Y�"�f�8e���2C���S�kb��<����G;��9V����>���4�<w���p��l�LxQ��.y`��{)��xU��In�w/#�6k!�P�8mȨ}C �q��	�fp�x��i��E� &��M�"�ӆ�û��sM%�O_\�s-����j���'�%UT�/@łVn�X�L��.���)�v⺽���zq���v���r�'��wE}\��*,J��ܲ`�t�o��8'��;�h#Yo~ϊ���l�ɭeb�ɭ�����.]�z�K���la�r�q�'���6�>�Q]p+�v�Rr�:�1�`���@OCW^cET�Eèc��͚/ #���H��K�h?���aI�g>�x�p�3zC�&묹��Φ��G�#8�B��
�VJ�u�V
W�e
���À�P�:��E��<VJR�Ӻ�0�-̈��8��a�NG	GtF(�QN�P'b�H��A�ή4��$$H�q��2����M,���j�n�%�q�>��Q	ѲJ�%;����'eD{ղinv+�X��!�륚�����ڂ�2B��0yx�Da�8*;!{�Z��Q$�e��ԋҘ��`�dWv�p0;�n���[�s8���4C"z��28Lf\����X��.�|�:�I99)�ΰ�U��p�W��qg�q~�5��FUDI�[S�f�׼�W��/`L�9�8S������6��i&T���y<W�mՒU��B�oGxK�(��~L��Dg�~F�x�3uʷc����ږ���u�
N'��;B�ME�X��]%ۊsx�aV#51*qsB��8u��"*�f��p6WsS�(�u�)wOuHw�����\�Q�`�gr�R�d�+7��하�)�o����m
����fP�ڱ�կ���"�w�hl'+�����fp�a�2�Zk?  ��*T�\k�řeb����"q�G�r����c`���T�,{�@2��ulL�\Ժ�0*^jbD�y)�X�rcCܯD�5 �;�vͼ�
�n��X���z���^Ty�N���H���*���3�����gۦF��ۺ}�,�=X�۵�x��&؋�<Evmx��X�V]��ҽ>����F8D[��M���yݾw�ޛۼ�0X��摞莀��r� ׆����jl�1�g+U/id���87���_%�9�K��q�5�*/#���Ej����U�P��*o��s�1U�p^��>[��wy:�KA%y-�A��*P)mP��1J�CՕ����J�M�ب�z��3YK�s�^νC�е�isU)�����K��&6dj{��f���v7�����L�*8RS�0�ob�`m�",.�k�UOG�b�Sn. ��:���RF�g�����T���ȯ{lڹ������P�5�U���V��^��`�t�1{�W3F�@]��γ)];\+��wP�d�`�����M����[[�@�������쬡�G���TM��J�ܺ9yJK�h����;x̀�N��.�JW���eK�2X;�����%t*�(�"�{�,�v0/J�wꪤ�痻x���GçW�G����Q��'���h��XG	��FgJ�6���ӨI���ߪ�[A�A�ז�p:/¹�s֝z��Ҳ;�^Xn���nj��wF�ٖ���Qq��_9��f��:��,}�d
5S�A��{��i�w�ȫ~�;������3�_��V c��A˫+�3^���utἂY��S+��}Ϲ�L����iyGKϭ�OTg��ؗ"(�]������o�i���J�'"0�T��F̻�DH��2԰x&��X����U�w2�ʬ������!�v�_�9׊��<�'�'!̜4���Ɲ��1��Yw��g-�����"䛓#Q©��ge�Qߵ��r ��R���4'ed]@����� 0��d>�΀��QjsI�f�e���{��oT�����UZf��D'<+� mǟ]bz��Ʒ��j_P9Sܱn��y���!&���\��z����Z�/3�dq@നC��k�Cr��5b�ܲ/�˥�j&&�d�v�W<M�p+6��M�,��ޒ�3�Q$��j��{��^3��w~�-�'+�e�:OQ��7y��������Sk&�:gi�����Nƚ�V^�HF�5����Ee�}$�	����9�ژ��>���q\��li�<G�c!(�B�p�2�t�\��V�27.�_	(m!g���}��1����nu���f�N0�܍c�Fk��R;�tB8����"���qbIqXs���s'��\���6�)]O���#w��Kvݩ��@��Ӊ��74�vӎ�vWX�ܮ��^�+���)�"0������ge�����f����8��55�V��uф'䨂����o�Њ�ȡ1;�O�<0:���2��hRۡ7b=��[ˋvO������ͩ�����Y�x6|�S`9(�xƷ7�PTi2��W����OS���6͋�l(�{a8g����pV�0E�}��FhFd# �ӊ��y��S����@$�����n�tM'9�Ď����E�Q����8*�ƽvra�^]�ĳ{�(0�L��z����
����o�>�'���ޙ�4"s�ι[D������yx������6htP#���[�̞�%�kT�N���ݷE���Qz���q��mӼ�4��\c�8�վ3���۴ki�A��{Ԅ�*��Wsp}����e*��2;ӽ�Ӡ�;�E�C^2��W�.:�$֮y�wa�51wa%�}���c��:��WXI��So��g<;�2&Զ��Kݓ��\{c%lWǰ�s�W΋^���=�
ӟ�,u����F�+�(�efO���F@;<�,��t��`���u9X�>wӳ�_����٨��.}]��Z�y-(%|i�5a��H\2%�͈��U�&���Vt�{��u{=�u�mr�U��)X��R��-�PdI�
t�ui`��>�'N�����-�����4K�ޢFqtziC!�e��rՍ;�7\zb�H&׆��z��:���n�[�O��}�D���"�֘�B4D����j,6��nQ]s��lE6��M�P�;�;������5�b)D8���Ϊ/ #���K��G�I�g>����D^���H#z"�����Q"��%�@z���
K(Wd�w۲9F�5���_r'E����ڦ�V�Xv+JNn w�(=H��"qE�e�5�=/��t�n+����P��u=�ZkXY~E�ҏx>�gaf����������Lg����L����-շ"a�7���},=���҈���gUmy���bad���
��0�1�5>�DIS�3+ޙ���'u������ԡ�[��ϫwe�Z5�kGV�NX{��.��@�̦�:'��|.�Z��ً+� �͛]:tⵗ{�u@v��Ȼi��)b��3�|��ݵ���IR�#���o�F(�dۢ��u�'(u�1�/
������fn�<ڼj�(�N�����M��r�Պk��l!>�6ֵ��|-�;��\u�jԥh���lQ�t2��)��l�e�ܳ�bp�~s��Ƙt�Z%W`N�,r���s�M��d�i_�gzЬ��	�
�4�Y6hc����Jrw����շّ�	Tx��#�<�;��TF}���o�c0T�P3�dzv�8��e���V�ob敜C�t&��C+ƥ�A����I�����X h��5b<{��3/���2�v��sg��x�)�X�q'@{�蘦����ӶˈˍQ�i��#����r���� n�/���{6�)F�.8��hy�y�3���H��0�3>ơ���.�q�����)E%\켉ا|1�Y4��ێ�4]\��N������D��p��sQX���kj�'��2�ă�z��}9�!��B5!8�j��n��^ff��m�n
�O��)�b;K��{��a�^�Q��0P/r|��-*CS�n׹y��=b�-h�U3�E��Dq�˦oc9�Rx�M���r:��@\y�F�;f�v�0�+��>�&��8+1g ��DZ.�|&W�ţ�'|�ަ%���TMgC2�����F������x��<��Ѯ.e�A\�8���j]����(A��[���(��I�F�:�wt�Hq��w�vU���8(%�(����ֲ�-I�q�-�ՙ9m���\^uޙQ������X�[Ҭ7�v�;�]��G���O:_]��n�P���c�KvmtR6�R�9`%���{n���*o ���VgV�S��7+����Jx�%tt��b���]��atm�b�I�YeV��e�y�>�.�.O{� $���q��� ��b)e�,�.�8�����v�76���lt�<�+���w��R��X,Ͷ�7F;�t�ݍ�G㝊���!SU@n��ȓ{�u�J*����� �\�w'�`�%Qi����j9+r����P�3_]��By��\�8j�2v��CH$��]8f�!�K�{;{2�VQ7���Y;���������8�rK.R��+]Fٷ���9�B	u����[6����wyZԫ��O;5^�1��ڿ	�ҥ�fc롙���r������+�M�P]@��`�/������I��$� �<���G��8�qPr�GIK�:�.��b��wY�Z*�O�@6w7������"�l���)����ćݸ\�gm�� T's@*�خ���u�mB�Z�Ыγ��-�G���q�{j�������Z���vS�	�g��1�7�	i'cv��X6Gb�Q�����ݦm���'��.�٠��r���a�q�f
�R�Qՠ.ͬ0�v�կW",i���(�)�W1E��s�k�S�֕u�]qr��Au�
_Մ֚4/��U���&xGʖ*2��dtZ�R���ە��N�إ�X�3����c�����7#�VJ�ŗZ[4b�����k�������ȧmᣭ#��x黦��DV��w�ũ�i�WWϘ�cC�-P��u@Չ�8��R�Ժ����,r
�f���n��0���hQ����; 8L���1���] ،[�R�feq�4�-�$��nW[�V7e_1��>��֒43B*��-J�،+\qdG\ѐLUZ�֞ӿ��ݮ
�U	���u(*R���N�IZ�3��XC	�����[m��7�W���J��ѫ�#��W+�[��9z�����L5Vfcu��z��"&gp��	�wv3s��o��7w�e*ɻ��Ϟm�B���y.Y�B��۵q��솦�0
�709y�U�Y�j�[�-�v䝭	`-7�P�b�v�	�z���N�3��l��U��f]
!N�T�Y��݃Cx��ވ��n*-�#:H�e]�:�.t�������+��Q�+���^C˼ԁf����L��y�Ḇ�ۏ�K��w�7g^�&���մ2hT�9��/"�I�8�@z&n�A뾷L;�6u#���UP�l���lP��	(��	yxV��PDԢ1���YUPEF���-mTb"�b����U�ʪ��1EQA����"[*+XV#V1*�**��U�IYm�Q"�Q�"�((���QeK1Ub��EUH��b*�*�H����)Ŋ�AT�QU
+QEQb21Pc���"����PTb����b�����QP`���H�F�
���T`�Պ*,cZ����Db-j ��U�X��(0Q�Q�e�*1*�j*1Tb"*��P��)*X嬭X��"�J//HzQ䮫��5V�z���fl�ׅ'�}���%�&i�25�^g	��z*�;���y�wA�;RC��T�[�O�T���v�Vسv�l!w�pS�5ʰ�5���u��b��f�\��J��X'�3�*�@��P��#�	�fķI�o����3�
:<��C(A����$��*���3l{��E\�`	N8�5H��z��V�Z괹��Px�@�� Ij�������wޫx�K&�)�7(�`8j�����u
.CyD0xm�X�{[��y���s�{k��H���j���om���iª4�����6��y��ۚ���a֯����1�=�8�O�h��Ҏ���ZJ���Q�Aҡ�r���<�.�fN��wX������|���|-_��v������q��әc�;��Vo�F{}crgu����eY�(��{�Ҭ�6��x�S����7B��u�)��Ooʬ�Ч~;[ٝ�� 1�(�ݚi�k�&,�;��+�Pua�YMg�F`�b-�Ҍ��z��7�X���*�XD���>��F�wS�g��'��ȗ��7���hawG�<��-Cs��=�:n��E��0Y�J�4ybta����5��@r/h$���"�pVĕn��SĄ'8��.݃B�6�f*��/a,�4�ptuX�xOhV+==Bc3�]�#W��җg�QQ�$g<���K�8ۓv����{�򏈮36���;�Up>�=1��/²Q{�kM�Ν��1JX�vl�G���e`E0G����c�����.$+׊�V�X>���u�L�	߲�`+�wU�0��s瑶ɍ�ـ��4>j�y_4�k+g����¬şa��+� h[�:�蔡�0Td�:���]�Ť�Ϙ�������G(Ӽ�Z1�8d�1�eze�(����lj�_N�g$�vȅӤ3��\b�qA�et����_%P{Y�k�zNB���y�=��n�&��c"TQG�M�jE��v��k���C���}���6�$����VV"���.{�f�gl9�8�U<B�S�t�߄Ѝ �)�N�ͅ�8ױ��9wi]\*�G��%..�Y��f_������ѢmD��k�]����Q~Qǌ�/�T
���d�2���:����ܟ��7|豪
h�7�S�#���BĞ-��d��{cx"���æX�]�����g��J�Qb2Q�5��PTi2+!�:*�֜�X��cor�J�md�Ν�V�q�WZd��M�;�`���F�kKO5E����
ƣ�M��E5jh�"p9��.���_��w�jv���<OC�}��p2��Yg�s3ax�㝫�+pT�������iV�˳9�}§U�~���2�5�d�2ι�SuFۆ}��Fkљ�x���/&oe��kR�7�t��d�@�,����bG'dg��8��7�� �,Z�ӾԬ�JQ 9�;�us��u��u�Mf�2; y9��9����!��^C�j����A^x��l�����b�Q�*�]at6_D��QqW�	��+��gJYZ�fZ��s1꽏S}�BP�YT}����lX�k�.�w��*�P�o��W/Q�s:�ziӜ�B�Q�x�}#�WE��LV�Xbzn����b����4j��+�]�V�4FL�f_-��7$o��
�Y��l��=��(�Z!g�ФV1�ǅX��Ykw�T�_u��rI	���d���K�BQ*Cs"�vۤc���L�������ݑ"�?!Ļ��'�K�t\O@*�i��#�SS�:m^���k���S�H�R��*-Ug�r?ov��F�?�¢'L��9MlzZ�o�"z�t$����;ʽ����mI�^������O7g@�Ѫ2�tj�R�&��e�u���/��'��O��8uX��(x��j�_>C�e�1W�W4�[�E��`t����oVu e�t*=B�*r���yGq��R:Qˬ|7ca>w�Sn��3���L|L��x�������%�ʼ����3��(WVSQf��<Q���^f؂";�!�Uf��_n���qF����9��(=HߧD≘.������P��!WU�:�u)�������ųҏ8Yz�+Ƀ1mχt#��G��~�/ ,�[k��^����T��*}IJQ��.�D�`��y�W�=�؇Y �*`�B �Ug�g��.�]�[z�oF�ۢUx5C�l��M��;�n��g���d�	��1��VL�W����77"%�S�5P1Ex�U�Nc�x�ug��D�f�t��18Y���������'G����<&h�=�u@�����N ӷK.���Y� ʃU��H�e���%|������p��[���j`�*\r�R����-��c+5�Vǥ���3�L���:��b)�aE3m�P�ȫ��Tٍ��34x>�{�6k�b�P3M*�p�5l\��I��Lfu�;�(��b,,��=��L5 �|bt�/��&Yȼ�����-W
4Ү���ݞI�f�*�������[o�*NO��%A�m�os1�,���;�/�i}S��o剈k��4i�U�p���^������i��h�	����u��1@�)�y����ۤZ��-�c�f�u��l���W�������7´\au�g/6�)F�)� �W�j� k���F���=�z���S��h��]7'h����a�C�^4���P��z]7����
�J��Xʣ��-��E����Imlr�}Y�B")���o��K�L��WT��HU�U��U�9a���;Y��i�<���r hnGؿ8hN�a�'���T�IFVt;���̪�k0�z����5�ܢ����G�M*�0�Xs<F�G�����N.!�6"n��le+�Mn�v�/O8��r�^νX�.����y��=�>�n�=w�v0�>M�o�
���(l�t�-��Sb�g��C��\��mJ�*�#��G_����tO.�V��� ��=(�z4��_���W:][w�h۳l�=ǹ�WV�Ѽ4�_-�A�0�dW���)����˂3�K�bJ��4Q��էl{&���WW"������C@��O�8��j��G�s�@XU;�������=)�����^n����N�)�7ޱaV�vL����PV���l��aWZ����|�������{��	���Y\�o��&A��~�	*L�8�;rE��S�X����n�:7�
+(�Qv�t��q`v���3u�k����Ƽ�u�1���ZS��Y�Sƶ$�B,s�Ss@�Y~l�I�x)����b��Q�t�ؗ��{�oIo'��[����Nvx]��CW�O�y���^�[�J}�1Ys�k�:�S�h����z${&��=Ё���~'&(57�,����^=>����{]<�:7̥�)��n.�uF�N���{Hf��0h&��X��w���^��J�,n�}�十O�V5�-'�Vzg��j��G��Vj���4[}X`��1��:�����J�Ǘ^�d�V*�,+:#j�.���)o]1������-���zw0�٘��7u����y�_�� |�����Bd�iϜ����]Ml��6*�$��(q�[���P���.�����*�:Gz7=x�:FD Ynfgov���^���Lj�2P�`�-�^n��R�p�8n�������p�ŎJ��c�F���_A�䨧R2.8�V��M�ֱ�#f��T:Ӡ�u��)�UR�Y��f�b���*U��:��{x��t:�;���lwc.�Շ56)���nn-�q!wY�#��0^ҳ:�h�sWZ�+.<;;�عN�Fi>j�e�(��U��h#,�]zD7K��o'��W-P͗�EN6/�pfi�����|x��׶�1�mK�cA���d-��nQ�����N�q�,�k�q뎢���ػ�Q֡��]=�������T�1aD��)FTV�U4EDj�p�
4�����oː��5m������\a�C�.�
���x;c��LN�,B�AGu����v�{Ns��ʵ;>��Zۡř�}h��W�>ȩUY�F������of��O:iF?E��:�����#�8]��Y��S���2���P�g�^;(�l��sm�<����߽�#wj�2�0�q�tM'-��9�"Í8�&*:��]!�(亭k{5o#�C!�:oJf�ְ5]���ׅd�O�J��#h�@�e�W\>�i!�^������.!^=��T�PU�B�x��aY�M�#%�I��)����G�d���m�ك���Ѱ���M��V�I�}9쌈
�@8YYc+�dZu[}�UO������s����f_u��M��ݍ뷈��v�+�h���+�O�l>�#!���}v���pv�}J��ܫ �wY�ݷ[��
���`\��z�5�����)aO_sڽ�k�<չx��v�eա�a��)�9��ͅw�1���{9]�ה9�|�D_V���}��s�^eowCV�<ܒ�W�Z�S�rt��v�ݢՕv���bHY�8!��,�Exo�\ʵ�e8=��y����
�R�e&y>�2�;���wغ!�nX4���D��tӆF�܊�{�U.?c�����X��0��wX�o۽�pO��8�|��倿�(ѿL&��M��ۯ]�9GTp���bJ�[]vtr���nh����:`�U5��j�|���v>��?(>����"e�c��7�#�*����}��n)G�
8�,-�|"��&)Z�س�6�8 ]:ĳ{�<��ؙ��k�L,AE�v��Yw��cF��6��֎��W����m�t�gU�ё��%�{z[A��<i���.ٵ��9m��\o�~�"����"�q�QM&�,��w�O��ݦ����&��K�y�]^�'�(�8Y ��U^�}St�nr��Z(q��쇵$�P��1����nv�G>~���*OV�!Xi��7k������=h�$3���̄��*���e��<đ����w���^;y�6�O딬%�9`�Y�ԼW��+�/�G����^m�#�����A�w7Ӽ>��?V
>���|�y{�8�g�g΋�+��Tz�:a+}5be���H����3@:Z��g#{�B`k;0[��Ԗ�Z5oy��v6
�XO)�*�ڗ�o�/-[�,7Z_̣�:x��ǆ��s�gw)�W�if�G�'���k��Ɠv�MX��V�Ytl8y7@�p\��2��i"c`�c#��||�G�50w�.8q|W��{�՛�;��~�"����Ml�!�}ڕ�Q���E_�X`�L����k�b>����J�=��RX /�/<@Y�N	^�=�<�Ω�Fق��t�^��l�6�0g�e��,���B��Tz������
D�SVa9�/�s�ʟ\K=y��J3`S�x�j�``qyO1�A��y�f������3O�܁�pJV�ea|F_��uf�X}���:��o�{µ/O�$�����\rN[!�����*�*]����V}`w����S�[�$J�����~���3j��{v�yFW�H�`�]CUN:��g�bvx�/#���C��$ˈ�9*��6B��b6��`*��|������$�W(��#��*P)_m�k�A]�ݬԗ����9�|�[��}<R �cR�w[ͣC��g����ĕd��M3p8"*.�*i��9yٍ��\��ur���d���Xhq:�cq��o犬p˾�8��]�;�Wu>k�I�$R<��ܾ��0�oU�r
��M8��D����]�Eyd��8�ܢ����ʧ��jWD"Њ�a��v�=Y����6���H�%�8)`k�D���F�e�"P��_[w�C�eB�ٲ"T�Y:����o��܃պ�?�_ux����{�|��	�,���0�Q��=A�T�i�fT�(7���Ʈ��O�������5�@����Y�H�0���zf�냇0}θM>j߅ß��0����΄Э�"	�N�;�ta�*��b�z�F�H��/إl�S�����sZ��!�����|U���Q=r�<����hY�w*W�2h���	Sn�2i9�~�
,��U�F��2"�����&�ݽ��S�M�/	����5�����o�ļ��,���C��q�}j��a�ǝ$��LИ S��v����P�U�^c�:V5�Vj��u9��sg��d[��Τ����EJ��uׄd�8��W���
�*�g`.ؕ������%�Vn̩P��6�'܌\c�)(��`���Q�;�:B����ٙY1n�૬�6���Q�WR�ޫ���m�fQ�l���oe��D�ə���A���#)g��|�D�\���sU�[\ ���w1�l��k�8z5��[5�iM����Kv^ܫ%��1|O��(k�ؾ�uwG�Y�/,:�\��oۈΦE�1#��ZƷ]y�ת�%�ԡ�J��7���`�X�u�Wma�  ��9V8nuE\5k|ڮAS�O�Wt�y�B|xV]f0d�Y�eKE�rW�qu<݊ЪKn��Ґ���a5�@PE8g
̫��L��X��h�h�,EƮ�"ۃ(�}���4��dO_$Q�R�V%Lo9��@�%e�y_gE���+X�U��M�r��x�Vfp��b��^��5PC�b��k/�����ɵx��@��_�)F.�}�N,_|���Y�f��T�o�0w�[G[�G)��
��C�f=�w�
��Թ;���b7��[�me���t�"���.���§���
�ٺ-��<6�Cs��á����(���
7�šT����Z�+���(����|	�t%�h �* t��]{�U�j�#q�!�!F�����u[|i��t�^�[N��;dR����Yy�kTޫ���������
�A}"�ģ��$̡wt6���m�gT'��������Rm[姻�>�9i����Өg7YeimP��(=�';:+O�]N�n�,�o�����kX���rQ�uu(vd��>��|�@�*�Xwo���+��Y�Do)YU��}j�-=0l=}]�nܼ-�\����Q8���0b��j�t�|��I+Gl��?�J�Of��b�7����8���K˟ZKm�Wʠ���R.���dp!Jdk6U*�$�Q5��oE"lҢR�*Lw"����J�ie^Q�'QQH}����Y��q.b�'FP�N]���4�JJR��"��̮Z�A�!7��E�#��@S3��*[���4or�������e;��-&=B�����YR�-tK�	Zi�c�^]���i��\lf^lr�<���Q���-"�jErb��L}�ٽH"9��+I#��.O�Ī2._Y����T:R�8s��Hַ�\۶-vm΢a����>g��X{�Z��*ej�u�b뽇9�1�.��O�[�������T�Ѣ�+��MA���昍��NN=Y-3][�F�"��{w.+��T��� ���Y� �r�р+`R40Ve�8CV����;C&.�|0jO�jS|i���yW�-Di)3TPW�J�*M��]�6��Pbm%�&V�Af�ڴn�3Xe#�2"��3h6ج�,��(֨cq�,[h�(�1�j�Qb(�n9�TL�U�TEa�*H�I�1�J����Q*!��`��*Ƶb�ʪ�Z�U�IZ�EV�ȫ*U��X�*"���Z��"T���[U��`�	DJ��Z&Z(�����1T���TD[j�(�(�("������R����RV��Z%�TD�-+-��-l�[R��ʮYR�F$V֍��V(VKj*�EZ�Qj"�F�`T��ĵ@�����մ[J"V���E���e��QV(�6Զ�m*(V\����ګ]�v�		�|b��q���z�37Pj�+��]y�f4��f�X;	��c�F�-��b��(U�NVH���Z�ik�&��[��L��u�������<�W�V�N��\�i��T�)���{SݳO����
�R�.Ӈ�<���z�w��5[���T���H��tT�ʰ�y�vX��;�.��g�_P(�mu�5�"�Q�0z9V8�8et�8b�Lo%P{X�5یVn�c���%�f����; #7h�R�\&�5n��3��:�u��k�U
�>>XT�r�޹2��ՍP���8φQΊ��B��m�F�@]�Y��r�#<Ve��hB�������۽�������ͩt��Q��6��Ek����&�uG����m.v9-ާ�&���UE���=��u�TAL�,�t!{��^1���S���5��9��6�;�����jG�#�3�w���&��1UpUMs#�\=��Dn�f��\��3����˥�
��o��{i�$Z��Q��f�'���	�iՙ"��>�b5�N�l��H˩ybD4�Y��N�7��D�s��#�9�!�T��#x� �z�D,6 Gwe�
GG���It���U��e��[��,�0�jS7�J��/a�$����3�@��(]�x����15{p�Z��zTD�v�ޭ,z�4�@1���b�^�w1ynp�6�\;Vr\)�_U�;v�hSu�{U8�kb�ӡD�+��xVxҤl_�޽`m����E�6��@�N`�k�/�Gq53'-Y�O��t�5꼙�����@U=�W5�8�P0ڜ�/a�i�R\V���.��8$޺��]�)8�P`�>ۢ�+Me{����M�Un����v�'$�np�+v%%�D�U�������eMZ�,ߛ���kjMy�V�SSf&d�d�~����.$[z�vr7�u���hd�,!���>`�^�E8�Ƿ�����>�H�'��N.VY�l�Z�.0�3�8T>�����<�QdH��j��w肔W���20y��[r.����?c� ��"�>$��]����g��5{�ҨgO���U)�u��ߢ$��[�mׯ3 X��T�#"i��>#՘�s;l�^�����m��t�鉮��RqW��?v>���#<\�#���Φ
V����n(�@�k8�E�8E	�
W�+��ME��î2�ļFmĪ��j���iO )�,�C<gر��=���OR�X������%wl\t#RE�����ڣR��)�7G~}�n�0����=�\vU���c�!ƴPrgh�|��&���t�*^�~�d�ë�' ���:�t����owP���z�Kt3o5��j((�wq��d�J��UJ�w-(�E*��9b��`j��"�Z���\i���~qԋ(��Z��Pq. �wJ17k���FEN+�|�c��c��u�kW�����v-�����sŞ����d��蚞�cL�8�����Q=X0΄hB;!X6]zs�	��DH��n�F���gp�sji�R���5u��:��F$1�0
%��Ô\I�(��qP�'2�;��V;�ǂVCiz�Y�3�ǨO}Jӱ�����B����p&rB11e8��h!��K�f�d�rz'�Sޮ�.bҢz1J6��9���]�c�Ls�t�Ë�h.�+�|��4�{+a��-G�ʧ�EZ���8��I��dC�����Oh/�l����5�鉕[O�ި�6`�G��2ŷzll7�CuH��LP{�蘦��$fQʵ��-�ܫ��q{��8����� ���ڲ�eH��z�i��f����m^l��U�[�`L܄�^e<k�.�^s!t��O����z�����=��Hᠺݳ�ά�]8���oDmD�O��U�ъ&R�g��e{'MW�a��mK�f�~��,�������9�9�M�scw�����u��M5�Q=������K��35@0,mL���h��;�E^��݉Z{$�˩�x1�k9��ڑ̵��h)���ء��_l���cx �U[�Xݭ>�w�;�"'�V�Md�=)������]l8�/t;vkS���D��*�iv6�0�aX�3dGv�Į��n8���q�l��{���1���ڙƪkjF�mR�
�ܳ�W��=J�Φ�v�TeU�
6�:�B&�èU�94W�f�Z��+�D�x��1W(F�\>�+<yרcT��u�����z��ToPئl2�U#��J����CT�w�U�W�M�S�nQ�+�z��<���\A9���zӌ�g��7�cF�D
=(Ս�ԋ�Q��'Kٕ}/9R���^��	���7v6���'�W�N�6-Ă,�������Ɏ�:�3xj1`��ɮNGv�5Ş6T�t'���U�:1�0N(�\�$�Υ�CP�]C�ɝ��֤)�?;Q��/9���NS69�*�uffr%
��	��|��C�[��[)�W�#T0��t���p(t	)��Cm9�pE����N[��>�z��A�ҨU�h\����*��M�R�Ѽ.������QQ�}��b��,~�蹢rL��ñ�s�සm�.S��t�g�f�M����ޮ�����I�Z݁#�c@�VQ͙�-�v�,N���t�%w#\$�Ɖ���y3rpΆ���+�^�IB(n�q�MTiӇ	*��;&�ͳRgU���'�5h��P~�8��$v�����<�X7�%5c�e8��sgM��dFl�Y�,�'�":��lK���N��;�gD�b겢O��e�� +��v�Ǡ�B���x�X�y�8ãz|��aJ{[{��T�᫯L	���E]Q�'�8��P/#M;)Z+o�~[�W)�mg����N�'��͆���¯;n��M*���6����D���E��=�+�Na<�v��}/�$��/�G��ĥbz��P��O��<Ù����{S഻�ZE;�[}7��9�c���
5㥃6��tȠxʎQ���_�N��m���ے����*�@���a��;��B��H��7j@FE��w2�0Sr7�c�F�t;:�r�z���[�:�uw<��U�ra�ӘS �Z:&����s������ؾ�|$�]����ߞ��ը��xt�Iiw��a��́Ɔ�Q~X��R�1�D���h�Qu��]YF���+tz=OJ�,�i[�δ��3����N����o�a�:#՘���2]<o�]"��5�q��.�R�pn���4��S����@���]H�{0��\V�0�9Ɋ���0��y�ݮ�(��o����rvt�Sj1���r섞RFT��aev��de����N���`����q��mS6{v}ֶ���^�+V�Q�`�.��G���Fi��&,�P����q�R8�.����u���e	�V�c�u��U#N�F�qU��_|�)ܟ����Y���\m�M2�48z�5�Ù�eZwfH�ˠ|�³�����(�>��噘̄vhJjp��̯eǷ�Js��#�'5��yN��iU���`�����O��8�G�+��X����{����:��P��1Ź3ٜc��y���
�ky�B�hD���
�@Ŏ�t�X�V���.�VD=3�I��S�ȭ�Q]�i�/�*��u�Sa��t@E+,߃���UxE
�W�Uoe�q'"�UUoyz���ꌁ���j�`78}^���Qy��V���ˆº9LsQ�S������򩞬�P є��!O�6����򥑾�W����J�'��WL����6�u�U����+�q�lAJD�dhni�mȮՍ;�C�(NP!���U�0�	�#�����jo�to����Hl�n����K���4��"=�����38�1�x�g������,�J�B�W��P�/n�&���r��&_d��7}��ˌ!M#���i<��H�qE|{�
�ơ�2t9��)X;Pk�j�A��aq* �S�6�xDIM� ��gwt��t��5��s�~ǒ���]�@6�w^/��xN�L�Qc��5���ςRiف5����5y����)��a靖�����F'q�"k��0�J�P��aTM:3��G^�僫���PY!�a:e�b����a���ޝ|"�W��P����;��w�����$o��#��m+��F|�kM<Y~��8�E�b�dAQ`9t����n\��z��ےP8`�F�*h�s���:=;�� �x�Ȱ�3V<Y�yƏ ���75�oMY�{��H(z��q,K߶�Bxo�&�@;�}Mgp�\q��k��LL�,x�#��w"�,3`��S �.v	�h����՗i��ڮ�,��c�*��7{��Igu�=b\�p9�N0DM�f<{L�4+(#S�HJLN��#b@0�\���/���r�|D!�/x[	�HNQf�:��c�LsF(R��l�+}�c}�۔V��CMfp��!k-S[f��� C+�\4�p>�F����o@ow�P������!`s�7Z��K��P�����ܟ!�:����V�5�ge��Y���(�fgՕ'C5�6*�V�*�əȓK�Y��oz���9eo1�v5�X5�#p��w�n���!��V�X���7�![o�n����o,��ޖxfdrE���;kU�$js���=`eKpj�}a�@�b��BKP.!���3<b�gpU����j67��-u6�J1!LL�SW@�fi�Ä YbԆ8W4>���=��Luڃ�úˣjb�P�NPӔL�t�K<lJx��[V:�t/i��`�ⅵ^8��j�ڐ��g�I۱+�P+/j'����� ���Ⱥٴ"��<F���-��"�r^{<���h��y<(�ǔ����aW�K�W��v����x���S��Hoxa�QM¤էh�v]�X��$Q�B�j���ĩ�(+US8`�s�6/�>��� z �յh��m񾵳�o�|��R!�MEº� ���z���Kt�v�|u$��c��Z+W#;�9�>>�O;#`ɧ�+B�V9�U�,ʵ���J.�:�cT��u��n�u�7���J�\���U3s��&A-B����
�U�Rɽ�q��D;+���^cQ�i�;uϫ]j��;�S��;.(�1�#^��X(�l�[��Xw�3��Wv�|�%Xҵ�����W�	ɫ��S���];p��τ���>�r[F�/L�Z��w�E�Ju��ت����Q��S��.x��Y���Ԟ�K3�/���J��/f�݇tN�4�4���=�ןW�}i�.������X;8���*��j�1[Q�0�`�[���Wu��r9^C	�N;}Q�^�6�R]�tATá
��̜QU�WS���k5q�p�6��Qn�z�Ү6�D�� n���ka� ��s��'�7F�����d�%5΍i�Ь�t}�O"VQ����.�}Ru�'��Ӫ�Lw���d��y�`� vz|z Sw���^��h+������S`�E�O���=C��Ӱ��n� ���f�����,�>��ݲ�_k��MX�N,�l<�^U^>��=�3�a�B;��tg鵅�)*�����{�^6)۫� ��!���b���^<_��>-�0�ל��r��I���֒�0[{�8���:nJ~Ub�z�B�!��l�_���7c;6�/+D&OlZWL��l:��Y�i�h�Y[�8t�f��¯��؜���b,�YZ��,�Ͷ�j���C�O�E�kw��-�~�!�ݍ�9R=����D҇��~�B�%���uл����V����9�!�0�&�b!��iH���^����Ӱt��e�L;�ȣN_[������Z�v��9��c��n�K��t�!7Xӱ��:(Yٜa���dϳ�(��R�n)�����==�2x��w	/-moQ��O0�bt�' �7�� ��Ծ���Y<xʎQ�ۋi�o�θ
�-SXgi��m=Ňf7z`�?��='!]Hυ��ec}������39cCRq����v�KBR-����ό��Z[㈚I��_j�|.�wB%��0k��D��A��r����]�k���>��A�D��j/���ud(�B
(.�k`�Y���hQ��5:��J(˩��T̓�GX[P
f`���b,�"�(�z�6g���	��Ҿȸ]T9�p���R��mH���w��>�5{e	�S�}��n�Z��jU��0ǌ-S$��4dVExJt6���6�%����j�qA��2������KCFNĕ�טW��y/6�s!�6�j ���7�I�b��v5Ev�C[ٔ��U���ɓ����(g�$p_N+���7o���g=t�s���N�(�"��,�n�#3y<f�����Љ�JS�!"�q�
���Ǻ��UDZyu"�����:�Q��J�Ž�87��am`iިC�{Y�c�kG���sw7�+'��{�cޕ�ٌ�[�������ֵ��3X���\���Wŵ��^.���//��P����6�mwX/0<C�[⬷H��jz��ۛcN��a�i�f�B,�����+�v;4ٜ�nt���7E݊K��BX4g�T|��+1�7�p����&^�7w�Z*�m�Ǝ�V��=���8
锫9�{�ջJ)̷}�������`J���y�޼�2�8��k뤴]7�ň�9Y|�8�Įм���*�56V��S�y�*	��I{S]e@9b�k��px�꽡h��#Hm������ [D*�˶�^U���«���a�/��.Nî�d�G�����z�b�{�?���{u���ꍗؕ�#�S�&�6��d�t������+r�J�b�K,��oJ��ƚ�C�+WU�t� �ׇ�/�ޮZV��}�0���ֶ<�!{�|/��u�ON�[yb� X��T�t��Lm�o7��N���6MJ&�+,<��]N	�)���̄���ߍ9��S�[2^ߩ[��G	]F���u��L�!����9��U:���z�+��������HE�d��Zeݕ�j���S��,���/,���fUt�Z���ϟd9Lwp�{J����5��K>8-���ݼ�śe���%�$_�j��\�+Z�\q@�T�/��J��&�σ�zST ]�jgW8��~��Q�>=��	�y�:���tT�n\}��1N��(u�{Nk�M�׿��B�u�+�ؖV�DX���9�.`UD��3�;��yg'����a�� 㮎��;7d��u���%	H�Y��n��·^�[jeX#f:�օ���ں�J* h��Ƕn�o�z�]�tS�c��Q�ݷ�]�a�ڬY��\8���:�DnW�4_f<��פki�չ>�>��*T�7\�0��\�wE\a��buf���`9ؕ�Sl�X˔�v�Q(U�H�л��T���3:GǸ�v��2.����v�y����v�l���0��Y�bf�T��0B\��*MB�b[U�,�Y�h�W[��s�\�ʙ�*�b�u�ݬ�QM��ZFTUt�]^��a[%q7�U�2���pǲ���u�Ԕ&�)��
a����yÇ�N�r�p��-�U�4�&7��8�7���X6�bVR�MA
2Z��Z,��ҳī͔��ޅ��'r�`�H��1�g�O�p�玡^�sNQ��X�^��D��]+���)��������&��R��V����Z�R����鍵V7�5�M�E�s�gH��B�|ja[�u�L�[��Z/��r3�,���>��ys-��y]:e��:�*�vg�X��V�=.��;r��%���l�z�L���=�)����VI�*V,�s��J8^Vד�}����H��6H��Նh��ף��R�8��.�Vch�IK�f�w �k��yR��:�XM:m�f��xC��k��X���rw�i����'N�߂�4`��V6¤Uj�E�Qj-eklJ+B��"��)Z���AFЬD��X#*���bUkV�˙X*֤R-ecQ��XʋDTUT��ZX�j�Dj�k#�P��#QF����Ubŭ-��b���-�kU*-G-�s
�і��ekD���� �V�U���+m�kX��J��VPH,��a����
��EZ�m�P�U�ʕP�P"��Q�`��J*cU1R����T�THQę�FZZ��6�YUE#����J�Җ���UQZѕ�e���U���(V��(bK���	mKl�)iR���m���j*�T�̸!T �K��ؓ����]�bh��[��6��A$X�鏇P&�$��܋��R��Wy��W�p��ó�ח��=���Gc��Z��X�u���U�w�X���qx���'F�)Y�up�Cn�e�58�K;�^�#�Σ"�t�TеvY�78}M-�6��T^x9����8�2q���ඒ�)BDK���0֩ä,0ϖ���8��m������0��؋�Ƙ��Z�,ٻϰ�/����8v�UADa@�ΔIJD�d?74��nE�`�$�{���[y�u��z5�ltBN���]�>c�U)�i���P���)�΅M��3��KI�r N�8}�KpR����-'ᾠgb:0T VOUB>ʹg.sHE_B�����@[\X�Z�h?M�����6�u�q��Dq�L�2�D
S�+E�[q8�f��k��L:͋7��@g�sǊ~*YGU���"#�ykᯆړ^݃������u»E�6�E8f����B��FB��4�,�p����W�ge_;$q�r�hc"�3�O`��bb�:�ѥ��[��,:)C��_�����3��g����Y�krWn�(�,vF]Ib氹�r�l�}�T�i�;�c�=G�6�Ѳ�֫	:��T�wXM�(�R�u�+��.c�[YW4Q��C�N�C�j*���TM�����r�b=��hoZչ�+��δ��M���Rgn�y��m<�]�K��j����nǬ=�ӫ�P�
"0�p�
�
��e�T;F�������{��n�a�8����jy��d���ĸ��2F(�1�s��V��Dˈ�mJｒ@�I�l�<
;0�l��#��sXY.�Î�\�+��,�W��k3|=�g`ӝ�\m�|��;�I�R�; ٓn�P~U]���7��L�K���V���La���h�YTY��Åy>��N"�u�L��s�j��G^��vg������xrG��Q��=�]����3PqB��,6�#%�kն�0����Rf�5a���������VS�,�J�:Q�z�L��ȳ��G�窺�N�̅��OZ]��[~ՋP�o�{Th��m�b�憩U�����s����niN�5yB%3^�A���&���^FC��̅���� �R}��6�|����د7�rÎ��皫J lö�^|�l�yW^[>�^�i�ޑ��"�*�z�!K���QN�d�,}�*�q-N�:��eiso��������Z�!�Ό���I�D�;���X�� ��o_u�T��J�=�ˀ�祗+vQVS��;:��v���
�1�\g�۠z� ��ԕ�m��t��x.�F����t�1J���jX��k�R���6��k�%m<�M����K�����������iۘ��a��<+��/�e�b���s4�P-珽��oɱ�\�ҁd'�D��'Ѱ���B�p���;J�u����U�m,���j5s�	���)l��1���i�ۺ���$(8�h���e;�r��v���Kx�v���#�Jd�������*Pt�;��xT3�す�Tb���dmV��h�-����ھ�s��׀��G�9��5/j毱9�`���{ڑ��ZȻ����i�z�w�r�[N]R�<5��s듘nq��&t=�U�ÏZȟe'4;��ɜs2�^�a�F��;l�^̱{Y`��vYS���Z�fL�q>�9�Zu�ݹ�����l�p=S�`4ī���xg�YuG�Gw�=In,���/�Ԁ{�U������;M�݁����y���\6���oR����%��Q��8�ފ� �V�Q���Y��Ba����wg%B���.��3c�����)_e�bD�=�{�u�M���4�YA�:�����1] g�(��댊�%'R��^$��ZZP�N�Xi��o�"^Q�ד��v5[Y��-�gǎ�g5.B&�κ�X�[��մ�1�紣5��Q�VQ�c&��MK݉
4;��wsz�S�CZ�~)O��M`n�[n���������m�T:�9uGl�z�	�3�*=+� U:m�ΰ�ڢ��;��x)��R����?,ܡ��zF
���}.��dnbo%�p;Glot��\�j�su[�]L]M���8�)㋌#���}�A��"��5t��r򁅥?xW$�Vr]ɕ�OV�Xmي�lO�9T`���9<��D����|�jq�K���-J^WwP���H\�[�,��dݧY�7���@�ݯe>yo��t���u�I�w��Z噢��,Z������&�p��7�&�x��wa�0V�&f���cCss���6>�Y��d�i�4�.�����㶳��8���3��ޫ%M,�uuew
�\���8P�`㶂�-��M+�U���u�0�bգ�8�Dr�͚�.�&u���+o�*��y39Ԏ�@eaopU�[�m���.��^=L�ȼ��e�t�^�Ɏ���uĉ�P��K"�=��)�YK�-�euWFFT����n���Λ�#��z��\48�]��Næ(� .�s~��Ü�`��++��Z���
o������МN��,�����m<�jR�����މʹ��#�&Bד@5YA�:���{X����tTΫzf�uv��:��J�2�9^�aEZ�M�-,�{6j�doh�7A��3s��5IwJ�Z��g:�r��3T�;Z���9�~k*�K��&�f��MΣx$O0�)b]yq/٨¥�j�S��c�=	Pe����w|������86�kO�<m�����3<�¶�gW��ug��J
T.�K"�k-U$�a[|�U�7���]�A�ol9�kOP��5z�V��|}�ɤG�	�_>}�sn�'v⠧;Z��X����F`-ta�����m�h+��:plL�\^�Z�s0dI��>�qe���K��܊�B���\э�N�s�C������Ĥ����som��*��Bm��⛵����r�^����e-Bi��Rk���vb>oj�v�Lϻ��bM.0t��{bȰc%wu�Y�G�-�*������M�ۀ:�
8���E�1'��C���AJ���$��<��>ᯔr�O�O/^=뉺�o_N^M.�����:���}�rؾKӍ)'���>������{'Cu.�(��O&Ȼ+C�lU���a�i���l�{��!z��X;�瑃p�����U�DP�F@8�#�W�����Ud�ۆ�e>�{���뫨JN�P�A�t�T3�8��T"C�w���9�D�H���6��!J`�fS���6��G���f7\��,��8���`��n���Z֬�&8(�'���(rN7�c:�:��κ��aWH�TuӺ-ш��ѹ���~�Բ�1S��L�.bG&K�ƫ!��{�]��a5�D��+�_�u{�v��e�W�1#���s��cv����ڮ)��Mb1���7�t��'�l�F3�Wv(�<5kVa������j�t�W[�A�A�;�ӌM��ҙ�l��5�##{�-������Ν�d���8d��^�����zj���x�JD^S�,�	��,���t���jL�wa�9-��"k�4�W�n�y���$Sղwko`��0�ﹿ-��ի�K^�ݸY��^R�}�h��j�L۞:E��ڪi!�7�SKN�'کϩ�v�۞U�h���qՄی�i�X��h�Eqz��{S�܂��ԕ�o��(:'8���I�Dl���5ٶ�vk��KFK�Hȵʼ���۞}q�C�V	�;�%b�ܦ�q7X��B��ʄh�������.[�˕�K�S�#2rb�溧��r\�B��-Q�c�,�4wIF���L�V*�cUvM.�
�h!��Ru����sͦ�nk�~Sꄅ �Y�v�	����r�^Շ]ٶ���Ʈ��J�s��\ԧ��߻j�8�xT5�B�]rvfg��6�v��hk����=�t���`��NՎB��0��V!�5+B��Zg��b(.�P!�֘�Pi��T�I��r[��ΤnwV�:WVJ,)_ hʴ[��W;��j鸹7d�:�9��)�G�����!BY7j:w�Q�-����Oh꽱��[j��.q�v
�6���#^��}�;��>s��5�{�JnR�*J�ᔽ���a�xYu����y�Sҋ���ܛ`�������:���b�z-dNSs@w!�4E9�{�d��]y'�*����~�Σ�x^NM{z���qGaŔ=8�	�Yc2�Ӂr��7WcwJ�U^�v�gC�o��ob^V�ך���n׋���B_�e
8�g�j�W�l�m滴%F�&��(_S�XZY�+С�^F��,c��(/��������r�ë��YAu7�5ӡm��R�v:-�9`��3�W�{����!�70[]��V$U��5v"�i��ol���$�K%�P�4^�9�����h�7m�[L8�ZG=�*�r�U6+!XJ�(����L����5���!�����nۣ+҂���ZFE��F5;YH�%n�A<Ol*)Y�O^S�:��İ5�w1hQ�%�6�W�f����vMfr+{�x	�s��c좓�,��~�=W$���;���i�#{�|�Y�i��h��vv[�s�U�����]ӌwv��wר%�i�;�`�[��5v����r�+z!�ZW��0!��*ި��9����Y�������w⻨�7��qJS"�r�F�N�X0������as����b[�sy�K;���V){��kHR�F���aW�	�&�\��.����O���!�����]�8�������SBC2����:0��N7�Gb�p:�o�����-#*,ӜȬ3"����9yv��n�U
�<1D]�!롃 ��Mޭ�m�.�޹:����5��l�Sm����:�:�v�*�:��(g0�BF�d��Oq������w�o9�Kk%�1z��Ê�q0C��q��3U]�ݼ��&<[�l9�7�&B�Zu�vS�A���i���;�k9d��}j�R������\���P�(�Z�M����^�
��r[+�W����mPgc�������T/)�̥��p����]�S��eh�ƪ���v�׎98�J�o�f���{y��S]Z�=�]���.�G���^ؾ��ڄ����X)v��MܔllW��u�Fg�MwJtjv�nl],f��wG�ܲ01�꫅m�X��j���w@-a��sN�YJ�5u����<�t�_*��cz�&�f��wD՘M	�$]�VR��7�g8Nm@�Q�{{���,4V���i]�[��lw��N�NZ����[ԧ`���.�l�5h77��P=-,�t��qvն��y�r�u��<�W<G�{����6rK��a�3��Չ\��_;{�6���:ҫ�8����	�6M���kz�,P��~���.ڜ��,��Iߏ>���r�o�_���{q����`���}r�<��Ѣ�L�WS�z��򠖥O+d�׃�#t���W������w�6(tr4v�D�n;j��ct��n!�â���6�VqY�VD�~��M�ix�Tr��d�U����}��D#{16��Y�PUoWr��ʹM��7�P�Q�9���`�{���l�M�s��+b�Y��㬽A�Uy����������f{U�k/U��G�;�=N��u�����rD(�P��z���p�h�{����3�j�7oD����q��1��gM&M��Ա}xm��Qӫ�J�Ҿ���U����,�d^��#{s��NYqɭ���;Ӧ�����ė��-����u��)Λy��3���h�2Z3bw�WN�%.�n3a�eE'g�Z
��*3�д>�Ϙ��ǝp�I	L��@�b���v�RXݭ@[g5m��vgM�F��6�7/m=�	��]�&�Sde�)^mՎ�5X�!���P���ѷp���r���Ύ�ᔱ
h$���Tݷpj
�_neMQl7s��wr��*�;3���2��R����yL�c3��eV5�['<T.uq���I3X7 ��$����Ā����x�\�ڪ�q�[iɛ���԰�ˈ�{��d�z�v[�&�ө�/�h�ƙ�Ó����U��7�r���'��F�C�qQeU9;��L!���n9��]s���b+r�pa|����%�M���o #��{[�hLf��&�E���#3v��k\�X�dS�n�=��H�*��Ub������R��3���V�j��N�u��kո-Ӯ�4ʳ�"(CQFp��Κ\���R$�d�,q�I[�a׭Y/#;���������d��ݙ�4��G��@S}�`ݡLr��/�����(�γ��!�����j�����i���8��:��O3-�h�e�;�9v�`��@!j�wjC8,0 �#��-
�2��O!J�. �X��3�Q+
�k�)�o9m��0G���gi�n�K.�ɴs��t�8��g!���w�JJ�i�t�u��X�I��4��k�/x�����0z>u
��f���ɢ�ma�mV5@g9����͜˥f�_,e˂4!2�ҥE�2�#lТr��2ٗ��bg���m�+M֧�	W?���ß<4�I�J�lT���5K~.�����MQ�e�P��5�:ڊ�T��I��o��8=#0�U�;���/�]�k.��wL�<�L��(�Ֆk& [���#3�VCk$��׮�5��nU�)�@3��u�*�k���Z>;m�d�ܘ5)�ŕ��Q���LU��ۦ����:)��Fa���yp���S���+K0D��4��kD��D�W�V���T�튍�k(�6�]����`��`���k:���<�>w��Э�0�8���s*�N���.���N�n��1A]\�v���'FG%]���[�a�`S,ڒf؇zg�p�7"@�Q2���u�Dm*ۚ7���� ��zr|�P��j�(���z/iƩ!
�]4�Y�V-SYĠ�K>g*�!��*�܊�
�ܬ
�V��X���Mk񁵴m�h�mR�jUk[mUijնT+T���`�m��Qak(�V�H�J���X�B�5�-h�s
TY�YU�E+
[*Q!r�LA�+*�QjT��5�JYiH��V�JŨ��Zʐ��j�3,�[`�HV��T�QAeJ��Z��R�F��
�Q`�"eB��B9AUE�mR�R��J���
B���)�������RTe�h�DE��DPQERc(�Q��)5�QXT+�B[bȢ"ª)PmT"��\f9l
��[L�dƉ*�!(Ԣ�hV"
2�ȰEb�[h�[fZ�֫F,���P�X�PK*�JءQVP���%R��UF
�AF��U��j��`�����G�P(�ݽ����Y[�� .q��:�l�́ ^��]V�@��,��M�fEP�����v,�V�n�v����s{P!񝮧oof�U�S���sV����뼽�N�k��x]���z��Y��9���&&����15��Fǅ��N�}�HW�3����b���=��fe-����W���~C+M��yy�F^))�����3�ݓ{��vJ���I�W-��ȧ�WY��8�⬛k/2����A�i�[��YV���PN��lq<�ڟ��w�t.59I�b��s��>��ܢ5*̘x��N��,4�m��M�zh9ݢ�kd����uqf T���x�ͼ�גL(ܮ�o�]:��ە��^K�ؙ�E�*leD�/j�m�F՘�+��mW��OYT�R�5�T�F��;��L��n�۾g/�i]�#���(<�_1I�����X
��$��{�M�k2��{y�A��S�:�OV��A,�K��f�$���K��v�v�hi$=��7v�i+n�%v�k��r���;�vƄn����RV�бv�=��F֕V:�x�{6v�f;[f�#�V���c�dk}#�����f�� �C�� ٯ"(�ZQ�Y�Ԧ�S��-y�;FX�ɘŜ�2K��γ� ��Ʈ^��Ժ�5?׮�tˡ�P��cE�zs���ɔs�=:z�q���C�==��'sN�
��Fw{�5���lGZڮ��Z�w<�Y�1+�MbOB�o�<��+�4�*�9��TR�YN7I�%C���0y�W��P�kX)wJp�������T����o�5�۸�����2�!�g��L�|2�fZ{GU��7�ھ�s�˰W<2�G*A�z9���=�~�p��j��<�R��5��[�ᾮ��r��0Zz!���i�M��Rz��J�u��{
�֮��Eo��^��h�Lv��~\��	 p6����95�!��:��S.���_y���˷�(h�ݺ^���g���$3ڱ��畱4՝vcv�}u��
:��1V��[�t�V�85i�,�^��Z¾�N�xi��`>���<�_x7�;��o��5C�F욘�DH:3��#܍��M���1��;�޾�� [��9�$B�B��|�)�����L|�Y��AjZ�C��c��r�^c��e)B�C�8;���U*YG�y�����+E��Z�/�����$�2�gwq��/����˸�����W;<�d,]-�{];n�C��[p��3������a������܈Sף�*;ԟ9r�Tq\l,i�����X�v��z��U�[F�&��@u{! RFq�:!>��,p�޸��Y\��Mۖ�sΖ��Y�n:����}=i9IT����{�y����z��M�WO�oZ�:����ƃ �p���<��5a�+;o�k͝P�I�zf�:-�_�I�+������Bdw+B�3�k���]�2���WT�Ѯ�k�K;����Ӿ�޵�.$V�wE�<q�[�)���g�`��WT��:���>K�r�����YI+{$�hK]��uk��Oûʊ+��7�;�)����Cw-�OeUһٮ]���t�����pB�8����9������i/@�7��Z��/D����_\9u�_�J���*R	�-Y��8���8#�Y�jهE�V9�5�:�.L�^��_j�K��V��v��I�&���vp6�2�
�˔((qH3.m�� Tg��&$��/��iѩ�������0���8�wvV�יfl�V��� �8�
�K
�,�`�6z���YJno
���<�c����9C����˜��'����ޯg��.���1�{:�:�v�)��TJ�ǳ3��dM͜�M�)��ع������8�\�(}�7>�jּe�^�9�=�-���SQ}ni�X�R1�H�a��c��1�䙵��3}�ߑ���/�������w��z�%54�˨κq<�s�Y�(�T��-���6�y��gA�����u<��Yrb����f��wKX}`c��*��7O�ݠ�_Iu�$���-�O4�W�n��0�	�$���R��DX�����T���w-��+i0�+m�+wp7��q�����AȞAU���jv��H,Q϶zk1�#����ǥ6��v6Z�ՙm��^9���~�����2�����૽�B���ncubW!���v�m���r�8���U��;��-IvQ��D�j���P��Ae�y��vy� �l�1�58�eM�_ڲ��M�ﮓ{e':�`ma��Th��v`sܫUo�SC�wYu�YT����ފ�eb��u �V�c|�`�Չ���q�7ݫ(�!`A�*kgr�6t��5�}�ɔ/UP�RZ�<��[F�>�ܙ�R��SWoۻ���pخ�F��U���ڙO���nrj��	~P�w4�ar	��~w�iV��4�~]](�b05^�ب�r6�/���4�[��yT5�{��yP�8!&��*�����J+����		'v��jvn�kE$�8i�m=�	�musl:�I�C=�w�XN��=�S�9���!��bS��LZȑ����(rghN��1X�μؼ=���I�|���0btc��j��f[�bؑ�i��sɓ}{�TUE$)���8�����e��F�Tuى����0+�t��dZyY�8뤬,�᪦]:�}�ғ�7h�9vM ��f�γ]���}F�h���f"��4#!���s�6�g'��к�M;a��[a��K�1��]y7�~ u7��č�����w��;I_���5u抚)��̲��.�o�#�aA����2ᶦ����b�)��V��G�)�7�(B����9v*yo���s���<.o2�Ո�����=}]`�}�ǰ��ܦw�c�K"	��gp�j]|O+7��2�W��8Z��o�/{���7��u|��t��ܭ��w��c�g��Z=W��G-}=��xP����:ҠzS֩�_7��S�vNԎ���]^�Ieq�{=ToT ���]�t&�ǩj��ޤ��ț����w��]v���ƫTW����;t_L��{%��2-r���g�a����J�v�y�:���\�Rz�G8�qʚ�/wF�Oy��7o
�f�5e�7V���m�������J-��9�s�f0���۫k,�w}=��5?GeP\��ӗ�z�|��� �$%Ƴ����t�rQNnor�m�$6�)ϣV���.I>�U�-uy;���α"HJFmS�SS{mB��K��M�Ŝ�Q!b��ohU����j�Ĺ�X�;~�q�*����<�.�$����t�Y����B2�t�����v��ru�_�Fbr�T]�y�+^�ʝ+�u�lk\��8�[�z�uABA̻�V_$��u�y-#h�A���t|U�Ӧ���^�@��}P9�u�!�*�GpX&����!��s��ot#Q<B�3��s��\{.������t�Qw,���L��z��J�:�5�zkX�VY��9Z�8����-���T\�\%�q�\�7�o��)Wi�J�K�b{R�\������~�y���(�.cy���jÛY�^�oƪ�{~���j]����=K^����8�^d��OXW:I��o�H��lOU�t�X�^�3����ְqm�z�d�B�Ud,]-�9o��Y�t����k=��k]�JO}S�;�v�W��r��\�ޤ�@t��=��#.��/���Ӵ�^�.o��}s��zf�#��v!���bs{�f�f�Q��Nu���Ͷ��}�K9[ω�^Ԩe=t��M^�郕����/�<�����t�j���`z�6�%�5v�Fx�������X	OC��M�z��R�V�U۝�4�����To[v┶"���'�(؍�͹1,65L�wt�D�v��sn�@ӝ��1��[�9�}����1EӼ�Ϝ�ס�2��:U�R�핪Cu:L��w�((�n�ۊ��ަ�;���M�4
'U:|@�#os�%�����v���D����'�Nz������d��+\Υb�f5U|�,�n���6�m�_^�3z2��56�v�oW3�[�|+����7�8�djk�mV��&�T�M��c��9+����%_��O�Tq�-�bܬ�OhW�I>35��d�gG=�y3X�u�%/}�pB�8�\3�w�b]���MT������֤�ZK���Rg:��M��'ѡ	����(u��ec]y0��a�o�`�������:l훳��[�_dH�oo�rf�9ɯ5Y�q�5y*x	ޕ��-O��Fz��c]�яbF�h.c�8:�"Z���|ͳۃ���}]�Ыo�2m�v�.;��ɺ����(��tk:5W
F����w�vfx��k�a�yc^F�hR��Y�s�(F<B�ǎ��Д�7��������/iY�N�߸7����]+�~�?UXu��t��l�1������?[E�I��9'#_w]�tRaɰPe�K]	.��9J�Z����"q��x��hIi�:e��iu�taMv7�N=�&y�̘n5��[]�j�P�8���M��]\_$E�/CӚ��dw_�M��ד4��OGM��A*ui;p�3C{�Ox��q�.�B9v�������N�:Ԑ��2J��M犦ҝ��ݻ��7�k6���=����5BӬ��1����/eд��M�J������v��aie���n4^�:||ҏ�i\�S�eV�3~��"G�����-���v>�E=A��e��e�gN>�Ʋ�w�R�I{z5�g6-�,�.Uw_�\�YD���[�1�f��7�b���G#@���t�T�a��.'�\���D��Z���c�t���9�oW�ݐ�c�P����5 H�M���fGNົ�|��N+���׆�yj���n��j�ߺj� ��!˘qY���Sx�P��$%*G�W����;q|ys�s��b�kƤ^i=�s�{��e�NQΪ��`��ډ��x��L�'8����#c4��X)������ng0�������8
�h׻v���v*@0��n�'�1�S��\�j[=�v���M�'�K�˵L�]�,�]v��f��:��������ikF\L!}���KN�V੨�t{��>썼���EZ��\ԧ"���zU��p�����ȥ�\�Rgެ5=P��;f-�d�{�R�ĕr%��rk�Ր��1=G���W�]TO����<��#��l��L��}iD!0�\$rVi�d���k.!���8�=9I�]I��53���Rbg�;��oSN�Xe���\N��c����oj�1	f0��<�V�-[��(\�v�]M��ж�ߜ��n�f���[r{4���"W8��3��!�جIf�!6�δ����պ���Z����$[Ef1n��ۼ�7Qܱ��@��aȾbm##/S��QT�9�T�]� �҇c9ܫwS��p*ҩGL������.�9}��b����b5����%Zk/X�v>��u/=y^S�
�Ѣ��2Һ�N����A�Js_r��+7�[�OLv��q�c�,�4tr�{«͝����ؙ-ՂJ`���k��ՑM��>��<-�
��G�R�+.-ιG���K%.�X���e��J��dVo<��46}����psܫ8Pr�lw{׍Q�c�����2�kss���d1r-J��JwV���Yv�z�n�����I��(hYiʰ�$I[���1R�1�tR���̬ΰu�{�V5���ڝw�:��R#-�D�����=��;!r�h����;5�Ў|��Rٴ�V��*�΃���L��"�F.����8���F��gG�7&�R�7D�}�ٌ�qW4uS��k��=!����`bVhlɠ���s��mRu�����o =�����c�	�Y��Tdަ�Q��� ܮacW���ԷD;�e.�������/a�*�GU�ʱu0vJJ���CN�g�f�'V�TMv��� -g���x�e$�-�;�9�V�q���k��6��		��a��"Ż�L|�!7C5Y��}��mԨ�Ko��
E9�6$��w��j�B���8�(�	y:���%HWgfk��!Z"EW,�;�{0ԉ��G�l�EP:��]mŏ�^E'��<�E7ԃ�@qܛL�����V���/���;�Q�oX���u�,�p��4�y�𗹹j땾�M��̵��S��Qoq��&]��e[U�^7
�������\��Yy��m�^���o�y2��OQ��|�6W֬_��h|�l���v��Wc����q/�t>wT"�!�!wt���
v��1�+L;Qr��k(ee��z����W�ØڼR��X<{����o�=B����!Z�\xԖ��($:�N�P�ҥv+�>���ɩU���J),�)�F���_\usH�]b�|X�����f�]���G500a0���ff�gYX�P�h�T����	]2�5r�&^���,��LdF�4�e���+YhgȻwI�!�I�CT��Q֢���K����5v�� �=�*�q����baX�x92mX�1�3]݊����X���ծ�+�wJއ����hU �k<�]�QCE�h1x��]ӄ3nI���)eԽ*� ��D��͘����Z��F����Ŝ4�y��[r��K#@��3��|r��ʤ�.����2ѥ��i��m�~�@���
a���)� ����J��K�u;i<F�����:��1)�U����[]pXA���g��l̋��J�ɡ
ǥ�+GD�W��ܻCe�ة9w��c�G2UV����+
��F�ItZܺ��iM�j�7HHk�Om!dY+!�� m�y2
+hP�/,n�B k!�lQNj���/%E���[*��*J2���m��Q���P(�ʅkiE�YR�"&Zȉ�T�DE��FXڵ
�*���e�
�Z����
J�1@���r�qF0DY���PX��W��(����,-�*%B��JШ"-J����b�m�E�9���F�E�DUH[X�*�3,��$����(XV(�`���"��b����
���*�Z֢�A@X�"�ER�S.ZX-�T��*��(˗�-��[b�*���%q�T�1�((����ł��"*���)m��Ь.fL�9X��lkE�Z"�DaR�Ԣ+�A-�iQEAk*�*�4rʉE(�e�A�TU�IYU�S(��b��Ab(�����e+P������*��([q*��"��QQ+[j�kDb��(ƶT����PZ�EP�!	yP�D
�o�7���QS�8\j3d�\K���[��x��z{y��k�.���鶢���r-�-�wغY���c�3{9��6w&���ڶd^��\n��Y�7a^��7ʃ�v1��B�xWFO�o0���o�U|$<u��5h��%��<��~������_�&���kB	����ϗ��6�K^1T���Q�	�u^X�o-�}y�� �
1��S<���3��tU�3�s���2���nt��R��u;Ϝk���Ը�n�cyV�f��;�p�X:�5�zk`e�<�)L��؛�w�4�r�q}�1ɛ�ӓA*�w��u�1<v��T����y�|�諌��2�v���T�(�a��3yٯ>�{׳V�5���{�����,i�����'g��8�/2�d<�(P��|�l>�����n��u��g9���������=�Cd�����:�����k������V7yj���|�ٷ;�e��f�;�ug����'����Ò�͒��-7˔
�g���%��<���m��^J��B���#}7{/��X��}��q��J�|+�N���bz��=|�'L��wC;nF���k�W9q��1�������yd�dn�Mnj.��]Fu�ֵj��w_Eg3�r�=�#}$X�{Xat����YS	0u@BKw.觼w��[�x"y
	O!m;�z��N��k^[�"��T�m/9z���rGrÉ�Z/�P@�y=�b�	��]�.�Z,Zn�V�y�����n�tq�c�T�8��)�Q�4���u.E�War�v�o�$����F�t�X};P@�bZ�F�Dzg��Tm�|�Ū�j��}���ʖwKu�-�\�z���!�9]��{\]tbj�:��gK=�Y�q���j�~��!��ί�I���vn��*jm6�D��?)�EP8������T\��TsDk�_N͊��at�-�Z.�#�o��sBZ�n,B�&�b�v�Q3����NvU���}.de[�^�M2������1��x��:��(u�\ʩ�s]mN6֊�~�mX�>wy)�����93�s���=='_�WM+�.�-��V��6�J��-ZQR�I�2Ƥֵ/0�eIH�6�+�\a�*�x�3���yҏ��O��$U�Wk���1iM	�z�M��x ��X�ۼ��[8�5ݔ$�I�1�5LY��N���ƞ�W9.-�}��|U�;��*b��Y����ܩ0��s�r�y�pl���3�h��w[�D��\�Ov�p�(�y�+�����\���5�/1�8������$r��`��Rb�ԭ�}:kC5m����pF+�j�2�E�gq��)S��S�s�<�gS��b��k��%*1��p�qt+�9I��X]^��Ը@H_:��]��0O4��b˰����&��=5�;�o0D�S���BN���mC��Ɵ�M�� w���9sM��/wp7�x�h�)j��cEzp�O7����ӕ�}�]�񈧧ZzSxU:m�--�T����5I_x�b4��Y6�)�빹�񃕤f�Tz�,����ro~˭�Tuc���w�z9�Y-Cg����=]�2����R�|�I���<�-��9�}�e���ّ�ʊa)Fw)���-+j������x,��4�z?q�l�ޘN?u��9N�nu�8lP��F�ɝ���b�z��a������{�%�i�
���b�E�P����G<�Ӟ5�����e#�ssm�<�0�=�On�9w����D�)�n���+ǽ�(���0�wwab$GB��N��>��gs�u�I�iv1�H�EP3�=x�wٓ��T.Z�
I�N}	��Yݭ� �\�OP��k��� �h��.��kV�+Et9���F�-=�dk��)�}n��;�,��*�2�u��U�sNcZ7���ѧ��z'(�+�`�����m��HW&v�w������Ի�r�qP�وL�O��&Ӭ�x�����c���`�;��a~Sm�����%��&=�zh5Yʣ���/�����[-nۜ�6�j�5s�&�+�9p���&���ɠ��&�Vu�X�סς��T��x��;��=�zy�R¯=����N�o���V��4�W�n�<d�E+���=���P�8�t')��k����y�t�N;1y�͘��* mʚ�h�z�-�=,t�vr8'��k��iW��Oq�t��Rr�LۡB]�@�N=��X�s729���:��w׫g�j�j��O+,��!�Cge���c��YҺ�/�<��������t4z�T���,��=�]>��W4^fu���r�*�w#��V��N�ؕ6t1�G9[�S���z6��Kh��7o\���3Շ��}핝9�����N�5��w�j�o�<�T(�k|�h��"PJ�)#Ɯ9�0s[�,+����S�c��|<��ϫԱ�����:9P��閖�W�r�u�Ҵ�λ����SƓ����޿b��y�b�G#n17N�!wlr��k����e�sEϵL�[K;��c��;х�K�v���a�i�����ڍ@c2v��r�F��N�]�s���:r{���m�vke��ۑ�kOUC*��d�*��`���q��GCw}�p��jbnq���{Q��'8*7'��g�3zE�@`ȵ�|���bi�VB��޽�E�褯�����^�vzOW��Jθ�:���,��DK6b	��=<�[>O۽yz�����}8�a��z�ۡ} ^ُ��/�,b���B{$�	8�͹�R��;��W���cq�{Ix(j9P�\��һ"��K(,�ٻ�z��1�a�Ÿ�q<s��p*����꺕����r�kWu[�#s{D��kS[�p��^���v�h���Bv��D��о�X��Ņ;��Q��k�vM#�Q�D����9:8v�=�٧7�pE'n�)�Fuק���!�{5��>k��؝W{b���c�R����^m��;�^i�PnS8��\�[���g'"�'l��7��i��\Ʈ�ב�o�X����y	���z{�^�h(�)�ʔ��+m%\k37�觼ol9�[���'��A�Uq#��}r�{�����>=+V��m ���Ll�K�Frc��u����["(�L��Z�"�u歧��;:��i�N��8��U�.l���ܓ�KrOc���kEOO������S�m&�]����Z���w+�[���*��*v�rg2��ts��E��jg�1U|�,��j3��)�pm�%�9�o_�5�"��c�3��Bgq]S����3l!�{���]֯����@����fWJ�'�/#�؉ǉ��8���5Y�#i:�|��n��� kj�w۴�d�{Z,w	�{�I�������a��̇�H����0E�v�hu8%#il鎺d��H�s����8�<ذ;���Y�Gw�nVN�V�R���{�^?.�G��Љ��0��><.�����(^N"��W4%�v����*��y�+��S�)=0F<P����ʗ��Z̢�펉M�w��l臠������!�t��me�R�ȋ�bk9ƍ�^J{��L��&�������훎�ՊL��'ˮNc1;G�ƤNb��c�{�����'ܙ:N� �
��@�9Gw�9�zԴ고�P7c��WBqڼ�7i�a^_I�R�ۄ�<�ݴ���3�v��d���&��^q�����{W{f�DbtD���v��fy{;�m׎� �e�kz�M�Շ�@(ݣW�"S2Z�n��٭�b�s�d5^z��r�Sj��^��zz��֞9T��Qs��A��Ċ1��K�u���ZCc�
[m�--�
�D�t���� ٽÞ֮�~��e�*��L���!4y 鋬�T"���>�]������t�!�+C;q[u�k�A�n�����(�b�z�Y��X�%��C�8�����ͨ����Z�J��o^��6��!O�-�\(��u�u��޽�@�7{��<7�A�=BPS}.�#6��Թ`=��7��4#b���������+��U��­Q^S��kE�	a*�놫)
���� �/J���V��U��>�>����V�R&ZWS�/Uw�Fw(�t_3�ɶq�粹�T�3���5����z�Q
���tr#i`���!�V��[�Oղw��T����2wRE�=����4���5�1��#��<�N^����0Й`Kn�S�!���}��'j楧A�ؕo>=�>���fkI���8Nfԇ��dz��:�ozm<VЗ)�q��Fs3x�ͬ�K^U�l앥���&sL�'���-dN;{}�^�V.LV��˯�kF����CT>?\��ד*��������/:[��Ge®���N�2��h]j�CS���:��{g`Md5p3��&�!��bα(>:���>�IZ��:W
Ww���Ȫ���Fg�����ƾ�a<��Y�ta�v��]M��oR�{���.�[��5����:@�k2='ld-dJ#��s�#�2M�ʂ���|'M=wXԗ�ޛO;/PQ��O��4��^���jλ��ck���K���HsJ�֊�~^����t��J������R���P��sY;�D<��=�fr��&=y�{���ֹ��NSoU{�ivCyn^���ܭ�VK��F�'�v�4`���'���׫پ1tj���)��B|-q��*=)����pÕ�X�Ρ���k��C^������s��$ZGS\�:0&��)n͸u-ޞ�-o�l�}�h{ލW�T(�|突�}@D���s��^#GyU���+wq�cx���r��x���}X��u�)*F�1����<2(^]�٪��(�-b�H���.�Y{.�M��.R�F�*PYhw�Y�*����Ē\�6J��W�3�\�����5�Agt��4��rY꺍҇u�5����c�Eh{�m��=��F��M.���� ��LU/L��E�e�i��a3#�{/[{�lu��9,������y��o�r��G��ǆ���q�F됬��:��-8!嫸��Q�Ю,��W\CUс��n�:�r%ڬK�T����}���L���[�	��c��EcD����Z��6i��{�"��G�$<T0e�q��fm��R�b��0�$噫�!��������#�)�%��j�w�R�������8�ba���Xuf�o2�O�������x��+:�@�{�\����
��<|Zȼ��^�˧ӓMVC�z��c�H�Dtl�4�jᲔ+�8Љμ�7(9|��FB�ɠ��&�w�����i?A�x���Ͼ��/y#�FC��(�|��GF��8>ӓ�Cz�d�ݛ�3���x����j
��u6˓��ٳ�6�{�y)3�{��-׵y(=�IN��N5�z˰@x��,"y٥9��U[��Uwm�����9��q�^5�B% ] ���s瞒:2��]�.]�~;o�+�.��.�
��rGn����������{� I?؁$ I?�H@�XB����$����$�xB����$��H@����$��	!I��IN@�$���$��$ I?�	!I��IO�H@�hB����$����$���$���e5��e:�e� ?�s2}p$����!@$�����T�AIR
% ���J$"��QPJHR�HU@������D�P���PT"H)AIU��$�@�mH��DJER�U*R!PBP�RREP �P���*�JH�D��PH-�� W}��(���*U$�R� �B��5 ��RU))AU�DQD��iP�Q��%;`��"UJ+Z�$B�   ��aN�jD�m�5�I��.�ۮ�4j�+N��e4������ݗ[u�3�.�0Q�*�T���k�ڴ�]�A�N�NR�T)J���   k�mVգ�N��eWb�ѱ6�cR
�r�5mJm;�ws]�MS ��lV��;�L蕃R�)V��lu��v꺺ݕAA5$�BIHJ"�H�Qx   ��uC�ݵ8k�k�Yĳ[]wm��kj�f�J�ڶڳ���ph�5�UZ��ui+[t7qΥr��B� ��C�.�B�HP�B���
 � HP��UP$��  �   �B�
(P�Gp�@(\;8�
$P�hm���8�A@P�B�s�r�Zڰf�;�W��YA��ڕ�9\��Z���WN��8�-0]��ۮr%)AE@�Ux  ��@
�Rj������ѣB�h `� 6 +D�P���#UP*Pk
$�Y�ڪ���j��I
��)Q%���� �� �-�:J�l���4�UJ�+m6��C�Ψ΃��`�PcD�)�T�U@�T5�B�T�c�J�  a���h[a#AV0ѧS]����-SJ��7N�K���;��jS 
�L� 5��*��8U$��£c���  cr�(��[�ZmQ���U�h�6�u�T�fq��ݸ�]إ�n����vڭ�ӻR�CT˳k��f)���s�ݺ���$�)J�D "�<  l��SC*����AU���� i�
L�n۲�4���gmҖ��6����R��K+)�[m�ہN�ݚ�d�kv�@�VT�N�ض���R�)$(%!^   �sM�Ԧ���Z���ٓV�XZekC*�¶�mQЬj�hkJ�S4a���v�wd���wmt:����:�:�*�Y��o 5= ʒ� 2 S�0���   �O�ңG��  S�A)J�� z�Ҫ� ɑ�M$D�T��♌�3���͂o'���bii
]LL	��)r݃�zfi@+$q��L<��I������$ I<��BC� IO�$ I?�	!H�B! �.2������T�Z�S))��1eXw=y��O R�h�{�Y��]D3J+�)а�s@�
V����&��BW톍ޖ*�M�opD�IFݣ�VB�96��42��4Tϖ�Q��[#�Ie-�P��V�'`a"��"�Ի�q�DZ�R}��@�X}e�۩�D+cl]bp,yy�׭a�0��-B��*�`��D�-R56�v���k�eܠ�b��ej�˻���DS-"��LJ�N��Z�]:�����dY��[�%6v���B�ڙD�ܵ�Y2+)R'���\wI[4.�Ņdb�&:�Ժٯ�A�O]kb��!=ҍ]	�6\����tl{Q�`��i���%�[�&J"�j�DW��-���%\�QB�4 �@�u1�&��.ƨ0S2�*�U�6wKs��lt�Fr$�ģQx���
d�z%��u�7) EYd�t���ي�8I�IY{�Ϊ����b���$�Mڪ�h�����/���v���T�!-���K{����M8�n��#v�	VX������&�����
G"��G��hnzP��Hi�`#r��RcH*��Tv�Rݬ�8�#w�[��v'��Q�/`Nl�h3yVP��N wXT����m1�J����L"ū�YL�$����Y�����bP,S�M*��,�`e⹍��&b0�y�BQѲi�LP�4JYwH�-�4tEσ�zȌ�B��2�g؆�Cp� �2�"l���&��(�)z�D��^�L�L�R����@b����d�Y�HS)e�� �h4Z�eVAz�=8�nA�l�X���D���^�s+E��%a(�or�ui��Eѫ(�p�d��l*mR��r=zN)�q�1Yb�"�e��r1L=[H�h�R�/�G5'(0���l��XNc�jc��g�-;����ɭ�팤Emt�1�z@ Y{��%�S3�%��28M1ZL�A�^8�b����j[�+.$ܙ-ܠ�bQ���"��t:E+.j̡LCa��)�V�HCY5��ʏR�t���6D�Xj�K�J�+GEe���Ua)�cJ&��IȎAȨ���8j�ʱL�ٲQJ�Yx�qE�ecê2n���	Q�-�o&<qm��C�P�Ia��/�c )Uӡzڧ@*�Y�Y֛{j�VYp]���^�+5H��R��}`T�e���鴷>IkpP�jKYngZ�d�*�I��z�Cq�4�6�E8t#WP�W�ɫvbcl'(n� ݭ+];��2��cV�.� �iZq&�
�|/	i�-e܋o.J�7XiM��Y�����c@���Z���5ḇn�5�a�Z�m�ԨH�j�76&6)��w+C����R�lcF�[:��]ڹ�	!?�^�Pf�32S��LbSZ�NEA�YyuF���5���1�Z6">w�q`vR�v^1��v����o.W7l��k�ҙx���{46V�7Ci��j�q����f��*����D�95ސ�]��Z��C8��������BU�f�6�"�-��B��ݑ�)7I��f�=O-G,�867
oF��1h@i�-5�]�c)個̀ƴ�4��	XYM�Vj��b����]<{��`'=��N�!X�0&<�jS�!z�)��&�S��B��Y¾2�g۵!��H�vF�DR�[�- `H1�����&�%ۀ�����iIn`��2��ML�	9���,@�5A�b3z��Cw~n�~C
e�{S��A^��m��0t���F���X��B�5�e#��%m�ҽ�q^�M�G���J���J�ݸ��N��(�ud"U�u�i�w���6z�����&�c`��l���4u<��j^N��e�l����5TY�,JST� �ͺd� �GlɷC�ĮS�ȓ�{�0��׶e*��e�c
 e^��[CXچ$�f�ʗ,�v�MJ/u�%Љ@Szv�m�ΈX��	� �D�6��*��k
ˉ�����	�e�`9b�B&\�AЬ,˰�ti��;t.��X`���c�%+4[j+�G.�ѪҒ���>�
�����e(/m�YX%c5kZ1���^137D���ߤ��j�ި(L`\� ���uv�%F�Z>r���,h��4�Xi���]�r�:#1&�"<"�7f�(�e^��1'Y������[V�e��j\���FI��o(��]��Y������+�5gU͹�c��@B<y��Y�j�(Q�L(�*��l`�G��P�{�n��oC��������.�|�"q�A�
ڲ�@��I��N��l�mMI�I�N�D�_*�f1Yt7&��-�b�!�/U��hfb�Z��ɛ�j�@I4���i��ũ�إm��]��)*&�]��P��d�3u�Ǚk6�[��6�b�f؉2<a]V}s\,<��ci�&���hD�t#��o3Sl�ף3���hH�Ŏ��zVnԺ;@�r��5���%*U{��B��!R������m����U�J��e��L&ʗ�q�QT�׭hGsS˄�ܚ�A�R�"�&�l��m�Ҥh��H5uMt ��(Qq�����y��뫢&)M��b3�0m�[b��kbS-�~�9𒊫Վ���ב,!2n��Lc�	0�ʬ�T"�k·L��,k��+p[�l2R���7V�O7p!��r[m�� ��`�ˡ��tbB�-�����K/{��XF��2��
lXT4`y�n1Kw�J�Щ��v�:A�FV���Cf�t(�$�n��uk�6�B�*�+6��2�t�fLs$�bZ�I�K~���[���Ȼ�u���ua
X��N�'Z��N�Lt�Vp���+p�i-էq�X+"f�l|��Č۳:��x���oh�4a����Y���@�0Ep�6�k�XqV( ��BF�e9!̹���c�V�q��< ޘ��vF�ߎ~jn�,�f�9����N���4�P_4Bܵ�)�Fʎ�4��a�S�GZ�V���a��/[ee$*U�VPW��Z��JSқ#yW�c*۩-^�qݧrn�b��e8�	�"�6�A >�:�FG���pR������e]A�b�&ڹ�]ёгi�iV���۬nD0*(^,nb��Y�����L 6�F�ی�^-�U�o%=О���R���us4j�Q6��dk&������7�v`V&ˠv<���0D�Rb�Α�V̎�U��ۥCe\
Q�h��ކ])C@9)����՚�L�v�y�*+�3��\L�S�!�.��}8�`@����ӻm]'��iLyqU������	hͅ���(�q�[�YPٻ�T�y�K���5�(�ăiD�	7n�U�(к
,�%h���a�z��!Z�������z�+V���Yec+[�X�	+`�Mҥ��ķ*l��b�x��YG�7�����;f3�0"�y���P&�rV������o^�74�`��z�c���+�V�^	kҴ䡀�{����m�SP����*RYyR���R�:��.ҭ/NaMw[��i�L-9�q+la��%�&�U�u���e��b'O�6b�Ζ�H_чZ!̋kA0f���D*1i*�Q�Z�L��ݙ�У�P ���X�օk6�L��{�V$)rQ�(GYkql����N�%Gm�SY-G&E�JQ�}���9[N�j�h�osec����QR��;��zޖ.)YIQL�!6k�l!�4nZ5`R{�t=��&��r�Ӆ���tT��kZ�.���k �4����ZV��Ʒ��K���*@4�-�-d�
�h�@j�H)��;4<x��jZ���dS�g2�\�N1W�4AR�A�s�W[X�d�X*�44c^�9���j��u.�A�ܭ��]�!S1���L�)�ss6-dmz����{p�/�cY�wl݅��b��ۂ=?@��l�() 'J�,��V[ `8E�[j��4�"�*�O��8VY�����17v>Ȫ� ��Ӵ��wA���\ȫ�vI	^f���Z�������zCݫ���?K7�k i��[6�r�0㊝LSF�aD�,Mn��t~�ah�n���G7ա����",P5��@�L/hefV��3L���{H������d	CvΪt�p��u�"*�`ٶ�9�;� �L�HD=ɴ��(uSn�Н�GSf$��j5\ܼ�lJ(���B<W���CC����D�G�PDul��ẳV�dVB� ^b��v5��ّ���=�Ϭ��D/y�㩣n��-���m�	���SJ���+�CkS�˽Z�eA���vдC��`��4��SVm�.�oTGe�I�Q�Uj;$h�W0֦c̳y���D��j�8�78�1�ڇt�w��.�7h�{o�	J}�n�k��a5�F��2�&���a�^Y� ő����B��%dL�����&�֥�l�h<����f��ki��$�j�)P��n����m�Tub�jP�P7���Y��3Z�A���Xu��SF�p���Ѳ�_������Ì�nfj�� )���Q���Z6ԄcV�JQ��4J�*��Yf��i�n䩡����$�x�(��t+z�SS*�������M,�sr���w4ҳc6�J"���i�_d�a �]3n��*����^ֵ!Vl�e`p�Iy���d� 0غB���V��y[�V��H(�ڛ�I$r�kӟ-JՉe(�`��^7mc�׫L5a,CE�Vd�N2���h �*�ݒ���U��,�f�B!M��N6�߂zW�����f�#7+�V��0LO#v�Kf�����4-H���h݋Q���U�l2�JɄ˲������0�Y�Y�Z+&C����Y+B4�D�vsܬƥ�A��Kbe�E(q]�Je�U�9a����F�����RY��f�(���Ż{Q軨�L}�XqK��]1��n�<%v��X��YC*չ�fm%+3u�σ�D(�JC񔭡�V�1��#��wZe�ѳ����t��!�����ݨ(n���ּ�����]=��E�Ia'IJ�v��hL�@���p�CWm��脲KB�U��m≐Z��ti�7(���ةE�/T!�Y������i��ݓHE�cp�M<�c+��t,�7\��n����ٖvۘ,Ő�ci%������2;m:6��%A�C�n���V��&-rem�ܘF�dHӔF!eÉ�1�;0��{�6��F�H�үu5W��Zgm଺�d�Щn����+S�b���.F٥.��5����L���hc�%KI0%�]`˥�툷!&QP�il9K[�#��]��m�m���6��p���<�#d:�]�`��@3L,H�f�)�q��Q��-�,
[q3F�/[N�����(70K#(�KtO����"�]$O
b��Cl�J��*a���#��I���Ed횼V�*�1���6����wM�lG]��AST���u��9Bm֝6-�֣�������ρW"w����]B�B���Mӕ�J+w1��ǪU�ԥ�w�4��WLȐ�H�櫚oT�a�17X�x�
q駘�e��yu��&��%ӕ�����{�hX捈5�
gj^��Y	�}d�ڊ�&�k�5T�J��*��kS�qɎ�eBW[�@U�#�x���V�
ZH��/t�8wF�Mm�V��e�"@��j�*̚" ,�/M� [�J�x�`ǘ������wlkl�M5�
FVkTN&+7!��MP�3�4T*���юVi#`�/RũN�Xqӻ�*)��q�x���H��$r���г0���f*�,MԞ��ƶVI�n�s�	LV`D%C5�ق�5�Dv����ޡ%[u��m\
\	D9e�l�7z�%l̤$Bn��G*�

x��:�I6K��J\����	ƛ��,��S��^}
�]�H̢m��-�o ����ݭ�m3cV�i�d��8)�e���ێ^�/F�����X�Y��˚f��`Ф�����s)p�6,ݘ.էokT��t�\��Ƨ$Nʖ���*�oeZ�kȟ<�3��i@�}+ĝ�Mv�$,b�e(��ZB���w2K�4(��B#Y6
.$]-��r�X2*u��kU�c@��n��M��<�2$�*�^��(��%�fּ�X/t�P���G�0++Z�q���Z��{��9`%�0=��ALTkr[�P�f�ǌ�tV�ubS�֜�s��Va�����X���0�3`�j�%W��*-�z��i��\��B�l��kNVS��7�N��f�:�F��2�q^��
��vvY\*���N�B#�\ȭ3uX��1��� U�,��qͥ��T&�
�6F��I�[%G0l e��o7T;�\D�u�m�:7@Y��
�kq��[܆+D�Ս|l@�`&�X*
����xd,h�+2V��ϭ�[�Xv,ذ��C���r���m�H���cEm�z��i�Gi��ʛ����7w X��\�oR�4��w�pfk
˒إZ�8ݑ��B��okcU�+M�B�Vv��&(�Ĳ��pÉSYy2[95X1�F]K;i�#53��9 m������r�٘2�]�Z�70[�)��=�gv��5����ax�ӄ=��Y.I[Z's2��gv�Ā�ْS��:l2���eX�	�u��f�n�^P�2�l�Y�B��t'�b�W{����k�`��Qj#��n��os,��t�
�.��dҫʓM����6M̥�s
z�`��/���;��Xۅ��X�.%ʹ;�5�ͤ�{7@ɛ[�[|(�E�(���"!��M�
��F�A���{z�L^��a�A�CrZǽs(r}�r�9H��W�H��R۩I�!��	:�;:������Z�0�/s��B��dy0��놅ܴ4����Q�)>4�l"�<�8D����3���R��w�����2�l4�+���0���Y�n� ���k��f�Q�ˢ���Uc�=��a6�����Z��ۂ:�Y[�|��^�,w:�NoGYy�o)�V��3�¬x���������Z/k�j- "=�Q�:�36�Z�
���*������|y�U�(3�6!\^�VF*Pk�]Ϩ�/u���Md���=�W�mo�Y�%L�|�݆7C��GOf��o��SSM�!AA�l�\�V̫CU�$�rW�Zx�߆K.�m��k�ͼI
6<�ضyB���YQ`k0s�Q�h5r�hҶ��j`Hdd`ͻEx:��U�O{��x<6���]��vv�E����2����^��u}��E4b�جJfb4:�`�V"#�`�#R]c��G#��Rޘc��;Oi�8䭺�V��7ٽ�co軓���m,��9�]��	P�bΝ���bz��h={�J	u(�k��R׽F�[�8�-,F������\\�*���w@j������XgI}����7)?��A.���n���D�����i�%˴��8+���0�s�4��6��rs;�2b��s�xI���z��'������q�����������X	Ԙ����4�|�L�|OeQ�$�����KD�lX�\\�nW'uίli8��B�Jeʗ�l ��L�Vu��]��҈YD��c����$Ġ�M��>:3��";GY������m���[�Z�S�u6������d5�bZ�_|���R�^>﷚5��K�ͅӸΑk�y��o�奚r�\W`,��� #�;�NI78�r�ɸ������s����V�TU(ד����}�
DnB���������r��RVj�W�
Ku7to*�V*��o�E48��72�Cw�<v�xl�� �H($g/Ts�Ib,gՁ����\M�u.��u�a�#Bc�B�lvE�u���Kr�K)v�'�P�Ȝ�
њ4�.UB�[��R����wU��V%ڡ|��ר$�� ��\��:,Vr[�roC,8�P㗫���څ�ϥ���	�]L��^��q�7}��Yw6Y������Ցt0QL:y�AЛǠ�2����̸˦Wl��u�-�>�u&N��sw|��T�lѾ��Ѣz-�W�]Dʳ��uz�vmkĊSr�`[��!�wK��B�j��a�r��ɡ�VQ��geX����]H��;$��U�T�OZ�o�f�[�2��j�^�����[�MG�=��0�$���p\�3�sl<�R�Ȗ����Gy�q�l��/�ֺ��2��yY+�m��3��6���j�:S$mUƺ<7J���m⚫�-3o6Ne2h倥�!�6�\`ɻY�C<��PP��wE]gs�j�W,�ҳz�^-�ح��J�����/�@���MC�Kʼ����C�R'}�u1���m�ڏ�o9�G%��O1\��ҷ�n���k�8˥���Vge^Ӻ��.�a�n�諟ן@�8�:2����睛îuv׌c�{���햹��Ы;��N��;���/'�ܕ3f�S������B�'*G�u�o���V��n'6�V˧��+�(����a��& ���]L�t�oP���cN��Oc����e>Y��lބ�	��GIe�a��ʉw\��s����{�7���o�V`!��P�H�n��mm���}��N�Iv�0��i5r�e��AGf��ɤ�+��r�1ud���]��p����E�4����U�����n���J�l{�c��IG�V�P���4��m��M�{n�:j=�	�"�t��%��WB��<��n�O,��ê�R.�GE[crqK<�X5[۝��r�70!M�Od��rfػMf+��}�,�jp۝[W<���|��ws�:�t���`)zc\m��A^���ʾ��͗XӺ�Y]u�-��.M�8�cX���Q
�'�klbk�]t��1��o:ѡo3(]�s,5t�<�u�0ؾ��%���]�-�2q�]j����؁��a�\��cZ�ٕ֩�/b����n��sH%R`q?%��	v�s�_t�<�ܼ����V�o&ˋy��Vl6��.m���B��F�[R��P�
� n��J1D��2���vJW�e)���qG1r!w^T%~>[��x��iK�q�y�oVT@�l�t+ ���jg!��iUd���ty�tE]hgL����X
��ف���4�rPRl��1j,�� �)B�_P2�7B�pZ��}��m�h��d��u+��
�{j�x)�}�A�v�}�]�x�N���\5O^Vk���l�l��ڸVa"v����t�xn��uh��*5�E�R���T&�p�ޱJ�5JG]j�e�m;�9l�wlPK��]\sv�{A�"���V#����.�	Q��i��V���M��G����s8��S��܆��Vv��k*d��8����gye^ҏBJ
��|^ۦٸ�s�WW}���H)��Jx/�9V���5������%��9-�hGY��c鵭e�LV��,>��=XB��鈗�;;vō��Is!�Wou��o:PG%�N�i�Y�_QZ���_L�z�=��-gq��(m>�#�\U�����n��7
K�܎r��զ�N���}h�H�<�z�Yڳ&�}�h�jl�V��a� f�/K�N����i�J����xR8*���ZT���Yw>�^�۴��0�V�������Hs��Y�d�}������+�������ڂ��u�N��胾β*����t�;oo���(Hڎ������� /V5���v���iAo4<�I3��j�}˔�]�R�y���gN����X�%�4�'yXX>倜�t3����ɾTٵ������j��'�B�r?E^�:1Ӆ����=.]<�J�1�S������X���﹆��[c�
�ݥz�3[k�ڴ�+�Y��shR�T�#�\Y�jː��Ù�.#�8��b*�B��l'���g^|&M�*��9Hq��[<v�k�}>�e_h��+nЈď(�D;f��&A����W��nv;Afc�Hu#�Y��mLff(�n���}]��y��$,;�DWJ�i��N�U�ǔ���U��ކP,�q!;�.�Tf:��j�r�D�r��sՐ`��lE�\Y.;���.�c;�
��ˮg~�^5Oo�r�S���^Nm�c&qe��t7�:�`eN�"r�@T��Q�����3oCX/��9����֗7*�qA�-��'��2ݝr�m*#�i�V3���Jۣ��\>˪y�_Kt	�6)d��B�����n�����/	����� 2�,I��԰m���7xf�.%�.���d �>�J���]v⻈ń>Z��EY���B���ĩǏ@-�iۧ=�_Lɱ�d���F�HK����n�(�d��Ra�߀�]��w#�2�<ޗd���!��hh�����w�WZ��+���
�z�G��n�/�"��4�7j
Ƴ��U�&ɾk�Z]��	�S���s�\�iAP�;�εwc�V½peZ�����XZe�s��FU��j�4tlю��ᇩ�ƭ@�~{kss0U�F�����-Mo:뭸�U�Uj�B;֢�2��CGq}B��m����ƶgG܍r�F�#�^��q�t�=i�V��4���R晲��[�!9
��K&<ǯ�f�Iu�zd��i��#��3m1��3�^BV1M����\H���ՑbՉ��t�~V^l�xul�9��K��G���kr�B�ܟY��K�B�y��n��D�*V�t&JUN�̷ܳS�9��+b���v<Mn�v2�K(>�٘W<Q��6-N+�d�����u�[��q⢼,�M^
�|��WW5� ����G�b"�p62u�(X�k�-����}BCY��q�W��f������)�(��)�5�Hb��͒����/U�)�OJ9���M�"˾��q�p�@KT�F����\�fͼ�k�[4.�6�}ST�;�_fXs���'M�ϻ2��s�;;��f���Z�³#��\�Eչ�n4)¢�&ۻ��c�j�D��%ht�CQ�T�����˒�Ή�/�o^���淌�������*V�xjV���g"+6�p���#~����+\��\��Pv��]�-���%Ec"���#�ݝ����^�f�hџ��^�1et̍�+��ff(Տ3q<�zv�N)-��LM�F�d�����=4�I�v�~���dͥ���^ ����q۶��9� q]�q2,N��ǃ��:�j��	u�s���l�w��I�ܼ��9$�j]^�+5R�+#Y��2�U��k;����v��L���˓Ju`�[�� X;�Ғ���غE���v�"�b�*ܥj�#j�8$�µ����Q���~]}AI,Wn�� a�W�P����\��*<F-��B8�����fPT*QK�+uf��H���Z�d�R�33Z���
o�ȥe�؂�4.����P�"�n+b��Fj��_�Ε=��ykO�٣�����ڴۺÓ���]_�"��V������u���J΃pSYǦ$�,���,]G]�Y	�$tT++��6�����G�A�h�a^��%�<�u��t�
�6�_�b���v�w.��-|�g(��Y�Q�M6m4�{[K�j��jƳs����r����0�b����"D�]���Cn����v�(��Y�f�X��������])rra�����(��cEͥ�]b�[��ʜ�57
��}��k�w*n�a)W�6X�3���Ϧ1�Z��3�vwj&�o-�N����-ʾ�B&��T5��wT��r��v�偔���'`[ۡ���[s���b�5d�ٳ9��#�-Ե��b��ev((jG�f�;V�Yqq���[uҐM��N�y��O�!X�����"�=yI�s��ǇfJ<�nMYy��m�]v2���|,���Ũ�����K�%,l#��2�5ڴ�-�,�0��Yܢt$�XB�I���Aa�c���l���TkI��\�36�vҠ�����*d�"-!j��SGzm^9�	��3O
�}���N�'t��:���鵼2���7%�),˵Ս'wv8:�|jf��H۬\�����#gki�Xe�����2�rqSn������?gs�65z��B��Yc�&8�'>ѭ�h��P�Բ�}i�k]�lD��r�j�\�z��%�E��"�ڰ�L�5���	.�K呞(�x��5�ku��1�)2J�C%�{Zw�FI� Dԁm�)Y�.�Z���y���s9S"D�F��7)ʴ/�]��z���Ѯ�p�0h6�iג���h�lk1�e�8��.�LXܾ���A�v>ъ�#���>C}L��m�D�*�qWZ�p	q��w
-���^��#~t�8h}�Ým.w�;U�F�c1�[��vIab�|�&�O(gJ�����Rۘ��R��^j����9�]Y�Hv�T�o��j�ҵ���f�i�0���v'5R�Xf���֩���oX�Wq`�l�ݬk���;a��NJ�1�S��}���
4S�[[A��;�j���,�9l@	�8uL�k���%k�hݎ\/1������Avn��SLC�3n�ig\\P�HU�\g,�5a�7(�lǜ�(���{9�:"˩wR��9�o��	Z
t�}�{/1$��81�c7Ri�ۥh
}���z���6t{\��36�G���z6�T'm�I�]�_m�*�����l�"�H�#��c�4���bJ�R{��vՓ�}��r;wE�Agc��bm��7��hmBg�k@� *b���tk�>�8�)�< �-E��.�l�Y����S̩��՛Pn�x�5)���D�.�0+짚{��%��}��d�8Q��R5�Q�/�\����j˘�1�jTz�h�={�<	���vv�Pz�W*&J�u�[�O��h�.^�wy��I�4vǷ�"]uw|;RSR9&_:2���,�=ֆy�m�MW ��\�B��"�&V!+Tݹ��b�#d�-�r�^�:�:����ޅg{l�*�KNes��2y\�;k*u)�=�V����*�.�ҭ�sE2|U@b���tn��>
vP��	}2_r�dN$�fG�+KM[]u��Xo[˛�١{D����ZMk�L��ش�t���ǫ>�m#(]*r���Z�fВw�^g�8;���:�Y�%.�xU�qK(��B�!Ɨ�}ymm[j1��$��,��Ɩ#;�l=eF�n�U�ֳ4�:�d���3K�p�����(�MK��Z��
�����L�A�ݹ#孍����c�yG���X��b|�nv����bb�lI�`筡mM�c
o86�P�Y��U������z�����!�ʝa�����{�1]����4JI<W`����R�ǚ���#s$w������R�����%]��E�$�jR=��*V��Bθ���O�&���T�\�7�e�o���}�7,��\)ɴ�}5�[X�bt;kt%s�_v�G;�ڝ�����6W]L��SZhĉ*�4�s�������;�T�gV+C.�Eë�H^��uu>���y=�:�/�
m�=ޫZ�}���W�~걄ʾ���&��/I�SM)�Z�&��:g����� ���$��=�������\��Օ�`;��i��77�
�����GX�� ��e]tyܕK��崫���O:=r����(�;ëV=��ǌ�[	��oz��W0Q��N��h|(so0j]W�%���Xьإ�G�b;�s*\U7��BV�٭�9���r�up�}Q���,�]�yڰ�&���'NA����KQ-�,n�������yg!���YX�I���B�Q"�bV�^���M?��]O��c|֊��z�nf�o��MX͔�La`s��L�-�|���3F=���9p;bmsb�����M���ҩ��L�%_2U��Ӆ��G���"�B��OEe��]��'`�>�.�]3`�r��hk�l6��E 9㊻�]���.źgb=�8��������H�}�،?�㻀�3@�Ksr+�ݬ=�1���d�hd�@t[K+���=����6�ݹ$ql�q��
ܜ�N��R�Zj�f�|\���V�;Qx�l���:�d��u/�	�*H��Ed����9����DZY�+�pvm�)־]�^�J��9��9wR��J�,��1b_c�Wմ\YyJj���7(���NV�%"6���O7Y(���b�v�m)�v	.��0�9��.�r�]ج���t�3�ojW����K��#v�PX̬'m���a�R�n�V]m]l�+Z! ��9��L�u�7O
�5��w�:�n�KP6�h�$&C)���*u�r%�q�Kcd�a��/�ToA!\V�LwN������������V�t�E�C6x��(�{JO���̳4gp��CXa�����)G��)e��� ��+�K�&���h8FI����p� [�v�H�yD�.��z��)һU�9�U��ܶ��X'�
Ø-�J��͒�R4�Y`�7x�ڈl�7���s�,��VC�z���Hc<�.�
��~���,�$����s7d������t[�� �6�빸��f������2WXU���O�z5�k��%��;sgO�
U�n�5y���u�Q��`��)-����]�R/F��,�*���5�:���e^+ƹ���n�Ҽ>���BZ���Ĕ���ۘ.��7E�MQ;ʬ�m���JŻ6�p��İl�[�n&��2H��X
QM�6�1����XJ��˕�!��F�Ug�l���؍uD�����]�K�"�xf7V+�e"�au��v���f��yu��ۮ��	��q�)r��vV��㗧D�f�o	��Ch,Uoz�ek���wX�Qjpܷ�r����Y��a55�����mLy类Td�W�l;m�J��.�Q�;n���hj�%6�.0�_C7�LY�=Ǔ)��@5Z�a-�]][�ǿr���2e�o���+��A3�334��L��FfHq��V��F5�A���Q�;�3��89�D�(�����v;߰�$��Eel�k)���T����c�I��U�sn.�������Y�K�T؁��bv��K#�bU�[u�VV3RQs��fg)�,�\��3�}D�7u��v8|�Ug�z5$�N�S5˧���{ـ`m�ou5���B��`�����o1Ǌ�i	ޢ��ٹ���+LR��c���Cz�խ^%T����e�*�#�p���Xv�u��
��W�	\�[[�����Ka��9��c�ٷ+��H�_A��q���6j�-X	"R]GU]���kpf��`;�U�o� ��pJ������P2��
��މX�nY�n��6���������]��!ă B�3�9������]-�`U�����an��	����N�+(M;:ܭ����ˊ�T���پ}�R=�B�2�wE"%��#[�X�~;j�Xc�ڋi�[KfrS��Jஷ�k���FH��)_j�P��^�/��|U#��n-��нU�V��k��Q��&w��,�u�+�G�k7).l��k�y�B������"*\ʻ�7��3(��A��� ���5����ܤ�v�ۙ�ˮ��n�Թ�Y��//1�� s���X+{<�3�\�S�3�]��B�j#�]�ű��T��1�K˃
�E,[Zŝ1WU����I-��lk�s�i�TfTdz�m�
P���LmI���XH�S7NL�����T���U����L����zmÈ�e�n]2��̤T2��X�sV�+�[6�&�*��1T��n�N��Y@�q�z�e�����	qt���z��T�����8o��[��ݵ� �eL%n��t��7z�)���
�u�P��*h���QV;z��\C릲�hҬ@��]�Y�Z�M�����0���IR�ҡ,���us�H��o{y�^
�onˑx�2�{vJ��jK���ɒ�b���'�fsO̊a2�;��ͪ81�TO�u�W�#�U�.fCI w6ݎ��������P��G3�MwV&�^ޫN���,j���ۮж��ra��C�;�@VL�*7|qAsm:=�{Ekǀe⒅�����(�6�ZV�$���O�.-�Qn���	7x��<��]ԟ[X��X���"�nTGr�v1���R�$�������w�;���+Klc��n��m:P�}n�=�0�PeC�;��B�u^����x�,Ԓ�PP�ydJ�� �y]7j�2����[Xh��3 ���
�wݗ���6ݜN�T�w�mݡwX��(-R�9�*�+4Y��Z.��/I��p��"�Ta��3SiԒ���wR"K[�5t�z��pGB���z�,�1:����1C��G�SFmn�}��g;��
���#�W�5^wk��"+�%@L��F�F�����t�"U��gSC �0�mm '�އ�>��}�E��vRw��딶� ��e$l>{@^��J��ޣ��wF\�]��.ɤ�&W7����f�7�����ui�������VGLR���&����Yz���v�u��%y��ґ9�u㧳-EIvر[�y�:6���G<7N��/F��52�����2�w<���:�>�R�X4�_e���U��:��*�5�nu�݊�\Z�}N7�0�\ߚ5��/�1����Z�{����x�bJqVǊ�6q[kV���d�j��`&�d�G�ti:�\�5��ed��ܥ���#9�=Wt�j@�TՁ.���^��B�V��P��k����(��(�)\V�"ڕ���[��Y���,l���j�܏�b�.��O����9��}���quƴQ��&p��9V�Y����w�ϧV�R}�vD��\р@��/^�i!�	m��a�R�ۂ2Mι6%Lj�ެ��A}�ٵK)p��a�i�G�5�-i���+^v�oY����8-^sYS׮�"��i	�h�7��CY�l:y�(*���r�S��K�OU�Z��7[��K������j�,|��[|�tЧ��N��]RV�>NWs!��}պm3�� 1�X�|�-�a�Ȥ^����%"��]J�X�q�q����|�û\�ѕep�,et*��E �C:у"��jj��Wd�\.�i���k�
t�꛶�&��J���u|k�c�QSB ��U��
�S�k?oE��S�s��J�*� �l�̇P������).��=��l���ݏ%�U/���b�2˗���9e\��!�B���+�(D3uIu��t�un0�VV#�%�k� ��4Za����ջ:�R�RO����z�\�Z�2[�ȗN��N�����|�`y�fIGu�O�ӷ�V�z�A�5�'/��]7��K(;���	����6/�����Y�V�Ұk4�ý�[�-(B-�t��)W覐��ҁl�dU�'����ћx��f�LqYj^oNw۶����t[��#��J��n΁����phZE�[���L�m�S$��H�/�w�:w�nT�C����L���&o���j�����w�sW:4�ݮ�{&����r����4dρ��(I@Nꂮ����av�]��\Y;�+	B_}�#��J��������ֻN�.�Ups).��_J\u���T�ʶU޺W�+1b�����_.5�Պ �1�W'�n�#�R�*N�kU+�R9JY"��2���]o[C �թ�q�U�+��/�Q�[2S��|�3Y�X����*C���A%:���#*Y7%�s酉�/u�Cl��뾫�'wN��0�9t�ʃ�,���3�cS ���;�Yis(D�I*�Z�5�w�xN/4�O�l!"�����j�SBJ����׌\ʕ.�8��i��Ȇ3!�&���c|0������B�9o"�)ܵu�C��Bg��#�:+�H��s�rٵ��g`����Î�}w.޸�ލ�r(+5�1)�Fl5�(��q�x��Z����Ve��ˣ��ӀYd��!�M��e����v�!�ue����:��3d�IN�}S]=umF���:�Q���=ޜHB����μm5��G��kI�>޺x����tݭy�~��������8ta�b��p�-u����U�
�������>�\���ͬ��dZ�����3$�J�����Y+cp/x�y�%ٸ6�9:WJ�V�ˊ
"��P��
D��wX��2ŀ8��嚇TfWNZ��S��/"���϶ȸ�����J,S�GCYnѠ�KH8��p�	���0��c"����
h�l���ڜ�bV�e-�]�j��jgg����j���=��z��y8�o\�6k�F��-��'��U�L6qNn���$��b����sj�	/�c��Gz��Ac0���,���e\�N�����F��gr�m�+�;Y��2 �������W+1m"�6���{]b�\�40o|�q寐�vH���1b��N(�<�%�\�)���Ey
���u$�7p��ٗ���Yc
#�����r�([�c���}�I�;�v��;ݹ�g'��:���Q
�(Í�r���"��%�nV�y��䣖��Ciܠ� �nҹNZ�Pe��[#;)�t�X��*�Ni�ikq�C:�G�\V~���.�c��:�1U��s���zCY��h�gС��2㳆�ڼ�er�[M٣Je�� �a[��R�$A�L|z�L��R�6�fرM�K,�r�sA�}�b6�LL[�������FٻRn%�˂��h��Ȼ��3��WΌ�twIy)�@�8K�VŅ�f��v�;�yT��A�rQ�����*%qھ����a���j�rk�z�t�z��U[b)���S���cR�N�#�mۭJ��NBa�hh=���+.��T�Fb��o��՟7K�ap���*`	oj�w�J���+�7w�u%(���g�e"���������u��Yw����]��7)Xq�LR�<X���+]�m�Z�;S�1�%sz]�R�,�����j�S��p�Yu��7��M�n� $�}�^j��y͡q���P���g+E�7��ܫ�f*e]�Ȇ�x�|��m��� Hzۀ��g:��V�, ,`/��f.��R�9���l<�x�6����-^�V���]�����呂�]��<B�M=`��!I����������u�y��be�����%�;�ݕvY|3��s�e�]|�fNoN^�uqR�	۫�m&��j�sB1l�ѣ�Nڭ&M��Rx��:��5��z�������ݡJ�6T�2�vk|�c�Yϣc��)X�&��|U^-�)gK�ۣ�m��j�II�Q��
 gD�'�H
f��`L�$� C��Β)Gq�7 ���
�ū�G��Aym����3f�[�	bn��ܠ��
v$˟^�ꡌr�-CU�(r��*��]��9B�j����MdO)ӻtg:״�����G@P�r���zj�AOA��[m�fAq}���X����u�����gY�]#Ƃ�m�Q�e���+mM�zֺ{WƖ��DQ�(��rT���߯�M1�;�/{����f��A,���V=E�9_ƳF�e�%ˁ�Vr٣):ݼR���`Ц�k&�B8��a*n{��*�.�GU�!-�:�E*U���̅Λ��1�0�Af�;8�u҈��]=�+���Fh큍��.�9�Yv��٠��v}�ZW[BQa���ai7�1�ü�ү���¬
�,�R<�%4�J����]��LDU���2}�f.�*`ކ�;�jL�%���>����Vp�r���,��]��(M�S��}�.��F��(X�r�QQu.e��V�!���}�iU�=t���-ٰyr�
��(%1��ũ56�-˫EVh�2�a��n��
5y�J�W1�,�) �/8�0+���i>�p��B@,��n�ѳ4ݚu{��z�:�� �։f�ݭ���C6R��+��8�ya�[F�q������!�l>R���ׂ��}Y�*�@���ww��Y����F��d���>ۍ����x78@��ah�r���e�9Z�����x=�E�f�2����`�-ˎ��oh�f�KQ����L��CnvtO�kZ��4���N���D^U�(_gU�±�ϫ{F�νwG+&r�\N�2��\����V��K
����w���b� �ط��-�1YV�݅͡�������,8f�:Yʌ�E��QO�����_g+&���xp�ukR�>ǎ�e���E�S�L����{D+��N�T{l�&w8�c6�ϓ��4nܬ�s
r� �6"��]��v���]�ڗS''�G-�;�Ԧ�|Q<N�U9)ٸ+3|K-\g������9:-!�xwZ;P���e�/�}U���� 3�b8@���0L���و�%nT�c_�40:�U��a��Y���sw#
�Sn�8�|՜�c��W��������[�Y[�m��$��t"�ʵu�0���9���e�e��1q�z���fHm�0K|h:���w�I]}el��`�ؘ˖�����Wk�C��(�ټ�6>������к��/�5BA��kL6O7�Ƚ���e�Еii�5�����q��+4�9}�6uõ# ��I�s'u�i�AVd��o ����hPg����tZ��ǥ<�{Yy����.�He�R8z��҅Ǘ���Yޟ���i�v�F,C�z'r�{�#��r�:i8F֭�U�
W�=���h�=��á�+�ŷڻ��Õe�Va�u��1ږ��\�_�r��ۧ�]CG��2�݀�i1N�ڼQ�z@���4�:���yn*�"5�����h
C7��ɓM�I��L���Jq��q��!x�]�Z�5�.Ӊ�I�pm�h]�N@J@| y��M&���e��:���MZkO$�J�Ջj�j�L�3䷺��2���(�4*{�N�Ǘ��	+w+����j��脹Oc��Gp�k5�x���J��w}�=#���w�Y@Z�]u66k��h���b#����N<ޗ�}���0��p��υttЛ�r�T-��3)�K��ki��N^�W�<g*���ۻO:Sl"C)N�o⻷�PJ
�c!B�*u�e�g���*{I���B�_�w�E�d�k��I�pK��y�+�2��q��
<�;9s��h*�=Υ�;�Ot��Y{0wk�
���Źj(���V-K��M�$� ��+Z�h�1F�!F��DKjffDQ�**�Z���KD[`��b�aRեB�-�1DF"҅��TX4e���mb"�[JQ+k�DeJ��F1�"�+j���X���j��Z�֨�T�X�Y-�*7�Q2�UF�,aZ�D*��T-
�iU��aZ�Ԫ �k�,���"*DX�����(��E�F��[c�������T�[J0Q-��6��lA�B�KQ�-��TDAB�UE�T���UV�cD\�,EDX�m��T�X6��QXVQV��R"�"����Eb4J ��$TX�j
)m#-�l��!l����60QĢ#F�m�QQ+(�%�Fԥ���Ub��(�."28�(�*�RPVڶ���X�+Z�D��F��#V�[%b�ET���@��jX(R�+m
��#[m�*�$X�����0i[ER�TU��jU��T*Ŋ��m+�q+klF�ր��"���Pkj""**�����~�?,9ں�T�����v�ʼ�pF�N�NR����c����P��pV�����;�v�������h�Y1n�7ӧh-sp����-q[�W��;=K���g[X�7�f�u�`l�r���Y6��;�[���k�kkZu.����D]mH�[k�X�(�tlث��?h�>v�es��5�PG^�!��2�ܸqal�B3��bZ����!��ui~˴����krU�K;6Xȣ�!�����p�h�ǟ%�|6�0��)�
fɋѩ��|��I֎����6w��|Wb��X�a��>�b�g�)������XUt���eM���:���V�:��W=Y�m�lJ��0$q&�G(V2B26@�5\F!�C"�n��";a�̰����"�c�n캧�ݙ.�]�\4.�2��S )��z�
Q��r�],M��ޭ�����t�v�Ey��Q~�$�U�qb��@�����]��zzA�؆��W%����8���.�Q}@ٵ�N<��A=+h~�ك���
3���k,�4p��y���y=��$��8c���+����s���U��/<��R���> v�U宽)*����\wD2+�Y���W�\*�N���b�*l�A��\9r�q�����d߀�����(�sV>�w�v4ݭ{��tf
��_��:!���b����#�+��)�]� J�*&.[�+�����r%_f%˳5+Et WMT0y׶8�{���3rK%��c�͒X��?lAAթ&�����A�=Ou�\ta�������g�)���Vb���Jx�_O�{z0R�v����]w�|�����[ઇW�Δv��#N2.�� Fx�M�9o�b.�(1�MYꓫ�Z.(���6}��~H��v騽�n��91U_�H�Hx�_.�ɞirԦ4� ς�p��$Q�z�U�8}>�a ������'/U���[��;x�� ��}�
�����k|=�\3���eGE��"���&�5����絮��O�6��̐��~�$H���c�O�t9���<r��t�afn��˵�	�Nxִ�M��b��M�"�~dU	���Ď1s,�ޟ�!��R�q�;�vgw��͸mL�Q5u-L�[\`:]o��zrb��b�	�B�^��Ȓ�n�b
���HB2M�}A���&�/Ӎzzknh�uw��y���@�������8Zԇs��]��f�;�`��}�D�\i^�@t���FszS�*���"�:����Z�ή�2n��٦�Zרq��s�^���[
�0�)wJ��<QY�m��nT/��U�W�
�n��}`�(>��F��\�~G�~�M��9��gK�[��7�j���JQc�4ۃQ�ڰ���&��$� �+}�h��t�$dovT��[V�1�(=^�=oH����d'a��lc�r����W��m����9;ڑw�Rv����6���xs��ǹ�c0�#__�������R���R��&���2����L�r�ݾP�^Ā��Qm�O�x�Bą���ylҍ�,�ȑdΙ��[!�wrҜ���U�$��2��0����l���o���lp�f*�^����a:�l�(��L���Ug��UǥFp�j&�ȳ��^jAjDD3�"��̫���ƾ�<\���o&Y��f�./Ǌi���G(S�H�9����[��ߜ��ݵ�"JB��?#7�زW�Ua�[+q�5>�o���yAQ�D�� �7肪YS�Vƛ�nQ]x�<����K��7b�
UY�����e�F���quS��ma���y�'vfۥ�yF_�,��B��{t�ot����I��ud��:���R1�nx����(�l���c	G�K�["j�]29#���n����ʋ��}7���_zE�׺��u�E����uPc��d]?^s9 ���+�w�Tj���=c7�M��<�T��]�,M:U�r��{4��L�Oz�jt�� ��G;�ˇySu�5�K�o����|�o��1n�wf�g�U{(���W�'a@��.����K].��u5%z�s�6�����6�*:-l����e�>���./�G�U�9�ɀ��v��=~�ۻ��݄�0�C�魡�9���z���j�rX�4���>��6I{��w��C�5y[v�V�8Z���`��:l��#��_�J#��h+9u;��L5湁�q�+i����T8o��'�}y��p�z��R�8�/��l��ܲ�Â�����T⊏b以�*���\��C!׭�]3�-�Y�nx�͇`���}T(>�����U�q�f�����m��C�*������ѱ�d�� +��dP.�p�k'��W5�n�_�����h���x��(�Ol3`�o�	��!^	����9�J.#����)���~���~�$�>s�2�� .��_����'n'FO�f�-�^]��j�u���^�e��Eϱkǰ.�	s��.��K����;P�G����:W��ۤ+�y��g5coz�ԋ�֔;�_�d�x�V=}״-c��->=�5֝;�oR���1wX�N4≊+?<&�=^�ȿR�����:�ͥ|���m�\�e�_A�m���+�qAg��$�
s&L�5T}�:.3ssZ���ʋ�'�l�z?gv����'�D8���a�����h9� �ز�9�'U�����|ڜ��ϳ�[#/�wJc'�k��_I�#��V���r�tE���q���'��x&X�JeJ�,M���'(Ӊ!��!�HD:,��]�qq9�p(o:�n����Xk�cђ��m{���4� �ܙ����q�vT��!n�P@Ϸ'�,�MK�Bj��fu,�.��c\�<�����A��40��Gkj��#\h�7��{	�#v�)nbQm�u�yٖO}~S��Ytz�&L6�~s8p�#=�x���vÄ'N.ѫ6_3�oG1�%Є[���'���4pZj_��r��5���[��wW��ƇL7�'���UK�fy@�WO}�>�z�\e8������j�����>:I�xVd�ӷ���
$��^�ҩc�hүk�9�\3��
�q=�K;�%�����{�fK7-	�xڈ�g��)�j�8�7 ����n�2��ӕ\�w���<=f<�Q��*X�5��n�[ƫu`4�"*oY�����l��Togu�Wf��� ���ӿ��
�a��S�R��t]��Q���'*f���fv�ӄ��۩G�=��%���԰Q��+������1I��'M��VW�v�<�ƢSys5���[�����6�l�P��v�:���m-�_��!ʑ|�)L��z�Q^��Q��U#�}���	�������Y-�:��6ۺ��%Ƕu�}��A>[�^������l������5���F��ʸ��J%E�4��8Ⱥ�4 �Ĕ�\�s1�v���$��>Pm>�;�R�-��:�[T8�߹S�g!ϱ���4���s �V�&r `��<���Y�k*$apꃱ�h	ӗw�F�t�@���8I�,�)�����h=���Oj��g��A~���W�vظ����*�G����'�m�`��lsbݻ�W���{�=�!?�hGL����1`�>y炥&�X�07v[�ݘ��.�rC�v�,��.��L�Y�1���u$Q㑙B�瘊�{C���Rm\�=�"��уw�&�m(�q��Ug����y`"�]3Ҝ�+*�(Mٿ�Ѳ�*й�(�Y7)wJ��(�Z�6�{k-�(���C;�A��"���DY���X����W���YX�`"-�z��hj�Ic7��\T��S��<�7 �WΛ+�������q�䒋��DN�<k�L��݆��L�pN\@5:��C�z���m���ü�a.��9��**��I3oX���9�.��ͽu��8��Toyȧv������]�[B�6*g\ag������ڧѮE>̖���:�Μ37O���Pp��Vb�8>5:	Sh�a���V�ixo�m�@����\q5�W���q�UfrTVF�YY����ٚѹ��3��@J �4fDt���̐΁���4ڋ��}9��9I�������]���
9�QA@%* �d�s>�u<_�XЉ���I���5�����+ey�m��0�97毬0�D�f	] �<��+"jڐ����kqK�(�����́�'kO\�N:�u�(��'"�H��Uˀ�b;�r���g���v��ʴ�ڡ�
Z<�Pv�G��{c0�61����v�we4f�`vQ8�܏Vcx��`3&m��(z��H
]�(Kk��^�rP��g��(�B�_pU��f� ��v*���;��eߝ�2j�����C�
�Q���.��ŝ���U��m�X��'{N��f	��U㪑>�n����+�{Z,x"M^�V��{5�	'v�vƕc��ze �mӦ�4p�EBΎ�������E`�le%�Ѭ�f8���:7vb���J��&܋�*����xwV.�,ͱ���A|����be���0u]Z�b��N��E��҅���o�ݘ��y�l�O>��n8X#���Y(8���Ɖ�ܜ5}�
�Oi�	��e����Y�򴸉��ʠ�ڥ�U:��̑-=ܗ�� �brg&�H����y�z�T��R#��d_��҉�4}Ç��������e^�@Z��z��7by_giy�i]mL !O��U�Y�"L�I/�h>����Fy��ݘ&�=E�N)+k��̭;�qX)���ۣ�4��ƣ\�e_���Эu���ģ9�S�����ԗ��P�U/6&3Vp�܂3_�nO�����k���JW2l�3<}^��X�2�����4��N��RxtZ��8�Cȱ�{cy�I*�
�J�AV:p�28�;���&Oa���a�ɋ �8�U�é��9��zݒ.`)n���ʘiʢ9��(�Ӊث}���s�Ku�6*}�͜!�����{P����-W��+�j�׊J�ڛ��>��佷�Wg;6DmE� C�2M�p0T"tL�a{��sǖk�v'�TQ������N=�t�NG�[(�p���7\"��ɴ]h�f��u��K3%��[IY��u^�:�[��^�Д����u��n����V8�+���:�f�;}������˂��3�V���[j��}�p͇��H�ƅ3I�Nb5f��;Pus-^�S���(T}�U8�����;�6dS4�f��6�Cq���a�Mˋx !
q���c��ʇn�K/n�|v�O��=2d���	%��|AZ�w��,
�맾��7I�|n6�[�y�eƘ�;lmt�$�D������VP��+q�A^n�p���V�Q6��$���]ү6��{ڕV��p#�3d�m�p�&`�˙��9�=�&���3;�;�a�K�	��=�ѫ5���8��ӗ��$-��Yȡ.x,�&S�s=!�^;Pڥtv��ږУ����Ɱ.\���{Ύŵ4r�9`סOdno�qr7&r~QON��꿝�$��5O�\NHy�p��uT��T�j/6��>ɵ��-�;}�:2��e��D���HwMW�s0(`�9W�@ex��7�|K���-�|f#Ӫl�$������A�S0y�tN�P��:�]E B�{(p-t~�7#�)��$�ۻ�1-p��|�uせs�HiT�,��F�j��+<D��.3�ko�p����|(��-��rd3nïv� ��)��lv�Dq�3����!g�,�jގ���KD�t����[�)���׍�tS�N޿�zx�V�r��H��;��n�y9�^��O�0Ƥ�os��ǚ�D��Y���d�E��:N��{\6
E���Y��A'cb�ސ0�;r��Ҫ�������k�����֫���ts��h�rB��#�,r��A��>�}�[��{Ұ
wL� =3 =bv�A� �*���.�C��3�z��fo4��k��读��Cz�S�e ܂f3���*C.܅�T��5E<�r[nz��s{�t�o!�����"B{N����(�@��;$Ϣ��H=�ꂲN֑Ҕ���M�L�97YcvGW��E�����v�[�h��E���>Ā��G�w� �oS��c�/uZ�W�l���t�ч��6\E���hsnwa� �q%t[��k�*`���]:9)Y�Q*�5�(:�$\�{N!Z�P͈s�s�d�w`��mE���5��\z�v\����hF̶׮�Y�'���{�ؐhÜ�Y'D����7#k�f���5����5��w}��������O�R�*�X�"Z<���];�2/�T�W�/%������ޮH��g�SDJw���y�ʕ*%*s��#�HF����A�vV_f��(�;.�
��[�t������QL�3�
���GHf_����{�YM�����K�n����B��
��3x�����\F:7Ǵ��>�F��2])7���ĭ����9�ி��c'u��@@Ʈ��t���ar��9����:�t��<��!���J��$M<`uwu��{�[Nڡ�>c���.�YX����h�F��`\U.�v$*ռs0�Kǫ�keizԷͷ�}ۥb�r�,�P����;N��cU݌��X�VN-p�6�6ի��"[�mJ�5vY�(q:�j�g��	��֒�xM�C��V�u{FKѧ����߼�+�^�*�O�L>�2�wV��{V*]%����0��Z�r�zVZ�OM���pB�3�#�b�C���Um�� �&���F�)P0�m��R�b�q4��ˑ^Z"=&�Xv4ۮ��L�����1x�5);�Ȏ|6�Ew������^����ƨ̸�ތm'��9��m	*�c/Ub,��ݘ:�b�s�'��pˬeέחZX�ѼT�mC P�5�(��4M���՛��w��f��������;���]�qgC�f�f�����C��A�fV�K6s���:_]ll��_�ԧ���K^b�ky��o%�Q7����x�����M��D���������Y�DJ��[�Y+�P��%��2�K��Ë�%
�4m�=vn:=�*�21�0ρj��y$�^;���
5hPla�0=N�O1i: Z)���M^m�7C4��b1%�`�X��cU����p��pw+f]L���V��c
�Y��X���z�K�v��,��j�QXR��o3 T,������j�1xVY�	<[����3�o+V��H�ov�ز��7@z^)^�Ab��rJ�aЎ�a�+��!53�UpeԠ�������R���/A����*V�N��OK��ՇK)`jعbD��*7/��smͻx#�&�l��q��D.Qe�4�-+w�ð��HQ�ׯ&�w�.R5� m�6�<ғ���Wr�nGD�.�
®�9�Ê����FA,�,R�;����`I�+^T� ӻ$�"������v�[�]����� �N
ИHA�f���̥Jk�aV�u���T�l��ے��<Ӻ+A��Y��IIf*`®��)SA�"�VѢ�����֝ە{�u�*��wFm�A���.^;�f�h8��.���ڗ1D�����|�S���y�b�����D���cZ�4��[--���S��%U�Ԣ�V��bQ��"(��VTlYTb���%����Ie�Q�#-�1F�$`�Ъ6�Ҫ� �b(��(�����(�2�ʕ��֢�`�Q�b#���J""**
���"5���EF4JV�J�j�Q��*�%Z(��TQD�`�1T-���D`��(���+�EX�h��EUX�&Z�S)jPX�X�UEAjc1EX�(�1H��V"�[[X�ŌF"*�#e��aTU`�cR�bETT�2�h��TZ�Q���l���2��b*��U ����TXŊ��,U2�UYj�G)Uph�U��E�1cb��Rڀ����P��QPQDE)Q������-�EUU���LKQb�e��Q�ѤTTLL�R�UR���I���AKE���X#l*(�
���X�\�6��F�kQAb��Uh�1QDTB�J��������*-��m�5+�*kB�+"��X�TUH�>��Q��G�T2
��ۙO`���2��/�˶8#'N�;f>�4^��m`��bl\舯%'p�PficR�:[O��o��#�k��v:��g��?�l|Y�_U`���y���X8J�,Q��8x�~���؍mj��~3��4�>�f�3�<a����pg���A�v��,�|	W�9�q>Q��E��ʥ�뼝�yB_�ͮYxG�#h9���sq����DZnfs�3wV�>���:nm+gV����`��VZ&���9�� �W]E�䟪�ܬ�O�������]1	l��!n�1R�q�g�zkb��<�� v��n��6bQ�[��|+\�g!k7���n�xݟ9Qi�9�R*�'ˉh\�<�k��p�-�.�F({S���>��~�s��Wn�(�"�6�"�T��,��Kޝ�Đ�b��B!f���<�w�#C���-�Q���]�����Q�
A�$�>��B����V�����*˺�A�c*�Q`S�"��x�w���iɸj�״z� ����;E�i����HH���,:y�� ld��!����QC���cSJ`o�bԈz�m�T[�Y���jP���#L�n�|��[�o[�c	<��a�-^d�=�p�xQ�]Dڼ�#�]V��Q�޶���r�웤���f\B�2�N�����;I��6�}+b���%���k�e���7;�ف �h�Me;l��R�m�UWYz��3��4�1r��	ېoE��݊��-B�8\Cb ^��x�+׵z|��Q��#�p�@汸����(寘�3Э��}�kB7Q>Z����,uל�N���c]2B��E��'kHLl�^>��<+�t0��5�����������9�$�j�}���M�I
�ʼuT�����
j��[����EXK��*r��?,3b��~C���Q��(�}!�Xl4r� ��Nh>��l�{��5��,�����R�2g?{he2�&�@��Av̨f^\�d�m��v�����������9�Uhxo�dv�W�V�g�zk�8���{=�Ç��y׆�8�Z(j�&�`e�� �꩗�FJ�1p��%�)�#<p�3p:iУ���u������o$<�ä́Oi��Dz�WL@K�{�n[��!z`*���`dp"r8�����8T���b1�uE�`uK#��J$�:<�j6Ғ�ɲ����Lk�� ����)���8�ږ��nq�9wV�y�%���V����&��v,�ki�<���Wl��:]��À^ ��ޢpc $3�ݘS�͜������8\u�/�u!���w�+�5�Vs��%�^U)�䫄��BZ���yV��V�U�J%Q�R ���q������if��g.����B��
Μ�پ��)fomS�Sq'�LwGO��f��S;�>gv-�d%�v+EL�W9H��o9RH\޿M�]�l(�\�PY �����u� ^���K�=T�NY���;:��F�҆E�)�o�j܍���/�e(l�&n�%��[�ZB�E���'��j��5��4���}w�X��P��j��F��GB��q�	%�т!t
:�݀���'^z�Q��4�,�#�#�y����\矬�)�8}�#Ƕ�C9�܌�@g&槪��}C!fHU��Q��,�%�t�]9��>f/&J1E��I˭�s���FsW��+��8G�zIz]Fܭ�J4:Ij�d)�q�|��>|��Vˁ3��|��bU�c��p�l�U���ӭ�1���z9`�±W.�J%wvGS�WDT���\U'Y���QnE�v�)uT�Al�1�+��B7`�z'&�J��A���.��Vθ�8��i�E��ϟE��Q�q�±D�Z��:�q��.倬� ү=�mG7�)��B=�٣8a�3i#����n�j�D3�K.����i�7�����[(ɼضj��X�3ô�h}�6C�X]�|	{��EpTn�t���
��B��.����K��pN�ܤ�}j����[�}����In����OFߝT@����8GX�1 �1(�(�=3�b�]Wr�T�������Mlq�܍4ٷ���X�0�OPm��S��}b��ˢox�����؎nP��FlQ�v"
�2�V���۰�ݱ^n}�j�c�2#O9�8[�5M��p�u;Gg4EGto��8��VL�P�Qi�q�PyCM ��_��й&�]Z�^s}����]�"gMLθ)�Q`dϚ�^�BS�+����YI4��>�^�vHY�^��껐W� �O}̓��ϖ:��� �k$q��	�iq�g_K�Y���T�ba�S9><B�Tn�:��	7�@�^�n��z<�/�y%yif����ZQ�9*8��n �*D�����U�Z��3�[k��7�*��-ї:�=Q�l�c4�z�g���G`n�ثsf0�)�%���>P8+͞�u��J?wRC�u�S��U!�W����h�%˵��W}1�K1ƀ�U���3<�Ѫ�m�__G-�Q�1"���A�<c{5��R�/7�[�
R�?�[ư���)��4j�H�8���S9Ókv�������w/�-��[c�i�Ğٸn<���.�i�^���:�*�F�M�~np���
Q/e]�<u��y�:��U�&�L�Aȸ�-�"��Y���jÁ[f��ݛ��Q��:-0�6)���\~�
�jz�ᇶ��=1�J��q����/��+f|:σ���ަM,>�j��ӎ|tk܅a��x��4;$�|���CQ F�Sә�Hg
���'��r"������obå�uT��k���ك��X�LË�dv�����n��d�n�M\��Foe�=��Ǵ6������ǜn�gD�� ����;�Z��߻{w}�zo&m��Z�LUW���_J���N��`�;~�=G(�{� lg�j�]�z�ɘd�������*��D��<5���@`L_:��M�JEo�3��������8�B$�z!��U!J����5Y'�-�!��q~�$�~�'T�s�J[�;վ�0�Ά7�'��s�[�ÈGlJ�!�"����u�ˉDP��y`ڒ9������ʜ�2�q�.���W3i�v�*ɗ�u�V�=��װ�ff��4\��3Leɛ}	���-s��c�wd��(++>���U˞�^�G~o;Y8^0���v��������V����lt9��}:��v�Y)�52[o�*X�Du��Փ�p�q���R�YN��7Y��Q�_��Pw(�U}Y�
8��!XU@*�"�̍���o�O_]�����9�hW��C��wvE��ߣ��E��Is�� ����������[Թlڊ%ԥ	g���Nt�nR�#S�Gth7q-۰��T�O��<�M�ڑ*g�Z��<ĺ�	�*���d��/!�[ZT@}�׸�x䜡n�	ƚ�4�|Q�KˡOň�W�o�^��^�w�I(��`D-ɿ"�v)��/D]�"ѳ}��g\�+|�Ԧ���������B��2H[0/Զ�	�X�,�,�t��b������)�Y�v�8D��2T�I�=EGY鲬m�fM�2+!棵F�r�2F&�7��������daj��N�}��	4����+�U"|2ƨ8O�c�O��ɴ�}X<�.���ܸ��'�Rϕ�G���6�tN8��ijf�F���~�mz]�Ϲ��R�Xq k5�[7� p�t��U*E��N�C0F��g��t-=;�<q�㛙4���j�J������W����@�°��Ej!XY�r]��P���JL)f�rг;�֕w[����00OP�\�x�vG,T[��G�"[XI�Aε\3-ɋ6c�*gU��%�i�8䤠���v�aJ�]�٘�G�n'љU�Nފ�Շf_/�W���Y���up W{q��e�K�;�kN���,:� 3"E_���:q�5�ʐ�V����ͩ�;��k���E��J/	��&���T�w#/Mzk]q����N���WHVx���r���Ʋ)^_k]s���d��E��БB�ez�3��I�	h��>�\z-tA��dT_0�l�+�y,�<��dѢN(�8��=����������ƶ�|����GD>S���3N�`Dq��#���Ua�j
��>gv,7,�Ko��s*q���/����ЗneL,\�%_�kxL�83槰d�,s���!=?Y}�f��	E=m�]��(��h\%�V%����U���-C�`��LŉJ	�C�t�V��g�:�A�T��\�8z�Q8�h��;d��l&��}T)gx}Ҙ�7��`�2Db�Z���i-�5p*3+Hj�F�ÓN�D�x����^D��g�m����)�O�>Rnb��N<��~���vTMa�ܽB�_R1J;u�-�v��984e����`Qý�Oc�ap�:>#x�\V/ί"�>w�L�t<� `����&�H�Xy�C��>V,���7{�r�;ؗ	���VgeMX$wÊ�b.�7J�B�n�Zl��ͥu����>N����Usn���S����쳮ZH�h�����������D����w�Y�lL�9�H�'ڶ��+n�`�8�E�6I��\�S.`���^d�Z��#`��c{Yk:*�K�(�)G#�#���z���B��Ȇ�A�$�k)����$D	ͽz�rʌC�l�+V*�-����y�Ԡ��GƮ�t_N	SG�!2Bgo��6�^�}5G�`�=eֵ�`!��j�zυL�`�V�y֩�jHU����u����W*�k#�5�Tw�9��½�(刓Zڮ���k���G~��MU�̥{�Þ��*u�!Z��8Zc��阼J�Nߞ�zM�����꠪;:}B����3��}��v��jI� Z� t�M��mŵT4�g
��n}��^9��ۙ׾��s��S(O'=�+1Mf�T��8q`�.G��`7���.47:B�>ˎ���؄]��Ig*/�3P�qI��7{~��v����]U"��dAX%�`)8G��Ӿ����G�����8� �+^$���5)K�x]D��ľ�J�^�Zh\[ߟ��5�9�8ٝye��!�ʔ��{�T߰l�/%�q��R4B��<Q�`9��!C��;3P�ğ����Ggr`ŨЕ�9"Ny��ڨ]{����x5]/{#q�[���T��8Y�5
�FȾ���4%�Q`V]6[�j=��iҜ��/�����?n�[��;N��3����>J(9�J�6MdbTT�xG8�����=����m�bi��"nҌ��c�������s��(׆@	EN�1��BJ߷��//�C.�ڹ�s[��bA�;�s���^�{ؘ��[G�LLB��hI-D�O�f$-��FC|�T{ˮqE��t����J;
l�����4-��19�����s��3םQ0ÿ1.�цV���v�Z��AF���>I��¼|�"g�#��%^u����Nh2J�y�J��Z�]��Iw��g¸;������3}[�s�������G���'��E���d�:��j�ԧʼ���J���{��tR�l���c�m�����߾�m�>ߟDW����U3�OlvΑ$u]���Qi����(��*&�a�:�A]T�lc�"$7@��=�1���S�ܨz0��2��O�	j�$�x.�Cq�F(ɴ�KE}�Lc�xjg�7,>PaḶv�v*O��m���e����oyא�ТDzH��
NwԶ�Y���.�f�*����J�VR�����uo6v8�=6��V1!�*f�+͢GGZJ/���ޏ�{��y��|�c��0�����U/c��R�Ont.�#JQ��Z�Obr��܎EgU�m��NGx�d�b�r�\X�$��l���n"pL���E����2�-p����$~��V��z�[>2�ƬWa��̢��L�� ��I�}RD�n}�ܾ�R�+�,��v�y��}�
*�g�]��u�Y
�%�]{"�ú����%�5gfoU��t<�w�rUV�"��Q���z}��s��R[��-d�w�H�m���+��&�Y�4��C8u8����݇�n��7u*/�9���ĢJ�z��\�k�ki.�u�^Q����/b�Q.0�����$n��n����'a�g�i��Kz���k�f�ۆ����j�T+���av�;R����{�61�9T��.e�wG����o�o��S]0,c�h�5X$��}���G�sӻ
�nO}n�U�t��O^kgb+r@a[S�+<"-H�Qnl�$=��Kha%8�$,�L�wħ��ΣO��=k6��4�=�U�m�<:^���Jv�g��9�H9�P�-},u�'nM%T�u��d��0J�;d��QYKz`)���N��T�>|^��wt����{���K	�I=�j��_�4�=Yr��"Vli�]�0��1ں�P�st�X�
��*?������[a����qVg�ZK�׭�!�\��=�5ɚ�j�"�Ku��B�"������L���7�ކ5M�3;��!�-�V����HW��ݰ�¶�4��hP��2���鮴VQ�(1y��beM�m=-��K@�U�Hn����������nٸo�
M;�2JL�r�������̅m]=��u���[�k����c1�����ͧ�^�B��r����\����l� ��k�����]��.����#�Z��{�+S�r���jҳס������Se����L$������k���va�ؔ�H�,M`u�D[p��7Eq��:+���"�~���9�����Fˮ\�> Fe�<��|���o�m=��%�+F}w9���ٶ�Hd��^4Ufs)٫�r#z�߼�8�g�Rzgv�u{�jY���&��:G7���9��V�v�^C��O��{zm*\��r�MҐ��@A�#�[͆��[J��M�G��rl������Mۆ�oj�itv��Hy Ӵ<&i�JA'��*�ė{���8�-*�U�j��h޷#��.k�Y;��ҺP���t�R���:`ͻ�)έn�1W-�}''4�h�Ӎ��w*=����,�Q�FP�6 Q���5yg�%%F+��q,"}Bl�����M�_ʿ��F̖�n0��M��"e�$N�B��j�^�@4@�1��n�Ys���L�E�J��!v�����,)����G��M��O�&G �t�#=:#Kv�+�h�5�w�]:�0Y�E�٧�12;f�i���-����T���&�w�S�k/%�E��[
�(43��\��h���{�۹����I�S�]b�RB�9ӵ�[xb�t��x�r�����H�o0�.�L�SZxhj�u��D�ǣr����֑��ѕq�y�>F�o\�N��)tG(��Ȗn}F�q
�8�GM��Uv�l�ͳ��/ͺ��~u��n�ԛ��\�j�w.ĕ����+�t��y�<[���ܙ���U�d�L$p��?,��bx������2��C���䐠.`�֭��v5ͫ��]�B���-��5s��8uvb�[S�N��`v�9C�jr��Z�6l��z�;�����ky���Z7�(��ݎ���A<��21��i}�X�S�#��o�:���R������^o�)���N�q��[6�TF��̂��'�r�Nkn�U��[W�A�;�]��q�e@�Uj�L�-�yrg��kN]��mt�h��쬧3�q�� �vC�3�;|���<�qv�s��p&�8�����l�-+<��x�d?agmj�qԠ��k���/
�ձg�@j�_.Z�
 ���&O,���c��u����׵�?oϽ�߷��Z)R�ZX�	m����Qb(�1UUEU2�"��1�X�Eq
���+D��eeVcr�
+�5��E��%�X1��,b����°PEV*" �E�%�V,QPYV1�Z�֕V*�*���b�m�DYmU(��U���(̶DU*�"+��PU%����h�J�#V[UAAb1j�������U�+DQF#��2ZQF-J��Q�Q�Q��Җ��UD��Eb�[D�6�DV1��DbƲ����j�V"*c
(��KlQ����
[b�"",Q
�X��b�X�ab,���4D�U�EF�%�-�KAS-EX�R*��Ԣ��*�*
�X�[eh��QU���0Tb
��Q`�V
�YU���Պ5�
,PU�����"�F
0Z�E�E�1��R0���b��ň�Q���Q2�""(�BQPm*%m��U��娊ETQ�cA����DDV#6�V
����+K,�aS��o�o�?iˊ��u�l�6�þk��v#Nu%ᮬ�X󕶥�a�pvPV�3���<�U�i\�u�F\b�{����c�)���Vl���ƒ���xV�iS�D�&|�2z;�c���E!�i�]KDw�F��E>̥��YP��*!
4��_`�XId�a=v*&E�Y�xo��#��Zy�;�;�S�ڳ�{#�#!�]F����q��p��Q���%�H��f5T7�^og-W�|+!�r8���E�k�K�YȎ��Ð�v�J�k��t�2A�C���R�oR��ν�m���l0�p�3s��c�Z�vvQ)MoC�e��*��Sh!n(�z|�Zb1	��=�Z��ݗ{�� �2�����Q8��x%�3�S�U3}<o���w�\��ꑏd`紐5uƸձl������@B���k����zf�Ըn���(P�_���8u�x*�F<wcu�Y���f��Dww�D��\��
�z��h�tɬU�2Jk�����9D��F�lۓF����nt��U����ܐ���h\�ZUˉ��C���p��}�0WC�7�j
����;�m�!�{+����2Lk���
��5��waC�1X�s.���ɋJ���ա\� Ҡ4F�{�N��v��#�������[���m䮤[C�vhX�[C{h�OV�#�:����oM��"N�$e��o%*�ǖtMN�ԫ�ի��N�A!�� �A���ُש��+����&���mVfj
��򊱓����^���2�w1�����O�E�b��T|����9���%(�9���&b�($�"��p���8��B��c� ��ܖ��4v���I���}A�q�ޡeLცL�w���P-���������9
�껠+_["�Q���&��(JE?y�P�R�hvo{d���r�i�5�m���ࠈ��C��J6:q���s���&�*�q�[����Q�^��NK+����Xo�k�E�_��I!oK�;
X/��q�ߋ ?Az/|��n�����m�ֈ�ԭ�
c�V�U�����.j��]�!O��t_M�'�pmA�/fsfco9���xgO>ӖxC ��s��!��̊+!�Cቯe"����3#d�rFy)�<�k|�:cN��9q$q9��ww��aNv�i����Q��IA�X٬�7�g8'�|��h�Չ��#�<��1`��b�~���������K�%B�����ǝ��xR��4�R���J��5H��k��W)����~)�d�zeI�B�J�nK���.�'��W�:�ν�H���F��r�iusb�o�y��2)���s���n�)ݕv����Ɍ�r�2p����x =�V�ںa�5�~(��(�e�q@wUml�V�n����+r��
k��0;>�|�2{9�kMXX�!�謆N)� �z�T�ۿtr��!���w�7Q�}ᩧZ��[V�O��|'�C:�v갬\C�M�ڕ�iٞ�mE��)�ݏ���{�vl�±u�/ANp��'�>�4��������fV>,���˦���ێc��E���G�Q��A�+Z�)k� � "��2�*��z���
�y��Q�]@f�"I`dZ)��D[�f�E��Un��Da�Q��\LA�
�yѱj�-׏9U��̡�b�a
���Q��%GpM��O6i�;��%QY���J�8٫K���[K+��'.wb�0�;:G��
�'���h�[�z*�قGL^�L�|y��o��OѾhW]�<�����qE�����*4���ˎ����j��`�%�5/z!����h]�θ%L) ���W�K;z%����T��җ�B��'vɳN�i���- �ޗ���F����#PzW_B�WQ���ݝ�x�̑y���V�;ƴ�+��MrʚӶn�)�4gd�F!1,�\�63-�Kά��Ǜ�M墺��Xܬ�q��K���sB��!���ϳ\�4����E�\r;��ݽ�{WOu�������):J��3�����1���bU\9~�C�xF�b��2�eE�Ed3ey�5�S�+��z�6�C_���s����
=S����<��Q�q��(*��K�y���sJ���{�NS�Υp���aZX��3*4/��L���{��wu����S*�s%��qZ1�G�71u��#�'�j���$��DM	�0�;���r�xv3�Y�=�>�¤eu1����d#���ǂ\�|0����wP�ʄ��x��M���v*Q��*�U�v����kX��!��\ѲΪ��N�\^����*�������o}��T^��uo��,�E�eGE�B؞j��+]r�Hp�������
���8g3ukǤ�Է��p����}u��Q�<3ڬ�W��C��Aʂ�Y)��Ȍ����؆u�d����<�n��ƌ\�#����oJ8�(��Tҹ��U���h���l}����R����!��9h*l�.7p�{L�8��Q���A���%%�N���8�]_}y�bwאS�����p�����D҅8o��~�|>M��7���*ʗ�V��k;�$�iԋ@�<3�-Љs�؇uj��n����]#Nu^���&�=:h�I0u���O�MLe8yݚof�4�n=�Aڔ!�c�E��
*.�c����� ��I��x��$��5���Ot.ͬ)E�Nt�nRgC�fk��.:�~�H�ի�w}�r(I~�I� ��N�$��F���[�\��ϴ��%��\�� 
�	��?�s���A����0�&�sN`X�����X�4L��ED-.��~���Vd2bgm���~ゟ�W��*ڜ�D��w��-́�$�{'mo=�d�I�/��~�{��n�����2܍#
�j�#��.h����g�K�''��� ��V+i�7��T���K�ݐ���2v�L0Q>�#�(�!Є�Q�y'D��
��NA2���E�{0�e�Ss�4_d~�ߵ�׺�i�?z�V��+���a�>�E��4V�kƷ9z�h�XU��-sȲb�o�]�>���
K�V�_�8���Wf?,ۭ��	r�P��M��*�K��v������ϲ�͞�X�l��D����$��U���Xvo��-��*���0خo��a���K�����=�D�V,?j0�*�ٮ8ݚ۩�L:�@_�o.��
�o}�m]�Q���s�\ �G�f���֥�)u�C�ñؕ7A�4r��!3��NlR^+˄�@���V�M�Ul�ZT!6�B>�ol#m�V��7�>ֈ<ye�� �K���,!�/X-e���Fju��J�[�ථ�6k#��z^�/xRӕK�G����U��R�ݛ�Ԍ���ޱ�MF�M'N�r
����=��<UU�����u�uu����'�d��T�[!�Ӽ��V�ndF��u^� �������5�b57�[Y�5s�oʥ���n��69�܅ᑅ+�(�3s�Ru��ONx���ʛ�����(I�Dm�S�d^He8��8�B�魡�����vV�CMq^c]��Ig��2���Vˉ�18��F
jozp��3���m��g����G��ǚ��b�K�ql���;5
$���"�1�jl�:�|,*Υ�tW���ֺ�szwo�{9��w#�1�Y
���H�y��[�`��b� B�
��*��/U1���fr��7�t�:p�C	���=���4Q�>��M�a�8�e��}����.8��d�v��Tq��0��[���dX.�Lu���uj�J>�5=^�@�M^f��w^`�9�dC�ݚ���q��V�Z-�.�xS�b���h��q�6I��˓`R�sr�q���`�꾪�a�o,�Z�0��:��,�A!N�;S��_Fz\�7=��h=Ni|�(���%;d�n�����cs^�5�{�+�k	���:���3U��3zf�@�)V��w�3R����u����d�f>����_}��Q����/[��G�^u���k��ϝ.^̾X<�k���"���7:���Zkqt9!O�Grg�ɚ����{C���潦Q,W����]g¯�[���*�nj�.''"^6�S���ŵU$P퐤���>�h�>��E!pւn�t���֬��y��W'{�{q��f����i3�N��Y�〈��<����~N^���Y�1�:��
쭊��4�o�ԫ�5�F?T�d��1Љ3�͸�uCM��p*��M��o*�G=2�0dd��5m$����$ɮ�.��H�TQY�S`'�z���<���
�ӏ4z�g���m(}8�H�F �՘��&.���*�7��$4S�^ҟt�;����}��b;"���*��O�ܦSyM����C]wKO\ Jb��1/L�y���׳�v��/��[�wŸ}�)���o%�4Qڨ��R�W��BbB$ÎQ�B�8ڇU�E-ž�ko�(+Vz_.�dz�.YGh:�E���>J+�e�Ѵ���h�5��Bk[X�n����R�����ʓã�m;c*0��s����js�@R�X��nH�
���JAT3$ �t��U+��*��y��<=K�!;G|��f_X�9pd-co��EVk<2ѹ��ḝ�j�>���B[鹨V����%+��eo��ꪡ�+q'�O�͎��9�*lU!rt�/s����p�*Qݚ{8΍�Q����ի7�R��Ki���ߊR��~GY��+�Nj��~v�Y��\�mRu>Ld�;��x�d�cz�ڤ�OSW�8| �	0|�/�u�b��\������{g��b��J���$��ֈ�����~�<�
E&3�~�:�<a�w��8�>a���偉8�z͜��m��PSfsO�J�1�a������(��{�tt�=���������������$I<7�4�1
���k�.䬬�4� T����AO�b���x���ʑ����
���œHJ����
�$�	#�B���c�d����wR�}�\��m��_�
�ϲi"�S��g;ݓ�~d�Xz=|v�Z��s6�é��Ak湀m%a���i���!��ɴ1*Aֳ�:͡�mg�ȼa�ε����5��]zkf�r(�^��\~"V(<',�����>�1�& x���`q�q�3}�N���{l/(b
E�����Ă�d��̞���VN3��7��N�̲y���|`T����Ă���s9���<�7�$�I��c��c�'��1Ӹj� ��:��
�`q����ٶi�La�?�O�m���g�?��M!PR/��?��Y3�
E�D�9��#'�}��
 �����DwȪ�'Won�ص_j�rp�#�@�����x�A�xL}B��Y6{f3�K�&:v��i�����bAz��+�)�*=�t��Y�z�p;p%H.&�w�R��1'��uw��}���~}�}�/�8�O��>��R(�	5�����i�P��\�01'P��e��R,P�~q>���2T���x��Z�f}��a�t�#�>UV|	��3�Vú��%E<US�I�֗M}� q�<	���U#O����T��w�?$�1'�g␯�=C\H�8Ԟk�&�̘��|�L:¿> c��Èi*[6�1"�S_���������<��f�+����'��4r&�jc\��F�,\��1,��+1�>�$|���~M9%���J��sDO�%��B��"�Kr-VW_*ŻR�	�s���(7����l]��s�w���k5���Ѯܛ��n�@j�����g��2����ѯ����M�b������!�L���1����������N3o�
��;��C�1!�Y�J�8��'���}d�1��k>Ci�&�SH.�V�{ԛf���Lg��2VW�q=����.<�{��t}��[H� A �>��?Ͻ�@)Ӟ`vΤ��~{�&�?%O�>�8�R~g��~׈���S�y��.2W�a�sZ��Y.Y6j��H/���O�Ă�3���_��q��u���c_>�$F� �}�>�γ��?ShJ�]�`i��C�c<�rM<C�1��;���m�Z��q�|Ɉ���̟�\�`b;�Cn03/y���
E�N��y!8�Y�X�ۖ#R���쏠�}�Ҧe'���P�}a�(i���ɧ�AC�X|�\H,��3h(z������Ru��a�9�m �a�y;�<v�`u��>��M<dę�/�|�)��oM�|��0�2=�I��a^|�P�a�0+*n�?2|��'������q1<݇Y����v�]$�8�'�ɦR=��#���G��>�'�ì槫�ޞ�̱7��;�{HG�8|>#��
�����%eg$��\�8��Y^3z���J�I���:���,<-P8��$뉿o��@�T�<��ώ0*N>e��O���?~��Y�58�/go�)�H�<}�G�) Q�0�1��;��Ă�ý�[���1 �=��
q
͞k�`|�q����*T�1���CHc�����>�xR,5�~���s�c>�߯�]��K7���4��@~�;C䗗�Os0<B��&e���&�R,P����/��d�7��羁�n$��|a��i���CM`T9�c�������h(z���|>���9-wv_�qX����Dz�����҆������,�R,5�����=OϬ���u�z���!XT<;���`()���uۦeL��Md�g�'��|`T�C�I��Tg\�y��^j��y�Q����h�
���a�R~f�a�|�i���Rq<����O�CmCI�_�:���I�9���+*~z���6��VJ���96�T*;�4��1�����~��:5��,`g�p8v��@þ�؝m:T�[\Y��!kK��.�����=m��N:�v��ۊڽ[jT��n�[�Y1�}�ռ���ٜ�>��;H6��y�(�䳿�vNA08��-�����U���#7�b����������e������Y�?�n��%@�Tٿ�'�o�a���i�'Ɏ�~f �_+����3��ji �C�3T�z�@�~�͚z��8�}@��>�궸�t~��|�'w�]�G���J�����
�N��6}��A~C��3�M$P8��_��g����w��?$�� {��N�Y��2�߿���X����Y�<��M��i�<;��k��sqj���]��8'���=���O�����ɦt��+�AM}�<M��8��߰�11� ��Wgs -I�1�OP�Ax���gZ�`s{�$��?2by�'L:¿:O'ԛI�+
�3��{���7��1��

O���h>a�X=>�6ɴ:��>�����3O�
���Oud����w�h4µ'�~q�Փ�*�����bAxɳ~a�}C
���@&τ.%����9�������r�w����%eO^3��@�����{�~gRbJ�O�C_������`q��;�u<g̕i�~ޏ̘�������2~L!�wy��_Y~jAg/���\3������?s�>�Od��4�_��K��x�I����eAN��SL5�ֻ����:��*7���+=C������d��YR,�O��h��|g+�1R^^$s��a�kw��~��߽������=B�L�.��0*
E���'yq ���?=t��yLt��X|�M>�`c�f�s:���ĞN~���u������Az���4ϸ� a���M$�.b�D�}�)��y���>�x�{����#�@�cĞC�͠z��W�j���!XzkXW�Af�T:��0/��1!�gl��C������b�7d�+�����Aa֤���>�17��ާ�*vr�Ϙ߼�q�O�c�F����e���i���~��C\a^ q�J��:��&�?%d٭d��q&$�Ӊ��9�}=�$Xk>M�C�g������������?]$huGmb��?*ǽ��!���̜>:�DP��!����ﻒ��_��f=jAgX?S=�i�i ����T�<f!ܤǨPR�C���i�g�
�<�!X)Գ���FsЩO?+��/6+�u��9���֜��!Ƿ|�� �)��yæI4����i�N����ӂ�oI
Ԫ�`�[W�	W�z����=�)�u�K<1�ޅ���[���:JI�O���d��b[�z�ob�z�e[ؒ���6p�n�����W�2'v�,��[(����=�}YMK���u��C�8��ޅ�M����5�n�V���q��ˌ��֜&�2;�B�̈����͕��<�q����C�Z�X��0p}�,�6RBarỷ���ʾz���A���*���]4�kfe�Fɋҍ�*P�%��Ax��l:v��6�C� �-���8Yt+%E*v!�揌
�C�R�Wd����(��L����tw쮫��WM�y��Yb��ͮ�@�%�?��B�i�3��lS0��4��=�k�nPZ�ˋ-��w��O��f�Xm��QNj<�B�r7.� .��e�z�$Vdv]f�� T���8��*���CA�ki�_v��qN�s�	u�Lp�����k����e9.A��C� ���:�N�M���wgT�y]�=�4�(�=g'ѓJ��,��7+~\;�$4�#ͮ�r��+�.�V�%Y���4�V�%7&����_jMR����=h��	O0���dż����)�h� �����="��	\z��J��l+//Y��:p�$�%a��حEX��Tv�s �,K�{`�E�,o_1Pj�K�]np�m����+o���}��v��f��ef\kE'�t�ho(,�͠�V����$��_D!"#��J��0 *�p�	�R��bhQ�Q{tĊ�.(e���R�O2�4�,8���I�J]�I�j�#o����O�x����/#vq]�20rՇs*�1��J���'�r|j^$e̻�F�W"#��-���4��dN���:�IX��L3,�*x��O�N>����wPBȖ��Ct^H@?�4����ސ��I��ܤ�c;B�x2��8]♟H�
��*+8Uċ�-PW�Ą�B�n�Z��6�Qŋ�%]?��l2�	��&�-
�P�'�}N�5i���TA�Ay�x)Q�W
ƫ�@`,�]D��l�o1
8EA�(�9x1��) ��T+9>�V�xD�u��)-&h�7|{Oj0���9�h0ҧ%P�MS��	#�wN�-�ѫZ!)0=�x���9\! )TJ�A�Y��1�h�.�*c&�d���ڣ�/�(䡕�VûV�A�7��"�yDD0Ò��4b�ʖ�@�	y�r�D�E_��x�ն�X��-|�����X���3p�l}D~6�
<#�.���+���VZu�&����5��˺�$�`�nGe	�݊EI+�@��رiѨ)3���cF�D��A�a;����MB�s�!��;&�i÷�Q�z>�M]0;�!:tը��-��bYQ���@0ﳲ�ǆ�(W\n�s*���-Z\��ּ�?E,U��Qk
1�b�h"5�Am�1��
�R�*#�F"�cJ��1� �(��EF(�A�lr�"�![jQ�AH���V##�*FF�ԣ�h��Qb�A(�(*��
k�ڌ.4�U�V2�X��Q(��QQQ������*+1-�������*�-�Vڈ��X�0AQe�c*Q�a�UUUfRQ��E�QV*Dm�X���V"�Z�$Pkm,�TV*�0"*�����EP"��
%h�"��`�A*�ň1Er؂�b(�Tc��AD�X��#U� �UX�Rң�
Ȋ
+��e�Um�E���U��`����e�Ub"�"�*��H�"*#b�X�DUTE-�b����"*ʅX����DEU1�+X�1EPU�Tb�H� �*�ʔUcZ���Z �PE�KeP�UE,D�1"�EDEV(��PD#�Y�ib�Z��(1Q���U@`Vȩ��vԗO���ް�`Ʌ���޵1�{���ES��D+��v�=��nb����˹r5}�ݳk^-�� ���=�"*�9�:�����w��T6�_1��"���h|�������w�E4��/׈{��T+?0��[�^0*
G}w.$y�ɉRq㤟�}�ی
�'�Si�
篟}ι���<��rb�����<�I���z��$�8�n���H/s�<gZ�C�܇�$��L~C�����g�M�{����$�<f!��P^�����K>�{}�?�^}9Y�4�����:z��P��:k���m��{��9�I_�*����zSI�IU��܇R���y9C�m��!�/(c�'S\C���񬕕;�|p�Y Q@���?k����v�^.>�����v�$ĕ̱H��':}�y�R,5�~ۄ��4�Xl��V濙<�M$����ϋR/���5��f������������ {���P�q�T���c8{���~�߳]���j/�B�+Y5�������f��
�$�V
a`~C�77�!��T�&'C�+�6ɟ��8�0/n���&�u
�ɸr�{���(}�y�Z�3����W�,Tmt}�lZ�iuF�����#��q��V&��;�i��0�x�H-@�3�PP�X|��=Ձ��3�i1 �I�{���z�07��0�gZ�`q�6�L}O4{�aܿp����{xl�ܸ� 
"�����> bO�_��a�V�Y��(u��}C�{��6�P����G��e|`W��!P��q��/�d������=t�YěޱgXz��^=���ǟ�¾��]��kX�>� �qd	 }�=/�N& ���i�ֲVh�Y6�& u*y�2f���La������������t���N$���%g��B�Ձ�_�<���b�&w�ѻ?s���i�j"����r�����~}`T��s$�iR>|����g���o0��z�<$�S��+��íf��1������A!Xs�a�C�������A'��2�!54�ygG��8�9�a�J��.��06��Vy�Z��4��q�i��%J���iX�
������q=H-a���6��R���ޔ���~f&��	����3𱥰�eugw��9��1
����: t��X��v%��α	�,�.�Q �����G�����9۽ÀO�b�F�Ӯ�cPQ��#c���S�o4�4/�뛃�m�1Af������LU����������rW9=��謟��G�K>����<N����4���q�<;�j�I�<�g̛@�V�����$�{�4�L+���T�u��'��$��%C��S��l�f>�wy�����?sF�ٽ�Yv��-��@S��AK'�Q ��T;9�m�8�Y�s�mY�>L`l繧����!����}d�b�k!��d٭4��Rb�d�c�8��,�H��'S[��?q���s_=�]��xl�� ��&��'g���^�&'>q�=�&�u
���oǌ
�����~�h֤�8ɞY1�i�xM<`6���s&�����9ijw���<��s-��Ú�����잺f��þ٤�A!Sg�bq!�s�s�*a��T�?<LC�+�z�k�
�Ĩ~Cgw���`bN�_s�=d��0+<��H�r�M����J�'k���_�r��?�쮜�z�'�������T/�~�z�'����	���a��'$q����%H/��!�x��c�a�a�1�ʇ=�`V�����d����0��h�Q�U�9�7�{[�.�Vo�17'��~���C�=q��ed�h��&�d��퇲�ĜC�d�~q���,��>���� ��r�J���c'�w���������H/���&'����l��� SS���n����,\:^a�c=t�6�a�J���I������?d�e"�F��~I��KL@�T��󏇿����B�g��O�
���1���k �����j�����&8GS�F����g����I߾�4�dR���p��<H.�k��He�X�Ϝ�Z�3�16w_h�6�^��X)�!�
/����R>��8����g���@�#�Z~��Ϙ�&$�f��'�~`W��M$X���y���'���R��z�� �Z��'SI��r��8���?d�m ��k�4��R����M��l�'�m%X���|�\N}�}�GƐ��W��<O��I�L���UC���3�9��m�a^�3�AH����;0++%w�d����q�힞o	��C�d�g�4��A ��Pڇ��>����|*�P��2��ghaݷm�ꤞwˠ=Y̲U������8�����Y��l���O������<'�z�����=�j������t����8�΀{x�v����%�9;ZҰ�%�*)��(�+Gٳz�N�.�?{��z��Z���މ��q�2G�#��=$��F�,6{a�Xz�0�N1H/Y:��
�`q����f٧�1��,�i����d��p�'�T��w�]��5�G����i��#�����x�����,OU���@D���6h�|�@����?&��
��J��_��+:�{d�OǷĂ�J��4���^��������8�@�8��g��� �T��w:~:�^�מo�>�w�߼�y"��ĝ���Cc�T7�a�5�Wf{���@�T5����'8o����̿�=AH�I�n'��d�S�x� �'�s�?#�(��r~��x+)��[W�ޟ��
���S�s'�u� �i�5����@��w�?3I1'�g␯�=C���H�8ԛטM��1���i�Xo/�
��Èi�a^��� <H����ffZfg6�>�����߳�;`VT����z����1��g;�`i'�Y6����,�;��������d�%T�Oɉ�w�i����f��6�^2xo�Av¾�˟
>}��='��t+�~��U_��J����7[G�F�z��G��
I�*E2~�'Y;�
E��tΤ��={�&�?%O�:�51������2bc����$\d��7U�O���1�IDQ���R��#����lĂ��� �P�<Cd���3��i��~04�N��1��!��eN�L�?2xs��u�8Ɉ%�SO*~�^P|��$|+��zg✋V��_M�uϿs�y�y������g5R<d��Z���Ajn�O�>O�i��l�L
���.�^�!�Ă�q����7�jN��=Nw�x�^�����#��|������)ή���{/��������=M?2bO-8��0�Ι;y�I�+
¼�4���C�}˴��C{�H|�ɝ�q?:|`T�C�Nnì���P]�w��q�q�+/�����+����	�j4ݿy;�n�+'�q!�
0}�"O��a����y��z�� z�0�+8�&;��|��Y^39I��
��3~N�}�%��`u�����HJ�'��>v���8�	�5�y$�o}o=E<��e,]G�lkW�o�y�j>+I�>A Nc汘�r�uk%k/^�=�����n��t������ߦJ9s!ђ�kU{Z�#����\��Tc�asQ�u�����ѴEࢺ(׼��d�V�W�Z��=�P\�8u���猷�ͮ9�۱ї��0\� �B�+��^�o���+2N{��֑��'f3�͆���8;TEm^��G��m��{��{މu��y�5�5��p��D�>���% ��	��1���a��0��=H.�9�f�:阐|�(�>B���XE�泌�_�6�R�h=�x�`�P�Nx�,����>��(\et���w��,Z�!�hi���1�;t��//X����
�̙��x�i��w����d��7�i8��Ak�w�6�a��i���q�P09�0q���x��.>�[�뽋�Ψ]�)�!�x�����&<I�1S�JH/z����2VZ����m<xɈ{�k�Ɍ:»t��6�J��{�{l ��m��� ��k��P�g�K!0�����T��������۝�lt�������d	Q�"�=��'x�y� q�}���2i���i�����Ì�d5>�'�0�ϲ�p�HE����.�{���?g�~���c'��~��M0=k:�����%@�T���������:��Wi<?Y����C��!����ϐ�SI���C[���b��W�`�q�:��lQ�^U�"��k�Ͼ��w�����g�i�I���Z�`��|͜�m �C�����:���O��&2i�b�^��}v��W�2��=��m �M'�<	��ٚ�M�p�T��W�����&�]$�y��6���(i�������a�m�!�<;�f!���;�jO��h�p���<��l�%`sˉ=B��Y17�'G���!
�{��p/�s��ߔԷ���4��+��iݰ���փ���S���d�Ci�Xzw�>g��I���>��&�_��`x�O���o��4�IU&��z��^2o~a�m��$�W�Pz�D��_}��|>{�F~aP��++<'O�6�Ĭ�5�ߵ��8�T*zj� �'Y=�;�&�k>C��_�%@�w�a�&8����y��+������m 'O�	�>��ן+�������O��^��OSI��y�kt>O�Ă�jN'��L5�ֻ��8Ρ�J���O���xH/�z�{v���Z��Oi��Ɍ/5�4-Ph������)��+,�>��U�Z-��*�N�X�㛅���v�X���oN��Y��>�nӣծ�,���J˧��7WejR�B�5�&w��諭����Gm�����U��h���3��&7�@����%��^��\S,ޣ�����ݐ����S0��I�W��л���;���8qJ�Ih��������}Ō��~i���˲��&�M��el���5����()���ǲ�Bp��e��`��q��}�}f�jRmn�,�����K��rϴ�=�*�#��y/P�q �żH�l����vSf�L�JX�#����i���ǖ�':�>���
�)E��<��5�F���V�S����x�ED.��d��w`.��Ȱ]Ƙ��:�Y��$���m�:e�{��|��!�X��=�n^t�sL9�# ״��Kw#M�0�]١��sg�ʋ~��&5�Ɍ찱r#�U{]q���Ym�=��Y߲��]�e>���~�[C�����d�
ldp;��g��e�{�Q� ��;�/ab����~�*�v�j9��_,�쬂�dB�CV����0n[=`��/�{HF�f��l��
k�L_$)?���4N�U���ڍ�j��OlԬfj��R�d��$�Xx���Nz�i�>���^,�eG]�]��;s��N�=D�hu���D[����c������ݘ�l۱Ƅ���ы��E���D� �"�eA��Q�{xF�%U�&gE�yK��ӑu<���x���t7��_�󷓕�7�;�W�p�:��m
vHsa���Ѭ��a�e��s$$�r�Ċ�,k�<Y-gp��#��bx�~�U�1��m[m.���lן���ѹ�n.��"}̹���H�j��8��>�&�S
np8�n�@�(���quݻN�s��[-{{-�S�D������]�#���|%���3Y���]��]�2�U����G�"s���#�rku6�aں[5
�Bg�Ϻ!=�x��x�dR��Cv��ݵ=��3O�돆/D�-�X�=�-���w�A�5׻���j��3��D4g	�QKj�n�Y����B7����b[�9��Gc�g��#�4Q
�B��(#����0�p�u��־��Zm
$�J���ɐ��n ������ݢQ�u\υ���Ac��K2_�ا��F��Ȣ3B��+�����&ʐK�N���!uUY
���(��J�61�8h�J4(h*���UGn�%�����	����Uc���\�ok�gmzxL�����w�n�Ϧ�I�tO�L`��Y��m�����.d!���{��O~�����E��̫G�=p�ݙ7:���H��R�0w�C���nq����Ї:�;	s*^�`�]��u0St��c���U����T�݁⽍�9�q$^w+��ge������b�uӝx�ͭ� ����1^		%���>E���v?�tӡ�.��Y�;~�1��K޾��F;�g(�`F͞�)����b�Ђk�ĕ�AȐ� ��#3���$��J�,�=���r�b1�u��y%M�Ms��]�:�hGUu�6hȎQ�v�C����ڶ~�lz�������l��0<'Ǘ��F��A�.Ѭ�U5P�tJ�HI��Y�|�1LBv�c��:���.#�Q�v�K�9&6��>���yi��{F�Oޛ��
3��PŃ�S�"�d�5����X@ɗ��u�GDC��}���)3�1�g��C��j�? �H��p�k�z��qb��88�ڱhM��~�g��4��/����R�΋�rb�nNt��+=�	�9^��.���vz���g����JTK������[뷙�6�,�z��Y��0k�!]�y��
�]>xخa����'�ej=�V�ٰ�)%�κ"�Q�ϯ���L�s��u	�g^�@�P���,�yF�wJ�m5cpj���H�Qv��!q�1�b�o!����ټU���塞�� ���m�W�p�o#��.���8�Z��fl�u��Mqr���JV=�@_`Kj�m곝a��ʮ7O''%�2�U�^<�$��]�#����V�'�����!��X��E�e,ڒ3��8��gl��(�tB���=AV�S�5��qc��t^�"�F���(�2$�k�΅��f���݅�,Ᵹ�U3�;��CIʙ�`8��x�D�~��{��2����H�n��[+���D�t�k��O5�E�>Rr(s�a�<�r�����Hy	�����o��\6�Kr2Pc���:�y�9�m̍P���Ȳ(ԺV%54��~��d��N�3�^�4.��MU��%�.OR�٭�����{c2��q�"��u��E7v&U>o���S���2w��5F�	�#��U��Q{�T�C3�[V���لp�2z��f皢�c])�Z��5QN��ɯTqɊ!��f�"����9��A'D��B�$��vv�_OL��j����G����Q��f��Y����+�Vt{PU׺��~���<�mJu��o^\��8�#Od͗���(A[o�״Ê�,WfS�;���[X��`(�Go�h��S�y�ot�*y1{ ���xȋf�wK�o!�3ׅ_�2=F���[��>ց��ȭ�)��p�b��6�vr�l�2�S.$�U��1����g���%��.fP��Zi	��!Vou��}���_!*�ڣ��L*�[H���U�sO����Ｆu�]2�g�fH�5u
-��E�
n�ۮ��²�_�)���f�I�Da�Q�ޙ.�6��s9_�K���5p� ��\��d@9��O@�j���>�+�=�ٱ�OǶ��Βq��&Ger�RWC_HG�H{ׯ5�8���a�9MYƺ��h��`Ī=�za��Qk��������TN�K&K5�;&�J#;��m��kU���9vfDa�GwR��T&x�D��
�F���d{ 2�X	�q�m�a\c�������zخ���R���\B۩0�MaE`U��g��a�"����)�{��9��N�������eq�:|��Zrȯ)����R�Wyy!�.`t��Oq��ܖ:�Vy�ڛ�`�4�
3�J�㚄��͐2_=�E`��"��)E�2���zM��=�R4��}�{��d3b��P}b�i
��{��bx��k�v�h���p*В���Y�ۄ�ۺo�c�K���= �<zb�_D�2Bw��
S#�.�LstNh�O"ND�Fcw*$k"���CV+<�,`ހ�ǫz*f5oy�
�)�cu�]̋��K��]����V�)˩c݈�b�k@aÓ�R|��WoT�s\��곳ip�}bW�%ԵVR������u�X��f�!O*�K�%'Z�Kwo������+�{u��TY�Ɣ:O8�+*MR�gp��0HDN���y$��>'[�	�������r9�K lˈJ~oQ�*�k��x���1���𖨏�T˺����`��{47p�C��x���	�V�*�W�Y�L���0lOW�6�*��B�v��at�NOTэeX�"}�"ڝ��@���X��"	��u/��!�ả�t���(V�[�+�f��8��8bk2�v"�]3$g��sa:��5���]�Z�u-t�:4/Ɵ����a�ڸm��X��'�j��N�G�������'�����,�9��v{}����F�mTGgO��R�n8/k�A#:Q&�,ӊj�qq��U�e+��l�c����S����-^�ԍ嚭"��p��� �z��������E�^KϨ�v_��؞�I�{�e�9��<y.!Z�#Ű�Ć�����իL��Z�ϳ9\���8�e����Z5�|��t1��+���3f�3/���y��w<�q��4��	r��09o0v�N,���Ζ��B,).�r-�;��Q�-����V�A�{�k1�]n�m�u�St]+���ȴ��9��+���:�3X�J�K���.]���o��vI�)�3�e�Y�V�`2'f)	�v*���pi�`�{�j���c��,>>��9Y�j=؜V���NF���IX5˛=���%b��mHe�;�q��T�uov��1���\�f<�N%h^�,vPA,��(C���mgٺV�x�(��or��ݠ`X:�1��`�1u����4L�*Ѥ=f��S�W@'](+m&�q_ƞ<�:v�9:!4
��L�ݩ�*�9���	ƹ�^@sm��Ǳ+|���,>���ǩ���X_XKA�w�[�WT̊��Z�U����8Xx�b��4#y� �H[�Y4�|�>��	Χ�q;ҳ�M+t��m�6�:];6ȹ�k�K$z�
b*-��eu؄WSY�Pe@�5�)[,�]]{kN&32�5�5��
�t�M#�c�����YԱ�{�e�]�iCz��4�7yY�C{^Ğ�O���o2f�ʜr���d�&�e�r?D�;��Í�׆�>/�NWj��.f��b���pb�sGsȱ������\� ���lN�&c�n�[�.�
�b��u��k�����}N�`X�����}�u�|��X���y��LW`�n���rjb��g1B�v;ǎ0Рkh���E�1���;e��,�]��R�n�щV����������t6�,�j�e.��0�O"ݓX� NfGo*+4���,妨	�賆ܷB(�#n<�0⅃n�M\�.�����ʑ����K8�b9�'J�"��Y���x�g��t�+�sn�<6�Y�d���``�.�N��/$�hA�I�VE�̐+���X��&d��51�L�*`7F^!h�v��̤�Ȁa՛I�DP�{�t�b417�Pv��QP��J�Rk�F+4@%P�zN�t����бM]�E�u.�� �
���i�A�l��)�$�iY��T�E��:��v�É
И-ͼ�n���"VΥ����Y�5��0�]���ɉ
�%�(S��ŋ$R�n�CKp��$�:O�[�rnlP:��U3z�/]��J�):�<���ձ\t�yDh�fi(>�EX��Ȓ�z������x ��.H�v�x�.�T�V娩�K*%yEK���a�U�Ւ�����[���U���_,T�<��]jn�H�*K�����%�I{����I��V+��t�\,ƨ���3e�W��LfZ�ӾΆH�#���A0A���"0D��A`�1Q-��VT(������Ul�[h����YUEY�(�����R(����",Dm��+YŁhڈ"�l*�ULh(��c*****��X�(*0EH��
��m`��dDb�(��UPDE�,T��Yj�j���UZ��*���\��b����mb�`֪��PQEPEDTX*�E�E�T@E���QUPA�j2*�,�
0UUU�(�0U�ER(
���U*��Eb0ĬF"�Qb�Eb����E ��J�����((�S)jX�`�""1�TE�h�"�`��TZ��*���QD"*�UT�F"#
���U"��E��(��E[e����+-���X�1�EF*�Ř�QT�¶��g۸��~����G�����ۚ��7e��H蓊�@cڝ*����p��ۆ�yh�aNZ�o.]=c7w��}U_}\����G�l��E�d���D׹�_����>}���5��\*���
"��:����q�T�nI7��R���WIc{����-ρ�7m���Lͻ��m.��2�8¨�4��%>��u� r}׬v�bΗˣk�b�jf����5����%�#�T4o�M���>�;��k�S=�T;��v�sk5��4��+�7Wy�5@\�6�ek���}��>�&�V+N�o]����.���m7qR���2F�V�O=���n&���/�eϵ<����؅b|۰^��x�V!⍩Xl���o�G�cͤ�f��L�ϜsӘŹOW�v�L�:!�|�����>Sz�D���_���%�3��]g1<�]��������n���w��/�N�Y���+]�ޱP���ǋ��� ����SSX��;V�Uz���[�b]1���j_l�Y��3�pbs'M��Į�� Q��ۛ���7Y#�|*��+�}�qbk�$��c5h4��r�'8���[8p�8�rgo:vi����j=E��}Y8�+9����<��� \�k�z�k
#�UlOK�K�_��U��X|��Ÿ�ƅ�<����7���9��r���c���{ny��7�vÓs�pr��R�j�É�S�����0by9#oX�ұ��}�ۼ]�]�|Vۜ�y[�MȆ#p���/;�������*x�κ{���F���Of��=����K�3m-Z�~}x�^K:�`5�9�|���.[�;���U�a�ͭ�wB}��ꓱc��*xuB���5�|���9�8���o2m�U:*vSs��7��Mc�U�YУ�AP�i!^3�,���7��בΐ;V;}�QY핸�ɾn�w��n��sBt��@�<w�M��|-R0/t�f�_w�>�p��򨎔KwB%���lmS��ۈ�!�d�S�ݺ�x�k(^]X�{�@���W�����M�T�(�h48�ZP�Y��0l	��e��S{[��4-4�o�%4~�R��7Yͫ�$�����5��&�.w��5.4zI�h�U9��Ҿ�l�F]�� �}�A�bo�)M��)�� ŕmk�1�
Ko�wEY�v�l��v�W�j�of+��v���3���<��K���
��S���{��.�5�HF����,��K�ǡit{�6ef�o<������n���&~Ws9��,��\�eϹm+ �n-�z���(���6��ז���w�P�	�iP�≗�8��+���=�����ǖ�ɍ���v���Z]Uè�c�t�JᲳ�G2���l%�ʙ|�=�{�E��������w��X������������X�|5����g%)�����O�:ɼ�.�r������] ���rzA�T&��!V7 v�V��6w�6�{�iN���Y������.�;a���xr������o&���D��d�s��}b��b�X�u�ұ��OR��4��������	�j<�Dg�'�z���[a�!�}Q��J��լWJX�;��8�V�P��ݝ�.{��˴�p�Y�+WYu�ְTj�p�_� _��:.n��4�.��'v�������s�jtRF5��=9�=�Vcg�7X׎��]HÌW�ͼiǗNRm彼�m;�ce����k�v��t�d��ƅ�U�a�aD��w�N�!p�Z:n����{����5�u������l-��Ok�k��� ��R
�ɩ��̥��ƞ���R��Lɵ�������~�1�ov'�V	O�p~��ځ.�hmF�U����Pg/EOj�iu	�]	6߫�P�H�]	Éu�!�7�"\�S��v��>��8�Z]8d�'S��B�í=͌�q�ޚ��]8�r�P�\TX<��7b���(
�^����Y��R2q�Yԯ9��ͨt��
9.����D�윔�E+����2�v��ŉ�s���<��VߋA�±!�B|ո���Y���MU�ն۶�ڭ�"�XŒ:OOl ��Cj�؆������LQ�k�UU����KTN&��O��� v�*��{V�my�qT����^SWJ�f��x���Z�0i�]ǆ齎�#������m���L�e\d��܋}W�t����0���3pZ1;�r��ݼ
b��Ϗ`VU0���I��|Bz����{��|���g6�t��ГP�����[;͜=t�%Zt�����q_D�����n�YqU�{��כ��uh���NW���K��?'�蟩-칔�fP�j�^ք_j˦�N��᝶�;j֡Թ�X��;@7�vܛ�&���|�-Ϲ5���3yc���v����*j�l�)���כ����z�!�]ǌs��'y �|�`n:��{7|�A��<Q����X�T�ҿ�~���ѧ�B�-�������b�ʜ��l��5l����}��a��t�UM�W.y�.�K눍�B_++w�܌AwX� �o؛�2�u��Z�m��Ȏw�s��U �#R�[]k����[Ǩ�n���k%�g!�mc�U���%�rѲD��@�u���uc�]��i������/�z�o��>���iW!�5C %Q�%k�+�dÇR�3�Fsb����u�^ˬ�p����z[BE:q@B�����-�PJ�Z�U9�p��s��;����'���*d�ФM��|���w9���m�=�Oxj��e����S��lWSg7�����X� ;tevv'��t��mr�[oZ�8\�l1����t��y�1��<O\s/8%�#�Dw	C��.W���5���/n��WS�ۜڵ�wr��k��>�ר�y)�zU��'_\�����lLW?M�H�Y41�Ւ:J��Z�1KG�GB����������uw.�����tv�f^xK�5���'���0�~�F��e�G������~�Z�i�%�Y�,7Z��.���ӹ�����bf$b6[�Pm�h���=����k^�[Vk*攇��PrP�Y6�_�'+�'��V ��f�u2��7���S���-�4�Sxwmɹ*��*�z�jX�U[Efհ��1�3��
v�
�Jǲ����C��+=v���Τ���I���=0T�K�P�y�k]���Y:��GuZ�aH�����-���kl{li-��tN�[t:������Iwj*`�6��؃��<�T4�)o�-���ġ�NLf]�y
���A@� Doio�9��r1ؗ;���ֵ�\�H�ϻɘ2��~qgO,�a�ܻ4w%�aup�K�颐f��G��Ι�>�6�zqj�n���V�oo�$�c���g�������9�@d�h���v�p�{����ˍ�;���Iq[��牺���Z��o?VCO;�p�[�v�t(�Z�!�{��]Gm{2	q������Ѿ.N4�Q��:�6:�����$*��m����VCO��,v���yuzw]z�7�V�p�S���zכ��9;|�g��*v���U�A�Woע�7��7c�^��4�}�6���b'}~��4��!o#�������q+r跔0+�V{��
���a��L�E��xa����Z�+jK�`���u8�e�MX�hW7�Us�ǻ-�{i�(�������7kiu�{��鹗�㴪s2�J{7�g'ؘN69�a�����1ԗ��^�sB3CS�捉�|��ߟA�u=�R���N��T��T5³	씷��Pyi�SMa�|Nۃ�㘨6miP��&�V(��Y���Q^و/DuGծyx��<���M7�Y��aef���>ݠH��V�^�L�8��!��Igu��~0zƫcҍݏ ���̼����0+n��M�O	 7���{bV����R�1���R�e��3���42���"Jq`�(!ZK��5��w������t�uՈ�bw*��/b�d�Z���>�>�78�t�!����C:V=��OR�Qaċ �b�0�D�����=�I��)̣�rq_�F�C�d41>S�Y�>��������ӏ>���%x`u�:�
��r�ҳ��r"��b���RR�9�U���߻�W���SPz�m+�MϢ7�/��Com%�"q�{�}��ns� ����fPmm��`��MC� �F�ՙ�BxV�c1�W��+98:�_uR�%�Aw_��x�Hn���앞��=0�Cv�4�b��k�ul'�e�:��J_v�C��t�����'�����T��1 �}70�/�9��v�~.���B���2Du2��(�(F糅p�~�`l~*��*�O��pL���r�g�&ef�X�g5����)�Tʗ �I���ƀ�.�~s�ѫ���-�r)#�o����x��PJ��>O6Wf���]z�$M��KOR{��[.�������$�O��َ�hӻNpkk'��ý�+��%n�{C�՜�S�m-90G�ʍ�]B�P�cy��w�NN���m>Z�N����-�\��n�E_�W>�;0��
ķPZ� ��E*���=;:+6�Cs�sX�ٮ���c���u�}~�7A�s�����r�PR�(:�K�M�jyG۝��:!�����%	�����=;a��h�V�eؼ���e	���J�{z�	�`l�'1��X��>��P�t�\���;5
jk�.���{{{,2`�K���}�u7�>������sA�#�>O�D�z����my�{T��M�9E�-��w����jY��_c͠�3�W�����
�i��w�A��~�W6�+�5^:�����f����E+�gXb��5{F.o'����=���6��J�6���^�5�U����{_*�'7>�ߢ��jU��X��v;{^�������z[�nN���@��׫���b,㶱�� ��{�1��w���*DB<��O�����,v'�@�6|�g=7�m�Y�˭U���쩚㩒�uA�i޶��֖l�K4Q[�q�.)q�q��q�#FV��m�ވ®V�U��B�>����v-e��+Y�זjܫ�+zqv�3�rzC��rjީc��������.��R솨���'�W��3upM,e����ۛ�i��?Q�u:9�%uB�#���ʄh�py��\�f>N��I��[k�R�4��V���JϷzh\��I;��2i���[�����r*��~C�8�zb�'�ƫ��������e��Кn�8#��ps�#���f�jy�x��z��f������d�o�X��O�v*8*��hp'N9Wd��j�<�+����$c����Y2�7��1K���޹��UM;̕��_"=NL>S�]|�Wv�]~O��K�9�>�m���y���ֲ�ӹk3P��7���w��}���iѮ��*������1v d���/r-�wv���ܳX]8��N6����/�̧%I�U6�]d��^�Vw[ ?A6,��z�.�t�T�z�]��佳xú����y:�[���.n�:y�f9��-�usZ��7��X;�DF��῀U����ڻ㯌�������� ojR��
E���ʳU�rmf/�
�ۼ�@��jq!b��:Gؐ��%�[g+qV��
�t�L��]���w`������<�Ae��S{G��L'�"�j����b�r�N���ĳ$�\���D+��L��/w�.�벟l�Dǃ���L4�=��Cp��cz�Ep����%�w�C������s=����F)'w���=��S�I��%���ޡ{�e�Dt�
2&����b{�M7��K-N�u�ei�ͫƸoӚ�l�nd�=���ؽ��nC"Wu�Z]�=:�.J�����f)��n�Z+z�K"�3�ڋ��w������� �͵YI.-�k�;������X�Ԡ�٣�3e�t���	����94')r�&�qV� ƾ�'1�J�hUp+� �ȸ�c᠝Z�E�������ۃ���zU���f�M��b$�N�ga���Q���N�T;��մv��YJ�i<ب�%m�����,Qw��\9du�;����F+�P���^h��ʳfl�'KͮT�l���*�6�t�!�wkfXM�|��"a}����Y7��C[u�^e����0U�~C�(U�vt�傥�=\skqK��W��aM�	�3�u����\W/*�A"v֊n�ٖ3���v�����ҹoj�P[+H(FݑLus���F��թ>Ŵ����P�ڦ��w�+�ԮVM��MB0���y]P5��͑��.$t^#�֎El�0�l�M7W��*̙�Ӝ���2]�bݰ�|zd;;���gI�%�F z]��0j��-�E�r���Vs�����F�SM�*�ڙE���|6�GZh���u˶���Y���͜���-��Kv�<�`MV�5|S����9�㻦U�KQA���5ٷ(b�3���ɺ�J|��g��v��Ai�ܳ�t���v�;k.E	����*̮����1g&�*X�;u���|�/�/��.ϙ4�m�m&e]��7w�1���ΗCU�b s�%V8�z��&����"��rٶ��_ul���c�oS�A:��w%-:*�W9�� �Wk^����_���E�au1x`�:�ȥ-����ƥ����V��4	6*d�u���"H��;zm��\��v�YĦ^9�*;z���v�f�^S�C��N�ܮ�g^A�\/J	qM$*��6ldWH��F��v�7Z�g�iQ3h��V�ʹ2�o:��A���ךh�s|5�^S�0eiX�Y�2�Y�Q���U��/T��x��"��
ѽ��z��BDDU�a���Y2�,��+��Yr��сM���Y&>�_��KU�7��B��ǋ�M�	
B��z�>8&ٗy�4�9��wۈ�B��};k�.��ٗ��3�s4��>�1._$׃��/INS�H0Er&�o`/q�i�z&[�"*�k���U�E��MK-�O�ᡗJ�n�H�e�}x���]o7�y+2��iv#Xؼip�gc1�m_!�/aca�ub��7���H+� �M�7]O+'o����|�t��'������K���߶;�D��X1#YT-��ѶE*�ŀ�XT����i*�-�QQ�*��\���"��*�i\Lʊ���U5��
��DU�bF
V��Z����(�R�����Hۙb�R(�X(�S��H��b��[*�U��AjJ*
�
����AQQF(�-���EPU�DX(#[J�X������bE+X�A���X*1b�(�F*�T��E""�Z��AEX��UEQU��EX�kUV�+X�m��mb�b1�amQb�,"�D�UB,UX��b�
6�*�"��#� 	��ީ�B�+9q&.;�q\��a��݆�=%J�׋.IG'vt�i6�Х�I�7�֡Ҏ����4=�s�8���oNS���v5Uʉ��3P�3��a1n�GE��z�S��}�W(~mܖ�h�� ��Ulґ��/���ٌ�����1�&<�:jX@�:ʴ��veQ���{}Pq��Uޒ����9ZV]����
��e8�b��wQ���ʆ\�`��@��ܭsf�F�q�v����t�D�ڣu0�D� �,�����OvI�l�)��w��"����Mv5p��uU�ݡ�!��r����k��S����-=�7�����mkc��=��(PQ�$+�����n^�;zf���qɹ���˦I�x��}׬v���� ����%Y�B�7�1#L�e��a�-o�Kf��Y��1�n����7�V1z��^�^|�������3"��mf+oo����� ������K[�xy������%=�JX���f"<�&�Ld3u�9��7r��<��\�er�ASq�sU���S��7.���&D�Ӵ�N��K��օr:J�� �++�4�f͛	� ʝA���;=���ٗV5V ��ov�̹-���Mg��*l��3�[�jh�ȣ�@ÉǇ�%��������5�u�{����������)�k�������-;F������ɲj�3�P��
�sȫ�A���W�Ӎ׾������Ս�����Oٸc�6S�مI%nЬk�'��ӓ�E�VFL�4f^���wڪn��>�����5;P���9�w&�xR���w0�3���q>{ױ�U�SE�)}9�=�0mjg}ʆ��^�o�\�t�騼�ujy��a�`<�,\t?j�X���<���Li��pvi���?Ql�T-�Og��W9mb��T�����';dT=3��gg2l0jk���g�ѯ=��b?_{�z�r���J*"w@�^�
�g;�J��ѫ�U��E��mmt�;�&����&��B�<������tU���u���%܍C��؃ݼc$7M��pxɾ�P��V��6��4��[>Y�d������*bZ9�~L|�'w9<I`���-�N݂�u Y����N��݄����"�b\�Ⱥ�U��z���(�,��\j�gح��h�eZ�n�*Ay!.��6��6R&���Jz����{�m�u�oU��H�C>����Ѻ�B}����ۈ]q9��=6�L�]qu�a5�Jr*��i��]�xS�E[bEdڭ���$�)R����X�ۭs� �O���٤�u>��,�+��i@K�ެ��ʹ�f���նv�_�7��T�R�h�ݵ��c@tY��C@�x��$�\��!n¹���r�E0����!3A}�4�����f����s;�s����i��ܵ�=���o��&_eG���>M�o��7}1wtm9QF��y*��$G�S�c*�zfx�8a�W����R���{X|���MY���$�*�8�szm�5���D��n��9B��K��{�7�}6������'��o��}1E�����1֡z(:��-ST���wE=�ֵ:������gs\�� ��VF��0�<)�]���A��#��������e���c��:����Y�	�Ӆ�h�Z\�ђJ��nW>.�����ש�?T���6�֞.���<��T�}��V�-7��+���z��J��/����dѮ�wώs2S,eQ�(������-LM��"q�UW����Bx[�߂���V�Og����m����R��h�~y0�yNs~����f�V�v�;�R1sy����oi'x�}Yҭ�(��mi=�r��ڞ+����0���Z9׮;�X�u������5�⤪1��Q��P��[�[{Ұ�k�n���Ѣ��3�|���7#]�1�j�F
#%��ƚ�4��Od�	q|:� *����w���k��O+���	�˔���Y�j����T-��U�˷4�P��A�"��y��>�n�{d0��]�9�N[�ޡW7|R�2iӊ�F�>�����&����4�&AG���mb���㛕����]B�V{���l7�BT�hC�����ӹ�K����Yb+�srher��+�̹����ۅa���d��lMס�􀾉a������"S��nwڲzJ���a�Î;��vv�F�[u�����еk��u��R'&�$�#�k�9��=���N7�Q���z��-��7�0J��3��1,�K����������n�G
�cv7y��[��QR���Z�=7Ӵ� 땹�DO �剋_tky�Z%F���*���s��Ԥ�V��}v����5�c���K����{i.*����ٍvv����~��O���U}�����x��9��2�1����t�'5�Wu���uv�-�e0S�g���m�Ďov��rxf,����)���=�<g�����b�ۥ��`}�/M�x�S�e��l�y+ �Eq��6k���=5������+�c������Eq���O�#�=����xF��5О�wQ��������.,h�xn�}"�U�s�ꌻO��]��^Sh�����zn_,$Wmn��mV]��N���{Jk��]���.��e��0f��j�5t��UĴd	f%�:�w�!�����an���Czd*��!�2�=:��U)�,�U�6͋�9�k^�uN-v�T1�ݼc���4ܮWu}���j�4�}E���Q�֮������t�2��V��?�DkTv�h�~�Y���,�8+� ^��uz���{
	X��5�s����9����z<z�㗆�1]�����<*[��-�Y�p��>��n5�l��t�kc�g�j�f7]OX�US�}`��w��Ix�	�u���~�9.��o�w�>�qW�d�|���b�
���w�=��F�/WX+������U�:�Zz[Ly_dd�%Q��d��ر������ڋ�[�a<�
�e�-�73���;^mVf:w��^�8��n�o�$����ľɯX�hVYӺ��VEٛw|�r���<֨�v�)`:+�[�6*_Q�Q�p�NuS$��~��d�+�v��P�Yh���6�.����w%�Q����a �0�v�S���mv����aR�{V9���]ԇ�����+h����fr�&�V�Ì�ڛ�vd���P�BD�y���l=ܔ"��:�A����L�͓��Lc3�
M�����t���:��z�t�{)��u�9��w[|9[��ҕ��=��c�	��b��{奊�y�̕����j�r���S֌�����v�д���7:�T�z���PJ�ٷ9�u���<�:���-qKk�͕(Ca��t@)gcݣ�N�	�=:��\F�*Vt��t�A�1�&Ρ:�M=o��d��9fN��)ǭs�ܙS��v�vkv���=K0�js(u�'Z���y�����Oaj���Ζ'��;#n�ɧێ��S]��C�hAH
Jbv�v=�#Y��y򝧘�&C��\w;U�����Z�F��v�P��g�]��bf��-�ɳ%ݰV���+��`����!�׈=��2|�7;by�1���es�睷��"9�΂RC�o����m���T!>��by[ۗn�=�r�1��g\eO�9QkܸdU��Z}8We^�n��V���T-l�Ʀ'4ei�B�7q
h5�r��q>Z�qN'n{:�kg��	��w�ܳ1�m���P���m�t3�YSeؘຼ�؝�T˥4+��*.�d�����K�s�E0��b@LАՖj9��L�=Ok����n�ϯ5l}?	K(D�ٷou�t�=��a�QXѱDl�v9�1�6��*[:P��/:*���л� ��t�$(���-��y2�����U��W�rT���'�}*�/�د�T���z�9r=�w��C͋&q��UbIԇ!��v�zt�4>b��c:��;nv�
ɦ$qӊ�K��nW	L�W�ޡ���a׻���le���e	x�Ƭ1 bs�Oz���%��ǔ�3|)f75���������RzNb����d�	��, Gkx6mN\:47��[�Z����[Kr�Cxr����Aip�fx��^7���9��0/�ss����s���^YN&G���)n�ú������Ue����q����OL��W��P������t��Ž����_w�!CO�mwQv�x���.)��Y�-Lh�~�ɺ$�9�Ŏ�]=䃴�q��I�>��/�ڻ����m��6��nDF��E�j�X��<�Y���SV�{|'g�$r�߁ۅ^�T��ѷ&
B�)��n@�v�N�C�w��S�,enr��4ٰ6g�V`H>�W�յY;�Q�Q�m���a���سzj%���S�V˥�]���%Y����N�$3�.��$�.��Δ)�ۥ�z��ｽGFf�sVS^���/C�����S4)5a20���������娏�g+���[��S������q���\�Wg��u � ���J����J�B�+���iP�S!�+��#z���h�m"d���[}lu,���[uo]��rH^3HTx;iܲ�xR邳���3�w	Tq�VR��ho(e���&Ƅ{�bMs�SZ�\�Z�us�wFc+�y�^1�M�P�*(z��r��2���U�WWvY]�ၹ��ж�T�s��[���y#��k2̹�����sp/H{q>�&�7�3B����Ҳ�zS�}�^i��v�����`��c�v�
�V��^̹��k9�j��IS���<�o���4�G�ܲ��,K��=N3/ ��hb���Z��;�����{uo0:1��Fh}?|�D������u�~�����kg��=�����J������g�t��f%�*��&6�}:r�[��^*{�g��ի�lũ�t5�+ە�^��O;%����9��dX\os�_�y��z��>��{������Ca[�`'�M_h�k��f���h��\GtS�~I_��!P���"��F1ʶ�n��}���p8;��úU����������xMe��^z�eL���K��o�d�>B�qBƞNv��B��TbQ�Tjw��`���:{9�W'oyu�oa���u��~þ����N���J{N#���CF/T���=�؍tC��ˉT���&��	��Yo�NŸ뛻]��N�����L{:�}���mgvU�~�R��@l-�*���2�;��9I;o�ӏ]��xc�x�'-��Aa	Q���_�Cz����]�1.��@�)tߟ9�b��[	�Xo8��S���kn�t�Y���7��HS�Ǻ���\uAZ��졁9��^��g�Lɾ2���I�`��D��k��P���1 ��cn$J��2�J��_\ռ�ށst��E�h;x�g5�v���b[v(T�Tg��	��}�X���E�VEf�X�����8�M�5@k��)Y�<�5�c?�݃@��EB�w�-���0��r��=�&#459M�p�g����Oy���S����|((���.�n.�+��?���@�S�ڮe|�zf���o��S���ɽ�'3�Z��̍c���\.� uH�� �++�S�J��R95��]G�I�ڤ��g;~&�T���Ԫ̬(����g�pɊ%�@̢�clw^��Pg���Z�彡ֵ����diu�mU�����ge 8����xyG&����HY�M�v��]�cz�]��;�c�����n��|��v:�����p �K���<}��5ӱ��ZAB��#1��{'ds�:sfq��ݶGJ����u���z����]�kU��S���������:�f4���\����wpƲ�A�����Ć!@t5}y�	]w .��uf.��(�P�q��X�(�81�A_wNv)��M�N@��&Q/"3M�Y����T�Ʌͨj�y�yDXivV�R�5d��|�O�!X�Jٮ�w������A7����vr"t�,�5�7**����n|V�c!������TE5K��\�%5�b���^�r�Ue?I�1�g�(��4�����VZ�N�qp�]|����VM�|ʧH,�4��i���6�u�ԸзnԢ���P\	�!��@���+Kk�P��$ �����쵘���0��(���uN4�Wס�\�W�]a����[6����+[��ύ��c��y���]�4XT�7a+}��&��v���.��V�j"�p�!ƗW�bu`�C��be��n��Î�Ō"ձ0��@Fص3R|�95��":O>�Wf*�B�q�r�Px�" ��yO/��[�e�iO��6q�Nл�cm�C���9L�U�0���.�v,|B�O$rb��VfS�AT���V������5v���M�80��(KۊJˬ`���%�ׇ���� ��K]�p��2QL|rژ �7)�]��ɀ�T2]Ы�/Yz��V�f�A�IQ�?F�m��<�t��:;�e'�mժeI2U��bT)u���[��*���l�B�`�q[b�he/��ԊPWBed?�S�N��&�F��e��M�l��45Kt$���NwfJ��n�����$�L�S�@W�eMé7Q������ �̷�tB뺌B�q�k`7A��SW<Ѧc� ���%1f"�p��r�<�t�8��b���ފ�Wz�)��jc6̗t�J������/�A�lԴr�K�ǸeK��7���	�iح5x����n�ъŶ�3�o*��¢���h�@U��PDTAb�(�"����bȱA�D�+l��+$X"(�X����1��Qb���"�A*UDX���DcUF(,U��1X�b#*�,QQR
����Qb1`��1Um�#"1,Q�DTQ��������"�2*
�F"��(�����*Ŋ(�Ŋ
E�`���R�UX��`��(�E�PEUTFbU1�������0X�TQE�V �R1�b��9B����E1��dD`�EQb)�TDV**�0QUG~~�[��v�r�Q��:�R79P� �ڳ]pe���t4��)�Qj��g<�}ܧ5������[{�N4V���F�V��u+��O�啌�_+i����#�+�ܩM�H�����q��9�/�p�������E�!^�m�{i�ݐ���ə'<�s�ҵ���vY�K���)�ǩ�~~����rH���ݽ�귨]��|��+�iqYw������5j��U�o$�(d�[׳���W�����}��}��f�)���!ٴe�N��sg��7x�氼����t�����y�cB
�RW�u�\�"���\�^�uU�����窷O,cu�ccy�
�a��W)��/����w4���r���'�z���<��-�A�w��Y�G���1�G#]��b�oo0]F�<!����+[]�D'݂���Y����u�Ld��,q�Ӛ^J�p�#D Oza���#�io���n��:���Ͷ�\��t�"Jp�V�uG݂�޶�69�kvr̃n��.�:qC��Vb�!w՝���<�O	�,�M=RuĲn��T��|�#k^Vv6\}@��b5]dZZu���;[�����YӖd�]�k]Zn�w,�{3���:qn��Kzj�=��.���2���J��A�#�A�е�dc9S&f�ma�yz6�cB#����UiX*ۋ�b|۸�%빁b�K��mJ=�#'c]�=���p�)t����
礬��w�[�W	lП5njuW�/+���u�*+���c{'���5䎒�bL=p���m{zzX��g>��`�V��<����Hq򏕌�]쩻��<]��`8�.܋y�)fj]}|�ǹ���=%�y�ᘢ���r��{d��ƒ�ˇC��Y�t��*u�\�f��Ó�pb�q�,��\���4Q����<��I�����h�)�����v��	Wk�{>��nM���8\�]�p�]C�{Qα�t/eׯP�t�{8��	�m���,��Tom9�����vcn�of\�]�\�\����:qsy�v�noh)��qw0�x��r�+gZԵq��hV�e���+�n�3��G�Wr�­L�]�>qYDT[:�S�ܻ�>��w�"�YZr��Rr��z�v�5��lզJ�65��#�n��7]t@��5P��j��q����������{>�wx�jë{yt�UsvT�)+�M�C�'��.v5X��<�w��˾�Q��nO#q1������*���Ո����m�׵��؝�yS3��՛�c���[��psM��^]�C��F��Ԅrh��ܖLKW�}s͞���km��m!����ĺ\)߼���
���=O�X�:�Rl���u���u�s���]CuL,{m�~��t�
r�-�y�s���m�����2���n�5�.uv_�졁>�z-�c�[=a�zM.�գ���.A[q>��4'��s����U��i�{���&o�g$������l��e\����[�5d���|�:��4�f�]�[B�F&2�Fk.m����@T���J��.�'W�M�+�2̓c�=�6]��S6���~��ܟ�����q^z���t3<r���ɊA]vd�\	\S�j�s������˱�l�a*\��1\�|Yspo���t�L;�pq�ynmk�
������8Z����)ّk�գ��'�*�Yi���b.ׂ��;I�+��C}�!�>mL�����`�lܽl�{���{�Si�J�qX��"k��vq���t;g��;a�Ć��z����DWko�f^;Z�T�0'�����bލB:P���Wm.[!���q�t��u��Y�i��9V�g�L]\���ԩ�/<Uޑd��A�hS�@	n��=X�<����`{�q0���
��dW���Nu+��S�����]7&��9���o'�)��7x�r�U�z�mQ���Ƶ~��e�8b��tT.{��ۄ?|��mT�zEJ�ה�e��	�%p
PU�nA�'c�3��k�0R����v�]�ǩ�Bwj�� �/؃ݶި��b{%gj�/�:W�]���O�-WE^����-uKơ�ۮ̫c���<��,Eiޘ�<w�z)����|���t��=�گB}��*�0Tz��[�}���V$�f���;^�8�0AXՕ�X�;uT-lfў}΁UuѹIh�fH���>�����޻�$U���II&�Y�:�ػ)C@���V[^Iv{���oE�_v�^���Zz3.��3�e����V���M5Z6���]C���6GJ����jo9��8��vٍne�ju��IQH���1�m���3��$1�T��4V@�Q��[�fS���[�*Ҟ��Z��{�T��iR����8˴��X�݊��r�:�|Z9�z,P �<�5�|�B�ֶ�h��2��B�d���$����2/��q�b����g_Dc���_�{��s����x��#�a�Ll�7��������+`���Ǎ^]M�[������H�#e��T˝�7�!�[	�v����K�ϟ��۞�|uI��9����u��1=��z���v�,�Ȩ��o�ǧ��6d�Nk'���ú��x�*���i�XB����0.w�7������LP�v�~ﻫ�_M�_{р�"*��ɏ����E�>G'���#�������[�V���y�z�+��J�Ƙ�<&�9='���<�n�W���<�Qh7w�M��v����e�zϝOq�
�1"ݿce����[�%2]�t��(/�mK�!�l�[]��m���D��'C/�<�V�SEZUs2����%��O	��w��Q�����ܝ����a�U;he���[У{��PT����kl<뾲�t6-gU���٠��w*�(:[rWL�|��1�����z����DI�����'��=׭�^���HN(fʌ^��t�I��cw�5���,�I��e��V.�9r�t��)�Ƌ��C��XBT�Cd���$J�@[]��eb%�*gRV���zj�OgD���+s���K�8�]��[���O�.�<f7�F�Q�ޤ��s���'w�4�+OO�
'��B�v�T��1DuD+������oV�ݤ���avO�+�Z�ҰU�!؟��	z�ɱK�8Tҍ�驅��7ל�%T+���ɠ1=��_AV7�+�1=��W��D,�s+o<��v\�V���̼��{)c���+��ޯ<CYk�JZ���b��S��h�q����g�x7��Inr�|l:I���9eƮ��o+튊���Mb�2���ӓ�szm�Y9��O��}vo��䊜Q��s:)�9�)R�]�ޱ�6�zĺ*73��������Z�^��y�u̾M��=���I�[<)�-=�{�c�l�E��Y��'��UgY�� ;�p���<�Q'$u���r��u�����Su�y��)�y�wq�_�yL)�v{�jͶ�ܠ����\gL��U�t��NӍ���W����X�v��N��s�M���2�y	��~BX��7��l	�{u�1�U�}��\�Uv?���!���3s��[s�*noն�c�̠c^I�z�--=8���;O�<���Mo ���.���C�Z�*���'I֤�Ekz�F �A�lLm������V������gn9�J�	��P	4�ک��;�fa�d6�J��|�{ch��.�l����3���ԕ��8�o$E�4��w���W^+ȼ͓�O�iT�:�&��c�al�JK�5�r��� �Zyu3���������T�Ƕ�qW�e7Q
��Xr��I9s����>�B���YU��@���v�[Jʶz�x�;�Q��l��<�8h�v�E�k�[\��]7��޺�7�i�y�9������⟁]���9�Y,�r6�޺Ե�4n�@|�w��ᶅ�v���)���Y��L����AO���X�A�� ߂��qr����:n���J��*�s3��8m�u�c��� �ݰ7�&�F��b��T=}5B�a�/ywen�o)a�{�����/s9²%˦�~=bD0����mĉ[���
�ݎ�BPp8]$�2^��W��h�q�'[�T�r8>���ә"Sɰ��qse�|��i\󷲏5�*�5����7M���D��mО̅�D��oh��Z���y6ﱌ�b�ꮠ7�W/>������N>'���u��u1�=�K���';)���Pn7}���Kڿ=��7eW��K��s�1
z�u�kL��j����M�묜�cB:P���Wm.���;E��ˋ8�e�x����n|s�M�+�>��!����$t��y�{�6{�ј�S��>���ӏ���]���2�A�YҪ��a*�I�����o7c\�Ky�Ak��ѯ��{�z4b���S�k��{�3��C�����:M��ۗy҄�s1�y��kht�e��Bx�\��6��f`��ȉ��L)�Uҹ1t���$�1,d�,�pff�B�+$鱬���x�Z�ç��c��0uû��d��8���*1�$
���/t�G�Ϟ^�&h���\^�v�{Ji����J�ڢ}��b*Y��]�U�)�w
�䲗C����[�WI����sȼ������F����R�Hׇ��F��n�s���sG>�O8��c�c����;�u{}��F����N��S�� �j�]��U�d��'=�I=�z�V
oC��*T
|����E�V�YO1,{k9oe˵O���ٌ����k�aSp�X�7L�*p*8.�8�nǷ/v\b"�;����26�Nry,Z͡��zK�7�RL=�VjlmS驗����D�D!Q�^��]?	]�%���N'9�V�i1���Ѱ����3�޽��]�虗���;���̠��{�B=��lB���X~�n��9�!�����?e�h���p����W��(!(;wdR���QgEx*l�R�Z�ڳf^9�@�I�:w���njK����u�	:��8]D�U�@�oB�3wB����_2=�[ۋyn�tj��Ϯ���I]9��OEV�CAK@칫����k7Prb���;w9�B��]���f���K�����Qf���x>û`97'1P���ը[Յ�i�nUZZ�3�z��e��ضp?I�{����[�6׷�vb��'"��������֚�]���z��V�b��Ǎ�K%l��v��
V�3ksw����`[���C�t�`*�n�ܟ�^>{ٱ��z�m�<�LK����A�2m��7'X�|�\&�ڮq��ٯ{���8}y���ɛ$�i)o�v}�0�ѵ D$*{��]�q�s좕��M��%�o��Z��s���¥�%A���	\�kq�9{JӮ��ͺ��zr���J���1�N�T=v�B]p5T! �}#�)ճ�.`@�]٬�Ύ�:{7u��䓬��}D�!��7)��Yw
ӕ���e�W+�U�WJ��״�u�+eiV˲�O�w*\�J�pԻɃ/M`���Ţq�߇<���D2��mn�z� :�|�zA�]��c�l��9l-[�w�|�qe`ݼ5vj���/r;/>@陴�����B�2�2r	lЃ",�R�`�L@M�4�6�f__7K���Q���#��ݬ��R�\��>�2�I�t%���E�"���0�����{���tyR����w��2%,��Q����S���9�����J�M�_1y���4�*���g�;5��m֌P$.�A�_W7tz�1�M�j�޽�B�
�g��^ެ�O[�B�+4�q�4�>�i�F���x��o�|/��}7*��&�:8X�o�[�R�E�����3T�|;#Kg3�Z��@a�	.]��l������]����Pq�E��KXy��4r��Y[)S��R����^��4�g2�ɝњ7����Y�3��:R��΍fs7[R�?�	���Ɛ[�g�Z��E&�!E*��5{QnR����l(������~�S�FJ=�����!.M̐���OhB$�]�V��Т{�[A�]D��5̹z�m�nn���b퀫��5�@���4[J��[{���g2G�ec^�ma՝#�Du��ٽ��e��C�n�1 ��R�� a���/�bh:j�K�����ݗ�԰��b���yV���
�H��Ƿ̱[%^A�]dN=`阩S��J�阻��V�O
�1\%��,􊱜�)�d'٘�JŖ��N\�]!�y�R͎S����J�wr���x 9k��������ڶ�ޚCu�M�j��u��R��I�5建Y��
���B��m��#���v�
�i���ͺ��[��Jq�0�X3-6�/�J���JÝ���3tyqn��XhM�}Y���w�2�agw�T|r*J^�\ƭ���ļ�,�s��2��/s���+^X[����Rͫ�b��&���eҺ�J`(��MA`��t�� ��HC�Ț�n�YmCw	ե]�Ӱ�ͫ������!���s�W�����ëx`ѕүj7���QO'=���:n3x��;d"!�޺}Eaq��R4@�A|�mdR�&��bE��S�-����/�Kv@���y���[��A���N��h�Q�Up0t�
��Y�������P*�S�3�V� s����4��,����;��ԕ���C�]N�ۖ�����k ����C/[��|fv�A݀ŎF�e����&X���#i�lKw4�{�wČ��b��%�bvn���s	\�S�F ��go��p��/�6p��wcg]w�`�.;�9�\��ݛ�=WȚY,���5^�ZJ�g�ۤ��Sz�p);V򜐎���k��ݠD-���Q�ep�V��(�h���w��ѽӳC
��J��l�˴��,'�L\��5�%%;R��V��K/�>/1Ϸ.P�h5H!�sB��n�'��euMa�r�q�T*�a	��t�Wi�[�;y��.�λ�^�qc\�kЗ��w`��=lΆc�$��uB��E��i�R
�*(�風������E*�cUF"�E���(���őT��E��� �,E#��*�"�QDU(�
�"���F(���SQce�E���b��QU�EX�Q1TR*
��c��U��
(��E+QQTU���1QE�DDb���#���1��D���Tb�b,\h"���UU�V+TE��1��0Tq�������֊��E+AEE-�(ƣlX�QTX��
(I5G��ye;�H�[�훖��+a��'m���\��.��r)��KM��&�\n�WK:�geВ݋EN��w+誧mZV����uf�2g�����ĉ]���\IS��Hv�'Uo:�׷�ls��S���u9�B{�cO��} 6n��7+0���'r���;\l�f�UӁ���4�$8�.6"�Ep́�ձz\ގ>O˦vʝ�sj���|O]'��*�x�VN<p��:۪w�μ��3
{�/��
-��9����OW3���ř��tCn��Y����[2�UQ��6�F�P�v�#��J3[��\Vx]�<+M�X�8gw��Z�^��Ê��R��m��֡���7ڟ'���\r���^f�)��NO+�uY|�d)�ě�v�nd�*z��=�NN;��(n#�����Ym�uc�	WI�u�<���cU�%X�\^vj���7ݞ|���� �Bm��J
�mȈHP��Jo�h>^�v��!{#u�6�v�+����536���y@t,m�u�oKbwì�����m�a�޲��1j�n��#�.�f�j��J�1NM:��w���8��|�=��:�
��Zr�d_91�q��rѕ�"���k��s���n��}�M�w\kz�a��l-��p{��m9��� ���N���3a�9�Ak��o��5��!�-�	�T94�X�W�ejv�P���H[UN��\��]��,ĺ�i�Wv�/�f>�ҵk�o4��2}M�%��6EL��]
|X@��y
�זFUs�߯��]���t{A��fi�Cu�6=�ɚ���{�����Ӻ�`X���.���$��N7D{��X��WD<��V�5ki�OUݭ�jB�`q2�2R�H��x�ic���ׅ�
�L9[/�ح�Z��,�fv�P�9h���	8tK���."P)S��lQgF���T����Eʕ۾]�TE�s�O'�`���wa_tԸ	~��P3�7���A�B���T����ÝQc9>x�8�>5C/ν+v�T�J��N2D��G{���q�ZϹAſ#�
w�b��(*[^+:��Sf�,R\u��TI�oK�g<���D5�d2pZꉣ��S��^V�몖dT�����@�L�<�����{6�Pُ��_&��i�������!ZQb���y�[w�s�t��h����8a��u��9�k#����������s�B��0�X�<��՛hA|�ogpS=�����R+X'�Ջ�YϹ�)P�5Μn�u�<����U^J.�O('����"���es�ͻz��[�)�����S�����s>�t�,d>�2�3�j9�����dv�ڴ�˴���cu�{�dv��;�4�5t!#R��K<F��ё��Os�Ҟ�8*�w[8�����aC}�A�?8N��-�W�7ے+�A���׹�|�.�gzgc�o,p��'uȱ0�;Ua�AR;�g��ņ�AM;�P�^�s��!Z��7a����ۼ�`n�4G�@�qw��S�jp�{�3��:j��`���#��R�}1����)ص<�J�����e+ѲL��8��B!�ᠺ4�Qe!��2+P�X������KzX>�n���}M�p+ք��#�.@����,P�j�]��Q>8��p?O{���6�Oޝ��,��1�[yėQGED�}^}#���|eR�h7��c��S��70Zp�j�Y�h@��Č"F�	lʎ�<h���%	WN`���8��<:�%��f������<��+���݉~M��D,���c6���]�[�44�P�"�v:.͈n�{]s�q'�zI�ڨ����ӑ�N���gpǣ�;�t�u��"V�7j_=��8�Xsw����H7�b �S{�TL��6��:���F�����9�<�啗�"@�<�u��>0]�9����,q���[S��.����ڕ�{]�s�f�վ�n��3\�۱N�-̫S�&��t����ޱ.8;�MM�K.��3��W���B❝��ٍ�	�\���]g®�`8�� ���|WMܿ�5��F�"��ֻkC�d{ï&�ej��{���V�a6%x� ��[\b�YSL7hʘ��-�X��(�/���+�&�uk������im��La��d[�|a�Z���M�/RO�s�z�s��#��'#A�I���8���Z{��N{2O���^�0 t�&�<�/{��Ls�Sw�C(�����j�ߕPG�fF���dv�&�(+��5���!N�YԳn�_�Sou2�<��W��W�$�Kqi�q���i���)Z_y[�@�����2p��{lcN���B����O,��ƣ.#�Պ��и���~�"2F<�#2�\���ƭ<«�>INGT9�!J�H�0'D��7(#S Z�,]������T��hz(0�@i\Ҁ�Zi�4U��S��0�=�L�	��I��2�S�P��l��U���!#B��I�y�OQ4V�.,�����U���˾��wbGGptsm�G���6��O	wYǤ6�<�.h�"A��Փ�p�aI���s���2��ˆI��Uj�GdR6p�(�2�gd��+�iuT�P��+�5uge�Mu����C�j���=^9'x�S&�oț� 7���_+@W��M����GA+���.Z���n��� g��s2Y
��P��o���i�|������3��+l"�В���?u.]�0�{c�9C�q)ҍ-���86���0�˵��S۴���y �"�)��ag�eĐ�0���^�G6f��;|G�|=�y�����*0���ӷ9Ļ�@�Z�A�*�6�+�ub��<f|+��?��J*]$	eu��{wn-#|�Ę�y�D�=Xѫ%�Y1��G#Xاi�h���KX�ɟv�洟.�<�:_��}Hm���΍�,��wG����Y���:�;GgJ7X�O��_���ms���m�h�유�y�4`3�j���q�h'@����nǴ�°�+���<�Λ���Ji��WJ�H��'��k�%ۛ	M�m�����jr�fJۈ��o*LV�a=`�P}���(�.��9�z�o�Or���\U���5I-�'ǖ��v+c���9�2���+�������|���z����R̓x��@H�Z7ZWph�,=�����x&`����ճ��qԜ�0|�.���7G^V6m�I��\Y������x(��:�t�tD�_s8�bm�O�J��
��0tV+c��1)�R�K�1}��r>EY�*�*�j'�̑�o�;�O�=�쬤�[B���c0�x<�N�L��.�ԃ�ۉC&׍m
(�F��YT�-�" �:��HI�%gcg&q�ǌ��}ʮ���݊���U��S���UpuѾKُ����O���4��.���8iz��靎,Da���DB���GH�fN4W�=�q(�-^�Ǩ�Y�2��X��5�R\n�����͈�Qj	%*.�%9�]�ʚ�.'^R���
�̀��-���=X)����s��99z���"K�&�[�w{=u���6h��`�,�l�`D}"�G�Vd����*�R)���dz���:�x�q�K)��������K�5���#�$F��ɸ"��[:���~�0�hS�H������{'-��L����Ѩ���:K�U^~����z�D>��@��Qo��^��x7B��P��ZYu�^�R=.:!8&�xM��d
�*w$ߥQqâ�cǁ<-k6�<�<���wUh����O���O�/��~���0v�P�:�T���}���w5N�%��>��٧�F<����i���a��	-����SLT~UЭaW�Ho9%�Tpߜ�g�Hp�]N�1�E���;�V+����wb��)ׄt� ��ˮ����j\���>_,ύ�]F�} �֥r2>\f�U\�7���d?C��62���[`m2�&��@O��t;j�H�%T��$=�1��m�����w���^�Gn@o,�}#�[\�W�9�;)']��J�>��y��v��|7�u_m[�:��&�^��<�d��gl�*U�\�q�5�<ا�_ /�4<�{�.u���wnl��v7ר]��,s�z�k/�59�9�
6�W��c�F�Aꐬ����èN ����;Ζ/���$ᡯ�����dv����ǲ#�{P ��A�N��yÅ�W<9�T����}QO^�@�����s��D�#��k�p9��O�n�䲤����zk�*͖u$�� ����2{�R���XkPT��>gv�G)�a��\j�K7g�Kv�^�\�1�-!����b�&U5��T�\5���5��%tw�2���ͥQJ��6�_N@�V��c�2)nf*v�w�%j�{J^�ҫ�+�{�p���qz�Q�P�^��K{����s;'H�B{����d�œvޜre@[v���*�[�|3�7�e�NǸ�dw��.VkT��{���f��s��N�n���L��R��{fQ#d�q�:���a�l����w/lT�Tӎ7촕�U��1۵�\��.h��n\@�ZZ�ْyt�/`���(��r��R�'y{����tr���]Ƙ�n���<�2lz!KR\,0O8�OeI����Z���㔆�9����];>�	��QA�L�P���E�$�o,��q��ՙU���z�|M#:�$��x�vf��^�ļ�54�lVz��=s�HR5S��JX-F	s��4Ir:jK�噈��U��rרGs�!���`�٭X�����4�+Ջ��"*}��)z8;����	t8e�i���'���;t��vO�Eg;Sd�ۓM	��Fx�u}^�y,�� �y<������jg(1��b�ha4Cf���5����N:k6�{)̸AR�Y�Rޥ'Iț�X��F6�3�ە�2�5��ڎ��:�864�&��;e�wD�j�1N�tn]��U��A�����_B<�i�y���V��ʃ��֝0o.Wށ����la�
Ȯ��L:�beޓ���];!JvkoF�(�ܻ��c��u���>��\�H�����O6�i�)QSvm�`,I0VlM��'U�r�U���+��J��n�;:����dv�!go*Q�\\�����v�r�g9@�*D��϶tܭ�~���ˮ����Jo�As˞cʨ#��n��[#�+��]༱6�Ob��F�m�&bV,J��؍,�먐�O�k��lQU��n1�q�yCJ�xTԨ��f&orB���eٲ�)
�b��B��K4�+�x��}��Y���=���,��=:�t'���N���.ͥCj9��O�«�E�jt�0(�3Je�%Pʘ��5����hL���v,�s���C���s��{�Ӈ'�ոg#�������%�zQ�@#{ҏ�S��a���<(�RUP�O;�	�Q�gK�2h7T�/ӊ�%>�w	{����)[6��rU�ħ~c:R%��{�v�̖B��7�E`m��lil��9D9<r�c얚������C�e�1��2�Dlgl�>�Mxа��lX��=�]/+�{G�4L{t�_L�<Z�bxLdH�\2J�����B��+إ���QΉ�Y�T���V�5jZ�N�桝��bvl\�,��"*U4#���YC�N���Y��9��~��q����N�K,�R�5,`����!9�=��Y�ֲ~t+;���:Y*�ӝ�LsH���o����~�����zfc�w[�y�7m�R'�C�q�N_4+M���,��p�W'`n��9u��U�wl�������j`�J�U��q�G�|Ĉ�y)ƽ��J坽�W1���V�D�`B�]4j�5�*z*�SPz(��s "B�uѧ��*��D}���DD�k3 �Q%���SF�^o��Lfz0���*�߷s'��U��s:�b��O �W{|C�Gѓ��\]��: �+�m��,�N��wVM��%=�q6���;O&��ύT�UVx�TD�nl%4F���v)��<���	�����ӲA��#��~b��j�����5A8p����D�U%�����Ǟ�Ӗ�>���:Q�ʉ�`��g��0�u���%SK�ϝ���]!(�Yn����Җ��wϞ�s�o)��Q�/�:َ6�A(�(��&�տ
��]e�W�����G��B�p�Ӽ�� P�$<��9�s�坿%w�4aF��"�T�F�g�7xn���}*�w>�Ķ-RԶ��$�58��#�Z��w��ë�͈�Qj	%'A�F�S���j֫Jwd��L��GQ�ɲ�:�t�NR�5�#T^99ҥ���OD�#Y*�,yT�̲�6U�S�!]���xq�t�3��At*��K�q�R�]���pX��}m&r��(��J�9Iҩ6��Һ�N(���/��j.�����lҜ
ț��X�E��v��曊��Qufr�dv9��n�
Y����iu
YY��%����@���w=&�f[��R5��g>
�V>��%%u�>}�dDDX5�[�؋j�}� &̦��P;�s��m��ohb�6.�g*��9��*b�K���XҮ�[�r�P�Şn������b�*�S�M�9����_	�b�k,�eh�N�ϣ�8��\V��p�N٬��e9�A
g�ح����u�Q�ܨpmc�2Q��[ˬ�k�}K{����A�Af�3ݲ9�NC����{eǁ��F�Et ,5[���XU|����%P�a�[r�'��˦0P�!K����C*�VQQj6��Y�)��{�5��ϼ3;��{Kx�)[3�"	�[�������<����sU=VNL��Ԙ��$^��t�̎���*I^2���Ͷ@Θ�R�L��]9땽�kB�-�`��n��&EtN�㮖����9�¹���:�����@�z�p�7\K��@r�S���uM���Ոn���1;lr��kf]�����}²�+��V�z�q���1�rĭ81E��3WV�F������ ܄%x�J���dSj�x^_e>�\m���'�VPy���k9�K���P�8[��T��87\:j�� \�n,�+�M�Y/��#b�O�1jX���Pr.�];B�b��ԁ��ì��:LH+Ȣ.��qVY��i���A1S�ĢFY#����4)�Y@b��*�`9>B9t$�(
[uy�%�ـ��C�R;8>U�Q�� ��e��b�B�
�݂�$��/���1R<4�8Xv�JW@Q� �)��6!P[,F�xn�"���(1vR�$�1�YXٰR�
"��6���pGI�ER��4�ZT�`��h��n:[�dy#��XO����E�V�L�K��J9,���˳��;iX���1Oe]X80��䴤"��F�- LthHjPwK99�+��%�
��	i�#Q
r0œy@���q%�+&HS�Q�l����d�ȣ+�H؊�+qʵ�a�Z����aXp3��.ݽ�Y�nE��~`�ճ�s�)u7h1-[ل*tS�"�80�V������A"�Xl0�;1�a��9-;�d�'�@�l���ڱwm j��r�!+y��� S0��A��^d�J�+6ُ�vh��ڨ����/�孲� �*�i�p�Pѭ{*�L� N��jp���%᥮�eYL�2�y�b�!�h�c)�����y!*��E$pҰ��!����Vc	���*=�ɭ�2�YX�A��\kdt!������*���0T١��`�V�9ĕ�ZM�Z>���QCƋ������[[Z�+Q����V%��U2ʢ������1DJ�4�k�QQ1�IU��(��X1Q*��%�Q�UX*T��n5���F��ȩi`�h҅Q���J(�2��*��Z�)lUaR�UeQ��*Q-�KZR�U�S)RؔDU�*���Z���ګm�pe-(ڥ����ZZ�2�YD(մm��(�E(Ѫ�kUAE���V�֬V�U+KF�JVYj�PD[ZV%k-������*��
��U�EjT�,�KQ*�Ѷ�0�1(5����iem��*�U��Tk-�]?�<}������6ԓ�N�>��n�r��5A�e��@�'w�������R�"�S[�X��2�Ӝ#n�Ww���\7/�1y/���*�3��40s��Hk�X#�7!��]\U�T�p�=�u�69�!Z��s���{��eĩ���B�-qDP�^�I��s�5�ʵfE�f:�t���u��f���4v#�N�'�IJ>o�P�{�<��(�Z�i��H��N6���!�Sۏ/�qq���6܍#�{V�L��`�%���*w$ܦ<vPt����sc�R������W�6�L1�F�{6�lX���5��I:%�B�8Y5�RR,L�=����"��p�׼[᷽f�]1�����X�ص������e�?���5��3㹓�s��Ͼ�2�2~Xs�v��H�~ɡ�.6C5;9��4�d��%l�����fqH����Of�Z��u��x�S��]#j�:��j��CJ7n�U\ºU
˜��j�3�Xw�+�+�<���h�q+g�{6�gr�/�SJu��5a�>�<E�+�J��n7f��R��Cnh؋8�J�A+�����z��kn
6.��K�`��kUu.�(oy�&�w:ù�W;�i�'C1��C��(��sFC۪�h_���n=��Y��Bw�?%}���oD�=����������Q�˙s���Y���;�&�86�·��@-����ENB��U���΀�Q)%��;���Y��7wc3l�f� ��͆P!O�L�kv�7�%�ێ�n�#��*:,-�V&ʮu�����o�T�&��`pT���di|�:$��[��8��т�F��$g��n��x�T���Fڽ������T������;���
���ݏ3�	�"e^d��:�K���S֌�mg��\e}�\��W��؀?���9�>��g�s��rVOnYq��/:s<�,v�sS�2;��"�EK�^XiwV�P�G
�[��<+���h2�M]Ejgs;X�K�y�24�cgJQi�q���ι���7. P�$�6̓ˠ�'�Ѫ�L��Cqi�ܲ/��!�0�v�V�~��Ȱ]Ƙ�ޓV��I�s��.q$�T�c��3�u�y�+}}z˨�q��V�X'��D�fC��26�G�-��zU�"=���O�Uc���={��q�,�$+�NnR��B\�"�'��E���䰵:l�W~�Q׃ڨ���Pڐ�Ve��K;Q�0���E�
����{��ט����{b��܇V-��E[�ڵ��Mw�S�]g��f^ҥԢ�uon�b�r��7#N�ܣ���ȳJ��LVeR�b�Q[����ǯuw݁�eaj�hܣ��gE���&������ݷټ��z
�uuF��:3�����e�4]�����n�Ϋ[�&�
���A�Yu�J`�n�양Y�Փ�nM4'{v�'U�����\:�ow-�/�UI�v��s�H[�t�lOpEhTn��C^�\�0,*���4��s�\��ل�Ɠ�.	�o*��W�[k��W�������:�9GgO�f.���y�W�kjU��#O+�#��W�5��2B<�kv8��)���9�ۂ�վ�@-�s�x�U�ٙ&��J�7�U�Y�E�'����|�2��ِ��퐹B�&�ӣ���{�k��N�f��8Lt٘s�!s'��B�*�P-�c����k�q��굂�y�i��Tx�O.D����JI,��ﷸ,Oj��9��7��^&6��Ib�K<
��	�<���<l�)�B���@����&$"MxOO8V�Rj��֥nk�����v� lQbc:aWg!,�8r|��,��Ȥl��C��0����^��y�:<���aڶ*F����}H[�N�a�*4��I�Eҙ4�L߱	%U
s9�́{K�ȗ�f��ݜ�Y���~����o�[[�mv�@b�(f���b�T������8tK��Ҩ����SX�sh��@�K��m
��|Nu���OT�����wal��v�*��1[=r���edy���\�b�"���F�]-Weق�	���
Sy���{r���+u7$�{{�N�/T�����Z�����t�_s�EЊ����u�oyZŘ�\�$�E�wEa�Ѷ6t�hNd�7q�tV��Ɩ������b|bw�'k���m�M&"=v��X�|��z�%N�� �=�~���pE(Ҏ��~�`
fX�\�y�Ny����MJQ�: :: ��^[r�tX�%�b�_/�<&}��֒���g�2m����n��D�	�(a�߽���Z��<�k�U5T���R�mG��&N9����I]5�>�*1�,����e�޲֗<߸�:��f��0��k�9�sw�q�D�P2�1�>N$tQf�mT���K3�ԟkF�M򛉌6c>�k���^�s�n{~��]��Æ�8��l dˀ��f���/�F\�nA�j�k��[7���vj�؈��"<�ю���Qy����{��m�b$�sa9�4�����T�En98�%�y�)��!�"7c˩��l(������r�y2p΅Z��|!���54y�,66����Mu�C4��5����5vA�^ǎ��Y�R���"u��,[�NdK�.v��W�b{�r4�U��F������z�Ĥ�'�B�ْ�j1"�f�&��`�-5j���[�uf�����H��w9�8����7�7\����	���`-�J4)]I�`���9���6����@���<_`�yP�����5훪9�DN���XOȰR�Z���(���VdpY��;|:dt��4�3j����7�#M{�Q����P�7s����>����t��a�F�%r.�%_�@�AB&��5yXWE�N�^��(�rH���ol����7�sZ���^��M�U�H{��Ҁ�a:8�&�9�!qC2Y���_�25�,�Wa����Jڷ6�U����,�Ċo,)OS:jW��*Z:,v�g�z�&�B"����b԰���9�Noj��޳�*#��i��6)�0�QJl9TE:�2]����l��̿l���x$nP��F}�j�d'D�.Y�z ��g&߇���>}�Vl%�<��Y�5�3����f<ΌE�gr^@�,M�U�Q�tN��UG&��jC�"�����u�]m��k�-�<��8�w���f��y�y_!�	��Rc^2����`�7�p�V$��P��VD��A��CXr�P;F:���1�VU�^�S��I��n�C����<��a9��8�4�r�]��p_q�}�)��g0�y���R�������\��KH�*k.�WjB^Rc��Sm5ܓ���oX��4�M�S�@�]����ʝ���V}T,W�����>8�4'r���3����� G�i�x��Uj��y3���5��uPЅo4x�{Q&�:��])�𮉻��q�J��u}��S��H�����w7�{+ݳ�,�c��d: ���Jq�5�<�11����3�,x{_�n��e��fN0;+�ar�Ԏ<q�V��V�"2�c���1�#���Y5��wmm�fy�)ɹ�q-E�O�gV�{K#���udaO��Z�$��Z�Ȍ;�i��{���%���2���6���M��/Hx������\6�j�l�c� �Ģ��=z��be���;
iU�VfGS�JQ�_}\:�Y��������Z�[�q�㸘��Me���eK�[*`A�Q+d�4R�1��6G^�p� �0��&+$�{��N&��ڱw�[x��T����2|�2+"�H��JQ�r��6K��g>:���l<6��ת����e�ya[�V��<|�8���$�;O.�	b3��	�D��Pr�{��	ŶB�txz� ��p�M��m���u3Κ��շ��zXy7	�x�y��9��V�ŋK���k��r�T���������G0M�t�\�e�����gA��]p��s�z���f�㔔��$���ֵd�=Z����� r�݀�Һ���~n���O"M�Nz�20p���q+�
E�����T����rܼs�V9�#5���(�D.�p#"�0}`/�����ͧi�fh�ΖSDy*��ӳ��[A����d|3����P�oS�����/v�*���\FR٩֗S͡� _��u�TO���[�b�R���倧X�{�"�{���;¸���;>~���|��{��{��?��'�'�0:��b#Ht#NdIY�qf&�`�K���R��o��AwvW��ܱA�1�������8m�g�X�#����`*��փs��V��ƝP�5@��d����q�j�ӯr�'G6�3����f�G�QVd�b�v&�����>r���=:@㭠���IӋ��n�5��X{��l�8>��ܰ����`�W�	Yf�H��'���Ȓ����*d#mϒ;�-�w%���=�$n��F��<��2��*+^Nx�Ć�p״��H��qn�
��G[���\�㳳���b��u:}�����y���2�GyX��tV��5<�:Q��Nb��7��ޫ�<պ{*Ȳ�6v�
�+J�U܎�.��U�Y�A3�)�[�����	뒨Ҝp��|�p��ؤ�r�9����+�{���iwsĉ�����c�ny�j�c��)�L_�R���H�=�tO���3�G�z����6�t��޼�:�:�x�V��t�X
����M��3~�U ��>�%���:[IVYʶɛ�ˑ��,�^�q�K;��M���Ўؤl>��D��Cʊڎ�n��]�����`iZ�H��Nfx�8:���ǟ$;�y�ܞ��$���WI���ح�$ͩ}~0�m���3Bwh+�A��C�؎�݃�������Ɇ�W�T� ұ��n�>u{�c͖�(}�w�XǓܞP�8�s�p�a�uj�(����x��;�=*p�r��~L����-�^�j����_��d��w�3��N��0	���8��>{��h6n������9�ݐ���R�mE���jɬs�'r��6�=�F}g������u���x��{�>5d��&z)̾�6EU�$-��A���l����^�YQ�LW��Hn'��5�U*,(��Ն�ϫ����UVv��i�{%ԓ�ɢNķ�,L�3Hd@)od��ICc#v*�G95u��כ6��ٚZܻ񵔟Z�kwz�o��y�Z�� ���W[O��ܮkOU��у�9ر�CZJ�8(ם��Wj�ìJ wD�3��v�X�m��w:��Ί��8��{ϑS�r��U�]F5��ٽ���.�ݛ^�_���r�'�5��K��|�����D��rDhf��;o��o>�U~9����A|P��M4�7��8Z�n��ǵ}�r�8�X�U���^nr#v/�/㔫��Y���3�a��L=;;p) �Y�Jr�2rݣ��]�c%ߛ&w��s�>a>�ז����P��<Շk]z<t�	T�� /?y��B0�S$p�u�ϴ
R�3�G�&��791�dx��YJ�]�i�;q�׸�#��];���؅>�^!�c�q��gmU_B8�[2� �"�*X�9[�rt�<Ĳ�
p��"g���Sܦ�D���7B��P�~��e�wzBȗ]A��݉,N����o��FOC �y�T�*�&@�\�ES�ٲ�N��Β�\�5D�ʨ��X��]����Vc�]t6� �zP2pk�[Q5�iЭ��=����8�궖�a��q�;��3�p'��'�Q�j��Ψ]
SJ`7����\�d�xT"E���uӤ�8R��
1f�����Y��Hj�8X��,u�(����2�ڳ�5t�yu��\����'�j����PP�q������/��u�F��ǒ�9�wl�;�*��f�1��8�8u��%պc���vL�v�=i�b��X�L��c�����k��`�;�UK�Η.o�P�X�S˙���M�+��F�Og3�����_�Fމ "�[V�!:%�z$Y-s� h�t"�����l���4W�oR�{��ܩF�:fMT3���s[AdP言���QI�/xB�8l87���L$�cn�(RL�W�g�֍�6�;��0p�_UP]�2����:{����	�S{��]��H�����.�DQ�J��Q�^M���XJǣħX��/:���q�u��Z�t͚��m���j)���;�N+� ky�Hb�YNK!p��7��A8�&Y涝�ZԮM�Kz�Β��c��GCꦡhk�MJ9d���a�,W�����]�Ƣ����1o��zeuJ��v���_o�+�aT�{#Om��Pk�8��0�۪�Fە��LMdSk6�v��SDi`��c�4VJ+Z��J垺�۴��*����h��Y�~�s`�Xar_�L�D�3Ԑ�ΑΆx�$�_)Ί3�8���8��=���{On�J#h��A6��&NuԸ�gmm]w%��}˵��r�Q#�+,�YaF��ڨ�':Gl�;[� =r��Li���^b�-�.X�G�M�o]&'gg4]�,�!�W���Ov�km�Ō^�Ư�,����xKh�F<��C���̛��q7CZ����9.=�l�o.F�ts��n��"������,SסѬ��-i��md��Ծ�qnnѤoQи(p�`7 �s�ˡ9���`��a��S�Aa�,f�;�7z��{p������}B �p䆳�9RPp��Ne��Ev��᫦��v`�n�ف�� �H"N:ӝ�۽��6Z����59]�v1�ʸ7j]gs#�(���+1.�z�2WvM�;�뎹���� �i�w�t�n�ybwf��V쨣��.8�5���JE��K9`��)F�[g��D�ĬeG�Y+�r�S�!��c�;q�- w�y#�t�vb'#ɵ�c�E����v�oQ�W=�N1��V鸒�����'f$��#�i|��Ub�gUi����B����")4��+�*�ź%&��Hٱ|Ɂ��]��Ecu�]�7���ř�C]��H6�xk{�BN�6��)�Ax�����fr������[t��5m�D�(��`덗�t�Z鄷S�d�U�M(�5�u1Q+:������j��S�뫫��6{�SKC���+x6+�G�\yӐ���wYo;\VYs���۴o�����H9�����J7�b�,�'!5Z��:�t@�S	Q���5wv٦څlD��
VP�.�ʙJ�Jj���e4B ���hk�iն��a|��w�*6Ȅ\��S�x�� Y�x�����I�5cܴ�C#f`����X�w%�.���2�%ڥUp]�]��PAO�����'1PdYh�XI��?b�q}fÅ"�U�99�%b��T����S��1j,���YQ�&!��#F�*�|D�����fd�.��e
x�̙P�V BRD(�i8׋��������^y�`sd�I)���Ɯ����a�:K)�F�2�c�WN���n�I�0��]=�kX�X�jʺ;p���z.�
7��@̕
��F���S0n
62��9l,#��3�1X�
�&$��j��f$Ƶ����Ō���ʵ!�Y&�˰U�A�v�\4N�"Iv=����c^���(�HmkӶ�-R���L�1��t50n������óv\��dbdD���K�)eد�j̶NABHj»xCT5� 㷙�jU趕�%�������Ӷ WB���O:̽R�����\�r�d���Ҫ�ҫ�be����-����ʂ�UQ*X�ƭ��A,@��E�[j%�����ڊ�e*aV�jR�6ڨRֶ�*VZ�h؉V�-���J���+X�TR�-A�+Ҳ��"VV�RҖ�U�Rխe`����Z�j�����*ZV��T�RҪ�jQ��*�mX�KIDkr� �UR���*X�ҕ��KF�Ib�eJ%EKBҬ��ek-�[*D��Eb���s-V
�Q��-*4aV�Q��[kR(��AAaQ��+FV*�"Ȱ�RҖ�[V�(���#J+lR����Tm�J����5�-Z�2�EKj�Q���Q-���im��ԭ���UkF�T[R�ʔkA����%-EV"�,AE�T��,Pkc[��-+ZR�m�X��YbZ�-�ZQV����,�����Z�{��|��7��ƥj����oT�r���;k]a�	c��{��ga���rf�έ4,ɘ��ٕ���L������Ѫܮ;�l�>��uc.�B��\{E�u���Ն����za�#`�J��^�#r�yD�v6v�ȵzQ���:�T,�F����0K��G��'p�l23W, �]�i��[�4`���G����l���!ｱט���Pɔ��e���4:��.w�6)j�^}Q�s�Au�i�JP�q�aU�%U�>����V�-E��<����
�_e>���ʷ]��"8�E��]�p���
Į�E��4�XޓB�<�2`�����#8��S�yڲ��Nı[�{�MS�Ӹ��P$"$k2[v�G@�(*��\�Z�mW(����>Lg��)*�k��ϼ%,����\�H����!N�9��c5���.��{J�P��wa���h�D��a�TĆF08D(ys鉠6���U���z�6,�)ٜ����Avȅ��9:�w�nex�{�<K�'Hz#NdUB�dl�L%����ى��͚P����(-��6�uGj�j�#�L���INb��e?5��o���52�\c�ǆ�\��3z�TN�U�:Vi[��c�:�VH���tӝPv�P9��=F˃���>����q�^Wvr�+.��::o
��A���Y�G>�jbQ��#T�H���wN+\�z�9jx�Q�+�E',Ώ�le��:g"�@�(��M('y�8��W�My��^���
[�G3��ܺ��{��r9گ20nY�M��T����ǲ9�(�^�H�]#����$F��FM�˼G8��]z�Z/�}�Zt�OR6+j�����'��Ax��t*��8��n1v���7����:*��p靛әB�X�X%4�Ǯ$G��^̕���q�r{��}o=���Z_nOp�sܲ��hԺ�@i�5|h�If�%?-㣁��W��g��ֵt�[�]��{�>����W�q�S�z�]�/�񲈦�C��3 ����L��j�}��Z]՜��Ir�(Y�����5\E��wa�m���n#����cD^c/LU�r�a����.[�ڤ�p�1��7R4�rum�Bu�{�{�i�*���ǟ$%��vZ{�ܲ�T0��x�@�d�6�\j�a ��ׯq��9�^�#�XW��0��w�VNu�1�C�0h}t�	��vegݴ8��;�Uc�;4�u���tZ	e����A�޸&�~������-�Q��#��J�_W"\�Fk��kJ�X+�5.�;�ںR���[LxAf��S��u�C;U��{1�OU���r�Be>�3Cr�]K�Es�9���T�9N;gp+�μ7@uӲ_2�!KǥN��I�\�Լ0����ۜ��8����|	��)�jǙȅmh]�]�b�׭��������)۽�E�=%��m剷�������u�j��A�b�q�:�ϥՙ|�fOK�w�Z���R�g!ϞŉSd�w"�U�d��	��
�e"�lX;Z��1X�O'5��𮳃�z�<���������>g�px u�^�+���+�U�r�k����yڪe�Od��ؿl�@HN8�g�fTpQ%���O�5�cx�]&�_!�1�6��Y������"j�B.6����y�t9M_L�Hs�W����_ K׌�6QG1�PSg�Y�I��"83v�Jv����� c���kڨ
�����͆l]�{89M����b����s����2�\a;=tH�|��+0.���iI��jvϡ=���7}��k�m��{�tT���'��+����Y�k�G����ETp�q}z^m[_f���[Ω"oss��){��#�&8�7[1���I�
��EuĽo�=%����c>��P;��Oǟ{)d
�F8��gg��������c��O�g��;�+���vuOp������0_]����%��.�D�}���@{���5�W!�f�juȮr�z�]�w���W��r��
"1�G�H�"g��.R��Ȓ4���V �q��V\wt��T���WG�G�ܹD��{ķX=Gn�C$��H��L� ҄M
�P�mAJ4�ru��λK��w��[�U٨^.��IȡnՅ��I�q�1W�I�9�!q��������z���}�~��ʉR�<���&�ٔ�qN�����P�Q*``k���<Tb��3½e��yat���.���m�%�4��E���4�؛�T�A�<)p5�˺����p����/{�y�x�˫��,�����!�Hd3>�j0Btvɖ��.\�-�q��O�T]�=�oz��A���.vtɓ��,���E�!P��t0�^2x�NM��D�����W��k�I�j��Tih�1A�<ǀ�Y����X��ײJ�[���m�
s]N���Y��ǁ~��o�8�2�߹�n}J��Q�^�����X�X���&��	��R~Ӽ��9�һ7U�g%3�hUQձ�;�";@�<hiF��GoºSV�u��<�s^�οK4Q�P{Gb^�꘎��"N��K���3��#�2�+WA��g��?	<`�UǷ�Y�b��paH�T��7����}x��.���w�l	+x-8+��]V�]H]���3	MS���gQ���[Ց�n�;��y����P�����(��f³��#��ݳ	_���3���\)/v,��x�Ww&��J�S]�k�Iy�N;ڒ�vW(&©�F�_����輄Eh"���x��I&�9�U>�ژْ��u{�!8�C�����
��QFǗ{|��κ�WM��*��
\7�A:�I�6j9��G8]\���HƩ��=�3�8���v<�wK�uҽ��T���i�MA�E�]f�J�$�)��fx���JE�)C�5VE&�y]1����H!�b[𮴇xuց�J���R���T��Z�V�;D���sS�9��Ԉ�)J�r�$ѳǟ:j��J�� cr�{��n�X皪r7C�Q6�mwޞ�͗�^v^��Il��GT0"4��fP}3�-�Y�	�������*bKS�o.Nv_%zt;��*�7i��]�L����=�u2�����
Į�E��4�Xn����P\�&�[3���73�H��U�]���0��&�
]Zt���!��x*s'����%�O��WV��,��w�cyFa��	�YB�K%�	�-(�TO�f)��̾
 gN�B�TV�CES��UoW^��$[H��F>�]s��M=�q��K��T�Τ�����<�ܫۺ��̯S#�a<U�fY�1��0�ܷ��\������>g���q^� ~ր/%Ld��_��;�&�9튽�����^���|��ovE���*w��yAq`�d����m1sA�@�@T2�a8z�v;@V��љ�|릘��yUO9�Piѝ�jh�׵B���R�,Di�ˁ���ʬQ��<|Z���.��lቯe2g6�C=�o��sa���~j�#���8`�.c0Kdx�c3�7޼�����U�5��"�S���ؕߵ:��W�m����V=�<?o��{�)R'�yf`F�ΟW��HV)�\Y��`϶�k��p�������or�N���pV���.��i׳]�#&���U�I�|p�yE�.us�GH��������iG�.���66{:隯DD�a<'���Z�6�x�$h������`��7BY�\P3Ce�w.�����謝8p�Γ�{C[~���Ї�x��sWƧ�(Kt��:W���M�tato�ϒ�Z��⎂�{Գ���g��E6�9�
e��)��{��)r�`V�eIG�u���Jܠwq���`�x�=#f�J�ya�DVr�}�J{�t����t�.�<c(��H[�0�\�ڋ�=���;��"#�M���5՝�oV�][K��Ǐ����8��o>�����Y��<�Nu�,-���K�tP�lI���nB<&@�AWc�������k�;�(��$E`}.sNT-�ʥ�-WV}�&Y:vA&��=R4�rL�! :�z�q�j���b[{�.��*��in7��Ē��(�N�3rU>��J6�t�Cy\������`�{L�{��I��P�S>��N<�v�����M�G���
5��{b�B9�0�Sf.��Zim�K7�{b��jyޗ�;�`�m�.$A8!WE=�
���}��+���=dȎa^�fv���`�9���s�~�6Kf�V9�lJ��ښ��߱�Y���-���a������r�j!�D�qI:$0�^� �v��p��gm��sCܧ=��Oh{��7[�w�����}�4G��\g<J�F>��Ҝn�-���k3/�`���,��:D�:p�^͊�C��fqiɷN��\��zזq�:�zĴEg��{��1�ײ�Ső���Zf�f�'�'v&B+�u��H�9XCK=W�m=�M�<�É����lJ��\0�7qPY��ȩ�[�W/��*��qq��_Q��s�zʹ�v�3hm=ǩ�P���#f� ����E��9���ڶ��}�A�ۼL�7��W��smM�3�_n��yN=k�Wc��9Vً�]"��W�8F��ȍ��S��׮�vz��<��pԭ���;ոHO�'ٷ���:�(}�gv(7��_�nM)�G>�5I~#e�U¼ț�|@y=6�#*�md�:X����L��RD��s�}�[Q�bL�i�N�c��l���M����]�I�q�]�Ҽ>�w���&�$�φR�7���x�qt|/�xtW/4�d�1�/~��X����u^i�����K�,\5K��2$�5�ЬAP�c���*(+k[��<tb�މ�Zv�k���Lׂ>���O..�%\υ(D�O'+�AJ%����;pL����'L���xY�����$���X0[F��>��#��.1��Vԕ\��t�r�!�]<U�dj��7^⍌rNZ瓂x W��hd��v�cx��},�v^�S��.�'�tǵ�{np9��b,��n@�ꄯ
UP�E�QJb�{ga3��5q�ﯻ:^��y�����LJ��C���C29�Z�����q�dp��$� 2��b�;�XqG��d�@�fki���*��l��)b&���zӮ�J����v��Q[K��W�����5����1bV��=�8�X�n�d�r���I�kGJ�]cӜ��ۘP樂~[��SNđq`ǏE%�(�͢�}t��\Upg�N_m�mb�f?��:Sׁ<-��C���3��G��<���0Zܒ%F{]�Mf���cF��ƴ�4�6PxG��O�,�r�:�HWm�]�n��r��v�޸Z�UNC������~fچW�@V��\�#��1b�=u����+�6��$]i�ӧ��W�wcYk�����NP��U�F
�]��0D7�
DD:�"3(+��BB�0���t0["|�]�&���m�)������&���ۈ6p�ؿ:�#]����uoj���uH��L�w�DP��R]���U#���X��Et^B3;s�\���/J��{Ŕ�L�dϮ\���R���X(�Ĕj�s���\;��x��W�W��a\�˙=����ͻrqK�*h��L��x|�0r��`�9�p,�9��N�=oq�]��&w`stŅW�7<��5u�����b�a��|�������9���ab�z�s�[�ՊM`�G�~e(�ȅ:�<;�=粦��d�.yDZEg>;���ͅkخs�L`�CV�ٞhGF]�$��xk�s���:.뫄�3��R�X6�z.|��=>=���Z��Sc��c�#�/r����Gg9����y����^�]`��!h@�{�v᭳��g�9�ؽ��ۛ��w�Ź�������������k���%tv���!��R�H�0�K��٧;����<�f�����U.�~Kk��wJ�{����Hl:퉔}-ˈ��^�d�Oq�����5S���v�{�e��uIҺ2!5bBq��[l�Ti����;��a�յoo3�&$���W��_dٯR�Ӡ�opHDk0�s'�3����|�Ox��&({��ݎ��|��-*��������p������*�q��ʎE}'�5�yD�cg����P-D8�t�D��WNc�=sA�@�
��5�R�w!<�8���&ΥOJv������|؁ڛrC%�g'Z�;m��i�(�Ŗx�	���[u٪�i�8�Mti\ቬ�L�f�3a,Y�Fx�{4�*��^�a��Z/_�8��y�~�Z�T��:��n�sf�7;%>٥���\`UzY�ͯ���FYE����0��k�+�]��:q�G�Տ�0V?��4�V��5�-��������B���IO� IO��$ I,	!I��IO�H@��	!I��IO�@�$��H@��	!I��IN@�$���$��$ I?�	!I��IO�H@�hB����$��H@�{H@���d�Mg���i~HAd����v@������x��`�� P PUDZZ� � �`5*�"W�"���Дh4��Wf��4�5��J�j@��T�JP�i *�"PR��#����u*�ͭ�f2���i�f��[j3����K�p��٥E&�b�bb��K	�Y6֛���T�R��pn��b��ؑ������`Ż�R���QSf� ݱ��̖إlU�xP
�ԪJ*�9�U*�{YJ��	%&�*��l1��Nv �)�X۸tv2t�٧@�P�I����� ��w2�w �
� uvͅ'`����w:t#q�l f�l�wp'wBl wn�9�Gesjհf���R� �S�����el�-,kX����ح��TB���ݴ[6��m��m��Tšk[$�%�2hj��� ��V��ͅQl�Y�m6�MSZ�7f��     T�L�JT��0@h4ɀCM OhaJRU�LCM�a2d��s �	������`���`E<��SP       "I0��he0��"d�#A���R="b%*i щ�� �&#vv�u���o�g�_��}X5��@��RQ��h4 l�*��6��$��T����?��g�?��i������%�T bQ ҇�H(�<�K$@�"�E�PDOW�;���o����i@]���M�k� �Lv= qT6|sd�$�j
h��'����>��V�Z�3-�Vp{!�vf�0��E��^����$r�1�.=����u��%Hnֻ��jkX��E"~�d:+UKR�]�-7����T��Z)�6vG��<���Lۮw�5���:4��\	K�s�)��e���m�ru��j�$Е���S�Ť�9D,�GM�om�5���X�#6�qC7.Z�3ol])+]�T` ��"�i�5n`Gs% j���zoI���p(2��e˻���.�FI����a�(�fѴ����8��N���n]���T�i����;{b�ʚ��HY�E�����!Z��1��XH�[gݲ�@n���7�=Z�*Lֈ���J*�i8J
��7�&��jIͭ�q��zqU�u�{1�t����3ÈY^4>�=�A��4�4�j�`�w�����T��TU&^Օ@Ij�K�(����)�e^�j�1�)i�snėf%�*j��T�e]�S
��(u%��;Y(f
R@�X��L#t��>�q9���)��#�m*ӧ+I��^��Vv�2�B2��14i�(E�O��xȊeY�dj��ڹ��B�ͣf���a����@Ҟ�{r��VX&[��B�N���x	�5�cE��b���H���w�������2��uP�����5L���$oA�����:m�W
ڶ��uZg�h-ܱ�.�A[7MQ�:���VX��v^n8Е6��f^��#�M�Z��[��rk6�̹6��NԧvD�@k'/�v�����������v�3�Մq2,��'v͠�A�[M�3���,��{j����M(ْ����N̥��b1B�r�eޫ���dc8�m�l,��kŇP�{X"ѭv]�&#�X�a+5��h�_ֱ��M3K$ӱ�a�m	b2�u&^���LfQ-<E��������=�2S7u%XB��ɀP�#q7/0P�S96�e��*�kY�����ȗB�4��ul��K���&J�Y�+,�q��}��������iy�`ZT�:��C5;�P{���e�v)0�<B��/h^�ɉj�ݝ��ɫ�d�0�x����Y ��<��噒�\F�Y�m�Ƶs�֕�N���4�l��Obc-"$��YzU���,�f�i"�]��Hpc/���~Lm�U܅vV��]nU�{�;)���,$.�̖�F�N�~+
�ŽY�Y��/��e�u��ӚV&�5��
�t?�\�obw��4mm��u�q`+h�:w��KX#�:B���Ҳm��(�������ԥ�hb��f�ܴChʅ��u��6)x�Y�࣍e���K��Udk�x�	�xQ��` �l�W�#�sA��j����5y���^kVNSܡ4��]������˨�8�>���v���1o�N�[<{���b�ѥ��&9��2)�؂�o��Zz�|�]K�&x ֚�/���!�\{,��u�,��J�>Ds��u�骳/v���"�(aے�ɶ�4��I��{�1ፒi[�v�VU"J��b8��H�Ek�֫�r�lh�d����LYù��v"e6>����lm���֌]E���6��NH��P�&�p��J蟎�e�zn�Qə��˅R42���ŵ��Ģx/$F�Ml`#!�lLL전���N�q��8�#c��i����-��X\��v���]M��Ѫȷ��%��Ooj
9��P.�����F��1_(W+��h*�����rr�Nm�w�X��Yw����;i�������6��v�����M�5�By��ѥ%$������*:��,�)�[�XKT����#�IQ��"��
��Lc���Ȏ�k�{�
��=%*�j�) 1�&�ߎ��f(�+<v%����u��]8@u㥗���9Yt�w�	v0R�����NA[���fC{Z.�ӗ[1�K� ��ⵔ
FY����@|�٘S�v����gj�5�sl:�6AT,{OO2�*�j/Wf����ݫ�i�:��t�!xj��n�I�8Z
]�j�t����=��+�J�o�;w��i���`�v] ic�@��i:�i�r�]#�nYv���L=��v^Uw�wt�nʪ؀Y6��;͍�z*� � �&!Kl�z�Pu���L���k$ڴ)6�b�����e��4K0�G5��?J�*�Ǜ��ɣI�J������!�n����lГ,ܬ �%�j;g.M���z��7��`�݀��61�����`��W7`���h�����;L����,�iV6���J�0^�3J�*7��x�K�N��Y�d!�/���یm��n�
����.��TM�P�*���4�*3r�=e�DCg
y�"�(�\Nf�ةfnn���Qp�J��Q����I�^����HT��&�],be)������j�̄4�B�/�w`�ƚU�0����
@����
�q�wb�NB>�����2��1ǹ��۳�bܓ&�	f�3ZH����,ԁé�T��ޜ�a�v�Y��������w*���Zr�㕋0�*W��X�Ys�Kϰ�]ce����C.-:�ux���̨	�����N��;��m��w:vv��68ѕwe�U��J�ᙯF������[�	2�����e��t�TĴ�۠n�7���z�I�s/��C5{E�i���ՠ�d�I<�B��g:���e�N�~��uR������H1���筭�2a��鵬Z��ݧS���UV�m�&�J&��Ww{�vt�6K��`7�R�F����5Cv�Yn���I%)%�4�M"
Β�{ہ���\:(��xnZV#Cp<�sQ�ܭt
5ĭ�Yu0f�H\G}�u�]��:�l���ǳ3�d�^ڽ}�
�1����[ێ����Ǡ��4��3��_q�-�ǲaTu:�H>��)Ü�^�V2P]%��6�1�v�mL�`� �-38;	���5%a�����XX7���+]�c�ԓ�Ea�\�����=w"�*���f��:`��a"��;w#<�2�ܕ�T�c��t��9����s[����@�妥�|��ݙ�����61ϒ�|c��x�5YA6���l��B���u,D���Sa�􂯑�6���
46�7[W����@�Fr���멎�h���@F<�w�2�[���-��U9���T���X"뺒�l^�2:��$���eÑ�Jv(�[1n䲙%�lM';��H��fo8��H46��eu
v�x�<�x�w\N']�i�t��e��&99��ޖ����z7o�q�*��)F���C�3G+u+�2�nf�{#�P��J&�	4�T�}�L����F��UH�>��؞<\�H-֑|#%�gV�9)m7\i�ز�\��4����/�t&���n͛�8J�X�Ӡ[
��7f�@�ɒU�7�%�;ʙ 2�e2��f�Fݣ����:��S\�fl��8��м�h"�;��b�[��� ����� p�F�h�׹i�j;T�.:��(*0�t��V�ؐt��;Wl��[Z.��
�V	�h�xm�u���xD����"��Q�ds��'`{�����^3�$�w����F�/�n�i�%,	:}>���GoQg�Zz�cd����7O2�S�	�9���F�f��F�[�֮�;��^���uޤ{�0yʀ�1����CUk��i�t��U�aM�"T!�m溞ojJ3>�t�2�n��`t�����7�[����>�l�v�/2�lTD0��?h�N�WXMm3J�^���|Ѷ{/���!zF�����*J}�@f�.t�ʺ|ʲ�`�r��Yx:>�t���Εv�!�u��|E��V�wpΣ}]n%A����u@�*�>޼n�{m<"�j��*k&��+pop�L�:sMd6xѤ�n(�'/;��h�`�wA!�grc5�ʽ|ĝ¥���|7�s�# �����0â�T�T򦆮�b|��>�F(�i ���e���n$���(uEc�m�|�2����K�ٳ�c�M ii�.�1�C��c]$����}�v�U��CŤKR-
�E�����V���x�VF7����[����>��ݹ\�J�@7.J��KB���g��e��2��>�.�Vj��'˚��l�"����s�`V`�S�9���� vں�ьV�ǻ�`
�N�|�s�����0W\N���aYU�>�.g].�1=�2�N �kV�U]�\�7k ��X��2�+��S�`�$�2e�rJ3'I��!-�yW0E��T�!]�ǒ��w�����i�xz|W>��w[�*��f"�ì��e�n�:�V���Bfک�^ڹH�A�^�ƌ�g�m :�]����_f�e�Փ�mp�	���
���yzf�u.�lm�7(�WŤC7Z�H�h�-��8w�w�9�4�p��Q^I�DV�*AG��tr�o��_V���&�#X�4�b�{�U�ӥ}��>WQ�e��E���n�yˍ��J�/�<H���[=�%�%6Zea��U��>K�zc�>�I�$G9E�+��T�G9^6��4!��k�������e�ͺ�8Rĕ쮕�^���˻[E����^>́������2BV��0�f�6p��p�ې��n_�q.ʊD��2���{�w�wǑ��rI���*v��l�r����U%Сhvor�d�P�2��L4�ix��M�3~�-V��9W�u�7�#�H���v�G�#��T0��{3�69��4��N˜�˜��]�P���51��̘�9uj�}�v�8�z�Y�H�5o���i��Yʕ D�f�^��H��\Y˾�k�k��{�K)b9��.V>�6�%���]�w����v�W+k��Y����v��9٩"�h�]�0�t��͕r��T�3ڮRw�|%�<�)�Y}��]s�ݭ�(K�y�:!%Ƶo���\�0Á�u4a$���	�2N'�D��ĝ�yg�e�bkD����HK�<�c����%Ye�˛���T���_F"S�j��l���n��OE
oH�/�Q�zE���6U��5�*���<qyת����*��O&k�^a���<��Ռ���䞠     l�c!���5㢱]&րU��     �0ؐ���:Ԃo�2�T�N�/S�� \�o3�H�_���P����4�JO�P&�{���%��k͕�I�c8���L��؛:ėL+k]�9rc�J�ݎ�BGbؾbm@T�I6�=ە��
�Ґ�t�����*�^^���i�R�97���҆�]��y���)Y+;������V    <ce�� �m�?35�^�Z *sڔ#޼�7exV��$!k�@�1!����``�Y�^ǌѦ� K4 �xx�ט1��0   �    �]���FO�u(k�YV�����}�ߍ��gS�s��;{:u1�=���  ۔�����DP��ʃ�C��I*t:|�����#���Nx��s�v�������!P5oS4@��wZ����g%��v�v�IC�F͓����F�4
�d��:��b�lə(fͫW�9uzmA|���Q�F2Lۅ�0dS�����P�Z�`;`!]-8\4iR����E�j�΄�Sf��90U]��T:v+�͵��Ĝ�P���n�$n�ȫ��Tp�{B���FQ�ajͳ*T��x��愭��*��]DP: /���7�@W=�s$tE\���tu��`XrJ��<�U�>�2�{ҷn�Wv�r�C-�Gi����[kB.�>�8�h
�q>h�Hn�s����YC�'��^��Η��)�N�|��ܶ���5�r�Y@�V�r�y����C�R��5k7n�ϛ�GJ����/l���:�)�k���0忴���Z�:��u!�V�^��wӜw��F��Q��,.i�����;Yku|0��mu'��rYz�;W�5�T;ib�`$
���VRT�%�ʲ�������6��dPn��NE}�;� _OE@�'Du �I@TB�u<�����7�LbmFyh�w�@~Vy�Y�˽�ΎR'��ZX���7\�I�9yCKY��w`�� ^8��ԎduŗyQ�h�dS}����"��p��,��Bj�G�^�型�mO�g̓��g��(.�Z�j����$c�`뗻�z��Hy�5�֛V4���p��,�H�����<ayQ7�Ф��,��̅�Օ+��x�m�c����k*Gdc�i���2��FL	M���e)G.�9L[��b!e��b>`t����}V('����B�l.;'�OE�z{]�ڳlE��ʗ�)	�r�Vw;��EM�g�z��n����Y��Ǘ:u�MR8^�l�ʇ*Q�l�����])"L|�/�Pڽє�=��CfS��s�d����8�,��r�L@
���1hi!D]*b�u*��JWZF����3~��{HZ�
շg�a]ؤ�.󵪲���W{e���I�F�E*¾�o�A�.,�r�Isq]hr�Ԗ�6+��D��e恳�M]G� ��)�g\|��0Pgn�Sq���E���-\&�*q�ͦ�,�ζ�
��"���f<�H@7�Z��.�e���RƤ7�\�5�d���v�lf�!\���TkRd!�J�b�-fXtv6�X�����W|�a���+��7C�6-�i���hY��^�9�����n��[��c�N�<sˬ�\���^���`(��E�ɕ{(X�FY7��d�o���꿯8�Ev��%m9Ӕ^m�����dv*��U)��:۝ݺX�4�̎��2�v�VaO��V�]\�����ֳpϷSB೯s7ghu��ˤ }���ë�ݲO^�ë�J�G��M�w�}iu��9���SD�+2�(T��.c$�v0�ܨ��ƯE�V&�K�$��C)�vb�Tr�7I���n��ۧ�h��ֱ�!��
��J�PO(��l��T�]AwWj�mv�q��JD�]r�6��
�CEգH��˻���7��_=x�x�BLm�v�zL�g/�N
CUH�F��qb��F=���SǄ�xj9\6�д�o�"���RVVt|ݬ\q[��y�]�L�1nM�mUپiR�Z�nn�XQ��d��b�v*y�#(.4���	��e��B�����doP���0�wxy�E
��'�z���=�1�3M�^N���dSK�=���:w�3����x������p@eo;Y.��������pBu.��v�v�f�X��Y��8^V�
z���Y���9���a]���@_����Z�g�@�[������;ԃS	��:��<�ΰn��-i۶*�IEX,T;��G_)Z�i�;�o�6ξ������)Zb]�[���j�D*�Zê�"�
'��<�g]�i�̾����|@�q5�-:E��U`���"�`��L�U��C�v�-�&�o�և�8�e�j��V=:Oe=�-��y�٨�[(�ݲ���ޭ7����e�͌��r��!�up�]6��c1�ٗZ��ed]W�V��V^`�q�R�*��1M�b��ʦKRڵ.�H���a,��fZu�T���v���zY�f����k2��3s���ʓ�Ao5�\A��2�T63V�QQ-=v	Pv
�-�NDEVeJ�maĴ�F+a�w"��Ӭp�j��WV1�5��u�+ҁ�Qڶ���Wu�k���P�ڗX._s�<����Znr�N���N��[b��{�����Rl�ֆ��civ��ݐ���Q�����Q�:OopQQ05v{�]^ЋV�l�u����p�Ҥ.����vm��Pn6�P͘Bh�hQ`��]�V�Y2*6�7H��{�!4mÅgi	Ig��.��k��[v�a��J��;6%r�	wdv^N�Ҏ�_e]ze>͘�SOƹ!r�"��1qTٻI�XZ�t�V��y;�!`�wv �(
��G�P�}�� >�j��B��ԅ�+rɂ(�_c᳹7n�j4�M���X��|�kD�G��� ��s6�,Lk:��,f���=8X����R�94�7�9�MdD�k���3Gz��/���H�C��R-Zzsj�uh\3�L]n^�D�y�Σ�)W!N�-}�;�uY�'!9s�TH�o	wq����5Z�2u_�o����9Yv����87.�;;�\S�k�J�U��PJ͗9�I�Y	n�ޙ�S;^լ�� �'ކ �I�w�	gW�T4D�o�_��{�gx�sA�;0�\��i�k�ݓ�[ݥ��3`��AբEI��8�и��h���ejKZ�ocЭ�J�gXɴOo1�w:�F}����2s�{��})A��H�*��Z�$`����s�闲��U�#˹R1������>6u�̩��S6,��a�^A�D��|�-vN�g/��kv`E��6�ݑ^�#O���N��SRA��z�4�s�iF�#2�QWC��� s��!)Z���ԯ2v�      }�G;n"� @-�TX�&F�4�q2���B
�p��$�)M�!"��i�kI,�L����0D���`��(�"T1��349j\ʉvɒ� S2�B�������5�͕ʉ"	.T��D�2�I
�����H��m�Ȋ#��JnTD��	���A�E	�1�c��v�&2#%��b�c�V�[�I�&Mf�;�~��nO�}_ݥV����o�5�(��P��F�=�6$��Q�]�������? ��R����<5{l����U&�GsqO[e�邖�۳G���\�A6zOB�2X�!�S{�縜�����[23'�;=넯z���������Gv�
�~9��۱ ;�?z�Ts��1w�W�z�ߔ�m��n��!>6s���n�նl�"�A�l����X�C=���y�v� �*�ٟ�z�r��ک�fX�=�^�����\%h���s����-A.�2��ui��{��W���wW��vy��$Z�viwov�p_�)){�gqNܞ�>�M�*<X*����9�f�T�v:���2d~��9��������Luaݏ5�+8��J�ު66��ϻ����f�B
������r��˫�\�}{�,�w����ιXqAF�;��G(Yyv�)��[໫�V��ٝ�U$1�$��M�&��ȭk=��'Oݙ�ʘ���'�)���I�v�lW�@���m�l/{8%f_��e�g�z�)��P>�Ѽ�_��E�^ܯ:� \�� 8��wz��Y�,��]i�YFvV�k��К�J�X~��+���5y��g�7����P��s�.����>VW�ϗ�ͺ�v���ڎ�mNlf���ך2��̺�����M\��7�HVm�q75�P�{�I$���FFèbח���K"�ܱA�L��sA��}�9�0�#
�2�c_���H`C����y�"١�Rr>�]��n�4(��U�9�;gͮ	߯�0�/.��V�������^_��k���]�=����w�XF4NQG4�ַ �w�VN�#�Ț�X�8_���a���ǝ�e#�����<@�?Lj�'׶<��V���y��fe��q���ˬ������NM�c ���"z�{��x�_]t��ܟ3�zܼn{f{hPf�O �����k�޶�-��/W�ލz�	R*�Z�{����}��L�Cx�`|�e�2���o-�Џc�h�O:��;�V��N�1�C�U��!́�6PĒ��Vn�|7�P�M��{��I�O��]�5z����I�,-0��rNW� ��9ṳnRS+2��w��P��/�G�)����l�B��f,�7Z,�*�Q3$�x��x������z�m��-c�{��ʮ�+nƬ��%�>X,����4������k�dly�g��b���y�v����4���rΐ�r;�
��l���ԧ�c5~�_�:�ע̱�}�WOre���� ��s>�:���'����,�my�sПx�{ݺU��&[�����{^Շ~=ٛE���nq��NڻSм�;���lDW���=ʐrf�r�lv6�[�:(��!#��!���n.'�9FU��W�u�����ԯ�QG�[oVy��I3p�uly�^�N�y�Uq5�vp����X���N����=
�/�6W��{]�Z��D�}�w}nH$"���]�L������k�N�N���;�]��g����x64wg�!�g��h�#ޚ����)^�w�&^w �`����*y�|-ݒ�5��j���]��#t7�+A9���갨����m������~���YpeύН�������C�+	���=�ݗ�I*���*�"���爿c~�W�Ty:b�^����^�f���h��$�ʞ_���'�h���\x��.'"�N�gn��n��B����������:������n��^�=ϲ��Λ�Wz���ʼKq�s�B/t���yO8���h�Y�^��ΫDq��N��V���ʹ��m�J��$�]�ے��ѹ%�IΞ�Ga=�&�B��vnS�:^���M�굯lLڹ�Y�mt�jy_�0���]&�����֧.L���MK���f���w�u�,�s�_�[��wZ{{�/���:�o�qØ|��_�9�Gj�5�{���2��[�Δw77G��w=Z/�l�R�2ץm+̔s���۝}͚F�x*�C�mu��ӓ��i��/.S�������~ @�wvp���Ȯ�~�W����R�CV���;����P�6=���n^����:|�U�u'Wk���X�郥�����&�-v��m܊�����ې����Fn���$��W���R��xTc��5p��df�=��u�s��,�LQ&#�;�{0�g���	���5f��99�m�i�������/��2������F����s�h�bt�e���և���uvz�z;�:�m�Z�Դ:��ky \�
����Mʳ��A�}y9��;A����[��G'v���K���ic,e�y����;P�{tSK��c��R��hhۣ�:�T�P���a5��X�|inQ��¥Z�R���B�c��u�����t.�fL������E`�ň�n�n�a�if[��uu�3��6:Tv�&��*�5�%X��[&O���K�י��׺��W��=�:��Vi�K(K�m�5��MB����6=�e�)�Cy��~���)����Jǐ�����勄R�	��uhmh�v�d�x�Z��}5�ȟ yl��a�T�W�ёD!��Ч;ť	|�u�E_�>�������d�CnSl�6rN�`.��v�&L�+�-G����M+r�u��G�b�FS���X��&6�m)�ekDS�[�ʳ,{=�D֣��:`X����H����mx�F\a*g�Hdۼ���o"���TS�M�*T�������FX���%�t0c �c4e
�U����M�`    @}�Τ��D� BIt�(��pP�L�	/D%"I�(&yL�4�!z�dIQ"IaM�j��E��@��	pIeMSn�Qd$�GM�#	*��{�Hq�$K|.k����K�
��iI	 c4�(�\i�r�D9JE �2�i��@�%�E4�m��L\'�H%�hQ�Yˣ����]�g��Ͳd[n*�m�����/g�����8U�`~3���<������~����ME���4�r�ۇߵdxY>P��[��?}��싛�9����DmM�Ǹ�}.��K��QQ�c�|�p�z�M�z��?���zy�E�%-�x׼��~Ѧ{V�Z�OI��W�dy���8x~jf~�~G�X�8��W:��v]�.�x�9�8&�����к�a���b�־f��}8�[�$�B�%,����s�k�k9�3t9�e��h"�Q�&�b`^�5������!u��6�*��!0�@n�+���H9]�N����F��?_���sJ��ab�w�~��n�O~��M��%m?O��)O�{i�8A�W�l��'Կ��g�͞�h.�;�=���?/M��V������Vj���EW���)�eꗷ��E�B��w�k�P�dގ��n5wVE��Ƚ���C+�h�w�\�Yxٹ�f�-e��Q+]��/��\���tkQ% ��Ӆ�\�)$S��4T��?�_��,N���n�}�e9�l�wN:-���g�n?x��v����M'��%�yG�Fn�b pp�?!�T�S�Z'���pZ�g��]O+��>�Ϋ>=w��+�/2`izQ���fLÆ�ydmr�LE���y7���sIa^g+8������R9l�D�t1d�0��^cm�Z����I+,O@�A;ۮ��a���]Q� -�o��,۞���pC��hB�X��A�Jd,�'��՛K<�7�zǋ|������bf*�J� ����=K�4k=�{�x�3�����r�h�,��q�=q�\�
���">X������o޹��/y�W^C�w��\[C�{���I|GsK:�͍���V�o{{�w���}	���Z���𾾲�����E�+�f�m��j)�uu֣�ؔD��J��v��/uk
V�$�oXT�X�5Cv�h~�l�ƽ���&�]�7K+`)�l�ɍ�$D�$Ds�;Eg�~#k5z
'��=��B!D�P>{����y>#�-o��F��Y�x�޺#��H+�|D�]]��p�&}���?O���^a;���{�L~ɇ=��Y��o�q����}�S�1�i%��t��
Q�ͽ�ۛ��vWLL���B}ÚN�E!�O`N�{l�=˜������-��?��.�z�����vʳ�e�A���ҡ]{�u��\U72Q�=v���D�6�����0`��kw{�����+��yK_�D�^~�o���#�W�_D��%jxt��W�s�e�^�6��=k#ՙz	$��xo��v/	�_2v��w������l��m���p`K���=:@�@��|��8>��{I��y"������/�x�}��G뚏d�����)'�B���0��<��:@��Փ���\+  _��?]�=]���n��
�6AOa郱9%��x�?�N�<��W�g��G�a��o͸�����n�_����z�=���pFAۨ��*̞y��˸#��a~���dp������݉�Aｺk�㘋����[��i�M�V�]4o���C{5}�t��Ϩ�𧼃}����gE�S=b��_��;�<¥zf���%��ܖ�r�y[A���0>�'�u�u�]�a�u���7X�(ӣ���ɋ?T��{s����F�5`z�
و�0'�Ź!�2����G�f��ml��f�5yS�^�PL��w'�s��^�0�X	�N�����z���R�dqW�y��W]َ-T�$2Su��y�w�;��Ւc���Q�<�g���ގ�ن��j>��gS-��􈬴>�+oC�޻�.���6�Ό�M+��fw��i5���e?���W�1fǥ��KWlR� ��j�
��B�X�>�Y��1r\�k�?������^y��ǐ��%6�05�$'x�������/��JI�R�� ZL��MK@�sv=��Q��
�<�<:v���;^yO��VxfW<�碼��uǩ�v�2{K��ϸ0��Q
$�*�\��z�p�H�Q"��/3�5ry>�lU�u��g�������wu���M��DW��%�긑���f�����2_��Z�k�{�>�g�K6�Rz��2nr�D��]������Z��Ry��͙�@��Ғ-߄1�l�DkI)����N��mM�֎y�����*t#n�`8z.�5J�1+"���I��3�~׽G|=�W����Λ�ǫ��5kd�w�����<��]���K�h����.畊���9�
�����\R|l?zz������z�F��@��1�r˃����͓�I���x��y^$�W����~g���T� �����z�S��;���k��EӁ�w�X���
�B�ҸF�� ���+7f�|��h)ƴ�V�*�]��vek�
�_�qe�a��7���wbt�Nj�.j��4]�9u���]La˥�ĘX�;Ϣ�S��(Z�d��R�)�f�9p ��%�9?�a����VC��h.�Ij�������P��j����q-����x�ݕϹe�rv�QQѠ�ƩU�4:���nTF�S�ʻ�2�1��V����y��"��܃�s��r�Z#hХ�ī-��[;�}k��]{�ް@��2Q�'E�U��kd;z����A����	�����7��O"P��R��F�	H7{E��b��v���aq�%u�a��܊�X6�&�m6�*r�ck�f�꤇	�]Xj����7Ab�]�8���M�)ǎ��S8[��\՜��[d��v�]�B�ue[�b�-�I�zM�@�!V"�zˑQ<�w|s �&�H�Hl���/3R�`��gJʝ�i�P���o������̘�&�|T���a%�����xx�K�dN�Oa��x3A�   �{��{ߖ~���Q���
I!2FO�@�S���lk�2'�;rQ 
� \�å$��BUL�l�UJ���RB�!�	O%H�!�14ܴ������"M:p�IK�R�(������hT*��&�t5I�әSBr)	M��p&1F$
�&�H�tL�]5�KM�8D���(LL�T�L�Ɠ�2$�v*#�k�	�)�� �H���3-�?2O�˛�z���=Ƚ��.�c����y��= ����"��=R��������U��w{�z:�y�N�k���#�G���y�u�Wo�a"zN������繧�c��KnD��7�X<�A����6E���\��͚Tӭ�ol�x1�>�ޘc����[�����c���P���E��勯+�S��+�zW��6M�i��f�>��|����佺l��nq}rB�x��Up��w�`�.��1�OS�����ٸ���Q��%�ocrO�}UH�I{��/_䛘;�����6�G�b�K��\���7��:D�h�7v$W��`��+�0��oՉ�2�I5�������O_�U�
�DtB��fHe�/�]*'��k�I����`ۢ���=���@� (޶�ܗ&m<qy����[��rv�fFKʎ���dB��;����ɞ�D��\<����|�ʒ��k���Ԭ���e#%�ύ���(�-����-1��DDF�IOT�w�*>��G��NF���_�A7�S��l���}�j��m�>f�4���xzxoI�}���_*+NG�5�޽�Z��񗮵�q�%���]
b�5��Wb�E{�nő�ԊW�<�z�n�[�*�y�u��<�xrߡ�Ħs�W�j�ةrO;��M��0�����s���f}�}ǽ�Ј��B��K�i�L3�,1�w7�Y�8PYF+�yq�Dl-oG�#b(�\�M�E�;\y3[�c5���""Ԕ��o��+Z���Ά�S˩{.�����9ږk��y[��}����,��<��/�ݸ�hi�,�@�/��vԧ��;~3$"���5���2[u⎯*u���՜�ww!�w<�Z|�lPM�L�Ḵ],�޻�y�F����U�������W���z�tϗs[�^��x=to��{l�D����$
��s�ʋ��� On\κpi�����W1D6F���Ǚ�n)�����m�~�""#�Z�������畻����T'���4�Aͤ���j^(�
��)�P��tGצ`�o>3��|�r	B=�������B�=v�nu�O��4/����~W�z�y��
|�>��9u��L��,WXhyp��/h�90lJ�{ Ȃ�^��7iȇrE,��������$�]��T�y��P'�q�
�W�}�#�v��n�ɝt���j�׳e�x�)X��K���[݉�XE����H[fI?W��}E$��~����*߇�������w+�%�z��{�KdUᏟo��F���b���T�霒�͚H��*%��t���?3�}D�<�xJ|�+3<��T���,�E�(B��{D=��޿/���)���Z0�W�x�,%Wb>S5�j��pۨۍ�������V�-�b�@�aD΢2�ɪ��
�ǃL3&�%&_=��(Wc�Ý ���"<��I78)h;j�G�lnI������"RY�صp#�������ff��,� �c~�:V4鳡��ϳE��G����Y$��җ�,��w�:�}�[1����}O�H�s �^���1�M��^��K~ѻkx^�M{�1�/�P�Q��wb��3�V�R�V7��xzoz|��^[/p�F��U����h�W���̟Z����Z�������&q�������a��E|`
�j�����x��
r1N�rd� � }�?~��ZIN.�T%ws1⫵��(+|fܛ k*�ѓȪg>u}���7��an�x{�vni4��[�H��q���T�J�co��;�`w�YQ�X�aoVo�rn犬.��R�Z󥬅���uL��sX���M6"��}ZVaY�0��㊎���l^F�_V���������X�>���ү6�v�C�%��ux���:���7�1�������L��N۳�iM]�K]�:Mj@D���"!B�������|r��Y�Wz�����C޺pU��ޫ�>ded�2x����Y;��iu�h�l$]��۹�S���c`Z_��y��Ӓ���g��`j�$��dqC����]�4*�����=�^ܶk�b/+��9錯����v8�K�}j��<�{��[��<7����W���2��5�3�n^=�%�ʒ˨@�/qXV��8�X�b
��رՐ�˦{f�QO�+����'$�����}��7���?�]�}��W�o�9v�����*!Q敝�0[>B�VAO�lݸo�ʪ�{1v�9j��u�Ҩ�yW^p�3n�{o�ۗ�<����۸�
[IY�>���5*_=8T�{ā~�p��<�UJ~@�Am� K�ne�[e^s�1#�|����Agw�*ۣ ���_~��?��}���OM1�ڦT�� X;���[c]��M���7�ѻ�sb���Y��/%u���G�q���KN\�����YÍ��O�m��Ozp�iԡ�p���I�u����t���}u��;�R�~�YޙS�j;��"�ͧ���2�T�6�иq+�2�WZ96�y �\'��n��S�]�o&٬��t�Y[�S+醙�T���ˮ&e�zj��L���3��L��3z��9
V�� Om=�M%L]���v�`G8�f+�t�eMD��Q�m���2F!&ڜg;�R�t�v�y�����r��c��Y��]؂�d6�A��ԾٓrS4,�f�[ck�=IT����Ԛ����8�y[��l�sc�����k�:vGj��m��k+���u�VJ���{]����W*-Wa�p�j��V�Q�'�ڼ�Y&�+�¡�$��¶u-�[�&%��
��4���2e
�]CrS���\�	�2�l��=<O�1�>�^�9�s4Ҩ�ei+xd"칼3.rL�����a�!�Wv� M�O���lk-�V$�񓕠&0 �  h��a~P�6A�rCn!��*p�Sh�S㙓��CN����RB�l&���#��UCr�`SiSMH��r�ǥK�K�A$UQ��pn�#��:o8�bb*���P17 6!�! M�D�MQS-�l�Hʩ�4���*Z���M�K dC��j�M�q�* �DKr B%�R��<ԔC"P��PE-�ʆBp�$J����D��6�Bi`L�!����MÁ�B�0%�R��Ki�i�52��H�6qn�&��t^V���f���Z �X��I)����?E�[3�5��w+9��Wg�$T����&�f��z��j$�\�o���ϥ�(�8o7b��my�=}�`�f[u���A�������}�'�,ޡ�B��y��|O����3��x�ח�{}eQ]�������!�t����3��>��+��0��}�<=�z�2�O|Ó-
�6����AV�e�NB�ɩj�!�^��q�eر�oq�mHX�K$��ڑ�Arx5�������(�C�����?9N~aA���\'����P���1N�^����z_t��9o�iv�����$��M�ѓޢax��Ϩde�vt�";^�g����G׼��\�K:��<KѺ���=>����{+��AOefv���ۧ3w��ӲX5外����n7��=�K��6ֻ��=�|�V.=t��8}X������
�P*	Ns��onX��6���}��e���vV���TVb���o�y'%c� ������ѭ$�+��%x�y��*�i�b��?[>�ˢ�Q��7�5���^N�a��h�f{�<��)����ol�C���x�YSz�P����6�l|��YU�����Uc�]y4L�������C��ZG]sa�x#�Y�~[�S�X@���󃺑�՝<��~�6���ᄀjzxz�e��v�Q�pz�T���5~<�z����eMI��[����q���m��2�����_���s���߿EI$��~����u�L(D�Y_���.�承�ӿL�F醶�ǻw��t��1^�amQ��_�:����W�xi>q�9�pW�,�/��2U��!�P؏�"�����`�~�t˄�d�|W'2��[��gs*Y��;���N*%c���ݸE��u/��w��6wz�J�%ύ��ֵͫ��F���p=���/*�*����*��4o�䈦ao�-�[
p[V�h�L(N&&6�\�WЭ��v{���������ߤB_cQ	�Db t�#���"��S��x-�.b��P�nx,���_HZ!�N b�+�]�ŀ�[f����f!~)P�/�<�LAs�-V�7���<p�Qb��6��-�j�����&о����mR;�-�	�F�����/�ߌ��QZ�*Z��+x�+x��������� �\`�t��痎ep���"$IN8�0�m��b%L@7�����QB\��k��y�{�T%"!{ZAo7�h!~iLD1-/�1 �S�	���睱{s}�*�ڃ\�1R�P3��MD�C1�Q3؂E�S��l^�s���i��.�1m�R�Ss�CQ�1BB�0� �0ő\E�M����s�
d��6��!�.�3�M�}�R�R`�zF�b��Ø�$�	h�/�|=3_xԬIx�_
�%LEy�b"�����)��X�	%R�G�%�8P�T���|��\m���{��U`�a������鬲�{ѐ怋ņ���w����g{��w����DDDs����P���Ɨ���ځ���M�)#����;l�%�)}��S��	i�/�����}è9��'��j%A@�P�s�EM�\��!PR@q�zH����������Q�(�$�Q"tGs
��D�MDu�S��M�UMB��<��}�{�|�u$���	 Q���b#��y�5C �-�o�q���!x��Z-����V8ߛ��5�-� 1�Q�D�)W8�� ����RD3A��	P�97󿾾sܿ��Q�J��j(H�"Eq���K�@e��XB�裤_�P�F��~/;� �x������x<Avx5�Z+���*ox��3��16��+���!-��T(^"��bP�Z�A%C�<�/��
b��K�2�M���<⹇u�z�D�T��V�b���/Rb�J�@��ys{=Ԓ����C[ҧ�����q9���1
לB�	pTB�!pJ#{]\s|����g��y<���^�&b�\2�Z�Z�j����=�K�[Ҥ�D��n�u5-�r8�\�.I�����I�����W�" �E�Cu65B��l����� j�i�m�KA��E6��R�6���Dh�"�X$���^.�A1�K��J�j�P�����s~s���ϏBd%���Q�@� ��[f��F�P-bµ.XB��P�J�K�]�o�jP��� �T����\�$�@"�(��&B@��IR��{$�k���	��v�q�l�7��Ц�5E6攼D�B�6�"��C0�
z��'�}��	|$
D��D�bK�<D*"fĨ�!�L�ͨD�E
�F	/f�z�mQ	�%��KGx�c����x�b��!�H�%�v\D&�i`��Q�<BXD+��8{���	1&xQ��"8'�{��֮��w7^�~����E��=�:��{�PL��ߐH+]Y�{�z8��`b]�{�#��(������!�.w{D�"�cU�ǌ�x��u���v&���{�Ĕ(�{��o�V�k�{*lG>��pE�խ\�n��i���&S�}j���J��o�������gq��u��zw��
��Gx(=.{=�՞稦�US��c�j�_KZO�~�Lj���6ݣ��(ໝ���:��-S���.�jϕC*{�ĺ<�g|n������ୱw�;҄�+ݵ��bB m!Aݴ�_�� �y!{*��Bҡ�mn�!+e�9�D]�J���3E-�@>���?BZ���~UQ����w,��y����E���x����Q���&��y�Wm��Z�.8]��d	�ʞ]�g�7\j|T"j^���O���ܪHWY�](QH�%��ӻ�3ҩ�m���1��]�9gt�0gG��}>hG\ƶ{y�������y/���c��>k��y ,���^���j��ח.��^��oi�U2��%��s��]�lE�4w���&ͻP9����0>�����ܒW���K�Mh�������!�~Y7�,4���3��*��� da�鏬���b�)�~;}~Eb�`�^���v����%���:ךQ�`B>l��+��Y����׀5���*���^�jM�{�[Z|٩��L��=7��������\i�����ݸ���k�E��_��A���&kj���dj��Lt�4f�� ���u�Ѫ�t
�e�� �M@���$#"�4'����ᛮ��Gҷf_b� �yK��6��p򵊻v�G:����µ��ⱛ:�ox�+�cʹ��?��8�}���)���g8������S����:ͽXK����|��%���s����%��.Ӻ��E��i=����u(WZY�R��r�ꏎ_(;R��@��3ܹW�Hj�"8�`�kхl��McXk(��-Ԇ��|=���+�ߦ&��U��ʀBR���e2���Dh�:s���]�m�NP��a���˥�{K����pIw��h��R^7�Z�;��Ƭ<��n�";;B��̭GF��
T]ZCvj�'��ٲ���U�X�حt�#��wa)4U��Y����fɎK�Шk띰c�mR�z��	ö����#6��!;���Or�aLL��\��8	B�y�g�ۏ��p1��.��ok�(�f�r��WО!Io�m�Jۮ��u��D^�\�����ǭ&g�c.� l4`���@��\�H(V��=+���   ���uL�ɩ������ b�B�L��nE3.T�� �4$���bY 6��l!�!rX��D6�.A�R�cl�8�!�|$��b8Cl�4�d53"����JN$�S;3>|TǃRӄp��S@�(M�I-2I!H	��r0@�L���4�L��r�	���Dr�m�A�3G�  �b�K� %\rB \n"�P��"kҥq�8CJ��0�ʡ%T' �N$r(��������?L�s4���sS![1 Z�ߣ5��z'�F�TL|xR���8|�
֯�~�7�b�=I�ۥ�|��^[���;۪��OJ�bX�bz�'�x��f�fAp�vO.c���ܩ�+J�8NjӼ�wit�&�(��ŋ
}t-��g���sON�=l�u�{�U*ɼ�_	�A�ڧ\����l��������錺�v��|�ON˘�;���P��3�ܫ����w���]�]m,��3�1
��ZN8VL�[��]�1�����`���ݷ��u���*�ew�2�� �VX���@���*r����p�{�Q�Y�S3/�b)�6{��oǜbLa2k5����4�����
~p�n�Z���q�~�����mt�i�0!x��vc���tX�5�z�rg�k�/�\!L��k�x���6{u����g��a�Xp����s39z�D�uͻc�u7�b��h��n/σU٬�/�<Q�q��8���E��X�h�.���V��W�3��resZ�q�4���ih���s\�ٌD�'\����|�Q����W_�T�D�]��|�|�XI��-�>k��[�wҦ޻���[�+��Qe�3L���4�ݯ]��OvWl� ]�HeeĨ��r �|�t)VXUz�bޙ�ϳq[��4�o6���ig����~���$�WW�8jv~Z�<�X�Re9mtVp^ڸ�o��;���֚+#��_^
�^"E-5�����s+-S�X%��.IZ�8�a�|�]﷘��oZ����t�r92�WוR��a=VMJ�_}�Q�O�	B�i3���m��s�nmw�;�km��5�vy
�0K��y�֬���j{�;7�q,㎱޺BX&G
W;��;��N�J���i�kw��J���3��ۅ�]z�8+���J��.��J�g�Փ�C#�~F�Z����~�>}���>���J��N�6 {��䍶K8�)��]���T��'�u(뭍��Y��]�mNׄ˒�}�{�D$�33
�	|.i��+ҹ��T��e�$gsuDnmԂ� �]]��������uGZ�;�!�D:xEn����=rxe@���²���y�5y}3�N	ۺk��g1��s�Ib�ڦ��K�U�fз�:��)xtVEo�KW�ӳ�fċ���R��0\���5Tr�}�����zT��8�%���2�^rM����J�]��6T���d��5�����c���K�r���`�Y'D-rYO�=Q�U�V]"i٦�Y>r����f	L.{�ӵ���;�Y��� }��r���CN�Т��dZ�M��
�*&�r���*pn�`}��F��YS�+�U���c�s~
���������^o�a��n4�A�4w��w�f��_N�8�귕v���V8}�>7Xa�'9�x�����֗EIѾqE�Y�%Q'��ޛ�ί8�4J�	�1���΁vˬ�ؕ��c��L��)ƁB���.d>�������gu��[��]�(�U��^Y������vBK0��q}�ѶՐ*ɏ9���Z�B��E�����ƬY�B�~NSu�j�͑4��U���r��-Y+����b��g>w�*m�U�ܳ���*������s�]Օ�J*�Jn�$k\��8�&K� Z`�?G�i%3Q3��^S�V,"E�K8qq��K�R�ɪ�É�蓂��[ݕ1��`�Xs�4e�>�Y��<���]c[�s��:��H��k����Y��Ɇb!S�1e�W��7=�t�9�X��mP��W�*���^\qu�㧌�����3�f�gJL�.7�uǽ��3�����13Kq#�蘎8N]�쩥�~��a}F�E���^#H�,8H�Q�=|~����_�/[ۛ'�:#l��s�+.�x}����O=~&�5oƕ��+�iDV5vl���=�r�p���	�
94ܩ��YkNu���d���e
���!.��y+�O@>���R_�������|ms��£�*q�_:4����)���z㤭i�Dn5�9�^p�ܣ|��u˾��0g*\pǤw��)T�=��;�<�̊�̩l��ۮ�u^���������TӔo��X� ��v)2���,�sy�uB�xU&�r׌��|.�p^1�V�Y�e*��8R�^ʧn��}n߳�`��:M�K�㗤Oj�[/��Luظڡ_�R�Y���W{�Ӫ�#�]P�p��)3� 
�����޶n��=�����o찂�[K˘*��]9�p�FiܥG�o;�*.�V�(�œ�P~vLD��M,�3���%4�2m6�c`G��i#�F�c_"|�ˍc�t$cI�)���&k_}��i�`�%N?�Ӟkw���p+�"��N�~�t*�}��}�'Җ;�3\{*Vx��ft���κ:tWy �Z�vtXt=�e�"��ٽ����>
GF�h2��T�m}<�V+,v�#���I#���};V�a�xw����'�FK�xYm.=9��W��J�����|~��cO��c��j��G-o�sӹ{sA�`�;'k�<0I�x\"��͛���w��F�<-3]�(��abʱ��?gyY���x�+�I_u�3��i69T}Wv� �3)^�(�Z0�]�sUj:���:���̓�B�y��^8�"��ӳ9��0���Y<��k�֋����(����㥞^[[��{Ϲ����]�Zz:֚$U��іEs;����n;oǆ$���yt�U������J5N�b��Vڨ�}M�5��yֺX��w�V�L��A�Ɔ�jžj֧�n��;���x�.DN���W�?d�:�ҧ��8轙<+b�Q�8�-	�vvoo'�'ǉ+�x^)mp�B�웓��s�T��q�<I��W�C�φ��7�Y�O/jiL�o0n��;w�V�R�AM%4�v��-�4�����Q�I��I�`�6C�~��%-ˮ��UC^+��]+��,X'ϧJ(TV^�����S��h�^��x�md����exؓ����&th��ًƝ��9�=�@.u����V=�z`�H�v��#�������PN��ܬ)
�aƓo����8w����u����,�خ���aF�E����4�u+�5m�z��kB~t-$���^��ӅgD�:�0]ĳ�ʞ̸�m�ltB�v�.�ZNԩB�5##��<b��:�;��yZr5{g�-�S10�psن��H�����O��;�g����@������:�9U�B��܇7�+	�]kvZ�p��Э��b'�w(w���F���k�p�V�5�Iy]vD5��!��������pWD�"�(���~�Yx�t΋jw� �Q��m)!r)uJ"U̺���q��}�x�JS����ux��^�YtC�4ZiC6evk�
L�^��-h���\^�ߞ����[�䩀N�=Q�[Q����j����{2��F�jg֌b��.�qYU�ɝX=�l������6_+8�'o���I�J�9`u|$���_�^(%�+��1�;3�s��߾���ڎ�Ag)�%Ek0n>bR���4��c�92�6\�V�ׂ�t��Fd��_u:��wNB�/E�$fM�fӷZm��E���� 8vr�io7K���ئ��9�;��o�$�G;���+��-�cx	�
��u�fnϖw�C�����ec�^�ap�� M?�,�F��8�Y��Y]u�:��R�{�P�Γ��r:��w���lŧnm_Kh�
��PGI�����` ` C�bld�] �Fy���@�� ��{�~�j?��9r�1!	��"h�-(� �p�D H\l@	 G�11p���c�����6���!q�B�\G��A 
GM�hT�ra��3(C��%�����WKE6�cB	8L�`�T"h� �D���褀Acv)�0-�s���\�έ���9�'k/�=:�592_�� ?�D~I��G�a�m~��e��RP����.��r��K�.���ҟ8�%��gl{�H�OM��AAL�z�נw�����4�O��צ.��E�5�dU�4���K�iD`�tM�{3���|W�w�i��Q���)[����u�(�]��]{�O*G>��;���3|e�쫻;��_��3ŕ.8��P��|�y;~�5����zF�mx�>k\�J<e�T�f��^<t^[��X�m���.�,vFK��[;�k�r�.�O��X`��^ـ�(Y�<�R�W���$5�����^�9��<$N�n�q7�a�s� &E�⠼�i&F��~��V��$Y�[��Ƙ����;.�fM5��L��C����W1�Y�`���R�2��G@��}����J��Fw,�ˀ�WBի8w��mc�%��s4^y[��B�L(��<u��+³q;%cZ��5��X�\*��1v�T�f��e�3gZ�b<o�����={��qi��:]���J~ia���f2��[\�p3!Y޹#�tx讯(�el�'5O���m�N�w͘G�yq��W�kU��z�Vr���=�E���,�묫��d̈�(��O���'��кB���^�+��G`� EJ���q�<����i��颽F��+ �G6�wH��W����x֌���v/��@��C�W_�뮺�X+�S�{�6���~��H����ye<j����.���aa1֬���_�|��k�.�gq�����
�O=:o�z5G�՜=*S��1;3��f������s�EX׵ŊNp�nۏ^������颥�wҴ��Zh�a'F�/���z���{�����Ե��<$Z^8[{��|:�y��ؗQG<�zeM���C�ٔ��{=���{^��4��K���b�vV�<-�9�Wd����륧ˏ�}6�J������w����V ��f��^%V�m�ۡ+�� F��B˼�3O���.pS�nB�4y�����1��`�hAӣ�َ��+��y�y<��N�p���(XX�p�Ǐ*���9��y�9�.��5�I7y+2/����?T�k�nJ�K��Ey/�WT�dR�;˨��<�*ڔל8��/��<����͹Q�s3x9�'	�㈎����E����+w
S�6@*�DHx����)��]�;X�/N�y�XE��#�IDu�y|�,���J�X+�2^ںZ�{�>�%gt������I>��*��+&Ԇ�z�|�O:���xb��o���	de�kj��%䀐E{��~Q���=_#�IJ�sZ�k���MS�/)�'�fwٹ��>������E�}.Z�6g�Z}��G;^-�5ߜH�sjT�xԌ�ųg��虛���qv�g��-����e*�w���<-^e2���Ɋ��B�vS����'�;m{"Q4͕}q�H��� ���$��\��LzҾ���<�\�y=^y7ҐC�����÷�J[�¼֔C캛��zJ��jq�'�2��}
��t�����Jɾ���	�p���8����)Q=��u���+tP'/�}xĐ��[b�v�P�*<)�<�a��^rw܍�1��{ߢ��c��땄f�<1p�3�8|}�([V�a�\��T5�,;�y�f�j�����3����Z�W�l�G���)�	@�R�Ù#��P�I�|���Muଆp�;�v���xR/���Ь�e�>v[Q�iy}�gB<c�ED:��`�D����f�Ynr�l�J�T�,�ҹ|8l��M�9o���W.�0�����³uD�E�5���SE�Q�O�����j9���y�s��yʀ��;*u����]72�Һ��e<�x���Q��q�g��&����Y��h���&cwWI��0���?BS�0}��]yƹ�>���-��~�nrso�"��J�l�#�k�<��H,�\�rreI��+,��y,���H\8t�s���v��x�Vu���\4b
8?8�լ���f�i��gvU.�0ô�Z3�:���]��߽��]��)d����e������z���]��}+�+�:/>�3�u�kᅐK�W����꛰�3{8D�0\��t��˳�x����y�mi�j�S¥���%�]���w�Ǘcg|�໎���+�0������&fm��sY�©;齣[k�#k5c�붮	�����%J]�1ԣl�3�Ȝ��_r%%{����he�n}+��.�7;7{���6x�"Jf��x|1g������y*W�௷��
pQ��6�i��C�mO�J�޼-P� k��ؽ�o]k��O�:�ʔr\��y�
����M#ig)��C�X�M/d��,-DQG}S�8�R�������3�ל=`��B��@����j_;���[}=���|X�$�-�S�=[��q{�=$�E
�zp�	k|��	;�<^��hi�N�S]q�aG^ܴ��v�+�C�*Z�f�m-K.fj*�W�01�P��3M¦�g��F�������V�@������a�D��P��#IE�g�,37�{;���n���*�Â���uǱ�P���#Y з9mm!CUܺ|��p��=9�[SWn��d��kg��oP���j1]^�˭�hq$�6�pamx\\�R%oӆTzU���������YSsD��E�~-KQ>��>�v��]�s�u-W��Ŕo��g;��o��Y�^"V\��<"^)�\i��g������dǥi��8���1j��[[���<`�����K��y�Jz�Ƹbɯ.�������_e���ħJݹ��<�oX4iR���]3!��v�{�R�b:䜊U��z�F�ԗO�SJ�1������SIfl��8�>0�_r6:�n6�N�E�4���^k}���|�F��âE'P��<(
S(���bg��k{VmL7�h��������8='.yUgk��w.W�ɣ��n0|}2y���ݩ��z=t��{���������:�l�vc��[S��La�H��+H|v<��E���۪�m����xՒ/.[�/������-�<�)mi��Mʟ4Ь���w˫Ӽ��W/�xN8z��x�8|k�X4
�n�����o&׺��	x3�һƯ�3���Yqiu�ȣ��t0t��S�[� ���J��`= l/�H�v5�б���ۯ�DV�PF[���R��zpާZ�YH�Y�i�j1�Y�b���F���o"Y}��b�Z�8%�>쫬 3Vj��|Gm����D��B>���M%pA���K��;]�rŷM�G��r�:��)�ő0:���|ng�|��辮ǂ�\�
�I'���M\�ĭQ`�\wWRٳu�qt����۫�U�RU��dCxHD�q#.e�Z8Z�#C }k퉣���h��*j=�����1��1��IgkY�I%@	ˁ��9f��p�ƓG�����C5x���4���S=�d\��ƪ�0�nњ�JT�RU�Y�y��ޓoa+�q����\�_��WIgx�Sp{�MT����(��7ʭ�r�iS�gt��>K�z���x1J�m�Z�l���y.eξ����b'�	�q�;g���]����zt��d\�{�Ĕ1jI��Ye]3@�� �	�M٘��u���D{�c   `  k����I4@" �q�]�2[q�#	�M�6*D�L�I�yJP��R�b!�`%M����`����P52%D4 � HC�b�� 
iT�N\D���!�H@�әI�RD�L��j\ˁ��C��92�.���1!$	�@D� �E6� M�#�r�.
�@bL 
Hb@ #��%���IKh ���@AM84$&$��ػ����£6�l�x��6��o��m���$��H�ܯ��p�0���E�Qٔ��7�\��p�4^�~zx�3[mz��vD��e�ݱ��ݏ
��k�����b�ZF��]!.v�:Y�M߯�-< �7Z���i�fl�R��M�@��q��k�k��O�*��]�O�/����*Dx�r&o�<+���jN�N��]��F���
8J��"�
n�oJ�m�J�<פuyȺ.1���2E]�w�������a���b�rxe)���y9�c�z�-3��_��ƼY�r�W���ɚ�7�8�����ʶ�+�n��M���1c�:Z�d}������0޽ �����~�jJH�W�}50�L���k��s]a��O���{S^��Q�|"|���>�vOo��yÝ����x�L�ms��^D�eI��vg/���빚���ǣ��c���v`���L��۾{;�bz�5c��9�3������	(XI~�'�W!�ii�֑u���Y���{�v�o���p�%�p���"��x������_,����N�MP�1���ؽ����W��E��ܛ0��n��F�钟/Ǫ䅚hwZ�>KZb��"���v���~z3E��Eq�6U���ε��S5�>�3���SG�" �R��kI�%��أØJ��L�,Z�������O��tw_<��	abjg��{W�.4VcvTs����5��ѵ�Jc�����Nb��|n��Z\%�namz���>{�-WvzQִ���J4q疞|���Iz!�^����tψ�VFU��&`�7+��s]�z�XxV.�g����HT	�Ǟ꽜��k^=��*�S�E�sdpVFi�z�fy��^
嬕�ҌVJ�5�}���L�6i��2m��r����]����6�e��[�b�D���=7��톳%�x�����WI�ڸ��=h��Rj�Ҁs���%2����F�INE}���1��UI��T�xԌ����w9�9f�7^�"}sӽxbB�p�P�L��'j��cܹ���gZ�M1�(�B��������]�|z׌B]0��^"��>��ۯe��<4p�|�-���x׺��e�	���{��in4�i���t�+qgM9��0�cs�e�a#����:��V:@PZ)\����	�y�v+;���	�p��#�8����^:��R�7�Q�&y�%�D�z�xq{d�3�r��K��S�o��P�f�wF�v�� U$#6�U������-���S��7zsjTcwwݩl���������vXe���@�'�n^f|@a�Ä���R�q6�~k���]W7��/[Z)��Q���+��ۍ�r�����9��ah�+���S7+¡Ye��7ޗ����Զb��.��J��yL��6,��K|�-g��c��E�Qڹ�[�YY�o.�̬�=��T�y�Y��W�XUrH���k��ц�Q�a�޽�3]�_�.�N#��(��X�o��kr���'���#��m]�S�J]�Ϻ]_�]����+�a���?@f�N�~ӱF�?h�+�%�'%ֺ2(��u�gkɗ���X�ѯRR�f>��^���0�^]O���.<rv�z{�z�W+g��Z,�ш��c��&c]��V�Yfӱ`������s�ƽN��pKO=����W�K.�Ůq��|��5$W,
<*�E�Dvy;zL�����@i�v�q×c~�E5��	�u"Z»r�XM��' ^�l�<:={1�}:2Ř�'Y*{�	�v]�A]�f�-;.Sqf�͚*Z�vV��z�B���묣P�I�qG	m=qs�åKY>r�6mb%��WE7�u&�״z�@׫�������Mp'�4�S�#��r}VS�1I���ww�~��<���?��ĸo��Vē.g�I��fJS}p�rc��B
�O�e�9�aֽN,Y����Ò�P�8�K��[��=�0^����>��0�k��h�+U8�9F���\q�P���=��`E�{��w3�J��[�X��v+:I��U\��N*@���B�D�z��͊E���S[��{�]�S*��5^qv����V�I�U����ى�8IDx����aʿtq�Y�i�[>�
���˳����=����߽^?'k�T=��nڇW�Q��a�K�{YY�]t��z����a�V�(d�����36��,�����R_58�x[�6b�W����'�*���_p���B���0Yk�K���2{�x��"�B��I��.[@���}�+i��g0Շ�����J�LJ�O�
�'�����������1A��c,)�߽��uj����f�{hS�=8�~(��T��i�VE`Eo�n2����1PM��N*����g�o.�ݍeU�]7� >V�����{����κ�k�Ct���.�LW�v���^��IJ�H�&c�q�a$d"�Ŭk-��;�ɒ� �����J��������*8���'���{rpg���j�C�{K��jO3�P���)s���|)��⚂>Xs�'�`�'������[�o��ʎ�{�i���;p����2c�a3�IdNv�;��u�z�9��!�k˳8o=��s|�l��At4?_�_����y�%<��5L����Q���W)���7��=�]���'�	Fn��,2T��iD31�."��9��M�Y#��$��E$/�V��H���_�^�<������W_ݢ�)�h�y�Ӯɉ.ղwWK���^v��*c��7��� Ӿ��@�%�;g��/MOog{;j݂��^S���{�Y[;ܽ�k���y�t�˂c:�5�+�u\~w���jXUq�Z{�~ӳ7v���o(m�`�_�����A�O�C+�ul��smKܺ��.�=�TEY����+��P�8�Pwg�hΖ�<�Vd� �*V��}�%N�p+~끻�P�=W V��'DԶ�M�^��t���0i�0e)�ϝ�wc#x�ہR�H)v���,��`���{��q�Y�����v\"�`�(h����b���s~����d���峢����pT�r�=�]��EJ7�gWR�d�K������!v���_R%��ބF������ƻ�ٽ8���R���x��n:Kc�m�aGxM�(�Ȗ�:_N��Vٛ�IC��F�7���m�g���Z�8����D�3q���dl�=��o��l9ٗkf�*S�gS�T@@܄�C���˹Ys3�-�"�\d��;����k�yQmo(*-�4��:M`�ݯ`�"�1��En{�y��8'\�</�.�t��IΜ�@[���h�X�P�^7�~L䏩��m,��q��v�����Υ�\儦�˴캌~^������l�I{QWA�a�  t6���m��x���3v��    @>�ș��lD [�Shu�� " @�
i4$ !!!qr�)$@�@�@�@  �@�$ T�L��HB�@  D�1	  �-��� � H &� A����#8&  �~�2�8���\1kI�.
e���H�  �B���l@ B �!��R�m �؛\$-5ne�i��m�!T��)-2Z�LM�$�$�n_&e��Ȗ�10A-�(�e��&����#=�%f	Ze��y�O꫙I�������έ8?+O+��t�1�{{%�xχ�W8v�7L����GN��E��vt$Uf�f/0���Sm�����^�)]yz�*�0�����U����ߧ��w{Km-1�m�^a�R������l�z(��R�Q+�u>��S<�z�S�j�o�q���b�Ù��^��ۜ;����N�N�ܩ���nJ6v)qO6��n��(�u7�1_gP�d����;�n�Q�[������}�!$��R��'���nśQ2x��g]�q �f]w��e��
Ds.�#��%W\����+ӥh�'�e�Ug�79H�2r�%�Ժ�]O���\��dvv�a��/��f_���p폭xQU��S�ź����Z��y�b�>~�&x��su��dא� ���Wuq��_�w�A��x�8]K{Y۞�.zC�(���VU�0�d�/yPI�gH�78���R��T�p[�H"�3^�>����R����T�̷D_i����\_Ow(���'�.����>"�~��y��	�OD���	�[�s�9�߅)�Q:�ߜ͍��Ud	��[��ٚ�Ο����g/;�¿(#�}�������S<P��T8�J,W�w�{�ho�;���tg1;I����.iFeo"1:��qB����ZR�k��T^�������<��}��1z�{S7�y����$rcNI?�W��Q,�7���즇�@-xM\�k�<��Z}���z,(�ݬ����m?��	�;M��ns��m�TtM���'3�{ǒ�۔�B|5��8�>Fyo_t�'�ݔ�ЯNN�vE�Y���dr&�M����JvP��F����:�OI��������ī%���n��#6�����h�c�J��1�g�|���<vh�q=�ue���%e&�m����U�	�ŷ���8`����������ݟ���y&lF�;q�o�WG|�?o�}/M{՚��O�"���X�՞�Ʈw=ީ��h��]��0{��7%=rW�m>���hsS�ÃC69�Wwo-�Y޹s]�R�v�U���oX>�3}wGS��4]�!�3i?{B��6�<{�����ހ'?]%�ŏ��2�;}:ȍ����q�����gJ��;���(�|;��l2'��ς�v]@w�<�M$��*',J���fty舅�$����\��v���龷�x����BJ����zj�{�O���茧�|���}��k����ӷ8���-�/����ǝ��}��W;�Zu��<����Ydw�~��Sy�^+�����:��n�B���k>���pt��^D�e��7����E~~K��`5�Wվ�9���}JW��c�m�g�L���&���oRݗ�s$���^��B�b ^߳5%3��nG�=֗����զc�^�u��[+��]�p��i��xo˼��xc�A^N�ž�?{%��m:�IٷAM��7�)��yxk+M y�^�Q��<z���N�-C�Ӟ��S��l?_����om�+��=���o׼'�[�|�p��
�.=�7K���Q�q-�]i%lȅ u����S]!5tY�9�0����ً2)l3e�x4���$�+���W���lm�?<��g�/ϕQX`>]XU��6�u����0���j���7��3�r���{�{㉈|����8�pT�'�g�7~$��\53��9\Pz镡3�yo�P=�9����������b��~۹�\�R��9F[��nr�����\L+Ş�k���PTb[v-!a�����wwO�����J5��5�3'h��8�)߄���舍i%/���K��xx�����ߩ����\�^D4�4�vѝ���Q�	G-Wp��}��;¨��,eL|���kİ�Ӝn�.��w�������Y�E��*�y��M��_���SXZ���m�����j�5�VזS���<4=�<bƜ^뼼j���Gق�ڲKu͵3iҖ�I�R��[�pԼ�
o����n��K� ���U}I�����<ף��A��ߕ!��Vk�!�:X��.;ޙ�ʨv��&L��j�5dWk~�����v�8+�yS�-�# �F���{_=�QL*J�|&�w��
;Ց8����5u�u��؛IԴu�ke��Z�N�y��{ӻɢ�.~�gVEG>a��bg�q�*<��Ћ�4h�f���xiy!��/.326�Hݗ�sV�mM�2��*uw�v��=-6���lX�6On�E��!S4/蘑���r@����B.�9��f̛�<��1��Ӕ�m��Y�[��m�T$@�@q)�������bÐ�5 �tQ}��T`A�q�N�#�[v�y��pܵ:c�}��YS)]�%�m����� �M�u��SB���K�U�V�_µ'��n�B�.oj��F�q��PQr�\�ޢ��m;� �Ԣl�6���z��r�{/l�\s��ȶ�;�Ԭ�p-$����S�]"B6�t�)U�@(��7H���vqNgE��.0��N\�Ԟ�>�5���y�mm�6��.��Yk��(͌��,N�3��Oӹ_��k�5(�禝�&0p��p�'%���q�G���z $���i�.�����	�owXsL�Z��S3V��cѝ�][�4R�k9>��/+���%��uM+����eDU�3-։� ;G	�3=c*K�4a�  e����$�6'$y� � `{�����{w  i�9�(@���A<��A\�(�H�D����5bS5!ʲW!P�G@(r�BI����! I6�EK�1*���!�#@��I"A$̕I4J�m��I�h@�8Y!  -�m��BB  W30B��(�� �E�� E	���� ( \!�ȋLR0 �	� +��_��7rx&b��%ʜ������n7�0?��?,�Iw4���=گ��^�3�W���<�y^
��s�(��y��Vh�;�YS����������z���{y�Pg�:�YS�ʫ	皹6����[����)p�q'#����ɋ4�_�m�����C���O>��v�􉻷Y��/�יl;�C��]�g�L������B�gy��X��Eۇϭ�{#�L>�Ur~`��Mٓ~���)S1 Zc�߷ZJg��*��t�k���;5m�G�����KZ���ʇ+�����a�����ZQt��5���wZ��Y�b�͑���y���>Y�GIb�җ���2p��G<a�غ�yv>���+��צ�^�~��q�y���?.�n/�W��V^��*}��\�oY�{~�Ͱ�y��z��낻��3�d'h�瓀�C�o}zg�ئ�3SD���I?�Wԑ)PۯߴhIȼ�v����V����|l�}�g_?@�~����S�>R8x�]}S�$^�˱^}�V�N��עQז��_��@��^��~�3/�_����|�gԢ�+�P�<��v��x����{(���d�/*m���V+�uwd��4�|[6�`��=��)��kl]��.ߵ�;���"E/��U��}�h����|������_��V
F���~�$�� ��x�{�2�S�˜�?͝W�A�Ӣ���v6���;�a�0�>��T�f�T��)s��t�����A��n��~�ںֻuIv��MC���2՝�\�j�(VJw�����G��u�/|U�ު }��G�趵򞜫�oie��=�I�x{Ο�=�ޥ����c��.�g�V]�(
q�z��]��r����:��갚���Βހ}���ڒJg���q쏞�Z�e�}�r���V7����;��~��n�??��g�}Q�����VMQ���[D(�N�\Z)���Y�g=��wzδ�W~�'��_�o�&o��tY�kO�L�g{��˭�ꜯYjzt�o�9�UkL�Okp��|kѯx:�b3�u�hɫ���z7B�I�ګ�DU�u,)`���E��.@QFە#f-�a(p,���~��bI#��?rt#8l�ċ�/d/!-�6/Ƴkئ�r2���k}�'�ٳ}�I	���̯(k�W5wu�QIL�j�AQ<��W<�M?���X{�_����@�A���k���/4H���;g+�L�A�N�b#E���������?����+bl�;��<Rɻ�x-z4qsX�N�vF��I�\���j����~ L �"#u��ﲶ�7޺��,�g~���]�},G��:x
z�[�/��k��6H3�����۴��p�o��L��-�j���)n_�x��AN�/K��z�+�^gޑXܛ��&zVs�� �8�90&�F�#tљB��Ë]u�S����z���YJ=1��hj5_o�E(}O�;��>��M�EZ��9(�y��A�=�'6���J���*���U�H!= ��|�r�������O�RN#%�}֝7��x�4^�	��d�����ݭ]��]_x�T�Z@��`�	�]��ө����3����׵y��|}���,�V�N�fx���p���J���-���|�/`~�K�^�o���].ʆùf�|=�=��%RU5�%XM�+Y�+~�3��&`�J���M�����ݛQ>^��v$f�R�g��D��ؘ��%?o��	�՛G��w�B_���A��g�e^���={��(��{�T�n�*���9"w�����{ciV{���/��Ȯd���Җ���@�"���2o^�u������AGT~��/"����~ӃuW��t��ᴕ�=��Oˑ�R}��f�^]��҇e/�X��o.��g)������Y���S���X[]H�f��6�Z�R�@$ހ""5$��<��P��"�#�~�R�QY>�#�����՚]�"e��Uen}
��V5ǥ�ۤ�牀��;�y��oH�v}��}�|ɏԽ���@�2*�y��3�p+��͊�&M�>��V
����s�[l�]�������ʜq̝������}�=�ٕ��O��_���T�*����]�^	�)�\Q'k���|r��Hz��n�\鳚�9����La�U�%|3�pjWG�%����7D�O��7{l�Es�[��Z½��I0�AD�x�]eAj΍������Ώ��t0�lj4P"����Yq�{*��Әb�n�
�QT7f�;cu����T��J��=Xm=m*��k��ࢉq�-�4�̵�Y����ta�!Wv��k]�0� :�z:�p5��,���^*͉�V�wQ�T�b��.�Vē�1��z��u�4����:؁��E;��ˠ*����:̸�&��Av�.�)�6T�,��V<c��x��B�ͅ:ja޾��7�Tw�Oó�۾V�6Y?bQ_ƻ5�=��3�9]���a��S�$u���n�l=�lf�f��Y��V�K�nsU�8���6��}�0���"#+i�/t�im���]yf\��9��ztS$���̓�0��	6Ē;%%�/)��K��|lD(剗[	��z��8�pU�=��T�w�`��Ԡ.�H�<�d�j�8F#X�3�2��0уl �~C!8�@F��&�p\���   �w��� P��p���%8�d$� PO�H M@$
�Dˀ��T&�#`��P�� Si+
 %�8��y)9p�VD��%� R9h"Ѕm���l�@��$�l�$ �Cm��1��p�M�fR��� k�U2�	"J08t�5$�   >n��Y^�G��k�m�B�=Arx4l�DD%��w�7~��+�+߶b���%���A��s<2h�p�sRA+����\b�\�)�%\`Q3��}������f�؍���}u�en��Wȧ���Ξ$��^�;�ފ��>谜,�uZ�Fo��^�Rƶ=��s�De����p���1^���r]���P9^�X2�}���xGx�NZ*ķt6�4x7+x\Wen�y�V��i�ݳ;ob���*��&[� ���kI)���@"=�����]��Z���^/uMɹy��>pj��ܓ�Q��T���3ի��b!I�TB�tX{n��yw��]��0�yA����|:�n��(���w�{�h^<Z�y�W�o�c|@𽛾�*�3�e?@�����(]Z�kO�
�����3�r:�J�o��y��3��ҥ���۠\�eתd,��Ya�M�Bl� G���=��������)����sj��)y*���;o�]����ǞX��ՙ����ߜIB\��6Q�U�1�y�A��p�����Ύ�w�
��z(��Z�˴���YD6l���d
�2gH������A��M�]�H�3s��R;Ҍ�C��=��I<�׬���z����n�vV(۩�wy��[^[��}���{�uINq$�ӝ�w2jHHB3r)0��V�)Jp���,�����ϛJ����[]_��h���x��%���t��������T��쨳�L|q��(#�����?ptQ��W�|�a��*ϼ��l��m!�g#�1��o}��w]�3�Z��o<�z	Oβ�c��@���oʃcۈ"���D����3dl`�"3�(� ����r�WP!�{�2/i�W�9�N�/�UH{��읽sF��~����@��?�Ȥ�����.��{�>�On��}G�%D�wYZ(���={��U)�A��Nu�zz�e�kqӮi��?r|�7/��0�s�Iq턤KB�v,U�)!`3�̮*��^����(�}���ڳ��g�� |@ܙ����H�]�h�vh��^�a�-�{Ɠ�]7��,�v��	���`��fyWWֽ.l|'c&l�y\H!V>n��Ҥ2���Rpu7-�r8�\�.HN�G��g���:�@���{3����&�j�4nϷ����g�ѠHw�52:�~wo�x�����LX	�s�*nny���t����a�Ш���7yb�0����lp��r�V�[�xD�g��˔n����q��L�r�xu�Ǵ��wG|�w�S��_�ߐ|!��b�� }�Ȓ�W{c^��7a�2hV^�e�
M�Z��z8��N �b�� ϧZJ[��k#�g��ک���Ri�K��i�]��sҙėom��k�f�L��f�k/��_}0��7l<۹�Ҿ��ʎ�==�w�,�А�֗��M/+R�rn�ja�q�I��Q�3�|�G*��[�+yqT�|GC�w���*�+�VK��{��u�Ry;�C�G��o����MSk�w�Gw ]v �;�ptյ�V��.�[sV֑��C �5jJO���-���s�#=����.����uF{���/���#;�$�U��1t���ۯj��Vxx�o�5=�����i�5V0�g��i�p��f=�V����Ԍap�ؿ�Kxe&�ډ��sw��X7V�y����3�VKIy*a�o? 5���yh����K�_����D&�t2dcN������1G�J Zٷjr�=0v6�3wdގ����)��v������{��ު���5�C�ſ){��zv��ד;�)t@�]�~���0A�{�c6��^���Z-�g��zB2��qѩ�{�t������;7jQc�Rb��v���x^��I���K���\��=^����}!T���yZ�j/������^A4f�з�T�Z�5�V'�[���e$�8��KL��X�f^��+oS![1 Z����O��i�f���ѭ�篯���&g�ள�u�X�q�M.��8�|Q� ��W��պ[���'�kl��O���Ci�go�E[���3�{�TH�w�ٝ\�&:���w>���J�]g��4�;��o5`��$&�*>���a��)�	��Q~1ߟF������_�W�����C�		$��$� j���AP�|P��@�jO����,\6i��ٶ��Rm1_@�6>{�m�!�)m�\�־KgdP�`�S!1A@t�%t�>a�����������X� � �H2vL�7�v���1�~C�C�;�!��(�-��p�؁g�H�b�!��1�͹,i����Y\�,X9�.�]�<"� �8���oW��_x*�"� �!  �?� I�Ǳ<?�m�'B��?�O��>�>�h�zX5�B��?7ѻ���FQ��AP�~�|�����$!��`�}��%� ����y�8P��t?QE�DJ�{l^��V7��z@�p�s]>^v}�a��d�r�T a���<1/����i���|%�T l�R�we�|6(.
3��\6���r?���� � �\)�H�w�5���~�z�	�B�V	����.C�@�{D�#�l������Z>���ϓ��GO!�� ��4����S������o�c�G���u �)ʇ��W���Ǐ��d�w-��W����v�+���ϑ�ru<�T {W�E�ׇ��0#���t�h�wAb��P{�פ(�P�v � �}�* ?�?X��n��y�$�;�ۿ1�鰺�0�p����ApvYP�:�$Hx6'Z�h{2"�I�� DN��0������`b�* �����+�4�Ѓh�Bn����fL�?qq ���=Ǽ��O  �O���b,���_'����C�㠟�x�?�;G� �~��^��3���,N��OW!�x���ڃo�uSo���4~��P
����_��;�I>HU�����O�@��pǵ�l����ø9����N�:=�6;��3��c�cd���lX�)i�A�vo��+�|7���N�O��'O��jɑ��6�'g��
�=~�|�������eyla4Cߐ����ܧo#���(ϯߢ�l�ܗD��b�@���6~�`;��<'�����O.�� >C�{�D������ن���m�YKZ��I@�A�R'�'A{���.�p� F*��