BZh91AY&SY{5ݗ_�`qg���#� ����bB�           q{lF5�e�)4�ie �m["���������JF�Ֆ�j�Q[J���SV�h�6��Fح��U4d���EP��[R^mv0�U����
�"��i�F��Del-+"�%�`��%��ѬU�"�h�q��M���s)M�Ѣֻ<�
z�V̊�-� ��P��N &��2�i���Mm��ڬ���j�`%L�i��ͩbZ��[&���,��mKi���5ZLԠ%D�Û��bafj @=P  c��m�BwWh�wfqݚ>� {ů{��=v��z^����di��CU�]}4�zQ�� ;A��J[iiLR�&�f���@ ��}�����T�T��N�nR� k7K��P���= ���:�@jν���B��y���P��^pP*�o�υAN�}�Y�5�fSwu��jQ���E$ ���


7��x5�: {���5� ҝ��=�z�=�Pi�^y�P���gE<�Mj^��*�=��z� �Z[�  c���H5��lZ�ѥ����$� �χ���x�z��@��'��:�B�;� ��o3� N��G�@�5���=+T�{� ){M�C ��z ]���$5�6,)Lڵ��T�1�`���5��m�( wZ�( k���@)J`]t%�@�m���.�^�=P���r��R�:�:��`�j��8�Z�*��Qa����o ��|�SL�� ���p�5B�S�*���t ҷT()Ї]� ���� �ގU[j��k�4 �R���R�lJ�,ѓS}� ��>�  ��wР�� &=�!�� ��z �9� �t� �:p [ݸ  ��T)�+f�fԼ��@:|� ���� �4�G@�  �p��ۀ -.�@�;ˁ��]� �T��T�2��JʐK�Ҡ�=�o�F�� �� n�t ��w� z7# �� w��  �p ۥ�  s�*zŪ4j�6T�+}� {�@ �`� fs�x �X �� �  o�1` w�� 6W��  J�(P@E � ����@~�	� �i�CC@��1))R����`�F�����R�j�     �*j�(`	��LCb4���HAJ�� 	�    "LjI F�MS�ޑ��I�OI���M?������O���'+�n�^m��
������m���f
�=Ns���UUz�����z���`
*}���� �*���?Q����O������U@X��$�gM 
�L���@TE��?������LZb���m��[`��6���m�l[alHŶ�m�lضĶl�lHŶl�%�b����m�l[b��6Ŷc`F-�m�l[b[�6���m�l[b�ض�-�l؅�`F�`��l`�-�l[d`���`�-�[�%2؅1bŶ!lؔ�ش�-�[��m�[ؑ��`�ضŶ-�b����m�[ضŶ!l[`���m�����m�lb�-�l[e��-�lBض��-�a�bŶ-�m�l[`���0m�lb�ض�-�lb[Ŷ-�b�ض�-�l��1K`Ŷ�m�l`Ŷ%�m�0�!L[b[ �lb�ض�-�l�؅�m�l[b�-�lؖ�0b� �lb��6���1m�l[`�؅�-�l`�ؖŶ1��m�lb�`[��Ŷl`�-�L[`��-�m�l[6Ŷ�m�l[b�ضŶ-�����Ŷ�m�l[`��!l`F�`�ض��-�m�l`FŶ�m�l[`��lb���0b�-�l[`��li�lZ`�-�l��m�l`Sb��6���m�l`�al�-1-�l[`��6Ŷ-�m�l�b���m�l`����m�lb��6Ŷ-�m�[ض�`�-�m�lBض��l�4�@S؅�m�lBض���m��# �%�m�l[`ŶlZm��lKb� ��m�l`���[؅�`�-�[�4��1m�lض�-�lm��)��
`�-�[ �!l��1Kb�-�[�l�alB؅�`��-�[��	lBإ�b6�m��)�[�lRإ�Kb��-�[�lRؖ��4�ش���-�lKb�ض�i��LT`��P�A`([B�� ���Vب�V؉lc؀�D�(��P-�lb [R� [ �V؈��*��@�"�P-�l K`��T�QKb[B�(�P�(��@m�	l`6�F1-�lDK`�[� �� �
�D-��F0 -�l@b [ ت� [`�lQm�%�B1� ���
�[`�l@` [[`+lm�Sb+L@b�l@b [[b�[ؠ�@�lPcؠ�@�(� -���� �P-�-�c[b�lUm�lE`�l`[[b�[B�"�-��*�� ��A-��lUm�-�c�1Q�*��@��P-�!l@K`[b�`�[B��P��ض��l`F�m�l[b�ض��-�m�lضŶ-�m�lb�ضƘŦl[`�ضŶ!l�S�0K`Ķ-�`� �1�l[`� �-�`� �-��`Ŷ-�`���m�Lm�L`Ŷ-�m�[�6�b[���-�lb�-�lc��m�[ �[1m�lb�1�-�m�[؅�m�[����K`Ŷl�6��K`Ŷ!l��m�[�lb�ضŶ%�m�l`S-�L`��6Ŷ�m�l[`��LbS�6Ŷ-���@��Ty�~��
?~����^�j�δ1u��Z�Se�=�1PY��y��H�x<�{��˴�ں�r�
� 7��E��U<$٫����}�Z`MT����/62v�j����kRUŮ��na���V�+�lؠ��l���������4��b���HSg�M���C%���[��3\�	v|��ŝ��4#�I��MwM�U�ccoY���$�JL���2�ZC����M�(hV��@�\�yqM�R�
��K����NP;P-�͹&ܡݧ��b����� ���٧/F��nC��A�uX5*�a֙*��u�6*]�Y�e��#���V��է4l�)��٭�1�
)j˚ڷ�zI�vb�N)���by(����Sӵdk�=$�
KP����p��c�)�+�� ��w�E,K܋!�� �	e[�y�ʚ+Y�K���P(�ڹ�^�a�U!��AF�����v6�˒�q��/�W���n�n^�	�s��8��tjm�O>;-,{(��*��v)�.Vݪp�,zV��n��Z5 �t�!l�4���U��AۦJV��v#0���-���	��[vek6�yf�qڔ���ct�f7�;ͼC.nH���[�;@���EU��P�X�]`����R�Ҭe�e���mSE�BV$ӈ��V�*֠�gw�jhCb��͝��*�W�a�;lå��]�$C@뽱��f"�,lV��t��N�ƭMJdr@lD�CcwE�z�Mii��R��a����KC,�1ܧ�����LV�DI�re�[F=�+�7���.��'X�{��z��6������+75�*P�;:- ��f:2\�u#���d�^5n��n]�*z��B<Y�M>��ܫ�������LUj��j(E������.
���L,�ԕ��Y�����&�i�uqe)�s)�����l:Ѻ��Z)]	U��[;��Il��QA�Ul]�q���.��x;�X�UE���>t4��o��y�w`M%c�����0]8�k %���i�%K	��v����7F0��/A�0��s%Ц�em衈� #cZd8
�Jz��
�*�,�.��#�WZl�T�K�r���$�i*�����*�G.ͻF�5���B��P�b���*�Lǎ��6̭8	�Eǹ�ֻtةq�{��:2� նE)Q(#��P�#%ז�w3c	㻹v_��Z�����	X2s�)T�h�1��B�f^۽5��ȴ�Ʋ���=@�,��}�d�&ۢ<��[��*f�Xc��Oo۳l�SJX�;ɐ�㫙�S8jB�Y� ݨ��G.�D<��6�&=W��4��c�<��7��n�&���RP֬�Ah��gv�ak7Z�6�$%CoXJ~[wNTR�ᵙ���;{I�d����paQC�i�^Q!��
{&����h��*d&8�KKqZ��'74\b��ִ����Xƃ41�էA�{-k��n	�ܹ2 ��XIު�!bȌ�av�:�7�]�w��/e�i�I�s"���[w."�a� �-�nb�E^G��2���l �o2�i�c���Ǜ�FH�(u+C%
2��n�{7s.[V�*ŵ�/f1�Tlf	*��m�"�L�SoĴ
@1`V
[�jӹ�S��U�!�l![�eVl4�wi���b1[a���TWf,+rZH �kۙL^���vΝ�8T�����W^��Im�a�ql*^��{�[@�݄sE�mZf���
6��4h�07����e�)
�r0ڠ�7��Kp�Ж5($v��tE�٘�b�c�<��^��ęZ&^X9v�+�N$�K�<�]Sݷ�VU�I����];qt`�A ���,��WCr�1zܧ�h�aiYg&j�c*P7E����i�7�n�ѫ��n�n=�6��`)�l^<m䀋��'�*a��4�����k����̰�����KB�ph;���n�B�g�w%������m�/e
���-*���k�y3THM���52Z"[��c.���s*� e �۩`'	�J �3c^��{��S�YRZ�XM�)��-^�T�f5{��Ļtj�=W��g=�$bJ�GV,tú5��B�w�;����%Zn
�ֆwr]�n@�R�tl{okvD�`f���P�bl4.݋��(�n�m1f�*֪���z�f��lH¨��-��{�+i��
���1�{D��ё5�V٢��VŖ�^h�+/!���8����n$jE�2e[L�([�*���-)��Kke���Y�֪��I1JQ�`�Q��͊�oE�)[5-�kX��0��h�!�f
��q�*ʎ���2U��/)��6��nQ�q*���	qSl�EB�
MMJ[Yv(ʕ��R�5)��:�m�S�L۹���VN��
�vN�Sj��zԅj{2����2�=�a)��`�<�^�'s3��d�ܩ{����gW�RC�l�p2UjY2Й,��+�M*�Ֆe��%\Q7�U�)�)Qt*jJ�"y!� ����GH����樉p�{��r�:��5�|Z�^�pп�c��M����q����I�k5^�(T@�ٱ�&��X��a�ͳ��p!X�L��oNꩲVB�t�R=�;�C2�2j61m��ը6�Zʎhzkuj��:CV�qn���%��U�i�4����9��t�)B��Cvٙ���E[��2�̼z&|��X6-��{�Q&�0��"�0�Gh��Q&�&!�n�`��鷵n�h&�5ph�y��uD`5�n�����Ȅ�JX����l2���b��8�i����� ��^e�w@2]��Fձ��f�&��ε�dd����t�Le�R�+eӨ�[%��2'DQ[�2W�٧���m5Q�2u,�g,^�i[�r�=�,�p�*��05L�
�Z���@wln�ӚN;����!
z5�Z@�"�%wm�����*Z�vqf�#B�,���v��4^��^��pyLn�ӊ��c�+�#7�R�X��v^�5{N�]A�IC7Af;*�L���H�54�8�R�Cx��<�5�ūժ�Hh(���U`�/\�*k��۷K$N��9������`���q�3��3F��"^Jyz5�az�ۻ;�^59�j�[��Զ�0S�J���(�ް���q˘����
Tr����V,ZÀbHڨm^'�
�D��$�tQ{�.���]Nt�a]m�3e�Ib��ը�qX������"^Z��F ���"���Z��km.��vK�Gn���Fl`Ly$�\�9Y7����@rې��(8�W�5���j��z2ΔI��ҸeܼVE���5ʱ�5�29�Ɯ8��M�!�i�n����R�@����PFP% �� n�emڅӦ�@n[�aQ�`l��Ȥn���� ӎ)&�A�{X[��0���7 �&\���ۍNVlb5Enn�4��W������f���R��ܸ -��Ȟ�5������d@� TJ��Sdk�{U�qZJ�*ͤ��x
w�dE���Sq@���)D�lOԕX��)0!�q�ዕ;LB!Z�,��v���mC"��nb��Zn��ٸQ/t�N�MY~�(�VN54�O)OFh�[eӢ�N��{�-=Ɖ)��Z)ɗ����3-���J�ݽ ���Ua�r��o6������-B޳h,�$�n��R�z��,�R�ި6�E�@@��,[{V�K�-���[���U�vv��e��Mq����dpշR���w�
�6��:��pH��r�6���ȥM�9��F�fzn�~�qݕ��m�Q�V�/j�C��1��&B^�z��f��ܸ�n�:#֔��vQL�\��j�̖�,bҗ�&�8l�&����W3
�H�ca,�cie �᥻t�o�)F���).6�kfu>YalSNmY{���q7��.��Mm���1r��3u)�u(K�f�/S�--�B	qzc��Ec�MT����&6���X�j�V��*��&⤴ G�k��ĲSj��/H���"ԛR��g/][�QNVǃ�Y���J%B]��Ӑ�L�H��L;�V�[���K�mQ�(���n�@�
ܬ�D&���z��ݛz}�N�Z�4ѳ.F�Я[fD�u�O�h.��HXZ��f�	�c���-Ӣ7@�fl�)�M�:������n�F8��Vܳ��`m�1#��A�i$�{2����Ƚ���i�t �Ex�1݆wIZ6ͫ��hە�[)J׀�y�`�A+�R�AH�Y�\"�e轑;��⹖���S��r�mA`Y4%��YƳK�5P�X��PDq���6����1�VIr������m�����������)�Ƒw7,SS*E0�t�ae��k�Z�<zY��D"���bݽ9Q`OP��e�M�a�hk�����ڹ���g���B�.:�5k�׫7�q��ҹL�`Q��բ�Y�-�4�!(j��mɮ���r�E^-kwn��oAՋ6�5.c���̼ڵub�T��m��.��	�+n�.ЪW�Ǘ�4�M�fE��c4���r����N�o�M��lm�Q*�hh�W5���$ã�c�y*L�*��.��vjK�Q㩏`��Gr�f��+��B�*�t�(���8%�Q'��X#�j��6�weL���*�e�{���p�z���Od�"m����,lZLVطSF�g0���g�U<��cTE��f&�%%3kVTz��IǬᕮ��7U�0f�7b�3Z�+I�)�t2�p`�5�j�ܷJ�5�����80S.��Z�<'	���ѻ�PH�#t�"�{pV֡�	JЩPM+�E����?XS���V�2��/e՗h�z�W�j
�5�����O��oQ[;5���.f�v)�K�zR�Zf ���I;m��K[B�i�Nb�V��\��l����#1r�e��=��<L�[t.ˠ��
'��K{!P�i����:�e�@ȑ�y�#Y�׌�	�C6�������D��C^0�fd�&֫���yu&�����{�H͘,����i�׸at�
�NR���D�뻻,II���b`;���B�^d�K�x�u�d����[�wv�6���2jtB��]5!��������c��dF�� �y����e$n�Nh�Oi�@Ev��)=��D���%J��A����r8w ��`��8�U6u��n�nV�@���v�Qe5���#*�M�c¥��t���hRNT:nkv�[o6���B)�6�E�HN��h�QU�v�S&6vfzQ�l:A{&\�I�mC3	�^�1d��-@��h���],����SH;Z�a�i���Ga*���eE{�,0��&���곬k"Z�DRF;��:���cT&9m�;H-t�:��]�%&<����A�F%������VIZ���5���Ж!D6� )Rw� V��ߢ٩HRB.�N�QLFe�f����l�}�5�mZfbY�	O%�^��s9N���in�h^_An-Sע�)S�h1[7�6����D������Ř����D�tn7�IM�t�OMƎ��g ��$u��n�R�TU�⻦a7��;�5��&�z�Pˌ9��+5�#30�v��c�����	͔�j�K0�6����D�9Kq�laئ�[����V���T�R��5��+�����:ܷ�A�<:�Z�Ŕ��nʼpNmJ/oI�m�b�*M[ae)[t�ol24��c�Vi��%�5��2F{�/!�p�f|��2�s��Z���ۄ�u���6Q}&�#xu�b��AY�E�.d�TP���K*���{nz�f��ZG��f��u���rG��q��e�	H�Vٺ���Y��O�Yd�q�qG��Rq�;	�Ql�%���Ⴏ7J�غ��f�.���<��q�n�j*Q�7����}���[6ȡ��%J�æC����͝$'O��$�	D���;��47�ׯn��'��������,�n�g�L�d(�L�qp�y�eP��"��S:�e���C-H¨J��!A7CI�M�d�z\%��Pp���I$�O&�T��|e�I,�*��l�N�|Z/	�0�E���Ca���	�Ʉ�	�#,�ݒь�;K<�.�q�G�Y�
	��r&��r�d�($�M�1�!�C�R.Ē��:�D����3%�%��g��o��Xa!�ۮj�x���zV��eqk�T��	G(DD/���m(��T$.�i��9�{��%"
$�$��s0�J�M���:H��\Q�-ipW=�}	�p�^$C��	�빻d�(a0����6K��!����X^A",�;e�zq�OP�B"(d3�I��|���C�PK;f�T�$Tط��	��0��I0�(�D�Qd�J;d���)�+	�aXE���n[��,,�AT���M,8�V��:l�N'J�6�&%��\�v�*�z�+۰��.DVe�O�FO�V��P\Q7BB!���l�E+�}N����L3$aH�wK$s�$I�����v�;�:\�1Ʉ�.�4QH�[<N��o�e�8��s��t�&ᐸMf��<�I�-H�E�:�!2�F" d���	�	�Iy~a�I8I%��m��U���5\�2$AIH�+
E��'H���6��I4ot���$P�:�m��0�
2�u�8ͽ�Ͳ��+_-p�;ӽ ˧+�i$ل�	CK:@�2j%%t���w&Ks�Zt�$���.�fB��#�ﻴ#	�sOP�N��ZmGY�YT�m�r���.��Bx�YX0��lu����b��p�]��eܒK}&�|��_��G����ō��`?����;�xN0��>o��Sٿ�I$�I$�I$�I ��gHg���\u1�-�D�ō��������x8�w�8�ʷ4u)3C�Y�8Dy7�w��N���y(l<dAt�Α	~x��{e`�E.젿�`=b�>��Fg?����$A���ÎL�b���βbbo.
�ǳ��ӋO]�R�w ���k�ׄ��$V
��,�بx��ե���5˯���ol���uIt��[4��y��og��$��e����t���)�J�ΫႲ�.�u�-�[������o*�Bś�v��%�4o�_ѧ_;�jn�_T�_+��!o��3��M�x�r�v��;�ά=�c:hu�ف\���Gn�9�[8��l���fG�{�s[���ֱ/���"p�hJ�eE2�]�gjX%�+l��B|���u\*���go1�͢v��Ag�骝�7EΈ�ʸ��z%�Zk]'(�,=F�N��\ ��ÏU,��zT�C �w1��-�n�Y�pV���V�.�0T�D��p�@(���5�f}�s�,�]k2�^��<��syķuz-�	G0>y�7���s\��g����8c������N�j�C�u0�.I!�F��)�݁a�P��)��7 ��Kqަ���G|���U���:�{�Xkl9`W��Y�kOL���+�46��M��:Yc�l�8�Ἡ����Z���i3Nhᣮ�{�ow��8�Ч��=��
�&���Nףz�Z΄\�Ŧ��
<�G��ٱ�ݻV�8�[CF\�٘�uwKc7:���r�EM7܂ޣl�F��:jl�a��qr�B���TʁSsy҂�����(\v�<n���<��HGz�\4;L�E5�5ef;��4FDJ��
�&�w<"&����@�L�gu*�6P�7�M9bK�Ϯ��Kq9P!��6�I'�W9w�d=u��SvU�����;6�+�`e;}�[&��%u�jU�V]�2�%+�"�ly��0B�d���3g\�2gQ�v�� 0�8�P��ט-�B�8Oqn 7�����(T��������H���魫R֪˓rV�z�N�˥2���/L&���7�r5����2�Xsr��+9p��dH-�B�VJW³�+(�*�����J@ �T&<�xe;��X��i!E��hS��x�w�[�b�s3�C�]�b1aYԜdwױpX֫�Gc�N)�h�j�:qا�0";�k^̖$��l�-H���C�Cwe���{�#uӥ3�Zl|�{�������'�mZ_I-��<�d�M��Run)�p��|����^�=��K�vH9�l�^s��s�=��T<wp��-�[�e���q@���5s'�"|}n�Zgb�]p�t���M�mb�#zI�E���
�z7���ሴ�+ 4�:�I��������*�wV9i]`�{ڲ�<���crh]3v�>�-k�M�pg\����������`�ɮhPZq�
3M��"��]*<2�ӎ�p�{���ܬÒ�[�}�Ԛ����vD��D��r�!�59F�sk�v�&��=v�˺HӬ|d��{�{CZvl-��pSf�4E��S�����^n�ǖ���8�C�ed�	�(�?�n#*qR�]��z����52RvԸ������7C��� Y�'yP�'w@c�`����y�lbo!���
�3�饣�� �L,�üȼ���* ��udѧn��EuS3v�#`�����uX�Y�w ΂���ዌ¯(n�<�݃N;5odi��Y�]>Zt��$N]�c5�1�q�����#�/&�z���f֗,���.�&A\�[f�|鼚J��&.!Hj�:�0��ddZ�-ܻ�WKoi'��LTGf�
�;��)	[%|�mu�[�kڃQP�ܙ�Pܩ�Ý[�0F�<shW=�:��?7�[�k�vwo4���)b�M.ĵ���5y��a��oD��Qu\5�cO�f���]�����o��#We�㻼�ua�5&�kIԇ���w��bD�sS2� ��K��I�]~�S#��E��'0��sV%��^Ӈ��Y��}���K�2k��r���cKn�Co��mJ�Jv�M�ɳ�����Ϯ��/4����Y�oqa���L���u�i�.u;��3�v��x��9��TO���RmΙ�v]v��6��|�n���XT"���L��ơ��Ӏ�ꃬ+r�ЮR��|fR����ld3�M��Y�g�z�F���#��"����֡�kF�7�Yl>��B�)Z�5��n��M���4tB��I�h𫻽�MX�X rf�mf�b�cqc��'��\���h�+��T˽�_v�@ȴ�pk�95L��$$K�O;]vvL�ooWv��6���[Q������1�{.���˫��g��6_vb`��}���������0�J�N8���:I*�ه��#0N�h�oo����J/��%f;����p{�CC$B�{2,�	�1��0�+���$�"J��ҹ�S�Jf� �k۠�v�&�0+6� �:s�]���*�%
"m����Oe_k��y��U�Sg�R�{Hܳd��V��lQ���dr�\�q�]p�V��e�\[x�s�\Y�'?6�7��Jl��թ'ypp�m�P�30*{,�C0My�q.�{��Ζ�_9���;�:��ۢ�P��ޙ;\M��;��&I��v�u���C]}�^^ԝУ�#;AC�{v����es��A"V���k��y�lسîvg5Ǯ�&ʹ�JU#b������U�L]E)��Ǥ�s��!��軨�Y��wS�b�nQK3k�1Gv&^zၐ�'f_Iw*�=�\�Ei��.�����9-X��3E��ze��M!�L�X���ۗ|&�R��L:��w��,�hi+%����Ν�1};�s�Ƈ�i�,{�~M����=�=:�V$E�ɽ��\�2큍�r���/w��3��;c��t�\��v���VM��9�`�Zr��yt�3{���r�{�ۺ2�;���Â:�F�Jw=$䷥�,��$�Y���c���P�O v9���u�y	j�d�]���=I2�a�;���F�b�z��W6��&��[�	i�Uj���$/z�]�٭h�w��������#÷`�`�X�Y��B�Ȗ���5��h2�^7K��[�Ҍ���Vs�L��;��۶�5����^7W�(ߺ{Ϧ�O�lsu��m&��H�Y�	�n�hu�&�Y�m�^*�1��3�b묾�\P�&�f#��\*�r�twt�ݮ��F��f�}�I���Yr�x�ܒ�q6lt��@��X���p`��%��
�]Y&^��O���l%�=ʏL��|�T5�O�U�Z\ZN2)��vR�:u7�c[�Xa{Nϟ����=]��-�9f�wt-,�r<m�k��:()z{�4���EJ���D�*�y���z�A��
dy��̱�5#���s�K��$�fqn�=�0��>V6Z3.n�;F������7�sk�n�̔
�C�6oV�R-��W����=i3{�긧W'B:��`�[+�)c�l��ĽYd�����i���[��n�����,�flDĺ�eʂ�'�ul/I.���pn�E�7�׶2��O��IL����9oӰn����O#e����us"I��LW��E}\�f���5�����[���`�B�v�¹��&ᗽ�t�jP�zvNg:X�\��*Rٜ����)�u���U�/u��]҅�򼷴t�s�f>�:l��J�3����n����A>��U����vu1����s��.1��9���Md>瘭���-$B�׮�ǭc�q��Rnsˎx�+��K)mf��ulFܷ�Yz�\'m$kD�����\٨t\ⶸX�vK�E;GH��}��Ž���Ͱ��k��u��;n����V��kJu��x��PBe���G+u1\;��>�ob]o]���s�˹KvO@���"}k�xbq�C�w9�Y�c��˾��3_lf)��IucD��T��fA��e-�������Uh»j��N���Yj����u��߃��w���d�q��-�1P���x5�s�fѹ�k:H�f�WQ���X����]�m����r�x9V���n����7hLp�+���4U��v�ӣWJ�V�1K�{��=��܆TWص���#U�x.KmF��N�!���B��}8�
�C3#T k�ZP\��7[{M�c7N:y��8L+0�c��`h&xQ�o�Z���]�K��]�0�ʫ�Q3��K:��:��y�]u-��ѻA�<D��pu�v��ܒ��QfN�jU�hr��k_RsS>�`�b�f����r`oz���C��Nc#T[t����t�s���@�&*���-�+�s��p劵����k�vވ�k��&=,��R���\�I�y��b45����P�c*�3�Y�k� @��΄Ә�P�hס�
�Y�t�m�1Cq���B%]�\��1��r)HH=�Ѝ[�i����Ku�N�eQ�o8� 4�t��pw��]��=E+�gP�dcv��ʱ���	>9xqb�1Ko0oB��D�l����W�����_>��x2츨�7�"J���:/5b�՜�k�d��5ᝣc��qL�I;9�M�/yo3����y�*+zj{��r��Lk7�ӷ�l=2p�w^ޙ��B��\w�����r��e���}�4^�fڃS�V�y�Grl�9&�ӸV�^ Y�-�Z۫������$�M����ES"���ʛ�>��j������_i��l�.-F�ӳv�	�o�=��
�Ay�Ѡ�S���
�ɇG^�`u�z�	�����(h��y9��udoy��$����e�5�	�܆.�4oP�C��#n��)�R��b`���n�yiT��Fc�7������>�u[ji���Ɍ76\��������(�z�F��>�o5���L�qn��`�n�>�Re`]������U��9wT�s]�ywu5�:��R+	]wA��N�.�7/��5Քʸ�3:�GT�wX�����L�]�q��%�jѡ:�	�q�`��Xp�{�*�Y��X<�q�g��)V��΢-�4��q��к��u�$T���lݫz��X���g�P�F�3G 4w�()Ճ�	��,z͎�6�q��j��i�cP��FZ�r�R���a��*p��1L8',Z��X����Ond+v���+�tQ�R^�mMp�ٕck7K�OȰ⼓����w:Vڄ�fb�S���f����Ò�R�71AD>����y��:��*≇u��lc웆fKD�ZdC����.�s�fA*p�R��C�t��$3/\��M�a쮧��Q�w�0-*�עw��V��;��,q������`�������M�|e���j������vM�ϓ���MGݫ�m�x]��W���ox,(-�q�F�X�E�S��I��ں���,6�k�
}�WQ��Z��9Z8Έ��V»e��wܜ�i]�����N�eQ�he�2�Ǭ��EYX{N����soB���ѷ�X˘g`�7��F���,R�="��X��Y��U��:ɹv��U0�=p����*rΥ;����v��Un>��z9[G5����b�b�E��)����uqn���� �/�(��
���gr��ib�#�rW@�۾�gᝣ���3:i�1����*�Ղ��Uu���Uf/�f��]B��rH˛(o9%�z"���V�K.��r9²��!�ie��j��l�i�
�-����y�qb����>Ӑ���o"��2R�wԆ'݄���t %8�-�ŒR,c����ť�UNA�k���m:u�ě�!A���d}P�t�:���}��':�����T���v�s�wwI'H�U�����$�%�r��W;���w/���j(yty5�5uٻ� ,���+����C��	�(��x	b��耿�G�h���vU75���o�T�j���A��_
��*
|���ȇ����*DOyg�C.�{ .�w�M@$�kZC*�����)p�N����Dw<���Y�����y�Y��W�wC������eMV�.��-:R�����O�mi��ڧ�x��59�,'��@��.��5��9T	�<��EJ��v!���R&��T���P��+�9T�s�վr�xkڶ@Z����7�^����D���>v�� ����(���������(*w��B}�>�����y�� (�������o���Z��<�<�����|���6+��e��]r��*�#�vJ�ؖ��Ƨ�%m�tU�v�@�mnE:��*�9�q:#0���G��}��;��pA�+kt`Jkp�!"KT��Z�y	���Ф��*�K���`�.��
hP��m���-ʕ܄�xS�[&�׋E��"<FY�l�It�V]7�l�6��X�}����U2�Ph���%�ɢfXv���V�����tS���kv�u��nv;V�-ڋ��CV����ō�n�� ݏ�.�i�����k!��	�M��r'۠�S%�r}�n��5%�[�Ɉ5�J疛�΢�g�N[���9�|<�3 �2έ*+}
����a��nR�j�\}j�l�~�0n�r�n�����r�J�F_��O`�q�lOj;�+r=0�[�zv�	p*}��ݮ{�C'WD �Lɩ�(�p�q�������H���˻kd�fP2o*�UL�X{#&�v��x�]��[�:붖�1���@���:.2��1�q�9-��&n)s�M��#c�]G��,ۭ�u�Nl��w,����{\O�Iu!z�wm�[��y7֡oy��6�ۏZq�q��q�N8�8��8��i�q�x�q�q��8�8�8ノ8�8�88�8�8ノ8�8�88�8�8��8�8�8��8�8�<qƜq�q�q��q�q�q�n8�8�8�q�qǮ8�8�8��8�8������8�8��q��q��q�qێ1�q�q냎8�8��i�t�Q�ni�0R�V`H��TwN��<T�D:����6+�F�b��O�l��N�����kQ�Θ�7��s��z��r�R;��U�ve�`Mg*�*Z^�΁>���>���yr۔��:���o�F�봩	/m�{��1f9�9)��k0�ιֳ8�M�h�4j�Cz����nrbLq݃�cUe-X�� b�)�u�6V�XǤ�{�uح���"�{w�N*�p߻��z�����7��*q����F��7���\��Һa���[�Ӡ�P����"�bo�vM�{�S5f;N��SxJ��]�"�S�e�l�S0��R��2CW�n�GxT�Y!*����2����N��iNgZ�n��&���}S2�\�-�VlM�g�F��n���QP��	ҙ4hسe:���Q�Rf+��p�A� %��1r:��2��W��\Ku��{s�θ-�7N���jyf�OZD��ӕd1h��r�/d����3^	1�r�X����5��R�!��7%��,�jl����I�|���Ã$&�B��lT��^ݠi �c+�u��y���0I�������Qy:��^���4�4n�}r5M�����t�v���o�ծZ��X2�y��F��v�����8�8�8�8�q�q�|q�t�8�q�qƜq�qǎ8�N8�8��pq�q�v�8ێ8�;q�q�q�8�8�8�q�8�8�\q�q�z�q�q��qӎ8���q�N8�:q�q��q�q�v�8�q�:t���m8�8�<qƜq�q��qӎ8㎜|q�v��8�8�=��w��7�i=�G/�C7l�����Н�λ6���|��빓ra�sb*����.��L+��n�dn��[w�����Y����&fH{�UK�6��o�����H]�]7���6��&E�v��r��Q�����Rf���wdm���8ƽ7pu�>�Q�5����6 �7Fr���NԄ���"*񭼺E��S�@w�FXr�(�+�� "��5�Β#W��pX�����%ŻB��YD0ٞE�np�e^�yi�F�L����������s��Ǭ�'[�Nd�9�N0�f�m����K�wMD2� {u��T�L��3{�o���/T��Dlō����Йh9�]��+���G�n�$���W��@h��Gj�pdUӃn�-l�<����YɋoL��V]ʻf-�ٷ2������l(=Hۥ0܋u�պ�)]X�Jز�6K�2Z*��zs2i]�v��y�uV�n�yh�Ev%H= 7|�r������ڮc�mi��'V^�ҋ#a� �P�],�ҥ��5�a(��:I�����I7Veax'��y��] ��չW�1�cݻb*��(X	ZF_Q?B
�TWi���odL��_Ws=���]2V�n6���n�,L�KQǋB�+v��|���~�?Ow����<qƜv�4�8�<pq�q�q�q�q�x�8�8��q��q�q��qӎ8�8��m�q�v�6�8㏎8�n1�q�q�8�8��q��q��q�qێ1�q�z�8�4ӏ\c�8�8��i�q�q�4�8�8��:|pq�q�q�q�q���q�qǎ8ӎ8㎜�{���o����x���6�a�v#E��nc��kr�ч���b�&��qMi��V2�����<����E]����;T��PA|�Q�[aP�t�b��`�S�k�>��zA��е��(X�Z5�̷Hc�I��ܛY��Jo^]����&���_n�+4+��U�s��f9��|�����rK��ww�����:��)�u�'|*@�4���Hh�.ޒ�$V)X�'N֔V)Y����8�]n;;�$���\v;���Z�:����g>�8�e�KV�M0�K����;��bB믋�i��gIO��X4�27�!]�Y�&巧x�#S�9��r3�>�}�kj��JMͰ![���q�g��5�]��T�qKsufN��d�}�E�{�Vۭ�d:2^2�C��ygU�,E�����Q�r�f�2WN�jA=+���Z���9W��F��̚,�V}~�w���}��|�v�T�;qu$J��V����ΰ�B�ؖ���5g�<�v�ZC����y(HkT���w���6gv��D@������Ć�=Ζg+an���늤�bݼ��% R?-�̽ÑG�5�d���	ƞ�aʕ������ݽp%�oSz�=�2�V;�B쎘9Q)
��{r��K��/��b�W��W� ���vmҾ83��1�$rh�T#��q</�j8U'��I*^�!Py��.ꤜ�z�rY�g#Y���Ηq�v+�օ�4v��f΅c�gq�/(�)�#M����ΤWr���Z�vw7��\��m�u��0b�ccq��j;�Ѕ]�Pݳ�D�"6��۸���L�	�cCsB9Z���M42z�]g2:�I���=��z�iat�B�5�An�}�[�u��4%�b�QZ.t�.�;���f�@�4���<��h��{�ٜ�[[���E�[����Ͻ��]m�^�DUs\�w�J\[
�S����e	�Y@����׈n��4�_�uk/i{��U��]�]׃����-\a9�5(��)���W���伫���cXA��s���.�&���jM�'��h��`�g�b�Ҭ*p�� Q��k�Dw��EU�\@��V��h���ܥ����j�pkz��Z�;9�'p�mbªV��7��H;��_�<僛Tp�˛���f�(��u&��pÂ�Dph�p���ʌ^M�������B(i��'��w^�ȱë����O-�4������h�W�R�{!���R�h�>R�N�!U�\�u��'d���� pUo�[�ᚻ{�C(f�L�o&>�t�۶�2��G;���Q=VJW��n;���g�Q�T���N�M�D�,��;��AD�g��*�Q��%7�
8*9UM�~{*������c�� ���Ic�M����n\U
;�'��KV!Yϭ��N\����{A�Ű��e��ʴj�i�GUs\q�Zu�4�#��uO�Wf�m)�=1��/w��jF�������C k��k�a�vD51��f�i�nr�`�\����	�hN�{ίs�/۽2����ؕ�WR�=���X���C[+]�Ż�,VȮt����J��	N�瘟Ԓ#y~�	D��k�vY����Ѻ\�u��ѻի+C��eA�BU�WW�F��K�,�R�UԙK����O�~kvrެ��!���Z�C��J=�j�,�F`��ǽ淏*W�#���Vd�WHśb_�
:fјPZ}	��eCo[���4�J�z��Up�d>:�;\'u����B�7�a���yH��[��eb	S��9t���������f4�ُ���o񣷀�|E`���Gb�(�ob�A=���;�&齧I�`]�Ն$uꦖU��.�Q4�]h�ST�ٸ\6�@&��%�}W�s7å���L�/2�%�-P-ફ��b1�*�p�����G�h#/&f����.�'��֫�$�}��8� ��"�xr���f
�m��R�*�WZ`T1+e��R.�@v���6�;Vy2�����Y��V�KC*�)t�F�r�.n����\縀G�
hW+�![
��\����n텓eJu{���ڭ�Gۊ�j9z����H�18�I���W:��[,^�.ew.�q7��f��+Ud_�}J���s�����m:�BN���:d�%v�{���+sq���
*�A�W�o�R��Μ�y�F5&�5��9)Ax��V�Y�S��,�Iw00�j:43ٳ�0у�Gȭ�s��L�|�f��^�ٺ�N��l��7�L��̒!�}��ڰv��2ȕS
Xu��T�#�=U��������y�u����5��S�(�qޘ8�F�mn�m=�/-�x�,�g(��z+��~L̂<��L�,�}�{�X�dE�;`3���="uE�)��}��t�h����Gz��̠�W326ޛf��ުV�ޱ|ٹ��GY ���]�z����ZӋ:�\x:+N�+�P,⇀�D@_	&E� �eoL�`�a<����A]6'��b&m�ޫʂ`+i-�7��ypR`�/�d�33f<A��ҦD�hQ��ޙG���-�K�R�ڧL�a�k�kyi}U���Z}TV�Q�U���b�����>��)��!���z�M8%<��1��	]��!;�q9}�Uг1��$߽T��S�Җ�x;=wg��]Xz~v۹�~�ʐ��y0����ȼgb�R4��a.s�w/^�SH��~��/l��F��v��5S�u��c����B�c�ZW����T�k]��r�cF����v����!}�N��W�sɮ��Зg]l�J���ݩ>���L*�a�{G�`c�|a�X��.��f{�Z�Z�&7Ʒs)��z��嶥��E�aƐvN��t�]���.��]�0��^9�ם�HǇ���y����7H�����#}b����K���TX��%y�I��0ڐn��g;�"A)�:^K�p�7P;��>�Ώ�lǬ$R�]��Ƴ(�Xw��6K��ۉS����8�#s������S���T�0/vZ`z��@����<�{pBP��%�Yz��Oh�]Rg�ߩIgB��h4;l��V)�r�-��yͻDqC\<��Q���gUo>;ci�&��{aC~*���*=��o��"z!���Œ�f$�6�'Ld���oMfv�8�W9�k���_��ܞ�x�n��Y*�ls��K8U��Qb��l�=��	pe8%��m�E��5�)W�I�9Y��B�Ծ�W�b���tT���kB�*R=��\�l�
���i��m"_��-n!2�2<<��	�k�@�Z�䝤j�82��Ko1���}zP�K���w�;x��E�BN#3�c��Q���C;*���1�<���i�u�}	#������ ��eӚ�����u�ӳ.޵m�5��K�EZH�#�ɦ��WiUؙ=��#�r��5ц:n ��ߵ�L�l��m�v�5�O&��Gy<�h�n��9���^f�f5�X�1 DG؎^�'ۻǇ�:,,8m��*��̺��ѝ+�S��9�P��ȭ�a�{���|V2x6t2x"�8�f���A��u$�@`N�����V�[��Z#o�ȁUjiJ���/��}v�og�O.@ǲp�yZ>Wr�5��S�2i8��7jsU5o<�wWQ������z�J�A�ktb��3��lt��ֻ��Mf�8��3�)�Ti^p�Rۺ�r�ք��u̱2 C�X���,�܇+an�@4ۢ��E���2h����u&2fb����=�Zz,o��\��J�] �9؄�r3��`���Ü�Z�У��v����l<*vA�k.�R-�֕ew��($ms�K�VN���t��ٖ��2�6��;�U��2�j��u4���0{ ٢���t�3Ve���J~h��Ӿ��7:^���i\�umaʓNT�.��c*���4[u��^�.�mm��
l
�����K�*���Бs7f{��/.������n�
��3�N$���{L��z-�>�r���6.��m�gG"$�G��6j�,�5�ٺ�S��jĐT�{үNŁ�S��9���p�1����b��BX�P}���G���Sӱ�R'���ڒ�򍡎k���R�,����|GX|���^�y�쉬fީbX�xh%���ܔx��I�j�lhݥ^���ξ���01�6s�����xrד��h�� ]9���fG�r
̮�{��%��6��$����Lǌ������݀�,��֮��[�/eNI�f�HΆ��Yv�]��1��pT�i�����6��Zl��6�F^^�8�v�Z]v��嗩����<��.�|䟫=��,�����7��k���`�;�9��B�����fT�w���4r�6h��oFk_��'� C��g��_��������������Tk�ε�5*�\� ���MK��2L(Ԣh��?��i(C,kB�S����A#���) D!�#��0�	!��"�1%��K�aFZ-�"8�J!S�bI�~,��^g�4QP��Q@�.c1D�#��A��b鴬+���G�Yp�
R�I�$d�M����H4�i��n[(�|p��,�[^"�x��m�QBg��L�f#��8�mC���	O�)1@ȍ"�P�4I4	i�D��$�_IjH�3г�Q�X�Q����o����BI/�v�p��i�e�Āg��Or�F�-�{��;����݉Ì$լC��X~���]��zEIy��w,�X� �q�.�EK�c1������/�f��Z|ATp�6�Fp�B*y؁����AIֆr�����	N����m��oeC�a݂A�M���[����=8���A|�َ)N`ż��׬]-�����_C��{�$�u&T��+��;W|���*9����ô�-� tf������kR���h�<��y�\'vI�{��;��[!�:lz�<���95B_,�a��U�q7�&�Yr�&�
t��]�|әK�wko�N8$(p���ޮ��F�l�o�̚�ٽ����$Uj-܉-��v�.ERl
��WO%�u�k���.�VV�j��i���;p�wjn<oQ����q�#^�v��>�մc�;�X�+i���c��O��&U�I�K���OwbݧE"��!Ïmu�Usx�gQ%.�E�ɻ�)�~��]�D�2�4��iP��:�i�%_d�w��׼�BX|$�*.�B{����0�Y�*'F�^ބ;6�h}�ol�.��O7���g^�b��IAd5q
	"�J�rF�$J(��$��T��II8�a�J�($�h�D����e�2cb$��(2`e�@m�*6BH�i�|�eO"e�[i�2 k���!Mi�B���Z1��,�EDP�UL��Ȍ��GB3NA���a�mE!&@�@����P4�a��؄��%y�K�HQ�ЁBڸ����%5#	?�
B�����q��ILR>>����J������gʘ��H�E�Fc#�%P0(S*|[-�|�� �h$�Q���N):��׭D"A��,�#.Ԍ[-���P��@�q�RN8"d��E�θ�F�:$ρ��%� Aۉ�K���LA�B�D�>JD
�!�(�q������)2j&�y��% # �Z4�D��'͙S��L��Ҕ�	7M�H 2�(�KRz$K�HXy���+INH�$�i��(2  p#�D# $	&Q'�&HFȁ�����"�(���-�1�"%�d"@נ%�0��Qd�A���7��h����w{�󋙄H&�����@�wӎ>=q��8�8�8���N>4���^���G�q3Q�%{��G:�\ܔ��4�㦑��:�$�42c/���6=z����8�=z�ӏ�>>:=BS$ȗ�gnL���&F"I�q}<x�1z�#���|ߛ�{ߛ�q���8�=z�ӏ�>>7�$ 2��.��""�\�NH�Թ&�O�K�@�)$��G�ǝ��� P�&�`&�H��vsWwt��x�ח"a.���u�t�˖w�^�z�w'wt��xw�Λ�o<�k ]ے�V���rj�˺�뻫��5�9�u�9��x��FJ��74���r��M����w3�ѻ��u˗uh�s�V��t���H��kn�n�ur���:����w.w�y^s��;���=��.tֽy������E"@�J�T؅����RJ�h��͓�w\��:���ݜ��wv�Z/7nu���4�G�o;W��wOns�֮4\���v"N�.��N��I���Br�N�#�:�wuu.�9��������Μ��]]���r�p�<�9�s�& �����wt7z�s�˹;��'D� �IwWw\^w&���Q��u��ˮ� �̣���iJ��!��4#)q�!0��$��"(dd��	��M��	I�>��%S,�?�j����Q
�G?^=���'���y�2�hS_'�t��:�+���.j6���Y۵�)���\ii�n�*7a�!"��1i&�1Z �gŘB6�@A���yQT����Ʉ���p*Rd��5��i&In���!$01$5
�E��$���$`1�h�"�a��������W�z��nq�}���,9�F�K�6��OY���lk{{�A�Y��Nٽ��^O?^m�{à������U�r�s=O[6�O	e���[���6�`��.�ȼ�!M��J�~�Y��M�e][փ����[R�rK�$]�
���P	%\ �F�[䊗ER*�������E���^T�h�Rg�<��+H�E�d"lk�PN�34KJ�M��c��𣹋ͳ��t�01��
a�Z�Q6��vxDC3�D��ƭٺZ�z�,:v��_�!�eB�e[3�W;w��kF��Dm���Nov0i���3��|��%��^�d[�sj>٘y�g�<K��ݙ��5�U�,N�bW�e�-��ѥ]U�o�ܖ���}i��1��>nbX�&���e�z��ь�����+�d7�k�&a�N����u�f���k_��Gf�{Ʈ_S�4f^��Ņ�ƶ��g$��e�7[�q̯r�ꏵ^�ڿ��T\&����:ar<��X���`��h�gZ��5�zM��os�w���K�Ț�*�k��e�Co��մ�'s^fTM,�y��7��Ӣ,�I�R�C 0N�.��.�W��[_/t���f�J���{�K�[H�\G��d63`��,�K�H*e�q�U�j�F C���!ka(����y��^_d�^�.d[.G������w>�v�X��''3���Z�h��^^��X���L)��;9��4#��x�v�8��V*�%u�$�`H�M�Qy�*�/vZ����BE/XF��@�&k D):��!���9�eU>F�L�����a�h\ۖ�
�
b�T:�V�Rȇ�V��4�,z[H!p��M\�`�RL�i�p�S�Sx!�*�3n�P_4ֺ��>&J�k�T�)7��}�ۧS��`i�zE��c�U\n�rDݕD�씋"�m����A6X�k ���+ˮz�(<�Eץe���Ғ��Wj'��'9�)����YB������y>�e���;���D�_J�$�
�| W\��ݓAp�e���߽޸x��f1�-�e�e��n.���x�J��q����5����@� ��z�K|/��#~:.G��tD��~�����8�ej��h�����RP���f��)���#��>��X����)�Z�R���6�cm`�c�p���c�63��{������o�68>͛�_yQ�e<M-��O��t��徺ܚg�2�!�>d���Nم(��t��;V��0V�WIl�1����A���?J��C5� �\㯤z'A�R���׋�Ζ�W�X&��
2h63@���mJ�������Z����Х��T	�@L�����m�b��q���-(�)�:̂芰^ƙ��I���3{���վ�j*�2��
O���{�{˅c�0ﺮ��T"OtQ*l�&�A�FxŴڙ*�T�k��]I�/��z���=2��� PJ<�S/GdU$���U�/
�����%�;�4�lՄ����f��U�^�{}��/�f/w���p��=�*bN���1��a?	��W/�KΨ��fIIu~dsdv�Ʋ�Mo�]F�,�۶ڢ�39�m�%�����o]眜5�d'B0#1S�V�*�m���֐SJF�n*%̌���������|�{*՜��+���M�F��$RR�Bٓ�s�O4� 2ݫ�ӏ!-kv"%T^-/1�+%��7��]z/)
M�^��:Iic�Z��t��Z}qv%��q����X��a�V�̄����Ͳ�$O�nS�cjA:���~��-��n=��zD$dE�)�zwc.�Z��e-g4XRײ�vJ����R��a�P�Z�-�F/�[�lNc���2��Q�h�Q�y)ѫc�J	V�D��"��@Cd��`�G�hL-�!as�K�8�(ʲTҬ5�^�E�0�a�V�lcݴ���csinTg�l�.p�uW��5U`��>��jӘ�4�X\�/)�y�l�*ʦ1���s9^�$�?��w=���A��YZ�Ό����N��4�-��ɲ�N��<C�����c^]wg��=Ϣ�-C��4���,��:�rP\�Իq��J����4wi4�Z��uL���n��.r��1�o\�̩ջ�ڒ��G����>>�ի)u��WQ��WR��vY�:,i:�"���Ժ�"`y�4�'���,��t�]<���P�t�^m�L�y��
��=���X��&�dN���P0�j�ʲ�"���ve]�v�d��^w�T��zx�I`��A�P2i38w��v,B��׭���]^�bIY�(�=I���;xs]�>�-����t�f���?�e�X�$�Z�*�);5�lDUB�)C���\���<�N���%.]�9MG��j#!�dH��U�&VV�@���rkVX�L�B��6�+R�B8v�^��U����56ዋ�е�,�-k��L��+��*������T���U�u1�L<+�g}D�(=��4�i�@��q�AYC)8܍'�M����pMk(hҡ�v"C8�\�S�R3���T�F0pj um��SQUr����/k���,�KT�XJ=�eh/*D�8Z���5�be�[W(��>�������nf�2P�tJں���l'F&��Y��Gz���<�ڰA*�WV�ܳsv�`XcG��{�UW�>*;܀��q�5;0iԦ�q�+{l�N������Au(j'�ye^�B]����8n��7�1��|�L�]�]{̿t��v$4��D�/�}h�m�*e;�{�lv�KӀ�󁂡���Z3$�[ Q�c99�^��ۉ֬���RM�Ccw�^��nO�,�B���>�Kh$MMR�]ѝ�&U�dޱG__�j�e��y��Ia��|�sU&FB���,l	�r_�M�Ь�oaEd��m��`���Yz�+�X��֚GjNƗT�j�}+�ە�Uǔ'��Q>U�?e�ʫ�+;,L����f�G�Et�����40jƞG8˦��2H$��8)���m\2��؀ J߅n���9��/��I���r�N��v�.s�	��Ƴ;���bGX�u�;U"��5�)	P
R8Ēbq{�k���%�jieXS��o���_�C�J�[[�):�غ�xݼ�A��:KK����U뷂\�G���sY�����<��u眧;�;�d��U;�w���N�'�DW@�A��sw��;�4�����Q�ۧ9�-ꥲs�&�5(ϛ�!Y�|�lsI��Y�3&�F����xxz��z�c|�>�b���6�ݻ��u4Q�P�)��t�EB��3����Z���B�n��ÖqW4�zd#t�c4� �Niӆ�^``�4��M:M�"�j'Y�В�2EN�ۍ�u#s� ���}T�T����Ɲ�G7�EN�ݏn�J����O���җ�]w_1`0h�҉u=o=��|/���*IB�϶�����e1�Jج��M-Vl,/����DH�:��n�k���O�B̪�c'-L�կE,�>��r!ݮ픨/��L�XM��Hvy�B�Y��z��j��-�?TǼJ�O3]X�'	�A,&kʧ�U�Sg��Fk��czړC��m�I��g�=���$�H�y�W��㛛ڸ�T[t��N��WҳD?juY��n�����ůw��۾̍-^9@os�v�5L�%���|%�������>�c+4n���J��RKX�y���솘�5�jQ*D.ipp�V���y�7�� {ۆ���[D�Wk�-Wu���tۧq(VV�y̖�sv_ [	yJ��z_���X�:9��U,z���
�x��B{�U�����}�ةE�|���N���c���St��֩^�
٭x�?�9�4R�<�5몝�	!-��{�,�Y�r�虙g{��Y�U�@k
�2�ED�"jYް���)*L�	�5U�}�?=���N�����x�+<�21�����Z�ػQ[�H��o�)���!H���;#(�ek���ʺ^�Dpl�@}��y�u�|����[�U@^�"���c�{ڍ��ƹ/�ddgu}/�}�-y�f�Fy^6"k��I.��|�s1�Z�%� =Sk1�7S��xH��,V�(�ov�g�V�iHl�U�˼�X��_\މӧJN�/h5��f
�:@l�)�zv=�s����d�S2E�f�ڌ�^���7��&�`�C�`���:��6�<]�9)
q��}�}�� ���~�w�.����mq��t�7�t���8o ��N�=�:�X�;_���!K4O_^^ߎ�{}z�����y}R�թқAk���ݴ�iޑrWP���T�Os���k�+���b�7;0�	�������+-�(V.�;�]���/W=��{ڷ�M�cTV���ql��\ʱ��;MB�Z�"db,f���l��u�u�HeM��h�9%�#O��D�mǒz%
�T�����e�<�//��T� �aj%�-9Y����0�Sb���i���[EP���se��V�ؖː<ɪƔ	Y��Yf�Ä`8;뚅im�&��{ݷP�~�GZ����5�M�P̍���� ��W�w�6���e#y�]�p3ZS,��*X"�#B��pJ���Wwʶ�"����}y��t.L����͝�(���24�KC_f�����I r��Efh,Cܭ`�H��OTq��e��!���F������jW(҄^��PUp��2׹�����F�L^-�:�>�3k�t��*�-TL�[=�+�W�{Woq�ݡy	\3��+J}g5��&��J���S�.md��}��ѩfݩ3���!�ՈM緘h�ȱQ����A
�D��&��x�יڅ����E\6s�c���n}&m��{�O��l֥+<9G#Й,]�=]	�.f-t���ٯ�M���'.����g��&�r�U+��`��o�����{��M^!Tl�J(��H|@Θę�L<f��jČ�љ%9��9o�Q�Y,o�L�)�6�]ia��M�n�qV2��j�l�E���������V���B�u����F�,ܑ����$cvR����w��F��>a��� �H�|0�e ���F��e�(��/�[�ib	+K�z�/Μj���C��嵢s�(3��ج���5@�b�Z��yx�2���0&-Xٔ)^�	g��2��=��y�,��E�
23gu-�$MI5�{�(�텳Z1"g�+�����k��sʄ�󆪝�#!`:�f-��jҖ�l�5(%(�x�G��A�r��cX�t�"�����-�f��r��r��ѷ#wpF�ϳ�#��S��� {�����T�V���u�e�L��lf��dn�JiZ�l�3�9xV������o"��i߹c7v:�(�).������R�Z�rN �e��v�=�h�\Wtyaw�pz��]kAD�T{�G�B����䵋d�W1%c��wKn��p�Nw>���2k#�_Yr�_Qkw0͎dM{L*\*�N��sx��[[�N	*Z�b��8�J�̸.�w3A��'�6Z�w;j�����U��\��0<�y�t��T%��Pl�V�'Bs�$�B{�M.����Xp`��ʸ�,�E�U��yllZE��S�vk�*�^ex��:on�+G�	7u�	ת�4�s����^%�[\4���G��`��ɴ�����b�l����ps\xk��畋�"\ѽ�{	Ujm����C���L�%����.��a���T�a�Fb��Z��s2,k;	v5�2o>}���9�:�,���c\1E0��W(�
��E'3���&�V�u��	ESS��ӽ�%!��Y�5�ɇ�_�87wٜI6˙C��f&8��9A�	f�Y��Kot(�螅wt��`��坬ӯ h`F,�e{����(蛷�s\���-��[�N��ggEJ�c��wnm�����%�_7م�]a�Qd���ǚ����.��םk�Ҷ��9� *±��`F�]��JȮ����6i	(�[�Z�B�9r��V!ED��1i����D�\��L����R. ���}M�Z�YشB�͋>�+�Ծ�vg���q�Ђ�B�)c6++��45pt����� �]�0�۟Nf�VxL�K���q�&Z�g��L��H��R�=ÝA��>"A�:���:X��4�s�-S.1�nq��]�&���8>�6��`q�wS�m
\8��PJ�]:�:�X�]���w跆LͲ�E��=���;���TM��]��ݚ�Lj��k�a�QWb������WGd&��jk�]�І]6���@�����"�n��|:}�=ݚ�w1եŊu2:�׳�':��k�l��fQ�h�hެv$�,]$}����p���F�r�ON�:�A�9S!��],N���K�[ܳ q�ޫ+ޠed��M�^�57�>}�6i{}eq/�ȓ����F�C��K$,%���
��V�6�0�%�c�|�=���L����o�yr��X�о���X���F
��eꨪ��0���vE��걼L��̖pMՓ{�1�n�(�3%��V/������3�5&�:���	Ot�}ϣ��0�K���㳑Mr��E姯:�n��t�J]����[Â>���un�B�9#�;h�n���L�6#��W3�e��Y׺���ɗyx����> ��-$�~�o.�x�L�g��}�D�ή��{tMѳ´I��o���}q�q�ǏG��m;vӭjRH�	B@�	"L���w2Jb��	3��!�$��$�%;����z��N8�8��Ǐ����v���$!$f�BFa#�]���2D��ݔҁ�BȒ���$���z�����׮4���8��Ǐ���ݶ�
�n�2H��}�2�qFIH���tWݷ]�I��\��M3l(�"D��Y���]$���#/K�'�^m����w] D	c	)�.eΡ���y܏��@��1&^u\e9�09��"�up��,��C&E�B2Ȑ��/�r]�	������r4"!'�^.B�����S��o1�F	+�F4J��@��bA�9W.2�nC��X���p�G�iȈ�^5t͔C eu�A J �`(�e��$��6��מn�b�B3�d��2��To�a��[P'/P��{�7;DPgS���2�w[{��nN�)٫�ަ�d�����SC�g|�u�����@?�(y��A�θ��� ��Hl��m^hl���
�D<*���}z�l��F�Y�\Lx��_]����;r��[�E���oJ�}V��q9��W>V�.�o"Ө�0�.`oS���<�uŒ_��{�ť�G���+��`�|��F<�)J�7�eك8�A�=}Ռd�qxl�z����W��*�|��9�C���υ;����,:O������j���7��k���uE�K�6NeU��w+���y�`d�}�)�>S�>��� z��z�fq�����"X\�7���ctq)�־�3I$�0�@���eם��U�d�'��[�&�s�t�Y�	�^]�3����'9�?��	z��ɗ�"����k[`p�P���AnO~1���|)��C�O5����oh[Ty�.܀�	�:i�i�<<>`8'�}��!���*5���\H&����̸�ou�Ԕbu���t{�����e�����p��UQ4��X"��=�^�<�~��C<��	�ºO�`��z�<����Gb�CV�}��ǽ�����)��G��h�9����p��f�x.6��Q�]��/�w<Y�Vm��W��gV��z�R�D� 2ua�j�N������c�;v�(.�.�����{in���e5zn
��b����Z=	ؓ{�/���'�wk���q���	��#���q]1�;M_PU}{�wf�8�i(c(V�~�U�u3����{�ጥ�9.:��y��xwƶv��?�/�A�<}���W�w�o��;�`F��I�W�}�{޼�[�()�(���V������4B����滳6�c;�C��9)�H��F�h�Ϟ�i��Hn}��k��[�{��&�9e��#���ўaȯ����fCST�N��{����nd�z67��K�|�/�d�r���`'3L(T�+�l�W,�S�{�9�%�欦��X{���<S����;�PP�d���_\�'-W�x���P��PJ@f|P���л�w�c�{��_?���'���&?�r�-���P�3�
�}�y�4]ʡ���9���u��;�o�~��X���Tl'~��
�\Fb�*�����N�=������~��U?I�t�W{�v�E?]5����>fJ �����|���<��^ͷQ�l��\��`N/�<���� ��:aX�R��/��� ë�"��h[ }ύ�����P�T3҃�$\�C�k��^�d��x�K��;��y����z-�^��[�FD¼�;��W�{�W��Y����V�R��]~rxD�f�X�+-%� NKqW'����U�ow���5�A����[��3��s��4u���'�Ը5]� �+ޣ�'��u|���%Tಌ�,W�6�>�,*�E���:��[��_�E3��"�-^����:�=�������J��Y5m&�|(|>
��r�<�&�w|��wV��3+y:o,ŷ���Zw�W�H��!W��+��2~��ܰZ�`鱀��Ľ�D����W�P���.e��N��*-a.�Ƕ
ޚ5���3A>�PX~7����g����_?�>��� @M�}�Ҝ�� ]�t�Kc�x���q5���{���{v ����0|���Ö�1�ω����s�+�-Ix�� ��>��E��v��Oy��5<�@%4�L�^�w����
�!��K��ޔa'���8,���]٘L��Ra&���p�s����H	��K�8�C�mz �b�1��/��O���=�O?Q� ��c{�/8�BzA�rJ��L��j��Wֽe�*�Z|^����dl��1�rp�m���'�2\�5��5�����T/��N(Fx��Г�X���GmH)z!DL��kCj�8wx��@`��3!�c��>C���]�L�۝��8ϥ�\��2�mS��t[.7����5�w��'��G�[pQ��S�g���?��ƈ��U߼���9�@Q~χ���#�kh��.��� Q�c��j�����T9�+򚀈���z~P5>V|)ӳ��SHi��}pQ�Yyz�ҁ�f�EJ�ĩ���<r�2*�6��h�ພ�j� ����bl��݌�j���B�on��;~�(P�eE(@o��K�_gkx�B��+c77�I��K�55#�^���R�� n�Z�rk]�7�����dc1����y����	��
�,ϖH<����e���%�eY���<�y�8n+1]�a�s���� ��xi���n���xj���?�p�T#��F��@�[SڡR����,r�O����>�8�S����\t]�'��+}^ӥHƫ0��@\�E��V8z�l�xoal����ΚNt��C�,�0G���坃���lud��i��k@�����W<F͢��	����\�.�fH��+�!��E=�� ��'�>�	O�G�h�1�>!%�r!�6,&ԫX�h�{�"�}q�M�y�W��˜]���z^��=J�s�!�3�)�eG��u�p��������X�J��1�z�������^Yw�r��?�A�/�gˈ��� _����Ds
��Յ}�Sk��<�n[�Ko.��
��"�'�b��x_*�O��7v��%A�MA�6�50qt�y�W�W�П���ژ�,�ԉTWC����c/@��r�Bdޮ0��P�榯eU����"��c�f��I�xN?��z��2`&8@�Ο�L�}�R+R�s)z��n���u\\3��jp��X|>�&�j����fѸ9M����v��_<4�A&�!���ᮻ��D����*w}Z*��=�[��;u�ڷ�&l8J��K^4��ް�e ����!̑d���.����]<��W/�|�����0c1�o^���s�ӻ1���;w��DHJ���mn�
=��x���vݩ�-ӳ�[���$�����'�Z/D�=�-:�4�n< ��(k�6`o���z�����:����ob�{��glcu��ڍX�=�7b�^>�t�_����(�[Q�`�v26G���;�i���7���Տ`ڠY=^B.���}� ����n{��ǥ�Ĉ(��W��d���kø��\��u믳)gQkr5#��F��;v��cx�K�o�^�m���v��;���3suwK��%�Cb*�����ݻ�� ���H��:L8	����޺������_�X��aCVHA�X���Z�s�)|c��5�w�Z���Zd5B������xS������Z��в�7E	��ծ���� ��5����Ƶ=끌�*E7��,8��fS��2=2:1�T.}�E��O5����6�x`@������ò'����xP�cս[�z���à\��>�o����7a������w_�5��[��p�Zax�%�p-r�n��B���b�i������3	����"�E��ß�C�e���B�1�g_���G���$�����X:�f%`��Z��qp)IV���3n�f鼁<	�U�>[or��]h���듮+-�So'9�A$d�b� �0ʉW"�!���A�n�
���z����o?�����`:�rg�K��V��A��a]��ן?O�Y7�xOݰ%�F@@57z>�p�tO|S�y��5�x�����>:�Q�:n	O���ʈ�]~c _���;�<�*}�N����S7���x�}	��������7�y��`����	��m�L;�t�����pz�]UkN������'%�'��y\d	�8�:,��;�p�`I�>��3�7>�[�����[Gr|��7�57����L�Iw 8�����75a�4'�^�:��ż���:�Ҵݱ�J��Z0��.��h�S�c>{��:���r<�U22����x�N��X@A�}Rʂ�x���{�1Oƿz�oĀ�3>0{�<��Ė��ϭ��E��S%�_-ǧhD��`�L�O�Lڎ�t��E74�;����\�ɵ#$nOs��'���qe4uMk�p&���:-��ǝ�gA��4q�K�=�؄�<�nlLxswVHlx9j+�m<�v��j�\�w0w��Mq��x��pA��C��^����İ0[�s��!鯝^G��tk�%K��[�0��EGY�hS�u	rΞ3��e��ӛr0�Kû9c����f�VLε��ڜ�f�X�z�1�/��~�:��x�R��z�kB���5P=ڥ,�]K3o���#�l�5���tH�^<�BI�ߦ1��4ƣLe,# r��;���_��!�e���wu��Q6'e�G���j�Ň�δ��tv���z�H`��m����2&]�>5��u��}�uP��zó�mY���-�K�3s@����S����	�wTiqB�870��Wr��{6�u���K�X&�;��:Lp�f9�q����	��7�ӄ���a5�㠜�Q�,�#X�J>����<~������,�|��D��n�Ϙ^����%�K�I\�<��^D�����w��
��XSPG'
|��$�T�Zx��c�0��ɪ~�x�����>S�m�D�5�[�r O?X�T:�t6�ָ�ǎ��ǼO��otdc	Y���q����~��hn�Tk��0 n����W�����̆r{�5�סG������ŗ���dL�>�/�|v��{����݁;ӓٌ���	�1��p�=���I��I�09�v����Ũ� ������G�9�n/"�Yԏ�-��6��+�>����[r��v��-���뻽��3�M ���Y�u惟~���6�S�֊x����Sy�KR~��Q~��j�����xv-Ժ�XJ{`5����)��j�.{�Ńԫ��;���W\Qо�oz���<�ǚ�V�9�X�Mr�6����L��}M��.)��桸yFrwYWe���2i<���/D���3�:�b��S���f�W\���w5w~o�����cAcLi�$ ��w�=���ϟ�p����>6x�?0�80k���c*Ԋ���7����Г�\� ��fc��c^;� �A�=����,$8p�f�p� ���{�uȩ-��}��@߂s5��i�Q���4�m��!Kl;Cy�W�z�n���d����;��=i�!��G�ؠN���>D{�g��cD�zt�K�Z/��	�-���r]���J< -L��gO���P���N���
����Ľ�{�*�˼���������ْp+�	)K����^���C%��!��D�a����w���U��ן�z*>�F��`.���� �Gu����S�:m��}޶�O���Okr=��h ���|�|��q>x���\~`�}�kׯ������^'eh�}��ͦ��ߟ|B�<�����zo��C�z�//N4��Hq���Z�?���F3{���<�tN{�1T�nÄ���1{���u�� ���ź{v�/v�nZfR���{���!y����z~Etcoo[c-.��^cu��� L�F����9�%�3������z���Mn�_�8�����cÙ�����T�����L\�+2�ks|��P�ͬ\9���m��\��?s�{EZ�&�7 T�����3�HW��A�&�f(c�k �-��{OLH��[�8�D8/����-�əe�>T����1�������ç��I�S��#cHƘ�EX �U���������|Bjr�h@���k��/ɽ�|b���P���v�c��s�C\@N.uFʀ�;�m�������,t=7��|T��I��O��c�O'�/�]��30mw�L�9�4�ʱ�� �`y�.���G5�Ǉ6ȳ"U���r<���Q|�:d�C����	~h�'��^��g�1�pǻ�㆟�� �/�G�C��� �����i�M~΂��@=l[�|6�F>lK�����;��I=����;ܽA��� g� �����8T��u��+Fj�mx� �t�K� ��9?��m�A���g�L�H�S�����L����T�`t���_Ne�}5�w�2逞�Cy�S�#Ӯ��շ>�������8?'�,s��~��ۈZ�X�x�t�\f��z�&߶���+���ú��<@�b��[��Y�:&Wvd,.�x	1���s���,� s�}X|͈���c�'�n)����N��K��)ǐʻ��3Wv�G_�����bY�`�hB�3�7s����zW���0�yJ��3P�<�AW!����:�5Ϝn5���֐��(�/y���c�;kמּ�<Яyq�{}��P�fs��[���V೏����՚���G�p�Crma��p��z3��08@����3�]ܸ�O�p������cJ<�Ǧ�Ŗ�D�O��* F��
hh��Ȁ�h���6�ب�j60Q@h��ϯ���������������W����T5���$?� _�����cϕhg�}@��lO�]�S?'��w��K�ip(1F)�2G'��#���X�����S���,?'b���m��E�GQ�U���D��I�x�h��*�}�x2�y��"y��:�3����D��1pXp�\0�BE�Ud�_�{�o	����{#d		�1,��P�/O*C���W�� �����%�]����m�?�� �Rc��Gc��s$����yۻ�Kq�\3[����ゲ{�;�[+[#Q~� e�S�t��@�pe5í��Ws�Qˬ1�M�[R×&{�(��/~N���k�T��'��c�$}=9���̬Lpe7��\�nAn�����6\��n��E�G�'���������|�ћo	J��E��t3Ɛ��D<77��LKm�'�����Z�%��� V>��D��?����o�S�Ljc���C�~���߻0��f��љ���k�/�2�a�2��I��as��d���Ey����exl[�y�]�{��Wa ����׳w/�y��K��>zJ�Z��l�k���k��ԘP,"/��̃�0N��B#u���o!��ӛ���bcn�q}1������.��GVd�QdYƟva�+n�{L��֞�/�F�r���f\��,K�q����˦�saeb�z);��WPg�<��3���'n5Cd�Y��&�r䣎��S+]�Tn�̲�;gEʻ�}�FJ�ŭ֛(V���Sf���q߈`�y����U��lL����Ww!B�RJ�5�>��3�[ڻ�%�O��%�8]�w��b=�r�U�85􏲳3S7��r�z$��[;��f��9�rܽ������#e.k�*	̊�ꨕ�����Y0��:�3����[�6<���.n�̷��_h��O#�&\�Z��$O�`T���}F��3���r�=yBc7�Q�/���L��&��	:%]�*�H��)\g_����ز1U�b�sm����Ӿ�H�|ww`^���eL7ϸSj~n���q��F�����Q-/���噥�}�a�f=
�WF�:ҁ�,2�lg@�5X�L����n!ɖ+i޸W\�.|B�"��n(�8P��&۫-U�<�֠�!�b�{)p�Z[��Ә3\���f��Ѽ7�Q�!fÒJ�5�b��M��9n(�/��|^�n���5}hܼaA�LEb����(��F �Z���KN�:�wT�$"��]����vR�:��L��p"�D&����DV�׻3�O#���8��Oic��3���
,&v�DԳ��[�b���ͦh�:�PW�Mwe�hf#,Fjo-ɋ�f�@$LVo����.����Cr�zI�b�G*kݝ��<��x1?��BЦ�&N�a[r+�#����zrE--�'I�M�H�{�<�3����b�<��K�] Z��X����Hws�|fIk�����X��wg�(w��W"��Ǐm��E���Pjoh|�;�pRZ�l�����3Z`+՜�ԛ�y�Z�dkϧrE��y�|p^�gbN ^T��ǂ���H�㭝�ع�u��,Jto�.�����l�qo�(��d���KI��[�ai�.��P'9I{���N�zAV���Յ�}6��6�_]��xn�V3*4�a�L�m�؋���7:�!�F���1vL�^-�q�g:�-��qɻ���ĢJe�u)5�s�΃4E�[�S�K0skF��:��#�i�J���8�O�Q���S�W��$�^��JR� �����mǏ)�+�ӻC�
�q������P��ܕ��S����8�{j�%&��(��o��n�x���;���9�`�5<NCg�:7[m$;4tK���}}��W�"�hT�Qz�����vMKy��:�$��HF2I/��$3(�۴̂,I�����������n�^���?___\z������n�7��љb @�a$��s#"A4i�/�� ��f%~o{���7���w�������ׯ^�q��۷n��%�L4b1!�ﮚ6P$1��y�D/]ٗ�v1��UQRHFCO__]�|x�덾����������v�a F!5*�!1��i2DM}������	���3��إ@�1C�t�!$|n%J(�ι]���"(ɒO�N��22����!�Z�� O]�����DE(Y {�d�)3�on(��tѢ&� ��
h"%
b�&4�A����)'���H�Q�۹q��J*2FFJd���2"�DS3H�
2e6-(h"�2T3��#�6�M�נPHK�@�Q��%�����h�R��() �(��%��)� B4! �����7y��vtƊ��#���<)v��p�RSt�_kŻ���Ӊn4�,�ZO`9�����x7r�FE(RF8A)�RM8C �L#.z2����I�C�ČHl�T�h�א�)�((���P%�LM�~�7����Q TT�x���8|�L�[��!7O��U�U�h�*4�
hiU���Z����/����^�/������˱P��RY��5+��M�Y9�����$��]���@}������$����Yk�D	�PS kH/�����Sg�w��xmok*m+���
����	�˞��۟-@͸�-�,��>إE�l6�V֚{^ì��]�&� 4���w��z^t�;]��H�D¿d��M�^��lx,РL)�Xm�mu�[�Z�h��x�웁�'���$�W�
���y��B���LLv�zk�W�<v�3�ހ�޻
J��� �V�^�^���I8��B�/�>O�<倊xY�q�@���5�����ɩJ�H�ٕ��Odd7xw�ئ�u�2�=�5.�����}���4���}��|� �ܗ{2a�L�E���02�v�p��	���9�S�-M��'����Fq�9�.b���Qp�f�"�eww�L�.'�S���Jz	�M��2#C+{a0
��P���,/�䭨��z�k�w�7	������.�[I� ,���y��Am}�>�q�DTscO�#���<�u�^��1��ݽuV�Iy�05�q]�xn=43�����?�à�"�X��Y����ʻ�os�a,g��p@��r���q�N�SV�^vk�9&�� ��ǘO{��ӱ���ٜ���ÄS���� \CGȎkؿ@����*/¾a��Y�-�㒮�0���9��4_ѝ�e�UH^���]�i�1������x�(������B�<� �"'��7�w�Ӟ��m���9��c"�����.�b��V?��Q�"����ɵg9*��F���u#���4�JSO�T�S�a(��?☎՞���
���w���pam~��ĲS=�Ө*���N�B$��i�,��_H��y��kff��,������~�t�#�u��in#��OX�Xc��K=��[���[�L��p(�|T�K�7��%���Xj{`5�ڄ�cY��;�`��n�������ߦ06�WQ�)�k��?'�`率���4�2�zi�'�[d��[s���0j켤����Q���Q9�mԞ�O��s��;��b���쾖�����޶�~�*�z�i�ɤ3�!�Bp� ��De��f\�d:�)�m^NJ��{����ZµD��P�|�.TxB�ʁ�l��y��tx7����{i�x�M<^]uui-����o$av��^����J�e�B���x��420Ԟ�2�fr�z�����B8��E�|�5����E�"�ێ�y\�!Z�y�\e�m��m�D��tf	{�{�M*�CL�p�BfGG7�˰�=�jv��&����²�U��١����A#ܯ5K/S�0]Դ1͍����wX�]0����$��/�K��+�Y��W3����gT�*,�xx��!�
hh)����*�H���q�Q�)�s`!2��K=��8?'"�i8%�����l��ej���q� m3�ebf���n�Y��� �P�E|�B������ۺ�W�i� s_�B��vP�g~�{�z��OL~��*�e��3�@Y��!��~^�iV֍����o�,���n���Fw�/�7�m��t��#��ԕ�l�����*x�2��������D�ˑ^���+��,ჳ������P=� �Ĳv�5mxt�g�������lN,y�&9��0im��?���A;���C����nGs�1\���zc�ɻ�^ ����¹���tngLo&�J鍧H�����w������~�j`&l���>��+� =|���/���� ި��OzZw���s�^�~`����妜L3��渍l��B�.�/��y�f�Vf;��'��<�p�\��/@�ɥ�
܏��`g�?4��y�s�~����������<sKo��L���t$�[����]b�����`�A�A�y�m~n�Xe�#���QV~�����)@�9�MM��`��Y1����b�y�+[X��:^�-	N�Զ�sx� P<Ŋemc˸i��Jܤ��z9��9��`��t0�˕�Mą7{Z��z�p<�
�g�<�7�z(>?�R�EhiE��������~���;��ul�E�y�Ɣ ff��J���	�3����f}��}�V�}Y;P�Ʃ��Z�M����U�J�9}���͵�0����?C��I*x;�����(�{R���*��F��û�uہ�@���+�U Zx����g2�����N���$����n��;�4Tg6�"�{�DT:�� CG��,C�n�Kս,�e]��l�e�CT��1{��]�b���ǥ;���M��i�'�*���>0·/�&zzr�Z�X��!9�Oy�Ӛ��:�87W�W��sX�F��綦tA�N�aŵ���w��?3M�n�uD�얙�k���2��Ĉ��s����<%5�3����v��\�;�G��F2�����3~:�䙛\�2a��EX���<0�X�\v�kC�h.(a�d�r�f�/O_�����C^���q�u�%��_>Uu*�'���ฺ_ИH���qN����̓�xO�wH���U�l�Z���~���,([�A����p�Ǡ'�#�C��*5�:}pK��Ws�Q�u��*-�=,���[}��;.�:S�3Q��v��H�7��\{k�׳�S=�o����#���A������pզs��-���L�&`�E̝|l�\�#9Yκ���tmr�―>Øpy)�*e��Ʀ��� N?CH�M*44
�$@����U�%Ϛ5ɭV�tW=�똹w��6�h��%0]�<加ިɼ�8I��Ù��#�b�G�C��^�!�n)�8}��y����4b�xG�cT����8��g�4Bx�#4�A0������s�N%��\�X�:�]JVGKO�B��S��ځ�C�wA.;���l�;n���\���D��9�?Z<�� E>��SW���o�-vvW8���7��=�Fy��Lڊ��j�>X_~.?��?|��2˼��D�`�m�v���%���g��LM
��7�=}�����2�S xvL>9�5]�x)j��r	`���3�a��,팓�۟$[�H���q��%�4�E&Rz�p��A$�n��M!=q�� `��с@���sw���r�
��3�؉ٕ.��՘�]�'{=����:~�|��ڭVT�P����
���r���Z��R�he��it�F�1˸n�x_%B(��p+ˠpi�!���8�+�]��K���fAN�5��4���&��7�>�kb��͝��3�p7r��/fۨ����v�3�`̦v��l0ɱ"��Be޳XN�_.ԧ tx5\��`>�}���st�Yķ���m��ro��Czm"�W1Ɩ�5Ԅ��Ƀ���&n�pM�����k�J��[��s<��+{�_�} �߃J�M"�44�"_��=3fk���G��_�{����-��k[n:	ͨ�ua+�gNm�`��Ɨ"إ��A5�3>��	�`��2r�����L���oA�����*��W4(�}ˑZ�T%t=���i�`[�o{kZ��!����&�{����)�C��"|Q�ǹp���+�0w�Q3�2���ޚ|Ԥ���-�-��e�C�8�>_|�~}�s�8[���w�G�cм8��srg����EW�;��P���zw�xa����0�v�ͱ�{��������%��%��RZw*O:O-��k�����6�3Eكkߝ韴v)i�����e6�(�/3-��=8�9��H�����,���>�rs��ʀ�T�8w�@c�׍.O\��)�ֻN��:va|Bg�Dm/B^=*:�H'#S�Ժ�
�2[��]k�Z�݌��y��w�37CŚK�~@��a������1��"��IN)#<^�놊�%����2�E�(�+pw��a v��P/ld�`C����k���"��EI`����N*��4��h)]� /)�ʚ J^ެ:3n�۝��r\΋�Jsj��=^S^c�Ӛ���~�����[s�Z�-�pcb��0��A$���{�Y��&���ɓW�t� ��Çg!z�KF�����&���k������iDi��C��p ���r���Y�Ӽk�����>f����Jz�Cg���9��R�@��2���2��vt�� ���f�7��(i�研3,t��<S��2���חx��.��N[�ܲ~��V9c�F�[��e��.�� $������Q���P� ���׊�A����7p��5P����I��ZŽ�]�/��ܮv|�T53%\�6U�N�/�ѽA��Gږw�j�G���e�4?���!}�c̕�0Y�=�}�W�C(<vb`�h�j����/�x��AW�������u�]ۢ���.��e5C�O>���ޱ��$��/����C��>����t�n���g�Х�3��bf
O֙��0|�7<���/ɅR 7A��f�0.���ލi�$�{LO?_t��#���[�fً|��~y�Jtj�{b��ƹߦ��}��{{#q����Ϥ˂Վ,p�>��=U�����{���C�W0`�q�w1�4�xu�;�^dk�G� c<�Bc�|۞{������u�o&�LR~a|�y?`/�C�P0;�U���GtU��2��,�wb�f����L� ���$^�����Hh�y<2��}Y2�U�@:��;�tx��;>�e��@ U!����ם	�m˹��ʲ��Y5h�S��q�Km]N��W�tT\�[j�6;������sk3l� �����F�Dw�����q쇶�`��١�!G���m��Ͷ`BÕ��l�0�Q|囕�ꍶ�~��ʚ����z�9t�~j�Yk���8�������x����)j��)1Ǔ��O��I׀î��=s̢�u/3%_/aܫ���u�G?0�-j��S�^�$��r����Dn�P��h0���ǧ�����pL��M��p��!p#�9N�5�d��M�c{Ǚ>�vj/K=�fM�;�.�~*}:��Ҷ�O�z�u��=�9}'����૗�|s�/�|��6��>�����$@9D׎��-��y臨�g�9�z� ���Y�������R��=6��s��.Cl�U�v�nץ'H8W���k�cE��m�<�Þ�?��a��y2΂	yO��|�&~�3-Oٓʮ��Bs��i�nr����V�P���k�w����� �׿:�V��*����|��3��Ƨҝ��\�zʹ�Ġ��E���.&����^�a�]�k|�~ٜ硏l��$ń,�?~O��f��XGZ�H� U��3�T��[ FٍV�h����Z��A���|n�M��N+�V����cX}�#�aɐ�>k{�8:�2؛=gb� �ү�U]wYZ�I�;ee�v�:'Q��xa}��y��ny�oZ���Px�
�44����	DD3/���{�f���"�W׏�=�nj�a�:۴�A6T��9��J$�G�b��=lB��P�j����7w���������o��o㨀,o�H|���~O�o�D���C���ɸ���d\W�Ĳ.�D�)�B�ͽ�<R��#Tɘژ����q|>V�!_�����cD�Ǘ��I��"S�t	n�ԥ���{M�b�#2D����1��-�;�L9�Q�:nx�&�{���f�JzJ�|P�Jc!�x�vvq�[i��"�}`q�a~/iF�m=�ÂP�sl9��Ӵݭ�*Q�:)��u7������;�1�g���OkQ�a �2{��+��qb�_��	q�-��tF�ןz��^�>�~��CqP��E�ڑ����K�u���̤�O;,�>�7��+/���_���`�/�Z��D������ݒՄ�s������S0/��V;�W�w�V�t[Z����>0�C�y�;)�sѻ�j��"��Ja��4���*��߂���Bn2c��ǈn���O)pT!��!���!��|nOBk���X�n�O����^=�	J>� B��.�ј�'��}�`�����ߛ�x�.��� �zr���lݫ��x����c2^؄ ��>��8T���Q�6�a�[�7�+;(�w���C����{K��) �^km�TkV��T�L���x�Ҡ�CB�M ���w�v������*�ެnb�؞���c�<Y����nn_�w`��^��m���wyF�o=���L ɫ�C0�Z���sdK��z2H����WPXn�f�X�z�P�')ٝ���<y��^�%;z��pi�Ɲ�=���y����3P��:}!�<���^c�^m��0"Ã��{��O��E5<��d�ˮx5w)7�m�`[?=E۫�j�y0��[`�Č�ܥ���?s�=��
�����G5�{r���$f��d��>��#(q��]8�t�H��� X���\
~�ni�Ɓ�+Ν�a�˛j�ޤ�;�{����pځ]7E������P���T�-�xBo@�R.��*c��n�iG�m&�O0��Kn?��sc�P�ҹ�؍�a;�m^3��m^��p�y�d�c�Z���������!����JdY�n\�Es� ��.�t����q�<��Uj�}�[x�d��}����'q"���m�:�&��+]'����`sO�S����p���>���գOE���Utʵ�l�1o�Plj�]��rPz䓖��0W-<Q�W����[���ŹcT�k0
S�h��Ss+��2�{u�FmZv;0L���:Y̽�;XE\��p�}�dP2��su^��:�Ψ; !�=��$���溹
m�n����b�'p[�{4��gd�j�/4(���N,f��2=e�P"hG��7nfdHT,кp�N1K���tp�q�Sgi�L�. y��v��5.CF-bN�k��e.7��ul[�U=gl�r��O�x �	i�I]���pʊ�)ҍ8{����2���,��T������^>ne�)5t)IN'e��x�J=�;��gS�3�o.D�W�tK�E{��Ò�N�|M�v�Ā4��BL�����,o���ǘ���r�� ��N'�|���c�ʛ����5���1�2��X���b�r�ķ
�y�u-��8X[uv�1��A/xK�X��=�����u�	K��L�^��q߶k{N�X<�5�G�_��<��V[}�:�5�x=�s�;�[�	��Boa�-��K��%Z������Ἦ���d��%�UN��̝��$��R�����o~�ь��*X6�BҊ���&�G7C��j��yM�ӱ�wy�N�wg�%�2�Q�7 A뤱*R�2<
8���  �b�%�e��!�eBDB$^�kQ��VX�b�0��Y�D���yr���A�fq�_��ڰ2����t��l�Ô,�ɍ�gl�����W �?�h��-�w__�W��ch�T� ��@Zb�[�S͗|�R�e��R�
���U��i�Wb���m'��oiu��;��sɘ��;��y)��Ḙ�qX�A�I�y{ܬ��^��^�$P�w-�a;�;)�6Ž{�0�LLˉf��٩ˤ�V<w5b��cf�'i^^�J�f4W�Ys�vP�]f4�;Y�6�:������TV�`�3��%-�W9��tz���R�y��+GU�E��{��dc��v�U��:6+��V�q^�@TSwuN3�}qo��s+U�G�� ��Z�ʆ	d�!G�Ѹ�݁�wfv̔�����h�9L\��e�n�_r�&���\%<I�e��3��c��L20{L����r,���Q�h�r�#p[�9�IstD��whA�=����{���Mi�ԕ��?"�"V=�)K���Ӛlh�`0V��tk���q�k@�[�	��^&�6
�y��3�w�E,�cl�LPrk�ٴݵԪk|��u��ݻ�qu���"���B{6���8��6�)��	�vh|"�j+�lw_V�Z���u��秳߷�������f�qQ�"�V�����۲4I��&�[��.���j�^�x���ǯ��㏯��8��o����|��E�e}�ݘS�5j�r02�$���d���G����z��Ǯ8��q��q���n�,��H�&
���RE	}wY΍(����)I�$��o����<x��8�>��:}}v��`\��h�F2!"1�������� &�Ha�TʃQQ���&��v5�u����J��o-K���0�<�`����w��\&$�B)~|�#(�F"�L�D�D�
���%AE&.k���5���|�y�c Q2��W��L�&H���_;](����	^�
2��_�]nW#j4i���{n����2TW�}����X2�Z��I�^�A�l�{m����(fE��/�������8�8�r�'s�n����:o��/\ԟ`��D���R�P9��{�����ʦO�����1���ṳ/�I9<�w�%�{us��ΙG����
Jw���X��:�D�;����fo1��Ȉ�^������S�K��W���������t8f�ܽ���YgL�C�P ���G�0r�(�U�1�ڑ]^1%8�Y�.,l�?E�	�e]��S�\���	[S���`�81�(��G�|�_�$��ݹ�%P����|�
 �0��#xs�Vł��Ӵ���ADҞ�:��7�����WFl��z�t�K8	�l/"�z�ٮ>q`�O^J�=$�1�
�"-��p-�>�;��Qm�Ջ�\M,u��������S�
QlU����>=��͜�$�����o�-5�Fra3{��}
���Ϲ�P����1���wJ�Y�VXm'���-<�B��5L��0��d2T�3�Ϲ{���-|k���V�����ՠ���2F!џ}��	�a�Q�]n��oPcǮ��r�68|ض.b��������Ŗ,|��`r�+?}��:�v�f��i��XJm����gG�w��g�zA�c6�[.��.9 �����J��tc��8ۚ�9�)��b+����h�1�,q�.7è\E�&��$��;��8A�Mq��g_MK�ۓUF$�����w1�w��S�B�	��~ q�PJhiQ)��@��\��]ͽ��9p��kd&�Α<�O-��XP��I�~�G�gG�C���dέ��x�mǷ�VG�iOmϚ'������O�|~+頓���};�VW�R��t}6�5B'�8P#Y٘?nN��L�@��Dџo��z�h/˟��q�r�aNbˉ~���&&s���l��ra�K� �����!�1����������yT�~�^)��;�T�v3U�ϻ��i�������:�TX�D��ǂ�Ƈ�k�����ٍ�:4�z3<*�9��F��vc�Ô&U��JZ�8���e��?64��udf�?��+�A*x0~�����~�Mg�vvw�Ǻ��_F�EwP%�v@,�=Q��t�����\�	L��K�-���wF�G;� C.�T�P���t$�NWd�����mỾ���0��ɞ�G�t땃�~�;c�L;1����=��6�^7�l>�w�%%��	�94!ۦV9���u��>�O��2�p�;�?�2~��-o-��>��s�hQP&��@h�5���e;��+eR��69���w��'g�wx=���^t�����Z� ^<��
հ]Z0K��	g�V�&ԧ�Y�Mp�c:��p=��u�wʁ�Nw�f=�՝҆�	}��v�p�ͷV�U�rj�����ҠSCJM
��Eރ���_�w[e�No]��.��(R�\8�����mdY�����tI��}����4_&��.!�__��
��N'��3��z���X����	tIr����VG�;q|��w
+ԩ�g��)x~�P�_��FX�����5ݘ4g	�S�'U�B��|M^�]�
�������Q�����8�]�/z8��O�-�v��Ō1��~��6Ú�w8MA�w��6�_Y�E���p8�ҭXlM�����5I���	7>������� x\C{�>7a�����]�u�y�zޭ�=c�4'��������8t
���� $�}����G��@��0ĲOes��h�	�B��y�"��z��/�"��[��r������!u����"�X�)����y�9��qN��oP��2�js�~jg��E��A�r.�������F��􏠷܄y7�Y��٣L�!*"wfeك�����;�1������R`��G�s��#���1ͷ0Ck�z�6-���n��)W�!�r�7!2�����ct��ڳ�C]0�UC�9K[�.,����U5M8	��D�����V�יt-�Tim-ǳi��P?|k�w��x�`}i.� ��u��̅bq�������ti�vq�>�{������әnr+o�����r�;+�GU�d�sG�o��w/�_�{�0� ��4�CH44�!�3��s�+�|�ߝ9G�����J^�egU
�S��W�C���K�taz��;ߣ�c��4����u�V��p�`��针���v7h��3���d����yUH�)�q���gYzâw;qa�A�>��?SЗ����[{��e0�	��̵�g��,���H}�I�(����� �i�"�C�3�08gBkL8E�\Q�r3%'�pfw���.�/*��l�NWq1�û�7��C����p~U��L���,`��Z6�fn�;�x�I��̭ܛ�K��F'���C&ԡ�@:"���ضs�!߃l�pY�(�N�������Hð��y�ݭ�9�\�c6R~�|x˴�ƾz/6��!��r��
$Dt�N]���'�"#)�����O-z;��(^��K�t5�!�b���Y��"���7����aO���K���@S��z��y���rOB�	e˓"��(Dm�YnFI�N_0}q��,���.��_Z����<�*,?-iĸ�������B=���C�T6֦�$��o�p�q�tm�A��W5�h��+>���vE� �33zg!�"�"=5Ӯ/�����pt#^�'��7���lz��쮄��s�<}f�(ƇXC'C�R��>t32�˓W���{��4�MM*-k�����{�w2�7[�o�R���[G�j'�9/m���5��R.��sϭ�w�����[���n�v�mn�G2N_}������]>�w�٦�\�ֵR�o@jm��p�2K�d�˨;M�gPj�cZ�=B��z��K�M�	���U�A�/N�o'2��j��a>X���fn�5&��'� �y	�2�FKHܩ<���i�?kݼ�7}�h���@wRGT��al�h,��!?}h��f����u�H�L�j|$���(���Z��r;�2��!��3��mscJvø�0���C��p�K����^� ��)��K�0����f�-g�<��=�h���=����x���Xv����3���Ӓ_�`�+bN��eNU�7�3��("tn�ӎ��D�{�=��Afi[S�E팘3!�g�{(��`;L��~\0��:U٢	�4NE_�&㫨+�SZ�yz|(ؕ@��	�'�ζ5{B���Y���c��ޅ�c���m �}�R�S�3U����'���󺇤�-,��hNr�dѳ_����6ѣ���:�ɻa�e��eOڳ����,N�[=��B�`�"t�^v��ٱ ���3^C�A�}���+!d�ʐ���A�/�t������S���#����
�۝����Ct�[��1�'p��xb���g��ihihi=�^��3ߝ�U_o�/��x�/��B�Gc��`Q��@]^:���y�
R�]������acqGSp�xe@�fp��28E��.;������1�]�O�� ����\�R�f�d��
c�͞��r�5�S��c��՞��."��W��}AFH���S��'YI��_�5��`ǅ���%+={6q���*k�?�9�v�y休�ahnk��S�8���c�O	MhǇ7u������ǫz����@���2ױJrKŽSk�-{��(��z`M�3�E�Ϝ$���~#�Sj�]B�ѳ����ǎw�+v�TvËÙ�Օ���Ŷ7̘	��c�3�y:,�˟��w*�𺅑���#��tf�o���˘/�,@P-ߘc\>�\�0;�O'b���O'���ݻ<�]����l+$W�)Z骢�{h�_���;Q��˞�����	�=F�muO���wo�_�E�BeC��r����}��`����"5��?*�i�2���d�������&J���zY;M��Qwi�h��rT���Yw ��U��u��(T�
���s���E����:7,���5���Z��p=]q��34��}����9+��8T��D:X��n���=�pJ組s]��k{�ֵ>�1�4!M
SCB�"�Y�˵��lf^���2pUc3L�b�K���*�ۙ�ҝ��$�U^8лG�K�>�Gt�1/�riOFA��X"�G��/���OD�Q�H�o}�k52���2�%���;�'�[=��
�#���V�T({���LC��s�9�H�9�y�n~i�;6�E1L����>7��z	AinF��;��L��]���S�v�����`D�#�ȇ��ɓ����Xk(nϿ/���7�@��f3�y�j݇5#� �z��Y�:X<�3����>1nVZa�;�L�	����}3�UŇ�,��d�_=�����M��v����/�8�].�_��ӑ��~�H/�V����dV�����`�K��*� ����	��%0���B�ω�W��ge����� ��*?�8t���O���Y:M#n�a0�zij�q��Ճ��c �^�a�@w#}� �6�2=Ѵ�N�'F�e.޾O2.��_7nA��������o�#��O6^������~R�4#�Ʈa�q�����٧I�k'1[�N��N����\؉an�����O�[� ��Ⱥ�Lx�J��%�UޜEl:�:��.ͺ�k�]J�:9�un+�LwRye�[��*�9�m�{⡒�������{Y}�U$��V:*�U�bNM̢4�I`�c�����՜��X1�4WEdp�{�u8ͧ��i�`W��� }�IM44�{�+����O~fo����Xh~VW�
V����	�����O�F���ky~�d������˳ɶ7K��ǤS��
���B��.�(������p�Cv��QaS��h;j��z�PsX(�z�����]`1�]�ޒ��J-;c���]��ty����`N?A�ʝ{��=�!�:~��յ�^�Q|���O�S�y�"X`&��aJ��kk�e�R���
0[���K�{bX�ΡUjx�PX�9����y��;��j��Y����]�_:9��ú�d����!����:�S[f4��nɎ�v<�c�}a�R�)�F��G�� `�XH��^D;s�ᵲ�	��/%��/ݯBƌ�����>�9��=���喽;���� ���Ȑ�?�|d��.�R7U�x�U�$D�FV�����4���TZS�M#�c)�|Q����ֻ�>y�_���	q���!��2�e��1<�
�d��i>8"��׶y�
w���3�]�L)��,�}���骮Rf]`���.��7R��M�ג��!�&��D6��,����x��i��� ��GX^��<��7�K��<.u]�)��Қ��{8�3��ۨ�Ǯp�T���	z���W�3��=�C�^q��{�*�6�X�C�8g޶�&/�魼���qw]B+6=)=����.Ҁ^�l��<v3�˄b�7NXpv�Պ����3��۵�E3���x���yu�	���Rb���&WKe�^.dk���\[:~ON��
z��<�ݜ�i�c���6ǜ�6۠�̻�`w��˱���a�m��m����oc	Ɋ�L=���>b���\��g�-a_|L��u�Չ}_�\/����i>�A�_��z���X��5E�27�E� S�<��B�u1��%N��WD��E�:�lvpq�c�7�B"�<ľ<���u�'�s�s��B�ƎQ����iZS���@�ˋ�$�G8��;Hj�T��f�t�-�&�Ȯz�*�y�Yz�o:��������;ÐPY��͸"�s�n�	�r������{�;F�a��OX��X��_-��v��Wt?|���9�ɰ�Pfl���p�����-�pN��:c#�I�W0���,m\�;<�e*��Q��W�q|�z�
�v)�L=y�ې���6 `��mO	������H���
�2�Zc.t��8ŦfS��L��s�͔���!�@���0v�+�՗1>���8,J�:��������]1Z���Km��&���4�����hű�n���GW�ڳ]o OM�g�['��vY�4HMs��<�]�n�p��J~���i����MK��;=L
�W�7��(��'�-!=%�`��!i^(~_���������.����e<O'9G�q{�]	=������7~{ >1����y���,Օӑ���)(��`�0Kg��,X<���٭MO0������k�P'i*�1�=-��S�g���-8�����K2�9q��ӂ7����n��T�t��vk�N�9���e�A(�ZYZ�kݚ)�����8}�5�S˽�p�b}��{aQQm˶Y��ȶ|� $�<��g�0�h1��6wr]�)ۻ[H��3�1�W��$�����̵�+�P~��8Pz����,��!��_���H�I*�M�[� �._Z�`���Ĉ��O�q�}gB�<EWeimL����F{�c�uZ�	*��p�l�'�:k�}i����i�DҊ��P�+w��΋�`�.Z��v��h���;
�Y4#�Bޭᩀ�vjݩm�L��,�i��ðpR� �]�8Ij�~����t�j�]B�ѳ�� 8����Ƨ�k$tC5���(�v���9���%'c9ڔ=��|׺a���5��.��Ң6�b���d<w3 ��}tp���S+T�&�  M+A�×x�\$\���H�!�����D�g��!�\ۣ��]������u�i���G�9��\�Ψ�m+�z�LmL�b8&����A�wMK�\5]���F�R�Q�9Le�I8�@��o)G\�S�ͻ�(-�i� qۦ��gC�1�XZXu���P���.�3z���)p�x5���fswq:���e�ث�8�
��b��[���T66v7���M,�����/(�|�l�LRۚ3F��'bMVK�� �����]���ܿI0ԍ���h��pX�Z4:S�F���w��� yy7{Z�1����w*Wpa���Z�S5���Ta�](P#:_G���� �5ڨ��oq��k�+���=k�j�V)�T��s2P���%ƯF����b%�%�S,%�qX_�Lz�T���jYiM����:��D�{fQ�k��aج����6���]���Uݢ�����ggd��__y6��$�Mr�g�j�b��l_S�ȶ��s��8��]өQ�/b��&X"�7<�$�����j����G�����6�����k�LY	���=����B,����	�ݷ�CI���t�X�cVE�����3{52�p���[}�s���{#P����������mٲ�-B���ޕ8�[�ŷ�vf�&r�	�Z+7�$:���x����sɽ�{�3)髩���9]���y��V��u�Mi�p�D�|�]EpyJ0�Υt�<������Is���sof1١��0K�Eh�n�J�7&r�d�I��b�T�C���i�3�WE��l�̵x/���GW�ۍ�����d�!��]��������>�#l���`-X�x��P��}/Tw�+rgbiF�#u�'kK �t˩�e͕f.�!�뷹�rHp�tQ��Ѡ(��f����5S���q@=��!z*��gi}�r�s��B>pZ��L���xI�8ʗ��P2�N�)����B�����Za��8脛���'�/�cљ}g������5]��c4��l7U�(>���pH�۲$n���X���R��h�+��Aw.�db��b�v��L�Q���6��y	�S�:d���
�a�|��j�^	����-���0r{����*��`>s�8%�S���z��P6�>[b���]��ڕ�s��^��3(�(đ��'LҼ��]��7xl�:�off^�*��IV�
 ����G�y�؁D[�nV)$jT!$��Ǯ�=t���t�8��q�}}v��.�"�T�$� ��7�j4��L����޼x�ӷ�\q��q��8��ݿ7���������������	�n�d=}x��o�㏎8���q���v�p��Q�kǍ&���-��35%_�^5p�Ѣ؍_�������%�D����UF�|Z�XɵQPb����Q���F"ƨ��\�(5���]-z�*!��r��p"�+��I��E���r�h�|��^_w<��'#I�� !3̗L¤�%� "(� ad�RI%I��BÅ��r+�lq,���������v��ϒYEv�bw�Ւ�S�r��YN�j	�E}zqT�o����Xj Ǡb/!�lE<J�2�D�8�eHd��GW�BHcB��D�DH� �`��ڐH[e bI�Q4!PR���$e�N �i��q�j��w��AM%44�����w+V�O/�#���rӃ�FkP����P*��eI�;n�t���/����S�!Ŵxc�|�O ��9�8ᢺ} ��N��K.{����s���t���i�%dhr��L�q�=��=k��yG�ȈL1�C)dt�$�	�O�0�,y@�xN�Ͻ��6�q��<S���5;���?��˃�������?��9�.MQW��ێ�S����|�t&T8ʇ��ߧ�B�_�_+Bӳ"Kݒ�
ۃRԧ_xQֈf~�FEp���q�v�R��}��	s� �iw���tk��o	�8׏]���u�V����	�c��l���/��7	=��8S0/FŰ�L��šƮӚ҆%�2�"��_y���`���?k�O�O~]x���״�5�W-�gWّVP���6ԢLp���� 3?�0�O>�����G��k-����bu�(���;�>G��4�l^�k�5z8+�oP6{���	G㿬4_&|�к�����#�Ncߧu�4�wl7��!��}P��|6V��,�z9=��;X/��ӑk7ҋ�c�������<Y��Y(V��Z��������2�DD7�t@�9V�$����X����o��n�s��w\�1���.�	�ȂA�m�cT{v	������p%ҵ��ӥV��cdN�V�hѺ�#��:��Aw��G�L�wy�?������y�?���hoG��������r=W["lf�a>�(!eJ�D
͌OI��q��S�����/�K��Mw�63�{�3n�z=	����#W�7P�a�^�[A�ٳ���l�"�d�i�Mx8�>%���J�	?��Q�~���d�R�?*�g!�vd�;"y���u�^�nf�~�6[_qc}R��V��V���.�D���^Gd��lr��%�w���Ş���8+c�rg��Ǆ�kN��<魟����T��.��0�q�_��ŵ'���ʹ��YswT���DO9��f��w*涱$G��&[��@Ǡ'��!�n���H�wX��ok����;D@�+�Qiĝ���N�ˆפR�wU�,��}|�<l[W��O��M-�q��}
��n��]1b��@Dך0ZF��z	E��� ���n�6�f��.�t���=W�mzJL9������^�a��Vg��Z�����K��g�׊(ܪ_�sz�����"ϳ�AX`�S�}�fUZ怘�"7h��������%�}�A]���{X�� f��Qb�7f���U{��?��^�H3�`S����|9�T��9�x�+�:%0���1Zk]w�b��M�#L�TuDgGE]\�U�#������fR�4%n�B�u�}�� Iz�mi�������^!����8�Cv%�{�ˑ�n�Y����0h)ݚ_��k^�R+�Ė�b��O[�s_R����w/'m��O�>��]��4��^�������%�&�<3s���6Wn盨���
�k��ǿ6��K�)�-J�`�̛Y2����T����|��T�?���}O��wK:`cY!����K�}*M %~�``<��{g26D��7�u�[������I$	!H��?{~ �U~6�޻�z������P�1��{�����.ɵ��%Z0�k�=W~
�a�8�fp0t	�8E�k{d�)�QMГ���5.���V$Q�t��4���\�&۫�������s�Cg9�>c��	m���m�Mm�Pb�td��{��w�k���C�<k��\\<â�=à[z}a�8�C�y��ԙ��z^b\�v��I��O�;�?k;���7�7U�P���,)������+�U��[>`�����3"��U���������w���q�+=)��^[��x��\�uGJ�q��'r-��8�nf��~�����������.�"��	^�6A�+-.E*Sr")06s�OZtU���T�|��Id�.���"\�R�%�����d� ��$@v���:�m�1Pz���z��{�)����o�;���[���ʐ�G[+\���Yg�`�R^�򏿕�|k��׏�3q�݋B�,q÷��C/��ke��ʮe�����Es� �1e�T�S#Yϕz.m7#�r��4֑ͮ�t�۴Q���ʓ�a(����c�,�4G;.8�Z��S�]�5�*�,e�C�"�W�e9�}�`�M+,~ax�>��
~e9�$������se���R��=�Yy��b�4�/��	��.��Z��א���@�)ᣜ�H!U�m��QB7N*.NgD����a�`�R�]k	Om�Z]�A��wvh��ɹ�u\�9����l�̭s�3�4���צ����ŀ��k�@�[�X���Bڝb�ĸ`C��d��sΟs�E8����l&ލ�ӓ�~��)�vl��O0n`��@ߓ�ֽ�v��c�+`&���%�4�9����ފ�H(��и��{�`}��_)�D������bS�A(fX��"n�T�A,��WϚIM��3���P�$t�G=�n���^BE��ٯK��ܔr���B��<s��!ێ��x��5�� �L�va�=�Ͼ��zj>��{ Vf�����X��K� vc'��J�5x9�oH�+ɳ�����fh%!?_|�}���i���v�����@�F>=�R��ث�{է,'Q.b��o��F�sQ}�YL	hmZ@3I�����HL�H�ʁ&�!��6h��+��ם�����B��\��x���lf���TK:�Y�g3:��L�\��"/&�{5i�����龳	�u��Z�y����-~6:<jj�/1bq~wr�%����𰟚�_0oօ�"�7zE�^��t ��p��8�=7S,�lK<p��g�sBv��e��P�����oK�>rs�V��T��γ"S����t�*�U�el�ߏ���9r��w�G���ـb|����.{�,W�΀�^|BKQȞ~]	�2�]B� &��9�0�f*_��!&�p�/��{KX�~��hKГϏ����"vG���.p�d�p�k{!�W�Ѷ��ކ��('��Z���&?1s��F�OY��2vMIy��K+�+#9n���=޺v��,�WzV�30b���쎀��{��09�㔆PT�+��u�r����988�˔�Ϡ7�|��,yĴ-����͌����Ó3v��9̪�wf���!��a0,q)�u)z���=R	r; ����x{��N�P��ǜ�|�n%c�a��~�Gs���mʙݻ�$�u ���{����U#1�{4Z���bv'�c�.�TW�+��~�;���l8zZ�N���g+��k�ܹ�[wQ�b}��2�h�����_/�I �uy@'ܦ].��-�km$�v=z�۽!5�A"tո�G�;���q_J\��c�p�\zwdI̩��op���o0�ν��v�7㿐 ؈p?�:�04NZ�Ώ�=CK>���������.�ڑn'#�=mò�Iz��p�CB��8G'�}�>'��n}���n9>����2N+��ܸj4x���7"ey*�tE1cAݯ7�ya����O�_�Gً݃(�t�@�y��������<�B���傗�7Mmc�|F���3�ں\v+�	���5���jO6�O����<�G��\�+ڤ����o&�^m�Y�e��3=K��{'��:ڛ�������?��*=ӝ�B�k0iA�
���;�l=��9ϙ=�խ��zMr}X��Ih&~��삒c<��,�z+��%B��7��k���nnǎw
�,h	�)�Vv�u�;��}��nF7^���1��?���iܯ�c�-�`,|9��W3<^��bf{�'T�c�ou[U�*]�{g禷{�]Ls
��y�,b�팷��;ϯ���Sو���[�r�kk��$�\?Q�?�(��A�9�����+�o�e���q��,#nb\���W��:������u,�iI��O�����a��5S���r�w*c*�uv�}�2���L8MNT��v$��q{�;�<��B-��\�҃9��gXP����ܮ�(�h��c�4��M�{��g�ߟ2�TO� `���pL������.��EW���
b�bz��׶g�M���3j�ˎ	aDoy�=5��zHg�p �s���-���M���!4���6��a�j��y��zf��8I�O�<�Z���q0�ݯBLKm{qP�����h�-_�st���I�skE���~.���:�8��ե��>��������|�h3��I���qyݏ�Ҏg����e��^�^���pmv�z��O��?|���=	}l�R+��c�C!5Ԣ	�Ά�xM����>��	�K:p6��C�m��K���=1j�8ܝ��P�]X;-S�����r:NL�@8��0���-�����0~T�^p���G���3�]B��������"ge��05�P�􊌃8��u�: ���&���-)���a���Hz��r6.��xް�����4h��^��N�-Iտ��ȃ�)?s���c�O��1�ء���=�8�<�¥!�����A�|+���\��=_�,��y�������6-gԜ������MKj`-wh}}sgj�(#%�'|
��*4��
���	�8r]C�T�ʦm�Y�P��l�)�sR':S�ْ��^Y�j�����m�C�-�l��ՄnJ��o��+"�ֹ
[�n;��Y�v��<�a�8��^N��1�Ӆ�C|�!�]�k�Κ^�80#���摻0}S�i�=�A������}�t��#o��57vG�hʀH�3҃�&�D}5P��ή���_�\��8C%4i��Svk�3;p�ց���t˭H�ޞ��[��@�\<�{g�����sj�&��hz�op�-�!�9�%�������\���a���4L:vz/�)�?g5J��Ml��xC��5��b�TO�@ݮ�e���M�6-�?w,��r�6�Tۗ��u��q�`�Q~w�L��g��	���_���j����`��Ξi�ʞO~�ܟ������.�}'�C��\8n��������Ӡ�<;�pam�����^�P����*kt��:���ο*;�O-��s��*ʑ|�Cq,V���6>;ɗ�}�+1���5�[9�rxF�Z�YE�v�G걷ZD��0T�A����|t����3Z�o�Ă�����jE1%8���{]	=�wz��je�@a6�����RC�˿�j�Me��3�u��n�×�%�^>�5�� g�U���]]�:�\�3A<��Z�D��p�W1oS;*��]��Sl�J<�Iխ�Η��.U��A�qy-��^=�v�]J�2��l�5�C�����u��ט�{��7�y��<�����_e��6f5��>=���SsZȸ�s36j3�r�ٮ~�?�<(�"OV
~���s\Wu�ā���w��A4����kn�E�):�7�H���@f��-?0��m����������S�P̱Ϣ�X��N�,�:ͤ�;�T���V���O�ƥm�"�)Em���`�q[��w�^��s���Q��ˤ�wq�iX"�Y��8f���x=������ަ�U�p/�m��(��]ٸ��8��6��B��^g�dn=���5B���G�~�j�&$h������;�ժ���[��筥clʅ����n}�8�E�T:�lS;��텚8;[���a��-0��Ƕ �G�n�<מ�b69�7dO9{�����n�whP��D�4lK�v����k;vҜK\������DtcH�Ij����)�6U�/#���]��nZXz��y3���JV�!`��ߣ���[�"�g��{];{�:!��u�[(h���׏�b���\�����s���#�d�	���C+� $wC��=�ݥ�/���]����Q��kWk#䦽��v�;��A�"��nM�E��ȓg@��� "�9�wY�=��Z��4.ǘ#�y����ݴzB1�O�:v�8:ad����fuoH��Fv;�K'6��*]���I�;vEN�� ����ǜ�?�4��6�t���z)?[�*����n�v�+
���MA�6�;�G��r#�g4s����:ا\��-b|ҸL�q"ʯQ��
��ֵЙqoBw,y�%��}�v㴲�e�0�U�X��޳o	M���$�M���Ms_���)k����ktWu^� �'�����].��̔պ��\�E��mf�^�����LK��cgi0'��}�Г�?Tz|�
�T<���FA�@���@�C���o���$N����v�r�lt�%�S�5���}�c�Q���3�����Ok��BD����^�n|�צ�f��<2��R|�,S��q�]x�nH@Y@#^�{D��U���������}�@��1V~�����x.�6�|~����@YV��wc�zH@S��}�� �gV��%��}ɂ�R�T�Ǝ铭J�5cf�����,S�=v��k��C6K	�B�R]���|Z�%���'��m<��ww�U`�C���/���~���)鳸��a��t���5�q��<#�j���GZ�^�<6��_�Q�#-f`ߣ�O��8�r���
lJə���ݠ�Lr���m�L��{mwW���&���g3��ϴ��x��:ӯ�%�7���I���,u���ԕFRV^�.+��[�tM��MM%�dw�{���&s
�J5r��
�Ge+Q�\o���;K�^��oQ��q�<�-�ƅ{X��X;�c7ОRӆ�V�).M�s:�W|]��{25nyܔ��*�c0�hɑޛx�Ļ�[�,�i V����z�X��E����"�����\�b��Ю��.{�=Nos'+�Z̫�}s��E�3/���"�8��M�탌n��/.g,�x���^L��5R����j�71H���Øk�_tۘ�a�L�4�=�ɦ�m�w�G$�y�ɛ�9Ҝ�R��[੬��I��޻z�&�ҷ�4�P���1�B�뜭���qLI΅�cpY;�)��3��ֲ�W�>���f�V���n{=��q7P,���v!���X�0}��7�:�X�#��Iy�>C��,Zq�,٧�n�T�b\�"��elۖ����
Ƈ#��
6�,v�z�az8 Vu2����j��Y�����j��(nE��&���gv=:���y.h�:���{V�5��sX�|E��:Xql3qb7;}R��c�QF�:�݄�_��
ѫo�&,!�����5V�N�)�p8��+�,��$�LB55�X�`�UP�^��B��8)���R�0�
h�T(�Nv��	��?u� ���-��5S=��jr�_����[���K16��\]�e6�	�v��Vtޖ��w�E�(eZ�)�u>�shm��wǡ�q�2Wwl�z�Cl�w[��k7id	˫ZpnK�d�h�h�\��*���y�Y��^�yF���bE's+rÐ.R]�ݳ�BC�n����e����jk8�q�סc�^�����.&�����U��(�ᯧRa�{}��[�z�����j�J��K<�j��ox�)�]�sW8�,��(��NT���2�Ǻ-�Jgc	g*���f�&ѩC��Y�F�K��O�h�=���5���84�-�\4Z�t0OÎu�g77F_$Ҳ�8�;%4�TS7Mj��$���a�֍h��n�̓��ᛳz����q�䓋����=�q�[4Ս�ٶ,��%��4���F���_S�8��I�@�f�N;�n���}�V��u��@�����%I��6Ze�s�^���8����f��}�s�_\ts!�\��M��ˢ�v�Z�{��N�*欋�huv����9�WP[�饆e���1�|+C���JvQ��E.�#`�K�Ӿ��
kz�n�D:z�ݙf�=K����wN�:�6�t��
0�]7��Y�y���D<�@z���$I$d �����o_\q��z���}q۷o4�B	'�*-N�7A�&���T"K��	����^6���q�n8���4��۷mY$"H,�j-C2�55<��@�UD�G]�z�oq�v�^���O�]�v�qd.5A��� o���ε�W�x6CW�vƵ�W�i�_����đm����E�(ش�Uݯg��J�FMoٹ�Q��ҽ/���1�����zڌb������K^�gw$��ܶ#h׮�y�b6�W4F��nr9ok��Q�I�>1yDδ�έ��Xܼ�4ct��5"U���4K#����^f�G�n�5�������*v-������W�^^C��x�G>:���&�Y@?৶~��BËk����������'�ю̈́��G�x��ΧGz���`Kݾz���ٟ�@��
��& $�; l�c*�,j}�V+y۬��퀱�?w)���]�.�>1jg��{w��s:qY1�
�o��L�E��[B�y��y��I˼'��L��W5��9ޡAld?'�qM���T³T�i�ٟ�����HE$W�怰r
|GO�	q ]]Ν�;�y�ߚ��i�b�OO��m|~�ɚ!r)�k(�a�AG���m� �n=��-"ܷ'����=��An��6j��rb8�#��.���+[ �`d1�a�ÐE�X�����P�'��R�nn�X��I��朄�x���j��������U�
!��^;D$^c}خdI~�0%�������Y�t�l�w\XN4����3sÎ]����u��W�*�>1�"����w��>hx�=/���c�vT9��G$f�%h[<�1<�kÞ5������F��yoA��Y�(h@�p���n}� ڇ&Q��;UݏhĠ�zՍ�M�ôugd��Jz��W�H��8*%�[2��ݺ{��{J�~�Z+I,��d�l�fSd��Ѫ��Tt���鰉7'�\��s������u�Z=��:��H��Hބ�}�xxW��y�����wܓm�z]���hoo7����bN��s4Mmy*->NY4�^��1�}��*U[�p���'a���{����闷���������LJzC�i�P� E�E��V.rw�oUbZ��,/�V|?Ab���z��?��6h��z2=wFDX���G�pj�s{_�L��ˢ�I2������Z)��m��'��{�nOsq隊h������r��Iqś;=���^�[�l���H��{6�W1e|��I1c���� j�Q�l~�c��u^F����&��0m�u�N�ӀqЗ��ʼ��g�}�+ֽ��}����à\��J�@���pWvk��,�̆���'-�=�#�}�W���j>�d}��\���ַ'���zj���rl��27�Ej8:�۾���&�0i�Q>�S�Sc�s K�x��P�ҹ��d��̱\.O[h؛��lt6�k�U7�H�E��?s��A�j��0#vz��g	�����⵳|YC��BIӅ�z�����"��?, �_����p�C��	o��r>�q��pt�x[��/��tr�)T���82�_8֢J��G�������ޑ��I�XϦ������׸T�n�Tֆwh���@�_X��tXL�	-��yh$���ȇ+�ɻ���n%���������6�S��c�W�)�Ӑ����<|G���+���(��vx#���C$T	:�I(R�hW�Eo�;��!�����t�o����_������_��Uǥ��u+�z��2+px��o\��{����&�����*ʝ��D�|{����l��ͥ�Finl/�y�ǧ�,짞�#�Gg@�K�֘_i����a��U{��lР~�Ď����_~���um�p$ü�"��`��)Q� ���/k� #+�0�8��POlb��؎umW���֔
9���l	��y^�eRXsO�;�Nf��}i�	P-S�[��\�c�JD��-!���!�����/���Z�_����'6��~#=��w��ƒ�Z�tյl�z=g���y�
����)��N2�s�E�����-��acs��?P���v�IJ7zY���OE@A�e�V��yxcy��(#�Zq>���+����m[�:/F����Ӿ���%��p��n9m�r���B������GmMU�N��Mϫ��[Yp׼l#8E��{�Ԋh��-�\�T�AIJ�GX���p�88�I	����3�ʋ������fC�yuG��N��?_0�}�oon�>��n�o<k��@M*ٷ�R���88�O��u8u	ܘ�����8����!,^�]F���|,���k��z�����q��߫�¼<+ӛ#ႊ-�Ä
l��^iO\���O����<D��H����l��W%@��@�,6[�
B�:K�M4����I�a���C�?~>'E|��	-��zw`S7.��ޫ��:��jD��i_���n�}�O����X��8����3я��k��ʡ�8Τ#��]��;���Wo��ܟ��q�s
s&]�s�y�	�3��S*��Đ��Cr��[����Q�䘩���9?y/�ڨ��6��;�/H����ۍ������g��U���{�6�遍�/dI���M�&��r˜��2��W8����e]	��֝����25�;4{�|���#�D<=�<����B��u)z�x��wo�z�[3%��nm�v�X�K��XV���_����z��/}J~�v�
'����Г�>�lY8Z)L�sN��A�OS��-���`�0ff2'������'���W������k���+^�D�Wf^yZ'�޻�G�^�r	f��ܨz`��x��_�i����n|�m���MUqh�$f�U� 1�c�����B��eo����+�2��]�{�ܛ˕�kή��z��I�~�Bu=Ŷɤ3�'hn-&u��=;7�5�nm�8�n,�y� |w�S.Qm^�
�������
"�n�br���<�a��{ը�3?��bw'���o�g˸�3����W��a����f���4<�Q&��Ee�GqsՏ���ײ�A���kݎOIx@R>�08e3��J#�P5=�x3@�>��wW�6�8;p��� �	z��~��[ё�)��W�Iwo4�E�Co!��f�0�C�.�:zaᵡ��r�'����|�N����ǟT�)�gwP�y7wE0�ټ-3����[�;�Γ昆k~>g���ߑ�e}�����a}�O;~���*����4׹��q�Q����w�K=ƥ��6�/�ܧXR1��oV�ny�8t�,.}~���7<�;>��S���]��:	�{z%����M7G)϶��{x�{w�HP9�P�z;�4U�mE��u[;��,yu�=�)����[u�]O>�d���\?�I�նܶ����Љ��&^b"^%��!��y�K��7��Ɨ�biWs�Q�u�����E��<&
q=�լ����EP��rK���F0�Tz�st���K<��'�X�ܝ'�r����Z��;sL�3��D� ����}�6���D��u���.��un���d���|맪����;�P�B�f(܂8�Q��^�\ W����a�=&�F�ä��Е-[�N��.`5�	է0च�y�=<	�ʎ=�5�=H��ǖv�߫��{��<�����zƗ�+�ɦ��.�(�<_���� �3���
�vO��a����Աߌ�H�7�Sl?{�=��7�?&���G��_j��ʑ2'_�`Kn+ܘ*��ʓ���-\7�s��O=_\�<��f�;�6;p}a�0���z�[��U�)��KGmȮ��M�����
3�
����^�k�
;=����?#v�	�f�4��僓v>/x�=�.��E�������[�6��S@Z����ɨ'��Ǉ��Svج�A��x����(<A�P�2�.[�u��Y�q�1v�*8�(]P���,�\5���gt��l���?ɏ������o�ҳ�:�{��+c6Jr�)��Ej�R�xۘG8�x˴�ƴ�ͼ*��0(?��`P��~�t�|�P]����s�9+,������z�c�sWvO�ܤ5�Mܠ[W�`���8�,?s�]���ʡ�S�V>(޶���I��W��I�O6���5�*H�3��7�k�Ɋ��6�z�cx�a7q��X��;���D�w1�.8*ZK:�vV'�.uz��;59�vH�*zw����ܳ��19�j5����5�+a��\��wts{y��:�����0p֎q�7׍t�/���Ϻ����� �؍8Y�����f�g.�����N9�^#��xxUf�z�(άO�o��TAG9N����J�S��c}Vz�]�ij�t�0N�vo�"�@��D��������|mi�����W_�X��뮲eŶ��P��bXWv��]N�Q.
�t7�����{`E��lf��%��O?X\�uGJ��Y�b[C�d��[@��	t[A��oG�=�O��q~wA�j5�i���=\��M�Q������yI�����M
�Q� !����	2y��gnm�מq��d�~���DV�3��<$\��j��)�?g����Ot#4^��kýC�gkg����%������_���Y���g����֢ycj��*�T�'��34K��~��w=6��՘���c�s�l,X�I�p-x�%��OH2IN-.��p�I�~�]i�� g*I��A�ܱuN`_}]���R�c�oc��1�c�Ln�{�<� v��'��r�B۝n�d���|���f) �v���ڜ0�X�38C���>'�vn�%�y=��.��v��"vu�a�Q̀��q��'�2�������=���x���Wb0	\�n��^���Z`���ې*�6^O[L��> �uk�~��y��$������F���w{�ʝ.��38N����������y���^���5p�,��/��oVJƄ�.2��G �֪Tν��4Utq8���Kxw~5xy�U���5�o�`�$�{��m[IiV_�C6�����V`\<(�חx�g�>�w��=��[�wIz��P �M��9I��S�?R=�B� S�{��" ,m#^)�8f�
�{N�E�k�'/9Ut�]ٟǩ?Kս5{h��熡�����!�ϛn2�[٨�y�Y�4�;�e��5��~M%h�8�S��5�r�:EH���mz�2�R
	J�Y��:�;+�^`��� ���8(��F��{
;���{n����'�����P�rK��<ЌJ�#sAv'M��3���E=��p1m)ĵ�zX:|�;�].��R��z",t\SM��m�Cq�o�zy����M����������S��� Z�0�~�^��Z�{?_׀���|�մg��ͩ�k��x�\��)�r�`C������s��va@����7t��槳�іIa�Xk�L�{��	�O�/����x�Su{�P4�㦠�����zl	�ջeGH<��S�Ұ�m@s��L�mH�q���T(z����m�t&U�z�{�K;��+�WQ7ϷP#�������m�8{#���شv���O;�t0�[1_��E;S"U�a���z�;+���ֲ�y�C��:8v]���]���=�V��rDcZkW[ںz�p�y2]v�Opk#jZ��'WJ��K�/��<|}�'i�9ߺ�pi��
�x�s+8`�=�J~�0����.�{�T�_/L����kا���/����������^��AP�������j�ϲK���mIad������ͺK[l�quQ�ni����2����+H��������h��;3���Ę�Rh�n]}Q-�t�K1�./�lwO�^�PYm@�������C�#���؝v'�mRh�
��ƫ��tb�%����'�\�i��&;ƍy�c���ϵ��<k�4r&������a�G+�/����V��y����^�g�!�ʶ��$�-'!P�,ϖ
^�������s�ϡ����4��u���<=���W�Ϯ�JS5�T�P�%�3�}̙�+y��G:s:�V&`�b�>0����·x�X�|D���<��,���I�.�.!����t��;��TAN{�#��y�k�[�l�@^�P�08Ɓ���D\zdŰJ�s���\r��)`7�8�k�<��㟸�0:�n���зf~�b%��1���f|ݓ��~S�0�t��XޮB��ս���T��2�G���fՋ�v�vX$�$SQ��aLc�C�I�sC�}�)j����X����Z����+�!�ν��V��v�"�n5n��cVa���.�b��w�Op�w��{<���o7���ۤ4�p͹�@�ͨ�I�#4Ǧ���*=pm�q�P�*�,��c�;ȩ���}݉c��a����; �
1�rT��������]u>�|/2_��n)����0 Y�7v�+�Ursr���^L����ޑd�2��1~(l*H�\�RF�տ�9����\����
a�vȂi�Om�R�=��}Д��ʓ:C��֜r�3ғhe��k��u�B�G:_��z��)��>�;s	���$k@�׽�>}��C��N����z�wf�xLq���={�qWhWZy����|��1���s�ɛ,�:��� ܨ��3������|
&�W����m�`��Ѵ)�������.�L��~�1��`,���-���2�	]	�j��NK�m�"��;w�[8'�������.��aH�� 6�f��W�3��g��Z5Z#P���x���c�aT���"e�o����܌�����K������5���](��7y,ܫƺ�}�6+͜����w������	�0����;�J��[GwC�j���en�wa�wR8eZ�xAZ*�j>�����ø/Y�93�e����w�je�Z�Ǜr�f�  ��9����0h��x�={iګz�� ������x�a֯�h9����ONjmp���wr�*�MFZlZ�2�o;'m�)�x�;��9η��M,(l�����"/��(SY�aYܫ|dC��Me��g7��]Y]�jEi�ru.�݃ǨPU�"�svJ�Q�Mـ^e	ʒ�&]��h����`�ٱ�[�h�f',c�r.���'K��9�H����罃/�W���+���PG����f:�9eu���%�u�ER�ɲLh�.<CP`���m�&l�V��'�۾��<��nW]IzX�j�E����û�3��kw��j��>6��Ӵ��m�^������S\�EE?��z�f���g,��Ud�B����Y�(Ԩ�s6�:{�+[~�g�##ܯ�8+�\Q��a�����E|�:��V�#\��̛dZ�Om<wr	[����2z��iG+{4��[�:�o^Ҏ���-^�\���s�a 6�Kj,v�Q{�g��Nc�稏lvx�4��3A�'W��&�3��9:�R��`���Z"���7\2WI*�m$�5(j��)���rdwpK兼c����U��Yx�r�a�6�0�lob�i%==��s_G�A��!-S��u���i �K�']Z)�G3D̜�a���涚��vU�.�O,koR���sj�ʲQR��\��&G}N�a�|�����s8Y�W���ʳon�m���i�[�jj���f'�
.��Q�e�YÞE�-�x�N҈��9W��WuXO����a�ճ��y��z���;����Kf��r�eEj�I���V:>�f��<}hN�5�^�Hz�wq1s-��rF�M4&�0�Ěnh�����Qy�E����r)�:u����*�������u	�r�@�5gH�V;z��׃��	�0��3#�D͙��`4�7*������9���}�ʣ&�{�l�W���<e�f����-��r���,�*��h�ȝhZ��&�<+���iXB�V{���)meؔp�ʒ���}Λ��'B��D��l���mY��vr��Hsy(:J]����k�o�jY�k�MNPu�_L�M�ͪ4b�2Rt����3j^d�4";)[����]F�|�&�#v�N��)��>��g�.2|��9]���|6m[z��۵xdF�<ˢ�{&_@A>$lco�����ms�o
I �4�>=x��<z�8�z���>�||j�2�j���Pz�o6�=v��;�\�Ź�@��n�_Zx��q�n8������[���ӷ~Ε⹤�%A��(4���ch��_[��߻��֞=q�qǎ=z��}v����"�U�Z�-����8T���x��F���f�Th�����؍��rK�nj#Wᖽ����V�u6��*+үJy�c]5�΍clh���X�k�-�[����~�x���絮_��xռk��U�x��E�	 �k"��zL�Dc@�H>A��8"i���@��,2\0�Jb45�����\E�qY�e�>3�R2�p�49��m֮b�ꐘqk�Pܼ�v/\�9
Ef��lap���F�M7yrF�A�a �i��Q�[E��D�b0Ƃ$BS��q+�h��@��D�����)��q'�����%#f4�m��D	� L�S�HT#r�d�������y�����h�KT�;�Q;V-��,����=����P�gr��"U���|�~_���:�(����ʬ�����?e*�j��-�%��:{��ù�0e;����t5�8Rk�X"��-M��Sy�
�$���j���8wup��D
�ot��~�-aM�j�7���l����[=ѝӹq�*��;EJH�j/l*%��mh�M����^5��z����<<���G/}{��P�J�J�/
��v>c;×E����t�"4惲�q�����Gs�(��?����7��%��$�.��<W=<��.ǉ�����7�q�� �`��5���|C̎����i��N�����Sz���eqR�;!��Χُ�>0��# r���xa9t�.*ˮ��vh��J�Z�Q+<_��>��>a�M``��!����feg<�R��ئ-��mW�P�}�8�8������x�U?/�mK���:�/�@/.��	95K����/?zQ�٣�E��qST�5�<7��߱�U;ϛ�-eZ�>6��l{��> wb��ܟ^(t��������ĺ�:_L'X�]<������x��P�3=�7�yڙ���osr}1�1��{�{��=�����#M�oj�\{�uOunϖ{6A�������7*7�4���aÅg���dCV���x�OiD��ܑ҇���2��L>����E�k���॓��J���F|����~g\Ջ��9���<b�I���I�e�sb���~�A���P�Y����I;gT͗�Ԝ��r��U�'��'U:�l4�T4b>P�{+n��;��� �~F��:�s�.�o"5����Ʀ�zU�?~�%���H|�ck�{q�Y��z�*�&;�v����{�#��yh��2�4wb�:w��u���q�wG�2VC�O�9M!�
>�J|��v�ު0�J?�Hac�2��ঀ~�jS��5�5������@���5���6�]���m2;k�!fN�܁SO�map;&�+�Z]���ro�Y�r��ׇ�]��������U��j�0*T��Û��.8�A���V����wSTj,#L;�,��<�(�����pÒ�v�4�EA���$��D� zԣ�%�i3=�Z���}M�\�Ս������<�a��z�g��ELn�>���F��]M^�w m7@�����r���7F�0�n���|,z��6k�$q�o�"���/׭�
�j��m�֍Qi��՛��W�R[�{�r�]e��;fY ���6��eUecu�#�4�9���GO��
אMv��J}ǜ�Ԑ_�Dh�:�ã��`|�=1��w�$���U�<�bqAk�97�-��(��Tgl(�<n2��Î�>��w�|�e�Iԭ�wa$q-H�&j�͙AS��܌j����ǡ��D0m���"�·����18A�1o����=�/&٣"<��]���~0���]�%�]5�.��~�kپl�=�_�32�H?���:�I�k��c����W��b��,I���x<+�}���ۢ�7R��Z�m�UB��D7z33��� h��&�$�����S�2��n g �ӵb��8�������Y���\C��/z��j<`�2v�x�44TF<�,r�^���)��?�3�����:�^��I���ś�-\ãx�cv�=sis���k���^���X����b2|a��z�����5rkּ���n�h�x{�����N�;�;,����S���8s���EA�>]���鿸�����{��Z5	#%�ơ+yq�k���tl�c�?��Z<�s=iK���y
;�Tf�̤�xHer����}h��s$\ө�3p�s�mB�먺��x�w�;@y@xe��U�xf�K�.�1,����H�e�w�1���[��js��B��k'�_��v��Qx]^K���˥:���m5}1qV]A)����D�j` '���z��ӓ��3�<=��x��l��;�T؍���֧�"Rӽ���n����,(�e�(q{�B�W��Lm��H���m��l޳QX�Ӆ�X-�WP�#�gp�n'�+`A�N��ict��v¼}:lRԶ&�wE{;��w��Pѕ�|��n�SV���/�n�/o���e�o��w����dc����i���v]tCn-&���s��ϳ~񪢉�}&�"�,�PIFK_"$%�.��r�D���;a���[r��y��˾c��vv�]�5ԷSr�x�W��xxy��h;5��kؕl�g�Z���m�ȍvC�����kCff^�V��h��p�_��r��x��׺��r���g~`�^*mG�n��h���x�y�R��. ��a�}�u���1����i���9����ct����@~���̥{}����*�M��RK(=�lE�Fç���F�q d7F�8A3�o���������t.�z��2��;��#�����p<���z�N����4Yg\�T�{��Yő����_H3۩�cI%!����}@Ż-�
P�@ܶQ6��װH�g����/�n �W
��~i��=�0�����P]J�bc��i��;�Zzk-4Vҵ'���o2i�E����al�������+�O�L�w*��9��)+t��Ju�=��b��*�mrcu	M<�V��Т}s�B��@���7����>+��r����]��i\HwvS2�E*Nvr�mQ5�s]�9{��U����L#��l�S��'3):��<O�1�m\`R��Y��[�1w��],���Ŋfo[�R�I:9b���1����S}���3F��P�q�1�7�w�9Z�=�gw��4���q�n��G�[��C�դE�O�l�xz�.��4��V ��u�3�!�vx�7���~����b�o�2L�����x��i+�8�+[���%�e�?��1�]�`����B�sw�ѧ0V���o�v���&���F&�wP�JK���;�����n{MMn�ZG�W��5��!7���=C���U����q�[/�6�و-fK�=0Ü�`�MǓt�`��iD�c�^E��9�:۵�O@���L�����U�7���{��9z�J�׽Ʃu�
�ݑOv��[-(�&jI{A9���40�
7��:a�,��9*�h��vWU�u8!��*ޠ���JS����E��S�����c�Pk��ޙ��p*�Ⲽ�ܰ�>Hɶ��ʇwg�P] 4�Q���+p%���;3����z��Z�f��S�l�6Z$�/��:���E�����.r-&�]C��T�oG�\H�%��y�'{RyZ��:8{��5�E=+s|�>�B�����;,�0�b�4%��c���O+9��������|C��x:�e��>Kz����n���W7B��ּ�h�w|��n!8ȭ��t׳Tèa�]��l;y��=����P�r��̽�-�l�ҥ-f���v���.ֻ��;�[�X���@�qA(r}�l,����f3���Q�w�N�Z�z8�m��e�~�Vρ\{�b���H(r�w�A9W���V��]٣P�H�	�\S�܍��N��r̛�ww[��Q��TI�[�@��=�O+�x]C�T�"�
l�]<s��
]�'9�R�F���=�E1$ǲ5)�m~	�����5o5I�̙����ųm��Q�B������í��B�UEk�3��!s��k�P�z�k7!�������;���oq���O@a�Fǝ�0N���T)&�����}[-�q�Zw�-���u�6B�*Z�</\v�W����P��A~�?���*�L����ӷ�艄_i�.۫yG��:��O��7y�e�Ѻ��t���{7����XY�v����Y���u���L��g�z��s����~2�I�R��Nb�/p6���,/�;o�͎�X:�� -^IV�7#�7����~��ֵS׏����hu/B�͞8|Áq��'���Х�K�s�t�GD=��L\n/c��x	���"�ה�vu3�,۳�ꩢf*��h��ٜ��e#f+��-�ݥ�il��t��I�l3��`���;��74K7�VKmح'C3y�B����<+�d{����v������Q~N
=�I�g�t2̇z�bQ"{�)�L3��g�Y��{����d��^~�ը���vQA�.��u���w��-.���������ȑ���*�3T�����ꙶf�7IA6Yf)�)�"f�ɰ��k���4�m����j��=ܜ��º7��i��O��k��d*���I�xds.%zE��TU��h�X��3[���v�
^���X�����\�j���?cF���H�]�9�:��A8��7P���u��s�u^��}^���!\w��	w����b�[����==ڝ=��K�E
�Q��tl�p͊�d�v�G��)w_�<?*����Tz��ږ�^.%� ��bZ��{��;+Q2d�
pS��H�t�>㼞E"v�{�p���r�t}�n��>����}���e����m����P���iJ�ߏVa�ʬ�۫8Wx_�M�w�|�����#�UG���'���ABoZ��*�ruӣ�h�)l�ڻ�����q������NoD<C]=]��Ow{*c���Î���>;*@'|�ep����3ҙ��<)���u�������7[���tWq;��vq����Ëp�=&\�|��~�]ً�r����I3��ٶ�Ob�ɍ�3�l��Y��b��6�"3��3�wu�qJ�]�Kgb)� ��
��Nb��,PLӃ���������!l?bU�+��ݴ\�0ck*�i�2�cZ<�e��D�V`�n�d6�0'�?Q�A+����n��繡����V7��s�  ��X���������Y@|-3���	$����u&��}gq�u� 9��o�zV��Z�]܆j؏C��]^��r:���4R�W�б��\��Ш����z�iG��4^F�Ζ6�*���ݨpVs��	�o��Ln�F����ҥ5T��g�LǕ��/���l�О��i�au�����^�AvP�S���2���"��۵�;S�1]�v�]�F�h;��0U�ysa�����o7�ҭ٭��������S���[�%��;�����{{�0m�r�5H-Ͳ�.�l��ӧE FkUG\^t�oaW���
���Idi�r�&������hSE�Bv.�����+�Y��}]]3x�B����֥Kl�`M��d��Н������2F�UāV���K�R}�"�y�=����w���1��x(���Ж�h����ߣ2�oّ�wbE�r��!�ZE���h>�z��V�$�~+���u.�>m�HT�Cr�B��4��rT�m�Q�အ�'��Z�ۓ�H�L_��ڟg�d�p�o4�t٘���VjX9���#��"��ZA�گF&�wWq2��H����,��n�rv=.W�|�&C�i�"96E���^'�W�f�M��ݸ�j�IFt3�t�P�1#����y��zX.U6mO)�n��Y�ϳM��9$�:��Qk1J7��үu<�D-�DNa��c��Z�`�B�����ۈ9a���{9v�a�mW �=Z>voP����v���tZ�.eH�1�\B�I7jcY�ST78ރ��ԫ�%��|��+H���}�i��z_PJ��lv`��$���pL� ���X�nfFI�E���L���@�܄UY3^,ш6�nPU�������m!##	t>ܫeeݬ�����+�N�&H���2��l�u�}u.En0�Sq����|�P��G�b�	k��W��l"�#9]���e����pX<�(�W(6�N�#�z�a���ݮn9s�M��u`��+�[+\��o��_'�N�]��b�L��pE�K�+l�t����5g�i
ާ����ut�Yh�04U�`��u�EE����4"onW5Z�e��K��Hc�y}�NC�5]���1t����� ��n0(���$��l�/i�ھ��(swm�K�W�y#���]b�B��e���t��r��|���p�d�k��_u�'�֥�%y����T��7��bΠ@��5�}nz���:w9>x�BOf�ĹU��
��)}t%�ל*��=Gy�"�%R��ͽܒ��N��� I&�/��/쫦��0���Q�wvRs�����Gj��bq�t��MlN��v��Z{P����`���<��8��߁ǲ�˔�Y�Xn��pC&�TsT[�Զ��r����Be��VW�F#� �Z�
�@�b�آ��ԝ�]��\��}�hil���o�q^c�E1/�`���p�Ʋ^Ʌ��.�_D^l:�݌=G_� ��^�6���C�dw/�2ٺ�����3�4�F�.ю� ���R·q�s���57��Z�	�Ѯi�E�M[wg��-̬�%����o���1�-���I�b����ꖑŹi$t�E�z�v�	ƤsV�fn�+��F��ŧ�r{��Я�[�k1�:Ӂ��--��N�/�5���cy���<���7�PZ��/���h\;	�`�
ţ�ەup�(�V�I�G�
����f�̝x;�����泻��b��=3��ݧ&M�.I�P}htU��W�#M�z��CS��Y^W�ດ+���t2l�8��9�UC"�F�m�"&;�5C�4�#Lu�{	Y�m겲�%��:����oWepڮ�{:>P��o;��՝Gy��B�X�dyn��}��oe�Բp�pj��Ƥ���"�EI�s�b	��;!\¼�/yb�6��5$2'8{�^�����p. q{�!ؗ�77 �\v����=z�8�z�������.6A
�� .)pdT��b�q��۷o�x��q�8��������IQ�$a*ơ�&�___���8�8�ǯ^�����p	*#.�+��&�E	�Z���!�b��m�\�Z�^5~�wj�oJ�kr�x��ݕr�kx�\���W�TU�-���ح�^u�V�[�+r�r���M�ƶ���J�-�h�ۅ�h��QPW�W��x�I���r�TF�h�}ڊ�h����z]��J��l��Wr��B>�#Ɛ_��c��~b0�u�uh�%�2u��G����c��N��D>��6���ޜ��&FW�L�Ǧ������1�c~�=��5�}�y������_K�uI�o�p��q�:��D�W��1f ���]OP̍('��&�gy#�ڕC��[�Ds>��y�09����6厫U��_���xi.&9��I�	3��H���{��v����cqm5��l@<euz*�W�c��y�	�wk��ܟ@�E1�7�U��1����C{�����>�1A7�E%1^��Ҽ�����6�4�:�\�����9����Y��$�R1O�3��t=ܪ�9����t/{�s���Z�!����JSCB��}y|Ā������z�ty�)O��d���f�6ڍ�á��@�^�ݵا�G,���K��*��(��e?�a%ҟ1�6��gl��87�c;5��tuCo8c�)��@G.������M¾u�un���X�6d��~�S����v`ċ��F�����*BEs8�O���嗤����;fE�Ft]h��W��8���)����- �k�P6�Ff�h�װJ����<)Y�~��77��:� N���i���m��rǸT��v����y��2k-��!�vV��f���S�N`���>�o�^hw����y�ި�Z_^�$e��˲ ��= xRP7d�r�]����;�m��r�"E���R@������!�vO�{myC� �[	�΋N�E8���ھy�3rp1�m;�d����Z�mF�d�#Y�P^;�'9U74l�n�������a�tPa�^0XT��uLu��T�Xv���$s�� ȉ�{]�u��{�{��Jd�g���H�� �0`a�+1�2���\N��6Q���{�=Kg^�N���}l-xϻ�>%�_}6������&25ps��0�+���[E����$��tQ��4��m�A��y÷���}�����ݶ��cQ$�)���]����PډDw�|��~p�:aﻪ*�W�����"���=��^��u;T"p�p�x%-�{�X90���lކ|����^^���Q?�~%��P*Y����K��&z6�N�;Ifnԓ[W�R����y�'1tZ�9֞r���-=���������Ӷ��/m�`�oD�ǯ��j�+���{�O��]�=�6�BN������~������e{7y���s�X���Л���������tr��v��;���0l�׏�������orƜ����
�X������ݘ���3��\%ou�f$:�p�<�Π����m�۳D�Z)��q��zpT����r�6?�z���F�0��7)�3!m�gVH�U��U0p��^���#�u:Q�{�e��,��K���3/���\�S��UK&ˆ`��2�]^�m�NGNoe�Lt�v8�b�e�ӘeQOJ֬٬�6L��K�ُm�xtc�[ A�LC�ֆnN��Ɣ1r�����=��Q�q�6��0�@��4��i��wzt�M�8��s ��F�ؑG������	ټ�mq���	�6�Agul�P�N3���*ARx��K�-�[�w{������]Ud�3@ؗ���$���Y�#���m����"3��Jz|c@5���Z&�B]�WT�k�v���2���5;K�X���x�0򳇆㬫+�{�C��N@;�{�$w��Y�
c;�^]
�ƃ[��X��VFS��WSn���^xۊ�Q6r��:~ý�[�����X%㜷�&�q������(�cvM��33p��y��aV�nN�% ߌ�A�7��y�s��������2�u���O�kT���8��ޅ���;eP�$|�_��X���f��zC1I�t[�	0䗀�{ܪT���|�+�%Y�P6�(���<w�5z�9ӭ�j�*�F�
��+���(�G���E��῟���%*��/�cю�C_�C��g5/m��ɟU �Ӭ=�B]Wޑ��$f�Nu�0q��/ m�
7��y�����晋zG@�p7��-4T�	n1�#�gq�6���c����gf̯�����[�2�z�e���UC
M.)�mܴIA��ә��$� �4�Ma�W1ݞ�!�nO]��ou��zպ}�s����G2*q��}�o�s#����ِ�oe��ij��c�f��|%��ㆧ̎&��]��yqC#45S��r{c�je��;�� oY�}��@檟���>$�[l4̣:��{�Nv*�_/oo
�F	����'��eCx'6��V���	�5�����c_oJT�jj����g��Rq������?���o7��/�muV;�7���2�E%����~��:@�>ς�3��D���F���Z�P#���8ǩ_�w9I.Y���ʮ���2��:�������D�t\��[|�r3��5�a7���|vң�|8A��y
��������S��0#M0.�q���Ϻ���KTu��BwZ��0f���bZ�
Xk�N�����A�І�3����mF�#��2�%Q�{����ὤ׹��{Td���q)E�3Xu>0"��qVTC�6���QK����sv�
��k��{(�R$$���Y�)y��2i�կ������s]b.ʯ`���[�3���A"�İK��ȟ$(�x��~Xff�1�g�q��dw������=���m��":�6����e�6�&y�����oz\��p��nc�ܲu3m�W}+�g	�5	[����b�|y���g޻�ć�+�Hj�x���r�Q����7$c�U�_C���tS����Q��F�
�>�����be;��&��-=��e�B���mZJ1P�|A�&���%�u;J��*�5�.\�ٛ΁�t�����_�������*ӽƥ�#xj�����_\K�,�)��ʽ"3��F�ol��Ut�U���jn6�
mC�RTs�v(�#�H[wQ.�����Ȼ�p�&���b��_��mgfo.�l
��a����ڑ����bd�M�4�ϛ=��Ӧ˾	6�pr��م:|(N�ΞJ�(q s��)��l�+Fe�W-ޖƆ�uM�����DB�`�j u� F�G�+�{��r�.���P��g�\p�!��sw%��
K4��>���h�<��8d5mI�6�k�
+^�
�|��l���ʺ�x��@L�*�0k��ǧJc#��W�}��,׀!�;�rOA��%��4\�ǉ�<����T�:3��n��8�=��9M\H�qW.�{���A5��._��*�<J� wg��n�1Y=����%���LKA�}��:�]t�@7���d��f�3�j�4�6�q	������ؠ����#��z�N���u�)�R��4X�/ ��{�mh�S!��7j	L[�����S�*�����n��{U��V4㫗�_%�:�J#�n_�(ִ�`���wհꅩ�S�����.w}��N�������|//��sf�}/ tv�o\���Y��TB��l��F'��a�P�:���Eu���"�6�\z�\��--1���']g�-b*&:`��x�"1��|�O�$��8�`��vs�v���p6輈�KY��˚��4��fx&�+Pq�'�����A߅r��c�+&ʚ�.�[t΋�E>�cy�+�hN��*�֨ŽNK=��Uɝt윜�Z"���iw�w�u�^<^��>J���cf�e�t�KǨ)�$��[��t�΄[R�]���{9U㕣��<:G\�Tz�;�f\K����uܗ��iYI�
b�u�G����q��1�@a��.^��s5����U�L����]nf������s�ȎU�]��GY�O�n�.*�Iەj��)���^˱H��:au
�<m�NB�NoH�>'j��1͸�:��gc��ȍ9�u��*��l��G��Kf>������}�W�q?։�缍�cL�j�n���E�}9rZ����(*�%E��eY��X5ʚ���E�0�����:k��T)/6/�n�"�.ʚ{^_"��sތڻ����p�C׋6>�0T��3x�Xv��%�\�6�|y��o7��ȣ�ԋ��Lm�R��2odyf�H�%�5�� 1�XP��Rm��+�DVL���Q�0E,��s��>�Y�޶��a����ߵ��_A�4Cz�0�-}�	��s�����׺�K���{'�x��M��zv����ia��#nt�[@���(��gy�o�Ѳ��5�[���0gp���P'ݖ�Y�m�fv�[V�-]#tҨ�b���ۼ��|���0KƐ�䑑��ه��[�W��<���{��=�t��}�	����M��:��Y��"!��[�/aH�e�pI���C?��,� �u���jg&���׵=$�A�7]wt�pc�b�
����s��g��w��-J��"*�ݭ����L33T�Imf�u��"��6�%a�5>����7��a�,r��Uz/�w����-EB�+wZb�?A��ۄ䚬_��JN>��<��)J�6]��Wl�U�Is��N���?��K�%!��M��m���!.q�v���6���䝀��b���j�I��|�gK�:��z�ɱ�0�rOR���H��#l���>�>>>�]N�9%߰��ڎ�-�v��s8A]�� -���}�B3B�={���*Fݽj�w���5�mNס�n�KĶ�F:�-�Qv�õ�!�鬼w�<�[�wr,눥˩����rߎfH���	���b�~�V�����ń�ϔawY~���h\@S�&��Sn�|��~��JI�[��ݝٴ����(�����<)⵻�j}��N-�����m��jp�kn�|�c���q�Q��Ò���1 R�U��^'*�ζ��]��,hKI~ �ak�>�;a�B#��F(��'�=
��r���n�s΍{(�t�>�1,�lp̀�_��~��Yk\p��t$ԑ��͌����$L����e����^r�׋��.�D>�ȫ[UczK���+�F��I��j�'�t-�����
�32�v�o*`���U�C�t�<7u�����\)�W�/]aRVȾ�Oۙ�n���Z�VQa��Cm�I�a�" �S�C�M��1zq�XI[{��E�)�,̝&��;���`*]h\*��]g������=��ٱ����j�j�B�+�&@ŰA':/�h�so� 1=���^�֊�u����v�����7��cm�x��I,?�?�.Ӎ��nb�3Fn�t+m*ޏ�"#E��.ktB��]�蚓^�{�^v��jؾ��X�^�шGcB���yKS봊��We�\�Z��W�M��;�U�R���������m5�,Ú�s\���q׎��H�4���P���ا�咶�ENz�^1{�����>���q��7(盃|"�@l�p�v�{�G.UB�|�}/��l�mǙ��YF����!Wg�S��$�gW��,�̂�+��,-�X܈!M����:�7Z�]>�,���w}G�*��R�����l&;�vK�60�/R�v�y��zC�{�;t�ٳ
Er� C�n��{�R��-���/����b�ҋ�\�.;Jn����pZ����oz��n�oI���{�R���(�;�T;���j�x&sL���l�(�ӣE1��h�4T�*i�&�f�8�IƆ-�h���wv�v�u�N��I�Rt3*,�{.4��m3�q%w�g҉v��`ݤZ�[����+]\�r��n���X��7+8�u��m����M����Lnsne�����ù�{��w9rf��]s)_,�R�l�7Zz �S���d����{Y��5�'o�g���߯�۫�X[�X��2]]3��~q�����۬z��n�b$��m��B4�Qpw����I^7��#%glQ�gs��s��|�#YE<//|�"X���
[��vNU����Au�]܍�ƉB��M֌�Oe�$��6!�η�/4v������)�NIWpY=5��-N����VM�.����Z~=�jk!�����ʥ�:����xq�ؕu��/mvE·���[�R<;y@&��[����m��u`V!����w�L˔Uu��XԹF.�/[��e�	�<Ԯ���Mb��w-᭠�t
�4O�@�]�/R�����h竫U��H�� �ʾ�7�]{�;��0ɑ��B�_�"��{�YxcN��3���h�V�B���ٓ�u�!�ܺ=�� �f�+.fw>���V���"��Ĩ�Y�D��#*!b����gOTQ
|.r<~G��,N]�m� �i���ѩGȎR�Ón��Dar-a�Y��02��l��Ѱu�0�wc�z�V|X؇lJ�\r�;���ɪ�!��ӕC���Qcw�U#�`��m.6�]���_�yf�b�Ypmĩ9���b�I��������}���R�گ^�`�o�ᣣeu]l�s[�*������Qd#lk�)m���ݐ�����9ʸ�����o!�'XT.�7O.޷�݋;�љ��Q8[�7ի�>��.b.�����/ns�S��3��Y�ȋ�c��W]�Or���Y����/�J��#�<DAe��u�.�䝢+9a�9X9���Kh�ϫ_=]��:�NPrU��]������/�T:�v�b�oe�e0�E�u��.���ͽm�>��r;����u#���C׷�)i�鷸�꼥Pj�4_e��z��Ƃs��۪����R�9\#"M7)�y���ol�p��%Bwwr�?^��87�z���0��a���-��7�Q�9Y1.f�ufb)��y���[,$�i�Y��l���nD2&07�b^ix�g�u>�l����8˂������'5Yy�!��t�sPrue��U��j�{�L��m�(v��JzB\P���K�����7(��\��9�Ec�ݻ�Sz�y�� ��	RA%P�a�#�H�PC����]�cǯ�q�8����>�||n�$���߯m���^���禍����!�*!*��������<}z=z�8�=z�������ҷ@�W-��#kZ��|߻�������q�q�ׯ__X�����F�oD�����ܮ���sj6����[��^���y,U�\6�5�X��ۖJ�{W�F������Tj�\���NF0^��Ϋ��e��b�s���cݿ|��D��\�f6�э7��Ƽ޾yx�up��ۆ�*��^��AE˛\6���wy�����x^u\��wj4wWO;\�m�_(��O;|���}zzцP��a�	��O�a�0���j"LD(�C"����eQ�+�����[��zk�ߞ�ٍH�k#h�eu�9�>Y��)S땜�iK�\i��qX*��Z�/�[e�)�MZ�RB�x�ф�FF̐�6?W���(�C�D	��s���a� �)8�,"%z��D�"D��-H�n�0ce��~0A<Jg?{�<<<<=T����$ZH����q��m�+�Թ�0�Ǵ\���b=ʯ7`L�k�A����7�7�s�5��-�c����FvC����wy�����U��L���KgV�3ʲ��[ʙ����a��qY�Eu�\`�j��@�5鍀��h�k�*�[��U�<s}����A��{M׍���#�8K�\Q�>��y�viQ�ڌ-��������Ku,}
,���t6�=y[郻0;)��v2�w�e:
�>{���l�m�}����3OwXoR�����.�#X�h�O}�bߎ8��~��yKr;{�JD֡�bB���M�˷�(ǝy7uB��Gv3�+�&i�Xn�J�{$Қ��P�Z岔�,�Nd�灁@$7~�U������<�;�9�e\,�(�R8�p���z�^����,i;���|��a���A�3��X:{�ik�5��o��]xt��U�#w[K`W5E�uf�=��"H-��o���'�5��t�@s]Y\ 5����T��VA��vԥ���3ۢ�7u
ԝb��R��d�v�{;���C�<U��Kd���L������)�],^�K%�R���7���� ?.q��� ��z��!�e�vã��
Ƿ#Ma��wG<M��/����]�&� ��A�~�V��tީ~QY� ��� r���m�6sb�x�����wvi�^+�Q��9� �?H�]{#�=B#Y��u	9ӎE׋�i��Ju�{T���&KͲ�#ƂX�6cǶ�u��B�E�뱌gutd�Y�S�F�:��ג�<8ǉ�OH�w��(l��[%S�{�YͲڵ`d
���A����#o�$=�lwa�;o@ǔ�͊��o�6�g}��W���X_z^y&���y����TOt���4�Klrػ5Ϣ<�>d�H�΁�����
S~�[����<u�_��۞��n	�L�]@��6�s'�·(u�W�ò,��v�C2�V�kFon>��u=C�-��Z��e~���h��Jwr��\��5oYyr��B�4�EҞ�;(M�`����2���Ս�jw7�����fCw���}˺꾧����Ė8Th}��jeY�7ۛ`�*3#�P�d���-�s)��ej׍��k� +�E#�n����1��������~�Q�A�ww��u���v:t�R��A�S;Lqۆx�R���7F�ZF����cn|�v�ee��s��K�<�����	��{���g��Ħ+��j! ���������$���
Wg
��"�q���jw�i�ՇX��Z{�5�OCz<�R_��f���T�Cf�G!�]�� �јz7��=�p}Q�s��=�d{(wP:���WO����SrxZZ���F��RP�B=U��I�{����z؎��%�t����y>'7��V��$��p�].��]�����'2E����2�wz��	�if�<��F��l�r�r������.�*GT���M��Z�N��E�)��	ٙ�����m��c�Z�����0�j�gL":��do &��Gd�ఎ0)F϶�Q�`�m?~K<>�-�e�����������.g95 �R1�n��d�8���e:��2��?iZ�O���{H��YyJ�H�~t��U��8#�/X��v���*PC��+'w���G,��<An�<�ڃ��������?eL�A�$C34��.��QN��D6�d����Љ�RF�lͼh�/��K�8vg���Ǩ	�un�
����f���W��{H� �	y��'~���IQ�rtϳsI Ol�-��N[|�:Nޚ�f��+[U�A����7'Ǌc�FJ'�_��2�ԓ��3=����d�s?Y���d�D+Rp�x��6	9Y�Z�KZ�RA�w�P���j<�ԨE_*1�wM��
��l�^Xײ�t.p�;%��!�CȔ<�H��tl���|�o=���{�F=����s���Qw�Ea��{$i�ז��F�P%=绕P��sn%l�W�������gf��Ih������S��{�Cn6���E��m��<O,� \y��8��˵W=�YU�4ꭶm��Q�\9N`6yTJ�^�ڣ�����Չb�]�<�����b!�*����c��7\�H���3�{���+�KM`'3�>.�b�h�p�v��7��t6h���Wa��_7����~�PQd�{7|��z�.��s|��|M�#�ѯr����&��r��+/z�f���Ī�櫓(��50�5s{��[�p��|x�-���}]�8_�BG��g��n�!�Md��s�o5�u�Yk3�g]ᇻj��D�ވ�%��.�~��F~Ȯׂ����[hu�'w��*�Z��iݘ*�K$C�S�G�"�A�=՚�bs����}�wD��^s)�Y��hA�-Ͱ��?�����fV��ˍ��Ȯ�����;0��<���n��N�{��)X�>��
v�+b���G>M��j��=�0��;������O!-�0l�j��:�S,l�
w��h�٫���WLA�sA�	�{�����u?���]�i�����m��������`[9[��d�lvkg^*v�Fg#��������}7��8�L�ޮ ���\!��rn���n�]����0E`|��n�;D��=�cy`�ƃc4p&0rg�V"���|�k��KC�sBU\q��Nf���e.�f9�2�9��ӛ��f7�j��X%Ѐ]��6��m������΢��u'�7���t^ȏ���u�TEL?cA+�í���X��8q225�5�+H�]��
�-��'ZKr�oZ+�|��zb¼��D���?y�xxU7��Y'��v�G�A@�'ѽ��.-���gL��c����h�"�f�uF`�@�N�a���ϯH�hH�Z*�������lZ�C7~GL�(��f�~���fa�.�`����ST�{�V���Ur�V�~���S�.�3�V�l�qm�)�'O�8��w֕]�!�H���)�W����L�LnayM:��NP�>ʞP;r*�܍5R�VJN�����f�v�N���s5B�ݪ��w���߱�*�M���]���BMb�1�l�JkM�	U�h����u*�r��7/ת>ˎ�t/��3�"�$(�347S�= y��p u����2ESl�	4�-��uì��r��ul�k��VV�a^���x�J �Ҧ�oW��������� �.#s,B/Z�]��N՛k$�����DrέZ��[Wg�{���Hz����������u�����n��~��{�V|��F��M�в5���+�rܼ���'6���2�7����WX<���HWq!?k��]:O�V�7bN��k�/I�(��u�+�-�䖅Z�wa]x��Wւ悝ȕ��v�g9�k˫><bF1���w��{����
���^(`�����}2I�P����/S�T�n������W�O~��hق4�\�6���jц�T�E��J����3U��� ���m��o���9l�k���!�l���(eի�L�g����{{_�,��kσ�0�҆�tv[֢o�s������gҨib�-pI�c����i�^b�x�����Å�r����/wE�PGr5����_���0���l*�7��ý�G���ϙ�QW2*�Չm{p��_	���z�L4������[��L���U��w7Qh���u;sf��l��0�B�,����ׁ!��d���q��n�bl:��(w=Q�U�;"yv�\<q�ڝ��H'Cj�XT�R��[�b^��?c�'�O�R�52�;=�ɨk|����~�5S�VZ��y�����:4��W����Cw��cwi&ƪ è�%q�66pÃI��W���96�-�1-��`4Kŭ��+E�Y� E��,`[�]i�+�����j�/���>>o7�F,dm�-�Kvw�R���o�㺻�K���2����o�a�9.�w&��n�wx���r�sG/���].�c=>\P���3X��Z��T���u>�����}d��~�l�	@�Kܞ���W��p����jN*��,r���Q:w�%	��7��Jt���n�n�)ӈ�;5D��8S���ʬú����g�l�}�!���j_к��Pʇ�x& [("�6����"V"���'���[��{ �?�8C6
��.�֙�g$�ooL���*��8î�N= �t�;�I]�u���F��p�S/=�Ns8�U%���qL��	fox�+�kx2�Q�T��"U8MWc�Y#�7%�y�<�:��wG�S�rU�eHH,���̪�U�%�>=�b��ĉ�[��w���9�Zg�W|��͐nd4�ӏ��`}�yW
mm[���n֊1�4:P��b枭�w��ۿ�,�\�M;���HJ����I���4� "�$i@��π> ��G֬���ݳ"���ɳ��9�\��v��ձOW��q�:����ܬ���=X܏+��Ug��xxxW�N
���W��G+'nT]#7��s;w�$�m�vrA��='hT8r��R�wjGiffSI�޼��&�y~�9��D{�\��uOhfl�Xvi�]^����iD��ƺEi�/�^R�b�5�;�%檄�b3"e�����=��n�^f."�)	k�,R�@�g�P]E�x}[ʐ��h�[4��O�{��U������a-�q���Tv�Vrh�ou��Wt�ə� K�kzg��r'�
� 6�gwV�� ��~�]Rz0C�1
��1���ؚg:�w^W��U:lgO+���g��Ϻ�NsferS׫9��lϚ��u�+�ȍ�kт�q褜y��c�:B��wj��]l@���>;@�Y1�\8����;�s%�(���N>0�fqt�h��|%�Y�/%���%0��k���h�iOҘ�bw}��;�ٓۂ��܈<Ȳ�O�K9�%��}�~���v$�L���&�%f�{����"�<�e	�7/��aoK�ΐj3q1�uÒ�/ ����<�9�p�znJ����\�+���%մ��\���)�=]�{vU����p5��Rv�daRnڌr����z�e��jw���o/U��_LH�3�<���*�q���/��Jb3�#�0�{������f�"��3a�m];hn��5��yL3��ˬ��il��j��(N��ܞ#68���04��u��n�u��0��m���5�o���͊h���������Wzֵ�%�D����vt	���j�_r/�c�C�ݚ�Ҙ�T��i���>d6�ȧ��j����=3�B*KL+�[$�T�g�9�ƺ�ފ�&yZ�E��k˜��Xi^��ہ���p:W,Ϭ%�[h��Uf??I���`�H�C���r�Vۛ}�|ْb�V������ZYꙇ4XF���JkF�ݗ�T;�}bs]E['��h���1������8���uy�4,7P(B��=��V,�*+�6O+�����g�(qhbS�̭�ާ�;0Q�u3�W��������Y+[�N�6PF􅥥Qs�����M�f�����
W[��,F] �˗b�j�Ƥԣ���5�l���j�+��XÍ���,�܁m�����Uu-m��	�ȗw�R)�`�Y9�k��I	O��ݱ�-U�70��N��,)Kxh��M�v�7W=��
';C��h��*t�8ۛ����4H����&���n�`V�X����o_+�lj����eŲ.ɲ_KD�z�.�,)��q����떉�P�����r-n��ˤ��6�����hJ����R0t^G���6u]l,�6+�+7�\���v�gD��ܻIp<�Y�]��1�tռv+��Ir�:h����q	�6��ȗE�ɉKE��:�v�S��z���u��>qf�B�:Pչ����Z�v�@��P�������e-+q-	�Ná.Ǯk�,����"Xx�l4��C4e��S-:�1�����kF��5�na/K�Ѩ'����-��%t�O��0�RD�>���_.yպ�e;��,쫏y
 �ɹ܎Ŧcpm��p
yg����M�9���q�+�fZ9�Vޮ|�"��� JN	����*��Zխ���_V��P*"ϰ2�m�ɛ-nᡂ�ႤO:�#ف��W9�9l�f�+(>�}.�_����	��O�v�P�T���ʉ]���f��㫍*<@knG�*�f����|F�4)C�O`^��\�7�����h������pҡ��� g�a���v�ϧ�R����*��򑨵�f]�^U����[�@��ߠe�x�����c��Q�bAm�A�~�=jF�wKy�ݖ :(�w�r�\��{��ՙZ��wu�S����!�𰌽0f���(i�[e,-s#T�O��uʵWs�����b�ɐrt���e�D�f�[��r��	΃�#Oqb��E��*����žz����YhInh�{�P��֞���jY�E��Ymv�d�t���g�<J#М�����R�`ܳ{*�N@.�}[���Â�W��_8�<��Z�S�Ԗ[�.�)`����5kv�eU���e/3� >U㾪���էipd"�5��&p����9E���3 �a��(��
6���Z�z�.�!�SV��Q:=!�ы��y�/��Ҡﴎ�ڷ��ע��MD��!���gJMp���z���*r/k[�v���8��ur�� 	�uv����w�v�G�G���۪����*��1Iˡq�F[��B��v���Μ+�;��+3�.�zG�����k�ނ�Œ:�и�xs��{{�PȞڳH�T<�nEh�>��e�2��*Em����f�y����ىp���@M���b5��Z�d��0�#ĒM~WU�-��^M��2����8���8�8�ׯ^�X����Z�	.\�*]�f߯h�6) �-�э{n2H�)�2^>�v��x��q�z�����>>>4�0$!B	��=u\(���1���=��/KǷ���&��߻�~��\q�q��z������������w���M�$�W�w�v��#)���b{��	C�v%Ižwm��o}t���k�m���z\��v�G�nI��co;pz�(����˞�͗��#�]�b ����	v��^-r�lg����i��Cz�݈��\��щ���e$"A�9А�:����t�z��������}b��&4�]�C*=7<������ˑ�2%5!$�i4RX�n����u�]��̽����u��;h��X}ӗ��E�
�,�Fu�!��k\��ٷ���u�aO˥L�]n�;����a�3aS�I,��h�g�6�U��U%��;�S�n��S���ϻ�����pX�{۪2Ւ%���0���)�TJW��nX�|��6���
<�+Nr�a��fT�P*=��e�Ҕ�(��_$���<���t7b�[M�1X�CAb��0cdm����+��%����3�,�t�9;����z'��kTv���"3�F�.U$�׳lGN�L���e:4M���z��L�<�3c�i`�\m�GLŹ�%��	��4�������&�ǎNH���m� AffnL������?U�������C�R�������Lq$alyI�^u��XF#�{a��\�	��=�b�>UTW�Whۣ�KTT�b� ����M1���w��UdIƢ���bbR��J����Ԥ�'Ө��|��}B�.<j�=f����A%�X��g��2�n�T�}���r�aVc�׵�_�3�w(�vq��󠋣�Cs�F��9TLS*��^56����ޭ��$��֦M���R�,�R״��7�t��7Җc�Q=>o7��xx+d�P�[J�Q��qn����`��𸇻�QW3T�W%�7V��<0s�Ga��&p�:%�s�{���`W�晅b,����ۀUı�;��In�:���xw�-\��IcHF��-c_�݇��n/��u��Q�'韝 ���wF����P:�v(��zV���ռM��[5m0�Ѩ�Z[ӛ;�1�{/Őy�4���_q��ǹs"�/�[����+o-�7]�k�4���/ �v!ui(�?q�H[��ry�;�k��2�0.0�ĳ�l�l���@���B�ӻ�n{�*����e(MF3gnt>�=��z}�w�A��<z�W��GTQ�;|�胊������g��B�)�_@��!����.M��l��t�&H�Κ��{d�Ʉ���<���{�e^��|����W �S�XVb!�{�!M3���Y�9n�2��s1�]�b̧�z�����х�S�6n��ǽ��"�{���m��EL����|�( ��Y����}����r�]���f�T�!zzKF���>٢^g[A����z�ۻg{���XUbZ�s���{�+p�Uʗ�1�b�/��s��Ԫ��d�z��򴸾}�\�7R}C��\Bt�8���[T���Cr�l����g�������D�X�[[[�!��V�X��Tֱ9#�r��=�\�%��_Vj{�v�2�U��y��n�X6/ ��������o�W淾G3 �lwV��1�t�mD��Mx�o�]�S�T;�:��*�ʆnSU��C�kWUcө�İvj�W��Tk˙��q��p�z�w:�d�]g��Щk��Wz��Y��$�0�O�-O�S��=��ueZ��f�aVI�[Eu7���Z� ���#m ^Z������l='�0���54��Z!���Sae�V�T��]��ܰ�#�y^�7��"�vf�3�p��B��r`u��+�b���ʺcבt#�w����v�&�y]܃L�U7��wr��Ѳ��I�����^���-����׫��Eyu9Ϟ�8ع����]�<=۫��[���ÇR`�;(r�u��"@�X�7�ݫ�e!�Y��.NcY�L�ڑc��Oݞ(�Ib[��
Y۫�F�v�6��X;)�^n�3I_�=�������ڢ�CA(�Ma�'J����,���7&D6{��Iݽ�bok1s>^liC��{�S���&��;��8�����i����s����3{�z���+�QE���3�j1e陛[Ѵ\=`n�B���Y��ģ�ߡD
f�Q������.O)nϕ�-�:D\���+��C-�������ףy����L�P�S�״!��:-3Q�ŵ�|�5�i�O�W�q�Ed
2�c�h;��XK�}��؜���q���Cd�p7�G��@�HGc�w�u�L�5GX�����d�9$��d�l`8�{��(�sIS���ّ[�0�y���O�K��@����l�M���e�����w�o{�S�j-���A�/=@EY������۟P�3���t�b��_�]�]���M5�l�i)l����iN��g3O1T�3����k��%�9x���=�ga�6���a�Ы��.��#|Y-��n�3|��X�5��-'G�2�M�Fl{Vj�˶�l��'s�|��vy��U}0#c �ޯ��9��N��R(\N0?��c�8U^X8��JEa
A��C�1�2�Y����4�'�VV�+�� s���S֌��w]y��_��R㠹T��z���^
�u��îÖK:�
���yOb_5�t��������O��|	����L-�S ����LS�C:E�a8,�;6zGD��Lf�.�X����O�n��K�z����ż��擶{7�vu�ݎ�m�=���)G��ٖ�w����Z���sqE���J��ψ�F���Gle������P;����~�q�#ns��7"����v���m��h�1ew0bT��ȫ뎨��tI��g`����M�-���Z��S�{��0l��/�q��=*�i�V��J1�U�q鑴�~`�d!��p��vS�h�h���_C��d�ug��.����jb�l�ʖ���0eG���k6���A�����V�K������t%�2:�Wu�V�t��%�ǚ��|�oo�x;lt�Δ-�ս��/��o�`��Y�w�Q{��©��7��{��.c)7l���]�ViD�B�99�۾���iڟʌ̎-�h�[�qF �cl��/>�VVy��~@6��F�Κ)�2U����2���vuJ�������S�
F�*Rp�I���cَ�%ꙫw3���ּ����t!��t���@^�s[�ݣ�yOt7���	Ţ��q^L>�e���踉��:#�)5r�D���#��vB��re=�c=��7XI����a�P<;�l0��b'�n(��.��W\�Dqܭ,����kJp��w���)	+i[qU�T0��
���z��s����6j2�a���n=y���Ĥ�*��R���Wl�����K��W����+=���T��0>�6*:^}�{�K�����[���14��uu��?{=�ox0�3��ޱZ��d.�dyl!d/�"&�=�C��Z�1׏*����HPx8����3 �Sᐦ,P�/f�QQ��t<t�h-@��B�V��"�e�L�q���n-�erW+�l��".�K�J�ޗy0ę\���N�oip$}�<<<<+��S�������Xw'\���T��o9D�-�on��5�Θi�RG{�������?d>��<*�M�6OLfM���o���3~2;V�[fXc��n`ˈ���0��#������8�wxo.��ݽ��h)��u��a�.x�ȧ�\��͐�e��/�.a+m)�Q�*�y�vU�4W���Ɪ�=��O!��go�m�A�0a��ʑ�7_M��ԉ�]Ka���ٝ�*|��ݦ����C�Ed?�(z�N��n���������s���m�`�^ΓcǸ*p42	��0�e��.�7�u��3qsJ��v�X[�U�ai�	H޷�����&a�/1�~���o���[̷hd�r�K�t#Q�O-I>Ί��/�42�s3
6����l���J���3�kM-���1�a�"����_,+�5+xK<7W��������4:�a{��.Q��*un\}��qP�W]���j,]�c�5�-2�N�
ځ5{k2�y�WA�2���1�>�^C�<OZ=��g>�5N��a��|���
�ŁڟbkZ���`�6XJ��������7����a��U�s�!�boO�-wCw8�:�i�6Ԍ���WO"��ET�'Yy�G�wC�GQ�i��u���%v�?o��R�3х��&T,��4���Rb�Q���sr�}����~��}����l�)E9��ގ����m�$
h
@���D��{D�R�s����)�þ�n窟��{m*R���:��YoƜuC��V1�0�FS�16-�.�Q݄�Or�c�wh �!5xm8� �K"�(T.�Q�k+M����p�����f�|f��ҝ����=��d#0u��`m`U����k(����ݝ�<�^��W'��O)nʾ~HUɉ�I�b;$諼�D����˨�2"3� ���$���ĩʫ��6�9��9�f�R�"���� ���������ek�*�NFK4
�R���@<h/��\P�\C��M�[](��˾�ݭzw/Ѭ�Ik�H�p�H�6��n��Jڶ�&�0J�Ԓ��t	�>���������= D��U��Hn���}��t�%v�k�`�Y�VEf�B::�1Wծ�ݏv�ѯ�<*����y�}���V���J��T�����.R��]P&���9z:�V�K������s�ߨic��`��l�A��p&=��K�T��_OcV$\ݨ���j��KL��!U�S����3����W3�����>���E]�U%�^#t9! ��ye��wr&�^j�V'@����w C8W��C?�Ҹȁ3ڍ�XB��EV-�2e�kr�i��1CW�ԙg9��U2�5o��y���6��˭g��63hi/�v��8��0��Tiю��M�{�w��mO�wg�ai/��!�=q��{��T���ʬT��N���Wsj4�KD�1n��EF%Lk8m�������v��wPK��t�������D=M�mk�ڠ���,(�oo۰���JA�V��Q���n�Ug8��[F~��w�)m�%�}]7���{jg�|�xz�����m�Wt���X�V@�r샥M�}�rg�u��b+��xOIܳle>���¤�:����(�&�+3F��h�
zn�mMIz5v�yx]��+Ξ��#1�����h�	��ƛ��^`��O�'��>�'��=��_�Zy����QZЕ�N��5p�Dv�mэ����؞/����n��v�Ѥ��aռ{NrlN�mu��;a�Kסs���v����'��}k�8�n�%�����
�V^�_��!7�)�f�Q�`���Y:�v�
�<N�iD������lG����CtX.-?g~2��}��~7.6���%�Uz�q~F�T'�)�P?����k�y�}����J��B�_�����0�l^�E�涢c�9g����M�)LL�=�}�H�2� g���u���B��̶�n�5��"l�kVm�Q�V4oe������w�f(��Q��3U>#�m���hR"��V���AjR�'�C�ʜV��#O��W�^y�����_����UH� �� P�����"!���P��PU�PQdPh<���I�A��1�֘ɖ�c36�1�5�fd��Y2����X��X��kFL�S%��,��f,�MKVjmS[SR֚���֦�Z�Sj��i�j��jjV���5+SS��ږ������MKjjkSSZ����mMJ��ڦ�Zmf�5*�R�5-���MMjjj��ښ��ԭM��MM�jkSR�55i�j���ԵMMjjU��[SSU5-�����jj[SSV��������6�ښ����MKjjU���jkSR�5-���M��MM�jkSSZ��TԫMJ�Զ���MJ���Tԭ���jkSR�5+SR�5*�SZ������H���"�AB!-SR�55���MM�5��U!�PD�1Qt�� � B����T�5���kU$"�R!J�B
 A6�Z��R�֪��ڪZ�j��mU-KZ�jU�.��!@ �A ����Z��R�֪����Z��RԫU-M�Uݭ]�U-J�R���KR�T�6�R�e��Z��T� B" Av[ZZ�jZ��jZ�ԫKSZ�L���ZjV�,�]�WMJ��զ,��R�,���Rژ�kMKZ00�@F��m�AR1f՚�l�f֖3m�K6��em�,ճ%���s2��[e��U2�Z�����1�jjm�c�ً-��L�k��k�0<�
7?�D@�U0QD�O�t+��_��_��߷����?�G����?������wg�~������_m���?p� �������hE��H��*����@��	�"��������Ȩ ��?��=�'�vZE����'�?�?�N�
��`~a��$���hQQ�U��"T���i�Z�i�J�Z�Z�����Z�����Қ��-��V�U4ڣV��������� ��j��j���EZ�5Zԛj*ԚښmR�h֦mR���Z��K-���J���M-���*V�R�56���M�Z�eZZkR�ښ��m�Zj�T��T���Ֆ��֦�kSZ���MZZ�jl�Q ����~���������'� V�mm��X�[Ej��� ���������~���� U��������o���?����HC����O��U p??Z~��/�NEW� �����=?x}��D]}��� " �� �?�(?�����,((?�+�G�tT}t�Ҩ �?i����k�U  �}�P�������k��?�'��0�A��W�?�U ~�}x?F��$O�u�R��	A��4�����@�;Љϻ�PW�܁�Д���@}��a��__����E��L
���@��-�����}x�����O�����)�� ��RP,�8(���1]�y��(R(!DD�J���H� �J�D "�R$�U*T*�D��TQ$�*EA"@�� D����(B�B(�T�	"RTEJ���
��D�UD�@��B*J�
H�R�E�Ԓ�P�U*�P"R�Q>��AI�IB%%�UR�
AJ��*��AP���E"H�����%JU(T��**�I(�"DU"��T�T�)w�   p/+˩�-��������\�ݳ6���t��(w��TV�eX����[vw\��v%�f;%Mt�V�����K-����W[V\�a��RB��@H��*��   0�CС�B���(]���<�cm�ض�Uؓ;�n$^�B��Уm�����j2�Q�V۳3�3�5Y%���UW:n�K@��7wmXdZ]-���mӻm��V;vke��%E(JR�"EHR�&�  ���Z����+-��;Vv])�lݲ�:���n�w*T���-��Q�ۺ:���ggjn�[M�mkmӭ�9�Wu���ֱ�ۑܻn���UQ).�D
�����  �׭e4��E�J㶮p��ڭ7mkΦ�A�)�k�F8��[5V�Ү�UR��F
WWG[�5UU��f�q�jꔢ��T
�PQ
x ���ki�Vpu�t��u��;NW-�;5:P�8�I�։:\�s]��ws�) ��Yڶ�Uv��,i��؁B�R���� 6{�v�m���wU�qB��V��Svq�ƢEŮ˵�eW`��:��ەt�WMq���bu�u�j.���lֻkGr��E�B�U
!)I*��� 1ުH(%�J
P�U��Q@:�9u���c����aҔ���]�JT9���Q]��c��n����A�C��T�*D*�P�^ =�JMkzN�; j��'u( ���i;vJ�8 w!ܢ��LTR��`:% ��($$;�á�қ��T%T���R�(�x � z+�����;��
�U]�r�٠wI��PpΊ��E�t 	u�:pr 4l�Ӯ�]0��:R�%	������+x  ��T ������V�������;\8�T�]�"��]�w@ (w*��JJ�f�`
n@S�7�"�����R4#MhE=�	)*��h�B)�d�h�  E?��  ��4JUOP OT�D�UH ��#
�5Ȍ�D��A1Ux+#��9)	�0�/e8�℺� Z�V��������ț�����ֶߺ�U[k��km�~�ֵ���[Z��U��m|��������g�<y��v�b4�;Xk�h��$r�v����jz���B��3���1��� ������-�*�"w�t[�Zr�K�e�d��=�V#$�a@S���l�XAN��68NiZH�#������Ebá2�;�Zf�`�r�ԥ��04^SY�X.�Un
h��x�s�+	4!�J����]kF"� U4�R3~5�Z>u��2�!�Y��R�K#�qZR=jƝ���˫$����+I&���cb�(���M��m���Q�j�q	��V;LJ�2��B��q�?\3d���6���΃n��b���،��Uu%�������f����L\�N�54m�oMm��lH7�pۼv�Ɲm]���l}ۉJqn�Դ"Zt%�ͫ"j�/�sF�NCR��'��r��I�U �	�[X��"����Y`<���I��S5X�4��钄ٻ��q@JVtM�*vϷdq[嫆��t�5���/�G7Ð?��ٍbS�s�gm�b�E'i1���4�����e)���/���W�aЦȱ��E֍F�ΛU���*�سq�-��}��Ѹ�xU
����x�T\zNYݬ[2�udi�I�ec�SPRˡ��dQWW{S�B����2n��,^J �J�)�o.���*0��Q5u����`��y��ݹs��T�n)�e���X���(+�J�T��Z����:S�֌��2�I圶�n��&��7���Ț2��0�u�6K�%�ܡj�X�۟h`%eTCD�ű<��eF�̀Q��lv��0��])�Am��̷v.��V��u��56�jɄ�ܿ�&I�WA#NѼ��s(�G�m��{�E�t�-�6��	�f�jJYi;A�l�4���ͽ2eJj�@�m�p�+RAr*�����T���$��W2j��c�][r�,mYa�&dY`�g٧��X݊��=0�XY1h�-���^�@�7��+u�M�|X�;!}/������dD,j0���Ŋ��4芋��$����f��m��V-a�t��t�۔dV�5nC���%���U%��M��zƅY�YL���]d��T�yyV�������4�ə��5��+��4KN�!cj��k�+�p�(���-�[Wt���I5�n��SS�ɤU�2Gj�ǵS�t�t	gM��n[؝h)�0:`�,���TDn`�_#z��-���$9wj�[��CA�ȣr9�Ry�v�U�[(�mЗ{W��^)%1LK��y��!0	h;?mf�@��=ť����JA�YTp�Շ����q����6)���5	�j�ǓX�Z,�#P���[{Y�%fᘨ�j�Vʑ\� F�*�^�Z?\!Sx4\���Uw�淲�Z��5[Yp�Wj)Z!VVPu�vu+ɸVJ3	X�YK��A٦6��n��Gڋusf�^��wS�'Ɲ�/F�V�HG���+!�ҥ
��R�Ҩ,�8E���Fm*�Ȍ�c�b˪ڬXb�_�ά�p�:G�,G"�`����x#oJ�b��؍��J)�Y�jD�]�+Q��bB�]�	�+F�,�O+����Q��Z��)Yy�X�(���ǆ)�9��i!n�)�V3�tkxC���s6�4���],kq,Z�_ǵ*-�ܘ�Zeҁ��2��ވ��2��5A�	C5U�� �2�n�3]�L�$�f�	�M͓�	��M�ľ�۱��j:ux7j���&f#w3r��;�G@-%��J:(�!�?����i`n�p� 4L���f�� VD�4�{lۧ����Q-���D[tҽ�Ų�NEi��w�^��f�P�M�pTLm�<�5� ۔б+D�F� �*e޲.��1(��%���f!p�n��������B��O{I��0^k����8�ZF��0�ܛH%�
��u�� /R���eDm``��v��Vn�c�"�Bh��rЭ�Jdl�8���0�+pGl0��ܬ�/X�K,a�lS��N�l0�f�Ȏb�-�A	��Ew�VSn�f��.�7B�H"��Wb�E��&��*
��t1�ql�@�Z�H��tnPǉU���J���I��*�-�
�� �M�V�mGU$��;�t��� Yә,Z���L�Q��D%�I��9����m��ŲYJZG1;�-{wb* e�
Ͷh�%1{NXi��@�	Z4:�i�Xŋ�,9��M�D��s�BwZj�r8��ݭ�cɫA����ԇ�4�-cէ-�@����Ƹ�n��A�%�Z�"�N(����6^PB��o3Hu*�(��R-�m�p�J ̬[�l��B$r��+X�`��Z��
2��:Ħm\AS��YQ�����mmc��J��4墌�ٵ�)�x̲ڰ�kK��W,\Ս�c�ODu����4Ǘ�*;k/�t�L@�7*AX2n��1ѥ��.Qfe1J�M�)�i�-u2�ɍ�&� ���0�OF-�+6��*��2�@3�W*�OM�Tl-�2��]n]���HDWd�@��Tؽ��BfV��+�E�h��X�G0�+�o��I��4��1k¶�Kۢ��0j�tO� �6#HJ6iبU�`K��n���(����Z7C��ٶڃk7Z�2bu���R�@"��r	&RV����3n�e��)[dF�3��X@8���B���{1���'u5Z/4�n�f������/ ��z/m<�b��3��l�'m`�Bz����16o6�V}qRl�F1��[�m�N�Edn3z�<xf����	�4ȆV��t��*�i�����U�wX�%31`��Z���e�ë��%�JnƠ��b�Ƌ��q���ĊӬ^}�/K���.�5��ʺ�0f�D(.�����[n��/�k!б]��W�Z�+��QC@�6l��n%�t��	���h��%ʱ���Ǳ@5]'��0-�������*c[���
{,����W���%�d�\*eм-%���j�q8����5i����a%q4V��^�	[,SS4����6�(1m�אL"�T���z��*Zj*�f�m���*��V��7A�]��ÚQbAt����zb;[�H�SbF�Ni*[��7卹��.opX�yf�W�����e�u�^��O��ܹX6��՗MF7�5�1A�z�5wnX�lʌ[���h�z�KY�
�1l<�����-m6��1�tL�N�S�P�j�.�aӤ6���ڻt�AZ�[�\���i�[Nb�O�ٹ[Q�����+u�w���|�"}vp�ؠO8լWv��nTc.:�f�]:��u�E
55g�L��Y'.�PR�˂�Ǖ�ż�C70�J�D���"�,�!I|�z���/�l��T+"5�Eb��R��{B�(�����GAm�����X�����Z{B�y�c(m��2���HV7A�Y�Y�5��Lm�&$%8�I�X���sZǈ���{��ӷ�T�kZe���'�u���7HFX�A�g7*�ʟ*Q3.����fl�Ih��mT��tYUa�@1Q^R�h��un�n�QW�ܺ�9�b�Ɋ���w@��J�X
��
-��w�9�$ e	D`#w�u����r��F:vn*'Uۡ��w[KW֕4	L���8�i��{&�eme V�
���{��������^}�"ܨ�8�5wF����	=Y�r�u�⊊�օ'}�,���y8U�a*�9Fh�9S�6��h�j
;L��@�*�j�6�,\[.^�R1��!"�i��Cҥ72�ge�4#�����$5V��j]�Z)F�b�@�d)wx�**&�\�7�Y�ef6k�f���hi�+�z���Gh�)mb��5��7�n�����ب��c�e۲jLp4�tsA��cE�5;�)Ѽ�ͱ�VĆčCR�����6RB�V�l��:jf�?4fC�J}zԳ0�ī�;�e��5�%��S1�QL�4�el�s`����X	i�0a-�*�����2�cE� �l���ں�rT���A��޸u�o"����u�����<3b��B���B�J8�ַY��-���O���i��+vĔ�8���wbO�d�˫�xjº�� ��A�[���F���sYw�369[sU�o�7��ъa�,zce���.kJ�M=�fԢ��c��{�R����х}��%�Pl��1��=��ڽ(ӌbգj�:�\1�������j�e`ʔq'B�n�zm=Jź�h6j�1`�tK����M�b5���U��Q�K,��`v���iZg0VJ%V3Pa�d���]d0{�Ȩ-%aa9�/�sr��w�r�1�Ҕ���l�d�ŧ^��#Vs���:o[���wR�_!���ʳ[L�����YM �t�uv�^��v�En��P�u�Ba`'�ͻ�/!W��NX���� �z��@0]��ѣiX���Y���a���X!�>�U{����#�$Ӈ.�R����_ Ȋ͋h��/	�2ou��[�@P��֍���Ka3Oz�!ʹK��6fْn[�lY��@�]`[m�Z�A�`�����ZꚷQjN�`�m��ʰ�^��ҫܔ����m,f#fK��ߚ�h�6^ZI�@�#���in=�!o�^j��X�×�u�"�[�zr��LU���6�n]!L���i�K�������jmE栫^�+^��V����`3�Fe�De"�d�yFn�Xf�{�Q+ 0�M�	d`��(�ƍ�ه�=�r�bf][�(�6�n�m��d�Zf����R�&+�Ks7j%�&һ5Afm�L4���\�gدF^����HU�1[H�Ц�Y&۴�B�GA��-�mP���aIh{��7�����h�p�����P�Tږ�m�iKSIT�60����[��l����	���.��uj���אF*2-�-
.�*�byq�[J�[z�^)�*�ct8�A�)�{ZB`��e)p(Z�S�4J�#!6/U�SenV��-�[/i*���915��J���*#������b�X ���3�&L��]
Z��2��֦�SK4�9��'�"d��v����˻؊��A�TC��;`Ptkq3/Q�׸�����Ec���Nħ��tn̏�h�P��z��������6���4) �Ss~1ѳC^�P���/b���qSHPt.��?�V"�}y˶N��XW��W+f��ct�ax	�U�O5�k�Y������cǋcwt����`��&��9�n����LU.%�b�B��63hh��ƙDXL�8ĝ�*5�^�1e��x��-�̋d�n�b���dQ"�[қ�Y�pM�yE�{-�N�B�n�T�rK�yOZجV��ֶ��~I|�4�B�+�� �ax���SgR�T�PD7���و*Y�5&Ă�^2�:��i��[d,^�J��]9W;8�@+���7s%Z0CR��6�$ۚ�H���H�O7Vԙ5X74��4.�l;#�o�Hl�Y���n�Z��pm� Pe�(��A/M-�b��iNŠ���ڭ+8��Yv��M�T�,��3r�B��ɑKb4�"I�)�u���ϴ� �HW�b����Y
��ɨ����q&r��f��x�l��1������:�/�%�{����Y,e���b�ǸaZ�h�Qڲցɸ�Ĳb��P��g-]Y&�],�)�"��ӄm^���TD!}�����r<�y���J�ЅVԔ)dJ=aʂ�e���՛����ݛ�#Ђ�Z���L`�	k9%IK5,�V�y+F�ow/’!+�~z4�!�\�wd�`.ˁ���բ^��G�k�I�DT�ƠR'/4�Q|�S��;�g[�u����A͖Vb�(����@��V�'L�[-V�P�X�I��~j�*GՐ+�Xfoʒ�\�u���-B�@��sd�w2 L�Z���Ì���CVEnnd�q�5�^��H�HC�f��`�f�[�zT핮��6�q��XX��&k���q7��(�J@y�b�N�2&�be�BGQ���f�v�h�1*'wz�T�7(Ŀ��M�ЯsV��:�7��У*mXWn�!9���q�U�E�����th�DҶ�
zڻ\�@X�尪'"�/NTG5�A����gw�S+Fj�p��\���I�ܺj�� !f]���5����ө��c�wR�ʸn�%�}���yor�ǈ��!��@q��̭M����Q p`B��K(T%IJ����ȓU{���Aw���5� ��7,�d�t����K��.=�����w��S����EC�$��[�Z[9�$��p�=��-
;�B�4�5�Ա���%˘"�wCVBFЎ�Jj�%l��R�.<j��� �e�fhP�3$�)����B��j�Kui��Tl�����2)Ԗ;Y{��hi[�7lP�D�!S+Sزf�'t��R�E �e��M�.2��U�V�D�F�V��^��^[���i�
�6�e� �� [jk�ܠ��b-` =(��B��3M�����ٶu��N�[b��Vc�֪�	���{�l/�R�K�A(s,,�n����lP֪Q�@��b;���H=:�mf �ܫ�#)�o+N�3e�Γ@e6,2����u�G�'2�5�T�T����n�z��j��vE���n9������5Ye��-�Ra�O�÷�#T,�ջͼ�E%O�5b�S4q�ւ�G/W�ˀ]�R�V�D̘S��.Yp+�̼��R���R�9�X�̒�^P[[F�Xz��{��-�T�2_S�Y�LN��zS.w1�VVܗŉW|T��2�nݾ��t�չ'x���\2֝��K��R�K�Z��3�4�`��;���Ŋ
�J�6������A-�nfL57�g�����1֚]���V��/���K�V�sM�ٮt�b��r�n�kwrR�j�e�z�Ǒ�::�rK��
�u��Yɍm�bu�.�/��ch��]�,��;i���bΈ���Ox~��/k~n��C�}�d9f��Ȋr[kr��g�O ���9���t��{Յ.��jج��ҫm@�Y��6�D7��
���
U�����A�C�tq5 7M��z�
f>jC��0�f�tHg��!_h���qf��fѥ%!��d.���Oi��਴Fl��Q�(�3O
��Z� ��8�a.$�`x��m�����0�Z�U���Ξ�iQǰW\}h>�����Q��Q�o%B�����D�#��V#H5]��f��޶��**_`j���]m�*��nsΉ7y�[+|��G��(:��u!ݑ�
��6\i��^��15�(�/!�s�μZtX착r��e���ysX%�JI��5ϵ�:�Ɋ�`���ܖrJa��Uй]�q��(�٪�G8�M�%6r��邻��*F�V����f��\���r�^<�j�Μv�X��t4h$��Ϯi�`��N{��ͫ������	�I,�v,���������� �RW������HYt���V�D��1��wM��N��x�w0f��b˧�{\[�J��%Oh�3z����91�B���=2����cV*��T��]�6�c�W�<����>�����U��y6�E�J߻6`݈}�#ټ]B�]��L+�.s�)��Pķ�ͼsZ)���j���S�w@��'3�1>dk�h[�WB�!�\I����{鮝�fL����<0���e�F���u�:���]��D/;V�ǔ��IeK�vk�-0g>�H1��$�`R^��1n�yv�h���.�;��W3s1�ύG:Tw��$�J��:�!#�Y��Ltc�8 �����QnˊL#6�R�baX�\)��=X��4��~�-٠���JI�"|����ܠ���=���¼]��'�P����L1�[�q(I���^4�A�B0j��$NFc��K{��O�%ԩq�����^�u�.#���U���Ɩf�]T�*gm�=����;�����{�`a��N����F-���%��LXh̔�[��]٣K��}r�A��[|�[�Uy�V�2�{ ��z��:�����
|�K���d�&��"�Yá$v�y����f?����vǶtt�:=�s��vڸ���
�;O��>��¥E���P�u��iC��&�N��Č�P�����[ƻ��Ч�sE'V3"����,W]�:ZY��%0"���eJb�@�e��{upH��ѳ���I�R��,v=�Y�7�76<6�N�ףWGw4��Q����.�,eeE(���$�S����n�n�����5�/���o��b��Vx�F���ur��ղ�]��u��xec,�p=��)HjQ��,$�
B�*�3�ɷ��\�|��� &�:j5&Z�*H_iQ_�PO�UdPk/��c���.��u�i������ZǎqظR��ً\��k���K��RZ9LMnfXIh��o4q!�oem�R�kB����&]
�d��W��u:�:���&uJ�cNh��]8u���ti퇣OIU�ko�/	�	y�'ψO�;�ؕ M��M�W�o����u1��X�Bc./x�y.��XE�����un�̜�y}�7�wζ!\�Py��a�U���IX�n��x�F�]�\��Sv����[v��嫖]��9%\����T]~�~v�:���r�ѕ�-��rqwv�L�H�t�h�4�+�i�]�=ƅ��N�<��9�s�,>���p^�误��+�>e�cF,���\hc1a
���5S��nX�����k_j3�`�oM1lM�=�hg42������ܕ
���{/�s;���K���� ����,�WW��l9cmlYû�*�VM]���e��n�ow@I3FY�Fe1��,s� ~J/�j���=J���39c�3&K���t��n�JV�d��.�l�]P�އ����}>�+
w3���j�C�sfYIF�!}��
��Ժ�n�5�mM�ۊ��n��nT��I��R�;-��fZ�	��tv�j���giҶüF�RY5ܕ�W�ƌG���+z3�{��k�s��=ͪ�X�yW��
�����TH���d�g�+�N�<Y˞K�9�_X3�G�/�S�����^I��
*�-���f٤�=u�()�5��[FZ�^��sv�ӡ��li��k�*���&.�w���;��v�Bl�Lͥ�D�,��k�q���v�Q���vΕ����o���]�*�ܙ S����Q�oH*¶��>��uaRR'����/*����ufĮ5�C�$R�޼���N[4V�#P��.�P׉���aT���%Yy�v���:������ڴ��kš��r%�FZ��k'D����k�J6��e쩦䎄�����~�.8e��i�2� �R<HNZs�E��:0��8&f����6� �q��,\ή,�*a�a˗�\p��lF�����K��病0�
I8�Ƅ��[�2��!�:#���L
���Z�먹���nC����MFp%^S�/�H6�6�e��V��T�0�k�����g�JNΡ<;��5iJ���x�}���۹��sے��ƕyS�#Ɛ�]}J;S.�M�+k�U
P-��3l�1t��:AN�]���x���y}�fe�����;���H3�F2T�W*P�X`[���44N�Z�"U�!pR���]ʰ̳��Ӕ�k|��{�fn�f��љ��ϊ��{WV����Ft�jy~�=��e@�����x��<���e�������v1�Z�S�X8������)�O-����X�oufD���:���`���+t�e�t�gh����U�ycv�n\�ɜ>ݵڈ�4�b�RN���ڠA�s�|�	�8��Wj�'&�]}�uMT�a��c�g�_ʽt�vٱ~��~�$�}Bf���`���i3q��
��"y�.����vn]��"��r�8,2��y��ͺ[|F��ݴ�S��YOD�m ��6,�,��ƭt4��_-�|����F][�N��������Zd�[�@ɣ8�lw
U�h�P���-��:�fsr47fQ�y#���L��#H��Q!���J�hR������ӈl�Aa��`8DYtZ�b���8P��`��J�`U�2#י�ېC\���w05E/�-��Gw��Āe�3AaV�73a�5��
qd8a���j���,X�L<�nu.��D�
�ET��N���:V�R��#���]�B�-Ϋ��;$,�����K��DU��Juj�{����V���S�c�s �X��r��ւ�3*WG]J��/�c�iQ\�;�oM��Sy��{��u���:76�&������޺�T��J�`�5iޕe��F3:�l�y)B~i6��\�Ķ��ԉ�Ҍ�gP���,�P]���Y�G�?��T��텯gw��N����*P�0ZhC��R�k$V�%��G��]f��=�/��L�5���e���ڄm�� ­���z��� ��8�����ΐ�������e�w3����b�{�@���5vbL���m�C�T;/5ج�����N�����ݍ�{��#��$�BMN�eLZ*8����p\�����óS��"<�y]��������56q��psl����s �ԝ-]Hʤy�N�K`�r�'yf<wZ��ZxI�΁v��ࢠ�,o\\g^���R-5��q}�F!�8�2��x QR�U8%�Zv� ���%��E�����d�r�C㈵�k�]�2w��Kˮ��k�X�X�,�Hq[7D>
������#%%vL[�mHn>�w�*P��RN�ڶU��W'J�%T/1���\�]{SR�6�I:6�y.���F���K���2!;����<E�n=������2_e.jage�F>.��#g�[�ð�E>,:B�WeM���jke�A"+�bγ94��T�=&�6�v�L��h#V�e�Xw�j�p��M�mM���Q-�Kd<��d�ݐyw�K�y��#+)�8���N��5]]o �B3�v��e3�6��gL�9�%�J<p���?<�F�U�ϸ���<A�[�<f��{�d�]ٲ����L����� ���7�#�+������Ki�R�{�k�1fʽv���#��*=��i0�u��;�V���W�pfN�T��]l]��E�[���2/�i#�e�Aһ@6K]c���Z�`W��z��N��k�7%�|�T�m4�=���maÊ+���rdtK/h5��k��Q.�6���A��6fu�����_jy;�;�(u`�Z�0BoI�Nہ�]��<U�fv+��4�� r��p����_��+�m_U��p���A�4�<b�^M�cPM�r|�ݓ�v�®d����pV��iuHȼ�D�� =f�zWrޜ�o4�;<5r�d��Nz�A'�&,�aΝ�l�Ȗ�Rʆ�:���qf��a�.�ZoZYU��]~��<-l�k���ۧn��]	qN���LX�DV�n�*��7��k���[�Iw9Y7`�c�/�� TY�!���k���r�U�fB���M�2�;����/��
F�f���P�Q��n��ZlB�����5�[�S�{KDj�掃Y%�l7�B�����r͗��o�W�IV��P(p4�VNF�!�l�Ɲo�w-�
`�X��W�r��M}�t�S7�X&Zϭ���,1=&��Ȣ���a�ٹI�*�I��m�n�7�[Z�ە���o���fK�B��x.JV��S�gou�t��+'�f6��@���+�3�Gw,+~��rڛ"�WKZ`k�A)��d'V˼��%ì��H��j�<?.]V/�3m�Avݪ�8vЖ�*n�]���L��.�U�V�Y6؎es��E��7-���x(��	׹���H�5�,�� ����n�� *��U��&�d$��Ւ�W�k�߭�+U9O%��.�ԥ�g	��]��*�S�wR��9��t����c/�wgu+U����H�ۏ�%6�Q���g)P��E��={M�
�V�obڔ ,_Z$D��>z,�a��ǝ��&LHl�t]Rv�-��s&d�:����\���rY{�"��� 4P̧y��1D8�=/��rJoM�Տ-�dD����d�r�b+4�ޜ��"�a�Y���Y�pl�Rk��]e���&�ҹ�:̇-A:9��rJ]�n���N�.�h\�,��Ʉgi<1.�[[�t��v_tdL��u�c�{!yxF���iIԏ`]�_*�����9��JNr���Xrk�򥫨���R��E�vg#��}������6Y�J���U���عAt!z��%�����W 9��&��'!��V>8-I94�:���4kߕ8/�Ft�[��@$;�u��fN���H_B0Ă���n�v��I	�-1^k���(�}���ws8`/��l��h��-�����TN�&��e9Ƅ?LL��u3XE�F��*�Cc�[�ڍc�W�^���^V��������gDO�i飅�V�AY���J�\���rL��h��eIWب��*��5�iMԓ8��,p���U��qI���-�ճgg:{J�C[���{�>��m�ƙÕ{�i�G2�=/�guQ��q&�"��ZyFn�V]B!2 =@Σ����W;;�����C͋I����_M�	+ ���&!c��4�9���Z�qC�^��_5Q�6�t;s{M�iȻo۲O7�BPt�6jB��/���n�zE��+��-�+O����'{�t]����'J�Aw�!�u���3ZN�W ��cÓqwgKU��� ���>��ڙ.�Ϯ*J���;8��e�q-;oM���$�0PB�bΧhd�kZ�2��K�yn����w\+䋊Q``B�����2�Ρ̭ǧ'�!�kp��ls��(�t$��0��V��������Y�r��T��nh�wxr�A���^P����<�˘������7��2sk
���(r��+
G,���n3mN�7[umw2e]#�9��>�'f���D��kjl�oN�;��c��P��6��=XUv �I��;u��m���>����%�����AF�ۭ;�k
'���Ȥ˭s-�:r�Æh��)5��+{���,oX���ָ������X�++�1�����,Q�p+a���}k��ٹ���et��Th�bZ~4s�:�������O�Ù�	f�9��� �X:���2��s�.���y�����!��\�O+v�>�Ɲ<����ft�U���>�5�H]C�wl����%n`��
P�:N-�/��s�H�':�Pk�P�t�V�>��;gA��S&P���o�
L�4��B�r��E.�t�������._S�����������p\߇s|1�UL��K�W�+|b]b�U���3I=�N��9%���`<��k��ޘ\28�śE��������Aӧi/kgU��޶+r��[t�K�Y\�V�����Y��^Q�oz=�ܽ�Ө��|����!�Kȅv��[vM�I�����3˻�:M�8�'9�E�K�n�7�i=�u�p����,����;��N�u^�`��?�"��η��ғ�����a;�z�]�#����}�(�9��=`n���{	]�Z[��L=�o� {[���KؐV�yj�f��B�	�j0�$�(ʚ����j�� >  >���}�����}���R��o��n���S��1�C6k�j������M�7�D�$i�h������ЇK1���F�N�W��+�q��ڦ`�G(�U�Ѐ�5�M[�˝��f��ï����Ix����	��
��LEq��㗌
�*��!K 9uø�`}է)P"�S�"�x��JQ�V<��L��m<g-e*�����Q8a�^�TE�Ո	z��mn�ڀ�>n��z(�����]��׻�xJOg'\�Y:�P!K<��D@\I��ĸRZ���m�4�nV ]L��J�J��J�5�n�u\e���P����Թc*]�E�\���ܙY{}�b�
��QA��)1&�%AoSڔ����B$a	�N'p�k$�Y���7ہ������=:��/3��Nk�? v�.@A8�g��yn�1O���]�P�Tj�<7�4,��V��L�d��{R,��k�m�f�>s��Z�C8��1#���]մ�l
��,�I]�~��,������aF���Z���SYvG&��d��J�q+@�壘*:�GA`�ֳ�w>�2|�)�))�Gŝ�!���n�(�v��E#w����XNP#*�·{lj��T����Ʒ�tZj��J}�e!ц2�<Gz]���p=$�&�4�.�Z�k�Qy��y�ж��4��0&	�5|�b�5VIې�9�"ͥ�6-���m�[���u���I�u��vwb��4�V����m��F��p3M��1���nr	bFk�,��59dK�Hrxlӣ��d���1��>���<9H���8�n�B%�V�+pm�wB��E������qI����'5�S�Ȯ�w,<fv"خT)���_h6��:1�y�x�%��Pf�ӓ�&B�p[Y+Wfɹϳ�LC-��웶p&E��lz�kʏD�|{A�2���b7p�[�^U��j��Y)K���,GD_e��e�a<�O>���F��Б*݌��㣎#/�&��0�)u]7��aK�M���-ﲅ�/��-S��X\^'6���M�Mn����51f���i1c�ذ�%����B�G��&J3Y�L����6�먣!t�Z�]������;)��G���Ky9+r���V�&-�ԣ�*�Xu�� GoJ�zJ�	�ُyb.�U�[T����k������*�:vRt�l�c�LĩgX2�l�$nr�hBv]3܂�����ݪ�EU�\��>nc�D�+y�b��ko��5f���-�c��e�+��q.��u�穴 �F�;W��F�V%���;V:�V��K�G\U�YjO�v�J�yeD�M�l?�-[�tgYׂ��+M�zLT̷M��^WM���1մu�Ħ1s����6Zx������/-�d��fթd˽�d+z�u=�P�WqI�>�5*�1^��.�I�G-"����X��Om��)Z�Nr���	R�p$����=�6���XP���J2�O�fq����*/6P���dj������w�i��s��cYN ��!t�
�B�g+Hj�1�\ ��0gbN�iG�,JM�8��4rpQR���ѵ�oZ��+���9��+�X�z;��Y��B9��}u��.��2K{�P���H)w���s�F��n�C��T�M�&Ϲn����i;�\n��U�(���&T�_i��<���2��q��'���r�-�ˮj����5{y�&x;5 YYqCk�?qX�"喷uZ�aꏙ�(�9̃��,�JR�`�f
[W��h
v`e�))|���(cy�f��/kS�U+xl�E g_9f��-�ƞ�bFiZ[���BĔ��yQ�K!���wk�����8{}�r����K��%Z�Yײ�gK��еg)c�6��Z��P�w�%�]��yx �J�X�K�n��g>�9�x�nT�OkE��|i!h�ejN����A�Y����p��C&��\Ьt㛸v�ãV�bb��:Xn	��`]'��d+���c)���NU�GnȚ �,��OR��L}�������ඕ�{���+�|�����뺦��k��s�&Tfn�mH�&RZ�۬�X}/�·�WH�%<��e^M�Y�;�5m��C�GZ�VѡrH�y� MLij�G
�Z|7��ڳI�o*�����[�t���;�/Ue=\nҬ�0�"�ưh�ktp���y�>_k �Ev��	
Jup�6��s��fm��b�l� �Zj-޻<Ev�G�wB兩��ӗ:�Q�z��
p�@V��T�}).٩RqX5t("vl%S��t�˕��qI�FQ۳�ςǇd�2������j�X��A�6~0Q!}A)l�Q��|Fql�A�i�Pb�.�}2�m$o v���9�oDzf�*��{��ݝSI�F>�;�M|��i�;NU�zF�k.�pEq��ǀT+�"���� kc�<�7O��P[��\���������ts��-I*V�l�o� '��o�-<8��3j�
���ޭ�hh�Gau�@�� =D�[y�(	8�E3w�t&��dB�O8*� ��I��1���5ʘ�;Q`�.���s�,����i;U�Wh-򂥛��:�V�LBނ��Ѯ�s�Cr�靁U��{C�K�y�vt�\�V�{��d+�B�Le+����r���)n�-��]�[͈�­�&���i��-�=Ԝ}���{���7��|�����s���s�:�hZ+���lXT�x��u֫;.�
Am�f��2L�w�j�`��RJ[Gxұ�of��@Le�n�)ָ�#���W�W:Ϸk�o#euJ��(B�ky�y��:��.PК��Nqe�S7�M{�3�����z=�c�:��5��P�ۧ
�SL�������oN'4�ھd�9�;A2�=�W�r��u���M�ж�PM���T%*f���k��ǩ"�'Ñ\�������r1,��阅��ro�î�$���]��E+��@�`�r�C�갥E�./_P�O���+��˂,�5wYs=N>���G)��;wG��vx���#�.g4>w�\�.�֎A�e�����۴�m��b���e-ڗO	+BX;z��M���-�v��l\��84Kէj�M�`��z�A�K\�Ԉ��6�ե>��Åv���E���5c��CnW$�@c���uY�o땚���._���m� �}����ﯕ�-�ʛ�vȹf'�%�E��wV��̞����y��I��J�A4�"����í�s�l�knV+�ȩ��7���ٰо���pǆ�
e���pN��qG��S,vS��x�v!���%�V�9?��ް��E��|�Pu�|.�9;a�/�l���nr���)������(`����Tȏ>��8�x]�,uvc《�Uƫeo�+Y�����9j;ڦ�]u�,狭�=Ss%�Q�ỶlP⳷oe_u5"Q_4���$�TsƟ+��:*�)��M���_���Ϊ�'��F�=tz�oW��]�x3CO-�@
��K��0_�r��[@��؟c�4�etٓ��,��d(�pF�9]q�5�:n^�ً��h���X�ίZ'.��0M�{I��zwj�=W�����j�y�:�,���R2�e*R���+3�J�,��)T,l!m�s�v\�y�Z�>��8��,�6����J��GL6����y�]�Q�N둥ݶ��s��'3�6s%)��p:y�:iM�E��F>j�����{"po+wWu1���6��y]m���1��pJQ�(���jt�����B[�i��(���*]�(:�ܥ��#�y��1��ӵ��h���|�e��[�1u\�5��I��$��0H�������i��c�ֱH�1I���z�ft�2J
�{N�a��c��`=[X�Û3�����f��0��5 �f���Q�ì�f��}[C熱�����R7M,.PDo6mi��Qf���v�m�� ��n��l��C��tCm�"v.v�3R�IԒۼ����7��&��oi���̓`��$�.�*vM][��Y\��5'U#�9V�-2�s_l���Nj�]׋&�d7Fm.�/�;&M���EM�"sn�X�;���v��b���e *�2>����as�t�ʇ[3v
���oU�Q��FP������]�l��E�"����,]��P7MG��v��� �=��ya�d���\�
]ՙ�m��َ��)ϋ��ku��$|$��#�>O[��U�]Gh�哃��Y������2�`�s��q�*mڼ�g0�:��5.<�ʘo��Qa��!Z���A*�
OU��b�����^�n���
{�B��0��]�,�p^!�ݮ5o#N�K-��IprCu��Η�m�(��-v��Yi.��Fvs��_2�6h�'W�ghkm�������Q��w۩bH
��f��X�;/5�p��-�څ]�6�*�&�5��٠��Y�ྚH;����X�X�B}\�*��Tz�2�'�Q�I��64Xy��e��+d��S;�C�Z����C�Mt��_$Y�ܦ1�)�ÜW[W�,8_*�ݍj�ؾ�0c2v]X�
�shkt��u�E^�
�S��-k�v�zW�a]oH�b���t�l4s"���*�ˍ�f�K]o�VZw[X����7�EU��[K3V�`j�7���J��nM�2�������VڡtE�w���M|u��u`�c�Wm�A���bXu�ZA\C�Ea����`�Y�W;%��f�5l�k�(i��Zo�ͅ:���&r8۫�dN�337oiI��a�'q�!#mZ�B-�w����r��T�x%'9��\�u(�OVTֶ��S�/�X��v� Y�v����6�}x�eeGm��s�[8���,�	�E
��j�s��o�L��x���A�\��c������\c���'6�[a
4y@���%Ϋ'ufjs�_e��@`Fi߄Ó��T�����K2����m��	p�W�1�iY�w�bf�r�0r�p4�6�^A���s��к<�뵷��.��-��]ȑ�� �Z��ʗ��UZ�Jرv��pcgYt�� 9��V5iF1V�nne���[朼�C���g9rQX�b8K�p��)�����'PYjE�.DD����Rf�Z5c"�{1�N��z���9��
}����(�ݑ�MX�v���b��X*X�-���V���o	OoW;��V�-PK�+��oE�n�H��y��6Y9���4+]f-������n���u�Wr���p�)�ρ�[�ܭA> �}��9�$ܛVc���3�^�S�v38���r�0�����R�#x��Ie�����m����FS_^�Y1Sޖ��{�h���e��3����-^���VMu�<����{ZS'�gH�vm]d�E؊�"�e�;W^h�L�&�S���]�[/>��;����d��^A��5[i
����l�	T�r��S��j�S�d��h�:��5���I�jq���we)��@�$�=`R@e�u�G�fԩ��SQ[Id jeZ{:�h��W�V���"�K�\^8�+\��V9s��++�Z���@c���б�z�������>�㴜fv'�#դn�AX��sJ�\U>D��p(��B�cC��B��z7�JQ�WFڱ��w�;$�P���dQ�6��#���6�p"���c�̽�:eҒ�h��8򻭵I٢CM�,�kF��
p	\S��G��8�:�I軁�Y:�;_*�P�|"�Y���7�øf�⳹6�ʅXu�pW�ˁ��c�}��`�o�Kvd�곖�������7�)�8�7������n�J�>S4�N�8	t�Pd֮ݮu%�����aY�6Cn�'D���x�Z��tn���7+E2���*��ǹU��:��Ыqe�v��B�U(Լm\�7������h�GO+(�G�+��nZ^+X#�V!|��V>z������Ox+��d�����=�l=�\Į�d5`P�ݻ�a�]Ʀ����r��K���є��X��aݕ���/qjw.��v�݅4 0X���ڋ����;�J�n�%�p]G���B��v��7��tb�ZZs0b��kv[�8;��r��������*����8��_0V9��^�GI�����#r8�f�{	�>�@]ѩJ�5]x��
�Sp�P�o3B��%����n����Z�f�Mt�C����p ju����.�
@qdX���h�9TWKM�T�UE����;W���G8�;Zv��9�rba�n�o=��Wp=��l�SE݃1siS��o|�p�b����]YͲ�s�ٱ.^�d�X:㕧N��}X]�]KHv�����t�tʛp���:Ņx{���OS��5�)�G���t�c��zˡf�wj��V:��0P%��m���l���]�9��EF�\狅M�V��� ��S� �efe�뙧�oA����&�DG9
B��*��O�J�X�D�aN�u�]B����l�6|���|�&é�cI�7`Dju)�ahu�LVh�D����=�/m��R�O�ی��C��6�������M!��4��mml��6.��f�ukz5�#ϝ��S9w��nvm̎j��(�B���#ku�M4v�Vh������=��@Ug��&e�
�]Jѭ��2��/M�@]�ǁv��CMϙ��E����Ӹ��&6��r>�]X+����u;��d�؈����щG�|�u�좭���7�J+�F��Vq����KV,NX9f����5x�����ڦ+g$;+N_��2�M�o Z�x��g�œw8<��5!��������yh���R91�<�|r�yCzՎ-WL��7gNq�������}_}���DƠ{Ȧ�t��0ڕb}����t�A%ɬ�Fm���t�c�!J�.v_)q�ua���RW!�sP��9+����;�|ӊ����:s�TN�ܞ(Oc�v�^���N����e�ͥwۚ�YC�3e�J�y�{��B�%9[������|U�w��n:�����3-���̶�4�5Ҙկ$Pq��&��,��(�-��k(�b�6pgN6�v��r�*�����>N�yX�X�/2�gT�U�N7�g.���������Q��Â��f���։H�w�M0�N<��.A:�a<�޷�j�5�U&wX�q�=��щ�x���̳��tz,}�P�<��
�}s)e`?F+�q�i���I#�B��zW4r�M�2� un|�6lw7�G\�D8�\Źup�K�l���f9q�<5}gzN�@��Ӳ�w5�ϝ�FR���ݫڼr�\� 高�3�*O�R%�X�uqt�Ly�\|�+]�����E�88��!���0�֑hm�N�X�t�+� ����'��h�X*���S��}���⧦�LgP%��Q����kR�n����:N�u�
V�c�L�N�++9T^����ꮨy��� X3z������m�[-�wn���0y�qM��V�~y,�k)AV��]��CF͉�U`_J�.�E������ڀ2��F����)��'��@� ���(|`$F�"0Y5?{�w�ng��$��sBcXH�EL���$4Y(.mp�ۛ���L(�#E�+λ�8�H��cox�sL�ix��uΖ"4��*Er��G�\�3	II*yۂ2$��cD]݈Z#��4���ܼt!)�v6�s�!$i1��� ����u#!��3%D������#	�ni�eDɠ�^u�c�"��a�]�r�W�E�Fk��`�h$�K�t�
#F���E$��7Bђ&r�D5˄�J1�$L�w'��%��3bb#"b3�4x��y݈�&�"��SDJf�t�.A���2s�f2�RQ.]C&JH# JJ��be�)61I�۔$�BL�
$�K�sE1��뤤H�"�$bwUٌ�����&���~�����ߟ���>'/��]9!��5aw�_pc�7���.�V��A��Ѵ.���0K|����Vm���c�DR�ލ���p;�����ݪ<f38�}Gq�2�����E+ιR�u�����wg_����=���Լ�v3��1��=Vh-�^G�?{K8�����(v3b�ڽPWW��G�P�����7a)��gw�� ��HOg�Ĥ�5�Z���k�t�������<�gVl�Ʊ�}H�.��r�����#���_0�(_4�z�	��"�x���	�6D\�p��s;��Y����vr��Џ���ig]��ȩŁ<�G��m���w���8a�3f��3Y�l,���T�{[�Yrr$}xp?��n+%<���:��3�kk��C^-����TVhĳ�Cb��o.���������o�ُ�
Vx n���:�d&n�f�QT�Uw�-�&�?�����N�T�qW���+�hS��φs��clG�j,o���{k�q>ڐP�o��e��;{EӠ���=��|�)��hT!��s��f��8H\��2�ݼ>jK/�!�M\1eM��'�iIL�F�����W�]����@I�X^FS�p!6xh���t8Ά|
�z�VP�Vg7���|����֌ғ��/(���`�����q��|�%Ƀ���Z��ҳ6��Ia8���+7�1�fS����� ���r�>[�]vu��uїË�\�kij�ʀ��lS��h�ٹ�3M֪���"ǅ�X�#�k��Y������.K)AUe��^�D �����j��^��`0c�e�5�
7��H�����F�ўn�I��;��&z~AFL�v���o5�]���Q�l�"����`�@TX�Y^ۂ�� ��#!���Q=�X�\�w���:��j�;�*��8?����F{�Q��7y���
C�K���;-��/���
p�`�E�1�%;�	Snd``v�O�{�_)zq���(��fZoAuwW�'�t�=��s̙7	�_���*6~�']Xu�(������BmZ�o�g�q;e�{��k��S��g�N�.�u#�I��+�y��&��V��RϹ�������m�C�W**:(����5a
r���]ZTPpb0I嘞��޲Q�Oz����٬ƫt����V�x<��*pJ��hȉ�[�U�7Ȳ��3'�k��ϻ\lOo='t�r�c�Ҋ�?��N�L ����UP��Q둚(z�R�y���}-C�0j�C�� �-޺*׮x��uug��x�޽�ѡ���笍-�R����vg�W��n�D*���^���N��iL�D�>h��tOp]��뇚۬�`;�'����Vtn�J�Ɵb�Sp��C��q�u1���o!��z�JF�; �<�}\ٰ4<Y���t~�{,��x(�c��Ć�Ɔ�ia��JxFٚ����J�x�K�Y�b��Ŵ���<�̯��оy��KGM:'�t�Қ^�\=k|����g9�sG��`��Y�'ţA�l���W�@�Ҁnzf�Ƀ�X�qR��.��J�0S��J�>�4!\at���-|�9Pڸ{����m
���!{�K�E �^���v	~��
�E��������������/L7�Q˂ƃ������N��(���n�1�f��~20D�ܢs�cK�=�K)wJ�+�~ӞÖ0�u�}���jsWy�)'��_����M&���( >�`�P#
gj,+�v��+	��+���vܧ�B���s7Y��4n�5�P&�D�Ѐ�'�j����Dv	��.��x�0#j�z�e�d���n	=��s1�d�%l3X�;�b/7D:Ԉ�pp�'Ļ�[w�ρ.�����B���������g���qB���B}i��,�|	�L�����Z�[��(s�6NVz������,�Sv��v����쇲��C*o�m���A�^�s�ZUw4s�\�]���eowrkr�ڎE��μ���
�LX�7&<z.¦�W��K�W$s7�R�^�u�ov��lcy�X�\&K����a�{�vj�ՉT��˔k������wt�W2η, ����_����腪�-�v��Q���\H�V�,�וٌ�f.e��+w�
��c�=��qV���D�\����D\d��P�j`'06��Am�tվ`���ҽ�	�z,(�%���R)�[����eA���Z�m'�=���И��(�g�i�+�Z�X˟�B���y���=5g��-)�ٔ˕�b8�:�_e��;*�Ȧ�9beŨ����o�oY�Uoc]����x��x�_==^{�B�\��T
����!�:~P3c|F�R-^�f�!I��+N��
>#�m�=�a����\	�gl&�A�-�*m�\m-�
y<�^�Yw<_�D@s������Ji{J�t$h��/:�x] �t=5%YT/(x:��pH��e��]`�%�8�'Q���A�4�\o���[��څ\n3W�.�������dkэ�@[�ѥ���f�� SRt>�$j��L��O�<Q���u�ygo=�-�w��8��Mx�*�]c�ӳ��Pӽ����y]�����^\=��m6&�tӾ�TM�%����-����P�+��9�ڱ�H��v�,�㍭�U�y^U�;;es�2��Q�QrT���r�R�\\�Џo�R���{K�L��n�ai�@��~w#���^fp
 ҉��j`R� �]lY��K[��Q`���[�!ܷM�pk'��E�t�M��U2��$��}��Q"���Q��t��v�W��C��$� ���VY���2i7EC�wܥG$�:��x�We{�	2��W$Fl� #F&�������Ag�m֒�>=�q}�*{�vF_WrÀT�h��XϫJ'�ώ�Mv�f3^�[�y��eos��57ep,R:߂���c��'8p\x���P��igZ��g���j��yh�$*W]���[�E��5��,/QMe�
���ؼ���*�/�\6|-}Η��*;=��������wi"�A�c�����vC�/��g���{$�r*'�2	�+�4QV���u���w��^N�OΗ+&�Z��m�����wy��g{>�]�d*3G0���O8�?�9��սR��/�UhT*�x:q;3���C��DOս[(N�v"�B��s�a���&���-P�X��M�C��y��evL"�vbh���#7�S�Z�ǓU}�u{�j*�сVF�q�ն^�3�U_$�ڙż
�kt%NA;��J� d�d�"RHM��ݷ%��f�9.�1o)�Ie�t��ח6heN s�qK}� ]]P��۱x�Cd�B������� =��~ Rz"7zu�Nݮ�1�D��׍CH�́nZq��9�|��ʘ۩�N�$�gW��b�(\ˍ���Pr"8;u��~�wb�g�1�P��-S�Yz.��j3����,P���M!���ҽ~y��~�[��M��Xbt�y;xZ%���CUl6����(�H#>�p��K�1"yNz���*f5J~!"Ň�;H�#�E���'P�;�>E�7w���]o�]�q�Ք:#e�g"�� ǖ��C�eT�<J]�>��ty��%yTNV\��0��$�ND�ͯ�U���i=΂���dՏt��b�t/��WC5:ȫ�;)>�9M����V)�W���&bB`�~ؾ�MG@ګϽy�msN���Qy���J�0E���'�̬�(q�'��2(A��Q��A�N��ъ�>�#Kt �f�3{��}=�������d�ߓt�3Xl�`N���g�^�`�m&�<����{�U�=Z�����yMص�3�)�ι[�m2�xn��)yw�kD2��':,gC�L9���)wo���bc�g��2ݠ��sp���Ӷ�W@��'0��l���8i�+N��
�%�6v����s8��N�:u_qv6��g>#T�#}��ӌ��xo}K#T�Wڝܘ�?"v� ��mQ�|4P/ORk����{#Y*��`�[���0�Z��EGEn��/9���r�}�Z�����na�쒯T��w��I��ﻐ'�����5�k�r��[���.:�>�`2���|��]z(��%
�.ѝ|�|�+=���q�=U�z�ey���V.x++��Q���J��7l�C&�k�
�R��}e��w��S}�D����������ec��?7����n��y	�N;��T��N���D)�����y�wT<U�tz�'L �\@���q�%�-0�Z�ͭ��kf#a!ƫ<�#�K-n[='���������z�:�����/�w'M��?XK�g�
��Z.�^�WS��<���9�o�0ʏ�W|Ub?MV!8af�yt�^^X�u6lĆ�X8��P���	:5�W�!J�<-�-�y%�]�> =ʹrT�XVm�C�����>0}[Ȫ��0.�_Xt�ޔ��k��Y��w�t�';U�)��ر��ab�B2����VWm[�[,���Ka��D�a�s$j�Rr���1Dd�f�@���MH��0:W!�Xk��fp�LW�Id<�s#T�Kp��wf�e�5ψ�+��Ы��o� �\yru 2U�?r��s.<�Φ�=Q��IG�r�oN��E�-�J��. ª��A�]��*�!�M�γ����}8R��y��`9���o�,v�{�����R'�֏j�㢊�y����y�{��P)��@�=�¯��h�cD0�ϙ+��dB歕- a}�&;ULCr܋� ��s��򋺨bzFD���B�e�F:�iRB��ndt,.j,�B����G`a��˒�韴F"dŌ�/Ƅ!~�k��Ԫ�Bdl�nX��'b��ג�[�6�27�ش!w]$vP���,���ve3½��A�8�V�U��Xok��y���dnƙՊ{Ɋ�THU�Q'_���0�:������ҵs�x��}P�MrOv�ω��L��p��!�9�'7�}��z�G���݄+o���Z�XR����f\��i�y���:M��P������Ǒ����/�*�l1~1�ἣ�	b�c�u"ls�b�K|if�,L�9�َ����c���Zȋ�t���M@���4����|�1J��w�u꘧[��9��M7Xo(W��6MHV{$���,u�G�ӳEB����T�](�҆���Y��M]sU���\����=�6}l���-@.�����%�zpE�&�F!1��
ӧ����t��n�ˍe:���75��05��Ij�_>�-t�.���+�=C����%�)��#����<���/��g|[�X���6��&9ŕ ���x�4j��iEk�>i{L|��ui��|�4g	-嚗�GEKX�7��x
�E;�t�s�o���P�N០��t��6�\o���WW.��K�mqhU-��l�FPx�v���lK����gĤ@�b$��:>��	�6uM����{k�S��꛹)D�6̮�^��� +_޿D.}����V)���$b�24�Gӭ8�&��T=(D<9Z�C�n�"��Oa��d�9_:�e�\�\mM��U��vPx�����X�2Az��Әc� �����I;AZ�ˀG�4���+�Ybc"G��+{Z�w�iL�t�G���kN%#�D����v�:(q�~A���Y�ں_����r�V�mb�z�`,���Q���iD�H֨��gY�N�p���;�2�5Q�G-�:�ڢ�*�/N������.<`k�rV�~�����G1���m���7�%��On��[8�K�l��3�? �~��ڎ��ǝ��l��{����5����X�h*w��{r�ǲfz��xY�W�Ss^�KGV[@��JU�Ю�m�m>�;�|���������qd���H��NB��,D�	^�V�8��;{ވՏV�@����9�rX�� bm(�ƣ&jW�Z�l�k�޾̀5�jZ�^�^�1�g�nt��185�~U&W����R�lcI����Ls!D�s��f��������)Ϸ�*���b����CD�ܸ���:4O%��汛�3��o�a�'c��K��w�O�Õ�I���ʀ��]
�<�ٟ>^:��)�[*u��H_Z����s���௪�|�W�[r������B�'m��� =�� ��� 6U�^����e�������v�T����m|�Ln�ZI��G����ѯib���'TP�x��k$�f�'Ie(�y1Y�c��s5){�����~��Ԧtu�� ���Rٝ��'��5������N���f�������CUo�M�����(�RAȿ%a���ׯ�m�� d�`y����cQ�J�!"��u�s\��oOև4qiŬ����^��L��8\( &�''^�{�P���X$\����6Όns	�}�"<�?Q���v��u),*���b������jMu����JTlU޾����lG6��X7	�Gg��#�ޚ���Ej�n���� �yO�Y�M��"o��]��ʻ4�����>�'E��-�B��9oU�3�r�>�c9*�s����X�f:r�g���YY����
�g�ۢ�)ז�r��Y�jU�K�w.�&��-D>CH¯�Ժ����vl��]����,�ԁ'r뷹�ԯ�mu��[Ǳ�^I�Afs��o;n�6��v�kMm[�;�_k��;!`���ù�T����t�tFP�/qb��Ԭ;X�\銶�"�=A�3��u'4k�A�Фm���N�WM�Z��|z�j��{R�ܭ��=w�Xq�b�W�K1��Щ��ٻNWP$е��*��������� S�԰9̍^�=��Xq�h���mH�tD�ǝ۹q\}X�0%�"���	ʙς�K��Kf����N�Z�^���#-R��+5moV@�@-�nN+p�\�vtb�ۦ��n��/
��N!Q��@{k8�� ���|���59;�k(�J��8��r΁]�<��\�; �0�9a�Li�z_Wt��k��wn71t4յǹԭ�޺IaL�Q\^�z�oD�ˇ����4i)�vvI�V�Yӧ3:��$��=L����;{��Z�hH�nU��6��cv뻲K�5'3��Ě2wO���y���%���ol��m@��2wv��j�4ќ;�Z�h�n�h�-5vl�٧(g&�'���ޭOoR�û��a
�Z@f�g�R��Z+�[&ŧ"�yg5���t,�Q4+z��4������z�x�Z@ۺϓ9:�q��{Z m�fC��i]�,�2�3k��{��GCw@��B�`\�Ǌ�G��];�.t4{#;\T���g.v-"��f�`(��q��7x�.�:
Z ����h��%�5�Τ3o��������YG�[��!v�H#S���u��J������fl�-Ēf���������2I�]e-Ȟą�ل]�2��֋/��!϶^�4��rW>�ᔃ¯�-}5�K�쒹�b����Vub������>�"Y�9}C4�lQ�e.�8�;P�7P[�7�m�b�<��@GBk�Led5���Ez�h��Z�wT�?�p�0OJ�(�i�~�M# �ު�l�ۘ�~��z�홝6r�+��W�У/c1eLI�1%2|u�ZEs��n��隥���f�뫙�/�����>��nb-%���C#]�W �0�=;K��aX�L2R����Օw�V�Q�B�՚ꀮ�ʕ�(��q�Ł��O����*gWS�41���n��]�ob��i��9\ِ�b�-�]�J�f�Ym��-��n����G�I_���EG9����]h0m��e3�[��:�$��%���yE/�؇6u�l�uaS��}7/�$\��WwWE\�4
'wb��	i$�s�H��h�т$�22	F�)^;)(6�;y�e�4����D��tD s�p�Ɛ�S")���(��f��WL@�a�Fi�e$DJH� 32&��� i`d�P�Z2f�ACBfFc2C1"6Y��H�$P4�.K3$dA�i�&E;�)4�RfM�����#%).\d��D�*F�"��Ȃ&e$�L���f"L�[��;�H��&�ԓ9v� Ɇ���L�J@�I��M�Nv����vX�,BH��2A�1�[@��%F4�D��`f��JM ���w6�q��H��*���S�sE]r�&�m���M�c��;�X�.���fHu�.P'G����	��Km�算�G���� ⮝ݚ1�������_P1�`�^�^��zZ�_�k�+��^-��W������\�����^u��m�W.W�:���}�|�uzZ|���������6�_/w�Ͼ���o��_>�|�l�9�{3�yA����h��"@�Dt������/=�>��k��wv����_W�ѽ��^���mϋ�.s�������j�W��z�����k�okſ7����k��[������������(p�]r�^ɳöp����,��m!��x���������ͻ��V����_����y�����W.o_>�_�Ͻk��~^�y��վ�=-?'op���^7���^��^�;��/j��{������܅�;�ʅ)z���S>���. ����j���7�����ּ^փ_�?��Kx�j�|�篝o��x���Ͻ���k����������\���y��j幽o�{W������^����ү���|��7E�ˆ��[s�,�F������~/_ݷ���u�������o���zo��5��~z߫�h����}�~5�ޗ�G������W��o~�����������+�W�Ϳ��_~y��v�*����+̨��ڰ�#�U�2) �Dsn�����+�����_���7�nU�^�.�6�x߭�z[������W����o���o�=yw����~�{�����Z7���6�ݷ<\�����z}r�������~^��$��a�H��#�E�~���_���W����yoM�Ƽ_�{���zZ�׾��~�ŧο/}zX���x�wu|\߭��ߪ��{{ z>��ܺ�������H��D2F{�XNe�ʡ��E��[��zU�����{m�o_�y�~����^ƣ|����^��n��}����zo�W��y��h�U��=�u�k����~+ſU�~������^/�~^���#�#�".�i�7���v��w>V�폾� t x-�>���0>0|~0ջ�6�/_�߾����_˥����ޛ��5�����^�ݷ��m��^-�ޞ-�����oſ7/�zZ7�{����G�c�
��eяM���I;��Nן��W���~v�?ݱ�����|�or����<ޛ��m�|�ޖ��m�����Z~���o�|���6��������m��6����_������sn� b�>1�l1�N�J�ތ�ݗr�=��j����)vȃ�|�q�[C6��	�u�t�87���wJT���ݎ'�,��JР�z��l�gb��Yr�,,�������H�e�Gn�>�]WD�=�<�TBoVM�-�^ēٜ��3��p���T(;��ɢ��;~ј��S�h�3A!�tY�����zZ?=�����������Ư�[����ӻW�?�z�_Z�}[������W�������o|���h����|�s���x����=|����%�����Hw_�ayV���}��#��r~�,}|[�ݼU+�6��ߛׯ5-�-�{��M����|U����r���ߍa�����nGG�|��B�T׍��/6�����a�����0>�쁐��\�w�[��x��{�ޕ�5�z����o|\�7��-���P�:Ǐ��[hd}��� 
��}�����3����D|w^-���G��:R�;!ǇDh��|����:z`鏣�ſ^=���+�ţ}~��y_����o��*"�����zZ�cr��||[ڮ\�{��[�|��x���z^���G�}C�@��Ωj�EW�Up�^S��SQu�|�x}�GC���,G6�x���Ͼ^�x��m�y����Z���d
�~ �>>Q�����@P+��׍ͻ�n|\�wj5��7�|d
���G�?l(���|&@��[U꤫=_��X�Z�x�?���_P!V>�+7<����W�>}�oo�|W��~��z��友�o?~��W�{o���_�~����K��~}��^�:�-�{�ץ鷏>u�/M��+�|G��|@Vu���"�f��ZU�؟Z�ct�������y��@���~��v�꿛�{������Ѿ!A�_\}��8�R�}�������_�o��x��~�潪�.k���|���z>�`P�@P>Q1�>K��dr��g�;n����^�� L��">���nU�����6�noM��o���o��P����z&�;yRG����/���/�{��ƾ�Ƽo��~�}ye �@�2~P>g���e�V�/7&��$�&�����"��?F�|�v�5��/����v����W�O>y�z�7�|^/��7��y�*����������Z-�\���|�����ֹ����'#���.��c���^hL���(}��?|E����F/\�{ZwW��<���/Mx�����^���5�޼��~��߮������j��%��=c�zE@�1�G������( 8>گ\^{�S��-��S�lY�zc�U�C��p֏ZY2>v�EV��<EnZ��2R\`ճ��\>�|�(��}����/N�<k��6�R��&����{�י��9���pePm��{)MԷX���3k���w\!Ѻ��^�(�fB�Y�ĳz��ﾮ&> }���@1��%�>�s{m��ޟ��߾j���p�������^����Kx�^+��}�~u�o��o�������o���o��ޏ����������  �#$����U�K�GYyy/�Yt0=��\��W��~��׭r��m⯟>�zW-����/߾��^��n����}���~��}��z�znoƿw��/j�w���x�ޏ�& 0. �#�c�M�ǫ��:�]�k�;*�=��F��DtY�����^7�x�?�W�b+��ޯ��{o�_޽om�����w����s~��_�߾[����~~��^��o��W�}��ο[x7��~}�����m�x��?��~���o���� 
����E����?{^~��~{��o]�?��~_��wm���_˖��w��������ŧu�z���_��}k��׿^o��F�_��}���_志�O_߿��:���z������b-���o�d�L|�}��?:�c�}\׊�.om~n��]�ͼU�s����޽�5����.m���[����{m�����|��ѹ�7W�.1#����}1���p�}�9v�H�{��E%���G��#�c��~����+�_�Ţ��|����ޚ�^5��r����b��[�^z����m�W���x׋��������r�|����oJ�-���~�����~��#�P��%W3��^U4����6�no��}����m��}�cQo��x����~���Z������~�k���m񹿚�x׍��W��h6"򻯫�^->v����7�żU�μm���3��Z�|z�6�}>�xt.7�_��A}�~�����o�x���y^���o�5�}�y{U�����������گ����������?��z~��y�,2��|I��@�@t}�$O� �� >}hژ�i��Jפt E��ux��{�׭_���k�����տ��a�i5�0:�c�6��񱾘�����wV����"��-�6P�U��+�����Æ"��hB���;
ֲ�n�"��Y=�ۑ���'+�UL��5��)?yp�x�Z(N�l^�]\9�v:ܱ�J��w�T�\�9���sV
�J�έ�*IH���-�$�M�� ^�!dTk1�;���R��t�;ʼr�0��D��^&92�=W��MDG:u]ޥм D�՗�K�*ʷܤ�˧��!�Y������h\R�c� ��wʾI�y�VY�#̜����J%�j��l��_Ћ�O��ejD{��F���(vWV��u��dӱT���Sͮ�⹤���Z��`/����\��3J'�a����x��ۮ��\�ZK��ZQNBS�� �뫓ᡂ5�`a~eFP,Y�C����P�-Y��NG�pfN�T�k��]����1�1�u_f�V;�!ɯ����m(�s2���D���F��0�ri���]N�^�l	Ցt�'/�Z����H�bm��\��t�:�:��֋Rl�*�������x]�5��j�Jj���+&�Z�t��E�%��汛�)��q9s�]�� ���V����C3��۱]k�W���q;3�|�vxSzh"-�z�F0e��V.�ZD^����5�Ǣ}^�ظ�6Od���U�����18�y�"�0Z���XV^�S���Db���M�p:���22�m|�;)�������A���4�q�D�L.�W�H�Z�6(f���BZ���P��.��c�:�5X��X� eL斂sS�d^o:tw:c�͠����EyW��Y�ة�������F�Y��������wp�h�"������ܬ�6�j�k_I��������b��3��ZU�9�UrX6P�`:�¸9���L�jX��V^��j��GA'I��u�vuwz&��W��+J��4�_ICQ�J3����RYxc!��>5�#��yU�w�:#3Wy=���F�t��սc"��t�*�*�M*���y�ҵ�¯��?{e]m��QN�R�:��cS<n&�eEI������*� �-��t
S|�!>�ݳ�\g���[�O�=3*�z:;�����%%Q8\@�s�'0Y@@k>	)Pvc��L,��m��;l)��juuF��7�꺡3yp�M��XddY(6�DP[��dLt/���҉�25���6�X3�:���/�q�;�~��BNa����_��hǀ���7+W�(غ�-���a��=sy�%�*N�����?8մBE2d�&�~f�
����j�9يu%���X�S$9�m�;�;���D���?�e�a@f���攑���%�9C](˦&p�|�쾝�W.���R@����A�́U�
��.�+��e8^���X�j Ɖ�N�b��i�;�i��W����>��"GQ��2p�	:�*�/�.�gf���\�g-;�����=n����X�ʡ���I�T��e���$��T������1J+.�p�ja����DwqB����/��2�Ai 5��{0��]l7}���}G����_�C���8F��A��&ϵ�R�c\�8,����:HzpGE������C��I/{��_(}�r��x����o�b�f�d�>}��U=��+�:�ۇ�'Y:�sI�^9���/S�"�!�]�N.ZC�(�8�ٰ�-�Z�lP-d�Uݏ��T����v�דĢ�&���8�U�}��������=��4�8�.�̠���IرW'Hf��ά�J�O:/ssO�{kי-`e4�#aY5g���%������}�Z�*�U�zd�䛽V��g v]>�� �+F�"�D�药o+��������:Cއ0�Ϧ5�ЛGv1*��Qɍ�*��g�i%a�AzP�aN�j-/`�Qb�T;��FN�iT)���!�rt��`�\��w��Q�j2 J@�r����# ~X�s�|���И�6QX%�<�8��Ә�1�h<�#��M'U.n $}��J�J��DF��}�j/oN'�Hl�ov��y���τ$}r��۹�hD��2I�s�����J�sց��0���2u��Յr
�t&��jR����̠��E�5����U�/�	��]�B^�&"�[�{dr���mo,��+)>�V󶤾�Ǹu'�rTRvַOe:�;;y�霧^%ݓ���Lav˹��NE.+�����~|=�n{�ݛ�#�O���;�zzh{�Im�}󙍇�m��!��C��TN�j�g;^ɕ��z��QI�1��*����lӳ̡���P=�I{�l9�-�M"(��oY�7��(7�,�/�u��C�H�`�4{A.^��p�|����%&y\��f���b^���J�_\/��B멓�۟D埐�7f��*2���L��|���-M�5P([j�.9ɠ�X���'P�P��1����i�}�{�%���*�F���]el_�Ló�� 8�-��uڨ�v���֢��%�v�D5
z��Ca�\�=	��i��&��I��;+x�\�ƛI��s�w�qVFG �qy�z<6�&�R�`c��ֶ�}�>�y>���Z��6u�؏ah�uA��6��m
L3:ct�\
��A�s�a���!�l��΀���\�O2Q[՚��kP���8�L{���4���"�p����QZ�Ji{J�vU�4o��ϥySU#�EoF��$/9WD��hd��7��Zζu��t�yݷ�j���J� .�'����jc�נ�&o��%��ښj���G�R̮,9�B���̫��t
u)��۵����{�HݸX���I�ѮoO���������nG<\plɕ�z">���j������G��}�� �����z� ,�r�Nџ��zk��gpU����nt�x;A]q��,_9t^ȶ#�����n]�Ά�zr o'T��[U�yxu����_;���x<5Ft�}�\I(m��1�|�v�b�:UǬ39>���9�D�[�c�.�a^� 1k���㢠�ªo�C���M��d��nFB��5�{��h�8·8�^��l�ǫ�k��l�@ՓCԦ�����?*������e����z�����f�P
��|K����iTQF\�$��@���MQXbj=(:�n܄$lN{�	�m�b��8~{��.�f\F������q�-�$�4v�B{V#A��^�b6�Em�u+��oR�=C��z�&����t0E7,/���.<`k�rV��_�&F ���:��H�+�Q�;F�Ǆ��C�ZVo��t�,���m(��d�>�+D�ﻂ�^�����dk��?k�WAOa8k�:�Z�����3x�q=�^����Kb�OV��1CX�2���<5���~��S����%��x`��+�3�sfı�א�ޠu=_Iy����n,j�m�Q���U�{���J�H��[̋.���\�Ckۗ�!*��@�\��  �Gf��l�<u%s��>����cp͛�,?��@��k���z5~??�+&�ָ	���Ї�UV�'X�h�6��V���:�:���_v�+�1xU�V+��e	�6TE)`��@M�yKbj^��m7OY�fn�C������t��y����l��E}�����ZW=�iu��2�M�[�_��P N7Z��C��])y������gdCn-$�h�Fu|�ob~��x�|���6+0GqW2��Tx�9��0Z�3ee�[�4Q�,9P��"_�Hd|zY�Wq�1rH��(j7	Fk����,�!��j�*|�$}?38�r��uo���&}��B�pCV����"kY���� {�����i�s{o����h<٨�Y̆����ڭ�.J* �Z� ���jt8VT�<�uY^�h��Nԅ5��.g����n�A�:nR��9��B"U@�1* i�e]����]�rq�}c�5a���t��ֲ,22,�k")�v	�1д���Hy�%h��bK�{�Z��v�+9-^���ik΃��.�E
~��Rތ�s�/u_X9����|/�:���v��htb+}�u���W��J��GV^uJ.i�ףY��5�����Y�qSt�Kx�Yx5@�d�˫9nwvsS�1�Y�\�p��(7���h?� ��7�=m�J��+=����C�w �M��]����\G4���ȯ��GePb�Y���|�����,�JsNQ��s5����[Dj)�E5 b3N���(�\�#
�C��Ԯ�Xmd�Q�E1�K���/y�vz�뎻��"1y�Ț���8����e�J��W�J���ط�1�� Ɖ!刑q��j��xQ�:�{}jM�U3�&v�rzq�wo\)j27">r6StuiQ�� N?����vk�5^��,v�xD��_Y�P̶�׏�ZYK��O\�}*�x��(��Z�;��e��ÊĲ��_�bg0{��w#��Lh ޭ�=*�<�}�h��=�|ּ~�ǁ�Y���U�O����Ɩm��%�� v�g�j��Y���tc��n��}'F�z�I�e���!�he{NpM��2��{dO����q��<� w�e�A�l��t�v������n�9��omϪ�V
<V��\5��p'V���׷��/,|�Hy�D�]��sk6�	�]m�Tȗ:�eۿ�0��$$idk��Ԭ�ȭ>�h��/��]S��ގ�},��a�.[%,i���e����̄�`����V��L\E�ҋy��]ʱ\Z�T4��*vV%j�{z�	N^��7��𸦺��,b!�1e�Q"�ȸ��r��=I7ҷF��S�㇙b�)Z������PX�ՄF���S���>�J��*�	U�d�9f�:�8m+����3����g�rrX9�D�S�p�kCN޵X��݋z	�� �V@/k+qA�k�h��t�Ե.��Wb\s�m��T��B��(t��(�����"�p�RYOn�a���ipM��W:��R�CnM�9&��fQ���Ç��4p��)+�Í_���v�Ѩm6��Sm��-�Yq�S�gv]�]]tɒ�SDF�v7M��7�Q��Ш��tIR�D�dn�jn�mڇ�����j�W��L3:��Rp�����m�1˷ޱ�@�&�[�/�V�J�/���$����`�هS�eS���N�p���Fp�ւE�#��[2�7[W����bn�{ne�������xS+�ng�;�\n��I�zڷ��5ΆJ�ѩ����1��[ؒ���o��ᖦf}�vk�O3vE���0"�����hf�z-�Ⱦ�m��DnD�|{�*�J_w;�j�/7��Y��)r`]�|9QT��vgvRH�>Ƿ+0����{q`��u*۫Wu]j�y K8�����{3�5�*K�#����.�T��.��-1:��B�妥'U�{2��������,eX|nwK����3���ћ%��ص���K��G�8ne�V+{�����Y\�젹�Y�h� U�{��{i@kV�\��nV��h}�
z��#�ʼ���l�����nU�b��w[����)>���.*6�}t:��5����F�]��c�Dr�j��TZ�O�٦���鸁����y��u�`�5�+�����R]��`�ZF�%6����F����0i:x�[�Ch�e;3;<�1�e� �(6����n����rïeu�u`�ִ�Wu;w��M+�������W�z�b�R�#��Jtvά#��N��[L<�S��s�z��r��=�Z��x�BC4�Z��M
�>�.���w%�v��L�}���У�*d-�;C�X��ﱷ[ⱙ�Ȝ�2Մ�
ݖ@uo+��ԲX����#wO�껡͇��P�[Olu}�7UE��b���oZ�i���u �����Ԣ�b�b�8����u�2���A�k)�NvZ� *z�Mۘu��mw��{�2�ؤ�����7�$6p5�C�C�'hf���F�ޓ �^iA�7��(�1�j�����Ǜ��z^�P��rڛ��d0��:��fU��[/7������tp@1^��|�.���j*X��f!0u�quf��jd��5#��Q�  � �d�!1K��iQ�L�F�IF��F2�"��P$"�#ZD˜� `4N]˲�9���9L��sv$d��#ww.ĢL��wp�B&E!��r��B�2h�I&	���H��D�J%,�%(M�i��H&��̔��F�I�C!Hb2�IR(��	L����$���wv��"@�F�1I����W)$�2����"!Hf�Ww(��[�4� � �̘�'.�M��n��2�T%F
P�$̂��aD%ˤ�FDl\��\9_�uU�NJõ%4:�qգ���_N殳�=�ҥ��S�w�Ubj5��WP�ι�*,Tԇ�Ze�W�
��NUћZ��_}��}�;ݎ�ӊ�(q���w�V#���B��J�8���q�]`	s��'yu��x��9��L:1�^��.�`k�b�IG��;w��<G��d`� �(�\�R�ݪ�.���Y�4z��n]	��Cc�������0E���Q	�K�D C��П|r�پ#���=:f*��ʃ����"ɱ�M��w#o��I�ʑ<%�rp���o�4ݻ����73 }�tW�G�|.���T/�u�m��s1�d�%hu���9FF
Z�UO^��lY�V��by alɇ�%Af�e����͢ZfLj�E��T�^�Z��g:�mw&`��=\]]?�����~FrDV��j.�V%R��.�r/]|�F�+���OFH�Ҷ�ܦ��0��f6er�!��g�1�B������B��^t�s���똽{�:�L�m\�\cub/��fCܶfk�{$�BC�_�9,5�^��=��}r�gk����E;�{��҅]et\vWsQ�i8����y������l�S�gn�,�X�S��8�l�Ř+I��*�s�1�lf73މ��WGU:���a�xNY�]&�9�CQsiV�Vk�[��x̔�)B3E����u�X�B� �0bk6W}�em��7n1�ǂ]Vxfosҧ^��w�u�=r6{m�)3�����>Z���&���,�g������' O(u��[�"ėƛI��Ǳ��X�1xݏζ:��^]jZ6o�p���ZQ�������
�����ֲ �M��J��}���&q�tD�a
O�v��^Հ邠��_�:�V�
�\��Zcۃ� ��׿o��|�7��Z�=����;`��m� D`��`��PS/M �bsw�e]�w��f-[��rl�C����yԫ��_�}���W�B�E$��za\���6b%��M����y2ne3q�l
3���`=��ǒc�跫�n]��4� 8��ws����O�p�=-��(}0,6j(�-�K��(o��%0�O�wS|�r���û���|G[mq�>Wi9�G��E���{id���n�W�F��(@�5�r�n�?B��:r2�9z#x���\����lp�Qz&۪�X����*��� ���|���<6���N�BN��,�WVW�;�d�iE�=�����6�*�M9:I	l	B�py�a��p�����^צ�S�L�V�)i��>|��ʆ��';�/�X�+�XėEoU��KKh	\�p�:�:�&�L5�}�5gX-Zn���g�OXŁ�VqO����X��s��s½�r��j��2��н��)4���}��܆���v���H�,�ә?���}��꛾t�(��l��[? �ZK�̸�v�q�8�t�h�d����A	�S �Ҍ��,��o��D�z�ՊW�s����eY��C�����,Y#ZOP�����@Ɉ�����Ȉҍ�4��D([���>0J��#(p�w6/��k��9���9[�H�p��c%_c\�\��	�0�+.���!�|��lcI��-l\L���f���2�h��G��H�b�!�f�#<~<a3mp
�����}�]rC.N���8�ޣ<��eac��;�5�a���PnDE���^���Vk�x�� �.���D=[������s}��Xi�_n�׋b��ڞ7P�=��ĢpV���*��a�v&ߚʭr�֫@?x������bs�������e��:Iӱ%"�nV��hk4&��S�~"<��C���ze��RG�����1q-S蕗��JrMh�鮦Uh��DFz�O$;uX p<��L�RP�l!(�G����IaY�u-ot5���X\���i�#2�brc�a��*�7����7oN[饷[�3N�^���IEͽ�x�8V��53+�W}��.\/��`�u����2	 ���XY��8�D��u��3Ӎ�۵���v��x�W���x�PTX��R�UҬj��������ǻT[�᷇c���H#�8����AL�f��_qqp���<�.pM����^����4�x~�7�pa�|gQy�V�B� �8�ڝ�M���R�irھ�٦1�4�,��gc9�a;�鉕?z�,�ȈT@�0L��~�2��{�ӽ\|�D-U:1� `^�1���WE�6���\Q8k"+��D�#���ۏ��F�q�G/���h�hp7C�F1�ǻi�M��_��hǀN���^s0�����bc7x�FR�����ǡ���80����{d�:�E�j#]�VD �м��ƼV\m,TS�c&i}1��X�b��"�~���Ö���r���T�V��$<�Y����֑����8%�7��F2w3�Ca�5���|X�^��<kp�V����o��l���o�peAڠ�Z�1L��Bl�n�	�_k��Jj���X3�,�zٹ�ZD��ť*.� ��NA����7��P����j���kd�ِ�c���o�ĥ��P<U5n��<&�ݏ8��&k�������v����A��w�s�g
ݔ��aV����E��wz÷^ۓ[�]���yj��"����Po��|�*�F���r)Y]��2%PT����;����$�����4��\���l|>�� ���z�q9C��N�;s oV�L�`�ǖϡ��q��|��I;�$�cDJx���2�^s�k*OV�AjXh"�B���@��Z��ʩ�az���w?]�.r�8�ҭ�)�q����`�[@u�õ2�E�����n:D_�x�Z4ܶzn���s�L�֋nۈ�����Ƚ/�p��)� �+�]�pik�^�W91]>����OY��ѥ1�c~��,*ȴ�8SNRj��*���0�}�'��`
�i�U���}�(.�^n�����t6�;bC�(x\BbZ1p�J8�l�N�8�9EF�3`�@J7��X�����޾�3��4�W��Tܥq��St��r���y�O���7�U?)�Y�oح����ϪYZUh�Zj#�v���t�d؄�s��m�S_:UD�Lm<�|�1���QM��ԟl�\��!ab��^���Gv��ndlͲy����۝۶�wuqPZ�{�k�X�[�jD{`�\��8m�v{���:|{KF���������?f@8��fݎ�0��XÈ�a���f��2ahe��[\E%>��o�LR�ڔ���K��\�Q�X`ˮ\���t[K)fQU��9��gR�q��w��9�VSB�u�NW]�1���P���jС��ȓOR��O�zkPڋ�%ܫ���&l�swNaF^�ǉ���a}�E���ӓC�LPq�����eQ�Hj��[�}/(9g��A���Ȇ�S-� M������������K�������"ks[�����֟|�֯jΙq[��_5�8�ss�ʀ��j`/��'P�P�؝t����fc	k�W�-�[�`\
������+�����Dm'���y�	���HJ���}#3r�ᜃ:�^'�]V6;og��40�i<��;+x�\�ƃi8o�$�Ɨ�{��Y�Q�������}��ˤ�t1}��l.#ط ��������qx6�+mpi���T
��'y���DX��2��3�	fDz%!�l��M�#ٮ��_v>},�����N�g�XN[;i�������ʝ6(�#G�H;(I/�(&6M4&�t�\�i�/�)�S#��W���z��:A�[���5��_/�@p߸@џWm��a��E�F+��]���\�l#.�3Ѽn��@__rvl=�����1�h[�Ѷ�s�O��'��4SqK��1z�n�p(����� �i��\�P\�$3DK�dŔ���xlJ�H�a`�u�XSQ��̏��eF�`�������A�����T����{,��^�pĈ�%��[�a�EuBN������xc��P�h�ǡU�ñe�5�"��R�\h]GFr�>��> *�o�A�xd���F�@��m���_u�Z��;�xv��<��~�D-��v./�-Xx��n�{
�Em������t��
��dV���i���7z:�kZxJ��H�c?�u�
�ѡ�%�*����;�LO�*��<7Dc�5�0E�~f+m�>�u��հ�,1l�ۯ�)��zS����##I�rPG��}u���t���mٌC\'�!��u���ZK`�1�"<�sN>]4�44�/M�Ji�Ũ��'|�����[Z=Z*Zŕ�I�}s�6J�������������Bإ1N�%%P��fM����'2|��o�l�����;C�6��u���}����� bm(��
t`�H��͂dz"Y�T`Tbѳ�k�+�k���O���Ƥ��iw�_�cS��R�fv��F�"q���q4hc�$Z�^�Z�����K��r�p
�뀯y����R6����X�xM��=�������N�X*���(�����L�W1/�Lp��"�K�C+3�2z���"�m�ޗ(�ߖ����������@�%��ʵ�����պ!g^_c�G�����N���jn�o�&�ꮨ�V����8�8����Ԯ͇CVz�2�oi�4�&�Wr��r��ͽ=,���]!Ů��_UUUP\�Y|ӗU7q���b��|�E���/���@g��5���B���� ������~�Mwbi�S��| �^(?n�����b�.�`�D5��<YhmŤ�4y$E%Enٓ;='\(�>+_Α����^��]��g0Y�\�t9�R�8�ֶ8_+Ϯ�eVWgP;���G��HX$�6��D�#�o���5N�CRYx}0B�U�=��^�z�{~9�^��!��p �8��@��A`��T��o��}���E��R�73�2��k[�T���ۑ�Y������.K*5�\''^��5*�Ή�j�0�������͛��;ھl�;6�I����	t��������ǹ������YxN�W�^u�]��!}@Å���/�6��a��d��Y��"c�i�����^j�F�0�^�F�E���[���(6��vYWq��(�N�XO����{��Pn��
�E��=��R����9���}���<�G{�`o�����#n�6h��ō�,�f�Y{�1>��+�{9%�;Uذ���L������bg��H6-�IjX��m='Յ��&mlSFD�����Bu�PE%Ye�ۻ¸CE*�2.�R���8��З�Q����V��ج���^T��.�Uk]�~^�ꯪ���{v=���X����~�%mX����>�ĥ�l�y�r�au�.W]wzFiK�h��8����ey���r��w�+���h�a��U�tk�l7��j|�Z���/��.*֫���vz�ٽ�;�1�aS���|����yJ́�`�B.~�>�vGR������\�;�aջ��&6
N6�t�������O\޹P����9�ҋ��l��2�[�e�����3cV���b���ڔ���Ek�G�X�u٣��6�ך�Q�!	��q��o9�u��z�9V:u<߯�͞7^�_t����f�sD�֚��
��D��w0����\W%�P�=/j<TM�ɰ�E�k��8�9�Ӣ���^KkC�ϛX]�h%���$U���{;��-�qӦυ�\��#���Z�׮��i��W��R������ ���wDh/����z/oD+��A�'�e[��N��>
�_j�����sΞ�s;�)��oe�S�{(�㎼�3����%b	�^+���Q;�S���\��k�����Z�4:M#|Y��[7L�R[C�X�:�k������evU�8��HѮ�Ù�|�t���Z:˛A�0�^4k�#Z�+�Wc�܏�u�)d.��_����菡ZkRA�ڬ������u�ϊ[�ƞ���^���k�J�%�+ucOV����57�w��}��,�x'���Gf}{���W�%�g<g��Nd��������l���x���+�{S�����G.�}A���-֊��p��cu�
E���z'])���n�+ntY�.�)fa�eN/�wv�rNW��8^n8tb�Ea����� �{��������p�������X�����>E}\����3k�/���p�����7}����G7u���V7��]*��u��/�eSL���Ŕ�۹��{)brw�.���Œ����k9Z�x�gP]��1з,�}��{3����d��o���72�X�.��D]��jm|'\]�<�;;;��$5oD�uv���5�B���m����7qw�ԁ��Sk�<�����~ǋSH�mCLY����t6��: ��N�T)���[AM%���\��e��@.W�IK_{�Cî��e;�r�D:��l wq��v��K�ڵ|E0a8&o����i ��ڎ�<i�r���Z�3�Xԙ���_h|�jO����%�YE(���|u�Lk|I]e��}DT7V-�}L�S�Я<�6�w����R�n�1sw��D����C*5�7r<[�:"�6�:�Q��`W�9H��a���5��Wv����|�j���vh��y��Q��vs�n�\r��D6��P�L��,���Ύ*l��A���+����s�L�^�ͤ�Ps�圧,��Ń��^����,k��"�yfT����}��dE�$��*����*w�+�zj�v�oiK}��"�V7/X���-�m��#n�^�E�恖����\�����5�u`��A���\CT�Q�|sl	N��R�W9�w5y�ϚW,a�e���ɳy#��$le�*X��`V��a1m3%خ�%��\����հ�u�IU�j�9Y�r�s&�������Xj��֐��N�c�.;�V��C�(�wڴ:,���3{E�]�p�Q*�"aD�V �ճ�%5U�n����m��+5�ut&)˨:�_�"}����es�z�*q����_�k�K�2�_��w���Ĥk��w��o]����ء��n�����R���t��j�=�!�c2���SfM��qD��Y�ZF晙�gg-L�ep�\���W��bh��Y��宭Z%�w:>�����w�K�wԥNv�[.�g�Vۄs9Y= �/K	5ҝ�����7��Uܵ^�ݯS��NKj�*4]1�f��v�zu_$wa�N���V_}�n���>����2��}�V���yX��A0��|O2�cc�D��b��A��T+�B�8tE������tF�qnQ������U��֦CI�^.a�&�۵B�N��c�7���7�����(i�ns�mr�#�Ҳ�j\�j}\�;��V���s{�(u�ќ�	[�CA
�д��E��	�Y+�v�06�.A�.wY��j�:�a�yw�h��hG)�<��oK�We�sR��O^]K;Җu9Le�ށ�L������4k*�3�{+���!���%Ȗz�jU�Ү��'���S�; �,W)�)CUl�8K�wq���b�r��V��ի����t4d�0�ՅǑ�Nڮa7����.�]53��0{0����;�A��DB��h���4������� ޖ�(��T�:���
3���	7t:�>��Ήr6<��t5𱂓� >yI��B�sb��r�g5+��wdY\�a��ka
=x��6��wXݪ�`T��U��� 89X�^`�K�����:֋Y�+�X�ݒ%Һj��:�Rxs���8^�uҸG�K�|���^
�F����	���&Y(��#I��݌��FLa)1�h���"(eAb(ؔ�!F��P�2e����R��.r��&(�2H���"BB�#bܹ�#6wsdB��#E!�Q���"�!$Q$�T0�H��)6H�Q��R��,�H�`�]ܢ��,D�	�&�fiw[�1�0�4lEF,�5��&H�D@���gw,@JQ��gu�21���$I�`HL؀�Y'w`Fd��)4;��$$�DR[�(��(���FB4lcb6(��9ʌ_�{�������`��\��^�Yĝ�<��J�8�i�	X��5�w��b��04^�W�:�}7L��]���9�s�U�W�|-oR]�|䘹��>�uy_7���b7&�5o���Y��l�^k܇�;ِڪ��xtOկy���z^��z�6��ց�lJS5I�b�w���Z�9�ܾ^��U|9�[���yG�z�a_mt����I��Nre�E�k�G�[R^�.�(_s��>��v!O{!�plE�!F	2�ֻ�M���]�q�rr�Djy��AK}%��c�dsm��z�o�Y��n��4�-K�B2�Q03^��Y7�m ��Py��c�SJ=3�7��=��Ϝ˔�Go��t�y��~F�P��!�5p�<�r�i��Cg	���a�j��FD9�4T�ZB��F�ϧe�b%��!d�]fou�QyR�����Ook:{�c��?'lW�m�}�=m�-���2��^Uj6�_ӛr�����or*�\c/=WWCːeQ����퇘��/Ȏ���ы���_A��:��p��1��q����WC���n��K������h�1�\Úƍ��䡶�������7V��W��&����$�;c��IF���U��9�q́�ϩ�k�1�0��#gj�b�6�P��~������daz�o޻@����M����^ƹeF��ֲ��{�M����MEWeD^Ki�ͬ3��SlYK�荑�}|]��j{��L�2�R,w�pM�9�j�^1�x�|�J�1��E���y������i���x,a���zι���7�w��m[�����̠]H{�MM�!����ܛˊ9{����;�� T�z'OWs�RO)<��kMſ=�����ys3Ґ���u,�s��������*&7V�>vڸ����X��â�m�I׾��Z9V�JW%mJ�^l(߯PNnonZzL����a]{ٙ9a�1��.����Q�v�Gu���O�|���a����RNiһ뎞1q�y�ey��g�Z�9n�*�;��/�LeKS��;�����'(Un1�o�����O�:o��ĎA	}��hmO���2!��e>�ԫ n��i%۶��j�x���Ԗ���3.��vn�XyWw'�c� �t��T�my�,�涮���^�>�X�&���v��K�:M�v���o�j��'ԑ֯h�Տ�U�k93��YhE�LI�U��X(���Y>���6�K��.Z0��O�׻_q���\o��8�K�s���� b�#�5��Ow^���iɆ���s��+f�=c!��Qm�|T��nm��Ŭu��sBg�#w��N��s�F���{�T%��6�;��0���Ssx�z�+6��zɛ���X^�z�b��ʗj唟�mT�~�޼z��,����o�ME���Č�B{���	���X3��q_)������R����켭ɏu�(sb1k�Ob��N؅آ�%y�f�r�_�1-y:dLS�op�gꮯ��m_0ʦ�����W5_cb�؋�W܄��X�(+�n�����8���kS��~"g;=�~4���/5�����9���TW�cM-����FT��&���F�l+^��h<ﵺ��y����A�Y�^���,#�]l�rj�jx=B�m�
�z�t��~Y ��Z�|(��!�k��������*��2�3v�-H�͖$e�V&�X��^{uٗ:�����덩��
�P,";�rX�H�����@A�DF��;���r��L���`���ŽJ>�8'ƕ\��w�j�j��F;'��ʘʇ�ӵի:���}UT [���+�����vTn��~��a����ێ=C\H|m�u�ǚV
�j_��ۉz��m|���+Dl�^ȃ�������S�op�%6���.oe<)���׮���W�\a�U��Ƞ��?%�;�l�b�.�������{�`1���7��ў��y����0��]��X��^m4��L�����d�a*�׊��>��s?l������;���A�6�it�2K�2�˚�6�U���hѷ�k������Gfn_ y�X���&�?�"�7B��n�Md�U���a�j%c������ֽW�%x'�qd���a�'�r��e}�;P�R�r������y��]�_]�t���6Nmt�>p�2ź����!�3�pF)=�w�!(�ST��QV����η��W1���>�V1��;p����?2wg��3hN=Av{0���P�����$�o �8��:V�:�j5
̶{��j6�x�ˣ��h� ���)-�w]#5��]y��nkS��,�S�����݅�|3y��r�r�bLG�h���K��qn�%���I���'3�l�e=�]<�/��  ս�k��V�әk����t��u����f��m��(�]��x�Zǆ1��@^�����I��b������u��V�yܞ�w�b�^�p�}�7A�h��|����?G�����F�Y�����;�/��Ό�����Z��(7��E���5���w��W�7��ڷV�I��k�id:��(���]^Po5|��W&��V�}�K}{W�G�ƣsK���ӛq���ks-��/^�=z�}�n+@д��r(c��Y5������;Ft�o�쳺�[�|9�}o�З�(�W<U2Q0��W�L:�S�!��[dk���┣䝼|���eE�Y�:-oI
��ʙ�n�<��W���ߵ�F�!�Q'S���j
[�K�i�䥓^PϳY��2�"22�h�L���:�}�~1�%�k��/^=�������U�符�Hr�\)8�@k\�5i��^]�iP�=2���xZ��`{b�\��G��x�|�2(�ܥ�^z�z{�w�v���4s�����1N�	?nq��]���1ME}C��T�I��� \+خAbO1�I���]�������͔�T�l.��Þ� �A��=c~�c^I�t�
�Oz^��VnW*ǲ��|�g{���6-��ÛrgѤ-��4���G�:�X�Y�V&�W�)H;jt����-�̱��Ӌ�5�u	Ol�P0e��Ӟ/��+�7k6�=�5r�O˧)4����-첦luI�ז��n�vWN����;v���*����]_f��|�3�
���4�t���Z���růԆ�t��z/�.��[��j�G7��Ǵ�Y&.\J�|��;W�/X�,�K���V�V��JK�=�V�]�`�p�Ȭ�<&���1�s�;�<e�>~�ix�^�P�ʫS�ù}}B��X�+D�ӝѵPb/V���\"�f���9��I[�s��۹*V�G�#�;�V����%��-��,�����7�Y�߹s�7���S��Ι\�|�^7Zx�q�\6Z}�fPbh�Z�³+��c�feq��ǯ�?ao��S�[!��U&��wV���"R5�Ξ]��5@vP�cV1��+l��O��iG&d�U�[V.̼<�]a�ʈ���*��l0�>�������֐	ǜ�}�+��%l�����Q����}g���s���fz^E�^8�9���-��t�#dC�BN�/T��y7�E�f}�F������{���}	���^n�x��h
`��CJ�N�j�$�`R{蝆�M#Vۄ�����7�[�0�4;����1�,�[b��u�yV��W#�.\��a	n�{�܄�A��̗��}���V*u5�v���	�LZ����+S�q�6��1��9�0�n���}��N�sP��#�P#Kf�g�a;�+"�[zg�;(�͏7lx՝�>X���4k�1i�0�����|%���b~:`�r�p��J�.��������c�lN1BC�ghBz�*Om�O;���[P�VU�j�f湋mJ���Ϸ�ߴ]/l'X}�w��'��%⯖ܭ�"�J`����0�br{����B���w�u����5:ZR���q��a��}����"�X�Yor�
�R����3fopj��m>�����l^��O��V�z.K���ZW��}%�$�zV<}x8<��oIG�n}���X�7;UF�W�;���m�/h_0��9_��W5X�\�=�qx活�S���P���;������륝z��1�Y�wY�:��ZqDZ�gK�E;9�ޘE�v�.�	��=ѫ��k\��T;ˢ�y9}�(M��v�����A�5՗\��P�`�.m}<�������5�sm��'g�2���#�x�{϶���~�roÍ[��A��>�{?5�i}�n ��v�v��
A��{6�{Kס^�k�C��UwM�� i쌡os�y���>�4����a�x��*O,�j�>
�h
~9�S�x�0�I�=]]�#�������s��A�x�-��r����)0XM�M�מ3�}�ȨQ�+_�AKv������P�Ϥ��&�ۜk��RC��b����Nυ1U}Օo�0�|����pSJ��H�,UƌV�M��f�^�u�3��OI���'_]M)��Zɶ��nN~�2�+��|�7:�|�cE,�ޫ�B��E�(uo3I�=��I�ec���,9f�t)ד{Fn� �h�jވp�!b�Ċ5s8��fǚ���j�y���K@�ev�V<
}�������@z�WʩMB��/��:��s���L�'|x�,�e�@�XS����z�{�M�0��L'Nk⥚���ʟ��5����C}�C24���K9�Geu�k�P���b����$>�W�a��H��ҀEٝ��^>Ѱξ�|	d�$Y�����;�mc��1���X����ܱ����&������Y\������z�0)�r��ی�5՘\��}Jpk���h~}w(�UV���l��կ���~�c�κ��FZpf�Qp���e������V���-.%U���Ծ;��*��q�˼Z�H���ܼ͠���^+���hx��jv�[�^��1bTw[ʕ:u��uU!�̅���so8K���^;�ct*�,4a1yk��X����7X��{q����no�����uc��ղ�V�� �V/���l�m�]K�~T(L�5�+�Q�ׄ�{MN�����f.�8�u�u�۱=־Ӡ|�S=_�k���n����Wc��m�:��,�fFp&�/)�yNC3���/a�t�<����u��v>��Ţĕ�b�R�c;Oe�:MЋ9W�}�޺�hʿ;jN�7�7E>]|9�|���y_��x�{7*�͂�7�Q"��v��۽)�H�zS���}޻zǁ{klY�m��#�-��&����{��K�Sr��Q'S��r�P�X��K�D�һ�Hc�2y�z����qP�w������Ggt��Y�q�e��w᳅'��_3Y�m�Bv�&��:d�߻d@��kɿ�&����mS�ԓ�ׅ��Oְ��&��2�;��0��g�m�E�F��a(z�%M�'˭�v\�=�6�>�y�e6��-�P�9ӈ.j���w1�d#��>��U,1ڄb��=�+�n�}r/��ȯ���m�kh�n9[�W��uO�ŉ�]=B�M	۴'�ʾ��\��k\6�{O��o<v�����r��z#�6�Ť�l�v������W��}��&��|sV�;�|�T�����ħ�L�R�W�
��=v0L����F�|�b1��;2mf�@t�6ơ�T����u�T�1}J���e�VL*R��5t͒]nӸf$	��u�IG��e���0��(f��B�#\��F�p[�"A�K=-Q���Z��N��-o�_w��|ɫye�͊�B¶��s�ԩn�<h�ןa�yܣ�/{E(E��YR��|M.���Κ�|�<%c��]�>;GҥI�W�V>��3�aƟA�[7s��BVie٧��>�4��d�������Y��y�B#1��7�R�N�U��t�*'FS�Y�y����f��MJfekbvV������S�*�]�[�ewm��v�}�N���s2��7;���Nj��+GY߶Ё9բ��ᰁZ�E��|��Ӎ��m!%��]��\(Y��ӛz*�V�2�Yu��kj#�U�:Qt����+�}��W���;sa+���VKܻ���Y��t�c�v9���b;��V����R��G+��9[J�9�h���G���En���%]N�x�+#:�4����J�ȥ���@ďKϦ[�u|�RB��ds��\Q�
>�hỦ�n�N퓘y�/�<��{n��on'>����ְ
�h��W�s���8*��3DMk�ZJ�:պ<z��v�՚#�ykK9��R���X2�[ǚ>��[�ԝ���S�:��Cǽ�hEq���x�J����MRf��p�`�!b�Eۺ��8���N�P�ew o�ﳶS�,�G�+�����|a�jt˚��4���Y\O.��o��4��=�a�`_����=��X/)wT��B��Y�
z�GG����@�ݑK��{[�u�[ɑI��5��b�*����2�^fQ�)���<B����ۖg_=�ElSUK��
�I뻭:6IVv�����(�]z)Ё�Q;��}�2��bp��c>��E1��t��}yb�Z9-s���Y9�XEv��N�L�����3]���f���1D�P[����J��~��2
��GCxM˻"Pz�ս�-.���|��]�:�V�.����s������v� 6�^�T��eE��A�)�(�,��_���b�֒k��i�r�aƓ���y�.؂�,��|v��W���;p�F�s�O$�.�/3T4t�p�
_�;��JE��/@*�t��d��Y�KU�����tB�>���l�[Ne=�K(�ᔌ/-c��̹I�'܌i��w�[����]Yj�َ�*l�ȹ��".+E	��Kr�,��b�4Z�no00�Ӹ,HNK���uW]���V�^��+��K��_����)����;m��ڷĝ�,-���b媓Muu(��[�ii.{qV�{��PJi�%�O7�Pm��\6��ŝPW]��\����t���W��F��/�%��`ŹAд�H�u���ŉ�[\�d�?���������E�2�
���r@Hئl��L'u�,F1��,c����%�#	�l�-�s���6R�Ɗ�h��6(��(�Lۺ�
�ATD6�V�W9b4�X�a�F�k��F��b ܮ��������cE�ԄZ �*,LRmd�$!�$Ӻ�ZwW1�����P�"FةF���nkFج�( �����Vr��h���w�Gg���ܹ�k)̾��k|�!�'WHU�����z�2��:��GfB�9foU�Q`���_W�.Ov}kL����ڶ�:ܳ�-�!ήk��/E�X�润A7v���(��oϽĐ%况I���e�w;}�^m��m}n�m���jI����f�2��h�e�Y�������"��^�_�}��f��y�t��h�g)�~�>Z��>L��+j%L߳��iz���'O��;��k�͕	�N�d�u��7�H���gæU��	/P���e���	��;���	��]�{��W܇&���q��{0rz��%�QJQ3T=ֻS��J�tSYú���_d>���v&���݌�K@CуtL�S��B����Ǜ��6�Ζ���7�k�k�x��M7_a�k�ތ�Vp�+�%��mu��]Y�.��;Y��vgq��7���A�ҹ�i��Q������k����'�r���
�M+�����6��!�&Mb��oܓ��j�#k
A8�uf�"��y�0l�g9��|\Ʀ֭��ja�y#i�z�r���Ֆv�ub�s����>u��y�G-�!��s9C/��x�5|/r�c��Wj��ԉ����:ь�1q�xƻ` �a
�G=��}����O������VU�#�C��F��J�z�'7�UBZ�CoC�T�9#SЈ�Q�(Z��`�y�8�����1Gc���*���{�����C�k��0��`�y��W����B��(Oϩ��ꌩ ��Оw9̷.���;�E�b���s&�j��֥\�؋��m=��'D�\]�n����B�T��}׏wՍ�~qe#��T�����M3��C]\�b.��Ou�I�I�H���t,������t��?	���y���xCT��,<np9�1�U���Y��4�P�Ir�8�'�m.�Fzx�잣C���(�E��f%�w\�Ҽs�X��y�r	0NXssط���_�ᝒ���K�N��t�Fn�/��]f7|�l�|F� �L�$�Bz����Kx�u&�6]]�Ja؛������y���V������4���V�>���g�#�1�-v�w������z
��R��J,]W3;>��H��+���!�}5&���]�R��-(�)w�Yٝ���"_V�f�3��>�GYҮ��L:J���J��U9Q]���rc4m`��{R@��g��}�^x���z�:g�Z߰�oV�7��m<�����*Zٛ��%�vZ��s�y�w[�^��~��nN?o��4���oG�:n�K�����o=4�-S"�N���|�W��Rud�;�8q���V:Rk�Ј�	��f�st||�VN"VB�T��0��ͅ���b	���э�dy�3�7���	��4���'�َ� a�{(Oc��5��Վ�JA�j�D�!���3��;�̓���v�I�啑xuN�)ڴ����/ᷳ{���E}�� ���6$}�P�t�0��F����[�؍ڍˣyR�܁z���܊�c�l[�5�ŉ�ڃmI�7����µ�EQ:&��X���B]���s�Ү�7Z��3NY��ͳAn}Y[�xg�Ʀز�ވ�z*��p�o��ҞË�	�^ vy'����0�S�,�Y�>R�!yp��`;O�;i���pS<��-e��1�*�4rtL;!�zT38�լR�Q��l_+�M����w������d�9N��]��f�Ζ�����ٳD��L�X�����h���U��:�.��ǳ�9G�V>�-t�=��/��߲~��.�)E�����MA1N)f�s:��s��yh[�����}*���Ej5`d���%�����ih�����[=�G6���|�kγ��7P�^f������p�S�,OK<�/n8_�}�ͦ�P��h��o��Ӧ��V�)>��U��`�@I�_O����"�_V�n���j_<���~��t|�^s��i<���t_Q�4��Iz��R��w�=b/�]zE^m*��4�)DxN�����>
�ڤ�݉����AwYC8�n�Ӎ)ɭ�r�V���lb�
n-4���������1�$Fk��c2Z=b��ɦjr�iɄ�������k;-��N��2��d�ϺeU�ݡ���=|d}x7�[8~f�
��V���1M��snj
�n>�|"ч>���2��Z��g���+��~����w�'Ïj[�	�SP8�|ld�s�;9���G?�j��4s ޺Dv;���˯
�����#v�3M#k{�\���؈�w�5dj�<1-��ۚ�ji��,N�Ŕ��o�}�&���v��e��!g���3f��{.P�s��@ok(�àc=�V՞[A�?'�<��7�J����`�7�{���~��ͥ���S�F����!T���S�-�.�o�sQa'���,t��	��Н�S��}}s��C�>���b��q6�T��ޫO�m=�K�3��]�wG�+��Є&o��mw��(O �^�_c�:�.�������ih��2.��/�+���i����)9H�~Pn��vV�����F=�>�W7M�fa�T�y㠢ЙŻ�������56��F�ol u�������y�1G���$P�"����2o,�Ygr�5B3hON������,�d�<ot�7�#t}��s���(um�li�~��w2�L��_�Ω��ԯ,�\u�L��7���L^����z��8컖�j�;pI���1��ﰁ�WTQW�7o���#�Z�$ʖ�^F�Pކ#���+�����en�$�ܙ.�=_�c�D���/��S{F�f.9�+�ˉ������+��f��t&$r�w7�����t�Z��u�DV���%�RzsEԹ������y��yk�}j�ࡱsy&�W��5뇁e6�_×�j���ﲃ�Ur\��m���1w�x�`]�B��_�{��KS~��k�n�����f��1u��S���w�iFܬl�v�4�-��A�8�K�VM�\����z��[�h�}X����ͅ���Z�W�7�������F����1����j��a�t�rai�#�=��V{О^�U	k'�Ys�%Q�R�;����o#��C�lO:qPU��-�H^r����6�2w�+�Jzjզ$�j|N8��F�4��ɸ�#bF1B~��2�=B2�۱�c.J���uR��/:���N�yMst6�b��{Eүl'_��z�栟^�S��9[���"5E�5�c^e�e#���g��ަj�3��f��ݯ{m�QMj��h�!y{wޫ}7�I�#�V���G:9ٮ�g�g����5S3�� �Zb����C=�t{%`�9������<��(�v��;P�ݢ6�	��cI�2xc��I�snbɻ{>	�n��
��6����̲��W"r�}v,:Ywzݧ�t)�]j��j�%�A��@�������ig66�r�1u�掝?��>nS����V�qX����dqʴ�r�Нq��Z��=:�����e@�R�"�d��t+��i^~~���a�@��:��˪M�*��H=��疏A���)�o�]f7}�|�� �7P=r*�/wAC!9�#$nW�ͫS*+_�s|V�ܸ��ۗ�l�m6����6hzb�żVކ�vC���� b��gN�R�-ݼz�xSi��^�x|{�n�u兏�ܾ��}W� ~7DN�H�����w[}����B�Ō�kp6:��l,8�7:�\+�f᡿k�p�`4�N���~5Rݴm�H/Q�v2S��5��x�����C�r�9-�Nυ1W�YV��+�1��4^u��i�ճ;o�˸��襉Xm���ҙ+je����雜���A����q}�=�2[�J���
�֭���>aX~��:sQ���;XN�o-���r|����V1���e��d*
-#Ϸ�o������Y5n*ో���g�
�<�&��<�AϦs,�Ȩ��cޝ��F�b���V�TP͓�X�e���h��J��%��^��k :�a��ܦ��dw:��ԝ:�ޖ2�+�\��}C���\ryU�>yr����-�E�p�2źlOØ�?k�1�+A�㳘c�|�̲�Uss��F�ܳirϔ���w"���ͱ���6��_j�8r��b.i��mY��j]��z�PιJ��Zھa�Bc�W��dn�/1�9�Q���F�S�"�Ӵ'�-֯c]ڍ��o���ik�+�O�O[�w�����xE�� E�)������z���sҷ�\��i+n����w�w����oԼV3�;l�����K��w�GWOC��G�����gK��������y��a�Q�4�r��]�Kv���%[wP���c�\�@Y����M��/^�={u��A�r�6��/g����lC��u�/P��}gu}�h���gm��"����n�
,�wպ^t6�����g�Ы��$CՑJQ��O�i�~�p˨��*}8�]>�,���w�"U��Z�ԥY��3.d��P[(����v���+�z˝"�;β�mQ��3��Z��2gJ�SEFUr�Kb�ǋoga���7���}�/�q֝]�uqe^�+nS]ͼN�#��j�+��I���g�^����
���zrE��cr�֬���g�_jßn��*�������\��.��8�E��ޮܾ���M.����mwӳ�N���,!B�6.�y��#�>�r���V�:-�S5��܄����߻0vϺ��p�"��4���AQq|d�[|��X�J�z�>b���4�uQ�Z���3�x=���;V�a��IYsi�aJ5k-�D2��B�ssc�'1��ÑA���V�4_M��9����?s�A���Dt�z����Q�{�x3��f���s�	��>�Ȗ�/f��GAe�^]~p��p@��f����P�e
lF ��b�ظ��M��s��-����Dp;��d]*���@�c��S7Ý\�1C�׽Wŝ����
oB里nk��k~]C�|D�v{��_��?3��:nB��L���D+~C<�Jr�<0����s����A:�'����3��<���5FT�)C/1FM��c���nr�{un��Lz������>Ȼ�c6�JY��Ty+N�hQ��/F���׼$��r�^��%s�sX��
�:�+8�k�gpN�Jʇ��ﾗ����\�%���H�|��Ж�o��[�z�t���������(�ˮ�d��a���{0�tz�!�%Ρ<��z�!�'OB�-�~͍���W��JKr�cw���-��=� �)/O���Ԡ��{K�l����[��hsoKO6
���7%]h0r��#v��W���׬��-z��)��a9�|�h{���YM��y��g��Z��էVz�7����d�"ݩ;�_.�(�t[��/W�ޛC�n��;<��}
:!��6��_a�	��(됱�	n�O<�opT?3��j^�{jI�L��Nx�=����ر��Y{�gښLV6Ie/7�x��8����a���MrC����V���e��7n���.��1���:J�`�{���f�>�ӎ��2���1H=�W����4F�4S�Ps�i���S�ǅ�-�$x�Wk�x��K�V.�Af�$��¶�Y�u�k;!+�b�Ⱥ���u,I:K��\�J�3C����:R�SBK�����&�޻Ώc��@eKH��=}-�W(�%]��䝁�{�%����ڂ�+�0��Z�,J���������@��{�A��L��0�#��M�	�l��i�{%E2.(���B��u���J���F�����	}B��R��clv�nvh㲈�[}(�+���:v��*[�n�[�q�k�\�]��5݀�us���G;��,�/`��/��v��]ӛQN���W�\����auwD��|��z�;��+x�} �����ܹ�����"��ڝ���X�N�k��J�:�2��\�u�K5����q�ٍA@(J㕷l*���؍�6+�,��3��� ���7����
�ԍ^Q) ���Îge�u��:�`����\#'1-��C�-��R��w�m����xPn﵍ȩ.�5U��+{g֢��f6������[.�J�.��N��L��S�Zv����̩6mpN�͋z)}��֦G�J�6Ql�@��wjfZ5K����(�U�aU� ��FV��Nsgci��_ue��t+�t���������!��;iޜ�W'�8���Z�Ix�MZhiL�J���W�]\�uڷ��F+uo#S�gt\fq�+y�V\�x��L`=�t|��g��xF�ێ��N�r�9k) ��]e�e�u�	��I�`��'`��5��ךl^!^�9l�Y������l]5����,|N&09��Z�ur�-���v�S6U��#�u8�͸�r��uq,����t�P:�����pdܗK�������:1�;�k�6u��2�2b��Wj|q�8�Ӡ0�f&!�f��
�B�V�-tK��'�r2�e�Nq�R�(|c<I�q1�	twKV�I�/�u�osfY��I7�c����+N��_p׽Vcs��d���fV]�eA��NQ��[{��V�\[�Z=P��`��ʛh�Hf��N�9��p,���uy���|�+��)ʉ�
:!�|o+nV]&�Ρ�(BwgS�x��l�Am@�T��]� +2�6��G��m�κ^�-U��9�M_^��80�>s{�=t.��d�)T�"��1�����!��d̺�wl�g =�������j>�D�D�̢�;j7��ԆR�O� ��Rh5�pf�}�u6p���Ƌv�}�(�*����{p�u���J�L�ih�[rZ�	A��s����S�h�ѝv-c�/z�[<*��ݣ��A����1��N����d�f(�v�+����Ϸ7)0�tá�� �h
}!"@D��V�]�WO.��R��i��:���q*|�f�A7�TX֊fƽ�åL�; 6�ݣ���u����S�;з��wMX��6���q�+��m�Ơ����IX�#l[��j*M�E���3Q\ܶ6��ҹQ��W+t��[���o�yՄ�Tll�/#�s�ƒ��F1X���Z66��W�x�(����Px�k���Ƣ4mF �k�6*4h�V-rۘ�Rj��1�k�`��#�#E�5%ssE�n���r�m�F�mr�Q�j�mʼso���F�X�Q?�<z�?ߟ��~�6�F�S�-R!u-Z*nݞ��NM�|q �Y� ���m�ʾ#�x&�d�a��,}��^m3N~���k�mz��Y�xr����F���&���b���Wڞ���;�b��sJ�Ы*��r������Z�+��lF!�m���'F����d^���x���۹������v�>ι�Uջ/h�B�g(79e\n���ͬP��752��Z��.����]b�_z��ë�J��7x�F��5r7����g�]��	_�U�ۇ�O\]K�==6��=�В�_�u�Rī�y��)�|��e{��Wƪ@����6��GbP�������a�]��xr1=P�K_��2��O֛�hq���W�=�C}cs�5�HJ{���.^�p[�ܶ����ר6�����AP��%Z�[z�/	���3��t�(���=���O�T�mAƑ�q
��`;�w͉�`UG(��U%*����ݴǁ{v�+E5���w�'����el�%�^��^ڶ	��̭��V����ޕZfL&�`t�+vf.�5t�F��_7d}��d�z�>w���e_�!5-�b#�@u�÷k��WR��mkR���{��,c�E9*���U��w&��v�tX̎�T�m���cnXm�����un��؇�D�CJ��ˊ��E-հT�:�wN���b�qMn����7N�MD'%���RcK�Og ,��.{e�ao᳅'��L�w_���m�U���rG�j�d��C��i�s�%���{g}�%�(e�vϘV�k����ྂ�c
�8�өj����=vd�=�*ۑ{������8t�덉�(^T�5QQ�q��U,1ڣ�e�}-ܯ��~�v�or(W1Ŷ-��o׺�<�������F��g/P��B]���EҮ����*m�6H���FZ��_5�(s�CX��؍��]�v��šz�F����zD�[Τ^Eu���˺���[�v���~�/;�.���ϭ.�8��-]p� �����Oq$��'��㳬P�����Ƕ�����.�@㋘�P�M���gE���"�ӟ]�N��Zi^u(P���Ն�Z�gGCv*]H�H�4VS9�@�Xqx�Bl��e�Bs92��E���瓔�a�����.=���l9(�ȑ,r�R=c!o/�.{;����Nͺf�%]����S�w�g��ǿN��|�텲��-��.�)�����/�=E����{��ʵ=@���ڄ��ö�ڎ6�[��6����z2���Z��ռ,�^e��=Gl�揠�В��|eO{E���F{�x���7�ۥ8���8�S�[C������}~���!%�R��v�0�x�x1҆�њ����ְ5�ʷ�.���*�_j����ݮ�/����a���8�ؽ��Y@�ۯ�u���c��n-��8�|;�����<Y�*�����u���˯e����u|�쿛܇l�4���'�푚�7���ؕ=��q_V}p��z�q��I4�zg�6�K�٠��Vn����}9eZ��֑�t+<r���_9���{Ym�<8�Z����X+1��TX�`q� c����e0�j��5���,��)?.��-��1���I5D����Cv�Sŷ+�T��h�I�G*v�FA (��Z%����W\���fYJH�|/�֞8�\9w�z P�~]�eX�a�nhO�Qx��9�H��P���۲Ba�jgLUy��J����q��0P�םt��j#˦9����}R6�n�u\���j�ŉ�NxK܌��n����`�ne�
خ��֤�mU�6����lF ���ZA�FȌ�Qw�yj���lxioY(�L�N�CV|�ʤt�٠_1���gh[�C�\�cw�qu�����7��iv������@�9����~�8�~�{�J,�t�����{Y��Eixq�S�w��+{a�X��K��q:��n�j1e�>y��>�/ga���BU5	�����^���^��g� �[&�P�m�1!1�'%履o�!2]�:e���uN�a����v�}|N��V��g����z_<ߏ^�}�z��l`_C�֬f�����z�!��'Վ&q+�R�y7���k��m<�+���P�"��m&M$�C/��bۨ��\R^5s���9�^��M��S4�)����K�1����9���F{�x��0e)6m,�ѷ�a��`��VV�Q�������Sإz�Ř��ũ���V{Q��(�<3BP�)��B��f�1��8����nT��Ph-׶`g�W�U/I5Z��\�S��QЫ }�.�٥	j�c��.��`75��/LV67��!�}�կ$�r�r
��{�~��xڙ��I������PŎaf^�U���u�6��h��>���a��C����r�Lr1ڄ�OeP�\,�P+5]3�g	���m�i�0и�'~����]�uV�?e�!���CmE<���P�M�?�旽�w�ľlc��Čb��́��<�����.�D+޳����8�s��+n4}X�ͥ�L�UR{qW1Ŷ"�sh=�8F�n	���F�V��vH����c�U�^g�� �Uջ/h_0ʦ��H������eX���]V5���jJ�Н�]�=�u����>t&s����P�뚇��#;m\���gW���X���9iv�Bz�]Hd�%g�be.SV)G�u�,��?P��x�i�����s�ոk=�}R1�OzzM����kV��p�u:�i˗R1|fAz�$;
���~�f�����-քa��R���wݽ�&���p�8\Թ���N=��u+;��~sWJ�f�R���a�ʝ��mpz̛8�M���i��!����k2��cA��r��,�f
j�ұqœxv������u��6l���8����l�ϷϘ��ܛC�+I	�S��.긾�jл}�Nv�&���.^���[���m��z��^��ak+�/o�.�7swaǯk�k4��Z�+j&V��R�}�S�}o!޷�%j�6�}�y쭔��3X���7@rs��_I�wJă��>�ؗnF
}��թ:��K1�6�x}Q���ag��Sr�`4�$�e-vO�1t��C"�x�X���
Y\ =�����mv�ͮ�O��J��Θ<Q�SI5�o��!��o�Q�wO���xWͳ�eϡL�Q�Ќ�)D��������l��ߦDﶫ�{���:�q���NP=,�okA�����,M���蓙�*{no�^�彨��p�0}>ਇ��A�f��r��++��͂��?˺��}}r/]��{�U�q�L�T��ο8�}�z_{4��MU� �L��&wҮ��}�N�N{)s}X�䵁-�U�����)��ԳήT�tᳫ�����2U�)7+^ �^ŶqB�u�߅�j��'�{�z��LJ��y�3�F���f�-J�Y9:CR�]�L���U:WfvU���}J�����KyVy-���i��t�'c�E)�qH͛�X������K���nsg��K��Y�ڴ�~����׾ȥ�!0�/�\$R�ȇ�N1���@���c�y�;}�0����]�����G[չ�aPF�v�k���OlZ�[�4��Zۗ�x�պ���.�{�r$�z��t��g ~�&�Ź�&�P�:]�OT�������n��g1�=ڧ�F୞&��5Q�9T�����W/U�}����0)Gu]��ea��'���g/P��;)��=���t�����gu�/̸��Rjb��Iu�/!E��o���w�����h0rz�K�^�^lJv��r����^
7�_�~�zǁ{b-��.ۿ�x�������'&�"�<�{��`���;9�����S|��;���ǝw��\�E�C�,�|��-�x���Xܭ�wFX�@ޥ�����]���]4��z�g��s��6-/1*�St֙ҹ����T��-��rʭ�h��Cs7��[ <C$�OWv��Ʌ���w��>z`�����R&�i32q�p�
�|�t}x�>����+^:����g^��!|�M'<��������[.�(l�>�p#���mo�_$Ҹe�vϘB���ӑ;�Fhou�7��mHç�ihF��5+.U�{����++��l�M�ݳ��W7��3�lO���=L���ѓ_�N�zӫ��(V���C�د�`G��Vo��(S�6�:����c']9�/]��ȒIfVe�_��-�X����H���ۊ�C7�U��(}M���=�����c7>�^�Ti�}ȍQz���略����ۥ�}|�;e��s��usP��4KZ/��h�I�{#���or�xz��Ry�v{"�s�A��e���Sc��פw�	]J���s��9jv�M�<�U�5�����˞�����r�r��塤E��s���^jy�v�]g�����yk�u{_����������|��spH�ov�M��.��.o������M�t��whLt1b�b���hm�'��"-�Y���}�pp�}�]_i�8ˏ�T�s6�=�N�����$&�cY\�Y p��J�w*��x��m;#17#�w��I.�<]�kֻ�Q������t���潪,;u�h[����	,s�<�z���i�����w3Ó㚅�+z9�6�Ծ{G�P��q��s*�������qi��0��ԗ���+\L�W�)F����z�xSk����huA���_�rqм�Sw2u_ND&l�cw����.�(�t��m����7#m�s!C��sj��b}�,c�~�'>J*k4�+4Rݴm�V)��-��
�z�BN����8�\�9.��O�0�J$b�7d�^�R�0id�͔&��f�G����x5~��c�r�L�Cf;~ʎ{'���/[�U��X'4:�k��ga�9�)���p�#�N�
��!ld�����`t���s�sn��K[ڊ�����>�©���+�4�_upH���|�ȥM��5t�r������3¹�(6�b�ٌ�k��eȽ�!�'r -׃�u��:iT�lՊK��.s�����]���aM����*2)LQ��Mъ��@�#J��u�-v�e��9��n����zFT�
�lyO������V!�*J?L�[�Ǽm��j7�#r�,v;&��ю4��U��b�K�o[ڴ���/&�e#��I��w�Ɣ���o+%-�S6b���q�S��J���/��{�����{�|��p���P˭��������Y��eD��z5Wg��\%{;}��Ϩ�V�Ӿ��GJv�L��x�\�_���ȿ���)v#��hzǔ�f"Ŀ-f�����|k��ɝ�oT��f��3��w���!W�;ye�oi�srЮ�'ݞ�,_aw�.���u��޸��w^��*QQgĤ#@�&|=M_!	�os7j׬�X�O�T�F����29o�]���_
�Guw=(v���N�� s{2�u_�C�{,����𣤖���2����R7S�:u!��ou�v����m���eͶx))\_e6����VSG��cI-���0yT9��S(w��N�*{��9�_�Onׅ׵G���ݩxT������Zo�T���]��i�%ېsQ'@����ȣ(�=I9�t�Y����s�9F�螉}}ǉ�+�<w���F_�ul����O�����6D6�_�d/=7�*{n�d�L�Jg Y��jIȳ�N�Y6m���ـ�����;��\������_���u�p�5%�i�|��];��� E�T�g;��i���]Ds��HS���X���hޝeHz��V�ӟ8��n���ݡǩ)� �Dc+�X*vQ�S��V�Kv+�3�\�I�)��!��;K�S���@��'X���ܤ�FF��3Z[*�!אJ� 4:�_u$�M���&���xؤ2gQD�GIvg�5����5v�nn�	 ��.�Ƀ���.)!e��i����F!Ϫ+Of�_fR�
�b-�Ur�5�[�c_Ѯ�})ŝv
8���6�9N���5�ژ�D������]H+�5�M��������f��L'����D�V��]5;�;���ۢS�O|�|�E�uKC�Z�oc|��N��bm:J!���n�2:p]�����ݺ%w.k�n.hmr密�$���,,��Y��R���ؕ\bQ(=U��X�0`Fw\��Gu�(۬{`*�[����.C�[�7J�`��aU�:�]�Q�Uۊ�n���(mM��x`��e�t�F�j�(,���1̷�֊b���]� �0S��f�*�aeBջ�$o���T�|sy�\�3QY���)ұb��C����X��rFnPѡ�Q8
s�fs�xa��=૱N�j�'��.ʜ�r�.`��1�O�mXtxY�nj�F'.����y+�7�acP��1�ɢ�٧$v�	X����e��wtN�v�+��؛��BnOJ{�,Y��VVʆ�RX�Lx(��{X[��k�%vr����2��=���F}�,��V Mb�M��!��r�,T�:�sr��5p-쥏�������er�6q�oIʀ� #���]9���{����ٌk\Ky�2V�ܬ��^�[W�(S�]|����ư�S"��%�v�1Dh�?�&ܱ|���ֺ�aGW�k��oGYy@��(h��/&;���j�7�[e�$�;�[�r���*m�t*\��9)T{@����_hg�.�!B���%�gZFz��>��-)$�o�+)���d�/�7�s�Pm�k�xeu�%\z7�7���m��33N��hl���Pԍ_P\/Z.�i��GhTu��ɵ�騬Գ�yv��`8ś��d�r�������{���ƞ�t��%m�s�-�m��7�v�<`;E=�&$���[n�`��1�U�v^vu9��ujr��:�T�^(m��u36�oZ�
נ�O���%�h+N��5���哉l�s���7�����X]FJ���v��m��ڶo&���Ԟ�.�tg�Pf����]���ϧ�>��fY��;.p3ul�F�B"��y�𮆞�/�]�,�@�$�<w[룪D�U���	"*U���l���s6Xw+�[}/%r+l^��#�͜W�KU�	��}ۄ��|��������
�s	�� ���f�j�v5�����3��-����������F�_��EEcIEO;x���6�F��ݪ�r�k�b�W9��(�cF��F�N[sh�FѢ�\Ʈ�$j1���wW5cZ�QIⷍ^#AN�ssk��*�D6ƢĚ5xںj��w9�\�6�IF�A��Z�����*��7#WwTF��ƮV6Şu���l�E�r��cy�F"y�\����.r5sk�܍��m?�?=��py�Q`�JCd��Z�n���3S�GO���
�5�r�D��F�����:��!}φ61���o
������ε��r�̡oVǬK�6E����}�;��uD����p�Y�RCLfK���x\�ܜ�N�uf��V\���3��x*Y�C��W��t����9ı�#�z��F�c��sv7*O��.��y̑�bhD��tn(��W��TbW!�M]�M�ό���As��[؎C��B���K�� ���7�/�}�<(g{+�c�U%n��c�{'�3Y��`��C��4�}�he�F\
��^��`�zF>���!��;��"8ȍ���o���C�}���>��:M���N���m���L��* �G��X�������W�4�΀8#��ӕoUT}<M���VV�랕�"�~|o<���~�~ߦ��?�N�,�_�zs��=�<���b�*U.)�'0�3���`�N�(�׌�;����޵�3��Zv�����$쉍qy1��u�./��}az��.�5����2���/�\��/旽�y�W�on3]�)W^˵�'�E��j|lQ�{����A��\o�rW�U
��9]�S7�=���[�he��*��~I���݃���y�����F�m@�X2���ƛ�p�`GY9jU�	��Q�Q\׌�7a��W7�XV'1��"�:��������m�7��ӣ��ү�T�嗙���}��bWz���v���cG'#���>گ>�����1�ad�a��/���^�D�j$�k�*���o�.f��&PSF��bp׷ל����Uخ��yH�:��ˈ�u�K� ���.���_L�9T;���oTWX��^��(�\����f�_a�)<^�v�goܮ�+����Ȗh0b9�gb:�Jy֮KX��;��
�*�`���S+�}��X&�%�C���h��;:�r��~�x���o� ���3_h��P�Fπ3�i��MMzck�.�==���{Lb����vu�������F���Ė� ��tWB��à@�S��Ixy�L5Q徐�|�.t��[�o�:��)��o�8	Q��0��]Zï?E\������/�d���/N*�~(gqA�w��G��h�׹�F��=�z��{�k��O��޾�]{�b���7�ٱR�d*
_�"�(Օ���[G1��w\G���ݹq����O�\L�������#�g˫éύ�lu������{��ąvٱԶ����Xim���W]�F>��7��z����g)>429I%gm��T���R �R����s5]��Q՚�wτ��\�=�fu��Pu�N���8��Gm��I]��^i� :���Ȼ�<��5�ۥkd��rѭ��G��
O����4f�3��7�a�r����7�gGo,aL]Y��6�K�hN��;:�}��j���Ό]R���,�7�'��.����ܽ�,~Q���^2�����v��榅G���q��G��+�Oq�n�����=J״�NrP�`	�����T�A�u��r�J���w�~�ʵ�������ku��{�p��#�Y�AҴ��E���q�_>����c�XQ'{+� �Of�*����.����]�kd��k$�ۙ�(:��������r-c_a35�=/����4�_k�Lϝ�6W����<�;�-I%T�
�Ά�d�]���]ee�վ�4���G��740ϏV� /�z�q�:��w�]b7�i�}�� ��G3�d�H�sc�4��{�,=�p;���R%�;惛�{�G!��z;h�����Y�9��h�X�:}��>��U`�UM�领_� $H�.[7�L���[~�"�[����̬�Tp��f��٘�als�������������,�"uc`��q��W׽�Kk�{��6�9��<y��v2ow\zg*{Ȯ�}Hi=�23���>����@�Cs�����Kb�#����ܮ���}砮X,i= ��Z���%@��<]����d��G:�ff��+;5�����Z�����U�ɫ�v�I�ַpk������ɋ��F>�����*��=H�VY�pض�y��|fk�I���C�§="j��+�Hl�=�}m�tϴ����{���q�uU%��RZ���6J����"��;��\�&�{M���=妡�j�M�O"x��s��3X>�q"�_����d��q�EF�Ϥm�JJ��{��G0��ea����_f�Hi��1����|��7�(`[�b,ju���v����N��Ԏ��!K쬋^�a���2�1]�0�UPQ���q�zרm6L�<��J71x{�`�^)�Lo�2U�.c���w�uf���۲Ǉ���IUr>�uh��]��R�`�g�U�;>���t/��|���neC��������~1taa�r<��׺�ފqKG�*�I}<3�ު�+ѝ�����}���N���?!�;�պ�k���.�
�`�跗��J'O|��>\��+�
_V���C6�g�'�3�m�;L�Y}��t���҅�:��ƅw�.��D5;X����u��^Wz�w�׬�kʔ,V�W�Zu�7J��|�}`��UfYb�Z2�enMW��^Lu�wWq^�����<�.e��U��I����3X�@��7X�P[��YOW3x73t�"�Y2�`��{��peIQ�u�����f>K��ħE�_W|�cV#��]H�^�'GpT�c���
�lRsԔ;k�#x��2���4��<O��Y7ECu8�wm�����@z�՘�Kv����F�2������U<�[�?@����h�g�ȭ��O}[]Z�xK���;��д�^R�zqk�x��F���A�F[4�z;�;�7.�iu.��8�k2�*��z!�s����zn#�T���|;A�-��# a��C���'ޜ���|��Y�3Xks����,�ⰾ#�{��F_�ul���<\ �ِ7�F�u��'zM����]Y�� ���+�҅���b_��/�{M��O��'=��Ux���R��n��Pb�ӾY���#�8����懫�x���d;m_8���L��<�Ak,7�P�U;��73^��sJM��9X�;�]F赓W�KQ��b�Wr-7\ON�W�Ec2�r�z3ݰ����Vs7}�=p+��}F�'��v�R�fE�⯱��ez�#7ʍ��cVv�w�Y��N�6y��{���C.}ν3*�>9>zs�>�����z�d��{ �Y�3��Ξ���q��U�F>�:MǺ��uHͅ�1)?s �tm~,x�;_��˳���qt��N�s��F���/��w��ݖ�iu�1Sٴ�?kX�/��ȫ���Gq��2e��pA�Ey��t9�]X�| �b�L���#ru��V��;8�O���IS�k�+����ʗU��'w`m��y����)F�3��b��i8pj;y{p�����o���t�	�����ߍq�;�� ��������˖ҭ6x��N��Q�V�'/'����0T�%��>��7�a����\K�V�V�tٹ�i�k�'v������zk�9�����'hr�w�9����uI��Գ7$eh��\/��*�}etW��O�d�P2�����I�C�ʡ�\atn���wk���Vk��w��������sې�(��}%��9��:���VտE��h��fT������1U���g\>S�����~���]Ô	(��r�o�6�����г�W�ݻ��}�R?8���S\f��>�'������{���A�����,ۂuQ㶗�+=~�7�e��6X0=�1�3���n�In���󭣟o�0���	��U2�s��P��-���v�|p�B��2���+㲹M{�X�.�r���3����
�O�D�Z�w�	l��EՏtO�u۸�ښ�n9P�4O�WT�����j���Hb���#��*j)@� ���>;�~^��'*V����gW+���c�wucd�˰���+�n��Wc@.]*h=,ʘK�L�z�{��4��̕]9�l��կz�]a��Y-�=����\����]��ܹ<Cz�YU
�����	vh�*h���:�ҏUi��+�d�i/����_t�7��鞂K�a����b�
�W��f\H����><�p���y��n;��=�5��'�>��\K�t�"O)�;6��UZ����I��N�;����:�?}��z�ܟ"��*;����5C.#z�K�éϠ��^�bU�Dh�>���s�+�������M<�У^S�,}�n=�����t2�63 ~�c`T)5���㐭-�_�ͱ��d�>Np���:��]�1䫗�������;i�wy�M�l�:��V�Qc�Yn�Ugx�7~2!�C��{M� �bq"��N.y:�'�=�,r�8o�nѝQq��y/�[T�6l���������a���=�מ�|�����)ye���:|�q����wehK��]�l��k$�ۙ�(Ρ���H<�#��Us�۾����Ы�.���.2�a��)����8��$�_L��6O��{��W���3T�S���EL�L]t��q�x�����^N�=G��u�㗏�q�g�i^1��y����)ԕ	���������7F�����n�G��֤����r��w@������5ܾ�gB�іi����ԃw��C=�9�'�ɠ���R0���dXw"�Q�S���#�VAA�T��i�7�Kb�<o�N����j�o8��"������Z����W`L�<$�C*��>���sx��0{��c=�mv���l[��1�ڧ3j��8|a����<�$��&H�G��u2��E��.[���y\�~�_{=+|�P���7�wV��'}q�Ӕx�"uc`L�
��3A
���NӬw�>Ҫ�-���^HUox#r��>�4��Ω}wlU���b#�P&4��!/O��32�bh�Uq��\�ǣ�m��x���x�����@��X�K�KSd����3<����{[wގX���p�朌�̡kMC�m_I�<���g8��5�T>�q"��zL��a����Rؼg=6d���@Ub���F��^5�/n����ܘ����4��7��{K��6�!��u�
׬d�/B1�t�Dwh��!/��-9����Ϊ�q}ުQ@[�3QqǕO��	��=���L�X� �}������B��OTT���C��f9S}n�Ӿ��S�t�4[X-o���h<�z��Ǻ�t����t-�*$�GeC�O#�E�8f{sٵ��H6}��<O��~�ͭ����#ۿ`F���c9&R�/(���n�]F�jJ���3uHM7�t�Lt�u�tG�-ۈ_V����އ��z���`�Yݗy�`k�mnO��X۱�%'@�[��:.��ښ3s6�h�h�l�m��*�B�PEUu����^��p�;�<'Vv���e�.��I�9'���{So�z�ˬ;D�y���D񡅈���=mJ���_��`{ֆm���my��-}�M�'�}��*<>�����=c;�2����8.)�Jo�<���.���u��޸���׬Ǘ����9^���Q>�t��gĮ�2ǫ�gO��F✆U�����y1�»����]H�l�ZK�ve�u/�ǘ��MwvT��Q%Q��ARǪe#uS�?[�?@������c�.jld�W��N��s�Q_S�}/)�9E�e]|f6�yT;�-���Aq�������s��yN뱰���t��z_�q�m��)���|;�g	v� ���Xn�u��@t/G`��.׭V܌�g�(�g֞\Mķi|�}�i|G���둝SL�C�<\ ��I_�4mym�����@����+��>[:���ُ}���t��7����wƇr��]!���򛰡�����RF+� l�54/�s�s��K6�m��t2�Y6�����?]p�o�J*Rd�%0�!:���syZ��e���:àJ8����}��XdK�eYΤ�ig]_FOK�;�Մzv�9�#6]���J�]��.�cH��޵W���]�c(��- T\�G��V0�k��`8��.�'+�wH�ٝ86�F��ߺzS�S�erD~��}��1�v'2X�ĮC	��>�q�~�]~����v�Y7�%�9��x�Ȅ�Ў�/#�q�}Ǝ�
^��a㊱�k�Ku��f���(l���c�z�M�{��sq�|�_�ʌ�E��fxB��Mà�ay^Y�{���ħ��i#���?1�c���G����7��;���G�k9#�7>���Q�iґ뾻��N��{����h˩�'go/n�Mv�7�[���\%{����;�5�O�>�?����;쇈�<�K�2p+��NY9q������*S�
_^3���/E�a�gr�y<|v??Ԍs�Uq�ߧIݺ*���8�Gi���+�__zp �]p8u�F~�d�YY�NQ�v�;�u׆���.;^ܣB�K~3��~���s��%�"�0�l%t&=���,�~5����K��\����ᾗ��sʐ�\�J5���A�P�(�#���fzU V�՛=�p�NᎬ\yHG�ѝp�L����g$�P$���:�wux~���.�8�W�s�ڤt��,:�r��hҎ��4�r���S����V�U�a�]�����sT?dY�8_�������YY]�q*ۮ��͙�d�4�$�A�V��v�v]=�4ʼ�K�����t�!!�Z�Sb��']y*�n�n���v���d^_����c�jQ7�4��p�B|{����X&���]<��B�Yu�`�_S톺�#��x��A����X7	��#�n�Q��TPX���&�;x�N\z�2:�Ed
\]]̫J�̕0�[@(sdO���S�Mq{#}Y'^����C���;�ڥ��ۻ���쫨mУӤ���Z�'�Т̃��^B�z ��R�W}SN��'4N��+��jT�^nvY�o�'��y����ۭ��kBϋ��w��̪�/D�� �n7Gm�.ɽ���c]%A�۠�H&imо׃����X�]�6��^ν���\�#}��g�ZF?W�K�T+}݀�������i�k�#u�a�M�]����Az���ߦ�Wj��ݵr���ԕ����/��v�/xcp��%JmWZ&��g6rj�0#,\�H�xG����.��y=�y|Mvڤ���#U�כ�	�D!������!��J�`�+�)wk{zq�qQT�E5�P]�d}���7��G�$�ǔ��ӭH��r'�v��5ci#�c4��0X��[�Ck������X�o��	4<n]��)�Ƒ����LW���p�n�x^�܅��]��-�-i٦\�Bʸ*r�Tr��ԩ��-Ѫmo��,EO�p#fs�Fޭ�huf�w��B�����a�ہ��os6�|Dc��n9o_k�[�j���qrT͍S��z�7�r��I�����e �^��b���5�<��bz�1ۙm��Jy�T����RVZ���]��`d��TN`�Q�xe�vLg �c��[�n��P��ٸ�%�Q������>�@�P:���z[�X��JpQtT4o(V`�*�{8f�f�p�(+��	�'	:T�W;�J��5��ע�T6؛�)⽜ȫtɺ�x��gX�!л+G1�558�K��
��24�R!chYŹyY�
���H���O�3{8��`` l=��M�8�/��ۮ�y��%�c�V�ܒs��m�$�/���d(>ǃ ��u������!�N��C����9��/ �o�,[�C�jݻ��<kw��C]���!b��2T�p ������d�\(T�XyR�No�v��� oUX��^ͮv��ov����!HnE|c�癋l z0<�Yz�����V۫r�w�Hzp���B���
[st�:V�kU<4wT[��mr���-�p���w܆�HL::@�v<�\���
�a�;7���N�]�z0�Eֈ����q�E���p���](��W�,����da���.�0nӏ��Z�U��]UP���ns�wc].nk�wW"���X�x�-�I��Qb�[����ܝ�Tm�<\���k�A�kŭ���k���\���Ak�ܣ�5�^8ZJ�k�;�#�^5ȷ���r<�^<�׍x�e�\�+�藀���N��מv�Z情���6�4ms\�X�5��x�wj6�뛕����#�׊K��k����&�V���U⹢�N��Q���K�O:�0nr)�Q��Ɗ�������??ߝ���f����L�@��BWa���ﴝ�[\̾�Z37�e#׆-H�7�wo#�Gl�z���by��]+�.v��}�(-s7NS3X�{����>��,���WGM�����,��-D���Nvn8G_�Lp\g ��Ē�OE�X&�C���h�oH®;:�q��'|q�Q2������=��q�o���td�����5�X�.�Os�=��5�Qí����O���Ѱ�h��z;��tۻwn����D�H�q%���0�G��C�P�;ӑ}<}~�5��޻�\I�`�;\Op>����<��KK�=��I�3�z��|�ӊ�����95x=/�ێ��d�=>�(:|���wR�q� oz����.��0�<�~;66��iSnn�j�y�T�����S�q}���C��Rz����q��������0��W�S�����#�r�{qm���׃x)�w�JÂ��_d�=��y��"��/I�/��}�1yWbp���)�M�3w�Mx���@�����w��~a٭�0����%[��^��?(�M�����XO�o43y�bχf������p��u��ސN`1�"st�{M� ���D��m8ڛ=�����5�}�i�9�N�V���olɟ�{pC��|���ٖ+n]��ᘴ�7e3�G��&��.z�^�]<�"�<�Ǜ��E��򳫫��Q��P}ǖ��vZ1��2�/�����D��/�B�'�$���+PBo�l�Sܦ�j�����c�ZN��dz�9�:�ZXi�{4uĐr�o�8�x�����xk2��ԙ�u����+B�˶и��[%z-�Icnf�gP��
�xI��^n�]Э�tGq���全�;����l���i�_����ك����h�Hsܪ׬˱�e����.�Bs��[��'E������Es���.���&j��x���r�>~f\���6z�H,�"ĕ(dUO'>���s�����:���,����S>��n+%�\��B�.�Q��㬢K�:��"�KfIAv�~� ���^��M?dۡ��9��S�{Ȯ��+�P������x�2 'Fc`Oź i\g x^��gCg�D�~�	�ܢ�66Q^y�q���;����t�͎��*�UOM�2 �5�4�Є(�r��~���*߳��ε�Ӌ�&9�=3���}�>��r:v��z��i�̖1T���,�\1M�uۺ�^�to�;&�x)l�e�>e�(:��}&���<x�q<���W���x�����Y^������ka��A�M��5y��׫{O��X8��Pf�KzfR�6=RTk��7�]�ϵ�����97�=��]n0�D��Sr�j�[��4s`v"lJ�vp�I�׉�dl�`������c�F#|��P*�aX��s��꾭�O֏１�k�Թ�TP^�¨d�(n�|�)#�y}��ow��U�)X�t�w����B�B}k��T���A}���aT2\b���]wA�t�O�O����i��`�3��t���7ѕ���d��\���C�NY�v}�58ȭc��W���nKU�6��e��Ad��ѝ�8�Ǻ�t���.�z����� �r#2a��i9Զ&��5*�.Q6{�<�g�mJ��'��p�;�<'Tgo�[�VQ�ӂp����f�	K��Zn�q���Mg1}N��-��<�\w��;���+�-�񟁯�̖	����WG�np���T	��T�8.��S���0���R��SeK���_}�8�3�T�VЮ@Y����4,��b�@3��'��C;�#��w Ty1�¸+���p�;��~Ԩ9���﫫�^�Ո�sʞ*,�J�1�ѕLI)��	�"��a���}�:�T��.�V��(-wm�}��i����NQf�D�Fcb$r�F[7۝���u��3�rf�Z�+R��e�xl3�S�I�ԕ3�4;�Ȳ3��V���SD��px��6�JAzj���ژyd)������L��I J� ~�;R��vt�Ja���|V��r��F��ܧd�EG���20�}t�V< (�E��;���[�A��_[���'��;h����U#.]��Di�%ېsQ'@�J/F���f�#ʳ���(�=�.&�H�o�H»:�{�i�]2%�yHI}��s򌦇�G3�L����P/ޞ�p^�/�l;�M�c�{M���'����}�$2��/�͓x��l�f�C���q�$r��H?���x��Y�C�m_=���?ou�Ӄ����*:p��Q�S���s]&�S$5bhD���7E����X�ĮC>��ۍkF���9zVf�b��9�9-�'��x�C7|�=p)w�����<��ۨ/q��{�{���V�ޭ�z.?���r�2u��zm�C�W&���sq��i�343��@�]^3*������~�{�t�v�I��X��窏��=�ƞÖ��r�q��_���m��3w�* �w�ky�V,t4hT�nk���Π�GyZq��'Gx����>�5��9�D��ʠ���w��#5:���{Í�_�/�i��KÝPŃҚ�pJ}<N_�,	���*S�
%��7M��3a	���ԲN(ә�.�]�t8_Ö���@���0��ǚ��Z7��ձ��z�B���ZS�4LY��Sz� su>}sqW3Z0*;�2E�c����(�D� Go��ޤ�vobc��Sݬ�o�V���Z��nh/nQ�5ҋ���=�ء�!}W�����g���(��->��s4��Nq�S��?v���_y� j�oQ�-�Ic��I6f��iy�y�W���]�{S��'���e|gPt��Nb7���7'y\���.��X}��u'�]sÔ�hc
�h��!QD�HzQ�P�;V���~\���}���G`6o��:�q�!�g\>S��\7�/-聳�[(Q�xom��Uzd�y�նй������1'�3�晛�����/O��K;q�W}��{{v9p�KY�u��1��l�����:"��ۘڙO���	�n���󭣑�#
��*����[���Ϻ';��Lo���ˀzd��l�Ger��,m}�ף��{���<|�щC�ߺ��{��霩�At>���uD�ꮨ��jY�������TIxy��P���N獮Y��'�����(Zj��z�=�3��q�ՠt�\Qs=3����F�����s��S5ˏgM��v��J�f�^�qC;���zM{�ގ5��3X>��%���g�d�\b��
~�΍�E{���j�Ȃq��5��΀q���o�6 �" O>�?t��ץ�;{<���f(͜O+���G��O6#���r�&d���5�s�pK���ϐ����&�}zw�,9�-��/$���衲���|�5|���K�o��e%i73�ڝ�&>��Eߪ<%��U�����+��eͥ'���ɾ�7��ޑ�]��i��g���=ᔧ��
�l�+����ep�.�v��{�K�~�h��A�
���K�Y�Y�=9�}G��%hَW���ชs�����Tg��J{n,��؛^����
�R�xk�Ϧ��c=Ai~�J�}��'2���0��+^�t�ˌ� ]~������_E!���NW^�������4;T�om`���]�'3k�����u�ia7��+[���lF^���u=(����jȸ��q�]pƧ;��/.�B�;]l��u�X�L�ƺ�O����Nk!oѺ��S,�P���r��B�k�f�A�֟�f���q^�[%~^��}�cH�[$�������Z��r���W��
�'e�����+�W;�I�J�vqo�h��zU��eOU���t�>�RATg@�Z,\T�Bd�s�nh9����`�:X�L���Bo[���{�Ok#e��7�ݷC�q�Cr���Q%��&H�G��qS(.�[~�#"o|�������>����� ��E�
t*~���cٔf�(��G�v����,Z���h �m���=��7��J�"�wr�/+���d3)�=S�ޜu�0�j"�l��gv�]�z`�=��4�:��\y5�v}�3g��.��QѲ%V�y�v5])�����es+���N��p����(�D���e� i\d§
��p� ��y(��=�}��W+A|����}�Hi7��#n:�ث��S�q�9�M`Q��hz�"~rIx7����[�õ^W��]�O���}����ӵ��u`�^�W�,Z��@9�5Ʊ�>~*\X�{ �7i
���{�_��P�}&�y��3�O{�k 1�5nl-.֯\�]�g���GD�R�)�9F�ON�WJ�X_�}��CMUI��7�h��7�`9f�_p�J5�
�$X��b�����\�+�N��D���Y��c�߃�>h-r'�"0��k'�����[�}�3o��:��|r#z2�Tr�̕�{bs9�������4��ڳ��݆R��/j��uSG�c�g�4:rw�hm���j.��"N���� �z��v��n��g��^S9��Qh�7�Y����L����﷪�J�����}Gغ�N����Я�#��^{SZh���'#f�p�Q�J7��>\�;�gx�Ju��;�Q�T��/�j�������?t�V�m(�Qֺ#i|!��^S�_���y
�{����V�F�;�x�H��؎�Ɔ�{\v��׼�_�z8NVט9�s�I�z9��,���̠������sV3�pp��mYu�껬�؇�����	��8Q߬�C��1���[�	�����[�gN��X�����S��n0�P��0:��.�n��'�|��ĸ��Q��*QQgĥfX�|�b�g���rXdr��� ��{�t��(�U{��
�|�k���WR��#�nx��(Fc�K��������bnx���Vvff�fC,�_h��k���gD�9��;n;���藋��qi�$��?r�{��_����h^��x]"s��I��5�0z%+�>���s���!鿻H�}wý�p�n@	���.�zTϺUef�v���=�B�.|��e�����	n���3~=��ŝ��L_��*et]ڙ�.&�.jŷ�6{�p�B�ꉐ6`wT
_J�^�/�l2��!�齦�zgb0���M�{����
j+�o�*(jJa�1�$���(�0�e���	+a���[/���I��d�qg�g4��ꌀ����\�ID�։��k��k�Y,ugL7��	P5�,�7x�gǤh�w#���3q�>���޾��'�؃���fye�t_�sސn��t�rGI\8��}+Z6���	[X_��Moq�����ɹM6�_�8�4�^i��P�����4/G�X��{z��cԯDĻB7�/z�s�A&���v��Nռ��!�B�J��u���ξ��d�l��aO���co+�Ř�7�njWr;�n���9���a7W&����upy342�����V���ɑ�G8Χ禟e~��-[��;�鱥��U�<�.�G����>���t6�]C&n��b�N�yw���H� �0������td����=⾬���OJ�a���>�:�������=���*�y����9f��A����C'��}Gҟ���&=}��=*��
�C,j[=:�����ק���:�z�οUi�8N`1��'b��Xn����,�����^�Jwf��{�ޱ<���x���{WE}�{S��'��2��A���q�}|��Ǆp=�>�o�厭̮�:��^@R�K�k�xrq]hp�D��.;�܅�Q%��윟1Q���2+���jF�Η�Fq��.f�ep3���HG��g�?t�^kѷ/+��7%Ⱥ���.��W{z��{���."D_�� �_�PS�L�2��7}���O��v�gn=����k�W �+��l�u���d��7��:��hnb�S���X&�[�0{����LeY��{�tm@��y�].�n%�N�/�3��݆Z5`a1����oj�oP��٘3�{H)B��v\vʸMK��w(�G�@�r]5��H32iu�͂�'Y�7�����}�:Ң�v�4��q��ѭ�kF������j��9ʺ������k��DG�i��D������7�td��l�4�S[��ח^�ٻ�k�ҟx��yw>�s�7>�Դ��θ�7w��̲�����q%���)�����B����='������|�;c��ԉ�����Z�u{�r�fђZ7�#Kv�w
�XSٿf�W���FG���2����#P�!5}&���@�	�r�k �޾�׺f7���ï�c)����k�\)~7�ic�,ׁ��������������C�s�&M{�#}a��b�<��g{�n򌙺b���H���6:N��K�𮌗��߮�5uޘ���+���3cRQ�v1��o*�v@>~��Tpؿ��J��X���"����?,''ظ~yrX�j��F�Ȗ�%�8{���3@��tj����\ez#:����+7��`��G�D��+^�A9�9w*�tU͹��=i=U� 赻|=�OS���oO##�eF����]�w���`���s�u�������.�7i�R}�g��J�`Oh��;�t��Ow��eh}��J���,m}�����@�*�l��m%lx����ׂ���0�v)�&���=��H��]���۫�<����mt���m0r��h��׎��v�1%k�ٽ�/)����d��|V>��Ӵ�_R�m�e��z���3dlza!9�@��r�Q��8���V� >\�� �T����`WK��������ti�V����׎�-q�3s�)+6r�j����w�� ����	\bc5c��T�YJ�m� Y��������`[�t�+�P���8)��˫:\5�t�+_D{4��� ������kf���R��}:L�/p��]�}��/2t���X:�D;@��T�;���Hէׅ5�.6�mvI��C�J}�oo���	��;�����A6eW ��)��v�[�����}u�!!�����q���VA��F�hΉ�oqA��Y�X���Aͣ�XQL���6���]��s����u��8��2t0v�4�KBL�ب��,�g�ee	]=��p_KA�Z)�y�p��}{O;v��Z9w���(f�U�_�
��<3";�N�� �wd!�C�]�rM��e&Z�w9�7$΋�m�Y>�7x�����2*'��h����K�5������� �t���s@�3�}Tj��P[B�w`EQ���Io�p�J�Gͫ�BT��� ��<���W���Ƨm"-����+Zh��eoXn��O�^
И!�v[�Xl�}&1'A�1%�Z>ror�{1�G���{\�Z�]��A��a�6�>�lX��V5���[T��8wy䛿i�";$���fi�u��rG��P�z�V�ι����p��R�ᙴs�P.]Ko��$W��	�V��p��.¡�U�s��9|��Τ@o���=W����ͥj3��Ff�����))�ʐ����?vvnS���{�r��fm��%���m�j�ƱڱN�R�-��D�3��grN���]�w�+y�Siڙ4���:��Hnef�9m��'��kP�ӷm�C��W;t1s��}J.��e{����-;һ�3�v��;t�g�����[:֯�Txt͞B����ӶԼ��d���R\�3t�gWwwtu�d�ȭ�E�vR���sn����v�FD��R��ZTt��r�^�:��wZXo#4�c��p��&�]:�sO�]k�m�٦Ҋ�7׸�mF��HoCz��%֞�Jt���V�jk��Y��u�Ǭ���!7�gnS3����o@P�t,��r�]x�P;W����%�:�KZ�H]�]��:��{h�x��*l^���_tZt�ˈ��YKt�*C�����	�L4f�K��Υ�d⶚����m��[�Z�g+
��gm<�7��sr�=���ңfj�'z��Vk-؀<Ŝ:p��vs�x���ze! �	(xʸ�jɌ���n2b�,@��}}5�ۻ��b��n\�f9�-ss�0cTQ�ww�[��;�tڹm��ۼ]�[�9�dwmr6���t����+��ۻ���H�hwr�����s�h�d�嫘�Q����r����mr�x�X�.j��7w64W.E�t���1��H�h�b��M�kㆊ��nV��#0Ć��[��`�+�����^+�rU���ɉ,Q���F�&��;�騬O��"��>�+��(n�����c�:1�y�l�R޵Y��<�����ZԤ��[��]����p�)|�V�t7��M��JJL�|�oI�3��u�H���=V@$�q�s	qO�3y�[�xs�����U	��\y�'��%��RI�aW�gGI<�2)�No�X���vY�>���+5d�PغʫnK���G:qU��b��x�-IT� r,z�RU<��"��sx��0M�q�z��l��5��r2rE�˨����o����u�Itg@���z[72���j�N��u���=bGD�w���+�\���ztO�}}C��Gƃ0#�24D��Fz�V���
=��w�݊�gN��Ī$����ϫ�܎�CI�Ω}wlS���d�r$wsl �m{}����x�����h��@�zj<��4��/�}���N�wu���s�-ꙿ _�V�G�'#�I� ��%���|�K4T6�t��<�����{��C��"�v�)��il#>�~�W� �ʓ��H�p6�w�����2^ޒ�j�Luo��ğ��l���h��/|Q�pF?0-� s��8�c�����z����c;�t~L��JE�����_c�W�?qԤ����YQKT�W�Տ�叻�L֋��n,�1묭N@C4�n漦T[�ӻ��m۾�V��㜃�kH��@\��'+y����]Jݳϓ�7�3�p��]v!*#u��)��r��|;���A��)`R��V�^��!l�����t/�wPs=ǀ9������ʁ��d��y�'0�>��gK����3�~��v{�o�\0Vz�hy*�G�����U���Gt���w��=�TI�Ñ��uC.�s����pKz�_x_�\��}��>�U�����xM���w���^���m�W�ֱ^��t*�+�^9{���E�K/�g�cGb��І�⬱}�C�Ԯ�~Z����hfϩ��j�o�����¡Ο9�S追�GN��7�L�u ���P�#��a`*���%ָ���Ts'׾R�<�����y���z�n��k"���J>�ωJ�2Ǩ����#,�W���7(�Up���u�7y�����닮�:�hW�Wq^��C�s�c�eOIރ1ȃ����qx�ǝK�C�èRݻ�~.���߯���u�gA�|㶈����]�C�8�4�KFF���c��}N潘��hd��{�����>�~�5)_q�9<�{d��v*�����3���׽-�4�}EI���]� l�I�$vT
�9L�E��ֻ.&�[��&��*H¯��FbQ7�*e��<L�q���v���E��xoa�Wr��}�Cvr����"�䶲�]�l�<�-��ym9$-`ޚ9v�[bR��`![�/������]6Ō�N	(L�/��V�78Z�r�=:��������VƆj���S���:VY�������u��eP�* E�� l�� ���+^�}�aܿSd_ޛ�l��;�c�B���
F�:O}��u�S4��)T����6~r��9�9�x*Y�C�7�gxw�k���z����r`�Чz�}�9Ŀ����늸�5�nɇ�"T	׫��E�J=ۡ��~�
N�tV����cu�H�˕܋��q=�#}a��~B��#�I�i1�!M�]y��˳�V;��{�*���by|sRTy� ���Oy���їtٙS�{.\�~��oؽ������>��Y�����^�_���}���~���#2�eo�ʗb��j�\s�	��3���:h�XV2pu�^�FW�^����5�P{=+�E�߂�N�9�0�y��Q��5�>�';�
�_���a��99Bg�pÐ�)�r)t�'+%�Lz�}o +7��LwD�!2)��N�Sw�Z�>�?J������+=yKM�zt�����n�,��>v�O�� ���u$\v^:���G[���;ݷ������u]�/+��t��i�{r�%-�3ƠΠ�(����t3�X��p2��x��tiY��x#@J�n�_�Q��*Z�p�i9ъh�ȶ2e��+�˚�L�}W���B,r�;�0^���q�θ�X�wS���'���u+Zf�%v�Y�QJ���=�'o
)ܤ��gv�ޢ2�5��&���횔�{���7ePa^@R�K�k#�\9���ᾉyh\w=��r�(�Y�Cz�H"��^����w��˨�#�Q�	���A\@ΫD#��)�W:ᾗ����gyՙ�
���U7]Rk��Z;";�t�[�'����38�w�i<V�Δ �-�~f��nN�����΂�Ȩ��<u�:��:"��y����S���Ku���{ܱM_��u�uG�r���}�#
���ˎ��a���;�td�� i\������ظ�MW!�L�����=b�D�V���=��%�Bp����R�q��������y���N7O���M�����ށ1μ��8\'���t�"{�g'�� ޯw���u]2�%�^�d-��H�b��'hߣ<�G��*�<��⃡ϫ��GwR�k��f�
�޾˞>��{�s��#T$ ��L�9���ٱR��U���x^��~��ܛ��ɸ��z��Ժ��ڜ���H����{�;�a�ç:nx+>u+	y<+~�xim���5u،{ND�"Mw��2���v��g���#ʖ
��-CMV��na+O8j�B�JWv��GV�v�㻽չ�u7\ 8%�@��a�u�\���WV�VD�0�}�wֵj���u`P�̡�uLp�rׯt��(`�u��!k����6����r�$�>� ��롗�����U@ɇ�+��Â⏸���>i�5l��������!�=�^�FwP�q��;�Q8w���Vl��8 {��!��3;�K�2�[�5��'�7�O+GGҫ�An{:_)���zl>�Us�'3��x偔��Wx������tOJ��qE"v�ɪ�+�q�]pƧ�ӃR�/�p��td�ӳ��O�$2�d��g� ���uB�����p6��*�K�qR�*_T{*z19}q�j�.�^&���9%�!K�gC���S�3^3�n<U@W�G����Ep�;�\����6s�ꅷ]{M�+L�H�P1��ȱu*��<��[�3m+u���j�d�[	zʨ�h!�GS�%�_w;��}�w��T�p��UD�'�y���l��^��J���U����U�t[^�"�_u��9�w��E��(O�����}�(��DTf2>Aˌzgٗ���^c���Ȏ�Z��_���s��w;�1�ꑷ�v�\>���B⑚�z9F���G���NHE�����-���/��;S�Ӣjʼ�@]˛6�Ix�V0�)\}�쨄��Nl��,
��G�l����{&�Ik��	��׏!9����
H�y�uo��c�mn�뵰��<lIv��J=RU��ъ��1y`����OA#��qt����>��GL�Kg>�Րh{ޡ���lT�z���kښ�ŧ����Jfd�vԞSpH0�+d���4T;��|/�y�m�� D��>��X��s�����ŗ��6�Hj�V(K��Q1�f�{��#h_�����~��g8�]�yI��K��Ǡ{�C5~Qf!y���G����W��
�Ő����Uܡ�g��������UB�HS=��m�����ѕ���QFh�����Ĕ|�f.q�m��:�hNu�裺V�#i�����r8�G��r{�hj�T���D�c�W�A�^���r[T��.>u_+N�dٸ�����UU�}�s�q�gUp������=v6�vxM-��L#�鞺+����.&Z(��:V��&2�[�A�ܥs1/�Y7jX�_�.k;�d�lQ�/����M❋�Qӷ2(Y��S�r('1�\D�:�W^���N���꾭rM�a�ש��z�n���l=��:o�6N��eP3�*'����!�4������>�)���۩U{J
�Y���3��������Vd�
Z��F��q�vVq����.�>:+�QՉewiB��6w{�wةf��ڷ����W�f�d��;�Kќ�wڜ4�\��c��w'ĵ�9�������Ue��:�"��E>�Ү ����	����W��^.����"F�w �=(��ƴΫ�G�G:��y틮�6�OE�c���~�y�>ڎ�����K��֜���(���=��/.�-��rC+�`s�g��L�L�02<��d�v�M��F\>�����b����_����R/�Mt9 oM}'@����FAҸ�ֻ.&�[�-���H��H�To`��X�i���ϺFuu^��>͸!S l��@;�D�+{z�?DK�lǼ��kz��ף��zg*o��};�������uU,�Ȁ�D	d�4.���1���Ҫ�������x�^t����t�q6�� S�늿��t�IA�u�u*�zZ��D\]�=վM{n�f�kO��v�Gj޹ۮ'�93C"��Bz����$��Qa~��7���O_(�^�r<��j���+��e8�椯9����O0d{7�.W�oy�6����C�G��i������a�a~5W���}���~��uW��}��o��/�˘a�(��v<�#=�/og�:@*�g"6��	︤�`��Ԭ���'+��m/Vz�q�RG�;�]��^��[.Е��cJ��P�hm�|�MM��� 6(�ҿ��K¹�������(�����0S[��1�����r��o�ԯ���wPɛ�N�(��@��+�\2�^��0�9�x��i���*��	��>ܧ��h�T<6;4�2��~�q=�k�q�/�N�,�����7�ล?��,��5S+ǌ��׏�_��C�+���g�����"�V�{ޜ'2̏Z9���W+�;���̔����Ծ���DH�u�`���9�Gz;��t�;����{r����_̷���*���ǒ�p�qtWE:�7�W�}�����5�����WZ��и�{r�x96c��{��@�i��%)LoD�Zn(���d�c:�Ȅ{���}\��P������oj�@eL��JrKEJ' ��C��e'�Q�SH��.��Ȟ,�HPvo��S��{�6QY�}�C����	f�:�΁!J�nb�eq�J�'�^Q�Jn��%oJq���E�!��k:�9�0��>�}v�?q�<n�3 �@�;+���x���fZ���Tx����b.
�hz�����ZM�vu��뺉���R�����	G���W��|��A�]-�9�Afy�M�x�+y(2��.PY;g8{�Я���|��J�x���+G�̞G�V{��U�F�~���Bw�n%�j�۳_��ʶS���kbCS�Z��b��[�������,U�������wqo��A:��0�c�}!�O����=�3��c��؊��aT������t��x��V�Yr���&��d���8�!���jj�J���ގ57��`U&\������k�3��%M��r�:j ��B^'
������� �&k��L�w� ���N3qڛ�*��j1w��ϕ�b�:V#�l.���/-�\7��O�"�&n�ߺ��&hKB:!.�Ro����T�r��
#��Ta�Go]��~a�Z�%����9P5?(�~W=Cz<��]/nc�o�t��Dw\-5���+6>�LF(#ܢj�yxW,�!ת��M���9��E9@��C���eS�����2��;+��{.�z;�I�G��Y��.&��v��ՐZ����ﲸ?yr��+�q�]pƧ#�+B�.�C���!���pv2��Y)��4e�͉91��A
�YP2�v��r�R�)Ւ��\c��Ỷ�`��=}o����J��E���gC���S�g<g���*�s���ӆxnI�,�F�TmL�z���=[Qޅ����W�����y���#U�R�����^E+wT��S�Y:Ae�qZH>W������kޖ��Q��7���!���i����3`�����y�@���N�A�p.�;ױ�q�ݓ��{k��<;����ʯi����,�ԐUD���y.*U!UO'&�z�hj�����-�!1s}��;�����u1���,��s���X!��=R�IZg@��yX;8��������+ȝ��|֫���^s�g}�E��(O�����Di�"�T_��R����㗯yS�{���eG��ȅ�/{�$��n{N71�=��1�I8Wp|}�[~66�"�r���h�NO" D���P(d�z��ӿymC���>�����}ӵ��S�^zC/��6ָ�J��/���UjJK���鈈��ؚ�Xxd�Vh�m��Q�{��W]��1��k'�Ig���{�ư�|c �WI�2CV6�TK��B���zW��o�����v9z���λ��Y��g11��}C�
���(G-�b�%�^1�M��v��%wB�,���V����g������G�G?\�V.c�x�YGo�2n����t�d�"7�A���G0�oS���H_۾^�`c���ӳﻦ����|5B�:�30r�������&�ߞ�-�m]we�n��:���j������w�51�ҏ����� +79��X����N�&X�H�|@�3�P	�&J�]��z�(�G6��3Dͽ��O��*�V�g��|�Y��y0,�s�x{6ۮ\���v�������M��U���w�~�e�*�u` �eMJ[��eNb�:�k�F��N��R�ְh3�=d��l���4�&u��1�o���QLQ���q��ؔ%�gS�s�u[M@6��@�q�X����U�|�Mh�N�E*t"33���lwIm�'.�67��v��W�VTۤ>��b�oZv��w�Z��gnЋ�X;������nf�}�)F7�V8ǈ^���1���f����B�L)���0T�Ǘ$:�|�㤧_e�yuz��K�qon࡝rg�k܉�ڻ3�{n��9Zo-��7J�2�z©k���$��Ѱ��Y�X1b�f����9�J�q�36�o	�#�5���e�0@�
�+r�)Β�S!i�w�/Y�6P����f�I��Am̮�6�3PWD��	��:!��Y(Օ]
HfnGW|˟5�V���֥���� 4�+�su�83��(m%���]ݦ�M_<w�iC�)H�Z��l�DYw6���Eq������O�PWn�ft��#�� �}/eᵉ�0��XfKC�V��ȭ�@'ОM��>�_�iS��V�CT��B���������WL�$�&�L[�Y{A�N�t5�e�u����:�z��l^g�:Wgf�����*h��R|~�Q��<�6�n��O1���5����҆�*v��e����9�e:�kf�N�G��Yܩ�i���{�ĳu,����m^{�XZ��c�=Y���5;���oU�����s{����1�e��!#ݠ�84���*t �]��"��U	�8��i��dd+���T:Һ�0��meWo*��xD�O*��:O�����s�w�����Ԩ ^J,7`��A嶾#]��2n��t�]�RA���]�
��ױ:i���`g��jM+(�T	u���t�pMɕ�4��]���ٻ�}ү,Ct�*Oq���t�',�e�~D�$T��`��{�x��t��:��aJ���L7����o�������&�	+��N���r��s���ກ�[r�/�9z�E)Z�K�bC�A%����B��� k%�3(������ټ�Z�]����ڸ�̑e�]Kwu��tja�l��ѱ'un�vV��-^�rK�J�:�t���Vs�EI_q�	d�K���ں�a!c�l)v8-��N����Z��N��)����ޒ��ɘ ���mXb�J�%&��m�R�7��܏u��((�ٕ;�g@p�Oz�:Uch���p��tニޚ4��Զ�0��E끝
��znħ��r�;8ɺ�ms�F�5�
ˣ�u��ܤ>�&	�)Vj��ZMR�t�F{BS�䐏� #�D��ҹ�F�U��$�wW7��wsh�(�;��W(ӻp����$�0P[��71���x�ú�a,QQ��DEb��\�h�С�l�h)1c@�b� ���\��Q���Es����-.�r(��0F1�2W�dň�H%�Q����\�$B���2�&d�U��6 ����4m&�wh�F"(�-�����7)M���b$��,�`3QDL6"$9�%�v���E(dI,b(����6H�I�Ƅd4TTlQ�]��r��&B<k�6ɨC`L��׎K)��$Ԇ� Z�h,�2+���.�d�@��^�5��n��`��4d�$���7e8�)`���E�s^ŏ/}���ǛZ�5NER3i*����%�Eq%�CF�bAZ�BK�l՞�B���,rK�o������N�^�n��>��t����r�����aZZf;��Yp/{j��L��;�y���Vټݰ�����Lǳ��8�t�*t{�{GN�f.~��Ю*z�	dr�G�*@��w/^ԯQf�w������/+�q����ز�O����P�Lg����������6%a�[�����e##7���+���Guw﫩^���c��H�:I�3I��W(��悴gK��S8̆�wA��VtO3��������D�JF��̨���SM�ҝ����q�=���P$h:�d�㢜��}����;cڌ=7�y�2�W��j
�z�е�
x7��8O\) .��:�0&JF��\}��ˉ-�ϸ�)g�F�\;n-;w�2����;��ˊu|_�\���g��
�w���V���hm{
��xf@82o'=��,����0�����w	���A�̲����f��9�8���='���"n��ڮ�;w���,����Kh��ɏ����9.�����_	�m�W9 �ӧJDq����۳2ܕ�7q��:�6hwpƤ@�t�ެ�m���1!]���r[���;z哐*u���J��\��{���(0EQɁ�ɵQ��{mK�t-�!Z}|X�������x�����z��%����L�����?��{	�;����®�G�����jD-[�"�u����<�������D.��v[�D۲,S�TͿY�u�,ϑ7��Ԃsk��}^�~9��l{��\���o��=�fhc��o�	�bQ�7Pz|�\�1�p��P^Y��/��/r�����?(�I���|�U1�z/7��T1�}�.�\F����j�(�A���N=8=�T�'�a\j3�뇛N$ww
�1�B���	c��Tm�����L�_�]�k�q_�>�8��a��*}��p�GH��iV&.�2�D��[���-fPq��{`�~��7Ҽw�}]�g�ҳ�p��f;�'`7�|7b|�e�=��{VힴO���ԥ�)�>N�"��\��<���	.�B���4,�������o{�m]+�xAٍ譪Fx���pV@$�wMu�K�3�9�����;�Y�{��y���x��Z4gj:��7E�L�d�p1�R����N�!No/ Ϸs�_�Ut�{ ���߶��x���*y.6�@�˗�����z%��L�9L�r�̢��v��s�z��F�.��eMYB����z�L���H�諵��:0oM]\tn�پ����j� ����|pE��!q3)SV9Y޶f.�K].��Nr�+-�����z"�J���'�ʡ�S=�(%��ا)��1����̅��I�a��jFNO�Y:s���o��q����RA`�� nbIK�eT�\�����9�M�=/��������U�+���\c�zO���A�~�o�:��wgH��Y��t裂0�U`��ڴ<��hnwR�n;:�t�]��|fx� r��>�B��w�ݾ�p} q-�����Hb�o������=��ta7�ZM��v���<�ݝS��5�����2��41�Kk���әb$?妡�6���t�{��0\��UoMG\cy`>�BS����z�7;^S1p�O)hz^�
��G(��^��P�5w%�rX�֧l�5��Cb&O>�_��Q�C�T.��"��6|*>�+S����$N6�3��iKʫ�[�x,뙯��I�n%�ﻧ��]t3��9N�0�2p9=��ݢ��ћ�m]ޛ��IUپV}�l�ʌ�߂�*���>��7�Mx�������^R��0M�#�B��B���+�m+����=r���;D�B0�����u��;����34�d��djU;���N���2���{\�*)x��;8k�_d�[ֺ(�r�ڵRE8�<{&>���5#+l��F79=�L���t�O�r�tG8����Ǌ�eY��W�5��v3�U��9�s'�����N�Cu������Y�X.{.�-Scwz߂U�>��+�����9�
��Xo�-��X�mp*gx���-���+B�X{�ˑ��R��I�Q`���I���v6���@Ρ���_"�y�.�.����S��e�A����K�Ъ�gBG:��7|�|����({���U�L��3��<�3�r��5�d/��t��.�j�]������Zvx�>}=�z�\r���#}���E� �3�@(��<�)�t�O���9�U�v�5��|��O�z�xz;GS�%�_w;��}�"��R�x�ѝ�<og�J��H�����t,��>S=��PN��	���_��v��tN���8�6�k.;�f??-]��g��@��\�n*f��ߥ��=�W#��F#q��#~���)�hY�ֶI��3�=��jS�@q��r�cL7"*6_�+!�C�v���q�>��˲(�Eq�.�hƃ�r둶s3%��T�� 6J��zxdG~Y���%��EF|��ilC/;`u���e��x琜���'�r^�ZZ�"5����2$<������n�G��{�84�<�{eЧ�SU�;��I���*o"rGw9���ٜ���Tcc�;R���]\6�ţIE�S��[:� ����
A�PYc��k��}�N��?6 ���3�K�>!�{��zNB�!�V*%��t�a�}�᳔*�e����{��s�ݻDm��w&}G�鞁��f�"��+�~����[w�)oh*��lk��<F�/�:"��5����<ۻ����q`cB�|z7�*;�����Q[4��޵Զ�g:1p��T�Q�/}��
�����]V���3~�ӳ�dgM���U�<��kHM�WHލtIT��@�!���E�8ha��em8�但��x�ٵ��7��=�����bs�緑]�X�X�(��(�3���t�-3�l���H���y�������QQs��okT	�Of:WV���Q��w�s���F��;L�-��t�9�s�R�w�Y�/�x�mک�Ԇ�]۠;;w�n_ZdE��^�s�C3G�[�P׵<n���@ˋPgK�x}�ްq�aOs3iOtM��8F�茚�:�3ɮ�
���+�ԇ/X�_s۔}Q%GR�N�������ԩ����=�U�IH�WH	�;����}���i�^����K���H�f�g�u����I�zQog+`�f�͒&���Lg7�o���(]0����h�W���#��ΛY�u*	�Sc������6r|�������V�E��n���o���٫��攻il���t��9��v�fm\�R��	#��O�����;�B/x�%�#DI�A���f�ϣ�����/x�)<�}�m��E�إ'�����\$���4���g	���9���L�@�l�E����Kv����5��*/xUnf��^)vuH��][/�:pOpB.�@ـ�@�WJ��q_j1��q�N�^6�|6p���5�G��������@{=Bv����E4��� k`Hv�c�:8���\�_��_o�����6����c�*<_�3�M����}qW����jd��;�zy	�5�p��-�֍8��V#0��̟CC;�C�k�GwJ'�q�{��`�ރ�{�љ��w�,�5�f��z�Z7��A}/V#_#�Y!���e8���Rj�W7�|��{�I���}���eF{k�����;�..�:���#ggåNx�;>F��`gU�v7�U���%\���-w'FU�l����Ϯ�\oPɛ��Dh�XW��������^����Jf�}����yKgtZ�;���=�{�o��Up�����W~��\|�H99L�
�N)��b��b���M��F�޲�1����"ۥ~�]���e<vX�Vwu���CD�1$�y�b�
th*^qӇ�S׍�����:�wtX��-R��G����;��s�ye�]١h�v�-p�e$^nMeow)�%����iec�]�5�z��]�5iZ:���vO"o�g@�_o�}*�}���o�x�o��3ה����Iݰdz�w�~���F�摖X+c)�>N�"�r�@s=�:��Gлi�׷(�{��Y���|�!��N0b��P�̣�N@�q��Q���N�t�}ޮ�ֆ��?A�0������lk5'�n�T��r�(Ԗ�A��wg���&w��c�*<�#�6;t�^l��Wt��-~97�ԝ�T#�	��v�藖��UmEJߦt�0䔦6��3���2қ'��8D�@�w�����.�#�d�x}�Y�|�;C���᳂Y��� �3�L(�y��~���u�&DrEo�`.��Y=�`������m�7�aW�v+��}w�;�r���:�΀�g�u����ns/�9	�ot�����p����"�[V������Wg\N��N���S�ކ�j+�nQw4����������`�*	�/��݈��Hb�o������ՠ]^IWh7�r��+n���H��E2}=���l��bu*7E����a���0���������~�~���T��V~勑���"�S�;+IV�3c��ͼZ�^[�ʈ�Y\���N�h��l3��N�48/�g;�N��csr���!�%-3�v���o_'��Ў��n���Bj_G�թy�J�fh��U��#R��h&Y]���u�N�r̭Yu��C���`9���o����dP��h��!/W�W�}��vs����#0B�����IԝӬ�<���C5�oH�M�������_K����`����=O�y���.p֪B����RE�	rx{��o��C/� r$��2a��2�:ႂ.^�w���+Q��6:�u҇�.��Ŏ��c�zf��k�v��Mw�)Y���'=~��N��*���&��;��Z;Np��c�g�m�J�zs����ң˦�{VA�D2%E�Dȳ*�~c���MG{Z�wl�1J��B��U�S O�+��T��DK���^��h��W��\��.<�ǚ���?o�$�N�ؙ�0vGO�8��5�#���
�/�D�>��MҼW΁�=�G:�H�E>������.#���B��V̱�:��)��r����6;�w���&�&����v�x6`^�(�=�=�z+�� ���wK�<}jH*��@�,�܊#$���G��O������nhs�������v�gw;�����P7*Y�Q%���MPq#ؕ����P��RW�Gc����������mjB�j�����e�V�N�F��Iսԅ-}&�9��#�$��hp;{;��Q���q	��?d�'���q7�T�dޜ����`2+]�S��[��������4�`�]1VG|�Qۙh��8"�H�]�o;��Y�g��T���-������;��,�����uG]������lة��r�v�b��|�� dh��D!��$�ßV�\M�k�3s���1]+\5���G��o�~�p_�/�ߤ��iK�f"9�Li��4�[�/�n}M��c�%emV8|�߂Ղg%��t�`7��u��32X�RZ��@ـ����zxg��n3�K�^�ݭ+ánQ�:��'�<x�2WG�*W�п��t�S$5cj�D��4:�f��4��V-��{�]
q�H��ܘ��}g���zw��ȧ�<@�s�Q1�P���WV����u�ҕ�F�,�}-m��+ƼxyF.�<ۻ�~}A��t��f�þ"7�D�#���.�Xb��"�̕��3n�l���أi��c#亭}#��M95���s~��{���/��2�ZrI[ �4neC��Wa�/	�xW��cbUWa+s�Og8��gۈ\���=�>�bW���-��(�u p�FbN>��!q>+�.����߄ƕ�A *2�ߠ�M�W��X�eX�w��&����e�)�0]�����C,��j=��h��=�+��������}���'��P�	&�c��ғ���2P�ʟo1;��R��ʐ��{!�k3@y�;���ꔥ�Y��f��w^	֭�ftc�EɫQ�5��&�����}�U��w�s���GvIÌ	�E��'��
m�����c�t,ss۫]�������H����\�w����V}޸��u�1v��F���,Z�h��g���{y�W=���s\n�Gy49`u g�]����T��ڋ�F/���*�P�fc�����W�f�3���S-�rw�T��3��z#K��9z���s����#�Zɬ��2�����nD�Fc`���.x&}���W�^��|�w}^�3���O�Ԯ[ف�#Èvy�������8K�r Nj$����-�������o.'�o�B���Ufߛt 6����)������ei�G��g\���e�N	�nE��2�@n�T��
��Y,���s^�%�>�J���ُt�m���uD���wƃ��g>P@j����{F�`.���I�t��}4'�t��aT,�!�7����g��'_u�����,�	��Ƽ�Wގ/s�>���g��b@����f;nV��^�LtV�Fmi.�2�6��_��������������:�ֵ���kkZ�v�ֵ���ֶ���Ͷ�ګ�������������v�����Z�ֶ���mk[o�-mk[o�[Z����ֵ��km��mk[o����m�뵵�m��kkZ���ֵ�����km�n�ֵ�����m��1AY&SY4}&�qfـ`P��3'� bE{�ǩ
���T���J�)D�RU�D��R��%JI"%��"�"�IR�D%(J��(�PPPTUB� ) !}����vʶ4�)UPU	UBJ�$[4�[e�d�#Y*Sf�5�*	A;j"�(:�B�EPQ*m���Ҋ%)���P�lJ�*���m%��$�����RTdkf�l�)"T�F�w\B�a����T	JE%CA��[iւ�me4Ԑ)(�H$�P��1�  'u��;:���C����ml6����t��ʪR�9w4�N���t��b��g$l��V�٦���uW5f�.�٨�Q"Q4�(��"�  n�$u��ts�ml�[;��J�u�袀 t ]  : t��B�  	��(�Q��:G���ǣ�4z4F���::(
 ����{޸�R(	J��u[2�Vve%�   ��N�3�F��P�q�gw�ZK�����R�҇v�ųmںp֫f[M���Յ[N��U������S������pv����ѣ*���mlƔ��$Qx   ��Q�jG��M���t�t��u������w0tɴw��ҳT�һY�۴ݪ���˛v�[��������ݍ:�K���ֻ5)Π�T�E�gM[[B�x   ;�4�Nٷr����+�:7*Ց�e�Gw6r�����1���㓳5e֪WL��2��ۡ�5N��F욲bY��5�U�%d�;S�ni"EU4h�i6jO  n�TԮ�k�A��U��C�v˥��;�ʶ;���k:�:U�u:��us��m[L�)�j�v�Ӛ�a�E��j����m�:;g0S�V�]8u$���n�t���]�  �y�eZ�v��f�)��3m����i�k��]��j;�(�lj�I�ҝ(��ӕv�Wc�H��U��RԚ�gm�:'Uc�v�����l��H�R��EQR�� �箌��9�7fݍ4��u5�n�v݊�����jWvҝv�u������wu� �
٭m���[q���n��R�9�pm����[ITUfډ�k�mm�ͯ  {2���˲n���UM����Q�aӧjt˹�n�'v�b�)iCNWn�l�gl�wPt]ek��m5:�w@��v;k��(���!UmYS�
;Iu���<  wM[m�λ���r��uݻ�]vT�R��p��s�n۹ݥ[)���N��t��5vg4:R�u.m�nլnfp��R�j���Y����fU)P  "�ф��@h  ��<�R4b  ���R�i�42j�ț%T��  iB���*@ ���sq�H�f&��`р�)pa+J�_~�fq���z���$����ILB!!��$�	'��IO�!$ I$ ��}��[��?�?�1��ӣ�Z6�(+�7�9�eX�E"��#�Ux22�az�+PL�A({͊�<x�%����q4¢��͛��n����U�w�^
j�?q��V�T�j�+6�n��,M��U���6��n ��4LN4a�^ұ����ze�r�˙HF	��Rp 6�,���[&�V�
n�����us>�Ty�e��	x]	 �khE�=��¥C2�d8���|M�H�KfĬ%�8]���b;_ �u�+R�f�K��Bƭʇ�>9'�ˍV$c�p����9��#�Z�M�#��}�UgJm�r�x̓l�N��աSv�b�[g5B�iܔZ��H*
���ۏ$&��3Sj�nn��Cl�(ʐ�`fB!Kl� (�* �{��tr{KP�Qu��Wpm�4+L�6mn�[�c��z�5�h���i=v�ث�4ψH�/P�*��z��q2.c����w��Q4�!�[zȼ���d3Av���y���i�Y�A�%�Ë2,�(��9��@��yB�6�U��B��1"h[�!J���UIM�@�`�lz+1nt �)m=H];�.(���J2�^�0�+.�Z�n��i'b�V���a�����HxTۧ��T�N����T\֩����mS�ff]�f �ݷ�XZ��)�{XE^&izͧ)2À4��䘓$4�B��G`��H�딞6�nky�7�7l�As0���u����ŕ�{Эk�z.���2f˧&ڬCb����ZF��Ò�e᫴��Q�.��p�bGQ���,\JT2�I6�ܰ��F��וt��͚�[0�lAN�XG��
�lF�=����9P��%R�^���<����8�˔�kk6����@��Q�Lc�6=ǡ�e��&�)H\��!y�ŻQ,q�I��E3����*ڣ!�1,J��E�5���JO)� ,�1�YS0*���xv�`�
�.<n��)������مfR�)��41��Ur�X?mi�:�4ڥ��
7U���R�ZrIOGȢ�"��S�"4�ec9���[�T�ی��a�=������j�'�F$�$ʂ���Zx�2E��	
�~G(+Ʊ��9�z7�!��7��)�,Ɔ��YO ��R�A��٘��f��-k�0��j��s;z������L0��-=�-��T�j��嫺�t-�ăK1�Obr��jA	�GmZYXF=�V�r�qb�-U�]l�YB�:ڷ�Ze�7��T�+0n�Sܷ�966�K��D�ܬi�Ө�� D�@*z���|�+o!�$ԋ3#�.��FD7N�����U����%mk�+�! �3m��K�[�{ w1+"bi��M����EV�jEj�!�h�M �Cb���!s����T=��ۅS�G;�R���������U��+-]�V�^L��JB�`Ձ�����e:J�F�L!n+P���-j�VS���qw�R��a$�Ѿ,����:���WK�q[���U%��m;6��bT&�7��7&�����2�[[@S�L����,��\�Yw�x�Wa�S/a�-�b�����9��ʗX(�i�!GA��nh��D(oP�?k�v�*�U��q��Rl�.�F-S�mU�)A2:P�ه/5J���5�S]k�����R�5NP�X���d��m�+�qѣE�γtP��On��7@�+a����L�76^
sHջJ�&�ʥ� ���h���	�۩��Җ����4櫫)�9Q��KW�-�r] Pƈ��c�
�k)]��ڵ��m
ю�����tť�����+��Pݥ�-�R�'���V2%���2�u��փNm[V���DԬ#.]-�u!��� ��^�gcv�����@X��u�@t��od��PۖAx�3���,e�q3�m��.4�	e�T��[����L��"���F��uzr����I�ZZ�Ħ� ���V˸���3Y.߅M�bm�S+ 0���:�p#v{2�b��X��Q�m�w"�z�];+Y`����*	-ա�A1d�5v�ݐ��7"��Qjpi��b1fn��["��w)�����5��i\"�m��Փ�B\�"�.�\{R4���[�ZԊG0h$:n�E�OJ�5*���]��Aޡ��b�X1R��f�ZS� M��qAf�7vµy�Q��QZ�;WQ�N�(4�ݠӺd�
Ź�O4[�lX��w-!4	�B��Ŋ��w�ɴ)�1�w��\ 5�S�SnA�7@��&�ܽň\ǳ`U"."b9������U�ej�ZP���C'Qˊ�f	M0�v��.���(�iA��L4��,;_!���nPl�o�ur��&�$n
�Gd�-�=�dŭ#�(eIj�۠mǶ��A5d\N����dXv,[���+a��W�E��5ET�dcy����4.�Ք&��Lc�Ժ��@4i�zhn�[�a�i6̧n�f�!�k�	��έ��3C��^h�3⮑We���k�V�|4�j۔�SU���W�����F�y�,IP!�DM�4�)YGXh�Z�m����hm%A��uŭkDb�c,��-�&�B w�~z�G5 ��.X�5滹�9AQ�G.M�����+�CF��4�*V/&?���j��o�MZ�&E��{�Fib�ެKê� �ˑ�V��fDh�-ҦD�E�6��U��@��VP45��k�M2������3oa�Ys I4�M(���%�v�G3p�e����Q�Z�k�`n��Z���Ϧ�u��c-�uz+f+n@��9˸(l�o[t��#c�K�6u��Qy+[T�B����D��=�����o�H�`۠/*Lb�\
��'qk���t%fe3�����{�A7y �t���/j(ݥJ���'5��,�2ލĐ
�+m5Gł��1i���1��	�NSɛ�uW��`XTGpT7�^t��IxsRۗ�D	�������%:
)�ѺJ�ܧ�`��n1��gp*w��h���e�a@��!5��i6)�6�T���ݝ ����YT�P���gkA.m�jP���*B�@B��iJJ�6�HVԲ�P�h�J�u��o�!�IVU-�	�:�2��V�i�"n�3(�+�)�<��T
¨��D�\T*�AX�S�V6|����H)A��$�5Y�0�,�^]�&5WiT�M�9ou�@ނ4���ٙ���G�n��aȯcG�[�v�h�v��P`���@�X�%'U��"V�cw�T���U.�^hF�Ձ�%��k5s�oD���Osp<"��H�M����v�f��+�V���\ʗQU����q����sl�����#�͉�Q��"iV��ZJ��T�L�®�`qfV�%�m�%�&�%P&]f-T�Mыe�yja�bm�qõ�@�gV�eL�UӶ�v�̱�ME��i;;��n�K��O�%.�(a�t�#�%�-Xυ�U�+~ ��^��5hK]dHЬ�rL^�4J��>4��4lt�J�����ב'��5��f�9H�ۑ@޼MyyiJ�DX�FF0֭`�yNZܣ�h4N���3j`�e �X���/��ְ�k\c�0�r�Ȇ++&���k	Xa��e@BgH��4�q��[к;����;�q;B�=w���r�edm�`5���E�WYux��ff��mf��tZ�-��@RT��T�o0-�����/���%`r�R��͹ssr[#B�
�X6��[[��H�ح82n�0��f�Պ�I����n��d+P�V�Z3,�Y:�MH�R��3�X��b$��WN��ojڵQQg,){�pj 2i�Pɐ���ʚ�Rm*�-�"�R6��l�%�鹋,�W^�"�sV8��d��Gb*��#bF�4�[� ���	�SI>E�Z�蜖�2�#��!N�̀,[��b7P3���+�c���V7��b�����o*b��,��^uE��e��������,���> �pIN�6�)�?������ӭ8�uu{P��B`��A-��:��73o+~���N�D�P�K[�Hi��t�
��څ��b�:�ĭz%��	�M�S�K�Z+^��p�2�������P�eQVcL<����(6s[r��F\B���H��V�k$k`Y���lZ�6ѽӆ$���8�Y�����܄L�?tḩu��ז5�-�E?�H�<?a��o*��-��)�R�kL��bzn�ȉ��r㼬ْ�,�	��1G^4�] ������Ue$A����WG�e�2x��t�XfY T�(=����9���[�g�,9��i�wzZ@���`�^��)(;Ѣ;J3��[d�Vz连�M��nbvS�sj�=�)�oF�j@4;�n�yJ�Қ��K�t5�R�	A��z2c��R"հ�l�+&��&����gfL�j��U�B�1�i�:�����t˚��w�Y�%fԺ#n�{IR�`;s[�H&�B�P4Mا�Z{�&K6�q��(���jBn�[����4�h��*��M��Ӽ2@�}�*Df,P���La
S8��*��NݜM�I����n��Һ�wd��o�V���1��r&��/6����l��̲t����L+ǭ2ژ2�/(�Q��ѻ��1�KR�(`�4�L��٣v�V�a�/@�P�Uv�J����YX�;7
E�:�4I3n����J�4v�ӋD�r�;��b��F�Уj��7r��&4^��[��.�T+,0��̳�
�6� M�x2nj�֧WM:�.���!c�l$lj[�e:;�[�cpD"Ɍ<�m<�ܫ�ߍYUn=�+�={m�CUjhM�i��YI]f�
T-��KX0P��cnm�Un�$�f,:��Ue�a)����h�{i�6��3Z��o"��n�ɢ�3+n��q`z�6��0S*�4�2�n��;�]�v�j챕�3�EwJ�еM�tp#PlP�/n�P�N�R�ŷm)��rf36�l[��;��\�j��	={n���퉋d庎$�j؂&�����0*�@kl�n�.1[��Pݺ-��,�Yw��p]1�RCR�iT�w�n�6�ɫ���؃
�إ��D&,�r���� U�L��IEH�e�j�A�����Z���n�Z%����2kZ̨���ڑ�V�f�{C�ډ� ����(���J��J
v�%H�
�9ki�8�IL�R��tEQb5	�&�˼Y����L�����]7Yf:ܠ�7X�T�e'����cY�!���wU��f|���r�0^�A�{�UM���lVܰ�	�課)kc5��X�T3*Ľ81��L^�@����5�S^�e՚D�4(���ʶ�ź
�2�)i�l��whZUc��b����Wj1�eV�C�F�)�'Mn��8j�*�c�u3���M�1�q��8ZЂy�[�����jdb�^�9��ր�y���e�:-V���`���`	X���
Է7�I�RWz��v��R�(�0`�C(hc��۶��uڔ���c5��Y�)nl��Oc!��3:m�7��$K1���J���[g��e�N�[�1��!��2Ȣ�H���t[b
ȯ�Vj�kT���oY��5x6��Y�Ӗf�L:ǵA�5AGp��5�"�2����kP�k��U�dXݬe6�"b�a@�=�i�rYa�j�i��n�W��F���l�ۡ�á�MeU�`Z�k`�N�--T��rғ�)b�_ۢԧ�����4³�#��w[[R��O/b��˹t1��V"��^M�?,�{�)[�2◕&�kUյ*����f�sJܷ�ɖ%��ঔt���m��:go�ڼX�qm�W��]*
9L`
����f��)Ie��f��zQ�#���X7"b���R�׻�K�w��:a�yv�����:���[{N����qޚ��b��]�wh�ն�mǪ1|���g�X�N�v�-Ge���#&=9Y��u�����P�E�[Ճ*m�ԝ�mJ���X��kTq��P�z�#-j��`��SI`>�]W�8�����66�Mc�h[��fk�藅`id�&m�)��d���M�Zzn�/n�7YT{5[�)&��H&���V��M��L@]]1׼��˨��-�D����S0�kC��M���gh$l�*[��KF;9I9h��c6�B�e�i���7D�f�9R�ȫY��J��.bާH�t'��j�d�I�թ�ϱ��<f]n��r*�V��@�����T��R=1�H�Ae�2�G�!6�C�ɓj�Ӣ�"fQ�u+E+�Å]�09����z5'U;�r��h<���������Sܩ��+�䣹s%�x�s)�.& u�0ÂV)fgE�v����Vi��:�9��2�I�ڠ�nL�l�Y�[��1��Q:��cKPHL�A��KU=xJҮ��;�\8���T%���N�uw�,!�:+i�F���/*e�Ê"U��Q��,eeN�N�+M�hT�Z[e��?a�n?�	Z(�-;(�?����[��d�.]eH7�f�JyJǷ�7�M��r��Ce��о���RAōŘ�7�^;���Ҳ��xV�����u��t�r�d�W'�t;�Ԙ�"�#�c+-�+J�Q:�k+x�R�I�n�'�UeZŋ�I���}nuG��]��H��]h��B�TuN����}����^'ْ�rw����.}�^�\�2���<��K�K.����$ǧÐ�B�ʲ�_�s��uU�ڎ���5�x�������稳R�`�8w�0K%'ՙ�w�98��ZoBX/%�A�+B̄��q�_f jgT�R�<'N�ė,|FvI7�J��f�	"�.�l���S/㓲K)ͬ�_b�{#hMͻ�T�q#E[�{uJ�y���S8�,��kW��(��^�Q�_u��Z6�����g���qD[�����V�]��Ǘ_Jhђ�yɊU˘:�֊�,WZ�0�4�p��P �`�w+f:7A��:#E�պ-T��P�Qtq���C#�5��4�5Y�8�
��`^WZ�P���xt�mv@������s����U���|��l1zy7��j�jS�wY;]���V��\���񼉕�b��
��K~ǜ�exY���t��X����z�z���1�|�����h�[�O���,V������U4-ĵ�5Z����_T��Y��\u>e�ad�<�	x��E�I��b�ڊR������2?����p�³�a�.�Ĝ�y2T0�ʘ�3MV�v��DP>�a)�:ݢ��,��-��,��Sx]�%u$�[�9
��<��F��]49�9��-�o�yp\�o������*v�rgXO7#�Ҵ�ww�<(Ȗ=x��<Y�B����+��][ӹǃ2(�/�]�n�B����Ql���Lmv�_0�++���m��7Omu���p�V��nr]!�,����H�m���V��-i2���ګot+�q#��k����$.����Yz�����ZlG;�,^�XZ�o�},^I �(㛠���l����}ʎ�.,<�b'e\�U�e��PlK&<~�u�/|�*�]!۳�F���-\�!���N�ھv�V[B�N�N�]f1R��%�݋�!��3!2Ď�b���{�Y����KD�9]@8M�-w-둇B�\-Է��p4��Z��3�%��NȠ�&��H�{���v��l]^r�yގam�׫�wj�O~F��,�`��O+0t��	g��O@h��nP�f�ǅ�1�N�O8\�l���z���n�5|�Y���ZD��y�t�^*��7Q�v�gO
:[Ē˽}1Zx����u�[��t=-�/.� :��:;�d��}���E�[�b�]��p��
�VBe	b�(��Y�.��Qi��!���	�y��[u-��F��\�n��8k�7�J�1|]�E�?�E?��ٹ�6�T�k��}�����jݨ���Xsix	�J�� yd�$Y[�}ȌJ�i��o�iAKo,h/`��^��C	�+�B'�wd��������E�>x�=�U�b:�#�:x@�qۣ��F�Ww$nowk����P����Ĝ�:q��u률>F��}��-���T��+b��}�Wt��B�6��f�YNm3���n�^֮&>�իSöԷ�J&�H�K#8��XK~s����|�.�}�>`qR�H���ܫ�"��]���r�ٕ�[��B�N
�����ȂP�]��r|7cڼ4�:��y�#؟=�Fܨ��{GR�a&&8!�Q)�:��A��glR%$LC��GWx�coLR�\���M����g1��g?�����.�W�T�{}a�\"�qי�O
�y[���N,���Jm[��$n����=��|��0f�;є{"i�n��<�a��X"e�!|�6�eϴ�w�V]�!̤Du�v������to4�.��Gm�IN�]��,����(�i�'��*����t���͛0jh=�|�#���s�-�[�� ����L�N���������>�N�u�Jٗ���Vd�ǔ�3J��,a��.�|������B��|B=tiou��Yzc���;n�e-�����S�ݍ���`X��U�HO'�����w�P=J�4�7�!n#�"�,��<���H�*kh<3S��2t��Z�ŅFD�diC$���w!y݀uu��f�j�*�n$�j��	�4(hy(�$��2SN������̳�GJ�x�.+l�8�
����f-�w|]����t� �����(鑊)d't��/n%V��e�C�S_u<�5;dG�oн��M�3��M��	Bi�����ۭ����j�P$���H�u���: b�{x1D����㾖���^H��d�3w/��ae``��-=�`4��Q��J�м��5�.�$�H�
�����8��y�B����rwd��"P���ٮx���X��-Sư,��n<���p��i�0���3�� ��a��
�Wy��ڱ\��'`=�Qr,T#��E��� f��7뿤����1�p΋L��1�l�"�l�5u���ZF^	Zy0x�=��(iE���w��Y<����c咲%ы]��Rԥ �n1��U^�y>a{p?hĖA��������d�Վ5)'hn)l��-e�5�v�-$8uդ5^�K*���0�7�a�5����x����/o��b)�3x�F����冯]�8`���KD�����t��
�;�ǧÑ�h�n"H����S+ܧ�FT}�Zr�����zD..��cy\����d�cb�N����z%���8_*��x�WÊn%oFelVF��ze"�����/J�U��刳n�[槕*�R5��k�Z,\�'~/�F8���Wv�Uҵ2s��fj_�Ֆ*P�T��,�	^�®[�0�����g���yKlq�6_g��KF�O9�h�C+7"m���cc�U����ɲ�Gan�G����������[�뫴�[-��N�wm���3�@IY���[2��b��5@�
Rhg"Wv���b�ٮ�bH%�eF�S��U�Q��䯖HF����#��e_S�6���\���^�s��v��p�&���1�$c�+��[��!���YV��ΐ7��5SHPJG�ܚ��8a����	��0!�:+�]݃GP���,�ܝ�ܮ-ڂ��4���ؚ�$@�DS�%I`\�aO@�H[8�L<]��5ڍm��췝�VD�`?m:���3��]���E�6��䩢��J��핓�j�0:_f�yD��u�[Wf�<�� k�^��7��U򶔶1�:ꂅi�m��[`�-�k�����/:���L����k�I*s���o)!^Y�;���4	BFp\heD%
HVn�؋k�vb�N-䱠:�R�nb�+{����}KN
�Z�J�(3B�{���t���ہޫ�>K�s�W��wD�7C#B��s�p^-�:�� ��%	 �ZO7x]��M����ц[��l[����_-�րU�����Cg���xaG�o:\J�2�z����
�㛕�^SxXw6�]���u��a�b�-pm�G�bbŦX�`	(����,��BM�DJo����l	>崺�|XC�i�x�ͩ�f��Qn�#�|ݚR�O��[�Gp��Uc���,n�WD{,hV�Ǉ7`� �ot_b�����`d;�j��4�f�3:�_\�ƕ�*Ʈ���uSn����r���]�A�3�q�!�������r\ꦅ�!T�;����� ��~�m��o��k[�NұWi��������-�2Ie�b��n�Ks�W�=�@H�mVc7:�Z�t�[�oc1s�AQs$����b��;#%�MԢ����[|ov;�2Ƌ.� pmi͇�>���ա�폞\L��D���^��1��AQ�nYv�Ȧ���¥��eS�������{��X��1�B���.�`�>��o3�����/o���;�/�u��>hw9�;R9��s���ְS��O�t���7��5R����n��[��ǌ�YQ[��"�:'��)���àT?KBN�HJ�U��}�r=�c�q��Iꕵ���ʞċ� J�t��y��{/��z{Cn޼޻�
:�hS���X�õ��)��d�]t��yȮ���5����9�
d$��QZ&�E{3��<���(��-E��.�ڒ B���/zr��hYΛ��3=4}���;�GeL<�6��=f�#C{ܾ�{��ǵ_#��;��ʲ��g�!�578��8����x�Xo770��'=v#�2��ݴ�f�F��Nu�,H25�ڴf(N�;9c�S��"M�Xo��WF���)�R KW�n���
]�m"��6dtb^����� ���fʽtf�]˚�vj�kQ㻆�_�^w�zJ>���3k}�+M��}��ư���s�j�!��Ә��no-r�Ф�lγ�,׊��{6n���P���{��HP.ޡB�<μ�.����$J=���]3������3�� �n�D,`FVn^6�f�����v�_�z!��Ȯ�0Tć�ֺ��_\K(!��K�
$�Z^��Vr*�z�N���Y)�YC��螔�Z�^f��%]t��գ���S$8��1ڍO�ԯ���>�wV��+�y_Q��}�%��͐��3.�����:s�q��*[��Z��.�jk���gu]v�J"H6�ו�s;c�L!�;S��n�}�EG;�]�J;
�����jv�=�ח**��جKƮp��w��.��b��CaqE.b��±4���Sj���+���cL�ɞ�+�� 0<�!���L�{)��	���\q�G*���m8W5�h�J�P�f�����L���*������v�����|y�r[I�]��ha��c���op�*�I���J<B𬦯���t�seڑ�تRD�sb�Ua��'��4H��RҶ,|���=�
����B�՗�g0�(v�z�a����2Nfnso��<��6˺����Q�
GRV�+T±*�tɪ���8�u��v*&:��pC](L[ld.�l=ky���vwU�Gp᳣���&�=��Р�(/_j�%�y	U�����rR��]�V,��)MӺTO9��-�jJ:L��Fn�"<͇z<�u
�9�n���8u6�*l���\��76�j���2��ͬ[8Q�8�X+�⭛w��.*
�)������/cG3��@]��;/i�DF��^�$[R��׎��nU�r�G�2D���u4:�a# 0��g+�ۜ��m�$���:ixS�p>�����]���v��+����`�(!V����c����Rc�T�]�F�88.P՘���CpٛJRux��Q�|F�Q����O��̺�����r�Vo;O�A�ykK���ڏ>�x��X��s0���-"���}���8,���u��Q�K���W`���e�P��&�����o7����ԍ�G+%#���ss�]��ۋ�S��V�{N�� ḷXb/��ά���N������Xc�U��y5�ū��ܵ�-����R 2���k�������{aV��Ad�SiT�+4a��O��A�g:��F46�v=�۴�@�����M�,`*Իܱ�u��P|z��˃h+���O�7�l�g:��j���Ҟ��P�C�SU�a��;s�Itݍ^ҭ����'b�V��aۓqK�ݫ	K�x��.��Y�c��X�L[[������g=���u��7&<�}Skg5ѩ5[ܧ�.������ؾd=�2wLtt�7OWCr�����uk���o������-c��c\��o*r�R�u��٩'\�c.�=�m���Zy�� l�
z]�ёc���q�qp��4�!���.�S���n�]s���9���&���q��v���BL�ۈ ��t�v�pe���+ib�or�	Q�D*�-�Pe��בd0�[{:�ܧ�Kgj�䵎J��m�����BɽO'�� ��1V�B��aluh}�Ĕ�T)����)��Gۖ��Y�[V��6�Z��Gs#��}�pz�(�k�C��e=4e)܎b��
6$9y���EA��K��0\��2�-��1i�KV%Z4;A2�7)g��_}ը!�L�*L7Բ���ݢ��KŶ�W�x"�پ�{
���KbQM���("���{�U���#�ޔ%��,���O!����T��"�E����嫢)�ǌ��H�7y�a�ճG`����v�#�����T�wa2\���j����+M>5��X�8K��e��J�c���7�����K��`47Vwpף��\�6fk�g�ЀpD��[;a���ݟo�C�z"���3
��+_Y�|�c$�ފ����)���}�k�\����Y���"�6��5罹��V�1��߅���&;�P<*ð̙�}:_{�}���md�
�\Ytt5�ܸ}�Z:�9IA@���'wZb#vYE^ޗ����eQ�hx�L_A+B��}��:cE�]'P�}���SڭiIY�|��t�)Z����g:ċ=�z6k�o3��� �s�����!s��iI�;<��
	%E���Yo��n�3ehO�y�h�VY��E}J+W���J�[�X���)`�Y�G�˩T(��6Y��O�/i��.�/p�8��츬s\�c<�����bbBޮzƷiލ�y��;��qSF�,f�4�KCH#6kk�r�d�q����7*-��!�ݎ}�}�WC"*�n0�%Q���Qu�Ù5+��O^��]�-��CiAoHy3Mhu9g;X#T|�;���&M#15X�<�_W\Jagx��)�Bn�[�+|jܱ�lZ㻛IsPp�mu���i������1�j��8�Sn��.���,��ѻ��\���+m�`��XDr��U���0S��� �q�1�U��ͩ���Z#��Q�[��
������I)����g���k9�9����������s�Ԝ/*&���D���@
�d�9����I! �����$�׷�g���_��/��M͈��^;&S���n����iu��NMk	6��I�.<�Qđ��� ҃ʗ29Eܧ�:�'4�!
���0af�=�Y`��׆����X���[��#�\(V-O`�:_�x�+fE)�a�:��;�
�{��ű�/�6����X���e`0�8�,V,�����hl=S[lg]��kEuI&6�B*�T��`���,�ESק�X� ���ۦU�%O���.��{�3]./�)nl��.�b}a�u�C��cI�hg�����)���rY�^�:�Z�S�\&[�Ȇϧ\�աA�+
��d����Ή�����s��"��"W�{���Ӊ���-�]��x���z��S��ww{1^�@���n�ia@Y)�}|r#���O��wyO��&�h�&��bلZt= ������J�XH����ub�4ۘb�� �WfZWNH@�Z�۲�X�U�7���9���f��6)]+*��ռ�j�չZd����2��.jl�RG�]3�Y�fΗ��R��:�(ћ�1���: 昜G�'�5��X�"�j�w���M۝]w(:�'�w��EUS��jp�*�c��7�V�A��2h��B[���.���7u�lQ-�m���}���;Qږ��ٝW�vNf�K�:�����J���ݔM�6!3�!����z$x�k�����-�{i�I�XA�m���N�3ie1���:��J�;�m�8� �w)���s�1V�v!x����0��@�oJp�4^5���]�ھ]��꺮�-�X�+�O�C+��Y�%r*�N�;�e!A7˳p�t�<4�vJ;�`s��+���r�&A�w�VP
�*���T�
��8�>ґ���V�u�H-5�=�$�u+;jS�-[ekU�[P�(^[��9B��[��T\[* �,Y��0���x+���2"}9AF+k��m+yX�w��79-�1�K6S�g�p�LK��P7N������Q�;�����ir3��Jks�W�t�1�ˮ�sx�e�*�R�W��'3-�j�٭���2�K��VoXcM7ut�*���v���8n�-,Y��|��
fI���8"��r�r�5V�����}�\��س�B|�	/�y��ƖVT`��Un��q	g89�C6��b7u˷TB.��z�5`r��;p<ll�������N����SF!��,�1$FF�;K�ؐ�}l�=��V-3�����e$+2�R��:.��g}W�ۓ��z��kp�|�Yr�uq��ζh��9�g��S�*
*ĵq����v{;o���/��C�ϕ*{vmMW(�oegU�^�,\��x������u4v��J�b�g��Ve�	�M�VVc���u��L9�0"������ܭ�f�l;5[�hR�ל�l��	���B;�6���t���
�LF��+���/��ၧ�ƥ�����oUqΥ��I����7 ��ݑv]貌�Z-��h3���ް����p v^r�F�+������.���{�U�;���n)��[ҹH|��z����+l!PV�M�˔�'�+v[���B��n�Q=�o�ak����ݔn��ɴlQ�-���M����R�w�xM���/N���@�����L��H ���ъ��Lg�6љh���	�KPT��������2v�
��쎶鶈��
������ӕÞ���x���;}�}�G�miU*��`t�Lh|�ε�+i�J]+k{lc5ɚ�u��j�$Gq}4T���.�ev�t�ڽ��ёV�|�	hy*�o�)�v8,�a6y�Z/K�f1�� {�B���o:�N)�x�^	.􉜴�}r۩Ue*��ql>RYrVJ�I+�sP�Ǒ�����]��vz�wN��d���3s��e�kҏ]a:m֑:�Z�ge��j�5�!������-�p.��FԬ�i�i�k�wj��"�R�|V�9���
Ź�լ+%B��cԩ,�#F^��j�<���A��jehHa�]|eJ{`�I���[�� �K�KZVnYJ��hƊAEiʻ��o:���;{�:��Hγ�kW=و�"^�KuCd�fG3�8v^��BK�5k����.
B��5h+t?��^[v�e�B�BXz�u]2���V�Ά�q�\냶T��n��p�/�6����r�'�W=�!D�#��q�J� ۱�b�ud��%�\�9���˭q+On����䨡`�Ԭ5�v�ıˣE��?�dQ��M�zM��p��n��{�$+e�9�)塡���TV� î�Δ�7|���U��S����(��c����8�&�[Z�P#.�9�,��p�ק��]�X�N<�'�^��E�Q^�������KuHi��ѷ	ƾ,�Y�����cV�[%=w5t�۾��m��ݬ<�N�U�,U�ݠ�0<-��oq%�	\ڮ�iȯl'ɫOC׸�bwEy6��k&\���>-�R�f��L�=��h���;���ޣ]�gs稳�f.�Mԫ�����\:2��)�Y
��j���u�U����Gcr�_M�˪5*" �^�V��=�s{i�����#���F�ģ�)4L����֮�C���*��߰\7��t��{.�T��u���/]nqD��eS7{K��LP��l�Ev۬|�gLrR	nc����u����w����W�-Uz�J�l�-�H�n�5��\�w��j�E�rn�C�u���"�E�w�@�+�X$M�g��Vg}�7{lU�`5h�)��}<˻7D��l�篭�I9'��j,��ܖn�#������t�����y
̾A`�f�gu$+��\T:f6�Ö�
vMN֗��
4��p;+�1^�M���;OZw���Z5�f�G�������wՏ��r�11ܺ�[ȳݘi��zy5P�25J��`�s����E�HA�Vd�ڦi\�q��`�!ئ�fbdR|�`�ԁ���̴#.��w(R�8�iPؖT��I#30j�4���(�����Kg.����^?�w� ���=��#��Q�J����	[�{�N���c�]�(js���|��u��]����,��4̧�T���hJx-�0aس�6x�%B�ǁb�xl|	vT�a �m�B�f�;Cticv���
���m�,�5�E�V���e��%�3P�]ݢB�^�"��[t�������M�eK��k��f�,�ۺ�Gj�#Qi"���v�-�����9Z�{A �q55�t������Z�
eV[\��&(����ү�͵��9�����.����R�c ;9h�cu�&մ���s��o��E�)�R���"b֦<fg*mK4h����$e���:t��圁��'Ku`ig+�k���l�ڕ��}���hFkB���`��P�ta��B�ژ;弪[�-g]��QK6��]B�Jy�]]�i7o�1j�+-	�����=�ݲ������r��v�3^��w�O�vv��R�ԧ3���%�+=�7xrƝ�:;�[:-��եfî��8�]nޔ�lo�EQ� ���v��
�w�ڑ$�.��ޠ��yJ�ZT3A�8�9�06Cj�lK��1y��p�Q��J��An�V�څ�fi���eM ����^$�>Y�ld����f�PC�PHZ��]�:�.�nً16���yO�9px�!��Jb�kN�e�}O&^ �����Qb����Gdc���y��`N�j�ol�Q:B����v�oM��K�������I��������sA$�GHǒ��}E��X5�H�,�9t��9��J�$h�n��L�ˮ������c�us�;m���ײ9y�H�!�i�Ӳ�=sh��uԐ���Ԡ*K8N%�wB\M�BZ��Rc�l�q��K�R6���F�������l����4�ۀ���_t
�e��2¬�f`��ڜ/�sAF�.�ctU��]U؈��ۻu��۩��o�9S�ei�8c��9���'�7GLH-�9�)n�v��p[�B�n_c�5�V^'�Q"��2Ő���Սn]�{�Y�=L���R���	��.�;q�JXC����k���WR�-
i8i:�m.�U�{��˫��<��%u5��X�&�T w9�3^��[�5�ЎZO���}�=��Ԛ��3�%�j�;���Ww�1��{�ަf_a��ڕ���)h��˷F�;���Y�S ܱ)�������b��w�W����W���._F(h[�P��f����6�������W�pL�������H1�W>����X��3K���eH��d;2�x!��`�u���7��I�i�Rq�6�,Ԁ�X�"���lԘ$��7h;�c\��ϊ��ɰ��:V�`�,\w��N�I�zs���������y������C���hX�v�v|� ��Er��bVm1+��͡���1�͉�]��ֻ����y%�����Os0�X��.�ǖP}{6�̅��9��OB�)��c �\�/��˩<���Ւ�D�8q;������Zɼ+]����vn�Y�8u����D�[C��n튂�ΔHkW���[BWpYJ_W���DPPa}�J���̌c"�,���ui<ce���3�n����+��4`�]��e��S�-�Ct�#��'�>��et�r<�P�а�-2�=���N��)_\Q�Ö��a�˷s�J�o�d=�YMسPd�C9�a���
�=w����3.�ofj4�\U��΁�Sp��EsJ��p��w]m��L��DY�R��a���w���1��kR��n���Y	ճ����Y�_��CxӾw�cv���a�H��;�D��`r�|õ{��gc㏻oH��R��h�s*��r��W4���b\nYxr��)/��'�]�f�1�=$U��r�`z"w�Z9f9��"�P
fS���@���ywzh���hR!�S�m�h���Ty]<,kGv�wC������V��A�\�/�s�6QPB�'>�T冸v����@�1�R��w8pHm*wB�rd)3,M��D��x%)Vݗ�'�m����WH��p����/�5{v��q�k����Jm�9���ڹ�+�2C{,\���S&����;���2�0��>��I��G4[MrJ��z�f��qƖ��� �H�n�w�@�W�ͺ��h����a8��	��P�d�5]' �Q��Mcc�����٥��B�L��5|5U���\"3�@Ko
y�hA-
A�cF'��v"_	�^Y��Q\�V�*A��^7�S^g��B�n�~G�p��#�jXvИ�[oE�V#=qNڴu7��θ�t�p$��O2e�(�f�k��Ӱ��ݒ�ћ�� �ɤ�{;K�-�F>�ڥ]o]�Σл��@�`��̺�&m2�KZWV�P�`��9u40� ��)���b��:��HRy�vf�3FG��&��S�ռ� {m4b}�5,�X�-X`����U�I*��Z0�m��@�/_gq�����s+��M�K�(�^WO�&ĉ	$g�L��[r�Q5�6)�D0�Շ��,Roe&V�CG�
,���
K\���m�1�շ��8��mJ�8c��.�ܻ����\7B��/p47�7Kwj�p-R0���Y�@�HW x;ݮ{č؞�{�Ve8�.��V�
rP7@ۧJi"��s/mI�����KsB��8�4����-�� �(�s���j��G�[7u�GT�n�@,GIoggc[o�X�S�L���S�@�R��Ł�Dg��\\�]�Q��� @�͖}�;�1)=�Z�Uh�n�
��[>X� ����C�c�=-:쥖xuu�e��]��94����")oc�ŭ�(E�v����9x�K%��e��۠�V5,H����gUU1DP�J�ʘp1��T.uE�c�7�+-����T򺥩`'(�[�@B�ǧ��'������@"R�3�Ι�@&�%	�,�t��Ғ��t�ۤ���auĩ�^����#�E��k��Á�
̾6;�̬�vkQ�Q��[I�Y��R��V�K�KpD]��-����RO���K|t�|�ș�8��¹+��7 Ź��B5'��.Ⱥ�e���ACr���7�Lȩ	�YEv�ИXy��X�*�	k��CwZ6{�Q*�:��K)�t�y���K[;]�4�FYS�)T� z���a���U����bzշ0������ILڦilx��u�J��Qo��I�uz��2[U��66'�U{ !�!�[��'!��ƫ���51�
�i��m�;�U�_Q�ݪ'���#NmVWr���G|�_umF�b��u�^� �9V�G��V�E��XF��ڶjk]Y[���5F�,d�֞J�M�8r��XܙQXe��7�$�ᜭ��:�
<��r�U}�P�w�@�p݇����:[F.㘹J�,�{�Xh���n�����ˋ��b�WO)�/1����(%6�S'Vf�o��2T�|���$*Ъ���ㄦ8R	�g�v��p����j�2{pmǂ��Cor��8��ݎʆ�}�#B�6���(pw��i����,��/q[���:D�i��^VՋ
K����L�z�ޮݢfS(�U�� �f��񧕋�s�"Wg�4+_q:���Q�!�k���1��ۄ���lU��9�i@�-���GW��ǥ�u���u��\��a���(�L���j��gQt;�Y���&�6d�ϞNQ��Aipw����*<2��2Yȡ�y�Z����������(k���Tf�gɓ�6
�V�����w&q�3x�*��/)H�o��X?ʾ�������|���v��-;n3�f>ù.���m�Cgn^Sl�sc����"g]0��G��[l�@�꣔�o�1e���u��g��-A�v7{�(n��ͱ�^oc��Nۻ5����&�����4��r����f��P��J�ҥ')B�O��4��ǉ�A���wv�{f0��K���[�Q�.�_b�E%���qHn�[�ԫ��E���!�g�������� ���w�f��۸���b]hԯsO]��i��}�QBQ����@y�*��ˏ*�塹\�]tNڶ���9�v�w�{��m C/rSe��K�se�c��lrz�ԥS)t��R^e�NwN�G�S�Y[�k]�.�\:����f��և��-,[����9Z7�P���˽��w�Ƚ#j��F>���L�]��(n(Y����x͔��[�ף�Z���a2K:�]��⍫���X�L췂��%;Q�2ŲS� ���w�jZ3��K2����@t��W��	��Gӳ#�|�Td"��ʲ���r�r����2N�d��SE�~�����)c���x~1��ո̍�
p�o�Ow��w�N��[���kvU}�%;J��ҍc�崳V_)�|b�bՍ:�.�#���m�OU�w����D����	��\������ʫ����5z��ӽR���U_0^P��b)Z��PYc+VڣQE��E�(�5�UԲ%V�DUJ�kk[*�*��Uh����mT-�P���h���Kh�cZ��h�Z�-mdKJ)Q��X�ѥIh�mEH�Z%B��5mF�V��Ԣƌ*((�(���,�hT�D[J�+mK�������mU�mR�#���TJ�+DE--�J�U�U ���2�m(�F�+R�mDX��V0RР�F�%m*�Q�[j[(�)P��hƔb��l--�EX�R�R��T�*����j��ki���E�+Z�"�R�c[lU��1Q�e-KJ
֥J1[AV�[X�J"��[Jխ���mm��iX��,U�UTDdT�(�V�������R���  �����W.���L{w�l�iih��pc�l4wXǉ�.���Fۚ/k�l"�ʅz��eϣ��u���a����sޡ���>�5d�T���_d�e���ίd]ڼ�����/���ù�oz��&b�tk���-SO 5�h@���8����t�}.�3���+�n�u��
��T�ҥ�9�Z�~�J]�N�����3C�f�3��/5�{�����\���)��kJ}<�]y�����^ϡ�>5R��
纏K=�7�:�n�㽞S̠�}P�׾Ms��F���J���k8b���,�6�X,r+<'��m6�����V=�uÖ́瞌�۳`�l�V_?kޢvxV��m�RQ�Ap:�؏����.�_Q��j�x�њ�pfѣ7�(J�6��x�g{�&/�LN�,������k2��r�{�On���v�L����Ӓ���6-kQ\0�������g8=p9sGG��Z��ħh�r�H�w��Mna�kIV q��D��i�Z��UG��S�� pL/��2�=�Yz0�U"�y�**�V�!�FkZ�ڲB�/iњ̒J�]������Ǟ�c��_h���q��ӽ�:��@s�wh0�cy9�jtа�<�	�wT�9�)s�Q��r�'au����~j9��<z�
�I�3�m��|�b����~ܩ$�|!~�'Z�|���^t~W��N�
�q�&u����S�[�}'9�s��~.�u�X��=�-�T"�'��	�&O>�}k��q�O7�����w`s�v=�A)�S{-?]d^痞̘���|�;�ǎ�cqo_s��wb�}����^��;�?��CK{{���(�Q�w���=��w��/����F�O�y�I)��Wu�ӿ`�{�[��[~�A���Uon��{պ�g��y�+�+绺z˜=/77.�ÆM�lph�cq����/�Րj��V�hݮ2��=."�t��6��X���=��z��Q�"muv�ǥ�0�T�lG�f�L̜�y�k�ɠ_��|�NS�_t�������pt+�9�F�
��v��^�E�A���)�Jz{2G�����}AK��]�b�k![A"��`��OV,=�V��D���t\48��}֝��|%zG*�=t���!y���z�`��������J;y|Ue�c���o��(�z�4�΢v��[ε��rc\b2\\���j<�����'J�;&�>��4ؓ����c2d�hO*^�vL�]k�W��+�ET�W���L{�sx��H�q��v�x4G�5o����+}٫:���PS��{I���f{s�ʙ�W�S���ޡ��)z���X����Z����ZWz��y��p�����l,����+�8wN{ro��~���x�9qQ������>�	`�x`BG��sgT3��p9���tί;�{͚�C�����D�5�-��~ݎ>Ĳg�M�.�t�U=�M�T��4L��:�B!þ[�n��]���3"���(���n	�>���v�z˛�N����A�)z�o�^�ߣ~����V�Y�Գ�-��#}c���{�:y^V*>f�R{�jnW�j��<�_�� �:����-�W���3���-�k��s(f>𷝐��;�X¡[g���u����,
�t"p�%4s���Jbxc`�(i��2R����R���N���v��%:w�e]�(�Ν۴�H��	M���8���G��Y��P�lf^��s.N�غ�1j� ���Ku�'����sRշ�S"_K�j���8_��Yz�}K����v�O_.�9����%m�y��"�2Q��_�Ƌ���k극f��v���A��u7��Sa������w�S�UK�)��W�ۼ��C+c���.�6���^�Y�{���HUS��r���^�s�+�S��-{�>e����U	
9�7|x��{~o��Ϋ������jd"���^�=i���箟��6��Z������
?f�}�=�,����G����J;ꜷ�u�ۤ���<��^���A��1��*�^׽�j΢����� 
���.M~�/6�S�,�v�?j�=ۛ7��f�T_�ґ���d;���Ar-��#��y����Ξ�o})Iۖ���z��w��
��y��OGL�'�������IEΌI����W����OX�)�ȃ��[!�:��� ���7�mҾ�cq��[�h�h�2+��Nߊ�uuX�m̌�KN�c[g.����+{��1�;��uhz#�ᒘfC�s�|���J�K�.d�k�ɘ�q�y^u=a�~��bd��*X���sْK�7o3Ҝ{�JO����Hew'�6?7:`s��3kA�L�~�eY�ݕ�=|}(�1V;e�v/�:_d��Q}1�?N����7������bY�ޓp�z�!U�{�C�i�ǞXfN�f`�(U�������|��V>�UW7_��iT��{�����l��[��o��EjɌ�,�3-g�>׸ܪ���z�쓞o|�]x�'M��¯���*�t�c�owx���+x9Z����u����=~��[-�*������^��oy�^,�qo�!����Ô�n�)�ͽ��/��]����%9��Rl�6<�(�`Aب͖��]b�U�/y��!���;�1%�zفwz=���W�2�}��p@��*
纏���~���c�˾���D���Y���>��FUt���1�d�^�����&�f��p�x��������]��=lfO&�^ڔ>������ݲ�u>F�s죢�G;~k>��^�X�T��� �*pL���:�~�4�Y*�81l])(v����H�Fa]��&��]}�2�.j#�k����ӥ��	���=��Ǟ��P~�9���������(��~��]XڰB���$�P��쌧��-��~]�����^�6yF}6�βn;:�̀x������R��1�ߩu�UY�)_���fSq�W��ng��J�0�9*�v�޾�'���j!c�r��c��=q���gF,�+�)��w����dy���}������_[���ç�=�����s����b�XǷ$���䊌�ѾF[D�_/-g�s�,���;��G���J�?{�ɓmWI�p��};Ǥ�*����ݭ堧��j��E���g]73&�S5�;^[t��s�v=�A9L[�{c��
'�J���:eҞ�^M�ao��w�I��\�.���ʖ:yt����\�����{�+b�Q����K��S���1{:5������1�^9+,b��쥗�:v�|�U�wr���:�unq%�P7�cjZ�L� �Ya��c�� �u�8�;D*��@UI��4�4;�.��oSyי�E)���]��p�@L���r���kj��Ǉ\�e�:y�����KK�:��CA�K:[��)����V��p׶w��ϩ�kV���Qu�7{�,��t��4��_��{7�~Kx=���M_T����5�^/e��׋�d���n뗾������v���s�
���4\��ֻ���Xa����b}�Nԣۉ�紌���;:Y�w����� ��<�,N�o���o�}���/��$�����7���/K�~]a�m^��8É�oJ���6��lz������)�F��{�T{.�=�{�]��~��K�׾ؖ�����m(����Osݪo�e�iZ�]�{ԯ��(,�Aay�ОӔC�;�2L�Qr^�,��N_�{�U��5�oYc�Sݪ�z�V?um�b�5��o(�[[���ޕyN�S�v�I۟[��6/ˋ�8_���8���Ez��gM`<w�	O��S��>��y;�{͟���qo�g*���$��}�C��*��S��i뗄%Iv	,���)�5�l�wi�"Օeb��5�Cԏ*�1���&c��q�;�|��!k�mU�VƉB`������>jY�;4f�}�]����4AN=#�k&�M�H��ق�k�u3�1��r�;�sn� ��-���6mI���<�v�{s���U�4���eU����w��
�P�j���_��{�o7�}noe8�1^�V�taSR�����ޗ�n����Y+jX�:���7����iVG�A=��q����^��4���D*��E�#]�[<���z�>��@���C�rc��z���*�D��90W��8Y{֭���9������*S�y��_��:}�����y��r.��yKʔ�ǆ���9'y�~�g�ߎ�x6V�1��pk��9��j�i95}/��m�;ݕ�|��y:.��yY�Es�W%���}����NS�Ҳn��Dg���s��/�7�
����<�2�\���w�[�
@d�<.m�Nz��"U��˫���S]��S�3Lx2oγn���U�k�{��$��|�{@����!j��6�5`�I1��e.r,��+�뫎���04�g)�Ï��GK,rd{��^Q�-Qz�+�D�a�v���d��
���C�%����3x�6[6�\�>��2:|7��Jt�qd#fq.�Giu�A��3�2��ZۉK󼱹<��2;=���A���(��^ߞ�j���];���c�\���L�T����^my�d~�8�]�򙒋����4��O��Q>v{Wz�,��?^�)�Bv����/w�ܛ��*��W�v��cy���$x�%��m!z�_rSgT���gk�o��OU�8h���u��>�|��}lfW[�g6�wMΔ�<^��G.-�Vwjz�r��o��b�hں]���\��c��N��&�J��gU��cw��\�v��ɻNT�:���}ޝ�wK�������jBI�^�F���8����7�W{�}��s�]ƺo�gi������ًf�t~P��y��'?u�{w6ۙS�{��/VS��}��>��6���igCQ�Ըr�^ז�v�E�����Kc S�c��3�A�|�[�� w[�]ҧ�j����&�6�zA��mTH!�]�(��u�;��<�\��]��e�nZ�P�i���DL�`�k�+�Z���P����M�9oV�V��n�t����j���[���Ċ���a�'[�<�Q��&]ߩ;�?b�9��j���+���T�ԴNz78>��G�#ϩy�ތ������C��B��K=]w��*��+99�W�0�^��>+t�V�j�^�Y�;����l��g���^��3�~쨖,6��q7�,jV[�U��_9磥{}1U��1�����}�o�{ǟmt��RmO{�״�����ޔ.��0�s�F}�V���W��3�gQb4x_�#���ȧ�z�ի'�S���w������s~�Q�i/4}�ٝ�����q�Fٞ�{ʷ���=%+�1�ש��=zOlg��1p�/?S�y|��=cQ��_�����Y���qA�� ][�����8�ǋ1>�gv�_s�Sް#��qK�_�/\���aj]mg�u=Z��^����Qw�ϙ��SC��9"�0�ѹ�-�v/�9;حR�<Hon|M�žj�@֭���u�R��6,Ay%K|�T�hR�=['p��;|m���:(q۔yU�QՇ���W��[c5����)G9D,�S����L���=&y7(�BW�U`���Y�e�~������&��r��#��*��A¸!��A����Xp�xWF��[t�hWmn�5ut�v��9�d�ټ�-w$����cg�K�Jͨ���aq��h�a�5��L��N&��7��D��f�yW��[�y�N�.�QH]����r!1���3;	"�OF����z���Rub,#櫭�׵�pgn�:�a51T�1U��JT�NΚ�>o*��_���]�z�˵&A��A�G;7��p�%��4�PV����v�_[W\6sO#}�`�0M�3��,n��׎c���e����0`n8�E��Mu}]��y'��*��pF�hm�:d]w/5�m�x�G\�W[\�uZ�V��[־��M� �oa QUz��E�7!U��[�a�Z��T�F��/+�/>&\���S����'j���5*]7qZ�S�gm�:K�If����j
cW^ev9J�j�t�4��?D,t�
��4v6-J���%D�.���5�A����9yP�:���9����ݸ��Z���o۹�Z2��Z��Ǔ�t�n�h�{�N�Ap�	]����'��=�R����B���]�s$�a�Nlwh����*�:��Hn�c�������T�s�jb�P�%���x�]3H��U0tٌms��I�ڐ�M
�xo<d�i�yǀ5f�V]�_r�s����D�!d�eu�z3��	�z��5����K^��k�[nO��d));��[Ǟ_ y��/�s{����Q�[�vW �j����)K�N���1�\�bUm��^sp�C�������(�"Le,N".TkC(�'U��XK���ط2���El:�ž�&�Z��^��^�j���t7����L͑vR���jf��a��u��|��|&�7t59jx2�2T��{�P�W+��ݛ��/�Z>S�.�-��T+&��o,êX/�5*[��� �f� �k.�+%T[������s��bQ��ס�^�-��9gys�7��([��"�.Ln����`�;��)�0�vN�0o9�yN���w�>k���Wu�)�f���W6�<zhw�_"�*a�[��x�>b�����|�����yR������z�[)K�Jv�0��\�Y��)��8�|�jZi��SB����iΨ�g���ݛ}��Zv��W㳥���/��pa����A�w׻ajH����4�5�d����N솺:�6T�q����ݼ
J5�D.�+|V�muX�;:f�|ČG�B\9|#\-7|l��<��ch�I�,���̭���(�x2�utuCo��{3��m��R����#�y~q��ڸ�Ʋ�+V�Ub�B�YV�UUDF1l��UR�+Q��Q+Q��[j"1+
"�+iV�b�Z�
�Q�TP`����2�*,#*Q�PAUQT��5QQ��Bֈ�(�B��b5�b�kKB��"�Z�e�Yh�eh��TX�bm
V���T�(���PUJ�UA�)���b�V��ʃZ��F*�b�Q�Ŷ��YkK"�h� ��`��%��`�E�*1m�����
�U`�*�Tb��
ZV ��)R���aJ1aZ��F�`��(�UkEU�"�����ڢ�֥b�l��"���)+V1�b��EF����PDK`�FТ)�UE"�PT[kE��#j����UT�[J2ڋ�J��H� 5xk�n�Џ�ŕ����ہwN�|�u�5�wD��v
�y��E�J|RɠN
���Zn�o`f��6�%�#���[���7��L{�\���}'<�;ۓ�yT�J����Ohn����a��kݾ}�I�r�1��+�f	��7�����ƕN��^�U���-c�Vw�_��ܰ�m�5��\�_��I��k���()�7�g�}��as��.��5Н�u���i����=~�
n��yS���=8s��yz��z���'��8x��_[�� wK���u���f�~����>�-��U�ޟt�����W��p�t{<��Q�u�����QN~iNS�ҽ��;Ҳh�}�6�9SE��k��>5��������=j��R~����痻nu�36��U��
s��;��󘊮�>��&�7�^>v�n5Y��]._�߾�\U]�F���X�
�ǣ*z��Q����[���T^��Z�3ò�So˦{T��G���Ҵ-K�����)�*��c�[�QȂ� ��3r��e�vb�鈜�mbt|WRUЀrvN�إ�_i&�t�M_q����u�<C/C ��4L�rX�^n��] ԸY#�Wl�I�Ѩ�;i�42�qي7w�n�����G��n"�5�k��{������$����
zߜ�a�3c��U���3ԯ����Aa)ʫ_��qe���a��6y�9�\Q�oNmV���+�+v�W������~UoyL�b��闣�KsQq<����;}JN��<ؼUG.#8���v	���L�f�S���Uc�󊋝���>w���5��T�d�Ӗ�^�{��O�	ȯiڜ/����OC����Ӻ��ɟ��?Z�;�Z����i�½P!^��.Z��:��#�dڈL֕[��`��]I�}�l����d����')�Oz�+jY�̏��7��!�cg��Ȳ�x��敹�8p׋��&��s<^�5��-��ț>X���v�;"��<}�>����*^S^򺞹hs��g1�����Fu��J�~A���a��d��;�򡹮K�觔���<��4S�(R�0n�$��h���<E�.�DL3Q.�-Cs=�I��%�^�V���^m3����ۭ~�U�V�5+6P�n�|��|]����DT�V>M�nV���'t'_\�r��;"��WvLc��o�56��mz��>���/��A��A읟3n�ծMU/��N�G9
�X��/u�˻~U�(y�߳��WndJ����*D�S��nn=L&����mu?=T���5���P��(�q���K<ߕ�:�F�S��֍&C�W�,�����;?{���ckܭx��_�G7��Ց�W�n���҄�s�Ĳ������.TL��Gǝ��z��߹�2V�|��{�*.�2��I��{�T�u�G����8�ҩ?j�=ە�z�}��t��9>����e�٤glN��z@��sG������w���z3U��;�	-�~�<�==&k�kQ](��|<����sa�E��=�����"�`��<��^���/߻������ٗ�9����$�&�l:��qά:�̬���N�u*h;�HVN��{��'�8�߽��c]��{}����{���5�x��N�Oo�T$��O��bN��f�{�d�$4[��|��6��$�4�d�!�ћ&Y'bé8����d�']�<֫�{������� ��;����J�kl�=�E�"ٜi�f�5�k�;˿	OqY��*h��_��m��{�)�h����/j|ws����\.��4��J�V�Y�. ��r��U:�)��6�.�>n�_T�������Ә�spn���c#YV�j�}�v;|sxo3ڳ��QU {_`��,�9�IǬ'�s��|ɨ{��&O���k2a�<�d��Hq�<�I�f��a�1��OƖJ`�������ΏN��p���W��8��hw��!�����,���>zɶM��!:�d׹��'P߳�*
|�P��Aa��:+�|�.�:��������מ�Wvt��N��=;C�d�M0�'?Y��̝I��6w8���h��q�M���{y4��O��!8�$﵀Y'��j��*���7�K{f�^O�؛��Iߵ�}�{)*O̩=1@�N2y5�O��P�Y'�&�>I]��}��$���s�0��v�y�L6���ĝM2q��=�O!��\}���_��j�[�����ϼ$�oy��I<�%I�VM�)<��'�̈́�ə����q�uC�+�C?}����jw�?$�I��q�,�a������:����O|��������gШi�h,���'�|ɩ��&�'�~��d�RLϯRVN~�*N�|��/�hN�8���i�	��Ci+�M!��d�+k<�ퟏ:���s8�?o:�a0���d�^� ��O�Y�{�d��~ɦI���&2O|s,��`fb���I��a	���v��N�����8�xǔYd�=ԻW���^��wU�~�}𿅆C}��IS<�2u��P���6ʇ�=�
O�2o߲i��&���J�{�E&���|�O�c���z���o?c�|���?k�>��ސ�!��q�d���v��e��/>�����<��*s�<�ĨO�&�u'̨{��M�|}���I�~�I]��L�_v�����]w��������M;`,?0�N�ݡ��BgT�2��I�ݓ�2����C�o���i�m����:�	���?$�'�R{��>d�g�<�>�{Vy��h��Ƃ|盧� Hoa�mV��.\�p}�Fӳ�k��R��K	�[�^��H�է:��Ksf�b������U�sD�M��ǀ�]���Y�8i8E�wU�ܤ�3�}�~�XY�z�N\��}i.Ԥb,�+��������������o�)��E'猚MbβM�fMP�N�2�C,�Ad��ɴ<��A��'u�'SL��?w�<����}�ta}����~������0ɖM�����>I���~�'�C�`�8I��eBm0���$�ʜ5C�,�?`<��M~��N��*jw��O0�G�_������U�����9�_���:��8�m���|��l'�{Y<�笛��$�|����I����+&X~CSC�e���S��<�3C�,�?P�'��3�y�v<����w���s�/?x�Iğ�S���B�|�ݧ�$�a���:���@�M�2~;�I�ɬ{�d�O$4Z2�|�hhŁ�2���)�I�N�:�7��mύ�^����>��\��6�d��(y�����N2{t?N��
��;���L���by'����8�o̟���d�O{8���C�l���,5�f���?w�|^5��*�}���Տ��I������P�'̂�Y8��P��d�����$�d�{��>x�i4�;�u4ɯsy�'�j�7�t�g�����]���t�	��y
����ğ$�50RN$�i�'Y�>d�����`:�ԛx�����4{��ԓ,��'��M0�����������>��g�I4�d�߰$�߷�T&NY�+'�g��'���u�ɐՇ�u�Շ�6���0u��_`�U�k���}��h��~��a��?<�����X��d�O�>�'��'�2�߰�i�^���:���T�&�)���Y3�R|���Fl'Y>L���XN��5aĕ�!߾���s�`��߾�}�}��o���ns�L$��������̓��\d�O�?�!P�'�,�}�!�&�����M��%J�f}z²|�@�b��O�=�k6��gs�ט��Ym�**���~�(�C"A'�u�2y�'8�'.��Ƨ��zb,/l�l�u���l��� �v{�H`���G�vZo�i�s{��va�VK�vU��%k߯>��zI6V[ۃZo��+�,#�J��g,5��e+��~�?|s��N<I4���RW�4�{�d�+��a�I�6a'PRw؂�Y>Ag}H)?$﵉���;�o2a+	�S��'��>|c>�~��uǎ��&Y?$�����:�N�N����y�(nox�$�Xg|��I\�I����AC��JÞ������ߍ�_e��e\9����9˷���S����L9I>|}dRu����08����:�`3M��4��?r��2��5ϱ��+}�Ad�2~�2u+!���~a�O�����ny���;oҸ��؜�����߾<�����~Y����e6rȤ�큛C��?>O�l4ì&CT�e��:��n��d��w�O�y�yO �����ٯ������~���������^?2e+!�|�~a�O��o���8ɮ{|ԓ���	�)�E&��2����iS:����5M�):�����hy��>���c���^k�}����ƽ	��C�>��i$������'R��N�y�n�p�ql�$�ﷂM�|}���I���d6ϙ4�1gY&ҦMXu$�z��z�"w�}��p�y존�A@��'P�'R�Fw��I�51�f�N�姙:�a8w���q�&}d��q��$����Jɔ���C�2�����N���������w^�a4�g�8��a�d�+��N0�'R�S��N���{�I�/py���O��@�M�I��Ğ`|����w�0ì���߽�v�o������o~���\�C�Y2���)��'SF)���y�� ��s��q+3�'y�����B�u��ﬓ�?�$�ԓ��q�6��y�q�������8~߸}�~���0�>N~�$�:�(|ʓ����2u*V�:���2�qы�q+�d�'��}߱!Y:�'c�&RzϽ1ﳝ�׵�>����fD�	�~qxK�Y!�b��;�^7�"�a_wг�����ȥoc��.�z{��u���EJ�ubف��.+��8���il��-܊.[�V���R�'�SG�bJ.�Ҝ,��e�y�D��������~�tN��e�,�K�Y?�}UL�5ޯ~l��R��Y����	�m��=���������PP����T�AH�8�̞M�$�N�uC��	�k<���C\��I�hL�~��m{�쀬t����6~����W����ē)4gؓ��O�2����O��Ms��0�y���PP�9gP��Jɐ��>d�k�q'�&�9l�����uCs�)�������7�W��A|x�1:��M�Cg��06�]�8��l8���bO&�8�/�߰�i�^�삒uO{y���39|��q+&f-UA�p����������z_o~������m�-�m��$�����$��;�i'�'=�,�a��}�y�I�~=��d�5�XO$��쒲��3ut_�����G��k���_�+�}�Ri��N�M��2|��˴��o�$��L��XJ�!���2N~��2����{�u'�,��`'�������`.�����U?R����W��u�w���&�dY>t���@�&ܦ0<�?PӴ��h?X�̚a��I+*�a�	���i��)(W�_��]��_��!9��������J���Ă�l�;��4�<���o2c��{��$Y8�@ɋ�8����!���|ɦI��i�O0�>�~: ����Ɠ�	[�=�K�y�eTIS]��O�R�I�M�a��`���L�����0ɩ��2]�'��Ri���l<��O���hi'XL�L�y�R<yO߽���L��7�~���q&�_o�$�0��py��5��y'YY{x��u��?w��O�4{y�$�&�����	&SS��O���ì&���G>��~�KE�����C�~���^�O)��'Y4~�m�y�w�O�y����L�l���:��j~��y���6k�h$��o<a>`}�}����*�V�5��O�C�2��wӪ�\�zv�(^�Pe�B��;pU`�D���D�;��q���#_��N�O7��
�~W��9JuFeg���}SB�%yR���di�x8/l������>ܕ��/Js�����ɯ֠��W~G�}�v?p��w���hmI�qC�'YS:��0��2y�s�hu��S��a����'�~���d�������d��M���<º��~�E���8)�7��J$�ƿ}_u�T�I��a�CCi�N�X��'��VAI13�̞A@��É:�ԩ߬'Xy�1�x�<���`�'�~����o��VO�;������>����̟�{y�ğ?����L$�CVÉY8�hkCl�N���|��:��q�ՇRy����É:�ԩ��
���gN�����x�����L���>I׬'��b�y&�2~�1'XN�X��ɆHj�|�������'Y���I�M��e�q�,:����U����E�����'r�T����ܿ�ObB�q��?0�d����N=a?Os��|ɣ�~�0�|��Y�8�)�+'Xn�C�O&�I�gu��y�\^�����/k��Uh��?U���9��h=�:��h{��!�o��d�}��=d�&��Bu4ɩ�o$�	�4o�̕	��:�d��G�w�r���������[8�UQ��2q<`�O�u�P�Y'L>d��!���u��6���>`y{�8�&�qf��<�d���^�'��;���y��Ow;���������%ABx��J���3�|���	�O��<�I�٫�Wl��Y�$���>a9��O2i��?�$�i��/�kk��ݴ���?l�߳�z�~��EV����dI�4}��J�$�/�T�edɊO2|��.��N�|��6��3�I]���N��<ü��y$��oƯ��=���:�ϋ�_���m�R����e��h9��2j{:ɦI����J�$�ש+'?X���'̞r�	�g�v�u��P�J��
��ޱ���B
c�k붐ݡn[��f*��.�GfU�֧Q|�4�mD	9��ۓE!7]���v�֜M�3w;��:�	(�c�7l�ű��V���\4EV��Y3�^��=��mZ>���h*OZt���<���>Ʌg�9��P'���m9o���[��	�o��5��������IR����I�	����N��;��m�s� ��&a�~ɦI����L?�'�s,��`d�'Y8����:��c;ӧ2����{���߾�9��>x��$�l�Y8���d���<��*fs�<������I�*�=�
O�7�`�	�O���%v�=���I����;~T�ꕛ�����x���ª�W���f�|�c4�:ɦI���'�_��	6�����$��wx<�ԨN���:�l�|{���O�>��ē_�v?]שZO��N%���{W�u��>�I��%��	�u�!��Bl�6̲y��m��0���w�O�u��&Y'�}��:�	���?$�'�R{q��5^w�t=O�ݯ��R��_�~���0�0?��'0�M~�)?<d�hŞd�J��P�N�3��2��ƠC̞Ay��'u�:�d�f/|�鯿{}��{���L�0��w�<�ߩ3��&�m�s�d����	�I�~�	��'�X���l��P�$���d�'�IԞeL�~��=������t�&��w �?�_e�����ge;�T���Y:���O$��N���<�ğ?���l��VL0�1d?&Y:�+$�&���$��z���y�t߹��\ǃl�J���&�q'SGw�
����<I<���by']����:��Nwؓ�'�F=�2a'�
2�|����<�Y:��v��Ǳ�ߵ�y���w�L�Hu<fé�I�P�'�7���<����;�$+'Xw�<��e'��by'���q�$��'��7�a�q4{�̕'�~w�|ݍ��s���o�~����VL���l�y���S'�8�a��$�P�'2�:��O~�߬�d�w�>x�e�F{��>x�i4��I��&No׿��h��{J�lymD雑*���Y�̩��g�.z�d�J��^X�՝ h�oc���E��������8{rͶ�(��¤�����
.��{"۫(�[�;c���7݃�� �ݛ[���eo\���'i�]��s�������c8λ�t��w;��d�g��Y%ABd��B�q�m�>I�j`��I��Շ,'YP��Ι�1��'Rm�;���=�ǩ&Y32~�l�����C����������_ն���,�=��I�5�o$�(L���VN%d�(I�N3X,'Y<�Շ�u����&ݲZu�䟞!�����]g�2g���޿���C�����i&�?s�'��N0��;�<��4{?�$����*V')���Y3�R|���Fl'Y>O�<��v�v㿵�݋:u%��wOZ�~��+����i���T��Og�d��L2y&�;�
�6�Ν�$<�̚�d�4^�̕*I����H1d�'̞�?cm���A��8c�ds���𿾗��>7믾�t~aԕ�&X|�:�*V�0u��'z�e'PR���Y6�ϧ}�
M��w߳4�y'o�I��'������vs���g[��ύ��|E��bɦN$��?f�����4�$�����&����2J��w�Ad����y'PR���Y?%a�=�
M����^���Q_��+W7G1��w��>�����Y����>dR|��08������3M��4��8���2y�>ǘO��4}�Ad�3��<�Ԩ��?w����_�7<s��<f)��.������JԅL��q}~]0{T��t��lw[����d�M^����X�q��Ǐu�oWOqS}�=�m���n�U��G��~���s�_�<�(��>�U���R~��5�2Ƿ��W��<Xms^�,����T�7Gƹ|��(�_ �e�]�}WO6Y�\)-؎>ň��;�XGS���tټҳ\�뇈j�z�X/��(��D`�>˶���s
��k�r�E&4��t�|���Xzh�P.#Ot)�z�p݃���M��W�O_
*#��h����U�pתֵ�	�+�(
F�m�o;jQt�"@ɔjsc�T�n�dĻD�4�fk�.�Z�k�����������˔bkJ��=n�f�mp�>*��a��0nl<Ú��n���5����d� ��ָ�>y˥=�Na��B��I+�;�Y¨}����h[�0�$�8@����Z������"�mFM���k����"G(e�`��%�YN֍|J���}K*��xY�ܳT���r�Fo��7�v+�b��]Qb}p��_\f��ֽ�#F��N�f�'V ¬x�`��L�D�)�L�|��ݓC2��8��J���h��7�����i���
�N�(n�;ʉ!MިoD�z��S��6!�`�2�XX��91��H�4�֪D���r���9LhfN��X�V]���::���1��L�p1�Z�w��6�[;��Y����&��\�l���u���F�w,@k9}���5ftW��,o���Ӈ���#{�Wb�B&۩���s��v��p�Q"1�h孝v��zm��幨47���n�,Uo��F滗��V�r��Q�R8�n����S�[��Oϴr�^t��8���Sx�1Pߑ0H⑆��b�����o���&ͽ��us�6,���AQ:Gu���]��K�څ� 봾,�U����i��=���_.�W��(>��^�7t��Q�Ѭ��fo2��n:����Wf�n�l��ڌbC5)U�B�"�����)n��+�Y�+��Mv�\U��2n�6KG(݁���z�3������+�v���f6d���2!���2#Q��PA�ι���U��SJ��_Kb�S��Z�3{�1��V��9V�/�{#� �h)U�t�K�F��r������c�r)0U�Jh�k���yφΈ�Oi{��g�#��K[-,b+5Ք+0��	��]�N^諧b�{|��A%/sׇ�A���L��V�h��bF��a[}��><�JR�>����	�DY��(J{ �1�k�:Ќ!<��qsCh�=/n�;�M��G��Opl���E!�ߏ�*��KwW[[Ș�:�Ӄ@ԕ*2j�����}��\�C�)��Z/^�C�t.S��]�U��}��Ҙ��Ҩ�n��2>�Z�WB��c�u}����v�z�dҗvJ�PEKUm��Ur�+�h:ؒ��.*"�����ٸ�Н1Gz�gz�s�#n�wj�^�A���P�g2���Ն��Nk��t;E���gP��^�Q�����A��X�Uqﯶ�ކ!l�{]���U�UX�������TU-*[*��,EADk(�+��F��`��h��U`�V4�"�b-J���1F
(*%�TEQV(*"���%jŭcm���K,V*J
(�#E��ZV**�V$X���*ZUUb���ƪ)Q(�*
�,QRҌQ�h�X�AEQb����b�(1�m�*��ĭF*��U�V
2"��T[ecUAT���֢��TX�)Z��,A�*�k*�*���E�DUU@J�DDUUQ�J!kh��+b��UDU
Z���iX����eVAQ����EQUb�"�����"���E��B�eVE�,-+#h�D����c,m,V�QUb "*�eaj��V
)+(����EX�����X�ETTb*T,X�b�*�

*�PDPYYYF,A�UlTEDEE��b�Z)1AEe�m���"�ʩ
��PX��QNC������gZ����)s�]�6���]s��뾳;mcG��w�8��ty\�ŭ+]�����!;ӭ���l�c��g�U}_}���t/��_ƼŁ�ޣ�)��==��=��=�=뒖;�"έ3���o��wN))���	��sc��_:S�:�h~�'����xw�JX����W9��p��A����G�zɳ���O0�V��{�l�����}��ů�B!ê�kD�0���u���M�(-û�Գ\��į%�[�0H�Gv�Ы����lF��/�v2�B�&�ռ|��֊�;�z�w�W���X;6�9����� �:_��!�#ݪ�U,>�����~^{�9�G���S��o��Ԥ]y�Ȕ����º�i�"t����ԚZX춴l\={�oz��y�Ϝ��*)�R�w�����%-c��TL��}w��U��(�����]��[^�����t=E]c�Q\�R�֟�Gpz���kb=����ry���U�p]\����9vs�k�wZ�E�@݋#'�^�W�A�w �V�Kr�g��sN"�"L�ҽ(�<�MG^~�6P�]vquY0+c�46��}H*��*���c�o8��YE���ꘔ���q�!�<��gv�{�Z,ZC�L�Ĺt���U_UW��zw����9_�.����?p@�Ԩs�Ь���y�23���v���~���ƥ|'��V9��6�>�=2���4s�{��*S) �Y��rw�{����y�Qt��~[��y����c6��?J�R �N��5�׎S����z��z1a{%�#���J�:s�|.{lN����K��ӼT�{d��Z�˹�4��𿓗K�Ҭ�_���fV��>�s�F��/:�]�o�2�fg�7� �;<��;%vsa�EΉS�/�|�Y�f���O.��M�);r������>��'b�\���7�z�1�QJ����sɢ{�6��1PѿM`k0�Kv�Ӓ�����zi;�T�|y��9�~y�|�������u=G�����{��s-�]��=�����/Q}�#��;���j�n�/S�*��ע>��ڱ����Y++�*�.A���Ԇ�V��z�D����Р��"���֎���m�*�I�0�l^pu
e�`a*�qS�h�K��.��\��	���^����kv*�.�,�������W�˺� 2�c�o�UUU}UW�ͳ����H����yl�������<�}��湎oK+�f-��ŷɰ�?z�u:�3]�&�T�׵���&j�'�{W��v�����-��n+�Tv�K�u�`,�vj�ؾ�5|�{����lr͏�'����Ϻ�URMRҙA��;�{o����{�V&蛪���o:����J��ΐ����'	��|<����v|x�y��y���>kܽ�'�/=�Y�����\�]s���z2�V�ޘ���=/����yL���p�u��6��/;���V��oх�z2?n�!b�Fz�.�z���Z�V�~|�j�y1��t���`����ął��{J\��jݚ���پS}��VD���/���t��Q�=�������J�m����}�����g���j�ɹ�=cU��C��oP���^2��6\��ov��N4�ӥ
EX����4kQ�q�m{\,��T��ӽ�E(w/ʜ��w�w<W�]Hv���wG�GQ}���YF�Lm ;l������In;VF�=Q��i��|�f�T��CC\b�u]�v3s.Z�a�A�o��Qɤ� ���\^���)���=�E�3���)�5ܛKk���:������J�#~kďR�vp��<}��~ʚ��|f���O�6��ק�oi���ބ�KT��:X�{&�S;S�rt��9��NF��>�~��w{���{�>J�����Tgb�c��oZ������DF(04��w5��W��O^hU�V�k����;1qo�Ϡ���+`���8��8R��bp��Sʽ�/+��u�ʣ5����^��%�;��Ɋӑj�틻r ��d��P����^|�%R�<)���_�nV��z��g����G��p�}:��p���{Iɪ��E�x��H5 ��X����Q���˓/��+n��T�}��<4	��v_3Kv���]��]t󓟒�赱l��2��W��̉W� �:�qҧ)��R�SR�Y��.����n�޾�oXS(ybd;
Xw/^���V�š��P��)���X𜾹z���N���\vj�h������uͅg���g��'�u�N����͂�� �<a
��Y'qAGa�x���!/mEqiO�W�}_}�.�^~l�O=T�l:<�>uR�ʡ�Q�b��#�y_S�����V��`s���Tz�t��U&yٯu<�^8_u�O�j�I�*�k�*�w�ڗ邦���~�cmr������adǺ�ac��+V!��}�~�gU����x�=���&�����Q�M��fs�,�n�y6k���=�fJ��b�����>�Z7ٽ�8s��@B���u?���ߙ��q��R��*߽F���Q�7���f�bܣ��p)G\Ÿ́����Ҝ��C�\ì,ƃ�{���)�w{d�P��:�?S3���\!����J��ꃮtW��&�{B\N����ʝ�ʤB!þ�~�y��_*/�>�f�SҀ���;��O0�˂�wm.����6��ö=.���)�Ps�ڋ�tþOS�ofr?V�k��!$]���*�y��K��^�U�,���6`?W��5�ض$l\q?]�����s����|�t�6��s܂�Õv�H�Ĉ>�y��bӷ{��p�	�Jh���~�g_�����c��<n�.�Mo
�r�K1Z�!�kʩtF뫒��2r�!�Ԩ�̋_��Q������r��%8���}�}�}UY�_�������)���yW��w�o�oR�u��2%�K�r`�_��|�a�m�b���gKW�c�^��w��77��*)�x(jy�
L���J]��V���K�����<���ޕ�#�y
���kպL��{v{^��u|���ER��kd�\wة.��σ�ės%_���ջ��Vg�R���Uҽt�)���R��
5�s���:�c�O�E�>�s������+\�u�:T�=]�P�f����ݟA��s�'��V{Ф9N>�Dz��>����N�e,�mF��|�o˽׿yvk�����߹�2%�qPڭ�ײ����m�������^2�G]~ƟE�8ì�v����tV��G����(���.n�W�V��U�:���X�y�q_���R����2gR�W��<��^7씛�/3�4�a��E�N�씆9*���=b)ꫵP�Q!{���GS0-pұm�%\Cͷ3؁�~9-��DW
3w嬬N���k�*"��KљPOf���+�8X2��X��7~g��\�:�w�k&��u)��̓���J ��rc5�wl#�Џ&�}<��dy-���Lyw� >  ���ֽS�I�֙���ތ�g!�W.-�Y;�򁫝W�)�����*E��J�u���M�9�f�7������.�z\�o������x��6��s��9������.�����^��/��-��8�qz���5��m�9pnd��Os�7^.�Ɣ�7MetёZo����ȫ�Q�����~>B�E{޶d���z��s��_u�7�����v�}�q爛�+^�z���S��`��_T_^אݝ�����{pq���Y�d��^��]���)�/)���U�pz�osü����VhVc���>������+RA/'���{�ڒz�����k�����h^��v`�M�lD�Y��:y�n��{���;��r���^�sc
��W`���F�':k��b�Ne�_fѻ�K�
���ys���5����Cҳ\Uw������m���@K��PZ8��6��{{҉Q�a�P
��~Rl���[�r�-�V�]�]�Ƣ�;��V��wh��O<{�-Rnk|��J0�U팤k|��\�.�c{���Y����M2gP4��/�뫛)��}o�}��UUU�ܔ�]Oͧx�l�W!F��z�auݾ�����0��=�E�S��0�1΋�؞����ƭf�+/��缅�w`��/��_�Mz2�9w��=�o�I���ͯs��'���6�ћ�W��+j�����9��6פ����5���s4�ލo�fy�zƣ�W�Ru4�nx/=�S�չ�%=p9sj�G�q�~�'n}o�|
��-�3�A��W��Ol�mi��U�5m�Όu?	qΘ�~Ϧ��Ϝ��%�!(�v�;S��uK'�����,q�*��o&��9�N��g���r��>y�����_������Ӱy��f}OCy�f�q�aҷ�:���r�3o��v9���]���`�/���ي���el�amiU<<�N��T�u��e�LԾ���¯��Q{»ʶ_V���z{���y�늟<Yyu�b����v���-O0�u9%n��F�%o�Q�"��?�󻗥վ�vR9�p�ZB�S�h�b��(%�)�t ���S��*�y��ٽ3�':o�te����KQ�w X���[Y(ua:��徜�0S�#ٸ���cC� �s���|>����^nI�1���Z��z������߹`����t�֧fPV�3�CR�o��zxl�bZc׻ۯ��#ʆ��8/i|�������7J��^�ر�i?v�}6��P3�H��ߏ����]Α�6�|�=��{V�f'^��F`f�S�Ԥ��b�-{�P�P��=>'۴������u	�����$ߓ�C┫`T���m�S}�a�_�Զ��yu��맯+x�h��c���>^��+�����r��OMxE4_��`VE�HnطO�j��<.�'<i�Ln�_�Sۜl���z{�ꓡ�z��I������&Lܶ7z��/�sU���͟fu�0��YS��@=~ؚnT<�X���U㢥]t'�U��Y+#R���qP���`yP۲���Ҷ�d�����2�UV4���#�DO�������>�'��;�ӦC�/��Yn{;��ڷ��:��f)n�˔	̄ɪ
E�ʞ�ۧa�!�`nx��2 %���*ٹ�v����O]Ё�-���Fp\t^.iQ�fy��r��)�/Fʋ��9�F����e��/w%��oCE��Ûl��˽�798V�� ]7�WV��=N�t��� q��ŷ���iG���La*��K��꯫����>^�ݎ}���̔�v����Ua�+Q抬�%(pX��`�ꝄO#j:~��0�̏�󮖳)���=��sz��D�Q�}A$W2�Q*�k���n@�2fT�n+���h߽�Ϲ�OsHr�[�)�ll�V8w�� %��
�����j}6�)L᷺�On�u�L��O���O2�kt�'���~���r��PlVhk�Y>�ׇz���m������=��V�doy[K�k[-:�1��>˰�Yػu�X�T�;���R=��~l�~�o��������v���ZX���.�܇Yb��9N�!�e�GFd~W��.���]*�l�N���].Z<���k�0�Y��]�#Ӕ�]d5�gIB���t�{3R��@����X�UD��0�צ��/�{N8�x�2͊e���l�"�;�r�{x�i^Q375�Xt��'e��f ϝ��S+�w�U�"x�GZ����YYO8����������F��U��J�=U�2Pʇr�`�z���?x+�~5�d3__�n�[�A�]��&Gv5���׭�T��x�Z�*�V�ٱa���mh��/�٠LHcQ�W�h\�v0��÷\3O�q�WÀ��Ud��t[�7W��w�󓥛>��|M�h�҅=�ӑ�3OaƩ���Wa�Oi�4�1�w���n�j�k�v06��g�(m�
�(�R�+OKg`�]q�\Ǵ#N٩�x�*�R���I|S�����R��Fփ'vvv
k)��,	f*������w�m$/��z�\혻�K��'k���"$�告�#��r;V-'�.�����eZ]tb�|����֠յ�ͻg�Nt�،��yz���k��tq���.��d�*�v��Ծҩ�Xr�K��(���P�Fg����~M��ȫeǭ�6�as���0�(���NK+V�'xQ0k���:��
()�����|����1Pɛ|'VN���%P9��r��i��zf��r��K��s8���4F�(��&������dД��Z�qQ�W�KX���޻�ntF��۲�;݁�`�3�������&��ta�Z����à[�����91L ��;��VoS��o%32�sl�/|�rƺ�N����]���
MՔ~r����4��]y�{'x"��R��7����q�9-�n^�v������с��m��Ŷ� Ia����P�����5�r���ܠ���,
�j�1�Dv�����`e[�3�֌��J���d�+l�z��,qd<ZpJ�e3�f�&�⥠�x;�"�%�2��]��Q���!۪�{��::�ʏŷ>�[1]�~���e�m����/<(���{B�Y��!�^�YFQU�q��PwZ�Y��1˄�cz �WK�Q�}�L�|��.弃wU|�K5ö�vT�T�sj>I];&�M�t��a�7�׭>�/p���^T�tJ��J�YwE�����!ݪ@���j'q��N����l֫�0G�W�\*gJ��0q��,�������DuEV�P��7�;���ڍܙt�I�a��rl�Kו���nn�7�7�-�TZ��E1r�9�~��Ò�)@���`�du�ۙK�^G���A�k�rȜ�n�g��W�h��X=T5ӏ2��KX��N8�U�Y%��//k���u�t`��W�Y�c�h�N���&�돥w:���Q�@C۰�B�P���ss+�G�dz;��-L�o��|�U�ҵ��>���i�Ώ.���Ķ����v�;s�IZ��GQl6�,4-�|����ne���`PR�j��Rn�_'8)�Y8nn�x���������aD=��7�}�CFK�@���5W�Wq�d]٠B�i�i�
nVd�:�*�ÛY=��*��3i�C�v�e
J�^7�@fҨU��F�<���te���(�m�\nT�Hp�����ْ����M�ƀ�E��&WZd=/��=+;	�z�q'�v���M�kxV+6���}�.b��Ep�*�
EU���P�TD"Ȉ"T���A�
�JʫZ�D��QAQ�1b���[D��Kh��QE
��ac ���[I�,+U��ȫQ��J��Dhւ��E)Z��`1QE��A
R����l�-)
�E���V�b��T���DT@�b��ZUTU�l�mQjQ%j*�����AB�V�EUVҬ)E��EH�*�VX����,��l��%���YQ�	YX"��"(1
�EEUb���VJ�F*� �E�1��""�-�E�DAF+U�eQTA�U"�TR(���R*�dX���"���`�,Z�aH�������cH�ED((���H�,��X"(���QQb��QV*��+UE����[���Z*"��U��Ȳ���Ȉ��Q�(�R*�D��PX��`
�,�(#PA����AdQb���ȳH���"[В�\͙�g�L,X�ڠ^����3f�䷶�N��􎤕uH�!��n��3�Ћ����1��S�}��W�U�z�~߇o]�����շ��O�EoJ�ͯ9���~�����н� JN����\�=87¨��y[��l��עB/o�����F/w�1�^쎙�ŕV�V�z�{ޔ�L��g�>�{�ȡ�<)#x��HVu��{K����&U��<̩�nW�ϼk�����fe^���׹.ޥ7գ'����vȨC>�(-�±�P� �|1gh�ޞJI�v������̺��y=/@ξ��{u0e)[�%�{(:�*o�y9J�g۵8�u_V��p00^�/��peS���N��*v0��n&/j�z��#�ɞ���G�I���7ہ�Wb�]�
p�{e����C*����1]Sp��{�|u�N�>��d�Κ��(	U���4�&��u����5�/�{��b�����4i��}��/C�ķeLֻH����4 d�Zbu3���P��N���R��.�Hy�6ț�������^O���aϪ`#��P����$���)��z�h��_���ҡw4bB	{�ֹX>T`G՜oǝ�r��{�m��4�J�"X�Lf3^��!�wO2E^���˕]����w��_U˕�Osi@Zlp��o��{��ҳ�e�_q�V�b�oF-�g+�Sݽ@��;;)����t0g�G랊�����t��췚;����!\F<PnT^�� �苣a��!��*}�=��W��绂i{z3廄�d�S���̤���Ahu �����^�B��vVXخ�f�� �w�qj��e�S<k�c	�yD�T��ET���|�z��<6Fw�~3��*��}R�꽏sd�+r,�*ƣҕ�ٛ�O����V�J��:	��:OB4��d�Syu�~�K���"y~��~�]�7����]b3�,�#�8,y�پ���KA\d�+��h/{_�C�b���Æmg�ۇJ��J2놋g�&C�{mX�x6��Ӫ^vJw$z���X��t�2�ޱ�}�E����^���U��q	A4�����Fx�->�.I1�g*������3Ӟ�A[����Nz&�.���}��F��*b����	�I3g���A�6�cg�	N6s2�ߋ�5�&A��g�>��������M�	7�<3;l���W�v�\ `��<��*��jc1=>��-���!��ag[��������V�sn�����(��&gi�%Y�%�˴���e�5V��	�wӍ�[7k7y�ap���)'2���}*��]t�F�
T��	��p�U״L��9��^dd�o��2VА��R�T�C����%I�mqJTRvs�UU�}�zM�.�9�P�� ~Ǜ|p���A�]�H^wO�)���ӽK�ҽ�If>�yW��ɷ�L�^��lҪd�*�0�����<�+h�k=���u־z/���*A�>ޏ�b�kNu�»ݖ'�ʹ����1¶��֩V�Y��Y#�b�YT�}���>j���]k���9��S�z���~ @��� �� _�F��+�$���nY빌NՓu�NsONK�{U-p��Ct�r�[�����/R���y=�ҬoY��@�V��N��v��ʡPL�t���Ѣ�~��2���J�c�Q��N2���}���t���;v@���I�4jx���+)N�x?V\;x2�Z$����t7�r�����d��"�:q~nR��1M}�� �+�E��xf�$�]"�X�"*��Nq�۬Q�Q^xh�Ғ��v�Q=UyK���u޷)M�E��u(���-���b���h�ڶ��Wz�^���X�f5�U�o��L/I��0)_�JBWv��>'�߮��5u���5����
'����pz_e4�Uͽ�۹}�,�l��b�˭�_��I掅�-�b��
��[޹+~�j��j�˶��+%J۠��9ٸ�[����iV'DR�,r���XsܣY����'K�U�b�ٶ�����,��nc���磌ꯪqo#^�^.�W������yW�bP��q2ro��ppѾ:�e�A��][�ب�/�o-��"x>R��۸+>��Z���0z�L���:2m�~=�h{
v�;5izj�>�Z �����ac@].�Ͻz _��ʾk)��b�`����o8<�UB�Ҷ�^�h�T�Lp��&�Cp���L����ͱ'֊'!��j���'r�Ö�Თ�ϸ�^�=��De|ɏ�P�˾�V;d�`�݄k�r��5��95)�퐥f���s��N7�?]���H�Q�}A��\��D���s��W�F����gI�:�v����x�|������S��8f��B�	;�I3�#�}�)2&�*5�=C�*o���9]wztw�<B႕ī��=*���K��joQG=���{�h�<�T�EJ�Hu������-V0\��}��]�*�=gW�H�)�(�y�mw���m-r��ԧnᠾ��d��_�(;ƀ~W��-,M��^P?B�p�����|�����XN�M/�ŏ��F���Ds���gϼ�Y>�	�_.aDG^�n�5�{�,�
�e��At-�"�[�3� �����)���>�ӫ�ofɏC֕ѭk7�R�����=I�|���o}U��}�.�Jqdm��#�?W��R�yJ�<�MkI,��¼xOn�戂�ܭ�:��K+��bx�b:x��t���v*^ �gU������I��T8�W����|����Ԟ�.�����Xt6��zNt@h�؃����]c�j����D���T�J&��\���Z��=��i�in�ZN}��Q�P�p1�+��l�e��
��!�Xܱ"����E���:;����,Ԡ�}fP�ע��ҕy�L���t�<<%��W �+�J��~���WG�����5��j�;��L��萌���	ج�s��Ȗ��5�5���C�ɔ3R��8���٣l�!.�hu���Tfht3�m�N-LN�η,s{���{d8}̾>�T�^����)��8��5�F�fЂ�z�T�l�0�3���a��xa�[qw8�̺�+鼞�R��jo�@,{n��f�gu���K��/M��1ee'�c��pïp�)θ:�������90ë�*�=g���3¶JN�On1�#kV��p��`��sܔ�R���Sǖ�F �iAq���r�4��+r��p�g�����r����ܶ%���3sE��0Ou���1�{D��f1����+��JR+��pgv8
�m�[
�Y/��?���UWމ��I�"Ǹ�p?��T&p>�N�l���� �˩����#iܱ!}����O<�4�E�Z�h�FY�áϮ�cH<���K��?
���N�d�dH�i�p(�&M�7�f��+%�Qzf
��z�g�ګ�b,�LY|+�W[Oǵ��?3SƐ
���"�Wy�)h�w��2�|}�
�u��B�}I�a��e=����:Κ���w��&�������v�ܕ[kGg��ã�#+��x�܋��WK<
�4�ϒ���	�O0�0��c�c��K�H�69��V#Y�?S)>>��� ��f=E�D/���1��S]�n-a+�Y�o�8��^g^��yU��/3veUSwt#��K�C������C鏳T���g��wڀ���n5��Rd��X���"O���T�'/��!�	���e�vvFڊ�=Ylz�D嚿 �v���*U�ҵ�x]n'�z��� �.�V�\�r��H7w^Mo;
���5&����|Pt3ǌ��JeP�Y��{mL��L�����K<��)o]n�YYr��v�ɳ]��i�+��-�4��J7�~�k��i(�2��]r=��ܔ�H?5H���^�~�Or��K_R���җY�*o˯�٩��d�z��O�b�Ƥ�/L/��75����W��r�����}Y�t��6��Q�(z���,���i��ݎ���N����֡e�ۊ��T�o�׷ �3�P)rݩJ;���6z���m_'���3Ӟ�A[��c0�`ǅ1d�>�86���S^u�v���f�'��b�a|x����a9� �oň��P}����g|9V���{7�n�~ȥ�/�^�gK���]p ��zL=P�51���N+Y����]�m�Ե�Y��qyBG���U���7��(�yw#��õOl���z���塎���=��9瘆%u=��z�Q�T򾖅@��OP�����y��B�,0��Nοgkhgv��>]�d������<2�3��WO�a,T��"f��r��ve*Įϟ�N���#��훞lͶ�ײ��T��R)��O.�N� �zx ��R���yz'��u��5�~}����A��{�>j_V�+hI����L<�(��(0OA�0���ݛ�N��2�n/nGf��^�X��pu΢Ӊ|41�/�Mze?}
U�)�(�9u4���at٢�P'=�V�nV�*=�Zn�9��q�tS��s�[v�L`s(Q5"�o��7�l>&�3�d��V*�y�֞�<;��a!M'��]�r=��_�F���yT�T�*?kڡ�<���L~��H6����$7�+����u!��������m�;��w|�i`��d�^�#l�墑<4!3�y�%���
N�[�} �6�	��{'��;��U��2�߫�&�/�=�`�E��xf�RLU��Xʡ�"��?	i:SC���hex�v���z�`yW����)UO�VN�a?�n-#� O��.��~�����onV �ݸ�>�μ�{����F��Z�^q�BazD�]�^,�Y��l��e��/p�O w;8���yi��U;v���z=X��;L�r�3�|7]�Â�|_M��De��w�c��y���^��g�pBr[�w½[B�aÁ>����0���;��=\:�x��]��'�K�r�~�tz�a<���C)j�]O0=^��D *�_�|�S�1M2h���-��b�Iw�=�顁�vˋy�f�뮳
��̸�.��p��c&T�ZjxV��ee�7ݲ�Ûy���8�5s��׸���=�ϋ�=WA�,"��]W-���0�l	��$sKپ�{�Ūl��5<�D�LM�m���O�D�� �O�+�;K�^\�H�[�5N��f7��u{h;��Z�c����1�a�Z��ӒV_�9��������Ǚ��z7;��s����j�{峝�[nD�Ç;^�;ra�
��ʴ�{�R-Gc�)��c���j[H^��p�#�׼e\vB>�?�U}U��س�����U�į�퉾��a*��\5�\���e�U�S�Y��X�f�<ߺ���cD�F������Rߎ��i�l�X�2�/�
�ə[�9�P^�i�лg���ٹ�Ew��x�JS�(+t�������5��י�����˰�V�6�;'��;�;�E���2��J�WM�A9d2U\�]��hgI�ե��~k�ik83 <m�7���/ZCt����\��)נ�d�y�i-r��)�uja�*�[\X�Fl�/+Xm�9�꛺��U+�c6�$���v*�x��W�*���&����=�og�̏�=��*�{�(��
�r��9�`c>��	�k�F������ܳnP�/G��R<<��y�}U�Q��i;ή�8�	4�@xn�vX��e��}�kↅdo�y�/}�o���R�m�0uf��m�2�>���*�Sٌ�^x� �o���phmi~iO73�\�=����Ǩ�j��G��L��¸�����"S�cҫ�ثM��m����	���_�<�*��_>�6�p�|�oY�>�K�u�Ϛ�.si<��#m�&z���A����T�3#��J��W:�2�����>O�0�k��)�����	�t��R��хP��[�0W�яW%���gCX55���꯫�2t�m��o�5�mv��/x��ޜ�Z�VtSeS~�sSB�Kq�`6����D�m���}���.���jn��9uF��=[�f�O��"�A�AC�x�3�_	��&E��OŎ'Ã�mN0y�U�7���U�@�Խ����<�%��JA�̕.���+�^��le�@�ӦO�����	�p�w3�/�nN�˞*{�1�2����׽5�b�Y��)%����'���x_�e���C>fg*��)y��;Zs+�z4���wj<�Ab�	���i�]�a��[Nm�C\"��r��}��9�F����~6�C����U:�y�Bh�fN�,V��L�+��P��N���R�2�#�I�������wp�ӃD�38/dOU	�j*�T(�Y>�/R�'���{L�e�/�<�n{f}���ީkG0b>#+��x��x�cj *륞UY�yeI��i݈�����<���e.��������)N2ck�j��0A��"6��&��b��Q�5��ԇ3�A��D��=��E®��[#�I����mGh�Zv������Z2ٜ8جwW�6��͖�Qs[ס�k�����rRU��:.<����"��������������h={�+����P�V�L̤���޾�9���+;�0����:'�Fs���XR���8�k/k��qM��ǰ�g�^�VM�è�5�ՇM>t��-N�Cl���E�!��q�w����m�n���*I]�q[��o~�������o�R�&����\e���h�*��>�'(;׌R��n@��Hl1�S�476�v0*DTW�q��P�Ͷ.�i�LY�\���y��X[��w݉�-�d��aV
�E�z�\mg+��%q��@�=��\�L�Ma�S#�ו/(!E�V�u0��f[����ԩgP������9G��ެ��+���N6��u���b���
Z"1���l<s;W7@Ʊ���B�e��3o�k��`(�E��.�31�eEl! �i>����.��o3�R4:ek�]WX�v&2�a�cn��v���r�����(՜�9\:c�r>*��i�p�^���"leS�����_U�	j�t���ms84�ϕt���;Rye�%�vs�ƪv�A��:��vj�;����������dI����������5e��N5%s�p�C���ݩ�����<��%|+E*�	��8
�O�T��
&Z�I�mQ�>�L������O6��Oo���)Q��������T�3�5�i��vR���"�p⹺K�G���ۊ���g�\�ۖ@ [3��S]��}��]��͝ǠW9vgU��"n�N8��R���	*͜`��wٔ��c�5k&�]+r:[Y(��r�OE�,�n�P��2Qse��s+��P{��ۈ�-����)�[���N|a�6E��
 .[���\��<�6�F;�WSY���u�ŕ��3�0&���npR�� �R�t�V�6r3����_G�y�͑�YU����eM"���`I�wu%!��x�b���c�ވ�,lz���X2��\��-	�k$�za���.u��P;%m!���$1��6ֆr���D�r�.���㏃�9	��I�X�*cŤo����(��
��F6x����[���罶��Q/#YL$Fr����Z�j���5���̺�imX�{�1 ���+b��P�Wi�P� x"=�2�����um5o�(�`K[QN���`�7e�P�Dt[7���������ٲ� ��dܡ� E�Dm���y�I��W�mK9����zr��^c��R����x��v�/�;j��6i��oD�KM��gK��.�\����(��1��_S��nx</��m�h�3�n���ծ�D��D�A]~ij��|�q�>�F(�b��(��"̰��� �1P��X"�������1�kX��D�Y�	Y	QED+
ĭJµ�X
�*֥����b�ő"�((b*Bڢ�)��X*�$YRTQ@,Qd
"�"���1U*���FAm,X�EQ��� �IF6¬dQE"�QV("*�R�PXVE`�,EAFEdX1 X��QUb2(�DX�lmb,P�(+mb�0Q���@m%hʐX*�VE �Z���X(*�YR� �EA@�
V�,F,F#`��`(��XU��TQEb�E�"�EYb�a""E@UPU�@D�+QV"EE"+UTKJ�b�%j�"���H�Ƞ��Em�TҢȠ�����E��DEX,�TX,QQ�dQU�`#"�PDV�UQ� �E�8�q��������.�o�)����,9e����2V1k��vp�&��)C0��K�ɸ|��PC&R,�+�l7-O��y���n{��g���j�9}�ܩ�z���ݙD��wt6���VW� 4<�(�u��>�f���vãح�9yP!�a��:�����`��+\�E8���=^��8��r����7�����x���|d�@^��wJ�V�������c�o��E_�]c���9˸���2j�'�y�_Oc��>5��B}VP�خY����2t��ŀju����jkt���z�(�7(�P��8����<�t��;�x�g����Y��A��fUYw��|��U�^��eY�����[/�_'�����j
�R��t����+��`��J�}�3}n���#��(c!mx\<p}/����ί��_�z�T|}2�;كt�C���-*�ز֏Uf���J��>Ih������<مC8�b[��N5��/>MmH�n��W���`��yJ*0��x���8������D�ć|��ϫ�Ո��f%Ǆs-os���N�V�����=k�4؜U��,U���"�yJ�,e\���r��]�Kzx���1�m]�$���o1I8!�q��/���H3���{EuG>��W�������5��E�W���2�v,��!K	��<��U�2LŃ�~�0`��msz�B��*��ޭ���.�bcBy�ʞ�1��Ғ�H�ͱ���UW�w�܋zF���Eo�h�Sۜ�9�9t�S��vUl�4)+� �� ����=��/�^o�^^�b�2�-���7����Rs�2��x���s��^����.�b>SQ�d���-R���eg�UY�t�\Pkږ�hp^;�0��Od2/R�G��镘�����˰/�`�6�2]v��x|5Y|v�n���ze?T)V�r�;K�:u�}��9�?��&Δ��U��Z2��2K��#lϗ��M.�c����}�Ȓ�i��_����f�媄��"����Ǌ��fTc�d�΋�0��ߒb��W���t��.;�t2ݜr���C��|A����M����K�e��S���Ց�=�i�����^��=z����sW��Uǣ��:2ϣ�4[�P!yǄ`�^���U�|ލ�Y�=�-P�0�V���n�<��_oO��3Y�u�����^��<y��ʛ��v��ÇC�����Þ1n���v^F���|�<0��r�u1�P�Y�]N�ʹ�����%dj㋁>���_���p�cu�W�"����ub��u�����g6l��3�R���il�\!�l��R��]P��홛P��ݍ�m�69w��O�s�;����z�\&ir���1�Gy�5�WQ��;��0x\g3�9������o+�=Ny�Y-�x�~�5���a�S�/L�O^� (K��d�5�5�miSi��f�$́�6w�VH�w�=�C�r���qp8`�����E�LL��A��~����jT+rX�
��=Ηk]C��w=���}Ĳz]�\>�hJ�(�Vk�y�t����1��v���D_O*�3��������a�Q��</� %�V�Ւ���??wZP�%u8{|�i���W��7�;�Os�3�.�����^���4����;�R>T��ğN���
ʕ��6����]o���ӵC�����e)�
�W#1%@c��:�=�wB|��!,����ϐ2��HK���+4����KN�����A�f�1	�U=�;��Ȭ��i��S�7	���Pw� �J�����v�Rz�gd��=�vε��~��k"#���u6�T��F�,�Q1|��ךXΡ��	N
���\�-ܡ�}��7*^;)�d�ޑ�`�UD���.�Q�=V_SY��wz}.5,/pٙ�T�2���k����h��ZV����ջ;��!b[�&�:�.ݽBX=�e�E\�s2�X�7�4�k9g�f��S�{�rJ2D}�Un\4:kq��b���i��<m�HRN2{M��	wմu=�0V��j��R��ūrs������q]��T�7cG�Ơ��ފ̭הO�8luB���r��9���(@�(�cW�vn�
��پ�}�eg���.ţַ�x��E/�݊���WG��(eT8ӕ� ��Ow��	9_��7�vD=ZlU��Ku{n�c~�J	���e�·��[H��ǀ��o���\��oJ����0=L;w��,�z=�4Ъ(gñ_��¬�L��^����_d��PC�m�k���,��b�g����}��3����7X�t.������G|7Q��\[����	��8��3�Q
���I��=}��w�j�
b �2��T]�����=c޶+=��b/���e�	��ב@��o�A�X�4W���\KS��猫��Ҭ���Zv�%.f٩N�5՟L��
����3�z���]E�/Su�E�<�|fW��WE��$��J�&:>'�j0��yu��9�n�!��ۏ��^COO\�+d2GS�:A�����k�m9�h���ݫ6ޫ�d[Y�n����c�']���ޭ2����I9�8e�+ĭ��וX��R�ٗ��*J���2�=*�]��{���}˨wu�ZP�z�X4�`o��[�X�3��skY�G%t�	�����Sz`\G���[��1mY˹۝\���:�;/�����{��f;���jt�-[%�4UT�"����"�BX�1:����(OX��z��Z���{��-Oϱؼ�wJipy/���KB�ᨨ�߽u(U�Ī����(����uޯ:ɻ�7O�vYS��{��h�na����5p{~��P�W]/��M����?=�n�ih�U!U��V;:UwE��7~��sOH-�س0@���a�B�'��ֽ}�'���`dp�L!���2��g�?1[�&C�{�%�V�iϛ��ē��vfm_�偁��bP�)�ь�5�Τ�c��c>�D���V��r�+���6|t�*=^�Me_������pk�',� �e�C��u��g��Uo�]�Vث{:���ԇ+�W�S Rs���>��5�^};p�A��:e�pʫ)�ifS�)�_+*%ޣ�U����2�oڷ��<2͵��,���l/�����*���8���Qgx��C��~�}�8?k��\I��½���<�O����GpW���t���p�[�[�-�'i�x0�듼d����y��^r-�l���v��y ���zx�xӦhr�����g}�oc*Tj����"��C-��\�V*���]V�.��+�9���H[�$W�^���{{r-�i�:�_��yߟ�������ŭj/�w�̻�I�F�K��Xy�s�k����ί5�4���ۃy/�X�)��]jY����n%a����g���u%Q��̎���.��a���Jbǌ��.��!�2�Ta_Q,��YU5�.J���W���J��l|�Ki���#&n�Rʣ�u��=kæ�9]��,U���"�D]�7x3�����N�_
ǶD8!�'9�FmK�����c�fa�H:R�==ѹy����睛���m��x��(5�T���9�.KxT�R��Ww��^W�y����ω���H�%�v, *Ʈ���jmg-ӕ����k���n�K�#����0wh��<�g6}��y�i�}�ŷcn�eR��R�F�J��BxbgPڕ��ĿvS�)V��3��R�{6l=�}��T��ً��޲M��~'����;7^�cYX7e�t�v1.��5gF�_^��l9^)u�dV�T��̨Ǯ��ޣ�Z��yt�
aY่y]�^ٗq�{_�Ŗ(��P�+�*���U5I��E�V�fd�Q�n xs�K
��N��팍�9*��-vv�g(��6� ���os��	��ݗX��ǜ��qwH,�#:�ò�^���d�T�K�_];���*���[ac�|�������'I^���?Y�k�N�2�X~���9�fy�b���"ì��Ek�w�z�HL�./)���Z��Ah��v�U�k������t@U�^��V2�ѹHwN^����q��y�O.���L����1�㨺�^U�q�C�W�L��ln�U�ÀXg��z�D�MI�Һ�!�`"We�A�!x�<0����1�P�gu:V�p9<M+��T[��zf5%A�ޠ����e�C�w��0=�q[ �v;�u�F}�� 
�|5���>ܽ&g�H��&^��/
�£�l��݌�
vH�}�K�AE���$EBک�\��zs�]�>�PR.vT�Ю�C���ջ�=���U�A�d�%\|�����^L^����3�Kbo���E<�D�L:�.o\~��@��}B��1�*�^x"��*<>�b�^fR�|N��g" s����4���'���Z6�|&�q��$����OK0�TѮq4�Wx��v�ztwOs�.u�X���'(;9���gծ���c+h9�$-u��ua�nm�1�&�z]٫1�wA�ι�R�L͠���9{��r���$,�7���Ηer�J�V��9��ZB����Ч���S{/���̶*�t��ք��Ew��й�����5�j��Wj�h�bֻpU����l%��������V]SZ��Y<Kn�f�K.y�)nk���U��sE�T��4$q&�%/�t*kI���S���ԥjܷ�׾a�r�ڼ�~���UK��P��P���T��E���&�Q:�K��w3q�'�ߞ��y����P���eu8T l�ޑ�`�TI
��
�WU��	�m5}��vF�x���jc=���7^Q+ے�B���ʷ���=�c�,�~R�v���\�(�{�N��ţ���L=��i�~s�hj�d�x�".�h�=�;�ޞz:j�٪Į>�1�ô �۴X��J���G���1�k���ZW����z��v�w@�|�>�����=�6�eQ�c����9��p{�ٮ��1�y������n���b��lc�O,��4��n=E�ttS*�^�1�n�J��)��y�R��G�J�m��S*���t�iףS���\���ѕ����q� {��>E�p=���?:���Z��%��9��s�`>�����ą�4���ˏ�>?w'm^m��v��sd@��O�Z���	�����k�1������:n��P~���KeV.BŌ��u-�Ľ�����t���y�Mi��ʎ�pgQ���"���]�ճ�)��,��]~�;�U�2r��1�8��qW�M����E�U)�����>,E��?��g�˓�]o ���E	B��+�C���0��pe;�����8�!G�
;f=���_e�	��Q�<B�`�I<;~��;J:7Bq�95l	���w�)��>��iq:otz����G�D6��2T8F����|q+�d����[R�1�Jwm�*�QC�&�o�M�,���/����]R͎hЖ=لU��%��bu3���P���ԷVtc7U�,����)�;{�dK�����H��+:����( ��&�3K��3M�qe�:9�\.z�<�=��;>RU;Z;��EFoH���7�| ����7]4�)�>G_���e���ٕ���%�*���c�COХ8��Pz�meH�>�|��R��ӕ˶�� ��D�,w��x|e�ݙD�Ϯ��x��xn�.s[	󜩭0?N�Z�3u���3��%��P��X:��e_*x�z̞�ѣ.��� �|0Q� X[o�N��EQ|��(�����d1ӯ���7�/9�U�~��2������u+#0��8�/;$�i�����v�u'5C��r跩�"���N�]F��[�.�����Z�γ3���6�r�N���,J�.TFNvז�|��ܚ��5m_��s�s�㬡��jU����uS�pm?"r�_ � f�.��`ሰ=}R����������Z�t�(��\�
z��9�݅U=�Sύg�І���&/�\������Ӈ��^�C�%��u�#��o���Cc�Ǆg��n�Gz;:k�p���9J���(-�����*I��V�e\T��1K���]T��3�����Nz5o�Qxn�3�����v{��,�[�:����i:�iJ�lg� ��%�8ڝ���)�1�}X�-,$B��f��1�P��OO�/\��J3��Ϫ��L�K� 0pl{fc|���0W���C�\������>�-���TaTO�9Wփ �{J$]�Mг`��N<�O{�Ų�}�痡�� ����zU<��@'��3��d�om^��z#�!��W��~!�)?Y�Oۜ��?h͗MS��v}�0�����?w�$���������9��+S]�.����+u�Ԝ����ˆg�� �}�ҽi�����ݼY70�a4�ر]|��[��uotP�e�a�R����T�1�p��#wE5@��(�#j�]p�T��H�Z��)V��wy�b�3���O���cRl�1��:�2����=�2ޠ�q��%5#v!ZY��l�jJ����}D�a�����Y]5��]�E �6��Nmgf���&�K��|Vq����#�j�+%�M��/{�Z�Te㲟�}ɇ�Q᳛X�nneb�|(N�&Y�<x�;<`�O45��B���b�2m�#W�SU�|2c!�R��[z8[�a)7���>��X�F��Y��z�{c��v�uB�:�V�&��t8�im.�����zl���6}v>�od���x����}�j�9
4���k=a�ݢ�.�Z�R��by��7�Uؒ+Ԩ�껹t�O�v,�>M�l�#.[�ܕ�|���Zdo�[!}�#Xjȭ��Vc�������AW���.�4�뤣�΁���S����|��U�VP5� ���S�q�M����[�n�bCnn��f�cs[�ik��E��j�FҾ���g�:�D(]d7Zjر=a�ش��YZ�r)�w��'^�vu�o�QP9�2R���F�>$;�|�!�3��(f&���aqP��h��V�|S#�3	 (K��)�u��t�4XV(���~ݫ�8ߡ\U_�Z�r� ���s��:���t���:��������zo�K��6�%q&�I�o'���G�X�m�H�7�{ ���fgw�ZJXY�9
z����0ޱ��;}�ˆ�C\���m�ϖ�a|k�kj�n�GwEZ)����������Wo��I�����7)�A�
�����j�ٝ�wwA۩�;X#1�Ԯ�L=�Y��	�ga>(0���*���0^�O�'��}�;P�3�]Xn�q���@YH��R����zM���v�gnb��y�HE%�9mC��ԍ˲d�7#��+�>��t�'f��Wepm�۹�-k,X�rkK�ܮ��!<�ra��S�IO6�jSe�:�Xx��v����"Nj�ғ�i�T~[C��QPD'wy���x�:�E=\:�ޮ�i݀�y\Y.!�`�sIn�c���Ts1�|K��{�:���V��8���B�^;�/��ݾ4��n���KWs@�T�2�o+���>� �nX���A�����)�-�KoN�XKE݂)��{��c��eҒ�a{b&L8�W��'��)[��l��W$�DgjgД �f�yδ�� �U�i��G��D�M��ww�I΋�_T��;��W(�S�;��]ꑰN����36��*�� ���q��Y�n�%��Iye]*��niM�LgvE|�ɽ��Nk8˛����ѧˠ�Ħ���G���]���3����ceJ1��QE �D��+YQQEDb2(+,UAEPb"�U�#TU�EUQE�H���J�ڌ"�T��X�1X(*1EFH�
ª)*��*�FA`�� ��)"�`)X�(,PY`�(��X���������X(*�,��
,*E-�k
�H��Ab�����(���R����Ŋ���`,PU� �V""�T6�X�AX�)A���EUbō��0b��� �����"��TUPET���
E���E�Q��)F1��X���$QA`*�@X(*�*$R�Q�H�"��Xpؿ���3y]�z��7��à�h<N'�i���_y�����;�{M��*��cO9vV�!~�UF$Sm��r����׺�ٹ���^�@B�ب�Ӆg��9n�������o�n�N9s-{��X�z{ݧ�I�//-'��A�x/��%UܠѺ��,bgU�ڕ���_�՘i�:)\������%��;l���F�3���I`>F��.N����f��0ö�T'X�˕u<��G�]rWd�7��Rt3�,����9�ʞ�uY2�uCs�-5��Q�7�ު>>�;��8 �ȯz"
�� *��dNU��˵�妰�O3�W�udC;�KK�T���cgU�U���ߋ�>��Ʀz�U���q�&��D]zf�X'Ə���Y;Z�K�i�mo�Z�� ���9�N�7\%Y�z�;u~3�>�aۉ��7Ɏ��q��}��ɲ{7��kG�!Wo�,.#6�����0mf�(A�u�8?�x�U���o����>�z�~�f&y��q�z�p�>ZkI�|5ρN��1�+ע .�M��?5��ű������oVT�1M>��=��"����6�)x�#�Al����R�5!��l��*�Qx����؜�i)}�#�8�U�P�W]���ݣ[j�a��|q��ͧ�,�wf�	M�W{�3���Q����/9 ӣ�N�v�w����17b+�EΗ��Ku�v[���������6�=�i�u���"[s`�1�;��U2)�Mwj����
E�ʞ�nM���sz��5�R~�p�B^R���N��7GW����=U�|���Uc�J�&��aT�c����g��z�<��Ww�;C�N��y�����14����Uy�}S��������S������ �Ċ�=��ӗj��=��_Ie��t��!԰Z"Z�~8Ґ�;M���9�~T���z@R����!�N���v���M�޴Eoӑ��]N�(!n�j�l�����^��o�L����i�5�FO��q�d���Db;�^�O>�p�NY������`�źm�c�\����?��c����Хz]Dz�F
ߥ�*���5﵋�W��[�z;�O�5s�E�<<=f���D6P���L��|@�K���ׄX穝S����P�M�n��{5A���Y�������A9V��}uZr{�g�SU	��V��<�&�V׾y��~?�z�x�u���ੇ���b�'7�*+�d��YK,pfO�{;-óLE&�c1G����o
li_���]X9/ي�ye��Uv��,M��+�nPx2P0��3ō���Q=�Ԙ���&�z�
��p���q�:dh�C�7ם�Wg����5���i:&�z�����\/u���_E��.�mus�+��<�ݻߜP���ѿ1a��S��}x�f���j�<+#[C��]��棏�~��븽�ut��	��_�w�?(r�t{0m�jv+�����O���%�"{l����wN�6Ⱦ��$+���]�C�2��R=�6ʡ.��� ���]�V���?l����o�C.U���_�w�������w7m�{�7գ*{��2Y�u2���o�wy���T�:G|y6��-w�g��g*�CU�8��3鼞����'������ԝ��'�F=^��+q-��{��`\J\0��7�]鞹]����W'��#�S{�E�v�Lp�\�PgǬ� �w��,����P�g�	����Z������3�ݬ��J�Dg'��d�]�s-����/�c�ʺ,EX���j�B�n���z��'�KIg��\!����,�s�ÿ*�u�MUzf�,���.�3E�CޛyR�3����f��d���x*�������2_3��Ւfp^Ȟ�2�E^��
������
�4F�m�C�ZbWr�.]Z��s�ny2�Y�W���Uj���Dz�4��J�L�յح<��-���xh �=yT�Zo7:�ۊ�r�'�������'p�CB�83�����Wd�Zα�{(WWdV5"h���p_��Ν#�%���լ=�뫁���,,�:Wt_o3~���:<#+�Ǌʋ�ߞ?'�/�K��@�ww^��u�~c��S���aVK:Wt\,e7~���Jq��[�|�,b���9{�1�^l۷�8V���3�]̕ҭi�����$�n�Z@g�T�������y�r�+�a����@hU#;��
B��s�V�ūݽFg�YD�8RD��K���֒o|:�b�N^�@U=��?"r���i����]u<��Κ΃g��ǣ^����2���ޘT�@9���K�9�^U��>*�PLU�Y��/��%��k�}��w�,�?x��k�h:ū�����8���E��U��p�<�T��!>:h}7�F���囗��?b�J\���)=o�O�zK����_'����NW�PV��;�ʊ�os��R�y5�c��e���M�]�,�4��WW��Aa�aƾp��ynt�����Ǽz�����|0o{$��'ˮX���q+��%������Xx6��V�X��#\�e�̦����!R�+)��k��1ht{; �PG��.��ʱ缵v�Luv��
�<䇙b��A�����x�u�:��٭���[�jӤ��9i�ev-����5�a��r�Dw1Yk��Rn�=�![�Y
�9�ǃ�Ə�+�%��-���!�3�Q<Ox��փ��>~lw��ɹ��KK��rw�Cѭ�"?]o�=�"~��B	��h;��O*Z ����3�K�m��fۛ~���a�vt=�}Te�Y�=D4���Ns�����;��lHЯ+���՚PU�y=��鶨X���Ce��F��8�(5�z>ꓞ!�E<W�����n�����Eݵ+=���70*���(J���x�	�o�1uyϥ���������K���S���e����:��umw��A�,�	J�E�����ZqV~VM;�&��4��;���\c����n�� �:3��9�XV���m�4�qrt��; ��o���7�i�i^��lLw�^�C���B���Y�#��eF=vL��9�=��Zp"�L�k��$���z*iL��0j+�h��y�;��	ʶ _t�<�Z���~5 ���v�y���XWgb~��t%�|�h��o�é����3>��4��<�Du	��9]������=���B|Q�E����,eovJ����Ȧp$2�:�·Xuu���Ԏov����mU,��-;����E�����AkiF;s)}ћ��/��o#"���8�f���(����8��R�;m����Y�J��\� owS�qp����H��^�N����OZ�i}��1�]u/*�9L��]��)��-�*����rq�<�N[8.w���M���f�ګ�4��ౚ�W�hA��p���_���Ye.�y�	��x�躷K6�:�V�#I��Bx�9U9������P{{��<�ޯ+��e�#����V��~f)��8{J��o|����|�ˋ�Z��X>������GhU~�o= �K��9ST���S�Lܛu�.o\��Og�t��>�=	.���Y'M����^�!d�f���V���U�9<=��[�7��a��&�^Qo�O�۠���Q"��J%O*��uvu��h�_}�8��S�䡯H���ә�s���ðl��Xc+f��,ЩN�!ԦH�]o�JC4������l���͉,fsR{~���]-������R��Ys���]N@�[�%����{��>w�/m��m�T�A�r��_K�VK�j�F#��S���p�Ŀ�_�(:��� �\���]�[/}�0�³�A�V��nჶw0�,c��2�6�c}5���9��<̀��;�oC�b��+K%�̋��[J�0N�o����iz{�Q5j��zzV��6r�u��{z-n���n|g_sO���_�Y�t����r�4�cxHj�t�.Ө�Fl��+��]���l���7��\�6K��P��[Q`���OY$X�I�[a�����Q���o���PE��,}�;�DD�w��f� g�|@�lI
��/]�i���_�N\�뉗w��G�z�w�״�Pg��Vf��'ڤ6:�A�T�[�q�/�e���SK����m�\����BW�0ץV���#᷊�g���<r����i��VP��Y�VH���f��W�Z��h���@0:���Bxث��C��WT���7��XϨh�2¬�2��7�*�i��E�M�	�x� 
��÷�7-�{0iE��^&������w�$پ��#>Z�&UF��g��Ͻ��r^�ʇ�td�]e���	�}&���vh�ej|W��C=�!8�12����tT�Կs��ϧ��m��]`��ӡ��5$��5�kQ��,�4���&�
�إ�u��^�"�jq���^7�����uONVKl���LSʞ��U+�R���<h�A�v�')���jU����o�� ��ڙ��0��en��PL�r0ם�^����P��bYvK�h�}�[�W����o�6L��|��whW���bfDx�`�Y]�x�m��p��U�.�vCv��L¥�W5t4���]���; ݦ�u�=z�N���q	{����/���q���\�ܼ���Eǔ��.'K$y�ϓ5�Xc*犀q<F�C�w�eR�ľ�
p�ŷ�fe[���[x^��Vv�C���)��U�72���H:���U� �u�C}ᡌ1O>���8G�m�����9�k�q{��f��	cݘEXf�Y�Ԧ퓹�S���ɝ�=A����xV	]q?ڦ�	����38/VD���F��EB�Oz��*���ko���,'�=`'\��0,�:Wt_o{�kGe3s�P��!����N����z�ŷ4J]�� ���
�,�+�4�ϒ��}���gO>N�Fs�|�dy{��/�Ł��7{#W������x_ǰ2�[	oۏ�qk��K�ߍ 3D+�߭-}[$�kJ_�b�FVLΡ��g�@`~1�	�ڳ� S���<=�&Ko�7�upO+�֗���]�~^�	U�R��qS���3����*�g�,e@!�S.�;>(N�̿{xt\K���;��b}�o��綡F	�� *����yo;��p�|k�!���Y[�׻!U�s�~��e��f!�8a���^V/�3c��e�9�Φ�ѓ��U�cۚ���-��0��%��t9C��3Ծ�6�㶷f��Y�Ef�A�bV�w{'�vǽ!��4g27%Je�;j�����):"+�u���)Nr���qM�[\X�%���7��׬�}�ë��n�B��}��^�U�}���A������f�6 ��:�wG��z,ϗXӈJ	�:���˃=mL����(�ܹx���β��<8{[��oj��s�r�(4���.�&��hAW���/��-�[o��%��ǣY���~0F`�QA���u��n|���$�z|��OW�J{R�M�5���=�2��w���g��g��OO�p�7���D�QQ�����a�x6�1k\�w����|�Ǟ>.����zHo&�(`�������y��*L'�N�i^ڂA����Ƽ��*��J�/�lVe|��L������{+�oދr���J� $�d�s��F��S���uu�V.E����S��ײ����"�+wI��	ED�������X�� *���!8�&�w�p5/�f�V�j#s�./������<�j��=B&���0eE�Pg�x/�x�WlWY���d
�;s^��9;�3�v���"���W�9�*������4$*j�/��F���e��ݾ�W}RoV�#����[|]nѬvV��jbt��ی�:��ݾ�Id���I�km'�p`R�ȗ���l]�6f֡�L�����SY��ޙC`)^j�y��k��渼n���.�o݂u$=Z'#gFN9�^� �d�t�;�._
�Wlv'�sh�C���{'����l����&�T):%�[AS�<\Īk:��3�E��*�8��Eh�υ�:�/|5���+Ō�`��z"
��N�2pR�������')w�V�*m��ζnn�F�h�2ݱ��Pxf�L��3���Uo)@���azO��J�iw��藼؜���ǫk/�O�٭3-<��S؜�W-��n��q�S
��;ɕ�]ҟ��,Ɖ�>�~�8p]/A�e�A�ĸa/�^������7�%ty<彌f�ʼ2�s+ޢ�pݞ�Ī<�\� ��Li�l�Y�s�[Ĭ��QdW�WR�#�G�p`��m�YO��4�p��d��[����}u�G��5{}1������4sδ���&[$o��NT�9T�
��<9��k�GV�\��#ܖ�^\�ܔ�̽�e��'½e��u&%(p�Y;^w�ȉ2���/W��m����P{y�	��C���Vj5��u���|yQߐ��4�
o�$��tr]g���%���ZV�s�"Ғ�St����ޕt"v:3Z�7�sRv������v�P�D�4S�k�ή���αs�Д�{B�b��v�rR�cJr �iJ=�b��*�PDۺ�l��Uٮ8ò�U�jG���9�]�����D�D�2]��d1����̭�w�&�LǮ�n�a�əQp]��»�c�!׹�@�1H��|^wm��^ ��z�=�'e�..�R����>��b&Ű�^�t��L�k+��O�jI#�8erGx`UIҜ�#�+��=����<V����7��^j3F4(9�Ae��`��+��}�r��uj�ʏ�5pi��֥b
4vE��m�@��� ����1圆�������������U�PmL��3�9���k�U���*��lR�9�Y"�{L�������Τ���\���-���͗D�î����6O
�����<�R5c6e�g���QVAI+<���:��fq����:-�,e��|��U^L
o��ڔ.��d�I��vj7��%k��q^-�o�(tT�K��bs8>�E�����,J�R[�]���bM:r��>h��k�����٥�����x��%j�õΎ�B4��O@�s�[�������Q�T�uz�,ۡi���W�-A� X�J��W`A״e���[U����X��-�����*��̳+��gx3� I������͞!UȣƮ���%�/${�W�4��tW�ͮ�=^y*1�5T
�t�R��¡�ˤ�����*X��a���:*ky�yI�n�5���*!E����})g@�"l�)tVe�W5EϜ�#��ݵ�%���1�(u�Z��,{t�9l������kb��R"#-k�%�uq���q����Eea�J���z[]�ř��fZ�祥]}�7w�-�?��~p��v�����O�1�bX��3�{o)��J���U8X��K�C[�G������Q �B�5��V��+S���::���V�v�%+4�هI4n�O��v�)w���fYe.Z4O.�,˴Zj�]��:�C�ôOb疨�꒹��'�������\�$ǒ��`u�r�S��>���9f��#���}�`�����Gso�����<��p�l�u��:��]���ե���Dѵ�iݣ� C�4��*+�>�2N�y5B�Q�`��.�:J$;t�F�fY`<��J���%����]�����W`W�����yҹt8G�,�FD,d��=Z�/Z��n0�if�U������߱bp+;;6�WX�ѓX�;-�+k_+8�s�a�[;ñ�K�M2/��j�N�w��lX-.N��f�1<2X�l���\���(ٗ+�UMR�d��y*��E�v�17����%.��u5�i[7�gw�V(��V,bE"��,H*����)8±E$PQ�dDE�H��((d*2,b���AV ��(�����(+U�����,�" "Ĉ��6�QEUEV �b0UcTQ�0DQb�(��� Ŋ�,Qb��XF1�,�(���1db�g�ʐP+YDPUV*�"�iQ������Q��6�QZ�1F�+�( ��*��F��(�U��Ub*AI)mEcY*��F2)1���+%d++Z��
T+*TX���,m�0�R)���"(�)+X�*�E�(�%�c渭���ٝ������`�C�l9��[S�Uf�QJmz�\�,L[2�$Swsm'��ö%K%���)���L��_oX�� G��D�̪Q*���X�����<C�\�ۚf���yr{��_e�*3��{cCE��,�Q��� �R�h�k���JC4�LM�=�b��^xθc��Wdo.�5�1t̮ß9�1�Y��Yd����Ϯ��k~�R�၉Z3�e��������JSִu�[�>^g�˰�]g����2M�A9d2L<���<�Bd9��w���GN�m_ᣄ�_|ה�
Pt5,��e�J^R���jy{6��s)>)�9�k�o�n��v\CX�7V��戙�s�@{H1�G/ak,�o3t�AR��I���K�����B��vҕ՗��ǵm�ـ�m�L;}V����+=kژ+�E��������,xNH�^�6,G��+g����^�
t߶�%�b�3¬>��3�k�������} ������V=>�!���+qp�����e�z���O�ӝo��g�'�襮R�g�f2s鷰�����,�{0m�j�د��\pr������[W�![�ч\�4�3� �;�W.�lX�x�i�z��/<׊i\�o�t��b�"�g^V�9>L����P��*!y�dZ&>����ۋ�D��W�y��L����[��WY��Ѽ��\��p��Z���7*K:�S�`���r�W�ϣHW���Fez9���K�0�G��-�r�c�+r/o�s�c�׈��F
f��9�ġ�.֦&U�����){����u������
5�W��C��*�y�,���
�|+=��9z��jq��\U��B����h���K-�a���;-���S�ö��<3�e)[�m�����u+��8&�xl�c���ڂ=�/:�b�W�K���Ӆ��ʝ�1�U�Q�<B�:N�cHV�K�ȱ+���:,>�{!�T���yt;g��p>�����苭��y����m\%�����}�ى��Z�O��?_���*���X��w�v�@�S��k�0�_qd�~UhӰ���_S�C����*Z"�d��¼u��{i��g����38/VD��	�jJBѮ�����^����ޥ	��zf�cՌ�;�}oz����ã�����Ͱ�xɧ��ߗ��O/`g�| ���xVf�YIS��-��K:UwE��7~���I/*Q'`��R�7\�Q�*�����r����=�Od[.Y�0J�,i�t�'9��z½t�r\,6ӺĘ7��jY�����,�	fPƆ�	|��@^l�6�fY���&etG�p�:f�,u3,�����۽+n��f�z��2���}䗭�|�={�x���hu ��9 ��µ�G�y��\�]a�f�#|�-��6����GT�͠J�b�o1��,3Վ 4(q1ߕ��u�X,1�}�+bk���� ���̛�mk>Gk��$����� ������6��9f� ��L�LttA�[κ~��T~��w�s�N�,�=q�C{� *��
Ny=����*�Cʇ�N�o��>K�r4�ѷ��hr��|��t*����LuG��J;�ŉ}���[���=���y�����nmozl�u�#���U��te�A}n�AW��t����6#~Ѵ�-5��=gmL��zf����Ԣ��>������o�[g�.�&����� �\<}a�̤�����{�����Q��̃������yE��~�}e�l�xF��^
?|��]]��_�C�)`W��=�
�ƦS1=>�-���)EFD�=�_Z'���}�R������ʜ/���RW���&�R��?ϏW8�s����(I�+�Թ{�\:��W�n���BEm_� ��B��������;(-����R�ݫ���=a��@�4~Gf,����I+��d4��uck'f�d-:�Kfe��he݌G(��r`6_)���N��h���t�jwZ��k��$)��i�d|��� �B��]C�#w:���d陰m�;D� N;�Eh��3�R��3�-�ǶC8!��~ћ.�=�]����m=�0{��vԍ
� ��4�F��b�Xʾ���(5���Rs�-���>�N�'�����ӻ�4��Ld8 �&��� ]
cy�p�Os����<<�Uj��l����]z0t�u�r�\��b���J��О'�w(4~���b:�)���}5�+�-p1�����~��FS�Q��N9�}f���6{���X e�5�z��RG=}����A����6�Z$�3�'C*K"���,x�=�S��� �7���zD�o�R�W���Ԕ"�`�"*��*�� U;��
��`].�/Ul i�z|x楳��8H�g����Զ˪^\/.���b��}fٙU���r�^q������z�o�Zt�|f(5 f]שB�e����L��~'�߭9�Ncu�Y�z��W�:m��v7�˸���52q��:��A�e�A�B�H�%�<���@��CB6��^���;u'�v�C����ܲT��߭�]N�nԖ����o�gpS�Ej����7v��r�:��\���Kơ��:��KU�������W}̮�?��(M�۩T�ƕt��dC��sj���twt�w�S�)D���=Q6������T2��SIq*�.J����?^��4�U�����7[�P���]r.��+"^.$;T�htB�w`�sՓ��u�=����=��d��z��у�X܉���r�Ɩp�1��/�������	�r�MPPs�N�nM���������g��yh�����שtԦ!^�����%��ּJP��|��QT�391x�N;jO�~M��ܼ1v�٪��h����'�5D��R����Iu|�{=��5����7[=���4��|eH-����5�`k�Y�e:�u/���x^5��r��q�ܑ�wx��4�����(+��2�9�1�1�۸9�A�8Bnuj�����8��}j�������Zu�,��a
�v.����E?��+��
JC9z]м������ҼJ����@u��|i�o_�����T����pR�yJ��Og�sz�E�]�A�{����d^N��	~Y���z�K4�{�B�f� d���O����q<�K�1o�X;vv�қK��k
�Ұ������vV��:��3�[8dt9��/�/Їt*���+C4��GGʺ�x��铴4�_�$�+�í�m�<���f[�7jV6�W_ǨZ��}�R���;��RɛS`zS[3�G���]�z� ���9��8����w1�O�
����D���
�g��a��M�=�<�!t��}`z�%�F���X�m��cآ�wN�Z�Sq��6�o;��d�>�Ey̔ A��h[=�	^6*Ǹ�s(�WN.l�.��Ȗ���q�픦�oF����'^�[ҕ.~��{��B���,�����U�G����dO@��c�<Lf�da𐆵xL����Q�Y��>;���W��ߩҫ�r܋�t��q��S��%E��p��x�KZ��nf{����ѩ�x��<c*����x�6���ɥO�}�X;��i5��<�$AU�{���a��EUmN0l�V]y�OիC�ޒ���.�J����(x_o�ug��R�[g��Pt-@��eq7Xy�|z8Y
����������{�>w3�����N�˞*=g��BI����V��Q����	����P�_�MG��wt�=N�Iԡ��w�ag� X�U}D�����V�x�]�QmFU��
��]g�P��D.��ݪo4���]ŗa�z�v!JPAe�ưMo�ܐ��j갩{�ȕ^�{�ǐ���hX�u�LK�سy����W�Q��������i��״�(Q��n��P���������x\��	�t�$g��/B:�T�eZ��z��"*�Y�W�a��d��4ͽ܋V�c{�����J2�����a���N�����֔���>�W�w�)|�XZ/�3b��+;��Q���UB�ԙ63K��x���d�{��n�c43`e�jm]Y�I�����b�Jk�`���D����.y/w�Bz������Z�ݭ�^bF�T)>>pZB=�f`�?#j��W�Xد>E�_{9��I!�������HLg����ݫ�G,3ՕN 4(q˼3~��+�\!u}EOZ�G���-v��s�i�̬�vY&��_8�n/3�ʯ��!}C���=��A�{B��Ց�xώ���7��,z�m2����@*s��>�{�;�9�\MN��r*Y-�,{�o��cD�_*����LuG���B���&����E�z�Z�V=i��<YOi��c�j�>U���oJs�')�i��U����_��K�u�m��¡��k�K/G�Az%b:���x�����~ѽ���m�ю��C�7l��H'$�����҆��p�Q�ݡN��q�#�4p�Ӭw����I8�f�fy�j����v%�m9���۠�lx#�K���A��=xg�yi�+�nSZ��<'��s�F����/�ꏗ���}�]�3.��VJ�\iЉ8%���_����\|r�ze[��{�'��0{^L���~���Q�>���	\ſ;�Q?w����0���ۀ�:�l¾�q���OO�cx�HtL�<l�K�����1�ai������jv�&�q�� ��$y�xu��?s�=\�9�z׺i��u��r�S���1��HJ&(*'t̳|&R��yu����RWc#��y40���� #����WO;��>�ޯR�Y<�v��
�(1H4�|�bh���x�]}[7����S�m�`]�hNw�	��Ɲ��=��O�L��w�
��� �� ]
cyQN7����;�(j�l�3�c{�ƅ��7Һ���f�r�SuE�}Y]�&�|�&�R�G�[�UWOu��"�n�_�G����C�ԭ�^����F|�v��U8�ʸ4�"J��Gx��h1�y�@��ێ����U�Å��go�OP�`yP��HH�P�,x���eN�� �U�d��*������\F8�����j�)T�� �]��joU�4�C��]J���W[��*ܹJ������k,�=���'s�7�b�=�7�� /H�5V%Jȷ�w����38wC�h8�6vu��:n�'][��)�����Y��&Z ;�:����i��v
B�X��U�DA[� ,�dr��w�E0��g6�?=[v�b�Y��ί�L,f�%��۬g+���0x�7�b�|��F�O�ŗǽ\�gi:E�gl��z�2R��d�>�/.x��P���? �uQ^�֮���zz�s�{k��g���_y����ct�����75X\Fz�U�NC\��={��)L��}�s2��a���fx�0�ݾ���e�<ý�)����C�on	������e���`�4e�7עUU�����=}��D����O�뛛^V� �y{}G�ԡp�G�a���\�k��Fy܄��*.vT`�y	�:]���t�ɣ_�������)�\5���+��l�R�e���<���$e�vnn�'	~�;���=���^�cC��L�4��}D��UR�W|N��fD��Z(�(&��,E�Ch���0L��C��8�7'{,pօ��YdPc��\�i�!�}��t��3�3�]�k$T��X.Z���u��}Ǯ�Rɛ��g��Y�\�&�l{�� y����n��he�.@�R�"þ���V�����v-V�;Ư�1�h&C��.�U�c�Q�H����QSh�;�޽�}e�3Ȇ�{7{^�M{t������A�k���>��3�l�;��0)�x�)�
��L��.x������Uw20��[Jd�n?��#��ml��u��e��R����1��>�]�*�ػ�$�4��*��x�T�9�ۖ��e\�]��4�W��-,M��^P?}
����u�+�� W��a��tŷ�1���MI�*ؔ�ךX�1��Pxl��|@��k&���X���>-��7�\"[T:��U���V_X�/�����
[���'Z]����X�ޛ#V�ڱ�6'�ATuoI����P��Q��nYnz�pĢ�X�ӫ|j^'æot�5��~�y�T[�P��Ɯ�hU�ȅP�*�Y~���9`Ӿt]j�d�2TSٕ+y�;�z����E*��J��L�s��B�O��]�����ʬ�~�ձ홪�x����6�6�>$!���3����Q�Y^�v�}%���m��z���Ṗ}��>����#�FsM���ې�R�be[��ާ=4��.#����IUX�񧚹�uo�e�C��T�w2ݫ&
f}�~��mJ��K��nI�MaCvPyK��2��PXQ������)_Q�GE �d�I�;A�7u���V^�˹/��A�ذ��9�%I��u����ز;&vV�2�l1�|��zC<��]�%tެ�Oc�����0�Nw9�]X��C��@f��
������!�9��q�z�k ,����Ѹ�*h��^ϑGt�H���g�8�T��Hd�
MK����]
��X�v���]���j�{��i���y�����Y����ɮ�%Oc����p4�wf�����
P����W�f��KE�U�`����e�~r�\�C��X�f;�*"_S��u���M�N4�� ��իkˍ
���0���\s�z%u��&ఄ�j\ʩ�.��j�Z�j���X��nس״][��0���b�W}ҬR�:��:�#��dTg��ԍG��׽�Y�C�(y4U]�O7�l:�ȶ�	�+�]��u�|�(%��RD��x������շE�|2|��"T�{�Z�\�������C�i�T������
S:��l�3d��nA.�q��JD��y�g�s��g.l6�ƭ6-&��]}���T7Ӈ��{ة�MK(�h77N�!���I!�O�4�ِLޅ-�̌�*f��G�Y���_��h�ݺG�	�м��j%A3�L�R���)�q}6���(`5�����e�MT���T��;�
��q��N]�ʼ�&x��f�+�vYk����u�|�ټB���)̘��0�G
qG��U����XOp�/�ӆ)�e��,	�v孬�����D �5�C-���:2���x���k��fM����Ά��Z�sawl8�o�S�շe�o:�[�2ȸih?5�h��t&n���i������@)����n=��Z�M�RE�7�Z�Y4�}Y��R���a���3���Sl�f�*�S+�k���]��^�*R�m̾�nѧʯ{�H��\��*�T�#��S�F�T	'\�{��5�8zvwU-�oT�nTFO�p�����r2�-�g	�*��7����C�|��Ƚf�c�~�����8"���h�%o�]��6�tH���~I�D2�r��N7³��Y,1�����F���'v�G�����%oK(1�&[N���[����U�r�K4YV�X�5kU�rV�n�30���x�@c��LF�K�c\<'��w*�i�ǖ�a�rq��74I}3���<�cA�I�e�[�¥1=���@��1˳�S�V�2��ƥ_b2��gm-{"YҠ�&��6��)-=	ً�]}1��ce�+HU�Xx�%�X��}�k0%-cl�0�l-�p�����,'"Fu	Np�l�����@�qjϵ�spU��7k�G��k��b)�VXTQEE"*�Q@b�c�Qd��*Ad���X�V[T`��$*,*,AV,U*�PR#�XEU��m+��Qb����(

��@��`-T"�`-B�YE�J�"��1e-��Ab"1ʑ�E�)hQ+J�,EIR�,�J2,�
Զ�`����YP��R�����*X�h�QU-���������XVUTXEKl��X�T�Q`�(��U�Ƞ��PR��FF�D�ET*�mYb� �J��YJ� ��m���TYm����ݭO���[���h�rٔ�0�8�Vm�F�>�@�148LM|ƭ��k7R�/�u���!���}՛�A��ޡ��~��*3���;?yA�	�gǕk�QW��%���r�-�9��e�����8t���f���[��Y����/���ޣ2��
A@�+�&Jn�smo�'�7���|g�냾w4_��:�⥚_�3%��B��ۚ�Zy�gJȽ�Y*�h*�hx{���z�t��}8_�M«rL��QvC�Ǳ{s�#�eH�x��2���>��"����?D&k�8��
�lh�R�,��Q�~�[=�DW}���VZu�R���"��X8�x{�ip��8+�I3���*�q�i95���U�B���b���R/�p �u�\OU�[V��Eٮ�gĚ�2�_���ܴ{��Kt1^�zd˃r/`A�
�K<	~J�O�,md��q�:��S8j��v�����Y�3]!Jq�����̨3��1[�}e����̀b>�K��DɎ��쬎�w��2�-�+jD��,3Ք�D
��؝]`RW���k���G�N�W��K��곱ȣ��P��̡ݺ���+����ݜ������S}.�B�*nkx��aj��k�(m�Fx#g%I�ٕ�!�ҍa-��	�qWo�s��)�Bu]�xZ�c��d�Ժn�N�
�R�=���z�K�R��YC�+�%�j�7e�]k���:�-�'�:�!%�}�4(K(���{Y와���@pGW�O�p4�z[���=�����wN��y���xǴ���o!��by��yCXg�m�Ya�b������͹F����L�����9���i�������U��5���(|�UG\)4���SǨd>w��۽~�Ƕ���|��y���Mxn���l��pǍfz�}Y��0L�뗲�1-V>�ȼ<+�t��/��ә���~58��E�=�q6p��>���y޼��8Z����h� !�0]=�3�Lf)��S���|$:[�,�=ƅ�]�\I�1�]� ���7�5�!W����{d4�;՟';��h��hE��;�]���w���:��3S҆�WC��&�E N�����q3�¯Kb����~�������o��c�����ۋ3=�q��v]��H��)��!���B��9_T�XĴ�se	��zT,��P�'��%�GB<��- w�֝#/��YC�D� ��Ν"3��Ja��T�o�	�wc�։�7g'BuY=�Z0�d�uf�
�s�D#u��S�.YD��q.��,�5*��F���\jj*�Y���ÞY��ݺ���݈b�O2�.w�Pz`�=\�,S�Հ^��>���FX�ו���xncf}���%�iϜ����{ ���A�x���x����|-��Ws2jԆr��Woϯk+D6ջ���צS�)V��-�.�����}Fy�R�@�P�>�}{�_��,z�Z*�Ѿ���a�mݱ
!IА�<+D�괏ÿ1⺟:|<�Q�·'D����yh�Ip�Tˇ��A�u.�a�m]��y<M��U���	O�KR��=������}�Y�_R�/�-�o���a��È�ۃA��J�w�t�"�o���^囔�����;�y�J��2R��2T�&&O�_�����&��{��1j)�T7���@�78z���i�e9l���Ɏ���2�/"j�D��r�/57������K��Hu��۲�[��L[^���i%�j�X�p���k���Fv�9{�T�g$G�˖�U�U�.�������<�����.x���iR^�����H�&��Z.�<6{^����>�,���&[n��i<ބ�ٻyj��0M@vD[��P��֬�\+��á^%�}�*���Nm�q�7�9]CΉ�R�oI�r�:��<0��K�_�ԥ��7D�]��rw���6��%�.덥�).X�p�>(Ϭ�,��;Yr����5�d&m���w�]ڄ�Wo��G�v�ތ̖��.5�iOs��yB0Hz����*�2�t4,���'T�Dw�}R����3tK2��(�xǾ�.k��t�K�"��|O
`
c*�%[�_-'����������#/���߽��xC
y��=_8-�ϧ{,p�ׁR�,�,p߅
�ϓ}��uj�g��~���A_�vL9��x��]�S���+ߜ��9NiLel�h*r�(�NNn�����s�y�<����H:ؼA�W��������i	��a�w��v9��Yޞ����7]l��f�ݲ!*��Wprˠ��I�ZX��漫����T���
8�:�a�N��SW=k�e\��h�U]_��M/���U[�bPw��������8O��8��O�I۵�^j^x�J���wPj���/���V{LYI1�f�2���7�M�,k�f�-�-���J򉙹���eA9V��KQ�P�>wgN#�ȯ,�G�2���eΜ��1��a��Xχ{;čTsWp���YGծs�-27:�TK�3�*/��q���
��gSơ�Î�]�����)�!f�c5	�d/�n���=�Ӷ��wrv�[+�"a4c�h�8��>�I�0�e��ss[�
����)QT��C!�ƞ���D*�7F�fY���7C�OrF�E~�6Ƿ�,����bi��A��[ҕ'�9N^�����隬o��l+V�{joo��wAd^]VA��g}e�� �B2��	�B��q�Y��^��[�QF��q���}\�h�xW�ǨB׸���Еx��>x�z.���7uԽ"x{۪���v��̫�S�qN�P������U����/���P /u�Y��K+'ft�"Q���B;x8J<�`�s���"����X��b�ܪ��a�tza�v�e�By�¦O�i��"�{lGq1�M�{�3����C������X�R����ڸ�e��ne���W^�F�6���c0s98_��p���L�ϕw�o}��w���Q�2�����;�ɭF��|>�^ܥS���Fnv^���Eia�a}^6�kb������1:����1J����mK�/D�u�����/6v�j����댵�U�����S�s��#=����:V|nPs�-����u��B��n��@�u���hKcC���W+Nm}w��Y�����kʲ��g_T}3�(����*W9��1i$+r�����Muv��WnLv�v��,�,�����t:�:�;�%�;G��( ��PE����0/��B��v�d���5�V��4���4�z[ͧ�+p�ⴹ��p�@8O R�#��c�u�_��W��^��<�N��o����a<edk�g��CN����V|`�W�fTE�")��
�u�nX�z��s*i-8�I�)��Gg�-f�0d=C�&*NU:�?�c>��=y��3ҁyy���d��+¬j=�ՙ��>f�d�9WFH��p��v�X�{ �ٸ�z��4�N� ~���0� �{.�߇�Eu��\��ݶ��<"ޘ_=P^�sy�^�to�9K���v<�%��a�y�Ɖ�Q�.���tJ��TG�g�x�ڕO�{a@D�k�]{&z��z�5�Լ��4�m6{�Sϗƫ��kOe��>^u��G\)SK�;����HV"�ŮJe�9S�MA���0�{�f2;���^��r�����}�e]���2�����qw���j��T�R�ۿ�ʾy�q��X��������� ���C���n
��W���칚߀ǧR�98~�=����z׹Kؓ)	��n�Z9�Z�G�-D&��}zH�m��-J���3�Z%���ոB���ݤ�#�C�Y��ε͚�ͣ���.�3u�7��i�g�3v��?�τΰ=�.� Xx6Sۂ	Ƨ|�SL�X����	��Ƴi�V'w&���/z�0�%��6�Vo��5�\d�3O�!����	��7��C���'�-��zgr���sf�R�вw��Y���"�}r�U�lVeS�C�󩋻�=���wk�!�~Ѱ��;.�z$h|�m  �W����>^^�+v3�{گ*^��Y����k�ʤ�g�E<T��߅@��� ��dt)��F���-�ݬX��͂O/=�9�=0˃�Ե�FIu�q˘yz���A�x�Oa��܊:L�;D��et�װS�*�A/8*CO���	���T໯	NZX⩧*/R���yt��K�Z����L��V�L�O�Q-�%�,k���b��`yP��eT�EmZ4���w�}�ۑ�%sr�����"i��2O�����K�FD�R�\<%<˻�Ay��N�G|������yc�䨈�< ����WO]���ߊ�l{|���)q�c>?|��/q��{e�c��t�DY�$���Up�lf�l�=ԾL{A�9�y�e��\w[r��j�#�Wxx�E�ts&�i���Љ�Y\�И���8z,�+S�&wh����%������K�9���{��gi[שwT�yC}�̵���{��h�Ѽ�"�N�@W��V=��ʮ"buD����<~��~[�I^�.�*3��ne����4?W��=S��^��<<�{�Ɏ�<4*�zT�ۖu�m�r���aK{"�Q�y��:[5'C�E:��>���|\,�U��;�~�'��}ǐ^r%϶�ˤ'�ݮ�����`/�Γ��-`���h�:uY�s������S�s1nZ�/ϟ鉝c[����gb��a��{Ƨ�|��ޛ��kʘʴ��9;^;mz �̳���MkÈ�{�=��De{��՛�L�I�г���	�V
q���Ǹ�N���
f��.v18�޺�R���Q<)����J����iX�3-���I.�V���;nM5*h C�\�����S�ٕb�5��w�L�y�$�]�%����]sĊ4z��8�;�
{�!s��{�]���𕞌��%�c��w9�ء�U)��A��`��+���y���/����#V:e�.t��(/�X<r��D=;j�L���]����s<������ߔWr�)C@��%Q�لi�z��{9�2��v��H*@4��`j[���v�k�P�����jn�7�v����[���]N �I���x�ԑz���{����O�JJ�@ŷc����}��&�'S.��@;W��-,M��5�]�S1A������/ng����yu��	��*��tD�Z��%�m%/�z�C��5�/���o�$6OA3�qozv�窼mq��-�R�Q$*���
�mª����& �ۃt�=M �[5goJ���}��M�%}7$6 ��o�U�9],gб�Ėk٨m��5��[:�o�Q�lg3l\�mz�a���ڻ�\�QM̔2�iΘ��Ȉ�#�4��˂�.�Gk��z�ø��r�{�շ����moJT���d㗰�
���Ӎ[ï4a�{��ޥ+�.b>�E�T��~U�^7}�B1j�݊��Q�\��y�v����[��VjC����vk����U�(u�7IFsM���2��/V�L��C�Ѭ��Һ*�k>�j>�o��W�ZU���#�1
@�(��f�)k ЯN�sq9�^��[qwz*��S��������X�Q�cr�Q��JL&x���݀_���#cV�pu4?n��,�A�ՅҎi��tc�v�=;�˷F�)o�G:sd��v[����/1�Y�t��U��+l�q��4L�
��F칂���Wkn�a�ȴ�8#F.&�*������v�)��ҹ��wm\�Ϩ��B�0��R�}W�t��}ۄ0��pc��Ϧ��=�9�1�<Tz��x�_VrV)m�o��߇���I8Wb���
�Pv]�<Uw�bA̺�/�ʦ�U�c���������{FY�<:�+�%�L	�T/�o���5�^\�q2�P�}�z�����H�K��^����Bi�v���,DxI�°.���rX<��M3��j�s�w~2��.�`u�^:�g\Â�~�( ��R/�b���/�ꦬ_)�..�㹗��[�V��s�z��+���i`L][�u� �+�����-���7U<L��L���,k��T�j]t��|��E�i�����A�eA���A��&`�ܙ@nL�x�B�q��5�~T�-{�Q%���J�I�Ϝ��V|�B�q3ԙy���9�J���:V��Ѓp�)\Vf�x�2��$���TT��N[K� x�οo$q�̩�-�Q��������˷x=�ng�t���xz�mC�G�[� 3��)Rd��� C����_\��ZWv_qUK����G�w4�CӋ_��-}�sm%��=�y2�bm����������rb�e%|�7��k��ڥm�����/��o�wM���y@�F��rkX�±N͠�Ng1��g�8\���·�vV�k�mm֥��w���\�$7���&۸�q�(SǃF=6S�>"��6͋SFg5��G\��N�P#֬��B��o��c�<�˃{x�	�6m�D��5۪��
{B��a�E:�W�7�ǌ!����ś��k7eZȘ�.!j��T�	�Dت�\����oP��� �{a+�4��U��Y��Y�))f�e�]�����ZS�%��u]�*�u�J��Ѭz�����_\�.擸oi��]:��ŝ�*0�Y��۽�ӽ(�r�����@ک����x��p��|�صǱU�ʹp�t�6��%Z��>H��1��w�'&.�-�X�%���[��{;]�J��"����n[�Pm��*n@��$��sy�\�8C���T������f"����M
S�b1���:�eͬf�y2�*gPܬ<*�h�|:�U�D���f7��3����Ν�Ŗ�k�H��k&&ow�sax-�fS�<|t���뛔����m8Q��V6�\�}Qnn�AKIJC��2�����Y��uC#a�OxVQ�G��Q-�I,��u�U-V��D�ma���lZ�T
S7��]�W�5(����plpzu�Ę�{�ӯ;Ú2P)R[����9�v���#�=���-D�*f�����B�3�S�^�[���f'�6Gif�Ѯ��pk�.�-�y76s��y�.�x�ԡNGL���Dz�WV1��%����m~�^��	I�l*�牮�Ը�᠋8Y�} :~�k5�KuSCg9�%����;�^�J/l�O�����u` ��+��o/��k9��.�2��YOef��j�-ZA������v9WF�>�N��+b��]��I3(�/�F�em$�a礕�(�M���s�"�7�������JYO,O���R��(v��{+� g�­��UӲ���I���Z�I%C&�N���YTe ������ �����P�/۔��乐Xz�ifg�G�ҩed8F�,�ىa��;����+��H{X��Ug��l6�PEi�"�f�힐�펵���%7=����9i��t��� �\8/�1-���]V�;tV��L*�,XO,.쎸�kp�	L�x�Cdٚx��sF�1�4wy�xAkv�mQ�{����Z&�y��rE5���(r�B�[�Y� �y]B1���Ywՙ̍Ȗ �8��<�ri�A��FdS���rH�*�D���5�Y�d�R�X�����N�ՙ��J�j��½)4e'�)z��o5n�K�U���iU�D�{l�έ�ml���Z��0�����hs��y��~��|�o8���+%eVT�(�B��A�*�l+"�h�*QQc[mdQ���,m� ڱJ�J���J��AB���b��b
�+(Z�iPR���*Ե*Q��E
4�jX#R�mUZ�R�V*�A-�ZQ*լYEIkV�BңUP�*���D��VV�,Ym�J���md�����@V����B�"��D�-YU*,��
�l�U��(*��	J���2�EYim���i[��
���V�)R�
��h�Y(�kQe@���\����h�D�V<\37	B��^17��U�ff�Ν��D��HF��yy�Y̳&�z�ab�����5r�
آ]W-]��wu�5��/��/_�5��d1�z��g��?�\X������ח�Y�d/v�8���"��y�^��6)^����+�i����������֞�]��{i�����@z�_���g�M�7^0U��Q�
=ݡ>��_/-*�L>�`aVF����[aw��5l� ��׷C�^����v�=W��fh�f������@NfJ�]sH�z������z��fY�W��ͽ];�v�Eʻ�\r�}�t�����g�L�4��iCD�i8�/o:���:'�.�7�,��Ū�.�r�2k��Bx���I�x����V7O&;-�K��$�^�sU׻��W�� BQ9g�+Ϛ�<"���˅C~�N�Nt󼎳�%Gm���:�]�g�q����+=!�N�
�
���F�n<gE�6t�9<HQo�nl�ԟ�}��S�޾�F�}'4�)�^���2��T�,tF���+]W(����}������%��h����Cld��R��q[^�܆i�b:�{ ��E�Pg�x=���^Sr�OC(�&t�:���,�:9�]�~�
 �(c�/f��Ĝ�>�'y ME�2F]���Xԏ�!��	2P�6�l �#+v��[�<��.�mp@�}�sS�����`}������:�OX�H1:���Le[<q���m�$G:3� ?fz��>v�[_#�֨xp{/�צS�)V��V��;M�j}��-�{�P[qF�f"O��Dhg�E'Ip�E������!C���):t���_�[��=3��"*�~��>ے�WZ$�oQ�.���'�]V�#����R]�Ǖ�~�Y�pk��m[�jĨʗ^����}���<��Ƨ�տW-�o�Jl�|�g��w�6x�N��I��c�a�z�Y�M�#�&Ut@W��V=��ϸ��D�ޞ�5�A��q�ƗzY�
���v�_���C�̡��d�W���0xhU�����Ֆ�r�g� 2n09�ޫ�kY�c�3n���N��S	�̯%N�7L�z�^�n��xcGn������f��u��RՀ�*�z��%U�UG��М�r�Z��#��w���n��g�}��A������+k��C�L��E��+v���ꞚN�^���y�^��$��=V(�"��.୫�o.~�i�k롗��6	���YY(fZ��b�ܗ0ۨ��.N�������^Ж���m�=�ՖT�is�)Hb�Ѱ1隻�[�q[����t��pEϘ!^a�&�D+9
�����M�ʃ�Ɍ8J�夆�`�j�z��+���=��_�{�kDr��V�0����g���꧕R��Q�}@�Ǻ,���)��b��w۾�ql�gW��į;bo�v�jÆ��������>�x*r�!���/Y�����1���6���B1n�fiߩ��}�1�+�2�U9�0R��^��xy{�����s�Ep�#ƪS�A[�%�^ �����T|�M��!R�}d�yG��鷋d�W���gz�G<�r�d���GD�5�ʚ�l<<=������ ��J�e.�1἗R��j��S)�~F
ڗ��}�&����U��|����"�X��mf��[��>����Y��vS6���[�3�u�� x���;���$��N�m�s���{�'�����2�UےXt5ʷ�>|����7]X"G�i���F�E�ټ/���=�>GCU�����:�-ب�t��nd�x�t�4-�DL㧄VE�B��/J���cg�aj�����/W���²5�,|,Or���~��F�G���~�m3�Q=o�fI�isY���[|4���E1�엚{�[ge4qv��Z�*r*�p!���hQ�Q�gg���G��l��.�(d��Ȇ�a.���2�j��G�v���S��.��6v����<�ˣs;��/Ǘ��j�τ���͵x萋��7����H��F���A3������د>�*���~�P;>�f�J�ٔ:��pE��+�{�bw\���c��	_{�k\���w��Q�zk>�j>�o��s}[Y�c7�|�"��R"
K�ڢ�*�_p��ԥ����������jK�5�OK܊ޥ7�)}Q�cs�Fja���ә�wcy��[ڂ���T�0�Ga㝸C��\�c���<�a�s�@ח�G,��z<���Q��FI=\���Q�����~E����]`�8ps���Ũګ��=A������Zzll���2�t���>��UX�.����劸}���Zi����#�׍�I�,�����)T�f�ä�uh�T�y�8�T�\���v{Lҫ<���]�A���k��J��
�$�Ց<#�����
��~;� �u�����˿@tɖ��Sͻ�f�c_ٲ����ã���.ʋ��C�*�#��G��w@pY ��b�Nc�	HM�����H��p����n�%�J�;�����j�<|�.�ͮ��t�tu2���1Y���e� -�=G��蓻�����[��!�J�(.�-�b繮�@&WS´z��'���2��ƽ��v�zy���O�����ܷN�"Y�O���x&6��U��@<%�ȹ����L��s�_F*Y�#�R�Ѷ��eZ��3veW���O>�'C)��9`xU�潸���m��V������x������ܪkG��d�׋<`��$��J��S�۹��R��W�����jpg	�_!���D%q�l�j,��;�<i��"�Wm�ka�>a��ޫ�~����,^ ɫ@��'��#O�j�rn(c��(����)�+�c(D��V^��;9i���Ӹt�^��j�hw�ڽ]�"׎RA���5<�VY���kxYy�=�î�?V��=��N�%���S>�P�^�)R��2�����fO�}t���l.��p��~�;�Jf�~��2�;G�y.�M��!l�u��K�e���c�q=5�|�do�69[�H,C=ޙ���V��O����|-��l�.� ���z�ۇ>�8��f)��]J�sw�����lv�$:7)EE��<Ox�6�f�LQ �e�H�4�x/�����EM�xF�<���ސ�ʺ���]3����N��$Sb@k���g�f����WT��|:-���e�^gj�Џ�>�������&��+K�gp���1�oc�٥�^c3+�)y؇5l(���4�	��d�g6.���y��y-#�[6�ku��#[����]�xt�bg+��`�Kd�3\R��O����3�n��}y~�W~��[>ֈ�Sۜ�Ns����N�x7��u(1H����3���)]=�鼱l̷�ķo�*[P=ڏ�T�<C>R)�<�c8�k�s� ��+��I��s�j��k�V�[3�ӕN�^�\4g�5^��.a���T�[�F����6�O�.�� @=Y���T)���S_e�ۭOu�^�OХZ2�����5�{�\S'�Jl�M�����[$��"4���Rt�,k��qA+3��:|�.�jm R�*{&j^Z�o���;�r/fT��$��t<��cK�]B���2�-��B���K��K��޳�L���JP�V�	�K��,��u_�O:�⪮[�%-^/a�ʹƏa��ݞ[��e�g��M�ϑ쭸4��^q�~'k���!u����u�^�f�'��+�(�4��{9d�窳O
�/v�j�S�5[q�<<�re��`��6_!\�u ����Uߜ�MZua����[�[C�<fu�@5��O�U4К)�c���0�Q�gWY�R���j.�Vp�9�Cj��gD�̣�Ѻ�;�j#�<ל�ɉ$��Ҡf�ް{����Ϛ]�Gn�_�[��!�X,*t;]������4���#L�^�喻	��o���e���[��X��U���A�Bo:_Sf�M+7����3(��_j~Z%	����_e��9���W���W뻘�_�v�K�Z�W�X��Oz	�ē6}{�0���.-�]��n�Q�>Fg�mp8]R됁�y܄�N��V�b�7��f�Z�
ܖ'
��<9���b�2��]�5(�Ua��y��=�߀����t1����P��K���T��A���'=���T�A�^J��	uą�r���蓯#�9��f&�n[\J����ꝄA<�!�S�\�N���c�V�	�`��/Omi�6w#��8D�B�p�k��ä��[��S���|+W�e<+0T	�ɗ��S��k��縍%�B�9��.��	`��+iJ�։i�a���U�Y�%�� �:>Ż��J��xr��*��p�T��_\�у���t�I�_ibo^Z'C���2�[���_[:�'��hn;�����^R�'�&���J�����;}zKCⲛ+&����HY��Y�f�KFu����2���o���7�ZE�gVQ	G+��R�մ��̐;�q�9�S@�1��lS��ԣ<O<Z\m�������b����g'j�w%�)bս���o`��� ��/���]7��rW=]��yn�3��R�1�ͦtzAk������P:/�*�a�/�W�8�W��'Ӻ-Rq��~g�֘X��@o�c��}
��*ޑ�]��0�|��5흊T��u��۳�<�VNhKD1��)"���>�:�-ب��Ε�73�g�Zq�Um<����M�K�7�8�[��i�V2W��>x���̋�m�2�}O�E-�J���c$�y�d��/g��Է�f�`{�h;�9g��᪖UX=�pʘ�����#�b ፌM���nq���º}�t�//��p5�@��d��u��Hb�^5u/V��g$�����wc��Ԥ���`��EOMez5^���wz��R�C���� ���ʋ٦/��*V�]C+��C�z��F=xg�54��Ƞ}�7�4eF-��2ɮ��k�������(z��/�a�o���;��\�'�Ӆ���2�wÖ��s�w����|fW�㤺\t$�vJ�&:>��<s��Osˬ�>7���gmj1
����^����-QO���s��9OU��Kq��fs��rۘUh�7���f�d���uf&=�[Tϰ,c�G\����Ʀ<콡����Jeh�J���s�Aj�`�Hn'��Ӻ%۵��4{�%=z����K	W��&�n3�1�j��.��*�S��2�:��ؙ_&�y�Z��)B�
c�S�{�����nr���4�_��߰�4g+�$hwOPE�h�va:)'�Y֩�y�[��ؼ�wq���J��x/dO	���T(W0x�}e��E��~��
��l�d�,�';zr�\_{�T�h�f��\V}O�ʋ��О��S�
~w�i�W�/��q��JU����t��%�D��fuZ!նY�A��|,�nf���7]���4Sª��c�yS�p���TI�nয়B���Xg� ���rM�u��D���'٨
����&Kb�g�=�}��~n:�<|_����2R���8�3܆޹�l>�j,�_g�	D/.�+��/�wb�K��įJ�O���c��n�ǵS�!��[�(k8�"��P���ѐ�D���y��H�[��HuOfܣ�U�О<�xFW��n�9z;��U��ҩ:v=�9����u�+�Z]���{R�׻y�y�"sK>ݜ&NHa�pK��3�I�J<�Lݹ�Y�M�y���y��#���ą��[�dm=�Ju�~H�K,��TU:�<�n8, �` �(;���3��=ۉ�۷���^�����SS���J��<������zA.��������|�:������t�����a�����UY���I���s�s���\�r���3���E�|�8OV��g�Ђ��>��|.�p�i1�W\OO�F`�W�ؿ{t�'W[����łGe�l��`�Ȁ\`Շ�`��p�Ʀ���r{����0�FN�1c�gApo	��MQeQ<Ox�6پ)D_e�H^wO��7�<Ϫb���<����FO�u���&��0v��k�4ؘ9]��X�%��)��-u�UO°�f�oj�so����2u�c�DOۜʤ�?hڨEFls��y��E}(1^%����!�K��ҭ{�Oo�z�>��#�-���q@�~���<C*��x�}<�fS� U^���f�o��e�� *��Vp���<w�qA�jZ�Gu�{�.a�1@���5N�����O1Ի��V��`���t��
�]
ኧ��qiĆ�&�����~�*Ѡ�e;����]�G��7Ŭ
W޲K�i�x襴�e��/Pfr>#��a2]j9y��[cAv�Y F�mt��M��S[]�3��_@P�1�}��G&��r���W��n��wV@������mh+y;�s��A��\F>i0��MĮu��Iۢ6 Hj�Tu�`�Qk�"TsxKH���u��̽�W�p�����` �r�v%=w�	�3{���ٵ]V@6���*M��x�R�<>ݩV���`�V��G�!yF��Y�1ƴ]��[ދ+��n�άḈz�]R�EkC/ܾ��w"�,���w	O��uw.�^�w8Z�TO`����^
��k�n�_`�+u"G��uܩ�;�We�kwM(eT�7�^-2Բ�*+��N�6�F�KLS�U��G&���ͫj�ۮc�v��oV0�@Q��J�y6���z�Y�G r�g��D�ks�R{w:H{x�d*���j\��Q��o:��0K\4Ju���H:��l�W�L�(rU�w�17hػVug1N�<�]�ūU��9v2*�O1�,�3	�4�x���z��V��!�@���%�v�������M�8�'Z[�@���:8��p���C����u�o���f�ծ��sK��ME���X泖�����9;����tA���[�f�6$3D+`�!Ïk~�W�j(!����%�<V�mp�K&��S��Q��-n^�ژ��X,�w�8.�!�Q�S1�*�@�y����R�&�eN����K�-$�r1
S��]��r⾵�l�ʖ�DІ���m[^u�Q*�NOT'{��}�ܬ̸��jۉ�sZ��Kj�bz+������@l�����}0���CZ�N�{�vDG/�A ����V�N�\�;�5���Xn�|-^	�m�?\��Sr���`�Y(�(�:A�jFX�օ�nwiO�@;2���5��'Q%v6�dB���&��T�4�p�,Q9�tO���
�'�4#ʑ�wo�ݸ~�b|Q�^�|�.^��̸�K�h������(��J��j��aa�jL�\t��h���n�k7+c�B�D�QER���*]���3��f���)�����-q�WΏ#Vͬ]��]�L����7�uo5L+#i������tf�s�E\���l����Y7�Ar;�p��༵��0qu��Wj�-�\��]���n1nf�}E�VJ�ذ)�Gn�3��\x�n�pܑ�oy�e���K��kk�!j������fb��D�ۀF��۵}���{Y��m���z;0Ԑ]Fks��T�m�{6N՝.����]�z�==�Ѻ��Ϟd-L���DƧL뙇�� ��c�ԭb�G��e`ztd��=���H'�v]�"�pG��v;H溲�NcDU�s�[o�(Zhr�]87�{,�Np��\�L��8aG8�K�+f렻���Η�-E'<���c��R̎��EӍ\���C+�m�DV�޺���h<°��*��T��6 ��UKj���VZ[JVڡm�VQ%�m�ikJ�V��Tm����iJ��ж��VR��*(+K`�d����k��U��l�m�%b�*��P��UPZ��Z�JJ�R�UX���EX�mX����F����ֶ�ZJ�V����e-h�(���E%`��db�����TZԭ[`QX(5�T��T�[V��iJ6b��m�jelX�Keeb�j%B�V5�c���eE����F�DUEX�j��k(�����Q�����QPU*R�R�KeR���
�����Z���ZUU�e�+[eB���Z�m���#��Ғ��Kl�-V*�֥�DDk-�ۏ�ˇC��A=�����S�@2S(j�\�-et2�X�q��v���Kvm�c$�[���J�9Ԭ����՜���.˙,��>)���߼R�	��*/fT�z�>������ю7B��@ �Iw2����{r>��^��g�5W��Ay.� 9E�7���NyeO3��j{�um��]��cq=o����.Sm[�ZD�#4��wy:/��<�/��DZ�f�Ϲ�5�:J�)zm�I���n��_X��ר�~��Ln�O�ͳ՟Wj��>�(x*��ƞ���Gn�f���%�2�_�W�J�C�#b��/ey�	������o�%Y�]O�n�}�7��	��3;i����u��=-���hlX���c�����w9��o���6�z  ��j���#� %��8v5��]#y8�M8{O�Eí�xo��h���wꋨ'�� X˨���O�`p�7�2�w�L�5"�eOB��r�ŸGS�3#K�=_x��)�M�ܬ�֚~�à��7��m)lC�7�]p�9���_��z�s� Tx_P���^���F��i�>�b�+!T�*�W������Dϒ9:2����T����O�l����mbK�䶆ߑu����nf�hSc$�c���k�L�iδ���3\O;F�Ep�OV�C(e�+��ZW�����=4LE�=U+C�Ku���X[�gh���Ѱɨ���p��꾧��Ҧ�}8dX�Į�oaR��g������c�{�pO��@��ѮQ�5���%�<X�0/�{�!��)t��Ü8���q�S���F���o�����,�d�b��]5F�z�]�5��Zu�&;A]����s_o�{֯O��5c�Îz�Lٸh',�J������ma6>e{֭V`��<���A]��~���3���#�2e�J^R��&�&�Al������:C�s,���8��t�g�CE1�DLw��m3��\D5�݊�vt�X����qa��ZD�^�O�ݺmr��߃٩��m�IW���RX�ʷ�gD�3
/[�V�W6�3�9�ݓ�zV�f�[+l?Yvm؂%�ʭ:�-ب��Ε�d���1�q_��W�M�<�W9��~�<��4ºW�2�{V=sڽ��c7�+���[B��u{�Nt�m�/�F/W-]���

�z����N�g��Y_X=2>�Z�i�p�&������[������{�H���~��� {�8
f��n��`C�}w�����L01r���-5C�5�I+��{W�]�Yb���r�v��}��*_e�Vm��S�%S]�Ւ�ӫ�ˬVi۵p�7���N� ���;�Ecz�� �˳d�9s���K��;�+[:��tm��6�ƞ��a`��o]o����Ok�7w��'��1jb���b��=o���3N��0iaV��Ы�����.竦ny(��g��!:�V�� �u��ji{�@��o�h�Zv�g�\�v��2v�6��K�f"�P�� �����.p	�D��\󸞟UN�������֓} qy<U��<o�E���U���u�iPw�QѱA�9��a�=�.��^w�f��}�zh+��{���׽��wf8#P]O� ���.]���A�O��,s�4�J�'H��تQn�eR�s�â��u�\�3\a,U�bu��
WX�,��8���%f�{�{f�
bW��x����g��&x/VD���F���P�\��H~=@���rr������9�G�<!��q.��޶��z���3s��ޔ��R�� �}��ً��ڡ��]�Fu�d�fZCt��]Y	ӭ��u��"{�S���VK�4� :e��/#����-���"+p�0kW������a�]�2�*����n�M��پԚT���v`E�[A���T������t� � +nM���j0P���m���LOu��<�q�vaXo]ױ��d�}�i����ڜ�^vI ����h}��H�X�qL٥U��z�˥K�!f&�G)�.bo�lG��u�y���yp.E�+vG���ya�Ы�m۽�tz�ܭ�}5P!�!�Mh�%��Ş07ȓ�0J��ߟw4���X@�CEFkL'8�>�\�p����Y<~vk�|�L,{g��+�4�po�\�绥�τӠ��0�z���OA�KV�vU�{̆6�WPLmb�o*���p~��Ig�J��_�ņ��P�j�{�Y�C�2r�xl�U�z����O�����ګ��f�t8��
�C�`^N���t����+}I��`����_����$}�)~�7ʳ�g[j���� ��C���ΐ����\�/�`�Cl�{׻�y�8J�Y����܊>'��ۖ��`z�u����q�r�o'��uv�yK2�-'E}��1���Htn|���Oa��փ ���.2@mzj�>�:Z}#=~]Y��Mo�?�&��0�]�{�lN*����J��#pd�� ��GW�؎F���{SaX����H��}�ə{y��S��vl�4)U+�xsN��K(��{bpr����/�+֩�y/jX�+���!&^���\˦r���f�ouց�v��<�kLG�݇���G6Dͭ>�i�I�:{Ik^dbT�\�k�G�j�&c�9���xz�d�)"'R�Ẹ�����b)ֱIuf�f��Oށܿ^zi��V.E���e����>U=��"�j��d�b�~�W��U+Y�6������ ��1�Q���8k�x�w�R5^��.a�_��Z�:V���<Z��ڵk�~����^6.�T�%U��W��5��mM��^�����bqm2v�H�r�\��̧~�=�c������޲M�F�7���+�_<9}��
SI���8d�����+(ʡ�`������ȭ����,��T�$�AS�N�Ҕ;�N�c������v#�o`�W�}�d�.� '*�WK��<����W�S�:������k�H2u_����Un�W��|2�|��ۃAU���xP�^��tWu�R�f���
���j�.�+�i��=�_'�ï-9�Ncu��G�7d9\e�'=<��M�u<2���g�E��{�ܷ~=�b���9zfZxOظg�����o�,`��V�q�����;]����n#��a�$�Ի�� ���S6��kI�/Ga,�*\�ڄg޽ ����n,*;�I[�0�u�	_*|[{��ዩvK��{�EؿN�&ŏLEEC!��9����Bo�?S����4��,I���Rc��(g8�M�1Vo_%E>4��q��IwM���iۺX*J�lla�'�w]nt.�ɏ�P�Na<s,�����H��Zi��T��m�x:4R��}g�)n��PPX��9�*�D��uS���m�:�.vT�3rmק59���{�=��]!꿨yo��\��s� �2�p�ns��Δ���V;d�;���E"�eQs��T�s]�=PO|��<,O��6Im�n�W㣝  ��Ċl�Ү�k�^w�};�O>�5̺�-���Z#���D=���W����Ɖ�A�Yd X�ѮQ�5�����ӵC�����wt��u*Ee㓸v}ر`�S{)��lw�1
��`@��t������*k]���fw"��W[���>���w�6����!S����;{�EN&�0���Wa�U�}Yb-yc}X�ײZ���,J�c���E壼�X;��#�2�\
�����H�ԡ6'R��4�۵��̽}�F϶�0*�C�w���k��L��="}^U�I
����.ݳ�OҚX��C~�9g�ޞr����c�^")/y���$62�A�T�[�2� 7��˩�[��t�JV"�HK��mB�b-�V4�;�qN6�ފ�2��'�{�=��ŶB!ĘƮH�aC]�f0"�s֥�^c��h�N�&'�q����,��.HZ>�{;t��=��^��RHl��A�44�u;=��m���^a�s��'g@m߾y��~:��ţ��^��Ek~� j�N���� ��Y�c�����}-^�0�`X�mȄ�c�P��o���y�B3�2�i�5�r�.�Kd붽�uSw9R^���?3���ڎ��j��ߓ;״^o���X�������7��7�_^I�55����d�e���};WYC+�|)+�o�,^��W��w�ӱlٻ4c��c�A�Ͻ�Ќ�Z��nfzEOMez5^佦�n�3y�s��a~�m�ݐ�zt�2�u�*�ܡ�X��p��ja�t���54�Ƞ}��cf���2W�v�l�վ�놺W^������퇉u��g>{�@��peS���������m����O5ܼ/����@�\�Pa�<w�8N�-*�����<pMFq��\�n�s]r����8�c����/��ʝ⫲L����ca]�*��L ���ݧ�ƅN7W��ZY{�V
9�JkWf���P��_�Z�҂r�B����l�y��/E<�̷b���k\��ȇѩu7,z*�W���N*5*;�U����+�j	Nn(�嬧e�}���hܝQ�{�iD�\Pek�NPA�����>�Y���>s�!�{,��B�Y�e�JI��!�-:C |���6�N�G�xw���-��]݉v�s_����ě��ۦvuʏť�Gk�Z�yi����*f/gF���B���V�!\�2v��.�ԝ��P��s�_f�YM�~T"Ι�v��KF��w��G}�3��Ǚ��U�03����y:]�;�S���/���>)R�ߖ�k&�Լ��ٵ�K����U3�"��W�W��/5�dM�z��f	uz��M�)�`E��kl_ӄ�X���o�}���{>S7.H�#�씚��w�z,{����U��0�~Ҷ�3J��=k������C�9���Q82z�gx��������K�Y1����]=���v����>����{ɽ��\<2]�=J�+��{�����g8����q�4���3+����������&��~��y[�+����XS�	��h=�/N�hG�A�v��)Ʀ��#�K��q��x�eK��&��H����q�v��o�P����z�ߛ'�����v�U�#�TB���-i`��Y�%���p0t��m�C0K�0����u$ީkM){kkqP�n���mt:'EZ+�+V9Sde�����;�������)e�]Ε�VΫ���7	^̭p��)_9�v��=�2�������NMܷ����G����W+�NxTO2�����L{�v��o&����&����<�BW����-�}�A���nU��E�!���&ԙ�����ݸv���
Nӑ`���v��Q~�h:�	���jz�s�3#��Ѿ�8�]݋�VS�v��J��-�g�&��렾�N�k�[�����O8}�$}�*ܷnC6V�]�l�I�����n�`��C��:@�j�\ϯ��YM����3h'�ޔy���2kR��:EՕ�yQ�k=E�~�xuH���~̝�T�<�ul��F5N��[R��ɪ^)O �]]�y�So9���̴39郛~�-Rq��3R��`]{�)��U9Oåg�s`�򯰫<�^���[��s����tDު�*�?_{w)�Ŷy1.jnŵ�s��J��+F��̓��\kW?aQM��:�g̚ΡZ%�h��t�u��Rˤ(�kwj>�v��]��l3�K��.�WP�D���O���W.�]�-��s��}!S6S=�U��v��ُ=뛳�kyк�8�����W�tɹ�@fWz�]���Z~�n��
5��K�}�[���zW��bA���LN���w�έ�l�5_�Q=�qA�y�3jQYsݪx_�d���d����sI����w�[��yF_�����	��}mAO6����xb�B����u�%[����3\{���mɾ/1�ҽ���/|�onD�#�X���4Gj�S~b�G�ru>ٿ3'�v������S�X�x
>G����(»͔N5W�֜Y͇�����扛ӛ�zտ�~�M���[�P���n�N�W/�|/~Ϟ�<��s�~鹘�d�.xI6[l���~ᝅ��.�JaSްC�[N�ꃻ�}^���מ�va5	(���j��%"��LʮdE�t�����*�s5��	!I��B�����$��	!IHIO�!$ I?̄��$��	!I��IO�HIO��$����$��$$�	'HIL�$��	!I�$$�	'�!$ I?�	!I�d$�	'���$��!$ I7!$ I?�b��L���L���"� � ����{ϻ ���©}�O�� ��A��� PP4(�B�mTրU�4 &Ɗ$�77%�T�cC5�m5��f��V�L�E�Z�m��kj�ڬ�͍U����Vm�ϳ���g�eX��jJ��$[kT�*I���2l�X�h&ѵ�Zck1���m*6�ʽ�](5p >�P y�N��sPtS�c@ij4��u�:SM��@E�,�hI��Δ��5�fjT��6��� <綐�Ц+mն� ���t� ���┠���S6	 �F�[m�i&� �    6    -�    ;�  �y�۲�:���7`�Og��U1��E;]�7[l�[5���l�� �����ॳL�Ъ(�� �e�k]�V�v��i��:��\�N�卭�FKZ[k�w��{u΀wg@��n���� n�(�4��֩l�mS� �)훌 ��GuwR�]wte�ֈ� T�(@i��4�ӋC"IP� ��F� 7s�, �`�nu�b�Z�(��'u�6�۪4��ڻf2׀x%��v�t��	���ٗN��s��Pu��@sq͘w	u6M�V�����颼�K��W:2��۸5��[��;��:�YA՝��umY�Ym�l6��< �����n�i�l6��8�ƺ-u`��k�GCT���%(T�� E7�©JPF�F���a��1JR���i�#!���J�L�i�&&��`  ф��?�%	�`�@`� � $�<��&Q�'���i�� 4b	4��)��)�z�<S&Q�hh�M�l�mṽ�UӅm�u���y�Ͳ�GZWu�M;zK�μ�O?L	$�1���0��	$ ���%	5	$�O�I $!?���7�_��?���H�!&����%C�d�I$�Ԓ��$P��$��������]MÎ�~v@���`V�"T��p(��dyc��U�  ����"#Y���%^��2��"�Ɏ�;�s"��]I5�Ĕ��:��J@��<c5��Z;X�9"���%��gM�����)ݼ�G��
�KVZLS����K�B�Ww�)Yt᧿gQ�4�x3Y�QT�of!���f�TDKʛ+N���:�^�<UCD���B.�V�ń䶤Wf�fT��*�ʴYr˒��kQf�[T�٘���v��Wn=li�{koNf7B]�v�R��1�z�3`�X��o1M.���k�˵s-��?�H�,d1n�"]Z�X7�a�b�� b���V,Z��2��F���=m��ϱ�vY��f��t�e��b<�wX�Z���$s4T)��	X��N�hL����C��~.ᐸ�ym�,bL�G�yq^>�%k�w���Ǒ�ݼ� �,���7�ի.�Y�!іIYwF�Dk`Q��H���mf��m�,҉[�u+o���[ �qE�h/l%�J�G �o,H�s(�����si1�;�P+��/K�-Ù6��O�˼	eHMU@����G-�-���}�X���5}ZDJ3`�l=�:r��y�
;�]���e6e-@�䐜����,��FÏPd=9X���37ܩZ��0�HڸshU�C���8��?��[b��dU,q�Dފ�Q�;�5�c����f�u�56������)˕+j[��:�#��:d��BN�iA�ZI2��F���i�a�w��5�Ȭ�E�+<���P'��Z!i�Ӏ���u�.���4݆f\4�z��2��M�͙WS0������ȣ5Wn��-���eI���ȩF3v��.�V
���mu��-��2�/u=�A�VFvh���hAb;f��]c����EsE�4Q�X���Y��0�'�|5�VOZ ��}F��8iodT�a�TPy2n���U0�2A��7�)�'4b��x���"1�Wn����6�Hܼ��:�aXbm�d<	;�N��GU�̋ܚE�"����nm���$^�DVeU�2^Z�5Z}��L<Ԭ�����t�VK5�m��ᬰ�ǰ<7+t���^�&�J)�1�U�56͗��V*
��Jn��TZ����*����j�4���s'���`�'�D!�nɡ�^Xc+6��[���iS愈�.F�e�
��lod�	u�ef�$�c&���<�P�����̽K{�j��^�QTz���\�*�!W��6�;��+�v��6e[�ZəAlh����1f�]�EY�*��>�X��0Ճ�
ʴ^��-n</L
����*�5��;�/-d�f���^�#�t�E27���įR�PT��^�ص�Sz�^Ǵ�aʥj�l���m�L�ٮ�Br�d����yӡ��[qѷPKED�*r�ұpf�NEXM
{�pqzE=x�kw�K��R��]ڳ��ڔ*���j�-V�	.�Z^�W��&т���v��jSke��Puv��͊�j�ى�F�b}� 5_n+���D��cB��T���v�JF�����e	bk��P�c�t��U��\�i�B5R�[��ZN�����۬�j�$��ha���,&MI��]�539U�c�K%l�!��Ci˖�S��ֽ��h�8�e-��	���;�)�ίww3G�'�����wY�xpƪam⡭��f6Y� ��{ψ���gl�Y�K]�]�,1��2��76-�Y��>WCe��*�SІ���x��Wx��xZ�O2^�Xi�YN�1H�y�jm�ċ�n�
m��n��6Ł����j�m����޲^#8���V�sL-�*���a�kt����_^�ocE���­�9PK-KC^Ь"�5U4풗�2�,����@u]�<�d�EieMO�6d�N�%�U�;��V[�X�R�MEQGW�X$H��p�h��靣�n�Լ��Z�zڻ7R�aҠ,��ܲ�.j�#k9�o��ԩ�u��l"SOF]u�@��#pn�+�W1�PzQH2��wxH���+�ر��r�7zAd���Ӧ�l�&Jن�+s2�`��b��BZhi:�]�
���z�j�h�I!x��F�k��Z�[z����ei[��Eef������nI���	J�%s.�r��X�De밍�c/!�b1��	mR43z�R����V�ݍ��r�BueG+(a��;j�.�Ml�M�"��pc��ۉMݻ�j=���j�m��{��=�c+���/us��eHn(���
���u�+�ݹxR��e%�I �L&�)b��H��X�*�w�kV�hՙq]ۙ�.b���N��]&�"�
l8��6}.�A���)��k�,ǇW_�N�i[z̽ȴ�D�
�s-+^�
v�f�4���߉t�w�,���3`n��+VҧX��x�w�7E�Z��%�hޑ�!���K���K1���7&v��4ȣ�WxC��J�R�u�.�;�
u�3YH5|q�Ya�AqV����Y�n�2�qa9m+-wB���5�W�Yb_�4�u���d�skVk��.�+���u���ж����@���5Zq�ۤEeT"���Ut��M�8��T.��ׄ�zm�\�'+�F�ҩV�܎�4�f�դ��j/�+i���,��R��V���
���nVDn��4���׷TV�B�Jn�8��H�+�.�j�m�]C�#�Mf:M�MX0�yceų)=�B�3�z��0�f0�k�w��m��Nª�W.��;��s^�(;H�r'/%�SLr��.-�[�5ՋVuf�Ө�n�7ἲ�1��@�3�3,���g*"�&�v+q�_C�f��g�q�wbJ���w�"��f!�uۖ�]B�5ï��hD\���dB��5�Ҧb*�-��ǥ!��W��@��B�S�,���re42�o��t��Ou���K�f�0�����5ۇ*��:���ݫR"�<��V�j���ա��nT`�M�'J���յx)�F��h �;�z��]�8ۻ��t
S*�����m�q���D���H���5�J��vj��(�U�Y��L��I*�+��Yg/eSE��d̡��Jj��qY2�ٵgoY�X�i��x��X��׶�b�JC���7�ڱ�T�1'uP$kfؤ3D�H�+�8��:F���DkVHP��:(P9o]M�Z��H��/j��u-�f����-Q͏��_ML)��R��|��EɁ�ͫˑ���T��:���j�Q�N��ʻ�c�Oj�o6�`dJ4Ѻ�z�E�1�n�gֆ�H��i��o�)K볶���S�ȶ\��W���GH��J�]�Yjl7r�5�ĺ�Q��m���%-�Ez���'��r�ݼ���ejt�Hg܂j��r��a9��v�!�V���,��;,^CS�/"�ϊ�����![i���N�"�P�W��6�f {�L)�9������f(B��]�p�+����T�tk�
٢��U���.]�کt��+*�B�ˁ�@F�xec�;�^4�h�x�TF��wS-A���D��Aæ�a������{v�<������a[���fS�*�s.
Ѩ��MU����s.�����1�-�%ʣWNnR&��v��5mS�6�zeũ�[��t�@bZ	���7L�Y/K���¬GW^+a��u�r�/������b�jZ��S�ZS[�'�t��C6`cMd�V�m���5BX���)����L�g,��y[7�w6�Y?u�"6�VZ����͌�"��t��$ٷ*��!�U��7xu[�7�eV��F���
;[{�YrSܼ��Z���E�D`f��"��3	�.�z��w�&j��t����[E��jQ(���u�c��*�H�0@U�aɊ���n��XKT����VRו�m�Ky�P��]��|�!o��h��YRw���r�j]75�����(eF&l5:��A�d��CBfdZՔ�9���qkfWI�ј�7yW��hಪ
OI��^hw*\K��J���]\&����T�<ډ�2���Hl]is�칷p���*cԕ0I$�Y׷*�&��o{��B�\8h����p�ک]p[.�؊��Tx��SP\=����a�<Dp�!շJ#�}���:����
v���.I]�<G^���*�<�§��V�N��K���$;f�o`;G���r��U5��a���U0�h���B�8`)5[V3N�lYzV�r�uF���n��wԲi<-�c�'�B���o��Ŏ(R�%n�мҰ�_lIa]�f�j����k�7���ö�+�}u�*��{|����zL��Q�2�^��<5l�f_>��ې(�O�v`�x�u�N��*K�-Fb�Y�A��!�x�4�.�k��6�r� �E��ua#Tqi����w�ݧ�h��Ձ��H�G~���-�kvnX����n.�3��X̬.�#�G^n)�@5�3����We���+���W�V�>�|�K��������	���pq��ĳ�f�o�b8U��feըu��&�U��]��"iaa�'�a�b�*'Qf��-�c[��̣�����ؑ�\7C���H�����ż��Q��X�ϜJ��}k5t�$�BO%���[��b�| ����0U����m�>�sk��Vf���o�����1^��)����H��ד"�5���7����V�Y٧�JwH� ����n��ݡV:�.�,�-�G��.l�N��}��S�-f���RCާ�K]*YvR7�����}i��/�sUj;�D���#/%Lvk�0��`UEѴ�z[�F0�h	��Du�W��:�;��+1p/���ޓv��1ŷ��8�"�-�b�[�pz@�9tms|;
m=�C�F�m�QoJC �sw[�u�����%JO�W�`!mN�iǛ��vv	Q:�V����Z�2��6�j��z�GY
�S1��z�]X�h�h�l��d�_F���q�fu���@X1�c�3|��5��ys�8+�hۋd�6�����2n��%��/dI�s��T�`��n�&*��9u�&���m���D0\GM�V�ѧ�4�p^�|Z�A��3"���Vv�"�#)�2�0�,��m�*K���\�T�f�+F�����v�P-'۔���΄�n�^YBnĩ��Z3;%I��o���di�ڦn"vhCw3m��b����~:$�p�GB�Y-��1+�f�W�ǈw�Z;"��Syt\�T�(�׎Q�]c�ajo��w~C.iGwYTw�suh���u�lV!0-xۗ���^T�R�2U���ilV����G���,���aL������#rV��Kv+���!�f�T.�gM�I����4�#:�Ym���9Z��ooA<U�]�VE�Vr�S&��)��;�[���y�9�����z�d���:�I�������sn�5�q��ubz�wHA"�`��7��}L,x������+Y��xn8}[��!�Y�5�|	�v���젩��Xl�B�?�<�Oz�ǫ
�ؖ*�R���eu����ڴdq�Cs#��	��0�b�c��i>[ZG�����KV�q�sW'���JK�E3�d�n�K�c��$�V�P��YRD��es*ͰE��
KS��M�͹+
9ٚ��]�,A�;�l��j��ͳ�d�y��������CL�cٌ��j�wN���Bp�Ўr�j���`M]i��5Wm�D���t`:��]�[!و�_J7w&N��i!0gR������,�_9Vj0�i+�;c2��f�|�s���]ܛ����:J�/X��� ��������vl��ﺕh�:��!]2�L��I%�d�j��)�x�s���)e�,�Xx�y��*��0�P�G-śGq�V(Juۅ-ی�0�5%�����8:���#�����극�--h��Tm�͋:ě�u���L�M�9˻�[m�5%�f�Oh�fo^��5�x�e1�-|켋�9m�oOj[U�[�;���QvV�
�X�KN�KrQ�{�iG�k��MggMq)�!zs%�ap���9���Uk���ڊ��Ữ䖭��;!pL7��*��-!-g�+A�tT�iG&��s��=w&�����޹�+s�+k5⋹i}yۉ���ge1K���:nZ]�5i79 ,�z�:�b��-�je-D\2��,�uE엺��ܨӫ5ō1�<��0r�d��V�u�8U��M[ȷ����a����/ᨎ��U�ɑ7r��TN��6. -�p�1�io��śzs�85�(��
q�Y�ot��.�0��,�OP�u�t&guZH��ѥ@ڗ[�h�L�D�0�ʦ��i�3me��U.�z�Ӯ�9��������h�cd_��fG)��AV���\��e�2��v+.�9n͠�bN	[P=��^��F416�Įni�]W֐�'S�\J�<���dx��҆tbe�)�B�w9�[�ҝoK�6nƱvI�]v���(z��sNq鉪i˳�-;�c�=.���N�V�U�0����!Y��\p��T؅�y�4f��	1N���A��]S�z#1��\�vr.�nM7��F�����*�Ftoz�����*«��u��.�5�(���d8ꭐ�=:k3^��خ�]U�n�(���7r��`ًc,��'b�_N���q7�h�{z��Q�Ӥ�ӹ���^����I͝�0���}u�v�*��96,S���ݜB���4ic�z�����Rń�U�*���Y.�O�J��RK��]\��E����k��EV�|�so�J��Z,,�oV7*���H��ɘ0W	��]&j>�ζL̏i����c�Ӌ�ڮ���6#N]c�j��b7N%/6�L�68)'��s5(�4��� ��ێ�:��xT.m�Y�N�s>�f�-x�dt����KD!]�#Fc���>��G��Q���y1��كָ�j��$α-iX�`c~t�7�f�7��tc=S�)᥺Ը*�(�����-�S���⋳+�j����������WolU����^bȝNŋu��ԲN�ZP2,�.���7�T��m����c.q��2�ɣg�����H}�e`ً[ݘ��N�t�x�ף�,тwC�.��1�.��t�6[DK�:cF�9O�Q�n4��.�ҥU���iԻ�v��a�=.�`KkR���P���Z�EG{�w�&���(.+Ň�^����۶�gz�E+�p�]���ڕ(/*K&cr#�v}i�P��=�Q:g���`�˺�%��5fε%1	B��V���j�c]Ȏ�em[M+Xr���uf�=JuM��"f@�)�eh��2e�{ڌ8�b�\���15B���o��Rje�V���$[�@�ł^�����_/�}�GJ츃9���W���ϫ��"�ǰ�x��#��W�K��Y�em���f�!�N��eNE��0�.�p�3�G2��LWx��rk���ae/��Z�u�Yu�neI��Y�W.L�ka��G��������#���Z��K�oLl����*b&�dƱͺ=:������n�ev�wOz��ނk�FRf��̙N�4�ܥZ�+^]�nh�8�svp�6<`Tm�R_\."���b��N53 �Z����ƹ�R�nnP�]�;�-���љ2+���P۾�4�\6�͑E(n�Jl�����H䑶�m��m��m��m��m��m�"�$�����)(��["r)�R��ؔ*�wK�˽a����6�Y*�o]>�_wLgs������4F<Cg|t,Н'*��D^�<��t]!�w���yh8�M{vn�\�b]{JSئ>�3*nw�E��q�zkp꼗�$�wS��#���M�"����a�L}9�I;Tdh5]A��Z�K�o����w��ם������ٷ�f��}G���B�7�Y��@��}߸����		!��0��v�)I)��>�D�+V6e)�����&��(��i���!X_*ٲ��<n����s���=����:șZQ���U[�v�e������+-�dj�2wӰ�.�54Q�9�8��R�S��Mou��LZ'W��5�GH\�M��|4jV=�:B�u7Oq�j���G۹�>z��gpD:�J��]��ȗy�.Ⱥ�ἷ]��$���`q9¥G)F���G����< ���E�_M�.VWP���3_[k�wEZ{r3y`i�<j��Y��#��y,{b3��^Cj�e���8R�l��[���Ђk�Ds�RZ����w+��w���+�AX�ɮqҫa֮k�=G��t%VKL�2�[r�7�N�#���%V�"�e�i�|�X&��$����iV�G�)%G&�ۡ׏�n.<Ŗ5��+
�8�a�U�5���^b�m1�.�x).�}	K�:Uu��cn��#qv��q�yiEA�,ʕ��&*-U�ж�m,iF�R62������&��7���k<��X�[�]��U�Ѭ�� �<�h]��}N7��fś.�:r,���!b�K��t(�o���Q`�:���=T���$�]H*�7�v�8�C䊪T��� �khqÁp�t,�9G�R�����te�]!ڭa(�������nnH�8O4{J=l���Z�8��8v5�I	YֲHn��^ë9dM�U([Z2`�Ku������<ڷ}����v��_+��o��]y��G�k!Lku;*�x-�{�_1��)C�,��� {^+�@Vq\��-�+�rc��ͽ$Px�g���2*5��)ge\�[{4����0�TD�X��e�V#��q�f�ٯ�]=8\|+�v�@���d+j���r:6Cq���:�Ҫ`�����,L�5�,��HfC�����fQ��E�0~t/��tU^@�0a��tc2�[�k���fɥ(�D�鯛g�Xj�]�<dn���=[dGF;~/��\;���Q�Q�� �����pV�p�Q��.�����7�u�<UK�^J��B�n�*���jIt�u�v��*�r$��m���>�u�m�R��N��3��l�Z�׹��V!Z2k�DX�G�����-E��U����Rl����g�P�7�Q�K\�5%=n�O*1M<����VԻ{ʛ2e3wcF+SQG��%X��5���8[4ЉӶ)ϡ�t�]���]��w������i-x'j���wm�B�� J (�Ԅ�39��ҁ�Zި��%����c�n�&/�S!���F�_t*.�7��4��W�b�= �t�v��ov�C�fÚ���4���9���u��SxΓ�mL�)��w�1;���2ݡ�ٹ�#
����s>�����uq�K�ءjß.�[k�m�{LnG�7{vn��ۘ�9u�P�ژ��iB62��:��k�
@�41z���lN�v����""��u�3a��/wf��5x�F1��ަ��U�R7#9�ׄ`�YP����MC]3�d�w�.�31K���B�1iKF��q ��k��{��]-�����Ƥ��S9X(M�j5��A]��c�"�v�+W!|�l��]����K�˟fd��t)NiKOrP[2��3����[��d�SV��V���/uh�vk_TV��n��7���d�w31��p��)�.L熯i�*7b-���ͫ���>+i]�N*IU�!s�"��Tk߯E�;b�r�[!L6mq�ېV9�#MP|��Yo�NP���!-�>�}wt�h�0�7��9ٸ�>���j�B�B�W���Т��R�f�[���C+�\����Eb�V�q��2�jb��ս��h�i�)��i�gH{W��I�D����)#�6�����n�l%����g�
fumw���,E��hj��V*�+�g��uz)R��N�݅[�Zг��aY�Z�f0��P��˱���� ''�2����]ZN����geks��AJ��'�k��t�%f,�)ݢ<A���@�%2f�ᇷb�]���gr�Ԏ���a7��[gP��)Q�3eV�)ٹ�wA��Ӭ�xSqs�1Z����!]��ӂw!j�	�7idw.b5�lH�qٳ�ֲ�Ђ�	�p-+i�\77�-uIBVgc~"AZ�ܙT�M�ʭ�<�xs�V�&i�:�2h�]3(��:��l��5�r���S�u�2�4�EUG1)���4d��;��<���fv;�+z��D��mc�8r;��M���5i�z�cZF�̜Mf]9��l�l��WYUp���a�tNTp3�e��1���s��2��2�20�9��k��\��xX �pb����g6��j�x�D���"�^��*mk&B��
k�'G^oA���s��4sC�˒�U�c�l�J6����)�魻} p�Z;N��4H���X0;�k�a����o8��;_m�hƃF��*��2 �C�	۷P3K��J�I���j��t�u!�T�V]ɜ�����.�c$�7f�Xm��Z��`�k^����{Wզh�)`Qǔf���Z��&l������˭�]-��YT�:���\����(�c��T�8�����y���PXW���J�-��F�p2�17�:�m5���`�
.ʀ���;t��[E���/��[��؃,�q/�Y�'!BH�A��C�ZE^�;XJ�� cxxJ���ST���X�,Ez�h�R��>͵�v�@H�
8+��]P̤>��5��[��h"����p��h�z��E�<�h��� C��SW��]CfkVJn�N��p���:6�b�R�u֒�h�A5�T]R�F�E�.���S_Cc�!ͻ�1�ɣ��+-�t������5��JUq�\8�N7f,����q5eb�w���ҫ��3@�.��t5`�M�u"/�1�k/��_K�b麉�w�k��G3�0.$.��)!}Kh���D+N$��鉳p�¾c��h��żf�mn�
L�fX��U�n�Dpa�\� ���S.�M��:��{Q��Z�ot-N��]$3�X���Fq��^"[Y�1�Y�����1��d�ַ�Z�U�j��J�f	󥝊�DQ���Yc_(9W0k�&��G~N0��,�;1�0A�J[&(󸩷,B�Z	�H�6;7��#A�tt�p�(�1Į6ӵ��^������Hⴲ��j&b��̴���G�Ь���-�3�jP˺uo6��2�4�G1QZ���%_6C�2�c�^�ۙ�v�Ą쥭A`��l�tp�kgb�Ė+=��]���qQ2^�m�w���=(��<!ZC���(\�K�R���ҳ$�h���P"ܤ�8~�"�p'x�jUB&��w�u�DmJ�)е���%L+�)���)Ch�UΪ+��C��E�rY�$�W���vi�;#��ܫ�����O�:3u\�BWY֑ܦIk[F��쮶�����l�gMn�wښ2|w&($6)3ve��e��B�O_=��� ���V�7��۪)���(oL�y�0�YY"	��-u���]*z��SV����2 �"v��f�W>Si-7�RG\RfeuͭJ��s%')ѺR�<�4!����B�
*�ַ3�f�jμm�]F(c�G�������2�z"�V<��L���Cv��R��᱖�4���oRP:8�R��Z�r��t�x-wCnZ�������7Sq���p��b��8�쫶U
�3.8���e��ɘud=��f|�©���z�S�h.Ƶ�2����gs��!���	���|��Y�uc���x!Y�aӼ�SB74�-�+��F��42�]�����s�I:�!������A��74�]�Wc��wn9kn��[��(�����N��v�XW.Fn�d:f��tk^��$�d_���2Cۼ�������}����
�
���h��އK4h�tv��R��eb�L�����nl�sG#2FRw�J���ݱl�腱���}�������b�&|����]�;:����<��N��Z2�&�)���V��,sX�uT�b[NA�c���[1��$FF	Lk��;fB��(��|�_=�pjSL��(0w��5��02�䫯�q\�B������u-Y�{��"��������h���5���k�����iv���j��`��42�&�V��5�P�U멮c(��i�vrU��қ�=���J)����4���$��'#ʷ)�ΰHi'X��Ωo��iKʝ�(��U�C�gj��ӷ9{�[�� k�`��c)#B����)ڎF�ycy9$��s�7]��ޱr^jV��,�4��((;J
Ī�J�b1AY��I��,+�+4�f9�+ Ts#Մ�:��5��6ֲf`�U�f�
LIXXTX1Z��LB�R��ɉR[B�)
��UB�i�q��Λ���TWVQ0˂6�km�J,���ci�dS��E$0E�YP�(ʘ�rѶ�"�%dmF�Y�VbE��$�¥B�Ԃ�i
������
����\[�S)Xm�RUE�q�-T�+�&1Ao��T �K�����,֮ɳ�ֽmw��2R�EZL�Oj��Ӑ���[�{9��������?���a�Ls>�������~�o��+�O��r�i�mo��_ -x�΁<"�����u��+�Q�ْ��ٻv<Yt�>��S�����C���q
����F��7�|0�ր��s��(��Ǘ��5�6�JϏɝV=���ޔ��"E�O�F�~\ra�,�Lf������,6��|��P��-�y�k��x�,j�~!̧�%Rʗy�f������#�ʅ�cǊ�V;��[�������;?Q'�fcV�c�yY?X�M���r��L����A�q`��p���҇/���C���w{/n������0��O�ŤP�򵔁5�;�̵���7T&/���L��<�nх�R���Q9}N<�^@s�vn����ݏ8��W%u��4V��m[���Ӯ���V��Ʒ�E���yY�6Gv�wF��e�b�!�"�Kz�7��;�kԼ]/�1�^٦��w��˦p<�蟝�r�3`XY���<��3���s���i���\����Џ��X����o�by�9T��}��>�0��{Ԧ��x�'�"yՄPJ�a/���)|���]n��
(��S����*z�����x�G������G�U��ڨ�/����Ѹ�#�Y��q�-�?o��h����� ������;��!��긻���G��{��v||�{�-_T[��r�X~o��ǁ�y(=�� �ԾD^zD���+4G��hGיn}���kBf����jIj��Z��cv9�^a/7l��u�7U�8�tG,��V��GY��<�����%�O��y��ɗȌE�wfc������֝,����5�[B�@�V;^��f/6n���K,;�v�x�?QM	Bc?W�}���f��Op{̛>0r��а�D�lQ��	<K`�+��p?d� 0�ab�&x����N�:mk�Z���{���$o��c����p�`Wk��~Cv��\y ��&]S�'���|���G�� +�����}Y���mx�#Z�"H#v<��KƏޯ���[|��+�����#�a�Nb�څ�fbg�5O�|+p(nMP[2L�T�>�7�T�����?H�[����:�ow�x�!�O�c����8t�!e����q�A޸}Kpf�{�d��f�+7J��H�G��vͽ���x�m�� vwk�8-�nA��v�=�`�r魜�"˱.��⇛,�f�i}�Ǡ��L_TO�CK��?����4�Rxz��m߶�0��A/��e:b�ٰ#Dq�ȭ�Nf��f/@�n/`��Uһн��c���%�
#�]��+����k?W!9���a��h�|�{s��Y;����_r���vb�(j���څb��'�����˽���<a?i����:ӧ����ӎ�'��!�fo�����u>]���g���x���/������jő�gr�}�E;��9��?�!�H�x}�r�w��J��,�ۺD;B$;ˌ1�����Y�fBn��ٞ�~�=^#ֆ���	}�ֱ���υz�WJLהb_]�t�[G+x�C!���XnU��f�|�A���:�f�zf��n{�]�[�5�N�+�����'-�K�Ȗ=\S��/�/�������o�l�F����D������)U1�j�^ut��>���f�Ŧ�����|N�!㾛DHӣQsB�� ���=��dbl��Q�H�+�c
͟a�c�Vw�X&���Ef�Z��|��o��C��x��I/s�|�*!%��ט��n�s��}D|����I��S� �
�����C=�_ 9�}�vngwu�c;�3da�,�yw)�}D4�ZD(|����p�!xJ�a;�]K�4=h�͂���zy!H�p����g����'���D�0��ھ憐������;6M�g��}Ò:��<�[��?`<x5�͞Nr��Í�7U�O:XGW_f9�����]����i�$b.���{bX�iU��J����L���(qH�����;U|�bkaI�����3���%�Ǘ���ځ���.��[ޯ#�@���-��(��.�����Up��ʶ��a��+�{х��_!��X�XF����>|u۩]^���ZX=�B�ҽ�O�b�b�+�(�X�i߂��G�<7^�d"\t#����&!�j��4Bmִk9�oo+��<6س�A��K������6X�����SZo�j�����hqb/��B��^#;9�~e�=�����'1���
4Q���.�
�:�>e.��=h�fv����ܧ!z� MO�����g/��c�V�yչ�3��FyQ�8�0��?����r�p��m��УM�%�[kC�7V[)�07��	A��ļ��gM�z�;�uae��Һ">��d=eV��&�i7Ҹ�����v�,r�jK�8��RƉ~�����Y�v�ty] @4���y~�x�=k�K�����Hm 3���N
����uW��Ȥp_�n{0�1/j�����`���Ǜ�ο8^W�����V��_}�s��|`Ь�Hqc�QI��z�;�e�CK��=bʥ���� �ˎ���ۙ�͓��E�X���9?YM	�P�;�cD�K��]�T~���65V��_qz$�B�Q���}U���ݯ=.a��ǅ���.�f_i� �M_
�;������ѣ�ǆ�Z��ǈ��M�c}]�aZ�t��4�י���av��V]���6���g9Q���{�Mc/�uB�\+c���W}�3]�_���էO�S�lk.Ҭ#�7a*�z��d�]�f���n+����n�Y���鶸
Y{g�K�f]�v�ϸ���#�cDhC�6�f�x�K�g�/=���vqN�,,�?�*?x�"�/�L��*\�2�D�����=�������Z�p�6ly?H�[}0�������k��!EyLCԾ�bӄYU���<�x�{;y�0�8t߫��&?�Pz��!]ek��B����zp���l����/��e�u��������Yy;�G���~�/���P�G�>�>�����k�����n�qd��^Rr�d4"��B!��h�H>P{����x�������q�}�@����>(���+?y`~����	menn���Y��(��>a�|�Pӧ�>/�K��Gp��nv�渊���,h����j�MCyF[��/�E�a�9=V8*�vڀ�ti�ӕ������\!�V��$X�ѵ�a��Ik�y,/�>�-��3���<}���ñy�Gv��i㇭Qę�/�??�,�f�]쪗�ŅnO�����D��d���$6��т����~t�Ⲟ̕N�����!��,\F���~�>�a�����fߩ��ՙ��V���3�y�����}�c�a���d��R�|���{�:�H���ϱ
�yjݟ}:�@^aG��zߩ_���*.?C���>�&<Ebk�bDyeq9ds~��<V!����4�>�1������}�򂏲A��2-{[{���*!|���g?ki�W�: ��}���~��~�P<_�m ����3�'�0"������
��H��ǒ�Q&�G۶��9�eY�5��ul-�)��9f�3��3�7�;oR�:��d	�X��87;_!% oZ�x�3Bۚ.Bz�j���g�����>"VF�ܸ���m�W�3���/�U��!��h>�R��?}�O]!H�p���aŋ��/���H�Λ_qG��s��o●��]��sR8{��F�.":b�Ӻ�y��.������^���p������OΏ�ք:��������I�C'�w�7{�0X�,?uO��?C@�Њ��Լ�&�ܫR��;������7u=��D/t�_�K=i�%�������k>(�2!~c�Z���s���#�1V��oѕ<�U�/Ǐ��ho��GF�cXǮΞ�HE]u���yQ%�B�iۦy��ԧ5�t�=�}������k�����'f��=��v\י�<mT7�#��3[��j��<f�u^]HN��V�L}�W��I���n�p�k�n7��v�C;�S*�X�>]�2KhYq��\�(���j&>o+ms�P��7�[(IS0ը{2k���rpǑ6x+D͖�+R��i�!������̒Z2�z�$�����z��g'����'g`Y�;ȳ��N�˪ۖ.ElBY��ǌ3���k�w�us\#�w7����cu�2���\s����8���Lh[}�h8��povݫۑŎ�A�"����^Xr�/q�nb�:�g"�Q�Sb����_��Vh̖�Ѓ���0�I��<[2k�p�~ޚ�=t.�o�Ӄ���[i�iaȯw����k��͔�2N��̴�8��q�Z�픱�F*�����4X��U����$��[�e'ck���G��-���$�fa����'i��7Ej*�Wڏ�q;�ZT�I6f���7X���ڤe�TJ�v���~�B�����y{K/[�er�(P�\5`�[Nl���l٘�m@��J�k�ڱ��|��ش���2��Yv�6��QV�J3��,1{Љ�/��x��K��_[���fp��%9H�Ā�bל���ɖ��2��r؋3+�e�n�MK�l��.�"����W��kv�s{'�i�`Fo^k%4﫝ZЭ#�z���9���kf�6�W1�3ln:� �w_ɓ3	2	�6nd�vS��@��c�'�sc�o~�ݮ��YbK�[-���G�;��}�ү ������떢/{Ej[�t�v�۠�ote�;R=�ܙ`�q�7��6F��Z73s��O��!��~�����`�`�Z2�j$�Le`��P(�4J���b����i�-r���AT��KK��X�Y&&V��j2��P���*9j�ʕ�PYPu���.�5�T�%�h��֑V,��3,�Z�b�6�TĨ��q%c�k
²�R*��bAaXR�M2�*����J�+D�(�X����J�*UUZ[�tܨ1��c�m�2��Uưb���Eb�[�L5�J�ʊ)YX�*
J�mm��E�����d�VAJ�UekD
���JY������ǿ������z���R˒9Z;��t�!+x��Ew���`�O�����W�������m44����U��^#q ���sjd^"�65}�I�	a���!�짶����g��Iˬ��xSC�|��
LF+��U�<��b�~�����Vf�Q���������5"�B��V$<Q~�\̙�;����`����۽g��^^DZ�Ъw�R�;Y3���`��}��5�bCk�`{����pb��ޗ��di��%G�K����z���+hW(��j��7�}��,� f,>���~zC�|t7Hqs4b���=�GZ�A������eR��?�k����Ӿ�%��x��W$��#/��B������K�F��
7P=�E�W�Y1L�#n4��ڛX����3��]��u;�K}:����&od��Gv?����;W�E<�ގ��sX�wC#˟u��B_�ؿRk��_�ˠ������z �&*��w�*Ց���(44��(� �}��欎vza#��R�H�[�?�"��4:��]�s��&�7;�����@x�T����o�V����:���-��(��=�jv��+����6�ft��oJE5��c=�>�U�Q��P$2���13��ޱ�������� ��YH
_u�><l�4tyk萄]i��Ù��~>~���?��ڄ��V!Ծ�l�CK�S��_����4(�Xzy���1�R����Ѭ�Ll��a��� ��ƊK�"�tŘ==j�c��G�o2�^v*��V�/>M��	�اv�%>�#��:_t���yю��ow��%4�nN���~|��ʲv#�yҌ�**%@�O#��%;�
��_��+����L����t1Y��|p�<=qbT�O{�/���(��b���W�N��p��"��Ol��Ly����=LF0��.c�����q�/�Y��.!�ǌP]�+¬VeKʁ�e�-�P+��(icW���ˬ.���ok}�t#�x%E�_���=4Q�B������c<�κ���<�F��4}a�kW���Q���[
��}n�{�!'JI�{��Y���AZ�Ck�0T���V�V��پ��h��ۻ �8��9hiX���������7{u�@߼Ǎ��7��bz��(�_n *,>�{Q>�+?��f�G��9o��C|����
��[�߱ڿ�����<5o����6�{a~>ad
�U��"���lY�'�d �{��.to��b��u��z۩}4����Êl��I�&���kg�f/QA���^!u�6t�"�)N�)��m�Õw��@��뮸����7��o�ϷM�5�އ���m���ǒ��C��~xg�l�?&����^��cHې1��z��_ھX����GGظ�z�׌+���o�n��{G�=VF�@�	!��z
�0��=�����
8~ڷ��9�Q���x�c�]�N��3�ݽ�ϐ'�|ǐ��\ZX��44�%���7;����~��a��.����^!R�b�|��|@�Rv׬/��xP<<�f�"����C�oJ.[x����'RE׽�۰uw�0�q�n���a�/��A���xV�A�;����]�o�cP[��
.f{�����+�x�|3?����vi�E������"ND�/�֩�+��V�~x�Fڔ���6N�Gx�~g�z�����	��(5?ű���Nf�BV����}ִ�jgA��_1�qS^��#�\>]It��▦�� �*z����><Z�p��!�=c�,5��uG��3%�څx/:\]/�1����[���ɗ7�w5y}ܙ�.S�m�^�����u�(�pR\��@�E�`{��E�1�O�.�8�*s��˽$�}�����>#���(u����B�A�!�TCK��C7�B�^m^����H�����fn1�a�vt�"�Q��1�+�B��=�o|~�K���ag���-�`�:w�~C�A/��mnx���e�E;q\�:Fcc]�;���7��y봿p �����s��]D7����y�@�o��2K��Us��=��?�_��`��w���̀E�-J榃�p��qU��Sn�i���yuqV�wP%�T!�6�8]�?�K�w� ЮPz�+����;������Aui��<��<���Y��1�;w�Č>B�a[<��4���jF���EAr"�x���w<�Yw�NC��\^�{T�����a�}U{���{��?NZx�GE�d�Z|~�Z$��3/s�k�������N���#>(�q��0b�&`�����m���\���Ζ/��GZ��ю"�砊h�� �w��͑u�N�lS���^v��ْ�>s�KĜ^��_�˽�^������y?(1#ZdC��f�U���y�l�����݊�b���X����:��C-X�Xg����:�c��"�]u ��يfʘ�8$c��	���Ͼ��B�-,<rd���̶jkט5�,�h73�_ѯ��y��s�G<P�"�,�l
?m�x�i��4��L��<gvv��y4�A���v�)>PV1־��F�8�SX�r�7h"���|p�����"|���G~�G�^��n]�nk�:D$��B�tř��F���({*������Ck������LF�@��@g��>;.��SMr���c���.	�ˢ��w�@����y?c5�_������@�����\{PVͯ���5������ZA����Q�[�ef�n������y�M�>�u-a���-|S��?zi��Z��g��S��U]�z����,��X�^_Pz�O�`R���:���sS��V���[U��tugs�GE�a�b��V�i-CU`A|j�"��e)t$���93�|�[Kw��{FD��tS���7/ֶ��U��\SeP���B�/ޢE��~|h��ב7�ǻW*������PكU�`i<���u��~�=W��u�δy(������3>��S�U��>Vn���-����^����.�Z/�E���:kG��б<Yvǖ5�������a�e&!������{��Yu�G��g�����(�+6U!��K�}�b��~]/8j�����pc�?eD$�7
��g�_�WK|��B�=�X���U$سZ�G�j�b�XHg��=�iOfo�g�Ҿ����_a�����\F�#�.�8 ��!�)�T��W����^��ZC��/�[�~O��\~c�ĕ�CB���3�I\W,�'�g��-q�Y�u���֌��ĳ�;��|eM��q)�̾7���k&�{%iٌ3`r��?���}@��o�F_��]1���H�����Bo�U�޺��z���+��,�˦<��^A�!q[<Å�U��u�����̓�{��E���q!ִ�����v;�[7*�����Ѕ\X v��Kx~�O����Y��RTHܗ��M���Q~��J�a`�;�n�쭵t�q8���|o���vt��Ȇ��8�5�����6�ҥ����n��Uha��><��@aU�]�6�������4l���`g�̺�?*�v����8s�k���ri��[(��5}X�Z��s���_Yr]w��-o��g)ɮK�uC�+D\�4��be�gXC������{�V��_���+D�h�|�{���He峰��Q�o�VK5{5+2^��
��wI
�iK��<�Ȱ�S�CI|��5�������\w�|`~�x1��C���n�z��	Q.:�>Yם碻^�~g�9hqs����8�j��3�eN�Ԋ3=�y����F�×����?�>?�ҕ�#N�7�ή/=�ێ{=��y��{��	�����t��Ʊ��jK],*�sjCM���J���V{��}pe1���VÉ^n2T�M�jƥ��x� f���/���H�\Ofb�^��޾�ǈ�C-چ���ݨYQe����>FWy��t���?| 9��M'����1�d�X]0�+4��S� �����*����Ƥ7ZB��6��ydĂ��T{��߼殾��{�=���i��Ă�Ւ�gi�H)Щ~7q�T�z���awE=I�+
��+�`{���
�*C�a���߯��x��׾y������o)!ݰ:j�+%Ld����t}�L6¤�dĨq%gL*,�eN"�!���yg̘�L*���g�{��u9�&��Vjٌ.W�r�ۙa0�,c��N��P㓝K�V�0�w�*-GysdAG��i��ג���}R����DS/.w�j�6M��հM��}UǪ�$��s9��LE�� ����� [R��"26sy�˹B�:��:^��u����6��V��v0^�z��$���x�u��u�%<dV�W��,n���Bk��Y.BtD�p�6m�b�9�	ŷm��ZwES���v�a��m���(��|��P�Y{�����`i$��pe����5�'��{iJ�w�����D��f��K��Ǧ�2Y� �mʮġ�+*sU)WL��EGKᕔ�l�F�-W�:�oؔ��V�O�gO����uXo)�ӈ�[i�0#�q�tlV	�Ӧ��h���np��
ø�|�H�Zp�5zNK��.��v���q��Q�%���+n�������1C�#���uҤ������q�2��z�6zD�p�������3��Y�(`ucn���u�S��}J'y}L�Z�j`Rt�#,�+�<�i�`W8����kjj�t�̀�n/���k�4��n�9'շ�-����ٜ������3�­��{%9���u���OY��KG�={���4+�S(����Z��T]�B��W��̥�:)�kJ��9]��VIÃb�ygY�<��k I��r:o�X��Z��ciذ-,M��d����U�W�l�h��;3XU�m-�>�04@Zi��W57$�к ����p-��Z3n�7�)>:&�O�1����R��;�Q��cT�g)�a�[�[('��}����2�.q�R9���{�]��;�����}u��Y�퀉ơY*J�F!�Lf0���b'� c��cT�*ê�`T�9d��+ ƨ�a�V�Y*%��(em��eeJ��X���(�b���Ƣ��
)�eKj,[�fXV[V(�Z�QW)UQ�X\���,+
j�Cժ�@A�-BQ&5Er�a�E��A�A-�*J��RҐ��C�ʕ�VA�J�Ta�t�&��*
��V�eq��IF[AH�r�"1aQaX��i���R,QACM1ana(���"�H?|��?���ݪ]bܕI�ǧ���#�^�*�`v��!��I��^u�Iu���7�?D$>IPS��vi*He�h��O����<�H.�<���@�'Rvu���6�T�
AIĽ�����ν�<�{������;a����.Xz�i��4�P��H(
)�v�hVv�wd�Vi��+:d��a ��\�iU �l�>L�����۸v�Ơ}>�wHVf���Y�& (���M0�1ԩvJ����i ��=C
M%E�L*z�ޮ�0�S�<�^��ۧ[����g�m��T8���+'L�
/��5��!��B�ua��wL`v��
�dی�ݓ�Si�`{�ۿ~������{y��P�%q����*v�w�M$Mufr�2cP�Ă�S�
���gl1:@���Y���!х��W�g̕ �Cg�y���>�~��o�O�H)�
2zʐ}�j��V*�jɉ&�CX56ͰĂ���a���w�H(q�Y������;IS�
�x}��U�5׻����c%݇�`��
�!�y�AHd��%UH)�Y�ã��!Xm���I �2z����2T�f$���wd��r��������<����¤�!������
���i ����a�4 W�aXT�ME<@�w�A����R
L뇞�9�y�|��>����PR������|���'L6¤�� i*a�
,�eO7E&$0��-��cS�Y����{���g��|߿k�S�
Ì*t�{�|yM0�
�����^'�1������e@�T�R�*�
�1E&O(2��������A���sn}-��k��̶�خ��m�|s)u00��;�ƴeB4ľ�^�֦k����s��5)˷+-��dW;�n�ū+�-��^o����� ����z��A����~,�
yI���TP�%OP:�Af�.��0�f��Xs�A@����%UH;����Y������'���U緂"�$� Y*��X��l�6��ḏa�
��Rq
�QH�Ì*z͟Xi ��v��
�l<.a����[�����^o��T��'h��)�B���j�YY+���*)+'���$���N&�m�C��L@�T8β�E�������>����}�z�J�S�P3�<d�l�Ă��T����O*z�Y�옝�_l:Ն�t½�q1 ����E �>�`��T�}�G|�y����u���a곎$��<B�(���LO�����ă�Pۦ�H(z��Y���J���bAf�;�\�
ö�k����;�>ֹ'��
O���J���T�`x���;�*��ϓ�����P6�s�4�l���(i�ņ�VL��I�!�����o��~{�ٮ �ö>��I���C_Q@�;gg)������a@Qx��ɤ���� �@���a�� �`v�;7CH)��9�����\��}��]�=La�
��P1*��Y<�s&��RT�Gy���&'���$���36�S����������w�];ߞk���\��=a]0�()�_Y*)��H6ʇV��!̰���`i �5�ĜB�(�H=g�1��*A�&������9�<�5���|���T�Ϗ�1<IS�q�$z�ș�!XxºL��YY*q%UIP��`<� �HWÔ6ϓ���^Rb�O�>�	��8Ǳ/����N�'�7�[�W�c�D��r���uP�O3T�[��s�(	*ױ�}`��}C�VV&�鬩���)����<�w��~s|I;a�~?���yN0�,=aXw�$���T���:@��auE��ɬ���N&$������
�{~�|�>���z�Ϸ��{���'>��0�,�q �<k���m�$M��@�cP�Ă��S����Xbz�N�IY4f$l��N�秾{�����^��CI�)!O,6��$8����&�v�C�Xm g�v�<a�P6���;��;��<���N!R�
v�bbH9a��!���{LC�*Av���dR6�����l�1�d�R�݁��J�n�����������6ԃ��n�Vx��SFP1Ĩk�LH)�,Ă���JŇ�*i����*Aa�s(��*A��Ͼs���oϡ�j�g��_X}�H(%}`T�����T��I�+�����X��I ��'H(i%�&0�gZ�y��;��o94�P6����%H,P��6�JÌ*A�a�i��*A~`T��*t�S�:�$�'�n��1�u偉Oz��>��?g�{�<����`VN2�@�'���I��xϕH,;�$��L�8Ͱ� �'�4����C����$4��oT�﹟}���T9�7HV~�3�Ne���Ă�2Utn�Ĩ<�㤃�M٦gn�A@�TP����Ă����k~��>��n�=�V,4'�V|nɉ������x��0��@�Ht�����I&Ohc�Ldۉm �>@�?h����Y�`�:������'���G��I�0]JTr��E��m1sn�ǥm�qs�8�I--5���APՌ���$HOus�W�W�U��$��}=PY?	�qE!��öN�H)��w@�c�
�P3)�|��)�ْ|ʜE%g^Y1 �ϙ�n�L;aP=J�R����~�~ֺ�Ͻ�ϼ�J�bLN}I���Chf�
��;q�R
t�^�*(T�4�FN}f$���j�H)����+�QH)�z�ns3�u}�o^k�w���f$��20��V}�&!�J��T;C���H,�ꐨxu{a�t��Rw��Si+ժAO*i��t<ߺ��.y�_^��^s�u�,<f&2p��H(&��E ��X|�$��g,���bAI�+��@Qf'�14�Rk��L/�Y:5t�� �y�w�s�k~��u�@� ���OX}ݚHn�����4ÙOP*Aa������*m�n$7�a��z¤
��T�os��������L�eN�I_�`bAݚ�̓���:�$M@QM�W���I8�#�!Xm<��>0+[��^2TSG�N�(�|����zߜ�|VbA�!�Xx�T��fRx�f�l�@լ2����ߗ���`�:w���C6�����qx��@y(E��h;_x�A"񱳺窐[η��xz>?��?����ң��>u/���^�����ڏ�?7�jxD�z_؂!�u��3�.x�ݭz`;�VP��˿dV�\w���9w���0T��Cxኊ�/;��J4w�ڨ��
��bigO��(���ǋX޿�W�UU6����Y����Hq�A�9p=�iy}څ�L2���~����ρEǎ��l��y<`p<t�ڳ��u����eׯx��y<B%�!GO��/4Q�x�V��/����p���3{�cQ�%z�@R��+�=?�D8��<�����3�y?l�J4t�+$����ǈ�y���~������M.U.�r��B�S��Hv�� �g��t-�/	��r����r�J�i��"�&�r�!��[�~�Z'�G������W��S�z�
��ա��1��s��1�g�P��e[�}K�F���i��vw�骺�m@���!��B��86(���*:���B��e�������W���D��ӓ��!\�p�nm%��yV��3����tm"�ɹ�;.	.'#������v��wa�_���
��{�Ug��@���� e���g����{0\y��d�����~��-X�D��E�tŚ}����י˷�^#�f�"�W��I���N�3��6�7{�J�V����8|t�������?1����A��)D��y��|��8�P~B����;���x��[���UY~�M���O�1f�ĞU���	T��C�������bG�P�U�6GtǾJ���{>^�Ŧy,^P���l�"�pe]+\=(W��_Y �m�{q�և��}���P� 4��^��j��!e�$,AZ�lm�پn�>��&.?Qg�Z��z�W�z���Әr*RwQ�7i?Iy���p�b^�J����r�2ɘ��#�t;;�ٺ���f)yH�oe,��:hء�.=J(��6�U��p��?�着����=�I���"Z��q��V8X��X��dQZ��v������0��ZQGܾ����Ho��<B���p�g-���R3�~=����x���E&!��k# �x'R������
�k�+V����R�Y��R��X��zj>?*��{�ax���"�Jq��9�Y��a��lS�y~�OC؝�r]/��tVr��cW��T���}
�Ӷ��'�B'!��wˍn0�\F�#�r�ywl��g����I��A�r�F���;*f�DtǼwbl࿼h�Z����5|ǐ��\Zx���m�ڞ�W������p�1/���m�O�t���z�����'�v�"&��?Xs8�=��W/��]e� ��c��W�1�]W՚�q-�&c�ffFo]�|3!�DZ	�e��w�����w�s�o�O�>>�3�������?4Z��bޔk(z�sw7:U���z��|������k�!�������������A�*���	��SP��;��z��y�����?Y��竍Zg�Lo��C�z���%�s���Ұz�_�BZ���]{�μ�R����2qc{J��=W�Et���(ED���\tG�����{�s���߳}���ҍyx���c�Ye�~H��������"u{ٮ8�lLT���s�V-"��^��&h��o�Oy�_���R���m�||�(>���$'��S��E��{%��U���|<�� ��ObF��P�07�$<���V�lb�z��'6	n������Kv����OVL]�6�9���4o�x�0nZ�$�K8�;����m��]Μ�����WI�xغ�L�Wda��}�erÂ./��v��L~�n��=^�:��yF���+�/QZ�5����ؠ�S�uC��ez��1�Ŝ!����������|�/�ճ�;���Z��7�C��Ә�5Sq���$�ܰ�N+>�C�z*zح�?�1�ρ�P����B�"�������͍,
��j��l��y<`s+��OjzS�gӮ��0p������/����^z/ʈ����;�mI��¾��:IV�R��	>S�!Nl�'���:&��}�C�bgڂ��"a����f$6��}�NWWUv{�|���Y�0�Nǘ�@Q�v��n�,:�*�Bt�߇K����Ҧ_qte�����7I;��]&D�;D��V'����3t���$,VM����Kz+930�:�n��
��UW��[K�zf��W�D�6)Y�*���_=O�������<KR^��`�ڿ���W�+�b���t	
��8�{\�x��������P���-}b����~\p{}�=5�<�������5������Q�����g�B�Y�������<�V� ,�1��1�8��گO�/��Ƶ�ٷ�R��!��S�<CNO0������a<w�˺��J�Gޗ4F��-�]4ϩ3�?��#	�<���Wb���gv郼�_x���~8QTo킟��6z�@F���J����%'�Ü��CN�>}��I��+.���E;�a��H�x�A���_�-�ed���;��ߍ��Y������
u3z���ֶ�`��-v�K��O"���ˏ_�ɉ�il;".�&f������ɭe���^v���-,�ǋ��h�_o��-z�\������T�ۺ�/�����r������m�*�1K�j���c<1�Dsև!e����?j�DB(���c�K�p�m�̅�P�B\�s��hȍ���vY]���*��I���f��vd�K�\���k&�en3�N��U��4l��Um� ���N->�ۿ��2u��x ��/	���pUc#�_U���'9��-ɬVWc�ku�ogSf�AQ�7%����0�Y����Q*U;���JOl�"Ԭͣ��$h���s�5�K/"��֖�kb���E-<]VCӕ_��F�Y��n��u��I{�-�/�.B7��3�%d�׋[y?_���5�Y\�ư�0w<(��j!B�<`��c��|�&/���7NHNig\'3��,�;/�Z�gZ�'���` ���qF�j[t�yD͐E���qCP5�a�&�p��k)�����9��T������9�.2)E�ܽt�	m���b�h����Y3�,`�
J�N���\�v���0���r�M�,(tY9XJ����owg;���	�1�U)���(�N�ZǱ��:-Q���ڷ�rT�C�ϑݬm�l�sW���>�`��i@���	�_�N��T�x���dT�Zֵcf+[���fGz��&����@ȁt�XF�2����5�.�f]���&�8�b�ɋ�ܘL�SYB�6�PVi����z�pL��N9'.I�<s;qx��Ԯ$�����꘬V*����*5�(
��+PFI�J�U�V,QDE��T#P��� .R��J��PX���Q�1�X
�#X(E��	��"�QUt�Qc0����bŊ���#E�EH��*
��U,U���d�4�Tb "�
,X�($UR+0��Q�UdQE��
*A�E��Lk���Ȫ((�H��F"��U$�~$�A~���o.���n�۬�P�u^<!9(�${��t�ǝ�Jɢ�a��������o��>a�C��ǟ��1iQ����?t�C�2�Fz������QAUӹ�P�A�xA�]r��Z�l���y�K��i�)�/��/�T�a��n�!]u���6�M\\M�(a�OA<���C�T_׽��#�-Pr~�B4��{�(񄟡���o��y�6~����X��q���+6�k���/��R��5��s�)��t�y��|Jl�+7<:�^;Z*��tW�����^?1b|G�4�ۚH�ޖXդag!��'Oږ���՟+�${zy���K��>����Jջ<>>�VP^�S�`�̉^U2���s�B���z9�sXe�_T�����^/�y�G��*CW@�s�R��6rٓ:�;e<>8n�u "�ޖ�X��)�����W�D��^�K:RipT��_��諭����)^�������������V���?�YA��z[N�=Ymw�� ��T�l����!����i�$�|ifg����?{W�����+>?(y����8}�j�W_�|��y!oA��5 0΅�ď'�*�ʜ����B�������{���H�O�?Y�C��f�N�o���{X��*"G��y;������;Xz�K��T��>>��uy-�и:�T��L]��&)ډT:�F�9�8��}�y|��-3�ʦ6y��!�=좃o/{�!���(�GbJ�!%�X�yײ�R���	��sqX�?UN|��L�+!���!�y����7wgiT8�5p�p�gpU[ϭ�]a�pK��[�͛��d1=W�q-=���JB�/��E{�OS�C�P��,�U�g⪫���������}�6|�zQ�\X��01�,�>��1K�-8�d�,���ۣ���+7T;t��p����^�����~Ӝpy�!�a�r�#Մz��wV�!z���Gw��P�XC	i�`ht���N}�c�÷�e�R�{�Ձ��Y���hS����g��X��e@�����ρ��'��a�s�������)-����J�)k�{�P��0�~�ң��fӯ]nl��z��-��=a��:GV�/�_c6i��o��9Q,:F�"P�<�׳�)z{�l��t���@��
<0\v�+���<�̮;��~�W���T��^�q ƽ<��3W����x\�y�pWݵՂ,hv.�c���L��pz�N$� �\xa5r�7.j�m�i�$�;�����������TKk�������(Fbt��ǍRgq3����~΋�/����%Z��+���?ǮG��}w��i"�CڷS<~��j'A���Y���_5���Z�̫�ާ���-�\���9����ڢ��cO{�w��������q��Vs�=��+�CHccP���=�����Y�l3�����yYÆ�54@.z���z�}Y�{�{�3>(�=t��|��(���x���w�����������^x
#��wP��?/L�a�a=$�gc9}�:tߐ��0����ן�9�����3x�}？��X��NB�!�'0�5�@�ҽ�����ݽM�0��ٛ0���m�+�iL{�wvY�rn�z#z3�W^u(��u(SN �1gN��U�Z�1o^Z|�SW�����u���?��c�_�����o,"�i��;<���!�:���������0>�!T/���8KV�Tş
�tH��MW����P��� ꯽�N_q��|���D5휯]u�v x{x�c���, �0����;n_�WL���y�7
X���q�CK.�ů�g��gV7r���sO�9����{�p_!�8e*8�5շ��ʜ̳��J�z�d��¼��A��!V���+�㜵1������)y�ޝ�L^?Qg��n��Ey��wT���f�G0����z7��y�,Z��3 ��k�hYε0��b��!�7C�V�>�2���ˁ�o�Z��;][���&l�Mɰ�R��M�z�Qi[��i�J�.�G�t8�X����YՏd⑜B�G!`pS�F��I�.�h�"�,�XA��=�[��ꪪ���S��t�Xo���?TC��尠Ϗ��t>�C��v礦��M�p��"~cVl�L��p���^{����g�{n	��.�ϥϷ�a��K��"%�1�U��3Z�Z�P����WK���~��|�K�o�w��.~T��s}���XHe���~�R���߄��(h���}�-��/7�!�z��h�FZ�<����(�9��/�6��w��9:B?i�e�HG����#Vv��{�a���4<B���s�j@Y�QH�o܇�gU����할w�0�:��~?3ǁ�;��O����{ލׯuA^��FZ."Gj�pCG�@���.��(��m��;��샳���4�-Ezq�J[��s�za�L�o_�զ��,(��k϶Q�y���L8���I��(��.����J{���7�?ʪ�꯭%=�/��7w���15�py�)������AL}�xe�>��>�!���?/-4Q�dT`���n5�ek+n���	�C>b��g"�j�HM�<�x�J��nv�gx1Y� {�Ҟ��\;�%3��8u�ۼ�H>�+(�\�L�����3Nv�9rCy�fN��Kh�Wc+�� ��s����%8{���ҁX�x��d�:�̞�8@���9B��\7�`p�҆�w��}�0��A����"�BUk�w\m�K֚�͵��@`�Q_����uC�ׅ�G�p������r�5OAi��-"���J�先i[#�]���r��i����d5�'Z��nwM+�1���Hd����UUW�:'"b/��k�Dk����;�Z�D8,p�e�%�p��;-�i/fi��e+Q��O9^�
�5V�[6�T�m%��r��(�&{:Uxa�m^Џ]*!�@�XH\z-��ޝ8eg�z7�9���3�}RX�Ҩ�י�&J1�_����^BT�i�'��z�q�W��8�7/n�c��`1�c�IEҼ��c��+��t#��)���1�O��cu�ک��&��]�����T�rH�s� ��ŕ�49���R�L��+β0�U����[�E\ȯ/�E�v����޷���U�ޛ;��|�)�L�7�E��,g��4��u�{��U}Tu��������!�rm���w�e����E�ԙ�5���C^"sII#94Ŝ#�o6O�r��|C��wi���y�c�v��8�.,K?����a�ʷRr��zo���[�13���cZk'�x,[�c�I],j���޾���1=�s^�a��]\��"�Ā�܁�`����]y}�Se��^��}/*�>Iuv���7M��rf>��i*G�_�)6W>�>��-x��Y��Ҵr���T�� ��+t��*�H1�6}R��IoA��_��{��"������u�"��b�/�č�D�yyr���n|�K���#���pyMǊS��bƅ�o�ꪧ|�I0o��7�+w��M/ɥ�iU�W6Ɔ�wO_�TЃ{��u����7v��^�^�9��G6���_�^T���sX�>OS��VI{gX�ot�v�7Z����P�II�kދ�n	���0��xk�s�*�xל=�+��}o����}�����gIe�)�zF�\��tP�;ހ��s�Q	F/.��"���Q�������;ћ�h}~~9�_G��W��|�����r[���zu�c�_MoL��e��uݱ���z���vCWGfyƙ�Txɤ�
w[w�_ʖ
	qNjk32� �U�ƈnb�	�o�k6�`�W�y�;��*��{��)S��R_q���SO�chO����f�VB�CI�uz5r8�
�Z�'e�A�L5�Z�
�F�/,9�e�r�)�ݵ��^R�k�D~��:T�˫�����d�R�Vn7�&�-�IуD�h��e�޴J��cC����Q�1tje��h�v$��\�±��$pn���y҉o#R�1�d1�B���!Pƞ�v�v�3p��2��HCv��W7{gI��:�B)&��7��:v���gk�N���_nn���W�Nݲ�׫���r�c�)̈́�Η5��r�8i.���",���ۨ�Y��/I�5+�C���S�KFS�쬊�;u�wU��\@��SN��n�Cut3���r��OQ��X�WQ#E���[��t����@�[Ȍ׸�!(gt�W��<������qS�B8�	��f:�qP-ʫ�xkx
�hw[���^�xje]_n�hS|RڳR7awdXW_�2Դs���1�O�+���s:�&Ys�T�b�=��C��9�w�R��os��u�Y�L���LA8ot��&��r,y1�Ei�vE&�fGL�J��|�۫żW��m�e�놮N�Q�)T���A5�u�w�8<�6���7����CX�wQ���<t"��d��3r�Τjd{sHG���h���=��%�̔����a���=0Htw�w��y���j� ��*ޝ�g4����ґ���̝K��\%nf9�utr��	�QPU`����X��(�X��b�A�Q��AT�h��T�"�E�H�a[b*�+"�TV*z�Y�(�)�dulT"��+����+""�̶E��*�AAY1�(�UX,PE���`�R,�U�+DPR,QH�,1AE�̥dD�a]3��
c%�Q���b6�b�T�X(i�1O�H-"@$F�qn��ڬ�'�e�[!�ޜ�ް�R��� �6���+�c�� _��de�W�b�5��dT�[`z =��ɫ����D���ru�Qۇ�K�ߖ�~n�7"�{Fe���P!Ix^��W��~�B5MV��_%4E>��q���Y�ȼ��ĸ�U�)��Zp8|pd�+�Q�gg�����MxǫX�4YO/�F֘l^z��zدW�ɫ�D!t�V�Yі\�p�8L�����M�&��[̤����뗷�O��<�,^�G�T�+�bd����J��r'5no̞7�8�����:v��+��*�d�#�\�a3�)��f:ۮr���}ݳ.'K�3%��M%;�M����\�]��8�ʹ��}U��rNP/e~��ȊӤ#�7�V�kp6����j�A�՗��Y����O���H�m�;]^b�xE�Og9�9)�p����j7�C4��Suc��C�S�2H�rK�P{U�����jxW�rfW@p�n%�'�׆�45�S�n��P%�|tfis�t�ja�Xq���݆���ҖN�K�L�NG8k���7Q��Gۣ��<4�x��gB�kѻ�w�}�aO�iԪDS���v_h�ǤN�t�����ތ��.��0;T%�X���.�����y��(2�����Ѿ��|O�W�U�����%E�����dwU��C����R&t>�&�U��UF)�����HI#q]���j{.�\�jW=�޵��Z����Ȼw59�M�h�t����1j�joty��63�ڇ^,3g}�{3щ����[��O�K���	��S��z�=S;���\䎕���p��];Ǹ��3�����O���O�����f}q`��^��G>�Q���VVd��$�q��7=�'ګ�q$����;��կݐT9#���-C�3�oY��v}��S> 3E���{��^�6�Njc�n����$A�Dya�q��x�sw6���K��	r�����Ȳ���)�(ɶ��}�f�J{˄�U��'���"٬;�Oc�T��\֕���I�A%���3V0�xn��t3�ʝp��aI����?z:���f%W�J���z%�|�H�`}�nXyx�-�Ǉw���j��~Mu r��3�᚞T��7%���Y]�ɯ�^񬬃�"S��z��Y��j�ﴽצW`���"�9�2�t��Z����I�X�{�����~���&i���wR�7.e�}��2�κ�m�g�R����+��[~Yi��~��$�sN��җ5IVI��Ż�=���֬TS���:6��N ����h�qN��(�j\ژ,u��s?�����?N�p�)~ӄ>S{��O���F� ���_�/ߨ��~�\7�����Ư�/���Yߋ�����W���C��}t���y�l���as��u��{�:9_Ғi��O�b�U���i}��X{S�ӹ钴�?3�Ǆ�Q�PIoo��O	�d�1[�+)��j���n��P����x���(Q���`��Tr�|�:ˇh�����d��
���[�%�ڝ��x}&��ݘt�p	!�yİ_�[�g=���&��<�#:xÖ��w0���u�U�K.�gcrg��h���/�0���=�'���qSK!��!��(�E�U�߭$2+�k��#�Yy�ݨ����N;��:U�v�W B����W���~n߫�7XU�ᚎKy��Zo>IKk�SN��q]l�:�v����Wi�B�a��ʲ���C�F�Y��ͣS��Й���r��6"�\8w6�|���]���%���m�;�,��6{<��b乥OE���n��jѻh����K�x{�I�IV���:r��ڼ�ߍjC]My�b�L�q���wC]�Be�L���`�O	yq�-���g^��R%�wIk�I:fDL_�\�MҼ����U�������@ל�O	]��p�Ir;$�� ��?ϻ�NN��n��/�7ʷ�<�a鵱=M�)����i�Ռ6���p]]����t��q���fפ���Ľ�fE5I�@j�W����w�B��:k���v-ynd��SA�UӍ���A��jA�y2��⊯�Z����o'��j�Y�r-v6�|!����x��ףA��{�z�*Q᱘}��:�
�'����=r��k�<�v�K��ze�V�j`h�:oH����K�r��3[@�w����=���,cH�Ы��L�u��^n���J��S�q���Z��[�l�V�s<��:���F`��m�X�#��qA��*[=�����z�_ʤ�2'�p����P�ox���dDSo��s�>��u����.Ӹ�#�.�֥>b~�����=�Q�VǄ'#����G���^5��
@z����we0G�(���/oT	ڿ��U�Xz_
wyK{�<-T1y%ݧ�c���Y�Me)p
�J������{�'fj�9{�׾;��1΄���%kF��xW5��OzB�3�bͻ�j��~Mz�IOk�m�|%J�w<�<��f���s��������8�Q��j�`Ώ�w�S���9�|�q�{�o��QO�,i���Z��o���K5ZIKj���o9i����>���V�.��g�+W'#�^ūl̐��Y�*i䢭2�Y;kuZ�>����c����#�u���:�M����o|�#�ܹ|'L�@t���BeW%52w�2��=<��V}�XS�ӄ>Fq�*��7�B�SS@�����E��K������2/ڵ�;� 
;Y�/�E_!�j��~�����NC<���ګ�v��5R�Q�x$�`��L�Ӷ����I5��*󬗗�6gD��2�c��^�<�hMkI��hS��G�|-sUfv3�s7�fZ�M��6��4����琡+3��o�����ɹ.va��_"�ܣ�l�Io��V6���k�U�ʒOE�?�ɔje5� ֮��&�{�SKm���V�>��O�"����L}΄�.�\��?�gtܯdZBj�����R_�v�DT�;�Kٯw��׷���*T�����W�e;��e�.�gf5=�'z���l����h��}���zFs.`۵�x�k�D�n�V�{�=CT&-�,_]�y�#�]iw=�圕�v�:.D)�7�5�̨��Ӥ+E���/���'K�J>]VtE^9p�a���U�>Y���*BH��C?��������ơe��oDhi���if�GFł6���%�8%�������<�_N$�X �aLU��w\+���ۓNC0�Cz�[���A�9X�.r�2W!-+m�ԧh�S����k�9bi![!��:)4�<����y�w@�%����{�tV���R��`L`6����)��KIM�w&�h�msKy�m㦲�tUԣ�Z�]��2	3�=N��N������dgu�JF����7_Q�w9 �v��Ь�Afhp]�:Q�k�y��"I�%d8�����Y7@�(�o?<�#̻���l�sg���M������2{)n��)��<���,��k���73	���:�V����]3aj¾j��y��d��WM�0:�Q��a�p�kܺ&e�7]�#���!��vEL䬣X�I!�w�ͨ�ޝ؅L�E��M�1�hLI��.ҷ���ME=�v,��Fo�PAS�,r=���gh�Qv��Qܢ��L,��{�bH��l���{1��{���X�.7��n�.i��:V�����H��Lf���HE����J�̢m3� ٩k�u�ʯuok,!��ymB�9�[Ҷ�+�)��ͥ33�]���6�a��oosA�wB���@�Ǫn7�Mg*!c�6���r�ʗ�}2m	�_T�
�^]��:�U�gV��>���Xy��jV�\��)g�!��6���^����n�]�Z��))yf�,�\29�\�����V1��*�<]'q����EurAǢ���k�\�/�jt%<z�0c]#�wW,�)k���׾;�{;ћ�W��ATD��PPX*+Ɗ�*��F(���"�T���Eb�*+T�����b��*�DX��Eb�������*��Z��D-U���Q",�����Dv�"�1T�b* ���E���b*(�Qb��(�X�&����V1QU����
(�(�T����� ����`����U���?+Kx�_�?�)|�ͫunx�J�J�T�����\3���ѹ�g_�?Ei���7]��h���Yӯxe���Y�֥YoH�mi��uE�ޜb/�eP�t��i���x�~�d����;���.W�湔��i��
[���2����W��=�U��/�7hj��ũ��gR:۵�r�5�-������e�f�1������7��`�:<��dM�~Ŷk��$uά����eK�^�E�c]L���k1�ʅ��RT��u�U�~ܛ���o�+N`��"�/�1]����(�*$�]��f/�<M.�-��z�fD�|�C㶰��ݶ����	�jp��*s*����z�㝕nQ� ��&^��ܾ�/���ʒg��~�7�۽�k$��֮�*�H�$��R���Xn�a�:�ɵ�O��1y)�b{��J�\E��y7��陷���xL�}2�E(o������U��1t�M�5Lһ�*�� ��6.<�t`I����qwV�X��Q"�o�zN�:YQ��o^��JU��ī��*n5XkM�T2<z��O�6�$u�d�^W�E�Lt����f�g�b�GҪu��aj�K>�,!��wϼ�`�7�M����2ުb��{Pӧ8�T�{l�v��nB��1+�.3[���vVJ$6��W�ӊ��y��G��,_���{�+�~<e�f��K|��1�Jq3�V.o���'�%{��8��N�J߽�d����C�7�΅�6/&��w[�T����"d������xs��yu�>�k-]��n-�o.,��N�{� v�gڅX5�\ �R�7$����x�^��\�ӻ.{��Ε�Ն<�':��j^!E��F�ΓəT9�[��ng�1\�a˾���s������G��!�!8ǫI{��:�[�=���`��؟��3v��Ѿ�d>�%��S;���M�F ��>�p�+԰�R9yYw��v0[�eX
�v,��ᗍ̰���״��Μ�Zە�5D��S���y�Փ7���U~�7�ߧY������~3�wS�x�-YO�9��z��}�k�Jδx-C8U���g��X|� z�F	�Z�)�K�9�6�q��s^� tZ�/ϵ
�wRs�TJ��M�ρ�����ǷpW�?CbW���^�>N�a�ghGQ}Ӕ���xi�
�����<.�i�e/,�"I�q�+ԏ�8�U�-�Q͸q^���ʥfu��H.��VV��E�}�ӹ17/5��NR�
O����^
T{kQtQ��`�K���[S]B�u^��z�]D�v}�y��T�����a��9��r0���T��ٜ���r�\�*{cN��k�}�Jr?~�ۖ2��2��Y��Kx��u��߹����k��8�9l}���ze�{��fc�n�RƖ�Z]m��I�mXr��~�.-�(����6�U��ۅx\'c`�2T��'���㧨zr�-'Wx��3���8��qN�-5�)jM<����$=H[]����D����79.�:��b�b߱;�'���"�q���*RB��.�\wJ�ӽYe�."��uF��)��� �WCP��;ʹ��Nv���Io�n`B)�f��}P1�TԞ:%�����rͪJ�J4.�n��)B1�_nlN�t�R�lU�|�x��|����Z�}~Z�}�Ȥ1�/U��G��ڦ���6�73�3i��p�'�u{TmQU���f�d�,1���,�y���඗���o�as)�n��fi�y�(;`�V�KW'3ş � ���V6�B5y �.|��j�yg���qg.�)X�W|jͅ�r�`�wp��͈��2"�p68K	�bz��-�uΓnE�4������Zb��wD[6�bi��zۤ��wXf���d�G6����s��E52�bX'W�aZ�^�,ٲ��o:�d\[�����9��[2囬�L����H�F�l3�o�=��/3����H,s��P�o�'5��4���'�km���I��_�ғt���W?v^�Fi���6��J���D�W�5�ݕC�4����h<���麭^F�a#�z��i_��"(��u+7z<j7WE�%���pV>s�lV�C42��5�߼�Q��{�����=�,�b���y�O�d�g�K{w1i.�Π۳E��к76ڮ���֫��M>y��WN�]��7�3Y�́C����Uxɀ�t���-"/Yy�>F�kyF��5��.j��}W�oi�+�5�*����e��b�P�y�E���J�ǝ��].4�%j�V�N�ٲ�j����R	��8�2ظm���lt�u�J���q~���:?/�#�V������g����St�٥�/��+YT	��\��n�g����+o�>��K}�dUt���Q�Y6�ӰŅ�O)͔��}
�uy]�U��.��uw�Z������%�!�P;B�e�7çyW�L��U�quѸ�~����{ϡY��gQ���ç-\�Z5�2b���0�/�%x�3�Q�7U�=v���k��}��!��:n��H}#N�Ph��g38���M_8'/e�mey�<4�X�l��s��kݎ�-�|�|x�d�*a��0���:e�W�r������"rf�����!���Io���
[��t��<�/�UT����4�W�r�0q��^�H{u_��L�RCWR�z�h�*u�N7O{B�'�9br������H�K6��L�]�Y��H2J��R��uu�+�G�"V�XY7��VnIx�e���EZ�5�-�ٽ�i�Z>r7|����zeė�\)>;���&���
Z(��׎�m�_}��힏�~��mHVҏɕ{����u��d�p��nh�ȼ)UN&n�o���Lx��cZ�{dn���x�Z��RL��Ԇm���ZDfYUg����]
>��8�\�J�^��Q��u\mc�����a�s�(E�녙h�|75��LCVL]��9�7���_U������
�(ɒ�]X�R>C�Nxbo}u'�������&+O���F��Ҡ�hRG~���m�gs_>#;�~!Ϳr��#wK����MƆқ���<Y���S�U���9d�O)cd����u�U��q�GUW������j���y��OQp[V�_B��q�=ҹ�P���'���C��:�����L�.���մ6�����e����.I%.N7pB�Z����^��n�&�x��Q{�(Dkv�]��]a{>TS�Sd:!�ⷳz�n,�x8+��u�� :�d��������Ѹ�J�(��|K�a�[4��Ǖq"��wIڬ�6�� ��(B�n�3l���scΥ���n¹c�y�1�޼�Er���v�U�*-��+`)k�z��q�1qD�����4e�̇%(��&;-���qx��te*�Q����K-џl��%��)��m�ʨ�8F���M�4�t��g0c��@�v�KAB���v�dW4Kw�IY��JJ�71�K�&��	�%}bs�Q��]�xd��>Ԑ=].�E4�9���+M��sp�B�*�[�F$���O�<]K)�S�3�nݣ,�=��Bns��]���+�<�@7B``�#4*�GHʳ>P��`�t��*����r�Dr�|Ѱn2�r���,l����Joq�8��&�4+�C%���c��cuL���d�G!��L�T�uQ����f5�N�R�ε��'W(ðP�j��;O��Za��V�,U���X��բ��m�a�!�����9 ���^ӹxy(/2n�l��.�j��2��^X�Ȋ�6t ɳ��YW��Tw��H�[=O����gN{Mb6�umgMЂ!��르�:�^�%%�c����96����v�J�]�U���	ъqG2��kI��U�bGl��Uf)�5�Qm�^�v��W^t��.N���-ޮ3��KFqAHs�{�ꊮ�w����;Ee3�C�
۔����Z��F�ukDzX���F�Y���	J��!,*x�C��k�r��N�\�N+���]�]g�Qb�Ȋ�ƊȨ�TX"+QQ�+
�"EEr�"���)E�V"(
���Pb�ZJ�U��TUn�QEDZ�X*(��.�� ��h��*EQZʪ��`����""TE��(*��Im/V^�DUEQ��5h��V�PD+b�-J���)�QH���d\�D��"�9���߹�7���
��ta�u4Vh|�7<�A��ȐK��B��}�}O�����%��5��4�q�|�T�L2Ι�=�V���r����[8�/h��fP*���6D�S(���I�-�i�v��O@nV����Çs�b&��͎�By{M,��:����#<�Z���C>�+<cF��>���&�V�]Y#�5�|�wpǘň��P�Q`�J�y��ζ�#��c������^�!i�栤�F����]+�+b�w�T*9׷��s�,�J�:�fG���,�
j�ޛ�r��Z-	0S�cI�z�u+���讀\��z\T�_X�r�YMKa�I4G��W̩m#��
|R2e�}_}_R���<X�_�
`t��&��w���O]-��i3`��D��z���
;�˻3�����3�`��/@��Xt{�Ꙇ!�>I�z�u}Ҷ;9�WKPF��x��P(��duڥ��u�º.R�W^��k��
F�(s[���O6xsS�F0�����
g��k�M�=8C#��+����}�i+���WXbp���{�n�D��o�g;p}H��r��]P9�fZE���Ǖe9�G�ծ�t����~�F���֯ʱ�4e���n�-�21�(ft��yuc��R���)�-8�M7�x�*3-z��wd�rK̴3�ؑ�{S�4��1-����`�6}_UU2q����߫�ٹ�-:��5����d1E��D{BwO(��&�
y�p��p�ɯ%:
힧=h�YM\���׵�q2�������]�:/m'��nB�WD���*65l"�k�l��Vi����z�f�
m����:`}<��=��^�/b���OW&��6��G�����흳����/$u|�����˜ayrP��JY�.V��e���d�\���Wu�p�$�V͉m��0Q�;'v�+^�S0=�?+u͇��&x��{4�*jn����ӻyKS���n:!�[�⺹�PJj�\7��h�&�ŝn!��k��Ժ�3�g��ɂ�?�鑯OZ�_���%���.��nq�8���z�2K�\�����M[W�f��Ϋ�{̖�2fA�#0�8&{GI�Ӑ�hO���?[o�IG|��s'}!X�	/��n��Zr�hvg�ں��{$���롰��'��0yÛ�� ��t=�HeÍ )<��(Q�']M�L�_�F��!�]� �|��텊ʂ�1��T���u8���<]�NZ������*߂j�C��֫��ʌ.������=8^��=�6z�\d+��{7ո��Pg��;�3M�~�p��=���Fnd��i�sy̌I 	wL��Py�����I4O۝t-~�G��s��U�٣S�7 *�}Z��W�nEX�t@6�knL��Q^k#��V�B5{�7WZ����Dmz����Wz�g{�~��J Ɯ�疺S�g�e�.�u��]Z�䟯��Q�j���,�o����gEy�X���ׅ�3zϯN�y���h�s}!W[�l!L���u6eڗ��:x�ޕSF_�9�t�~�6�����;�x�e n5n��Z���T��izjOV9=�8�P�Y���n��[�t.��W	�Vq1QX��-O��{�t)v�@��ZFt�J����I�x���ͯ)�ٟ�m�zwjZ�ĩ�#��O�3���p��լ��/*�%b�(&Ug>����_����czC�W�1�[\]�T��ΐ��>������˜�^x���e���xjT�7��G���v��J���v����[��DR�W{T��x{7a�jf9���9􋼾�n���Â4���$�͓o�����D>������ېx��S��۔��e^����\��u�.�/��7-y�-m�s����4.�׹;���Ԟ���Z9D;�J���]�s�"Jئ]��xX'��P��HJĲ�g<��uٛ�xor�t%ш�v�ݻZ�-dL}�3�7{����9<W���D!���9~Ԍ�m\�WGx{޺ebp�7{�f��O-e�7	٥E���?[����7\�����$�ۈ\��Z'����L���D���z,V-9k�>�Z5�8���٦w9՗��չ��������c¦���+���~k��Ƙ~���<�rv���Ut�gh�[A�T4e�o/����8�oΣ������
z�kQ�w�U��+�j���ӫ��ؖ��^m�<���[3�<V^�T�cK*_W.�O�mc���[U���4g�����&ڀ�@�ە�Y�]�q�>���.��eYܽ�z�����~�7��[���3��*���'ْ��l&eH���zvB���Jr � ��n�e���d�*_(��Ӑ8YJ=���}����׽���C}��p�9vWd;��;�}4�3-r�%L�p�hwި��(�j�����jy���:��ͺDV��f���Ś���q3'�yP�кek�l5�����|q�.nQ�L�U{���k��R�Lƪd���=9ś��x�/�`<��zrm�{Y�&��N�=��g�
��^89�|s&$G#����ĉ�roW>3����r��2[��vK��/_-y���f��MŪI��z�`aY��'o��!��קbo5�����hb7IF�/v��G��5�6T���J��|R�'{y��I�=�:}�
^+��ej���c�Į�=�oâ���%�5Y+��>䛏{�όu����e�\�P�N��z)Eױ%����ׅvŇrN;�z<�J}�
.b���DR�ʡ���^��#JԐ��]u�zx�Z+7����v�n��}�s�9�gݱ�-��4���S-=�Zv���;OBM����ݩ^�2(��Q����#�pf%箐�u�/7Y�Ip�0�e��y����wu0&��m8Ya��Ž�]��$7�//�U�7{7�U�!n�3Vv]o��U�W�yrg����L֧�R���*�{����ҭ�B(#�	�DZ��lT#���2�s�;啦�=���sf"I9�����j~C+V}�f�%g�=�����[��S��i����Z���kz�F�z��+h���9{/Dj�ss�oN{"�N�|P�߯y
�,fE���ۼ[mM�z[�5n�x�ȅ@w�������ۆ���do΁�z��7�.���]Wwiq�0"f�܇(�V�6�3;�P3���XP^&a6���kT����բ�s���m�{��X
�B�Z��N�@sӄ6f��͞�)��w�ZH@��)Ғ�Į��w�}A�����*ь�=w���$�5�&���Q��:
ޕv���Tu}%0[�h�w?	^֌�=x�ɔjeU����X샧=ڷ���V5u����M�бh�U�����WS�vX �v�ȩ�c�RJ뻫mb=�*M�b�X֭`��ܛE\�e�d@���$Δ�n�V&�r�j2��X+l��Wn�J��u�$4u��,�Ĝ�u���b�s�8u�as�"q���z��2O\6{l8e{ywV��I��=^Ί=B�W�
����A���
"����̳*����h<�G5�S�Fv��z�Yn
��{��]?p�"W2�ہ��]+�ޫ��{�/\o��8�1�5���"ؠ��v��Cx��ʲ�F:W�v�Q^�E�!�/]����$�p���Y�6���"�XM�סM���wyT���#;m��t���q���jU���}!�����R�;3$��\�Ԛ�u��w� Kz"�첗<'��_u��m
��*�26�K]̎�����ǔ.H/�w�-�2�/��/yhv�,�xlo3
m��ތ��
!nԾ�G�\J|sf|몡qqw�bb�(�
�ZS��k�/��8���њ*o\`ۻ��}}�@�9٭K�I���U}6m%�7�*;�b`��ְo$3#x2t�	��}I7F�b�n*�b�MxR����R�`�u�}j��[F�I;��I�_D�[��\�rpٹ2+�$��"�]�:���h��TE���b�YE��TAPeac�Q��ň�EEV**"e�����EH�Ȫ,P�QR�e�D(�"�1QT!F(����e�0U���A\q2�D`��0SMEU������Vj���V-W-b�d��U�1r��F�����JV� �TR��X"���Vf���Y����1�Q�.W3+�%m�V�52�d�9E�Q�Z�c�7���3���s�OfmAkF���:���3�=R�ƶ�-y��ܥ�ϱR�G����̐�%#�|��l��j�P�XJ�cT4�9���w�s�^4sq�^+wQ��U�sQ;-�����v|�Gt�u�˞G�u���Έz,�ň��s�n���5��juy׆a�n�\�=����~�z�U�ػ{M։${�;���h����|tJ亟�*�ӣ��&oe�T[�q+F�}�1�[�S�&���l�[B���FF�<�i��I7�<�R�V{��{Y�0����SN��mT`Ԩ����tFk� ���_DB�u�&Y�Ӻ��r�TM�DqK�Q4����
5�+jJ5��%G]>�����b�Q|�E+.^y5V��?H�j�Ev�%�`z�'����%;z�*.�I�W/-)�.ox��^�QS��4���
�w���<�جG.�*�Z��v���)�j�D޲�9A{k�d;��S*�1#�w�4@�t.g	R��sۯ1�0<ߤU|����D����|��}��{춫7a�ev��VޖܤT�n��i���a���g��0�s�̝����p68M2�I|bvK�����лu�et[�Վ�\ً���%��g�=עdZ��:�剄��(�}��m3}y�X�O2��{����.I���4����ͤK9f�+����H�dk]�qC#)�N��w�<"oDX�YUϥ���y��<��*�Y7���;��z��
�����,��c�^����y��?n���O��U���`�Vv~�y<�֒�vj��w�[}T9�� g��,D�4�ygHզMZ�����h6���f9g1�=����,�U���5ҿ!E(u}՘L\L�FU��~�"�VV�=�G��;#�' �Ht�>�$�mV��i��M%d��Ӵ��]�ϗG�Ypx*���ɦ�R	R�|5�f�vB6ז�+��xj���A��\�r���޳�6E�[3�L�R%�)K��1%rAӴa*��P����7�)�Ń���*Zo���ؚEv[�ҽ�Vgǆ�g"�6�j>8>���~N�7�
(���X\����닷��ώ��8g8#{�9���^<��¹��Q���LڍÃ]�0y��˝qM6CƎ�x��]�:+��W���8�=��v��޹P��v�E� �����8���9���
sQ�[V��F�{8�t΋d��eX�ɤ#Uˮ[�ƪN��6FDK:B_��������jcAnJ�]%��x��Q�ͣmYIG�ܗ�v��AK���m�ۛ^֧��3� F�ܤ��i��t�볔V>�q����73sM\�ګ�`�>k��#��C6�ò�~+�^|i�5<������K��&<h(�AT��j�k��>��Љ�q̮S����i�r�pDX̝I� ���)�d��j�WK�R4]Uڊ����7f�)�W���sܘG���`���)9��oobdU�]��Q!`̮ިC�a�9p9mF������n`ѷ�u ^n�J>2�9]��7&��Z}�X{���*^s�xɡaK���h5�/�D�V�*�滇^�%ӗe{�Y�qBE�S�mi������^���2���to�����xa^�j1o;�u���tl�g?�/��~��׶8�����v�ǖ��MB�J�2���������L������=�x�5z�v����l�,C�l}�K~F�0��U�������({�,�-�uc�����c�Q�p:�������'i���rN。��M+�W���[t}7�+mB�RtѢ+�t���{��<V`�:������y����
��|t�H"K��J˲^�0�]Z_�4뮚z��S���1�<�qѯ]s�,��M��X�=�������*��@}�m������5��d����&��En4 ������3\����l�hf����/��Y�^��d&D�Q�)�
kyo�d�xͳ�H�=��H1�F#�j����mV������idvx�-��Ϯ��[� ���g��^L��|l��V�K�q]�g;'���{�V�Þ[�s+�$��ܫ��nPJ��dK|�Z�ޫ��2�u�Jo���h�L���ɼ�R�ԯ ���_���K�}[uk�fx�x^�}�����1鮬����6j)�멽z���-�n�Y=W-C�0��J��u4}za�į��a�+T~n��,���A�%��3��w/m2qu�hsyu�^����F]ܘ�V�)�����32�!Z�89B
�{�s�9�r��8�5�s.o=�ǜizN��W�le5=��_��ޘ}���hp� �߰V�Z�Tk|�T���[}е���jTݵ_���>�?��o���i�weW�5s��	��Z�����^���Q33�Muu�z�B���k�G9��6�U��x�͙*ĬϜY����[��b��}VW��^���$�0���O|Wo�.�/b�zyf��\��`EU�[���z(���T��:���Wۑd~ϏE�\�S����U�^�e]i3p�f��H�����DZ�Ϛ��{��=��ե�6^�oΤuFk���U�l�z^�ҁh�)�*t�W�梛;�r����[8}�Zֳ��㲥ɻ������9������2��崸�u�6+4��K<ә��@
�%��j�.�v�Z�=Q��>�K��aQVG�g��7�}5���}��t�f�F*N^8H�>�4b4����������L�*il`��.^qX�D�d^IԠnRt��4X{s���-��}{�%~�J���R�~�-�!P�=>�*�]���;�b�����sܘ�G¥��gr���͎�wk��_��EZY���y�Ytݼ�^#.���$Yռ�^q,�_^���s\�qW���0�Q��Q'����͹�ι��%y��ɬs��;~/#�#v0֬� SE���#�y�"�"��ǆ�VPܞ쎙��՝I�b���-��M��n�B2�k��O"pu��S�me�=ͬ��.��_vTB��zx��p}uh�$��3��7��V&�ɭ���+���{R���{?=����ɕ��8��W<��y5�}ĩ/%yP�!)���5Yy�F���L	�����F����/��ށ�ZB��
�p�'d�0��ug{r���@�L���U/���/fy��r��Kj�����������Jъ\۱כ��7��aWy��"=�)e�w*p�M�����W�	�5C����K�� �4q{ʏnO9��kaYy<kÒ7c�&EPaƭ�x�[:�	܈UӮSe��j@�#�Y-Xx5��Z���
�q-���Yj_jlȮ��I�MnUw�5u:2�w2�<I��0�\��nVNVce^�9Z�Y\,M�zDJ����u���E-](����TGlZk�=ȅ�;����4Cڝ�6G Qj�^��������Yͥ2�7z ��s/E(��<��a)���0�I���8uԡ�8+{m�����m�A��w�����#�Z�[]�h���5s��$�� j#�R�SZߥ��;��}�:m��5���!H��VN�3����=�C����(ܗ�n������ͬ�N�)�K�E��V1��C95��u����-k��J꟔�k�VN
�rRl�Ji�j>��:�����;gE<�{Lx����E���%�i��<�ٓ,:�#�g.o3P�;���c$��5v3�-+��{'VeBs�f�ܐ�+̪+�e�B֮�
�k A�@_sW����9��T��j���;�ٺc��CPL��c��ID��^B��v�b�N�.껌aEf��Q��6�'>����nVj�� ��F��Bʒ���C��2��i*�8��r���xЩ���UZ��,�qgۿk�l�Wk��)X�	(( 3K�W3/����h-���!�����hj�N���K�zƮ-#���e]����'n�������"=-��^���fJ�*e[���h���&9�3P�7�������l9��'���M=*���E�ܳ�Fd���
wuwK��DmK� �-E�TaiAV,���TPm�Eb5��2ɂ
��Q�aECUAA`�T�C0�iP�,Z�V�c�Q��amF��ADm�V�2�,�iVdPR�e5�c(��PQkF����d-
E�E�D�����4�Le��	R4h�*2V
�k4�
E4�դF�E*���z۱~t�r��	J�N��'Aߎrt��t�s��c�.�[no#-N�Ҽ1�Ok�Cҝ<�M<���W&�G=~�t�;���ui~�]��/"W�8�+�3'�ł�>�j�ɵ�:_l�o���)׵;u��L�L�S�N4�)���$�@�f��.�>�7夲ᗝE�7���n�[���x}��+6���~y��7�u�b���m�u���w=�{�zv�H���ΞЮ�Dk)>�yp*Ŵ�8oU�*����=�����b�$�2�w>��h�B�Ad�}ئϖ{�mzUλF,8	L��.��23��uy�D���L'��^�Z��2�û( Ht�*YG^���H�G�}���r���{j)޳]Hg���u�d`�<=$J����3W]Y�5ۧ���{Iܞ2�Iu���gT�xۡ���_��&��S��U��>}v�UҌ��n���)���F�a�~�j��]/@�ذ�%�sz�F�z}ּ*5�|B=;;�.�it��"Q���ؗn��ؼg��=���<+��mW8p'�{��Tw�*^��-��d�Դ��g�5��<�A+����E�縱�b�1�Z��>�zM2�ђ]���K.m��õh��에���Œ������rk�� Q_:�28"�1T�1�8J�[x(�#�8��I4�W�z �Y��N'��{��ǖQP��I-���sţ�\�&�e�=���t�Ew9��2{@ʆ����IYc5��s�y�%�S��G��{�eu���9=�ͳܹS^��������)$v�lS�e/C����ծ������7��׌��r�����ƚ52R�����H��O�Ø5�ڈ����x�ƶ���8��y^�խK�����Jl��;�2K�%��<�I� �pտ��¢���,����Y�[#�T�5��|L��,�l���|f�G��K����"�FT��f=�	�=�$du��*R:�,��	�r��V�q�c}:D��ڲ��]*��ЌR����oTɲ��Jf`����luʽ�?��U��9��`���{T�`8낭���]{w�Z
���M���.{X��"������𰱖��{�'����̊6=�s�W����U�gHJ�T�y��
�pu�	���K}#N�x�8(�dһ��[��E�ڊ~Ώ�{�#��~-һ�2.˥���XgƢ�p�[X�/[�ڙ9�O`w��tM���B���[�F\4�+z�D��}n������v��W����^PYY��uYe4;���nqy毲�[~ƚ]��a�ÄVҙ6��	R^n��c[Qb��(4N�}�xg�G�}��5�p{��-�ZB�F�P����ߪ0z��������>p,�����j�I=�N�O7��;K	L�R�*�r7�CT�o��
>6;��<zd�jPAPȢ��t�O5�+٢���s���������ꥡ�V��b���U��k�z�fu�-�T�V��D�U���_ӎ��i��<P`ܯjv�j�˛�gw	/�J3�T>x
���TX�/�\�ѲɉL��Y�7���l�VKԞx�Ѩ=����Y��T��IZ��`<X����y���aLe,%�FԲ9�:����+�[�,ˑ�/�%Km�yG� �ᇛ4�R'n? r���4�Ǩ��~[��*3!��)R߷(.��?v�4}Cd��։^gv���W~+͛��kV����+>���/���琫�d�dI+�}&���^�Y�g��g��=�l�R�t�M���^��jK����c�]Y�n!Sܦ$[�H+|���-�otjҰ���V�_9�%��I��5��)��IE��;�����z��sC�0�1�_A���gq�����Ԟ*=�
#*��/F@Ԧ�G�՜|҆�i�5�K
R�Y�4�h8X��2�l��o�RY3)�8f5��f-Y0"c�{-���)��-0#����n\��̧/z���ʊ���>:���wuƻ��7	�e�4��W������M�2���ˑ���59�ݏcʩ;�+2���)��6�w��Y���qZ�i�]c�4��Υ�������*�2�;�,����7�ؗZ��˘Y�Uκ�'����_aٯI���R\�5��<�X"�s;�`���A�;!No�[�w���c��Pӽ���L��������
+5'��D[u=��.���G�m].�%���s�pO޷�w���UvFC�0l��BI�>������9[���8f���(������]��6F^����y��ǽ!�ܗ16�-M�ػ�/���X�<�����V����D�;������)UE�5����f�c�΃Xl��I}�O;J�UԞ��[��5�!Eʝ=�ו��}�k�~�*��w�N��P����Ќ|���K�M�NhJ�N"�J�J�ujX�2�wRS�qq\h:��^[R�\w��Z�Ʌ���RY=,ߘ1k畋�"��Ǵ�{(�$���mxnyl�������>�<r����g��r�w3)0V�λ�<���Ѯ�4W��Oعq���Slhm���Jϭ�`��,r��>���M�-`�=Y�V>����`DE��殆MD��3iYs�s��m�$8���>M��WlG���jW�o�C���W���l�Xmt��.�r�9N~���=�66����&~^2w��E���?��x�5���Y�j�[}��zaNp�1Sc�O;�C�z���c`��j�)Йh����=Y�43~�.��+�y����/��X ���T�ƺ��s�=Y>�z��hƮm��n�&W�px�[��<g��S�7q�Z��+���B��В�Oh	�:��yd�^�<�޾S�ҟ��b}Hv�l�X���Sk��������Πq-��yظ��L�#X�u3��9�KR�xW��'�](��Q��(���r�0�u�w�v4C
�<���&W�8IS����,R�����)�y.麔����
7� boWWj^(����-�Ceg�����/Tv�+U�L��j��,�3��5��]��I�V����+H�!�~�� �9�V�۫'D��Q�%Ԇ����X�Y�3�g���Ĕ��[�M��~>����S*�f?}|��.>O�d�a��y�ѥ��a��n�"��s����i;������U����~��$D`~�[Y��וTE��7����Y��f�&Y<8�J�@wA��#E��x�u���a�F�nC1���xNJ��jt��!�՛:+QjL��ޘ[�j�z�<��w|���z-��4e������b��s�4�j;�j$"SOy9�W�4�s��*�r��]�#����u��"��<����X�O��CV�J�P{���s
��V�z�.���Mv�FM�N���M�x�����7S����v!{g'em҈�"�"v�k�Ovm+�Dv���,�Эa2Nf���� k珒�Yґ�xy|k���#�w6��1�éX�mg0%���T�	�)�������;�i7Y H"'vYF����"x%�6-��t3���U���J�1_
�tN���P���K0�j��tA�ee���q"I�}:��6���z��哋�jWc��cK��j1������[aL;Gj�%_'�v�'���H�6�]☶e���Xr���i�T#�c6Hѥٽaf�^�ies�L*1ô�a
N�/GWz�,�c:�u�|��y���.���c���a8a�6��fƤ2��#yִo����n��1��G[��wd��:�8��[��}���]���lh���ĸbQj�	��j����ar�������5�3N�t�4N7u�-��r
�@�Sb$��h�ɕ��ڨU#4^��2�7.6�Ž,�rQ��DKj3Ɔ7�)��p��2,�5���49�fk�T��%��8^_v�|{e���]f7nm㒂D�ó\�1��,�8n��\����'#b<����M�JX�Hݚܻ\�Υ�>�aR��H,�AIRVQ
�sTҦ���8�X��AI�E�1���	[�0d"�IY5iIe����1��VTY0RE�`bLʡI�M0��J�Ek
��%I+
��AB�%I�J�J��IFLdӎ2k(QP�1	1RV�\�eC-VV+ �k2����������4���y7ң�����]M�G
T�0����K���À���!�Pc��Kxۮ�)p���y���^�>�[5��3��������	�0�S�ș�}P���m���,��v���,N�ey4�%�^���׾s���͗�8�^JTV��v��q��>播��27o� �ܒ��_�K�iW+�*magd,t�S/-�U���&����WwǓ�bqm[��~5y�������$cp�:�+WG�{� 9�X�V8�1�⨜����ԙ��5ܼ@�r���j�b������'�Հ����ʕ̲Y�c85Z���@������}�*��>n�C{{��qK�T �4{���(D��U�a����x,��/s�ߡ��#^6�ɱ=rf\����)ģ�w+�\�u�On��E�޺°���kѨ���DcQ/^N��ì#����5�����n��J��@�:�Ť.g�<�r-��9{x�8�5��!����u���"����|«��	�:*
f�������ֹ3T��Jl�P)\`���z���.ʝ���a��@�zk���Y��g4�=���i�&GJ�?�(�=�Qz�;2��-8\�'�V��7y˱�y���=C�<�^u����E�&���ze���Ss�fJs<��)U��:T'Z�K,G%tI^iI2��6[53=:�-��{�ۂ0�&s����+��_!V&E�yް�7�R�2`I�PJ�׆�v�v��KB�Ҍ��rҲ���O��y]b��2��VN�Pu����݌��R�{}������
��+�ƍx�}�եF�'!_�}Ր��꿋=3�Z��c��kQ؟s��������#ЛmL�Eڒ�QL)��5O+8=�ry��b(���]�-�j=>�κ�3�@�F�o��^�J��ާ��`fY�.�1�<����h-C*
r��XK�3���*��{XlD�i�����ˮ-�p�2C�.�dx�����{ vZ��I]޷�E�td��=D�⬶f"����F�f�4=M�$��4����i�{Aܝ)����(�ү{\���^?F�B��w�J��a3�T��mQ�Z�V9{q��@2�$��[�j������o�1V'���{r^�j���ֺ�B��[����u30m��m�ߌ���1�O��=�k��֗R�������.�q�N*뫏=fD��mI��z`J��ӞW��YT*k���;7�P9}5�V��~,��`^��3���7c"�]�ٷ��wûLZ�
���W�$�RዚF󚷐��%�®�S�i{��E��_u`�M!柼���:��d�+��9�G�A�?�fl�6LwYe��#�y�K3��}喤1�o�}z���n'g�5xǴ���?T�WK��
G$w���g����撄����^�0uh�B��ug-o"�OE[n3;�)�5���{O��P�؝~��Mˢ��ҥ�+lF�{4����p��3}&�j���ͻ�D 8��3�%S�-i<�u=�<��үZ�>q�0��3�~������n�K��cC!�;����ǡ]������5go+ɉ��d�n�Q��sc|����IJJH��Y�q�S�Jo<�z�͝$��߫�M��{����G&�`��佶�YR�'[L#:<�>���Z��~5rv�tpIIޝJ"�Խ�:�;W�p	:�v6�n/)�TT���c{���˘[�.˜ʲd���N[�n|2�������e����u�a�˾�o�i�������@i�ܢ1�G�R��?m���8�a��6�N۷��-}�n��ZW]O<�	�c�ې��w�eS��ŧ�]�쇲���('�Q�x�\� kka���~v��ׇ;�f��6�u�+5�����޼��Uƹ�%�9[C�2e��	ޡ��"����R��� چiDT�ӌ�c�e��$r&)�W�G�E�wq�7B��j[�rI.}��TvƵ�n��w��Ir.�z���ȟ�P ���kr�T�эS^l�#�^��R�o�r�����rc�������H/z���wU�)��N��w��Zc1bT��5=��ѕ������Z�j�����x�������a&y
q����!���Y�y�G�R$�9�]W�Vl9G��&Vu��Gl<Y�P�m�l�';܂ٜ��Pъa8N��O���	�ו0�0�XEz�՜��{c�5��v��]o)o�!�ި6��O80��Ë�rP�7��vq7��'/
�C��a�Y�Nkq�N8�孓��4E�,�s�54^�+yq�8������(%D4��041�L3�_(��_�c�w�~��~����k�6F��dec�I��A
��逿{�o�>��\g���5���N�z�F�4�)+��Cּ9��xWh;[���>�kH����=0�pyq��#�7������ݝ����f_W�O�"��
��<�#�w��aÔ9e�{����|@���!�|t7Hq��ЙOnd�/��[�4_�;[r�|+�.Hq�@*<0yq�D�V����o�M^���0x�:I�+�~���ٟ;�|%�O���T���9�m[��@���5�az�l[R��I�B�Ѱ�z��={�s#�x�0�c���_i�5]�۴��|��S�S!J�웥v��N�gLU	�F����9(�k�_�m5���e����{1�Ɔ��%���qN*m�Kfq����J�U�̊��hqq�>���Wl�OS��o -ߌO���;g���vd�O��"Z!_@j��g�d�u[G@�'��VG���|�f��0��o��3י��"Sp�u{�A!�W~�)�G�L8��([ ��4����o��J}���i��l�K萄Z��@g��;TE]�I�'�5
� �)���7f}�NeV?����<kƸU�+;��6���|�������7Kbkbry���t�����{�͞$�di��`���n�\)��l�$vC�ļ��Q1o���|p���.6Q��[�����e�|<�Q1|��H'�a�a���Ӵ>�&ｵ���6�D����ι��>��%ܥ�ڙt�K\���:����� Ω���c/�G�m]W*Ǔ�����v�����Ip=̼F-d�S���L<{Πc����=z��g����y�\����i�q�Bp�z��bX�pD�[W�1�U��3��������ψk���.� Q��:�;���W��7������<n�墇�~z�T�RL�̄��Q�C<��Ꞃ��ƭQb���㑜ڻ������#�~�+Xb,���x��j����|�y��:�r���z�������b�r_׎�zĬ$������'և�8t�����8~���3���Y�J�}��q��}k܃��0�\C�(�c�4�+�)���}��g���&M�k�d�ڼ�IZXH�,�HU�q����?]+UQUrB�?��@����%��	! ��{�/�3+��S:���0�F{�O[4���H��	I$��B�hXr��48�~�M��wC����!$ f���Ń�~�T���Kh�:��*�Sd�#jay%o���ի<�+�-�4C#�a���xk͐����Nw�����<� ��~�HI�&�!$ ���XE�����s:#��b
%�JC=��_����?��?g���
~��	! ������?��t ����!ْ����'R>���+&��A�UI�s�.�|F�v��v�(o�	?���@	!�	 @��}<a���������!  �tl*�o�S��0.g����i�?�������읤/�;���g��������dY��Xg�F���K�̧xs� ����}B���,I����~��a����?�?w�����룅q@�o��ත������8 ��Is+������!$ ;���w	C��}�����=��'�w""�I! �p~p!$ �t�D�O_ܓ�hY?V��Ŀ����B�����;��B���8�1�0P�?�zO��@ �2ud��@?Q��a��ٲ']V����r���'}����0���GZ����?�tBB��?a��g ?\?`����	�����z�G�2��؏�Z6%!�-3����K3���\�}��u3D�vd{��v$�������O��a� BH@?l���u���a�O�'���?�='�N�&|��h;C�#�l�zhb!���_���w ��lXa_00��i��Z
����{� BH@m4$�����ՠ�vs��k�3��PD9z��_��c�Ԓ������2$$���,� a�� ~����<���BBH@?l���������?o��:�{'�N��?}�D�����q@7��Gg���H�
|��